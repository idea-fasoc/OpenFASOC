* NGSPICE file created from diff_pair_sample_0474.ext - technology: sky130A

.subckt diff_pair_sample_0474 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=2.19615 pd=13.64 as=5.1909 ps=27.4 w=13.31 l=1.16
X1 VTAIL.t4 VP.t0 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=5.1909 pd=27.4 as=2.19615 ps=13.64 w=13.31 l=1.16
X2 VDD1.t2 VP.t1 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.19615 pd=13.64 as=5.1909 ps=27.4 w=13.31 l=1.16
X3 VTAIL.t2 VN.t1 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=5.1909 pd=27.4 as=2.19615 ps=13.64 w=13.31 l=1.16
X4 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=5.1909 pd=27.4 as=0 ps=0 w=13.31 l=1.16
X5 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=5.1909 pd=27.4 as=0 ps=0 w=13.31 l=1.16
X6 VTAIL.t6 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=5.1909 pd=27.4 as=2.19615 ps=13.64 w=13.31 l=1.16
X7 VDD2.t1 VN.t2 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.19615 pd=13.64 as=5.1909 ps=27.4 w=13.31 l=1.16
X8 VTAIL.t1 VN.t3 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.1909 pd=27.4 as=2.19615 ps=13.64 w=13.31 l=1.16
X9 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=5.1909 pd=27.4 as=0 ps=0 w=13.31 l=1.16
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.1909 pd=27.4 as=0 ps=0 w=13.31 l=1.16
X11 VDD1.t0 VP.t3 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.19615 pd=13.64 as=5.1909 ps=27.4 w=13.31 l=1.16
R0 VN.n0 VN.t3 312.007
R1 VN.n1 VN.t2 312.007
R2 VN.n0 VN.t0 311.791
R3 VN.n1 VN.t1 311.791
R4 VN VN.n1 61.8135
R5 VN VN.n0 18.7188
R6 VTAIL.n570 VTAIL.n504 214.453
R7 VTAIL.n66 VTAIL.n0 214.453
R8 VTAIL.n138 VTAIL.n72 214.453
R9 VTAIL.n210 VTAIL.n144 214.453
R10 VTAIL.n498 VTAIL.n432 214.453
R11 VTAIL.n426 VTAIL.n360 214.453
R12 VTAIL.n354 VTAIL.n288 214.453
R13 VTAIL.n282 VTAIL.n216 214.453
R14 VTAIL.n529 VTAIL.n528 185
R15 VTAIL.n531 VTAIL.n530 185
R16 VTAIL.n524 VTAIL.n523 185
R17 VTAIL.n537 VTAIL.n536 185
R18 VTAIL.n539 VTAIL.n538 185
R19 VTAIL.n520 VTAIL.n519 185
R20 VTAIL.n545 VTAIL.n544 185
R21 VTAIL.n547 VTAIL.n546 185
R22 VTAIL.n516 VTAIL.n515 185
R23 VTAIL.n553 VTAIL.n552 185
R24 VTAIL.n555 VTAIL.n554 185
R25 VTAIL.n512 VTAIL.n511 185
R26 VTAIL.n561 VTAIL.n560 185
R27 VTAIL.n563 VTAIL.n562 185
R28 VTAIL.n508 VTAIL.n507 185
R29 VTAIL.n569 VTAIL.n568 185
R30 VTAIL.n571 VTAIL.n570 185
R31 VTAIL.n25 VTAIL.n24 185
R32 VTAIL.n27 VTAIL.n26 185
R33 VTAIL.n20 VTAIL.n19 185
R34 VTAIL.n33 VTAIL.n32 185
R35 VTAIL.n35 VTAIL.n34 185
R36 VTAIL.n16 VTAIL.n15 185
R37 VTAIL.n41 VTAIL.n40 185
R38 VTAIL.n43 VTAIL.n42 185
R39 VTAIL.n12 VTAIL.n11 185
R40 VTAIL.n49 VTAIL.n48 185
R41 VTAIL.n51 VTAIL.n50 185
R42 VTAIL.n8 VTAIL.n7 185
R43 VTAIL.n57 VTAIL.n56 185
R44 VTAIL.n59 VTAIL.n58 185
R45 VTAIL.n4 VTAIL.n3 185
R46 VTAIL.n65 VTAIL.n64 185
R47 VTAIL.n67 VTAIL.n66 185
R48 VTAIL.n97 VTAIL.n96 185
R49 VTAIL.n99 VTAIL.n98 185
R50 VTAIL.n92 VTAIL.n91 185
R51 VTAIL.n105 VTAIL.n104 185
R52 VTAIL.n107 VTAIL.n106 185
R53 VTAIL.n88 VTAIL.n87 185
R54 VTAIL.n113 VTAIL.n112 185
R55 VTAIL.n115 VTAIL.n114 185
R56 VTAIL.n84 VTAIL.n83 185
R57 VTAIL.n121 VTAIL.n120 185
R58 VTAIL.n123 VTAIL.n122 185
R59 VTAIL.n80 VTAIL.n79 185
R60 VTAIL.n129 VTAIL.n128 185
R61 VTAIL.n131 VTAIL.n130 185
R62 VTAIL.n76 VTAIL.n75 185
R63 VTAIL.n137 VTAIL.n136 185
R64 VTAIL.n139 VTAIL.n138 185
R65 VTAIL.n169 VTAIL.n168 185
R66 VTAIL.n171 VTAIL.n170 185
R67 VTAIL.n164 VTAIL.n163 185
R68 VTAIL.n177 VTAIL.n176 185
R69 VTAIL.n179 VTAIL.n178 185
R70 VTAIL.n160 VTAIL.n159 185
R71 VTAIL.n185 VTAIL.n184 185
R72 VTAIL.n187 VTAIL.n186 185
R73 VTAIL.n156 VTAIL.n155 185
R74 VTAIL.n193 VTAIL.n192 185
R75 VTAIL.n195 VTAIL.n194 185
R76 VTAIL.n152 VTAIL.n151 185
R77 VTAIL.n201 VTAIL.n200 185
R78 VTAIL.n203 VTAIL.n202 185
R79 VTAIL.n148 VTAIL.n147 185
R80 VTAIL.n209 VTAIL.n208 185
R81 VTAIL.n211 VTAIL.n210 185
R82 VTAIL.n499 VTAIL.n498 185
R83 VTAIL.n497 VTAIL.n496 185
R84 VTAIL.n436 VTAIL.n435 185
R85 VTAIL.n491 VTAIL.n490 185
R86 VTAIL.n489 VTAIL.n488 185
R87 VTAIL.n440 VTAIL.n439 185
R88 VTAIL.n483 VTAIL.n482 185
R89 VTAIL.n481 VTAIL.n480 185
R90 VTAIL.n444 VTAIL.n443 185
R91 VTAIL.n475 VTAIL.n474 185
R92 VTAIL.n473 VTAIL.n472 185
R93 VTAIL.n448 VTAIL.n447 185
R94 VTAIL.n467 VTAIL.n466 185
R95 VTAIL.n465 VTAIL.n464 185
R96 VTAIL.n452 VTAIL.n451 185
R97 VTAIL.n459 VTAIL.n458 185
R98 VTAIL.n457 VTAIL.n456 185
R99 VTAIL.n427 VTAIL.n426 185
R100 VTAIL.n425 VTAIL.n424 185
R101 VTAIL.n364 VTAIL.n363 185
R102 VTAIL.n419 VTAIL.n418 185
R103 VTAIL.n417 VTAIL.n416 185
R104 VTAIL.n368 VTAIL.n367 185
R105 VTAIL.n411 VTAIL.n410 185
R106 VTAIL.n409 VTAIL.n408 185
R107 VTAIL.n372 VTAIL.n371 185
R108 VTAIL.n403 VTAIL.n402 185
R109 VTAIL.n401 VTAIL.n400 185
R110 VTAIL.n376 VTAIL.n375 185
R111 VTAIL.n395 VTAIL.n394 185
R112 VTAIL.n393 VTAIL.n392 185
R113 VTAIL.n380 VTAIL.n379 185
R114 VTAIL.n387 VTAIL.n386 185
R115 VTAIL.n385 VTAIL.n384 185
R116 VTAIL.n355 VTAIL.n354 185
R117 VTAIL.n353 VTAIL.n352 185
R118 VTAIL.n292 VTAIL.n291 185
R119 VTAIL.n347 VTAIL.n346 185
R120 VTAIL.n345 VTAIL.n344 185
R121 VTAIL.n296 VTAIL.n295 185
R122 VTAIL.n339 VTAIL.n338 185
R123 VTAIL.n337 VTAIL.n336 185
R124 VTAIL.n300 VTAIL.n299 185
R125 VTAIL.n331 VTAIL.n330 185
R126 VTAIL.n329 VTAIL.n328 185
R127 VTAIL.n304 VTAIL.n303 185
R128 VTAIL.n323 VTAIL.n322 185
R129 VTAIL.n321 VTAIL.n320 185
R130 VTAIL.n308 VTAIL.n307 185
R131 VTAIL.n315 VTAIL.n314 185
R132 VTAIL.n313 VTAIL.n312 185
R133 VTAIL.n283 VTAIL.n282 185
R134 VTAIL.n281 VTAIL.n280 185
R135 VTAIL.n220 VTAIL.n219 185
R136 VTAIL.n275 VTAIL.n274 185
R137 VTAIL.n273 VTAIL.n272 185
R138 VTAIL.n224 VTAIL.n223 185
R139 VTAIL.n267 VTAIL.n266 185
R140 VTAIL.n265 VTAIL.n264 185
R141 VTAIL.n228 VTAIL.n227 185
R142 VTAIL.n259 VTAIL.n258 185
R143 VTAIL.n257 VTAIL.n256 185
R144 VTAIL.n232 VTAIL.n231 185
R145 VTAIL.n251 VTAIL.n250 185
R146 VTAIL.n249 VTAIL.n248 185
R147 VTAIL.n236 VTAIL.n235 185
R148 VTAIL.n243 VTAIL.n242 185
R149 VTAIL.n241 VTAIL.n240 185
R150 VTAIL.n527 VTAIL.t0 147.659
R151 VTAIL.n23 VTAIL.t1 147.659
R152 VTAIL.n95 VTAIL.t5 147.659
R153 VTAIL.n167 VTAIL.t4 147.659
R154 VTAIL.n455 VTAIL.t7 147.659
R155 VTAIL.n383 VTAIL.t6 147.659
R156 VTAIL.n311 VTAIL.t3 147.659
R157 VTAIL.n239 VTAIL.t2 147.659
R158 VTAIL.n530 VTAIL.n529 104.615
R159 VTAIL.n530 VTAIL.n523 104.615
R160 VTAIL.n537 VTAIL.n523 104.615
R161 VTAIL.n538 VTAIL.n537 104.615
R162 VTAIL.n538 VTAIL.n519 104.615
R163 VTAIL.n545 VTAIL.n519 104.615
R164 VTAIL.n546 VTAIL.n545 104.615
R165 VTAIL.n546 VTAIL.n515 104.615
R166 VTAIL.n553 VTAIL.n515 104.615
R167 VTAIL.n554 VTAIL.n553 104.615
R168 VTAIL.n554 VTAIL.n511 104.615
R169 VTAIL.n561 VTAIL.n511 104.615
R170 VTAIL.n562 VTAIL.n561 104.615
R171 VTAIL.n562 VTAIL.n507 104.615
R172 VTAIL.n569 VTAIL.n507 104.615
R173 VTAIL.n570 VTAIL.n569 104.615
R174 VTAIL.n26 VTAIL.n25 104.615
R175 VTAIL.n26 VTAIL.n19 104.615
R176 VTAIL.n33 VTAIL.n19 104.615
R177 VTAIL.n34 VTAIL.n33 104.615
R178 VTAIL.n34 VTAIL.n15 104.615
R179 VTAIL.n41 VTAIL.n15 104.615
R180 VTAIL.n42 VTAIL.n41 104.615
R181 VTAIL.n42 VTAIL.n11 104.615
R182 VTAIL.n49 VTAIL.n11 104.615
R183 VTAIL.n50 VTAIL.n49 104.615
R184 VTAIL.n50 VTAIL.n7 104.615
R185 VTAIL.n57 VTAIL.n7 104.615
R186 VTAIL.n58 VTAIL.n57 104.615
R187 VTAIL.n58 VTAIL.n3 104.615
R188 VTAIL.n65 VTAIL.n3 104.615
R189 VTAIL.n66 VTAIL.n65 104.615
R190 VTAIL.n98 VTAIL.n97 104.615
R191 VTAIL.n98 VTAIL.n91 104.615
R192 VTAIL.n105 VTAIL.n91 104.615
R193 VTAIL.n106 VTAIL.n105 104.615
R194 VTAIL.n106 VTAIL.n87 104.615
R195 VTAIL.n113 VTAIL.n87 104.615
R196 VTAIL.n114 VTAIL.n113 104.615
R197 VTAIL.n114 VTAIL.n83 104.615
R198 VTAIL.n121 VTAIL.n83 104.615
R199 VTAIL.n122 VTAIL.n121 104.615
R200 VTAIL.n122 VTAIL.n79 104.615
R201 VTAIL.n129 VTAIL.n79 104.615
R202 VTAIL.n130 VTAIL.n129 104.615
R203 VTAIL.n130 VTAIL.n75 104.615
R204 VTAIL.n137 VTAIL.n75 104.615
R205 VTAIL.n138 VTAIL.n137 104.615
R206 VTAIL.n170 VTAIL.n169 104.615
R207 VTAIL.n170 VTAIL.n163 104.615
R208 VTAIL.n177 VTAIL.n163 104.615
R209 VTAIL.n178 VTAIL.n177 104.615
R210 VTAIL.n178 VTAIL.n159 104.615
R211 VTAIL.n185 VTAIL.n159 104.615
R212 VTAIL.n186 VTAIL.n185 104.615
R213 VTAIL.n186 VTAIL.n155 104.615
R214 VTAIL.n193 VTAIL.n155 104.615
R215 VTAIL.n194 VTAIL.n193 104.615
R216 VTAIL.n194 VTAIL.n151 104.615
R217 VTAIL.n201 VTAIL.n151 104.615
R218 VTAIL.n202 VTAIL.n201 104.615
R219 VTAIL.n202 VTAIL.n147 104.615
R220 VTAIL.n209 VTAIL.n147 104.615
R221 VTAIL.n210 VTAIL.n209 104.615
R222 VTAIL.n498 VTAIL.n497 104.615
R223 VTAIL.n497 VTAIL.n435 104.615
R224 VTAIL.n490 VTAIL.n435 104.615
R225 VTAIL.n490 VTAIL.n489 104.615
R226 VTAIL.n489 VTAIL.n439 104.615
R227 VTAIL.n482 VTAIL.n439 104.615
R228 VTAIL.n482 VTAIL.n481 104.615
R229 VTAIL.n481 VTAIL.n443 104.615
R230 VTAIL.n474 VTAIL.n443 104.615
R231 VTAIL.n474 VTAIL.n473 104.615
R232 VTAIL.n473 VTAIL.n447 104.615
R233 VTAIL.n466 VTAIL.n447 104.615
R234 VTAIL.n466 VTAIL.n465 104.615
R235 VTAIL.n465 VTAIL.n451 104.615
R236 VTAIL.n458 VTAIL.n451 104.615
R237 VTAIL.n458 VTAIL.n457 104.615
R238 VTAIL.n426 VTAIL.n425 104.615
R239 VTAIL.n425 VTAIL.n363 104.615
R240 VTAIL.n418 VTAIL.n363 104.615
R241 VTAIL.n418 VTAIL.n417 104.615
R242 VTAIL.n417 VTAIL.n367 104.615
R243 VTAIL.n410 VTAIL.n367 104.615
R244 VTAIL.n410 VTAIL.n409 104.615
R245 VTAIL.n409 VTAIL.n371 104.615
R246 VTAIL.n402 VTAIL.n371 104.615
R247 VTAIL.n402 VTAIL.n401 104.615
R248 VTAIL.n401 VTAIL.n375 104.615
R249 VTAIL.n394 VTAIL.n375 104.615
R250 VTAIL.n394 VTAIL.n393 104.615
R251 VTAIL.n393 VTAIL.n379 104.615
R252 VTAIL.n386 VTAIL.n379 104.615
R253 VTAIL.n386 VTAIL.n385 104.615
R254 VTAIL.n354 VTAIL.n353 104.615
R255 VTAIL.n353 VTAIL.n291 104.615
R256 VTAIL.n346 VTAIL.n291 104.615
R257 VTAIL.n346 VTAIL.n345 104.615
R258 VTAIL.n345 VTAIL.n295 104.615
R259 VTAIL.n338 VTAIL.n295 104.615
R260 VTAIL.n338 VTAIL.n337 104.615
R261 VTAIL.n337 VTAIL.n299 104.615
R262 VTAIL.n330 VTAIL.n299 104.615
R263 VTAIL.n330 VTAIL.n329 104.615
R264 VTAIL.n329 VTAIL.n303 104.615
R265 VTAIL.n322 VTAIL.n303 104.615
R266 VTAIL.n322 VTAIL.n321 104.615
R267 VTAIL.n321 VTAIL.n307 104.615
R268 VTAIL.n314 VTAIL.n307 104.615
R269 VTAIL.n314 VTAIL.n313 104.615
R270 VTAIL.n282 VTAIL.n281 104.615
R271 VTAIL.n281 VTAIL.n219 104.615
R272 VTAIL.n274 VTAIL.n219 104.615
R273 VTAIL.n274 VTAIL.n273 104.615
R274 VTAIL.n273 VTAIL.n223 104.615
R275 VTAIL.n266 VTAIL.n223 104.615
R276 VTAIL.n266 VTAIL.n265 104.615
R277 VTAIL.n265 VTAIL.n227 104.615
R278 VTAIL.n258 VTAIL.n227 104.615
R279 VTAIL.n258 VTAIL.n257 104.615
R280 VTAIL.n257 VTAIL.n231 104.615
R281 VTAIL.n250 VTAIL.n231 104.615
R282 VTAIL.n250 VTAIL.n249 104.615
R283 VTAIL.n249 VTAIL.n235 104.615
R284 VTAIL.n242 VTAIL.n235 104.615
R285 VTAIL.n242 VTAIL.n241 104.615
R286 VTAIL.n529 VTAIL.t0 52.3082
R287 VTAIL.n25 VTAIL.t1 52.3082
R288 VTAIL.n97 VTAIL.t5 52.3082
R289 VTAIL.n169 VTAIL.t4 52.3082
R290 VTAIL.n457 VTAIL.t7 52.3082
R291 VTAIL.n385 VTAIL.t6 52.3082
R292 VTAIL.n313 VTAIL.t3 52.3082
R293 VTAIL.n241 VTAIL.t2 52.3082
R294 VTAIL.n575 VTAIL.n574 34.3187
R295 VTAIL.n71 VTAIL.n70 34.3187
R296 VTAIL.n143 VTAIL.n142 34.3187
R297 VTAIL.n215 VTAIL.n214 34.3187
R298 VTAIL.n503 VTAIL.n502 34.3187
R299 VTAIL.n431 VTAIL.n430 34.3187
R300 VTAIL.n359 VTAIL.n358 34.3187
R301 VTAIL.n287 VTAIL.n286 34.3187
R302 VTAIL.n575 VTAIL.n503 25.1255
R303 VTAIL.n287 VTAIL.n215 25.1255
R304 VTAIL.n528 VTAIL.n527 15.6677
R305 VTAIL.n24 VTAIL.n23 15.6677
R306 VTAIL.n96 VTAIL.n95 15.6677
R307 VTAIL.n168 VTAIL.n167 15.6677
R308 VTAIL.n456 VTAIL.n455 15.6677
R309 VTAIL.n384 VTAIL.n383 15.6677
R310 VTAIL.n312 VTAIL.n311 15.6677
R311 VTAIL.n240 VTAIL.n239 15.6677
R312 VTAIL.n531 VTAIL.n526 12.8005
R313 VTAIL.n572 VTAIL.n571 12.8005
R314 VTAIL.n27 VTAIL.n22 12.8005
R315 VTAIL.n68 VTAIL.n67 12.8005
R316 VTAIL.n99 VTAIL.n94 12.8005
R317 VTAIL.n140 VTAIL.n139 12.8005
R318 VTAIL.n171 VTAIL.n166 12.8005
R319 VTAIL.n212 VTAIL.n211 12.8005
R320 VTAIL.n500 VTAIL.n499 12.8005
R321 VTAIL.n459 VTAIL.n454 12.8005
R322 VTAIL.n428 VTAIL.n427 12.8005
R323 VTAIL.n387 VTAIL.n382 12.8005
R324 VTAIL.n356 VTAIL.n355 12.8005
R325 VTAIL.n315 VTAIL.n310 12.8005
R326 VTAIL.n284 VTAIL.n283 12.8005
R327 VTAIL.n243 VTAIL.n238 12.8005
R328 VTAIL.n532 VTAIL.n524 12.0247
R329 VTAIL.n568 VTAIL.n506 12.0247
R330 VTAIL.n28 VTAIL.n20 12.0247
R331 VTAIL.n64 VTAIL.n2 12.0247
R332 VTAIL.n100 VTAIL.n92 12.0247
R333 VTAIL.n136 VTAIL.n74 12.0247
R334 VTAIL.n172 VTAIL.n164 12.0247
R335 VTAIL.n208 VTAIL.n146 12.0247
R336 VTAIL.n496 VTAIL.n434 12.0247
R337 VTAIL.n460 VTAIL.n452 12.0247
R338 VTAIL.n424 VTAIL.n362 12.0247
R339 VTAIL.n388 VTAIL.n380 12.0247
R340 VTAIL.n352 VTAIL.n290 12.0247
R341 VTAIL.n316 VTAIL.n308 12.0247
R342 VTAIL.n280 VTAIL.n218 12.0247
R343 VTAIL.n244 VTAIL.n236 12.0247
R344 VTAIL.n536 VTAIL.n535 11.249
R345 VTAIL.n567 VTAIL.n508 11.249
R346 VTAIL.n32 VTAIL.n31 11.249
R347 VTAIL.n63 VTAIL.n4 11.249
R348 VTAIL.n104 VTAIL.n103 11.249
R349 VTAIL.n135 VTAIL.n76 11.249
R350 VTAIL.n176 VTAIL.n175 11.249
R351 VTAIL.n207 VTAIL.n148 11.249
R352 VTAIL.n495 VTAIL.n436 11.249
R353 VTAIL.n464 VTAIL.n463 11.249
R354 VTAIL.n423 VTAIL.n364 11.249
R355 VTAIL.n392 VTAIL.n391 11.249
R356 VTAIL.n351 VTAIL.n292 11.249
R357 VTAIL.n320 VTAIL.n319 11.249
R358 VTAIL.n279 VTAIL.n220 11.249
R359 VTAIL.n248 VTAIL.n247 11.249
R360 VTAIL.n539 VTAIL.n522 10.4732
R361 VTAIL.n564 VTAIL.n563 10.4732
R362 VTAIL.n35 VTAIL.n18 10.4732
R363 VTAIL.n60 VTAIL.n59 10.4732
R364 VTAIL.n107 VTAIL.n90 10.4732
R365 VTAIL.n132 VTAIL.n131 10.4732
R366 VTAIL.n179 VTAIL.n162 10.4732
R367 VTAIL.n204 VTAIL.n203 10.4732
R368 VTAIL.n492 VTAIL.n491 10.4732
R369 VTAIL.n467 VTAIL.n450 10.4732
R370 VTAIL.n420 VTAIL.n419 10.4732
R371 VTAIL.n395 VTAIL.n378 10.4732
R372 VTAIL.n348 VTAIL.n347 10.4732
R373 VTAIL.n323 VTAIL.n306 10.4732
R374 VTAIL.n276 VTAIL.n275 10.4732
R375 VTAIL.n251 VTAIL.n234 10.4732
R376 VTAIL.n540 VTAIL.n520 9.69747
R377 VTAIL.n560 VTAIL.n510 9.69747
R378 VTAIL.n36 VTAIL.n16 9.69747
R379 VTAIL.n56 VTAIL.n6 9.69747
R380 VTAIL.n108 VTAIL.n88 9.69747
R381 VTAIL.n128 VTAIL.n78 9.69747
R382 VTAIL.n180 VTAIL.n160 9.69747
R383 VTAIL.n200 VTAIL.n150 9.69747
R384 VTAIL.n488 VTAIL.n438 9.69747
R385 VTAIL.n468 VTAIL.n448 9.69747
R386 VTAIL.n416 VTAIL.n366 9.69747
R387 VTAIL.n396 VTAIL.n376 9.69747
R388 VTAIL.n344 VTAIL.n294 9.69747
R389 VTAIL.n324 VTAIL.n304 9.69747
R390 VTAIL.n272 VTAIL.n222 9.69747
R391 VTAIL.n252 VTAIL.n232 9.69747
R392 VTAIL.n574 VTAIL.n573 9.45567
R393 VTAIL.n70 VTAIL.n69 9.45567
R394 VTAIL.n142 VTAIL.n141 9.45567
R395 VTAIL.n214 VTAIL.n213 9.45567
R396 VTAIL.n502 VTAIL.n501 9.45567
R397 VTAIL.n430 VTAIL.n429 9.45567
R398 VTAIL.n358 VTAIL.n357 9.45567
R399 VTAIL.n286 VTAIL.n285 9.45567
R400 VTAIL.n549 VTAIL.n548 9.3005
R401 VTAIL.n518 VTAIL.n517 9.3005
R402 VTAIL.n543 VTAIL.n542 9.3005
R403 VTAIL.n541 VTAIL.n540 9.3005
R404 VTAIL.n522 VTAIL.n521 9.3005
R405 VTAIL.n535 VTAIL.n534 9.3005
R406 VTAIL.n533 VTAIL.n532 9.3005
R407 VTAIL.n526 VTAIL.n525 9.3005
R408 VTAIL.n551 VTAIL.n550 9.3005
R409 VTAIL.n514 VTAIL.n513 9.3005
R410 VTAIL.n557 VTAIL.n556 9.3005
R411 VTAIL.n559 VTAIL.n558 9.3005
R412 VTAIL.n510 VTAIL.n509 9.3005
R413 VTAIL.n565 VTAIL.n564 9.3005
R414 VTAIL.n567 VTAIL.n566 9.3005
R415 VTAIL.n506 VTAIL.n505 9.3005
R416 VTAIL.n573 VTAIL.n572 9.3005
R417 VTAIL.n45 VTAIL.n44 9.3005
R418 VTAIL.n14 VTAIL.n13 9.3005
R419 VTAIL.n39 VTAIL.n38 9.3005
R420 VTAIL.n37 VTAIL.n36 9.3005
R421 VTAIL.n18 VTAIL.n17 9.3005
R422 VTAIL.n31 VTAIL.n30 9.3005
R423 VTAIL.n29 VTAIL.n28 9.3005
R424 VTAIL.n22 VTAIL.n21 9.3005
R425 VTAIL.n47 VTAIL.n46 9.3005
R426 VTAIL.n10 VTAIL.n9 9.3005
R427 VTAIL.n53 VTAIL.n52 9.3005
R428 VTAIL.n55 VTAIL.n54 9.3005
R429 VTAIL.n6 VTAIL.n5 9.3005
R430 VTAIL.n61 VTAIL.n60 9.3005
R431 VTAIL.n63 VTAIL.n62 9.3005
R432 VTAIL.n2 VTAIL.n1 9.3005
R433 VTAIL.n69 VTAIL.n68 9.3005
R434 VTAIL.n117 VTAIL.n116 9.3005
R435 VTAIL.n86 VTAIL.n85 9.3005
R436 VTAIL.n111 VTAIL.n110 9.3005
R437 VTAIL.n109 VTAIL.n108 9.3005
R438 VTAIL.n90 VTAIL.n89 9.3005
R439 VTAIL.n103 VTAIL.n102 9.3005
R440 VTAIL.n101 VTAIL.n100 9.3005
R441 VTAIL.n94 VTAIL.n93 9.3005
R442 VTAIL.n119 VTAIL.n118 9.3005
R443 VTAIL.n82 VTAIL.n81 9.3005
R444 VTAIL.n125 VTAIL.n124 9.3005
R445 VTAIL.n127 VTAIL.n126 9.3005
R446 VTAIL.n78 VTAIL.n77 9.3005
R447 VTAIL.n133 VTAIL.n132 9.3005
R448 VTAIL.n135 VTAIL.n134 9.3005
R449 VTAIL.n74 VTAIL.n73 9.3005
R450 VTAIL.n141 VTAIL.n140 9.3005
R451 VTAIL.n189 VTAIL.n188 9.3005
R452 VTAIL.n158 VTAIL.n157 9.3005
R453 VTAIL.n183 VTAIL.n182 9.3005
R454 VTAIL.n181 VTAIL.n180 9.3005
R455 VTAIL.n162 VTAIL.n161 9.3005
R456 VTAIL.n175 VTAIL.n174 9.3005
R457 VTAIL.n173 VTAIL.n172 9.3005
R458 VTAIL.n166 VTAIL.n165 9.3005
R459 VTAIL.n191 VTAIL.n190 9.3005
R460 VTAIL.n154 VTAIL.n153 9.3005
R461 VTAIL.n197 VTAIL.n196 9.3005
R462 VTAIL.n199 VTAIL.n198 9.3005
R463 VTAIL.n150 VTAIL.n149 9.3005
R464 VTAIL.n205 VTAIL.n204 9.3005
R465 VTAIL.n207 VTAIL.n206 9.3005
R466 VTAIL.n146 VTAIL.n145 9.3005
R467 VTAIL.n213 VTAIL.n212 9.3005
R468 VTAIL.n442 VTAIL.n441 9.3005
R469 VTAIL.n485 VTAIL.n484 9.3005
R470 VTAIL.n487 VTAIL.n486 9.3005
R471 VTAIL.n438 VTAIL.n437 9.3005
R472 VTAIL.n493 VTAIL.n492 9.3005
R473 VTAIL.n495 VTAIL.n494 9.3005
R474 VTAIL.n434 VTAIL.n433 9.3005
R475 VTAIL.n501 VTAIL.n500 9.3005
R476 VTAIL.n479 VTAIL.n478 9.3005
R477 VTAIL.n477 VTAIL.n476 9.3005
R478 VTAIL.n446 VTAIL.n445 9.3005
R479 VTAIL.n471 VTAIL.n470 9.3005
R480 VTAIL.n469 VTAIL.n468 9.3005
R481 VTAIL.n450 VTAIL.n449 9.3005
R482 VTAIL.n463 VTAIL.n462 9.3005
R483 VTAIL.n461 VTAIL.n460 9.3005
R484 VTAIL.n454 VTAIL.n453 9.3005
R485 VTAIL.n370 VTAIL.n369 9.3005
R486 VTAIL.n413 VTAIL.n412 9.3005
R487 VTAIL.n415 VTAIL.n414 9.3005
R488 VTAIL.n366 VTAIL.n365 9.3005
R489 VTAIL.n421 VTAIL.n420 9.3005
R490 VTAIL.n423 VTAIL.n422 9.3005
R491 VTAIL.n362 VTAIL.n361 9.3005
R492 VTAIL.n429 VTAIL.n428 9.3005
R493 VTAIL.n407 VTAIL.n406 9.3005
R494 VTAIL.n405 VTAIL.n404 9.3005
R495 VTAIL.n374 VTAIL.n373 9.3005
R496 VTAIL.n399 VTAIL.n398 9.3005
R497 VTAIL.n397 VTAIL.n396 9.3005
R498 VTAIL.n378 VTAIL.n377 9.3005
R499 VTAIL.n391 VTAIL.n390 9.3005
R500 VTAIL.n389 VTAIL.n388 9.3005
R501 VTAIL.n382 VTAIL.n381 9.3005
R502 VTAIL.n298 VTAIL.n297 9.3005
R503 VTAIL.n341 VTAIL.n340 9.3005
R504 VTAIL.n343 VTAIL.n342 9.3005
R505 VTAIL.n294 VTAIL.n293 9.3005
R506 VTAIL.n349 VTAIL.n348 9.3005
R507 VTAIL.n351 VTAIL.n350 9.3005
R508 VTAIL.n290 VTAIL.n289 9.3005
R509 VTAIL.n357 VTAIL.n356 9.3005
R510 VTAIL.n335 VTAIL.n334 9.3005
R511 VTAIL.n333 VTAIL.n332 9.3005
R512 VTAIL.n302 VTAIL.n301 9.3005
R513 VTAIL.n327 VTAIL.n326 9.3005
R514 VTAIL.n325 VTAIL.n324 9.3005
R515 VTAIL.n306 VTAIL.n305 9.3005
R516 VTAIL.n319 VTAIL.n318 9.3005
R517 VTAIL.n317 VTAIL.n316 9.3005
R518 VTAIL.n310 VTAIL.n309 9.3005
R519 VTAIL.n226 VTAIL.n225 9.3005
R520 VTAIL.n269 VTAIL.n268 9.3005
R521 VTAIL.n271 VTAIL.n270 9.3005
R522 VTAIL.n222 VTAIL.n221 9.3005
R523 VTAIL.n277 VTAIL.n276 9.3005
R524 VTAIL.n279 VTAIL.n278 9.3005
R525 VTAIL.n218 VTAIL.n217 9.3005
R526 VTAIL.n285 VTAIL.n284 9.3005
R527 VTAIL.n263 VTAIL.n262 9.3005
R528 VTAIL.n261 VTAIL.n260 9.3005
R529 VTAIL.n230 VTAIL.n229 9.3005
R530 VTAIL.n255 VTAIL.n254 9.3005
R531 VTAIL.n253 VTAIL.n252 9.3005
R532 VTAIL.n234 VTAIL.n233 9.3005
R533 VTAIL.n247 VTAIL.n246 9.3005
R534 VTAIL.n245 VTAIL.n244 9.3005
R535 VTAIL.n238 VTAIL.n237 9.3005
R536 VTAIL.n544 VTAIL.n543 8.92171
R537 VTAIL.n559 VTAIL.n512 8.92171
R538 VTAIL.n40 VTAIL.n39 8.92171
R539 VTAIL.n55 VTAIL.n8 8.92171
R540 VTAIL.n112 VTAIL.n111 8.92171
R541 VTAIL.n127 VTAIL.n80 8.92171
R542 VTAIL.n184 VTAIL.n183 8.92171
R543 VTAIL.n199 VTAIL.n152 8.92171
R544 VTAIL.n487 VTAIL.n440 8.92171
R545 VTAIL.n472 VTAIL.n471 8.92171
R546 VTAIL.n415 VTAIL.n368 8.92171
R547 VTAIL.n400 VTAIL.n399 8.92171
R548 VTAIL.n343 VTAIL.n296 8.92171
R549 VTAIL.n328 VTAIL.n327 8.92171
R550 VTAIL.n271 VTAIL.n224 8.92171
R551 VTAIL.n256 VTAIL.n255 8.92171
R552 VTAIL.n574 VTAIL.n504 8.2187
R553 VTAIL.n70 VTAIL.n0 8.2187
R554 VTAIL.n142 VTAIL.n72 8.2187
R555 VTAIL.n214 VTAIL.n144 8.2187
R556 VTAIL.n502 VTAIL.n432 8.2187
R557 VTAIL.n430 VTAIL.n360 8.2187
R558 VTAIL.n358 VTAIL.n288 8.2187
R559 VTAIL.n286 VTAIL.n216 8.2187
R560 VTAIL.n547 VTAIL.n518 8.14595
R561 VTAIL.n556 VTAIL.n555 8.14595
R562 VTAIL.n43 VTAIL.n14 8.14595
R563 VTAIL.n52 VTAIL.n51 8.14595
R564 VTAIL.n115 VTAIL.n86 8.14595
R565 VTAIL.n124 VTAIL.n123 8.14595
R566 VTAIL.n187 VTAIL.n158 8.14595
R567 VTAIL.n196 VTAIL.n195 8.14595
R568 VTAIL.n484 VTAIL.n483 8.14595
R569 VTAIL.n475 VTAIL.n446 8.14595
R570 VTAIL.n412 VTAIL.n411 8.14595
R571 VTAIL.n403 VTAIL.n374 8.14595
R572 VTAIL.n340 VTAIL.n339 8.14595
R573 VTAIL.n331 VTAIL.n302 8.14595
R574 VTAIL.n268 VTAIL.n267 8.14595
R575 VTAIL.n259 VTAIL.n230 8.14595
R576 VTAIL.n548 VTAIL.n516 7.3702
R577 VTAIL.n552 VTAIL.n514 7.3702
R578 VTAIL.n44 VTAIL.n12 7.3702
R579 VTAIL.n48 VTAIL.n10 7.3702
R580 VTAIL.n116 VTAIL.n84 7.3702
R581 VTAIL.n120 VTAIL.n82 7.3702
R582 VTAIL.n188 VTAIL.n156 7.3702
R583 VTAIL.n192 VTAIL.n154 7.3702
R584 VTAIL.n480 VTAIL.n442 7.3702
R585 VTAIL.n476 VTAIL.n444 7.3702
R586 VTAIL.n408 VTAIL.n370 7.3702
R587 VTAIL.n404 VTAIL.n372 7.3702
R588 VTAIL.n336 VTAIL.n298 7.3702
R589 VTAIL.n332 VTAIL.n300 7.3702
R590 VTAIL.n264 VTAIL.n226 7.3702
R591 VTAIL.n260 VTAIL.n228 7.3702
R592 VTAIL.n551 VTAIL.n516 6.59444
R593 VTAIL.n552 VTAIL.n551 6.59444
R594 VTAIL.n47 VTAIL.n12 6.59444
R595 VTAIL.n48 VTAIL.n47 6.59444
R596 VTAIL.n119 VTAIL.n84 6.59444
R597 VTAIL.n120 VTAIL.n119 6.59444
R598 VTAIL.n191 VTAIL.n156 6.59444
R599 VTAIL.n192 VTAIL.n191 6.59444
R600 VTAIL.n480 VTAIL.n479 6.59444
R601 VTAIL.n479 VTAIL.n444 6.59444
R602 VTAIL.n408 VTAIL.n407 6.59444
R603 VTAIL.n407 VTAIL.n372 6.59444
R604 VTAIL.n336 VTAIL.n335 6.59444
R605 VTAIL.n335 VTAIL.n300 6.59444
R606 VTAIL.n264 VTAIL.n263 6.59444
R607 VTAIL.n263 VTAIL.n228 6.59444
R608 VTAIL.n548 VTAIL.n547 5.81868
R609 VTAIL.n555 VTAIL.n514 5.81868
R610 VTAIL.n44 VTAIL.n43 5.81868
R611 VTAIL.n51 VTAIL.n10 5.81868
R612 VTAIL.n116 VTAIL.n115 5.81868
R613 VTAIL.n123 VTAIL.n82 5.81868
R614 VTAIL.n188 VTAIL.n187 5.81868
R615 VTAIL.n195 VTAIL.n154 5.81868
R616 VTAIL.n483 VTAIL.n442 5.81868
R617 VTAIL.n476 VTAIL.n475 5.81868
R618 VTAIL.n411 VTAIL.n370 5.81868
R619 VTAIL.n404 VTAIL.n403 5.81868
R620 VTAIL.n339 VTAIL.n298 5.81868
R621 VTAIL.n332 VTAIL.n331 5.81868
R622 VTAIL.n267 VTAIL.n226 5.81868
R623 VTAIL.n260 VTAIL.n259 5.81868
R624 VTAIL.n572 VTAIL.n504 5.3904
R625 VTAIL.n68 VTAIL.n0 5.3904
R626 VTAIL.n140 VTAIL.n72 5.3904
R627 VTAIL.n212 VTAIL.n144 5.3904
R628 VTAIL.n500 VTAIL.n432 5.3904
R629 VTAIL.n428 VTAIL.n360 5.3904
R630 VTAIL.n356 VTAIL.n288 5.3904
R631 VTAIL.n284 VTAIL.n216 5.3904
R632 VTAIL.n544 VTAIL.n518 5.04292
R633 VTAIL.n556 VTAIL.n512 5.04292
R634 VTAIL.n40 VTAIL.n14 5.04292
R635 VTAIL.n52 VTAIL.n8 5.04292
R636 VTAIL.n112 VTAIL.n86 5.04292
R637 VTAIL.n124 VTAIL.n80 5.04292
R638 VTAIL.n184 VTAIL.n158 5.04292
R639 VTAIL.n196 VTAIL.n152 5.04292
R640 VTAIL.n484 VTAIL.n440 5.04292
R641 VTAIL.n472 VTAIL.n446 5.04292
R642 VTAIL.n412 VTAIL.n368 5.04292
R643 VTAIL.n400 VTAIL.n374 5.04292
R644 VTAIL.n340 VTAIL.n296 5.04292
R645 VTAIL.n328 VTAIL.n302 5.04292
R646 VTAIL.n268 VTAIL.n224 5.04292
R647 VTAIL.n256 VTAIL.n230 5.04292
R648 VTAIL.n527 VTAIL.n525 4.38563
R649 VTAIL.n23 VTAIL.n21 4.38563
R650 VTAIL.n95 VTAIL.n93 4.38563
R651 VTAIL.n167 VTAIL.n165 4.38563
R652 VTAIL.n455 VTAIL.n453 4.38563
R653 VTAIL.n383 VTAIL.n381 4.38563
R654 VTAIL.n311 VTAIL.n309 4.38563
R655 VTAIL.n239 VTAIL.n237 4.38563
R656 VTAIL.n543 VTAIL.n520 4.26717
R657 VTAIL.n560 VTAIL.n559 4.26717
R658 VTAIL.n39 VTAIL.n16 4.26717
R659 VTAIL.n56 VTAIL.n55 4.26717
R660 VTAIL.n111 VTAIL.n88 4.26717
R661 VTAIL.n128 VTAIL.n127 4.26717
R662 VTAIL.n183 VTAIL.n160 4.26717
R663 VTAIL.n200 VTAIL.n199 4.26717
R664 VTAIL.n488 VTAIL.n487 4.26717
R665 VTAIL.n471 VTAIL.n448 4.26717
R666 VTAIL.n416 VTAIL.n415 4.26717
R667 VTAIL.n399 VTAIL.n376 4.26717
R668 VTAIL.n344 VTAIL.n343 4.26717
R669 VTAIL.n327 VTAIL.n304 4.26717
R670 VTAIL.n272 VTAIL.n271 4.26717
R671 VTAIL.n255 VTAIL.n232 4.26717
R672 VTAIL.n540 VTAIL.n539 3.49141
R673 VTAIL.n563 VTAIL.n510 3.49141
R674 VTAIL.n36 VTAIL.n35 3.49141
R675 VTAIL.n59 VTAIL.n6 3.49141
R676 VTAIL.n108 VTAIL.n107 3.49141
R677 VTAIL.n131 VTAIL.n78 3.49141
R678 VTAIL.n180 VTAIL.n179 3.49141
R679 VTAIL.n203 VTAIL.n150 3.49141
R680 VTAIL.n491 VTAIL.n438 3.49141
R681 VTAIL.n468 VTAIL.n467 3.49141
R682 VTAIL.n419 VTAIL.n366 3.49141
R683 VTAIL.n396 VTAIL.n395 3.49141
R684 VTAIL.n347 VTAIL.n294 3.49141
R685 VTAIL.n324 VTAIL.n323 3.49141
R686 VTAIL.n275 VTAIL.n222 3.49141
R687 VTAIL.n252 VTAIL.n251 3.49141
R688 VTAIL.n536 VTAIL.n522 2.71565
R689 VTAIL.n564 VTAIL.n508 2.71565
R690 VTAIL.n32 VTAIL.n18 2.71565
R691 VTAIL.n60 VTAIL.n4 2.71565
R692 VTAIL.n104 VTAIL.n90 2.71565
R693 VTAIL.n132 VTAIL.n76 2.71565
R694 VTAIL.n176 VTAIL.n162 2.71565
R695 VTAIL.n204 VTAIL.n148 2.71565
R696 VTAIL.n492 VTAIL.n436 2.71565
R697 VTAIL.n464 VTAIL.n450 2.71565
R698 VTAIL.n420 VTAIL.n364 2.71565
R699 VTAIL.n392 VTAIL.n378 2.71565
R700 VTAIL.n348 VTAIL.n292 2.71565
R701 VTAIL.n320 VTAIL.n306 2.71565
R702 VTAIL.n276 VTAIL.n220 2.71565
R703 VTAIL.n248 VTAIL.n234 2.71565
R704 VTAIL.n535 VTAIL.n524 1.93989
R705 VTAIL.n568 VTAIL.n567 1.93989
R706 VTAIL.n31 VTAIL.n20 1.93989
R707 VTAIL.n64 VTAIL.n63 1.93989
R708 VTAIL.n103 VTAIL.n92 1.93989
R709 VTAIL.n136 VTAIL.n135 1.93989
R710 VTAIL.n175 VTAIL.n164 1.93989
R711 VTAIL.n208 VTAIL.n207 1.93989
R712 VTAIL.n496 VTAIL.n495 1.93989
R713 VTAIL.n463 VTAIL.n452 1.93989
R714 VTAIL.n424 VTAIL.n423 1.93989
R715 VTAIL.n391 VTAIL.n380 1.93989
R716 VTAIL.n352 VTAIL.n351 1.93989
R717 VTAIL.n319 VTAIL.n308 1.93989
R718 VTAIL.n280 VTAIL.n279 1.93989
R719 VTAIL.n247 VTAIL.n236 1.93989
R720 VTAIL.n359 VTAIL.n287 1.28498
R721 VTAIL.n503 VTAIL.n431 1.28498
R722 VTAIL.n215 VTAIL.n143 1.28498
R723 VTAIL.n532 VTAIL.n531 1.16414
R724 VTAIL.n571 VTAIL.n506 1.16414
R725 VTAIL.n28 VTAIL.n27 1.16414
R726 VTAIL.n67 VTAIL.n2 1.16414
R727 VTAIL.n100 VTAIL.n99 1.16414
R728 VTAIL.n139 VTAIL.n74 1.16414
R729 VTAIL.n172 VTAIL.n171 1.16414
R730 VTAIL.n211 VTAIL.n146 1.16414
R731 VTAIL.n499 VTAIL.n434 1.16414
R732 VTAIL.n460 VTAIL.n459 1.16414
R733 VTAIL.n427 VTAIL.n362 1.16414
R734 VTAIL.n388 VTAIL.n387 1.16414
R735 VTAIL.n355 VTAIL.n290 1.16414
R736 VTAIL.n316 VTAIL.n315 1.16414
R737 VTAIL.n283 VTAIL.n218 1.16414
R738 VTAIL.n244 VTAIL.n243 1.16414
R739 VTAIL VTAIL.n71 0.700931
R740 VTAIL VTAIL.n575 0.584552
R741 VTAIL.n431 VTAIL.n359 0.470328
R742 VTAIL.n143 VTAIL.n71 0.470328
R743 VTAIL.n528 VTAIL.n526 0.388379
R744 VTAIL.n24 VTAIL.n22 0.388379
R745 VTAIL.n96 VTAIL.n94 0.388379
R746 VTAIL.n168 VTAIL.n166 0.388379
R747 VTAIL.n456 VTAIL.n454 0.388379
R748 VTAIL.n384 VTAIL.n382 0.388379
R749 VTAIL.n312 VTAIL.n310 0.388379
R750 VTAIL.n240 VTAIL.n238 0.388379
R751 VTAIL.n533 VTAIL.n525 0.155672
R752 VTAIL.n534 VTAIL.n533 0.155672
R753 VTAIL.n534 VTAIL.n521 0.155672
R754 VTAIL.n541 VTAIL.n521 0.155672
R755 VTAIL.n542 VTAIL.n541 0.155672
R756 VTAIL.n542 VTAIL.n517 0.155672
R757 VTAIL.n549 VTAIL.n517 0.155672
R758 VTAIL.n550 VTAIL.n549 0.155672
R759 VTAIL.n550 VTAIL.n513 0.155672
R760 VTAIL.n557 VTAIL.n513 0.155672
R761 VTAIL.n558 VTAIL.n557 0.155672
R762 VTAIL.n558 VTAIL.n509 0.155672
R763 VTAIL.n565 VTAIL.n509 0.155672
R764 VTAIL.n566 VTAIL.n565 0.155672
R765 VTAIL.n566 VTAIL.n505 0.155672
R766 VTAIL.n573 VTAIL.n505 0.155672
R767 VTAIL.n29 VTAIL.n21 0.155672
R768 VTAIL.n30 VTAIL.n29 0.155672
R769 VTAIL.n30 VTAIL.n17 0.155672
R770 VTAIL.n37 VTAIL.n17 0.155672
R771 VTAIL.n38 VTAIL.n37 0.155672
R772 VTAIL.n38 VTAIL.n13 0.155672
R773 VTAIL.n45 VTAIL.n13 0.155672
R774 VTAIL.n46 VTAIL.n45 0.155672
R775 VTAIL.n46 VTAIL.n9 0.155672
R776 VTAIL.n53 VTAIL.n9 0.155672
R777 VTAIL.n54 VTAIL.n53 0.155672
R778 VTAIL.n54 VTAIL.n5 0.155672
R779 VTAIL.n61 VTAIL.n5 0.155672
R780 VTAIL.n62 VTAIL.n61 0.155672
R781 VTAIL.n62 VTAIL.n1 0.155672
R782 VTAIL.n69 VTAIL.n1 0.155672
R783 VTAIL.n101 VTAIL.n93 0.155672
R784 VTAIL.n102 VTAIL.n101 0.155672
R785 VTAIL.n102 VTAIL.n89 0.155672
R786 VTAIL.n109 VTAIL.n89 0.155672
R787 VTAIL.n110 VTAIL.n109 0.155672
R788 VTAIL.n110 VTAIL.n85 0.155672
R789 VTAIL.n117 VTAIL.n85 0.155672
R790 VTAIL.n118 VTAIL.n117 0.155672
R791 VTAIL.n118 VTAIL.n81 0.155672
R792 VTAIL.n125 VTAIL.n81 0.155672
R793 VTAIL.n126 VTAIL.n125 0.155672
R794 VTAIL.n126 VTAIL.n77 0.155672
R795 VTAIL.n133 VTAIL.n77 0.155672
R796 VTAIL.n134 VTAIL.n133 0.155672
R797 VTAIL.n134 VTAIL.n73 0.155672
R798 VTAIL.n141 VTAIL.n73 0.155672
R799 VTAIL.n173 VTAIL.n165 0.155672
R800 VTAIL.n174 VTAIL.n173 0.155672
R801 VTAIL.n174 VTAIL.n161 0.155672
R802 VTAIL.n181 VTAIL.n161 0.155672
R803 VTAIL.n182 VTAIL.n181 0.155672
R804 VTAIL.n182 VTAIL.n157 0.155672
R805 VTAIL.n189 VTAIL.n157 0.155672
R806 VTAIL.n190 VTAIL.n189 0.155672
R807 VTAIL.n190 VTAIL.n153 0.155672
R808 VTAIL.n197 VTAIL.n153 0.155672
R809 VTAIL.n198 VTAIL.n197 0.155672
R810 VTAIL.n198 VTAIL.n149 0.155672
R811 VTAIL.n205 VTAIL.n149 0.155672
R812 VTAIL.n206 VTAIL.n205 0.155672
R813 VTAIL.n206 VTAIL.n145 0.155672
R814 VTAIL.n213 VTAIL.n145 0.155672
R815 VTAIL.n501 VTAIL.n433 0.155672
R816 VTAIL.n494 VTAIL.n433 0.155672
R817 VTAIL.n494 VTAIL.n493 0.155672
R818 VTAIL.n493 VTAIL.n437 0.155672
R819 VTAIL.n486 VTAIL.n437 0.155672
R820 VTAIL.n486 VTAIL.n485 0.155672
R821 VTAIL.n485 VTAIL.n441 0.155672
R822 VTAIL.n478 VTAIL.n441 0.155672
R823 VTAIL.n478 VTAIL.n477 0.155672
R824 VTAIL.n477 VTAIL.n445 0.155672
R825 VTAIL.n470 VTAIL.n445 0.155672
R826 VTAIL.n470 VTAIL.n469 0.155672
R827 VTAIL.n469 VTAIL.n449 0.155672
R828 VTAIL.n462 VTAIL.n449 0.155672
R829 VTAIL.n462 VTAIL.n461 0.155672
R830 VTAIL.n461 VTAIL.n453 0.155672
R831 VTAIL.n429 VTAIL.n361 0.155672
R832 VTAIL.n422 VTAIL.n361 0.155672
R833 VTAIL.n422 VTAIL.n421 0.155672
R834 VTAIL.n421 VTAIL.n365 0.155672
R835 VTAIL.n414 VTAIL.n365 0.155672
R836 VTAIL.n414 VTAIL.n413 0.155672
R837 VTAIL.n413 VTAIL.n369 0.155672
R838 VTAIL.n406 VTAIL.n369 0.155672
R839 VTAIL.n406 VTAIL.n405 0.155672
R840 VTAIL.n405 VTAIL.n373 0.155672
R841 VTAIL.n398 VTAIL.n373 0.155672
R842 VTAIL.n398 VTAIL.n397 0.155672
R843 VTAIL.n397 VTAIL.n377 0.155672
R844 VTAIL.n390 VTAIL.n377 0.155672
R845 VTAIL.n390 VTAIL.n389 0.155672
R846 VTAIL.n389 VTAIL.n381 0.155672
R847 VTAIL.n357 VTAIL.n289 0.155672
R848 VTAIL.n350 VTAIL.n289 0.155672
R849 VTAIL.n350 VTAIL.n349 0.155672
R850 VTAIL.n349 VTAIL.n293 0.155672
R851 VTAIL.n342 VTAIL.n293 0.155672
R852 VTAIL.n342 VTAIL.n341 0.155672
R853 VTAIL.n341 VTAIL.n297 0.155672
R854 VTAIL.n334 VTAIL.n297 0.155672
R855 VTAIL.n334 VTAIL.n333 0.155672
R856 VTAIL.n333 VTAIL.n301 0.155672
R857 VTAIL.n326 VTAIL.n301 0.155672
R858 VTAIL.n326 VTAIL.n325 0.155672
R859 VTAIL.n325 VTAIL.n305 0.155672
R860 VTAIL.n318 VTAIL.n305 0.155672
R861 VTAIL.n318 VTAIL.n317 0.155672
R862 VTAIL.n317 VTAIL.n309 0.155672
R863 VTAIL.n285 VTAIL.n217 0.155672
R864 VTAIL.n278 VTAIL.n217 0.155672
R865 VTAIL.n278 VTAIL.n277 0.155672
R866 VTAIL.n277 VTAIL.n221 0.155672
R867 VTAIL.n270 VTAIL.n221 0.155672
R868 VTAIL.n270 VTAIL.n269 0.155672
R869 VTAIL.n269 VTAIL.n225 0.155672
R870 VTAIL.n262 VTAIL.n225 0.155672
R871 VTAIL.n262 VTAIL.n261 0.155672
R872 VTAIL.n261 VTAIL.n229 0.155672
R873 VTAIL.n254 VTAIL.n229 0.155672
R874 VTAIL.n254 VTAIL.n253 0.155672
R875 VTAIL.n253 VTAIL.n233 0.155672
R876 VTAIL.n246 VTAIL.n233 0.155672
R877 VTAIL.n246 VTAIL.n245 0.155672
R878 VTAIL.n245 VTAIL.n237 0.155672
R879 VDD2.n2 VDD2.n0 102.296
R880 VDD2.n2 VDD2.n1 63.2528
R881 VDD2.n1 VDD2.t2 1.4881
R882 VDD2.n1 VDD2.t1 1.4881
R883 VDD2.n0 VDD2.t0 1.4881
R884 VDD2.n0 VDD2.t3 1.4881
R885 VDD2 VDD2.n2 0.0586897
R886 B.n681 B.n680 585
R887 B.n294 B.n91 585
R888 B.n293 B.n292 585
R889 B.n291 B.n290 585
R890 B.n289 B.n288 585
R891 B.n287 B.n286 585
R892 B.n285 B.n284 585
R893 B.n283 B.n282 585
R894 B.n281 B.n280 585
R895 B.n279 B.n278 585
R896 B.n277 B.n276 585
R897 B.n275 B.n274 585
R898 B.n273 B.n272 585
R899 B.n271 B.n270 585
R900 B.n269 B.n268 585
R901 B.n267 B.n266 585
R902 B.n265 B.n264 585
R903 B.n263 B.n262 585
R904 B.n261 B.n260 585
R905 B.n259 B.n258 585
R906 B.n257 B.n256 585
R907 B.n255 B.n254 585
R908 B.n253 B.n252 585
R909 B.n251 B.n250 585
R910 B.n249 B.n248 585
R911 B.n247 B.n246 585
R912 B.n245 B.n244 585
R913 B.n243 B.n242 585
R914 B.n241 B.n240 585
R915 B.n239 B.n238 585
R916 B.n237 B.n236 585
R917 B.n235 B.n234 585
R918 B.n233 B.n232 585
R919 B.n231 B.n230 585
R920 B.n229 B.n228 585
R921 B.n227 B.n226 585
R922 B.n225 B.n224 585
R923 B.n223 B.n222 585
R924 B.n221 B.n220 585
R925 B.n219 B.n218 585
R926 B.n217 B.n216 585
R927 B.n215 B.n214 585
R928 B.n213 B.n212 585
R929 B.n211 B.n210 585
R930 B.n209 B.n208 585
R931 B.n206 B.n205 585
R932 B.n204 B.n203 585
R933 B.n202 B.n201 585
R934 B.n200 B.n199 585
R935 B.n198 B.n197 585
R936 B.n196 B.n195 585
R937 B.n194 B.n193 585
R938 B.n192 B.n191 585
R939 B.n190 B.n189 585
R940 B.n188 B.n187 585
R941 B.n185 B.n184 585
R942 B.n183 B.n182 585
R943 B.n181 B.n180 585
R944 B.n179 B.n178 585
R945 B.n177 B.n176 585
R946 B.n175 B.n174 585
R947 B.n173 B.n172 585
R948 B.n171 B.n170 585
R949 B.n169 B.n168 585
R950 B.n167 B.n166 585
R951 B.n165 B.n164 585
R952 B.n163 B.n162 585
R953 B.n161 B.n160 585
R954 B.n159 B.n158 585
R955 B.n157 B.n156 585
R956 B.n155 B.n154 585
R957 B.n153 B.n152 585
R958 B.n151 B.n150 585
R959 B.n149 B.n148 585
R960 B.n147 B.n146 585
R961 B.n145 B.n144 585
R962 B.n143 B.n142 585
R963 B.n141 B.n140 585
R964 B.n139 B.n138 585
R965 B.n137 B.n136 585
R966 B.n135 B.n134 585
R967 B.n133 B.n132 585
R968 B.n131 B.n130 585
R969 B.n129 B.n128 585
R970 B.n127 B.n126 585
R971 B.n125 B.n124 585
R972 B.n123 B.n122 585
R973 B.n121 B.n120 585
R974 B.n119 B.n118 585
R975 B.n117 B.n116 585
R976 B.n115 B.n114 585
R977 B.n113 B.n112 585
R978 B.n111 B.n110 585
R979 B.n109 B.n108 585
R980 B.n107 B.n106 585
R981 B.n105 B.n104 585
R982 B.n103 B.n102 585
R983 B.n101 B.n100 585
R984 B.n99 B.n98 585
R985 B.n97 B.n96 585
R986 B.n679 B.n41 585
R987 B.n684 B.n41 585
R988 B.n678 B.n40 585
R989 B.n685 B.n40 585
R990 B.n677 B.n676 585
R991 B.n676 B.n36 585
R992 B.n675 B.n35 585
R993 B.n691 B.n35 585
R994 B.n674 B.n34 585
R995 B.n692 B.n34 585
R996 B.n673 B.n33 585
R997 B.n693 B.n33 585
R998 B.n672 B.n671 585
R999 B.n671 B.n29 585
R1000 B.n670 B.n28 585
R1001 B.n699 B.n28 585
R1002 B.n669 B.n27 585
R1003 B.n700 B.n27 585
R1004 B.n668 B.n26 585
R1005 B.n701 B.n26 585
R1006 B.n667 B.n666 585
R1007 B.n666 B.n22 585
R1008 B.n665 B.n21 585
R1009 B.n707 B.n21 585
R1010 B.n664 B.n20 585
R1011 B.n708 B.n20 585
R1012 B.n663 B.n19 585
R1013 B.n709 B.n19 585
R1014 B.n662 B.n661 585
R1015 B.n661 B.n15 585
R1016 B.n660 B.n14 585
R1017 B.n715 B.n14 585
R1018 B.n659 B.n13 585
R1019 B.n716 B.n13 585
R1020 B.n658 B.n12 585
R1021 B.n717 B.n12 585
R1022 B.n657 B.n656 585
R1023 B.n656 B.n8 585
R1024 B.n655 B.n7 585
R1025 B.n723 B.n7 585
R1026 B.n654 B.n6 585
R1027 B.n724 B.n6 585
R1028 B.n653 B.n5 585
R1029 B.n725 B.n5 585
R1030 B.n652 B.n651 585
R1031 B.n651 B.n4 585
R1032 B.n650 B.n295 585
R1033 B.n650 B.n649 585
R1034 B.n640 B.n296 585
R1035 B.n297 B.n296 585
R1036 B.n642 B.n641 585
R1037 B.n643 B.n642 585
R1038 B.n639 B.n302 585
R1039 B.n302 B.n301 585
R1040 B.n638 B.n637 585
R1041 B.n637 B.n636 585
R1042 B.n304 B.n303 585
R1043 B.n305 B.n304 585
R1044 B.n629 B.n628 585
R1045 B.n630 B.n629 585
R1046 B.n627 B.n309 585
R1047 B.n313 B.n309 585
R1048 B.n626 B.n625 585
R1049 B.n625 B.n624 585
R1050 B.n311 B.n310 585
R1051 B.n312 B.n311 585
R1052 B.n617 B.n616 585
R1053 B.n618 B.n617 585
R1054 B.n615 B.n318 585
R1055 B.n318 B.n317 585
R1056 B.n614 B.n613 585
R1057 B.n613 B.n612 585
R1058 B.n320 B.n319 585
R1059 B.n321 B.n320 585
R1060 B.n605 B.n604 585
R1061 B.n606 B.n605 585
R1062 B.n603 B.n326 585
R1063 B.n326 B.n325 585
R1064 B.n602 B.n601 585
R1065 B.n601 B.n600 585
R1066 B.n328 B.n327 585
R1067 B.n329 B.n328 585
R1068 B.n593 B.n592 585
R1069 B.n594 B.n593 585
R1070 B.n591 B.n334 585
R1071 B.n334 B.n333 585
R1072 B.n586 B.n585 585
R1073 B.n584 B.n386 585
R1074 B.n583 B.n385 585
R1075 B.n588 B.n385 585
R1076 B.n582 B.n581 585
R1077 B.n580 B.n579 585
R1078 B.n578 B.n577 585
R1079 B.n576 B.n575 585
R1080 B.n574 B.n573 585
R1081 B.n572 B.n571 585
R1082 B.n570 B.n569 585
R1083 B.n568 B.n567 585
R1084 B.n566 B.n565 585
R1085 B.n564 B.n563 585
R1086 B.n562 B.n561 585
R1087 B.n560 B.n559 585
R1088 B.n558 B.n557 585
R1089 B.n556 B.n555 585
R1090 B.n554 B.n553 585
R1091 B.n552 B.n551 585
R1092 B.n550 B.n549 585
R1093 B.n548 B.n547 585
R1094 B.n546 B.n545 585
R1095 B.n544 B.n543 585
R1096 B.n542 B.n541 585
R1097 B.n540 B.n539 585
R1098 B.n538 B.n537 585
R1099 B.n536 B.n535 585
R1100 B.n534 B.n533 585
R1101 B.n532 B.n531 585
R1102 B.n530 B.n529 585
R1103 B.n528 B.n527 585
R1104 B.n526 B.n525 585
R1105 B.n524 B.n523 585
R1106 B.n522 B.n521 585
R1107 B.n520 B.n519 585
R1108 B.n518 B.n517 585
R1109 B.n516 B.n515 585
R1110 B.n514 B.n513 585
R1111 B.n512 B.n511 585
R1112 B.n510 B.n509 585
R1113 B.n508 B.n507 585
R1114 B.n506 B.n505 585
R1115 B.n504 B.n503 585
R1116 B.n502 B.n501 585
R1117 B.n500 B.n499 585
R1118 B.n498 B.n497 585
R1119 B.n496 B.n495 585
R1120 B.n494 B.n493 585
R1121 B.n492 B.n491 585
R1122 B.n490 B.n489 585
R1123 B.n488 B.n487 585
R1124 B.n486 B.n485 585
R1125 B.n484 B.n483 585
R1126 B.n482 B.n481 585
R1127 B.n480 B.n479 585
R1128 B.n478 B.n477 585
R1129 B.n476 B.n475 585
R1130 B.n474 B.n473 585
R1131 B.n472 B.n471 585
R1132 B.n470 B.n469 585
R1133 B.n468 B.n467 585
R1134 B.n466 B.n465 585
R1135 B.n464 B.n463 585
R1136 B.n462 B.n461 585
R1137 B.n460 B.n459 585
R1138 B.n458 B.n457 585
R1139 B.n456 B.n455 585
R1140 B.n454 B.n453 585
R1141 B.n452 B.n451 585
R1142 B.n450 B.n449 585
R1143 B.n448 B.n447 585
R1144 B.n446 B.n445 585
R1145 B.n444 B.n443 585
R1146 B.n442 B.n441 585
R1147 B.n440 B.n439 585
R1148 B.n438 B.n437 585
R1149 B.n436 B.n435 585
R1150 B.n434 B.n433 585
R1151 B.n432 B.n431 585
R1152 B.n430 B.n429 585
R1153 B.n428 B.n427 585
R1154 B.n426 B.n425 585
R1155 B.n424 B.n423 585
R1156 B.n422 B.n421 585
R1157 B.n420 B.n419 585
R1158 B.n418 B.n417 585
R1159 B.n416 B.n415 585
R1160 B.n414 B.n413 585
R1161 B.n412 B.n411 585
R1162 B.n410 B.n409 585
R1163 B.n408 B.n407 585
R1164 B.n406 B.n405 585
R1165 B.n404 B.n403 585
R1166 B.n402 B.n401 585
R1167 B.n400 B.n399 585
R1168 B.n398 B.n397 585
R1169 B.n396 B.n395 585
R1170 B.n394 B.n393 585
R1171 B.n336 B.n335 585
R1172 B.n590 B.n589 585
R1173 B.n589 B.n588 585
R1174 B.n332 B.n331 585
R1175 B.n333 B.n332 585
R1176 B.n596 B.n595 585
R1177 B.n595 B.n594 585
R1178 B.n597 B.n330 585
R1179 B.n330 B.n329 585
R1180 B.n599 B.n598 585
R1181 B.n600 B.n599 585
R1182 B.n324 B.n323 585
R1183 B.n325 B.n324 585
R1184 B.n608 B.n607 585
R1185 B.n607 B.n606 585
R1186 B.n609 B.n322 585
R1187 B.n322 B.n321 585
R1188 B.n611 B.n610 585
R1189 B.n612 B.n611 585
R1190 B.n316 B.n315 585
R1191 B.n317 B.n316 585
R1192 B.n620 B.n619 585
R1193 B.n619 B.n618 585
R1194 B.n621 B.n314 585
R1195 B.n314 B.n312 585
R1196 B.n623 B.n622 585
R1197 B.n624 B.n623 585
R1198 B.n308 B.n307 585
R1199 B.n313 B.n308 585
R1200 B.n632 B.n631 585
R1201 B.n631 B.n630 585
R1202 B.n633 B.n306 585
R1203 B.n306 B.n305 585
R1204 B.n635 B.n634 585
R1205 B.n636 B.n635 585
R1206 B.n300 B.n299 585
R1207 B.n301 B.n300 585
R1208 B.n645 B.n644 585
R1209 B.n644 B.n643 585
R1210 B.n646 B.n298 585
R1211 B.n298 B.n297 585
R1212 B.n648 B.n647 585
R1213 B.n649 B.n648 585
R1214 B.n2 B.n0 585
R1215 B.n4 B.n2 585
R1216 B.n3 B.n1 585
R1217 B.n724 B.n3 585
R1218 B.n722 B.n721 585
R1219 B.n723 B.n722 585
R1220 B.n720 B.n9 585
R1221 B.n9 B.n8 585
R1222 B.n719 B.n718 585
R1223 B.n718 B.n717 585
R1224 B.n11 B.n10 585
R1225 B.n716 B.n11 585
R1226 B.n714 B.n713 585
R1227 B.n715 B.n714 585
R1228 B.n712 B.n16 585
R1229 B.n16 B.n15 585
R1230 B.n711 B.n710 585
R1231 B.n710 B.n709 585
R1232 B.n18 B.n17 585
R1233 B.n708 B.n18 585
R1234 B.n706 B.n705 585
R1235 B.n707 B.n706 585
R1236 B.n704 B.n23 585
R1237 B.n23 B.n22 585
R1238 B.n703 B.n702 585
R1239 B.n702 B.n701 585
R1240 B.n25 B.n24 585
R1241 B.n700 B.n25 585
R1242 B.n698 B.n697 585
R1243 B.n699 B.n698 585
R1244 B.n696 B.n30 585
R1245 B.n30 B.n29 585
R1246 B.n695 B.n694 585
R1247 B.n694 B.n693 585
R1248 B.n32 B.n31 585
R1249 B.n692 B.n32 585
R1250 B.n690 B.n689 585
R1251 B.n691 B.n690 585
R1252 B.n688 B.n37 585
R1253 B.n37 B.n36 585
R1254 B.n687 B.n686 585
R1255 B.n686 B.n685 585
R1256 B.n39 B.n38 585
R1257 B.n684 B.n39 585
R1258 B.n727 B.n726 585
R1259 B.n726 B.n725 585
R1260 B.n586 B.n332 583.793
R1261 B.n96 B.n39 583.793
R1262 B.n589 B.n334 583.793
R1263 B.n681 B.n41 583.793
R1264 B.n390 B.t4 480.43
R1265 B.n387 B.t8 480.43
R1266 B.n94 B.t15 480.43
R1267 B.n92 B.t11 480.43
R1268 B.n390 B.t7 333.361
R1269 B.n92 B.t13 333.361
R1270 B.n387 B.t10 333.361
R1271 B.n94 B.t16 333.361
R1272 B.n391 B.t6 304.464
R1273 B.n93 B.t14 304.464
R1274 B.n388 B.t9 304.464
R1275 B.n95 B.t17 304.464
R1276 B.n683 B.n682 256.663
R1277 B.n683 B.n90 256.663
R1278 B.n683 B.n89 256.663
R1279 B.n683 B.n88 256.663
R1280 B.n683 B.n87 256.663
R1281 B.n683 B.n86 256.663
R1282 B.n683 B.n85 256.663
R1283 B.n683 B.n84 256.663
R1284 B.n683 B.n83 256.663
R1285 B.n683 B.n82 256.663
R1286 B.n683 B.n81 256.663
R1287 B.n683 B.n80 256.663
R1288 B.n683 B.n79 256.663
R1289 B.n683 B.n78 256.663
R1290 B.n683 B.n77 256.663
R1291 B.n683 B.n76 256.663
R1292 B.n683 B.n75 256.663
R1293 B.n683 B.n74 256.663
R1294 B.n683 B.n73 256.663
R1295 B.n683 B.n72 256.663
R1296 B.n683 B.n71 256.663
R1297 B.n683 B.n70 256.663
R1298 B.n683 B.n69 256.663
R1299 B.n683 B.n68 256.663
R1300 B.n683 B.n67 256.663
R1301 B.n683 B.n66 256.663
R1302 B.n683 B.n65 256.663
R1303 B.n683 B.n64 256.663
R1304 B.n683 B.n63 256.663
R1305 B.n683 B.n62 256.663
R1306 B.n683 B.n61 256.663
R1307 B.n683 B.n60 256.663
R1308 B.n683 B.n59 256.663
R1309 B.n683 B.n58 256.663
R1310 B.n683 B.n57 256.663
R1311 B.n683 B.n56 256.663
R1312 B.n683 B.n55 256.663
R1313 B.n683 B.n54 256.663
R1314 B.n683 B.n53 256.663
R1315 B.n683 B.n52 256.663
R1316 B.n683 B.n51 256.663
R1317 B.n683 B.n50 256.663
R1318 B.n683 B.n49 256.663
R1319 B.n683 B.n48 256.663
R1320 B.n683 B.n47 256.663
R1321 B.n683 B.n46 256.663
R1322 B.n683 B.n45 256.663
R1323 B.n683 B.n44 256.663
R1324 B.n683 B.n43 256.663
R1325 B.n683 B.n42 256.663
R1326 B.n588 B.n587 256.663
R1327 B.n588 B.n337 256.663
R1328 B.n588 B.n338 256.663
R1329 B.n588 B.n339 256.663
R1330 B.n588 B.n340 256.663
R1331 B.n588 B.n341 256.663
R1332 B.n588 B.n342 256.663
R1333 B.n588 B.n343 256.663
R1334 B.n588 B.n344 256.663
R1335 B.n588 B.n345 256.663
R1336 B.n588 B.n346 256.663
R1337 B.n588 B.n347 256.663
R1338 B.n588 B.n348 256.663
R1339 B.n588 B.n349 256.663
R1340 B.n588 B.n350 256.663
R1341 B.n588 B.n351 256.663
R1342 B.n588 B.n352 256.663
R1343 B.n588 B.n353 256.663
R1344 B.n588 B.n354 256.663
R1345 B.n588 B.n355 256.663
R1346 B.n588 B.n356 256.663
R1347 B.n588 B.n357 256.663
R1348 B.n588 B.n358 256.663
R1349 B.n588 B.n359 256.663
R1350 B.n588 B.n360 256.663
R1351 B.n588 B.n361 256.663
R1352 B.n588 B.n362 256.663
R1353 B.n588 B.n363 256.663
R1354 B.n588 B.n364 256.663
R1355 B.n588 B.n365 256.663
R1356 B.n588 B.n366 256.663
R1357 B.n588 B.n367 256.663
R1358 B.n588 B.n368 256.663
R1359 B.n588 B.n369 256.663
R1360 B.n588 B.n370 256.663
R1361 B.n588 B.n371 256.663
R1362 B.n588 B.n372 256.663
R1363 B.n588 B.n373 256.663
R1364 B.n588 B.n374 256.663
R1365 B.n588 B.n375 256.663
R1366 B.n588 B.n376 256.663
R1367 B.n588 B.n377 256.663
R1368 B.n588 B.n378 256.663
R1369 B.n588 B.n379 256.663
R1370 B.n588 B.n380 256.663
R1371 B.n588 B.n381 256.663
R1372 B.n588 B.n382 256.663
R1373 B.n588 B.n383 256.663
R1374 B.n588 B.n384 256.663
R1375 B.n595 B.n332 163.367
R1376 B.n595 B.n330 163.367
R1377 B.n599 B.n330 163.367
R1378 B.n599 B.n324 163.367
R1379 B.n607 B.n324 163.367
R1380 B.n607 B.n322 163.367
R1381 B.n611 B.n322 163.367
R1382 B.n611 B.n316 163.367
R1383 B.n619 B.n316 163.367
R1384 B.n619 B.n314 163.367
R1385 B.n623 B.n314 163.367
R1386 B.n623 B.n308 163.367
R1387 B.n631 B.n308 163.367
R1388 B.n631 B.n306 163.367
R1389 B.n635 B.n306 163.367
R1390 B.n635 B.n300 163.367
R1391 B.n644 B.n300 163.367
R1392 B.n644 B.n298 163.367
R1393 B.n648 B.n298 163.367
R1394 B.n648 B.n2 163.367
R1395 B.n726 B.n2 163.367
R1396 B.n726 B.n3 163.367
R1397 B.n722 B.n3 163.367
R1398 B.n722 B.n9 163.367
R1399 B.n718 B.n9 163.367
R1400 B.n718 B.n11 163.367
R1401 B.n714 B.n11 163.367
R1402 B.n714 B.n16 163.367
R1403 B.n710 B.n16 163.367
R1404 B.n710 B.n18 163.367
R1405 B.n706 B.n18 163.367
R1406 B.n706 B.n23 163.367
R1407 B.n702 B.n23 163.367
R1408 B.n702 B.n25 163.367
R1409 B.n698 B.n25 163.367
R1410 B.n698 B.n30 163.367
R1411 B.n694 B.n30 163.367
R1412 B.n694 B.n32 163.367
R1413 B.n690 B.n32 163.367
R1414 B.n690 B.n37 163.367
R1415 B.n686 B.n37 163.367
R1416 B.n686 B.n39 163.367
R1417 B.n386 B.n385 163.367
R1418 B.n581 B.n385 163.367
R1419 B.n579 B.n578 163.367
R1420 B.n575 B.n574 163.367
R1421 B.n571 B.n570 163.367
R1422 B.n567 B.n566 163.367
R1423 B.n563 B.n562 163.367
R1424 B.n559 B.n558 163.367
R1425 B.n555 B.n554 163.367
R1426 B.n551 B.n550 163.367
R1427 B.n547 B.n546 163.367
R1428 B.n543 B.n542 163.367
R1429 B.n539 B.n538 163.367
R1430 B.n535 B.n534 163.367
R1431 B.n531 B.n530 163.367
R1432 B.n527 B.n526 163.367
R1433 B.n523 B.n522 163.367
R1434 B.n519 B.n518 163.367
R1435 B.n515 B.n514 163.367
R1436 B.n511 B.n510 163.367
R1437 B.n507 B.n506 163.367
R1438 B.n503 B.n502 163.367
R1439 B.n499 B.n498 163.367
R1440 B.n495 B.n494 163.367
R1441 B.n491 B.n490 163.367
R1442 B.n487 B.n486 163.367
R1443 B.n483 B.n482 163.367
R1444 B.n479 B.n478 163.367
R1445 B.n475 B.n474 163.367
R1446 B.n471 B.n470 163.367
R1447 B.n467 B.n466 163.367
R1448 B.n463 B.n462 163.367
R1449 B.n459 B.n458 163.367
R1450 B.n455 B.n454 163.367
R1451 B.n451 B.n450 163.367
R1452 B.n447 B.n446 163.367
R1453 B.n443 B.n442 163.367
R1454 B.n439 B.n438 163.367
R1455 B.n435 B.n434 163.367
R1456 B.n431 B.n430 163.367
R1457 B.n427 B.n426 163.367
R1458 B.n423 B.n422 163.367
R1459 B.n419 B.n418 163.367
R1460 B.n415 B.n414 163.367
R1461 B.n411 B.n410 163.367
R1462 B.n407 B.n406 163.367
R1463 B.n403 B.n402 163.367
R1464 B.n399 B.n398 163.367
R1465 B.n395 B.n394 163.367
R1466 B.n589 B.n336 163.367
R1467 B.n593 B.n334 163.367
R1468 B.n593 B.n328 163.367
R1469 B.n601 B.n328 163.367
R1470 B.n601 B.n326 163.367
R1471 B.n605 B.n326 163.367
R1472 B.n605 B.n320 163.367
R1473 B.n613 B.n320 163.367
R1474 B.n613 B.n318 163.367
R1475 B.n617 B.n318 163.367
R1476 B.n617 B.n311 163.367
R1477 B.n625 B.n311 163.367
R1478 B.n625 B.n309 163.367
R1479 B.n629 B.n309 163.367
R1480 B.n629 B.n304 163.367
R1481 B.n637 B.n304 163.367
R1482 B.n637 B.n302 163.367
R1483 B.n642 B.n302 163.367
R1484 B.n642 B.n296 163.367
R1485 B.n650 B.n296 163.367
R1486 B.n651 B.n650 163.367
R1487 B.n651 B.n5 163.367
R1488 B.n6 B.n5 163.367
R1489 B.n7 B.n6 163.367
R1490 B.n656 B.n7 163.367
R1491 B.n656 B.n12 163.367
R1492 B.n13 B.n12 163.367
R1493 B.n14 B.n13 163.367
R1494 B.n661 B.n14 163.367
R1495 B.n661 B.n19 163.367
R1496 B.n20 B.n19 163.367
R1497 B.n21 B.n20 163.367
R1498 B.n666 B.n21 163.367
R1499 B.n666 B.n26 163.367
R1500 B.n27 B.n26 163.367
R1501 B.n28 B.n27 163.367
R1502 B.n671 B.n28 163.367
R1503 B.n671 B.n33 163.367
R1504 B.n34 B.n33 163.367
R1505 B.n35 B.n34 163.367
R1506 B.n676 B.n35 163.367
R1507 B.n676 B.n40 163.367
R1508 B.n41 B.n40 163.367
R1509 B.n100 B.n99 163.367
R1510 B.n104 B.n103 163.367
R1511 B.n108 B.n107 163.367
R1512 B.n112 B.n111 163.367
R1513 B.n116 B.n115 163.367
R1514 B.n120 B.n119 163.367
R1515 B.n124 B.n123 163.367
R1516 B.n128 B.n127 163.367
R1517 B.n132 B.n131 163.367
R1518 B.n136 B.n135 163.367
R1519 B.n140 B.n139 163.367
R1520 B.n144 B.n143 163.367
R1521 B.n148 B.n147 163.367
R1522 B.n152 B.n151 163.367
R1523 B.n156 B.n155 163.367
R1524 B.n160 B.n159 163.367
R1525 B.n164 B.n163 163.367
R1526 B.n168 B.n167 163.367
R1527 B.n172 B.n171 163.367
R1528 B.n176 B.n175 163.367
R1529 B.n180 B.n179 163.367
R1530 B.n184 B.n183 163.367
R1531 B.n189 B.n188 163.367
R1532 B.n193 B.n192 163.367
R1533 B.n197 B.n196 163.367
R1534 B.n201 B.n200 163.367
R1535 B.n205 B.n204 163.367
R1536 B.n210 B.n209 163.367
R1537 B.n214 B.n213 163.367
R1538 B.n218 B.n217 163.367
R1539 B.n222 B.n221 163.367
R1540 B.n226 B.n225 163.367
R1541 B.n230 B.n229 163.367
R1542 B.n234 B.n233 163.367
R1543 B.n238 B.n237 163.367
R1544 B.n242 B.n241 163.367
R1545 B.n246 B.n245 163.367
R1546 B.n250 B.n249 163.367
R1547 B.n254 B.n253 163.367
R1548 B.n258 B.n257 163.367
R1549 B.n262 B.n261 163.367
R1550 B.n266 B.n265 163.367
R1551 B.n270 B.n269 163.367
R1552 B.n274 B.n273 163.367
R1553 B.n278 B.n277 163.367
R1554 B.n282 B.n281 163.367
R1555 B.n286 B.n285 163.367
R1556 B.n290 B.n289 163.367
R1557 B.n292 B.n91 163.367
R1558 B.n588 B.n333 83.4549
R1559 B.n684 B.n683 83.4549
R1560 B.n587 B.n586 71.676
R1561 B.n581 B.n337 71.676
R1562 B.n578 B.n338 71.676
R1563 B.n574 B.n339 71.676
R1564 B.n570 B.n340 71.676
R1565 B.n566 B.n341 71.676
R1566 B.n562 B.n342 71.676
R1567 B.n558 B.n343 71.676
R1568 B.n554 B.n344 71.676
R1569 B.n550 B.n345 71.676
R1570 B.n546 B.n346 71.676
R1571 B.n542 B.n347 71.676
R1572 B.n538 B.n348 71.676
R1573 B.n534 B.n349 71.676
R1574 B.n530 B.n350 71.676
R1575 B.n526 B.n351 71.676
R1576 B.n522 B.n352 71.676
R1577 B.n518 B.n353 71.676
R1578 B.n514 B.n354 71.676
R1579 B.n510 B.n355 71.676
R1580 B.n506 B.n356 71.676
R1581 B.n502 B.n357 71.676
R1582 B.n498 B.n358 71.676
R1583 B.n494 B.n359 71.676
R1584 B.n490 B.n360 71.676
R1585 B.n486 B.n361 71.676
R1586 B.n482 B.n362 71.676
R1587 B.n478 B.n363 71.676
R1588 B.n474 B.n364 71.676
R1589 B.n470 B.n365 71.676
R1590 B.n466 B.n366 71.676
R1591 B.n462 B.n367 71.676
R1592 B.n458 B.n368 71.676
R1593 B.n454 B.n369 71.676
R1594 B.n450 B.n370 71.676
R1595 B.n446 B.n371 71.676
R1596 B.n442 B.n372 71.676
R1597 B.n438 B.n373 71.676
R1598 B.n434 B.n374 71.676
R1599 B.n430 B.n375 71.676
R1600 B.n426 B.n376 71.676
R1601 B.n422 B.n377 71.676
R1602 B.n418 B.n378 71.676
R1603 B.n414 B.n379 71.676
R1604 B.n410 B.n380 71.676
R1605 B.n406 B.n381 71.676
R1606 B.n402 B.n382 71.676
R1607 B.n398 B.n383 71.676
R1608 B.n394 B.n384 71.676
R1609 B.n96 B.n42 71.676
R1610 B.n100 B.n43 71.676
R1611 B.n104 B.n44 71.676
R1612 B.n108 B.n45 71.676
R1613 B.n112 B.n46 71.676
R1614 B.n116 B.n47 71.676
R1615 B.n120 B.n48 71.676
R1616 B.n124 B.n49 71.676
R1617 B.n128 B.n50 71.676
R1618 B.n132 B.n51 71.676
R1619 B.n136 B.n52 71.676
R1620 B.n140 B.n53 71.676
R1621 B.n144 B.n54 71.676
R1622 B.n148 B.n55 71.676
R1623 B.n152 B.n56 71.676
R1624 B.n156 B.n57 71.676
R1625 B.n160 B.n58 71.676
R1626 B.n164 B.n59 71.676
R1627 B.n168 B.n60 71.676
R1628 B.n172 B.n61 71.676
R1629 B.n176 B.n62 71.676
R1630 B.n180 B.n63 71.676
R1631 B.n184 B.n64 71.676
R1632 B.n189 B.n65 71.676
R1633 B.n193 B.n66 71.676
R1634 B.n197 B.n67 71.676
R1635 B.n201 B.n68 71.676
R1636 B.n205 B.n69 71.676
R1637 B.n210 B.n70 71.676
R1638 B.n214 B.n71 71.676
R1639 B.n218 B.n72 71.676
R1640 B.n222 B.n73 71.676
R1641 B.n226 B.n74 71.676
R1642 B.n230 B.n75 71.676
R1643 B.n234 B.n76 71.676
R1644 B.n238 B.n77 71.676
R1645 B.n242 B.n78 71.676
R1646 B.n246 B.n79 71.676
R1647 B.n250 B.n80 71.676
R1648 B.n254 B.n81 71.676
R1649 B.n258 B.n82 71.676
R1650 B.n262 B.n83 71.676
R1651 B.n266 B.n84 71.676
R1652 B.n270 B.n85 71.676
R1653 B.n274 B.n86 71.676
R1654 B.n278 B.n87 71.676
R1655 B.n282 B.n88 71.676
R1656 B.n286 B.n89 71.676
R1657 B.n290 B.n90 71.676
R1658 B.n682 B.n91 71.676
R1659 B.n682 B.n681 71.676
R1660 B.n292 B.n90 71.676
R1661 B.n289 B.n89 71.676
R1662 B.n285 B.n88 71.676
R1663 B.n281 B.n87 71.676
R1664 B.n277 B.n86 71.676
R1665 B.n273 B.n85 71.676
R1666 B.n269 B.n84 71.676
R1667 B.n265 B.n83 71.676
R1668 B.n261 B.n82 71.676
R1669 B.n257 B.n81 71.676
R1670 B.n253 B.n80 71.676
R1671 B.n249 B.n79 71.676
R1672 B.n245 B.n78 71.676
R1673 B.n241 B.n77 71.676
R1674 B.n237 B.n76 71.676
R1675 B.n233 B.n75 71.676
R1676 B.n229 B.n74 71.676
R1677 B.n225 B.n73 71.676
R1678 B.n221 B.n72 71.676
R1679 B.n217 B.n71 71.676
R1680 B.n213 B.n70 71.676
R1681 B.n209 B.n69 71.676
R1682 B.n204 B.n68 71.676
R1683 B.n200 B.n67 71.676
R1684 B.n196 B.n66 71.676
R1685 B.n192 B.n65 71.676
R1686 B.n188 B.n64 71.676
R1687 B.n183 B.n63 71.676
R1688 B.n179 B.n62 71.676
R1689 B.n175 B.n61 71.676
R1690 B.n171 B.n60 71.676
R1691 B.n167 B.n59 71.676
R1692 B.n163 B.n58 71.676
R1693 B.n159 B.n57 71.676
R1694 B.n155 B.n56 71.676
R1695 B.n151 B.n55 71.676
R1696 B.n147 B.n54 71.676
R1697 B.n143 B.n53 71.676
R1698 B.n139 B.n52 71.676
R1699 B.n135 B.n51 71.676
R1700 B.n131 B.n50 71.676
R1701 B.n127 B.n49 71.676
R1702 B.n123 B.n48 71.676
R1703 B.n119 B.n47 71.676
R1704 B.n115 B.n46 71.676
R1705 B.n111 B.n45 71.676
R1706 B.n107 B.n44 71.676
R1707 B.n103 B.n43 71.676
R1708 B.n99 B.n42 71.676
R1709 B.n587 B.n386 71.676
R1710 B.n579 B.n337 71.676
R1711 B.n575 B.n338 71.676
R1712 B.n571 B.n339 71.676
R1713 B.n567 B.n340 71.676
R1714 B.n563 B.n341 71.676
R1715 B.n559 B.n342 71.676
R1716 B.n555 B.n343 71.676
R1717 B.n551 B.n344 71.676
R1718 B.n547 B.n345 71.676
R1719 B.n543 B.n346 71.676
R1720 B.n539 B.n347 71.676
R1721 B.n535 B.n348 71.676
R1722 B.n531 B.n349 71.676
R1723 B.n527 B.n350 71.676
R1724 B.n523 B.n351 71.676
R1725 B.n519 B.n352 71.676
R1726 B.n515 B.n353 71.676
R1727 B.n511 B.n354 71.676
R1728 B.n507 B.n355 71.676
R1729 B.n503 B.n356 71.676
R1730 B.n499 B.n357 71.676
R1731 B.n495 B.n358 71.676
R1732 B.n491 B.n359 71.676
R1733 B.n487 B.n360 71.676
R1734 B.n483 B.n361 71.676
R1735 B.n479 B.n362 71.676
R1736 B.n475 B.n363 71.676
R1737 B.n471 B.n364 71.676
R1738 B.n467 B.n365 71.676
R1739 B.n463 B.n366 71.676
R1740 B.n459 B.n367 71.676
R1741 B.n455 B.n368 71.676
R1742 B.n451 B.n369 71.676
R1743 B.n447 B.n370 71.676
R1744 B.n443 B.n371 71.676
R1745 B.n439 B.n372 71.676
R1746 B.n435 B.n373 71.676
R1747 B.n431 B.n374 71.676
R1748 B.n427 B.n375 71.676
R1749 B.n423 B.n376 71.676
R1750 B.n419 B.n377 71.676
R1751 B.n415 B.n378 71.676
R1752 B.n411 B.n379 71.676
R1753 B.n407 B.n380 71.676
R1754 B.n403 B.n381 71.676
R1755 B.n399 B.n382 71.676
R1756 B.n395 B.n383 71.676
R1757 B.n384 B.n336 71.676
R1758 B.n392 B.n391 59.5399
R1759 B.n389 B.n388 59.5399
R1760 B.n186 B.n95 59.5399
R1761 B.n207 B.n93 59.5399
R1762 B.n594 B.n333 40.248
R1763 B.n594 B.n329 40.248
R1764 B.n600 B.n329 40.248
R1765 B.n600 B.n325 40.248
R1766 B.n606 B.n325 40.248
R1767 B.n612 B.n321 40.248
R1768 B.n612 B.n317 40.248
R1769 B.n618 B.n317 40.248
R1770 B.n618 B.n312 40.248
R1771 B.n624 B.n312 40.248
R1772 B.n624 B.n313 40.248
R1773 B.n630 B.n305 40.248
R1774 B.n636 B.n305 40.248
R1775 B.n636 B.n301 40.248
R1776 B.n643 B.n301 40.248
R1777 B.n649 B.n297 40.248
R1778 B.n649 B.n4 40.248
R1779 B.n725 B.n4 40.248
R1780 B.n725 B.n724 40.248
R1781 B.n724 B.n723 40.248
R1782 B.n723 B.n8 40.248
R1783 B.n717 B.n716 40.248
R1784 B.n716 B.n715 40.248
R1785 B.n715 B.n15 40.248
R1786 B.n709 B.n15 40.248
R1787 B.n708 B.n707 40.248
R1788 B.n707 B.n22 40.248
R1789 B.n701 B.n22 40.248
R1790 B.n701 B.n700 40.248
R1791 B.n700 B.n699 40.248
R1792 B.n699 B.n29 40.248
R1793 B.n693 B.n692 40.248
R1794 B.n692 B.n691 40.248
R1795 B.n691 B.n36 40.248
R1796 B.n685 B.n36 40.248
R1797 B.n685 B.n684 40.248
R1798 B.n97 B.n38 37.9322
R1799 B.n680 B.n679 37.9322
R1800 B.n591 B.n590 37.9322
R1801 B.n585 B.n331 37.9322
R1802 B.n313 B.t2 33.1455
R1803 B.t3 B.n708 33.1455
R1804 B.t1 B.n297 31.9618
R1805 B.t0 B.n8 31.9618
R1806 B.t5 B.n321 30.778
R1807 B.t12 B.n29 30.778
R1808 B.n391 B.n390 28.8975
R1809 B.n388 B.n387 28.8975
R1810 B.n95 B.n94 28.8975
R1811 B.n93 B.n92 28.8975
R1812 B B.n727 18.0485
R1813 B.n98 B.n97 10.6151
R1814 B.n101 B.n98 10.6151
R1815 B.n102 B.n101 10.6151
R1816 B.n105 B.n102 10.6151
R1817 B.n106 B.n105 10.6151
R1818 B.n109 B.n106 10.6151
R1819 B.n110 B.n109 10.6151
R1820 B.n113 B.n110 10.6151
R1821 B.n114 B.n113 10.6151
R1822 B.n117 B.n114 10.6151
R1823 B.n118 B.n117 10.6151
R1824 B.n121 B.n118 10.6151
R1825 B.n122 B.n121 10.6151
R1826 B.n125 B.n122 10.6151
R1827 B.n126 B.n125 10.6151
R1828 B.n129 B.n126 10.6151
R1829 B.n130 B.n129 10.6151
R1830 B.n133 B.n130 10.6151
R1831 B.n134 B.n133 10.6151
R1832 B.n137 B.n134 10.6151
R1833 B.n138 B.n137 10.6151
R1834 B.n141 B.n138 10.6151
R1835 B.n142 B.n141 10.6151
R1836 B.n145 B.n142 10.6151
R1837 B.n146 B.n145 10.6151
R1838 B.n149 B.n146 10.6151
R1839 B.n150 B.n149 10.6151
R1840 B.n153 B.n150 10.6151
R1841 B.n154 B.n153 10.6151
R1842 B.n157 B.n154 10.6151
R1843 B.n158 B.n157 10.6151
R1844 B.n161 B.n158 10.6151
R1845 B.n162 B.n161 10.6151
R1846 B.n165 B.n162 10.6151
R1847 B.n166 B.n165 10.6151
R1848 B.n169 B.n166 10.6151
R1849 B.n170 B.n169 10.6151
R1850 B.n173 B.n170 10.6151
R1851 B.n174 B.n173 10.6151
R1852 B.n177 B.n174 10.6151
R1853 B.n178 B.n177 10.6151
R1854 B.n181 B.n178 10.6151
R1855 B.n182 B.n181 10.6151
R1856 B.n185 B.n182 10.6151
R1857 B.n190 B.n187 10.6151
R1858 B.n191 B.n190 10.6151
R1859 B.n194 B.n191 10.6151
R1860 B.n195 B.n194 10.6151
R1861 B.n198 B.n195 10.6151
R1862 B.n199 B.n198 10.6151
R1863 B.n202 B.n199 10.6151
R1864 B.n203 B.n202 10.6151
R1865 B.n206 B.n203 10.6151
R1866 B.n211 B.n208 10.6151
R1867 B.n212 B.n211 10.6151
R1868 B.n215 B.n212 10.6151
R1869 B.n216 B.n215 10.6151
R1870 B.n219 B.n216 10.6151
R1871 B.n220 B.n219 10.6151
R1872 B.n223 B.n220 10.6151
R1873 B.n224 B.n223 10.6151
R1874 B.n227 B.n224 10.6151
R1875 B.n228 B.n227 10.6151
R1876 B.n231 B.n228 10.6151
R1877 B.n232 B.n231 10.6151
R1878 B.n235 B.n232 10.6151
R1879 B.n236 B.n235 10.6151
R1880 B.n239 B.n236 10.6151
R1881 B.n240 B.n239 10.6151
R1882 B.n243 B.n240 10.6151
R1883 B.n244 B.n243 10.6151
R1884 B.n247 B.n244 10.6151
R1885 B.n248 B.n247 10.6151
R1886 B.n251 B.n248 10.6151
R1887 B.n252 B.n251 10.6151
R1888 B.n255 B.n252 10.6151
R1889 B.n256 B.n255 10.6151
R1890 B.n259 B.n256 10.6151
R1891 B.n260 B.n259 10.6151
R1892 B.n263 B.n260 10.6151
R1893 B.n264 B.n263 10.6151
R1894 B.n267 B.n264 10.6151
R1895 B.n268 B.n267 10.6151
R1896 B.n271 B.n268 10.6151
R1897 B.n272 B.n271 10.6151
R1898 B.n275 B.n272 10.6151
R1899 B.n276 B.n275 10.6151
R1900 B.n279 B.n276 10.6151
R1901 B.n280 B.n279 10.6151
R1902 B.n283 B.n280 10.6151
R1903 B.n284 B.n283 10.6151
R1904 B.n287 B.n284 10.6151
R1905 B.n288 B.n287 10.6151
R1906 B.n291 B.n288 10.6151
R1907 B.n293 B.n291 10.6151
R1908 B.n294 B.n293 10.6151
R1909 B.n680 B.n294 10.6151
R1910 B.n592 B.n591 10.6151
R1911 B.n592 B.n327 10.6151
R1912 B.n602 B.n327 10.6151
R1913 B.n603 B.n602 10.6151
R1914 B.n604 B.n603 10.6151
R1915 B.n604 B.n319 10.6151
R1916 B.n614 B.n319 10.6151
R1917 B.n615 B.n614 10.6151
R1918 B.n616 B.n615 10.6151
R1919 B.n616 B.n310 10.6151
R1920 B.n626 B.n310 10.6151
R1921 B.n627 B.n626 10.6151
R1922 B.n628 B.n627 10.6151
R1923 B.n628 B.n303 10.6151
R1924 B.n638 B.n303 10.6151
R1925 B.n639 B.n638 10.6151
R1926 B.n641 B.n639 10.6151
R1927 B.n641 B.n640 10.6151
R1928 B.n640 B.n295 10.6151
R1929 B.n652 B.n295 10.6151
R1930 B.n653 B.n652 10.6151
R1931 B.n654 B.n653 10.6151
R1932 B.n655 B.n654 10.6151
R1933 B.n657 B.n655 10.6151
R1934 B.n658 B.n657 10.6151
R1935 B.n659 B.n658 10.6151
R1936 B.n660 B.n659 10.6151
R1937 B.n662 B.n660 10.6151
R1938 B.n663 B.n662 10.6151
R1939 B.n664 B.n663 10.6151
R1940 B.n665 B.n664 10.6151
R1941 B.n667 B.n665 10.6151
R1942 B.n668 B.n667 10.6151
R1943 B.n669 B.n668 10.6151
R1944 B.n670 B.n669 10.6151
R1945 B.n672 B.n670 10.6151
R1946 B.n673 B.n672 10.6151
R1947 B.n674 B.n673 10.6151
R1948 B.n675 B.n674 10.6151
R1949 B.n677 B.n675 10.6151
R1950 B.n678 B.n677 10.6151
R1951 B.n679 B.n678 10.6151
R1952 B.n585 B.n584 10.6151
R1953 B.n584 B.n583 10.6151
R1954 B.n583 B.n582 10.6151
R1955 B.n582 B.n580 10.6151
R1956 B.n580 B.n577 10.6151
R1957 B.n577 B.n576 10.6151
R1958 B.n576 B.n573 10.6151
R1959 B.n573 B.n572 10.6151
R1960 B.n572 B.n569 10.6151
R1961 B.n569 B.n568 10.6151
R1962 B.n568 B.n565 10.6151
R1963 B.n565 B.n564 10.6151
R1964 B.n564 B.n561 10.6151
R1965 B.n561 B.n560 10.6151
R1966 B.n560 B.n557 10.6151
R1967 B.n557 B.n556 10.6151
R1968 B.n556 B.n553 10.6151
R1969 B.n553 B.n552 10.6151
R1970 B.n552 B.n549 10.6151
R1971 B.n549 B.n548 10.6151
R1972 B.n548 B.n545 10.6151
R1973 B.n545 B.n544 10.6151
R1974 B.n544 B.n541 10.6151
R1975 B.n541 B.n540 10.6151
R1976 B.n540 B.n537 10.6151
R1977 B.n537 B.n536 10.6151
R1978 B.n536 B.n533 10.6151
R1979 B.n533 B.n532 10.6151
R1980 B.n532 B.n529 10.6151
R1981 B.n529 B.n528 10.6151
R1982 B.n528 B.n525 10.6151
R1983 B.n525 B.n524 10.6151
R1984 B.n524 B.n521 10.6151
R1985 B.n521 B.n520 10.6151
R1986 B.n520 B.n517 10.6151
R1987 B.n517 B.n516 10.6151
R1988 B.n516 B.n513 10.6151
R1989 B.n513 B.n512 10.6151
R1990 B.n512 B.n509 10.6151
R1991 B.n509 B.n508 10.6151
R1992 B.n508 B.n505 10.6151
R1993 B.n505 B.n504 10.6151
R1994 B.n504 B.n501 10.6151
R1995 B.n501 B.n500 10.6151
R1996 B.n497 B.n496 10.6151
R1997 B.n496 B.n493 10.6151
R1998 B.n493 B.n492 10.6151
R1999 B.n492 B.n489 10.6151
R2000 B.n489 B.n488 10.6151
R2001 B.n488 B.n485 10.6151
R2002 B.n485 B.n484 10.6151
R2003 B.n484 B.n481 10.6151
R2004 B.n481 B.n480 10.6151
R2005 B.n477 B.n476 10.6151
R2006 B.n476 B.n473 10.6151
R2007 B.n473 B.n472 10.6151
R2008 B.n472 B.n469 10.6151
R2009 B.n469 B.n468 10.6151
R2010 B.n468 B.n465 10.6151
R2011 B.n465 B.n464 10.6151
R2012 B.n464 B.n461 10.6151
R2013 B.n461 B.n460 10.6151
R2014 B.n460 B.n457 10.6151
R2015 B.n457 B.n456 10.6151
R2016 B.n456 B.n453 10.6151
R2017 B.n453 B.n452 10.6151
R2018 B.n452 B.n449 10.6151
R2019 B.n449 B.n448 10.6151
R2020 B.n448 B.n445 10.6151
R2021 B.n445 B.n444 10.6151
R2022 B.n444 B.n441 10.6151
R2023 B.n441 B.n440 10.6151
R2024 B.n440 B.n437 10.6151
R2025 B.n437 B.n436 10.6151
R2026 B.n436 B.n433 10.6151
R2027 B.n433 B.n432 10.6151
R2028 B.n432 B.n429 10.6151
R2029 B.n429 B.n428 10.6151
R2030 B.n428 B.n425 10.6151
R2031 B.n425 B.n424 10.6151
R2032 B.n424 B.n421 10.6151
R2033 B.n421 B.n420 10.6151
R2034 B.n420 B.n417 10.6151
R2035 B.n417 B.n416 10.6151
R2036 B.n416 B.n413 10.6151
R2037 B.n413 B.n412 10.6151
R2038 B.n412 B.n409 10.6151
R2039 B.n409 B.n408 10.6151
R2040 B.n408 B.n405 10.6151
R2041 B.n405 B.n404 10.6151
R2042 B.n404 B.n401 10.6151
R2043 B.n401 B.n400 10.6151
R2044 B.n400 B.n397 10.6151
R2045 B.n397 B.n396 10.6151
R2046 B.n396 B.n393 10.6151
R2047 B.n393 B.n335 10.6151
R2048 B.n590 B.n335 10.6151
R2049 B.n596 B.n331 10.6151
R2050 B.n597 B.n596 10.6151
R2051 B.n598 B.n597 10.6151
R2052 B.n598 B.n323 10.6151
R2053 B.n608 B.n323 10.6151
R2054 B.n609 B.n608 10.6151
R2055 B.n610 B.n609 10.6151
R2056 B.n610 B.n315 10.6151
R2057 B.n620 B.n315 10.6151
R2058 B.n621 B.n620 10.6151
R2059 B.n622 B.n621 10.6151
R2060 B.n622 B.n307 10.6151
R2061 B.n632 B.n307 10.6151
R2062 B.n633 B.n632 10.6151
R2063 B.n634 B.n633 10.6151
R2064 B.n634 B.n299 10.6151
R2065 B.n645 B.n299 10.6151
R2066 B.n646 B.n645 10.6151
R2067 B.n647 B.n646 10.6151
R2068 B.n647 B.n0 10.6151
R2069 B.n721 B.n1 10.6151
R2070 B.n721 B.n720 10.6151
R2071 B.n720 B.n719 10.6151
R2072 B.n719 B.n10 10.6151
R2073 B.n713 B.n10 10.6151
R2074 B.n713 B.n712 10.6151
R2075 B.n712 B.n711 10.6151
R2076 B.n711 B.n17 10.6151
R2077 B.n705 B.n17 10.6151
R2078 B.n705 B.n704 10.6151
R2079 B.n704 B.n703 10.6151
R2080 B.n703 B.n24 10.6151
R2081 B.n697 B.n24 10.6151
R2082 B.n697 B.n696 10.6151
R2083 B.n696 B.n695 10.6151
R2084 B.n695 B.n31 10.6151
R2085 B.n689 B.n31 10.6151
R2086 B.n689 B.n688 10.6151
R2087 B.n688 B.n687 10.6151
R2088 B.n687 B.n38 10.6151
R2089 B.n606 B.t5 9.4705
R2090 B.n693 B.t12 9.4705
R2091 B.n186 B.n185 9.36635
R2092 B.n208 B.n207 9.36635
R2093 B.n500 B.n389 9.36635
R2094 B.n477 B.n392 9.36635
R2095 B.n643 B.t1 8.28675
R2096 B.n717 B.t0 8.28675
R2097 B.n630 B.t2 7.103
R2098 B.n709 B.t3 7.103
R2099 B.n727 B.n0 2.81026
R2100 B.n727 B.n1 2.81026
R2101 B.n187 B.n186 1.24928
R2102 B.n207 B.n206 1.24928
R2103 B.n497 B.n389 1.24928
R2104 B.n480 B.n392 1.24928
R2105 VP.n2 VP.t2 312.007
R2106 VP.n2 VP.t1 311.791
R2107 VP.n3 VP.t0 276.527
R2108 VP.n9 VP.t3 276.527
R2109 VP.n4 VP.n3 173.779
R2110 VP.n10 VP.n9 173.779
R2111 VP.n8 VP.n0 161.3
R2112 VP.n7 VP.n6 161.3
R2113 VP.n5 VP.n1 161.3
R2114 VP.n4 VP.n2 61.4328
R2115 VP.n7 VP.n1 40.4934
R2116 VP.n8 VP.n7 40.4934
R2117 VP.n3 VP.n1 11.9893
R2118 VP.n9 VP.n8 11.9893
R2119 VP.n5 VP.n4 0.189894
R2120 VP.n6 VP.n5 0.189894
R2121 VP.n6 VP.n0 0.189894
R2122 VP.n10 VP.n0 0.189894
R2123 VP VP.n10 0.0516364
R2124 VDD1 VDD1.n1 102.82
R2125 VDD1 VDD1.n0 63.311
R2126 VDD1.n0 VDD1.t1 1.4881
R2127 VDD1.n0 VDD1.t2 1.4881
R2128 VDD1.n1 VDD1.t3 1.4881
R2129 VDD1.n1 VDD1.t0 1.4881
C0 VTAIL VN 3.88628f
C1 VDD1 VN 0.147511f
C2 VP VN 5.39961f
C3 VDD2 VN 4.25473f
C4 VDD1 VTAIL 6.26785f
C5 VTAIL VP 3.90038f
C6 VTAIL VDD2 6.3124f
C7 VDD1 VP 4.40933f
C8 VDD1 VDD2 0.674754f
C9 VP VDD2 0.302488f
C10 VDD2 B 3.059945f
C11 VDD1 B 6.91453f
C12 VTAIL B 9.904902f
C13 VN B 8.571321f
C14 VP B 5.963175f
C15 VDD1.t1 B 0.284693f
C16 VDD1.t2 B 0.284693f
C17 VDD1.n0 B 2.56116f
C18 VDD1.t3 B 0.284693f
C19 VDD1.t0 B 0.284693f
C20 VDD1.n1 B 3.22581f
C21 VP.n0 B 0.040455f
C22 VP.t3 B 1.70662f
C23 VP.n1 B 0.061418f
C24 VP.t2 B 1.79121f
C25 VP.t1 B 1.79066f
C26 VP.n2 B 2.67561f
C27 VP.t0 B 1.70662f
C28 VP.n3 B 0.684125f
C29 VP.n4 B 2.33502f
C30 VP.n5 B 0.040455f
C31 VP.n6 B 0.040455f
C32 VP.n7 B 0.032704f
C33 VP.n8 B 0.061418f
C34 VP.n9 B 0.684125f
C35 VP.n10 B 0.036257f
C36 VDD2.t0 B 0.284692f
C37 VDD2.t3 B 0.284692f
C38 VDD2.n0 B 3.19956f
C39 VDD2.t2 B 0.284692f
C40 VDD2.t1 B 0.284692f
C41 VDD2.n1 B 2.56083f
C42 VDD2.n2 B 3.58298f
C43 VTAIL.n0 B 0.021104f
C44 VTAIL.n1 B 0.015722f
C45 VTAIL.n2 B 0.008448f
C46 VTAIL.n3 B 0.019969f
C47 VTAIL.n4 B 0.008945f
C48 VTAIL.n5 B 0.015722f
C49 VTAIL.n6 B 0.008448f
C50 VTAIL.n7 B 0.019969f
C51 VTAIL.n8 B 0.008945f
C52 VTAIL.n9 B 0.015722f
C53 VTAIL.n10 B 0.008448f
C54 VTAIL.n11 B 0.019969f
C55 VTAIL.n12 B 0.008945f
C56 VTAIL.n13 B 0.015722f
C57 VTAIL.n14 B 0.008448f
C58 VTAIL.n15 B 0.019969f
C59 VTAIL.n16 B 0.008945f
C60 VTAIL.n17 B 0.015722f
C61 VTAIL.n18 B 0.008448f
C62 VTAIL.n19 B 0.019969f
C63 VTAIL.n20 B 0.008945f
C64 VTAIL.n21 B 0.901119f
C65 VTAIL.n22 B 0.008448f
C66 VTAIL.t1 B 0.032835f
C67 VTAIL.n23 B 0.09588f
C68 VTAIL.n24 B 0.011796f
C69 VTAIL.n25 B 0.014977f
C70 VTAIL.n26 B 0.019969f
C71 VTAIL.n27 B 0.008945f
C72 VTAIL.n28 B 0.008448f
C73 VTAIL.n29 B 0.015722f
C74 VTAIL.n30 B 0.015722f
C75 VTAIL.n31 B 0.008448f
C76 VTAIL.n32 B 0.008945f
C77 VTAIL.n33 B 0.019969f
C78 VTAIL.n34 B 0.019969f
C79 VTAIL.n35 B 0.008945f
C80 VTAIL.n36 B 0.008448f
C81 VTAIL.n37 B 0.015722f
C82 VTAIL.n38 B 0.015722f
C83 VTAIL.n39 B 0.008448f
C84 VTAIL.n40 B 0.008945f
C85 VTAIL.n41 B 0.019969f
C86 VTAIL.n42 B 0.019969f
C87 VTAIL.n43 B 0.008945f
C88 VTAIL.n44 B 0.008448f
C89 VTAIL.n45 B 0.015722f
C90 VTAIL.n46 B 0.015722f
C91 VTAIL.n47 B 0.008448f
C92 VTAIL.n48 B 0.008945f
C93 VTAIL.n49 B 0.019969f
C94 VTAIL.n50 B 0.019969f
C95 VTAIL.n51 B 0.008945f
C96 VTAIL.n52 B 0.008448f
C97 VTAIL.n53 B 0.015722f
C98 VTAIL.n54 B 0.015722f
C99 VTAIL.n55 B 0.008448f
C100 VTAIL.n56 B 0.008945f
C101 VTAIL.n57 B 0.019969f
C102 VTAIL.n58 B 0.019969f
C103 VTAIL.n59 B 0.008945f
C104 VTAIL.n60 B 0.008448f
C105 VTAIL.n61 B 0.015722f
C106 VTAIL.n62 B 0.015722f
C107 VTAIL.n63 B 0.008448f
C108 VTAIL.n64 B 0.008945f
C109 VTAIL.n65 B 0.019969f
C110 VTAIL.n66 B 0.040476f
C111 VTAIL.n67 B 0.008945f
C112 VTAIL.n68 B 0.016519f
C113 VTAIL.n69 B 0.038703f
C114 VTAIL.n70 B 0.041247f
C115 VTAIL.n71 B 0.074048f
C116 VTAIL.n72 B 0.021104f
C117 VTAIL.n73 B 0.015722f
C118 VTAIL.n74 B 0.008448f
C119 VTAIL.n75 B 0.019969f
C120 VTAIL.n76 B 0.008945f
C121 VTAIL.n77 B 0.015722f
C122 VTAIL.n78 B 0.008448f
C123 VTAIL.n79 B 0.019969f
C124 VTAIL.n80 B 0.008945f
C125 VTAIL.n81 B 0.015722f
C126 VTAIL.n82 B 0.008448f
C127 VTAIL.n83 B 0.019969f
C128 VTAIL.n84 B 0.008945f
C129 VTAIL.n85 B 0.015722f
C130 VTAIL.n86 B 0.008448f
C131 VTAIL.n87 B 0.019969f
C132 VTAIL.n88 B 0.008945f
C133 VTAIL.n89 B 0.015722f
C134 VTAIL.n90 B 0.008448f
C135 VTAIL.n91 B 0.019969f
C136 VTAIL.n92 B 0.008945f
C137 VTAIL.n93 B 0.901119f
C138 VTAIL.n94 B 0.008448f
C139 VTAIL.t5 B 0.032835f
C140 VTAIL.n95 B 0.09588f
C141 VTAIL.n96 B 0.011796f
C142 VTAIL.n97 B 0.014977f
C143 VTAIL.n98 B 0.019969f
C144 VTAIL.n99 B 0.008945f
C145 VTAIL.n100 B 0.008448f
C146 VTAIL.n101 B 0.015722f
C147 VTAIL.n102 B 0.015722f
C148 VTAIL.n103 B 0.008448f
C149 VTAIL.n104 B 0.008945f
C150 VTAIL.n105 B 0.019969f
C151 VTAIL.n106 B 0.019969f
C152 VTAIL.n107 B 0.008945f
C153 VTAIL.n108 B 0.008448f
C154 VTAIL.n109 B 0.015722f
C155 VTAIL.n110 B 0.015722f
C156 VTAIL.n111 B 0.008448f
C157 VTAIL.n112 B 0.008945f
C158 VTAIL.n113 B 0.019969f
C159 VTAIL.n114 B 0.019969f
C160 VTAIL.n115 B 0.008945f
C161 VTAIL.n116 B 0.008448f
C162 VTAIL.n117 B 0.015722f
C163 VTAIL.n118 B 0.015722f
C164 VTAIL.n119 B 0.008448f
C165 VTAIL.n120 B 0.008945f
C166 VTAIL.n121 B 0.019969f
C167 VTAIL.n122 B 0.019969f
C168 VTAIL.n123 B 0.008945f
C169 VTAIL.n124 B 0.008448f
C170 VTAIL.n125 B 0.015722f
C171 VTAIL.n126 B 0.015722f
C172 VTAIL.n127 B 0.008448f
C173 VTAIL.n128 B 0.008945f
C174 VTAIL.n129 B 0.019969f
C175 VTAIL.n130 B 0.019969f
C176 VTAIL.n131 B 0.008945f
C177 VTAIL.n132 B 0.008448f
C178 VTAIL.n133 B 0.015722f
C179 VTAIL.n134 B 0.015722f
C180 VTAIL.n135 B 0.008448f
C181 VTAIL.n136 B 0.008945f
C182 VTAIL.n137 B 0.019969f
C183 VTAIL.n138 B 0.040476f
C184 VTAIL.n139 B 0.008945f
C185 VTAIL.n140 B 0.016519f
C186 VTAIL.n141 B 0.038703f
C187 VTAIL.n142 B 0.041247f
C188 VTAIL.n143 B 0.103636f
C189 VTAIL.n144 B 0.021104f
C190 VTAIL.n145 B 0.015722f
C191 VTAIL.n146 B 0.008448f
C192 VTAIL.n147 B 0.019969f
C193 VTAIL.n148 B 0.008945f
C194 VTAIL.n149 B 0.015722f
C195 VTAIL.n150 B 0.008448f
C196 VTAIL.n151 B 0.019969f
C197 VTAIL.n152 B 0.008945f
C198 VTAIL.n153 B 0.015722f
C199 VTAIL.n154 B 0.008448f
C200 VTAIL.n155 B 0.019969f
C201 VTAIL.n156 B 0.008945f
C202 VTAIL.n157 B 0.015722f
C203 VTAIL.n158 B 0.008448f
C204 VTAIL.n159 B 0.019969f
C205 VTAIL.n160 B 0.008945f
C206 VTAIL.n161 B 0.015722f
C207 VTAIL.n162 B 0.008448f
C208 VTAIL.n163 B 0.019969f
C209 VTAIL.n164 B 0.008945f
C210 VTAIL.n165 B 0.901119f
C211 VTAIL.n166 B 0.008448f
C212 VTAIL.t4 B 0.032835f
C213 VTAIL.n167 B 0.09588f
C214 VTAIL.n168 B 0.011796f
C215 VTAIL.n169 B 0.014977f
C216 VTAIL.n170 B 0.019969f
C217 VTAIL.n171 B 0.008945f
C218 VTAIL.n172 B 0.008448f
C219 VTAIL.n173 B 0.015722f
C220 VTAIL.n174 B 0.015722f
C221 VTAIL.n175 B 0.008448f
C222 VTAIL.n176 B 0.008945f
C223 VTAIL.n177 B 0.019969f
C224 VTAIL.n178 B 0.019969f
C225 VTAIL.n179 B 0.008945f
C226 VTAIL.n180 B 0.008448f
C227 VTAIL.n181 B 0.015722f
C228 VTAIL.n182 B 0.015722f
C229 VTAIL.n183 B 0.008448f
C230 VTAIL.n184 B 0.008945f
C231 VTAIL.n185 B 0.019969f
C232 VTAIL.n186 B 0.019969f
C233 VTAIL.n187 B 0.008945f
C234 VTAIL.n188 B 0.008448f
C235 VTAIL.n189 B 0.015722f
C236 VTAIL.n190 B 0.015722f
C237 VTAIL.n191 B 0.008448f
C238 VTAIL.n192 B 0.008945f
C239 VTAIL.n193 B 0.019969f
C240 VTAIL.n194 B 0.019969f
C241 VTAIL.n195 B 0.008945f
C242 VTAIL.n196 B 0.008448f
C243 VTAIL.n197 B 0.015722f
C244 VTAIL.n198 B 0.015722f
C245 VTAIL.n199 B 0.008448f
C246 VTAIL.n200 B 0.008945f
C247 VTAIL.n201 B 0.019969f
C248 VTAIL.n202 B 0.019969f
C249 VTAIL.n203 B 0.008945f
C250 VTAIL.n204 B 0.008448f
C251 VTAIL.n205 B 0.015722f
C252 VTAIL.n206 B 0.015722f
C253 VTAIL.n207 B 0.008448f
C254 VTAIL.n208 B 0.008945f
C255 VTAIL.n209 B 0.019969f
C256 VTAIL.n210 B 0.040476f
C257 VTAIL.n211 B 0.008945f
C258 VTAIL.n212 B 0.016519f
C259 VTAIL.n213 B 0.038703f
C260 VTAIL.n214 B 0.041247f
C261 VTAIL.n215 B 0.939743f
C262 VTAIL.n216 B 0.021104f
C263 VTAIL.n217 B 0.015722f
C264 VTAIL.n218 B 0.008448f
C265 VTAIL.n219 B 0.019969f
C266 VTAIL.n220 B 0.008945f
C267 VTAIL.n221 B 0.015722f
C268 VTAIL.n222 B 0.008448f
C269 VTAIL.n223 B 0.019969f
C270 VTAIL.n224 B 0.008945f
C271 VTAIL.n225 B 0.015722f
C272 VTAIL.n226 B 0.008448f
C273 VTAIL.n227 B 0.019969f
C274 VTAIL.n228 B 0.008945f
C275 VTAIL.n229 B 0.015722f
C276 VTAIL.n230 B 0.008448f
C277 VTAIL.n231 B 0.019969f
C278 VTAIL.n232 B 0.008945f
C279 VTAIL.n233 B 0.015722f
C280 VTAIL.n234 B 0.008448f
C281 VTAIL.n235 B 0.019969f
C282 VTAIL.n236 B 0.008945f
C283 VTAIL.n237 B 0.901119f
C284 VTAIL.n238 B 0.008448f
C285 VTAIL.t2 B 0.032835f
C286 VTAIL.n239 B 0.09588f
C287 VTAIL.n240 B 0.011796f
C288 VTAIL.n241 B 0.014977f
C289 VTAIL.n242 B 0.019969f
C290 VTAIL.n243 B 0.008945f
C291 VTAIL.n244 B 0.008448f
C292 VTAIL.n245 B 0.015722f
C293 VTAIL.n246 B 0.015722f
C294 VTAIL.n247 B 0.008448f
C295 VTAIL.n248 B 0.008945f
C296 VTAIL.n249 B 0.019969f
C297 VTAIL.n250 B 0.019969f
C298 VTAIL.n251 B 0.008945f
C299 VTAIL.n252 B 0.008448f
C300 VTAIL.n253 B 0.015722f
C301 VTAIL.n254 B 0.015722f
C302 VTAIL.n255 B 0.008448f
C303 VTAIL.n256 B 0.008945f
C304 VTAIL.n257 B 0.019969f
C305 VTAIL.n258 B 0.019969f
C306 VTAIL.n259 B 0.008945f
C307 VTAIL.n260 B 0.008448f
C308 VTAIL.n261 B 0.015722f
C309 VTAIL.n262 B 0.015722f
C310 VTAIL.n263 B 0.008448f
C311 VTAIL.n264 B 0.008945f
C312 VTAIL.n265 B 0.019969f
C313 VTAIL.n266 B 0.019969f
C314 VTAIL.n267 B 0.008945f
C315 VTAIL.n268 B 0.008448f
C316 VTAIL.n269 B 0.015722f
C317 VTAIL.n270 B 0.015722f
C318 VTAIL.n271 B 0.008448f
C319 VTAIL.n272 B 0.008945f
C320 VTAIL.n273 B 0.019969f
C321 VTAIL.n274 B 0.019969f
C322 VTAIL.n275 B 0.008945f
C323 VTAIL.n276 B 0.008448f
C324 VTAIL.n277 B 0.015722f
C325 VTAIL.n278 B 0.015722f
C326 VTAIL.n279 B 0.008448f
C327 VTAIL.n280 B 0.008945f
C328 VTAIL.n281 B 0.019969f
C329 VTAIL.n282 B 0.040476f
C330 VTAIL.n283 B 0.008945f
C331 VTAIL.n284 B 0.016519f
C332 VTAIL.n285 B 0.038703f
C333 VTAIL.n286 B 0.041247f
C334 VTAIL.n287 B 0.939743f
C335 VTAIL.n288 B 0.021104f
C336 VTAIL.n289 B 0.015722f
C337 VTAIL.n290 B 0.008448f
C338 VTAIL.n291 B 0.019969f
C339 VTAIL.n292 B 0.008945f
C340 VTAIL.n293 B 0.015722f
C341 VTAIL.n294 B 0.008448f
C342 VTAIL.n295 B 0.019969f
C343 VTAIL.n296 B 0.008945f
C344 VTAIL.n297 B 0.015722f
C345 VTAIL.n298 B 0.008448f
C346 VTAIL.n299 B 0.019969f
C347 VTAIL.n300 B 0.008945f
C348 VTAIL.n301 B 0.015722f
C349 VTAIL.n302 B 0.008448f
C350 VTAIL.n303 B 0.019969f
C351 VTAIL.n304 B 0.008945f
C352 VTAIL.n305 B 0.015722f
C353 VTAIL.n306 B 0.008448f
C354 VTAIL.n307 B 0.019969f
C355 VTAIL.n308 B 0.008945f
C356 VTAIL.n309 B 0.901119f
C357 VTAIL.n310 B 0.008448f
C358 VTAIL.t3 B 0.032835f
C359 VTAIL.n311 B 0.09588f
C360 VTAIL.n312 B 0.011796f
C361 VTAIL.n313 B 0.014977f
C362 VTAIL.n314 B 0.019969f
C363 VTAIL.n315 B 0.008945f
C364 VTAIL.n316 B 0.008448f
C365 VTAIL.n317 B 0.015722f
C366 VTAIL.n318 B 0.015722f
C367 VTAIL.n319 B 0.008448f
C368 VTAIL.n320 B 0.008945f
C369 VTAIL.n321 B 0.019969f
C370 VTAIL.n322 B 0.019969f
C371 VTAIL.n323 B 0.008945f
C372 VTAIL.n324 B 0.008448f
C373 VTAIL.n325 B 0.015722f
C374 VTAIL.n326 B 0.015722f
C375 VTAIL.n327 B 0.008448f
C376 VTAIL.n328 B 0.008945f
C377 VTAIL.n329 B 0.019969f
C378 VTAIL.n330 B 0.019969f
C379 VTAIL.n331 B 0.008945f
C380 VTAIL.n332 B 0.008448f
C381 VTAIL.n333 B 0.015722f
C382 VTAIL.n334 B 0.015722f
C383 VTAIL.n335 B 0.008448f
C384 VTAIL.n336 B 0.008945f
C385 VTAIL.n337 B 0.019969f
C386 VTAIL.n338 B 0.019969f
C387 VTAIL.n339 B 0.008945f
C388 VTAIL.n340 B 0.008448f
C389 VTAIL.n341 B 0.015722f
C390 VTAIL.n342 B 0.015722f
C391 VTAIL.n343 B 0.008448f
C392 VTAIL.n344 B 0.008945f
C393 VTAIL.n345 B 0.019969f
C394 VTAIL.n346 B 0.019969f
C395 VTAIL.n347 B 0.008945f
C396 VTAIL.n348 B 0.008448f
C397 VTAIL.n349 B 0.015722f
C398 VTAIL.n350 B 0.015722f
C399 VTAIL.n351 B 0.008448f
C400 VTAIL.n352 B 0.008945f
C401 VTAIL.n353 B 0.019969f
C402 VTAIL.n354 B 0.040476f
C403 VTAIL.n355 B 0.008945f
C404 VTAIL.n356 B 0.016519f
C405 VTAIL.n357 B 0.038703f
C406 VTAIL.n358 B 0.041247f
C407 VTAIL.n359 B 0.103636f
C408 VTAIL.n360 B 0.021104f
C409 VTAIL.n361 B 0.015722f
C410 VTAIL.n362 B 0.008448f
C411 VTAIL.n363 B 0.019969f
C412 VTAIL.n364 B 0.008945f
C413 VTAIL.n365 B 0.015722f
C414 VTAIL.n366 B 0.008448f
C415 VTAIL.n367 B 0.019969f
C416 VTAIL.n368 B 0.008945f
C417 VTAIL.n369 B 0.015722f
C418 VTAIL.n370 B 0.008448f
C419 VTAIL.n371 B 0.019969f
C420 VTAIL.n372 B 0.008945f
C421 VTAIL.n373 B 0.015722f
C422 VTAIL.n374 B 0.008448f
C423 VTAIL.n375 B 0.019969f
C424 VTAIL.n376 B 0.008945f
C425 VTAIL.n377 B 0.015722f
C426 VTAIL.n378 B 0.008448f
C427 VTAIL.n379 B 0.019969f
C428 VTAIL.n380 B 0.008945f
C429 VTAIL.n381 B 0.901119f
C430 VTAIL.n382 B 0.008448f
C431 VTAIL.t6 B 0.032835f
C432 VTAIL.n383 B 0.09588f
C433 VTAIL.n384 B 0.011796f
C434 VTAIL.n385 B 0.014977f
C435 VTAIL.n386 B 0.019969f
C436 VTAIL.n387 B 0.008945f
C437 VTAIL.n388 B 0.008448f
C438 VTAIL.n389 B 0.015722f
C439 VTAIL.n390 B 0.015722f
C440 VTAIL.n391 B 0.008448f
C441 VTAIL.n392 B 0.008945f
C442 VTAIL.n393 B 0.019969f
C443 VTAIL.n394 B 0.019969f
C444 VTAIL.n395 B 0.008945f
C445 VTAIL.n396 B 0.008448f
C446 VTAIL.n397 B 0.015722f
C447 VTAIL.n398 B 0.015722f
C448 VTAIL.n399 B 0.008448f
C449 VTAIL.n400 B 0.008945f
C450 VTAIL.n401 B 0.019969f
C451 VTAIL.n402 B 0.019969f
C452 VTAIL.n403 B 0.008945f
C453 VTAIL.n404 B 0.008448f
C454 VTAIL.n405 B 0.015722f
C455 VTAIL.n406 B 0.015722f
C456 VTAIL.n407 B 0.008448f
C457 VTAIL.n408 B 0.008945f
C458 VTAIL.n409 B 0.019969f
C459 VTAIL.n410 B 0.019969f
C460 VTAIL.n411 B 0.008945f
C461 VTAIL.n412 B 0.008448f
C462 VTAIL.n413 B 0.015722f
C463 VTAIL.n414 B 0.015722f
C464 VTAIL.n415 B 0.008448f
C465 VTAIL.n416 B 0.008945f
C466 VTAIL.n417 B 0.019969f
C467 VTAIL.n418 B 0.019969f
C468 VTAIL.n419 B 0.008945f
C469 VTAIL.n420 B 0.008448f
C470 VTAIL.n421 B 0.015722f
C471 VTAIL.n422 B 0.015722f
C472 VTAIL.n423 B 0.008448f
C473 VTAIL.n424 B 0.008945f
C474 VTAIL.n425 B 0.019969f
C475 VTAIL.n426 B 0.040476f
C476 VTAIL.n427 B 0.008945f
C477 VTAIL.n428 B 0.016519f
C478 VTAIL.n429 B 0.038703f
C479 VTAIL.n430 B 0.041247f
C480 VTAIL.n431 B 0.103636f
C481 VTAIL.n432 B 0.021104f
C482 VTAIL.n433 B 0.015722f
C483 VTAIL.n434 B 0.008448f
C484 VTAIL.n435 B 0.019969f
C485 VTAIL.n436 B 0.008945f
C486 VTAIL.n437 B 0.015722f
C487 VTAIL.n438 B 0.008448f
C488 VTAIL.n439 B 0.019969f
C489 VTAIL.n440 B 0.008945f
C490 VTAIL.n441 B 0.015722f
C491 VTAIL.n442 B 0.008448f
C492 VTAIL.n443 B 0.019969f
C493 VTAIL.n444 B 0.008945f
C494 VTAIL.n445 B 0.015722f
C495 VTAIL.n446 B 0.008448f
C496 VTAIL.n447 B 0.019969f
C497 VTAIL.n448 B 0.008945f
C498 VTAIL.n449 B 0.015722f
C499 VTAIL.n450 B 0.008448f
C500 VTAIL.n451 B 0.019969f
C501 VTAIL.n452 B 0.008945f
C502 VTAIL.n453 B 0.901119f
C503 VTAIL.n454 B 0.008448f
C504 VTAIL.t7 B 0.032835f
C505 VTAIL.n455 B 0.09588f
C506 VTAIL.n456 B 0.011796f
C507 VTAIL.n457 B 0.014977f
C508 VTAIL.n458 B 0.019969f
C509 VTAIL.n459 B 0.008945f
C510 VTAIL.n460 B 0.008448f
C511 VTAIL.n461 B 0.015722f
C512 VTAIL.n462 B 0.015722f
C513 VTAIL.n463 B 0.008448f
C514 VTAIL.n464 B 0.008945f
C515 VTAIL.n465 B 0.019969f
C516 VTAIL.n466 B 0.019969f
C517 VTAIL.n467 B 0.008945f
C518 VTAIL.n468 B 0.008448f
C519 VTAIL.n469 B 0.015722f
C520 VTAIL.n470 B 0.015722f
C521 VTAIL.n471 B 0.008448f
C522 VTAIL.n472 B 0.008945f
C523 VTAIL.n473 B 0.019969f
C524 VTAIL.n474 B 0.019969f
C525 VTAIL.n475 B 0.008945f
C526 VTAIL.n476 B 0.008448f
C527 VTAIL.n477 B 0.015722f
C528 VTAIL.n478 B 0.015722f
C529 VTAIL.n479 B 0.008448f
C530 VTAIL.n480 B 0.008945f
C531 VTAIL.n481 B 0.019969f
C532 VTAIL.n482 B 0.019969f
C533 VTAIL.n483 B 0.008945f
C534 VTAIL.n484 B 0.008448f
C535 VTAIL.n485 B 0.015722f
C536 VTAIL.n486 B 0.015722f
C537 VTAIL.n487 B 0.008448f
C538 VTAIL.n488 B 0.008945f
C539 VTAIL.n489 B 0.019969f
C540 VTAIL.n490 B 0.019969f
C541 VTAIL.n491 B 0.008945f
C542 VTAIL.n492 B 0.008448f
C543 VTAIL.n493 B 0.015722f
C544 VTAIL.n494 B 0.015722f
C545 VTAIL.n495 B 0.008448f
C546 VTAIL.n496 B 0.008945f
C547 VTAIL.n497 B 0.019969f
C548 VTAIL.n498 B 0.040476f
C549 VTAIL.n499 B 0.008945f
C550 VTAIL.n500 B 0.016519f
C551 VTAIL.n501 B 0.038703f
C552 VTAIL.n502 B 0.041247f
C553 VTAIL.n503 B 0.939743f
C554 VTAIL.n504 B 0.021104f
C555 VTAIL.n505 B 0.015722f
C556 VTAIL.n506 B 0.008448f
C557 VTAIL.n507 B 0.019969f
C558 VTAIL.n508 B 0.008945f
C559 VTAIL.n509 B 0.015722f
C560 VTAIL.n510 B 0.008448f
C561 VTAIL.n511 B 0.019969f
C562 VTAIL.n512 B 0.008945f
C563 VTAIL.n513 B 0.015722f
C564 VTAIL.n514 B 0.008448f
C565 VTAIL.n515 B 0.019969f
C566 VTAIL.n516 B 0.008945f
C567 VTAIL.n517 B 0.015722f
C568 VTAIL.n518 B 0.008448f
C569 VTAIL.n519 B 0.019969f
C570 VTAIL.n520 B 0.008945f
C571 VTAIL.n521 B 0.015722f
C572 VTAIL.n522 B 0.008448f
C573 VTAIL.n523 B 0.019969f
C574 VTAIL.n524 B 0.008945f
C575 VTAIL.n525 B 0.901119f
C576 VTAIL.n526 B 0.008448f
C577 VTAIL.t0 B 0.032835f
C578 VTAIL.n527 B 0.09588f
C579 VTAIL.n528 B 0.011796f
C580 VTAIL.n529 B 0.014977f
C581 VTAIL.n530 B 0.019969f
C582 VTAIL.n531 B 0.008945f
C583 VTAIL.n532 B 0.008448f
C584 VTAIL.n533 B 0.015722f
C585 VTAIL.n534 B 0.015722f
C586 VTAIL.n535 B 0.008448f
C587 VTAIL.n536 B 0.008945f
C588 VTAIL.n537 B 0.019969f
C589 VTAIL.n538 B 0.019969f
C590 VTAIL.n539 B 0.008945f
C591 VTAIL.n540 B 0.008448f
C592 VTAIL.n541 B 0.015722f
C593 VTAIL.n542 B 0.015722f
C594 VTAIL.n543 B 0.008448f
C595 VTAIL.n544 B 0.008945f
C596 VTAIL.n545 B 0.019969f
C597 VTAIL.n546 B 0.019969f
C598 VTAIL.n547 B 0.008945f
C599 VTAIL.n548 B 0.008448f
C600 VTAIL.n549 B 0.015722f
C601 VTAIL.n550 B 0.015722f
C602 VTAIL.n551 B 0.008448f
C603 VTAIL.n552 B 0.008945f
C604 VTAIL.n553 B 0.019969f
C605 VTAIL.n554 B 0.019969f
C606 VTAIL.n555 B 0.008945f
C607 VTAIL.n556 B 0.008448f
C608 VTAIL.n557 B 0.015722f
C609 VTAIL.n558 B 0.015722f
C610 VTAIL.n559 B 0.008448f
C611 VTAIL.n560 B 0.008945f
C612 VTAIL.n561 B 0.019969f
C613 VTAIL.n562 B 0.019969f
C614 VTAIL.n563 B 0.008945f
C615 VTAIL.n564 B 0.008448f
C616 VTAIL.n565 B 0.015722f
C617 VTAIL.n566 B 0.015722f
C618 VTAIL.n567 B 0.008448f
C619 VTAIL.n568 B 0.008945f
C620 VTAIL.n569 B 0.019969f
C621 VTAIL.n570 B 0.040476f
C622 VTAIL.n571 B 0.008945f
C623 VTAIL.n572 B 0.016519f
C624 VTAIL.n573 B 0.038703f
C625 VTAIL.n574 B 0.041247f
C626 VTAIL.n575 B 0.90426f
C627 VN.t3 B 1.77078f
C628 VN.t0 B 1.77024f
C629 VN.n0 B 1.34223f
C630 VN.t2 B 1.77078f
C631 VN.t1 B 1.77024f
C632 VN.n1 B 2.66691f
.ends

