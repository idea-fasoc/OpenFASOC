* NGSPICE file created from diff_pair_sample_1507.ext - technology: sky130A

.subckt diff_pair_sample_1507 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t6 w_n2032_n1696# sky130_fd_pr__pfet_01v8 ad=0.6006 pd=3.97 as=1.4196 ps=8.06 w=3.64 l=1.44
X1 B.t11 B.t9 B.t10 w_n2032_n1696# sky130_fd_pr__pfet_01v8 ad=1.4196 pd=8.06 as=0 ps=0 w=3.64 l=1.44
X2 VTAIL.t1 VN.t0 VDD2.t3 w_n2032_n1696# sky130_fd_pr__pfet_01v8 ad=1.4196 pd=8.06 as=0.6006 ps=3.97 w=3.64 l=1.44
X3 VDD2.t2 VN.t1 VTAIL.t2 w_n2032_n1696# sky130_fd_pr__pfet_01v8 ad=0.6006 pd=3.97 as=1.4196 ps=8.06 w=3.64 l=1.44
X4 VTAIL.t7 VP.t1 VDD1.t2 w_n2032_n1696# sky130_fd_pr__pfet_01v8 ad=1.4196 pd=8.06 as=0.6006 ps=3.97 w=3.64 l=1.44
X5 VTAIL.t4 VP.t2 VDD1.t1 w_n2032_n1696# sky130_fd_pr__pfet_01v8 ad=1.4196 pd=8.06 as=0.6006 ps=3.97 w=3.64 l=1.44
X6 B.t8 B.t6 B.t7 w_n2032_n1696# sky130_fd_pr__pfet_01v8 ad=1.4196 pd=8.06 as=0 ps=0 w=3.64 l=1.44
X7 VDD2.t1 VN.t2 VTAIL.t0 w_n2032_n1696# sky130_fd_pr__pfet_01v8 ad=0.6006 pd=3.97 as=1.4196 ps=8.06 w=3.64 l=1.44
X8 B.t5 B.t3 B.t4 w_n2032_n1696# sky130_fd_pr__pfet_01v8 ad=1.4196 pd=8.06 as=0 ps=0 w=3.64 l=1.44
X9 B.t2 B.t0 B.t1 w_n2032_n1696# sky130_fd_pr__pfet_01v8 ad=1.4196 pd=8.06 as=0 ps=0 w=3.64 l=1.44
X10 VDD1.t0 VP.t3 VTAIL.t5 w_n2032_n1696# sky130_fd_pr__pfet_01v8 ad=0.6006 pd=3.97 as=1.4196 ps=8.06 w=3.64 l=1.44
X11 VTAIL.t3 VN.t3 VDD2.t0 w_n2032_n1696# sky130_fd_pr__pfet_01v8 ad=1.4196 pd=8.06 as=0.6006 ps=3.97 w=3.64 l=1.44
R0 VP.n4 VP.n3 179.071
R1 VP.n12 VP.n11 179.071
R2 VP.n10 VP.n0 161.3
R3 VP.n9 VP.n8 161.3
R4 VP.n7 VP.n1 161.3
R5 VP.n6 VP.n5 161.3
R6 VP.n2 VP.t2 96.317
R7 VP.n2 VP.t3 96.0064
R8 VP.n4 VP.t1 60.9199
R9 VP.n11 VP.t0 60.9199
R10 VP.n9 VP.n1 56.4773
R11 VP.n3 VP.n2 49.558
R12 VP.n5 VP.n1 24.3439
R13 VP.n10 VP.n9 24.3439
R14 VP.n5 VP.n4 6.57323
R15 VP.n11 VP.n10 6.57323
R16 VP.n6 VP.n3 0.189894
R17 VP.n7 VP.n6 0.189894
R18 VP.n8 VP.n7 0.189894
R19 VP.n8 VP.n0 0.189894
R20 VP.n12 VP.n0 0.189894
R21 VP VP.n12 0.0516364
R22 VTAIL.n5 VTAIL.t4 115.263
R23 VTAIL.n4 VTAIL.t0 115.263
R24 VTAIL.n3 VTAIL.t3 115.263
R25 VTAIL.n7 VTAIL.t2 115.263
R26 VTAIL.n0 VTAIL.t1 115.263
R27 VTAIL.n1 VTAIL.t6 115.263
R28 VTAIL.n2 VTAIL.t7 115.263
R29 VTAIL.n6 VTAIL.t5 115.263
R30 VTAIL.n7 VTAIL.n6 17.0307
R31 VTAIL.n3 VTAIL.n2 17.0307
R32 VTAIL.n4 VTAIL.n3 1.52636
R33 VTAIL.n6 VTAIL.n5 1.52636
R34 VTAIL.n2 VTAIL.n1 1.52636
R35 VTAIL VTAIL.n0 0.821621
R36 VTAIL VTAIL.n7 0.705241
R37 VTAIL.n5 VTAIL.n4 0.470328
R38 VTAIL.n1 VTAIL.n0 0.470328
R39 VDD1 VDD1.n1 154.966
R40 VDD1 VDD1.n0 123.07
R41 VDD1.n0 VDD1.t1 8.93044
R42 VDD1.n0 VDD1.t0 8.93044
R43 VDD1.n1 VDD1.t2 8.93044
R44 VDD1.n1 VDD1.t3 8.93044
R45 B.n201 B.n64 585
R46 B.n200 B.n199 585
R47 B.n198 B.n65 585
R48 B.n197 B.n196 585
R49 B.n195 B.n66 585
R50 B.n194 B.n193 585
R51 B.n192 B.n67 585
R52 B.n191 B.n190 585
R53 B.n189 B.n68 585
R54 B.n188 B.n187 585
R55 B.n186 B.n69 585
R56 B.n185 B.n184 585
R57 B.n183 B.n70 585
R58 B.n182 B.n181 585
R59 B.n180 B.n71 585
R60 B.n179 B.n178 585
R61 B.n177 B.n72 585
R62 B.n176 B.n175 585
R63 B.n171 B.n73 585
R64 B.n170 B.n169 585
R65 B.n168 B.n74 585
R66 B.n167 B.n166 585
R67 B.n165 B.n75 585
R68 B.n164 B.n163 585
R69 B.n162 B.n76 585
R70 B.n161 B.n160 585
R71 B.n159 B.n77 585
R72 B.n157 B.n156 585
R73 B.n155 B.n80 585
R74 B.n154 B.n153 585
R75 B.n152 B.n81 585
R76 B.n151 B.n150 585
R77 B.n149 B.n82 585
R78 B.n148 B.n147 585
R79 B.n146 B.n83 585
R80 B.n145 B.n144 585
R81 B.n143 B.n84 585
R82 B.n142 B.n141 585
R83 B.n140 B.n85 585
R84 B.n139 B.n138 585
R85 B.n137 B.n86 585
R86 B.n136 B.n135 585
R87 B.n134 B.n87 585
R88 B.n133 B.n132 585
R89 B.n203 B.n202 585
R90 B.n204 B.n63 585
R91 B.n206 B.n205 585
R92 B.n207 B.n62 585
R93 B.n209 B.n208 585
R94 B.n210 B.n61 585
R95 B.n212 B.n211 585
R96 B.n213 B.n60 585
R97 B.n215 B.n214 585
R98 B.n216 B.n59 585
R99 B.n218 B.n217 585
R100 B.n219 B.n58 585
R101 B.n221 B.n220 585
R102 B.n222 B.n57 585
R103 B.n224 B.n223 585
R104 B.n225 B.n56 585
R105 B.n227 B.n226 585
R106 B.n228 B.n55 585
R107 B.n230 B.n229 585
R108 B.n231 B.n54 585
R109 B.n233 B.n232 585
R110 B.n234 B.n53 585
R111 B.n236 B.n235 585
R112 B.n237 B.n52 585
R113 B.n239 B.n238 585
R114 B.n240 B.n51 585
R115 B.n242 B.n241 585
R116 B.n243 B.n50 585
R117 B.n245 B.n244 585
R118 B.n246 B.n49 585
R119 B.n248 B.n247 585
R120 B.n249 B.n48 585
R121 B.n251 B.n250 585
R122 B.n252 B.n47 585
R123 B.n254 B.n253 585
R124 B.n255 B.n46 585
R125 B.n257 B.n256 585
R126 B.n258 B.n45 585
R127 B.n260 B.n259 585
R128 B.n261 B.n44 585
R129 B.n263 B.n262 585
R130 B.n264 B.n43 585
R131 B.n266 B.n265 585
R132 B.n267 B.n42 585
R133 B.n269 B.n268 585
R134 B.n270 B.n41 585
R135 B.n272 B.n271 585
R136 B.n273 B.n40 585
R137 B.n341 B.n340 585
R138 B.n339 B.n14 585
R139 B.n338 B.n337 585
R140 B.n336 B.n15 585
R141 B.n335 B.n334 585
R142 B.n333 B.n16 585
R143 B.n332 B.n331 585
R144 B.n330 B.n17 585
R145 B.n329 B.n328 585
R146 B.n327 B.n18 585
R147 B.n326 B.n325 585
R148 B.n324 B.n19 585
R149 B.n323 B.n322 585
R150 B.n321 B.n20 585
R151 B.n320 B.n319 585
R152 B.n318 B.n21 585
R153 B.n317 B.n316 585
R154 B.n315 B.n314 585
R155 B.n313 B.n25 585
R156 B.n312 B.n311 585
R157 B.n310 B.n26 585
R158 B.n309 B.n308 585
R159 B.n307 B.n27 585
R160 B.n306 B.n305 585
R161 B.n304 B.n28 585
R162 B.n303 B.n302 585
R163 B.n301 B.n29 585
R164 B.n299 B.n298 585
R165 B.n297 B.n32 585
R166 B.n296 B.n295 585
R167 B.n294 B.n33 585
R168 B.n293 B.n292 585
R169 B.n291 B.n34 585
R170 B.n290 B.n289 585
R171 B.n288 B.n35 585
R172 B.n287 B.n286 585
R173 B.n285 B.n36 585
R174 B.n284 B.n283 585
R175 B.n282 B.n37 585
R176 B.n281 B.n280 585
R177 B.n279 B.n38 585
R178 B.n278 B.n277 585
R179 B.n276 B.n39 585
R180 B.n275 B.n274 585
R181 B.n342 B.n13 585
R182 B.n344 B.n343 585
R183 B.n345 B.n12 585
R184 B.n347 B.n346 585
R185 B.n348 B.n11 585
R186 B.n350 B.n349 585
R187 B.n351 B.n10 585
R188 B.n353 B.n352 585
R189 B.n354 B.n9 585
R190 B.n356 B.n355 585
R191 B.n357 B.n8 585
R192 B.n359 B.n358 585
R193 B.n360 B.n7 585
R194 B.n362 B.n361 585
R195 B.n363 B.n6 585
R196 B.n365 B.n364 585
R197 B.n366 B.n5 585
R198 B.n368 B.n367 585
R199 B.n369 B.n4 585
R200 B.n371 B.n370 585
R201 B.n372 B.n3 585
R202 B.n374 B.n373 585
R203 B.n375 B.n0 585
R204 B.n2 B.n1 585
R205 B.n100 B.n99 585
R206 B.n101 B.n98 585
R207 B.n103 B.n102 585
R208 B.n104 B.n97 585
R209 B.n106 B.n105 585
R210 B.n107 B.n96 585
R211 B.n109 B.n108 585
R212 B.n110 B.n95 585
R213 B.n112 B.n111 585
R214 B.n113 B.n94 585
R215 B.n115 B.n114 585
R216 B.n116 B.n93 585
R217 B.n118 B.n117 585
R218 B.n119 B.n92 585
R219 B.n121 B.n120 585
R220 B.n122 B.n91 585
R221 B.n124 B.n123 585
R222 B.n125 B.n90 585
R223 B.n127 B.n126 585
R224 B.n128 B.n89 585
R225 B.n130 B.n129 585
R226 B.n131 B.n88 585
R227 B.n132 B.n131 506.916
R228 B.n202 B.n201 506.916
R229 B.n274 B.n273 506.916
R230 B.n340 B.n13 506.916
R231 B.n172 B.t0 266.772
R232 B.n30 B.t3 266.772
R233 B.n78 B.t9 266.291
R234 B.n22 B.t6 266.291
R235 B.n377 B.n376 256.663
R236 B.n376 B.n375 235.042
R237 B.n376 B.n2 235.042
R238 B.n172 B.t1 165.174
R239 B.n30 B.t5 165.174
R240 B.n78 B.t10 165.172
R241 B.n22 B.t8 165.172
R242 B.n132 B.n87 163.367
R243 B.n136 B.n87 163.367
R244 B.n137 B.n136 163.367
R245 B.n138 B.n137 163.367
R246 B.n138 B.n85 163.367
R247 B.n142 B.n85 163.367
R248 B.n143 B.n142 163.367
R249 B.n144 B.n143 163.367
R250 B.n144 B.n83 163.367
R251 B.n148 B.n83 163.367
R252 B.n149 B.n148 163.367
R253 B.n150 B.n149 163.367
R254 B.n150 B.n81 163.367
R255 B.n154 B.n81 163.367
R256 B.n155 B.n154 163.367
R257 B.n156 B.n155 163.367
R258 B.n156 B.n77 163.367
R259 B.n161 B.n77 163.367
R260 B.n162 B.n161 163.367
R261 B.n163 B.n162 163.367
R262 B.n163 B.n75 163.367
R263 B.n167 B.n75 163.367
R264 B.n168 B.n167 163.367
R265 B.n169 B.n168 163.367
R266 B.n169 B.n73 163.367
R267 B.n176 B.n73 163.367
R268 B.n177 B.n176 163.367
R269 B.n178 B.n177 163.367
R270 B.n178 B.n71 163.367
R271 B.n182 B.n71 163.367
R272 B.n183 B.n182 163.367
R273 B.n184 B.n183 163.367
R274 B.n184 B.n69 163.367
R275 B.n188 B.n69 163.367
R276 B.n189 B.n188 163.367
R277 B.n190 B.n189 163.367
R278 B.n190 B.n67 163.367
R279 B.n194 B.n67 163.367
R280 B.n195 B.n194 163.367
R281 B.n196 B.n195 163.367
R282 B.n196 B.n65 163.367
R283 B.n200 B.n65 163.367
R284 B.n201 B.n200 163.367
R285 B.n273 B.n272 163.367
R286 B.n272 B.n41 163.367
R287 B.n268 B.n41 163.367
R288 B.n268 B.n267 163.367
R289 B.n267 B.n266 163.367
R290 B.n266 B.n43 163.367
R291 B.n262 B.n43 163.367
R292 B.n262 B.n261 163.367
R293 B.n261 B.n260 163.367
R294 B.n260 B.n45 163.367
R295 B.n256 B.n45 163.367
R296 B.n256 B.n255 163.367
R297 B.n255 B.n254 163.367
R298 B.n254 B.n47 163.367
R299 B.n250 B.n47 163.367
R300 B.n250 B.n249 163.367
R301 B.n249 B.n248 163.367
R302 B.n248 B.n49 163.367
R303 B.n244 B.n49 163.367
R304 B.n244 B.n243 163.367
R305 B.n243 B.n242 163.367
R306 B.n242 B.n51 163.367
R307 B.n238 B.n51 163.367
R308 B.n238 B.n237 163.367
R309 B.n237 B.n236 163.367
R310 B.n236 B.n53 163.367
R311 B.n232 B.n53 163.367
R312 B.n232 B.n231 163.367
R313 B.n231 B.n230 163.367
R314 B.n230 B.n55 163.367
R315 B.n226 B.n55 163.367
R316 B.n226 B.n225 163.367
R317 B.n225 B.n224 163.367
R318 B.n224 B.n57 163.367
R319 B.n220 B.n57 163.367
R320 B.n220 B.n219 163.367
R321 B.n219 B.n218 163.367
R322 B.n218 B.n59 163.367
R323 B.n214 B.n59 163.367
R324 B.n214 B.n213 163.367
R325 B.n213 B.n212 163.367
R326 B.n212 B.n61 163.367
R327 B.n208 B.n61 163.367
R328 B.n208 B.n207 163.367
R329 B.n207 B.n206 163.367
R330 B.n206 B.n63 163.367
R331 B.n202 B.n63 163.367
R332 B.n340 B.n339 163.367
R333 B.n339 B.n338 163.367
R334 B.n338 B.n15 163.367
R335 B.n334 B.n15 163.367
R336 B.n334 B.n333 163.367
R337 B.n333 B.n332 163.367
R338 B.n332 B.n17 163.367
R339 B.n328 B.n17 163.367
R340 B.n328 B.n327 163.367
R341 B.n327 B.n326 163.367
R342 B.n326 B.n19 163.367
R343 B.n322 B.n19 163.367
R344 B.n322 B.n321 163.367
R345 B.n321 B.n320 163.367
R346 B.n320 B.n21 163.367
R347 B.n316 B.n21 163.367
R348 B.n316 B.n315 163.367
R349 B.n315 B.n25 163.367
R350 B.n311 B.n25 163.367
R351 B.n311 B.n310 163.367
R352 B.n310 B.n309 163.367
R353 B.n309 B.n27 163.367
R354 B.n305 B.n27 163.367
R355 B.n305 B.n304 163.367
R356 B.n304 B.n303 163.367
R357 B.n303 B.n29 163.367
R358 B.n298 B.n29 163.367
R359 B.n298 B.n297 163.367
R360 B.n297 B.n296 163.367
R361 B.n296 B.n33 163.367
R362 B.n292 B.n33 163.367
R363 B.n292 B.n291 163.367
R364 B.n291 B.n290 163.367
R365 B.n290 B.n35 163.367
R366 B.n286 B.n35 163.367
R367 B.n286 B.n285 163.367
R368 B.n285 B.n284 163.367
R369 B.n284 B.n37 163.367
R370 B.n280 B.n37 163.367
R371 B.n280 B.n279 163.367
R372 B.n279 B.n278 163.367
R373 B.n278 B.n39 163.367
R374 B.n274 B.n39 163.367
R375 B.n344 B.n13 163.367
R376 B.n345 B.n344 163.367
R377 B.n346 B.n345 163.367
R378 B.n346 B.n11 163.367
R379 B.n350 B.n11 163.367
R380 B.n351 B.n350 163.367
R381 B.n352 B.n351 163.367
R382 B.n352 B.n9 163.367
R383 B.n356 B.n9 163.367
R384 B.n357 B.n356 163.367
R385 B.n358 B.n357 163.367
R386 B.n358 B.n7 163.367
R387 B.n362 B.n7 163.367
R388 B.n363 B.n362 163.367
R389 B.n364 B.n363 163.367
R390 B.n364 B.n5 163.367
R391 B.n368 B.n5 163.367
R392 B.n369 B.n368 163.367
R393 B.n370 B.n369 163.367
R394 B.n370 B.n3 163.367
R395 B.n374 B.n3 163.367
R396 B.n375 B.n374 163.367
R397 B.n100 B.n2 163.367
R398 B.n101 B.n100 163.367
R399 B.n102 B.n101 163.367
R400 B.n102 B.n97 163.367
R401 B.n106 B.n97 163.367
R402 B.n107 B.n106 163.367
R403 B.n108 B.n107 163.367
R404 B.n108 B.n95 163.367
R405 B.n112 B.n95 163.367
R406 B.n113 B.n112 163.367
R407 B.n114 B.n113 163.367
R408 B.n114 B.n93 163.367
R409 B.n118 B.n93 163.367
R410 B.n119 B.n118 163.367
R411 B.n120 B.n119 163.367
R412 B.n120 B.n91 163.367
R413 B.n124 B.n91 163.367
R414 B.n125 B.n124 163.367
R415 B.n126 B.n125 163.367
R416 B.n126 B.n89 163.367
R417 B.n130 B.n89 163.367
R418 B.n131 B.n130 163.367
R419 B.n173 B.t2 130.847
R420 B.n31 B.t4 130.847
R421 B.n79 B.t11 130.845
R422 B.n23 B.t7 130.845
R423 B.n158 B.n79 59.5399
R424 B.n174 B.n173 59.5399
R425 B.n300 B.n31 59.5399
R426 B.n24 B.n23 59.5399
R427 B.n79 B.n78 34.3278
R428 B.n173 B.n172 34.3278
R429 B.n31 B.n30 34.3278
R430 B.n23 B.n22 34.3278
R431 B.n342 B.n341 32.9371
R432 B.n275 B.n40 32.9371
R433 B.n203 B.n64 32.9371
R434 B.n133 B.n88 32.9371
R435 B B.n377 18.0485
R436 B.n343 B.n342 10.6151
R437 B.n343 B.n12 10.6151
R438 B.n347 B.n12 10.6151
R439 B.n348 B.n347 10.6151
R440 B.n349 B.n348 10.6151
R441 B.n349 B.n10 10.6151
R442 B.n353 B.n10 10.6151
R443 B.n354 B.n353 10.6151
R444 B.n355 B.n354 10.6151
R445 B.n355 B.n8 10.6151
R446 B.n359 B.n8 10.6151
R447 B.n360 B.n359 10.6151
R448 B.n361 B.n360 10.6151
R449 B.n361 B.n6 10.6151
R450 B.n365 B.n6 10.6151
R451 B.n366 B.n365 10.6151
R452 B.n367 B.n366 10.6151
R453 B.n367 B.n4 10.6151
R454 B.n371 B.n4 10.6151
R455 B.n372 B.n371 10.6151
R456 B.n373 B.n372 10.6151
R457 B.n373 B.n0 10.6151
R458 B.n341 B.n14 10.6151
R459 B.n337 B.n14 10.6151
R460 B.n337 B.n336 10.6151
R461 B.n336 B.n335 10.6151
R462 B.n335 B.n16 10.6151
R463 B.n331 B.n16 10.6151
R464 B.n331 B.n330 10.6151
R465 B.n330 B.n329 10.6151
R466 B.n329 B.n18 10.6151
R467 B.n325 B.n18 10.6151
R468 B.n325 B.n324 10.6151
R469 B.n324 B.n323 10.6151
R470 B.n323 B.n20 10.6151
R471 B.n319 B.n20 10.6151
R472 B.n319 B.n318 10.6151
R473 B.n318 B.n317 10.6151
R474 B.n314 B.n313 10.6151
R475 B.n313 B.n312 10.6151
R476 B.n312 B.n26 10.6151
R477 B.n308 B.n26 10.6151
R478 B.n308 B.n307 10.6151
R479 B.n307 B.n306 10.6151
R480 B.n306 B.n28 10.6151
R481 B.n302 B.n28 10.6151
R482 B.n302 B.n301 10.6151
R483 B.n299 B.n32 10.6151
R484 B.n295 B.n32 10.6151
R485 B.n295 B.n294 10.6151
R486 B.n294 B.n293 10.6151
R487 B.n293 B.n34 10.6151
R488 B.n289 B.n34 10.6151
R489 B.n289 B.n288 10.6151
R490 B.n288 B.n287 10.6151
R491 B.n287 B.n36 10.6151
R492 B.n283 B.n36 10.6151
R493 B.n283 B.n282 10.6151
R494 B.n282 B.n281 10.6151
R495 B.n281 B.n38 10.6151
R496 B.n277 B.n38 10.6151
R497 B.n277 B.n276 10.6151
R498 B.n276 B.n275 10.6151
R499 B.n271 B.n40 10.6151
R500 B.n271 B.n270 10.6151
R501 B.n270 B.n269 10.6151
R502 B.n269 B.n42 10.6151
R503 B.n265 B.n42 10.6151
R504 B.n265 B.n264 10.6151
R505 B.n264 B.n263 10.6151
R506 B.n263 B.n44 10.6151
R507 B.n259 B.n44 10.6151
R508 B.n259 B.n258 10.6151
R509 B.n258 B.n257 10.6151
R510 B.n257 B.n46 10.6151
R511 B.n253 B.n46 10.6151
R512 B.n253 B.n252 10.6151
R513 B.n252 B.n251 10.6151
R514 B.n251 B.n48 10.6151
R515 B.n247 B.n48 10.6151
R516 B.n247 B.n246 10.6151
R517 B.n246 B.n245 10.6151
R518 B.n245 B.n50 10.6151
R519 B.n241 B.n50 10.6151
R520 B.n241 B.n240 10.6151
R521 B.n240 B.n239 10.6151
R522 B.n239 B.n52 10.6151
R523 B.n235 B.n52 10.6151
R524 B.n235 B.n234 10.6151
R525 B.n234 B.n233 10.6151
R526 B.n233 B.n54 10.6151
R527 B.n229 B.n54 10.6151
R528 B.n229 B.n228 10.6151
R529 B.n228 B.n227 10.6151
R530 B.n227 B.n56 10.6151
R531 B.n223 B.n56 10.6151
R532 B.n223 B.n222 10.6151
R533 B.n222 B.n221 10.6151
R534 B.n221 B.n58 10.6151
R535 B.n217 B.n58 10.6151
R536 B.n217 B.n216 10.6151
R537 B.n216 B.n215 10.6151
R538 B.n215 B.n60 10.6151
R539 B.n211 B.n60 10.6151
R540 B.n211 B.n210 10.6151
R541 B.n210 B.n209 10.6151
R542 B.n209 B.n62 10.6151
R543 B.n205 B.n62 10.6151
R544 B.n205 B.n204 10.6151
R545 B.n204 B.n203 10.6151
R546 B.n99 B.n1 10.6151
R547 B.n99 B.n98 10.6151
R548 B.n103 B.n98 10.6151
R549 B.n104 B.n103 10.6151
R550 B.n105 B.n104 10.6151
R551 B.n105 B.n96 10.6151
R552 B.n109 B.n96 10.6151
R553 B.n110 B.n109 10.6151
R554 B.n111 B.n110 10.6151
R555 B.n111 B.n94 10.6151
R556 B.n115 B.n94 10.6151
R557 B.n116 B.n115 10.6151
R558 B.n117 B.n116 10.6151
R559 B.n117 B.n92 10.6151
R560 B.n121 B.n92 10.6151
R561 B.n122 B.n121 10.6151
R562 B.n123 B.n122 10.6151
R563 B.n123 B.n90 10.6151
R564 B.n127 B.n90 10.6151
R565 B.n128 B.n127 10.6151
R566 B.n129 B.n128 10.6151
R567 B.n129 B.n88 10.6151
R568 B.n134 B.n133 10.6151
R569 B.n135 B.n134 10.6151
R570 B.n135 B.n86 10.6151
R571 B.n139 B.n86 10.6151
R572 B.n140 B.n139 10.6151
R573 B.n141 B.n140 10.6151
R574 B.n141 B.n84 10.6151
R575 B.n145 B.n84 10.6151
R576 B.n146 B.n145 10.6151
R577 B.n147 B.n146 10.6151
R578 B.n147 B.n82 10.6151
R579 B.n151 B.n82 10.6151
R580 B.n152 B.n151 10.6151
R581 B.n153 B.n152 10.6151
R582 B.n153 B.n80 10.6151
R583 B.n157 B.n80 10.6151
R584 B.n160 B.n159 10.6151
R585 B.n160 B.n76 10.6151
R586 B.n164 B.n76 10.6151
R587 B.n165 B.n164 10.6151
R588 B.n166 B.n165 10.6151
R589 B.n166 B.n74 10.6151
R590 B.n170 B.n74 10.6151
R591 B.n171 B.n170 10.6151
R592 B.n175 B.n171 10.6151
R593 B.n179 B.n72 10.6151
R594 B.n180 B.n179 10.6151
R595 B.n181 B.n180 10.6151
R596 B.n181 B.n70 10.6151
R597 B.n185 B.n70 10.6151
R598 B.n186 B.n185 10.6151
R599 B.n187 B.n186 10.6151
R600 B.n187 B.n68 10.6151
R601 B.n191 B.n68 10.6151
R602 B.n192 B.n191 10.6151
R603 B.n193 B.n192 10.6151
R604 B.n193 B.n66 10.6151
R605 B.n197 B.n66 10.6151
R606 B.n198 B.n197 10.6151
R607 B.n199 B.n198 10.6151
R608 B.n199 B.n64 10.6151
R609 B.n317 B.n24 9.52245
R610 B.n300 B.n299 9.52245
R611 B.n158 B.n157 9.52245
R612 B.n174 B.n72 9.52245
R613 B.n377 B.n0 8.11757
R614 B.n377 B.n1 8.11757
R615 B.n314 B.n24 1.09318
R616 B.n301 B.n300 1.09318
R617 B.n159 B.n158 1.09318
R618 B.n175 B.n174 1.09318
R619 VN.n0 VN.t0 96.317
R620 VN.n1 VN.t2 96.317
R621 VN.n0 VN.t1 96.0064
R622 VN.n1 VN.t3 96.0064
R623 VN VN.n1 49.9386
R624 VN VN.n0 13.2985
R625 VDD2.n2 VDD2.n0 154.441
R626 VDD2.n2 VDD2.n1 123.011
R627 VDD2.n1 VDD2.t0 8.93044
R628 VDD2.n1 VDD2.t1 8.93044
R629 VDD2.n0 VDD2.t3 8.93044
R630 VDD2.n0 VDD2.t2 8.93044
R631 VDD2 VDD2.n2 0.0586897
C0 VDD2 VN 1.46532f
C1 VP VN 3.81889f
C2 VTAIL VDD1 3.00157f
C3 VDD2 VDD1 0.744985f
C4 VP VDD1 1.63738f
C5 VDD2 VTAIL 3.048f
C6 VTAIL VP 1.6614f
C7 B w_n2032_n1696# 5.48786f
C8 VDD2 VP 0.3252f
C9 w_n2032_n1696# VN 3.07467f
C10 w_n2032_n1696# VDD1 0.998684f
C11 VTAIL w_n2032_n1696# 2.00008f
C12 VDD2 w_n2032_n1696# 1.02855f
C13 VP w_n2032_n1696# 3.3316f
C14 B VN 0.789552f
C15 B VDD1 0.831699f
C16 VTAIL B 1.81163f
C17 VDD1 VN 0.152219f
C18 VDD2 B 0.865038f
C19 VP B 1.2125f
C20 VTAIL VN 1.64729f
C21 VDD2 VSUBS 0.518256f
C22 VDD1 VSUBS 2.751466f
C23 VTAIL VSUBS 0.441715f
C24 VN VSUBS 3.99681f
C25 VP VSUBS 1.225851f
C26 B VSUBS 2.437396f
C27 w_n2032_n1696# VSUBS 43.4767f
C28 VDD2.t3 VSUBS 0.052048f
C29 VDD2.t2 VSUBS 0.052048f
C30 VDD2.n0 VSUBS 0.459376f
C31 VDD2.t0 VSUBS 0.052048f
C32 VDD2.t1 VSUBS 0.052048f
C33 VDD2.n1 VSUBS 0.294083f
C34 VDD2.n2 VSUBS 1.94549f
C35 VN.t0 VSUBS 0.677878f
C36 VN.t1 VSUBS 0.676575f
C37 VN.n0 VSUBS 0.547392f
C38 VN.t2 VSUBS 0.677878f
C39 VN.t3 VSUBS 0.676575f
C40 VN.n1 VSUBS 1.66888f
C41 B.n0 VSUBS 0.00662f
C42 B.n1 VSUBS 0.00662f
C43 B.n2 VSUBS 0.009791f
C44 B.n3 VSUBS 0.007503f
C45 B.n4 VSUBS 0.007503f
C46 B.n5 VSUBS 0.007503f
C47 B.n6 VSUBS 0.007503f
C48 B.n7 VSUBS 0.007503f
C49 B.n8 VSUBS 0.007503f
C50 B.n9 VSUBS 0.007503f
C51 B.n10 VSUBS 0.007503f
C52 B.n11 VSUBS 0.007503f
C53 B.n12 VSUBS 0.007503f
C54 B.n13 VSUBS 0.016935f
C55 B.n14 VSUBS 0.007503f
C56 B.n15 VSUBS 0.007503f
C57 B.n16 VSUBS 0.007503f
C58 B.n17 VSUBS 0.007503f
C59 B.n18 VSUBS 0.007503f
C60 B.n19 VSUBS 0.007503f
C61 B.n20 VSUBS 0.007503f
C62 B.n21 VSUBS 0.007503f
C63 B.t7 VSUBS 0.099513f
C64 B.t8 VSUBS 0.11133f
C65 B.t6 VSUBS 0.264561f
C66 B.n22 VSUBS 0.084176f
C67 B.n23 VSUBS 0.067564f
C68 B.n24 VSUBS 0.017383f
C69 B.n25 VSUBS 0.007503f
C70 B.n26 VSUBS 0.007503f
C71 B.n27 VSUBS 0.007503f
C72 B.n28 VSUBS 0.007503f
C73 B.n29 VSUBS 0.007503f
C74 B.t4 VSUBS 0.099513f
C75 B.t5 VSUBS 0.11133f
C76 B.t3 VSUBS 0.264592f
C77 B.n30 VSUBS 0.084146f
C78 B.n31 VSUBS 0.067564f
C79 B.n32 VSUBS 0.007503f
C80 B.n33 VSUBS 0.007503f
C81 B.n34 VSUBS 0.007503f
C82 B.n35 VSUBS 0.007503f
C83 B.n36 VSUBS 0.007503f
C84 B.n37 VSUBS 0.007503f
C85 B.n38 VSUBS 0.007503f
C86 B.n39 VSUBS 0.007503f
C87 B.n40 VSUBS 0.016935f
C88 B.n41 VSUBS 0.007503f
C89 B.n42 VSUBS 0.007503f
C90 B.n43 VSUBS 0.007503f
C91 B.n44 VSUBS 0.007503f
C92 B.n45 VSUBS 0.007503f
C93 B.n46 VSUBS 0.007503f
C94 B.n47 VSUBS 0.007503f
C95 B.n48 VSUBS 0.007503f
C96 B.n49 VSUBS 0.007503f
C97 B.n50 VSUBS 0.007503f
C98 B.n51 VSUBS 0.007503f
C99 B.n52 VSUBS 0.007503f
C100 B.n53 VSUBS 0.007503f
C101 B.n54 VSUBS 0.007503f
C102 B.n55 VSUBS 0.007503f
C103 B.n56 VSUBS 0.007503f
C104 B.n57 VSUBS 0.007503f
C105 B.n58 VSUBS 0.007503f
C106 B.n59 VSUBS 0.007503f
C107 B.n60 VSUBS 0.007503f
C108 B.n61 VSUBS 0.007503f
C109 B.n62 VSUBS 0.007503f
C110 B.n63 VSUBS 0.007503f
C111 B.n64 VSUBS 0.017493f
C112 B.n65 VSUBS 0.007503f
C113 B.n66 VSUBS 0.007503f
C114 B.n67 VSUBS 0.007503f
C115 B.n68 VSUBS 0.007503f
C116 B.n69 VSUBS 0.007503f
C117 B.n70 VSUBS 0.007503f
C118 B.n71 VSUBS 0.007503f
C119 B.n72 VSUBS 0.007117f
C120 B.n73 VSUBS 0.007503f
C121 B.n74 VSUBS 0.007503f
C122 B.n75 VSUBS 0.007503f
C123 B.n76 VSUBS 0.007503f
C124 B.n77 VSUBS 0.007503f
C125 B.t11 VSUBS 0.099513f
C126 B.t10 VSUBS 0.11133f
C127 B.t9 VSUBS 0.264561f
C128 B.n78 VSUBS 0.084176f
C129 B.n79 VSUBS 0.067564f
C130 B.n80 VSUBS 0.007503f
C131 B.n81 VSUBS 0.007503f
C132 B.n82 VSUBS 0.007503f
C133 B.n83 VSUBS 0.007503f
C134 B.n84 VSUBS 0.007503f
C135 B.n85 VSUBS 0.007503f
C136 B.n86 VSUBS 0.007503f
C137 B.n87 VSUBS 0.007503f
C138 B.n88 VSUBS 0.016935f
C139 B.n89 VSUBS 0.007503f
C140 B.n90 VSUBS 0.007503f
C141 B.n91 VSUBS 0.007503f
C142 B.n92 VSUBS 0.007503f
C143 B.n93 VSUBS 0.007503f
C144 B.n94 VSUBS 0.007503f
C145 B.n95 VSUBS 0.007503f
C146 B.n96 VSUBS 0.007503f
C147 B.n97 VSUBS 0.007503f
C148 B.n98 VSUBS 0.007503f
C149 B.n99 VSUBS 0.007503f
C150 B.n100 VSUBS 0.007503f
C151 B.n101 VSUBS 0.007503f
C152 B.n102 VSUBS 0.007503f
C153 B.n103 VSUBS 0.007503f
C154 B.n104 VSUBS 0.007503f
C155 B.n105 VSUBS 0.007503f
C156 B.n106 VSUBS 0.007503f
C157 B.n107 VSUBS 0.007503f
C158 B.n108 VSUBS 0.007503f
C159 B.n109 VSUBS 0.007503f
C160 B.n110 VSUBS 0.007503f
C161 B.n111 VSUBS 0.007503f
C162 B.n112 VSUBS 0.007503f
C163 B.n113 VSUBS 0.007503f
C164 B.n114 VSUBS 0.007503f
C165 B.n115 VSUBS 0.007503f
C166 B.n116 VSUBS 0.007503f
C167 B.n117 VSUBS 0.007503f
C168 B.n118 VSUBS 0.007503f
C169 B.n119 VSUBS 0.007503f
C170 B.n120 VSUBS 0.007503f
C171 B.n121 VSUBS 0.007503f
C172 B.n122 VSUBS 0.007503f
C173 B.n123 VSUBS 0.007503f
C174 B.n124 VSUBS 0.007503f
C175 B.n125 VSUBS 0.007503f
C176 B.n126 VSUBS 0.007503f
C177 B.n127 VSUBS 0.007503f
C178 B.n128 VSUBS 0.007503f
C179 B.n129 VSUBS 0.007503f
C180 B.n130 VSUBS 0.007503f
C181 B.n131 VSUBS 0.016935f
C182 B.n132 VSUBS 0.018372f
C183 B.n133 VSUBS 0.018372f
C184 B.n134 VSUBS 0.007503f
C185 B.n135 VSUBS 0.007503f
C186 B.n136 VSUBS 0.007503f
C187 B.n137 VSUBS 0.007503f
C188 B.n138 VSUBS 0.007503f
C189 B.n139 VSUBS 0.007503f
C190 B.n140 VSUBS 0.007503f
C191 B.n141 VSUBS 0.007503f
C192 B.n142 VSUBS 0.007503f
C193 B.n143 VSUBS 0.007503f
C194 B.n144 VSUBS 0.007503f
C195 B.n145 VSUBS 0.007503f
C196 B.n146 VSUBS 0.007503f
C197 B.n147 VSUBS 0.007503f
C198 B.n148 VSUBS 0.007503f
C199 B.n149 VSUBS 0.007503f
C200 B.n150 VSUBS 0.007503f
C201 B.n151 VSUBS 0.007503f
C202 B.n152 VSUBS 0.007503f
C203 B.n153 VSUBS 0.007503f
C204 B.n154 VSUBS 0.007503f
C205 B.n155 VSUBS 0.007503f
C206 B.n156 VSUBS 0.007503f
C207 B.n157 VSUBS 0.007117f
C208 B.n158 VSUBS 0.017383f
C209 B.n159 VSUBS 0.004138f
C210 B.n160 VSUBS 0.007503f
C211 B.n161 VSUBS 0.007503f
C212 B.n162 VSUBS 0.007503f
C213 B.n163 VSUBS 0.007503f
C214 B.n164 VSUBS 0.007503f
C215 B.n165 VSUBS 0.007503f
C216 B.n166 VSUBS 0.007503f
C217 B.n167 VSUBS 0.007503f
C218 B.n168 VSUBS 0.007503f
C219 B.n169 VSUBS 0.007503f
C220 B.n170 VSUBS 0.007503f
C221 B.n171 VSUBS 0.007503f
C222 B.t2 VSUBS 0.099513f
C223 B.t1 VSUBS 0.11133f
C224 B.t0 VSUBS 0.264592f
C225 B.n172 VSUBS 0.084146f
C226 B.n173 VSUBS 0.067564f
C227 B.n174 VSUBS 0.017383f
C228 B.n175 VSUBS 0.004138f
C229 B.n176 VSUBS 0.007503f
C230 B.n177 VSUBS 0.007503f
C231 B.n178 VSUBS 0.007503f
C232 B.n179 VSUBS 0.007503f
C233 B.n180 VSUBS 0.007503f
C234 B.n181 VSUBS 0.007503f
C235 B.n182 VSUBS 0.007503f
C236 B.n183 VSUBS 0.007503f
C237 B.n184 VSUBS 0.007503f
C238 B.n185 VSUBS 0.007503f
C239 B.n186 VSUBS 0.007503f
C240 B.n187 VSUBS 0.007503f
C241 B.n188 VSUBS 0.007503f
C242 B.n189 VSUBS 0.007503f
C243 B.n190 VSUBS 0.007503f
C244 B.n191 VSUBS 0.007503f
C245 B.n192 VSUBS 0.007503f
C246 B.n193 VSUBS 0.007503f
C247 B.n194 VSUBS 0.007503f
C248 B.n195 VSUBS 0.007503f
C249 B.n196 VSUBS 0.007503f
C250 B.n197 VSUBS 0.007503f
C251 B.n198 VSUBS 0.007503f
C252 B.n199 VSUBS 0.007503f
C253 B.n200 VSUBS 0.007503f
C254 B.n201 VSUBS 0.018372f
C255 B.n202 VSUBS 0.016935f
C256 B.n203 VSUBS 0.017814f
C257 B.n204 VSUBS 0.007503f
C258 B.n205 VSUBS 0.007503f
C259 B.n206 VSUBS 0.007503f
C260 B.n207 VSUBS 0.007503f
C261 B.n208 VSUBS 0.007503f
C262 B.n209 VSUBS 0.007503f
C263 B.n210 VSUBS 0.007503f
C264 B.n211 VSUBS 0.007503f
C265 B.n212 VSUBS 0.007503f
C266 B.n213 VSUBS 0.007503f
C267 B.n214 VSUBS 0.007503f
C268 B.n215 VSUBS 0.007503f
C269 B.n216 VSUBS 0.007503f
C270 B.n217 VSUBS 0.007503f
C271 B.n218 VSUBS 0.007503f
C272 B.n219 VSUBS 0.007503f
C273 B.n220 VSUBS 0.007503f
C274 B.n221 VSUBS 0.007503f
C275 B.n222 VSUBS 0.007503f
C276 B.n223 VSUBS 0.007503f
C277 B.n224 VSUBS 0.007503f
C278 B.n225 VSUBS 0.007503f
C279 B.n226 VSUBS 0.007503f
C280 B.n227 VSUBS 0.007503f
C281 B.n228 VSUBS 0.007503f
C282 B.n229 VSUBS 0.007503f
C283 B.n230 VSUBS 0.007503f
C284 B.n231 VSUBS 0.007503f
C285 B.n232 VSUBS 0.007503f
C286 B.n233 VSUBS 0.007503f
C287 B.n234 VSUBS 0.007503f
C288 B.n235 VSUBS 0.007503f
C289 B.n236 VSUBS 0.007503f
C290 B.n237 VSUBS 0.007503f
C291 B.n238 VSUBS 0.007503f
C292 B.n239 VSUBS 0.007503f
C293 B.n240 VSUBS 0.007503f
C294 B.n241 VSUBS 0.007503f
C295 B.n242 VSUBS 0.007503f
C296 B.n243 VSUBS 0.007503f
C297 B.n244 VSUBS 0.007503f
C298 B.n245 VSUBS 0.007503f
C299 B.n246 VSUBS 0.007503f
C300 B.n247 VSUBS 0.007503f
C301 B.n248 VSUBS 0.007503f
C302 B.n249 VSUBS 0.007503f
C303 B.n250 VSUBS 0.007503f
C304 B.n251 VSUBS 0.007503f
C305 B.n252 VSUBS 0.007503f
C306 B.n253 VSUBS 0.007503f
C307 B.n254 VSUBS 0.007503f
C308 B.n255 VSUBS 0.007503f
C309 B.n256 VSUBS 0.007503f
C310 B.n257 VSUBS 0.007503f
C311 B.n258 VSUBS 0.007503f
C312 B.n259 VSUBS 0.007503f
C313 B.n260 VSUBS 0.007503f
C314 B.n261 VSUBS 0.007503f
C315 B.n262 VSUBS 0.007503f
C316 B.n263 VSUBS 0.007503f
C317 B.n264 VSUBS 0.007503f
C318 B.n265 VSUBS 0.007503f
C319 B.n266 VSUBS 0.007503f
C320 B.n267 VSUBS 0.007503f
C321 B.n268 VSUBS 0.007503f
C322 B.n269 VSUBS 0.007503f
C323 B.n270 VSUBS 0.007503f
C324 B.n271 VSUBS 0.007503f
C325 B.n272 VSUBS 0.007503f
C326 B.n273 VSUBS 0.016935f
C327 B.n274 VSUBS 0.018372f
C328 B.n275 VSUBS 0.018372f
C329 B.n276 VSUBS 0.007503f
C330 B.n277 VSUBS 0.007503f
C331 B.n278 VSUBS 0.007503f
C332 B.n279 VSUBS 0.007503f
C333 B.n280 VSUBS 0.007503f
C334 B.n281 VSUBS 0.007503f
C335 B.n282 VSUBS 0.007503f
C336 B.n283 VSUBS 0.007503f
C337 B.n284 VSUBS 0.007503f
C338 B.n285 VSUBS 0.007503f
C339 B.n286 VSUBS 0.007503f
C340 B.n287 VSUBS 0.007503f
C341 B.n288 VSUBS 0.007503f
C342 B.n289 VSUBS 0.007503f
C343 B.n290 VSUBS 0.007503f
C344 B.n291 VSUBS 0.007503f
C345 B.n292 VSUBS 0.007503f
C346 B.n293 VSUBS 0.007503f
C347 B.n294 VSUBS 0.007503f
C348 B.n295 VSUBS 0.007503f
C349 B.n296 VSUBS 0.007503f
C350 B.n297 VSUBS 0.007503f
C351 B.n298 VSUBS 0.007503f
C352 B.n299 VSUBS 0.007117f
C353 B.n300 VSUBS 0.017383f
C354 B.n301 VSUBS 0.004138f
C355 B.n302 VSUBS 0.007503f
C356 B.n303 VSUBS 0.007503f
C357 B.n304 VSUBS 0.007503f
C358 B.n305 VSUBS 0.007503f
C359 B.n306 VSUBS 0.007503f
C360 B.n307 VSUBS 0.007503f
C361 B.n308 VSUBS 0.007503f
C362 B.n309 VSUBS 0.007503f
C363 B.n310 VSUBS 0.007503f
C364 B.n311 VSUBS 0.007503f
C365 B.n312 VSUBS 0.007503f
C366 B.n313 VSUBS 0.007503f
C367 B.n314 VSUBS 0.004138f
C368 B.n315 VSUBS 0.007503f
C369 B.n316 VSUBS 0.007503f
C370 B.n317 VSUBS 0.007117f
C371 B.n318 VSUBS 0.007503f
C372 B.n319 VSUBS 0.007503f
C373 B.n320 VSUBS 0.007503f
C374 B.n321 VSUBS 0.007503f
C375 B.n322 VSUBS 0.007503f
C376 B.n323 VSUBS 0.007503f
C377 B.n324 VSUBS 0.007503f
C378 B.n325 VSUBS 0.007503f
C379 B.n326 VSUBS 0.007503f
C380 B.n327 VSUBS 0.007503f
C381 B.n328 VSUBS 0.007503f
C382 B.n329 VSUBS 0.007503f
C383 B.n330 VSUBS 0.007503f
C384 B.n331 VSUBS 0.007503f
C385 B.n332 VSUBS 0.007503f
C386 B.n333 VSUBS 0.007503f
C387 B.n334 VSUBS 0.007503f
C388 B.n335 VSUBS 0.007503f
C389 B.n336 VSUBS 0.007503f
C390 B.n337 VSUBS 0.007503f
C391 B.n338 VSUBS 0.007503f
C392 B.n339 VSUBS 0.007503f
C393 B.n340 VSUBS 0.018372f
C394 B.n341 VSUBS 0.018372f
C395 B.n342 VSUBS 0.016935f
C396 B.n343 VSUBS 0.007503f
C397 B.n344 VSUBS 0.007503f
C398 B.n345 VSUBS 0.007503f
C399 B.n346 VSUBS 0.007503f
C400 B.n347 VSUBS 0.007503f
C401 B.n348 VSUBS 0.007503f
C402 B.n349 VSUBS 0.007503f
C403 B.n350 VSUBS 0.007503f
C404 B.n351 VSUBS 0.007503f
C405 B.n352 VSUBS 0.007503f
C406 B.n353 VSUBS 0.007503f
C407 B.n354 VSUBS 0.007503f
C408 B.n355 VSUBS 0.007503f
C409 B.n356 VSUBS 0.007503f
C410 B.n357 VSUBS 0.007503f
C411 B.n358 VSUBS 0.007503f
C412 B.n359 VSUBS 0.007503f
C413 B.n360 VSUBS 0.007503f
C414 B.n361 VSUBS 0.007503f
C415 B.n362 VSUBS 0.007503f
C416 B.n363 VSUBS 0.007503f
C417 B.n364 VSUBS 0.007503f
C418 B.n365 VSUBS 0.007503f
C419 B.n366 VSUBS 0.007503f
C420 B.n367 VSUBS 0.007503f
C421 B.n368 VSUBS 0.007503f
C422 B.n369 VSUBS 0.007503f
C423 B.n370 VSUBS 0.007503f
C424 B.n371 VSUBS 0.007503f
C425 B.n372 VSUBS 0.007503f
C426 B.n373 VSUBS 0.007503f
C427 B.n374 VSUBS 0.007503f
C428 B.n375 VSUBS 0.009791f
C429 B.n376 VSUBS 0.01043f
C430 B.n377 VSUBS 0.02074f
C431 VDD1.t1 VSUBS 0.050913f
C432 VDD1.t0 VSUBS 0.050913f
C433 VDD1.n0 VSUBS 0.287835f
C434 VDD1.t2 VSUBS 0.050913f
C435 VDD1.t3 VSUBS 0.050913f
C436 VDD1.n1 VSUBS 0.458979f
C437 VTAIL.t1 VSUBS 0.363681f
C438 VTAIL.n0 VSUBS 0.355725f
C439 VTAIL.t6 VSUBS 0.363681f
C440 VTAIL.n1 VSUBS 0.396003f
C441 VTAIL.t7 VSUBS 0.363681f
C442 VTAIL.n2 VSUBS 0.876635f
C443 VTAIL.t3 VSUBS 0.363683f
C444 VTAIL.n3 VSUBS 0.876633f
C445 VTAIL.t0 VSUBS 0.363683f
C446 VTAIL.n4 VSUBS 0.396001f
C447 VTAIL.t4 VSUBS 0.363683f
C448 VTAIL.n5 VSUBS 0.396001f
C449 VTAIL.t5 VSUBS 0.363681f
C450 VTAIL.n6 VSUBS 0.876635f
C451 VTAIL.t2 VSUBS 0.363681f
C452 VTAIL.n7 VSUBS 0.829706f
C453 VP.n0 VSUBS 0.041665f
C454 VP.t0 VSUBS 0.554864f
C455 VP.n1 VSUBS 0.061088f
C456 VP.t2 VSUBS 0.703281f
C457 VP.t3 VSUBS 0.701929f
C458 VP.n2 VSUBS 1.70795f
C459 VP.n3 VSUBS 1.79698f
C460 VP.t1 VSUBS 0.554864f
C461 VP.n4 VSUBS 0.318046f
C462 VP.n5 VSUBS 0.049913f
C463 VP.n6 VSUBS 0.041665f
C464 VP.n7 VSUBS 0.041665f
C465 VP.n8 VSUBS 0.041665f
C466 VP.n9 VSUBS 0.061088f
C467 VP.n10 VSUBS 0.049913f
C468 VP.n11 VSUBS 0.318046f
C469 VP.n12 VSUBS 0.040607f
.ends

