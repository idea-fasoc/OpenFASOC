* NGSPICE file created from diff_pair_sample_0428.ext - technology: sky130A

.subckt diff_pair_sample_0428 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 w_n1734_n3764# sky130_fd_pr__pfet_01v8 ad=5.4522 pd=28.74 as=5.4522 ps=28.74 w=13.98 l=1.58
X1 VDD1.t1 VP.t0 VTAIL.t1 w_n1734_n3764# sky130_fd_pr__pfet_01v8 ad=5.4522 pd=28.74 as=5.4522 ps=28.74 w=13.98 l=1.58
X2 VDD1.t0 VP.t1 VTAIL.t0 w_n1734_n3764# sky130_fd_pr__pfet_01v8 ad=5.4522 pd=28.74 as=5.4522 ps=28.74 w=13.98 l=1.58
X3 B.t11 B.t9 B.t10 w_n1734_n3764# sky130_fd_pr__pfet_01v8 ad=5.4522 pd=28.74 as=0 ps=0 w=13.98 l=1.58
X4 VDD2.t0 VN.t1 VTAIL.t3 w_n1734_n3764# sky130_fd_pr__pfet_01v8 ad=5.4522 pd=28.74 as=5.4522 ps=28.74 w=13.98 l=1.58
X5 B.t8 B.t6 B.t7 w_n1734_n3764# sky130_fd_pr__pfet_01v8 ad=5.4522 pd=28.74 as=0 ps=0 w=13.98 l=1.58
X6 B.t5 B.t3 B.t4 w_n1734_n3764# sky130_fd_pr__pfet_01v8 ad=5.4522 pd=28.74 as=0 ps=0 w=13.98 l=1.58
X7 B.t2 B.t0 B.t1 w_n1734_n3764# sky130_fd_pr__pfet_01v8 ad=5.4522 pd=28.74 as=0 ps=0 w=13.98 l=1.58
R0 VN VN.t1 362.748
R1 VN VN.t0 319.156
R2 VTAIL.n306 VTAIL.n234 756.745
R3 VTAIL.n72 VTAIL.n0 756.745
R4 VTAIL.n228 VTAIL.n156 756.745
R5 VTAIL.n150 VTAIL.n78 756.745
R6 VTAIL.n258 VTAIL.n257 585
R7 VTAIL.n263 VTAIL.n262 585
R8 VTAIL.n265 VTAIL.n264 585
R9 VTAIL.n254 VTAIL.n253 585
R10 VTAIL.n271 VTAIL.n270 585
R11 VTAIL.n273 VTAIL.n272 585
R12 VTAIL.n250 VTAIL.n249 585
R13 VTAIL.n279 VTAIL.n278 585
R14 VTAIL.n281 VTAIL.n280 585
R15 VTAIL.n246 VTAIL.n245 585
R16 VTAIL.n287 VTAIL.n286 585
R17 VTAIL.n289 VTAIL.n288 585
R18 VTAIL.n242 VTAIL.n241 585
R19 VTAIL.n295 VTAIL.n294 585
R20 VTAIL.n297 VTAIL.n296 585
R21 VTAIL.n238 VTAIL.n237 585
R22 VTAIL.n304 VTAIL.n303 585
R23 VTAIL.n305 VTAIL.n236 585
R24 VTAIL.n307 VTAIL.n306 585
R25 VTAIL.n24 VTAIL.n23 585
R26 VTAIL.n29 VTAIL.n28 585
R27 VTAIL.n31 VTAIL.n30 585
R28 VTAIL.n20 VTAIL.n19 585
R29 VTAIL.n37 VTAIL.n36 585
R30 VTAIL.n39 VTAIL.n38 585
R31 VTAIL.n16 VTAIL.n15 585
R32 VTAIL.n45 VTAIL.n44 585
R33 VTAIL.n47 VTAIL.n46 585
R34 VTAIL.n12 VTAIL.n11 585
R35 VTAIL.n53 VTAIL.n52 585
R36 VTAIL.n55 VTAIL.n54 585
R37 VTAIL.n8 VTAIL.n7 585
R38 VTAIL.n61 VTAIL.n60 585
R39 VTAIL.n63 VTAIL.n62 585
R40 VTAIL.n4 VTAIL.n3 585
R41 VTAIL.n70 VTAIL.n69 585
R42 VTAIL.n71 VTAIL.n2 585
R43 VTAIL.n73 VTAIL.n72 585
R44 VTAIL.n229 VTAIL.n228 585
R45 VTAIL.n227 VTAIL.n158 585
R46 VTAIL.n226 VTAIL.n225 585
R47 VTAIL.n161 VTAIL.n159 585
R48 VTAIL.n220 VTAIL.n219 585
R49 VTAIL.n218 VTAIL.n217 585
R50 VTAIL.n165 VTAIL.n164 585
R51 VTAIL.n212 VTAIL.n211 585
R52 VTAIL.n210 VTAIL.n209 585
R53 VTAIL.n169 VTAIL.n168 585
R54 VTAIL.n204 VTAIL.n203 585
R55 VTAIL.n202 VTAIL.n201 585
R56 VTAIL.n173 VTAIL.n172 585
R57 VTAIL.n196 VTAIL.n195 585
R58 VTAIL.n194 VTAIL.n193 585
R59 VTAIL.n177 VTAIL.n176 585
R60 VTAIL.n188 VTAIL.n187 585
R61 VTAIL.n186 VTAIL.n185 585
R62 VTAIL.n181 VTAIL.n180 585
R63 VTAIL.n151 VTAIL.n150 585
R64 VTAIL.n149 VTAIL.n80 585
R65 VTAIL.n148 VTAIL.n147 585
R66 VTAIL.n83 VTAIL.n81 585
R67 VTAIL.n142 VTAIL.n141 585
R68 VTAIL.n140 VTAIL.n139 585
R69 VTAIL.n87 VTAIL.n86 585
R70 VTAIL.n134 VTAIL.n133 585
R71 VTAIL.n132 VTAIL.n131 585
R72 VTAIL.n91 VTAIL.n90 585
R73 VTAIL.n126 VTAIL.n125 585
R74 VTAIL.n124 VTAIL.n123 585
R75 VTAIL.n95 VTAIL.n94 585
R76 VTAIL.n118 VTAIL.n117 585
R77 VTAIL.n116 VTAIL.n115 585
R78 VTAIL.n99 VTAIL.n98 585
R79 VTAIL.n110 VTAIL.n109 585
R80 VTAIL.n108 VTAIL.n107 585
R81 VTAIL.n103 VTAIL.n102 585
R82 VTAIL.n259 VTAIL.t2 327.466
R83 VTAIL.n25 VTAIL.t1 327.466
R84 VTAIL.n182 VTAIL.t0 327.466
R85 VTAIL.n104 VTAIL.t3 327.466
R86 VTAIL.n263 VTAIL.n257 171.744
R87 VTAIL.n264 VTAIL.n263 171.744
R88 VTAIL.n264 VTAIL.n253 171.744
R89 VTAIL.n271 VTAIL.n253 171.744
R90 VTAIL.n272 VTAIL.n271 171.744
R91 VTAIL.n272 VTAIL.n249 171.744
R92 VTAIL.n279 VTAIL.n249 171.744
R93 VTAIL.n280 VTAIL.n279 171.744
R94 VTAIL.n280 VTAIL.n245 171.744
R95 VTAIL.n287 VTAIL.n245 171.744
R96 VTAIL.n288 VTAIL.n287 171.744
R97 VTAIL.n288 VTAIL.n241 171.744
R98 VTAIL.n295 VTAIL.n241 171.744
R99 VTAIL.n296 VTAIL.n295 171.744
R100 VTAIL.n296 VTAIL.n237 171.744
R101 VTAIL.n304 VTAIL.n237 171.744
R102 VTAIL.n305 VTAIL.n304 171.744
R103 VTAIL.n306 VTAIL.n305 171.744
R104 VTAIL.n29 VTAIL.n23 171.744
R105 VTAIL.n30 VTAIL.n29 171.744
R106 VTAIL.n30 VTAIL.n19 171.744
R107 VTAIL.n37 VTAIL.n19 171.744
R108 VTAIL.n38 VTAIL.n37 171.744
R109 VTAIL.n38 VTAIL.n15 171.744
R110 VTAIL.n45 VTAIL.n15 171.744
R111 VTAIL.n46 VTAIL.n45 171.744
R112 VTAIL.n46 VTAIL.n11 171.744
R113 VTAIL.n53 VTAIL.n11 171.744
R114 VTAIL.n54 VTAIL.n53 171.744
R115 VTAIL.n54 VTAIL.n7 171.744
R116 VTAIL.n61 VTAIL.n7 171.744
R117 VTAIL.n62 VTAIL.n61 171.744
R118 VTAIL.n62 VTAIL.n3 171.744
R119 VTAIL.n70 VTAIL.n3 171.744
R120 VTAIL.n71 VTAIL.n70 171.744
R121 VTAIL.n72 VTAIL.n71 171.744
R122 VTAIL.n228 VTAIL.n227 171.744
R123 VTAIL.n227 VTAIL.n226 171.744
R124 VTAIL.n226 VTAIL.n159 171.744
R125 VTAIL.n219 VTAIL.n159 171.744
R126 VTAIL.n219 VTAIL.n218 171.744
R127 VTAIL.n218 VTAIL.n164 171.744
R128 VTAIL.n211 VTAIL.n164 171.744
R129 VTAIL.n211 VTAIL.n210 171.744
R130 VTAIL.n210 VTAIL.n168 171.744
R131 VTAIL.n203 VTAIL.n168 171.744
R132 VTAIL.n203 VTAIL.n202 171.744
R133 VTAIL.n202 VTAIL.n172 171.744
R134 VTAIL.n195 VTAIL.n172 171.744
R135 VTAIL.n195 VTAIL.n194 171.744
R136 VTAIL.n194 VTAIL.n176 171.744
R137 VTAIL.n187 VTAIL.n176 171.744
R138 VTAIL.n187 VTAIL.n186 171.744
R139 VTAIL.n186 VTAIL.n180 171.744
R140 VTAIL.n150 VTAIL.n149 171.744
R141 VTAIL.n149 VTAIL.n148 171.744
R142 VTAIL.n148 VTAIL.n81 171.744
R143 VTAIL.n141 VTAIL.n81 171.744
R144 VTAIL.n141 VTAIL.n140 171.744
R145 VTAIL.n140 VTAIL.n86 171.744
R146 VTAIL.n133 VTAIL.n86 171.744
R147 VTAIL.n133 VTAIL.n132 171.744
R148 VTAIL.n132 VTAIL.n90 171.744
R149 VTAIL.n125 VTAIL.n90 171.744
R150 VTAIL.n125 VTAIL.n124 171.744
R151 VTAIL.n124 VTAIL.n94 171.744
R152 VTAIL.n117 VTAIL.n94 171.744
R153 VTAIL.n117 VTAIL.n116 171.744
R154 VTAIL.n116 VTAIL.n98 171.744
R155 VTAIL.n109 VTAIL.n98 171.744
R156 VTAIL.n109 VTAIL.n108 171.744
R157 VTAIL.n108 VTAIL.n102 171.744
R158 VTAIL.t2 VTAIL.n257 85.8723
R159 VTAIL.t1 VTAIL.n23 85.8723
R160 VTAIL.t0 VTAIL.n180 85.8723
R161 VTAIL.t3 VTAIL.n102 85.8723
R162 VTAIL.n311 VTAIL.n310 33.349
R163 VTAIL.n77 VTAIL.n76 33.349
R164 VTAIL.n233 VTAIL.n232 33.349
R165 VTAIL.n155 VTAIL.n154 33.349
R166 VTAIL.n155 VTAIL.n77 27.7117
R167 VTAIL.n311 VTAIL.n233 26.0652
R168 VTAIL.n259 VTAIL.n258 16.3895
R169 VTAIL.n25 VTAIL.n24 16.3895
R170 VTAIL.n182 VTAIL.n181 16.3895
R171 VTAIL.n104 VTAIL.n103 16.3895
R172 VTAIL.n307 VTAIL.n236 13.1884
R173 VTAIL.n73 VTAIL.n2 13.1884
R174 VTAIL.n229 VTAIL.n158 13.1884
R175 VTAIL.n151 VTAIL.n80 13.1884
R176 VTAIL.n262 VTAIL.n261 12.8005
R177 VTAIL.n303 VTAIL.n302 12.8005
R178 VTAIL.n308 VTAIL.n234 12.8005
R179 VTAIL.n28 VTAIL.n27 12.8005
R180 VTAIL.n69 VTAIL.n68 12.8005
R181 VTAIL.n74 VTAIL.n0 12.8005
R182 VTAIL.n230 VTAIL.n156 12.8005
R183 VTAIL.n225 VTAIL.n160 12.8005
R184 VTAIL.n185 VTAIL.n184 12.8005
R185 VTAIL.n152 VTAIL.n78 12.8005
R186 VTAIL.n147 VTAIL.n82 12.8005
R187 VTAIL.n107 VTAIL.n106 12.8005
R188 VTAIL.n265 VTAIL.n256 12.0247
R189 VTAIL.n301 VTAIL.n238 12.0247
R190 VTAIL.n31 VTAIL.n22 12.0247
R191 VTAIL.n67 VTAIL.n4 12.0247
R192 VTAIL.n224 VTAIL.n161 12.0247
R193 VTAIL.n188 VTAIL.n179 12.0247
R194 VTAIL.n146 VTAIL.n83 12.0247
R195 VTAIL.n110 VTAIL.n101 12.0247
R196 VTAIL.n266 VTAIL.n254 11.249
R197 VTAIL.n298 VTAIL.n297 11.249
R198 VTAIL.n32 VTAIL.n20 11.249
R199 VTAIL.n64 VTAIL.n63 11.249
R200 VTAIL.n221 VTAIL.n220 11.249
R201 VTAIL.n189 VTAIL.n177 11.249
R202 VTAIL.n143 VTAIL.n142 11.249
R203 VTAIL.n111 VTAIL.n99 11.249
R204 VTAIL.n270 VTAIL.n269 10.4732
R205 VTAIL.n294 VTAIL.n240 10.4732
R206 VTAIL.n36 VTAIL.n35 10.4732
R207 VTAIL.n60 VTAIL.n6 10.4732
R208 VTAIL.n217 VTAIL.n163 10.4732
R209 VTAIL.n193 VTAIL.n192 10.4732
R210 VTAIL.n139 VTAIL.n85 10.4732
R211 VTAIL.n115 VTAIL.n114 10.4732
R212 VTAIL.n273 VTAIL.n252 9.69747
R213 VTAIL.n293 VTAIL.n242 9.69747
R214 VTAIL.n39 VTAIL.n18 9.69747
R215 VTAIL.n59 VTAIL.n8 9.69747
R216 VTAIL.n216 VTAIL.n165 9.69747
R217 VTAIL.n196 VTAIL.n175 9.69747
R218 VTAIL.n138 VTAIL.n87 9.69747
R219 VTAIL.n118 VTAIL.n97 9.69747
R220 VTAIL.n310 VTAIL.n309 9.45567
R221 VTAIL.n76 VTAIL.n75 9.45567
R222 VTAIL.n232 VTAIL.n231 9.45567
R223 VTAIL.n154 VTAIL.n153 9.45567
R224 VTAIL.n309 VTAIL.n308 9.3005
R225 VTAIL.n248 VTAIL.n247 9.3005
R226 VTAIL.n277 VTAIL.n276 9.3005
R227 VTAIL.n275 VTAIL.n274 9.3005
R228 VTAIL.n252 VTAIL.n251 9.3005
R229 VTAIL.n269 VTAIL.n268 9.3005
R230 VTAIL.n267 VTAIL.n266 9.3005
R231 VTAIL.n256 VTAIL.n255 9.3005
R232 VTAIL.n261 VTAIL.n260 9.3005
R233 VTAIL.n283 VTAIL.n282 9.3005
R234 VTAIL.n285 VTAIL.n284 9.3005
R235 VTAIL.n244 VTAIL.n243 9.3005
R236 VTAIL.n291 VTAIL.n290 9.3005
R237 VTAIL.n293 VTAIL.n292 9.3005
R238 VTAIL.n240 VTAIL.n239 9.3005
R239 VTAIL.n299 VTAIL.n298 9.3005
R240 VTAIL.n301 VTAIL.n300 9.3005
R241 VTAIL.n302 VTAIL.n235 9.3005
R242 VTAIL.n75 VTAIL.n74 9.3005
R243 VTAIL.n14 VTAIL.n13 9.3005
R244 VTAIL.n43 VTAIL.n42 9.3005
R245 VTAIL.n41 VTAIL.n40 9.3005
R246 VTAIL.n18 VTAIL.n17 9.3005
R247 VTAIL.n35 VTAIL.n34 9.3005
R248 VTAIL.n33 VTAIL.n32 9.3005
R249 VTAIL.n22 VTAIL.n21 9.3005
R250 VTAIL.n27 VTAIL.n26 9.3005
R251 VTAIL.n49 VTAIL.n48 9.3005
R252 VTAIL.n51 VTAIL.n50 9.3005
R253 VTAIL.n10 VTAIL.n9 9.3005
R254 VTAIL.n57 VTAIL.n56 9.3005
R255 VTAIL.n59 VTAIL.n58 9.3005
R256 VTAIL.n6 VTAIL.n5 9.3005
R257 VTAIL.n65 VTAIL.n64 9.3005
R258 VTAIL.n67 VTAIL.n66 9.3005
R259 VTAIL.n68 VTAIL.n1 9.3005
R260 VTAIL.n208 VTAIL.n207 9.3005
R261 VTAIL.n167 VTAIL.n166 9.3005
R262 VTAIL.n214 VTAIL.n213 9.3005
R263 VTAIL.n216 VTAIL.n215 9.3005
R264 VTAIL.n163 VTAIL.n162 9.3005
R265 VTAIL.n222 VTAIL.n221 9.3005
R266 VTAIL.n224 VTAIL.n223 9.3005
R267 VTAIL.n160 VTAIL.n157 9.3005
R268 VTAIL.n231 VTAIL.n230 9.3005
R269 VTAIL.n206 VTAIL.n205 9.3005
R270 VTAIL.n171 VTAIL.n170 9.3005
R271 VTAIL.n200 VTAIL.n199 9.3005
R272 VTAIL.n198 VTAIL.n197 9.3005
R273 VTAIL.n175 VTAIL.n174 9.3005
R274 VTAIL.n192 VTAIL.n191 9.3005
R275 VTAIL.n190 VTAIL.n189 9.3005
R276 VTAIL.n179 VTAIL.n178 9.3005
R277 VTAIL.n184 VTAIL.n183 9.3005
R278 VTAIL.n130 VTAIL.n129 9.3005
R279 VTAIL.n89 VTAIL.n88 9.3005
R280 VTAIL.n136 VTAIL.n135 9.3005
R281 VTAIL.n138 VTAIL.n137 9.3005
R282 VTAIL.n85 VTAIL.n84 9.3005
R283 VTAIL.n144 VTAIL.n143 9.3005
R284 VTAIL.n146 VTAIL.n145 9.3005
R285 VTAIL.n82 VTAIL.n79 9.3005
R286 VTAIL.n153 VTAIL.n152 9.3005
R287 VTAIL.n128 VTAIL.n127 9.3005
R288 VTAIL.n93 VTAIL.n92 9.3005
R289 VTAIL.n122 VTAIL.n121 9.3005
R290 VTAIL.n120 VTAIL.n119 9.3005
R291 VTAIL.n97 VTAIL.n96 9.3005
R292 VTAIL.n114 VTAIL.n113 9.3005
R293 VTAIL.n112 VTAIL.n111 9.3005
R294 VTAIL.n101 VTAIL.n100 9.3005
R295 VTAIL.n106 VTAIL.n105 9.3005
R296 VTAIL.n274 VTAIL.n250 8.92171
R297 VTAIL.n290 VTAIL.n289 8.92171
R298 VTAIL.n40 VTAIL.n16 8.92171
R299 VTAIL.n56 VTAIL.n55 8.92171
R300 VTAIL.n213 VTAIL.n212 8.92171
R301 VTAIL.n197 VTAIL.n173 8.92171
R302 VTAIL.n135 VTAIL.n134 8.92171
R303 VTAIL.n119 VTAIL.n95 8.92171
R304 VTAIL.n278 VTAIL.n277 8.14595
R305 VTAIL.n286 VTAIL.n244 8.14595
R306 VTAIL.n44 VTAIL.n43 8.14595
R307 VTAIL.n52 VTAIL.n10 8.14595
R308 VTAIL.n209 VTAIL.n167 8.14595
R309 VTAIL.n201 VTAIL.n200 8.14595
R310 VTAIL.n131 VTAIL.n89 8.14595
R311 VTAIL.n123 VTAIL.n122 8.14595
R312 VTAIL.n281 VTAIL.n248 7.3702
R313 VTAIL.n285 VTAIL.n246 7.3702
R314 VTAIL.n47 VTAIL.n14 7.3702
R315 VTAIL.n51 VTAIL.n12 7.3702
R316 VTAIL.n208 VTAIL.n169 7.3702
R317 VTAIL.n204 VTAIL.n171 7.3702
R318 VTAIL.n130 VTAIL.n91 7.3702
R319 VTAIL.n126 VTAIL.n93 7.3702
R320 VTAIL.n282 VTAIL.n281 6.59444
R321 VTAIL.n282 VTAIL.n246 6.59444
R322 VTAIL.n48 VTAIL.n47 6.59444
R323 VTAIL.n48 VTAIL.n12 6.59444
R324 VTAIL.n205 VTAIL.n169 6.59444
R325 VTAIL.n205 VTAIL.n204 6.59444
R326 VTAIL.n127 VTAIL.n91 6.59444
R327 VTAIL.n127 VTAIL.n126 6.59444
R328 VTAIL.n278 VTAIL.n248 5.81868
R329 VTAIL.n286 VTAIL.n285 5.81868
R330 VTAIL.n44 VTAIL.n14 5.81868
R331 VTAIL.n52 VTAIL.n51 5.81868
R332 VTAIL.n209 VTAIL.n208 5.81868
R333 VTAIL.n201 VTAIL.n171 5.81868
R334 VTAIL.n131 VTAIL.n130 5.81868
R335 VTAIL.n123 VTAIL.n93 5.81868
R336 VTAIL.n277 VTAIL.n250 5.04292
R337 VTAIL.n289 VTAIL.n244 5.04292
R338 VTAIL.n43 VTAIL.n16 5.04292
R339 VTAIL.n55 VTAIL.n10 5.04292
R340 VTAIL.n212 VTAIL.n167 5.04292
R341 VTAIL.n200 VTAIL.n173 5.04292
R342 VTAIL.n134 VTAIL.n89 5.04292
R343 VTAIL.n122 VTAIL.n95 5.04292
R344 VTAIL.n274 VTAIL.n273 4.26717
R345 VTAIL.n290 VTAIL.n242 4.26717
R346 VTAIL.n40 VTAIL.n39 4.26717
R347 VTAIL.n56 VTAIL.n8 4.26717
R348 VTAIL.n213 VTAIL.n165 4.26717
R349 VTAIL.n197 VTAIL.n196 4.26717
R350 VTAIL.n135 VTAIL.n87 4.26717
R351 VTAIL.n119 VTAIL.n118 4.26717
R352 VTAIL.n260 VTAIL.n259 3.70982
R353 VTAIL.n26 VTAIL.n25 3.70982
R354 VTAIL.n183 VTAIL.n182 3.70982
R355 VTAIL.n105 VTAIL.n104 3.70982
R356 VTAIL.n270 VTAIL.n252 3.49141
R357 VTAIL.n294 VTAIL.n293 3.49141
R358 VTAIL.n36 VTAIL.n18 3.49141
R359 VTAIL.n60 VTAIL.n59 3.49141
R360 VTAIL.n217 VTAIL.n216 3.49141
R361 VTAIL.n193 VTAIL.n175 3.49141
R362 VTAIL.n139 VTAIL.n138 3.49141
R363 VTAIL.n115 VTAIL.n97 3.49141
R364 VTAIL.n269 VTAIL.n254 2.71565
R365 VTAIL.n297 VTAIL.n240 2.71565
R366 VTAIL.n35 VTAIL.n20 2.71565
R367 VTAIL.n63 VTAIL.n6 2.71565
R368 VTAIL.n220 VTAIL.n163 2.71565
R369 VTAIL.n192 VTAIL.n177 2.71565
R370 VTAIL.n142 VTAIL.n85 2.71565
R371 VTAIL.n114 VTAIL.n99 2.71565
R372 VTAIL.n266 VTAIL.n265 1.93989
R373 VTAIL.n298 VTAIL.n238 1.93989
R374 VTAIL.n32 VTAIL.n31 1.93989
R375 VTAIL.n64 VTAIL.n4 1.93989
R376 VTAIL.n221 VTAIL.n161 1.93989
R377 VTAIL.n189 VTAIL.n188 1.93989
R378 VTAIL.n143 VTAIL.n83 1.93989
R379 VTAIL.n111 VTAIL.n110 1.93989
R380 VTAIL.n233 VTAIL.n155 1.2936
R381 VTAIL.n262 VTAIL.n256 1.16414
R382 VTAIL.n303 VTAIL.n301 1.16414
R383 VTAIL.n310 VTAIL.n234 1.16414
R384 VTAIL.n28 VTAIL.n22 1.16414
R385 VTAIL.n69 VTAIL.n67 1.16414
R386 VTAIL.n76 VTAIL.n0 1.16414
R387 VTAIL.n232 VTAIL.n156 1.16414
R388 VTAIL.n225 VTAIL.n224 1.16414
R389 VTAIL.n185 VTAIL.n179 1.16414
R390 VTAIL.n154 VTAIL.n78 1.16414
R391 VTAIL.n147 VTAIL.n146 1.16414
R392 VTAIL.n107 VTAIL.n101 1.16414
R393 VTAIL VTAIL.n77 0.940155
R394 VTAIL.n261 VTAIL.n258 0.388379
R395 VTAIL.n302 VTAIL.n236 0.388379
R396 VTAIL.n308 VTAIL.n307 0.388379
R397 VTAIL.n27 VTAIL.n24 0.388379
R398 VTAIL.n68 VTAIL.n2 0.388379
R399 VTAIL.n74 VTAIL.n73 0.388379
R400 VTAIL.n230 VTAIL.n229 0.388379
R401 VTAIL.n160 VTAIL.n158 0.388379
R402 VTAIL.n184 VTAIL.n181 0.388379
R403 VTAIL.n152 VTAIL.n151 0.388379
R404 VTAIL.n82 VTAIL.n80 0.388379
R405 VTAIL.n106 VTAIL.n103 0.388379
R406 VTAIL VTAIL.n311 0.353948
R407 VTAIL.n260 VTAIL.n255 0.155672
R408 VTAIL.n267 VTAIL.n255 0.155672
R409 VTAIL.n268 VTAIL.n267 0.155672
R410 VTAIL.n268 VTAIL.n251 0.155672
R411 VTAIL.n275 VTAIL.n251 0.155672
R412 VTAIL.n276 VTAIL.n275 0.155672
R413 VTAIL.n276 VTAIL.n247 0.155672
R414 VTAIL.n283 VTAIL.n247 0.155672
R415 VTAIL.n284 VTAIL.n283 0.155672
R416 VTAIL.n284 VTAIL.n243 0.155672
R417 VTAIL.n291 VTAIL.n243 0.155672
R418 VTAIL.n292 VTAIL.n291 0.155672
R419 VTAIL.n292 VTAIL.n239 0.155672
R420 VTAIL.n299 VTAIL.n239 0.155672
R421 VTAIL.n300 VTAIL.n299 0.155672
R422 VTAIL.n300 VTAIL.n235 0.155672
R423 VTAIL.n309 VTAIL.n235 0.155672
R424 VTAIL.n26 VTAIL.n21 0.155672
R425 VTAIL.n33 VTAIL.n21 0.155672
R426 VTAIL.n34 VTAIL.n33 0.155672
R427 VTAIL.n34 VTAIL.n17 0.155672
R428 VTAIL.n41 VTAIL.n17 0.155672
R429 VTAIL.n42 VTAIL.n41 0.155672
R430 VTAIL.n42 VTAIL.n13 0.155672
R431 VTAIL.n49 VTAIL.n13 0.155672
R432 VTAIL.n50 VTAIL.n49 0.155672
R433 VTAIL.n50 VTAIL.n9 0.155672
R434 VTAIL.n57 VTAIL.n9 0.155672
R435 VTAIL.n58 VTAIL.n57 0.155672
R436 VTAIL.n58 VTAIL.n5 0.155672
R437 VTAIL.n65 VTAIL.n5 0.155672
R438 VTAIL.n66 VTAIL.n65 0.155672
R439 VTAIL.n66 VTAIL.n1 0.155672
R440 VTAIL.n75 VTAIL.n1 0.155672
R441 VTAIL.n231 VTAIL.n157 0.155672
R442 VTAIL.n223 VTAIL.n157 0.155672
R443 VTAIL.n223 VTAIL.n222 0.155672
R444 VTAIL.n222 VTAIL.n162 0.155672
R445 VTAIL.n215 VTAIL.n162 0.155672
R446 VTAIL.n215 VTAIL.n214 0.155672
R447 VTAIL.n214 VTAIL.n166 0.155672
R448 VTAIL.n207 VTAIL.n166 0.155672
R449 VTAIL.n207 VTAIL.n206 0.155672
R450 VTAIL.n206 VTAIL.n170 0.155672
R451 VTAIL.n199 VTAIL.n170 0.155672
R452 VTAIL.n199 VTAIL.n198 0.155672
R453 VTAIL.n198 VTAIL.n174 0.155672
R454 VTAIL.n191 VTAIL.n174 0.155672
R455 VTAIL.n191 VTAIL.n190 0.155672
R456 VTAIL.n190 VTAIL.n178 0.155672
R457 VTAIL.n183 VTAIL.n178 0.155672
R458 VTAIL.n153 VTAIL.n79 0.155672
R459 VTAIL.n145 VTAIL.n79 0.155672
R460 VTAIL.n145 VTAIL.n144 0.155672
R461 VTAIL.n144 VTAIL.n84 0.155672
R462 VTAIL.n137 VTAIL.n84 0.155672
R463 VTAIL.n137 VTAIL.n136 0.155672
R464 VTAIL.n136 VTAIL.n88 0.155672
R465 VTAIL.n129 VTAIL.n88 0.155672
R466 VTAIL.n129 VTAIL.n128 0.155672
R467 VTAIL.n128 VTAIL.n92 0.155672
R468 VTAIL.n121 VTAIL.n92 0.155672
R469 VTAIL.n121 VTAIL.n120 0.155672
R470 VTAIL.n120 VTAIL.n96 0.155672
R471 VTAIL.n113 VTAIL.n96 0.155672
R472 VTAIL.n113 VTAIL.n112 0.155672
R473 VTAIL.n112 VTAIL.n100 0.155672
R474 VTAIL.n105 VTAIL.n100 0.155672
R475 VDD2.n149 VDD2.n77 756.745
R476 VDD2.n72 VDD2.n0 756.745
R477 VDD2.n150 VDD2.n149 585
R478 VDD2.n148 VDD2.n79 585
R479 VDD2.n147 VDD2.n146 585
R480 VDD2.n82 VDD2.n80 585
R481 VDD2.n141 VDD2.n140 585
R482 VDD2.n139 VDD2.n138 585
R483 VDD2.n86 VDD2.n85 585
R484 VDD2.n133 VDD2.n132 585
R485 VDD2.n131 VDD2.n130 585
R486 VDD2.n90 VDD2.n89 585
R487 VDD2.n125 VDD2.n124 585
R488 VDD2.n123 VDD2.n122 585
R489 VDD2.n94 VDD2.n93 585
R490 VDD2.n117 VDD2.n116 585
R491 VDD2.n115 VDD2.n114 585
R492 VDD2.n98 VDD2.n97 585
R493 VDD2.n109 VDD2.n108 585
R494 VDD2.n107 VDD2.n106 585
R495 VDD2.n102 VDD2.n101 585
R496 VDD2.n24 VDD2.n23 585
R497 VDD2.n29 VDD2.n28 585
R498 VDD2.n31 VDD2.n30 585
R499 VDD2.n20 VDD2.n19 585
R500 VDD2.n37 VDD2.n36 585
R501 VDD2.n39 VDD2.n38 585
R502 VDD2.n16 VDD2.n15 585
R503 VDD2.n45 VDD2.n44 585
R504 VDD2.n47 VDD2.n46 585
R505 VDD2.n12 VDD2.n11 585
R506 VDD2.n53 VDD2.n52 585
R507 VDD2.n55 VDD2.n54 585
R508 VDD2.n8 VDD2.n7 585
R509 VDD2.n61 VDD2.n60 585
R510 VDD2.n63 VDD2.n62 585
R511 VDD2.n4 VDD2.n3 585
R512 VDD2.n70 VDD2.n69 585
R513 VDD2.n71 VDD2.n2 585
R514 VDD2.n73 VDD2.n72 585
R515 VDD2.n103 VDD2.t0 327.466
R516 VDD2.n25 VDD2.t1 327.466
R517 VDD2.n149 VDD2.n148 171.744
R518 VDD2.n148 VDD2.n147 171.744
R519 VDD2.n147 VDD2.n80 171.744
R520 VDD2.n140 VDD2.n80 171.744
R521 VDD2.n140 VDD2.n139 171.744
R522 VDD2.n139 VDD2.n85 171.744
R523 VDD2.n132 VDD2.n85 171.744
R524 VDD2.n132 VDD2.n131 171.744
R525 VDD2.n131 VDD2.n89 171.744
R526 VDD2.n124 VDD2.n89 171.744
R527 VDD2.n124 VDD2.n123 171.744
R528 VDD2.n123 VDD2.n93 171.744
R529 VDD2.n116 VDD2.n93 171.744
R530 VDD2.n116 VDD2.n115 171.744
R531 VDD2.n115 VDD2.n97 171.744
R532 VDD2.n108 VDD2.n97 171.744
R533 VDD2.n108 VDD2.n107 171.744
R534 VDD2.n107 VDD2.n101 171.744
R535 VDD2.n29 VDD2.n23 171.744
R536 VDD2.n30 VDD2.n29 171.744
R537 VDD2.n30 VDD2.n19 171.744
R538 VDD2.n37 VDD2.n19 171.744
R539 VDD2.n38 VDD2.n37 171.744
R540 VDD2.n38 VDD2.n15 171.744
R541 VDD2.n45 VDD2.n15 171.744
R542 VDD2.n46 VDD2.n45 171.744
R543 VDD2.n46 VDD2.n11 171.744
R544 VDD2.n53 VDD2.n11 171.744
R545 VDD2.n54 VDD2.n53 171.744
R546 VDD2.n54 VDD2.n7 171.744
R547 VDD2.n61 VDD2.n7 171.744
R548 VDD2.n62 VDD2.n61 171.744
R549 VDD2.n62 VDD2.n3 171.744
R550 VDD2.n70 VDD2.n3 171.744
R551 VDD2.n71 VDD2.n70 171.744
R552 VDD2.n72 VDD2.n71 171.744
R553 VDD2.n154 VDD2.n76 89.0321
R554 VDD2.t0 VDD2.n101 85.8723
R555 VDD2.t1 VDD2.n23 85.8723
R556 VDD2.n154 VDD2.n153 50.0278
R557 VDD2.n103 VDD2.n102 16.3895
R558 VDD2.n25 VDD2.n24 16.3895
R559 VDD2.n150 VDD2.n79 13.1884
R560 VDD2.n73 VDD2.n2 13.1884
R561 VDD2.n151 VDD2.n77 12.8005
R562 VDD2.n146 VDD2.n81 12.8005
R563 VDD2.n106 VDD2.n105 12.8005
R564 VDD2.n28 VDD2.n27 12.8005
R565 VDD2.n69 VDD2.n68 12.8005
R566 VDD2.n74 VDD2.n0 12.8005
R567 VDD2.n145 VDD2.n82 12.0247
R568 VDD2.n109 VDD2.n100 12.0247
R569 VDD2.n31 VDD2.n22 12.0247
R570 VDD2.n67 VDD2.n4 12.0247
R571 VDD2.n142 VDD2.n141 11.249
R572 VDD2.n110 VDD2.n98 11.249
R573 VDD2.n32 VDD2.n20 11.249
R574 VDD2.n64 VDD2.n63 11.249
R575 VDD2.n138 VDD2.n84 10.4732
R576 VDD2.n114 VDD2.n113 10.4732
R577 VDD2.n36 VDD2.n35 10.4732
R578 VDD2.n60 VDD2.n6 10.4732
R579 VDD2.n137 VDD2.n86 9.69747
R580 VDD2.n117 VDD2.n96 9.69747
R581 VDD2.n39 VDD2.n18 9.69747
R582 VDD2.n59 VDD2.n8 9.69747
R583 VDD2.n153 VDD2.n152 9.45567
R584 VDD2.n76 VDD2.n75 9.45567
R585 VDD2.n129 VDD2.n128 9.3005
R586 VDD2.n88 VDD2.n87 9.3005
R587 VDD2.n135 VDD2.n134 9.3005
R588 VDD2.n137 VDD2.n136 9.3005
R589 VDD2.n84 VDD2.n83 9.3005
R590 VDD2.n143 VDD2.n142 9.3005
R591 VDD2.n145 VDD2.n144 9.3005
R592 VDD2.n81 VDD2.n78 9.3005
R593 VDD2.n152 VDD2.n151 9.3005
R594 VDD2.n127 VDD2.n126 9.3005
R595 VDD2.n92 VDD2.n91 9.3005
R596 VDD2.n121 VDD2.n120 9.3005
R597 VDD2.n119 VDD2.n118 9.3005
R598 VDD2.n96 VDD2.n95 9.3005
R599 VDD2.n113 VDD2.n112 9.3005
R600 VDD2.n111 VDD2.n110 9.3005
R601 VDD2.n100 VDD2.n99 9.3005
R602 VDD2.n105 VDD2.n104 9.3005
R603 VDD2.n75 VDD2.n74 9.3005
R604 VDD2.n14 VDD2.n13 9.3005
R605 VDD2.n43 VDD2.n42 9.3005
R606 VDD2.n41 VDD2.n40 9.3005
R607 VDD2.n18 VDD2.n17 9.3005
R608 VDD2.n35 VDD2.n34 9.3005
R609 VDD2.n33 VDD2.n32 9.3005
R610 VDD2.n22 VDD2.n21 9.3005
R611 VDD2.n27 VDD2.n26 9.3005
R612 VDD2.n49 VDD2.n48 9.3005
R613 VDD2.n51 VDD2.n50 9.3005
R614 VDD2.n10 VDD2.n9 9.3005
R615 VDD2.n57 VDD2.n56 9.3005
R616 VDD2.n59 VDD2.n58 9.3005
R617 VDD2.n6 VDD2.n5 9.3005
R618 VDD2.n65 VDD2.n64 9.3005
R619 VDD2.n67 VDD2.n66 9.3005
R620 VDD2.n68 VDD2.n1 9.3005
R621 VDD2.n134 VDD2.n133 8.92171
R622 VDD2.n118 VDD2.n94 8.92171
R623 VDD2.n40 VDD2.n16 8.92171
R624 VDD2.n56 VDD2.n55 8.92171
R625 VDD2.n130 VDD2.n88 8.14595
R626 VDD2.n122 VDD2.n121 8.14595
R627 VDD2.n44 VDD2.n43 8.14595
R628 VDD2.n52 VDD2.n10 8.14595
R629 VDD2.n129 VDD2.n90 7.3702
R630 VDD2.n125 VDD2.n92 7.3702
R631 VDD2.n47 VDD2.n14 7.3702
R632 VDD2.n51 VDD2.n12 7.3702
R633 VDD2.n126 VDD2.n90 6.59444
R634 VDD2.n126 VDD2.n125 6.59444
R635 VDD2.n48 VDD2.n47 6.59444
R636 VDD2.n48 VDD2.n12 6.59444
R637 VDD2.n130 VDD2.n129 5.81868
R638 VDD2.n122 VDD2.n92 5.81868
R639 VDD2.n44 VDD2.n14 5.81868
R640 VDD2.n52 VDD2.n51 5.81868
R641 VDD2.n133 VDD2.n88 5.04292
R642 VDD2.n121 VDD2.n94 5.04292
R643 VDD2.n43 VDD2.n16 5.04292
R644 VDD2.n55 VDD2.n10 5.04292
R645 VDD2.n134 VDD2.n86 4.26717
R646 VDD2.n118 VDD2.n117 4.26717
R647 VDD2.n40 VDD2.n39 4.26717
R648 VDD2.n56 VDD2.n8 4.26717
R649 VDD2.n104 VDD2.n103 3.70982
R650 VDD2.n26 VDD2.n25 3.70982
R651 VDD2.n138 VDD2.n137 3.49141
R652 VDD2.n114 VDD2.n96 3.49141
R653 VDD2.n36 VDD2.n18 3.49141
R654 VDD2.n60 VDD2.n59 3.49141
R655 VDD2.n141 VDD2.n84 2.71565
R656 VDD2.n113 VDD2.n98 2.71565
R657 VDD2.n35 VDD2.n20 2.71565
R658 VDD2.n63 VDD2.n6 2.71565
R659 VDD2.n142 VDD2.n82 1.93989
R660 VDD2.n110 VDD2.n109 1.93989
R661 VDD2.n32 VDD2.n31 1.93989
R662 VDD2.n64 VDD2.n4 1.93989
R663 VDD2.n153 VDD2.n77 1.16414
R664 VDD2.n146 VDD2.n145 1.16414
R665 VDD2.n106 VDD2.n100 1.16414
R666 VDD2.n28 VDD2.n22 1.16414
R667 VDD2.n69 VDD2.n67 1.16414
R668 VDD2.n76 VDD2.n0 1.16414
R669 VDD2 VDD2.n154 0.470328
R670 VDD2.n151 VDD2.n150 0.388379
R671 VDD2.n81 VDD2.n79 0.388379
R672 VDD2.n105 VDD2.n102 0.388379
R673 VDD2.n27 VDD2.n24 0.388379
R674 VDD2.n68 VDD2.n2 0.388379
R675 VDD2.n74 VDD2.n73 0.388379
R676 VDD2.n152 VDD2.n78 0.155672
R677 VDD2.n144 VDD2.n78 0.155672
R678 VDD2.n144 VDD2.n143 0.155672
R679 VDD2.n143 VDD2.n83 0.155672
R680 VDD2.n136 VDD2.n83 0.155672
R681 VDD2.n136 VDD2.n135 0.155672
R682 VDD2.n135 VDD2.n87 0.155672
R683 VDD2.n128 VDD2.n87 0.155672
R684 VDD2.n128 VDD2.n127 0.155672
R685 VDD2.n127 VDD2.n91 0.155672
R686 VDD2.n120 VDD2.n91 0.155672
R687 VDD2.n120 VDD2.n119 0.155672
R688 VDD2.n119 VDD2.n95 0.155672
R689 VDD2.n112 VDD2.n95 0.155672
R690 VDD2.n112 VDD2.n111 0.155672
R691 VDD2.n111 VDD2.n99 0.155672
R692 VDD2.n104 VDD2.n99 0.155672
R693 VDD2.n26 VDD2.n21 0.155672
R694 VDD2.n33 VDD2.n21 0.155672
R695 VDD2.n34 VDD2.n33 0.155672
R696 VDD2.n34 VDD2.n17 0.155672
R697 VDD2.n41 VDD2.n17 0.155672
R698 VDD2.n42 VDD2.n41 0.155672
R699 VDD2.n42 VDD2.n13 0.155672
R700 VDD2.n49 VDD2.n13 0.155672
R701 VDD2.n50 VDD2.n49 0.155672
R702 VDD2.n50 VDD2.n9 0.155672
R703 VDD2.n57 VDD2.n9 0.155672
R704 VDD2.n58 VDD2.n57 0.155672
R705 VDD2.n58 VDD2.n5 0.155672
R706 VDD2.n65 VDD2.n5 0.155672
R707 VDD2.n66 VDD2.n65 0.155672
R708 VDD2.n66 VDD2.n1 0.155672
R709 VDD2.n75 VDD2.n1 0.155672
R710 VP.n0 VP.t1 362.462
R711 VP.n0 VP.t0 319.01
R712 VP VP.n0 0.146778
R713 VDD1.n72 VDD1.n0 756.745
R714 VDD1.n149 VDD1.n77 756.745
R715 VDD1.n73 VDD1.n72 585
R716 VDD1.n71 VDD1.n2 585
R717 VDD1.n70 VDD1.n69 585
R718 VDD1.n5 VDD1.n3 585
R719 VDD1.n64 VDD1.n63 585
R720 VDD1.n62 VDD1.n61 585
R721 VDD1.n9 VDD1.n8 585
R722 VDD1.n56 VDD1.n55 585
R723 VDD1.n54 VDD1.n53 585
R724 VDD1.n13 VDD1.n12 585
R725 VDD1.n48 VDD1.n47 585
R726 VDD1.n46 VDD1.n45 585
R727 VDD1.n17 VDD1.n16 585
R728 VDD1.n40 VDD1.n39 585
R729 VDD1.n38 VDD1.n37 585
R730 VDD1.n21 VDD1.n20 585
R731 VDD1.n32 VDD1.n31 585
R732 VDD1.n30 VDD1.n29 585
R733 VDD1.n25 VDD1.n24 585
R734 VDD1.n101 VDD1.n100 585
R735 VDD1.n106 VDD1.n105 585
R736 VDD1.n108 VDD1.n107 585
R737 VDD1.n97 VDD1.n96 585
R738 VDD1.n114 VDD1.n113 585
R739 VDD1.n116 VDD1.n115 585
R740 VDD1.n93 VDD1.n92 585
R741 VDD1.n122 VDD1.n121 585
R742 VDD1.n124 VDD1.n123 585
R743 VDD1.n89 VDD1.n88 585
R744 VDD1.n130 VDD1.n129 585
R745 VDD1.n132 VDD1.n131 585
R746 VDD1.n85 VDD1.n84 585
R747 VDD1.n138 VDD1.n137 585
R748 VDD1.n140 VDD1.n139 585
R749 VDD1.n81 VDD1.n80 585
R750 VDD1.n147 VDD1.n146 585
R751 VDD1.n148 VDD1.n79 585
R752 VDD1.n150 VDD1.n149 585
R753 VDD1.n26 VDD1.t0 327.466
R754 VDD1.n102 VDD1.t1 327.466
R755 VDD1.n72 VDD1.n71 171.744
R756 VDD1.n71 VDD1.n70 171.744
R757 VDD1.n70 VDD1.n3 171.744
R758 VDD1.n63 VDD1.n3 171.744
R759 VDD1.n63 VDD1.n62 171.744
R760 VDD1.n62 VDD1.n8 171.744
R761 VDD1.n55 VDD1.n8 171.744
R762 VDD1.n55 VDD1.n54 171.744
R763 VDD1.n54 VDD1.n12 171.744
R764 VDD1.n47 VDD1.n12 171.744
R765 VDD1.n47 VDD1.n46 171.744
R766 VDD1.n46 VDD1.n16 171.744
R767 VDD1.n39 VDD1.n16 171.744
R768 VDD1.n39 VDD1.n38 171.744
R769 VDD1.n38 VDD1.n20 171.744
R770 VDD1.n31 VDD1.n20 171.744
R771 VDD1.n31 VDD1.n30 171.744
R772 VDD1.n30 VDD1.n24 171.744
R773 VDD1.n106 VDD1.n100 171.744
R774 VDD1.n107 VDD1.n106 171.744
R775 VDD1.n107 VDD1.n96 171.744
R776 VDD1.n114 VDD1.n96 171.744
R777 VDD1.n115 VDD1.n114 171.744
R778 VDD1.n115 VDD1.n92 171.744
R779 VDD1.n122 VDD1.n92 171.744
R780 VDD1.n123 VDD1.n122 171.744
R781 VDD1.n123 VDD1.n88 171.744
R782 VDD1.n130 VDD1.n88 171.744
R783 VDD1.n131 VDD1.n130 171.744
R784 VDD1.n131 VDD1.n84 171.744
R785 VDD1.n138 VDD1.n84 171.744
R786 VDD1.n139 VDD1.n138 171.744
R787 VDD1.n139 VDD1.n80 171.744
R788 VDD1.n147 VDD1.n80 171.744
R789 VDD1.n148 VDD1.n147 171.744
R790 VDD1.n149 VDD1.n148 171.744
R791 VDD1 VDD1.n153 89.9685
R792 VDD1.t0 VDD1.n24 85.8723
R793 VDD1.t1 VDD1.n100 85.8723
R794 VDD1 VDD1.n76 50.4976
R795 VDD1.n26 VDD1.n25 16.3895
R796 VDD1.n102 VDD1.n101 16.3895
R797 VDD1.n73 VDD1.n2 13.1884
R798 VDD1.n150 VDD1.n79 13.1884
R799 VDD1.n74 VDD1.n0 12.8005
R800 VDD1.n69 VDD1.n4 12.8005
R801 VDD1.n29 VDD1.n28 12.8005
R802 VDD1.n105 VDD1.n104 12.8005
R803 VDD1.n146 VDD1.n145 12.8005
R804 VDD1.n151 VDD1.n77 12.8005
R805 VDD1.n68 VDD1.n5 12.0247
R806 VDD1.n32 VDD1.n23 12.0247
R807 VDD1.n108 VDD1.n99 12.0247
R808 VDD1.n144 VDD1.n81 12.0247
R809 VDD1.n65 VDD1.n64 11.249
R810 VDD1.n33 VDD1.n21 11.249
R811 VDD1.n109 VDD1.n97 11.249
R812 VDD1.n141 VDD1.n140 11.249
R813 VDD1.n61 VDD1.n7 10.4732
R814 VDD1.n37 VDD1.n36 10.4732
R815 VDD1.n113 VDD1.n112 10.4732
R816 VDD1.n137 VDD1.n83 10.4732
R817 VDD1.n60 VDD1.n9 9.69747
R818 VDD1.n40 VDD1.n19 9.69747
R819 VDD1.n116 VDD1.n95 9.69747
R820 VDD1.n136 VDD1.n85 9.69747
R821 VDD1.n76 VDD1.n75 9.45567
R822 VDD1.n153 VDD1.n152 9.45567
R823 VDD1.n52 VDD1.n51 9.3005
R824 VDD1.n11 VDD1.n10 9.3005
R825 VDD1.n58 VDD1.n57 9.3005
R826 VDD1.n60 VDD1.n59 9.3005
R827 VDD1.n7 VDD1.n6 9.3005
R828 VDD1.n66 VDD1.n65 9.3005
R829 VDD1.n68 VDD1.n67 9.3005
R830 VDD1.n4 VDD1.n1 9.3005
R831 VDD1.n75 VDD1.n74 9.3005
R832 VDD1.n50 VDD1.n49 9.3005
R833 VDD1.n15 VDD1.n14 9.3005
R834 VDD1.n44 VDD1.n43 9.3005
R835 VDD1.n42 VDD1.n41 9.3005
R836 VDD1.n19 VDD1.n18 9.3005
R837 VDD1.n36 VDD1.n35 9.3005
R838 VDD1.n34 VDD1.n33 9.3005
R839 VDD1.n23 VDD1.n22 9.3005
R840 VDD1.n28 VDD1.n27 9.3005
R841 VDD1.n152 VDD1.n151 9.3005
R842 VDD1.n91 VDD1.n90 9.3005
R843 VDD1.n120 VDD1.n119 9.3005
R844 VDD1.n118 VDD1.n117 9.3005
R845 VDD1.n95 VDD1.n94 9.3005
R846 VDD1.n112 VDD1.n111 9.3005
R847 VDD1.n110 VDD1.n109 9.3005
R848 VDD1.n99 VDD1.n98 9.3005
R849 VDD1.n104 VDD1.n103 9.3005
R850 VDD1.n126 VDD1.n125 9.3005
R851 VDD1.n128 VDD1.n127 9.3005
R852 VDD1.n87 VDD1.n86 9.3005
R853 VDD1.n134 VDD1.n133 9.3005
R854 VDD1.n136 VDD1.n135 9.3005
R855 VDD1.n83 VDD1.n82 9.3005
R856 VDD1.n142 VDD1.n141 9.3005
R857 VDD1.n144 VDD1.n143 9.3005
R858 VDD1.n145 VDD1.n78 9.3005
R859 VDD1.n57 VDD1.n56 8.92171
R860 VDD1.n41 VDD1.n17 8.92171
R861 VDD1.n117 VDD1.n93 8.92171
R862 VDD1.n133 VDD1.n132 8.92171
R863 VDD1.n53 VDD1.n11 8.14595
R864 VDD1.n45 VDD1.n44 8.14595
R865 VDD1.n121 VDD1.n120 8.14595
R866 VDD1.n129 VDD1.n87 8.14595
R867 VDD1.n52 VDD1.n13 7.3702
R868 VDD1.n48 VDD1.n15 7.3702
R869 VDD1.n124 VDD1.n91 7.3702
R870 VDD1.n128 VDD1.n89 7.3702
R871 VDD1.n49 VDD1.n13 6.59444
R872 VDD1.n49 VDD1.n48 6.59444
R873 VDD1.n125 VDD1.n124 6.59444
R874 VDD1.n125 VDD1.n89 6.59444
R875 VDD1.n53 VDD1.n52 5.81868
R876 VDD1.n45 VDD1.n15 5.81868
R877 VDD1.n121 VDD1.n91 5.81868
R878 VDD1.n129 VDD1.n128 5.81868
R879 VDD1.n56 VDD1.n11 5.04292
R880 VDD1.n44 VDD1.n17 5.04292
R881 VDD1.n120 VDD1.n93 5.04292
R882 VDD1.n132 VDD1.n87 5.04292
R883 VDD1.n57 VDD1.n9 4.26717
R884 VDD1.n41 VDD1.n40 4.26717
R885 VDD1.n117 VDD1.n116 4.26717
R886 VDD1.n133 VDD1.n85 4.26717
R887 VDD1.n27 VDD1.n26 3.70982
R888 VDD1.n103 VDD1.n102 3.70982
R889 VDD1.n61 VDD1.n60 3.49141
R890 VDD1.n37 VDD1.n19 3.49141
R891 VDD1.n113 VDD1.n95 3.49141
R892 VDD1.n137 VDD1.n136 3.49141
R893 VDD1.n64 VDD1.n7 2.71565
R894 VDD1.n36 VDD1.n21 2.71565
R895 VDD1.n112 VDD1.n97 2.71565
R896 VDD1.n140 VDD1.n83 2.71565
R897 VDD1.n65 VDD1.n5 1.93989
R898 VDD1.n33 VDD1.n32 1.93989
R899 VDD1.n109 VDD1.n108 1.93989
R900 VDD1.n141 VDD1.n81 1.93989
R901 VDD1.n76 VDD1.n0 1.16414
R902 VDD1.n69 VDD1.n68 1.16414
R903 VDD1.n29 VDD1.n23 1.16414
R904 VDD1.n105 VDD1.n99 1.16414
R905 VDD1.n146 VDD1.n144 1.16414
R906 VDD1.n153 VDD1.n77 1.16414
R907 VDD1.n74 VDD1.n73 0.388379
R908 VDD1.n4 VDD1.n2 0.388379
R909 VDD1.n28 VDD1.n25 0.388379
R910 VDD1.n104 VDD1.n101 0.388379
R911 VDD1.n145 VDD1.n79 0.388379
R912 VDD1.n151 VDD1.n150 0.388379
R913 VDD1.n75 VDD1.n1 0.155672
R914 VDD1.n67 VDD1.n1 0.155672
R915 VDD1.n67 VDD1.n66 0.155672
R916 VDD1.n66 VDD1.n6 0.155672
R917 VDD1.n59 VDD1.n6 0.155672
R918 VDD1.n59 VDD1.n58 0.155672
R919 VDD1.n58 VDD1.n10 0.155672
R920 VDD1.n51 VDD1.n10 0.155672
R921 VDD1.n51 VDD1.n50 0.155672
R922 VDD1.n50 VDD1.n14 0.155672
R923 VDD1.n43 VDD1.n14 0.155672
R924 VDD1.n43 VDD1.n42 0.155672
R925 VDD1.n42 VDD1.n18 0.155672
R926 VDD1.n35 VDD1.n18 0.155672
R927 VDD1.n35 VDD1.n34 0.155672
R928 VDD1.n34 VDD1.n22 0.155672
R929 VDD1.n27 VDD1.n22 0.155672
R930 VDD1.n103 VDD1.n98 0.155672
R931 VDD1.n110 VDD1.n98 0.155672
R932 VDD1.n111 VDD1.n110 0.155672
R933 VDD1.n111 VDD1.n94 0.155672
R934 VDD1.n118 VDD1.n94 0.155672
R935 VDD1.n119 VDD1.n118 0.155672
R936 VDD1.n119 VDD1.n90 0.155672
R937 VDD1.n126 VDD1.n90 0.155672
R938 VDD1.n127 VDD1.n126 0.155672
R939 VDD1.n127 VDD1.n86 0.155672
R940 VDD1.n134 VDD1.n86 0.155672
R941 VDD1.n135 VDD1.n134 0.155672
R942 VDD1.n135 VDD1.n82 0.155672
R943 VDD1.n142 VDD1.n82 0.155672
R944 VDD1.n143 VDD1.n142 0.155672
R945 VDD1.n143 VDD1.n78 0.155672
R946 VDD1.n152 VDD1.n78 0.155672
R947 B.n337 B.n88 585
R948 B.n336 B.n335 585
R949 B.n334 B.n89 585
R950 B.n333 B.n332 585
R951 B.n331 B.n90 585
R952 B.n330 B.n329 585
R953 B.n328 B.n91 585
R954 B.n327 B.n326 585
R955 B.n325 B.n92 585
R956 B.n324 B.n323 585
R957 B.n322 B.n93 585
R958 B.n321 B.n320 585
R959 B.n319 B.n94 585
R960 B.n318 B.n317 585
R961 B.n316 B.n95 585
R962 B.n315 B.n314 585
R963 B.n313 B.n96 585
R964 B.n312 B.n311 585
R965 B.n310 B.n97 585
R966 B.n309 B.n308 585
R967 B.n307 B.n98 585
R968 B.n306 B.n305 585
R969 B.n304 B.n99 585
R970 B.n303 B.n302 585
R971 B.n301 B.n100 585
R972 B.n300 B.n299 585
R973 B.n298 B.n101 585
R974 B.n297 B.n296 585
R975 B.n295 B.n102 585
R976 B.n294 B.n293 585
R977 B.n292 B.n103 585
R978 B.n291 B.n290 585
R979 B.n289 B.n104 585
R980 B.n288 B.n287 585
R981 B.n286 B.n105 585
R982 B.n285 B.n284 585
R983 B.n283 B.n106 585
R984 B.n282 B.n281 585
R985 B.n280 B.n107 585
R986 B.n279 B.n278 585
R987 B.n277 B.n108 585
R988 B.n276 B.n275 585
R989 B.n274 B.n109 585
R990 B.n273 B.n272 585
R991 B.n271 B.n110 585
R992 B.n270 B.n269 585
R993 B.n268 B.n111 585
R994 B.n266 B.n265 585
R995 B.n264 B.n114 585
R996 B.n263 B.n262 585
R997 B.n261 B.n115 585
R998 B.n260 B.n259 585
R999 B.n258 B.n116 585
R1000 B.n257 B.n256 585
R1001 B.n255 B.n117 585
R1002 B.n254 B.n253 585
R1003 B.n252 B.n118 585
R1004 B.n251 B.n250 585
R1005 B.n246 B.n119 585
R1006 B.n245 B.n244 585
R1007 B.n243 B.n120 585
R1008 B.n242 B.n241 585
R1009 B.n240 B.n121 585
R1010 B.n239 B.n238 585
R1011 B.n237 B.n122 585
R1012 B.n236 B.n235 585
R1013 B.n234 B.n123 585
R1014 B.n233 B.n232 585
R1015 B.n231 B.n124 585
R1016 B.n230 B.n229 585
R1017 B.n228 B.n125 585
R1018 B.n227 B.n226 585
R1019 B.n225 B.n126 585
R1020 B.n224 B.n223 585
R1021 B.n222 B.n127 585
R1022 B.n221 B.n220 585
R1023 B.n219 B.n128 585
R1024 B.n218 B.n217 585
R1025 B.n216 B.n129 585
R1026 B.n215 B.n214 585
R1027 B.n213 B.n130 585
R1028 B.n212 B.n211 585
R1029 B.n210 B.n131 585
R1030 B.n209 B.n208 585
R1031 B.n207 B.n132 585
R1032 B.n206 B.n205 585
R1033 B.n204 B.n133 585
R1034 B.n203 B.n202 585
R1035 B.n201 B.n134 585
R1036 B.n200 B.n199 585
R1037 B.n198 B.n135 585
R1038 B.n197 B.n196 585
R1039 B.n195 B.n136 585
R1040 B.n194 B.n193 585
R1041 B.n192 B.n137 585
R1042 B.n191 B.n190 585
R1043 B.n189 B.n138 585
R1044 B.n188 B.n187 585
R1045 B.n186 B.n139 585
R1046 B.n185 B.n184 585
R1047 B.n183 B.n140 585
R1048 B.n182 B.n181 585
R1049 B.n180 B.n141 585
R1050 B.n179 B.n178 585
R1051 B.n339 B.n338 585
R1052 B.n340 B.n87 585
R1053 B.n342 B.n341 585
R1054 B.n343 B.n86 585
R1055 B.n345 B.n344 585
R1056 B.n346 B.n85 585
R1057 B.n348 B.n347 585
R1058 B.n349 B.n84 585
R1059 B.n351 B.n350 585
R1060 B.n352 B.n83 585
R1061 B.n354 B.n353 585
R1062 B.n355 B.n82 585
R1063 B.n357 B.n356 585
R1064 B.n358 B.n81 585
R1065 B.n360 B.n359 585
R1066 B.n361 B.n80 585
R1067 B.n363 B.n362 585
R1068 B.n364 B.n79 585
R1069 B.n366 B.n365 585
R1070 B.n367 B.n78 585
R1071 B.n369 B.n368 585
R1072 B.n370 B.n77 585
R1073 B.n372 B.n371 585
R1074 B.n373 B.n76 585
R1075 B.n375 B.n374 585
R1076 B.n376 B.n75 585
R1077 B.n378 B.n377 585
R1078 B.n379 B.n74 585
R1079 B.n381 B.n380 585
R1080 B.n382 B.n73 585
R1081 B.n384 B.n383 585
R1082 B.n385 B.n72 585
R1083 B.n387 B.n386 585
R1084 B.n388 B.n71 585
R1085 B.n390 B.n389 585
R1086 B.n391 B.n70 585
R1087 B.n393 B.n392 585
R1088 B.n394 B.n69 585
R1089 B.n396 B.n395 585
R1090 B.n397 B.n68 585
R1091 B.n555 B.n554 585
R1092 B.n553 B.n12 585
R1093 B.n552 B.n551 585
R1094 B.n550 B.n13 585
R1095 B.n549 B.n548 585
R1096 B.n547 B.n14 585
R1097 B.n546 B.n545 585
R1098 B.n544 B.n15 585
R1099 B.n543 B.n542 585
R1100 B.n541 B.n16 585
R1101 B.n540 B.n539 585
R1102 B.n538 B.n17 585
R1103 B.n537 B.n536 585
R1104 B.n535 B.n18 585
R1105 B.n534 B.n533 585
R1106 B.n532 B.n19 585
R1107 B.n531 B.n530 585
R1108 B.n529 B.n20 585
R1109 B.n528 B.n527 585
R1110 B.n526 B.n21 585
R1111 B.n525 B.n524 585
R1112 B.n523 B.n22 585
R1113 B.n522 B.n521 585
R1114 B.n520 B.n23 585
R1115 B.n519 B.n518 585
R1116 B.n517 B.n24 585
R1117 B.n516 B.n515 585
R1118 B.n514 B.n25 585
R1119 B.n513 B.n512 585
R1120 B.n511 B.n26 585
R1121 B.n510 B.n509 585
R1122 B.n508 B.n27 585
R1123 B.n507 B.n506 585
R1124 B.n505 B.n28 585
R1125 B.n504 B.n503 585
R1126 B.n502 B.n29 585
R1127 B.n501 B.n500 585
R1128 B.n499 B.n30 585
R1129 B.n498 B.n497 585
R1130 B.n496 B.n31 585
R1131 B.n495 B.n494 585
R1132 B.n493 B.n32 585
R1133 B.n492 B.n491 585
R1134 B.n490 B.n33 585
R1135 B.n489 B.n488 585
R1136 B.n487 B.n34 585
R1137 B.n486 B.n485 585
R1138 B.n483 B.n35 585
R1139 B.n482 B.n481 585
R1140 B.n480 B.n38 585
R1141 B.n479 B.n478 585
R1142 B.n477 B.n39 585
R1143 B.n476 B.n475 585
R1144 B.n474 B.n40 585
R1145 B.n473 B.n472 585
R1146 B.n471 B.n41 585
R1147 B.n470 B.n469 585
R1148 B.n468 B.n467 585
R1149 B.n466 B.n45 585
R1150 B.n465 B.n464 585
R1151 B.n463 B.n46 585
R1152 B.n462 B.n461 585
R1153 B.n460 B.n47 585
R1154 B.n459 B.n458 585
R1155 B.n457 B.n48 585
R1156 B.n456 B.n455 585
R1157 B.n454 B.n49 585
R1158 B.n453 B.n452 585
R1159 B.n451 B.n50 585
R1160 B.n450 B.n449 585
R1161 B.n448 B.n51 585
R1162 B.n447 B.n446 585
R1163 B.n445 B.n52 585
R1164 B.n444 B.n443 585
R1165 B.n442 B.n53 585
R1166 B.n441 B.n440 585
R1167 B.n439 B.n54 585
R1168 B.n438 B.n437 585
R1169 B.n436 B.n55 585
R1170 B.n435 B.n434 585
R1171 B.n433 B.n56 585
R1172 B.n432 B.n431 585
R1173 B.n430 B.n57 585
R1174 B.n429 B.n428 585
R1175 B.n427 B.n58 585
R1176 B.n426 B.n425 585
R1177 B.n424 B.n59 585
R1178 B.n423 B.n422 585
R1179 B.n421 B.n60 585
R1180 B.n420 B.n419 585
R1181 B.n418 B.n61 585
R1182 B.n417 B.n416 585
R1183 B.n415 B.n62 585
R1184 B.n414 B.n413 585
R1185 B.n412 B.n63 585
R1186 B.n411 B.n410 585
R1187 B.n409 B.n64 585
R1188 B.n408 B.n407 585
R1189 B.n406 B.n65 585
R1190 B.n405 B.n404 585
R1191 B.n403 B.n66 585
R1192 B.n402 B.n401 585
R1193 B.n400 B.n67 585
R1194 B.n399 B.n398 585
R1195 B.n556 B.n11 585
R1196 B.n558 B.n557 585
R1197 B.n559 B.n10 585
R1198 B.n561 B.n560 585
R1199 B.n562 B.n9 585
R1200 B.n564 B.n563 585
R1201 B.n565 B.n8 585
R1202 B.n567 B.n566 585
R1203 B.n568 B.n7 585
R1204 B.n570 B.n569 585
R1205 B.n571 B.n6 585
R1206 B.n573 B.n572 585
R1207 B.n574 B.n5 585
R1208 B.n576 B.n575 585
R1209 B.n577 B.n4 585
R1210 B.n579 B.n578 585
R1211 B.n580 B.n3 585
R1212 B.n582 B.n581 585
R1213 B.n583 B.n0 585
R1214 B.n2 B.n1 585
R1215 B.n152 B.n151 585
R1216 B.n153 B.n150 585
R1217 B.n155 B.n154 585
R1218 B.n156 B.n149 585
R1219 B.n158 B.n157 585
R1220 B.n159 B.n148 585
R1221 B.n161 B.n160 585
R1222 B.n162 B.n147 585
R1223 B.n164 B.n163 585
R1224 B.n165 B.n146 585
R1225 B.n167 B.n166 585
R1226 B.n168 B.n145 585
R1227 B.n170 B.n169 585
R1228 B.n171 B.n144 585
R1229 B.n173 B.n172 585
R1230 B.n174 B.n143 585
R1231 B.n176 B.n175 585
R1232 B.n177 B.n142 585
R1233 B.n178 B.n177 511.721
R1234 B.n338 B.n337 511.721
R1235 B.n398 B.n397 511.721
R1236 B.n554 B.n11 511.721
R1237 B.n112 B.t7 448.151
R1238 B.n42 B.t5 448.151
R1239 B.n247 B.t10 448.151
R1240 B.n36 B.t2 448.151
R1241 B.n247 B.t9 418.964
R1242 B.n112 B.t6 418.964
R1243 B.n42 B.t3 418.964
R1244 B.n36 B.t0 418.964
R1245 B.n113 B.t8 411.108
R1246 B.n43 B.t4 411.108
R1247 B.n248 B.t11 411.108
R1248 B.n37 B.t1 411.108
R1249 B.n585 B.n584 256.663
R1250 B.n584 B.n583 235.042
R1251 B.n584 B.n2 235.042
R1252 B.n178 B.n141 163.367
R1253 B.n182 B.n141 163.367
R1254 B.n183 B.n182 163.367
R1255 B.n184 B.n183 163.367
R1256 B.n184 B.n139 163.367
R1257 B.n188 B.n139 163.367
R1258 B.n189 B.n188 163.367
R1259 B.n190 B.n189 163.367
R1260 B.n190 B.n137 163.367
R1261 B.n194 B.n137 163.367
R1262 B.n195 B.n194 163.367
R1263 B.n196 B.n195 163.367
R1264 B.n196 B.n135 163.367
R1265 B.n200 B.n135 163.367
R1266 B.n201 B.n200 163.367
R1267 B.n202 B.n201 163.367
R1268 B.n202 B.n133 163.367
R1269 B.n206 B.n133 163.367
R1270 B.n207 B.n206 163.367
R1271 B.n208 B.n207 163.367
R1272 B.n208 B.n131 163.367
R1273 B.n212 B.n131 163.367
R1274 B.n213 B.n212 163.367
R1275 B.n214 B.n213 163.367
R1276 B.n214 B.n129 163.367
R1277 B.n218 B.n129 163.367
R1278 B.n219 B.n218 163.367
R1279 B.n220 B.n219 163.367
R1280 B.n220 B.n127 163.367
R1281 B.n224 B.n127 163.367
R1282 B.n225 B.n224 163.367
R1283 B.n226 B.n225 163.367
R1284 B.n226 B.n125 163.367
R1285 B.n230 B.n125 163.367
R1286 B.n231 B.n230 163.367
R1287 B.n232 B.n231 163.367
R1288 B.n232 B.n123 163.367
R1289 B.n236 B.n123 163.367
R1290 B.n237 B.n236 163.367
R1291 B.n238 B.n237 163.367
R1292 B.n238 B.n121 163.367
R1293 B.n242 B.n121 163.367
R1294 B.n243 B.n242 163.367
R1295 B.n244 B.n243 163.367
R1296 B.n244 B.n119 163.367
R1297 B.n251 B.n119 163.367
R1298 B.n252 B.n251 163.367
R1299 B.n253 B.n252 163.367
R1300 B.n253 B.n117 163.367
R1301 B.n257 B.n117 163.367
R1302 B.n258 B.n257 163.367
R1303 B.n259 B.n258 163.367
R1304 B.n259 B.n115 163.367
R1305 B.n263 B.n115 163.367
R1306 B.n264 B.n263 163.367
R1307 B.n265 B.n264 163.367
R1308 B.n265 B.n111 163.367
R1309 B.n270 B.n111 163.367
R1310 B.n271 B.n270 163.367
R1311 B.n272 B.n271 163.367
R1312 B.n272 B.n109 163.367
R1313 B.n276 B.n109 163.367
R1314 B.n277 B.n276 163.367
R1315 B.n278 B.n277 163.367
R1316 B.n278 B.n107 163.367
R1317 B.n282 B.n107 163.367
R1318 B.n283 B.n282 163.367
R1319 B.n284 B.n283 163.367
R1320 B.n284 B.n105 163.367
R1321 B.n288 B.n105 163.367
R1322 B.n289 B.n288 163.367
R1323 B.n290 B.n289 163.367
R1324 B.n290 B.n103 163.367
R1325 B.n294 B.n103 163.367
R1326 B.n295 B.n294 163.367
R1327 B.n296 B.n295 163.367
R1328 B.n296 B.n101 163.367
R1329 B.n300 B.n101 163.367
R1330 B.n301 B.n300 163.367
R1331 B.n302 B.n301 163.367
R1332 B.n302 B.n99 163.367
R1333 B.n306 B.n99 163.367
R1334 B.n307 B.n306 163.367
R1335 B.n308 B.n307 163.367
R1336 B.n308 B.n97 163.367
R1337 B.n312 B.n97 163.367
R1338 B.n313 B.n312 163.367
R1339 B.n314 B.n313 163.367
R1340 B.n314 B.n95 163.367
R1341 B.n318 B.n95 163.367
R1342 B.n319 B.n318 163.367
R1343 B.n320 B.n319 163.367
R1344 B.n320 B.n93 163.367
R1345 B.n324 B.n93 163.367
R1346 B.n325 B.n324 163.367
R1347 B.n326 B.n325 163.367
R1348 B.n326 B.n91 163.367
R1349 B.n330 B.n91 163.367
R1350 B.n331 B.n330 163.367
R1351 B.n332 B.n331 163.367
R1352 B.n332 B.n89 163.367
R1353 B.n336 B.n89 163.367
R1354 B.n337 B.n336 163.367
R1355 B.n397 B.n396 163.367
R1356 B.n396 B.n69 163.367
R1357 B.n392 B.n69 163.367
R1358 B.n392 B.n391 163.367
R1359 B.n391 B.n390 163.367
R1360 B.n390 B.n71 163.367
R1361 B.n386 B.n71 163.367
R1362 B.n386 B.n385 163.367
R1363 B.n385 B.n384 163.367
R1364 B.n384 B.n73 163.367
R1365 B.n380 B.n73 163.367
R1366 B.n380 B.n379 163.367
R1367 B.n379 B.n378 163.367
R1368 B.n378 B.n75 163.367
R1369 B.n374 B.n75 163.367
R1370 B.n374 B.n373 163.367
R1371 B.n373 B.n372 163.367
R1372 B.n372 B.n77 163.367
R1373 B.n368 B.n77 163.367
R1374 B.n368 B.n367 163.367
R1375 B.n367 B.n366 163.367
R1376 B.n366 B.n79 163.367
R1377 B.n362 B.n79 163.367
R1378 B.n362 B.n361 163.367
R1379 B.n361 B.n360 163.367
R1380 B.n360 B.n81 163.367
R1381 B.n356 B.n81 163.367
R1382 B.n356 B.n355 163.367
R1383 B.n355 B.n354 163.367
R1384 B.n354 B.n83 163.367
R1385 B.n350 B.n83 163.367
R1386 B.n350 B.n349 163.367
R1387 B.n349 B.n348 163.367
R1388 B.n348 B.n85 163.367
R1389 B.n344 B.n85 163.367
R1390 B.n344 B.n343 163.367
R1391 B.n343 B.n342 163.367
R1392 B.n342 B.n87 163.367
R1393 B.n338 B.n87 163.367
R1394 B.n554 B.n553 163.367
R1395 B.n553 B.n552 163.367
R1396 B.n552 B.n13 163.367
R1397 B.n548 B.n13 163.367
R1398 B.n548 B.n547 163.367
R1399 B.n547 B.n546 163.367
R1400 B.n546 B.n15 163.367
R1401 B.n542 B.n15 163.367
R1402 B.n542 B.n541 163.367
R1403 B.n541 B.n540 163.367
R1404 B.n540 B.n17 163.367
R1405 B.n536 B.n17 163.367
R1406 B.n536 B.n535 163.367
R1407 B.n535 B.n534 163.367
R1408 B.n534 B.n19 163.367
R1409 B.n530 B.n19 163.367
R1410 B.n530 B.n529 163.367
R1411 B.n529 B.n528 163.367
R1412 B.n528 B.n21 163.367
R1413 B.n524 B.n21 163.367
R1414 B.n524 B.n523 163.367
R1415 B.n523 B.n522 163.367
R1416 B.n522 B.n23 163.367
R1417 B.n518 B.n23 163.367
R1418 B.n518 B.n517 163.367
R1419 B.n517 B.n516 163.367
R1420 B.n516 B.n25 163.367
R1421 B.n512 B.n25 163.367
R1422 B.n512 B.n511 163.367
R1423 B.n511 B.n510 163.367
R1424 B.n510 B.n27 163.367
R1425 B.n506 B.n27 163.367
R1426 B.n506 B.n505 163.367
R1427 B.n505 B.n504 163.367
R1428 B.n504 B.n29 163.367
R1429 B.n500 B.n29 163.367
R1430 B.n500 B.n499 163.367
R1431 B.n499 B.n498 163.367
R1432 B.n498 B.n31 163.367
R1433 B.n494 B.n31 163.367
R1434 B.n494 B.n493 163.367
R1435 B.n493 B.n492 163.367
R1436 B.n492 B.n33 163.367
R1437 B.n488 B.n33 163.367
R1438 B.n488 B.n487 163.367
R1439 B.n487 B.n486 163.367
R1440 B.n486 B.n35 163.367
R1441 B.n481 B.n35 163.367
R1442 B.n481 B.n480 163.367
R1443 B.n480 B.n479 163.367
R1444 B.n479 B.n39 163.367
R1445 B.n475 B.n39 163.367
R1446 B.n475 B.n474 163.367
R1447 B.n474 B.n473 163.367
R1448 B.n473 B.n41 163.367
R1449 B.n469 B.n41 163.367
R1450 B.n469 B.n468 163.367
R1451 B.n468 B.n45 163.367
R1452 B.n464 B.n45 163.367
R1453 B.n464 B.n463 163.367
R1454 B.n463 B.n462 163.367
R1455 B.n462 B.n47 163.367
R1456 B.n458 B.n47 163.367
R1457 B.n458 B.n457 163.367
R1458 B.n457 B.n456 163.367
R1459 B.n456 B.n49 163.367
R1460 B.n452 B.n49 163.367
R1461 B.n452 B.n451 163.367
R1462 B.n451 B.n450 163.367
R1463 B.n450 B.n51 163.367
R1464 B.n446 B.n51 163.367
R1465 B.n446 B.n445 163.367
R1466 B.n445 B.n444 163.367
R1467 B.n444 B.n53 163.367
R1468 B.n440 B.n53 163.367
R1469 B.n440 B.n439 163.367
R1470 B.n439 B.n438 163.367
R1471 B.n438 B.n55 163.367
R1472 B.n434 B.n55 163.367
R1473 B.n434 B.n433 163.367
R1474 B.n433 B.n432 163.367
R1475 B.n432 B.n57 163.367
R1476 B.n428 B.n57 163.367
R1477 B.n428 B.n427 163.367
R1478 B.n427 B.n426 163.367
R1479 B.n426 B.n59 163.367
R1480 B.n422 B.n59 163.367
R1481 B.n422 B.n421 163.367
R1482 B.n421 B.n420 163.367
R1483 B.n420 B.n61 163.367
R1484 B.n416 B.n61 163.367
R1485 B.n416 B.n415 163.367
R1486 B.n415 B.n414 163.367
R1487 B.n414 B.n63 163.367
R1488 B.n410 B.n63 163.367
R1489 B.n410 B.n409 163.367
R1490 B.n409 B.n408 163.367
R1491 B.n408 B.n65 163.367
R1492 B.n404 B.n65 163.367
R1493 B.n404 B.n403 163.367
R1494 B.n403 B.n402 163.367
R1495 B.n402 B.n67 163.367
R1496 B.n398 B.n67 163.367
R1497 B.n558 B.n11 163.367
R1498 B.n559 B.n558 163.367
R1499 B.n560 B.n559 163.367
R1500 B.n560 B.n9 163.367
R1501 B.n564 B.n9 163.367
R1502 B.n565 B.n564 163.367
R1503 B.n566 B.n565 163.367
R1504 B.n566 B.n7 163.367
R1505 B.n570 B.n7 163.367
R1506 B.n571 B.n570 163.367
R1507 B.n572 B.n571 163.367
R1508 B.n572 B.n5 163.367
R1509 B.n576 B.n5 163.367
R1510 B.n577 B.n576 163.367
R1511 B.n578 B.n577 163.367
R1512 B.n578 B.n3 163.367
R1513 B.n582 B.n3 163.367
R1514 B.n583 B.n582 163.367
R1515 B.n152 B.n2 163.367
R1516 B.n153 B.n152 163.367
R1517 B.n154 B.n153 163.367
R1518 B.n154 B.n149 163.367
R1519 B.n158 B.n149 163.367
R1520 B.n159 B.n158 163.367
R1521 B.n160 B.n159 163.367
R1522 B.n160 B.n147 163.367
R1523 B.n164 B.n147 163.367
R1524 B.n165 B.n164 163.367
R1525 B.n166 B.n165 163.367
R1526 B.n166 B.n145 163.367
R1527 B.n170 B.n145 163.367
R1528 B.n171 B.n170 163.367
R1529 B.n172 B.n171 163.367
R1530 B.n172 B.n143 163.367
R1531 B.n176 B.n143 163.367
R1532 B.n177 B.n176 163.367
R1533 B.n249 B.n248 59.5399
R1534 B.n267 B.n113 59.5399
R1535 B.n44 B.n43 59.5399
R1536 B.n484 B.n37 59.5399
R1537 B.n248 B.n247 37.0429
R1538 B.n113 B.n112 37.0429
R1539 B.n43 B.n42 37.0429
R1540 B.n37 B.n36 37.0429
R1541 B.n556 B.n555 33.2493
R1542 B.n399 B.n68 33.2493
R1543 B.n339 B.n88 33.2493
R1544 B.n179 B.n142 33.2493
R1545 B B.n585 18.0485
R1546 B.n557 B.n556 10.6151
R1547 B.n557 B.n10 10.6151
R1548 B.n561 B.n10 10.6151
R1549 B.n562 B.n561 10.6151
R1550 B.n563 B.n562 10.6151
R1551 B.n563 B.n8 10.6151
R1552 B.n567 B.n8 10.6151
R1553 B.n568 B.n567 10.6151
R1554 B.n569 B.n568 10.6151
R1555 B.n569 B.n6 10.6151
R1556 B.n573 B.n6 10.6151
R1557 B.n574 B.n573 10.6151
R1558 B.n575 B.n574 10.6151
R1559 B.n575 B.n4 10.6151
R1560 B.n579 B.n4 10.6151
R1561 B.n580 B.n579 10.6151
R1562 B.n581 B.n580 10.6151
R1563 B.n581 B.n0 10.6151
R1564 B.n555 B.n12 10.6151
R1565 B.n551 B.n12 10.6151
R1566 B.n551 B.n550 10.6151
R1567 B.n550 B.n549 10.6151
R1568 B.n549 B.n14 10.6151
R1569 B.n545 B.n14 10.6151
R1570 B.n545 B.n544 10.6151
R1571 B.n544 B.n543 10.6151
R1572 B.n543 B.n16 10.6151
R1573 B.n539 B.n16 10.6151
R1574 B.n539 B.n538 10.6151
R1575 B.n538 B.n537 10.6151
R1576 B.n537 B.n18 10.6151
R1577 B.n533 B.n18 10.6151
R1578 B.n533 B.n532 10.6151
R1579 B.n532 B.n531 10.6151
R1580 B.n531 B.n20 10.6151
R1581 B.n527 B.n20 10.6151
R1582 B.n527 B.n526 10.6151
R1583 B.n526 B.n525 10.6151
R1584 B.n525 B.n22 10.6151
R1585 B.n521 B.n22 10.6151
R1586 B.n521 B.n520 10.6151
R1587 B.n520 B.n519 10.6151
R1588 B.n519 B.n24 10.6151
R1589 B.n515 B.n24 10.6151
R1590 B.n515 B.n514 10.6151
R1591 B.n514 B.n513 10.6151
R1592 B.n513 B.n26 10.6151
R1593 B.n509 B.n26 10.6151
R1594 B.n509 B.n508 10.6151
R1595 B.n508 B.n507 10.6151
R1596 B.n507 B.n28 10.6151
R1597 B.n503 B.n28 10.6151
R1598 B.n503 B.n502 10.6151
R1599 B.n502 B.n501 10.6151
R1600 B.n501 B.n30 10.6151
R1601 B.n497 B.n30 10.6151
R1602 B.n497 B.n496 10.6151
R1603 B.n496 B.n495 10.6151
R1604 B.n495 B.n32 10.6151
R1605 B.n491 B.n32 10.6151
R1606 B.n491 B.n490 10.6151
R1607 B.n490 B.n489 10.6151
R1608 B.n489 B.n34 10.6151
R1609 B.n485 B.n34 10.6151
R1610 B.n483 B.n482 10.6151
R1611 B.n482 B.n38 10.6151
R1612 B.n478 B.n38 10.6151
R1613 B.n478 B.n477 10.6151
R1614 B.n477 B.n476 10.6151
R1615 B.n476 B.n40 10.6151
R1616 B.n472 B.n40 10.6151
R1617 B.n472 B.n471 10.6151
R1618 B.n471 B.n470 10.6151
R1619 B.n467 B.n466 10.6151
R1620 B.n466 B.n465 10.6151
R1621 B.n465 B.n46 10.6151
R1622 B.n461 B.n46 10.6151
R1623 B.n461 B.n460 10.6151
R1624 B.n460 B.n459 10.6151
R1625 B.n459 B.n48 10.6151
R1626 B.n455 B.n48 10.6151
R1627 B.n455 B.n454 10.6151
R1628 B.n454 B.n453 10.6151
R1629 B.n453 B.n50 10.6151
R1630 B.n449 B.n50 10.6151
R1631 B.n449 B.n448 10.6151
R1632 B.n448 B.n447 10.6151
R1633 B.n447 B.n52 10.6151
R1634 B.n443 B.n52 10.6151
R1635 B.n443 B.n442 10.6151
R1636 B.n442 B.n441 10.6151
R1637 B.n441 B.n54 10.6151
R1638 B.n437 B.n54 10.6151
R1639 B.n437 B.n436 10.6151
R1640 B.n436 B.n435 10.6151
R1641 B.n435 B.n56 10.6151
R1642 B.n431 B.n56 10.6151
R1643 B.n431 B.n430 10.6151
R1644 B.n430 B.n429 10.6151
R1645 B.n429 B.n58 10.6151
R1646 B.n425 B.n58 10.6151
R1647 B.n425 B.n424 10.6151
R1648 B.n424 B.n423 10.6151
R1649 B.n423 B.n60 10.6151
R1650 B.n419 B.n60 10.6151
R1651 B.n419 B.n418 10.6151
R1652 B.n418 B.n417 10.6151
R1653 B.n417 B.n62 10.6151
R1654 B.n413 B.n62 10.6151
R1655 B.n413 B.n412 10.6151
R1656 B.n412 B.n411 10.6151
R1657 B.n411 B.n64 10.6151
R1658 B.n407 B.n64 10.6151
R1659 B.n407 B.n406 10.6151
R1660 B.n406 B.n405 10.6151
R1661 B.n405 B.n66 10.6151
R1662 B.n401 B.n66 10.6151
R1663 B.n401 B.n400 10.6151
R1664 B.n400 B.n399 10.6151
R1665 B.n395 B.n68 10.6151
R1666 B.n395 B.n394 10.6151
R1667 B.n394 B.n393 10.6151
R1668 B.n393 B.n70 10.6151
R1669 B.n389 B.n70 10.6151
R1670 B.n389 B.n388 10.6151
R1671 B.n388 B.n387 10.6151
R1672 B.n387 B.n72 10.6151
R1673 B.n383 B.n72 10.6151
R1674 B.n383 B.n382 10.6151
R1675 B.n382 B.n381 10.6151
R1676 B.n381 B.n74 10.6151
R1677 B.n377 B.n74 10.6151
R1678 B.n377 B.n376 10.6151
R1679 B.n376 B.n375 10.6151
R1680 B.n375 B.n76 10.6151
R1681 B.n371 B.n76 10.6151
R1682 B.n371 B.n370 10.6151
R1683 B.n370 B.n369 10.6151
R1684 B.n369 B.n78 10.6151
R1685 B.n365 B.n78 10.6151
R1686 B.n365 B.n364 10.6151
R1687 B.n364 B.n363 10.6151
R1688 B.n363 B.n80 10.6151
R1689 B.n359 B.n80 10.6151
R1690 B.n359 B.n358 10.6151
R1691 B.n358 B.n357 10.6151
R1692 B.n357 B.n82 10.6151
R1693 B.n353 B.n82 10.6151
R1694 B.n353 B.n352 10.6151
R1695 B.n352 B.n351 10.6151
R1696 B.n351 B.n84 10.6151
R1697 B.n347 B.n84 10.6151
R1698 B.n347 B.n346 10.6151
R1699 B.n346 B.n345 10.6151
R1700 B.n345 B.n86 10.6151
R1701 B.n341 B.n86 10.6151
R1702 B.n341 B.n340 10.6151
R1703 B.n340 B.n339 10.6151
R1704 B.n151 B.n1 10.6151
R1705 B.n151 B.n150 10.6151
R1706 B.n155 B.n150 10.6151
R1707 B.n156 B.n155 10.6151
R1708 B.n157 B.n156 10.6151
R1709 B.n157 B.n148 10.6151
R1710 B.n161 B.n148 10.6151
R1711 B.n162 B.n161 10.6151
R1712 B.n163 B.n162 10.6151
R1713 B.n163 B.n146 10.6151
R1714 B.n167 B.n146 10.6151
R1715 B.n168 B.n167 10.6151
R1716 B.n169 B.n168 10.6151
R1717 B.n169 B.n144 10.6151
R1718 B.n173 B.n144 10.6151
R1719 B.n174 B.n173 10.6151
R1720 B.n175 B.n174 10.6151
R1721 B.n175 B.n142 10.6151
R1722 B.n180 B.n179 10.6151
R1723 B.n181 B.n180 10.6151
R1724 B.n181 B.n140 10.6151
R1725 B.n185 B.n140 10.6151
R1726 B.n186 B.n185 10.6151
R1727 B.n187 B.n186 10.6151
R1728 B.n187 B.n138 10.6151
R1729 B.n191 B.n138 10.6151
R1730 B.n192 B.n191 10.6151
R1731 B.n193 B.n192 10.6151
R1732 B.n193 B.n136 10.6151
R1733 B.n197 B.n136 10.6151
R1734 B.n198 B.n197 10.6151
R1735 B.n199 B.n198 10.6151
R1736 B.n199 B.n134 10.6151
R1737 B.n203 B.n134 10.6151
R1738 B.n204 B.n203 10.6151
R1739 B.n205 B.n204 10.6151
R1740 B.n205 B.n132 10.6151
R1741 B.n209 B.n132 10.6151
R1742 B.n210 B.n209 10.6151
R1743 B.n211 B.n210 10.6151
R1744 B.n211 B.n130 10.6151
R1745 B.n215 B.n130 10.6151
R1746 B.n216 B.n215 10.6151
R1747 B.n217 B.n216 10.6151
R1748 B.n217 B.n128 10.6151
R1749 B.n221 B.n128 10.6151
R1750 B.n222 B.n221 10.6151
R1751 B.n223 B.n222 10.6151
R1752 B.n223 B.n126 10.6151
R1753 B.n227 B.n126 10.6151
R1754 B.n228 B.n227 10.6151
R1755 B.n229 B.n228 10.6151
R1756 B.n229 B.n124 10.6151
R1757 B.n233 B.n124 10.6151
R1758 B.n234 B.n233 10.6151
R1759 B.n235 B.n234 10.6151
R1760 B.n235 B.n122 10.6151
R1761 B.n239 B.n122 10.6151
R1762 B.n240 B.n239 10.6151
R1763 B.n241 B.n240 10.6151
R1764 B.n241 B.n120 10.6151
R1765 B.n245 B.n120 10.6151
R1766 B.n246 B.n245 10.6151
R1767 B.n250 B.n246 10.6151
R1768 B.n254 B.n118 10.6151
R1769 B.n255 B.n254 10.6151
R1770 B.n256 B.n255 10.6151
R1771 B.n256 B.n116 10.6151
R1772 B.n260 B.n116 10.6151
R1773 B.n261 B.n260 10.6151
R1774 B.n262 B.n261 10.6151
R1775 B.n262 B.n114 10.6151
R1776 B.n266 B.n114 10.6151
R1777 B.n269 B.n268 10.6151
R1778 B.n269 B.n110 10.6151
R1779 B.n273 B.n110 10.6151
R1780 B.n274 B.n273 10.6151
R1781 B.n275 B.n274 10.6151
R1782 B.n275 B.n108 10.6151
R1783 B.n279 B.n108 10.6151
R1784 B.n280 B.n279 10.6151
R1785 B.n281 B.n280 10.6151
R1786 B.n281 B.n106 10.6151
R1787 B.n285 B.n106 10.6151
R1788 B.n286 B.n285 10.6151
R1789 B.n287 B.n286 10.6151
R1790 B.n287 B.n104 10.6151
R1791 B.n291 B.n104 10.6151
R1792 B.n292 B.n291 10.6151
R1793 B.n293 B.n292 10.6151
R1794 B.n293 B.n102 10.6151
R1795 B.n297 B.n102 10.6151
R1796 B.n298 B.n297 10.6151
R1797 B.n299 B.n298 10.6151
R1798 B.n299 B.n100 10.6151
R1799 B.n303 B.n100 10.6151
R1800 B.n304 B.n303 10.6151
R1801 B.n305 B.n304 10.6151
R1802 B.n305 B.n98 10.6151
R1803 B.n309 B.n98 10.6151
R1804 B.n310 B.n309 10.6151
R1805 B.n311 B.n310 10.6151
R1806 B.n311 B.n96 10.6151
R1807 B.n315 B.n96 10.6151
R1808 B.n316 B.n315 10.6151
R1809 B.n317 B.n316 10.6151
R1810 B.n317 B.n94 10.6151
R1811 B.n321 B.n94 10.6151
R1812 B.n322 B.n321 10.6151
R1813 B.n323 B.n322 10.6151
R1814 B.n323 B.n92 10.6151
R1815 B.n327 B.n92 10.6151
R1816 B.n328 B.n327 10.6151
R1817 B.n329 B.n328 10.6151
R1818 B.n329 B.n90 10.6151
R1819 B.n333 B.n90 10.6151
R1820 B.n334 B.n333 10.6151
R1821 B.n335 B.n334 10.6151
R1822 B.n335 B.n88 10.6151
R1823 B.n485 B.n484 9.36635
R1824 B.n467 B.n44 9.36635
R1825 B.n250 B.n249 9.36635
R1826 B.n268 B.n267 9.36635
R1827 B.n585 B.n0 8.11757
R1828 B.n585 B.n1 8.11757
R1829 B.n484 B.n483 1.24928
R1830 B.n470 B.n44 1.24928
R1831 B.n249 B.n118 1.24928
R1832 B.n267 B.n266 1.24928
C0 w_n1734_n3764# VDD2 1.8221f
C1 VTAIL B 3.60156f
C2 VN VTAIL 2.41965f
C3 VP VDD2 0.290218f
C4 VN B 0.897844f
C5 VTAIL VDD2 5.67128f
C6 B VDD2 1.73324f
C7 VDD1 w_n1734_n3764# 1.80844f
C8 VN VDD2 2.90643f
C9 VDD1 VP 3.0456f
C10 VTAIL VDD1 5.62973f
C11 w_n1734_n3764# VP 2.55389f
C12 VDD1 B 1.71217f
C13 VN VDD1 0.14732f
C14 VTAIL w_n1734_n3764# 3.0852f
C15 w_n1734_n3764# B 8.261451f
C16 VTAIL VP 2.43411f
C17 VDD1 VDD2 0.555516f
C18 VN w_n1734_n3764# 2.33521f
C19 VP B 1.25327f
C20 VN VP 5.34241f
C21 VDD2 VSUBS 0.873244f
C22 VDD1 VSUBS 3.575196f
C23 VTAIL VSUBS 0.964877f
C24 VN VSUBS 7.90498f
C25 VP VSUBS 1.447657f
C26 B VSUBS 3.306309f
C27 w_n1734_n3764# VSUBS 80.1316f
C28 B.n0 VSUBS 0.005666f
C29 B.n1 VSUBS 0.005666f
C30 B.n2 VSUBS 0.00838f
C31 B.n3 VSUBS 0.006421f
C32 B.n4 VSUBS 0.006421f
C33 B.n5 VSUBS 0.006421f
C34 B.n6 VSUBS 0.006421f
C35 B.n7 VSUBS 0.006421f
C36 B.n8 VSUBS 0.006421f
C37 B.n9 VSUBS 0.006421f
C38 B.n10 VSUBS 0.006421f
C39 B.n11 VSUBS 0.015085f
C40 B.n12 VSUBS 0.006421f
C41 B.n13 VSUBS 0.006421f
C42 B.n14 VSUBS 0.006421f
C43 B.n15 VSUBS 0.006421f
C44 B.n16 VSUBS 0.006421f
C45 B.n17 VSUBS 0.006421f
C46 B.n18 VSUBS 0.006421f
C47 B.n19 VSUBS 0.006421f
C48 B.n20 VSUBS 0.006421f
C49 B.n21 VSUBS 0.006421f
C50 B.n22 VSUBS 0.006421f
C51 B.n23 VSUBS 0.006421f
C52 B.n24 VSUBS 0.006421f
C53 B.n25 VSUBS 0.006421f
C54 B.n26 VSUBS 0.006421f
C55 B.n27 VSUBS 0.006421f
C56 B.n28 VSUBS 0.006421f
C57 B.n29 VSUBS 0.006421f
C58 B.n30 VSUBS 0.006421f
C59 B.n31 VSUBS 0.006421f
C60 B.n32 VSUBS 0.006421f
C61 B.n33 VSUBS 0.006421f
C62 B.n34 VSUBS 0.006421f
C63 B.n35 VSUBS 0.006421f
C64 B.t1 VSUBS 0.234582f
C65 B.t2 VSUBS 0.254639f
C66 B.t0 VSUBS 0.880437f
C67 B.n36 VSUBS 0.37918f
C68 B.n37 VSUBS 0.25181f
C69 B.n38 VSUBS 0.006421f
C70 B.n39 VSUBS 0.006421f
C71 B.n40 VSUBS 0.006421f
C72 B.n41 VSUBS 0.006421f
C73 B.t4 VSUBS 0.234585f
C74 B.t5 VSUBS 0.254641f
C75 B.t3 VSUBS 0.880437f
C76 B.n42 VSUBS 0.379178f
C77 B.n43 VSUBS 0.251807f
C78 B.n44 VSUBS 0.014878f
C79 B.n45 VSUBS 0.006421f
C80 B.n46 VSUBS 0.006421f
C81 B.n47 VSUBS 0.006421f
C82 B.n48 VSUBS 0.006421f
C83 B.n49 VSUBS 0.006421f
C84 B.n50 VSUBS 0.006421f
C85 B.n51 VSUBS 0.006421f
C86 B.n52 VSUBS 0.006421f
C87 B.n53 VSUBS 0.006421f
C88 B.n54 VSUBS 0.006421f
C89 B.n55 VSUBS 0.006421f
C90 B.n56 VSUBS 0.006421f
C91 B.n57 VSUBS 0.006421f
C92 B.n58 VSUBS 0.006421f
C93 B.n59 VSUBS 0.006421f
C94 B.n60 VSUBS 0.006421f
C95 B.n61 VSUBS 0.006421f
C96 B.n62 VSUBS 0.006421f
C97 B.n63 VSUBS 0.006421f
C98 B.n64 VSUBS 0.006421f
C99 B.n65 VSUBS 0.006421f
C100 B.n66 VSUBS 0.006421f
C101 B.n67 VSUBS 0.006421f
C102 B.n68 VSUBS 0.015085f
C103 B.n69 VSUBS 0.006421f
C104 B.n70 VSUBS 0.006421f
C105 B.n71 VSUBS 0.006421f
C106 B.n72 VSUBS 0.006421f
C107 B.n73 VSUBS 0.006421f
C108 B.n74 VSUBS 0.006421f
C109 B.n75 VSUBS 0.006421f
C110 B.n76 VSUBS 0.006421f
C111 B.n77 VSUBS 0.006421f
C112 B.n78 VSUBS 0.006421f
C113 B.n79 VSUBS 0.006421f
C114 B.n80 VSUBS 0.006421f
C115 B.n81 VSUBS 0.006421f
C116 B.n82 VSUBS 0.006421f
C117 B.n83 VSUBS 0.006421f
C118 B.n84 VSUBS 0.006421f
C119 B.n85 VSUBS 0.006421f
C120 B.n86 VSUBS 0.006421f
C121 B.n87 VSUBS 0.006421f
C122 B.n88 VSUBS 0.014576f
C123 B.n89 VSUBS 0.006421f
C124 B.n90 VSUBS 0.006421f
C125 B.n91 VSUBS 0.006421f
C126 B.n92 VSUBS 0.006421f
C127 B.n93 VSUBS 0.006421f
C128 B.n94 VSUBS 0.006421f
C129 B.n95 VSUBS 0.006421f
C130 B.n96 VSUBS 0.006421f
C131 B.n97 VSUBS 0.006421f
C132 B.n98 VSUBS 0.006421f
C133 B.n99 VSUBS 0.006421f
C134 B.n100 VSUBS 0.006421f
C135 B.n101 VSUBS 0.006421f
C136 B.n102 VSUBS 0.006421f
C137 B.n103 VSUBS 0.006421f
C138 B.n104 VSUBS 0.006421f
C139 B.n105 VSUBS 0.006421f
C140 B.n106 VSUBS 0.006421f
C141 B.n107 VSUBS 0.006421f
C142 B.n108 VSUBS 0.006421f
C143 B.n109 VSUBS 0.006421f
C144 B.n110 VSUBS 0.006421f
C145 B.n111 VSUBS 0.006421f
C146 B.t8 VSUBS 0.234585f
C147 B.t7 VSUBS 0.254641f
C148 B.t6 VSUBS 0.880437f
C149 B.n112 VSUBS 0.379178f
C150 B.n113 VSUBS 0.251807f
C151 B.n114 VSUBS 0.006421f
C152 B.n115 VSUBS 0.006421f
C153 B.n116 VSUBS 0.006421f
C154 B.n117 VSUBS 0.006421f
C155 B.n118 VSUBS 0.003588f
C156 B.n119 VSUBS 0.006421f
C157 B.n120 VSUBS 0.006421f
C158 B.n121 VSUBS 0.006421f
C159 B.n122 VSUBS 0.006421f
C160 B.n123 VSUBS 0.006421f
C161 B.n124 VSUBS 0.006421f
C162 B.n125 VSUBS 0.006421f
C163 B.n126 VSUBS 0.006421f
C164 B.n127 VSUBS 0.006421f
C165 B.n128 VSUBS 0.006421f
C166 B.n129 VSUBS 0.006421f
C167 B.n130 VSUBS 0.006421f
C168 B.n131 VSUBS 0.006421f
C169 B.n132 VSUBS 0.006421f
C170 B.n133 VSUBS 0.006421f
C171 B.n134 VSUBS 0.006421f
C172 B.n135 VSUBS 0.006421f
C173 B.n136 VSUBS 0.006421f
C174 B.n137 VSUBS 0.006421f
C175 B.n138 VSUBS 0.006421f
C176 B.n139 VSUBS 0.006421f
C177 B.n140 VSUBS 0.006421f
C178 B.n141 VSUBS 0.006421f
C179 B.n142 VSUBS 0.015085f
C180 B.n143 VSUBS 0.006421f
C181 B.n144 VSUBS 0.006421f
C182 B.n145 VSUBS 0.006421f
C183 B.n146 VSUBS 0.006421f
C184 B.n147 VSUBS 0.006421f
C185 B.n148 VSUBS 0.006421f
C186 B.n149 VSUBS 0.006421f
C187 B.n150 VSUBS 0.006421f
C188 B.n151 VSUBS 0.006421f
C189 B.n152 VSUBS 0.006421f
C190 B.n153 VSUBS 0.006421f
C191 B.n154 VSUBS 0.006421f
C192 B.n155 VSUBS 0.006421f
C193 B.n156 VSUBS 0.006421f
C194 B.n157 VSUBS 0.006421f
C195 B.n158 VSUBS 0.006421f
C196 B.n159 VSUBS 0.006421f
C197 B.n160 VSUBS 0.006421f
C198 B.n161 VSUBS 0.006421f
C199 B.n162 VSUBS 0.006421f
C200 B.n163 VSUBS 0.006421f
C201 B.n164 VSUBS 0.006421f
C202 B.n165 VSUBS 0.006421f
C203 B.n166 VSUBS 0.006421f
C204 B.n167 VSUBS 0.006421f
C205 B.n168 VSUBS 0.006421f
C206 B.n169 VSUBS 0.006421f
C207 B.n170 VSUBS 0.006421f
C208 B.n171 VSUBS 0.006421f
C209 B.n172 VSUBS 0.006421f
C210 B.n173 VSUBS 0.006421f
C211 B.n174 VSUBS 0.006421f
C212 B.n175 VSUBS 0.006421f
C213 B.n176 VSUBS 0.006421f
C214 B.n177 VSUBS 0.015085f
C215 B.n178 VSUBS 0.015322f
C216 B.n179 VSUBS 0.015322f
C217 B.n180 VSUBS 0.006421f
C218 B.n181 VSUBS 0.006421f
C219 B.n182 VSUBS 0.006421f
C220 B.n183 VSUBS 0.006421f
C221 B.n184 VSUBS 0.006421f
C222 B.n185 VSUBS 0.006421f
C223 B.n186 VSUBS 0.006421f
C224 B.n187 VSUBS 0.006421f
C225 B.n188 VSUBS 0.006421f
C226 B.n189 VSUBS 0.006421f
C227 B.n190 VSUBS 0.006421f
C228 B.n191 VSUBS 0.006421f
C229 B.n192 VSUBS 0.006421f
C230 B.n193 VSUBS 0.006421f
C231 B.n194 VSUBS 0.006421f
C232 B.n195 VSUBS 0.006421f
C233 B.n196 VSUBS 0.006421f
C234 B.n197 VSUBS 0.006421f
C235 B.n198 VSUBS 0.006421f
C236 B.n199 VSUBS 0.006421f
C237 B.n200 VSUBS 0.006421f
C238 B.n201 VSUBS 0.006421f
C239 B.n202 VSUBS 0.006421f
C240 B.n203 VSUBS 0.006421f
C241 B.n204 VSUBS 0.006421f
C242 B.n205 VSUBS 0.006421f
C243 B.n206 VSUBS 0.006421f
C244 B.n207 VSUBS 0.006421f
C245 B.n208 VSUBS 0.006421f
C246 B.n209 VSUBS 0.006421f
C247 B.n210 VSUBS 0.006421f
C248 B.n211 VSUBS 0.006421f
C249 B.n212 VSUBS 0.006421f
C250 B.n213 VSUBS 0.006421f
C251 B.n214 VSUBS 0.006421f
C252 B.n215 VSUBS 0.006421f
C253 B.n216 VSUBS 0.006421f
C254 B.n217 VSUBS 0.006421f
C255 B.n218 VSUBS 0.006421f
C256 B.n219 VSUBS 0.006421f
C257 B.n220 VSUBS 0.006421f
C258 B.n221 VSUBS 0.006421f
C259 B.n222 VSUBS 0.006421f
C260 B.n223 VSUBS 0.006421f
C261 B.n224 VSUBS 0.006421f
C262 B.n225 VSUBS 0.006421f
C263 B.n226 VSUBS 0.006421f
C264 B.n227 VSUBS 0.006421f
C265 B.n228 VSUBS 0.006421f
C266 B.n229 VSUBS 0.006421f
C267 B.n230 VSUBS 0.006421f
C268 B.n231 VSUBS 0.006421f
C269 B.n232 VSUBS 0.006421f
C270 B.n233 VSUBS 0.006421f
C271 B.n234 VSUBS 0.006421f
C272 B.n235 VSUBS 0.006421f
C273 B.n236 VSUBS 0.006421f
C274 B.n237 VSUBS 0.006421f
C275 B.n238 VSUBS 0.006421f
C276 B.n239 VSUBS 0.006421f
C277 B.n240 VSUBS 0.006421f
C278 B.n241 VSUBS 0.006421f
C279 B.n242 VSUBS 0.006421f
C280 B.n243 VSUBS 0.006421f
C281 B.n244 VSUBS 0.006421f
C282 B.n245 VSUBS 0.006421f
C283 B.n246 VSUBS 0.006421f
C284 B.t11 VSUBS 0.234582f
C285 B.t10 VSUBS 0.254639f
C286 B.t9 VSUBS 0.880437f
C287 B.n247 VSUBS 0.37918f
C288 B.n248 VSUBS 0.25181f
C289 B.n249 VSUBS 0.014878f
C290 B.n250 VSUBS 0.006044f
C291 B.n251 VSUBS 0.006421f
C292 B.n252 VSUBS 0.006421f
C293 B.n253 VSUBS 0.006421f
C294 B.n254 VSUBS 0.006421f
C295 B.n255 VSUBS 0.006421f
C296 B.n256 VSUBS 0.006421f
C297 B.n257 VSUBS 0.006421f
C298 B.n258 VSUBS 0.006421f
C299 B.n259 VSUBS 0.006421f
C300 B.n260 VSUBS 0.006421f
C301 B.n261 VSUBS 0.006421f
C302 B.n262 VSUBS 0.006421f
C303 B.n263 VSUBS 0.006421f
C304 B.n264 VSUBS 0.006421f
C305 B.n265 VSUBS 0.006421f
C306 B.n266 VSUBS 0.003588f
C307 B.n267 VSUBS 0.014878f
C308 B.n268 VSUBS 0.006044f
C309 B.n269 VSUBS 0.006421f
C310 B.n270 VSUBS 0.006421f
C311 B.n271 VSUBS 0.006421f
C312 B.n272 VSUBS 0.006421f
C313 B.n273 VSUBS 0.006421f
C314 B.n274 VSUBS 0.006421f
C315 B.n275 VSUBS 0.006421f
C316 B.n276 VSUBS 0.006421f
C317 B.n277 VSUBS 0.006421f
C318 B.n278 VSUBS 0.006421f
C319 B.n279 VSUBS 0.006421f
C320 B.n280 VSUBS 0.006421f
C321 B.n281 VSUBS 0.006421f
C322 B.n282 VSUBS 0.006421f
C323 B.n283 VSUBS 0.006421f
C324 B.n284 VSUBS 0.006421f
C325 B.n285 VSUBS 0.006421f
C326 B.n286 VSUBS 0.006421f
C327 B.n287 VSUBS 0.006421f
C328 B.n288 VSUBS 0.006421f
C329 B.n289 VSUBS 0.006421f
C330 B.n290 VSUBS 0.006421f
C331 B.n291 VSUBS 0.006421f
C332 B.n292 VSUBS 0.006421f
C333 B.n293 VSUBS 0.006421f
C334 B.n294 VSUBS 0.006421f
C335 B.n295 VSUBS 0.006421f
C336 B.n296 VSUBS 0.006421f
C337 B.n297 VSUBS 0.006421f
C338 B.n298 VSUBS 0.006421f
C339 B.n299 VSUBS 0.006421f
C340 B.n300 VSUBS 0.006421f
C341 B.n301 VSUBS 0.006421f
C342 B.n302 VSUBS 0.006421f
C343 B.n303 VSUBS 0.006421f
C344 B.n304 VSUBS 0.006421f
C345 B.n305 VSUBS 0.006421f
C346 B.n306 VSUBS 0.006421f
C347 B.n307 VSUBS 0.006421f
C348 B.n308 VSUBS 0.006421f
C349 B.n309 VSUBS 0.006421f
C350 B.n310 VSUBS 0.006421f
C351 B.n311 VSUBS 0.006421f
C352 B.n312 VSUBS 0.006421f
C353 B.n313 VSUBS 0.006421f
C354 B.n314 VSUBS 0.006421f
C355 B.n315 VSUBS 0.006421f
C356 B.n316 VSUBS 0.006421f
C357 B.n317 VSUBS 0.006421f
C358 B.n318 VSUBS 0.006421f
C359 B.n319 VSUBS 0.006421f
C360 B.n320 VSUBS 0.006421f
C361 B.n321 VSUBS 0.006421f
C362 B.n322 VSUBS 0.006421f
C363 B.n323 VSUBS 0.006421f
C364 B.n324 VSUBS 0.006421f
C365 B.n325 VSUBS 0.006421f
C366 B.n326 VSUBS 0.006421f
C367 B.n327 VSUBS 0.006421f
C368 B.n328 VSUBS 0.006421f
C369 B.n329 VSUBS 0.006421f
C370 B.n330 VSUBS 0.006421f
C371 B.n331 VSUBS 0.006421f
C372 B.n332 VSUBS 0.006421f
C373 B.n333 VSUBS 0.006421f
C374 B.n334 VSUBS 0.006421f
C375 B.n335 VSUBS 0.006421f
C376 B.n336 VSUBS 0.006421f
C377 B.n337 VSUBS 0.015322f
C378 B.n338 VSUBS 0.015085f
C379 B.n339 VSUBS 0.015831f
C380 B.n340 VSUBS 0.006421f
C381 B.n341 VSUBS 0.006421f
C382 B.n342 VSUBS 0.006421f
C383 B.n343 VSUBS 0.006421f
C384 B.n344 VSUBS 0.006421f
C385 B.n345 VSUBS 0.006421f
C386 B.n346 VSUBS 0.006421f
C387 B.n347 VSUBS 0.006421f
C388 B.n348 VSUBS 0.006421f
C389 B.n349 VSUBS 0.006421f
C390 B.n350 VSUBS 0.006421f
C391 B.n351 VSUBS 0.006421f
C392 B.n352 VSUBS 0.006421f
C393 B.n353 VSUBS 0.006421f
C394 B.n354 VSUBS 0.006421f
C395 B.n355 VSUBS 0.006421f
C396 B.n356 VSUBS 0.006421f
C397 B.n357 VSUBS 0.006421f
C398 B.n358 VSUBS 0.006421f
C399 B.n359 VSUBS 0.006421f
C400 B.n360 VSUBS 0.006421f
C401 B.n361 VSUBS 0.006421f
C402 B.n362 VSUBS 0.006421f
C403 B.n363 VSUBS 0.006421f
C404 B.n364 VSUBS 0.006421f
C405 B.n365 VSUBS 0.006421f
C406 B.n366 VSUBS 0.006421f
C407 B.n367 VSUBS 0.006421f
C408 B.n368 VSUBS 0.006421f
C409 B.n369 VSUBS 0.006421f
C410 B.n370 VSUBS 0.006421f
C411 B.n371 VSUBS 0.006421f
C412 B.n372 VSUBS 0.006421f
C413 B.n373 VSUBS 0.006421f
C414 B.n374 VSUBS 0.006421f
C415 B.n375 VSUBS 0.006421f
C416 B.n376 VSUBS 0.006421f
C417 B.n377 VSUBS 0.006421f
C418 B.n378 VSUBS 0.006421f
C419 B.n379 VSUBS 0.006421f
C420 B.n380 VSUBS 0.006421f
C421 B.n381 VSUBS 0.006421f
C422 B.n382 VSUBS 0.006421f
C423 B.n383 VSUBS 0.006421f
C424 B.n384 VSUBS 0.006421f
C425 B.n385 VSUBS 0.006421f
C426 B.n386 VSUBS 0.006421f
C427 B.n387 VSUBS 0.006421f
C428 B.n388 VSUBS 0.006421f
C429 B.n389 VSUBS 0.006421f
C430 B.n390 VSUBS 0.006421f
C431 B.n391 VSUBS 0.006421f
C432 B.n392 VSUBS 0.006421f
C433 B.n393 VSUBS 0.006421f
C434 B.n394 VSUBS 0.006421f
C435 B.n395 VSUBS 0.006421f
C436 B.n396 VSUBS 0.006421f
C437 B.n397 VSUBS 0.015085f
C438 B.n398 VSUBS 0.015322f
C439 B.n399 VSUBS 0.015322f
C440 B.n400 VSUBS 0.006421f
C441 B.n401 VSUBS 0.006421f
C442 B.n402 VSUBS 0.006421f
C443 B.n403 VSUBS 0.006421f
C444 B.n404 VSUBS 0.006421f
C445 B.n405 VSUBS 0.006421f
C446 B.n406 VSUBS 0.006421f
C447 B.n407 VSUBS 0.006421f
C448 B.n408 VSUBS 0.006421f
C449 B.n409 VSUBS 0.006421f
C450 B.n410 VSUBS 0.006421f
C451 B.n411 VSUBS 0.006421f
C452 B.n412 VSUBS 0.006421f
C453 B.n413 VSUBS 0.006421f
C454 B.n414 VSUBS 0.006421f
C455 B.n415 VSUBS 0.006421f
C456 B.n416 VSUBS 0.006421f
C457 B.n417 VSUBS 0.006421f
C458 B.n418 VSUBS 0.006421f
C459 B.n419 VSUBS 0.006421f
C460 B.n420 VSUBS 0.006421f
C461 B.n421 VSUBS 0.006421f
C462 B.n422 VSUBS 0.006421f
C463 B.n423 VSUBS 0.006421f
C464 B.n424 VSUBS 0.006421f
C465 B.n425 VSUBS 0.006421f
C466 B.n426 VSUBS 0.006421f
C467 B.n427 VSUBS 0.006421f
C468 B.n428 VSUBS 0.006421f
C469 B.n429 VSUBS 0.006421f
C470 B.n430 VSUBS 0.006421f
C471 B.n431 VSUBS 0.006421f
C472 B.n432 VSUBS 0.006421f
C473 B.n433 VSUBS 0.006421f
C474 B.n434 VSUBS 0.006421f
C475 B.n435 VSUBS 0.006421f
C476 B.n436 VSUBS 0.006421f
C477 B.n437 VSUBS 0.006421f
C478 B.n438 VSUBS 0.006421f
C479 B.n439 VSUBS 0.006421f
C480 B.n440 VSUBS 0.006421f
C481 B.n441 VSUBS 0.006421f
C482 B.n442 VSUBS 0.006421f
C483 B.n443 VSUBS 0.006421f
C484 B.n444 VSUBS 0.006421f
C485 B.n445 VSUBS 0.006421f
C486 B.n446 VSUBS 0.006421f
C487 B.n447 VSUBS 0.006421f
C488 B.n448 VSUBS 0.006421f
C489 B.n449 VSUBS 0.006421f
C490 B.n450 VSUBS 0.006421f
C491 B.n451 VSUBS 0.006421f
C492 B.n452 VSUBS 0.006421f
C493 B.n453 VSUBS 0.006421f
C494 B.n454 VSUBS 0.006421f
C495 B.n455 VSUBS 0.006421f
C496 B.n456 VSUBS 0.006421f
C497 B.n457 VSUBS 0.006421f
C498 B.n458 VSUBS 0.006421f
C499 B.n459 VSUBS 0.006421f
C500 B.n460 VSUBS 0.006421f
C501 B.n461 VSUBS 0.006421f
C502 B.n462 VSUBS 0.006421f
C503 B.n463 VSUBS 0.006421f
C504 B.n464 VSUBS 0.006421f
C505 B.n465 VSUBS 0.006421f
C506 B.n466 VSUBS 0.006421f
C507 B.n467 VSUBS 0.006044f
C508 B.n468 VSUBS 0.006421f
C509 B.n469 VSUBS 0.006421f
C510 B.n470 VSUBS 0.003588f
C511 B.n471 VSUBS 0.006421f
C512 B.n472 VSUBS 0.006421f
C513 B.n473 VSUBS 0.006421f
C514 B.n474 VSUBS 0.006421f
C515 B.n475 VSUBS 0.006421f
C516 B.n476 VSUBS 0.006421f
C517 B.n477 VSUBS 0.006421f
C518 B.n478 VSUBS 0.006421f
C519 B.n479 VSUBS 0.006421f
C520 B.n480 VSUBS 0.006421f
C521 B.n481 VSUBS 0.006421f
C522 B.n482 VSUBS 0.006421f
C523 B.n483 VSUBS 0.003588f
C524 B.n484 VSUBS 0.014878f
C525 B.n485 VSUBS 0.006044f
C526 B.n486 VSUBS 0.006421f
C527 B.n487 VSUBS 0.006421f
C528 B.n488 VSUBS 0.006421f
C529 B.n489 VSUBS 0.006421f
C530 B.n490 VSUBS 0.006421f
C531 B.n491 VSUBS 0.006421f
C532 B.n492 VSUBS 0.006421f
C533 B.n493 VSUBS 0.006421f
C534 B.n494 VSUBS 0.006421f
C535 B.n495 VSUBS 0.006421f
C536 B.n496 VSUBS 0.006421f
C537 B.n497 VSUBS 0.006421f
C538 B.n498 VSUBS 0.006421f
C539 B.n499 VSUBS 0.006421f
C540 B.n500 VSUBS 0.006421f
C541 B.n501 VSUBS 0.006421f
C542 B.n502 VSUBS 0.006421f
C543 B.n503 VSUBS 0.006421f
C544 B.n504 VSUBS 0.006421f
C545 B.n505 VSUBS 0.006421f
C546 B.n506 VSUBS 0.006421f
C547 B.n507 VSUBS 0.006421f
C548 B.n508 VSUBS 0.006421f
C549 B.n509 VSUBS 0.006421f
C550 B.n510 VSUBS 0.006421f
C551 B.n511 VSUBS 0.006421f
C552 B.n512 VSUBS 0.006421f
C553 B.n513 VSUBS 0.006421f
C554 B.n514 VSUBS 0.006421f
C555 B.n515 VSUBS 0.006421f
C556 B.n516 VSUBS 0.006421f
C557 B.n517 VSUBS 0.006421f
C558 B.n518 VSUBS 0.006421f
C559 B.n519 VSUBS 0.006421f
C560 B.n520 VSUBS 0.006421f
C561 B.n521 VSUBS 0.006421f
C562 B.n522 VSUBS 0.006421f
C563 B.n523 VSUBS 0.006421f
C564 B.n524 VSUBS 0.006421f
C565 B.n525 VSUBS 0.006421f
C566 B.n526 VSUBS 0.006421f
C567 B.n527 VSUBS 0.006421f
C568 B.n528 VSUBS 0.006421f
C569 B.n529 VSUBS 0.006421f
C570 B.n530 VSUBS 0.006421f
C571 B.n531 VSUBS 0.006421f
C572 B.n532 VSUBS 0.006421f
C573 B.n533 VSUBS 0.006421f
C574 B.n534 VSUBS 0.006421f
C575 B.n535 VSUBS 0.006421f
C576 B.n536 VSUBS 0.006421f
C577 B.n537 VSUBS 0.006421f
C578 B.n538 VSUBS 0.006421f
C579 B.n539 VSUBS 0.006421f
C580 B.n540 VSUBS 0.006421f
C581 B.n541 VSUBS 0.006421f
C582 B.n542 VSUBS 0.006421f
C583 B.n543 VSUBS 0.006421f
C584 B.n544 VSUBS 0.006421f
C585 B.n545 VSUBS 0.006421f
C586 B.n546 VSUBS 0.006421f
C587 B.n547 VSUBS 0.006421f
C588 B.n548 VSUBS 0.006421f
C589 B.n549 VSUBS 0.006421f
C590 B.n550 VSUBS 0.006421f
C591 B.n551 VSUBS 0.006421f
C592 B.n552 VSUBS 0.006421f
C593 B.n553 VSUBS 0.006421f
C594 B.n554 VSUBS 0.015322f
C595 B.n555 VSUBS 0.015322f
C596 B.n556 VSUBS 0.015085f
C597 B.n557 VSUBS 0.006421f
C598 B.n558 VSUBS 0.006421f
C599 B.n559 VSUBS 0.006421f
C600 B.n560 VSUBS 0.006421f
C601 B.n561 VSUBS 0.006421f
C602 B.n562 VSUBS 0.006421f
C603 B.n563 VSUBS 0.006421f
C604 B.n564 VSUBS 0.006421f
C605 B.n565 VSUBS 0.006421f
C606 B.n566 VSUBS 0.006421f
C607 B.n567 VSUBS 0.006421f
C608 B.n568 VSUBS 0.006421f
C609 B.n569 VSUBS 0.006421f
C610 B.n570 VSUBS 0.006421f
C611 B.n571 VSUBS 0.006421f
C612 B.n572 VSUBS 0.006421f
C613 B.n573 VSUBS 0.006421f
C614 B.n574 VSUBS 0.006421f
C615 B.n575 VSUBS 0.006421f
C616 B.n576 VSUBS 0.006421f
C617 B.n577 VSUBS 0.006421f
C618 B.n578 VSUBS 0.006421f
C619 B.n579 VSUBS 0.006421f
C620 B.n580 VSUBS 0.006421f
C621 B.n581 VSUBS 0.006421f
C622 B.n582 VSUBS 0.006421f
C623 B.n583 VSUBS 0.00838f
C624 B.n584 VSUBS 0.008926f
C625 B.n585 VSUBS 0.017751f
C626 VDD1.n0 VSUBS 0.020362f
C627 VDD1.n1 VSUBS 0.019996f
C628 VDD1.n2 VSUBS 0.011061f
C629 VDD1.n3 VSUBS 0.025397f
C630 VDD1.n4 VSUBS 0.010745f
C631 VDD1.n5 VSUBS 0.011377f
C632 VDD1.n6 VSUBS 0.019996f
C633 VDD1.n7 VSUBS 0.010745f
C634 VDD1.n8 VSUBS 0.025397f
C635 VDD1.n9 VSUBS 0.011377f
C636 VDD1.n10 VSUBS 0.019996f
C637 VDD1.n11 VSUBS 0.010745f
C638 VDD1.n12 VSUBS 0.025397f
C639 VDD1.n13 VSUBS 0.011377f
C640 VDD1.n14 VSUBS 0.019996f
C641 VDD1.n15 VSUBS 0.010745f
C642 VDD1.n16 VSUBS 0.025397f
C643 VDD1.n17 VSUBS 0.011377f
C644 VDD1.n18 VSUBS 0.019996f
C645 VDD1.n19 VSUBS 0.010745f
C646 VDD1.n20 VSUBS 0.025397f
C647 VDD1.n21 VSUBS 0.011377f
C648 VDD1.n22 VSUBS 0.019996f
C649 VDD1.n23 VSUBS 0.010745f
C650 VDD1.n24 VSUBS 0.019048f
C651 VDD1.n25 VSUBS 0.016157f
C652 VDD1.t0 VSUBS 0.05432f
C653 VDD1.n26 VSUBS 0.134939f
C654 VDD1.n27 VSUBS 1.18419f
C655 VDD1.n28 VSUBS 0.010745f
C656 VDD1.n29 VSUBS 0.011377f
C657 VDD1.n30 VSUBS 0.025397f
C658 VDD1.n31 VSUBS 0.025397f
C659 VDD1.n32 VSUBS 0.011377f
C660 VDD1.n33 VSUBS 0.010745f
C661 VDD1.n34 VSUBS 0.019996f
C662 VDD1.n35 VSUBS 0.019996f
C663 VDD1.n36 VSUBS 0.010745f
C664 VDD1.n37 VSUBS 0.011377f
C665 VDD1.n38 VSUBS 0.025397f
C666 VDD1.n39 VSUBS 0.025397f
C667 VDD1.n40 VSUBS 0.011377f
C668 VDD1.n41 VSUBS 0.010745f
C669 VDD1.n42 VSUBS 0.019996f
C670 VDD1.n43 VSUBS 0.019996f
C671 VDD1.n44 VSUBS 0.010745f
C672 VDD1.n45 VSUBS 0.011377f
C673 VDD1.n46 VSUBS 0.025397f
C674 VDD1.n47 VSUBS 0.025397f
C675 VDD1.n48 VSUBS 0.011377f
C676 VDD1.n49 VSUBS 0.010745f
C677 VDD1.n50 VSUBS 0.019996f
C678 VDD1.n51 VSUBS 0.019996f
C679 VDD1.n52 VSUBS 0.010745f
C680 VDD1.n53 VSUBS 0.011377f
C681 VDD1.n54 VSUBS 0.025397f
C682 VDD1.n55 VSUBS 0.025397f
C683 VDD1.n56 VSUBS 0.011377f
C684 VDD1.n57 VSUBS 0.010745f
C685 VDD1.n58 VSUBS 0.019996f
C686 VDD1.n59 VSUBS 0.019996f
C687 VDD1.n60 VSUBS 0.010745f
C688 VDD1.n61 VSUBS 0.011377f
C689 VDD1.n62 VSUBS 0.025397f
C690 VDD1.n63 VSUBS 0.025397f
C691 VDD1.n64 VSUBS 0.011377f
C692 VDD1.n65 VSUBS 0.010745f
C693 VDD1.n66 VSUBS 0.019996f
C694 VDD1.n67 VSUBS 0.019996f
C695 VDD1.n68 VSUBS 0.010745f
C696 VDD1.n69 VSUBS 0.011377f
C697 VDD1.n70 VSUBS 0.025397f
C698 VDD1.n71 VSUBS 0.025397f
C699 VDD1.n72 VSUBS 0.056002f
C700 VDD1.n73 VSUBS 0.011061f
C701 VDD1.n74 VSUBS 0.010745f
C702 VDD1.n75 VSUBS 0.047859f
C703 VDD1.n76 VSUBS 0.042412f
C704 VDD1.n77 VSUBS 0.020362f
C705 VDD1.n78 VSUBS 0.019996f
C706 VDD1.n79 VSUBS 0.011061f
C707 VDD1.n80 VSUBS 0.025397f
C708 VDD1.n81 VSUBS 0.011377f
C709 VDD1.n82 VSUBS 0.019996f
C710 VDD1.n83 VSUBS 0.010745f
C711 VDD1.n84 VSUBS 0.025397f
C712 VDD1.n85 VSUBS 0.011377f
C713 VDD1.n86 VSUBS 0.019996f
C714 VDD1.n87 VSUBS 0.010745f
C715 VDD1.n88 VSUBS 0.025397f
C716 VDD1.n89 VSUBS 0.011377f
C717 VDD1.n90 VSUBS 0.019996f
C718 VDD1.n91 VSUBS 0.010745f
C719 VDD1.n92 VSUBS 0.025397f
C720 VDD1.n93 VSUBS 0.011377f
C721 VDD1.n94 VSUBS 0.019996f
C722 VDD1.n95 VSUBS 0.010745f
C723 VDD1.n96 VSUBS 0.025397f
C724 VDD1.n97 VSUBS 0.011377f
C725 VDD1.n98 VSUBS 0.019996f
C726 VDD1.n99 VSUBS 0.010745f
C727 VDD1.n100 VSUBS 0.019048f
C728 VDD1.n101 VSUBS 0.016157f
C729 VDD1.t1 VSUBS 0.05432f
C730 VDD1.n102 VSUBS 0.134939f
C731 VDD1.n103 VSUBS 1.18419f
C732 VDD1.n104 VSUBS 0.010745f
C733 VDD1.n105 VSUBS 0.011377f
C734 VDD1.n106 VSUBS 0.025397f
C735 VDD1.n107 VSUBS 0.025397f
C736 VDD1.n108 VSUBS 0.011377f
C737 VDD1.n109 VSUBS 0.010745f
C738 VDD1.n110 VSUBS 0.019996f
C739 VDD1.n111 VSUBS 0.019996f
C740 VDD1.n112 VSUBS 0.010745f
C741 VDD1.n113 VSUBS 0.011377f
C742 VDD1.n114 VSUBS 0.025397f
C743 VDD1.n115 VSUBS 0.025397f
C744 VDD1.n116 VSUBS 0.011377f
C745 VDD1.n117 VSUBS 0.010745f
C746 VDD1.n118 VSUBS 0.019996f
C747 VDD1.n119 VSUBS 0.019996f
C748 VDD1.n120 VSUBS 0.010745f
C749 VDD1.n121 VSUBS 0.011377f
C750 VDD1.n122 VSUBS 0.025397f
C751 VDD1.n123 VSUBS 0.025397f
C752 VDD1.n124 VSUBS 0.011377f
C753 VDD1.n125 VSUBS 0.010745f
C754 VDD1.n126 VSUBS 0.019996f
C755 VDD1.n127 VSUBS 0.019996f
C756 VDD1.n128 VSUBS 0.010745f
C757 VDD1.n129 VSUBS 0.011377f
C758 VDD1.n130 VSUBS 0.025397f
C759 VDD1.n131 VSUBS 0.025397f
C760 VDD1.n132 VSUBS 0.011377f
C761 VDD1.n133 VSUBS 0.010745f
C762 VDD1.n134 VSUBS 0.019996f
C763 VDD1.n135 VSUBS 0.019996f
C764 VDD1.n136 VSUBS 0.010745f
C765 VDD1.n137 VSUBS 0.011377f
C766 VDD1.n138 VSUBS 0.025397f
C767 VDD1.n139 VSUBS 0.025397f
C768 VDD1.n140 VSUBS 0.011377f
C769 VDD1.n141 VSUBS 0.010745f
C770 VDD1.n142 VSUBS 0.019996f
C771 VDD1.n143 VSUBS 0.019996f
C772 VDD1.n144 VSUBS 0.010745f
C773 VDD1.n145 VSUBS 0.010745f
C774 VDD1.n146 VSUBS 0.011377f
C775 VDD1.n147 VSUBS 0.025397f
C776 VDD1.n148 VSUBS 0.025397f
C777 VDD1.n149 VSUBS 0.056002f
C778 VDD1.n150 VSUBS 0.011061f
C779 VDD1.n151 VSUBS 0.010745f
C780 VDD1.n152 VSUBS 0.047859f
C781 VDD1.n153 VSUBS 0.614126f
C782 VP.t1 VSUBS 3.85025f
C783 VP.t0 VSUBS 3.47174f
C784 VP.n0 VSUBS 5.92329f
C785 VDD2.n0 VSUBS 0.020538f
C786 VDD2.n1 VSUBS 0.020169f
C787 VDD2.n2 VSUBS 0.011157f
C788 VDD2.n3 VSUBS 0.025617f
C789 VDD2.n4 VSUBS 0.011476f
C790 VDD2.n5 VSUBS 0.020169f
C791 VDD2.n6 VSUBS 0.010838f
C792 VDD2.n7 VSUBS 0.025617f
C793 VDD2.n8 VSUBS 0.011476f
C794 VDD2.n9 VSUBS 0.020169f
C795 VDD2.n10 VSUBS 0.010838f
C796 VDD2.n11 VSUBS 0.025617f
C797 VDD2.n12 VSUBS 0.011476f
C798 VDD2.n13 VSUBS 0.020169f
C799 VDD2.n14 VSUBS 0.010838f
C800 VDD2.n15 VSUBS 0.025617f
C801 VDD2.n16 VSUBS 0.011476f
C802 VDD2.n17 VSUBS 0.020169f
C803 VDD2.n18 VSUBS 0.010838f
C804 VDD2.n19 VSUBS 0.025617f
C805 VDD2.n20 VSUBS 0.011476f
C806 VDD2.n21 VSUBS 0.020169f
C807 VDD2.n22 VSUBS 0.010838f
C808 VDD2.n23 VSUBS 0.019213f
C809 VDD2.n24 VSUBS 0.016296f
C810 VDD2.t1 VSUBS 0.05479f
C811 VDD2.n25 VSUBS 0.136107f
C812 VDD2.n26 VSUBS 1.19445f
C813 VDD2.n27 VSUBS 0.010838f
C814 VDD2.n28 VSUBS 0.011476f
C815 VDD2.n29 VSUBS 0.025617f
C816 VDD2.n30 VSUBS 0.025617f
C817 VDD2.n31 VSUBS 0.011476f
C818 VDD2.n32 VSUBS 0.010838f
C819 VDD2.n33 VSUBS 0.020169f
C820 VDD2.n34 VSUBS 0.020169f
C821 VDD2.n35 VSUBS 0.010838f
C822 VDD2.n36 VSUBS 0.011476f
C823 VDD2.n37 VSUBS 0.025617f
C824 VDD2.n38 VSUBS 0.025617f
C825 VDD2.n39 VSUBS 0.011476f
C826 VDD2.n40 VSUBS 0.010838f
C827 VDD2.n41 VSUBS 0.020169f
C828 VDD2.n42 VSUBS 0.020169f
C829 VDD2.n43 VSUBS 0.010838f
C830 VDD2.n44 VSUBS 0.011476f
C831 VDD2.n45 VSUBS 0.025617f
C832 VDD2.n46 VSUBS 0.025617f
C833 VDD2.n47 VSUBS 0.011476f
C834 VDD2.n48 VSUBS 0.010838f
C835 VDD2.n49 VSUBS 0.020169f
C836 VDD2.n50 VSUBS 0.020169f
C837 VDD2.n51 VSUBS 0.010838f
C838 VDD2.n52 VSUBS 0.011476f
C839 VDD2.n53 VSUBS 0.025617f
C840 VDD2.n54 VSUBS 0.025617f
C841 VDD2.n55 VSUBS 0.011476f
C842 VDD2.n56 VSUBS 0.010838f
C843 VDD2.n57 VSUBS 0.020169f
C844 VDD2.n58 VSUBS 0.020169f
C845 VDD2.n59 VSUBS 0.010838f
C846 VDD2.n60 VSUBS 0.011476f
C847 VDD2.n61 VSUBS 0.025617f
C848 VDD2.n62 VSUBS 0.025617f
C849 VDD2.n63 VSUBS 0.011476f
C850 VDD2.n64 VSUBS 0.010838f
C851 VDD2.n65 VSUBS 0.020169f
C852 VDD2.n66 VSUBS 0.020169f
C853 VDD2.n67 VSUBS 0.010838f
C854 VDD2.n68 VSUBS 0.010838f
C855 VDD2.n69 VSUBS 0.011476f
C856 VDD2.n70 VSUBS 0.025617f
C857 VDD2.n71 VSUBS 0.025617f
C858 VDD2.n72 VSUBS 0.056487f
C859 VDD2.n73 VSUBS 0.011157f
C860 VDD2.n74 VSUBS 0.010838f
C861 VDD2.n75 VSUBS 0.048273f
C862 VDD2.n76 VSUBS 0.586144f
C863 VDD2.n77 VSUBS 0.020538f
C864 VDD2.n78 VSUBS 0.020169f
C865 VDD2.n79 VSUBS 0.011157f
C866 VDD2.n80 VSUBS 0.025617f
C867 VDD2.n81 VSUBS 0.010838f
C868 VDD2.n82 VSUBS 0.011476f
C869 VDD2.n83 VSUBS 0.020169f
C870 VDD2.n84 VSUBS 0.010838f
C871 VDD2.n85 VSUBS 0.025617f
C872 VDD2.n86 VSUBS 0.011476f
C873 VDD2.n87 VSUBS 0.020169f
C874 VDD2.n88 VSUBS 0.010838f
C875 VDD2.n89 VSUBS 0.025617f
C876 VDD2.n90 VSUBS 0.011476f
C877 VDD2.n91 VSUBS 0.020169f
C878 VDD2.n92 VSUBS 0.010838f
C879 VDD2.n93 VSUBS 0.025617f
C880 VDD2.n94 VSUBS 0.011476f
C881 VDD2.n95 VSUBS 0.020169f
C882 VDD2.n96 VSUBS 0.010838f
C883 VDD2.n97 VSUBS 0.025617f
C884 VDD2.n98 VSUBS 0.011476f
C885 VDD2.n99 VSUBS 0.020169f
C886 VDD2.n100 VSUBS 0.010838f
C887 VDD2.n101 VSUBS 0.019213f
C888 VDD2.n102 VSUBS 0.016296f
C889 VDD2.t0 VSUBS 0.05479f
C890 VDD2.n103 VSUBS 0.136107f
C891 VDD2.n104 VSUBS 1.19445f
C892 VDD2.n105 VSUBS 0.010838f
C893 VDD2.n106 VSUBS 0.011476f
C894 VDD2.n107 VSUBS 0.025617f
C895 VDD2.n108 VSUBS 0.025617f
C896 VDD2.n109 VSUBS 0.011476f
C897 VDD2.n110 VSUBS 0.010838f
C898 VDD2.n111 VSUBS 0.020169f
C899 VDD2.n112 VSUBS 0.020169f
C900 VDD2.n113 VSUBS 0.010838f
C901 VDD2.n114 VSUBS 0.011476f
C902 VDD2.n115 VSUBS 0.025617f
C903 VDD2.n116 VSUBS 0.025617f
C904 VDD2.n117 VSUBS 0.011476f
C905 VDD2.n118 VSUBS 0.010838f
C906 VDD2.n119 VSUBS 0.020169f
C907 VDD2.n120 VSUBS 0.020169f
C908 VDD2.n121 VSUBS 0.010838f
C909 VDD2.n122 VSUBS 0.011476f
C910 VDD2.n123 VSUBS 0.025617f
C911 VDD2.n124 VSUBS 0.025617f
C912 VDD2.n125 VSUBS 0.011476f
C913 VDD2.n126 VSUBS 0.010838f
C914 VDD2.n127 VSUBS 0.020169f
C915 VDD2.n128 VSUBS 0.020169f
C916 VDD2.n129 VSUBS 0.010838f
C917 VDD2.n130 VSUBS 0.011476f
C918 VDD2.n131 VSUBS 0.025617f
C919 VDD2.n132 VSUBS 0.025617f
C920 VDD2.n133 VSUBS 0.011476f
C921 VDD2.n134 VSUBS 0.010838f
C922 VDD2.n135 VSUBS 0.020169f
C923 VDD2.n136 VSUBS 0.020169f
C924 VDD2.n137 VSUBS 0.010838f
C925 VDD2.n138 VSUBS 0.011476f
C926 VDD2.n139 VSUBS 0.025617f
C927 VDD2.n140 VSUBS 0.025617f
C928 VDD2.n141 VSUBS 0.011476f
C929 VDD2.n142 VSUBS 0.010838f
C930 VDD2.n143 VSUBS 0.020169f
C931 VDD2.n144 VSUBS 0.020169f
C932 VDD2.n145 VSUBS 0.010838f
C933 VDD2.n146 VSUBS 0.011476f
C934 VDD2.n147 VSUBS 0.025617f
C935 VDD2.n148 VSUBS 0.025617f
C936 VDD2.n149 VSUBS 0.056487f
C937 VDD2.n150 VSUBS 0.011157f
C938 VDD2.n151 VSUBS 0.010838f
C939 VDD2.n152 VSUBS 0.048273f
C940 VDD2.n153 VSUBS 0.042125f
C941 VDD2.n154 VSUBS 2.47641f
C942 VTAIL.n0 VSUBS 0.028881f
C943 VTAIL.n1 VSUBS 0.028362f
C944 VTAIL.n2 VSUBS 0.015689f
C945 VTAIL.n3 VSUBS 0.036023f
C946 VTAIL.n4 VSUBS 0.016137f
C947 VTAIL.n5 VSUBS 0.028362f
C948 VTAIL.n6 VSUBS 0.01524f
C949 VTAIL.n7 VSUBS 0.036023f
C950 VTAIL.n8 VSUBS 0.016137f
C951 VTAIL.n9 VSUBS 0.028362f
C952 VTAIL.n10 VSUBS 0.01524f
C953 VTAIL.n11 VSUBS 0.036023f
C954 VTAIL.n12 VSUBS 0.016137f
C955 VTAIL.n13 VSUBS 0.028362f
C956 VTAIL.n14 VSUBS 0.01524f
C957 VTAIL.n15 VSUBS 0.036023f
C958 VTAIL.n16 VSUBS 0.016137f
C959 VTAIL.n17 VSUBS 0.028362f
C960 VTAIL.n18 VSUBS 0.01524f
C961 VTAIL.n19 VSUBS 0.036023f
C962 VTAIL.n20 VSUBS 0.016137f
C963 VTAIL.n21 VSUBS 0.028362f
C964 VTAIL.n22 VSUBS 0.01524f
C965 VTAIL.n23 VSUBS 0.027017f
C966 VTAIL.n24 VSUBS 0.022916f
C967 VTAIL.t1 VSUBS 0.077046f
C968 VTAIL.n25 VSUBS 0.191393f
C969 VTAIL.n26 VSUBS 1.67963f
C970 VTAIL.n27 VSUBS 0.01524f
C971 VTAIL.n28 VSUBS 0.016137f
C972 VTAIL.n29 VSUBS 0.036023f
C973 VTAIL.n30 VSUBS 0.036023f
C974 VTAIL.n31 VSUBS 0.016137f
C975 VTAIL.n32 VSUBS 0.01524f
C976 VTAIL.n33 VSUBS 0.028362f
C977 VTAIL.n34 VSUBS 0.028362f
C978 VTAIL.n35 VSUBS 0.01524f
C979 VTAIL.n36 VSUBS 0.016137f
C980 VTAIL.n37 VSUBS 0.036023f
C981 VTAIL.n38 VSUBS 0.036023f
C982 VTAIL.n39 VSUBS 0.016137f
C983 VTAIL.n40 VSUBS 0.01524f
C984 VTAIL.n41 VSUBS 0.028362f
C985 VTAIL.n42 VSUBS 0.028362f
C986 VTAIL.n43 VSUBS 0.01524f
C987 VTAIL.n44 VSUBS 0.016137f
C988 VTAIL.n45 VSUBS 0.036023f
C989 VTAIL.n46 VSUBS 0.036023f
C990 VTAIL.n47 VSUBS 0.016137f
C991 VTAIL.n48 VSUBS 0.01524f
C992 VTAIL.n49 VSUBS 0.028362f
C993 VTAIL.n50 VSUBS 0.028362f
C994 VTAIL.n51 VSUBS 0.01524f
C995 VTAIL.n52 VSUBS 0.016137f
C996 VTAIL.n53 VSUBS 0.036023f
C997 VTAIL.n54 VSUBS 0.036023f
C998 VTAIL.n55 VSUBS 0.016137f
C999 VTAIL.n56 VSUBS 0.01524f
C1000 VTAIL.n57 VSUBS 0.028362f
C1001 VTAIL.n58 VSUBS 0.028362f
C1002 VTAIL.n59 VSUBS 0.01524f
C1003 VTAIL.n60 VSUBS 0.016137f
C1004 VTAIL.n61 VSUBS 0.036023f
C1005 VTAIL.n62 VSUBS 0.036023f
C1006 VTAIL.n63 VSUBS 0.016137f
C1007 VTAIL.n64 VSUBS 0.01524f
C1008 VTAIL.n65 VSUBS 0.028362f
C1009 VTAIL.n66 VSUBS 0.028362f
C1010 VTAIL.n67 VSUBS 0.01524f
C1011 VTAIL.n68 VSUBS 0.01524f
C1012 VTAIL.n69 VSUBS 0.016137f
C1013 VTAIL.n70 VSUBS 0.036023f
C1014 VTAIL.n71 VSUBS 0.036023f
C1015 VTAIL.n72 VSUBS 0.079432f
C1016 VTAIL.n73 VSUBS 0.015689f
C1017 VTAIL.n74 VSUBS 0.01524f
C1018 VTAIL.n75 VSUBS 0.067882f
C1019 VTAIL.n76 VSUBS 0.039671f
C1020 VTAIL.n77 VSUBS 1.899f
C1021 VTAIL.n78 VSUBS 0.028881f
C1022 VTAIL.n79 VSUBS 0.028362f
C1023 VTAIL.n80 VSUBS 0.015689f
C1024 VTAIL.n81 VSUBS 0.036023f
C1025 VTAIL.n82 VSUBS 0.01524f
C1026 VTAIL.n83 VSUBS 0.016137f
C1027 VTAIL.n84 VSUBS 0.028362f
C1028 VTAIL.n85 VSUBS 0.01524f
C1029 VTAIL.n86 VSUBS 0.036023f
C1030 VTAIL.n87 VSUBS 0.016137f
C1031 VTAIL.n88 VSUBS 0.028362f
C1032 VTAIL.n89 VSUBS 0.01524f
C1033 VTAIL.n90 VSUBS 0.036023f
C1034 VTAIL.n91 VSUBS 0.016137f
C1035 VTAIL.n92 VSUBS 0.028362f
C1036 VTAIL.n93 VSUBS 0.01524f
C1037 VTAIL.n94 VSUBS 0.036023f
C1038 VTAIL.n95 VSUBS 0.016137f
C1039 VTAIL.n96 VSUBS 0.028362f
C1040 VTAIL.n97 VSUBS 0.01524f
C1041 VTAIL.n98 VSUBS 0.036023f
C1042 VTAIL.n99 VSUBS 0.016137f
C1043 VTAIL.n100 VSUBS 0.028362f
C1044 VTAIL.n101 VSUBS 0.01524f
C1045 VTAIL.n102 VSUBS 0.027017f
C1046 VTAIL.n103 VSUBS 0.022916f
C1047 VTAIL.t3 VSUBS 0.077046f
C1048 VTAIL.n104 VSUBS 0.191393f
C1049 VTAIL.n105 VSUBS 1.67963f
C1050 VTAIL.n106 VSUBS 0.01524f
C1051 VTAIL.n107 VSUBS 0.016137f
C1052 VTAIL.n108 VSUBS 0.036023f
C1053 VTAIL.n109 VSUBS 0.036023f
C1054 VTAIL.n110 VSUBS 0.016137f
C1055 VTAIL.n111 VSUBS 0.01524f
C1056 VTAIL.n112 VSUBS 0.028362f
C1057 VTAIL.n113 VSUBS 0.028362f
C1058 VTAIL.n114 VSUBS 0.01524f
C1059 VTAIL.n115 VSUBS 0.016137f
C1060 VTAIL.n116 VSUBS 0.036023f
C1061 VTAIL.n117 VSUBS 0.036023f
C1062 VTAIL.n118 VSUBS 0.016137f
C1063 VTAIL.n119 VSUBS 0.01524f
C1064 VTAIL.n120 VSUBS 0.028362f
C1065 VTAIL.n121 VSUBS 0.028362f
C1066 VTAIL.n122 VSUBS 0.01524f
C1067 VTAIL.n123 VSUBS 0.016137f
C1068 VTAIL.n124 VSUBS 0.036023f
C1069 VTAIL.n125 VSUBS 0.036023f
C1070 VTAIL.n126 VSUBS 0.016137f
C1071 VTAIL.n127 VSUBS 0.01524f
C1072 VTAIL.n128 VSUBS 0.028362f
C1073 VTAIL.n129 VSUBS 0.028362f
C1074 VTAIL.n130 VSUBS 0.01524f
C1075 VTAIL.n131 VSUBS 0.016137f
C1076 VTAIL.n132 VSUBS 0.036023f
C1077 VTAIL.n133 VSUBS 0.036023f
C1078 VTAIL.n134 VSUBS 0.016137f
C1079 VTAIL.n135 VSUBS 0.01524f
C1080 VTAIL.n136 VSUBS 0.028362f
C1081 VTAIL.n137 VSUBS 0.028362f
C1082 VTAIL.n138 VSUBS 0.01524f
C1083 VTAIL.n139 VSUBS 0.016137f
C1084 VTAIL.n140 VSUBS 0.036023f
C1085 VTAIL.n141 VSUBS 0.036023f
C1086 VTAIL.n142 VSUBS 0.016137f
C1087 VTAIL.n143 VSUBS 0.01524f
C1088 VTAIL.n144 VSUBS 0.028362f
C1089 VTAIL.n145 VSUBS 0.028362f
C1090 VTAIL.n146 VSUBS 0.01524f
C1091 VTAIL.n147 VSUBS 0.016137f
C1092 VTAIL.n148 VSUBS 0.036023f
C1093 VTAIL.n149 VSUBS 0.036023f
C1094 VTAIL.n150 VSUBS 0.079432f
C1095 VTAIL.n151 VSUBS 0.015689f
C1096 VTAIL.n152 VSUBS 0.01524f
C1097 VTAIL.n153 VSUBS 0.067882f
C1098 VTAIL.n154 VSUBS 0.039671f
C1099 VTAIL.n155 VSUBS 1.9313f
C1100 VTAIL.n156 VSUBS 0.028881f
C1101 VTAIL.n157 VSUBS 0.028362f
C1102 VTAIL.n158 VSUBS 0.015689f
C1103 VTAIL.n159 VSUBS 0.036023f
C1104 VTAIL.n160 VSUBS 0.01524f
C1105 VTAIL.n161 VSUBS 0.016137f
C1106 VTAIL.n162 VSUBS 0.028362f
C1107 VTAIL.n163 VSUBS 0.01524f
C1108 VTAIL.n164 VSUBS 0.036023f
C1109 VTAIL.n165 VSUBS 0.016137f
C1110 VTAIL.n166 VSUBS 0.028362f
C1111 VTAIL.n167 VSUBS 0.01524f
C1112 VTAIL.n168 VSUBS 0.036023f
C1113 VTAIL.n169 VSUBS 0.016137f
C1114 VTAIL.n170 VSUBS 0.028362f
C1115 VTAIL.n171 VSUBS 0.01524f
C1116 VTAIL.n172 VSUBS 0.036023f
C1117 VTAIL.n173 VSUBS 0.016137f
C1118 VTAIL.n174 VSUBS 0.028362f
C1119 VTAIL.n175 VSUBS 0.01524f
C1120 VTAIL.n176 VSUBS 0.036023f
C1121 VTAIL.n177 VSUBS 0.016137f
C1122 VTAIL.n178 VSUBS 0.028362f
C1123 VTAIL.n179 VSUBS 0.01524f
C1124 VTAIL.n180 VSUBS 0.027017f
C1125 VTAIL.n181 VSUBS 0.022916f
C1126 VTAIL.t0 VSUBS 0.077046f
C1127 VTAIL.n182 VSUBS 0.191393f
C1128 VTAIL.n183 VSUBS 1.67963f
C1129 VTAIL.n184 VSUBS 0.01524f
C1130 VTAIL.n185 VSUBS 0.016137f
C1131 VTAIL.n186 VSUBS 0.036023f
C1132 VTAIL.n187 VSUBS 0.036023f
C1133 VTAIL.n188 VSUBS 0.016137f
C1134 VTAIL.n189 VSUBS 0.01524f
C1135 VTAIL.n190 VSUBS 0.028362f
C1136 VTAIL.n191 VSUBS 0.028362f
C1137 VTAIL.n192 VSUBS 0.01524f
C1138 VTAIL.n193 VSUBS 0.016137f
C1139 VTAIL.n194 VSUBS 0.036023f
C1140 VTAIL.n195 VSUBS 0.036023f
C1141 VTAIL.n196 VSUBS 0.016137f
C1142 VTAIL.n197 VSUBS 0.01524f
C1143 VTAIL.n198 VSUBS 0.028362f
C1144 VTAIL.n199 VSUBS 0.028362f
C1145 VTAIL.n200 VSUBS 0.01524f
C1146 VTAIL.n201 VSUBS 0.016137f
C1147 VTAIL.n202 VSUBS 0.036023f
C1148 VTAIL.n203 VSUBS 0.036023f
C1149 VTAIL.n204 VSUBS 0.016137f
C1150 VTAIL.n205 VSUBS 0.01524f
C1151 VTAIL.n206 VSUBS 0.028362f
C1152 VTAIL.n207 VSUBS 0.028362f
C1153 VTAIL.n208 VSUBS 0.01524f
C1154 VTAIL.n209 VSUBS 0.016137f
C1155 VTAIL.n210 VSUBS 0.036023f
C1156 VTAIL.n211 VSUBS 0.036023f
C1157 VTAIL.n212 VSUBS 0.016137f
C1158 VTAIL.n213 VSUBS 0.01524f
C1159 VTAIL.n214 VSUBS 0.028362f
C1160 VTAIL.n215 VSUBS 0.028362f
C1161 VTAIL.n216 VSUBS 0.01524f
C1162 VTAIL.n217 VSUBS 0.016137f
C1163 VTAIL.n218 VSUBS 0.036023f
C1164 VTAIL.n219 VSUBS 0.036023f
C1165 VTAIL.n220 VSUBS 0.016137f
C1166 VTAIL.n221 VSUBS 0.01524f
C1167 VTAIL.n222 VSUBS 0.028362f
C1168 VTAIL.n223 VSUBS 0.028362f
C1169 VTAIL.n224 VSUBS 0.01524f
C1170 VTAIL.n225 VSUBS 0.016137f
C1171 VTAIL.n226 VSUBS 0.036023f
C1172 VTAIL.n227 VSUBS 0.036023f
C1173 VTAIL.n228 VSUBS 0.079432f
C1174 VTAIL.n229 VSUBS 0.015689f
C1175 VTAIL.n230 VSUBS 0.01524f
C1176 VTAIL.n231 VSUBS 0.067882f
C1177 VTAIL.n232 VSUBS 0.039671f
C1178 VTAIL.n233 VSUBS 1.78083f
C1179 VTAIL.n234 VSUBS 0.028881f
C1180 VTAIL.n235 VSUBS 0.028362f
C1181 VTAIL.n236 VSUBS 0.015689f
C1182 VTAIL.n237 VSUBS 0.036023f
C1183 VTAIL.n238 VSUBS 0.016137f
C1184 VTAIL.n239 VSUBS 0.028362f
C1185 VTAIL.n240 VSUBS 0.01524f
C1186 VTAIL.n241 VSUBS 0.036023f
C1187 VTAIL.n242 VSUBS 0.016137f
C1188 VTAIL.n243 VSUBS 0.028362f
C1189 VTAIL.n244 VSUBS 0.01524f
C1190 VTAIL.n245 VSUBS 0.036023f
C1191 VTAIL.n246 VSUBS 0.016137f
C1192 VTAIL.n247 VSUBS 0.028362f
C1193 VTAIL.n248 VSUBS 0.01524f
C1194 VTAIL.n249 VSUBS 0.036023f
C1195 VTAIL.n250 VSUBS 0.016137f
C1196 VTAIL.n251 VSUBS 0.028362f
C1197 VTAIL.n252 VSUBS 0.01524f
C1198 VTAIL.n253 VSUBS 0.036023f
C1199 VTAIL.n254 VSUBS 0.016137f
C1200 VTAIL.n255 VSUBS 0.028362f
C1201 VTAIL.n256 VSUBS 0.01524f
C1202 VTAIL.n257 VSUBS 0.027017f
C1203 VTAIL.n258 VSUBS 0.022916f
C1204 VTAIL.t2 VSUBS 0.077046f
C1205 VTAIL.n259 VSUBS 0.191393f
C1206 VTAIL.n260 VSUBS 1.67963f
C1207 VTAIL.n261 VSUBS 0.01524f
C1208 VTAIL.n262 VSUBS 0.016137f
C1209 VTAIL.n263 VSUBS 0.036023f
C1210 VTAIL.n264 VSUBS 0.036023f
C1211 VTAIL.n265 VSUBS 0.016137f
C1212 VTAIL.n266 VSUBS 0.01524f
C1213 VTAIL.n267 VSUBS 0.028362f
C1214 VTAIL.n268 VSUBS 0.028362f
C1215 VTAIL.n269 VSUBS 0.01524f
C1216 VTAIL.n270 VSUBS 0.016137f
C1217 VTAIL.n271 VSUBS 0.036023f
C1218 VTAIL.n272 VSUBS 0.036023f
C1219 VTAIL.n273 VSUBS 0.016137f
C1220 VTAIL.n274 VSUBS 0.01524f
C1221 VTAIL.n275 VSUBS 0.028362f
C1222 VTAIL.n276 VSUBS 0.028362f
C1223 VTAIL.n277 VSUBS 0.01524f
C1224 VTAIL.n278 VSUBS 0.016137f
C1225 VTAIL.n279 VSUBS 0.036023f
C1226 VTAIL.n280 VSUBS 0.036023f
C1227 VTAIL.n281 VSUBS 0.016137f
C1228 VTAIL.n282 VSUBS 0.01524f
C1229 VTAIL.n283 VSUBS 0.028362f
C1230 VTAIL.n284 VSUBS 0.028362f
C1231 VTAIL.n285 VSUBS 0.01524f
C1232 VTAIL.n286 VSUBS 0.016137f
C1233 VTAIL.n287 VSUBS 0.036023f
C1234 VTAIL.n288 VSUBS 0.036023f
C1235 VTAIL.n289 VSUBS 0.016137f
C1236 VTAIL.n290 VSUBS 0.01524f
C1237 VTAIL.n291 VSUBS 0.028362f
C1238 VTAIL.n292 VSUBS 0.028362f
C1239 VTAIL.n293 VSUBS 0.01524f
C1240 VTAIL.n294 VSUBS 0.016137f
C1241 VTAIL.n295 VSUBS 0.036023f
C1242 VTAIL.n296 VSUBS 0.036023f
C1243 VTAIL.n297 VSUBS 0.016137f
C1244 VTAIL.n298 VSUBS 0.01524f
C1245 VTAIL.n299 VSUBS 0.028362f
C1246 VTAIL.n300 VSUBS 0.028362f
C1247 VTAIL.n301 VSUBS 0.01524f
C1248 VTAIL.n302 VSUBS 0.01524f
C1249 VTAIL.n303 VSUBS 0.016137f
C1250 VTAIL.n304 VSUBS 0.036023f
C1251 VTAIL.n305 VSUBS 0.036023f
C1252 VTAIL.n306 VSUBS 0.079432f
C1253 VTAIL.n307 VSUBS 0.015689f
C1254 VTAIL.n308 VSUBS 0.01524f
C1255 VTAIL.n309 VSUBS 0.067882f
C1256 VTAIL.n310 VSUBS 0.039671f
C1257 VTAIL.n311 VSUBS 1.69496f
C1258 VN.t0 VSUBS 3.34993f
C1259 VN.t1 VSUBS 3.72007f
.ends

