* NGSPICE file created from diff_pair_sample_1643.ext - technology: sky130A

.subckt diff_pair_sample_1643 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4883 pd=9.35 as=3.5178 ps=18.82 w=9.02 l=0.65
X1 VDD1.t2 VP.t1 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.4883 pd=9.35 as=3.5178 ps=18.82 w=9.02 l=0.65
X2 VTAIL.t1 VN.t0 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.5178 pd=18.82 as=1.4883 ps=9.35 w=9.02 l=0.65
X3 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=3.5178 pd=18.82 as=0 ps=0 w=9.02 l=0.65
X4 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=3.5178 pd=18.82 as=0 ps=0 w=9.02 l=0.65
X5 VTAIL.t7 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.5178 pd=18.82 as=1.4883 ps=9.35 w=9.02 l=0.65
X6 VTAIL.t5 VP.t3 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=3.5178 pd=18.82 as=1.4883 ps=9.35 w=9.02 l=0.65
X7 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.5178 pd=18.82 as=0 ps=0 w=9.02 l=0.65
X8 VTAIL.t2 VN.t1 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.5178 pd=18.82 as=1.4883 ps=9.35 w=9.02 l=0.65
X9 VDD2.t1 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4883 pd=9.35 as=3.5178 ps=18.82 w=9.02 l=0.65
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.5178 pd=18.82 as=0 ps=0 w=9.02 l=0.65
X11 VDD2.t0 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.4883 pd=9.35 as=3.5178 ps=18.82 w=9.02 l=0.65
R0 VP.n1 VP.t3 415.865
R1 VP.n1 VP.t1 415.817
R2 VP.n3 VP.t2 394.87
R3 VP.n5 VP.t0 394.87
R4 VP.n6 VP.n5 161.3
R5 VP.n4 VP.n0 161.3
R6 VP.n3 VP.n2 161.3
R7 VP.n2 VP.n1 82.6242
R8 VP.n4 VP.n3 24.1005
R9 VP.n5 VP.n4 24.1005
R10 VP.n2 VP.n0 0.189894
R11 VP.n6 VP.n0 0.189894
R12 VP VP.n6 0.0516364
R13 VTAIL.n5 VTAIL.t5 51.4418
R14 VTAIL.n4 VTAIL.t3 51.4418
R15 VTAIL.n3 VTAIL.t1 51.4418
R16 VTAIL.n7 VTAIL.t0 51.4416
R17 VTAIL.n0 VTAIL.t2 51.4416
R18 VTAIL.n1 VTAIL.t4 51.4416
R19 VTAIL.n2 VTAIL.t7 51.4416
R20 VTAIL.n6 VTAIL.t6 51.4416
R21 VTAIL.n7 VTAIL.n6 20.9876
R22 VTAIL.n3 VTAIL.n2 20.9876
R23 VTAIL.n4 VTAIL.n3 0.845328
R24 VTAIL.n6 VTAIL.n5 0.845328
R25 VTAIL.n2 VTAIL.n1 0.845328
R26 VTAIL VTAIL.n0 0.481103
R27 VTAIL.n5 VTAIL.n4 0.470328
R28 VTAIL.n1 VTAIL.n0 0.470328
R29 VTAIL VTAIL.n7 0.364724
R30 VDD1 VDD1.n1 100.475
R31 VDD1 VDD1.n0 65.9835
R32 VDD1.n0 VDD1.t0 2.19562
R33 VDD1.n0 VDD1.t2 2.19562
R34 VDD1.n1 VDD1.t1 2.19562
R35 VDD1.n1 VDD1.t3 2.19562
R36 B.n519 B.n518 585
R37 B.n520 B.n519 585
R38 B.n223 B.n72 585
R39 B.n222 B.n221 585
R40 B.n220 B.n219 585
R41 B.n218 B.n217 585
R42 B.n216 B.n215 585
R43 B.n214 B.n213 585
R44 B.n212 B.n211 585
R45 B.n210 B.n209 585
R46 B.n208 B.n207 585
R47 B.n206 B.n205 585
R48 B.n204 B.n203 585
R49 B.n202 B.n201 585
R50 B.n200 B.n199 585
R51 B.n198 B.n197 585
R52 B.n196 B.n195 585
R53 B.n194 B.n193 585
R54 B.n192 B.n191 585
R55 B.n190 B.n189 585
R56 B.n188 B.n187 585
R57 B.n186 B.n185 585
R58 B.n184 B.n183 585
R59 B.n182 B.n181 585
R60 B.n180 B.n179 585
R61 B.n178 B.n177 585
R62 B.n176 B.n175 585
R63 B.n174 B.n173 585
R64 B.n172 B.n171 585
R65 B.n170 B.n169 585
R66 B.n168 B.n167 585
R67 B.n166 B.n165 585
R68 B.n164 B.n163 585
R69 B.n162 B.n161 585
R70 B.n160 B.n159 585
R71 B.n158 B.n157 585
R72 B.n156 B.n155 585
R73 B.n154 B.n153 585
R74 B.n152 B.n151 585
R75 B.n150 B.n149 585
R76 B.n148 B.n147 585
R77 B.n146 B.n145 585
R78 B.n144 B.n143 585
R79 B.n141 B.n140 585
R80 B.n139 B.n138 585
R81 B.n137 B.n136 585
R82 B.n135 B.n134 585
R83 B.n133 B.n132 585
R84 B.n131 B.n130 585
R85 B.n129 B.n128 585
R86 B.n127 B.n126 585
R87 B.n125 B.n124 585
R88 B.n123 B.n122 585
R89 B.n121 B.n120 585
R90 B.n119 B.n118 585
R91 B.n117 B.n116 585
R92 B.n115 B.n114 585
R93 B.n113 B.n112 585
R94 B.n111 B.n110 585
R95 B.n109 B.n108 585
R96 B.n107 B.n106 585
R97 B.n105 B.n104 585
R98 B.n103 B.n102 585
R99 B.n101 B.n100 585
R100 B.n99 B.n98 585
R101 B.n97 B.n96 585
R102 B.n95 B.n94 585
R103 B.n93 B.n92 585
R104 B.n91 B.n90 585
R105 B.n89 B.n88 585
R106 B.n87 B.n86 585
R107 B.n85 B.n84 585
R108 B.n83 B.n82 585
R109 B.n81 B.n80 585
R110 B.n79 B.n78 585
R111 B.n33 B.n32 585
R112 B.n517 B.n34 585
R113 B.n521 B.n34 585
R114 B.n516 B.n515 585
R115 B.n515 B.n30 585
R116 B.n514 B.n29 585
R117 B.n527 B.n29 585
R118 B.n513 B.n28 585
R119 B.n528 B.n28 585
R120 B.n512 B.n27 585
R121 B.n529 B.n27 585
R122 B.n511 B.n510 585
R123 B.n510 B.n23 585
R124 B.n509 B.n22 585
R125 B.n535 B.n22 585
R126 B.n508 B.n21 585
R127 B.n536 B.n21 585
R128 B.n507 B.n20 585
R129 B.n537 B.n20 585
R130 B.n506 B.n505 585
R131 B.n505 B.n16 585
R132 B.n504 B.n15 585
R133 B.n543 B.n15 585
R134 B.n503 B.n14 585
R135 B.n544 B.n14 585
R136 B.n502 B.n13 585
R137 B.n545 B.n13 585
R138 B.n501 B.n500 585
R139 B.n500 B.n12 585
R140 B.n499 B.n498 585
R141 B.n499 B.n8 585
R142 B.n497 B.n7 585
R143 B.n552 B.n7 585
R144 B.n496 B.n6 585
R145 B.n553 B.n6 585
R146 B.n495 B.n5 585
R147 B.n554 B.n5 585
R148 B.n494 B.n493 585
R149 B.n493 B.n4 585
R150 B.n492 B.n224 585
R151 B.n492 B.n491 585
R152 B.n481 B.n225 585
R153 B.n484 B.n225 585
R154 B.n483 B.n482 585
R155 B.n485 B.n483 585
R156 B.n480 B.n230 585
R157 B.n230 B.n229 585
R158 B.n479 B.n478 585
R159 B.n478 B.n477 585
R160 B.n232 B.n231 585
R161 B.n233 B.n232 585
R162 B.n470 B.n469 585
R163 B.n471 B.n470 585
R164 B.n468 B.n238 585
R165 B.n238 B.n237 585
R166 B.n467 B.n466 585
R167 B.n466 B.n465 585
R168 B.n240 B.n239 585
R169 B.n241 B.n240 585
R170 B.n458 B.n457 585
R171 B.n459 B.n458 585
R172 B.n456 B.n246 585
R173 B.n246 B.n245 585
R174 B.n455 B.n454 585
R175 B.n454 B.n453 585
R176 B.n248 B.n247 585
R177 B.n249 B.n248 585
R178 B.n446 B.n445 585
R179 B.n447 B.n446 585
R180 B.n252 B.n251 585
R181 B.n298 B.n297 585
R182 B.n299 B.n295 585
R183 B.n295 B.n253 585
R184 B.n301 B.n300 585
R185 B.n303 B.n294 585
R186 B.n306 B.n305 585
R187 B.n307 B.n293 585
R188 B.n309 B.n308 585
R189 B.n311 B.n292 585
R190 B.n314 B.n313 585
R191 B.n315 B.n291 585
R192 B.n317 B.n316 585
R193 B.n319 B.n290 585
R194 B.n322 B.n321 585
R195 B.n323 B.n289 585
R196 B.n325 B.n324 585
R197 B.n327 B.n288 585
R198 B.n330 B.n329 585
R199 B.n331 B.n287 585
R200 B.n333 B.n332 585
R201 B.n335 B.n286 585
R202 B.n338 B.n337 585
R203 B.n339 B.n285 585
R204 B.n341 B.n340 585
R205 B.n343 B.n284 585
R206 B.n346 B.n345 585
R207 B.n347 B.n283 585
R208 B.n349 B.n348 585
R209 B.n351 B.n282 585
R210 B.n354 B.n353 585
R211 B.n355 B.n281 585
R212 B.n357 B.n356 585
R213 B.n359 B.n280 585
R214 B.n362 B.n361 585
R215 B.n363 B.n276 585
R216 B.n365 B.n364 585
R217 B.n367 B.n275 585
R218 B.n370 B.n369 585
R219 B.n371 B.n274 585
R220 B.n373 B.n372 585
R221 B.n375 B.n273 585
R222 B.n378 B.n377 585
R223 B.n380 B.n270 585
R224 B.n382 B.n381 585
R225 B.n384 B.n269 585
R226 B.n387 B.n386 585
R227 B.n388 B.n268 585
R228 B.n390 B.n389 585
R229 B.n392 B.n267 585
R230 B.n395 B.n394 585
R231 B.n396 B.n266 585
R232 B.n398 B.n397 585
R233 B.n400 B.n265 585
R234 B.n403 B.n402 585
R235 B.n404 B.n264 585
R236 B.n406 B.n405 585
R237 B.n408 B.n263 585
R238 B.n411 B.n410 585
R239 B.n412 B.n262 585
R240 B.n414 B.n413 585
R241 B.n416 B.n261 585
R242 B.n419 B.n418 585
R243 B.n420 B.n260 585
R244 B.n422 B.n421 585
R245 B.n424 B.n259 585
R246 B.n427 B.n426 585
R247 B.n428 B.n258 585
R248 B.n430 B.n429 585
R249 B.n432 B.n257 585
R250 B.n435 B.n434 585
R251 B.n436 B.n256 585
R252 B.n438 B.n437 585
R253 B.n440 B.n255 585
R254 B.n443 B.n442 585
R255 B.n444 B.n254 585
R256 B.n449 B.n448 585
R257 B.n448 B.n447 585
R258 B.n450 B.n250 585
R259 B.n250 B.n249 585
R260 B.n452 B.n451 585
R261 B.n453 B.n452 585
R262 B.n244 B.n243 585
R263 B.n245 B.n244 585
R264 B.n461 B.n460 585
R265 B.n460 B.n459 585
R266 B.n462 B.n242 585
R267 B.n242 B.n241 585
R268 B.n464 B.n463 585
R269 B.n465 B.n464 585
R270 B.n236 B.n235 585
R271 B.n237 B.n236 585
R272 B.n473 B.n472 585
R273 B.n472 B.n471 585
R274 B.n474 B.n234 585
R275 B.n234 B.n233 585
R276 B.n476 B.n475 585
R277 B.n477 B.n476 585
R278 B.n228 B.n227 585
R279 B.n229 B.n228 585
R280 B.n487 B.n486 585
R281 B.n486 B.n485 585
R282 B.n488 B.n226 585
R283 B.n484 B.n226 585
R284 B.n490 B.n489 585
R285 B.n491 B.n490 585
R286 B.n3 B.n0 585
R287 B.n4 B.n3 585
R288 B.n551 B.n1 585
R289 B.n552 B.n551 585
R290 B.n550 B.n549 585
R291 B.n550 B.n8 585
R292 B.n548 B.n9 585
R293 B.n12 B.n9 585
R294 B.n547 B.n546 585
R295 B.n546 B.n545 585
R296 B.n11 B.n10 585
R297 B.n544 B.n11 585
R298 B.n542 B.n541 585
R299 B.n543 B.n542 585
R300 B.n540 B.n17 585
R301 B.n17 B.n16 585
R302 B.n539 B.n538 585
R303 B.n538 B.n537 585
R304 B.n19 B.n18 585
R305 B.n536 B.n19 585
R306 B.n534 B.n533 585
R307 B.n535 B.n534 585
R308 B.n532 B.n24 585
R309 B.n24 B.n23 585
R310 B.n531 B.n530 585
R311 B.n530 B.n529 585
R312 B.n26 B.n25 585
R313 B.n528 B.n26 585
R314 B.n526 B.n525 585
R315 B.n527 B.n526 585
R316 B.n524 B.n31 585
R317 B.n31 B.n30 585
R318 B.n523 B.n522 585
R319 B.n522 B.n521 585
R320 B.n555 B.n554 585
R321 B.n553 B.n2 585
R322 B.n522 B.n33 564.573
R323 B.n519 B.n34 564.573
R324 B.n446 B.n254 564.573
R325 B.n448 B.n252 564.573
R326 B.n76 B.t12 538.062
R327 B.n73 B.t4 538.062
R328 B.n271 B.t15 538.062
R329 B.n277 B.t8 538.062
R330 B.n520 B.n71 256.663
R331 B.n520 B.n70 256.663
R332 B.n520 B.n69 256.663
R333 B.n520 B.n68 256.663
R334 B.n520 B.n67 256.663
R335 B.n520 B.n66 256.663
R336 B.n520 B.n65 256.663
R337 B.n520 B.n64 256.663
R338 B.n520 B.n63 256.663
R339 B.n520 B.n62 256.663
R340 B.n520 B.n61 256.663
R341 B.n520 B.n60 256.663
R342 B.n520 B.n59 256.663
R343 B.n520 B.n58 256.663
R344 B.n520 B.n57 256.663
R345 B.n520 B.n56 256.663
R346 B.n520 B.n55 256.663
R347 B.n520 B.n54 256.663
R348 B.n520 B.n53 256.663
R349 B.n520 B.n52 256.663
R350 B.n520 B.n51 256.663
R351 B.n520 B.n50 256.663
R352 B.n520 B.n49 256.663
R353 B.n520 B.n48 256.663
R354 B.n520 B.n47 256.663
R355 B.n520 B.n46 256.663
R356 B.n520 B.n45 256.663
R357 B.n520 B.n44 256.663
R358 B.n520 B.n43 256.663
R359 B.n520 B.n42 256.663
R360 B.n520 B.n41 256.663
R361 B.n520 B.n40 256.663
R362 B.n520 B.n39 256.663
R363 B.n520 B.n38 256.663
R364 B.n520 B.n37 256.663
R365 B.n520 B.n36 256.663
R366 B.n520 B.n35 256.663
R367 B.n296 B.n253 256.663
R368 B.n302 B.n253 256.663
R369 B.n304 B.n253 256.663
R370 B.n310 B.n253 256.663
R371 B.n312 B.n253 256.663
R372 B.n318 B.n253 256.663
R373 B.n320 B.n253 256.663
R374 B.n326 B.n253 256.663
R375 B.n328 B.n253 256.663
R376 B.n334 B.n253 256.663
R377 B.n336 B.n253 256.663
R378 B.n342 B.n253 256.663
R379 B.n344 B.n253 256.663
R380 B.n350 B.n253 256.663
R381 B.n352 B.n253 256.663
R382 B.n358 B.n253 256.663
R383 B.n360 B.n253 256.663
R384 B.n366 B.n253 256.663
R385 B.n368 B.n253 256.663
R386 B.n374 B.n253 256.663
R387 B.n376 B.n253 256.663
R388 B.n383 B.n253 256.663
R389 B.n385 B.n253 256.663
R390 B.n391 B.n253 256.663
R391 B.n393 B.n253 256.663
R392 B.n399 B.n253 256.663
R393 B.n401 B.n253 256.663
R394 B.n407 B.n253 256.663
R395 B.n409 B.n253 256.663
R396 B.n415 B.n253 256.663
R397 B.n417 B.n253 256.663
R398 B.n423 B.n253 256.663
R399 B.n425 B.n253 256.663
R400 B.n431 B.n253 256.663
R401 B.n433 B.n253 256.663
R402 B.n439 B.n253 256.663
R403 B.n441 B.n253 256.663
R404 B.n557 B.n556 256.663
R405 B.n80 B.n79 163.367
R406 B.n84 B.n83 163.367
R407 B.n88 B.n87 163.367
R408 B.n92 B.n91 163.367
R409 B.n96 B.n95 163.367
R410 B.n100 B.n99 163.367
R411 B.n104 B.n103 163.367
R412 B.n108 B.n107 163.367
R413 B.n112 B.n111 163.367
R414 B.n116 B.n115 163.367
R415 B.n120 B.n119 163.367
R416 B.n124 B.n123 163.367
R417 B.n128 B.n127 163.367
R418 B.n132 B.n131 163.367
R419 B.n136 B.n135 163.367
R420 B.n140 B.n139 163.367
R421 B.n145 B.n144 163.367
R422 B.n149 B.n148 163.367
R423 B.n153 B.n152 163.367
R424 B.n157 B.n156 163.367
R425 B.n161 B.n160 163.367
R426 B.n165 B.n164 163.367
R427 B.n169 B.n168 163.367
R428 B.n173 B.n172 163.367
R429 B.n177 B.n176 163.367
R430 B.n181 B.n180 163.367
R431 B.n185 B.n184 163.367
R432 B.n189 B.n188 163.367
R433 B.n193 B.n192 163.367
R434 B.n197 B.n196 163.367
R435 B.n201 B.n200 163.367
R436 B.n205 B.n204 163.367
R437 B.n209 B.n208 163.367
R438 B.n213 B.n212 163.367
R439 B.n217 B.n216 163.367
R440 B.n221 B.n220 163.367
R441 B.n519 B.n72 163.367
R442 B.n446 B.n248 163.367
R443 B.n454 B.n248 163.367
R444 B.n454 B.n246 163.367
R445 B.n458 B.n246 163.367
R446 B.n458 B.n240 163.367
R447 B.n466 B.n240 163.367
R448 B.n466 B.n238 163.367
R449 B.n470 B.n238 163.367
R450 B.n470 B.n232 163.367
R451 B.n478 B.n232 163.367
R452 B.n478 B.n230 163.367
R453 B.n483 B.n230 163.367
R454 B.n483 B.n225 163.367
R455 B.n492 B.n225 163.367
R456 B.n493 B.n492 163.367
R457 B.n493 B.n5 163.367
R458 B.n6 B.n5 163.367
R459 B.n7 B.n6 163.367
R460 B.n499 B.n7 163.367
R461 B.n500 B.n499 163.367
R462 B.n500 B.n13 163.367
R463 B.n14 B.n13 163.367
R464 B.n15 B.n14 163.367
R465 B.n505 B.n15 163.367
R466 B.n505 B.n20 163.367
R467 B.n21 B.n20 163.367
R468 B.n22 B.n21 163.367
R469 B.n510 B.n22 163.367
R470 B.n510 B.n27 163.367
R471 B.n28 B.n27 163.367
R472 B.n29 B.n28 163.367
R473 B.n515 B.n29 163.367
R474 B.n515 B.n34 163.367
R475 B.n297 B.n295 163.367
R476 B.n301 B.n295 163.367
R477 B.n305 B.n303 163.367
R478 B.n309 B.n293 163.367
R479 B.n313 B.n311 163.367
R480 B.n317 B.n291 163.367
R481 B.n321 B.n319 163.367
R482 B.n325 B.n289 163.367
R483 B.n329 B.n327 163.367
R484 B.n333 B.n287 163.367
R485 B.n337 B.n335 163.367
R486 B.n341 B.n285 163.367
R487 B.n345 B.n343 163.367
R488 B.n349 B.n283 163.367
R489 B.n353 B.n351 163.367
R490 B.n357 B.n281 163.367
R491 B.n361 B.n359 163.367
R492 B.n365 B.n276 163.367
R493 B.n369 B.n367 163.367
R494 B.n373 B.n274 163.367
R495 B.n377 B.n375 163.367
R496 B.n382 B.n270 163.367
R497 B.n386 B.n384 163.367
R498 B.n390 B.n268 163.367
R499 B.n394 B.n392 163.367
R500 B.n398 B.n266 163.367
R501 B.n402 B.n400 163.367
R502 B.n406 B.n264 163.367
R503 B.n410 B.n408 163.367
R504 B.n414 B.n262 163.367
R505 B.n418 B.n416 163.367
R506 B.n422 B.n260 163.367
R507 B.n426 B.n424 163.367
R508 B.n430 B.n258 163.367
R509 B.n434 B.n432 163.367
R510 B.n438 B.n256 163.367
R511 B.n442 B.n440 163.367
R512 B.n448 B.n250 163.367
R513 B.n452 B.n250 163.367
R514 B.n452 B.n244 163.367
R515 B.n460 B.n244 163.367
R516 B.n460 B.n242 163.367
R517 B.n464 B.n242 163.367
R518 B.n464 B.n236 163.367
R519 B.n472 B.n236 163.367
R520 B.n472 B.n234 163.367
R521 B.n476 B.n234 163.367
R522 B.n476 B.n228 163.367
R523 B.n486 B.n228 163.367
R524 B.n486 B.n226 163.367
R525 B.n490 B.n226 163.367
R526 B.n490 B.n3 163.367
R527 B.n555 B.n3 163.367
R528 B.n551 B.n2 163.367
R529 B.n551 B.n550 163.367
R530 B.n550 B.n9 163.367
R531 B.n546 B.n9 163.367
R532 B.n546 B.n11 163.367
R533 B.n542 B.n11 163.367
R534 B.n542 B.n17 163.367
R535 B.n538 B.n17 163.367
R536 B.n538 B.n19 163.367
R537 B.n534 B.n19 163.367
R538 B.n534 B.n24 163.367
R539 B.n530 B.n24 163.367
R540 B.n530 B.n26 163.367
R541 B.n526 B.n26 163.367
R542 B.n526 B.n31 163.367
R543 B.n522 B.n31 163.367
R544 B.n447 B.n253 108.499
R545 B.n521 B.n520 108.499
R546 B.n73 B.t6 90.8277
R547 B.n271 B.t17 90.8277
R548 B.n76 B.t13 90.8169
R549 B.n277 B.t11 90.8169
R550 B.n74 B.t7 71.8216
R551 B.n272 B.t16 71.8216
R552 B.n77 B.t14 71.8108
R553 B.n278 B.t10 71.8108
R554 B.n35 B.n33 71.676
R555 B.n80 B.n36 71.676
R556 B.n84 B.n37 71.676
R557 B.n88 B.n38 71.676
R558 B.n92 B.n39 71.676
R559 B.n96 B.n40 71.676
R560 B.n100 B.n41 71.676
R561 B.n104 B.n42 71.676
R562 B.n108 B.n43 71.676
R563 B.n112 B.n44 71.676
R564 B.n116 B.n45 71.676
R565 B.n120 B.n46 71.676
R566 B.n124 B.n47 71.676
R567 B.n128 B.n48 71.676
R568 B.n132 B.n49 71.676
R569 B.n136 B.n50 71.676
R570 B.n140 B.n51 71.676
R571 B.n145 B.n52 71.676
R572 B.n149 B.n53 71.676
R573 B.n153 B.n54 71.676
R574 B.n157 B.n55 71.676
R575 B.n161 B.n56 71.676
R576 B.n165 B.n57 71.676
R577 B.n169 B.n58 71.676
R578 B.n173 B.n59 71.676
R579 B.n177 B.n60 71.676
R580 B.n181 B.n61 71.676
R581 B.n185 B.n62 71.676
R582 B.n189 B.n63 71.676
R583 B.n193 B.n64 71.676
R584 B.n197 B.n65 71.676
R585 B.n201 B.n66 71.676
R586 B.n205 B.n67 71.676
R587 B.n209 B.n68 71.676
R588 B.n213 B.n69 71.676
R589 B.n217 B.n70 71.676
R590 B.n221 B.n71 71.676
R591 B.n72 B.n71 71.676
R592 B.n220 B.n70 71.676
R593 B.n216 B.n69 71.676
R594 B.n212 B.n68 71.676
R595 B.n208 B.n67 71.676
R596 B.n204 B.n66 71.676
R597 B.n200 B.n65 71.676
R598 B.n196 B.n64 71.676
R599 B.n192 B.n63 71.676
R600 B.n188 B.n62 71.676
R601 B.n184 B.n61 71.676
R602 B.n180 B.n60 71.676
R603 B.n176 B.n59 71.676
R604 B.n172 B.n58 71.676
R605 B.n168 B.n57 71.676
R606 B.n164 B.n56 71.676
R607 B.n160 B.n55 71.676
R608 B.n156 B.n54 71.676
R609 B.n152 B.n53 71.676
R610 B.n148 B.n52 71.676
R611 B.n144 B.n51 71.676
R612 B.n139 B.n50 71.676
R613 B.n135 B.n49 71.676
R614 B.n131 B.n48 71.676
R615 B.n127 B.n47 71.676
R616 B.n123 B.n46 71.676
R617 B.n119 B.n45 71.676
R618 B.n115 B.n44 71.676
R619 B.n111 B.n43 71.676
R620 B.n107 B.n42 71.676
R621 B.n103 B.n41 71.676
R622 B.n99 B.n40 71.676
R623 B.n95 B.n39 71.676
R624 B.n91 B.n38 71.676
R625 B.n87 B.n37 71.676
R626 B.n83 B.n36 71.676
R627 B.n79 B.n35 71.676
R628 B.n296 B.n252 71.676
R629 B.n302 B.n301 71.676
R630 B.n305 B.n304 71.676
R631 B.n310 B.n309 71.676
R632 B.n313 B.n312 71.676
R633 B.n318 B.n317 71.676
R634 B.n321 B.n320 71.676
R635 B.n326 B.n325 71.676
R636 B.n329 B.n328 71.676
R637 B.n334 B.n333 71.676
R638 B.n337 B.n336 71.676
R639 B.n342 B.n341 71.676
R640 B.n345 B.n344 71.676
R641 B.n350 B.n349 71.676
R642 B.n353 B.n352 71.676
R643 B.n358 B.n357 71.676
R644 B.n361 B.n360 71.676
R645 B.n366 B.n365 71.676
R646 B.n369 B.n368 71.676
R647 B.n374 B.n373 71.676
R648 B.n377 B.n376 71.676
R649 B.n383 B.n382 71.676
R650 B.n386 B.n385 71.676
R651 B.n391 B.n390 71.676
R652 B.n394 B.n393 71.676
R653 B.n399 B.n398 71.676
R654 B.n402 B.n401 71.676
R655 B.n407 B.n406 71.676
R656 B.n410 B.n409 71.676
R657 B.n415 B.n414 71.676
R658 B.n418 B.n417 71.676
R659 B.n423 B.n422 71.676
R660 B.n426 B.n425 71.676
R661 B.n431 B.n430 71.676
R662 B.n434 B.n433 71.676
R663 B.n439 B.n438 71.676
R664 B.n442 B.n441 71.676
R665 B.n297 B.n296 71.676
R666 B.n303 B.n302 71.676
R667 B.n304 B.n293 71.676
R668 B.n311 B.n310 71.676
R669 B.n312 B.n291 71.676
R670 B.n319 B.n318 71.676
R671 B.n320 B.n289 71.676
R672 B.n327 B.n326 71.676
R673 B.n328 B.n287 71.676
R674 B.n335 B.n334 71.676
R675 B.n336 B.n285 71.676
R676 B.n343 B.n342 71.676
R677 B.n344 B.n283 71.676
R678 B.n351 B.n350 71.676
R679 B.n352 B.n281 71.676
R680 B.n359 B.n358 71.676
R681 B.n360 B.n276 71.676
R682 B.n367 B.n366 71.676
R683 B.n368 B.n274 71.676
R684 B.n375 B.n374 71.676
R685 B.n376 B.n270 71.676
R686 B.n384 B.n383 71.676
R687 B.n385 B.n268 71.676
R688 B.n392 B.n391 71.676
R689 B.n393 B.n266 71.676
R690 B.n400 B.n399 71.676
R691 B.n401 B.n264 71.676
R692 B.n408 B.n407 71.676
R693 B.n409 B.n262 71.676
R694 B.n416 B.n415 71.676
R695 B.n417 B.n260 71.676
R696 B.n424 B.n423 71.676
R697 B.n425 B.n258 71.676
R698 B.n432 B.n431 71.676
R699 B.n433 B.n256 71.676
R700 B.n440 B.n439 71.676
R701 B.n441 B.n254 71.676
R702 B.n556 B.n555 71.676
R703 B.n556 B.n2 71.676
R704 B.n142 B.n77 59.5399
R705 B.n75 B.n74 59.5399
R706 B.n379 B.n272 59.5399
R707 B.n279 B.n278 59.5399
R708 B.n447 B.n249 52.3265
R709 B.n453 B.n249 52.3265
R710 B.n453 B.n245 52.3265
R711 B.n459 B.n245 52.3265
R712 B.n465 B.n241 52.3265
R713 B.n465 B.n237 52.3265
R714 B.n471 B.n237 52.3265
R715 B.n471 B.n233 52.3265
R716 B.n477 B.n233 52.3265
R717 B.n485 B.n229 52.3265
R718 B.n485 B.n484 52.3265
R719 B.n491 B.n4 52.3265
R720 B.n554 B.n4 52.3265
R721 B.n554 B.n553 52.3265
R722 B.n553 B.n552 52.3265
R723 B.n552 B.n8 52.3265
R724 B.n545 B.n12 52.3265
R725 B.n545 B.n544 52.3265
R726 B.n543 B.n16 52.3265
R727 B.n537 B.n16 52.3265
R728 B.n537 B.n536 52.3265
R729 B.n536 B.n535 52.3265
R730 B.n535 B.n23 52.3265
R731 B.n529 B.n528 52.3265
R732 B.n528 B.n527 52.3265
R733 B.n527 B.n30 52.3265
R734 B.n521 B.n30 52.3265
R735 B.n449 B.n251 36.6834
R736 B.n445 B.n444 36.6834
R737 B.n518 B.n517 36.6834
R738 B.n523 B.n32 36.6834
R739 B.n477 B.t1 30.011
R740 B.t0 B.n543 30.011
R741 B.n491 B.t3 28.472
R742 B.t2 B.n8 28.472
R743 B.t9 B.n241 26.933
R744 B.t5 B.n23 26.933
R745 B.n459 B.t9 25.394
R746 B.n529 B.t5 25.394
R747 B.n484 B.t3 23.855
R748 B.n12 B.t2 23.855
R749 B.t1 B.n229 22.316
R750 B.n544 B.t0 22.316
R751 B.n77 B.n76 19.0066
R752 B.n74 B.n73 19.0066
R753 B.n272 B.n271 19.0066
R754 B.n278 B.n277 19.0066
R755 B B.n557 18.0485
R756 B.n450 B.n449 10.6151
R757 B.n451 B.n450 10.6151
R758 B.n451 B.n243 10.6151
R759 B.n461 B.n243 10.6151
R760 B.n462 B.n461 10.6151
R761 B.n463 B.n462 10.6151
R762 B.n463 B.n235 10.6151
R763 B.n473 B.n235 10.6151
R764 B.n474 B.n473 10.6151
R765 B.n475 B.n474 10.6151
R766 B.n475 B.n227 10.6151
R767 B.n487 B.n227 10.6151
R768 B.n488 B.n487 10.6151
R769 B.n489 B.n488 10.6151
R770 B.n489 B.n0 10.6151
R771 B.n298 B.n251 10.6151
R772 B.n299 B.n298 10.6151
R773 B.n300 B.n299 10.6151
R774 B.n300 B.n294 10.6151
R775 B.n306 B.n294 10.6151
R776 B.n307 B.n306 10.6151
R777 B.n308 B.n307 10.6151
R778 B.n308 B.n292 10.6151
R779 B.n314 B.n292 10.6151
R780 B.n315 B.n314 10.6151
R781 B.n316 B.n315 10.6151
R782 B.n316 B.n290 10.6151
R783 B.n322 B.n290 10.6151
R784 B.n323 B.n322 10.6151
R785 B.n324 B.n323 10.6151
R786 B.n324 B.n288 10.6151
R787 B.n330 B.n288 10.6151
R788 B.n331 B.n330 10.6151
R789 B.n332 B.n331 10.6151
R790 B.n332 B.n286 10.6151
R791 B.n338 B.n286 10.6151
R792 B.n339 B.n338 10.6151
R793 B.n340 B.n339 10.6151
R794 B.n340 B.n284 10.6151
R795 B.n346 B.n284 10.6151
R796 B.n347 B.n346 10.6151
R797 B.n348 B.n347 10.6151
R798 B.n348 B.n282 10.6151
R799 B.n354 B.n282 10.6151
R800 B.n355 B.n354 10.6151
R801 B.n356 B.n355 10.6151
R802 B.n356 B.n280 10.6151
R803 B.n363 B.n362 10.6151
R804 B.n364 B.n363 10.6151
R805 B.n364 B.n275 10.6151
R806 B.n370 B.n275 10.6151
R807 B.n371 B.n370 10.6151
R808 B.n372 B.n371 10.6151
R809 B.n372 B.n273 10.6151
R810 B.n378 B.n273 10.6151
R811 B.n381 B.n380 10.6151
R812 B.n381 B.n269 10.6151
R813 B.n387 B.n269 10.6151
R814 B.n388 B.n387 10.6151
R815 B.n389 B.n388 10.6151
R816 B.n389 B.n267 10.6151
R817 B.n395 B.n267 10.6151
R818 B.n396 B.n395 10.6151
R819 B.n397 B.n396 10.6151
R820 B.n397 B.n265 10.6151
R821 B.n403 B.n265 10.6151
R822 B.n404 B.n403 10.6151
R823 B.n405 B.n404 10.6151
R824 B.n405 B.n263 10.6151
R825 B.n411 B.n263 10.6151
R826 B.n412 B.n411 10.6151
R827 B.n413 B.n412 10.6151
R828 B.n413 B.n261 10.6151
R829 B.n419 B.n261 10.6151
R830 B.n420 B.n419 10.6151
R831 B.n421 B.n420 10.6151
R832 B.n421 B.n259 10.6151
R833 B.n427 B.n259 10.6151
R834 B.n428 B.n427 10.6151
R835 B.n429 B.n428 10.6151
R836 B.n429 B.n257 10.6151
R837 B.n435 B.n257 10.6151
R838 B.n436 B.n435 10.6151
R839 B.n437 B.n436 10.6151
R840 B.n437 B.n255 10.6151
R841 B.n443 B.n255 10.6151
R842 B.n444 B.n443 10.6151
R843 B.n445 B.n247 10.6151
R844 B.n455 B.n247 10.6151
R845 B.n456 B.n455 10.6151
R846 B.n457 B.n456 10.6151
R847 B.n457 B.n239 10.6151
R848 B.n467 B.n239 10.6151
R849 B.n468 B.n467 10.6151
R850 B.n469 B.n468 10.6151
R851 B.n469 B.n231 10.6151
R852 B.n479 B.n231 10.6151
R853 B.n480 B.n479 10.6151
R854 B.n482 B.n480 10.6151
R855 B.n482 B.n481 10.6151
R856 B.n481 B.n224 10.6151
R857 B.n494 B.n224 10.6151
R858 B.n495 B.n494 10.6151
R859 B.n496 B.n495 10.6151
R860 B.n497 B.n496 10.6151
R861 B.n498 B.n497 10.6151
R862 B.n501 B.n498 10.6151
R863 B.n502 B.n501 10.6151
R864 B.n503 B.n502 10.6151
R865 B.n504 B.n503 10.6151
R866 B.n506 B.n504 10.6151
R867 B.n507 B.n506 10.6151
R868 B.n508 B.n507 10.6151
R869 B.n509 B.n508 10.6151
R870 B.n511 B.n509 10.6151
R871 B.n512 B.n511 10.6151
R872 B.n513 B.n512 10.6151
R873 B.n514 B.n513 10.6151
R874 B.n516 B.n514 10.6151
R875 B.n517 B.n516 10.6151
R876 B.n549 B.n1 10.6151
R877 B.n549 B.n548 10.6151
R878 B.n548 B.n547 10.6151
R879 B.n547 B.n10 10.6151
R880 B.n541 B.n10 10.6151
R881 B.n541 B.n540 10.6151
R882 B.n540 B.n539 10.6151
R883 B.n539 B.n18 10.6151
R884 B.n533 B.n18 10.6151
R885 B.n533 B.n532 10.6151
R886 B.n532 B.n531 10.6151
R887 B.n531 B.n25 10.6151
R888 B.n525 B.n25 10.6151
R889 B.n525 B.n524 10.6151
R890 B.n524 B.n523 10.6151
R891 B.n78 B.n32 10.6151
R892 B.n81 B.n78 10.6151
R893 B.n82 B.n81 10.6151
R894 B.n85 B.n82 10.6151
R895 B.n86 B.n85 10.6151
R896 B.n89 B.n86 10.6151
R897 B.n90 B.n89 10.6151
R898 B.n93 B.n90 10.6151
R899 B.n94 B.n93 10.6151
R900 B.n97 B.n94 10.6151
R901 B.n98 B.n97 10.6151
R902 B.n101 B.n98 10.6151
R903 B.n102 B.n101 10.6151
R904 B.n105 B.n102 10.6151
R905 B.n106 B.n105 10.6151
R906 B.n109 B.n106 10.6151
R907 B.n110 B.n109 10.6151
R908 B.n113 B.n110 10.6151
R909 B.n114 B.n113 10.6151
R910 B.n117 B.n114 10.6151
R911 B.n118 B.n117 10.6151
R912 B.n121 B.n118 10.6151
R913 B.n122 B.n121 10.6151
R914 B.n125 B.n122 10.6151
R915 B.n126 B.n125 10.6151
R916 B.n129 B.n126 10.6151
R917 B.n130 B.n129 10.6151
R918 B.n133 B.n130 10.6151
R919 B.n134 B.n133 10.6151
R920 B.n137 B.n134 10.6151
R921 B.n138 B.n137 10.6151
R922 B.n141 B.n138 10.6151
R923 B.n146 B.n143 10.6151
R924 B.n147 B.n146 10.6151
R925 B.n150 B.n147 10.6151
R926 B.n151 B.n150 10.6151
R927 B.n154 B.n151 10.6151
R928 B.n155 B.n154 10.6151
R929 B.n158 B.n155 10.6151
R930 B.n159 B.n158 10.6151
R931 B.n163 B.n162 10.6151
R932 B.n166 B.n163 10.6151
R933 B.n167 B.n166 10.6151
R934 B.n170 B.n167 10.6151
R935 B.n171 B.n170 10.6151
R936 B.n174 B.n171 10.6151
R937 B.n175 B.n174 10.6151
R938 B.n178 B.n175 10.6151
R939 B.n179 B.n178 10.6151
R940 B.n182 B.n179 10.6151
R941 B.n183 B.n182 10.6151
R942 B.n186 B.n183 10.6151
R943 B.n187 B.n186 10.6151
R944 B.n190 B.n187 10.6151
R945 B.n191 B.n190 10.6151
R946 B.n194 B.n191 10.6151
R947 B.n195 B.n194 10.6151
R948 B.n198 B.n195 10.6151
R949 B.n199 B.n198 10.6151
R950 B.n202 B.n199 10.6151
R951 B.n203 B.n202 10.6151
R952 B.n206 B.n203 10.6151
R953 B.n207 B.n206 10.6151
R954 B.n210 B.n207 10.6151
R955 B.n211 B.n210 10.6151
R956 B.n214 B.n211 10.6151
R957 B.n215 B.n214 10.6151
R958 B.n218 B.n215 10.6151
R959 B.n219 B.n218 10.6151
R960 B.n222 B.n219 10.6151
R961 B.n223 B.n222 10.6151
R962 B.n518 B.n223 10.6151
R963 B.n557 B.n0 8.11757
R964 B.n557 B.n1 8.11757
R965 B.n362 B.n279 6.5566
R966 B.n379 B.n378 6.5566
R967 B.n143 B.n142 6.5566
R968 B.n159 B.n75 6.5566
R969 B.n280 B.n279 4.05904
R970 B.n380 B.n379 4.05904
R971 B.n142 B.n141 4.05904
R972 B.n162 B.n75 4.05904
R973 VN.n0 VN.t1 415.865
R974 VN.n1 VN.t2 415.865
R975 VN.n0 VN.t3 415.817
R976 VN.n1 VN.t0 415.817
R977 VN VN.n1 83.0049
R978 VN VN.n0 44.7132
R979 VDD2.n2 VDD2.n0 99.9504
R980 VDD2.n2 VDD2.n1 65.9253
R981 VDD2.n1 VDD2.t3 2.19562
R982 VDD2.n1 VDD2.t1 2.19562
R983 VDD2.n0 VDD2.t2 2.19562
R984 VDD2.n0 VDD2.t0 2.19562
R985 VDD2 VDD2.n2 0.0586897
C0 VTAIL VDD1 5.59947f
C1 VDD2 VN 2.36834f
C2 VP VDD1 2.49109f
C3 VP VTAIL 2.09349f
C4 VDD2 VDD1 0.555011f
C5 VDD2 VTAIL 5.6406f
C6 VP VDD2 0.270363f
C7 VDD1 VN 0.147377f
C8 VTAIL VN 2.07938f
C9 VP VN 4.23527f
C10 VDD2 B 2.437639f
C11 VDD1 B 5.76593f
C12 VTAIL B 7.054526f
C13 VN B 7.64907f
C14 VP B 4.592678f
C15 VDD2.t2 B 0.201762f
C16 VDD2.t0 B 0.201762f
C17 VDD2.n0 B 2.24855f
C18 VDD2.t3 B 0.201762f
C19 VDD2.t1 B 0.201762f
C20 VDD2.n1 B 1.76533f
C21 VDD2.n2 B 3.09592f
C22 VN.t1 B 0.870975f
C23 VN.t3 B 0.870924f
C24 VN.n0 B 0.685264f
C25 VN.t2 B 0.870975f
C26 VN.t0 B 0.870924f
C27 VN.n1 B 1.56129f
C28 VDD1.t0 B 0.201648f
C29 VDD1.t2 B 0.201648f
C30 VDD1.n0 B 1.76462f
C31 VDD1.t1 B 0.201648f
C32 VDD1.t3 B 0.201648f
C33 VDD1.n1 B 2.27205f
C34 VTAIL.t2 B 1.30068f
C35 VTAIL.n0 B 0.263668f
C36 VTAIL.t4 B 1.30068f
C37 VTAIL.n1 B 0.283731f
C38 VTAIL.t7 B 1.30068f
C39 VTAIL.n2 B 0.964917f
C40 VTAIL.t1 B 1.30068f
C41 VTAIL.n3 B 0.964914f
C42 VTAIL.t3 B 1.30068f
C43 VTAIL.n4 B 0.283728f
C44 VTAIL.t5 B 1.30068f
C45 VTAIL.n5 B 0.283728f
C46 VTAIL.t6 B 1.30068f
C47 VTAIL.n6 B 0.964917f
C48 VTAIL.t0 B 1.30068f
C49 VTAIL.n7 B 0.938444f
C50 VP.n0 B 0.051733f
C51 VP.t1 B 0.888215f
C52 VP.t3 B 0.888266f
C53 VP.n1 B 1.57179f
C54 VP.n2 B 2.86928f
C55 VP.t2 B 0.869804f
C56 VP.n3 B 0.361749f
C57 VP.n4 B 0.011739f
C58 VP.t0 B 0.869804f
C59 VP.n5 B 0.361749f
C60 VP.n6 B 0.040091f
.ends

