* NGSPICE file created from diff_pair_sample_0009.ext - technology: sky130A

.subckt diff_pair_sample_0009 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t12 VN.t0 VDD2.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=1.73745 pd=10.86 as=1.73745 ps=10.86 w=10.53 l=0.42
X1 VDD2.t2 VN.t1 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=1.73745 pd=10.86 as=1.73745 ps=10.86 w=10.53 l=0.42
X2 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=4.1067 pd=21.84 as=0 ps=0 w=10.53 l=0.42
X3 VTAIL.t10 VN.t2 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.73745 pd=10.86 as=1.73745 ps=10.86 w=10.53 l=0.42
X4 VTAIL.t9 VN.t3 VDD2.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=4.1067 pd=21.84 as=1.73745 ps=10.86 w=10.53 l=0.42
X5 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=4.1067 pd=21.84 as=0 ps=0 w=10.53 l=0.42
X6 VTAIL.t3 VP.t0 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=4.1067 pd=21.84 as=1.73745 ps=10.86 w=10.53 l=0.42
X7 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.1067 pd=21.84 as=0 ps=0 w=10.53 l=0.42
X8 VTAIL.t8 VN.t4 VDD2.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=4.1067 pd=21.84 as=1.73745 ps=10.86 w=10.53 l=0.42
X9 VTAIL.t14 VP.t1 VDD1.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=4.1067 pd=21.84 as=1.73745 ps=10.86 w=10.53 l=0.42
X10 VTAIL.t4 VP.t2 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=1.73745 pd=10.86 as=1.73745 ps=10.86 w=10.53 l=0.42
X11 VTAIL.t13 VP.t3 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=1.73745 pd=10.86 as=1.73745 ps=10.86 w=10.53 l=0.42
X12 VDD1.t3 VP.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.73745 pd=10.86 as=1.73745 ps=10.86 w=10.53 l=0.42
X13 VDD2.t0 VN.t5 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=1.73745 pd=10.86 as=4.1067 ps=21.84 w=10.53 l=0.42
X14 VDD2.t1 VN.t6 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=1.73745 pd=10.86 as=1.73745 ps=10.86 w=10.53 l=0.42
X15 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.1067 pd=21.84 as=0 ps=0 w=10.53 l=0.42
X16 VDD2.t5 VN.t7 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.73745 pd=10.86 as=4.1067 ps=21.84 w=10.53 l=0.42
X17 VDD1.t2 VP.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.73745 pd=10.86 as=1.73745 ps=10.86 w=10.53 l=0.42
X18 VDD1.t1 VP.t6 VTAIL.t15 B.t5 sky130_fd_pr__nfet_01v8 ad=1.73745 pd=10.86 as=4.1067 ps=21.84 w=10.53 l=0.42
X19 VDD1.t0 VP.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.73745 pd=10.86 as=4.1067 ps=21.84 w=10.53 l=0.42
R0 VN.n2 VN.t4 719.308
R1 VN.n10 VN.t5 719.308
R2 VN.n1 VN.t1 698.327
R3 VN.n5 VN.t2 698.327
R4 VN.n6 VN.t7 698.327
R5 VN.n9 VN.t0 698.327
R6 VN.n13 VN.t6 698.327
R7 VN.n14 VN.t3 698.327
R8 VN.n7 VN.n6 161.3
R9 VN.n15 VN.n14 161.3
R10 VN.n13 VN.n8 161.3
R11 VN.n12 VN.n11 161.3
R12 VN.n5 VN.n0 161.3
R13 VN.n4 VN.n3 161.3
R14 VN.n11 VN.n10 70.4033
R15 VN.n3 VN.n2 70.4033
R16 VN.n6 VN.n5 48.2005
R17 VN.n14 VN.n13 48.2005
R18 VN VN.n15 39.9418
R19 VN.n4 VN.n1 24.1005
R20 VN.n5 VN.n4 24.1005
R21 VN.n13 VN.n12 24.1005
R22 VN.n12 VN.n9 24.1005
R23 VN.n10 VN.n9 20.9576
R24 VN.n2 VN.n1 20.9576
R25 VN.n15 VN.n8 0.189894
R26 VN.n11 VN.n8 0.189894
R27 VN.n3 VN.n0 0.189894
R28 VN.n7 VN.n0 0.189894
R29 VN VN.n7 0.0516364
R30 VDD2.n2 VDD2.n1 66.8234
R31 VDD2.n2 VDD2.n0 66.8234
R32 VDD2 VDD2.n5 66.8206
R33 VDD2.n4 VDD2.n3 66.5557
R34 VDD2.n4 VDD2.n2 35.7024
R35 VDD2.n5 VDD2.t3 1.88084
R36 VDD2.n5 VDD2.t0 1.88084
R37 VDD2.n3 VDD2.t7 1.88084
R38 VDD2.n3 VDD2.t1 1.88084
R39 VDD2.n1 VDD2.t4 1.88084
R40 VDD2.n1 VDD2.t5 1.88084
R41 VDD2.n0 VDD2.t6 1.88084
R42 VDD2.n0 VDD2.t2 1.88084
R43 VDD2 VDD2.n4 0.381966
R44 VTAIL.n11 VTAIL.t14 51.7573
R45 VTAIL.n10 VTAIL.t7 51.7573
R46 VTAIL.n7 VTAIL.t9 51.7573
R47 VTAIL.n14 VTAIL.t0 51.757
R48 VTAIL.n15 VTAIL.t5 51.757
R49 VTAIL.n2 VTAIL.t8 51.757
R50 VTAIL.n3 VTAIL.t15 51.757
R51 VTAIL.n6 VTAIL.t3 51.757
R52 VTAIL.n13 VTAIL.n12 49.8769
R53 VTAIL.n9 VTAIL.n8 49.8769
R54 VTAIL.n1 VTAIL.n0 49.8767
R55 VTAIL.n5 VTAIL.n4 49.8767
R56 VTAIL.n15 VTAIL.n14 22.091
R57 VTAIL.n7 VTAIL.n6 22.091
R58 VTAIL.n0 VTAIL.t11 1.88084
R59 VTAIL.n0 VTAIL.t10 1.88084
R60 VTAIL.n4 VTAIL.t1 1.88084
R61 VTAIL.n4 VTAIL.t13 1.88084
R62 VTAIL.n12 VTAIL.t2 1.88084
R63 VTAIL.n12 VTAIL.t4 1.88084
R64 VTAIL.n8 VTAIL.t6 1.88084
R65 VTAIL.n8 VTAIL.t12 1.88084
R66 VTAIL.n9 VTAIL.n7 0.647052
R67 VTAIL.n10 VTAIL.n9 0.647052
R68 VTAIL.n13 VTAIL.n11 0.647052
R69 VTAIL.n14 VTAIL.n13 0.647052
R70 VTAIL.n6 VTAIL.n5 0.647052
R71 VTAIL.n5 VTAIL.n3 0.647052
R72 VTAIL.n2 VTAIL.n1 0.647052
R73 VTAIL VTAIL.n15 0.588862
R74 VTAIL.n11 VTAIL.n10 0.470328
R75 VTAIL.n3 VTAIL.n2 0.470328
R76 VTAIL VTAIL.n1 0.0586897
R77 B.n330 B.t16 812.924
R78 B.n327 B.t12 812.924
R79 B.n84 B.t19 812.924
R80 B.n82 B.t8 812.924
R81 B.n582 B.n581 585
R82 B.n248 B.n80 585
R83 B.n247 B.n246 585
R84 B.n245 B.n244 585
R85 B.n243 B.n242 585
R86 B.n241 B.n240 585
R87 B.n239 B.n238 585
R88 B.n237 B.n236 585
R89 B.n235 B.n234 585
R90 B.n233 B.n232 585
R91 B.n231 B.n230 585
R92 B.n229 B.n228 585
R93 B.n227 B.n226 585
R94 B.n225 B.n224 585
R95 B.n223 B.n222 585
R96 B.n221 B.n220 585
R97 B.n219 B.n218 585
R98 B.n217 B.n216 585
R99 B.n215 B.n214 585
R100 B.n213 B.n212 585
R101 B.n211 B.n210 585
R102 B.n209 B.n208 585
R103 B.n207 B.n206 585
R104 B.n205 B.n204 585
R105 B.n203 B.n202 585
R106 B.n201 B.n200 585
R107 B.n199 B.n198 585
R108 B.n197 B.n196 585
R109 B.n195 B.n194 585
R110 B.n193 B.n192 585
R111 B.n191 B.n190 585
R112 B.n189 B.n188 585
R113 B.n187 B.n186 585
R114 B.n185 B.n184 585
R115 B.n183 B.n182 585
R116 B.n181 B.n180 585
R117 B.n179 B.n178 585
R118 B.n176 B.n175 585
R119 B.n174 B.n173 585
R120 B.n172 B.n171 585
R121 B.n170 B.n169 585
R122 B.n168 B.n167 585
R123 B.n166 B.n165 585
R124 B.n164 B.n163 585
R125 B.n162 B.n161 585
R126 B.n160 B.n159 585
R127 B.n158 B.n157 585
R128 B.n155 B.n154 585
R129 B.n153 B.n152 585
R130 B.n151 B.n150 585
R131 B.n149 B.n148 585
R132 B.n147 B.n146 585
R133 B.n145 B.n144 585
R134 B.n143 B.n142 585
R135 B.n141 B.n140 585
R136 B.n139 B.n138 585
R137 B.n137 B.n136 585
R138 B.n135 B.n134 585
R139 B.n133 B.n132 585
R140 B.n131 B.n130 585
R141 B.n129 B.n128 585
R142 B.n127 B.n126 585
R143 B.n125 B.n124 585
R144 B.n123 B.n122 585
R145 B.n121 B.n120 585
R146 B.n119 B.n118 585
R147 B.n117 B.n116 585
R148 B.n115 B.n114 585
R149 B.n113 B.n112 585
R150 B.n111 B.n110 585
R151 B.n109 B.n108 585
R152 B.n107 B.n106 585
R153 B.n105 B.n104 585
R154 B.n103 B.n102 585
R155 B.n101 B.n100 585
R156 B.n99 B.n98 585
R157 B.n97 B.n96 585
R158 B.n95 B.n94 585
R159 B.n93 B.n92 585
R160 B.n91 B.n90 585
R161 B.n89 B.n88 585
R162 B.n87 B.n86 585
R163 B.n39 B.n38 585
R164 B.n587 B.n586 585
R165 B.n580 B.n81 585
R166 B.n81 B.n36 585
R167 B.n579 B.n35 585
R168 B.n591 B.n35 585
R169 B.n578 B.n34 585
R170 B.n592 B.n34 585
R171 B.n577 B.n33 585
R172 B.n593 B.n33 585
R173 B.n576 B.n575 585
R174 B.n575 B.n32 585
R175 B.n574 B.n28 585
R176 B.n599 B.n28 585
R177 B.n573 B.n27 585
R178 B.n600 B.n27 585
R179 B.n572 B.n26 585
R180 B.n601 B.n26 585
R181 B.n571 B.n570 585
R182 B.n570 B.n22 585
R183 B.n569 B.n21 585
R184 B.n607 B.n21 585
R185 B.n568 B.n20 585
R186 B.n608 B.n20 585
R187 B.n567 B.n19 585
R188 B.n609 B.n19 585
R189 B.n566 B.n565 585
R190 B.n565 B.n15 585
R191 B.n564 B.n14 585
R192 B.n615 B.n14 585
R193 B.n563 B.n13 585
R194 B.n616 B.n13 585
R195 B.n562 B.n12 585
R196 B.n617 B.n12 585
R197 B.n561 B.n560 585
R198 B.n560 B.n11 585
R199 B.n559 B.n7 585
R200 B.n623 B.n7 585
R201 B.n558 B.n6 585
R202 B.n624 B.n6 585
R203 B.n557 B.n5 585
R204 B.n625 B.n5 585
R205 B.n556 B.n555 585
R206 B.n555 B.n4 585
R207 B.n554 B.n249 585
R208 B.n554 B.n553 585
R209 B.n543 B.n250 585
R210 B.n546 B.n250 585
R211 B.n545 B.n544 585
R212 B.n547 B.n545 585
R213 B.n542 B.n254 585
R214 B.n258 B.n254 585
R215 B.n541 B.n540 585
R216 B.n540 B.n539 585
R217 B.n256 B.n255 585
R218 B.n257 B.n256 585
R219 B.n532 B.n531 585
R220 B.n533 B.n532 585
R221 B.n530 B.n263 585
R222 B.n263 B.n262 585
R223 B.n529 B.n528 585
R224 B.n528 B.n527 585
R225 B.n265 B.n264 585
R226 B.n266 B.n265 585
R227 B.n520 B.n519 585
R228 B.n521 B.n520 585
R229 B.n518 B.n271 585
R230 B.n271 B.n270 585
R231 B.n517 B.n516 585
R232 B.n516 B.n515 585
R233 B.n273 B.n272 585
R234 B.n508 B.n273 585
R235 B.n507 B.n506 585
R236 B.n509 B.n507 585
R237 B.n505 B.n278 585
R238 B.n278 B.n277 585
R239 B.n504 B.n503 585
R240 B.n503 B.n502 585
R241 B.n280 B.n279 585
R242 B.n281 B.n280 585
R243 B.n498 B.n497 585
R244 B.n284 B.n283 585
R245 B.n494 B.n493 585
R246 B.n495 B.n494 585
R247 B.n492 B.n326 585
R248 B.n491 B.n490 585
R249 B.n489 B.n488 585
R250 B.n487 B.n486 585
R251 B.n485 B.n484 585
R252 B.n483 B.n482 585
R253 B.n481 B.n480 585
R254 B.n479 B.n478 585
R255 B.n477 B.n476 585
R256 B.n475 B.n474 585
R257 B.n473 B.n472 585
R258 B.n471 B.n470 585
R259 B.n469 B.n468 585
R260 B.n467 B.n466 585
R261 B.n465 B.n464 585
R262 B.n463 B.n462 585
R263 B.n461 B.n460 585
R264 B.n459 B.n458 585
R265 B.n457 B.n456 585
R266 B.n455 B.n454 585
R267 B.n453 B.n452 585
R268 B.n451 B.n450 585
R269 B.n449 B.n448 585
R270 B.n447 B.n446 585
R271 B.n445 B.n444 585
R272 B.n443 B.n442 585
R273 B.n441 B.n440 585
R274 B.n439 B.n438 585
R275 B.n437 B.n436 585
R276 B.n435 B.n434 585
R277 B.n433 B.n432 585
R278 B.n431 B.n430 585
R279 B.n429 B.n428 585
R280 B.n427 B.n426 585
R281 B.n425 B.n424 585
R282 B.n423 B.n422 585
R283 B.n421 B.n420 585
R284 B.n419 B.n418 585
R285 B.n417 B.n416 585
R286 B.n415 B.n414 585
R287 B.n413 B.n412 585
R288 B.n411 B.n410 585
R289 B.n409 B.n408 585
R290 B.n407 B.n406 585
R291 B.n405 B.n404 585
R292 B.n403 B.n402 585
R293 B.n401 B.n400 585
R294 B.n399 B.n398 585
R295 B.n397 B.n396 585
R296 B.n395 B.n394 585
R297 B.n393 B.n392 585
R298 B.n391 B.n390 585
R299 B.n389 B.n388 585
R300 B.n387 B.n386 585
R301 B.n385 B.n384 585
R302 B.n383 B.n382 585
R303 B.n381 B.n380 585
R304 B.n379 B.n378 585
R305 B.n377 B.n376 585
R306 B.n375 B.n374 585
R307 B.n373 B.n372 585
R308 B.n371 B.n370 585
R309 B.n369 B.n368 585
R310 B.n367 B.n366 585
R311 B.n365 B.n364 585
R312 B.n363 B.n362 585
R313 B.n361 B.n360 585
R314 B.n359 B.n358 585
R315 B.n357 B.n356 585
R316 B.n355 B.n354 585
R317 B.n353 B.n352 585
R318 B.n351 B.n350 585
R319 B.n349 B.n348 585
R320 B.n347 B.n346 585
R321 B.n345 B.n344 585
R322 B.n343 B.n342 585
R323 B.n341 B.n340 585
R324 B.n339 B.n338 585
R325 B.n337 B.n336 585
R326 B.n335 B.n334 585
R327 B.n333 B.n325 585
R328 B.n495 B.n325 585
R329 B.n499 B.n282 585
R330 B.n282 B.n281 585
R331 B.n501 B.n500 585
R332 B.n502 B.n501 585
R333 B.n276 B.n275 585
R334 B.n277 B.n276 585
R335 B.n511 B.n510 585
R336 B.n510 B.n509 585
R337 B.n512 B.n274 585
R338 B.n508 B.n274 585
R339 B.n514 B.n513 585
R340 B.n515 B.n514 585
R341 B.n269 B.n268 585
R342 B.n270 B.n269 585
R343 B.n523 B.n522 585
R344 B.n522 B.n521 585
R345 B.n524 B.n267 585
R346 B.n267 B.n266 585
R347 B.n526 B.n525 585
R348 B.n527 B.n526 585
R349 B.n261 B.n260 585
R350 B.n262 B.n261 585
R351 B.n535 B.n534 585
R352 B.n534 B.n533 585
R353 B.n536 B.n259 585
R354 B.n259 B.n257 585
R355 B.n538 B.n537 585
R356 B.n539 B.n538 585
R357 B.n253 B.n252 585
R358 B.n258 B.n253 585
R359 B.n549 B.n548 585
R360 B.n548 B.n547 585
R361 B.n550 B.n251 585
R362 B.n546 B.n251 585
R363 B.n552 B.n551 585
R364 B.n553 B.n552 585
R365 B.n2 B.n0 585
R366 B.n4 B.n2 585
R367 B.n3 B.n1 585
R368 B.n624 B.n3 585
R369 B.n622 B.n621 585
R370 B.n623 B.n622 585
R371 B.n620 B.n8 585
R372 B.n11 B.n8 585
R373 B.n619 B.n618 585
R374 B.n618 B.n617 585
R375 B.n10 B.n9 585
R376 B.n616 B.n10 585
R377 B.n614 B.n613 585
R378 B.n615 B.n614 585
R379 B.n612 B.n16 585
R380 B.n16 B.n15 585
R381 B.n611 B.n610 585
R382 B.n610 B.n609 585
R383 B.n18 B.n17 585
R384 B.n608 B.n18 585
R385 B.n606 B.n605 585
R386 B.n607 B.n606 585
R387 B.n604 B.n23 585
R388 B.n23 B.n22 585
R389 B.n603 B.n602 585
R390 B.n602 B.n601 585
R391 B.n25 B.n24 585
R392 B.n600 B.n25 585
R393 B.n598 B.n597 585
R394 B.n599 B.n598 585
R395 B.n596 B.n29 585
R396 B.n32 B.n29 585
R397 B.n595 B.n594 585
R398 B.n594 B.n593 585
R399 B.n31 B.n30 585
R400 B.n592 B.n31 585
R401 B.n590 B.n589 585
R402 B.n591 B.n590 585
R403 B.n588 B.n37 585
R404 B.n37 B.n36 585
R405 B.n627 B.n626 585
R406 B.n626 B.n625 585
R407 B.n497 B.n282 535.745
R408 B.n586 B.n37 535.745
R409 B.n325 B.n280 535.745
R410 B.n582 B.n81 535.745
R411 B.n584 B.n583 256.663
R412 B.n584 B.n79 256.663
R413 B.n584 B.n78 256.663
R414 B.n584 B.n77 256.663
R415 B.n584 B.n76 256.663
R416 B.n584 B.n75 256.663
R417 B.n584 B.n74 256.663
R418 B.n584 B.n73 256.663
R419 B.n584 B.n72 256.663
R420 B.n584 B.n71 256.663
R421 B.n584 B.n70 256.663
R422 B.n584 B.n69 256.663
R423 B.n584 B.n68 256.663
R424 B.n584 B.n67 256.663
R425 B.n584 B.n66 256.663
R426 B.n584 B.n65 256.663
R427 B.n584 B.n64 256.663
R428 B.n584 B.n63 256.663
R429 B.n584 B.n62 256.663
R430 B.n584 B.n61 256.663
R431 B.n584 B.n60 256.663
R432 B.n584 B.n59 256.663
R433 B.n584 B.n58 256.663
R434 B.n584 B.n57 256.663
R435 B.n584 B.n56 256.663
R436 B.n584 B.n55 256.663
R437 B.n584 B.n54 256.663
R438 B.n584 B.n53 256.663
R439 B.n584 B.n52 256.663
R440 B.n584 B.n51 256.663
R441 B.n584 B.n50 256.663
R442 B.n584 B.n49 256.663
R443 B.n584 B.n48 256.663
R444 B.n584 B.n47 256.663
R445 B.n584 B.n46 256.663
R446 B.n584 B.n45 256.663
R447 B.n584 B.n44 256.663
R448 B.n584 B.n43 256.663
R449 B.n584 B.n42 256.663
R450 B.n584 B.n41 256.663
R451 B.n584 B.n40 256.663
R452 B.n585 B.n584 256.663
R453 B.n496 B.n495 256.663
R454 B.n495 B.n285 256.663
R455 B.n495 B.n286 256.663
R456 B.n495 B.n287 256.663
R457 B.n495 B.n288 256.663
R458 B.n495 B.n289 256.663
R459 B.n495 B.n290 256.663
R460 B.n495 B.n291 256.663
R461 B.n495 B.n292 256.663
R462 B.n495 B.n293 256.663
R463 B.n495 B.n294 256.663
R464 B.n495 B.n295 256.663
R465 B.n495 B.n296 256.663
R466 B.n495 B.n297 256.663
R467 B.n495 B.n298 256.663
R468 B.n495 B.n299 256.663
R469 B.n495 B.n300 256.663
R470 B.n495 B.n301 256.663
R471 B.n495 B.n302 256.663
R472 B.n495 B.n303 256.663
R473 B.n495 B.n304 256.663
R474 B.n495 B.n305 256.663
R475 B.n495 B.n306 256.663
R476 B.n495 B.n307 256.663
R477 B.n495 B.n308 256.663
R478 B.n495 B.n309 256.663
R479 B.n495 B.n310 256.663
R480 B.n495 B.n311 256.663
R481 B.n495 B.n312 256.663
R482 B.n495 B.n313 256.663
R483 B.n495 B.n314 256.663
R484 B.n495 B.n315 256.663
R485 B.n495 B.n316 256.663
R486 B.n495 B.n317 256.663
R487 B.n495 B.n318 256.663
R488 B.n495 B.n319 256.663
R489 B.n495 B.n320 256.663
R490 B.n495 B.n321 256.663
R491 B.n495 B.n322 256.663
R492 B.n495 B.n323 256.663
R493 B.n495 B.n324 256.663
R494 B.n501 B.n282 163.367
R495 B.n501 B.n276 163.367
R496 B.n510 B.n276 163.367
R497 B.n510 B.n274 163.367
R498 B.n514 B.n274 163.367
R499 B.n514 B.n269 163.367
R500 B.n522 B.n269 163.367
R501 B.n522 B.n267 163.367
R502 B.n526 B.n267 163.367
R503 B.n526 B.n261 163.367
R504 B.n534 B.n261 163.367
R505 B.n534 B.n259 163.367
R506 B.n538 B.n259 163.367
R507 B.n538 B.n253 163.367
R508 B.n548 B.n253 163.367
R509 B.n548 B.n251 163.367
R510 B.n552 B.n251 163.367
R511 B.n552 B.n2 163.367
R512 B.n626 B.n2 163.367
R513 B.n626 B.n3 163.367
R514 B.n622 B.n3 163.367
R515 B.n622 B.n8 163.367
R516 B.n618 B.n8 163.367
R517 B.n618 B.n10 163.367
R518 B.n614 B.n10 163.367
R519 B.n614 B.n16 163.367
R520 B.n610 B.n16 163.367
R521 B.n610 B.n18 163.367
R522 B.n606 B.n18 163.367
R523 B.n606 B.n23 163.367
R524 B.n602 B.n23 163.367
R525 B.n602 B.n25 163.367
R526 B.n598 B.n25 163.367
R527 B.n598 B.n29 163.367
R528 B.n594 B.n29 163.367
R529 B.n594 B.n31 163.367
R530 B.n590 B.n31 163.367
R531 B.n590 B.n37 163.367
R532 B.n494 B.n284 163.367
R533 B.n494 B.n326 163.367
R534 B.n490 B.n489 163.367
R535 B.n486 B.n485 163.367
R536 B.n482 B.n481 163.367
R537 B.n478 B.n477 163.367
R538 B.n474 B.n473 163.367
R539 B.n470 B.n469 163.367
R540 B.n466 B.n465 163.367
R541 B.n462 B.n461 163.367
R542 B.n458 B.n457 163.367
R543 B.n454 B.n453 163.367
R544 B.n450 B.n449 163.367
R545 B.n446 B.n445 163.367
R546 B.n442 B.n441 163.367
R547 B.n438 B.n437 163.367
R548 B.n434 B.n433 163.367
R549 B.n430 B.n429 163.367
R550 B.n426 B.n425 163.367
R551 B.n422 B.n421 163.367
R552 B.n418 B.n417 163.367
R553 B.n414 B.n413 163.367
R554 B.n410 B.n409 163.367
R555 B.n406 B.n405 163.367
R556 B.n402 B.n401 163.367
R557 B.n398 B.n397 163.367
R558 B.n394 B.n393 163.367
R559 B.n390 B.n389 163.367
R560 B.n386 B.n385 163.367
R561 B.n382 B.n381 163.367
R562 B.n378 B.n377 163.367
R563 B.n374 B.n373 163.367
R564 B.n370 B.n369 163.367
R565 B.n366 B.n365 163.367
R566 B.n362 B.n361 163.367
R567 B.n358 B.n357 163.367
R568 B.n354 B.n353 163.367
R569 B.n350 B.n349 163.367
R570 B.n346 B.n345 163.367
R571 B.n342 B.n341 163.367
R572 B.n338 B.n337 163.367
R573 B.n334 B.n325 163.367
R574 B.n503 B.n280 163.367
R575 B.n503 B.n278 163.367
R576 B.n507 B.n278 163.367
R577 B.n507 B.n273 163.367
R578 B.n516 B.n273 163.367
R579 B.n516 B.n271 163.367
R580 B.n520 B.n271 163.367
R581 B.n520 B.n265 163.367
R582 B.n528 B.n265 163.367
R583 B.n528 B.n263 163.367
R584 B.n532 B.n263 163.367
R585 B.n532 B.n256 163.367
R586 B.n540 B.n256 163.367
R587 B.n540 B.n254 163.367
R588 B.n545 B.n254 163.367
R589 B.n545 B.n250 163.367
R590 B.n554 B.n250 163.367
R591 B.n555 B.n554 163.367
R592 B.n555 B.n5 163.367
R593 B.n6 B.n5 163.367
R594 B.n7 B.n6 163.367
R595 B.n560 B.n7 163.367
R596 B.n560 B.n12 163.367
R597 B.n13 B.n12 163.367
R598 B.n14 B.n13 163.367
R599 B.n565 B.n14 163.367
R600 B.n565 B.n19 163.367
R601 B.n20 B.n19 163.367
R602 B.n21 B.n20 163.367
R603 B.n570 B.n21 163.367
R604 B.n570 B.n26 163.367
R605 B.n27 B.n26 163.367
R606 B.n28 B.n27 163.367
R607 B.n575 B.n28 163.367
R608 B.n575 B.n33 163.367
R609 B.n34 B.n33 163.367
R610 B.n35 B.n34 163.367
R611 B.n81 B.n35 163.367
R612 B.n86 B.n39 163.367
R613 B.n90 B.n89 163.367
R614 B.n94 B.n93 163.367
R615 B.n98 B.n97 163.367
R616 B.n102 B.n101 163.367
R617 B.n106 B.n105 163.367
R618 B.n110 B.n109 163.367
R619 B.n114 B.n113 163.367
R620 B.n118 B.n117 163.367
R621 B.n122 B.n121 163.367
R622 B.n126 B.n125 163.367
R623 B.n130 B.n129 163.367
R624 B.n134 B.n133 163.367
R625 B.n138 B.n137 163.367
R626 B.n142 B.n141 163.367
R627 B.n146 B.n145 163.367
R628 B.n150 B.n149 163.367
R629 B.n154 B.n153 163.367
R630 B.n159 B.n158 163.367
R631 B.n163 B.n162 163.367
R632 B.n167 B.n166 163.367
R633 B.n171 B.n170 163.367
R634 B.n175 B.n174 163.367
R635 B.n180 B.n179 163.367
R636 B.n184 B.n183 163.367
R637 B.n188 B.n187 163.367
R638 B.n192 B.n191 163.367
R639 B.n196 B.n195 163.367
R640 B.n200 B.n199 163.367
R641 B.n204 B.n203 163.367
R642 B.n208 B.n207 163.367
R643 B.n212 B.n211 163.367
R644 B.n216 B.n215 163.367
R645 B.n220 B.n219 163.367
R646 B.n224 B.n223 163.367
R647 B.n228 B.n227 163.367
R648 B.n232 B.n231 163.367
R649 B.n236 B.n235 163.367
R650 B.n240 B.n239 163.367
R651 B.n244 B.n243 163.367
R652 B.n246 B.n80 163.367
R653 B.n495 B.n281 92.5661
R654 B.n584 B.n36 92.5661
R655 B.n330 B.t18 88.9632
R656 B.n82 B.t10 88.9632
R657 B.n327 B.t15 88.9505
R658 B.n84 B.t20 88.9505
R659 B.n331 B.t17 74.4178
R660 B.n83 B.t11 74.4178
R661 B.n328 B.t14 74.405
R662 B.n85 B.t21 74.405
R663 B.n497 B.n496 71.676
R664 B.n326 B.n285 71.676
R665 B.n489 B.n286 71.676
R666 B.n485 B.n287 71.676
R667 B.n481 B.n288 71.676
R668 B.n477 B.n289 71.676
R669 B.n473 B.n290 71.676
R670 B.n469 B.n291 71.676
R671 B.n465 B.n292 71.676
R672 B.n461 B.n293 71.676
R673 B.n457 B.n294 71.676
R674 B.n453 B.n295 71.676
R675 B.n449 B.n296 71.676
R676 B.n445 B.n297 71.676
R677 B.n441 B.n298 71.676
R678 B.n437 B.n299 71.676
R679 B.n433 B.n300 71.676
R680 B.n429 B.n301 71.676
R681 B.n425 B.n302 71.676
R682 B.n421 B.n303 71.676
R683 B.n417 B.n304 71.676
R684 B.n413 B.n305 71.676
R685 B.n409 B.n306 71.676
R686 B.n405 B.n307 71.676
R687 B.n401 B.n308 71.676
R688 B.n397 B.n309 71.676
R689 B.n393 B.n310 71.676
R690 B.n389 B.n311 71.676
R691 B.n385 B.n312 71.676
R692 B.n381 B.n313 71.676
R693 B.n377 B.n314 71.676
R694 B.n373 B.n315 71.676
R695 B.n369 B.n316 71.676
R696 B.n365 B.n317 71.676
R697 B.n361 B.n318 71.676
R698 B.n357 B.n319 71.676
R699 B.n353 B.n320 71.676
R700 B.n349 B.n321 71.676
R701 B.n345 B.n322 71.676
R702 B.n341 B.n323 71.676
R703 B.n337 B.n324 71.676
R704 B.n586 B.n585 71.676
R705 B.n86 B.n40 71.676
R706 B.n90 B.n41 71.676
R707 B.n94 B.n42 71.676
R708 B.n98 B.n43 71.676
R709 B.n102 B.n44 71.676
R710 B.n106 B.n45 71.676
R711 B.n110 B.n46 71.676
R712 B.n114 B.n47 71.676
R713 B.n118 B.n48 71.676
R714 B.n122 B.n49 71.676
R715 B.n126 B.n50 71.676
R716 B.n130 B.n51 71.676
R717 B.n134 B.n52 71.676
R718 B.n138 B.n53 71.676
R719 B.n142 B.n54 71.676
R720 B.n146 B.n55 71.676
R721 B.n150 B.n56 71.676
R722 B.n154 B.n57 71.676
R723 B.n159 B.n58 71.676
R724 B.n163 B.n59 71.676
R725 B.n167 B.n60 71.676
R726 B.n171 B.n61 71.676
R727 B.n175 B.n62 71.676
R728 B.n180 B.n63 71.676
R729 B.n184 B.n64 71.676
R730 B.n188 B.n65 71.676
R731 B.n192 B.n66 71.676
R732 B.n196 B.n67 71.676
R733 B.n200 B.n68 71.676
R734 B.n204 B.n69 71.676
R735 B.n208 B.n70 71.676
R736 B.n212 B.n71 71.676
R737 B.n216 B.n72 71.676
R738 B.n220 B.n73 71.676
R739 B.n224 B.n74 71.676
R740 B.n228 B.n75 71.676
R741 B.n232 B.n76 71.676
R742 B.n236 B.n77 71.676
R743 B.n240 B.n78 71.676
R744 B.n244 B.n79 71.676
R745 B.n583 B.n80 71.676
R746 B.n583 B.n582 71.676
R747 B.n246 B.n79 71.676
R748 B.n243 B.n78 71.676
R749 B.n239 B.n77 71.676
R750 B.n235 B.n76 71.676
R751 B.n231 B.n75 71.676
R752 B.n227 B.n74 71.676
R753 B.n223 B.n73 71.676
R754 B.n219 B.n72 71.676
R755 B.n215 B.n71 71.676
R756 B.n211 B.n70 71.676
R757 B.n207 B.n69 71.676
R758 B.n203 B.n68 71.676
R759 B.n199 B.n67 71.676
R760 B.n195 B.n66 71.676
R761 B.n191 B.n65 71.676
R762 B.n187 B.n64 71.676
R763 B.n183 B.n63 71.676
R764 B.n179 B.n62 71.676
R765 B.n174 B.n61 71.676
R766 B.n170 B.n60 71.676
R767 B.n166 B.n59 71.676
R768 B.n162 B.n58 71.676
R769 B.n158 B.n57 71.676
R770 B.n153 B.n56 71.676
R771 B.n149 B.n55 71.676
R772 B.n145 B.n54 71.676
R773 B.n141 B.n53 71.676
R774 B.n137 B.n52 71.676
R775 B.n133 B.n51 71.676
R776 B.n129 B.n50 71.676
R777 B.n125 B.n49 71.676
R778 B.n121 B.n48 71.676
R779 B.n117 B.n47 71.676
R780 B.n113 B.n46 71.676
R781 B.n109 B.n45 71.676
R782 B.n105 B.n44 71.676
R783 B.n101 B.n43 71.676
R784 B.n97 B.n42 71.676
R785 B.n93 B.n41 71.676
R786 B.n89 B.n40 71.676
R787 B.n585 B.n39 71.676
R788 B.n496 B.n284 71.676
R789 B.n490 B.n285 71.676
R790 B.n486 B.n286 71.676
R791 B.n482 B.n287 71.676
R792 B.n478 B.n288 71.676
R793 B.n474 B.n289 71.676
R794 B.n470 B.n290 71.676
R795 B.n466 B.n291 71.676
R796 B.n462 B.n292 71.676
R797 B.n458 B.n293 71.676
R798 B.n454 B.n294 71.676
R799 B.n450 B.n295 71.676
R800 B.n446 B.n296 71.676
R801 B.n442 B.n297 71.676
R802 B.n438 B.n298 71.676
R803 B.n434 B.n299 71.676
R804 B.n430 B.n300 71.676
R805 B.n426 B.n301 71.676
R806 B.n422 B.n302 71.676
R807 B.n418 B.n303 71.676
R808 B.n414 B.n304 71.676
R809 B.n410 B.n305 71.676
R810 B.n406 B.n306 71.676
R811 B.n402 B.n307 71.676
R812 B.n398 B.n308 71.676
R813 B.n394 B.n309 71.676
R814 B.n390 B.n310 71.676
R815 B.n386 B.n311 71.676
R816 B.n382 B.n312 71.676
R817 B.n378 B.n313 71.676
R818 B.n374 B.n314 71.676
R819 B.n370 B.n315 71.676
R820 B.n366 B.n316 71.676
R821 B.n362 B.n317 71.676
R822 B.n358 B.n318 71.676
R823 B.n354 B.n319 71.676
R824 B.n350 B.n320 71.676
R825 B.n346 B.n321 71.676
R826 B.n342 B.n322 71.676
R827 B.n338 B.n323 71.676
R828 B.n334 B.n324 71.676
R829 B.n332 B.n331 59.5399
R830 B.n329 B.n328 59.5399
R831 B.n156 B.n85 59.5399
R832 B.n177 B.n83 59.5399
R833 B.n502 B.n281 47.3273
R834 B.n502 B.n277 47.3273
R835 B.n509 B.n277 47.3273
R836 B.n509 B.n508 47.3273
R837 B.n515 B.n270 47.3273
R838 B.n521 B.n270 47.3273
R839 B.n521 B.n266 47.3273
R840 B.n527 B.n266 47.3273
R841 B.n533 B.n262 47.3273
R842 B.n539 B.n257 47.3273
R843 B.n539 B.n258 47.3273
R844 B.n547 B.n546 47.3273
R845 B.n553 B.n4 47.3273
R846 B.n625 B.n4 47.3273
R847 B.n625 B.n624 47.3273
R848 B.n624 B.n623 47.3273
R849 B.n617 B.n11 47.3273
R850 B.n616 B.n615 47.3273
R851 B.n615 B.n15 47.3273
R852 B.n609 B.n608 47.3273
R853 B.n607 B.n22 47.3273
R854 B.n601 B.n22 47.3273
R855 B.n601 B.n600 47.3273
R856 B.n600 B.n599 47.3273
R857 B.n593 B.n32 47.3273
R858 B.n593 B.n592 47.3273
R859 B.n592 B.n591 47.3273
R860 B.n591 B.n36 47.3273
R861 B.n547 B.t7 43.1514
R862 B.n617 B.t2 43.1514
R863 B.n533 B.t1 41.7594
R864 B.n609 B.t4 41.7594
R865 B.n588 B.n587 34.8103
R866 B.n581 B.n580 34.8103
R867 B.n333 B.n279 34.8103
R868 B.n499 B.n498 34.8103
R869 B.n515 B.t13 34.7996
R870 B.n599 B.t9 34.7996
R871 B.n553 B.t5 33.4077
R872 B.n623 B.t6 33.4077
R873 B.n527 B.t3 32.0157
R874 B.t0 B.n607 32.0157
R875 B B.n627 18.0485
R876 B.t3 B.n262 15.3121
R877 B.n608 B.t0 15.3121
R878 B.n331 B.n330 14.546
R879 B.n328 B.n327 14.546
R880 B.n85 B.n84 14.546
R881 B.n83 B.n82 14.546
R882 B.n546 B.t5 13.9201
R883 B.n11 B.t6 13.9201
R884 B.n508 B.t13 12.5282
R885 B.n32 B.t9 12.5282
R886 B.n587 B.n38 10.6151
R887 B.n87 B.n38 10.6151
R888 B.n88 B.n87 10.6151
R889 B.n91 B.n88 10.6151
R890 B.n92 B.n91 10.6151
R891 B.n95 B.n92 10.6151
R892 B.n96 B.n95 10.6151
R893 B.n99 B.n96 10.6151
R894 B.n100 B.n99 10.6151
R895 B.n103 B.n100 10.6151
R896 B.n104 B.n103 10.6151
R897 B.n107 B.n104 10.6151
R898 B.n108 B.n107 10.6151
R899 B.n111 B.n108 10.6151
R900 B.n112 B.n111 10.6151
R901 B.n115 B.n112 10.6151
R902 B.n116 B.n115 10.6151
R903 B.n119 B.n116 10.6151
R904 B.n120 B.n119 10.6151
R905 B.n123 B.n120 10.6151
R906 B.n124 B.n123 10.6151
R907 B.n127 B.n124 10.6151
R908 B.n128 B.n127 10.6151
R909 B.n131 B.n128 10.6151
R910 B.n132 B.n131 10.6151
R911 B.n135 B.n132 10.6151
R912 B.n136 B.n135 10.6151
R913 B.n139 B.n136 10.6151
R914 B.n140 B.n139 10.6151
R915 B.n143 B.n140 10.6151
R916 B.n144 B.n143 10.6151
R917 B.n147 B.n144 10.6151
R918 B.n148 B.n147 10.6151
R919 B.n151 B.n148 10.6151
R920 B.n152 B.n151 10.6151
R921 B.n155 B.n152 10.6151
R922 B.n160 B.n157 10.6151
R923 B.n161 B.n160 10.6151
R924 B.n164 B.n161 10.6151
R925 B.n165 B.n164 10.6151
R926 B.n168 B.n165 10.6151
R927 B.n169 B.n168 10.6151
R928 B.n172 B.n169 10.6151
R929 B.n173 B.n172 10.6151
R930 B.n176 B.n173 10.6151
R931 B.n181 B.n178 10.6151
R932 B.n182 B.n181 10.6151
R933 B.n185 B.n182 10.6151
R934 B.n186 B.n185 10.6151
R935 B.n189 B.n186 10.6151
R936 B.n190 B.n189 10.6151
R937 B.n193 B.n190 10.6151
R938 B.n194 B.n193 10.6151
R939 B.n197 B.n194 10.6151
R940 B.n198 B.n197 10.6151
R941 B.n201 B.n198 10.6151
R942 B.n202 B.n201 10.6151
R943 B.n205 B.n202 10.6151
R944 B.n206 B.n205 10.6151
R945 B.n209 B.n206 10.6151
R946 B.n210 B.n209 10.6151
R947 B.n213 B.n210 10.6151
R948 B.n214 B.n213 10.6151
R949 B.n217 B.n214 10.6151
R950 B.n218 B.n217 10.6151
R951 B.n221 B.n218 10.6151
R952 B.n222 B.n221 10.6151
R953 B.n225 B.n222 10.6151
R954 B.n226 B.n225 10.6151
R955 B.n229 B.n226 10.6151
R956 B.n230 B.n229 10.6151
R957 B.n233 B.n230 10.6151
R958 B.n234 B.n233 10.6151
R959 B.n237 B.n234 10.6151
R960 B.n238 B.n237 10.6151
R961 B.n241 B.n238 10.6151
R962 B.n242 B.n241 10.6151
R963 B.n245 B.n242 10.6151
R964 B.n247 B.n245 10.6151
R965 B.n248 B.n247 10.6151
R966 B.n581 B.n248 10.6151
R967 B.n504 B.n279 10.6151
R968 B.n505 B.n504 10.6151
R969 B.n506 B.n505 10.6151
R970 B.n506 B.n272 10.6151
R971 B.n517 B.n272 10.6151
R972 B.n518 B.n517 10.6151
R973 B.n519 B.n518 10.6151
R974 B.n519 B.n264 10.6151
R975 B.n529 B.n264 10.6151
R976 B.n530 B.n529 10.6151
R977 B.n531 B.n530 10.6151
R978 B.n531 B.n255 10.6151
R979 B.n541 B.n255 10.6151
R980 B.n542 B.n541 10.6151
R981 B.n544 B.n542 10.6151
R982 B.n544 B.n543 10.6151
R983 B.n543 B.n249 10.6151
R984 B.n556 B.n249 10.6151
R985 B.n557 B.n556 10.6151
R986 B.n558 B.n557 10.6151
R987 B.n559 B.n558 10.6151
R988 B.n561 B.n559 10.6151
R989 B.n562 B.n561 10.6151
R990 B.n563 B.n562 10.6151
R991 B.n564 B.n563 10.6151
R992 B.n566 B.n564 10.6151
R993 B.n567 B.n566 10.6151
R994 B.n568 B.n567 10.6151
R995 B.n569 B.n568 10.6151
R996 B.n571 B.n569 10.6151
R997 B.n572 B.n571 10.6151
R998 B.n573 B.n572 10.6151
R999 B.n574 B.n573 10.6151
R1000 B.n576 B.n574 10.6151
R1001 B.n577 B.n576 10.6151
R1002 B.n578 B.n577 10.6151
R1003 B.n579 B.n578 10.6151
R1004 B.n580 B.n579 10.6151
R1005 B.n498 B.n283 10.6151
R1006 B.n493 B.n283 10.6151
R1007 B.n493 B.n492 10.6151
R1008 B.n492 B.n491 10.6151
R1009 B.n491 B.n488 10.6151
R1010 B.n488 B.n487 10.6151
R1011 B.n487 B.n484 10.6151
R1012 B.n484 B.n483 10.6151
R1013 B.n483 B.n480 10.6151
R1014 B.n480 B.n479 10.6151
R1015 B.n479 B.n476 10.6151
R1016 B.n476 B.n475 10.6151
R1017 B.n475 B.n472 10.6151
R1018 B.n472 B.n471 10.6151
R1019 B.n471 B.n468 10.6151
R1020 B.n468 B.n467 10.6151
R1021 B.n467 B.n464 10.6151
R1022 B.n464 B.n463 10.6151
R1023 B.n463 B.n460 10.6151
R1024 B.n460 B.n459 10.6151
R1025 B.n459 B.n456 10.6151
R1026 B.n456 B.n455 10.6151
R1027 B.n455 B.n452 10.6151
R1028 B.n452 B.n451 10.6151
R1029 B.n451 B.n448 10.6151
R1030 B.n448 B.n447 10.6151
R1031 B.n447 B.n444 10.6151
R1032 B.n444 B.n443 10.6151
R1033 B.n443 B.n440 10.6151
R1034 B.n440 B.n439 10.6151
R1035 B.n439 B.n436 10.6151
R1036 B.n436 B.n435 10.6151
R1037 B.n435 B.n432 10.6151
R1038 B.n432 B.n431 10.6151
R1039 B.n431 B.n428 10.6151
R1040 B.n428 B.n427 10.6151
R1041 B.n424 B.n423 10.6151
R1042 B.n423 B.n420 10.6151
R1043 B.n420 B.n419 10.6151
R1044 B.n419 B.n416 10.6151
R1045 B.n416 B.n415 10.6151
R1046 B.n415 B.n412 10.6151
R1047 B.n412 B.n411 10.6151
R1048 B.n411 B.n408 10.6151
R1049 B.n408 B.n407 10.6151
R1050 B.n404 B.n403 10.6151
R1051 B.n403 B.n400 10.6151
R1052 B.n400 B.n399 10.6151
R1053 B.n399 B.n396 10.6151
R1054 B.n396 B.n395 10.6151
R1055 B.n395 B.n392 10.6151
R1056 B.n392 B.n391 10.6151
R1057 B.n391 B.n388 10.6151
R1058 B.n388 B.n387 10.6151
R1059 B.n387 B.n384 10.6151
R1060 B.n384 B.n383 10.6151
R1061 B.n383 B.n380 10.6151
R1062 B.n380 B.n379 10.6151
R1063 B.n379 B.n376 10.6151
R1064 B.n376 B.n375 10.6151
R1065 B.n375 B.n372 10.6151
R1066 B.n372 B.n371 10.6151
R1067 B.n371 B.n368 10.6151
R1068 B.n368 B.n367 10.6151
R1069 B.n367 B.n364 10.6151
R1070 B.n364 B.n363 10.6151
R1071 B.n363 B.n360 10.6151
R1072 B.n360 B.n359 10.6151
R1073 B.n359 B.n356 10.6151
R1074 B.n356 B.n355 10.6151
R1075 B.n355 B.n352 10.6151
R1076 B.n352 B.n351 10.6151
R1077 B.n351 B.n348 10.6151
R1078 B.n348 B.n347 10.6151
R1079 B.n347 B.n344 10.6151
R1080 B.n344 B.n343 10.6151
R1081 B.n343 B.n340 10.6151
R1082 B.n340 B.n339 10.6151
R1083 B.n339 B.n336 10.6151
R1084 B.n336 B.n335 10.6151
R1085 B.n335 B.n333 10.6151
R1086 B.n500 B.n499 10.6151
R1087 B.n500 B.n275 10.6151
R1088 B.n511 B.n275 10.6151
R1089 B.n512 B.n511 10.6151
R1090 B.n513 B.n512 10.6151
R1091 B.n513 B.n268 10.6151
R1092 B.n523 B.n268 10.6151
R1093 B.n524 B.n523 10.6151
R1094 B.n525 B.n524 10.6151
R1095 B.n525 B.n260 10.6151
R1096 B.n535 B.n260 10.6151
R1097 B.n536 B.n535 10.6151
R1098 B.n537 B.n536 10.6151
R1099 B.n537 B.n252 10.6151
R1100 B.n549 B.n252 10.6151
R1101 B.n550 B.n549 10.6151
R1102 B.n551 B.n550 10.6151
R1103 B.n551 B.n0 10.6151
R1104 B.n621 B.n1 10.6151
R1105 B.n621 B.n620 10.6151
R1106 B.n620 B.n619 10.6151
R1107 B.n619 B.n9 10.6151
R1108 B.n613 B.n9 10.6151
R1109 B.n613 B.n612 10.6151
R1110 B.n612 B.n611 10.6151
R1111 B.n611 B.n17 10.6151
R1112 B.n605 B.n17 10.6151
R1113 B.n605 B.n604 10.6151
R1114 B.n604 B.n603 10.6151
R1115 B.n603 B.n24 10.6151
R1116 B.n597 B.n24 10.6151
R1117 B.n597 B.n596 10.6151
R1118 B.n596 B.n595 10.6151
R1119 B.n595 B.n30 10.6151
R1120 B.n589 B.n30 10.6151
R1121 B.n589 B.n588 10.6151
R1122 B.n156 B.n155 9.36635
R1123 B.n178 B.n177 9.36635
R1124 B.n427 B.n329 9.36635
R1125 B.n404 B.n332 9.36635
R1126 B.t1 B.n257 5.56836
R1127 B.t4 B.n15 5.56836
R1128 B.n258 B.t7 4.17639
R1129 B.t2 B.n616 4.17639
R1130 B.n627 B.n0 2.81026
R1131 B.n627 B.n1 2.81026
R1132 B.n157 B.n156 1.24928
R1133 B.n177 B.n176 1.24928
R1134 B.n424 B.n329 1.24928
R1135 B.n407 B.n332 1.24928
R1136 VP.n4 VP.t1 719.308
R1137 VP.n10 VP.t0 698.327
R1138 VP.n1 VP.t4 698.327
R1139 VP.n15 VP.t3 698.327
R1140 VP.n16 VP.t6 698.327
R1141 VP.n8 VP.t7 698.327
R1142 VP.n7 VP.t2 698.327
R1143 VP.n3 VP.t5 698.327
R1144 VP.n17 VP.n16 161.3
R1145 VP.n6 VP.n5 161.3
R1146 VP.n7 VP.n2 161.3
R1147 VP.n9 VP.n8 161.3
R1148 VP.n15 VP.n0 161.3
R1149 VP.n14 VP.n13 161.3
R1150 VP.n12 VP.n1 161.3
R1151 VP.n11 VP.n10 161.3
R1152 VP.n5 VP.n4 70.4033
R1153 VP.n10 VP.n1 48.2005
R1154 VP.n16 VP.n15 48.2005
R1155 VP.n8 VP.n7 48.2005
R1156 VP.n11 VP.n9 39.5611
R1157 VP.n14 VP.n1 24.1005
R1158 VP.n15 VP.n14 24.1005
R1159 VP.n6 VP.n3 24.1005
R1160 VP.n7 VP.n6 24.1005
R1161 VP.n4 VP.n3 20.9576
R1162 VP.n5 VP.n2 0.189894
R1163 VP.n9 VP.n2 0.189894
R1164 VP.n12 VP.n11 0.189894
R1165 VP.n13 VP.n12 0.189894
R1166 VP.n13 VP.n0 0.189894
R1167 VP.n17 VP.n0 0.189894
R1168 VP VP.n17 0.0516364
R1169 VDD1 VDD1.n0 66.9372
R1170 VDD1.n3 VDD1.n2 66.8234
R1171 VDD1.n3 VDD1.n1 66.8234
R1172 VDD1.n5 VDD1.n4 66.5556
R1173 VDD1.n5 VDD1.n3 36.2854
R1174 VDD1.n4 VDD1.t5 1.88084
R1175 VDD1.n4 VDD1.t0 1.88084
R1176 VDD1.n0 VDD1.t6 1.88084
R1177 VDD1.n0 VDD1.t2 1.88084
R1178 VDD1.n2 VDD1.t4 1.88084
R1179 VDD1.n2 VDD1.t1 1.88084
R1180 VDD1.n1 VDD1.t7 1.88084
R1181 VDD1.n1 VDD1.t3 1.88084
R1182 VDD1 VDD1.n5 0.265586
C0 VDD1 VTAIL 12.5554f
C1 VDD1 VDD2 0.689803f
C2 VDD1 VP 3.79561f
C3 VTAIL VN 3.3608f
C4 VDD2 VN 3.65599f
C5 VP VN 4.72715f
C6 VTAIL VDD2 12.595201f
C7 VP VTAIL 3.37491f
C8 VP VDD2 0.28773f
C9 VDD1 VN 0.147821f
C10 VDD2 B 3.123835f
C11 VDD1 B 3.329986f
C12 VTAIL B 7.81226f
C13 VN B 7.49325f
C14 VP B 5.437992f
C15 VDD1.t6 B 0.253721f
C16 VDD1.t2 B 0.253721f
C17 VDD1.n0 B 2.24812f
C18 VDD1.t7 B 0.253721f
C19 VDD1.t3 B 0.253721f
C20 VDD1.n1 B 2.24748f
C21 VDD1.t4 B 0.253721f
C22 VDD1.t1 B 0.253721f
C23 VDD1.n2 B 2.24748f
C24 VDD1.n3 B 2.39571f
C25 VDD1.t5 B 0.253721f
C26 VDD1.t0 B 0.253721f
C27 VDD1.n4 B 2.24607f
C28 VDD1.n5 B 2.56492f
C29 VP.n0 B 0.052241f
C30 VP.t4 B 0.660608f
C31 VP.n1 B 0.280142f
C32 VP.n2 B 0.052241f
C33 VP.t7 B 0.660608f
C34 VP.t2 B 0.660608f
C35 VP.t5 B 0.660608f
C36 VP.n3 B 0.280142f
C37 VP.t1 B 0.668626f
C38 VP.n4 B 0.267172f
C39 VP.n5 B 0.161836f
C40 VP.n6 B 0.011855f
C41 VP.n7 B 0.280142f
C42 VP.n8 B 0.274827f
C43 VP.n9 B 1.9476f
C44 VP.t0 B 0.660608f
C45 VP.n10 B 0.274827f
C46 VP.n11 B 1.99507f
C47 VP.n12 B 0.052241f
C48 VP.n13 B 0.052241f
C49 VP.n14 B 0.011855f
C50 VP.t3 B 0.660608f
C51 VP.n15 B 0.280142f
C52 VP.t6 B 0.660608f
C53 VP.n16 B 0.274827f
C54 VP.n17 B 0.040485f
C55 VTAIL.t11 B 0.186009f
C56 VTAIL.t10 B 0.186009f
C57 VTAIL.n0 B 1.58783f
C58 VTAIL.n1 B 0.259328f
C59 VTAIL.t8 B 2.02577f
C60 VTAIL.n2 B 0.358338f
C61 VTAIL.t15 B 2.02577f
C62 VTAIL.n3 B 0.358338f
C63 VTAIL.t1 B 0.186009f
C64 VTAIL.t13 B 0.186009f
C65 VTAIL.n4 B 1.58783f
C66 VTAIL.n5 B 0.301708f
C67 VTAIL.t3 B 2.02577f
C68 VTAIL.n6 B 1.32857f
C69 VTAIL.t9 B 2.02577f
C70 VTAIL.n7 B 1.32856f
C71 VTAIL.t6 B 0.186009f
C72 VTAIL.t12 B 0.186009f
C73 VTAIL.n8 B 1.58784f
C74 VTAIL.n9 B 0.301703f
C75 VTAIL.t7 B 2.02577f
C76 VTAIL.n10 B 0.358333f
C77 VTAIL.t14 B 2.02577f
C78 VTAIL.n11 B 0.358333f
C79 VTAIL.t2 B 0.186009f
C80 VTAIL.t4 B 0.186009f
C81 VTAIL.n12 B 1.58784f
C82 VTAIL.n13 B 0.301703f
C83 VTAIL.t0 B 2.02577f
C84 VTAIL.n14 B 1.32857f
C85 VTAIL.t5 B 2.02577f
C86 VTAIL.n15 B 1.32437f
C87 VDD2.t6 B 0.253918f
C88 VDD2.t2 B 0.253918f
C89 VDD2.n0 B 2.24922f
C90 VDD2.t4 B 0.253918f
C91 VDD2.t5 B 0.253918f
C92 VDD2.n1 B 2.24922f
C93 VDD2.n2 B 2.33207f
C94 VDD2.t7 B 0.253918f
C95 VDD2.t1 B 0.253918f
C96 VDD2.n3 B 2.24781f
C97 VDD2.n4 B 2.53113f
C98 VDD2.t3 B 0.253918f
C99 VDD2.t0 B 0.253918f
C100 VDD2.n5 B 2.24919f
C101 VN.n0 B 0.051485f
C102 VN.t1 B 0.651039f
C103 VN.n1 B 0.276084f
C104 VN.t4 B 0.658941f
C105 VN.n2 B 0.263302f
C106 VN.n3 B 0.159492f
C107 VN.n4 B 0.011683f
C108 VN.t2 B 0.651039f
C109 VN.n5 B 0.276084f
C110 VN.t7 B 0.651039f
C111 VN.n6 B 0.270846f
C112 VN.n7 B 0.039899f
C113 VN.n8 B 0.051485f
C114 VN.t0 B 0.651039f
C115 VN.n9 B 0.276084f
C116 VN.t5 B 0.658941f
C117 VN.n10 B 0.263302f
C118 VN.n11 B 0.159492f
C119 VN.n12 B 0.011683f
C120 VN.t6 B 0.651039f
C121 VN.n13 B 0.276084f
C122 VN.t3 B 0.651039f
C123 VN.n14 B 0.270846f
C124 VN.n15 B 1.95332f
.ends

