* NGSPICE file created from diff_pair_sample_0460.ext - technology: sky130A

.subckt diff_pair_sample_0460 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6575 pd=9.28 as=0 ps=0 w=4.25 l=0.77
X1 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=1.6575 pd=9.28 as=0 ps=0 w=4.25 l=0.77
X2 VTAIL.t7 VP.t0 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6575 pd=9.28 as=0.70125 ps=4.58 w=4.25 l=0.77
X3 VDD2.t3 VN.t0 VTAIL.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.70125 pd=4.58 as=1.6575 ps=9.28 w=4.25 l=0.77
X4 VTAIL.t3 VN.t1 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6575 pd=9.28 as=0.70125 ps=4.58 w=4.25 l=0.77
X5 VTAIL.t6 VP.t1 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6575 pd=9.28 as=0.70125 ps=4.58 w=4.25 l=0.77
X6 VDD2.t1 VN.t2 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.70125 pd=4.58 as=1.6575 ps=9.28 w=4.25 l=0.77
X7 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.6575 pd=9.28 as=0 ps=0 w=4.25 l=0.77
X8 VTAIL.t1 VN.t3 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6575 pd=9.28 as=0.70125 ps=4.58 w=4.25 l=0.77
X9 VDD1.t2 VP.t2 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.70125 pd=4.58 as=1.6575 ps=9.28 w=4.25 l=0.77
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6575 pd=9.28 as=0 ps=0 w=4.25 l=0.77
X11 VDD1.t1 VP.t3 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.70125 pd=4.58 as=1.6575 ps=9.28 w=4.25 l=0.77
R0 B.n300 B.n299 585
R1 B.n300 B.n36 585
R2 B.n303 B.n302 585
R3 B.n304 B.n64 585
R4 B.n306 B.n305 585
R5 B.n308 B.n63 585
R6 B.n311 B.n310 585
R7 B.n312 B.n62 585
R8 B.n314 B.n313 585
R9 B.n316 B.n61 585
R10 B.n319 B.n318 585
R11 B.n320 B.n60 585
R12 B.n322 B.n321 585
R13 B.n324 B.n59 585
R14 B.n327 B.n326 585
R15 B.n328 B.n58 585
R16 B.n330 B.n329 585
R17 B.n332 B.n57 585
R18 B.n335 B.n334 585
R19 B.n336 B.n54 585
R20 B.n339 B.n338 585
R21 B.n341 B.n53 585
R22 B.n344 B.n343 585
R23 B.n345 B.n52 585
R24 B.n347 B.n346 585
R25 B.n349 B.n51 585
R26 B.n352 B.n351 585
R27 B.n353 B.n47 585
R28 B.n355 B.n354 585
R29 B.n357 B.n46 585
R30 B.n360 B.n359 585
R31 B.n361 B.n45 585
R32 B.n363 B.n362 585
R33 B.n365 B.n44 585
R34 B.n368 B.n367 585
R35 B.n369 B.n43 585
R36 B.n371 B.n370 585
R37 B.n373 B.n42 585
R38 B.n376 B.n375 585
R39 B.n377 B.n41 585
R40 B.n379 B.n378 585
R41 B.n381 B.n40 585
R42 B.n384 B.n383 585
R43 B.n385 B.n39 585
R44 B.n387 B.n386 585
R45 B.n389 B.n38 585
R46 B.n392 B.n391 585
R47 B.n393 B.n37 585
R48 B.n298 B.n35 585
R49 B.n396 B.n35 585
R50 B.n297 B.n34 585
R51 B.n397 B.n34 585
R52 B.n296 B.n33 585
R53 B.n398 B.n33 585
R54 B.n295 B.n294 585
R55 B.n294 B.n29 585
R56 B.n293 B.n28 585
R57 B.n404 B.n28 585
R58 B.n292 B.n27 585
R59 B.n405 B.n27 585
R60 B.n291 B.n26 585
R61 B.n406 B.n26 585
R62 B.n290 B.n289 585
R63 B.n289 B.n22 585
R64 B.n288 B.n21 585
R65 B.n412 B.n21 585
R66 B.n287 B.n20 585
R67 B.n413 B.n20 585
R68 B.n286 B.n19 585
R69 B.n414 B.n19 585
R70 B.n285 B.n284 585
R71 B.n284 B.n18 585
R72 B.n283 B.n14 585
R73 B.n420 B.n14 585
R74 B.n282 B.n13 585
R75 B.n421 B.n13 585
R76 B.n281 B.n12 585
R77 B.n422 B.n12 585
R78 B.n280 B.n279 585
R79 B.n279 B.n8 585
R80 B.n278 B.n7 585
R81 B.n428 B.n7 585
R82 B.n277 B.n6 585
R83 B.n429 B.n6 585
R84 B.n276 B.n5 585
R85 B.n430 B.n5 585
R86 B.n275 B.n274 585
R87 B.n274 B.n4 585
R88 B.n273 B.n65 585
R89 B.n273 B.n272 585
R90 B.n263 B.n66 585
R91 B.n67 B.n66 585
R92 B.n265 B.n264 585
R93 B.n266 B.n265 585
R94 B.n262 B.n72 585
R95 B.n72 B.n71 585
R96 B.n261 B.n260 585
R97 B.n260 B.n259 585
R98 B.n74 B.n73 585
R99 B.n252 B.n74 585
R100 B.n251 B.n250 585
R101 B.n253 B.n251 585
R102 B.n249 B.n79 585
R103 B.n79 B.n78 585
R104 B.n248 B.n247 585
R105 B.n247 B.n246 585
R106 B.n81 B.n80 585
R107 B.n82 B.n81 585
R108 B.n239 B.n238 585
R109 B.n240 B.n239 585
R110 B.n237 B.n86 585
R111 B.n90 B.n86 585
R112 B.n236 B.n235 585
R113 B.n235 B.n234 585
R114 B.n88 B.n87 585
R115 B.n89 B.n88 585
R116 B.n227 B.n226 585
R117 B.n228 B.n227 585
R118 B.n225 B.n95 585
R119 B.n95 B.n94 585
R120 B.n224 B.n223 585
R121 B.n223 B.n222 585
R122 B.n219 B.n99 585
R123 B.n218 B.n217 585
R124 B.n215 B.n100 585
R125 B.n215 B.n98 585
R126 B.n214 B.n213 585
R127 B.n212 B.n211 585
R128 B.n210 B.n102 585
R129 B.n208 B.n207 585
R130 B.n206 B.n103 585
R131 B.n205 B.n204 585
R132 B.n202 B.n104 585
R133 B.n200 B.n199 585
R134 B.n198 B.n105 585
R135 B.n197 B.n196 585
R136 B.n194 B.n106 585
R137 B.n192 B.n191 585
R138 B.n190 B.n107 585
R139 B.n189 B.n188 585
R140 B.n186 B.n108 585
R141 B.n184 B.n183 585
R142 B.n181 B.n109 585
R143 B.n180 B.n179 585
R144 B.n177 B.n112 585
R145 B.n175 B.n174 585
R146 B.n173 B.n113 585
R147 B.n172 B.n171 585
R148 B.n169 B.n114 585
R149 B.n167 B.n166 585
R150 B.n165 B.n115 585
R151 B.n163 B.n162 585
R152 B.n160 B.n118 585
R153 B.n158 B.n157 585
R154 B.n156 B.n119 585
R155 B.n155 B.n154 585
R156 B.n152 B.n120 585
R157 B.n150 B.n149 585
R158 B.n148 B.n121 585
R159 B.n147 B.n146 585
R160 B.n144 B.n122 585
R161 B.n142 B.n141 585
R162 B.n140 B.n123 585
R163 B.n139 B.n138 585
R164 B.n136 B.n124 585
R165 B.n134 B.n133 585
R166 B.n132 B.n125 585
R167 B.n131 B.n130 585
R168 B.n128 B.n126 585
R169 B.n97 B.n96 585
R170 B.n221 B.n220 585
R171 B.n222 B.n221 585
R172 B.n93 B.n92 585
R173 B.n94 B.n93 585
R174 B.n230 B.n229 585
R175 B.n229 B.n228 585
R176 B.n231 B.n91 585
R177 B.n91 B.n89 585
R178 B.n233 B.n232 585
R179 B.n234 B.n233 585
R180 B.n85 B.n84 585
R181 B.n90 B.n85 585
R182 B.n242 B.n241 585
R183 B.n241 B.n240 585
R184 B.n243 B.n83 585
R185 B.n83 B.n82 585
R186 B.n245 B.n244 585
R187 B.n246 B.n245 585
R188 B.n77 B.n76 585
R189 B.n78 B.n77 585
R190 B.n255 B.n254 585
R191 B.n254 B.n253 585
R192 B.n256 B.n75 585
R193 B.n252 B.n75 585
R194 B.n258 B.n257 585
R195 B.n259 B.n258 585
R196 B.n70 B.n69 585
R197 B.n71 B.n70 585
R198 B.n268 B.n267 585
R199 B.n267 B.n266 585
R200 B.n269 B.n68 585
R201 B.n68 B.n67 585
R202 B.n271 B.n270 585
R203 B.n272 B.n271 585
R204 B.n2 B.n0 585
R205 B.n4 B.n2 585
R206 B.n3 B.n1 585
R207 B.n429 B.n3 585
R208 B.n427 B.n426 585
R209 B.n428 B.n427 585
R210 B.n425 B.n9 585
R211 B.n9 B.n8 585
R212 B.n424 B.n423 585
R213 B.n423 B.n422 585
R214 B.n11 B.n10 585
R215 B.n421 B.n11 585
R216 B.n419 B.n418 585
R217 B.n420 B.n419 585
R218 B.n417 B.n15 585
R219 B.n18 B.n15 585
R220 B.n416 B.n415 585
R221 B.n415 B.n414 585
R222 B.n17 B.n16 585
R223 B.n413 B.n17 585
R224 B.n411 B.n410 585
R225 B.n412 B.n411 585
R226 B.n409 B.n23 585
R227 B.n23 B.n22 585
R228 B.n408 B.n407 585
R229 B.n407 B.n406 585
R230 B.n25 B.n24 585
R231 B.n405 B.n25 585
R232 B.n403 B.n402 585
R233 B.n404 B.n403 585
R234 B.n401 B.n30 585
R235 B.n30 B.n29 585
R236 B.n400 B.n399 585
R237 B.n399 B.n398 585
R238 B.n32 B.n31 585
R239 B.n397 B.n32 585
R240 B.n395 B.n394 585
R241 B.n396 B.n395 585
R242 B.n432 B.n431 585
R243 B.n431 B.n430 585
R244 B.n221 B.n99 487.695
R245 B.n395 B.n37 487.695
R246 B.n223 B.n97 487.695
R247 B.n300 B.n35 487.695
R248 B.n116 B.t4 335.202
R249 B.n110 B.t15 335.202
R250 B.n48 B.t12 335.202
R251 B.n55 B.t8 335.202
R252 B.n301 B.n36 256.663
R253 B.n307 B.n36 256.663
R254 B.n309 B.n36 256.663
R255 B.n315 B.n36 256.663
R256 B.n317 B.n36 256.663
R257 B.n323 B.n36 256.663
R258 B.n325 B.n36 256.663
R259 B.n331 B.n36 256.663
R260 B.n333 B.n36 256.663
R261 B.n340 B.n36 256.663
R262 B.n342 B.n36 256.663
R263 B.n348 B.n36 256.663
R264 B.n350 B.n36 256.663
R265 B.n356 B.n36 256.663
R266 B.n358 B.n36 256.663
R267 B.n364 B.n36 256.663
R268 B.n366 B.n36 256.663
R269 B.n372 B.n36 256.663
R270 B.n374 B.n36 256.663
R271 B.n380 B.n36 256.663
R272 B.n382 B.n36 256.663
R273 B.n388 B.n36 256.663
R274 B.n390 B.n36 256.663
R275 B.n216 B.n98 256.663
R276 B.n101 B.n98 256.663
R277 B.n209 B.n98 256.663
R278 B.n203 B.n98 256.663
R279 B.n201 B.n98 256.663
R280 B.n195 B.n98 256.663
R281 B.n193 B.n98 256.663
R282 B.n187 B.n98 256.663
R283 B.n185 B.n98 256.663
R284 B.n178 B.n98 256.663
R285 B.n176 B.n98 256.663
R286 B.n170 B.n98 256.663
R287 B.n168 B.n98 256.663
R288 B.n161 B.n98 256.663
R289 B.n159 B.n98 256.663
R290 B.n153 B.n98 256.663
R291 B.n151 B.n98 256.663
R292 B.n145 B.n98 256.663
R293 B.n143 B.n98 256.663
R294 B.n137 B.n98 256.663
R295 B.n135 B.n98 256.663
R296 B.n129 B.n98 256.663
R297 B.n127 B.n98 256.663
R298 B.n221 B.n93 163.367
R299 B.n229 B.n93 163.367
R300 B.n229 B.n91 163.367
R301 B.n233 B.n91 163.367
R302 B.n233 B.n85 163.367
R303 B.n241 B.n85 163.367
R304 B.n241 B.n83 163.367
R305 B.n245 B.n83 163.367
R306 B.n245 B.n77 163.367
R307 B.n254 B.n77 163.367
R308 B.n254 B.n75 163.367
R309 B.n258 B.n75 163.367
R310 B.n258 B.n70 163.367
R311 B.n267 B.n70 163.367
R312 B.n267 B.n68 163.367
R313 B.n271 B.n68 163.367
R314 B.n271 B.n2 163.367
R315 B.n431 B.n2 163.367
R316 B.n431 B.n3 163.367
R317 B.n427 B.n3 163.367
R318 B.n427 B.n9 163.367
R319 B.n423 B.n9 163.367
R320 B.n423 B.n11 163.367
R321 B.n419 B.n11 163.367
R322 B.n419 B.n15 163.367
R323 B.n415 B.n15 163.367
R324 B.n415 B.n17 163.367
R325 B.n411 B.n17 163.367
R326 B.n411 B.n23 163.367
R327 B.n407 B.n23 163.367
R328 B.n407 B.n25 163.367
R329 B.n403 B.n25 163.367
R330 B.n403 B.n30 163.367
R331 B.n399 B.n30 163.367
R332 B.n399 B.n32 163.367
R333 B.n395 B.n32 163.367
R334 B.n217 B.n215 163.367
R335 B.n215 B.n214 163.367
R336 B.n211 B.n210 163.367
R337 B.n208 B.n103 163.367
R338 B.n204 B.n202 163.367
R339 B.n200 B.n105 163.367
R340 B.n196 B.n194 163.367
R341 B.n192 B.n107 163.367
R342 B.n188 B.n186 163.367
R343 B.n184 B.n109 163.367
R344 B.n179 B.n177 163.367
R345 B.n175 B.n113 163.367
R346 B.n171 B.n169 163.367
R347 B.n167 B.n115 163.367
R348 B.n162 B.n160 163.367
R349 B.n158 B.n119 163.367
R350 B.n154 B.n152 163.367
R351 B.n150 B.n121 163.367
R352 B.n146 B.n144 163.367
R353 B.n142 B.n123 163.367
R354 B.n138 B.n136 163.367
R355 B.n134 B.n125 163.367
R356 B.n130 B.n128 163.367
R357 B.n223 B.n95 163.367
R358 B.n227 B.n95 163.367
R359 B.n227 B.n88 163.367
R360 B.n235 B.n88 163.367
R361 B.n235 B.n86 163.367
R362 B.n239 B.n86 163.367
R363 B.n239 B.n81 163.367
R364 B.n247 B.n81 163.367
R365 B.n247 B.n79 163.367
R366 B.n251 B.n79 163.367
R367 B.n251 B.n74 163.367
R368 B.n260 B.n74 163.367
R369 B.n260 B.n72 163.367
R370 B.n265 B.n72 163.367
R371 B.n265 B.n66 163.367
R372 B.n273 B.n66 163.367
R373 B.n274 B.n273 163.367
R374 B.n274 B.n5 163.367
R375 B.n6 B.n5 163.367
R376 B.n7 B.n6 163.367
R377 B.n279 B.n7 163.367
R378 B.n279 B.n12 163.367
R379 B.n13 B.n12 163.367
R380 B.n14 B.n13 163.367
R381 B.n284 B.n14 163.367
R382 B.n284 B.n19 163.367
R383 B.n20 B.n19 163.367
R384 B.n21 B.n20 163.367
R385 B.n289 B.n21 163.367
R386 B.n289 B.n26 163.367
R387 B.n27 B.n26 163.367
R388 B.n28 B.n27 163.367
R389 B.n294 B.n28 163.367
R390 B.n294 B.n33 163.367
R391 B.n34 B.n33 163.367
R392 B.n35 B.n34 163.367
R393 B.n391 B.n389 163.367
R394 B.n387 B.n39 163.367
R395 B.n383 B.n381 163.367
R396 B.n379 B.n41 163.367
R397 B.n375 B.n373 163.367
R398 B.n371 B.n43 163.367
R399 B.n367 B.n365 163.367
R400 B.n363 B.n45 163.367
R401 B.n359 B.n357 163.367
R402 B.n355 B.n47 163.367
R403 B.n351 B.n349 163.367
R404 B.n347 B.n52 163.367
R405 B.n343 B.n341 163.367
R406 B.n339 B.n54 163.367
R407 B.n334 B.n332 163.367
R408 B.n330 B.n58 163.367
R409 B.n326 B.n324 163.367
R410 B.n322 B.n60 163.367
R411 B.n318 B.n316 163.367
R412 B.n314 B.n62 163.367
R413 B.n310 B.n308 163.367
R414 B.n306 B.n64 163.367
R415 B.n302 B.n300 163.367
R416 B.n222 B.n98 128.19
R417 B.n396 B.n36 128.19
R418 B.n116 B.t7 95.7036
R419 B.n55 B.t10 95.7036
R420 B.n110 B.t17 95.6998
R421 B.n48 B.t13 95.6998
R422 B.n222 B.n94 78.5307
R423 B.n228 B.n94 78.5307
R424 B.n228 B.n89 78.5307
R425 B.n234 B.n89 78.5307
R426 B.n234 B.n90 78.5307
R427 B.n240 B.n82 78.5307
R428 B.n246 B.n82 78.5307
R429 B.n246 B.n78 78.5307
R430 B.n253 B.n78 78.5307
R431 B.n253 B.n252 78.5307
R432 B.n259 B.n71 78.5307
R433 B.n266 B.n71 78.5307
R434 B.n272 B.n67 78.5307
R435 B.n272 B.n4 78.5307
R436 B.n430 B.n4 78.5307
R437 B.n430 B.n429 78.5307
R438 B.n429 B.n428 78.5307
R439 B.n428 B.n8 78.5307
R440 B.n422 B.n421 78.5307
R441 B.n421 B.n420 78.5307
R442 B.n414 B.n18 78.5307
R443 B.n414 B.n413 78.5307
R444 B.n413 B.n412 78.5307
R445 B.n412 B.n22 78.5307
R446 B.n406 B.n22 78.5307
R447 B.n405 B.n404 78.5307
R448 B.n404 B.n29 78.5307
R449 B.n398 B.n29 78.5307
R450 B.n398 B.n397 78.5307
R451 B.n397 B.n396 78.5307
R452 B.n117 B.t6 74.3703
R453 B.n56 B.t11 74.3703
R454 B.n111 B.t16 74.3664
R455 B.n49 B.t14 74.3664
R456 B.n216 B.n99 71.676
R457 B.n214 B.n101 71.676
R458 B.n210 B.n209 71.676
R459 B.n203 B.n103 71.676
R460 B.n202 B.n201 71.676
R461 B.n195 B.n105 71.676
R462 B.n194 B.n193 71.676
R463 B.n187 B.n107 71.676
R464 B.n186 B.n185 71.676
R465 B.n178 B.n109 71.676
R466 B.n177 B.n176 71.676
R467 B.n170 B.n113 71.676
R468 B.n169 B.n168 71.676
R469 B.n161 B.n115 71.676
R470 B.n160 B.n159 71.676
R471 B.n153 B.n119 71.676
R472 B.n152 B.n151 71.676
R473 B.n145 B.n121 71.676
R474 B.n144 B.n143 71.676
R475 B.n137 B.n123 71.676
R476 B.n136 B.n135 71.676
R477 B.n129 B.n125 71.676
R478 B.n128 B.n127 71.676
R479 B.n390 B.n37 71.676
R480 B.n389 B.n388 71.676
R481 B.n382 B.n39 71.676
R482 B.n381 B.n380 71.676
R483 B.n374 B.n41 71.676
R484 B.n373 B.n372 71.676
R485 B.n366 B.n43 71.676
R486 B.n365 B.n364 71.676
R487 B.n358 B.n45 71.676
R488 B.n357 B.n356 71.676
R489 B.n350 B.n47 71.676
R490 B.n349 B.n348 71.676
R491 B.n342 B.n52 71.676
R492 B.n341 B.n340 71.676
R493 B.n333 B.n54 71.676
R494 B.n332 B.n331 71.676
R495 B.n325 B.n58 71.676
R496 B.n324 B.n323 71.676
R497 B.n317 B.n60 71.676
R498 B.n316 B.n315 71.676
R499 B.n309 B.n62 71.676
R500 B.n308 B.n307 71.676
R501 B.n301 B.n64 71.676
R502 B.n302 B.n301 71.676
R503 B.n307 B.n306 71.676
R504 B.n310 B.n309 71.676
R505 B.n315 B.n314 71.676
R506 B.n318 B.n317 71.676
R507 B.n323 B.n322 71.676
R508 B.n326 B.n325 71.676
R509 B.n331 B.n330 71.676
R510 B.n334 B.n333 71.676
R511 B.n340 B.n339 71.676
R512 B.n343 B.n342 71.676
R513 B.n348 B.n347 71.676
R514 B.n351 B.n350 71.676
R515 B.n356 B.n355 71.676
R516 B.n359 B.n358 71.676
R517 B.n364 B.n363 71.676
R518 B.n367 B.n366 71.676
R519 B.n372 B.n371 71.676
R520 B.n375 B.n374 71.676
R521 B.n380 B.n379 71.676
R522 B.n383 B.n382 71.676
R523 B.n388 B.n387 71.676
R524 B.n391 B.n390 71.676
R525 B.n217 B.n216 71.676
R526 B.n211 B.n101 71.676
R527 B.n209 B.n208 71.676
R528 B.n204 B.n203 71.676
R529 B.n201 B.n200 71.676
R530 B.n196 B.n195 71.676
R531 B.n193 B.n192 71.676
R532 B.n188 B.n187 71.676
R533 B.n185 B.n184 71.676
R534 B.n179 B.n178 71.676
R535 B.n176 B.n175 71.676
R536 B.n171 B.n170 71.676
R537 B.n168 B.n167 71.676
R538 B.n162 B.n161 71.676
R539 B.n159 B.n158 71.676
R540 B.n154 B.n153 71.676
R541 B.n151 B.n150 71.676
R542 B.n146 B.n145 71.676
R543 B.n143 B.n142 71.676
R544 B.n138 B.n137 71.676
R545 B.n135 B.n134 71.676
R546 B.n130 B.n129 71.676
R547 B.n127 B.n97 71.676
R548 B.n240 B.t5 70.4467
R549 B.n406 B.t9 70.4467
R550 B.n266 B.t1 61.2078
R551 B.n422 B.t0 61.2078
R552 B.n164 B.n117 59.5399
R553 B.n182 B.n111 59.5399
R554 B.n50 B.n49 59.5399
R555 B.n337 B.n56 59.5399
R556 B.n252 B.t3 42.7302
R557 B.n18 B.t2 42.7302
R558 B.n259 B.t3 35.801
R559 B.n420 B.t2 35.801
R560 B.n394 B.n393 31.6883
R561 B.n299 B.n298 31.6883
R562 B.n224 B.n96 31.6883
R563 B.n220 B.n219 31.6883
R564 B.n117 B.n116 21.3338
R565 B.n111 B.n110 21.3338
R566 B.n49 B.n48 21.3338
R567 B.n56 B.n55 21.3338
R568 B B.n432 18.0485
R569 B.t1 B.n67 17.3233
R570 B.t0 B.n8 17.3233
R571 B.n393 B.n392 10.6151
R572 B.n392 B.n38 10.6151
R573 B.n386 B.n38 10.6151
R574 B.n386 B.n385 10.6151
R575 B.n385 B.n384 10.6151
R576 B.n384 B.n40 10.6151
R577 B.n378 B.n40 10.6151
R578 B.n378 B.n377 10.6151
R579 B.n377 B.n376 10.6151
R580 B.n376 B.n42 10.6151
R581 B.n370 B.n42 10.6151
R582 B.n370 B.n369 10.6151
R583 B.n369 B.n368 10.6151
R584 B.n368 B.n44 10.6151
R585 B.n362 B.n44 10.6151
R586 B.n362 B.n361 10.6151
R587 B.n361 B.n360 10.6151
R588 B.n360 B.n46 10.6151
R589 B.n354 B.n353 10.6151
R590 B.n353 B.n352 10.6151
R591 B.n352 B.n51 10.6151
R592 B.n346 B.n51 10.6151
R593 B.n346 B.n345 10.6151
R594 B.n345 B.n344 10.6151
R595 B.n344 B.n53 10.6151
R596 B.n338 B.n53 10.6151
R597 B.n336 B.n335 10.6151
R598 B.n335 B.n57 10.6151
R599 B.n329 B.n57 10.6151
R600 B.n329 B.n328 10.6151
R601 B.n328 B.n327 10.6151
R602 B.n327 B.n59 10.6151
R603 B.n321 B.n59 10.6151
R604 B.n321 B.n320 10.6151
R605 B.n320 B.n319 10.6151
R606 B.n319 B.n61 10.6151
R607 B.n313 B.n61 10.6151
R608 B.n313 B.n312 10.6151
R609 B.n312 B.n311 10.6151
R610 B.n311 B.n63 10.6151
R611 B.n305 B.n63 10.6151
R612 B.n305 B.n304 10.6151
R613 B.n304 B.n303 10.6151
R614 B.n303 B.n299 10.6151
R615 B.n225 B.n224 10.6151
R616 B.n226 B.n225 10.6151
R617 B.n226 B.n87 10.6151
R618 B.n236 B.n87 10.6151
R619 B.n237 B.n236 10.6151
R620 B.n238 B.n237 10.6151
R621 B.n238 B.n80 10.6151
R622 B.n248 B.n80 10.6151
R623 B.n249 B.n248 10.6151
R624 B.n250 B.n249 10.6151
R625 B.n250 B.n73 10.6151
R626 B.n261 B.n73 10.6151
R627 B.n262 B.n261 10.6151
R628 B.n264 B.n262 10.6151
R629 B.n264 B.n263 10.6151
R630 B.n263 B.n65 10.6151
R631 B.n275 B.n65 10.6151
R632 B.n276 B.n275 10.6151
R633 B.n277 B.n276 10.6151
R634 B.n278 B.n277 10.6151
R635 B.n280 B.n278 10.6151
R636 B.n281 B.n280 10.6151
R637 B.n282 B.n281 10.6151
R638 B.n283 B.n282 10.6151
R639 B.n285 B.n283 10.6151
R640 B.n286 B.n285 10.6151
R641 B.n287 B.n286 10.6151
R642 B.n288 B.n287 10.6151
R643 B.n290 B.n288 10.6151
R644 B.n291 B.n290 10.6151
R645 B.n292 B.n291 10.6151
R646 B.n293 B.n292 10.6151
R647 B.n295 B.n293 10.6151
R648 B.n296 B.n295 10.6151
R649 B.n297 B.n296 10.6151
R650 B.n298 B.n297 10.6151
R651 B.n219 B.n218 10.6151
R652 B.n218 B.n100 10.6151
R653 B.n213 B.n100 10.6151
R654 B.n213 B.n212 10.6151
R655 B.n212 B.n102 10.6151
R656 B.n207 B.n102 10.6151
R657 B.n207 B.n206 10.6151
R658 B.n206 B.n205 10.6151
R659 B.n205 B.n104 10.6151
R660 B.n199 B.n104 10.6151
R661 B.n199 B.n198 10.6151
R662 B.n198 B.n197 10.6151
R663 B.n197 B.n106 10.6151
R664 B.n191 B.n106 10.6151
R665 B.n191 B.n190 10.6151
R666 B.n190 B.n189 10.6151
R667 B.n189 B.n108 10.6151
R668 B.n183 B.n108 10.6151
R669 B.n181 B.n180 10.6151
R670 B.n180 B.n112 10.6151
R671 B.n174 B.n112 10.6151
R672 B.n174 B.n173 10.6151
R673 B.n173 B.n172 10.6151
R674 B.n172 B.n114 10.6151
R675 B.n166 B.n114 10.6151
R676 B.n166 B.n165 10.6151
R677 B.n163 B.n118 10.6151
R678 B.n157 B.n118 10.6151
R679 B.n157 B.n156 10.6151
R680 B.n156 B.n155 10.6151
R681 B.n155 B.n120 10.6151
R682 B.n149 B.n120 10.6151
R683 B.n149 B.n148 10.6151
R684 B.n148 B.n147 10.6151
R685 B.n147 B.n122 10.6151
R686 B.n141 B.n122 10.6151
R687 B.n141 B.n140 10.6151
R688 B.n140 B.n139 10.6151
R689 B.n139 B.n124 10.6151
R690 B.n133 B.n124 10.6151
R691 B.n133 B.n132 10.6151
R692 B.n132 B.n131 10.6151
R693 B.n131 B.n126 10.6151
R694 B.n126 B.n96 10.6151
R695 B.n220 B.n92 10.6151
R696 B.n230 B.n92 10.6151
R697 B.n231 B.n230 10.6151
R698 B.n232 B.n231 10.6151
R699 B.n232 B.n84 10.6151
R700 B.n242 B.n84 10.6151
R701 B.n243 B.n242 10.6151
R702 B.n244 B.n243 10.6151
R703 B.n244 B.n76 10.6151
R704 B.n255 B.n76 10.6151
R705 B.n256 B.n255 10.6151
R706 B.n257 B.n256 10.6151
R707 B.n257 B.n69 10.6151
R708 B.n268 B.n69 10.6151
R709 B.n269 B.n268 10.6151
R710 B.n270 B.n269 10.6151
R711 B.n270 B.n0 10.6151
R712 B.n426 B.n1 10.6151
R713 B.n426 B.n425 10.6151
R714 B.n425 B.n424 10.6151
R715 B.n424 B.n10 10.6151
R716 B.n418 B.n10 10.6151
R717 B.n418 B.n417 10.6151
R718 B.n417 B.n416 10.6151
R719 B.n416 B.n16 10.6151
R720 B.n410 B.n16 10.6151
R721 B.n410 B.n409 10.6151
R722 B.n409 B.n408 10.6151
R723 B.n408 B.n24 10.6151
R724 B.n402 B.n24 10.6151
R725 B.n402 B.n401 10.6151
R726 B.n401 B.n400 10.6151
R727 B.n400 B.n31 10.6151
R728 B.n394 B.n31 10.6151
R729 B.n90 B.t5 8.08449
R730 B.t9 B.n405 8.08449
R731 B.n354 B.n50 6.5566
R732 B.n338 B.n337 6.5566
R733 B.n182 B.n181 6.5566
R734 B.n165 B.n164 6.5566
R735 B.n50 B.n46 4.05904
R736 B.n337 B.n336 4.05904
R737 B.n183 B.n182 4.05904
R738 B.n164 B.n163 4.05904
R739 B.n432 B.n0 2.81026
R740 B.n432 B.n1 2.81026
R741 VP.n1 VP.t1 205.346
R742 VP.n1 VP.t2 205.297
R743 VP.n3 VP.t0 184.35
R744 VP.n5 VP.t3 184.35
R745 VP.n6 VP.n5 161.3
R746 VP.n4 VP.n0 161.3
R747 VP.n3 VP.n2 161.3
R748 VP.n2 VP.n1 79.4651
R749 VP.n4 VP.n3 24.1005
R750 VP.n5 VP.n4 24.1005
R751 VP.n2 VP.n0 0.189894
R752 VP.n6 VP.n0 0.189894
R753 VP VP.n6 0.0516364
R754 VDD1 VDD1.n1 103.636
R755 VDD1 VDD1.n0 72.9462
R756 VDD1.n0 VDD1.t0 4.65932
R757 VDD1.n0 VDD1.t2 4.65932
R758 VDD1.n1 VDD1.t3 4.65932
R759 VDD1.n1 VDD1.t1 4.65932
R760 VTAIL.n5 VTAIL.t6 60.8682
R761 VTAIL.n4 VTAIL.t2 60.8682
R762 VTAIL.n3 VTAIL.t3 60.8682
R763 VTAIL.n7 VTAIL.t0 60.868
R764 VTAIL.n0 VTAIL.t1 60.868
R765 VTAIL.n1 VTAIL.t4 60.868
R766 VTAIL.n2 VTAIL.t7 60.868
R767 VTAIL.n6 VTAIL.t5 60.868
R768 VTAIL.n7 VTAIL.n6 16.9789
R769 VTAIL.n3 VTAIL.n2 16.9789
R770 VTAIL.n4 VTAIL.n3 0.948776
R771 VTAIL.n6 VTAIL.n5 0.948776
R772 VTAIL.n2 VTAIL.n1 0.948776
R773 VTAIL VTAIL.n0 0.532828
R774 VTAIL.n5 VTAIL.n4 0.470328
R775 VTAIL.n1 VTAIL.n0 0.470328
R776 VTAIL VTAIL.n7 0.416448
R777 VN.n0 VN.t3 205.346
R778 VN.n1 VN.t2 205.346
R779 VN.n0 VN.t0 205.297
R780 VN.n1 VN.t1 205.297
R781 VN VN.n1 79.8458
R782 VN VN.n0 44.7132
R783 VDD2.n2 VDD2.n0 103.112
R784 VDD2.n2 VDD2.n1 72.888
R785 VDD2.n1 VDD2.t2 4.65932
R786 VDD2.n1 VDD2.t1 4.65932
R787 VDD2.n0 VDD2.t0 4.65932
R788 VDD2.n0 VDD2.t3 4.65932
R789 VDD2 VDD2.n2 0.0586897
C0 VP VDD1 1.48826f
C1 VTAIL VN 1.3519f
C2 VDD2 VN 1.35802f
C3 VDD1 VN 0.151274f
C4 VTAIL VDD2 3.34044f
C5 VTAIL VDD1 3.2985f
C6 VDD2 VDD1 0.582539f
C7 VP VN 3.44241f
C8 VTAIL VP 1.36601f
C9 VP VDD2 0.28211f
C10 VDD2 B 2.096888f
C11 VDD1 B 4.00312f
C12 VTAIL B 4.288809f
C13 VN B 5.92598f
C14 VP B 4.407461f
C15 VDD2.t0 B 0.06482f
C16 VDD2.t3 B 0.06482f
C17 VDD2.n0 B 0.735841f
C18 VDD2.t2 B 0.06482f
C19 VDD2.t1 B 0.06482f
C20 VDD2.n1 B 0.514838f
C21 VDD2.n2 B 1.72691f
C22 VN.t3 B 0.277479f
C23 VN.t0 B 0.277438f
C24 VN.n0 B 0.243901f
C25 VN.t2 B 0.277479f
C26 VN.t1 B 0.277438f
C27 VN.n1 B 0.634264f
C28 VTAIL.t1 B 0.427385f
C29 VTAIL.n0 B 0.19517f
C30 VTAIL.t4 B 0.427385f
C31 VTAIL.n1 B 0.213496f
C32 VTAIL.t7 B 0.427385f
C33 VTAIL.n2 B 0.581734f
C34 VTAIL.t3 B 0.427386f
C35 VTAIL.n3 B 0.581733f
C36 VTAIL.t2 B 0.427386f
C37 VTAIL.n4 B 0.213494f
C38 VTAIL.t6 B 0.427386f
C39 VTAIL.n5 B 0.213494f
C40 VTAIL.t5 B 0.427385f
C41 VTAIL.n6 B 0.581734f
C42 VTAIL.t0 B 0.427385f
C43 VTAIL.n7 B 0.558281f
C44 VDD1.t0 B 0.063449f
C45 VDD1.t2 B 0.063449f
C46 VDD1.n0 B 0.504125f
C47 VDD1.t3 B 0.063449f
C48 VDD1.t1 B 0.063449f
C49 VDD1.n1 B 0.73447f
C50 VP.n0 B 0.027695f
C51 VP.t2 B 0.280615f
C52 VP.t1 B 0.280656f
C53 VP.n1 B 0.63106f
C54 VP.n2 B 1.33829f
C55 VP.t0 B 0.266744f
C56 VP.n3 B 0.133951f
C57 VP.n4 B 0.006285f
C58 VP.t3 B 0.266744f
C59 VP.n5 B 0.133951f
C60 VP.n6 B 0.021463f
.ends

