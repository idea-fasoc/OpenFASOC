* NGSPICE file created from diff_pair_sample_1252.ext - technology: sky130A

.subckt diff_pair_sample_1252 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3170_n1974# sky130_fd_pr__pfet_01v8 ad=1.9617 pd=10.84 as=0 ps=0 w=5.03 l=1.87
X1 VDD1.t7 VP.t0 VTAIL.t10 w_n3170_n1974# sky130_fd_pr__pfet_01v8 ad=0.82995 pd=5.36 as=1.9617 ps=10.84 w=5.03 l=1.87
X2 VTAIL.t4 VP.t1 VDD1.t6 w_n3170_n1974# sky130_fd_pr__pfet_01v8 ad=0.82995 pd=5.36 as=0.82995 ps=5.36 w=5.03 l=1.87
X3 VTAIL.t12 VN.t0 VDD2.t7 w_n3170_n1974# sky130_fd_pr__pfet_01v8 ad=1.9617 pd=10.84 as=0.82995 ps=5.36 w=5.03 l=1.87
X4 VDD1.t5 VP.t2 VTAIL.t5 w_n3170_n1974# sky130_fd_pr__pfet_01v8 ad=0.82995 pd=5.36 as=1.9617 ps=10.84 w=5.03 l=1.87
X5 VDD2.t6 VN.t1 VTAIL.t13 w_n3170_n1974# sky130_fd_pr__pfet_01v8 ad=0.82995 pd=5.36 as=0.82995 ps=5.36 w=5.03 l=1.87
X6 VTAIL.t6 VP.t3 VDD1.t4 w_n3170_n1974# sky130_fd_pr__pfet_01v8 ad=1.9617 pd=10.84 as=0.82995 ps=5.36 w=5.03 l=1.87
X7 B.t8 B.t6 B.t7 w_n3170_n1974# sky130_fd_pr__pfet_01v8 ad=1.9617 pd=10.84 as=0 ps=0 w=5.03 l=1.87
X8 VTAIL.t15 VN.t2 VDD2.t5 w_n3170_n1974# sky130_fd_pr__pfet_01v8 ad=0.82995 pd=5.36 as=0.82995 ps=5.36 w=5.03 l=1.87
X9 B.t5 B.t3 B.t4 w_n3170_n1974# sky130_fd_pr__pfet_01v8 ad=1.9617 pd=10.84 as=0 ps=0 w=5.03 l=1.87
X10 VDD2.t4 VN.t3 VTAIL.t14 w_n3170_n1974# sky130_fd_pr__pfet_01v8 ad=0.82995 pd=5.36 as=0.82995 ps=5.36 w=5.03 l=1.87
X11 VDD1.t3 VP.t4 VTAIL.t8 w_n3170_n1974# sky130_fd_pr__pfet_01v8 ad=0.82995 pd=5.36 as=0.82995 ps=5.36 w=5.03 l=1.87
X12 VDD2.t3 VN.t4 VTAIL.t11 w_n3170_n1974# sky130_fd_pr__pfet_01v8 ad=0.82995 pd=5.36 as=1.9617 ps=10.84 w=5.03 l=1.87
X13 B.t2 B.t0 B.t1 w_n3170_n1974# sky130_fd_pr__pfet_01v8 ad=1.9617 pd=10.84 as=0 ps=0 w=5.03 l=1.87
X14 VTAIL.t1 VN.t5 VDD2.t2 w_n3170_n1974# sky130_fd_pr__pfet_01v8 ad=1.9617 pd=10.84 as=0.82995 ps=5.36 w=5.03 l=1.87
X15 VDD1.t2 VP.t5 VTAIL.t3 w_n3170_n1974# sky130_fd_pr__pfet_01v8 ad=0.82995 pd=5.36 as=0.82995 ps=5.36 w=5.03 l=1.87
X16 VTAIL.t9 VP.t6 VDD1.t1 w_n3170_n1974# sky130_fd_pr__pfet_01v8 ad=1.9617 pd=10.84 as=0.82995 ps=5.36 w=5.03 l=1.87
X17 VTAIL.t7 VP.t7 VDD1.t0 w_n3170_n1974# sky130_fd_pr__pfet_01v8 ad=0.82995 pd=5.36 as=0.82995 ps=5.36 w=5.03 l=1.87
X18 VDD2.t1 VN.t6 VTAIL.t0 w_n3170_n1974# sky130_fd_pr__pfet_01v8 ad=0.82995 pd=5.36 as=1.9617 ps=10.84 w=5.03 l=1.87
X19 VTAIL.t2 VN.t7 VDD2.t0 w_n3170_n1974# sky130_fd_pr__pfet_01v8 ad=0.82995 pd=5.36 as=0.82995 ps=5.36 w=5.03 l=1.87
R0 B.n281 B.n94 585
R1 B.n280 B.n279 585
R2 B.n278 B.n95 585
R3 B.n277 B.n276 585
R4 B.n275 B.n96 585
R5 B.n274 B.n273 585
R6 B.n272 B.n97 585
R7 B.n271 B.n270 585
R8 B.n269 B.n98 585
R9 B.n268 B.n267 585
R10 B.n266 B.n99 585
R11 B.n265 B.n264 585
R12 B.n263 B.n100 585
R13 B.n262 B.n261 585
R14 B.n260 B.n101 585
R15 B.n259 B.n258 585
R16 B.n257 B.n102 585
R17 B.n256 B.n255 585
R18 B.n254 B.n103 585
R19 B.n253 B.n252 585
R20 B.n251 B.n104 585
R21 B.n249 B.n248 585
R22 B.n247 B.n107 585
R23 B.n246 B.n245 585
R24 B.n244 B.n108 585
R25 B.n243 B.n242 585
R26 B.n241 B.n109 585
R27 B.n240 B.n239 585
R28 B.n238 B.n110 585
R29 B.n237 B.n236 585
R30 B.n235 B.n111 585
R31 B.n234 B.n233 585
R32 B.n229 B.n112 585
R33 B.n228 B.n227 585
R34 B.n226 B.n113 585
R35 B.n225 B.n224 585
R36 B.n223 B.n114 585
R37 B.n222 B.n221 585
R38 B.n220 B.n115 585
R39 B.n219 B.n218 585
R40 B.n217 B.n116 585
R41 B.n216 B.n215 585
R42 B.n214 B.n117 585
R43 B.n213 B.n212 585
R44 B.n211 B.n118 585
R45 B.n210 B.n209 585
R46 B.n208 B.n119 585
R47 B.n207 B.n206 585
R48 B.n205 B.n120 585
R49 B.n204 B.n203 585
R50 B.n202 B.n121 585
R51 B.n201 B.n200 585
R52 B.n283 B.n282 585
R53 B.n284 B.n93 585
R54 B.n286 B.n285 585
R55 B.n287 B.n92 585
R56 B.n289 B.n288 585
R57 B.n290 B.n91 585
R58 B.n292 B.n291 585
R59 B.n293 B.n90 585
R60 B.n295 B.n294 585
R61 B.n296 B.n89 585
R62 B.n298 B.n297 585
R63 B.n299 B.n88 585
R64 B.n301 B.n300 585
R65 B.n302 B.n87 585
R66 B.n304 B.n303 585
R67 B.n305 B.n86 585
R68 B.n307 B.n306 585
R69 B.n308 B.n85 585
R70 B.n310 B.n309 585
R71 B.n311 B.n84 585
R72 B.n313 B.n312 585
R73 B.n314 B.n83 585
R74 B.n316 B.n315 585
R75 B.n317 B.n82 585
R76 B.n319 B.n318 585
R77 B.n320 B.n81 585
R78 B.n322 B.n321 585
R79 B.n323 B.n80 585
R80 B.n325 B.n324 585
R81 B.n326 B.n79 585
R82 B.n328 B.n327 585
R83 B.n329 B.n78 585
R84 B.n331 B.n330 585
R85 B.n332 B.n77 585
R86 B.n334 B.n333 585
R87 B.n335 B.n76 585
R88 B.n337 B.n336 585
R89 B.n338 B.n75 585
R90 B.n340 B.n339 585
R91 B.n341 B.n74 585
R92 B.n343 B.n342 585
R93 B.n344 B.n73 585
R94 B.n346 B.n345 585
R95 B.n347 B.n72 585
R96 B.n349 B.n348 585
R97 B.n350 B.n71 585
R98 B.n352 B.n351 585
R99 B.n353 B.n70 585
R100 B.n355 B.n354 585
R101 B.n356 B.n69 585
R102 B.n358 B.n357 585
R103 B.n359 B.n68 585
R104 B.n361 B.n360 585
R105 B.n362 B.n67 585
R106 B.n364 B.n363 585
R107 B.n365 B.n66 585
R108 B.n367 B.n366 585
R109 B.n368 B.n65 585
R110 B.n370 B.n369 585
R111 B.n371 B.n64 585
R112 B.n373 B.n372 585
R113 B.n374 B.n63 585
R114 B.n376 B.n375 585
R115 B.n377 B.n62 585
R116 B.n379 B.n378 585
R117 B.n380 B.n61 585
R118 B.n382 B.n381 585
R119 B.n383 B.n60 585
R120 B.n385 B.n384 585
R121 B.n386 B.n59 585
R122 B.n388 B.n387 585
R123 B.n389 B.n58 585
R124 B.n391 B.n390 585
R125 B.n392 B.n57 585
R126 B.n394 B.n393 585
R127 B.n395 B.n56 585
R128 B.n397 B.n396 585
R129 B.n398 B.n55 585
R130 B.n400 B.n399 585
R131 B.n401 B.n54 585
R132 B.n403 B.n402 585
R133 B.n404 B.n53 585
R134 B.n483 B.n22 585
R135 B.n482 B.n481 585
R136 B.n480 B.n23 585
R137 B.n479 B.n478 585
R138 B.n477 B.n24 585
R139 B.n476 B.n475 585
R140 B.n474 B.n25 585
R141 B.n473 B.n472 585
R142 B.n471 B.n26 585
R143 B.n470 B.n469 585
R144 B.n468 B.n27 585
R145 B.n467 B.n466 585
R146 B.n465 B.n28 585
R147 B.n464 B.n463 585
R148 B.n462 B.n29 585
R149 B.n461 B.n460 585
R150 B.n459 B.n30 585
R151 B.n458 B.n457 585
R152 B.n456 B.n31 585
R153 B.n455 B.n454 585
R154 B.n453 B.n32 585
R155 B.n452 B.n451 585
R156 B.n450 B.n33 585
R157 B.n449 B.n448 585
R158 B.n447 B.n37 585
R159 B.n446 B.n445 585
R160 B.n444 B.n38 585
R161 B.n443 B.n442 585
R162 B.n441 B.n39 585
R163 B.n440 B.n439 585
R164 B.n438 B.n40 585
R165 B.n436 B.n435 585
R166 B.n434 B.n43 585
R167 B.n433 B.n432 585
R168 B.n431 B.n44 585
R169 B.n430 B.n429 585
R170 B.n428 B.n45 585
R171 B.n427 B.n426 585
R172 B.n425 B.n46 585
R173 B.n424 B.n423 585
R174 B.n422 B.n47 585
R175 B.n421 B.n420 585
R176 B.n419 B.n48 585
R177 B.n418 B.n417 585
R178 B.n416 B.n49 585
R179 B.n415 B.n414 585
R180 B.n413 B.n50 585
R181 B.n412 B.n411 585
R182 B.n410 B.n51 585
R183 B.n409 B.n408 585
R184 B.n407 B.n52 585
R185 B.n406 B.n405 585
R186 B.n485 B.n484 585
R187 B.n486 B.n21 585
R188 B.n488 B.n487 585
R189 B.n489 B.n20 585
R190 B.n491 B.n490 585
R191 B.n492 B.n19 585
R192 B.n494 B.n493 585
R193 B.n495 B.n18 585
R194 B.n497 B.n496 585
R195 B.n498 B.n17 585
R196 B.n500 B.n499 585
R197 B.n501 B.n16 585
R198 B.n503 B.n502 585
R199 B.n504 B.n15 585
R200 B.n506 B.n505 585
R201 B.n507 B.n14 585
R202 B.n509 B.n508 585
R203 B.n510 B.n13 585
R204 B.n512 B.n511 585
R205 B.n513 B.n12 585
R206 B.n515 B.n514 585
R207 B.n516 B.n11 585
R208 B.n518 B.n517 585
R209 B.n519 B.n10 585
R210 B.n521 B.n520 585
R211 B.n522 B.n9 585
R212 B.n524 B.n523 585
R213 B.n525 B.n8 585
R214 B.n527 B.n526 585
R215 B.n528 B.n7 585
R216 B.n530 B.n529 585
R217 B.n531 B.n6 585
R218 B.n533 B.n532 585
R219 B.n534 B.n5 585
R220 B.n536 B.n535 585
R221 B.n537 B.n4 585
R222 B.n539 B.n538 585
R223 B.n540 B.n3 585
R224 B.n542 B.n541 585
R225 B.n543 B.n0 585
R226 B.n2 B.n1 585
R227 B.n142 B.n141 585
R228 B.n144 B.n143 585
R229 B.n145 B.n140 585
R230 B.n147 B.n146 585
R231 B.n148 B.n139 585
R232 B.n150 B.n149 585
R233 B.n151 B.n138 585
R234 B.n153 B.n152 585
R235 B.n154 B.n137 585
R236 B.n156 B.n155 585
R237 B.n157 B.n136 585
R238 B.n159 B.n158 585
R239 B.n160 B.n135 585
R240 B.n162 B.n161 585
R241 B.n163 B.n134 585
R242 B.n165 B.n164 585
R243 B.n166 B.n133 585
R244 B.n168 B.n167 585
R245 B.n169 B.n132 585
R246 B.n171 B.n170 585
R247 B.n172 B.n131 585
R248 B.n174 B.n173 585
R249 B.n175 B.n130 585
R250 B.n177 B.n176 585
R251 B.n178 B.n129 585
R252 B.n180 B.n179 585
R253 B.n181 B.n128 585
R254 B.n183 B.n182 585
R255 B.n184 B.n127 585
R256 B.n186 B.n185 585
R257 B.n187 B.n126 585
R258 B.n189 B.n188 585
R259 B.n190 B.n125 585
R260 B.n192 B.n191 585
R261 B.n193 B.n124 585
R262 B.n195 B.n194 585
R263 B.n196 B.n123 585
R264 B.n198 B.n197 585
R265 B.n199 B.n122 585
R266 B.n201 B.n122 478.086
R267 B.n283 B.n94 478.086
R268 B.n405 B.n404 478.086
R269 B.n484 B.n483 478.086
R270 B.n230 B.t6 271.421
R271 B.n105 B.t3 271.421
R272 B.n41 B.t9 271.421
R273 B.n34 B.t0 271.421
R274 B.n545 B.n544 256.663
R275 B.n544 B.n543 235.042
R276 B.n544 B.n2 235.042
R277 B.n202 B.n201 163.367
R278 B.n203 B.n202 163.367
R279 B.n203 B.n120 163.367
R280 B.n207 B.n120 163.367
R281 B.n208 B.n207 163.367
R282 B.n209 B.n208 163.367
R283 B.n209 B.n118 163.367
R284 B.n213 B.n118 163.367
R285 B.n214 B.n213 163.367
R286 B.n215 B.n214 163.367
R287 B.n215 B.n116 163.367
R288 B.n219 B.n116 163.367
R289 B.n220 B.n219 163.367
R290 B.n221 B.n220 163.367
R291 B.n221 B.n114 163.367
R292 B.n225 B.n114 163.367
R293 B.n226 B.n225 163.367
R294 B.n227 B.n226 163.367
R295 B.n227 B.n112 163.367
R296 B.n234 B.n112 163.367
R297 B.n235 B.n234 163.367
R298 B.n236 B.n235 163.367
R299 B.n236 B.n110 163.367
R300 B.n240 B.n110 163.367
R301 B.n241 B.n240 163.367
R302 B.n242 B.n241 163.367
R303 B.n242 B.n108 163.367
R304 B.n246 B.n108 163.367
R305 B.n247 B.n246 163.367
R306 B.n248 B.n247 163.367
R307 B.n248 B.n104 163.367
R308 B.n253 B.n104 163.367
R309 B.n254 B.n253 163.367
R310 B.n255 B.n254 163.367
R311 B.n255 B.n102 163.367
R312 B.n259 B.n102 163.367
R313 B.n260 B.n259 163.367
R314 B.n261 B.n260 163.367
R315 B.n261 B.n100 163.367
R316 B.n265 B.n100 163.367
R317 B.n266 B.n265 163.367
R318 B.n267 B.n266 163.367
R319 B.n267 B.n98 163.367
R320 B.n271 B.n98 163.367
R321 B.n272 B.n271 163.367
R322 B.n273 B.n272 163.367
R323 B.n273 B.n96 163.367
R324 B.n277 B.n96 163.367
R325 B.n278 B.n277 163.367
R326 B.n279 B.n278 163.367
R327 B.n279 B.n94 163.367
R328 B.n404 B.n403 163.367
R329 B.n403 B.n54 163.367
R330 B.n399 B.n54 163.367
R331 B.n399 B.n398 163.367
R332 B.n398 B.n397 163.367
R333 B.n397 B.n56 163.367
R334 B.n393 B.n56 163.367
R335 B.n393 B.n392 163.367
R336 B.n392 B.n391 163.367
R337 B.n391 B.n58 163.367
R338 B.n387 B.n58 163.367
R339 B.n387 B.n386 163.367
R340 B.n386 B.n385 163.367
R341 B.n385 B.n60 163.367
R342 B.n381 B.n60 163.367
R343 B.n381 B.n380 163.367
R344 B.n380 B.n379 163.367
R345 B.n379 B.n62 163.367
R346 B.n375 B.n62 163.367
R347 B.n375 B.n374 163.367
R348 B.n374 B.n373 163.367
R349 B.n373 B.n64 163.367
R350 B.n369 B.n64 163.367
R351 B.n369 B.n368 163.367
R352 B.n368 B.n367 163.367
R353 B.n367 B.n66 163.367
R354 B.n363 B.n66 163.367
R355 B.n363 B.n362 163.367
R356 B.n362 B.n361 163.367
R357 B.n361 B.n68 163.367
R358 B.n357 B.n68 163.367
R359 B.n357 B.n356 163.367
R360 B.n356 B.n355 163.367
R361 B.n355 B.n70 163.367
R362 B.n351 B.n70 163.367
R363 B.n351 B.n350 163.367
R364 B.n350 B.n349 163.367
R365 B.n349 B.n72 163.367
R366 B.n345 B.n72 163.367
R367 B.n345 B.n344 163.367
R368 B.n344 B.n343 163.367
R369 B.n343 B.n74 163.367
R370 B.n339 B.n74 163.367
R371 B.n339 B.n338 163.367
R372 B.n338 B.n337 163.367
R373 B.n337 B.n76 163.367
R374 B.n333 B.n76 163.367
R375 B.n333 B.n332 163.367
R376 B.n332 B.n331 163.367
R377 B.n331 B.n78 163.367
R378 B.n327 B.n78 163.367
R379 B.n327 B.n326 163.367
R380 B.n326 B.n325 163.367
R381 B.n325 B.n80 163.367
R382 B.n321 B.n80 163.367
R383 B.n321 B.n320 163.367
R384 B.n320 B.n319 163.367
R385 B.n319 B.n82 163.367
R386 B.n315 B.n82 163.367
R387 B.n315 B.n314 163.367
R388 B.n314 B.n313 163.367
R389 B.n313 B.n84 163.367
R390 B.n309 B.n84 163.367
R391 B.n309 B.n308 163.367
R392 B.n308 B.n307 163.367
R393 B.n307 B.n86 163.367
R394 B.n303 B.n86 163.367
R395 B.n303 B.n302 163.367
R396 B.n302 B.n301 163.367
R397 B.n301 B.n88 163.367
R398 B.n297 B.n88 163.367
R399 B.n297 B.n296 163.367
R400 B.n296 B.n295 163.367
R401 B.n295 B.n90 163.367
R402 B.n291 B.n90 163.367
R403 B.n291 B.n290 163.367
R404 B.n290 B.n289 163.367
R405 B.n289 B.n92 163.367
R406 B.n285 B.n92 163.367
R407 B.n285 B.n284 163.367
R408 B.n284 B.n283 163.367
R409 B.n483 B.n482 163.367
R410 B.n482 B.n23 163.367
R411 B.n478 B.n23 163.367
R412 B.n478 B.n477 163.367
R413 B.n477 B.n476 163.367
R414 B.n476 B.n25 163.367
R415 B.n472 B.n25 163.367
R416 B.n472 B.n471 163.367
R417 B.n471 B.n470 163.367
R418 B.n470 B.n27 163.367
R419 B.n466 B.n27 163.367
R420 B.n466 B.n465 163.367
R421 B.n465 B.n464 163.367
R422 B.n464 B.n29 163.367
R423 B.n460 B.n29 163.367
R424 B.n460 B.n459 163.367
R425 B.n459 B.n458 163.367
R426 B.n458 B.n31 163.367
R427 B.n454 B.n31 163.367
R428 B.n454 B.n453 163.367
R429 B.n453 B.n452 163.367
R430 B.n452 B.n33 163.367
R431 B.n448 B.n33 163.367
R432 B.n448 B.n447 163.367
R433 B.n447 B.n446 163.367
R434 B.n446 B.n38 163.367
R435 B.n442 B.n38 163.367
R436 B.n442 B.n441 163.367
R437 B.n441 B.n440 163.367
R438 B.n440 B.n40 163.367
R439 B.n435 B.n40 163.367
R440 B.n435 B.n434 163.367
R441 B.n434 B.n433 163.367
R442 B.n433 B.n44 163.367
R443 B.n429 B.n44 163.367
R444 B.n429 B.n428 163.367
R445 B.n428 B.n427 163.367
R446 B.n427 B.n46 163.367
R447 B.n423 B.n46 163.367
R448 B.n423 B.n422 163.367
R449 B.n422 B.n421 163.367
R450 B.n421 B.n48 163.367
R451 B.n417 B.n48 163.367
R452 B.n417 B.n416 163.367
R453 B.n416 B.n415 163.367
R454 B.n415 B.n50 163.367
R455 B.n411 B.n50 163.367
R456 B.n411 B.n410 163.367
R457 B.n410 B.n409 163.367
R458 B.n409 B.n52 163.367
R459 B.n405 B.n52 163.367
R460 B.n484 B.n21 163.367
R461 B.n488 B.n21 163.367
R462 B.n489 B.n488 163.367
R463 B.n490 B.n489 163.367
R464 B.n490 B.n19 163.367
R465 B.n494 B.n19 163.367
R466 B.n495 B.n494 163.367
R467 B.n496 B.n495 163.367
R468 B.n496 B.n17 163.367
R469 B.n500 B.n17 163.367
R470 B.n501 B.n500 163.367
R471 B.n502 B.n501 163.367
R472 B.n502 B.n15 163.367
R473 B.n506 B.n15 163.367
R474 B.n507 B.n506 163.367
R475 B.n508 B.n507 163.367
R476 B.n508 B.n13 163.367
R477 B.n512 B.n13 163.367
R478 B.n513 B.n512 163.367
R479 B.n514 B.n513 163.367
R480 B.n514 B.n11 163.367
R481 B.n518 B.n11 163.367
R482 B.n519 B.n518 163.367
R483 B.n520 B.n519 163.367
R484 B.n520 B.n9 163.367
R485 B.n524 B.n9 163.367
R486 B.n525 B.n524 163.367
R487 B.n526 B.n525 163.367
R488 B.n526 B.n7 163.367
R489 B.n530 B.n7 163.367
R490 B.n531 B.n530 163.367
R491 B.n532 B.n531 163.367
R492 B.n532 B.n5 163.367
R493 B.n536 B.n5 163.367
R494 B.n537 B.n536 163.367
R495 B.n538 B.n537 163.367
R496 B.n538 B.n3 163.367
R497 B.n542 B.n3 163.367
R498 B.n543 B.n542 163.367
R499 B.n142 B.n2 163.367
R500 B.n143 B.n142 163.367
R501 B.n143 B.n140 163.367
R502 B.n147 B.n140 163.367
R503 B.n148 B.n147 163.367
R504 B.n149 B.n148 163.367
R505 B.n149 B.n138 163.367
R506 B.n153 B.n138 163.367
R507 B.n154 B.n153 163.367
R508 B.n155 B.n154 163.367
R509 B.n155 B.n136 163.367
R510 B.n159 B.n136 163.367
R511 B.n160 B.n159 163.367
R512 B.n161 B.n160 163.367
R513 B.n161 B.n134 163.367
R514 B.n165 B.n134 163.367
R515 B.n166 B.n165 163.367
R516 B.n167 B.n166 163.367
R517 B.n167 B.n132 163.367
R518 B.n171 B.n132 163.367
R519 B.n172 B.n171 163.367
R520 B.n173 B.n172 163.367
R521 B.n173 B.n130 163.367
R522 B.n177 B.n130 163.367
R523 B.n178 B.n177 163.367
R524 B.n179 B.n178 163.367
R525 B.n179 B.n128 163.367
R526 B.n183 B.n128 163.367
R527 B.n184 B.n183 163.367
R528 B.n185 B.n184 163.367
R529 B.n185 B.n126 163.367
R530 B.n189 B.n126 163.367
R531 B.n190 B.n189 163.367
R532 B.n191 B.n190 163.367
R533 B.n191 B.n124 163.367
R534 B.n195 B.n124 163.367
R535 B.n196 B.n195 163.367
R536 B.n197 B.n196 163.367
R537 B.n197 B.n122 163.367
R538 B.n105 B.t4 162.383
R539 B.n41 B.t11 162.383
R540 B.n230 B.t7 162.38
R541 B.n34 B.t2 162.38
R542 B.n106 B.t5 119.718
R543 B.n42 B.t10 119.718
R544 B.n231 B.t8 119.713
R545 B.n35 B.t1 119.713
R546 B.n232 B.n231 59.5399
R547 B.n250 B.n106 59.5399
R548 B.n437 B.n42 59.5399
R549 B.n36 B.n35 59.5399
R550 B.n231 B.n230 42.6672
R551 B.n106 B.n105 42.6672
R552 B.n42 B.n41 42.6672
R553 B.n35 B.n34 42.6672
R554 B.n485 B.n22 31.0639
R555 B.n406 B.n53 31.0639
R556 B.n282 B.n281 31.0639
R557 B.n200 B.n199 31.0639
R558 B B.n545 18.0485
R559 B.n486 B.n485 10.6151
R560 B.n487 B.n486 10.6151
R561 B.n487 B.n20 10.6151
R562 B.n491 B.n20 10.6151
R563 B.n492 B.n491 10.6151
R564 B.n493 B.n492 10.6151
R565 B.n493 B.n18 10.6151
R566 B.n497 B.n18 10.6151
R567 B.n498 B.n497 10.6151
R568 B.n499 B.n498 10.6151
R569 B.n499 B.n16 10.6151
R570 B.n503 B.n16 10.6151
R571 B.n504 B.n503 10.6151
R572 B.n505 B.n504 10.6151
R573 B.n505 B.n14 10.6151
R574 B.n509 B.n14 10.6151
R575 B.n510 B.n509 10.6151
R576 B.n511 B.n510 10.6151
R577 B.n511 B.n12 10.6151
R578 B.n515 B.n12 10.6151
R579 B.n516 B.n515 10.6151
R580 B.n517 B.n516 10.6151
R581 B.n517 B.n10 10.6151
R582 B.n521 B.n10 10.6151
R583 B.n522 B.n521 10.6151
R584 B.n523 B.n522 10.6151
R585 B.n523 B.n8 10.6151
R586 B.n527 B.n8 10.6151
R587 B.n528 B.n527 10.6151
R588 B.n529 B.n528 10.6151
R589 B.n529 B.n6 10.6151
R590 B.n533 B.n6 10.6151
R591 B.n534 B.n533 10.6151
R592 B.n535 B.n534 10.6151
R593 B.n535 B.n4 10.6151
R594 B.n539 B.n4 10.6151
R595 B.n540 B.n539 10.6151
R596 B.n541 B.n540 10.6151
R597 B.n541 B.n0 10.6151
R598 B.n481 B.n22 10.6151
R599 B.n481 B.n480 10.6151
R600 B.n480 B.n479 10.6151
R601 B.n479 B.n24 10.6151
R602 B.n475 B.n24 10.6151
R603 B.n475 B.n474 10.6151
R604 B.n474 B.n473 10.6151
R605 B.n473 B.n26 10.6151
R606 B.n469 B.n26 10.6151
R607 B.n469 B.n468 10.6151
R608 B.n468 B.n467 10.6151
R609 B.n467 B.n28 10.6151
R610 B.n463 B.n28 10.6151
R611 B.n463 B.n462 10.6151
R612 B.n462 B.n461 10.6151
R613 B.n461 B.n30 10.6151
R614 B.n457 B.n30 10.6151
R615 B.n457 B.n456 10.6151
R616 B.n456 B.n455 10.6151
R617 B.n455 B.n32 10.6151
R618 B.n451 B.n450 10.6151
R619 B.n450 B.n449 10.6151
R620 B.n449 B.n37 10.6151
R621 B.n445 B.n37 10.6151
R622 B.n445 B.n444 10.6151
R623 B.n444 B.n443 10.6151
R624 B.n443 B.n39 10.6151
R625 B.n439 B.n39 10.6151
R626 B.n439 B.n438 10.6151
R627 B.n436 B.n43 10.6151
R628 B.n432 B.n43 10.6151
R629 B.n432 B.n431 10.6151
R630 B.n431 B.n430 10.6151
R631 B.n430 B.n45 10.6151
R632 B.n426 B.n45 10.6151
R633 B.n426 B.n425 10.6151
R634 B.n425 B.n424 10.6151
R635 B.n424 B.n47 10.6151
R636 B.n420 B.n47 10.6151
R637 B.n420 B.n419 10.6151
R638 B.n419 B.n418 10.6151
R639 B.n418 B.n49 10.6151
R640 B.n414 B.n49 10.6151
R641 B.n414 B.n413 10.6151
R642 B.n413 B.n412 10.6151
R643 B.n412 B.n51 10.6151
R644 B.n408 B.n51 10.6151
R645 B.n408 B.n407 10.6151
R646 B.n407 B.n406 10.6151
R647 B.n402 B.n53 10.6151
R648 B.n402 B.n401 10.6151
R649 B.n401 B.n400 10.6151
R650 B.n400 B.n55 10.6151
R651 B.n396 B.n55 10.6151
R652 B.n396 B.n395 10.6151
R653 B.n395 B.n394 10.6151
R654 B.n394 B.n57 10.6151
R655 B.n390 B.n57 10.6151
R656 B.n390 B.n389 10.6151
R657 B.n389 B.n388 10.6151
R658 B.n388 B.n59 10.6151
R659 B.n384 B.n59 10.6151
R660 B.n384 B.n383 10.6151
R661 B.n383 B.n382 10.6151
R662 B.n382 B.n61 10.6151
R663 B.n378 B.n61 10.6151
R664 B.n378 B.n377 10.6151
R665 B.n377 B.n376 10.6151
R666 B.n376 B.n63 10.6151
R667 B.n372 B.n63 10.6151
R668 B.n372 B.n371 10.6151
R669 B.n371 B.n370 10.6151
R670 B.n370 B.n65 10.6151
R671 B.n366 B.n65 10.6151
R672 B.n366 B.n365 10.6151
R673 B.n365 B.n364 10.6151
R674 B.n364 B.n67 10.6151
R675 B.n360 B.n67 10.6151
R676 B.n360 B.n359 10.6151
R677 B.n359 B.n358 10.6151
R678 B.n358 B.n69 10.6151
R679 B.n354 B.n69 10.6151
R680 B.n354 B.n353 10.6151
R681 B.n353 B.n352 10.6151
R682 B.n352 B.n71 10.6151
R683 B.n348 B.n71 10.6151
R684 B.n348 B.n347 10.6151
R685 B.n347 B.n346 10.6151
R686 B.n346 B.n73 10.6151
R687 B.n342 B.n73 10.6151
R688 B.n342 B.n341 10.6151
R689 B.n341 B.n340 10.6151
R690 B.n340 B.n75 10.6151
R691 B.n336 B.n75 10.6151
R692 B.n336 B.n335 10.6151
R693 B.n335 B.n334 10.6151
R694 B.n334 B.n77 10.6151
R695 B.n330 B.n77 10.6151
R696 B.n330 B.n329 10.6151
R697 B.n329 B.n328 10.6151
R698 B.n328 B.n79 10.6151
R699 B.n324 B.n79 10.6151
R700 B.n324 B.n323 10.6151
R701 B.n323 B.n322 10.6151
R702 B.n322 B.n81 10.6151
R703 B.n318 B.n81 10.6151
R704 B.n318 B.n317 10.6151
R705 B.n317 B.n316 10.6151
R706 B.n316 B.n83 10.6151
R707 B.n312 B.n83 10.6151
R708 B.n312 B.n311 10.6151
R709 B.n311 B.n310 10.6151
R710 B.n310 B.n85 10.6151
R711 B.n306 B.n85 10.6151
R712 B.n306 B.n305 10.6151
R713 B.n305 B.n304 10.6151
R714 B.n304 B.n87 10.6151
R715 B.n300 B.n87 10.6151
R716 B.n300 B.n299 10.6151
R717 B.n299 B.n298 10.6151
R718 B.n298 B.n89 10.6151
R719 B.n294 B.n89 10.6151
R720 B.n294 B.n293 10.6151
R721 B.n293 B.n292 10.6151
R722 B.n292 B.n91 10.6151
R723 B.n288 B.n91 10.6151
R724 B.n288 B.n287 10.6151
R725 B.n287 B.n286 10.6151
R726 B.n286 B.n93 10.6151
R727 B.n282 B.n93 10.6151
R728 B.n141 B.n1 10.6151
R729 B.n144 B.n141 10.6151
R730 B.n145 B.n144 10.6151
R731 B.n146 B.n145 10.6151
R732 B.n146 B.n139 10.6151
R733 B.n150 B.n139 10.6151
R734 B.n151 B.n150 10.6151
R735 B.n152 B.n151 10.6151
R736 B.n152 B.n137 10.6151
R737 B.n156 B.n137 10.6151
R738 B.n157 B.n156 10.6151
R739 B.n158 B.n157 10.6151
R740 B.n158 B.n135 10.6151
R741 B.n162 B.n135 10.6151
R742 B.n163 B.n162 10.6151
R743 B.n164 B.n163 10.6151
R744 B.n164 B.n133 10.6151
R745 B.n168 B.n133 10.6151
R746 B.n169 B.n168 10.6151
R747 B.n170 B.n169 10.6151
R748 B.n170 B.n131 10.6151
R749 B.n174 B.n131 10.6151
R750 B.n175 B.n174 10.6151
R751 B.n176 B.n175 10.6151
R752 B.n176 B.n129 10.6151
R753 B.n180 B.n129 10.6151
R754 B.n181 B.n180 10.6151
R755 B.n182 B.n181 10.6151
R756 B.n182 B.n127 10.6151
R757 B.n186 B.n127 10.6151
R758 B.n187 B.n186 10.6151
R759 B.n188 B.n187 10.6151
R760 B.n188 B.n125 10.6151
R761 B.n192 B.n125 10.6151
R762 B.n193 B.n192 10.6151
R763 B.n194 B.n193 10.6151
R764 B.n194 B.n123 10.6151
R765 B.n198 B.n123 10.6151
R766 B.n199 B.n198 10.6151
R767 B.n200 B.n121 10.6151
R768 B.n204 B.n121 10.6151
R769 B.n205 B.n204 10.6151
R770 B.n206 B.n205 10.6151
R771 B.n206 B.n119 10.6151
R772 B.n210 B.n119 10.6151
R773 B.n211 B.n210 10.6151
R774 B.n212 B.n211 10.6151
R775 B.n212 B.n117 10.6151
R776 B.n216 B.n117 10.6151
R777 B.n217 B.n216 10.6151
R778 B.n218 B.n217 10.6151
R779 B.n218 B.n115 10.6151
R780 B.n222 B.n115 10.6151
R781 B.n223 B.n222 10.6151
R782 B.n224 B.n223 10.6151
R783 B.n224 B.n113 10.6151
R784 B.n228 B.n113 10.6151
R785 B.n229 B.n228 10.6151
R786 B.n233 B.n229 10.6151
R787 B.n237 B.n111 10.6151
R788 B.n238 B.n237 10.6151
R789 B.n239 B.n238 10.6151
R790 B.n239 B.n109 10.6151
R791 B.n243 B.n109 10.6151
R792 B.n244 B.n243 10.6151
R793 B.n245 B.n244 10.6151
R794 B.n245 B.n107 10.6151
R795 B.n249 B.n107 10.6151
R796 B.n252 B.n251 10.6151
R797 B.n252 B.n103 10.6151
R798 B.n256 B.n103 10.6151
R799 B.n257 B.n256 10.6151
R800 B.n258 B.n257 10.6151
R801 B.n258 B.n101 10.6151
R802 B.n262 B.n101 10.6151
R803 B.n263 B.n262 10.6151
R804 B.n264 B.n263 10.6151
R805 B.n264 B.n99 10.6151
R806 B.n268 B.n99 10.6151
R807 B.n269 B.n268 10.6151
R808 B.n270 B.n269 10.6151
R809 B.n270 B.n97 10.6151
R810 B.n274 B.n97 10.6151
R811 B.n275 B.n274 10.6151
R812 B.n276 B.n275 10.6151
R813 B.n276 B.n95 10.6151
R814 B.n280 B.n95 10.6151
R815 B.n281 B.n280 10.6151
R816 B.n36 B.n32 9.36635
R817 B.n437 B.n436 9.36635
R818 B.n233 B.n232 9.36635
R819 B.n251 B.n250 9.36635
R820 B.n545 B.n0 8.11757
R821 B.n545 B.n1 8.11757
R822 B.n451 B.n36 1.24928
R823 B.n438 B.n437 1.24928
R824 B.n232 B.n111 1.24928
R825 B.n250 B.n249 1.24928
R826 VP.n31 VP.n7 183.321
R827 VP.n56 VP.n55 183.321
R828 VP.n30 VP.n29 183.321
R829 VP.n15 VP.n12 161.3
R830 VP.n17 VP.n16 161.3
R831 VP.n18 VP.n11 161.3
R832 VP.n20 VP.n19 161.3
R833 VP.n22 VP.n10 161.3
R834 VP.n24 VP.n23 161.3
R835 VP.n25 VP.n9 161.3
R836 VP.n27 VP.n26 161.3
R837 VP.n28 VP.n8 161.3
R838 VP.n54 VP.n0 161.3
R839 VP.n53 VP.n52 161.3
R840 VP.n51 VP.n1 161.3
R841 VP.n50 VP.n49 161.3
R842 VP.n48 VP.n2 161.3
R843 VP.n46 VP.n45 161.3
R844 VP.n44 VP.n3 161.3
R845 VP.n43 VP.n42 161.3
R846 VP.n41 VP.n4 161.3
R847 VP.n39 VP.n38 161.3
R848 VP.n37 VP.n5 161.3
R849 VP.n36 VP.n35 161.3
R850 VP.n34 VP.n6 161.3
R851 VP.n33 VP.n32 161.3
R852 VP.n13 VP.t6 98.2057
R853 VP.n7 VP.t3 64.8256
R854 VP.n40 VP.t5 64.8256
R855 VP.n47 VP.t7 64.8256
R856 VP.n55 VP.t0 64.8256
R857 VP.n29 VP.t2 64.8256
R858 VP.n21 VP.t1 64.8256
R859 VP.n14 VP.t4 64.8256
R860 VP.n42 VP.n3 56.5193
R861 VP.n16 VP.n11 56.5193
R862 VP.n14 VP.n13 52.6042
R863 VP.n35 VP.n5 45.3497
R864 VP.n49 VP.n1 45.3497
R865 VP.n23 VP.n9 45.3497
R866 VP.n31 VP.n30 42.099
R867 VP.n35 VP.n34 35.6371
R868 VP.n53 VP.n1 35.6371
R869 VP.n27 VP.n9 35.6371
R870 VP.n34 VP.n33 24.4675
R871 VP.n39 VP.n5 24.4675
R872 VP.n42 VP.n41 24.4675
R873 VP.n46 VP.n3 24.4675
R874 VP.n49 VP.n48 24.4675
R875 VP.n54 VP.n53 24.4675
R876 VP.n28 VP.n27 24.4675
R877 VP.n20 VP.n11 24.4675
R878 VP.n23 VP.n22 24.4675
R879 VP.n16 VP.n15 24.4675
R880 VP.n41 VP.n40 17.1274
R881 VP.n47 VP.n46 17.1274
R882 VP.n21 VP.n20 17.1274
R883 VP.n15 VP.n14 17.1274
R884 VP.n13 VP.n12 12.4054
R885 VP.n40 VP.n39 7.3406
R886 VP.n48 VP.n47 7.3406
R887 VP.n22 VP.n21 7.3406
R888 VP.n33 VP.n7 2.4472
R889 VP.n55 VP.n54 2.4472
R890 VP.n29 VP.n28 2.4472
R891 VP.n17 VP.n12 0.189894
R892 VP.n18 VP.n17 0.189894
R893 VP.n19 VP.n18 0.189894
R894 VP.n19 VP.n10 0.189894
R895 VP.n24 VP.n10 0.189894
R896 VP.n25 VP.n24 0.189894
R897 VP.n26 VP.n25 0.189894
R898 VP.n26 VP.n8 0.189894
R899 VP.n30 VP.n8 0.189894
R900 VP.n32 VP.n31 0.189894
R901 VP.n32 VP.n6 0.189894
R902 VP.n36 VP.n6 0.189894
R903 VP.n37 VP.n36 0.189894
R904 VP.n38 VP.n37 0.189894
R905 VP.n38 VP.n4 0.189894
R906 VP.n43 VP.n4 0.189894
R907 VP.n44 VP.n43 0.189894
R908 VP.n45 VP.n44 0.189894
R909 VP.n45 VP.n2 0.189894
R910 VP.n50 VP.n2 0.189894
R911 VP.n51 VP.n50 0.189894
R912 VP.n52 VP.n51 0.189894
R913 VP.n52 VP.n0 0.189894
R914 VP.n56 VP.n0 0.189894
R915 VP VP.n56 0.0516364
R916 VTAIL.n11 VTAIL.t9 92.3575
R917 VTAIL.n10 VTAIL.t11 92.3575
R918 VTAIL.n7 VTAIL.t12 92.3575
R919 VTAIL.n15 VTAIL.t0 92.3574
R920 VTAIL.n2 VTAIL.t1 92.3574
R921 VTAIL.n3 VTAIL.t10 92.3574
R922 VTAIL.n6 VTAIL.t6 92.3574
R923 VTAIL.n14 VTAIL.t5 92.3574
R924 VTAIL.n13 VTAIL.n12 85.8953
R925 VTAIL.n9 VTAIL.n8 85.8953
R926 VTAIL.n1 VTAIL.n0 85.8951
R927 VTAIL.n5 VTAIL.n4 85.8951
R928 VTAIL.n15 VTAIL.n14 18.5996
R929 VTAIL.n7 VTAIL.n6 18.5996
R930 VTAIL.n0 VTAIL.t13 6.46273
R931 VTAIL.n0 VTAIL.t2 6.46273
R932 VTAIL.n4 VTAIL.t3 6.46273
R933 VTAIL.n4 VTAIL.t7 6.46273
R934 VTAIL.n12 VTAIL.t8 6.46273
R935 VTAIL.n12 VTAIL.t4 6.46273
R936 VTAIL.n8 VTAIL.t14 6.46273
R937 VTAIL.n8 VTAIL.t15 6.46273
R938 VTAIL.n9 VTAIL.n7 1.89705
R939 VTAIL.n10 VTAIL.n9 1.89705
R940 VTAIL.n13 VTAIL.n11 1.89705
R941 VTAIL.n14 VTAIL.n13 1.89705
R942 VTAIL.n6 VTAIL.n5 1.89705
R943 VTAIL.n5 VTAIL.n3 1.89705
R944 VTAIL.n2 VTAIL.n1 1.89705
R945 VTAIL VTAIL.n15 1.83886
R946 VTAIL.n11 VTAIL.n10 0.470328
R947 VTAIL.n3 VTAIL.n2 0.470328
R948 VTAIL VTAIL.n1 0.0586897
R949 VDD1 VDD1.n0 103.581
R950 VDD1.n3 VDD1.n2 103.466
R951 VDD1.n3 VDD1.n1 103.466
R952 VDD1.n5 VDD1.n4 102.573
R953 VDD1.n5 VDD1.n3 37.169
R954 VDD1.n4 VDD1.t6 6.46273
R955 VDD1.n4 VDD1.t5 6.46273
R956 VDD1.n0 VDD1.t1 6.46273
R957 VDD1.n0 VDD1.t3 6.46273
R958 VDD1.n2 VDD1.t0 6.46273
R959 VDD1.n2 VDD1.t7 6.46273
R960 VDD1.n1 VDD1.t4 6.46273
R961 VDD1.n1 VDD1.t2 6.46273
R962 VDD1 VDD1.n5 0.890586
R963 VN.n22 VN.n21 183.321
R964 VN.n45 VN.n44 183.321
R965 VN.n43 VN.n23 161.3
R966 VN.n42 VN.n41 161.3
R967 VN.n40 VN.n24 161.3
R968 VN.n39 VN.n38 161.3
R969 VN.n37 VN.n25 161.3
R970 VN.n35 VN.n34 161.3
R971 VN.n33 VN.n26 161.3
R972 VN.n32 VN.n31 161.3
R973 VN.n30 VN.n27 161.3
R974 VN.n20 VN.n0 161.3
R975 VN.n19 VN.n18 161.3
R976 VN.n17 VN.n1 161.3
R977 VN.n16 VN.n15 161.3
R978 VN.n14 VN.n2 161.3
R979 VN.n12 VN.n11 161.3
R980 VN.n10 VN.n3 161.3
R981 VN.n9 VN.n8 161.3
R982 VN.n7 VN.n4 161.3
R983 VN.n5 VN.t5 98.2057
R984 VN.n28 VN.t4 98.2057
R985 VN.n6 VN.t1 64.8256
R986 VN.n13 VN.t7 64.8256
R987 VN.n21 VN.t6 64.8256
R988 VN.n29 VN.t2 64.8256
R989 VN.n36 VN.t3 64.8256
R990 VN.n44 VN.t0 64.8256
R991 VN.n8 VN.n3 56.5193
R992 VN.n31 VN.n26 56.5193
R993 VN.n6 VN.n5 52.6042
R994 VN.n29 VN.n28 52.6042
R995 VN.n15 VN.n1 45.3497
R996 VN.n38 VN.n24 45.3497
R997 VN VN.n45 42.4797
R998 VN.n19 VN.n1 35.6371
R999 VN.n42 VN.n24 35.6371
R1000 VN.n8 VN.n7 24.4675
R1001 VN.n12 VN.n3 24.4675
R1002 VN.n15 VN.n14 24.4675
R1003 VN.n20 VN.n19 24.4675
R1004 VN.n31 VN.n30 24.4675
R1005 VN.n38 VN.n37 24.4675
R1006 VN.n35 VN.n26 24.4675
R1007 VN.n43 VN.n42 24.4675
R1008 VN.n7 VN.n6 17.1274
R1009 VN.n13 VN.n12 17.1274
R1010 VN.n30 VN.n29 17.1274
R1011 VN.n36 VN.n35 17.1274
R1012 VN.n28 VN.n27 12.4054
R1013 VN.n5 VN.n4 12.4054
R1014 VN.n14 VN.n13 7.3406
R1015 VN.n37 VN.n36 7.3406
R1016 VN.n21 VN.n20 2.4472
R1017 VN.n44 VN.n43 2.4472
R1018 VN.n45 VN.n23 0.189894
R1019 VN.n41 VN.n23 0.189894
R1020 VN.n41 VN.n40 0.189894
R1021 VN.n40 VN.n39 0.189894
R1022 VN.n39 VN.n25 0.189894
R1023 VN.n34 VN.n25 0.189894
R1024 VN.n34 VN.n33 0.189894
R1025 VN.n33 VN.n32 0.189894
R1026 VN.n32 VN.n27 0.189894
R1027 VN.n9 VN.n4 0.189894
R1028 VN.n10 VN.n9 0.189894
R1029 VN.n11 VN.n10 0.189894
R1030 VN.n11 VN.n2 0.189894
R1031 VN.n16 VN.n2 0.189894
R1032 VN.n17 VN.n16 0.189894
R1033 VN.n18 VN.n17 0.189894
R1034 VN.n18 VN.n0 0.189894
R1035 VN.n22 VN.n0 0.189894
R1036 VN VN.n22 0.0516364
R1037 VDD2.n2 VDD2.n1 103.466
R1038 VDD2.n2 VDD2.n0 103.466
R1039 VDD2 VDD2.n5 103.465
R1040 VDD2.n4 VDD2.n3 102.575
R1041 VDD2.n4 VDD2.n2 36.586
R1042 VDD2.n5 VDD2.t5 6.46273
R1043 VDD2.n5 VDD2.t3 6.46273
R1044 VDD2.n3 VDD2.t7 6.46273
R1045 VDD2.n3 VDD2.t4 6.46273
R1046 VDD2.n1 VDD2.t0 6.46273
R1047 VDD2.n1 VDD2.t1 6.46273
R1048 VDD2.n0 VDD2.t2 6.46273
R1049 VDD2.n0 VDD2.t6 6.46273
R1050 VDD2 VDD2.n4 1.00697
C0 VP VDD1 3.92798f
C1 VN VTAIL 4.221839f
C2 w_n3170_n1974# VP 6.53044f
C3 VP B 1.67776f
C4 VDD2 VTAIL 5.38214f
C5 VDD2 VN 3.63752f
C6 VTAIL VDD1 5.33262f
C7 w_n3170_n1974# VTAIL 2.54811f
C8 VTAIL B 2.43003f
C9 VN VDD1 0.150065f
C10 VN w_n3170_n1974# 6.12114f
C11 VN B 0.995451f
C12 VDD2 VDD1 1.39516f
C13 VDD2 w_n3170_n1974# 1.60724f
C14 VDD2 B 1.31296f
C15 VP VTAIL 4.23595f
C16 w_n3170_n1974# VDD1 1.52342f
C17 VDD1 B 1.23982f
C18 VN VP 5.47801f
C19 w_n3170_n1974# B 7.05147f
C20 VDD2 VP 0.445826f
C21 VDD2 VSUBS 1.345845f
C22 VDD1 VSUBS 1.869803f
C23 VTAIL VSUBS 0.609278f
C24 VN VSUBS 5.45993f
C25 VP VSUBS 2.3749f
C26 B VSUBS 3.407136f
C27 w_n3170_n1974# VSUBS 78.4004f
C28 VDD2.t2 VSUBS 0.097247f
C29 VDD2.t6 VSUBS 0.097247f
C30 VDD2.n0 VSUBS 0.618546f
C31 VDD2.t0 VSUBS 0.097247f
C32 VDD2.t1 VSUBS 0.097247f
C33 VDD2.n1 VSUBS 0.618546f
C34 VDD2.n2 VSUBS 2.72555f
C35 VDD2.t7 VSUBS 0.097247f
C36 VDD2.t4 VSUBS 0.097247f
C37 VDD2.n3 VSUBS 0.613331f
C38 VDD2.n4 VSUBS 2.27943f
C39 VDD2.t5 VSUBS 0.097247f
C40 VDD2.t3 VSUBS 0.097247f
C41 VDD2.n5 VSUBS 0.618522f
C42 VN.n0 VSUBS 0.043974f
C43 VN.t6 VSUBS 1.08235f
C44 VN.n1 VSUBS 0.036981f
C45 VN.n2 VSUBS 0.043974f
C46 VN.t7 VSUBS 1.08235f
C47 VN.n3 VSUBS 0.064194f
C48 VN.n4 VSUBS 0.325547f
C49 VN.t1 VSUBS 1.08235f
C50 VN.t5 VSUBS 1.30009f
C51 VN.n5 VSUBS 0.521337f
C52 VN.n6 VSUBS 0.535094f
C53 VN.n7 VSUBS 0.069817f
C54 VN.n8 VSUBS 0.064194f
C55 VN.n9 VSUBS 0.043974f
C56 VN.n10 VSUBS 0.043974f
C57 VN.n11 VSUBS 0.043974f
C58 VN.n12 VSUBS 0.069817f
C59 VN.n13 VSUBS 0.42685f
C60 VN.n14 VSUBS 0.053633f
C61 VN.n15 VSUBS 0.084561f
C62 VN.n16 VSUBS 0.043974f
C63 VN.n17 VSUBS 0.043974f
C64 VN.n18 VSUBS 0.043974f
C65 VN.n19 VSUBS 0.088801f
C66 VN.n20 VSUBS 0.04554f
C67 VN.n21 VSUBS 0.528868f
C68 VN.n22 VSUBS 0.048005f
C69 VN.n23 VSUBS 0.043974f
C70 VN.t0 VSUBS 1.08235f
C71 VN.n24 VSUBS 0.036981f
C72 VN.n25 VSUBS 0.043974f
C73 VN.t3 VSUBS 1.08235f
C74 VN.n26 VSUBS 0.064194f
C75 VN.n27 VSUBS 0.325547f
C76 VN.t2 VSUBS 1.08235f
C77 VN.t4 VSUBS 1.30009f
C78 VN.n28 VSUBS 0.521337f
C79 VN.n29 VSUBS 0.535094f
C80 VN.n30 VSUBS 0.069817f
C81 VN.n31 VSUBS 0.064194f
C82 VN.n32 VSUBS 0.043974f
C83 VN.n33 VSUBS 0.043974f
C84 VN.n34 VSUBS 0.043974f
C85 VN.n35 VSUBS 0.069817f
C86 VN.n36 VSUBS 0.42685f
C87 VN.n37 VSUBS 0.053633f
C88 VN.n38 VSUBS 0.084561f
C89 VN.n39 VSUBS 0.043974f
C90 VN.n40 VSUBS 0.043974f
C91 VN.n41 VSUBS 0.043974f
C92 VN.n42 VSUBS 0.088801f
C93 VN.n43 VSUBS 0.04554f
C94 VN.n44 VSUBS 0.528868f
C95 VN.n45 VSUBS 1.86502f
C96 VDD1.t1 VSUBS 0.09842f
C97 VDD1.t3 VSUBS 0.09842f
C98 VDD1.n0 VSUBS 0.626756f
C99 VDD1.t4 VSUBS 0.09842f
C100 VDD1.t2 VSUBS 0.09842f
C101 VDD1.n1 VSUBS 0.626007f
C102 VDD1.t0 VSUBS 0.09842f
C103 VDD1.t7 VSUBS 0.09842f
C104 VDD1.n2 VSUBS 0.626007f
C105 VDD1.n3 VSUBS 2.81064f
C106 VDD1.t6 VSUBS 0.09842f
C107 VDD1.t5 VSUBS 0.09842f
C108 VDD1.n4 VSUBS 0.620725f
C109 VDD1.n5 VSUBS 2.33687f
C110 VTAIL.t13 VSUBS 0.115617f
C111 VTAIL.t2 VSUBS 0.115617f
C112 VTAIL.n0 VSUBS 0.643866f
C113 VTAIL.n1 VSUBS 0.673939f
C114 VTAIL.t1 VSUBS 0.900161f
C115 VTAIL.n2 VSUBS 0.771545f
C116 VTAIL.t10 VSUBS 0.900161f
C117 VTAIL.n3 VSUBS 0.771545f
C118 VTAIL.t3 VSUBS 0.115617f
C119 VTAIL.t7 VSUBS 0.115617f
C120 VTAIL.n4 VSUBS 0.643866f
C121 VTAIL.n5 VSUBS 0.84624f
C122 VTAIL.t6 VSUBS 0.900161f
C123 VTAIL.n6 VSUBS 1.70679f
C124 VTAIL.t12 VSUBS 0.900166f
C125 VTAIL.n7 VSUBS 1.70679f
C126 VTAIL.t14 VSUBS 0.115617f
C127 VTAIL.t15 VSUBS 0.115617f
C128 VTAIL.n8 VSUBS 0.643869f
C129 VTAIL.n9 VSUBS 0.846236f
C130 VTAIL.t11 VSUBS 0.900166f
C131 VTAIL.n10 VSUBS 0.77154f
C132 VTAIL.t9 VSUBS 0.900166f
C133 VTAIL.n11 VSUBS 0.77154f
C134 VTAIL.t8 VSUBS 0.115617f
C135 VTAIL.t4 VSUBS 0.115617f
C136 VTAIL.n12 VSUBS 0.643869f
C137 VTAIL.n13 VSUBS 0.846236f
C138 VTAIL.t5 VSUBS 0.900161f
C139 VTAIL.n14 VSUBS 1.70679f
C140 VTAIL.t0 VSUBS 0.900161f
C141 VTAIL.n15 VSUBS 1.70134f
C142 VP.n0 VSUBS 0.045706f
C143 VP.t0 VSUBS 1.12499f
C144 VP.n1 VSUBS 0.038438f
C145 VP.n2 VSUBS 0.045706f
C146 VP.t7 VSUBS 1.12499f
C147 VP.n3 VSUBS 0.066723f
C148 VP.n4 VSUBS 0.045706f
C149 VP.t5 VSUBS 1.12499f
C150 VP.n5 VSUBS 0.087892f
C151 VP.n6 VSUBS 0.045706f
C152 VP.t3 VSUBS 1.12499f
C153 VP.n7 VSUBS 0.549702f
C154 VP.n8 VSUBS 0.045706f
C155 VP.t2 VSUBS 1.12499f
C156 VP.n9 VSUBS 0.038438f
C157 VP.n10 VSUBS 0.045706f
C158 VP.t1 VSUBS 1.12499f
C159 VP.n11 VSUBS 0.066723f
C160 VP.n12 VSUBS 0.338371f
C161 VP.t4 VSUBS 1.12499f
C162 VP.t6 VSUBS 1.35131f
C163 VP.n13 VSUBS 0.541874f
C164 VP.n14 VSUBS 0.556174f
C165 VP.n15 VSUBS 0.072568f
C166 VP.n16 VSUBS 0.066723f
C167 VP.n17 VSUBS 0.045706f
C168 VP.n18 VSUBS 0.045706f
C169 VP.n19 VSUBS 0.045706f
C170 VP.n20 VSUBS 0.072568f
C171 VP.n21 VSUBS 0.443666f
C172 VP.n22 VSUBS 0.055746f
C173 VP.n23 VSUBS 0.087892f
C174 VP.n24 VSUBS 0.045706f
C175 VP.n25 VSUBS 0.045706f
C176 VP.n26 VSUBS 0.045706f
C177 VP.n27 VSUBS 0.0923f
C178 VP.n28 VSUBS 0.047334f
C179 VP.n29 VSUBS 0.549702f
C180 VP.n30 VSUBS 1.9085f
C181 VP.n31 VSUBS 1.94752f
C182 VP.n32 VSUBS 0.045706f
C183 VP.n33 VSUBS 0.047334f
C184 VP.n34 VSUBS 0.0923f
C185 VP.n35 VSUBS 0.038438f
C186 VP.n36 VSUBS 0.045706f
C187 VP.n37 VSUBS 0.045706f
C188 VP.n38 VSUBS 0.045706f
C189 VP.n39 VSUBS 0.055746f
C190 VP.n40 VSUBS 0.443666f
C191 VP.n41 VSUBS 0.072568f
C192 VP.n42 VSUBS 0.066723f
C193 VP.n43 VSUBS 0.045706f
C194 VP.n44 VSUBS 0.045706f
C195 VP.n45 VSUBS 0.045706f
C196 VP.n46 VSUBS 0.072568f
C197 VP.n47 VSUBS 0.443666f
C198 VP.n48 VSUBS 0.055746f
C199 VP.n49 VSUBS 0.087892f
C200 VP.n50 VSUBS 0.045706f
C201 VP.n51 VSUBS 0.045706f
C202 VP.n52 VSUBS 0.045706f
C203 VP.n53 VSUBS 0.0923f
C204 VP.n54 VSUBS 0.047334f
C205 VP.n55 VSUBS 0.549702f
C206 VP.n56 VSUBS 0.049896f
C207 B.n0 VSUBS 0.007757f
C208 B.n1 VSUBS 0.007757f
C209 B.n2 VSUBS 0.011473f
C210 B.n3 VSUBS 0.008792f
C211 B.n4 VSUBS 0.008792f
C212 B.n5 VSUBS 0.008792f
C213 B.n6 VSUBS 0.008792f
C214 B.n7 VSUBS 0.008792f
C215 B.n8 VSUBS 0.008792f
C216 B.n9 VSUBS 0.008792f
C217 B.n10 VSUBS 0.008792f
C218 B.n11 VSUBS 0.008792f
C219 B.n12 VSUBS 0.008792f
C220 B.n13 VSUBS 0.008792f
C221 B.n14 VSUBS 0.008792f
C222 B.n15 VSUBS 0.008792f
C223 B.n16 VSUBS 0.008792f
C224 B.n17 VSUBS 0.008792f
C225 B.n18 VSUBS 0.008792f
C226 B.n19 VSUBS 0.008792f
C227 B.n20 VSUBS 0.008792f
C228 B.n21 VSUBS 0.008792f
C229 B.n22 VSUBS 0.020483f
C230 B.n23 VSUBS 0.008792f
C231 B.n24 VSUBS 0.008792f
C232 B.n25 VSUBS 0.008792f
C233 B.n26 VSUBS 0.008792f
C234 B.n27 VSUBS 0.008792f
C235 B.n28 VSUBS 0.008792f
C236 B.n29 VSUBS 0.008792f
C237 B.n30 VSUBS 0.008792f
C238 B.n31 VSUBS 0.008792f
C239 B.n32 VSUBS 0.008275f
C240 B.n33 VSUBS 0.008792f
C241 B.t1 VSUBS 0.176491f
C242 B.t2 VSUBS 0.19541f
C243 B.t0 VSUBS 0.554227f
C244 B.n34 VSUBS 0.121846f
C245 B.n35 VSUBS 0.084541f
C246 B.n36 VSUBS 0.020369f
C247 B.n37 VSUBS 0.008792f
C248 B.n38 VSUBS 0.008792f
C249 B.n39 VSUBS 0.008792f
C250 B.n40 VSUBS 0.008792f
C251 B.t10 VSUBS 0.176491f
C252 B.t11 VSUBS 0.19541f
C253 B.t9 VSUBS 0.554227f
C254 B.n41 VSUBS 0.121847f
C255 B.n42 VSUBS 0.084541f
C256 B.n43 VSUBS 0.008792f
C257 B.n44 VSUBS 0.008792f
C258 B.n45 VSUBS 0.008792f
C259 B.n46 VSUBS 0.008792f
C260 B.n47 VSUBS 0.008792f
C261 B.n48 VSUBS 0.008792f
C262 B.n49 VSUBS 0.008792f
C263 B.n50 VSUBS 0.008792f
C264 B.n51 VSUBS 0.008792f
C265 B.n52 VSUBS 0.008792f
C266 B.n53 VSUBS 0.019338f
C267 B.n54 VSUBS 0.008792f
C268 B.n55 VSUBS 0.008792f
C269 B.n56 VSUBS 0.008792f
C270 B.n57 VSUBS 0.008792f
C271 B.n58 VSUBS 0.008792f
C272 B.n59 VSUBS 0.008792f
C273 B.n60 VSUBS 0.008792f
C274 B.n61 VSUBS 0.008792f
C275 B.n62 VSUBS 0.008792f
C276 B.n63 VSUBS 0.008792f
C277 B.n64 VSUBS 0.008792f
C278 B.n65 VSUBS 0.008792f
C279 B.n66 VSUBS 0.008792f
C280 B.n67 VSUBS 0.008792f
C281 B.n68 VSUBS 0.008792f
C282 B.n69 VSUBS 0.008792f
C283 B.n70 VSUBS 0.008792f
C284 B.n71 VSUBS 0.008792f
C285 B.n72 VSUBS 0.008792f
C286 B.n73 VSUBS 0.008792f
C287 B.n74 VSUBS 0.008792f
C288 B.n75 VSUBS 0.008792f
C289 B.n76 VSUBS 0.008792f
C290 B.n77 VSUBS 0.008792f
C291 B.n78 VSUBS 0.008792f
C292 B.n79 VSUBS 0.008792f
C293 B.n80 VSUBS 0.008792f
C294 B.n81 VSUBS 0.008792f
C295 B.n82 VSUBS 0.008792f
C296 B.n83 VSUBS 0.008792f
C297 B.n84 VSUBS 0.008792f
C298 B.n85 VSUBS 0.008792f
C299 B.n86 VSUBS 0.008792f
C300 B.n87 VSUBS 0.008792f
C301 B.n88 VSUBS 0.008792f
C302 B.n89 VSUBS 0.008792f
C303 B.n90 VSUBS 0.008792f
C304 B.n91 VSUBS 0.008792f
C305 B.n92 VSUBS 0.008792f
C306 B.n93 VSUBS 0.008792f
C307 B.n94 VSUBS 0.020483f
C308 B.n95 VSUBS 0.008792f
C309 B.n96 VSUBS 0.008792f
C310 B.n97 VSUBS 0.008792f
C311 B.n98 VSUBS 0.008792f
C312 B.n99 VSUBS 0.008792f
C313 B.n100 VSUBS 0.008792f
C314 B.n101 VSUBS 0.008792f
C315 B.n102 VSUBS 0.008792f
C316 B.n103 VSUBS 0.008792f
C317 B.n104 VSUBS 0.008792f
C318 B.t5 VSUBS 0.176491f
C319 B.t4 VSUBS 0.19541f
C320 B.t3 VSUBS 0.554227f
C321 B.n105 VSUBS 0.121847f
C322 B.n106 VSUBS 0.084541f
C323 B.n107 VSUBS 0.008792f
C324 B.n108 VSUBS 0.008792f
C325 B.n109 VSUBS 0.008792f
C326 B.n110 VSUBS 0.008792f
C327 B.n111 VSUBS 0.004913f
C328 B.n112 VSUBS 0.008792f
C329 B.n113 VSUBS 0.008792f
C330 B.n114 VSUBS 0.008792f
C331 B.n115 VSUBS 0.008792f
C332 B.n116 VSUBS 0.008792f
C333 B.n117 VSUBS 0.008792f
C334 B.n118 VSUBS 0.008792f
C335 B.n119 VSUBS 0.008792f
C336 B.n120 VSUBS 0.008792f
C337 B.n121 VSUBS 0.008792f
C338 B.n122 VSUBS 0.019338f
C339 B.n123 VSUBS 0.008792f
C340 B.n124 VSUBS 0.008792f
C341 B.n125 VSUBS 0.008792f
C342 B.n126 VSUBS 0.008792f
C343 B.n127 VSUBS 0.008792f
C344 B.n128 VSUBS 0.008792f
C345 B.n129 VSUBS 0.008792f
C346 B.n130 VSUBS 0.008792f
C347 B.n131 VSUBS 0.008792f
C348 B.n132 VSUBS 0.008792f
C349 B.n133 VSUBS 0.008792f
C350 B.n134 VSUBS 0.008792f
C351 B.n135 VSUBS 0.008792f
C352 B.n136 VSUBS 0.008792f
C353 B.n137 VSUBS 0.008792f
C354 B.n138 VSUBS 0.008792f
C355 B.n139 VSUBS 0.008792f
C356 B.n140 VSUBS 0.008792f
C357 B.n141 VSUBS 0.008792f
C358 B.n142 VSUBS 0.008792f
C359 B.n143 VSUBS 0.008792f
C360 B.n144 VSUBS 0.008792f
C361 B.n145 VSUBS 0.008792f
C362 B.n146 VSUBS 0.008792f
C363 B.n147 VSUBS 0.008792f
C364 B.n148 VSUBS 0.008792f
C365 B.n149 VSUBS 0.008792f
C366 B.n150 VSUBS 0.008792f
C367 B.n151 VSUBS 0.008792f
C368 B.n152 VSUBS 0.008792f
C369 B.n153 VSUBS 0.008792f
C370 B.n154 VSUBS 0.008792f
C371 B.n155 VSUBS 0.008792f
C372 B.n156 VSUBS 0.008792f
C373 B.n157 VSUBS 0.008792f
C374 B.n158 VSUBS 0.008792f
C375 B.n159 VSUBS 0.008792f
C376 B.n160 VSUBS 0.008792f
C377 B.n161 VSUBS 0.008792f
C378 B.n162 VSUBS 0.008792f
C379 B.n163 VSUBS 0.008792f
C380 B.n164 VSUBS 0.008792f
C381 B.n165 VSUBS 0.008792f
C382 B.n166 VSUBS 0.008792f
C383 B.n167 VSUBS 0.008792f
C384 B.n168 VSUBS 0.008792f
C385 B.n169 VSUBS 0.008792f
C386 B.n170 VSUBS 0.008792f
C387 B.n171 VSUBS 0.008792f
C388 B.n172 VSUBS 0.008792f
C389 B.n173 VSUBS 0.008792f
C390 B.n174 VSUBS 0.008792f
C391 B.n175 VSUBS 0.008792f
C392 B.n176 VSUBS 0.008792f
C393 B.n177 VSUBS 0.008792f
C394 B.n178 VSUBS 0.008792f
C395 B.n179 VSUBS 0.008792f
C396 B.n180 VSUBS 0.008792f
C397 B.n181 VSUBS 0.008792f
C398 B.n182 VSUBS 0.008792f
C399 B.n183 VSUBS 0.008792f
C400 B.n184 VSUBS 0.008792f
C401 B.n185 VSUBS 0.008792f
C402 B.n186 VSUBS 0.008792f
C403 B.n187 VSUBS 0.008792f
C404 B.n188 VSUBS 0.008792f
C405 B.n189 VSUBS 0.008792f
C406 B.n190 VSUBS 0.008792f
C407 B.n191 VSUBS 0.008792f
C408 B.n192 VSUBS 0.008792f
C409 B.n193 VSUBS 0.008792f
C410 B.n194 VSUBS 0.008792f
C411 B.n195 VSUBS 0.008792f
C412 B.n196 VSUBS 0.008792f
C413 B.n197 VSUBS 0.008792f
C414 B.n198 VSUBS 0.008792f
C415 B.n199 VSUBS 0.019338f
C416 B.n200 VSUBS 0.020483f
C417 B.n201 VSUBS 0.020483f
C418 B.n202 VSUBS 0.008792f
C419 B.n203 VSUBS 0.008792f
C420 B.n204 VSUBS 0.008792f
C421 B.n205 VSUBS 0.008792f
C422 B.n206 VSUBS 0.008792f
C423 B.n207 VSUBS 0.008792f
C424 B.n208 VSUBS 0.008792f
C425 B.n209 VSUBS 0.008792f
C426 B.n210 VSUBS 0.008792f
C427 B.n211 VSUBS 0.008792f
C428 B.n212 VSUBS 0.008792f
C429 B.n213 VSUBS 0.008792f
C430 B.n214 VSUBS 0.008792f
C431 B.n215 VSUBS 0.008792f
C432 B.n216 VSUBS 0.008792f
C433 B.n217 VSUBS 0.008792f
C434 B.n218 VSUBS 0.008792f
C435 B.n219 VSUBS 0.008792f
C436 B.n220 VSUBS 0.008792f
C437 B.n221 VSUBS 0.008792f
C438 B.n222 VSUBS 0.008792f
C439 B.n223 VSUBS 0.008792f
C440 B.n224 VSUBS 0.008792f
C441 B.n225 VSUBS 0.008792f
C442 B.n226 VSUBS 0.008792f
C443 B.n227 VSUBS 0.008792f
C444 B.n228 VSUBS 0.008792f
C445 B.n229 VSUBS 0.008792f
C446 B.t8 VSUBS 0.176491f
C447 B.t7 VSUBS 0.19541f
C448 B.t6 VSUBS 0.554227f
C449 B.n230 VSUBS 0.121846f
C450 B.n231 VSUBS 0.084541f
C451 B.n232 VSUBS 0.020369f
C452 B.n233 VSUBS 0.008275f
C453 B.n234 VSUBS 0.008792f
C454 B.n235 VSUBS 0.008792f
C455 B.n236 VSUBS 0.008792f
C456 B.n237 VSUBS 0.008792f
C457 B.n238 VSUBS 0.008792f
C458 B.n239 VSUBS 0.008792f
C459 B.n240 VSUBS 0.008792f
C460 B.n241 VSUBS 0.008792f
C461 B.n242 VSUBS 0.008792f
C462 B.n243 VSUBS 0.008792f
C463 B.n244 VSUBS 0.008792f
C464 B.n245 VSUBS 0.008792f
C465 B.n246 VSUBS 0.008792f
C466 B.n247 VSUBS 0.008792f
C467 B.n248 VSUBS 0.008792f
C468 B.n249 VSUBS 0.004913f
C469 B.n250 VSUBS 0.020369f
C470 B.n251 VSUBS 0.008275f
C471 B.n252 VSUBS 0.008792f
C472 B.n253 VSUBS 0.008792f
C473 B.n254 VSUBS 0.008792f
C474 B.n255 VSUBS 0.008792f
C475 B.n256 VSUBS 0.008792f
C476 B.n257 VSUBS 0.008792f
C477 B.n258 VSUBS 0.008792f
C478 B.n259 VSUBS 0.008792f
C479 B.n260 VSUBS 0.008792f
C480 B.n261 VSUBS 0.008792f
C481 B.n262 VSUBS 0.008792f
C482 B.n263 VSUBS 0.008792f
C483 B.n264 VSUBS 0.008792f
C484 B.n265 VSUBS 0.008792f
C485 B.n266 VSUBS 0.008792f
C486 B.n267 VSUBS 0.008792f
C487 B.n268 VSUBS 0.008792f
C488 B.n269 VSUBS 0.008792f
C489 B.n270 VSUBS 0.008792f
C490 B.n271 VSUBS 0.008792f
C491 B.n272 VSUBS 0.008792f
C492 B.n273 VSUBS 0.008792f
C493 B.n274 VSUBS 0.008792f
C494 B.n275 VSUBS 0.008792f
C495 B.n276 VSUBS 0.008792f
C496 B.n277 VSUBS 0.008792f
C497 B.n278 VSUBS 0.008792f
C498 B.n279 VSUBS 0.008792f
C499 B.n280 VSUBS 0.008792f
C500 B.n281 VSUBS 0.019391f
C501 B.n282 VSUBS 0.02043f
C502 B.n283 VSUBS 0.019338f
C503 B.n284 VSUBS 0.008792f
C504 B.n285 VSUBS 0.008792f
C505 B.n286 VSUBS 0.008792f
C506 B.n287 VSUBS 0.008792f
C507 B.n288 VSUBS 0.008792f
C508 B.n289 VSUBS 0.008792f
C509 B.n290 VSUBS 0.008792f
C510 B.n291 VSUBS 0.008792f
C511 B.n292 VSUBS 0.008792f
C512 B.n293 VSUBS 0.008792f
C513 B.n294 VSUBS 0.008792f
C514 B.n295 VSUBS 0.008792f
C515 B.n296 VSUBS 0.008792f
C516 B.n297 VSUBS 0.008792f
C517 B.n298 VSUBS 0.008792f
C518 B.n299 VSUBS 0.008792f
C519 B.n300 VSUBS 0.008792f
C520 B.n301 VSUBS 0.008792f
C521 B.n302 VSUBS 0.008792f
C522 B.n303 VSUBS 0.008792f
C523 B.n304 VSUBS 0.008792f
C524 B.n305 VSUBS 0.008792f
C525 B.n306 VSUBS 0.008792f
C526 B.n307 VSUBS 0.008792f
C527 B.n308 VSUBS 0.008792f
C528 B.n309 VSUBS 0.008792f
C529 B.n310 VSUBS 0.008792f
C530 B.n311 VSUBS 0.008792f
C531 B.n312 VSUBS 0.008792f
C532 B.n313 VSUBS 0.008792f
C533 B.n314 VSUBS 0.008792f
C534 B.n315 VSUBS 0.008792f
C535 B.n316 VSUBS 0.008792f
C536 B.n317 VSUBS 0.008792f
C537 B.n318 VSUBS 0.008792f
C538 B.n319 VSUBS 0.008792f
C539 B.n320 VSUBS 0.008792f
C540 B.n321 VSUBS 0.008792f
C541 B.n322 VSUBS 0.008792f
C542 B.n323 VSUBS 0.008792f
C543 B.n324 VSUBS 0.008792f
C544 B.n325 VSUBS 0.008792f
C545 B.n326 VSUBS 0.008792f
C546 B.n327 VSUBS 0.008792f
C547 B.n328 VSUBS 0.008792f
C548 B.n329 VSUBS 0.008792f
C549 B.n330 VSUBS 0.008792f
C550 B.n331 VSUBS 0.008792f
C551 B.n332 VSUBS 0.008792f
C552 B.n333 VSUBS 0.008792f
C553 B.n334 VSUBS 0.008792f
C554 B.n335 VSUBS 0.008792f
C555 B.n336 VSUBS 0.008792f
C556 B.n337 VSUBS 0.008792f
C557 B.n338 VSUBS 0.008792f
C558 B.n339 VSUBS 0.008792f
C559 B.n340 VSUBS 0.008792f
C560 B.n341 VSUBS 0.008792f
C561 B.n342 VSUBS 0.008792f
C562 B.n343 VSUBS 0.008792f
C563 B.n344 VSUBS 0.008792f
C564 B.n345 VSUBS 0.008792f
C565 B.n346 VSUBS 0.008792f
C566 B.n347 VSUBS 0.008792f
C567 B.n348 VSUBS 0.008792f
C568 B.n349 VSUBS 0.008792f
C569 B.n350 VSUBS 0.008792f
C570 B.n351 VSUBS 0.008792f
C571 B.n352 VSUBS 0.008792f
C572 B.n353 VSUBS 0.008792f
C573 B.n354 VSUBS 0.008792f
C574 B.n355 VSUBS 0.008792f
C575 B.n356 VSUBS 0.008792f
C576 B.n357 VSUBS 0.008792f
C577 B.n358 VSUBS 0.008792f
C578 B.n359 VSUBS 0.008792f
C579 B.n360 VSUBS 0.008792f
C580 B.n361 VSUBS 0.008792f
C581 B.n362 VSUBS 0.008792f
C582 B.n363 VSUBS 0.008792f
C583 B.n364 VSUBS 0.008792f
C584 B.n365 VSUBS 0.008792f
C585 B.n366 VSUBS 0.008792f
C586 B.n367 VSUBS 0.008792f
C587 B.n368 VSUBS 0.008792f
C588 B.n369 VSUBS 0.008792f
C589 B.n370 VSUBS 0.008792f
C590 B.n371 VSUBS 0.008792f
C591 B.n372 VSUBS 0.008792f
C592 B.n373 VSUBS 0.008792f
C593 B.n374 VSUBS 0.008792f
C594 B.n375 VSUBS 0.008792f
C595 B.n376 VSUBS 0.008792f
C596 B.n377 VSUBS 0.008792f
C597 B.n378 VSUBS 0.008792f
C598 B.n379 VSUBS 0.008792f
C599 B.n380 VSUBS 0.008792f
C600 B.n381 VSUBS 0.008792f
C601 B.n382 VSUBS 0.008792f
C602 B.n383 VSUBS 0.008792f
C603 B.n384 VSUBS 0.008792f
C604 B.n385 VSUBS 0.008792f
C605 B.n386 VSUBS 0.008792f
C606 B.n387 VSUBS 0.008792f
C607 B.n388 VSUBS 0.008792f
C608 B.n389 VSUBS 0.008792f
C609 B.n390 VSUBS 0.008792f
C610 B.n391 VSUBS 0.008792f
C611 B.n392 VSUBS 0.008792f
C612 B.n393 VSUBS 0.008792f
C613 B.n394 VSUBS 0.008792f
C614 B.n395 VSUBS 0.008792f
C615 B.n396 VSUBS 0.008792f
C616 B.n397 VSUBS 0.008792f
C617 B.n398 VSUBS 0.008792f
C618 B.n399 VSUBS 0.008792f
C619 B.n400 VSUBS 0.008792f
C620 B.n401 VSUBS 0.008792f
C621 B.n402 VSUBS 0.008792f
C622 B.n403 VSUBS 0.008792f
C623 B.n404 VSUBS 0.019338f
C624 B.n405 VSUBS 0.020483f
C625 B.n406 VSUBS 0.020483f
C626 B.n407 VSUBS 0.008792f
C627 B.n408 VSUBS 0.008792f
C628 B.n409 VSUBS 0.008792f
C629 B.n410 VSUBS 0.008792f
C630 B.n411 VSUBS 0.008792f
C631 B.n412 VSUBS 0.008792f
C632 B.n413 VSUBS 0.008792f
C633 B.n414 VSUBS 0.008792f
C634 B.n415 VSUBS 0.008792f
C635 B.n416 VSUBS 0.008792f
C636 B.n417 VSUBS 0.008792f
C637 B.n418 VSUBS 0.008792f
C638 B.n419 VSUBS 0.008792f
C639 B.n420 VSUBS 0.008792f
C640 B.n421 VSUBS 0.008792f
C641 B.n422 VSUBS 0.008792f
C642 B.n423 VSUBS 0.008792f
C643 B.n424 VSUBS 0.008792f
C644 B.n425 VSUBS 0.008792f
C645 B.n426 VSUBS 0.008792f
C646 B.n427 VSUBS 0.008792f
C647 B.n428 VSUBS 0.008792f
C648 B.n429 VSUBS 0.008792f
C649 B.n430 VSUBS 0.008792f
C650 B.n431 VSUBS 0.008792f
C651 B.n432 VSUBS 0.008792f
C652 B.n433 VSUBS 0.008792f
C653 B.n434 VSUBS 0.008792f
C654 B.n435 VSUBS 0.008792f
C655 B.n436 VSUBS 0.008275f
C656 B.n437 VSUBS 0.020369f
C657 B.n438 VSUBS 0.004913f
C658 B.n439 VSUBS 0.008792f
C659 B.n440 VSUBS 0.008792f
C660 B.n441 VSUBS 0.008792f
C661 B.n442 VSUBS 0.008792f
C662 B.n443 VSUBS 0.008792f
C663 B.n444 VSUBS 0.008792f
C664 B.n445 VSUBS 0.008792f
C665 B.n446 VSUBS 0.008792f
C666 B.n447 VSUBS 0.008792f
C667 B.n448 VSUBS 0.008792f
C668 B.n449 VSUBS 0.008792f
C669 B.n450 VSUBS 0.008792f
C670 B.n451 VSUBS 0.004913f
C671 B.n452 VSUBS 0.008792f
C672 B.n453 VSUBS 0.008792f
C673 B.n454 VSUBS 0.008792f
C674 B.n455 VSUBS 0.008792f
C675 B.n456 VSUBS 0.008792f
C676 B.n457 VSUBS 0.008792f
C677 B.n458 VSUBS 0.008792f
C678 B.n459 VSUBS 0.008792f
C679 B.n460 VSUBS 0.008792f
C680 B.n461 VSUBS 0.008792f
C681 B.n462 VSUBS 0.008792f
C682 B.n463 VSUBS 0.008792f
C683 B.n464 VSUBS 0.008792f
C684 B.n465 VSUBS 0.008792f
C685 B.n466 VSUBS 0.008792f
C686 B.n467 VSUBS 0.008792f
C687 B.n468 VSUBS 0.008792f
C688 B.n469 VSUBS 0.008792f
C689 B.n470 VSUBS 0.008792f
C690 B.n471 VSUBS 0.008792f
C691 B.n472 VSUBS 0.008792f
C692 B.n473 VSUBS 0.008792f
C693 B.n474 VSUBS 0.008792f
C694 B.n475 VSUBS 0.008792f
C695 B.n476 VSUBS 0.008792f
C696 B.n477 VSUBS 0.008792f
C697 B.n478 VSUBS 0.008792f
C698 B.n479 VSUBS 0.008792f
C699 B.n480 VSUBS 0.008792f
C700 B.n481 VSUBS 0.008792f
C701 B.n482 VSUBS 0.008792f
C702 B.n483 VSUBS 0.020483f
C703 B.n484 VSUBS 0.019338f
C704 B.n485 VSUBS 0.019338f
C705 B.n486 VSUBS 0.008792f
C706 B.n487 VSUBS 0.008792f
C707 B.n488 VSUBS 0.008792f
C708 B.n489 VSUBS 0.008792f
C709 B.n490 VSUBS 0.008792f
C710 B.n491 VSUBS 0.008792f
C711 B.n492 VSUBS 0.008792f
C712 B.n493 VSUBS 0.008792f
C713 B.n494 VSUBS 0.008792f
C714 B.n495 VSUBS 0.008792f
C715 B.n496 VSUBS 0.008792f
C716 B.n497 VSUBS 0.008792f
C717 B.n498 VSUBS 0.008792f
C718 B.n499 VSUBS 0.008792f
C719 B.n500 VSUBS 0.008792f
C720 B.n501 VSUBS 0.008792f
C721 B.n502 VSUBS 0.008792f
C722 B.n503 VSUBS 0.008792f
C723 B.n504 VSUBS 0.008792f
C724 B.n505 VSUBS 0.008792f
C725 B.n506 VSUBS 0.008792f
C726 B.n507 VSUBS 0.008792f
C727 B.n508 VSUBS 0.008792f
C728 B.n509 VSUBS 0.008792f
C729 B.n510 VSUBS 0.008792f
C730 B.n511 VSUBS 0.008792f
C731 B.n512 VSUBS 0.008792f
C732 B.n513 VSUBS 0.008792f
C733 B.n514 VSUBS 0.008792f
C734 B.n515 VSUBS 0.008792f
C735 B.n516 VSUBS 0.008792f
C736 B.n517 VSUBS 0.008792f
C737 B.n518 VSUBS 0.008792f
C738 B.n519 VSUBS 0.008792f
C739 B.n520 VSUBS 0.008792f
C740 B.n521 VSUBS 0.008792f
C741 B.n522 VSUBS 0.008792f
C742 B.n523 VSUBS 0.008792f
C743 B.n524 VSUBS 0.008792f
C744 B.n525 VSUBS 0.008792f
C745 B.n526 VSUBS 0.008792f
C746 B.n527 VSUBS 0.008792f
C747 B.n528 VSUBS 0.008792f
C748 B.n529 VSUBS 0.008792f
C749 B.n530 VSUBS 0.008792f
C750 B.n531 VSUBS 0.008792f
C751 B.n532 VSUBS 0.008792f
C752 B.n533 VSUBS 0.008792f
C753 B.n534 VSUBS 0.008792f
C754 B.n535 VSUBS 0.008792f
C755 B.n536 VSUBS 0.008792f
C756 B.n537 VSUBS 0.008792f
C757 B.n538 VSUBS 0.008792f
C758 B.n539 VSUBS 0.008792f
C759 B.n540 VSUBS 0.008792f
C760 B.n541 VSUBS 0.008792f
C761 B.n542 VSUBS 0.008792f
C762 B.n543 VSUBS 0.011473f
C763 B.n544 VSUBS 0.012221f
C764 B.n545 VSUBS 0.024303f
.ends

