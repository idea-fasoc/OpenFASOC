* NGSPICE file created from diff_pair_sample_0969.ext - technology: sky130A

.subckt diff_pair_sample_0969 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=1.3926 pd=8.77 as=1.3926 ps=8.77 w=8.44 l=1.11
X1 VTAIL.t5 VN.t0 VDD2.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=1.3926 pd=8.77 as=1.3926 ps=8.77 w=8.44 l=1.11
X2 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=3.2916 pd=17.66 as=0 ps=0 w=8.44 l=1.11
X3 VDD2.t6 VN.t1 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.3926 pd=8.77 as=1.3926 ps=8.77 w=8.44 l=1.11
X4 VTAIL.t9 VP.t1 VDD1.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3926 pd=8.77 as=1.3926 ps=8.77 w=8.44 l=1.11
X5 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=3.2916 pd=17.66 as=0 ps=0 w=8.44 l=1.11
X6 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=3.2916 pd=17.66 as=0 ps=0 w=8.44 l=1.11
X7 VTAIL.t13 VP.t2 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=3.2916 pd=17.66 as=1.3926 ps=8.77 w=8.44 l=1.11
X8 VDD2.t5 VN.t2 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.3926 pd=8.77 as=3.2916 ps=17.66 w=8.44 l=1.11
X9 VDD2.t4 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3926 pd=8.77 as=3.2916 ps=17.66 w=8.44 l=1.11
X10 VTAIL.t0 VN.t4 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3926 pd=8.77 as=1.3926 ps=8.77 w=8.44 l=1.11
X11 VDD1.t4 VP.t3 VTAIL.t12 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3926 pd=8.77 as=3.2916 ps=17.66 w=8.44 l=1.11
X12 VDD2.t2 VN.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.3926 pd=8.77 as=1.3926 ps=8.77 w=8.44 l=1.11
X13 VTAIL.t1 VN.t6 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2916 pd=17.66 as=1.3926 ps=8.77 w=8.44 l=1.11
X14 VDD1.t3 VP.t4 VTAIL.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.3926 pd=8.77 as=3.2916 ps=17.66 w=8.44 l=1.11
X15 VDD1.t2 VP.t5 VTAIL.t15 B.t6 sky130_fd_pr__nfet_01v8 ad=1.3926 pd=8.77 as=1.3926 ps=8.77 w=8.44 l=1.11
X16 VTAIL.t14 VP.t6 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2916 pd=17.66 as=1.3926 ps=8.77 w=8.44 l=1.11
X17 VTAIL.t2 VN.t7 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=3.2916 pd=17.66 as=1.3926 ps=8.77 w=8.44 l=1.11
X18 VTAIL.t11 VP.t7 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=1.3926 pd=8.77 as=1.3926 ps=8.77 w=8.44 l=1.11
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.2916 pd=17.66 as=0 ps=0 w=8.44 l=1.11
R0 VP.n7 VP.t6 241.387
R1 VP.n17 VP.t2 218.637
R2 VP.n29 VP.t3 218.637
R3 VP.n15 VP.t4 218.637
R4 VP.n22 VP.t0 183.248
R5 VP.n1 VP.t1 183.248
R6 VP.n5 VP.t7 183.248
R7 VP.n8 VP.t5 183.248
R8 VP.n9 VP.n6 161.3
R9 VP.n11 VP.n10 161.3
R10 VP.n13 VP.n12 161.3
R11 VP.n14 VP.n4 161.3
R12 VP.n28 VP.n0 161.3
R13 VP.n27 VP.n26 161.3
R14 VP.n25 VP.n24 161.3
R15 VP.n23 VP.n2 161.3
R16 VP.n21 VP.n20 161.3
R17 VP.n19 VP.n3 161.3
R18 VP.n16 VP.n15 80.6037
R19 VP.n30 VP.n29 80.6037
R20 VP.n18 VP.n17 80.6037
R21 VP.n24 VP.n23 56.5617
R22 VP.n10 VP.n9 56.5617
R23 VP.n17 VP.n3 49.4301
R24 VP.n29 VP.n28 49.4301
R25 VP.n15 VP.n14 49.4301
R26 VP.n18 VP.n16 41.4029
R27 VP.n8 VP.n7 33.9241
R28 VP.n7 VP.n6 28.263
R29 VP.n21 VP.n3 24.5923
R30 VP.n28 VP.n27 24.5923
R31 VP.n14 VP.n13 24.5923
R32 VP.n23 VP.n22 23.1168
R33 VP.n24 VP.n1 23.1168
R34 VP.n10 VP.n5 23.1168
R35 VP.n9 VP.n8 23.1168
R36 VP.n22 VP.n21 1.47601
R37 VP.n27 VP.n1 1.47601
R38 VP.n13 VP.n5 1.47601
R39 VP.n16 VP.n4 0.285035
R40 VP.n19 VP.n18 0.285035
R41 VP.n30 VP.n0 0.285035
R42 VP.n11 VP.n6 0.189894
R43 VP.n12 VP.n11 0.189894
R44 VP.n12 VP.n4 0.189894
R45 VP.n20 VP.n19 0.189894
R46 VP.n20 VP.n2 0.189894
R47 VP.n25 VP.n2 0.189894
R48 VP.n26 VP.n25 0.189894
R49 VP.n26 VP.n0 0.189894
R50 VP VP.n30 0.146778
R51 VTAIL.n11 VTAIL.t14 48.3217
R52 VTAIL.n10 VTAIL.t3 48.3217
R53 VTAIL.n7 VTAIL.t2 48.3217
R54 VTAIL.n14 VTAIL.t8 48.3217
R55 VTAIL.n15 VTAIL.t7 48.3215
R56 VTAIL.n2 VTAIL.t1 48.3215
R57 VTAIL.n3 VTAIL.t12 48.3215
R58 VTAIL.n6 VTAIL.t13 48.3215
R59 VTAIL.n13 VTAIL.n12 45.9758
R60 VTAIL.n9 VTAIL.n8 45.9758
R61 VTAIL.n1 VTAIL.n0 45.9757
R62 VTAIL.n5 VTAIL.n4 45.9757
R63 VTAIL.n15 VTAIL.n14 20.8841
R64 VTAIL.n7 VTAIL.n6 20.8841
R65 VTAIL.n0 VTAIL.t6 2.34647
R66 VTAIL.n0 VTAIL.t5 2.34647
R67 VTAIL.n4 VTAIL.t10 2.34647
R68 VTAIL.n4 VTAIL.t9 2.34647
R69 VTAIL.n12 VTAIL.t15 2.34647
R70 VTAIL.n12 VTAIL.t11 2.34647
R71 VTAIL.n8 VTAIL.t4 2.34647
R72 VTAIL.n8 VTAIL.t0 2.34647
R73 VTAIL.n9 VTAIL.n7 1.24188
R74 VTAIL.n10 VTAIL.n9 1.24188
R75 VTAIL.n13 VTAIL.n11 1.24188
R76 VTAIL.n14 VTAIL.n13 1.24188
R77 VTAIL.n6 VTAIL.n5 1.24188
R78 VTAIL.n5 VTAIL.n3 1.24188
R79 VTAIL.n2 VTAIL.n1 1.24188
R80 VTAIL VTAIL.n15 1.18369
R81 VTAIL.n11 VTAIL.n10 0.470328
R82 VTAIL.n3 VTAIL.n2 0.470328
R83 VTAIL VTAIL.n1 0.0586897
R84 VDD1 VDD1.n0 63.3334
R85 VDD1.n3 VDD1.n2 63.2199
R86 VDD1.n3 VDD1.n1 63.2199
R87 VDD1.n5 VDD1.n4 62.6545
R88 VDD1.n5 VDD1.n3 37.1604
R89 VDD1.n4 VDD1.t0 2.34647
R90 VDD1.n4 VDD1.t3 2.34647
R91 VDD1.n0 VDD1.t1 2.34647
R92 VDD1.n0 VDD1.t2 2.34647
R93 VDD1.n2 VDD1.t6 2.34647
R94 VDD1.n2 VDD1.t4 2.34647
R95 VDD1.n1 VDD1.t5 2.34647
R96 VDD1.n1 VDD1.t7 2.34647
R97 VDD1 VDD1.n5 0.563
R98 B.n605 B.n604 585
R99 B.n238 B.n91 585
R100 B.n237 B.n236 585
R101 B.n235 B.n234 585
R102 B.n233 B.n232 585
R103 B.n231 B.n230 585
R104 B.n229 B.n228 585
R105 B.n227 B.n226 585
R106 B.n225 B.n224 585
R107 B.n223 B.n222 585
R108 B.n221 B.n220 585
R109 B.n219 B.n218 585
R110 B.n217 B.n216 585
R111 B.n215 B.n214 585
R112 B.n213 B.n212 585
R113 B.n211 B.n210 585
R114 B.n209 B.n208 585
R115 B.n207 B.n206 585
R116 B.n205 B.n204 585
R117 B.n203 B.n202 585
R118 B.n201 B.n200 585
R119 B.n199 B.n198 585
R120 B.n197 B.n196 585
R121 B.n195 B.n194 585
R122 B.n193 B.n192 585
R123 B.n191 B.n190 585
R124 B.n189 B.n188 585
R125 B.n187 B.n186 585
R126 B.n185 B.n184 585
R127 B.n183 B.n182 585
R128 B.n181 B.n180 585
R129 B.n178 B.n177 585
R130 B.n176 B.n175 585
R131 B.n174 B.n173 585
R132 B.n172 B.n171 585
R133 B.n170 B.n169 585
R134 B.n168 B.n167 585
R135 B.n166 B.n165 585
R136 B.n164 B.n163 585
R137 B.n162 B.n161 585
R138 B.n160 B.n159 585
R139 B.n157 B.n156 585
R140 B.n155 B.n154 585
R141 B.n153 B.n152 585
R142 B.n151 B.n150 585
R143 B.n149 B.n148 585
R144 B.n147 B.n146 585
R145 B.n145 B.n144 585
R146 B.n143 B.n142 585
R147 B.n141 B.n140 585
R148 B.n139 B.n138 585
R149 B.n137 B.n136 585
R150 B.n135 B.n134 585
R151 B.n133 B.n132 585
R152 B.n131 B.n130 585
R153 B.n129 B.n128 585
R154 B.n127 B.n126 585
R155 B.n125 B.n124 585
R156 B.n123 B.n122 585
R157 B.n121 B.n120 585
R158 B.n119 B.n118 585
R159 B.n117 B.n116 585
R160 B.n115 B.n114 585
R161 B.n113 B.n112 585
R162 B.n111 B.n110 585
R163 B.n109 B.n108 585
R164 B.n107 B.n106 585
R165 B.n105 B.n104 585
R166 B.n103 B.n102 585
R167 B.n101 B.n100 585
R168 B.n99 B.n98 585
R169 B.n97 B.n96 585
R170 B.n603 B.n55 585
R171 B.n608 B.n55 585
R172 B.n602 B.n54 585
R173 B.n609 B.n54 585
R174 B.n601 B.n600 585
R175 B.n600 B.n50 585
R176 B.n599 B.n49 585
R177 B.n615 B.n49 585
R178 B.n598 B.n48 585
R179 B.n616 B.n48 585
R180 B.n597 B.n47 585
R181 B.n617 B.n47 585
R182 B.n596 B.n595 585
R183 B.n595 B.n43 585
R184 B.n594 B.n42 585
R185 B.n623 B.n42 585
R186 B.n593 B.n41 585
R187 B.n624 B.n41 585
R188 B.n592 B.n40 585
R189 B.n625 B.n40 585
R190 B.n591 B.n590 585
R191 B.n590 B.n36 585
R192 B.n589 B.n35 585
R193 B.n631 B.n35 585
R194 B.n588 B.n34 585
R195 B.n632 B.n34 585
R196 B.n587 B.n33 585
R197 B.n633 B.n33 585
R198 B.n586 B.n585 585
R199 B.n585 B.n29 585
R200 B.n584 B.n28 585
R201 B.n639 B.n28 585
R202 B.n583 B.n27 585
R203 B.n640 B.n27 585
R204 B.n582 B.n26 585
R205 B.n641 B.n26 585
R206 B.n581 B.n580 585
R207 B.n580 B.n22 585
R208 B.n579 B.n21 585
R209 B.n647 B.n21 585
R210 B.n578 B.n20 585
R211 B.n648 B.n20 585
R212 B.n577 B.n19 585
R213 B.n649 B.n19 585
R214 B.n576 B.n575 585
R215 B.n575 B.n15 585
R216 B.n574 B.n14 585
R217 B.n655 B.n14 585
R218 B.n573 B.n13 585
R219 B.n656 B.n13 585
R220 B.n572 B.n12 585
R221 B.n657 B.n12 585
R222 B.n571 B.n570 585
R223 B.n570 B.n8 585
R224 B.n569 B.n7 585
R225 B.n663 B.n7 585
R226 B.n568 B.n6 585
R227 B.n664 B.n6 585
R228 B.n567 B.n5 585
R229 B.n665 B.n5 585
R230 B.n566 B.n565 585
R231 B.n565 B.n4 585
R232 B.n564 B.n239 585
R233 B.n564 B.n563 585
R234 B.n554 B.n240 585
R235 B.n241 B.n240 585
R236 B.n556 B.n555 585
R237 B.n557 B.n556 585
R238 B.n553 B.n246 585
R239 B.n246 B.n245 585
R240 B.n552 B.n551 585
R241 B.n551 B.n550 585
R242 B.n248 B.n247 585
R243 B.n249 B.n248 585
R244 B.n543 B.n542 585
R245 B.n544 B.n543 585
R246 B.n541 B.n254 585
R247 B.n254 B.n253 585
R248 B.n540 B.n539 585
R249 B.n539 B.n538 585
R250 B.n256 B.n255 585
R251 B.n257 B.n256 585
R252 B.n531 B.n530 585
R253 B.n532 B.n531 585
R254 B.n529 B.n261 585
R255 B.n265 B.n261 585
R256 B.n528 B.n527 585
R257 B.n527 B.n526 585
R258 B.n263 B.n262 585
R259 B.n264 B.n263 585
R260 B.n519 B.n518 585
R261 B.n520 B.n519 585
R262 B.n517 B.n269 585
R263 B.n273 B.n269 585
R264 B.n516 B.n515 585
R265 B.n515 B.n514 585
R266 B.n271 B.n270 585
R267 B.n272 B.n271 585
R268 B.n507 B.n506 585
R269 B.n508 B.n507 585
R270 B.n505 B.n278 585
R271 B.n278 B.n277 585
R272 B.n504 B.n503 585
R273 B.n503 B.n502 585
R274 B.n280 B.n279 585
R275 B.n281 B.n280 585
R276 B.n495 B.n494 585
R277 B.n496 B.n495 585
R278 B.n493 B.n286 585
R279 B.n286 B.n285 585
R280 B.n492 B.n491 585
R281 B.n491 B.n490 585
R282 B.n288 B.n287 585
R283 B.n289 B.n288 585
R284 B.n483 B.n482 585
R285 B.n484 B.n483 585
R286 B.n481 B.n294 585
R287 B.n294 B.n293 585
R288 B.n476 B.n475 585
R289 B.n474 B.n332 585
R290 B.n473 B.n331 585
R291 B.n478 B.n331 585
R292 B.n472 B.n471 585
R293 B.n470 B.n469 585
R294 B.n468 B.n467 585
R295 B.n466 B.n465 585
R296 B.n464 B.n463 585
R297 B.n462 B.n461 585
R298 B.n460 B.n459 585
R299 B.n458 B.n457 585
R300 B.n456 B.n455 585
R301 B.n454 B.n453 585
R302 B.n452 B.n451 585
R303 B.n450 B.n449 585
R304 B.n448 B.n447 585
R305 B.n446 B.n445 585
R306 B.n444 B.n443 585
R307 B.n442 B.n441 585
R308 B.n440 B.n439 585
R309 B.n438 B.n437 585
R310 B.n436 B.n435 585
R311 B.n434 B.n433 585
R312 B.n432 B.n431 585
R313 B.n430 B.n429 585
R314 B.n428 B.n427 585
R315 B.n426 B.n425 585
R316 B.n424 B.n423 585
R317 B.n422 B.n421 585
R318 B.n420 B.n419 585
R319 B.n418 B.n417 585
R320 B.n416 B.n415 585
R321 B.n414 B.n413 585
R322 B.n412 B.n411 585
R323 B.n410 B.n409 585
R324 B.n408 B.n407 585
R325 B.n406 B.n405 585
R326 B.n404 B.n403 585
R327 B.n402 B.n401 585
R328 B.n400 B.n399 585
R329 B.n398 B.n397 585
R330 B.n396 B.n395 585
R331 B.n394 B.n393 585
R332 B.n392 B.n391 585
R333 B.n390 B.n389 585
R334 B.n388 B.n387 585
R335 B.n386 B.n385 585
R336 B.n384 B.n383 585
R337 B.n382 B.n381 585
R338 B.n380 B.n379 585
R339 B.n378 B.n377 585
R340 B.n376 B.n375 585
R341 B.n374 B.n373 585
R342 B.n372 B.n371 585
R343 B.n370 B.n369 585
R344 B.n368 B.n367 585
R345 B.n366 B.n365 585
R346 B.n364 B.n363 585
R347 B.n362 B.n361 585
R348 B.n360 B.n359 585
R349 B.n358 B.n357 585
R350 B.n356 B.n355 585
R351 B.n354 B.n353 585
R352 B.n352 B.n351 585
R353 B.n350 B.n349 585
R354 B.n348 B.n347 585
R355 B.n346 B.n345 585
R356 B.n344 B.n343 585
R357 B.n342 B.n341 585
R358 B.n340 B.n339 585
R359 B.n296 B.n295 585
R360 B.n480 B.n479 585
R361 B.n479 B.n478 585
R362 B.n292 B.n291 585
R363 B.n293 B.n292 585
R364 B.n486 B.n485 585
R365 B.n485 B.n484 585
R366 B.n487 B.n290 585
R367 B.n290 B.n289 585
R368 B.n489 B.n488 585
R369 B.n490 B.n489 585
R370 B.n284 B.n283 585
R371 B.n285 B.n284 585
R372 B.n498 B.n497 585
R373 B.n497 B.n496 585
R374 B.n499 B.n282 585
R375 B.n282 B.n281 585
R376 B.n501 B.n500 585
R377 B.n502 B.n501 585
R378 B.n276 B.n275 585
R379 B.n277 B.n276 585
R380 B.n510 B.n509 585
R381 B.n509 B.n508 585
R382 B.n511 B.n274 585
R383 B.n274 B.n272 585
R384 B.n513 B.n512 585
R385 B.n514 B.n513 585
R386 B.n268 B.n267 585
R387 B.n273 B.n268 585
R388 B.n522 B.n521 585
R389 B.n521 B.n520 585
R390 B.n523 B.n266 585
R391 B.n266 B.n264 585
R392 B.n525 B.n524 585
R393 B.n526 B.n525 585
R394 B.n260 B.n259 585
R395 B.n265 B.n260 585
R396 B.n534 B.n533 585
R397 B.n533 B.n532 585
R398 B.n535 B.n258 585
R399 B.n258 B.n257 585
R400 B.n537 B.n536 585
R401 B.n538 B.n537 585
R402 B.n252 B.n251 585
R403 B.n253 B.n252 585
R404 B.n546 B.n545 585
R405 B.n545 B.n544 585
R406 B.n547 B.n250 585
R407 B.n250 B.n249 585
R408 B.n549 B.n548 585
R409 B.n550 B.n549 585
R410 B.n244 B.n243 585
R411 B.n245 B.n244 585
R412 B.n559 B.n558 585
R413 B.n558 B.n557 585
R414 B.n560 B.n242 585
R415 B.n242 B.n241 585
R416 B.n562 B.n561 585
R417 B.n563 B.n562 585
R418 B.n2 B.n0 585
R419 B.n4 B.n2 585
R420 B.n3 B.n1 585
R421 B.n664 B.n3 585
R422 B.n662 B.n661 585
R423 B.n663 B.n662 585
R424 B.n660 B.n9 585
R425 B.n9 B.n8 585
R426 B.n659 B.n658 585
R427 B.n658 B.n657 585
R428 B.n11 B.n10 585
R429 B.n656 B.n11 585
R430 B.n654 B.n653 585
R431 B.n655 B.n654 585
R432 B.n652 B.n16 585
R433 B.n16 B.n15 585
R434 B.n651 B.n650 585
R435 B.n650 B.n649 585
R436 B.n18 B.n17 585
R437 B.n648 B.n18 585
R438 B.n646 B.n645 585
R439 B.n647 B.n646 585
R440 B.n644 B.n23 585
R441 B.n23 B.n22 585
R442 B.n643 B.n642 585
R443 B.n642 B.n641 585
R444 B.n25 B.n24 585
R445 B.n640 B.n25 585
R446 B.n638 B.n637 585
R447 B.n639 B.n638 585
R448 B.n636 B.n30 585
R449 B.n30 B.n29 585
R450 B.n635 B.n634 585
R451 B.n634 B.n633 585
R452 B.n32 B.n31 585
R453 B.n632 B.n32 585
R454 B.n630 B.n629 585
R455 B.n631 B.n630 585
R456 B.n628 B.n37 585
R457 B.n37 B.n36 585
R458 B.n627 B.n626 585
R459 B.n626 B.n625 585
R460 B.n39 B.n38 585
R461 B.n624 B.n39 585
R462 B.n622 B.n621 585
R463 B.n623 B.n622 585
R464 B.n620 B.n44 585
R465 B.n44 B.n43 585
R466 B.n619 B.n618 585
R467 B.n618 B.n617 585
R468 B.n46 B.n45 585
R469 B.n616 B.n46 585
R470 B.n614 B.n613 585
R471 B.n615 B.n614 585
R472 B.n612 B.n51 585
R473 B.n51 B.n50 585
R474 B.n611 B.n610 585
R475 B.n610 B.n609 585
R476 B.n53 B.n52 585
R477 B.n608 B.n53 585
R478 B.n667 B.n666 585
R479 B.n666 B.n665 585
R480 B.n476 B.n292 535.745
R481 B.n96 B.n53 535.745
R482 B.n479 B.n294 535.745
R483 B.n605 B.n55 535.745
R484 B.n336 B.t8 386.866
R485 B.n333 B.t12 386.866
R486 B.n94 B.t15 386.866
R487 B.n92 B.t19 386.866
R488 B.n607 B.n606 256.663
R489 B.n607 B.n90 256.663
R490 B.n607 B.n89 256.663
R491 B.n607 B.n88 256.663
R492 B.n607 B.n87 256.663
R493 B.n607 B.n86 256.663
R494 B.n607 B.n85 256.663
R495 B.n607 B.n84 256.663
R496 B.n607 B.n83 256.663
R497 B.n607 B.n82 256.663
R498 B.n607 B.n81 256.663
R499 B.n607 B.n80 256.663
R500 B.n607 B.n79 256.663
R501 B.n607 B.n78 256.663
R502 B.n607 B.n77 256.663
R503 B.n607 B.n76 256.663
R504 B.n607 B.n75 256.663
R505 B.n607 B.n74 256.663
R506 B.n607 B.n73 256.663
R507 B.n607 B.n72 256.663
R508 B.n607 B.n71 256.663
R509 B.n607 B.n70 256.663
R510 B.n607 B.n69 256.663
R511 B.n607 B.n68 256.663
R512 B.n607 B.n67 256.663
R513 B.n607 B.n66 256.663
R514 B.n607 B.n65 256.663
R515 B.n607 B.n64 256.663
R516 B.n607 B.n63 256.663
R517 B.n607 B.n62 256.663
R518 B.n607 B.n61 256.663
R519 B.n607 B.n60 256.663
R520 B.n607 B.n59 256.663
R521 B.n607 B.n58 256.663
R522 B.n607 B.n57 256.663
R523 B.n607 B.n56 256.663
R524 B.n478 B.n477 256.663
R525 B.n478 B.n297 256.663
R526 B.n478 B.n298 256.663
R527 B.n478 B.n299 256.663
R528 B.n478 B.n300 256.663
R529 B.n478 B.n301 256.663
R530 B.n478 B.n302 256.663
R531 B.n478 B.n303 256.663
R532 B.n478 B.n304 256.663
R533 B.n478 B.n305 256.663
R534 B.n478 B.n306 256.663
R535 B.n478 B.n307 256.663
R536 B.n478 B.n308 256.663
R537 B.n478 B.n309 256.663
R538 B.n478 B.n310 256.663
R539 B.n478 B.n311 256.663
R540 B.n478 B.n312 256.663
R541 B.n478 B.n313 256.663
R542 B.n478 B.n314 256.663
R543 B.n478 B.n315 256.663
R544 B.n478 B.n316 256.663
R545 B.n478 B.n317 256.663
R546 B.n478 B.n318 256.663
R547 B.n478 B.n319 256.663
R548 B.n478 B.n320 256.663
R549 B.n478 B.n321 256.663
R550 B.n478 B.n322 256.663
R551 B.n478 B.n323 256.663
R552 B.n478 B.n324 256.663
R553 B.n478 B.n325 256.663
R554 B.n478 B.n326 256.663
R555 B.n478 B.n327 256.663
R556 B.n478 B.n328 256.663
R557 B.n478 B.n329 256.663
R558 B.n478 B.n330 256.663
R559 B.n485 B.n292 163.367
R560 B.n485 B.n290 163.367
R561 B.n489 B.n290 163.367
R562 B.n489 B.n284 163.367
R563 B.n497 B.n284 163.367
R564 B.n497 B.n282 163.367
R565 B.n501 B.n282 163.367
R566 B.n501 B.n276 163.367
R567 B.n509 B.n276 163.367
R568 B.n509 B.n274 163.367
R569 B.n513 B.n274 163.367
R570 B.n513 B.n268 163.367
R571 B.n521 B.n268 163.367
R572 B.n521 B.n266 163.367
R573 B.n525 B.n266 163.367
R574 B.n525 B.n260 163.367
R575 B.n533 B.n260 163.367
R576 B.n533 B.n258 163.367
R577 B.n537 B.n258 163.367
R578 B.n537 B.n252 163.367
R579 B.n545 B.n252 163.367
R580 B.n545 B.n250 163.367
R581 B.n549 B.n250 163.367
R582 B.n549 B.n244 163.367
R583 B.n558 B.n244 163.367
R584 B.n558 B.n242 163.367
R585 B.n562 B.n242 163.367
R586 B.n562 B.n2 163.367
R587 B.n666 B.n2 163.367
R588 B.n666 B.n3 163.367
R589 B.n662 B.n3 163.367
R590 B.n662 B.n9 163.367
R591 B.n658 B.n9 163.367
R592 B.n658 B.n11 163.367
R593 B.n654 B.n11 163.367
R594 B.n654 B.n16 163.367
R595 B.n650 B.n16 163.367
R596 B.n650 B.n18 163.367
R597 B.n646 B.n18 163.367
R598 B.n646 B.n23 163.367
R599 B.n642 B.n23 163.367
R600 B.n642 B.n25 163.367
R601 B.n638 B.n25 163.367
R602 B.n638 B.n30 163.367
R603 B.n634 B.n30 163.367
R604 B.n634 B.n32 163.367
R605 B.n630 B.n32 163.367
R606 B.n630 B.n37 163.367
R607 B.n626 B.n37 163.367
R608 B.n626 B.n39 163.367
R609 B.n622 B.n39 163.367
R610 B.n622 B.n44 163.367
R611 B.n618 B.n44 163.367
R612 B.n618 B.n46 163.367
R613 B.n614 B.n46 163.367
R614 B.n614 B.n51 163.367
R615 B.n610 B.n51 163.367
R616 B.n610 B.n53 163.367
R617 B.n332 B.n331 163.367
R618 B.n471 B.n331 163.367
R619 B.n469 B.n468 163.367
R620 B.n465 B.n464 163.367
R621 B.n461 B.n460 163.367
R622 B.n457 B.n456 163.367
R623 B.n453 B.n452 163.367
R624 B.n449 B.n448 163.367
R625 B.n445 B.n444 163.367
R626 B.n441 B.n440 163.367
R627 B.n437 B.n436 163.367
R628 B.n433 B.n432 163.367
R629 B.n429 B.n428 163.367
R630 B.n425 B.n424 163.367
R631 B.n421 B.n420 163.367
R632 B.n417 B.n416 163.367
R633 B.n413 B.n412 163.367
R634 B.n409 B.n408 163.367
R635 B.n405 B.n404 163.367
R636 B.n401 B.n400 163.367
R637 B.n397 B.n396 163.367
R638 B.n393 B.n392 163.367
R639 B.n389 B.n388 163.367
R640 B.n385 B.n384 163.367
R641 B.n381 B.n380 163.367
R642 B.n377 B.n376 163.367
R643 B.n373 B.n372 163.367
R644 B.n369 B.n368 163.367
R645 B.n365 B.n364 163.367
R646 B.n361 B.n360 163.367
R647 B.n357 B.n356 163.367
R648 B.n353 B.n352 163.367
R649 B.n349 B.n348 163.367
R650 B.n345 B.n344 163.367
R651 B.n341 B.n340 163.367
R652 B.n479 B.n296 163.367
R653 B.n483 B.n294 163.367
R654 B.n483 B.n288 163.367
R655 B.n491 B.n288 163.367
R656 B.n491 B.n286 163.367
R657 B.n495 B.n286 163.367
R658 B.n495 B.n280 163.367
R659 B.n503 B.n280 163.367
R660 B.n503 B.n278 163.367
R661 B.n507 B.n278 163.367
R662 B.n507 B.n271 163.367
R663 B.n515 B.n271 163.367
R664 B.n515 B.n269 163.367
R665 B.n519 B.n269 163.367
R666 B.n519 B.n263 163.367
R667 B.n527 B.n263 163.367
R668 B.n527 B.n261 163.367
R669 B.n531 B.n261 163.367
R670 B.n531 B.n256 163.367
R671 B.n539 B.n256 163.367
R672 B.n539 B.n254 163.367
R673 B.n543 B.n254 163.367
R674 B.n543 B.n248 163.367
R675 B.n551 B.n248 163.367
R676 B.n551 B.n246 163.367
R677 B.n556 B.n246 163.367
R678 B.n556 B.n240 163.367
R679 B.n564 B.n240 163.367
R680 B.n565 B.n564 163.367
R681 B.n565 B.n5 163.367
R682 B.n6 B.n5 163.367
R683 B.n7 B.n6 163.367
R684 B.n570 B.n7 163.367
R685 B.n570 B.n12 163.367
R686 B.n13 B.n12 163.367
R687 B.n14 B.n13 163.367
R688 B.n575 B.n14 163.367
R689 B.n575 B.n19 163.367
R690 B.n20 B.n19 163.367
R691 B.n21 B.n20 163.367
R692 B.n580 B.n21 163.367
R693 B.n580 B.n26 163.367
R694 B.n27 B.n26 163.367
R695 B.n28 B.n27 163.367
R696 B.n585 B.n28 163.367
R697 B.n585 B.n33 163.367
R698 B.n34 B.n33 163.367
R699 B.n35 B.n34 163.367
R700 B.n590 B.n35 163.367
R701 B.n590 B.n40 163.367
R702 B.n41 B.n40 163.367
R703 B.n42 B.n41 163.367
R704 B.n595 B.n42 163.367
R705 B.n595 B.n47 163.367
R706 B.n48 B.n47 163.367
R707 B.n49 B.n48 163.367
R708 B.n600 B.n49 163.367
R709 B.n600 B.n54 163.367
R710 B.n55 B.n54 163.367
R711 B.n100 B.n99 163.367
R712 B.n104 B.n103 163.367
R713 B.n108 B.n107 163.367
R714 B.n112 B.n111 163.367
R715 B.n116 B.n115 163.367
R716 B.n120 B.n119 163.367
R717 B.n124 B.n123 163.367
R718 B.n128 B.n127 163.367
R719 B.n132 B.n131 163.367
R720 B.n136 B.n135 163.367
R721 B.n140 B.n139 163.367
R722 B.n144 B.n143 163.367
R723 B.n148 B.n147 163.367
R724 B.n152 B.n151 163.367
R725 B.n156 B.n155 163.367
R726 B.n161 B.n160 163.367
R727 B.n165 B.n164 163.367
R728 B.n169 B.n168 163.367
R729 B.n173 B.n172 163.367
R730 B.n177 B.n176 163.367
R731 B.n182 B.n181 163.367
R732 B.n186 B.n185 163.367
R733 B.n190 B.n189 163.367
R734 B.n194 B.n193 163.367
R735 B.n198 B.n197 163.367
R736 B.n202 B.n201 163.367
R737 B.n206 B.n205 163.367
R738 B.n210 B.n209 163.367
R739 B.n214 B.n213 163.367
R740 B.n218 B.n217 163.367
R741 B.n222 B.n221 163.367
R742 B.n226 B.n225 163.367
R743 B.n230 B.n229 163.367
R744 B.n234 B.n233 163.367
R745 B.n236 B.n91 163.367
R746 B.n478 B.n293 114.692
R747 B.n608 B.n607 114.692
R748 B.n336 B.t11 101.838
R749 B.n92 B.t20 101.838
R750 B.n333 B.t14 101.829
R751 B.n94 B.t17 101.829
R752 B.n337 B.t10 73.9112
R753 B.n93 B.t21 73.9112
R754 B.n334 B.t13 73.9014
R755 B.n95 B.t18 73.9014
R756 B.n477 B.n476 71.676
R757 B.n471 B.n297 71.676
R758 B.n468 B.n298 71.676
R759 B.n464 B.n299 71.676
R760 B.n460 B.n300 71.676
R761 B.n456 B.n301 71.676
R762 B.n452 B.n302 71.676
R763 B.n448 B.n303 71.676
R764 B.n444 B.n304 71.676
R765 B.n440 B.n305 71.676
R766 B.n436 B.n306 71.676
R767 B.n432 B.n307 71.676
R768 B.n428 B.n308 71.676
R769 B.n424 B.n309 71.676
R770 B.n420 B.n310 71.676
R771 B.n416 B.n311 71.676
R772 B.n412 B.n312 71.676
R773 B.n408 B.n313 71.676
R774 B.n404 B.n314 71.676
R775 B.n400 B.n315 71.676
R776 B.n396 B.n316 71.676
R777 B.n392 B.n317 71.676
R778 B.n388 B.n318 71.676
R779 B.n384 B.n319 71.676
R780 B.n380 B.n320 71.676
R781 B.n376 B.n321 71.676
R782 B.n372 B.n322 71.676
R783 B.n368 B.n323 71.676
R784 B.n364 B.n324 71.676
R785 B.n360 B.n325 71.676
R786 B.n356 B.n326 71.676
R787 B.n352 B.n327 71.676
R788 B.n348 B.n328 71.676
R789 B.n344 B.n329 71.676
R790 B.n340 B.n330 71.676
R791 B.n96 B.n56 71.676
R792 B.n100 B.n57 71.676
R793 B.n104 B.n58 71.676
R794 B.n108 B.n59 71.676
R795 B.n112 B.n60 71.676
R796 B.n116 B.n61 71.676
R797 B.n120 B.n62 71.676
R798 B.n124 B.n63 71.676
R799 B.n128 B.n64 71.676
R800 B.n132 B.n65 71.676
R801 B.n136 B.n66 71.676
R802 B.n140 B.n67 71.676
R803 B.n144 B.n68 71.676
R804 B.n148 B.n69 71.676
R805 B.n152 B.n70 71.676
R806 B.n156 B.n71 71.676
R807 B.n161 B.n72 71.676
R808 B.n165 B.n73 71.676
R809 B.n169 B.n74 71.676
R810 B.n173 B.n75 71.676
R811 B.n177 B.n76 71.676
R812 B.n182 B.n77 71.676
R813 B.n186 B.n78 71.676
R814 B.n190 B.n79 71.676
R815 B.n194 B.n80 71.676
R816 B.n198 B.n81 71.676
R817 B.n202 B.n82 71.676
R818 B.n206 B.n83 71.676
R819 B.n210 B.n84 71.676
R820 B.n214 B.n85 71.676
R821 B.n218 B.n86 71.676
R822 B.n222 B.n87 71.676
R823 B.n226 B.n88 71.676
R824 B.n230 B.n89 71.676
R825 B.n234 B.n90 71.676
R826 B.n606 B.n91 71.676
R827 B.n606 B.n605 71.676
R828 B.n236 B.n90 71.676
R829 B.n233 B.n89 71.676
R830 B.n229 B.n88 71.676
R831 B.n225 B.n87 71.676
R832 B.n221 B.n86 71.676
R833 B.n217 B.n85 71.676
R834 B.n213 B.n84 71.676
R835 B.n209 B.n83 71.676
R836 B.n205 B.n82 71.676
R837 B.n201 B.n81 71.676
R838 B.n197 B.n80 71.676
R839 B.n193 B.n79 71.676
R840 B.n189 B.n78 71.676
R841 B.n185 B.n77 71.676
R842 B.n181 B.n76 71.676
R843 B.n176 B.n75 71.676
R844 B.n172 B.n74 71.676
R845 B.n168 B.n73 71.676
R846 B.n164 B.n72 71.676
R847 B.n160 B.n71 71.676
R848 B.n155 B.n70 71.676
R849 B.n151 B.n69 71.676
R850 B.n147 B.n68 71.676
R851 B.n143 B.n67 71.676
R852 B.n139 B.n66 71.676
R853 B.n135 B.n65 71.676
R854 B.n131 B.n64 71.676
R855 B.n127 B.n63 71.676
R856 B.n123 B.n62 71.676
R857 B.n119 B.n61 71.676
R858 B.n115 B.n60 71.676
R859 B.n111 B.n59 71.676
R860 B.n107 B.n58 71.676
R861 B.n103 B.n57 71.676
R862 B.n99 B.n56 71.676
R863 B.n477 B.n332 71.676
R864 B.n469 B.n297 71.676
R865 B.n465 B.n298 71.676
R866 B.n461 B.n299 71.676
R867 B.n457 B.n300 71.676
R868 B.n453 B.n301 71.676
R869 B.n449 B.n302 71.676
R870 B.n445 B.n303 71.676
R871 B.n441 B.n304 71.676
R872 B.n437 B.n305 71.676
R873 B.n433 B.n306 71.676
R874 B.n429 B.n307 71.676
R875 B.n425 B.n308 71.676
R876 B.n421 B.n309 71.676
R877 B.n417 B.n310 71.676
R878 B.n413 B.n311 71.676
R879 B.n409 B.n312 71.676
R880 B.n405 B.n313 71.676
R881 B.n401 B.n314 71.676
R882 B.n397 B.n315 71.676
R883 B.n393 B.n316 71.676
R884 B.n389 B.n317 71.676
R885 B.n385 B.n318 71.676
R886 B.n381 B.n319 71.676
R887 B.n377 B.n320 71.676
R888 B.n373 B.n321 71.676
R889 B.n369 B.n322 71.676
R890 B.n365 B.n323 71.676
R891 B.n361 B.n324 71.676
R892 B.n357 B.n325 71.676
R893 B.n353 B.n326 71.676
R894 B.n349 B.n327 71.676
R895 B.n345 B.n328 71.676
R896 B.n341 B.n329 71.676
R897 B.n330 B.n296 71.676
R898 B.n338 B.n337 59.5399
R899 B.n335 B.n334 59.5399
R900 B.n158 B.n95 59.5399
R901 B.n179 B.n93 59.5399
R902 B.n484 B.n293 54.5393
R903 B.n484 B.n289 54.5393
R904 B.n490 B.n289 54.5393
R905 B.n490 B.n285 54.5393
R906 B.n496 B.n285 54.5393
R907 B.n502 B.n281 54.5393
R908 B.n502 B.n277 54.5393
R909 B.n508 B.n277 54.5393
R910 B.n508 B.n272 54.5393
R911 B.n514 B.n272 54.5393
R912 B.n514 B.n273 54.5393
R913 B.n520 B.n264 54.5393
R914 B.n526 B.n264 54.5393
R915 B.n526 B.n265 54.5393
R916 B.n532 B.n257 54.5393
R917 B.n538 B.n257 54.5393
R918 B.n538 B.n253 54.5393
R919 B.n544 B.n253 54.5393
R920 B.n550 B.n249 54.5393
R921 B.n550 B.n245 54.5393
R922 B.n557 B.n245 54.5393
R923 B.n563 B.n241 54.5393
R924 B.n563 B.n4 54.5393
R925 B.n665 B.n4 54.5393
R926 B.n665 B.n664 54.5393
R927 B.n664 B.n663 54.5393
R928 B.n663 B.n8 54.5393
R929 B.n657 B.n656 54.5393
R930 B.n656 B.n655 54.5393
R931 B.n655 B.n15 54.5393
R932 B.n649 B.n648 54.5393
R933 B.n648 B.n647 54.5393
R934 B.n647 B.n22 54.5393
R935 B.n641 B.n22 54.5393
R936 B.n640 B.n639 54.5393
R937 B.n639 B.n29 54.5393
R938 B.n633 B.n29 54.5393
R939 B.n632 B.n631 54.5393
R940 B.n631 B.n36 54.5393
R941 B.n625 B.n36 54.5393
R942 B.n625 B.n624 54.5393
R943 B.n624 B.n623 54.5393
R944 B.n623 B.n43 54.5393
R945 B.n617 B.n616 54.5393
R946 B.n616 B.n615 54.5393
R947 B.n615 B.n50 54.5393
R948 B.n609 B.n50 54.5393
R949 B.n609 B.n608 54.5393
R950 B.t0 B.n249 52.1332
R951 B.t6 B.n15 52.1332
R952 B.t9 B.n281 47.321
R953 B.t16 B.n43 47.321
R954 B.n265 B.t4 44.1128
R955 B.t5 B.n640 44.1128
R956 B.t3 B.n241 39.3005
R957 B.t1 B.n8 39.3005
R958 B.n97 B.n52 34.8103
R959 B.n604 B.n603 34.8103
R960 B.n481 B.n480 34.8103
R961 B.n475 B.n291 34.8103
R962 B.n273 B.t2 31.2801
R963 B.t7 B.n632 31.2801
R964 B.n337 B.n336 27.9278
R965 B.n334 B.n333 27.9278
R966 B.n95 B.n94 27.9278
R967 B.n93 B.n92 27.9278
R968 B.n520 B.t2 23.2597
R969 B.n633 B.t7 23.2597
R970 B B.n667 18.0485
R971 B.n557 B.t3 15.2393
R972 B.n657 B.t1 15.2393
R973 B.n98 B.n97 10.6151
R974 B.n101 B.n98 10.6151
R975 B.n102 B.n101 10.6151
R976 B.n105 B.n102 10.6151
R977 B.n106 B.n105 10.6151
R978 B.n109 B.n106 10.6151
R979 B.n110 B.n109 10.6151
R980 B.n113 B.n110 10.6151
R981 B.n114 B.n113 10.6151
R982 B.n117 B.n114 10.6151
R983 B.n118 B.n117 10.6151
R984 B.n121 B.n118 10.6151
R985 B.n122 B.n121 10.6151
R986 B.n125 B.n122 10.6151
R987 B.n126 B.n125 10.6151
R988 B.n129 B.n126 10.6151
R989 B.n130 B.n129 10.6151
R990 B.n133 B.n130 10.6151
R991 B.n134 B.n133 10.6151
R992 B.n137 B.n134 10.6151
R993 B.n138 B.n137 10.6151
R994 B.n141 B.n138 10.6151
R995 B.n142 B.n141 10.6151
R996 B.n145 B.n142 10.6151
R997 B.n146 B.n145 10.6151
R998 B.n149 B.n146 10.6151
R999 B.n150 B.n149 10.6151
R1000 B.n153 B.n150 10.6151
R1001 B.n154 B.n153 10.6151
R1002 B.n157 B.n154 10.6151
R1003 B.n162 B.n159 10.6151
R1004 B.n163 B.n162 10.6151
R1005 B.n166 B.n163 10.6151
R1006 B.n167 B.n166 10.6151
R1007 B.n170 B.n167 10.6151
R1008 B.n171 B.n170 10.6151
R1009 B.n174 B.n171 10.6151
R1010 B.n175 B.n174 10.6151
R1011 B.n178 B.n175 10.6151
R1012 B.n183 B.n180 10.6151
R1013 B.n184 B.n183 10.6151
R1014 B.n187 B.n184 10.6151
R1015 B.n188 B.n187 10.6151
R1016 B.n191 B.n188 10.6151
R1017 B.n192 B.n191 10.6151
R1018 B.n195 B.n192 10.6151
R1019 B.n196 B.n195 10.6151
R1020 B.n199 B.n196 10.6151
R1021 B.n200 B.n199 10.6151
R1022 B.n203 B.n200 10.6151
R1023 B.n204 B.n203 10.6151
R1024 B.n207 B.n204 10.6151
R1025 B.n208 B.n207 10.6151
R1026 B.n211 B.n208 10.6151
R1027 B.n212 B.n211 10.6151
R1028 B.n215 B.n212 10.6151
R1029 B.n216 B.n215 10.6151
R1030 B.n219 B.n216 10.6151
R1031 B.n220 B.n219 10.6151
R1032 B.n223 B.n220 10.6151
R1033 B.n224 B.n223 10.6151
R1034 B.n227 B.n224 10.6151
R1035 B.n228 B.n227 10.6151
R1036 B.n231 B.n228 10.6151
R1037 B.n232 B.n231 10.6151
R1038 B.n235 B.n232 10.6151
R1039 B.n237 B.n235 10.6151
R1040 B.n238 B.n237 10.6151
R1041 B.n604 B.n238 10.6151
R1042 B.n482 B.n481 10.6151
R1043 B.n482 B.n287 10.6151
R1044 B.n492 B.n287 10.6151
R1045 B.n493 B.n492 10.6151
R1046 B.n494 B.n493 10.6151
R1047 B.n494 B.n279 10.6151
R1048 B.n504 B.n279 10.6151
R1049 B.n505 B.n504 10.6151
R1050 B.n506 B.n505 10.6151
R1051 B.n506 B.n270 10.6151
R1052 B.n516 B.n270 10.6151
R1053 B.n517 B.n516 10.6151
R1054 B.n518 B.n517 10.6151
R1055 B.n518 B.n262 10.6151
R1056 B.n528 B.n262 10.6151
R1057 B.n529 B.n528 10.6151
R1058 B.n530 B.n529 10.6151
R1059 B.n530 B.n255 10.6151
R1060 B.n540 B.n255 10.6151
R1061 B.n541 B.n540 10.6151
R1062 B.n542 B.n541 10.6151
R1063 B.n542 B.n247 10.6151
R1064 B.n552 B.n247 10.6151
R1065 B.n553 B.n552 10.6151
R1066 B.n555 B.n553 10.6151
R1067 B.n555 B.n554 10.6151
R1068 B.n554 B.n239 10.6151
R1069 B.n566 B.n239 10.6151
R1070 B.n567 B.n566 10.6151
R1071 B.n568 B.n567 10.6151
R1072 B.n569 B.n568 10.6151
R1073 B.n571 B.n569 10.6151
R1074 B.n572 B.n571 10.6151
R1075 B.n573 B.n572 10.6151
R1076 B.n574 B.n573 10.6151
R1077 B.n576 B.n574 10.6151
R1078 B.n577 B.n576 10.6151
R1079 B.n578 B.n577 10.6151
R1080 B.n579 B.n578 10.6151
R1081 B.n581 B.n579 10.6151
R1082 B.n582 B.n581 10.6151
R1083 B.n583 B.n582 10.6151
R1084 B.n584 B.n583 10.6151
R1085 B.n586 B.n584 10.6151
R1086 B.n587 B.n586 10.6151
R1087 B.n588 B.n587 10.6151
R1088 B.n589 B.n588 10.6151
R1089 B.n591 B.n589 10.6151
R1090 B.n592 B.n591 10.6151
R1091 B.n593 B.n592 10.6151
R1092 B.n594 B.n593 10.6151
R1093 B.n596 B.n594 10.6151
R1094 B.n597 B.n596 10.6151
R1095 B.n598 B.n597 10.6151
R1096 B.n599 B.n598 10.6151
R1097 B.n601 B.n599 10.6151
R1098 B.n602 B.n601 10.6151
R1099 B.n603 B.n602 10.6151
R1100 B.n475 B.n474 10.6151
R1101 B.n474 B.n473 10.6151
R1102 B.n473 B.n472 10.6151
R1103 B.n472 B.n470 10.6151
R1104 B.n470 B.n467 10.6151
R1105 B.n467 B.n466 10.6151
R1106 B.n466 B.n463 10.6151
R1107 B.n463 B.n462 10.6151
R1108 B.n462 B.n459 10.6151
R1109 B.n459 B.n458 10.6151
R1110 B.n458 B.n455 10.6151
R1111 B.n455 B.n454 10.6151
R1112 B.n454 B.n451 10.6151
R1113 B.n451 B.n450 10.6151
R1114 B.n450 B.n447 10.6151
R1115 B.n447 B.n446 10.6151
R1116 B.n446 B.n443 10.6151
R1117 B.n443 B.n442 10.6151
R1118 B.n442 B.n439 10.6151
R1119 B.n439 B.n438 10.6151
R1120 B.n438 B.n435 10.6151
R1121 B.n435 B.n434 10.6151
R1122 B.n434 B.n431 10.6151
R1123 B.n431 B.n430 10.6151
R1124 B.n430 B.n427 10.6151
R1125 B.n427 B.n426 10.6151
R1126 B.n426 B.n423 10.6151
R1127 B.n423 B.n422 10.6151
R1128 B.n422 B.n419 10.6151
R1129 B.n419 B.n418 10.6151
R1130 B.n415 B.n414 10.6151
R1131 B.n414 B.n411 10.6151
R1132 B.n411 B.n410 10.6151
R1133 B.n410 B.n407 10.6151
R1134 B.n407 B.n406 10.6151
R1135 B.n406 B.n403 10.6151
R1136 B.n403 B.n402 10.6151
R1137 B.n402 B.n399 10.6151
R1138 B.n399 B.n398 10.6151
R1139 B.n395 B.n394 10.6151
R1140 B.n394 B.n391 10.6151
R1141 B.n391 B.n390 10.6151
R1142 B.n390 B.n387 10.6151
R1143 B.n387 B.n386 10.6151
R1144 B.n386 B.n383 10.6151
R1145 B.n383 B.n382 10.6151
R1146 B.n382 B.n379 10.6151
R1147 B.n379 B.n378 10.6151
R1148 B.n378 B.n375 10.6151
R1149 B.n375 B.n374 10.6151
R1150 B.n374 B.n371 10.6151
R1151 B.n371 B.n370 10.6151
R1152 B.n370 B.n367 10.6151
R1153 B.n367 B.n366 10.6151
R1154 B.n366 B.n363 10.6151
R1155 B.n363 B.n362 10.6151
R1156 B.n362 B.n359 10.6151
R1157 B.n359 B.n358 10.6151
R1158 B.n358 B.n355 10.6151
R1159 B.n355 B.n354 10.6151
R1160 B.n354 B.n351 10.6151
R1161 B.n351 B.n350 10.6151
R1162 B.n350 B.n347 10.6151
R1163 B.n347 B.n346 10.6151
R1164 B.n346 B.n343 10.6151
R1165 B.n343 B.n342 10.6151
R1166 B.n342 B.n339 10.6151
R1167 B.n339 B.n295 10.6151
R1168 B.n480 B.n295 10.6151
R1169 B.n486 B.n291 10.6151
R1170 B.n487 B.n486 10.6151
R1171 B.n488 B.n487 10.6151
R1172 B.n488 B.n283 10.6151
R1173 B.n498 B.n283 10.6151
R1174 B.n499 B.n498 10.6151
R1175 B.n500 B.n499 10.6151
R1176 B.n500 B.n275 10.6151
R1177 B.n510 B.n275 10.6151
R1178 B.n511 B.n510 10.6151
R1179 B.n512 B.n511 10.6151
R1180 B.n512 B.n267 10.6151
R1181 B.n522 B.n267 10.6151
R1182 B.n523 B.n522 10.6151
R1183 B.n524 B.n523 10.6151
R1184 B.n524 B.n259 10.6151
R1185 B.n534 B.n259 10.6151
R1186 B.n535 B.n534 10.6151
R1187 B.n536 B.n535 10.6151
R1188 B.n536 B.n251 10.6151
R1189 B.n546 B.n251 10.6151
R1190 B.n547 B.n546 10.6151
R1191 B.n548 B.n547 10.6151
R1192 B.n548 B.n243 10.6151
R1193 B.n559 B.n243 10.6151
R1194 B.n560 B.n559 10.6151
R1195 B.n561 B.n560 10.6151
R1196 B.n561 B.n0 10.6151
R1197 B.n661 B.n1 10.6151
R1198 B.n661 B.n660 10.6151
R1199 B.n660 B.n659 10.6151
R1200 B.n659 B.n10 10.6151
R1201 B.n653 B.n10 10.6151
R1202 B.n653 B.n652 10.6151
R1203 B.n652 B.n651 10.6151
R1204 B.n651 B.n17 10.6151
R1205 B.n645 B.n17 10.6151
R1206 B.n645 B.n644 10.6151
R1207 B.n644 B.n643 10.6151
R1208 B.n643 B.n24 10.6151
R1209 B.n637 B.n24 10.6151
R1210 B.n637 B.n636 10.6151
R1211 B.n636 B.n635 10.6151
R1212 B.n635 B.n31 10.6151
R1213 B.n629 B.n31 10.6151
R1214 B.n629 B.n628 10.6151
R1215 B.n628 B.n627 10.6151
R1216 B.n627 B.n38 10.6151
R1217 B.n621 B.n38 10.6151
R1218 B.n621 B.n620 10.6151
R1219 B.n620 B.n619 10.6151
R1220 B.n619 B.n45 10.6151
R1221 B.n613 B.n45 10.6151
R1222 B.n613 B.n612 10.6151
R1223 B.n612 B.n611 10.6151
R1224 B.n611 B.n52 10.6151
R1225 B.n532 B.t4 10.427
R1226 B.n641 B.t5 10.427
R1227 B.n158 B.n157 9.36635
R1228 B.n180 B.n179 9.36635
R1229 B.n418 B.n335 9.36635
R1230 B.n395 B.n338 9.36635
R1231 B.n496 B.t9 7.21887
R1232 B.n617 B.t16 7.21887
R1233 B.n667 B.n0 2.81026
R1234 B.n667 B.n1 2.81026
R1235 B.n544 B.t0 2.40662
R1236 B.n649 B.t6 2.40662
R1237 B.n159 B.n158 1.24928
R1238 B.n179 B.n178 1.24928
R1239 B.n415 B.n335 1.24928
R1240 B.n398 B.n338 1.24928
R1241 VN.n3 VN.t6 241.387
R1242 VN.n16 VN.t3 241.387
R1243 VN.n11 VN.t2 218.637
R1244 VN.n24 VN.t7 218.637
R1245 VN.n4 VN.t1 183.248
R1246 VN.n1 VN.t0 183.248
R1247 VN.n17 VN.t4 183.248
R1248 VN.n14 VN.t5 183.248
R1249 VN.n23 VN.n13 161.3
R1250 VN.n22 VN.n21 161.3
R1251 VN.n20 VN.n19 161.3
R1252 VN.n18 VN.n15 161.3
R1253 VN.n10 VN.n0 161.3
R1254 VN.n9 VN.n8 161.3
R1255 VN.n7 VN.n6 161.3
R1256 VN.n5 VN.n2 161.3
R1257 VN.n25 VN.n24 80.6037
R1258 VN.n12 VN.n11 80.6037
R1259 VN.n6 VN.n5 56.5617
R1260 VN.n19 VN.n18 56.5617
R1261 VN.n11 VN.n10 49.4301
R1262 VN.n24 VN.n23 49.4301
R1263 VN VN.n25 41.6884
R1264 VN.n4 VN.n3 33.9241
R1265 VN.n17 VN.n16 33.9241
R1266 VN.n16 VN.n15 28.263
R1267 VN.n3 VN.n2 28.263
R1268 VN.n10 VN.n9 24.5923
R1269 VN.n23 VN.n22 24.5923
R1270 VN.n5 VN.n4 23.1168
R1271 VN.n6 VN.n1 23.1168
R1272 VN.n18 VN.n17 23.1168
R1273 VN.n19 VN.n14 23.1168
R1274 VN.n9 VN.n1 1.47601
R1275 VN.n22 VN.n14 1.47601
R1276 VN.n25 VN.n13 0.285035
R1277 VN.n12 VN.n0 0.285035
R1278 VN.n21 VN.n13 0.189894
R1279 VN.n21 VN.n20 0.189894
R1280 VN.n20 VN.n15 0.189894
R1281 VN.n7 VN.n2 0.189894
R1282 VN.n8 VN.n7 0.189894
R1283 VN.n8 VN.n0 0.189894
R1284 VN VN.n12 0.146778
R1285 VDD2.n2 VDD2.n1 63.2199
R1286 VDD2.n2 VDD2.n0 63.2199
R1287 VDD2 VDD2.n5 63.217
R1288 VDD2.n4 VDD2.n3 62.6545
R1289 VDD2.n4 VDD2.n2 36.5774
R1290 VDD2.n5 VDD2.t3 2.34647
R1291 VDD2.n5 VDD2.t4 2.34647
R1292 VDD2.n3 VDD2.t0 2.34647
R1293 VDD2.n3 VDD2.t2 2.34647
R1294 VDD2.n1 VDD2.t7 2.34647
R1295 VDD2.n1 VDD2.t5 2.34647
R1296 VDD2.n0 VDD2.t1 2.34647
R1297 VDD2.n0 VDD2.t6 2.34647
R1298 VDD2 VDD2.n4 0.679379
C0 VTAIL VDD2 7.28102f
C1 VN VDD2 4.89457f
C2 VTAIL VN 4.94818f
C3 VDD2 VP 0.361507f
C4 VTAIL VP 4.96229f
C5 VDD2 VDD1 1.03155f
C6 VN VP 5.17645f
C7 VTAIL VDD1 7.236589f
C8 VN VDD1 0.149422f
C9 VP VDD1 5.10601f
C10 VDD2 B 3.616516f
C11 VDD1 B 3.892128f
C12 VTAIL B 7.281541f
C13 VN B 9.62362f
C14 VP B 8.008044f
C15 VDD2.t1 B 0.17053f
C16 VDD2.t6 B 0.17053f
C17 VDD2.n0 B 1.47604f
C18 VDD2.t7 B 0.17053f
C19 VDD2.t5 B 0.17053f
C20 VDD2.n1 B 1.47604f
C21 VDD2.n2 B 2.25378f
C22 VDD2.t0 B 0.17053f
C23 VDD2.t2 B 0.17053f
C24 VDD2.n3 B 1.47269f
C25 VDD2.n4 B 2.20834f
C26 VDD2.t3 B 0.17053f
C27 VDD2.t4 B 0.17053f
C28 VDD2.n5 B 1.47601f
C29 VN.n0 B 0.049062f
C30 VN.t0 B 0.927202f
C31 VN.n1 B 0.355436f
C32 VN.n2 B 0.191786f
C33 VN.t1 B 0.927202f
C34 VN.t6 B 1.02963f
C35 VN.n3 B 0.404029f
C36 VN.n4 B 0.41312f
C37 VN.n5 B 0.051428f
C38 VN.n6 B 0.051428f
C39 VN.n7 B 0.036768f
C40 VN.n8 B 0.036768f
C41 VN.n9 B 0.036542f
C42 VN.n10 B 0.045141f
C43 VN.t2 B 0.989346f
C44 VN.n11 B 0.418516f
C45 VN.n12 B 0.034435f
C46 VN.n13 B 0.049062f
C47 VN.t5 B 0.927202f
C48 VN.n14 B 0.355436f
C49 VN.n15 B 0.191786f
C50 VN.t4 B 0.927202f
C51 VN.t3 B 1.02963f
C52 VN.n16 B 0.404029f
C53 VN.n17 B 0.41312f
C54 VN.n18 B 0.051428f
C55 VN.n19 B 0.051428f
C56 VN.n20 B 0.036768f
C57 VN.n21 B 0.036768f
C58 VN.n22 B 0.036542f
C59 VN.n23 B 0.045141f
C60 VN.t7 B 0.989346f
C61 VN.n24 B 0.418516f
C62 VN.n25 B 1.51542f
C63 VDD1.t1 B 0.170607f
C64 VDD1.t2 B 0.170607f
C65 VDD1.n0 B 1.47747f
C66 VDD1.t5 B 0.170607f
C67 VDD1.t7 B 0.170607f
C68 VDD1.n1 B 1.47671f
C69 VDD1.t6 B 0.170607f
C70 VDD1.t4 B 0.170607f
C71 VDD1.n2 B 1.47671f
C72 VDD1.n3 B 2.30922f
C73 VDD1.t0 B 0.170607f
C74 VDD1.t3 B 0.170607f
C75 VDD1.n4 B 1.47335f
C76 VDD1.n5 B 2.23981f
C77 VTAIL.t6 B 0.134626f
C78 VTAIL.t5 B 0.134626f
C79 VTAIL.n0 B 1.10244f
C80 VTAIL.n1 B 0.286999f
C81 VTAIL.t1 B 1.40479f
C82 VTAIL.n2 B 0.378589f
C83 VTAIL.t12 B 1.40479f
C84 VTAIL.n3 B 0.378589f
C85 VTAIL.t10 B 0.134626f
C86 VTAIL.t9 B 0.134626f
C87 VTAIL.n4 B 1.10244f
C88 VTAIL.n5 B 0.363955f
C89 VTAIL.t13 B 1.40479f
C90 VTAIL.n6 B 1.17619f
C91 VTAIL.t2 B 1.40479f
C92 VTAIL.n7 B 1.17619f
C93 VTAIL.t4 B 0.134626f
C94 VTAIL.t0 B 0.134626f
C95 VTAIL.n8 B 1.10244f
C96 VTAIL.n9 B 0.363953f
C97 VTAIL.t3 B 1.40479f
C98 VTAIL.n10 B 0.378583f
C99 VTAIL.t14 B 1.40479f
C100 VTAIL.n11 B 0.378583f
C101 VTAIL.t15 B 0.134626f
C102 VTAIL.t11 B 0.134626f
C103 VTAIL.n12 B 1.10244f
C104 VTAIL.n13 B 0.363953f
C105 VTAIL.t8 B 1.40479f
C106 VTAIL.n14 B 1.17619f
C107 VTAIL.t7 B 1.40479f
C108 VTAIL.n15 B 1.17241f
C109 VP.n0 B 0.050216f
C110 VP.t1 B 0.949016f
C111 VP.n1 B 0.363798f
C112 VP.n2 B 0.037633f
C113 VP.t0 B 0.949016f
C114 VP.n3 B 0.046203f
C115 VP.n4 B 0.050216f
C116 VP.t4 B 1.01262f
C117 VP.t7 B 0.949016f
C118 VP.n5 B 0.363798f
C119 VP.n6 B 0.196299f
C120 VP.t5 B 0.949016f
C121 VP.t6 B 1.05386f
C122 VP.n7 B 0.413534f
C123 VP.n8 B 0.42284f
C124 VP.n9 B 0.052638f
C125 VP.n10 B 0.052638f
C126 VP.n11 B 0.037633f
C127 VP.n12 B 0.037633f
C128 VP.n13 B 0.037402f
C129 VP.n14 B 0.046203f
C130 VP.n15 B 0.428362f
C131 VP.n16 B 1.52991f
C132 VP.t2 B 1.01262f
C133 VP.n17 B 0.428362f
C134 VP.n18 B 1.56268f
C135 VP.n19 B 0.050216f
C136 VP.n20 B 0.037633f
C137 VP.n21 B 0.037402f
C138 VP.n22 B 0.363798f
C139 VP.n23 B 0.052638f
C140 VP.n24 B 0.052638f
C141 VP.n25 B 0.037633f
C142 VP.n26 B 0.037633f
C143 VP.n27 B 0.037402f
C144 VP.n28 B 0.046203f
C145 VP.t3 B 1.01262f
C146 VP.n29 B 0.428362f
C147 VP.n30 B 0.035245f
.ends

