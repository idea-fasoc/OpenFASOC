* NGSPICE file created from diff_pair_sample_0535.ext - technology: sky130A

.subckt diff_pair_sample_0535 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=1.8369 pd=10.2 as=0 ps=0 w=4.71 l=0.26
X1 VDD2.t9 VN.t0 VTAIL.t17 B.t4 sky130_fd_pr__nfet_01v8 ad=1.8369 pd=10.2 as=0.77715 ps=5.04 w=4.71 l=0.26
X2 VTAIL.t13 VN.t1 VDD2.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=0.77715 ps=5.04 w=4.71 l=0.26
X3 VDD1.t9 VP.t0 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=1.8369 ps=10.2 w=4.71 l=0.26
X4 VDD2.t7 VN.t2 VTAIL.t18 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8369 pd=10.2 as=0.77715 ps=5.04 w=4.71 l=0.26
X5 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=1.8369 pd=10.2 as=0 ps=0 w=4.71 l=0.26
X6 VDD2.t6 VN.t3 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=0.77715 ps=5.04 w=4.71 l=0.26
X7 VDD1.t8 VP.t1 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8369 pd=10.2 as=0.77715 ps=5.04 w=4.71 l=0.26
X8 VTAIL.t0 VP.t2 VDD1.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=0.77715 ps=5.04 w=4.71 l=0.26
X9 VTAIL.t9 VN.t4 VDD2.t5 B.t9 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=0.77715 ps=5.04 w=4.71 l=0.26
X10 VTAIL.t14 VN.t5 VDD2.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=0.77715 ps=5.04 w=4.71 l=0.26
X11 VDD1.t6 VP.t3 VTAIL.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=0.77715 ps=5.04 w=4.71 l=0.26
X12 VDD1.t5 VP.t4 VTAIL.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=1.8369 pd=10.2 as=0.77715 ps=5.04 w=4.71 l=0.26
X13 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=1.8369 pd=10.2 as=0 ps=0 w=4.71 l=0.26
X14 VDD2.t3 VN.t6 VTAIL.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=1.8369 ps=10.2 w=4.71 l=0.26
X15 VDD1.t4 VP.t5 VTAIL.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=1.8369 ps=10.2 w=4.71 l=0.26
X16 VTAIL.t8 VP.t6 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=0.77715 ps=5.04 w=4.71 l=0.26
X17 VTAIL.t19 VP.t7 VDD1.t2 B.t9 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=0.77715 ps=5.04 w=4.71 l=0.26
X18 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.8369 pd=10.2 as=0 ps=0 w=4.71 l=0.26
X19 VDD2.t2 VN.t7 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=0.77715 ps=5.04 w=4.71 l=0.26
X20 VDD2.t1 VN.t8 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=1.8369 ps=10.2 w=4.71 l=0.26
X21 VTAIL.t12 VN.t9 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=0.77715 ps=5.04 w=4.71 l=0.26
X22 VDD1.t1 VP.t8 VTAIL.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=0.77715 ps=5.04 w=4.71 l=0.26
X23 VTAIL.t3 VP.t9 VDD1.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=0.77715 ps=5.04 w=4.71 l=0.26
R0 B.n68 B.t10 659.028
R1 B.n65 B.t21 659.028
R2 B.n220 B.t18 659.028
R3 B.n212 B.t14 659.028
R4 B.n409 B.n408 585
R5 B.n165 B.n64 585
R6 B.n164 B.n163 585
R7 B.n162 B.n161 585
R8 B.n160 B.n159 585
R9 B.n158 B.n157 585
R10 B.n156 B.n155 585
R11 B.n154 B.n153 585
R12 B.n152 B.n151 585
R13 B.n150 B.n149 585
R14 B.n148 B.n147 585
R15 B.n146 B.n145 585
R16 B.n144 B.n143 585
R17 B.n142 B.n141 585
R18 B.n140 B.n139 585
R19 B.n138 B.n137 585
R20 B.n136 B.n135 585
R21 B.n134 B.n133 585
R22 B.n132 B.n131 585
R23 B.n130 B.n129 585
R24 B.n128 B.n127 585
R25 B.n126 B.n125 585
R26 B.n124 B.n123 585
R27 B.n122 B.n121 585
R28 B.n120 B.n119 585
R29 B.n118 B.n117 585
R30 B.n116 B.n115 585
R31 B.n114 B.n113 585
R32 B.n112 B.n111 585
R33 B.n110 B.n109 585
R34 B.n108 B.n107 585
R35 B.n106 B.n105 585
R36 B.n104 B.n103 585
R37 B.n102 B.n101 585
R38 B.n100 B.n99 585
R39 B.n98 B.n97 585
R40 B.n96 B.n95 585
R41 B.n94 B.n93 585
R42 B.n92 B.n91 585
R43 B.n90 B.n89 585
R44 B.n88 B.n87 585
R45 B.n86 B.n85 585
R46 B.n84 B.n83 585
R47 B.n82 B.n81 585
R48 B.n80 B.n79 585
R49 B.n78 B.n77 585
R50 B.n76 B.n75 585
R51 B.n74 B.n73 585
R52 B.n72 B.n71 585
R53 B.n38 B.n37 585
R54 B.n407 B.n39 585
R55 B.n412 B.n39 585
R56 B.n406 B.n405 585
R57 B.n405 B.n35 585
R58 B.n404 B.n34 585
R59 B.n418 B.n34 585
R60 B.n403 B.n33 585
R61 B.n419 B.n33 585
R62 B.n402 B.n32 585
R63 B.n420 B.n32 585
R64 B.n401 B.n400 585
R65 B.n400 B.n28 585
R66 B.n399 B.n27 585
R67 B.n426 B.n27 585
R68 B.n398 B.n26 585
R69 B.n427 B.n26 585
R70 B.n397 B.n25 585
R71 B.n428 B.n25 585
R72 B.n396 B.n395 585
R73 B.n395 B.n24 585
R74 B.n394 B.n20 585
R75 B.n434 B.n20 585
R76 B.n393 B.n19 585
R77 B.n435 B.n19 585
R78 B.n392 B.n18 585
R79 B.n436 B.n18 585
R80 B.n391 B.n390 585
R81 B.n390 B.n13 585
R82 B.n389 B.n12 585
R83 B.n442 B.n12 585
R84 B.n388 B.n11 585
R85 B.n443 B.n11 585
R86 B.n387 B.n10 585
R87 B.n444 B.n10 585
R88 B.n386 B.n7 585
R89 B.n447 B.n7 585
R90 B.n385 B.n6 585
R91 B.n448 B.n6 585
R92 B.n384 B.n5 585
R93 B.n449 B.n5 585
R94 B.n383 B.n382 585
R95 B.n382 B.n4 585
R96 B.n381 B.n166 585
R97 B.n381 B.n380 585
R98 B.n371 B.n167 585
R99 B.n168 B.n167 585
R100 B.n373 B.n372 585
R101 B.n374 B.n373 585
R102 B.n370 B.n173 585
R103 B.n173 B.n172 585
R104 B.n369 B.n368 585
R105 B.n368 B.n367 585
R106 B.n175 B.n174 585
R107 B.n176 B.n175 585
R108 B.n360 B.n359 585
R109 B.n361 B.n360 585
R110 B.n358 B.n180 585
R111 B.n184 B.n180 585
R112 B.n357 B.n356 585
R113 B.n356 B.n355 585
R114 B.n182 B.n181 585
R115 B.n183 B.n182 585
R116 B.n348 B.n347 585
R117 B.n349 B.n348 585
R118 B.n346 B.n189 585
R119 B.n189 B.n188 585
R120 B.n345 B.n344 585
R121 B.n344 B.n343 585
R122 B.n191 B.n190 585
R123 B.n192 B.n191 585
R124 B.n336 B.n335 585
R125 B.n337 B.n336 585
R126 B.n334 B.n197 585
R127 B.n197 B.n196 585
R128 B.n333 B.n332 585
R129 B.n332 B.n331 585
R130 B.n328 B.n201 585
R131 B.n327 B.n326 585
R132 B.n324 B.n202 585
R133 B.n324 B.n200 585
R134 B.n323 B.n322 585
R135 B.n321 B.n320 585
R136 B.n319 B.n204 585
R137 B.n317 B.n316 585
R138 B.n315 B.n205 585
R139 B.n314 B.n313 585
R140 B.n311 B.n206 585
R141 B.n309 B.n308 585
R142 B.n307 B.n207 585
R143 B.n306 B.n305 585
R144 B.n303 B.n208 585
R145 B.n301 B.n300 585
R146 B.n299 B.n209 585
R147 B.n298 B.n297 585
R148 B.n295 B.n210 585
R149 B.n293 B.n292 585
R150 B.n291 B.n211 585
R151 B.n289 B.n288 585
R152 B.n286 B.n214 585
R153 B.n284 B.n283 585
R154 B.n282 B.n215 585
R155 B.n281 B.n280 585
R156 B.n278 B.n216 585
R157 B.n276 B.n275 585
R158 B.n274 B.n217 585
R159 B.n273 B.n272 585
R160 B.n270 B.n218 585
R161 B.n268 B.n267 585
R162 B.n266 B.n219 585
R163 B.n265 B.n264 585
R164 B.n262 B.n223 585
R165 B.n260 B.n259 585
R166 B.n258 B.n224 585
R167 B.n257 B.n256 585
R168 B.n254 B.n225 585
R169 B.n252 B.n251 585
R170 B.n250 B.n226 585
R171 B.n249 B.n248 585
R172 B.n246 B.n227 585
R173 B.n244 B.n243 585
R174 B.n242 B.n228 585
R175 B.n241 B.n240 585
R176 B.n238 B.n229 585
R177 B.n236 B.n235 585
R178 B.n234 B.n230 585
R179 B.n233 B.n232 585
R180 B.n199 B.n198 585
R181 B.n200 B.n199 585
R182 B.n330 B.n329 585
R183 B.n331 B.n330 585
R184 B.n195 B.n194 585
R185 B.n196 B.n195 585
R186 B.n339 B.n338 585
R187 B.n338 B.n337 585
R188 B.n340 B.n193 585
R189 B.n193 B.n192 585
R190 B.n342 B.n341 585
R191 B.n343 B.n342 585
R192 B.n187 B.n186 585
R193 B.n188 B.n187 585
R194 B.n351 B.n350 585
R195 B.n350 B.n349 585
R196 B.n352 B.n185 585
R197 B.n185 B.n183 585
R198 B.n354 B.n353 585
R199 B.n355 B.n354 585
R200 B.n179 B.n178 585
R201 B.n184 B.n179 585
R202 B.n363 B.n362 585
R203 B.n362 B.n361 585
R204 B.n364 B.n177 585
R205 B.n177 B.n176 585
R206 B.n366 B.n365 585
R207 B.n367 B.n366 585
R208 B.n171 B.n170 585
R209 B.n172 B.n171 585
R210 B.n376 B.n375 585
R211 B.n375 B.n374 585
R212 B.n377 B.n169 585
R213 B.n169 B.n168 585
R214 B.n379 B.n378 585
R215 B.n380 B.n379 585
R216 B.n3 B.n0 585
R217 B.n4 B.n3 585
R218 B.n446 B.n1 585
R219 B.n447 B.n446 585
R220 B.n445 B.n9 585
R221 B.n445 B.n444 585
R222 B.n15 B.n8 585
R223 B.n443 B.n8 585
R224 B.n441 B.n440 585
R225 B.n442 B.n441 585
R226 B.n439 B.n14 585
R227 B.n14 B.n13 585
R228 B.n438 B.n437 585
R229 B.n437 B.n436 585
R230 B.n17 B.n16 585
R231 B.n435 B.n17 585
R232 B.n433 B.n432 585
R233 B.n434 B.n433 585
R234 B.n431 B.n21 585
R235 B.n24 B.n21 585
R236 B.n430 B.n429 585
R237 B.n429 B.n428 585
R238 B.n23 B.n22 585
R239 B.n427 B.n23 585
R240 B.n425 B.n424 585
R241 B.n426 B.n425 585
R242 B.n423 B.n29 585
R243 B.n29 B.n28 585
R244 B.n422 B.n421 585
R245 B.n421 B.n420 585
R246 B.n31 B.n30 585
R247 B.n419 B.n31 585
R248 B.n417 B.n416 585
R249 B.n418 B.n417 585
R250 B.n415 B.n36 585
R251 B.n36 B.n35 585
R252 B.n414 B.n413 585
R253 B.n413 B.n412 585
R254 B.n450 B.n449 585
R255 B.n448 B.n2 585
R256 B.n413 B.n38 497.305
R257 B.n409 B.n39 497.305
R258 B.n332 B.n199 497.305
R259 B.n330 B.n201 497.305
R260 B.n411 B.n410 256.663
R261 B.n411 B.n63 256.663
R262 B.n411 B.n62 256.663
R263 B.n411 B.n61 256.663
R264 B.n411 B.n60 256.663
R265 B.n411 B.n59 256.663
R266 B.n411 B.n58 256.663
R267 B.n411 B.n57 256.663
R268 B.n411 B.n56 256.663
R269 B.n411 B.n55 256.663
R270 B.n411 B.n54 256.663
R271 B.n411 B.n53 256.663
R272 B.n411 B.n52 256.663
R273 B.n411 B.n51 256.663
R274 B.n411 B.n50 256.663
R275 B.n411 B.n49 256.663
R276 B.n411 B.n48 256.663
R277 B.n411 B.n47 256.663
R278 B.n411 B.n46 256.663
R279 B.n411 B.n45 256.663
R280 B.n411 B.n44 256.663
R281 B.n411 B.n43 256.663
R282 B.n411 B.n42 256.663
R283 B.n411 B.n41 256.663
R284 B.n411 B.n40 256.663
R285 B.n325 B.n200 256.663
R286 B.n203 B.n200 256.663
R287 B.n318 B.n200 256.663
R288 B.n312 B.n200 256.663
R289 B.n310 B.n200 256.663
R290 B.n304 B.n200 256.663
R291 B.n302 B.n200 256.663
R292 B.n296 B.n200 256.663
R293 B.n294 B.n200 256.663
R294 B.n287 B.n200 256.663
R295 B.n285 B.n200 256.663
R296 B.n279 B.n200 256.663
R297 B.n277 B.n200 256.663
R298 B.n271 B.n200 256.663
R299 B.n269 B.n200 256.663
R300 B.n263 B.n200 256.663
R301 B.n261 B.n200 256.663
R302 B.n255 B.n200 256.663
R303 B.n253 B.n200 256.663
R304 B.n247 B.n200 256.663
R305 B.n245 B.n200 256.663
R306 B.n239 B.n200 256.663
R307 B.n237 B.n200 256.663
R308 B.n231 B.n200 256.663
R309 B.n452 B.n451 256.663
R310 B.n65 B.t22 168.607
R311 B.n220 B.t20 168.607
R312 B.n68 B.t12 168.607
R313 B.n212 B.t17 168.607
R314 B.n73 B.n72 163.367
R315 B.n77 B.n76 163.367
R316 B.n81 B.n80 163.367
R317 B.n85 B.n84 163.367
R318 B.n89 B.n88 163.367
R319 B.n93 B.n92 163.367
R320 B.n97 B.n96 163.367
R321 B.n101 B.n100 163.367
R322 B.n105 B.n104 163.367
R323 B.n109 B.n108 163.367
R324 B.n113 B.n112 163.367
R325 B.n117 B.n116 163.367
R326 B.n121 B.n120 163.367
R327 B.n125 B.n124 163.367
R328 B.n129 B.n128 163.367
R329 B.n133 B.n132 163.367
R330 B.n137 B.n136 163.367
R331 B.n141 B.n140 163.367
R332 B.n145 B.n144 163.367
R333 B.n149 B.n148 163.367
R334 B.n153 B.n152 163.367
R335 B.n157 B.n156 163.367
R336 B.n161 B.n160 163.367
R337 B.n163 B.n64 163.367
R338 B.n332 B.n197 163.367
R339 B.n336 B.n197 163.367
R340 B.n336 B.n191 163.367
R341 B.n344 B.n191 163.367
R342 B.n344 B.n189 163.367
R343 B.n348 B.n189 163.367
R344 B.n348 B.n182 163.367
R345 B.n356 B.n182 163.367
R346 B.n356 B.n180 163.367
R347 B.n360 B.n180 163.367
R348 B.n360 B.n175 163.367
R349 B.n368 B.n175 163.367
R350 B.n368 B.n173 163.367
R351 B.n373 B.n173 163.367
R352 B.n373 B.n167 163.367
R353 B.n381 B.n167 163.367
R354 B.n382 B.n381 163.367
R355 B.n382 B.n5 163.367
R356 B.n6 B.n5 163.367
R357 B.n7 B.n6 163.367
R358 B.n10 B.n7 163.367
R359 B.n11 B.n10 163.367
R360 B.n12 B.n11 163.367
R361 B.n390 B.n12 163.367
R362 B.n390 B.n18 163.367
R363 B.n19 B.n18 163.367
R364 B.n20 B.n19 163.367
R365 B.n395 B.n20 163.367
R366 B.n395 B.n25 163.367
R367 B.n26 B.n25 163.367
R368 B.n27 B.n26 163.367
R369 B.n400 B.n27 163.367
R370 B.n400 B.n32 163.367
R371 B.n33 B.n32 163.367
R372 B.n34 B.n33 163.367
R373 B.n405 B.n34 163.367
R374 B.n405 B.n39 163.367
R375 B.n326 B.n324 163.367
R376 B.n324 B.n323 163.367
R377 B.n320 B.n319 163.367
R378 B.n317 B.n205 163.367
R379 B.n313 B.n311 163.367
R380 B.n309 B.n207 163.367
R381 B.n305 B.n303 163.367
R382 B.n301 B.n209 163.367
R383 B.n297 B.n295 163.367
R384 B.n293 B.n211 163.367
R385 B.n288 B.n286 163.367
R386 B.n284 B.n215 163.367
R387 B.n280 B.n278 163.367
R388 B.n276 B.n217 163.367
R389 B.n272 B.n270 163.367
R390 B.n268 B.n219 163.367
R391 B.n264 B.n262 163.367
R392 B.n260 B.n224 163.367
R393 B.n256 B.n254 163.367
R394 B.n252 B.n226 163.367
R395 B.n248 B.n246 163.367
R396 B.n244 B.n228 163.367
R397 B.n240 B.n238 163.367
R398 B.n236 B.n230 163.367
R399 B.n232 B.n199 163.367
R400 B.n330 B.n195 163.367
R401 B.n338 B.n195 163.367
R402 B.n338 B.n193 163.367
R403 B.n342 B.n193 163.367
R404 B.n342 B.n187 163.367
R405 B.n350 B.n187 163.367
R406 B.n350 B.n185 163.367
R407 B.n354 B.n185 163.367
R408 B.n354 B.n179 163.367
R409 B.n362 B.n179 163.367
R410 B.n362 B.n177 163.367
R411 B.n366 B.n177 163.367
R412 B.n366 B.n171 163.367
R413 B.n375 B.n171 163.367
R414 B.n375 B.n169 163.367
R415 B.n379 B.n169 163.367
R416 B.n379 B.n3 163.367
R417 B.n450 B.n3 163.367
R418 B.n446 B.n2 163.367
R419 B.n446 B.n445 163.367
R420 B.n445 B.n8 163.367
R421 B.n441 B.n8 163.367
R422 B.n441 B.n14 163.367
R423 B.n437 B.n14 163.367
R424 B.n437 B.n17 163.367
R425 B.n433 B.n17 163.367
R426 B.n433 B.n21 163.367
R427 B.n429 B.n21 163.367
R428 B.n429 B.n23 163.367
R429 B.n425 B.n23 163.367
R430 B.n425 B.n29 163.367
R431 B.n421 B.n29 163.367
R432 B.n421 B.n31 163.367
R433 B.n417 B.n31 163.367
R434 B.n417 B.n36 163.367
R435 B.n413 B.n36 163.367
R436 B.n66 B.t23 157.163
R437 B.n221 B.t19 157.163
R438 B.n69 B.t13 157.163
R439 B.n213 B.t16 157.163
R440 B.n331 B.n200 137.708
R441 B.n412 B.n411 137.708
R442 B.n331 B.n196 74.9129
R443 B.n337 B.n196 74.9129
R444 B.n337 B.n192 74.9129
R445 B.n343 B.n192 74.9129
R446 B.n349 B.n188 74.9129
R447 B.n349 B.n183 74.9129
R448 B.n355 B.n183 74.9129
R449 B.n355 B.n184 74.9129
R450 B.n367 B.n176 74.9129
R451 B.n374 B.n172 74.9129
R452 B.n380 B.n168 74.9129
R453 B.n449 B.n4 74.9129
R454 B.n449 B.n448 74.9129
R455 B.n448 B.n447 74.9129
R456 B.n444 B.n443 74.9129
R457 B.n442 B.n13 74.9129
R458 B.n436 B.n435 74.9129
R459 B.n428 B.n24 74.9129
R460 B.n428 B.n427 74.9129
R461 B.n427 B.n426 74.9129
R462 B.n426 B.n28 74.9129
R463 B.n420 B.n419 74.9129
R464 B.n419 B.n418 74.9129
R465 B.n418 B.n35 74.9129
R466 B.n412 B.n35 74.9129
R467 B.t8 B.n4 72.7096
R468 B.n447 B.t4 72.7096
R469 B.n40 B.n38 71.676
R470 B.n73 B.n41 71.676
R471 B.n77 B.n42 71.676
R472 B.n81 B.n43 71.676
R473 B.n85 B.n44 71.676
R474 B.n89 B.n45 71.676
R475 B.n93 B.n46 71.676
R476 B.n97 B.n47 71.676
R477 B.n101 B.n48 71.676
R478 B.n105 B.n49 71.676
R479 B.n109 B.n50 71.676
R480 B.n113 B.n51 71.676
R481 B.n117 B.n52 71.676
R482 B.n121 B.n53 71.676
R483 B.n125 B.n54 71.676
R484 B.n129 B.n55 71.676
R485 B.n133 B.n56 71.676
R486 B.n137 B.n57 71.676
R487 B.n141 B.n58 71.676
R488 B.n145 B.n59 71.676
R489 B.n149 B.n60 71.676
R490 B.n153 B.n61 71.676
R491 B.n157 B.n62 71.676
R492 B.n161 B.n63 71.676
R493 B.n410 B.n64 71.676
R494 B.n410 B.n409 71.676
R495 B.n163 B.n63 71.676
R496 B.n160 B.n62 71.676
R497 B.n156 B.n61 71.676
R498 B.n152 B.n60 71.676
R499 B.n148 B.n59 71.676
R500 B.n144 B.n58 71.676
R501 B.n140 B.n57 71.676
R502 B.n136 B.n56 71.676
R503 B.n132 B.n55 71.676
R504 B.n128 B.n54 71.676
R505 B.n124 B.n53 71.676
R506 B.n120 B.n52 71.676
R507 B.n116 B.n51 71.676
R508 B.n112 B.n50 71.676
R509 B.n108 B.n49 71.676
R510 B.n104 B.n48 71.676
R511 B.n100 B.n47 71.676
R512 B.n96 B.n46 71.676
R513 B.n92 B.n45 71.676
R514 B.n88 B.n44 71.676
R515 B.n84 B.n43 71.676
R516 B.n80 B.n42 71.676
R517 B.n76 B.n41 71.676
R518 B.n72 B.n40 71.676
R519 B.n325 B.n201 71.676
R520 B.n323 B.n203 71.676
R521 B.n319 B.n318 71.676
R522 B.n312 B.n205 71.676
R523 B.n311 B.n310 71.676
R524 B.n304 B.n207 71.676
R525 B.n303 B.n302 71.676
R526 B.n296 B.n209 71.676
R527 B.n295 B.n294 71.676
R528 B.n287 B.n211 71.676
R529 B.n286 B.n285 71.676
R530 B.n279 B.n215 71.676
R531 B.n278 B.n277 71.676
R532 B.n271 B.n217 71.676
R533 B.n270 B.n269 71.676
R534 B.n263 B.n219 71.676
R535 B.n262 B.n261 71.676
R536 B.n255 B.n224 71.676
R537 B.n254 B.n253 71.676
R538 B.n247 B.n226 71.676
R539 B.n246 B.n245 71.676
R540 B.n239 B.n228 71.676
R541 B.n238 B.n237 71.676
R542 B.n231 B.n230 71.676
R543 B.n326 B.n325 71.676
R544 B.n320 B.n203 71.676
R545 B.n318 B.n317 71.676
R546 B.n313 B.n312 71.676
R547 B.n310 B.n309 71.676
R548 B.n305 B.n304 71.676
R549 B.n302 B.n301 71.676
R550 B.n297 B.n296 71.676
R551 B.n294 B.n293 71.676
R552 B.n288 B.n287 71.676
R553 B.n285 B.n284 71.676
R554 B.n280 B.n279 71.676
R555 B.n277 B.n276 71.676
R556 B.n272 B.n271 71.676
R557 B.n269 B.n268 71.676
R558 B.n264 B.n263 71.676
R559 B.n261 B.n260 71.676
R560 B.n256 B.n255 71.676
R561 B.n253 B.n252 71.676
R562 B.n248 B.n247 71.676
R563 B.n245 B.n244 71.676
R564 B.n240 B.n239 71.676
R565 B.n237 B.n236 71.676
R566 B.n232 B.n231 71.676
R567 B.n451 B.n450 71.676
R568 B.n451 B.n2 71.676
R569 B.n361 B.t5 68.303
R570 B.n434 B.t0 68.303
R571 B.t15 B.n188 63.8963
R572 B.t11 B.n28 63.8963
R573 B.n361 B.t6 61.693
R574 B.t1 B.n434 61.693
R575 B.n70 B.n69 59.5399
R576 B.n67 B.n66 59.5399
R577 B.n222 B.n221 59.5399
R578 B.n290 B.n213 59.5399
R579 B.t9 B.n168 52.8798
R580 B.n443 B.t3 52.8798
R581 B.n367 B.t7 41.8633
R582 B.n436 B.t2 41.8633
R583 B.t7 B.n172 33.0501
R584 B.t2 B.n13 33.0501
R585 B.n329 B.n328 32.3127
R586 B.n333 B.n198 32.3127
R587 B.n408 B.n407 32.3127
R588 B.n414 B.n37 32.3127
R589 B.n374 B.t9 22.0335
R590 B.t3 B.n442 22.0335
R591 B B.n452 18.0485
R592 B.t6 B.n176 13.2203
R593 B.n435 B.t1 13.2203
R594 B.n69 B.n68 11.4429
R595 B.n66 B.n65 11.4429
R596 B.n221 B.n220 11.4429
R597 B.n213 B.n212 11.4429
R598 B.n343 B.t15 11.017
R599 B.n420 B.t11 11.017
R600 B.n329 B.n194 10.6151
R601 B.n339 B.n194 10.6151
R602 B.n340 B.n339 10.6151
R603 B.n341 B.n340 10.6151
R604 B.n341 B.n186 10.6151
R605 B.n351 B.n186 10.6151
R606 B.n352 B.n351 10.6151
R607 B.n353 B.n352 10.6151
R608 B.n353 B.n178 10.6151
R609 B.n363 B.n178 10.6151
R610 B.n364 B.n363 10.6151
R611 B.n365 B.n364 10.6151
R612 B.n365 B.n170 10.6151
R613 B.n376 B.n170 10.6151
R614 B.n377 B.n376 10.6151
R615 B.n378 B.n377 10.6151
R616 B.n378 B.n0 10.6151
R617 B.n328 B.n327 10.6151
R618 B.n327 B.n202 10.6151
R619 B.n322 B.n202 10.6151
R620 B.n322 B.n321 10.6151
R621 B.n321 B.n204 10.6151
R622 B.n316 B.n204 10.6151
R623 B.n316 B.n315 10.6151
R624 B.n315 B.n314 10.6151
R625 B.n314 B.n206 10.6151
R626 B.n308 B.n206 10.6151
R627 B.n308 B.n307 10.6151
R628 B.n307 B.n306 10.6151
R629 B.n306 B.n208 10.6151
R630 B.n300 B.n208 10.6151
R631 B.n300 B.n299 10.6151
R632 B.n299 B.n298 10.6151
R633 B.n298 B.n210 10.6151
R634 B.n292 B.n210 10.6151
R635 B.n292 B.n291 10.6151
R636 B.n289 B.n214 10.6151
R637 B.n283 B.n214 10.6151
R638 B.n283 B.n282 10.6151
R639 B.n282 B.n281 10.6151
R640 B.n281 B.n216 10.6151
R641 B.n275 B.n216 10.6151
R642 B.n275 B.n274 10.6151
R643 B.n274 B.n273 10.6151
R644 B.n273 B.n218 10.6151
R645 B.n267 B.n266 10.6151
R646 B.n266 B.n265 10.6151
R647 B.n265 B.n223 10.6151
R648 B.n259 B.n223 10.6151
R649 B.n259 B.n258 10.6151
R650 B.n258 B.n257 10.6151
R651 B.n257 B.n225 10.6151
R652 B.n251 B.n225 10.6151
R653 B.n251 B.n250 10.6151
R654 B.n250 B.n249 10.6151
R655 B.n249 B.n227 10.6151
R656 B.n243 B.n227 10.6151
R657 B.n243 B.n242 10.6151
R658 B.n242 B.n241 10.6151
R659 B.n241 B.n229 10.6151
R660 B.n235 B.n229 10.6151
R661 B.n235 B.n234 10.6151
R662 B.n234 B.n233 10.6151
R663 B.n233 B.n198 10.6151
R664 B.n334 B.n333 10.6151
R665 B.n335 B.n334 10.6151
R666 B.n335 B.n190 10.6151
R667 B.n345 B.n190 10.6151
R668 B.n346 B.n345 10.6151
R669 B.n347 B.n346 10.6151
R670 B.n347 B.n181 10.6151
R671 B.n357 B.n181 10.6151
R672 B.n358 B.n357 10.6151
R673 B.n359 B.n358 10.6151
R674 B.n359 B.n174 10.6151
R675 B.n369 B.n174 10.6151
R676 B.n370 B.n369 10.6151
R677 B.n372 B.n370 10.6151
R678 B.n372 B.n371 10.6151
R679 B.n371 B.n166 10.6151
R680 B.n383 B.n166 10.6151
R681 B.n384 B.n383 10.6151
R682 B.n385 B.n384 10.6151
R683 B.n386 B.n385 10.6151
R684 B.n387 B.n386 10.6151
R685 B.n388 B.n387 10.6151
R686 B.n389 B.n388 10.6151
R687 B.n391 B.n389 10.6151
R688 B.n392 B.n391 10.6151
R689 B.n393 B.n392 10.6151
R690 B.n394 B.n393 10.6151
R691 B.n396 B.n394 10.6151
R692 B.n397 B.n396 10.6151
R693 B.n398 B.n397 10.6151
R694 B.n399 B.n398 10.6151
R695 B.n401 B.n399 10.6151
R696 B.n402 B.n401 10.6151
R697 B.n403 B.n402 10.6151
R698 B.n404 B.n403 10.6151
R699 B.n406 B.n404 10.6151
R700 B.n407 B.n406 10.6151
R701 B.n9 B.n1 10.6151
R702 B.n15 B.n9 10.6151
R703 B.n440 B.n15 10.6151
R704 B.n440 B.n439 10.6151
R705 B.n439 B.n438 10.6151
R706 B.n438 B.n16 10.6151
R707 B.n432 B.n16 10.6151
R708 B.n432 B.n431 10.6151
R709 B.n431 B.n430 10.6151
R710 B.n430 B.n22 10.6151
R711 B.n424 B.n22 10.6151
R712 B.n424 B.n423 10.6151
R713 B.n423 B.n422 10.6151
R714 B.n422 B.n30 10.6151
R715 B.n416 B.n30 10.6151
R716 B.n416 B.n415 10.6151
R717 B.n415 B.n414 10.6151
R718 B.n71 B.n37 10.6151
R719 B.n74 B.n71 10.6151
R720 B.n75 B.n74 10.6151
R721 B.n78 B.n75 10.6151
R722 B.n79 B.n78 10.6151
R723 B.n82 B.n79 10.6151
R724 B.n83 B.n82 10.6151
R725 B.n86 B.n83 10.6151
R726 B.n87 B.n86 10.6151
R727 B.n90 B.n87 10.6151
R728 B.n91 B.n90 10.6151
R729 B.n94 B.n91 10.6151
R730 B.n95 B.n94 10.6151
R731 B.n98 B.n95 10.6151
R732 B.n99 B.n98 10.6151
R733 B.n102 B.n99 10.6151
R734 B.n103 B.n102 10.6151
R735 B.n106 B.n103 10.6151
R736 B.n107 B.n106 10.6151
R737 B.n111 B.n110 10.6151
R738 B.n114 B.n111 10.6151
R739 B.n115 B.n114 10.6151
R740 B.n118 B.n115 10.6151
R741 B.n119 B.n118 10.6151
R742 B.n122 B.n119 10.6151
R743 B.n123 B.n122 10.6151
R744 B.n126 B.n123 10.6151
R745 B.n127 B.n126 10.6151
R746 B.n131 B.n130 10.6151
R747 B.n134 B.n131 10.6151
R748 B.n135 B.n134 10.6151
R749 B.n138 B.n135 10.6151
R750 B.n139 B.n138 10.6151
R751 B.n142 B.n139 10.6151
R752 B.n143 B.n142 10.6151
R753 B.n146 B.n143 10.6151
R754 B.n147 B.n146 10.6151
R755 B.n150 B.n147 10.6151
R756 B.n151 B.n150 10.6151
R757 B.n154 B.n151 10.6151
R758 B.n155 B.n154 10.6151
R759 B.n158 B.n155 10.6151
R760 B.n159 B.n158 10.6151
R761 B.n162 B.n159 10.6151
R762 B.n164 B.n162 10.6151
R763 B.n165 B.n164 10.6151
R764 B.n408 B.n165 10.6151
R765 B.n291 B.n290 9.36635
R766 B.n267 B.n222 9.36635
R767 B.n107 B.n70 9.36635
R768 B.n130 B.n67 9.36635
R769 B.n452 B.n0 8.11757
R770 B.n452 B.n1 8.11757
R771 B.n184 B.t5 6.61042
R772 B.n24 B.t0 6.61042
R773 B.n380 B.t8 2.20381
R774 B.n444 B.t4 2.20381
R775 B.n290 B.n289 1.24928
R776 B.n222 B.n218 1.24928
R777 B.n110 B.n70 1.24928
R778 B.n127 B.n67 1.24928
R779 VN.n9 VN.t8 584.299
R780 VN.n3 VN.t0 584.299
R781 VN.n20 VN.t2 584.299
R782 VN.n14 VN.t6 584.299
R783 VN.n6 VN.t7 558.009
R784 VN.n8 VN.t9 558.009
R785 VN.n2 VN.t5 558.009
R786 VN.n17 VN.t3 558.009
R787 VN.n19 VN.t1 558.009
R788 VN.n13 VN.t4 558.009
R789 VN.n15 VN.n14 161.489
R790 VN.n4 VN.n3 161.489
R791 VN.n10 VN.n9 161.3
R792 VN.n21 VN.n20 161.3
R793 VN.n18 VN.n11 161.3
R794 VN.n17 VN.n16 161.3
R795 VN.n15 VN.n12 161.3
R796 VN.n7 VN.n0 161.3
R797 VN.n6 VN.n5 161.3
R798 VN.n4 VN.n1 161.3
R799 VN.n6 VN.n1 73.0308
R800 VN.n7 VN.n6 73.0308
R801 VN.n18 VN.n17 73.0308
R802 VN.n17 VN.n12 73.0308
R803 VN.n3 VN.n2 59.8853
R804 VN.n9 VN.n8 59.8853
R805 VN.n20 VN.n19 59.8853
R806 VN.n14 VN.n13 59.8853
R807 VN VN.n21 35.2335
R808 VN.n2 VN.n1 13.146
R809 VN.n8 VN.n7 13.146
R810 VN.n19 VN.n18 13.146
R811 VN.n13 VN.n12 13.146
R812 VN.n21 VN.n11 0.189894
R813 VN.n16 VN.n11 0.189894
R814 VN.n16 VN.n15 0.189894
R815 VN.n5 VN.n4 0.189894
R816 VN.n5 VN.n0 0.189894
R817 VN.n10 VN.n0 0.189894
R818 VN VN.n10 0.0516364
R819 VTAIL.n104 VTAIL.n86 289.615
R820 VTAIL.n20 VTAIL.n2 289.615
R821 VTAIL.n80 VTAIL.n62 289.615
R822 VTAIL.n52 VTAIL.n34 289.615
R823 VTAIL.n95 VTAIL.n94 185
R824 VTAIL.n97 VTAIL.n96 185
R825 VTAIL.n90 VTAIL.n89 185
R826 VTAIL.n103 VTAIL.n102 185
R827 VTAIL.n105 VTAIL.n104 185
R828 VTAIL.n11 VTAIL.n10 185
R829 VTAIL.n13 VTAIL.n12 185
R830 VTAIL.n6 VTAIL.n5 185
R831 VTAIL.n19 VTAIL.n18 185
R832 VTAIL.n21 VTAIL.n20 185
R833 VTAIL.n81 VTAIL.n80 185
R834 VTAIL.n79 VTAIL.n78 185
R835 VTAIL.n66 VTAIL.n65 185
R836 VTAIL.n73 VTAIL.n72 185
R837 VTAIL.n71 VTAIL.n70 185
R838 VTAIL.n53 VTAIL.n52 185
R839 VTAIL.n51 VTAIL.n50 185
R840 VTAIL.n38 VTAIL.n37 185
R841 VTAIL.n45 VTAIL.n44 185
R842 VTAIL.n43 VTAIL.n42 185
R843 VTAIL.n93 VTAIL.t10 147.714
R844 VTAIL.n9 VTAIL.t5 147.714
R845 VTAIL.n69 VTAIL.t6 147.714
R846 VTAIL.n41 VTAIL.t16 147.714
R847 VTAIL.n96 VTAIL.n95 104.615
R848 VTAIL.n96 VTAIL.n89 104.615
R849 VTAIL.n103 VTAIL.n89 104.615
R850 VTAIL.n104 VTAIL.n103 104.615
R851 VTAIL.n12 VTAIL.n11 104.615
R852 VTAIL.n12 VTAIL.n5 104.615
R853 VTAIL.n19 VTAIL.n5 104.615
R854 VTAIL.n20 VTAIL.n19 104.615
R855 VTAIL.n80 VTAIL.n79 104.615
R856 VTAIL.n79 VTAIL.n65 104.615
R857 VTAIL.n72 VTAIL.n65 104.615
R858 VTAIL.n72 VTAIL.n71 104.615
R859 VTAIL.n52 VTAIL.n51 104.615
R860 VTAIL.n51 VTAIL.n37 104.615
R861 VTAIL.n44 VTAIL.n37 104.615
R862 VTAIL.n44 VTAIL.n43 104.615
R863 VTAIL.n61 VTAIL.n60 56.8721
R864 VTAIL.n59 VTAIL.n58 56.8721
R865 VTAIL.n33 VTAIL.n32 56.8721
R866 VTAIL.n31 VTAIL.n30 56.8721
R867 VTAIL.n111 VTAIL.n110 56.8719
R868 VTAIL.n1 VTAIL.n0 56.8719
R869 VTAIL.n27 VTAIL.n26 56.8719
R870 VTAIL.n29 VTAIL.n28 56.8719
R871 VTAIL.n95 VTAIL.t10 52.3082
R872 VTAIL.n11 VTAIL.t5 52.3082
R873 VTAIL.n71 VTAIL.t6 52.3082
R874 VTAIL.n43 VTAIL.t16 52.3082
R875 VTAIL.n109 VTAIL.n108 35.0944
R876 VTAIL.n25 VTAIL.n24 35.0944
R877 VTAIL.n85 VTAIL.n84 35.0944
R878 VTAIL.n57 VTAIL.n56 35.0944
R879 VTAIL.n31 VTAIL.n29 17.4445
R880 VTAIL.n109 VTAIL.n85 16.9358
R881 VTAIL.n94 VTAIL.n93 15.6631
R882 VTAIL.n10 VTAIL.n9 15.6631
R883 VTAIL.n70 VTAIL.n69 15.6631
R884 VTAIL.n42 VTAIL.n41 15.6631
R885 VTAIL.n97 VTAIL.n92 12.8005
R886 VTAIL.n13 VTAIL.n8 12.8005
R887 VTAIL.n73 VTAIL.n68 12.8005
R888 VTAIL.n45 VTAIL.n40 12.8005
R889 VTAIL.n98 VTAIL.n90 12.0247
R890 VTAIL.n14 VTAIL.n6 12.0247
R891 VTAIL.n74 VTAIL.n66 12.0247
R892 VTAIL.n46 VTAIL.n38 12.0247
R893 VTAIL.n102 VTAIL.n101 11.249
R894 VTAIL.n18 VTAIL.n17 11.249
R895 VTAIL.n78 VTAIL.n77 11.249
R896 VTAIL.n50 VTAIL.n49 11.249
R897 VTAIL.n105 VTAIL.n88 10.4732
R898 VTAIL.n21 VTAIL.n4 10.4732
R899 VTAIL.n81 VTAIL.n64 10.4732
R900 VTAIL.n53 VTAIL.n36 10.4732
R901 VTAIL.n106 VTAIL.n86 9.69747
R902 VTAIL.n22 VTAIL.n2 9.69747
R903 VTAIL.n82 VTAIL.n62 9.69747
R904 VTAIL.n54 VTAIL.n34 9.69747
R905 VTAIL.n108 VTAIL.n107 9.45567
R906 VTAIL.n24 VTAIL.n23 9.45567
R907 VTAIL.n84 VTAIL.n83 9.45567
R908 VTAIL.n56 VTAIL.n55 9.45567
R909 VTAIL.n107 VTAIL.n106 9.3005
R910 VTAIL.n88 VTAIL.n87 9.3005
R911 VTAIL.n101 VTAIL.n100 9.3005
R912 VTAIL.n99 VTAIL.n98 9.3005
R913 VTAIL.n92 VTAIL.n91 9.3005
R914 VTAIL.n23 VTAIL.n22 9.3005
R915 VTAIL.n4 VTAIL.n3 9.3005
R916 VTAIL.n17 VTAIL.n16 9.3005
R917 VTAIL.n15 VTAIL.n14 9.3005
R918 VTAIL.n8 VTAIL.n7 9.3005
R919 VTAIL.n83 VTAIL.n82 9.3005
R920 VTAIL.n64 VTAIL.n63 9.3005
R921 VTAIL.n77 VTAIL.n76 9.3005
R922 VTAIL.n75 VTAIL.n74 9.3005
R923 VTAIL.n68 VTAIL.n67 9.3005
R924 VTAIL.n55 VTAIL.n54 9.3005
R925 VTAIL.n36 VTAIL.n35 9.3005
R926 VTAIL.n49 VTAIL.n48 9.3005
R927 VTAIL.n47 VTAIL.n46 9.3005
R928 VTAIL.n40 VTAIL.n39 9.3005
R929 VTAIL.n93 VTAIL.n91 4.39059
R930 VTAIL.n9 VTAIL.n7 4.39059
R931 VTAIL.n69 VTAIL.n67 4.39059
R932 VTAIL.n41 VTAIL.n39 4.39059
R933 VTAIL.n108 VTAIL.n86 4.26717
R934 VTAIL.n24 VTAIL.n2 4.26717
R935 VTAIL.n84 VTAIL.n62 4.26717
R936 VTAIL.n56 VTAIL.n34 4.26717
R937 VTAIL.n110 VTAIL.t11 4.20432
R938 VTAIL.n110 VTAIL.t12 4.20432
R939 VTAIL.n0 VTAIL.t17 4.20432
R940 VTAIL.n0 VTAIL.t14 4.20432
R941 VTAIL.n26 VTAIL.t4 4.20432
R942 VTAIL.n26 VTAIL.t19 4.20432
R943 VTAIL.n28 VTAIL.t7 4.20432
R944 VTAIL.n28 VTAIL.t3 4.20432
R945 VTAIL.n60 VTAIL.t1 4.20432
R946 VTAIL.n60 VTAIL.t0 4.20432
R947 VTAIL.n58 VTAIL.t2 4.20432
R948 VTAIL.n58 VTAIL.t8 4.20432
R949 VTAIL.n32 VTAIL.t15 4.20432
R950 VTAIL.n32 VTAIL.t9 4.20432
R951 VTAIL.n30 VTAIL.t18 4.20432
R952 VTAIL.n30 VTAIL.t13 4.20432
R953 VTAIL.n106 VTAIL.n105 3.49141
R954 VTAIL.n22 VTAIL.n21 3.49141
R955 VTAIL.n82 VTAIL.n81 3.49141
R956 VTAIL.n54 VTAIL.n53 3.49141
R957 VTAIL.n102 VTAIL.n88 2.71565
R958 VTAIL.n18 VTAIL.n4 2.71565
R959 VTAIL.n78 VTAIL.n64 2.71565
R960 VTAIL.n50 VTAIL.n36 2.71565
R961 VTAIL.n101 VTAIL.n90 1.93989
R962 VTAIL.n17 VTAIL.n6 1.93989
R963 VTAIL.n77 VTAIL.n66 1.93989
R964 VTAIL.n49 VTAIL.n38 1.93989
R965 VTAIL.n98 VTAIL.n97 1.16414
R966 VTAIL.n14 VTAIL.n13 1.16414
R967 VTAIL.n74 VTAIL.n73 1.16414
R968 VTAIL.n46 VTAIL.n45 1.16414
R969 VTAIL.n59 VTAIL.n57 0.724638
R970 VTAIL.n25 VTAIL.n1 0.724638
R971 VTAIL.n33 VTAIL.n31 0.509121
R972 VTAIL.n57 VTAIL.n33 0.509121
R973 VTAIL.n61 VTAIL.n59 0.509121
R974 VTAIL.n85 VTAIL.n61 0.509121
R975 VTAIL.n29 VTAIL.n27 0.509121
R976 VTAIL.n27 VTAIL.n25 0.509121
R977 VTAIL.n111 VTAIL.n109 0.509121
R978 VTAIL VTAIL.n1 0.440155
R979 VTAIL.n94 VTAIL.n92 0.388379
R980 VTAIL.n10 VTAIL.n8 0.388379
R981 VTAIL.n70 VTAIL.n68 0.388379
R982 VTAIL.n42 VTAIL.n40 0.388379
R983 VTAIL.n99 VTAIL.n91 0.155672
R984 VTAIL.n100 VTAIL.n99 0.155672
R985 VTAIL.n100 VTAIL.n87 0.155672
R986 VTAIL.n107 VTAIL.n87 0.155672
R987 VTAIL.n15 VTAIL.n7 0.155672
R988 VTAIL.n16 VTAIL.n15 0.155672
R989 VTAIL.n16 VTAIL.n3 0.155672
R990 VTAIL.n23 VTAIL.n3 0.155672
R991 VTAIL.n83 VTAIL.n63 0.155672
R992 VTAIL.n76 VTAIL.n63 0.155672
R993 VTAIL.n76 VTAIL.n75 0.155672
R994 VTAIL.n75 VTAIL.n67 0.155672
R995 VTAIL.n55 VTAIL.n35 0.155672
R996 VTAIL.n48 VTAIL.n35 0.155672
R997 VTAIL.n48 VTAIL.n47 0.155672
R998 VTAIL.n47 VTAIL.n39 0.155672
R999 VTAIL VTAIL.n111 0.0694655
R1000 VDD2.n45 VDD2.n27 289.615
R1001 VDD2.n18 VDD2.n0 289.615
R1002 VDD2.n46 VDD2.n45 185
R1003 VDD2.n44 VDD2.n43 185
R1004 VDD2.n31 VDD2.n30 185
R1005 VDD2.n38 VDD2.n37 185
R1006 VDD2.n36 VDD2.n35 185
R1007 VDD2.n9 VDD2.n8 185
R1008 VDD2.n11 VDD2.n10 185
R1009 VDD2.n4 VDD2.n3 185
R1010 VDD2.n17 VDD2.n16 185
R1011 VDD2.n19 VDD2.n18 185
R1012 VDD2.n34 VDD2.t7 147.714
R1013 VDD2.n7 VDD2.t9 147.714
R1014 VDD2.n45 VDD2.n44 104.615
R1015 VDD2.n44 VDD2.n30 104.615
R1016 VDD2.n37 VDD2.n30 104.615
R1017 VDD2.n37 VDD2.n36 104.615
R1018 VDD2.n10 VDD2.n9 104.615
R1019 VDD2.n10 VDD2.n3 104.615
R1020 VDD2.n17 VDD2.n3 104.615
R1021 VDD2.n18 VDD2.n17 104.615
R1022 VDD2.n26 VDD2.n25 73.8769
R1023 VDD2 VDD2.n53 73.874
R1024 VDD2.n52 VDD2.n51 73.5509
R1025 VDD2.n24 VDD2.n23 73.5507
R1026 VDD2.n36 VDD2.t7 52.3082
R1027 VDD2.n9 VDD2.t9 52.3082
R1028 VDD2.n24 VDD2.n22 52.2818
R1029 VDD2.n50 VDD2.n49 51.7732
R1030 VDD2.n50 VDD2.n26 30.1916
R1031 VDD2.n35 VDD2.n34 15.6631
R1032 VDD2.n8 VDD2.n7 15.6631
R1033 VDD2.n38 VDD2.n33 12.8005
R1034 VDD2.n11 VDD2.n6 12.8005
R1035 VDD2.n39 VDD2.n31 12.0247
R1036 VDD2.n12 VDD2.n4 12.0247
R1037 VDD2.n43 VDD2.n42 11.249
R1038 VDD2.n16 VDD2.n15 11.249
R1039 VDD2.n46 VDD2.n29 10.4732
R1040 VDD2.n19 VDD2.n2 10.4732
R1041 VDD2.n47 VDD2.n27 9.69747
R1042 VDD2.n20 VDD2.n0 9.69747
R1043 VDD2.n49 VDD2.n48 9.45567
R1044 VDD2.n22 VDD2.n21 9.45567
R1045 VDD2.n48 VDD2.n47 9.3005
R1046 VDD2.n29 VDD2.n28 9.3005
R1047 VDD2.n42 VDD2.n41 9.3005
R1048 VDD2.n40 VDD2.n39 9.3005
R1049 VDD2.n33 VDD2.n32 9.3005
R1050 VDD2.n21 VDD2.n20 9.3005
R1051 VDD2.n2 VDD2.n1 9.3005
R1052 VDD2.n15 VDD2.n14 9.3005
R1053 VDD2.n13 VDD2.n12 9.3005
R1054 VDD2.n6 VDD2.n5 9.3005
R1055 VDD2.n34 VDD2.n32 4.39059
R1056 VDD2.n7 VDD2.n5 4.39059
R1057 VDD2.n49 VDD2.n27 4.26717
R1058 VDD2.n22 VDD2.n0 4.26717
R1059 VDD2.n53 VDD2.t5 4.20432
R1060 VDD2.n53 VDD2.t3 4.20432
R1061 VDD2.n51 VDD2.t8 4.20432
R1062 VDD2.n51 VDD2.t6 4.20432
R1063 VDD2.n25 VDD2.t0 4.20432
R1064 VDD2.n25 VDD2.t1 4.20432
R1065 VDD2.n23 VDD2.t4 4.20432
R1066 VDD2.n23 VDD2.t2 4.20432
R1067 VDD2.n47 VDD2.n46 3.49141
R1068 VDD2.n20 VDD2.n19 3.49141
R1069 VDD2.n43 VDD2.n29 2.71565
R1070 VDD2.n16 VDD2.n2 2.71565
R1071 VDD2.n42 VDD2.n31 1.93989
R1072 VDD2.n15 VDD2.n4 1.93989
R1073 VDD2.n39 VDD2.n38 1.16414
R1074 VDD2.n12 VDD2.n11 1.16414
R1075 VDD2.n52 VDD2.n50 0.509121
R1076 VDD2.n35 VDD2.n33 0.388379
R1077 VDD2.n8 VDD2.n6 0.388379
R1078 VDD2 VDD2.n52 0.185845
R1079 VDD2.n48 VDD2.n28 0.155672
R1080 VDD2.n41 VDD2.n28 0.155672
R1081 VDD2.n41 VDD2.n40 0.155672
R1082 VDD2.n40 VDD2.n32 0.155672
R1083 VDD2.n13 VDD2.n5 0.155672
R1084 VDD2.n14 VDD2.n13 0.155672
R1085 VDD2.n14 VDD2.n1 0.155672
R1086 VDD2.n21 VDD2.n1 0.155672
R1087 VDD2.n26 VDD2.n24 0.0723091
R1088 VP.n21 VP.t5 584.299
R1089 VP.n14 VP.t1 584.299
R1090 VP.n5 VP.t4 584.299
R1091 VP.n11 VP.t0 584.299
R1092 VP.n18 VP.t8 558.009
R1093 VP.n20 VP.t7 558.009
R1094 VP.n13 VP.t9 558.009
R1095 VP.n8 VP.t3 558.009
R1096 VP.n4 VP.t6 558.009
R1097 VP.n10 VP.t2 558.009
R1098 VP.n6 VP.n5 161.489
R1099 VP.n22 VP.n21 161.3
R1100 VP.n6 VP.n3 161.3
R1101 VP.n8 VP.n7 161.3
R1102 VP.n9 VP.n2 161.3
R1103 VP.n12 VP.n11 161.3
R1104 VP.n19 VP.n0 161.3
R1105 VP.n18 VP.n17 161.3
R1106 VP.n16 VP.n1 161.3
R1107 VP.n15 VP.n14 161.3
R1108 VP.n18 VP.n1 73.0308
R1109 VP.n19 VP.n18 73.0308
R1110 VP.n8 VP.n3 73.0308
R1111 VP.n9 VP.n8 73.0308
R1112 VP.n14 VP.n13 59.8853
R1113 VP.n21 VP.n20 59.8853
R1114 VP.n5 VP.n4 59.8853
R1115 VP.n11 VP.n10 59.8853
R1116 VP.n15 VP.n12 34.8528
R1117 VP.n13 VP.n1 13.146
R1118 VP.n20 VP.n19 13.146
R1119 VP.n4 VP.n3 13.146
R1120 VP.n10 VP.n9 13.146
R1121 VP.n7 VP.n6 0.189894
R1122 VP.n7 VP.n2 0.189894
R1123 VP.n12 VP.n2 0.189894
R1124 VP.n16 VP.n15 0.189894
R1125 VP.n17 VP.n16 0.189894
R1126 VP.n17 VP.n0 0.189894
R1127 VP.n22 VP.n0 0.189894
R1128 VP VP.n22 0.0516364
R1129 VDD1.n18 VDD1.n0 289.615
R1130 VDD1.n43 VDD1.n25 289.615
R1131 VDD1.n19 VDD1.n18 185
R1132 VDD1.n17 VDD1.n16 185
R1133 VDD1.n4 VDD1.n3 185
R1134 VDD1.n11 VDD1.n10 185
R1135 VDD1.n9 VDD1.n8 185
R1136 VDD1.n34 VDD1.n33 185
R1137 VDD1.n36 VDD1.n35 185
R1138 VDD1.n29 VDD1.n28 185
R1139 VDD1.n42 VDD1.n41 185
R1140 VDD1.n44 VDD1.n43 185
R1141 VDD1.n7 VDD1.t5 147.714
R1142 VDD1.n32 VDD1.t8 147.714
R1143 VDD1.n18 VDD1.n17 104.615
R1144 VDD1.n17 VDD1.n3 104.615
R1145 VDD1.n10 VDD1.n3 104.615
R1146 VDD1.n10 VDD1.n9 104.615
R1147 VDD1.n35 VDD1.n34 104.615
R1148 VDD1.n35 VDD1.n28 104.615
R1149 VDD1.n42 VDD1.n28 104.615
R1150 VDD1.n43 VDD1.n42 104.615
R1151 VDD1.n51 VDD1.n50 73.8769
R1152 VDD1.n24 VDD1.n23 73.5509
R1153 VDD1.n53 VDD1.n52 73.5507
R1154 VDD1.n49 VDD1.n48 73.5507
R1155 VDD1.n9 VDD1.t5 52.3082
R1156 VDD1.n34 VDD1.t8 52.3082
R1157 VDD1.n24 VDD1.n22 52.2818
R1158 VDD1.n49 VDD1.n47 52.2818
R1159 VDD1.n53 VDD1.n51 31.0289
R1160 VDD1.n8 VDD1.n7 15.6631
R1161 VDD1.n33 VDD1.n32 15.6631
R1162 VDD1.n11 VDD1.n6 12.8005
R1163 VDD1.n36 VDD1.n31 12.8005
R1164 VDD1.n12 VDD1.n4 12.0247
R1165 VDD1.n37 VDD1.n29 12.0247
R1166 VDD1.n16 VDD1.n15 11.249
R1167 VDD1.n41 VDD1.n40 11.249
R1168 VDD1.n19 VDD1.n2 10.4732
R1169 VDD1.n44 VDD1.n27 10.4732
R1170 VDD1.n20 VDD1.n0 9.69747
R1171 VDD1.n45 VDD1.n25 9.69747
R1172 VDD1.n22 VDD1.n21 9.45567
R1173 VDD1.n47 VDD1.n46 9.45567
R1174 VDD1.n21 VDD1.n20 9.3005
R1175 VDD1.n2 VDD1.n1 9.3005
R1176 VDD1.n15 VDD1.n14 9.3005
R1177 VDD1.n13 VDD1.n12 9.3005
R1178 VDD1.n6 VDD1.n5 9.3005
R1179 VDD1.n46 VDD1.n45 9.3005
R1180 VDD1.n27 VDD1.n26 9.3005
R1181 VDD1.n40 VDD1.n39 9.3005
R1182 VDD1.n38 VDD1.n37 9.3005
R1183 VDD1.n31 VDD1.n30 9.3005
R1184 VDD1.n7 VDD1.n5 4.39059
R1185 VDD1.n32 VDD1.n30 4.39059
R1186 VDD1.n22 VDD1.n0 4.26717
R1187 VDD1.n47 VDD1.n25 4.26717
R1188 VDD1.n52 VDD1.t7 4.20432
R1189 VDD1.n52 VDD1.t9 4.20432
R1190 VDD1.n23 VDD1.t3 4.20432
R1191 VDD1.n23 VDD1.t6 4.20432
R1192 VDD1.n50 VDD1.t2 4.20432
R1193 VDD1.n50 VDD1.t4 4.20432
R1194 VDD1.n48 VDD1.t0 4.20432
R1195 VDD1.n48 VDD1.t1 4.20432
R1196 VDD1.n20 VDD1.n19 3.49141
R1197 VDD1.n45 VDD1.n44 3.49141
R1198 VDD1.n16 VDD1.n2 2.71565
R1199 VDD1.n41 VDD1.n27 2.71565
R1200 VDD1.n15 VDD1.n4 1.93989
R1201 VDD1.n40 VDD1.n29 1.93989
R1202 VDD1.n12 VDD1.n11 1.16414
R1203 VDD1.n37 VDD1.n36 1.16414
R1204 VDD1.n8 VDD1.n6 0.388379
R1205 VDD1.n33 VDD1.n31 0.388379
R1206 VDD1 VDD1.n53 0.323776
R1207 VDD1 VDD1.n24 0.185845
R1208 VDD1.n21 VDD1.n1 0.155672
R1209 VDD1.n14 VDD1.n1 0.155672
R1210 VDD1.n14 VDD1.n13 0.155672
R1211 VDD1.n13 VDD1.n5 0.155672
R1212 VDD1.n38 VDD1.n30 0.155672
R1213 VDD1.n39 VDD1.n38 0.155672
R1214 VDD1.n39 VDD1.n26 0.155672
R1215 VDD1.n46 VDD1.n26 0.155672
R1216 VDD1.n51 VDD1.n49 0.0723091
C0 VDD1 VP 1.78617f
C1 VDD1 VDD2 0.69965f
C2 VN VTAIL 1.59448f
C3 VDD2 VP 0.288631f
C4 VN VDD1 0.151962f
C5 VDD1 VTAIL 9.98386f
C6 VN VP 3.60236f
C7 VN VDD2 1.65199f
C8 VTAIL VP 1.60885f
C9 VTAIL VDD2 10.018401f
C10 VDD2 B 3.122467f
C11 VDD1 B 3.031991f
C12 VTAIL B 3.381487f
C13 VN B 5.781529f
C14 VP B 4.811124f
C15 VDD1.n0 B 0.037392f
C16 VDD1.n1 B 0.025738f
C17 VDD1.n2 B 0.01383f
C18 VDD1.n3 B 0.03269f
C19 VDD1.n4 B 0.014644f
C20 VDD1.n5 B 0.458466f
C21 VDD1.n6 B 0.01383f
C22 VDD1.t5 B 0.053787f
C23 VDD1.n7 B 0.102988f
C24 VDD1.n8 B 0.019292f
C25 VDD1.n9 B 0.024517f
C26 VDD1.n10 B 0.03269f
C27 VDD1.n11 B 0.014644f
C28 VDD1.n12 B 0.01383f
C29 VDD1.n13 B 0.025738f
C30 VDD1.n14 B 0.025738f
C31 VDD1.n15 B 0.01383f
C32 VDD1.n16 B 0.014644f
C33 VDD1.n17 B 0.03269f
C34 VDD1.n18 B 0.072918f
C35 VDD1.n19 B 0.014644f
C36 VDD1.n20 B 0.01383f
C37 VDD1.n21 B 0.064766f
C38 VDD1.n22 B 0.059833f
C39 VDD1.t3 B 0.095796f
C40 VDD1.t6 B 0.095796f
C41 VDD1.n23 B 0.773078f
C42 VDD1.n24 B 0.355314f
C43 VDD1.n25 B 0.037392f
C44 VDD1.n26 B 0.025738f
C45 VDD1.n27 B 0.01383f
C46 VDD1.n28 B 0.03269f
C47 VDD1.n29 B 0.014644f
C48 VDD1.n30 B 0.458466f
C49 VDD1.n31 B 0.01383f
C50 VDD1.t8 B 0.053787f
C51 VDD1.n32 B 0.102988f
C52 VDD1.n33 B 0.019292f
C53 VDD1.n34 B 0.024517f
C54 VDD1.n35 B 0.03269f
C55 VDD1.n36 B 0.014644f
C56 VDD1.n37 B 0.01383f
C57 VDD1.n38 B 0.025738f
C58 VDD1.n39 B 0.025738f
C59 VDD1.n40 B 0.01383f
C60 VDD1.n41 B 0.014644f
C61 VDD1.n42 B 0.03269f
C62 VDD1.n43 B 0.072918f
C63 VDD1.n44 B 0.014644f
C64 VDD1.n45 B 0.01383f
C65 VDD1.n46 B 0.064766f
C66 VDD1.n47 B 0.059833f
C67 VDD1.t0 B 0.095796f
C68 VDD1.t1 B 0.095796f
C69 VDD1.n48 B 0.773074f
C70 VDD1.n49 B 0.354212f
C71 VDD1.t2 B 0.095796f
C72 VDD1.t4 B 0.095796f
C73 VDD1.n50 B 0.774334f
C74 VDD1.n51 B 1.33211f
C75 VDD1.t7 B 0.095796f
C76 VDD1.t9 B 0.095796f
C77 VDD1.n52 B 0.773074f
C78 VDD1.n53 B 1.66232f
C79 VP.n0 B 0.028874f
C80 VP.t7 B 0.101266f
C81 VP.t8 B 0.101266f
C82 VP.n1 B 0.011181f
C83 VP.n2 B 0.028874f
C84 VP.t2 B 0.101266f
C85 VP.t3 B 0.101266f
C86 VP.n3 B 0.011181f
C87 VP.t4 B 0.103518f
C88 VP.t6 B 0.101266f
C89 VP.n4 B 0.051119f
C90 VP.n5 B 0.059015f
C91 VP.n6 B 0.059847f
C92 VP.n7 B 0.028874f
C93 VP.n8 B 0.060697f
C94 VP.n9 B 0.011181f
C95 VP.n10 B 0.051119f
C96 VP.t0 B 0.103518f
C97 VP.n11 B 0.058979f
C98 VP.n12 B 0.85339f
C99 VP.t1 B 0.103518f
C100 VP.t9 B 0.101266f
C101 VP.n13 B 0.051119f
C102 VP.n14 B 0.058979f
C103 VP.n15 B 0.88317f
C104 VP.n16 B 0.028874f
C105 VP.n17 B 0.028874f
C106 VP.n18 B 0.060697f
C107 VP.n19 B 0.011181f
C108 VP.n20 B 0.051119f
C109 VP.t5 B 0.103518f
C110 VP.n21 B 0.058979f
C111 VP.n22 B 0.022376f
C112 VDD2.n0 B 0.037751f
C113 VDD2.n1 B 0.025985f
C114 VDD2.n2 B 0.013963f
C115 VDD2.n3 B 0.033004f
C116 VDD2.n4 B 0.014784f
C117 VDD2.n5 B 0.462866f
C118 VDD2.n6 B 0.013963f
C119 VDD2.t9 B 0.054303f
C120 VDD2.n7 B 0.103976f
C121 VDD2.n8 B 0.019477f
C122 VDD2.n9 B 0.024753f
C123 VDD2.n10 B 0.033004f
C124 VDD2.n11 B 0.014784f
C125 VDD2.n12 B 0.013963f
C126 VDD2.n13 B 0.025985f
C127 VDD2.n14 B 0.025985f
C128 VDD2.n15 B 0.013963f
C129 VDD2.n16 B 0.014784f
C130 VDD2.n17 B 0.033004f
C131 VDD2.n18 B 0.073618f
C132 VDD2.n19 B 0.014784f
C133 VDD2.n20 B 0.013963f
C134 VDD2.n21 B 0.065387f
C135 VDD2.n22 B 0.060407f
C136 VDD2.t4 B 0.096715f
C137 VDD2.t2 B 0.096715f
C138 VDD2.n23 B 0.780494f
C139 VDD2.n24 B 0.357611f
C140 VDD2.t0 B 0.096715f
C141 VDD2.t1 B 0.096715f
C142 VDD2.n25 B 0.781766f
C143 VDD2.n26 B 1.2773f
C144 VDD2.n27 B 0.037751f
C145 VDD2.n28 B 0.025985f
C146 VDD2.n29 B 0.013963f
C147 VDD2.n30 B 0.033004f
C148 VDD2.n31 B 0.014784f
C149 VDD2.n32 B 0.462866f
C150 VDD2.n33 B 0.013963f
C151 VDD2.t7 B 0.054303f
C152 VDD2.n34 B 0.103976f
C153 VDD2.n35 B 0.019477f
C154 VDD2.n36 B 0.024753f
C155 VDD2.n37 B 0.033004f
C156 VDD2.n38 B 0.014784f
C157 VDD2.n39 B 0.013963f
C158 VDD2.n40 B 0.025985f
C159 VDD2.n41 B 0.025985f
C160 VDD2.n42 B 0.013963f
C161 VDD2.n43 B 0.014784f
C162 VDD2.n44 B 0.033004f
C163 VDD2.n45 B 0.073618f
C164 VDD2.n46 B 0.014784f
C165 VDD2.n47 B 0.013963f
C166 VDD2.n48 B 0.065387f
C167 VDD2.n49 B 0.059476f
C168 VDD2.n50 B 1.45957f
C169 VDD2.t8 B 0.096715f
C170 VDD2.t6 B 0.096715f
C171 VDD2.n51 B 0.780497f
C172 VDD2.n52 B 0.263984f
C173 VDD2.t5 B 0.096715f
C174 VDD2.t3 B 0.096715f
C175 VDD2.n53 B 0.781745f
C176 VTAIL.t17 B 0.107662f
C177 VTAIL.t14 B 0.107662f
C178 VTAIL.n0 B 0.803239f
C179 VTAIL.n1 B 0.363942f
C180 VTAIL.n2 B 0.042024f
C181 VTAIL.n3 B 0.028926f
C182 VTAIL.n4 B 0.015544f
C183 VTAIL.n5 B 0.036739f
C184 VTAIL.n6 B 0.016458f
C185 VTAIL.n7 B 0.515258f
C186 VTAIL.n8 B 0.015544f
C187 VTAIL.t5 B 0.060449f
C188 VTAIL.n9 B 0.115745f
C189 VTAIL.n10 B 0.021681f
C190 VTAIL.n11 B 0.027555f
C191 VTAIL.n12 B 0.036739f
C192 VTAIL.n13 B 0.016458f
C193 VTAIL.n14 B 0.015544f
C194 VTAIL.n15 B 0.028926f
C195 VTAIL.n16 B 0.028926f
C196 VTAIL.n17 B 0.015544f
C197 VTAIL.n18 B 0.016458f
C198 VTAIL.n19 B 0.036739f
C199 VTAIL.n20 B 0.08195f
C200 VTAIL.n21 B 0.016458f
C201 VTAIL.n22 B 0.015544f
C202 VTAIL.n23 B 0.072788f
C203 VTAIL.n24 B 0.046278f
C204 VTAIL.n25 B 0.142958f
C205 VTAIL.t4 B 0.107662f
C206 VTAIL.t19 B 0.107662f
C207 VTAIL.n26 B 0.803239f
C208 VTAIL.n27 B 0.350282f
C209 VTAIL.t7 B 0.107662f
C210 VTAIL.t3 B 0.107662f
C211 VTAIL.n28 B 0.803239f
C212 VTAIL.n29 B 1.16906f
C213 VTAIL.t18 B 0.107662f
C214 VTAIL.t13 B 0.107662f
C215 VTAIL.n30 B 0.803244f
C216 VTAIL.n31 B 1.16906f
C217 VTAIL.t15 B 0.107662f
C218 VTAIL.t9 B 0.107662f
C219 VTAIL.n32 B 0.803244f
C220 VTAIL.n33 B 0.350277f
C221 VTAIL.n34 B 0.042024f
C222 VTAIL.n35 B 0.028926f
C223 VTAIL.n36 B 0.015544f
C224 VTAIL.n37 B 0.036739f
C225 VTAIL.n38 B 0.016458f
C226 VTAIL.n39 B 0.515258f
C227 VTAIL.n40 B 0.015544f
C228 VTAIL.t16 B 0.060449f
C229 VTAIL.n41 B 0.115745f
C230 VTAIL.n42 B 0.021681f
C231 VTAIL.n43 B 0.027555f
C232 VTAIL.n44 B 0.036739f
C233 VTAIL.n45 B 0.016458f
C234 VTAIL.n46 B 0.015544f
C235 VTAIL.n47 B 0.028926f
C236 VTAIL.n48 B 0.028926f
C237 VTAIL.n49 B 0.015544f
C238 VTAIL.n50 B 0.016458f
C239 VTAIL.n51 B 0.036739f
C240 VTAIL.n52 B 0.08195f
C241 VTAIL.n53 B 0.016458f
C242 VTAIL.n54 B 0.015544f
C243 VTAIL.n55 B 0.072788f
C244 VTAIL.n56 B 0.046278f
C245 VTAIL.n57 B 0.142958f
C246 VTAIL.t2 B 0.107662f
C247 VTAIL.t8 B 0.107662f
C248 VTAIL.n58 B 0.803244f
C249 VTAIL.n59 B 0.370365f
C250 VTAIL.t1 B 0.107662f
C251 VTAIL.t0 B 0.107662f
C252 VTAIL.n60 B 0.803244f
C253 VTAIL.n61 B 0.350277f
C254 VTAIL.n62 B 0.042024f
C255 VTAIL.n63 B 0.028926f
C256 VTAIL.n64 B 0.015544f
C257 VTAIL.n65 B 0.036739f
C258 VTAIL.n66 B 0.016458f
C259 VTAIL.n67 B 0.515258f
C260 VTAIL.n68 B 0.015544f
C261 VTAIL.t6 B 0.060449f
C262 VTAIL.n69 B 0.115745f
C263 VTAIL.n70 B 0.021681f
C264 VTAIL.n71 B 0.027555f
C265 VTAIL.n72 B 0.036739f
C266 VTAIL.n73 B 0.016458f
C267 VTAIL.n74 B 0.015544f
C268 VTAIL.n75 B 0.028926f
C269 VTAIL.n76 B 0.028926f
C270 VTAIL.n77 B 0.015544f
C271 VTAIL.n78 B 0.016458f
C272 VTAIL.n79 B 0.036739f
C273 VTAIL.n80 B 0.08195f
C274 VTAIL.n81 B 0.016458f
C275 VTAIL.n82 B 0.015544f
C276 VTAIL.n83 B 0.072788f
C277 VTAIL.n84 B 0.046278f
C278 VTAIL.n85 B 0.894244f
C279 VTAIL.n86 B 0.042024f
C280 VTAIL.n87 B 0.028926f
C281 VTAIL.n88 B 0.015544f
C282 VTAIL.n89 B 0.036739f
C283 VTAIL.n90 B 0.016458f
C284 VTAIL.n91 B 0.515258f
C285 VTAIL.n92 B 0.015544f
C286 VTAIL.t10 B 0.060449f
C287 VTAIL.n93 B 0.115745f
C288 VTAIL.n94 B 0.021681f
C289 VTAIL.n95 B 0.027555f
C290 VTAIL.n96 B 0.036739f
C291 VTAIL.n97 B 0.016458f
C292 VTAIL.n98 B 0.015544f
C293 VTAIL.n99 B 0.028926f
C294 VTAIL.n100 B 0.028926f
C295 VTAIL.n101 B 0.015544f
C296 VTAIL.n102 B 0.016458f
C297 VTAIL.n103 B 0.036739f
C298 VTAIL.n104 B 0.08195f
C299 VTAIL.n105 B 0.016458f
C300 VTAIL.n106 B 0.015544f
C301 VTAIL.n107 B 0.072788f
C302 VTAIL.n108 B 0.046278f
C303 VTAIL.n109 B 0.894244f
C304 VTAIL.t11 B 0.107662f
C305 VTAIL.t12 B 0.107662f
C306 VTAIL.n110 B 0.803239f
C307 VTAIL.n111 B 0.309304f
C308 VN.n0 B 0.028552f
C309 VN.t9 B 0.100137f
C310 VN.t7 B 0.100137f
C311 VN.n1 B 0.011056f
C312 VN.t0 B 0.102364f
C313 VN.t5 B 0.100137f
C314 VN.n2 B 0.050549f
C315 VN.n3 B 0.058357f
C316 VN.n4 B 0.05918f
C317 VN.n5 B 0.028552f
C318 VN.n6 B 0.06002f
C319 VN.n7 B 0.011056f
C320 VN.n8 B 0.050549f
C321 VN.t8 B 0.102364f
C322 VN.n9 B 0.058322f
C323 VN.n10 B 0.022127f
C324 VN.n11 B 0.028552f
C325 VN.t2 B 0.102364f
C326 VN.t1 B 0.100137f
C327 VN.t3 B 0.100137f
C328 VN.n12 B 0.011056f
C329 VN.t4 B 0.100137f
C330 VN.n13 B 0.050549f
C331 VN.t6 B 0.102364f
C332 VN.n14 B 0.058357f
C333 VN.n15 B 0.05918f
C334 VN.n16 B 0.028552f
C335 VN.n17 B 0.06002f
C336 VN.n18 B 0.011056f
C337 VN.n19 B 0.050549f
C338 VN.n20 B 0.058322f
C339 VN.n21 B 0.862859f
.ends

