* NGSPICE file created from diff_pair_sample_0812.ext - technology: sky130A

.subckt diff_pair_sample_0812 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t12 w_n4190_n4774# sky130_fd_pr__pfet_01v8 ad=3.13995 pd=19.36 as=3.13995 ps=19.36 w=19.03 l=2.89
X1 VTAIL.t7 VN.t0 VDD2.t7 w_n4190_n4774# sky130_fd_pr__pfet_01v8 ad=3.13995 pd=19.36 as=3.13995 ps=19.36 w=19.03 l=2.89
X2 VTAIL.t6 VN.t1 VDD2.t6 w_n4190_n4774# sky130_fd_pr__pfet_01v8 ad=7.4217 pd=38.84 as=3.13995 ps=19.36 w=19.03 l=2.89
X3 VDD2.t5 VN.t2 VTAIL.t0 w_n4190_n4774# sky130_fd_pr__pfet_01v8 ad=3.13995 pd=19.36 as=7.4217 ps=38.84 w=19.03 l=2.89
X4 VTAIL.t11 VP.t1 VDD1.t6 w_n4190_n4774# sky130_fd_pr__pfet_01v8 ad=7.4217 pd=38.84 as=3.13995 ps=19.36 w=19.03 l=2.89
X5 VDD1.t5 VP.t2 VTAIL.t14 w_n4190_n4774# sky130_fd_pr__pfet_01v8 ad=3.13995 pd=19.36 as=7.4217 ps=38.84 w=19.03 l=2.89
X6 VTAIL.t3 VN.t3 VDD2.t4 w_n4190_n4774# sky130_fd_pr__pfet_01v8 ad=3.13995 pd=19.36 as=3.13995 ps=19.36 w=19.03 l=2.89
X7 VTAIL.t9 VP.t3 VDD1.t4 w_n4190_n4774# sky130_fd_pr__pfet_01v8 ad=3.13995 pd=19.36 as=3.13995 ps=19.36 w=19.03 l=2.89
X8 VDD2.t3 VN.t4 VTAIL.t4 w_n4190_n4774# sky130_fd_pr__pfet_01v8 ad=3.13995 pd=19.36 as=7.4217 ps=38.84 w=19.03 l=2.89
X9 VDD1.t3 VP.t4 VTAIL.t10 w_n4190_n4774# sky130_fd_pr__pfet_01v8 ad=3.13995 pd=19.36 as=3.13995 ps=19.36 w=19.03 l=2.89
X10 VDD2.t2 VN.t5 VTAIL.t1 w_n4190_n4774# sky130_fd_pr__pfet_01v8 ad=3.13995 pd=19.36 as=3.13995 ps=19.36 w=19.03 l=2.89
X11 VDD1.t2 VP.t5 VTAIL.t8 w_n4190_n4774# sky130_fd_pr__pfet_01v8 ad=3.13995 pd=19.36 as=7.4217 ps=38.84 w=19.03 l=2.89
X12 B.t11 B.t9 B.t10 w_n4190_n4774# sky130_fd_pr__pfet_01v8 ad=7.4217 pd=38.84 as=0 ps=0 w=19.03 l=2.89
X13 VDD2.t1 VN.t6 VTAIL.t2 w_n4190_n4774# sky130_fd_pr__pfet_01v8 ad=3.13995 pd=19.36 as=3.13995 ps=19.36 w=19.03 l=2.89
X14 VTAIL.t5 VN.t7 VDD2.t0 w_n4190_n4774# sky130_fd_pr__pfet_01v8 ad=7.4217 pd=38.84 as=3.13995 ps=19.36 w=19.03 l=2.89
X15 B.t8 B.t6 B.t7 w_n4190_n4774# sky130_fd_pr__pfet_01v8 ad=7.4217 pd=38.84 as=0 ps=0 w=19.03 l=2.89
X16 VTAIL.t13 VP.t6 VDD1.t1 w_n4190_n4774# sky130_fd_pr__pfet_01v8 ad=7.4217 pd=38.84 as=3.13995 ps=19.36 w=19.03 l=2.89
X17 B.t5 B.t3 B.t4 w_n4190_n4774# sky130_fd_pr__pfet_01v8 ad=7.4217 pd=38.84 as=0 ps=0 w=19.03 l=2.89
X18 VTAIL.t15 VP.t7 VDD1.t0 w_n4190_n4774# sky130_fd_pr__pfet_01v8 ad=3.13995 pd=19.36 as=3.13995 ps=19.36 w=19.03 l=2.89
X19 B.t2 B.t0 B.t1 w_n4190_n4774# sky130_fd_pr__pfet_01v8 ad=7.4217 pd=38.84 as=0 ps=0 w=19.03 l=2.89
R0 VP.n17 VP.t6 192.218
R1 VP.n19 VP.n16 161.3
R2 VP.n21 VP.n20 161.3
R3 VP.n22 VP.n15 161.3
R4 VP.n24 VP.n23 161.3
R5 VP.n25 VP.n14 161.3
R6 VP.n28 VP.n27 161.3
R7 VP.n29 VP.n13 161.3
R8 VP.n31 VP.n30 161.3
R9 VP.n32 VP.n12 161.3
R10 VP.n34 VP.n33 161.3
R11 VP.n35 VP.n11 161.3
R12 VP.n37 VP.n36 161.3
R13 VP.n38 VP.n10 161.3
R14 VP.n74 VP.n0 161.3
R15 VP.n73 VP.n72 161.3
R16 VP.n71 VP.n1 161.3
R17 VP.n70 VP.n69 161.3
R18 VP.n68 VP.n2 161.3
R19 VP.n67 VP.n66 161.3
R20 VP.n65 VP.n3 161.3
R21 VP.n64 VP.n63 161.3
R22 VP.n61 VP.n4 161.3
R23 VP.n60 VP.n59 161.3
R24 VP.n58 VP.n5 161.3
R25 VP.n57 VP.n56 161.3
R26 VP.n55 VP.n6 161.3
R27 VP.n53 VP.n52 161.3
R28 VP.n51 VP.n7 161.3
R29 VP.n50 VP.n49 161.3
R30 VP.n48 VP.n8 161.3
R31 VP.n47 VP.n46 161.3
R32 VP.n45 VP.n9 161.3
R33 VP.n44 VP.n43 161.3
R34 VP.n42 VP.t1 158.694
R35 VP.n54 VP.t0 158.694
R36 VP.n62 VP.t7 158.694
R37 VP.n75 VP.t5 158.694
R38 VP.n39 VP.t2 158.694
R39 VP.n26 VP.t3 158.694
R40 VP.n18 VP.t4 158.694
R41 VP.n42 VP.n41 106.841
R42 VP.n76 VP.n75 106.841
R43 VP.n40 VP.n39 106.841
R44 VP.n41 VP.n40 57.5753
R45 VP.n60 VP.n5 56.5193
R46 VP.n24 VP.n15 56.5193
R47 VP.n18 VP.n17 56.0641
R48 VP.n49 VP.n48 43.4072
R49 VP.n69 VP.n68 43.4072
R50 VP.n33 VP.n32 43.4072
R51 VP.n48 VP.n47 37.5796
R52 VP.n69 VP.n1 37.5796
R53 VP.n33 VP.n11 37.5796
R54 VP.n43 VP.n9 24.4675
R55 VP.n47 VP.n9 24.4675
R56 VP.n49 VP.n7 24.4675
R57 VP.n53 VP.n7 24.4675
R58 VP.n56 VP.n55 24.4675
R59 VP.n56 VP.n5 24.4675
R60 VP.n61 VP.n60 24.4675
R61 VP.n63 VP.n61 24.4675
R62 VP.n67 VP.n3 24.4675
R63 VP.n68 VP.n67 24.4675
R64 VP.n73 VP.n1 24.4675
R65 VP.n74 VP.n73 24.4675
R66 VP.n37 VP.n11 24.4675
R67 VP.n38 VP.n37 24.4675
R68 VP.n25 VP.n24 24.4675
R69 VP.n27 VP.n25 24.4675
R70 VP.n31 VP.n13 24.4675
R71 VP.n32 VP.n31 24.4675
R72 VP.n20 VP.n19 24.4675
R73 VP.n20 VP.n15 24.4675
R74 VP.n55 VP.n54 17.6167
R75 VP.n63 VP.n62 17.6167
R76 VP.n27 VP.n26 17.6167
R77 VP.n19 VP.n18 17.6167
R78 VP.n54 VP.n53 6.85126
R79 VP.n62 VP.n3 6.85126
R80 VP.n26 VP.n13 6.85126
R81 VP.n17 VP.n16 5.02778
R82 VP.n43 VP.n42 3.91522
R83 VP.n75 VP.n74 3.91522
R84 VP.n39 VP.n38 3.91522
R85 VP.n40 VP.n10 0.278367
R86 VP.n44 VP.n41 0.278367
R87 VP.n76 VP.n0 0.278367
R88 VP.n21 VP.n16 0.189894
R89 VP.n22 VP.n21 0.189894
R90 VP.n23 VP.n22 0.189894
R91 VP.n23 VP.n14 0.189894
R92 VP.n28 VP.n14 0.189894
R93 VP.n29 VP.n28 0.189894
R94 VP.n30 VP.n29 0.189894
R95 VP.n30 VP.n12 0.189894
R96 VP.n34 VP.n12 0.189894
R97 VP.n35 VP.n34 0.189894
R98 VP.n36 VP.n35 0.189894
R99 VP.n36 VP.n10 0.189894
R100 VP.n45 VP.n44 0.189894
R101 VP.n46 VP.n45 0.189894
R102 VP.n46 VP.n8 0.189894
R103 VP.n50 VP.n8 0.189894
R104 VP.n51 VP.n50 0.189894
R105 VP.n52 VP.n51 0.189894
R106 VP.n52 VP.n6 0.189894
R107 VP.n57 VP.n6 0.189894
R108 VP.n58 VP.n57 0.189894
R109 VP.n59 VP.n58 0.189894
R110 VP.n59 VP.n4 0.189894
R111 VP.n64 VP.n4 0.189894
R112 VP.n65 VP.n64 0.189894
R113 VP.n66 VP.n65 0.189894
R114 VP.n66 VP.n2 0.189894
R115 VP.n70 VP.n2 0.189894
R116 VP.n71 VP.n70 0.189894
R117 VP.n72 VP.n71 0.189894
R118 VP.n72 VP.n0 0.189894
R119 VP VP.n76 0.153454
R120 VTAIL.n850 VTAIL.n750 756.745
R121 VTAIL.n102 VTAIL.n2 756.745
R122 VTAIL.n208 VTAIL.n108 756.745
R123 VTAIL.n316 VTAIL.n216 756.745
R124 VTAIL.n744 VTAIL.n644 756.745
R125 VTAIL.n636 VTAIL.n536 756.745
R126 VTAIL.n530 VTAIL.n430 756.745
R127 VTAIL.n422 VTAIL.n322 756.745
R128 VTAIL.n785 VTAIL.n784 585
R129 VTAIL.n782 VTAIL.n781 585
R130 VTAIL.n791 VTAIL.n790 585
R131 VTAIL.n793 VTAIL.n792 585
R132 VTAIL.n778 VTAIL.n777 585
R133 VTAIL.n799 VTAIL.n798 585
R134 VTAIL.n801 VTAIL.n800 585
R135 VTAIL.n774 VTAIL.n773 585
R136 VTAIL.n807 VTAIL.n806 585
R137 VTAIL.n809 VTAIL.n808 585
R138 VTAIL.n770 VTAIL.n769 585
R139 VTAIL.n815 VTAIL.n814 585
R140 VTAIL.n817 VTAIL.n816 585
R141 VTAIL.n766 VTAIL.n765 585
R142 VTAIL.n823 VTAIL.n822 585
R143 VTAIL.n826 VTAIL.n825 585
R144 VTAIL.n824 VTAIL.n762 585
R145 VTAIL.n831 VTAIL.n761 585
R146 VTAIL.n833 VTAIL.n832 585
R147 VTAIL.n835 VTAIL.n834 585
R148 VTAIL.n758 VTAIL.n757 585
R149 VTAIL.n841 VTAIL.n840 585
R150 VTAIL.n843 VTAIL.n842 585
R151 VTAIL.n754 VTAIL.n753 585
R152 VTAIL.n849 VTAIL.n848 585
R153 VTAIL.n851 VTAIL.n850 585
R154 VTAIL.n37 VTAIL.n36 585
R155 VTAIL.n34 VTAIL.n33 585
R156 VTAIL.n43 VTAIL.n42 585
R157 VTAIL.n45 VTAIL.n44 585
R158 VTAIL.n30 VTAIL.n29 585
R159 VTAIL.n51 VTAIL.n50 585
R160 VTAIL.n53 VTAIL.n52 585
R161 VTAIL.n26 VTAIL.n25 585
R162 VTAIL.n59 VTAIL.n58 585
R163 VTAIL.n61 VTAIL.n60 585
R164 VTAIL.n22 VTAIL.n21 585
R165 VTAIL.n67 VTAIL.n66 585
R166 VTAIL.n69 VTAIL.n68 585
R167 VTAIL.n18 VTAIL.n17 585
R168 VTAIL.n75 VTAIL.n74 585
R169 VTAIL.n78 VTAIL.n77 585
R170 VTAIL.n76 VTAIL.n14 585
R171 VTAIL.n83 VTAIL.n13 585
R172 VTAIL.n85 VTAIL.n84 585
R173 VTAIL.n87 VTAIL.n86 585
R174 VTAIL.n10 VTAIL.n9 585
R175 VTAIL.n93 VTAIL.n92 585
R176 VTAIL.n95 VTAIL.n94 585
R177 VTAIL.n6 VTAIL.n5 585
R178 VTAIL.n101 VTAIL.n100 585
R179 VTAIL.n103 VTAIL.n102 585
R180 VTAIL.n143 VTAIL.n142 585
R181 VTAIL.n140 VTAIL.n139 585
R182 VTAIL.n149 VTAIL.n148 585
R183 VTAIL.n151 VTAIL.n150 585
R184 VTAIL.n136 VTAIL.n135 585
R185 VTAIL.n157 VTAIL.n156 585
R186 VTAIL.n159 VTAIL.n158 585
R187 VTAIL.n132 VTAIL.n131 585
R188 VTAIL.n165 VTAIL.n164 585
R189 VTAIL.n167 VTAIL.n166 585
R190 VTAIL.n128 VTAIL.n127 585
R191 VTAIL.n173 VTAIL.n172 585
R192 VTAIL.n175 VTAIL.n174 585
R193 VTAIL.n124 VTAIL.n123 585
R194 VTAIL.n181 VTAIL.n180 585
R195 VTAIL.n184 VTAIL.n183 585
R196 VTAIL.n182 VTAIL.n120 585
R197 VTAIL.n189 VTAIL.n119 585
R198 VTAIL.n191 VTAIL.n190 585
R199 VTAIL.n193 VTAIL.n192 585
R200 VTAIL.n116 VTAIL.n115 585
R201 VTAIL.n199 VTAIL.n198 585
R202 VTAIL.n201 VTAIL.n200 585
R203 VTAIL.n112 VTAIL.n111 585
R204 VTAIL.n207 VTAIL.n206 585
R205 VTAIL.n209 VTAIL.n208 585
R206 VTAIL.n251 VTAIL.n250 585
R207 VTAIL.n248 VTAIL.n247 585
R208 VTAIL.n257 VTAIL.n256 585
R209 VTAIL.n259 VTAIL.n258 585
R210 VTAIL.n244 VTAIL.n243 585
R211 VTAIL.n265 VTAIL.n264 585
R212 VTAIL.n267 VTAIL.n266 585
R213 VTAIL.n240 VTAIL.n239 585
R214 VTAIL.n273 VTAIL.n272 585
R215 VTAIL.n275 VTAIL.n274 585
R216 VTAIL.n236 VTAIL.n235 585
R217 VTAIL.n281 VTAIL.n280 585
R218 VTAIL.n283 VTAIL.n282 585
R219 VTAIL.n232 VTAIL.n231 585
R220 VTAIL.n289 VTAIL.n288 585
R221 VTAIL.n292 VTAIL.n291 585
R222 VTAIL.n290 VTAIL.n228 585
R223 VTAIL.n297 VTAIL.n227 585
R224 VTAIL.n299 VTAIL.n298 585
R225 VTAIL.n301 VTAIL.n300 585
R226 VTAIL.n224 VTAIL.n223 585
R227 VTAIL.n307 VTAIL.n306 585
R228 VTAIL.n309 VTAIL.n308 585
R229 VTAIL.n220 VTAIL.n219 585
R230 VTAIL.n315 VTAIL.n314 585
R231 VTAIL.n317 VTAIL.n316 585
R232 VTAIL.n745 VTAIL.n744 585
R233 VTAIL.n743 VTAIL.n742 585
R234 VTAIL.n648 VTAIL.n647 585
R235 VTAIL.n737 VTAIL.n736 585
R236 VTAIL.n735 VTAIL.n734 585
R237 VTAIL.n652 VTAIL.n651 585
R238 VTAIL.n729 VTAIL.n728 585
R239 VTAIL.n727 VTAIL.n726 585
R240 VTAIL.n725 VTAIL.n655 585
R241 VTAIL.n659 VTAIL.n656 585
R242 VTAIL.n720 VTAIL.n719 585
R243 VTAIL.n718 VTAIL.n717 585
R244 VTAIL.n661 VTAIL.n660 585
R245 VTAIL.n712 VTAIL.n711 585
R246 VTAIL.n710 VTAIL.n709 585
R247 VTAIL.n665 VTAIL.n664 585
R248 VTAIL.n704 VTAIL.n703 585
R249 VTAIL.n702 VTAIL.n701 585
R250 VTAIL.n669 VTAIL.n668 585
R251 VTAIL.n696 VTAIL.n695 585
R252 VTAIL.n694 VTAIL.n693 585
R253 VTAIL.n673 VTAIL.n672 585
R254 VTAIL.n688 VTAIL.n687 585
R255 VTAIL.n686 VTAIL.n685 585
R256 VTAIL.n677 VTAIL.n676 585
R257 VTAIL.n680 VTAIL.n679 585
R258 VTAIL.n637 VTAIL.n636 585
R259 VTAIL.n635 VTAIL.n634 585
R260 VTAIL.n540 VTAIL.n539 585
R261 VTAIL.n629 VTAIL.n628 585
R262 VTAIL.n627 VTAIL.n626 585
R263 VTAIL.n544 VTAIL.n543 585
R264 VTAIL.n621 VTAIL.n620 585
R265 VTAIL.n619 VTAIL.n618 585
R266 VTAIL.n617 VTAIL.n547 585
R267 VTAIL.n551 VTAIL.n548 585
R268 VTAIL.n612 VTAIL.n611 585
R269 VTAIL.n610 VTAIL.n609 585
R270 VTAIL.n553 VTAIL.n552 585
R271 VTAIL.n604 VTAIL.n603 585
R272 VTAIL.n602 VTAIL.n601 585
R273 VTAIL.n557 VTAIL.n556 585
R274 VTAIL.n596 VTAIL.n595 585
R275 VTAIL.n594 VTAIL.n593 585
R276 VTAIL.n561 VTAIL.n560 585
R277 VTAIL.n588 VTAIL.n587 585
R278 VTAIL.n586 VTAIL.n585 585
R279 VTAIL.n565 VTAIL.n564 585
R280 VTAIL.n580 VTAIL.n579 585
R281 VTAIL.n578 VTAIL.n577 585
R282 VTAIL.n569 VTAIL.n568 585
R283 VTAIL.n572 VTAIL.n571 585
R284 VTAIL.n531 VTAIL.n530 585
R285 VTAIL.n529 VTAIL.n528 585
R286 VTAIL.n434 VTAIL.n433 585
R287 VTAIL.n523 VTAIL.n522 585
R288 VTAIL.n521 VTAIL.n520 585
R289 VTAIL.n438 VTAIL.n437 585
R290 VTAIL.n515 VTAIL.n514 585
R291 VTAIL.n513 VTAIL.n512 585
R292 VTAIL.n511 VTAIL.n441 585
R293 VTAIL.n445 VTAIL.n442 585
R294 VTAIL.n506 VTAIL.n505 585
R295 VTAIL.n504 VTAIL.n503 585
R296 VTAIL.n447 VTAIL.n446 585
R297 VTAIL.n498 VTAIL.n497 585
R298 VTAIL.n496 VTAIL.n495 585
R299 VTAIL.n451 VTAIL.n450 585
R300 VTAIL.n490 VTAIL.n489 585
R301 VTAIL.n488 VTAIL.n487 585
R302 VTAIL.n455 VTAIL.n454 585
R303 VTAIL.n482 VTAIL.n481 585
R304 VTAIL.n480 VTAIL.n479 585
R305 VTAIL.n459 VTAIL.n458 585
R306 VTAIL.n474 VTAIL.n473 585
R307 VTAIL.n472 VTAIL.n471 585
R308 VTAIL.n463 VTAIL.n462 585
R309 VTAIL.n466 VTAIL.n465 585
R310 VTAIL.n423 VTAIL.n422 585
R311 VTAIL.n421 VTAIL.n420 585
R312 VTAIL.n326 VTAIL.n325 585
R313 VTAIL.n415 VTAIL.n414 585
R314 VTAIL.n413 VTAIL.n412 585
R315 VTAIL.n330 VTAIL.n329 585
R316 VTAIL.n407 VTAIL.n406 585
R317 VTAIL.n405 VTAIL.n404 585
R318 VTAIL.n403 VTAIL.n333 585
R319 VTAIL.n337 VTAIL.n334 585
R320 VTAIL.n398 VTAIL.n397 585
R321 VTAIL.n396 VTAIL.n395 585
R322 VTAIL.n339 VTAIL.n338 585
R323 VTAIL.n390 VTAIL.n389 585
R324 VTAIL.n388 VTAIL.n387 585
R325 VTAIL.n343 VTAIL.n342 585
R326 VTAIL.n382 VTAIL.n381 585
R327 VTAIL.n380 VTAIL.n379 585
R328 VTAIL.n347 VTAIL.n346 585
R329 VTAIL.n374 VTAIL.n373 585
R330 VTAIL.n372 VTAIL.n371 585
R331 VTAIL.n351 VTAIL.n350 585
R332 VTAIL.n366 VTAIL.n365 585
R333 VTAIL.n364 VTAIL.n363 585
R334 VTAIL.n355 VTAIL.n354 585
R335 VTAIL.n358 VTAIL.n357 585
R336 VTAIL.t14 VTAIL.n678 327.466
R337 VTAIL.t13 VTAIL.n570 327.466
R338 VTAIL.t4 VTAIL.n464 327.466
R339 VTAIL.t6 VTAIL.n356 327.466
R340 VTAIL.t0 VTAIL.n783 327.466
R341 VTAIL.t5 VTAIL.n35 327.466
R342 VTAIL.t8 VTAIL.n141 327.466
R343 VTAIL.t11 VTAIL.n249 327.466
R344 VTAIL.n784 VTAIL.n781 171.744
R345 VTAIL.n791 VTAIL.n781 171.744
R346 VTAIL.n792 VTAIL.n791 171.744
R347 VTAIL.n792 VTAIL.n777 171.744
R348 VTAIL.n799 VTAIL.n777 171.744
R349 VTAIL.n800 VTAIL.n799 171.744
R350 VTAIL.n800 VTAIL.n773 171.744
R351 VTAIL.n807 VTAIL.n773 171.744
R352 VTAIL.n808 VTAIL.n807 171.744
R353 VTAIL.n808 VTAIL.n769 171.744
R354 VTAIL.n815 VTAIL.n769 171.744
R355 VTAIL.n816 VTAIL.n815 171.744
R356 VTAIL.n816 VTAIL.n765 171.744
R357 VTAIL.n823 VTAIL.n765 171.744
R358 VTAIL.n825 VTAIL.n823 171.744
R359 VTAIL.n825 VTAIL.n824 171.744
R360 VTAIL.n824 VTAIL.n761 171.744
R361 VTAIL.n833 VTAIL.n761 171.744
R362 VTAIL.n834 VTAIL.n833 171.744
R363 VTAIL.n834 VTAIL.n757 171.744
R364 VTAIL.n841 VTAIL.n757 171.744
R365 VTAIL.n842 VTAIL.n841 171.744
R366 VTAIL.n842 VTAIL.n753 171.744
R367 VTAIL.n849 VTAIL.n753 171.744
R368 VTAIL.n850 VTAIL.n849 171.744
R369 VTAIL.n36 VTAIL.n33 171.744
R370 VTAIL.n43 VTAIL.n33 171.744
R371 VTAIL.n44 VTAIL.n43 171.744
R372 VTAIL.n44 VTAIL.n29 171.744
R373 VTAIL.n51 VTAIL.n29 171.744
R374 VTAIL.n52 VTAIL.n51 171.744
R375 VTAIL.n52 VTAIL.n25 171.744
R376 VTAIL.n59 VTAIL.n25 171.744
R377 VTAIL.n60 VTAIL.n59 171.744
R378 VTAIL.n60 VTAIL.n21 171.744
R379 VTAIL.n67 VTAIL.n21 171.744
R380 VTAIL.n68 VTAIL.n67 171.744
R381 VTAIL.n68 VTAIL.n17 171.744
R382 VTAIL.n75 VTAIL.n17 171.744
R383 VTAIL.n77 VTAIL.n75 171.744
R384 VTAIL.n77 VTAIL.n76 171.744
R385 VTAIL.n76 VTAIL.n13 171.744
R386 VTAIL.n85 VTAIL.n13 171.744
R387 VTAIL.n86 VTAIL.n85 171.744
R388 VTAIL.n86 VTAIL.n9 171.744
R389 VTAIL.n93 VTAIL.n9 171.744
R390 VTAIL.n94 VTAIL.n93 171.744
R391 VTAIL.n94 VTAIL.n5 171.744
R392 VTAIL.n101 VTAIL.n5 171.744
R393 VTAIL.n102 VTAIL.n101 171.744
R394 VTAIL.n142 VTAIL.n139 171.744
R395 VTAIL.n149 VTAIL.n139 171.744
R396 VTAIL.n150 VTAIL.n149 171.744
R397 VTAIL.n150 VTAIL.n135 171.744
R398 VTAIL.n157 VTAIL.n135 171.744
R399 VTAIL.n158 VTAIL.n157 171.744
R400 VTAIL.n158 VTAIL.n131 171.744
R401 VTAIL.n165 VTAIL.n131 171.744
R402 VTAIL.n166 VTAIL.n165 171.744
R403 VTAIL.n166 VTAIL.n127 171.744
R404 VTAIL.n173 VTAIL.n127 171.744
R405 VTAIL.n174 VTAIL.n173 171.744
R406 VTAIL.n174 VTAIL.n123 171.744
R407 VTAIL.n181 VTAIL.n123 171.744
R408 VTAIL.n183 VTAIL.n181 171.744
R409 VTAIL.n183 VTAIL.n182 171.744
R410 VTAIL.n182 VTAIL.n119 171.744
R411 VTAIL.n191 VTAIL.n119 171.744
R412 VTAIL.n192 VTAIL.n191 171.744
R413 VTAIL.n192 VTAIL.n115 171.744
R414 VTAIL.n199 VTAIL.n115 171.744
R415 VTAIL.n200 VTAIL.n199 171.744
R416 VTAIL.n200 VTAIL.n111 171.744
R417 VTAIL.n207 VTAIL.n111 171.744
R418 VTAIL.n208 VTAIL.n207 171.744
R419 VTAIL.n250 VTAIL.n247 171.744
R420 VTAIL.n257 VTAIL.n247 171.744
R421 VTAIL.n258 VTAIL.n257 171.744
R422 VTAIL.n258 VTAIL.n243 171.744
R423 VTAIL.n265 VTAIL.n243 171.744
R424 VTAIL.n266 VTAIL.n265 171.744
R425 VTAIL.n266 VTAIL.n239 171.744
R426 VTAIL.n273 VTAIL.n239 171.744
R427 VTAIL.n274 VTAIL.n273 171.744
R428 VTAIL.n274 VTAIL.n235 171.744
R429 VTAIL.n281 VTAIL.n235 171.744
R430 VTAIL.n282 VTAIL.n281 171.744
R431 VTAIL.n282 VTAIL.n231 171.744
R432 VTAIL.n289 VTAIL.n231 171.744
R433 VTAIL.n291 VTAIL.n289 171.744
R434 VTAIL.n291 VTAIL.n290 171.744
R435 VTAIL.n290 VTAIL.n227 171.744
R436 VTAIL.n299 VTAIL.n227 171.744
R437 VTAIL.n300 VTAIL.n299 171.744
R438 VTAIL.n300 VTAIL.n223 171.744
R439 VTAIL.n307 VTAIL.n223 171.744
R440 VTAIL.n308 VTAIL.n307 171.744
R441 VTAIL.n308 VTAIL.n219 171.744
R442 VTAIL.n315 VTAIL.n219 171.744
R443 VTAIL.n316 VTAIL.n315 171.744
R444 VTAIL.n744 VTAIL.n743 171.744
R445 VTAIL.n743 VTAIL.n647 171.744
R446 VTAIL.n736 VTAIL.n647 171.744
R447 VTAIL.n736 VTAIL.n735 171.744
R448 VTAIL.n735 VTAIL.n651 171.744
R449 VTAIL.n728 VTAIL.n651 171.744
R450 VTAIL.n728 VTAIL.n727 171.744
R451 VTAIL.n727 VTAIL.n655 171.744
R452 VTAIL.n659 VTAIL.n655 171.744
R453 VTAIL.n719 VTAIL.n659 171.744
R454 VTAIL.n719 VTAIL.n718 171.744
R455 VTAIL.n718 VTAIL.n660 171.744
R456 VTAIL.n711 VTAIL.n660 171.744
R457 VTAIL.n711 VTAIL.n710 171.744
R458 VTAIL.n710 VTAIL.n664 171.744
R459 VTAIL.n703 VTAIL.n664 171.744
R460 VTAIL.n703 VTAIL.n702 171.744
R461 VTAIL.n702 VTAIL.n668 171.744
R462 VTAIL.n695 VTAIL.n668 171.744
R463 VTAIL.n695 VTAIL.n694 171.744
R464 VTAIL.n694 VTAIL.n672 171.744
R465 VTAIL.n687 VTAIL.n672 171.744
R466 VTAIL.n687 VTAIL.n686 171.744
R467 VTAIL.n686 VTAIL.n676 171.744
R468 VTAIL.n679 VTAIL.n676 171.744
R469 VTAIL.n636 VTAIL.n635 171.744
R470 VTAIL.n635 VTAIL.n539 171.744
R471 VTAIL.n628 VTAIL.n539 171.744
R472 VTAIL.n628 VTAIL.n627 171.744
R473 VTAIL.n627 VTAIL.n543 171.744
R474 VTAIL.n620 VTAIL.n543 171.744
R475 VTAIL.n620 VTAIL.n619 171.744
R476 VTAIL.n619 VTAIL.n547 171.744
R477 VTAIL.n551 VTAIL.n547 171.744
R478 VTAIL.n611 VTAIL.n551 171.744
R479 VTAIL.n611 VTAIL.n610 171.744
R480 VTAIL.n610 VTAIL.n552 171.744
R481 VTAIL.n603 VTAIL.n552 171.744
R482 VTAIL.n603 VTAIL.n602 171.744
R483 VTAIL.n602 VTAIL.n556 171.744
R484 VTAIL.n595 VTAIL.n556 171.744
R485 VTAIL.n595 VTAIL.n594 171.744
R486 VTAIL.n594 VTAIL.n560 171.744
R487 VTAIL.n587 VTAIL.n560 171.744
R488 VTAIL.n587 VTAIL.n586 171.744
R489 VTAIL.n586 VTAIL.n564 171.744
R490 VTAIL.n579 VTAIL.n564 171.744
R491 VTAIL.n579 VTAIL.n578 171.744
R492 VTAIL.n578 VTAIL.n568 171.744
R493 VTAIL.n571 VTAIL.n568 171.744
R494 VTAIL.n530 VTAIL.n529 171.744
R495 VTAIL.n529 VTAIL.n433 171.744
R496 VTAIL.n522 VTAIL.n433 171.744
R497 VTAIL.n522 VTAIL.n521 171.744
R498 VTAIL.n521 VTAIL.n437 171.744
R499 VTAIL.n514 VTAIL.n437 171.744
R500 VTAIL.n514 VTAIL.n513 171.744
R501 VTAIL.n513 VTAIL.n441 171.744
R502 VTAIL.n445 VTAIL.n441 171.744
R503 VTAIL.n505 VTAIL.n445 171.744
R504 VTAIL.n505 VTAIL.n504 171.744
R505 VTAIL.n504 VTAIL.n446 171.744
R506 VTAIL.n497 VTAIL.n446 171.744
R507 VTAIL.n497 VTAIL.n496 171.744
R508 VTAIL.n496 VTAIL.n450 171.744
R509 VTAIL.n489 VTAIL.n450 171.744
R510 VTAIL.n489 VTAIL.n488 171.744
R511 VTAIL.n488 VTAIL.n454 171.744
R512 VTAIL.n481 VTAIL.n454 171.744
R513 VTAIL.n481 VTAIL.n480 171.744
R514 VTAIL.n480 VTAIL.n458 171.744
R515 VTAIL.n473 VTAIL.n458 171.744
R516 VTAIL.n473 VTAIL.n472 171.744
R517 VTAIL.n472 VTAIL.n462 171.744
R518 VTAIL.n465 VTAIL.n462 171.744
R519 VTAIL.n422 VTAIL.n421 171.744
R520 VTAIL.n421 VTAIL.n325 171.744
R521 VTAIL.n414 VTAIL.n325 171.744
R522 VTAIL.n414 VTAIL.n413 171.744
R523 VTAIL.n413 VTAIL.n329 171.744
R524 VTAIL.n406 VTAIL.n329 171.744
R525 VTAIL.n406 VTAIL.n405 171.744
R526 VTAIL.n405 VTAIL.n333 171.744
R527 VTAIL.n337 VTAIL.n333 171.744
R528 VTAIL.n397 VTAIL.n337 171.744
R529 VTAIL.n397 VTAIL.n396 171.744
R530 VTAIL.n396 VTAIL.n338 171.744
R531 VTAIL.n389 VTAIL.n338 171.744
R532 VTAIL.n389 VTAIL.n388 171.744
R533 VTAIL.n388 VTAIL.n342 171.744
R534 VTAIL.n381 VTAIL.n342 171.744
R535 VTAIL.n381 VTAIL.n380 171.744
R536 VTAIL.n380 VTAIL.n346 171.744
R537 VTAIL.n373 VTAIL.n346 171.744
R538 VTAIL.n373 VTAIL.n372 171.744
R539 VTAIL.n372 VTAIL.n350 171.744
R540 VTAIL.n365 VTAIL.n350 171.744
R541 VTAIL.n365 VTAIL.n364 171.744
R542 VTAIL.n364 VTAIL.n354 171.744
R543 VTAIL.n357 VTAIL.n354 171.744
R544 VTAIL.n784 VTAIL.t0 85.8723
R545 VTAIL.n36 VTAIL.t5 85.8723
R546 VTAIL.n142 VTAIL.t8 85.8723
R547 VTAIL.n250 VTAIL.t11 85.8723
R548 VTAIL.n679 VTAIL.t14 85.8723
R549 VTAIL.n571 VTAIL.t13 85.8723
R550 VTAIL.n465 VTAIL.t4 85.8723
R551 VTAIL.n357 VTAIL.t6 85.8723
R552 VTAIL.n1 VTAIL.n0 53.0637
R553 VTAIL.n215 VTAIL.n214 53.0637
R554 VTAIL.n643 VTAIL.n642 53.0637
R555 VTAIL.n429 VTAIL.n428 53.0637
R556 VTAIL.n855 VTAIL.n854 33.5429
R557 VTAIL.n107 VTAIL.n106 33.5429
R558 VTAIL.n213 VTAIL.n212 33.5429
R559 VTAIL.n321 VTAIL.n320 33.5429
R560 VTAIL.n749 VTAIL.n748 33.5429
R561 VTAIL.n641 VTAIL.n640 33.5429
R562 VTAIL.n535 VTAIL.n534 33.5429
R563 VTAIL.n427 VTAIL.n426 33.5429
R564 VTAIL.n855 VTAIL.n749 31.5479
R565 VTAIL.n427 VTAIL.n321 31.5479
R566 VTAIL.n785 VTAIL.n783 16.3895
R567 VTAIL.n37 VTAIL.n35 16.3895
R568 VTAIL.n143 VTAIL.n141 16.3895
R569 VTAIL.n251 VTAIL.n249 16.3895
R570 VTAIL.n680 VTAIL.n678 16.3895
R571 VTAIL.n572 VTAIL.n570 16.3895
R572 VTAIL.n466 VTAIL.n464 16.3895
R573 VTAIL.n358 VTAIL.n356 16.3895
R574 VTAIL.n832 VTAIL.n831 13.1884
R575 VTAIL.n84 VTAIL.n83 13.1884
R576 VTAIL.n190 VTAIL.n189 13.1884
R577 VTAIL.n298 VTAIL.n297 13.1884
R578 VTAIL.n726 VTAIL.n725 13.1884
R579 VTAIL.n618 VTAIL.n617 13.1884
R580 VTAIL.n512 VTAIL.n511 13.1884
R581 VTAIL.n404 VTAIL.n403 13.1884
R582 VTAIL.n786 VTAIL.n782 12.8005
R583 VTAIL.n830 VTAIL.n762 12.8005
R584 VTAIL.n835 VTAIL.n760 12.8005
R585 VTAIL.n38 VTAIL.n34 12.8005
R586 VTAIL.n82 VTAIL.n14 12.8005
R587 VTAIL.n87 VTAIL.n12 12.8005
R588 VTAIL.n144 VTAIL.n140 12.8005
R589 VTAIL.n188 VTAIL.n120 12.8005
R590 VTAIL.n193 VTAIL.n118 12.8005
R591 VTAIL.n252 VTAIL.n248 12.8005
R592 VTAIL.n296 VTAIL.n228 12.8005
R593 VTAIL.n301 VTAIL.n226 12.8005
R594 VTAIL.n729 VTAIL.n654 12.8005
R595 VTAIL.n724 VTAIL.n656 12.8005
R596 VTAIL.n681 VTAIL.n677 12.8005
R597 VTAIL.n621 VTAIL.n546 12.8005
R598 VTAIL.n616 VTAIL.n548 12.8005
R599 VTAIL.n573 VTAIL.n569 12.8005
R600 VTAIL.n515 VTAIL.n440 12.8005
R601 VTAIL.n510 VTAIL.n442 12.8005
R602 VTAIL.n467 VTAIL.n463 12.8005
R603 VTAIL.n407 VTAIL.n332 12.8005
R604 VTAIL.n402 VTAIL.n334 12.8005
R605 VTAIL.n359 VTAIL.n355 12.8005
R606 VTAIL.n790 VTAIL.n789 12.0247
R607 VTAIL.n827 VTAIL.n826 12.0247
R608 VTAIL.n836 VTAIL.n758 12.0247
R609 VTAIL.n42 VTAIL.n41 12.0247
R610 VTAIL.n79 VTAIL.n78 12.0247
R611 VTAIL.n88 VTAIL.n10 12.0247
R612 VTAIL.n148 VTAIL.n147 12.0247
R613 VTAIL.n185 VTAIL.n184 12.0247
R614 VTAIL.n194 VTAIL.n116 12.0247
R615 VTAIL.n256 VTAIL.n255 12.0247
R616 VTAIL.n293 VTAIL.n292 12.0247
R617 VTAIL.n302 VTAIL.n224 12.0247
R618 VTAIL.n730 VTAIL.n652 12.0247
R619 VTAIL.n721 VTAIL.n720 12.0247
R620 VTAIL.n685 VTAIL.n684 12.0247
R621 VTAIL.n622 VTAIL.n544 12.0247
R622 VTAIL.n613 VTAIL.n612 12.0247
R623 VTAIL.n577 VTAIL.n576 12.0247
R624 VTAIL.n516 VTAIL.n438 12.0247
R625 VTAIL.n507 VTAIL.n506 12.0247
R626 VTAIL.n471 VTAIL.n470 12.0247
R627 VTAIL.n408 VTAIL.n330 12.0247
R628 VTAIL.n399 VTAIL.n398 12.0247
R629 VTAIL.n363 VTAIL.n362 12.0247
R630 VTAIL.n793 VTAIL.n780 11.249
R631 VTAIL.n822 VTAIL.n764 11.249
R632 VTAIL.n840 VTAIL.n839 11.249
R633 VTAIL.n45 VTAIL.n32 11.249
R634 VTAIL.n74 VTAIL.n16 11.249
R635 VTAIL.n92 VTAIL.n91 11.249
R636 VTAIL.n151 VTAIL.n138 11.249
R637 VTAIL.n180 VTAIL.n122 11.249
R638 VTAIL.n198 VTAIL.n197 11.249
R639 VTAIL.n259 VTAIL.n246 11.249
R640 VTAIL.n288 VTAIL.n230 11.249
R641 VTAIL.n306 VTAIL.n305 11.249
R642 VTAIL.n734 VTAIL.n733 11.249
R643 VTAIL.n717 VTAIL.n658 11.249
R644 VTAIL.n688 VTAIL.n675 11.249
R645 VTAIL.n626 VTAIL.n625 11.249
R646 VTAIL.n609 VTAIL.n550 11.249
R647 VTAIL.n580 VTAIL.n567 11.249
R648 VTAIL.n520 VTAIL.n519 11.249
R649 VTAIL.n503 VTAIL.n444 11.249
R650 VTAIL.n474 VTAIL.n461 11.249
R651 VTAIL.n412 VTAIL.n411 11.249
R652 VTAIL.n395 VTAIL.n336 11.249
R653 VTAIL.n366 VTAIL.n353 11.249
R654 VTAIL.n794 VTAIL.n778 10.4732
R655 VTAIL.n821 VTAIL.n766 10.4732
R656 VTAIL.n843 VTAIL.n756 10.4732
R657 VTAIL.n46 VTAIL.n30 10.4732
R658 VTAIL.n73 VTAIL.n18 10.4732
R659 VTAIL.n95 VTAIL.n8 10.4732
R660 VTAIL.n152 VTAIL.n136 10.4732
R661 VTAIL.n179 VTAIL.n124 10.4732
R662 VTAIL.n201 VTAIL.n114 10.4732
R663 VTAIL.n260 VTAIL.n244 10.4732
R664 VTAIL.n287 VTAIL.n232 10.4732
R665 VTAIL.n309 VTAIL.n222 10.4732
R666 VTAIL.n737 VTAIL.n650 10.4732
R667 VTAIL.n716 VTAIL.n661 10.4732
R668 VTAIL.n689 VTAIL.n673 10.4732
R669 VTAIL.n629 VTAIL.n542 10.4732
R670 VTAIL.n608 VTAIL.n553 10.4732
R671 VTAIL.n581 VTAIL.n565 10.4732
R672 VTAIL.n523 VTAIL.n436 10.4732
R673 VTAIL.n502 VTAIL.n447 10.4732
R674 VTAIL.n475 VTAIL.n459 10.4732
R675 VTAIL.n415 VTAIL.n328 10.4732
R676 VTAIL.n394 VTAIL.n339 10.4732
R677 VTAIL.n367 VTAIL.n351 10.4732
R678 VTAIL.n798 VTAIL.n797 9.69747
R679 VTAIL.n818 VTAIL.n817 9.69747
R680 VTAIL.n844 VTAIL.n754 9.69747
R681 VTAIL.n50 VTAIL.n49 9.69747
R682 VTAIL.n70 VTAIL.n69 9.69747
R683 VTAIL.n96 VTAIL.n6 9.69747
R684 VTAIL.n156 VTAIL.n155 9.69747
R685 VTAIL.n176 VTAIL.n175 9.69747
R686 VTAIL.n202 VTAIL.n112 9.69747
R687 VTAIL.n264 VTAIL.n263 9.69747
R688 VTAIL.n284 VTAIL.n283 9.69747
R689 VTAIL.n310 VTAIL.n220 9.69747
R690 VTAIL.n738 VTAIL.n648 9.69747
R691 VTAIL.n713 VTAIL.n712 9.69747
R692 VTAIL.n693 VTAIL.n692 9.69747
R693 VTAIL.n630 VTAIL.n540 9.69747
R694 VTAIL.n605 VTAIL.n604 9.69747
R695 VTAIL.n585 VTAIL.n584 9.69747
R696 VTAIL.n524 VTAIL.n434 9.69747
R697 VTAIL.n499 VTAIL.n498 9.69747
R698 VTAIL.n479 VTAIL.n478 9.69747
R699 VTAIL.n416 VTAIL.n326 9.69747
R700 VTAIL.n391 VTAIL.n390 9.69747
R701 VTAIL.n371 VTAIL.n370 9.69747
R702 VTAIL.n854 VTAIL.n853 9.45567
R703 VTAIL.n106 VTAIL.n105 9.45567
R704 VTAIL.n212 VTAIL.n211 9.45567
R705 VTAIL.n320 VTAIL.n319 9.45567
R706 VTAIL.n748 VTAIL.n747 9.45567
R707 VTAIL.n640 VTAIL.n639 9.45567
R708 VTAIL.n534 VTAIL.n533 9.45567
R709 VTAIL.n426 VTAIL.n425 9.45567
R710 VTAIL.n752 VTAIL.n751 9.3005
R711 VTAIL.n847 VTAIL.n846 9.3005
R712 VTAIL.n845 VTAIL.n844 9.3005
R713 VTAIL.n756 VTAIL.n755 9.3005
R714 VTAIL.n839 VTAIL.n838 9.3005
R715 VTAIL.n837 VTAIL.n836 9.3005
R716 VTAIL.n760 VTAIL.n759 9.3005
R717 VTAIL.n805 VTAIL.n804 9.3005
R718 VTAIL.n803 VTAIL.n802 9.3005
R719 VTAIL.n776 VTAIL.n775 9.3005
R720 VTAIL.n797 VTAIL.n796 9.3005
R721 VTAIL.n795 VTAIL.n794 9.3005
R722 VTAIL.n780 VTAIL.n779 9.3005
R723 VTAIL.n789 VTAIL.n788 9.3005
R724 VTAIL.n787 VTAIL.n786 9.3005
R725 VTAIL.n772 VTAIL.n771 9.3005
R726 VTAIL.n811 VTAIL.n810 9.3005
R727 VTAIL.n813 VTAIL.n812 9.3005
R728 VTAIL.n768 VTAIL.n767 9.3005
R729 VTAIL.n819 VTAIL.n818 9.3005
R730 VTAIL.n821 VTAIL.n820 9.3005
R731 VTAIL.n764 VTAIL.n763 9.3005
R732 VTAIL.n828 VTAIL.n827 9.3005
R733 VTAIL.n830 VTAIL.n829 9.3005
R734 VTAIL.n853 VTAIL.n852 9.3005
R735 VTAIL.n4 VTAIL.n3 9.3005
R736 VTAIL.n99 VTAIL.n98 9.3005
R737 VTAIL.n97 VTAIL.n96 9.3005
R738 VTAIL.n8 VTAIL.n7 9.3005
R739 VTAIL.n91 VTAIL.n90 9.3005
R740 VTAIL.n89 VTAIL.n88 9.3005
R741 VTAIL.n12 VTAIL.n11 9.3005
R742 VTAIL.n57 VTAIL.n56 9.3005
R743 VTAIL.n55 VTAIL.n54 9.3005
R744 VTAIL.n28 VTAIL.n27 9.3005
R745 VTAIL.n49 VTAIL.n48 9.3005
R746 VTAIL.n47 VTAIL.n46 9.3005
R747 VTAIL.n32 VTAIL.n31 9.3005
R748 VTAIL.n41 VTAIL.n40 9.3005
R749 VTAIL.n39 VTAIL.n38 9.3005
R750 VTAIL.n24 VTAIL.n23 9.3005
R751 VTAIL.n63 VTAIL.n62 9.3005
R752 VTAIL.n65 VTAIL.n64 9.3005
R753 VTAIL.n20 VTAIL.n19 9.3005
R754 VTAIL.n71 VTAIL.n70 9.3005
R755 VTAIL.n73 VTAIL.n72 9.3005
R756 VTAIL.n16 VTAIL.n15 9.3005
R757 VTAIL.n80 VTAIL.n79 9.3005
R758 VTAIL.n82 VTAIL.n81 9.3005
R759 VTAIL.n105 VTAIL.n104 9.3005
R760 VTAIL.n110 VTAIL.n109 9.3005
R761 VTAIL.n205 VTAIL.n204 9.3005
R762 VTAIL.n203 VTAIL.n202 9.3005
R763 VTAIL.n114 VTAIL.n113 9.3005
R764 VTAIL.n197 VTAIL.n196 9.3005
R765 VTAIL.n195 VTAIL.n194 9.3005
R766 VTAIL.n118 VTAIL.n117 9.3005
R767 VTAIL.n163 VTAIL.n162 9.3005
R768 VTAIL.n161 VTAIL.n160 9.3005
R769 VTAIL.n134 VTAIL.n133 9.3005
R770 VTAIL.n155 VTAIL.n154 9.3005
R771 VTAIL.n153 VTAIL.n152 9.3005
R772 VTAIL.n138 VTAIL.n137 9.3005
R773 VTAIL.n147 VTAIL.n146 9.3005
R774 VTAIL.n145 VTAIL.n144 9.3005
R775 VTAIL.n130 VTAIL.n129 9.3005
R776 VTAIL.n169 VTAIL.n168 9.3005
R777 VTAIL.n171 VTAIL.n170 9.3005
R778 VTAIL.n126 VTAIL.n125 9.3005
R779 VTAIL.n177 VTAIL.n176 9.3005
R780 VTAIL.n179 VTAIL.n178 9.3005
R781 VTAIL.n122 VTAIL.n121 9.3005
R782 VTAIL.n186 VTAIL.n185 9.3005
R783 VTAIL.n188 VTAIL.n187 9.3005
R784 VTAIL.n211 VTAIL.n210 9.3005
R785 VTAIL.n218 VTAIL.n217 9.3005
R786 VTAIL.n313 VTAIL.n312 9.3005
R787 VTAIL.n311 VTAIL.n310 9.3005
R788 VTAIL.n222 VTAIL.n221 9.3005
R789 VTAIL.n305 VTAIL.n304 9.3005
R790 VTAIL.n303 VTAIL.n302 9.3005
R791 VTAIL.n226 VTAIL.n225 9.3005
R792 VTAIL.n271 VTAIL.n270 9.3005
R793 VTAIL.n269 VTAIL.n268 9.3005
R794 VTAIL.n242 VTAIL.n241 9.3005
R795 VTAIL.n263 VTAIL.n262 9.3005
R796 VTAIL.n261 VTAIL.n260 9.3005
R797 VTAIL.n246 VTAIL.n245 9.3005
R798 VTAIL.n255 VTAIL.n254 9.3005
R799 VTAIL.n253 VTAIL.n252 9.3005
R800 VTAIL.n238 VTAIL.n237 9.3005
R801 VTAIL.n277 VTAIL.n276 9.3005
R802 VTAIL.n279 VTAIL.n278 9.3005
R803 VTAIL.n234 VTAIL.n233 9.3005
R804 VTAIL.n285 VTAIL.n284 9.3005
R805 VTAIL.n287 VTAIL.n286 9.3005
R806 VTAIL.n230 VTAIL.n229 9.3005
R807 VTAIL.n294 VTAIL.n293 9.3005
R808 VTAIL.n296 VTAIL.n295 9.3005
R809 VTAIL.n319 VTAIL.n318 9.3005
R810 VTAIL.n706 VTAIL.n705 9.3005
R811 VTAIL.n708 VTAIL.n707 9.3005
R812 VTAIL.n663 VTAIL.n662 9.3005
R813 VTAIL.n714 VTAIL.n713 9.3005
R814 VTAIL.n716 VTAIL.n715 9.3005
R815 VTAIL.n658 VTAIL.n657 9.3005
R816 VTAIL.n722 VTAIL.n721 9.3005
R817 VTAIL.n724 VTAIL.n723 9.3005
R818 VTAIL.n747 VTAIL.n746 9.3005
R819 VTAIL.n646 VTAIL.n645 9.3005
R820 VTAIL.n741 VTAIL.n740 9.3005
R821 VTAIL.n739 VTAIL.n738 9.3005
R822 VTAIL.n650 VTAIL.n649 9.3005
R823 VTAIL.n733 VTAIL.n732 9.3005
R824 VTAIL.n731 VTAIL.n730 9.3005
R825 VTAIL.n654 VTAIL.n653 9.3005
R826 VTAIL.n667 VTAIL.n666 9.3005
R827 VTAIL.n700 VTAIL.n699 9.3005
R828 VTAIL.n698 VTAIL.n697 9.3005
R829 VTAIL.n671 VTAIL.n670 9.3005
R830 VTAIL.n692 VTAIL.n691 9.3005
R831 VTAIL.n690 VTAIL.n689 9.3005
R832 VTAIL.n675 VTAIL.n674 9.3005
R833 VTAIL.n684 VTAIL.n683 9.3005
R834 VTAIL.n682 VTAIL.n681 9.3005
R835 VTAIL.n598 VTAIL.n597 9.3005
R836 VTAIL.n600 VTAIL.n599 9.3005
R837 VTAIL.n555 VTAIL.n554 9.3005
R838 VTAIL.n606 VTAIL.n605 9.3005
R839 VTAIL.n608 VTAIL.n607 9.3005
R840 VTAIL.n550 VTAIL.n549 9.3005
R841 VTAIL.n614 VTAIL.n613 9.3005
R842 VTAIL.n616 VTAIL.n615 9.3005
R843 VTAIL.n639 VTAIL.n638 9.3005
R844 VTAIL.n538 VTAIL.n537 9.3005
R845 VTAIL.n633 VTAIL.n632 9.3005
R846 VTAIL.n631 VTAIL.n630 9.3005
R847 VTAIL.n542 VTAIL.n541 9.3005
R848 VTAIL.n625 VTAIL.n624 9.3005
R849 VTAIL.n623 VTAIL.n622 9.3005
R850 VTAIL.n546 VTAIL.n545 9.3005
R851 VTAIL.n559 VTAIL.n558 9.3005
R852 VTAIL.n592 VTAIL.n591 9.3005
R853 VTAIL.n590 VTAIL.n589 9.3005
R854 VTAIL.n563 VTAIL.n562 9.3005
R855 VTAIL.n584 VTAIL.n583 9.3005
R856 VTAIL.n582 VTAIL.n581 9.3005
R857 VTAIL.n567 VTAIL.n566 9.3005
R858 VTAIL.n576 VTAIL.n575 9.3005
R859 VTAIL.n574 VTAIL.n573 9.3005
R860 VTAIL.n492 VTAIL.n491 9.3005
R861 VTAIL.n494 VTAIL.n493 9.3005
R862 VTAIL.n449 VTAIL.n448 9.3005
R863 VTAIL.n500 VTAIL.n499 9.3005
R864 VTAIL.n502 VTAIL.n501 9.3005
R865 VTAIL.n444 VTAIL.n443 9.3005
R866 VTAIL.n508 VTAIL.n507 9.3005
R867 VTAIL.n510 VTAIL.n509 9.3005
R868 VTAIL.n533 VTAIL.n532 9.3005
R869 VTAIL.n432 VTAIL.n431 9.3005
R870 VTAIL.n527 VTAIL.n526 9.3005
R871 VTAIL.n525 VTAIL.n524 9.3005
R872 VTAIL.n436 VTAIL.n435 9.3005
R873 VTAIL.n519 VTAIL.n518 9.3005
R874 VTAIL.n517 VTAIL.n516 9.3005
R875 VTAIL.n440 VTAIL.n439 9.3005
R876 VTAIL.n453 VTAIL.n452 9.3005
R877 VTAIL.n486 VTAIL.n485 9.3005
R878 VTAIL.n484 VTAIL.n483 9.3005
R879 VTAIL.n457 VTAIL.n456 9.3005
R880 VTAIL.n478 VTAIL.n477 9.3005
R881 VTAIL.n476 VTAIL.n475 9.3005
R882 VTAIL.n461 VTAIL.n460 9.3005
R883 VTAIL.n470 VTAIL.n469 9.3005
R884 VTAIL.n468 VTAIL.n467 9.3005
R885 VTAIL.n384 VTAIL.n383 9.3005
R886 VTAIL.n386 VTAIL.n385 9.3005
R887 VTAIL.n341 VTAIL.n340 9.3005
R888 VTAIL.n392 VTAIL.n391 9.3005
R889 VTAIL.n394 VTAIL.n393 9.3005
R890 VTAIL.n336 VTAIL.n335 9.3005
R891 VTAIL.n400 VTAIL.n399 9.3005
R892 VTAIL.n402 VTAIL.n401 9.3005
R893 VTAIL.n425 VTAIL.n424 9.3005
R894 VTAIL.n324 VTAIL.n323 9.3005
R895 VTAIL.n419 VTAIL.n418 9.3005
R896 VTAIL.n417 VTAIL.n416 9.3005
R897 VTAIL.n328 VTAIL.n327 9.3005
R898 VTAIL.n411 VTAIL.n410 9.3005
R899 VTAIL.n409 VTAIL.n408 9.3005
R900 VTAIL.n332 VTAIL.n331 9.3005
R901 VTAIL.n345 VTAIL.n344 9.3005
R902 VTAIL.n378 VTAIL.n377 9.3005
R903 VTAIL.n376 VTAIL.n375 9.3005
R904 VTAIL.n349 VTAIL.n348 9.3005
R905 VTAIL.n370 VTAIL.n369 9.3005
R906 VTAIL.n368 VTAIL.n367 9.3005
R907 VTAIL.n353 VTAIL.n352 9.3005
R908 VTAIL.n362 VTAIL.n361 9.3005
R909 VTAIL.n360 VTAIL.n359 9.3005
R910 VTAIL.n801 VTAIL.n776 8.92171
R911 VTAIL.n814 VTAIL.n768 8.92171
R912 VTAIL.n848 VTAIL.n847 8.92171
R913 VTAIL.n53 VTAIL.n28 8.92171
R914 VTAIL.n66 VTAIL.n20 8.92171
R915 VTAIL.n100 VTAIL.n99 8.92171
R916 VTAIL.n159 VTAIL.n134 8.92171
R917 VTAIL.n172 VTAIL.n126 8.92171
R918 VTAIL.n206 VTAIL.n205 8.92171
R919 VTAIL.n267 VTAIL.n242 8.92171
R920 VTAIL.n280 VTAIL.n234 8.92171
R921 VTAIL.n314 VTAIL.n313 8.92171
R922 VTAIL.n742 VTAIL.n741 8.92171
R923 VTAIL.n709 VTAIL.n663 8.92171
R924 VTAIL.n696 VTAIL.n671 8.92171
R925 VTAIL.n634 VTAIL.n633 8.92171
R926 VTAIL.n601 VTAIL.n555 8.92171
R927 VTAIL.n588 VTAIL.n563 8.92171
R928 VTAIL.n528 VTAIL.n527 8.92171
R929 VTAIL.n495 VTAIL.n449 8.92171
R930 VTAIL.n482 VTAIL.n457 8.92171
R931 VTAIL.n420 VTAIL.n419 8.92171
R932 VTAIL.n387 VTAIL.n341 8.92171
R933 VTAIL.n374 VTAIL.n349 8.92171
R934 VTAIL.n802 VTAIL.n774 8.14595
R935 VTAIL.n813 VTAIL.n770 8.14595
R936 VTAIL.n851 VTAIL.n752 8.14595
R937 VTAIL.n54 VTAIL.n26 8.14595
R938 VTAIL.n65 VTAIL.n22 8.14595
R939 VTAIL.n103 VTAIL.n4 8.14595
R940 VTAIL.n160 VTAIL.n132 8.14595
R941 VTAIL.n171 VTAIL.n128 8.14595
R942 VTAIL.n209 VTAIL.n110 8.14595
R943 VTAIL.n268 VTAIL.n240 8.14595
R944 VTAIL.n279 VTAIL.n236 8.14595
R945 VTAIL.n317 VTAIL.n218 8.14595
R946 VTAIL.n745 VTAIL.n646 8.14595
R947 VTAIL.n708 VTAIL.n665 8.14595
R948 VTAIL.n697 VTAIL.n669 8.14595
R949 VTAIL.n637 VTAIL.n538 8.14595
R950 VTAIL.n600 VTAIL.n557 8.14595
R951 VTAIL.n589 VTAIL.n561 8.14595
R952 VTAIL.n531 VTAIL.n432 8.14595
R953 VTAIL.n494 VTAIL.n451 8.14595
R954 VTAIL.n483 VTAIL.n455 8.14595
R955 VTAIL.n423 VTAIL.n324 8.14595
R956 VTAIL.n386 VTAIL.n343 8.14595
R957 VTAIL.n375 VTAIL.n347 8.14595
R958 VTAIL.n806 VTAIL.n805 7.3702
R959 VTAIL.n810 VTAIL.n809 7.3702
R960 VTAIL.n852 VTAIL.n750 7.3702
R961 VTAIL.n58 VTAIL.n57 7.3702
R962 VTAIL.n62 VTAIL.n61 7.3702
R963 VTAIL.n104 VTAIL.n2 7.3702
R964 VTAIL.n164 VTAIL.n163 7.3702
R965 VTAIL.n168 VTAIL.n167 7.3702
R966 VTAIL.n210 VTAIL.n108 7.3702
R967 VTAIL.n272 VTAIL.n271 7.3702
R968 VTAIL.n276 VTAIL.n275 7.3702
R969 VTAIL.n318 VTAIL.n216 7.3702
R970 VTAIL.n746 VTAIL.n644 7.3702
R971 VTAIL.n705 VTAIL.n704 7.3702
R972 VTAIL.n701 VTAIL.n700 7.3702
R973 VTAIL.n638 VTAIL.n536 7.3702
R974 VTAIL.n597 VTAIL.n596 7.3702
R975 VTAIL.n593 VTAIL.n592 7.3702
R976 VTAIL.n532 VTAIL.n430 7.3702
R977 VTAIL.n491 VTAIL.n490 7.3702
R978 VTAIL.n487 VTAIL.n486 7.3702
R979 VTAIL.n424 VTAIL.n322 7.3702
R980 VTAIL.n383 VTAIL.n382 7.3702
R981 VTAIL.n379 VTAIL.n378 7.3702
R982 VTAIL.n806 VTAIL.n772 6.59444
R983 VTAIL.n809 VTAIL.n772 6.59444
R984 VTAIL.n854 VTAIL.n750 6.59444
R985 VTAIL.n58 VTAIL.n24 6.59444
R986 VTAIL.n61 VTAIL.n24 6.59444
R987 VTAIL.n106 VTAIL.n2 6.59444
R988 VTAIL.n164 VTAIL.n130 6.59444
R989 VTAIL.n167 VTAIL.n130 6.59444
R990 VTAIL.n212 VTAIL.n108 6.59444
R991 VTAIL.n272 VTAIL.n238 6.59444
R992 VTAIL.n275 VTAIL.n238 6.59444
R993 VTAIL.n320 VTAIL.n216 6.59444
R994 VTAIL.n748 VTAIL.n644 6.59444
R995 VTAIL.n704 VTAIL.n667 6.59444
R996 VTAIL.n701 VTAIL.n667 6.59444
R997 VTAIL.n640 VTAIL.n536 6.59444
R998 VTAIL.n596 VTAIL.n559 6.59444
R999 VTAIL.n593 VTAIL.n559 6.59444
R1000 VTAIL.n534 VTAIL.n430 6.59444
R1001 VTAIL.n490 VTAIL.n453 6.59444
R1002 VTAIL.n487 VTAIL.n453 6.59444
R1003 VTAIL.n426 VTAIL.n322 6.59444
R1004 VTAIL.n382 VTAIL.n345 6.59444
R1005 VTAIL.n379 VTAIL.n345 6.59444
R1006 VTAIL.n805 VTAIL.n774 5.81868
R1007 VTAIL.n810 VTAIL.n770 5.81868
R1008 VTAIL.n852 VTAIL.n851 5.81868
R1009 VTAIL.n57 VTAIL.n26 5.81868
R1010 VTAIL.n62 VTAIL.n22 5.81868
R1011 VTAIL.n104 VTAIL.n103 5.81868
R1012 VTAIL.n163 VTAIL.n132 5.81868
R1013 VTAIL.n168 VTAIL.n128 5.81868
R1014 VTAIL.n210 VTAIL.n209 5.81868
R1015 VTAIL.n271 VTAIL.n240 5.81868
R1016 VTAIL.n276 VTAIL.n236 5.81868
R1017 VTAIL.n318 VTAIL.n317 5.81868
R1018 VTAIL.n746 VTAIL.n745 5.81868
R1019 VTAIL.n705 VTAIL.n665 5.81868
R1020 VTAIL.n700 VTAIL.n669 5.81868
R1021 VTAIL.n638 VTAIL.n637 5.81868
R1022 VTAIL.n597 VTAIL.n557 5.81868
R1023 VTAIL.n592 VTAIL.n561 5.81868
R1024 VTAIL.n532 VTAIL.n531 5.81868
R1025 VTAIL.n491 VTAIL.n451 5.81868
R1026 VTAIL.n486 VTAIL.n455 5.81868
R1027 VTAIL.n424 VTAIL.n423 5.81868
R1028 VTAIL.n383 VTAIL.n343 5.81868
R1029 VTAIL.n378 VTAIL.n347 5.81868
R1030 VTAIL.n802 VTAIL.n801 5.04292
R1031 VTAIL.n814 VTAIL.n813 5.04292
R1032 VTAIL.n848 VTAIL.n752 5.04292
R1033 VTAIL.n54 VTAIL.n53 5.04292
R1034 VTAIL.n66 VTAIL.n65 5.04292
R1035 VTAIL.n100 VTAIL.n4 5.04292
R1036 VTAIL.n160 VTAIL.n159 5.04292
R1037 VTAIL.n172 VTAIL.n171 5.04292
R1038 VTAIL.n206 VTAIL.n110 5.04292
R1039 VTAIL.n268 VTAIL.n267 5.04292
R1040 VTAIL.n280 VTAIL.n279 5.04292
R1041 VTAIL.n314 VTAIL.n218 5.04292
R1042 VTAIL.n742 VTAIL.n646 5.04292
R1043 VTAIL.n709 VTAIL.n708 5.04292
R1044 VTAIL.n697 VTAIL.n696 5.04292
R1045 VTAIL.n634 VTAIL.n538 5.04292
R1046 VTAIL.n601 VTAIL.n600 5.04292
R1047 VTAIL.n589 VTAIL.n588 5.04292
R1048 VTAIL.n528 VTAIL.n432 5.04292
R1049 VTAIL.n495 VTAIL.n494 5.04292
R1050 VTAIL.n483 VTAIL.n482 5.04292
R1051 VTAIL.n420 VTAIL.n324 5.04292
R1052 VTAIL.n387 VTAIL.n386 5.04292
R1053 VTAIL.n375 VTAIL.n374 5.04292
R1054 VTAIL.n798 VTAIL.n776 4.26717
R1055 VTAIL.n817 VTAIL.n768 4.26717
R1056 VTAIL.n847 VTAIL.n754 4.26717
R1057 VTAIL.n50 VTAIL.n28 4.26717
R1058 VTAIL.n69 VTAIL.n20 4.26717
R1059 VTAIL.n99 VTAIL.n6 4.26717
R1060 VTAIL.n156 VTAIL.n134 4.26717
R1061 VTAIL.n175 VTAIL.n126 4.26717
R1062 VTAIL.n205 VTAIL.n112 4.26717
R1063 VTAIL.n264 VTAIL.n242 4.26717
R1064 VTAIL.n283 VTAIL.n234 4.26717
R1065 VTAIL.n313 VTAIL.n220 4.26717
R1066 VTAIL.n741 VTAIL.n648 4.26717
R1067 VTAIL.n712 VTAIL.n663 4.26717
R1068 VTAIL.n693 VTAIL.n671 4.26717
R1069 VTAIL.n633 VTAIL.n540 4.26717
R1070 VTAIL.n604 VTAIL.n555 4.26717
R1071 VTAIL.n585 VTAIL.n563 4.26717
R1072 VTAIL.n527 VTAIL.n434 4.26717
R1073 VTAIL.n498 VTAIL.n449 4.26717
R1074 VTAIL.n479 VTAIL.n457 4.26717
R1075 VTAIL.n419 VTAIL.n326 4.26717
R1076 VTAIL.n390 VTAIL.n341 4.26717
R1077 VTAIL.n371 VTAIL.n349 4.26717
R1078 VTAIL.n787 VTAIL.n783 3.70982
R1079 VTAIL.n39 VTAIL.n35 3.70982
R1080 VTAIL.n145 VTAIL.n141 3.70982
R1081 VTAIL.n253 VTAIL.n249 3.70982
R1082 VTAIL.n682 VTAIL.n678 3.70982
R1083 VTAIL.n574 VTAIL.n570 3.70982
R1084 VTAIL.n468 VTAIL.n464 3.70982
R1085 VTAIL.n360 VTAIL.n356 3.70982
R1086 VTAIL.n797 VTAIL.n778 3.49141
R1087 VTAIL.n818 VTAIL.n766 3.49141
R1088 VTAIL.n844 VTAIL.n843 3.49141
R1089 VTAIL.n49 VTAIL.n30 3.49141
R1090 VTAIL.n70 VTAIL.n18 3.49141
R1091 VTAIL.n96 VTAIL.n95 3.49141
R1092 VTAIL.n155 VTAIL.n136 3.49141
R1093 VTAIL.n176 VTAIL.n124 3.49141
R1094 VTAIL.n202 VTAIL.n201 3.49141
R1095 VTAIL.n263 VTAIL.n244 3.49141
R1096 VTAIL.n284 VTAIL.n232 3.49141
R1097 VTAIL.n310 VTAIL.n309 3.49141
R1098 VTAIL.n738 VTAIL.n737 3.49141
R1099 VTAIL.n713 VTAIL.n661 3.49141
R1100 VTAIL.n692 VTAIL.n673 3.49141
R1101 VTAIL.n630 VTAIL.n629 3.49141
R1102 VTAIL.n605 VTAIL.n553 3.49141
R1103 VTAIL.n584 VTAIL.n565 3.49141
R1104 VTAIL.n524 VTAIL.n523 3.49141
R1105 VTAIL.n499 VTAIL.n447 3.49141
R1106 VTAIL.n478 VTAIL.n459 3.49141
R1107 VTAIL.n416 VTAIL.n415 3.49141
R1108 VTAIL.n391 VTAIL.n339 3.49141
R1109 VTAIL.n370 VTAIL.n351 3.49141
R1110 VTAIL.n429 VTAIL.n427 2.77636
R1111 VTAIL.n535 VTAIL.n429 2.77636
R1112 VTAIL.n643 VTAIL.n641 2.77636
R1113 VTAIL.n749 VTAIL.n643 2.77636
R1114 VTAIL.n321 VTAIL.n215 2.77636
R1115 VTAIL.n215 VTAIL.n213 2.77636
R1116 VTAIL.n107 VTAIL.n1 2.77636
R1117 VTAIL VTAIL.n855 2.71817
R1118 VTAIL.n794 VTAIL.n793 2.71565
R1119 VTAIL.n822 VTAIL.n821 2.71565
R1120 VTAIL.n840 VTAIL.n756 2.71565
R1121 VTAIL.n46 VTAIL.n45 2.71565
R1122 VTAIL.n74 VTAIL.n73 2.71565
R1123 VTAIL.n92 VTAIL.n8 2.71565
R1124 VTAIL.n152 VTAIL.n151 2.71565
R1125 VTAIL.n180 VTAIL.n179 2.71565
R1126 VTAIL.n198 VTAIL.n114 2.71565
R1127 VTAIL.n260 VTAIL.n259 2.71565
R1128 VTAIL.n288 VTAIL.n287 2.71565
R1129 VTAIL.n306 VTAIL.n222 2.71565
R1130 VTAIL.n734 VTAIL.n650 2.71565
R1131 VTAIL.n717 VTAIL.n716 2.71565
R1132 VTAIL.n689 VTAIL.n688 2.71565
R1133 VTAIL.n626 VTAIL.n542 2.71565
R1134 VTAIL.n609 VTAIL.n608 2.71565
R1135 VTAIL.n581 VTAIL.n580 2.71565
R1136 VTAIL.n520 VTAIL.n436 2.71565
R1137 VTAIL.n503 VTAIL.n502 2.71565
R1138 VTAIL.n475 VTAIL.n474 2.71565
R1139 VTAIL.n412 VTAIL.n328 2.71565
R1140 VTAIL.n395 VTAIL.n394 2.71565
R1141 VTAIL.n367 VTAIL.n366 2.71565
R1142 VTAIL.n790 VTAIL.n780 1.93989
R1143 VTAIL.n826 VTAIL.n764 1.93989
R1144 VTAIL.n839 VTAIL.n758 1.93989
R1145 VTAIL.n42 VTAIL.n32 1.93989
R1146 VTAIL.n78 VTAIL.n16 1.93989
R1147 VTAIL.n91 VTAIL.n10 1.93989
R1148 VTAIL.n148 VTAIL.n138 1.93989
R1149 VTAIL.n184 VTAIL.n122 1.93989
R1150 VTAIL.n197 VTAIL.n116 1.93989
R1151 VTAIL.n256 VTAIL.n246 1.93989
R1152 VTAIL.n292 VTAIL.n230 1.93989
R1153 VTAIL.n305 VTAIL.n224 1.93989
R1154 VTAIL.n733 VTAIL.n652 1.93989
R1155 VTAIL.n720 VTAIL.n658 1.93989
R1156 VTAIL.n685 VTAIL.n675 1.93989
R1157 VTAIL.n625 VTAIL.n544 1.93989
R1158 VTAIL.n612 VTAIL.n550 1.93989
R1159 VTAIL.n577 VTAIL.n567 1.93989
R1160 VTAIL.n519 VTAIL.n438 1.93989
R1161 VTAIL.n506 VTAIL.n444 1.93989
R1162 VTAIL.n471 VTAIL.n461 1.93989
R1163 VTAIL.n411 VTAIL.n330 1.93989
R1164 VTAIL.n398 VTAIL.n336 1.93989
R1165 VTAIL.n363 VTAIL.n353 1.93989
R1166 VTAIL.n0 VTAIL.t2 1.70859
R1167 VTAIL.n0 VTAIL.t7 1.70859
R1168 VTAIL.n214 VTAIL.t12 1.70859
R1169 VTAIL.n214 VTAIL.t15 1.70859
R1170 VTAIL.n642 VTAIL.t10 1.70859
R1171 VTAIL.n642 VTAIL.t9 1.70859
R1172 VTAIL.n428 VTAIL.t1 1.70859
R1173 VTAIL.n428 VTAIL.t3 1.70859
R1174 VTAIL.n789 VTAIL.n782 1.16414
R1175 VTAIL.n827 VTAIL.n762 1.16414
R1176 VTAIL.n836 VTAIL.n835 1.16414
R1177 VTAIL.n41 VTAIL.n34 1.16414
R1178 VTAIL.n79 VTAIL.n14 1.16414
R1179 VTAIL.n88 VTAIL.n87 1.16414
R1180 VTAIL.n147 VTAIL.n140 1.16414
R1181 VTAIL.n185 VTAIL.n120 1.16414
R1182 VTAIL.n194 VTAIL.n193 1.16414
R1183 VTAIL.n255 VTAIL.n248 1.16414
R1184 VTAIL.n293 VTAIL.n228 1.16414
R1185 VTAIL.n302 VTAIL.n301 1.16414
R1186 VTAIL.n730 VTAIL.n729 1.16414
R1187 VTAIL.n721 VTAIL.n656 1.16414
R1188 VTAIL.n684 VTAIL.n677 1.16414
R1189 VTAIL.n622 VTAIL.n621 1.16414
R1190 VTAIL.n613 VTAIL.n548 1.16414
R1191 VTAIL.n576 VTAIL.n569 1.16414
R1192 VTAIL.n516 VTAIL.n515 1.16414
R1193 VTAIL.n507 VTAIL.n442 1.16414
R1194 VTAIL.n470 VTAIL.n463 1.16414
R1195 VTAIL.n408 VTAIL.n407 1.16414
R1196 VTAIL.n399 VTAIL.n334 1.16414
R1197 VTAIL.n362 VTAIL.n355 1.16414
R1198 VTAIL.n641 VTAIL.n535 0.470328
R1199 VTAIL.n213 VTAIL.n107 0.470328
R1200 VTAIL.n786 VTAIL.n785 0.388379
R1201 VTAIL.n831 VTAIL.n830 0.388379
R1202 VTAIL.n832 VTAIL.n760 0.388379
R1203 VTAIL.n38 VTAIL.n37 0.388379
R1204 VTAIL.n83 VTAIL.n82 0.388379
R1205 VTAIL.n84 VTAIL.n12 0.388379
R1206 VTAIL.n144 VTAIL.n143 0.388379
R1207 VTAIL.n189 VTAIL.n188 0.388379
R1208 VTAIL.n190 VTAIL.n118 0.388379
R1209 VTAIL.n252 VTAIL.n251 0.388379
R1210 VTAIL.n297 VTAIL.n296 0.388379
R1211 VTAIL.n298 VTAIL.n226 0.388379
R1212 VTAIL.n726 VTAIL.n654 0.388379
R1213 VTAIL.n725 VTAIL.n724 0.388379
R1214 VTAIL.n681 VTAIL.n680 0.388379
R1215 VTAIL.n618 VTAIL.n546 0.388379
R1216 VTAIL.n617 VTAIL.n616 0.388379
R1217 VTAIL.n573 VTAIL.n572 0.388379
R1218 VTAIL.n512 VTAIL.n440 0.388379
R1219 VTAIL.n511 VTAIL.n510 0.388379
R1220 VTAIL.n467 VTAIL.n466 0.388379
R1221 VTAIL.n404 VTAIL.n332 0.388379
R1222 VTAIL.n403 VTAIL.n402 0.388379
R1223 VTAIL.n359 VTAIL.n358 0.388379
R1224 VTAIL.n788 VTAIL.n787 0.155672
R1225 VTAIL.n788 VTAIL.n779 0.155672
R1226 VTAIL.n795 VTAIL.n779 0.155672
R1227 VTAIL.n796 VTAIL.n795 0.155672
R1228 VTAIL.n796 VTAIL.n775 0.155672
R1229 VTAIL.n803 VTAIL.n775 0.155672
R1230 VTAIL.n804 VTAIL.n803 0.155672
R1231 VTAIL.n804 VTAIL.n771 0.155672
R1232 VTAIL.n811 VTAIL.n771 0.155672
R1233 VTAIL.n812 VTAIL.n811 0.155672
R1234 VTAIL.n812 VTAIL.n767 0.155672
R1235 VTAIL.n819 VTAIL.n767 0.155672
R1236 VTAIL.n820 VTAIL.n819 0.155672
R1237 VTAIL.n820 VTAIL.n763 0.155672
R1238 VTAIL.n828 VTAIL.n763 0.155672
R1239 VTAIL.n829 VTAIL.n828 0.155672
R1240 VTAIL.n829 VTAIL.n759 0.155672
R1241 VTAIL.n837 VTAIL.n759 0.155672
R1242 VTAIL.n838 VTAIL.n837 0.155672
R1243 VTAIL.n838 VTAIL.n755 0.155672
R1244 VTAIL.n845 VTAIL.n755 0.155672
R1245 VTAIL.n846 VTAIL.n845 0.155672
R1246 VTAIL.n846 VTAIL.n751 0.155672
R1247 VTAIL.n853 VTAIL.n751 0.155672
R1248 VTAIL.n40 VTAIL.n39 0.155672
R1249 VTAIL.n40 VTAIL.n31 0.155672
R1250 VTAIL.n47 VTAIL.n31 0.155672
R1251 VTAIL.n48 VTAIL.n47 0.155672
R1252 VTAIL.n48 VTAIL.n27 0.155672
R1253 VTAIL.n55 VTAIL.n27 0.155672
R1254 VTAIL.n56 VTAIL.n55 0.155672
R1255 VTAIL.n56 VTAIL.n23 0.155672
R1256 VTAIL.n63 VTAIL.n23 0.155672
R1257 VTAIL.n64 VTAIL.n63 0.155672
R1258 VTAIL.n64 VTAIL.n19 0.155672
R1259 VTAIL.n71 VTAIL.n19 0.155672
R1260 VTAIL.n72 VTAIL.n71 0.155672
R1261 VTAIL.n72 VTAIL.n15 0.155672
R1262 VTAIL.n80 VTAIL.n15 0.155672
R1263 VTAIL.n81 VTAIL.n80 0.155672
R1264 VTAIL.n81 VTAIL.n11 0.155672
R1265 VTAIL.n89 VTAIL.n11 0.155672
R1266 VTAIL.n90 VTAIL.n89 0.155672
R1267 VTAIL.n90 VTAIL.n7 0.155672
R1268 VTAIL.n97 VTAIL.n7 0.155672
R1269 VTAIL.n98 VTAIL.n97 0.155672
R1270 VTAIL.n98 VTAIL.n3 0.155672
R1271 VTAIL.n105 VTAIL.n3 0.155672
R1272 VTAIL.n146 VTAIL.n145 0.155672
R1273 VTAIL.n146 VTAIL.n137 0.155672
R1274 VTAIL.n153 VTAIL.n137 0.155672
R1275 VTAIL.n154 VTAIL.n153 0.155672
R1276 VTAIL.n154 VTAIL.n133 0.155672
R1277 VTAIL.n161 VTAIL.n133 0.155672
R1278 VTAIL.n162 VTAIL.n161 0.155672
R1279 VTAIL.n162 VTAIL.n129 0.155672
R1280 VTAIL.n169 VTAIL.n129 0.155672
R1281 VTAIL.n170 VTAIL.n169 0.155672
R1282 VTAIL.n170 VTAIL.n125 0.155672
R1283 VTAIL.n177 VTAIL.n125 0.155672
R1284 VTAIL.n178 VTAIL.n177 0.155672
R1285 VTAIL.n178 VTAIL.n121 0.155672
R1286 VTAIL.n186 VTAIL.n121 0.155672
R1287 VTAIL.n187 VTAIL.n186 0.155672
R1288 VTAIL.n187 VTAIL.n117 0.155672
R1289 VTAIL.n195 VTAIL.n117 0.155672
R1290 VTAIL.n196 VTAIL.n195 0.155672
R1291 VTAIL.n196 VTAIL.n113 0.155672
R1292 VTAIL.n203 VTAIL.n113 0.155672
R1293 VTAIL.n204 VTAIL.n203 0.155672
R1294 VTAIL.n204 VTAIL.n109 0.155672
R1295 VTAIL.n211 VTAIL.n109 0.155672
R1296 VTAIL.n254 VTAIL.n253 0.155672
R1297 VTAIL.n254 VTAIL.n245 0.155672
R1298 VTAIL.n261 VTAIL.n245 0.155672
R1299 VTAIL.n262 VTAIL.n261 0.155672
R1300 VTAIL.n262 VTAIL.n241 0.155672
R1301 VTAIL.n269 VTAIL.n241 0.155672
R1302 VTAIL.n270 VTAIL.n269 0.155672
R1303 VTAIL.n270 VTAIL.n237 0.155672
R1304 VTAIL.n277 VTAIL.n237 0.155672
R1305 VTAIL.n278 VTAIL.n277 0.155672
R1306 VTAIL.n278 VTAIL.n233 0.155672
R1307 VTAIL.n285 VTAIL.n233 0.155672
R1308 VTAIL.n286 VTAIL.n285 0.155672
R1309 VTAIL.n286 VTAIL.n229 0.155672
R1310 VTAIL.n294 VTAIL.n229 0.155672
R1311 VTAIL.n295 VTAIL.n294 0.155672
R1312 VTAIL.n295 VTAIL.n225 0.155672
R1313 VTAIL.n303 VTAIL.n225 0.155672
R1314 VTAIL.n304 VTAIL.n303 0.155672
R1315 VTAIL.n304 VTAIL.n221 0.155672
R1316 VTAIL.n311 VTAIL.n221 0.155672
R1317 VTAIL.n312 VTAIL.n311 0.155672
R1318 VTAIL.n312 VTAIL.n217 0.155672
R1319 VTAIL.n319 VTAIL.n217 0.155672
R1320 VTAIL.n747 VTAIL.n645 0.155672
R1321 VTAIL.n740 VTAIL.n645 0.155672
R1322 VTAIL.n740 VTAIL.n739 0.155672
R1323 VTAIL.n739 VTAIL.n649 0.155672
R1324 VTAIL.n732 VTAIL.n649 0.155672
R1325 VTAIL.n732 VTAIL.n731 0.155672
R1326 VTAIL.n731 VTAIL.n653 0.155672
R1327 VTAIL.n723 VTAIL.n653 0.155672
R1328 VTAIL.n723 VTAIL.n722 0.155672
R1329 VTAIL.n722 VTAIL.n657 0.155672
R1330 VTAIL.n715 VTAIL.n657 0.155672
R1331 VTAIL.n715 VTAIL.n714 0.155672
R1332 VTAIL.n714 VTAIL.n662 0.155672
R1333 VTAIL.n707 VTAIL.n662 0.155672
R1334 VTAIL.n707 VTAIL.n706 0.155672
R1335 VTAIL.n706 VTAIL.n666 0.155672
R1336 VTAIL.n699 VTAIL.n666 0.155672
R1337 VTAIL.n699 VTAIL.n698 0.155672
R1338 VTAIL.n698 VTAIL.n670 0.155672
R1339 VTAIL.n691 VTAIL.n670 0.155672
R1340 VTAIL.n691 VTAIL.n690 0.155672
R1341 VTAIL.n690 VTAIL.n674 0.155672
R1342 VTAIL.n683 VTAIL.n674 0.155672
R1343 VTAIL.n683 VTAIL.n682 0.155672
R1344 VTAIL.n639 VTAIL.n537 0.155672
R1345 VTAIL.n632 VTAIL.n537 0.155672
R1346 VTAIL.n632 VTAIL.n631 0.155672
R1347 VTAIL.n631 VTAIL.n541 0.155672
R1348 VTAIL.n624 VTAIL.n541 0.155672
R1349 VTAIL.n624 VTAIL.n623 0.155672
R1350 VTAIL.n623 VTAIL.n545 0.155672
R1351 VTAIL.n615 VTAIL.n545 0.155672
R1352 VTAIL.n615 VTAIL.n614 0.155672
R1353 VTAIL.n614 VTAIL.n549 0.155672
R1354 VTAIL.n607 VTAIL.n549 0.155672
R1355 VTAIL.n607 VTAIL.n606 0.155672
R1356 VTAIL.n606 VTAIL.n554 0.155672
R1357 VTAIL.n599 VTAIL.n554 0.155672
R1358 VTAIL.n599 VTAIL.n598 0.155672
R1359 VTAIL.n598 VTAIL.n558 0.155672
R1360 VTAIL.n591 VTAIL.n558 0.155672
R1361 VTAIL.n591 VTAIL.n590 0.155672
R1362 VTAIL.n590 VTAIL.n562 0.155672
R1363 VTAIL.n583 VTAIL.n562 0.155672
R1364 VTAIL.n583 VTAIL.n582 0.155672
R1365 VTAIL.n582 VTAIL.n566 0.155672
R1366 VTAIL.n575 VTAIL.n566 0.155672
R1367 VTAIL.n575 VTAIL.n574 0.155672
R1368 VTAIL.n533 VTAIL.n431 0.155672
R1369 VTAIL.n526 VTAIL.n431 0.155672
R1370 VTAIL.n526 VTAIL.n525 0.155672
R1371 VTAIL.n525 VTAIL.n435 0.155672
R1372 VTAIL.n518 VTAIL.n435 0.155672
R1373 VTAIL.n518 VTAIL.n517 0.155672
R1374 VTAIL.n517 VTAIL.n439 0.155672
R1375 VTAIL.n509 VTAIL.n439 0.155672
R1376 VTAIL.n509 VTAIL.n508 0.155672
R1377 VTAIL.n508 VTAIL.n443 0.155672
R1378 VTAIL.n501 VTAIL.n443 0.155672
R1379 VTAIL.n501 VTAIL.n500 0.155672
R1380 VTAIL.n500 VTAIL.n448 0.155672
R1381 VTAIL.n493 VTAIL.n448 0.155672
R1382 VTAIL.n493 VTAIL.n492 0.155672
R1383 VTAIL.n492 VTAIL.n452 0.155672
R1384 VTAIL.n485 VTAIL.n452 0.155672
R1385 VTAIL.n485 VTAIL.n484 0.155672
R1386 VTAIL.n484 VTAIL.n456 0.155672
R1387 VTAIL.n477 VTAIL.n456 0.155672
R1388 VTAIL.n477 VTAIL.n476 0.155672
R1389 VTAIL.n476 VTAIL.n460 0.155672
R1390 VTAIL.n469 VTAIL.n460 0.155672
R1391 VTAIL.n469 VTAIL.n468 0.155672
R1392 VTAIL.n425 VTAIL.n323 0.155672
R1393 VTAIL.n418 VTAIL.n323 0.155672
R1394 VTAIL.n418 VTAIL.n417 0.155672
R1395 VTAIL.n417 VTAIL.n327 0.155672
R1396 VTAIL.n410 VTAIL.n327 0.155672
R1397 VTAIL.n410 VTAIL.n409 0.155672
R1398 VTAIL.n409 VTAIL.n331 0.155672
R1399 VTAIL.n401 VTAIL.n331 0.155672
R1400 VTAIL.n401 VTAIL.n400 0.155672
R1401 VTAIL.n400 VTAIL.n335 0.155672
R1402 VTAIL.n393 VTAIL.n335 0.155672
R1403 VTAIL.n393 VTAIL.n392 0.155672
R1404 VTAIL.n392 VTAIL.n340 0.155672
R1405 VTAIL.n385 VTAIL.n340 0.155672
R1406 VTAIL.n385 VTAIL.n384 0.155672
R1407 VTAIL.n384 VTAIL.n344 0.155672
R1408 VTAIL.n377 VTAIL.n344 0.155672
R1409 VTAIL.n377 VTAIL.n376 0.155672
R1410 VTAIL.n376 VTAIL.n348 0.155672
R1411 VTAIL.n369 VTAIL.n348 0.155672
R1412 VTAIL.n369 VTAIL.n368 0.155672
R1413 VTAIL.n368 VTAIL.n352 0.155672
R1414 VTAIL.n361 VTAIL.n352 0.155672
R1415 VTAIL.n361 VTAIL.n360 0.155672
R1416 VTAIL VTAIL.n1 0.0586897
R1417 VDD1 VDD1.n0 71.1886
R1418 VDD1.n3 VDD1.n2 71.0751
R1419 VDD1.n3 VDD1.n1 71.0751
R1420 VDD1.n5 VDD1.n4 69.7423
R1421 VDD1.n5 VDD1.n3 53.1949
R1422 VDD1.n4 VDD1.t4 1.70859
R1423 VDD1.n4 VDD1.t5 1.70859
R1424 VDD1.n0 VDD1.t1 1.70859
R1425 VDD1.n0 VDD1.t3 1.70859
R1426 VDD1.n2 VDD1.t0 1.70859
R1427 VDD1.n2 VDD1.t2 1.70859
R1428 VDD1.n1 VDD1.t6 1.70859
R1429 VDD1.n1 VDD1.t7 1.70859
R1430 VDD1 VDD1.n5 1.33024
R1431 VN.n7 VN.t7 192.218
R1432 VN.n39 VN.t4 192.218
R1433 VN.n59 VN.n31 161.3
R1434 VN.n58 VN.n57 161.3
R1435 VN.n56 VN.n32 161.3
R1436 VN.n55 VN.n54 161.3
R1437 VN.n53 VN.n33 161.3
R1438 VN.n52 VN.n51 161.3
R1439 VN.n50 VN.n34 161.3
R1440 VN.n49 VN.n48 161.3
R1441 VN.n47 VN.n35 161.3
R1442 VN.n46 VN.n45 161.3
R1443 VN.n44 VN.n37 161.3
R1444 VN.n43 VN.n42 161.3
R1445 VN.n41 VN.n38 161.3
R1446 VN.n28 VN.n0 161.3
R1447 VN.n27 VN.n26 161.3
R1448 VN.n25 VN.n1 161.3
R1449 VN.n24 VN.n23 161.3
R1450 VN.n22 VN.n2 161.3
R1451 VN.n21 VN.n20 161.3
R1452 VN.n19 VN.n3 161.3
R1453 VN.n18 VN.n17 161.3
R1454 VN.n15 VN.n4 161.3
R1455 VN.n14 VN.n13 161.3
R1456 VN.n12 VN.n5 161.3
R1457 VN.n11 VN.n10 161.3
R1458 VN.n9 VN.n6 161.3
R1459 VN.n8 VN.t6 158.694
R1460 VN.n16 VN.t0 158.694
R1461 VN.n29 VN.t2 158.694
R1462 VN.n40 VN.t3 158.694
R1463 VN.n36 VN.t5 158.694
R1464 VN.n60 VN.t1 158.694
R1465 VN.n30 VN.n29 106.841
R1466 VN.n61 VN.n60 106.841
R1467 VN VN.n61 57.8542
R1468 VN.n14 VN.n5 56.5193
R1469 VN.n46 VN.n37 56.5193
R1470 VN.n8 VN.n7 56.0641
R1471 VN.n40 VN.n39 56.0641
R1472 VN.n23 VN.n22 43.4072
R1473 VN.n54 VN.n53 43.4072
R1474 VN.n23 VN.n1 37.5796
R1475 VN.n54 VN.n32 37.5796
R1476 VN.n10 VN.n9 24.4675
R1477 VN.n10 VN.n5 24.4675
R1478 VN.n15 VN.n14 24.4675
R1479 VN.n17 VN.n15 24.4675
R1480 VN.n21 VN.n3 24.4675
R1481 VN.n22 VN.n21 24.4675
R1482 VN.n27 VN.n1 24.4675
R1483 VN.n28 VN.n27 24.4675
R1484 VN.n42 VN.n37 24.4675
R1485 VN.n42 VN.n41 24.4675
R1486 VN.n53 VN.n52 24.4675
R1487 VN.n52 VN.n34 24.4675
R1488 VN.n48 VN.n47 24.4675
R1489 VN.n47 VN.n46 24.4675
R1490 VN.n59 VN.n58 24.4675
R1491 VN.n58 VN.n32 24.4675
R1492 VN.n9 VN.n8 17.6167
R1493 VN.n17 VN.n16 17.6167
R1494 VN.n41 VN.n40 17.6167
R1495 VN.n48 VN.n36 17.6167
R1496 VN.n16 VN.n3 6.85126
R1497 VN.n36 VN.n34 6.85126
R1498 VN.n39 VN.n38 5.02778
R1499 VN.n7 VN.n6 5.02778
R1500 VN.n29 VN.n28 3.91522
R1501 VN.n60 VN.n59 3.91522
R1502 VN.n61 VN.n31 0.278367
R1503 VN.n30 VN.n0 0.278367
R1504 VN.n57 VN.n31 0.189894
R1505 VN.n57 VN.n56 0.189894
R1506 VN.n56 VN.n55 0.189894
R1507 VN.n55 VN.n33 0.189894
R1508 VN.n51 VN.n33 0.189894
R1509 VN.n51 VN.n50 0.189894
R1510 VN.n50 VN.n49 0.189894
R1511 VN.n49 VN.n35 0.189894
R1512 VN.n45 VN.n35 0.189894
R1513 VN.n45 VN.n44 0.189894
R1514 VN.n44 VN.n43 0.189894
R1515 VN.n43 VN.n38 0.189894
R1516 VN.n11 VN.n6 0.189894
R1517 VN.n12 VN.n11 0.189894
R1518 VN.n13 VN.n12 0.189894
R1519 VN.n13 VN.n4 0.189894
R1520 VN.n18 VN.n4 0.189894
R1521 VN.n19 VN.n18 0.189894
R1522 VN.n20 VN.n19 0.189894
R1523 VN.n20 VN.n2 0.189894
R1524 VN.n24 VN.n2 0.189894
R1525 VN.n25 VN.n24 0.189894
R1526 VN.n26 VN.n25 0.189894
R1527 VN.n26 VN.n0 0.189894
R1528 VN VN.n30 0.153454
R1529 VDD2.n2 VDD2.n1 71.0751
R1530 VDD2.n2 VDD2.n0 71.0751
R1531 VDD2 VDD2.n5 71.072
R1532 VDD2.n4 VDD2.n3 69.7425
R1533 VDD2.n4 VDD2.n2 52.6118
R1534 VDD2.n5 VDD2.t4 1.70859
R1535 VDD2.n5 VDD2.t3 1.70859
R1536 VDD2.n3 VDD2.t6 1.70859
R1537 VDD2.n3 VDD2.t2 1.70859
R1538 VDD2.n1 VDD2.t7 1.70859
R1539 VDD2.n1 VDD2.t5 1.70859
R1540 VDD2.n0 VDD2.t0 1.70859
R1541 VDD2.n0 VDD2.t1 1.70859
R1542 VDD2 VDD2.n4 1.44662
R1543 B.n539 B.n538 585
R1544 B.n537 B.n158 585
R1545 B.n536 B.n535 585
R1546 B.n534 B.n159 585
R1547 B.n533 B.n532 585
R1548 B.n531 B.n160 585
R1549 B.n530 B.n529 585
R1550 B.n528 B.n161 585
R1551 B.n527 B.n526 585
R1552 B.n525 B.n162 585
R1553 B.n524 B.n523 585
R1554 B.n522 B.n163 585
R1555 B.n521 B.n520 585
R1556 B.n519 B.n164 585
R1557 B.n518 B.n517 585
R1558 B.n516 B.n165 585
R1559 B.n515 B.n514 585
R1560 B.n513 B.n166 585
R1561 B.n512 B.n511 585
R1562 B.n510 B.n167 585
R1563 B.n509 B.n508 585
R1564 B.n507 B.n168 585
R1565 B.n506 B.n505 585
R1566 B.n504 B.n169 585
R1567 B.n503 B.n502 585
R1568 B.n501 B.n170 585
R1569 B.n500 B.n499 585
R1570 B.n498 B.n171 585
R1571 B.n497 B.n496 585
R1572 B.n495 B.n172 585
R1573 B.n494 B.n493 585
R1574 B.n492 B.n173 585
R1575 B.n491 B.n490 585
R1576 B.n489 B.n174 585
R1577 B.n488 B.n487 585
R1578 B.n486 B.n175 585
R1579 B.n485 B.n484 585
R1580 B.n483 B.n176 585
R1581 B.n482 B.n481 585
R1582 B.n480 B.n177 585
R1583 B.n479 B.n478 585
R1584 B.n477 B.n178 585
R1585 B.n476 B.n475 585
R1586 B.n474 B.n179 585
R1587 B.n473 B.n472 585
R1588 B.n471 B.n180 585
R1589 B.n470 B.n469 585
R1590 B.n468 B.n181 585
R1591 B.n467 B.n466 585
R1592 B.n465 B.n182 585
R1593 B.n464 B.n463 585
R1594 B.n462 B.n183 585
R1595 B.n461 B.n460 585
R1596 B.n459 B.n184 585
R1597 B.n458 B.n457 585
R1598 B.n456 B.n185 585
R1599 B.n455 B.n454 585
R1600 B.n453 B.n186 585
R1601 B.n452 B.n451 585
R1602 B.n450 B.n187 585
R1603 B.n449 B.n448 585
R1604 B.n447 B.n188 585
R1605 B.n445 B.n444 585
R1606 B.n443 B.n191 585
R1607 B.n442 B.n441 585
R1608 B.n440 B.n192 585
R1609 B.n439 B.n438 585
R1610 B.n437 B.n193 585
R1611 B.n436 B.n435 585
R1612 B.n434 B.n194 585
R1613 B.n433 B.n432 585
R1614 B.n431 B.n195 585
R1615 B.n430 B.n429 585
R1616 B.n425 B.n196 585
R1617 B.n424 B.n423 585
R1618 B.n422 B.n197 585
R1619 B.n421 B.n420 585
R1620 B.n419 B.n198 585
R1621 B.n418 B.n417 585
R1622 B.n416 B.n199 585
R1623 B.n415 B.n414 585
R1624 B.n413 B.n200 585
R1625 B.n412 B.n411 585
R1626 B.n410 B.n201 585
R1627 B.n409 B.n408 585
R1628 B.n407 B.n202 585
R1629 B.n406 B.n405 585
R1630 B.n404 B.n203 585
R1631 B.n403 B.n402 585
R1632 B.n401 B.n204 585
R1633 B.n400 B.n399 585
R1634 B.n398 B.n205 585
R1635 B.n397 B.n396 585
R1636 B.n395 B.n206 585
R1637 B.n394 B.n393 585
R1638 B.n392 B.n207 585
R1639 B.n391 B.n390 585
R1640 B.n389 B.n208 585
R1641 B.n388 B.n387 585
R1642 B.n386 B.n209 585
R1643 B.n385 B.n384 585
R1644 B.n383 B.n210 585
R1645 B.n382 B.n381 585
R1646 B.n380 B.n211 585
R1647 B.n379 B.n378 585
R1648 B.n377 B.n212 585
R1649 B.n376 B.n375 585
R1650 B.n374 B.n213 585
R1651 B.n373 B.n372 585
R1652 B.n371 B.n214 585
R1653 B.n370 B.n369 585
R1654 B.n368 B.n215 585
R1655 B.n367 B.n366 585
R1656 B.n365 B.n216 585
R1657 B.n364 B.n363 585
R1658 B.n362 B.n217 585
R1659 B.n361 B.n360 585
R1660 B.n359 B.n218 585
R1661 B.n358 B.n357 585
R1662 B.n356 B.n219 585
R1663 B.n355 B.n354 585
R1664 B.n353 B.n220 585
R1665 B.n352 B.n351 585
R1666 B.n350 B.n221 585
R1667 B.n349 B.n348 585
R1668 B.n347 B.n222 585
R1669 B.n346 B.n345 585
R1670 B.n344 B.n223 585
R1671 B.n343 B.n342 585
R1672 B.n341 B.n224 585
R1673 B.n340 B.n339 585
R1674 B.n338 B.n225 585
R1675 B.n337 B.n336 585
R1676 B.n335 B.n226 585
R1677 B.n540 B.n157 585
R1678 B.n542 B.n541 585
R1679 B.n543 B.n156 585
R1680 B.n545 B.n544 585
R1681 B.n546 B.n155 585
R1682 B.n548 B.n547 585
R1683 B.n549 B.n154 585
R1684 B.n551 B.n550 585
R1685 B.n552 B.n153 585
R1686 B.n554 B.n553 585
R1687 B.n555 B.n152 585
R1688 B.n557 B.n556 585
R1689 B.n558 B.n151 585
R1690 B.n560 B.n559 585
R1691 B.n561 B.n150 585
R1692 B.n563 B.n562 585
R1693 B.n564 B.n149 585
R1694 B.n566 B.n565 585
R1695 B.n567 B.n148 585
R1696 B.n569 B.n568 585
R1697 B.n570 B.n147 585
R1698 B.n572 B.n571 585
R1699 B.n573 B.n146 585
R1700 B.n575 B.n574 585
R1701 B.n576 B.n145 585
R1702 B.n578 B.n577 585
R1703 B.n579 B.n144 585
R1704 B.n581 B.n580 585
R1705 B.n582 B.n143 585
R1706 B.n584 B.n583 585
R1707 B.n585 B.n142 585
R1708 B.n587 B.n586 585
R1709 B.n588 B.n141 585
R1710 B.n590 B.n589 585
R1711 B.n591 B.n140 585
R1712 B.n593 B.n592 585
R1713 B.n594 B.n139 585
R1714 B.n596 B.n595 585
R1715 B.n597 B.n138 585
R1716 B.n599 B.n598 585
R1717 B.n600 B.n137 585
R1718 B.n602 B.n601 585
R1719 B.n603 B.n136 585
R1720 B.n605 B.n604 585
R1721 B.n606 B.n135 585
R1722 B.n608 B.n607 585
R1723 B.n609 B.n134 585
R1724 B.n611 B.n610 585
R1725 B.n612 B.n133 585
R1726 B.n614 B.n613 585
R1727 B.n615 B.n132 585
R1728 B.n617 B.n616 585
R1729 B.n618 B.n131 585
R1730 B.n620 B.n619 585
R1731 B.n621 B.n130 585
R1732 B.n623 B.n622 585
R1733 B.n624 B.n129 585
R1734 B.n626 B.n625 585
R1735 B.n627 B.n128 585
R1736 B.n629 B.n628 585
R1737 B.n630 B.n127 585
R1738 B.n632 B.n631 585
R1739 B.n633 B.n126 585
R1740 B.n635 B.n634 585
R1741 B.n636 B.n125 585
R1742 B.n638 B.n637 585
R1743 B.n639 B.n124 585
R1744 B.n641 B.n640 585
R1745 B.n642 B.n123 585
R1746 B.n644 B.n643 585
R1747 B.n645 B.n122 585
R1748 B.n647 B.n646 585
R1749 B.n648 B.n121 585
R1750 B.n650 B.n649 585
R1751 B.n651 B.n120 585
R1752 B.n653 B.n652 585
R1753 B.n654 B.n119 585
R1754 B.n656 B.n655 585
R1755 B.n657 B.n118 585
R1756 B.n659 B.n658 585
R1757 B.n660 B.n117 585
R1758 B.n662 B.n661 585
R1759 B.n663 B.n116 585
R1760 B.n665 B.n664 585
R1761 B.n666 B.n115 585
R1762 B.n668 B.n667 585
R1763 B.n669 B.n114 585
R1764 B.n671 B.n670 585
R1765 B.n672 B.n113 585
R1766 B.n674 B.n673 585
R1767 B.n675 B.n112 585
R1768 B.n677 B.n676 585
R1769 B.n678 B.n111 585
R1770 B.n680 B.n679 585
R1771 B.n681 B.n110 585
R1772 B.n683 B.n682 585
R1773 B.n684 B.n109 585
R1774 B.n686 B.n685 585
R1775 B.n687 B.n108 585
R1776 B.n689 B.n688 585
R1777 B.n690 B.n107 585
R1778 B.n692 B.n691 585
R1779 B.n693 B.n106 585
R1780 B.n695 B.n694 585
R1781 B.n696 B.n105 585
R1782 B.n698 B.n697 585
R1783 B.n699 B.n104 585
R1784 B.n701 B.n700 585
R1785 B.n702 B.n103 585
R1786 B.n704 B.n703 585
R1787 B.n705 B.n102 585
R1788 B.n707 B.n706 585
R1789 B.n909 B.n908 585
R1790 B.n907 B.n30 585
R1791 B.n906 B.n905 585
R1792 B.n904 B.n31 585
R1793 B.n903 B.n902 585
R1794 B.n901 B.n32 585
R1795 B.n900 B.n899 585
R1796 B.n898 B.n33 585
R1797 B.n897 B.n896 585
R1798 B.n895 B.n34 585
R1799 B.n894 B.n893 585
R1800 B.n892 B.n35 585
R1801 B.n891 B.n890 585
R1802 B.n889 B.n36 585
R1803 B.n888 B.n887 585
R1804 B.n886 B.n37 585
R1805 B.n885 B.n884 585
R1806 B.n883 B.n38 585
R1807 B.n882 B.n881 585
R1808 B.n880 B.n39 585
R1809 B.n879 B.n878 585
R1810 B.n877 B.n40 585
R1811 B.n876 B.n875 585
R1812 B.n874 B.n41 585
R1813 B.n873 B.n872 585
R1814 B.n871 B.n42 585
R1815 B.n870 B.n869 585
R1816 B.n868 B.n43 585
R1817 B.n867 B.n866 585
R1818 B.n865 B.n44 585
R1819 B.n864 B.n863 585
R1820 B.n862 B.n45 585
R1821 B.n861 B.n860 585
R1822 B.n859 B.n46 585
R1823 B.n858 B.n857 585
R1824 B.n856 B.n47 585
R1825 B.n855 B.n854 585
R1826 B.n853 B.n48 585
R1827 B.n852 B.n851 585
R1828 B.n850 B.n49 585
R1829 B.n849 B.n848 585
R1830 B.n847 B.n50 585
R1831 B.n846 B.n845 585
R1832 B.n844 B.n51 585
R1833 B.n843 B.n842 585
R1834 B.n841 B.n52 585
R1835 B.n840 B.n839 585
R1836 B.n838 B.n53 585
R1837 B.n837 B.n836 585
R1838 B.n835 B.n54 585
R1839 B.n834 B.n833 585
R1840 B.n832 B.n55 585
R1841 B.n831 B.n830 585
R1842 B.n829 B.n56 585
R1843 B.n828 B.n827 585
R1844 B.n826 B.n57 585
R1845 B.n825 B.n824 585
R1846 B.n823 B.n58 585
R1847 B.n822 B.n821 585
R1848 B.n820 B.n59 585
R1849 B.n819 B.n818 585
R1850 B.n817 B.n60 585
R1851 B.n816 B.n815 585
R1852 B.n814 B.n61 585
R1853 B.n813 B.n812 585
R1854 B.n811 B.n65 585
R1855 B.n810 B.n809 585
R1856 B.n808 B.n66 585
R1857 B.n807 B.n806 585
R1858 B.n805 B.n67 585
R1859 B.n804 B.n803 585
R1860 B.n802 B.n68 585
R1861 B.n800 B.n799 585
R1862 B.n798 B.n71 585
R1863 B.n797 B.n796 585
R1864 B.n795 B.n72 585
R1865 B.n794 B.n793 585
R1866 B.n792 B.n73 585
R1867 B.n791 B.n790 585
R1868 B.n789 B.n74 585
R1869 B.n788 B.n787 585
R1870 B.n786 B.n75 585
R1871 B.n785 B.n784 585
R1872 B.n783 B.n76 585
R1873 B.n782 B.n781 585
R1874 B.n780 B.n77 585
R1875 B.n779 B.n778 585
R1876 B.n777 B.n78 585
R1877 B.n776 B.n775 585
R1878 B.n774 B.n79 585
R1879 B.n773 B.n772 585
R1880 B.n771 B.n80 585
R1881 B.n770 B.n769 585
R1882 B.n768 B.n81 585
R1883 B.n767 B.n766 585
R1884 B.n765 B.n82 585
R1885 B.n764 B.n763 585
R1886 B.n762 B.n83 585
R1887 B.n761 B.n760 585
R1888 B.n759 B.n84 585
R1889 B.n758 B.n757 585
R1890 B.n756 B.n85 585
R1891 B.n755 B.n754 585
R1892 B.n753 B.n86 585
R1893 B.n752 B.n751 585
R1894 B.n750 B.n87 585
R1895 B.n749 B.n748 585
R1896 B.n747 B.n88 585
R1897 B.n746 B.n745 585
R1898 B.n744 B.n89 585
R1899 B.n743 B.n742 585
R1900 B.n741 B.n90 585
R1901 B.n740 B.n739 585
R1902 B.n738 B.n91 585
R1903 B.n737 B.n736 585
R1904 B.n735 B.n92 585
R1905 B.n734 B.n733 585
R1906 B.n732 B.n93 585
R1907 B.n731 B.n730 585
R1908 B.n729 B.n94 585
R1909 B.n728 B.n727 585
R1910 B.n726 B.n95 585
R1911 B.n725 B.n724 585
R1912 B.n723 B.n96 585
R1913 B.n722 B.n721 585
R1914 B.n720 B.n97 585
R1915 B.n719 B.n718 585
R1916 B.n717 B.n98 585
R1917 B.n716 B.n715 585
R1918 B.n714 B.n99 585
R1919 B.n713 B.n712 585
R1920 B.n711 B.n100 585
R1921 B.n710 B.n709 585
R1922 B.n708 B.n101 585
R1923 B.n910 B.n29 585
R1924 B.n912 B.n911 585
R1925 B.n913 B.n28 585
R1926 B.n915 B.n914 585
R1927 B.n916 B.n27 585
R1928 B.n918 B.n917 585
R1929 B.n919 B.n26 585
R1930 B.n921 B.n920 585
R1931 B.n922 B.n25 585
R1932 B.n924 B.n923 585
R1933 B.n925 B.n24 585
R1934 B.n927 B.n926 585
R1935 B.n928 B.n23 585
R1936 B.n930 B.n929 585
R1937 B.n931 B.n22 585
R1938 B.n933 B.n932 585
R1939 B.n934 B.n21 585
R1940 B.n936 B.n935 585
R1941 B.n937 B.n20 585
R1942 B.n939 B.n938 585
R1943 B.n940 B.n19 585
R1944 B.n942 B.n941 585
R1945 B.n943 B.n18 585
R1946 B.n945 B.n944 585
R1947 B.n946 B.n17 585
R1948 B.n948 B.n947 585
R1949 B.n949 B.n16 585
R1950 B.n951 B.n950 585
R1951 B.n952 B.n15 585
R1952 B.n954 B.n953 585
R1953 B.n955 B.n14 585
R1954 B.n957 B.n956 585
R1955 B.n958 B.n13 585
R1956 B.n960 B.n959 585
R1957 B.n961 B.n12 585
R1958 B.n963 B.n962 585
R1959 B.n964 B.n11 585
R1960 B.n966 B.n965 585
R1961 B.n967 B.n10 585
R1962 B.n969 B.n968 585
R1963 B.n970 B.n9 585
R1964 B.n972 B.n971 585
R1965 B.n973 B.n8 585
R1966 B.n975 B.n974 585
R1967 B.n976 B.n7 585
R1968 B.n978 B.n977 585
R1969 B.n979 B.n6 585
R1970 B.n981 B.n980 585
R1971 B.n982 B.n5 585
R1972 B.n984 B.n983 585
R1973 B.n985 B.n4 585
R1974 B.n987 B.n986 585
R1975 B.n988 B.n3 585
R1976 B.n990 B.n989 585
R1977 B.n991 B.n0 585
R1978 B.n2 B.n1 585
R1979 B.n254 B.n253 585
R1980 B.n256 B.n255 585
R1981 B.n257 B.n252 585
R1982 B.n259 B.n258 585
R1983 B.n260 B.n251 585
R1984 B.n262 B.n261 585
R1985 B.n263 B.n250 585
R1986 B.n265 B.n264 585
R1987 B.n266 B.n249 585
R1988 B.n268 B.n267 585
R1989 B.n269 B.n248 585
R1990 B.n271 B.n270 585
R1991 B.n272 B.n247 585
R1992 B.n274 B.n273 585
R1993 B.n275 B.n246 585
R1994 B.n277 B.n276 585
R1995 B.n278 B.n245 585
R1996 B.n280 B.n279 585
R1997 B.n281 B.n244 585
R1998 B.n283 B.n282 585
R1999 B.n284 B.n243 585
R2000 B.n286 B.n285 585
R2001 B.n287 B.n242 585
R2002 B.n289 B.n288 585
R2003 B.n290 B.n241 585
R2004 B.n292 B.n291 585
R2005 B.n293 B.n240 585
R2006 B.n295 B.n294 585
R2007 B.n296 B.n239 585
R2008 B.n298 B.n297 585
R2009 B.n299 B.n238 585
R2010 B.n301 B.n300 585
R2011 B.n302 B.n237 585
R2012 B.n304 B.n303 585
R2013 B.n305 B.n236 585
R2014 B.n307 B.n306 585
R2015 B.n308 B.n235 585
R2016 B.n310 B.n309 585
R2017 B.n311 B.n234 585
R2018 B.n313 B.n312 585
R2019 B.n314 B.n233 585
R2020 B.n316 B.n315 585
R2021 B.n317 B.n232 585
R2022 B.n319 B.n318 585
R2023 B.n320 B.n231 585
R2024 B.n322 B.n321 585
R2025 B.n323 B.n230 585
R2026 B.n325 B.n324 585
R2027 B.n326 B.n229 585
R2028 B.n328 B.n327 585
R2029 B.n329 B.n228 585
R2030 B.n331 B.n330 585
R2031 B.n332 B.n227 585
R2032 B.n334 B.n333 585
R2033 B.n189 B.t10 564.919
R2034 B.n69 B.t5 564.919
R2035 B.n426 B.t7 564.918
R2036 B.n62 B.t2 564.918
R2037 B.n333 B.n226 506.916
R2038 B.n540 B.n539 506.916
R2039 B.n708 B.n707 506.916
R2040 B.n908 B.n29 506.916
R2041 B.n190 B.t11 502.471
R2042 B.n70 B.t4 502.471
R2043 B.n427 B.t8 502.471
R2044 B.n63 B.t1 502.471
R2045 B.n426 B.t6 367.139
R2046 B.n189 B.t9 367.139
R2047 B.n69 B.t3 367.139
R2048 B.n62 B.t0 367.139
R2049 B.n993 B.n992 256.663
R2050 B.n992 B.n991 235.042
R2051 B.n992 B.n2 235.042
R2052 B.n337 B.n226 163.367
R2053 B.n338 B.n337 163.367
R2054 B.n339 B.n338 163.367
R2055 B.n339 B.n224 163.367
R2056 B.n343 B.n224 163.367
R2057 B.n344 B.n343 163.367
R2058 B.n345 B.n344 163.367
R2059 B.n345 B.n222 163.367
R2060 B.n349 B.n222 163.367
R2061 B.n350 B.n349 163.367
R2062 B.n351 B.n350 163.367
R2063 B.n351 B.n220 163.367
R2064 B.n355 B.n220 163.367
R2065 B.n356 B.n355 163.367
R2066 B.n357 B.n356 163.367
R2067 B.n357 B.n218 163.367
R2068 B.n361 B.n218 163.367
R2069 B.n362 B.n361 163.367
R2070 B.n363 B.n362 163.367
R2071 B.n363 B.n216 163.367
R2072 B.n367 B.n216 163.367
R2073 B.n368 B.n367 163.367
R2074 B.n369 B.n368 163.367
R2075 B.n369 B.n214 163.367
R2076 B.n373 B.n214 163.367
R2077 B.n374 B.n373 163.367
R2078 B.n375 B.n374 163.367
R2079 B.n375 B.n212 163.367
R2080 B.n379 B.n212 163.367
R2081 B.n380 B.n379 163.367
R2082 B.n381 B.n380 163.367
R2083 B.n381 B.n210 163.367
R2084 B.n385 B.n210 163.367
R2085 B.n386 B.n385 163.367
R2086 B.n387 B.n386 163.367
R2087 B.n387 B.n208 163.367
R2088 B.n391 B.n208 163.367
R2089 B.n392 B.n391 163.367
R2090 B.n393 B.n392 163.367
R2091 B.n393 B.n206 163.367
R2092 B.n397 B.n206 163.367
R2093 B.n398 B.n397 163.367
R2094 B.n399 B.n398 163.367
R2095 B.n399 B.n204 163.367
R2096 B.n403 B.n204 163.367
R2097 B.n404 B.n403 163.367
R2098 B.n405 B.n404 163.367
R2099 B.n405 B.n202 163.367
R2100 B.n409 B.n202 163.367
R2101 B.n410 B.n409 163.367
R2102 B.n411 B.n410 163.367
R2103 B.n411 B.n200 163.367
R2104 B.n415 B.n200 163.367
R2105 B.n416 B.n415 163.367
R2106 B.n417 B.n416 163.367
R2107 B.n417 B.n198 163.367
R2108 B.n421 B.n198 163.367
R2109 B.n422 B.n421 163.367
R2110 B.n423 B.n422 163.367
R2111 B.n423 B.n196 163.367
R2112 B.n430 B.n196 163.367
R2113 B.n431 B.n430 163.367
R2114 B.n432 B.n431 163.367
R2115 B.n432 B.n194 163.367
R2116 B.n436 B.n194 163.367
R2117 B.n437 B.n436 163.367
R2118 B.n438 B.n437 163.367
R2119 B.n438 B.n192 163.367
R2120 B.n442 B.n192 163.367
R2121 B.n443 B.n442 163.367
R2122 B.n444 B.n443 163.367
R2123 B.n444 B.n188 163.367
R2124 B.n449 B.n188 163.367
R2125 B.n450 B.n449 163.367
R2126 B.n451 B.n450 163.367
R2127 B.n451 B.n186 163.367
R2128 B.n455 B.n186 163.367
R2129 B.n456 B.n455 163.367
R2130 B.n457 B.n456 163.367
R2131 B.n457 B.n184 163.367
R2132 B.n461 B.n184 163.367
R2133 B.n462 B.n461 163.367
R2134 B.n463 B.n462 163.367
R2135 B.n463 B.n182 163.367
R2136 B.n467 B.n182 163.367
R2137 B.n468 B.n467 163.367
R2138 B.n469 B.n468 163.367
R2139 B.n469 B.n180 163.367
R2140 B.n473 B.n180 163.367
R2141 B.n474 B.n473 163.367
R2142 B.n475 B.n474 163.367
R2143 B.n475 B.n178 163.367
R2144 B.n479 B.n178 163.367
R2145 B.n480 B.n479 163.367
R2146 B.n481 B.n480 163.367
R2147 B.n481 B.n176 163.367
R2148 B.n485 B.n176 163.367
R2149 B.n486 B.n485 163.367
R2150 B.n487 B.n486 163.367
R2151 B.n487 B.n174 163.367
R2152 B.n491 B.n174 163.367
R2153 B.n492 B.n491 163.367
R2154 B.n493 B.n492 163.367
R2155 B.n493 B.n172 163.367
R2156 B.n497 B.n172 163.367
R2157 B.n498 B.n497 163.367
R2158 B.n499 B.n498 163.367
R2159 B.n499 B.n170 163.367
R2160 B.n503 B.n170 163.367
R2161 B.n504 B.n503 163.367
R2162 B.n505 B.n504 163.367
R2163 B.n505 B.n168 163.367
R2164 B.n509 B.n168 163.367
R2165 B.n510 B.n509 163.367
R2166 B.n511 B.n510 163.367
R2167 B.n511 B.n166 163.367
R2168 B.n515 B.n166 163.367
R2169 B.n516 B.n515 163.367
R2170 B.n517 B.n516 163.367
R2171 B.n517 B.n164 163.367
R2172 B.n521 B.n164 163.367
R2173 B.n522 B.n521 163.367
R2174 B.n523 B.n522 163.367
R2175 B.n523 B.n162 163.367
R2176 B.n527 B.n162 163.367
R2177 B.n528 B.n527 163.367
R2178 B.n529 B.n528 163.367
R2179 B.n529 B.n160 163.367
R2180 B.n533 B.n160 163.367
R2181 B.n534 B.n533 163.367
R2182 B.n535 B.n534 163.367
R2183 B.n535 B.n158 163.367
R2184 B.n539 B.n158 163.367
R2185 B.n707 B.n102 163.367
R2186 B.n703 B.n102 163.367
R2187 B.n703 B.n702 163.367
R2188 B.n702 B.n701 163.367
R2189 B.n701 B.n104 163.367
R2190 B.n697 B.n104 163.367
R2191 B.n697 B.n696 163.367
R2192 B.n696 B.n695 163.367
R2193 B.n695 B.n106 163.367
R2194 B.n691 B.n106 163.367
R2195 B.n691 B.n690 163.367
R2196 B.n690 B.n689 163.367
R2197 B.n689 B.n108 163.367
R2198 B.n685 B.n108 163.367
R2199 B.n685 B.n684 163.367
R2200 B.n684 B.n683 163.367
R2201 B.n683 B.n110 163.367
R2202 B.n679 B.n110 163.367
R2203 B.n679 B.n678 163.367
R2204 B.n678 B.n677 163.367
R2205 B.n677 B.n112 163.367
R2206 B.n673 B.n112 163.367
R2207 B.n673 B.n672 163.367
R2208 B.n672 B.n671 163.367
R2209 B.n671 B.n114 163.367
R2210 B.n667 B.n114 163.367
R2211 B.n667 B.n666 163.367
R2212 B.n666 B.n665 163.367
R2213 B.n665 B.n116 163.367
R2214 B.n661 B.n116 163.367
R2215 B.n661 B.n660 163.367
R2216 B.n660 B.n659 163.367
R2217 B.n659 B.n118 163.367
R2218 B.n655 B.n118 163.367
R2219 B.n655 B.n654 163.367
R2220 B.n654 B.n653 163.367
R2221 B.n653 B.n120 163.367
R2222 B.n649 B.n120 163.367
R2223 B.n649 B.n648 163.367
R2224 B.n648 B.n647 163.367
R2225 B.n647 B.n122 163.367
R2226 B.n643 B.n122 163.367
R2227 B.n643 B.n642 163.367
R2228 B.n642 B.n641 163.367
R2229 B.n641 B.n124 163.367
R2230 B.n637 B.n124 163.367
R2231 B.n637 B.n636 163.367
R2232 B.n636 B.n635 163.367
R2233 B.n635 B.n126 163.367
R2234 B.n631 B.n126 163.367
R2235 B.n631 B.n630 163.367
R2236 B.n630 B.n629 163.367
R2237 B.n629 B.n128 163.367
R2238 B.n625 B.n128 163.367
R2239 B.n625 B.n624 163.367
R2240 B.n624 B.n623 163.367
R2241 B.n623 B.n130 163.367
R2242 B.n619 B.n130 163.367
R2243 B.n619 B.n618 163.367
R2244 B.n618 B.n617 163.367
R2245 B.n617 B.n132 163.367
R2246 B.n613 B.n132 163.367
R2247 B.n613 B.n612 163.367
R2248 B.n612 B.n611 163.367
R2249 B.n611 B.n134 163.367
R2250 B.n607 B.n134 163.367
R2251 B.n607 B.n606 163.367
R2252 B.n606 B.n605 163.367
R2253 B.n605 B.n136 163.367
R2254 B.n601 B.n136 163.367
R2255 B.n601 B.n600 163.367
R2256 B.n600 B.n599 163.367
R2257 B.n599 B.n138 163.367
R2258 B.n595 B.n138 163.367
R2259 B.n595 B.n594 163.367
R2260 B.n594 B.n593 163.367
R2261 B.n593 B.n140 163.367
R2262 B.n589 B.n140 163.367
R2263 B.n589 B.n588 163.367
R2264 B.n588 B.n587 163.367
R2265 B.n587 B.n142 163.367
R2266 B.n583 B.n142 163.367
R2267 B.n583 B.n582 163.367
R2268 B.n582 B.n581 163.367
R2269 B.n581 B.n144 163.367
R2270 B.n577 B.n144 163.367
R2271 B.n577 B.n576 163.367
R2272 B.n576 B.n575 163.367
R2273 B.n575 B.n146 163.367
R2274 B.n571 B.n146 163.367
R2275 B.n571 B.n570 163.367
R2276 B.n570 B.n569 163.367
R2277 B.n569 B.n148 163.367
R2278 B.n565 B.n148 163.367
R2279 B.n565 B.n564 163.367
R2280 B.n564 B.n563 163.367
R2281 B.n563 B.n150 163.367
R2282 B.n559 B.n150 163.367
R2283 B.n559 B.n558 163.367
R2284 B.n558 B.n557 163.367
R2285 B.n557 B.n152 163.367
R2286 B.n553 B.n152 163.367
R2287 B.n553 B.n552 163.367
R2288 B.n552 B.n551 163.367
R2289 B.n551 B.n154 163.367
R2290 B.n547 B.n154 163.367
R2291 B.n547 B.n546 163.367
R2292 B.n546 B.n545 163.367
R2293 B.n545 B.n156 163.367
R2294 B.n541 B.n156 163.367
R2295 B.n541 B.n540 163.367
R2296 B.n908 B.n907 163.367
R2297 B.n907 B.n906 163.367
R2298 B.n906 B.n31 163.367
R2299 B.n902 B.n31 163.367
R2300 B.n902 B.n901 163.367
R2301 B.n901 B.n900 163.367
R2302 B.n900 B.n33 163.367
R2303 B.n896 B.n33 163.367
R2304 B.n896 B.n895 163.367
R2305 B.n895 B.n894 163.367
R2306 B.n894 B.n35 163.367
R2307 B.n890 B.n35 163.367
R2308 B.n890 B.n889 163.367
R2309 B.n889 B.n888 163.367
R2310 B.n888 B.n37 163.367
R2311 B.n884 B.n37 163.367
R2312 B.n884 B.n883 163.367
R2313 B.n883 B.n882 163.367
R2314 B.n882 B.n39 163.367
R2315 B.n878 B.n39 163.367
R2316 B.n878 B.n877 163.367
R2317 B.n877 B.n876 163.367
R2318 B.n876 B.n41 163.367
R2319 B.n872 B.n41 163.367
R2320 B.n872 B.n871 163.367
R2321 B.n871 B.n870 163.367
R2322 B.n870 B.n43 163.367
R2323 B.n866 B.n43 163.367
R2324 B.n866 B.n865 163.367
R2325 B.n865 B.n864 163.367
R2326 B.n864 B.n45 163.367
R2327 B.n860 B.n45 163.367
R2328 B.n860 B.n859 163.367
R2329 B.n859 B.n858 163.367
R2330 B.n858 B.n47 163.367
R2331 B.n854 B.n47 163.367
R2332 B.n854 B.n853 163.367
R2333 B.n853 B.n852 163.367
R2334 B.n852 B.n49 163.367
R2335 B.n848 B.n49 163.367
R2336 B.n848 B.n847 163.367
R2337 B.n847 B.n846 163.367
R2338 B.n846 B.n51 163.367
R2339 B.n842 B.n51 163.367
R2340 B.n842 B.n841 163.367
R2341 B.n841 B.n840 163.367
R2342 B.n840 B.n53 163.367
R2343 B.n836 B.n53 163.367
R2344 B.n836 B.n835 163.367
R2345 B.n835 B.n834 163.367
R2346 B.n834 B.n55 163.367
R2347 B.n830 B.n55 163.367
R2348 B.n830 B.n829 163.367
R2349 B.n829 B.n828 163.367
R2350 B.n828 B.n57 163.367
R2351 B.n824 B.n57 163.367
R2352 B.n824 B.n823 163.367
R2353 B.n823 B.n822 163.367
R2354 B.n822 B.n59 163.367
R2355 B.n818 B.n59 163.367
R2356 B.n818 B.n817 163.367
R2357 B.n817 B.n816 163.367
R2358 B.n816 B.n61 163.367
R2359 B.n812 B.n61 163.367
R2360 B.n812 B.n811 163.367
R2361 B.n811 B.n810 163.367
R2362 B.n810 B.n66 163.367
R2363 B.n806 B.n66 163.367
R2364 B.n806 B.n805 163.367
R2365 B.n805 B.n804 163.367
R2366 B.n804 B.n68 163.367
R2367 B.n799 B.n68 163.367
R2368 B.n799 B.n798 163.367
R2369 B.n798 B.n797 163.367
R2370 B.n797 B.n72 163.367
R2371 B.n793 B.n72 163.367
R2372 B.n793 B.n792 163.367
R2373 B.n792 B.n791 163.367
R2374 B.n791 B.n74 163.367
R2375 B.n787 B.n74 163.367
R2376 B.n787 B.n786 163.367
R2377 B.n786 B.n785 163.367
R2378 B.n785 B.n76 163.367
R2379 B.n781 B.n76 163.367
R2380 B.n781 B.n780 163.367
R2381 B.n780 B.n779 163.367
R2382 B.n779 B.n78 163.367
R2383 B.n775 B.n78 163.367
R2384 B.n775 B.n774 163.367
R2385 B.n774 B.n773 163.367
R2386 B.n773 B.n80 163.367
R2387 B.n769 B.n80 163.367
R2388 B.n769 B.n768 163.367
R2389 B.n768 B.n767 163.367
R2390 B.n767 B.n82 163.367
R2391 B.n763 B.n82 163.367
R2392 B.n763 B.n762 163.367
R2393 B.n762 B.n761 163.367
R2394 B.n761 B.n84 163.367
R2395 B.n757 B.n84 163.367
R2396 B.n757 B.n756 163.367
R2397 B.n756 B.n755 163.367
R2398 B.n755 B.n86 163.367
R2399 B.n751 B.n86 163.367
R2400 B.n751 B.n750 163.367
R2401 B.n750 B.n749 163.367
R2402 B.n749 B.n88 163.367
R2403 B.n745 B.n88 163.367
R2404 B.n745 B.n744 163.367
R2405 B.n744 B.n743 163.367
R2406 B.n743 B.n90 163.367
R2407 B.n739 B.n90 163.367
R2408 B.n739 B.n738 163.367
R2409 B.n738 B.n737 163.367
R2410 B.n737 B.n92 163.367
R2411 B.n733 B.n92 163.367
R2412 B.n733 B.n732 163.367
R2413 B.n732 B.n731 163.367
R2414 B.n731 B.n94 163.367
R2415 B.n727 B.n94 163.367
R2416 B.n727 B.n726 163.367
R2417 B.n726 B.n725 163.367
R2418 B.n725 B.n96 163.367
R2419 B.n721 B.n96 163.367
R2420 B.n721 B.n720 163.367
R2421 B.n720 B.n719 163.367
R2422 B.n719 B.n98 163.367
R2423 B.n715 B.n98 163.367
R2424 B.n715 B.n714 163.367
R2425 B.n714 B.n713 163.367
R2426 B.n713 B.n100 163.367
R2427 B.n709 B.n100 163.367
R2428 B.n709 B.n708 163.367
R2429 B.n912 B.n29 163.367
R2430 B.n913 B.n912 163.367
R2431 B.n914 B.n913 163.367
R2432 B.n914 B.n27 163.367
R2433 B.n918 B.n27 163.367
R2434 B.n919 B.n918 163.367
R2435 B.n920 B.n919 163.367
R2436 B.n920 B.n25 163.367
R2437 B.n924 B.n25 163.367
R2438 B.n925 B.n924 163.367
R2439 B.n926 B.n925 163.367
R2440 B.n926 B.n23 163.367
R2441 B.n930 B.n23 163.367
R2442 B.n931 B.n930 163.367
R2443 B.n932 B.n931 163.367
R2444 B.n932 B.n21 163.367
R2445 B.n936 B.n21 163.367
R2446 B.n937 B.n936 163.367
R2447 B.n938 B.n937 163.367
R2448 B.n938 B.n19 163.367
R2449 B.n942 B.n19 163.367
R2450 B.n943 B.n942 163.367
R2451 B.n944 B.n943 163.367
R2452 B.n944 B.n17 163.367
R2453 B.n948 B.n17 163.367
R2454 B.n949 B.n948 163.367
R2455 B.n950 B.n949 163.367
R2456 B.n950 B.n15 163.367
R2457 B.n954 B.n15 163.367
R2458 B.n955 B.n954 163.367
R2459 B.n956 B.n955 163.367
R2460 B.n956 B.n13 163.367
R2461 B.n960 B.n13 163.367
R2462 B.n961 B.n960 163.367
R2463 B.n962 B.n961 163.367
R2464 B.n962 B.n11 163.367
R2465 B.n966 B.n11 163.367
R2466 B.n967 B.n966 163.367
R2467 B.n968 B.n967 163.367
R2468 B.n968 B.n9 163.367
R2469 B.n972 B.n9 163.367
R2470 B.n973 B.n972 163.367
R2471 B.n974 B.n973 163.367
R2472 B.n974 B.n7 163.367
R2473 B.n978 B.n7 163.367
R2474 B.n979 B.n978 163.367
R2475 B.n980 B.n979 163.367
R2476 B.n980 B.n5 163.367
R2477 B.n984 B.n5 163.367
R2478 B.n985 B.n984 163.367
R2479 B.n986 B.n985 163.367
R2480 B.n986 B.n3 163.367
R2481 B.n990 B.n3 163.367
R2482 B.n991 B.n990 163.367
R2483 B.n254 B.n2 163.367
R2484 B.n255 B.n254 163.367
R2485 B.n255 B.n252 163.367
R2486 B.n259 B.n252 163.367
R2487 B.n260 B.n259 163.367
R2488 B.n261 B.n260 163.367
R2489 B.n261 B.n250 163.367
R2490 B.n265 B.n250 163.367
R2491 B.n266 B.n265 163.367
R2492 B.n267 B.n266 163.367
R2493 B.n267 B.n248 163.367
R2494 B.n271 B.n248 163.367
R2495 B.n272 B.n271 163.367
R2496 B.n273 B.n272 163.367
R2497 B.n273 B.n246 163.367
R2498 B.n277 B.n246 163.367
R2499 B.n278 B.n277 163.367
R2500 B.n279 B.n278 163.367
R2501 B.n279 B.n244 163.367
R2502 B.n283 B.n244 163.367
R2503 B.n284 B.n283 163.367
R2504 B.n285 B.n284 163.367
R2505 B.n285 B.n242 163.367
R2506 B.n289 B.n242 163.367
R2507 B.n290 B.n289 163.367
R2508 B.n291 B.n290 163.367
R2509 B.n291 B.n240 163.367
R2510 B.n295 B.n240 163.367
R2511 B.n296 B.n295 163.367
R2512 B.n297 B.n296 163.367
R2513 B.n297 B.n238 163.367
R2514 B.n301 B.n238 163.367
R2515 B.n302 B.n301 163.367
R2516 B.n303 B.n302 163.367
R2517 B.n303 B.n236 163.367
R2518 B.n307 B.n236 163.367
R2519 B.n308 B.n307 163.367
R2520 B.n309 B.n308 163.367
R2521 B.n309 B.n234 163.367
R2522 B.n313 B.n234 163.367
R2523 B.n314 B.n313 163.367
R2524 B.n315 B.n314 163.367
R2525 B.n315 B.n232 163.367
R2526 B.n319 B.n232 163.367
R2527 B.n320 B.n319 163.367
R2528 B.n321 B.n320 163.367
R2529 B.n321 B.n230 163.367
R2530 B.n325 B.n230 163.367
R2531 B.n326 B.n325 163.367
R2532 B.n327 B.n326 163.367
R2533 B.n327 B.n228 163.367
R2534 B.n331 B.n228 163.367
R2535 B.n332 B.n331 163.367
R2536 B.n333 B.n332 163.367
R2537 B.n427 B.n426 62.449
R2538 B.n190 B.n189 62.449
R2539 B.n70 B.n69 62.449
R2540 B.n63 B.n62 62.449
R2541 B.n428 B.n427 59.5399
R2542 B.n446 B.n190 59.5399
R2543 B.n801 B.n70 59.5399
R2544 B.n64 B.n63 59.5399
R2545 B.n910 B.n909 32.9371
R2546 B.n706 B.n101 32.9371
R2547 B.n538 B.n157 32.9371
R2548 B.n335 B.n334 32.9371
R2549 B B.n993 18.0485
R2550 B.n911 B.n910 10.6151
R2551 B.n911 B.n28 10.6151
R2552 B.n915 B.n28 10.6151
R2553 B.n916 B.n915 10.6151
R2554 B.n917 B.n916 10.6151
R2555 B.n917 B.n26 10.6151
R2556 B.n921 B.n26 10.6151
R2557 B.n922 B.n921 10.6151
R2558 B.n923 B.n922 10.6151
R2559 B.n923 B.n24 10.6151
R2560 B.n927 B.n24 10.6151
R2561 B.n928 B.n927 10.6151
R2562 B.n929 B.n928 10.6151
R2563 B.n929 B.n22 10.6151
R2564 B.n933 B.n22 10.6151
R2565 B.n934 B.n933 10.6151
R2566 B.n935 B.n934 10.6151
R2567 B.n935 B.n20 10.6151
R2568 B.n939 B.n20 10.6151
R2569 B.n940 B.n939 10.6151
R2570 B.n941 B.n940 10.6151
R2571 B.n941 B.n18 10.6151
R2572 B.n945 B.n18 10.6151
R2573 B.n946 B.n945 10.6151
R2574 B.n947 B.n946 10.6151
R2575 B.n947 B.n16 10.6151
R2576 B.n951 B.n16 10.6151
R2577 B.n952 B.n951 10.6151
R2578 B.n953 B.n952 10.6151
R2579 B.n953 B.n14 10.6151
R2580 B.n957 B.n14 10.6151
R2581 B.n958 B.n957 10.6151
R2582 B.n959 B.n958 10.6151
R2583 B.n959 B.n12 10.6151
R2584 B.n963 B.n12 10.6151
R2585 B.n964 B.n963 10.6151
R2586 B.n965 B.n964 10.6151
R2587 B.n965 B.n10 10.6151
R2588 B.n969 B.n10 10.6151
R2589 B.n970 B.n969 10.6151
R2590 B.n971 B.n970 10.6151
R2591 B.n971 B.n8 10.6151
R2592 B.n975 B.n8 10.6151
R2593 B.n976 B.n975 10.6151
R2594 B.n977 B.n976 10.6151
R2595 B.n977 B.n6 10.6151
R2596 B.n981 B.n6 10.6151
R2597 B.n982 B.n981 10.6151
R2598 B.n983 B.n982 10.6151
R2599 B.n983 B.n4 10.6151
R2600 B.n987 B.n4 10.6151
R2601 B.n988 B.n987 10.6151
R2602 B.n989 B.n988 10.6151
R2603 B.n989 B.n0 10.6151
R2604 B.n909 B.n30 10.6151
R2605 B.n905 B.n30 10.6151
R2606 B.n905 B.n904 10.6151
R2607 B.n904 B.n903 10.6151
R2608 B.n903 B.n32 10.6151
R2609 B.n899 B.n32 10.6151
R2610 B.n899 B.n898 10.6151
R2611 B.n898 B.n897 10.6151
R2612 B.n897 B.n34 10.6151
R2613 B.n893 B.n34 10.6151
R2614 B.n893 B.n892 10.6151
R2615 B.n892 B.n891 10.6151
R2616 B.n891 B.n36 10.6151
R2617 B.n887 B.n36 10.6151
R2618 B.n887 B.n886 10.6151
R2619 B.n886 B.n885 10.6151
R2620 B.n885 B.n38 10.6151
R2621 B.n881 B.n38 10.6151
R2622 B.n881 B.n880 10.6151
R2623 B.n880 B.n879 10.6151
R2624 B.n879 B.n40 10.6151
R2625 B.n875 B.n40 10.6151
R2626 B.n875 B.n874 10.6151
R2627 B.n874 B.n873 10.6151
R2628 B.n873 B.n42 10.6151
R2629 B.n869 B.n42 10.6151
R2630 B.n869 B.n868 10.6151
R2631 B.n868 B.n867 10.6151
R2632 B.n867 B.n44 10.6151
R2633 B.n863 B.n44 10.6151
R2634 B.n863 B.n862 10.6151
R2635 B.n862 B.n861 10.6151
R2636 B.n861 B.n46 10.6151
R2637 B.n857 B.n46 10.6151
R2638 B.n857 B.n856 10.6151
R2639 B.n856 B.n855 10.6151
R2640 B.n855 B.n48 10.6151
R2641 B.n851 B.n48 10.6151
R2642 B.n851 B.n850 10.6151
R2643 B.n850 B.n849 10.6151
R2644 B.n849 B.n50 10.6151
R2645 B.n845 B.n50 10.6151
R2646 B.n845 B.n844 10.6151
R2647 B.n844 B.n843 10.6151
R2648 B.n843 B.n52 10.6151
R2649 B.n839 B.n52 10.6151
R2650 B.n839 B.n838 10.6151
R2651 B.n838 B.n837 10.6151
R2652 B.n837 B.n54 10.6151
R2653 B.n833 B.n54 10.6151
R2654 B.n833 B.n832 10.6151
R2655 B.n832 B.n831 10.6151
R2656 B.n831 B.n56 10.6151
R2657 B.n827 B.n56 10.6151
R2658 B.n827 B.n826 10.6151
R2659 B.n826 B.n825 10.6151
R2660 B.n825 B.n58 10.6151
R2661 B.n821 B.n58 10.6151
R2662 B.n821 B.n820 10.6151
R2663 B.n820 B.n819 10.6151
R2664 B.n819 B.n60 10.6151
R2665 B.n815 B.n814 10.6151
R2666 B.n814 B.n813 10.6151
R2667 B.n813 B.n65 10.6151
R2668 B.n809 B.n65 10.6151
R2669 B.n809 B.n808 10.6151
R2670 B.n808 B.n807 10.6151
R2671 B.n807 B.n67 10.6151
R2672 B.n803 B.n67 10.6151
R2673 B.n803 B.n802 10.6151
R2674 B.n800 B.n71 10.6151
R2675 B.n796 B.n71 10.6151
R2676 B.n796 B.n795 10.6151
R2677 B.n795 B.n794 10.6151
R2678 B.n794 B.n73 10.6151
R2679 B.n790 B.n73 10.6151
R2680 B.n790 B.n789 10.6151
R2681 B.n789 B.n788 10.6151
R2682 B.n788 B.n75 10.6151
R2683 B.n784 B.n75 10.6151
R2684 B.n784 B.n783 10.6151
R2685 B.n783 B.n782 10.6151
R2686 B.n782 B.n77 10.6151
R2687 B.n778 B.n77 10.6151
R2688 B.n778 B.n777 10.6151
R2689 B.n777 B.n776 10.6151
R2690 B.n776 B.n79 10.6151
R2691 B.n772 B.n79 10.6151
R2692 B.n772 B.n771 10.6151
R2693 B.n771 B.n770 10.6151
R2694 B.n770 B.n81 10.6151
R2695 B.n766 B.n81 10.6151
R2696 B.n766 B.n765 10.6151
R2697 B.n765 B.n764 10.6151
R2698 B.n764 B.n83 10.6151
R2699 B.n760 B.n83 10.6151
R2700 B.n760 B.n759 10.6151
R2701 B.n759 B.n758 10.6151
R2702 B.n758 B.n85 10.6151
R2703 B.n754 B.n85 10.6151
R2704 B.n754 B.n753 10.6151
R2705 B.n753 B.n752 10.6151
R2706 B.n752 B.n87 10.6151
R2707 B.n748 B.n87 10.6151
R2708 B.n748 B.n747 10.6151
R2709 B.n747 B.n746 10.6151
R2710 B.n746 B.n89 10.6151
R2711 B.n742 B.n89 10.6151
R2712 B.n742 B.n741 10.6151
R2713 B.n741 B.n740 10.6151
R2714 B.n740 B.n91 10.6151
R2715 B.n736 B.n91 10.6151
R2716 B.n736 B.n735 10.6151
R2717 B.n735 B.n734 10.6151
R2718 B.n734 B.n93 10.6151
R2719 B.n730 B.n93 10.6151
R2720 B.n730 B.n729 10.6151
R2721 B.n729 B.n728 10.6151
R2722 B.n728 B.n95 10.6151
R2723 B.n724 B.n95 10.6151
R2724 B.n724 B.n723 10.6151
R2725 B.n723 B.n722 10.6151
R2726 B.n722 B.n97 10.6151
R2727 B.n718 B.n97 10.6151
R2728 B.n718 B.n717 10.6151
R2729 B.n717 B.n716 10.6151
R2730 B.n716 B.n99 10.6151
R2731 B.n712 B.n99 10.6151
R2732 B.n712 B.n711 10.6151
R2733 B.n711 B.n710 10.6151
R2734 B.n710 B.n101 10.6151
R2735 B.n706 B.n705 10.6151
R2736 B.n705 B.n704 10.6151
R2737 B.n704 B.n103 10.6151
R2738 B.n700 B.n103 10.6151
R2739 B.n700 B.n699 10.6151
R2740 B.n699 B.n698 10.6151
R2741 B.n698 B.n105 10.6151
R2742 B.n694 B.n105 10.6151
R2743 B.n694 B.n693 10.6151
R2744 B.n693 B.n692 10.6151
R2745 B.n692 B.n107 10.6151
R2746 B.n688 B.n107 10.6151
R2747 B.n688 B.n687 10.6151
R2748 B.n687 B.n686 10.6151
R2749 B.n686 B.n109 10.6151
R2750 B.n682 B.n109 10.6151
R2751 B.n682 B.n681 10.6151
R2752 B.n681 B.n680 10.6151
R2753 B.n680 B.n111 10.6151
R2754 B.n676 B.n111 10.6151
R2755 B.n676 B.n675 10.6151
R2756 B.n675 B.n674 10.6151
R2757 B.n674 B.n113 10.6151
R2758 B.n670 B.n113 10.6151
R2759 B.n670 B.n669 10.6151
R2760 B.n669 B.n668 10.6151
R2761 B.n668 B.n115 10.6151
R2762 B.n664 B.n115 10.6151
R2763 B.n664 B.n663 10.6151
R2764 B.n663 B.n662 10.6151
R2765 B.n662 B.n117 10.6151
R2766 B.n658 B.n117 10.6151
R2767 B.n658 B.n657 10.6151
R2768 B.n657 B.n656 10.6151
R2769 B.n656 B.n119 10.6151
R2770 B.n652 B.n119 10.6151
R2771 B.n652 B.n651 10.6151
R2772 B.n651 B.n650 10.6151
R2773 B.n650 B.n121 10.6151
R2774 B.n646 B.n121 10.6151
R2775 B.n646 B.n645 10.6151
R2776 B.n645 B.n644 10.6151
R2777 B.n644 B.n123 10.6151
R2778 B.n640 B.n123 10.6151
R2779 B.n640 B.n639 10.6151
R2780 B.n639 B.n638 10.6151
R2781 B.n638 B.n125 10.6151
R2782 B.n634 B.n125 10.6151
R2783 B.n634 B.n633 10.6151
R2784 B.n633 B.n632 10.6151
R2785 B.n632 B.n127 10.6151
R2786 B.n628 B.n127 10.6151
R2787 B.n628 B.n627 10.6151
R2788 B.n627 B.n626 10.6151
R2789 B.n626 B.n129 10.6151
R2790 B.n622 B.n129 10.6151
R2791 B.n622 B.n621 10.6151
R2792 B.n621 B.n620 10.6151
R2793 B.n620 B.n131 10.6151
R2794 B.n616 B.n131 10.6151
R2795 B.n616 B.n615 10.6151
R2796 B.n615 B.n614 10.6151
R2797 B.n614 B.n133 10.6151
R2798 B.n610 B.n133 10.6151
R2799 B.n610 B.n609 10.6151
R2800 B.n609 B.n608 10.6151
R2801 B.n608 B.n135 10.6151
R2802 B.n604 B.n135 10.6151
R2803 B.n604 B.n603 10.6151
R2804 B.n603 B.n602 10.6151
R2805 B.n602 B.n137 10.6151
R2806 B.n598 B.n137 10.6151
R2807 B.n598 B.n597 10.6151
R2808 B.n597 B.n596 10.6151
R2809 B.n596 B.n139 10.6151
R2810 B.n592 B.n139 10.6151
R2811 B.n592 B.n591 10.6151
R2812 B.n591 B.n590 10.6151
R2813 B.n590 B.n141 10.6151
R2814 B.n586 B.n141 10.6151
R2815 B.n586 B.n585 10.6151
R2816 B.n585 B.n584 10.6151
R2817 B.n584 B.n143 10.6151
R2818 B.n580 B.n143 10.6151
R2819 B.n580 B.n579 10.6151
R2820 B.n579 B.n578 10.6151
R2821 B.n578 B.n145 10.6151
R2822 B.n574 B.n145 10.6151
R2823 B.n574 B.n573 10.6151
R2824 B.n573 B.n572 10.6151
R2825 B.n572 B.n147 10.6151
R2826 B.n568 B.n147 10.6151
R2827 B.n568 B.n567 10.6151
R2828 B.n567 B.n566 10.6151
R2829 B.n566 B.n149 10.6151
R2830 B.n562 B.n149 10.6151
R2831 B.n562 B.n561 10.6151
R2832 B.n561 B.n560 10.6151
R2833 B.n560 B.n151 10.6151
R2834 B.n556 B.n151 10.6151
R2835 B.n556 B.n555 10.6151
R2836 B.n555 B.n554 10.6151
R2837 B.n554 B.n153 10.6151
R2838 B.n550 B.n153 10.6151
R2839 B.n550 B.n549 10.6151
R2840 B.n549 B.n548 10.6151
R2841 B.n548 B.n155 10.6151
R2842 B.n544 B.n155 10.6151
R2843 B.n544 B.n543 10.6151
R2844 B.n543 B.n542 10.6151
R2845 B.n542 B.n157 10.6151
R2846 B.n253 B.n1 10.6151
R2847 B.n256 B.n253 10.6151
R2848 B.n257 B.n256 10.6151
R2849 B.n258 B.n257 10.6151
R2850 B.n258 B.n251 10.6151
R2851 B.n262 B.n251 10.6151
R2852 B.n263 B.n262 10.6151
R2853 B.n264 B.n263 10.6151
R2854 B.n264 B.n249 10.6151
R2855 B.n268 B.n249 10.6151
R2856 B.n269 B.n268 10.6151
R2857 B.n270 B.n269 10.6151
R2858 B.n270 B.n247 10.6151
R2859 B.n274 B.n247 10.6151
R2860 B.n275 B.n274 10.6151
R2861 B.n276 B.n275 10.6151
R2862 B.n276 B.n245 10.6151
R2863 B.n280 B.n245 10.6151
R2864 B.n281 B.n280 10.6151
R2865 B.n282 B.n281 10.6151
R2866 B.n282 B.n243 10.6151
R2867 B.n286 B.n243 10.6151
R2868 B.n287 B.n286 10.6151
R2869 B.n288 B.n287 10.6151
R2870 B.n288 B.n241 10.6151
R2871 B.n292 B.n241 10.6151
R2872 B.n293 B.n292 10.6151
R2873 B.n294 B.n293 10.6151
R2874 B.n294 B.n239 10.6151
R2875 B.n298 B.n239 10.6151
R2876 B.n299 B.n298 10.6151
R2877 B.n300 B.n299 10.6151
R2878 B.n300 B.n237 10.6151
R2879 B.n304 B.n237 10.6151
R2880 B.n305 B.n304 10.6151
R2881 B.n306 B.n305 10.6151
R2882 B.n306 B.n235 10.6151
R2883 B.n310 B.n235 10.6151
R2884 B.n311 B.n310 10.6151
R2885 B.n312 B.n311 10.6151
R2886 B.n312 B.n233 10.6151
R2887 B.n316 B.n233 10.6151
R2888 B.n317 B.n316 10.6151
R2889 B.n318 B.n317 10.6151
R2890 B.n318 B.n231 10.6151
R2891 B.n322 B.n231 10.6151
R2892 B.n323 B.n322 10.6151
R2893 B.n324 B.n323 10.6151
R2894 B.n324 B.n229 10.6151
R2895 B.n328 B.n229 10.6151
R2896 B.n329 B.n328 10.6151
R2897 B.n330 B.n329 10.6151
R2898 B.n330 B.n227 10.6151
R2899 B.n334 B.n227 10.6151
R2900 B.n336 B.n335 10.6151
R2901 B.n336 B.n225 10.6151
R2902 B.n340 B.n225 10.6151
R2903 B.n341 B.n340 10.6151
R2904 B.n342 B.n341 10.6151
R2905 B.n342 B.n223 10.6151
R2906 B.n346 B.n223 10.6151
R2907 B.n347 B.n346 10.6151
R2908 B.n348 B.n347 10.6151
R2909 B.n348 B.n221 10.6151
R2910 B.n352 B.n221 10.6151
R2911 B.n353 B.n352 10.6151
R2912 B.n354 B.n353 10.6151
R2913 B.n354 B.n219 10.6151
R2914 B.n358 B.n219 10.6151
R2915 B.n359 B.n358 10.6151
R2916 B.n360 B.n359 10.6151
R2917 B.n360 B.n217 10.6151
R2918 B.n364 B.n217 10.6151
R2919 B.n365 B.n364 10.6151
R2920 B.n366 B.n365 10.6151
R2921 B.n366 B.n215 10.6151
R2922 B.n370 B.n215 10.6151
R2923 B.n371 B.n370 10.6151
R2924 B.n372 B.n371 10.6151
R2925 B.n372 B.n213 10.6151
R2926 B.n376 B.n213 10.6151
R2927 B.n377 B.n376 10.6151
R2928 B.n378 B.n377 10.6151
R2929 B.n378 B.n211 10.6151
R2930 B.n382 B.n211 10.6151
R2931 B.n383 B.n382 10.6151
R2932 B.n384 B.n383 10.6151
R2933 B.n384 B.n209 10.6151
R2934 B.n388 B.n209 10.6151
R2935 B.n389 B.n388 10.6151
R2936 B.n390 B.n389 10.6151
R2937 B.n390 B.n207 10.6151
R2938 B.n394 B.n207 10.6151
R2939 B.n395 B.n394 10.6151
R2940 B.n396 B.n395 10.6151
R2941 B.n396 B.n205 10.6151
R2942 B.n400 B.n205 10.6151
R2943 B.n401 B.n400 10.6151
R2944 B.n402 B.n401 10.6151
R2945 B.n402 B.n203 10.6151
R2946 B.n406 B.n203 10.6151
R2947 B.n407 B.n406 10.6151
R2948 B.n408 B.n407 10.6151
R2949 B.n408 B.n201 10.6151
R2950 B.n412 B.n201 10.6151
R2951 B.n413 B.n412 10.6151
R2952 B.n414 B.n413 10.6151
R2953 B.n414 B.n199 10.6151
R2954 B.n418 B.n199 10.6151
R2955 B.n419 B.n418 10.6151
R2956 B.n420 B.n419 10.6151
R2957 B.n420 B.n197 10.6151
R2958 B.n424 B.n197 10.6151
R2959 B.n425 B.n424 10.6151
R2960 B.n429 B.n425 10.6151
R2961 B.n433 B.n195 10.6151
R2962 B.n434 B.n433 10.6151
R2963 B.n435 B.n434 10.6151
R2964 B.n435 B.n193 10.6151
R2965 B.n439 B.n193 10.6151
R2966 B.n440 B.n439 10.6151
R2967 B.n441 B.n440 10.6151
R2968 B.n441 B.n191 10.6151
R2969 B.n445 B.n191 10.6151
R2970 B.n448 B.n447 10.6151
R2971 B.n448 B.n187 10.6151
R2972 B.n452 B.n187 10.6151
R2973 B.n453 B.n452 10.6151
R2974 B.n454 B.n453 10.6151
R2975 B.n454 B.n185 10.6151
R2976 B.n458 B.n185 10.6151
R2977 B.n459 B.n458 10.6151
R2978 B.n460 B.n459 10.6151
R2979 B.n460 B.n183 10.6151
R2980 B.n464 B.n183 10.6151
R2981 B.n465 B.n464 10.6151
R2982 B.n466 B.n465 10.6151
R2983 B.n466 B.n181 10.6151
R2984 B.n470 B.n181 10.6151
R2985 B.n471 B.n470 10.6151
R2986 B.n472 B.n471 10.6151
R2987 B.n472 B.n179 10.6151
R2988 B.n476 B.n179 10.6151
R2989 B.n477 B.n476 10.6151
R2990 B.n478 B.n477 10.6151
R2991 B.n478 B.n177 10.6151
R2992 B.n482 B.n177 10.6151
R2993 B.n483 B.n482 10.6151
R2994 B.n484 B.n483 10.6151
R2995 B.n484 B.n175 10.6151
R2996 B.n488 B.n175 10.6151
R2997 B.n489 B.n488 10.6151
R2998 B.n490 B.n489 10.6151
R2999 B.n490 B.n173 10.6151
R3000 B.n494 B.n173 10.6151
R3001 B.n495 B.n494 10.6151
R3002 B.n496 B.n495 10.6151
R3003 B.n496 B.n171 10.6151
R3004 B.n500 B.n171 10.6151
R3005 B.n501 B.n500 10.6151
R3006 B.n502 B.n501 10.6151
R3007 B.n502 B.n169 10.6151
R3008 B.n506 B.n169 10.6151
R3009 B.n507 B.n506 10.6151
R3010 B.n508 B.n507 10.6151
R3011 B.n508 B.n167 10.6151
R3012 B.n512 B.n167 10.6151
R3013 B.n513 B.n512 10.6151
R3014 B.n514 B.n513 10.6151
R3015 B.n514 B.n165 10.6151
R3016 B.n518 B.n165 10.6151
R3017 B.n519 B.n518 10.6151
R3018 B.n520 B.n519 10.6151
R3019 B.n520 B.n163 10.6151
R3020 B.n524 B.n163 10.6151
R3021 B.n525 B.n524 10.6151
R3022 B.n526 B.n525 10.6151
R3023 B.n526 B.n161 10.6151
R3024 B.n530 B.n161 10.6151
R3025 B.n531 B.n530 10.6151
R3026 B.n532 B.n531 10.6151
R3027 B.n532 B.n159 10.6151
R3028 B.n536 B.n159 10.6151
R3029 B.n537 B.n536 10.6151
R3030 B.n538 B.n537 10.6151
R3031 B.n64 B.n60 9.36635
R3032 B.n801 B.n800 9.36635
R3033 B.n429 B.n428 9.36635
R3034 B.n447 B.n446 9.36635
R3035 B.n993 B.n0 8.11757
R3036 B.n993 B.n1 8.11757
R3037 B.n815 B.n64 1.24928
R3038 B.n802 B.n801 1.24928
R3039 B.n428 B.n195 1.24928
R3040 B.n446 B.n445 1.24928
C0 VP VTAIL 13.9868f
C1 B w_n4190_n4774# 12.530701f
C2 VTAIL VDD2 10.443501f
C3 w_n4190_n4774# VDD1 2.23132f
C4 VP w_n4190_n4774# 9.28115f
C5 w_n4190_n4774# VDD2 2.35819f
C6 B VDD1 1.92651f
C7 B VP 2.29008f
C8 VP VDD1 14.201f
C9 B VDD2 2.03166f
C10 VDD1 VDD2 1.92577f
C11 VP VDD2 0.55015f
C12 VN VTAIL 13.9727f
C13 w_n4190_n4774# VN 8.736341f
C14 w_n4190_n4774# VTAIL 5.80219f
C15 B VN 1.37525f
C16 VN VDD1 0.151873f
C17 B VTAIL 7.45626f
C18 VP VN 9.31742f
C19 VTAIL VDD1 10.3872f
C20 VN VDD2 13.8043f
C21 VDD2 VSUBS 2.22222f
C22 VDD1 VSUBS 2.83364f
C23 VTAIL VSUBS 1.702503f
C24 VN VSUBS 7.38771f
C25 VP VSUBS 4.133156f
C26 B VSUBS 5.922937f
C27 w_n4190_n4774# VSUBS 0.244411p
C28 B.n0 VSUBS 0.006258f
C29 B.n1 VSUBS 0.006258f
C30 B.n2 VSUBS 0.009255f
C31 B.n3 VSUBS 0.007092f
C32 B.n4 VSUBS 0.007092f
C33 B.n5 VSUBS 0.007092f
C34 B.n6 VSUBS 0.007092f
C35 B.n7 VSUBS 0.007092f
C36 B.n8 VSUBS 0.007092f
C37 B.n9 VSUBS 0.007092f
C38 B.n10 VSUBS 0.007092f
C39 B.n11 VSUBS 0.007092f
C40 B.n12 VSUBS 0.007092f
C41 B.n13 VSUBS 0.007092f
C42 B.n14 VSUBS 0.007092f
C43 B.n15 VSUBS 0.007092f
C44 B.n16 VSUBS 0.007092f
C45 B.n17 VSUBS 0.007092f
C46 B.n18 VSUBS 0.007092f
C47 B.n19 VSUBS 0.007092f
C48 B.n20 VSUBS 0.007092f
C49 B.n21 VSUBS 0.007092f
C50 B.n22 VSUBS 0.007092f
C51 B.n23 VSUBS 0.007092f
C52 B.n24 VSUBS 0.007092f
C53 B.n25 VSUBS 0.007092f
C54 B.n26 VSUBS 0.007092f
C55 B.n27 VSUBS 0.007092f
C56 B.n28 VSUBS 0.007092f
C57 B.n29 VSUBS 0.016373f
C58 B.n30 VSUBS 0.007092f
C59 B.n31 VSUBS 0.007092f
C60 B.n32 VSUBS 0.007092f
C61 B.n33 VSUBS 0.007092f
C62 B.n34 VSUBS 0.007092f
C63 B.n35 VSUBS 0.007092f
C64 B.n36 VSUBS 0.007092f
C65 B.n37 VSUBS 0.007092f
C66 B.n38 VSUBS 0.007092f
C67 B.n39 VSUBS 0.007092f
C68 B.n40 VSUBS 0.007092f
C69 B.n41 VSUBS 0.007092f
C70 B.n42 VSUBS 0.007092f
C71 B.n43 VSUBS 0.007092f
C72 B.n44 VSUBS 0.007092f
C73 B.n45 VSUBS 0.007092f
C74 B.n46 VSUBS 0.007092f
C75 B.n47 VSUBS 0.007092f
C76 B.n48 VSUBS 0.007092f
C77 B.n49 VSUBS 0.007092f
C78 B.n50 VSUBS 0.007092f
C79 B.n51 VSUBS 0.007092f
C80 B.n52 VSUBS 0.007092f
C81 B.n53 VSUBS 0.007092f
C82 B.n54 VSUBS 0.007092f
C83 B.n55 VSUBS 0.007092f
C84 B.n56 VSUBS 0.007092f
C85 B.n57 VSUBS 0.007092f
C86 B.n58 VSUBS 0.007092f
C87 B.n59 VSUBS 0.007092f
C88 B.n60 VSUBS 0.006675f
C89 B.n61 VSUBS 0.007092f
C90 B.t1 VSUBS 0.381283f
C91 B.t2 VSUBS 0.418458f
C92 B.t0 VSUBS 2.48169f
C93 B.n62 VSUBS 0.648033f
C94 B.n63 VSUBS 0.346405f
C95 B.n64 VSUBS 0.016432f
C96 B.n65 VSUBS 0.007092f
C97 B.n66 VSUBS 0.007092f
C98 B.n67 VSUBS 0.007092f
C99 B.n68 VSUBS 0.007092f
C100 B.t4 VSUBS 0.381287f
C101 B.t5 VSUBS 0.418461f
C102 B.t3 VSUBS 2.48169f
C103 B.n69 VSUBS 0.64803f
C104 B.n70 VSUBS 0.346402f
C105 B.n71 VSUBS 0.007092f
C106 B.n72 VSUBS 0.007092f
C107 B.n73 VSUBS 0.007092f
C108 B.n74 VSUBS 0.007092f
C109 B.n75 VSUBS 0.007092f
C110 B.n76 VSUBS 0.007092f
C111 B.n77 VSUBS 0.007092f
C112 B.n78 VSUBS 0.007092f
C113 B.n79 VSUBS 0.007092f
C114 B.n80 VSUBS 0.007092f
C115 B.n81 VSUBS 0.007092f
C116 B.n82 VSUBS 0.007092f
C117 B.n83 VSUBS 0.007092f
C118 B.n84 VSUBS 0.007092f
C119 B.n85 VSUBS 0.007092f
C120 B.n86 VSUBS 0.007092f
C121 B.n87 VSUBS 0.007092f
C122 B.n88 VSUBS 0.007092f
C123 B.n89 VSUBS 0.007092f
C124 B.n90 VSUBS 0.007092f
C125 B.n91 VSUBS 0.007092f
C126 B.n92 VSUBS 0.007092f
C127 B.n93 VSUBS 0.007092f
C128 B.n94 VSUBS 0.007092f
C129 B.n95 VSUBS 0.007092f
C130 B.n96 VSUBS 0.007092f
C131 B.n97 VSUBS 0.007092f
C132 B.n98 VSUBS 0.007092f
C133 B.n99 VSUBS 0.007092f
C134 B.n100 VSUBS 0.007092f
C135 B.n101 VSUBS 0.017002f
C136 B.n102 VSUBS 0.007092f
C137 B.n103 VSUBS 0.007092f
C138 B.n104 VSUBS 0.007092f
C139 B.n105 VSUBS 0.007092f
C140 B.n106 VSUBS 0.007092f
C141 B.n107 VSUBS 0.007092f
C142 B.n108 VSUBS 0.007092f
C143 B.n109 VSUBS 0.007092f
C144 B.n110 VSUBS 0.007092f
C145 B.n111 VSUBS 0.007092f
C146 B.n112 VSUBS 0.007092f
C147 B.n113 VSUBS 0.007092f
C148 B.n114 VSUBS 0.007092f
C149 B.n115 VSUBS 0.007092f
C150 B.n116 VSUBS 0.007092f
C151 B.n117 VSUBS 0.007092f
C152 B.n118 VSUBS 0.007092f
C153 B.n119 VSUBS 0.007092f
C154 B.n120 VSUBS 0.007092f
C155 B.n121 VSUBS 0.007092f
C156 B.n122 VSUBS 0.007092f
C157 B.n123 VSUBS 0.007092f
C158 B.n124 VSUBS 0.007092f
C159 B.n125 VSUBS 0.007092f
C160 B.n126 VSUBS 0.007092f
C161 B.n127 VSUBS 0.007092f
C162 B.n128 VSUBS 0.007092f
C163 B.n129 VSUBS 0.007092f
C164 B.n130 VSUBS 0.007092f
C165 B.n131 VSUBS 0.007092f
C166 B.n132 VSUBS 0.007092f
C167 B.n133 VSUBS 0.007092f
C168 B.n134 VSUBS 0.007092f
C169 B.n135 VSUBS 0.007092f
C170 B.n136 VSUBS 0.007092f
C171 B.n137 VSUBS 0.007092f
C172 B.n138 VSUBS 0.007092f
C173 B.n139 VSUBS 0.007092f
C174 B.n140 VSUBS 0.007092f
C175 B.n141 VSUBS 0.007092f
C176 B.n142 VSUBS 0.007092f
C177 B.n143 VSUBS 0.007092f
C178 B.n144 VSUBS 0.007092f
C179 B.n145 VSUBS 0.007092f
C180 B.n146 VSUBS 0.007092f
C181 B.n147 VSUBS 0.007092f
C182 B.n148 VSUBS 0.007092f
C183 B.n149 VSUBS 0.007092f
C184 B.n150 VSUBS 0.007092f
C185 B.n151 VSUBS 0.007092f
C186 B.n152 VSUBS 0.007092f
C187 B.n153 VSUBS 0.007092f
C188 B.n154 VSUBS 0.007092f
C189 B.n155 VSUBS 0.007092f
C190 B.n156 VSUBS 0.007092f
C191 B.n157 VSUBS 0.017204f
C192 B.n158 VSUBS 0.007092f
C193 B.n159 VSUBS 0.007092f
C194 B.n160 VSUBS 0.007092f
C195 B.n161 VSUBS 0.007092f
C196 B.n162 VSUBS 0.007092f
C197 B.n163 VSUBS 0.007092f
C198 B.n164 VSUBS 0.007092f
C199 B.n165 VSUBS 0.007092f
C200 B.n166 VSUBS 0.007092f
C201 B.n167 VSUBS 0.007092f
C202 B.n168 VSUBS 0.007092f
C203 B.n169 VSUBS 0.007092f
C204 B.n170 VSUBS 0.007092f
C205 B.n171 VSUBS 0.007092f
C206 B.n172 VSUBS 0.007092f
C207 B.n173 VSUBS 0.007092f
C208 B.n174 VSUBS 0.007092f
C209 B.n175 VSUBS 0.007092f
C210 B.n176 VSUBS 0.007092f
C211 B.n177 VSUBS 0.007092f
C212 B.n178 VSUBS 0.007092f
C213 B.n179 VSUBS 0.007092f
C214 B.n180 VSUBS 0.007092f
C215 B.n181 VSUBS 0.007092f
C216 B.n182 VSUBS 0.007092f
C217 B.n183 VSUBS 0.007092f
C218 B.n184 VSUBS 0.007092f
C219 B.n185 VSUBS 0.007092f
C220 B.n186 VSUBS 0.007092f
C221 B.n187 VSUBS 0.007092f
C222 B.n188 VSUBS 0.007092f
C223 B.t11 VSUBS 0.381287f
C224 B.t10 VSUBS 0.418461f
C225 B.t9 VSUBS 2.48169f
C226 B.n189 VSUBS 0.64803f
C227 B.n190 VSUBS 0.346402f
C228 B.n191 VSUBS 0.007092f
C229 B.n192 VSUBS 0.007092f
C230 B.n193 VSUBS 0.007092f
C231 B.n194 VSUBS 0.007092f
C232 B.n195 VSUBS 0.003963f
C233 B.n196 VSUBS 0.007092f
C234 B.n197 VSUBS 0.007092f
C235 B.n198 VSUBS 0.007092f
C236 B.n199 VSUBS 0.007092f
C237 B.n200 VSUBS 0.007092f
C238 B.n201 VSUBS 0.007092f
C239 B.n202 VSUBS 0.007092f
C240 B.n203 VSUBS 0.007092f
C241 B.n204 VSUBS 0.007092f
C242 B.n205 VSUBS 0.007092f
C243 B.n206 VSUBS 0.007092f
C244 B.n207 VSUBS 0.007092f
C245 B.n208 VSUBS 0.007092f
C246 B.n209 VSUBS 0.007092f
C247 B.n210 VSUBS 0.007092f
C248 B.n211 VSUBS 0.007092f
C249 B.n212 VSUBS 0.007092f
C250 B.n213 VSUBS 0.007092f
C251 B.n214 VSUBS 0.007092f
C252 B.n215 VSUBS 0.007092f
C253 B.n216 VSUBS 0.007092f
C254 B.n217 VSUBS 0.007092f
C255 B.n218 VSUBS 0.007092f
C256 B.n219 VSUBS 0.007092f
C257 B.n220 VSUBS 0.007092f
C258 B.n221 VSUBS 0.007092f
C259 B.n222 VSUBS 0.007092f
C260 B.n223 VSUBS 0.007092f
C261 B.n224 VSUBS 0.007092f
C262 B.n225 VSUBS 0.007092f
C263 B.n226 VSUBS 0.017002f
C264 B.n227 VSUBS 0.007092f
C265 B.n228 VSUBS 0.007092f
C266 B.n229 VSUBS 0.007092f
C267 B.n230 VSUBS 0.007092f
C268 B.n231 VSUBS 0.007092f
C269 B.n232 VSUBS 0.007092f
C270 B.n233 VSUBS 0.007092f
C271 B.n234 VSUBS 0.007092f
C272 B.n235 VSUBS 0.007092f
C273 B.n236 VSUBS 0.007092f
C274 B.n237 VSUBS 0.007092f
C275 B.n238 VSUBS 0.007092f
C276 B.n239 VSUBS 0.007092f
C277 B.n240 VSUBS 0.007092f
C278 B.n241 VSUBS 0.007092f
C279 B.n242 VSUBS 0.007092f
C280 B.n243 VSUBS 0.007092f
C281 B.n244 VSUBS 0.007092f
C282 B.n245 VSUBS 0.007092f
C283 B.n246 VSUBS 0.007092f
C284 B.n247 VSUBS 0.007092f
C285 B.n248 VSUBS 0.007092f
C286 B.n249 VSUBS 0.007092f
C287 B.n250 VSUBS 0.007092f
C288 B.n251 VSUBS 0.007092f
C289 B.n252 VSUBS 0.007092f
C290 B.n253 VSUBS 0.007092f
C291 B.n254 VSUBS 0.007092f
C292 B.n255 VSUBS 0.007092f
C293 B.n256 VSUBS 0.007092f
C294 B.n257 VSUBS 0.007092f
C295 B.n258 VSUBS 0.007092f
C296 B.n259 VSUBS 0.007092f
C297 B.n260 VSUBS 0.007092f
C298 B.n261 VSUBS 0.007092f
C299 B.n262 VSUBS 0.007092f
C300 B.n263 VSUBS 0.007092f
C301 B.n264 VSUBS 0.007092f
C302 B.n265 VSUBS 0.007092f
C303 B.n266 VSUBS 0.007092f
C304 B.n267 VSUBS 0.007092f
C305 B.n268 VSUBS 0.007092f
C306 B.n269 VSUBS 0.007092f
C307 B.n270 VSUBS 0.007092f
C308 B.n271 VSUBS 0.007092f
C309 B.n272 VSUBS 0.007092f
C310 B.n273 VSUBS 0.007092f
C311 B.n274 VSUBS 0.007092f
C312 B.n275 VSUBS 0.007092f
C313 B.n276 VSUBS 0.007092f
C314 B.n277 VSUBS 0.007092f
C315 B.n278 VSUBS 0.007092f
C316 B.n279 VSUBS 0.007092f
C317 B.n280 VSUBS 0.007092f
C318 B.n281 VSUBS 0.007092f
C319 B.n282 VSUBS 0.007092f
C320 B.n283 VSUBS 0.007092f
C321 B.n284 VSUBS 0.007092f
C322 B.n285 VSUBS 0.007092f
C323 B.n286 VSUBS 0.007092f
C324 B.n287 VSUBS 0.007092f
C325 B.n288 VSUBS 0.007092f
C326 B.n289 VSUBS 0.007092f
C327 B.n290 VSUBS 0.007092f
C328 B.n291 VSUBS 0.007092f
C329 B.n292 VSUBS 0.007092f
C330 B.n293 VSUBS 0.007092f
C331 B.n294 VSUBS 0.007092f
C332 B.n295 VSUBS 0.007092f
C333 B.n296 VSUBS 0.007092f
C334 B.n297 VSUBS 0.007092f
C335 B.n298 VSUBS 0.007092f
C336 B.n299 VSUBS 0.007092f
C337 B.n300 VSUBS 0.007092f
C338 B.n301 VSUBS 0.007092f
C339 B.n302 VSUBS 0.007092f
C340 B.n303 VSUBS 0.007092f
C341 B.n304 VSUBS 0.007092f
C342 B.n305 VSUBS 0.007092f
C343 B.n306 VSUBS 0.007092f
C344 B.n307 VSUBS 0.007092f
C345 B.n308 VSUBS 0.007092f
C346 B.n309 VSUBS 0.007092f
C347 B.n310 VSUBS 0.007092f
C348 B.n311 VSUBS 0.007092f
C349 B.n312 VSUBS 0.007092f
C350 B.n313 VSUBS 0.007092f
C351 B.n314 VSUBS 0.007092f
C352 B.n315 VSUBS 0.007092f
C353 B.n316 VSUBS 0.007092f
C354 B.n317 VSUBS 0.007092f
C355 B.n318 VSUBS 0.007092f
C356 B.n319 VSUBS 0.007092f
C357 B.n320 VSUBS 0.007092f
C358 B.n321 VSUBS 0.007092f
C359 B.n322 VSUBS 0.007092f
C360 B.n323 VSUBS 0.007092f
C361 B.n324 VSUBS 0.007092f
C362 B.n325 VSUBS 0.007092f
C363 B.n326 VSUBS 0.007092f
C364 B.n327 VSUBS 0.007092f
C365 B.n328 VSUBS 0.007092f
C366 B.n329 VSUBS 0.007092f
C367 B.n330 VSUBS 0.007092f
C368 B.n331 VSUBS 0.007092f
C369 B.n332 VSUBS 0.007092f
C370 B.n333 VSUBS 0.016373f
C371 B.n334 VSUBS 0.016373f
C372 B.n335 VSUBS 0.017002f
C373 B.n336 VSUBS 0.007092f
C374 B.n337 VSUBS 0.007092f
C375 B.n338 VSUBS 0.007092f
C376 B.n339 VSUBS 0.007092f
C377 B.n340 VSUBS 0.007092f
C378 B.n341 VSUBS 0.007092f
C379 B.n342 VSUBS 0.007092f
C380 B.n343 VSUBS 0.007092f
C381 B.n344 VSUBS 0.007092f
C382 B.n345 VSUBS 0.007092f
C383 B.n346 VSUBS 0.007092f
C384 B.n347 VSUBS 0.007092f
C385 B.n348 VSUBS 0.007092f
C386 B.n349 VSUBS 0.007092f
C387 B.n350 VSUBS 0.007092f
C388 B.n351 VSUBS 0.007092f
C389 B.n352 VSUBS 0.007092f
C390 B.n353 VSUBS 0.007092f
C391 B.n354 VSUBS 0.007092f
C392 B.n355 VSUBS 0.007092f
C393 B.n356 VSUBS 0.007092f
C394 B.n357 VSUBS 0.007092f
C395 B.n358 VSUBS 0.007092f
C396 B.n359 VSUBS 0.007092f
C397 B.n360 VSUBS 0.007092f
C398 B.n361 VSUBS 0.007092f
C399 B.n362 VSUBS 0.007092f
C400 B.n363 VSUBS 0.007092f
C401 B.n364 VSUBS 0.007092f
C402 B.n365 VSUBS 0.007092f
C403 B.n366 VSUBS 0.007092f
C404 B.n367 VSUBS 0.007092f
C405 B.n368 VSUBS 0.007092f
C406 B.n369 VSUBS 0.007092f
C407 B.n370 VSUBS 0.007092f
C408 B.n371 VSUBS 0.007092f
C409 B.n372 VSUBS 0.007092f
C410 B.n373 VSUBS 0.007092f
C411 B.n374 VSUBS 0.007092f
C412 B.n375 VSUBS 0.007092f
C413 B.n376 VSUBS 0.007092f
C414 B.n377 VSUBS 0.007092f
C415 B.n378 VSUBS 0.007092f
C416 B.n379 VSUBS 0.007092f
C417 B.n380 VSUBS 0.007092f
C418 B.n381 VSUBS 0.007092f
C419 B.n382 VSUBS 0.007092f
C420 B.n383 VSUBS 0.007092f
C421 B.n384 VSUBS 0.007092f
C422 B.n385 VSUBS 0.007092f
C423 B.n386 VSUBS 0.007092f
C424 B.n387 VSUBS 0.007092f
C425 B.n388 VSUBS 0.007092f
C426 B.n389 VSUBS 0.007092f
C427 B.n390 VSUBS 0.007092f
C428 B.n391 VSUBS 0.007092f
C429 B.n392 VSUBS 0.007092f
C430 B.n393 VSUBS 0.007092f
C431 B.n394 VSUBS 0.007092f
C432 B.n395 VSUBS 0.007092f
C433 B.n396 VSUBS 0.007092f
C434 B.n397 VSUBS 0.007092f
C435 B.n398 VSUBS 0.007092f
C436 B.n399 VSUBS 0.007092f
C437 B.n400 VSUBS 0.007092f
C438 B.n401 VSUBS 0.007092f
C439 B.n402 VSUBS 0.007092f
C440 B.n403 VSUBS 0.007092f
C441 B.n404 VSUBS 0.007092f
C442 B.n405 VSUBS 0.007092f
C443 B.n406 VSUBS 0.007092f
C444 B.n407 VSUBS 0.007092f
C445 B.n408 VSUBS 0.007092f
C446 B.n409 VSUBS 0.007092f
C447 B.n410 VSUBS 0.007092f
C448 B.n411 VSUBS 0.007092f
C449 B.n412 VSUBS 0.007092f
C450 B.n413 VSUBS 0.007092f
C451 B.n414 VSUBS 0.007092f
C452 B.n415 VSUBS 0.007092f
C453 B.n416 VSUBS 0.007092f
C454 B.n417 VSUBS 0.007092f
C455 B.n418 VSUBS 0.007092f
C456 B.n419 VSUBS 0.007092f
C457 B.n420 VSUBS 0.007092f
C458 B.n421 VSUBS 0.007092f
C459 B.n422 VSUBS 0.007092f
C460 B.n423 VSUBS 0.007092f
C461 B.n424 VSUBS 0.007092f
C462 B.n425 VSUBS 0.007092f
C463 B.t8 VSUBS 0.381283f
C464 B.t7 VSUBS 0.418458f
C465 B.t6 VSUBS 2.48169f
C466 B.n426 VSUBS 0.648033f
C467 B.n427 VSUBS 0.346405f
C468 B.n428 VSUBS 0.016432f
C469 B.n429 VSUBS 0.006675f
C470 B.n430 VSUBS 0.007092f
C471 B.n431 VSUBS 0.007092f
C472 B.n432 VSUBS 0.007092f
C473 B.n433 VSUBS 0.007092f
C474 B.n434 VSUBS 0.007092f
C475 B.n435 VSUBS 0.007092f
C476 B.n436 VSUBS 0.007092f
C477 B.n437 VSUBS 0.007092f
C478 B.n438 VSUBS 0.007092f
C479 B.n439 VSUBS 0.007092f
C480 B.n440 VSUBS 0.007092f
C481 B.n441 VSUBS 0.007092f
C482 B.n442 VSUBS 0.007092f
C483 B.n443 VSUBS 0.007092f
C484 B.n444 VSUBS 0.007092f
C485 B.n445 VSUBS 0.003963f
C486 B.n446 VSUBS 0.016432f
C487 B.n447 VSUBS 0.006675f
C488 B.n448 VSUBS 0.007092f
C489 B.n449 VSUBS 0.007092f
C490 B.n450 VSUBS 0.007092f
C491 B.n451 VSUBS 0.007092f
C492 B.n452 VSUBS 0.007092f
C493 B.n453 VSUBS 0.007092f
C494 B.n454 VSUBS 0.007092f
C495 B.n455 VSUBS 0.007092f
C496 B.n456 VSUBS 0.007092f
C497 B.n457 VSUBS 0.007092f
C498 B.n458 VSUBS 0.007092f
C499 B.n459 VSUBS 0.007092f
C500 B.n460 VSUBS 0.007092f
C501 B.n461 VSUBS 0.007092f
C502 B.n462 VSUBS 0.007092f
C503 B.n463 VSUBS 0.007092f
C504 B.n464 VSUBS 0.007092f
C505 B.n465 VSUBS 0.007092f
C506 B.n466 VSUBS 0.007092f
C507 B.n467 VSUBS 0.007092f
C508 B.n468 VSUBS 0.007092f
C509 B.n469 VSUBS 0.007092f
C510 B.n470 VSUBS 0.007092f
C511 B.n471 VSUBS 0.007092f
C512 B.n472 VSUBS 0.007092f
C513 B.n473 VSUBS 0.007092f
C514 B.n474 VSUBS 0.007092f
C515 B.n475 VSUBS 0.007092f
C516 B.n476 VSUBS 0.007092f
C517 B.n477 VSUBS 0.007092f
C518 B.n478 VSUBS 0.007092f
C519 B.n479 VSUBS 0.007092f
C520 B.n480 VSUBS 0.007092f
C521 B.n481 VSUBS 0.007092f
C522 B.n482 VSUBS 0.007092f
C523 B.n483 VSUBS 0.007092f
C524 B.n484 VSUBS 0.007092f
C525 B.n485 VSUBS 0.007092f
C526 B.n486 VSUBS 0.007092f
C527 B.n487 VSUBS 0.007092f
C528 B.n488 VSUBS 0.007092f
C529 B.n489 VSUBS 0.007092f
C530 B.n490 VSUBS 0.007092f
C531 B.n491 VSUBS 0.007092f
C532 B.n492 VSUBS 0.007092f
C533 B.n493 VSUBS 0.007092f
C534 B.n494 VSUBS 0.007092f
C535 B.n495 VSUBS 0.007092f
C536 B.n496 VSUBS 0.007092f
C537 B.n497 VSUBS 0.007092f
C538 B.n498 VSUBS 0.007092f
C539 B.n499 VSUBS 0.007092f
C540 B.n500 VSUBS 0.007092f
C541 B.n501 VSUBS 0.007092f
C542 B.n502 VSUBS 0.007092f
C543 B.n503 VSUBS 0.007092f
C544 B.n504 VSUBS 0.007092f
C545 B.n505 VSUBS 0.007092f
C546 B.n506 VSUBS 0.007092f
C547 B.n507 VSUBS 0.007092f
C548 B.n508 VSUBS 0.007092f
C549 B.n509 VSUBS 0.007092f
C550 B.n510 VSUBS 0.007092f
C551 B.n511 VSUBS 0.007092f
C552 B.n512 VSUBS 0.007092f
C553 B.n513 VSUBS 0.007092f
C554 B.n514 VSUBS 0.007092f
C555 B.n515 VSUBS 0.007092f
C556 B.n516 VSUBS 0.007092f
C557 B.n517 VSUBS 0.007092f
C558 B.n518 VSUBS 0.007092f
C559 B.n519 VSUBS 0.007092f
C560 B.n520 VSUBS 0.007092f
C561 B.n521 VSUBS 0.007092f
C562 B.n522 VSUBS 0.007092f
C563 B.n523 VSUBS 0.007092f
C564 B.n524 VSUBS 0.007092f
C565 B.n525 VSUBS 0.007092f
C566 B.n526 VSUBS 0.007092f
C567 B.n527 VSUBS 0.007092f
C568 B.n528 VSUBS 0.007092f
C569 B.n529 VSUBS 0.007092f
C570 B.n530 VSUBS 0.007092f
C571 B.n531 VSUBS 0.007092f
C572 B.n532 VSUBS 0.007092f
C573 B.n533 VSUBS 0.007092f
C574 B.n534 VSUBS 0.007092f
C575 B.n535 VSUBS 0.007092f
C576 B.n536 VSUBS 0.007092f
C577 B.n537 VSUBS 0.007092f
C578 B.n538 VSUBS 0.016171f
C579 B.n539 VSUBS 0.017002f
C580 B.n540 VSUBS 0.016373f
C581 B.n541 VSUBS 0.007092f
C582 B.n542 VSUBS 0.007092f
C583 B.n543 VSUBS 0.007092f
C584 B.n544 VSUBS 0.007092f
C585 B.n545 VSUBS 0.007092f
C586 B.n546 VSUBS 0.007092f
C587 B.n547 VSUBS 0.007092f
C588 B.n548 VSUBS 0.007092f
C589 B.n549 VSUBS 0.007092f
C590 B.n550 VSUBS 0.007092f
C591 B.n551 VSUBS 0.007092f
C592 B.n552 VSUBS 0.007092f
C593 B.n553 VSUBS 0.007092f
C594 B.n554 VSUBS 0.007092f
C595 B.n555 VSUBS 0.007092f
C596 B.n556 VSUBS 0.007092f
C597 B.n557 VSUBS 0.007092f
C598 B.n558 VSUBS 0.007092f
C599 B.n559 VSUBS 0.007092f
C600 B.n560 VSUBS 0.007092f
C601 B.n561 VSUBS 0.007092f
C602 B.n562 VSUBS 0.007092f
C603 B.n563 VSUBS 0.007092f
C604 B.n564 VSUBS 0.007092f
C605 B.n565 VSUBS 0.007092f
C606 B.n566 VSUBS 0.007092f
C607 B.n567 VSUBS 0.007092f
C608 B.n568 VSUBS 0.007092f
C609 B.n569 VSUBS 0.007092f
C610 B.n570 VSUBS 0.007092f
C611 B.n571 VSUBS 0.007092f
C612 B.n572 VSUBS 0.007092f
C613 B.n573 VSUBS 0.007092f
C614 B.n574 VSUBS 0.007092f
C615 B.n575 VSUBS 0.007092f
C616 B.n576 VSUBS 0.007092f
C617 B.n577 VSUBS 0.007092f
C618 B.n578 VSUBS 0.007092f
C619 B.n579 VSUBS 0.007092f
C620 B.n580 VSUBS 0.007092f
C621 B.n581 VSUBS 0.007092f
C622 B.n582 VSUBS 0.007092f
C623 B.n583 VSUBS 0.007092f
C624 B.n584 VSUBS 0.007092f
C625 B.n585 VSUBS 0.007092f
C626 B.n586 VSUBS 0.007092f
C627 B.n587 VSUBS 0.007092f
C628 B.n588 VSUBS 0.007092f
C629 B.n589 VSUBS 0.007092f
C630 B.n590 VSUBS 0.007092f
C631 B.n591 VSUBS 0.007092f
C632 B.n592 VSUBS 0.007092f
C633 B.n593 VSUBS 0.007092f
C634 B.n594 VSUBS 0.007092f
C635 B.n595 VSUBS 0.007092f
C636 B.n596 VSUBS 0.007092f
C637 B.n597 VSUBS 0.007092f
C638 B.n598 VSUBS 0.007092f
C639 B.n599 VSUBS 0.007092f
C640 B.n600 VSUBS 0.007092f
C641 B.n601 VSUBS 0.007092f
C642 B.n602 VSUBS 0.007092f
C643 B.n603 VSUBS 0.007092f
C644 B.n604 VSUBS 0.007092f
C645 B.n605 VSUBS 0.007092f
C646 B.n606 VSUBS 0.007092f
C647 B.n607 VSUBS 0.007092f
C648 B.n608 VSUBS 0.007092f
C649 B.n609 VSUBS 0.007092f
C650 B.n610 VSUBS 0.007092f
C651 B.n611 VSUBS 0.007092f
C652 B.n612 VSUBS 0.007092f
C653 B.n613 VSUBS 0.007092f
C654 B.n614 VSUBS 0.007092f
C655 B.n615 VSUBS 0.007092f
C656 B.n616 VSUBS 0.007092f
C657 B.n617 VSUBS 0.007092f
C658 B.n618 VSUBS 0.007092f
C659 B.n619 VSUBS 0.007092f
C660 B.n620 VSUBS 0.007092f
C661 B.n621 VSUBS 0.007092f
C662 B.n622 VSUBS 0.007092f
C663 B.n623 VSUBS 0.007092f
C664 B.n624 VSUBS 0.007092f
C665 B.n625 VSUBS 0.007092f
C666 B.n626 VSUBS 0.007092f
C667 B.n627 VSUBS 0.007092f
C668 B.n628 VSUBS 0.007092f
C669 B.n629 VSUBS 0.007092f
C670 B.n630 VSUBS 0.007092f
C671 B.n631 VSUBS 0.007092f
C672 B.n632 VSUBS 0.007092f
C673 B.n633 VSUBS 0.007092f
C674 B.n634 VSUBS 0.007092f
C675 B.n635 VSUBS 0.007092f
C676 B.n636 VSUBS 0.007092f
C677 B.n637 VSUBS 0.007092f
C678 B.n638 VSUBS 0.007092f
C679 B.n639 VSUBS 0.007092f
C680 B.n640 VSUBS 0.007092f
C681 B.n641 VSUBS 0.007092f
C682 B.n642 VSUBS 0.007092f
C683 B.n643 VSUBS 0.007092f
C684 B.n644 VSUBS 0.007092f
C685 B.n645 VSUBS 0.007092f
C686 B.n646 VSUBS 0.007092f
C687 B.n647 VSUBS 0.007092f
C688 B.n648 VSUBS 0.007092f
C689 B.n649 VSUBS 0.007092f
C690 B.n650 VSUBS 0.007092f
C691 B.n651 VSUBS 0.007092f
C692 B.n652 VSUBS 0.007092f
C693 B.n653 VSUBS 0.007092f
C694 B.n654 VSUBS 0.007092f
C695 B.n655 VSUBS 0.007092f
C696 B.n656 VSUBS 0.007092f
C697 B.n657 VSUBS 0.007092f
C698 B.n658 VSUBS 0.007092f
C699 B.n659 VSUBS 0.007092f
C700 B.n660 VSUBS 0.007092f
C701 B.n661 VSUBS 0.007092f
C702 B.n662 VSUBS 0.007092f
C703 B.n663 VSUBS 0.007092f
C704 B.n664 VSUBS 0.007092f
C705 B.n665 VSUBS 0.007092f
C706 B.n666 VSUBS 0.007092f
C707 B.n667 VSUBS 0.007092f
C708 B.n668 VSUBS 0.007092f
C709 B.n669 VSUBS 0.007092f
C710 B.n670 VSUBS 0.007092f
C711 B.n671 VSUBS 0.007092f
C712 B.n672 VSUBS 0.007092f
C713 B.n673 VSUBS 0.007092f
C714 B.n674 VSUBS 0.007092f
C715 B.n675 VSUBS 0.007092f
C716 B.n676 VSUBS 0.007092f
C717 B.n677 VSUBS 0.007092f
C718 B.n678 VSUBS 0.007092f
C719 B.n679 VSUBS 0.007092f
C720 B.n680 VSUBS 0.007092f
C721 B.n681 VSUBS 0.007092f
C722 B.n682 VSUBS 0.007092f
C723 B.n683 VSUBS 0.007092f
C724 B.n684 VSUBS 0.007092f
C725 B.n685 VSUBS 0.007092f
C726 B.n686 VSUBS 0.007092f
C727 B.n687 VSUBS 0.007092f
C728 B.n688 VSUBS 0.007092f
C729 B.n689 VSUBS 0.007092f
C730 B.n690 VSUBS 0.007092f
C731 B.n691 VSUBS 0.007092f
C732 B.n692 VSUBS 0.007092f
C733 B.n693 VSUBS 0.007092f
C734 B.n694 VSUBS 0.007092f
C735 B.n695 VSUBS 0.007092f
C736 B.n696 VSUBS 0.007092f
C737 B.n697 VSUBS 0.007092f
C738 B.n698 VSUBS 0.007092f
C739 B.n699 VSUBS 0.007092f
C740 B.n700 VSUBS 0.007092f
C741 B.n701 VSUBS 0.007092f
C742 B.n702 VSUBS 0.007092f
C743 B.n703 VSUBS 0.007092f
C744 B.n704 VSUBS 0.007092f
C745 B.n705 VSUBS 0.007092f
C746 B.n706 VSUBS 0.016373f
C747 B.n707 VSUBS 0.016373f
C748 B.n708 VSUBS 0.017002f
C749 B.n709 VSUBS 0.007092f
C750 B.n710 VSUBS 0.007092f
C751 B.n711 VSUBS 0.007092f
C752 B.n712 VSUBS 0.007092f
C753 B.n713 VSUBS 0.007092f
C754 B.n714 VSUBS 0.007092f
C755 B.n715 VSUBS 0.007092f
C756 B.n716 VSUBS 0.007092f
C757 B.n717 VSUBS 0.007092f
C758 B.n718 VSUBS 0.007092f
C759 B.n719 VSUBS 0.007092f
C760 B.n720 VSUBS 0.007092f
C761 B.n721 VSUBS 0.007092f
C762 B.n722 VSUBS 0.007092f
C763 B.n723 VSUBS 0.007092f
C764 B.n724 VSUBS 0.007092f
C765 B.n725 VSUBS 0.007092f
C766 B.n726 VSUBS 0.007092f
C767 B.n727 VSUBS 0.007092f
C768 B.n728 VSUBS 0.007092f
C769 B.n729 VSUBS 0.007092f
C770 B.n730 VSUBS 0.007092f
C771 B.n731 VSUBS 0.007092f
C772 B.n732 VSUBS 0.007092f
C773 B.n733 VSUBS 0.007092f
C774 B.n734 VSUBS 0.007092f
C775 B.n735 VSUBS 0.007092f
C776 B.n736 VSUBS 0.007092f
C777 B.n737 VSUBS 0.007092f
C778 B.n738 VSUBS 0.007092f
C779 B.n739 VSUBS 0.007092f
C780 B.n740 VSUBS 0.007092f
C781 B.n741 VSUBS 0.007092f
C782 B.n742 VSUBS 0.007092f
C783 B.n743 VSUBS 0.007092f
C784 B.n744 VSUBS 0.007092f
C785 B.n745 VSUBS 0.007092f
C786 B.n746 VSUBS 0.007092f
C787 B.n747 VSUBS 0.007092f
C788 B.n748 VSUBS 0.007092f
C789 B.n749 VSUBS 0.007092f
C790 B.n750 VSUBS 0.007092f
C791 B.n751 VSUBS 0.007092f
C792 B.n752 VSUBS 0.007092f
C793 B.n753 VSUBS 0.007092f
C794 B.n754 VSUBS 0.007092f
C795 B.n755 VSUBS 0.007092f
C796 B.n756 VSUBS 0.007092f
C797 B.n757 VSUBS 0.007092f
C798 B.n758 VSUBS 0.007092f
C799 B.n759 VSUBS 0.007092f
C800 B.n760 VSUBS 0.007092f
C801 B.n761 VSUBS 0.007092f
C802 B.n762 VSUBS 0.007092f
C803 B.n763 VSUBS 0.007092f
C804 B.n764 VSUBS 0.007092f
C805 B.n765 VSUBS 0.007092f
C806 B.n766 VSUBS 0.007092f
C807 B.n767 VSUBS 0.007092f
C808 B.n768 VSUBS 0.007092f
C809 B.n769 VSUBS 0.007092f
C810 B.n770 VSUBS 0.007092f
C811 B.n771 VSUBS 0.007092f
C812 B.n772 VSUBS 0.007092f
C813 B.n773 VSUBS 0.007092f
C814 B.n774 VSUBS 0.007092f
C815 B.n775 VSUBS 0.007092f
C816 B.n776 VSUBS 0.007092f
C817 B.n777 VSUBS 0.007092f
C818 B.n778 VSUBS 0.007092f
C819 B.n779 VSUBS 0.007092f
C820 B.n780 VSUBS 0.007092f
C821 B.n781 VSUBS 0.007092f
C822 B.n782 VSUBS 0.007092f
C823 B.n783 VSUBS 0.007092f
C824 B.n784 VSUBS 0.007092f
C825 B.n785 VSUBS 0.007092f
C826 B.n786 VSUBS 0.007092f
C827 B.n787 VSUBS 0.007092f
C828 B.n788 VSUBS 0.007092f
C829 B.n789 VSUBS 0.007092f
C830 B.n790 VSUBS 0.007092f
C831 B.n791 VSUBS 0.007092f
C832 B.n792 VSUBS 0.007092f
C833 B.n793 VSUBS 0.007092f
C834 B.n794 VSUBS 0.007092f
C835 B.n795 VSUBS 0.007092f
C836 B.n796 VSUBS 0.007092f
C837 B.n797 VSUBS 0.007092f
C838 B.n798 VSUBS 0.007092f
C839 B.n799 VSUBS 0.007092f
C840 B.n800 VSUBS 0.006675f
C841 B.n801 VSUBS 0.016432f
C842 B.n802 VSUBS 0.003963f
C843 B.n803 VSUBS 0.007092f
C844 B.n804 VSUBS 0.007092f
C845 B.n805 VSUBS 0.007092f
C846 B.n806 VSUBS 0.007092f
C847 B.n807 VSUBS 0.007092f
C848 B.n808 VSUBS 0.007092f
C849 B.n809 VSUBS 0.007092f
C850 B.n810 VSUBS 0.007092f
C851 B.n811 VSUBS 0.007092f
C852 B.n812 VSUBS 0.007092f
C853 B.n813 VSUBS 0.007092f
C854 B.n814 VSUBS 0.007092f
C855 B.n815 VSUBS 0.003963f
C856 B.n816 VSUBS 0.007092f
C857 B.n817 VSUBS 0.007092f
C858 B.n818 VSUBS 0.007092f
C859 B.n819 VSUBS 0.007092f
C860 B.n820 VSUBS 0.007092f
C861 B.n821 VSUBS 0.007092f
C862 B.n822 VSUBS 0.007092f
C863 B.n823 VSUBS 0.007092f
C864 B.n824 VSUBS 0.007092f
C865 B.n825 VSUBS 0.007092f
C866 B.n826 VSUBS 0.007092f
C867 B.n827 VSUBS 0.007092f
C868 B.n828 VSUBS 0.007092f
C869 B.n829 VSUBS 0.007092f
C870 B.n830 VSUBS 0.007092f
C871 B.n831 VSUBS 0.007092f
C872 B.n832 VSUBS 0.007092f
C873 B.n833 VSUBS 0.007092f
C874 B.n834 VSUBS 0.007092f
C875 B.n835 VSUBS 0.007092f
C876 B.n836 VSUBS 0.007092f
C877 B.n837 VSUBS 0.007092f
C878 B.n838 VSUBS 0.007092f
C879 B.n839 VSUBS 0.007092f
C880 B.n840 VSUBS 0.007092f
C881 B.n841 VSUBS 0.007092f
C882 B.n842 VSUBS 0.007092f
C883 B.n843 VSUBS 0.007092f
C884 B.n844 VSUBS 0.007092f
C885 B.n845 VSUBS 0.007092f
C886 B.n846 VSUBS 0.007092f
C887 B.n847 VSUBS 0.007092f
C888 B.n848 VSUBS 0.007092f
C889 B.n849 VSUBS 0.007092f
C890 B.n850 VSUBS 0.007092f
C891 B.n851 VSUBS 0.007092f
C892 B.n852 VSUBS 0.007092f
C893 B.n853 VSUBS 0.007092f
C894 B.n854 VSUBS 0.007092f
C895 B.n855 VSUBS 0.007092f
C896 B.n856 VSUBS 0.007092f
C897 B.n857 VSUBS 0.007092f
C898 B.n858 VSUBS 0.007092f
C899 B.n859 VSUBS 0.007092f
C900 B.n860 VSUBS 0.007092f
C901 B.n861 VSUBS 0.007092f
C902 B.n862 VSUBS 0.007092f
C903 B.n863 VSUBS 0.007092f
C904 B.n864 VSUBS 0.007092f
C905 B.n865 VSUBS 0.007092f
C906 B.n866 VSUBS 0.007092f
C907 B.n867 VSUBS 0.007092f
C908 B.n868 VSUBS 0.007092f
C909 B.n869 VSUBS 0.007092f
C910 B.n870 VSUBS 0.007092f
C911 B.n871 VSUBS 0.007092f
C912 B.n872 VSUBS 0.007092f
C913 B.n873 VSUBS 0.007092f
C914 B.n874 VSUBS 0.007092f
C915 B.n875 VSUBS 0.007092f
C916 B.n876 VSUBS 0.007092f
C917 B.n877 VSUBS 0.007092f
C918 B.n878 VSUBS 0.007092f
C919 B.n879 VSUBS 0.007092f
C920 B.n880 VSUBS 0.007092f
C921 B.n881 VSUBS 0.007092f
C922 B.n882 VSUBS 0.007092f
C923 B.n883 VSUBS 0.007092f
C924 B.n884 VSUBS 0.007092f
C925 B.n885 VSUBS 0.007092f
C926 B.n886 VSUBS 0.007092f
C927 B.n887 VSUBS 0.007092f
C928 B.n888 VSUBS 0.007092f
C929 B.n889 VSUBS 0.007092f
C930 B.n890 VSUBS 0.007092f
C931 B.n891 VSUBS 0.007092f
C932 B.n892 VSUBS 0.007092f
C933 B.n893 VSUBS 0.007092f
C934 B.n894 VSUBS 0.007092f
C935 B.n895 VSUBS 0.007092f
C936 B.n896 VSUBS 0.007092f
C937 B.n897 VSUBS 0.007092f
C938 B.n898 VSUBS 0.007092f
C939 B.n899 VSUBS 0.007092f
C940 B.n900 VSUBS 0.007092f
C941 B.n901 VSUBS 0.007092f
C942 B.n902 VSUBS 0.007092f
C943 B.n903 VSUBS 0.007092f
C944 B.n904 VSUBS 0.007092f
C945 B.n905 VSUBS 0.007092f
C946 B.n906 VSUBS 0.007092f
C947 B.n907 VSUBS 0.007092f
C948 B.n908 VSUBS 0.017002f
C949 B.n909 VSUBS 0.017002f
C950 B.n910 VSUBS 0.016373f
C951 B.n911 VSUBS 0.007092f
C952 B.n912 VSUBS 0.007092f
C953 B.n913 VSUBS 0.007092f
C954 B.n914 VSUBS 0.007092f
C955 B.n915 VSUBS 0.007092f
C956 B.n916 VSUBS 0.007092f
C957 B.n917 VSUBS 0.007092f
C958 B.n918 VSUBS 0.007092f
C959 B.n919 VSUBS 0.007092f
C960 B.n920 VSUBS 0.007092f
C961 B.n921 VSUBS 0.007092f
C962 B.n922 VSUBS 0.007092f
C963 B.n923 VSUBS 0.007092f
C964 B.n924 VSUBS 0.007092f
C965 B.n925 VSUBS 0.007092f
C966 B.n926 VSUBS 0.007092f
C967 B.n927 VSUBS 0.007092f
C968 B.n928 VSUBS 0.007092f
C969 B.n929 VSUBS 0.007092f
C970 B.n930 VSUBS 0.007092f
C971 B.n931 VSUBS 0.007092f
C972 B.n932 VSUBS 0.007092f
C973 B.n933 VSUBS 0.007092f
C974 B.n934 VSUBS 0.007092f
C975 B.n935 VSUBS 0.007092f
C976 B.n936 VSUBS 0.007092f
C977 B.n937 VSUBS 0.007092f
C978 B.n938 VSUBS 0.007092f
C979 B.n939 VSUBS 0.007092f
C980 B.n940 VSUBS 0.007092f
C981 B.n941 VSUBS 0.007092f
C982 B.n942 VSUBS 0.007092f
C983 B.n943 VSUBS 0.007092f
C984 B.n944 VSUBS 0.007092f
C985 B.n945 VSUBS 0.007092f
C986 B.n946 VSUBS 0.007092f
C987 B.n947 VSUBS 0.007092f
C988 B.n948 VSUBS 0.007092f
C989 B.n949 VSUBS 0.007092f
C990 B.n950 VSUBS 0.007092f
C991 B.n951 VSUBS 0.007092f
C992 B.n952 VSUBS 0.007092f
C993 B.n953 VSUBS 0.007092f
C994 B.n954 VSUBS 0.007092f
C995 B.n955 VSUBS 0.007092f
C996 B.n956 VSUBS 0.007092f
C997 B.n957 VSUBS 0.007092f
C998 B.n958 VSUBS 0.007092f
C999 B.n959 VSUBS 0.007092f
C1000 B.n960 VSUBS 0.007092f
C1001 B.n961 VSUBS 0.007092f
C1002 B.n962 VSUBS 0.007092f
C1003 B.n963 VSUBS 0.007092f
C1004 B.n964 VSUBS 0.007092f
C1005 B.n965 VSUBS 0.007092f
C1006 B.n966 VSUBS 0.007092f
C1007 B.n967 VSUBS 0.007092f
C1008 B.n968 VSUBS 0.007092f
C1009 B.n969 VSUBS 0.007092f
C1010 B.n970 VSUBS 0.007092f
C1011 B.n971 VSUBS 0.007092f
C1012 B.n972 VSUBS 0.007092f
C1013 B.n973 VSUBS 0.007092f
C1014 B.n974 VSUBS 0.007092f
C1015 B.n975 VSUBS 0.007092f
C1016 B.n976 VSUBS 0.007092f
C1017 B.n977 VSUBS 0.007092f
C1018 B.n978 VSUBS 0.007092f
C1019 B.n979 VSUBS 0.007092f
C1020 B.n980 VSUBS 0.007092f
C1021 B.n981 VSUBS 0.007092f
C1022 B.n982 VSUBS 0.007092f
C1023 B.n983 VSUBS 0.007092f
C1024 B.n984 VSUBS 0.007092f
C1025 B.n985 VSUBS 0.007092f
C1026 B.n986 VSUBS 0.007092f
C1027 B.n987 VSUBS 0.007092f
C1028 B.n988 VSUBS 0.007092f
C1029 B.n989 VSUBS 0.007092f
C1030 B.n990 VSUBS 0.007092f
C1031 B.n991 VSUBS 0.009255f
C1032 B.n992 VSUBS 0.009859f
C1033 B.n993 VSUBS 0.019605f
C1034 VDD2.t0 VSUBS 0.429851f
C1035 VDD2.t1 VSUBS 0.429851f
C1036 VDD2.n0 VSUBS 3.61853f
C1037 VDD2.t7 VSUBS 0.429851f
C1038 VDD2.t5 VSUBS 0.429851f
C1039 VDD2.n1 VSUBS 3.61853f
C1040 VDD2.n2 VSUBS 5.09408f
C1041 VDD2.t6 VSUBS 0.429851f
C1042 VDD2.t2 VSUBS 0.429851f
C1043 VDD2.n3 VSUBS 3.60068f
C1044 VDD2.n4 VSUBS 4.42121f
C1045 VDD2.t4 VSUBS 0.429851f
C1046 VDD2.t3 VSUBS 0.429851f
C1047 VDD2.n5 VSUBS 3.61847f
C1048 VN.n0 VSUBS 0.031904f
C1049 VN.t2 VSUBS 3.66443f
C1050 VN.n1 VSUBS 0.048674f
C1051 VN.n2 VSUBS 0.024199f
C1052 VN.n3 VSUBS 0.029069f
C1053 VN.n4 VSUBS 0.024199f
C1054 VN.n5 VSUBS 0.035327f
C1055 VN.n6 VSUBS 0.256404f
C1056 VN.t6 VSUBS 3.66443f
C1057 VN.t7 VSUBS 3.91393f
C1058 VN.n7 VSUBS 1.302f
C1059 VN.n8 VSUBS 1.34589f
C1060 VN.n9 VSUBS 0.038867f
C1061 VN.n10 VSUBS 0.045102f
C1062 VN.n11 VSUBS 0.024199f
C1063 VN.n12 VSUBS 0.024199f
C1064 VN.n13 VSUBS 0.024199f
C1065 VN.n14 VSUBS 0.035327f
C1066 VN.n15 VSUBS 0.045102f
C1067 VN.t0 VSUBS 3.66443f
C1068 VN.n16 VSUBS 1.26552f
C1069 VN.n17 VSUBS 0.038867f
C1070 VN.n18 VSUBS 0.024199f
C1071 VN.n19 VSUBS 0.024199f
C1072 VN.n20 VSUBS 0.024199f
C1073 VN.n21 VSUBS 0.045102f
C1074 VN.n22 VSUBS 0.047237f
C1075 VN.n23 VSUBS 0.019844f
C1076 VN.n24 VSUBS 0.024199f
C1077 VN.n25 VSUBS 0.024199f
C1078 VN.n26 VSUBS 0.024199f
C1079 VN.n27 VSUBS 0.045102f
C1080 VN.n28 VSUBS 0.026397f
C1081 VN.n29 VSUBS 1.34787f
C1082 VN.n30 VSUBS 0.045443f
C1083 VN.n31 VSUBS 0.031904f
C1084 VN.t1 VSUBS 3.66443f
C1085 VN.n32 VSUBS 0.048674f
C1086 VN.n33 VSUBS 0.024199f
C1087 VN.n34 VSUBS 0.029069f
C1088 VN.n35 VSUBS 0.024199f
C1089 VN.t5 VSUBS 3.66443f
C1090 VN.n36 VSUBS 1.26552f
C1091 VN.n37 VSUBS 0.035327f
C1092 VN.n38 VSUBS 0.256404f
C1093 VN.t3 VSUBS 3.66443f
C1094 VN.t4 VSUBS 3.91393f
C1095 VN.n39 VSUBS 1.302f
C1096 VN.n40 VSUBS 1.34589f
C1097 VN.n41 VSUBS 0.038867f
C1098 VN.n42 VSUBS 0.045102f
C1099 VN.n43 VSUBS 0.024199f
C1100 VN.n44 VSUBS 0.024199f
C1101 VN.n45 VSUBS 0.024199f
C1102 VN.n46 VSUBS 0.035327f
C1103 VN.n47 VSUBS 0.045102f
C1104 VN.n48 VSUBS 0.038867f
C1105 VN.n49 VSUBS 0.024199f
C1106 VN.n50 VSUBS 0.024199f
C1107 VN.n51 VSUBS 0.024199f
C1108 VN.n52 VSUBS 0.045102f
C1109 VN.n53 VSUBS 0.047237f
C1110 VN.n54 VSUBS 0.019844f
C1111 VN.n55 VSUBS 0.024199f
C1112 VN.n56 VSUBS 0.024199f
C1113 VN.n57 VSUBS 0.024199f
C1114 VN.n58 VSUBS 0.045102f
C1115 VN.n59 VSUBS 0.026397f
C1116 VN.n60 VSUBS 1.34787f
C1117 VN.n61 VSUBS 1.66515f
C1118 VDD1.t1 VSUBS 0.401316f
C1119 VDD1.t3 VSUBS 0.401316f
C1120 VDD1.n0 VSUBS 3.37991f
C1121 VDD1.t6 VSUBS 0.401316f
C1122 VDD1.t7 VSUBS 0.401316f
C1123 VDD1.n1 VSUBS 3.37832f
C1124 VDD1.t0 VSUBS 0.401316f
C1125 VDD1.t2 VSUBS 0.401316f
C1126 VDD1.n2 VSUBS 3.37832f
C1127 VDD1.n3 VSUBS 4.81103f
C1128 VDD1.t4 VSUBS 0.401316f
C1129 VDD1.t5 VSUBS 0.401316f
C1130 VDD1.n4 VSUBS 3.36164f
C1131 VDD1.n5 VSUBS 4.16118f
C1132 VTAIL.t2 VSUBS 0.355023f
C1133 VTAIL.t7 VSUBS 0.355023f
C1134 VTAIL.n0 VSUBS 2.82935f
C1135 VTAIL.n1 VSUBS 0.792327f
C1136 VTAIL.n2 VSUBS 0.026943f
C1137 VTAIL.n3 VSUBS 0.023608f
C1138 VTAIL.n4 VSUBS 0.012686f
C1139 VTAIL.n5 VSUBS 0.029985f
C1140 VTAIL.n6 VSUBS 0.013432f
C1141 VTAIL.n7 VSUBS 0.023608f
C1142 VTAIL.n8 VSUBS 0.012686f
C1143 VTAIL.n9 VSUBS 0.029985f
C1144 VTAIL.n10 VSUBS 0.013432f
C1145 VTAIL.n11 VSUBS 0.023608f
C1146 VTAIL.n12 VSUBS 0.012686f
C1147 VTAIL.n13 VSUBS 0.029985f
C1148 VTAIL.n14 VSUBS 0.013432f
C1149 VTAIL.n15 VSUBS 0.023608f
C1150 VTAIL.n16 VSUBS 0.012686f
C1151 VTAIL.n17 VSUBS 0.029985f
C1152 VTAIL.n18 VSUBS 0.013432f
C1153 VTAIL.n19 VSUBS 0.023608f
C1154 VTAIL.n20 VSUBS 0.012686f
C1155 VTAIL.n21 VSUBS 0.029985f
C1156 VTAIL.n22 VSUBS 0.013432f
C1157 VTAIL.n23 VSUBS 0.023608f
C1158 VTAIL.n24 VSUBS 0.012686f
C1159 VTAIL.n25 VSUBS 0.029985f
C1160 VTAIL.n26 VSUBS 0.013432f
C1161 VTAIL.n27 VSUBS 0.023608f
C1162 VTAIL.n28 VSUBS 0.012686f
C1163 VTAIL.n29 VSUBS 0.029985f
C1164 VTAIL.n30 VSUBS 0.013432f
C1165 VTAIL.n31 VSUBS 0.023608f
C1166 VTAIL.n32 VSUBS 0.012686f
C1167 VTAIL.n33 VSUBS 0.029985f
C1168 VTAIL.n34 VSUBS 0.013432f
C1169 VTAIL.n35 VSUBS 0.194481f
C1170 VTAIL.t5 VSUBS 0.064429f
C1171 VTAIL.n36 VSUBS 0.022489f
C1172 VTAIL.n37 VSUBS 0.019075f
C1173 VTAIL.n38 VSUBS 0.012686f
C1174 VTAIL.n39 VSUBS 1.93935f
C1175 VTAIL.n40 VSUBS 0.023608f
C1176 VTAIL.n41 VSUBS 0.012686f
C1177 VTAIL.n42 VSUBS 0.013432f
C1178 VTAIL.n43 VSUBS 0.029985f
C1179 VTAIL.n44 VSUBS 0.029985f
C1180 VTAIL.n45 VSUBS 0.013432f
C1181 VTAIL.n46 VSUBS 0.012686f
C1182 VTAIL.n47 VSUBS 0.023608f
C1183 VTAIL.n48 VSUBS 0.023608f
C1184 VTAIL.n49 VSUBS 0.012686f
C1185 VTAIL.n50 VSUBS 0.013432f
C1186 VTAIL.n51 VSUBS 0.029985f
C1187 VTAIL.n52 VSUBS 0.029985f
C1188 VTAIL.n53 VSUBS 0.013432f
C1189 VTAIL.n54 VSUBS 0.012686f
C1190 VTAIL.n55 VSUBS 0.023608f
C1191 VTAIL.n56 VSUBS 0.023608f
C1192 VTAIL.n57 VSUBS 0.012686f
C1193 VTAIL.n58 VSUBS 0.013432f
C1194 VTAIL.n59 VSUBS 0.029985f
C1195 VTAIL.n60 VSUBS 0.029985f
C1196 VTAIL.n61 VSUBS 0.013432f
C1197 VTAIL.n62 VSUBS 0.012686f
C1198 VTAIL.n63 VSUBS 0.023608f
C1199 VTAIL.n64 VSUBS 0.023608f
C1200 VTAIL.n65 VSUBS 0.012686f
C1201 VTAIL.n66 VSUBS 0.013432f
C1202 VTAIL.n67 VSUBS 0.029985f
C1203 VTAIL.n68 VSUBS 0.029985f
C1204 VTAIL.n69 VSUBS 0.013432f
C1205 VTAIL.n70 VSUBS 0.012686f
C1206 VTAIL.n71 VSUBS 0.023608f
C1207 VTAIL.n72 VSUBS 0.023608f
C1208 VTAIL.n73 VSUBS 0.012686f
C1209 VTAIL.n74 VSUBS 0.013432f
C1210 VTAIL.n75 VSUBS 0.029985f
C1211 VTAIL.n76 VSUBS 0.029985f
C1212 VTAIL.n77 VSUBS 0.029985f
C1213 VTAIL.n78 VSUBS 0.013432f
C1214 VTAIL.n79 VSUBS 0.012686f
C1215 VTAIL.n80 VSUBS 0.023608f
C1216 VTAIL.n81 VSUBS 0.023608f
C1217 VTAIL.n82 VSUBS 0.012686f
C1218 VTAIL.n83 VSUBS 0.013059f
C1219 VTAIL.n84 VSUBS 0.013059f
C1220 VTAIL.n85 VSUBS 0.029985f
C1221 VTAIL.n86 VSUBS 0.029985f
C1222 VTAIL.n87 VSUBS 0.013432f
C1223 VTAIL.n88 VSUBS 0.012686f
C1224 VTAIL.n89 VSUBS 0.023608f
C1225 VTAIL.n90 VSUBS 0.023608f
C1226 VTAIL.n91 VSUBS 0.012686f
C1227 VTAIL.n92 VSUBS 0.013432f
C1228 VTAIL.n93 VSUBS 0.029985f
C1229 VTAIL.n94 VSUBS 0.029985f
C1230 VTAIL.n95 VSUBS 0.013432f
C1231 VTAIL.n96 VSUBS 0.012686f
C1232 VTAIL.n97 VSUBS 0.023608f
C1233 VTAIL.n98 VSUBS 0.023608f
C1234 VTAIL.n99 VSUBS 0.012686f
C1235 VTAIL.n100 VSUBS 0.013432f
C1236 VTAIL.n101 VSUBS 0.029985f
C1237 VTAIL.n102 VSUBS 0.076005f
C1238 VTAIL.n103 VSUBS 0.013432f
C1239 VTAIL.n104 VSUBS 0.012686f
C1240 VTAIL.n105 VSUBS 0.056827f
C1241 VTAIL.n106 VSUBS 0.038442f
C1242 VTAIL.n107 VSUBS 0.268342f
C1243 VTAIL.n108 VSUBS 0.026943f
C1244 VTAIL.n109 VSUBS 0.023608f
C1245 VTAIL.n110 VSUBS 0.012686f
C1246 VTAIL.n111 VSUBS 0.029985f
C1247 VTAIL.n112 VSUBS 0.013432f
C1248 VTAIL.n113 VSUBS 0.023608f
C1249 VTAIL.n114 VSUBS 0.012686f
C1250 VTAIL.n115 VSUBS 0.029985f
C1251 VTAIL.n116 VSUBS 0.013432f
C1252 VTAIL.n117 VSUBS 0.023608f
C1253 VTAIL.n118 VSUBS 0.012686f
C1254 VTAIL.n119 VSUBS 0.029985f
C1255 VTAIL.n120 VSUBS 0.013432f
C1256 VTAIL.n121 VSUBS 0.023608f
C1257 VTAIL.n122 VSUBS 0.012686f
C1258 VTAIL.n123 VSUBS 0.029985f
C1259 VTAIL.n124 VSUBS 0.013432f
C1260 VTAIL.n125 VSUBS 0.023608f
C1261 VTAIL.n126 VSUBS 0.012686f
C1262 VTAIL.n127 VSUBS 0.029985f
C1263 VTAIL.n128 VSUBS 0.013432f
C1264 VTAIL.n129 VSUBS 0.023608f
C1265 VTAIL.n130 VSUBS 0.012686f
C1266 VTAIL.n131 VSUBS 0.029985f
C1267 VTAIL.n132 VSUBS 0.013432f
C1268 VTAIL.n133 VSUBS 0.023608f
C1269 VTAIL.n134 VSUBS 0.012686f
C1270 VTAIL.n135 VSUBS 0.029985f
C1271 VTAIL.n136 VSUBS 0.013432f
C1272 VTAIL.n137 VSUBS 0.023608f
C1273 VTAIL.n138 VSUBS 0.012686f
C1274 VTAIL.n139 VSUBS 0.029985f
C1275 VTAIL.n140 VSUBS 0.013432f
C1276 VTAIL.n141 VSUBS 0.194481f
C1277 VTAIL.t8 VSUBS 0.064429f
C1278 VTAIL.n142 VSUBS 0.022489f
C1279 VTAIL.n143 VSUBS 0.019075f
C1280 VTAIL.n144 VSUBS 0.012686f
C1281 VTAIL.n145 VSUBS 1.93935f
C1282 VTAIL.n146 VSUBS 0.023608f
C1283 VTAIL.n147 VSUBS 0.012686f
C1284 VTAIL.n148 VSUBS 0.013432f
C1285 VTAIL.n149 VSUBS 0.029985f
C1286 VTAIL.n150 VSUBS 0.029985f
C1287 VTAIL.n151 VSUBS 0.013432f
C1288 VTAIL.n152 VSUBS 0.012686f
C1289 VTAIL.n153 VSUBS 0.023608f
C1290 VTAIL.n154 VSUBS 0.023608f
C1291 VTAIL.n155 VSUBS 0.012686f
C1292 VTAIL.n156 VSUBS 0.013432f
C1293 VTAIL.n157 VSUBS 0.029985f
C1294 VTAIL.n158 VSUBS 0.029985f
C1295 VTAIL.n159 VSUBS 0.013432f
C1296 VTAIL.n160 VSUBS 0.012686f
C1297 VTAIL.n161 VSUBS 0.023608f
C1298 VTAIL.n162 VSUBS 0.023608f
C1299 VTAIL.n163 VSUBS 0.012686f
C1300 VTAIL.n164 VSUBS 0.013432f
C1301 VTAIL.n165 VSUBS 0.029985f
C1302 VTAIL.n166 VSUBS 0.029985f
C1303 VTAIL.n167 VSUBS 0.013432f
C1304 VTAIL.n168 VSUBS 0.012686f
C1305 VTAIL.n169 VSUBS 0.023608f
C1306 VTAIL.n170 VSUBS 0.023608f
C1307 VTAIL.n171 VSUBS 0.012686f
C1308 VTAIL.n172 VSUBS 0.013432f
C1309 VTAIL.n173 VSUBS 0.029985f
C1310 VTAIL.n174 VSUBS 0.029985f
C1311 VTAIL.n175 VSUBS 0.013432f
C1312 VTAIL.n176 VSUBS 0.012686f
C1313 VTAIL.n177 VSUBS 0.023608f
C1314 VTAIL.n178 VSUBS 0.023608f
C1315 VTAIL.n179 VSUBS 0.012686f
C1316 VTAIL.n180 VSUBS 0.013432f
C1317 VTAIL.n181 VSUBS 0.029985f
C1318 VTAIL.n182 VSUBS 0.029985f
C1319 VTAIL.n183 VSUBS 0.029985f
C1320 VTAIL.n184 VSUBS 0.013432f
C1321 VTAIL.n185 VSUBS 0.012686f
C1322 VTAIL.n186 VSUBS 0.023608f
C1323 VTAIL.n187 VSUBS 0.023608f
C1324 VTAIL.n188 VSUBS 0.012686f
C1325 VTAIL.n189 VSUBS 0.013059f
C1326 VTAIL.n190 VSUBS 0.013059f
C1327 VTAIL.n191 VSUBS 0.029985f
C1328 VTAIL.n192 VSUBS 0.029985f
C1329 VTAIL.n193 VSUBS 0.013432f
C1330 VTAIL.n194 VSUBS 0.012686f
C1331 VTAIL.n195 VSUBS 0.023608f
C1332 VTAIL.n196 VSUBS 0.023608f
C1333 VTAIL.n197 VSUBS 0.012686f
C1334 VTAIL.n198 VSUBS 0.013432f
C1335 VTAIL.n199 VSUBS 0.029985f
C1336 VTAIL.n200 VSUBS 0.029985f
C1337 VTAIL.n201 VSUBS 0.013432f
C1338 VTAIL.n202 VSUBS 0.012686f
C1339 VTAIL.n203 VSUBS 0.023608f
C1340 VTAIL.n204 VSUBS 0.023608f
C1341 VTAIL.n205 VSUBS 0.012686f
C1342 VTAIL.n206 VSUBS 0.013432f
C1343 VTAIL.n207 VSUBS 0.029985f
C1344 VTAIL.n208 VSUBS 0.076005f
C1345 VTAIL.n209 VSUBS 0.013432f
C1346 VTAIL.n210 VSUBS 0.012686f
C1347 VTAIL.n211 VSUBS 0.056827f
C1348 VTAIL.n212 VSUBS 0.038442f
C1349 VTAIL.n213 VSUBS 0.268342f
C1350 VTAIL.t12 VSUBS 0.355023f
C1351 VTAIL.t15 VSUBS 0.355023f
C1352 VTAIL.n214 VSUBS 2.82935f
C1353 VTAIL.n215 VSUBS 0.999063f
C1354 VTAIL.n216 VSUBS 0.026943f
C1355 VTAIL.n217 VSUBS 0.023608f
C1356 VTAIL.n218 VSUBS 0.012686f
C1357 VTAIL.n219 VSUBS 0.029985f
C1358 VTAIL.n220 VSUBS 0.013432f
C1359 VTAIL.n221 VSUBS 0.023608f
C1360 VTAIL.n222 VSUBS 0.012686f
C1361 VTAIL.n223 VSUBS 0.029985f
C1362 VTAIL.n224 VSUBS 0.013432f
C1363 VTAIL.n225 VSUBS 0.023608f
C1364 VTAIL.n226 VSUBS 0.012686f
C1365 VTAIL.n227 VSUBS 0.029985f
C1366 VTAIL.n228 VSUBS 0.013432f
C1367 VTAIL.n229 VSUBS 0.023608f
C1368 VTAIL.n230 VSUBS 0.012686f
C1369 VTAIL.n231 VSUBS 0.029985f
C1370 VTAIL.n232 VSUBS 0.013432f
C1371 VTAIL.n233 VSUBS 0.023608f
C1372 VTAIL.n234 VSUBS 0.012686f
C1373 VTAIL.n235 VSUBS 0.029985f
C1374 VTAIL.n236 VSUBS 0.013432f
C1375 VTAIL.n237 VSUBS 0.023608f
C1376 VTAIL.n238 VSUBS 0.012686f
C1377 VTAIL.n239 VSUBS 0.029985f
C1378 VTAIL.n240 VSUBS 0.013432f
C1379 VTAIL.n241 VSUBS 0.023608f
C1380 VTAIL.n242 VSUBS 0.012686f
C1381 VTAIL.n243 VSUBS 0.029985f
C1382 VTAIL.n244 VSUBS 0.013432f
C1383 VTAIL.n245 VSUBS 0.023608f
C1384 VTAIL.n246 VSUBS 0.012686f
C1385 VTAIL.n247 VSUBS 0.029985f
C1386 VTAIL.n248 VSUBS 0.013432f
C1387 VTAIL.n249 VSUBS 0.194481f
C1388 VTAIL.t11 VSUBS 0.064429f
C1389 VTAIL.n250 VSUBS 0.022489f
C1390 VTAIL.n251 VSUBS 0.019075f
C1391 VTAIL.n252 VSUBS 0.012686f
C1392 VTAIL.n253 VSUBS 1.93935f
C1393 VTAIL.n254 VSUBS 0.023608f
C1394 VTAIL.n255 VSUBS 0.012686f
C1395 VTAIL.n256 VSUBS 0.013432f
C1396 VTAIL.n257 VSUBS 0.029985f
C1397 VTAIL.n258 VSUBS 0.029985f
C1398 VTAIL.n259 VSUBS 0.013432f
C1399 VTAIL.n260 VSUBS 0.012686f
C1400 VTAIL.n261 VSUBS 0.023608f
C1401 VTAIL.n262 VSUBS 0.023608f
C1402 VTAIL.n263 VSUBS 0.012686f
C1403 VTAIL.n264 VSUBS 0.013432f
C1404 VTAIL.n265 VSUBS 0.029985f
C1405 VTAIL.n266 VSUBS 0.029985f
C1406 VTAIL.n267 VSUBS 0.013432f
C1407 VTAIL.n268 VSUBS 0.012686f
C1408 VTAIL.n269 VSUBS 0.023608f
C1409 VTAIL.n270 VSUBS 0.023608f
C1410 VTAIL.n271 VSUBS 0.012686f
C1411 VTAIL.n272 VSUBS 0.013432f
C1412 VTAIL.n273 VSUBS 0.029985f
C1413 VTAIL.n274 VSUBS 0.029985f
C1414 VTAIL.n275 VSUBS 0.013432f
C1415 VTAIL.n276 VSUBS 0.012686f
C1416 VTAIL.n277 VSUBS 0.023608f
C1417 VTAIL.n278 VSUBS 0.023608f
C1418 VTAIL.n279 VSUBS 0.012686f
C1419 VTAIL.n280 VSUBS 0.013432f
C1420 VTAIL.n281 VSUBS 0.029985f
C1421 VTAIL.n282 VSUBS 0.029985f
C1422 VTAIL.n283 VSUBS 0.013432f
C1423 VTAIL.n284 VSUBS 0.012686f
C1424 VTAIL.n285 VSUBS 0.023608f
C1425 VTAIL.n286 VSUBS 0.023608f
C1426 VTAIL.n287 VSUBS 0.012686f
C1427 VTAIL.n288 VSUBS 0.013432f
C1428 VTAIL.n289 VSUBS 0.029985f
C1429 VTAIL.n290 VSUBS 0.029985f
C1430 VTAIL.n291 VSUBS 0.029985f
C1431 VTAIL.n292 VSUBS 0.013432f
C1432 VTAIL.n293 VSUBS 0.012686f
C1433 VTAIL.n294 VSUBS 0.023608f
C1434 VTAIL.n295 VSUBS 0.023608f
C1435 VTAIL.n296 VSUBS 0.012686f
C1436 VTAIL.n297 VSUBS 0.013059f
C1437 VTAIL.n298 VSUBS 0.013059f
C1438 VTAIL.n299 VSUBS 0.029985f
C1439 VTAIL.n300 VSUBS 0.029985f
C1440 VTAIL.n301 VSUBS 0.013432f
C1441 VTAIL.n302 VSUBS 0.012686f
C1442 VTAIL.n303 VSUBS 0.023608f
C1443 VTAIL.n304 VSUBS 0.023608f
C1444 VTAIL.n305 VSUBS 0.012686f
C1445 VTAIL.n306 VSUBS 0.013432f
C1446 VTAIL.n307 VSUBS 0.029985f
C1447 VTAIL.n308 VSUBS 0.029985f
C1448 VTAIL.n309 VSUBS 0.013432f
C1449 VTAIL.n310 VSUBS 0.012686f
C1450 VTAIL.n311 VSUBS 0.023608f
C1451 VTAIL.n312 VSUBS 0.023608f
C1452 VTAIL.n313 VSUBS 0.012686f
C1453 VTAIL.n314 VSUBS 0.013432f
C1454 VTAIL.n315 VSUBS 0.029985f
C1455 VTAIL.n316 VSUBS 0.076005f
C1456 VTAIL.n317 VSUBS 0.013432f
C1457 VTAIL.n318 VSUBS 0.012686f
C1458 VTAIL.n319 VSUBS 0.056827f
C1459 VTAIL.n320 VSUBS 0.038442f
C1460 VTAIL.n321 VSUBS 2.01242f
C1461 VTAIL.n322 VSUBS 0.026943f
C1462 VTAIL.n323 VSUBS 0.023608f
C1463 VTAIL.n324 VSUBS 0.012686f
C1464 VTAIL.n325 VSUBS 0.029985f
C1465 VTAIL.n326 VSUBS 0.013432f
C1466 VTAIL.n327 VSUBS 0.023608f
C1467 VTAIL.n328 VSUBS 0.012686f
C1468 VTAIL.n329 VSUBS 0.029985f
C1469 VTAIL.n330 VSUBS 0.013432f
C1470 VTAIL.n331 VSUBS 0.023608f
C1471 VTAIL.n332 VSUBS 0.012686f
C1472 VTAIL.n333 VSUBS 0.029985f
C1473 VTAIL.n334 VSUBS 0.013432f
C1474 VTAIL.n335 VSUBS 0.023608f
C1475 VTAIL.n336 VSUBS 0.012686f
C1476 VTAIL.n337 VSUBS 0.029985f
C1477 VTAIL.n338 VSUBS 0.029985f
C1478 VTAIL.n339 VSUBS 0.013432f
C1479 VTAIL.n340 VSUBS 0.023608f
C1480 VTAIL.n341 VSUBS 0.012686f
C1481 VTAIL.n342 VSUBS 0.029985f
C1482 VTAIL.n343 VSUBS 0.013432f
C1483 VTAIL.n344 VSUBS 0.023608f
C1484 VTAIL.n345 VSUBS 0.012686f
C1485 VTAIL.n346 VSUBS 0.029985f
C1486 VTAIL.n347 VSUBS 0.013432f
C1487 VTAIL.n348 VSUBS 0.023608f
C1488 VTAIL.n349 VSUBS 0.012686f
C1489 VTAIL.n350 VSUBS 0.029985f
C1490 VTAIL.n351 VSUBS 0.013432f
C1491 VTAIL.n352 VSUBS 0.023608f
C1492 VTAIL.n353 VSUBS 0.012686f
C1493 VTAIL.n354 VSUBS 0.029985f
C1494 VTAIL.n355 VSUBS 0.013432f
C1495 VTAIL.n356 VSUBS 0.194481f
C1496 VTAIL.t6 VSUBS 0.064429f
C1497 VTAIL.n357 VSUBS 0.022489f
C1498 VTAIL.n358 VSUBS 0.019075f
C1499 VTAIL.n359 VSUBS 0.012686f
C1500 VTAIL.n360 VSUBS 1.93935f
C1501 VTAIL.n361 VSUBS 0.023608f
C1502 VTAIL.n362 VSUBS 0.012686f
C1503 VTAIL.n363 VSUBS 0.013432f
C1504 VTAIL.n364 VSUBS 0.029985f
C1505 VTAIL.n365 VSUBS 0.029985f
C1506 VTAIL.n366 VSUBS 0.013432f
C1507 VTAIL.n367 VSUBS 0.012686f
C1508 VTAIL.n368 VSUBS 0.023608f
C1509 VTAIL.n369 VSUBS 0.023608f
C1510 VTAIL.n370 VSUBS 0.012686f
C1511 VTAIL.n371 VSUBS 0.013432f
C1512 VTAIL.n372 VSUBS 0.029985f
C1513 VTAIL.n373 VSUBS 0.029985f
C1514 VTAIL.n374 VSUBS 0.013432f
C1515 VTAIL.n375 VSUBS 0.012686f
C1516 VTAIL.n376 VSUBS 0.023608f
C1517 VTAIL.n377 VSUBS 0.023608f
C1518 VTAIL.n378 VSUBS 0.012686f
C1519 VTAIL.n379 VSUBS 0.013432f
C1520 VTAIL.n380 VSUBS 0.029985f
C1521 VTAIL.n381 VSUBS 0.029985f
C1522 VTAIL.n382 VSUBS 0.013432f
C1523 VTAIL.n383 VSUBS 0.012686f
C1524 VTAIL.n384 VSUBS 0.023608f
C1525 VTAIL.n385 VSUBS 0.023608f
C1526 VTAIL.n386 VSUBS 0.012686f
C1527 VTAIL.n387 VSUBS 0.013432f
C1528 VTAIL.n388 VSUBS 0.029985f
C1529 VTAIL.n389 VSUBS 0.029985f
C1530 VTAIL.n390 VSUBS 0.013432f
C1531 VTAIL.n391 VSUBS 0.012686f
C1532 VTAIL.n392 VSUBS 0.023608f
C1533 VTAIL.n393 VSUBS 0.023608f
C1534 VTAIL.n394 VSUBS 0.012686f
C1535 VTAIL.n395 VSUBS 0.013432f
C1536 VTAIL.n396 VSUBS 0.029985f
C1537 VTAIL.n397 VSUBS 0.029985f
C1538 VTAIL.n398 VSUBS 0.013432f
C1539 VTAIL.n399 VSUBS 0.012686f
C1540 VTAIL.n400 VSUBS 0.023608f
C1541 VTAIL.n401 VSUBS 0.023608f
C1542 VTAIL.n402 VSUBS 0.012686f
C1543 VTAIL.n403 VSUBS 0.013059f
C1544 VTAIL.n404 VSUBS 0.013059f
C1545 VTAIL.n405 VSUBS 0.029985f
C1546 VTAIL.n406 VSUBS 0.029985f
C1547 VTAIL.n407 VSUBS 0.013432f
C1548 VTAIL.n408 VSUBS 0.012686f
C1549 VTAIL.n409 VSUBS 0.023608f
C1550 VTAIL.n410 VSUBS 0.023608f
C1551 VTAIL.n411 VSUBS 0.012686f
C1552 VTAIL.n412 VSUBS 0.013432f
C1553 VTAIL.n413 VSUBS 0.029985f
C1554 VTAIL.n414 VSUBS 0.029985f
C1555 VTAIL.n415 VSUBS 0.013432f
C1556 VTAIL.n416 VSUBS 0.012686f
C1557 VTAIL.n417 VSUBS 0.023608f
C1558 VTAIL.n418 VSUBS 0.023608f
C1559 VTAIL.n419 VSUBS 0.012686f
C1560 VTAIL.n420 VSUBS 0.013432f
C1561 VTAIL.n421 VSUBS 0.029985f
C1562 VTAIL.n422 VSUBS 0.076005f
C1563 VTAIL.n423 VSUBS 0.013432f
C1564 VTAIL.n424 VSUBS 0.012686f
C1565 VTAIL.n425 VSUBS 0.056827f
C1566 VTAIL.n426 VSUBS 0.038442f
C1567 VTAIL.n427 VSUBS 2.01242f
C1568 VTAIL.t1 VSUBS 0.355023f
C1569 VTAIL.t3 VSUBS 0.355023f
C1570 VTAIL.n428 VSUBS 2.82936f
C1571 VTAIL.n429 VSUBS 0.999054f
C1572 VTAIL.n430 VSUBS 0.026943f
C1573 VTAIL.n431 VSUBS 0.023608f
C1574 VTAIL.n432 VSUBS 0.012686f
C1575 VTAIL.n433 VSUBS 0.029985f
C1576 VTAIL.n434 VSUBS 0.013432f
C1577 VTAIL.n435 VSUBS 0.023608f
C1578 VTAIL.n436 VSUBS 0.012686f
C1579 VTAIL.n437 VSUBS 0.029985f
C1580 VTAIL.n438 VSUBS 0.013432f
C1581 VTAIL.n439 VSUBS 0.023608f
C1582 VTAIL.n440 VSUBS 0.012686f
C1583 VTAIL.n441 VSUBS 0.029985f
C1584 VTAIL.n442 VSUBS 0.013432f
C1585 VTAIL.n443 VSUBS 0.023608f
C1586 VTAIL.n444 VSUBS 0.012686f
C1587 VTAIL.n445 VSUBS 0.029985f
C1588 VTAIL.n446 VSUBS 0.029985f
C1589 VTAIL.n447 VSUBS 0.013432f
C1590 VTAIL.n448 VSUBS 0.023608f
C1591 VTAIL.n449 VSUBS 0.012686f
C1592 VTAIL.n450 VSUBS 0.029985f
C1593 VTAIL.n451 VSUBS 0.013432f
C1594 VTAIL.n452 VSUBS 0.023608f
C1595 VTAIL.n453 VSUBS 0.012686f
C1596 VTAIL.n454 VSUBS 0.029985f
C1597 VTAIL.n455 VSUBS 0.013432f
C1598 VTAIL.n456 VSUBS 0.023608f
C1599 VTAIL.n457 VSUBS 0.012686f
C1600 VTAIL.n458 VSUBS 0.029985f
C1601 VTAIL.n459 VSUBS 0.013432f
C1602 VTAIL.n460 VSUBS 0.023608f
C1603 VTAIL.n461 VSUBS 0.012686f
C1604 VTAIL.n462 VSUBS 0.029985f
C1605 VTAIL.n463 VSUBS 0.013432f
C1606 VTAIL.n464 VSUBS 0.194481f
C1607 VTAIL.t4 VSUBS 0.064429f
C1608 VTAIL.n465 VSUBS 0.022489f
C1609 VTAIL.n466 VSUBS 0.019075f
C1610 VTAIL.n467 VSUBS 0.012686f
C1611 VTAIL.n468 VSUBS 1.93935f
C1612 VTAIL.n469 VSUBS 0.023608f
C1613 VTAIL.n470 VSUBS 0.012686f
C1614 VTAIL.n471 VSUBS 0.013432f
C1615 VTAIL.n472 VSUBS 0.029985f
C1616 VTAIL.n473 VSUBS 0.029985f
C1617 VTAIL.n474 VSUBS 0.013432f
C1618 VTAIL.n475 VSUBS 0.012686f
C1619 VTAIL.n476 VSUBS 0.023608f
C1620 VTAIL.n477 VSUBS 0.023608f
C1621 VTAIL.n478 VSUBS 0.012686f
C1622 VTAIL.n479 VSUBS 0.013432f
C1623 VTAIL.n480 VSUBS 0.029985f
C1624 VTAIL.n481 VSUBS 0.029985f
C1625 VTAIL.n482 VSUBS 0.013432f
C1626 VTAIL.n483 VSUBS 0.012686f
C1627 VTAIL.n484 VSUBS 0.023608f
C1628 VTAIL.n485 VSUBS 0.023608f
C1629 VTAIL.n486 VSUBS 0.012686f
C1630 VTAIL.n487 VSUBS 0.013432f
C1631 VTAIL.n488 VSUBS 0.029985f
C1632 VTAIL.n489 VSUBS 0.029985f
C1633 VTAIL.n490 VSUBS 0.013432f
C1634 VTAIL.n491 VSUBS 0.012686f
C1635 VTAIL.n492 VSUBS 0.023608f
C1636 VTAIL.n493 VSUBS 0.023608f
C1637 VTAIL.n494 VSUBS 0.012686f
C1638 VTAIL.n495 VSUBS 0.013432f
C1639 VTAIL.n496 VSUBS 0.029985f
C1640 VTAIL.n497 VSUBS 0.029985f
C1641 VTAIL.n498 VSUBS 0.013432f
C1642 VTAIL.n499 VSUBS 0.012686f
C1643 VTAIL.n500 VSUBS 0.023608f
C1644 VTAIL.n501 VSUBS 0.023608f
C1645 VTAIL.n502 VSUBS 0.012686f
C1646 VTAIL.n503 VSUBS 0.013432f
C1647 VTAIL.n504 VSUBS 0.029985f
C1648 VTAIL.n505 VSUBS 0.029985f
C1649 VTAIL.n506 VSUBS 0.013432f
C1650 VTAIL.n507 VSUBS 0.012686f
C1651 VTAIL.n508 VSUBS 0.023608f
C1652 VTAIL.n509 VSUBS 0.023608f
C1653 VTAIL.n510 VSUBS 0.012686f
C1654 VTAIL.n511 VSUBS 0.013059f
C1655 VTAIL.n512 VSUBS 0.013059f
C1656 VTAIL.n513 VSUBS 0.029985f
C1657 VTAIL.n514 VSUBS 0.029985f
C1658 VTAIL.n515 VSUBS 0.013432f
C1659 VTAIL.n516 VSUBS 0.012686f
C1660 VTAIL.n517 VSUBS 0.023608f
C1661 VTAIL.n518 VSUBS 0.023608f
C1662 VTAIL.n519 VSUBS 0.012686f
C1663 VTAIL.n520 VSUBS 0.013432f
C1664 VTAIL.n521 VSUBS 0.029985f
C1665 VTAIL.n522 VSUBS 0.029985f
C1666 VTAIL.n523 VSUBS 0.013432f
C1667 VTAIL.n524 VSUBS 0.012686f
C1668 VTAIL.n525 VSUBS 0.023608f
C1669 VTAIL.n526 VSUBS 0.023608f
C1670 VTAIL.n527 VSUBS 0.012686f
C1671 VTAIL.n528 VSUBS 0.013432f
C1672 VTAIL.n529 VSUBS 0.029985f
C1673 VTAIL.n530 VSUBS 0.076005f
C1674 VTAIL.n531 VSUBS 0.013432f
C1675 VTAIL.n532 VSUBS 0.012686f
C1676 VTAIL.n533 VSUBS 0.056827f
C1677 VTAIL.n534 VSUBS 0.038442f
C1678 VTAIL.n535 VSUBS 0.268342f
C1679 VTAIL.n536 VSUBS 0.026943f
C1680 VTAIL.n537 VSUBS 0.023608f
C1681 VTAIL.n538 VSUBS 0.012686f
C1682 VTAIL.n539 VSUBS 0.029985f
C1683 VTAIL.n540 VSUBS 0.013432f
C1684 VTAIL.n541 VSUBS 0.023608f
C1685 VTAIL.n542 VSUBS 0.012686f
C1686 VTAIL.n543 VSUBS 0.029985f
C1687 VTAIL.n544 VSUBS 0.013432f
C1688 VTAIL.n545 VSUBS 0.023608f
C1689 VTAIL.n546 VSUBS 0.012686f
C1690 VTAIL.n547 VSUBS 0.029985f
C1691 VTAIL.n548 VSUBS 0.013432f
C1692 VTAIL.n549 VSUBS 0.023608f
C1693 VTAIL.n550 VSUBS 0.012686f
C1694 VTAIL.n551 VSUBS 0.029985f
C1695 VTAIL.n552 VSUBS 0.029985f
C1696 VTAIL.n553 VSUBS 0.013432f
C1697 VTAIL.n554 VSUBS 0.023608f
C1698 VTAIL.n555 VSUBS 0.012686f
C1699 VTAIL.n556 VSUBS 0.029985f
C1700 VTAIL.n557 VSUBS 0.013432f
C1701 VTAIL.n558 VSUBS 0.023608f
C1702 VTAIL.n559 VSUBS 0.012686f
C1703 VTAIL.n560 VSUBS 0.029985f
C1704 VTAIL.n561 VSUBS 0.013432f
C1705 VTAIL.n562 VSUBS 0.023608f
C1706 VTAIL.n563 VSUBS 0.012686f
C1707 VTAIL.n564 VSUBS 0.029985f
C1708 VTAIL.n565 VSUBS 0.013432f
C1709 VTAIL.n566 VSUBS 0.023608f
C1710 VTAIL.n567 VSUBS 0.012686f
C1711 VTAIL.n568 VSUBS 0.029985f
C1712 VTAIL.n569 VSUBS 0.013432f
C1713 VTAIL.n570 VSUBS 0.194481f
C1714 VTAIL.t13 VSUBS 0.064429f
C1715 VTAIL.n571 VSUBS 0.022489f
C1716 VTAIL.n572 VSUBS 0.019075f
C1717 VTAIL.n573 VSUBS 0.012686f
C1718 VTAIL.n574 VSUBS 1.93935f
C1719 VTAIL.n575 VSUBS 0.023608f
C1720 VTAIL.n576 VSUBS 0.012686f
C1721 VTAIL.n577 VSUBS 0.013432f
C1722 VTAIL.n578 VSUBS 0.029985f
C1723 VTAIL.n579 VSUBS 0.029985f
C1724 VTAIL.n580 VSUBS 0.013432f
C1725 VTAIL.n581 VSUBS 0.012686f
C1726 VTAIL.n582 VSUBS 0.023608f
C1727 VTAIL.n583 VSUBS 0.023608f
C1728 VTAIL.n584 VSUBS 0.012686f
C1729 VTAIL.n585 VSUBS 0.013432f
C1730 VTAIL.n586 VSUBS 0.029985f
C1731 VTAIL.n587 VSUBS 0.029985f
C1732 VTAIL.n588 VSUBS 0.013432f
C1733 VTAIL.n589 VSUBS 0.012686f
C1734 VTAIL.n590 VSUBS 0.023608f
C1735 VTAIL.n591 VSUBS 0.023608f
C1736 VTAIL.n592 VSUBS 0.012686f
C1737 VTAIL.n593 VSUBS 0.013432f
C1738 VTAIL.n594 VSUBS 0.029985f
C1739 VTAIL.n595 VSUBS 0.029985f
C1740 VTAIL.n596 VSUBS 0.013432f
C1741 VTAIL.n597 VSUBS 0.012686f
C1742 VTAIL.n598 VSUBS 0.023608f
C1743 VTAIL.n599 VSUBS 0.023608f
C1744 VTAIL.n600 VSUBS 0.012686f
C1745 VTAIL.n601 VSUBS 0.013432f
C1746 VTAIL.n602 VSUBS 0.029985f
C1747 VTAIL.n603 VSUBS 0.029985f
C1748 VTAIL.n604 VSUBS 0.013432f
C1749 VTAIL.n605 VSUBS 0.012686f
C1750 VTAIL.n606 VSUBS 0.023608f
C1751 VTAIL.n607 VSUBS 0.023608f
C1752 VTAIL.n608 VSUBS 0.012686f
C1753 VTAIL.n609 VSUBS 0.013432f
C1754 VTAIL.n610 VSUBS 0.029985f
C1755 VTAIL.n611 VSUBS 0.029985f
C1756 VTAIL.n612 VSUBS 0.013432f
C1757 VTAIL.n613 VSUBS 0.012686f
C1758 VTAIL.n614 VSUBS 0.023608f
C1759 VTAIL.n615 VSUBS 0.023608f
C1760 VTAIL.n616 VSUBS 0.012686f
C1761 VTAIL.n617 VSUBS 0.013059f
C1762 VTAIL.n618 VSUBS 0.013059f
C1763 VTAIL.n619 VSUBS 0.029985f
C1764 VTAIL.n620 VSUBS 0.029985f
C1765 VTAIL.n621 VSUBS 0.013432f
C1766 VTAIL.n622 VSUBS 0.012686f
C1767 VTAIL.n623 VSUBS 0.023608f
C1768 VTAIL.n624 VSUBS 0.023608f
C1769 VTAIL.n625 VSUBS 0.012686f
C1770 VTAIL.n626 VSUBS 0.013432f
C1771 VTAIL.n627 VSUBS 0.029985f
C1772 VTAIL.n628 VSUBS 0.029985f
C1773 VTAIL.n629 VSUBS 0.013432f
C1774 VTAIL.n630 VSUBS 0.012686f
C1775 VTAIL.n631 VSUBS 0.023608f
C1776 VTAIL.n632 VSUBS 0.023608f
C1777 VTAIL.n633 VSUBS 0.012686f
C1778 VTAIL.n634 VSUBS 0.013432f
C1779 VTAIL.n635 VSUBS 0.029985f
C1780 VTAIL.n636 VSUBS 0.076005f
C1781 VTAIL.n637 VSUBS 0.013432f
C1782 VTAIL.n638 VSUBS 0.012686f
C1783 VTAIL.n639 VSUBS 0.056827f
C1784 VTAIL.n640 VSUBS 0.038442f
C1785 VTAIL.n641 VSUBS 0.268342f
C1786 VTAIL.t10 VSUBS 0.355023f
C1787 VTAIL.t9 VSUBS 0.355023f
C1788 VTAIL.n642 VSUBS 2.82936f
C1789 VTAIL.n643 VSUBS 0.999054f
C1790 VTAIL.n644 VSUBS 0.026943f
C1791 VTAIL.n645 VSUBS 0.023608f
C1792 VTAIL.n646 VSUBS 0.012686f
C1793 VTAIL.n647 VSUBS 0.029985f
C1794 VTAIL.n648 VSUBS 0.013432f
C1795 VTAIL.n649 VSUBS 0.023608f
C1796 VTAIL.n650 VSUBS 0.012686f
C1797 VTAIL.n651 VSUBS 0.029985f
C1798 VTAIL.n652 VSUBS 0.013432f
C1799 VTAIL.n653 VSUBS 0.023608f
C1800 VTAIL.n654 VSUBS 0.012686f
C1801 VTAIL.n655 VSUBS 0.029985f
C1802 VTAIL.n656 VSUBS 0.013432f
C1803 VTAIL.n657 VSUBS 0.023608f
C1804 VTAIL.n658 VSUBS 0.012686f
C1805 VTAIL.n659 VSUBS 0.029985f
C1806 VTAIL.n660 VSUBS 0.029985f
C1807 VTAIL.n661 VSUBS 0.013432f
C1808 VTAIL.n662 VSUBS 0.023608f
C1809 VTAIL.n663 VSUBS 0.012686f
C1810 VTAIL.n664 VSUBS 0.029985f
C1811 VTAIL.n665 VSUBS 0.013432f
C1812 VTAIL.n666 VSUBS 0.023608f
C1813 VTAIL.n667 VSUBS 0.012686f
C1814 VTAIL.n668 VSUBS 0.029985f
C1815 VTAIL.n669 VSUBS 0.013432f
C1816 VTAIL.n670 VSUBS 0.023608f
C1817 VTAIL.n671 VSUBS 0.012686f
C1818 VTAIL.n672 VSUBS 0.029985f
C1819 VTAIL.n673 VSUBS 0.013432f
C1820 VTAIL.n674 VSUBS 0.023608f
C1821 VTAIL.n675 VSUBS 0.012686f
C1822 VTAIL.n676 VSUBS 0.029985f
C1823 VTAIL.n677 VSUBS 0.013432f
C1824 VTAIL.n678 VSUBS 0.194481f
C1825 VTAIL.t14 VSUBS 0.064429f
C1826 VTAIL.n679 VSUBS 0.022489f
C1827 VTAIL.n680 VSUBS 0.019075f
C1828 VTAIL.n681 VSUBS 0.012686f
C1829 VTAIL.n682 VSUBS 1.93935f
C1830 VTAIL.n683 VSUBS 0.023608f
C1831 VTAIL.n684 VSUBS 0.012686f
C1832 VTAIL.n685 VSUBS 0.013432f
C1833 VTAIL.n686 VSUBS 0.029985f
C1834 VTAIL.n687 VSUBS 0.029985f
C1835 VTAIL.n688 VSUBS 0.013432f
C1836 VTAIL.n689 VSUBS 0.012686f
C1837 VTAIL.n690 VSUBS 0.023608f
C1838 VTAIL.n691 VSUBS 0.023608f
C1839 VTAIL.n692 VSUBS 0.012686f
C1840 VTAIL.n693 VSUBS 0.013432f
C1841 VTAIL.n694 VSUBS 0.029985f
C1842 VTAIL.n695 VSUBS 0.029985f
C1843 VTAIL.n696 VSUBS 0.013432f
C1844 VTAIL.n697 VSUBS 0.012686f
C1845 VTAIL.n698 VSUBS 0.023608f
C1846 VTAIL.n699 VSUBS 0.023608f
C1847 VTAIL.n700 VSUBS 0.012686f
C1848 VTAIL.n701 VSUBS 0.013432f
C1849 VTAIL.n702 VSUBS 0.029985f
C1850 VTAIL.n703 VSUBS 0.029985f
C1851 VTAIL.n704 VSUBS 0.013432f
C1852 VTAIL.n705 VSUBS 0.012686f
C1853 VTAIL.n706 VSUBS 0.023608f
C1854 VTAIL.n707 VSUBS 0.023608f
C1855 VTAIL.n708 VSUBS 0.012686f
C1856 VTAIL.n709 VSUBS 0.013432f
C1857 VTAIL.n710 VSUBS 0.029985f
C1858 VTAIL.n711 VSUBS 0.029985f
C1859 VTAIL.n712 VSUBS 0.013432f
C1860 VTAIL.n713 VSUBS 0.012686f
C1861 VTAIL.n714 VSUBS 0.023608f
C1862 VTAIL.n715 VSUBS 0.023608f
C1863 VTAIL.n716 VSUBS 0.012686f
C1864 VTAIL.n717 VSUBS 0.013432f
C1865 VTAIL.n718 VSUBS 0.029985f
C1866 VTAIL.n719 VSUBS 0.029985f
C1867 VTAIL.n720 VSUBS 0.013432f
C1868 VTAIL.n721 VSUBS 0.012686f
C1869 VTAIL.n722 VSUBS 0.023608f
C1870 VTAIL.n723 VSUBS 0.023608f
C1871 VTAIL.n724 VSUBS 0.012686f
C1872 VTAIL.n725 VSUBS 0.013059f
C1873 VTAIL.n726 VSUBS 0.013059f
C1874 VTAIL.n727 VSUBS 0.029985f
C1875 VTAIL.n728 VSUBS 0.029985f
C1876 VTAIL.n729 VSUBS 0.013432f
C1877 VTAIL.n730 VSUBS 0.012686f
C1878 VTAIL.n731 VSUBS 0.023608f
C1879 VTAIL.n732 VSUBS 0.023608f
C1880 VTAIL.n733 VSUBS 0.012686f
C1881 VTAIL.n734 VSUBS 0.013432f
C1882 VTAIL.n735 VSUBS 0.029985f
C1883 VTAIL.n736 VSUBS 0.029985f
C1884 VTAIL.n737 VSUBS 0.013432f
C1885 VTAIL.n738 VSUBS 0.012686f
C1886 VTAIL.n739 VSUBS 0.023608f
C1887 VTAIL.n740 VSUBS 0.023608f
C1888 VTAIL.n741 VSUBS 0.012686f
C1889 VTAIL.n742 VSUBS 0.013432f
C1890 VTAIL.n743 VSUBS 0.029985f
C1891 VTAIL.n744 VSUBS 0.076005f
C1892 VTAIL.n745 VSUBS 0.013432f
C1893 VTAIL.n746 VSUBS 0.012686f
C1894 VTAIL.n747 VSUBS 0.056827f
C1895 VTAIL.n748 VSUBS 0.038442f
C1896 VTAIL.n749 VSUBS 2.01242f
C1897 VTAIL.n750 VSUBS 0.026943f
C1898 VTAIL.n751 VSUBS 0.023608f
C1899 VTAIL.n752 VSUBS 0.012686f
C1900 VTAIL.n753 VSUBS 0.029985f
C1901 VTAIL.n754 VSUBS 0.013432f
C1902 VTAIL.n755 VSUBS 0.023608f
C1903 VTAIL.n756 VSUBS 0.012686f
C1904 VTAIL.n757 VSUBS 0.029985f
C1905 VTAIL.n758 VSUBS 0.013432f
C1906 VTAIL.n759 VSUBS 0.023608f
C1907 VTAIL.n760 VSUBS 0.012686f
C1908 VTAIL.n761 VSUBS 0.029985f
C1909 VTAIL.n762 VSUBS 0.013432f
C1910 VTAIL.n763 VSUBS 0.023608f
C1911 VTAIL.n764 VSUBS 0.012686f
C1912 VTAIL.n765 VSUBS 0.029985f
C1913 VTAIL.n766 VSUBS 0.013432f
C1914 VTAIL.n767 VSUBS 0.023608f
C1915 VTAIL.n768 VSUBS 0.012686f
C1916 VTAIL.n769 VSUBS 0.029985f
C1917 VTAIL.n770 VSUBS 0.013432f
C1918 VTAIL.n771 VSUBS 0.023608f
C1919 VTAIL.n772 VSUBS 0.012686f
C1920 VTAIL.n773 VSUBS 0.029985f
C1921 VTAIL.n774 VSUBS 0.013432f
C1922 VTAIL.n775 VSUBS 0.023608f
C1923 VTAIL.n776 VSUBS 0.012686f
C1924 VTAIL.n777 VSUBS 0.029985f
C1925 VTAIL.n778 VSUBS 0.013432f
C1926 VTAIL.n779 VSUBS 0.023608f
C1927 VTAIL.n780 VSUBS 0.012686f
C1928 VTAIL.n781 VSUBS 0.029985f
C1929 VTAIL.n782 VSUBS 0.013432f
C1930 VTAIL.n783 VSUBS 0.194481f
C1931 VTAIL.t0 VSUBS 0.064429f
C1932 VTAIL.n784 VSUBS 0.022489f
C1933 VTAIL.n785 VSUBS 0.019075f
C1934 VTAIL.n786 VSUBS 0.012686f
C1935 VTAIL.n787 VSUBS 1.93935f
C1936 VTAIL.n788 VSUBS 0.023608f
C1937 VTAIL.n789 VSUBS 0.012686f
C1938 VTAIL.n790 VSUBS 0.013432f
C1939 VTAIL.n791 VSUBS 0.029985f
C1940 VTAIL.n792 VSUBS 0.029985f
C1941 VTAIL.n793 VSUBS 0.013432f
C1942 VTAIL.n794 VSUBS 0.012686f
C1943 VTAIL.n795 VSUBS 0.023608f
C1944 VTAIL.n796 VSUBS 0.023608f
C1945 VTAIL.n797 VSUBS 0.012686f
C1946 VTAIL.n798 VSUBS 0.013432f
C1947 VTAIL.n799 VSUBS 0.029985f
C1948 VTAIL.n800 VSUBS 0.029985f
C1949 VTAIL.n801 VSUBS 0.013432f
C1950 VTAIL.n802 VSUBS 0.012686f
C1951 VTAIL.n803 VSUBS 0.023608f
C1952 VTAIL.n804 VSUBS 0.023608f
C1953 VTAIL.n805 VSUBS 0.012686f
C1954 VTAIL.n806 VSUBS 0.013432f
C1955 VTAIL.n807 VSUBS 0.029985f
C1956 VTAIL.n808 VSUBS 0.029985f
C1957 VTAIL.n809 VSUBS 0.013432f
C1958 VTAIL.n810 VSUBS 0.012686f
C1959 VTAIL.n811 VSUBS 0.023608f
C1960 VTAIL.n812 VSUBS 0.023608f
C1961 VTAIL.n813 VSUBS 0.012686f
C1962 VTAIL.n814 VSUBS 0.013432f
C1963 VTAIL.n815 VSUBS 0.029985f
C1964 VTAIL.n816 VSUBS 0.029985f
C1965 VTAIL.n817 VSUBS 0.013432f
C1966 VTAIL.n818 VSUBS 0.012686f
C1967 VTAIL.n819 VSUBS 0.023608f
C1968 VTAIL.n820 VSUBS 0.023608f
C1969 VTAIL.n821 VSUBS 0.012686f
C1970 VTAIL.n822 VSUBS 0.013432f
C1971 VTAIL.n823 VSUBS 0.029985f
C1972 VTAIL.n824 VSUBS 0.029985f
C1973 VTAIL.n825 VSUBS 0.029985f
C1974 VTAIL.n826 VSUBS 0.013432f
C1975 VTAIL.n827 VSUBS 0.012686f
C1976 VTAIL.n828 VSUBS 0.023608f
C1977 VTAIL.n829 VSUBS 0.023608f
C1978 VTAIL.n830 VSUBS 0.012686f
C1979 VTAIL.n831 VSUBS 0.013059f
C1980 VTAIL.n832 VSUBS 0.013059f
C1981 VTAIL.n833 VSUBS 0.029985f
C1982 VTAIL.n834 VSUBS 0.029985f
C1983 VTAIL.n835 VSUBS 0.013432f
C1984 VTAIL.n836 VSUBS 0.012686f
C1985 VTAIL.n837 VSUBS 0.023608f
C1986 VTAIL.n838 VSUBS 0.023608f
C1987 VTAIL.n839 VSUBS 0.012686f
C1988 VTAIL.n840 VSUBS 0.013432f
C1989 VTAIL.n841 VSUBS 0.029985f
C1990 VTAIL.n842 VSUBS 0.029985f
C1991 VTAIL.n843 VSUBS 0.013432f
C1992 VTAIL.n844 VSUBS 0.012686f
C1993 VTAIL.n845 VSUBS 0.023608f
C1994 VTAIL.n846 VSUBS 0.023608f
C1995 VTAIL.n847 VSUBS 0.012686f
C1996 VTAIL.n848 VSUBS 0.013432f
C1997 VTAIL.n849 VSUBS 0.029985f
C1998 VTAIL.n850 VSUBS 0.076005f
C1999 VTAIL.n851 VSUBS 0.013432f
C2000 VTAIL.n852 VSUBS 0.012686f
C2001 VTAIL.n853 VSUBS 0.056827f
C2002 VTAIL.n854 VSUBS 0.038442f
C2003 VTAIL.n855 VSUBS 2.00799f
C2004 VP.n0 VSUBS 0.034229f
C2005 VP.t5 VSUBS 3.93138f
C2006 VP.n1 VSUBS 0.05222f
C2007 VP.n2 VSUBS 0.025962f
C2008 VP.n3 VSUBS 0.031187f
C2009 VP.n4 VSUBS 0.025962f
C2010 VP.n5 VSUBS 0.0379f
C2011 VP.n6 VSUBS 0.025962f
C2012 VP.t0 VSUBS 3.93138f
C2013 VP.n7 VSUBS 0.048387f
C2014 VP.n8 VSUBS 0.025962f
C2015 VP.n9 VSUBS 0.048387f
C2016 VP.n10 VSUBS 0.034229f
C2017 VP.t2 VSUBS 3.93138f
C2018 VP.n11 VSUBS 0.05222f
C2019 VP.n12 VSUBS 0.025962f
C2020 VP.n13 VSUBS 0.031187f
C2021 VP.n14 VSUBS 0.025962f
C2022 VP.n15 VSUBS 0.0379f
C2023 VP.n16 VSUBS 0.275083f
C2024 VP.t4 VSUBS 3.93138f
C2025 VP.t6 VSUBS 4.19906f
C2026 VP.n17 VSUBS 1.39685f
C2027 VP.n18 VSUBS 1.44394f
C2028 VP.n19 VSUBS 0.041698f
C2029 VP.n20 VSUBS 0.048387f
C2030 VP.n21 VSUBS 0.025962f
C2031 VP.n22 VSUBS 0.025962f
C2032 VP.n23 VSUBS 0.025962f
C2033 VP.n24 VSUBS 0.0379f
C2034 VP.n25 VSUBS 0.048387f
C2035 VP.t3 VSUBS 3.93138f
C2036 VP.n26 VSUBS 1.35771f
C2037 VP.n27 VSUBS 0.041698f
C2038 VP.n28 VSUBS 0.025962f
C2039 VP.n29 VSUBS 0.025962f
C2040 VP.n30 VSUBS 0.025962f
C2041 VP.n31 VSUBS 0.048387f
C2042 VP.n32 VSUBS 0.050678f
C2043 VP.n33 VSUBS 0.02129f
C2044 VP.n34 VSUBS 0.025962f
C2045 VP.n35 VSUBS 0.025962f
C2046 VP.n36 VSUBS 0.025962f
C2047 VP.n37 VSUBS 0.048387f
C2048 VP.n38 VSUBS 0.02832f
C2049 VP.n39 VSUBS 1.44606f
C2050 VP.n40 VSUBS 1.7728f
C2051 VP.n41 VSUBS 1.78901f
C2052 VP.t1 VSUBS 3.93138f
C2053 VP.n42 VSUBS 1.44606f
C2054 VP.n43 VSUBS 0.02832f
C2055 VP.n44 VSUBS 0.034229f
C2056 VP.n45 VSUBS 0.025962f
C2057 VP.n46 VSUBS 0.025962f
C2058 VP.n47 VSUBS 0.05222f
C2059 VP.n48 VSUBS 0.02129f
C2060 VP.n49 VSUBS 0.050678f
C2061 VP.n50 VSUBS 0.025962f
C2062 VP.n51 VSUBS 0.025962f
C2063 VP.n52 VSUBS 0.025962f
C2064 VP.n53 VSUBS 0.031187f
C2065 VP.n54 VSUBS 1.35771f
C2066 VP.n55 VSUBS 0.041698f
C2067 VP.n56 VSUBS 0.048387f
C2068 VP.n57 VSUBS 0.025962f
C2069 VP.n58 VSUBS 0.025962f
C2070 VP.n59 VSUBS 0.025962f
C2071 VP.n60 VSUBS 0.0379f
C2072 VP.n61 VSUBS 0.048387f
C2073 VP.t7 VSUBS 3.93138f
C2074 VP.n62 VSUBS 1.35771f
C2075 VP.n63 VSUBS 0.041698f
C2076 VP.n64 VSUBS 0.025962f
C2077 VP.n65 VSUBS 0.025962f
C2078 VP.n66 VSUBS 0.025962f
C2079 VP.n67 VSUBS 0.048387f
C2080 VP.n68 VSUBS 0.050678f
C2081 VP.n69 VSUBS 0.02129f
C2082 VP.n70 VSUBS 0.025962f
C2083 VP.n71 VSUBS 0.025962f
C2084 VP.n72 VSUBS 0.025962f
C2085 VP.n73 VSUBS 0.048387f
C2086 VP.n74 VSUBS 0.02832f
C2087 VP.n75 VSUBS 1.44606f
C2088 VP.n76 VSUBS 0.048754f
.ends

