* NGSPICE file created from diff_pair_sample_1529.ext - technology: sky130A

.subckt diff_pair_sample_1529 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t9 VN.t0 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=2.4717 pd=15.31 as=2.4717 ps=15.31 w=14.98 l=1.37
X1 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=5.8422 pd=30.74 as=0 ps=0 w=14.98 l=1.37
X2 VDD2.t1 VN.t1 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=5.8422 pd=30.74 as=2.4717 ps=15.31 w=14.98 l=1.37
X3 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=5.8422 pd=30.74 as=0 ps=0 w=14.98 l=1.37
X4 VDD1.t5 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=5.8422 pd=30.74 as=2.4717 ps=15.31 w=14.98 l=1.37
X5 VDD1.t4 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.4717 pd=15.31 as=5.8422 ps=30.74 w=14.98 l=1.37
X6 VTAIL.t11 VP.t2 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=2.4717 pd=15.31 as=2.4717 ps=15.31 w=14.98 l=1.37
X7 VDD2.t3 VN.t2 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=5.8422 pd=30.74 as=2.4717 ps=15.31 w=14.98 l=1.37
X8 VTAIL.t10 VP.t3 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.4717 pd=15.31 as=2.4717 ps=15.31 w=14.98 l=1.37
X9 VDD1.t1 VP.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.8422 pd=30.74 as=2.4717 ps=15.31 w=14.98 l=1.37
X10 VDD2.t5 VN.t3 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=2.4717 pd=15.31 as=5.8422 ps=30.74 w=14.98 l=1.37
X11 VTAIL.t5 VN.t4 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=2.4717 pd=15.31 as=2.4717 ps=15.31 w=14.98 l=1.37
X12 VDD1.t0 VP.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.4717 pd=15.31 as=5.8422 ps=30.74 w=14.98 l=1.37
X13 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.8422 pd=30.74 as=0 ps=0 w=14.98 l=1.37
X14 VDD2.t2 VN.t5 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=2.4717 pd=15.31 as=5.8422 ps=30.74 w=14.98 l=1.37
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.8422 pd=30.74 as=0 ps=0 w=14.98 l=1.37
R0 VN.n3 VN.t2 297.433
R1 VN.n13 VN.t3 297.433
R2 VN.n2 VN.t0 263.517
R3 VN.n8 VN.t5 263.517
R4 VN.n12 VN.t4 263.517
R5 VN.n18 VN.t1 263.517
R6 VN.n9 VN.n8 176.055
R7 VN.n19 VN.n18 176.055
R8 VN.n17 VN.n10 161.3
R9 VN.n16 VN.n15 161.3
R10 VN.n14 VN.n11 161.3
R11 VN.n7 VN.n0 161.3
R12 VN.n6 VN.n5 161.3
R13 VN.n4 VN.n1 161.3
R14 VN.n6 VN.n1 55.1086
R15 VN.n16 VN.n11 55.1086
R16 VN VN.n19 46.3812
R17 VN.n3 VN.n2 41.862
R18 VN.n13 VN.n12 41.862
R19 VN.n7 VN.n6 26.0455
R20 VN.n17 VN.n16 26.0455
R21 VN.n2 VN.n1 24.5923
R22 VN.n12 VN.n11 24.5923
R23 VN.n14 VN.n13 17.7677
R24 VN.n4 VN.n3 17.7677
R25 VN.n8 VN.n7 9.83723
R26 VN.n18 VN.n17 9.83723
R27 VN.n19 VN.n10 0.189894
R28 VN.n15 VN.n10 0.189894
R29 VN.n15 VN.n14 0.189894
R30 VN.n5 VN.n4 0.189894
R31 VN.n5 VN.n0 0.189894
R32 VN.n9 VN.n0 0.189894
R33 VN VN.n9 0.0516364
R34 VDD2.n1 VDD2.t3 62.8572
R35 VDD2.n2 VDD2.t1 61.8137
R36 VDD2.n1 VDD2.n0 60.8027
R37 VDD2 VDD2.n3 60.7999
R38 VDD2.n2 VDD2.n1 41.392
R39 VDD2.n3 VDD2.t0 1.32226
R40 VDD2.n3 VDD2.t5 1.32226
R41 VDD2.n0 VDD2.t4 1.32226
R42 VDD2.n0 VDD2.t2 1.32226
R43 VDD2 VDD2.n2 1.15783
R44 VTAIL.n7 VTAIL.t6 45.1349
R45 VTAIL.n11 VTAIL.t4 45.1347
R46 VTAIL.n2 VTAIL.t0 45.1347
R47 VTAIL.n10 VTAIL.t2 45.1347
R48 VTAIL.n9 VTAIL.n8 43.8131
R49 VTAIL.n6 VTAIL.n5 43.8131
R50 VTAIL.n1 VTAIL.n0 43.8129
R51 VTAIL.n4 VTAIL.n3 43.8129
R52 VTAIL.n6 VTAIL.n4 28.2117
R53 VTAIL.n11 VTAIL.n10 26.7462
R54 VTAIL.n7 VTAIL.n6 1.46602
R55 VTAIL.n10 VTAIL.n9 1.46602
R56 VTAIL.n4 VTAIL.n2 1.46602
R57 VTAIL.n0 VTAIL.t7 1.32226
R58 VTAIL.n0 VTAIL.t9 1.32226
R59 VTAIL.n3 VTAIL.t1 1.32226
R60 VTAIL.n3 VTAIL.t10 1.32226
R61 VTAIL.n8 VTAIL.t3 1.32226
R62 VTAIL.n8 VTAIL.t11 1.32226
R63 VTAIL.n5 VTAIL.t8 1.32226
R64 VTAIL.n5 VTAIL.t5 1.32226
R65 VTAIL.n9 VTAIL.n7 1.20309
R66 VTAIL.n2 VTAIL.n1 1.20309
R67 VTAIL VTAIL.n11 1.04145
R68 VTAIL VTAIL.n1 0.425069
R69 B.n786 B.n785 585
R70 B.n330 B.n109 585
R71 B.n329 B.n328 585
R72 B.n327 B.n326 585
R73 B.n325 B.n324 585
R74 B.n323 B.n322 585
R75 B.n321 B.n320 585
R76 B.n319 B.n318 585
R77 B.n317 B.n316 585
R78 B.n315 B.n314 585
R79 B.n313 B.n312 585
R80 B.n311 B.n310 585
R81 B.n309 B.n308 585
R82 B.n307 B.n306 585
R83 B.n305 B.n304 585
R84 B.n303 B.n302 585
R85 B.n301 B.n300 585
R86 B.n299 B.n298 585
R87 B.n297 B.n296 585
R88 B.n295 B.n294 585
R89 B.n293 B.n292 585
R90 B.n291 B.n290 585
R91 B.n289 B.n288 585
R92 B.n287 B.n286 585
R93 B.n285 B.n284 585
R94 B.n283 B.n282 585
R95 B.n281 B.n280 585
R96 B.n279 B.n278 585
R97 B.n277 B.n276 585
R98 B.n275 B.n274 585
R99 B.n273 B.n272 585
R100 B.n271 B.n270 585
R101 B.n269 B.n268 585
R102 B.n267 B.n266 585
R103 B.n265 B.n264 585
R104 B.n263 B.n262 585
R105 B.n261 B.n260 585
R106 B.n259 B.n258 585
R107 B.n257 B.n256 585
R108 B.n255 B.n254 585
R109 B.n253 B.n252 585
R110 B.n251 B.n250 585
R111 B.n249 B.n248 585
R112 B.n247 B.n246 585
R113 B.n245 B.n244 585
R114 B.n243 B.n242 585
R115 B.n241 B.n240 585
R116 B.n239 B.n238 585
R117 B.n237 B.n236 585
R118 B.n235 B.n234 585
R119 B.n233 B.n232 585
R120 B.n231 B.n230 585
R121 B.n229 B.n228 585
R122 B.n227 B.n226 585
R123 B.n225 B.n224 585
R124 B.n223 B.n222 585
R125 B.n221 B.n220 585
R126 B.n219 B.n218 585
R127 B.n217 B.n216 585
R128 B.n215 B.n214 585
R129 B.n213 B.n212 585
R130 B.n211 B.n210 585
R131 B.n209 B.n208 585
R132 B.n207 B.n206 585
R133 B.n205 B.n204 585
R134 B.n203 B.n202 585
R135 B.n201 B.n200 585
R136 B.n199 B.n198 585
R137 B.n197 B.n196 585
R138 B.n195 B.n194 585
R139 B.n193 B.n192 585
R140 B.n191 B.n190 585
R141 B.n189 B.n188 585
R142 B.n187 B.n186 585
R143 B.n185 B.n184 585
R144 B.n183 B.n182 585
R145 B.n181 B.n180 585
R146 B.n179 B.n178 585
R147 B.n177 B.n176 585
R148 B.n175 B.n174 585
R149 B.n173 B.n172 585
R150 B.n171 B.n170 585
R151 B.n169 B.n168 585
R152 B.n167 B.n166 585
R153 B.n165 B.n164 585
R154 B.n163 B.n162 585
R155 B.n161 B.n160 585
R156 B.n159 B.n158 585
R157 B.n157 B.n156 585
R158 B.n155 B.n154 585
R159 B.n153 B.n152 585
R160 B.n151 B.n150 585
R161 B.n149 B.n148 585
R162 B.n147 B.n146 585
R163 B.n145 B.n144 585
R164 B.n143 B.n142 585
R165 B.n141 B.n140 585
R166 B.n139 B.n138 585
R167 B.n137 B.n136 585
R168 B.n135 B.n134 585
R169 B.n133 B.n132 585
R170 B.n131 B.n130 585
R171 B.n129 B.n128 585
R172 B.n127 B.n126 585
R173 B.n125 B.n124 585
R174 B.n123 B.n122 585
R175 B.n121 B.n120 585
R176 B.n119 B.n118 585
R177 B.n117 B.n116 585
R178 B.n53 B.n52 585
R179 B.n784 B.n54 585
R180 B.n789 B.n54 585
R181 B.n783 B.n782 585
R182 B.n782 B.n50 585
R183 B.n781 B.n49 585
R184 B.n795 B.n49 585
R185 B.n780 B.n48 585
R186 B.n796 B.n48 585
R187 B.n779 B.n47 585
R188 B.n797 B.n47 585
R189 B.n778 B.n777 585
R190 B.n777 B.n46 585
R191 B.n776 B.n42 585
R192 B.n803 B.n42 585
R193 B.n775 B.n41 585
R194 B.n804 B.n41 585
R195 B.n774 B.n40 585
R196 B.n805 B.n40 585
R197 B.n773 B.n772 585
R198 B.n772 B.n36 585
R199 B.n771 B.n35 585
R200 B.n811 B.n35 585
R201 B.n770 B.n34 585
R202 B.n812 B.n34 585
R203 B.n769 B.n33 585
R204 B.n813 B.n33 585
R205 B.n768 B.n767 585
R206 B.n767 B.n32 585
R207 B.n766 B.n28 585
R208 B.n819 B.n28 585
R209 B.n765 B.n27 585
R210 B.n820 B.n27 585
R211 B.n764 B.n26 585
R212 B.n821 B.n26 585
R213 B.n763 B.n762 585
R214 B.n762 B.n22 585
R215 B.n761 B.n21 585
R216 B.n827 B.n21 585
R217 B.n760 B.n20 585
R218 B.n828 B.n20 585
R219 B.n759 B.n19 585
R220 B.n829 B.n19 585
R221 B.n758 B.n757 585
R222 B.n757 B.n15 585
R223 B.n756 B.n14 585
R224 B.n835 B.n14 585
R225 B.n755 B.n13 585
R226 B.n836 B.n13 585
R227 B.n754 B.n12 585
R228 B.n837 B.n12 585
R229 B.n753 B.n752 585
R230 B.n752 B.n8 585
R231 B.n751 B.n7 585
R232 B.n843 B.n7 585
R233 B.n750 B.n6 585
R234 B.n844 B.n6 585
R235 B.n749 B.n5 585
R236 B.n845 B.n5 585
R237 B.n748 B.n747 585
R238 B.n747 B.n4 585
R239 B.n746 B.n331 585
R240 B.n746 B.n745 585
R241 B.n736 B.n332 585
R242 B.n333 B.n332 585
R243 B.n738 B.n737 585
R244 B.n739 B.n738 585
R245 B.n735 B.n337 585
R246 B.n341 B.n337 585
R247 B.n734 B.n733 585
R248 B.n733 B.n732 585
R249 B.n339 B.n338 585
R250 B.n340 B.n339 585
R251 B.n725 B.n724 585
R252 B.n726 B.n725 585
R253 B.n723 B.n346 585
R254 B.n346 B.n345 585
R255 B.n722 B.n721 585
R256 B.n721 B.n720 585
R257 B.n348 B.n347 585
R258 B.n349 B.n348 585
R259 B.n713 B.n712 585
R260 B.n714 B.n713 585
R261 B.n711 B.n354 585
R262 B.n354 B.n353 585
R263 B.n710 B.n709 585
R264 B.n709 B.n708 585
R265 B.n356 B.n355 585
R266 B.n701 B.n356 585
R267 B.n700 B.n699 585
R268 B.n702 B.n700 585
R269 B.n698 B.n361 585
R270 B.n361 B.n360 585
R271 B.n697 B.n696 585
R272 B.n696 B.n695 585
R273 B.n363 B.n362 585
R274 B.n364 B.n363 585
R275 B.n688 B.n687 585
R276 B.n689 B.n688 585
R277 B.n686 B.n369 585
R278 B.n369 B.n368 585
R279 B.n685 B.n684 585
R280 B.n684 B.n683 585
R281 B.n371 B.n370 585
R282 B.n676 B.n371 585
R283 B.n675 B.n674 585
R284 B.n677 B.n675 585
R285 B.n673 B.n376 585
R286 B.n376 B.n375 585
R287 B.n672 B.n671 585
R288 B.n671 B.n670 585
R289 B.n378 B.n377 585
R290 B.n379 B.n378 585
R291 B.n663 B.n662 585
R292 B.n664 B.n663 585
R293 B.n382 B.n381 585
R294 B.n443 B.n441 585
R295 B.n444 B.n440 585
R296 B.n444 B.n383 585
R297 B.n447 B.n446 585
R298 B.n448 B.n439 585
R299 B.n450 B.n449 585
R300 B.n452 B.n438 585
R301 B.n455 B.n454 585
R302 B.n456 B.n437 585
R303 B.n458 B.n457 585
R304 B.n460 B.n436 585
R305 B.n463 B.n462 585
R306 B.n464 B.n435 585
R307 B.n466 B.n465 585
R308 B.n468 B.n434 585
R309 B.n471 B.n470 585
R310 B.n472 B.n433 585
R311 B.n474 B.n473 585
R312 B.n476 B.n432 585
R313 B.n479 B.n478 585
R314 B.n480 B.n431 585
R315 B.n482 B.n481 585
R316 B.n484 B.n430 585
R317 B.n487 B.n486 585
R318 B.n488 B.n429 585
R319 B.n490 B.n489 585
R320 B.n492 B.n428 585
R321 B.n495 B.n494 585
R322 B.n496 B.n427 585
R323 B.n498 B.n497 585
R324 B.n500 B.n426 585
R325 B.n503 B.n502 585
R326 B.n504 B.n425 585
R327 B.n506 B.n505 585
R328 B.n508 B.n424 585
R329 B.n511 B.n510 585
R330 B.n512 B.n423 585
R331 B.n514 B.n513 585
R332 B.n516 B.n422 585
R333 B.n519 B.n518 585
R334 B.n520 B.n421 585
R335 B.n522 B.n521 585
R336 B.n524 B.n420 585
R337 B.n527 B.n526 585
R338 B.n528 B.n419 585
R339 B.n530 B.n529 585
R340 B.n532 B.n418 585
R341 B.n535 B.n534 585
R342 B.n536 B.n417 585
R343 B.n541 B.n540 585
R344 B.n543 B.n416 585
R345 B.n546 B.n545 585
R346 B.n547 B.n415 585
R347 B.n549 B.n548 585
R348 B.n551 B.n414 585
R349 B.n554 B.n553 585
R350 B.n555 B.n413 585
R351 B.n557 B.n556 585
R352 B.n559 B.n412 585
R353 B.n562 B.n561 585
R354 B.n564 B.n409 585
R355 B.n566 B.n565 585
R356 B.n568 B.n408 585
R357 B.n571 B.n570 585
R358 B.n572 B.n407 585
R359 B.n574 B.n573 585
R360 B.n576 B.n406 585
R361 B.n579 B.n578 585
R362 B.n580 B.n405 585
R363 B.n582 B.n581 585
R364 B.n584 B.n404 585
R365 B.n587 B.n586 585
R366 B.n588 B.n403 585
R367 B.n590 B.n589 585
R368 B.n592 B.n402 585
R369 B.n595 B.n594 585
R370 B.n596 B.n401 585
R371 B.n598 B.n597 585
R372 B.n600 B.n400 585
R373 B.n603 B.n602 585
R374 B.n604 B.n399 585
R375 B.n606 B.n605 585
R376 B.n608 B.n398 585
R377 B.n611 B.n610 585
R378 B.n612 B.n397 585
R379 B.n614 B.n613 585
R380 B.n616 B.n396 585
R381 B.n619 B.n618 585
R382 B.n620 B.n395 585
R383 B.n622 B.n621 585
R384 B.n624 B.n394 585
R385 B.n627 B.n626 585
R386 B.n628 B.n393 585
R387 B.n630 B.n629 585
R388 B.n632 B.n392 585
R389 B.n635 B.n634 585
R390 B.n636 B.n391 585
R391 B.n638 B.n637 585
R392 B.n640 B.n390 585
R393 B.n643 B.n642 585
R394 B.n644 B.n389 585
R395 B.n646 B.n645 585
R396 B.n648 B.n388 585
R397 B.n651 B.n650 585
R398 B.n652 B.n387 585
R399 B.n654 B.n653 585
R400 B.n656 B.n386 585
R401 B.n657 B.n385 585
R402 B.n660 B.n659 585
R403 B.n661 B.n384 585
R404 B.n384 B.n383 585
R405 B.n666 B.n665 585
R406 B.n665 B.n664 585
R407 B.n667 B.n380 585
R408 B.n380 B.n379 585
R409 B.n669 B.n668 585
R410 B.n670 B.n669 585
R411 B.n374 B.n373 585
R412 B.n375 B.n374 585
R413 B.n679 B.n678 585
R414 B.n678 B.n677 585
R415 B.n680 B.n372 585
R416 B.n676 B.n372 585
R417 B.n682 B.n681 585
R418 B.n683 B.n682 585
R419 B.n367 B.n366 585
R420 B.n368 B.n367 585
R421 B.n691 B.n690 585
R422 B.n690 B.n689 585
R423 B.n692 B.n365 585
R424 B.n365 B.n364 585
R425 B.n694 B.n693 585
R426 B.n695 B.n694 585
R427 B.n359 B.n358 585
R428 B.n360 B.n359 585
R429 B.n704 B.n703 585
R430 B.n703 B.n702 585
R431 B.n705 B.n357 585
R432 B.n701 B.n357 585
R433 B.n707 B.n706 585
R434 B.n708 B.n707 585
R435 B.n352 B.n351 585
R436 B.n353 B.n352 585
R437 B.n716 B.n715 585
R438 B.n715 B.n714 585
R439 B.n717 B.n350 585
R440 B.n350 B.n349 585
R441 B.n719 B.n718 585
R442 B.n720 B.n719 585
R443 B.n344 B.n343 585
R444 B.n345 B.n344 585
R445 B.n728 B.n727 585
R446 B.n727 B.n726 585
R447 B.n729 B.n342 585
R448 B.n342 B.n340 585
R449 B.n731 B.n730 585
R450 B.n732 B.n731 585
R451 B.n336 B.n335 585
R452 B.n341 B.n336 585
R453 B.n741 B.n740 585
R454 B.n740 B.n739 585
R455 B.n742 B.n334 585
R456 B.n334 B.n333 585
R457 B.n744 B.n743 585
R458 B.n745 B.n744 585
R459 B.n2 B.n0 585
R460 B.n4 B.n2 585
R461 B.n3 B.n1 585
R462 B.n844 B.n3 585
R463 B.n842 B.n841 585
R464 B.n843 B.n842 585
R465 B.n840 B.n9 585
R466 B.n9 B.n8 585
R467 B.n839 B.n838 585
R468 B.n838 B.n837 585
R469 B.n11 B.n10 585
R470 B.n836 B.n11 585
R471 B.n834 B.n833 585
R472 B.n835 B.n834 585
R473 B.n832 B.n16 585
R474 B.n16 B.n15 585
R475 B.n831 B.n830 585
R476 B.n830 B.n829 585
R477 B.n18 B.n17 585
R478 B.n828 B.n18 585
R479 B.n826 B.n825 585
R480 B.n827 B.n826 585
R481 B.n824 B.n23 585
R482 B.n23 B.n22 585
R483 B.n823 B.n822 585
R484 B.n822 B.n821 585
R485 B.n25 B.n24 585
R486 B.n820 B.n25 585
R487 B.n818 B.n817 585
R488 B.n819 B.n818 585
R489 B.n816 B.n29 585
R490 B.n32 B.n29 585
R491 B.n815 B.n814 585
R492 B.n814 B.n813 585
R493 B.n31 B.n30 585
R494 B.n812 B.n31 585
R495 B.n810 B.n809 585
R496 B.n811 B.n810 585
R497 B.n808 B.n37 585
R498 B.n37 B.n36 585
R499 B.n807 B.n806 585
R500 B.n806 B.n805 585
R501 B.n39 B.n38 585
R502 B.n804 B.n39 585
R503 B.n802 B.n801 585
R504 B.n803 B.n802 585
R505 B.n800 B.n43 585
R506 B.n46 B.n43 585
R507 B.n799 B.n798 585
R508 B.n798 B.n797 585
R509 B.n45 B.n44 585
R510 B.n796 B.n45 585
R511 B.n794 B.n793 585
R512 B.n795 B.n794 585
R513 B.n792 B.n51 585
R514 B.n51 B.n50 585
R515 B.n791 B.n790 585
R516 B.n790 B.n789 585
R517 B.n847 B.n846 585
R518 B.n846 B.n845 585
R519 B.n665 B.n382 545.355
R520 B.n790 B.n53 545.355
R521 B.n663 B.n384 545.355
R522 B.n786 B.n54 545.355
R523 B.n410 B.t14 468.438
R524 B.n537 B.t10 468.438
R525 B.n113 B.t17 468.438
R526 B.n110 B.t6 468.438
R527 B.n788 B.n787 256.663
R528 B.n788 B.n108 256.663
R529 B.n788 B.n107 256.663
R530 B.n788 B.n106 256.663
R531 B.n788 B.n105 256.663
R532 B.n788 B.n104 256.663
R533 B.n788 B.n103 256.663
R534 B.n788 B.n102 256.663
R535 B.n788 B.n101 256.663
R536 B.n788 B.n100 256.663
R537 B.n788 B.n99 256.663
R538 B.n788 B.n98 256.663
R539 B.n788 B.n97 256.663
R540 B.n788 B.n96 256.663
R541 B.n788 B.n95 256.663
R542 B.n788 B.n94 256.663
R543 B.n788 B.n93 256.663
R544 B.n788 B.n92 256.663
R545 B.n788 B.n91 256.663
R546 B.n788 B.n90 256.663
R547 B.n788 B.n89 256.663
R548 B.n788 B.n88 256.663
R549 B.n788 B.n87 256.663
R550 B.n788 B.n86 256.663
R551 B.n788 B.n85 256.663
R552 B.n788 B.n84 256.663
R553 B.n788 B.n83 256.663
R554 B.n788 B.n82 256.663
R555 B.n788 B.n81 256.663
R556 B.n788 B.n80 256.663
R557 B.n788 B.n79 256.663
R558 B.n788 B.n78 256.663
R559 B.n788 B.n77 256.663
R560 B.n788 B.n76 256.663
R561 B.n788 B.n75 256.663
R562 B.n788 B.n74 256.663
R563 B.n788 B.n73 256.663
R564 B.n788 B.n72 256.663
R565 B.n788 B.n71 256.663
R566 B.n788 B.n70 256.663
R567 B.n788 B.n69 256.663
R568 B.n788 B.n68 256.663
R569 B.n788 B.n67 256.663
R570 B.n788 B.n66 256.663
R571 B.n788 B.n65 256.663
R572 B.n788 B.n64 256.663
R573 B.n788 B.n63 256.663
R574 B.n788 B.n62 256.663
R575 B.n788 B.n61 256.663
R576 B.n788 B.n60 256.663
R577 B.n788 B.n59 256.663
R578 B.n788 B.n58 256.663
R579 B.n788 B.n57 256.663
R580 B.n788 B.n56 256.663
R581 B.n788 B.n55 256.663
R582 B.n442 B.n383 256.663
R583 B.n445 B.n383 256.663
R584 B.n451 B.n383 256.663
R585 B.n453 B.n383 256.663
R586 B.n459 B.n383 256.663
R587 B.n461 B.n383 256.663
R588 B.n467 B.n383 256.663
R589 B.n469 B.n383 256.663
R590 B.n475 B.n383 256.663
R591 B.n477 B.n383 256.663
R592 B.n483 B.n383 256.663
R593 B.n485 B.n383 256.663
R594 B.n491 B.n383 256.663
R595 B.n493 B.n383 256.663
R596 B.n499 B.n383 256.663
R597 B.n501 B.n383 256.663
R598 B.n507 B.n383 256.663
R599 B.n509 B.n383 256.663
R600 B.n515 B.n383 256.663
R601 B.n517 B.n383 256.663
R602 B.n523 B.n383 256.663
R603 B.n525 B.n383 256.663
R604 B.n531 B.n383 256.663
R605 B.n533 B.n383 256.663
R606 B.n542 B.n383 256.663
R607 B.n544 B.n383 256.663
R608 B.n550 B.n383 256.663
R609 B.n552 B.n383 256.663
R610 B.n558 B.n383 256.663
R611 B.n560 B.n383 256.663
R612 B.n567 B.n383 256.663
R613 B.n569 B.n383 256.663
R614 B.n575 B.n383 256.663
R615 B.n577 B.n383 256.663
R616 B.n583 B.n383 256.663
R617 B.n585 B.n383 256.663
R618 B.n591 B.n383 256.663
R619 B.n593 B.n383 256.663
R620 B.n599 B.n383 256.663
R621 B.n601 B.n383 256.663
R622 B.n607 B.n383 256.663
R623 B.n609 B.n383 256.663
R624 B.n615 B.n383 256.663
R625 B.n617 B.n383 256.663
R626 B.n623 B.n383 256.663
R627 B.n625 B.n383 256.663
R628 B.n631 B.n383 256.663
R629 B.n633 B.n383 256.663
R630 B.n639 B.n383 256.663
R631 B.n641 B.n383 256.663
R632 B.n647 B.n383 256.663
R633 B.n649 B.n383 256.663
R634 B.n655 B.n383 256.663
R635 B.n658 B.n383 256.663
R636 B.n665 B.n380 163.367
R637 B.n669 B.n380 163.367
R638 B.n669 B.n374 163.367
R639 B.n678 B.n374 163.367
R640 B.n678 B.n372 163.367
R641 B.n682 B.n372 163.367
R642 B.n682 B.n367 163.367
R643 B.n690 B.n367 163.367
R644 B.n690 B.n365 163.367
R645 B.n694 B.n365 163.367
R646 B.n694 B.n359 163.367
R647 B.n703 B.n359 163.367
R648 B.n703 B.n357 163.367
R649 B.n707 B.n357 163.367
R650 B.n707 B.n352 163.367
R651 B.n715 B.n352 163.367
R652 B.n715 B.n350 163.367
R653 B.n719 B.n350 163.367
R654 B.n719 B.n344 163.367
R655 B.n727 B.n344 163.367
R656 B.n727 B.n342 163.367
R657 B.n731 B.n342 163.367
R658 B.n731 B.n336 163.367
R659 B.n740 B.n336 163.367
R660 B.n740 B.n334 163.367
R661 B.n744 B.n334 163.367
R662 B.n744 B.n2 163.367
R663 B.n846 B.n2 163.367
R664 B.n846 B.n3 163.367
R665 B.n842 B.n3 163.367
R666 B.n842 B.n9 163.367
R667 B.n838 B.n9 163.367
R668 B.n838 B.n11 163.367
R669 B.n834 B.n11 163.367
R670 B.n834 B.n16 163.367
R671 B.n830 B.n16 163.367
R672 B.n830 B.n18 163.367
R673 B.n826 B.n18 163.367
R674 B.n826 B.n23 163.367
R675 B.n822 B.n23 163.367
R676 B.n822 B.n25 163.367
R677 B.n818 B.n25 163.367
R678 B.n818 B.n29 163.367
R679 B.n814 B.n29 163.367
R680 B.n814 B.n31 163.367
R681 B.n810 B.n31 163.367
R682 B.n810 B.n37 163.367
R683 B.n806 B.n37 163.367
R684 B.n806 B.n39 163.367
R685 B.n802 B.n39 163.367
R686 B.n802 B.n43 163.367
R687 B.n798 B.n43 163.367
R688 B.n798 B.n45 163.367
R689 B.n794 B.n45 163.367
R690 B.n794 B.n51 163.367
R691 B.n790 B.n51 163.367
R692 B.n444 B.n443 163.367
R693 B.n446 B.n444 163.367
R694 B.n450 B.n439 163.367
R695 B.n454 B.n452 163.367
R696 B.n458 B.n437 163.367
R697 B.n462 B.n460 163.367
R698 B.n466 B.n435 163.367
R699 B.n470 B.n468 163.367
R700 B.n474 B.n433 163.367
R701 B.n478 B.n476 163.367
R702 B.n482 B.n431 163.367
R703 B.n486 B.n484 163.367
R704 B.n490 B.n429 163.367
R705 B.n494 B.n492 163.367
R706 B.n498 B.n427 163.367
R707 B.n502 B.n500 163.367
R708 B.n506 B.n425 163.367
R709 B.n510 B.n508 163.367
R710 B.n514 B.n423 163.367
R711 B.n518 B.n516 163.367
R712 B.n522 B.n421 163.367
R713 B.n526 B.n524 163.367
R714 B.n530 B.n419 163.367
R715 B.n534 B.n532 163.367
R716 B.n541 B.n417 163.367
R717 B.n545 B.n543 163.367
R718 B.n549 B.n415 163.367
R719 B.n553 B.n551 163.367
R720 B.n557 B.n413 163.367
R721 B.n561 B.n559 163.367
R722 B.n566 B.n409 163.367
R723 B.n570 B.n568 163.367
R724 B.n574 B.n407 163.367
R725 B.n578 B.n576 163.367
R726 B.n582 B.n405 163.367
R727 B.n586 B.n584 163.367
R728 B.n590 B.n403 163.367
R729 B.n594 B.n592 163.367
R730 B.n598 B.n401 163.367
R731 B.n602 B.n600 163.367
R732 B.n606 B.n399 163.367
R733 B.n610 B.n608 163.367
R734 B.n614 B.n397 163.367
R735 B.n618 B.n616 163.367
R736 B.n622 B.n395 163.367
R737 B.n626 B.n624 163.367
R738 B.n630 B.n393 163.367
R739 B.n634 B.n632 163.367
R740 B.n638 B.n391 163.367
R741 B.n642 B.n640 163.367
R742 B.n646 B.n389 163.367
R743 B.n650 B.n648 163.367
R744 B.n654 B.n387 163.367
R745 B.n657 B.n656 163.367
R746 B.n659 B.n384 163.367
R747 B.n663 B.n378 163.367
R748 B.n671 B.n378 163.367
R749 B.n671 B.n376 163.367
R750 B.n675 B.n376 163.367
R751 B.n675 B.n371 163.367
R752 B.n684 B.n371 163.367
R753 B.n684 B.n369 163.367
R754 B.n688 B.n369 163.367
R755 B.n688 B.n363 163.367
R756 B.n696 B.n363 163.367
R757 B.n696 B.n361 163.367
R758 B.n700 B.n361 163.367
R759 B.n700 B.n356 163.367
R760 B.n709 B.n356 163.367
R761 B.n709 B.n354 163.367
R762 B.n713 B.n354 163.367
R763 B.n713 B.n348 163.367
R764 B.n721 B.n348 163.367
R765 B.n721 B.n346 163.367
R766 B.n725 B.n346 163.367
R767 B.n725 B.n339 163.367
R768 B.n733 B.n339 163.367
R769 B.n733 B.n337 163.367
R770 B.n738 B.n337 163.367
R771 B.n738 B.n332 163.367
R772 B.n746 B.n332 163.367
R773 B.n747 B.n746 163.367
R774 B.n747 B.n5 163.367
R775 B.n6 B.n5 163.367
R776 B.n7 B.n6 163.367
R777 B.n752 B.n7 163.367
R778 B.n752 B.n12 163.367
R779 B.n13 B.n12 163.367
R780 B.n14 B.n13 163.367
R781 B.n757 B.n14 163.367
R782 B.n757 B.n19 163.367
R783 B.n20 B.n19 163.367
R784 B.n21 B.n20 163.367
R785 B.n762 B.n21 163.367
R786 B.n762 B.n26 163.367
R787 B.n27 B.n26 163.367
R788 B.n28 B.n27 163.367
R789 B.n767 B.n28 163.367
R790 B.n767 B.n33 163.367
R791 B.n34 B.n33 163.367
R792 B.n35 B.n34 163.367
R793 B.n772 B.n35 163.367
R794 B.n772 B.n40 163.367
R795 B.n41 B.n40 163.367
R796 B.n42 B.n41 163.367
R797 B.n777 B.n42 163.367
R798 B.n777 B.n47 163.367
R799 B.n48 B.n47 163.367
R800 B.n49 B.n48 163.367
R801 B.n782 B.n49 163.367
R802 B.n782 B.n54 163.367
R803 B.n118 B.n117 163.367
R804 B.n122 B.n121 163.367
R805 B.n126 B.n125 163.367
R806 B.n130 B.n129 163.367
R807 B.n134 B.n133 163.367
R808 B.n138 B.n137 163.367
R809 B.n142 B.n141 163.367
R810 B.n146 B.n145 163.367
R811 B.n150 B.n149 163.367
R812 B.n154 B.n153 163.367
R813 B.n158 B.n157 163.367
R814 B.n162 B.n161 163.367
R815 B.n166 B.n165 163.367
R816 B.n170 B.n169 163.367
R817 B.n174 B.n173 163.367
R818 B.n178 B.n177 163.367
R819 B.n182 B.n181 163.367
R820 B.n186 B.n185 163.367
R821 B.n190 B.n189 163.367
R822 B.n194 B.n193 163.367
R823 B.n198 B.n197 163.367
R824 B.n202 B.n201 163.367
R825 B.n206 B.n205 163.367
R826 B.n210 B.n209 163.367
R827 B.n214 B.n213 163.367
R828 B.n218 B.n217 163.367
R829 B.n222 B.n221 163.367
R830 B.n226 B.n225 163.367
R831 B.n230 B.n229 163.367
R832 B.n234 B.n233 163.367
R833 B.n238 B.n237 163.367
R834 B.n242 B.n241 163.367
R835 B.n246 B.n245 163.367
R836 B.n250 B.n249 163.367
R837 B.n254 B.n253 163.367
R838 B.n258 B.n257 163.367
R839 B.n262 B.n261 163.367
R840 B.n266 B.n265 163.367
R841 B.n270 B.n269 163.367
R842 B.n274 B.n273 163.367
R843 B.n278 B.n277 163.367
R844 B.n282 B.n281 163.367
R845 B.n286 B.n285 163.367
R846 B.n290 B.n289 163.367
R847 B.n294 B.n293 163.367
R848 B.n298 B.n297 163.367
R849 B.n302 B.n301 163.367
R850 B.n306 B.n305 163.367
R851 B.n310 B.n309 163.367
R852 B.n314 B.n313 163.367
R853 B.n318 B.n317 163.367
R854 B.n322 B.n321 163.367
R855 B.n326 B.n325 163.367
R856 B.n328 B.n109 163.367
R857 B.n410 B.t16 100.823
R858 B.n110 B.t8 100.823
R859 B.n537 B.t13 100.803
R860 B.n113 B.t18 100.803
R861 B.n442 B.n382 71.676
R862 B.n446 B.n445 71.676
R863 B.n451 B.n450 71.676
R864 B.n454 B.n453 71.676
R865 B.n459 B.n458 71.676
R866 B.n462 B.n461 71.676
R867 B.n467 B.n466 71.676
R868 B.n470 B.n469 71.676
R869 B.n475 B.n474 71.676
R870 B.n478 B.n477 71.676
R871 B.n483 B.n482 71.676
R872 B.n486 B.n485 71.676
R873 B.n491 B.n490 71.676
R874 B.n494 B.n493 71.676
R875 B.n499 B.n498 71.676
R876 B.n502 B.n501 71.676
R877 B.n507 B.n506 71.676
R878 B.n510 B.n509 71.676
R879 B.n515 B.n514 71.676
R880 B.n518 B.n517 71.676
R881 B.n523 B.n522 71.676
R882 B.n526 B.n525 71.676
R883 B.n531 B.n530 71.676
R884 B.n534 B.n533 71.676
R885 B.n542 B.n541 71.676
R886 B.n545 B.n544 71.676
R887 B.n550 B.n549 71.676
R888 B.n553 B.n552 71.676
R889 B.n558 B.n557 71.676
R890 B.n561 B.n560 71.676
R891 B.n567 B.n566 71.676
R892 B.n570 B.n569 71.676
R893 B.n575 B.n574 71.676
R894 B.n578 B.n577 71.676
R895 B.n583 B.n582 71.676
R896 B.n586 B.n585 71.676
R897 B.n591 B.n590 71.676
R898 B.n594 B.n593 71.676
R899 B.n599 B.n598 71.676
R900 B.n602 B.n601 71.676
R901 B.n607 B.n606 71.676
R902 B.n610 B.n609 71.676
R903 B.n615 B.n614 71.676
R904 B.n618 B.n617 71.676
R905 B.n623 B.n622 71.676
R906 B.n626 B.n625 71.676
R907 B.n631 B.n630 71.676
R908 B.n634 B.n633 71.676
R909 B.n639 B.n638 71.676
R910 B.n642 B.n641 71.676
R911 B.n647 B.n646 71.676
R912 B.n650 B.n649 71.676
R913 B.n655 B.n654 71.676
R914 B.n658 B.n657 71.676
R915 B.n55 B.n53 71.676
R916 B.n118 B.n56 71.676
R917 B.n122 B.n57 71.676
R918 B.n126 B.n58 71.676
R919 B.n130 B.n59 71.676
R920 B.n134 B.n60 71.676
R921 B.n138 B.n61 71.676
R922 B.n142 B.n62 71.676
R923 B.n146 B.n63 71.676
R924 B.n150 B.n64 71.676
R925 B.n154 B.n65 71.676
R926 B.n158 B.n66 71.676
R927 B.n162 B.n67 71.676
R928 B.n166 B.n68 71.676
R929 B.n170 B.n69 71.676
R930 B.n174 B.n70 71.676
R931 B.n178 B.n71 71.676
R932 B.n182 B.n72 71.676
R933 B.n186 B.n73 71.676
R934 B.n190 B.n74 71.676
R935 B.n194 B.n75 71.676
R936 B.n198 B.n76 71.676
R937 B.n202 B.n77 71.676
R938 B.n206 B.n78 71.676
R939 B.n210 B.n79 71.676
R940 B.n214 B.n80 71.676
R941 B.n218 B.n81 71.676
R942 B.n222 B.n82 71.676
R943 B.n226 B.n83 71.676
R944 B.n230 B.n84 71.676
R945 B.n234 B.n85 71.676
R946 B.n238 B.n86 71.676
R947 B.n242 B.n87 71.676
R948 B.n246 B.n88 71.676
R949 B.n250 B.n89 71.676
R950 B.n254 B.n90 71.676
R951 B.n258 B.n91 71.676
R952 B.n262 B.n92 71.676
R953 B.n266 B.n93 71.676
R954 B.n270 B.n94 71.676
R955 B.n274 B.n95 71.676
R956 B.n278 B.n96 71.676
R957 B.n282 B.n97 71.676
R958 B.n286 B.n98 71.676
R959 B.n290 B.n99 71.676
R960 B.n294 B.n100 71.676
R961 B.n298 B.n101 71.676
R962 B.n302 B.n102 71.676
R963 B.n306 B.n103 71.676
R964 B.n310 B.n104 71.676
R965 B.n314 B.n105 71.676
R966 B.n318 B.n106 71.676
R967 B.n322 B.n107 71.676
R968 B.n326 B.n108 71.676
R969 B.n787 B.n109 71.676
R970 B.n787 B.n786 71.676
R971 B.n328 B.n108 71.676
R972 B.n325 B.n107 71.676
R973 B.n321 B.n106 71.676
R974 B.n317 B.n105 71.676
R975 B.n313 B.n104 71.676
R976 B.n309 B.n103 71.676
R977 B.n305 B.n102 71.676
R978 B.n301 B.n101 71.676
R979 B.n297 B.n100 71.676
R980 B.n293 B.n99 71.676
R981 B.n289 B.n98 71.676
R982 B.n285 B.n97 71.676
R983 B.n281 B.n96 71.676
R984 B.n277 B.n95 71.676
R985 B.n273 B.n94 71.676
R986 B.n269 B.n93 71.676
R987 B.n265 B.n92 71.676
R988 B.n261 B.n91 71.676
R989 B.n257 B.n90 71.676
R990 B.n253 B.n89 71.676
R991 B.n249 B.n88 71.676
R992 B.n245 B.n87 71.676
R993 B.n241 B.n86 71.676
R994 B.n237 B.n85 71.676
R995 B.n233 B.n84 71.676
R996 B.n229 B.n83 71.676
R997 B.n225 B.n82 71.676
R998 B.n221 B.n81 71.676
R999 B.n217 B.n80 71.676
R1000 B.n213 B.n79 71.676
R1001 B.n209 B.n78 71.676
R1002 B.n205 B.n77 71.676
R1003 B.n201 B.n76 71.676
R1004 B.n197 B.n75 71.676
R1005 B.n193 B.n74 71.676
R1006 B.n189 B.n73 71.676
R1007 B.n185 B.n72 71.676
R1008 B.n181 B.n71 71.676
R1009 B.n177 B.n70 71.676
R1010 B.n173 B.n69 71.676
R1011 B.n169 B.n68 71.676
R1012 B.n165 B.n67 71.676
R1013 B.n161 B.n66 71.676
R1014 B.n157 B.n65 71.676
R1015 B.n153 B.n64 71.676
R1016 B.n149 B.n63 71.676
R1017 B.n145 B.n62 71.676
R1018 B.n141 B.n61 71.676
R1019 B.n137 B.n60 71.676
R1020 B.n133 B.n59 71.676
R1021 B.n129 B.n58 71.676
R1022 B.n125 B.n57 71.676
R1023 B.n121 B.n56 71.676
R1024 B.n117 B.n55 71.676
R1025 B.n443 B.n442 71.676
R1026 B.n445 B.n439 71.676
R1027 B.n452 B.n451 71.676
R1028 B.n453 B.n437 71.676
R1029 B.n460 B.n459 71.676
R1030 B.n461 B.n435 71.676
R1031 B.n468 B.n467 71.676
R1032 B.n469 B.n433 71.676
R1033 B.n476 B.n475 71.676
R1034 B.n477 B.n431 71.676
R1035 B.n484 B.n483 71.676
R1036 B.n485 B.n429 71.676
R1037 B.n492 B.n491 71.676
R1038 B.n493 B.n427 71.676
R1039 B.n500 B.n499 71.676
R1040 B.n501 B.n425 71.676
R1041 B.n508 B.n507 71.676
R1042 B.n509 B.n423 71.676
R1043 B.n516 B.n515 71.676
R1044 B.n517 B.n421 71.676
R1045 B.n524 B.n523 71.676
R1046 B.n525 B.n419 71.676
R1047 B.n532 B.n531 71.676
R1048 B.n533 B.n417 71.676
R1049 B.n543 B.n542 71.676
R1050 B.n544 B.n415 71.676
R1051 B.n551 B.n550 71.676
R1052 B.n552 B.n413 71.676
R1053 B.n559 B.n558 71.676
R1054 B.n560 B.n409 71.676
R1055 B.n568 B.n567 71.676
R1056 B.n569 B.n407 71.676
R1057 B.n576 B.n575 71.676
R1058 B.n577 B.n405 71.676
R1059 B.n584 B.n583 71.676
R1060 B.n585 B.n403 71.676
R1061 B.n592 B.n591 71.676
R1062 B.n593 B.n401 71.676
R1063 B.n600 B.n599 71.676
R1064 B.n601 B.n399 71.676
R1065 B.n608 B.n607 71.676
R1066 B.n609 B.n397 71.676
R1067 B.n616 B.n615 71.676
R1068 B.n617 B.n395 71.676
R1069 B.n624 B.n623 71.676
R1070 B.n625 B.n393 71.676
R1071 B.n632 B.n631 71.676
R1072 B.n633 B.n391 71.676
R1073 B.n640 B.n639 71.676
R1074 B.n641 B.n389 71.676
R1075 B.n648 B.n647 71.676
R1076 B.n649 B.n387 71.676
R1077 B.n656 B.n655 71.676
R1078 B.n659 B.n658 71.676
R1079 B.n664 B.n383 71.1434
R1080 B.n789 B.n788 71.1434
R1081 B.n411 B.t15 67.854
R1082 B.n111 B.t9 67.854
R1083 B.n538 B.t12 67.8343
R1084 B.n114 B.t19 67.8343
R1085 B.n563 B.n411 59.5399
R1086 B.n539 B.n538 59.5399
R1087 B.n115 B.n114 59.5399
R1088 B.n112 B.n111 59.5399
R1089 B.n664 B.n379 36.9297
R1090 B.n670 B.n379 36.9297
R1091 B.n670 B.n375 36.9297
R1092 B.n677 B.n375 36.9297
R1093 B.n677 B.n676 36.9297
R1094 B.n683 B.n368 36.9297
R1095 B.n689 B.n368 36.9297
R1096 B.n689 B.n364 36.9297
R1097 B.n695 B.n364 36.9297
R1098 B.n695 B.n360 36.9297
R1099 B.n702 B.n360 36.9297
R1100 B.n702 B.n701 36.9297
R1101 B.n708 B.n353 36.9297
R1102 B.n714 B.n353 36.9297
R1103 B.n714 B.n349 36.9297
R1104 B.n720 B.n349 36.9297
R1105 B.n726 B.n345 36.9297
R1106 B.n726 B.n340 36.9297
R1107 B.n732 B.n340 36.9297
R1108 B.n732 B.n341 36.9297
R1109 B.n739 B.n333 36.9297
R1110 B.n745 B.n333 36.9297
R1111 B.n745 B.n4 36.9297
R1112 B.n845 B.n4 36.9297
R1113 B.n845 B.n844 36.9297
R1114 B.n844 B.n843 36.9297
R1115 B.n843 B.n8 36.9297
R1116 B.n837 B.n8 36.9297
R1117 B.n836 B.n835 36.9297
R1118 B.n835 B.n15 36.9297
R1119 B.n829 B.n15 36.9297
R1120 B.n829 B.n828 36.9297
R1121 B.n827 B.n22 36.9297
R1122 B.n821 B.n22 36.9297
R1123 B.n821 B.n820 36.9297
R1124 B.n820 B.n819 36.9297
R1125 B.n813 B.n32 36.9297
R1126 B.n813 B.n812 36.9297
R1127 B.n812 B.n811 36.9297
R1128 B.n811 B.n36 36.9297
R1129 B.n805 B.n36 36.9297
R1130 B.n805 B.n804 36.9297
R1131 B.n804 B.n803 36.9297
R1132 B.n797 B.n46 36.9297
R1133 B.n797 B.n796 36.9297
R1134 B.n796 B.n795 36.9297
R1135 B.n795 B.n50 36.9297
R1136 B.n789 B.n50 36.9297
R1137 B.n791 B.n52 35.4346
R1138 B.n662 B.n661 35.4346
R1139 B.n666 B.n381 35.4346
R1140 B.n785 B.n784 35.4346
R1141 B.n701 B.t1 33.1281
R1142 B.n720 B.t4 33.1281
R1143 B.n341 B.t0 33.1281
R1144 B.t3 B.n836 33.1281
R1145 B.t5 B.n827 33.1281
R1146 B.n32 B.t2 33.1281
R1147 B.n411 B.n410 32.9702
R1148 B.n538 B.n537 32.9702
R1149 B.n114 B.n113 32.9702
R1150 B.n111 B.n110 32.9702
R1151 B.n676 B.t11 25.5251
R1152 B.n46 B.t7 25.5251
R1153 B B.n847 18.0485
R1154 B.n683 B.t11 11.4051
R1155 B.n803 B.t7 11.4051
R1156 B.n116 B.n52 10.6151
R1157 B.n119 B.n116 10.6151
R1158 B.n120 B.n119 10.6151
R1159 B.n123 B.n120 10.6151
R1160 B.n124 B.n123 10.6151
R1161 B.n127 B.n124 10.6151
R1162 B.n128 B.n127 10.6151
R1163 B.n131 B.n128 10.6151
R1164 B.n132 B.n131 10.6151
R1165 B.n135 B.n132 10.6151
R1166 B.n136 B.n135 10.6151
R1167 B.n139 B.n136 10.6151
R1168 B.n140 B.n139 10.6151
R1169 B.n143 B.n140 10.6151
R1170 B.n144 B.n143 10.6151
R1171 B.n147 B.n144 10.6151
R1172 B.n148 B.n147 10.6151
R1173 B.n151 B.n148 10.6151
R1174 B.n152 B.n151 10.6151
R1175 B.n155 B.n152 10.6151
R1176 B.n156 B.n155 10.6151
R1177 B.n159 B.n156 10.6151
R1178 B.n160 B.n159 10.6151
R1179 B.n163 B.n160 10.6151
R1180 B.n164 B.n163 10.6151
R1181 B.n167 B.n164 10.6151
R1182 B.n168 B.n167 10.6151
R1183 B.n171 B.n168 10.6151
R1184 B.n172 B.n171 10.6151
R1185 B.n175 B.n172 10.6151
R1186 B.n176 B.n175 10.6151
R1187 B.n179 B.n176 10.6151
R1188 B.n180 B.n179 10.6151
R1189 B.n183 B.n180 10.6151
R1190 B.n184 B.n183 10.6151
R1191 B.n187 B.n184 10.6151
R1192 B.n188 B.n187 10.6151
R1193 B.n191 B.n188 10.6151
R1194 B.n192 B.n191 10.6151
R1195 B.n195 B.n192 10.6151
R1196 B.n196 B.n195 10.6151
R1197 B.n199 B.n196 10.6151
R1198 B.n200 B.n199 10.6151
R1199 B.n203 B.n200 10.6151
R1200 B.n204 B.n203 10.6151
R1201 B.n207 B.n204 10.6151
R1202 B.n208 B.n207 10.6151
R1203 B.n211 B.n208 10.6151
R1204 B.n212 B.n211 10.6151
R1205 B.n216 B.n215 10.6151
R1206 B.n219 B.n216 10.6151
R1207 B.n220 B.n219 10.6151
R1208 B.n223 B.n220 10.6151
R1209 B.n224 B.n223 10.6151
R1210 B.n227 B.n224 10.6151
R1211 B.n228 B.n227 10.6151
R1212 B.n231 B.n228 10.6151
R1213 B.n232 B.n231 10.6151
R1214 B.n236 B.n235 10.6151
R1215 B.n239 B.n236 10.6151
R1216 B.n240 B.n239 10.6151
R1217 B.n243 B.n240 10.6151
R1218 B.n244 B.n243 10.6151
R1219 B.n247 B.n244 10.6151
R1220 B.n248 B.n247 10.6151
R1221 B.n251 B.n248 10.6151
R1222 B.n252 B.n251 10.6151
R1223 B.n255 B.n252 10.6151
R1224 B.n256 B.n255 10.6151
R1225 B.n259 B.n256 10.6151
R1226 B.n260 B.n259 10.6151
R1227 B.n263 B.n260 10.6151
R1228 B.n264 B.n263 10.6151
R1229 B.n267 B.n264 10.6151
R1230 B.n268 B.n267 10.6151
R1231 B.n271 B.n268 10.6151
R1232 B.n272 B.n271 10.6151
R1233 B.n275 B.n272 10.6151
R1234 B.n276 B.n275 10.6151
R1235 B.n279 B.n276 10.6151
R1236 B.n280 B.n279 10.6151
R1237 B.n283 B.n280 10.6151
R1238 B.n284 B.n283 10.6151
R1239 B.n287 B.n284 10.6151
R1240 B.n288 B.n287 10.6151
R1241 B.n291 B.n288 10.6151
R1242 B.n292 B.n291 10.6151
R1243 B.n295 B.n292 10.6151
R1244 B.n296 B.n295 10.6151
R1245 B.n299 B.n296 10.6151
R1246 B.n300 B.n299 10.6151
R1247 B.n303 B.n300 10.6151
R1248 B.n304 B.n303 10.6151
R1249 B.n307 B.n304 10.6151
R1250 B.n308 B.n307 10.6151
R1251 B.n311 B.n308 10.6151
R1252 B.n312 B.n311 10.6151
R1253 B.n315 B.n312 10.6151
R1254 B.n316 B.n315 10.6151
R1255 B.n319 B.n316 10.6151
R1256 B.n320 B.n319 10.6151
R1257 B.n323 B.n320 10.6151
R1258 B.n324 B.n323 10.6151
R1259 B.n327 B.n324 10.6151
R1260 B.n329 B.n327 10.6151
R1261 B.n330 B.n329 10.6151
R1262 B.n785 B.n330 10.6151
R1263 B.n662 B.n377 10.6151
R1264 B.n672 B.n377 10.6151
R1265 B.n673 B.n672 10.6151
R1266 B.n674 B.n673 10.6151
R1267 B.n674 B.n370 10.6151
R1268 B.n685 B.n370 10.6151
R1269 B.n686 B.n685 10.6151
R1270 B.n687 B.n686 10.6151
R1271 B.n687 B.n362 10.6151
R1272 B.n697 B.n362 10.6151
R1273 B.n698 B.n697 10.6151
R1274 B.n699 B.n698 10.6151
R1275 B.n699 B.n355 10.6151
R1276 B.n710 B.n355 10.6151
R1277 B.n711 B.n710 10.6151
R1278 B.n712 B.n711 10.6151
R1279 B.n712 B.n347 10.6151
R1280 B.n722 B.n347 10.6151
R1281 B.n723 B.n722 10.6151
R1282 B.n724 B.n723 10.6151
R1283 B.n724 B.n338 10.6151
R1284 B.n734 B.n338 10.6151
R1285 B.n735 B.n734 10.6151
R1286 B.n737 B.n735 10.6151
R1287 B.n737 B.n736 10.6151
R1288 B.n736 B.n331 10.6151
R1289 B.n748 B.n331 10.6151
R1290 B.n749 B.n748 10.6151
R1291 B.n750 B.n749 10.6151
R1292 B.n751 B.n750 10.6151
R1293 B.n753 B.n751 10.6151
R1294 B.n754 B.n753 10.6151
R1295 B.n755 B.n754 10.6151
R1296 B.n756 B.n755 10.6151
R1297 B.n758 B.n756 10.6151
R1298 B.n759 B.n758 10.6151
R1299 B.n760 B.n759 10.6151
R1300 B.n761 B.n760 10.6151
R1301 B.n763 B.n761 10.6151
R1302 B.n764 B.n763 10.6151
R1303 B.n765 B.n764 10.6151
R1304 B.n766 B.n765 10.6151
R1305 B.n768 B.n766 10.6151
R1306 B.n769 B.n768 10.6151
R1307 B.n770 B.n769 10.6151
R1308 B.n771 B.n770 10.6151
R1309 B.n773 B.n771 10.6151
R1310 B.n774 B.n773 10.6151
R1311 B.n775 B.n774 10.6151
R1312 B.n776 B.n775 10.6151
R1313 B.n778 B.n776 10.6151
R1314 B.n779 B.n778 10.6151
R1315 B.n780 B.n779 10.6151
R1316 B.n781 B.n780 10.6151
R1317 B.n783 B.n781 10.6151
R1318 B.n784 B.n783 10.6151
R1319 B.n441 B.n381 10.6151
R1320 B.n441 B.n440 10.6151
R1321 B.n447 B.n440 10.6151
R1322 B.n448 B.n447 10.6151
R1323 B.n449 B.n448 10.6151
R1324 B.n449 B.n438 10.6151
R1325 B.n455 B.n438 10.6151
R1326 B.n456 B.n455 10.6151
R1327 B.n457 B.n456 10.6151
R1328 B.n457 B.n436 10.6151
R1329 B.n463 B.n436 10.6151
R1330 B.n464 B.n463 10.6151
R1331 B.n465 B.n464 10.6151
R1332 B.n465 B.n434 10.6151
R1333 B.n471 B.n434 10.6151
R1334 B.n472 B.n471 10.6151
R1335 B.n473 B.n472 10.6151
R1336 B.n473 B.n432 10.6151
R1337 B.n479 B.n432 10.6151
R1338 B.n480 B.n479 10.6151
R1339 B.n481 B.n480 10.6151
R1340 B.n481 B.n430 10.6151
R1341 B.n487 B.n430 10.6151
R1342 B.n488 B.n487 10.6151
R1343 B.n489 B.n488 10.6151
R1344 B.n489 B.n428 10.6151
R1345 B.n495 B.n428 10.6151
R1346 B.n496 B.n495 10.6151
R1347 B.n497 B.n496 10.6151
R1348 B.n497 B.n426 10.6151
R1349 B.n503 B.n426 10.6151
R1350 B.n504 B.n503 10.6151
R1351 B.n505 B.n504 10.6151
R1352 B.n505 B.n424 10.6151
R1353 B.n511 B.n424 10.6151
R1354 B.n512 B.n511 10.6151
R1355 B.n513 B.n512 10.6151
R1356 B.n513 B.n422 10.6151
R1357 B.n519 B.n422 10.6151
R1358 B.n520 B.n519 10.6151
R1359 B.n521 B.n520 10.6151
R1360 B.n521 B.n420 10.6151
R1361 B.n527 B.n420 10.6151
R1362 B.n528 B.n527 10.6151
R1363 B.n529 B.n528 10.6151
R1364 B.n529 B.n418 10.6151
R1365 B.n535 B.n418 10.6151
R1366 B.n536 B.n535 10.6151
R1367 B.n540 B.n536 10.6151
R1368 B.n546 B.n416 10.6151
R1369 B.n547 B.n546 10.6151
R1370 B.n548 B.n547 10.6151
R1371 B.n548 B.n414 10.6151
R1372 B.n554 B.n414 10.6151
R1373 B.n555 B.n554 10.6151
R1374 B.n556 B.n555 10.6151
R1375 B.n556 B.n412 10.6151
R1376 B.n562 B.n412 10.6151
R1377 B.n565 B.n564 10.6151
R1378 B.n565 B.n408 10.6151
R1379 B.n571 B.n408 10.6151
R1380 B.n572 B.n571 10.6151
R1381 B.n573 B.n572 10.6151
R1382 B.n573 B.n406 10.6151
R1383 B.n579 B.n406 10.6151
R1384 B.n580 B.n579 10.6151
R1385 B.n581 B.n580 10.6151
R1386 B.n581 B.n404 10.6151
R1387 B.n587 B.n404 10.6151
R1388 B.n588 B.n587 10.6151
R1389 B.n589 B.n588 10.6151
R1390 B.n589 B.n402 10.6151
R1391 B.n595 B.n402 10.6151
R1392 B.n596 B.n595 10.6151
R1393 B.n597 B.n596 10.6151
R1394 B.n597 B.n400 10.6151
R1395 B.n603 B.n400 10.6151
R1396 B.n604 B.n603 10.6151
R1397 B.n605 B.n604 10.6151
R1398 B.n605 B.n398 10.6151
R1399 B.n611 B.n398 10.6151
R1400 B.n612 B.n611 10.6151
R1401 B.n613 B.n612 10.6151
R1402 B.n613 B.n396 10.6151
R1403 B.n619 B.n396 10.6151
R1404 B.n620 B.n619 10.6151
R1405 B.n621 B.n620 10.6151
R1406 B.n621 B.n394 10.6151
R1407 B.n627 B.n394 10.6151
R1408 B.n628 B.n627 10.6151
R1409 B.n629 B.n628 10.6151
R1410 B.n629 B.n392 10.6151
R1411 B.n635 B.n392 10.6151
R1412 B.n636 B.n635 10.6151
R1413 B.n637 B.n636 10.6151
R1414 B.n637 B.n390 10.6151
R1415 B.n643 B.n390 10.6151
R1416 B.n644 B.n643 10.6151
R1417 B.n645 B.n644 10.6151
R1418 B.n645 B.n388 10.6151
R1419 B.n651 B.n388 10.6151
R1420 B.n652 B.n651 10.6151
R1421 B.n653 B.n652 10.6151
R1422 B.n653 B.n386 10.6151
R1423 B.n386 B.n385 10.6151
R1424 B.n660 B.n385 10.6151
R1425 B.n661 B.n660 10.6151
R1426 B.n667 B.n666 10.6151
R1427 B.n668 B.n667 10.6151
R1428 B.n668 B.n373 10.6151
R1429 B.n679 B.n373 10.6151
R1430 B.n680 B.n679 10.6151
R1431 B.n681 B.n680 10.6151
R1432 B.n681 B.n366 10.6151
R1433 B.n691 B.n366 10.6151
R1434 B.n692 B.n691 10.6151
R1435 B.n693 B.n692 10.6151
R1436 B.n693 B.n358 10.6151
R1437 B.n704 B.n358 10.6151
R1438 B.n705 B.n704 10.6151
R1439 B.n706 B.n705 10.6151
R1440 B.n706 B.n351 10.6151
R1441 B.n716 B.n351 10.6151
R1442 B.n717 B.n716 10.6151
R1443 B.n718 B.n717 10.6151
R1444 B.n718 B.n343 10.6151
R1445 B.n728 B.n343 10.6151
R1446 B.n729 B.n728 10.6151
R1447 B.n730 B.n729 10.6151
R1448 B.n730 B.n335 10.6151
R1449 B.n741 B.n335 10.6151
R1450 B.n742 B.n741 10.6151
R1451 B.n743 B.n742 10.6151
R1452 B.n743 B.n0 10.6151
R1453 B.n841 B.n1 10.6151
R1454 B.n841 B.n840 10.6151
R1455 B.n840 B.n839 10.6151
R1456 B.n839 B.n10 10.6151
R1457 B.n833 B.n10 10.6151
R1458 B.n833 B.n832 10.6151
R1459 B.n832 B.n831 10.6151
R1460 B.n831 B.n17 10.6151
R1461 B.n825 B.n17 10.6151
R1462 B.n825 B.n824 10.6151
R1463 B.n824 B.n823 10.6151
R1464 B.n823 B.n24 10.6151
R1465 B.n817 B.n24 10.6151
R1466 B.n817 B.n816 10.6151
R1467 B.n816 B.n815 10.6151
R1468 B.n815 B.n30 10.6151
R1469 B.n809 B.n30 10.6151
R1470 B.n809 B.n808 10.6151
R1471 B.n808 B.n807 10.6151
R1472 B.n807 B.n38 10.6151
R1473 B.n801 B.n38 10.6151
R1474 B.n801 B.n800 10.6151
R1475 B.n800 B.n799 10.6151
R1476 B.n799 B.n44 10.6151
R1477 B.n793 B.n44 10.6151
R1478 B.n793 B.n792 10.6151
R1479 B.n792 B.n791 10.6151
R1480 B.n212 B.n115 9.36635
R1481 B.n235 B.n112 9.36635
R1482 B.n540 B.n539 9.36635
R1483 B.n564 B.n563 9.36635
R1484 B.n708 B.t1 3.80203
R1485 B.t4 B.n345 3.80203
R1486 B.n739 B.t0 3.80203
R1487 B.n837 B.t3 3.80203
R1488 B.n828 B.t5 3.80203
R1489 B.n819 B.t2 3.80203
R1490 B.n847 B.n0 2.81026
R1491 B.n847 B.n1 2.81026
R1492 B.n215 B.n115 1.24928
R1493 B.n232 B.n112 1.24928
R1494 B.n539 B.n416 1.24928
R1495 B.n563 B.n562 1.24928
R1496 VP.n7 VP.t0 297.433
R1497 VP.n20 VP.t3 263.517
R1498 VP.n14 VP.t4 263.517
R1499 VP.n26 VP.t5 263.517
R1500 VP.n6 VP.t2 263.517
R1501 VP.n12 VP.t1 263.517
R1502 VP.n15 VP.n14 176.055
R1503 VP.n27 VP.n26 176.055
R1504 VP.n13 VP.n12 176.055
R1505 VP.n8 VP.n5 161.3
R1506 VP.n10 VP.n9 161.3
R1507 VP.n11 VP.n4 161.3
R1508 VP.n25 VP.n0 161.3
R1509 VP.n24 VP.n23 161.3
R1510 VP.n22 VP.n1 161.3
R1511 VP.n21 VP.n20 161.3
R1512 VP.n19 VP.n2 161.3
R1513 VP.n18 VP.n17 161.3
R1514 VP.n16 VP.n3 161.3
R1515 VP.n19 VP.n18 55.1086
R1516 VP.n24 VP.n1 55.1086
R1517 VP.n10 VP.n5 55.1086
R1518 VP.n15 VP.n13 46.0005
R1519 VP.n7 VP.n6 41.862
R1520 VP.n18 VP.n3 26.0455
R1521 VP.n25 VP.n24 26.0455
R1522 VP.n11 VP.n10 26.0455
R1523 VP.n20 VP.n19 24.5923
R1524 VP.n20 VP.n1 24.5923
R1525 VP.n6 VP.n5 24.5923
R1526 VP.n8 VP.n7 17.7677
R1527 VP.n14 VP.n3 9.83723
R1528 VP.n26 VP.n25 9.83723
R1529 VP.n12 VP.n11 9.83723
R1530 VP.n9 VP.n8 0.189894
R1531 VP.n9 VP.n4 0.189894
R1532 VP.n13 VP.n4 0.189894
R1533 VP.n16 VP.n15 0.189894
R1534 VP.n17 VP.n16 0.189894
R1535 VP.n17 VP.n2 0.189894
R1536 VP.n21 VP.n2 0.189894
R1537 VP.n22 VP.n21 0.189894
R1538 VP.n23 VP.n22 0.189894
R1539 VP.n23 VP.n0 0.189894
R1540 VP.n27 VP.n0 0.189894
R1541 VP VP.n27 0.0516364
R1542 VDD1 VDD1.t5 62.971
R1543 VDD1.n1 VDD1.t1 62.8572
R1544 VDD1.n1 VDD1.n0 60.8027
R1545 VDD1.n3 VDD1.n2 60.4918
R1546 VDD1.n3 VDD1.n1 42.7078
R1547 VDD1.n2 VDD1.t3 1.32226
R1548 VDD1.n2 VDD1.t4 1.32226
R1549 VDD1.n0 VDD1.t2 1.32226
R1550 VDD1.n0 VDD1.t0 1.32226
R1551 VDD1 VDD1.n3 0.30869
C0 VDD2 VDD1 0.959029f
C1 VN VDD2 7.04068f
C2 VDD2 VTAIL 9.59412f
C3 VP VDD1 7.24157f
C4 VN VP 6.28166f
C5 VP VTAIL 6.81241f
C6 VN VDD1 0.14942f
C7 VTAIL VDD1 9.554669f
C8 VN VTAIL 6.79788f
C9 VP VDD2 0.354907f
C10 VDD2 B 5.544674f
C11 VDD1 B 5.811231f
C12 VTAIL B 8.079161f
C13 VN B 9.729481f
C14 VP B 7.984685f
C15 VDD1.t5 B 2.99479f
C16 VDD1.t1 B 2.99408f
C17 VDD1.t2 B 0.259128f
C18 VDD1.t0 B 0.259128f
C19 VDD1.n0 B 2.34327f
C20 VDD1.n1 B 2.3238f
C21 VDD1.t3 B 0.259128f
C22 VDD1.t4 B 0.259128f
C23 VDD1.n2 B 2.34165f
C24 VDD1.n3 B 2.33882f
C25 VP.n0 B 0.033984f
C26 VP.t5 B 1.91103f
C27 VP.n1 B 0.05854f
C28 VP.n2 B 0.033984f
C29 VP.t3 B 1.91103f
C30 VP.n3 B 0.045984f
C31 VP.n4 B 0.033984f
C32 VP.t1 B 1.91103f
C33 VP.n5 B 0.05854f
C34 VP.t0 B 2.0027f
C35 VP.t2 B 1.91103f
C36 VP.n6 B 0.758402f
C37 VP.n7 B 0.755543f
C38 VP.n8 B 0.21162f
C39 VP.n9 B 0.033984f
C40 VP.n10 B 0.038629f
C41 VP.n11 B 0.045984f
C42 VP.n12 B 0.744347f
C43 VP.n13 B 1.63089f
C44 VP.t4 B 1.91103f
C45 VP.n14 B 0.744347f
C46 VP.n15 B 1.65752f
C47 VP.n16 B 0.033984f
C48 VP.n17 B 0.033984f
C49 VP.n18 B 0.038629f
C50 VP.n19 B 0.05854f
C51 VP.n20 B 0.714527f
C52 VP.n21 B 0.033984f
C53 VP.n22 B 0.033984f
C54 VP.n23 B 0.033984f
C55 VP.n24 B 0.038629f
C56 VP.n25 B 0.045984f
C57 VP.n26 B 0.744347f
C58 VP.n27 B 0.031983f
C59 VTAIL.t7 B 0.270234f
C60 VTAIL.t9 B 0.270234f
C61 VTAIL.n0 B 2.37234f
C62 VTAIL.n1 B 0.345725f
C63 VTAIL.t0 B 3.0262f
C64 VTAIL.n2 B 0.505439f
C65 VTAIL.t1 B 0.270234f
C66 VTAIL.t10 B 0.270234f
C67 VTAIL.n3 B 2.37234f
C68 VTAIL.n4 B 1.80945f
C69 VTAIL.t8 B 0.270234f
C70 VTAIL.t5 B 0.270234f
C71 VTAIL.n5 B 2.37235f
C72 VTAIL.n6 B 1.80944f
C73 VTAIL.t6 B 3.02621f
C74 VTAIL.n7 B 0.505435f
C75 VTAIL.t3 B 0.270234f
C76 VTAIL.t11 B 0.270234f
C77 VTAIL.n8 B 2.37235f
C78 VTAIL.n9 B 0.422292f
C79 VTAIL.t2 B 3.0262f
C80 VTAIL.n10 B 1.78479f
C81 VTAIL.t4 B 3.0262f
C82 VTAIL.n11 B 1.75356f
C83 VDD2.t3 B 2.97274f
C84 VDD2.t4 B 0.257281f
C85 VDD2.t2 B 0.257281f
C86 VDD2.n0 B 2.32657f
C87 VDD2.n1 B 2.22511f
C88 VDD2.t1 B 2.96743f
C89 VDD2.n2 B 2.34005f
C90 VDD2.t0 B 0.257281f
C91 VDD2.t5 B 0.257281f
C92 VDD2.n3 B 2.32654f
C93 VN.n0 B 0.03357f
C94 VN.t5 B 1.88776f
C95 VN.n1 B 0.057827f
C96 VN.t2 B 1.97831f
C97 VN.t0 B 1.88776f
C98 VN.n2 B 0.749167f
C99 VN.n3 B 0.746343f
C100 VN.n4 B 0.209043f
C101 VN.n5 B 0.03357f
C102 VN.n6 B 0.038158f
C103 VN.n7 B 0.045424f
C104 VN.n8 B 0.735283f
C105 VN.n9 B 0.031593f
C106 VN.n10 B 0.03357f
C107 VN.t1 B 1.88776f
C108 VN.n11 B 0.057827f
C109 VN.t3 B 1.97831f
C110 VN.t4 B 1.88776f
C111 VN.n12 B 0.749167f
C112 VN.n13 B 0.746343f
C113 VN.n14 B 0.209043f
C114 VN.n15 B 0.03357f
C115 VN.n16 B 0.038158f
C116 VN.n17 B 0.045424f
C117 VN.n18 B 0.735283f
C118 VN.n19 B 1.63295f
.ends

