* NGSPICE file created from diff_pair_sample_1239.ext - technology: sky130A

.subckt diff_pair_sample_1239 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=0.94215 pd=6.04 as=2.2269 ps=12.2 w=5.71 l=2.12
X1 VDD1.t3 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.94215 pd=6.04 as=2.2269 ps=12.2 w=5.71 l=2.12
X2 VDD1.t2 VP.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.94215 pd=6.04 as=2.2269 ps=12.2 w=5.71 l=2.12
X3 VTAIL.t7 VN.t1 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.2269 pd=12.2 as=0.94215 ps=6.04 w=5.71 l=2.12
X4 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=2.2269 pd=12.2 as=0 ps=0 w=5.71 l=2.12
X5 VTAIL.t6 VN.t2 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2269 pd=12.2 as=0.94215 ps=6.04 w=5.71 l=2.12
X6 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=2.2269 pd=12.2 as=0 ps=0 w=5.71 l=2.12
X7 VTAIL.t0 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.2269 pd=12.2 as=0.94215 ps=6.04 w=5.71 l=2.12
X8 VDD2.t0 VN.t3 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.94215 pd=6.04 as=2.2269 ps=12.2 w=5.71 l=2.12
X9 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.2269 pd=12.2 as=0 ps=0 w=5.71 l=2.12
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.2269 pd=12.2 as=0 ps=0 w=5.71 l=2.12
X11 VTAIL.t1 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2269 pd=12.2 as=0.94215 ps=6.04 w=5.71 l=2.12
R0 VN.n0 VN.t1 101.112
R1 VN.n1 VN.t3 101.112
R2 VN.n0 VN.t0 100.561
R3 VN.n1 VN.t2 100.561
R4 VN VN.n1 47.2374
R5 VN VN.n0 6.83209
R6 VTAIL.n5 VTAIL.t0 56.0164
R7 VTAIL.n4 VTAIL.t4 56.0164
R8 VTAIL.n3 VTAIL.t6 56.0164
R9 VTAIL.n7 VTAIL.t5 56.0162
R10 VTAIL.n0 VTAIL.t7 56.0162
R11 VTAIL.n1 VTAIL.t2 56.0162
R12 VTAIL.n2 VTAIL.t1 56.0162
R13 VTAIL.n6 VTAIL.t3 56.0162
R14 VTAIL.n7 VTAIL.n6 19.4014
R15 VTAIL.n3 VTAIL.n2 19.4014
R16 VTAIL.n4 VTAIL.n3 2.11257
R17 VTAIL.n6 VTAIL.n5 2.11257
R18 VTAIL.n2 VTAIL.n1 2.11257
R19 VTAIL VTAIL.n0 1.11472
R20 VTAIL VTAIL.n7 0.998345
R21 VTAIL.n5 VTAIL.n4 0.470328
R22 VTAIL.n1 VTAIL.n0 0.470328
R23 VDD2.n2 VDD2.n0 104.201
R24 VDD2.n2 VDD2.n1 69.2274
R25 VDD2.n1 VDD2.t1 3.4681
R26 VDD2.n1 VDD2.t0 3.4681
R27 VDD2.n0 VDD2.t2 3.4681
R28 VDD2.n0 VDD2.t3 3.4681
R29 VDD2 VDD2.n2 0.0586897
R30 B.n528 B.n527 585
R31 B.n199 B.n84 585
R32 B.n198 B.n197 585
R33 B.n196 B.n195 585
R34 B.n194 B.n193 585
R35 B.n192 B.n191 585
R36 B.n190 B.n189 585
R37 B.n188 B.n187 585
R38 B.n186 B.n185 585
R39 B.n184 B.n183 585
R40 B.n182 B.n181 585
R41 B.n180 B.n179 585
R42 B.n178 B.n177 585
R43 B.n176 B.n175 585
R44 B.n174 B.n173 585
R45 B.n172 B.n171 585
R46 B.n170 B.n169 585
R47 B.n168 B.n167 585
R48 B.n166 B.n165 585
R49 B.n164 B.n163 585
R50 B.n162 B.n161 585
R51 B.n160 B.n159 585
R52 B.n158 B.n157 585
R53 B.n155 B.n154 585
R54 B.n153 B.n152 585
R55 B.n151 B.n150 585
R56 B.n149 B.n148 585
R57 B.n147 B.n146 585
R58 B.n145 B.n144 585
R59 B.n143 B.n142 585
R60 B.n141 B.n140 585
R61 B.n139 B.n138 585
R62 B.n137 B.n136 585
R63 B.n134 B.n133 585
R64 B.n132 B.n131 585
R65 B.n130 B.n129 585
R66 B.n128 B.n127 585
R67 B.n126 B.n125 585
R68 B.n124 B.n123 585
R69 B.n122 B.n121 585
R70 B.n120 B.n119 585
R71 B.n118 B.n117 585
R72 B.n116 B.n115 585
R73 B.n114 B.n113 585
R74 B.n112 B.n111 585
R75 B.n110 B.n109 585
R76 B.n108 B.n107 585
R77 B.n106 B.n105 585
R78 B.n104 B.n103 585
R79 B.n102 B.n101 585
R80 B.n100 B.n99 585
R81 B.n98 B.n97 585
R82 B.n96 B.n95 585
R83 B.n94 B.n93 585
R84 B.n92 B.n91 585
R85 B.n90 B.n89 585
R86 B.n526 B.n56 585
R87 B.n531 B.n56 585
R88 B.n525 B.n55 585
R89 B.n532 B.n55 585
R90 B.n524 B.n523 585
R91 B.n523 B.n51 585
R92 B.n522 B.n50 585
R93 B.n538 B.n50 585
R94 B.n521 B.n49 585
R95 B.n539 B.n49 585
R96 B.n520 B.n48 585
R97 B.n540 B.n48 585
R98 B.n519 B.n518 585
R99 B.n518 B.n47 585
R100 B.n517 B.n43 585
R101 B.n546 B.n43 585
R102 B.n516 B.n42 585
R103 B.n547 B.n42 585
R104 B.n515 B.n41 585
R105 B.n548 B.n41 585
R106 B.n514 B.n513 585
R107 B.n513 B.n37 585
R108 B.n512 B.n36 585
R109 B.n554 B.n36 585
R110 B.n511 B.n35 585
R111 B.n555 B.n35 585
R112 B.n510 B.n34 585
R113 B.n556 B.n34 585
R114 B.n509 B.n508 585
R115 B.n508 B.n30 585
R116 B.n507 B.n29 585
R117 B.n562 B.n29 585
R118 B.n506 B.n28 585
R119 B.n563 B.n28 585
R120 B.n505 B.n27 585
R121 B.n564 B.n27 585
R122 B.n504 B.n503 585
R123 B.n503 B.n23 585
R124 B.n502 B.n22 585
R125 B.n570 B.n22 585
R126 B.n501 B.n21 585
R127 B.n571 B.n21 585
R128 B.n500 B.n20 585
R129 B.n572 B.n20 585
R130 B.n499 B.n498 585
R131 B.n498 B.n16 585
R132 B.n497 B.n15 585
R133 B.n578 B.n15 585
R134 B.n496 B.n14 585
R135 B.n579 B.n14 585
R136 B.n495 B.n13 585
R137 B.n580 B.n13 585
R138 B.n494 B.n493 585
R139 B.n493 B.n12 585
R140 B.n492 B.n491 585
R141 B.n492 B.n8 585
R142 B.n490 B.n7 585
R143 B.n587 B.n7 585
R144 B.n489 B.n6 585
R145 B.n588 B.n6 585
R146 B.n488 B.n5 585
R147 B.n589 B.n5 585
R148 B.n487 B.n486 585
R149 B.n486 B.n4 585
R150 B.n485 B.n200 585
R151 B.n485 B.n484 585
R152 B.n475 B.n201 585
R153 B.n202 B.n201 585
R154 B.n477 B.n476 585
R155 B.n478 B.n477 585
R156 B.n474 B.n206 585
R157 B.n210 B.n206 585
R158 B.n473 B.n472 585
R159 B.n472 B.n471 585
R160 B.n208 B.n207 585
R161 B.n209 B.n208 585
R162 B.n464 B.n463 585
R163 B.n465 B.n464 585
R164 B.n462 B.n215 585
R165 B.n215 B.n214 585
R166 B.n461 B.n460 585
R167 B.n460 B.n459 585
R168 B.n217 B.n216 585
R169 B.n218 B.n217 585
R170 B.n452 B.n451 585
R171 B.n453 B.n452 585
R172 B.n450 B.n223 585
R173 B.n223 B.n222 585
R174 B.n449 B.n448 585
R175 B.n448 B.n447 585
R176 B.n225 B.n224 585
R177 B.n226 B.n225 585
R178 B.n440 B.n439 585
R179 B.n441 B.n440 585
R180 B.n438 B.n231 585
R181 B.n231 B.n230 585
R182 B.n437 B.n436 585
R183 B.n436 B.n435 585
R184 B.n233 B.n232 585
R185 B.n234 B.n233 585
R186 B.n428 B.n427 585
R187 B.n429 B.n428 585
R188 B.n426 B.n239 585
R189 B.n239 B.n238 585
R190 B.n425 B.n424 585
R191 B.n424 B.n423 585
R192 B.n241 B.n240 585
R193 B.n416 B.n241 585
R194 B.n415 B.n414 585
R195 B.n417 B.n415 585
R196 B.n413 B.n246 585
R197 B.n246 B.n245 585
R198 B.n412 B.n411 585
R199 B.n411 B.n410 585
R200 B.n248 B.n247 585
R201 B.n249 B.n248 585
R202 B.n403 B.n402 585
R203 B.n404 B.n403 585
R204 B.n401 B.n254 585
R205 B.n254 B.n253 585
R206 B.n396 B.n395 585
R207 B.n394 B.n284 585
R208 B.n393 B.n283 585
R209 B.n398 B.n283 585
R210 B.n392 B.n391 585
R211 B.n390 B.n389 585
R212 B.n388 B.n387 585
R213 B.n386 B.n385 585
R214 B.n384 B.n383 585
R215 B.n382 B.n381 585
R216 B.n380 B.n379 585
R217 B.n378 B.n377 585
R218 B.n376 B.n375 585
R219 B.n374 B.n373 585
R220 B.n372 B.n371 585
R221 B.n370 B.n369 585
R222 B.n368 B.n367 585
R223 B.n366 B.n365 585
R224 B.n364 B.n363 585
R225 B.n362 B.n361 585
R226 B.n360 B.n359 585
R227 B.n358 B.n357 585
R228 B.n356 B.n355 585
R229 B.n354 B.n353 585
R230 B.n352 B.n351 585
R231 B.n350 B.n349 585
R232 B.n348 B.n347 585
R233 B.n346 B.n345 585
R234 B.n344 B.n343 585
R235 B.n342 B.n341 585
R236 B.n340 B.n339 585
R237 B.n338 B.n337 585
R238 B.n336 B.n335 585
R239 B.n334 B.n333 585
R240 B.n332 B.n331 585
R241 B.n330 B.n329 585
R242 B.n328 B.n327 585
R243 B.n326 B.n325 585
R244 B.n324 B.n323 585
R245 B.n322 B.n321 585
R246 B.n320 B.n319 585
R247 B.n318 B.n317 585
R248 B.n316 B.n315 585
R249 B.n314 B.n313 585
R250 B.n312 B.n311 585
R251 B.n310 B.n309 585
R252 B.n308 B.n307 585
R253 B.n306 B.n305 585
R254 B.n304 B.n303 585
R255 B.n302 B.n301 585
R256 B.n300 B.n299 585
R257 B.n298 B.n297 585
R258 B.n296 B.n295 585
R259 B.n294 B.n293 585
R260 B.n292 B.n291 585
R261 B.n256 B.n255 585
R262 B.n400 B.n399 585
R263 B.n399 B.n398 585
R264 B.n252 B.n251 585
R265 B.n253 B.n252 585
R266 B.n406 B.n405 585
R267 B.n405 B.n404 585
R268 B.n407 B.n250 585
R269 B.n250 B.n249 585
R270 B.n409 B.n408 585
R271 B.n410 B.n409 585
R272 B.n244 B.n243 585
R273 B.n245 B.n244 585
R274 B.n419 B.n418 585
R275 B.n418 B.n417 585
R276 B.n420 B.n242 585
R277 B.n416 B.n242 585
R278 B.n422 B.n421 585
R279 B.n423 B.n422 585
R280 B.n237 B.n236 585
R281 B.n238 B.n237 585
R282 B.n431 B.n430 585
R283 B.n430 B.n429 585
R284 B.n432 B.n235 585
R285 B.n235 B.n234 585
R286 B.n434 B.n433 585
R287 B.n435 B.n434 585
R288 B.n229 B.n228 585
R289 B.n230 B.n229 585
R290 B.n443 B.n442 585
R291 B.n442 B.n441 585
R292 B.n444 B.n227 585
R293 B.n227 B.n226 585
R294 B.n446 B.n445 585
R295 B.n447 B.n446 585
R296 B.n221 B.n220 585
R297 B.n222 B.n221 585
R298 B.n455 B.n454 585
R299 B.n454 B.n453 585
R300 B.n456 B.n219 585
R301 B.n219 B.n218 585
R302 B.n458 B.n457 585
R303 B.n459 B.n458 585
R304 B.n213 B.n212 585
R305 B.n214 B.n213 585
R306 B.n467 B.n466 585
R307 B.n466 B.n465 585
R308 B.n468 B.n211 585
R309 B.n211 B.n209 585
R310 B.n470 B.n469 585
R311 B.n471 B.n470 585
R312 B.n205 B.n204 585
R313 B.n210 B.n205 585
R314 B.n480 B.n479 585
R315 B.n479 B.n478 585
R316 B.n481 B.n203 585
R317 B.n203 B.n202 585
R318 B.n483 B.n482 585
R319 B.n484 B.n483 585
R320 B.n3 B.n0 585
R321 B.n4 B.n3 585
R322 B.n586 B.n1 585
R323 B.n587 B.n586 585
R324 B.n585 B.n584 585
R325 B.n585 B.n8 585
R326 B.n583 B.n9 585
R327 B.n12 B.n9 585
R328 B.n582 B.n581 585
R329 B.n581 B.n580 585
R330 B.n11 B.n10 585
R331 B.n579 B.n11 585
R332 B.n577 B.n576 585
R333 B.n578 B.n577 585
R334 B.n575 B.n17 585
R335 B.n17 B.n16 585
R336 B.n574 B.n573 585
R337 B.n573 B.n572 585
R338 B.n19 B.n18 585
R339 B.n571 B.n19 585
R340 B.n569 B.n568 585
R341 B.n570 B.n569 585
R342 B.n567 B.n24 585
R343 B.n24 B.n23 585
R344 B.n566 B.n565 585
R345 B.n565 B.n564 585
R346 B.n26 B.n25 585
R347 B.n563 B.n26 585
R348 B.n561 B.n560 585
R349 B.n562 B.n561 585
R350 B.n559 B.n31 585
R351 B.n31 B.n30 585
R352 B.n558 B.n557 585
R353 B.n557 B.n556 585
R354 B.n33 B.n32 585
R355 B.n555 B.n33 585
R356 B.n553 B.n552 585
R357 B.n554 B.n553 585
R358 B.n551 B.n38 585
R359 B.n38 B.n37 585
R360 B.n550 B.n549 585
R361 B.n549 B.n548 585
R362 B.n40 B.n39 585
R363 B.n547 B.n40 585
R364 B.n545 B.n544 585
R365 B.n546 B.n545 585
R366 B.n543 B.n44 585
R367 B.n47 B.n44 585
R368 B.n542 B.n541 585
R369 B.n541 B.n540 585
R370 B.n46 B.n45 585
R371 B.n539 B.n46 585
R372 B.n537 B.n536 585
R373 B.n538 B.n537 585
R374 B.n535 B.n52 585
R375 B.n52 B.n51 585
R376 B.n534 B.n533 585
R377 B.n533 B.n532 585
R378 B.n54 B.n53 585
R379 B.n531 B.n54 585
R380 B.n590 B.n589 585
R381 B.n588 B.n2 585
R382 B.n89 B.n54 521.33
R383 B.n528 B.n56 521.33
R384 B.n399 B.n254 521.33
R385 B.n396 B.n252 521.33
R386 B.n87 B.t12 272.098
R387 B.n85 B.t4 272.098
R388 B.n288 B.t15 272.098
R389 B.n285 B.t8 272.098
R390 B.n530 B.n529 256.663
R391 B.n530 B.n83 256.663
R392 B.n530 B.n82 256.663
R393 B.n530 B.n81 256.663
R394 B.n530 B.n80 256.663
R395 B.n530 B.n79 256.663
R396 B.n530 B.n78 256.663
R397 B.n530 B.n77 256.663
R398 B.n530 B.n76 256.663
R399 B.n530 B.n75 256.663
R400 B.n530 B.n74 256.663
R401 B.n530 B.n73 256.663
R402 B.n530 B.n72 256.663
R403 B.n530 B.n71 256.663
R404 B.n530 B.n70 256.663
R405 B.n530 B.n69 256.663
R406 B.n530 B.n68 256.663
R407 B.n530 B.n67 256.663
R408 B.n530 B.n66 256.663
R409 B.n530 B.n65 256.663
R410 B.n530 B.n64 256.663
R411 B.n530 B.n63 256.663
R412 B.n530 B.n62 256.663
R413 B.n530 B.n61 256.663
R414 B.n530 B.n60 256.663
R415 B.n530 B.n59 256.663
R416 B.n530 B.n58 256.663
R417 B.n530 B.n57 256.663
R418 B.n398 B.n397 256.663
R419 B.n398 B.n257 256.663
R420 B.n398 B.n258 256.663
R421 B.n398 B.n259 256.663
R422 B.n398 B.n260 256.663
R423 B.n398 B.n261 256.663
R424 B.n398 B.n262 256.663
R425 B.n398 B.n263 256.663
R426 B.n398 B.n264 256.663
R427 B.n398 B.n265 256.663
R428 B.n398 B.n266 256.663
R429 B.n398 B.n267 256.663
R430 B.n398 B.n268 256.663
R431 B.n398 B.n269 256.663
R432 B.n398 B.n270 256.663
R433 B.n398 B.n271 256.663
R434 B.n398 B.n272 256.663
R435 B.n398 B.n273 256.663
R436 B.n398 B.n274 256.663
R437 B.n398 B.n275 256.663
R438 B.n398 B.n276 256.663
R439 B.n398 B.n277 256.663
R440 B.n398 B.n278 256.663
R441 B.n398 B.n279 256.663
R442 B.n398 B.n280 256.663
R443 B.n398 B.n281 256.663
R444 B.n398 B.n282 256.663
R445 B.n592 B.n591 256.663
R446 B.n93 B.n92 163.367
R447 B.n97 B.n96 163.367
R448 B.n101 B.n100 163.367
R449 B.n105 B.n104 163.367
R450 B.n109 B.n108 163.367
R451 B.n113 B.n112 163.367
R452 B.n117 B.n116 163.367
R453 B.n121 B.n120 163.367
R454 B.n125 B.n124 163.367
R455 B.n129 B.n128 163.367
R456 B.n133 B.n132 163.367
R457 B.n138 B.n137 163.367
R458 B.n142 B.n141 163.367
R459 B.n146 B.n145 163.367
R460 B.n150 B.n149 163.367
R461 B.n154 B.n153 163.367
R462 B.n159 B.n158 163.367
R463 B.n163 B.n162 163.367
R464 B.n167 B.n166 163.367
R465 B.n171 B.n170 163.367
R466 B.n175 B.n174 163.367
R467 B.n179 B.n178 163.367
R468 B.n183 B.n182 163.367
R469 B.n187 B.n186 163.367
R470 B.n191 B.n190 163.367
R471 B.n195 B.n194 163.367
R472 B.n197 B.n84 163.367
R473 B.n403 B.n254 163.367
R474 B.n403 B.n248 163.367
R475 B.n411 B.n248 163.367
R476 B.n411 B.n246 163.367
R477 B.n415 B.n246 163.367
R478 B.n415 B.n241 163.367
R479 B.n424 B.n241 163.367
R480 B.n424 B.n239 163.367
R481 B.n428 B.n239 163.367
R482 B.n428 B.n233 163.367
R483 B.n436 B.n233 163.367
R484 B.n436 B.n231 163.367
R485 B.n440 B.n231 163.367
R486 B.n440 B.n225 163.367
R487 B.n448 B.n225 163.367
R488 B.n448 B.n223 163.367
R489 B.n452 B.n223 163.367
R490 B.n452 B.n217 163.367
R491 B.n460 B.n217 163.367
R492 B.n460 B.n215 163.367
R493 B.n464 B.n215 163.367
R494 B.n464 B.n208 163.367
R495 B.n472 B.n208 163.367
R496 B.n472 B.n206 163.367
R497 B.n477 B.n206 163.367
R498 B.n477 B.n201 163.367
R499 B.n485 B.n201 163.367
R500 B.n486 B.n485 163.367
R501 B.n486 B.n5 163.367
R502 B.n6 B.n5 163.367
R503 B.n7 B.n6 163.367
R504 B.n492 B.n7 163.367
R505 B.n493 B.n492 163.367
R506 B.n493 B.n13 163.367
R507 B.n14 B.n13 163.367
R508 B.n15 B.n14 163.367
R509 B.n498 B.n15 163.367
R510 B.n498 B.n20 163.367
R511 B.n21 B.n20 163.367
R512 B.n22 B.n21 163.367
R513 B.n503 B.n22 163.367
R514 B.n503 B.n27 163.367
R515 B.n28 B.n27 163.367
R516 B.n29 B.n28 163.367
R517 B.n508 B.n29 163.367
R518 B.n508 B.n34 163.367
R519 B.n35 B.n34 163.367
R520 B.n36 B.n35 163.367
R521 B.n513 B.n36 163.367
R522 B.n513 B.n41 163.367
R523 B.n42 B.n41 163.367
R524 B.n43 B.n42 163.367
R525 B.n518 B.n43 163.367
R526 B.n518 B.n48 163.367
R527 B.n49 B.n48 163.367
R528 B.n50 B.n49 163.367
R529 B.n523 B.n50 163.367
R530 B.n523 B.n55 163.367
R531 B.n56 B.n55 163.367
R532 B.n284 B.n283 163.367
R533 B.n391 B.n283 163.367
R534 B.n389 B.n388 163.367
R535 B.n385 B.n384 163.367
R536 B.n381 B.n380 163.367
R537 B.n377 B.n376 163.367
R538 B.n373 B.n372 163.367
R539 B.n369 B.n368 163.367
R540 B.n365 B.n364 163.367
R541 B.n361 B.n360 163.367
R542 B.n357 B.n356 163.367
R543 B.n353 B.n352 163.367
R544 B.n349 B.n348 163.367
R545 B.n345 B.n344 163.367
R546 B.n341 B.n340 163.367
R547 B.n337 B.n336 163.367
R548 B.n333 B.n332 163.367
R549 B.n329 B.n328 163.367
R550 B.n325 B.n324 163.367
R551 B.n321 B.n320 163.367
R552 B.n317 B.n316 163.367
R553 B.n313 B.n312 163.367
R554 B.n309 B.n308 163.367
R555 B.n305 B.n304 163.367
R556 B.n301 B.n300 163.367
R557 B.n297 B.n296 163.367
R558 B.n293 B.n292 163.367
R559 B.n399 B.n256 163.367
R560 B.n405 B.n252 163.367
R561 B.n405 B.n250 163.367
R562 B.n409 B.n250 163.367
R563 B.n409 B.n244 163.367
R564 B.n418 B.n244 163.367
R565 B.n418 B.n242 163.367
R566 B.n422 B.n242 163.367
R567 B.n422 B.n237 163.367
R568 B.n430 B.n237 163.367
R569 B.n430 B.n235 163.367
R570 B.n434 B.n235 163.367
R571 B.n434 B.n229 163.367
R572 B.n442 B.n229 163.367
R573 B.n442 B.n227 163.367
R574 B.n446 B.n227 163.367
R575 B.n446 B.n221 163.367
R576 B.n454 B.n221 163.367
R577 B.n454 B.n219 163.367
R578 B.n458 B.n219 163.367
R579 B.n458 B.n213 163.367
R580 B.n466 B.n213 163.367
R581 B.n466 B.n211 163.367
R582 B.n470 B.n211 163.367
R583 B.n470 B.n205 163.367
R584 B.n479 B.n205 163.367
R585 B.n479 B.n203 163.367
R586 B.n483 B.n203 163.367
R587 B.n483 B.n3 163.367
R588 B.n590 B.n3 163.367
R589 B.n586 B.n2 163.367
R590 B.n586 B.n585 163.367
R591 B.n585 B.n9 163.367
R592 B.n581 B.n9 163.367
R593 B.n581 B.n11 163.367
R594 B.n577 B.n11 163.367
R595 B.n577 B.n17 163.367
R596 B.n573 B.n17 163.367
R597 B.n573 B.n19 163.367
R598 B.n569 B.n19 163.367
R599 B.n569 B.n24 163.367
R600 B.n565 B.n24 163.367
R601 B.n565 B.n26 163.367
R602 B.n561 B.n26 163.367
R603 B.n561 B.n31 163.367
R604 B.n557 B.n31 163.367
R605 B.n557 B.n33 163.367
R606 B.n553 B.n33 163.367
R607 B.n553 B.n38 163.367
R608 B.n549 B.n38 163.367
R609 B.n549 B.n40 163.367
R610 B.n545 B.n40 163.367
R611 B.n545 B.n44 163.367
R612 B.n541 B.n44 163.367
R613 B.n541 B.n46 163.367
R614 B.n537 B.n46 163.367
R615 B.n537 B.n52 163.367
R616 B.n533 B.n52 163.367
R617 B.n533 B.n54 163.367
R618 B.n398 B.n253 139.19
R619 B.n531 B.n530 139.19
R620 B.n85 B.t6 122.383
R621 B.n288 B.t17 122.383
R622 B.n87 B.t13 122.377
R623 B.n285 B.t11 122.377
R624 B.n86 B.t7 74.8683
R625 B.n289 B.t16 74.8683
R626 B.n88 B.t14 74.8625
R627 B.n286 B.t10 74.8625
R628 B.n89 B.n57 71.676
R629 B.n93 B.n58 71.676
R630 B.n97 B.n59 71.676
R631 B.n101 B.n60 71.676
R632 B.n105 B.n61 71.676
R633 B.n109 B.n62 71.676
R634 B.n113 B.n63 71.676
R635 B.n117 B.n64 71.676
R636 B.n121 B.n65 71.676
R637 B.n125 B.n66 71.676
R638 B.n129 B.n67 71.676
R639 B.n133 B.n68 71.676
R640 B.n138 B.n69 71.676
R641 B.n142 B.n70 71.676
R642 B.n146 B.n71 71.676
R643 B.n150 B.n72 71.676
R644 B.n154 B.n73 71.676
R645 B.n159 B.n74 71.676
R646 B.n163 B.n75 71.676
R647 B.n167 B.n76 71.676
R648 B.n171 B.n77 71.676
R649 B.n175 B.n78 71.676
R650 B.n179 B.n79 71.676
R651 B.n183 B.n80 71.676
R652 B.n187 B.n81 71.676
R653 B.n191 B.n82 71.676
R654 B.n195 B.n83 71.676
R655 B.n529 B.n84 71.676
R656 B.n529 B.n528 71.676
R657 B.n197 B.n83 71.676
R658 B.n194 B.n82 71.676
R659 B.n190 B.n81 71.676
R660 B.n186 B.n80 71.676
R661 B.n182 B.n79 71.676
R662 B.n178 B.n78 71.676
R663 B.n174 B.n77 71.676
R664 B.n170 B.n76 71.676
R665 B.n166 B.n75 71.676
R666 B.n162 B.n74 71.676
R667 B.n158 B.n73 71.676
R668 B.n153 B.n72 71.676
R669 B.n149 B.n71 71.676
R670 B.n145 B.n70 71.676
R671 B.n141 B.n69 71.676
R672 B.n137 B.n68 71.676
R673 B.n132 B.n67 71.676
R674 B.n128 B.n66 71.676
R675 B.n124 B.n65 71.676
R676 B.n120 B.n64 71.676
R677 B.n116 B.n63 71.676
R678 B.n112 B.n62 71.676
R679 B.n108 B.n61 71.676
R680 B.n104 B.n60 71.676
R681 B.n100 B.n59 71.676
R682 B.n96 B.n58 71.676
R683 B.n92 B.n57 71.676
R684 B.n397 B.n396 71.676
R685 B.n391 B.n257 71.676
R686 B.n388 B.n258 71.676
R687 B.n384 B.n259 71.676
R688 B.n380 B.n260 71.676
R689 B.n376 B.n261 71.676
R690 B.n372 B.n262 71.676
R691 B.n368 B.n263 71.676
R692 B.n364 B.n264 71.676
R693 B.n360 B.n265 71.676
R694 B.n356 B.n266 71.676
R695 B.n352 B.n267 71.676
R696 B.n348 B.n268 71.676
R697 B.n344 B.n269 71.676
R698 B.n340 B.n270 71.676
R699 B.n336 B.n271 71.676
R700 B.n332 B.n272 71.676
R701 B.n328 B.n273 71.676
R702 B.n324 B.n274 71.676
R703 B.n320 B.n275 71.676
R704 B.n316 B.n276 71.676
R705 B.n312 B.n277 71.676
R706 B.n308 B.n278 71.676
R707 B.n304 B.n279 71.676
R708 B.n300 B.n280 71.676
R709 B.n296 B.n281 71.676
R710 B.n292 B.n282 71.676
R711 B.n397 B.n284 71.676
R712 B.n389 B.n257 71.676
R713 B.n385 B.n258 71.676
R714 B.n381 B.n259 71.676
R715 B.n377 B.n260 71.676
R716 B.n373 B.n261 71.676
R717 B.n369 B.n262 71.676
R718 B.n365 B.n263 71.676
R719 B.n361 B.n264 71.676
R720 B.n357 B.n265 71.676
R721 B.n353 B.n266 71.676
R722 B.n349 B.n267 71.676
R723 B.n345 B.n268 71.676
R724 B.n341 B.n269 71.676
R725 B.n337 B.n270 71.676
R726 B.n333 B.n271 71.676
R727 B.n329 B.n272 71.676
R728 B.n325 B.n273 71.676
R729 B.n321 B.n274 71.676
R730 B.n317 B.n275 71.676
R731 B.n313 B.n276 71.676
R732 B.n309 B.n277 71.676
R733 B.n305 B.n278 71.676
R734 B.n301 B.n279 71.676
R735 B.n297 B.n280 71.676
R736 B.n293 B.n281 71.676
R737 B.n282 B.n256 71.676
R738 B.n591 B.n590 71.676
R739 B.n591 B.n2 71.676
R740 B.n404 B.n253 68.0933
R741 B.n404 B.n249 68.0933
R742 B.n410 B.n249 68.0933
R743 B.n410 B.n245 68.0933
R744 B.n417 B.n245 68.0933
R745 B.n417 B.n416 68.0933
R746 B.n423 B.n238 68.0933
R747 B.n429 B.n238 68.0933
R748 B.n429 B.n234 68.0933
R749 B.n435 B.n234 68.0933
R750 B.n435 B.n230 68.0933
R751 B.n441 B.n230 68.0933
R752 B.n441 B.n226 68.0933
R753 B.n447 B.n226 68.0933
R754 B.n447 B.n222 68.0933
R755 B.n453 B.n222 68.0933
R756 B.n459 B.n218 68.0933
R757 B.n459 B.n214 68.0933
R758 B.n465 B.n214 68.0933
R759 B.n465 B.n209 68.0933
R760 B.n471 B.n209 68.0933
R761 B.n471 B.n210 68.0933
R762 B.n478 B.n202 68.0933
R763 B.n484 B.n202 68.0933
R764 B.n484 B.n4 68.0933
R765 B.n589 B.n4 68.0933
R766 B.n589 B.n588 68.0933
R767 B.n588 B.n587 68.0933
R768 B.n587 B.n8 68.0933
R769 B.n12 B.n8 68.0933
R770 B.n580 B.n12 68.0933
R771 B.n579 B.n578 68.0933
R772 B.n578 B.n16 68.0933
R773 B.n572 B.n16 68.0933
R774 B.n572 B.n571 68.0933
R775 B.n571 B.n570 68.0933
R776 B.n570 B.n23 68.0933
R777 B.n564 B.n563 68.0933
R778 B.n563 B.n562 68.0933
R779 B.n562 B.n30 68.0933
R780 B.n556 B.n30 68.0933
R781 B.n556 B.n555 68.0933
R782 B.n555 B.n554 68.0933
R783 B.n554 B.n37 68.0933
R784 B.n548 B.n37 68.0933
R785 B.n548 B.n547 68.0933
R786 B.n547 B.n546 68.0933
R787 B.n540 B.n47 68.0933
R788 B.n540 B.n539 68.0933
R789 B.n539 B.n538 68.0933
R790 B.n538 B.n51 68.0933
R791 B.n532 B.n51 68.0933
R792 B.n532 B.n531 68.0933
R793 B.t1 B.n218 62.0852
R794 B.t3 B.n23 62.0852
R795 B.n135 B.n88 59.5399
R796 B.n156 B.n86 59.5399
R797 B.n290 B.n289 59.5399
R798 B.n287 B.n286 59.5399
R799 B.n478 B.t2 48.066
R800 B.n580 B.t0 48.066
R801 B.n88 B.n87 47.5157
R802 B.n86 B.n85 47.5157
R803 B.n289 B.n288 47.5157
R804 B.n286 B.n285 47.5157
R805 B.n416 B.t9 46.0633
R806 B.n47 B.t5 46.0633
R807 B.n395 B.n251 33.8737
R808 B.n401 B.n400 33.8737
R809 B.n527 B.n526 33.8737
R810 B.n90 B.n53 33.8737
R811 B.n423 B.t9 22.0305
R812 B.n546 B.t5 22.0305
R813 B.n210 B.t2 20.0278
R814 B.t0 B.n579 20.0278
R815 B B.n592 18.0485
R816 B.n406 B.n251 10.6151
R817 B.n407 B.n406 10.6151
R818 B.n408 B.n407 10.6151
R819 B.n408 B.n243 10.6151
R820 B.n419 B.n243 10.6151
R821 B.n420 B.n419 10.6151
R822 B.n421 B.n420 10.6151
R823 B.n421 B.n236 10.6151
R824 B.n431 B.n236 10.6151
R825 B.n432 B.n431 10.6151
R826 B.n433 B.n432 10.6151
R827 B.n433 B.n228 10.6151
R828 B.n443 B.n228 10.6151
R829 B.n444 B.n443 10.6151
R830 B.n445 B.n444 10.6151
R831 B.n445 B.n220 10.6151
R832 B.n455 B.n220 10.6151
R833 B.n456 B.n455 10.6151
R834 B.n457 B.n456 10.6151
R835 B.n457 B.n212 10.6151
R836 B.n467 B.n212 10.6151
R837 B.n468 B.n467 10.6151
R838 B.n469 B.n468 10.6151
R839 B.n469 B.n204 10.6151
R840 B.n480 B.n204 10.6151
R841 B.n481 B.n480 10.6151
R842 B.n482 B.n481 10.6151
R843 B.n482 B.n0 10.6151
R844 B.n395 B.n394 10.6151
R845 B.n394 B.n393 10.6151
R846 B.n393 B.n392 10.6151
R847 B.n392 B.n390 10.6151
R848 B.n390 B.n387 10.6151
R849 B.n387 B.n386 10.6151
R850 B.n386 B.n383 10.6151
R851 B.n383 B.n382 10.6151
R852 B.n382 B.n379 10.6151
R853 B.n379 B.n378 10.6151
R854 B.n378 B.n375 10.6151
R855 B.n375 B.n374 10.6151
R856 B.n374 B.n371 10.6151
R857 B.n371 B.n370 10.6151
R858 B.n370 B.n367 10.6151
R859 B.n367 B.n366 10.6151
R860 B.n366 B.n363 10.6151
R861 B.n363 B.n362 10.6151
R862 B.n362 B.n359 10.6151
R863 B.n359 B.n358 10.6151
R864 B.n358 B.n355 10.6151
R865 B.n355 B.n354 10.6151
R866 B.n351 B.n350 10.6151
R867 B.n350 B.n347 10.6151
R868 B.n347 B.n346 10.6151
R869 B.n346 B.n343 10.6151
R870 B.n343 B.n342 10.6151
R871 B.n342 B.n339 10.6151
R872 B.n339 B.n338 10.6151
R873 B.n338 B.n335 10.6151
R874 B.n335 B.n334 10.6151
R875 B.n331 B.n330 10.6151
R876 B.n330 B.n327 10.6151
R877 B.n327 B.n326 10.6151
R878 B.n326 B.n323 10.6151
R879 B.n323 B.n322 10.6151
R880 B.n322 B.n319 10.6151
R881 B.n319 B.n318 10.6151
R882 B.n318 B.n315 10.6151
R883 B.n315 B.n314 10.6151
R884 B.n314 B.n311 10.6151
R885 B.n311 B.n310 10.6151
R886 B.n310 B.n307 10.6151
R887 B.n307 B.n306 10.6151
R888 B.n306 B.n303 10.6151
R889 B.n303 B.n302 10.6151
R890 B.n302 B.n299 10.6151
R891 B.n299 B.n298 10.6151
R892 B.n298 B.n295 10.6151
R893 B.n295 B.n294 10.6151
R894 B.n294 B.n291 10.6151
R895 B.n291 B.n255 10.6151
R896 B.n400 B.n255 10.6151
R897 B.n402 B.n401 10.6151
R898 B.n402 B.n247 10.6151
R899 B.n412 B.n247 10.6151
R900 B.n413 B.n412 10.6151
R901 B.n414 B.n413 10.6151
R902 B.n414 B.n240 10.6151
R903 B.n425 B.n240 10.6151
R904 B.n426 B.n425 10.6151
R905 B.n427 B.n426 10.6151
R906 B.n427 B.n232 10.6151
R907 B.n437 B.n232 10.6151
R908 B.n438 B.n437 10.6151
R909 B.n439 B.n438 10.6151
R910 B.n439 B.n224 10.6151
R911 B.n449 B.n224 10.6151
R912 B.n450 B.n449 10.6151
R913 B.n451 B.n450 10.6151
R914 B.n451 B.n216 10.6151
R915 B.n461 B.n216 10.6151
R916 B.n462 B.n461 10.6151
R917 B.n463 B.n462 10.6151
R918 B.n463 B.n207 10.6151
R919 B.n473 B.n207 10.6151
R920 B.n474 B.n473 10.6151
R921 B.n476 B.n474 10.6151
R922 B.n476 B.n475 10.6151
R923 B.n475 B.n200 10.6151
R924 B.n487 B.n200 10.6151
R925 B.n488 B.n487 10.6151
R926 B.n489 B.n488 10.6151
R927 B.n490 B.n489 10.6151
R928 B.n491 B.n490 10.6151
R929 B.n494 B.n491 10.6151
R930 B.n495 B.n494 10.6151
R931 B.n496 B.n495 10.6151
R932 B.n497 B.n496 10.6151
R933 B.n499 B.n497 10.6151
R934 B.n500 B.n499 10.6151
R935 B.n501 B.n500 10.6151
R936 B.n502 B.n501 10.6151
R937 B.n504 B.n502 10.6151
R938 B.n505 B.n504 10.6151
R939 B.n506 B.n505 10.6151
R940 B.n507 B.n506 10.6151
R941 B.n509 B.n507 10.6151
R942 B.n510 B.n509 10.6151
R943 B.n511 B.n510 10.6151
R944 B.n512 B.n511 10.6151
R945 B.n514 B.n512 10.6151
R946 B.n515 B.n514 10.6151
R947 B.n516 B.n515 10.6151
R948 B.n517 B.n516 10.6151
R949 B.n519 B.n517 10.6151
R950 B.n520 B.n519 10.6151
R951 B.n521 B.n520 10.6151
R952 B.n522 B.n521 10.6151
R953 B.n524 B.n522 10.6151
R954 B.n525 B.n524 10.6151
R955 B.n526 B.n525 10.6151
R956 B.n584 B.n1 10.6151
R957 B.n584 B.n583 10.6151
R958 B.n583 B.n582 10.6151
R959 B.n582 B.n10 10.6151
R960 B.n576 B.n10 10.6151
R961 B.n576 B.n575 10.6151
R962 B.n575 B.n574 10.6151
R963 B.n574 B.n18 10.6151
R964 B.n568 B.n18 10.6151
R965 B.n568 B.n567 10.6151
R966 B.n567 B.n566 10.6151
R967 B.n566 B.n25 10.6151
R968 B.n560 B.n25 10.6151
R969 B.n560 B.n559 10.6151
R970 B.n559 B.n558 10.6151
R971 B.n558 B.n32 10.6151
R972 B.n552 B.n32 10.6151
R973 B.n552 B.n551 10.6151
R974 B.n551 B.n550 10.6151
R975 B.n550 B.n39 10.6151
R976 B.n544 B.n39 10.6151
R977 B.n544 B.n543 10.6151
R978 B.n543 B.n542 10.6151
R979 B.n542 B.n45 10.6151
R980 B.n536 B.n45 10.6151
R981 B.n536 B.n535 10.6151
R982 B.n535 B.n534 10.6151
R983 B.n534 B.n53 10.6151
R984 B.n91 B.n90 10.6151
R985 B.n94 B.n91 10.6151
R986 B.n95 B.n94 10.6151
R987 B.n98 B.n95 10.6151
R988 B.n99 B.n98 10.6151
R989 B.n102 B.n99 10.6151
R990 B.n103 B.n102 10.6151
R991 B.n106 B.n103 10.6151
R992 B.n107 B.n106 10.6151
R993 B.n110 B.n107 10.6151
R994 B.n111 B.n110 10.6151
R995 B.n114 B.n111 10.6151
R996 B.n115 B.n114 10.6151
R997 B.n118 B.n115 10.6151
R998 B.n119 B.n118 10.6151
R999 B.n122 B.n119 10.6151
R1000 B.n123 B.n122 10.6151
R1001 B.n126 B.n123 10.6151
R1002 B.n127 B.n126 10.6151
R1003 B.n130 B.n127 10.6151
R1004 B.n131 B.n130 10.6151
R1005 B.n134 B.n131 10.6151
R1006 B.n139 B.n136 10.6151
R1007 B.n140 B.n139 10.6151
R1008 B.n143 B.n140 10.6151
R1009 B.n144 B.n143 10.6151
R1010 B.n147 B.n144 10.6151
R1011 B.n148 B.n147 10.6151
R1012 B.n151 B.n148 10.6151
R1013 B.n152 B.n151 10.6151
R1014 B.n155 B.n152 10.6151
R1015 B.n160 B.n157 10.6151
R1016 B.n161 B.n160 10.6151
R1017 B.n164 B.n161 10.6151
R1018 B.n165 B.n164 10.6151
R1019 B.n168 B.n165 10.6151
R1020 B.n169 B.n168 10.6151
R1021 B.n172 B.n169 10.6151
R1022 B.n173 B.n172 10.6151
R1023 B.n176 B.n173 10.6151
R1024 B.n177 B.n176 10.6151
R1025 B.n180 B.n177 10.6151
R1026 B.n181 B.n180 10.6151
R1027 B.n184 B.n181 10.6151
R1028 B.n185 B.n184 10.6151
R1029 B.n188 B.n185 10.6151
R1030 B.n189 B.n188 10.6151
R1031 B.n192 B.n189 10.6151
R1032 B.n193 B.n192 10.6151
R1033 B.n196 B.n193 10.6151
R1034 B.n198 B.n196 10.6151
R1035 B.n199 B.n198 10.6151
R1036 B.n527 B.n199 10.6151
R1037 B.n354 B.n287 9.36635
R1038 B.n331 B.n290 9.36635
R1039 B.n135 B.n134 9.36635
R1040 B.n157 B.n156 9.36635
R1041 B.n592 B.n0 8.11757
R1042 B.n592 B.n1 8.11757
R1043 B.n453 B.t1 6.00869
R1044 B.n564 B.t3 6.00869
R1045 B.n351 B.n287 1.24928
R1046 B.n334 B.n290 1.24928
R1047 B.n136 B.n135 1.24928
R1048 B.n156 B.n155 1.24928
R1049 VP.n10 VP.n0 161.3
R1050 VP.n9 VP.n8 161.3
R1051 VP.n7 VP.n1 161.3
R1052 VP.n6 VP.n5 161.3
R1053 VP.n2 VP.t2 101.112
R1054 VP.n2 VP.t1 100.561
R1055 VP.n4 VP.n3 87.5128
R1056 VP.n12 VP.n11 87.5128
R1057 VP.n4 VP.t3 64.9114
R1058 VP.n11 VP.t0 64.9114
R1059 VP.n9 VP.n1 56.5193
R1060 VP.n3 VP.n2 46.9585
R1061 VP.n5 VP.n1 24.4675
R1062 VP.n10 VP.n9 24.4675
R1063 VP.n5 VP.n4 23.2442
R1064 VP.n11 VP.n10 23.2442
R1065 VP.n6 VP.n3 0.278367
R1066 VP.n12 VP.n0 0.278367
R1067 VP.n7 VP.n6 0.189894
R1068 VP.n8 VP.n7 0.189894
R1069 VP.n8 VP.n0 0.189894
R1070 VP VP.n12 0.153454
R1071 VDD1 VDD1.n1 104.725
R1072 VDD1 VDD1.n0 69.2856
R1073 VDD1.n0 VDD1.t1 3.4681
R1074 VDD1.n0 VDD1.t2 3.4681
R1075 VDD1.n1 VDD1.t0 3.4681
R1076 VDD1.n1 VDD1.t3 3.4681
C0 VDD2 VN 2.33356f
C1 VDD1 VTAIL 3.74937f
C2 VDD2 VP 0.36389f
C3 VDD1 VN 0.148694f
C4 VDD1 VP 2.54814f
C5 VN VTAIL 2.54903f
C6 VDD1 VDD2 0.913864f
C7 VTAIL VP 2.56314f
C8 VDD2 VTAIL 3.80036f
C9 VN VP 4.6776f
C10 VDD2 B 3.00275f
C11 VDD1 B 6.29714f
C12 VTAIL B 5.829346f
C13 VN B 9.189349f
C14 VP B 7.377882f
C15 VDD1.t1 B 0.122643f
C16 VDD1.t2 B 0.122643f
C17 VDD1.n0 B 1.01731f
C18 VDD1.t0 B 0.122643f
C19 VDD1.t3 B 0.122643f
C20 VDD1.n1 B 1.45606f
C21 VP.n0 B 0.043465f
C22 VP.t0 B 1.05313f
C23 VP.n1 B 0.048127f
C24 VP.t1 B 1.26142f
C25 VP.t2 B 1.26454f
C26 VP.n2 B 2.14321f
C27 VP.n3 B 1.53926f
C28 VP.t3 B 1.05313f
C29 VP.n4 B 0.51752f
C30 VP.n5 B 0.059926f
C31 VP.n6 B 0.043465f
C32 VP.n7 B 0.032968f
C33 VP.n8 B 0.032968f
C34 VP.n9 B 0.048127f
C35 VP.n10 B 0.059926f
C36 VP.n11 B 0.51752f
C37 VP.n12 B 0.036863f
C38 VDD2.t2 B 0.122651f
C39 VDD2.t3 B 0.122651f
C40 VDD2.n0 B 1.43337f
C41 VDD2.t1 B 0.122651f
C42 VDD2.t0 B 0.122651f
C43 VDD2.n1 B 1.01702f
C44 VDD2.n2 B 2.96816f
C45 VTAIL.t7 B 0.85505f
C46 VTAIL.n0 B 0.325141f
C47 VTAIL.t2 B 0.85505f
C48 VTAIL.n1 B 0.386812f
C49 VTAIL.t1 B 0.85505f
C50 VTAIL.n2 B 1.05309f
C51 VTAIL.t6 B 0.855054f
C52 VTAIL.n3 B 1.05308f
C53 VTAIL.t4 B 0.855054f
C54 VTAIL.n4 B 0.386809f
C55 VTAIL.t0 B 0.855054f
C56 VTAIL.n5 B 0.386809f
C57 VTAIL.t3 B 0.85505f
C58 VTAIL.n6 B 1.05309f
C59 VTAIL.t5 B 0.85505f
C60 VTAIL.n7 B 0.984222f
C61 VN.t1 B 1.22006f
C62 VN.t0 B 1.21705f
C63 VN.n0 B 0.815935f
C64 VN.t3 B 1.22006f
C65 VN.t2 B 1.21705f
C66 VN.n1 B 2.08429f
.ends

