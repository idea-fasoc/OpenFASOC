* NGSPICE file created from diff_pair_sample_0583.ext - technology: sky130A

.subckt diff_pair_sample_0583 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t15 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=2.0046 pd=11.06 as=0.8481 ps=5.47 w=5.14 l=0.63
X1 VDD1.t9 VP.t0 VTAIL.t3 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=0.8481 pd=5.47 as=0.8481 ps=5.47 w=5.14 l=0.63
X2 B.t11 B.t9 B.t10 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=2.0046 pd=11.06 as=0 ps=0 w=5.14 l=0.63
X3 B.t8 B.t6 B.t7 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=2.0046 pd=11.06 as=0 ps=0 w=5.14 l=0.63
X4 VDD1.t8 VP.t1 VTAIL.t8 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=0.8481 pd=5.47 as=2.0046 ps=11.06 w=5.14 l=0.63
X5 VTAIL.t10 VN.t1 VDD2.t8 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=0.8481 pd=5.47 as=0.8481 ps=5.47 w=5.14 l=0.63
X6 VDD2.t7 VN.t2 VTAIL.t13 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=0.8481 pd=5.47 as=2.0046 ps=11.06 w=5.14 l=0.63
X7 VTAIL.t18 VN.t3 VDD2.t6 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=0.8481 pd=5.47 as=0.8481 ps=5.47 w=5.14 l=0.63
X8 VDD2.t5 VN.t4 VTAIL.t16 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=0.8481 pd=5.47 as=0.8481 ps=5.47 w=5.14 l=0.63
X9 VDD2.t4 VN.t5 VTAIL.t19 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=2.0046 pd=11.06 as=0.8481 ps=5.47 w=5.14 l=0.63
X10 VTAIL.t17 VN.t6 VDD2.t3 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=0.8481 pd=5.47 as=0.8481 ps=5.47 w=5.14 l=0.63
X11 VTAIL.t12 VN.t7 VDD2.t2 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=0.8481 pd=5.47 as=0.8481 ps=5.47 w=5.14 l=0.63
X12 VTAIL.t5 VP.t2 VDD1.t7 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=0.8481 pd=5.47 as=0.8481 ps=5.47 w=5.14 l=0.63
X13 VDD1.t6 VP.t3 VTAIL.t6 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=0.8481 pd=5.47 as=2.0046 ps=11.06 w=5.14 l=0.63
X14 VTAIL.t4 VP.t4 VDD1.t5 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=0.8481 pd=5.47 as=0.8481 ps=5.47 w=5.14 l=0.63
X15 VDD1.t4 VP.t5 VTAIL.t9 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=0.8481 pd=5.47 as=0.8481 ps=5.47 w=5.14 l=0.63
X16 VDD1.t3 VP.t6 VTAIL.t7 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=2.0046 pd=11.06 as=0.8481 ps=5.47 w=5.14 l=0.63
X17 VTAIL.t0 VP.t7 VDD1.t2 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=0.8481 pd=5.47 as=0.8481 ps=5.47 w=5.14 l=0.63
X18 VTAIL.t1 VP.t8 VDD1.t1 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=0.8481 pd=5.47 as=0.8481 ps=5.47 w=5.14 l=0.63
X19 VDD2.t1 VN.t8 VTAIL.t14 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=0.8481 pd=5.47 as=2.0046 ps=11.06 w=5.14 l=0.63
X20 VDD2.t0 VN.t9 VTAIL.t11 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=0.8481 pd=5.47 as=0.8481 ps=5.47 w=5.14 l=0.63
X21 VDD1.t0 VP.t9 VTAIL.t2 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=2.0046 pd=11.06 as=0.8481 ps=5.47 w=5.14 l=0.63
X22 B.t5 B.t3 B.t4 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=2.0046 pd=11.06 as=0 ps=0 w=5.14 l=0.63
X23 B.t2 B.t0 B.t1 w_n2122_n1996# sky130_fd_pr__pfet_01v8 ad=2.0046 pd=11.06 as=0 ps=0 w=5.14 l=0.63
R0 VN.n2 VN.t0 285.8
R1 VN.n10 VN.t2 285.8
R2 VN.n1 VN.t7 258.979
R3 VN.n4 VN.t9 258.979
R4 VN.n5 VN.t1 258.979
R5 VN.n6 VN.t8 258.979
R6 VN.n9 VN.t3 258.979
R7 VN.n12 VN.t4 258.979
R8 VN.n13 VN.t6 258.979
R9 VN.n14 VN.t5 258.979
R10 VN.n7 VN.n6 161.3
R11 VN.n15 VN.n14 161.3
R12 VN.n13 VN.n8 80.6037
R13 VN.n12 VN.n11 80.6037
R14 VN.n5 VN.n0 80.6037
R15 VN.n4 VN.n3 80.6037
R16 VN.n4 VN.n1 48.2005
R17 VN.n5 VN.n4 48.2005
R18 VN.n6 VN.n5 48.2005
R19 VN.n12 VN.n9 48.2005
R20 VN.n13 VN.n12 48.2005
R21 VN.n14 VN.n13 48.2005
R22 VN.n11 VN.n10 45.2318
R23 VN.n3 VN.n2 45.2318
R24 VN VN.n15 37.6539
R25 VN.n10 VN.n9 13.3799
R26 VN.n2 VN.n1 13.3799
R27 VN.n11 VN.n8 0.380177
R28 VN.n3 VN.n0 0.380177
R29 VN.n15 VN.n8 0.285035
R30 VN.n7 VN.n0 0.285035
R31 VN VN.n7 0.0516364
R32 VTAIL.n116 VTAIL.n115 756.745
R33 VTAIL.n26 VTAIL.n25 756.745
R34 VTAIL.n90 VTAIL.n89 756.745
R35 VTAIL.n60 VTAIL.n59 756.745
R36 VTAIL.n101 VTAIL.n100 585
R37 VTAIL.n98 VTAIL.n97 585
R38 VTAIL.n107 VTAIL.n106 585
R39 VTAIL.n109 VTAIL.n108 585
R40 VTAIL.n94 VTAIL.n93 585
R41 VTAIL.n115 VTAIL.n114 585
R42 VTAIL.n11 VTAIL.n10 585
R43 VTAIL.n8 VTAIL.n7 585
R44 VTAIL.n17 VTAIL.n16 585
R45 VTAIL.n19 VTAIL.n18 585
R46 VTAIL.n4 VTAIL.n3 585
R47 VTAIL.n25 VTAIL.n24 585
R48 VTAIL.n89 VTAIL.n88 585
R49 VTAIL.n68 VTAIL.n67 585
R50 VTAIL.n83 VTAIL.n82 585
R51 VTAIL.n81 VTAIL.n80 585
R52 VTAIL.n72 VTAIL.n71 585
R53 VTAIL.n75 VTAIL.n74 585
R54 VTAIL.n59 VTAIL.n58 585
R55 VTAIL.n38 VTAIL.n37 585
R56 VTAIL.n53 VTAIL.n52 585
R57 VTAIL.n51 VTAIL.n50 585
R58 VTAIL.n42 VTAIL.n41 585
R59 VTAIL.n45 VTAIL.n44 585
R60 VTAIL.t6 VTAIL.n73 329.435
R61 VTAIL.t14 VTAIL.n99 329.435
R62 VTAIL.t8 VTAIL.n9 329.435
R63 VTAIL.t13 VTAIL.n43 329.435
R64 VTAIL.n100 VTAIL.n97 171.744
R65 VTAIL.n107 VTAIL.n97 171.744
R66 VTAIL.n108 VTAIL.n107 171.744
R67 VTAIL.n108 VTAIL.n93 171.744
R68 VTAIL.n115 VTAIL.n93 171.744
R69 VTAIL.n10 VTAIL.n7 171.744
R70 VTAIL.n17 VTAIL.n7 171.744
R71 VTAIL.n18 VTAIL.n17 171.744
R72 VTAIL.n18 VTAIL.n3 171.744
R73 VTAIL.n25 VTAIL.n3 171.744
R74 VTAIL.n89 VTAIL.n67 171.744
R75 VTAIL.n82 VTAIL.n67 171.744
R76 VTAIL.n82 VTAIL.n81 171.744
R77 VTAIL.n81 VTAIL.n71 171.744
R78 VTAIL.n74 VTAIL.n71 171.744
R79 VTAIL.n59 VTAIL.n37 171.744
R80 VTAIL.n52 VTAIL.n37 171.744
R81 VTAIL.n52 VTAIL.n51 171.744
R82 VTAIL.n51 VTAIL.n41 171.744
R83 VTAIL.n44 VTAIL.n41 171.744
R84 VTAIL.n100 VTAIL.t14 85.8723
R85 VTAIL.n10 VTAIL.t8 85.8723
R86 VTAIL.n74 VTAIL.t6 85.8723
R87 VTAIL.n44 VTAIL.t13 85.8723
R88 VTAIL.n65 VTAIL.n64 84.0869
R89 VTAIL.n63 VTAIL.n62 84.0869
R90 VTAIL.n35 VTAIL.n34 84.0869
R91 VTAIL.n33 VTAIL.n32 84.0869
R92 VTAIL.n119 VTAIL.n118 84.0868
R93 VTAIL.n1 VTAIL.n0 84.0868
R94 VTAIL.n29 VTAIL.n28 84.0868
R95 VTAIL.n31 VTAIL.n30 84.0868
R96 VTAIL.n117 VTAIL.n116 34.5126
R97 VTAIL.n27 VTAIL.n26 34.5126
R98 VTAIL.n91 VTAIL.n90 34.5126
R99 VTAIL.n61 VTAIL.n60 34.5126
R100 VTAIL.n33 VTAIL.n31 18.4531
R101 VTAIL.n117 VTAIL.n91 17.6255
R102 VTAIL.n114 VTAIL.n92 11.249
R103 VTAIL.n24 VTAIL.n2 11.249
R104 VTAIL.n88 VTAIL.n66 11.249
R105 VTAIL.n58 VTAIL.n36 11.249
R106 VTAIL.n101 VTAIL.n99 10.7185
R107 VTAIL.n11 VTAIL.n9 10.7185
R108 VTAIL.n75 VTAIL.n73 10.7185
R109 VTAIL.n45 VTAIL.n43 10.7185
R110 VTAIL.n113 VTAIL.n94 10.4732
R111 VTAIL.n23 VTAIL.n4 10.4732
R112 VTAIL.n87 VTAIL.n68 10.4732
R113 VTAIL.n57 VTAIL.n38 10.4732
R114 VTAIL.n110 VTAIL.n109 9.69747
R115 VTAIL.n20 VTAIL.n19 9.69747
R116 VTAIL.n84 VTAIL.n83 9.69747
R117 VTAIL.n54 VTAIL.n53 9.69747
R118 VTAIL.n112 VTAIL.n92 9.45567
R119 VTAIL.n22 VTAIL.n2 9.45567
R120 VTAIL.n86 VTAIL.n66 9.45567
R121 VTAIL.n56 VTAIL.n36 9.45567
R122 VTAIL.n103 VTAIL.n102 9.3005
R123 VTAIL.n105 VTAIL.n104 9.3005
R124 VTAIL.n96 VTAIL.n95 9.3005
R125 VTAIL.n111 VTAIL.n110 9.3005
R126 VTAIL.n113 VTAIL.n112 9.3005
R127 VTAIL.n13 VTAIL.n12 9.3005
R128 VTAIL.n15 VTAIL.n14 9.3005
R129 VTAIL.n6 VTAIL.n5 9.3005
R130 VTAIL.n21 VTAIL.n20 9.3005
R131 VTAIL.n23 VTAIL.n22 9.3005
R132 VTAIL.n87 VTAIL.n86 9.3005
R133 VTAIL.n85 VTAIL.n84 9.3005
R134 VTAIL.n70 VTAIL.n69 9.3005
R135 VTAIL.n79 VTAIL.n78 9.3005
R136 VTAIL.n77 VTAIL.n76 9.3005
R137 VTAIL.n49 VTAIL.n48 9.3005
R138 VTAIL.n40 VTAIL.n39 9.3005
R139 VTAIL.n55 VTAIL.n54 9.3005
R140 VTAIL.n57 VTAIL.n56 9.3005
R141 VTAIL.n47 VTAIL.n46 9.3005
R142 VTAIL.n106 VTAIL.n96 8.92171
R143 VTAIL.n16 VTAIL.n6 8.92171
R144 VTAIL.n80 VTAIL.n70 8.92171
R145 VTAIL.n50 VTAIL.n40 8.92171
R146 VTAIL.n105 VTAIL.n98 8.14595
R147 VTAIL.n15 VTAIL.n8 8.14595
R148 VTAIL.n79 VTAIL.n72 8.14595
R149 VTAIL.n49 VTAIL.n42 8.14595
R150 VTAIL.n102 VTAIL.n101 7.3702
R151 VTAIL.n12 VTAIL.n11 7.3702
R152 VTAIL.n76 VTAIL.n75 7.3702
R153 VTAIL.n46 VTAIL.n45 7.3702
R154 VTAIL.n118 VTAIL.t11 6.32443
R155 VTAIL.n118 VTAIL.t10 6.32443
R156 VTAIL.n0 VTAIL.t15 6.32443
R157 VTAIL.n0 VTAIL.t12 6.32443
R158 VTAIL.n28 VTAIL.t3 6.32443
R159 VTAIL.n28 VTAIL.t0 6.32443
R160 VTAIL.n30 VTAIL.t2 6.32443
R161 VTAIL.n30 VTAIL.t5 6.32443
R162 VTAIL.n64 VTAIL.t9 6.32443
R163 VTAIL.n64 VTAIL.t4 6.32443
R164 VTAIL.n62 VTAIL.t7 6.32443
R165 VTAIL.n62 VTAIL.t1 6.32443
R166 VTAIL.n34 VTAIL.t16 6.32443
R167 VTAIL.n34 VTAIL.t18 6.32443
R168 VTAIL.n32 VTAIL.t19 6.32443
R169 VTAIL.n32 VTAIL.t17 6.32443
R170 VTAIL.n102 VTAIL.n98 5.81868
R171 VTAIL.n12 VTAIL.n8 5.81868
R172 VTAIL.n76 VTAIL.n72 5.81868
R173 VTAIL.n46 VTAIL.n42 5.81868
R174 VTAIL.n106 VTAIL.n105 5.04292
R175 VTAIL.n16 VTAIL.n15 5.04292
R176 VTAIL.n80 VTAIL.n79 5.04292
R177 VTAIL.n50 VTAIL.n49 5.04292
R178 VTAIL.n109 VTAIL.n96 4.26717
R179 VTAIL.n19 VTAIL.n6 4.26717
R180 VTAIL.n83 VTAIL.n70 4.26717
R181 VTAIL.n53 VTAIL.n40 4.26717
R182 VTAIL.n110 VTAIL.n94 3.49141
R183 VTAIL.n20 VTAIL.n4 3.49141
R184 VTAIL.n84 VTAIL.n68 3.49141
R185 VTAIL.n54 VTAIL.n38 3.49141
R186 VTAIL.n114 VTAIL.n113 2.71565
R187 VTAIL.n24 VTAIL.n23 2.71565
R188 VTAIL.n88 VTAIL.n87 2.71565
R189 VTAIL.n58 VTAIL.n57 2.71565
R190 VTAIL.n103 VTAIL.n99 2.41827
R191 VTAIL.n13 VTAIL.n9 2.41827
R192 VTAIL.n77 VTAIL.n73 2.41827
R193 VTAIL.n47 VTAIL.n43 2.41827
R194 VTAIL.n116 VTAIL.n92 1.93989
R195 VTAIL.n26 VTAIL.n2 1.93989
R196 VTAIL.n90 VTAIL.n66 1.93989
R197 VTAIL.n60 VTAIL.n36 1.93989
R198 VTAIL.n63 VTAIL.n61 0.884121
R199 VTAIL.n27 VTAIL.n1 0.884121
R200 VTAIL.n35 VTAIL.n33 0.828086
R201 VTAIL.n61 VTAIL.n35 0.828086
R202 VTAIL.n65 VTAIL.n63 0.828086
R203 VTAIL.n91 VTAIL.n65 0.828086
R204 VTAIL.n31 VTAIL.n29 0.828086
R205 VTAIL.n29 VTAIL.n27 0.828086
R206 VTAIL.n119 VTAIL.n117 0.828086
R207 VTAIL VTAIL.n1 0.679379
R208 VTAIL.n104 VTAIL.n103 0.155672
R209 VTAIL.n104 VTAIL.n95 0.155672
R210 VTAIL.n111 VTAIL.n95 0.155672
R211 VTAIL.n112 VTAIL.n111 0.155672
R212 VTAIL.n14 VTAIL.n13 0.155672
R213 VTAIL.n14 VTAIL.n5 0.155672
R214 VTAIL.n21 VTAIL.n5 0.155672
R215 VTAIL.n22 VTAIL.n21 0.155672
R216 VTAIL.n86 VTAIL.n85 0.155672
R217 VTAIL.n85 VTAIL.n69 0.155672
R218 VTAIL.n78 VTAIL.n69 0.155672
R219 VTAIL.n78 VTAIL.n77 0.155672
R220 VTAIL.n56 VTAIL.n55 0.155672
R221 VTAIL.n55 VTAIL.n39 0.155672
R222 VTAIL.n48 VTAIL.n39 0.155672
R223 VTAIL.n48 VTAIL.n47 0.155672
R224 VTAIL VTAIL.n119 0.149207
R225 VDD2.n53 VDD2.n52 756.745
R226 VDD2.n24 VDD2.n23 756.745
R227 VDD2.n52 VDD2.n51 585
R228 VDD2.n31 VDD2.n30 585
R229 VDD2.n46 VDD2.n45 585
R230 VDD2.n44 VDD2.n43 585
R231 VDD2.n35 VDD2.n34 585
R232 VDD2.n38 VDD2.n37 585
R233 VDD2.n9 VDD2.n8 585
R234 VDD2.n6 VDD2.n5 585
R235 VDD2.n15 VDD2.n14 585
R236 VDD2.n17 VDD2.n16 585
R237 VDD2.n2 VDD2.n1 585
R238 VDD2.n23 VDD2.n22 585
R239 VDD2.t4 VDD2.n36 329.435
R240 VDD2.t9 VDD2.n7 329.435
R241 VDD2.n52 VDD2.n30 171.744
R242 VDD2.n45 VDD2.n30 171.744
R243 VDD2.n45 VDD2.n44 171.744
R244 VDD2.n44 VDD2.n34 171.744
R245 VDD2.n37 VDD2.n34 171.744
R246 VDD2.n8 VDD2.n5 171.744
R247 VDD2.n15 VDD2.n5 171.744
R248 VDD2.n16 VDD2.n15 171.744
R249 VDD2.n16 VDD2.n1 171.744
R250 VDD2.n23 VDD2.n1 171.744
R251 VDD2.n28 VDD2.n27 101.331
R252 VDD2 VDD2.n57 101.328
R253 VDD2.n56 VDD2.n55 100.766
R254 VDD2.n26 VDD2.n25 100.766
R255 VDD2.n37 VDD2.t4 85.8723
R256 VDD2.n8 VDD2.t9 85.8723
R257 VDD2.n26 VDD2.n24 52.019
R258 VDD2.n54 VDD2.n53 51.1914
R259 VDD2.n54 VDD2.n28 32.0774
R260 VDD2.n51 VDD2.n29 11.249
R261 VDD2.n22 VDD2.n0 11.249
R262 VDD2.n38 VDD2.n36 10.7185
R263 VDD2.n9 VDD2.n7 10.7185
R264 VDD2.n50 VDD2.n31 10.4732
R265 VDD2.n21 VDD2.n2 10.4732
R266 VDD2.n47 VDD2.n46 9.69747
R267 VDD2.n18 VDD2.n17 9.69747
R268 VDD2.n49 VDD2.n29 9.45567
R269 VDD2.n20 VDD2.n0 9.45567
R270 VDD2.n42 VDD2.n41 9.3005
R271 VDD2.n33 VDD2.n32 9.3005
R272 VDD2.n48 VDD2.n47 9.3005
R273 VDD2.n50 VDD2.n49 9.3005
R274 VDD2.n40 VDD2.n39 9.3005
R275 VDD2.n11 VDD2.n10 9.3005
R276 VDD2.n13 VDD2.n12 9.3005
R277 VDD2.n4 VDD2.n3 9.3005
R278 VDD2.n19 VDD2.n18 9.3005
R279 VDD2.n21 VDD2.n20 9.3005
R280 VDD2.n43 VDD2.n33 8.92171
R281 VDD2.n14 VDD2.n4 8.92171
R282 VDD2.n42 VDD2.n35 8.14595
R283 VDD2.n13 VDD2.n6 8.14595
R284 VDD2.n39 VDD2.n38 7.3702
R285 VDD2.n10 VDD2.n9 7.3702
R286 VDD2.n57 VDD2.t6 6.32443
R287 VDD2.n57 VDD2.t7 6.32443
R288 VDD2.n55 VDD2.t3 6.32443
R289 VDD2.n55 VDD2.t5 6.32443
R290 VDD2.n27 VDD2.t8 6.32443
R291 VDD2.n27 VDD2.t1 6.32443
R292 VDD2.n25 VDD2.t2 6.32443
R293 VDD2.n25 VDD2.t0 6.32443
R294 VDD2.n39 VDD2.n35 5.81868
R295 VDD2.n10 VDD2.n6 5.81868
R296 VDD2.n43 VDD2.n42 5.04292
R297 VDD2.n14 VDD2.n13 5.04292
R298 VDD2.n46 VDD2.n33 4.26717
R299 VDD2.n17 VDD2.n4 4.26717
R300 VDD2.n47 VDD2.n31 3.49141
R301 VDD2.n18 VDD2.n2 3.49141
R302 VDD2.n51 VDD2.n50 2.71565
R303 VDD2.n22 VDD2.n21 2.71565
R304 VDD2.n40 VDD2.n36 2.41827
R305 VDD2.n11 VDD2.n7 2.41827
R306 VDD2.n53 VDD2.n29 1.93989
R307 VDD2.n24 VDD2.n0 1.93989
R308 VDD2.n56 VDD2.n54 0.828086
R309 VDD2 VDD2.n56 0.265586
R310 VDD2.n49 VDD2.n48 0.155672
R311 VDD2.n48 VDD2.n32 0.155672
R312 VDD2.n41 VDD2.n32 0.155672
R313 VDD2.n41 VDD2.n40 0.155672
R314 VDD2.n12 VDD2.n11 0.155672
R315 VDD2.n12 VDD2.n3 0.155672
R316 VDD2.n19 VDD2.n3 0.155672
R317 VDD2.n20 VDD2.n19 0.155672
R318 VDD2.n28 VDD2.n26 0.152051
R319 VP.n4 VP.t6 285.8
R320 VP.n10 VP.t9 258.979
R321 VP.n1 VP.t2 258.979
R322 VP.n14 VP.t0 258.979
R323 VP.n15 VP.t7 258.979
R324 VP.n16 VP.t1 258.979
R325 VP.n8 VP.t3 258.979
R326 VP.n7 VP.t4 258.979
R327 VP.n6 VP.t5 258.979
R328 VP.n5 VP.t8 258.979
R329 VP.n17 VP.n16 161.3
R330 VP.n9 VP.n8 161.3
R331 VP.n11 VP.n10 161.3
R332 VP.n6 VP.n3 80.6037
R333 VP.n7 VP.n2 80.6037
R334 VP.n15 VP.n0 80.6037
R335 VP.n14 VP.n13 80.6037
R336 VP.n12 VP.n1 80.6037
R337 VP.n10 VP.n1 48.2005
R338 VP.n14 VP.n1 48.2005
R339 VP.n15 VP.n14 48.2005
R340 VP.n16 VP.n15 48.2005
R341 VP.n8 VP.n7 48.2005
R342 VP.n7 VP.n6 48.2005
R343 VP.n6 VP.n5 48.2005
R344 VP.n4 VP.n3 45.2318
R345 VP.n11 VP.n9 37.2732
R346 VP.n5 VP.n4 13.3799
R347 VP.n3 VP.n2 0.380177
R348 VP.n13 VP.n12 0.380177
R349 VP.n13 VP.n0 0.380177
R350 VP.n9 VP.n2 0.285035
R351 VP.n12 VP.n11 0.285035
R352 VP.n17 VP.n0 0.285035
R353 VP VP.n17 0.0516364
R354 VDD1.n24 VDD1.n23 756.745
R355 VDD1.n51 VDD1.n50 756.745
R356 VDD1.n23 VDD1.n22 585
R357 VDD1.n2 VDD1.n1 585
R358 VDD1.n17 VDD1.n16 585
R359 VDD1.n15 VDD1.n14 585
R360 VDD1.n6 VDD1.n5 585
R361 VDD1.n9 VDD1.n8 585
R362 VDD1.n36 VDD1.n35 585
R363 VDD1.n33 VDD1.n32 585
R364 VDD1.n42 VDD1.n41 585
R365 VDD1.n44 VDD1.n43 585
R366 VDD1.n29 VDD1.n28 585
R367 VDD1.n50 VDD1.n49 585
R368 VDD1.t3 VDD1.n7 329.435
R369 VDD1.t0 VDD1.n34 329.435
R370 VDD1.n23 VDD1.n1 171.744
R371 VDD1.n16 VDD1.n1 171.744
R372 VDD1.n16 VDD1.n15 171.744
R373 VDD1.n15 VDD1.n5 171.744
R374 VDD1.n8 VDD1.n5 171.744
R375 VDD1.n35 VDD1.n32 171.744
R376 VDD1.n42 VDD1.n32 171.744
R377 VDD1.n43 VDD1.n42 171.744
R378 VDD1.n43 VDD1.n28 171.744
R379 VDD1.n50 VDD1.n28 171.744
R380 VDD1.n55 VDD1.n54 101.331
R381 VDD1.n26 VDD1.n25 100.766
R382 VDD1.n53 VDD1.n52 100.766
R383 VDD1.n57 VDD1.n56 100.764
R384 VDD1.n8 VDD1.t3 85.8723
R385 VDD1.n35 VDD1.t0 85.8723
R386 VDD1.n26 VDD1.n24 52.019
R387 VDD1.n53 VDD1.n51 52.019
R388 VDD1.n57 VDD1.n55 33.0742
R389 VDD1.n22 VDD1.n0 11.249
R390 VDD1.n49 VDD1.n27 11.249
R391 VDD1.n9 VDD1.n7 10.7185
R392 VDD1.n36 VDD1.n34 10.7185
R393 VDD1.n21 VDD1.n2 10.4732
R394 VDD1.n48 VDD1.n29 10.4732
R395 VDD1.n18 VDD1.n17 9.69747
R396 VDD1.n45 VDD1.n44 9.69747
R397 VDD1.n20 VDD1.n0 9.45567
R398 VDD1.n47 VDD1.n27 9.45567
R399 VDD1.n13 VDD1.n12 9.3005
R400 VDD1.n4 VDD1.n3 9.3005
R401 VDD1.n19 VDD1.n18 9.3005
R402 VDD1.n21 VDD1.n20 9.3005
R403 VDD1.n11 VDD1.n10 9.3005
R404 VDD1.n38 VDD1.n37 9.3005
R405 VDD1.n40 VDD1.n39 9.3005
R406 VDD1.n31 VDD1.n30 9.3005
R407 VDD1.n46 VDD1.n45 9.3005
R408 VDD1.n48 VDD1.n47 9.3005
R409 VDD1.n14 VDD1.n4 8.92171
R410 VDD1.n41 VDD1.n31 8.92171
R411 VDD1.n13 VDD1.n6 8.14595
R412 VDD1.n40 VDD1.n33 8.14595
R413 VDD1.n10 VDD1.n9 7.3702
R414 VDD1.n37 VDD1.n36 7.3702
R415 VDD1.n56 VDD1.t5 6.32443
R416 VDD1.n56 VDD1.t6 6.32443
R417 VDD1.n25 VDD1.t1 6.32443
R418 VDD1.n25 VDD1.t4 6.32443
R419 VDD1.n54 VDD1.t2 6.32443
R420 VDD1.n54 VDD1.t8 6.32443
R421 VDD1.n52 VDD1.t7 6.32443
R422 VDD1.n52 VDD1.t9 6.32443
R423 VDD1.n10 VDD1.n6 5.81868
R424 VDD1.n37 VDD1.n33 5.81868
R425 VDD1.n14 VDD1.n13 5.04292
R426 VDD1.n41 VDD1.n40 5.04292
R427 VDD1.n17 VDD1.n4 4.26717
R428 VDD1.n44 VDD1.n31 4.26717
R429 VDD1.n18 VDD1.n2 3.49141
R430 VDD1.n45 VDD1.n29 3.49141
R431 VDD1.n22 VDD1.n21 2.71565
R432 VDD1.n49 VDD1.n48 2.71565
R433 VDD1.n11 VDD1.n7 2.41827
R434 VDD1.n38 VDD1.n34 2.41827
R435 VDD1.n24 VDD1.n0 1.93989
R436 VDD1.n51 VDD1.n27 1.93989
R437 VDD1 VDD1.n57 0.563
R438 VDD1 VDD1.n26 0.265586
R439 VDD1.n20 VDD1.n19 0.155672
R440 VDD1.n19 VDD1.n3 0.155672
R441 VDD1.n12 VDD1.n3 0.155672
R442 VDD1.n12 VDD1.n11 0.155672
R443 VDD1.n39 VDD1.n38 0.155672
R444 VDD1.n39 VDD1.n30 0.155672
R445 VDD1.n46 VDD1.n30 0.155672
R446 VDD1.n47 VDD1.n46 0.155672
R447 VDD1.n55 VDD1.n53 0.152051
R448 B.n306 B.n305 585
R449 B.n307 B.n44 585
R450 B.n309 B.n308 585
R451 B.n310 B.n43 585
R452 B.n312 B.n311 585
R453 B.n313 B.n42 585
R454 B.n315 B.n314 585
R455 B.n316 B.n41 585
R456 B.n318 B.n317 585
R457 B.n319 B.n40 585
R458 B.n321 B.n320 585
R459 B.n322 B.n39 585
R460 B.n324 B.n323 585
R461 B.n325 B.n38 585
R462 B.n327 B.n326 585
R463 B.n328 B.n37 585
R464 B.n330 B.n329 585
R465 B.n331 B.n36 585
R466 B.n333 B.n332 585
R467 B.n334 B.n35 585
R468 B.n336 B.n335 585
R469 B.n338 B.n337 585
R470 B.n339 B.n31 585
R471 B.n341 B.n340 585
R472 B.n342 B.n30 585
R473 B.n344 B.n343 585
R474 B.n345 B.n29 585
R475 B.n347 B.n346 585
R476 B.n348 B.n28 585
R477 B.n350 B.n349 585
R478 B.n351 B.n25 585
R479 B.n354 B.n353 585
R480 B.n355 B.n24 585
R481 B.n357 B.n356 585
R482 B.n358 B.n23 585
R483 B.n360 B.n359 585
R484 B.n361 B.n22 585
R485 B.n363 B.n362 585
R486 B.n364 B.n21 585
R487 B.n366 B.n365 585
R488 B.n367 B.n20 585
R489 B.n369 B.n368 585
R490 B.n370 B.n19 585
R491 B.n372 B.n371 585
R492 B.n373 B.n18 585
R493 B.n375 B.n374 585
R494 B.n376 B.n17 585
R495 B.n378 B.n377 585
R496 B.n379 B.n16 585
R497 B.n381 B.n380 585
R498 B.n382 B.n15 585
R499 B.n384 B.n383 585
R500 B.n304 B.n45 585
R501 B.n303 B.n302 585
R502 B.n301 B.n46 585
R503 B.n300 B.n299 585
R504 B.n298 B.n47 585
R505 B.n297 B.n296 585
R506 B.n295 B.n48 585
R507 B.n294 B.n293 585
R508 B.n292 B.n49 585
R509 B.n291 B.n290 585
R510 B.n289 B.n50 585
R511 B.n288 B.n287 585
R512 B.n286 B.n51 585
R513 B.n285 B.n284 585
R514 B.n283 B.n52 585
R515 B.n282 B.n281 585
R516 B.n280 B.n53 585
R517 B.n279 B.n278 585
R518 B.n277 B.n54 585
R519 B.n276 B.n275 585
R520 B.n274 B.n55 585
R521 B.n273 B.n272 585
R522 B.n271 B.n56 585
R523 B.n270 B.n269 585
R524 B.n268 B.n57 585
R525 B.n267 B.n266 585
R526 B.n265 B.n58 585
R527 B.n264 B.n263 585
R528 B.n262 B.n59 585
R529 B.n261 B.n260 585
R530 B.n259 B.n60 585
R531 B.n258 B.n257 585
R532 B.n256 B.n61 585
R533 B.n255 B.n254 585
R534 B.n253 B.n62 585
R535 B.n252 B.n251 585
R536 B.n250 B.n63 585
R537 B.n249 B.n248 585
R538 B.n247 B.n64 585
R539 B.n246 B.n245 585
R540 B.n244 B.n65 585
R541 B.n243 B.n242 585
R542 B.n241 B.n66 585
R543 B.n240 B.n239 585
R544 B.n238 B.n67 585
R545 B.n237 B.n236 585
R546 B.n235 B.n68 585
R547 B.n234 B.n233 585
R548 B.n232 B.n69 585
R549 B.n231 B.n230 585
R550 B.n229 B.n70 585
R551 B.n150 B.n149 585
R552 B.n151 B.n100 585
R553 B.n153 B.n152 585
R554 B.n154 B.n99 585
R555 B.n156 B.n155 585
R556 B.n157 B.n98 585
R557 B.n159 B.n158 585
R558 B.n160 B.n97 585
R559 B.n162 B.n161 585
R560 B.n163 B.n96 585
R561 B.n165 B.n164 585
R562 B.n166 B.n95 585
R563 B.n168 B.n167 585
R564 B.n169 B.n94 585
R565 B.n171 B.n170 585
R566 B.n172 B.n93 585
R567 B.n174 B.n173 585
R568 B.n175 B.n92 585
R569 B.n177 B.n176 585
R570 B.n178 B.n91 585
R571 B.n180 B.n179 585
R572 B.n182 B.n181 585
R573 B.n183 B.n87 585
R574 B.n185 B.n184 585
R575 B.n186 B.n86 585
R576 B.n188 B.n187 585
R577 B.n189 B.n85 585
R578 B.n191 B.n190 585
R579 B.n192 B.n84 585
R580 B.n194 B.n193 585
R581 B.n195 B.n81 585
R582 B.n198 B.n197 585
R583 B.n199 B.n80 585
R584 B.n201 B.n200 585
R585 B.n202 B.n79 585
R586 B.n204 B.n203 585
R587 B.n205 B.n78 585
R588 B.n207 B.n206 585
R589 B.n208 B.n77 585
R590 B.n210 B.n209 585
R591 B.n211 B.n76 585
R592 B.n213 B.n212 585
R593 B.n214 B.n75 585
R594 B.n216 B.n215 585
R595 B.n217 B.n74 585
R596 B.n219 B.n218 585
R597 B.n220 B.n73 585
R598 B.n222 B.n221 585
R599 B.n223 B.n72 585
R600 B.n225 B.n224 585
R601 B.n226 B.n71 585
R602 B.n228 B.n227 585
R603 B.n148 B.n101 585
R604 B.n147 B.n146 585
R605 B.n145 B.n102 585
R606 B.n144 B.n143 585
R607 B.n142 B.n103 585
R608 B.n141 B.n140 585
R609 B.n139 B.n104 585
R610 B.n138 B.n137 585
R611 B.n136 B.n105 585
R612 B.n135 B.n134 585
R613 B.n133 B.n106 585
R614 B.n132 B.n131 585
R615 B.n130 B.n107 585
R616 B.n129 B.n128 585
R617 B.n127 B.n108 585
R618 B.n126 B.n125 585
R619 B.n124 B.n109 585
R620 B.n123 B.n122 585
R621 B.n121 B.n110 585
R622 B.n120 B.n119 585
R623 B.n118 B.n111 585
R624 B.n117 B.n116 585
R625 B.n115 B.n112 585
R626 B.n114 B.n113 585
R627 B.n2 B.n0 585
R628 B.n421 B.n1 585
R629 B.n420 B.n419 585
R630 B.n418 B.n3 585
R631 B.n417 B.n416 585
R632 B.n415 B.n4 585
R633 B.n414 B.n413 585
R634 B.n412 B.n5 585
R635 B.n411 B.n410 585
R636 B.n409 B.n6 585
R637 B.n408 B.n407 585
R638 B.n406 B.n7 585
R639 B.n405 B.n404 585
R640 B.n403 B.n8 585
R641 B.n402 B.n401 585
R642 B.n400 B.n9 585
R643 B.n399 B.n398 585
R644 B.n397 B.n10 585
R645 B.n396 B.n395 585
R646 B.n394 B.n11 585
R647 B.n393 B.n392 585
R648 B.n391 B.n12 585
R649 B.n390 B.n389 585
R650 B.n388 B.n13 585
R651 B.n387 B.n386 585
R652 B.n385 B.n14 585
R653 B.n423 B.n422 585
R654 B.n150 B.n101 545.355
R655 B.n385 B.n384 545.355
R656 B.n229 B.n228 545.355
R657 B.n306 B.n45 545.355
R658 B.n82 B.t3 400.546
R659 B.n88 B.t6 400.546
R660 B.n26 B.t9 400.546
R661 B.n32 B.t0 400.546
R662 B.n82 B.t5 271.551
R663 B.n32 B.t1 271.551
R664 B.n88 B.t8 271.551
R665 B.n26 B.t10 271.551
R666 B.n83 B.t4 252.934
R667 B.n33 B.t2 252.934
R668 B.n89 B.t7 252.934
R669 B.n27 B.t11 252.934
R670 B.n146 B.n101 163.367
R671 B.n146 B.n145 163.367
R672 B.n145 B.n144 163.367
R673 B.n144 B.n103 163.367
R674 B.n140 B.n103 163.367
R675 B.n140 B.n139 163.367
R676 B.n139 B.n138 163.367
R677 B.n138 B.n105 163.367
R678 B.n134 B.n105 163.367
R679 B.n134 B.n133 163.367
R680 B.n133 B.n132 163.367
R681 B.n132 B.n107 163.367
R682 B.n128 B.n107 163.367
R683 B.n128 B.n127 163.367
R684 B.n127 B.n126 163.367
R685 B.n126 B.n109 163.367
R686 B.n122 B.n109 163.367
R687 B.n122 B.n121 163.367
R688 B.n121 B.n120 163.367
R689 B.n120 B.n111 163.367
R690 B.n116 B.n111 163.367
R691 B.n116 B.n115 163.367
R692 B.n115 B.n114 163.367
R693 B.n114 B.n2 163.367
R694 B.n422 B.n2 163.367
R695 B.n422 B.n421 163.367
R696 B.n421 B.n420 163.367
R697 B.n420 B.n3 163.367
R698 B.n416 B.n3 163.367
R699 B.n416 B.n415 163.367
R700 B.n415 B.n414 163.367
R701 B.n414 B.n5 163.367
R702 B.n410 B.n5 163.367
R703 B.n410 B.n409 163.367
R704 B.n409 B.n408 163.367
R705 B.n408 B.n7 163.367
R706 B.n404 B.n7 163.367
R707 B.n404 B.n403 163.367
R708 B.n403 B.n402 163.367
R709 B.n402 B.n9 163.367
R710 B.n398 B.n9 163.367
R711 B.n398 B.n397 163.367
R712 B.n397 B.n396 163.367
R713 B.n396 B.n11 163.367
R714 B.n392 B.n11 163.367
R715 B.n392 B.n391 163.367
R716 B.n391 B.n390 163.367
R717 B.n390 B.n13 163.367
R718 B.n386 B.n13 163.367
R719 B.n386 B.n385 163.367
R720 B.n151 B.n150 163.367
R721 B.n152 B.n151 163.367
R722 B.n152 B.n99 163.367
R723 B.n156 B.n99 163.367
R724 B.n157 B.n156 163.367
R725 B.n158 B.n157 163.367
R726 B.n158 B.n97 163.367
R727 B.n162 B.n97 163.367
R728 B.n163 B.n162 163.367
R729 B.n164 B.n163 163.367
R730 B.n164 B.n95 163.367
R731 B.n168 B.n95 163.367
R732 B.n169 B.n168 163.367
R733 B.n170 B.n169 163.367
R734 B.n170 B.n93 163.367
R735 B.n174 B.n93 163.367
R736 B.n175 B.n174 163.367
R737 B.n176 B.n175 163.367
R738 B.n176 B.n91 163.367
R739 B.n180 B.n91 163.367
R740 B.n181 B.n180 163.367
R741 B.n181 B.n87 163.367
R742 B.n185 B.n87 163.367
R743 B.n186 B.n185 163.367
R744 B.n187 B.n186 163.367
R745 B.n187 B.n85 163.367
R746 B.n191 B.n85 163.367
R747 B.n192 B.n191 163.367
R748 B.n193 B.n192 163.367
R749 B.n193 B.n81 163.367
R750 B.n198 B.n81 163.367
R751 B.n199 B.n198 163.367
R752 B.n200 B.n199 163.367
R753 B.n200 B.n79 163.367
R754 B.n204 B.n79 163.367
R755 B.n205 B.n204 163.367
R756 B.n206 B.n205 163.367
R757 B.n206 B.n77 163.367
R758 B.n210 B.n77 163.367
R759 B.n211 B.n210 163.367
R760 B.n212 B.n211 163.367
R761 B.n212 B.n75 163.367
R762 B.n216 B.n75 163.367
R763 B.n217 B.n216 163.367
R764 B.n218 B.n217 163.367
R765 B.n218 B.n73 163.367
R766 B.n222 B.n73 163.367
R767 B.n223 B.n222 163.367
R768 B.n224 B.n223 163.367
R769 B.n224 B.n71 163.367
R770 B.n228 B.n71 163.367
R771 B.n230 B.n229 163.367
R772 B.n230 B.n69 163.367
R773 B.n234 B.n69 163.367
R774 B.n235 B.n234 163.367
R775 B.n236 B.n235 163.367
R776 B.n236 B.n67 163.367
R777 B.n240 B.n67 163.367
R778 B.n241 B.n240 163.367
R779 B.n242 B.n241 163.367
R780 B.n242 B.n65 163.367
R781 B.n246 B.n65 163.367
R782 B.n247 B.n246 163.367
R783 B.n248 B.n247 163.367
R784 B.n248 B.n63 163.367
R785 B.n252 B.n63 163.367
R786 B.n253 B.n252 163.367
R787 B.n254 B.n253 163.367
R788 B.n254 B.n61 163.367
R789 B.n258 B.n61 163.367
R790 B.n259 B.n258 163.367
R791 B.n260 B.n259 163.367
R792 B.n260 B.n59 163.367
R793 B.n264 B.n59 163.367
R794 B.n265 B.n264 163.367
R795 B.n266 B.n265 163.367
R796 B.n266 B.n57 163.367
R797 B.n270 B.n57 163.367
R798 B.n271 B.n270 163.367
R799 B.n272 B.n271 163.367
R800 B.n272 B.n55 163.367
R801 B.n276 B.n55 163.367
R802 B.n277 B.n276 163.367
R803 B.n278 B.n277 163.367
R804 B.n278 B.n53 163.367
R805 B.n282 B.n53 163.367
R806 B.n283 B.n282 163.367
R807 B.n284 B.n283 163.367
R808 B.n284 B.n51 163.367
R809 B.n288 B.n51 163.367
R810 B.n289 B.n288 163.367
R811 B.n290 B.n289 163.367
R812 B.n290 B.n49 163.367
R813 B.n294 B.n49 163.367
R814 B.n295 B.n294 163.367
R815 B.n296 B.n295 163.367
R816 B.n296 B.n47 163.367
R817 B.n300 B.n47 163.367
R818 B.n301 B.n300 163.367
R819 B.n302 B.n301 163.367
R820 B.n302 B.n45 163.367
R821 B.n384 B.n15 163.367
R822 B.n380 B.n15 163.367
R823 B.n380 B.n379 163.367
R824 B.n379 B.n378 163.367
R825 B.n378 B.n17 163.367
R826 B.n374 B.n17 163.367
R827 B.n374 B.n373 163.367
R828 B.n373 B.n372 163.367
R829 B.n372 B.n19 163.367
R830 B.n368 B.n19 163.367
R831 B.n368 B.n367 163.367
R832 B.n367 B.n366 163.367
R833 B.n366 B.n21 163.367
R834 B.n362 B.n21 163.367
R835 B.n362 B.n361 163.367
R836 B.n361 B.n360 163.367
R837 B.n360 B.n23 163.367
R838 B.n356 B.n23 163.367
R839 B.n356 B.n355 163.367
R840 B.n355 B.n354 163.367
R841 B.n354 B.n25 163.367
R842 B.n349 B.n25 163.367
R843 B.n349 B.n348 163.367
R844 B.n348 B.n347 163.367
R845 B.n347 B.n29 163.367
R846 B.n343 B.n29 163.367
R847 B.n343 B.n342 163.367
R848 B.n342 B.n341 163.367
R849 B.n341 B.n31 163.367
R850 B.n337 B.n31 163.367
R851 B.n337 B.n336 163.367
R852 B.n336 B.n35 163.367
R853 B.n332 B.n35 163.367
R854 B.n332 B.n331 163.367
R855 B.n331 B.n330 163.367
R856 B.n330 B.n37 163.367
R857 B.n326 B.n37 163.367
R858 B.n326 B.n325 163.367
R859 B.n325 B.n324 163.367
R860 B.n324 B.n39 163.367
R861 B.n320 B.n39 163.367
R862 B.n320 B.n319 163.367
R863 B.n319 B.n318 163.367
R864 B.n318 B.n41 163.367
R865 B.n314 B.n41 163.367
R866 B.n314 B.n313 163.367
R867 B.n313 B.n312 163.367
R868 B.n312 B.n43 163.367
R869 B.n308 B.n43 163.367
R870 B.n308 B.n307 163.367
R871 B.n307 B.n306 163.367
R872 B.n196 B.n83 59.5399
R873 B.n90 B.n89 59.5399
R874 B.n352 B.n27 59.5399
R875 B.n34 B.n33 59.5399
R876 B.n383 B.n14 35.4346
R877 B.n305 B.n304 35.4346
R878 B.n227 B.n70 35.4346
R879 B.n149 B.n148 35.4346
R880 B.n83 B.n82 18.6187
R881 B.n89 B.n88 18.6187
R882 B.n27 B.n26 18.6187
R883 B.n33 B.n32 18.6187
R884 B B.n423 18.0485
R885 B.n383 B.n382 10.6151
R886 B.n382 B.n381 10.6151
R887 B.n381 B.n16 10.6151
R888 B.n377 B.n16 10.6151
R889 B.n377 B.n376 10.6151
R890 B.n376 B.n375 10.6151
R891 B.n375 B.n18 10.6151
R892 B.n371 B.n18 10.6151
R893 B.n371 B.n370 10.6151
R894 B.n370 B.n369 10.6151
R895 B.n369 B.n20 10.6151
R896 B.n365 B.n20 10.6151
R897 B.n365 B.n364 10.6151
R898 B.n364 B.n363 10.6151
R899 B.n363 B.n22 10.6151
R900 B.n359 B.n22 10.6151
R901 B.n359 B.n358 10.6151
R902 B.n358 B.n357 10.6151
R903 B.n357 B.n24 10.6151
R904 B.n353 B.n24 10.6151
R905 B.n351 B.n350 10.6151
R906 B.n350 B.n28 10.6151
R907 B.n346 B.n28 10.6151
R908 B.n346 B.n345 10.6151
R909 B.n345 B.n344 10.6151
R910 B.n344 B.n30 10.6151
R911 B.n340 B.n30 10.6151
R912 B.n340 B.n339 10.6151
R913 B.n339 B.n338 10.6151
R914 B.n335 B.n334 10.6151
R915 B.n334 B.n333 10.6151
R916 B.n333 B.n36 10.6151
R917 B.n329 B.n36 10.6151
R918 B.n329 B.n328 10.6151
R919 B.n328 B.n327 10.6151
R920 B.n327 B.n38 10.6151
R921 B.n323 B.n38 10.6151
R922 B.n323 B.n322 10.6151
R923 B.n322 B.n321 10.6151
R924 B.n321 B.n40 10.6151
R925 B.n317 B.n40 10.6151
R926 B.n317 B.n316 10.6151
R927 B.n316 B.n315 10.6151
R928 B.n315 B.n42 10.6151
R929 B.n311 B.n42 10.6151
R930 B.n311 B.n310 10.6151
R931 B.n310 B.n309 10.6151
R932 B.n309 B.n44 10.6151
R933 B.n305 B.n44 10.6151
R934 B.n231 B.n70 10.6151
R935 B.n232 B.n231 10.6151
R936 B.n233 B.n232 10.6151
R937 B.n233 B.n68 10.6151
R938 B.n237 B.n68 10.6151
R939 B.n238 B.n237 10.6151
R940 B.n239 B.n238 10.6151
R941 B.n239 B.n66 10.6151
R942 B.n243 B.n66 10.6151
R943 B.n244 B.n243 10.6151
R944 B.n245 B.n244 10.6151
R945 B.n245 B.n64 10.6151
R946 B.n249 B.n64 10.6151
R947 B.n250 B.n249 10.6151
R948 B.n251 B.n250 10.6151
R949 B.n251 B.n62 10.6151
R950 B.n255 B.n62 10.6151
R951 B.n256 B.n255 10.6151
R952 B.n257 B.n256 10.6151
R953 B.n257 B.n60 10.6151
R954 B.n261 B.n60 10.6151
R955 B.n262 B.n261 10.6151
R956 B.n263 B.n262 10.6151
R957 B.n263 B.n58 10.6151
R958 B.n267 B.n58 10.6151
R959 B.n268 B.n267 10.6151
R960 B.n269 B.n268 10.6151
R961 B.n269 B.n56 10.6151
R962 B.n273 B.n56 10.6151
R963 B.n274 B.n273 10.6151
R964 B.n275 B.n274 10.6151
R965 B.n275 B.n54 10.6151
R966 B.n279 B.n54 10.6151
R967 B.n280 B.n279 10.6151
R968 B.n281 B.n280 10.6151
R969 B.n281 B.n52 10.6151
R970 B.n285 B.n52 10.6151
R971 B.n286 B.n285 10.6151
R972 B.n287 B.n286 10.6151
R973 B.n287 B.n50 10.6151
R974 B.n291 B.n50 10.6151
R975 B.n292 B.n291 10.6151
R976 B.n293 B.n292 10.6151
R977 B.n293 B.n48 10.6151
R978 B.n297 B.n48 10.6151
R979 B.n298 B.n297 10.6151
R980 B.n299 B.n298 10.6151
R981 B.n299 B.n46 10.6151
R982 B.n303 B.n46 10.6151
R983 B.n304 B.n303 10.6151
R984 B.n149 B.n100 10.6151
R985 B.n153 B.n100 10.6151
R986 B.n154 B.n153 10.6151
R987 B.n155 B.n154 10.6151
R988 B.n155 B.n98 10.6151
R989 B.n159 B.n98 10.6151
R990 B.n160 B.n159 10.6151
R991 B.n161 B.n160 10.6151
R992 B.n161 B.n96 10.6151
R993 B.n165 B.n96 10.6151
R994 B.n166 B.n165 10.6151
R995 B.n167 B.n166 10.6151
R996 B.n167 B.n94 10.6151
R997 B.n171 B.n94 10.6151
R998 B.n172 B.n171 10.6151
R999 B.n173 B.n172 10.6151
R1000 B.n173 B.n92 10.6151
R1001 B.n177 B.n92 10.6151
R1002 B.n178 B.n177 10.6151
R1003 B.n179 B.n178 10.6151
R1004 B.n183 B.n182 10.6151
R1005 B.n184 B.n183 10.6151
R1006 B.n184 B.n86 10.6151
R1007 B.n188 B.n86 10.6151
R1008 B.n189 B.n188 10.6151
R1009 B.n190 B.n189 10.6151
R1010 B.n190 B.n84 10.6151
R1011 B.n194 B.n84 10.6151
R1012 B.n195 B.n194 10.6151
R1013 B.n197 B.n80 10.6151
R1014 B.n201 B.n80 10.6151
R1015 B.n202 B.n201 10.6151
R1016 B.n203 B.n202 10.6151
R1017 B.n203 B.n78 10.6151
R1018 B.n207 B.n78 10.6151
R1019 B.n208 B.n207 10.6151
R1020 B.n209 B.n208 10.6151
R1021 B.n209 B.n76 10.6151
R1022 B.n213 B.n76 10.6151
R1023 B.n214 B.n213 10.6151
R1024 B.n215 B.n214 10.6151
R1025 B.n215 B.n74 10.6151
R1026 B.n219 B.n74 10.6151
R1027 B.n220 B.n219 10.6151
R1028 B.n221 B.n220 10.6151
R1029 B.n221 B.n72 10.6151
R1030 B.n225 B.n72 10.6151
R1031 B.n226 B.n225 10.6151
R1032 B.n227 B.n226 10.6151
R1033 B.n148 B.n147 10.6151
R1034 B.n147 B.n102 10.6151
R1035 B.n143 B.n102 10.6151
R1036 B.n143 B.n142 10.6151
R1037 B.n142 B.n141 10.6151
R1038 B.n141 B.n104 10.6151
R1039 B.n137 B.n104 10.6151
R1040 B.n137 B.n136 10.6151
R1041 B.n136 B.n135 10.6151
R1042 B.n135 B.n106 10.6151
R1043 B.n131 B.n106 10.6151
R1044 B.n131 B.n130 10.6151
R1045 B.n130 B.n129 10.6151
R1046 B.n129 B.n108 10.6151
R1047 B.n125 B.n108 10.6151
R1048 B.n125 B.n124 10.6151
R1049 B.n124 B.n123 10.6151
R1050 B.n123 B.n110 10.6151
R1051 B.n119 B.n110 10.6151
R1052 B.n119 B.n118 10.6151
R1053 B.n118 B.n117 10.6151
R1054 B.n117 B.n112 10.6151
R1055 B.n113 B.n112 10.6151
R1056 B.n113 B.n0 10.6151
R1057 B.n419 B.n1 10.6151
R1058 B.n419 B.n418 10.6151
R1059 B.n418 B.n417 10.6151
R1060 B.n417 B.n4 10.6151
R1061 B.n413 B.n4 10.6151
R1062 B.n413 B.n412 10.6151
R1063 B.n412 B.n411 10.6151
R1064 B.n411 B.n6 10.6151
R1065 B.n407 B.n6 10.6151
R1066 B.n407 B.n406 10.6151
R1067 B.n406 B.n405 10.6151
R1068 B.n405 B.n8 10.6151
R1069 B.n401 B.n8 10.6151
R1070 B.n401 B.n400 10.6151
R1071 B.n400 B.n399 10.6151
R1072 B.n399 B.n10 10.6151
R1073 B.n395 B.n10 10.6151
R1074 B.n395 B.n394 10.6151
R1075 B.n394 B.n393 10.6151
R1076 B.n393 B.n12 10.6151
R1077 B.n389 B.n12 10.6151
R1078 B.n389 B.n388 10.6151
R1079 B.n388 B.n387 10.6151
R1080 B.n387 B.n14 10.6151
R1081 B.n353 B.n352 9.36635
R1082 B.n335 B.n34 9.36635
R1083 B.n179 B.n90 9.36635
R1084 B.n197 B.n196 9.36635
R1085 B.n423 B.n0 2.81026
R1086 B.n423 B.n1 2.81026
R1087 B.n352 B.n351 1.24928
R1088 B.n338 B.n34 1.24928
R1089 B.n182 B.n90 1.24928
R1090 B.n196 B.n195 1.24928
C0 VDD1 VN 0.149316f
C1 VDD1 VDD2 0.927715f
C2 VN VDD2 2.94682f
C3 w_n2122_n1996# B 5.31506f
C4 w_n2122_n1996# VP 4.06511f
C5 B VTAIL 1.47142f
C6 VP VTAIL 3.10111f
C7 w_n2122_n1996# VDD1 1.50382f
C8 VDD1 VTAIL 7.77255f
C9 w_n2122_n1996# VN 3.79501f
C10 w_n2122_n1996# VDD2 1.54455f
C11 VN VTAIL 3.08677f
C12 VTAIL VDD2 7.80995f
C13 B VP 1.15478f
C14 VDD1 B 1.17624f
C15 VDD1 VP 3.12717f
C16 B VN 0.711334f
C17 B VDD2 1.2179f
C18 VN VP 4.21865f
C19 VP VDD2 0.336127f
C20 w_n2122_n1996# VTAIL 1.9433f
C21 VDD2 VSUBS 1.066474f
C22 VDD1 VSUBS 0.910633f
C23 VTAIL VSUBS 0.400994f
C24 VN VSUBS 4.327651f
C25 VP VSUBS 1.385643f
C26 B VSUBS 2.238369f
C27 w_n2122_n1996# VSUBS 53.0415f
C28 B.n0 VSUBS 0.004321f
C29 B.n1 VSUBS 0.004321f
C30 B.n2 VSUBS 0.006833f
C31 B.n3 VSUBS 0.006833f
C32 B.n4 VSUBS 0.006833f
C33 B.n5 VSUBS 0.006833f
C34 B.n6 VSUBS 0.006833f
C35 B.n7 VSUBS 0.006833f
C36 B.n8 VSUBS 0.006833f
C37 B.n9 VSUBS 0.006833f
C38 B.n10 VSUBS 0.006833f
C39 B.n11 VSUBS 0.006833f
C40 B.n12 VSUBS 0.006833f
C41 B.n13 VSUBS 0.006833f
C42 B.n14 VSUBS 0.016636f
C43 B.n15 VSUBS 0.006833f
C44 B.n16 VSUBS 0.006833f
C45 B.n17 VSUBS 0.006833f
C46 B.n18 VSUBS 0.006833f
C47 B.n19 VSUBS 0.006833f
C48 B.n20 VSUBS 0.006833f
C49 B.n21 VSUBS 0.006833f
C50 B.n22 VSUBS 0.006833f
C51 B.n23 VSUBS 0.006833f
C52 B.n24 VSUBS 0.006833f
C53 B.n25 VSUBS 0.006833f
C54 B.t11 VSUBS 0.072867f
C55 B.t10 VSUBS 0.081034f
C56 B.t9 VSUBS 0.137375f
C57 B.n26 VSUBS 0.145406f
C58 B.n27 VSUBS 0.12887f
C59 B.n28 VSUBS 0.006833f
C60 B.n29 VSUBS 0.006833f
C61 B.n30 VSUBS 0.006833f
C62 B.n31 VSUBS 0.006833f
C63 B.t2 VSUBS 0.072868f
C64 B.t1 VSUBS 0.081036f
C65 B.t0 VSUBS 0.137375f
C66 B.n32 VSUBS 0.145405f
C67 B.n33 VSUBS 0.128869f
C68 B.n34 VSUBS 0.015831f
C69 B.n35 VSUBS 0.006833f
C70 B.n36 VSUBS 0.006833f
C71 B.n37 VSUBS 0.006833f
C72 B.n38 VSUBS 0.006833f
C73 B.n39 VSUBS 0.006833f
C74 B.n40 VSUBS 0.006833f
C75 B.n41 VSUBS 0.006833f
C76 B.n42 VSUBS 0.006833f
C77 B.n43 VSUBS 0.006833f
C78 B.n44 VSUBS 0.006833f
C79 B.n45 VSUBS 0.016636f
C80 B.n46 VSUBS 0.006833f
C81 B.n47 VSUBS 0.006833f
C82 B.n48 VSUBS 0.006833f
C83 B.n49 VSUBS 0.006833f
C84 B.n50 VSUBS 0.006833f
C85 B.n51 VSUBS 0.006833f
C86 B.n52 VSUBS 0.006833f
C87 B.n53 VSUBS 0.006833f
C88 B.n54 VSUBS 0.006833f
C89 B.n55 VSUBS 0.006833f
C90 B.n56 VSUBS 0.006833f
C91 B.n57 VSUBS 0.006833f
C92 B.n58 VSUBS 0.006833f
C93 B.n59 VSUBS 0.006833f
C94 B.n60 VSUBS 0.006833f
C95 B.n61 VSUBS 0.006833f
C96 B.n62 VSUBS 0.006833f
C97 B.n63 VSUBS 0.006833f
C98 B.n64 VSUBS 0.006833f
C99 B.n65 VSUBS 0.006833f
C100 B.n66 VSUBS 0.006833f
C101 B.n67 VSUBS 0.006833f
C102 B.n68 VSUBS 0.006833f
C103 B.n69 VSUBS 0.006833f
C104 B.n70 VSUBS 0.016636f
C105 B.n71 VSUBS 0.006833f
C106 B.n72 VSUBS 0.006833f
C107 B.n73 VSUBS 0.006833f
C108 B.n74 VSUBS 0.006833f
C109 B.n75 VSUBS 0.006833f
C110 B.n76 VSUBS 0.006833f
C111 B.n77 VSUBS 0.006833f
C112 B.n78 VSUBS 0.006833f
C113 B.n79 VSUBS 0.006833f
C114 B.n80 VSUBS 0.006833f
C115 B.n81 VSUBS 0.006833f
C116 B.t4 VSUBS 0.072868f
C117 B.t5 VSUBS 0.081036f
C118 B.t3 VSUBS 0.137375f
C119 B.n82 VSUBS 0.145405f
C120 B.n83 VSUBS 0.128869f
C121 B.n84 VSUBS 0.006833f
C122 B.n85 VSUBS 0.006833f
C123 B.n86 VSUBS 0.006833f
C124 B.n87 VSUBS 0.006833f
C125 B.t7 VSUBS 0.072867f
C126 B.t8 VSUBS 0.081034f
C127 B.t6 VSUBS 0.137375f
C128 B.n88 VSUBS 0.145406f
C129 B.n89 VSUBS 0.12887f
C130 B.n90 VSUBS 0.015831f
C131 B.n91 VSUBS 0.006833f
C132 B.n92 VSUBS 0.006833f
C133 B.n93 VSUBS 0.006833f
C134 B.n94 VSUBS 0.006833f
C135 B.n95 VSUBS 0.006833f
C136 B.n96 VSUBS 0.006833f
C137 B.n97 VSUBS 0.006833f
C138 B.n98 VSUBS 0.006833f
C139 B.n99 VSUBS 0.006833f
C140 B.n100 VSUBS 0.006833f
C141 B.n101 VSUBS 0.016636f
C142 B.n102 VSUBS 0.006833f
C143 B.n103 VSUBS 0.006833f
C144 B.n104 VSUBS 0.006833f
C145 B.n105 VSUBS 0.006833f
C146 B.n106 VSUBS 0.006833f
C147 B.n107 VSUBS 0.006833f
C148 B.n108 VSUBS 0.006833f
C149 B.n109 VSUBS 0.006833f
C150 B.n110 VSUBS 0.006833f
C151 B.n111 VSUBS 0.006833f
C152 B.n112 VSUBS 0.006833f
C153 B.n113 VSUBS 0.006833f
C154 B.n114 VSUBS 0.006833f
C155 B.n115 VSUBS 0.006833f
C156 B.n116 VSUBS 0.006833f
C157 B.n117 VSUBS 0.006833f
C158 B.n118 VSUBS 0.006833f
C159 B.n119 VSUBS 0.006833f
C160 B.n120 VSUBS 0.006833f
C161 B.n121 VSUBS 0.006833f
C162 B.n122 VSUBS 0.006833f
C163 B.n123 VSUBS 0.006833f
C164 B.n124 VSUBS 0.006833f
C165 B.n125 VSUBS 0.006833f
C166 B.n126 VSUBS 0.006833f
C167 B.n127 VSUBS 0.006833f
C168 B.n128 VSUBS 0.006833f
C169 B.n129 VSUBS 0.006833f
C170 B.n130 VSUBS 0.006833f
C171 B.n131 VSUBS 0.006833f
C172 B.n132 VSUBS 0.006833f
C173 B.n133 VSUBS 0.006833f
C174 B.n134 VSUBS 0.006833f
C175 B.n135 VSUBS 0.006833f
C176 B.n136 VSUBS 0.006833f
C177 B.n137 VSUBS 0.006833f
C178 B.n138 VSUBS 0.006833f
C179 B.n139 VSUBS 0.006833f
C180 B.n140 VSUBS 0.006833f
C181 B.n141 VSUBS 0.006833f
C182 B.n142 VSUBS 0.006833f
C183 B.n143 VSUBS 0.006833f
C184 B.n144 VSUBS 0.006833f
C185 B.n145 VSUBS 0.006833f
C186 B.n146 VSUBS 0.006833f
C187 B.n147 VSUBS 0.006833f
C188 B.n148 VSUBS 0.016636f
C189 B.n149 VSUBS 0.017126f
C190 B.n150 VSUBS 0.017126f
C191 B.n151 VSUBS 0.006833f
C192 B.n152 VSUBS 0.006833f
C193 B.n153 VSUBS 0.006833f
C194 B.n154 VSUBS 0.006833f
C195 B.n155 VSUBS 0.006833f
C196 B.n156 VSUBS 0.006833f
C197 B.n157 VSUBS 0.006833f
C198 B.n158 VSUBS 0.006833f
C199 B.n159 VSUBS 0.006833f
C200 B.n160 VSUBS 0.006833f
C201 B.n161 VSUBS 0.006833f
C202 B.n162 VSUBS 0.006833f
C203 B.n163 VSUBS 0.006833f
C204 B.n164 VSUBS 0.006833f
C205 B.n165 VSUBS 0.006833f
C206 B.n166 VSUBS 0.006833f
C207 B.n167 VSUBS 0.006833f
C208 B.n168 VSUBS 0.006833f
C209 B.n169 VSUBS 0.006833f
C210 B.n170 VSUBS 0.006833f
C211 B.n171 VSUBS 0.006833f
C212 B.n172 VSUBS 0.006833f
C213 B.n173 VSUBS 0.006833f
C214 B.n174 VSUBS 0.006833f
C215 B.n175 VSUBS 0.006833f
C216 B.n176 VSUBS 0.006833f
C217 B.n177 VSUBS 0.006833f
C218 B.n178 VSUBS 0.006833f
C219 B.n179 VSUBS 0.006431f
C220 B.n180 VSUBS 0.006833f
C221 B.n181 VSUBS 0.006833f
C222 B.n182 VSUBS 0.003818f
C223 B.n183 VSUBS 0.006833f
C224 B.n184 VSUBS 0.006833f
C225 B.n185 VSUBS 0.006833f
C226 B.n186 VSUBS 0.006833f
C227 B.n187 VSUBS 0.006833f
C228 B.n188 VSUBS 0.006833f
C229 B.n189 VSUBS 0.006833f
C230 B.n190 VSUBS 0.006833f
C231 B.n191 VSUBS 0.006833f
C232 B.n192 VSUBS 0.006833f
C233 B.n193 VSUBS 0.006833f
C234 B.n194 VSUBS 0.006833f
C235 B.n195 VSUBS 0.003818f
C236 B.n196 VSUBS 0.015831f
C237 B.n197 VSUBS 0.006431f
C238 B.n198 VSUBS 0.006833f
C239 B.n199 VSUBS 0.006833f
C240 B.n200 VSUBS 0.006833f
C241 B.n201 VSUBS 0.006833f
C242 B.n202 VSUBS 0.006833f
C243 B.n203 VSUBS 0.006833f
C244 B.n204 VSUBS 0.006833f
C245 B.n205 VSUBS 0.006833f
C246 B.n206 VSUBS 0.006833f
C247 B.n207 VSUBS 0.006833f
C248 B.n208 VSUBS 0.006833f
C249 B.n209 VSUBS 0.006833f
C250 B.n210 VSUBS 0.006833f
C251 B.n211 VSUBS 0.006833f
C252 B.n212 VSUBS 0.006833f
C253 B.n213 VSUBS 0.006833f
C254 B.n214 VSUBS 0.006833f
C255 B.n215 VSUBS 0.006833f
C256 B.n216 VSUBS 0.006833f
C257 B.n217 VSUBS 0.006833f
C258 B.n218 VSUBS 0.006833f
C259 B.n219 VSUBS 0.006833f
C260 B.n220 VSUBS 0.006833f
C261 B.n221 VSUBS 0.006833f
C262 B.n222 VSUBS 0.006833f
C263 B.n223 VSUBS 0.006833f
C264 B.n224 VSUBS 0.006833f
C265 B.n225 VSUBS 0.006833f
C266 B.n226 VSUBS 0.006833f
C267 B.n227 VSUBS 0.017126f
C268 B.n228 VSUBS 0.017126f
C269 B.n229 VSUBS 0.016636f
C270 B.n230 VSUBS 0.006833f
C271 B.n231 VSUBS 0.006833f
C272 B.n232 VSUBS 0.006833f
C273 B.n233 VSUBS 0.006833f
C274 B.n234 VSUBS 0.006833f
C275 B.n235 VSUBS 0.006833f
C276 B.n236 VSUBS 0.006833f
C277 B.n237 VSUBS 0.006833f
C278 B.n238 VSUBS 0.006833f
C279 B.n239 VSUBS 0.006833f
C280 B.n240 VSUBS 0.006833f
C281 B.n241 VSUBS 0.006833f
C282 B.n242 VSUBS 0.006833f
C283 B.n243 VSUBS 0.006833f
C284 B.n244 VSUBS 0.006833f
C285 B.n245 VSUBS 0.006833f
C286 B.n246 VSUBS 0.006833f
C287 B.n247 VSUBS 0.006833f
C288 B.n248 VSUBS 0.006833f
C289 B.n249 VSUBS 0.006833f
C290 B.n250 VSUBS 0.006833f
C291 B.n251 VSUBS 0.006833f
C292 B.n252 VSUBS 0.006833f
C293 B.n253 VSUBS 0.006833f
C294 B.n254 VSUBS 0.006833f
C295 B.n255 VSUBS 0.006833f
C296 B.n256 VSUBS 0.006833f
C297 B.n257 VSUBS 0.006833f
C298 B.n258 VSUBS 0.006833f
C299 B.n259 VSUBS 0.006833f
C300 B.n260 VSUBS 0.006833f
C301 B.n261 VSUBS 0.006833f
C302 B.n262 VSUBS 0.006833f
C303 B.n263 VSUBS 0.006833f
C304 B.n264 VSUBS 0.006833f
C305 B.n265 VSUBS 0.006833f
C306 B.n266 VSUBS 0.006833f
C307 B.n267 VSUBS 0.006833f
C308 B.n268 VSUBS 0.006833f
C309 B.n269 VSUBS 0.006833f
C310 B.n270 VSUBS 0.006833f
C311 B.n271 VSUBS 0.006833f
C312 B.n272 VSUBS 0.006833f
C313 B.n273 VSUBS 0.006833f
C314 B.n274 VSUBS 0.006833f
C315 B.n275 VSUBS 0.006833f
C316 B.n276 VSUBS 0.006833f
C317 B.n277 VSUBS 0.006833f
C318 B.n278 VSUBS 0.006833f
C319 B.n279 VSUBS 0.006833f
C320 B.n280 VSUBS 0.006833f
C321 B.n281 VSUBS 0.006833f
C322 B.n282 VSUBS 0.006833f
C323 B.n283 VSUBS 0.006833f
C324 B.n284 VSUBS 0.006833f
C325 B.n285 VSUBS 0.006833f
C326 B.n286 VSUBS 0.006833f
C327 B.n287 VSUBS 0.006833f
C328 B.n288 VSUBS 0.006833f
C329 B.n289 VSUBS 0.006833f
C330 B.n290 VSUBS 0.006833f
C331 B.n291 VSUBS 0.006833f
C332 B.n292 VSUBS 0.006833f
C333 B.n293 VSUBS 0.006833f
C334 B.n294 VSUBS 0.006833f
C335 B.n295 VSUBS 0.006833f
C336 B.n296 VSUBS 0.006833f
C337 B.n297 VSUBS 0.006833f
C338 B.n298 VSUBS 0.006833f
C339 B.n299 VSUBS 0.006833f
C340 B.n300 VSUBS 0.006833f
C341 B.n301 VSUBS 0.006833f
C342 B.n302 VSUBS 0.006833f
C343 B.n303 VSUBS 0.006833f
C344 B.n304 VSUBS 0.01738f
C345 B.n305 VSUBS 0.016382f
C346 B.n306 VSUBS 0.017126f
C347 B.n307 VSUBS 0.006833f
C348 B.n308 VSUBS 0.006833f
C349 B.n309 VSUBS 0.006833f
C350 B.n310 VSUBS 0.006833f
C351 B.n311 VSUBS 0.006833f
C352 B.n312 VSUBS 0.006833f
C353 B.n313 VSUBS 0.006833f
C354 B.n314 VSUBS 0.006833f
C355 B.n315 VSUBS 0.006833f
C356 B.n316 VSUBS 0.006833f
C357 B.n317 VSUBS 0.006833f
C358 B.n318 VSUBS 0.006833f
C359 B.n319 VSUBS 0.006833f
C360 B.n320 VSUBS 0.006833f
C361 B.n321 VSUBS 0.006833f
C362 B.n322 VSUBS 0.006833f
C363 B.n323 VSUBS 0.006833f
C364 B.n324 VSUBS 0.006833f
C365 B.n325 VSUBS 0.006833f
C366 B.n326 VSUBS 0.006833f
C367 B.n327 VSUBS 0.006833f
C368 B.n328 VSUBS 0.006833f
C369 B.n329 VSUBS 0.006833f
C370 B.n330 VSUBS 0.006833f
C371 B.n331 VSUBS 0.006833f
C372 B.n332 VSUBS 0.006833f
C373 B.n333 VSUBS 0.006833f
C374 B.n334 VSUBS 0.006833f
C375 B.n335 VSUBS 0.006431f
C376 B.n336 VSUBS 0.006833f
C377 B.n337 VSUBS 0.006833f
C378 B.n338 VSUBS 0.003818f
C379 B.n339 VSUBS 0.006833f
C380 B.n340 VSUBS 0.006833f
C381 B.n341 VSUBS 0.006833f
C382 B.n342 VSUBS 0.006833f
C383 B.n343 VSUBS 0.006833f
C384 B.n344 VSUBS 0.006833f
C385 B.n345 VSUBS 0.006833f
C386 B.n346 VSUBS 0.006833f
C387 B.n347 VSUBS 0.006833f
C388 B.n348 VSUBS 0.006833f
C389 B.n349 VSUBS 0.006833f
C390 B.n350 VSUBS 0.006833f
C391 B.n351 VSUBS 0.003818f
C392 B.n352 VSUBS 0.015831f
C393 B.n353 VSUBS 0.006431f
C394 B.n354 VSUBS 0.006833f
C395 B.n355 VSUBS 0.006833f
C396 B.n356 VSUBS 0.006833f
C397 B.n357 VSUBS 0.006833f
C398 B.n358 VSUBS 0.006833f
C399 B.n359 VSUBS 0.006833f
C400 B.n360 VSUBS 0.006833f
C401 B.n361 VSUBS 0.006833f
C402 B.n362 VSUBS 0.006833f
C403 B.n363 VSUBS 0.006833f
C404 B.n364 VSUBS 0.006833f
C405 B.n365 VSUBS 0.006833f
C406 B.n366 VSUBS 0.006833f
C407 B.n367 VSUBS 0.006833f
C408 B.n368 VSUBS 0.006833f
C409 B.n369 VSUBS 0.006833f
C410 B.n370 VSUBS 0.006833f
C411 B.n371 VSUBS 0.006833f
C412 B.n372 VSUBS 0.006833f
C413 B.n373 VSUBS 0.006833f
C414 B.n374 VSUBS 0.006833f
C415 B.n375 VSUBS 0.006833f
C416 B.n376 VSUBS 0.006833f
C417 B.n377 VSUBS 0.006833f
C418 B.n378 VSUBS 0.006833f
C419 B.n379 VSUBS 0.006833f
C420 B.n380 VSUBS 0.006833f
C421 B.n381 VSUBS 0.006833f
C422 B.n382 VSUBS 0.006833f
C423 B.n383 VSUBS 0.017126f
C424 B.n384 VSUBS 0.017126f
C425 B.n385 VSUBS 0.016636f
C426 B.n386 VSUBS 0.006833f
C427 B.n387 VSUBS 0.006833f
C428 B.n388 VSUBS 0.006833f
C429 B.n389 VSUBS 0.006833f
C430 B.n390 VSUBS 0.006833f
C431 B.n391 VSUBS 0.006833f
C432 B.n392 VSUBS 0.006833f
C433 B.n393 VSUBS 0.006833f
C434 B.n394 VSUBS 0.006833f
C435 B.n395 VSUBS 0.006833f
C436 B.n396 VSUBS 0.006833f
C437 B.n397 VSUBS 0.006833f
C438 B.n398 VSUBS 0.006833f
C439 B.n399 VSUBS 0.006833f
C440 B.n400 VSUBS 0.006833f
C441 B.n401 VSUBS 0.006833f
C442 B.n402 VSUBS 0.006833f
C443 B.n403 VSUBS 0.006833f
C444 B.n404 VSUBS 0.006833f
C445 B.n405 VSUBS 0.006833f
C446 B.n406 VSUBS 0.006833f
C447 B.n407 VSUBS 0.006833f
C448 B.n408 VSUBS 0.006833f
C449 B.n409 VSUBS 0.006833f
C450 B.n410 VSUBS 0.006833f
C451 B.n411 VSUBS 0.006833f
C452 B.n412 VSUBS 0.006833f
C453 B.n413 VSUBS 0.006833f
C454 B.n414 VSUBS 0.006833f
C455 B.n415 VSUBS 0.006833f
C456 B.n416 VSUBS 0.006833f
C457 B.n417 VSUBS 0.006833f
C458 B.n418 VSUBS 0.006833f
C459 B.n419 VSUBS 0.006833f
C460 B.n420 VSUBS 0.006833f
C461 B.n421 VSUBS 0.006833f
C462 B.n422 VSUBS 0.006833f
C463 B.n423 VSUBS 0.015472f
C464 VDD1.n0 VSUBS 0.014141f
C465 VDD1.n1 VSUBS 0.031831f
C466 VDD1.n2 VSUBS 0.014259f
C467 VDD1.n3 VSUBS 0.025061f
C468 VDD1.n4 VSUBS 0.013467f
C469 VDD1.n5 VSUBS 0.031831f
C470 VDD1.n6 VSUBS 0.014259f
C471 VDD1.n7 VSUBS 0.120276f
C472 VDD1.t3 VSUBS 0.068824f
C473 VDD1.n8 VSUBS 0.023873f
C474 VDD1.n9 VSUBS 0.023915f
C475 VDD1.n10 VSUBS 0.013467f
C476 VDD1.n11 VSUBS 0.476623f
C477 VDD1.n12 VSUBS 0.025061f
C478 VDD1.n13 VSUBS 0.013467f
C479 VDD1.n14 VSUBS 0.014259f
C480 VDD1.n15 VSUBS 0.031831f
C481 VDD1.n16 VSUBS 0.031831f
C482 VDD1.n17 VSUBS 0.014259f
C483 VDD1.n18 VSUBS 0.013467f
C484 VDD1.n19 VSUBS 0.025061f
C485 VDD1.n20 VSUBS 0.06546f
C486 VDD1.n21 VSUBS 0.013467f
C487 VDD1.n22 VSUBS 0.014259f
C488 VDD1.n23 VSUBS 0.070188f
C489 VDD1.n24 VSUBS 0.066881f
C490 VDD1.t1 VSUBS 0.101793f
C491 VDD1.t4 VSUBS 0.101793f
C492 VDD1.n25 VSUBS 0.661944f
C493 VDD1.n26 VSUBS 0.574208f
C494 VDD1.n27 VSUBS 0.014141f
C495 VDD1.n28 VSUBS 0.031831f
C496 VDD1.n29 VSUBS 0.014259f
C497 VDD1.n30 VSUBS 0.025061f
C498 VDD1.n31 VSUBS 0.013467f
C499 VDD1.n32 VSUBS 0.031831f
C500 VDD1.n33 VSUBS 0.014259f
C501 VDD1.n34 VSUBS 0.120276f
C502 VDD1.t0 VSUBS 0.068824f
C503 VDD1.n35 VSUBS 0.023873f
C504 VDD1.n36 VSUBS 0.023915f
C505 VDD1.n37 VSUBS 0.013467f
C506 VDD1.n38 VSUBS 0.476623f
C507 VDD1.n39 VSUBS 0.025061f
C508 VDD1.n40 VSUBS 0.013467f
C509 VDD1.n41 VSUBS 0.014259f
C510 VDD1.n42 VSUBS 0.031831f
C511 VDD1.n43 VSUBS 0.031831f
C512 VDD1.n44 VSUBS 0.014259f
C513 VDD1.n45 VSUBS 0.013467f
C514 VDD1.n46 VSUBS 0.025061f
C515 VDD1.n47 VSUBS 0.06546f
C516 VDD1.n48 VSUBS 0.013467f
C517 VDD1.n49 VSUBS 0.014259f
C518 VDD1.n50 VSUBS 0.070188f
C519 VDD1.n51 VSUBS 0.066881f
C520 VDD1.t7 VSUBS 0.101793f
C521 VDD1.t9 VSUBS 0.101793f
C522 VDD1.n52 VSUBS 0.661941f
C523 VDD1.n53 VSUBS 0.568877f
C524 VDD1.t2 VSUBS 0.101793f
C525 VDD1.t8 VSUBS 0.101793f
C526 VDD1.n54 VSUBS 0.664697f
C527 VDD1.n55 VSUBS 1.70024f
C528 VDD1.t5 VSUBS 0.101793f
C529 VDD1.t6 VSUBS 0.101793f
C530 VDD1.n56 VSUBS 0.66194f
C531 VDD1.n57 VSUBS 1.98235f
C532 VP.n0 VSUBS 0.107619f
C533 VP.t2 VSUBS 0.610306f
C534 VP.n1 VSUBS 0.311852f
C535 VP.n2 VSUBS 0.107619f
C536 VP.t3 VSUBS 0.610306f
C537 VP.t4 VSUBS 0.610306f
C538 VP.t5 VSUBS 0.610306f
C539 VP.n3 VSUBS 0.339815f
C540 VP.t8 VSUBS 0.610306f
C541 VP.t6 VSUBS 0.638213f
C542 VP.n4 VSUBS 0.27125f
C543 VP.n5 VSUBS 0.311852f
C544 VP.n6 VSUBS 0.311852f
C545 VP.n7 VSUBS 0.311852f
C546 VP.n8 VSUBS 0.29719f
C547 VP.n9 VSUBS 2.18789f
C548 VP.t9 VSUBS 0.610306f
C549 VP.n10 VSUBS 0.29719f
C550 VP.n11 VSUBS 2.25038f
C551 VP.n12 VSUBS 0.107619f
C552 VP.n13 VSUBS 0.129224f
C553 VP.t0 VSUBS 0.610306f
C554 VP.n14 VSUBS 0.311852f
C555 VP.t7 VSUBS 0.610306f
C556 VP.n15 VSUBS 0.311852f
C557 VP.t1 VSUBS 0.610306f
C558 VP.n16 VSUBS 0.29719f
C559 VP.n17 VSUBS 0.071676f
C560 VDD2.n0 VSUBS 0.014f
C561 VDD2.n1 VSUBS 0.031514f
C562 VDD2.n2 VSUBS 0.014117f
C563 VDD2.n3 VSUBS 0.024812f
C564 VDD2.n4 VSUBS 0.013333f
C565 VDD2.n5 VSUBS 0.031514f
C566 VDD2.n6 VSUBS 0.014117f
C567 VDD2.n7 VSUBS 0.119081f
C568 VDD2.t9 VSUBS 0.06814f
C569 VDD2.n8 VSUBS 0.023636f
C570 VDD2.n9 VSUBS 0.023678f
C571 VDD2.n10 VSUBS 0.013333f
C572 VDD2.n11 VSUBS 0.471885f
C573 VDD2.n12 VSUBS 0.024812f
C574 VDD2.n13 VSUBS 0.013333f
C575 VDD2.n14 VSUBS 0.014117f
C576 VDD2.n15 VSUBS 0.031514f
C577 VDD2.n16 VSUBS 0.031514f
C578 VDD2.n17 VSUBS 0.014117f
C579 VDD2.n18 VSUBS 0.013333f
C580 VDD2.n19 VSUBS 0.024812f
C581 VDD2.n20 VSUBS 0.064809f
C582 VDD2.n21 VSUBS 0.013333f
C583 VDD2.n22 VSUBS 0.014117f
C584 VDD2.n23 VSUBS 0.06949f
C585 VDD2.n24 VSUBS 0.066216f
C586 VDD2.t2 VSUBS 0.100781f
C587 VDD2.t0 VSUBS 0.100781f
C588 VDD2.n25 VSUBS 0.655361f
C589 VDD2.n26 VSUBS 0.563221f
C590 VDD2.t8 VSUBS 0.100781f
C591 VDD2.t1 VSUBS 0.100781f
C592 VDD2.n27 VSUBS 0.65809f
C593 VDD2.n28 VSUBS 1.61123f
C594 VDD2.n29 VSUBS 0.014f
C595 VDD2.n30 VSUBS 0.031514f
C596 VDD2.n31 VSUBS 0.014117f
C597 VDD2.n32 VSUBS 0.024812f
C598 VDD2.n33 VSUBS 0.013333f
C599 VDD2.n34 VSUBS 0.031514f
C600 VDD2.n35 VSUBS 0.014117f
C601 VDD2.n36 VSUBS 0.119081f
C602 VDD2.t4 VSUBS 0.06814f
C603 VDD2.n37 VSUBS 0.023636f
C604 VDD2.n38 VSUBS 0.023678f
C605 VDD2.n39 VSUBS 0.013333f
C606 VDD2.n40 VSUBS 0.471885f
C607 VDD2.n41 VSUBS 0.024812f
C608 VDD2.n42 VSUBS 0.013333f
C609 VDD2.n43 VSUBS 0.014117f
C610 VDD2.n44 VSUBS 0.031514f
C611 VDD2.n45 VSUBS 0.031514f
C612 VDD2.n46 VSUBS 0.014117f
C613 VDD2.n47 VSUBS 0.013333f
C614 VDD2.n48 VSUBS 0.024812f
C615 VDD2.n49 VSUBS 0.064809f
C616 VDD2.n50 VSUBS 0.013333f
C617 VDD2.n51 VSUBS 0.014117f
C618 VDD2.n52 VSUBS 0.06949f
C619 VDD2.n53 VSUBS 0.064367f
C620 VDD2.n54 VSUBS 1.57152f
C621 VDD2.t3 VSUBS 0.100781f
C622 VDD2.t5 VSUBS 0.100781f
C623 VDD2.n55 VSUBS 0.655363f
C624 VDD2.n56 VSUBS 0.454078f
C625 VDD2.t6 VSUBS 0.100781f
C626 VDD2.t7 VSUBS 0.100781f
C627 VDD2.n57 VSUBS 0.658068f
C628 VTAIL.t15 VSUBS 0.115174f
C629 VTAIL.t12 VSUBS 0.115174f
C630 VTAIL.n0 VSUBS 0.6669f
C631 VTAIL.n1 VSUBS 0.605376f
C632 VTAIL.n2 VSUBS 0.016f
C633 VTAIL.n3 VSUBS 0.036015f
C634 VTAIL.n4 VSUBS 0.016133f
C635 VTAIL.n5 VSUBS 0.028356f
C636 VTAIL.n6 VSUBS 0.015237f
C637 VTAIL.n7 VSUBS 0.036015f
C638 VTAIL.n8 VSUBS 0.016133f
C639 VTAIL.n9 VSUBS 0.136087f
C640 VTAIL.t8 VSUBS 0.077871f
C641 VTAIL.n10 VSUBS 0.027011f
C642 VTAIL.n11 VSUBS 0.027059f
C643 VTAIL.n12 VSUBS 0.015237f
C644 VTAIL.n13 VSUBS 0.539278f
C645 VTAIL.n14 VSUBS 0.028356f
C646 VTAIL.n15 VSUBS 0.015237f
C647 VTAIL.n16 VSUBS 0.016133f
C648 VTAIL.n17 VSUBS 0.036015f
C649 VTAIL.n18 VSUBS 0.036015f
C650 VTAIL.n19 VSUBS 0.016133f
C651 VTAIL.n20 VSUBS 0.015237f
C652 VTAIL.n21 VSUBS 0.028356f
C653 VTAIL.n22 VSUBS 0.074065f
C654 VTAIL.n23 VSUBS 0.015237f
C655 VTAIL.n24 VSUBS 0.016133f
C656 VTAIL.n25 VSUBS 0.079415f
C657 VTAIL.n26 VSUBS 0.054014f
C658 VTAIL.n27 VSUBS 0.183196f
C659 VTAIL.t3 VSUBS 0.115174f
C660 VTAIL.t0 VSUBS 0.115174f
C661 VTAIL.n28 VSUBS 0.6669f
C662 VTAIL.n29 VSUBS 0.613844f
C663 VTAIL.t2 VSUBS 0.115174f
C664 VTAIL.t5 VSUBS 0.115174f
C665 VTAIL.n30 VSUBS 0.6669f
C666 VTAIL.n31 VSUBS 1.47949f
C667 VTAIL.t19 VSUBS 0.115174f
C668 VTAIL.t17 VSUBS 0.115174f
C669 VTAIL.n32 VSUBS 0.666903f
C670 VTAIL.n33 VSUBS 1.47949f
C671 VTAIL.t16 VSUBS 0.115174f
C672 VTAIL.t18 VSUBS 0.115174f
C673 VTAIL.n34 VSUBS 0.666903f
C674 VTAIL.n35 VSUBS 0.61384f
C675 VTAIL.n36 VSUBS 0.016f
C676 VTAIL.n37 VSUBS 0.036015f
C677 VTAIL.n38 VSUBS 0.016133f
C678 VTAIL.n39 VSUBS 0.028356f
C679 VTAIL.n40 VSUBS 0.015237f
C680 VTAIL.n41 VSUBS 0.036015f
C681 VTAIL.n42 VSUBS 0.016133f
C682 VTAIL.n43 VSUBS 0.136087f
C683 VTAIL.t13 VSUBS 0.077871f
C684 VTAIL.n44 VSUBS 0.027011f
C685 VTAIL.n45 VSUBS 0.027059f
C686 VTAIL.n46 VSUBS 0.015237f
C687 VTAIL.n47 VSUBS 0.539278f
C688 VTAIL.n48 VSUBS 0.028356f
C689 VTAIL.n49 VSUBS 0.015237f
C690 VTAIL.n50 VSUBS 0.016133f
C691 VTAIL.n51 VSUBS 0.036015f
C692 VTAIL.n52 VSUBS 0.036015f
C693 VTAIL.n53 VSUBS 0.016133f
C694 VTAIL.n54 VSUBS 0.015237f
C695 VTAIL.n55 VSUBS 0.028356f
C696 VTAIL.n56 VSUBS 0.074065f
C697 VTAIL.n57 VSUBS 0.015237f
C698 VTAIL.n58 VSUBS 0.016133f
C699 VTAIL.n59 VSUBS 0.079415f
C700 VTAIL.n60 VSUBS 0.054014f
C701 VTAIL.n61 VSUBS 0.183196f
C702 VTAIL.t7 VSUBS 0.115174f
C703 VTAIL.t1 VSUBS 0.115174f
C704 VTAIL.n62 VSUBS 0.666903f
C705 VTAIL.n63 VSUBS 0.61896f
C706 VTAIL.t9 VSUBS 0.115174f
C707 VTAIL.t4 VSUBS 0.115174f
C708 VTAIL.n64 VSUBS 0.666903f
C709 VTAIL.n65 VSUBS 0.61384f
C710 VTAIL.n66 VSUBS 0.016f
C711 VTAIL.n67 VSUBS 0.036015f
C712 VTAIL.n68 VSUBS 0.016133f
C713 VTAIL.n69 VSUBS 0.028356f
C714 VTAIL.n70 VSUBS 0.015237f
C715 VTAIL.n71 VSUBS 0.036015f
C716 VTAIL.n72 VSUBS 0.016133f
C717 VTAIL.n73 VSUBS 0.136087f
C718 VTAIL.t6 VSUBS 0.077871f
C719 VTAIL.n74 VSUBS 0.027011f
C720 VTAIL.n75 VSUBS 0.027059f
C721 VTAIL.n76 VSUBS 0.015237f
C722 VTAIL.n77 VSUBS 0.539278f
C723 VTAIL.n78 VSUBS 0.028356f
C724 VTAIL.n79 VSUBS 0.015237f
C725 VTAIL.n80 VSUBS 0.016133f
C726 VTAIL.n81 VSUBS 0.036015f
C727 VTAIL.n82 VSUBS 0.036015f
C728 VTAIL.n83 VSUBS 0.016133f
C729 VTAIL.n84 VSUBS 0.015237f
C730 VTAIL.n85 VSUBS 0.028356f
C731 VTAIL.n86 VSUBS 0.074065f
C732 VTAIL.n87 VSUBS 0.015237f
C733 VTAIL.n88 VSUBS 0.016133f
C734 VTAIL.n89 VSUBS 0.079415f
C735 VTAIL.n90 VSUBS 0.054014f
C736 VTAIL.n91 VSUBS 0.968109f
C737 VTAIL.n92 VSUBS 0.016f
C738 VTAIL.n93 VSUBS 0.036015f
C739 VTAIL.n94 VSUBS 0.016133f
C740 VTAIL.n95 VSUBS 0.028356f
C741 VTAIL.n96 VSUBS 0.015237f
C742 VTAIL.n97 VSUBS 0.036015f
C743 VTAIL.n98 VSUBS 0.016133f
C744 VTAIL.n99 VSUBS 0.136087f
C745 VTAIL.t14 VSUBS 0.077871f
C746 VTAIL.n100 VSUBS 0.027011f
C747 VTAIL.n101 VSUBS 0.027059f
C748 VTAIL.n102 VSUBS 0.015237f
C749 VTAIL.n103 VSUBS 0.539278f
C750 VTAIL.n104 VSUBS 0.028356f
C751 VTAIL.n105 VSUBS 0.015237f
C752 VTAIL.n106 VSUBS 0.016133f
C753 VTAIL.n107 VSUBS 0.036015f
C754 VTAIL.n108 VSUBS 0.036015f
C755 VTAIL.n109 VSUBS 0.016133f
C756 VTAIL.n110 VSUBS 0.015237f
C757 VTAIL.n111 VSUBS 0.028356f
C758 VTAIL.n112 VSUBS 0.074065f
C759 VTAIL.n113 VSUBS 0.015237f
C760 VTAIL.n114 VSUBS 0.016133f
C761 VTAIL.n115 VSUBS 0.079415f
C762 VTAIL.n116 VSUBS 0.054014f
C763 VTAIL.n117 VSUBS 0.968109f
C764 VTAIL.t11 VSUBS 0.115174f
C765 VTAIL.t10 VSUBS 0.115174f
C766 VTAIL.n118 VSUBS 0.6669f
C767 VTAIL.n119 VSUBS 0.551816f
C768 VN.n0 VSUBS 0.103261f
C769 VN.t7 VSUBS 0.585593f
C770 VN.n1 VSUBS 0.299224f
C771 VN.t0 VSUBS 0.61237f
C772 VN.n2 VSUBS 0.260266f
C773 VN.n3 VSUBS 0.326055f
C774 VN.t9 VSUBS 0.585593f
C775 VN.n4 VSUBS 0.299224f
C776 VN.t1 VSUBS 0.585593f
C777 VN.n5 VSUBS 0.299224f
C778 VN.t8 VSUBS 0.585593f
C779 VN.n6 VSUBS 0.285156f
C780 VN.n7 VSUBS 0.068774f
C781 VN.n8 VSUBS 0.103261f
C782 VN.t3 VSUBS 0.585593f
C783 VN.n9 VSUBS 0.299224f
C784 VN.t4 VSUBS 0.585593f
C785 VN.t2 VSUBS 0.61237f
C786 VN.n10 VSUBS 0.260266f
C787 VN.n11 VSUBS 0.326055f
C788 VN.n12 VSUBS 0.299224f
C789 VN.t6 VSUBS 0.585593f
C790 VN.n13 VSUBS 0.299224f
C791 VN.t5 VSUBS 0.585593f
C792 VN.n14 VSUBS 0.285156f
C793 VN.n15 VSUBS 2.14031f
.ends

