* NGSPICE file created from diff_pair_sample_1077.ext - technology: sky130A

.subckt diff_pair_sample_1077 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 w_n2090_n3756# sky130_fd_pr__pfet_01v8 ad=5.4366 pd=28.66 as=5.4366 ps=28.66 w=13.94 l=2.47
X1 B.t11 B.t9 B.t10 w_n2090_n3756# sky130_fd_pr__pfet_01v8 ad=5.4366 pd=28.66 as=0 ps=0 w=13.94 l=2.47
X2 B.t8 B.t6 B.t7 w_n2090_n3756# sky130_fd_pr__pfet_01v8 ad=5.4366 pd=28.66 as=0 ps=0 w=13.94 l=2.47
X3 VDD2.t1 VN.t0 VTAIL.t1 w_n2090_n3756# sky130_fd_pr__pfet_01v8 ad=5.4366 pd=28.66 as=5.4366 ps=28.66 w=13.94 l=2.47
X4 B.t5 B.t3 B.t4 w_n2090_n3756# sky130_fd_pr__pfet_01v8 ad=5.4366 pd=28.66 as=0 ps=0 w=13.94 l=2.47
X5 B.t2 B.t0 B.t1 w_n2090_n3756# sky130_fd_pr__pfet_01v8 ad=5.4366 pd=28.66 as=0 ps=0 w=13.94 l=2.47
X6 VDD1.t0 VP.t1 VTAIL.t2 w_n2090_n3756# sky130_fd_pr__pfet_01v8 ad=5.4366 pd=28.66 as=5.4366 ps=28.66 w=13.94 l=2.47
X7 VDD2.t0 VN.t1 VTAIL.t0 w_n2090_n3756# sky130_fd_pr__pfet_01v8 ad=5.4366 pd=28.66 as=5.4366 ps=28.66 w=13.94 l=2.47
R0 VP.n0 VP.t1 231.011
R1 VP.n0 VP.t0 185.23
R2 VP VP.n0 0.336784
R3 VTAIL.n2 VTAIL.t2 57.988
R4 VTAIL.n1 VTAIL.t1 57.988
R5 VTAIL.n3 VTAIL.t0 57.9878
R6 VTAIL.n0 VTAIL.t3 57.9878
R7 VTAIL.n1 VTAIL.n0 29.2117
R8 VTAIL.n3 VTAIL.n2 26.7979
R9 VTAIL.n2 VTAIL.n1 1.67722
R10 VTAIL VTAIL.n0 1.13197
R11 VTAIL VTAIL.n3 0.545759
R12 VDD1 VDD1.t1 116.299
R13 VDD1 VDD1.t0 75.3285
R14 B.n355 B.n96 585
R15 B.n354 B.n353 585
R16 B.n352 B.n97 585
R17 B.n351 B.n350 585
R18 B.n349 B.n98 585
R19 B.n348 B.n347 585
R20 B.n346 B.n99 585
R21 B.n345 B.n344 585
R22 B.n343 B.n100 585
R23 B.n342 B.n341 585
R24 B.n340 B.n101 585
R25 B.n339 B.n338 585
R26 B.n337 B.n102 585
R27 B.n336 B.n335 585
R28 B.n334 B.n103 585
R29 B.n333 B.n332 585
R30 B.n331 B.n104 585
R31 B.n330 B.n329 585
R32 B.n328 B.n105 585
R33 B.n327 B.n326 585
R34 B.n325 B.n106 585
R35 B.n324 B.n323 585
R36 B.n322 B.n107 585
R37 B.n321 B.n320 585
R38 B.n319 B.n108 585
R39 B.n318 B.n317 585
R40 B.n316 B.n109 585
R41 B.n315 B.n314 585
R42 B.n313 B.n110 585
R43 B.n312 B.n311 585
R44 B.n310 B.n111 585
R45 B.n309 B.n308 585
R46 B.n307 B.n112 585
R47 B.n306 B.n305 585
R48 B.n304 B.n113 585
R49 B.n303 B.n302 585
R50 B.n301 B.n114 585
R51 B.n300 B.n299 585
R52 B.n298 B.n115 585
R53 B.n297 B.n296 585
R54 B.n295 B.n116 585
R55 B.n294 B.n293 585
R56 B.n292 B.n117 585
R57 B.n291 B.n290 585
R58 B.n289 B.n118 585
R59 B.n288 B.n287 585
R60 B.n286 B.n119 585
R61 B.n285 B.n284 585
R62 B.n280 B.n120 585
R63 B.n279 B.n278 585
R64 B.n277 B.n121 585
R65 B.n276 B.n275 585
R66 B.n274 B.n122 585
R67 B.n273 B.n272 585
R68 B.n271 B.n123 585
R69 B.n270 B.n269 585
R70 B.n268 B.n124 585
R71 B.n266 B.n265 585
R72 B.n264 B.n127 585
R73 B.n263 B.n262 585
R74 B.n261 B.n128 585
R75 B.n260 B.n259 585
R76 B.n258 B.n129 585
R77 B.n257 B.n256 585
R78 B.n255 B.n130 585
R79 B.n254 B.n253 585
R80 B.n252 B.n131 585
R81 B.n251 B.n250 585
R82 B.n249 B.n132 585
R83 B.n248 B.n247 585
R84 B.n246 B.n133 585
R85 B.n245 B.n244 585
R86 B.n243 B.n134 585
R87 B.n242 B.n241 585
R88 B.n240 B.n135 585
R89 B.n239 B.n238 585
R90 B.n237 B.n136 585
R91 B.n236 B.n235 585
R92 B.n234 B.n137 585
R93 B.n233 B.n232 585
R94 B.n231 B.n138 585
R95 B.n230 B.n229 585
R96 B.n228 B.n139 585
R97 B.n227 B.n226 585
R98 B.n225 B.n140 585
R99 B.n224 B.n223 585
R100 B.n222 B.n141 585
R101 B.n221 B.n220 585
R102 B.n219 B.n142 585
R103 B.n218 B.n217 585
R104 B.n216 B.n143 585
R105 B.n215 B.n214 585
R106 B.n213 B.n144 585
R107 B.n212 B.n211 585
R108 B.n210 B.n145 585
R109 B.n209 B.n208 585
R110 B.n207 B.n146 585
R111 B.n206 B.n205 585
R112 B.n204 B.n147 585
R113 B.n203 B.n202 585
R114 B.n201 B.n148 585
R115 B.n200 B.n199 585
R116 B.n198 B.n149 585
R117 B.n197 B.n196 585
R118 B.n357 B.n356 585
R119 B.n358 B.n95 585
R120 B.n360 B.n359 585
R121 B.n361 B.n94 585
R122 B.n363 B.n362 585
R123 B.n364 B.n93 585
R124 B.n366 B.n365 585
R125 B.n367 B.n92 585
R126 B.n369 B.n368 585
R127 B.n370 B.n91 585
R128 B.n372 B.n371 585
R129 B.n373 B.n90 585
R130 B.n375 B.n374 585
R131 B.n376 B.n89 585
R132 B.n378 B.n377 585
R133 B.n379 B.n88 585
R134 B.n381 B.n380 585
R135 B.n382 B.n87 585
R136 B.n384 B.n383 585
R137 B.n385 B.n86 585
R138 B.n387 B.n386 585
R139 B.n388 B.n85 585
R140 B.n390 B.n389 585
R141 B.n391 B.n84 585
R142 B.n393 B.n392 585
R143 B.n394 B.n83 585
R144 B.n396 B.n395 585
R145 B.n397 B.n82 585
R146 B.n399 B.n398 585
R147 B.n400 B.n81 585
R148 B.n402 B.n401 585
R149 B.n403 B.n80 585
R150 B.n405 B.n404 585
R151 B.n406 B.n79 585
R152 B.n408 B.n407 585
R153 B.n409 B.n78 585
R154 B.n411 B.n410 585
R155 B.n412 B.n77 585
R156 B.n414 B.n413 585
R157 B.n415 B.n76 585
R158 B.n417 B.n416 585
R159 B.n418 B.n75 585
R160 B.n420 B.n419 585
R161 B.n421 B.n74 585
R162 B.n423 B.n422 585
R163 B.n424 B.n73 585
R164 B.n426 B.n425 585
R165 B.n427 B.n72 585
R166 B.n429 B.n428 585
R167 B.n430 B.n71 585
R168 B.n587 B.n14 585
R169 B.n586 B.n585 585
R170 B.n584 B.n15 585
R171 B.n583 B.n582 585
R172 B.n581 B.n16 585
R173 B.n580 B.n579 585
R174 B.n578 B.n17 585
R175 B.n577 B.n576 585
R176 B.n575 B.n18 585
R177 B.n574 B.n573 585
R178 B.n572 B.n19 585
R179 B.n571 B.n570 585
R180 B.n569 B.n20 585
R181 B.n568 B.n567 585
R182 B.n566 B.n21 585
R183 B.n565 B.n564 585
R184 B.n563 B.n22 585
R185 B.n562 B.n561 585
R186 B.n560 B.n23 585
R187 B.n559 B.n558 585
R188 B.n557 B.n24 585
R189 B.n556 B.n555 585
R190 B.n554 B.n25 585
R191 B.n553 B.n552 585
R192 B.n551 B.n26 585
R193 B.n550 B.n549 585
R194 B.n548 B.n27 585
R195 B.n547 B.n546 585
R196 B.n545 B.n28 585
R197 B.n544 B.n543 585
R198 B.n542 B.n29 585
R199 B.n541 B.n540 585
R200 B.n539 B.n30 585
R201 B.n538 B.n537 585
R202 B.n536 B.n31 585
R203 B.n535 B.n534 585
R204 B.n533 B.n32 585
R205 B.n532 B.n531 585
R206 B.n530 B.n33 585
R207 B.n529 B.n528 585
R208 B.n527 B.n34 585
R209 B.n526 B.n525 585
R210 B.n524 B.n35 585
R211 B.n523 B.n522 585
R212 B.n521 B.n36 585
R213 B.n520 B.n519 585
R214 B.n518 B.n37 585
R215 B.n516 B.n515 585
R216 B.n514 B.n40 585
R217 B.n513 B.n512 585
R218 B.n511 B.n41 585
R219 B.n510 B.n509 585
R220 B.n508 B.n42 585
R221 B.n507 B.n506 585
R222 B.n505 B.n43 585
R223 B.n504 B.n503 585
R224 B.n502 B.n44 585
R225 B.n501 B.n500 585
R226 B.n499 B.n45 585
R227 B.n498 B.n497 585
R228 B.n496 B.n49 585
R229 B.n495 B.n494 585
R230 B.n493 B.n50 585
R231 B.n492 B.n491 585
R232 B.n490 B.n51 585
R233 B.n489 B.n488 585
R234 B.n487 B.n52 585
R235 B.n486 B.n485 585
R236 B.n484 B.n53 585
R237 B.n483 B.n482 585
R238 B.n481 B.n54 585
R239 B.n480 B.n479 585
R240 B.n478 B.n55 585
R241 B.n477 B.n476 585
R242 B.n475 B.n56 585
R243 B.n474 B.n473 585
R244 B.n472 B.n57 585
R245 B.n471 B.n470 585
R246 B.n469 B.n58 585
R247 B.n468 B.n467 585
R248 B.n466 B.n59 585
R249 B.n465 B.n464 585
R250 B.n463 B.n60 585
R251 B.n462 B.n461 585
R252 B.n460 B.n61 585
R253 B.n459 B.n458 585
R254 B.n457 B.n62 585
R255 B.n456 B.n455 585
R256 B.n454 B.n63 585
R257 B.n453 B.n452 585
R258 B.n451 B.n64 585
R259 B.n450 B.n449 585
R260 B.n448 B.n65 585
R261 B.n447 B.n446 585
R262 B.n445 B.n66 585
R263 B.n444 B.n443 585
R264 B.n442 B.n67 585
R265 B.n441 B.n440 585
R266 B.n439 B.n68 585
R267 B.n438 B.n437 585
R268 B.n436 B.n69 585
R269 B.n435 B.n434 585
R270 B.n433 B.n70 585
R271 B.n432 B.n431 585
R272 B.n589 B.n588 585
R273 B.n590 B.n13 585
R274 B.n592 B.n591 585
R275 B.n593 B.n12 585
R276 B.n595 B.n594 585
R277 B.n596 B.n11 585
R278 B.n598 B.n597 585
R279 B.n599 B.n10 585
R280 B.n601 B.n600 585
R281 B.n602 B.n9 585
R282 B.n604 B.n603 585
R283 B.n605 B.n8 585
R284 B.n607 B.n606 585
R285 B.n608 B.n7 585
R286 B.n610 B.n609 585
R287 B.n611 B.n6 585
R288 B.n613 B.n612 585
R289 B.n614 B.n5 585
R290 B.n616 B.n615 585
R291 B.n617 B.n4 585
R292 B.n619 B.n618 585
R293 B.n620 B.n3 585
R294 B.n622 B.n621 585
R295 B.n623 B.n0 585
R296 B.n2 B.n1 585
R297 B.n162 B.n161 585
R298 B.n164 B.n163 585
R299 B.n165 B.n160 585
R300 B.n167 B.n166 585
R301 B.n168 B.n159 585
R302 B.n170 B.n169 585
R303 B.n171 B.n158 585
R304 B.n173 B.n172 585
R305 B.n174 B.n157 585
R306 B.n176 B.n175 585
R307 B.n177 B.n156 585
R308 B.n179 B.n178 585
R309 B.n180 B.n155 585
R310 B.n182 B.n181 585
R311 B.n183 B.n154 585
R312 B.n185 B.n184 585
R313 B.n186 B.n153 585
R314 B.n188 B.n187 585
R315 B.n189 B.n152 585
R316 B.n191 B.n190 585
R317 B.n192 B.n151 585
R318 B.n194 B.n193 585
R319 B.n195 B.n150 585
R320 B.n197 B.n150 530.939
R321 B.n357 B.n96 530.939
R322 B.n431 B.n430 530.939
R323 B.n588 B.n587 530.939
R324 B.n125 B.t3 343.856
R325 B.n281 B.t6 343.856
R326 B.n46 B.t0 343.856
R327 B.n38 B.t9 343.856
R328 B.n625 B.n624 256.663
R329 B.n624 B.n623 235.042
R330 B.n624 B.n2 235.042
R331 B.n281 B.t7 167.623
R332 B.n46 B.t2 167.623
R333 B.n125 B.t4 167.606
R334 B.n38 B.t11 167.606
R335 B.n198 B.n197 163.367
R336 B.n199 B.n198 163.367
R337 B.n199 B.n148 163.367
R338 B.n203 B.n148 163.367
R339 B.n204 B.n203 163.367
R340 B.n205 B.n204 163.367
R341 B.n205 B.n146 163.367
R342 B.n209 B.n146 163.367
R343 B.n210 B.n209 163.367
R344 B.n211 B.n210 163.367
R345 B.n211 B.n144 163.367
R346 B.n215 B.n144 163.367
R347 B.n216 B.n215 163.367
R348 B.n217 B.n216 163.367
R349 B.n217 B.n142 163.367
R350 B.n221 B.n142 163.367
R351 B.n222 B.n221 163.367
R352 B.n223 B.n222 163.367
R353 B.n223 B.n140 163.367
R354 B.n227 B.n140 163.367
R355 B.n228 B.n227 163.367
R356 B.n229 B.n228 163.367
R357 B.n229 B.n138 163.367
R358 B.n233 B.n138 163.367
R359 B.n234 B.n233 163.367
R360 B.n235 B.n234 163.367
R361 B.n235 B.n136 163.367
R362 B.n239 B.n136 163.367
R363 B.n240 B.n239 163.367
R364 B.n241 B.n240 163.367
R365 B.n241 B.n134 163.367
R366 B.n245 B.n134 163.367
R367 B.n246 B.n245 163.367
R368 B.n247 B.n246 163.367
R369 B.n247 B.n132 163.367
R370 B.n251 B.n132 163.367
R371 B.n252 B.n251 163.367
R372 B.n253 B.n252 163.367
R373 B.n253 B.n130 163.367
R374 B.n257 B.n130 163.367
R375 B.n258 B.n257 163.367
R376 B.n259 B.n258 163.367
R377 B.n259 B.n128 163.367
R378 B.n263 B.n128 163.367
R379 B.n264 B.n263 163.367
R380 B.n265 B.n264 163.367
R381 B.n265 B.n124 163.367
R382 B.n270 B.n124 163.367
R383 B.n271 B.n270 163.367
R384 B.n272 B.n271 163.367
R385 B.n272 B.n122 163.367
R386 B.n276 B.n122 163.367
R387 B.n277 B.n276 163.367
R388 B.n278 B.n277 163.367
R389 B.n278 B.n120 163.367
R390 B.n285 B.n120 163.367
R391 B.n286 B.n285 163.367
R392 B.n287 B.n286 163.367
R393 B.n287 B.n118 163.367
R394 B.n291 B.n118 163.367
R395 B.n292 B.n291 163.367
R396 B.n293 B.n292 163.367
R397 B.n293 B.n116 163.367
R398 B.n297 B.n116 163.367
R399 B.n298 B.n297 163.367
R400 B.n299 B.n298 163.367
R401 B.n299 B.n114 163.367
R402 B.n303 B.n114 163.367
R403 B.n304 B.n303 163.367
R404 B.n305 B.n304 163.367
R405 B.n305 B.n112 163.367
R406 B.n309 B.n112 163.367
R407 B.n310 B.n309 163.367
R408 B.n311 B.n310 163.367
R409 B.n311 B.n110 163.367
R410 B.n315 B.n110 163.367
R411 B.n316 B.n315 163.367
R412 B.n317 B.n316 163.367
R413 B.n317 B.n108 163.367
R414 B.n321 B.n108 163.367
R415 B.n322 B.n321 163.367
R416 B.n323 B.n322 163.367
R417 B.n323 B.n106 163.367
R418 B.n327 B.n106 163.367
R419 B.n328 B.n327 163.367
R420 B.n329 B.n328 163.367
R421 B.n329 B.n104 163.367
R422 B.n333 B.n104 163.367
R423 B.n334 B.n333 163.367
R424 B.n335 B.n334 163.367
R425 B.n335 B.n102 163.367
R426 B.n339 B.n102 163.367
R427 B.n340 B.n339 163.367
R428 B.n341 B.n340 163.367
R429 B.n341 B.n100 163.367
R430 B.n345 B.n100 163.367
R431 B.n346 B.n345 163.367
R432 B.n347 B.n346 163.367
R433 B.n347 B.n98 163.367
R434 B.n351 B.n98 163.367
R435 B.n352 B.n351 163.367
R436 B.n353 B.n352 163.367
R437 B.n353 B.n96 163.367
R438 B.n430 B.n429 163.367
R439 B.n429 B.n72 163.367
R440 B.n425 B.n72 163.367
R441 B.n425 B.n424 163.367
R442 B.n424 B.n423 163.367
R443 B.n423 B.n74 163.367
R444 B.n419 B.n74 163.367
R445 B.n419 B.n418 163.367
R446 B.n418 B.n417 163.367
R447 B.n417 B.n76 163.367
R448 B.n413 B.n76 163.367
R449 B.n413 B.n412 163.367
R450 B.n412 B.n411 163.367
R451 B.n411 B.n78 163.367
R452 B.n407 B.n78 163.367
R453 B.n407 B.n406 163.367
R454 B.n406 B.n405 163.367
R455 B.n405 B.n80 163.367
R456 B.n401 B.n80 163.367
R457 B.n401 B.n400 163.367
R458 B.n400 B.n399 163.367
R459 B.n399 B.n82 163.367
R460 B.n395 B.n82 163.367
R461 B.n395 B.n394 163.367
R462 B.n394 B.n393 163.367
R463 B.n393 B.n84 163.367
R464 B.n389 B.n84 163.367
R465 B.n389 B.n388 163.367
R466 B.n388 B.n387 163.367
R467 B.n387 B.n86 163.367
R468 B.n383 B.n86 163.367
R469 B.n383 B.n382 163.367
R470 B.n382 B.n381 163.367
R471 B.n381 B.n88 163.367
R472 B.n377 B.n88 163.367
R473 B.n377 B.n376 163.367
R474 B.n376 B.n375 163.367
R475 B.n375 B.n90 163.367
R476 B.n371 B.n90 163.367
R477 B.n371 B.n370 163.367
R478 B.n370 B.n369 163.367
R479 B.n369 B.n92 163.367
R480 B.n365 B.n92 163.367
R481 B.n365 B.n364 163.367
R482 B.n364 B.n363 163.367
R483 B.n363 B.n94 163.367
R484 B.n359 B.n94 163.367
R485 B.n359 B.n358 163.367
R486 B.n358 B.n357 163.367
R487 B.n587 B.n586 163.367
R488 B.n586 B.n15 163.367
R489 B.n582 B.n15 163.367
R490 B.n582 B.n581 163.367
R491 B.n581 B.n580 163.367
R492 B.n580 B.n17 163.367
R493 B.n576 B.n17 163.367
R494 B.n576 B.n575 163.367
R495 B.n575 B.n574 163.367
R496 B.n574 B.n19 163.367
R497 B.n570 B.n19 163.367
R498 B.n570 B.n569 163.367
R499 B.n569 B.n568 163.367
R500 B.n568 B.n21 163.367
R501 B.n564 B.n21 163.367
R502 B.n564 B.n563 163.367
R503 B.n563 B.n562 163.367
R504 B.n562 B.n23 163.367
R505 B.n558 B.n23 163.367
R506 B.n558 B.n557 163.367
R507 B.n557 B.n556 163.367
R508 B.n556 B.n25 163.367
R509 B.n552 B.n25 163.367
R510 B.n552 B.n551 163.367
R511 B.n551 B.n550 163.367
R512 B.n550 B.n27 163.367
R513 B.n546 B.n27 163.367
R514 B.n546 B.n545 163.367
R515 B.n545 B.n544 163.367
R516 B.n544 B.n29 163.367
R517 B.n540 B.n29 163.367
R518 B.n540 B.n539 163.367
R519 B.n539 B.n538 163.367
R520 B.n538 B.n31 163.367
R521 B.n534 B.n31 163.367
R522 B.n534 B.n533 163.367
R523 B.n533 B.n532 163.367
R524 B.n532 B.n33 163.367
R525 B.n528 B.n33 163.367
R526 B.n528 B.n527 163.367
R527 B.n527 B.n526 163.367
R528 B.n526 B.n35 163.367
R529 B.n522 B.n35 163.367
R530 B.n522 B.n521 163.367
R531 B.n521 B.n520 163.367
R532 B.n520 B.n37 163.367
R533 B.n515 B.n37 163.367
R534 B.n515 B.n514 163.367
R535 B.n514 B.n513 163.367
R536 B.n513 B.n41 163.367
R537 B.n509 B.n41 163.367
R538 B.n509 B.n508 163.367
R539 B.n508 B.n507 163.367
R540 B.n507 B.n43 163.367
R541 B.n503 B.n43 163.367
R542 B.n503 B.n502 163.367
R543 B.n502 B.n501 163.367
R544 B.n501 B.n45 163.367
R545 B.n497 B.n45 163.367
R546 B.n497 B.n496 163.367
R547 B.n496 B.n495 163.367
R548 B.n495 B.n50 163.367
R549 B.n491 B.n50 163.367
R550 B.n491 B.n490 163.367
R551 B.n490 B.n489 163.367
R552 B.n489 B.n52 163.367
R553 B.n485 B.n52 163.367
R554 B.n485 B.n484 163.367
R555 B.n484 B.n483 163.367
R556 B.n483 B.n54 163.367
R557 B.n479 B.n54 163.367
R558 B.n479 B.n478 163.367
R559 B.n478 B.n477 163.367
R560 B.n477 B.n56 163.367
R561 B.n473 B.n56 163.367
R562 B.n473 B.n472 163.367
R563 B.n472 B.n471 163.367
R564 B.n471 B.n58 163.367
R565 B.n467 B.n58 163.367
R566 B.n467 B.n466 163.367
R567 B.n466 B.n465 163.367
R568 B.n465 B.n60 163.367
R569 B.n461 B.n60 163.367
R570 B.n461 B.n460 163.367
R571 B.n460 B.n459 163.367
R572 B.n459 B.n62 163.367
R573 B.n455 B.n62 163.367
R574 B.n455 B.n454 163.367
R575 B.n454 B.n453 163.367
R576 B.n453 B.n64 163.367
R577 B.n449 B.n64 163.367
R578 B.n449 B.n448 163.367
R579 B.n448 B.n447 163.367
R580 B.n447 B.n66 163.367
R581 B.n443 B.n66 163.367
R582 B.n443 B.n442 163.367
R583 B.n442 B.n441 163.367
R584 B.n441 B.n68 163.367
R585 B.n437 B.n68 163.367
R586 B.n437 B.n436 163.367
R587 B.n436 B.n435 163.367
R588 B.n435 B.n70 163.367
R589 B.n431 B.n70 163.367
R590 B.n588 B.n13 163.367
R591 B.n592 B.n13 163.367
R592 B.n593 B.n592 163.367
R593 B.n594 B.n593 163.367
R594 B.n594 B.n11 163.367
R595 B.n598 B.n11 163.367
R596 B.n599 B.n598 163.367
R597 B.n600 B.n599 163.367
R598 B.n600 B.n9 163.367
R599 B.n604 B.n9 163.367
R600 B.n605 B.n604 163.367
R601 B.n606 B.n605 163.367
R602 B.n606 B.n7 163.367
R603 B.n610 B.n7 163.367
R604 B.n611 B.n610 163.367
R605 B.n612 B.n611 163.367
R606 B.n612 B.n5 163.367
R607 B.n616 B.n5 163.367
R608 B.n617 B.n616 163.367
R609 B.n618 B.n617 163.367
R610 B.n618 B.n3 163.367
R611 B.n622 B.n3 163.367
R612 B.n623 B.n622 163.367
R613 B.n162 B.n2 163.367
R614 B.n163 B.n162 163.367
R615 B.n163 B.n160 163.367
R616 B.n167 B.n160 163.367
R617 B.n168 B.n167 163.367
R618 B.n169 B.n168 163.367
R619 B.n169 B.n158 163.367
R620 B.n173 B.n158 163.367
R621 B.n174 B.n173 163.367
R622 B.n175 B.n174 163.367
R623 B.n175 B.n156 163.367
R624 B.n179 B.n156 163.367
R625 B.n180 B.n179 163.367
R626 B.n181 B.n180 163.367
R627 B.n181 B.n154 163.367
R628 B.n185 B.n154 163.367
R629 B.n186 B.n185 163.367
R630 B.n187 B.n186 163.367
R631 B.n187 B.n152 163.367
R632 B.n191 B.n152 163.367
R633 B.n192 B.n191 163.367
R634 B.n193 B.n192 163.367
R635 B.n193 B.n150 163.367
R636 B.n282 B.t8 113.32
R637 B.n47 B.t1 113.32
R638 B.n126 B.t5 113.302
R639 B.n39 B.t10 113.302
R640 B.n267 B.n126 59.5399
R641 B.n283 B.n282 59.5399
R642 B.n48 B.n47 59.5399
R643 B.n517 B.n39 59.5399
R644 B.n126 B.n125 54.3035
R645 B.n282 B.n281 54.3035
R646 B.n47 B.n46 54.3035
R647 B.n39 B.n38 54.3035
R648 B.n589 B.n14 34.4981
R649 B.n432 B.n71 34.4981
R650 B.n356 B.n355 34.4981
R651 B.n196 B.n195 34.4981
R652 B B.n625 18.0485
R653 B.n590 B.n589 10.6151
R654 B.n591 B.n590 10.6151
R655 B.n591 B.n12 10.6151
R656 B.n595 B.n12 10.6151
R657 B.n596 B.n595 10.6151
R658 B.n597 B.n596 10.6151
R659 B.n597 B.n10 10.6151
R660 B.n601 B.n10 10.6151
R661 B.n602 B.n601 10.6151
R662 B.n603 B.n602 10.6151
R663 B.n603 B.n8 10.6151
R664 B.n607 B.n8 10.6151
R665 B.n608 B.n607 10.6151
R666 B.n609 B.n608 10.6151
R667 B.n609 B.n6 10.6151
R668 B.n613 B.n6 10.6151
R669 B.n614 B.n613 10.6151
R670 B.n615 B.n614 10.6151
R671 B.n615 B.n4 10.6151
R672 B.n619 B.n4 10.6151
R673 B.n620 B.n619 10.6151
R674 B.n621 B.n620 10.6151
R675 B.n621 B.n0 10.6151
R676 B.n585 B.n14 10.6151
R677 B.n585 B.n584 10.6151
R678 B.n584 B.n583 10.6151
R679 B.n583 B.n16 10.6151
R680 B.n579 B.n16 10.6151
R681 B.n579 B.n578 10.6151
R682 B.n578 B.n577 10.6151
R683 B.n577 B.n18 10.6151
R684 B.n573 B.n18 10.6151
R685 B.n573 B.n572 10.6151
R686 B.n572 B.n571 10.6151
R687 B.n571 B.n20 10.6151
R688 B.n567 B.n20 10.6151
R689 B.n567 B.n566 10.6151
R690 B.n566 B.n565 10.6151
R691 B.n565 B.n22 10.6151
R692 B.n561 B.n22 10.6151
R693 B.n561 B.n560 10.6151
R694 B.n560 B.n559 10.6151
R695 B.n559 B.n24 10.6151
R696 B.n555 B.n24 10.6151
R697 B.n555 B.n554 10.6151
R698 B.n554 B.n553 10.6151
R699 B.n553 B.n26 10.6151
R700 B.n549 B.n26 10.6151
R701 B.n549 B.n548 10.6151
R702 B.n548 B.n547 10.6151
R703 B.n547 B.n28 10.6151
R704 B.n543 B.n28 10.6151
R705 B.n543 B.n542 10.6151
R706 B.n542 B.n541 10.6151
R707 B.n541 B.n30 10.6151
R708 B.n537 B.n30 10.6151
R709 B.n537 B.n536 10.6151
R710 B.n536 B.n535 10.6151
R711 B.n535 B.n32 10.6151
R712 B.n531 B.n32 10.6151
R713 B.n531 B.n530 10.6151
R714 B.n530 B.n529 10.6151
R715 B.n529 B.n34 10.6151
R716 B.n525 B.n34 10.6151
R717 B.n525 B.n524 10.6151
R718 B.n524 B.n523 10.6151
R719 B.n523 B.n36 10.6151
R720 B.n519 B.n36 10.6151
R721 B.n519 B.n518 10.6151
R722 B.n516 B.n40 10.6151
R723 B.n512 B.n40 10.6151
R724 B.n512 B.n511 10.6151
R725 B.n511 B.n510 10.6151
R726 B.n510 B.n42 10.6151
R727 B.n506 B.n42 10.6151
R728 B.n506 B.n505 10.6151
R729 B.n505 B.n504 10.6151
R730 B.n504 B.n44 10.6151
R731 B.n500 B.n499 10.6151
R732 B.n499 B.n498 10.6151
R733 B.n498 B.n49 10.6151
R734 B.n494 B.n49 10.6151
R735 B.n494 B.n493 10.6151
R736 B.n493 B.n492 10.6151
R737 B.n492 B.n51 10.6151
R738 B.n488 B.n51 10.6151
R739 B.n488 B.n487 10.6151
R740 B.n487 B.n486 10.6151
R741 B.n486 B.n53 10.6151
R742 B.n482 B.n53 10.6151
R743 B.n482 B.n481 10.6151
R744 B.n481 B.n480 10.6151
R745 B.n480 B.n55 10.6151
R746 B.n476 B.n55 10.6151
R747 B.n476 B.n475 10.6151
R748 B.n475 B.n474 10.6151
R749 B.n474 B.n57 10.6151
R750 B.n470 B.n57 10.6151
R751 B.n470 B.n469 10.6151
R752 B.n469 B.n468 10.6151
R753 B.n468 B.n59 10.6151
R754 B.n464 B.n59 10.6151
R755 B.n464 B.n463 10.6151
R756 B.n463 B.n462 10.6151
R757 B.n462 B.n61 10.6151
R758 B.n458 B.n61 10.6151
R759 B.n458 B.n457 10.6151
R760 B.n457 B.n456 10.6151
R761 B.n456 B.n63 10.6151
R762 B.n452 B.n63 10.6151
R763 B.n452 B.n451 10.6151
R764 B.n451 B.n450 10.6151
R765 B.n450 B.n65 10.6151
R766 B.n446 B.n65 10.6151
R767 B.n446 B.n445 10.6151
R768 B.n445 B.n444 10.6151
R769 B.n444 B.n67 10.6151
R770 B.n440 B.n67 10.6151
R771 B.n440 B.n439 10.6151
R772 B.n439 B.n438 10.6151
R773 B.n438 B.n69 10.6151
R774 B.n434 B.n69 10.6151
R775 B.n434 B.n433 10.6151
R776 B.n433 B.n432 10.6151
R777 B.n428 B.n71 10.6151
R778 B.n428 B.n427 10.6151
R779 B.n427 B.n426 10.6151
R780 B.n426 B.n73 10.6151
R781 B.n422 B.n73 10.6151
R782 B.n422 B.n421 10.6151
R783 B.n421 B.n420 10.6151
R784 B.n420 B.n75 10.6151
R785 B.n416 B.n75 10.6151
R786 B.n416 B.n415 10.6151
R787 B.n415 B.n414 10.6151
R788 B.n414 B.n77 10.6151
R789 B.n410 B.n77 10.6151
R790 B.n410 B.n409 10.6151
R791 B.n409 B.n408 10.6151
R792 B.n408 B.n79 10.6151
R793 B.n404 B.n79 10.6151
R794 B.n404 B.n403 10.6151
R795 B.n403 B.n402 10.6151
R796 B.n402 B.n81 10.6151
R797 B.n398 B.n81 10.6151
R798 B.n398 B.n397 10.6151
R799 B.n397 B.n396 10.6151
R800 B.n396 B.n83 10.6151
R801 B.n392 B.n83 10.6151
R802 B.n392 B.n391 10.6151
R803 B.n391 B.n390 10.6151
R804 B.n390 B.n85 10.6151
R805 B.n386 B.n85 10.6151
R806 B.n386 B.n385 10.6151
R807 B.n385 B.n384 10.6151
R808 B.n384 B.n87 10.6151
R809 B.n380 B.n87 10.6151
R810 B.n380 B.n379 10.6151
R811 B.n379 B.n378 10.6151
R812 B.n378 B.n89 10.6151
R813 B.n374 B.n89 10.6151
R814 B.n374 B.n373 10.6151
R815 B.n373 B.n372 10.6151
R816 B.n372 B.n91 10.6151
R817 B.n368 B.n91 10.6151
R818 B.n368 B.n367 10.6151
R819 B.n367 B.n366 10.6151
R820 B.n366 B.n93 10.6151
R821 B.n362 B.n93 10.6151
R822 B.n362 B.n361 10.6151
R823 B.n361 B.n360 10.6151
R824 B.n360 B.n95 10.6151
R825 B.n356 B.n95 10.6151
R826 B.n161 B.n1 10.6151
R827 B.n164 B.n161 10.6151
R828 B.n165 B.n164 10.6151
R829 B.n166 B.n165 10.6151
R830 B.n166 B.n159 10.6151
R831 B.n170 B.n159 10.6151
R832 B.n171 B.n170 10.6151
R833 B.n172 B.n171 10.6151
R834 B.n172 B.n157 10.6151
R835 B.n176 B.n157 10.6151
R836 B.n177 B.n176 10.6151
R837 B.n178 B.n177 10.6151
R838 B.n178 B.n155 10.6151
R839 B.n182 B.n155 10.6151
R840 B.n183 B.n182 10.6151
R841 B.n184 B.n183 10.6151
R842 B.n184 B.n153 10.6151
R843 B.n188 B.n153 10.6151
R844 B.n189 B.n188 10.6151
R845 B.n190 B.n189 10.6151
R846 B.n190 B.n151 10.6151
R847 B.n194 B.n151 10.6151
R848 B.n195 B.n194 10.6151
R849 B.n196 B.n149 10.6151
R850 B.n200 B.n149 10.6151
R851 B.n201 B.n200 10.6151
R852 B.n202 B.n201 10.6151
R853 B.n202 B.n147 10.6151
R854 B.n206 B.n147 10.6151
R855 B.n207 B.n206 10.6151
R856 B.n208 B.n207 10.6151
R857 B.n208 B.n145 10.6151
R858 B.n212 B.n145 10.6151
R859 B.n213 B.n212 10.6151
R860 B.n214 B.n213 10.6151
R861 B.n214 B.n143 10.6151
R862 B.n218 B.n143 10.6151
R863 B.n219 B.n218 10.6151
R864 B.n220 B.n219 10.6151
R865 B.n220 B.n141 10.6151
R866 B.n224 B.n141 10.6151
R867 B.n225 B.n224 10.6151
R868 B.n226 B.n225 10.6151
R869 B.n226 B.n139 10.6151
R870 B.n230 B.n139 10.6151
R871 B.n231 B.n230 10.6151
R872 B.n232 B.n231 10.6151
R873 B.n232 B.n137 10.6151
R874 B.n236 B.n137 10.6151
R875 B.n237 B.n236 10.6151
R876 B.n238 B.n237 10.6151
R877 B.n238 B.n135 10.6151
R878 B.n242 B.n135 10.6151
R879 B.n243 B.n242 10.6151
R880 B.n244 B.n243 10.6151
R881 B.n244 B.n133 10.6151
R882 B.n248 B.n133 10.6151
R883 B.n249 B.n248 10.6151
R884 B.n250 B.n249 10.6151
R885 B.n250 B.n131 10.6151
R886 B.n254 B.n131 10.6151
R887 B.n255 B.n254 10.6151
R888 B.n256 B.n255 10.6151
R889 B.n256 B.n129 10.6151
R890 B.n260 B.n129 10.6151
R891 B.n261 B.n260 10.6151
R892 B.n262 B.n261 10.6151
R893 B.n262 B.n127 10.6151
R894 B.n266 B.n127 10.6151
R895 B.n269 B.n268 10.6151
R896 B.n269 B.n123 10.6151
R897 B.n273 B.n123 10.6151
R898 B.n274 B.n273 10.6151
R899 B.n275 B.n274 10.6151
R900 B.n275 B.n121 10.6151
R901 B.n279 B.n121 10.6151
R902 B.n280 B.n279 10.6151
R903 B.n284 B.n280 10.6151
R904 B.n288 B.n119 10.6151
R905 B.n289 B.n288 10.6151
R906 B.n290 B.n289 10.6151
R907 B.n290 B.n117 10.6151
R908 B.n294 B.n117 10.6151
R909 B.n295 B.n294 10.6151
R910 B.n296 B.n295 10.6151
R911 B.n296 B.n115 10.6151
R912 B.n300 B.n115 10.6151
R913 B.n301 B.n300 10.6151
R914 B.n302 B.n301 10.6151
R915 B.n302 B.n113 10.6151
R916 B.n306 B.n113 10.6151
R917 B.n307 B.n306 10.6151
R918 B.n308 B.n307 10.6151
R919 B.n308 B.n111 10.6151
R920 B.n312 B.n111 10.6151
R921 B.n313 B.n312 10.6151
R922 B.n314 B.n313 10.6151
R923 B.n314 B.n109 10.6151
R924 B.n318 B.n109 10.6151
R925 B.n319 B.n318 10.6151
R926 B.n320 B.n319 10.6151
R927 B.n320 B.n107 10.6151
R928 B.n324 B.n107 10.6151
R929 B.n325 B.n324 10.6151
R930 B.n326 B.n325 10.6151
R931 B.n326 B.n105 10.6151
R932 B.n330 B.n105 10.6151
R933 B.n331 B.n330 10.6151
R934 B.n332 B.n331 10.6151
R935 B.n332 B.n103 10.6151
R936 B.n336 B.n103 10.6151
R937 B.n337 B.n336 10.6151
R938 B.n338 B.n337 10.6151
R939 B.n338 B.n101 10.6151
R940 B.n342 B.n101 10.6151
R941 B.n343 B.n342 10.6151
R942 B.n344 B.n343 10.6151
R943 B.n344 B.n99 10.6151
R944 B.n348 B.n99 10.6151
R945 B.n349 B.n348 10.6151
R946 B.n350 B.n349 10.6151
R947 B.n350 B.n97 10.6151
R948 B.n354 B.n97 10.6151
R949 B.n355 B.n354 10.6151
R950 B.n518 B.n517 9.36635
R951 B.n500 B.n48 9.36635
R952 B.n267 B.n266 9.36635
R953 B.n283 B.n119 9.36635
R954 B.n625 B.n0 8.11757
R955 B.n625 B.n1 8.11757
R956 B.n517 B.n516 1.24928
R957 B.n48 B.n44 1.24928
R958 B.n268 B.n267 1.24928
R959 B.n284 B.n283 1.24928
R960 VN VN.t0 231.107
R961 VN VN.t1 185.565
R962 VDD2.n0 VDD2.t0 115.171
R963 VDD2.n0 VDD2.t1 74.6668
R964 VDD2 VDD2.n0 0.662138
C0 VDD1 VTAIL 5.56712f
C1 B VN 1.05442f
C2 VDD2 VN 3.16338f
C3 VP VN 5.74955f
C4 B VDD2 1.86937f
C5 VP B 1.49113f
C6 VP VDD2 0.328106f
C7 w_n2090_n3756# VN 2.90903f
C8 w_n2090_n3756# B 9.2128f
C9 VDD1 VN 0.148396f
C10 w_n2090_n3756# VDD2 1.9259f
C11 B VDD1 1.84044f
C12 VP w_n2090_n3756# 3.17498f
C13 VDD1 VDD2 0.659266f
C14 VP VDD1 3.34013f
C15 w_n2090_n3756# VDD1 1.90158f
C16 VTAIL VN 2.73025f
C17 B VTAIL 4.03527f
C18 VDD2 VTAIL 5.61624f
C19 VP VTAIL 2.74458f
C20 w_n2090_n3756# VTAIL 3.03808f
C21 VDD2 VSUBS 0.938425f
C22 VDD1 VSUBS 4.67326f
C23 VTAIL VSUBS 1.06614f
C24 VN VSUBS 8.17465f
C25 VP VSUBS 1.717026f
C26 B VSUBS 3.977321f
C27 w_n2090_n3756# VSUBS 96.38239f
C28 VDD2.t0 VSUBS 2.92704f
C29 VDD2.t1 VSUBS 2.31413f
C30 VDD2.n0 VSUBS 3.4369f
C31 VN.t1 VSUBS 4.07509f
C32 VN.t0 VSUBS 4.6977f
C33 B.n0 VSUBS 0.005165f
C34 B.n1 VSUBS 0.005165f
C35 B.n2 VSUBS 0.007638f
C36 B.n3 VSUBS 0.005853f
C37 B.n4 VSUBS 0.005853f
C38 B.n5 VSUBS 0.005853f
C39 B.n6 VSUBS 0.005853f
C40 B.n7 VSUBS 0.005853f
C41 B.n8 VSUBS 0.005853f
C42 B.n9 VSUBS 0.005853f
C43 B.n10 VSUBS 0.005853f
C44 B.n11 VSUBS 0.005853f
C45 B.n12 VSUBS 0.005853f
C46 B.n13 VSUBS 0.005853f
C47 B.n14 VSUBS 0.014499f
C48 B.n15 VSUBS 0.005853f
C49 B.n16 VSUBS 0.005853f
C50 B.n17 VSUBS 0.005853f
C51 B.n18 VSUBS 0.005853f
C52 B.n19 VSUBS 0.005853f
C53 B.n20 VSUBS 0.005853f
C54 B.n21 VSUBS 0.005853f
C55 B.n22 VSUBS 0.005853f
C56 B.n23 VSUBS 0.005853f
C57 B.n24 VSUBS 0.005853f
C58 B.n25 VSUBS 0.005853f
C59 B.n26 VSUBS 0.005853f
C60 B.n27 VSUBS 0.005853f
C61 B.n28 VSUBS 0.005853f
C62 B.n29 VSUBS 0.005853f
C63 B.n30 VSUBS 0.005853f
C64 B.n31 VSUBS 0.005853f
C65 B.n32 VSUBS 0.005853f
C66 B.n33 VSUBS 0.005853f
C67 B.n34 VSUBS 0.005853f
C68 B.n35 VSUBS 0.005853f
C69 B.n36 VSUBS 0.005853f
C70 B.n37 VSUBS 0.005853f
C71 B.t10 VSUBS 0.385564f
C72 B.t11 VSUBS 0.402195f
C73 B.t9 VSUBS 1.2943f
C74 B.n38 VSUBS 0.21017f
C75 B.n39 VSUBS 0.059682f
C76 B.n40 VSUBS 0.005853f
C77 B.n41 VSUBS 0.005853f
C78 B.n42 VSUBS 0.005853f
C79 B.n43 VSUBS 0.005853f
C80 B.n44 VSUBS 0.003271f
C81 B.n45 VSUBS 0.005853f
C82 B.t1 VSUBS 0.385554f
C83 B.t2 VSUBS 0.402188f
C84 B.t0 VSUBS 1.2943f
C85 B.n46 VSUBS 0.210178f
C86 B.n47 VSUBS 0.059692f
C87 B.n48 VSUBS 0.013562f
C88 B.n49 VSUBS 0.005853f
C89 B.n50 VSUBS 0.005853f
C90 B.n51 VSUBS 0.005853f
C91 B.n52 VSUBS 0.005853f
C92 B.n53 VSUBS 0.005853f
C93 B.n54 VSUBS 0.005853f
C94 B.n55 VSUBS 0.005853f
C95 B.n56 VSUBS 0.005853f
C96 B.n57 VSUBS 0.005853f
C97 B.n58 VSUBS 0.005853f
C98 B.n59 VSUBS 0.005853f
C99 B.n60 VSUBS 0.005853f
C100 B.n61 VSUBS 0.005853f
C101 B.n62 VSUBS 0.005853f
C102 B.n63 VSUBS 0.005853f
C103 B.n64 VSUBS 0.005853f
C104 B.n65 VSUBS 0.005853f
C105 B.n66 VSUBS 0.005853f
C106 B.n67 VSUBS 0.005853f
C107 B.n68 VSUBS 0.005853f
C108 B.n69 VSUBS 0.005853f
C109 B.n70 VSUBS 0.005853f
C110 B.n71 VSUBS 0.013908f
C111 B.n72 VSUBS 0.005853f
C112 B.n73 VSUBS 0.005853f
C113 B.n74 VSUBS 0.005853f
C114 B.n75 VSUBS 0.005853f
C115 B.n76 VSUBS 0.005853f
C116 B.n77 VSUBS 0.005853f
C117 B.n78 VSUBS 0.005853f
C118 B.n79 VSUBS 0.005853f
C119 B.n80 VSUBS 0.005853f
C120 B.n81 VSUBS 0.005853f
C121 B.n82 VSUBS 0.005853f
C122 B.n83 VSUBS 0.005853f
C123 B.n84 VSUBS 0.005853f
C124 B.n85 VSUBS 0.005853f
C125 B.n86 VSUBS 0.005853f
C126 B.n87 VSUBS 0.005853f
C127 B.n88 VSUBS 0.005853f
C128 B.n89 VSUBS 0.005853f
C129 B.n90 VSUBS 0.005853f
C130 B.n91 VSUBS 0.005853f
C131 B.n92 VSUBS 0.005853f
C132 B.n93 VSUBS 0.005853f
C133 B.n94 VSUBS 0.005853f
C134 B.n95 VSUBS 0.005853f
C135 B.n96 VSUBS 0.014499f
C136 B.n97 VSUBS 0.005853f
C137 B.n98 VSUBS 0.005853f
C138 B.n99 VSUBS 0.005853f
C139 B.n100 VSUBS 0.005853f
C140 B.n101 VSUBS 0.005853f
C141 B.n102 VSUBS 0.005853f
C142 B.n103 VSUBS 0.005853f
C143 B.n104 VSUBS 0.005853f
C144 B.n105 VSUBS 0.005853f
C145 B.n106 VSUBS 0.005853f
C146 B.n107 VSUBS 0.005853f
C147 B.n108 VSUBS 0.005853f
C148 B.n109 VSUBS 0.005853f
C149 B.n110 VSUBS 0.005853f
C150 B.n111 VSUBS 0.005853f
C151 B.n112 VSUBS 0.005853f
C152 B.n113 VSUBS 0.005853f
C153 B.n114 VSUBS 0.005853f
C154 B.n115 VSUBS 0.005853f
C155 B.n116 VSUBS 0.005853f
C156 B.n117 VSUBS 0.005853f
C157 B.n118 VSUBS 0.005853f
C158 B.n119 VSUBS 0.005509f
C159 B.n120 VSUBS 0.005853f
C160 B.n121 VSUBS 0.005853f
C161 B.n122 VSUBS 0.005853f
C162 B.n123 VSUBS 0.005853f
C163 B.n124 VSUBS 0.005853f
C164 B.t5 VSUBS 0.385564f
C165 B.t4 VSUBS 0.402195f
C166 B.t3 VSUBS 1.2943f
C167 B.n125 VSUBS 0.21017f
C168 B.n126 VSUBS 0.059682f
C169 B.n127 VSUBS 0.005853f
C170 B.n128 VSUBS 0.005853f
C171 B.n129 VSUBS 0.005853f
C172 B.n130 VSUBS 0.005853f
C173 B.n131 VSUBS 0.005853f
C174 B.n132 VSUBS 0.005853f
C175 B.n133 VSUBS 0.005853f
C176 B.n134 VSUBS 0.005853f
C177 B.n135 VSUBS 0.005853f
C178 B.n136 VSUBS 0.005853f
C179 B.n137 VSUBS 0.005853f
C180 B.n138 VSUBS 0.005853f
C181 B.n139 VSUBS 0.005853f
C182 B.n140 VSUBS 0.005853f
C183 B.n141 VSUBS 0.005853f
C184 B.n142 VSUBS 0.005853f
C185 B.n143 VSUBS 0.005853f
C186 B.n144 VSUBS 0.005853f
C187 B.n145 VSUBS 0.005853f
C188 B.n146 VSUBS 0.005853f
C189 B.n147 VSUBS 0.005853f
C190 B.n148 VSUBS 0.005853f
C191 B.n149 VSUBS 0.005853f
C192 B.n150 VSUBS 0.013908f
C193 B.n151 VSUBS 0.005853f
C194 B.n152 VSUBS 0.005853f
C195 B.n153 VSUBS 0.005853f
C196 B.n154 VSUBS 0.005853f
C197 B.n155 VSUBS 0.005853f
C198 B.n156 VSUBS 0.005853f
C199 B.n157 VSUBS 0.005853f
C200 B.n158 VSUBS 0.005853f
C201 B.n159 VSUBS 0.005853f
C202 B.n160 VSUBS 0.005853f
C203 B.n161 VSUBS 0.005853f
C204 B.n162 VSUBS 0.005853f
C205 B.n163 VSUBS 0.005853f
C206 B.n164 VSUBS 0.005853f
C207 B.n165 VSUBS 0.005853f
C208 B.n166 VSUBS 0.005853f
C209 B.n167 VSUBS 0.005853f
C210 B.n168 VSUBS 0.005853f
C211 B.n169 VSUBS 0.005853f
C212 B.n170 VSUBS 0.005853f
C213 B.n171 VSUBS 0.005853f
C214 B.n172 VSUBS 0.005853f
C215 B.n173 VSUBS 0.005853f
C216 B.n174 VSUBS 0.005853f
C217 B.n175 VSUBS 0.005853f
C218 B.n176 VSUBS 0.005853f
C219 B.n177 VSUBS 0.005853f
C220 B.n178 VSUBS 0.005853f
C221 B.n179 VSUBS 0.005853f
C222 B.n180 VSUBS 0.005853f
C223 B.n181 VSUBS 0.005853f
C224 B.n182 VSUBS 0.005853f
C225 B.n183 VSUBS 0.005853f
C226 B.n184 VSUBS 0.005853f
C227 B.n185 VSUBS 0.005853f
C228 B.n186 VSUBS 0.005853f
C229 B.n187 VSUBS 0.005853f
C230 B.n188 VSUBS 0.005853f
C231 B.n189 VSUBS 0.005853f
C232 B.n190 VSUBS 0.005853f
C233 B.n191 VSUBS 0.005853f
C234 B.n192 VSUBS 0.005853f
C235 B.n193 VSUBS 0.005853f
C236 B.n194 VSUBS 0.005853f
C237 B.n195 VSUBS 0.013908f
C238 B.n196 VSUBS 0.014499f
C239 B.n197 VSUBS 0.014499f
C240 B.n198 VSUBS 0.005853f
C241 B.n199 VSUBS 0.005853f
C242 B.n200 VSUBS 0.005853f
C243 B.n201 VSUBS 0.005853f
C244 B.n202 VSUBS 0.005853f
C245 B.n203 VSUBS 0.005853f
C246 B.n204 VSUBS 0.005853f
C247 B.n205 VSUBS 0.005853f
C248 B.n206 VSUBS 0.005853f
C249 B.n207 VSUBS 0.005853f
C250 B.n208 VSUBS 0.005853f
C251 B.n209 VSUBS 0.005853f
C252 B.n210 VSUBS 0.005853f
C253 B.n211 VSUBS 0.005853f
C254 B.n212 VSUBS 0.005853f
C255 B.n213 VSUBS 0.005853f
C256 B.n214 VSUBS 0.005853f
C257 B.n215 VSUBS 0.005853f
C258 B.n216 VSUBS 0.005853f
C259 B.n217 VSUBS 0.005853f
C260 B.n218 VSUBS 0.005853f
C261 B.n219 VSUBS 0.005853f
C262 B.n220 VSUBS 0.005853f
C263 B.n221 VSUBS 0.005853f
C264 B.n222 VSUBS 0.005853f
C265 B.n223 VSUBS 0.005853f
C266 B.n224 VSUBS 0.005853f
C267 B.n225 VSUBS 0.005853f
C268 B.n226 VSUBS 0.005853f
C269 B.n227 VSUBS 0.005853f
C270 B.n228 VSUBS 0.005853f
C271 B.n229 VSUBS 0.005853f
C272 B.n230 VSUBS 0.005853f
C273 B.n231 VSUBS 0.005853f
C274 B.n232 VSUBS 0.005853f
C275 B.n233 VSUBS 0.005853f
C276 B.n234 VSUBS 0.005853f
C277 B.n235 VSUBS 0.005853f
C278 B.n236 VSUBS 0.005853f
C279 B.n237 VSUBS 0.005853f
C280 B.n238 VSUBS 0.005853f
C281 B.n239 VSUBS 0.005853f
C282 B.n240 VSUBS 0.005853f
C283 B.n241 VSUBS 0.005853f
C284 B.n242 VSUBS 0.005853f
C285 B.n243 VSUBS 0.005853f
C286 B.n244 VSUBS 0.005853f
C287 B.n245 VSUBS 0.005853f
C288 B.n246 VSUBS 0.005853f
C289 B.n247 VSUBS 0.005853f
C290 B.n248 VSUBS 0.005853f
C291 B.n249 VSUBS 0.005853f
C292 B.n250 VSUBS 0.005853f
C293 B.n251 VSUBS 0.005853f
C294 B.n252 VSUBS 0.005853f
C295 B.n253 VSUBS 0.005853f
C296 B.n254 VSUBS 0.005853f
C297 B.n255 VSUBS 0.005853f
C298 B.n256 VSUBS 0.005853f
C299 B.n257 VSUBS 0.005853f
C300 B.n258 VSUBS 0.005853f
C301 B.n259 VSUBS 0.005853f
C302 B.n260 VSUBS 0.005853f
C303 B.n261 VSUBS 0.005853f
C304 B.n262 VSUBS 0.005853f
C305 B.n263 VSUBS 0.005853f
C306 B.n264 VSUBS 0.005853f
C307 B.n265 VSUBS 0.005853f
C308 B.n266 VSUBS 0.005509f
C309 B.n267 VSUBS 0.013562f
C310 B.n268 VSUBS 0.003271f
C311 B.n269 VSUBS 0.005853f
C312 B.n270 VSUBS 0.005853f
C313 B.n271 VSUBS 0.005853f
C314 B.n272 VSUBS 0.005853f
C315 B.n273 VSUBS 0.005853f
C316 B.n274 VSUBS 0.005853f
C317 B.n275 VSUBS 0.005853f
C318 B.n276 VSUBS 0.005853f
C319 B.n277 VSUBS 0.005853f
C320 B.n278 VSUBS 0.005853f
C321 B.n279 VSUBS 0.005853f
C322 B.n280 VSUBS 0.005853f
C323 B.t8 VSUBS 0.385554f
C324 B.t7 VSUBS 0.402188f
C325 B.t6 VSUBS 1.2943f
C326 B.n281 VSUBS 0.210178f
C327 B.n282 VSUBS 0.059692f
C328 B.n283 VSUBS 0.013562f
C329 B.n284 VSUBS 0.003271f
C330 B.n285 VSUBS 0.005853f
C331 B.n286 VSUBS 0.005853f
C332 B.n287 VSUBS 0.005853f
C333 B.n288 VSUBS 0.005853f
C334 B.n289 VSUBS 0.005853f
C335 B.n290 VSUBS 0.005853f
C336 B.n291 VSUBS 0.005853f
C337 B.n292 VSUBS 0.005853f
C338 B.n293 VSUBS 0.005853f
C339 B.n294 VSUBS 0.005853f
C340 B.n295 VSUBS 0.005853f
C341 B.n296 VSUBS 0.005853f
C342 B.n297 VSUBS 0.005853f
C343 B.n298 VSUBS 0.005853f
C344 B.n299 VSUBS 0.005853f
C345 B.n300 VSUBS 0.005853f
C346 B.n301 VSUBS 0.005853f
C347 B.n302 VSUBS 0.005853f
C348 B.n303 VSUBS 0.005853f
C349 B.n304 VSUBS 0.005853f
C350 B.n305 VSUBS 0.005853f
C351 B.n306 VSUBS 0.005853f
C352 B.n307 VSUBS 0.005853f
C353 B.n308 VSUBS 0.005853f
C354 B.n309 VSUBS 0.005853f
C355 B.n310 VSUBS 0.005853f
C356 B.n311 VSUBS 0.005853f
C357 B.n312 VSUBS 0.005853f
C358 B.n313 VSUBS 0.005853f
C359 B.n314 VSUBS 0.005853f
C360 B.n315 VSUBS 0.005853f
C361 B.n316 VSUBS 0.005853f
C362 B.n317 VSUBS 0.005853f
C363 B.n318 VSUBS 0.005853f
C364 B.n319 VSUBS 0.005853f
C365 B.n320 VSUBS 0.005853f
C366 B.n321 VSUBS 0.005853f
C367 B.n322 VSUBS 0.005853f
C368 B.n323 VSUBS 0.005853f
C369 B.n324 VSUBS 0.005853f
C370 B.n325 VSUBS 0.005853f
C371 B.n326 VSUBS 0.005853f
C372 B.n327 VSUBS 0.005853f
C373 B.n328 VSUBS 0.005853f
C374 B.n329 VSUBS 0.005853f
C375 B.n330 VSUBS 0.005853f
C376 B.n331 VSUBS 0.005853f
C377 B.n332 VSUBS 0.005853f
C378 B.n333 VSUBS 0.005853f
C379 B.n334 VSUBS 0.005853f
C380 B.n335 VSUBS 0.005853f
C381 B.n336 VSUBS 0.005853f
C382 B.n337 VSUBS 0.005853f
C383 B.n338 VSUBS 0.005853f
C384 B.n339 VSUBS 0.005853f
C385 B.n340 VSUBS 0.005853f
C386 B.n341 VSUBS 0.005853f
C387 B.n342 VSUBS 0.005853f
C388 B.n343 VSUBS 0.005853f
C389 B.n344 VSUBS 0.005853f
C390 B.n345 VSUBS 0.005853f
C391 B.n346 VSUBS 0.005853f
C392 B.n347 VSUBS 0.005853f
C393 B.n348 VSUBS 0.005853f
C394 B.n349 VSUBS 0.005853f
C395 B.n350 VSUBS 0.005853f
C396 B.n351 VSUBS 0.005853f
C397 B.n352 VSUBS 0.005853f
C398 B.n353 VSUBS 0.005853f
C399 B.n354 VSUBS 0.005853f
C400 B.n355 VSUBS 0.013844f
C401 B.n356 VSUBS 0.014562f
C402 B.n357 VSUBS 0.013908f
C403 B.n358 VSUBS 0.005853f
C404 B.n359 VSUBS 0.005853f
C405 B.n360 VSUBS 0.005853f
C406 B.n361 VSUBS 0.005853f
C407 B.n362 VSUBS 0.005853f
C408 B.n363 VSUBS 0.005853f
C409 B.n364 VSUBS 0.005853f
C410 B.n365 VSUBS 0.005853f
C411 B.n366 VSUBS 0.005853f
C412 B.n367 VSUBS 0.005853f
C413 B.n368 VSUBS 0.005853f
C414 B.n369 VSUBS 0.005853f
C415 B.n370 VSUBS 0.005853f
C416 B.n371 VSUBS 0.005853f
C417 B.n372 VSUBS 0.005853f
C418 B.n373 VSUBS 0.005853f
C419 B.n374 VSUBS 0.005853f
C420 B.n375 VSUBS 0.005853f
C421 B.n376 VSUBS 0.005853f
C422 B.n377 VSUBS 0.005853f
C423 B.n378 VSUBS 0.005853f
C424 B.n379 VSUBS 0.005853f
C425 B.n380 VSUBS 0.005853f
C426 B.n381 VSUBS 0.005853f
C427 B.n382 VSUBS 0.005853f
C428 B.n383 VSUBS 0.005853f
C429 B.n384 VSUBS 0.005853f
C430 B.n385 VSUBS 0.005853f
C431 B.n386 VSUBS 0.005853f
C432 B.n387 VSUBS 0.005853f
C433 B.n388 VSUBS 0.005853f
C434 B.n389 VSUBS 0.005853f
C435 B.n390 VSUBS 0.005853f
C436 B.n391 VSUBS 0.005853f
C437 B.n392 VSUBS 0.005853f
C438 B.n393 VSUBS 0.005853f
C439 B.n394 VSUBS 0.005853f
C440 B.n395 VSUBS 0.005853f
C441 B.n396 VSUBS 0.005853f
C442 B.n397 VSUBS 0.005853f
C443 B.n398 VSUBS 0.005853f
C444 B.n399 VSUBS 0.005853f
C445 B.n400 VSUBS 0.005853f
C446 B.n401 VSUBS 0.005853f
C447 B.n402 VSUBS 0.005853f
C448 B.n403 VSUBS 0.005853f
C449 B.n404 VSUBS 0.005853f
C450 B.n405 VSUBS 0.005853f
C451 B.n406 VSUBS 0.005853f
C452 B.n407 VSUBS 0.005853f
C453 B.n408 VSUBS 0.005853f
C454 B.n409 VSUBS 0.005853f
C455 B.n410 VSUBS 0.005853f
C456 B.n411 VSUBS 0.005853f
C457 B.n412 VSUBS 0.005853f
C458 B.n413 VSUBS 0.005853f
C459 B.n414 VSUBS 0.005853f
C460 B.n415 VSUBS 0.005853f
C461 B.n416 VSUBS 0.005853f
C462 B.n417 VSUBS 0.005853f
C463 B.n418 VSUBS 0.005853f
C464 B.n419 VSUBS 0.005853f
C465 B.n420 VSUBS 0.005853f
C466 B.n421 VSUBS 0.005853f
C467 B.n422 VSUBS 0.005853f
C468 B.n423 VSUBS 0.005853f
C469 B.n424 VSUBS 0.005853f
C470 B.n425 VSUBS 0.005853f
C471 B.n426 VSUBS 0.005853f
C472 B.n427 VSUBS 0.005853f
C473 B.n428 VSUBS 0.005853f
C474 B.n429 VSUBS 0.005853f
C475 B.n430 VSUBS 0.013908f
C476 B.n431 VSUBS 0.014499f
C477 B.n432 VSUBS 0.014499f
C478 B.n433 VSUBS 0.005853f
C479 B.n434 VSUBS 0.005853f
C480 B.n435 VSUBS 0.005853f
C481 B.n436 VSUBS 0.005853f
C482 B.n437 VSUBS 0.005853f
C483 B.n438 VSUBS 0.005853f
C484 B.n439 VSUBS 0.005853f
C485 B.n440 VSUBS 0.005853f
C486 B.n441 VSUBS 0.005853f
C487 B.n442 VSUBS 0.005853f
C488 B.n443 VSUBS 0.005853f
C489 B.n444 VSUBS 0.005853f
C490 B.n445 VSUBS 0.005853f
C491 B.n446 VSUBS 0.005853f
C492 B.n447 VSUBS 0.005853f
C493 B.n448 VSUBS 0.005853f
C494 B.n449 VSUBS 0.005853f
C495 B.n450 VSUBS 0.005853f
C496 B.n451 VSUBS 0.005853f
C497 B.n452 VSUBS 0.005853f
C498 B.n453 VSUBS 0.005853f
C499 B.n454 VSUBS 0.005853f
C500 B.n455 VSUBS 0.005853f
C501 B.n456 VSUBS 0.005853f
C502 B.n457 VSUBS 0.005853f
C503 B.n458 VSUBS 0.005853f
C504 B.n459 VSUBS 0.005853f
C505 B.n460 VSUBS 0.005853f
C506 B.n461 VSUBS 0.005853f
C507 B.n462 VSUBS 0.005853f
C508 B.n463 VSUBS 0.005853f
C509 B.n464 VSUBS 0.005853f
C510 B.n465 VSUBS 0.005853f
C511 B.n466 VSUBS 0.005853f
C512 B.n467 VSUBS 0.005853f
C513 B.n468 VSUBS 0.005853f
C514 B.n469 VSUBS 0.005853f
C515 B.n470 VSUBS 0.005853f
C516 B.n471 VSUBS 0.005853f
C517 B.n472 VSUBS 0.005853f
C518 B.n473 VSUBS 0.005853f
C519 B.n474 VSUBS 0.005853f
C520 B.n475 VSUBS 0.005853f
C521 B.n476 VSUBS 0.005853f
C522 B.n477 VSUBS 0.005853f
C523 B.n478 VSUBS 0.005853f
C524 B.n479 VSUBS 0.005853f
C525 B.n480 VSUBS 0.005853f
C526 B.n481 VSUBS 0.005853f
C527 B.n482 VSUBS 0.005853f
C528 B.n483 VSUBS 0.005853f
C529 B.n484 VSUBS 0.005853f
C530 B.n485 VSUBS 0.005853f
C531 B.n486 VSUBS 0.005853f
C532 B.n487 VSUBS 0.005853f
C533 B.n488 VSUBS 0.005853f
C534 B.n489 VSUBS 0.005853f
C535 B.n490 VSUBS 0.005853f
C536 B.n491 VSUBS 0.005853f
C537 B.n492 VSUBS 0.005853f
C538 B.n493 VSUBS 0.005853f
C539 B.n494 VSUBS 0.005853f
C540 B.n495 VSUBS 0.005853f
C541 B.n496 VSUBS 0.005853f
C542 B.n497 VSUBS 0.005853f
C543 B.n498 VSUBS 0.005853f
C544 B.n499 VSUBS 0.005853f
C545 B.n500 VSUBS 0.005509f
C546 B.n501 VSUBS 0.005853f
C547 B.n502 VSUBS 0.005853f
C548 B.n503 VSUBS 0.005853f
C549 B.n504 VSUBS 0.005853f
C550 B.n505 VSUBS 0.005853f
C551 B.n506 VSUBS 0.005853f
C552 B.n507 VSUBS 0.005853f
C553 B.n508 VSUBS 0.005853f
C554 B.n509 VSUBS 0.005853f
C555 B.n510 VSUBS 0.005853f
C556 B.n511 VSUBS 0.005853f
C557 B.n512 VSUBS 0.005853f
C558 B.n513 VSUBS 0.005853f
C559 B.n514 VSUBS 0.005853f
C560 B.n515 VSUBS 0.005853f
C561 B.n516 VSUBS 0.003271f
C562 B.n517 VSUBS 0.013562f
C563 B.n518 VSUBS 0.005509f
C564 B.n519 VSUBS 0.005853f
C565 B.n520 VSUBS 0.005853f
C566 B.n521 VSUBS 0.005853f
C567 B.n522 VSUBS 0.005853f
C568 B.n523 VSUBS 0.005853f
C569 B.n524 VSUBS 0.005853f
C570 B.n525 VSUBS 0.005853f
C571 B.n526 VSUBS 0.005853f
C572 B.n527 VSUBS 0.005853f
C573 B.n528 VSUBS 0.005853f
C574 B.n529 VSUBS 0.005853f
C575 B.n530 VSUBS 0.005853f
C576 B.n531 VSUBS 0.005853f
C577 B.n532 VSUBS 0.005853f
C578 B.n533 VSUBS 0.005853f
C579 B.n534 VSUBS 0.005853f
C580 B.n535 VSUBS 0.005853f
C581 B.n536 VSUBS 0.005853f
C582 B.n537 VSUBS 0.005853f
C583 B.n538 VSUBS 0.005853f
C584 B.n539 VSUBS 0.005853f
C585 B.n540 VSUBS 0.005853f
C586 B.n541 VSUBS 0.005853f
C587 B.n542 VSUBS 0.005853f
C588 B.n543 VSUBS 0.005853f
C589 B.n544 VSUBS 0.005853f
C590 B.n545 VSUBS 0.005853f
C591 B.n546 VSUBS 0.005853f
C592 B.n547 VSUBS 0.005853f
C593 B.n548 VSUBS 0.005853f
C594 B.n549 VSUBS 0.005853f
C595 B.n550 VSUBS 0.005853f
C596 B.n551 VSUBS 0.005853f
C597 B.n552 VSUBS 0.005853f
C598 B.n553 VSUBS 0.005853f
C599 B.n554 VSUBS 0.005853f
C600 B.n555 VSUBS 0.005853f
C601 B.n556 VSUBS 0.005853f
C602 B.n557 VSUBS 0.005853f
C603 B.n558 VSUBS 0.005853f
C604 B.n559 VSUBS 0.005853f
C605 B.n560 VSUBS 0.005853f
C606 B.n561 VSUBS 0.005853f
C607 B.n562 VSUBS 0.005853f
C608 B.n563 VSUBS 0.005853f
C609 B.n564 VSUBS 0.005853f
C610 B.n565 VSUBS 0.005853f
C611 B.n566 VSUBS 0.005853f
C612 B.n567 VSUBS 0.005853f
C613 B.n568 VSUBS 0.005853f
C614 B.n569 VSUBS 0.005853f
C615 B.n570 VSUBS 0.005853f
C616 B.n571 VSUBS 0.005853f
C617 B.n572 VSUBS 0.005853f
C618 B.n573 VSUBS 0.005853f
C619 B.n574 VSUBS 0.005853f
C620 B.n575 VSUBS 0.005853f
C621 B.n576 VSUBS 0.005853f
C622 B.n577 VSUBS 0.005853f
C623 B.n578 VSUBS 0.005853f
C624 B.n579 VSUBS 0.005853f
C625 B.n580 VSUBS 0.005853f
C626 B.n581 VSUBS 0.005853f
C627 B.n582 VSUBS 0.005853f
C628 B.n583 VSUBS 0.005853f
C629 B.n584 VSUBS 0.005853f
C630 B.n585 VSUBS 0.005853f
C631 B.n586 VSUBS 0.005853f
C632 B.n587 VSUBS 0.014499f
C633 B.n588 VSUBS 0.013908f
C634 B.n589 VSUBS 0.013908f
C635 B.n590 VSUBS 0.005853f
C636 B.n591 VSUBS 0.005853f
C637 B.n592 VSUBS 0.005853f
C638 B.n593 VSUBS 0.005853f
C639 B.n594 VSUBS 0.005853f
C640 B.n595 VSUBS 0.005853f
C641 B.n596 VSUBS 0.005853f
C642 B.n597 VSUBS 0.005853f
C643 B.n598 VSUBS 0.005853f
C644 B.n599 VSUBS 0.005853f
C645 B.n600 VSUBS 0.005853f
C646 B.n601 VSUBS 0.005853f
C647 B.n602 VSUBS 0.005853f
C648 B.n603 VSUBS 0.005853f
C649 B.n604 VSUBS 0.005853f
C650 B.n605 VSUBS 0.005853f
C651 B.n606 VSUBS 0.005853f
C652 B.n607 VSUBS 0.005853f
C653 B.n608 VSUBS 0.005853f
C654 B.n609 VSUBS 0.005853f
C655 B.n610 VSUBS 0.005853f
C656 B.n611 VSUBS 0.005853f
C657 B.n612 VSUBS 0.005853f
C658 B.n613 VSUBS 0.005853f
C659 B.n614 VSUBS 0.005853f
C660 B.n615 VSUBS 0.005853f
C661 B.n616 VSUBS 0.005853f
C662 B.n617 VSUBS 0.005853f
C663 B.n618 VSUBS 0.005853f
C664 B.n619 VSUBS 0.005853f
C665 B.n620 VSUBS 0.005853f
C666 B.n621 VSUBS 0.005853f
C667 B.n622 VSUBS 0.005853f
C668 B.n623 VSUBS 0.007638f
C669 B.n624 VSUBS 0.008137f
C670 B.n625 VSUBS 0.016181f
C671 VDD1.t0 VSUBS 2.32526f
C672 VDD1.t1 VSUBS 2.97059f
C673 VTAIL.t3 VSUBS 3.11175f
C674 VTAIL.n0 VSUBS 2.84948f
C675 VTAIL.t1 VSUBS 3.11177f
C676 VTAIL.n1 VSUBS 2.89992f
C677 VTAIL.t2 VSUBS 3.11177f
C678 VTAIL.n2 VSUBS 2.67654f
C679 VTAIL.t0 VSUBS 3.11175f
C680 VTAIL.n3 VSUBS 2.57184f
C681 VP.t1 VSUBS 4.841721f
C682 VP.t0 VSUBS 4.20095f
C683 VP.n0 VSUBS 5.766f
.ends

