* NGSPICE file created from diff_pair_sample_0552.ext - technology: sky130A

.subckt diff_pair_sample_0552 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=0.585 pd=3.78 as=0.2475 ps=1.83 w=1.5 l=0.27
X1 VDD1.t5 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.585 ps=3.78 w=1.5 l=0.27
X2 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=0.585 pd=3.78 as=0 ps=0 w=1.5 l=0.27
X3 VTAIL.t4 VP.t1 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.2475 ps=1.83 w=1.5 l=0.27
X4 VTAIL.t5 VP.t2 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.2475 ps=1.83 w=1.5 l=0.27
X5 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=0.585 pd=3.78 as=0 ps=0 w=1.5 l=0.27
X6 VDD1.t2 VP.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.585 pd=3.78 as=0.2475 ps=1.83 w=1.5 l=0.27
X7 VDD1.t1 VP.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.585 ps=3.78 w=1.5 l=0.27
X8 VDD2.t4 VN.t1 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.585 ps=3.78 w=1.5 l=0.27
X9 VTAIL.t9 VN.t2 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.2475 ps=1.83 w=1.5 l=0.27
X10 VTAIL.t7 VN.t3 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.2475 ps=1.83 w=1.5 l=0.27
X11 VDD2.t1 VN.t4 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.585 pd=3.78 as=0.2475 ps=1.83 w=1.5 l=0.27
X12 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=0.585 pd=3.78 as=0 ps=0 w=1.5 l=0.27
X13 VDD1.t0 VP.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.585 pd=3.78 as=0.2475 ps=1.83 w=1.5 l=0.27
X14 VDD2.t0 VN.t5 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.585 ps=3.78 w=1.5 l=0.27
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.585 pd=3.78 as=0 ps=0 w=1.5 l=0.27
R0 VN.n2 VN.t5 301.048
R1 VN.n0 VN.t4 301.048
R2 VN.n6 VN.t0 301.048
R3 VN.n4 VN.t1 301.048
R4 VN.n1 VN.t2 249.927
R5 VN.n5 VN.t3 249.927
R6 VN.n7 VN.n4 161.489
R7 VN.n3 VN.n0 161.489
R8 VN.n3 VN.n2 161.3
R9 VN.n7 VN.n6 161.3
R10 VN.n1 VN.n0 36.5157
R11 VN.n2 VN.n1 36.5157
R12 VN.n6 VN.n5 36.5157
R13 VN.n5 VN.n4 36.5157
R14 VN VN.n7 32.0782
R15 VN VN.n3 0.0516364
R16 VTAIL.n7 VTAIL.t10 114.085
R17 VTAIL.n11 VTAIL.t8 114.085
R18 VTAIL.n2 VTAIL.t3 114.085
R19 VTAIL.n10 VTAIL.t1 114.085
R20 VTAIL.n9 VTAIL.n8 100.885
R21 VTAIL.n6 VTAIL.n5 100.885
R22 VTAIL.n1 VTAIL.n0 100.885
R23 VTAIL.n4 VTAIL.n3 100.885
R24 VTAIL.n6 VTAIL.n4 14.6945
R25 VTAIL.n11 VTAIL.n10 14.1772
R26 VTAIL.n0 VTAIL.t6 13.2005
R27 VTAIL.n0 VTAIL.t9 13.2005
R28 VTAIL.n3 VTAIL.t2 13.2005
R29 VTAIL.n3 VTAIL.t5 13.2005
R30 VTAIL.n8 VTAIL.t0 13.2005
R31 VTAIL.n8 VTAIL.t4 13.2005
R32 VTAIL.n5 VTAIL.t11 13.2005
R33 VTAIL.n5 VTAIL.t7 13.2005
R34 VTAIL.n9 VTAIL.n7 0.728948
R35 VTAIL.n2 VTAIL.n1 0.728948
R36 VTAIL.n7 VTAIL.n6 0.517741
R37 VTAIL.n10 VTAIL.n9 0.517741
R38 VTAIL.n4 VTAIL.n2 0.517741
R39 VTAIL VTAIL.n11 0.330241
R40 VTAIL VTAIL.n1 0.188
R41 VDD2.n1 VDD2.t1 131.096
R42 VDD2.n2 VDD2.t5 130.764
R43 VDD2.n1 VDD2.n0 117.638
R44 VDD2 VDD2.n3 117.635
R45 VDD2.n2 VDD2.n1 26.6894
R46 VDD2.n3 VDD2.t2 13.2005
R47 VDD2.n3 VDD2.t4 13.2005
R48 VDD2.n0 VDD2.t3 13.2005
R49 VDD2.n0 VDD2.t0 13.2005
R50 VDD2 VDD2.n2 0.446621
R51 B.n286 B.n285 585
R52 B.n287 B.n286 585
R53 B.n109 B.n47 585
R54 B.n108 B.n107 585
R55 B.n106 B.n105 585
R56 B.n104 B.n103 585
R57 B.n102 B.n101 585
R58 B.n100 B.n99 585
R59 B.n98 B.n97 585
R60 B.n96 B.n95 585
R61 B.n94 B.n93 585
R62 B.n92 B.n91 585
R63 B.n90 B.n89 585
R64 B.n88 B.n87 585
R65 B.n86 B.n85 585
R66 B.n84 B.n83 585
R67 B.n82 B.n81 585
R68 B.n80 B.n79 585
R69 B.n78 B.n77 585
R70 B.n76 B.n75 585
R71 B.n74 B.n73 585
R72 B.n71 B.n70 585
R73 B.n69 B.n68 585
R74 B.n67 B.n66 585
R75 B.n65 B.n64 585
R76 B.n63 B.n62 585
R77 B.n61 B.n60 585
R78 B.n59 B.n58 585
R79 B.n57 B.n56 585
R80 B.n55 B.n54 585
R81 B.n32 B.n31 585
R82 B.n290 B.n289 585
R83 B.n284 B.n48 585
R84 B.n48 B.n29 585
R85 B.n283 B.n28 585
R86 B.n294 B.n28 585
R87 B.n282 B.n27 585
R88 B.n295 B.n27 585
R89 B.n281 B.n26 585
R90 B.n296 B.n26 585
R91 B.n280 B.n279 585
R92 B.n279 B.n25 585
R93 B.n278 B.n21 585
R94 B.n302 B.n21 585
R95 B.n277 B.n20 585
R96 B.n303 B.n20 585
R97 B.n276 B.n19 585
R98 B.n304 B.n19 585
R99 B.n275 B.n274 585
R100 B.n274 B.n18 585
R101 B.n273 B.n14 585
R102 B.n310 B.n14 585
R103 B.n272 B.n13 585
R104 B.n311 B.n13 585
R105 B.n271 B.n12 585
R106 B.n312 B.n12 585
R107 B.n270 B.n269 585
R108 B.n269 B.n11 585
R109 B.n268 B.n7 585
R110 B.n318 B.n7 585
R111 B.n267 B.n6 585
R112 B.n319 B.n6 585
R113 B.n266 B.n5 585
R114 B.n320 B.n5 585
R115 B.n265 B.n264 585
R116 B.n264 B.n4 585
R117 B.n263 B.n110 585
R118 B.n263 B.n262 585
R119 B.n252 B.n111 585
R120 B.n255 B.n111 585
R121 B.n254 B.n253 585
R122 B.n256 B.n254 585
R123 B.n251 B.n115 585
R124 B.n118 B.n115 585
R125 B.n250 B.n249 585
R126 B.n249 B.n248 585
R127 B.n117 B.n116 585
R128 B.n241 B.n117 585
R129 B.n240 B.n239 585
R130 B.n242 B.n240 585
R131 B.n238 B.n123 585
R132 B.n123 B.n122 585
R133 B.n237 B.n236 585
R134 B.n236 B.n235 585
R135 B.n125 B.n124 585
R136 B.n228 B.n125 585
R137 B.n227 B.n226 585
R138 B.n229 B.n227 585
R139 B.n225 B.n130 585
R140 B.n130 B.n129 585
R141 B.n224 B.n223 585
R142 B.n223 B.n222 585
R143 B.n132 B.n131 585
R144 B.n133 B.n132 585
R145 B.n218 B.n217 585
R146 B.n136 B.n135 585
R147 B.n214 B.n213 585
R148 B.n215 B.n214 585
R149 B.n212 B.n151 585
R150 B.n211 B.n210 585
R151 B.n209 B.n208 585
R152 B.n207 B.n206 585
R153 B.n205 B.n204 585
R154 B.n203 B.n202 585
R155 B.n201 B.n200 585
R156 B.n199 B.n198 585
R157 B.n197 B.n196 585
R158 B.n195 B.n194 585
R159 B.n193 B.n192 585
R160 B.n191 B.n190 585
R161 B.n189 B.n188 585
R162 B.n187 B.n186 585
R163 B.n185 B.n184 585
R164 B.n183 B.n182 585
R165 B.n181 B.n180 585
R166 B.n178 B.n177 585
R167 B.n176 B.n175 585
R168 B.n174 B.n173 585
R169 B.n172 B.n171 585
R170 B.n170 B.n169 585
R171 B.n168 B.n167 585
R172 B.n166 B.n165 585
R173 B.n164 B.n163 585
R174 B.n162 B.n161 585
R175 B.n160 B.n159 585
R176 B.n158 B.n157 585
R177 B.n219 B.n134 585
R178 B.n134 B.n133 585
R179 B.n221 B.n220 585
R180 B.n222 B.n221 585
R181 B.n128 B.n127 585
R182 B.n129 B.n128 585
R183 B.n231 B.n230 585
R184 B.n230 B.n229 585
R185 B.n232 B.n126 585
R186 B.n228 B.n126 585
R187 B.n234 B.n233 585
R188 B.n235 B.n234 585
R189 B.n121 B.n120 585
R190 B.n122 B.n121 585
R191 B.n244 B.n243 585
R192 B.n243 B.n242 585
R193 B.n245 B.n119 585
R194 B.n241 B.n119 585
R195 B.n247 B.n246 585
R196 B.n248 B.n247 585
R197 B.n114 B.n113 585
R198 B.n118 B.n114 585
R199 B.n258 B.n257 585
R200 B.n257 B.n256 585
R201 B.n259 B.n112 585
R202 B.n255 B.n112 585
R203 B.n261 B.n260 585
R204 B.n262 B.n261 585
R205 B.n2 B.n0 585
R206 B.n4 B.n2 585
R207 B.n3 B.n1 585
R208 B.n319 B.n3 585
R209 B.n317 B.n316 585
R210 B.n318 B.n317 585
R211 B.n315 B.n8 585
R212 B.n11 B.n8 585
R213 B.n314 B.n313 585
R214 B.n313 B.n312 585
R215 B.n10 B.n9 585
R216 B.n311 B.n10 585
R217 B.n309 B.n308 585
R218 B.n310 B.n309 585
R219 B.n307 B.n15 585
R220 B.n18 B.n15 585
R221 B.n306 B.n305 585
R222 B.n305 B.n304 585
R223 B.n17 B.n16 585
R224 B.n303 B.n17 585
R225 B.n301 B.n300 585
R226 B.n302 B.n301 585
R227 B.n299 B.n22 585
R228 B.n25 B.n22 585
R229 B.n298 B.n297 585
R230 B.n297 B.n296 585
R231 B.n24 B.n23 585
R232 B.n295 B.n24 585
R233 B.n293 B.n292 585
R234 B.n294 B.n293 585
R235 B.n291 B.n30 585
R236 B.n30 B.n29 585
R237 B.n322 B.n321 585
R238 B.n321 B.n320 585
R239 B.n217 B.n134 530.939
R240 B.n289 B.n30 530.939
R241 B.n157 B.n132 530.939
R242 B.n286 B.n48 530.939
R243 B.n155 B.t10 354.618
R244 B.n152 B.t6 354.618
R245 B.n52 B.t17 354.618
R246 B.n49 B.t13 354.618
R247 B.n287 B.n46 256.663
R248 B.n287 B.n45 256.663
R249 B.n287 B.n44 256.663
R250 B.n287 B.n43 256.663
R251 B.n287 B.n42 256.663
R252 B.n287 B.n41 256.663
R253 B.n287 B.n40 256.663
R254 B.n287 B.n39 256.663
R255 B.n287 B.n38 256.663
R256 B.n287 B.n37 256.663
R257 B.n287 B.n36 256.663
R258 B.n287 B.n35 256.663
R259 B.n287 B.n34 256.663
R260 B.n287 B.n33 256.663
R261 B.n288 B.n287 256.663
R262 B.n216 B.n215 256.663
R263 B.n215 B.n137 256.663
R264 B.n215 B.n138 256.663
R265 B.n215 B.n139 256.663
R266 B.n215 B.n140 256.663
R267 B.n215 B.n141 256.663
R268 B.n215 B.n142 256.663
R269 B.n215 B.n143 256.663
R270 B.n215 B.n144 256.663
R271 B.n215 B.n145 256.663
R272 B.n215 B.n146 256.663
R273 B.n215 B.n147 256.663
R274 B.n215 B.n148 256.663
R275 B.n215 B.n149 256.663
R276 B.n215 B.n150 256.663
R277 B.n215 B.n133 219.189
R278 B.n287 B.n29 219.189
R279 B.n221 B.n134 163.367
R280 B.n221 B.n128 163.367
R281 B.n230 B.n128 163.367
R282 B.n230 B.n126 163.367
R283 B.n234 B.n126 163.367
R284 B.n234 B.n121 163.367
R285 B.n243 B.n121 163.367
R286 B.n243 B.n119 163.367
R287 B.n247 B.n119 163.367
R288 B.n247 B.n114 163.367
R289 B.n257 B.n114 163.367
R290 B.n257 B.n112 163.367
R291 B.n261 B.n112 163.367
R292 B.n261 B.n2 163.367
R293 B.n321 B.n2 163.367
R294 B.n321 B.n3 163.367
R295 B.n317 B.n3 163.367
R296 B.n317 B.n8 163.367
R297 B.n313 B.n8 163.367
R298 B.n313 B.n10 163.367
R299 B.n309 B.n10 163.367
R300 B.n309 B.n15 163.367
R301 B.n305 B.n15 163.367
R302 B.n305 B.n17 163.367
R303 B.n301 B.n17 163.367
R304 B.n301 B.n22 163.367
R305 B.n297 B.n22 163.367
R306 B.n297 B.n24 163.367
R307 B.n293 B.n24 163.367
R308 B.n293 B.n30 163.367
R309 B.n214 B.n136 163.367
R310 B.n214 B.n151 163.367
R311 B.n210 B.n209 163.367
R312 B.n206 B.n205 163.367
R313 B.n202 B.n201 163.367
R314 B.n198 B.n197 163.367
R315 B.n194 B.n193 163.367
R316 B.n190 B.n189 163.367
R317 B.n186 B.n185 163.367
R318 B.n182 B.n181 163.367
R319 B.n177 B.n176 163.367
R320 B.n173 B.n172 163.367
R321 B.n169 B.n168 163.367
R322 B.n165 B.n164 163.367
R323 B.n161 B.n160 163.367
R324 B.n223 B.n132 163.367
R325 B.n223 B.n130 163.367
R326 B.n227 B.n130 163.367
R327 B.n227 B.n125 163.367
R328 B.n236 B.n125 163.367
R329 B.n236 B.n123 163.367
R330 B.n240 B.n123 163.367
R331 B.n240 B.n117 163.367
R332 B.n249 B.n117 163.367
R333 B.n249 B.n115 163.367
R334 B.n254 B.n115 163.367
R335 B.n254 B.n111 163.367
R336 B.n263 B.n111 163.367
R337 B.n264 B.n263 163.367
R338 B.n264 B.n5 163.367
R339 B.n6 B.n5 163.367
R340 B.n7 B.n6 163.367
R341 B.n269 B.n7 163.367
R342 B.n269 B.n12 163.367
R343 B.n13 B.n12 163.367
R344 B.n14 B.n13 163.367
R345 B.n274 B.n14 163.367
R346 B.n274 B.n19 163.367
R347 B.n20 B.n19 163.367
R348 B.n21 B.n20 163.367
R349 B.n279 B.n21 163.367
R350 B.n279 B.n26 163.367
R351 B.n27 B.n26 163.367
R352 B.n28 B.n27 163.367
R353 B.n48 B.n28 163.367
R354 B.n54 B.n32 163.367
R355 B.n58 B.n57 163.367
R356 B.n62 B.n61 163.367
R357 B.n66 B.n65 163.367
R358 B.n70 B.n69 163.367
R359 B.n75 B.n74 163.367
R360 B.n79 B.n78 163.367
R361 B.n83 B.n82 163.367
R362 B.n87 B.n86 163.367
R363 B.n91 B.n90 163.367
R364 B.n95 B.n94 163.367
R365 B.n99 B.n98 163.367
R366 B.n103 B.n102 163.367
R367 B.n107 B.n106 163.367
R368 B.n286 B.n47 163.367
R369 B.n155 B.t12 118.975
R370 B.n49 B.t15 118.975
R371 B.n152 B.t9 118.975
R372 B.n52 B.t18 118.975
R373 B.n222 B.n133 110.406
R374 B.n222 B.n129 110.406
R375 B.n229 B.n129 110.406
R376 B.n229 B.n228 110.406
R377 B.n235 B.n122 110.406
R378 B.n242 B.n122 110.406
R379 B.n242 B.n241 110.406
R380 B.n248 B.n118 110.406
R381 B.n256 B.n255 110.406
R382 B.n262 B.n4 110.406
R383 B.n320 B.n4 110.406
R384 B.n320 B.n319 110.406
R385 B.n319 B.n318 110.406
R386 B.n312 B.n11 110.406
R387 B.n311 B.n310 110.406
R388 B.n304 B.n18 110.406
R389 B.n304 B.n303 110.406
R390 B.n303 B.n302 110.406
R391 B.n296 B.n25 110.406
R392 B.n296 B.n295 110.406
R393 B.n295 B.n294 110.406
R394 B.n294 B.n29 110.406
R395 B.n235 B.t7 108.782
R396 B.n241 B.t2 108.782
R397 B.n18 B.t1 108.782
R398 B.n302 B.t14 108.782
R399 B.n156 B.t11 107.34
R400 B.n50 B.t16 107.34
R401 B.n153 B.t8 107.338
R402 B.n53 B.t19 107.338
R403 B.n118 B.t5 82.8049
R404 B.t4 B.n311 82.8049
R405 B.n217 B.n216 71.676
R406 B.n151 B.n137 71.676
R407 B.n209 B.n138 71.676
R408 B.n205 B.n139 71.676
R409 B.n201 B.n140 71.676
R410 B.n197 B.n141 71.676
R411 B.n193 B.n142 71.676
R412 B.n189 B.n143 71.676
R413 B.n185 B.n144 71.676
R414 B.n181 B.n145 71.676
R415 B.n176 B.n146 71.676
R416 B.n172 B.n147 71.676
R417 B.n168 B.n148 71.676
R418 B.n164 B.n149 71.676
R419 B.n160 B.n150 71.676
R420 B.n289 B.n288 71.676
R421 B.n54 B.n33 71.676
R422 B.n58 B.n34 71.676
R423 B.n62 B.n35 71.676
R424 B.n66 B.n36 71.676
R425 B.n70 B.n37 71.676
R426 B.n75 B.n38 71.676
R427 B.n79 B.n39 71.676
R428 B.n83 B.n40 71.676
R429 B.n87 B.n41 71.676
R430 B.n91 B.n42 71.676
R431 B.n95 B.n43 71.676
R432 B.n99 B.n44 71.676
R433 B.n103 B.n45 71.676
R434 B.n107 B.n46 71.676
R435 B.n47 B.n46 71.676
R436 B.n106 B.n45 71.676
R437 B.n102 B.n44 71.676
R438 B.n98 B.n43 71.676
R439 B.n94 B.n42 71.676
R440 B.n90 B.n41 71.676
R441 B.n86 B.n40 71.676
R442 B.n82 B.n39 71.676
R443 B.n78 B.n38 71.676
R444 B.n74 B.n37 71.676
R445 B.n69 B.n36 71.676
R446 B.n65 B.n35 71.676
R447 B.n61 B.n34 71.676
R448 B.n57 B.n33 71.676
R449 B.n288 B.n32 71.676
R450 B.n216 B.n136 71.676
R451 B.n210 B.n137 71.676
R452 B.n206 B.n138 71.676
R453 B.n202 B.n139 71.676
R454 B.n198 B.n140 71.676
R455 B.n194 B.n141 71.676
R456 B.n190 B.n142 71.676
R457 B.n186 B.n143 71.676
R458 B.n182 B.n144 71.676
R459 B.n177 B.n145 71.676
R460 B.n173 B.n146 71.676
R461 B.n169 B.n147 71.676
R462 B.n165 B.n148 71.676
R463 B.n161 B.n149 71.676
R464 B.n157 B.n150 71.676
R465 B.n179 B.n156 59.5399
R466 B.n154 B.n153 59.5399
R467 B.n72 B.n53 59.5399
R468 B.n51 B.n50 59.5399
R469 B.n255 B.t3 56.8271
R470 B.n11 B.t0 56.8271
R471 B.n262 B.t3 53.5798
R472 B.n318 B.t0 53.5798
R473 B.n291 B.n290 34.4981
R474 B.n285 B.n284 34.4981
R475 B.n158 B.n131 34.4981
R476 B.n219 B.n218 34.4981
R477 B.n256 B.t5 27.602
R478 B.n312 B.t4 27.602
R479 B B.n322 18.0485
R480 B.n156 B.n155 11.6369
R481 B.n153 B.n152 11.6369
R482 B.n53 B.n52 11.6369
R483 B.n50 B.n49 11.6369
R484 B.n290 B.n31 10.6151
R485 B.n55 B.n31 10.6151
R486 B.n56 B.n55 10.6151
R487 B.n59 B.n56 10.6151
R488 B.n60 B.n59 10.6151
R489 B.n63 B.n60 10.6151
R490 B.n64 B.n63 10.6151
R491 B.n67 B.n64 10.6151
R492 B.n68 B.n67 10.6151
R493 B.n71 B.n68 10.6151
R494 B.n76 B.n73 10.6151
R495 B.n77 B.n76 10.6151
R496 B.n80 B.n77 10.6151
R497 B.n81 B.n80 10.6151
R498 B.n84 B.n81 10.6151
R499 B.n85 B.n84 10.6151
R500 B.n88 B.n85 10.6151
R501 B.n89 B.n88 10.6151
R502 B.n93 B.n92 10.6151
R503 B.n96 B.n93 10.6151
R504 B.n97 B.n96 10.6151
R505 B.n100 B.n97 10.6151
R506 B.n101 B.n100 10.6151
R507 B.n104 B.n101 10.6151
R508 B.n105 B.n104 10.6151
R509 B.n108 B.n105 10.6151
R510 B.n109 B.n108 10.6151
R511 B.n285 B.n109 10.6151
R512 B.n224 B.n131 10.6151
R513 B.n225 B.n224 10.6151
R514 B.n226 B.n225 10.6151
R515 B.n226 B.n124 10.6151
R516 B.n237 B.n124 10.6151
R517 B.n238 B.n237 10.6151
R518 B.n239 B.n238 10.6151
R519 B.n239 B.n116 10.6151
R520 B.n250 B.n116 10.6151
R521 B.n251 B.n250 10.6151
R522 B.n253 B.n251 10.6151
R523 B.n253 B.n252 10.6151
R524 B.n252 B.n110 10.6151
R525 B.n265 B.n110 10.6151
R526 B.n266 B.n265 10.6151
R527 B.n267 B.n266 10.6151
R528 B.n268 B.n267 10.6151
R529 B.n270 B.n268 10.6151
R530 B.n271 B.n270 10.6151
R531 B.n272 B.n271 10.6151
R532 B.n273 B.n272 10.6151
R533 B.n275 B.n273 10.6151
R534 B.n276 B.n275 10.6151
R535 B.n277 B.n276 10.6151
R536 B.n278 B.n277 10.6151
R537 B.n280 B.n278 10.6151
R538 B.n281 B.n280 10.6151
R539 B.n282 B.n281 10.6151
R540 B.n283 B.n282 10.6151
R541 B.n284 B.n283 10.6151
R542 B.n218 B.n135 10.6151
R543 B.n213 B.n135 10.6151
R544 B.n213 B.n212 10.6151
R545 B.n212 B.n211 10.6151
R546 B.n211 B.n208 10.6151
R547 B.n208 B.n207 10.6151
R548 B.n207 B.n204 10.6151
R549 B.n204 B.n203 10.6151
R550 B.n203 B.n200 10.6151
R551 B.n200 B.n199 10.6151
R552 B.n196 B.n195 10.6151
R553 B.n195 B.n192 10.6151
R554 B.n192 B.n191 10.6151
R555 B.n191 B.n188 10.6151
R556 B.n188 B.n187 10.6151
R557 B.n187 B.n184 10.6151
R558 B.n184 B.n183 10.6151
R559 B.n183 B.n180 10.6151
R560 B.n178 B.n175 10.6151
R561 B.n175 B.n174 10.6151
R562 B.n174 B.n171 10.6151
R563 B.n171 B.n170 10.6151
R564 B.n170 B.n167 10.6151
R565 B.n167 B.n166 10.6151
R566 B.n166 B.n163 10.6151
R567 B.n163 B.n162 10.6151
R568 B.n162 B.n159 10.6151
R569 B.n159 B.n158 10.6151
R570 B.n220 B.n219 10.6151
R571 B.n220 B.n127 10.6151
R572 B.n231 B.n127 10.6151
R573 B.n232 B.n231 10.6151
R574 B.n233 B.n232 10.6151
R575 B.n233 B.n120 10.6151
R576 B.n244 B.n120 10.6151
R577 B.n245 B.n244 10.6151
R578 B.n246 B.n245 10.6151
R579 B.n246 B.n113 10.6151
R580 B.n258 B.n113 10.6151
R581 B.n259 B.n258 10.6151
R582 B.n260 B.n259 10.6151
R583 B.n260 B.n0 10.6151
R584 B.n316 B.n1 10.6151
R585 B.n316 B.n315 10.6151
R586 B.n315 B.n314 10.6151
R587 B.n314 B.n9 10.6151
R588 B.n308 B.n9 10.6151
R589 B.n308 B.n307 10.6151
R590 B.n307 B.n306 10.6151
R591 B.n306 B.n16 10.6151
R592 B.n300 B.n16 10.6151
R593 B.n300 B.n299 10.6151
R594 B.n299 B.n298 10.6151
R595 B.n298 B.n23 10.6151
R596 B.n292 B.n23 10.6151
R597 B.n292 B.n291 10.6151
R598 B.n73 B.n72 6.5566
R599 B.n89 B.n51 6.5566
R600 B.n196 B.n154 6.5566
R601 B.n180 B.n179 6.5566
R602 B.n72 B.n71 4.05904
R603 B.n92 B.n51 4.05904
R604 B.n199 B.n154 4.05904
R605 B.n179 B.n178 4.05904
R606 B.n322 B.n0 2.81026
R607 B.n322 B.n1 2.81026
R608 B.n228 B.t7 1.62412
R609 B.n248 B.t2 1.62412
R610 B.n310 B.t1 1.62412
R611 B.n25 B.t14 1.62412
R612 VP.n7 VP.t0 301.048
R613 VP.n5 VP.t3 301.048
R614 VP.n0 VP.t5 301.048
R615 VP.n2 VP.t4 301.048
R616 VP.n6 VP.t2 249.927
R617 VP.n1 VP.t1 249.927
R618 VP.n3 VP.n0 161.489
R619 VP.n8 VP.n7 161.3
R620 VP.n3 VP.n2 161.3
R621 VP.n5 VP.n4 161.3
R622 VP.n6 VP.n5 36.5157
R623 VP.n7 VP.n6 36.5157
R624 VP.n1 VP.n0 36.5157
R625 VP.n2 VP.n1 36.5157
R626 VP.n4 VP.n3 31.6975
R627 VP.n8 VP.n4 0.189894
R628 VP VP.n8 0.0516364
R629 VDD1 VDD1.t0 131.21
R630 VDD1.n1 VDD1.t2 131.096
R631 VDD1.n1 VDD1.n0 117.638
R632 VDD1.n3 VDD1.n2 117.564
R633 VDD1.n3 VDD1.n1 27.5311
R634 VDD1.n2 VDD1.t4 13.2005
R635 VDD1.n2 VDD1.t1 13.2005
R636 VDD1.n0 VDD1.t3 13.2005
R637 VDD1.n0 VDD1.t5 13.2005
R638 VDD1 VDD1.n3 0.0716207
C0 VDD2 VN 0.589163f
C1 VDD2 VTAIL 3.23542f
C2 VN VTAIL 0.660793f
C3 VDD2 VDD1 0.555588f
C4 VDD1 VN 0.154746f
C5 VDD1 VTAIL 3.19863f
C6 VDD2 VP 0.267485f
C7 VP VN 2.72194f
C8 VP VTAIL 0.674983f
C9 VP VDD1 0.700363f
C10 VDD2 B 2.177107f
C11 VDD1 B 2.330162f
C12 VTAIL B 2.089009f
C13 VN B 4.69216f
C14 VP B 3.599071f
C15 VDD1.t0 B 0.201435f
C16 VDD1.t2 B 0.20124f
C17 VDD1.t3 B 0.025588f
C18 VDD1.t5 B 0.025588f
C19 VDD1.n0 B 0.150739f
C20 VDD1.n1 B 1.07527f
C21 VDD1.t4 B 0.025588f
C22 VDD1.t1 B 0.025588f
C23 VDD1.n2 B 0.15061f
C24 VDD1.n3 B 1.0759f
C25 VP.t5 B 0.055679f
C26 VP.n0 B 0.05181f
C27 VP.t1 B 0.048304f
C28 VP.n1 B 0.040477f
C29 VP.t4 B 0.055679f
C30 VP.n2 B 0.05175f
C31 VP.n3 B 1.02361f
C32 VP.n4 B 1.01759f
C33 VP.t2 B 0.048304f
C34 VP.t3 B 0.055679f
C35 VP.n5 B 0.05175f
C36 VP.n6 B 0.040477f
C37 VP.t0 B 0.055679f
C38 VP.n7 B 0.05175f
C39 VP.n8 B 0.03092f
C40 VDD2.t1 B 0.206382f
C41 VDD2.t3 B 0.026242f
C42 VDD2.t0 B 0.026242f
C43 VDD2.n0 B 0.154591f
C44 VDD2.n1 B 1.04621f
C45 VDD2.t5 B 0.20586f
C46 VDD2.n2 B 1.08818f
C47 VDD2.t2 B 0.026242f
C48 VDD2.t4 B 0.026242f
C49 VDD2.n3 B 0.154581f
C50 VTAIL.t6 B 0.03359f
C51 VTAIL.t9 B 0.03359f
C52 VTAIL.n0 B 0.166528f
C53 VTAIL.n1 B 0.270305f
C54 VTAIL.t3 B 0.232155f
C55 VTAIL.n2 B 0.326395f
C56 VTAIL.t2 B 0.03359f
C57 VTAIL.t5 B 0.03359f
C58 VTAIL.n3 B 0.166528f
C59 VTAIL.n4 B 0.831359f
C60 VTAIL.t11 B 0.03359f
C61 VTAIL.t7 B 0.03359f
C62 VTAIL.n5 B 0.166528f
C63 VTAIL.n6 B 0.831358f
C64 VTAIL.t10 B 0.232155f
C65 VTAIL.n7 B 0.326394f
C66 VTAIL.t0 B 0.03359f
C67 VTAIL.t4 B 0.03359f
C68 VTAIL.n8 B 0.166528f
C69 VTAIL.n9 B 0.300413f
C70 VTAIL.t1 B 0.232155f
C71 VTAIL.n10 B 0.81011f
C72 VTAIL.t8 B 0.232155f
C73 VTAIL.n11 B 0.79299f
C74 VN.t4 B 0.054546f
C75 VN.n0 B 0.050756f
C76 VN.t2 B 0.047321f
C77 VN.n1 B 0.039653f
C78 VN.t5 B 0.054546f
C79 VN.n2 B 0.050697f
C80 VN.n3 B 0.080645f
C81 VN.t1 B 0.054546f
C82 VN.n4 B 0.050756f
C83 VN.t0 B 0.054546f
C84 VN.t3 B 0.047321f
C85 VN.n5 B 0.039653f
C86 VN.n6 B 0.050697f
C87 VN.n7 B 1.02897f
.ends

