* NGSPICE file created from diff_pair_sample_0632.ext - technology: sky130A

.subckt diff_pair_sample_0632 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=1.55595 pd=9.76 as=3.6777 ps=19.64 w=9.43 l=1.42
X1 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=3.6777 pd=19.64 as=0 ps=0 w=9.43 l=1.42
X2 VTAIL.t6 VN.t1 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.55595 pd=9.76 as=1.55595 ps=9.76 w=9.43 l=1.42
X3 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=3.6777 pd=19.64 as=0 ps=0 w=9.43 l=1.42
X4 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.6777 pd=19.64 as=0 ps=0 w=9.43 l=1.42
X5 VDD1.t5 VP.t0 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=1.55595 pd=9.76 as=3.6777 ps=19.64 w=9.43 l=1.42
X6 VTAIL.t9 VN.t2 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.55595 pd=9.76 as=1.55595 ps=9.76 w=9.43 l=1.42
X7 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.6777 pd=19.64 as=0 ps=0 w=9.43 l=1.42
X8 VDD2.t2 VN.t3 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=3.6777 pd=19.64 as=1.55595 ps=9.76 w=9.43 l=1.42
X9 VDD2.t1 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.55595 pd=9.76 as=3.6777 ps=19.64 w=9.43 l=1.42
X10 VDD1.t4 VP.t1 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=1.55595 pd=9.76 as=3.6777 ps=19.64 w=9.43 l=1.42
X11 VTAIL.t1 VP.t2 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.55595 pd=9.76 as=1.55595 ps=9.76 w=9.43 l=1.42
X12 VDD2.t0 VN.t5 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=3.6777 pd=19.64 as=1.55595 ps=9.76 w=9.43 l=1.42
X13 VDD1.t2 VP.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.6777 pd=19.64 as=1.55595 ps=9.76 w=9.43 l=1.42
X14 VDD1.t1 VP.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.6777 pd=19.64 as=1.55595 ps=9.76 w=9.43 l=1.42
X15 VTAIL.t0 VP.t5 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.55595 pd=9.76 as=1.55595 ps=9.76 w=9.43 l=1.42
R0 VN.n3 VN.t5 195.463
R1 VN.n13 VN.t4 195.463
R2 VN.n9 VN.n8 173.534
R3 VN.n19 VN.n18 173.534
R4 VN.n17 VN.n10 161.3
R5 VN.n16 VN.n15 161.3
R6 VN.n14 VN.n11 161.3
R7 VN.n7 VN.n0 161.3
R8 VN.n6 VN.n5 161.3
R9 VN.n4 VN.n1 161.3
R10 VN.n2 VN.t1 160.044
R11 VN.n8 VN.t0 160.044
R12 VN.n12 VN.t2 160.044
R13 VN.n18 VN.t3 160.044
R14 VN.n6 VN.n1 52.6342
R15 VN.n16 VN.n11 52.6342
R16 VN VN.n19 42.4229
R17 VN.n3 VN.n2 41.826
R18 VN.n13 VN.n12 41.826
R19 VN.n7 VN.n6 28.3526
R20 VN.n17 VN.n16 28.3526
R21 VN.n2 VN.n1 24.4675
R22 VN.n12 VN.n11 24.4675
R23 VN.n14 VN.n13 17.5327
R24 VN.n4 VN.n3 17.5327
R25 VN.n8 VN.n7 12.234
R26 VN.n18 VN.n17 12.234
R27 VN.n19 VN.n10 0.189894
R28 VN.n15 VN.n10 0.189894
R29 VN.n15 VN.n14 0.189894
R30 VN.n5 VN.n4 0.189894
R31 VN.n5 VN.n0 0.189894
R32 VN.n9 VN.n0 0.189894
R33 VN VN.n9 0.0516364
R34 VTAIL.n202 VTAIL.n158 289.615
R35 VTAIL.n46 VTAIL.n2 289.615
R36 VTAIL.n152 VTAIL.n108 289.615
R37 VTAIL.n100 VTAIL.n56 289.615
R38 VTAIL.n175 VTAIL.n174 185
R39 VTAIL.n177 VTAIL.n176 185
R40 VTAIL.n170 VTAIL.n169 185
R41 VTAIL.n183 VTAIL.n182 185
R42 VTAIL.n185 VTAIL.n184 185
R43 VTAIL.n166 VTAIL.n165 185
R44 VTAIL.n192 VTAIL.n191 185
R45 VTAIL.n193 VTAIL.n164 185
R46 VTAIL.n195 VTAIL.n194 185
R47 VTAIL.n162 VTAIL.n161 185
R48 VTAIL.n201 VTAIL.n200 185
R49 VTAIL.n203 VTAIL.n202 185
R50 VTAIL.n19 VTAIL.n18 185
R51 VTAIL.n21 VTAIL.n20 185
R52 VTAIL.n14 VTAIL.n13 185
R53 VTAIL.n27 VTAIL.n26 185
R54 VTAIL.n29 VTAIL.n28 185
R55 VTAIL.n10 VTAIL.n9 185
R56 VTAIL.n36 VTAIL.n35 185
R57 VTAIL.n37 VTAIL.n8 185
R58 VTAIL.n39 VTAIL.n38 185
R59 VTAIL.n6 VTAIL.n5 185
R60 VTAIL.n45 VTAIL.n44 185
R61 VTAIL.n47 VTAIL.n46 185
R62 VTAIL.n153 VTAIL.n152 185
R63 VTAIL.n151 VTAIL.n150 185
R64 VTAIL.n112 VTAIL.n111 185
R65 VTAIL.n116 VTAIL.n114 185
R66 VTAIL.n145 VTAIL.n144 185
R67 VTAIL.n143 VTAIL.n142 185
R68 VTAIL.n118 VTAIL.n117 185
R69 VTAIL.n137 VTAIL.n136 185
R70 VTAIL.n135 VTAIL.n134 185
R71 VTAIL.n122 VTAIL.n121 185
R72 VTAIL.n129 VTAIL.n128 185
R73 VTAIL.n127 VTAIL.n126 185
R74 VTAIL.n101 VTAIL.n100 185
R75 VTAIL.n99 VTAIL.n98 185
R76 VTAIL.n60 VTAIL.n59 185
R77 VTAIL.n64 VTAIL.n62 185
R78 VTAIL.n93 VTAIL.n92 185
R79 VTAIL.n91 VTAIL.n90 185
R80 VTAIL.n66 VTAIL.n65 185
R81 VTAIL.n85 VTAIL.n84 185
R82 VTAIL.n83 VTAIL.n82 185
R83 VTAIL.n70 VTAIL.n69 185
R84 VTAIL.n77 VTAIL.n76 185
R85 VTAIL.n75 VTAIL.n74 185
R86 VTAIL.n173 VTAIL.t8 149.524
R87 VTAIL.n17 VTAIL.t11 149.524
R88 VTAIL.n125 VTAIL.t10 149.524
R89 VTAIL.n73 VTAIL.t4 149.524
R90 VTAIL.n176 VTAIL.n175 104.615
R91 VTAIL.n176 VTAIL.n169 104.615
R92 VTAIL.n183 VTAIL.n169 104.615
R93 VTAIL.n184 VTAIL.n183 104.615
R94 VTAIL.n184 VTAIL.n165 104.615
R95 VTAIL.n192 VTAIL.n165 104.615
R96 VTAIL.n193 VTAIL.n192 104.615
R97 VTAIL.n194 VTAIL.n193 104.615
R98 VTAIL.n194 VTAIL.n161 104.615
R99 VTAIL.n201 VTAIL.n161 104.615
R100 VTAIL.n202 VTAIL.n201 104.615
R101 VTAIL.n20 VTAIL.n19 104.615
R102 VTAIL.n20 VTAIL.n13 104.615
R103 VTAIL.n27 VTAIL.n13 104.615
R104 VTAIL.n28 VTAIL.n27 104.615
R105 VTAIL.n28 VTAIL.n9 104.615
R106 VTAIL.n36 VTAIL.n9 104.615
R107 VTAIL.n37 VTAIL.n36 104.615
R108 VTAIL.n38 VTAIL.n37 104.615
R109 VTAIL.n38 VTAIL.n5 104.615
R110 VTAIL.n45 VTAIL.n5 104.615
R111 VTAIL.n46 VTAIL.n45 104.615
R112 VTAIL.n152 VTAIL.n151 104.615
R113 VTAIL.n151 VTAIL.n111 104.615
R114 VTAIL.n116 VTAIL.n111 104.615
R115 VTAIL.n144 VTAIL.n116 104.615
R116 VTAIL.n144 VTAIL.n143 104.615
R117 VTAIL.n143 VTAIL.n117 104.615
R118 VTAIL.n136 VTAIL.n117 104.615
R119 VTAIL.n136 VTAIL.n135 104.615
R120 VTAIL.n135 VTAIL.n121 104.615
R121 VTAIL.n128 VTAIL.n121 104.615
R122 VTAIL.n128 VTAIL.n127 104.615
R123 VTAIL.n100 VTAIL.n99 104.615
R124 VTAIL.n99 VTAIL.n59 104.615
R125 VTAIL.n64 VTAIL.n59 104.615
R126 VTAIL.n92 VTAIL.n64 104.615
R127 VTAIL.n92 VTAIL.n91 104.615
R128 VTAIL.n91 VTAIL.n65 104.615
R129 VTAIL.n84 VTAIL.n65 104.615
R130 VTAIL.n84 VTAIL.n83 104.615
R131 VTAIL.n83 VTAIL.n69 104.615
R132 VTAIL.n76 VTAIL.n69 104.615
R133 VTAIL.n76 VTAIL.n75 104.615
R134 VTAIL.n175 VTAIL.t8 52.3082
R135 VTAIL.n19 VTAIL.t11 52.3082
R136 VTAIL.n127 VTAIL.t10 52.3082
R137 VTAIL.n75 VTAIL.t4 52.3082
R138 VTAIL.n107 VTAIL.n106 50.0081
R139 VTAIL.n55 VTAIL.n54 50.0081
R140 VTAIL.n1 VTAIL.n0 50.0079
R141 VTAIL.n53 VTAIL.n52 50.0079
R142 VTAIL.n207 VTAIL.n206 35.8702
R143 VTAIL.n51 VTAIL.n50 35.8702
R144 VTAIL.n157 VTAIL.n156 35.8702
R145 VTAIL.n105 VTAIL.n104 35.8702
R146 VTAIL.n55 VTAIL.n53 23.5134
R147 VTAIL.n207 VTAIL.n157 22.0048
R148 VTAIL.n195 VTAIL.n162 13.1884
R149 VTAIL.n39 VTAIL.n6 13.1884
R150 VTAIL.n114 VTAIL.n112 13.1884
R151 VTAIL.n62 VTAIL.n60 13.1884
R152 VTAIL.n196 VTAIL.n164 12.8005
R153 VTAIL.n200 VTAIL.n199 12.8005
R154 VTAIL.n40 VTAIL.n8 12.8005
R155 VTAIL.n44 VTAIL.n43 12.8005
R156 VTAIL.n150 VTAIL.n149 12.8005
R157 VTAIL.n146 VTAIL.n145 12.8005
R158 VTAIL.n98 VTAIL.n97 12.8005
R159 VTAIL.n94 VTAIL.n93 12.8005
R160 VTAIL.n191 VTAIL.n190 12.0247
R161 VTAIL.n203 VTAIL.n160 12.0247
R162 VTAIL.n35 VTAIL.n34 12.0247
R163 VTAIL.n47 VTAIL.n4 12.0247
R164 VTAIL.n153 VTAIL.n110 12.0247
R165 VTAIL.n142 VTAIL.n115 12.0247
R166 VTAIL.n101 VTAIL.n58 12.0247
R167 VTAIL.n90 VTAIL.n63 12.0247
R168 VTAIL.n189 VTAIL.n166 11.249
R169 VTAIL.n204 VTAIL.n158 11.249
R170 VTAIL.n33 VTAIL.n10 11.249
R171 VTAIL.n48 VTAIL.n2 11.249
R172 VTAIL.n154 VTAIL.n108 11.249
R173 VTAIL.n141 VTAIL.n118 11.249
R174 VTAIL.n102 VTAIL.n56 11.249
R175 VTAIL.n89 VTAIL.n66 11.249
R176 VTAIL.n186 VTAIL.n185 10.4732
R177 VTAIL.n30 VTAIL.n29 10.4732
R178 VTAIL.n138 VTAIL.n137 10.4732
R179 VTAIL.n86 VTAIL.n85 10.4732
R180 VTAIL.n174 VTAIL.n173 10.2747
R181 VTAIL.n18 VTAIL.n17 10.2747
R182 VTAIL.n126 VTAIL.n125 10.2747
R183 VTAIL.n74 VTAIL.n73 10.2747
R184 VTAIL.n182 VTAIL.n168 9.69747
R185 VTAIL.n26 VTAIL.n12 9.69747
R186 VTAIL.n134 VTAIL.n120 9.69747
R187 VTAIL.n82 VTAIL.n68 9.69747
R188 VTAIL.n206 VTAIL.n205 9.45567
R189 VTAIL.n50 VTAIL.n49 9.45567
R190 VTAIL.n156 VTAIL.n155 9.45567
R191 VTAIL.n104 VTAIL.n103 9.45567
R192 VTAIL.n205 VTAIL.n204 9.3005
R193 VTAIL.n160 VTAIL.n159 9.3005
R194 VTAIL.n199 VTAIL.n198 9.3005
R195 VTAIL.n172 VTAIL.n171 9.3005
R196 VTAIL.n179 VTAIL.n178 9.3005
R197 VTAIL.n181 VTAIL.n180 9.3005
R198 VTAIL.n168 VTAIL.n167 9.3005
R199 VTAIL.n187 VTAIL.n186 9.3005
R200 VTAIL.n189 VTAIL.n188 9.3005
R201 VTAIL.n190 VTAIL.n163 9.3005
R202 VTAIL.n197 VTAIL.n196 9.3005
R203 VTAIL.n49 VTAIL.n48 9.3005
R204 VTAIL.n4 VTAIL.n3 9.3005
R205 VTAIL.n43 VTAIL.n42 9.3005
R206 VTAIL.n16 VTAIL.n15 9.3005
R207 VTAIL.n23 VTAIL.n22 9.3005
R208 VTAIL.n25 VTAIL.n24 9.3005
R209 VTAIL.n12 VTAIL.n11 9.3005
R210 VTAIL.n31 VTAIL.n30 9.3005
R211 VTAIL.n33 VTAIL.n32 9.3005
R212 VTAIL.n34 VTAIL.n7 9.3005
R213 VTAIL.n41 VTAIL.n40 9.3005
R214 VTAIL.n124 VTAIL.n123 9.3005
R215 VTAIL.n131 VTAIL.n130 9.3005
R216 VTAIL.n133 VTAIL.n132 9.3005
R217 VTAIL.n120 VTAIL.n119 9.3005
R218 VTAIL.n139 VTAIL.n138 9.3005
R219 VTAIL.n141 VTAIL.n140 9.3005
R220 VTAIL.n115 VTAIL.n113 9.3005
R221 VTAIL.n147 VTAIL.n146 9.3005
R222 VTAIL.n155 VTAIL.n154 9.3005
R223 VTAIL.n110 VTAIL.n109 9.3005
R224 VTAIL.n149 VTAIL.n148 9.3005
R225 VTAIL.n72 VTAIL.n71 9.3005
R226 VTAIL.n79 VTAIL.n78 9.3005
R227 VTAIL.n81 VTAIL.n80 9.3005
R228 VTAIL.n68 VTAIL.n67 9.3005
R229 VTAIL.n87 VTAIL.n86 9.3005
R230 VTAIL.n89 VTAIL.n88 9.3005
R231 VTAIL.n63 VTAIL.n61 9.3005
R232 VTAIL.n95 VTAIL.n94 9.3005
R233 VTAIL.n103 VTAIL.n102 9.3005
R234 VTAIL.n58 VTAIL.n57 9.3005
R235 VTAIL.n97 VTAIL.n96 9.3005
R236 VTAIL.n181 VTAIL.n170 8.92171
R237 VTAIL.n25 VTAIL.n14 8.92171
R238 VTAIL.n133 VTAIL.n122 8.92171
R239 VTAIL.n81 VTAIL.n70 8.92171
R240 VTAIL.n178 VTAIL.n177 8.14595
R241 VTAIL.n22 VTAIL.n21 8.14595
R242 VTAIL.n130 VTAIL.n129 8.14595
R243 VTAIL.n78 VTAIL.n77 8.14595
R244 VTAIL.n174 VTAIL.n172 7.3702
R245 VTAIL.n18 VTAIL.n16 7.3702
R246 VTAIL.n126 VTAIL.n124 7.3702
R247 VTAIL.n74 VTAIL.n72 7.3702
R248 VTAIL.n177 VTAIL.n172 5.81868
R249 VTAIL.n21 VTAIL.n16 5.81868
R250 VTAIL.n129 VTAIL.n124 5.81868
R251 VTAIL.n77 VTAIL.n72 5.81868
R252 VTAIL.n178 VTAIL.n170 5.04292
R253 VTAIL.n22 VTAIL.n14 5.04292
R254 VTAIL.n130 VTAIL.n122 5.04292
R255 VTAIL.n78 VTAIL.n70 5.04292
R256 VTAIL.n182 VTAIL.n181 4.26717
R257 VTAIL.n26 VTAIL.n25 4.26717
R258 VTAIL.n134 VTAIL.n133 4.26717
R259 VTAIL.n82 VTAIL.n81 4.26717
R260 VTAIL.n185 VTAIL.n168 3.49141
R261 VTAIL.n29 VTAIL.n12 3.49141
R262 VTAIL.n137 VTAIL.n120 3.49141
R263 VTAIL.n85 VTAIL.n68 3.49141
R264 VTAIL.n173 VTAIL.n171 2.84303
R265 VTAIL.n17 VTAIL.n15 2.84303
R266 VTAIL.n125 VTAIL.n123 2.84303
R267 VTAIL.n73 VTAIL.n71 2.84303
R268 VTAIL.n186 VTAIL.n166 2.71565
R269 VTAIL.n206 VTAIL.n158 2.71565
R270 VTAIL.n30 VTAIL.n10 2.71565
R271 VTAIL.n50 VTAIL.n2 2.71565
R272 VTAIL.n156 VTAIL.n108 2.71565
R273 VTAIL.n138 VTAIL.n118 2.71565
R274 VTAIL.n104 VTAIL.n56 2.71565
R275 VTAIL.n86 VTAIL.n66 2.71565
R276 VTAIL.n0 VTAIL.t7 2.10018
R277 VTAIL.n0 VTAIL.t6 2.10018
R278 VTAIL.n52 VTAIL.t2 2.10018
R279 VTAIL.n52 VTAIL.t0 2.10018
R280 VTAIL.n106 VTAIL.t3 2.10018
R281 VTAIL.n106 VTAIL.t1 2.10018
R282 VTAIL.n54 VTAIL.t5 2.10018
R283 VTAIL.n54 VTAIL.t9 2.10018
R284 VTAIL.n191 VTAIL.n189 1.93989
R285 VTAIL.n204 VTAIL.n203 1.93989
R286 VTAIL.n35 VTAIL.n33 1.93989
R287 VTAIL.n48 VTAIL.n47 1.93989
R288 VTAIL.n154 VTAIL.n153 1.93989
R289 VTAIL.n142 VTAIL.n141 1.93989
R290 VTAIL.n102 VTAIL.n101 1.93989
R291 VTAIL.n90 VTAIL.n89 1.93989
R292 VTAIL.n105 VTAIL.n55 1.50912
R293 VTAIL.n157 VTAIL.n107 1.50912
R294 VTAIL.n53 VTAIL.n51 1.50912
R295 VTAIL.n107 VTAIL.n105 1.22464
R296 VTAIL.n51 VTAIL.n1 1.22464
R297 VTAIL.n190 VTAIL.n164 1.16414
R298 VTAIL.n200 VTAIL.n160 1.16414
R299 VTAIL.n34 VTAIL.n8 1.16414
R300 VTAIL.n44 VTAIL.n4 1.16414
R301 VTAIL.n150 VTAIL.n110 1.16414
R302 VTAIL.n145 VTAIL.n115 1.16414
R303 VTAIL.n98 VTAIL.n58 1.16414
R304 VTAIL.n93 VTAIL.n63 1.16414
R305 VTAIL VTAIL.n207 1.07378
R306 VTAIL VTAIL.n1 0.435845
R307 VTAIL.n196 VTAIL.n195 0.388379
R308 VTAIL.n199 VTAIL.n162 0.388379
R309 VTAIL.n40 VTAIL.n39 0.388379
R310 VTAIL.n43 VTAIL.n6 0.388379
R311 VTAIL.n149 VTAIL.n112 0.388379
R312 VTAIL.n146 VTAIL.n114 0.388379
R313 VTAIL.n97 VTAIL.n60 0.388379
R314 VTAIL.n94 VTAIL.n62 0.388379
R315 VTAIL.n179 VTAIL.n171 0.155672
R316 VTAIL.n180 VTAIL.n179 0.155672
R317 VTAIL.n180 VTAIL.n167 0.155672
R318 VTAIL.n187 VTAIL.n167 0.155672
R319 VTAIL.n188 VTAIL.n187 0.155672
R320 VTAIL.n188 VTAIL.n163 0.155672
R321 VTAIL.n197 VTAIL.n163 0.155672
R322 VTAIL.n198 VTAIL.n197 0.155672
R323 VTAIL.n198 VTAIL.n159 0.155672
R324 VTAIL.n205 VTAIL.n159 0.155672
R325 VTAIL.n23 VTAIL.n15 0.155672
R326 VTAIL.n24 VTAIL.n23 0.155672
R327 VTAIL.n24 VTAIL.n11 0.155672
R328 VTAIL.n31 VTAIL.n11 0.155672
R329 VTAIL.n32 VTAIL.n31 0.155672
R330 VTAIL.n32 VTAIL.n7 0.155672
R331 VTAIL.n41 VTAIL.n7 0.155672
R332 VTAIL.n42 VTAIL.n41 0.155672
R333 VTAIL.n42 VTAIL.n3 0.155672
R334 VTAIL.n49 VTAIL.n3 0.155672
R335 VTAIL.n155 VTAIL.n109 0.155672
R336 VTAIL.n148 VTAIL.n109 0.155672
R337 VTAIL.n148 VTAIL.n147 0.155672
R338 VTAIL.n147 VTAIL.n113 0.155672
R339 VTAIL.n140 VTAIL.n113 0.155672
R340 VTAIL.n140 VTAIL.n139 0.155672
R341 VTAIL.n139 VTAIL.n119 0.155672
R342 VTAIL.n132 VTAIL.n119 0.155672
R343 VTAIL.n132 VTAIL.n131 0.155672
R344 VTAIL.n131 VTAIL.n123 0.155672
R345 VTAIL.n103 VTAIL.n57 0.155672
R346 VTAIL.n96 VTAIL.n57 0.155672
R347 VTAIL.n96 VTAIL.n95 0.155672
R348 VTAIL.n95 VTAIL.n61 0.155672
R349 VTAIL.n88 VTAIL.n61 0.155672
R350 VTAIL.n88 VTAIL.n87 0.155672
R351 VTAIL.n87 VTAIL.n67 0.155672
R352 VTAIL.n80 VTAIL.n67 0.155672
R353 VTAIL.n80 VTAIL.n79 0.155672
R354 VTAIL.n79 VTAIL.n71 0.155672
R355 VDD2.n95 VDD2.n51 289.615
R356 VDD2.n44 VDD2.n0 289.615
R357 VDD2.n96 VDD2.n95 185
R358 VDD2.n94 VDD2.n93 185
R359 VDD2.n55 VDD2.n54 185
R360 VDD2.n59 VDD2.n57 185
R361 VDD2.n88 VDD2.n87 185
R362 VDD2.n86 VDD2.n85 185
R363 VDD2.n61 VDD2.n60 185
R364 VDD2.n80 VDD2.n79 185
R365 VDD2.n78 VDD2.n77 185
R366 VDD2.n65 VDD2.n64 185
R367 VDD2.n72 VDD2.n71 185
R368 VDD2.n70 VDD2.n69 185
R369 VDD2.n17 VDD2.n16 185
R370 VDD2.n19 VDD2.n18 185
R371 VDD2.n12 VDD2.n11 185
R372 VDD2.n25 VDD2.n24 185
R373 VDD2.n27 VDD2.n26 185
R374 VDD2.n8 VDD2.n7 185
R375 VDD2.n34 VDD2.n33 185
R376 VDD2.n35 VDD2.n6 185
R377 VDD2.n37 VDD2.n36 185
R378 VDD2.n4 VDD2.n3 185
R379 VDD2.n43 VDD2.n42 185
R380 VDD2.n45 VDD2.n44 185
R381 VDD2.n68 VDD2.t2 149.524
R382 VDD2.n15 VDD2.t0 149.524
R383 VDD2.n95 VDD2.n94 104.615
R384 VDD2.n94 VDD2.n54 104.615
R385 VDD2.n59 VDD2.n54 104.615
R386 VDD2.n87 VDD2.n59 104.615
R387 VDD2.n87 VDD2.n86 104.615
R388 VDD2.n86 VDD2.n60 104.615
R389 VDD2.n79 VDD2.n60 104.615
R390 VDD2.n79 VDD2.n78 104.615
R391 VDD2.n78 VDD2.n64 104.615
R392 VDD2.n71 VDD2.n64 104.615
R393 VDD2.n71 VDD2.n70 104.615
R394 VDD2.n18 VDD2.n17 104.615
R395 VDD2.n18 VDD2.n11 104.615
R396 VDD2.n25 VDD2.n11 104.615
R397 VDD2.n26 VDD2.n25 104.615
R398 VDD2.n26 VDD2.n7 104.615
R399 VDD2.n34 VDD2.n7 104.615
R400 VDD2.n35 VDD2.n34 104.615
R401 VDD2.n36 VDD2.n35 104.615
R402 VDD2.n36 VDD2.n3 104.615
R403 VDD2.n43 VDD2.n3 104.615
R404 VDD2.n44 VDD2.n43 104.615
R405 VDD2.n50 VDD2.n49 67.0085
R406 VDD2 VDD2.n101 67.0057
R407 VDD2.n50 VDD2.n48 53.6251
R408 VDD2.n100 VDD2.n99 52.549
R409 VDD2.n70 VDD2.t2 52.3082
R410 VDD2.n17 VDD2.t0 52.3082
R411 VDD2.n100 VDD2.n50 36.7476
R412 VDD2.n57 VDD2.n55 13.1884
R413 VDD2.n37 VDD2.n4 13.1884
R414 VDD2.n93 VDD2.n92 12.8005
R415 VDD2.n89 VDD2.n88 12.8005
R416 VDD2.n38 VDD2.n6 12.8005
R417 VDD2.n42 VDD2.n41 12.8005
R418 VDD2.n96 VDD2.n53 12.0247
R419 VDD2.n85 VDD2.n58 12.0247
R420 VDD2.n33 VDD2.n32 12.0247
R421 VDD2.n45 VDD2.n2 12.0247
R422 VDD2.n97 VDD2.n51 11.249
R423 VDD2.n84 VDD2.n61 11.249
R424 VDD2.n31 VDD2.n8 11.249
R425 VDD2.n46 VDD2.n0 11.249
R426 VDD2.n81 VDD2.n80 10.4732
R427 VDD2.n28 VDD2.n27 10.4732
R428 VDD2.n69 VDD2.n68 10.2747
R429 VDD2.n16 VDD2.n15 10.2747
R430 VDD2.n77 VDD2.n63 9.69747
R431 VDD2.n24 VDD2.n10 9.69747
R432 VDD2.n99 VDD2.n98 9.45567
R433 VDD2.n48 VDD2.n47 9.45567
R434 VDD2.n67 VDD2.n66 9.3005
R435 VDD2.n74 VDD2.n73 9.3005
R436 VDD2.n76 VDD2.n75 9.3005
R437 VDD2.n63 VDD2.n62 9.3005
R438 VDD2.n82 VDD2.n81 9.3005
R439 VDD2.n84 VDD2.n83 9.3005
R440 VDD2.n58 VDD2.n56 9.3005
R441 VDD2.n90 VDD2.n89 9.3005
R442 VDD2.n98 VDD2.n97 9.3005
R443 VDD2.n53 VDD2.n52 9.3005
R444 VDD2.n92 VDD2.n91 9.3005
R445 VDD2.n47 VDD2.n46 9.3005
R446 VDD2.n2 VDD2.n1 9.3005
R447 VDD2.n41 VDD2.n40 9.3005
R448 VDD2.n14 VDD2.n13 9.3005
R449 VDD2.n21 VDD2.n20 9.3005
R450 VDD2.n23 VDD2.n22 9.3005
R451 VDD2.n10 VDD2.n9 9.3005
R452 VDD2.n29 VDD2.n28 9.3005
R453 VDD2.n31 VDD2.n30 9.3005
R454 VDD2.n32 VDD2.n5 9.3005
R455 VDD2.n39 VDD2.n38 9.3005
R456 VDD2.n76 VDD2.n65 8.92171
R457 VDD2.n23 VDD2.n12 8.92171
R458 VDD2.n73 VDD2.n72 8.14595
R459 VDD2.n20 VDD2.n19 8.14595
R460 VDD2.n69 VDD2.n67 7.3702
R461 VDD2.n16 VDD2.n14 7.3702
R462 VDD2.n72 VDD2.n67 5.81868
R463 VDD2.n19 VDD2.n14 5.81868
R464 VDD2.n73 VDD2.n65 5.04292
R465 VDD2.n20 VDD2.n12 5.04292
R466 VDD2.n77 VDD2.n76 4.26717
R467 VDD2.n24 VDD2.n23 4.26717
R468 VDD2.n80 VDD2.n63 3.49141
R469 VDD2.n27 VDD2.n10 3.49141
R470 VDD2.n68 VDD2.n66 2.84303
R471 VDD2.n15 VDD2.n13 2.84303
R472 VDD2.n99 VDD2.n51 2.71565
R473 VDD2.n81 VDD2.n61 2.71565
R474 VDD2.n28 VDD2.n8 2.71565
R475 VDD2.n48 VDD2.n0 2.71565
R476 VDD2.n101 VDD2.t3 2.10018
R477 VDD2.n101 VDD2.t1 2.10018
R478 VDD2.n49 VDD2.t4 2.10018
R479 VDD2.n49 VDD2.t5 2.10018
R480 VDD2.n97 VDD2.n96 1.93989
R481 VDD2.n85 VDD2.n84 1.93989
R482 VDD2.n33 VDD2.n31 1.93989
R483 VDD2.n46 VDD2.n45 1.93989
R484 VDD2 VDD2.n100 1.19016
R485 VDD2.n93 VDD2.n53 1.16414
R486 VDD2.n88 VDD2.n58 1.16414
R487 VDD2.n32 VDD2.n6 1.16414
R488 VDD2.n42 VDD2.n2 1.16414
R489 VDD2.n92 VDD2.n55 0.388379
R490 VDD2.n89 VDD2.n57 0.388379
R491 VDD2.n38 VDD2.n37 0.388379
R492 VDD2.n41 VDD2.n4 0.388379
R493 VDD2.n98 VDD2.n52 0.155672
R494 VDD2.n91 VDD2.n52 0.155672
R495 VDD2.n91 VDD2.n90 0.155672
R496 VDD2.n90 VDD2.n56 0.155672
R497 VDD2.n83 VDD2.n56 0.155672
R498 VDD2.n83 VDD2.n82 0.155672
R499 VDD2.n82 VDD2.n62 0.155672
R500 VDD2.n75 VDD2.n62 0.155672
R501 VDD2.n75 VDD2.n74 0.155672
R502 VDD2.n74 VDD2.n66 0.155672
R503 VDD2.n21 VDD2.n13 0.155672
R504 VDD2.n22 VDD2.n21 0.155672
R505 VDD2.n22 VDD2.n9 0.155672
R506 VDD2.n29 VDD2.n9 0.155672
R507 VDD2.n30 VDD2.n29 0.155672
R508 VDD2.n30 VDD2.n5 0.155672
R509 VDD2.n39 VDD2.n5 0.155672
R510 VDD2.n40 VDD2.n39 0.155672
R511 VDD2.n40 VDD2.n1 0.155672
R512 VDD2.n47 VDD2.n1 0.155672
R513 B.n629 B.n628 585
R514 B.n250 B.n93 585
R515 B.n249 B.n248 585
R516 B.n247 B.n246 585
R517 B.n245 B.n244 585
R518 B.n243 B.n242 585
R519 B.n241 B.n240 585
R520 B.n239 B.n238 585
R521 B.n237 B.n236 585
R522 B.n235 B.n234 585
R523 B.n233 B.n232 585
R524 B.n231 B.n230 585
R525 B.n229 B.n228 585
R526 B.n227 B.n226 585
R527 B.n225 B.n224 585
R528 B.n223 B.n222 585
R529 B.n221 B.n220 585
R530 B.n219 B.n218 585
R531 B.n217 B.n216 585
R532 B.n215 B.n214 585
R533 B.n213 B.n212 585
R534 B.n211 B.n210 585
R535 B.n209 B.n208 585
R536 B.n207 B.n206 585
R537 B.n205 B.n204 585
R538 B.n203 B.n202 585
R539 B.n201 B.n200 585
R540 B.n199 B.n198 585
R541 B.n197 B.n196 585
R542 B.n195 B.n194 585
R543 B.n193 B.n192 585
R544 B.n191 B.n190 585
R545 B.n189 B.n188 585
R546 B.n187 B.n186 585
R547 B.n185 B.n184 585
R548 B.n183 B.n182 585
R549 B.n181 B.n180 585
R550 B.n179 B.n178 585
R551 B.n177 B.n176 585
R552 B.n175 B.n174 585
R553 B.n173 B.n172 585
R554 B.n171 B.n170 585
R555 B.n169 B.n168 585
R556 B.n167 B.n166 585
R557 B.n165 B.n164 585
R558 B.n163 B.n162 585
R559 B.n161 B.n160 585
R560 B.n159 B.n158 585
R561 B.n157 B.n156 585
R562 B.n155 B.n154 585
R563 B.n153 B.n152 585
R564 B.n151 B.n150 585
R565 B.n149 B.n148 585
R566 B.n147 B.n146 585
R567 B.n145 B.n144 585
R568 B.n143 B.n142 585
R569 B.n141 B.n140 585
R570 B.n139 B.n138 585
R571 B.n137 B.n136 585
R572 B.n135 B.n134 585
R573 B.n133 B.n132 585
R574 B.n131 B.n130 585
R575 B.n129 B.n128 585
R576 B.n127 B.n126 585
R577 B.n125 B.n124 585
R578 B.n123 B.n122 585
R579 B.n121 B.n120 585
R580 B.n119 B.n118 585
R581 B.n117 B.n116 585
R582 B.n115 B.n114 585
R583 B.n113 B.n112 585
R584 B.n111 B.n110 585
R585 B.n109 B.n108 585
R586 B.n107 B.n106 585
R587 B.n105 B.n104 585
R588 B.n103 B.n102 585
R589 B.n101 B.n100 585
R590 B.n53 B.n52 585
R591 B.n627 B.n54 585
R592 B.n632 B.n54 585
R593 B.n626 B.n625 585
R594 B.n625 B.n50 585
R595 B.n624 B.n49 585
R596 B.n638 B.n49 585
R597 B.n623 B.n48 585
R598 B.n639 B.n48 585
R599 B.n622 B.n47 585
R600 B.n640 B.n47 585
R601 B.n621 B.n620 585
R602 B.n620 B.n46 585
R603 B.n619 B.n42 585
R604 B.n646 B.n42 585
R605 B.n618 B.n41 585
R606 B.n647 B.n41 585
R607 B.n617 B.n40 585
R608 B.n648 B.n40 585
R609 B.n616 B.n615 585
R610 B.n615 B.n36 585
R611 B.n614 B.n35 585
R612 B.n654 B.n35 585
R613 B.n613 B.n34 585
R614 B.n655 B.n34 585
R615 B.n612 B.n33 585
R616 B.n656 B.n33 585
R617 B.n611 B.n610 585
R618 B.n610 B.n29 585
R619 B.n609 B.n28 585
R620 B.n662 B.n28 585
R621 B.n608 B.n27 585
R622 B.n663 B.n27 585
R623 B.n607 B.n26 585
R624 B.n664 B.n26 585
R625 B.n606 B.n605 585
R626 B.n605 B.n22 585
R627 B.n604 B.n21 585
R628 B.n670 B.n21 585
R629 B.n603 B.n20 585
R630 B.n671 B.n20 585
R631 B.n602 B.n19 585
R632 B.n672 B.n19 585
R633 B.n601 B.n600 585
R634 B.n600 B.n15 585
R635 B.n599 B.n14 585
R636 B.n678 B.n14 585
R637 B.n598 B.n13 585
R638 B.n679 B.n13 585
R639 B.n597 B.n12 585
R640 B.n680 B.n12 585
R641 B.n596 B.n595 585
R642 B.n595 B.n594 585
R643 B.n593 B.n592 585
R644 B.n593 B.n8 585
R645 B.n591 B.n7 585
R646 B.n687 B.n7 585
R647 B.n590 B.n6 585
R648 B.n688 B.n6 585
R649 B.n589 B.n5 585
R650 B.n689 B.n5 585
R651 B.n588 B.n587 585
R652 B.n587 B.n4 585
R653 B.n586 B.n251 585
R654 B.n586 B.n585 585
R655 B.n576 B.n252 585
R656 B.n253 B.n252 585
R657 B.n578 B.n577 585
R658 B.n579 B.n578 585
R659 B.n575 B.n258 585
R660 B.n258 B.n257 585
R661 B.n574 B.n573 585
R662 B.n573 B.n572 585
R663 B.n260 B.n259 585
R664 B.n261 B.n260 585
R665 B.n565 B.n564 585
R666 B.n566 B.n565 585
R667 B.n563 B.n265 585
R668 B.n269 B.n265 585
R669 B.n562 B.n561 585
R670 B.n561 B.n560 585
R671 B.n267 B.n266 585
R672 B.n268 B.n267 585
R673 B.n553 B.n552 585
R674 B.n554 B.n553 585
R675 B.n551 B.n274 585
R676 B.n274 B.n273 585
R677 B.n550 B.n549 585
R678 B.n549 B.n548 585
R679 B.n276 B.n275 585
R680 B.n277 B.n276 585
R681 B.n541 B.n540 585
R682 B.n542 B.n541 585
R683 B.n539 B.n282 585
R684 B.n282 B.n281 585
R685 B.n538 B.n537 585
R686 B.n537 B.n536 585
R687 B.n284 B.n283 585
R688 B.n285 B.n284 585
R689 B.n529 B.n528 585
R690 B.n530 B.n529 585
R691 B.n527 B.n290 585
R692 B.n290 B.n289 585
R693 B.n526 B.n525 585
R694 B.n525 B.n524 585
R695 B.n292 B.n291 585
R696 B.n517 B.n292 585
R697 B.n516 B.n515 585
R698 B.n518 B.n516 585
R699 B.n514 B.n297 585
R700 B.n297 B.n296 585
R701 B.n513 B.n512 585
R702 B.n512 B.n511 585
R703 B.n299 B.n298 585
R704 B.n300 B.n299 585
R705 B.n504 B.n503 585
R706 B.n505 B.n504 585
R707 B.n303 B.n302 585
R708 B.n348 B.n346 585
R709 B.n349 B.n345 585
R710 B.n349 B.n304 585
R711 B.n352 B.n351 585
R712 B.n353 B.n344 585
R713 B.n355 B.n354 585
R714 B.n357 B.n343 585
R715 B.n360 B.n359 585
R716 B.n361 B.n342 585
R717 B.n363 B.n362 585
R718 B.n365 B.n341 585
R719 B.n368 B.n367 585
R720 B.n369 B.n340 585
R721 B.n371 B.n370 585
R722 B.n373 B.n339 585
R723 B.n376 B.n375 585
R724 B.n377 B.n338 585
R725 B.n379 B.n378 585
R726 B.n381 B.n337 585
R727 B.n384 B.n383 585
R728 B.n385 B.n336 585
R729 B.n387 B.n386 585
R730 B.n389 B.n335 585
R731 B.n392 B.n391 585
R732 B.n393 B.n334 585
R733 B.n395 B.n394 585
R734 B.n397 B.n333 585
R735 B.n400 B.n399 585
R736 B.n401 B.n332 585
R737 B.n403 B.n402 585
R738 B.n405 B.n331 585
R739 B.n408 B.n407 585
R740 B.n409 B.n330 585
R741 B.n414 B.n413 585
R742 B.n416 B.n329 585
R743 B.n419 B.n418 585
R744 B.n420 B.n328 585
R745 B.n422 B.n421 585
R746 B.n424 B.n327 585
R747 B.n427 B.n426 585
R748 B.n428 B.n326 585
R749 B.n430 B.n429 585
R750 B.n432 B.n325 585
R751 B.n435 B.n434 585
R752 B.n437 B.n322 585
R753 B.n439 B.n438 585
R754 B.n441 B.n321 585
R755 B.n444 B.n443 585
R756 B.n445 B.n320 585
R757 B.n447 B.n446 585
R758 B.n449 B.n319 585
R759 B.n452 B.n451 585
R760 B.n453 B.n318 585
R761 B.n455 B.n454 585
R762 B.n457 B.n317 585
R763 B.n460 B.n459 585
R764 B.n461 B.n316 585
R765 B.n463 B.n462 585
R766 B.n465 B.n315 585
R767 B.n468 B.n467 585
R768 B.n469 B.n314 585
R769 B.n471 B.n470 585
R770 B.n473 B.n313 585
R771 B.n476 B.n475 585
R772 B.n477 B.n312 585
R773 B.n479 B.n478 585
R774 B.n481 B.n311 585
R775 B.n484 B.n483 585
R776 B.n485 B.n310 585
R777 B.n487 B.n486 585
R778 B.n489 B.n309 585
R779 B.n492 B.n491 585
R780 B.n493 B.n308 585
R781 B.n495 B.n494 585
R782 B.n497 B.n307 585
R783 B.n498 B.n306 585
R784 B.n501 B.n500 585
R785 B.n502 B.n305 585
R786 B.n305 B.n304 585
R787 B.n507 B.n506 585
R788 B.n506 B.n505 585
R789 B.n508 B.n301 585
R790 B.n301 B.n300 585
R791 B.n510 B.n509 585
R792 B.n511 B.n510 585
R793 B.n295 B.n294 585
R794 B.n296 B.n295 585
R795 B.n520 B.n519 585
R796 B.n519 B.n518 585
R797 B.n521 B.n293 585
R798 B.n517 B.n293 585
R799 B.n523 B.n522 585
R800 B.n524 B.n523 585
R801 B.n288 B.n287 585
R802 B.n289 B.n288 585
R803 B.n532 B.n531 585
R804 B.n531 B.n530 585
R805 B.n533 B.n286 585
R806 B.n286 B.n285 585
R807 B.n535 B.n534 585
R808 B.n536 B.n535 585
R809 B.n280 B.n279 585
R810 B.n281 B.n280 585
R811 B.n544 B.n543 585
R812 B.n543 B.n542 585
R813 B.n545 B.n278 585
R814 B.n278 B.n277 585
R815 B.n547 B.n546 585
R816 B.n548 B.n547 585
R817 B.n272 B.n271 585
R818 B.n273 B.n272 585
R819 B.n556 B.n555 585
R820 B.n555 B.n554 585
R821 B.n557 B.n270 585
R822 B.n270 B.n268 585
R823 B.n559 B.n558 585
R824 B.n560 B.n559 585
R825 B.n264 B.n263 585
R826 B.n269 B.n264 585
R827 B.n568 B.n567 585
R828 B.n567 B.n566 585
R829 B.n569 B.n262 585
R830 B.n262 B.n261 585
R831 B.n571 B.n570 585
R832 B.n572 B.n571 585
R833 B.n256 B.n255 585
R834 B.n257 B.n256 585
R835 B.n581 B.n580 585
R836 B.n580 B.n579 585
R837 B.n582 B.n254 585
R838 B.n254 B.n253 585
R839 B.n584 B.n583 585
R840 B.n585 B.n584 585
R841 B.n3 B.n0 585
R842 B.n4 B.n3 585
R843 B.n686 B.n1 585
R844 B.n687 B.n686 585
R845 B.n685 B.n684 585
R846 B.n685 B.n8 585
R847 B.n683 B.n9 585
R848 B.n594 B.n9 585
R849 B.n682 B.n681 585
R850 B.n681 B.n680 585
R851 B.n11 B.n10 585
R852 B.n679 B.n11 585
R853 B.n677 B.n676 585
R854 B.n678 B.n677 585
R855 B.n675 B.n16 585
R856 B.n16 B.n15 585
R857 B.n674 B.n673 585
R858 B.n673 B.n672 585
R859 B.n18 B.n17 585
R860 B.n671 B.n18 585
R861 B.n669 B.n668 585
R862 B.n670 B.n669 585
R863 B.n667 B.n23 585
R864 B.n23 B.n22 585
R865 B.n666 B.n665 585
R866 B.n665 B.n664 585
R867 B.n25 B.n24 585
R868 B.n663 B.n25 585
R869 B.n661 B.n660 585
R870 B.n662 B.n661 585
R871 B.n659 B.n30 585
R872 B.n30 B.n29 585
R873 B.n658 B.n657 585
R874 B.n657 B.n656 585
R875 B.n32 B.n31 585
R876 B.n655 B.n32 585
R877 B.n653 B.n652 585
R878 B.n654 B.n653 585
R879 B.n651 B.n37 585
R880 B.n37 B.n36 585
R881 B.n650 B.n649 585
R882 B.n649 B.n648 585
R883 B.n39 B.n38 585
R884 B.n647 B.n39 585
R885 B.n645 B.n644 585
R886 B.n646 B.n645 585
R887 B.n643 B.n43 585
R888 B.n46 B.n43 585
R889 B.n642 B.n641 585
R890 B.n641 B.n640 585
R891 B.n45 B.n44 585
R892 B.n639 B.n45 585
R893 B.n637 B.n636 585
R894 B.n638 B.n637 585
R895 B.n635 B.n51 585
R896 B.n51 B.n50 585
R897 B.n634 B.n633 585
R898 B.n633 B.n632 585
R899 B.n690 B.n689 585
R900 B.n688 B.n2 585
R901 B.n633 B.n53 506.916
R902 B.n629 B.n54 506.916
R903 B.n504 B.n305 506.916
R904 B.n506 B.n303 506.916
R905 B.n97 B.t17 365.173
R906 B.n94 B.t6 365.173
R907 B.n323 B.t10 365.173
R908 B.n410 B.t14 365.173
R909 B.n94 B.t8 272.009
R910 B.n323 B.t13 272.009
R911 B.n97 B.t18 272.009
R912 B.n410 B.t16 272.009
R913 B.n631 B.n630 256.663
R914 B.n631 B.n92 256.663
R915 B.n631 B.n91 256.663
R916 B.n631 B.n90 256.663
R917 B.n631 B.n89 256.663
R918 B.n631 B.n88 256.663
R919 B.n631 B.n87 256.663
R920 B.n631 B.n86 256.663
R921 B.n631 B.n85 256.663
R922 B.n631 B.n84 256.663
R923 B.n631 B.n83 256.663
R924 B.n631 B.n82 256.663
R925 B.n631 B.n81 256.663
R926 B.n631 B.n80 256.663
R927 B.n631 B.n79 256.663
R928 B.n631 B.n78 256.663
R929 B.n631 B.n77 256.663
R930 B.n631 B.n76 256.663
R931 B.n631 B.n75 256.663
R932 B.n631 B.n74 256.663
R933 B.n631 B.n73 256.663
R934 B.n631 B.n72 256.663
R935 B.n631 B.n71 256.663
R936 B.n631 B.n70 256.663
R937 B.n631 B.n69 256.663
R938 B.n631 B.n68 256.663
R939 B.n631 B.n67 256.663
R940 B.n631 B.n66 256.663
R941 B.n631 B.n65 256.663
R942 B.n631 B.n64 256.663
R943 B.n631 B.n63 256.663
R944 B.n631 B.n62 256.663
R945 B.n631 B.n61 256.663
R946 B.n631 B.n60 256.663
R947 B.n631 B.n59 256.663
R948 B.n631 B.n58 256.663
R949 B.n631 B.n57 256.663
R950 B.n631 B.n56 256.663
R951 B.n631 B.n55 256.663
R952 B.n347 B.n304 256.663
R953 B.n350 B.n304 256.663
R954 B.n356 B.n304 256.663
R955 B.n358 B.n304 256.663
R956 B.n364 B.n304 256.663
R957 B.n366 B.n304 256.663
R958 B.n372 B.n304 256.663
R959 B.n374 B.n304 256.663
R960 B.n380 B.n304 256.663
R961 B.n382 B.n304 256.663
R962 B.n388 B.n304 256.663
R963 B.n390 B.n304 256.663
R964 B.n396 B.n304 256.663
R965 B.n398 B.n304 256.663
R966 B.n404 B.n304 256.663
R967 B.n406 B.n304 256.663
R968 B.n415 B.n304 256.663
R969 B.n417 B.n304 256.663
R970 B.n423 B.n304 256.663
R971 B.n425 B.n304 256.663
R972 B.n431 B.n304 256.663
R973 B.n433 B.n304 256.663
R974 B.n440 B.n304 256.663
R975 B.n442 B.n304 256.663
R976 B.n448 B.n304 256.663
R977 B.n450 B.n304 256.663
R978 B.n456 B.n304 256.663
R979 B.n458 B.n304 256.663
R980 B.n464 B.n304 256.663
R981 B.n466 B.n304 256.663
R982 B.n472 B.n304 256.663
R983 B.n474 B.n304 256.663
R984 B.n480 B.n304 256.663
R985 B.n482 B.n304 256.663
R986 B.n488 B.n304 256.663
R987 B.n490 B.n304 256.663
R988 B.n496 B.n304 256.663
R989 B.n499 B.n304 256.663
R990 B.n692 B.n691 256.663
R991 B.n95 B.t9 238.069
R992 B.n324 B.t12 238.069
R993 B.n98 B.t19 238.069
R994 B.n411 B.t15 238.069
R995 B.n102 B.n101 163.367
R996 B.n106 B.n105 163.367
R997 B.n110 B.n109 163.367
R998 B.n114 B.n113 163.367
R999 B.n118 B.n117 163.367
R1000 B.n122 B.n121 163.367
R1001 B.n126 B.n125 163.367
R1002 B.n130 B.n129 163.367
R1003 B.n134 B.n133 163.367
R1004 B.n138 B.n137 163.367
R1005 B.n142 B.n141 163.367
R1006 B.n146 B.n145 163.367
R1007 B.n150 B.n149 163.367
R1008 B.n154 B.n153 163.367
R1009 B.n158 B.n157 163.367
R1010 B.n162 B.n161 163.367
R1011 B.n166 B.n165 163.367
R1012 B.n170 B.n169 163.367
R1013 B.n174 B.n173 163.367
R1014 B.n178 B.n177 163.367
R1015 B.n182 B.n181 163.367
R1016 B.n186 B.n185 163.367
R1017 B.n190 B.n189 163.367
R1018 B.n194 B.n193 163.367
R1019 B.n198 B.n197 163.367
R1020 B.n202 B.n201 163.367
R1021 B.n206 B.n205 163.367
R1022 B.n210 B.n209 163.367
R1023 B.n214 B.n213 163.367
R1024 B.n218 B.n217 163.367
R1025 B.n222 B.n221 163.367
R1026 B.n226 B.n225 163.367
R1027 B.n230 B.n229 163.367
R1028 B.n234 B.n233 163.367
R1029 B.n238 B.n237 163.367
R1030 B.n242 B.n241 163.367
R1031 B.n246 B.n245 163.367
R1032 B.n248 B.n93 163.367
R1033 B.n504 B.n299 163.367
R1034 B.n512 B.n299 163.367
R1035 B.n512 B.n297 163.367
R1036 B.n516 B.n297 163.367
R1037 B.n516 B.n292 163.367
R1038 B.n525 B.n292 163.367
R1039 B.n525 B.n290 163.367
R1040 B.n529 B.n290 163.367
R1041 B.n529 B.n284 163.367
R1042 B.n537 B.n284 163.367
R1043 B.n537 B.n282 163.367
R1044 B.n541 B.n282 163.367
R1045 B.n541 B.n276 163.367
R1046 B.n549 B.n276 163.367
R1047 B.n549 B.n274 163.367
R1048 B.n553 B.n274 163.367
R1049 B.n553 B.n267 163.367
R1050 B.n561 B.n267 163.367
R1051 B.n561 B.n265 163.367
R1052 B.n565 B.n265 163.367
R1053 B.n565 B.n260 163.367
R1054 B.n573 B.n260 163.367
R1055 B.n573 B.n258 163.367
R1056 B.n578 B.n258 163.367
R1057 B.n578 B.n252 163.367
R1058 B.n586 B.n252 163.367
R1059 B.n587 B.n586 163.367
R1060 B.n587 B.n5 163.367
R1061 B.n6 B.n5 163.367
R1062 B.n7 B.n6 163.367
R1063 B.n593 B.n7 163.367
R1064 B.n595 B.n593 163.367
R1065 B.n595 B.n12 163.367
R1066 B.n13 B.n12 163.367
R1067 B.n14 B.n13 163.367
R1068 B.n600 B.n14 163.367
R1069 B.n600 B.n19 163.367
R1070 B.n20 B.n19 163.367
R1071 B.n21 B.n20 163.367
R1072 B.n605 B.n21 163.367
R1073 B.n605 B.n26 163.367
R1074 B.n27 B.n26 163.367
R1075 B.n28 B.n27 163.367
R1076 B.n610 B.n28 163.367
R1077 B.n610 B.n33 163.367
R1078 B.n34 B.n33 163.367
R1079 B.n35 B.n34 163.367
R1080 B.n615 B.n35 163.367
R1081 B.n615 B.n40 163.367
R1082 B.n41 B.n40 163.367
R1083 B.n42 B.n41 163.367
R1084 B.n620 B.n42 163.367
R1085 B.n620 B.n47 163.367
R1086 B.n48 B.n47 163.367
R1087 B.n49 B.n48 163.367
R1088 B.n625 B.n49 163.367
R1089 B.n625 B.n54 163.367
R1090 B.n349 B.n348 163.367
R1091 B.n351 B.n349 163.367
R1092 B.n355 B.n344 163.367
R1093 B.n359 B.n357 163.367
R1094 B.n363 B.n342 163.367
R1095 B.n367 B.n365 163.367
R1096 B.n371 B.n340 163.367
R1097 B.n375 B.n373 163.367
R1098 B.n379 B.n338 163.367
R1099 B.n383 B.n381 163.367
R1100 B.n387 B.n336 163.367
R1101 B.n391 B.n389 163.367
R1102 B.n395 B.n334 163.367
R1103 B.n399 B.n397 163.367
R1104 B.n403 B.n332 163.367
R1105 B.n407 B.n405 163.367
R1106 B.n414 B.n330 163.367
R1107 B.n418 B.n416 163.367
R1108 B.n422 B.n328 163.367
R1109 B.n426 B.n424 163.367
R1110 B.n430 B.n326 163.367
R1111 B.n434 B.n432 163.367
R1112 B.n439 B.n322 163.367
R1113 B.n443 B.n441 163.367
R1114 B.n447 B.n320 163.367
R1115 B.n451 B.n449 163.367
R1116 B.n455 B.n318 163.367
R1117 B.n459 B.n457 163.367
R1118 B.n463 B.n316 163.367
R1119 B.n467 B.n465 163.367
R1120 B.n471 B.n314 163.367
R1121 B.n475 B.n473 163.367
R1122 B.n479 B.n312 163.367
R1123 B.n483 B.n481 163.367
R1124 B.n487 B.n310 163.367
R1125 B.n491 B.n489 163.367
R1126 B.n495 B.n308 163.367
R1127 B.n498 B.n497 163.367
R1128 B.n500 B.n305 163.367
R1129 B.n506 B.n301 163.367
R1130 B.n510 B.n301 163.367
R1131 B.n510 B.n295 163.367
R1132 B.n519 B.n295 163.367
R1133 B.n519 B.n293 163.367
R1134 B.n523 B.n293 163.367
R1135 B.n523 B.n288 163.367
R1136 B.n531 B.n288 163.367
R1137 B.n531 B.n286 163.367
R1138 B.n535 B.n286 163.367
R1139 B.n535 B.n280 163.367
R1140 B.n543 B.n280 163.367
R1141 B.n543 B.n278 163.367
R1142 B.n547 B.n278 163.367
R1143 B.n547 B.n272 163.367
R1144 B.n555 B.n272 163.367
R1145 B.n555 B.n270 163.367
R1146 B.n559 B.n270 163.367
R1147 B.n559 B.n264 163.367
R1148 B.n567 B.n264 163.367
R1149 B.n567 B.n262 163.367
R1150 B.n571 B.n262 163.367
R1151 B.n571 B.n256 163.367
R1152 B.n580 B.n256 163.367
R1153 B.n580 B.n254 163.367
R1154 B.n584 B.n254 163.367
R1155 B.n584 B.n3 163.367
R1156 B.n690 B.n3 163.367
R1157 B.n686 B.n2 163.367
R1158 B.n686 B.n685 163.367
R1159 B.n685 B.n9 163.367
R1160 B.n681 B.n9 163.367
R1161 B.n681 B.n11 163.367
R1162 B.n677 B.n11 163.367
R1163 B.n677 B.n16 163.367
R1164 B.n673 B.n16 163.367
R1165 B.n673 B.n18 163.367
R1166 B.n669 B.n18 163.367
R1167 B.n669 B.n23 163.367
R1168 B.n665 B.n23 163.367
R1169 B.n665 B.n25 163.367
R1170 B.n661 B.n25 163.367
R1171 B.n661 B.n30 163.367
R1172 B.n657 B.n30 163.367
R1173 B.n657 B.n32 163.367
R1174 B.n653 B.n32 163.367
R1175 B.n653 B.n37 163.367
R1176 B.n649 B.n37 163.367
R1177 B.n649 B.n39 163.367
R1178 B.n645 B.n39 163.367
R1179 B.n645 B.n43 163.367
R1180 B.n641 B.n43 163.367
R1181 B.n641 B.n45 163.367
R1182 B.n637 B.n45 163.367
R1183 B.n637 B.n51 163.367
R1184 B.n633 B.n51 163.367
R1185 B.n505 B.n304 102.483
R1186 B.n632 B.n631 102.483
R1187 B.n55 B.n53 71.676
R1188 B.n102 B.n56 71.676
R1189 B.n106 B.n57 71.676
R1190 B.n110 B.n58 71.676
R1191 B.n114 B.n59 71.676
R1192 B.n118 B.n60 71.676
R1193 B.n122 B.n61 71.676
R1194 B.n126 B.n62 71.676
R1195 B.n130 B.n63 71.676
R1196 B.n134 B.n64 71.676
R1197 B.n138 B.n65 71.676
R1198 B.n142 B.n66 71.676
R1199 B.n146 B.n67 71.676
R1200 B.n150 B.n68 71.676
R1201 B.n154 B.n69 71.676
R1202 B.n158 B.n70 71.676
R1203 B.n162 B.n71 71.676
R1204 B.n166 B.n72 71.676
R1205 B.n170 B.n73 71.676
R1206 B.n174 B.n74 71.676
R1207 B.n178 B.n75 71.676
R1208 B.n182 B.n76 71.676
R1209 B.n186 B.n77 71.676
R1210 B.n190 B.n78 71.676
R1211 B.n194 B.n79 71.676
R1212 B.n198 B.n80 71.676
R1213 B.n202 B.n81 71.676
R1214 B.n206 B.n82 71.676
R1215 B.n210 B.n83 71.676
R1216 B.n214 B.n84 71.676
R1217 B.n218 B.n85 71.676
R1218 B.n222 B.n86 71.676
R1219 B.n226 B.n87 71.676
R1220 B.n230 B.n88 71.676
R1221 B.n234 B.n89 71.676
R1222 B.n238 B.n90 71.676
R1223 B.n242 B.n91 71.676
R1224 B.n246 B.n92 71.676
R1225 B.n630 B.n93 71.676
R1226 B.n630 B.n629 71.676
R1227 B.n248 B.n92 71.676
R1228 B.n245 B.n91 71.676
R1229 B.n241 B.n90 71.676
R1230 B.n237 B.n89 71.676
R1231 B.n233 B.n88 71.676
R1232 B.n229 B.n87 71.676
R1233 B.n225 B.n86 71.676
R1234 B.n221 B.n85 71.676
R1235 B.n217 B.n84 71.676
R1236 B.n213 B.n83 71.676
R1237 B.n209 B.n82 71.676
R1238 B.n205 B.n81 71.676
R1239 B.n201 B.n80 71.676
R1240 B.n197 B.n79 71.676
R1241 B.n193 B.n78 71.676
R1242 B.n189 B.n77 71.676
R1243 B.n185 B.n76 71.676
R1244 B.n181 B.n75 71.676
R1245 B.n177 B.n74 71.676
R1246 B.n173 B.n73 71.676
R1247 B.n169 B.n72 71.676
R1248 B.n165 B.n71 71.676
R1249 B.n161 B.n70 71.676
R1250 B.n157 B.n69 71.676
R1251 B.n153 B.n68 71.676
R1252 B.n149 B.n67 71.676
R1253 B.n145 B.n66 71.676
R1254 B.n141 B.n65 71.676
R1255 B.n137 B.n64 71.676
R1256 B.n133 B.n63 71.676
R1257 B.n129 B.n62 71.676
R1258 B.n125 B.n61 71.676
R1259 B.n121 B.n60 71.676
R1260 B.n117 B.n59 71.676
R1261 B.n113 B.n58 71.676
R1262 B.n109 B.n57 71.676
R1263 B.n105 B.n56 71.676
R1264 B.n101 B.n55 71.676
R1265 B.n347 B.n303 71.676
R1266 B.n351 B.n350 71.676
R1267 B.n356 B.n355 71.676
R1268 B.n359 B.n358 71.676
R1269 B.n364 B.n363 71.676
R1270 B.n367 B.n366 71.676
R1271 B.n372 B.n371 71.676
R1272 B.n375 B.n374 71.676
R1273 B.n380 B.n379 71.676
R1274 B.n383 B.n382 71.676
R1275 B.n388 B.n387 71.676
R1276 B.n391 B.n390 71.676
R1277 B.n396 B.n395 71.676
R1278 B.n399 B.n398 71.676
R1279 B.n404 B.n403 71.676
R1280 B.n407 B.n406 71.676
R1281 B.n415 B.n414 71.676
R1282 B.n418 B.n417 71.676
R1283 B.n423 B.n422 71.676
R1284 B.n426 B.n425 71.676
R1285 B.n431 B.n430 71.676
R1286 B.n434 B.n433 71.676
R1287 B.n440 B.n439 71.676
R1288 B.n443 B.n442 71.676
R1289 B.n448 B.n447 71.676
R1290 B.n451 B.n450 71.676
R1291 B.n456 B.n455 71.676
R1292 B.n459 B.n458 71.676
R1293 B.n464 B.n463 71.676
R1294 B.n467 B.n466 71.676
R1295 B.n472 B.n471 71.676
R1296 B.n475 B.n474 71.676
R1297 B.n480 B.n479 71.676
R1298 B.n483 B.n482 71.676
R1299 B.n488 B.n487 71.676
R1300 B.n491 B.n490 71.676
R1301 B.n496 B.n495 71.676
R1302 B.n499 B.n498 71.676
R1303 B.n348 B.n347 71.676
R1304 B.n350 B.n344 71.676
R1305 B.n357 B.n356 71.676
R1306 B.n358 B.n342 71.676
R1307 B.n365 B.n364 71.676
R1308 B.n366 B.n340 71.676
R1309 B.n373 B.n372 71.676
R1310 B.n374 B.n338 71.676
R1311 B.n381 B.n380 71.676
R1312 B.n382 B.n336 71.676
R1313 B.n389 B.n388 71.676
R1314 B.n390 B.n334 71.676
R1315 B.n397 B.n396 71.676
R1316 B.n398 B.n332 71.676
R1317 B.n405 B.n404 71.676
R1318 B.n406 B.n330 71.676
R1319 B.n416 B.n415 71.676
R1320 B.n417 B.n328 71.676
R1321 B.n424 B.n423 71.676
R1322 B.n425 B.n326 71.676
R1323 B.n432 B.n431 71.676
R1324 B.n433 B.n322 71.676
R1325 B.n441 B.n440 71.676
R1326 B.n442 B.n320 71.676
R1327 B.n449 B.n448 71.676
R1328 B.n450 B.n318 71.676
R1329 B.n457 B.n456 71.676
R1330 B.n458 B.n316 71.676
R1331 B.n465 B.n464 71.676
R1332 B.n466 B.n314 71.676
R1333 B.n473 B.n472 71.676
R1334 B.n474 B.n312 71.676
R1335 B.n481 B.n480 71.676
R1336 B.n482 B.n310 71.676
R1337 B.n489 B.n488 71.676
R1338 B.n490 B.n308 71.676
R1339 B.n497 B.n496 71.676
R1340 B.n500 B.n499 71.676
R1341 B.n691 B.n690 71.676
R1342 B.n691 B.n2 71.676
R1343 B.n99 B.n98 59.5399
R1344 B.n96 B.n95 59.5399
R1345 B.n436 B.n324 59.5399
R1346 B.n412 B.n411 59.5399
R1347 B.n505 B.n300 50.8676
R1348 B.n511 B.n300 50.8676
R1349 B.n511 B.n296 50.8676
R1350 B.n518 B.n296 50.8676
R1351 B.n518 B.n517 50.8676
R1352 B.n524 B.n289 50.8676
R1353 B.n530 B.n289 50.8676
R1354 B.n530 B.n285 50.8676
R1355 B.n536 B.n285 50.8676
R1356 B.n536 B.n281 50.8676
R1357 B.n542 B.n281 50.8676
R1358 B.n542 B.n277 50.8676
R1359 B.n548 B.n277 50.8676
R1360 B.n554 B.n273 50.8676
R1361 B.n554 B.n268 50.8676
R1362 B.n560 B.n268 50.8676
R1363 B.n560 B.n269 50.8676
R1364 B.n566 B.n261 50.8676
R1365 B.n572 B.n261 50.8676
R1366 B.n572 B.n257 50.8676
R1367 B.n579 B.n257 50.8676
R1368 B.n585 B.n253 50.8676
R1369 B.n585 B.n4 50.8676
R1370 B.n689 B.n4 50.8676
R1371 B.n689 B.n688 50.8676
R1372 B.n688 B.n687 50.8676
R1373 B.n687 B.n8 50.8676
R1374 B.n594 B.n8 50.8676
R1375 B.n680 B.n679 50.8676
R1376 B.n679 B.n678 50.8676
R1377 B.n678 B.n15 50.8676
R1378 B.n672 B.n15 50.8676
R1379 B.n671 B.n670 50.8676
R1380 B.n670 B.n22 50.8676
R1381 B.n664 B.n22 50.8676
R1382 B.n664 B.n663 50.8676
R1383 B.n662 B.n29 50.8676
R1384 B.n656 B.n29 50.8676
R1385 B.n656 B.n655 50.8676
R1386 B.n655 B.n654 50.8676
R1387 B.n654 B.n36 50.8676
R1388 B.n648 B.n36 50.8676
R1389 B.n648 B.n647 50.8676
R1390 B.n647 B.n646 50.8676
R1391 B.n640 B.n46 50.8676
R1392 B.n640 B.n639 50.8676
R1393 B.n639 B.n638 50.8676
R1394 B.n638 B.n50 50.8676
R1395 B.n632 B.n50 50.8676
R1396 B.t2 B.n273 49.3715
R1397 B.n663 B.t5 49.3715
R1398 B.n566 B.t0 41.891
R1399 B.n672 B.t1 41.891
R1400 B.n517 B.t11 34.4106
R1401 B.t4 B.n253 34.4106
R1402 B.n594 B.t3 34.4106
R1403 B.n46 B.t7 34.4106
R1404 B.n98 B.n97 33.9399
R1405 B.n95 B.n94 33.9399
R1406 B.n324 B.n323 33.9399
R1407 B.n411 B.n410 33.9399
R1408 B.n507 B.n302 32.9371
R1409 B.n503 B.n502 32.9371
R1410 B.n628 B.n627 32.9371
R1411 B.n634 B.n52 32.9371
R1412 B B.n692 18.0485
R1413 B.n524 B.t11 16.4575
R1414 B.n579 B.t4 16.4575
R1415 B.n680 B.t3 16.4575
R1416 B.n646 B.t7 16.4575
R1417 B.n508 B.n507 10.6151
R1418 B.n509 B.n508 10.6151
R1419 B.n509 B.n294 10.6151
R1420 B.n520 B.n294 10.6151
R1421 B.n521 B.n520 10.6151
R1422 B.n522 B.n521 10.6151
R1423 B.n522 B.n287 10.6151
R1424 B.n532 B.n287 10.6151
R1425 B.n533 B.n532 10.6151
R1426 B.n534 B.n533 10.6151
R1427 B.n534 B.n279 10.6151
R1428 B.n544 B.n279 10.6151
R1429 B.n545 B.n544 10.6151
R1430 B.n546 B.n545 10.6151
R1431 B.n546 B.n271 10.6151
R1432 B.n556 B.n271 10.6151
R1433 B.n557 B.n556 10.6151
R1434 B.n558 B.n557 10.6151
R1435 B.n558 B.n263 10.6151
R1436 B.n568 B.n263 10.6151
R1437 B.n569 B.n568 10.6151
R1438 B.n570 B.n569 10.6151
R1439 B.n570 B.n255 10.6151
R1440 B.n581 B.n255 10.6151
R1441 B.n582 B.n581 10.6151
R1442 B.n583 B.n582 10.6151
R1443 B.n583 B.n0 10.6151
R1444 B.n346 B.n302 10.6151
R1445 B.n346 B.n345 10.6151
R1446 B.n352 B.n345 10.6151
R1447 B.n353 B.n352 10.6151
R1448 B.n354 B.n353 10.6151
R1449 B.n354 B.n343 10.6151
R1450 B.n360 B.n343 10.6151
R1451 B.n361 B.n360 10.6151
R1452 B.n362 B.n361 10.6151
R1453 B.n362 B.n341 10.6151
R1454 B.n368 B.n341 10.6151
R1455 B.n369 B.n368 10.6151
R1456 B.n370 B.n369 10.6151
R1457 B.n370 B.n339 10.6151
R1458 B.n376 B.n339 10.6151
R1459 B.n377 B.n376 10.6151
R1460 B.n378 B.n377 10.6151
R1461 B.n378 B.n337 10.6151
R1462 B.n384 B.n337 10.6151
R1463 B.n385 B.n384 10.6151
R1464 B.n386 B.n385 10.6151
R1465 B.n386 B.n335 10.6151
R1466 B.n392 B.n335 10.6151
R1467 B.n393 B.n392 10.6151
R1468 B.n394 B.n393 10.6151
R1469 B.n394 B.n333 10.6151
R1470 B.n400 B.n333 10.6151
R1471 B.n401 B.n400 10.6151
R1472 B.n402 B.n401 10.6151
R1473 B.n402 B.n331 10.6151
R1474 B.n408 B.n331 10.6151
R1475 B.n409 B.n408 10.6151
R1476 B.n413 B.n409 10.6151
R1477 B.n419 B.n329 10.6151
R1478 B.n420 B.n419 10.6151
R1479 B.n421 B.n420 10.6151
R1480 B.n421 B.n327 10.6151
R1481 B.n427 B.n327 10.6151
R1482 B.n428 B.n427 10.6151
R1483 B.n429 B.n428 10.6151
R1484 B.n429 B.n325 10.6151
R1485 B.n435 B.n325 10.6151
R1486 B.n438 B.n437 10.6151
R1487 B.n438 B.n321 10.6151
R1488 B.n444 B.n321 10.6151
R1489 B.n445 B.n444 10.6151
R1490 B.n446 B.n445 10.6151
R1491 B.n446 B.n319 10.6151
R1492 B.n452 B.n319 10.6151
R1493 B.n453 B.n452 10.6151
R1494 B.n454 B.n453 10.6151
R1495 B.n454 B.n317 10.6151
R1496 B.n460 B.n317 10.6151
R1497 B.n461 B.n460 10.6151
R1498 B.n462 B.n461 10.6151
R1499 B.n462 B.n315 10.6151
R1500 B.n468 B.n315 10.6151
R1501 B.n469 B.n468 10.6151
R1502 B.n470 B.n469 10.6151
R1503 B.n470 B.n313 10.6151
R1504 B.n476 B.n313 10.6151
R1505 B.n477 B.n476 10.6151
R1506 B.n478 B.n477 10.6151
R1507 B.n478 B.n311 10.6151
R1508 B.n484 B.n311 10.6151
R1509 B.n485 B.n484 10.6151
R1510 B.n486 B.n485 10.6151
R1511 B.n486 B.n309 10.6151
R1512 B.n492 B.n309 10.6151
R1513 B.n493 B.n492 10.6151
R1514 B.n494 B.n493 10.6151
R1515 B.n494 B.n307 10.6151
R1516 B.n307 B.n306 10.6151
R1517 B.n501 B.n306 10.6151
R1518 B.n502 B.n501 10.6151
R1519 B.n503 B.n298 10.6151
R1520 B.n513 B.n298 10.6151
R1521 B.n514 B.n513 10.6151
R1522 B.n515 B.n514 10.6151
R1523 B.n515 B.n291 10.6151
R1524 B.n526 B.n291 10.6151
R1525 B.n527 B.n526 10.6151
R1526 B.n528 B.n527 10.6151
R1527 B.n528 B.n283 10.6151
R1528 B.n538 B.n283 10.6151
R1529 B.n539 B.n538 10.6151
R1530 B.n540 B.n539 10.6151
R1531 B.n540 B.n275 10.6151
R1532 B.n550 B.n275 10.6151
R1533 B.n551 B.n550 10.6151
R1534 B.n552 B.n551 10.6151
R1535 B.n552 B.n266 10.6151
R1536 B.n562 B.n266 10.6151
R1537 B.n563 B.n562 10.6151
R1538 B.n564 B.n563 10.6151
R1539 B.n564 B.n259 10.6151
R1540 B.n574 B.n259 10.6151
R1541 B.n575 B.n574 10.6151
R1542 B.n577 B.n575 10.6151
R1543 B.n577 B.n576 10.6151
R1544 B.n576 B.n251 10.6151
R1545 B.n588 B.n251 10.6151
R1546 B.n589 B.n588 10.6151
R1547 B.n590 B.n589 10.6151
R1548 B.n591 B.n590 10.6151
R1549 B.n592 B.n591 10.6151
R1550 B.n596 B.n592 10.6151
R1551 B.n597 B.n596 10.6151
R1552 B.n598 B.n597 10.6151
R1553 B.n599 B.n598 10.6151
R1554 B.n601 B.n599 10.6151
R1555 B.n602 B.n601 10.6151
R1556 B.n603 B.n602 10.6151
R1557 B.n604 B.n603 10.6151
R1558 B.n606 B.n604 10.6151
R1559 B.n607 B.n606 10.6151
R1560 B.n608 B.n607 10.6151
R1561 B.n609 B.n608 10.6151
R1562 B.n611 B.n609 10.6151
R1563 B.n612 B.n611 10.6151
R1564 B.n613 B.n612 10.6151
R1565 B.n614 B.n613 10.6151
R1566 B.n616 B.n614 10.6151
R1567 B.n617 B.n616 10.6151
R1568 B.n618 B.n617 10.6151
R1569 B.n619 B.n618 10.6151
R1570 B.n621 B.n619 10.6151
R1571 B.n622 B.n621 10.6151
R1572 B.n623 B.n622 10.6151
R1573 B.n624 B.n623 10.6151
R1574 B.n626 B.n624 10.6151
R1575 B.n627 B.n626 10.6151
R1576 B.n684 B.n1 10.6151
R1577 B.n684 B.n683 10.6151
R1578 B.n683 B.n682 10.6151
R1579 B.n682 B.n10 10.6151
R1580 B.n676 B.n10 10.6151
R1581 B.n676 B.n675 10.6151
R1582 B.n675 B.n674 10.6151
R1583 B.n674 B.n17 10.6151
R1584 B.n668 B.n17 10.6151
R1585 B.n668 B.n667 10.6151
R1586 B.n667 B.n666 10.6151
R1587 B.n666 B.n24 10.6151
R1588 B.n660 B.n24 10.6151
R1589 B.n660 B.n659 10.6151
R1590 B.n659 B.n658 10.6151
R1591 B.n658 B.n31 10.6151
R1592 B.n652 B.n31 10.6151
R1593 B.n652 B.n651 10.6151
R1594 B.n651 B.n650 10.6151
R1595 B.n650 B.n38 10.6151
R1596 B.n644 B.n38 10.6151
R1597 B.n644 B.n643 10.6151
R1598 B.n643 B.n642 10.6151
R1599 B.n642 B.n44 10.6151
R1600 B.n636 B.n44 10.6151
R1601 B.n636 B.n635 10.6151
R1602 B.n635 B.n634 10.6151
R1603 B.n100 B.n52 10.6151
R1604 B.n103 B.n100 10.6151
R1605 B.n104 B.n103 10.6151
R1606 B.n107 B.n104 10.6151
R1607 B.n108 B.n107 10.6151
R1608 B.n111 B.n108 10.6151
R1609 B.n112 B.n111 10.6151
R1610 B.n115 B.n112 10.6151
R1611 B.n116 B.n115 10.6151
R1612 B.n119 B.n116 10.6151
R1613 B.n120 B.n119 10.6151
R1614 B.n123 B.n120 10.6151
R1615 B.n124 B.n123 10.6151
R1616 B.n127 B.n124 10.6151
R1617 B.n128 B.n127 10.6151
R1618 B.n131 B.n128 10.6151
R1619 B.n132 B.n131 10.6151
R1620 B.n135 B.n132 10.6151
R1621 B.n136 B.n135 10.6151
R1622 B.n139 B.n136 10.6151
R1623 B.n140 B.n139 10.6151
R1624 B.n143 B.n140 10.6151
R1625 B.n144 B.n143 10.6151
R1626 B.n147 B.n144 10.6151
R1627 B.n148 B.n147 10.6151
R1628 B.n151 B.n148 10.6151
R1629 B.n152 B.n151 10.6151
R1630 B.n155 B.n152 10.6151
R1631 B.n156 B.n155 10.6151
R1632 B.n159 B.n156 10.6151
R1633 B.n160 B.n159 10.6151
R1634 B.n163 B.n160 10.6151
R1635 B.n164 B.n163 10.6151
R1636 B.n168 B.n167 10.6151
R1637 B.n171 B.n168 10.6151
R1638 B.n172 B.n171 10.6151
R1639 B.n175 B.n172 10.6151
R1640 B.n176 B.n175 10.6151
R1641 B.n179 B.n176 10.6151
R1642 B.n180 B.n179 10.6151
R1643 B.n183 B.n180 10.6151
R1644 B.n184 B.n183 10.6151
R1645 B.n188 B.n187 10.6151
R1646 B.n191 B.n188 10.6151
R1647 B.n192 B.n191 10.6151
R1648 B.n195 B.n192 10.6151
R1649 B.n196 B.n195 10.6151
R1650 B.n199 B.n196 10.6151
R1651 B.n200 B.n199 10.6151
R1652 B.n203 B.n200 10.6151
R1653 B.n204 B.n203 10.6151
R1654 B.n207 B.n204 10.6151
R1655 B.n208 B.n207 10.6151
R1656 B.n211 B.n208 10.6151
R1657 B.n212 B.n211 10.6151
R1658 B.n215 B.n212 10.6151
R1659 B.n216 B.n215 10.6151
R1660 B.n219 B.n216 10.6151
R1661 B.n220 B.n219 10.6151
R1662 B.n223 B.n220 10.6151
R1663 B.n224 B.n223 10.6151
R1664 B.n227 B.n224 10.6151
R1665 B.n228 B.n227 10.6151
R1666 B.n231 B.n228 10.6151
R1667 B.n232 B.n231 10.6151
R1668 B.n235 B.n232 10.6151
R1669 B.n236 B.n235 10.6151
R1670 B.n239 B.n236 10.6151
R1671 B.n240 B.n239 10.6151
R1672 B.n243 B.n240 10.6151
R1673 B.n244 B.n243 10.6151
R1674 B.n247 B.n244 10.6151
R1675 B.n249 B.n247 10.6151
R1676 B.n250 B.n249 10.6151
R1677 B.n628 B.n250 10.6151
R1678 B.n413 B.n412 9.36635
R1679 B.n437 B.n436 9.36635
R1680 B.n164 B.n99 9.36635
R1681 B.n187 B.n96 9.36635
R1682 B.n269 B.t0 8.97704
R1683 B.t1 B.n671 8.97704
R1684 B.n692 B.n0 8.11757
R1685 B.n692 B.n1 8.11757
R1686 B.n548 B.t2 1.49659
R1687 B.t5 B.n662 1.49659
R1688 B.n412 B.n329 1.24928
R1689 B.n436 B.n435 1.24928
R1690 B.n167 B.n99 1.24928
R1691 B.n184 B.n96 1.24928
R1692 VP.n7 VP.t4 195.463
R1693 VP.n15 VP.n14 173.534
R1694 VP.n27 VP.n26 173.534
R1695 VP.n13 VP.n12 173.534
R1696 VP.n8 VP.n5 161.3
R1697 VP.n10 VP.n9 161.3
R1698 VP.n11 VP.n4 161.3
R1699 VP.n25 VP.n0 161.3
R1700 VP.n24 VP.n23 161.3
R1701 VP.n22 VP.n1 161.3
R1702 VP.n21 VP.n20 161.3
R1703 VP.n19 VP.n2 161.3
R1704 VP.n18 VP.n17 161.3
R1705 VP.n16 VP.n3 161.3
R1706 VP.n20 VP.t5 160.044
R1707 VP.n14 VP.t3 160.044
R1708 VP.n26 VP.t0 160.044
R1709 VP.n6 VP.t2 160.044
R1710 VP.n12 VP.t1 160.044
R1711 VP.n19 VP.n18 52.6342
R1712 VP.n24 VP.n1 52.6342
R1713 VP.n10 VP.n5 52.6342
R1714 VP.n15 VP.n13 42.0422
R1715 VP.n7 VP.n6 41.826
R1716 VP.n18 VP.n3 28.3526
R1717 VP.n25 VP.n24 28.3526
R1718 VP.n11 VP.n10 28.3526
R1719 VP.n20 VP.n19 24.4675
R1720 VP.n20 VP.n1 24.4675
R1721 VP.n6 VP.n5 24.4675
R1722 VP.n8 VP.n7 17.5327
R1723 VP.n14 VP.n3 12.234
R1724 VP.n26 VP.n25 12.234
R1725 VP.n12 VP.n11 12.234
R1726 VP.n9 VP.n8 0.189894
R1727 VP.n9 VP.n4 0.189894
R1728 VP.n13 VP.n4 0.189894
R1729 VP.n16 VP.n15 0.189894
R1730 VP.n17 VP.n16 0.189894
R1731 VP.n17 VP.n2 0.189894
R1732 VP.n21 VP.n2 0.189894
R1733 VP.n22 VP.n21 0.189894
R1734 VP.n23 VP.n22 0.189894
R1735 VP.n23 VP.n0 0.189894
R1736 VP.n27 VP.n0 0.189894
R1737 VP VP.n27 0.0516364
R1738 VDD1.n44 VDD1.n0 289.615
R1739 VDD1.n93 VDD1.n49 289.615
R1740 VDD1.n45 VDD1.n44 185
R1741 VDD1.n43 VDD1.n42 185
R1742 VDD1.n4 VDD1.n3 185
R1743 VDD1.n8 VDD1.n6 185
R1744 VDD1.n37 VDD1.n36 185
R1745 VDD1.n35 VDD1.n34 185
R1746 VDD1.n10 VDD1.n9 185
R1747 VDD1.n29 VDD1.n28 185
R1748 VDD1.n27 VDD1.n26 185
R1749 VDD1.n14 VDD1.n13 185
R1750 VDD1.n21 VDD1.n20 185
R1751 VDD1.n19 VDD1.n18 185
R1752 VDD1.n66 VDD1.n65 185
R1753 VDD1.n68 VDD1.n67 185
R1754 VDD1.n61 VDD1.n60 185
R1755 VDD1.n74 VDD1.n73 185
R1756 VDD1.n76 VDD1.n75 185
R1757 VDD1.n57 VDD1.n56 185
R1758 VDD1.n83 VDD1.n82 185
R1759 VDD1.n84 VDD1.n55 185
R1760 VDD1.n86 VDD1.n85 185
R1761 VDD1.n53 VDD1.n52 185
R1762 VDD1.n92 VDD1.n91 185
R1763 VDD1.n94 VDD1.n93 185
R1764 VDD1.n17 VDD1.t1 149.524
R1765 VDD1.n64 VDD1.t2 149.524
R1766 VDD1.n44 VDD1.n43 104.615
R1767 VDD1.n43 VDD1.n3 104.615
R1768 VDD1.n8 VDD1.n3 104.615
R1769 VDD1.n36 VDD1.n8 104.615
R1770 VDD1.n36 VDD1.n35 104.615
R1771 VDD1.n35 VDD1.n9 104.615
R1772 VDD1.n28 VDD1.n9 104.615
R1773 VDD1.n28 VDD1.n27 104.615
R1774 VDD1.n27 VDD1.n13 104.615
R1775 VDD1.n20 VDD1.n13 104.615
R1776 VDD1.n20 VDD1.n19 104.615
R1777 VDD1.n67 VDD1.n66 104.615
R1778 VDD1.n67 VDD1.n60 104.615
R1779 VDD1.n74 VDD1.n60 104.615
R1780 VDD1.n75 VDD1.n74 104.615
R1781 VDD1.n75 VDD1.n56 104.615
R1782 VDD1.n83 VDD1.n56 104.615
R1783 VDD1.n84 VDD1.n83 104.615
R1784 VDD1.n85 VDD1.n84 104.615
R1785 VDD1.n85 VDD1.n52 104.615
R1786 VDD1.n92 VDD1.n52 104.615
R1787 VDD1.n93 VDD1.n92 104.615
R1788 VDD1.n99 VDD1.n98 67.0085
R1789 VDD1.n101 VDD1.n100 66.6867
R1790 VDD1 VDD1.n48 53.7386
R1791 VDD1.n99 VDD1.n97 53.6251
R1792 VDD1.n19 VDD1.t1 52.3082
R1793 VDD1.n66 VDD1.t2 52.3082
R1794 VDD1.n101 VDD1.n99 38.0849
R1795 VDD1.n6 VDD1.n4 13.1884
R1796 VDD1.n86 VDD1.n53 13.1884
R1797 VDD1.n42 VDD1.n41 12.8005
R1798 VDD1.n38 VDD1.n37 12.8005
R1799 VDD1.n87 VDD1.n55 12.8005
R1800 VDD1.n91 VDD1.n90 12.8005
R1801 VDD1.n45 VDD1.n2 12.0247
R1802 VDD1.n34 VDD1.n7 12.0247
R1803 VDD1.n82 VDD1.n81 12.0247
R1804 VDD1.n94 VDD1.n51 12.0247
R1805 VDD1.n46 VDD1.n0 11.249
R1806 VDD1.n33 VDD1.n10 11.249
R1807 VDD1.n80 VDD1.n57 11.249
R1808 VDD1.n95 VDD1.n49 11.249
R1809 VDD1.n30 VDD1.n29 10.4732
R1810 VDD1.n77 VDD1.n76 10.4732
R1811 VDD1.n18 VDD1.n17 10.2747
R1812 VDD1.n65 VDD1.n64 10.2747
R1813 VDD1.n26 VDD1.n12 9.69747
R1814 VDD1.n73 VDD1.n59 9.69747
R1815 VDD1.n48 VDD1.n47 9.45567
R1816 VDD1.n97 VDD1.n96 9.45567
R1817 VDD1.n16 VDD1.n15 9.3005
R1818 VDD1.n23 VDD1.n22 9.3005
R1819 VDD1.n25 VDD1.n24 9.3005
R1820 VDD1.n12 VDD1.n11 9.3005
R1821 VDD1.n31 VDD1.n30 9.3005
R1822 VDD1.n33 VDD1.n32 9.3005
R1823 VDD1.n7 VDD1.n5 9.3005
R1824 VDD1.n39 VDD1.n38 9.3005
R1825 VDD1.n47 VDD1.n46 9.3005
R1826 VDD1.n2 VDD1.n1 9.3005
R1827 VDD1.n41 VDD1.n40 9.3005
R1828 VDD1.n96 VDD1.n95 9.3005
R1829 VDD1.n51 VDD1.n50 9.3005
R1830 VDD1.n90 VDD1.n89 9.3005
R1831 VDD1.n63 VDD1.n62 9.3005
R1832 VDD1.n70 VDD1.n69 9.3005
R1833 VDD1.n72 VDD1.n71 9.3005
R1834 VDD1.n59 VDD1.n58 9.3005
R1835 VDD1.n78 VDD1.n77 9.3005
R1836 VDD1.n80 VDD1.n79 9.3005
R1837 VDD1.n81 VDD1.n54 9.3005
R1838 VDD1.n88 VDD1.n87 9.3005
R1839 VDD1.n25 VDD1.n14 8.92171
R1840 VDD1.n72 VDD1.n61 8.92171
R1841 VDD1.n22 VDD1.n21 8.14595
R1842 VDD1.n69 VDD1.n68 8.14595
R1843 VDD1.n18 VDD1.n16 7.3702
R1844 VDD1.n65 VDD1.n63 7.3702
R1845 VDD1.n21 VDD1.n16 5.81868
R1846 VDD1.n68 VDD1.n63 5.81868
R1847 VDD1.n22 VDD1.n14 5.04292
R1848 VDD1.n69 VDD1.n61 5.04292
R1849 VDD1.n26 VDD1.n25 4.26717
R1850 VDD1.n73 VDD1.n72 4.26717
R1851 VDD1.n29 VDD1.n12 3.49141
R1852 VDD1.n76 VDD1.n59 3.49141
R1853 VDD1.n17 VDD1.n15 2.84303
R1854 VDD1.n64 VDD1.n62 2.84303
R1855 VDD1.n48 VDD1.n0 2.71565
R1856 VDD1.n30 VDD1.n10 2.71565
R1857 VDD1.n77 VDD1.n57 2.71565
R1858 VDD1.n97 VDD1.n49 2.71565
R1859 VDD1.n100 VDD1.t3 2.10018
R1860 VDD1.n100 VDD1.t4 2.10018
R1861 VDD1.n98 VDD1.t0 2.10018
R1862 VDD1.n98 VDD1.t5 2.10018
R1863 VDD1.n46 VDD1.n45 1.93989
R1864 VDD1.n34 VDD1.n33 1.93989
R1865 VDD1.n82 VDD1.n80 1.93989
R1866 VDD1.n95 VDD1.n94 1.93989
R1867 VDD1.n42 VDD1.n2 1.16414
R1868 VDD1.n37 VDD1.n7 1.16414
R1869 VDD1.n81 VDD1.n55 1.16414
R1870 VDD1.n91 VDD1.n51 1.16414
R1871 VDD1.n41 VDD1.n4 0.388379
R1872 VDD1.n38 VDD1.n6 0.388379
R1873 VDD1.n87 VDD1.n86 0.388379
R1874 VDD1.n90 VDD1.n53 0.388379
R1875 VDD1 VDD1.n101 0.319466
R1876 VDD1.n47 VDD1.n1 0.155672
R1877 VDD1.n40 VDD1.n1 0.155672
R1878 VDD1.n40 VDD1.n39 0.155672
R1879 VDD1.n39 VDD1.n5 0.155672
R1880 VDD1.n32 VDD1.n5 0.155672
R1881 VDD1.n32 VDD1.n31 0.155672
R1882 VDD1.n31 VDD1.n11 0.155672
R1883 VDD1.n24 VDD1.n11 0.155672
R1884 VDD1.n24 VDD1.n23 0.155672
R1885 VDD1.n23 VDD1.n15 0.155672
R1886 VDD1.n70 VDD1.n62 0.155672
R1887 VDD1.n71 VDD1.n70 0.155672
R1888 VDD1.n71 VDD1.n58 0.155672
R1889 VDD1.n78 VDD1.n58 0.155672
R1890 VDD1.n79 VDD1.n78 0.155672
R1891 VDD1.n79 VDD1.n54 0.155672
R1892 VDD1.n88 VDD1.n54 0.155672
R1893 VDD1.n89 VDD1.n88 0.155672
R1894 VDD1.n89 VDD1.n50 0.155672
R1895 VDD1.n96 VDD1.n50 0.155672
C0 VP VDD1 4.82197f
C1 VN VDD1 0.149112f
C2 VP VDD2 0.358107f
C3 VN VDD2 4.61607f
C4 VP VTAIL 4.61957f
C5 VN VTAIL 4.60521f
C6 VDD2 VDD1 0.976436f
C7 VN VP 5.30359f
C8 VDD1 VTAIL 6.86552f
C9 VDD2 VTAIL 6.90757f
C10 VDD2 B 4.588096f
C11 VDD1 B 4.661616f
C12 VTAIL B 5.990814f
C13 VN B 9.301741f
C14 VP B 7.758371f
C15 VDD1.n0 B 0.031477f
C16 VDD1.n1 B 0.022076f
C17 VDD1.n2 B 0.011863f
C18 VDD1.n3 B 0.028039f
C19 VDD1.n4 B 0.012212f
C20 VDD1.n5 B 0.022076f
C21 VDD1.n6 B 0.012212f
C22 VDD1.n7 B 0.011863f
C23 VDD1.n8 B 0.028039f
C24 VDD1.n9 B 0.028039f
C25 VDD1.n10 B 0.012561f
C26 VDD1.n11 B 0.022076f
C27 VDD1.n12 B 0.011863f
C28 VDD1.n13 B 0.028039f
C29 VDD1.n14 B 0.012561f
C30 VDD1.n15 B 0.861344f
C31 VDD1.n16 B 0.011863f
C32 VDD1.t1 B 0.047056f
C33 VDD1.n17 B 0.137394f
C34 VDD1.n18 B 0.019822f
C35 VDD1.n19 B 0.02103f
C36 VDD1.n20 B 0.028039f
C37 VDD1.n21 B 0.012561f
C38 VDD1.n22 B 0.011863f
C39 VDD1.n23 B 0.022076f
C40 VDD1.n24 B 0.022076f
C41 VDD1.n25 B 0.011863f
C42 VDD1.n26 B 0.012561f
C43 VDD1.n27 B 0.028039f
C44 VDD1.n28 B 0.028039f
C45 VDD1.n29 B 0.012561f
C46 VDD1.n30 B 0.011863f
C47 VDD1.n31 B 0.022076f
C48 VDD1.n32 B 0.022076f
C49 VDD1.n33 B 0.011863f
C50 VDD1.n34 B 0.012561f
C51 VDD1.n35 B 0.028039f
C52 VDD1.n36 B 0.028039f
C53 VDD1.n37 B 0.012561f
C54 VDD1.n38 B 0.011863f
C55 VDD1.n39 B 0.022076f
C56 VDD1.n40 B 0.022076f
C57 VDD1.n41 B 0.011863f
C58 VDD1.n42 B 0.012561f
C59 VDD1.n43 B 0.028039f
C60 VDD1.n44 B 0.061491f
C61 VDD1.n45 B 0.012561f
C62 VDD1.n46 B 0.011863f
C63 VDD1.n47 B 0.056758f
C64 VDD1.n48 B 0.052746f
C65 VDD1.n49 B 0.031477f
C66 VDD1.n50 B 0.022076f
C67 VDD1.n51 B 0.011863f
C68 VDD1.n52 B 0.028039f
C69 VDD1.n53 B 0.012212f
C70 VDD1.n54 B 0.022076f
C71 VDD1.n55 B 0.012561f
C72 VDD1.n56 B 0.028039f
C73 VDD1.n57 B 0.012561f
C74 VDD1.n58 B 0.022076f
C75 VDD1.n59 B 0.011863f
C76 VDD1.n60 B 0.028039f
C77 VDD1.n61 B 0.012561f
C78 VDD1.n62 B 0.861344f
C79 VDD1.n63 B 0.011863f
C80 VDD1.t2 B 0.047056f
C81 VDD1.n64 B 0.137394f
C82 VDD1.n65 B 0.019822f
C83 VDD1.n66 B 0.02103f
C84 VDD1.n67 B 0.028039f
C85 VDD1.n68 B 0.012561f
C86 VDD1.n69 B 0.011863f
C87 VDD1.n70 B 0.022076f
C88 VDD1.n71 B 0.022076f
C89 VDD1.n72 B 0.011863f
C90 VDD1.n73 B 0.012561f
C91 VDD1.n74 B 0.028039f
C92 VDD1.n75 B 0.028039f
C93 VDD1.n76 B 0.012561f
C94 VDD1.n77 B 0.011863f
C95 VDD1.n78 B 0.022076f
C96 VDD1.n79 B 0.022076f
C97 VDD1.n80 B 0.011863f
C98 VDD1.n81 B 0.011863f
C99 VDD1.n82 B 0.012561f
C100 VDD1.n83 B 0.028039f
C101 VDD1.n84 B 0.028039f
C102 VDD1.n85 B 0.028039f
C103 VDD1.n86 B 0.012212f
C104 VDD1.n87 B 0.011863f
C105 VDD1.n88 B 0.022076f
C106 VDD1.n89 B 0.022076f
C107 VDD1.n90 B 0.011863f
C108 VDD1.n91 B 0.012561f
C109 VDD1.n92 B 0.028039f
C110 VDD1.n93 B 0.061491f
C111 VDD1.n94 B 0.012561f
C112 VDD1.n95 B 0.011863f
C113 VDD1.n96 B 0.056758f
C114 VDD1.n97 B 0.052324f
C115 VDD1.t0 B 0.16451f
C116 VDD1.t5 B 0.16451f
C117 VDD1.n98 B 1.44632f
C118 VDD1.n99 B 1.85587f
C119 VDD1.t3 B 0.16451f
C120 VDD1.t4 B 0.16451f
C121 VDD1.n100 B 1.44479f
C122 VDD1.n101 B 1.98824f
C123 VP.n0 B 0.034529f
C124 VP.t0 B 1.24996f
C125 VP.n1 B 0.061633f
C126 VP.n2 B 0.034529f
C127 VP.t5 B 1.24996f
C128 VP.n3 B 0.052125f
C129 VP.n4 B 0.034529f
C130 VP.t1 B 1.24996f
C131 VP.n5 B 0.061633f
C132 VP.t4 B 1.35744f
C133 VP.t2 B 1.24996f
C134 VP.n6 B 0.542712f
C135 VP.n7 B 0.532688f
C136 VP.n8 B 0.217648f
C137 VP.n9 B 0.034529f
C138 VP.n10 B 0.035529f
C139 VP.n11 B 0.052125f
C140 VP.n12 B 0.533551f
C141 VP.n13 B 1.43294f
C142 VP.t3 B 1.24996f
C143 VP.n14 B 0.533551f
C144 VP.n15 B 1.46246f
C145 VP.n16 B 0.034529f
C146 VP.n17 B 0.034529f
C147 VP.n18 B 0.035529f
C148 VP.n19 B 0.061633f
C149 VP.n20 B 0.496275f
C150 VP.n21 B 0.034529f
C151 VP.n22 B 0.034529f
C152 VP.n23 B 0.034529f
C153 VP.n24 B 0.035529f
C154 VP.n25 B 0.052125f
C155 VP.n26 B 0.533551f
C156 VP.n27 B 0.032057f
C157 VDD2.n0 B 0.031156f
C158 VDD2.n1 B 0.021851f
C159 VDD2.n2 B 0.011742f
C160 VDD2.n3 B 0.027754f
C161 VDD2.n4 B 0.012087f
C162 VDD2.n5 B 0.021851f
C163 VDD2.n6 B 0.012433f
C164 VDD2.n7 B 0.027754f
C165 VDD2.n8 B 0.012433f
C166 VDD2.n9 B 0.021851f
C167 VDD2.n10 B 0.011742f
C168 VDD2.n11 B 0.027754f
C169 VDD2.n12 B 0.012433f
C170 VDD2.n13 B 0.852561f
C171 VDD2.n14 B 0.011742f
C172 VDD2.t0 B 0.046576f
C173 VDD2.n15 B 0.135993f
C174 VDD2.n16 B 0.01962f
C175 VDD2.n17 B 0.020815f
C176 VDD2.n18 B 0.027754f
C177 VDD2.n19 B 0.012433f
C178 VDD2.n20 B 0.011742f
C179 VDD2.n21 B 0.021851f
C180 VDD2.n22 B 0.021851f
C181 VDD2.n23 B 0.011742f
C182 VDD2.n24 B 0.012433f
C183 VDD2.n25 B 0.027754f
C184 VDD2.n26 B 0.027754f
C185 VDD2.n27 B 0.012433f
C186 VDD2.n28 B 0.011742f
C187 VDD2.n29 B 0.021851f
C188 VDD2.n30 B 0.021851f
C189 VDD2.n31 B 0.011742f
C190 VDD2.n32 B 0.011742f
C191 VDD2.n33 B 0.012433f
C192 VDD2.n34 B 0.027754f
C193 VDD2.n35 B 0.027754f
C194 VDD2.n36 B 0.027754f
C195 VDD2.n37 B 0.012087f
C196 VDD2.n38 B 0.011742f
C197 VDD2.n39 B 0.021851f
C198 VDD2.n40 B 0.021851f
C199 VDD2.n41 B 0.011742f
C200 VDD2.n42 B 0.012433f
C201 VDD2.n43 B 0.027754f
C202 VDD2.n44 B 0.060864f
C203 VDD2.n45 B 0.012433f
C204 VDD2.n46 B 0.011742f
C205 VDD2.n47 B 0.05618f
C206 VDD2.n48 B 0.05179f
C207 VDD2.t4 B 0.162832f
C208 VDD2.t5 B 0.162832f
C209 VDD2.n49 B 1.43157f
C210 VDD2.n50 B 1.75583f
C211 VDD2.n51 B 0.031156f
C212 VDD2.n52 B 0.021851f
C213 VDD2.n53 B 0.011742f
C214 VDD2.n54 B 0.027754f
C215 VDD2.n55 B 0.012087f
C216 VDD2.n56 B 0.021851f
C217 VDD2.n57 B 0.012087f
C218 VDD2.n58 B 0.011742f
C219 VDD2.n59 B 0.027754f
C220 VDD2.n60 B 0.027754f
C221 VDD2.n61 B 0.012433f
C222 VDD2.n62 B 0.021851f
C223 VDD2.n63 B 0.011742f
C224 VDD2.n64 B 0.027754f
C225 VDD2.n65 B 0.012433f
C226 VDD2.n66 B 0.852561f
C227 VDD2.n67 B 0.011742f
C228 VDD2.t2 B 0.046576f
C229 VDD2.n68 B 0.135993f
C230 VDD2.n69 B 0.01962f
C231 VDD2.n70 B 0.020815f
C232 VDD2.n71 B 0.027754f
C233 VDD2.n72 B 0.012433f
C234 VDD2.n73 B 0.011742f
C235 VDD2.n74 B 0.021851f
C236 VDD2.n75 B 0.021851f
C237 VDD2.n76 B 0.011742f
C238 VDD2.n77 B 0.012433f
C239 VDD2.n78 B 0.027754f
C240 VDD2.n79 B 0.027754f
C241 VDD2.n80 B 0.012433f
C242 VDD2.n81 B 0.011742f
C243 VDD2.n82 B 0.021851f
C244 VDD2.n83 B 0.021851f
C245 VDD2.n84 B 0.011742f
C246 VDD2.n85 B 0.012433f
C247 VDD2.n86 B 0.027754f
C248 VDD2.n87 B 0.027754f
C249 VDD2.n88 B 0.012433f
C250 VDD2.n89 B 0.011742f
C251 VDD2.n90 B 0.021851f
C252 VDD2.n91 B 0.021851f
C253 VDD2.n92 B 0.011742f
C254 VDD2.n93 B 0.012433f
C255 VDD2.n94 B 0.027754f
C256 VDD2.n95 B 0.060864f
C257 VDD2.n96 B 0.012433f
C258 VDD2.n97 B 0.011742f
C259 VDD2.n98 B 0.05618f
C260 VDD2.n99 B 0.049351f
C261 VDD2.n100 B 1.78507f
C262 VDD2.t3 B 0.162832f
C263 VDD2.t1 B 0.162832f
C264 VDD2.n101 B 1.43155f
C265 VTAIL.t7 B 0.178426f
C266 VTAIL.t6 B 0.178426f
C267 VTAIL.n0 B 1.50461f
C268 VTAIL.n1 B 0.349555f
C269 VTAIL.n2 B 0.03414f
C270 VTAIL.n3 B 0.023944f
C271 VTAIL.n4 B 0.012866f
C272 VTAIL.n5 B 0.030411f
C273 VTAIL.n6 B 0.013245f
C274 VTAIL.n7 B 0.023944f
C275 VTAIL.n8 B 0.013623f
C276 VTAIL.n9 B 0.030411f
C277 VTAIL.n10 B 0.013623f
C278 VTAIL.n11 B 0.023944f
C279 VTAIL.n12 B 0.012866f
C280 VTAIL.n13 B 0.030411f
C281 VTAIL.n14 B 0.013623f
C282 VTAIL.n15 B 0.934208f
C283 VTAIL.n16 B 0.012866f
C284 VTAIL.t11 B 0.051036f
C285 VTAIL.n17 B 0.149016f
C286 VTAIL.n18 B 0.021498f
C287 VTAIL.n19 B 0.022808f
C288 VTAIL.n20 B 0.030411f
C289 VTAIL.n21 B 0.013623f
C290 VTAIL.n22 B 0.012866f
C291 VTAIL.n23 B 0.023944f
C292 VTAIL.n24 B 0.023944f
C293 VTAIL.n25 B 0.012866f
C294 VTAIL.n26 B 0.013623f
C295 VTAIL.n27 B 0.030411f
C296 VTAIL.n28 B 0.030411f
C297 VTAIL.n29 B 0.013623f
C298 VTAIL.n30 B 0.012866f
C299 VTAIL.n31 B 0.023944f
C300 VTAIL.n32 B 0.023944f
C301 VTAIL.n33 B 0.012866f
C302 VTAIL.n34 B 0.012866f
C303 VTAIL.n35 B 0.013623f
C304 VTAIL.n36 B 0.030411f
C305 VTAIL.n37 B 0.030411f
C306 VTAIL.n38 B 0.030411f
C307 VTAIL.n39 B 0.013245f
C308 VTAIL.n40 B 0.012866f
C309 VTAIL.n41 B 0.023944f
C310 VTAIL.n42 B 0.023944f
C311 VTAIL.n43 B 0.012866f
C312 VTAIL.n44 B 0.013623f
C313 VTAIL.n45 B 0.030411f
C314 VTAIL.n46 B 0.066693f
C315 VTAIL.n47 B 0.013623f
C316 VTAIL.n48 B 0.012866f
C317 VTAIL.n49 B 0.06156f
C318 VTAIL.n50 B 0.037587f
C319 VTAIL.n51 B 0.234805f
C320 VTAIL.t2 B 0.178426f
C321 VTAIL.t0 B 0.178426f
C322 VTAIL.n52 B 1.50461f
C323 VTAIL.n53 B 1.52315f
C324 VTAIL.t5 B 0.178426f
C325 VTAIL.t9 B 0.178426f
C326 VTAIL.n54 B 1.50462f
C327 VTAIL.n55 B 1.52314f
C328 VTAIL.n56 B 0.03414f
C329 VTAIL.n57 B 0.023944f
C330 VTAIL.n58 B 0.012866f
C331 VTAIL.n59 B 0.030411f
C332 VTAIL.n60 B 0.013245f
C333 VTAIL.n61 B 0.023944f
C334 VTAIL.n62 B 0.013245f
C335 VTAIL.n63 B 0.012866f
C336 VTAIL.n64 B 0.030411f
C337 VTAIL.n65 B 0.030411f
C338 VTAIL.n66 B 0.013623f
C339 VTAIL.n67 B 0.023944f
C340 VTAIL.n68 B 0.012866f
C341 VTAIL.n69 B 0.030411f
C342 VTAIL.n70 B 0.013623f
C343 VTAIL.n71 B 0.934208f
C344 VTAIL.n72 B 0.012866f
C345 VTAIL.t4 B 0.051036f
C346 VTAIL.n73 B 0.149016f
C347 VTAIL.n74 B 0.021498f
C348 VTAIL.n75 B 0.022808f
C349 VTAIL.n76 B 0.030411f
C350 VTAIL.n77 B 0.013623f
C351 VTAIL.n78 B 0.012866f
C352 VTAIL.n79 B 0.023944f
C353 VTAIL.n80 B 0.023944f
C354 VTAIL.n81 B 0.012866f
C355 VTAIL.n82 B 0.013623f
C356 VTAIL.n83 B 0.030411f
C357 VTAIL.n84 B 0.030411f
C358 VTAIL.n85 B 0.013623f
C359 VTAIL.n86 B 0.012866f
C360 VTAIL.n87 B 0.023944f
C361 VTAIL.n88 B 0.023944f
C362 VTAIL.n89 B 0.012866f
C363 VTAIL.n90 B 0.013623f
C364 VTAIL.n91 B 0.030411f
C365 VTAIL.n92 B 0.030411f
C366 VTAIL.n93 B 0.013623f
C367 VTAIL.n94 B 0.012866f
C368 VTAIL.n95 B 0.023944f
C369 VTAIL.n96 B 0.023944f
C370 VTAIL.n97 B 0.012866f
C371 VTAIL.n98 B 0.013623f
C372 VTAIL.n99 B 0.030411f
C373 VTAIL.n100 B 0.066693f
C374 VTAIL.n101 B 0.013623f
C375 VTAIL.n102 B 0.012866f
C376 VTAIL.n103 B 0.06156f
C377 VTAIL.n104 B 0.037587f
C378 VTAIL.n105 B 0.234805f
C379 VTAIL.t3 B 0.178426f
C380 VTAIL.t1 B 0.178426f
C381 VTAIL.n106 B 1.50462f
C382 VTAIL.n107 B 0.432352f
C383 VTAIL.n108 B 0.03414f
C384 VTAIL.n109 B 0.023944f
C385 VTAIL.n110 B 0.012866f
C386 VTAIL.n111 B 0.030411f
C387 VTAIL.n112 B 0.013245f
C388 VTAIL.n113 B 0.023944f
C389 VTAIL.n114 B 0.013245f
C390 VTAIL.n115 B 0.012866f
C391 VTAIL.n116 B 0.030411f
C392 VTAIL.n117 B 0.030411f
C393 VTAIL.n118 B 0.013623f
C394 VTAIL.n119 B 0.023944f
C395 VTAIL.n120 B 0.012866f
C396 VTAIL.n121 B 0.030411f
C397 VTAIL.n122 B 0.013623f
C398 VTAIL.n123 B 0.934208f
C399 VTAIL.n124 B 0.012866f
C400 VTAIL.t10 B 0.051036f
C401 VTAIL.n125 B 0.149016f
C402 VTAIL.n126 B 0.021498f
C403 VTAIL.n127 B 0.022808f
C404 VTAIL.n128 B 0.030411f
C405 VTAIL.n129 B 0.013623f
C406 VTAIL.n130 B 0.012866f
C407 VTAIL.n131 B 0.023944f
C408 VTAIL.n132 B 0.023944f
C409 VTAIL.n133 B 0.012866f
C410 VTAIL.n134 B 0.013623f
C411 VTAIL.n135 B 0.030411f
C412 VTAIL.n136 B 0.030411f
C413 VTAIL.n137 B 0.013623f
C414 VTAIL.n138 B 0.012866f
C415 VTAIL.n139 B 0.023944f
C416 VTAIL.n140 B 0.023944f
C417 VTAIL.n141 B 0.012866f
C418 VTAIL.n142 B 0.013623f
C419 VTAIL.n143 B 0.030411f
C420 VTAIL.n144 B 0.030411f
C421 VTAIL.n145 B 0.013623f
C422 VTAIL.n146 B 0.012866f
C423 VTAIL.n147 B 0.023944f
C424 VTAIL.n148 B 0.023944f
C425 VTAIL.n149 B 0.012866f
C426 VTAIL.n150 B 0.013623f
C427 VTAIL.n151 B 0.030411f
C428 VTAIL.n152 B 0.066693f
C429 VTAIL.n153 B 0.013623f
C430 VTAIL.n154 B 0.012866f
C431 VTAIL.n155 B 0.06156f
C432 VTAIL.n156 B 0.037587f
C433 VTAIL.n157 B 1.2092f
C434 VTAIL.n158 B 0.03414f
C435 VTAIL.n159 B 0.023944f
C436 VTAIL.n160 B 0.012866f
C437 VTAIL.n161 B 0.030411f
C438 VTAIL.n162 B 0.013245f
C439 VTAIL.n163 B 0.023944f
C440 VTAIL.n164 B 0.013623f
C441 VTAIL.n165 B 0.030411f
C442 VTAIL.n166 B 0.013623f
C443 VTAIL.n167 B 0.023944f
C444 VTAIL.n168 B 0.012866f
C445 VTAIL.n169 B 0.030411f
C446 VTAIL.n170 B 0.013623f
C447 VTAIL.n171 B 0.934208f
C448 VTAIL.n172 B 0.012866f
C449 VTAIL.t8 B 0.051036f
C450 VTAIL.n173 B 0.149016f
C451 VTAIL.n174 B 0.021498f
C452 VTAIL.n175 B 0.022808f
C453 VTAIL.n176 B 0.030411f
C454 VTAIL.n177 B 0.013623f
C455 VTAIL.n178 B 0.012866f
C456 VTAIL.n179 B 0.023944f
C457 VTAIL.n180 B 0.023944f
C458 VTAIL.n181 B 0.012866f
C459 VTAIL.n182 B 0.013623f
C460 VTAIL.n183 B 0.030411f
C461 VTAIL.n184 B 0.030411f
C462 VTAIL.n185 B 0.013623f
C463 VTAIL.n186 B 0.012866f
C464 VTAIL.n187 B 0.023944f
C465 VTAIL.n188 B 0.023944f
C466 VTAIL.n189 B 0.012866f
C467 VTAIL.n190 B 0.012866f
C468 VTAIL.n191 B 0.013623f
C469 VTAIL.n192 B 0.030411f
C470 VTAIL.n193 B 0.030411f
C471 VTAIL.n194 B 0.030411f
C472 VTAIL.n195 B 0.013245f
C473 VTAIL.n196 B 0.012866f
C474 VTAIL.n197 B 0.023944f
C475 VTAIL.n198 B 0.023944f
C476 VTAIL.n199 B 0.012866f
C477 VTAIL.n200 B 0.013623f
C478 VTAIL.n201 B 0.030411f
C479 VTAIL.n202 B 0.066693f
C480 VTAIL.n203 B 0.013623f
C481 VTAIL.n204 B 0.012866f
C482 VTAIL.n205 B 0.06156f
C483 VTAIL.n206 B 0.037587f
C484 VTAIL.n207 B 1.17561f
C485 VN.n0 B 0.033947f
C486 VN.t0 B 1.2289f
C487 VN.n1 B 0.060594f
C488 VN.t5 B 1.33456f
C489 VN.t1 B 1.2289f
C490 VN.n2 B 0.533567f
C491 VN.n3 B 0.523711f
C492 VN.n4 B 0.21398f
C493 VN.n5 B 0.033947f
C494 VN.n6 B 0.03493f
C495 VN.n7 B 0.051246f
C496 VN.n8 B 0.524559f
C497 VN.n9 B 0.031517f
C498 VN.n10 B 0.033947f
C499 VN.t3 B 1.2289f
C500 VN.n11 B 0.060594f
C501 VN.t4 B 1.33456f
C502 VN.t2 B 1.2289f
C503 VN.n12 B 0.533567f
C504 VN.n13 B 0.523711f
C505 VN.n14 B 0.21398f
C506 VN.n15 B 0.033947f
C507 VN.n16 B 0.03493f
C508 VN.n17 B 0.051246f
C509 VN.n18 B 0.524559f
C510 VN.n19 B 1.43107f
.ends

