* NGSPICE file created from diff_pair_sample_1590.ext - technology: sky130A

.subckt diff_pair_sample_1590 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=4.8906 pd=25.86 as=2.0691 ps=12.87 w=12.54 l=3.97
X1 VDD1.t3 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.0691 pd=12.87 as=4.8906 ps=25.86 w=12.54 l=3.97
X2 VTAIL.t1 VP.t1 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=4.8906 pd=25.86 as=2.0691 ps=12.87 w=12.54 l=3.97
X3 VTAIL.t2 VP.t2 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=4.8906 pd=25.86 as=2.0691 ps=12.87 w=12.54 l=3.97
X4 VDD1.t0 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.0691 pd=12.87 as=4.8906 ps=25.86 w=12.54 l=3.97
X5 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=4.8906 pd=25.86 as=0 ps=0 w=12.54 l=3.97
X6 VDD2.t0 VN.t1 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=2.0691 pd=12.87 as=4.8906 ps=25.86 w=12.54 l=3.97
X7 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=4.8906 pd=25.86 as=0 ps=0 w=12.54 l=3.97
X8 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.8906 pd=25.86 as=0 ps=0 w=12.54 l=3.97
X9 VDD2.t3 VN.t2 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.0691 pd=12.87 as=4.8906 ps=25.86 w=12.54 l=3.97
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=4.8906 pd=25.86 as=0 ps=0 w=12.54 l=3.97
X11 VTAIL.t4 VN.t3 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=4.8906 pd=25.86 as=2.0691 ps=12.87 w=12.54 l=3.97
R0 VN.n0 VN.t3 110.007
R1 VN.n1 VN.t1 110.007
R2 VN.n0 VN.t2 108.569
R3 VN.n1 VN.t0 108.569
R4 VN VN.n1 52.8154
R5 VN VN.n0 1.74345
R6 VDD2.n2 VDD2.n0 108.597
R7 VDD2.n2 VDD2.n1 62.951
R8 VDD2.n1 VDD2.t1 1.57945
R9 VDD2.n1 VDD2.t0 1.57945
R10 VDD2.n0 VDD2.t2 1.57945
R11 VDD2.n0 VDD2.t3 1.57945
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t1 47.8513
R14 VTAIL.n4 VTAIL.t6 47.8513
R15 VTAIL.n3 VTAIL.t7 47.8513
R16 VTAIL.n7 VTAIL.t5 47.8511
R17 VTAIL.n0 VTAIL.t4 47.8511
R18 VTAIL.n1 VTAIL.t0 47.8511
R19 VTAIL.n2 VTAIL.t2 47.8511
R20 VTAIL.n6 VTAIL.t3 47.8511
R21 VTAIL.n7 VTAIL.n6 26.8841
R22 VTAIL.n3 VTAIL.n2 26.8841
R23 VTAIL.n4 VTAIL.n3 3.7074
R24 VTAIL.n6 VTAIL.n5 3.7074
R25 VTAIL.n2 VTAIL.n1 3.7074
R26 VTAIL VTAIL.n0 1.91214
R27 VTAIL VTAIL.n7 1.79576
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 B.n671 B.n670 585
R31 B.n673 B.n138 585
R32 B.n676 B.n675 585
R33 B.n677 B.n137 585
R34 B.n679 B.n678 585
R35 B.n681 B.n136 585
R36 B.n684 B.n683 585
R37 B.n685 B.n135 585
R38 B.n687 B.n686 585
R39 B.n689 B.n134 585
R40 B.n692 B.n691 585
R41 B.n693 B.n133 585
R42 B.n695 B.n694 585
R43 B.n697 B.n132 585
R44 B.n700 B.n699 585
R45 B.n701 B.n131 585
R46 B.n703 B.n702 585
R47 B.n705 B.n130 585
R48 B.n708 B.n707 585
R49 B.n709 B.n129 585
R50 B.n711 B.n710 585
R51 B.n713 B.n128 585
R52 B.n716 B.n715 585
R53 B.n717 B.n127 585
R54 B.n719 B.n718 585
R55 B.n721 B.n126 585
R56 B.n724 B.n723 585
R57 B.n725 B.n125 585
R58 B.n727 B.n726 585
R59 B.n729 B.n124 585
R60 B.n732 B.n731 585
R61 B.n733 B.n123 585
R62 B.n735 B.n734 585
R63 B.n737 B.n122 585
R64 B.n740 B.n739 585
R65 B.n741 B.n121 585
R66 B.n743 B.n742 585
R67 B.n745 B.n120 585
R68 B.n748 B.n747 585
R69 B.n749 B.n119 585
R70 B.n751 B.n750 585
R71 B.n753 B.n118 585
R72 B.n756 B.n755 585
R73 B.n758 B.n115 585
R74 B.n760 B.n759 585
R75 B.n762 B.n114 585
R76 B.n765 B.n764 585
R77 B.n766 B.n113 585
R78 B.n768 B.n767 585
R79 B.n770 B.n112 585
R80 B.n773 B.n772 585
R81 B.n774 B.n108 585
R82 B.n776 B.n775 585
R83 B.n778 B.n107 585
R84 B.n781 B.n780 585
R85 B.n782 B.n106 585
R86 B.n784 B.n783 585
R87 B.n786 B.n105 585
R88 B.n789 B.n788 585
R89 B.n790 B.n104 585
R90 B.n792 B.n791 585
R91 B.n794 B.n103 585
R92 B.n797 B.n796 585
R93 B.n798 B.n102 585
R94 B.n800 B.n799 585
R95 B.n802 B.n101 585
R96 B.n805 B.n804 585
R97 B.n806 B.n100 585
R98 B.n808 B.n807 585
R99 B.n810 B.n99 585
R100 B.n813 B.n812 585
R101 B.n814 B.n98 585
R102 B.n816 B.n815 585
R103 B.n818 B.n97 585
R104 B.n821 B.n820 585
R105 B.n822 B.n96 585
R106 B.n824 B.n823 585
R107 B.n826 B.n95 585
R108 B.n829 B.n828 585
R109 B.n830 B.n94 585
R110 B.n832 B.n831 585
R111 B.n834 B.n93 585
R112 B.n837 B.n836 585
R113 B.n838 B.n92 585
R114 B.n840 B.n839 585
R115 B.n842 B.n91 585
R116 B.n845 B.n844 585
R117 B.n846 B.n90 585
R118 B.n848 B.n847 585
R119 B.n850 B.n89 585
R120 B.n853 B.n852 585
R121 B.n854 B.n88 585
R122 B.n856 B.n855 585
R123 B.n858 B.n87 585
R124 B.n861 B.n860 585
R125 B.n862 B.n86 585
R126 B.n669 B.n84 585
R127 B.n865 B.n84 585
R128 B.n668 B.n83 585
R129 B.n866 B.n83 585
R130 B.n667 B.n82 585
R131 B.n867 B.n82 585
R132 B.n666 B.n665 585
R133 B.n665 B.n78 585
R134 B.n664 B.n77 585
R135 B.n873 B.n77 585
R136 B.n663 B.n76 585
R137 B.n874 B.n76 585
R138 B.n662 B.n75 585
R139 B.n875 B.n75 585
R140 B.n661 B.n660 585
R141 B.n660 B.n71 585
R142 B.n659 B.n70 585
R143 B.n881 B.n70 585
R144 B.n658 B.n69 585
R145 B.n882 B.n69 585
R146 B.n657 B.n68 585
R147 B.n883 B.n68 585
R148 B.n656 B.n655 585
R149 B.n655 B.n64 585
R150 B.n654 B.n63 585
R151 B.n889 B.n63 585
R152 B.n653 B.n62 585
R153 B.n890 B.n62 585
R154 B.n652 B.n61 585
R155 B.n891 B.n61 585
R156 B.n651 B.n650 585
R157 B.n650 B.n57 585
R158 B.n649 B.n56 585
R159 B.n897 B.n56 585
R160 B.n648 B.n55 585
R161 B.n898 B.n55 585
R162 B.n647 B.n54 585
R163 B.n899 B.n54 585
R164 B.n646 B.n645 585
R165 B.n645 B.n50 585
R166 B.n644 B.n49 585
R167 B.n905 B.n49 585
R168 B.n643 B.n48 585
R169 B.n906 B.n48 585
R170 B.n642 B.n47 585
R171 B.n907 B.n47 585
R172 B.n641 B.n640 585
R173 B.n640 B.n43 585
R174 B.n639 B.n42 585
R175 B.n913 B.n42 585
R176 B.n638 B.n41 585
R177 B.n914 B.n41 585
R178 B.n637 B.n40 585
R179 B.n915 B.n40 585
R180 B.n636 B.n635 585
R181 B.n635 B.n36 585
R182 B.n634 B.n35 585
R183 B.n921 B.n35 585
R184 B.n633 B.n34 585
R185 B.n922 B.n34 585
R186 B.n632 B.n33 585
R187 B.n923 B.n33 585
R188 B.n631 B.n630 585
R189 B.n630 B.n29 585
R190 B.n629 B.n28 585
R191 B.n929 B.n28 585
R192 B.n628 B.n27 585
R193 B.n930 B.n27 585
R194 B.n627 B.n26 585
R195 B.n931 B.n26 585
R196 B.n626 B.n625 585
R197 B.n625 B.n22 585
R198 B.n624 B.n21 585
R199 B.n937 B.n21 585
R200 B.n623 B.n20 585
R201 B.n938 B.n20 585
R202 B.n622 B.n19 585
R203 B.n939 B.n19 585
R204 B.n621 B.n620 585
R205 B.n620 B.n15 585
R206 B.n619 B.n14 585
R207 B.n945 B.n14 585
R208 B.n618 B.n13 585
R209 B.n946 B.n13 585
R210 B.n617 B.n12 585
R211 B.n947 B.n12 585
R212 B.n616 B.n615 585
R213 B.n615 B.n8 585
R214 B.n614 B.n7 585
R215 B.n953 B.n7 585
R216 B.n613 B.n6 585
R217 B.n954 B.n6 585
R218 B.n612 B.n5 585
R219 B.n955 B.n5 585
R220 B.n611 B.n610 585
R221 B.n610 B.n4 585
R222 B.n609 B.n139 585
R223 B.n609 B.n608 585
R224 B.n599 B.n140 585
R225 B.n141 B.n140 585
R226 B.n601 B.n600 585
R227 B.n602 B.n601 585
R228 B.n598 B.n146 585
R229 B.n146 B.n145 585
R230 B.n597 B.n596 585
R231 B.n596 B.n595 585
R232 B.n148 B.n147 585
R233 B.n149 B.n148 585
R234 B.n588 B.n587 585
R235 B.n589 B.n588 585
R236 B.n586 B.n154 585
R237 B.n154 B.n153 585
R238 B.n585 B.n584 585
R239 B.n584 B.n583 585
R240 B.n156 B.n155 585
R241 B.n157 B.n156 585
R242 B.n576 B.n575 585
R243 B.n577 B.n576 585
R244 B.n574 B.n162 585
R245 B.n162 B.n161 585
R246 B.n573 B.n572 585
R247 B.n572 B.n571 585
R248 B.n164 B.n163 585
R249 B.n165 B.n164 585
R250 B.n564 B.n563 585
R251 B.n565 B.n564 585
R252 B.n562 B.n170 585
R253 B.n170 B.n169 585
R254 B.n561 B.n560 585
R255 B.n560 B.n559 585
R256 B.n172 B.n171 585
R257 B.n173 B.n172 585
R258 B.n552 B.n551 585
R259 B.n553 B.n552 585
R260 B.n550 B.n177 585
R261 B.n181 B.n177 585
R262 B.n549 B.n548 585
R263 B.n548 B.n547 585
R264 B.n179 B.n178 585
R265 B.n180 B.n179 585
R266 B.n540 B.n539 585
R267 B.n541 B.n540 585
R268 B.n538 B.n186 585
R269 B.n186 B.n185 585
R270 B.n537 B.n536 585
R271 B.n536 B.n535 585
R272 B.n188 B.n187 585
R273 B.n189 B.n188 585
R274 B.n528 B.n527 585
R275 B.n529 B.n528 585
R276 B.n526 B.n194 585
R277 B.n194 B.n193 585
R278 B.n525 B.n524 585
R279 B.n524 B.n523 585
R280 B.n196 B.n195 585
R281 B.n197 B.n196 585
R282 B.n516 B.n515 585
R283 B.n517 B.n516 585
R284 B.n514 B.n202 585
R285 B.n202 B.n201 585
R286 B.n513 B.n512 585
R287 B.n512 B.n511 585
R288 B.n204 B.n203 585
R289 B.n205 B.n204 585
R290 B.n504 B.n503 585
R291 B.n505 B.n504 585
R292 B.n502 B.n209 585
R293 B.n213 B.n209 585
R294 B.n501 B.n500 585
R295 B.n500 B.n499 585
R296 B.n211 B.n210 585
R297 B.n212 B.n211 585
R298 B.n492 B.n491 585
R299 B.n493 B.n492 585
R300 B.n490 B.n218 585
R301 B.n218 B.n217 585
R302 B.n489 B.n488 585
R303 B.n488 B.n487 585
R304 B.n220 B.n219 585
R305 B.n221 B.n220 585
R306 B.n480 B.n479 585
R307 B.n481 B.n480 585
R308 B.n478 B.n226 585
R309 B.n226 B.n225 585
R310 B.n477 B.n476 585
R311 B.n476 B.n475 585
R312 B.n472 B.n230 585
R313 B.n471 B.n470 585
R314 B.n468 B.n231 585
R315 B.n468 B.n229 585
R316 B.n467 B.n466 585
R317 B.n465 B.n464 585
R318 B.n463 B.n233 585
R319 B.n461 B.n460 585
R320 B.n459 B.n234 585
R321 B.n458 B.n457 585
R322 B.n455 B.n235 585
R323 B.n453 B.n452 585
R324 B.n451 B.n236 585
R325 B.n450 B.n449 585
R326 B.n447 B.n237 585
R327 B.n445 B.n444 585
R328 B.n443 B.n238 585
R329 B.n442 B.n441 585
R330 B.n439 B.n239 585
R331 B.n437 B.n436 585
R332 B.n435 B.n240 585
R333 B.n434 B.n433 585
R334 B.n431 B.n241 585
R335 B.n429 B.n428 585
R336 B.n427 B.n242 585
R337 B.n426 B.n425 585
R338 B.n423 B.n243 585
R339 B.n421 B.n420 585
R340 B.n419 B.n244 585
R341 B.n418 B.n417 585
R342 B.n415 B.n245 585
R343 B.n413 B.n412 585
R344 B.n411 B.n246 585
R345 B.n410 B.n409 585
R346 B.n407 B.n247 585
R347 B.n405 B.n404 585
R348 B.n403 B.n248 585
R349 B.n402 B.n401 585
R350 B.n399 B.n249 585
R351 B.n397 B.n396 585
R352 B.n395 B.n250 585
R353 B.n394 B.n393 585
R354 B.n391 B.n251 585
R355 B.n389 B.n388 585
R356 B.n386 B.n252 585
R357 B.n385 B.n384 585
R358 B.n382 B.n255 585
R359 B.n380 B.n379 585
R360 B.n378 B.n256 585
R361 B.n377 B.n376 585
R362 B.n374 B.n257 585
R363 B.n372 B.n371 585
R364 B.n370 B.n258 585
R365 B.n369 B.n368 585
R366 B.n366 B.n365 585
R367 B.n364 B.n363 585
R368 B.n362 B.n263 585
R369 B.n360 B.n359 585
R370 B.n358 B.n264 585
R371 B.n357 B.n356 585
R372 B.n354 B.n265 585
R373 B.n352 B.n351 585
R374 B.n350 B.n266 585
R375 B.n349 B.n348 585
R376 B.n346 B.n267 585
R377 B.n344 B.n343 585
R378 B.n342 B.n268 585
R379 B.n341 B.n340 585
R380 B.n338 B.n269 585
R381 B.n336 B.n335 585
R382 B.n334 B.n270 585
R383 B.n333 B.n332 585
R384 B.n330 B.n271 585
R385 B.n328 B.n327 585
R386 B.n326 B.n272 585
R387 B.n325 B.n324 585
R388 B.n322 B.n273 585
R389 B.n320 B.n319 585
R390 B.n318 B.n274 585
R391 B.n317 B.n316 585
R392 B.n314 B.n275 585
R393 B.n312 B.n311 585
R394 B.n310 B.n276 585
R395 B.n309 B.n308 585
R396 B.n306 B.n277 585
R397 B.n304 B.n303 585
R398 B.n302 B.n278 585
R399 B.n301 B.n300 585
R400 B.n298 B.n279 585
R401 B.n296 B.n295 585
R402 B.n294 B.n280 585
R403 B.n293 B.n292 585
R404 B.n290 B.n281 585
R405 B.n288 B.n287 585
R406 B.n286 B.n282 585
R407 B.n285 B.n284 585
R408 B.n228 B.n227 585
R409 B.n229 B.n228 585
R410 B.n474 B.n473 585
R411 B.n475 B.n474 585
R412 B.n224 B.n223 585
R413 B.n225 B.n224 585
R414 B.n483 B.n482 585
R415 B.n482 B.n481 585
R416 B.n484 B.n222 585
R417 B.n222 B.n221 585
R418 B.n486 B.n485 585
R419 B.n487 B.n486 585
R420 B.n216 B.n215 585
R421 B.n217 B.n216 585
R422 B.n495 B.n494 585
R423 B.n494 B.n493 585
R424 B.n496 B.n214 585
R425 B.n214 B.n212 585
R426 B.n498 B.n497 585
R427 B.n499 B.n498 585
R428 B.n208 B.n207 585
R429 B.n213 B.n208 585
R430 B.n507 B.n506 585
R431 B.n506 B.n505 585
R432 B.n508 B.n206 585
R433 B.n206 B.n205 585
R434 B.n510 B.n509 585
R435 B.n511 B.n510 585
R436 B.n200 B.n199 585
R437 B.n201 B.n200 585
R438 B.n519 B.n518 585
R439 B.n518 B.n517 585
R440 B.n520 B.n198 585
R441 B.n198 B.n197 585
R442 B.n522 B.n521 585
R443 B.n523 B.n522 585
R444 B.n192 B.n191 585
R445 B.n193 B.n192 585
R446 B.n531 B.n530 585
R447 B.n530 B.n529 585
R448 B.n532 B.n190 585
R449 B.n190 B.n189 585
R450 B.n534 B.n533 585
R451 B.n535 B.n534 585
R452 B.n184 B.n183 585
R453 B.n185 B.n184 585
R454 B.n543 B.n542 585
R455 B.n542 B.n541 585
R456 B.n544 B.n182 585
R457 B.n182 B.n180 585
R458 B.n546 B.n545 585
R459 B.n547 B.n546 585
R460 B.n176 B.n175 585
R461 B.n181 B.n176 585
R462 B.n555 B.n554 585
R463 B.n554 B.n553 585
R464 B.n556 B.n174 585
R465 B.n174 B.n173 585
R466 B.n558 B.n557 585
R467 B.n559 B.n558 585
R468 B.n168 B.n167 585
R469 B.n169 B.n168 585
R470 B.n567 B.n566 585
R471 B.n566 B.n565 585
R472 B.n568 B.n166 585
R473 B.n166 B.n165 585
R474 B.n570 B.n569 585
R475 B.n571 B.n570 585
R476 B.n160 B.n159 585
R477 B.n161 B.n160 585
R478 B.n579 B.n578 585
R479 B.n578 B.n577 585
R480 B.n580 B.n158 585
R481 B.n158 B.n157 585
R482 B.n582 B.n581 585
R483 B.n583 B.n582 585
R484 B.n152 B.n151 585
R485 B.n153 B.n152 585
R486 B.n591 B.n590 585
R487 B.n590 B.n589 585
R488 B.n592 B.n150 585
R489 B.n150 B.n149 585
R490 B.n594 B.n593 585
R491 B.n595 B.n594 585
R492 B.n144 B.n143 585
R493 B.n145 B.n144 585
R494 B.n604 B.n603 585
R495 B.n603 B.n602 585
R496 B.n605 B.n142 585
R497 B.n142 B.n141 585
R498 B.n607 B.n606 585
R499 B.n608 B.n607 585
R500 B.n2 B.n0 585
R501 B.n4 B.n2 585
R502 B.n3 B.n1 585
R503 B.n954 B.n3 585
R504 B.n952 B.n951 585
R505 B.n953 B.n952 585
R506 B.n950 B.n9 585
R507 B.n9 B.n8 585
R508 B.n949 B.n948 585
R509 B.n948 B.n947 585
R510 B.n11 B.n10 585
R511 B.n946 B.n11 585
R512 B.n944 B.n943 585
R513 B.n945 B.n944 585
R514 B.n942 B.n16 585
R515 B.n16 B.n15 585
R516 B.n941 B.n940 585
R517 B.n940 B.n939 585
R518 B.n18 B.n17 585
R519 B.n938 B.n18 585
R520 B.n936 B.n935 585
R521 B.n937 B.n936 585
R522 B.n934 B.n23 585
R523 B.n23 B.n22 585
R524 B.n933 B.n932 585
R525 B.n932 B.n931 585
R526 B.n25 B.n24 585
R527 B.n930 B.n25 585
R528 B.n928 B.n927 585
R529 B.n929 B.n928 585
R530 B.n926 B.n30 585
R531 B.n30 B.n29 585
R532 B.n925 B.n924 585
R533 B.n924 B.n923 585
R534 B.n32 B.n31 585
R535 B.n922 B.n32 585
R536 B.n920 B.n919 585
R537 B.n921 B.n920 585
R538 B.n918 B.n37 585
R539 B.n37 B.n36 585
R540 B.n917 B.n916 585
R541 B.n916 B.n915 585
R542 B.n39 B.n38 585
R543 B.n914 B.n39 585
R544 B.n912 B.n911 585
R545 B.n913 B.n912 585
R546 B.n910 B.n44 585
R547 B.n44 B.n43 585
R548 B.n909 B.n908 585
R549 B.n908 B.n907 585
R550 B.n46 B.n45 585
R551 B.n906 B.n46 585
R552 B.n904 B.n903 585
R553 B.n905 B.n904 585
R554 B.n902 B.n51 585
R555 B.n51 B.n50 585
R556 B.n901 B.n900 585
R557 B.n900 B.n899 585
R558 B.n53 B.n52 585
R559 B.n898 B.n53 585
R560 B.n896 B.n895 585
R561 B.n897 B.n896 585
R562 B.n894 B.n58 585
R563 B.n58 B.n57 585
R564 B.n893 B.n892 585
R565 B.n892 B.n891 585
R566 B.n60 B.n59 585
R567 B.n890 B.n60 585
R568 B.n888 B.n887 585
R569 B.n889 B.n888 585
R570 B.n886 B.n65 585
R571 B.n65 B.n64 585
R572 B.n885 B.n884 585
R573 B.n884 B.n883 585
R574 B.n67 B.n66 585
R575 B.n882 B.n67 585
R576 B.n880 B.n879 585
R577 B.n881 B.n880 585
R578 B.n878 B.n72 585
R579 B.n72 B.n71 585
R580 B.n877 B.n876 585
R581 B.n876 B.n875 585
R582 B.n74 B.n73 585
R583 B.n874 B.n74 585
R584 B.n872 B.n871 585
R585 B.n873 B.n872 585
R586 B.n870 B.n79 585
R587 B.n79 B.n78 585
R588 B.n869 B.n868 585
R589 B.n868 B.n867 585
R590 B.n81 B.n80 585
R591 B.n866 B.n81 585
R592 B.n864 B.n863 585
R593 B.n865 B.n864 585
R594 B.n957 B.n956 585
R595 B.n956 B.n955 585
R596 B.n474 B.n230 506.916
R597 B.n864 B.n86 506.916
R598 B.n476 B.n228 506.916
R599 B.n671 B.n84 506.916
R600 B.n259 B.t4 285.594
R601 B.n253 B.t15 285.594
R602 B.n109 B.t12 285.594
R603 B.n116 B.t8 285.594
R604 B.n672 B.n85 256.663
R605 B.n674 B.n85 256.663
R606 B.n680 B.n85 256.663
R607 B.n682 B.n85 256.663
R608 B.n688 B.n85 256.663
R609 B.n690 B.n85 256.663
R610 B.n696 B.n85 256.663
R611 B.n698 B.n85 256.663
R612 B.n704 B.n85 256.663
R613 B.n706 B.n85 256.663
R614 B.n712 B.n85 256.663
R615 B.n714 B.n85 256.663
R616 B.n720 B.n85 256.663
R617 B.n722 B.n85 256.663
R618 B.n728 B.n85 256.663
R619 B.n730 B.n85 256.663
R620 B.n736 B.n85 256.663
R621 B.n738 B.n85 256.663
R622 B.n744 B.n85 256.663
R623 B.n746 B.n85 256.663
R624 B.n752 B.n85 256.663
R625 B.n754 B.n85 256.663
R626 B.n761 B.n85 256.663
R627 B.n763 B.n85 256.663
R628 B.n769 B.n85 256.663
R629 B.n771 B.n85 256.663
R630 B.n777 B.n85 256.663
R631 B.n779 B.n85 256.663
R632 B.n785 B.n85 256.663
R633 B.n787 B.n85 256.663
R634 B.n793 B.n85 256.663
R635 B.n795 B.n85 256.663
R636 B.n801 B.n85 256.663
R637 B.n803 B.n85 256.663
R638 B.n809 B.n85 256.663
R639 B.n811 B.n85 256.663
R640 B.n817 B.n85 256.663
R641 B.n819 B.n85 256.663
R642 B.n825 B.n85 256.663
R643 B.n827 B.n85 256.663
R644 B.n833 B.n85 256.663
R645 B.n835 B.n85 256.663
R646 B.n841 B.n85 256.663
R647 B.n843 B.n85 256.663
R648 B.n849 B.n85 256.663
R649 B.n851 B.n85 256.663
R650 B.n857 B.n85 256.663
R651 B.n859 B.n85 256.663
R652 B.n469 B.n229 256.663
R653 B.n232 B.n229 256.663
R654 B.n462 B.n229 256.663
R655 B.n456 B.n229 256.663
R656 B.n454 B.n229 256.663
R657 B.n448 B.n229 256.663
R658 B.n446 B.n229 256.663
R659 B.n440 B.n229 256.663
R660 B.n438 B.n229 256.663
R661 B.n432 B.n229 256.663
R662 B.n430 B.n229 256.663
R663 B.n424 B.n229 256.663
R664 B.n422 B.n229 256.663
R665 B.n416 B.n229 256.663
R666 B.n414 B.n229 256.663
R667 B.n408 B.n229 256.663
R668 B.n406 B.n229 256.663
R669 B.n400 B.n229 256.663
R670 B.n398 B.n229 256.663
R671 B.n392 B.n229 256.663
R672 B.n390 B.n229 256.663
R673 B.n383 B.n229 256.663
R674 B.n381 B.n229 256.663
R675 B.n375 B.n229 256.663
R676 B.n373 B.n229 256.663
R677 B.n367 B.n229 256.663
R678 B.n262 B.n229 256.663
R679 B.n361 B.n229 256.663
R680 B.n355 B.n229 256.663
R681 B.n353 B.n229 256.663
R682 B.n347 B.n229 256.663
R683 B.n345 B.n229 256.663
R684 B.n339 B.n229 256.663
R685 B.n337 B.n229 256.663
R686 B.n331 B.n229 256.663
R687 B.n329 B.n229 256.663
R688 B.n323 B.n229 256.663
R689 B.n321 B.n229 256.663
R690 B.n315 B.n229 256.663
R691 B.n313 B.n229 256.663
R692 B.n307 B.n229 256.663
R693 B.n305 B.n229 256.663
R694 B.n299 B.n229 256.663
R695 B.n297 B.n229 256.663
R696 B.n291 B.n229 256.663
R697 B.n289 B.n229 256.663
R698 B.n283 B.n229 256.663
R699 B.n474 B.n224 163.367
R700 B.n482 B.n224 163.367
R701 B.n482 B.n222 163.367
R702 B.n486 B.n222 163.367
R703 B.n486 B.n216 163.367
R704 B.n494 B.n216 163.367
R705 B.n494 B.n214 163.367
R706 B.n498 B.n214 163.367
R707 B.n498 B.n208 163.367
R708 B.n506 B.n208 163.367
R709 B.n506 B.n206 163.367
R710 B.n510 B.n206 163.367
R711 B.n510 B.n200 163.367
R712 B.n518 B.n200 163.367
R713 B.n518 B.n198 163.367
R714 B.n522 B.n198 163.367
R715 B.n522 B.n192 163.367
R716 B.n530 B.n192 163.367
R717 B.n530 B.n190 163.367
R718 B.n534 B.n190 163.367
R719 B.n534 B.n184 163.367
R720 B.n542 B.n184 163.367
R721 B.n542 B.n182 163.367
R722 B.n546 B.n182 163.367
R723 B.n546 B.n176 163.367
R724 B.n554 B.n176 163.367
R725 B.n554 B.n174 163.367
R726 B.n558 B.n174 163.367
R727 B.n558 B.n168 163.367
R728 B.n566 B.n168 163.367
R729 B.n566 B.n166 163.367
R730 B.n570 B.n166 163.367
R731 B.n570 B.n160 163.367
R732 B.n578 B.n160 163.367
R733 B.n578 B.n158 163.367
R734 B.n582 B.n158 163.367
R735 B.n582 B.n152 163.367
R736 B.n590 B.n152 163.367
R737 B.n590 B.n150 163.367
R738 B.n594 B.n150 163.367
R739 B.n594 B.n144 163.367
R740 B.n603 B.n144 163.367
R741 B.n603 B.n142 163.367
R742 B.n607 B.n142 163.367
R743 B.n607 B.n2 163.367
R744 B.n956 B.n2 163.367
R745 B.n956 B.n3 163.367
R746 B.n952 B.n3 163.367
R747 B.n952 B.n9 163.367
R748 B.n948 B.n9 163.367
R749 B.n948 B.n11 163.367
R750 B.n944 B.n11 163.367
R751 B.n944 B.n16 163.367
R752 B.n940 B.n16 163.367
R753 B.n940 B.n18 163.367
R754 B.n936 B.n18 163.367
R755 B.n936 B.n23 163.367
R756 B.n932 B.n23 163.367
R757 B.n932 B.n25 163.367
R758 B.n928 B.n25 163.367
R759 B.n928 B.n30 163.367
R760 B.n924 B.n30 163.367
R761 B.n924 B.n32 163.367
R762 B.n920 B.n32 163.367
R763 B.n920 B.n37 163.367
R764 B.n916 B.n37 163.367
R765 B.n916 B.n39 163.367
R766 B.n912 B.n39 163.367
R767 B.n912 B.n44 163.367
R768 B.n908 B.n44 163.367
R769 B.n908 B.n46 163.367
R770 B.n904 B.n46 163.367
R771 B.n904 B.n51 163.367
R772 B.n900 B.n51 163.367
R773 B.n900 B.n53 163.367
R774 B.n896 B.n53 163.367
R775 B.n896 B.n58 163.367
R776 B.n892 B.n58 163.367
R777 B.n892 B.n60 163.367
R778 B.n888 B.n60 163.367
R779 B.n888 B.n65 163.367
R780 B.n884 B.n65 163.367
R781 B.n884 B.n67 163.367
R782 B.n880 B.n67 163.367
R783 B.n880 B.n72 163.367
R784 B.n876 B.n72 163.367
R785 B.n876 B.n74 163.367
R786 B.n872 B.n74 163.367
R787 B.n872 B.n79 163.367
R788 B.n868 B.n79 163.367
R789 B.n868 B.n81 163.367
R790 B.n864 B.n81 163.367
R791 B.n470 B.n468 163.367
R792 B.n468 B.n467 163.367
R793 B.n464 B.n463 163.367
R794 B.n461 B.n234 163.367
R795 B.n457 B.n455 163.367
R796 B.n453 B.n236 163.367
R797 B.n449 B.n447 163.367
R798 B.n445 B.n238 163.367
R799 B.n441 B.n439 163.367
R800 B.n437 B.n240 163.367
R801 B.n433 B.n431 163.367
R802 B.n429 B.n242 163.367
R803 B.n425 B.n423 163.367
R804 B.n421 B.n244 163.367
R805 B.n417 B.n415 163.367
R806 B.n413 B.n246 163.367
R807 B.n409 B.n407 163.367
R808 B.n405 B.n248 163.367
R809 B.n401 B.n399 163.367
R810 B.n397 B.n250 163.367
R811 B.n393 B.n391 163.367
R812 B.n389 B.n252 163.367
R813 B.n384 B.n382 163.367
R814 B.n380 B.n256 163.367
R815 B.n376 B.n374 163.367
R816 B.n372 B.n258 163.367
R817 B.n368 B.n366 163.367
R818 B.n363 B.n362 163.367
R819 B.n360 B.n264 163.367
R820 B.n356 B.n354 163.367
R821 B.n352 B.n266 163.367
R822 B.n348 B.n346 163.367
R823 B.n344 B.n268 163.367
R824 B.n340 B.n338 163.367
R825 B.n336 B.n270 163.367
R826 B.n332 B.n330 163.367
R827 B.n328 B.n272 163.367
R828 B.n324 B.n322 163.367
R829 B.n320 B.n274 163.367
R830 B.n316 B.n314 163.367
R831 B.n312 B.n276 163.367
R832 B.n308 B.n306 163.367
R833 B.n304 B.n278 163.367
R834 B.n300 B.n298 163.367
R835 B.n296 B.n280 163.367
R836 B.n292 B.n290 163.367
R837 B.n288 B.n282 163.367
R838 B.n284 B.n228 163.367
R839 B.n476 B.n226 163.367
R840 B.n480 B.n226 163.367
R841 B.n480 B.n220 163.367
R842 B.n488 B.n220 163.367
R843 B.n488 B.n218 163.367
R844 B.n492 B.n218 163.367
R845 B.n492 B.n211 163.367
R846 B.n500 B.n211 163.367
R847 B.n500 B.n209 163.367
R848 B.n504 B.n209 163.367
R849 B.n504 B.n204 163.367
R850 B.n512 B.n204 163.367
R851 B.n512 B.n202 163.367
R852 B.n516 B.n202 163.367
R853 B.n516 B.n196 163.367
R854 B.n524 B.n196 163.367
R855 B.n524 B.n194 163.367
R856 B.n528 B.n194 163.367
R857 B.n528 B.n188 163.367
R858 B.n536 B.n188 163.367
R859 B.n536 B.n186 163.367
R860 B.n540 B.n186 163.367
R861 B.n540 B.n179 163.367
R862 B.n548 B.n179 163.367
R863 B.n548 B.n177 163.367
R864 B.n552 B.n177 163.367
R865 B.n552 B.n172 163.367
R866 B.n560 B.n172 163.367
R867 B.n560 B.n170 163.367
R868 B.n564 B.n170 163.367
R869 B.n564 B.n164 163.367
R870 B.n572 B.n164 163.367
R871 B.n572 B.n162 163.367
R872 B.n576 B.n162 163.367
R873 B.n576 B.n156 163.367
R874 B.n584 B.n156 163.367
R875 B.n584 B.n154 163.367
R876 B.n588 B.n154 163.367
R877 B.n588 B.n148 163.367
R878 B.n596 B.n148 163.367
R879 B.n596 B.n146 163.367
R880 B.n601 B.n146 163.367
R881 B.n601 B.n140 163.367
R882 B.n609 B.n140 163.367
R883 B.n610 B.n609 163.367
R884 B.n610 B.n5 163.367
R885 B.n6 B.n5 163.367
R886 B.n7 B.n6 163.367
R887 B.n615 B.n7 163.367
R888 B.n615 B.n12 163.367
R889 B.n13 B.n12 163.367
R890 B.n14 B.n13 163.367
R891 B.n620 B.n14 163.367
R892 B.n620 B.n19 163.367
R893 B.n20 B.n19 163.367
R894 B.n21 B.n20 163.367
R895 B.n625 B.n21 163.367
R896 B.n625 B.n26 163.367
R897 B.n27 B.n26 163.367
R898 B.n28 B.n27 163.367
R899 B.n630 B.n28 163.367
R900 B.n630 B.n33 163.367
R901 B.n34 B.n33 163.367
R902 B.n35 B.n34 163.367
R903 B.n635 B.n35 163.367
R904 B.n635 B.n40 163.367
R905 B.n41 B.n40 163.367
R906 B.n42 B.n41 163.367
R907 B.n640 B.n42 163.367
R908 B.n640 B.n47 163.367
R909 B.n48 B.n47 163.367
R910 B.n49 B.n48 163.367
R911 B.n645 B.n49 163.367
R912 B.n645 B.n54 163.367
R913 B.n55 B.n54 163.367
R914 B.n56 B.n55 163.367
R915 B.n650 B.n56 163.367
R916 B.n650 B.n61 163.367
R917 B.n62 B.n61 163.367
R918 B.n63 B.n62 163.367
R919 B.n655 B.n63 163.367
R920 B.n655 B.n68 163.367
R921 B.n69 B.n68 163.367
R922 B.n70 B.n69 163.367
R923 B.n660 B.n70 163.367
R924 B.n660 B.n75 163.367
R925 B.n76 B.n75 163.367
R926 B.n77 B.n76 163.367
R927 B.n665 B.n77 163.367
R928 B.n665 B.n82 163.367
R929 B.n83 B.n82 163.367
R930 B.n84 B.n83 163.367
R931 B.n860 B.n858 163.367
R932 B.n856 B.n88 163.367
R933 B.n852 B.n850 163.367
R934 B.n848 B.n90 163.367
R935 B.n844 B.n842 163.367
R936 B.n840 B.n92 163.367
R937 B.n836 B.n834 163.367
R938 B.n832 B.n94 163.367
R939 B.n828 B.n826 163.367
R940 B.n824 B.n96 163.367
R941 B.n820 B.n818 163.367
R942 B.n816 B.n98 163.367
R943 B.n812 B.n810 163.367
R944 B.n808 B.n100 163.367
R945 B.n804 B.n802 163.367
R946 B.n800 B.n102 163.367
R947 B.n796 B.n794 163.367
R948 B.n792 B.n104 163.367
R949 B.n788 B.n786 163.367
R950 B.n784 B.n106 163.367
R951 B.n780 B.n778 163.367
R952 B.n776 B.n108 163.367
R953 B.n772 B.n770 163.367
R954 B.n768 B.n113 163.367
R955 B.n764 B.n762 163.367
R956 B.n760 B.n115 163.367
R957 B.n755 B.n753 163.367
R958 B.n751 B.n119 163.367
R959 B.n747 B.n745 163.367
R960 B.n743 B.n121 163.367
R961 B.n739 B.n737 163.367
R962 B.n735 B.n123 163.367
R963 B.n731 B.n729 163.367
R964 B.n727 B.n125 163.367
R965 B.n723 B.n721 163.367
R966 B.n719 B.n127 163.367
R967 B.n715 B.n713 163.367
R968 B.n711 B.n129 163.367
R969 B.n707 B.n705 163.367
R970 B.n703 B.n131 163.367
R971 B.n699 B.n697 163.367
R972 B.n695 B.n133 163.367
R973 B.n691 B.n689 163.367
R974 B.n687 B.n135 163.367
R975 B.n683 B.n681 163.367
R976 B.n679 B.n137 163.367
R977 B.n675 B.n673 163.367
R978 B.n259 B.t7 156.931
R979 B.n116 B.t10 156.931
R980 B.n253 B.t17 156.916
R981 B.n109 B.t13 156.916
R982 B.n260 B.n259 83.3944
R983 B.n254 B.n253 83.3944
R984 B.n110 B.n109 83.3944
R985 B.n117 B.n116 83.3944
R986 B.n475 B.n229 78.4176
R987 B.n865 B.n85 78.4176
R988 B.n260 B.t6 73.5375
R989 B.n117 B.t11 73.5375
R990 B.n254 B.t16 73.5218
R991 B.n110 B.t14 73.5218
R992 B.n469 B.n230 71.676
R993 B.n467 B.n232 71.676
R994 B.n463 B.n462 71.676
R995 B.n456 B.n234 71.676
R996 B.n455 B.n454 71.676
R997 B.n448 B.n236 71.676
R998 B.n447 B.n446 71.676
R999 B.n440 B.n238 71.676
R1000 B.n439 B.n438 71.676
R1001 B.n432 B.n240 71.676
R1002 B.n431 B.n430 71.676
R1003 B.n424 B.n242 71.676
R1004 B.n423 B.n422 71.676
R1005 B.n416 B.n244 71.676
R1006 B.n415 B.n414 71.676
R1007 B.n408 B.n246 71.676
R1008 B.n407 B.n406 71.676
R1009 B.n400 B.n248 71.676
R1010 B.n399 B.n398 71.676
R1011 B.n392 B.n250 71.676
R1012 B.n391 B.n390 71.676
R1013 B.n383 B.n252 71.676
R1014 B.n382 B.n381 71.676
R1015 B.n375 B.n256 71.676
R1016 B.n374 B.n373 71.676
R1017 B.n367 B.n258 71.676
R1018 B.n366 B.n262 71.676
R1019 B.n362 B.n361 71.676
R1020 B.n355 B.n264 71.676
R1021 B.n354 B.n353 71.676
R1022 B.n347 B.n266 71.676
R1023 B.n346 B.n345 71.676
R1024 B.n339 B.n268 71.676
R1025 B.n338 B.n337 71.676
R1026 B.n331 B.n270 71.676
R1027 B.n330 B.n329 71.676
R1028 B.n323 B.n272 71.676
R1029 B.n322 B.n321 71.676
R1030 B.n315 B.n274 71.676
R1031 B.n314 B.n313 71.676
R1032 B.n307 B.n276 71.676
R1033 B.n306 B.n305 71.676
R1034 B.n299 B.n278 71.676
R1035 B.n298 B.n297 71.676
R1036 B.n291 B.n280 71.676
R1037 B.n290 B.n289 71.676
R1038 B.n283 B.n282 71.676
R1039 B.n859 B.n86 71.676
R1040 B.n858 B.n857 71.676
R1041 B.n851 B.n88 71.676
R1042 B.n850 B.n849 71.676
R1043 B.n843 B.n90 71.676
R1044 B.n842 B.n841 71.676
R1045 B.n835 B.n92 71.676
R1046 B.n834 B.n833 71.676
R1047 B.n827 B.n94 71.676
R1048 B.n826 B.n825 71.676
R1049 B.n819 B.n96 71.676
R1050 B.n818 B.n817 71.676
R1051 B.n811 B.n98 71.676
R1052 B.n810 B.n809 71.676
R1053 B.n803 B.n100 71.676
R1054 B.n802 B.n801 71.676
R1055 B.n795 B.n102 71.676
R1056 B.n794 B.n793 71.676
R1057 B.n787 B.n104 71.676
R1058 B.n786 B.n785 71.676
R1059 B.n779 B.n106 71.676
R1060 B.n778 B.n777 71.676
R1061 B.n771 B.n108 71.676
R1062 B.n770 B.n769 71.676
R1063 B.n763 B.n113 71.676
R1064 B.n762 B.n761 71.676
R1065 B.n754 B.n115 71.676
R1066 B.n753 B.n752 71.676
R1067 B.n746 B.n119 71.676
R1068 B.n745 B.n744 71.676
R1069 B.n738 B.n121 71.676
R1070 B.n737 B.n736 71.676
R1071 B.n730 B.n123 71.676
R1072 B.n729 B.n728 71.676
R1073 B.n722 B.n125 71.676
R1074 B.n721 B.n720 71.676
R1075 B.n714 B.n127 71.676
R1076 B.n713 B.n712 71.676
R1077 B.n706 B.n129 71.676
R1078 B.n705 B.n704 71.676
R1079 B.n698 B.n131 71.676
R1080 B.n697 B.n696 71.676
R1081 B.n690 B.n133 71.676
R1082 B.n689 B.n688 71.676
R1083 B.n682 B.n135 71.676
R1084 B.n681 B.n680 71.676
R1085 B.n674 B.n137 71.676
R1086 B.n673 B.n672 71.676
R1087 B.n672 B.n671 71.676
R1088 B.n675 B.n674 71.676
R1089 B.n680 B.n679 71.676
R1090 B.n683 B.n682 71.676
R1091 B.n688 B.n687 71.676
R1092 B.n691 B.n690 71.676
R1093 B.n696 B.n695 71.676
R1094 B.n699 B.n698 71.676
R1095 B.n704 B.n703 71.676
R1096 B.n707 B.n706 71.676
R1097 B.n712 B.n711 71.676
R1098 B.n715 B.n714 71.676
R1099 B.n720 B.n719 71.676
R1100 B.n723 B.n722 71.676
R1101 B.n728 B.n727 71.676
R1102 B.n731 B.n730 71.676
R1103 B.n736 B.n735 71.676
R1104 B.n739 B.n738 71.676
R1105 B.n744 B.n743 71.676
R1106 B.n747 B.n746 71.676
R1107 B.n752 B.n751 71.676
R1108 B.n755 B.n754 71.676
R1109 B.n761 B.n760 71.676
R1110 B.n764 B.n763 71.676
R1111 B.n769 B.n768 71.676
R1112 B.n772 B.n771 71.676
R1113 B.n777 B.n776 71.676
R1114 B.n780 B.n779 71.676
R1115 B.n785 B.n784 71.676
R1116 B.n788 B.n787 71.676
R1117 B.n793 B.n792 71.676
R1118 B.n796 B.n795 71.676
R1119 B.n801 B.n800 71.676
R1120 B.n804 B.n803 71.676
R1121 B.n809 B.n808 71.676
R1122 B.n812 B.n811 71.676
R1123 B.n817 B.n816 71.676
R1124 B.n820 B.n819 71.676
R1125 B.n825 B.n824 71.676
R1126 B.n828 B.n827 71.676
R1127 B.n833 B.n832 71.676
R1128 B.n836 B.n835 71.676
R1129 B.n841 B.n840 71.676
R1130 B.n844 B.n843 71.676
R1131 B.n849 B.n848 71.676
R1132 B.n852 B.n851 71.676
R1133 B.n857 B.n856 71.676
R1134 B.n860 B.n859 71.676
R1135 B.n470 B.n469 71.676
R1136 B.n464 B.n232 71.676
R1137 B.n462 B.n461 71.676
R1138 B.n457 B.n456 71.676
R1139 B.n454 B.n453 71.676
R1140 B.n449 B.n448 71.676
R1141 B.n446 B.n445 71.676
R1142 B.n441 B.n440 71.676
R1143 B.n438 B.n437 71.676
R1144 B.n433 B.n432 71.676
R1145 B.n430 B.n429 71.676
R1146 B.n425 B.n424 71.676
R1147 B.n422 B.n421 71.676
R1148 B.n417 B.n416 71.676
R1149 B.n414 B.n413 71.676
R1150 B.n409 B.n408 71.676
R1151 B.n406 B.n405 71.676
R1152 B.n401 B.n400 71.676
R1153 B.n398 B.n397 71.676
R1154 B.n393 B.n392 71.676
R1155 B.n390 B.n389 71.676
R1156 B.n384 B.n383 71.676
R1157 B.n381 B.n380 71.676
R1158 B.n376 B.n375 71.676
R1159 B.n373 B.n372 71.676
R1160 B.n368 B.n367 71.676
R1161 B.n363 B.n262 71.676
R1162 B.n361 B.n360 71.676
R1163 B.n356 B.n355 71.676
R1164 B.n353 B.n352 71.676
R1165 B.n348 B.n347 71.676
R1166 B.n345 B.n344 71.676
R1167 B.n340 B.n339 71.676
R1168 B.n337 B.n336 71.676
R1169 B.n332 B.n331 71.676
R1170 B.n329 B.n328 71.676
R1171 B.n324 B.n323 71.676
R1172 B.n321 B.n320 71.676
R1173 B.n316 B.n315 71.676
R1174 B.n313 B.n312 71.676
R1175 B.n308 B.n307 71.676
R1176 B.n305 B.n304 71.676
R1177 B.n300 B.n299 71.676
R1178 B.n297 B.n296 71.676
R1179 B.n292 B.n291 71.676
R1180 B.n289 B.n288 71.676
R1181 B.n284 B.n283 71.676
R1182 B.n261 B.n260 59.5399
R1183 B.n387 B.n254 59.5399
R1184 B.n111 B.n110 59.5399
R1185 B.n757 B.n117 59.5399
R1186 B.n475 B.n225 41.9876
R1187 B.n481 B.n225 41.9876
R1188 B.n481 B.n221 41.9876
R1189 B.n487 B.n221 41.9876
R1190 B.n487 B.n217 41.9876
R1191 B.n493 B.n217 41.9876
R1192 B.n493 B.n212 41.9876
R1193 B.n499 B.n212 41.9876
R1194 B.n499 B.n213 41.9876
R1195 B.n505 B.n205 41.9876
R1196 B.n511 B.n205 41.9876
R1197 B.n511 B.n201 41.9876
R1198 B.n517 B.n201 41.9876
R1199 B.n517 B.n197 41.9876
R1200 B.n523 B.n197 41.9876
R1201 B.n523 B.n193 41.9876
R1202 B.n529 B.n193 41.9876
R1203 B.n529 B.n189 41.9876
R1204 B.n535 B.n189 41.9876
R1205 B.n535 B.n185 41.9876
R1206 B.n541 B.n185 41.9876
R1207 B.n541 B.n180 41.9876
R1208 B.n547 B.n180 41.9876
R1209 B.n547 B.n181 41.9876
R1210 B.n553 B.n173 41.9876
R1211 B.n559 B.n173 41.9876
R1212 B.n559 B.n169 41.9876
R1213 B.n565 B.n169 41.9876
R1214 B.n565 B.n165 41.9876
R1215 B.n571 B.n165 41.9876
R1216 B.n571 B.n161 41.9876
R1217 B.n577 B.n161 41.9876
R1218 B.n577 B.n157 41.9876
R1219 B.n583 B.n157 41.9876
R1220 B.n583 B.n153 41.9876
R1221 B.n589 B.n153 41.9876
R1222 B.n595 B.n149 41.9876
R1223 B.n595 B.n145 41.9876
R1224 B.n602 B.n145 41.9876
R1225 B.n602 B.n141 41.9876
R1226 B.n608 B.n141 41.9876
R1227 B.n608 B.n4 41.9876
R1228 B.n955 B.n4 41.9876
R1229 B.n955 B.n954 41.9876
R1230 B.n954 B.n953 41.9876
R1231 B.n953 B.n8 41.9876
R1232 B.n947 B.n8 41.9876
R1233 B.n947 B.n946 41.9876
R1234 B.n946 B.n945 41.9876
R1235 B.n945 B.n15 41.9876
R1236 B.n939 B.n938 41.9876
R1237 B.n938 B.n937 41.9876
R1238 B.n937 B.n22 41.9876
R1239 B.n931 B.n22 41.9876
R1240 B.n931 B.n930 41.9876
R1241 B.n930 B.n929 41.9876
R1242 B.n929 B.n29 41.9876
R1243 B.n923 B.n29 41.9876
R1244 B.n923 B.n922 41.9876
R1245 B.n922 B.n921 41.9876
R1246 B.n921 B.n36 41.9876
R1247 B.n915 B.n36 41.9876
R1248 B.n914 B.n913 41.9876
R1249 B.n913 B.n43 41.9876
R1250 B.n907 B.n43 41.9876
R1251 B.n907 B.n906 41.9876
R1252 B.n906 B.n905 41.9876
R1253 B.n905 B.n50 41.9876
R1254 B.n899 B.n50 41.9876
R1255 B.n899 B.n898 41.9876
R1256 B.n898 B.n897 41.9876
R1257 B.n897 B.n57 41.9876
R1258 B.n891 B.n57 41.9876
R1259 B.n891 B.n890 41.9876
R1260 B.n890 B.n889 41.9876
R1261 B.n889 B.n64 41.9876
R1262 B.n883 B.n64 41.9876
R1263 B.n882 B.n881 41.9876
R1264 B.n881 B.n71 41.9876
R1265 B.n875 B.n71 41.9876
R1266 B.n875 B.n874 41.9876
R1267 B.n874 B.n873 41.9876
R1268 B.n873 B.n78 41.9876
R1269 B.n867 B.n78 41.9876
R1270 B.n867 B.n866 41.9876
R1271 B.n866 B.n865 41.9876
R1272 B.t0 B.n149 38.9003
R1273 B.t1 B.n15 38.9003
R1274 B.n863 B.n862 32.9371
R1275 B.n670 B.n669 32.9371
R1276 B.n477 B.n227 32.9371
R1277 B.n473 B.n472 32.9371
R1278 B.n213 B.t5 24.0813
R1279 B.n553 B.t2 24.0813
R1280 B.n915 B.t3 24.0813
R1281 B.t9 B.n882 24.0813
R1282 B B.n957 18.0485
R1283 B.n505 B.t5 17.9068
R1284 B.n181 B.t2 17.9068
R1285 B.t3 B.n914 17.9068
R1286 B.n883 B.t9 17.9068
R1287 B.n862 B.n861 10.6151
R1288 B.n861 B.n87 10.6151
R1289 B.n855 B.n87 10.6151
R1290 B.n855 B.n854 10.6151
R1291 B.n854 B.n853 10.6151
R1292 B.n853 B.n89 10.6151
R1293 B.n847 B.n89 10.6151
R1294 B.n847 B.n846 10.6151
R1295 B.n846 B.n845 10.6151
R1296 B.n845 B.n91 10.6151
R1297 B.n839 B.n91 10.6151
R1298 B.n839 B.n838 10.6151
R1299 B.n838 B.n837 10.6151
R1300 B.n837 B.n93 10.6151
R1301 B.n831 B.n93 10.6151
R1302 B.n831 B.n830 10.6151
R1303 B.n830 B.n829 10.6151
R1304 B.n829 B.n95 10.6151
R1305 B.n823 B.n95 10.6151
R1306 B.n823 B.n822 10.6151
R1307 B.n822 B.n821 10.6151
R1308 B.n821 B.n97 10.6151
R1309 B.n815 B.n97 10.6151
R1310 B.n815 B.n814 10.6151
R1311 B.n814 B.n813 10.6151
R1312 B.n813 B.n99 10.6151
R1313 B.n807 B.n99 10.6151
R1314 B.n807 B.n806 10.6151
R1315 B.n806 B.n805 10.6151
R1316 B.n805 B.n101 10.6151
R1317 B.n799 B.n101 10.6151
R1318 B.n799 B.n798 10.6151
R1319 B.n798 B.n797 10.6151
R1320 B.n797 B.n103 10.6151
R1321 B.n791 B.n103 10.6151
R1322 B.n791 B.n790 10.6151
R1323 B.n790 B.n789 10.6151
R1324 B.n789 B.n105 10.6151
R1325 B.n783 B.n105 10.6151
R1326 B.n783 B.n782 10.6151
R1327 B.n782 B.n781 10.6151
R1328 B.n781 B.n107 10.6151
R1329 B.n775 B.n774 10.6151
R1330 B.n774 B.n773 10.6151
R1331 B.n773 B.n112 10.6151
R1332 B.n767 B.n112 10.6151
R1333 B.n767 B.n766 10.6151
R1334 B.n766 B.n765 10.6151
R1335 B.n765 B.n114 10.6151
R1336 B.n759 B.n114 10.6151
R1337 B.n759 B.n758 10.6151
R1338 B.n756 B.n118 10.6151
R1339 B.n750 B.n118 10.6151
R1340 B.n750 B.n749 10.6151
R1341 B.n749 B.n748 10.6151
R1342 B.n748 B.n120 10.6151
R1343 B.n742 B.n120 10.6151
R1344 B.n742 B.n741 10.6151
R1345 B.n741 B.n740 10.6151
R1346 B.n740 B.n122 10.6151
R1347 B.n734 B.n122 10.6151
R1348 B.n734 B.n733 10.6151
R1349 B.n733 B.n732 10.6151
R1350 B.n732 B.n124 10.6151
R1351 B.n726 B.n124 10.6151
R1352 B.n726 B.n725 10.6151
R1353 B.n725 B.n724 10.6151
R1354 B.n724 B.n126 10.6151
R1355 B.n718 B.n126 10.6151
R1356 B.n718 B.n717 10.6151
R1357 B.n717 B.n716 10.6151
R1358 B.n716 B.n128 10.6151
R1359 B.n710 B.n128 10.6151
R1360 B.n710 B.n709 10.6151
R1361 B.n709 B.n708 10.6151
R1362 B.n708 B.n130 10.6151
R1363 B.n702 B.n130 10.6151
R1364 B.n702 B.n701 10.6151
R1365 B.n701 B.n700 10.6151
R1366 B.n700 B.n132 10.6151
R1367 B.n694 B.n132 10.6151
R1368 B.n694 B.n693 10.6151
R1369 B.n693 B.n692 10.6151
R1370 B.n692 B.n134 10.6151
R1371 B.n686 B.n134 10.6151
R1372 B.n686 B.n685 10.6151
R1373 B.n685 B.n684 10.6151
R1374 B.n684 B.n136 10.6151
R1375 B.n678 B.n136 10.6151
R1376 B.n678 B.n677 10.6151
R1377 B.n677 B.n676 10.6151
R1378 B.n676 B.n138 10.6151
R1379 B.n670 B.n138 10.6151
R1380 B.n478 B.n477 10.6151
R1381 B.n479 B.n478 10.6151
R1382 B.n479 B.n219 10.6151
R1383 B.n489 B.n219 10.6151
R1384 B.n490 B.n489 10.6151
R1385 B.n491 B.n490 10.6151
R1386 B.n491 B.n210 10.6151
R1387 B.n501 B.n210 10.6151
R1388 B.n502 B.n501 10.6151
R1389 B.n503 B.n502 10.6151
R1390 B.n503 B.n203 10.6151
R1391 B.n513 B.n203 10.6151
R1392 B.n514 B.n513 10.6151
R1393 B.n515 B.n514 10.6151
R1394 B.n515 B.n195 10.6151
R1395 B.n525 B.n195 10.6151
R1396 B.n526 B.n525 10.6151
R1397 B.n527 B.n526 10.6151
R1398 B.n527 B.n187 10.6151
R1399 B.n537 B.n187 10.6151
R1400 B.n538 B.n537 10.6151
R1401 B.n539 B.n538 10.6151
R1402 B.n539 B.n178 10.6151
R1403 B.n549 B.n178 10.6151
R1404 B.n550 B.n549 10.6151
R1405 B.n551 B.n550 10.6151
R1406 B.n551 B.n171 10.6151
R1407 B.n561 B.n171 10.6151
R1408 B.n562 B.n561 10.6151
R1409 B.n563 B.n562 10.6151
R1410 B.n563 B.n163 10.6151
R1411 B.n573 B.n163 10.6151
R1412 B.n574 B.n573 10.6151
R1413 B.n575 B.n574 10.6151
R1414 B.n575 B.n155 10.6151
R1415 B.n585 B.n155 10.6151
R1416 B.n586 B.n585 10.6151
R1417 B.n587 B.n586 10.6151
R1418 B.n587 B.n147 10.6151
R1419 B.n597 B.n147 10.6151
R1420 B.n598 B.n597 10.6151
R1421 B.n600 B.n598 10.6151
R1422 B.n600 B.n599 10.6151
R1423 B.n599 B.n139 10.6151
R1424 B.n611 B.n139 10.6151
R1425 B.n612 B.n611 10.6151
R1426 B.n613 B.n612 10.6151
R1427 B.n614 B.n613 10.6151
R1428 B.n616 B.n614 10.6151
R1429 B.n617 B.n616 10.6151
R1430 B.n618 B.n617 10.6151
R1431 B.n619 B.n618 10.6151
R1432 B.n621 B.n619 10.6151
R1433 B.n622 B.n621 10.6151
R1434 B.n623 B.n622 10.6151
R1435 B.n624 B.n623 10.6151
R1436 B.n626 B.n624 10.6151
R1437 B.n627 B.n626 10.6151
R1438 B.n628 B.n627 10.6151
R1439 B.n629 B.n628 10.6151
R1440 B.n631 B.n629 10.6151
R1441 B.n632 B.n631 10.6151
R1442 B.n633 B.n632 10.6151
R1443 B.n634 B.n633 10.6151
R1444 B.n636 B.n634 10.6151
R1445 B.n637 B.n636 10.6151
R1446 B.n638 B.n637 10.6151
R1447 B.n639 B.n638 10.6151
R1448 B.n641 B.n639 10.6151
R1449 B.n642 B.n641 10.6151
R1450 B.n643 B.n642 10.6151
R1451 B.n644 B.n643 10.6151
R1452 B.n646 B.n644 10.6151
R1453 B.n647 B.n646 10.6151
R1454 B.n648 B.n647 10.6151
R1455 B.n649 B.n648 10.6151
R1456 B.n651 B.n649 10.6151
R1457 B.n652 B.n651 10.6151
R1458 B.n653 B.n652 10.6151
R1459 B.n654 B.n653 10.6151
R1460 B.n656 B.n654 10.6151
R1461 B.n657 B.n656 10.6151
R1462 B.n658 B.n657 10.6151
R1463 B.n659 B.n658 10.6151
R1464 B.n661 B.n659 10.6151
R1465 B.n662 B.n661 10.6151
R1466 B.n663 B.n662 10.6151
R1467 B.n664 B.n663 10.6151
R1468 B.n666 B.n664 10.6151
R1469 B.n667 B.n666 10.6151
R1470 B.n668 B.n667 10.6151
R1471 B.n669 B.n668 10.6151
R1472 B.n472 B.n471 10.6151
R1473 B.n471 B.n231 10.6151
R1474 B.n466 B.n231 10.6151
R1475 B.n466 B.n465 10.6151
R1476 B.n465 B.n233 10.6151
R1477 B.n460 B.n233 10.6151
R1478 B.n460 B.n459 10.6151
R1479 B.n459 B.n458 10.6151
R1480 B.n458 B.n235 10.6151
R1481 B.n452 B.n235 10.6151
R1482 B.n452 B.n451 10.6151
R1483 B.n451 B.n450 10.6151
R1484 B.n450 B.n237 10.6151
R1485 B.n444 B.n237 10.6151
R1486 B.n444 B.n443 10.6151
R1487 B.n443 B.n442 10.6151
R1488 B.n442 B.n239 10.6151
R1489 B.n436 B.n239 10.6151
R1490 B.n436 B.n435 10.6151
R1491 B.n435 B.n434 10.6151
R1492 B.n434 B.n241 10.6151
R1493 B.n428 B.n241 10.6151
R1494 B.n428 B.n427 10.6151
R1495 B.n427 B.n426 10.6151
R1496 B.n426 B.n243 10.6151
R1497 B.n420 B.n243 10.6151
R1498 B.n420 B.n419 10.6151
R1499 B.n419 B.n418 10.6151
R1500 B.n418 B.n245 10.6151
R1501 B.n412 B.n245 10.6151
R1502 B.n412 B.n411 10.6151
R1503 B.n411 B.n410 10.6151
R1504 B.n410 B.n247 10.6151
R1505 B.n404 B.n247 10.6151
R1506 B.n404 B.n403 10.6151
R1507 B.n403 B.n402 10.6151
R1508 B.n402 B.n249 10.6151
R1509 B.n396 B.n249 10.6151
R1510 B.n396 B.n395 10.6151
R1511 B.n395 B.n394 10.6151
R1512 B.n394 B.n251 10.6151
R1513 B.n388 B.n251 10.6151
R1514 B.n386 B.n385 10.6151
R1515 B.n385 B.n255 10.6151
R1516 B.n379 B.n255 10.6151
R1517 B.n379 B.n378 10.6151
R1518 B.n378 B.n377 10.6151
R1519 B.n377 B.n257 10.6151
R1520 B.n371 B.n257 10.6151
R1521 B.n371 B.n370 10.6151
R1522 B.n370 B.n369 10.6151
R1523 B.n365 B.n364 10.6151
R1524 B.n364 B.n263 10.6151
R1525 B.n359 B.n263 10.6151
R1526 B.n359 B.n358 10.6151
R1527 B.n358 B.n357 10.6151
R1528 B.n357 B.n265 10.6151
R1529 B.n351 B.n265 10.6151
R1530 B.n351 B.n350 10.6151
R1531 B.n350 B.n349 10.6151
R1532 B.n349 B.n267 10.6151
R1533 B.n343 B.n267 10.6151
R1534 B.n343 B.n342 10.6151
R1535 B.n342 B.n341 10.6151
R1536 B.n341 B.n269 10.6151
R1537 B.n335 B.n269 10.6151
R1538 B.n335 B.n334 10.6151
R1539 B.n334 B.n333 10.6151
R1540 B.n333 B.n271 10.6151
R1541 B.n327 B.n271 10.6151
R1542 B.n327 B.n326 10.6151
R1543 B.n326 B.n325 10.6151
R1544 B.n325 B.n273 10.6151
R1545 B.n319 B.n273 10.6151
R1546 B.n319 B.n318 10.6151
R1547 B.n318 B.n317 10.6151
R1548 B.n317 B.n275 10.6151
R1549 B.n311 B.n275 10.6151
R1550 B.n311 B.n310 10.6151
R1551 B.n310 B.n309 10.6151
R1552 B.n309 B.n277 10.6151
R1553 B.n303 B.n277 10.6151
R1554 B.n303 B.n302 10.6151
R1555 B.n302 B.n301 10.6151
R1556 B.n301 B.n279 10.6151
R1557 B.n295 B.n279 10.6151
R1558 B.n295 B.n294 10.6151
R1559 B.n294 B.n293 10.6151
R1560 B.n293 B.n281 10.6151
R1561 B.n287 B.n281 10.6151
R1562 B.n287 B.n286 10.6151
R1563 B.n286 B.n285 10.6151
R1564 B.n285 B.n227 10.6151
R1565 B.n473 B.n223 10.6151
R1566 B.n483 B.n223 10.6151
R1567 B.n484 B.n483 10.6151
R1568 B.n485 B.n484 10.6151
R1569 B.n485 B.n215 10.6151
R1570 B.n495 B.n215 10.6151
R1571 B.n496 B.n495 10.6151
R1572 B.n497 B.n496 10.6151
R1573 B.n497 B.n207 10.6151
R1574 B.n507 B.n207 10.6151
R1575 B.n508 B.n507 10.6151
R1576 B.n509 B.n508 10.6151
R1577 B.n509 B.n199 10.6151
R1578 B.n519 B.n199 10.6151
R1579 B.n520 B.n519 10.6151
R1580 B.n521 B.n520 10.6151
R1581 B.n521 B.n191 10.6151
R1582 B.n531 B.n191 10.6151
R1583 B.n532 B.n531 10.6151
R1584 B.n533 B.n532 10.6151
R1585 B.n533 B.n183 10.6151
R1586 B.n543 B.n183 10.6151
R1587 B.n544 B.n543 10.6151
R1588 B.n545 B.n544 10.6151
R1589 B.n545 B.n175 10.6151
R1590 B.n555 B.n175 10.6151
R1591 B.n556 B.n555 10.6151
R1592 B.n557 B.n556 10.6151
R1593 B.n557 B.n167 10.6151
R1594 B.n567 B.n167 10.6151
R1595 B.n568 B.n567 10.6151
R1596 B.n569 B.n568 10.6151
R1597 B.n569 B.n159 10.6151
R1598 B.n579 B.n159 10.6151
R1599 B.n580 B.n579 10.6151
R1600 B.n581 B.n580 10.6151
R1601 B.n581 B.n151 10.6151
R1602 B.n591 B.n151 10.6151
R1603 B.n592 B.n591 10.6151
R1604 B.n593 B.n592 10.6151
R1605 B.n593 B.n143 10.6151
R1606 B.n604 B.n143 10.6151
R1607 B.n605 B.n604 10.6151
R1608 B.n606 B.n605 10.6151
R1609 B.n606 B.n0 10.6151
R1610 B.n951 B.n1 10.6151
R1611 B.n951 B.n950 10.6151
R1612 B.n950 B.n949 10.6151
R1613 B.n949 B.n10 10.6151
R1614 B.n943 B.n10 10.6151
R1615 B.n943 B.n942 10.6151
R1616 B.n942 B.n941 10.6151
R1617 B.n941 B.n17 10.6151
R1618 B.n935 B.n17 10.6151
R1619 B.n935 B.n934 10.6151
R1620 B.n934 B.n933 10.6151
R1621 B.n933 B.n24 10.6151
R1622 B.n927 B.n24 10.6151
R1623 B.n927 B.n926 10.6151
R1624 B.n926 B.n925 10.6151
R1625 B.n925 B.n31 10.6151
R1626 B.n919 B.n31 10.6151
R1627 B.n919 B.n918 10.6151
R1628 B.n918 B.n917 10.6151
R1629 B.n917 B.n38 10.6151
R1630 B.n911 B.n38 10.6151
R1631 B.n911 B.n910 10.6151
R1632 B.n910 B.n909 10.6151
R1633 B.n909 B.n45 10.6151
R1634 B.n903 B.n45 10.6151
R1635 B.n903 B.n902 10.6151
R1636 B.n902 B.n901 10.6151
R1637 B.n901 B.n52 10.6151
R1638 B.n895 B.n52 10.6151
R1639 B.n895 B.n894 10.6151
R1640 B.n894 B.n893 10.6151
R1641 B.n893 B.n59 10.6151
R1642 B.n887 B.n59 10.6151
R1643 B.n887 B.n886 10.6151
R1644 B.n886 B.n885 10.6151
R1645 B.n885 B.n66 10.6151
R1646 B.n879 B.n66 10.6151
R1647 B.n879 B.n878 10.6151
R1648 B.n878 B.n877 10.6151
R1649 B.n877 B.n73 10.6151
R1650 B.n871 B.n73 10.6151
R1651 B.n871 B.n870 10.6151
R1652 B.n870 B.n869 10.6151
R1653 B.n869 B.n80 10.6151
R1654 B.n863 B.n80 10.6151
R1655 B.n111 B.n107 9.36635
R1656 B.n757 B.n756 9.36635
R1657 B.n388 B.n387 9.36635
R1658 B.n365 B.n261 9.36635
R1659 B.n589 B.t0 3.08779
R1660 B.n939 B.t1 3.08779
R1661 B.n957 B.n0 2.81026
R1662 B.n957 B.n1 2.81026
R1663 B.n775 B.n111 1.24928
R1664 B.n758 B.n757 1.24928
R1665 B.n387 B.n386 1.24928
R1666 B.n369 B.n261 1.24928
R1667 VP.n18 VP.n0 161.3
R1668 VP.n17 VP.n16 161.3
R1669 VP.n15 VP.n1 161.3
R1670 VP.n14 VP.n13 161.3
R1671 VP.n12 VP.n2 161.3
R1672 VP.n11 VP.n10 161.3
R1673 VP.n9 VP.n3 161.3
R1674 VP.n8 VP.n7 161.3
R1675 VP.n4 VP.t1 110.007
R1676 VP.n4 VP.t0 108.569
R1677 VP.n6 VP.t2 76.1249
R1678 VP.n19 VP.t3 76.1249
R1679 VP.n6 VP.n5 62.7064
R1680 VP.n20 VP.n19 62.7064
R1681 VP.n13 VP.n12 56.5617
R1682 VP.n5 VP.n4 52.7776
R1683 VP.n7 VP.n3 24.5923
R1684 VP.n11 VP.n3 24.5923
R1685 VP.n12 VP.n11 24.5923
R1686 VP.n13 VP.n1 24.5923
R1687 VP.n17 VP.n1 24.5923
R1688 VP.n18 VP.n17 24.5923
R1689 VP.n7 VP.n6 19.674
R1690 VP.n19 VP.n18 19.674
R1691 VP.n8 VP.n5 0.417304
R1692 VP.n20 VP.n0 0.417304
R1693 VP VP.n20 0.394524
R1694 VP.n9 VP.n8 0.189894
R1695 VP.n10 VP.n9 0.189894
R1696 VP.n10 VP.n2 0.189894
R1697 VP.n14 VP.n2 0.189894
R1698 VP.n15 VP.n14 0.189894
R1699 VP.n16 VP.n15 0.189894
R1700 VP.n16 VP.n0 0.189894
R1701 VDD1 VDD1.n1 109.121
R1702 VDD1 VDD1.n0 63.0092
R1703 VDD1.n0 VDD1.t2 1.57945
R1704 VDD1.n0 VDD1.t3 1.57945
R1705 VDD1.n1 VDD1.t1 1.57945
R1706 VDD1.n1 VDD1.t0 1.57945
C0 VTAIL VDD1 5.92431f
C1 VN VP 7.27639f
C2 VTAIL VDD2 5.9877f
C3 VDD1 VDD2 1.3641f
C4 VN VTAIL 5.36103f
C5 VN VDD1 0.15073f
C6 VTAIL VP 5.37514f
C7 VN VDD2 5.26967f
C8 VP VDD1 5.59983f
C9 VP VDD2 0.481973f
C10 VDD2 B 4.583461f
C11 VDD1 B 9.29675f
C12 VTAIL B 11.148631f
C13 VN B 13.419359f
C14 VP B 11.903472f
C15 VDD1.t2 B 0.273909f
C16 VDD1.t3 B 0.273909f
C17 VDD1.n0 B 2.44872f
C18 VDD1.t1 B 0.273909f
C19 VDD1.t0 B 0.273909f
C20 VDD1.n1 B 3.25674f
C21 VP.n0 B 0.036956f
C22 VP.t3 B 2.66899f
C23 VP.n1 B 0.036444f
C24 VP.n2 B 0.019652f
C25 VP.n3 B 0.036444f
C26 VP.t0 B 2.99253f
C27 VP.t1 B 3.00618f
C28 VP.n4 B 3.10788f
C29 VP.n5 B 1.24077f
C30 VP.t2 B 2.66899f
C31 VP.n6 B 1.01662f
C32 VP.n7 B 0.032846f
C33 VP.n8 B 0.036956f
C34 VP.n9 B 0.019652f
C35 VP.n10 B 0.019652f
C36 VP.n11 B 0.036444f
C37 VP.n12 B 0.028568f
C38 VP.n13 B 0.028568f
C39 VP.n14 B 0.019652f
C40 VP.n15 B 0.019652f
C41 VP.n16 B 0.019652f
C42 VP.n17 B 0.036444f
C43 VP.n18 B 0.032846f
C44 VP.n19 B 1.01662f
C45 VP.n20 B 0.063235f
C46 VTAIL.t4 B 1.87518f
C47 VTAIL.n0 B 0.358246f
C48 VTAIL.t0 B 1.87518f
C49 VTAIL.n1 B 0.457495f
C50 VTAIL.t2 B 1.87518f
C51 VTAIL.n2 B 1.46715f
C52 VTAIL.t7 B 1.87519f
C53 VTAIL.n3 B 1.46714f
C54 VTAIL.t6 B 1.87519f
C55 VTAIL.n4 B 0.457483f
C56 VTAIL.t1 B 1.87519f
C57 VTAIL.n5 B 0.457483f
C58 VTAIL.t3 B 1.87518f
C59 VTAIL.n6 B 1.46715f
C60 VTAIL.t5 B 1.87518f
C61 VTAIL.n7 B 1.36147f
C62 VDD2.t2 B 0.271556f
C63 VDD2.t3 B 0.271556f
C64 VDD2.n0 B 3.20087f
C65 VDD2.t1 B 0.271556f
C66 VDD2.t0 B 0.271556f
C67 VDD2.n1 B 2.42716f
C68 VDD2.n2 B 4.25253f
C69 VN.t3 B 2.95244f
C70 VN.t2 B 2.93904f
C71 VN.n0 B 1.75163f
C72 VN.t1 B 2.95244f
C73 VN.t0 B 2.93904f
C74 VN.n1 B 3.05716f
.ends

