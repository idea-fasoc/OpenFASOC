* NGSPICE file created from diff_pair_sample_1131.ext - technology: sky130A

.subckt diff_pair_sample_1131 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t5 VP.t0 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.8578 pd=30.82 as=2.4783 ps=15.35 w=15.02 l=1.47
X1 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=5.8578 pd=30.82 as=0 ps=0 w=15.02 l=1.47
X2 VDD1.t3 VP.t1 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.4783 pd=15.35 as=5.8578 ps=30.82 w=15.02 l=1.47
X3 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=5.8578 pd=30.82 as=0 ps=0 w=15.02 l=1.47
X4 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.8578 pd=30.82 as=0 ps=0 w=15.02 l=1.47
X5 VTAIL.t1 VN.t0 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=5.8578 pd=30.82 as=2.4783 ps=15.35 w=15.02 l=1.47
X6 VDD1.t0 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.4783 pd=15.35 as=5.8578 ps=30.82 w=15.02 l=1.47
X7 VTAIL.t7 VN.t1 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=5.8578 pd=30.82 as=2.4783 ps=15.35 w=15.02 l=1.47
X8 VTAIL.t2 VP.t3 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=5.8578 pd=30.82 as=2.4783 ps=15.35 w=15.02 l=1.47
X9 VDD2.t1 VN.t2 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.4783 pd=15.35 as=5.8578 ps=30.82 w=15.02 l=1.47
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.8578 pd=30.82 as=0 ps=0 w=15.02 l=1.47
X11 VDD2.t0 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.4783 pd=15.35 as=5.8578 ps=30.82 w=15.02 l=1.47
R0 VP.n2 VP.t3 282.248
R1 VP.n2 VP.t1 281.933
R2 VP.n4 VP.t0 246.246
R3 VP.n11 VP.t2 246.246
R4 VP.n4 VP.n3 178.514
R5 VP.n12 VP.n11 178.514
R6 VP.n10 VP.n0 161.3
R7 VP.n9 VP.n8 161.3
R8 VP.n7 VP.n1 161.3
R9 VP.n6 VP.n5 161.3
R10 VP.n3 VP.n2 58.1439
R11 VP.n9 VP.n1 56.5617
R12 VP.n5 VP.n1 24.5923
R13 VP.n10 VP.n9 24.5923
R14 VP.n5 VP.n4 7.37805
R15 VP.n11 VP.n10 7.37805
R16 VP.n6 VP.n3 0.189894
R17 VP.n7 VP.n6 0.189894
R18 VP.n8 VP.n7 0.189894
R19 VP.n8 VP.n0 0.189894
R20 VP.n12 VP.n0 0.189894
R21 VP VP.n12 0.0516364
R22 VDD1 VDD1.n1 103.111
R23 VDD1 VDD1.n0 61.3257
R24 VDD1.n0 VDD1.t2 1.31874
R25 VDD1.n0 VDD1.t3 1.31874
R26 VDD1.n1 VDD1.t1 1.31874
R27 VDD1.n1 VDD1.t0 1.31874
R28 VTAIL.n5 VTAIL.t2 45.9071
R29 VTAIL.n4 VTAIL.t6 45.9071
R30 VTAIL.n3 VTAIL.t1 45.9071
R31 VTAIL.n7 VTAIL.t0 45.9069
R32 VTAIL.n0 VTAIL.t7 45.9069
R33 VTAIL.n1 VTAIL.t3 45.9069
R34 VTAIL.n2 VTAIL.t5 45.9069
R35 VTAIL.n6 VTAIL.t4 45.9069
R36 VTAIL.n7 VTAIL.n6 26.8669
R37 VTAIL.n3 VTAIL.n2 26.8669
R38 VTAIL.n4 VTAIL.n3 1.55222
R39 VTAIL.n6 VTAIL.n5 1.55222
R40 VTAIL.n2 VTAIL.n1 1.55222
R41 VTAIL VTAIL.n0 0.834552
R42 VTAIL VTAIL.n7 0.718172
R43 VTAIL.n5 VTAIL.n4 0.470328
R44 VTAIL.n1 VTAIL.n0 0.470328
R45 B.n760 B.n759 585
R46 B.n761 B.n760 585
R47 B.n326 B.n103 585
R48 B.n325 B.n324 585
R49 B.n323 B.n322 585
R50 B.n321 B.n320 585
R51 B.n319 B.n318 585
R52 B.n317 B.n316 585
R53 B.n315 B.n314 585
R54 B.n313 B.n312 585
R55 B.n311 B.n310 585
R56 B.n309 B.n308 585
R57 B.n307 B.n306 585
R58 B.n305 B.n304 585
R59 B.n303 B.n302 585
R60 B.n301 B.n300 585
R61 B.n299 B.n298 585
R62 B.n297 B.n296 585
R63 B.n295 B.n294 585
R64 B.n293 B.n292 585
R65 B.n291 B.n290 585
R66 B.n289 B.n288 585
R67 B.n287 B.n286 585
R68 B.n285 B.n284 585
R69 B.n283 B.n282 585
R70 B.n281 B.n280 585
R71 B.n279 B.n278 585
R72 B.n277 B.n276 585
R73 B.n275 B.n274 585
R74 B.n273 B.n272 585
R75 B.n271 B.n270 585
R76 B.n269 B.n268 585
R77 B.n267 B.n266 585
R78 B.n265 B.n264 585
R79 B.n263 B.n262 585
R80 B.n261 B.n260 585
R81 B.n259 B.n258 585
R82 B.n257 B.n256 585
R83 B.n255 B.n254 585
R84 B.n253 B.n252 585
R85 B.n251 B.n250 585
R86 B.n249 B.n248 585
R87 B.n247 B.n246 585
R88 B.n245 B.n244 585
R89 B.n243 B.n242 585
R90 B.n241 B.n240 585
R91 B.n239 B.n238 585
R92 B.n237 B.n236 585
R93 B.n235 B.n234 585
R94 B.n233 B.n232 585
R95 B.n231 B.n230 585
R96 B.n229 B.n228 585
R97 B.n227 B.n226 585
R98 B.n225 B.n224 585
R99 B.n223 B.n222 585
R100 B.n221 B.n220 585
R101 B.n219 B.n218 585
R102 B.n217 B.n216 585
R103 B.n215 B.n214 585
R104 B.n213 B.n212 585
R105 B.n211 B.n210 585
R106 B.n208 B.n207 585
R107 B.n206 B.n205 585
R108 B.n204 B.n203 585
R109 B.n202 B.n201 585
R110 B.n200 B.n199 585
R111 B.n198 B.n197 585
R112 B.n196 B.n195 585
R113 B.n194 B.n193 585
R114 B.n192 B.n191 585
R115 B.n190 B.n189 585
R116 B.n188 B.n187 585
R117 B.n186 B.n185 585
R118 B.n184 B.n183 585
R119 B.n182 B.n181 585
R120 B.n180 B.n179 585
R121 B.n178 B.n177 585
R122 B.n176 B.n175 585
R123 B.n174 B.n173 585
R124 B.n172 B.n171 585
R125 B.n170 B.n169 585
R126 B.n168 B.n167 585
R127 B.n166 B.n165 585
R128 B.n164 B.n163 585
R129 B.n162 B.n161 585
R130 B.n160 B.n159 585
R131 B.n158 B.n157 585
R132 B.n156 B.n155 585
R133 B.n154 B.n153 585
R134 B.n152 B.n151 585
R135 B.n150 B.n149 585
R136 B.n148 B.n147 585
R137 B.n146 B.n145 585
R138 B.n144 B.n143 585
R139 B.n142 B.n141 585
R140 B.n140 B.n139 585
R141 B.n138 B.n137 585
R142 B.n136 B.n135 585
R143 B.n134 B.n133 585
R144 B.n132 B.n131 585
R145 B.n130 B.n129 585
R146 B.n128 B.n127 585
R147 B.n126 B.n125 585
R148 B.n124 B.n123 585
R149 B.n122 B.n121 585
R150 B.n120 B.n119 585
R151 B.n118 B.n117 585
R152 B.n116 B.n115 585
R153 B.n114 B.n113 585
R154 B.n112 B.n111 585
R155 B.n110 B.n109 585
R156 B.n46 B.n45 585
R157 B.n758 B.n47 585
R158 B.n762 B.n47 585
R159 B.n757 B.n756 585
R160 B.n756 B.n43 585
R161 B.n755 B.n42 585
R162 B.n768 B.n42 585
R163 B.n754 B.n41 585
R164 B.n769 B.n41 585
R165 B.n753 B.n40 585
R166 B.n770 B.n40 585
R167 B.n752 B.n751 585
R168 B.n751 B.n39 585
R169 B.n750 B.n35 585
R170 B.n776 B.n35 585
R171 B.n749 B.n34 585
R172 B.n777 B.n34 585
R173 B.n748 B.n33 585
R174 B.n778 B.n33 585
R175 B.n747 B.n746 585
R176 B.n746 B.n29 585
R177 B.n745 B.n28 585
R178 B.n784 B.n28 585
R179 B.n744 B.n27 585
R180 B.n785 B.n27 585
R181 B.n743 B.n26 585
R182 B.n786 B.n26 585
R183 B.n742 B.n741 585
R184 B.n741 B.n22 585
R185 B.n740 B.n21 585
R186 B.n792 B.n21 585
R187 B.n739 B.n20 585
R188 B.n793 B.n20 585
R189 B.n738 B.n19 585
R190 B.n794 B.n19 585
R191 B.n737 B.n736 585
R192 B.n736 B.n15 585
R193 B.n735 B.n14 585
R194 B.n800 B.n14 585
R195 B.n734 B.n13 585
R196 B.n801 B.n13 585
R197 B.n733 B.n12 585
R198 B.n802 B.n12 585
R199 B.n732 B.n731 585
R200 B.n731 B.n8 585
R201 B.n730 B.n7 585
R202 B.n808 B.n7 585
R203 B.n729 B.n6 585
R204 B.n809 B.n6 585
R205 B.n728 B.n5 585
R206 B.n810 B.n5 585
R207 B.n727 B.n726 585
R208 B.n726 B.n4 585
R209 B.n725 B.n327 585
R210 B.n725 B.n724 585
R211 B.n715 B.n328 585
R212 B.n329 B.n328 585
R213 B.n717 B.n716 585
R214 B.n718 B.n717 585
R215 B.n714 B.n333 585
R216 B.n337 B.n333 585
R217 B.n713 B.n712 585
R218 B.n712 B.n711 585
R219 B.n335 B.n334 585
R220 B.n336 B.n335 585
R221 B.n704 B.n703 585
R222 B.n705 B.n704 585
R223 B.n702 B.n342 585
R224 B.n342 B.n341 585
R225 B.n701 B.n700 585
R226 B.n700 B.n699 585
R227 B.n344 B.n343 585
R228 B.n345 B.n344 585
R229 B.n692 B.n691 585
R230 B.n693 B.n692 585
R231 B.n690 B.n350 585
R232 B.n350 B.n349 585
R233 B.n689 B.n688 585
R234 B.n688 B.n687 585
R235 B.n352 B.n351 585
R236 B.n353 B.n352 585
R237 B.n680 B.n679 585
R238 B.n681 B.n680 585
R239 B.n678 B.n358 585
R240 B.n358 B.n357 585
R241 B.n677 B.n676 585
R242 B.n676 B.n675 585
R243 B.n360 B.n359 585
R244 B.n668 B.n360 585
R245 B.n667 B.n666 585
R246 B.n669 B.n667 585
R247 B.n665 B.n365 585
R248 B.n365 B.n364 585
R249 B.n664 B.n663 585
R250 B.n663 B.n662 585
R251 B.n367 B.n366 585
R252 B.n368 B.n367 585
R253 B.n655 B.n654 585
R254 B.n656 B.n655 585
R255 B.n371 B.n370 585
R256 B.n432 B.n431 585
R257 B.n433 B.n429 585
R258 B.n429 B.n372 585
R259 B.n435 B.n434 585
R260 B.n437 B.n428 585
R261 B.n440 B.n439 585
R262 B.n441 B.n427 585
R263 B.n443 B.n442 585
R264 B.n445 B.n426 585
R265 B.n448 B.n447 585
R266 B.n449 B.n425 585
R267 B.n451 B.n450 585
R268 B.n453 B.n424 585
R269 B.n456 B.n455 585
R270 B.n457 B.n423 585
R271 B.n459 B.n458 585
R272 B.n461 B.n422 585
R273 B.n464 B.n463 585
R274 B.n465 B.n421 585
R275 B.n467 B.n466 585
R276 B.n469 B.n420 585
R277 B.n472 B.n471 585
R278 B.n473 B.n419 585
R279 B.n475 B.n474 585
R280 B.n477 B.n418 585
R281 B.n480 B.n479 585
R282 B.n481 B.n417 585
R283 B.n483 B.n482 585
R284 B.n485 B.n416 585
R285 B.n488 B.n487 585
R286 B.n489 B.n415 585
R287 B.n491 B.n490 585
R288 B.n493 B.n414 585
R289 B.n496 B.n495 585
R290 B.n497 B.n413 585
R291 B.n499 B.n498 585
R292 B.n501 B.n412 585
R293 B.n504 B.n503 585
R294 B.n505 B.n411 585
R295 B.n507 B.n506 585
R296 B.n509 B.n410 585
R297 B.n512 B.n511 585
R298 B.n513 B.n409 585
R299 B.n515 B.n514 585
R300 B.n517 B.n408 585
R301 B.n520 B.n519 585
R302 B.n521 B.n407 585
R303 B.n523 B.n522 585
R304 B.n525 B.n406 585
R305 B.n528 B.n527 585
R306 B.n529 B.n403 585
R307 B.n532 B.n531 585
R308 B.n534 B.n402 585
R309 B.n537 B.n536 585
R310 B.n538 B.n401 585
R311 B.n540 B.n539 585
R312 B.n542 B.n400 585
R313 B.n545 B.n544 585
R314 B.n546 B.n399 585
R315 B.n551 B.n550 585
R316 B.n553 B.n398 585
R317 B.n556 B.n555 585
R318 B.n557 B.n397 585
R319 B.n559 B.n558 585
R320 B.n561 B.n396 585
R321 B.n564 B.n563 585
R322 B.n565 B.n395 585
R323 B.n567 B.n566 585
R324 B.n569 B.n394 585
R325 B.n572 B.n571 585
R326 B.n573 B.n393 585
R327 B.n575 B.n574 585
R328 B.n577 B.n392 585
R329 B.n580 B.n579 585
R330 B.n581 B.n391 585
R331 B.n583 B.n582 585
R332 B.n585 B.n390 585
R333 B.n588 B.n587 585
R334 B.n589 B.n389 585
R335 B.n591 B.n590 585
R336 B.n593 B.n388 585
R337 B.n596 B.n595 585
R338 B.n597 B.n387 585
R339 B.n599 B.n598 585
R340 B.n601 B.n386 585
R341 B.n604 B.n603 585
R342 B.n605 B.n385 585
R343 B.n607 B.n606 585
R344 B.n609 B.n384 585
R345 B.n612 B.n611 585
R346 B.n613 B.n383 585
R347 B.n615 B.n614 585
R348 B.n617 B.n382 585
R349 B.n620 B.n619 585
R350 B.n621 B.n381 585
R351 B.n623 B.n622 585
R352 B.n625 B.n380 585
R353 B.n628 B.n627 585
R354 B.n629 B.n379 585
R355 B.n631 B.n630 585
R356 B.n633 B.n378 585
R357 B.n636 B.n635 585
R358 B.n637 B.n377 585
R359 B.n639 B.n638 585
R360 B.n641 B.n376 585
R361 B.n644 B.n643 585
R362 B.n645 B.n375 585
R363 B.n647 B.n646 585
R364 B.n649 B.n374 585
R365 B.n652 B.n651 585
R366 B.n653 B.n373 585
R367 B.n658 B.n657 585
R368 B.n657 B.n656 585
R369 B.n659 B.n369 585
R370 B.n369 B.n368 585
R371 B.n661 B.n660 585
R372 B.n662 B.n661 585
R373 B.n363 B.n362 585
R374 B.n364 B.n363 585
R375 B.n671 B.n670 585
R376 B.n670 B.n669 585
R377 B.n672 B.n361 585
R378 B.n668 B.n361 585
R379 B.n674 B.n673 585
R380 B.n675 B.n674 585
R381 B.n356 B.n355 585
R382 B.n357 B.n356 585
R383 B.n683 B.n682 585
R384 B.n682 B.n681 585
R385 B.n684 B.n354 585
R386 B.n354 B.n353 585
R387 B.n686 B.n685 585
R388 B.n687 B.n686 585
R389 B.n348 B.n347 585
R390 B.n349 B.n348 585
R391 B.n695 B.n694 585
R392 B.n694 B.n693 585
R393 B.n696 B.n346 585
R394 B.n346 B.n345 585
R395 B.n698 B.n697 585
R396 B.n699 B.n698 585
R397 B.n340 B.n339 585
R398 B.n341 B.n340 585
R399 B.n707 B.n706 585
R400 B.n706 B.n705 585
R401 B.n708 B.n338 585
R402 B.n338 B.n336 585
R403 B.n710 B.n709 585
R404 B.n711 B.n710 585
R405 B.n332 B.n331 585
R406 B.n337 B.n332 585
R407 B.n720 B.n719 585
R408 B.n719 B.n718 585
R409 B.n721 B.n330 585
R410 B.n330 B.n329 585
R411 B.n723 B.n722 585
R412 B.n724 B.n723 585
R413 B.n2 B.n0 585
R414 B.n4 B.n2 585
R415 B.n3 B.n1 585
R416 B.n809 B.n3 585
R417 B.n807 B.n806 585
R418 B.n808 B.n807 585
R419 B.n805 B.n9 585
R420 B.n9 B.n8 585
R421 B.n804 B.n803 585
R422 B.n803 B.n802 585
R423 B.n11 B.n10 585
R424 B.n801 B.n11 585
R425 B.n799 B.n798 585
R426 B.n800 B.n799 585
R427 B.n797 B.n16 585
R428 B.n16 B.n15 585
R429 B.n796 B.n795 585
R430 B.n795 B.n794 585
R431 B.n18 B.n17 585
R432 B.n793 B.n18 585
R433 B.n791 B.n790 585
R434 B.n792 B.n791 585
R435 B.n789 B.n23 585
R436 B.n23 B.n22 585
R437 B.n788 B.n787 585
R438 B.n787 B.n786 585
R439 B.n25 B.n24 585
R440 B.n785 B.n25 585
R441 B.n783 B.n782 585
R442 B.n784 B.n783 585
R443 B.n781 B.n30 585
R444 B.n30 B.n29 585
R445 B.n780 B.n779 585
R446 B.n779 B.n778 585
R447 B.n32 B.n31 585
R448 B.n777 B.n32 585
R449 B.n775 B.n774 585
R450 B.n776 B.n775 585
R451 B.n773 B.n36 585
R452 B.n39 B.n36 585
R453 B.n772 B.n771 585
R454 B.n771 B.n770 585
R455 B.n38 B.n37 585
R456 B.n769 B.n38 585
R457 B.n767 B.n766 585
R458 B.n768 B.n767 585
R459 B.n765 B.n44 585
R460 B.n44 B.n43 585
R461 B.n764 B.n763 585
R462 B.n763 B.n762 585
R463 B.n812 B.n811 585
R464 B.n811 B.n810 585
R465 B.n657 B.n371 463.671
R466 B.n763 B.n46 463.671
R467 B.n655 B.n373 463.671
R468 B.n760 B.n47 463.671
R469 B.n547 B.t15 451.572
R470 B.n404 B.t4 451.572
R471 B.n107 B.t8 451.572
R472 B.n104 B.t12 451.572
R473 B.n761 B.n102 256.663
R474 B.n761 B.n101 256.663
R475 B.n761 B.n100 256.663
R476 B.n761 B.n99 256.663
R477 B.n761 B.n98 256.663
R478 B.n761 B.n97 256.663
R479 B.n761 B.n96 256.663
R480 B.n761 B.n95 256.663
R481 B.n761 B.n94 256.663
R482 B.n761 B.n93 256.663
R483 B.n761 B.n92 256.663
R484 B.n761 B.n91 256.663
R485 B.n761 B.n90 256.663
R486 B.n761 B.n89 256.663
R487 B.n761 B.n88 256.663
R488 B.n761 B.n87 256.663
R489 B.n761 B.n86 256.663
R490 B.n761 B.n85 256.663
R491 B.n761 B.n84 256.663
R492 B.n761 B.n83 256.663
R493 B.n761 B.n82 256.663
R494 B.n761 B.n81 256.663
R495 B.n761 B.n80 256.663
R496 B.n761 B.n79 256.663
R497 B.n761 B.n78 256.663
R498 B.n761 B.n77 256.663
R499 B.n761 B.n76 256.663
R500 B.n761 B.n75 256.663
R501 B.n761 B.n74 256.663
R502 B.n761 B.n73 256.663
R503 B.n761 B.n72 256.663
R504 B.n761 B.n71 256.663
R505 B.n761 B.n70 256.663
R506 B.n761 B.n69 256.663
R507 B.n761 B.n68 256.663
R508 B.n761 B.n67 256.663
R509 B.n761 B.n66 256.663
R510 B.n761 B.n65 256.663
R511 B.n761 B.n64 256.663
R512 B.n761 B.n63 256.663
R513 B.n761 B.n62 256.663
R514 B.n761 B.n61 256.663
R515 B.n761 B.n60 256.663
R516 B.n761 B.n59 256.663
R517 B.n761 B.n58 256.663
R518 B.n761 B.n57 256.663
R519 B.n761 B.n56 256.663
R520 B.n761 B.n55 256.663
R521 B.n761 B.n54 256.663
R522 B.n761 B.n53 256.663
R523 B.n761 B.n52 256.663
R524 B.n761 B.n51 256.663
R525 B.n761 B.n50 256.663
R526 B.n761 B.n49 256.663
R527 B.n761 B.n48 256.663
R528 B.n430 B.n372 256.663
R529 B.n436 B.n372 256.663
R530 B.n438 B.n372 256.663
R531 B.n444 B.n372 256.663
R532 B.n446 B.n372 256.663
R533 B.n452 B.n372 256.663
R534 B.n454 B.n372 256.663
R535 B.n460 B.n372 256.663
R536 B.n462 B.n372 256.663
R537 B.n468 B.n372 256.663
R538 B.n470 B.n372 256.663
R539 B.n476 B.n372 256.663
R540 B.n478 B.n372 256.663
R541 B.n484 B.n372 256.663
R542 B.n486 B.n372 256.663
R543 B.n492 B.n372 256.663
R544 B.n494 B.n372 256.663
R545 B.n500 B.n372 256.663
R546 B.n502 B.n372 256.663
R547 B.n508 B.n372 256.663
R548 B.n510 B.n372 256.663
R549 B.n516 B.n372 256.663
R550 B.n518 B.n372 256.663
R551 B.n524 B.n372 256.663
R552 B.n526 B.n372 256.663
R553 B.n533 B.n372 256.663
R554 B.n535 B.n372 256.663
R555 B.n541 B.n372 256.663
R556 B.n543 B.n372 256.663
R557 B.n552 B.n372 256.663
R558 B.n554 B.n372 256.663
R559 B.n560 B.n372 256.663
R560 B.n562 B.n372 256.663
R561 B.n568 B.n372 256.663
R562 B.n570 B.n372 256.663
R563 B.n576 B.n372 256.663
R564 B.n578 B.n372 256.663
R565 B.n584 B.n372 256.663
R566 B.n586 B.n372 256.663
R567 B.n592 B.n372 256.663
R568 B.n594 B.n372 256.663
R569 B.n600 B.n372 256.663
R570 B.n602 B.n372 256.663
R571 B.n608 B.n372 256.663
R572 B.n610 B.n372 256.663
R573 B.n616 B.n372 256.663
R574 B.n618 B.n372 256.663
R575 B.n624 B.n372 256.663
R576 B.n626 B.n372 256.663
R577 B.n632 B.n372 256.663
R578 B.n634 B.n372 256.663
R579 B.n640 B.n372 256.663
R580 B.n642 B.n372 256.663
R581 B.n648 B.n372 256.663
R582 B.n650 B.n372 256.663
R583 B.n657 B.n369 163.367
R584 B.n661 B.n369 163.367
R585 B.n661 B.n363 163.367
R586 B.n670 B.n363 163.367
R587 B.n670 B.n361 163.367
R588 B.n674 B.n361 163.367
R589 B.n674 B.n356 163.367
R590 B.n682 B.n356 163.367
R591 B.n682 B.n354 163.367
R592 B.n686 B.n354 163.367
R593 B.n686 B.n348 163.367
R594 B.n694 B.n348 163.367
R595 B.n694 B.n346 163.367
R596 B.n698 B.n346 163.367
R597 B.n698 B.n340 163.367
R598 B.n706 B.n340 163.367
R599 B.n706 B.n338 163.367
R600 B.n710 B.n338 163.367
R601 B.n710 B.n332 163.367
R602 B.n719 B.n332 163.367
R603 B.n719 B.n330 163.367
R604 B.n723 B.n330 163.367
R605 B.n723 B.n2 163.367
R606 B.n811 B.n2 163.367
R607 B.n811 B.n3 163.367
R608 B.n807 B.n3 163.367
R609 B.n807 B.n9 163.367
R610 B.n803 B.n9 163.367
R611 B.n803 B.n11 163.367
R612 B.n799 B.n11 163.367
R613 B.n799 B.n16 163.367
R614 B.n795 B.n16 163.367
R615 B.n795 B.n18 163.367
R616 B.n791 B.n18 163.367
R617 B.n791 B.n23 163.367
R618 B.n787 B.n23 163.367
R619 B.n787 B.n25 163.367
R620 B.n783 B.n25 163.367
R621 B.n783 B.n30 163.367
R622 B.n779 B.n30 163.367
R623 B.n779 B.n32 163.367
R624 B.n775 B.n32 163.367
R625 B.n775 B.n36 163.367
R626 B.n771 B.n36 163.367
R627 B.n771 B.n38 163.367
R628 B.n767 B.n38 163.367
R629 B.n767 B.n44 163.367
R630 B.n763 B.n44 163.367
R631 B.n431 B.n429 163.367
R632 B.n435 B.n429 163.367
R633 B.n439 B.n437 163.367
R634 B.n443 B.n427 163.367
R635 B.n447 B.n445 163.367
R636 B.n451 B.n425 163.367
R637 B.n455 B.n453 163.367
R638 B.n459 B.n423 163.367
R639 B.n463 B.n461 163.367
R640 B.n467 B.n421 163.367
R641 B.n471 B.n469 163.367
R642 B.n475 B.n419 163.367
R643 B.n479 B.n477 163.367
R644 B.n483 B.n417 163.367
R645 B.n487 B.n485 163.367
R646 B.n491 B.n415 163.367
R647 B.n495 B.n493 163.367
R648 B.n499 B.n413 163.367
R649 B.n503 B.n501 163.367
R650 B.n507 B.n411 163.367
R651 B.n511 B.n509 163.367
R652 B.n515 B.n409 163.367
R653 B.n519 B.n517 163.367
R654 B.n523 B.n407 163.367
R655 B.n527 B.n525 163.367
R656 B.n532 B.n403 163.367
R657 B.n536 B.n534 163.367
R658 B.n540 B.n401 163.367
R659 B.n544 B.n542 163.367
R660 B.n551 B.n399 163.367
R661 B.n555 B.n553 163.367
R662 B.n559 B.n397 163.367
R663 B.n563 B.n561 163.367
R664 B.n567 B.n395 163.367
R665 B.n571 B.n569 163.367
R666 B.n575 B.n393 163.367
R667 B.n579 B.n577 163.367
R668 B.n583 B.n391 163.367
R669 B.n587 B.n585 163.367
R670 B.n591 B.n389 163.367
R671 B.n595 B.n593 163.367
R672 B.n599 B.n387 163.367
R673 B.n603 B.n601 163.367
R674 B.n607 B.n385 163.367
R675 B.n611 B.n609 163.367
R676 B.n615 B.n383 163.367
R677 B.n619 B.n617 163.367
R678 B.n623 B.n381 163.367
R679 B.n627 B.n625 163.367
R680 B.n631 B.n379 163.367
R681 B.n635 B.n633 163.367
R682 B.n639 B.n377 163.367
R683 B.n643 B.n641 163.367
R684 B.n647 B.n375 163.367
R685 B.n651 B.n649 163.367
R686 B.n655 B.n367 163.367
R687 B.n663 B.n367 163.367
R688 B.n663 B.n365 163.367
R689 B.n667 B.n365 163.367
R690 B.n667 B.n360 163.367
R691 B.n676 B.n360 163.367
R692 B.n676 B.n358 163.367
R693 B.n680 B.n358 163.367
R694 B.n680 B.n352 163.367
R695 B.n688 B.n352 163.367
R696 B.n688 B.n350 163.367
R697 B.n692 B.n350 163.367
R698 B.n692 B.n344 163.367
R699 B.n700 B.n344 163.367
R700 B.n700 B.n342 163.367
R701 B.n704 B.n342 163.367
R702 B.n704 B.n335 163.367
R703 B.n712 B.n335 163.367
R704 B.n712 B.n333 163.367
R705 B.n717 B.n333 163.367
R706 B.n717 B.n328 163.367
R707 B.n725 B.n328 163.367
R708 B.n726 B.n725 163.367
R709 B.n726 B.n5 163.367
R710 B.n6 B.n5 163.367
R711 B.n7 B.n6 163.367
R712 B.n731 B.n7 163.367
R713 B.n731 B.n12 163.367
R714 B.n13 B.n12 163.367
R715 B.n14 B.n13 163.367
R716 B.n736 B.n14 163.367
R717 B.n736 B.n19 163.367
R718 B.n20 B.n19 163.367
R719 B.n21 B.n20 163.367
R720 B.n741 B.n21 163.367
R721 B.n741 B.n26 163.367
R722 B.n27 B.n26 163.367
R723 B.n28 B.n27 163.367
R724 B.n746 B.n28 163.367
R725 B.n746 B.n33 163.367
R726 B.n34 B.n33 163.367
R727 B.n35 B.n34 163.367
R728 B.n751 B.n35 163.367
R729 B.n751 B.n40 163.367
R730 B.n41 B.n40 163.367
R731 B.n42 B.n41 163.367
R732 B.n756 B.n42 163.367
R733 B.n756 B.n47 163.367
R734 B.n111 B.n110 163.367
R735 B.n115 B.n114 163.367
R736 B.n119 B.n118 163.367
R737 B.n123 B.n122 163.367
R738 B.n127 B.n126 163.367
R739 B.n131 B.n130 163.367
R740 B.n135 B.n134 163.367
R741 B.n139 B.n138 163.367
R742 B.n143 B.n142 163.367
R743 B.n147 B.n146 163.367
R744 B.n151 B.n150 163.367
R745 B.n155 B.n154 163.367
R746 B.n159 B.n158 163.367
R747 B.n163 B.n162 163.367
R748 B.n167 B.n166 163.367
R749 B.n171 B.n170 163.367
R750 B.n175 B.n174 163.367
R751 B.n179 B.n178 163.367
R752 B.n183 B.n182 163.367
R753 B.n187 B.n186 163.367
R754 B.n191 B.n190 163.367
R755 B.n195 B.n194 163.367
R756 B.n199 B.n198 163.367
R757 B.n203 B.n202 163.367
R758 B.n207 B.n206 163.367
R759 B.n212 B.n211 163.367
R760 B.n216 B.n215 163.367
R761 B.n220 B.n219 163.367
R762 B.n224 B.n223 163.367
R763 B.n228 B.n227 163.367
R764 B.n232 B.n231 163.367
R765 B.n236 B.n235 163.367
R766 B.n240 B.n239 163.367
R767 B.n244 B.n243 163.367
R768 B.n248 B.n247 163.367
R769 B.n252 B.n251 163.367
R770 B.n256 B.n255 163.367
R771 B.n260 B.n259 163.367
R772 B.n264 B.n263 163.367
R773 B.n268 B.n267 163.367
R774 B.n272 B.n271 163.367
R775 B.n276 B.n275 163.367
R776 B.n280 B.n279 163.367
R777 B.n284 B.n283 163.367
R778 B.n288 B.n287 163.367
R779 B.n292 B.n291 163.367
R780 B.n296 B.n295 163.367
R781 B.n300 B.n299 163.367
R782 B.n304 B.n303 163.367
R783 B.n308 B.n307 163.367
R784 B.n312 B.n311 163.367
R785 B.n316 B.n315 163.367
R786 B.n320 B.n319 163.367
R787 B.n324 B.n323 163.367
R788 B.n760 B.n103 163.367
R789 B.n547 B.t17 103.535
R790 B.n104 B.t13 103.535
R791 B.n404 B.t7 103.516
R792 B.n107 B.t10 103.516
R793 B.n430 B.n371 71.676
R794 B.n436 B.n435 71.676
R795 B.n439 B.n438 71.676
R796 B.n444 B.n443 71.676
R797 B.n447 B.n446 71.676
R798 B.n452 B.n451 71.676
R799 B.n455 B.n454 71.676
R800 B.n460 B.n459 71.676
R801 B.n463 B.n462 71.676
R802 B.n468 B.n467 71.676
R803 B.n471 B.n470 71.676
R804 B.n476 B.n475 71.676
R805 B.n479 B.n478 71.676
R806 B.n484 B.n483 71.676
R807 B.n487 B.n486 71.676
R808 B.n492 B.n491 71.676
R809 B.n495 B.n494 71.676
R810 B.n500 B.n499 71.676
R811 B.n503 B.n502 71.676
R812 B.n508 B.n507 71.676
R813 B.n511 B.n510 71.676
R814 B.n516 B.n515 71.676
R815 B.n519 B.n518 71.676
R816 B.n524 B.n523 71.676
R817 B.n527 B.n526 71.676
R818 B.n533 B.n532 71.676
R819 B.n536 B.n535 71.676
R820 B.n541 B.n540 71.676
R821 B.n544 B.n543 71.676
R822 B.n552 B.n551 71.676
R823 B.n555 B.n554 71.676
R824 B.n560 B.n559 71.676
R825 B.n563 B.n562 71.676
R826 B.n568 B.n567 71.676
R827 B.n571 B.n570 71.676
R828 B.n576 B.n575 71.676
R829 B.n579 B.n578 71.676
R830 B.n584 B.n583 71.676
R831 B.n587 B.n586 71.676
R832 B.n592 B.n591 71.676
R833 B.n595 B.n594 71.676
R834 B.n600 B.n599 71.676
R835 B.n603 B.n602 71.676
R836 B.n608 B.n607 71.676
R837 B.n611 B.n610 71.676
R838 B.n616 B.n615 71.676
R839 B.n619 B.n618 71.676
R840 B.n624 B.n623 71.676
R841 B.n627 B.n626 71.676
R842 B.n632 B.n631 71.676
R843 B.n635 B.n634 71.676
R844 B.n640 B.n639 71.676
R845 B.n643 B.n642 71.676
R846 B.n648 B.n647 71.676
R847 B.n651 B.n650 71.676
R848 B.n48 B.n46 71.676
R849 B.n111 B.n49 71.676
R850 B.n115 B.n50 71.676
R851 B.n119 B.n51 71.676
R852 B.n123 B.n52 71.676
R853 B.n127 B.n53 71.676
R854 B.n131 B.n54 71.676
R855 B.n135 B.n55 71.676
R856 B.n139 B.n56 71.676
R857 B.n143 B.n57 71.676
R858 B.n147 B.n58 71.676
R859 B.n151 B.n59 71.676
R860 B.n155 B.n60 71.676
R861 B.n159 B.n61 71.676
R862 B.n163 B.n62 71.676
R863 B.n167 B.n63 71.676
R864 B.n171 B.n64 71.676
R865 B.n175 B.n65 71.676
R866 B.n179 B.n66 71.676
R867 B.n183 B.n67 71.676
R868 B.n187 B.n68 71.676
R869 B.n191 B.n69 71.676
R870 B.n195 B.n70 71.676
R871 B.n199 B.n71 71.676
R872 B.n203 B.n72 71.676
R873 B.n207 B.n73 71.676
R874 B.n212 B.n74 71.676
R875 B.n216 B.n75 71.676
R876 B.n220 B.n76 71.676
R877 B.n224 B.n77 71.676
R878 B.n228 B.n78 71.676
R879 B.n232 B.n79 71.676
R880 B.n236 B.n80 71.676
R881 B.n240 B.n81 71.676
R882 B.n244 B.n82 71.676
R883 B.n248 B.n83 71.676
R884 B.n252 B.n84 71.676
R885 B.n256 B.n85 71.676
R886 B.n260 B.n86 71.676
R887 B.n264 B.n87 71.676
R888 B.n268 B.n88 71.676
R889 B.n272 B.n89 71.676
R890 B.n276 B.n90 71.676
R891 B.n280 B.n91 71.676
R892 B.n284 B.n92 71.676
R893 B.n288 B.n93 71.676
R894 B.n292 B.n94 71.676
R895 B.n296 B.n95 71.676
R896 B.n300 B.n96 71.676
R897 B.n304 B.n97 71.676
R898 B.n308 B.n98 71.676
R899 B.n312 B.n99 71.676
R900 B.n316 B.n100 71.676
R901 B.n320 B.n101 71.676
R902 B.n324 B.n102 71.676
R903 B.n103 B.n102 71.676
R904 B.n323 B.n101 71.676
R905 B.n319 B.n100 71.676
R906 B.n315 B.n99 71.676
R907 B.n311 B.n98 71.676
R908 B.n307 B.n97 71.676
R909 B.n303 B.n96 71.676
R910 B.n299 B.n95 71.676
R911 B.n295 B.n94 71.676
R912 B.n291 B.n93 71.676
R913 B.n287 B.n92 71.676
R914 B.n283 B.n91 71.676
R915 B.n279 B.n90 71.676
R916 B.n275 B.n89 71.676
R917 B.n271 B.n88 71.676
R918 B.n267 B.n87 71.676
R919 B.n263 B.n86 71.676
R920 B.n259 B.n85 71.676
R921 B.n255 B.n84 71.676
R922 B.n251 B.n83 71.676
R923 B.n247 B.n82 71.676
R924 B.n243 B.n81 71.676
R925 B.n239 B.n80 71.676
R926 B.n235 B.n79 71.676
R927 B.n231 B.n78 71.676
R928 B.n227 B.n77 71.676
R929 B.n223 B.n76 71.676
R930 B.n219 B.n75 71.676
R931 B.n215 B.n74 71.676
R932 B.n211 B.n73 71.676
R933 B.n206 B.n72 71.676
R934 B.n202 B.n71 71.676
R935 B.n198 B.n70 71.676
R936 B.n194 B.n69 71.676
R937 B.n190 B.n68 71.676
R938 B.n186 B.n67 71.676
R939 B.n182 B.n66 71.676
R940 B.n178 B.n65 71.676
R941 B.n174 B.n64 71.676
R942 B.n170 B.n63 71.676
R943 B.n166 B.n62 71.676
R944 B.n162 B.n61 71.676
R945 B.n158 B.n60 71.676
R946 B.n154 B.n59 71.676
R947 B.n150 B.n58 71.676
R948 B.n146 B.n57 71.676
R949 B.n142 B.n56 71.676
R950 B.n138 B.n55 71.676
R951 B.n134 B.n54 71.676
R952 B.n130 B.n53 71.676
R953 B.n126 B.n52 71.676
R954 B.n122 B.n51 71.676
R955 B.n118 B.n50 71.676
R956 B.n114 B.n49 71.676
R957 B.n110 B.n48 71.676
R958 B.n431 B.n430 71.676
R959 B.n437 B.n436 71.676
R960 B.n438 B.n427 71.676
R961 B.n445 B.n444 71.676
R962 B.n446 B.n425 71.676
R963 B.n453 B.n452 71.676
R964 B.n454 B.n423 71.676
R965 B.n461 B.n460 71.676
R966 B.n462 B.n421 71.676
R967 B.n469 B.n468 71.676
R968 B.n470 B.n419 71.676
R969 B.n477 B.n476 71.676
R970 B.n478 B.n417 71.676
R971 B.n485 B.n484 71.676
R972 B.n486 B.n415 71.676
R973 B.n493 B.n492 71.676
R974 B.n494 B.n413 71.676
R975 B.n501 B.n500 71.676
R976 B.n502 B.n411 71.676
R977 B.n509 B.n508 71.676
R978 B.n510 B.n409 71.676
R979 B.n517 B.n516 71.676
R980 B.n518 B.n407 71.676
R981 B.n525 B.n524 71.676
R982 B.n526 B.n403 71.676
R983 B.n534 B.n533 71.676
R984 B.n535 B.n401 71.676
R985 B.n542 B.n541 71.676
R986 B.n543 B.n399 71.676
R987 B.n553 B.n552 71.676
R988 B.n554 B.n397 71.676
R989 B.n561 B.n560 71.676
R990 B.n562 B.n395 71.676
R991 B.n569 B.n568 71.676
R992 B.n570 B.n393 71.676
R993 B.n577 B.n576 71.676
R994 B.n578 B.n391 71.676
R995 B.n585 B.n584 71.676
R996 B.n586 B.n389 71.676
R997 B.n593 B.n592 71.676
R998 B.n594 B.n387 71.676
R999 B.n601 B.n600 71.676
R1000 B.n602 B.n385 71.676
R1001 B.n609 B.n608 71.676
R1002 B.n610 B.n383 71.676
R1003 B.n617 B.n616 71.676
R1004 B.n618 B.n381 71.676
R1005 B.n625 B.n624 71.676
R1006 B.n626 B.n379 71.676
R1007 B.n633 B.n632 71.676
R1008 B.n634 B.n377 71.676
R1009 B.n641 B.n640 71.676
R1010 B.n642 B.n375 71.676
R1011 B.n649 B.n648 71.676
R1012 B.n650 B.n373 71.676
R1013 B.n548 B.t16 68.6263
R1014 B.n105 B.t14 68.6263
R1015 B.n405 B.t6 68.6065
R1016 B.n108 B.t11 68.6065
R1017 B.n656 B.n372 66.6672
R1018 B.n762 B.n761 66.6672
R1019 B.n549 B.n548 59.5399
R1020 B.n530 B.n405 59.5399
R1021 B.n209 B.n108 59.5399
R1022 B.n106 B.n105 59.5399
R1023 B.n656 B.n368 36.8569
R1024 B.n662 B.n368 36.8569
R1025 B.n662 B.n364 36.8569
R1026 B.n669 B.n364 36.8569
R1027 B.n669 B.n668 36.8569
R1028 B.n675 B.n357 36.8569
R1029 B.n681 B.n357 36.8569
R1030 B.n681 B.n353 36.8569
R1031 B.n687 B.n353 36.8569
R1032 B.n687 B.n349 36.8569
R1033 B.n693 B.n349 36.8569
R1034 B.n693 B.n345 36.8569
R1035 B.n699 B.n345 36.8569
R1036 B.n705 B.n341 36.8569
R1037 B.n705 B.n336 36.8569
R1038 B.n711 B.n336 36.8569
R1039 B.n711 B.n337 36.8569
R1040 B.n718 B.n329 36.8569
R1041 B.n724 B.n329 36.8569
R1042 B.n724 B.n4 36.8569
R1043 B.n810 B.n4 36.8569
R1044 B.n810 B.n809 36.8569
R1045 B.n809 B.n808 36.8569
R1046 B.n808 B.n8 36.8569
R1047 B.n802 B.n8 36.8569
R1048 B.n801 B.n800 36.8569
R1049 B.n800 B.n15 36.8569
R1050 B.n794 B.n15 36.8569
R1051 B.n794 B.n793 36.8569
R1052 B.n792 B.n22 36.8569
R1053 B.n786 B.n22 36.8569
R1054 B.n786 B.n785 36.8569
R1055 B.n785 B.n784 36.8569
R1056 B.n784 B.n29 36.8569
R1057 B.n778 B.n29 36.8569
R1058 B.n778 B.n777 36.8569
R1059 B.n777 B.n776 36.8569
R1060 B.n770 B.n39 36.8569
R1061 B.n770 B.n769 36.8569
R1062 B.n769 B.n768 36.8569
R1063 B.n768 B.n43 36.8569
R1064 B.n762 B.n43 36.8569
R1065 B.n668 B.t5 35.2309
R1066 B.n39 B.t9 35.2309
R1067 B.n548 B.n547 34.9096
R1068 B.n405 B.n404 34.9096
R1069 B.n108 B.n107 34.9096
R1070 B.n105 B.n104 34.9096
R1071 B.n759 B.n758 30.1273
R1072 B.n764 B.n45 30.1273
R1073 B.n654 B.n653 30.1273
R1074 B.n658 B.n370 30.1273
R1075 B.n337 B.t3 27.6428
R1076 B.t2 B.n801 27.6428
R1077 B.t1 B.n341 20.0547
R1078 B.n793 B.t0 20.0547
R1079 B B.n812 18.0485
R1080 B.n699 B.t1 16.8027
R1081 B.t0 B.n792 16.8027
R1082 B.n109 B.n45 10.6151
R1083 B.n112 B.n109 10.6151
R1084 B.n113 B.n112 10.6151
R1085 B.n116 B.n113 10.6151
R1086 B.n117 B.n116 10.6151
R1087 B.n120 B.n117 10.6151
R1088 B.n121 B.n120 10.6151
R1089 B.n124 B.n121 10.6151
R1090 B.n125 B.n124 10.6151
R1091 B.n128 B.n125 10.6151
R1092 B.n129 B.n128 10.6151
R1093 B.n132 B.n129 10.6151
R1094 B.n133 B.n132 10.6151
R1095 B.n136 B.n133 10.6151
R1096 B.n137 B.n136 10.6151
R1097 B.n140 B.n137 10.6151
R1098 B.n141 B.n140 10.6151
R1099 B.n144 B.n141 10.6151
R1100 B.n145 B.n144 10.6151
R1101 B.n148 B.n145 10.6151
R1102 B.n149 B.n148 10.6151
R1103 B.n152 B.n149 10.6151
R1104 B.n153 B.n152 10.6151
R1105 B.n156 B.n153 10.6151
R1106 B.n157 B.n156 10.6151
R1107 B.n160 B.n157 10.6151
R1108 B.n161 B.n160 10.6151
R1109 B.n164 B.n161 10.6151
R1110 B.n165 B.n164 10.6151
R1111 B.n168 B.n165 10.6151
R1112 B.n169 B.n168 10.6151
R1113 B.n172 B.n169 10.6151
R1114 B.n173 B.n172 10.6151
R1115 B.n176 B.n173 10.6151
R1116 B.n177 B.n176 10.6151
R1117 B.n180 B.n177 10.6151
R1118 B.n181 B.n180 10.6151
R1119 B.n184 B.n181 10.6151
R1120 B.n185 B.n184 10.6151
R1121 B.n188 B.n185 10.6151
R1122 B.n189 B.n188 10.6151
R1123 B.n192 B.n189 10.6151
R1124 B.n193 B.n192 10.6151
R1125 B.n196 B.n193 10.6151
R1126 B.n197 B.n196 10.6151
R1127 B.n200 B.n197 10.6151
R1128 B.n201 B.n200 10.6151
R1129 B.n204 B.n201 10.6151
R1130 B.n205 B.n204 10.6151
R1131 B.n208 B.n205 10.6151
R1132 B.n213 B.n210 10.6151
R1133 B.n214 B.n213 10.6151
R1134 B.n217 B.n214 10.6151
R1135 B.n218 B.n217 10.6151
R1136 B.n221 B.n218 10.6151
R1137 B.n222 B.n221 10.6151
R1138 B.n225 B.n222 10.6151
R1139 B.n226 B.n225 10.6151
R1140 B.n230 B.n229 10.6151
R1141 B.n233 B.n230 10.6151
R1142 B.n234 B.n233 10.6151
R1143 B.n237 B.n234 10.6151
R1144 B.n238 B.n237 10.6151
R1145 B.n241 B.n238 10.6151
R1146 B.n242 B.n241 10.6151
R1147 B.n245 B.n242 10.6151
R1148 B.n246 B.n245 10.6151
R1149 B.n249 B.n246 10.6151
R1150 B.n250 B.n249 10.6151
R1151 B.n253 B.n250 10.6151
R1152 B.n254 B.n253 10.6151
R1153 B.n257 B.n254 10.6151
R1154 B.n258 B.n257 10.6151
R1155 B.n261 B.n258 10.6151
R1156 B.n262 B.n261 10.6151
R1157 B.n265 B.n262 10.6151
R1158 B.n266 B.n265 10.6151
R1159 B.n269 B.n266 10.6151
R1160 B.n270 B.n269 10.6151
R1161 B.n273 B.n270 10.6151
R1162 B.n274 B.n273 10.6151
R1163 B.n277 B.n274 10.6151
R1164 B.n278 B.n277 10.6151
R1165 B.n281 B.n278 10.6151
R1166 B.n282 B.n281 10.6151
R1167 B.n285 B.n282 10.6151
R1168 B.n286 B.n285 10.6151
R1169 B.n289 B.n286 10.6151
R1170 B.n290 B.n289 10.6151
R1171 B.n293 B.n290 10.6151
R1172 B.n294 B.n293 10.6151
R1173 B.n297 B.n294 10.6151
R1174 B.n298 B.n297 10.6151
R1175 B.n301 B.n298 10.6151
R1176 B.n302 B.n301 10.6151
R1177 B.n305 B.n302 10.6151
R1178 B.n306 B.n305 10.6151
R1179 B.n309 B.n306 10.6151
R1180 B.n310 B.n309 10.6151
R1181 B.n313 B.n310 10.6151
R1182 B.n314 B.n313 10.6151
R1183 B.n317 B.n314 10.6151
R1184 B.n318 B.n317 10.6151
R1185 B.n321 B.n318 10.6151
R1186 B.n322 B.n321 10.6151
R1187 B.n325 B.n322 10.6151
R1188 B.n326 B.n325 10.6151
R1189 B.n759 B.n326 10.6151
R1190 B.n654 B.n366 10.6151
R1191 B.n664 B.n366 10.6151
R1192 B.n665 B.n664 10.6151
R1193 B.n666 B.n665 10.6151
R1194 B.n666 B.n359 10.6151
R1195 B.n677 B.n359 10.6151
R1196 B.n678 B.n677 10.6151
R1197 B.n679 B.n678 10.6151
R1198 B.n679 B.n351 10.6151
R1199 B.n689 B.n351 10.6151
R1200 B.n690 B.n689 10.6151
R1201 B.n691 B.n690 10.6151
R1202 B.n691 B.n343 10.6151
R1203 B.n701 B.n343 10.6151
R1204 B.n702 B.n701 10.6151
R1205 B.n703 B.n702 10.6151
R1206 B.n703 B.n334 10.6151
R1207 B.n713 B.n334 10.6151
R1208 B.n714 B.n713 10.6151
R1209 B.n716 B.n714 10.6151
R1210 B.n716 B.n715 10.6151
R1211 B.n715 B.n327 10.6151
R1212 B.n727 B.n327 10.6151
R1213 B.n728 B.n727 10.6151
R1214 B.n729 B.n728 10.6151
R1215 B.n730 B.n729 10.6151
R1216 B.n732 B.n730 10.6151
R1217 B.n733 B.n732 10.6151
R1218 B.n734 B.n733 10.6151
R1219 B.n735 B.n734 10.6151
R1220 B.n737 B.n735 10.6151
R1221 B.n738 B.n737 10.6151
R1222 B.n739 B.n738 10.6151
R1223 B.n740 B.n739 10.6151
R1224 B.n742 B.n740 10.6151
R1225 B.n743 B.n742 10.6151
R1226 B.n744 B.n743 10.6151
R1227 B.n745 B.n744 10.6151
R1228 B.n747 B.n745 10.6151
R1229 B.n748 B.n747 10.6151
R1230 B.n749 B.n748 10.6151
R1231 B.n750 B.n749 10.6151
R1232 B.n752 B.n750 10.6151
R1233 B.n753 B.n752 10.6151
R1234 B.n754 B.n753 10.6151
R1235 B.n755 B.n754 10.6151
R1236 B.n757 B.n755 10.6151
R1237 B.n758 B.n757 10.6151
R1238 B.n432 B.n370 10.6151
R1239 B.n433 B.n432 10.6151
R1240 B.n434 B.n433 10.6151
R1241 B.n434 B.n428 10.6151
R1242 B.n440 B.n428 10.6151
R1243 B.n441 B.n440 10.6151
R1244 B.n442 B.n441 10.6151
R1245 B.n442 B.n426 10.6151
R1246 B.n448 B.n426 10.6151
R1247 B.n449 B.n448 10.6151
R1248 B.n450 B.n449 10.6151
R1249 B.n450 B.n424 10.6151
R1250 B.n456 B.n424 10.6151
R1251 B.n457 B.n456 10.6151
R1252 B.n458 B.n457 10.6151
R1253 B.n458 B.n422 10.6151
R1254 B.n464 B.n422 10.6151
R1255 B.n465 B.n464 10.6151
R1256 B.n466 B.n465 10.6151
R1257 B.n466 B.n420 10.6151
R1258 B.n472 B.n420 10.6151
R1259 B.n473 B.n472 10.6151
R1260 B.n474 B.n473 10.6151
R1261 B.n474 B.n418 10.6151
R1262 B.n480 B.n418 10.6151
R1263 B.n481 B.n480 10.6151
R1264 B.n482 B.n481 10.6151
R1265 B.n482 B.n416 10.6151
R1266 B.n488 B.n416 10.6151
R1267 B.n489 B.n488 10.6151
R1268 B.n490 B.n489 10.6151
R1269 B.n490 B.n414 10.6151
R1270 B.n496 B.n414 10.6151
R1271 B.n497 B.n496 10.6151
R1272 B.n498 B.n497 10.6151
R1273 B.n498 B.n412 10.6151
R1274 B.n504 B.n412 10.6151
R1275 B.n505 B.n504 10.6151
R1276 B.n506 B.n505 10.6151
R1277 B.n506 B.n410 10.6151
R1278 B.n512 B.n410 10.6151
R1279 B.n513 B.n512 10.6151
R1280 B.n514 B.n513 10.6151
R1281 B.n514 B.n408 10.6151
R1282 B.n520 B.n408 10.6151
R1283 B.n521 B.n520 10.6151
R1284 B.n522 B.n521 10.6151
R1285 B.n522 B.n406 10.6151
R1286 B.n528 B.n406 10.6151
R1287 B.n529 B.n528 10.6151
R1288 B.n531 B.n402 10.6151
R1289 B.n537 B.n402 10.6151
R1290 B.n538 B.n537 10.6151
R1291 B.n539 B.n538 10.6151
R1292 B.n539 B.n400 10.6151
R1293 B.n545 B.n400 10.6151
R1294 B.n546 B.n545 10.6151
R1295 B.n550 B.n546 10.6151
R1296 B.n556 B.n398 10.6151
R1297 B.n557 B.n556 10.6151
R1298 B.n558 B.n557 10.6151
R1299 B.n558 B.n396 10.6151
R1300 B.n564 B.n396 10.6151
R1301 B.n565 B.n564 10.6151
R1302 B.n566 B.n565 10.6151
R1303 B.n566 B.n394 10.6151
R1304 B.n572 B.n394 10.6151
R1305 B.n573 B.n572 10.6151
R1306 B.n574 B.n573 10.6151
R1307 B.n574 B.n392 10.6151
R1308 B.n580 B.n392 10.6151
R1309 B.n581 B.n580 10.6151
R1310 B.n582 B.n581 10.6151
R1311 B.n582 B.n390 10.6151
R1312 B.n588 B.n390 10.6151
R1313 B.n589 B.n588 10.6151
R1314 B.n590 B.n589 10.6151
R1315 B.n590 B.n388 10.6151
R1316 B.n596 B.n388 10.6151
R1317 B.n597 B.n596 10.6151
R1318 B.n598 B.n597 10.6151
R1319 B.n598 B.n386 10.6151
R1320 B.n604 B.n386 10.6151
R1321 B.n605 B.n604 10.6151
R1322 B.n606 B.n605 10.6151
R1323 B.n606 B.n384 10.6151
R1324 B.n612 B.n384 10.6151
R1325 B.n613 B.n612 10.6151
R1326 B.n614 B.n613 10.6151
R1327 B.n614 B.n382 10.6151
R1328 B.n620 B.n382 10.6151
R1329 B.n621 B.n620 10.6151
R1330 B.n622 B.n621 10.6151
R1331 B.n622 B.n380 10.6151
R1332 B.n628 B.n380 10.6151
R1333 B.n629 B.n628 10.6151
R1334 B.n630 B.n629 10.6151
R1335 B.n630 B.n378 10.6151
R1336 B.n636 B.n378 10.6151
R1337 B.n637 B.n636 10.6151
R1338 B.n638 B.n637 10.6151
R1339 B.n638 B.n376 10.6151
R1340 B.n644 B.n376 10.6151
R1341 B.n645 B.n644 10.6151
R1342 B.n646 B.n645 10.6151
R1343 B.n646 B.n374 10.6151
R1344 B.n652 B.n374 10.6151
R1345 B.n653 B.n652 10.6151
R1346 B.n659 B.n658 10.6151
R1347 B.n660 B.n659 10.6151
R1348 B.n660 B.n362 10.6151
R1349 B.n671 B.n362 10.6151
R1350 B.n672 B.n671 10.6151
R1351 B.n673 B.n672 10.6151
R1352 B.n673 B.n355 10.6151
R1353 B.n683 B.n355 10.6151
R1354 B.n684 B.n683 10.6151
R1355 B.n685 B.n684 10.6151
R1356 B.n685 B.n347 10.6151
R1357 B.n695 B.n347 10.6151
R1358 B.n696 B.n695 10.6151
R1359 B.n697 B.n696 10.6151
R1360 B.n697 B.n339 10.6151
R1361 B.n707 B.n339 10.6151
R1362 B.n708 B.n707 10.6151
R1363 B.n709 B.n708 10.6151
R1364 B.n709 B.n331 10.6151
R1365 B.n720 B.n331 10.6151
R1366 B.n721 B.n720 10.6151
R1367 B.n722 B.n721 10.6151
R1368 B.n722 B.n0 10.6151
R1369 B.n806 B.n1 10.6151
R1370 B.n806 B.n805 10.6151
R1371 B.n805 B.n804 10.6151
R1372 B.n804 B.n10 10.6151
R1373 B.n798 B.n10 10.6151
R1374 B.n798 B.n797 10.6151
R1375 B.n797 B.n796 10.6151
R1376 B.n796 B.n17 10.6151
R1377 B.n790 B.n17 10.6151
R1378 B.n790 B.n789 10.6151
R1379 B.n789 B.n788 10.6151
R1380 B.n788 B.n24 10.6151
R1381 B.n782 B.n24 10.6151
R1382 B.n782 B.n781 10.6151
R1383 B.n781 B.n780 10.6151
R1384 B.n780 B.n31 10.6151
R1385 B.n774 B.n31 10.6151
R1386 B.n774 B.n773 10.6151
R1387 B.n773 B.n772 10.6151
R1388 B.n772 B.n37 10.6151
R1389 B.n766 B.n37 10.6151
R1390 B.n766 B.n765 10.6151
R1391 B.n765 B.n764 10.6151
R1392 B.n718 B.t3 9.21459
R1393 B.n802 B.t2 9.21459
R1394 B.n210 B.n209 6.5566
R1395 B.n226 B.n106 6.5566
R1396 B.n531 B.n530 6.5566
R1397 B.n550 B.n549 6.5566
R1398 B.n209 B.n208 4.05904
R1399 B.n229 B.n106 4.05904
R1400 B.n530 B.n529 4.05904
R1401 B.n549 B.n398 4.05904
R1402 B.n812 B.n0 2.81026
R1403 B.n812 B.n1 2.81026
R1404 B.n675 B.t5 1.62652
R1405 B.n776 B.t9 1.62652
R1406 VN.n0 VN.t1 282.248
R1407 VN.n1 VN.t2 282.248
R1408 VN.n0 VN.t3 281.933
R1409 VN.n1 VN.t0 281.933
R1410 VN VN.n1 58.5245
R1411 VN VN.n0 13.1495
R1412 VDD2.n2 VDD2.n0 102.585
R1413 VDD2.n2 VDD2.n1 61.2675
R1414 VDD2.n1 VDD2.t3 1.31874
R1415 VDD2.n1 VDD2.t1 1.31874
R1416 VDD2.n0 VDD2.t2 1.31874
R1417 VDD2.n0 VDD2.t0 1.31874
R1418 VDD2 VDD2.n2 0.0586897
C0 VP VN 5.93481f
C1 VDD1 VDD2 0.752352f
C2 VDD1 VN 0.148429f
C3 VP VTAIL 4.76263f
C4 VDD2 VN 5.13046f
C5 VDD1 VTAIL 6.46911f
C6 VDD1 VP 5.30443f
C7 VTAIL VDD2 6.51574f
C8 VTAIL VN 4.74852f
C9 VP VDD2 0.322852f
C10 VDD2 B 3.369412f
C11 VDD1 B 7.46927f
C12 VTAIL B 11.161695f
C13 VN B 9.089221f
C14 VP B 6.729236f
C15 VDD2.t2 B 0.315395f
C16 VDD2.t0 B 0.315395f
C17 VDD2.n0 B 3.56873f
C18 VDD2.t3 B 0.315395f
C19 VDD2.t1 B 0.315395f
C20 VDD2.n1 B 2.85145f
C21 VDD2.n2 B 3.77966f
C22 VN.t1 B 2.2133f
C23 VN.t3 B 2.21229f
C24 VN.n0 B 1.59116f
C25 VN.t2 B 2.2133f
C26 VN.t0 B 2.21229f
C27 VN.n1 B 3.00182f
C28 VTAIL.t7 B 2.05242f
C29 VTAIL.n0 B 0.271161f
C30 VTAIL.t3 B 2.05242f
C31 VTAIL.n1 B 0.306817f
C32 VTAIL.t5 B 2.05242f
C33 VTAIL.n2 B 1.21334f
C34 VTAIL.t1 B 2.05242f
C35 VTAIL.n3 B 1.21334f
C36 VTAIL.t6 B 2.05242f
C37 VTAIL.n4 B 0.306815f
C38 VTAIL.t2 B 2.05242f
C39 VTAIL.n5 B 0.306815f
C40 VTAIL.t4 B 2.05242f
C41 VTAIL.n6 B 1.21334f
C42 VTAIL.t0 B 2.05242f
C43 VTAIL.n7 B 1.1719f
C44 VDD1.t2 B 0.318141f
C45 VDD1.t3 B 0.318141f
C46 VDD1.n0 B 2.87663f
C47 VDD1.t1 B 0.318141f
C48 VDD1.t0 B 0.318141f
C49 VDD1.n1 B 3.627f
C50 VP.n0 B 0.035492f
C51 VP.t2 B 2.14741f
C52 VP.n1 B 0.051593f
C53 VP.t3 B 2.26263f
C54 VP.t1 B 2.2616f
C55 VP.n2 B 3.04802f
C56 VP.n3 B 2.09102f
C57 VP.t0 B 2.14741f
C58 VP.n4 B 0.831058f
C59 VP.n5 B 0.043073f
C60 VP.n6 B 0.035492f
C61 VP.n7 B 0.035492f
C62 VP.n8 B 0.035492f
C63 VP.n9 B 0.051593f
C64 VP.n10 B 0.043073f
C65 VP.n11 B 0.831058f
C66 VP.n12 B 0.034604f
.ends

