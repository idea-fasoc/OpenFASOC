* NGSPICE file created from diff_pair_sample_0936.ext - technology: sky130A

.subckt diff_pair_sample_0936 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2212_n3270# sky130_fd_pr__pfet_01v8 ad=4.4889 pd=23.8 as=0 ps=0 w=11.51 l=1.74
X1 VDD1.t3 VP.t0 VTAIL.t6 w_n2212_n3270# sky130_fd_pr__pfet_01v8 ad=1.89915 pd=11.84 as=4.4889 ps=23.8 w=11.51 l=1.74
X2 VTAIL.t3 VN.t0 VDD2.t3 w_n2212_n3270# sky130_fd_pr__pfet_01v8 ad=4.4889 pd=23.8 as=1.89915 ps=11.84 w=11.51 l=1.74
X3 VDD2.t2 VN.t1 VTAIL.t2 w_n2212_n3270# sky130_fd_pr__pfet_01v8 ad=1.89915 pd=11.84 as=4.4889 ps=23.8 w=11.51 l=1.74
X4 B.t8 B.t6 B.t7 w_n2212_n3270# sky130_fd_pr__pfet_01v8 ad=4.4889 pd=23.8 as=0 ps=0 w=11.51 l=1.74
X5 VDD2.t1 VN.t2 VTAIL.t1 w_n2212_n3270# sky130_fd_pr__pfet_01v8 ad=1.89915 pd=11.84 as=4.4889 ps=23.8 w=11.51 l=1.74
X6 VDD1.t2 VP.t1 VTAIL.t5 w_n2212_n3270# sky130_fd_pr__pfet_01v8 ad=1.89915 pd=11.84 as=4.4889 ps=23.8 w=11.51 l=1.74
X7 VTAIL.t0 VN.t3 VDD2.t0 w_n2212_n3270# sky130_fd_pr__pfet_01v8 ad=4.4889 pd=23.8 as=1.89915 ps=11.84 w=11.51 l=1.74
X8 B.t5 B.t3 B.t4 w_n2212_n3270# sky130_fd_pr__pfet_01v8 ad=4.4889 pd=23.8 as=0 ps=0 w=11.51 l=1.74
X9 B.t2 B.t0 B.t1 w_n2212_n3270# sky130_fd_pr__pfet_01v8 ad=4.4889 pd=23.8 as=0 ps=0 w=11.51 l=1.74
X10 VTAIL.t4 VP.t2 VDD1.t1 w_n2212_n3270# sky130_fd_pr__pfet_01v8 ad=4.4889 pd=23.8 as=1.89915 ps=11.84 w=11.51 l=1.74
X11 VTAIL.t7 VP.t3 VDD1.t0 w_n2212_n3270# sky130_fd_pr__pfet_01v8 ad=4.4889 pd=23.8 as=1.89915 ps=11.84 w=11.51 l=1.74
R0 B.n327 B.n326 585
R1 B.n325 B.n92 585
R2 B.n324 B.n323 585
R3 B.n322 B.n93 585
R4 B.n321 B.n320 585
R5 B.n319 B.n94 585
R6 B.n318 B.n317 585
R7 B.n316 B.n95 585
R8 B.n315 B.n314 585
R9 B.n313 B.n96 585
R10 B.n312 B.n311 585
R11 B.n310 B.n97 585
R12 B.n309 B.n308 585
R13 B.n307 B.n98 585
R14 B.n306 B.n305 585
R15 B.n304 B.n99 585
R16 B.n303 B.n302 585
R17 B.n301 B.n100 585
R18 B.n300 B.n299 585
R19 B.n298 B.n101 585
R20 B.n297 B.n296 585
R21 B.n295 B.n102 585
R22 B.n294 B.n293 585
R23 B.n292 B.n103 585
R24 B.n291 B.n290 585
R25 B.n289 B.n104 585
R26 B.n288 B.n287 585
R27 B.n286 B.n105 585
R28 B.n285 B.n284 585
R29 B.n283 B.n106 585
R30 B.n282 B.n281 585
R31 B.n280 B.n107 585
R32 B.n279 B.n278 585
R33 B.n277 B.n108 585
R34 B.n276 B.n275 585
R35 B.n274 B.n109 585
R36 B.n273 B.n272 585
R37 B.n271 B.n110 585
R38 B.n270 B.n269 585
R39 B.n268 B.n111 585
R40 B.n266 B.n265 585
R41 B.n264 B.n114 585
R42 B.n263 B.n262 585
R43 B.n261 B.n115 585
R44 B.n260 B.n259 585
R45 B.n258 B.n116 585
R46 B.n257 B.n256 585
R47 B.n255 B.n117 585
R48 B.n254 B.n253 585
R49 B.n252 B.n118 585
R50 B.n251 B.n250 585
R51 B.n246 B.n119 585
R52 B.n245 B.n244 585
R53 B.n243 B.n120 585
R54 B.n242 B.n241 585
R55 B.n240 B.n121 585
R56 B.n239 B.n238 585
R57 B.n237 B.n122 585
R58 B.n236 B.n235 585
R59 B.n234 B.n123 585
R60 B.n233 B.n232 585
R61 B.n231 B.n124 585
R62 B.n230 B.n229 585
R63 B.n228 B.n125 585
R64 B.n227 B.n226 585
R65 B.n225 B.n126 585
R66 B.n224 B.n223 585
R67 B.n222 B.n127 585
R68 B.n221 B.n220 585
R69 B.n219 B.n128 585
R70 B.n218 B.n217 585
R71 B.n216 B.n129 585
R72 B.n215 B.n214 585
R73 B.n213 B.n130 585
R74 B.n212 B.n211 585
R75 B.n210 B.n131 585
R76 B.n209 B.n208 585
R77 B.n207 B.n132 585
R78 B.n206 B.n205 585
R79 B.n204 B.n133 585
R80 B.n203 B.n202 585
R81 B.n201 B.n134 585
R82 B.n200 B.n199 585
R83 B.n198 B.n135 585
R84 B.n197 B.n196 585
R85 B.n195 B.n136 585
R86 B.n194 B.n193 585
R87 B.n192 B.n137 585
R88 B.n191 B.n190 585
R89 B.n189 B.n138 585
R90 B.n328 B.n91 585
R91 B.n330 B.n329 585
R92 B.n331 B.n90 585
R93 B.n333 B.n332 585
R94 B.n334 B.n89 585
R95 B.n336 B.n335 585
R96 B.n337 B.n88 585
R97 B.n339 B.n338 585
R98 B.n340 B.n87 585
R99 B.n342 B.n341 585
R100 B.n343 B.n86 585
R101 B.n345 B.n344 585
R102 B.n346 B.n85 585
R103 B.n348 B.n347 585
R104 B.n349 B.n84 585
R105 B.n351 B.n350 585
R106 B.n352 B.n83 585
R107 B.n354 B.n353 585
R108 B.n355 B.n82 585
R109 B.n357 B.n356 585
R110 B.n358 B.n81 585
R111 B.n360 B.n359 585
R112 B.n361 B.n80 585
R113 B.n363 B.n362 585
R114 B.n364 B.n79 585
R115 B.n366 B.n365 585
R116 B.n367 B.n78 585
R117 B.n369 B.n368 585
R118 B.n370 B.n77 585
R119 B.n372 B.n371 585
R120 B.n373 B.n76 585
R121 B.n375 B.n374 585
R122 B.n376 B.n75 585
R123 B.n378 B.n377 585
R124 B.n379 B.n74 585
R125 B.n381 B.n380 585
R126 B.n382 B.n73 585
R127 B.n384 B.n383 585
R128 B.n385 B.n72 585
R129 B.n387 B.n386 585
R130 B.n388 B.n71 585
R131 B.n390 B.n389 585
R132 B.n391 B.n70 585
R133 B.n393 B.n392 585
R134 B.n394 B.n69 585
R135 B.n396 B.n395 585
R136 B.n397 B.n68 585
R137 B.n399 B.n398 585
R138 B.n400 B.n67 585
R139 B.n402 B.n401 585
R140 B.n403 B.n66 585
R141 B.n405 B.n404 585
R142 B.n406 B.n65 585
R143 B.n408 B.n407 585
R144 B.n544 B.n15 585
R145 B.n543 B.n542 585
R146 B.n541 B.n16 585
R147 B.n540 B.n539 585
R148 B.n538 B.n17 585
R149 B.n537 B.n536 585
R150 B.n535 B.n18 585
R151 B.n534 B.n533 585
R152 B.n532 B.n19 585
R153 B.n531 B.n530 585
R154 B.n529 B.n20 585
R155 B.n528 B.n527 585
R156 B.n526 B.n21 585
R157 B.n525 B.n524 585
R158 B.n523 B.n22 585
R159 B.n522 B.n521 585
R160 B.n520 B.n23 585
R161 B.n519 B.n518 585
R162 B.n517 B.n24 585
R163 B.n516 B.n515 585
R164 B.n514 B.n25 585
R165 B.n513 B.n512 585
R166 B.n511 B.n26 585
R167 B.n510 B.n509 585
R168 B.n508 B.n27 585
R169 B.n507 B.n506 585
R170 B.n505 B.n28 585
R171 B.n504 B.n503 585
R172 B.n502 B.n29 585
R173 B.n501 B.n500 585
R174 B.n499 B.n30 585
R175 B.n498 B.n497 585
R176 B.n496 B.n31 585
R177 B.n495 B.n494 585
R178 B.n493 B.n32 585
R179 B.n492 B.n491 585
R180 B.n490 B.n33 585
R181 B.n489 B.n488 585
R182 B.n487 B.n34 585
R183 B.n486 B.n485 585
R184 B.n483 B.n35 585
R185 B.n482 B.n481 585
R186 B.n480 B.n38 585
R187 B.n479 B.n478 585
R188 B.n477 B.n39 585
R189 B.n476 B.n475 585
R190 B.n474 B.n40 585
R191 B.n473 B.n472 585
R192 B.n471 B.n41 585
R193 B.n470 B.n469 585
R194 B.n468 B.n467 585
R195 B.n466 B.n45 585
R196 B.n465 B.n464 585
R197 B.n463 B.n46 585
R198 B.n462 B.n461 585
R199 B.n460 B.n47 585
R200 B.n459 B.n458 585
R201 B.n457 B.n48 585
R202 B.n456 B.n455 585
R203 B.n454 B.n49 585
R204 B.n453 B.n452 585
R205 B.n451 B.n50 585
R206 B.n450 B.n449 585
R207 B.n448 B.n51 585
R208 B.n447 B.n446 585
R209 B.n445 B.n52 585
R210 B.n444 B.n443 585
R211 B.n442 B.n53 585
R212 B.n441 B.n440 585
R213 B.n439 B.n54 585
R214 B.n438 B.n437 585
R215 B.n436 B.n55 585
R216 B.n435 B.n434 585
R217 B.n433 B.n56 585
R218 B.n432 B.n431 585
R219 B.n430 B.n57 585
R220 B.n429 B.n428 585
R221 B.n427 B.n58 585
R222 B.n426 B.n425 585
R223 B.n424 B.n59 585
R224 B.n423 B.n422 585
R225 B.n421 B.n60 585
R226 B.n420 B.n419 585
R227 B.n418 B.n61 585
R228 B.n417 B.n416 585
R229 B.n415 B.n62 585
R230 B.n414 B.n413 585
R231 B.n412 B.n63 585
R232 B.n411 B.n410 585
R233 B.n409 B.n64 585
R234 B.n546 B.n545 585
R235 B.n547 B.n14 585
R236 B.n549 B.n548 585
R237 B.n550 B.n13 585
R238 B.n552 B.n551 585
R239 B.n553 B.n12 585
R240 B.n555 B.n554 585
R241 B.n556 B.n11 585
R242 B.n558 B.n557 585
R243 B.n559 B.n10 585
R244 B.n561 B.n560 585
R245 B.n562 B.n9 585
R246 B.n564 B.n563 585
R247 B.n565 B.n8 585
R248 B.n567 B.n566 585
R249 B.n568 B.n7 585
R250 B.n570 B.n569 585
R251 B.n571 B.n6 585
R252 B.n573 B.n572 585
R253 B.n574 B.n5 585
R254 B.n576 B.n575 585
R255 B.n577 B.n4 585
R256 B.n579 B.n578 585
R257 B.n580 B.n3 585
R258 B.n582 B.n581 585
R259 B.n583 B.n0 585
R260 B.n2 B.n1 585
R261 B.n152 B.n151 585
R262 B.n153 B.n150 585
R263 B.n155 B.n154 585
R264 B.n156 B.n149 585
R265 B.n158 B.n157 585
R266 B.n159 B.n148 585
R267 B.n161 B.n160 585
R268 B.n162 B.n147 585
R269 B.n164 B.n163 585
R270 B.n165 B.n146 585
R271 B.n167 B.n166 585
R272 B.n168 B.n145 585
R273 B.n170 B.n169 585
R274 B.n171 B.n144 585
R275 B.n173 B.n172 585
R276 B.n174 B.n143 585
R277 B.n176 B.n175 585
R278 B.n177 B.n142 585
R279 B.n179 B.n178 585
R280 B.n180 B.n141 585
R281 B.n182 B.n181 585
R282 B.n183 B.n140 585
R283 B.n185 B.n184 585
R284 B.n186 B.n139 585
R285 B.n188 B.n187 585
R286 B.n189 B.n188 473.281
R287 B.n326 B.n91 473.281
R288 B.n409 B.n408 473.281
R289 B.n546 B.n15 473.281
R290 B.n112 B.t4 407.115
R291 B.n42 B.t2 407.115
R292 B.n247 B.t10 407.115
R293 B.n36 B.t8 407.115
R294 B.n113 B.t5 366.969
R295 B.n43 B.t1 366.969
R296 B.n248 B.t11 366.969
R297 B.n37 B.t7 366.969
R298 B.n247 B.t9 365.654
R299 B.n112 B.t3 365.654
R300 B.n42 B.t0 365.654
R301 B.n36 B.t6 365.654
R302 B.n585 B.n584 256.663
R303 B.n584 B.n583 235.042
R304 B.n584 B.n2 235.042
R305 B.n190 B.n189 163.367
R306 B.n190 B.n137 163.367
R307 B.n194 B.n137 163.367
R308 B.n195 B.n194 163.367
R309 B.n196 B.n195 163.367
R310 B.n196 B.n135 163.367
R311 B.n200 B.n135 163.367
R312 B.n201 B.n200 163.367
R313 B.n202 B.n201 163.367
R314 B.n202 B.n133 163.367
R315 B.n206 B.n133 163.367
R316 B.n207 B.n206 163.367
R317 B.n208 B.n207 163.367
R318 B.n208 B.n131 163.367
R319 B.n212 B.n131 163.367
R320 B.n213 B.n212 163.367
R321 B.n214 B.n213 163.367
R322 B.n214 B.n129 163.367
R323 B.n218 B.n129 163.367
R324 B.n219 B.n218 163.367
R325 B.n220 B.n219 163.367
R326 B.n220 B.n127 163.367
R327 B.n224 B.n127 163.367
R328 B.n225 B.n224 163.367
R329 B.n226 B.n225 163.367
R330 B.n226 B.n125 163.367
R331 B.n230 B.n125 163.367
R332 B.n231 B.n230 163.367
R333 B.n232 B.n231 163.367
R334 B.n232 B.n123 163.367
R335 B.n236 B.n123 163.367
R336 B.n237 B.n236 163.367
R337 B.n238 B.n237 163.367
R338 B.n238 B.n121 163.367
R339 B.n242 B.n121 163.367
R340 B.n243 B.n242 163.367
R341 B.n244 B.n243 163.367
R342 B.n244 B.n119 163.367
R343 B.n251 B.n119 163.367
R344 B.n252 B.n251 163.367
R345 B.n253 B.n252 163.367
R346 B.n253 B.n117 163.367
R347 B.n257 B.n117 163.367
R348 B.n258 B.n257 163.367
R349 B.n259 B.n258 163.367
R350 B.n259 B.n115 163.367
R351 B.n263 B.n115 163.367
R352 B.n264 B.n263 163.367
R353 B.n265 B.n264 163.367
R354 B.n265 B.n111 163.367
R355 B.n270 B.n111 163.367
R356 B.n271 B.n270 163.367
R357 B.n272 B.n271 163.367
R358 B.n272 B.n109 163.367
R359 B.n276 B.n109 163.367
R360 B.n277 B.n276 163.367
R361 B.n278 B.n277 163.367
R362 B.n278 B.n107 163.367
R363 B.n282 B.n107 163.367
R364 B.n283 B.n282 163.367
R365 B.n284 B.n283 163.367
R366 B.n284 B.n105 163.367
R367 B.n288 B.n105 163.367
R368 B.n289 B.n288 163.367
R369 B.n290 B.n289 163.367
R370 B.n290 B.n103 163.367
R371 B.n294 B.n103 163.367
R372 B.n295 B.n294 163.367
R373 B.n296 B.n295 163.367
R374 B.n296 B.n101 163.367
R375 B.n300 B.n101 163.367
R376 B.n301 B.n300 163.367
R377 B.n302 B.n301 163.367
R378 B.n302 B.n99 163.367
R379 B.n306 B.n99 163.367
R380 B.n307 B.n306 163.367
R381 B.n308 B.n307 163.367
R382 B.n308 B.n97 163.367
R383 B.n312 B.n97 163.367
R384 B.n313 B.n312 163.367
R385 B.n314 B.n313 163.367
R386 B.n314 B.n95 163.367
R387 B.n318 B.n95 163.367
R388 B.n319 B.n318 163.367
R389 B.n320 B.n319 163.367
R390 B.n320 B.n93 163.367
R391 B.n324 B.n93 163.367
R392 B.n325 B.n324 163.367
R393 B.n326 B.n325 163.367
R394 B.n408 B.n65 163.367
R395 B.n404 B.n65 163.367
R396 B.n404 B.n403 163.367
R397 B.n403 B.n402 163.367
R398 B.n402 B.n67 163.367
R399 B.n398 B.n67 163.367
R400 B.n398 B.n397 163.367
R401 B.n397 B.n396 163.367
R402 B.n396 B.n69 163.367
R403 B.n392 B.n69 163.367
R404 B.n392 B.n391 163.367
R405 B.n391 B.n390 163.367
R406 B.n390 B.n71 163.367
R407 B.n386 B.n71 163.367
R408 B.n386 B.n385 163.367
R409 B.n385 B.n384 163.367
R410 B.n384 B.n73 163.367
R411 B.n380 B.n73 163.367
R412 B.n380 B.n379 163.367
R413 B.n379 B.n378 163.367
R414 B.n378 B.n75 163.367
R415 B.n374 B.n75 163.367
R416 B.n374 B.n373 163.367
R417 B.n373 B.n372 163.367
R418 B.n372 B.n77 163.367
R419 B.n368 B.n77 163.367
R420 B.n368 B.n367 163.367
R421 B.n367 B.n366 163.367
R422 B.n366 B.n79 163.367
R423 B.n362 B.n79 163.367
R424 B.n362 B.n361 163.367
R425 B.n361 B.n360 163.367
R426 B.n360 B.n81 163.367
R427 B.n356 B.n81 163.367
R428 B.n356 B.n355 163.367
R429 B.n355 B.n354 163.367
R430 B.n354 B.n83 163.367
R431 B.n350 B.n83 163.367
R432 B.n350 B.n349 163.367
R433 B.n349 B.n348 163.367
R434 B.n348 B.n85 163.367
R435 B.n344 B.n85 163.367
R436 B.n344 B.n343 163.367
R437 B.n343 B.n342 163.367
R438 B.n342 B.n87 163.367
R439 B.n338 B.n87 163.367
R440 B.n338 B.n337 163.367
R441 B.n337 B.n336 163.367
R442 B.n336 B.n89 163.367
R443 B.n332 B.n89 163.367
R444 B.n332 B.n331 163.367
R445 B.n331 B.n330 163.367
R446 B.n330 B.n91 163.367
R447 B.n542 B.n15 163.367
R448 B.n542 B.n541 163.367
R449 B.n541 B.n540 163.367
R450 B.n540 B.n17 163.367
R451 B.n536 B.n17 163.367
R452 B.n536 B.n535 163.367
R453 B.n535 B.n534 163.367
R454 B.n534 B.n19 163.367
R455 B.n530 B.n19 163.367
R456 B.n530 B.n529 163.367
R457 B.n529 B.n528 163.367
R458 B.n528 B.n21 163.367
R459 B.n524 B.n21 163.367
R460 B.n524 B.n523 163.367
R461 B.n523 B.n522 163.367
R462 B.n522 B.n23 163.367
R463 B.n518 B.n23 163.367
R464 B.n518 B.n517 163.367
R465 B.n517 B.n516 163.367
R466 B.n516 B.n25 163.367
R467 B.n512 B.n25 163.367
R468 B.n512 B.n511 163.367
R469 B.n511 B.n510 163.367
R470 B.n510 B.n27 163.367
R471 B.n506 B.n27 163.367
R472 B.n506 B.n505 163.367
R473 B.n505 B.n504 163.367
R474 B.n504 B.n29 163.367
R475 B.n500 B.n29 163.367
R476 B.n500 B.n499 163.367
R477 B.n499 B.n498 163.367
R478 B.n498 B.n31 163.367
R479 B.n494 B.n31 163.367
R480 B.n494 B.n493 163.367
R481 B.n493 B.n492 163.367
R482 B.n492 B.n33 163.367
R483 B.n488 B.n33 163.367
R484 B.n488 B.n487 163.367
R485 B.n487 B.n486 163.367
R486 B.n486 B.n35 163.367
R487 B.n481 B.n35 163.367
R488 B.n481 B.n480 163.367
R489 B.n480 B.n479 163.367
R490 B.n479 B.n39 163.367
R491 B.n475 B.n39 163.367
R492 B.n475 B.n474 163.367
R493 B.n474 B.n473 163.367
R494 B.n473 B.n41 163.367
R495 B.n469 B.n41 163.367
R496 B.n469 B.n468 163.367
R497 B.n468 B.n45 163.367
R498 B.n464 B.n45 163.367
R499 B.n464 B.n463 163.367
R500 B.n463 B.n462 163.367
R501 B.n462 B.n47 163.367
R502 B.n458 B.n47 163.367
R503 B.n458 B.n457 163.367
R504 B.n457 B.n456 163.367
R505 B.n456 B.n49 163.367
R506 B.n452 B.n49 163.367
R507 B.n452 B.n451 163.367
R508 B.n451 B.n450 163.367
R509 B.n450 B.n51 163.367
R510 B.n446 B.n51 163.367
R511 B.n446 B.n445 163.367
R512 B.n445 B.n444 163.367
R513 B.n444 B.n53 163.367
R514 B.n440 B.n53 163.367
R515 B.n440 B.n439 163.367
R516 B.n439 B.n438 163.367
R517 B.n438 B.n55 163.367
R518 B.n434 B.n55 163.367
R519 B.n434 B.n433 163.367
R520 B.n433 B.n432 163.367
R521 B.n432 B.n57 163.367
R522 B.n428 B.n57 163.367
R523 B.n428 B.n427 163.367
R524 B.n427 B.n426 163.367
R525 B.n426 B.n59 163.367
R526 B.n422 B.n59 163.367
R527 B.n422 B.n421 163.367
R528 B.n421 B.n420 163.367
R529 B.n420 B.n61 163.367
R530 B.n416 B.n61 163.367
R531 B.n416 B.n415 163.367
R532 B.n415 B.n414 163.367
R533 B.n414 B.n63 163.367
R534 B.n410 B.n63 163.367
R535 B.n410 B.n409 163.367
R536 B.n547 B.n546 163.367
R537 B.n548 B.n547 163.367
R538 B.n548 B.n13 163.367
R539 B.n552 B.n13 163.367
R540 B.n553 B.n552 163.367
R541 B.n554 B.n553 163.367
R542 B.n554 B.n11 163.367
R543 B.n558 B.n11 163.367
R544 B.n559 B.n558 163.367
R545 B.n560 B.n559 163.367
R546 B.n560 B.n9 163.367
R547 B.n564 B.n9 163.367
R548 B.n565 B.n564 163.367
R549 B.n566 B.n565 163.367
R550 B.n566 B.n7 163.367
R551 B.n570 B.n7 163.367
R552 B.n571 B.n570 163.367
R553 B.n572 B.n571 163.367
R554 B.n572 B.n5 163.367
R555 B.n576 B.n5 163.367
R556 B.n577 B.n576 163.367
R557 B.n578 B.n577 163.367
R558 B.n578 B.n3 163.367
R559 B.n582 B.n3 163.367
R560 B.n583 B.n582 163.367
R561 B.n152 B.n2 163.367
R562 B.n153 B.n152 163.367
R563 B.n154 B.n153 163.367
R564 B.n154 B.n149 163.367
R565 B.n158 B.n149 163.367
R566 B.n159 B.n158 163.367
R567 B.n160 B.n159 163.367
R568 B.n160 B.n147 163.367
R569 B.n164 B.n147 163.367
R570 B.n165 B.n164 163.367
R571 B.n166 B.n165 163.367
R572 B.n166 B.n145 163.367
R573 B.n170 B.n145 163.367
R574 B.n171 B.n170 163.367
R575 B.n172 B.n171 163.367
R576 B.n172 B.n143 163.367
R577 B.n176 B.n143 163.367
R578 B.n177 B.n176 163.367
R579 B.n178 B.n177 163.367
R580 B.n178 B.n141 163.367
R581 B.n182 B.n141 163.367
R582 B.n183 B.n182 163.367
R583 B.n184 B.n183 163.367
R584 B.n184 B.n139 163.367
R585 B.n188 B.n139 163.367
R586 B.n249 B.n248 59.5399
R587 B.n267 B.n113 59.5399
R588 B.n44 B.n43 59.5399
R589 B.n484 B.n37 59.5399
R590 B.n248 B.n247 40.146
R591 B.n113 B.n112 40.146
R592 B.n43 B.n42 40.146
R593 B.n37 B.n36 40.146
R594 B.n545 B.n544 30.7517
R595 B.n407 B.n64 30.7517
R596 B.n328 B.n327 30.7517
R597 B.n187 B.n138 30.7517
R598 B B.n585 18.0485
R599 B.n545 B.n14 10.6151
R600 B.n549 B.n14 10.6151
R601 B.n550 B.n549 10.6151
R602 B.n551 B.n550 10.6151
R603 B.n551 B.n12 10.6151
R604 B.n555 B.n12 10.6151
R605 B.n556 B.n555 10.6151
R606 B.n557 B.n556 10.6151
R607 B.n557 B.n10 10.6151
R608 B.n561 B.n10 10.6151
R609 B.n562 B.n561 10.6151
R610 B.n563 B.n562 10.6151
R611 B.n563 B.n8 10.6151
R612 B.n567 B.n8 10.6151
R613 B.n568 B.n567 10.6151
R614 B.n569 B.n568 10.6151
R615 B.n569 B.n6 10.6151
R616 B.n573 B.n6 10.6151
R617 B.n574 B.n573 10.6151
R618 B.n575 B.n574 10.6151
R619 B.n575 B.n4 10.6151
R620 B.n579 B.n4 10.6151
R621 B.n580 B.n579 10.6151
R622 B.n581 B.n580 10.6151
R623 B.n581 B.n0 10.6151
R624 B.n544 B.n543 10.6151
R625 B.n543 B.n16 10.6151
R626 B.n539 B.n16 10.6151
R627 B.n539 B.n538 10.6151
R628 B.n538 B.n537 10.6151
R629 B.n537 B.n18 10.6151
R630 B.n533 B.n18 10.6151
R631 B.n533 B.n532 10.6151
R632 B.n532 B.n531 10.6151
R633 B.n531 B.n20 10.6151
R634 B.n527 B.n20 10.6151
R635 B.n527 B.n526 10.6151
R636 B.n526 B.n525 10.6151
R637 B.n525 B.n22 10.6151
R638 B.n521 B.n22 10.6151
R639 B.n521 B.n520 10.6151
R640 B.n520 B.n519 10.6151
R641 B.n519 B.n24 10.6151
R642 B.n515 B.n24 10.6151
R643 B.n515 B.n514 10.6151
R644 B.n514 B.n513 10.6151
R645 B.n513 B.n26 10.6151
R646 B.n509 B.n26 10.6151
R647 B.n509 B.n508 10.6151
R648 B.n508 B.n507 10.6151
R649 B.n507 B.n28 10.6151
R650 B.n503 B.n28 10.6151
R651 B.n503 B.n502 10.6151
R652 B.n502 B.n501 10.6151
R653 B.n501 B.n30 10.6151
R654 B.n497 B.n30 10.6151
R655 B.n497 B.n496 10.6151
R656 B.n496 B.n495 10.6151
R657 B.n495 B.n32 10.6151
R658 B.n491 B.n32 10.6151
R659 B.n491 B.n490 10.6151
R660 B.n490 B.n489 10.6151
R661 B.n489 B.n34 10.6151
R662 B.n485 B.n34 10.6151
R663 B.n483 B.n482 10.6151
R664 B.n482 B.n38 10.6151
R665 B.n478 B.n38 10.6151
R666 B.n478 B.n477 10.6151
R667 B.n477 B.n476 10.6151
R668 B.n476 B.n40 10.6151
R669 B.n472 B.n40 10.6151
R670 B.n472 B.n471 10.6151
R671 B.n471 B.n470 10.6151
R672 B.n467 B.n466 10.6151
R673 B.n466 B.n465 10.6151
R674 B.n465 B.n46 10.6151
R675 B.n461 B.n46 10.6151
R676 B.n461 B.n460 10.6151
R677 B.n460 B.n459 10.6151
R678 B.n459 B.n48 10.6151
R679 B.n455 B.n48 10.6151
R680 B.n455 B.n454 10.6151
R681 B.n454 B.n453 10.6151
R682 B.n453 B.n50 10.6151
R683 B.n449 B.n50 10.6151
R684 B.n449 B.n448 10.6151
R685 B.n448 B.n447 10.6151
R686 B.n447 B.n52 10.6151
R687 B.n443 B.n52 10.6151
R688 B.n443 B.n442 10.6151
R689 B.n442 B.n441 10.6151
R690 B.n441 B.n54 10.6151
R691 B.n437 B.n54 10.6151
R692 B.n437 B.n436 10.6151
R693 B.n436 B.n435 10.6151
R694 B.n435 B.n56 10.6151
R695 B.n431 B.n56 10.6151
R696 B.n431 B.n430 10.6151
R697 B.n430 B.n429 10.6151
R698 B.n429 B.n58 10.6151
R699 B.n425 B.n58 10.6151
R700 B.n425 B.n424 10.6151
R701 B.n424 B.n423 10.6151
R702 B.n423 B.n60 10.6151
R703 B.n419 B.n60 10.6151
R704 B.n419 B.n418 10.6151
R705 B.n418 B.n417 10.6151
R706 B.n417 B.n62 10.6151
R707 B.n413 B.n62 10.6151
R708 B.n413 B.n412 10.6151
R709 B.n412 B.n411 10.6151
R710 B.n411 B.n64 10.6151
R711 B.n407 B.n406 10.6151
R712 B.n406 B.n405 10.6151
R713 B.n405 B.n66 10.6151
R714 B.n401 B.n66 10.6151
R715 B.n401 B.n400 10.6151
R716 B.n400 B.n399 10.6151
R717 B.n399 B.n68 10.6151
R718 B.n395 B.n68 10.6151
R719 B.n395 B.n394 10.6151
R720 B.n394 B.n393 10.6151
R721 B.n393 B.n70 10.6151
R722 B.n389 B.n70 10.6151
R723 B.n389 B.n388 10.6151
R724 B.n388 B.n387 10.6151
R725 B.n387 B.n72 10.6151
R726 B.n383 B.n72 10.6151
R727 B.n383 B.n382 10.6151
R728 B.n382 B.n381 10.6151
R729 B.n381 B.n74 10.6151
R730 B.n377 B.n74 10.6151
R731 B.n377 B.n376 10.6151
R732 B.n376 B.n375 10.6151
R733 B.n375 B.n76 10.6151
R734 B.n371 B.n76 10.6151
R735 B.n371 B.n370 10.6151
R736 B.n370 B.n369 10.6151
R737 B.n369 B.n78 10.6151
R738 B.n365 B.n78 10.6151
R739 B.n365 B.n364 10.6151
R740 B.n364 B.n363 10.6151
R741 B.n363 B.n80 10.6151
R742 B.n359 B.n80 10.6151
R743 B.n359 B.n358 10.6151
R744 B.n358 B.n357 10.6151
R745 B.n357 B.n82 10.6151
R746 B.n353 B.n82 10.6151
R747 B.n353 B.n352 10.6151
R748 B.n352 B.n351 10.6151
R749 B.n351 B.n84 10.6151
R750 B.n347 B.n84 10.6151
R751 B.n347 B.n346 10.6151
R752 B.n346 B.n345 10.6151
R753 B.n345 B.n86 10.6151
R754 B.n341 B.n86 10.6151
R755 B.n341 B.n340 10.6151
R756 B.n340 B.n339 10.6151
R757 B.n339 B.n88 10.6151
R758 B.n335 B.n88 10.6151
R759 B.n335 B.n334 10.6151
R760 B.n334 B.n333 10.6151
R761 B.n333 B.n90 10.6151
R762 B.n329 B.n90 10.6151
R763 B.n329 B.n328 10.6151
R764 B.n151 B.n1 10.6151
R765 B.n151 B.n150 10.6151
R766 B.n155 B.n150 10.6151
R767 B.n156 B.n155 10.6151
R768 B.n157 B.n156 10.6151
R769 B.n157 B.n148 10.6151
R770 B.n161 B.n148 10.6151
R771 B.n162 B.n161 10.6151
R772 B.n163 B.n162 10.6151
R773 B.n163 B.n146 10.6151
R774 B.n167 B.n146 10.6151
R775 B.n168 B.n167 10.6151
R776 B.n169 B.n168 10.6151
R777 B.n169 B.n144 10.6151
R778 B.n173 B.n144 10.6151
R779 B.n174 B.n173 10.6151
R780 B.n175 B.n174 10.6151
R781 B.n175 B.n142 10.6151
R782 B.n179 B.n142 10.6151
R783 B.n180 B.n179 10.6151
R784 B.n181 B.n180 10.6151
R785 B.n181 B.n140 10.6151
R786 B.n185 B.n140 10.6151
R787 B.n186 B.n185 10.6151
R788 B.n187 B.n186 10.6151
R789 B.n191 B.n138 10.6151
R790 B.n192 B.n191 10.6151
R791 B.n193 B.n192 10.6151
R792 B.n193 B.n136 10.6151
R793 B.n197 B.n136 10.6151
R794 B.n198 B.n197 10.6151
R795 B.n199 B.n198 10.6151
R796 B.n199 B.n134 10.6151
R797 B.n203 B.n134 10.6151
R798 B.n204 B.n203 10.6151
R799 B.n205 B.n204 10.6151
R800 B.n205 B.n132 10.6151
R801 B.n209 B.n132 10.6151
R802 B.n210 B.n209 10.6151
R803 B.n211 B.n210 10.6151
R804 B.n211 B.n130 10.6151
R805 B.n215 B.n130 10.6151
R806 B.n216 B.n215 10.6151
R807 B.n217 B.n216 10.6151
R808 B.n217 B.n128 10.6151
R809 B.n221 B.n128 10.6151
R810 B.n222 B.n221 10.6151
R811 B.n223 B.n222 10.6151
R812 B.n223 B.n126 10.6151
R813 B.n227 B.n126 10.6151
R814 B.n228 B.n227 10.6151
R815 B.n229 B.n228 10.6151
R816 B.n229 B.n124 10.6151
R817 B.n233 B.n124 10.6151
R818 B.n234 B.n233 10.6151
R819 B.n235 B.n234 10.6151
R820 B.n235 B.n122 10.6151
R821 B.n239 B.n122 10.6151
R822 B.n240 B.n239 10.6151
R823 B.n241 B.n240 10.6151
R824 B.n241 B.n120 10.6151
R825 B.n245 B.n120 10.6151
R826 B.n246 B.n245 10.6151
R827 B.n250 B.n246 10.6151
R828 B.n254 B.n118 10.6151
R829 B.n255 B.n254 10.6151
R830 B.n256 B.n255 10.6151
R831 B.n256 B.n116 10.6151
R832 B.n260 B.n116 10.6151
R833 B.n261 B.n260 10.6151
R834 B.n262 B.n261 10.6151
R835 B.n262 B.n114 10.6151
R836 B.n266 B.n114 10.6151
R837 B.n269 B.n268 10.6151
R838 B.n269 B.n110 10.6151
R839 B.n273 B.n110 10.6151
R840 B.n274 B.n273 10.6151
R841 B.n275 B.n274 10.6151
R842 B.n275 B.n108 10.6151
R843 B.n279 B.n108 10.6151
R844 B.n280 B.n279 10.6151
R845 B.n281 B.n280 10.6151
R846 B.n281 B.n106 10.6151
R847 B.n285 B.n106 10.6151
R848 B.n286 B.n285 10.6151
R849 B.n287 B.n286 10.6151
R850 B.n287 B.n104 10.6151
R851 B.n291 B.n104 10.6151
R852 B.n292 B.n291 10.6151
R853 B.n293 B.n292 10.6151
R854 B.n293 B.n102 10.6151
R855 B.n297 B.n102 10.6151
R856 B.n298 B.n297 10.6151
R857 B.n299 B.n298 10.6151
R858 B.n299 B.n100 10.6151
R859 B.n303 B.n100 10.6151
R860 B.n304 B.n303 10.6151
R861 B.n305 B.n304 10.6151
R862 B.n305 B.n98 10.6151
R863 B.n309 B.n98 10.6151
R864 B.n310 B.n309 10.6151
R865 B.n311 B.n310 10.6151
R866 B.n311 B.n96 10.6151
R867 B.n315 B.n96 10.6151
R868 B.n316 B.n315 10.6151
R869 B.n317 B.n316 10.6151
R870 B.n317 B.n94 10.6151
R871 B.n321 B.n94 10.6151
R872 B.n322 B.n321 10.6151
R873 B.n323 B.n322 10.6151
R874 B.n323 B.n92 10.6151
R875 B.n327 B.n92 10.6151
R876 B.n485 B.n484 9.36635
R877 B.n467 B.n44 9.36635
R878 B.n250 B.n249 9.36635
R879 B.n268 B.n267 9.36635
R880 B.n585 B.n0 8.11757
R881 B.n585 B.n1 8.11757
R882 B.n484 B.n483 1.24928
R883 B.n470 B.n44 1.24928
R884 B.n249 B.n118 1.24928
R885 B.n267 B.n266 1.24928
R886 VP.n3 VP.t2 195.065
R887 VP.n3 VP.t0 194.641
R888 VP.n5 VP.n4 184.054
R889 VP.n14 VP.n13 184.054
R890 VP.n12 VP.n0 161.3
R891 VP.n11 VP.n10 161.3
R892 VP.n9 VP.n1 161.3
R893 VP.n8 VP.n7 161.3
R894 VP.n6 VP.n2 161.3
R895 VP.n5 VP.t3 159.421
R896 VP.n13 VP.t1 159.421
R897 VP.n4 VP.n3 52.6329
R898 VP.n7 VP.n1 40.4934
R899 VP.n11 VP.n1 40.4934
R900 VP.n7 VP.n6 24.4675
R901 VP.n12 VP.n11 24.4675
R902 VP.n6 VP.n5 1.71319
R903 VP.n13 VP.n12 1.71319
R904 VP.n4 VP.n2 0.189894
R905 VP.n8 VP.n2 0.189894
R906 VP.n9 VP.n8 0.189894
R907 VP.n10 VP.n9 0.189894
R908 VP.n10 VP.n0 0.189894
R909 VP.n14 VP.n0 0.189894
R910 VP VP.n14 0.0516364
R911 VTAIL.n490 VTAIL.n434 756.745
R912 VTAIL.n56 VTAIL.n0 756.745
R913 VTAIL.n118 VTAIL.n62 756.745
R914 VTAIL.n180 VTAIL.n124 756.745
R915 VTAIL.n428 VTAIL.n372 756.745
R916 VTAIL.n366 VTAIL.n310 756.745
R917 VTAIL.n304 VTAIL.n248 756.745
R918 VTAIL.n242 VTAIL.n186 756.745
R919 VTAIL.n455 VTAIL.n454 585
R920 VTAIL.n457 VTAIL.n456 585
R921 VTAIL.n450 VTAIL.n449 585
R922 VTAIL.n463 VTAIL.n462 585
R923 VTAIL.n465 VTAIL.n464 585
R924 VTAIL.n446 VTAIL.n445 585
R925 VTAIL.n472 VTAIL.n471 585
R926 VTAIL.n473 VTAIL.n444 585
R927 VTAIL.n475 VTAIL.n474 585
R928 VTAIL.n442 VTAIL.n441 585
R929 VTAIL.n481 VTAIL.n480 585
R930 VTAIL.n483 VTAIL.n482 585
R931 VTAIL.n438 VTAIL.n437 585
R932 VTAIL.n489 VTAIL.n488 585
R933 VTAIL.n491 VTAIL.n490 585
R934 VTAIL.n21 VTAIL.n20 585
R935 VTAIL.n23 VTAIL.n22 585
R936 VTAIL.n16 VTAIL.n15 585
R937 VTAIL.n29 VTAIL.n28 585
R938 VTAIL.n31 VTAIL.n30 585
R939 VTAIL.n12 VTAIL.n11 585
R940 VTAIL.n38 VTAIL.n37 585
R941 VTAIL.n39 VTAIL.n10 585
R942 VTAIL.n41 VTAIL.n40 585
R943 VTAIL.n8 VTAIL.n7 585
R944 VTAIL.n47 VTAIL.n46 585
R945 VTAIL.n49 VTAIL.n48 585
R946 VTAIL.n4 VTAIL.n3 585
R947 VTAIL.n55 VTAIL.n54 585
R948 VTAIL.n57 VTAIL.n56 585
R949 VTAIL.n83 VTAIL.n82 585
R950 VTAIL.n85 VTAIL.n84 585
R951 VTAIL.n78 VTAIL.n77 585
R952 VTAIL.n91 VTAIL.n90 585
R953 VTAIL.n93 VTAIL.n92 585
R954 VTAIL.n74 VTAIL.n73 585
R955 VTAIL.n100 VTAIL.n99 585
R956 VTAIL.n101 VTAIL.n72 585
R957 VTAIL.n103 VTAIL.n102 585
R958 VTAIL.n70 VTAIL.n69 585
R959 VTAIL.n109 VTAIL.n108 585
R960 VTAIL.n111 VTAIL.n110 585
R961 VTAIL.n66 VTAIL.n65 585
R962 VTAIL.n117 VTAIL.n116 585
R963 VTAIL.n119 VTAIL.n118 585
R964 VTAIL.n145 VTAIL.n144 585
R965 VTAIL.n147 VTAIL.n146 585
R966 VTAIL.n140 VTAIL.n139 585
R967 VTAIL.n153 VTAIL.n152 585
R968 VTAIL.n155 VTAIL.n154 585
R969 VTAIL.n136 VTAIL.n135 585
R970 VTAIL.n162 VTAIL.n161 585
R971 VTAIL.n163 VTAIL.n134 585
R972 VTAIL.n165 VTAIL.n164 585
R973 VTAIL.n132 VTAIL.n131 585
R974 VTAIL.n171 VTAIL.n170 585
R975 VTAIL.n173 VTAIL.n172 585
R976 VTAIL.n128 VTAIL.n127 585
R977 VTAIL.n179 VTAIL.n178 585
R978 VTAIL.n181 VTAIL.n180 585
R979 VTAIL.n429 VTAIL.n428 585
R980 VTAIL.n427 VTAIL.n426 585
R981 VTAIL.n376 VTAIL.n375 585
R982 VTAIL.n421 VTAIL.n420 585
R983 VTAIL.n419 VTAIL.n418 585
R984 VTAIL.n380 VTAIL.n379 585
R985 VTAIL.n384 VTAIL.n382 585
R986 VTAIL.n413 VTAIL.n412 585
R987 VTAIL.n411 VTAIL.n410 585
R988 VTAIL.n386 VTAIL.n385 585
R989 VTAIL.n405 VTAIL.n404 585
R990 VTAIL.n403 VTAIL.n402 585
R991 VTAIL.n390 VTAIL.n389 585
R992 VTAIL.n397 VTAIL.n396 585
R993 VTAIL.n395 VTAIL.n394 585
R994 VTAIL.n367 VTAIL.n366 585
R995 VTAIL.n365 VTAIL.n364 585
R996 VTAIL.n314 VTAIL.n313 585
R997 VTAIL.n359 VTAIL.n358 585
R998 VTAIL.n357 VTAIL.n356 585
R999 VTAIL.n318 VTAIL.n317 585
R1000 VTAIL.n322 VTAIL.n320 585
R1001 VTAIL.n351 VTAIL.n350 585
R1002 VTAIL.n349 VTAIL.n348 585
R1003 VTAIL.n324 VTAIL.n323 585
R1004 VTAIL.n343 VTAIL.n342 585
R1005 VTAIL.n341 VTAIL.n340 585
R1006 VTAIL.n328 VTAIL.n327 585
R1007 VTAIL.n335 VTAIL.n334 585
R1008 VTAIL.n333 VTAIL.n332 585
R1009 VTAIL.n305 VTAIL.n304 585
R1010 VTAIL.n303 VTAIL.n302 585
R1011 VTAIL.n252 VTAIL.n251 585
R1012 VTAIL.n297 VTAIL.n296 585
R1013 VTAIL.n295 VTAIL.n294 585
R1014 VTAIL.n256 VTAIL.n255 585
R1015 VTAIL.n260 VTAIL.n258 585
R1016 VTAIL.n289 VTAIL.n288 585
R1017 VTAIL.n287 VTAIL.n286 585
R1018 VTAIL.n262 VTAIL.n261 585
R1019 VTAIL.n281 VTAIL.n280 585
R1020 VTAIL.n279 VTAIL.n278 585
R1021 VTAIL.n266 VTAIL.n265 585
R1022 VTAIL.n273 VTAIL.n272 585
R1023 VTAIL.n271 VTAIL.n270 585
R1024 VTAIL.n243 VTAIL.n242 585
R1025 VTAIL.n241 VTAIL.n240 585
R1026 VTAIL.n190 VTAIL.n189 585
R1027 VTAIL.n235 VTAIL.n234 585
R1028 VTAIL.n233 VTAIL.n232 585
R1029 VTAIL.n194 VTAIL.n193 585
R1030 VTAIL.n198 VTAIL.n196 585
R1031 VTAIL.n227 VTAIL.n226 585
R1032 VTAIL.n225 VTAIL.n224 585
R1033 VTAIL.n200 VTAIL.n199 585
R1034 VTAIL.n219 VTAIL.n218 585
R1035 VTAIL.n217 VTAIL.n216 585
R1036 VTAIL.n204 VTAIL.n203 585
R1037 VTAIL.n211 VTAIL.n210 585
R1038 VTAIL.n209 VTAIL.n208 585
R1039 VTAIL.n453 VTAIL.t1 329.036
R1040 VTAIL.n19 VTAIL.t3 329.036
R1041 VTAIL.n81 VTAIL.t5 329.036
R1042 VTAIL.n143 VTAIL.t7 329.036
R1043 VTAIL.n393 VTAIL.t6 329.036
R1044 VTAIL.n331 VTAIL.t4 329.036
R1045 VTAIL.n269 VTAIL.t2 329.036
R1046 VTAIL.n207 VTAIL.t0 329.036
R1047 VTAIL.n456 VTAIL.n455 171.744
R1048 VTAIL.n456 VTAIL.n449 171.744
R1049 VTAIL.n463 VTAIL.n449 171.744
R1050 VTAIL.n464 VTAIL.n463 171.744
R1051 VTAIL.n464 VTAIL.n445 171.744
R1052 VTAIL.n472 VTAIL.n445 171.744
R1053 VTAIL.n473 VTAIL.n472 171.744
R1054 VTAIL.n474 VTAIL.n473 171.744
R1055 VTAIL.n474 VTAIL.n441 171.744
R1056 VTAIL.n481 VTAIL.n441 171.744
R1057 VTAIL.n482 VTAIL.n481 171.744
R1058 VTAIL.n482 VTAIL.n437 171.744
R1059 VTAIL.n489 VTAIL.n437 171.744
R1060 VTAIL.n490 VTAIL.n489 171.744
R1061 VTAIL.n22 VTAIL.n21 171.744
R1062 VTAIL.n22 VTAIL.n15 171.744
R1063 VTAIL.n29 VTAIL.n15 171.744
R1064 VTAIL.n30 VTAIL.n29 171.744
R1065 VTAIL.n30 VTAIL.n11 171.744
R1066 VTAIL.n38 VTAIL.n11 171.744
R1067 VTAIL.n39 VTAIL.n38 171.744
R1068 VTAIL.n40 VTAIL.n39 171.744
R1069 VTAIL.n40 VTAIL.n7 171.744
R1070 VTAIL.n47 VTAIL.n7 171.744
R1071 VTAIL.n48 VTAIL.n47 171.744
R1072 VTAIL.n48 VTAIL.n3 171.744
R1073 VTAIL.n55 VTAIL.n3 171.744
R1074 VTAIL.n56 VTAIL.n55 171.744
R1075 VTAIL.n84 VTAIL.n83 171.744
R1076 VTAIL.n84 VTAIL.n77 171.744
R1077 VTAIL.n91 VTAIL.n77 171.744
R1078 VTAIL.n92 VTAIL.n91 171.744
R1079 VTAIL.n92 VTAIL.n73 171.744
R1080 VTAIL.n100 VTAIL.n73 171.744
R1081 VTAIL.n101 VTAIL.n100 171.744
R1082 VTAIL.n102 VTAIL.n101 171.744
R1083 VTAIL.n102 VTAIL.n69 171.744
R1084 VTAIL.n109 VTAIL.n69 171.744
R1085 VTAIL.n110 VTAIL.n109 171.744
R1086 VTAIL.n110 VTAIL.n65 171.744
R1087 VTAIL.n117 VTAIL.n65 171.744
R1088 VTAIL.n118 VTAIL.n117 171.744
R1089 VTAIL.n146 VTAIL.n145 171.744
R1090 VTAIL.n146 VTAIL.n139 171.744
R1091 VTAIL.n153 VTAIL.n139 171.744
R1092 VTAIL.n154 VTAIL.n153 171.744
R1093 VTAIL.n154 VTAIL.n135 171.744
R1094 VTAIL.n162 VTAIL.n135 171.744
R1095 VTAIL.n163 VTAIL.n162 171.744
R1096 VTAIL.n164 VTAIL.n163 171.744
R1097 VTAIL.n164 VTAIL.n131 171.744
R1098 VTAIL.n171 VTAIL.n131 171.744
R1099 VTAIL.n172 VTAIL.n171 171.744
R1100 VTAIL.n172 VTAIL.n127 171.744
R1101 VTAIL.n179 VTAIL.n127 171.744
R1102 VTAIL.n180 VTAIL.n179 171.744
R1103 VTAIL.n428 VTAIL.n427 171.744
R1104 VTAIL.n427 VTAIL.n375 171.744
R1105 VTAIL.n420 VTAIL.n375 171.744
R1106 VTAIL.n420 VTAIL.n419 171.744
R1107 VTAIL.n419 VTAIL.n379 171.744
R1108 VTAIL.n384 VTAIL.n379 171.744
R1109 VTAIL.n412 VTAIL.n384 171.744
R1110 VTAIL.n412 VTAIL.n411 171.744
R1111 VTAIL.n411 VTAIL.n385 171.744
R1112 VTAIL.n404 VTAIL.n385 171.744
R1113 VTAIL.n404 VTAIL.n403 171.744
R1114 VTAIL.n403 VTAIL.n389 171.744
R1115 VTAIL.n396 VTAIL.n389 171.744
R1116 VTAIL.n396 VTAIL.n395 171.744
R1117 VTAIL.n366 VTAIL.n365 171.744
R1118 VTAIL.n365 VTAIL.n313 171.744
R1119 VTAIL.n358 VTAIL.n313 171.744
R1120 VTAIL.n358 VTAIL.n357 171.744
R1121 VTAIL.n357 VTAIL.n317 171.744
R1122 VTAIL.n322 VTAIL.n317 171.744
R1123 VTAIL.n350 VTAIL.n322 171.744
R1124 VTAIL.n350 VTAIL.n349 171.744
R1125 VTAIL.n349 VTAIL.n323 171.744
R1126 VTAIL.n342 VTAIL.n323 171.744
R1127 VTAIL.n342 VTAIL.n341 171.744
R1128 VTAIL.n341 VTAIL.n327 171.744
R1129 VTAIL.n334 VTAIL.n327 171.744
R1130 VTAIL.n334 VTAIL.n333 171.744
R1131 VTAIL.n304 VTAIL.n303 171.744
R1132 VTAIL.n303 VTAIL.n251 171.744
R1133 VTAIL.n296 VTAIL.n251 171.744
R1134 VTAIL.n296 VTAIL.n295 171.744
R1135 VTAIL.n295 VTAIL.n255 171.744
R1136 VTAIL.n260 VTAIL.n255 171.744
R1137 VTAIL.n288 VTAIL.n260 171.744
R1138 VTAIL.n288 VTAIL.n287 171.744
R1139 VTAIL.n287 VTAIL.n261 171.744
R1140 VTAIL.n280 VTAIL.n261 171.744
R1141 VTAIL.n280 VTAIL.n279 171.744
R1142 VTAIL.n279 VTAIL.n265 171.744
R1143 VTAIL.n272 VTAIL.n265 171.744
R1144 VTAIL.n272 VTAIL.n271 171.744
R1145 VTAIL.n242 VTAIL.n241 171.744
R1146 VTAIL.n241 VTAIL.n189 171.744
R1147 VTAIL.n234 VTAIL.n189 171.744
R1148 VTAIL.n234 VTAIL.n233 171.744
R1149 VTAIL.n233 VTAIL.n193 171.744
R1150 VTAIL.n198 VTAIL.n193 171.744
R1151 VTAIL.n226 VTAIL.n198 171.744
R1152 VTAIL.n226 VTAIL.n225 171.744
R1153 VTAIL.n225 VTAIL.n199 171.744
R1154 VTAIL.n218 VTAIL.n199 171.744
R1155 VTAIL.n218 VTAIL.n217 171.744
R1156 VTAIL.n217 VTAIL.n203 171.744
R1157 VTAIL.n210 VTAIL.n203 171.744
R1158 VTAIL.n210 VTAIL.n209 171.744
R1159 VTAIL.n455 VTAIL.t1 85.8723
R1160 VTAIL.n21 VTAIL.t3 85.8723
R1161 VTAIL.n83 VTAIL.t5 85.8723
R1162 VTAIL.n145 VTAIL.t7 85.8723
R1163 VTAIL.n395 VTAIL.t6 85.8723
R1164 VTAIL.n333 VTAIL.t4 85.8723
R1165 VTAIL.n271 VTAIL.t2 85.8723
R1166 VTAIL.n209 VTAIL.t0 85.8723
R1167 VTAIL.n495 VTAIL.n494 34.3187
R1168 VTAIL.n61 VTAIL.n60 34.3187
R1169 VTAIL.n123 VTAIL.n122 34.3187
R1170 VTAIL.n185 VTAIL.n184 34.3187
R1171 VTAIL.n433 VTAIL.n432 34.3187
R1172 VTAIL.n371 VTAIL.n370 34.3187
R1173 VTAIL.n309 VTAIL.n308 34.3187
R1174 VTAIL.n247 VTAIL.n246 34.3187
R1175 VTAIL.n495 VTAIL.n433 24.0738
R1176 VTAIL.n247 VTAIL.n185 24.0738
R1177 VTAIL.n475 VTAIL.n442 13.1884
R1178 VTAIL.n41 VTAIL.n8 13.1884
R1179 VTAIL.n103 VTAIL.n70 13.1884
R1180 VTAIL.n165 VTAIL.n132 13.1884
R1181 VTAIL.n382 VTAIL.n380 13.1884
R1182 VTAIL.n320 VTAIL.n318 13.1884
R1183 VTAIL.n258 VTAIL.n256 13.1884
R1184 VTAIL.n196 VTAIL.n194 13.1884
R1185 VTAIL.n476 VTAIL.n444 12.8005
R1186 VTAIL.n480 VTAIL.n479 12.8005
R1187 VTAIL.n42 VTAIL.n10 12.8005
R1188 VTAIL.n46 VTAIL.n45 12.8005
R1189 VTAIL.n104 VTAIL.n72 12.8005
R1190 VTAIL.n108 VTAIL.n107 12.8005
R1191 VTAIL.n166 VTAIL.n134 12.8005
R1192 VTAIL.n170 VTAIL.n169 12.8005
R1193 VTAIL.n418 VTAIL.n417 12.8005
R1194 VTAIL.n414 VTAIL.n413 12.8005
R1195 VTAIL.n356 VTAIL.n355 12.8005
R1196 VTAIL.n352 VTAIL.n351 12.8005
R1197 VTAIL.n294 VTAIL.n293 12.8005
R1198 VTAIL.n290 VTAIL.n289 12.8005
R1199 VTAIL.n232 VTAIL.n231 12.8005
R1200 VTAIL.n228 VTAIL.n227 12.8005
R1201 VTAIL.n471 VTAIL.n470 12.0247
R1202 VTAIL.n483 VTAIL.n440 12.0247
R1203 VTAIL.n37 VTAIL.n36 12.0247
R1204 VTAIL.n49 VTAIL.n6 12.0247
R1205 VTAIL.n99 VTAIL.n98 12.0247
R1206 VTAIL.n111 VTAIL.n68 12.0247
R1207 VTAIL.n161 VTAIL.n160 12.0247
R1208 VTAIL.n173 VTAIL.n130 12.0247
R1209 VTAIL.n421 VTAIL.n378 12.0247
R1210 VTAIL.n410 VTAIL.n383 12.0247
R1211 VTAIL.n359 VTAIL.n316 12.0247
R1212 VTAIL.n348 VTAIL.n321 12.0247
R1213 VTAIL.n297 VTAIL.n254 12.0247
R1214 VTAIL.n286 VTAIL.n259 12.0247
R1215 VTAIL.n235 VTAIL.n192 12.0247
R1216 VTAIL.n224 VTAIL.n197 12.0247
R1217 VTAIL.n469 VTAIL.n446 11.249
R1218 VTAIL.n484 VTAIL.n438 11.249
R1219 VTAIL.n35 VTAIL.n12 11.249
R1220 VTAIL.n50 VTAIL.n4 11.249
R1221 VTAIL.n97 VTAIL.n74 11.249
R1222 VTAIL.n112 VTAIL.n66 11.249
R1223 VTAIL.n159 VTAIL.n136 11.249
R1224 VTAIL.n174 VTAIL.n128 11.249
R1225 VTAIL.n422 VTAIL.n376 11.249
R1226 VTAIL.n409 VTAIL.n386 11.249
R1227 VTAIL.n360 VTAIL.n314 11.249
R1228 VTAIL.n347 VTAIL.n324 11.249
R1229 VTAIL.n298 VTAIL.n252 11.249
R1230 VTAIL.n285 VTAIL.n262 11.249
R1231 VTAIL.n236 VTAIL.n190 11.249
R1232 VTAIL.n223 VTAIL.n200 11.249
R1233 VTAIL.n454 VTAIL.n453 10.7239
R1234 VTAIL.n20 VTAIL.n19 10.7239
R1235 VTAIL.n82 VTAIL.n81 10.7239
R1236 VTAIL.n144 VTAIL.n143 10.7239
R1237 VTAIL.n394 VTAIL.n393 10.7239
R1238 VTAIL.n332 VTAIL.n331 10.7239
R1239 VTAIL.n270 VTAIL.n269 10.7239
R1240 VTAIL.n208 VTAIL.n207 10.7239
R1241 VTAIL.n466 VTAIL.n465 10.4732
R1242 VTAIL.n488 VTAIL.n487 10.4732
R1243 VTAIL.n32 VTAIL.n31 10.4732
R1244 VTAIL.n54 VTAIL.n53 10.4732
R1245 VTAIL.n94 VTAIL.n93 10.4732
R1246 VTAIL.n116 VTAIL.n115 10.4732
R1247 VTAIL.n156 VTAIL.n155 10.4732
R1248 VTAIL.n178 VTAIL.n177 10.4732
R1249 VTAIL.n426 VTAIL.n425 10.4732
R1250 VTAIL.n406 VTAIL.n405 10.4732
R1251 VTAIL.n364 VTAIL.n363 10.4732
R1252 VTAIL.n344 VTAIL.n343 10.4732
R1253 VTAIL.n302 VTAIL.n301 10.4732
R1254 VTAIL.n282 VTAIL.n281 10.4732
R1255 VTAIL.n240 VTAIL.n239 10.4732
R1256 VTAIL.n220 VTAIL.n219 10.4732
R1257 VTAIL.n462 VTAIL.n448 9.69747
R1258 VTAIL.n491 VTAIL.n436 9.69747
R1259 VTAIL.n28 VTAIL.n14 9.69747
R1260 VTAIL.n57 VTAIL.n2 9.69747
R1261 VTAIL.n90 VTAIL.n76 9.69747
R1262 VTAIL.n119 VTAIL.n64 9.69747
R1263 VTAIL.n152 VTAIL.n138 9.69747
R1264 VTAIL.n181 VTAIL.n126 9.69747
R1265 VTAIL.n429 VTAIL.n374 9.69747
R1266 VTAIL.n402 VTAIL.n388 9.69747
R1267 VTAIL.n367 VTAIL.n312 9.69747
R1268 VTAIL.n340 VTAIL.n326 9.69747
R1269 VTAIL.n305 VTAIL.n250 9.69747
R1270 VTAIL.n278 VTAIL.n264 9.69747
R1271 VTAIL.n243 VTAIL.n188 9.69747
R1272 VTAIL.n216 VTAIL.n202 9.69747
R1273 VTAIL.n494 VTAIL.n493 9.45567
R1274 VTAIL.n60 VTAIL.n59 9.45567
R1275 VTAIL.n122 VTAIL.n121 9.45567
R1276 VTAIL.n184 VTAIL.n183 9.45567
R1277 VTAIL.n432 VTAIL.n431 9.45567
R1278 VTAIL.n370 VTAIL.n369 9.45567
R1279 VTAIL.n308 VTAIL.n307 9.45567
R1280 VTAIL.n246 VTAIL.n245 9.45567
R1281 VTAIL.n493 VTAIL.n492 9.3005
R1282 VTAIL.n436 VTAIL.n435 9.3005
R1283 VTAIL.n487 VTAIL.n486 9.3005
R1284 VTAIL.n485 VTAIL.n484 9.3005
R1285 VTAIL.n440 VTAIL.n439 9.3005
R1286 VTAIL.n479 VTAIL.n478 9.3005
R1287 VTAIL.n452 VTAIL.n451 9.3005
R1288 VTAIL.n459 VTAIL.n458 9.3005
R1289 VTAIL.n461 VTAIL.n460 9.3005
R1290 VTAIL.n448 VTAIL.n447 9.3005
R1291 VTAIL.n467 VTAIL.n466 9.3005
R1292 VTAIL.n469 VTAIL.n468 9.3005
R1293 VTAIL.n470 VTAIL.n443 9.3005
R1294 VTAIL.n477 VTAIL.n476 9.3005
R1295 VTAIL.n59 VTAIL.n58 9.3005
R1296 VTAIL.n2 VTAIL.n1 9.3005
R1297 VTAIL.n53 VTAIL.n52 9.3005
R1298 VTAIL.n51 VTAIL.n50 9.3005
R1299 VTAIL.n6 VTAIL.n5 9.3005
R1300 VTAIL.n45 VTAIL.n44 9.3005
R1301 VTAIL.n18 VTAIL.n17 9.3005
R1302 VTAIL.n25 VTAIL.n24 9.3005
R1303 VTAIL.n27 VTAIL.n26 9.3005
R1304 VTAIL.n14 VTAIL.n13 9.3005
R1305 VTAIL.n33 VTAIL.n32 9.3005
R1306 VTAIL.n35 VTAIL.n34 9.3005
R1307 VTAIL.n36 VTAIL.n9 9.3005
R1308 VTAIL.n43 VTAIL.n42 9.3005
R1309 VTAIL.n121 VTAIL.n120 9.3005
R1310 VTAIL.n64 VTAIL.n63 9.3005
R1311 VTAIL.n115 VTAIL.n114 9.3005
R1312 VTAIL.n113 VTAIL.n112 9.3005
R1313 VTAIL.n68 VTAIL.n67 9.3005
R1314 VTAIL.n107 VTAIL.n106 9.3005
R1315 VTAIL.n80 VTAIL.n79 9.3005
R1316 VTAIL.n87 VTAIL.n86 9.3005
R1317 VTAIL.n89 VTAIL.n88 9.3005
R1318 VTAIL.n76 VTAIL.n75 9.3005
R1319 VTAIL.n95 VTAIL.n94 9.3005
R1320 VTAIL.n97 VTAIL.n96 9.3005
R1321 VTAIL.n98 VTAIL.n71 9.3005
R1322 VTAIL.n105 VTAIL.n104 9.3005
R1323 VTAIL.n183 VTAIL.n182 9.3005
R1324 VTAIL.n126 VTAIL.n125 9.3005
R1325 VTAIL.n177 VTAIL.n176 9.3005
R1326 VTAIL.n175 VTAIL.n174 9.3005
R1327 VTAIL.n130 VTAIL.n129 9.3005
R1328 VTAIL.n169 VTAIL.n168 9.3005
R1329 VTAIL.n142 VTAIL.n141 9.3005
R1330 VTAIL.n149 VTAIL.n148 9.3005
R1331 VTAIL.n151 VTAIL.n150 9.3005
R1332 VTAIL.n138 VTAIL.n137 9.3005
R1333 VTAIL.n157 VTAIL.n156 9.3005
R1334 VTAIL.n159 VTAIL.n158 9.3005
R1335 VTAIL.n160 VTAIL.n133 9.3005
R1336 VTAIL.n167 VTAIL.n166 9.3005
R1337 VTAIL.n392 VTAIL.n391 9.3005
R1338 VTAIL.n399 VTAIL.n398 9.3005
R1339 VTAIL.n401 VTAIL.n400 9.3005
R1340 VTAIL.n388 VTAIL.n387 9.3005
R1341 VTAIL.n407 VTAIL.n406 9.3005
R1342 VTAIL.n409 VTAIL.n408 9.3005
R1343 VTAIL.n383 VTAIL.n381 9.3005
R1344 VTAIL.n415 VTAIL.n414 9.3005
R1345 VTAIL.n431 VTAIL.n430 9.3005
R1346 VTAIL.n374 VTAIL.n373 9.3005
R1347 VTAIL.n425 VTAIL.n424 9.3005
R1348 VTAIL.n423 VTAIL.n422 9.3005
R1349 VTAIL.n378 VTAIL.n377 9.3005
R1350 VTAIL.n417 VTAIL.n416 9.3005
R1351 VTAIL.n330 VTAIL.n329 9.3005
R1352 VTAIL.n337 VTAIL.n336 9.3005
R1353 VTAIL.n339 VTAIL.n338 9.3005
R1354 VTAIL.n326 VTAIL.n325 9.3005
R1355 VTAIL.n345 VTAIL.n344 9.3005
R1356 VTAIL.n347 VTAIL.n346 9.3005
R1357 VTAIL.n321 VTAIL.n319 9.3005
R1358 VTAIL.n353 VTAIL.n352 9.3005
R1359 VTAIL.n369 VTAIL.n368 9.3005
R1360 VTAIL.n312 VTAIL.n311 9.3005
R1361 VTAIL.n363 VTAIL.n362 9.3005
R1362 VTAIL.n361 VTAIL.n360 9.3005
R1363 VTAIL.n316 VTAIL.n315 9.3005
R1364 VTAIL.n355 VTAIL.n354 9.3005
R1365 VTAIL.n268 VTAIL.n267 9.3005
R1366 VTAIL.n275 VTAIL.n274 9.3005
R1367 VTAIL.n277 VTAIL.n276 9.3005
R1368 VTAIL.n264 VTAIL.n263 9.3005
R1369 VTAIL.n283 VTAIL.n282 9.3005
R1370 VTAIL.n285 VTAIL.n284 9.3005
R1371 VTAIL.n259 VTAIL.n257 9.3005
R1372 VTAIL.n291 VTAIL.n290 9.3005
R1373 VTAIL.n307 VTAIL.n306 9.3005
R1374 VTAIL.n250 VTAIL.n249 9.3005
R1375 VTAIL.n301 VTAIL.n300 9.3005
R1376 VTAIL.n299 VTAIL.n298 9.3005
R1377 VTAIL.n254 VTAIL.n253 9.3005
R1378 VTAIL.n293 VTAIL.n292 9.3005
R1379 VTAIL.n206 VTAIL.n205 9.3005
R1380 VTAIL.n213 VTAIL.n212 9.3005
R1381 VTAIL.n215 VTAIL.n214 9.3005
R1382 VTAIL.n202 VTAIL.n201 9.3005
R1383 VTAIL.n221 VTAIL.n220 9.3005
R1384 VTAIL.n223 VTAIL.n222 9.3005
R1385 VTAIL.n197 VTAIL.n195 9.3005
R1386 VTAIL.n229 VTAIL.n228 9.3005
R1387 VTAIL.n245 VTAIL.n244 9.3005
R1388 VTAIL.n188 VTAIL.n187 9.3005
R1389 VTAIL.n239 VTAIL.n238 9.3005
R1390 VTAIL.n237 VTAIL.n236 9.3005
R1391 VTAIL.n192 VTAIL.n191 9.3005
R1392 VTAIL.n231 VTAIL.n230 9.3005
R1393 VTAIL.n461 VTAIL.n450 8.92171
R1394 VTAIL.n492 VTAIL.n434 8.92171
R1395 VTAIL.n27 VTAIL.n16 8.92171
R1396 VTAIL.n58 VTAIL.n0 8.92171
R1397 VTAIL.n89 VTAIL.n78 8.92171
R1398 VTAIL.n120 VTAIL.n62 8.92171
R1399 VTAIL.n151 VTAIL.n140 8.92171
R1400 VTAIL.n182 VTAIL.n124 8.92171
R1401 VTAIL.n430 VTAIL.n372 8.92171
R1402 VTAIL.n401 VTAIL.n390 8.92171
R1403 VTAIL.n368 VTAIL.n310 8.92171
R1404 VTAIL.n339 VTAIL.n328 8.92171
R1405 VTAIL.n306 VTAIL.n248 8.92171
R1406 VTAIL.n277 VTAIL.n266 8.92171
R1407 VTAIL.n244 VTAIL.n186 8.92171
R1408 VTAIL.n215 VTAIL.n204 8.92171
R1409 VTAIL.n458 VTAIL.n457 8.14595
R1410 VTAIL.n24 VTAIL.n23 8.14595
R1411 VTAIL.n86 VTAIL.n85 8.14595
R1412 VTAIL.n148 VTAIL.n147 8.14595
R1413 VTAIL.n398 VTAIL.n397 8.14595
R1414 VTAIL.n336 VTAIL.n335 8.14595
R1415 VTAIL.n274 VTAIL.n273 8.14595
R1416 VTAIL.n212 VTAIL.n211 8.14595
R1417 VTAIL.n454 VTAIL.n452 7.3702
R1418 VTAIL.n20 VTAIL.n18 7.3702
R1419 VTAIL.n82 VTAIL.n80 7.3702
R1420 VTAIL.n144 VTAIL.n142 7.3702
R1421 VTAIL.n394 VTAIL.n392 7.3702
R1422 VTAIL.n332 VTAIL.n330 7.3702
R1423 VTAIL.n270 VTAIL.n268 7.3702
R1424 VTAIL.n208 VTAIL.n206 7.3702
R1425 VTAIL.n457 VTAIL.n452 5.81868
R1426 VTAIL.n23 VTAIL.n18 5.81868
R1427 VTAIL.n85 VTAIL.n80 5.81868
R1428 VTAIL.n147 VTAIL.n142 5.81868
R1429 VTAIL.n397 VTAIL.n392 5.81868
R1430 VTAIL.n335 VTAIL.n330 5.81868
R1431 VTAIL.n273 VTAIL.n268 5.81868
R1432 VTAIL.n211 VTAIL.n206 5.81868
R1433 VTAIL.n458 VTAIL.n450 5.04292
R1434 VTAIL.n494 VTAIL.n434 5.04292
R1435 VTAIL.n24 VTAIL.n16 5.04292
R1436 VTAIL.n60 VTAIL.n0 5.04292
R1437 VTAIL.n86 VTAIL.n78 5.04292
R1438 VTAIL.n122 VTAIL.n62 5.04292
R1439 VTAIL.n148 VTAIL.n140 5.04292
R1440 VTAIL.n184 VTAIL.n124 5.04292
R1441 VTAIL.n432 VTAIL.n372 5.04292
R1442 VTAIL.n398 VTAIL.n390 5.04292
R1443 VTAIL.n370 VTAIL.n310 5.04292
R1444 VTAIL.n336 VTAIL.n328 5.04292
R1445 VTAIL.n308 VTAIL.n248 5.04292
R1446 VTAIL.n274 VTAIL.n266 5.04292
R1447 VTAIL.n246 VTAIL.n186 5.04292
R1448 VTAIL.n212 VTAIL.n204 5.04292
R1449 VTAIL.n462 VTAIL.n461 4.26717
R1450 VTAIL.n492 VTAIL.n491 4.26717
R1451 VTAIL.n28 VTAIL.n27 4.26717
R1452 VTAIL.n58 VTAIL.n57 4.26717
R1453 VTAIL.n90 VTAIL.n89 4.26717
R1454 VTAIL.n120 VTAIL.n119 4.26717
R1455 VTAIL.n152 VTAIL.n151 4.26717
R1456 VTAIL.n182 VTAIL.n181 4.26717
R1457 VTAIL.n430 VTAIL.n429 4.26717
R1458 VTAIL.n402 VTAIL.n401 4.26717
R1459 VTAIL.n368 VTAIL.n367 4.26717
R1460 VTAIL.n340 VTAIL.n339 4.26717
R1461 VTAIL.n306 VTAIL.n305 4.26717
R1462 VTAIL.n278 VTAIL.n277 4.26717
R1463 VTAIL.n244 VTAIL.n243 4.26717
R1464 VTAIL.n216 VTAIL.n215 4.26717
R1465 VTAIL.n465 VTAIL.n448 3.49141
R1466 VTAIL.n488 VTAIL.n436 3.49141
R1467 VTAIL.n31 VTAIL.n14 3.49141
R1468 VTAIL.n54 VTAIL.n2 3.49141
R1469 VTAIL.n93 VTAIL.n76 3.49141
R1470 VTAIL.n116 VTAIL.n64 3.49141
R1471 VTAIL.n155 VTAIL.n138 3.49141
R1472 VTAIL.n178 VTAIL.n126 3.49141
R1473 VTAIL.n426 VTAIL.n374 3.49141
R1474 VTAIL.n405 VTAIL.n388 3.49141
R1475 VTAIL.n364 VTAIL.n312 3.49141
R1476 VTAIL.n343 VTAIL.n326 3.49141
R1477 VTAIL.n302 VTAIL.n250 3.49141
R1478 VTAIL.n281 VTAIL.n264 3.49141
R1479 VTAIL.n240 VTAIL.n188 3.49141
R1480 VTAIL.n219 VTAIL.n202 3.49141
R1481 VTAIL.n466 VTAIL.n446 2.71565
R1482 VTAIL.n487 VTAIL.n438 2.71565
R1483 VTAIL.n32 VTAIL.n12 2.71565
R1484 VTAIL.n53 VTAIL.n4 2.71565
R1485 VTAIL.n94 VTAIL.n74 2.71565
R1486 VTAIL.n115 VTAIL.n66 2.71565
R1487 VTAIL.n156 VTAIL.n136 2.71565
R1488 VTAIL.n177 VTAIL.n128 2.71565
R1489 VTAIL.n425 VTAIL.n376 2.71565
R1490 VTAIL.n406 VTAIL.n386 2.71565
R1491 VTAIL.n363 VTAIL.n314 2.71565
R1492 VTAIL.n344 VTAIL.n324 2.71565
R1493 VTAIL.n301 VTAIL.n252 2.71565
R1494 VTAIL.n282 VTAIL.n262 2.71565
R1495 VTAIL.n239 VTAIL.n190 2.71565
R1496 VTAIL.n220 VTAIL.n200 2.71565
R1497 VTAIL.n453 VTAIL.n451 2.41282
R1498 VTAIL.n19 VTAIL.n17 2.41282
R1499 VTAIL.n81 VTAIL.n79 2.41282
R1500 VTAIL.n143 VTAIL.n141 2.41282
R1501 VTAIL.n393 VTAIL.n391 2.41282
R1502 VTAIL.n331 VTAIL.n329 2.41282
R1503 VTAIL.n269 VTAIL.n267 2.41282
R1504 VTAIL.n207 VTAIL.n205 2.41282
R1505 VTAIL.n471 VTAIL.n469 1.93989
R1506 VTAIL.n484 VTAIL.n483 1.93989
R1507 VTAIL.n37 VTAIL.n35 1.93989
R1508 VTAIL.n50 VTAIL.n49 1.93989
R1509 VTAIL.n99 VTAIL.n97 1.93989
R1510 VTAIL.n112 VTAIL.n111 1.93989
R1511 VTAIL.n161 VTAIL.n159 1.93989
R1512 VTAIL.n174 VTAIL.n173 1.93989
R1513 VTAIL.n422 VTAIL.n421 1.93989
R1514 VTAIL.n410 VTAIL.n409 1.93989
R1515 VTAIL.n360 VTAIL.n359 1.93989
R1516 VTAIL.n348 VTAIL.n347 1.93989
R1517 VTAIL.n298 VTAIL.n297 1.93989
R1518 VTAIL.n286 VTAIL.n285 1.93989
R1519 VTAIL.n236 VTAIL.n235 1.93989
R1520 VTAIL.n224 VTAIL.n223 1.93989
R1521 VTAIL.n309 VTAIL.n247 1.78498
R1522 VTAIL.n433 VTAIL.n371 1.78498
R1523 VTAIL.n185 VTAIL.n123 1.78498
R1524 VTAIL.n470 VTAIL.n444 1.16414
R1525 VTAIL.n480 VTAIL.n440 1.16414
R1526 VTAIL.n36 VTAIL.n10 1.16414
R1527 VTAIL.n46 VTAIL.n6 1.16414
R1528 VTAIL.n98 VTAIL.n72 1.16414
R1529 VTAIL.n108 VTAIL.n68 1.16414
R1530 VTAIL.n160 VTAIL.n134 1.16414
R1531 VTAIL.n170 VTAIL.n130 1.16414
R1532 VTAIL.n418 VTAIL.n378 1.16414
R1533 VTAIL.n413 VTAIL.n383 1.16414
R1534 VTAIL.n356 VTAIL.n316 1.16414
R1535 VTAIL.n351 VTAIL.n321 1.16414
R1536 VTAIL.n294 VTAIL.n254 1.16414
R1537 VTAIL.n289 VTAIL.n259 1.16414
R1538 VTAIL.n232 VTAIL.n192 1.16414
R1539 VTAIL.n227 VTAIL.n197 1.16414
R1540 VTAIL VTAIL.n61 0.950931
R1541 VTAIL VTAIL.n495 0.834552
R1542 VTAIL.n371 VTAIL.n309 0.470328
R1543 VTAIL.n123 VTAIL.n61 0.470328
R1544 VTAIL.n476 VTAIL.n475 0.388379
R1545 VTAIL.n479 VTAIL.n442 0.388379
R1546 VTAIL.n42 VTAIL.n41 0.388379
R1547 VTAIL.n45 VTAIL.n8 0.388379
R1548 VTAIL.n104 VTAIL.n103 0.388379
R1549 VTAIL.n107 VTAIL.n70 0.388379
R1550 VTAIL.n166 VTAIL.n165 0.388379
R1551 VTAIL.n169 VTAIL.n132 0.388379
R1552 VTAIL.n417 VTAIL.n380 0.388379
R1553 VTAIL.n414 VTAIL.n382 0.388379
R1554 VTAIL.n355 VTAIL.n318 0.388379
R1555 VTAIL.n352 VTAIL.n320 0.388379
R1556 VTAIL.n293 VTAIL.n256 0.388379
R1557 VTAIL.n290 VTAIL.n258 0.388379
R1558 VTAIL.n231 VTAIL.n194 0.388379
R1559 VTAIL.n228 VTAIL.n196 0.388379
R1560 VTAIL.n459 VTAIL.n451 0.155672
R1561 VTAIL.n460 VTAIL.n459 0.155672
R1562 VTAIL.n460 VTAIL.n447 0.155672
R1563 VTAIL.n467 VTAIL.n447 0.155672
R1564 VTAIL.n468 VTAIL.n467 0.155672
R1565 VTAIL.n468 VTAIL.n443 0.155672
R1566 VTAIL.n477 VTAIL.n443 0.155672
R1567 VTAIL.n478 VTAIL.n477 0.155672
R1568 VTAIL.n478 VTAIL.n439 0.155672
R1569 VTAIL.n485 VTAIL.n439 0.155672
R1570 VTAIL.n486 VTAIL.n485 0.155672
R1571 VTAIL.n486 VTAIL.n435 0.155672
R1572 VTAIL.n493 VTAIL.n435 0.155672
R1573 VTAIL.n25 VTAIL.n17 0.155672
R1574 VTAIL.n26 VTAIL.n25 0.155672
R1575 VTAIL.n26 VTAIL.n13 0.155672
R1576 VTAIL.n33 VTAIL.n13 0.155672
R1577 VTAIL.n34 VTAIL.n33 0.155672
R1578 VTAIL.n34 VTAIL.n9 0.155672
R1579 VTAIL.n43 VTAIL.n9 0.155672
R1580 VTAIL.n44 VTAIL.n43 0.155672
R1581 VTAIL.n44 VTAIL.n5 0.155672
R1582 VTAIL.n51 VTAIL.n5 0.155672
R1583 VTAIL.n52 VTAIL.n51 0.155672
R1584 VTAIL.n52 VTAIL.n1 0.155672
R1585 VTAIL.n59 VTAIL.n1 0.155672
R1586 VTAIL.n87 VTAIL.n79 0.155672
R1587 VTAIL.n88 VTAIL.n87 0.155672
R1588 VTAIL.n88 VTAIL.n75 0.155672
R1589 VTAIL.n95 VTAIL.n75 0.155672
R1590 VTAIL.n96 VTAIL.n95 0.155672
R1591 VTAIL.n96 VTAIL.n71 0.155672
R1592 VTAIL.n105 VTAIL.n71 0.155672
R1593 VTAIL.n106 VTAIL.n105 0.155672
R1594 VTAIL.n106 VTAIL.n67 0.155672
R1595 VTAIL.n113 VTAIL.n67 0.155672
R1596 VTAIL.n114 VTAIL.n113 0.155672
R1597 VTAIL.n114 VTAIL.n63 0.155672
R1598 VTAIL.n121 VTAIL.n63 0.155672
R1599 VTAIL.n149 VTAIL.n141 0.155672
R1600 VTAIL.n150 VTAIL.n149 0.155672
R1601 VTAIL.n150 VTAIL.n137 0.155672
R1602 VTAIL.n157 VTAIL.n137 0.155672
R1603 VTAIL.n158 VTAIL.n157 0.155672
R1604 VTAIL.n158 VTAIL.n133 0.155672
R1605 VTAIL.n167 VTAIL.n133 0.155672
R1606 VTAIL.n168 VTAIL.n167 0.155672
R1607 VTAIL.n168 VTAIL.n129 0.155672
R1608 VTAIL.n175 VTAIL.n129 0.155672
R1609 VTAIL.n176 VTAIL.n175 0.155672
R1610 VTAIL.n176 VTAIL.n125 0.155672
R1611 VTAIL.n183 VTAIL.n125 0.155672
R1612 VTAIL.n431 VTAIL.n373 0.155672
R1613 VTAIL.n424 VTAIL.n373 0.155672
R1614 VTAIL.n424 VTAIL.n423 0.155672
R1615 VTAIL.n423 VTAIL.n377 0.155672
R1616 VTAIL.n416 VTAIL.n377 0.155672
R1617 VTAIL.n416 VTAIL.n415 0.155672
R1618 VTAIL.n415 VTAIL.n381 0.155672
R1619 VTAIL.n408 VTAIL.n381 0.155672
R1620 VTAIL.n408 VTAIL.n407 0.155672
R1621 VTAIL.n407 VTAIL.n387 0.155672
R1622 VTAIL.n400 VTAIL.n387 0.155672
R1623 VTAIL.n400 VTAIL.n399 0.155672
R1624 VTAIL.n399 VTAIL.n391 0.155672
R1625 VTAIL.n369 VTAIL.n311 0.155672
R1626 VTAIL.n362 VTAIL.n311 0.155672
R1627 VTAIL.n362 VTAIL.n361 0.155672
R1628 VTAIL.n361 VTAIL.n315 0.155672
R1629 VTAIL.n354 VTAIL.n315 0.155672
R1630 VTAIL.n354 VTAIL.n353 0.155672
R1631 VTAIL.n353 VTAIL.n319 0.155672
R1632 VTAIL.n346 VTAIL.n319 0.155672
R1633 VTAIL.n346 VTAIL.n345 0.155672
R1634 VTAIL.n345 VTAIL.n325 0.155672
R1635 VTAIL.n338 VTAIL.n325 0.155672
R1636 VTAIL.n338 VTAIL.n337 0.155672
R1637 VTAIL.n337 VTAIL.n329 0.155672
R1638 VTAIL.n307 VTAIL.n249 0.155672
R1639 VTAIL.n300 VTAIL.n249 0.155672
R1640 VTAIL.n300 VTAIL.n299 0.155672
R1641 VTAIL.n299 VTAIL.n253 0.155672
R1642 VTAIL.n292 VTAIL.n253 0.155672
R1643 VTAIL.n292 VTAIL.n291 0.155672
R1644 VTAIL.n291 VTAIL.n257 0.155672
R1645 VTAIL.n284 VTAIL.n257 0.155672
R1646 VTAIL.n284 VTAIL.n283 0.155672
R1647 VTAIL.n283 VTAIL.n263 0.155672
R1648 VTAIL.n276 VTAIL.n263 0.155672
R1649 VTAIL.n276 VTAIL.n275 0.155672
R1650 VTAIL.n275 VTAIL.n267 0.155672
R1651 VTAIL.n245 VTAIL.n187 0.155672
R1652 VTAIL.n238 VTAIL.n187 0.155672
R1653 VTAIL.n238 VTAIL.n237 0.155672
R1654 VTAIL.n237 VTAIL.n191 0.155672
R1655 VTAIL.n230 VTAIL.n191 0.155672
R1656 VTAIL.n230 VTAIL.n229 0.155672
R1657 VTAIL.n229 VTAIL.n195 0.155672
R1658 VTAIL.n222 VTAIL.n195 0.155672
R1659 VTAIL.n222 VTAIL.n221 0.155672
R1660 VTAIL.n221 VTAIL.n201 0.155672
R1661 VTAIL.n214 VTAIL.n201 0.155672
R1662 VTAIL.n214 VTAIL.n213 0.155672
R1663 VTAIL.n213 VTAIL.n205 0.155672
R1664 VDD1 VDD1.n1 116.431
R1665 VDD1 VDD1.n0 76.9743
R1666 VDD1.n0 VDD1.t1 2.82457
R1667 VDD1.n0 VDD1.t3 2.82457
R1668 VDD1.n1 VDD1.t0 2.82457
R1669 VDD1.n1 VDD1.t2 2.82457
R1670 VN.n0 VN.t0 195.065
R1671 VN.n1 VN.t1 195.065
R1672 VN.n0 VN.t2 194.641
R1673 VN.n1 VN.t3 194.641
R1674 VN VN.n1 53.0136
R1675 VN VN.n0 9.46438
R1676 VDD2.n2 VDD2.n0 115.906
R1677 VDD2.n2 VDD2.n1 76.9161
R1678 VDD2.n1 VDD2.t0 2.82457
R1679 VDD2.n1 VDD2.t2 2.82457
R1680 VDD2.n0 VDD2.t3 2.82457
R1681 VDD2.n0 VDD2.t1 2.82457
R1682 VDD2 VDD2.n2 0.0586897
C0 B VN 0.9398f
C1 VP VN 5.48196f
C2 VN w_n2212_n3270# 3.58448f
C3 VP B 1.40407f
C4 VTAIL VN 4.00207f
C5 VN VDD2 4.19523f
C6 B w_n2212_n3270# 8.05f
C7 VP w_n2212_n3270# 3.86667f
C8 VTAIL B 4.36371f
C9 VN VDD1 0.148044f
C10 VTAIL VP 4.01618f
C11 B VDD2 1.1356f
C12 VP VDD2 0.339403f
C13 VTAIL w_n2212_n3270# 3.86451f
C14 B VDD1 1.0975f
C15 VP VDD1 4.38607f
C16 VDD2 w_n2212_n3270# 1.30522f
C17 VTAIL VDD2 5.3426f
C18 VDD1 w_n2212_n3270# 1.26834f
C19 VTAIL VDD1 5.29416f
C20 VDD1 VDD2 0.816882f
C21 VDD2 VSUBS 0.799774f
C22 VDD1 VSUBS 5.211009f
C23 VTAIL VSUBS 1.06317f
C24 VN VSUBS 5.13196f
C25 VP VSUBS 1.798134f
C26 B VSUBS 3.489973f
C27 w_n2212_n3270# VSUBS 89.10821f
C28 VDD2.t3 VSUBS 0.242097f
C29 VDD2.t1 VSUBS 0.242097f
C30 VDD2.n0 VSUBS 2.50175f
C31 VDD2.t0 VSUBS 0.242097f
C32 VDD2.t2 VSUBS 0.242097f
C33 VDD2.n1 VSUBS 1.88271f
C34 VDD2.n2 VSUBS 3.98838f
C35 VN.t0 VSUBS 2.42379f
C36 VN.t2 VSUBS 2.42158f
C37 VN.n0 VSUBS 1.71053f
C38 VN.t1 VSUBS 2.42379f
C39 VN.t3 VSUBS 2.42158f
C40 VN.n1 VSUBS 3.41685f
C41 VDD1.t1 VSUBS 0.244662f
C42 VDD1.t3 VSUBS 0.244662f
C43 VDD1.n0 VSUBS 1.90315f
C44 VDD1.t0 VSUBS 0.244662f
C45 VDD1.t2 VSUBS 0.244662f
C46 VDD1.n1 VSUBS 2.55215f
C47 VTAIL.n0 VSUBS 0.026126f
C48 VTAIL.n1 VSUBS 0.023238f
C49 VTAIL.n2 VSUBS 0.012487f
C50 VTAIL.n3 VSUBS 0.029515f
C51 VTAIL.n4 VSUBS 0.013222f
C52 VTAIL.n5 VSUBS 0.023238f
C53 VTAIL.n6 VSUBS 0.012487f
C54 VTAIL.n7 VSUBS 0.029515f
C55 VTAIL.n8 VSUBS 0.012854f
C56 VTAIL.n9 VSUBS 0.023238f
C57 VTAIL.n10 VSUBS 0.013222f
C58 VTAIL.n11 VSUBS 0.029515f
C59 VTAIL.n12 VSUBS 0.013222f
C60 VTAIL.n13 VSUBS 0.023238f
C61 VTAIL.n14 VSUBS 0.012487f
C62 VTAIL.n15 VSUBS 0.029515f
C63 VTAIL.n16 VSUBS 0.013222f
C64 VTAIL.n17 VSUBS 1.09187f
C65 VTAIL.n18 VSUBS 0.012487f
C66 VTAIL.t3 VSUBS 0.063569f
C67 VTAIL.n19 VSUBS 0.177871f
C68 VTAIL.n20 VSUBS 0.022203f
C69 VTAIL.n21 VSUBS 0.022136f
C70 VTAIL.n22 VSUBS 0.029515f
C71 VTAIL.n23 VSUBS 0.013222f
C72 VTAIL.n24 VSUBS 0.012487f
C73 VTAIL.n25 VSUBS 0.023238f
C74 VTAIL.n26 VSUBS 0.023238f
C75 VTAIL.n27 VSUBS 0.012487f
C76 VTAIL.n28 VSUBS 0.013222f
C77 VTAIL.n29 VSUBS 0.029515f
C78 VTAIL.n30 VSUBS 0.029515f
C79 VTAIL.n31 VSUBS 0.013222f
C80 VTAIL.n32 VSUBS 0.012487f
C81 VTAIL.n33 VSUBS 0.023238f
C82 VTAIL.n34 VSUBS 0.023238f
C83 VTAIL.n35 VSUBS 0.012487f
C84 VTAIL.n36 VSUBS 0.012487f
C85 VTAIL.n37 VSUBS 0.013222f
C86 VTAIL.n38 VSUBS 0.029515f
C87 VTAIL.n39 VSUBS 0.029515f
C88 VTAIL.n40 VSUBS 0.029515f
C89 VTAIL.n41 VSUBS 0.012854f
C90 VTAIL.n42 VSUBS 0.012487f
C91 VTAIL.n43 VSUBS 0.023238f
C92 VTAIL.n44 VSUBS 0.023238f
C93 VTAIL.n45 VSUBS 0.012487f
C94 VTAIL.n46 VSUBS 0.013222f
C95 VTAIL.n47 VSUBS 0.029515f
C96 VTAIL.n48 VSUBS 0.029515f
C97 VTAIL.n49 VSUBS 0.013222f
C98 VTAIL.n50 VSUBS 0.012487f
C99 VTAIL.n51 VSUBS 0.023238f
C100 VTAIL.n52 VSUBS 0.023238f
C101 VTAIL.n53 VSUBS 0.012487f
C102 VTAIL.n54 VSUBS 0.013222f
C103 VTAIL.n55 VSUBS 0.029515f
C104 VTAIL.n56 VSUBS 0.073471f
C105 VTAIL.n57 VSUBS 0.013222f
C106 VTAIL.n58 VSUBS 0.012487f
C107 VTAIL.n59 VSUBS 0.057206f
C108 VTAIL.n60 VSUBS 0.037142f
C109 VTAIL.n61 VSUBS 0.128168f
C110 VTAIL.n62 VSUBS 0.026126f
C111 VTAIL.n63 VSUBS 0.023238f
C112 VTAIL.n64 VSUBS 0.012487f
C113 VTAIL.n65 VSUBS 0.029515f
C114 VTAIL.n66 VSUBS 0.013222f
C115 VTAIL.n67 VSUBS 0.023238f
C116 VTAIL.n68 VSUBS 0.012487f
C117 VTAIL.n69 VSUBS 0.029515f
C118 VTAIL.n70 VSUBS 0.012854f
C119 VTAIL.n71 VSUBS 0.023238f
C120 VTAIL.n72 VSUBS 0.013222f
C121 VTAIL.n73 VSUBS 0.029515f
C122 VTAIL.n74 VSUBS 0.013222f
C123 VTAIL.n75 VSUBS 0.023238f
C124 VTAIL.n76 VSUBS 0.012487f
C125 VTAIL.n77 VSUBS 0.029515f
C126 VTAIL.n78 VSUBS 0.013222f
C127 VTAIL.n79 VSUBS 1.09187f
C128 VTAIL.n80 VSUBS 0.012487f
C129 VTAIL.t5 VSUBS 0.063569f
C130 VTAIL.n81 VSUBS 0.177871f
C131 VTAIL.n82 VSUBS 0.022203f
C132 VTAIL.n83 VSUBS 0.022136f
C133 VTAIL.n84 VSUBS 0.029515f
C134 VTAIL.n85 VSUBS 0.013222f
C135 VTAIL.n86 VSUBS 0.012487f
C136 VTAIL.n87 VSUBS 0.023238f
C137 VTAIL.n88 VSUBS 0.023238f
C138 VTAIL.n89 VSUBS 0.012487f
C139 VTAIL.n90 VSUBS 0.013222f
C140 VTAIL.n91 VSUBS 0.029515f
C141 VTAIL.n92 VSUBS 0.029515f
C142 VTAIL.n93 VSUBS 0.013222f
C143 VTAIL.n94 VSUBS 0.012487f
C144 VTAIL.n95 VSUBS 0.023238f
C145 VTAIL.n96 VSUBS 0.023238f
C146 VTAIL.n97 VSUBS 0.012487f
C147 VTAIL.n98 VSUBS 0.012487f
C148 VTAIL.n99 VSUBS 0.013222f
C149 VTAIL.n100 VSUBS 0.029515f
C150 VTAIL.n101 VSUBS 0.029515f
C151 VTAIL.n102 VSUBS 0.029515f
C152 VTAIL.n103 VSUBS 0.012854f
C153 VTAIL.n104 VSUBS 0.012487f
C154 VTAIL.n105 VSUBS 0.023238f
C155 VTAIL.n106 VSUBS 0.023238f
C156 VTAIL.n107 VSUBS 0.012487f
C157 VTAIL.n108 VSUBS 0.013222f
C158 VTAIL.n109 VSUBS 0.029515f
C159 VTAIL.n110 VSUBS 0.029515f
C160 VTAIL.n111 VSUBS 0.013222f
C161 VTAIL.n112 VSUBS 0.012487f
C162 VTAIL.n113 VSUBS 0.023238f
C163 VTAIL.n114 VSUBS 0.023238f
C164 VTAIL.n115 VSUBS 0.012487f
C165 VTAIL.n116 VSUBS 0.013222f
C166 VTAIL.n117 VSUBS 0.029515f
C167 VTAIL.n118 VSUBS 0.073471f
C168 VTAIL.n119 VSUBS 0.013222f
C169 VTAIL.n120 VSUBS 0.012487f
C170 VTAIL.n121 VSUBS 0.057206f
C171 VTAIL.n122 VSUBS 0.037142f
C172 VTAIL.n123 VSUBS 0.190621f
C173 VTAIL.n124 VSUBS 0.026126f
C174 VTAIL.n125 VSUBS 0.023238f
C175 VTAIL.n126 VSUBS 0.012487f
C176 VTAIL.n127 VSUBS 0.029515f
C177 VTAIL.n128 VSUBS 0.013222f
C178 VTAIL.n129 VSUBS 0.023238f
C179 VTAIL.n130 VSUBS 0.012487f
C180 VTAIL.n131 VSUBS 0.029515f
C181 VTAIL.n132 VSUBS 0.012854f
C182 VTAIL.n133 VSUBS 0.023238f
C183 VTAIL.n134 VSUBS 0.013222f
C184 VTAIL.n135 VSUBS 0.029515f
C185 VTAIL.n136 VSUBS 0.013222f
C186 VTAIL.n137 VSUBS 0.023238f
C187 VTAIL.n138 VSUBS 0.012487f
C188 VTAIL.n139 VSUBS 0.029515f
C189 VTAIL.n140 VSUBS 0.013222f
C190 VTAIL.n141 VSUBS 1.09187f
C191 VTAIL.n142 VSUBS 0.012487f
C192 VTAIL.t7 VSUBS 0.063569f
C193 VTAIL.n143 VSUBS 0.177871f
C194 VTAIL.n144 VSUBS 0.022203f
C195 VTAIL.n145 VSUBS 0.022136f
C196 VTAIL.n146 VSUBS 0.029515f
C197 VTAIL.n147 VSUBS 0.013222f
C198 VTAIL.n148 VSUBS 0.012487f
C199 VTAIL.n149 VSUBS 0.023238f
C200 VTAIL.n150 VSUBS 0.023238f
C201 VTAIL.n151 VSUBS 0.012487f
C202 VTAIL.n152 VSUBS 0.013222f
C203 VTAIL.n153 VSUBS 0.029515f
C204 VTAIL.n154 VSUBS 0.029515f
C205 VTAIL.n155 VSUBS 0.013222f
C206 VTAIL.n156 VSUBS 0.012487f
C207 VTAIL.n157 VSUBS 0.023238f
C208 VTAIL.n158 VSUBS 0.023238f
C209 VTAIL.n159 VSUBS 0.012487f
C210 VTAIL.n160 VSUBS 0.012487f
C211 VTAIL.n161 VSUBS 0.013222f
C212 VTAIL.n162 VSUBS 0.029515f
C213 VTAIL.n163 VSUBS 0.029515f
C214 VTAIL.n164 VSUBS 0.029515f
C215 VTAIL.n165 VSUBS 0.012854f
C216 VTAIL.n166 VSUBS 0.012487f
C217 VTAIL.n167 VSUBS 0.023238f
C218 VTAIL.n168 VSUBS 0.023238f
C219 VTAIL.n169 VSUBS 0.012487f
C220 VTAIL.n170 VSUBS 0.013222f
C221 VTAIL.n171 VSUBS 0.029515f
C222 VTAIL.n172 VSUBS 0.029515f
C223 VTAIL.n173 VSUBS 0.013222f
C224 VTAIL.n174 VSUBS 0.012487f
C225 VTAIL.n175 VSUBS 0.023238f
C226 VTAIL.n176 VSUBS 0.023238f
C227 VTAIL.n177 VSUBS 0.012487f
C228 VTAIL.n178 VSUBS 0.013222f
C229 VTAIL.n179 VSUBS 0.029515f
C230 VTAIL.n180 VSUBS 0.073471f
C231 VTAIL.n181 VSUBS 0.013222f
C232 VTAIL.n182 VSUBS 0.012487f
C233 VTAIL.n183 VSUBS 0.057206f
C234 VTAIL.n184 VSUBS 0.037142f
C235 VTAIL.n185 VSUBS 1.3477f
C236 VTAIL.n186 VSUBS 0.026126f
C237 VTAIL.n187 VSUBS 0.023238f
C238 VTAIL.n188 VSUBS 0.012487f
C239 VTAIL.n189 VSUBS 0.029515f
C240 VTAIL.n190 VSUBS 0.013222f
C241 VTAIL.n191 VSUBS 0.023238f
C242 VTAIL.n192 VSUBS 0.012487f
C243 VTAIL.n193 VSUBS 0.029515f
C244 VTAIL.n194 VSUBS 0.012854f
C245 VTAIL.n195 VSUBS 0.023238f
C246 VTAIL.n196 VSUBS 0.012854f
C247 VTAIL.n197 VSUBS 0.012487f
C248 VTAIL.n198 VSUBS 0.029515f
C249 VTAIL.n199 VSUBS 0.029515f
C250 VTAIL.n200 VSUBS 0.013222f
C251 VTAIL.n201 VSUBS 0.023238f
C252 VTAIL.n202 VSUBS 0.012487f
C253 VTAIL.n203 VSUBS 0.029515f
C254 VTAIL.n204 VSUBS 0.013222f
C255 VTAIL.n205 VSUBS 1.09187f
C256 VTAIL.n206 VSUBS 0.012487f
C257 VTAIL.t0 VSUBS 0.063569f
C258 VTAIL.n207 VSUBS 0.177871f
C259 VTAIL.n208 VSUBS 0.022203f
C260 VTAIL.n209 VSUBS 0.022136f
C261 VTAIL.n210 VSUBS 0.029515f
C262 VTAIL.n211 VSUBS 0.013222f
C263 VTAIL.n212 VSUBS 0.012487f
C264 VTAIL.n213 VSUBS 0.023238f
C265 VTAIL.n214 VSUBS 0.023238f
C266 VTAIL.n215 VSUBS 0.012487f
C267 VTAIL.n216 VSUBS 0.013222f
C268 VTAIL.n217 VSUBS 0.029515f
C269 VTAIL.n218 VSUBS 0.029515f
C270 VTAIL.n219 VSUBS 0.013222f
C271 VTAIL.n220 VSUBS 0.012487f
C272 VTAIL.n221 VSUBS 0.023238f
C273 VTAIL.n222 VSUBS 0.023238f
C274 VTAIL.n223 VSUBS 0.012487f
C275 VTAIL.n224 VSUBS 0.013222f
C276 VTAIL.n225 VSUBS 0.029515f
C277 VTAIL.n226 VSUBS 0.029515f
C278 VTAIL.n227 VSUBS 0.013222f
C279 VTAIL.n228 VSUBS 0.012487f
C280 VTAIL.n229 VSUBS 0.023238f
C281 VTAIL.n230 VSUBS 0.023238f
C282 VTAIL.n231 VSUBS 0.012487f
C283 VTAIL.n232 VSUBS 0.013222f
C284 VTAIL.n233 VSUBS 0.029515f
C285 VTAIL.n234 VSUBS 0.029515f
C286 VTAIL.n235 VSUBS 0.013222f
C287 VTAIL.n236 VSUBS 0.012487f
C288 VTAIL.n237 VSUBS 0.023238f
C289 VTAIL.n238 VSUBS 0.023238f
C290 VTAIL.n239 VSUBS 0.012487f
C291 VTAIL.n240 VSUBS 0.013222f
C292 VTAIL.n241 VSUBS 0.029515f
C293 VTAIL.n242 VSUBS 0.073471f
C294 VTAIL.n243 VSUBS 0.013222f
C295 VTAIL.n244 VSUBS 0.012487f
C296 VTAIL.n245 VSUBS 0.057206f
C297 VTAIL.n246 VSUBS 0.037142f
C298 VTAIL.n247 VSUBS 1.3477f
C299 VTAIL.n248 VSUBS 0.026126f
C300 VTAIL.n249 VSUBS 0.023238f
C301 VTAIL.n250 VSUBS 0.012487f
C302 VTAIL.n251 VSUBS 0.029515f
C303 VTAIL.n252 VSUBS 0.013222f
C304 VTAIL.n253 VSUBS 0.023238f
C305 VTAIL.n254 VSUBS 0.012487f
C306 VTAIL.n255 VSUBS 0.029515f
C307 VTAIL.n256 VSUBS 0.012854f
C308 VTAIL.n257 VSUBS 0.023238f
C309 VTAIL.n258 VSUBS 0.012854f
C310 VTAIL.n259 VSUBS 0.012487f
C311 VTAIL.n260 VSUBS 0.029515f
C312 VTAIL.n261 VSUBS 0.029515f
C313 VTAIL.n262 VSUBS 0.013222f
C314 VTAIL.n263 VSUBS 0.023238f
C315 VTAIL.n264 VSUBS 0.012487f
C316 VTAIL.n265 VSUBS 0.029515f
C317 VTAIL.n266 VSUBS 0.013222f
C318 VTAIL.n267 VSUBS 1.09187f
C319 VTAIL.n268 VSUBS 0.012487f
C320 VTAIL.t2 VSUBS 0.063569f
C321 VTAIL.n269 VSUBS 0.177871f
C322 VTAIL.n270 VSUBS 0.022203f
C323 VTAIL.n271 VSUBS 0.022136f
C324 VTAIL.n272 VSUBS 0.029515f
C325 VTAIL.n273 VSUBS 0.013222f
C326 VTAIL.n274 VSUBS 0.012487f
C327 VTAIL.n275 VSUBS 0.023238f
C328 VTAIL.n276 VSUBS 0.023238f
C329 VTAIL.n277 VSUBS 0.012487f
C330 VTAIL.n278 VSUBS 0.013222f
C331 VTAIL.n279 VSUBS 0.029515f
C332 VTAIL.n280 VSUBS 0.029515f
C333 VTAIL.n281 VSUBS 0.013222f
C334 VTAIL.n282 VSUBS 0.012487f
C335 VTAIL.n283 VSUBS 0.023238f
C336 VTAIL.n284 VSUBS 0.023238f
C337 VTAIL.n285 VSUBS 0.012487f
C338 VTAIL.n286 VSUBS 0.013222f
C339 VTAIL.n287 VSUBS 0.029515f
C340 VTAIL.n288 VSUBS 0.029515f
C341 VTAIL.n289 VSUBS 0.013222f
C342 VTAIL.n290 VSUBS 0.012487f
C343 VTAIL.n291 VSUBS 0.023238f
C344 VTAIL.n292 VSUBS 0.023238f
C345 VTAIL.n293 VSUBS 0.012487f
C346 VTAIL.n294 VSUBS 0.013222f
C347 VTAIL.n295 VSUBS 0.029515f
C348 VTAIL.n296 VSUBS 0.029515f
C349 VTAIL.n297 VSUBS 0.013222f
C350 VTAIL.n298 VSUBS 0.012487f
C351 VTAIL.n299 VSUBS 0.023238f
C352 VTAIL.n300 VSUBS 0.023238f
C353 VTAIL.n301 VSUBS 0.012487f
C354 VTAIL.n302 VSUBS 0.013222f
C355 VTAIL.n303 VSUBS 0.029515f
C356 VTAIL.n304 VSUBS 0.073471f
C357 VTAIL.n305 VSUBS 0.013222f
C358 VTAIL.n306 VSUBS 0.012487f
C359 VTAIL.n307 VSUBS 0.057206f
C360 VTAIL.n308 VSUBS 0.037142f
C361 VTAIL.n309 VSUBS 0.190621f
C362 VTAIL.n310 VSUBS 0.026126f
C363 VTAIL.n311 VSUBS 0.023238f
C364 VTAIL.n312 VSUBS 0.012487f
C365 VTAIL.n313 VSUBS 0.029515f
C366 VTAIL.n314 VSUBS 0.013222f
C367 VTAIL.n315 VSUBS 0.023238f
C368 VTAIL.n316 VSUBS 0.012487f
C369 VTAIL.n317 VSUBS 0.029515f
C370 VTAIL.n318 VSUBS 0.012854f
C371 VTAIL.n319 VSUBS 0.023238f
C372 VTAIL.n320 VSUBS 0.012854f
C373 VTAIL.n321 VSUBS 0.012487f
C374 VTAIL.n322 VSUBS 0.029515f
C375 VTAIL.n323 VSUBS 0.029515f
C376 VTAIL.n324 VSUBS 0.013222f
C377 VTAIL.n325 VSUBS 0.023238f
C378 VTAIL.n326 VSUBS 0.012487f
C379 VTAIL.n327 VSUBS 0.029515f
C380 VTAIL.n328 VSUBS 0.013222f
C381 VTAIL.n329 VSUBS 1.09187f
C382 VTAIL.n330 VSUBS 0.012487f
C383 VTAIL.t4 VSUBS 0.063569f
C384 VTAIL.n331 VSUBS 0.177871f
C385 VTAIL.n332 VSUBS 0.022203f
C386 VTAIL.n333 VSUBS 0.022136f
C387 VTAIL.n334 VSUBS 0.029515f
C388 VTAIL.n335 VSUBS 0.013222f
C389 VTAIL.n336 VSUBS 0.012487f
C390 VTAIL.n337 VSUBS 0.023238f
C391 VTAIL.n338 VSUBS 0.023238f
C392 VTAIL.n339 VSUBS 0.012487f
C393 VTAIL.n340 VSUBS 0.013222f
C394 VTAIL.n341 VSUBS 0.029515f
C395 VTAIL.n342 VSUBS 0.029515f
C396 VTAIL.n343 VSUBS 0.013222f
C397 VTAIL.n344 VSUBS 0.012487f
C398 VTAIL.n345 VSUBS 0.023238f
C399 VTAIL.n346 VSUBS 0.023238f
C400 VTAIL.n347 VSUBS 0.012487f
C401 VTAIL.n348 VSUBS 0.013222f
C402 VTAIL.n349 VSUBS 0.029515f
C403 VTAIL.n350 VSUBS 0.029515f
C404 VTAIL.n351 VSUBS 0.013222f
C405 VTAIL.n352 VSUBS 0.012487f
C406 VTAIL.n353 VSUBS 0.023238f
C407 VTAIL.n354 VSUBS 0.023238f
C408 VTAIL.n355 VSUBS 0.012487f
C409 VTAIL.n356 VSUBS 0.013222f
C410 VTAIL.n357 VSUBS 0.029515f
C411 VTAIL.n358 VSUBS 0.029515f
C412 VTAIL.n359 VSUBS 0.013222f
C413 VTAIL.n360 VSUBS 0.012487f
C414 VTAIL.n361 VSUBS 0.023238f
C415 VTAIL.n362 VSUBS 0.023238f
C416 VTAIL.n363 VSUBS 0.012487f
C417 VTAIL.n364 VSUBS 0.013222f
C418 VTAIL.n365 VSUBS 0.029515f
C419 VTAIL.n366 VSUBS 0.073471f
C420 VTAIL.n367 VSUBS 0.013222f
C421 VTAIL.n368 VSUBS 0.012487f
C422 VTAIL.n369 VSUBS 0.057206f
C423 VTAIL.n370 VSUBS 0.037142f
C424 VTAIL.n371 VSUBS 0.190621f
C425 VTAIL.n372 VSUBS 0.026126f
C426 VTAIL.n373 VSUBS 0.023238f
C427 VTAIL.n374 VSUBS 0.012487f
C428 VTAIL.n375 VSUBS 0.029515f
C429 VTAIL.n376 VSUBS 0.013222f
C430 VTAIL.n377 VSUBS 0.023238f
C431 VTAIL.n378 VSUBS 0.012487f
C432 VTAIL.n379 VSUBS 0.029515f
C433 VTAIL.n380 VSUBS 0.012854f
C434 VTAIL.n381 VSUBS 0.023238f
C435 VTAIL.n382 VSUBS 0.012854f
C436 VTAIL.n383 VSUBS 0.012487f
C437 VTAIL.n384 VSUBS 0.029515f
C438 VTAIL.n385 VSUBS 0.029515f
C439 VTAIL.n386 VSUBS 0.013222f
C440 VTAIL.n387 VSUBS 0.023238f
C441 VTAIL.n388 VSUBS 0.012487f
C442 VTAIL.n389 VSUBS 0.029515f
C443 VTAIL.n390 VSUBS 0.013222f
C444 VTAIL.n391 VSUBS 1.09187f
C445 VTAIL.n392 VSUBS 0.012487f
C446 VTAIL.t6 VSUBS 0.063569f
C447 VTAIL.n393 VSUBS 0.177871f
C448 VTAIL.n394 VSUBS 0.022203f
C449 VTAIL.n395 VSUBS 0.022136f
C450 VTAIL.n396 VSUBS 0.029515f
C451 VTAIL.n397 VSUBS 0.013222f
C452 VTAIL.n398 VSUBS 0.012487f
C453 VTAIL.n399 VSUBS 0.023238f
C454 VTAIL.n400 VSUBS 0.023238f
C455 VTAIL.n401 VSUBS 0.012487f
C456 VTAIL.n402 VSUBS 0.013222f
C457 VTAIL.n403 VSUBS 0.029515f
C458 VTAIL.n404 VSUBS 0.029515f
C459 VTAIL.n405 VSUBS 0.013222f
C460 VTAIL.n406 VSUBS 0.012487f
C461 VTAIL.n407 VSUBS 0.023238f
C462 VTAIL.n408 VSUBS 0.023238f
C463 VTAIL.n409 VSUBS 0.012487f
C464 VTAIL.n410 VSUBS 0.013222f
C465 VTAIL.n411 VSUBS 0.029515f
C466 VTAIL.n412 VSUBS 0.029515f
C467 VTAIL.n413 VSUBS 0.013222f
C468 VTAIL.n414 VSUBS 0.012487f
C469 VTAIL.n415 VSUBS 0.023238f
C470 VTAIL.n416 VSUBS 0.023238f
C471 VTAIL.n417 VSUBS 0.012487f
C472 VTAIL.n418 VSUBS 0.013222f
C473 VTAIL.n419 VSUBS 0.029515f
C474 VTAIL.n420 VSUBS 0.029515f
C475 VTAIL.n421 VSUBS 0.013222f
C476 VTAIL.n422 VSUBS 0.012487f
C477 VTAIL.n423 VSUBS 0.023238f
C478 VTAIL.n424 VSUBS 0.023238f
C479 VTAIL.n425 VSUBS 0.012487f
C480 VTAIL.n426 VSUBS 0.013222f
C481 VTAIL.n427 VSUBS 0.029515f
C482 VTAIL.n428 VSUBS 0.073471f
C483 VTAIL.n429 VSUBS 0.013222f
C484 VTAIL.n430 VSUBS 0.012487f
C485 VTAIL.n431 VSUBS 0.057206f
C486 VTAIL.n432 VSUBS 0.037142f
C487 VTAIL.n433 VSUBS 1.3477f
C488 VTAIL.n434 VSUBS 0.026126f
C489 VTAIL.n435 VSUBS 0.023238f
C490 VTAIL.n436 VSUBS 0.012487f
C491 VTAIL.n437 VSUBS 0.029515f
C492 VTAIL.n438 VSUBS 0.013222f
C493 VTAIL.n439 VSUBS 0.023238f
C494 VTAIL.n440 VSUBS 0.012487f
C495 VTAIL.n441 VSUBS 0.029515f
C496 VTAIL.n442 VSUBS 0.012854f
C497 VTAIL.n443 VSUBS 0.023238f
C498 VTAIL.n444 VSUBS 0.013222f
C499 VTAIL.n445 VSUBS 0.029515f
C500 VTAIL.n446 VSUBS 0.013222f
C501 VTAIL.n447 VSUBS 0.023238f
C502 VTAIL.n448 VSUBS 0.012487f
C503 VTAIL.n449 VSUBS 0.029515f
C504 VTAIL.n450 VSUBS 0.013222f
C505 VTAIL.n451 VSUBS 1.09187f
C506 VTAIL.n452 VSUBS 0.012487f
C507 VTAIL.t1 VSUBS 0.063569f
C508 VTAIL.n453 VSUBS 0.177871f
C509 VTAIL.n454 VSUBS 0.022203f
C510 VTAIL.n455 VSUBS 0.022136f
C511 VTAIL.n456 VSUBS 0.029515f
C512 VTAIL.n457 VSUBS 0.013222f
C513 VTAIL.n458 VSUBS 0.012487f
C514 VTAIL.n459 VSUBS 0.023238f
C515 VTAIL.n460 VSUBS 0.023238f
C516 VTAIL.n461 VSUBS 0.012487f
C517 VTAIL.n462 VSUBS 0.013222f
C518 VTAIL.n463 VSUBS 0.029515f
C519 VTAIL.n464 VSUBS 0.029515f
C520 VTAIL.n465 VSUBS 0.013222f
C521 VTAIL.n466 VSUBS 0.012487f
C522 VTAIL.n467 VSUBS 0.023238f
C523 VTAIL.n468 VSUBS 0.023238f
C524 VTAIL.n469 VSUBS 0.012487f
C525 VTAIL.n470 VSUBS 0.012487f
C526 VTAIL.n471 VSUBS 0.013222f
C527 VTAIL.n472 VSUBS 0.029515f
C528 VTAIL.n473 VSUBS 0.029515f
C529 VTAIL.n474 VSUBS 0.029515f
C530 VTAIL.n475 VSUBS 0.012854f
C531 VTAIL.n476 VSUBS 0.012487f
C532 VTAIL.n477 VSUBS 0.023238f
C533 VTAIL.n478 VSUBS 0.023238f
C534 VTAIL.n479 VSUBS 0.012487f
C535 VTAIL.n480 VSUBS 0.013222f
C536 VTAIL.n481 VSUBS 0.029515f
C537 VTAIL.n482 VSUBS 0.029515f
C538 VTAIL.n483 VSUBS 0.013222f
C539 VTAIL.n484 VSUBS 0.012487f
C540 VTAIL.n485 VSUBS 0.023238f
C541 VTAIL.n486 VSUBS 0.023238f
C542 VTAIL.n487 VSUBS 0.012487f
C543 VTAIL.n488 VSUBS 0.013222f
C544 VTAIL.n489 VSUBS 0.029515f
C545 VTAIL.n490 VSUBS 0.073471f
C546 VTAIL.n491 VSUBS 0.013222f
C547 VTAIL.n492 VSUBS 0.012487f
C548 VTAIL.n493 VSUBS 0.057206f
C549 VTAIL.n494 VSUBS 0.037142f
C550 VTAIL.n495 VSUBS 1.27654f
C551 VP.n0 VSUBS 0.042446f
C552 VP.t1 VSUBS 2.31332f
C553 VP.n1 VSUBS 0.034313f
C554 VP.n2 VSUBS 0.042446f
C555 VP.t3 VSUBS 2.31332f
C556 VP.t2 VSUBS 2.5022f
C557 VP.t0 VSUBS 2.49992f
C558 VP.n3 VSUBS 3.5018f
C559 VP.n4 VSUBS 2.26301f
C560 VP.n5 VSUBS 0.921307f
C561 VP.n6 VSUBS 0.042784f
C562 VP.n7 VSUBS 0.08436f
C563 VP.n8 VSUBS 0.042446f
C564 VP.n9 VSUBS 0.042446f
C565 VP.n10 VSUBS 0.042446f
C566 VP.n11 VSUBS 0.08436f
C567 VP.n12 VSUBS 0.042784f
C568 VP.n13 VSUBS 0.921307f
C569 VP.n14 VSUBS 0.045329f
C570 B.n0 VSUBS 0.00652f
C571 B.n1 VSUBS 0.00652f
C572 B.n2 VSUBS 0.009643f
C573 B.n3 VSUBS 0.007389f
C574 B.n4 VSUBS 0.007389f
C575 B.n5 VSUBS 0.007389f
C576 B.n6 VSUBS 0.007389f
C577 B.n7 VSUBS 0.007389f
C578 B.n8 VSUBS 0.007389f
C579 B.n9 VSUBS 0.007389f
C580 B.n10 VSUBS 0.007389f
C581 B.n11 VSUBS 0.007389f
C582 B.n12 VSUBS 0.007389f
C583 B.n13 VSUBS 0.007389f
C584 B.n14 VSUBS 0.007389f
C585 B.n15 VSUBS 0.016999f
C586 B.n16 VSUBS 0.007389f
C587 B.n17 VSUBS 0.007389f
C588 B.n18 VSUBS 0.007389f
C589 B.n19 VSUBS 0.007389f
C590 B.n20 VSUBS 0.007389f
C591 B.n21 VSUBS 0.007389f
C592 B.n22 VSUBS 0.007389f
C593 B.n23 VSUBS 0.007389f
C594 B.n24 VSUBS 0.007389f
C595 B.n25 VSUBS 0.007389f
C596 B.n26 VSUBS 0.007389f
C597 B.n27 VSUBS 0.007389f
C598 B.n28 VSUBS 0.007389f
C599 B.n29 VSUBS 0.007389f
C600 B.n30 VSUBS 0.007389f
C601 B.n31 VSUBS 0.007389f
C602 B.n32 VSUBS 0.007389f
C603 B.n33 VSUBS 0.007389f
C604 B.n34 VSUBS 0.007389f
C605 B.n35 VSUBS 0.007389f
C606 B.t7 VSUBS 0.211509f
C607 B.t8 VSUBS 0.235579f
C608 B.t6 VSUBS 0.938037f
C609 B.n36 VSUBS 0.367486f
C610 B.n37 VSUBS 0.254634f
C611 B.n38 VSUBS 0.007389f
C612 B.n39 VSUBS 0.007389f
C613 B.n40 VSUBS 0.007389f
C614 B.n41 VSUBS 0.007389f
C615 B.t1 VSUBS 0.211512f
C616 B.t2 VSUBS 0.235582f
C617 B.t0 VSUBS 0.938037f
C618 B.n42 VSUBS 0.367483f
C619 B.n43 VSUBS 0.254631f
C620 B.n44 VSUBS 0.01712f
C621 B.n45 VSUBS 0.007389f
C622 B.n46 VSUBS 0.007389f
C623 B.n47 VSUBS 0.007389f
C624 B.n48 VSUBS 0.007389f
C625 B.n49 VSUBS 0.007389f
C626 B.n50 VSUBS 0.007389f
C627 B.n51 VSUBS 0.007389f
C628 B.n52 VSUBS 0.007389f
C629 B.n53 VSUBS 0.007389f
C630 B.n54 VSUBS 0.007389f
C631 B.n55 VSUBS 0.007389f
C632 B.n56 VSUBS 0.007389f
C633 B.n57 VSUBS 0.007389f
C634 B.n58 VSUBS 0.007389f
C635 B.n59 VSUBS 0.007389f
C636 B.n60 VSUBS 0.007389f
C637 B.n61 VSUBS 0.007389f
C638 B.n62 VSUBS 0.007389f
C639 B.n63 VSUBS 0.007389f
C640 B.n64 VSUBS 0.016999f
C641 B.n65 VSUBS 0.007389f
C642 B.n66 VSUBS 0.007389f
C643 B.n67 VSUBS 0.007389f
C644 B.n68 VSUBS 0.007389f
C645 B.n69 VSUBS 0.007389f
C646 B.n70 VSUBS 0.007389f
C647 B.n71 VSUBS 0.007389f
C648 B.n72 VSUBS 0.007389f
C649 B.n73 VSUBS 0.007389f
C650 B.n74 VSUBS 0.007389f
C651 B.n75 VSUBS 0.007389f
C652 B.n76 VSUBS 0.007389f
C653 B.n77 VSUBS 0.007389f
C654 B.n78 VSUBS 0.007389f
C655 B.n79 VSUBS 0.007389f
C656 B.n80 VSUBS 0.007389f
C657 B.n81 VSUBS 0.007389f
C658 B.n82 VSUBS 0.007389f
C659 B.n83 VSUBS 0.007389f
C660 B.n84 VSUBS 0.007389f
C661 B.n85 VSUBS 0.007389f
C662 B.n86 VSUBS 0.007389f
C663 B.n87 VSUBS 0.007389f
C664 B.n88 VSUBS 0.007389f
C665 B.n89 VSUBS 0.007389f
C666 B.n90 VSUBS 0.007389f
C667 B.n91 VSUBS 0.016253f
C668 B.n92 VSUBS 0.007389f
C669 B.n93 VSUBS 0.007389f
C670 B.n94 VSUBS 0.007389f
C671 B.n95 VSUBS 0.007389f
C672 B.n96 VSUBS 0.007389f
C673 B.n97 VSUBS 0.007389f
C674 B.n98 VSUBS 0.007389f
C675 B.n99 VSUBS 0.007389f
C676 B.n100 VSUBS 0.007389f
C677 B.n101 VSUBS 0.007389f
C678 B.n102 VSUBS 0.007389f
C679 B.n103 VSUBS 0.007389f
C680 B.n104 VSUBS 0.007389f
C681 B.n105 VSUBS 0.007389f
C682 B.n106 VSUBS 0.007389f
C683 B.n107 VSUBS 0.007389f
C684 B.n108 VSUBS 0.007389f
C685 B.n109 VSUBS 0.007389f
C686 B.n110 VSUBS 0.007389f
C687 B.n111 VSUBS 0.007389f
C688 B.t5 VSUBS 0.211512f
C689 B.t4 VSUBS 0.235582f
C690 B.t3 VSUBS 0.938037f
C691 B.n112 VSUBS 0.367483f
C692 B.n113 VSUBS 0.254631f
C693 B.n114 VSUBS 0.007389f
C694 B.n115 VSUBS 0.007389f
C695 B.n116 VSUBS 0.007389f
C696 B.n117 VSUBS 0.007389f
C697 B.n118 VSUBS 0.004129f
C698 B.n119 VSUBS 0.007389f
C699 B.n120 VSUBS 0.007389f
C700 B.n121 VSUBS 0.007389f
C701 B.n122 VSUBS 0.007389f
C702 B.n123 VSUBS 0.007389f
C703 B.n124 VSUBS 0.007389f
C704 B.n125 VSUBS 0.007389f
C705 B.n126 VSUBS 0.007389f
C706 B.n127 VSUBS 0.007389f
C707 B.n128 VSUBS 0.007389f
C708 B.n129 VSUBS 0.007389f
C709 B.n130 VSUBS 0.007389f
C710 B.n131 VSUBS 0.007389f
C711 B.n132 VSUBS 0.007389f
C712 B.n133 VSUBS 0.007389f
C713 B.n134 VSUBS 0.007389f
C714 B.n135 VSUBS 0.007389f
C715 B.n136 VSUBS 0.007389f
C716 B.n137 VSUBS 0.007389f
C717 B.n138 VSUBS 0.016999f
C718 B.n139 VSUBS 0.007389f
C719 B.n140 VSUBS 0.007389f
C720 B.n141 VSUBS 0.007389f
C721 B.n142 VSUBS 0.007389f
C722 B.n143 VSUBS 0.007389f
C723 B.n144 VSUBS 0.007389f
C724 B.n145 VSUBS 0.007389f
C725 B.n146 VSUBS 0.007389f
C726 B.n147 VSUBS 0.007389f
C727 B.n148 VSUBS 0.007389f
C728 B.n149 VSUBS 0.007389f
C729 B.n150 VSUBS 0.007389f
C730 B.n151 VSUBS 0.007389f
C731 B.n152 VSUBS 0.007389f
C732 B.n153 VSUBS 0.007389f
C733 B.n154 VSUBS 0.007389f
C734 B.n155 VSUBS 0.007389f
C735 B.n156 VSUBS 0.007389f
C736 B.n157 VSUBS 0.007389f
C737 B.n158 VSUBS 0.007389f
C738 B.n159 VSUBS 0.007389f
C739 B.n160 VSUBS 0.007389f
C740 B.n161 VSUBS 0.007389f
C741 B.n162 VSUBS 0.007389f
C742 B.n163 VSUBS 0.007389f
C743 B.n164 VSUBS 0.007389f
C744 B.n165 VSUBS 0.007389f
C745 B.n166 VSUBS 0.007389f
C746 B.n167 VSUBS 0.007389f
C747 B.n168 VSUBS 0.007389f
C748 B.n169 VSUBS 0.007389f
C749 B.n170 VSUBS 0.007389f
C750 B.n171 VSUBS 0.007389f
C751 B.n172 VSUBS 0.007389f
C752 B.n173 VSUBS 0.007389f
C753 B.n174 VSUBS 0.007389f
C754 B.n175 VSUBS 0.007389f
C755 B.n176 VSUBS 0.007389f
C756 B.n177 VSUBS 0.007389f
C757 B.n178 VSUBS 0.007389f
C758 B.n179 VSUBS 0.007389f
C759 B.n180 VSUBS 0.007389f
C760 B.n181 VSUBS 0.007389f
C761 B.n182 VSUBS 0.007389f
C762 B.n183 VSUBS 0.007389f
C763 B.n184 VSUBS 0.007389f
C764 B.n185 VSUBS 0.007389f
C765 B.n186 VSUBS 0.007389f
C766 B.n187 VSUBS 0.016253f
C767 B.n188 VSUBS 0.016253f
C768 B.n189 VSUBS 0.016999f
C769 B.n190 VSUBS 0.007389f
C770 B.n191 VSUBS 0.007389f
C771 B.n192 VSUBS 0.007389f
C772 B.n193 VSUBS 0.007389f
C773 B.n194 VSUBS 0.007389f
C774 B.n195 VSUBS 0.007389f
C775 B.n196 VSUBS 0.007389f
C776 B.n197 VSUBS 0.007389f
C777 B.n198 VSUBS 0.007389f
C778 B.n199 VSUBS 0.007389f
C779 B.n200 VSUBS 0.007389f
C780 B.n201 VSUBS 0.007389f
C781 B.n202 VSUBS 0.007389f
C782 B.n203 VSUBS 0.007389f
C783 B.n204 VSUBS 0.007389f
C784 B.n205 VSUBS 0.007389f
C785 B.n206 VSUBS 0.007389f
C786 B.n207 VSUBS 0.007389f
C787 B.n208 VSUBS 0.007389f
C788 B.n209 VSUBS 0.007389f
C789 B.n210 VSUBS 0.007389f
C790 B.n211 VSUBS 0.007389f
C791 B.n212 VSUBS 0.007389f
C792 B.n213 VSUBS 0.007389f
C793 B.n214 VSUBS 0.007389f
C794 B.n215 VSUBS 0.007389f
C795 B.n216 VSUBS 0.007389f
C796 B.n217 VSUBS 0.007389f
C797 B.n218 VSUBS 0.007389f
C798 B.n219 VSUBS 0.007389f
C799 B.n220 VSUBS 0.007389f
C800 B.n221 VSUBS 0.007389f
C801 B.n222 VSUBS 0.007389f
C802 B.n223 VSUBS 0.007389f
C803 B.n224 VSUBS 0.007389f
C804 B.n225 VSUBS 0.007389f
C805 B.n226 VSUBS 0.007389f
C806 B.n227 VSUBS 0.007389f
C807 B.n228 VSUBS 0.007389f
C808 B.n229 VSUBS 0.007389f
C809 B.n230 VSUBS 0.007389f
C810 B.n231 VSUBS 0.007389f
C811 B.n232 VSUBS 0.007389f
C812 B.n233 VSUBS 0.007389f
C813 B.n234 VSUBS 0.007389f
C814 B.n235 VSUBS 0.007389f
C815 B.n236 VSUBS 0.007389f
C816 B.n237 VSUBS 0.007389f
C817 B.n238 VSUBS 0.007389f
C818 B.n239 VSUBS 0.007389f
C819 B.n240 VSUBS 0.007389f
C820 B.n241 VSUBS 0.007389f
C821 B.n242 VSUBS 0.007389f
C822 B.n243 VSUBS 0.007389f
C823 B.n244 VSUBS 0.007389f
C824 B.n245 VSUBS 0.007389f
C825 B.n246 VSUBS 0.007389f
C826 B.t11 VSUBS 0.211509f
C827 B.t10 VSUBS 0.235579f
C828 B.t9 VSUBS 0.938037f
C829 B.n247 VSUBS 0.367486f
C830 B.n248 VSUBS 0.254634f
C831 B.n249 VSUBS 0.01712f
C832 B.n250 VSUBS 0.006955f
C833 B.n251 VSUBS 0.007389f
C834 B.n252 VSUBS 0.007389f
C835 B.n253 VSUBS 0.007389f
C836 B.n254 VSUBS 0.007389f
C837 B.n255 VSUBS 0.007389f
C838 B.n256 VSUBS 0.007389f
C839 B.n257 VSUBS 0.007389f
C840 B.n258 VSUBS 0.007389f
C841 B.n259 VSUBS 0.007389f
C842 B.n260 VSUBS 0.007389f
C843 B.n261 VSUBS 0.007389f
C844 B.n262 VSUBS 0.007389f
C845 B.n263 VSUBS 0.007389f
C846 B.n264 VSUBS 0.007389f
C847 B.n265 VSUBS 0.007389f
C848 B.n266 VSUBS 0.004129f
C849 B.n267 VSUBS 0.01712f
C850 B.n268 VSUBS 0.006955f
C851 B.n269 VSUBS 0.007389f
C852 B.n270 VSUBS 0.007389f
C853 B.n271 VSUBS 0.007389f
C854 B.n272 VSUBS 0.007389f
C855 B.n273 VSUBS 0.007389f
C856 B.n274 VSUBS 0.007389f
C857 B.n275 VSUBS 0.007389f
C858 B.n276 VSUBS 0.007389f
C859 B.n277 VSUBS 0.007389f
C860 B.n278 VSUBS 0.007389f
C861 B.n279 VSUBS 0.007389f
C862 B.n280 VSUBS 0.007389f
C863 B.n281 VSUBS 0.007389f
C864 B.n282 VSUBS 0.007389f
C865 B.n283 VSUBS 0.007389f
C866 B.n284 VSUBS 0.007389f
C867 B.n285 VSUBS 0.007389f
C868 B.n286 VSUBS 0.007389f
C869 B.n287 VSUBS 0.007389f
C870 B.n288 VSUBS 0.007389f
C871 B.n289 VSUBS 0.007389f
C872 B.n290 VSUBS 0.007389f
C873 B.n291 VSUBS 0.007389f
C874 B.n292 VSUBS 0.007389f
C875 B.n293 VSUBS 0.007389f
C876 B.n294 VSUBS 0.007389f
C877 B.n295 VSUBS 0.007389f
C878 B.n296 VSUBS 0.007389f
C879 B.n297 VSUBS 0.007389f
C880 B.n298 VSUBS 0.007389f
C881 B.n299 VSUBS 0.007389f
C882 B.n300 VSUBS 0.007389f
C883 B.n301 VSUBS 0.007389f
C884 B.n302 VSUBS 0.007389f
C885 B.n303 VSUBS 0.007389f
C886 B.n304 VSUBS 0.007389f
C887 B.n305 VSUBS 0.007389f
C888 B.n306 VSUBS 0.007389f
C889 B.n307 VSUBS 0.007389f
C890 B.n308 VSUBS 0.007389f
C891 B.n309 VSUBS 0.007389f
C892 B.n310 VSUBS 0.007389f
C893 B.n311 VSUBS 0.007389f
C894 B.n312 VSUBS 0.007389f
C895 B.n313 VSUBS 0.007389f
C896 B.n314 VSUBS 0.007389f
C897 B.n315 VSUBS 0.007389f
C898 B.n316 VSUBS 0.007389f
C899 B.n317 VSUBS 0.007389f
C900 B.n318 VSUBS 0.007389f
C901 B.n319 VSUBS 0.007389f
C902 B.n320 VSUBS 0.007389f
C903 B.n321 VSUBS 0.007389f
C904 B.n322 VSUBS 0.007389f
C905 B.n323 VSUBS 0.007389f
C906 B.n324 VSUBS 0.007389f
C907 B.n325 VSUBS 0.007389f
C908 B.n326 VSUBS 0.016999f
C909 B.n327 VSUBS 0.016072f
C910 B.n328 VSUBS 0.01718f
C911 B.n329 VSUBS 0.007389f
C912 B.n330 VSUBS 0.007389f
C913 B.n331 VSUBS 0.007389f
C914 B.n332 VSUBS 0.007389f
C915 B.n333 VSUBS 0.007389f
C916 B.n334 VSUBS 0.007389f
C917 B.n335 VSUBS 0.007389f
C918 B.n336 VSUBS 0.007389f
C919 B.n337 VSUBS 0.007389f
C920 B.n338 VSUBS 0.007389f
C921 B.n339 VSUBS 0.007389f
C922 B.n340 VSUBS 0.007389f
C923 B.n341 VSUBS 0.007389f
C924 B.n342 VSUBS 0.007389f
C925 B.n343 VSUBS 0.007389f
C926 B.n344 VSUBS 0.007389f
C927 B.n345 VSUBS 0.007389f
C928 B.n346 VSUBS 0.007389f
C929 B.n347 VSUBS 0.007389f
C930 B.n348 VSUBS 0.007389f
C931 B.n349 VSUBS 0.007389f
C932 B.n350 VSUBS 0.007389f
C933 B.n351 VSUBS 0.007389f
C934 B.n352 VSUBS 0.007389f
C935 B.n353 VSUBS 0.007389f
C936 B.n354 VSUBS 0.007389f
C937 B.n355 VSUBS 0.007389f
C938 B.n356 VSUBS 0.007389f
C939 B.n357 VSUBS 0.007389f
C940 B.n358 VSUBS 0.007389f
C941 B.n359 VSUBS 0.007389f
C942 B.n360 VSUBS 0.007389f
C943 B.n361 VSUBS 0.007389f
C944 B.n362 VSUBS 0.007389f
C945 B.n363 VSUBS 0.007389f
C946 B.n364 VSUBS 0.007389f
C947 B.n365 VSUBS 0.007389f
C948 B.n366 VSUBS 0.007389f
C949 B.n367 VSUBS 0.007389f
C950 B.n368 VSUBS 0.007389f
C951 B.n369 VSUBS 0.007389f
C952 B.n370 VSUBS 0.007389f
C953 B.n371 VSUBS 0.007389f
C954 B.n372 VSUBS 0.007389f
C955 B.n373 VSUBS 0.007389f
C956 B.n374 VSUBS 0.007389f
C957 B.n375 VSUBS 0.007389f
C958 B.n376 VSUBS 0.007389f
C959 B.n377 VSUBS 0.007389f
C960 B.n378 VSUBS 0.007389f
C961 B.n379 VSUBS 0.007389f
C962 B.n380 VSUBS 0.007389f
C963 B.n381 VSUBS 0.007389f
C964 B.n382 VSUBS 0.007389f
C965 B.n383 VSUBS 0.007389f
C966 B.n384 VSUBS 0.007389f
C967 B.n385 VSUBS 0.007389f
C968 B.n386 VSUBS 0.007389f
C969 B.n387 VSUBS 0.007389f
C970 B.n388 VSUBS 0.007389f
C971 B.n389 VSUBS 0.007389f
C972 B.n390 VSUBS 0.007389f
C973 B.n391 VSUBS 0.007389f
C974 B.n392 VSUBS 0.007389f
C975 B.n393 VSUBS 0.007389f
C976 B.n394 VSUBS 0.007389f
C977 B.n395 VSUBS 0.007389f
C978 B.n396 VSUBS 0.007389f
C979 B.n397 VSUBS 0.007389f
C980 B.n398 VSUBS 0.007389f
C981 B.n399 VSUBS 0.007389f
C982 B.n400 VSUBS 0.007389f
C983 B.n401 VSUBS 0.007389f
C984 B.n402 VSUBS 0.007389f
C985 B.n403 VSUBS 0.007389f
C986 B.n404 VSUBS 0.007389f
C987 B.n405 VSUBS 0.007389f
C988 B.n406 VSUBS 0.007389f
C989 B.n407 VSUBS 0.016253f
C990 B.n408 VSUBS 0.016253f
C991 B.n409 VSUBS 0.016999f
C992 B.n410 VSUBS 0.007389f
C993 B.n411 VSUBS 0.007389f
C994 B.n412 VSUBS 0.007389f
C995 B.n413 VSUBS 0.007389f
C996 B.n414 VSUBS 0.007389f
C997 B.n415 VSUBS 0.007389f
C998 B.n416 VSUBS 0.007389f
C999 B.n417 VSUBS 0.007389f
C1000 B.n418 VSUBS 0.007389f
C1001 B.n419 VSUBS 0.007389f
C1002 B.n420 VSUBS 0.007389f
C1003 B.n421 VSUBS 0.007389f
C1004 B.n422 VSUBS 0.007389f
C1005 B.n423 VSUBS 0.007389f
C1006 B.n424 VSUBS 0.007389f
C1007 B.n425 VSUBS 0.007389f
C1008 B.n426 VSUBS 0.007389f
C1009 B.n427 VSUBS 0.007389f
C1010 B.n428 VSUBS 0.007389f
C1011 B.n429 VSUBS 0.007389f
C1012 B.n430 VSUBS 0.007389f
C1013 B.n431 VSUBS 0.007389f
C1014 B.n432 VSUBS 0.007389f
C1015 B.n433 VSUBS 0.007389f
C1016 B.n434 VSUBS 0.007389f
C1017 B.n435 VSUBS 0.007389f
C1018 B.n436 VSUBS 0.007389f
C1019 B.n437 VSUBS 0.007389f
C1020 B.n438 VSUBS 0.007389f
C1021 B.n439 VSUBS 0.007389f
C1022 B.n440 VSUBS 0.007389f
C1023 B.n441 VSUBS 0.007389f
C1024 B.n442 VSUBS 0.007389f
C1025 B.n443 VSUBS 0.007389f
C1026 B.n444 VSUBS 0.007389f
C1027 B.n445 VSUBS 0.007389f
C1028 B.n446 VSUBS 0.007389f
C1029 B.n447 VSUBS 0.007389f
C1030 B.n448 VSUBS 0.007389f
C1031 B.n449 VSUBS 0.007389f
C1032 B.n450 VSUBS 0.007389f
C1033 B.n451 VSUBS 0.007389f
C1034 B.n452 VSUBS 0.007389f
C1035 B.n453 VSUBS 0.007389f
C1036 B.n454 VSUBS 0.007389f
C1037 B.n455 VSUBS 0.007389f
C1038 B.n456 VSUBS 0.007389f
C1039 B.n457 VSUBS 0.007389f
C1040 B.n458 VSUBS 0.007389f
C1041 B.n459 VSUBS 0.007389f
C1042 B.n460 VSUBS 0.007389f
C1043 B.n461 VSUBS 0.007389f
C1044 B.n462 VSUBS 0.007389f
C1045 B.n463 VSUBS 0.007389f
C1046 B.n464 VSUBS 0.007389f
C1047 B.n465 VSUBS 0.007389f
C1048 B.n466 VSUBS 0.007389f
C1049 B.n467 VSUBS 0.006955f
C1050 B.n468 VSUBS 0.007389f
C1051 B.n469 VSUBS 0.007389f
C1052 B.n470 VSUBS 0.004129f
C1053 B.n471 VSUBS 0.007389f
C1054 B.n472 VSUBS 0.007389f
C1055 B.n473 VSUBS 0.007389f
C1056 B.n474 VSUBS 0.007389f
C1057 B.n475 VSUBS 0.007389f
C1058 B.n476 VSUBS 0.007389f
C1059 B.n477 VSUBS 0.007389f
C1060 B.n478 VSUBS 0.007389f
C1061 B.n479 VSUBS 0.007389f
C1062 B.n480 VSUBS 0.007389f
C1063 B.n481 VSUBS 0.007389f
C1064 B.n482 VSUBS 0.007389f
C1065 B.n483 VSUBS 0.004129f
C1066 B.n484 VSUBS 0.01712f
C1067 B.n485 VSUBS 0.006955f
C1068 B.n486 VSUBS 0.007389f
C1069 B.n487 VSUBS 0.007389f
C1070 B.n488 VSUBS 0.007389f
C1071 B.n489 VSUBS 0.007389f
C1072 B.n490 VSUBS 0.007389f
C1073 B.n491 VSUBS 0.007389f
C1074 B.n492 VSUBS 0.007389f
C1075 B.n493 VSUBS 0.007389f
C1076 B.n494 VSUBS 0.007389f
C1077 B.n495 VSUBS 0.007389f
C1078 B.n496 VSUBS 0.007389f
C1079 B.n497 VSUBS 0.007389f
C1080 B.n498 VSUBS 0.007389f
C1081 B.n499 VSUBS 0.007389f
C1082 B.n500 VSUBS 0.007389f
C1083 B.n501 VSUBS 0.007389f
C1084 B.n502 VSUBS 0.007389f
C1085 B.n503 VSUBS 0.007389f
C1086 B.n504 VSUBS 0.007389f
C1087 B.n505 VSUBS 0.007389f
C1088 B.n506 VSUBS 0.007389f
C1089 B.n507 VSUBS 0.007389f
C1090 B.n508 VSUBS 0.007389f
C1091 B.n509 VSUBS 0.007389f
C1092 B.n510 VSUBS 0.007389f
C1093 B.n511 VSUBS 0.007389f
C1094 B.n512 VSUBS 0.007389f
C1095 B.n513 VSUBS 0.007389f
C1096 B.n514 VSUBS 0.007389f
C1097 B.n515 VSUBS 0.007389f
C1098 B.n516 VSUBS 0.007389f
C1099 B.n517 VSUBS 0.007389f
C1100 B.n518 VSUBS 0.007389f
C1101 B.n519 VSUBS 0.007389f
C1102 B.n520 VSUBS 0.007389f
C1103 B.n521 VSUBS 0.007389f
C1104 B.n522 VSUBS 0.007389f
C1105 B.n523 VSUBS 0.007389f
C1106 B.n524 VSUBS 0.007389f
C1107 B.n525 VSUBS 0.007389f
C1108 B.n526 VSUBS 0.007389f
C1109 B.n527 VSUBS 0.007389f
C1110 B.n528 VSUBS 0.007389f
C1111 B.n529 VSUBS 0.007389f
C1112 B.n530 VSUBS 0.007389f
C1113 B.n531 VSUBS 0.007389f
C1114 B.n532 VSUBS 0.007389f
C1115 B.n533 VSUBS 0.007389f
C1116 B.n534 VSUBS 0.007389f
C1117 B.n535 VSUBS 0.007389f
C1118 B.n536 VSUBS 0.007389f
C1119 B.n537 VSUBS 0.007389f
C1120 B.n538 VSUBS 0.007389f
C1121 B.n539 VSUBS 0.007389f
C1122 B.n540 VSUBS 0.007389f
C1123 B.n541 VSUBS 0.007389f
C1124 B.n542 VSUBS 0.007389f
C1125 B.n543 VSUBS 0.007389f
C1126 B.n544 VSUBS 0.016999f
C1127 B.n545 VSUBS 0.016253f
C1128 B.n546 VSUBS 0.016253f
C1129 B.n547 VSUBS 0.007389f
C1130 B.n548 VSUBS 0.007389f
C1131 B.n549 VSUBS 0.007389f
C1132 B.n550 VSUBS 0.007389f
C1133 B.n551 VSUBS 0.007389f
C1134 B.n552 VSUBS 0.007389f
C1135 B.n553 VSUBS 0.007389f
C1136 B.n554 VSUBS 0.007389f
C1137 B.n555 VSUBS 0.007389f
C1138 B.n556 VSUBS 0.007389f
C1139 B.n557 VSUBS 0.007389f
C1140 B.n558 VSUBS 0.007389f
C1141 B.n559 VSUBS 0.007389f
C1142 B.n560 VSUBS 0.007389f
C1143 B.n561 VSUBS 0.007389f
C1144 B.n562 VSUBS 0.007389f
C1145 B.n563 VSUBS 0.007389f
C1146 B.n564 VSUBS 0.007389f
C1147 B.n565 VSUBS 0.007389f
C1148 B.n566 VSUBS 0.007389f
C1149 B.n567 VSUBS 0.007389f
C1150 B.n568 VSUBS 0.007389f
C1151 B.n569 VSUBS 0.007389f
C1152 B.n570 VSUBS 0.007389f
C1153 B.n571 VSUBS 0.007389f
C1154 B.n572 VSUBS 0.007389f
C1155 B.n573 VSUBS 0.007389f
C1156 B.n574 VSUBS 0.007389f
C1157 B.n575 VSUBS 0.007389f
C1158 B.n576 VSUBS 0.007389f
C1159 B.n577 VSUBS 0.007389f
C1160 B.n578 VSUBS 0.007389f
C1161 B.n579 VSUBS 0.007389f
C1162 B.n580 VSUBS 0.007389f
C1163 B.n581 VSUBS 0.007389f
C1164 B.n582 VSUBS 0.007389f
C1165 B.n583 VSUBS 0.009643f
C1166 B.n584 VSUBS 0.010272f
C1167 B.n585 VSUBS 0.020427f
.ends

