* NGSPICE file created from diff_pair_sample_0655.ext - technology: sky130A

.subckt diff_pair_sample_0655 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=3.00465 pd=18.54 as=7.1019 ps=37.2 w=18.21 l=0.84
X1 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=7.1019 pd=37.2 as=0 ps=0 w=18.21 l=0.84
X2 VDD2.t5 VN.t0 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=7.1019 pd=37.2 as=3.00465 ps=18.54 w=18.21 l=0.84
X3 VDD1.t4 VP.t1 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=7.1019 pd=37.2 as=3.00465 ps=18.54 w=18.21 l=0.84
X4 VTAIL.t8 VP.t2 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=3.00465 pd=18.54 as=3.00465 ps=18.54 w=18.21 l=0.84
X5 VDD1.t2 VP.t3 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=7.1019 pd=37.2 as=3.00465 ps=18.54 w=18.21 l=0.84
X6 VDD1.t1 VP.t4 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=3.00465 pd=18.54 as=7.1019 ps=37.2 w=18.21 l=0.84
X7 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=7.1019 pd=37.2 as=0 ps=0 w=18.21 l=0.84
X8 VDD2.t4 VN.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=7.1019 pd=37.2 as=3.00465 ps=18.54 w=18.21 l=0.84
X9 VDD2.t3 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.00465 pd=18.54 as=7.1019 ps=37.2 w=18.21 l=0.84
X10 VTAIL.t9 VP.t5 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=3.00465 pd=18.54 as=3.00465 ps=18.54 w=18.21 l=0.84
X11 VDD2.t2 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.00465 pd=18.54 as=7.1019 ps=37.2 w=18.21 l=0.84
X12 VTAIL.t3 VN.t4 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=3.00465 pd=18.54 as=3.00465 ps=18.54 w=18.21 l=0.84
X13 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.1019 pd=37.2 as=0 ps=0 w=18.21 l=0.84
X14 VTAIL.t0 VN.t5 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.00465 pd=18.54 as=3.00465 ps=18.54 w=18.21 l=0.84
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.1019 pd=37.2 as=0 ps=0 w=18.21 l=0.84
R0 VP.n3 VP.t1 584.812
R1 VP.n1 VP.t3 569.506
R2 VP.n13 VP.t4 569.506
R3 VP.n6 VP.t0 569.506
R4 VP.n11 VP.t2 522.455
R5 VP.n4 VP.t5 522.455
R6 VP.n5 VP.n2 161.3
R7 VP.n12 VP.n0 161.3
R8 VP.n10 VP.n9 161.3
R9 VP.n7 VP.n6 80.6037
R10 VP.n14 VP.n13 80.6037
R11 VP.n8 VP.n1 80.6037
R12 VP.n10 VP.n1 56.5193
R13 VP.n13 VP.n12 56.5193
R14 VP.n6 VP.n5 56.5193
R15 VP.n8 VP.n7 46.5961
R16 VP.n3 VP.n2 43.8693
R17 VP.n4 VP.n3 42.7544
R18 VP.n11 VP.n10 12.234
R19 VP.n12 VP.n11 12.234
R20 VP.n5 VP.n4 12.234
R21 VP.n7 VP.n2 0.285035
R22 VP.n9 VP.n8 0.285035
R23 VP.n14 VP.n0 0.285035
R24 VP.n9 VP.n0 0.189894
R25 VP VP.n14 0.146778
R26 VTAIL.n410 VTAIL.n314 289.615
R27 VTAIL.n98 VTAIL.n2 289.615
R28 VTAIL.n308 VTAIL.n212 289.615
R29 VTAIL.n204 VTAIL.n108 289.615
R30 VTAIL.n346 VTAIL.n345 185
R31 VTAIL.n351 VTAIL.n350 185
R32 VTAIL.n353 VTAIL.n352 185
R33 VTAIL.n342 VTAIL.n341 185
R34 VTAIL.n359 VTAIL.n358 185
R35 VTAIL.n361 VTAIL.n360 185
R36 VTAIL.n338 VTAIL.n337 185
R37 VTAIL.n367 VTAIL.n366 185
R38 VTAIL.n369 VTAIL.n368 185
R39 VTAIL.n334 VTAIL.n333 185
R40 VTAIL.n375 VTAIL.n374 185
R41 VTAIL.n377 VTAIL.n376 185
R42 VTAIL.n330 VTAIL.n329 185
R43 VTAIL.n383 VTAIL.n382 185
R44 VTAIL.n385 VTAIL.n384 185
R45 VTAIL.n326 VTAIL.n325 185
R46 VTAIL.n392 VTAIL.n391 185
R47 VTAIL.n393 VTAIL.n324 185
R48 VTAIL.n395 VTAIL.n394 185
R49 VTAIL.n322 VTAIL.n321 185
R50 VTAIL.n401 VTAIL.n400 185
R51 VTAIL.n403 VTAIL.n402 185
R52 VTAIL.n318 VTAIL.n317 185
R53 VTAIL.n409 VTAIL.n408 185
R54 VTAIL.n411 VTAIL.n410 185
R55 VTAIL.n34 VTAIL.n33 185
R56 VTAIL.n39 VTAIL.n38 185
R57 VTAIL.n41 VTAIL.n40 185
R58 VTAIL.n30 VTAIL.n29 185
R59 VTAIL.n47 VTAIL.n46 185
R60 VTAIL.n49 VTAIL.n48 185
R61 VTAIL.n26 VTAIL.n25 185
R62 VTAIL.n55 VTAIL.n54 185
R63 VTAIL.n57 VTAIL.n56 185
R64 VTAIL.n22 VTAIL.n21 185
R65 VTAIL.n63 VTAIL.n62 185
R66 VTAIL.n65 VTAIL.n64 185
R67 VTAIL.n18 VTAIL.n17 185
R68 VTAIL.n71 VTAIL.n70 185
R69 VTAIL.n73 VTAIL.n72 185
R70 VTAIL.n14 VTAIL.n13 185
R71 VTAIL.n80 VTAIL.n79 185
R72 VTAIL.n81 VTAIL.n12 185
R73 VTAIL.n83 VTAIL.n82 185
R74 VTAIL.n10 VTAIL.n9 185
R75 VTAIL.n89 VTAIL.n88 185
R76 VTAIL.n91 VTAIL.n90 185
R77 VTAIL.n6 VTAIL.n5 185
R78 VTAIL.n97 VTAIL.n96 185
R79 VTAIL.n99 VTAIL.n98 185
R80 VTAIL.n309 VTAIL.n308 185
R81 VTAIL.n307 VTAIL.n306 185
R82 VTAIL.n216 VTAIL.n215 185
R83 VTAIL.n301 VTAIL.n300 185
R84 VTAIL.n299 VTAIL.n298 185
R85 VTAIL.n220 VTAIL.n219 185
R86 VTAIL.n293 VTAIL.n292 185
R87 VTAIL.n291 VTAIL.n222 185
R88 VTAIL.n290 VTAIL.n289 185
R89 VTAIL.n225 VTAIL.n223 185
R90 VTAIL.n284 VTAIL.n283 185
R91 VTAIL.n282 VTAIL.n281 185
R92 VTAIL.n229 VTAIL.n228 185
R93 VTAIL.n276 VTAIL.n275 185
R94 VTAIL.n274 VTAIL.n273 185
R95 VTAIL.n233 VTAIL.n232 185
R96 VTAIL.n268 VTAIL.n267 185
R97 VTAIL.n266 VTAIL.n265 185
R98 VTAIL.n237 VTAIL.n236 185
R99 VTAIL.n260 VTAIL.n259 185
R100 VTAIL.n258 VTAIL.n257 185
R101 VTAIL.n241 VTAIL.n240 185
R102 VTAIL.n252 VTAIL.n251 185
R103 VTAIL.n250 VTAIL.n249 185
R104 VTAIL.n245 VTAIL.n244 185
R105 VTAIL.n205 VTAIL.n204 185
R106 VTAIL.n203 VTAIL.n202 185
R107 VTAIL.n112 VTAIL.n111 185
R108 VTAIL.n197 VTAIL.n196 185
R109 VTAIL.n195 VTAIL.n194 185
R110 VTAIL.n116 VTAIL.n115 185
R111 VTAIL.n189 VTAIL.n188 185
R112 VTAIL.n187 VTAIL.n118 185
R113 VTAIL.n186 VTAIL.n185 185
R114 VTAIL.n121 VTAIL.n119 185
R115 VTAIL.n180 VTAIL.n179 185
R116 VTAIL.n178 VTAIL.n177 185
R117 VTAIL.n125 VTAIL.n124 185
R118 VTAIL.n172 VTAIL.n171 185
R119 VTAIL.n170 VTAIL.n169 185
R120 VTAIL.n129 VTAIL.n128 185
R121 VTAIL.n164 VTAIL.n163 185
R122 VTAIL.n162 VTAIL.n161 185
R123 VTAIL.n133 VTAIL.n132 185
R124 VTAIL.n156 VTAIL.n155 185
R125 VTAIL.n154 VTAIL.n153 185
R126 VTAIL.n137 VTAIL.n136 185
R127 VTAIL.n148 VTAIL.n147 185
R128 VTAIL.n146 VTAIL.n145 185
R129 VTAIL.n141 VTAIL.n140 185
R130 VTAIL.n347 VTAIL.t2 147.659
R131 VTAIL.n35 VTAIL.t6 147.659
R132 VTAIL.n246 VTAIL.t10 147.659
R133 VTAIL.n142 VTAIL.t1 147.659
R134 VTAIL.n351 VTAIL.n345 104.615
R135 VTAIL.n352 VTAIL.n351 104.615
R136 VTAIL.n352 VTAIL.n341 104.615
R137 VTAIL.n359 VTAIL.n341 104.615
R138 VTAIL.n360 VTAIL.n359 104.615
R139 VTAIL.n360 VTAIL.n337 104.615
R140 VTAIL.n367 VTAIL.n337 104.615
R141 VTAIL.n368 VTAIL.n367 104.615
R142 VTAIL.n368 VTAIL.n333 104.615
R143 VTAIL.n375 VTAIL.n333 104.615
R144 VTAIL.n376 VTAIL.n375 104.615
R145 VTAIL.n376 VTAIL.n329 104.615
R146 VTAIL.n383 VTAIL.n329 104.615
R147 VTAIL.n384 VTAIL.n383 104.615
R148 VTAIL.n384 VTAIL.n325 104.615
R149 VTAIL.n392 VTAIL.n325 104.615
R150 VTAIL.n393 VTAIL.n392 104.615
R151 VTAIL.n394 VTAIL.n393 104.615
R152 VTAIL.n394 VTAIL.n321 104.615
R153 VTAIL.n401 VTAIL.n321 104.615
R154 VTAIL.n402 VTAIL.n401 104.615
R155 VTAIL.n402 VTAIL.n317 104.615
R156 VTAIL.n409 VTAIL.n317 104.615
R157 VTAIL.n410 VTAIL.n409 104.615
R158 VTAIL.n39 VTAIL.n33 104.615
R159 VTAIL.n40 VTAIL.n39 104.615
R160 VTAIL.n40 VTAIL.n29 104.615
R161 VTAIL.n47 VTAIL.n29 104.615
R162 VTAIL.n48 VTAIL.n47 104.615
R163 VTAIL.n48 VTAIL.n25 104.615
R164 VTAIL.n55 VTAIL.n25 104.615
R165 VTAIL.n56 VTAIL.n55 104.615
R166 VTAIL.n56 VTAIL.n21 104.615
R167 VTAIL.n63 VTAIL.n21 104.615
R168 VTAIL.n64 VTAIL.n63 104.615
R169 VTAIL.n64 VTAIL.n17 104.615
R170 VTAIL.n71 VTAIL.n17 104.615
R171 VTAIL.n72 VTAIL.n71 104.615
R172 VTAIL.n72 VTAIL.n13 104.615
R173 VTAIL.n80 VTAIL.n13 104.615
R174 VTAIL.n81 VTAIL.n80 104.615
R175 VTAIL.n82 VTAIL.n81 104.615
R176 VTAIL.n82 VTAIL.n9 104.615
R177 VTAIL.n89 VTAIL.n9 104.615
R178 VTAIL.n90 VTAIL.n89 104.615
R179 VTAIL.n90 VTAIL.n5 104.615
R180 VTAIL.n97 VTAIL.n5 104.615
R181 VTAIL.n98 VTAIL.n97 104.615
R182 VTAIL.n308 VTAIL.n307 104.615
R183 VTAIL.n307 VTAIL.n215 104.615
R184 VTAIL.n300 VTAIL.n215 104.615
R185 VTAIL.n300 VTAIL.n299 104.615
R186 VTAIL.n299 VTAIL.n219 104.615
R187 VTAIL.n292 VTAIL.n219 104.615
R188 VTAIL.n292 VTAIL.n291 104.615
R189 VTAIL.n291 VTAIL.n290 104.615
R190 VTAIL.n290 VTAIL.n223 104.615
R191 VTAIL.n283 VTAIL.n223 104.615
R192 VTAIL.n283 VTAIL.n282 104.615
R193 VTAIL.n282 VTAIL.n228 104.615
R194 VTAIL.n275 VTAIL.n228 104.615
R195 VTAIL.n275 VTAIL.n274 104.615
R196 VTAIL.n274 VTAIL.n232 104.615
R197 VTAIL.n267 VTAIL.n232 104.615
R198 VTAIL.n267 VTAIL.n266 104.615
R199 VTAIL.n266 VTAIL.n236 104.615
R200 VTAIL.n259 VTAIL.n236 104.615
R201 VTAIL.n259 VTAIL.n258 104.615
R202 VTAIL.n258 VTAIL.n240 104.615
R203 VTAIL.n251 VTAIL.n240 104.615
R204 VTAIL.n251 VTAIL.n250 104.615
R205 VTAIL.n250 VTAIL.n244 104.615
R206 VTAIL.n204 VTAIL.n203 104.615
R207 VTAIL.n203 VTAIL.n111 104.615
R208 VTAIL.n196 VTAIL.n111 104.615
R209 VTAIL.n196 VTAIL.n195 104.615
R210 VTAIL.n195 VTAIL.n115 104.615
R211 VTAIL.n188 VTAIL.n115 104.615
R212 VTAIL.n188 VTAIL.n187 104.615
R213 VTAIL.n187 VTAIL.n186 104.615
R214 VTAIL.n186 VTAIL.n119 104.615
R215 VTAIL.n179 VTAIL.n119 104.615
R216 VTAIL.n179 VTAIL.n178 104.615
R217 VTAIL.n178 VTAIL.n124 104.615
R218 VTAIL.n171 VTAIL.n124 104.615
R219 VTAIL.n171 VTAIL.n170 104.615
R220 VTAIL.n170 VTAIL.n128 104.615
R221 VTAIL.n163 VTAIL.n128 104.615
R222 VTAIL.n163 VTAIL.n162 104.615
R223 VTAIL.n162 VTAIL.n132 104.615
R224 VTAIL.n155 VTAIL.n132 104.615
R225 VTAIL.n155 VTAIL.n154 104.615
R226 VTAIL.n154 VTAIL.n136 104.615
R227 VTAIL.n147 VTAIL.n136 104.615
R228 VTAIL.n147 VTAIL.n146 104.615
R229 VTAIL.n146 VTAIL.n140 104.615
R230 VTAIL.t2 VTAIL.n345 52.3082
R231 VTAIL.t6 VTAIL.n33 52.3082
R232 VTAIL.t10 VTAIL.n244 52.3082
R233 VTAIL.t1 VTAIL.n140 52.3082
R234 VTAIL.n211 VTAIL.n210 43.3877
R235 VTAIL.n107 VTAIL.n106 43.3877
R236 VTAIL.n1 VTAIL.n0 43.3875
R237 VTAIL.n105 VTAIL.n104 43.3875
R238 VTAIL.n415 VTAIL.n414 31.6035
R239 VTAIL.n103 VTAIL.n102 31.6035
R240 VTAIL.n313 VTAIL.n312 31.6035
R241 VTAIL.n209 VTAIL.n208 31.6035
R242 VTAIL.n107 VTAIL.n105 30.0824
R243 VTAIL.n415 VTAIL.n313 29.0738
R244 VTAIL.n347 VTAIL.n346 15.6677
R245 VTAIL.n35 VTAIL.n34 15.6677
R246 VTAIL.n246 VTAIL.n245 15.6677
R247 VTAIL.n142 VTAIL.n141 15.6677
R248 VTAIL.n395 VTAIL.n324 13.1884
R249 VTAIL.n83 VTAIL.n12 13.1884
R250 VTAIL.n293 VTAIL.n222 13.1884
R251 VTAIL.n189 VTAIL.n118 13.1884
R252 VTAIL.n350 VTAIL.n349 12.8005
R253 VTAIL.n391 VTAIL.n390 12.8005
R254 VTAIL.n396 VTAIL.n322 12.8005
R255 VTAIL.n38 VTAIL.n37 12.8005
R256 VTAIL.n79 VTAIL.n78 12.8005
R257 VTAIL.n84 VTAIL.n10 12.8005
R258 VTAIL.n294 VTAIL.n220 12.8005
R259 VTAIL.n289 VTAIL.n224 12.8005
R260 VTAIL.n249 VTAIL.n248 12.8005
R261 VTAIL.n190 VTAIL.n116 12.8005
R262 VTAIL.n185 VTAIL.n120 12.8005
R263 VTAIL.n145 VTAIL.n144 12.8005
R264 VTAIL.n353 VTAIL.n344 12.0247
R265 VTAIL.n389 VTAIL.n326 12.0247
R266 VTAIL.n400 VTAIL.n399 12.0247
R267 VTAIL.n41 VTAIL.n32 12.0247
R268 VTAIL.n77 VTAIL.n14 12.0247
R269 VTAIL.n88 VTAIL.n87 12.0247
R270 VTAIL.n298 VTAIL.n297 12.0247
R271 VTAIL.n288 VTAIL.n225 12.0247
R272 VTAIL.n252 VTAIL.n243 12.0247
R273 VTAIL.n194 VTAIL.n193 12.0247
R274 VTAIL.n184 VTAIL.n121 12.0247
R275 VTAIL.n148 VTAIL.n139 12.0247
R276 VTAIL.n354 VTAIL.n342 11.249
R277 VTAIL.n386 VTAIL.n385 11.249
R278 VTAIL.n403 VTAIL.n320 11.249
R279 VTAIL.n42 VTAIL.n30 11.249
R280 VTAIL.n74 VTAIL.n73 11.249
R281 VTAIL.n91 VTAIL.n8 11.249
R282 VTAIL.n301 VTAIL.n218 11.249
R283 VTAIL.n285 VTAIL.n284 11.249
R284 VTAIL.n253 VTAIL.n241 11.249
R285 VTAIL.n197 VTAIL.n114 11.249
R286 VTAIL.n181 VTAIL.n180 11.249
R287 VTAIL.n149 VTAIL.n137 11.249
R288 VTAIL.n358 VTAIL.n357 10.4732
R289 VTAIL.n382 VTAIL.n328 10.4732
R290 VTAIL.n404 VTAIL.n318 10.4732
R291 VTAIL.n46 VTAIL.n45 10.4732
R292 VTAIL.n70 VTAIL.n16 10.4732
R293 VTAIL.n92 VTAIL.n6 10.4732
R294 VTAIL.n302 VTAIL.n216 10.4732
R295 VTAIL.n281 VTAIL.n227 10.4732
R296 VTAIL.n257 VTAIL.n256 10.4732
R297 VTAIL.n198 VTAIL.n112 10.4732
R298 VTAIL.n177 VTAIL.n123 10.4732
R299 VTAIL.n153 VTAIL.n152 10.4732
R300 VTAIL.n361 VTAIL.n340 9.69747
R301 VTAIL.n381 VTAIL.n330 9.69747
R302 VTAIL.n408 VTAIL.n407 9.69747
R303 VTAIL.n49 VTAIL.n28 9.69747
R304 VTAIL.n69 VTAIL.n18 9.69747
R305 VTAIL.n96 VTAIL.n95 9.69747
R306 VTAIL.n306 VTAIL.n305 9.69747
R307 VTAIL.n280 VTAIL.n229 9.69747
R308 VTAIL.n260 VTAIL.n239 9.69747
R309 VTAIL.n202 VTAIL.n201 9.69747
R310 VTAIL.n176 VTAIL.n125 9.69747
R311 VTAIL.n156 VTAIL.n135 9.69747
R312 VTAIL.n414 VTAIL.n413 9.45567
R313 VTAIL.n102 VTAIL.n101 9.45567
R314 VTAIL.n312 VTAIL.n311 9.45567
R315 VTAIL.n208 VTAIL.n207 9.45567
R316 VTAIL.n413 VTAIL.n412 9.3005
R317 VTAIL.n316 VTAIL.n315 9.3005
R318 VTAIL.n407 VTAIL.n406 9.3005
R319 VTAIL.n405 VTAIL.n404 9.3005
R320 VTAIL.n320 VTAIL.n319 9.3005
R321 VTAIL.n399 VTAIL.n398 9.3005
R322 VTAIL.n397 VTAIL.n396 9.3005
R323 VTAIL.n336 VTAIL.n335 9.3005
R324 VTAIL.n365 VTAIL.n364 9.3005
R325 VTAIL.n363 VTAIL.n362 9.3005
R326 VTAIL.n340 VTAIL.n339 9.3005
R327 VTAIL.n357 VTAIL.n356 9.3005
R328 VTAIL.n355 VTAIL.n354 9.3005
R329 VTAIL.n344 VTAIL.n343 9.3005
R330 VTAIL.n349 VTAIL.n348 9.3005
R331 VTAIL.n371 VTAIL.n370 9.3005
R332 VTAIL.n373 VTAIL.n372 9.3005
R333 VTAIL.n332 VTAIL.n331 9.3005
R334 VTAIL.n379 VTAIL.n378 9.3005
R335 VTAIL.n381 VTAIL.n380 9.3005
R336 VTAIL.n328 VTAIL.n327 9.3005
R337 VTAIL.n387 VTAIL.n386 9.3005
R338 VTAIL.n389 VTAIL.n388 9.3005
R339 VTAIL.n390 VTAIL.n323 9.3005
R340 VTAIL.n101 VTAIL.n100 9.3005
R341 VTAIL.n4 VTAIL.n3 9.3005
R342 VTAIL.n95 VTAIL.n94 9.3005
R343 VTAIL.n93 VTAIL.n92 9.3005
R344 VTAIL.n8 VTAIL.n7 9.3005
R345 VTAIL.n87 VTAIL.n86 9.3005
R346 VTAIL.n85 VTAIL.n84 9.3005
R347 VTAIL.n24 VTAIL.n23 9.3005
R348 VTAIL.n53 VTAIL.n52 9.3005
R349 VTAIL.n51 VTAIL.n50 9.3005
R350 VTAIL.n28 VTAIL.n27 9.3005
R351 VTAIL.n45 VTAIL.n44 9.3005
R352 VTAIL.n43 VTAIL.n42 9.3005
R353 VTAIL.n32 VTAIL.n31 9.3005
R354 VTAIL.n37 VTAIL.n36 9.3005
R355 VTAIL.n59 VTAIL.n58 9.3005
R356 VTAIL.n61 VTAIL.n60 9.3005
R357 VTAIL.n20 VTAIL.n19 9.3005
R358 VTAIL.n67 VTAIL.n66 9.3005
R359 VTAIL.n69 VTAIL.n68 9.3005
R360 VTAIL.n16 VTAIL.n15 9.3005
R361 VTAIL.n75 VTAIL.n74 9.3005
R362 VTAIL.n77 VTAIL.n76 9.3005
R363 VTAIL.n78 VTAIL.n11 9.3005
R364 VTAIL.n272 VTAIL.n271 9.3005
R365 VTAIL.n231 VTAIL.n230 9.3005
R366 VTAIL.n278 VTAIL.n277 9.3005
R367 VTAIL.n280 VTAIL.n279 9.3005
R368 VTAIL.n227 VTAIL.n226 9.3005
R369 VTAIL.n286 VTAIL.n285 9.3005
R370 VTAIL.n288 VTAIL.n287 9.3005
R371 VTAIL.n224 VTAIL.n221 9.3005
R372 VTAIL.n311 VTAIL.n310 9.3005
R373 VTAIL.n214 VTAIL.n213 9.3005
R374 VTAIL.n305 VTAIL.n304 9.3005
R375 VTAIL.n303 VTAIL.n302 9.3005
R376 VTAIL.n218 VTAIL.n217 9.3005
R377 VTAIL.n297 VTAIL.n296 9.3005
R378 VTAIL.n295 VTAIL.n294 9.3005
R379 VTAIL.n270 VTAIL.n269 9.3005
R380 VTAIL.n235 VTAIL.n234 9.3005
R381 VTAIL.n264 VTAIL.n263 9.3005
R382 VTAIL.n262 VTAIL.n261 9.3005
R383 VTAIL.n239 VTAIL.n238 9.3005
R384 VTAIL.n256 VTAIL.n255 9.3005
R385 VTAIL.n254 VTAIL.n253 9.3005
R386 VTAIL.n243 VTAIL.n242 9.3005
R387 VTAIL.n248 VTAIL.n247 9.3005
R388 VTAIL.n168 VTAIL.n167 9.3005
R389 VTAIL.n127 VTAIL.n126 9.3005
R390 VTAIL.n174 VTAIL.n173 9.3005
R391 VTAIL.n176 VTAIL.n175 9.3005
R392 VTAIL.n123 VTAIL.n122 9.3005
R393 VTAIL.n182 VTAIL.n181 9.3005
R394 VTAIL.n184 VTAIL.n183 9.3005
R395 VTAIL.n120 VTAIL.n117 9.3005
R396 VTAIL.n207 VTAIL.n206 9.3005
R397 VTAIL.n110 VTAIL.n109 9.3005
R398 VTAIL.n201 VTAIL.n200 9.3005
R399 VTAIL.n199 VTAIL.n198 9.3005
R400 VTAIL.n114 VTAIL.n113 9.3005
R401 VTAIL.n193 VTAIL.n192 9.3005
R402 VTAIL.n191 VTAIL.n190 9.3005
R403 VTAIL.n166 VTAIL.n165 9.3005
R404 VTAIL.n131 VTAIL.n130 9.3005
R405 VTAIL.n160 VTAIL.n159 9.3005
R406 VTAIL.n158 VTAIL.n157 9.3005
R407 VTAIL.n135 VTAIL.n134 9.3005
R408 VTAIL.n152 VTAIL.n151 9.3005
R409 VTAIL.n150 VTAIL.n149 9.3005
R410 VTAIL.n139 VTAIL.n138 9.3005
R411 VTAIL.n144 VTAIL.n143 9.3005
R412 VTAIL.n362 VTAIL.n338 8.92171
R413 VTAIL.n378 VTAIL.n377 8.92171
R414 VTAIL.n411 VTAIL.n316 8.92171
R415 VTAIL.n50 VTAIL.n26 8.92171
R416 VTAIL.n66 VTAIL.n65 8.92171
R417 VTAIL.n99 VTAIL.n4 8.92171
R418 VTAIL.n309 VTAIL.n214 8.92171
R419 VTAIL.n277 VTAIL.n276 8.92171
R420 VTAIL.n261 VTAIL.n237 8.92171
R421 VTAIL.n205 VTAIL.n110 8.92171
R422 VTAIL.n173 VTAIL.n172 8.92171
R423 VTAIL.n157 VTAIL.n133 8.92171
R424 VTAIL.n366 VTAIL.n365 8.14595
R425 VTAIL.n374 VTAIL.n332 8.14595
R426 VTAIL.n412 VTAIL.n314 8.14595
R427 VTAIL.n54 VTAIL.n53 8.14595
R428 VTAIL.n62 VTAIL.n20 8.14595
R429 VTAIL.n100 VTAIL.n2 8.14595
R430 VTAIL.n310 VTAIL.n212 8.14595
R431 VTAIL.n273 VTAIL.n231 8.14595
R432 VTAIL.n265 VTAIL.n264 8.14595
R433 VTAIL.n206 VTAIL.n108 8.14595
R434 VTAIL.n169 VTAIL.n127 8.14595
R435 VTAIL.n161 VTAIL.n160 8.14595
R436 VTAIL.n369 VTAIL.n336 7.3702
R437 VTAIL.n373 VTAIL.n334 7.3702
R438 VTAIL.n57 VTAIL.n24 7.3702
R439 VTAIL.n61 VTAIL.n22 7.3702
R440 VTAIL.n272 VTAIL.n233 7.3702
R441 VTAIL.n268 VTAIL.n235 7.3702
R442 VTAIL.n168 VTAIL.n129 7.3702
R443 VTAIL.n164 VTAIL.n131 7.3702
R444 VTAIL.n370 VTAIL.n369 6.59444
R445 VTAIL.n370 VTAIL.n334 6.59444
R446 VTAIL.n58 VTAIL.n57 6.59444
R447 VTAIL.n58 VTAIL.n22 6.59444
R448 VTAIL.n269 VTAIL.n233 6.59444
R449 VTAIL.n269 VTAIL.n268 6.59444
R450 VTAIL.n165 VTAIL.n129 6.59444
R451 VTAIL.n165 VTAIL.n164 6.59444
R452 VTAIL.n366 VTAIL.n336 5.81868
R453 VTAIL.n374 VTAIL.n373 5.81868
R454 VTAIL.n414 VTAIL.n314 5.81868
R455 VTAIL.n54 VTAIL.n24 5.81868
R456 VTAIL.n62 VTAIL.n61 5.81868
R457 VTAIL.n102 VTAIL.n2 5.81868
R458 VTAIL.n312 VTAIL.n212 5.81868
R459 VTAIL.n273 VTAIL.n272 5.81868
R460 VTAIL.n265 VTAIL.n235 5.81868
R461 VTAIL.n208 VTAIL.n108 5.81868
R462 VTAIL.n169 VTAIL.n168 5.81868
R463 VTAIL.n161 VTAIL.n131 5.81868
R464 VTAIL.n365 VTAIL.n338 5.04292
R465 VTAIL.n377 VTAIL.n332 5.04292
R466 VTAIL.n412 VTAIL.n411 5.04292
R467 VTAIL.n53 VTAIL.n26 5.04292
R468 VTAIL.n65 VTAIL.n20 5.04292
R469 VTAIL.n100 VTAIL.n99 5.04292
R470 VTAIL.n310 VTAIL.n309 5.04292
R471 VTAIL.n276 VTAIL.n231 5.04292
R472 VTAIL.n264 VTAIL.n237 5.04292
R473 VTAIL.n206 VTAIL.n205 5.04292
R474 VTAIL.n172 VTAIL.n127 5.04292
R475 VTAIL.n160 VTAIL.n133 5.04292
R476 VTAIL.n348 VTAIL.n347 4.38563
R477 VTAIL.n36 VTAIL.n35 4.38563
R478 VTAIL.n247 VTAIL.n246 4.38563
R479 VTAIL.n143 VTAIL.n142 4.38563
R480 VTAIL.n362 VTAIL.n361 4.26717
R481 VTAIL.n378 VTAIL.n330 4.26717
R482 VTAIL.n408 VTAIL.n316 4.26717
R483 VTAIL.n50 VTAIL.n49 4.26717
R484 VTAIL.n66 VTAIL.n18 4.26717
R485 VTAIL.n96 VTAIL.n4 4.26717
R486 VTAIL.n306 VTAIL.n214 4.26717
R487 VTAIL.n277 VTAIL.n229 4.26717
R488 VTAIL.n261 VTAIL.n260 4.26717
R489 VTAIL.n202 VTAIL.n110 4.26717
R490 VTAIL.n173 VTAIL.n125 4.26717
R491 VTAIL.n157 VTAIL.n156 4.26717
R492 VTAIL.n358 VTAIL.n340 3.49141
R493 VTAIL.n382 VTAIL.n381 3.49141
R494 VTAIL.n407 VTAIL.n318 3.49141
R495 VTAIL.n46 VTAIL.n28 3.49141
R496 VTAIL.n70 VTAIL.n69 3.49141
R497 VTAIL.n95 VTAIL.n6 3.49141
R498 VTAIL.n305 VTAIL.n216 3.49141
R499 VTAIL.n281 VTAIL.n280 3.49141
R500 VTAIL.n257 VTAIL.n239 3.49141
R501 VTAIL.n201 VTAIL.n112 3.49141
R502 VTAIL.n177 VTAIL.n176 3.49141
R503 VTAIL.n153 VTAIL.n135 3.49141
R504 VTAIL.n357 VTAIL.n342 2.71565
R505 VTAIL.n385 VTAIL.n328 2.71565
R506 VTAIL.n404 VTAIL.n403 2.71565
R507 VTAIL.n45 VTAIL.n30 2.71565
R508 VTAIL.n73 VTAIL.n16 2.71565
R509 VTAIL.n92 VTAIL.n91 2.71565
R510 VTAIL.n302 VTAIL.n301 2.71565
R511 VTAIL.n284 VTAIL.n227 2.71565
R512 VTAIL.n256 VTAIL.n241 2.71565
R513 VTAIL.n198 VTAIL.n197 2.71565
R514 VTAIL.n180 VTAIL.n123 2.71565
R515 VTAIL.n152 VTAIL.n137 2.71565
R516 VTAIL.n354 VTAIL.n353 1.93989
R517 VTAIL.n386 VTAIL.n326 1.93989
R518 VTAIL.n400 VTAIL.n320 1.93989
R519 VTAIL.n42 VTAIL.n41 1.93989
R520 VTAIL.n74 VTAIL.n14 1.93989
R521 VTAIL.n88 VTAIL.n8 1.93989
R522 VTAIL.n298 VTAIL.n218 1.93989
R523 VTAIL.n285 VTAIL.n225 1.93989
R524 VTAIL.n253 VTAIL.n252 1.93989
R525 VTAIL.n194 VTAIL.n114 1.93989
R526 VTAIL.n181 VTAIL.n121 1.93989
R527 VTAIL.n149 VTAIL.n148 1.93989
R528 VTAIL.n350 VTAIL.n344 1.16414
R529 VTAIL.n391 VTAIL.n389 1.16414
R530 VTAIL.n399 VTAIL.n322 1.16414
R531 VTAIL.n38 VTAIL.n32 1.16414
R532 VTAIL.n79 VTAIL.n77 1.16414
R533 VTAIL.n87 VTAIL.n10 1.16414
R534 VTAIL.n297 VTAIL.n220 1.16414
R535 VTAIL.n289 VTAIL.n288 1.16414
R536 VTAIL.n249 VTAIL.n243 1.16414
R537 VTAIL.n193 VTAIL.n116 1.16414
R538 VTAIL.n185 VTAIL.n184 1.16414
R539 VTAIL.n145 VTAIL.n139 1.16414
R540 VTAIL.n0 VTAIL.t5 1.08781
R541 VTAIL.n0 VTAIL.t3 1.08781
R542 VTAIL.n104 VTAIL.t7 1.08781
R543 VTAIL.n104 VTAIL.t8 1.08781
R544 VTAIL.n210 VTAIL.t11 1.08781
R545 VTAIL.n210 VTAIL.t9 1.08781
R546 VTAIL.n106 VTAIL.t4 1.08781
R547 VTAIL.n106 VTAIL.t0 1.08781
R548 VTAIL.n209 VTAIL.n107 1.00912
R549 VTAIL.n313 VTAIL.n211 1.00912
R550 VTAIL.n105 VTAIL.n103 1.00912
R551 VTAIL.n211 VTAIL.n209 0.974638
R552 VTAIL.n103 VTAIL.n1 0.974638
R553 VTAIL VTAIL.n415 0.698776
R554 VTAIL.n349 VTAIL.n346 0.388379
R555 VTAIL.n390 VTAIL.n324 0.388379
R556 VTAIL.n396 VTAIL.n395 0.388379
R557 VTAIL.n37 VTAIL.n34 0.388379
R558 VTAIL.n78 VTAIL.n12 0.388379
R559 VTAIL.n84 VTAIL.n83 0.388379
R560 VTAIL.n294 VTAIL.n293 0.388379
R561 VTAIL.n224 VTAIL.n222 0.388379
R562 VTAIL.n248 VTAIL.n245 0.388379
R563 VTAIL.n190 VTAIL.n189 0.388379
R564 VTAIL.n120 VTAIL.n118 0.388379
R565 VTAIL.n144 VTAIL.n141 0.388379
R566 VTAIL VTAIL.n1 0.310845
R567 VTAIL.n348 VTAIL.n343 0.155672
R568 VTAIL.n355 VTAIL.n343 0.155672
R569 VTAIL.n356 VTAIL.n355 0.155672
R570 VTAIL.n356 VTAIL.n339 0.155672
R571 VTAIL.n363 VTAIL.n339 0.155672
R572 VTAIL.n364 VTAIL.n363 0.155672
R573 VTAIL.n364 VTAIL.n335 0.155672
R574 VTAIL.n371 VTAIL.n335 0.155672
R575 VTAIL.n372 VTAIL.n371 0.155672
R576 VTAIL.n372 VTAIL.n331 0.155672
R577 VTAIL.n379 VTAIL.n331 0.155672
R578 VTAIL.n380 VTAIL.n379 0.155672
R579 VTAIL.n380 VTAIL.n327 0.155672
R580 VTAIL.n387 VTAIL.n327 0.155672
R581 VTAIL.n388 VTAIL.n387 0.155672
R582 VTAIL.n388 VTAIL.n323 0.155672
R583 VTAIL.n397 VTAIL.n323 0.155672
R584 VTAIL.n398 VTAIL.n397 0.155672
R585 VTAIL.n398 VTAIL.n319 0.155672
R586 VTAIL.n405 VTAIL.n319 0.155672
R587 VTAIL.n406 VTAIL.n405 0.155672
R588 VTAIL.n406 VTAIL.n315 0.155672
R589 VTAIL.n413 VTAIL.n315 0.155672
R590 VTAIL.n36 VTAIL.n31 0.155672
R591 VTAIL.n43 VTAIL.n31 0.155672
R592 VTAIL.n44 VTAIL.n43 0.155672
R593 VTAIL.n44 VTAIL.n27 0.155672
R594 VTAIL.n51 VTAIL.n27 0.155672
R595 VTAIL.n52 VTAIL.n51 0.155672
R596 VTAIL.n52 VTAIL.n23 0.155672
R597 VTAIL.n59 VTAIL.n23 0.155672
R598 VTAIL.n60 VTAIL.n59 0.155672
R599 VTAIL.n60 VTAIL.n19 0.155672
R600 VTAIL.n67 VTAIL.n19 0.155672
R601 VTAIL.n68 VTAIL.n67 0.155672
R602 VTAIL.n68 VTAIL.n15 0.155672
R603 VTAIL.n75 VTAIL.n15 0.155672
R604 VTAIL.n76 VTAIL.n75 0.155672
R605 VTAIL.n76 VTAIL.n11 0.155672
R606 VTAIL.n85 VTAIL.n11 0.155672
R607 VTAIL.n86 VTAIL.n85 0.155672
R608 VTAIL.n86 VTAIL.n7 0.155672
R609 VTAIL.n93 VTAIL.n7 0.155672
R610 VTAIL.n94 VTAIL.n93 0.155672
R611 VTAIL.n94 VTAIL.n3 0.155672
R612 VTAIL.n101 VTAIL.n3 0.155672
R613 VTAIL.n311 VTAIL.n213 0.155672
R614 VTAIL.n304 VTAIL.n213 0.155672
R615 VTAIL.n304 VTAIL.n303 0.155672
R616 VTAIL.n303 VTAIL.n217 0.155672
R617 VTAIL.n296 VTAIL.n217 0.155672
R618 VTAIL.n296 VTAIL.n295 0.155672
R619 VTAIL.n295 VTAIL.n221 0.155672
R620 VTAIL.n287 VTAIL.n221 0.155672
R621 VTAIL.n287 VTAIL.n286 0.155672
R622 VTAIL.n286 VTAIL.n226 0.155672
R623 VTAIL.n279 VTAIL.n226 0.155672
R624 VTAIL.n279 VTAIL.n278 0.155672
R625 VTAIL.n278 VTAIL.n230 0.155672
R626 VTAIL.n271 VTAIL.n230 0.155672
R627 VTAIL.n271 VTAIL.n270 0.155672
R628 VTAIL.n270 VTAIL.n234 0.155672
R629 VTAIL.n263 VTAIL.n234 0.155672
R630 VTAIL.n263 VTAIL.n262 0.155672
R631 VTAIL.n262 VTAIL.n238 0.155672
R632 VTAIL.n255 VTAIL.n238 0.155672
R633 VTAIL.n255 VTAIL.n254 0.155672
R634 VTAIL.n254 VTAIL.n242 0.155672
R635 VTAIL.n247 VTAIL.n242 0.155672
R636 VTAIL.n207 VTAIL.n109 0.155672
R637 VTAIL.n200 VTAIL.n109 0.155672
R638 VTAIL.n200 VTAIL.n199 0.155672
R639 VTAIL.n199 VTAIL.n113 0.155672
R640 VTAIL.n192 VTAIL.n113 0.155672
R641 VTAIL.n192 VTAIL.n191 0.155672
R642 VTAIL.n191 VTAIL.n117 0.155672
R643 VTAIL.n183 VTAIL.n117 0.155672
R644 VTAIL.n183 VTAIL.n182 0.155672
R645 VTAIL.n182 VTAIL.n122 0.155672
R646 VTAIL.n175 VTAIL.n122 0.155672
R647 VTAIL.n175 VTAIL.n174 0.155672
R648 VTAIL.n174 VTAIL.n126 0.155672
R649 VTAIL.n167 VTAIL.n126 0.155672
R650 VTAIL.n167 VTAIL.n166 0.155672
R651 VTAIL.n166 VTAIL.n130 0.155672
R652 VTAIL.n159 VTAIL.n130 0.155672
R653 VTAIL.n159 VTAIL.n158 0.155672
R654 VTAIL.n158 VTAIL.n134 0.155672
R655 VTAIL.n151 VTAIL.n134 0.155672
R656 VTAIL.n151 VTAIL.n150 0.155672
R657 VTAIL.n150 VTAIL.n138 0.155672
R658 VTAIL.n143 VTAIL.n138 0.155672
R659 VDD1.n96 VDD1.n0 289.615
R660 VDD1.n197 VDD1.n101 289.615
R661 VDD1.n97 VDD1.n96 185
R662 VDD1.n95 VDD1.n94 185
R663 VDD1.n4 VDD1.n3 185
R664 VDD1.n89 VDD1.n88 185
R665 VDD1.n87 VDD1.n86 185
R666 VDD1.n8 VDD1.n7 185
R667 VDD1.n81 VDD1.n80 185
R668 VDD1.n79 VDD1.n10 185
R669 VDD1.n78 VDD1.n77 185
R670 VDD1.n13 VDD1.n11 185
R671 VDD1.n72 VDD1.n71 185
R672 VDD1.n70 VDD1.n69 185
R673 VDD1.n17 VDD1.n16 185
R674 VDD1.n64 VDD1.n63 185
R675 VDD1.n62 VDD1.n61 185
R676 VDD1.n21 VDD1.n20 185
R677 VDD1.n56 VDD1.n55 185
R678 VDD1.n54 VDD1.n53 185
R679 VDD1.n25 VDD1.n24 185
R680 VDD1.n48 VDD1.n47 185
R681 VDD1.n46 VDD1.n45 185
R682 VDD1.n29 VDD1.n28 185
R683 VDD1.n40 VDD1.n39 185
R684 VDD1.n38 VDD1.n37 185
R685 VDD1.n33 VDD1.n32 185
R686 VDD1.n133 VDD1.n132 185
R687 VDD1.n138 VDD1.n137 185
R688 VDD1.n140 VDD1.n139 185
R689 VDD1.n129 VDD1.n128 185
R690 VDD1.n146 VDD1.n145 185
R691 VDD1.n148 VDD1.n147 185
R692 VDD1.n125 VDD1.n124 185
R693 VDD1.n154 VDD1.n153 185
R694 VDD1.n156 VDD1.n155 185
R695 VDD1.n121 VDD1.n120 185
R696 VDD1.n162 VDD1.n161 185
R697 VDD1.n164 VDD1.n163 185
R698 VDD1.n117 VDD1.n116 185
R699 VDD1.n170 VDD1.n169 185
R700 VDD1.n172 VDD1.n171 185
R701 VDD1.n113 VDD1.n112 185
R702 VDD1.n179 VDD1.n178 185
R703 VDD1.n180 VDD1.n111 185
R704 VDD1.n182 VDD1.n181 185
R705 VDD1.n109 VDD1.n108 185
R706 VDD1.n188 VDD1.n187 185
R707 VDD1.n190 VDD1.n189 185
R708 VDD1.n105 VDD1.n104 185
R709 VDD1.n196 VDD1.n195 185
R710 VDD1.n198 VDD1.n197 185
R711 VDD1.n34 VDD1.t4 147.659
R712 VDD1.n134 VDD1.t2 147.659
R713 VDD1.n96 VDD1.n95 104.615
R714 VDD1.n95 VDD1.n3 104.615
R715 VDD1.n88 VDD1.n3 104.615
R716 VDD1.n88 VDD1.n87 104.615
R717 VDD1.n87 VDD1.n7 104.615
R718 VDD1.n80 VDD1.n7 104.615
R719 VDD1.n80 VDD1.n79 104.615
R720 VDD1.n79 VDD1.n78 104.615
R721 VDD1.n78 VDD1.n11 104.615
R722 VDD1.n71 VDD1.n11 104.615
R723 VDD1.n71 VDD1.n70 104.615
R724 VDD1.n70 VDD1.n16 104.615
R725 VDD1.n63 VDD1.n16 104.615
R726 VDD1.n63 VDD1.n62 104.615
R727 VDD1.n62 VDD1.n20 104.615
R728 VDD1.n55 VDD1.n20 104.615
R729 VDD1.n55 VDD1.n54 104.615
R730 VDD1.n54 VDD1.n24 104.615
R731 VDD1.n47 VDD1.n24 104.615
R732 VDD1.n47 VDD1.n46 104.615
R733 VDD1.n46 VDD1.n28 104.615
R734 VDD1.n39 VDD1.n28 104.615
R735 VDD1.n39 VDD1.n38 104.615
R736 VDD1.n38 VDD1.n32 104.615
R737 VDD1.n138 VDD1.n132 104.615
R738 VDD1.n139 VDD1.n138 104.615
R739 VDD1.n139 VDD1.n128 104.615
R740 VDD1.n146 VDD1.n128 104.615
R741 VDD1.n147 VDD1.n146 104.615
R742 VDD1.n147 VDD1.n124 104.615
R743 VDD1.n154 VDD1.n124 104.615
R744 VDD1.n155 VDD1.n154 104.615
R745 VDD1.n155 VDD1.n120 104.615
R746 VDD1.n162 VDD1.n120 104.615
R747 VDD1.n163 VDD1.n162 104.615
R748 VDD1.n163 VDD1.n116 104.615
R749 VDD1.n170 VDD1.n116 104.615
R750 VDD1.n171 VDD1.n170 104.615
R751 VDD1.n171 VDD1.n112 104.615
R752 VDD1.n179 VDD1.n112 104.615
R753 VDD1.n180 VDD1.n179 104.615
R754 VDD1.n181 VDD1.n180 104.615
R755 VDD1.n181 VDD1.n108 104.615
R756 VDD1.n188 VDD1.n108 104.615
R757 VDD1.n189 VDD1.n188 104.615
R758 VDD1.n189 VDD1.n104 104.615
R759 VDD1.n196 VDD1.n104 104.615
R760 VDD1.n197 VDD1.n196 104.615
R761 VDD1.n203 VDD1.n202 60.2631
R762 VDD1.n205 VDD1.n204 60.0663
R763 VDD1.t4 VDD1.n32 52.3082
R764 VDD1.t2 VDD1.n132 52.3082
R765 VDD1 VDD1.n100 49.097
R766 VDD1.n203 VDD1.n201 48.9834
R767 VDD1.n205 VDD1.n203 43.7789
R768 VDD1.n34 VDD1.n33 15.6677
R769 VDD1.n134 VDD1.n133 15.6677
R770 VDD1.n81 VDD1.n10 13.1884
R771 VDD1.n182 VDD1.n111 13.1884
R772 VDD1.n82 VDD1.n8 12.8005
R773 VDD1.n77 VDD1.n12 12.8005
R774 VDD1.n37 VDD1.n36 12.8005
R775 VDD1.n137 VDD1.n136 12.8005
R776 VDD1.n178 VDD1.n177 12.8005
R777 VDD1.n183 VDD1.n109 12.8005
R778 VDD1.n86 VDD1.n85 12.0247
R779 VDD1.n76 VDD1.n13 12.0247
R780 VDD1.n40 VDD1.n31 12.0247
R781 VDD1.n140 VDD1.n131 12.0247
R782 VDD1.n176 VDD1.n113 12.0247
R783 VDD1.n187 VDD1.n186 12.0247
R784 VDD1.n89 VDD1.n6 11.249
R785 VDD1.n73 VDD1.n72 11.249
R786 VDD1.n41 VDD1.n29 11.249
R787 VDD1.n141 VDD1.n129 11.249
R788 VDD1.n173 VDD1.n172 11.249
R789 VDD1.n190 VDD1.n107 11.249
R790 VDD1.n90 VDD1.n4 10.4732
R791 VDD1.n69 VDD1.n15 10.4732
R792 VDD1.n45 VDD1.n44 10.4732
R793 VDD1.n145 VDD1.n144 10.4732
R794 VDD1.n169 VDD1.n115 10.4732
R795 VDD1.n191 VDD1.n105 10.4732
R796 VDD1.n94 VDD1.n93 9.69747
R797 VDD1.n68 VDD1.n17 9.69747
R798 VDD1.n48 VDD1.n27 9.69747
R799 VDD1.n148 VDD1.n127 9.69747
R800 VDD1.n168 VDD1.n117 9.69747
R801 VDD1.n195 VDD1.n194 9.69747
R802 VDD1.n100 VDD1.n99 9.45567
R803 VDD1.n201 VDD1.n200 9.45567
R804 VDD1.n60 VDD1.n59 9.3005
R805 VDD1.n19 VDD1.n18 9.3005
R806 VDD1.n66 VDD1.n65 9.3005
R807 VDD1.n68 VDD1.n67 9.3005
R808 VDD1.n15 VDD1.n14 9.3005
R809 VDD1.n74 VDD1.n73 9.3005
R810 VDD1.n76 VDD1.n75 9.3005
R811 VDD1.n12 VDD1.n9 9.3005
R812 VDD1.n99 VDD1.n98 9.3005
R813 VDD1.n2 VDD1.n1 9.3005
R814 VDD1.n93 VDD1.n92 9.3005
R815 VDD1.n91 VDD1.n90 9.3005
R816 VDD1.n6 VDD1.n5 9.3005
R817 VDD1.n85 VDD1.n84 9.3005
R818 VDD1.n83 VDD1.n82 9.3005
R819 VDD1.n58 VDD1.n57 9.3005
R820 VDD1.n23 VDD1.n22 9.3005
R821 VDD1.n52 VDD1.n51 9.3005
R822 VDD1.n50 VDD1.n49 9.3005
R823 VDD1.n27 VDD1.n26 9.3005
R824 VDD1.n44 VDD1.n43 9.3005
R825 VDD1.n42 VDD1.n41 9.3005
R826 VDD1.n31 VDD1.n30 9.3005
R827 VDD1.n36 VDD1.n35 9.3005
R828 VDD1.n200 VDD1.n199 9.3005
R829 VDD1.n103 VDD1.n102 9.3005
R830 VDD1.n194 VDD1.n193 9.3005
R831 VDD1.n192 VDD1.n191 9.3005
R832 VDD1.n107 VDD1.n106 9.3005
R833 VDD1.n186 VDD1.n185 9.3005
R834 VDD1.n184 VDD1.n183 9.3005
R835 VDD1.n123 VDD1.n122 9.3005
R836 VDD1.n152 VDD1.n151 9.3005
R837 VDD1.n150 VDD1.n149 9.3005
R838 VDD1.n127 VDD1.n126 9.3005
R839 VDD1.n144 VDD1.n143 9.3005
R840 VDD1.n142 VDD1.n141 9.3005
R841 VDD1.n131 VDD1.n130 9.3005
R842 VDD1.n136 VDD1.n135 9.3005
R843 VDD1.n158 VDD1.n157 9.3005
R844 VDD1.n160 VDD1.n159 9.3005
R845 VDD1.n119 VDD1.n118 9.3005
R846 VDD1.n166 VDD1.n165 9.3005
R847 VDD1.n168 VDD1.n167 9.3005
R848 VDD1.n115 VDD1.n114 9.3005
R849 VDD1.n174 VDD1.n173 9.3005
R850 VDD1.n176 VDD1.n175 9.3005
R851 VDD1.n177 VDD1.n110 9.3005
R852 VDD1.n97 VDD1.n2 8.92171
R853 VDD1.n65 VDD1.n64 8.92171
R854 VDD1.n49 VDD1.n25 8.92171
R855 VDD1.n149 VDD1.n125 8.92171
R856 VDD1.n165 VDD1.n164 8.92171
R857 VDD1.n198 VDD1.n103 8.92171
R858 VDD1.n98 VDD1.n0 8.14595
R859 VDD1.n61 VDD1.n19 8.14595
R860 VDD1.n53 VDD1.n52 8.14595
R861 VDD1.n153 VDD1.n152 8.14595
R862 VDD1.n161 VDD1.n119 8.14595
R863 VDD1.n199 VDD1.n101 8.14595
R864 VDD1.n60 VDD1.n21 7.3702
R865 VDD1.n56 VDD1.n23 7.3702
R866 VDD1.n156 VDD1.n123 7.3702
R867 VDD1.n160 VDD1.n121 7.3702
R868 VDD1.n57 VDD1.n21 6.59444
R869 VDD1.n57 VDD1.n56 6.59444
R870 VDD1.n157 VDD1.n156 6.59444
R871 VDD1.n157 VDD1.n121 6.59444
R872 VDD1.n100 VDD1.n0 5.81868
R873 VDD1.n61 VDD1.n60 5.81868
R874 VDD1.n53 VDD1.n23 5.81868
R875 VDD1.n153 VDD1.n123 5.81868
R876 VDD1.n161 VDD1.n160 5.81868
R877 VDD1.n201 VDD1.n101 5.81868
R878 VDD1.n98 VDD1.n97 5.04292
R879 VDD1.n64 VDD1.n19 5.04292
R880 VDD1.n52 VDD1.n25 5.04292
R881 VDD1.n152 VDD1.n125 5.04292
R882 VDD1.n164 VDD1.n119 5.04292
R883 VDD1.n199 VDD1.n198 5.04292
R884 VDD1.n35 VDD1.n34 4.38563
R885 VDD1.n135 VDD1.n134 4.38563
R886 VDD1.n94 VDD1.n2 4.26717
R887 VDD1.n65 VDD1.n17 4.26717
R888 VDD1.n49 VDD1.n48 4.26717
R889 VDD1.n149 VDD1.n148 4.26717
R890 VDD1.n165 VDD1.n117 4.26717
R891 VDD1.n195 VDD1.n103 4.26717
R892 VDD1.n93 VDD1.n4 3.49141
R893 VDD1.n69 VDD1.n68 3.49141
R894 VDD1.n45 VDD1.n27 3.49141
R895 VDD1.n145 VDD1.n127 3.49141
R896 VDD1.n169 VDD1.n168 3.49141
R897 VDD1.n194 VDD1.n105 3.49141
R898 VDD1.n90 VDD1.n89 2.71565
R899 VDD1.n72 VDD1.n15 2.71565
R900 VDD1.n44 VDD1.n29 2.71565
R901 VDD1.n144 VDD1.n129 2.71565
R902 VDD1.n172 VDD1.n115 2.71565
R903 VDD1.n191 VDD1.n190 2.71565
R904 VDD1.n86 VDD1.n6 1.93989
R905 VDD1.n73 VDD1.n13 1.93989
R906 VDD1.n41 VDD1.n40 1.93989
R907 VDD1.n141 VDD1.n140 1.93989
R908 VDD1.n173 VDD1.n113 1.93989
R909 VDD1.n187 VDD1.n107 1.93989
R910 VDD1.n85 VDD1.n8 1.16414
R911 VDD1.n77 VDD1.n76 1.16414
R912 VDD1.n37 VDD1.n31 1.16414
R913 VDD1.n137 VDD1.n131 1.16414
R914 VDD1.n178 VDD1.n176 1.16414
R915 VDD1.n186 VDD1.n109 1.16414
R916 VDD1.n204 VDD1.t0 1.08781
R917 VDD1.n204 VDD1.t5 1.08781
R918 VDD1.n202 VDD1.t3 1.08781
R919 VDD1.n202 VDD1.t1 1.08781
R920 VDD1.n82 VDD1.n81 0.388379
R921 VDD1.n12 VDD1.n10 0.388379
R922 VDD1.n36 VDD1.n33 0.388379
R923 VDD1.n136 VDD1.n133 0.388379
R924 VDD1.n177 VDD1.n111 0.388379
R925 VDD1.n183 VDD1.n182 0.388379
R926 VDD1 VDD1.n205 0.194466
R927 VDD1.n99 VDD1.n1 0.155672
R928 VDD1.n92 VDD1.n1 0.155672
R929 VDD1.n92 VDD1.n91 0.155672
R930 VDD1.n91 VDD1.n5 0.155672
R931 VDD1.n84 VDD1.n5 0.155672
R932 VDD1.n84 VDD1.n83 0.155672
R933 VDD1.n83 VDD1.n9 0.155672
R934 VDD1.n75 VDD1.n9 0.155672
R935 VDD1.n75 VDD1.n74 0.155672
R936 VDD1.n74 VDD1.n14 0.155672
R937 VDD1.n67 VDD1.n14 0.155672
R938 VDD1.n67 VDD1.n66 0.155672
R939 VDD1.n66 VDD1.n18 0.155672
R940 VDD1.n59 VDD1.n18 0.155672
R941 VDD1.n59 VDD1.n58 0.155672
R942 VDD1.n58 VDD1.n22 0.155672
R943 VDD1.n51 VDD1.n22 0.155672
R944 VDD1.n51 VDD1.n50 0.155672
R945 VDD1.n50 VDD1.n26 0.155672
R946 VDD1.n43 VDD1.n26 0.155672
R947 VDD1.n43 VDD1.n42 0.155672
R948 VDD1.n42 VDD1.n30 0.155672
R949 VDD1.n35 VDD1.n30 0.155672
R950 VDD1.n135 VDD1.n130 0.155672
R951 VDD1.n142 VDD1.n130 0.155672
R952 VDD1.n143 VDD1.n142 0.155672
R953 VDD1.n143 VDD1.n126 0.155672
R954 VDD1.n150 VDD1.n126 0.155672
R955 VDD1.n151 VDD1.n150 0.155672
R956 VDD1.n151 VDD1.n122 0.155672
R957 VDD1.n158 VDD1.n122 0.155672
R958 VDD1.n159 VDD1.n158 0.155672
R959 VDD1.n159 VDD1.n118 0.155672
R960 VDD1.n166 VDD1.n118 0.155672
R961 VDD1.n167 VDD1.n166 0.155672
R962 VDD1.n167 VDD1.n114 0.155672
R963 VDD1.n174 VDD1.n114 0.155672
R964 VDD1.n175 VDD1.n174 0.155672
R965 VDD1.n175 VDD1.n110 0.155672
R966 VDD1.n184 VDD1.n110 0.155672
R967 VDD1.n185 VDD1.n184 0.155672
R968 VDD1.n185 VDD1.n106 0.155672
R969 VDD1.n192 VDD1.n106 0.155672
R970 VDD1.n193 VDD1.n192 0.155672
R971 VDD1.n193 VDD1.n102 0.155672
R972 VDD1.n200 VDD1.n102 0.155672
R973 B.n191 B.t6 724.155
R974 B.n185 B.t14 724.155
R975 B.n75 B.t17 724.155
R976 B.n81 B.t10 724.155
R977 B.n577 B.n112 585
R978 B.n112 B.n43 585
R979 B.n579 B.n578 585
R980 B.n581 B.n111 585
R981 B.n584 B.n583 585
R982 B.n585 B.n110 585
R983 B.n587 B.n586 585
R984 B.n589 B.n109 585
R985 B.n592 B.n591 585
R986 B.n593 B.n108 585
R987 B.n595 B.n594 585
R988 B.n597 B.n107 585
R989 B.n600 B.n599 585
R990 B.n601 B.n106 585
R991 B.n603 B.n602 585
R992 B.n605 B.n105 585
R993 B.n608 B.n607 585
R994 B.n609 B.n104 585
R995 B.n611 B.n610 585
R996 B.n613 B.n103 585
R997 B.n616 B.n615 585
R998 B.n617 B.n102 585
R999 B.n619 B.n618 585
R1000 B.n621 B.n101 585
R1001 B.n624 B.n623 585
R1002 B.n625 B.n100 585
R1003 B.n627 B.n626 585
R1004 B.n629 B.n99 585
R1005 B.n632 B.n631 585
R1006 B.n633 B.n98 585
R1007 B.n635 B.n634 585
R1008 B.n637 B.n97 585
R1009 B.n640 B.n639 585
R1010 B.n641 B.n96 585
R1011 B.n643 B.n642 585
R1012 B.n645 B.n95 585
R1013 B.n648 B.n647 585
R1014 B.n649 B.n94 585
R1015 B.n651 B.n650 585
R1016 B.n653 B.n93 585
R1017 B.n656 B.n655 585
R1018 B.n657 B.n92 585
R1019 B.n659 B.n658 585
R1020 B.n661 B.n91 585
R1021 B.n664 B.n663 585
R1022 B.n665 B.n90 585
R1023 B.n667 B.n666 585
R1024 B.n669 B.n89 585
R1025 B.n672 B.n671 585
R1026 B.n673 B.n88 585
R1027 B.n675 B.n674 585
R1028 B.n677 B.n87 585
R1029 B.n680 B.n679 585
R1030 B.n681 B.n86 585
R1031 B.n683 B.n682 585
R1032 B.n685 B.n85 585
R1033 B.n688 B.n687 585
R1034 B.n689 B.n84 585
R1035 B.n691 B.n690 585
R1036 B.n693 B.n83 585
R1037 B.n696 B.n695 585
R1038 B.n698 B.n80 585
R1039 B.n700 B.n699 585
R1040 B.n702 B.n79 585
R1041 B.n705 B.n704 585
R1042 B.n706 B.n78 585
R1043 B.n708 B.n707 585
R1044 B.n710 B.n77 585
R1045 B.n713 B.n712 585
R1046 B.n714 B.n74 585
R1047 B.n717 B.n716 585
R1048 B.n719 B.n73 585
R1049 B.n722 B.n721 585
R1050 B.n723 B.n72 585
R1051 B.n725 B.n724 585
R1052 B.n727 B.n71 585
R1053 B.n730 B.n729 585
R1054 B.n731 B.n70 585
R1055 B.n733 B.n732 585
R1056 B.n735 B.n69 585
R1057 B.n738 B.n737 585
R1058 B.n739 B.n68 585
R1059 B.n741 B.n740 585
R1060 B.n743 B.n67 585
R1061 B.n746 B.n745 585
R1062 B.n747 B.n66 585
R1063 B.n749 B.n748 585
R1064 B.n751 B.n65 585
R1065 B.n754 B.n753 585
R1066 B.n755 B.n64 585
R1067 B.n757 B.n756 585
R1068 B.n759 B.n63 585
R1069 B.n762 B.n761 585
R1070 B.n763 B.n62 585
R1071 B.n765 B.n764 585
R1072 B.n767 B.n61 585
R1073 B.n770 B.n769 585
R1074 B.n771 B.n60 585
R1075 B.n773 B.n772 585
R1076 B.n775 B.n59 585
R1077 B.n778 B.n777 585
R1078 B.n779 B.n58 585
R1079 B.n781 B.n780 585
R1080 B.n783 B.n57 585
R1081 B.n786 B.n785 585
R1082 B.n787 B.n56 585
R1083 B.n789 B.n788 585
R1084 B.n791 B.n55 585
R1085 B.n794 B.n793 585
R1086 B.n795 B.n54 585
R1087 B.n797 B.n796 585
R1088 B.n799 B.n53 585
R1089 B.n802 B.n801 585
R1090 B.n803 B.n52 585
R1091 B.n805 B.n804 585
R1092 B.n807 B.n51 585
R1093 B.n810 B.n809 585
R1094 B.n811 B.n50 585
R1095 B.n813 B.n812 585
R1096 B.n815 B.n49 585
R1097 B.n818 B.n817 585
R1098 B.n819 B.n48 585
R1099 B.n821 B.n820 585
R1100 B.n823 B.n47 585
R1101 B.n826 B.n825 585
R1102 B.n827 B.n46 585
R1103 B.n829 B.n828 585
R1104 B.n831 B.n45 585
R1105 B.n834 B.n833 585
R1106 B.n835 B.n44 585
R1107 B.n576 B.n42 585
R1108 B.n838 B.n42 585
R1109 B.n575 B.n41 585
R1110 B.n839 B.n41 585
R1111 B.n574 B.n40 585
R1112 B.n840 B.n40 585
R1113 B.n573 B.n572 585
R1114 B.n572 B.n36 585
R1115 B.n571 B.n35 585
R1116 B.n846 B.n35 585
R1117 B.n570 B.n34 585
R1118 B.n847 B.n34 585
R1119 B.n569 B.n33 585
R1120 B.n848 B.n33 585
R1121 B.n568 B.n567 585
R1122 B.n567 B.n29 585
R1123 B.n566 B.n28 585
R1124 B.n854 B.n28 585
R1125 B.n565 B.n27 585
R1126 B.n855 B.n27 585
R1127 B.n564 B.n26 585
R1128 B.n856 B.n26 585
R1129 B.n563 B.n562 585
R1130 B.n562 B.n25 585
R1131 B.n561 B.n21 585
R1132 B.n862 B.n21 585
R1133 B.n560 B.n20 585
R1134 B.n863 B.n20 585
R1135 B.n559 B.n19 585
R1136 B.n864 B.n19 585
R1137 B.n558 B.n557 585
R1138 B.n557 B.n18 585
R1139 B.n556 B.n14 585
R1140 B.n870 B.n14 585
R1141 B.n555 B.n13 585
R1142 B.n871 B.n13 585
R1143 B.n554 B.n12 585
R1144 B.n872 B.n12 585
R1145 B.n553 B.n552 585
R1146 B.n552 B.n8 585
R1147 B.n551 B.n7 585
R1148 B.n878 B.n7 585
R1149 B.n550 B.n6 585
R1150 B.n879 B.n6 585
R1151 B.n549 B.n5 585
R1152 B.n880 B.n5 585
R1153 B.n548 B.n547 585
R1154 B.n547 B.n4 585
R1155 B.n546 B.n113 585
R1156 B.n546 B.n545 585
R1157 B.n536 B.n114 585
R1158 B.n115 B.n114 585
R1159 B.n538 B.n537 585
R1160 B.n539 B.n538 585
R1161 B.n535 B.n120 585
R1162 B.n120 B.n119 585
R1163 B.n534 B.n533 585
R1164 B.n533 B.n532 585
R1165 B.n122 B.n121 585
R1166 B.n525 B.n122 585
R1167 B.n524 B.n523 585
R1168 B.n526 B.n524 585
R1169 B.n522 B.n127 585
R1170 B.n127 B.n126 585
R1171 B.n521 B.n520 585
R1172 B.n520 B.n519 585
R1173 B.n129 B.n128 585
R1174 B.n512 B.n129 585
R1175 B.n511 B.n510 585
R1176 B.n513 B.n511 585
R1177 B.n509 B.n134 585
R1178 B.n134 B.n133 585
R1179 B.n508 B.n507 585
R1180 B.n507 B.n506 585
R1181 B.n136 B.n135 585
R1182 B.n137 B.n136 585
R1183 B.n499 B.n498 585
R1184 B.n500 B.n499 585
R1185 B.n497 B.n141 585
R1186 B.n145 B.n141 585
R1187 B.n496 B.n495 585
R1188 B.n495 B.n494 585
R1189 B.n143 B.n142 585
R1190 B.n144 B.n143 585
R1191 B.n487 B.n486 585
R1192 B.n488 B.n487 585
R1193 B.n485 B.n150 585
R1194 B.n150 B.n149 585
R1195 B.n484 B.n483 585
R1196 B.n483 B.n482 585
R1197 B.n479 B.n154 585
R1198 B.n478 B.n477 585
R1199 B.n475 B.n155 585
R1200 B.n475 B.n153 585
R1201 B.n474 B.n473 585
R1202 B.n472 B.n471 585
R1203 B.n470 B.n157 585
R1204 B.n468 B.n467 585
R1205 B.n466 B.n158 585
R1206 B.n465 B.n464 585
R1207 B.n462 B.n159 585
R1208 B.n460 B.n459 585
R1209 B.n458 B.n160 585
R1210 B.n457 B.n456 585
R1211 B.n454 B.n161 585
R1212 B.n452 B.n451 585
R1213 B.n450 B.n162 585
R1214 B.n449 B.n448 585
R1215 B.n446 B.n163 585
R1216 B.n444 B.n443 585
R1217 B.n442 B.n164 585
R1218 B.n441 B.n440 585
R1219 B.n438 B.n165 585
R1220 B.n436 B.n435 585
R1221 B.n434 B.n166 585
R1222 B.n433 B.n432 585
R1223 B.n430 B.n167 585
R1224 B.n428 B.n427 585
R1225 B.n426 B.n168 585
R1226 B.n425 B.n424 585
R1227 B.n422 B.n169 585
R1228 B.n420 B.n419 585
R1229 B.n418 B.n170 585
R1230 B.n417 B.n416 585
R1231 B.n414 B.n171 585
R1232 B.n412 B.n411 585
R1233 B.n410 B.n172 585
R1234 B.n409 B.n408 585
R1235 B.n406 B.n173 585
R1236 B.n404 B.n403 585
R1237 B.n402 B.n174 585
R1238 B.n401 B.n400 585
R1239 B.n398 B.n175 585
R1240 B.n396 B.n395 585
R1241 B.n394 B.n176 585
R1242 B.n393 B.n392 585
R1243 B.n390 B.n177 585
R1244 B.n388 B.n387 585
R1245 B.n386 B.n178 585
R1246 B.n385 B.n384 585
R1247 B.n382 B.n179 585
R1248 B.n380 B.n379 585
R1249 B.n378 B.n180 585
R1250 B.n377 B.n376 585
R1251 B.n374 B.n181 585
R1252 B.n372 B.n371 585
R1253 B.n370 B.n182 585
R1254 B.n369 B.n368 585
R1255 B.n366 B.n183 585
R1256 B.n364 B.n363 585
R1257 B.n362 B.n184 585
R1258 B.n360 B.n359 585
R1259 B.n357 B.n187 585
R1260 B.n355 B.n354 585
R1261 B.n353 B.n188 585
R1262 B.n352 B.n351 585
R1263 B.n349 B.n189 585
R1264 B.n347 B.n346 585
R1265 B.n345 B.n190 585
R1266 B.n344 B.n343 585
R1267 B.n341 B.n340 585
R1268 B.n339 B.n338 585
R1269 B.n337 B.n195 585
R1270 B.n335 B.n334 585
R1271 B.n333 B.n196 585
R1272 B.n332 B.n331 585
R1273 B.n329 B.n197 585
R1274 B.n327 B.n326 585
R1275 B.n325 B.n198 585
R1276 B.n324 B.n323 585
R1277 B.n321 B.n199 585
R1278 B.n319 B.n318 585
R1279 B.n317 B.n200 585
R1280 B.n316 B.n315 585
R1281 B.n313 B.n201 585
R1282 B.n311 B.n310 585
R1283 B.n309 B.n202 585
R1284 B.n308 B.n307 585
R1285 B.n305 B.n203 585
R1286 B.n303 B.n302 585
R1287 B.n301 B.n204 585
R1288 B.n300 B.n299 585
R1289 B.n297 B.n205 585
R1290 B.n295 B.n294 585
R1291 B.n293 B.n206 585
R1292 B.n292 B.n291 585
R1293 B.n289 B.n207 585
R1294 B.n287 B.n286 585
R1295 B.n285 B.n208 585
R1296 B.n284 B.n283 585
R1297 B.n281 B.n209 585
R1298 B.n279 B.n278 585
R1299 B.n277 B.n210 585
R1300 B.n276 B.n275 585
R1301 B.n273 B.n211 585
R1302 B.n271 B.n270 585
R1303 B.n269 B.n212 585
R1304 B.n268 B.n267 585
R1305 B.n265 B.n213 585
R1306 B.n263 B.n262 585
R1307 B.n261 B.n214 585
R1308 B.n260 B.n259 585
R1309 B.n257 B.n215 585
R1310 B.n255 B.n254 585
R1311 B.n253 B.n216 585
R1312 B.n252 B.n251 585
R1313 B.n249 B.n217 585
R1314 B.n247 B.n246 585
R1315 B.n245 B.n218 585
R1316 B.n244 B.n243 585
R1317 B.n241 B.n219 585
R1318 B.n239 B.n238 585
R1319 B.n237 B.n220 585
R1320 B.n236 B.n235 585
R1321 B.n233 B.n221 585
R1322 B.n231 B.n230 585
R1323 B.n229 B.n222 585
R1324 B.n228 B.n227 585
R1325 B.n225 B.n223 585
R1326 B.n152 B.n151 585
R1327 B.n481 B.n480 585
R1328 B.n482 B.n481 585
R1329 B.n148 B.n147 585
R1330 B.n149 B.n148 585
R1331 B.n490 B.n489 585
R1332 B.n489 B.n488 585
R1333 B.n491 B.n146 585
R1334 B.n146 B.n144 585
R1335 B.n493 B.n492 585
R1336 B.n494 B.n493 585
R1337 B.n140 B.n139 585
R1338 B.n145 B.n140 585
R1339 B.n502 B.n501 585
R1340 B.n501 B.n500 585
R1341 B.n503 B.n138 585
R1342 B.n138 B.n137 585
R1343 B.n505 B.n504 585
R1344 B.n506 B.n505 585
R1345 B.n132 B.n131 585
R1346 B.n133 B.n132 585
R1347 B.n515 B.n514 585
R1348 B.n514 B.n513 585
R1349 B.n516 B.n130 585
R1350 B.n512 B.n130 585
R1351 B.n518 B.n517 585
R1352 B.n519 B.n518 585
R1353 B.n125 B.n124 585
R1354 B.n126 B.n125 585
R1355 B.n528 B.n527 585
R1356 B.n527 B.n526 585
R1357 B.n529 B.n123 585
R1358 B.n525 B.n123 585
R1359 B.n531 B.n530 585
R1360 B.n532 B.n531 585
R1361 B.n118 B.n117 585
R1362 B.n119 B.n118 585
R1363 B.n541 B.n540 585
R1364 B.n540 B.n539 585
R1365 B.n542 B.n116 585
R1366 B.n116 B.n115 585
R1367 B.n544 B.n543 585
R1368 B.n545 B.n544 585
R1369 B.n2 B.n0 585
R1370 B.n4 B.n2 585
R1371 B.n3 B.n1 585
R1372 B.n879 B.n3 585
R1373 B.n877 B.n876 585
R1374 B.n878 B.n877 585
R1375 B.n875 B.n9 585
R1376 B.n9 B.n8 585
R1377 B.n874 B.n873 585
R1378 B.n873 B.n872 585
R1379 B.n11 B.n10 585
R1380 B.n871 B.n11 585
R1381 B.n869 B.n868 585
R1382 B.n870 B.n869 585
R1383 B.n867 B.n15 585
R1384 B.n18 B.n15 585
R1385 B.n866 B.n865 585
R1386 B.n865 B.n864 585
R1387 B.n17 B.n16 585
R1388 B.n863 B.n17 585
R1389 B.n861 B.n860 585
R1390 B.n862 B.n861 585
R1391 B.n859 B.n22 585
R1392 B.n25 B.n22 585
R1393 B.n858 B.n857 585
R1394 B.n857 B.n856 585
R1395 B.n24 B.n23 585
R1396 B.n855 B.n24 585
R1397 B.n853 B.n852 585
R1398 B.n854 B.n853 585
R1399 B.n851 B.n30 585
R1400 B.n30 B.n29 585
R1401 B.n850 B.n849 585
R1402 B.n849 B.n848 585
R1403 B.n32 B.n31 585
R1404 B.n847 B.n32 585
R1405 B.n845 B.n844 585
R1406 B.n846 B.n845 585
R1407 B.n843 B.n37 585
R1408 B.n37 B.n36 585
R1409 B.n842 B.n841 585
R1410 B.n841 B.n840 585
R1411 B.n39 B.n38 585
R1412 B.n839 B.n39 585
R1413 B.n837 B.n836 585
R1414 B.n838 B.n837 585
R1415 B.n882 B.n881 585
R1416 B.n881 B.n880 585
R1417 B.n481 B.n154 506.916
R1418 B.n837 B.n44 506.916
R1419 B.n483 B.n152 506.916
R1420 B.n112 B.n42 506.916
R1421 B.n191 B.t9 411.856
R1422 B.n81 B.t12 411.856
R1423 B.n185 B.t16 411.856
R1424 B.n75 B.t18 411.856
R1425 B.n192 B.t8 389.166
R1426 B.n82 B.t13 389.166
R1427 B.n186 B.t15 389.166
R1428 B.n76 B.t19 389.166
R1429 B.n580 B.n43 256.663
R1430 B.n582 B.n43 256.663
R1431 B.n588 B.n43 256.663
R1432 B.n590 B.n43 256.663
R1433 B.n596 B.n43 256.663
R1434 B.n598 B.n43 256.663
R1435 B.n604 B.n43 256.663
R1436 B.n606 B.n43 256.663
R1437 B.n612 B.n43 256.663
R1438 B.n614 B.n43 256.663
R1439 B.n620 B.n43 256.663
R1440 B.n622 B.n43 256.663
R1441 B.n628 B.n43 256.663
R1442 B.n630 B.n43 256.663
R1443 B.n636 B.n43 256.663
R1444 B.n638 B.n43 256.663
R1445 B.n644 B.n43 256.663
R1446 B.n646 B.n43 256.663
R1447 B.n652 B.n43 256.663
R1448 B.n654 B.n43 256.663
R1449 B.n660 B.n43 256.663
R1450 B.n662 B.n43 256.663
R1451 B.n668 B.n43 256.663
R1452 B.n670 B.n43 256.663
R1453 B.n676 B.n43 256.663
R1454 B.n678 B.n43 256.663
R1455 B.n684 B.n43 256.663
R1456 B.n686 B.n43 256.663
R1457 B.n692 B.n43 256.663
R1458 B.n694 B.n43 256.663
R1459 B.n701 B.n43 256.663
R1460 B.n703 B.n43 256.663
R1461 B.n709 B.n43 256.663
R1462 B.n711 B.n43 256.663
R1463 B.n718 B.n43 256.663
R1464 B.n720 B.n43 256.663
R1465 B.n726 B.n43 256.663
R1466 B.n728 B.n43 256.663
R1467 B.n734 B.n43 256.663
R1468 B.n736 B.n43 256.663
R1469 B.n742 B.n43 256.663
R1470 B.n744 B.n43 256.663
R1471 B.n750 B.n43 256.663
R1472 B.n752 B.n43 256.663
R1473 B.n758 B.n43 256.663
R1474 B.n760 B.n43 256.663
R1475 B.n766 B.n43 256.663
R1476 B.n768 B.n43 256.663
R1477 B.n774 B.n43 256.663
R1478 B.n776 B.n43 256.663
R1479 B.n782 B.n43 256.663
R1480 B.n784 B.n43 256.663
R1481 B.n790 B.n43 256.663
R1482 B.n792 B.n43 256.663
R1483 B.n798 B.n43 256.663
R1484 B.n800 B.n43 256.663
R1485 B.n806 B.n43 256.663
R1486 B.n808 B.n43 256.663
R1487 B.n814 B.n43 256.663
R1488 B.n816 B.n43 256.663
R1489 B.n822 B.n43 256.663
R1490 B.n824 B.n43 256.663
R1491 B.n830 B.n43 256.663
R1492 B.n832 B.n43 256.663
R1493 B.n476 B.n153 256.663
R1494 B.n156 B.n153 256.663
R1495 B.n469 B.n153 256.663
R1496 B.n463 B.n153 256.663
R1497 B.n461 B.n153 256.663
R1498 B.n455 B.n153 256.663
R1499 B.n453 B.n153 256.663
R1500 B.n447 B.n153 256.663
R1501 B.n445 B.n153 256.663
R1502 B.n439 B.n153 256.663
R1503 B.n437 B.n153 256.663
R1504 B.n431 B.n153 256.663
R1505 B.n429 B.n153 256.663
R1506 B.n423 B.n153 256.663
R1507 B.n421 B.n153 256.663
R1508 B.n415 B.n153 256.663
R1509 B.n413 B.n153 256.663
R1510 B.n407 B.n153 256.663
R1511 B.n405 B.n153 256.663
R1512 B.n399 B.n153 256.663
R1513 B.n397 B.n153 256.663
R1514 B.n391 B.n153 256.663
R1515 B.n389 B.n153 256.663
R1516 B.n383 B.n153 256.663
R1517 B.n381 B.n153 256.663
R1518 B.n375 B.n153 256.663
R1519 B.n373 B.n153 256.663
R1520 B.n367 B.n153 256.663
R1521 B.n365 B.n153 256.663
R1522 B.n358 B.n153 256.663
R1523 B.n356 B.n153 256.663
R1524 B.n350 B.n153 256.663
R1525 B.n348 B.n153 256.663
R1526 B.n342 B.n153 256.663
R1527 B.n194 B.n153 256.663
R1528 B.n336 B.n153 256.663
R1529 B.n330 B.n153 256.663
R1530 B.n328 B.n153 256.663
R1531 B.n322 B.n153 256.663
R1532 B.n320 B.n153 256.663
R1533 B.n314 B.n153 256.663
R1534 B.n312 B.n153 256.663
R1535 B.n306 B.n153 256.663
R1536 B.n304 B.n153 256.663
R1537 B.n298 B.n153 256.663
R1538 B.n296 B.n153 256.663
R1539 B.n290 B.n153 256.663
R1540 B.n288 B.n153 256.663
R1541 B.n282 B.n153 256.663
R1542 B.n280 B.n153 256.663
R1543 B.n274 B.n153 256.663
R1544 B.n272 B.n153 256.663
R1545 B.n266 B.n153 256.663
R1546 B.n264 B.n153 256.663
R1547 B.n258 B.n153 256.663
R1548 B.n256 B.n153 256.663
R1549 B.n250 B.n153 256.663
R1550 B.n248 B.n153 256.663
R1551 B.n242 B.n153 256.663
R1552 B.n240 B.n153 256.663
R1553 B.n234 B.n153 256.663
R1554 B.n232 B.n153 256.663
R1555 B.n226 B.n153 256.663
R1556 B.n224 B.n153 256.663
R1557 B.n481 B.n148 163.367
R1558 B.n489 B.n148 163.367
R1559 B.n489 B.n146 163.367
R1560 B.n493 B.n146 163.367
R1561 B.n493 B.n140 163.367
R1562 B.n501 B.n140 163.367
R1563 B.n501 B.n138 163.367
R1564 B.n505 B.n138 163.367
R1565 B.n505 B.n132 163.367
R1566 B.n514 B.n132 163.367
R1567 B.n514 B.n130 163.367
R1568 B.n518 B.n130 163.367
R1569 B.n518 B.n125 163.367
R1570 B.n527 B.n125 163.367
R1571 B.n527 B.n123 163.367
R1572 B.n531 B.n123 163.367
R1573 B.n531 B.n118 163.367
R1574 B.n540 B.n118 163.367
R1575 B.n540 B.n116 163.367
R1576 B.n544 B.n116 163.367
R1577 B.n544 B.n2 163.367
R1578 B.n881 B.n2 163.367
R1579 B.n881 B.n3 163.367
R1580 B.n877 B.n3 163.367
R1581 B.n877 B.n9 163.367
R1582 B.n873 B.n9 163.367
R1583 B.n873 B.n11 163.367
R1584 B.n869 B.n11 163.367
R1585 B.n869 B.n15 163.367
R1586 B.n865 B.n15 163.367
R1587 B.n865 B.n17 163.367
R1588 B.n861 B.n17 163.367
R1589 B.n861 B.n22 163.367
R1590 B.n857 B.n22 163.367
R1591 B.n857 B.n24 163.367
R1592 B.n853 B.n24 163.367
R1593 B.n853 B.n30 163.367
R1594 B.n849 B.n30 163.367
R1595 B.n849 B.n32 163.367
R1596 B.n845 B.n32 163.367
R1597 B.n845 B.n37 163.367
R1598 B.n841 B.n37 163.367
R1599 B.n841 B.n39 163.367
R1600 B.n837 B.n39 163.367
R1601 B.n477 B.n475 163.367
R1602 B.n475 B.n474 163.367
R1603 B.n471 B.n470 163.367
R1604 B.n468 B.n158 163.367
R1605 B.n464 B.n462 163.367
R1606 B.n460 B.n160 163.367
R1607 B.n456 B.n454 163.367
R1608 B.n452 B.n162 163.367
R1609 B.n448 B.n446 163.367
R1610 B.n444 B.n164 163.367
R1611 B.n440 B.n438 163.367
R1612 B.n436 B.n166 163.367
R1613 B.n432 B.n430 163.367
R1614 B.n428 B.n168 163.367
R1615 B.n424 B.n422 163.367
R1616 B.n420 B.n170 163.367
R1617 B.n416 B.n414 163.367
R1618 B.n412 B.n172 163.367
R1619 B.n408 B.n406 163.367
R1620 B.n404 B.n174 163.367
R1621 B.n400 B.n398 163.367
R1622 B.n396 B.n176 163.367
R1623 B.n392 B.n390 163.367
R1624 B.n388 B.n178 163.367
R1625 B.n384 B.n382 163.367
R1626 B.n380 B.n180 163.367
R1627 B.n376 B.n374 163.367
R1628 B.n372 B.n182 163.367
R1629 B.n368 B.n366 163.367
R1630 B.n364 B.n184 163.367
R1631 B.n359 B.n357 163.367
R1632 B.n355 B.n188 163.367
R1633 B.n351 B.n349 163.367
R1634 B.n347 B.n190 163.367
R1635 B.n343 B.n341 163.367
R1636 B.n338 B.n337 163.367
R1637 B.n335 B.n196 163.367
R1638 B.n331 B.n329 163.367
R1639 B.n327 B.n198 163.367
R1640 B.n323 B.n321 163.367
R1641 B.n319 B.n200 163.367
R1642 B.n315 B.n313 163.367
R1643 B.n311 B.n202 163.367
R1644 B.n307 B.n305 163.367
R1645 B.n303 B.n204 163.367
R1646 B.n299 B.n297 163.367
R1647 B.n295 B.n206 163.367
R1648 B.n291 B.n289 163.367
R1649 B.n287 B.n208 163.367
R1650 B.n283 B.n281 163.367
R1651 B.n279 B.n210 163.367
R1652 B.n275 B.n273 163.367
R1653 B.n271 B.n212 163.367
R1654 B.n267 B.n265 163.367
R1655 B.n263 B.n214 163.367
R1656 B.n259 B.n257 163.367
R1657 B.n255 B.n216 163.367
R1658 B.n251 B.n249 163.367
R1659 B.n247 B.n218 163.367
R1660 B.n243 B.n241 163.367
R1661 B.n239 B.n220 163.367
R1662 B.n235 B.n233 163.367
R1663 B.n231 B.n222 163.367
R1664 B.n227 B.n225 163.367
R1665 B.n483 B.n150 163.367
R1666 B.n487 B.n150 163.367
R1667 B.n487 B.n143 163.367
R1668 B.n495 B.n143 163.367
R1669 B.n495 B.n141 163.367
R1670 B.n499 B.n141 163.367
R1671 B.n499 B.n136 163.367
R1672 B.n507 B.n136 163.367
R1673 B.n507 B.n134 163.367
R1674 B.n511 B.n134 163.367
R1675 B.n511 B.n129 163.367
R1676 B.n520 B.n129 163.367
R1677 B.n520 B.n127 163.367
R1678 B.n524 B.n127 163.367
R1679 B.n524 B.n122 163.367
R1680 B.n533 B.n122 163.367
R1681 B.n533 B.n120 163.367
R1682 B.n538 B.n120 163.367
R1683 B.n538 B.n114 163.367
R1684 B.n546 B.n114 163.367
R1685 B.n547 B.n546 163.367
R1686 B.n547 B.n5 163.367
R1687 B.n6 B.n5 163.367
R1688 B.n7 B.n6 163.367
R1689 B.n552 B.n7 163.367
R1690 B.n552 B.n12 163.367
R1691 B.n13 B.n12 163.367
R1692 B.n14 B.n13 163.367
R1693 B.n557 B.n14 163.367
R1694 B.n557 B.n19 163.367
R1695 B.n20 B.n19 163.367
R1696 B.n21 B.n20 163.367
R1697 B.n562 B.n21 163.367
R1698 B.n562 B.n26 163.367
R1699 B.n27 B.n26 163.367
R1700 B.n28 B.n27 163.367
R1701 B.n567 B.n28 163.367
R1702 B.n567 B.n33 163.367
R1703 B.n34 B.n33 163.367
R1704 B.n35 B.n34 163.367
R1705 B.n572 B.n35 163.367
R1706 B.n572 B.n40 163.367
R1707 B.n41 B.n40 163.367
R1708 B.n42 B.n41 163.367
R1709 B.n833 B.n831 163.367
R1710 B.n829 B.n46 163.367
R1711 B.n825 B.n823 163.367
R1712 B.n821 B.n48 163.367
R1713 B.n817 B.n815 163.367
R1714 B.n813 B.n50 163.367
R1715 B.n809 B.n807 163.367
R1716 B.n805 B.n52 163.367
R1717 B.n801 B.n799 163.367
R1718 B.n797 B.n54 163.367
R1719 B.n793 B.n791 163.367
R1720 B.n789 B.n56 163.367
R1721 B.n785 B.n783 163.367
R1722 B.n781 B.n58 163.367
R1723 B.n777 B.n775 163.367
R1724 B.n773 B.n60 163.367
R1725 B.n769 B.n767 163.367
R1726 B.n765 B.n62 163.367
R1727 B.n761 B.n759 163.367
R1728 B.n757 B.n64 163.367
R1729 B.n753 B.n751 163.367
R1730 B.n749 B.n66 163.367
R1731 B.n745 B.n743 163.367
R1732 B.n741 B.n68 163.367
R1733 B.n737 B.n735 163.367
R1734 B.n733 B.n70 163.367
R1735 B.n729 B.n727 163.367
R1736 B.n725 B.n72 163.367
R1737 B.n721 B.n719 163.367
R1738 B.n717 B.n74 163.367
R1739 B.n712 B.n710 163.367
R1740 B.n708 B.n78 163.367
R1741 B.n704 B.n702 163.367
R1742 B.n700 B.n80 163.367
R1743 B.n695 B.n693 163.367
R1744 B.n691 B.n84 163.367
R1745 B.n687 B.n685 163.367
R1746 B.n683 B.n86 163.367
R1747 B.n679 B.n677 163.367
R1748 B.n675 B.n88 163.367
R1749 B.n671 B.n669 163.367
R1750 B.n667 B.n90 163.367
R1751 B.n663 B.n661 163.367
R1752 B.n659 B.n92 163.367
R1753 B.n655 B.n653 163.367
R1754 B.n651 B.n94 163.367
R1755 B.n647 B.n645 163.367
R1756 B.n643 B.n96 163.367
R1757 B.n639 B.n637 163.367
R1758 B.n635 B.n98 163.367
R1759 B.n631 B.n629 163.367
R1760 B.n627 B.n100 163.367
R1761 B.n623 B.n621 163.367
R1762 B.n619 B.n102 163.367
R1763 B.n615 B.n613 163.367
R1764 B.n611 B.n104 163.367
R1765 B.n607 B.n605 163.367
R1766 B.n603 B.n106 163.367
R1767 B.n599 B.n597 163.367
R1768 B.n595 B.n108 163.367
R1769 B.n591 B.n589 163.367
R1770 B.n587 B.n110 163.367
R1771 B.n583 B.n581 163.367
R1772 B.n579 B.n112 163.367
R1773 B.n476 B.n154 71.676
R1774 B.n474 B.n156 71.676
R1775 B.n470 B.n469 71.676
R1776 B.n463 B.n158 71.676
R1777 B.n462 B.n461 71.676
R1778 B.n455 B.n160 71.676
R1779 B.n454 B.n453 71.676
R1780 B.n447 B.n162 71.676
R1781 B.n446 B.n445 71.676
R1782 B.n439 B.n164 71.676
R1783 B.n438 B.n437 71.676
R1784 B.n431 B.n166 71.676
R1785 B.n430 B.n429 71.676
R1786 B.n423 B.n168 71.676
R1787 B.n422 B.n421 71.676
R1788 B.n415 B.n170 71.676
R1789 B.n414 B.n413 71.676
R1790 B.n407 B.n172 71.676
R1791 B.n406 B.n405 71.676
R1792 B.n399 B.n174 71.676
R1793 B.n398 B.n397 71.676
R1794 B.n391 B.n176 71.676
R1795 B.n390 B.n389 71.676
R1796 B.n383 B.n178 71.676
R1797 B.n382 B.n381 71.676
R1798 B.n375 B.n180 71.676
R1799 B.n374 B.n373 71.676
R1800 B.n367 B.n182 71.676
R1801 B.n366 B.n365 71.676
R1802 B.n358 B.n184 71.676
R1803 B.n357 B.n356 71.676
R1804 B.n350 B.n188 71.676
R1805 B.n349 B.n348 71.676
R1806 B.n342 B.n190 71.676
R1807 B.n341 B.n194 71.676
R1808 B.n337 B.n336 71.676
R1809 B.n330 B.n196 71.676
R1810 B.n329 B.n328 71.676
R1811 B.n322 B.n198 71.676
R1812 B.n321 B.n320 71.676
R1813 B.n314 B.n200 71.676
R1814 B.n313 B.n312 71.676
R1815 B.n306 B.n202 71.676
R1816 B.n305 B.n304 71.676
R1817 B.n298 B.n204 71.676
R1818 B.n297 B.n296 71.676
R1819 B.n290 B.n206 71.676
R1820 B.n289 B.n288 71.676
R1821 B.n282 B.n208 71.676
R1822 B.n281 B.n280 71.676
R1823 B.n274 B.n210 71.676
R1824 B.n273 B.n272 71.676
R1825 B.n266 B.n212 71.676
R1826 B.n265 B.n264 71.676
R1827 B.n258 B.n214 71.676
R1828 B.n257 B.n256 71.676
R1829 B.n250 B.n216 71.676
R1830 B.n249 B.n248 71.676
R1831 B.n242 B.n218 71.676
R1832 B.n241 B.n240 71.676
R1833 B.n234 B.n220 71.676
R1834 B.n233 B.n232 71.676
R1835 B.n226 B.n222 71.676
R1836 B.n225 B.n224 71.676
R1837 B.n832 B.n44 71.676
R1838 B.n831 B.n830 71.676
R1839 B.n824 B.n46 71.676
R1840 B.n823 B.n822 71.676
R1841 B.n816 B.n48 71.676
R1842 B.n815 B.n814 71.676
R1843 B.n808 B.n50 71.676
R1844 B.n807 B.n806 71.676
R1845 B.n800 B.n52 71.676
R1846 B.n799 B.n798 71.676
R1847 B.n792 B.n54 71.676
R1848 B.n791 B.n790 71.676
R1849 B.n784 B.n56 71.676
R1850 B.n783 B.n782 71.676
R1851 B.n776 B.n58 71.676
R1852 B.n775 B.n774 71.676
R1853 B.n768 B.n60 71.676
R1854 B.n767 B.n766 71.676
R1855 B.n760 B.n62 71.676
R1856 B.n759 B.n758 71.676
R1857 B.n752 B.n64 71.676
R1858 B.n751 B.n750 71.676
R1859 B.n744 B.n66 71.676
R1860 B.n743 B.n742 71.676
R1861 B.n736 B.n68 71.676
R1862 B.n735 B.n734 71.676
R1863 B.n728 B.n70 71.676
R1864 B.n727 B.n726 71.676
R1865 B.n720 B.n72 71.676
R1866 B.n719 B.n718 71.676
R1867 B.n711 B.n74 71.676
R1868 B.n710 B.n709 71.676
R1869 B.n703 B.n78 71.676
R1870 B.n702 B.n701 71.676
R1871 B.n694 B.n80 71.676
R1872 B.n693 B.n692 71.676
R1873 B.n686 B.n84 71.676
R1874 B.n685 B.n684 71.676
R1875 B.n678 B.n86 71.676
R1876 B.n677 B.n676 71.676
R1877 B.n670 B.n88 71.676
R1878 B.n669 B.n668 71.676
R1879 B.n662 B.n90 71.676
R1880 B.n661 B.n660 71.676
R1881 B.n654 B.n92 71.676
R1882 B.n653 B.n652 71.676
R1883 B.n646 B.n94 71.676
R1884 B.n645 B.n644 71.676
R1885 B.n638 B.n96 71.676
R1886 B.n637 B.n636 71.676
R1887 B.n630 B.n98 71.676
R1888 B.n629 B.n628 71.676
R1889 B.n622 B.n100 71.676
R1890 B.n621 B.n620 71.676
R1891 B.n614 B.n102 71.676
R1892 B.n613 B.n612 71.676
R1893 B.n606 B.n104 71.676
R1894 B.n605 B.n604 71.676
R1895 B.n598 B.n106 71.676
R1896 B.n597 B.n596 71.676
R1897 B.n590 B.n108 71.676
R1898 B.n589 B.n588 71.676
R1899 B.n582 B.n110 71.676
R1900 B.n581 B.n580 71.676
R1901 B.n580 B.n579 71.676
R1902 B.n583 B.n582 71.676
R1903 B.n588 B.n587 71.676
R1904 B.n591 B.n590 71.676
R1905 B.n596 B.n595 71.676
R1906 B.n599 B.n598 71.676
R1907 B.n604 B.n603 71.676
R1908 B.n607 B.n606 71.676
R1909 B.n612 B.n611 71.676
R1910 B.n615 B.n614 71.676
R1911 B.n620 B.n619 71.676
R1912 B.n623 B.n622 71.676
R1913 B.n628 B.n627 71.676
R1914 B.n631 B.n630 71.676
R1915 B.n636 B.n635 71.676
R1916 B.n639 B.n638 71.676
R1917 B.n644 B.n643 71.676
R1918 B.n647 B.n646 71.676
R1919 B.n652 B.n651 71.676
R1920 B.n655 B.n654 71.676
R1921 B.n660 B.n659 71.676
R1922 B.n663 B.n662 71.676
R1923 B.n668 B.n667 71.676
R1924 B.n671 B.n670 71.676
R1925 B.n676 B.n675 71.676
R1926 B.n679 B.n678 71.676
R1927 B.n684 B.n683 71.676
R1928 B.n687 B.n686 71.676
R1929 B.n692 B.n691 71.676
R1930 B.n695 B.n694 71.676
R1931 B.n701 B.n700 71.676
R1932 B.n704 B.n703 71.676
R1933 B.n709 B.n708 71.676
R1934 B.n712 B.n711 71.676
R1935 B.n718 B.n717 71.676
R1936 B.n721 B.n720 71.676
R1937 B.n726 B.n725 71.676
R1938 B.n729 B.n728 71.676
R1939 B.n734 B.n733 71.676
R1940 B.n737 B.n736 71.676
R1941 B.n742 B.n741 71.676
R1942 B.n745 B.n744 71.676
R1943 B.n750 B.n749 71.676
R1944 B.n753 B.n752 71.676
R1945 B.n758 B.n757 71.676
R1946 B.n761 B.n760 71.676
R1947 B.n766 B.n765 71.676
R1948 B.n769 B.n768 71.676
R1949 B.n774 B.n773 71.676
R1950 B.n777 B.n776 71.676
R1951 B.n782 B.n781 71.676
R1952 B.n785 B.n784 71.676
R1953 B.n790 B.n789 71.676
R1954 B.n793 B.n792 71.676
R1955 B.n798 B.n797 71.676
R1956 B.n801 B.n800 71.676
R1957 B.n806 B.n805 71.676
R1958 B.n809 B.n808 71.676
R1959 B.n814 B.n813 71.676
R1960 B.n817 B.n816 71.676
R1961 B.n822 B.n821 71.676
R1962 B.n825 B.n824 71.676
R1963 B.n830 B.n829 71.676
R1964 B.n833 B.n832 71.676
R1965 B.n477 B.n476 71.676
R1966 B.n471 B.n156 71.676
R1967 B.n469 B.n468 71.676
R1968 B.n464 B.n463 71.676
R1969 B.n461 B.n460 71.676
R1970 B.n456 B.n455 71.676
R1971 B.n453 B.n452 71.676
R1972 B.n448 B.n447 71.676
R1973 B.n445 B.n444 71.676
R1974 B.n440 B.n439 71.676
R1975 B.n437 B.n436 71.676
R1976 B.n432 B.n431 71.676
R1977 B.n429 B.n428 71.676
R1978 B.n424 B.n423 71.676
R1979 B.n421 B.n420 71.676
R1980 B.n416 B.n415 71.676
R1981 B.n413 B.n412 71.676
R1982 B.n408 B.n407 71.676
R1983 B.n405 B.n404 71.676
R1984 B.n400 B.n399 71.676
R1985 B.n397 B.n396 71.676
R1986 B.n392 B.n391 71.676
R1987 B.n389 B.n388 71.676
R1988 B.n384 B.n383 71.676
R1989 B.n381 B.n380 71.676
R1990 B.n376 B.n375 71.676
R1991 B.n373 B.n372 71.676
R1992 B.n368 B.n367 71.676
R1993 B.n365 B.n364 71.676
R1994 B.n359 B.n358 71.676
R1995 B.n356 B.n355 71.676
R1996 B.n351 B.n350 71.676
R1997 B.n348 B.n347 71.676
R1998 B.n343 B.n342 71.676
R1999 B.n338 B.n194 71.676
R2000 B.n336 B.n335 71.676
R2001 B.n331 B.n330 71.676
R2002 B.n328 B.n327 71.676
R2003 B.n323 B.n322 71.676
R2004 B.n320 B.n319 71.676
R2005 B.n315 B.n314 71.676
R2006 B.n312 B.n311 71.676
R2007 B.n307 B.n306 71.676
R2008 B.n304 B.n303 71.676
R2009 B.n299 B.n298 71.676
R2010 B.n296 B.n295 71.676
R2011 B.n291 B.n290 71.676
R2012 B.n288 B.n287 71.676
R2013 B.n283 B.n282 71.676
R2014 B.n280 B.n279 71.676
R2015 B.n275 B.n274 71.676
R2016 B.n272 B.n271 71.676
R2017 B.n267 B.n266 71.676
R2018 B.n264 B.n263 71.676
R2019 B.n259 B.n258 71.676
R2020 B.n256 B.n255 71.676
R2021 B.n251 B.n250 71.676
R2022 B.n248 B.n247 71.676
R2023 B.n243 B.n242 71.676
R2024 B.n240 B.n239 71.676
R2025 B.n235 B.n234 71.676
R2026 B.n232 B.n231 71.676
R2027 B.n227 B.n226 71.676
R2028 B.n224 B.n152 71.676
R2029 B.n193 B.n192 59.5399
R2030 B.n361 B.n186 59.5399
R2031 B.n715 B.n76 59.5399
R2032 B.n697 B.n82 59.5399
R2033 B.n482 B.n153 53.8647
R2034 B.n838 B.n43 53.8647
R2035 B.n836 B.n835 32.9371
R2036 B.n577 B.n576 32.9371
R2037 B.n484 B.n151 32.9371
R2038 B.n480 B.n479 32.9371
R2039 B.n482 B.n149 31.8506
R2040 B.n488 B.n149 31.8506
R2041 B.n488 B.n144 31.8506
R2042 B.n494 B.n144 31.8506
R2043 B.n494 B.n145 31.8506
R2044 B.n500 B.n137 31.8506
R2045 B.n506 B.n137 31.8506
R2046 B.n506 B.n133 31.8506
R2047 B.n513 B.n133 31.8506
R2048 B.n513 B.n512 31.8506
R2049 B.n519 B.n126 31.8506
R2050 B.n526 B.n126 31.8506
R2051 B.n526 B.n525 31.8506
R2052 B.n532 B.n119 31.8506
R2053 B.n539 B.n119 31.8506
R2054 B.n545 B.n115 31.8506
R2055 B.n545 B.n4 31.8506
R2056 B.n880 B.n4 31.8506
R2057 B.n880 B.n879 31.8506
R2058 B.n879 B.n878 31.8506
R2059 B.n878 B.n8 31.8506
R2060 B.n872 B.n871 31.8506
R2061 B.n871 B.n870 31.8506
R2062 B.n864 B.n18 31.8506
R2063 B.n864 B.n863 31.8506
R2064 B.n863 B.n862 31.8506
R2065 B.n856 B.n25 31.8506
R2066 B.n856 B.n855 31.8506
R2067 B.n855 B.n854 31.8506
R2068 B.n854 B.n29 31.8506
R2069 B.n848 B.n29 31.8506
R2070 B.n847 B.n846 31.8506
R2071 B.n846 B.n36 31.8506
R2072 B.n840 B.n36 31.8506
R2073 B.n840 B.n839 31.8506
R2074 B.n839 B.n838 31.8506
R2075 B.n500 B.t7 27.1668
R2076 B.n848 B.t11 27.1668
R2077 B.n512 B.t4 25.2932
R2078 B.n25 B.t2 25.2932
R2079 B.n532 B.t0 24.3565
R2080 B.n870 B.t3 24.3565
R2081 B.n192 B.n191 22.6914
R2082 B.n186 B.n185 22.6914
R2083 B.n76 B.n75 22.6914
R2084 B.n82 B.n81 22.6914
R2085 B.n539 B.t1 21.5462
R2086 B.n872 B.t5 21.5462
R2087 B B.n882 18.0485
R2088 B.n835 B.n834 10.6151
R2089 B.n834 B.n45 10.6151
R2090 B.n828 B.n45 10.6151
R2091 B.n828 B.n827 10.6151
R2092 B.n827 B.n826 10.6151
R2093 B.n826 B.n47 10.6151
R2094 B.n820 B.n47 10.6151
R2095 B.n820 B.n819 10.6151
R2096 B.n819 B.n818 10.6151
R2097 B.n818 B.n49 10.6151
R2098 B.n812 B.n49 10.6151
R2099 B.n812 B.n811 10.6151
R2100 B.n811 B.n810 10.6151
R2101 B.n810 B.n51 10.6151
R2102 B.n804 B.n51 10.6151
R2103 B.n804 B.n803 10.6151
R2104 B.n803 B.n802 10.6151
R2105 B.n802 B.n53 10.6151
R2106 B.n796 B.n53 10.6151
R2107 B.n796 B.n795 10.6151
R2108 B.n795 B.n794 10.6151
R2109 B.n794 B.n55 10.6151
R2110 B.n788 B.n55 10.6151
R2111 B.n788 B.n787 10.6151
R2112 B.n787 B.n786 10.6151
R2113 B.n786 B.n57 10.6151
R2114 B.n780 B.n57 10.6151
R2115 B.n780 B.n779 10.6151
R2116 B.n779 B.n778 10.6151
R2117 B.n778 B.n59 10.6151
R2118 B.n772 B.n59 10.6151
R2119 B.n772 B.n771 10.6151
R2120 B.n771 B.n770 10.6151
R2121 B.n770 B.n61 10.6151
R2122 B.n764 B.n61 10.6151
R2123 B.n764 B.n763 10.6151
R2124 B.n763 B.n762 10.6151
R2125 B.n762 B.n63 10.6151
R2126 B.n756 B.n63 10.6151
R2127 B.n756 B.n755 10.6151
R2128 B.n755 B.n754 10.6151
R2129 B.n754 B.n65 10.6151
R2130 B.n748 B.n65 10.6151
R2131 B.n748 B.n747 10.6151
R2132 B.n747 B.n746 10.6151
R2133 B.n746 B.n67 10.6151
R2134 B.n740 B.n67 10.6151
R2135 B.n740 B.n739 10.6151
R2136 B.n739 B.n738 10.6151
R2137 B.n738 B.n69 10.6151
R2138 B.n732 B.n69 10.6151
R2139 B.n732 B.n731 10.6151
R2140 B.n731 B.n730 10.6151
R2141 B.n730 B.n71 10.6151
R2142 B.n724 B.n71 10.6151
R2143 B.n724 B.n723 10.6151
R2144 B.n723 B.n722 10.6151
R2145 B.n722 B.n73 10.6151
R2146 B.n716 B.n73 10.6151
R2147 B.n714 B.n713 10.6151
R2148 B.n713 B.n77 10.6151
R2149 B.n707 B.n77 10.6151
R2150 B.n707 B.n706 10.6151
R2151 B.n706 B.n705 10.6151
R2152 B.n705 B.n79 10.6151
R2153 B.n699 B.n79 10.6151
R2154 B.n699 B.n698 10.6151
R2155 B.n696 B.n83 10.6151
R2156 B.n690 B.n83 10.6151
R2157 B.n690 B.n689 10.6151
R2158 B.n689 B.n688 10.6151
R2159 B.n688 B.n85 10.6151
R2160 B.n682 B.n85 10.6151
R2161 B.n682 B.n681 10.6151
R2162 B.n681 B.n680 10.6151
R2163 B.n680 B.n87 10.6151
R2164 B.n674 B.n87 10.6151
R2165 B.n674 B.n673 10.6151
R2166 B.n673 B.n672 10.6151
R2167 B.n672 B.n89 10.6151
R2168 B.n666 B.n89 10.6151
R2169 B.n666 B.n665 10.6151
R2170 B.n665 B.n664 10.6151
R2171 B.n664 B.n91 10.6151
R2172 B.n658 B.n91 10.6151
R2173 B.n658 B.n657 10.6151
R2174 B.n657 B.n656 10.6151
R2175 B.n656 B.n93 10.6151
R2176 B.n650 B.n93 10.6151
R2177 B.n650 B.n649 10.6151
R2178 B.n649 B.n648 10.6151
R2179 B.n648 B.n95 10.6151
R2180 B.n642 B.n95 10.6151
R2181 B.n642 B.n641 10.6151
R2182 B.n641 B.n640 10.6151
R2183 B.n640 B.n97 10.6151
R2184 B.n634 B.n97 10.6151
R2185 B.n634 B.n633 10.6151
R2186 B.n633 B.n632 10.6151
R2187 B.n632 B.n99 10.6151
R2188 B.n626 B.n99 10.6151
R2189 B.n626 B.n625 10.6151
R2190 B.n625 B.n624 10.6151
R2191 B.n624 B.n101 10.6151
R2192 B.n618 B.n101 10.6151
R2193 B.n618 B.n617 10.6151
R2194 B.n617 B.n616 10.6151
R2195 B.n616 B.n103 10.6151
R2196 B.n610 B.n103 10.6151
R2197 B.n610 B.n609 10.6151
R2198 B.n609 B.n608 10.6151
R2199 B.n608 B.n105 10.6151
R2200 B.n602 B.n105 10.6151
R2201 B.n602 B.n601 10.6151
R2202 B.n601 B.n600 10.6151
R2203 B.n600 B.n107 10.6151
R2204 B.n594 B.n107 10.6151
R2205 B.n594 B.n593 10.6151
R2206 B.n593 B.n592 10.6151
R2207 B.n592 B.n109 10.6151
R2208 B.n586 B.n109 10.6151
R2209 B.n586 B.n585 10.6151
R2210 B.n585 B.n584 10.6151
R2211 B.n584 B.n111 10.6151
R2212 B.n578 B.n111 10.6151
R2213 B.n578 B.n577 10.6151
R2214 B.n485 B.n484 10.6151
R2215 B.n486 B.n485 10.6151
R2216 B.n486 B.n142 10.6151
R2217 B.n496 B.n142 10.6151
R2218 B.n497 B.n496 10.6151
R2219 B.n498 B.n497 10.6151
R2220 B.n498 B.n135 10.6151
R2221 B.n508 B.n135 10.6151
R2222 B.n509 B.n508 10.6151
R2223 B.n510 B.n509 10.6151
R2224 B.n510 B.n128 10.6151
R2225 B.n521 B.n128 10.6151
R2226 B.n522 B.n521 10.6151
R2227 B.n523 B.n522 10.6151
R2228 B.n523 B.n121 10.6151
R2229 B.n534 B.n121 10.6151
R2230 B.n535 B.n534 10.6151
R2231 B.n537 B.n535 10.6151
R2232 B.n537 B.n536 10.6151
R2233 B.n536 B.n113 10.6151
R2234 B.n548 B.n113 10.6151
R2235 B.n549 B.n548 10.6151
R2236 B.n550 B.n549 10.6151
R2237 B.n551 B.n550 10.6151
R2238 B.n553 B.n551 10.6151
R2239 B.n554 B.n553 10.6151
R2240 B.n555 B.n554 10.6151
R2241 B.n556 B.n555 10.6151
R2242 B.n558 B.n556 10.6151
R2243 B.n559 B.n558 10.6151
R2244 B.n560 B.n559 10.6151
R2245 B.n561 B.n560 10.6151
R2246 B.n563 B.n561 10.6151
R2247 B.n564 B.n563 10.6151
R2248 B.n565 B.n564 10.6151
R2249 B.n566 B.n565 10.6151
R2250 B.n568 B.n566 10.6151
R2251 B.n569 B.n568 10.6151
R2252 B.n570 B.n569 10.6151
R2253 B.n571 B.n570 10.6151
R2254 B.n573 B.n571 10.6151
R2255 B.n574 B.n573 10.6151
R2256 B.n575 B.n574 10.6151
R2257 B.n576 B.n575 10.6151
R2258 B.n479 B.n478 10.6151
R2259 B.n478 B.n155 10.6151
R2260 B.n473 B.n155 10.6151
R2261 B.n473 B.n472 10.6151
R2262 B.n472 B.n157 10.6151
R2263 B.n467 B.n157 10.6151
R2264 B.n467 B.n466 10.6151
R2265 B.n466 B.n465 10.6151
R2266 B.n465 B.n159 10.6151
R2267 B.n459 B.n159 10.6151
R2268 B.n459 B.n458 10.6151
R2269 B.n458 B.n457 10.6151
R2270 B.n457 B.n161 10.6151
R2271 B.n451 B.n161 10.6151
R2272 B.n451 B.n450 10.6151
R2273 B.n450 B.n449 10.6151
R2274 B.n449 B.n163 10.6151
R2275 B.n443 B.n163 10.6151
R2276 B.n443 B.n442 10.6151
R2277 B.n442 B.n441 10.6151
R2278 B.n441 B.n165 10.6151
R2279 B.n435 B.n165 10.6151
R2280 B.n435 B.n434 10.6151
R2281 B.n434 B.n433 10.6151
R2282 B.n433 B.n167 10.6151
R2283 B.n427 B.n167 10.6151
R2284 B.n427 B.n426 10.6151
R2285 B.n426 B.n425 10.6151
R2286 B.n425 B.n169 10.6151
R2287 B.n419 B.n169 10.6151
R2288 B.n419 B.n418 10.6151
R2289 B.n418 B.n417 10.6151
R2290 B.n417 B.n171 10.6151
R2291 B.n411 B.n171 10.6151
R2292 B.n411 B.n410 10.6151
R2293 B.n410 B.n409 10.6151
R2294 B.n409 B.n173 10.6151
R2295 B.n403 B.n173 10.6151
R2296 B.n403 B.n402 10.6151
R2297 B.n402 B.n401 10.6151
R2298 B.n401 B.n175 10.6151
R2299 B.n395 B.n175 10.6151
R2300 B.n395 B.n394 10.6151
R2301 B.n394 B.n393 10.6151
R2302 B.n393 B.n177 10.6151
R2303 B.n387 B.n177 10.6151
R2304 B.n387 B.n386 10.6151
R2305 B.n386 B.n385 10.6151
R2306 B.n385 B.n179 10.6151
R2307 B.n379 B.n179 10.6151
R2308 B.n379 B.n378 10.6151
R2309 B.n378 B.n377 10.6151
R2310 B.n377 B.n181 10.6151
R2311 B.n371 B.n181 10.6151
R2312 B.n371 B.n370 10.6151
R2313 B.n370 B.n369 10.6151
R2314 B.n369 B.n183 10.6151
R2315 B.n363 B.n183 10.6151
R2316 B.n363 B.n362 10.6151
R2317 B.n360 B.n187 10.6151
R2318 B.n354 B.n187 10.6151
R2319 B.n354 B.n353 10.6151
R2320 B.n353 B.n352 10.6151
R2321 B.n352 B.n189 10.6151
R2322 B.n346 B.n189 10.6151
R2323 B.n346 B.n345 10.6151
R2324 B.n345 B.n344 10.6151
R2325 B.n340 B.n339 10.6151
R2326 B.n339 B.n195 10.6151
R2327 B.n334 B.n195 10.6151
R2328 B.n334 B.n333 10.6151
R2329 B.n333 B.n332 10.6151
R2330 B.n332 B.n197 10.6151
R2331 B.n326 B.n197 10.6151
R2332 B.n326 B.n325 10.6151
R2333 B.n325 B.n324 10.6151
R2334 B.n324 B.n199 10.6151
R2335 B.n318 B.n199 10.6151
R2336 B.n318 B.n317 10.6151
R2337 B.n317 B.n316 10.6151
R2338 B.n316 B.n201 10.6151
R2339 B.n310 B.n201 10.6151
R2340 B.n310 B.n309 10.6151
R2341 B.n309 B.n308 10.6151
R2342 B.n308 B.n203 10.6151
R2343 B.n302 B.n203 10.6151
R2344 B.n302 B.n301 10.6151
R2345 B.n301 B.n300 10.6151
R2346 B.n300 B.n205 10.6151
R2347 B.n294 B.n205 10.6151
R2348 B.n294 B.n293 10.6151
R2349 B.n293 B.n292 10.6151
R2350 B.n292 B.n207 10.6151
R2351 B.n286 B.n207 10.6151
R2352 B.n286 B.n285 10.6151
R2353 B.n285 B.n284 10.6151
R2354 B.n284 B.n209 10.6151
R2355 B.n278 B.n209 10.6151
R2356 B.n278 B.n277 10.6151
R2357 B.n277 B.n276 10.6151
R2358 B.n276 B.n211 10.6151
R2359 B.n270 B.n211 10.6151
R2360 B.n270 B.n269 10.6151
R2361 B.n269 B.n268 10.6151
R2362 B.n268 B.n213 10.6151
R2363 B.n262 B.n213 10.6151
R2364 B.n262 B.n261 10.6151
R2365 B.n261 B.n260 10.6151
R2366 B.n260 B.n215 10.6151
R2367 B.n254 B.n215 10.6151
R2368 B.n254 B.n253 10.6151
R2369 B.n253 B.n252 10.6151
R2370 B.n252 B.n217 10.6151
R2371 B.n246 B.n217 10.6151
R2372 B.n246 B.n245 10.6151
R2373 B.n245 B.n244 10.6151
R2374 B.n244 B.n219 10.6151
R2375 B.n238 B.n219 10.6151
R2376 B.n238 B.n237 10.6151
R2377 B.n237 B.n236 10.6151
R2378 B.n236 B.n221 10.6151
R2379 B.n230 B.n221 10.6151
R2380 B.n230 B.n229 10.6151
R2381 B.n229 B.n228 10.6151
R2382 B.n228 B.n223 10.6151
R2383 B.n223 B.n151 10.6151
R2384 B.n480 B.n147 10.6151
R2385 B.n490 B.n147 10.6151
R2386 B.n491 B.n490 10.6151
R2387 B.n492 B.n491 10.6151
R2388 B.n492 B.n139 10.6151
R2389 B.n502 B.n139 10.6151
R2390 B.n503 B.n502 10.6151
R2391 B.n504 B.n503 10.6151
R2392 B.n504 B.n131 10.6151
R2393 B.n515 B.n131 10.6151
R2394 B.n516 B.n515 10.6151
R2395 B.n517 B.n516 10.6151
R2396 B.n517 B.n124 10.6151
R2397 B.n528 B.n124 10.6151
R2398 B.n529 B.n528 10.6151
R2399 B.n530 B.n529 10.6151
R2400 B.n530 B.n117 10.6151
R2401 B.n541 B.n117 10.6151
R2402 B.n542 B.n541 10.6151
R2403 B.n543 B.n542 10.6151
R2404 B.n543 B.n0 10.6151
R2405 B.n876 B.n1 10.6151
R2406 B.n876 B.n875 10.6151
R2407 B.n875 B.n874 10.6151
R2408 B.n874 B.n10 10.6151
R2409 B.n868 B.n10 10.6151
R2410 B.n868 B.n867 10.6151
R2411 B.n867 B.n866 10.6151
R2412 B.n866 B.n16 10.6151
R2413 B.n860 B.n16 10.6151
R2414 B.n860 B.n859 10.6151
R2415 B.n859 B.n858 10.6151
R2416 B.n858 B.n23 10.6151
R2417 B.n852 B.n23 10.6151
R2418 B.n852 B.n851 10.6151
R2419 B.n851 B.n850 10.6151
R2420 B.n850 B.n31 10.6151
R2421 B.n844 B.n31 10.6151
R2422 B.n844 B.n843 10.6151
R2423 B.n843 B.n842 10.6151
R2424 B.n842 B.n38 10.6151
R2425 B.n836 B.n38 10.6151
R2426 B.t1 B.n115 10.3049
R2427 B.t5 B.n8 10.3049
R2428 B.n525 B.t0 7.49464
R2429 B.n18 B.t3 7.49464
R2430 B.n519 B.t4 6.55788
R2431 B.n862 B.t2 6.55788
R2432 B.n715 B.n714 6.5566
R2433 B.n698 B.n697 6.5566
R2434 B.n361 B.n360 6.5566
R2435 B.n344 B.n193 6.5566
R2436 B.n145 B.t7 4.68434
R2437 B.t11 B.n847 4.68434
R2438 B.n716 B.n715 4.05904
R2439 B.n697 B.n696 4.05904
R2440 B.n362 B.n361 4.05904
R2441 B.n340 B.n193 4.05904
R2442 B.n882 B.n0 2.81026
R2443 B.n882 B.n1 2.81026
R2444 VN.n1 VN.t0 584.812
R2445 VN.n7 VN.t2 584.812
R2446 VN.n4 VN.t3 569.506
R2447 VN.n10 VN.t1 569.506
R2448 VN.n2 VN.t4 522.455
R2449 VN.n8 VN.t5 522.455
R2450 VN.n9 VN.n6 161.3
R2451 VN.n3 VN.n0 161.3
R2452 VN.n11 VN.n10 80.6037
R2453 VN.n5 VN.n4 80.6037
R2454 VN.n4 VN.n3 56.5193
R2455 VN.n10 VN.n9 56.5193
R2456 VN VN.n11 46.8816
R2457 VN.n7 VN.n6 43.8694
R2458 VN.n1 VN.n0 43.8694
R2459 VN.n2 VN.n1 42.7544
R2460 VN.n8 VN.n7 42.7544
R2461 VN.n3 VN.n2 12.234
R2462 VN.n9 VN.n8 12.234
R2463 VN.n11 VN.n6 0.285035
R2464 VN.n5 VN.n0 0.285035
R2465 VN VN.n5 0.146778
R2466 VDD2.n199 VDD2.n103 289.615
R2467 VDD2.n96 VDD2.n0 289.615
R2468 VDD2.n200 VDD2.n199 185
R2469 VDD2.n198 VDD2.n197 185
R2470 VDD2.n107 VDD2.n106 185
R2471 VDD2.n192 VDD2.n191 185
R2472 VDD2.n190 VDD2.n189 185
R2473 VDD2.n111 VDD2.n110 185
R2474 VDD2.n184 VDD2.n183 185
R2475 VDD2.n182 VDD2.n113 185
R2476 VDD2.n181 VDD2.n180 185
R2477 VDD2.n116 VDD2.n114 185
R2478 VDD2.n175 VDD2.n174 185
R2479 VDD2.n173 VDD2.n172 185
R2480 VDD2.n120 VDD2.n119 185
R2481 VDD2.n167 VDD2.n166 185
R2482 VDD2.n165 VDD2.n164 185
R2483 VDD2.n124 VDD2.n123 185
R2484 VDD2.n159 VDD2.n158 185
R2485 VDD2.n157 VDD2.n156 185
R2486 VDD2.n128 VDD2.n127 185
R2487 VDD2.n151 VDD2.n150 185
R2488 VDD2.n149 VDD2.n148 185
R2489 VDD2.n132 VDD2.n131 185
R2490 VDD2.n143 VDD2.n142 185
R2491 VDD2.n141 VDD2.n140 185
R2492 VDD2.n136 VDD2.n135 185
R2493 VDD2.n32 VDD2.n31 185
R2494 VDD2.n37 VDD2.n36 185
R2495 VDD2.n39 VDD2.n38 185
R2496 VDD2.n28 VDD2.n27 185
R2497 VDD2.n45 VDD2.n44 185
R2498 VDD2.n47 VDD2.n46 185
R2499 VDD2.n24 VDD2.n23 185
R2500 VDD2.n53 VDD2.n52 185
R2501 VDD2.n55 VDD2.n54 185
R2502 VDD2.n20 VDD2.n19 185
R2503 VDD2.n61 VDD2.n60 185
R2504 VDD2.n63 VDD2.n62 185
R2505 VDD2.n16 VDD2.n15 185
R2506 VDD2.n69 VDD2.n68 185
R2507 VDD2.n71 VDD2.n70 185
R2508 VDD2.n12 VDD2.n11 185
R2509 VDD2.n78 VDD2.n77 185
R2510 VDD2.n79 VDD2.n10 185
R2511 VDD2.n81 VDD2.n80 185
R2512 VDD2.n8 VDD2.n7 185
R2513 VDD2.n87 VDD2.n86 185
R2514 VDD2.n89 VDD2.n88 185
R2515 VDD2.n4 VDD2.n3 185
R2516 VDD2.n95 VDD2.n94 185
R2517 VDD2.n97 VDD2.n96 185
R2518 VDD2.n137 VDD2.t4 147.659
R2519 VDD2.n33 VDD2.t5 147.659
R2520 VDD2.n199 VDD2.n198 104.615
R2521 VDD2.n198 VDD2.n106 104.615
R2522 VDD2.n191 VDD2.n106 104.615
R2523 VDD2.n191 VDD2.n190 104.615
R2524 VDD2.n190 VDD2.n110 104.615
R2525 VDD2.n183 VDD2.n110 104.615
R2526 VDD2.n183 VDD2.n182 104.615
R2527 VDD2.n182 VDD2.n181 104.615
R2528 VDD2.n181 VDD2.n114 104.615
R2529 VDD2.n174 VDD2.n114 104.615
R2530 VDD2.n174 VDD2.n173 104.615
R2531 VDD2.n173 VDD2.n119 104.615
R2532 VDD2.n166 VDD2.n119 104.615
R2533 VDD2.n166 VDD2.n165 104.615
R2534 VDD2.n165 VDD2.n123 104.615
R2535 VDD2.n158 VDD2.n123 104.615
R2536 VDD2.n158 VDD2.n157 104.615
R2537 VDD2.n157 VDD2.n127 104.615
R2538 VDD2.n150 VDD2.n127 104.615
R2539 VDD2.n150 VDD2.n149 104.615
R2540 VDD2.n149 VDD2.n131 104.615
R2541 VDD2.n142 VDD2.n131 104.615
R2542 VDD2.n142 VDD2.n141 104.615
R2543 VDD2.n141 VDD2.n135 104.615
R2544 VDD2.n37 VDD2.n31 104.615
R2545 VDD2.n38 VDD2.n37 104.615
R2546 VDD2.n38 VDD2.n27 104.615
R2547 VDD2.n45 VDD2.n27 104.615
R2548 VDD2.n46 VDD2.n45 104.615
R2549 VDD2.n46 VDD2.n23 104.615
R2550 VDD2.n53 VDD2.n23 104.615
R2551 VDD2.n54 VDD2.n53 104.615
R2552 VDD2.n54 VDD2.n19 104.615
R2553 VDD2.n61 VDD2.n19 104.615
R2554 VDD2.n62 VDD2.n61 104.615
R2555 VDD2.n62 VDD2.n15 104.615
R2556 VDD2.n69 VDD2.n15 104.615
R2557 VDD2.n70 VDD2.n69 104.615
R2558 VDD2.n70 VDD2.n11 104.615
R2559 VDD2.n78 VDD2.n11 104.615
R2560 VDD2.n79 VDD2.n78 104.615
R2561 VDD2.n80 VDD2.n79 104.615
R2562 VDD2.n80 VDD2.n7 104.615
R2563 VDD2.n87 VDD2.n7 104.615
R2564 VDD2.n88 VDD2.n87 104.615
R2565 VDD2.n88 VDD2.n3 104.615
R2566 VDD2.n95 VDD2.n3 104.615
R2567 VDD2.n96 VDD2.n95 104.615
R2568 VDD2.n102 VDD2.n101 60.2631
R2569 VDD2 VDD2.n205 60.2603
R2570 VDD2.t4 VDD2.n135 52.3082
R2571 VDD2.t5 VDD2.n31 52.3082
R2572 VDD2.n102 VDD2.n100 48.9834
R2573 VDD2.n204 VDD2.n203 48.2823
R2574 VDD2.n204 VDD2.n102 42.6916
R2575 VDD2.n137 VDD2.n136 15.6677
R2576 VDD2.n33 VDD2.n32 15.6677
R2577 VDD2.n184 VDD2.n113 13.1884
R2578 VDD2.n81 VDD2.n10 13.1884
R2579 VDD2.n185 VDD2.n111 12.8005
R2580 VDD2.n180 VDD2.n115 12.8005
R2581 VDD2.n140 VDD2.n139 12.8005
R2582 VDD2.n36 VDD2.n35 12.8005
R2583 VDD2.n77 VDD2.n76 12.8005
R2584 VDD2.n82 VDD2.n8 12.8005
R2585 VDD2.n189 VDD2.n188 12.0247
R2586 VDD2.n179 VDD2.n116 12.0247
R2587 VDD2.n143 VDD2.n134 12.0247
R2588 VDD2.n39 VDD2.n30 12.0247
R2589 VDD2.n75 VDD2.n12 12.0247
R2590 VDD2.n86 VDD2.n85 12.0247
R2591 VDD2.n192 VDD2.n109 11.249
R2592 VDD2.n176 VDD2.n175 11.249
R2593 VDD2.n144 VDD2.n132 11.249
R2594 VDD2.n40 VDD2.n28 11.249
R2595 VDD2.n72 VDD2.n71 11.249
R2596 VDD2.n89 VDD2.n6 11.249
R2597 VDD2.n193 VDD2.n107 10.4732
R2598 VDD2.n172 VDD2.n118 10.4732
R2599 VDD2.n148 VDD2.n147 10.4732
R2600 VDD2.n44 VDD2.n43 10.4732
R2601 VDD2.n68 VDD2.n14 10.4732
R2602 VDD2.n90 VDD2.n4 10.4732
R2603 VDD2.n197 VDD2.n196 9.69747
R2604 VDD2.n171 VDD2.n120 9.69747
R2605 VDD2.n151 VDD2.n130 9.69747
R2606 VDD2.n47 VDD2.n26 9.69747
R2607 VDD2.n67 VDD2.n16 9.69747
R2608 VDD2.n94 VDD2.n93 9.69747
R2609 VDD2.n203 VDD2.n202 9.45567
R2610 VDD2.n100 VDD2.n99 9.45567
R2611 VDD2.n163 VDD2.n162 9.3005
R2612 VDD2.n122 VDD2.n121 9.3005
R2613 VDD2.n169 VDD2.n168 9.3005
R2614 VDD2.n171 VDD2.n170 9.3005
R2615 VDD2.n118 VDD2.n117 9.3005
R2616 VDD2.n177 VDD2.n176 9.3005
R2617 VDD2.n179 VDD2.n178 9.3005
R2618 VDD2.n115 VDD2.n112 9.3005
R2619 VDD2.n202 VDD2.n201 9.3005
R2620 VDD2.n105 VDD2.n104 9.3005
R2621 VDD2.n196 VDD2.n195 9.3005
R2622 VDD2.n194 VDD2.n193 9.3005
R2623 VDD2.n109 VDD2.n108 9.3005
R2624 VDD2.n188 VDD2.n187 9.3005
R2625 VDD2.n186 VDD2.n185 9.3005
R2626 VDD2.n161 VDD2.n160 9.3005
R2627 VDD2.n126 VDD2.n125 9.3005
R2628 VDD2.n155 VDD2.n154 9.3005
R2629 VDD2.n153 VDD2.n152 9.3005
R2630 VDD2.n130 VDD2.n129 9.3005
R2631 VDD2.n147 VDD2.n146 9.3005
R2632 VDD2.n145 VDD2.n144 9.3005
R2633 VDD2.n134 VDD2.n133 9.3005
R2634 VDD2.n139 VDD2.n138 9.3005
R2635 VDD2.n99 VDD2.n98 9.3005
R2636 VDD2.n2 VDD2.n1 9.3005
R2637 VDD2.n93 VDD2.n92 9.3005
R2638 VDD2.n91 VDD2.n90 9.3005
R2639 VDD2.n6 VDD2.n5 9.3005
R2640 VDD2.n85 VDD2.n84 9.3005
R2641 VDD2.n83 VDD2.n82 9.3005
R2642 VDD2.n22 VDD2.n21 9.3005
R2643 VDD2.n51 VDD2.n50 9.3005
R2644 VDD2.n49 VDD2.n48 9.3005
R2645 VDD2.n26 VDD2.n25 9.3005
R2646 VDD2.n43 VDD2.n42 9.3005
R2647 VDD2.n41 VDD2.n40 9.3005
R2648 VDD2.n30 VDD2.n29 9.3005
R2649 VDD2.n35 VDD2.n34 9.3005
R2650 VDD2.n57 VDD2.n56 9.3005
R2651 VDD2.n59 VDD2.n58 9.3005
R2652 VDD2.n18 VDD2.n17 9.3005
R2653 VDD2.n65 VDD2.n64 9.3005
R2654 VDD2.n67 VDD2.n66 9.3005
R2655 VDD2.n14 VDD2.n13 9.3005
R2656 VDD2.n73 VDD2.n72 9.3005
R2657 VDD2.n75 VDD2.n74 9.3005
R2658 VDD2.n76 VDD2.n9 9.3005
R2659 VDD2.n200 VDD2.n105 8.92171
R2660 VDD2.n168 VDD2.n167 8.92171
R2661 VDD2.n152 VDD2.n128 8.92171
R2662 VDD2.n48 VDD2.n24 8.92171
R2663 VDD2.n64 VDD2.n63 8.92171
R2664 VDD2.n97 VDD2.n2 8.92171
R2665 VDD2.n201 VDD2.n103 8.14595
R2666 VDD2.n164 VDD2.n122 8.14595
R2667 VDD2.n156 VDD2.n155 8.14595
R2668 VDD2.n52 VDD2.n51 8.14595
R2669 VDD2.n60 VDD2.n18 8.14595
R2670 VDD2.n98 VDD2.n0 8.14595
R2671 VDD2.n163 VDD2.n124 7.3702
R2672 VDD2.n159 VDD2.n126 7.3702
R2673 VDD2.n55 VDD2.n22 7.3702
R2674 VDD2.n59 VDD2.n20 7.3702
R2675 VDD2.n160 VDD2.n124 6.59444
R2676 VDD2.n160 VDD2.n159 6.59444
R2677 VDD2.n56 VDD2.n55 6.59444
R2678 VDD2.n56 VDD2.n20 6.59444
R2679 VDD2.n203 VDD2.n103 5.81868
R2680 VDD2.n164 VDD2.n163 5.81868
R2681 VDD2.n156 VDD2.n126 5.81868
R2682 VDD2.n52 VDD2.n22 5.81868
R2683 VDD2.n60 VDD2.n59 5.81868
R2684 VDD2.n100 VDD2.n0 5.81868
R2685 VDD2.n201 VDD2.n200 5.04292
R2686 VDD2.n167 VDD2.n122 5.04292
R2687 VDD2.n155 VDD2.n128 5.04292
R2688 VDD2.n51 VDD2.n24 5.04292
R2689 VDD2.n63 VDD2.n18 5.04292
R2690 VDD2.n98 VDD2.n97 5.04292
R2691 VDD2.n138 VDD2.n137 4.38563
R2692 VDD2.n34 VDD2.n33 4.38563
R2693 VDD2.n197 VDD2.n105 4.26717
R2694 VDD2.n168 VDD2.n120 4.26717
R2695 VDD2.n152 VDD2.n151 4.26717
R2696 VDD2.n48 VDD2.n47 4.26717
R2697 VDD2.n64 VDD2.n16 4.26717
R2698 VDD2.n94 VDD2.n2 4.26717
R2699 VDD2.n196 VDD2.n107 3.49141
R2700 VDD2.n172 VDD2.n171 3.49141
R2701 VDD2.n148 VDD2.n130 3.49141
R2702 VDD2.n44 VDD2.n26 3.49141
R2703 VDD2.n68 VDD2.n67 3.49141
R2704 VDD2.n93 VDD2.n4 3.49141
R2705 VDD2.n193 VDD2.n192 2.71565
R2706 VDD2.n175 VDD2.n118 2.71565
R2707 VDD2.n147 VDD2.n132 2.71565
R2708 VDD2.n43 VDD2.n28 2.71565
R2709 VDD2.n71 VDD2.n14 2.71565
R2710 VDD2.n90 VDD2.n89 2.71565
R2711 VDD2.n189 VDD2.n109 1.93989
R2712 VDD2.n176 VDD2.n116 1.93989
R2713 VDD2.n144 VDD2.n143 1.93989
R2714 VDD2.n40 VDD2.n39 1.93989
R2715 VDD2.n72 VDD2.n12 1.93989
R2716 VDD2.n86 VDD2.n6 1.93989
R2717 VDD2.n188 VDD2.n111 1.16414
R2718 VDD2.n180 VDD2.n179 1.16414
R2719 VDD2.n140 VDD2.n134 1.16414
R2720 VDD2.n36 VDD2.n30 1.16414
R2721 VDD2.n77 VDD2.n75 1.16414
R2722 VDD2.n85 VDD2.n8 1.16414
R2723 VDD2.n205 VDD2.t0 1.08781
R2724 VDD2.n205 VDD2.t3 1.08781
R2725 VDD2.n101 VDD2.t1 1.08781
R2726 VDD2.n101 VDD2.t2 1.08781
R2727 VDD2 VDD2.n204 0.815155
R2728 VDD2.n185 VDD2.n184 0.388379
R2729 VDD2.n115 VDD2.n113 0.388379
R2730 VDD2.n139 VDD2.n136 0.388379
R2731 VDD2.n35 VDD2.n32 0.388379
R2732 VDD2.n76 VDD2.n10 0.388379
R2733 VDD2.n82 VDD2.n81 0.388379
R2734 VDD2.n202 VDD2.n104 0.155672
R2735 VDD2.n195 VDD2.n104 0.155672
R2736 VDD2.n195 VDD2.n194 0.155672
R2737 VDD2.n194 VDD2.n108 0.155672
R2738 VDD2.n187 VDD2.n108 0.155672
R2739 VDD2.n187 VDD2.n186 0.155672
R2740 VDD2.n186 VDD2.n112 0.155672
R2741 VDD2.n178 VDD2.n112 0.155672
R2742 VDD2.n178 VDD2.n177 0.155672
R2743 VDD2.n177 VDD2.n117 0.155672
R2744 VDD2.n170 VDD2.n117 0.155672
R2745 VDD2.n170 VDD2.n169 0.155672
R2746 VDD2.n169 VDD2.n121 0.155672
R2747 VDD2.n162 VDD2.n121 0.155672
R2748 VDD2.n162 VDD2.n161 0.155672
R2749 VDD2.n161 VDD2.n125 0.155672
R2750 VDD2.n154 VDD2.n125 0.155672
R2751 VDD2.n154 VDD2.n153 0.155672
R2752 VDD2.n153 VDD2.n129 0.155672
R2753 VDD2.n146 VDD2.n129 0.155672
R2754 VDD2.n146 VDD2.n145 0.155672
R2755 VDD2.n145 VDD2.n133 0.155672
R2756 VDD2.n138 VDD2.n133 0.155672
R2757 VDD2.n34 VDD2.n29 0.155672
R2758 VDD2.n41 VDD2.n29 0.155672
R2759 VDD2.n42 VDD2.n41 0.155672
R2760 VDD2.n42 VDD2.n25 0.155672
R2761 VDD2.n49 VDD2.n25 0.155672
R2762 VDD2.n50 VDD2.n49 0.155672
R2763 VDD2.n50 VDD2.n21 0.155672
R2764 VDD2.n57 VDD2.n21 0.155672
R2765 VDD2.n58 VDD2.n57 0.155672
R2766 VDD2.n58 VDD2.n17 0.155672
R2767 VDD2.n65 VDD2.n17 0.155672
R2768 VDD2.n66 VDD2.n65 0.155672
R2769 VDD2.n66 VDD2.n13 0.155672
R2770 VDD2.n73 VDD2.n13 0.155672
R2771 VDD2.n74 VDD2.n73 0.155672
R2772 VDD2.n74 VDD2.n9 0.155672
R2773 VDD2.n83 VDD2.n9 0.155672
R2774 VDD2.n84 VDD2.n83 0.155672
R2775 VDD2.n84 VDD2.n5 0.155672
R2776 VDD2.n91 VDD2.n5 0.155672
R2777 VDD2.n92 VDD2.n91 0.155672
R2778 VDD2.n92 VDD2.n1 0.155672
R2779 VDD2.n99 VDD2.n1 0.155672
C0 VN VP 6.36946f
C1 VP VDD2 0.310377f
C2 VTAIL VP 6.48523f
C3 VN VDD2 6.99314f
C4 VN VTAIL 6.47043f
C5 VP VDD1 7.14877f
C6 VTAIL VDD2 13.1361f
C7 VN VDD1 0.148383f
C8 VDD1 VDD2 0.763569f
C9 VTAIL VDD1 13.103701f
C10 VDD2 B 5.716596f
C11 VDD1 B 5.742146f
C12 VTAIL B 8.826838f
C13 VN B 8.826429f
C14 VP B 6.629613f
C15 VDD2.n0 B 0.031478f
C16 VDD2.n1 B 0.022722f
C17 VDD2.n2 B 0.01221f
C18 VDD2.n3 B 0.02886f
C19 VDD2.n4 B 0.012928f
C20 VDD2.n5 B 0.022722f
C21 VDD2.n6 B 0.01221f
C22 VDD2.n7 B 0.02886f
C23 VDD2.n8 B 0.012928f
C24 VDD2.n9 B 0.022722f
C25 VDD2.n10 B 0.012569f
C26 VDD2.n11 B 0.02886f
C27 VDD2.n12 B 0.012928f
C28 VDD2.n13 B 0.022722f
C29 VDD2.n14 B 0.01221f
C30 VDD2.n15 B 0.02886f
C31 VDD2.n16 B 0.012928f
C32 VDD2.n17 B 0.022722f
C33 VDD2.n18 B 0.01221f
C34 VDD2.n19 B 0.02886f
C35 VDD2.n20 B 0.012928f
C36 VDD2.n21 B 0.022722f
C37 VDD2.n22 B 0.01221f
C38 VDD2.n23 B 0.02886f
C39 VDD2.n24 B 0.012928f
C40 VDD2.n25 B 0.022722f
C41 VDD2.n26 B 0.01221f
C42 VDD2.n27 B 0.02886f
C43 VDD2.n28 B 0.012928f
C44 VDD2.n29 B 0.022722f
C45 VDD2.n30 B 0.01221f
C46 VDD2.n31 B 0.021645f
C47 VDD2.n32 B 0.017048f
C48 VDD2.t5 B 0.047837f
C49 VDD2.n33 B 0.166487f
C50 VDD2.n34 B 1.81262f
C51 VDD2.n35 B 0.01221f
C52 VDD2.n36 B 0.012928f
C53 VDD2.n37 B 0.02886f
C54 VDD2.n38 B 0.02886f
C55 VDD2.n39 B 0.012928f
C56 VDD2.n40 B 0.01221f
C57 VDD2.n41 B 0.022722f
C58 VDD2.n42 B 0.022722f
C59 VDD2.n43 B 0.01221f
C60 VDD2.n44 B 0.012928f
C61 VDD2.n45 B 0.02886f
C62 VDD2.n46 B 0.02886f
C63 VDD2.n47 B 0.012928f
C64 VDD2.n48 B 0.01221f
C65 VDD2.n49 B 0.022722f
C66 VDD2.n50 B 0.022722f
C67 VDD2.n51 B 0.01221f
C68 VDD2.n52 B 0.012928f
C69 VDD2.n53 B 0.02886f
C70 VDD2.n54 B 0.02886f
C71 VDD2.n55 B 0.012928f
C72 VDD2.n56 B 0.01221f
C73 VDD2.n57 B 0.022722f
C74 VDD2.n58 B 0.022722f
C75 VDD2.n59 B 0.01221f
C76 VDD2.n60 B 0.012928f
C77 VDD2.n61 B 0.02886f
C78 VDD2.n62 B 0.02886f
C79 VDD2.n63 B 0.012928f
C80 VDD2.n64 B 0.01221f
C81 VDD2.n65 B 0.022722f
C82 VDD2.n66 B 0.022722f
C83 VDD2.n67 B 0.01221f
C84 VDD2.n68 B 0.012928f
C85 VDD2.n69 B 0.02886f
C86 VDD2.n70 B 0.02886f
C87 VDD2.n71 B 0.012928f
C88 VDD2.n72 B 0.01221f
C89 VDD2.n73 B 0.022722f
C90 VDD2.n74 B 0.022722f
C91 VDD2.n75 B 0.01221f
C92 VDD2.n76 B 0.01221f
C93 VDD2.n77 B 0.012928f
C94 VDD2.n78 B 0.02886f
C95 VDD2.n79 B 0.02886f
C96 VDD2.n80 B 0.02886f
C97 VDD2.n81 B 0.012569f
C98 VDD2.n82 B 0.01221f
C99 VDD2.n83 B 0.022722f
C100 VDD2.n84 B 0.022722f
C101 VDD2.n85 B 0.01221f
C102 VDD2.n86 B 0.012928f
C103 VDD2.n87 B 0.02886f
C104 VDD2.n88 B 0.02886f
C105 VDD2.n89 B 0.012928f
C106 VDD2.n90 B 0.01221f
C107 VDD2.n91 B 0.022722f
C108 VDD2.n92 B 0.022722f
C109 VDD2.n93 B 0.01221f
C110 VDD2.n94 B 0.012928f
C111 VDD2.n95 B 0.02886f
C112 VDD2.n96 B 0.061663f
C113 VDD2.n97 B 0.012928f
C114 VDD2.n98 B 0.01221f
C115 VDD2.n99 B 0.05159f
C116 VDD2.n100 B 0.051452f
C117 VDD2.t1 B 0.326975f
C118 VDD2.t2 B 0.326975f
C119 VDD2.n101 B 2.98003f
C120 VDD2.n102 B 2.09094f
C121 VDD2.n103 B 0.031478f
C122 VDD2.n104 B 0.022722f
C123 VDD2.n105 B 0.01221f
C124 VDD2.n106 B 0.02886f
C125 VDD2.n107 B 0.012928f
C126 VDD2.n108 B 0.022722f
C127 VDD2.n109 B 0.01221f
C128 VDD2.n110 B 0.02886f
C129 VDD2.n111 B 0.012928f
C130 VDD2.n112 B 0.022722f
C131 VDD2.n113 B 0.012569f
C132 VDD2.n114 B 0.02886f
C133 VDD2.n115 B 0.01221f
C134 VDD2.n116 B 0.012928f
C135 VDD2.n117 B 0.022722f
C136 VDD2.n118 B 0.01221f
C137 VDD2.n119 B 0.02886f
C138 VDD2.n120 B 0.012928f
C139 VDD2.n121 B 0.022722f
C140 VDD2.n122 B 0.01221f
C141 VDD2.n123 B 0.02886f
C142 VDD2.n124 B 0.012928f
C143 VDD2.n125 B 0.022722f
C144 VDD2.n126 B 0.01221f
C145 VDD2.n127 B 0.02886f
C146 VDD2.n128 B 0.012928f
C147 VDD2.n129 B 0.022722f
C148 VDD2.n130 B 0.01221f
C149 VDD2.n131 B 0.02886f
C150 VDD2.n132 B 0.012928f
C151 VDD2.n133 B 0.022722f
C152 VDD2.n134 B 0.01221f
C153 VDD2.n135 B 0.021645f
C154 VDD2.n136 B 0.017048f
C155 VDD2.t4 B 0.047837f
C156 VDD2.n137 B 0.166487f
C157 VDD2.n138 B 1.81262f
C158 VDD2.n139 B 0.01221f
C159 VDD2.n140 B 0.012928f
C160 VDD2.n141 B 0.02886f
C161 VDD2.n142 B 0.02886f
C162 VDD2.n143 B 0.012928f
C163 VDD2.n144 B 0.01221f
C164 VDD2.n145 B 0.022722f
C165 VDD2.n146 B 0.022722f
C166 VDD2.n147 B 0.01221f
C167 VDD2.n148 B 0.012928f
C168 VDD2.n149 B 0.02886f
C169 VDD2.n150 B 0.02886f
C170 VDD2.n151 B 0.012928f
C171 VDD2.n152 B 0.01221f
C172 VDD2.n153 B 0.022722f
C173 VDD2.n154 B 0.022722f
C174 VDD2.n155 B 0.01221f
C175 VDD2.n156 B 0.012928f
C176 VDD2.n157 B 0.02886f
C177 VDD2.n158 B 0.02886f
C178 VDD2.n159 B 0.012928f
C179 VDD2.n160 B 0.01221f
C180 VDD2.n161 B 0.022722f
C181 VDD2.n162 B 0.022722f
C182 VDD2.n163 B 0.01221f
C183 VDD2.n164 B 0.012928f
C184 VDD2.n165 B 0.02886f
C185 VDD2.n166 B 0.02886f
C186 VDD2.n167 B 0.012928f
C187 VDD2.n168 B 0.01221f
C188 VDD2.n169 B 0.022722f
C189 VDD2.n170 B 0.022722f
C190 VDD2.n171 B 0.01221f
C191 VDD2.n172 B 0.012928f
C192 VDD2.n173 B 0.02886f
C193 VDD2.n174 B 0.02886f
C194 VDD2.n175 B 0.012928f
C195 VDD2.n176 B 0.01221f
C196 VDD2.n177 B 0.022722f
C197 VDD2.n178 B 0.022722f
C198 VDD2.n179 B 0.01221f
C199 VDD2.n180 B 0.012928f
C200 VDD2.n181 B 0.02886f
C201 VDD2.n182 B 0.02886f
C202 VDD2.n183 B 0.02886f
C203 VDD2.n184 B 0.012569f
C204 VDD2.n185 B 0.01221f
C205 VDD2.n186 B 0.022722f
C206 VDD2.n187 B 0.022722f
C207 VDD2.n188 B 0.01221f
C208 VDD2.n189 B 0.012928f
C209 VDD2.n190 B 0.02886f
C210 VDD2.n191 B 0.02886f
C211 VDD2.n192 B 0.012928f
C212 VDD2.n193 B 0.01221f
C213 VDD2.n194 B 0.022722f
C214 VDD2.n195 B 0.022722f
C215 VDD2.n196 B 0.01221f
C216 VDD2.n197 B 0.012928f
C217 VDD2.n198 B 0.02886f
C218 VDD2.n199 B 0.061663f
C219 VDD2.n200 B 0.012928f
C220 VDD2.n201 B 0.01221f
C221 VDD2.n202 B 0.05159f
C222 VDD2.n203 B 0.050087f
C223 VDD2.n204 B 2.32626f
C224 VDD2.t0 B 0.326975f
C225 VDD2.t3 B 0.326975f
C226 VDD2.n205 B 2.98f
C227 VN.n0 B 0.188158f
C228 VN.t4 B 1.78915f
C229 VN.t0 B 1.86214f
C230 VN.n1 B 0.695712f
C231 VN.n2 B 0.684157f
C232 VN.n3 B 0.052578f
C233 VN.t3 B 1.84386f
C234 VN.n4 B 0.698109f
C235 VN.n5 B 0.039817f
C236 VN.n6 B 0.188158f
C237 VN.t5 B 1.78915f
C238 VN.t2 B 1.86214f
C239 VN.n7 B 0.695712f
C240 VN.n8 B 0.684157f
C241 VN.n9 B 0.052578f
C242 VN.t1 B 1.84386f
C243 VN.n10 B 0.698109f
C244 VN.n11 B 2.1133f
C245 VDD1.n0 B 0.031503f
C246 VDD1.n1 B 0.02274f
C247 VDD1.n2 B 0.01222f
C248 VDD1.n3 B 0.028883f
C249 VDD1.n4 B 0.012939f
C250 VDD1.n5 B 0.02274f
C251 VDD1.n6 B 0.01222f
C252 VDD1.n7 B 0.028883f
C253 VDD1.n8 B 0.012939f
C254 VDD1.n9 B 0.02274f
C255 VDD1.n10 B 0.012579f
C256 VDD1.n11 B 0.028883f
C257 VDD1.n12 B 0.01222f
C258 VDD1.n13 B 0.012939f
C259 VDD1.n14 B 0.02274f
C260 VDD1.n15 B 0.01222f
C261 VDD1.n16 B 0.028883f
C262 VDD1.n17 B 0.012939f
C263 VDD1.n18 B 0.02274f
C264 VDD1.n19 B 0.01222f
C265 VDD1.n20 B 0.028883f
C266 VDD1.n21 B 0.012939f
C267 VDD1.n22 B 0.02274f
C268 VDD1.n23 B 0.01222f
C269 VDD1.n24 B 0.028883f
C270 VDD1.n25 B 0.012939f
C271 VDD1.n26 B 0.02274f
C272 VDD1.n27 B 0.01222f
C273 VDD1.n28 B 0.028883f
C274 VDD1.n29 B 0.012939f
C275 VDD1.n30 B 0.02274f
C276 VDD1.n31 B 0.01222f
C277 VDD1.n32 B 0.021662f
C278 VDD1.n33 B 0.017062f
C279 VDD1.t4 B 0.047875f
C280 VDD1.n34 B 0.166619f
C281 VDD1.n35 B 1.81406f
C282 VDD1.n36 B 0.01222f
C283 VDD1.n37 B 0.012939f
C284 VDD1.n38 B 0.028883f
C285 VDD1.n39 B 0.028883f
C286 VDD1.n40 B 0.012939f
C287 VDD1.n41 B 0.01222f
C288 VDD1.n42 B 0.02274f
C289 VDD1.n43 B 0.02274f
C290 VDD1.n44 B 0.01222f
C291 VDD1.n45 B 0.012939f
C292 VDD1.n46 B 0.028883f
C293 VDD1.n47 B 0.028883f
C294 VDD1.n48 B 0.012939f
C295 VDD1.n49 B 0.01222f
C296 VDD1.n50 B 0.02274f
C297 VDD1.n51 B 0.02274f
C298 VDD1.n52 B 0.01222f
C299 VDD1.n53 B 0.012939f
C300 VDD1.n54 B 0.028883f
C301 VDD1.n55 B 0.028883f
C302 VDD1.n56 B 0.012939f
C303 VDD1.n57 B 0.01222f
C304 VDD1.n58 B 0.02274f
C305 VDD1.n59 B 0.02274f
C306 VDD1.n60 B 0.01222f
C307 VDD1.n61 B 0.012939f
C308 VDD1.n62 B 0.028883f
C309 VDD1.n63 B 0.028883f
C310 VDD1.n64 B 0.012939f
C311 VDD1.n65 B 0.01222f
C312 VDD1.n66 B 0.02274f
C313 VDD1.n67 B 0.02274f
C314 VDD1.n68 B 0.01222f
C315 VDD1.n69 B 0.012939f
C316 VDD1.n70 B 0.028883f
C317 VDD1.n71 B 0.028883f
C318 VDD1.n72 B 0.012939f
C319 VDD1.n73 B 0.01222f
C320 VDD1.n74 B 0.02274f
C321 VDD1.n75 B 0.02274f
C322 VDD1.n76 B 0.01222f
C323 VDD1.n77 B 0.012939f
C324 VDD1.n78 B 0.028883f
C325 VDD1.n79 B 0.028883f
C326 VDD1.n80 B 0.028883f
C327 VDD1.n81 B 0.012579f
C328 VDD1.n82 B 0.01222f
C329 VDD1.n83 B 0.02274f
C330 VDD1.n84 B 0.02274f
C331 VDD1.n85 B 0.01222f
C332 VDD1.n86 B 0.012939f
C333 VDD1.n87 B 0.028883f
C334 VDD1.n88 B 0.028883f
C335 VDD1.n89 B 0.012939f
C336 VDD1.n90 B 0.01222f
C337 VDD1.n91 B 0.02274f
C338 VDD1.n92 B 0.02274f
C339 VDD1.n93 B 0.01222f
C340 VDD1.n94 B 0.012939f
C341 VDD1.n95 B 0.028883f
C342 VDD1.n96 B 0.061713f
C343 VDD1.n97 B 0.012939f
C344 VDD1.n98 B 0.01222f
C345 VDD1.n99 B 0.051631f
C346 VDD1.n100 B 0.051835f
C347 VDD1.n101 B 0.031503f
C348 VDD1.n102 B 0.02274f
C349 VDD1.n103 B 0.01222f
C350 VDD1.n104 B 0.028883f
C351 VDD1.n105 B 0.012939f
C352 VDD1.n106 B 0.02274f
C353 VDD1.n107 B 0.01222f
C354 VDD1.n108 B 0.028883f
C355 VDD1.n109 B 0.012939f
C356 VDD1.n110 B 0.02274f
C357 VDD1.n111 B 0.012579f
C358 VDD1.n112 B 0.028883f
C359 VDD1.n113 B 0.012939f
C360 VDD1.n114 B 0.02274f
C361 VDD1.n115 B 0.01222f
C362 VDD1.n116 B 0.028883f
C363 VDD1.n117 B 0.012939f
C364 VDD1.n118 B 0.02274f
C365 VDD1.n119 B 0.01222f
C366 VDD1.n120 B 0.028883f
C367 VDD1.n121 B 0.012939f
C368 VDD1.n122 B 0.02274f
C369 VDD1.n123 B 0.01222f
C370 VDD1.n124 B 0.028883f
C371 VDD1.n125 B 0.012939f
C372 VDD1.n126 B 0.02274f
C373 VDD1.n127 B 0.01222f
C374 VDD1.n128 B 0.028883f
C375 VDD1.n129 B 0.012939f
C376 VDD1.n130 B 0.02274f
C377 VDD1.n131 B 0.01222f
C378 VDD1.n132 B 0.021662f
C379 VDD1.n133 B 0.017062f
C380 VDD1.t2 B 0.047875f
C381 VDD1.n134 B 0.166619f
C382 VDD1.n135 B 1.81406f
C383 VDD1.n136 B 0.01222f
C384 VDD1.n137 B 0.012939f
C385 VDD1.n138 B 0.028883f
C386 VDD1.n139 B 0.028883f
C387 VDD1.n140 B 0.012939f
C388 VDD1.n141 B 0.01222f
C389 VDD1.n142 B 0.02274f
C390 VDD1.n143 B 0.02274f
C391 VDD1.n144 B 0.01222f
C392 VDD1.n145 B 0.012939f
C393 VDD1.n146 B 0.028883f
C394 VDD1.n147 B 0.028883f
C395 VDD1.n148 B 0.012939f
C396 VDD1.n149 B 0.01222f
C397 VDD1.n150 B 0.02274f
C398 VDD1.n151 B 0.02274f
C399 VDD1.n152 B 0.01222f
C400 VDD1.n153 B 0.012939f
C401 VDD1.n154 B 0.028883f
C402 VDD1.n155 B 0.028883f
C403 VDD1.n156 B 0.012939f
C404 VDD1.n157 B 0.01222f
C405 VDD1.n158 B 0.02274f
C406 VDD1.n159 B 0.02274f
C407 VDD1.n160 B 0.01222f
C408 VDD1.n161 B 0.012939f
C409 VDD1.n162 B 0.028883f
C410 VDD1.n163 B 0.028883f
C411 VDD1.n164 B 0.012939f
C412 VDD1.n165 B 0.01222f
C413 VDD1.n166 B 0.02274f
C414 VDD1.n167 B 0.02274f
C415 VDD1.n168 B 0.01222f
C416 VDD1.n169 B 0.012939f
C417 VDD1.n170 B 0.028883f
C418 VDD1.n171 B 0.028883f
C419 VDD1.n172 B 0.012939f
C420 VDD1.n173 B 0.01222f
C421 VDD1.n174 B 0.02274f
C422 VDD1.n175 B 0.02274f
C423 VDD1.n176 B 0.01222f
C424 VDD1.n177 B 0.01222f
C425 VDD1.n178 B 0.012939f
C426 VDD1.n179 B 0.028883f
C427 VDD1.n180 B 0.028883f
C428 VDD1.n181 B 0.028883f
C429 VDD1.n182 B 0.012579f
C430 VDD1.n183 B 0.01222f
C431 VDD1.n184 B 0.02274f
C432 VDD1.n185 B 0.02274f
C433 VDD1.n186 B 0.01222f
C434 VDD1.n187 B 0.012939f
C435 VDD1.n188 B 0.028883f
C436 VDD1.n189 B 0.028883f
C437 VDD1.n190 B 0.012939f
C438 VDD1.n191 B 0.01222f
C439 VDD1.n192 B 0.02274f
C440 VDD1.n193 B 0.02274f
C441 VDD1.n194 B 0.01222f
C442 VDD1.n195 B 0.012939f
C443 VDD1.n196 B 0.028883f
C444 VDD1.n197 B 0.061713f
C445 VDD1.n198 B 0.012939f
C446 VDD1.n199 B 0.01222f
C447 VDD1.n200 B 0.051631f
C448 VDD1.n201 B 0.051492f
C449 VDD1.t3 B 0.327235f
C450 VDD1.t1 B 0.327235f
C451 VDD1.n202 B 2.9824f
C452 VDD1.n203 B 2.1674f
C453 VDD1.t0 B 0.327235f
C454 VDD1.t5 B 0.327235f
C455 VDD1.n204 B 2.98145f
C456 VDD1.n205 B 2.52174f
C457 VTAIL.t5 B 0.333446f
C458 VTAIL.t3 B 0.333446f
C459 VTAIL.n0 B 2.96527f
C460 VTAIL.n1 B 0.330893f
C461 VTAIL.n2 B 0.032101f
C462 VTAIL.n3 B 0.023172f
C463 VTAIL.n4 B 0.012452f
C464 VTAIL.n5 B 0.029431f
C465 VTAIL.n6 B 0.013184f
C466 VTAIL.n7 B 0.023172f
C467 VTAIL.n8 B 0.012452f
C468 VTAIL.n9 B 0.029431f
C469 VTAIL.n10 B 0.013184f
C470 VTAIL.n11 B 0.023172f
C471 VTAIL.n12 B 0.012818f
C472 VTAIL.n13 B 0.029431f
C473 VTAIL.n14 B 0.013184f
C474 VTAIL.n15 B 0.023172f
C475 VTAIL.n16 B 0.012452f
C476 VTAIL.n17 B 0.029431f
C477 VTAIL.n18 B 0.013184f
C478 VTAIL.n19 B 0.023172f
C479 VTAIL.n20 B 0.012452f
C480 VTAIL.n21 B 0.029431f
C481 VTAIL.n22 B 0.013184f
C482 VTAIL.n23 B 0.023172f
C483 VTAIL.n24 B 0.012452f
C484 VTAIL.n25 B 0.029431f
C485 VTAIL.n26 B 0.013184f
C486 VTAIL.n27 B 0.023172f
C487 VTAIL.n28 B 0.012452f
C488 VTAIL.n29 B 0.029431f
C489 VTAIL.n30 B 0.013184f
C490 VTAIL.n31 B 0.023172f
C491 VTAIL.n32 B 0.012452f
C492 VTAIL.n33 B 0.022073f
C493 VTAIL.n34 B 0.017386f
C494 VTAIL.t6 B 0.048783f
C495 VTAIL.n35 B 0.169782f
C496 VTAIL.n36 B 1.84849f
C497 VTAIL.n37 B 0.012452f
C498 VTAIL.n38 B 0.013184f
C499 VTAIL.n39 B 0.029431f
C500 VTAIL.n40 B 0.029431f
C501 VTAIL.n41 B 0.013184f
C502 VTAIL.n42 B 0.012452f
C503 VTAIL.n43 B 0.023172f
C504 VTAIL.n44 B 0.023172f
C505 VTAIL.n45 B 0.012452f
C506 VTAIL.n46 B 0.013184f
C507 VTAIL.n47 B 0.029431f
C508 VTAIL.n48 B 0.029431f
C509 VTAIL.n49 B 0.013184f
C510 VTAIL.n50 B 0.012452f
C511 VTAIL.n51 B 0.023172f
C512 VTAIL.n52 B 0.023172f
C513 VTAIL.n53 B 0.012452f
C514 VTAIL.n54 B 0.013184f
C515 VTAIL.n55 B 0.029431f
C516 VTAIL.n56 B 0.029431f
C517 VTAIL.n57 B 0.013184f
C518 VTAIL.n58 B 0.012452f
C519 VTAIL.n59 B 0.023172f
C520 VTAIL.n60 B 0.023172f
C521 VTAIL.n61 B 0.012452f
C522 VTAIL.n62 B 0.013184f
C523 VTAIL.n63 B 0.029431f
C524 VTAIL.n64 B 0.029431f
C525 VTAIL.n65 B 0.013184f
C526 VTAIL.n66 B 0.012452f
C527 VTAIL.n67 B 0.023172f
C528 VTAIL.n68 B 0.023172f
C529 VTAIL.n69 B 0.012452f
C530 VTAIL.n70 B 0.013184f
C531 VTAIL.n71 B 0.029431f
C532 VTAIL.n72 B 0.029431f
C533 VTAIL.n73 B 0.013184f
C534 VTAIL.n74 B 0.012452f
C535 VTAIL.n75 B 0.023172f
C536 VTAIL.n76 B 0.023172f
C537 VTAIL.n77 B 0.012452f
C538 VTAIL.n78 B 0.012452f
C539 VTAIL.n79 B 0.013184f
C540 VTAIL.n80 B 0.029431f
C541 VTAIL.n81 B 0.029431f
C542 VTAIL.n82 B 0.029431f
C543 VTAIL.n83 B 0.012818f
C544 VTAIL.n84 B 0.012452f
C545 VTAIL.n85 B 0.023172f
C546 VTAIL.n86 B 0.023172f
C547 VTAIL.n87 B 0.012452f
C548 VTAIL.n88 B 0.013184f
C549 VTAIL.n89 B 0.029431f
C550 VTAIL.n90 B 0.029431f
C551 VTAIL.n91 B 0.013184f
C552 VTAIL.n92 B 0.012452f
C553 VTAIL.n93 B 0.023172f
C554 VTAIL.n94 B 0.023172f
C555 VTAIL.n95 B 0.012452f
C556 VTAIL.n96 B 0.013184f
C557 VTAIL.n97 B 0.029431f
C558 VTAIL.n98 B 0.062884f
C559 VTAIL.n99 B 0.013184f
C560 VTAIL.n100 B 0.012452f
C561 VTAIL.n101 B 0.052611f
C562 VTAIL.n102 B 0.035071f
C563 VTAIL.n103 B 0.167298f
C564 VTAIL.t7 B 0.333446f
C565 VTAIL.t8 B 0.333446f
C566 VTAIL.n104 B 2.96527f
C567 VTAIL.n105 B 1.94779f
C568 VTAIL.t4 B 0.333446f
C569 VTAIL.t0 B 0.333446f
C570 VTAIL.n106 B 2.96529f
C571 VTAIL.n107 B 1.94778f
C572 VTAIL.n108 B 0.032101f
C573 VTAIL.n109 B 0.023172f
C574 VTAIL.n110 B 0.012452f
C575 VTAIL.n111 B 0.029431f
C576 VTAIL.n112 B 0.013184f
C577 VTAIL.n113 B 0.023172f
C578 VTAIL.n114 B 0.012452f
C579 VTAIL.n115 B 0.029431f
C580 VTAIL.n116 B 0.013184f
C581 VTAIL.n117 B 0.023172f
C582 VTAIL.n118 B 0.012818f
C583 VTAIL.n119 B 0.029431f
C584 VTAIL.n120 B 0.012452f
C585 VTAIL.n121 B 0.013184f
C586 VTAIL.n122 B 0.023172f
C587 VTAIL.n123 B 0.012452f
C588 VTAIL.n124 B 0.029431f
C589 VTAIL.n125 B 0.013184f
C590 VTAIL.n126 B 0.023172f
C591 VTAIL.n127 B 0.012452f
C592 VTAIL.n128 B 0.029431f
C593 VTAIL.n129 B 0.013184f
C594 VTAIL.n130 B 0.023172f
C595 VTAIL.n131 B 0.012452f
C596 VTAIL.n132 B 0.029431f
C597 VTAIL.n133 B 0.013184f
C598 VTAIL.n134 B 0.023172f
C599 VTAIL.n135 B 0.012452f
C600 VTAIL.n136 B 0.029431f
C601 VTAIL.n137 B 0.013184f
C602 VTAIL.n138 B 0.023172f
C603 VTAIL.n139 B 0.012452f
C604 VTAIL.n140 B 0.022073f
C605 VTAIL.n141 B 0.017386f
C606 VTAIL.t1 B 0.048783f
C607 VTAIL.n142 B 0.169782f
C608 VTAIL.n143 B 1.84849f
C609 VTAIL.n144 B 0.012452f
C610 VTAIL.n145 B 0.013184f
C611 VTAIL.n146 B 0.029431f
C612 VTAIL.n147 B 0.029431f
C613 VTAIL.n148 B 0.013184f
C614 VTAIL.n149 B 0.012452f
C615 VTAIL.n150 B 0.023172f
C616 VTAIL.n151 B 0.023172f
C617 VTAIL.n152 B 0.012452f
C618 VTAIL.n153 B 0.013184f
C619 VTAIL.n154 B 0.029431f
C620 VTAIL.n155 B 0.029431f
C621 VTAIL.n156 B 0.013184f
C622 VTAIL.n157 B 0.012452f
C623 VTAIL.n158 B 0.023172f
C624 VTAIL.n159 B 0.023172f
C625 VTAIL.n160 B 0.012452f
C626 VTAIL.n161 B 0.013184f
C627 VTAIL.n162 B 0.029431f
C628 VTAIL.n163 B 0.029431f
C629 VTAIL.n164 B 0.013184f
C630 VTAIL.n165 B 0.012452f
C631 VTAIL.n166 B 0.023172f
C632 VTAIL.n167 B 0.023172f
C633 VTAIL.n168 B 0.012452f
C634 VTAIL.n169 B 0.013184f
C635 VTAIL.n170 B 0.029431f
C636 VTAIL.n171 B 0.029431f
C637 VTAIL.n172 B 0.013184f
C638 VTAIL.n173 B 0.012452f
C639 VTAIL.n174 B 0.023172f
C640 VTAIL.n175 B 0.023172f
C641 VTAIL.n176 B 0.012452f
C642 VTAIL.n177 B 0.013184f
C643 VTAIL.n178 B 0.029431f
C644 VTAIL.n179 B 0.029431f
C645 VTAIL.n180 B 0.013184f
C646 VTAIL.n181 B 0.012452f
C647 VTAIL.n182 B 0.023172f
C648 VTAIL.n183 B 0.023172f
C649 VTAIL.n184 B 0.012452f
C650 VTAIL.n185 B 0.013184f
C651 VTAIL.n186 B 0.029431f
C652 VTAIL.n187 B 0.029431f
C653 VTAIL.n188 B 0.029431f
C654 VTAIL.n189 B 0.012818f
C655 VTAIL.n190 B 0.012452f
C656 VTAIL.n191 B 0.023172f
C657 VTAIL.n192 B 0.023172f
C658 VTAIL.n193 B 0.012452f
C659 VTAIL.n194 B 0.013184f
C660 VTAIL.n195 B 0.029431f
C661 VTAIL.n196 B 0.029431f
C662 VTAIL.n197 B 0.013184f
C663 VTAIL.n198 B 0.012452f
C664 VTAIL.n199 B 0.023172f
C665 VTAIL.n200 B 0.023172f
C666 VTAIL.n201 B 0.012452f
C667 VTAIL.n202 B 0.013184f
C668 VTAIL.n203 B 0.029431f
C669 VTAIL.n204 B 0.062884f
C670 VTAIL.n205 B 0.013184f
C671 VTAIL.n206 B 0.012452f
C672 VTAIL.n207 B 0.052611f
C673 VTAIL.n208 B 0.035071f
C674 VTAIL.n209 B 0.167298f
C675 VTAIL.t11 B 0.333446f
C676 VTAIL.t9 B 0.333446f
C677 VTAIL.n210 B 2.96529f
C678 VTAIL.n211 B 0.383016f
C679 VTAIL.n212 B 0.032101f
C680 VTAIL.n213 B 0.023172f
C681 VTAIL.n214 B 0.012452f
C682 VTAIL.n215 B 0.029431f
C683 VTAIL.n216 B 0.013184f
C684 VTAIL.n217 B 0.023172f
C685 VTAIL.n218 B 0.012452f
C686 VTAIL.n219 B 0.029431f
C687 VTAIL.n220 B 0.013184f
C688 VTAIL.n221 B 0.023172f
C689 VTAIL.n222 B 0.012818f
C690 VTAIL.n223 B 0.029431f
C691 VTAIL.n224 B 0.012452f
C692 VTAIL.n225 B 0.013184f
C693 VTAIL.n226 B 0.023172f
C694 VTAIL.n227 B 0.012452f
C695 VTAIL.n228 B 0.029431f
C696 VTAIL.n229 B 0.013184f
C697 VTAIL.n230 B 0.023172f
C698 VTAIL.n231 B 0.012452f
C699 VTAIL.n232 B 0.029431f
C700 VTAIL.n233 B 0.013184f
C701 VTAIL.n234 B 0.023172f
C702 VTAIL.n235 B 0.012452f
C703 VTAIL.n236 B 0.029431f
C704 VTAIL.n237 B 0.013184f
C705 VTAIL.n238 B 0.023172f
C706 VTAIL.n239 B 0.012452f
C707 VTAIL.n240 B 0.029431f
C708 VTAIL.n241 B 0.013184f
C709 VTAIL.n242 B 0.023172f
C710 VTAIL.n243 B 0.012452f
C711 VTAIL.n244 B 0.022073f
C712 VTAIL.n245 B 0.017386f
C713 VTAIL.t10 B 0.048783f
C714 VTAIL.n246 B 0.169782f
C715 VTAIL.n247 B 1.84849f
C716 VTAIL.n248 B 0.012452f
C717 VTAIL.n249 B 0.013184f
C718 VTAIL.n250 B 0.029431f
C719 VTAIL.n251 B 0.029431f
C720 VTAIL.n252 B 0.013184f
C721 VTAIL.n253 B 0.012452f
C722 VTAIL.n254 B 0.023172f
C723 VTAIL.n255 B 0.023172f
C724 VTAIL.n256 B 0.012452f
C725 VTAIL.n257 B 0.013184f
C726 VTAIL.n258 B 0.029431f
C727 VTAIL.n259 B 0.029431f
C728 VTAIL.n260 B 0.013184f
C729 VTAIL.n261 B 0.012452f
C730 VTAIL.n262 B 0.023172f
C731 VTAIL.n263 B 0.023172f
C732 VTAIL.n264 B 0.012452f
C733 VTAIL.n265 B 0.013184f
C734 VTAIL.n266 B 0.029431f
C735 VTAIL.n267 B 0.029431f
C736 VTAIL.n268 B 0.013184f
C737 VTAIL.n269 B 0.012452f
C738 VTAIL.n270 B 0.023172f
C739 VTAIL.n271 B 0.023172f
C740 VTAIL.n272 B 0.012452f
C741 VTAIL.n273 B 0.013184f
C742 VTAIL.n274 B 0.029431f
C743 VTAIL.n275 B 0.029431f
C744 VTAIL.n276 B 0.013184f
C745 VTAIL.n277 B 0.012452f
C746 VTAIL.n278 B 0.023172f
C747 VTAIL.n279 B 0.023172f
C748 VTAIL.n280 B 0.012452f
C749 VTAIL.n281 B 0.013184f
C750 VTAIL.n282 B 0.029431f
C751 VTAIL.n283 B 0.029431f
C752 VTAIL.n284 B 0.013184f
C753 VTAIL.n285 B 0.012452f
C754 VTAIL.n286 B 0.023172f
C755 VTAIL.n287 B 0.023172f
C756 VTAIL.n288 B 0.012452f
C757 VTAIL.n289 B 0.013184f
C758 VTAIL.n290 B 0.029431f
C759 VTAIL.n291 B 0.029431f
C760 VTAIL.n292 B 0.029431f
C761 VTAIL.n293 B 0.012818f
C762 VTAIL.n294 B 0.012452f
C763 VTAIL.n295 B 0.023172f
C764 VTAIL.n296 B 0.023172f
C765 VTAIL.n297 B 0.012452f
C766 VTAIL.n298 B 0.013184f
C767 VTAIL.n299 B 0.029431f
C768 VTAIL.n300 B 0.029431f
C769 VTAIL.n301 B 0.013184f
C770 VTAIL.n302 B 0.012452f
C771 VTAIL.n303 B 0.023172f
C772 VTAIL.n304 B 0.023172f
C773 VTAIL.n305 B 0.012452f
C774 VTAIL.n306 B 0.013184f
C775 VTAIL.n307 B 0.029431f
C776 VTAIL.n308 B 0.062884f
C777 VTAIL.n309 B 0.013184f
C778 VTAIL.n310 B 0.012452f
C779 VTAIL.n311 B 0.052611f
C780 VTAIL.n312 B 0.035071f
C781 VTAIL.n313 B 1.65675f
C782 VTAIL.n314 B 0.032101f
C783 VTAIL.n315 B 0.023172f
C784 VTAIL.n316 B 0.012452f
C785 VTAIL.n317 B 0.029431f
C786 VTAIL.n318 B 0.013184f
C787 VTAIL.n319 B 0.023172f
C788 VTAIL.n320 B 0.012452f
C789 VTAIL.n321 B 0.029431f
C790 VTAIL.n322 B 0.013184f
C791 VTAIL.n323 B 0.023172f
C792 VTAIL.n324 B 0.012818f
C793 VTAIL.n325 B 0.029431f
C794 VTAIL.n326 B 0.013184f
C795 VTAIL.n327 B 0.023172f
C796 VTAIL.n328 B 0.012452f
C797 VTAIL.n329 B 0.029431f
C798 VTAIL.n330 B 0.013184f
C799 VTAIL.n331 B 0.023172f
C800 VTAIL.n332 B 0.012452f
C801 VTAIL.n333 B 0.029431f
C802 VTAIL.n334 B 0.013184f
C803 VTAIL.n335 B 0.023172f
C804 VTAIL.n336 B 0.012452f
C805 VTAIL.n337 B 0.029431f
C806 VTAIL.n338 B 0.013184f
C807 VTAIL.n339 B 0.023172f
C808 VTAIL.n340 B 0.012452f
C809 VTAIL.n341 B 0.029431f
C810 VTAIL.n342 B 0.013184f
C811 VTAIL.n343 B 0.023172f
C812 VTAIL.n344 B 0.012452f
C813 VTAIL.n345 B 0.022073f
C814 VTAIL.n346 B 0.017386f
C815 VTAIL.t2 B 0.048783f
C816 VTAIL.n347 B 0.169782f
C817 VTAIL.n348 B 1.84849f
C818 VTAIL.n349 B 0.012452f
C819 VTAIL.n350 B 0.013184f
C820 VTAIL.n351 B 0.029431f
C821 VTAIL.n352 B 0.029431f
C822 VTAIL.n353 B 0.013184f
C823 VTAIL.n354 B 0.012452f
C824 VTAIL.n355 B 0.023172f
C825 VTAIL.n356 B 0.023172f
C826 VTAIL.n357 B 0.012452f
C827 VTAIL.n358 B 0.013184f
C828 VTAIL.n359 B 0.029431f
C829 VTAIL.n360 B 0.029431f
C830 VTAIL.n361 B 0.013184f
C831 VTAIL.n362 B 0.012452f
C832 VTAIL.n363 B 0.023172f
C833 VTAIL.n364 B 0.023172f
C834 VTAIL.n365 B 0.012452f
C835 VTAIL.n366 B 0.013184f
C836 VTAIL.n367 B 0.029431f
C837 VTAIL.n368 B 0.029431f
C838 VTAIL.n369 B 0.013184f
C839 VTAIL.n370 B 0.012452f
C840 VTAIL.n371 B 0.023172f
C841 VTAIL.n372 B 0.023172f
C842 VTAIL.n373 B 0.012452f
C843 VTAIL.n374 B 0.013184f
C844 VTAIL.n375 B 0.029431f
C845 VTAIL.n376 B 0.029431f
C846 VTAIL.n377 B 0.013184f
C847 VTAIL.n378 B 0.012452f
C848 VTAIL.n379 B 0.023172f
C849 VTAIL.n380 B 0.023172f
C850 VTAIL.n381 B 0.012452f
C851 VTAIL.n382 B 0.013184f
C852 VTAIL.n383 B 0.029431f
C853 VTAIL.n384 B 0.029431f
C854 VTAIL.n385 B 0.013184f
C855 VTAIL.n386 B 0.012452f
C856 VTAIL.n387 B 0.023172f
C857 VTAIL.n388 B 0.023172f
C858 VTAIL.n389 B 0.012452f
C859 VTAIL.n390 B 0.012452f
C860 VTAIL.n391 B 0.013184f
C861 VTAIL.n392 B 0.029431f
C862 VTAIL.n393 B 0.029431f
C863 VTAIL.n394 B 0.029431f
C864 VTAIL.n395 B 0.012818f
C865 VTAIL.n396 B 0.012452f
C866 VTAIL.n397 B 0.023172f
C867 VTAIL.n398 B 0.023172f
C868 VTAIL.n399 B 0.012452f
C869 VTAIL.n400 B 0.013184f
C870 VTAIL.n401 B 0.029431f
C871 VTAIL.n402 B 0.029431f
C872 VTAIL.n403 B 0.013184f
C873 VTAIL.n404 B 0.012452f
C874 VTAIL.n405 B 0.023172f
C875 VTAIL.n406 B 0.023172f
C876 VTAIL.n407 B 0.012452f
C877 VTAIL.n408 B 0.013184f
C878 VTAIL.n409 B 0.029431f
C879 VTAIL.n410 B 0.062884f
C880 VTAIL.n411 B 0.013184f
C881 VTAIL.n412 B 0.012452f
C882 VTAIL.n413 B 0.052611f
C883 VTAIL.n414 B 0.035071f
C884 VTAIL.n415 B 1.63358f
C885 VP.n0 B 0.057188f
C886 VP.t2 B 1.80356f
C887 VP.t3 B 1.85871f
C888 VP.n1 B 0.703731f
C889 VP.n2 B 0.189673f
C890 VP.t0 B 1.85871f
C891 VP.t5 B 1.80356f
C892 VP.t1 B 1.87713f
C893 VP.n3 B 0.701314f
C894 VP.n4 B 0.689666f
C895 VP.n5 B 0.053001f
C896 VP.n6 B 0.703731f
C897 VP.n7 B 2.10668f
C898 VP.n8 B 2.13975f
C899 VP.n9 B 0.057188f
C900 VP.n10 B 0.053001f
C901 VP.n11 B 0.65183f
C902 VP.n12 B 0.053001f
C903 VP.t4 B 1.85871f
C904 VP.n13 B 0.703731f
C905 VP.n14 B 0.040137f
.ends

