* NGSPICE file created from diff_pair_sample_0063.ext - technology: sky130A

.subckt diff_pair_sample_0063 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=6.3024 pd=33.1 as=0 ps=0 w=16.16 l=1.94
X1 VDD1.t9 VP.t0 VTAIL.t18 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=6.3024 pd=33.1 as=2.6664 ps=16.49 w=16.16 l=1.94
X2 B.t8 B.t6 B.t7 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=6.3024 pd=33.1 as=0 ps=0 w=16.16 l=1.94
X3 VDD1.t8 VP.t1 VTAIL.t17 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=2.6664 pd=16.49 as=2.6664 ps=16.49 w=16.16 l=1.94
X4 VDD1.t7 VP.t2 VTAIL.t12 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=2.6664 pd=16.49 as=6.3024 ps=33.1 w=16.16 l=1.94
X5 VDD2.t9 VN.t0 VTAIL.t3 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=2.6664 pd=16.49 as=2.6664 ps=16.49 w=16.16 l=1.94
X6 VTAIL.t9 VP.t3 VDD1.t6 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=2.6664 pd=16.49 as=2.6664 ps=16.49 w=16.16 l=1.94
X7 VTAIL.t6 VN.t1 VDD2.t8 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=2.6664 pd=16.49 as=2.6664 ps=16.49 w=16.16 l=1.94
X8 VDD2.t7 VN.t2 VTAIL.t7 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=2.6664 pd=16.49 as=2.6664 ps=16.49 w=16.16 l=1.94
X9 VDD2.t6 VN.t3 VTAIL.t0 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=2.6664 pd=16.49 as=6.3024 ps=33.1 w=16.16 l=1.94
X10 VDD1.t5 VP.t4 VTAIL.t13 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=2.6664 pd=16.49 as=2.6664 ps=16.49 w=16.16 l=1.94
X11 VTAIL.t4 VN.t4 VDD2.t5 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=2.6664 pd=16.49 as=2.6664 ps=16.49 w=16.16 l=1.94
X12 VTAIL.t10 VP.t5 VDD1.t4 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=2.6664 pd=16.49 as=2.6664 ps=16.49 w=16.16 l=1.94
X13 VTAIL.t1 VN.t5 VDD2.t4 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=2.6664 pd=16.49 as=2.6664 ps=16.49 w=16.16 l=1.94
X14 B.t5 B.t3 B.t4 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=6.3024 pd=33.1 as=0 ps=0 w=16.16 l=1.94
X15 VDD2.t3 VN.t6 VTAIL.t8 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=2.6664 pd=16.49 as=6.3024 ps=33.1 w=16.16 l=1.94
X16 VTAIL.t5 VN.t7 VDD2.t2 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=2.6664 pd=16.49 as=2.6664 ps=16.49 w=16.16 l=1.94
X17 VDD1.t3 VP.t6 VTAIL.t11 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=2.6664 pd=16.49 as=6.3024 ps=33.1 w=16.16 l=1.94
X18 VDD2.t1 VN.t8 VTAIL.t19 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=6.3024 pd=33.1 as=2.6664 ps=16.49 w=16.16 l=1.94
X19 VTAIL.t15 VP.t7 VDD1.t2 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=2.6664 pd=16.49 as=2.6664 ps=16.49 w=16.16 l=1.94
X20 B.t2 B.t0 B.t1 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=6.3024 pd=33.1 as=0 ps=0 w=16.16 l=1.94
X21 VDD1.t1 VP.t8 VTAIL.t14 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=6.3024 pd=33.1 as=2.6664 ps=16.49 w=16.16 l=1.94
X22 VDD2.t0 VN.t9 VTAIL.t2 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=6.3024 pd=33.1 as=2.6664 ps=16.49 w=16.16 l=1.94
X23 VTAIL.t16 VP.t9 VDD1.t0 w_n3694_n4200# sky130_fd_pr__pfet_01v8 ad=2.6664 pd=16.49 as=2.6664 ps=16.49 w=16.16 l=1.94
R0 B.n617 B.n88 585
R1 B.n619 B.n618 585
R2 B.n620 B.n87 585
R3 B.n622 B.n621 585
R4 B.n623 B.n86 585
R5 B.n625 B.n624 585
R6 B.n626 B.n85 585
R7 B.n628 B.n627 585
R8 B.n629 B.n84 585
R9 B.n631 B.n630 585
R10 B.n632 B.n83 585
R11 B.n634 B.n633 585
R12 B.n635 B.n82 585
R13 B.n637 B.n636 585
R14 B.n638 B.n81 585
R15 B.n640 B.n639 585
R16 B.n641 B.n80 585
R17 B.n643 B.n642 585
R18 B.n644 B.n79 585
R19 B.n646 B.n645 585
R20 B.n647 B.n78 585
R21 B.n649 B.n648 585
R22 B.n650 B.n77 585
R23 B.n652 B.n651 585
R24 B.n653 B.n76 585
R25 B.n655 B.n654 585
R26 B.n656 B.n75 585
R27 B.n658 B.n657 585
R28 B.n659 B.n74 585
R29 B.n661 B.n660 585
R30 B.n662 B.n73 585
R31 B.n664 B.n663 585
R32 B.n665 B.n72 585
R33 B.n667 B.n666 585
R34 B.n668 B.n71 585
R35 B.n670 B.n669 585
R36 B.n671 B.n70 585
R37 B.n673 B.n672 585
R38 B.n674 B.n69 585
R39 B.n676 B.n675 585
R40 B.n677 B.n68 585
R41 B.n679 B.n678 585
R42 B.n680 B.n67 585
R43 B.n682 B.n681 585
R44 B.n683 B.n66 585
R45 B.n685 B.n684 585
R46 B.n686 B.n65 585
R47 B.n688 B.n687 585
R48 B.n689 B.n64 585
R49 B.n691 B.n690 585
R50 B.n692 B.n63 585
R51 B.n694 B.n693 585
R52 B.n695 B.n62 585
R53 B.n697 B.n696 585
R54 B.n699 B.n59 585
R55 B.n701 B.n700 585
R56 B.n702 B.n58 585
R57 B.n704 B.n703 585
R58 B.n705 B.n57 585
R59 B.n707 B.n706 585
R60 B.n708 B.n56 585
R61 B.n710 B.n709 585
R62 B.n711 B.n53 585
R63 B.n714 B.n713 585
R64 B.n715 B.n52 585
R65 B.n717 B.n716 585
R66 B.n718 B.n51 585
R67 B.n720 B.n719 585
R68 B.n721 B.n50 585
R69 B.n723 B.n722 585
R70 B.n724 B.n49 585
R71 B.n726 B.n725 585
R72 B.n727 B.n48 585
R73 B.n729 B.n728 585
R74 B.n730 B.n47 585
R75 B.n732 B.n731 585
R76 B.n733 B.n46 585
R77 B.n735 B.n734 585
R78 B.n736 B.n45 585
R79 B.n738 B.n737 585
R80 B.n739 B.n44 585
R81 B.n741 B.n740 585
R82 B.n742 B.n43 585
R83 B.n744 B.n743 585
R84 B.n745 B.n42 585
R85 B.n747 B.n746 585
R86 B.n748 B.n41 585
R87 B.n750 B.n749 585
R88 B.n751 B.n40 585
R89 B.n753 B.n752 585
R90 B.n754 B.n39 585
R91 B.n756 B.n755 585
R92 B.n757 B.n38 585
R93 B.n759 B.n758 585
R94 B.n760 B.n37 585
R95 B.n762 B.n761 585
R96 B.n763 B.n36 585
R97 B.n765 B.n764 585
R98 B.n766 B.n35 585
R99 B.n768 B.n767 585
R100 B.n769 B.n34 585
R101 B.n771 B.n770 585
R102 B.n772 B.n33 585
R103 B.n774 B.n773 585
R104 B.n775 B.n32 585
R105 B.n777 B.n776 585
R106 B.n778 B.n31 585
R107 B.n780 B.n779 585
R108 B.n781 B.n30 585
R109 B.n783 B.n782 585
R110 B.n784 B.n29 585
R111 B.n786 B.n785 585
R112 B.n787 B.n28 585
R113 B.n789 B.n788 585
R114 B.n790 B.n27 585
R115 B.n792 B.n791 585
R116 B.n793 B.n26 585
R117 B.n616 B.n615 585
R118 B.n614 B.n89 585
R119 B.n613 B.n612 585
R120 B.n611 B.n90 585
R121 B.n610 B.n609 585
R122 B.n608 B.n91 585
R123 B.n607 B.n606 585
R124 B.n605 B.n92 585
R125 B.n604 B.n603 585
R126 B.n602 B.n93 585
R127 B.n601 B.n600 585
R128 B.n599 B.n94 585
R129 B.n598 B.n597 585
R130 B.n596 B.n95 585
R131 B.n595 B.n594 585
R132 B.n593 B.n96 585
R133 B.n592 B.n591 585
R134 B.n590 B.n97 585
R135 B.n589 B.n588 585
R136 B.n587 B.n98 585
R137 B.n586 B.n585 585
R138 B.n584 B.n99 585
R139 B.n583 B.n582 585
R140 B.n581 B.n100 585
R141 B.n580 B.n579 585
R142 B.n578 B.n101 585
R143 B.n577 B.n576 585
R144 B.n575 B.n102 585
R145 B.n574 B.n573 585
R146 B.n572 B.n103 585
R147 B.n571 B.n570 585
R148 B.n569 B.n104 585
R149 B.n568 B.n567 585
R150 B.n566 B.n105 585
R151 B.n565 B.n564 585
R152 B.n563 B.n106 585
R153 B.n562 B.n561 585
R154 B.n560 B.n107 585
R155 B.n559 B.n558 585
R156 B.n557 B.n108 585
R157 B.n556 B.n555 585
R158 B.n554 B.n109 585
R159 B.n553 B.n552 585
R160 B.n551 B.n110 585
R161 B.n550 B.n549 585
R162 B.n548 B.n111 585
R163 B.n547 B.n546 585
R164 B.n545 B.n112 585
R165 B.n544 B.n543 585
R166 B.n542 B.n113 585
R167 B.n541 B.n540 585
R168 B.n539 B.n114 585
R169 B.n538 B.n537 585
R170 B.n536 B.n115 585
R171 B.n535 B.n534 585
R172 B.n533 B.n116 585
R173 B.n532 B.n531 585
R174 B.n530 B.n117 585
R175 B.n529 B.n528 585
R176 B.n527 B.n118 585
R177 B.n526 B.n525 585
R178 B.n524 B.n119 585
R179 B.n523 B.n522 585
R180 B.n521 B.n120 585
R181 B.n520 B.n519 585
R182 B.n518 B.n121 585
R183 B.n517 B.n516 585
R184 B.n515 B.n122 585
R185 B.n514 B.n513 585
R186 B.n512 B.n123 585
R187 B.n511 B.n510 585
R188 B.n509 B.n124 585
R189 B.n508 B.n507 585
R190 B.n506 B.n125 585
R191 B.n505 B.n504 585
R192 B.n503 B.n126 585
R193 B.n502 B.n501 585
R194 B.n500 B.n127 585
R195 B.n499 B.n498 585
R196 B.n497 B.n128 585
R197 B.n496 B.n495 585
R198 B.n494 B.n129 585
R199 B.n493 B.n492 585
R200 B.n491 B.n130 585
R201 B.n490 B.n489 585
R202 B.n488 B.n131 585
R203 B.n487 B.n486 585
R204 B.n485 B.n132 585
R205 B.n484 B.n483 585
R206 B.n482 B.n133 585
R207 B.n481 B.n480 585
R208 B.n479 B.n134 585
R209 B.n478 B.n477 585
R210 B.n476 B.n135 585
R211 B.n475 B.n474 585
R212 B.n473 B.n136 585
R213 B.n472 B.n471 585
R214 B.n295 B.n294 585
R215 B.n296 B.n199 585
R216 B.n298 B.n297 585
R217 B.n299 B.n198 585
R218 B.n301 B.n300 585
R219 B.n302 B.n197 585
R220 B.n304 B.n303 585
R221 B.n305 B.n196 585
R222 B.n307 B.n306 585
R223 B.n308 B.n195 585
R224 B.n310 B.n309 585
R225 B.n311 B.n194 585
R226 B.n313 B.n312 585
R227 B.n314 B.n193 585
R228 B.n316 B.n315 585
R229 B.n317 B.n192 585
R230 B.n319 B.n318 585
R231 B.n320 B.n191 585
R232 B.n322 B.n321 585
R233 B.n323 B.n190 585
R234 B.n325 B.n324 585
R235 B.n326 B.n189 585
R236 B.n328 B.n327 585
R237 B.n329 B.n188 585
R238 B.n331 B.n330 585
R239 B.n332 B.n187 585
R240 B.n334 B.n333 585
R241 B.n335 B.n186 585
R242 B.n337 B.n336 585
R243 B.n338 B.n185 585
R244 B.n340 B.n339 585
R245 B.n341 B.n184 585
R246 B.n343 B.n342 585
R247 B.n344 B.n183 585
R248 B.n346 B.n345 585
R249 B.n347 B.n182 585
R250 B.n349 B.n348 585
R251 B.n350 B.n181 585
R252 B.n352 B.n351 585
R253 B.n353 B.n180 585
R254 B.n355 B.n354 585
R255 B.n356 B.n179 585
R256 B.n358 B.n357 585
R257 B.n359 B.n178 585
R258 B.n361 B.n360 585
R259 B.n362 B.n177 585
R260 B.n364 B.n363 585
R261 B.n365 B.n176 585
R262 B.n367 B.n366 585
R263 B.n368 B.n175 585
R264 B.n370 B.n369 585
R265 B.n371 B.n174 585
R266 B.n373 B.n372 585
R267 B.n374 B.n171 585
R268 B.n377 B.n376 585
R269 B.n378 B.n170 585
R270 B.n380 B.n379 585
R271 B.n381 B.n169 585
R272 B.n383 B.n382 585
R273 B.n384 B.n168 585
R274 B.n386 B.n385 585
R275 B.n387 B.n167 585
R276 B.n389 B.n388 585
R277 B.n391 B.n390 585
R278 B.n392 B.n163 585
R279 B.n394 B.n393 585
R280 B.n395 B.n162 585
R281 B.n397 B.n396 585
R282 B.n398 B.n161 585
R283 B.n400 B.n399 585
R284 B.n401 B.n160 585
R285 B.n403 B.n402 585
R286 B.n404 B.n159 585
R287 B.n406 B.n405 585
R288 B.n407 B.n158 585
R289 B.n409 B.n408 585
R290 B.n410 B.n157 585
R291 B.n412 B.n411 585
R292 B.n413 B.n156 585
R293 B.n415 B.n414 585
R294 B.n416 B.n155 585
R295 B.n418 B.n417 585
R296 B.n419 B.n154 585
R297 B.n421 B.n420 585
R298 B.n422 B.n153 585
R299 B.n424 B.n423 585
R300 B.n425 B.n152 585
R301 B.n427 B.n426 585
R302 B.n428 B.n151 585
R303 B.n430 B.n429 585
R304 B.n431 B.n150 585
R305 B.n433 B.n432 585
R306 B.n434 B.n149 585
R307 B.n436 B.n435 585
R308 B.n437 B.n148 585
R309 B.n439 B.n438 585
R310 B.n440 B.n147 585
R311 B.n442 B.n441 585
R312 B.n443 B.n146 585
R313 B.n445 B.n444 585
R314 B.n446 B.n145 585
R315 B.n448 B.n447 585
R316 B.n449 B.n144 585
R317 B.n451 B.n450 585
R318 B.n452 B.n143 585
R319 B.n454 B.n453 585
R320 B.n455 B.n142 585
R321 B.n457 B.n456 585
R322 B.n458 B.n141 585
R323 B.n460 B.n459 585
R324 B.n461 B.n140 585
R325 B.n463 B.n462 585
R326 B.n464 B.n139 585
R327 B.n466 B.n465 585
R328 B.n467 B.n138 585
R329 B.n469 B.n468 585
R330 B.n470 B.n137 585
R331 B.n293 B.n200 585
R332 B.n292 B.n291 585
R333 B.n290 B.n201 585
R334 B.n289 B.n288 585
R335 B.n287 B.n202 585
R336 B.n286 B.n285 585
R337 B.n284 B.n203 585
R338 B.n283 B.n282 585
R339 B.n281 B.n204 585
R340 B.n280 B.n279 585
R341 B.n278 B.n205 585
R342 B.n277 B.n276 585
R343 B.n275 B.n206 585
R344 B.n274 B.n273 585
R345 B.n272 B.n207 585
R346 B.n271 B.n270 585
R347 B.n269 B.n208 585
R348 B.n268 B.n267 585
R349 B.n266 B.n209 585
R350 B.n265 B.n264 585
R351 B.n263 B.n210 585
R352 B.n262 B.n261 585
R353 B.n260 B.n211 585
R354 B.n259 B.n258 585
R355 B.n257 B.n212 585
R356 B.n256 B.n255 585
R357 B.n254 B.n213 585
R358 B.n253 B.n252 585
R359 B.n251 B.n214 585
R360 B.n250 B.n249 585
R361 B.n248 B.n215 585
R362 B.n247 B.n246 585
R363 B.n245 B.n216 585
R364 B.n244 B.n243 585
R365 B.n242 B.n217 585
R366 B.n241 B.n240 585
R367 B.n239 B.n218 585
R368 B.n238 B.n237 585
R369 B.n236 B.n219 585
R370 B.n235 B.n234 585
R371 B.n233 B.n220 585
R372 B.n232 B.n231 585
R373 B.n230 B.n221 585
R374 B.n229 B.n228 585
R375 B.n227 B.n222 585
R376 B.n226 B.n225 585
R377 B.n224 B.n223 585
R378 B.n2 B.n0 585
R379 B.n865 B.n1 585
R380 B.n864 B.n863 585
R381 B.n862 B.n3 585
R382 B.n861 B.n860 585
R383 B.n859 B.n4 585
R384 B.n858 B.n857 585
R385 B.n856 B.n5 585
R386 B.n855 B.n854 585
R387 B.n853 B.n6 585
R388 B.n852 B.n851 585
R389 B.n850 B.n7 585
R390 B.n849 B.n848 585
R391 B.n847 B.n8 585
R392 B.n846 B.n845 585
R393 B.n844 B.n9 585
R394 B.n843 B.n842 585
R395 B.n841 B.n10 585
R396 B.n840 B.n839 585
R397 B.n838 B.n11 585
R398 B.n837 B.n836 585
R399 B.n835 B.n12 585
R400 B.n834 B.n833 585
R401 B.n832 B.n13 585
R402 B.n831 B.n830 585
R403 B.n829 B.n14 585
R404 B.n828 B.n827 585
R405 B.n826 B.n15 585
R406 B.n825 B.n824 585
R407 B.n823 B.n16 585
R408 B.n822 B.n821 585
R409 B.n820 B.n17 585
R410 B.n819 B.n818 585
R411 B.n817 B.n18 585
R412 B.n816 B.n815 585
R413 B.n814 B.n19 585
R414 B.n813 B.n812 585
R415 B.n811 B.n20 585
R416 B.n810 B.n809 585
R417 B.n808 B.n21 585
R418 B.n807 B.n806 585
R419 B.n805 B.n22 585
R420 B.n804 B.n803 585
R421 B.n802 B.n23 585
R422 B.n801 B.n800 585
R423 B.n799 B.n24 585
R424 B.n798 B.n797 585
R425 B.n796 B.n25 585
R426 B.n795 B.n794 585
R427 B.n867 B.n866 585
R428 B.n294 B.n293 550.159
R429 B.n794 B.n793 550.159
R430 B.n472 B.n137 550.159
R431 B.n617 B.n616 550.159
R432 B.n164 B.t11 494.592
R433 B.n60 B.t7 494.592
R434 B.n172 B.t5 494.592
R435 B.n54 B.t1 494.592
R436 B.n165 B.t10 450.568
R437 B.n61 B.t8 450.568
R438 B.n173 B.t4 450.568
R439 B.n55 B.t2 450.568
R440 B.n164 B.t9 407.524
R441 B.n172 B.t3 407.524
R442 B.n54 B.t0 407.524
R443 B.n60 B.t6 407.524
R444 B.n293 B.n292 163.367
R445 B.n292 B.n201 163.367
R446 B.n288 B.n201 163.367
R447 B.n288 B.n287 163.367
R448 B.n287 B.n286 163.367
R449 B.n286 B.n203 163.367
R450 B.n282 B.n203 163.367
R451 B.n282 B.n281 163.367
R452 B.n281 B.n280 163.367
R453 B.n280 B.n205 163.367
R454 B.n276 B.n205 163.367
R455 B.n276 B.n275 163.367
R456 B.n275 B.n274 163.367
R457 B.n274 B.n207 163.367
R458 B.n270 B.n207 163.367
R459 B.n270 B.n269 163.367
R460 B.n269 B.n268 163.367
R461 B.n268 B.n209 163.367
R462 B.n264 B.n209 163.367
R463 B.n264 B.n263 163.367
R464 B.n263 B.n262 163.367
R465 B.n262 B.n211 163.367
R466 B.n258 B.n211 163.367
R467 B.n258 B.n257 163.367
R468 B.n257 B.n256 163.367
R469 B.n256 B.n213 163.367
R470 B.n252 B.n213 163.367
R471 B.n252 B.n251 163.367
R472 B.n251 B.n250 163.367
R473 B.n250 B.n215 163.367
R474 B.n246 B.n215 163.367
R475 B.n246 B.n245 163.367
R476 B.n245 B.n244 163.367
R477 B.n244 B.n217 163.367
R478 B.n240 B.n217 163.367
R479 B.n240 B.n239 163.367
R480 B.n239 B.n238 163.367
R481 B.n238 B.n219 163.367
R482 B.n234 B.n219 163.367
R483 B.n234 B.n233 163.367
R484 B.n233 B.n232 163.367
R485 B.n232 B.n221 163.367
R486 B.n228 B.n221 163.367
R487 B.n228 B.n227 163.367
R488 B.n227 B.n226 163.367
R489 B.n226 B.n223 163.367
R490 B.n223 B.n2 163.367
R491 B.n866 B.n2 163.367
R492 B.n866 B.n865 163.367
R493 B.n865 B.n864 163.367
R494 B.n864 B.n3 163.367
R495 B.n860 B.n3 163.367
R496 B.n860 B.n859 163.367
R497 B.n859 B.n858 163.367
R498 B.n858 B.n5 163.367
R499 B.n854 B.n5 163.367
R500 B.n854 B.n853 163.367
R501 B.n853 B.n852 163.367
R502 B.n852 B.n7 163.367
R503 B.n848 B.n7 163.367
R504 B.n848 B.n847 163.367
R505 B.n847 B.n846 163.367
R506 B.n846 B.n9 163.367
R507 B.n842 B.n9 163.367
R508 B.n842 B.n841 163.367
R509 B.n841 B.n840 163.367
R510 B.n840 B.n11 163.367
R511 B.n836 B.n11 163.367
R512 B.n836 B.n835 163.367
R513 B.n835 B.n834 163.367
R514 B.n834 B.n13 163.367
R515 B.n830 B.n13 163.367
R516 B.n830 B.n829 163.367
R517 B.n829 B.n828 163.367
R518 B.n828 B.n15 163.367
R519 B.n824 B.n15 163.367
R520 B.n824 B.n823 163.367
R521 B.n823 B.n822 163.367
R522 B.n822 B.n17 163.367
R523 B.n818 B.n17 163.367
R524 B.n818 B.n817 163.367
R525 B.n817 B.n816 163.367
R526 B.n816 B.n19 163.367
R527 B.n812 B.n19 163.367
R528 B.n812 B.n811 163.367
R529 B.n811 B.n810 163.367
R530 B.n810 B.n21 163.367
R531 B.n806 B.n21 163.367
R532 B.n806 B.n805 163.367
R533 B.n805 B.n804 163.367
R534 B.n804 B.n23 163.367
R535 B.n800 B.n23 163.367
R536 B.n800 B.n799 163.367
R537 B.n799 B.n798 163.367
R538 B.n798 B.n25 163.367
R539 B.n794 B.n25 163.367
R540 B.n294 B.n199 163.367
R541 B.n298 B.n199 163.367
R542 B.n299 B.n298 163.367
R543 B.n300 B.n299 163.367
R544 B.n300 B.n197 163.367
R545 B.n304 B.n197 163.367
R546 B.n305 B.n304 163.367
R547 B.n306 B.n305 163.367
R548 B.n306 B.n195 163.367
R549 B.n310 B.n195 163.367
R550 B.n311 B.n310 163.367
R551 B.n312 B.n311 163.367
R552 B.n312 B.n193 163.367
R553 B.n316 B.n193 163.367
R554 B.n317 B.n316 163.367
R555 B.n318 B.n317 163.367
R556 B.n318 B.n191 163.367
R557 B.n322 B.n191 163.367
R558 B.n323 B.n322 163.367
R559 B.n324 B.n323 163.367
R560 B.n324 B.n189 163.367
R561 B.n328 B.n189 163.367
R562 B.n329 B.n328 163.367
R563 B.n330 B.n329 163.367
R564 B.n330 B.n187 163.367
R565 B.n334 B.n187 163.367
R566 B.n335 B.n334 163.367
R567 B.n336 B.n335 163.367
R568 B.n336 B.n185 163.367
R569 B.n340 B.n185 163.367
R570 B.n341 B.n340 163.367
R571 B.n342 B.n341 163.367
R572 B.n342 B.n183 163.367
R573 B.n346 B.n183 163.367
R574 B.n347 B.n346 163.367
R575 B.n348 B.n347 163.367
R576 B.n348 B.n181 163.367
R577 B.n352 B.n181 163.367
R578 B.n353 B.n352 163.367
R579 B.n354 B.n353 163.367
R580 B.n354 B.n179 163.367
R581 B.n358 B.n179 163.367
R582 B.n359 B.n358 163.367
R583 B.n360 B.n359 163.367
R584 B.n360 B.n177 163.367
R585 B.n364 B.n177 163.367
R586 B.n365 B.n364 163.367
R587 B.n366 B.n365 163.367
R588 B.n366 B.n175 163.367
R589 B.n370 B.n175 163.367
R590 B.n371 B.n370 163.367
R591 B.n372 B.n371 163.367
R592 B.n372 B.n171 163.367
R593 B.n377 B.n171 163.367
R594 B.n378 B.n377 163.367
R595 B.n379 B.n378 163.367
R596 B.n379 B.n169 163.367
R597 B.n383 B.n169 163.367
R598 B.n384 B.n383 163.367
R599 B.n385 B.n384 163.367
R600 B.n385 B.n167 163.367
R601 B.n389 B.n167 163.367
R602 B.n390 B.n389 163.367
R603 B.n390 B.n163 163.367
R604 B.n394 B.n163 163.367
R605 B.n395 B.n394 163.367
R606 B.n396 B.n395 163.367
R607 B.n396 B.n161 163.367
R608 B.n400 B.n161 163.367
R609 B.n401 B.n400 163.367
R610 B.n402 B.n401 163.367
R611 B.n402 B.n159 163.367
R612 B.n406 B.n159 163.367
R613 B.n407 B.n406 163.367
R614 B.n408 B.n407 163.367
R615 B.n408 B.n157 163.367
R616 B.n412 B.n157 163.367
R617 B.n413 B.n412 163.367
R618 B.n414 B.n413 163.367
R619 B.n414 B.n155 163.367
R620 B.n418 B.n155 163.367
R621 B.n419 B.n418 163.367
R622 B.n420 B.n419 163.367
R623 B.n420 B.n153 163.367
R624 B.n424 B.n153 163.367
R625 B.n425 B.n424 163.367
R626 B.n426 B.n425 163.367
R627 B.n426 B.n151 163.367
R628 B.n430 B.n151 163.367
R629 B.n431 B.n430 163.367
R630 B.n432 B.n431 163.367
R631 B.n432 B.n149 163.367
R632 B.n436 B.n149 163.367
R633 B.n437 B.n436 163.367
R634 B.n438 B.n437 163.367
R635 B.n438 B.n147 163.367
R636 B.n442 B.n147 163.367
R637 B.n443 B.n442 163.367
R638 B.n444 B.n443 163.367
R639 B.n444 B.n145 163.367
R640 B.n448 B.n145 163.367
R641 B.n449 B.n448 163.367
R642 B.n450 B.n449 163.367
R643 B.n450 B.n143 163.367
R644 B.n454 B.n143 163.367
R645 B.n455 B.n454 163.367
R646 B.n456 B.n455 163.367
R647 B.n456 B.n141 163.367
R648 B.n460 B.n141 163.367
R649 B.n461 B.n460 163.367
R650 B.n462 B.n461 163.367
R651 B.n462 B.n139 163.367
R652 B.n466 B.n139 163.367
R653 B.n467 B.n466 163.367
R654 B.n468 B.n467 163.367
R655 B.n468 B.n137 163.367
R656 B.n473 B.n472 163.367
R657 B.n474 B.n473 163.367
R658 B.n474 B.n135 163.367
R659 B.n478 B.n135 163.367
R660 B.n479 B.n478 163.367
R661 B.n480 B.n479 163.367
R662 B.n480 B.n133 163.367
R663 B.n484 B.n133 163.367
R664 B.n485 B.n484 163.367
R665 B.n486 B.n485 163.367
R666 B.n486 B.n131 163.367
R667 B.n490 B.n131 163.367
R668 B.n491 B.n490 163.367
R669 B.n492 B.n491 163.367
R670 B.n492 B.n129 163.367
R671 B.n496 B.n129 163.367
R672 B.n497 B.n496 163.367
R673 B.n498 B.n497 163.367
R674 B.n498 B.n127 163.367
R675 B.n502 B.n127 163.367
R676 B.n503 B.n502 163.367
R677 B.n504 B.n503 163.367
R678 B.n504 B.n125 163.367
R679 B.n508 B.n125 163.367
R680 B.n509 B.n508 163.367
R681 B.n510 B.n509 163.367
R682 B.n510 B.n123 163.367
R683 B.n514 B.n123 163.367
R684 B.n515 B.n514 163.367
R685 B.n516 B.n515 163.367
R686 B.n516 B.n121 163.367
R687 B.n520 B.n121 163.367
R688 B.n521 B.n520 163.367
R689 B.n522 B.n521 163.367
R690 B.n522 B.n119 163.367
R691 B.n526 B.n119 163.367
R692 B.n527 B.n526 163.367
R693 B.n528 B.n527 163.367
R694 B.n528 B.n117 163.367
R695 B.n532 B.n117 163.367
R696 B.n533 B.n532 163.367
R697 B.n534 B.n533 163.367
R698 B.n534 B.n115 163.367
R699 B.n538 B.n115 163.367
R700 B.n539 B.n538 163.367
R701 B.n540 B.n539 163.367
R702 B.n540 B.n113 163.367
R703 B.n544 B.n113 163.367
R704 B.n545 B.n544 163.367
R705 B.n546 B.n545 163.367
R706 B.n546 B.n111 163.367
R707 B.n550 B.n111 163.367
R708 B.n551 B.n550 163.367
R709 B.n552 B.n551 163.367
R710 B.n552 B.n109 163.367
R711 B.n556 B.n109 163.367
R712 B.n557 B.n556 163.367
R713 B.n558 B.n557 163.367
R714 B.n558 B.n107 163.367
R715 B.n562 B.n107 163.367
R716 B.n563 B.n562 163.367
R717 B.n564 B.n563 163.367
R718 B.n564 B.n105 163.367
R719 B.n568 B.n105 163.367
R720 B.n569 B.n568 163.367
R721 B.n570 B.n569 163.367
R722 B.n570 B.n103 163.367
R723 B.n574 B.n103 163.367
R724 B.n575 B.n574 163.367
R725 B.n576 B.n575 163.367
R726 B.n576 B.n101 163.367
R727 B.n580 B.n101 163.367
R728 B.n581 B.n580 163.367
R729 B.n582 B.n581 163.367
R730 B.n582 B.n99 163.367
R731 B.n586 B.n99 163.367
R732 B.n587 B.n586 163.367
R733 B.n588 B.n587 163.367
R734 B.n588 B.n97 163.367
R735 B.n592 B.n97 163.367
R736 B.n593 B.n592 163.367
R737 B.n594 B.n593 163.367
R738 B.n594 B.n95 163.367
R739 B.n598 B.n95 163.367
R740 B.n599 B.n598 163.367
R741 B.n600 B.n599 163.367
R742 B.n600 B.n93 163.367
R743 B.n604 B.n93 163.367
R744 B.n605 B.n604 163.367
R745 B.n606 B.n605 163.367
R746 B.n606 B.n91 163.367
R747 B.n610 B.n91 163.367
R748 B.n611 B.n610 163.367
R749 B.n612 B.n611 163.367
R750 B.n612 B.n89 163.367
R751 B.n616 B.n89 163.367
R752 B.n793 B.n792 163.367
R753 B.n792 B.n27 163.367
R754 B.n788 B.n27 163.367
R755 B.n788 B.n787 163.367
R756 B.n787 B.n786 163.367
R757 B.n786 B.n29 163.367
R758 B.n782 B.n29 163.367
R759 B.n782 B.n781 163.367
R760 B.n781 B.n780 163.367
R761 B.n780 B.n31 163.367
R762 B.n776 B.n31 163.367
R763 B.n776 B.n775 163.367
R764 B.n775 B.n774 163.367
R765 B.n774 B.n33 163.367
R766 B.n770 B.n33 163.367
R767 B.n770 B.n769 163.367
R768 B.n769 B.n768 163.367
R769 B.n768 B.n35 163.367
R770 B.n764 B.n35 163.367
R771 B.n764 B.n763 163.367
R772 B.n763 B.n762 163.367
R773 B.n762 B.n37 163.367
R774 B.n758 B.n37 163.367
R775 B.n758 B.n757 163.367
R776 B.n757 B.n756 163.367
R777 B.n756 B.n39 163.367
R778 B.n752 B.n39 163.367
R779 B.n752 B.n751 163.367
R780 B.n751 B.n750 163.367
R781 B.n750 B.n41 163.367
R782 B.n746 B.n41 163.367
R783 B.n746 B.n745 163.367
R784 B.n745 B.n744 163.367
R785 B.n744 B.n43 163.367
R786 B.n740 B.n43 163.367
R787 B.n740 B.n739 163.367
R788 B.n739 B.n738 163.367
R789 B.n738 B.n45 163.367
R790 B.n734 B.n45 163.367
R791 B.n734 B.n733 163.367
R792 B.n733 B.n732 163.367
R793 B.n732 B.n47 163.367
R794 B.n728 B.n47 163.367
R795 B.n728 B.n727 163.367
R796 B.n727 B.n726 163.367
R797 B.n726 B.n49 163.367
R798 B.n722 B.n49 163.367
R799 B.n722 B.n721 163.367
R800 B.n721 B.n720 163.367
R801 B.n720 B.n51 163.367
R802 B.n716 B.n51 163.367
R803 B.n716 B.n715 163.367
R804 B.n715 B.n714 163.367
R805 B.n714 B.n53 163.367
R806 B.n709 B.n53 163.367
R807 B.n709 B.n708 163.367
R808 B.n708 B.n707 163.367
R809 B.n707 B.n57 163.367
R810 B.n703 B.n57 163.367
R811 B.n703 B.n702 163.367
R812 B.n702 B.n701 163.367
R813 B.n701 B.n59 163.367
R814 B.n696 B.n59 163.367
R815 B.n696 B.n695 163.367
R816 B.n695 B.n694 163.367
R817 B.n694 B.n63 163.367
R818 B.n690 B.n63 163.367
R819 B.n690 B.n689 163.367
R820 B.n689 B.n688 163.367
R821 B.n688 B.n65 163.367
R822 B.n684 B.n65 163.367
R823 B.n684 B.n683 163.367
R824 B.n683 B.n682 163.367
R825 B.n682 B.n67 163.367
R826 B.n678 B.n67 163.367
R827 B.n678 B.n677 163.367
R828 B.n677 B.n676 163.367
R829 B.n676 B.n69 163.367
R830 B.n672 B.n69 163.367
R831 B.n672 B.n671 163.367
R832 B.n671 B.n670 163.367
R833 B.n670 B.n71 163.367
R834 B.n666 B.n71 163.367
R835 B.n666 B.n665 163.367
R836 B.n665 B.n664 163.367
R837 B.n664 B.n73 163.367
R838 B.n660 B.n73 163.367
R839 B.n660 B.n659 163.367
R840 B.n659 B.n658 163.367
R841 B.n658 B.n75 163.367
R842 B.n654 B.n75 163.367
R843 B.n654 B.n653 163.367
R844 B.n653 B.n652 163.367
R845 B.n652 B.n77 163.367
R846 B.n648 B.n77 163.367
R847 B.n648 B.n647 163.367
R848 B.n647 B.n646 163.367
R849 B.n646 B.n79 163.367
R850 B.n642 B.n79 163.367
R851 B.n642 B.n641 163.367
R852 B.n641 B.n640 163.367
R853 B.n640 B.n81 163.367
R854 B.n636 B.n81 163.367
R855 B.n636 B.n635 163.367
R856 B.n635 B.n634 163.367
R857 B.n634 B.n83 163.367
R858 B.n630 B.n83 163.367
R859 B.n630 B.n629 163.367
R860 B.n629 B.n628 163.367
R861 B.n628 B.n85 163.367
R862 B.n624 B.n85 163.367
R863 B.n624 B.n623 163.367
R864 B.n623 B.n622 163.367
R865 B.n622 B.n87 163.367
R866 B.n618 B.n87 163.367
R867 B.n618 B.n617 163.367
R868 B.n166 B.n165 59.5399
R869 B.n375 B.n173 59.5399
R870 B.n712 B.n55 59.5399
R871 B.n698 B.n61 59.5399
R872 B.n165 B.n164 44.0247
R873 B.n173 B.n172 44.0247
R874 B.n55 B.n54 44.0247
R875 B.n61 B.n60 44.0247
R876 B.n795 B.n26 35.7468
R877 B.n615 B.n88 35.7468
R878 B.n471 B.n470 35.7468
R879 B.n295 B.n200 35.7468
R880 B B.n867 18.0485
R881 B.n791 B.n26 10.6151
R882 B.n791 B.n790 10.6151
R883 B.n790 B.n789 10.6151
R884 B.n789 B.n28 10.6151
R885 B.n785 B.n28 10.6151
R886 B.n785 B.n784 10.6151
R887 B.n784 B.n783 10.6151
R888 B.n783 B.n30 10.6151
R889 B.n779 B.n30 10.6151
R890 B.n779 B.n778 10.6151
R891 B.n778 B.n777 10.6151
R892 B.n777 B.n32 10.6151
R893 B.n773 B.n32 10.6151
R894 B.n773 B.n772 10.6151
R895 B.n772 B.n771 10.6151
R896 B.n771 B.n34 10.6151
R897 B.n767 B.n34 10.6151
R898 B.n767 B.n766 10.6151
R899 B.n766 B.n765 10.6151
R900 B.n765 B.n36 10.6151
R901 B.n761 B.n36 10.6151
R902 B.n761 B.n760 10.6151
R903 B.n760 B.n759 10.6151
R904 B.n759 B.n38 10.6151
R905 B.n755 B.n38 10.6151
R906 B.n755 B.n754 10.6151
R907 B.n754 B.n753 10.6151
R908 B.n753 B.n40 10.6151
R909 B.n749 B.n40 10.6151
R910 B.n749 B.n748 10.6151
R911 B.n748 B.n747 10.6151
R912 B.n747 B.n42 10.6151
R913 B.n743 B.n42 10.6151
R914 B.n743 B.n742 10.6151
R915 B.n742 B.n741 10.6151
R916 B.n741 B.n44 10.6151
R917 B.n737 B.n44 10.6151
R918 B.n737 B.n736 10.6151
R919 B.n736 B.n735 10.6151
R920 B.n735 B.n46 10.6151
R921 B.n731 B.n46 10.6151
R922 B.n731 B.n730 10.6151
R923 B.n730 B.n729 10.6151
R924 B.n729 B.n48 10.6151
R925 B.n725 B.n48 10.6151
R926 B.n725 B.n724 10.6151
R927 B.n724 B.n723 10.6151
R928 B.n723 B.n50 10.6151
R929 B.n719 B.n50 10.6151
R930 B.n719 B.n718 10.6151
R931 B.n718 B.n717 10.6151
R932 B.n717 B.n52 10.6151
R933 B.n713 B.n52 10.6151
R934 B.n711 B.n710 10.6151
R935 B.n710 B.n56 10.6151
R936 B.n706 B.n56 10.6151
R937 B.n706 B.n705 10.6151
R938 B.n705 B.n704 10.6151
R939 B.n704 B.n58 10.6151
R940 B.n700 B.n58 10.6151
R941 B.n700 B.n699 10.6151
R942 B.n697 B.n62 10.6151
R943 B.n693 B.n62 10.6151
R944 B.n693 B.n692 10.6151
R945 B.n692 B.n691 10.6151
R946 B.n691 B.n64 10.6151
R947 B.n687 B.n64 10.6151
R948 B.n687 B.n686 10.6151
R949 B.n686 B.n685 10.6151
R950 B.n685 B.n66 10.6151
R951 B.n681 B.n66 10.6151
R952 B.n681 B.n680 10.6151
R953 B.n680 B.n679 10.6151
R954 B.n679 B.n68 10.6151
R955 B.n675 B.n68 10.6151
R956 B.n675 B.n674 10.6151
R957 B.n674 B.n673 10.6151
R958 B.n673 B.n70 10.6151
R959 B.n669 B.n70 10.6151
R960 B.n669 B.n668 10.6151
R961 B.n668 B.n667 10.6151
R962 B.n667 B.n72 10.6151
R963 B.n663 B.n72 10.6151
R964 B.n663 B.n662 10.6151
R965 B.n662 B.n661 10.6151
R966 B.n661 B.n74 10.6151
R967 B.n657 B.n74 10.6151
R968 B.n657 B.n656 10.6151
R969 B.n656 B.n655 10.6151
R970 B.n655 B.n76 10.6151
R971 B.n651 B.n76 10.6151
R972 B.n651 B.n650 10.6151
R973 B.n650 B.n649 10.6151
R974 B.n649 B.n78 10.6151
R975 B.n645 B.n78 10.6151
R976 B.n645 B.n644 10.6151
R977 B.n644 B.n643 10.6151
R978 B.n643 B.n80 10.6151
R979 B.n639 B.n80 10.6151
R980 B.n639 B.n638 10.6151
R981 B.n638 B.n637 10.6151
R982 B.n637 B.n82 10.6151
R983 B.n633 B.n82 10.6151
R984 B.n633 B.n632 10.6151
R985 B.n632 B.n631 10.6151
R986 B.n631 B.n84 10.6151
R987 B.n627 B.n84 10.6151
R988 B.n627 B.n626 10.6151
R989 B.n626 B.n625 10.6151
R990 B.n625 B.n86 10.6151
R991 B.n621 B.n86 10.6151
R992 B.n621 B.n620 10.6151
R993 B.n620 B.n619 10.6151
R994 B.n619 B.n88 10.6151
R995 B.n471 B.n136 10.6151
R996 B.n475 B.n136 10.6151
R997 B.n476 B.n475 10.6151
R998 B.n477 B.n476 10.6151
R999 B.n477 B.n134 10.6151
R1000 B.n481 B.n134 10.6151
R1001 B.n482 B.n481 10.6151
R1002 B.n483 B.n482 10.6151
R1003 B.n483 B.n132 10.6151
R1004 B.n487 B.n132 10.6151
R1005 B.n488 B.n487 10.6151
R1006 B.n489 B.n488 10.6151
R1007 B.n489 B.n130 10.6151
R1008 B.n493 B.n130 10.6151
R1009 B.n494 B.n493 10.6151
R1010 B.n495 B.n494 10.6151
R1011 B.n495 B.n128 10.6151
R1012 B.n499 B.n128 10.6151
R1013 B.n500 B.n499 10.6151
R1014 B.n501 B.n500 10.6151
R1015 B.n501 B.n126 10.6151
R1016 B.n505 B.n126 10.6151
R1017 B.n506 B.n505 10.6151
R1018 B.n507 B.n506 10.6151
R1019 B.n507 B.n124 10.6151
R1020 B.n511 B.n124 10.6151
R1021 B.n512 B.n511 10.6151
R1022 B.n513 B.n512 10.6151
R1023 B.n513 B.n122 10.6151
R1024 B.n517 B.n122 10.6151
R1025 B.n518 B.n517 10.6151
R1026 B.n519 B.n518 10.6151
R1027 B.n519 B.n120 10.6151
R1028 B.n523 B.n120 10.6151
R1029 B.n524 B.n523 10.6151
R1030 B.n525 B.n524 10.6151
R1031 B.n525 B.n118 10.6151
R1032 B.n529 B.n118 10.6151
R1033 B.n530 B.n529 10.6151
R1034 B.n531 B.n530 10.6151
R1035 B.n531 B.n116 10.6151
R1036 B.n535 B.n116 10.6151
R1037 B.n536 B.n535 10.6151
R1038 B.n537 B.n536 10.6151
R1039 B.n537 B.n114 10.6151
R1040 B.n541 B.n114 10.6151
R1041 B.n542 B.n541 10.6151
R1042 B.n543 B.n542 10.6151
R1043 B.n543 B.n112 10.6151
R1044 B.n547 B.n112 10.6151
R1045 B.n548 B.n547 10.6151
R1046 B.n549 B.n548 10.6151
R1047 B.n549 B.n110 10.6151
R1048 B.n553 B.n110 10.6151
R1049 B.n554 B.n553 10.6151
R1050 B.n555 B.n554 10.6151
R1051 B.n555 B.n108 10.6151
R1052 B.n559 B.n108 10.6151
R1053 B.n560 B.n559 10.6151
R1054 B.n561 B.n560 10.6151
R1055 B.n561 B.n106 10.6151
R1056 B.n565 B.n106 10.6151
R1057 B.n566 B.n565 10.6151
R1058 B.n567 B.n566 10.6151
R1059 B.n567 B.n104 10.6151
R1060 B.n571 B.n104 10.6151
R1061 B.n572 B.n571 10.6151
R1062 B.n573 B.n572 10.6151
R1063 B.n573 B.n102 10.6151
R1064 B.n577 B.n102 10.6151
R1065 B.n578 B.n577 10.6151
R1066 B.n579 B.n578 10.6151
R1067 B.n579 B.n100 10.6151
R1068 B.n583 B.n100 10.6151
R1069 B.n584 B.n583 10.6151
R1070 B.n585 B.n584 10.6151
R1071 B.n585 B.n98 10.6151
R1072 B.n589 B.n98 10.6151
R1073 B.n590 B.n589 10.6151
R1074 B.n591 B.n590 10.6151
R1075 B.n591 B.n96 10.6151
R1076 B.n595 B.n96 10.6151
R1077 B.n596 B.n595 10.6151
R1078 B.n597 B.n596 10.6151
R1079 B.n597 B.n94 10.6151
R1080 B.n601 B.n94 10.6151
R1081 B.n602 B.n601 10.6151
R1082 B.n603 B.n602 10.6151
R1083 B.n603 B.n92 10.6151
R1084 B.n607 B.n92 10.6151
R1085 B.n608 B.n607 10.6151
R1086 B.n609 B.n608 10.6151
R1087 B.n609 B.n90 10.6151
R1088 B.n613 B.n90 10.6151
R1089 B.n614 B.n613 10.6151
R1090 B.n615 B.n614 10.6151
R1091 B.n296 B.n295 10.6151
R1092 B.n297 B.n296 10.6151
R1093 B.n297 B.n198 10.6151
R1094 B.n301 B.n198 10.6151
R1095 B.n302 B.n301 10.6151
R1096 B.n303 B.n302 10.6151
R1097 B.n303 B.n196 10.6151
R1098 B.n307 B.n196 10.6151
R1099 B.n308 B.n307 10.6151
R1100 B.n309 B.n308 10.6151
R1101 B.n309 B.n194 10.6151
R1102 B.n313 B.n194 10.6151
R1103 B.n314 B.n313 10.6151
R1104 B.n315 B.n314 10.6151
R1105 B.n315 B.n192 10.6151
R1106 B.n319 B.n192 10.6151
R1107 B.n320 B.n319 10.6151
R1108 B.n321 B.n320 10.6151
R1109 B.n321 B.n190 10.6151
R1110 B.n325 B.n190 10.6151
R1111 B.n326 B.n325 10.6151
R1112 B.n327 B.n326 10.6151
R1113 B.n327 B.n188 10.6151
R1114 B.n331 B.n188 10.6151
R1115 B.n332 B.n331 10.6151
R1116 B.n333 B.n332 10.6151
R1117 B.n333 B.n186 10.6151
R1118 B.n337 B.n186 10.6151
R1119 B.n338 B.n337 10.6151
R1120 B.n339 B.n338 10.6151
R1121 B.n339 B.n184 10.6151
R1122 B.n343 B.n184 10.6151
R1123 B.n344 B.n343 10.6151
R1124 B.n345 B.n344 10.6151
R1125 B.n345 B.n182 10.6151
R1126 B.n349 B.n182 10.6151
R1127 B.n350 B.n349 10.6151
R1128 B.n351 B.n350 10.6151
R1129 B.n351 B.n180 10.6151
R1130 B.n355 B.n180 10.6151
R1131 B.n356 B.n355 10.6151
R1132 B.n357 B.n356 10.6151
R1133 B.n357 B.n178 10.6151
R1134 B.n361 B.n178 10.6151
R1135 B.n362 B.n361 10.6151
R1136 B.n363 B.n362 10.6151
R1137 B.n363 B.n176 10.6151
R1138 B.n367 B.n176 10.6151
R1139 B.n368 B.n367 10.6151
R1140 B.n369 B.n368 10.6151
R1141 B.n369 B.n174 10.6151
R1142 B.n373 B.n174 10.6151
R1143 B.n374 B.n373 10.6151
R1144 B.n376 B.n170 10.6151
R1145 B.n380 B.n170 10.6151
R1146 B.n381 B.n380 10.6151
R1147 B.n382 B.n381 10.6151
R1148 B.n382 B.n168 10.6151
R1149 B.n386 B.n168 10.6151
R1150 B.n387 B.n386 10.6151
R1151 B.n388 B.n387 10.6151
R1152 B.n392 B.n391 10.6151
R1153 B.n393 B.n392 10.6151
R1154 B.n393 B.n162 10.6151
R1155 B.n397 B.n162 10.6151
R1156 B.n398 B.n397 10.6151
R1157 B.n399 B.n398 10.6151
R1158 B.n399 B.n160 10.6151
R1159 B.n403 B.n160 10.6151
R1160 B.n404 B.n403 10.6151
R1161 B.n405 B.n404 10.6151
R1162 B.n405 B.n158 10.6151
R1163 B.n409 B.n158 10.6151
R1164 B.n410 B.n409 10.6151
R1165 B.n411 B.n410 10.6151
R1166 B.n411 B.n156 10.6151
R1167 B.n415 B.n156 10.6151
R1168 B.n416 B.n415 10.6151
R1169 B.n417 B.n416 10.6151
R1170 B.n417 B.n154 10.6151
R1171 B.n421 B.n154 10.6151
R1172 B.n422 B.n421 10.6151
R1173 B.n423 B.n422 10.6151
R1174 B.n423 B.n152 10.6151
R1175 B.n427 B.n152 10.6151
R1176 B.n428 B.n427 10.6151
R1177 B.n429 B.n428 10.6151
R1178 B.n429 B.n150 10.6151
R1179 B.n433 B.n150 10.6151
R1180 B.n434 B.n433 10.6151
R1181 B.n435 B.n434 10.6151
R1182 B.n435 B.n148 10.6151
R1183 B.n439 B.n148 10.6151
R1184 B.n440 B.n439 10.6151
R1185 B.n441 B.n440 10.6151
R1186 B.n441 B.n146 10.6151
R1187 B.n445 B.n146 10.6151
R1188 B.n446 B.n445 10.6151
R1189 B.n447 B.n446 10.6151
R1190 B.n447 B.n144 10.6151
R1191 B.n451 B.n144 10.6151
R1192 B.n452 B.n451 10.6151
R1193 B.n453 B.n452 10.6151
R1194 B.n453 B.n142 10.6151
R1195 B.n457 B.n142 10.6151
R1196 B.n458 B.n457 10.6151
R1197 B.n459 B.n458 10.6151
R1198 B.n459 B.n140 10.6151
R1199 B.n463 B.n140 10.6151
R1200 B.n464 B.n463 10.6151
R1201 B.n465 B.n464 10.6151
R1202 B.n465 B.n138 10.6151
R1203 B.n469 B.n138 10.6151
R1204 B.n470 B.n469 10.6151
R1205 B.n291 B.n200 10.6151
R1206 B.n291 B.n290 10.6151
R1207 B.n290 B.n289 10.6151
R1208 B.n289 B.n202 10.6151
R1209 B.n285 B.n202 10.6151
R1210 B.n285 B.n284 10.6151
R1211 B.n284 B.n283 10.6151
R1212 B.n283 B.n204 10.6151
R1213 B.n279 B.n204 10.6151
R1214 B.n279 B.n278 10.6151
R1215 B.n278 B.n277 10.6151
R1216 B.n277 B.n206 10.6151
R1217 B.n273 B.n206 10.6151
R1218 B.n273 B.n272 10.6151
R1219 B.n272 B.n271 10.6151
R1220 B.n271 B.n208 10.6151
R1221 B.n267 B.n208 10.6151
R1222 B.n267 B.n266 10.6151
R1223 B.n266 B.n265 10.6151
R1224 B.n265 B.n210 10.6151
R1225 B.n261 B.n210 10.6151
R1226 B.n261 B.n260 10.6151
R1227 B.n260 B.n259 10.6151
R1228 B.n259 B.n212 10.6151
R1229 B.n255 B.n212 10.6151
R1230 B.n255 B.n254 10.6151
R1231 B.n254 B.n253 10.6151
R1232 B.n253 B.n214 10.6151
R1233 B.n249 B.n214 10.6151
R1234 B.n249 B.n248 10.6151
R1235 B.n248 B.n247 10.6151
R1236 B.n247 B.n216 10.6151
R1237 B.n243 B.n216 10.6151
R1238 B.n243 B.n242 10.6151
R1239 B.n242 B.n241 10.6151
R1240 B.n241 B.n218 10.6151
R1241 B.n237 B.n218 10.6151
R1242 B.n237 B.n236 10.6151
R1243 B.n236 B.n235 10.6151
R1244 B.n235 B.n220 10.6151
R1245 B.n231 B.n220 10.6151
R1246 B.n231 B.n230 10.6151
R1247 B.n230 B.n229 10.6151
R1248 B.n229 B.n222 10.6151
R1249 B.n225 B.n222 10.6151
R1250 B.n225 B.n224 10.6151
R1251 B.n224 B.n0 10.6151
R1252 B.n863 B.n1 10.6151
R1253 B.n863 B.n862 10.6151
R1254 B.n862 B.n861 10.6151
R1255 B.n861 B.n4 10.6151
R1256 B.n857 B.n4 10.6151
R1257 B.n857 B.n856 10.6151
R1258 B.n856 B.n855 10.6151
R1259 B.n855 B.n6 10.6151
R1260 B.n851 B.n6 10.6151
R1261 B.n851 B.n850 10.6151
R1262 B.n850 B.n849 10.6151
R1263 B.n849 B.n8 10.6151
R1264 B.n845 B.n8 10.6151
R1265 B.n845 B.n844 10.6151
R1266 B.n844 B.n843 10.6151
R1267 B.n843 B.n10 10.6151
R1268 B.n839 B.n10 10.6151
R1269 B.n839 B.n838 10.6151
R1270 B.n838 B.n837 10.6151
R1271 B.n837 B.n12 10.6151
R1272 B.n833 B.n12 10.6151
R1273 B.n833 B.n832 10.6151
R1274 B.n832 B.n831 10.6151
R1275 B.n831 B.n14 10.6151
R1276 B.n827 B.n14 10.6151
R1277 B.n827 B.n826 10.6151
R1278 B.n826 B.n825 10.6151
R1279 B.n825 B.n16 10.6151
R1280 B.n821 B.n16 10.6151
R1281 B.n821 B.n820 10.6151
R1282 B.n820 B.n819 10.6151
R1283 B.n819 B.n18 10.6151
R1284 B.n815 B.n18 10.6151
R1285 B.n815 B.n814 10.6151
R1286 B.n814 B.n813 10.6151
R1287 B.n813 B.n20 10.6151
R1288 B.n809 B.n20 10.6151
R1289 B.n809 B.n808 10.6151
R1290 B.n808 B.n807 10.6151
R1291 B.n807 B.n22 10.6151
R1292 B.n803 B.n22 10.6151
R1293 B.n803 B.n802 10.6151
R1294 B.n802 B.n801 10.6151
R1295 B.n801 B.n24 10.6151
R1296 B.n797 B.n24 10.6151
R1297 B.n797 B.n796 10.6151
R1298 B.n796 B.n795 10.6151
R1299 B.n712 B.n711 6.5566
R1300 B.n699 B.n698 6.5566
R1301 B.n376 B.n375 6.5566
R1302 B.n388 B.n166 6.5566
R1303 B.n713 B.n712 4.05904
R1304 B.n698 B.n697 4.05904
R1305 B.n375 B.n374 4.05904
R1306 B.n391 B.n166 4.05904
R1307 B.n867 B.n0 2.81026
R1308 B.n867 B.n1 2.81026
R1309 VP.n18 VP.t0 233.626
R1310 VP.n60 VP.t1 200.751
R1311 VP.n44 VP.t8 200.751
R1312 VP.n7 VP.t5 200.751
R1313 VP.n67 VP.t9 200.751
R1314 VP.n75 VP.t6 200.751
R1315 VP.n26 VP.t4 200.751
R1316 VP.n41 VP.t2 200.751
R1317 VP.n33 VP.t7 200.751
R1318 VP.n17 VP.t3 200.751
R1319 VP.n44 VP.n43 183.924
R1320 VP.n76 VP.n75 183.924
R1321 VP.n42 VP.n41 183.924
R1322 VP.n20 VP.n19 161.3
R1323 VP.n21 VP.n16 161.3
R1324 VP.n23 VP.n22 161.3
R1325 VP.n24 VP.n15 161.3
R1326 VP.n26 VP.n25 161.3
R1327 VP.n27 VP.n14 161.3
R1328 VP.n29 VP.n28 161.3
R1329 VP.n30 VP.n13 161.3
R1330 VP.n32 VP.n31 161.3
R1331 VP.n34 VP.n12 161.3
R1332 VP.n36 VP.n35 161.3
R1333 VP.n37 VP.n11 161.3
R1334 VP.n39 VP.n38 161.3
R1335 VP.n40 VP.n10 161.3
R1336 VP.n74 VP.n0 161.3
R1337 VP.n73 VP.n72 161.3
R1338 VP.n71 VP.n1 161.3
R1339 VP.n70 VP.n69 161.3
R1340 VP.n68 VP.n2 161.3
R1341 VP.n66 VP.n65 161.3
R1342 VP.n64 VP.n3 161.3
R1343 VP.n63 VP.n62 161.3
R1344 VP.n61 VP.n4 161.3
R1345 VP.n60 VP.n59 161.3
R1346 VP.n58 VP.n5 161.3
R1347 VP.n57 VP.n56 161.3
R1348 VP.n55 VP.n6 161.3
R1349 VP.n54 VP.n53 161.3
R1350 VP.n52 VP.n51 161.3
R1351 VP.n50 VP.n8 161.3
R1352 VP.n49 VP.n48 161.3
R1353 VP.n47 VP.n9 161.3
R1354 VP.n46 VP.n45 161.3
R1355 VP.n18 VP.n17 56.9995
R1356 VP.n56 VP.n55 53.6554
R1357 VP.n62 VP.n3 53.6554
R1358 VP.n28 VP.n13 53.6554
R1359 VP.n22 VP.n21 53.6554
R1360 VP.n43 VP.n42 52.5876
R1361 VP.n50 VP.n49 49.7803
R1362 VP.n69 VP.n1 49.7803
R1363 VP.n35 VP.n11 49.7803
R1364 VP.n49 VP.n9 31.3737
R1365 VP.n73 VP.n1 31.3737
R1366 VP.n39 VP.n11 31.3737
R1367 VP.n56 VP.n5 27.4986
R1368 VP.n62 VP.n61 27.4986
R1369 VP.n28 VP.n27 27.4986
R1370 VP.n22 VP.n15 27.4986
R1371 VP.n45 VP.n9 24.5923
R1372 VP.n51 VP.n50 24.5923
R1373 VP.n55 VP.n54 24.5923
R1374 VP.n60 VP.n5 24.5923
R1375 VP.n61 VP.n60 24.5923
R1376 VP.n66 VP.n3 24.5923
R1377 VP.n69 VP.n68 24.5923
R1378 VP.n74 VP.n73 24.5923
R1379 VP.n40 VP.n39 24.5923
R1380 VP.n32 VP.n13 24.5923
R1381 VP.n35 VP.n34 24.5923
R1382 VP.n26 VP.n15 24.5923
R1383 VP.n27 VP.n26 24.5923
R1384 VP.n21 VP.n20 24.5923
R1385 VP.n54 VP.n7 13.2801
R1386 VP.n67 VP.n66 13.2801
R1387 VP.n33 VP.n32 13.2801
R1388 VP.n20 VP.n17 13.2801
R1389 VP.n19 VP.n18 12.447
R1390 VP.n51 VP.n7 11.3127
R1391 VP.n68 VP.n67 11.3127
R1392 VP.n34 VP.n33 11.3127
R1393 VP.n45 VP.n44 1.96785
R1394 VP.n75 VP.n74 1.96785
R1395 VP.n41 VP.n40 1.96785
R1396 VP.n19 VP.n16 0.189894
R1397 VP.n23 VP.n16 0.189894
R1398 VP.n24 VP.n23 0.189894
R1399 VP.n25 VP.n24 0.189894
R1400 VP.n25 VP.n14 0.189894
R1401 VP.n29 VP.n14 0.189894
R1402 VP.n30 VP.n29 0.189894
R1403 VP.n31 VP.n30 0.189894
R1404 VP.n31 VP.n12 0.189894
R1405 VP.n36 VP.n12 0.189894
R1406 VP.n37 VP.n36 0.189894
R1407 VP.n38 VP.n37 0.189894
R1408 VP.n38 VP.n10 0.189894
R1409 VP.n42 VP.n10 0.189894
R1410 VP.n46 VP.n43 0.189894
R1411 VP.n47 VP.n46 0.189894
R1412 VP.n48 VP.n47 0.189894
R1413 VP.n48 VP.n8 0.189894
R1414 VP.n52 VP.n8 0.189894
R1415 VP.n53 VP.n52 0.189894
R1416 VP.n53 VP.n6 0.189894
R1417 VP.n57 VP.n6 0.189894
R1418 VP.n58 VP.n57 0.189894
R1419 VP.n59 VP.n58 0.189894
R1420 VP.n59 VP.n4 0.189894
R1421 VP.n63 VP.n4 0.189894
R1422 VP.n64 VP.n63 0.189894
R1423 VP.n65 VP.n64 0.189894
R1424 VP.n65 VP.n2 0.189894
R1425 VP.n70 VP.n2 0.189894
R1426 VP.n71 VP.n70 0.189894
R1427 VP.n72 VP.n71 0.189894
R1428 VP.n72 VP.n0 0.189894
R1429 VP.n76 VP.n0 0.189894
R1430 VP VP.n76 0.0516364
R1431 VTAIL.n368 VTAIL.n284 756.745
R1432 VTAIL.n86 VTAIL.n2 756.745
R1433 VTAIL.n278 VTAIL.n194 756.745
R1434 VTAIL.n184 VTAIL.n100 756.745
R1435 VTAIL.n312 VTAIL.n311 585
R1436 VTAIL.n317 VTAIL.n316 585
R1437 VTAIL.n319 VTAIL.n318 585
R1438 VTAIL.n308 VTAIL.n307 585
R1439 VTAIL.n325 VTAIL.n324 585
R1440 VTAIL.n327 VTAIL.n326 585
R1441 VTAIL.n304 VTAIL.n303 585
R1442 VTAIL.n333 VTAIL.n332 585
R1443 VTAIL.n335 VTAIL.n334 585
R1444 VTAIL.n300 VTAIL.n299 585
R1445 VTAIL.n341 VTAIL.n340 585
R1446 VTAIL.n343 VTAIL.n342 585
R1447 VTAIL.n296 VTAIL.n295 585
R1448 VTAIL.n349 VTAIL.n348 585
R1449 VTAIL.n351 VTAIL.n350 585
R1450 VTAIL.n292 VTAIL.n291 585
R1451 VTAIL.n358 VTAIL.n357 585
R1452 VTAIL.n359 VTAIL.n290 585
R1453 VTAIL.n361 VTAIL.n360 585
R1454 VTAIL.n288 VTAIL.n287 585
R1455 VTAIL.n367 VTAIL.n366 585
R1456 VTAIL.n369 VTAIL.n368 585
R1457 VTAIL.n30 VTAIL.n29 585
R1458 VTAIL.n35 VTAIL.n34 585
R1459 VTAIL.n37 VTAIL.n36 585
R1460 VTAIL.n26 VTAIL.n25 585
R1461 VTAIL.n43 VTAIL.n42 585
R1462 VTAIL.n45 VTAIL.n44 585
R1463 VTAIL.n22 VTAIL.n21 585
R1464 VTAIL.n51 VTAIL.n50 585
R1465 VTAIL.n53 VTAIL.n52 585
R1466 VTAIL.n18 VTAIL.n17 585
R1467 VTAIL.n59 VTAIL.n58 585
R1468 VTAIL.n61 VTAIL.n60 585
R1469 VTAIL.n14 VTAIL.n13 585
R1470 VTAIL.n67 VTAIL.n66 585
R1471 VTAIL.n69 VTAIL.n68 585
R1472 VTAIL.n10 VTAIL.n9 585
R1473 VTAIL.n76 VTAIL.n75 585
R1474 VTAIL.n77 VTAIL.n8 585
R1475 VTAIL.n79 VTAIL.n78 585
R1476 VTAIL.n6 VTAIL.n5 585
R1477 VTAIL.n85 VTAIL.n84 585
R1478 VTAIL.n87 VTAIL.n86 585
R1479 VTAIL.n279 VTAIL.n278 585
R1480 VTAIL.n277 VTAIL.n276 585
R1481 VTAIL.n198 VTAIL.n197 585
R1482 VTAIL.n271 VTAIL.n270 585
R1483 VTAIL.n269 VTAIL.n200 585
R1484 VTAIL.n268 VTAIL.n267 585
R1485 VTAIL.n203 VTAIL.n201 585
R1486 VTAIL.n262 VTAIL.n261 585
R1487 VTAIL.n260 VTAIL.n259 585
R1488 VTAIL.n207 VTAIL.n206 585
R1489 VTAIL.n254 VTAIL.n253 585
R1490 VTAIL.n252 VTAIL.n251 585
R1491 VTAIL.n211 VTAIL.n210 585
R1492 VTAIL.n246 VTAIL.n245 585
R1493 VTAIL.n244 VTAIL.n243 585
R1494 VTAIL.n215 VTAIL.n214 585
R1495 VTAIL.n238 VTAIL.n237 585
R1496 VTAIL.n236 VTAIL.n235 585
R1497 VTAIL.n219 VTAIL.n218 585
R1498 VTAIL.n230 VTAIL.n229 585
R1499 VTAIL.n228 VTAIL.n227 585
R1500 VTAIL.n223 VTAIL.n222 585
R1501 VTAIL.n185 VTAIL.n184 585
R1502 VTAIL.n183 VTAIL.n182 585
R1503 VTAIL.n104 VTAIL.n103 585
R1504 VTAIL.n177 VTAIL.n176 585
R1505 VTAIL.n175 VTAIL.n106 585
R1506 VTAIL.n174 VTAIL.n173 585
R1507 VTAIL.n109 VTAIL.n107 585
R1508 VTAIL.n168 VTAIL.n167 585
R1509 VTAIL.n166 VTAIL.n165 585
R1510 VTAIL.n113 VTAIL.n112 585
R1511 VTAIL.n160 VTAIL.n159 585
R1512 VTAIL.n158 VTAIL.n157 585
R1513 VTAIL.n117 VTAIL.n116 585
R1514 VTAIL.n152 VTAIL.n151 585
R1515 VTAIL.n150 VTAIL.n149 585
R1516 VTAIL.n121 VTAIL.n120 585
R1517 VTAIL.n144 VTAIL.n143 585
R1518 VTAIL.n142 VTAIL.n141 585
R1519 VTAIL.n125 VTAIL.n124 585
R1520 VTAIL.n136 VTAIL.n135 585
R1521 VTAIL.n134 VTAIL.n133 585
R1522 VTAIL.n129 VTAIL.n128 585
R1523 VTAIL.n313 VTAIL.t8 327.466
R1524 VTAIL.n31 VTAIL.t11 327.466
R1525 VTAIL.n224 VTAIL.t12 327.466
R1526 VTAIL.n130 VTAIL.t0 327.466
R1527 VTAIL.n317 VTAIL.n311 171.744
R1528 VTAIL.n318 VTAIL.n317 171.744
R1529 VTAIL.n318 VTAIL.n307 171.744
R1530 VTAIL.n325 VTAIL.n307 171.744
R1531 VTAIL.n326 VTAIL.n325 171.744
R1532 VTAIL.n326 VTAIL.n303 171.744
R1533 VTAIL.n333 VTAIL.n303 171.744
R1534 VTAIL.n334 VTAIL.n333 171.744
R1535 VTAIL.n334 VTAIL.n299 171.744
R1536 VTAIL.n341 VTAIL.n299 171.744
R1537 VTAIL.n342 VTAIL.n341 171.744
R1538 VTAIL.n342 VTAIL.n295 171.744
R1539 VTAIL.n349 VTAIL.n295 171.744
R1540 VTAIL.n350 VTAIL.n349 171.744
R1541 VTAIL.n350 VTAIL.n291 171.744
R1542 VTAIL.n358 VTAIL.n291 171.744
R1543 VTAIL.n359 VTAIL.n358 171.744
R1544 VTAIL.n360 VTAIL.n359 171.744
R1545 VTAIL.n360 VTAIL.n287 171.744
R1546 VTAIL.n367 VTAIL.n287 171.744
R1547 VTAIL.n368 VTAIL.n367 171.744
R1548 VTAIL.n35 VTAIL.n29 171.744
R1549 VTAIL.n36 VTAIL.n35 171.744
R1550 VTAIL.n36 VTAIL.n25 171.744
R1551 VTAIL.n43 VTAIL.n25 171.744
R1552 VTAIL.n44 VTAIL.n43 171.744
R1553 VTAIL.n44 VTAIL.n21 171.744
R1554 VTAIL.n51 VTAIL.n21 171.744
R1555 VTAIL.n52 VTAIL.n51 171.744
R1556 VTAIL.n52 VTAIL.n17 171.744
R1557 VTAIL.n59 VTAIL.n17 171.744
R1558 VTAIL.n60 VTAIL.n59 171.744
R1559 VTAIL.n60 VTAIL.n13 171.744
R1560 VTAIL.n67 VTAIL.n13 171.744
R1561 VTAIL.n68 VTAIL.n67 171.744
R1562 VTAIL.n68 VTAIL.n9 171.744
R1563 VTAIL.n76 VTAIL.n9 171.744
R1564 VTAIL.n77 VTAIL.n76 171.744
R1565 VTAIL.n78 VTAIL.n77 171.744
R1566 VTAIL.n78 VTAIL.n5 171.744
R1567 VTAIL.n85 VTAIL.n5 171.744
R1568 VTAIL.n86 VTAIL.n85 171.744
R1569 VTAIL.n278 VTAIL.n277 171.744
R1570 VTAIL.n277 VTAIL.n197 171.744
R1571 VTAIL.n270 VTAIL.n197 171.744
R1572 VTAIL.n270 VTAIL.n269 171.744
R1573 VTAIL.n269 VTAIL.n268 171.744
R1574 VTAIL.n268 VTAIL.n201 171.744
R1575 VTAIL.n261 VTAIL.n201 171.744
R1576 VTAIL.n261 VTAIL.n260 171.744
R1577 VTAIL.n260 VTAIL.n206 171.744
R1578 VTAIL.n253 VTAIL.n206 171.744
R1579 VTAIL.n253 VTAIL.n252 171.744
R1580 VTAIL.n252 VTAIL.n210 171.744
R1581 VTAIL.n245 VTAIL.n210 171.744
R1582 VTAIL.n245 VTAIL.n244 171.744
R1583 VTAIL.n244 VTAIL.n214 171.744
R1584 VTAIL.n237 VTAIL.n214 171.744
R1585 VTAIL.n237 VTAIL.n236 171.744
R1586 VTAIL.n236 VTAIL.n218 171.744
R1587 VTAIL.n229 VTAIL.n218 171.744
R1588 VTAIL.n229 VTAIL.n228 171.744
R1589 VTAIL.n228 VTAIL.n222 171.744
R1590 VTAIL.n184 VTAIL.n183 171.744
R1591 VTAIL.n183 VTAIL.n103 171.744
R1592 VTAIL.n176 VTAIL.n103 171.744
R1593 VTAIL.n176 VTAIL.n175 171.744
R1594 VTAIL.n175 VTAIL.n174 171.744
R1595 VTAIL.n174 VTAIL.n107 171.744
R1596 VTAIL.n167 VTAIL.n107 171.744
R1597 VTAIL.n167 VTAIL.n166 171.744
R1598 VTAIL.n166 VTAIL.n112 171.744
R1599 VTAIL.n159 VTAIL.n112 171.744
R1600 VTAIL.n159 VTAIL.n158 171.744
R1601 VTAIL.n158 VTAIL.n116 171.744
R1602 VTAIL.n151 VTAIL.n116 171.744
R1603 VTAIL.n151 VTAIL.n150 171.744
R1604 VTAIL.n150 VTAIL.n120 171.744
R1605 VTAIL.n143 VTAIL.n120 171.744
R1606 VTAIL.n143 VTAIL.n142 171.744
R1607 VTAIL.n142 VTAIL.n124 171.744
R1608 VTAIL.n135 VTAIL.n124 171.744
R1609 VTAIL.n135 VTAIL.n134 171.744
R1610 VTAIL.n134 VTAIL.n128 171.744
R1611 VTAIL.t8 VTAIL.n311 85.8723
R1612 VTAIL.t11 VTAIL.n29 85.8723
R1613 VTAIL.t12 VTAIL.n222 85.8723
R1614 VTAIL.t0 VTAIL.n128 85.8723
R1615 VTAIL.n193 VTAIL.n192 54.6749
R1616 VTAIL.n191 VTAIL.n190 54.6749
R1617 VTAIL.n99 VTAIL.n98 54.6749
R1618 VTAIL.n97 VTAIL.n96 54.6749
R1619 VTAIL.n375 VTAIL.n374 54.6747
R1620 VTAIL.n1 VTAIL.n0 54.6747
R1621 VTAIL.n93 VTAIL.n92 54.6747
R1622 VTAIL.n95 VTAIL.n94 54.6747
R1623 VTAIL.n373 VTAIL.n372 33.7369
R1624 VTAIL.n91 VTAIL.n90 33.7369
R1625 VTAIL.n283 VTAIL.n282 33.7369
R1626 VTAIL.n189 VTAIL.n188 33.7369
R1627 VTAIL.n97 VTAIL.n95 30.2117
R1628 VTAIL.n373 VTAIL.n283 28.2548
R1629 VTAIL.n313 VTAIL.n312 16.3895
R1630 VTAIL.n31 VTAIL.n30 16.3895
R1631 VTAIL.n224 VTAIL.n223 16.3895
R1632 VTAIL.n130 VTAIL.n129 16.3895
R1633 VTAIL.n361 VTAIL.n290 13.1884
R1634 VTAIL.n79 VTAIL.n8 13.1884
R1635 VTAIL.n271 VTAIL.n200 13.1884
R1636 VTAIL.n177 VTAIL.n106 13.1884
R1637 VTAIL.n316 VTAIL.n315 12.8005
R1638 VTAIL.n357 VTAIL.n356 12.8005
R1639 VTAIL.n362 VTAIL.n288 12.8005
R1640 VTAIL.n34 VTAIL.n33 12.8005
R1641 VTAIL.n75 VTAIL.n74 12.8005
R1642 VTAIL.n80 VTAIL.n6 12.8005
R1643 VTAIL.n272 VTAIL.n198 12.8005
R1644 VTAIL.n267 VTAIL.n202 12.8005
R1645 VTAIL.n227 VTAIL.n226 12.8005
R1646 VTAIL.n178 VTAIL.n104 12.8005
R1647 VTAIL.n173 VTAIL.n108 12.8005
R1648 VTAIL.n133 VTAIL.n132 12.8005
R1649 VTAIL.n319 VTAIL.n310 12.0247
R1650 VTAIL.n355 VTAIL.n292 12.0247
R1651 VTAIL.n366 VTAIL.n365 12.0247
R1652 VTAIL.n37 VTAIL.n28 12.0247
R1653 VTAIL.n73 VTAIL.n10 12.0247
R1654 VTAIL.n84 VTAIL.n83 12.0247
R1655 VTAIL.n276 VTAIL.n275 12.0247
R1656 VTAIL.n266 VTAIL.n203 12.0247
R1657 VTAIL.n230 VTAIL.n221 12.0247
R1658 VTAIL.n182 VTAIL.n181 12.0247
R1659 VTAIL.n172 VTAIL.n109 12.0247
R1660 VTAIL.n136 VTAIL.n127 12.0247
R1661 VTAIL.n320 VTAIL.n308 11.249
R1662 VTAIL.n352 VTAIL.n351 11.249
R1663 VTAIL.n369 VTAIL.n286 11.249
R1664 VTAIL.n38 VTAIL.n26 11.249
R1665 VTAIL.n70 VTAIL.n69 11.249
R1666 VTAIL.n87 VTAIL.n4 11.249
R1667 VTAIL.n279 VTAIL.n196 11.249
R1668 VTAIL.n263 VTAIL.n262 11.249
R1669 VTAIL.n231 VTAIL.n219 11.249
R1670 VTAIL.n185 VTAIL.n102 11.249
R1671 VTAIL.n169 VTAIL.n168 11.249
R1672 VTAIL.n137 VTAIL.n125 11.249
R1673 VTAIL.n324 VTAIL.n323 10.4732
R1674 VTAIL.n348 VTAIL.n294 10.4732
R1675 VTAIL.n370 VTAIL.n284 10.4732
R1676 VTAIL.n42 VTAIL.n41 10.4732
R1677 VTAIL.n66 VTAIL.n12 10.4732
R1678 VTAIL.n88 VTAIL.n2 10.4732
R1679 VTAIL.n280 VTAIL.n194 10.4732
R1680 VTAIL.n259 VTAIL.n205 10.4732
R1681 VTAIL.n235 VTAIL.n234 10.4732
R1682 VTAIL.n186 VTAIL.n100 10.4732
R1683 VTAIL.n165 VTAIL.n111 10.4732
R1684 VTAIL.n141 VTAIL.n140 10.4732
R1685 VTAIL.n327 VTAIL.n306 9.69747
R1686 VTAIL.n347 VTAIL.n296 9.69747
R1687 VTAIL.n45 VTAIL.n24 9.69747
R1688 VTAIL.n65 VTAIL.n14 9.69747
R1689 VTAIL.n258 VTAIL.n207 9.69747
R1690 VTAIL.n238 VTAIL.n217 9.69747
R1691 VTAIL.n164 VTAIL.n113 9.69747
R1692 VTAIL.n144 VTAIL.n123 9.69747
R1693 VTAIL.n372 VTAIL.n371 9.45567
R1694 VTAIL.n90 VTAIL.n89 9.45567
R1695 VTAIL.n282 VTAIL.n281 9.45567
R1696 VTAIL.n188 VTAIL.n187 9.45567
R1697 VTAIL.n371 VTAIL.n370 9.3005
R1698 VTAIL.n286 VTAIL.n285 9.3005
R1699 VTAIL.n365 VTAIL.n364 9.3005
R1700 VTAIL.n363 VTAIL.n362 9.3005
R1701 VTAIL.n302 VTAIL.n301 9.3005
R1702 VTAIL.n331 VTAIL.n330 9.3005
R1703 VTAIL.n329 VTAIL.n328 9.3005
R1704 VTAIL.n306 VTAIL.n305 9.3005
R1705 VTAIL.n323 VTAIL.n322 9.3005
R1706 VTAIL.n321 VTAIL.n320 9.3005
R1707 VTAIL.n310 VTAIL.n309 9.3005
R1708 VTAIL.n315 VTAIL.n314 9.3005
R1709 VTAIL.n337 VTAIL.n336 9.3005
R1710 VTAIL.n339 VTAIL.n338 9.3005
R1711 VTAIL.n298 VTAIL.n297 9.3005
R1712 VTAIL.n345 VTAIL.n344 9.3005
R1713 VTAIL.n347 VTAIL.n346 9.3005
R1714 VTAIL.n294 VTAIL.n293 9.3005
R1715 VTAIL.n353 VTAIL.n352 9.3005
R1716 VTAIL.n355 VTAIL.n354 9.3005
R1717 VTAIL.n356 VTAIL.n289 9.3005
R1718 VTAIL.n89 VTAIL.n88 9.3005
R1719 VTAIL.n4 VTAIL.n3 9.3005
R1720 VTAIL.n83 VTAIL.n82 9.3005
R1721 VTAIL.n81 VTAIL.n80 9.3005
R1722 VTAIL.n20 VTAIL.n19 9.3005
R1723 VTAIL.n49 VTAIL.n48 9.3005
R1724 VTAIL.n47 VTAIL.n46 9.3005
R1725 VTAIL.n24 VTAIL.n23 9.3005
R1726 VTAIL.n41 VTAIL.n40 9.3005
R1727 VTAIL.n39 VTAIL.n38 9.3005
R1728 VTAIL.n28 VTAIL.n27 9.3005
R1729 VTAIL.n33 VTAIL.n32 9.3005
R1730 VTAIL.n55 VTAIL.n54 9.3005
R1731 VTAIL.n57 VTAIL.n56 9.3005
R1732 VTAIL.n16 VTAIL.n15 9.3005
R1733 VTAIL.n63 VTAIL.n62 9.3005
R1734 VTAIL.n65 VTAIL.n64 9.3005
R1735 VTAIL.n12 VTAIL.n11 9.3005
R1736 VTAIL.n71 VTAIL.n70 9.3005
R1737 VTAIL.n73 VTAIL.n72 9.3005
R1738 VTAIL.n74 VTAIL.n7 9.3005
R1739 VTAIL.n250 VTAIL.n249 9.3005
R1740 VTAIL.n209 VTAIL.n208 9.3005
R1741 VTAIL.n256 VTAIL.n255 9.3005
R1742 VTAIL.n258 VTAIL.n257 9.3005
R1743 VTAIL.n205 VTAIL.n204 9.3005
R1744 VTAIL.n264 VTAIL.n263 9.3005
R1745 VTAIL.n266 VTAIL.n265 9.3005
R1746 VTAIL.n202 VTAIL.n199 9.3005
R1747 VTAIL.n281 VTAIL.n280 9.3005
R1748 VTAIL.n196 VTAIL.n195 9.3005
R1749 VTAIL.n275 VTAIL.n274 9.3005
R1750 VTAIL.n273 VTAIL.n272 9.3005
R1751 VTAIL.n248 VTAIL.n247 9.3005
R1752 VTAIL.n213 VTAIL.n212 9.3005
R1753 VTAIL.n242 VTAIL.n241 9.3005
R1754 VTAIL.n240 VTAIL.n239 9.3005
R1755 VTAIL.n217 VTAIL.n216 9.3005
R1756 VTAIL.n234 VTAIL.n233 9.3005
R1757 VTAIL.n232 VTAIL.n231 9.3005
R1758 VTAIL.n221 VTAIL.n220 9.3005
R1759 VTAIL.n226 VTAIL.n225 9.3005
R1760 VTAIL.n156 VTAIL.n155 9.3005
R1761 VTAIL.n115 VTAIL.n114 9.3005
R1762 VTAIL.n162 VTAIL.n161 9.3005
R1763 VTAIL.n164 VTAIL.n163 9.3005
R1764 VTAIL.n111 VTAIL.n110 9.3005
R1765 VTAIL.n170 VTAIL.n169 9.3005
R1766 VTAIL.n172 VTAIL.n171 9.3005
R1767 VTAIL.n108 VTAIL.n105 9.3005
R1768 VTAIL.n187 VTAIL.n186 9.3005
R1769 VTAIL.n102 VTAIL.n101 9.3005
R1770 VTAIL.n181 VTAIL.n180 9.3005
R1771 VTAIL.n179 VTAIL.n178 9.3005
R1772 VTAIL.n154 VTAIL.n153 9.3005
R1773 VTAIL.n119 VTAIL.n118 9.3005
R1774 VTAIL.n148 VTAIL.n147 9.3005
R1775 VTAIL.n146 VTAIL.n145 9.3005
R1776 VTAIL.n123 VTAIL.n122 9.3005
R1777 VTAIL.n140 VTAIL.n139 9.3005
R1778 VTAIL.n138 VTAIL.n137 9.3005
R1779 VTAIL.n127 VTAIL.n126 9.3005
R1780 VTAIL.n132 VTAIL.n131 9.3005
R1781 VTAIL.n328 VTAIL.n304 8.92171
R1782 VTAIL.n344 VTAIL.n343 8.92171
R1783 VTAIL.n46 VTAIL.n22 8.92171
R1784 VTAIL.n62 VTAIL.n61 8.92171
R1785 VTAIL.n255 VTAIL.n254 8.92171
R1786 VTAIL.n239 VTAIL.n215 8.92171
R1787 VTAIL.n161 VTAIL.n160 8.92171
R1788 VTAIL.n145 VTAIL.n121 8.92171
R1789 VTAIL.n332 VTAIL.n331 8.14595
R1790 VTAIL.n340 VTAIL.n298 8.14595
R1791 VTAIL.n50 VTAIL.n49 8.14595
R1792 VTAIL.n58 VTAIL.n16 8.14595
R1793 VTAIL.n251 VTAIL.n209 8.14595
R1794 VTAIL.n243 VTAIL.n242 8.14595
R1795 VTAIL.n157 VTAIL.n115 8.14595
R1796 VTAIL.n149 VTAIL.n148 8.14595
R1797 VTAIL.n335 VTAIL.n302 7.3702
R1798 VTAIL.n339 VTAIL.n300 7.3702
R1799 VTAIL.n53 VTAIL.n20 7.3702
R1800 VTAIL.n57 VTAIL.n18 7.3702
R1801 VTAIL.n250 VTAIL.n211 7.3702
R1802 VTAIL.n246 VTAIL.n213 7.3702
R1803 VTAIL.n156 VTAIL.n117 7.3702
R1804 VTAIL.n152 VTAIL.n119 7.3702
R1805 VTAIL.n336 VTAIL.n335 6.59444
R1806 VTAIL.n336 VTAIL.n300 6.59444
R1807 VTAIL.n54 VTAIL.n53 6.59444
R1808 VTAIL.n54 VTAIL.n18 6.59444
R1809 VTAIL.n247 VTAIL.n211 6.59444
R1810 VTAIL.n247 VTAIL.n246 6.59444
R1811 VTAIL.n153 VTAIL.n117 6.59444
R1812 VTAIL.n153 VTAIL.n152 6.59444
R1813 VTAIL.n332 VTAIL.n302 5.81868
R1814 VTAIL.n340 VTAIL.n339 5.81868
R1815 VTAIL.n50 VTAIL.n20 5.81868
R1816 VTAIL.n58 VTAIL.n57 5.81868
R1817 VTAIL.n251 VTAIL.n250 5.81868
R1818 VTAIL.n243 VTAIL.n213 5.81868
R1819 VTAIL.n157 VTAIL.n156 5.81868
R1820 VTAIL.n149 VTAIL.n119 5.81868
R1821 VTAIL.n331 VTAIL.n304 5.04292
R1822 VTAIL.n343 VTAIL.n298 5.04292
R1823 VTAIL.n49 VTAIL.n22 5.04292
R1824 VTAIL.n61 VTAIL.n16 5.04292
R1825 VTAIL.n254 VTAIL.n209 5.04292
R1826 VTAIL.n242 VTAIL.n215 5.04292
R1827 VTAIL.n160 VTAIL.n115 5.04292
R1828 VTAIL.n148 VTAIL.n121 5.04292
R1829 VTAIL.n328 VTAIL.n327 4.26717
R1830 VTAIL.n344 VTAIL.n296 4.26717
R1831 VTAIL.n46 VTAIL.n45 4.26717
R1832 VTAIL.n62 VTAIL.n14 4.26717
R1833 VTAIL.n255 VTAIL.n207 4.26717
R1834 VTAIL.n239 VTAIL.n238 4.26717
R1835 VTAIL.n161 VTAIL.n113 4.26717
R1836 VTAIL.n145 VTAIL.n144 4.26717
R1837 VTAIL.n314 VTAIL.n313 3.70982
R1838 VTAIL.n32 VTAIL.n31 3.70982
R1839 VTAIL.n225 VTAIL.n224 3.70982
R1840 VTAIL.n131 VTAIL.n130 3.70982
R1841 VTAIL.n324 VTAIL.n306 3.49141
R1842 VTAIL.n348 VTAIL.n347 3.49141
R1843 VTAIL.n372 VTAIL.n284 3.49141
R1844 VTAIL.n42 VTAIL.n24 3.49141
R1845 VTAIL.n66 VTAIL.n65 3.49141
R1846 VTAIL.n90 VTAIL.n2 3.49141
R1847 VTAIL.n282 VTAIL.n194 3.49141
R1848 VTAIL.n259 VTAIL.n258 3.49141
R1849 VTAIL.n235 VTAIL.n217 3.49141
R1850 VTAIL.n188 VTAIL.n100 3.49141
R1851 VTAIL.n165 VTAIL.n164 3.49141
R1852 VTAIL.n141 VTAIL.n123 3.49141
R1853 VTAIL.n323 VTAIL.n308 2.71565
R1854 VTAIL.n351 VTAIL.n294 2.71565
R1855 VTAIL.n370 VTAIL.n369 2.71565
R1856 VTAIL.n41 VTAIL.n26 2.71565
R1857 VTAIL.n69 VTAIL.n12 2.71565
R1858 VTAIL.n88 VTAIL.n87 2.71565
R1859 VTAIL.n280 VTAIL.n279 2.71565
R1860 VTAIL.n262 VTAIL.n205 2.71565
R1861 VTAIL.n234 VTAIL.n219 2.71565
R1862 VTAIL.n186 VTAIL.n185 2.71565
R1863 VTAIL.n168 VTAIL.n111 2.71565
R1864 VTAIL.n140 VTAIL.n125 2.71565
R1865 VTAIL.n374 VTAIL.t7 2.01195
R1866 VTAIL.n374 VTAIL.t6 2.01195
R1867 VTAIL.n0 VTAIL.t19 2.01195
R1868 VTAIL.n0 VTAIL.t5 2.01195
R1869 VTAIL.n92 VTAIL.t17 2.01195
R1870 VTAIL.n92 VTAIL.t16 2.01195
R1871 VTAIL.n94 VTAIL.t14 2.01195
R1872 VTAIL.n94 VTAIL.t10 2.01195
R1873 VTAIL.n192 VTAIL.t13 2.01195
R1874 VTAIL.n192 VTAIL.t15 2.01195
R1875 VTAIL.n190 VTAIL.t18 2.01195
R1876 VTAIL.n190 VTAIL.t9 2.01195
R1877 VTAIL.n98 VTAIL.t3 2.01195
R1878 VTAIL.n98 VTAIL.t4 2.01195
R1879 VTAIL.n96 VTAIL.t2 2.01195
R1880 VTAIL.n96 VTAIL.t1 2.01195
R1881 VTAIL.n99 VTAIL.n97 1.9574
R1882 VTAIL.n189 VTAIL.n99 1.9574
R1883 VTAIL.n193 VTAIL.n191 1.9574
R1884 VTAIL.n283 VTAIL.n193 1.9574
R1885 VTAIL.n95 VTAIL.n93 1.9574
R1886 VTAIL.n93 VTAIL.n91 1.9574
R1887 VTAIL.n375 VTAIL.n373 1.9574
R1888 VTAIL.n320 VTAIL.n319 1.93989
R1889 VTAIL.n352 VTAIL.n292 1.93989
R1890 VTAIL.n366 VTAIL.n286 1.93989
R1891 VTAIL.n38 VTAIL.n37 1.93989
R1892 VTAIL.n70 VTAIL.n10 1.93989
R1893 VTAIL.n84 VTAIL.n4 1.93989
R1894 VTAIL.n276 VTAIL.n196 1.93989
R1895 VTAIL.n263 VTAIL.n203 1.93989
R1896 VTAIL.n231 VTAIL.n230 1.93989
R1897 VTAIL.n182 VTAIL.n102 1.93989
R1898 VTAIL.n169 VTAIL.n109 1.93989
R1899 VTAIL.n137 VTAIL.n136 1.93989
R1900 VTAIL VTAIL.n1 1.52636
R1901 VTAIL.n191 VTAIL.n189 1.44878
R1902 VTAIL.n91 VTAIL.n1 1.44878
R1903 VTAIL.n316 VTAIL.n310 1.16414
R1904 VTAIL.n357 VTAIL.n355 1.16414
R1905 VTAIL.n365 VTAIL.n288 1.16414
R1906 VTAIL.n34 VTAIL.n28 1.16414
R1907 VTAIL.n75 VTAIL.n73 1.16414
R1908 VTAIL.n83 VTAIL.n6 1.16414
R1909 VTAIL.n275 VTAIL.n198 1.16414
R1910 VTAIL.n267 VTAIL.n266 1.16414
R1911 VTAIL.n227 VTAIL.n221 1.16414
R1912 VTAIL.n181 VTAIL.n104 1.16414
R1913 VTAIL.n173 VTAIL.n172 1.16414
R1914 VTAIL.n133 VTAIL.n127 1.16414
R1915 VTAIL VTAIL.n375 0.431534
R1916 VTAIL.n315 VTAIL.n312 0.388379
R1917 VTAIL.n356 VTAIL.n290 0.388379
R1918 VTAIL.n362 VTAIL.n361 0.388379
R1919 VTAIL.n33 VTAIL.n30 0.388379
R1920 VTAIL.n74 VTAIL.n8 0.388379
R1921 VTAIL.n80 VTAIL.n79 0.388379
R1922 VTAIL.n272 VTAIL.n271 0.388379
R1923 VTAIL.n202 VTAIL.n200 0.388379
R1924 VTAIL.n226 VTAIL.n223 0.388379
R1925 VTAIL.n178 VTAIL.n177 0.388379
R1926 VTAIL.n108 VTAIL.n106 0.388379
R1927 VTAIL.n132 VTAIL.n129 0.388379
R1928 VTAIL.n314 VTAIL.n309 0.155672
R1929 VTAIL.n321 VTAIL.n309 0.155672
R1930 VTAIL.n322 VTAIL.n321 0.155672
R1931 VTAIL.n322 VTAIL.n305 0.155672
R1932 VTAIL.n329 VTAIL.n305 0.155672
R1933 VTAIL.n330 VTAIL.n329 0.155672
R1934 VTAIL.n330 VTAIL.n301 0.155672
R1935 VTAIL.n337 VTAIL.n301 0.155672
R1936 VTAIL.n338 VTAIL.n337 0.155672
R1937 VTAIL.n338 VTAIL.n297 0.155672
R1938 VTAIL.n345 VTAIL.n297 0.155672
R1939 VTAIL.n346 VTAIL.n345 0.155672
R1940 VTAIL.n346 VTAIL.n293 0.155672
R1941 VTAIL.n353 VTAIL.n293 0.155672
R1942 VTAIL.n354 VTAIL.n353 0.155672
R1943 VTAIL.n354 VTAIL.n289 0.155672
R1944 VTAIL.n363 VTAIL.n289 0.155672
R1945 VTAIL.n364 VTAIL.n363 0.155672
R1946 VTAIL.n364 VTAIL.n285 0.155672
R1947 VTAIL.n371 VTAIL.n285 0.155672
R1948 VTAIL.n32 VTAIL.n27 0.155672
R1949 VTAIL.n39 VTAIL.n27 0.155672
R1950 VTAIL.n40 VTAIL.n39 0.155672
R1951 VTAIL.n40 VTAIL.n23 0.155672
R1952 VTAIL.n47 VTAIL.n23 0.155672
R1953 VTAIL.n48 VTAIL.n47 0.155672
R1954 VTAIL.n48 VTAIL.n19 0.155672
R1955 VTAIL.n55 VTAIL.n19 0.155672
R1956 VTAIL.n56 VTAIL.n55 0.155672
R1957 VTAIL.n56 VTAIL.n15 0.155672
R1958 VTAIL.n63 VTAIL.n15 0.155672
R1959 VTAIL.n64 VTAIL.n63 0.155672
R1960 VTAIL.n64 VTAIL.n11 0.155672
R1961 VTAIL.n71 VTAIL.n11 0.155672
R1962 VTAIL.n72 VTAIL.n71 0.155672
R1963 VTAIL.n72 VTAIL.n7 0.155672
R1964 VTAIL.n81 VTAIL.n7 0.155672
R1965 VTAIL.n82 VTAIL.n81 0.155672
R1966 VTAIL.n82 VTAIL.n3 0.155672
R1967 VTAIL.n89 VTAIL.n3 0.155672
R1968 VTAIL.n281 VTAIL.n195 0.155672
R1969 VTAIL.n274 VTAIL.n195 0.155672
R1970 VTAIL.n274 VTAIL.n273 0.155672
R1971 VTAIL.n273 VTAIL.n199 0.155672
R1972 VTAIL.n265 VTAIL.n199 0.155672
R1973 VTAIL.n265 VTAIL.n264 0.155672
R1974 VTAIL.n264 VTAIL.n204 0.155672
R1975 VTAIL.n257 VTAIL.n204 0.155672
R1976 VTAIL.n257 VTAIL.n256 0.155672
R1977 VTAIL.n256 VTAIL.n208 0.155672
R1978 VTAIL.n249 VTAIL.n208 0.155672
R1979 VTAIL.n249 VTAIL.n248 0.155672
R1980 VTAIL.n248 VTAIL.n212 0.155672
R1981 VTAIL.n241 VTAIL.n212 0.155672
R1982 VTAIL.n241 VTAIL.n240 0.155672
R1983 VTAIL.n240 VTAIL.n216 0.155672
R1984 VTAIL.n233 VTAIL.n216 0.155672
R1985 VTAIL.n233 VTAIL.n232 0.155672
R1986 VTAIL.n232 VTAIL.n220 0.155672
R1987 VTAIL.n225 VTAIL.n220 0.155672
R1988 VTAIL.n187 VTAIL.n101 0.155672
R1989 VTAIL.n180 VTAIL.n101 0.155672
R1990 VTAIL.n180 VTAIL.n179 0.155672
R1991 VTAIL.n179 VTAIL.n105 0.155672
R1992 VTAIL.n171 VTAIL.n105 0.155672
R1993 VTAIL.n171 VTAIL.n170 0.155672
R1994 VTAIL.n170 VTAIL.n110 0.155672
R1995 VTAIL.n163 VTAIL.n110 0.155672
R1996 VTAIL.n163 VTAIL.n162 0.155672
R1997 VTAIL.n162 VTAIL.n114 0.155672
R1998 VTAIL.n155 VTAIL.n114 0.155672
R1999 VTAIL.n155 VTAIL.n154 0.155672
R2000 VTAIL.n154 VTAIL.n118 0.155672
R2001 VTAIL.n147 VTAIL.n118 0.155672
R2002 VTAIL.n147 VTAIL.n146 0.155672
R2003 VTAIL.n146 VTAIL.n122 0.155672
R2004 VTAIL.n139 VTAIL.n122 0.155672
R2005 VTAIL.n139 VTAIL.n138 0.155672
R2006 VTAIL.n138 VTAIL.n126 0.155672
R2007 VTAIL.n131 VTAIL.n126 0.155672
R2008 VDD1.n84 VDD1.n0 756.745
R2009 VDD1.n175 VDD1.n91 756.745
R2010 VDD1.n85 VDD1.n84 585
R2011 VDD1.n83 VDD1.n82 585
R2012 VDD1.n4 VDD1.n3 585
R2013 VDD1.n77 VDD1.n76 585
R2014 VDD1.n75 VDD1.n6 585
R2015 VDD1.n74 VDD1.n73 585
R2016 VDD1.n9 VDD1.n7 585
R2017 VDD1.n68 VDD1.n67 585
R2018 VDD1.n66 VDD1.n65 585
R2019 VDD1.n13 VDD1.n12 585
R2020 VDD1.n60 VDD1.n59 585
R2021 VDD1.n58 VDD1.n57 585
R2022 VDD1.n17 VDD1.n16 585
R2023 VDD1.n52 VDD1.n51 585
R2024 VDD1.n50 VDD1.n49 585
R2025 VDD1.n21 VDD1.n20 585
R2026 VDD1.n44 VDD1.n43 585
R2027 VDD1.n42 VDD1.n41 585
R2028 VDD1.n25 VDD1.n24 585
R2029 VDD1.n36 VDD1.n35 585
R2030 VDD1.n34 VDD1.n33 585
R2031 VDD1.n29 VDD1.n28 585
R2032 VDD1.n119 VDD1.n118 585
R2033 VDD1.n124 VDD1.n123 585
R2034 VDD1.n126 VDD1.n125 585
R2035 VDD1.n115 VDD1.n114 585
R2036 VDD1.n132 VDD1.n131 585
R2037 VDD1.n134 VDD1.n133 585
R2038 VDD1.n111 VDD1.n110 585
R2039 VDD1.n140 VDD1.n139 585
R2040 VDD1.n142 VDD1.n141 585
R2041 VDD1.n107 VDD1.n106 585
R2042 VDD1.n148 VDD1.n147 585
R2043 VDD1.n150 VDD1.n149 585
R2044 VDD1.n103 VDD1.n102 585
R2045 VDD1.n156 VDD1.n155 585
R2046 VDD1.n158 VDD1.n157 585
R2047 VDD1.n99 VDD1.n98 585
R2048 VDD1.n165 VDD1.n164 585
R2049 VDD1.n166 VDD1.n97 585
R2050 VDD1.n168 VDD1.n167 585
R2051 VDD1.n95 VDD1.n94 585
R2052 VDD1.n174 VDD1.n173 585
R2053 VDD1.n176 VDD1.n175 585
R2054 VDD1.n30 VDD1.t9 327.466
R2055 VDD1.n120 VDD1.t1 327.466
R2056 VDD1.n84 VDD1.n83 171.744
R2057 VDD1.n83 VDD1.n3 171.744
R2058 VDD1.n76 VDD1.n3 171.744
R2059 VDD1.n76 VDD1.n75 171.744
R2060 VDD1.n75 VDD1.n74 171.744
R2061 VDD1.n74 VDD1.n7 171.744
R2062 VDD1.n67 VDD1.n7 171.744
R2063 VDD1.n67 VDD1.n66 171.744
R2064 VDD1.n66 VDD1.n12 171.744
R2065 VDD1.n59 VDD1.n12 171.744
R2066 VDD1.n59 VDD1.n58 171.744
R2067 VDD1.n58 VDD1.n16 171.744
R2068 VDD1.n51 VDD1.n16 171.744
R2069 VDD1.n51 VDD1.n50 171.744
R2070 VDD1.n50 VDD1.n20 171.744
R2071 VDD1.n43 VDD1.n20 171.744
R2072 VDD1.n43 VDD1.n42 171.744
R2073 VDD1.n42 VDD1.n24 171.744
R2074 VDD1.n35 VDD1.n24 171.744
R2075 VDD1.n35 VDD1.n34 171.744
R2076 VDD1.n34 VDD1.n28 171.744
R2077 VDD1.n124 VDD1.n118 171.744
R2078 VDD1.n125 VDD1.n124 171.744
R2079 VDD1.n125 VDD1.n114 171.744
R2080 VDD1.n132 VDD1.n114 171.744
R2081 VDD1.n133 VDD1.n132 171.744
R2082 VDD1.n133 VDD1.n110 171.744
R2083 VDD1.n140 VDD1.n110 171.744
R2084 VDD1.n141 VDD1.n140 171.744
R2085 VDD1.n141 VDD1.n106 171.744
R2086 VDD1.n148 VDD1.n106 171.744
R2087 VDD1.n149 VDD1.n148 171.744
R2088 VDD1.n149 VDD1.n102 171.744
R2089 VDD1.n156 VDD1.n102 171.744
R2090 VDD1.n157 VDD1.n156 171.744
R2091 VDD1.n157 VDD1.n98 171.744
R2092 VDD1.n165 VDD1.n98 171.744
R2093 VDD1.n166 VDD1.n165 171.744
R2094 VDD1.n167 VDD1.n166 171.744
R2095 VDD1.n167 VDD1.n94 171.744
R2096 VDD1.n174 VDD1.n94 171.744
R2097 VDD1.n175 VDD1.n174 171.744
R2098 VDD1.t9 VDD1.n28 85.8723
R2099 VDD1.t1 VDD1.n118 85.8723
R2100 VDD1.n183 VDD1.n182 72.7658
R2101 VDD1.n90 VDD1.n89 71.3537
R2102 VDD1.n185 VDD1.n184 71.3535
R2103 VDD1.n181 VDD1.n180 71.3535
R2104 VDD1.n90 VDD1.n88 52.3725
R2105 VDD1.n181 VDD1.n179 52.3725
R2106 VDD1.n185 VDD1.n183 48.5031
R2107 VDD1.n30 VDD1.n29 16.3895
R2108 VDD1.n120 VDD1.n119 16.3895
R2109 VDD1.n77 VDD1.n6 13.1884
R2110 VDD1.n168 VDD1.n97 13.1884
R2111 VDD1.n78 VDD1.n4 12.8005
R2112 VDD1.n73 VDD1.n8 12.8005
R2113 VDD1.n33 VDD1.n32 12.8005
R2114 VDD1.n123 VDD1.n122 12.8005
R2115 VDD1.n164 VDD1.n163 12.8005
R2116 VDD1.n169 VDD1.n95 12.8005
R2117 VDD1.n82 VDD1.n81 12.0247
R2118 VDD1.n72 VDD1.n9 12.0247
R2119 VDD1.n36 VDD1.n27 12.0247
R2120 VDD1.n126 VDD1.n117 12.0247
R2121 VDD1.n162 VDD1.n99 12.0247
R2122 VDD1.n173 VDD1.n172 12.0247
R2123 VDD1.n85 VDD1.n2 11.249
R2124 VDD1.n69 VDD1.n68 11.249
R2125 VDD1.n37 VDD1.n25 11.249
R2126 VDD1.n127 VDD1.n115 11.249
R2127 VDD1.n159 VDD1.n158 11.249
R2128 VDD1.n176 VDD1.n93 11.249
R2129 VDD1.n86 VDD1.n0 10.4732
R2130 VDD1.n65 VDD1.n11 10.4732
R2131 VDD1.n41 VDD1.n40 10.4732
R2132 VDD1.n131 VDD1.n130 10.4732
R2133 VDD1.n155 VDD1.n101 10.4732
R2134 VDD1.n177 VDD1.n91 10.4732
R2135 VDD1.n64 VDD1.n13 9.69747
R2136 VDD1.n44 VDD1.n23 9.69747
R2137 VDD1.n134 VDD1.n113 9.69747
R2138 VDD1.n154 VDD1.n103 9.69747
R2139 VDD1.n88 VDD1.n87 9.45567
R2140 VDD1.n179 VDD1.n178 9.45567
R2141 VDD1.n56 VDD1.n55 9.3005
R2142 VDD1.n15 VDD1.n14 9.3005
R2143 VDD1.n62 VDD1.n61 9.3005
R2144 VDD1.n64 VDD1.n63 9.3005
R2145 VDD1.n11 VDD1.n10 9.3005
R2146 VDD1.n70 VDD1.n69 9.3005
R2147 VDD1.n72 VDD1.n71 9.3005
R2148 VDD1.n8 VDD1.n5 9.3005
R2149 VDD1.n87 VDD1.n86 9.3005
R2150 VDD1.n2 VDD1.n1 9.3005
R2151 VDD1.n81 VDD1.n80 9.3005
R2152 VDD1.n79 VDD1.n78 9.3005
R2153 VDD1.n54 VDD1.n53 9.3005
R2154 VDD1.n19 VDD1.n18 9.3005
R2155 VDD1.n48 VDD1.n47 9.3005
R2156 VDD1.n46 VDD1.n45 9.3005
R2157 VDD1.n23 VDD1.n22 9.3005
R2158 VDD1.n40 VDD1.n39 9.3005
R2159 VDD1.n38 VDD1.n37 9.3005
R2160 VDD1.n27 VDD1.n26 9.3005
R2161 VDD1.n32 VDD1.n31 9.3005
R2162 VDD1.n178 VDD1.n177 9.3005
R2163 VDD1.n93 VDD1.n92 9.3005
R2164 VDD1.n172 VDD1.n171 9.3005
R2165 VDD1.n170 VDD1.n169 9.3005
R2166 VDD1.n109 VDD1.n108 9.3005
R2167 VDD1.n138 VDD1.n137 9.3005
R2168 VDD1.n136 VDD1.n135 9.3005
R2169 VDD1.n113 VDD1.n112 9.3005
R2170 VDD1.n130 VDD1.n129 9.3005
R2171 VDD1.n128 VDD1.n127 9.3005
R2172 VDD1.n117 VDD1.n116 9.3005
R2173 VDD1.n122 VDD1.n121 9.3005
R2174 VDD1.n144 VDD1.n143 9.3005
R2175 VDD1.n146 VDD1.n145 9.3005
R2176 VDD1.n105 VDD1.n104 9.3005
R2177 VDD1.n152 VDD1.n151 9.3005
R2178 VDD1.n154 VDD1.n153 9.3005
R2179 VDD1.n101 VDD1.n100 9.3005
R2180 VDD1.n160 VDD1.n159 9.3005
R2181 VDD1.n162 VDD1.n161 9.3005
R2182 VDD1.n163 VDD1.n96 9.3005
R2183 VDD1.n61 VDD1.n60 8.92171
R2184 VDD1.n45 VDD1.n21 8.92171
R2185 VDD1.n135 VDD1.n111 8.92171
R2186 VDD1.n151 VDD1.n150 8.92171
R2187 VDD1.n57 VDD1.n15 8.14595
R2188 VDD1.n49 VDD1.n48 8.14595
R2189 VDD1.n139 VDD1.n138 8.14595
R2190 VDD1.n147 VDD1.n105 8.14595
R2191 VDD1.n56 VDD1.n17 7.3702
R2192 VDD1.n52 VDD1.n19 7.3702
R2193 VDD1.n142 VDD1.n109 7.3702
R2194 VDD1.n146 VDD1.n107 7.3702
R2195 VDD1.n53 VDD1.n17 6.59444
R2196 VDD1.n53 VDD1.n52 6.59444
R2197 VDD1.n143 VDD1.n142 6.59444
R2198 VDD1.n143 VDD1.n107 6.59444
R2199 VDD1.n57 VDD1.n56 5.81868
R2200 VDD1.n49 VDD1.n19 5.81868
R2201 VDD1.n139 VDD1.n109 5.81868
R2202 VDD1.n147 VDD1.n146 5.81868
R2203 VDD1.n60 VDD1.n15 5.04292
R2204 VDD1.n48 VDD1.n21 5.04292
R2205 VDD1.n138 VDD1.n111 5.04292
R2206 VDD1.n150 VDD1.n105 5.04292
R2207 VDD1.n61 VDD1.n13 4.26717
R2208 VDD1.n45 VDD1.n44 4.26717
R2209 VDD1.n135 VDD1.n134 4.26717
R2210 VDD1.n151 VDD1.n103 4.26717
R2211 VDD1.n31 VDD1.n30 3.70982
R2212 VDD1.n121 VDD1.n120 3.70982
R2213 VDD1.n88 VDD1.n0 3.49141
R2214 VDD1.n65 VDD1.n64 3.49141
R2215 VDD1.n41 VDD1.n23 3.49141
R2216 VDD1.n131 VDD1.n113 3.49141
R2217 VDD1.n155 VDD1.n154 3.49141
R2218 VDD1.n179 VDD1.n91 3.49141
R2219 VDD1.n86 VDD1.n85 2.71565
R2220 VDD1.n68 VDD1.n11 2.71565
R2221 VDD1.n40 VDD1.n25 2.71565
R2222 VDD1.n130 VDD1.n115 2.71565
R2223 VDD1.n158 VDD1.n101 2.71565
R2224 VDD1.n177 VDD1.n176 2.71565
R2225 VDD1.n184 VDD1.t2 2.01195
R2226 VDD1.n184 VDD1.t7 2.01195
R2227 VDD1.n89 VDD1.t6 2.01195
R2228 VDD1.n89 VDD1.t5 2.01195
R2229 VDD1.n182 VDD1.t0 2.01195
R2230 VDD1.n182 VDD1.t3 2.01195
R2231 VDD1.n180 VDD1.t4 2.01195
R2232 VDD1.n180 VDD1.t8 2.01195
R2233 VDD1.n82 VDD1.n2 1.93989
R2234 VDD1.n69 VDD1.n9 1.93989
R2235 VDD1.n37 VDD1.n36 1.93989
R2236 VDD1.n127 VDD1.n126 1.93989
R2237 VDD1.n159 VDD1.n99 1.93989
R2238 VDD1.n173 VDD1.n93 1.93989
R2239 VDD1 VDD1.n185 1.40998
R2240 VDD1.n81 VDD1.n4 1.16414
R2241 VDD1.n73 VDD1.n72 1.16414
R2242 VDD1.n33 VDD1.n27 1.16414
R2243 VDD1.n123 VDD1.n117 1.16414
R2244 VDD1.n164 VDD1.n162 1.16414
R2245 VDD1.n172 VDD1.n95 1.16414
R2246 VDD1 VDD1.n90 0.547914
R2247 VDD1.n183 VDD1.n181 0.434378
R2248 VDD1.n78 VDD1.n77 0.388379
R2249 VDD1.n8 VDD1.n6 0.388379
R2250 VDD1.n32 VDD1.n29 0.388379
R2251 VDD1.n122 VDD1.n119 0.388379
R2252 VDD1.n163 VDD1.n97 0.388379
R2253 VDD1.n169 VDD1.n168 0.388379
R2254 VDD1.n87 VDD1.n1 0.155672
R2255 VDD1.n80 VDD1.n1 0.155672
R2256 VDD1.n80 VDD1.n79 0.155672
R2257 VDD1.n79 VDD1.n5 0.155672
R2258 VDD1.n71 VDD1.n5 0.155672
R2259 VDD1.n71 VDD1.n70 0.155672
R2260 VDD1.n70 VDD1.n10 0.155672
R2261 VDD1.n63 VDD1.n10 0.155672
R2262 VDD1.n63 VDD1.n62 0.155672
R2263 VDD1.n62 VDD1.n14 0.155672
R2264 VDD1.n55 VDD1.n14 0.155672
R2265 VDD1.n55 VDD1.n54 0.155672
R2266 VDD1.n54 VDD1.n18 0.155672
R2267 VDD1.n47 VDD1.n18 0.155672
R2268 VDD1.n47 VDD1.n46 0.155672
R2269 VDD1.n46 VDD1.n22 0.155672
R2270 VDD1.n39 VDD1.n22 0.155672
R2271 VDD1.n39 VDD1.n38 0.155672
R2272 VDD1.n38 VDD1.n26 0.155672
R2273 VDD1.n31 VDD1.n26 0.155672
R2274 VDD1.n121 VDD1.n116 0.155672
R2275 VDD1.n128 VDD1.n116 0.155672
R2276 VDD1.n129 VDD1.n128 0.155672
R2277 VDD1.n129 VDD1.n112 0.155672
R2278 VDD1.n136 VDD1.n112 0.155672
R2279 VDD1.n137 VDD1.n136 0.155672
R2280 VDD1.n137 VDD1.n108 0.155672
R2281 VDD1.n144 VDD1.n108 0.155672
R2282 VDD1.n145 VDD1.n144 0.155672
R2283 VDD1.n145 VDD1.n104 0.155672
R2284 VDD1.n152 VDD1.n104 0.155672
R2285 VDD1.n153 VDD1.n152 0.155672
R2286 VDD1.n153 VDD1.n100 0.155672
R2287 VDD1.n160 VDD1.n100 0.155672
R2288 VDD1.n161 VDD1.n160 0.155672
R2289 VDD1.n161 VDD1.n96 0.155672
R2290 VDD1.n170 VDD1.n96 0.155672
R2291 VDD1.n171 VDD1.n170 0.155672
R2292 VDD1.n171 VDD1.n92 0.155672
R2293 VDD1.n178 VDD1.n92 0.155672
R2294 VN.n8 VN.t8 233.626
R2295 VN.n41 VN.t3 233.626
R2296 VN.n16 VN.t2 200.751
R2297 VN.n7 VN.t7 200.751
R2298 VN.n23 VN.t1 200.751
R2299 VN.n31 VN.t6 200.751
R2300 VN.n49 VN.t0 200.751
R2301 VN.n40 VN.t4 200.751
R2302 VN.n56 VN.t5 200.751
R2303 VN.n64 VN.t9 200.751
R2304 VN.n32 VN.n31 183.924
R2305 VN.n65 VN.n64 183.924
R2306 VN.n63 VN.n33 161.3
R2307 VN.n62 VN.n61 161.3
R2308 VN.n60 VN.n34 161.3
R2309 VN.n59 VN.n58 161.3
R2310 VN.n57 VN.n35 161.3
R2311 VN.n55 VN.n54 161.3
R2312 VN.n53 VN.n36 161.3
R2313 VN.n52 VN.n51 161.3
R2314 VN.n50 VN.n37 161.3
R2315 VN.n49 VN.n48 161.3
R2316 VN.n47 VN.n38 161.3
R2317 VN.n46 VN.n45 161.3
R2318 VN.n44 VN.n39 161.3
R2319 VN.n43 VN.n42 161.3
R2320 VN.n30 VN.n0 161.3
R2321 VN.n29 VN.n28 161.3
R2322 VN.n27 VN.n1 161.3
R2323 VN.n26 VN.n25 161.3
R2324 VN.n24 VN.n2 161.3
R2325 VN.n22 VN.n21 161.3
R2326 VN.n20 VN.n3 161.3
R2327 VN.n19 VN.n18 161.3
R2328 VN.n17 VN.n4 161.3
R2329 VN.n16 VN.n15 161.3
R2330 VN.n14 VN.n5 161.3
R2331 VN.n13 VN.n12 161.3
R2332 VN.n11 VN.n6 161.3
R2333 VN.n10 VN.n9 161.3
R2334 VN.n8 VN.n7 56.9995
R2335 VN.n41 VN.n40 56.9995
R2336 VN.n12 VN.n11 53.6554
R2337 VN.n18 VN.n3 53.6554
R2338 VN.n45 VN.n44 53.6554
R2339 VN.n51 VN.n36 53.6554
R2340 VN VN.n65 52.9683
R2341 VN.n25 VN.n1 49.7803
R2342 VN.n58 VN.n34 49.7803
R2343 VN.n29 VN.n1 31.3737
R2344 VN.n62 VN.n34 31.3737
R2345 VN.n12 VN.n5 27.4986
R2346 VN.n18 VN.n17 27.4986
R2347 VN.n45 VN.n38 27.4986
R2348 VN.n51 VN.n50 27.4986
R2349 VN.n11 VN.n10 24.5923
R2350 VN.n16 VN.n5 24.5923
R2351 VN.n17 VN.n16 24.5923
R2352 VN.n22 VN.n3 24.5923
R2353 VN.n25 VN.n24 24.5923
R2354 VN.n30 VN.n29 24.5923
R2355 VN.n44 VN.n43 24.5923
R2356 VN.n50 VN.n49 24.5923
R2357 VN.n49 VN.n38 24.5923
R2358 VN.n58 VN.n57 24.5923
R2359 VN.n55 VN.n36 24.5923
R2360 VN.n63 VN.n62 24.5923
R2361 VN.n10 VN.n7 13.2801
R2362 VN.n23 VN.n22 13.2801
R2363 VN.n43 VN.n40 13.2801
R2364 VN.n56 VN.n55 13.2801
R2365 VN.n42 VN.n41 12.447
R2366 VN.n9 VN.n8 12.447
R2367 VN.n24 VN.n23 11.3127
R2368 VN.n57 VN.n56 11.3127
R2369 VN.n31 VN.n30 1.96785
R2370 VN.n64 VN.n63 1.96785
R2371 VN.n65 VN.n33 0.189894
R2372 VN.n61 VN.n33 0.189894
R2373 VN.n61 VN.n60 0.189894
R2374 VN.n60 VN.n59 0.189894
R2375 VN.n59 VN.n35 0.189894
R2376 VN.n54 VN.n35 0.189894
R2377 VN.n54 VN.n53 0.189894
R2378 VN.n53 VN.n52 0.189894
R2379 VN.n52 VN.n37 0.189894
R2380 VN.n48 VN.n37 0.189894
R2381 VN.n48 VN.n47 0.189894
R2382 VN.n47 VN.n46 0.189894
R2383 VN.n46 VN.n39 0.189894
R2384 VN.n42 VN.n39 0.189894
R2385 VN.n9 VN.n6 0.189894
R2386 VN.n13 VN.n6 0.189894
R2387 VN.n14 VN.n13 0.189894
R2388 VN.n15 VN.n14 0.189894
R2389 VN.n15 VN.n4 0.189894
R2390 VN.n19 VN.n4 0.189894
R2391 VN.n20 VN.n19 0.189894
R2392 VN.n21 VN.n20 0.189894
R2393 VN.n21 VN.n2 0.189894
R2394 VN.n26 VN.n2 0.189894
R2395 VN.n27 VN.n26 0.189894
R2396 VN.n28 VN.n27 0.189894
R2397 VN.n28 VN.n0 0.189894
R2398 VN.n32 VN.n0 0.189894
R2399 VN VN.n32 0.0516364
R2400 VDD2.n177 VDD2.n93 756.745
R2401 VDD2.n84 VDD2.n0 756.745
R2402 VDD2.n178 VDD2.n177 585
R2403 VDD2.n176 VDD2.n175 585
R2404 VDD2.n97 VDD2.n96 585
R2405 VDD2.n170 VDD2.n169 585
R2406 VDD2.n168 VDD2.n99 585
R2407 VDD2.n167 VDD2.n166 585
R2408 VDD2.n102 VDD2.n100 585
R2409 VDD2.n161 VDD2.n160 585
R2410 VDD2.n159 VDD2.n158 585
R2411 VDD2.n106 VDD2.n105 585
R2412 VDD2.n153 VDD2.n152 585
R2413 VDD2.n151 VDD2.n150 585
R2414 VDD2.n110 VDD2.n109 585
R2415 VDD2.n145 VDD2.n144 585
R2416 VDD2.n143 VDD2.n142 585
R2417 VDD2.n114 VDD2.n113 585
R2418 VDD2.n137 VDD2.n136 585
R2419 VDD2.n135 VDD2.n134 585
R2420 VDD2.n118 VDD2.n117 585
R2421 VDD2.n129 VDD2.n128 585
R2422 VDD2.n127 VDD2.n126 585
R2423 VDD2.n122 VDD2.n121 585
R2424 VDD2.n28 VDD2.n27 585
R2425 VDD2.n33 VDD2.n32 585
R2426 VDD2.n35 VDD2.n34 585
R2427 VDD2.n24 VDD2.n23 585
R2428 VDD2.n41 VDD2.n40 585
R2429 VDD2.n43 VDD2.n42 585
R2430 VDD2.n20 VDD2.n19 585
R2431 VDD2.n49 VDD2.n48 585
R2432 VDD2.n51 VDD2.n50 585
R2433 VDD2.n16 VDD2.n15 585
R2434 VDD2.n57 VDD2.n56 585
R2435 VDD2.n59 VDD2.n58 585
R2436 VDD2.n12 VDD2.n11 585
R2437 VDD2.n65 VDD2.n64 585
R2438 VDD2.n67 VDD2.n66 585
R2439 VDD2.n8 VDD2.n7 585
R2440 VDD2.n74 VDD2.n73 585
R2441 VDD2.n75 VDD2.n6 585
R2442 VDD2.n77 VDD2.n76 585
R2443 VDD2.n4 VDD2.n3 585
R2444 VDD2.n83 VDD2.n82 585
R2445 VDD2.n85 VDD2.n84 585
R2446 VDD2.n123 VDD2.t0 327.466
R2447 VDD2.n29 VDD2.t1 327.466
R2448 VDD2.n177 VDD2.n176 171.744
R2449 VDD2.n176 VDD2.n96 171.744
R2450 VDD2.n169 VDD2.n96 171.744
R2451 VDD2.n169 VDD2.n168 171.744
R2452 VDD2.n168 VDD2.n167 171.744
R2453 VDD2.n167 VDD2.n100 171.744
R2454 VDD2.n160 VDD2.n100 171.744
R2455 VDD2.n160 VDD2.n159 171.744
R2456 VDD2.n159 VDD2.n105 171.744
R2457 VDD2.n152 VDD2.n105 171.744
R2458 VDD2.n152 VDD2.n151 171.744
R2459 VDD2.n151 VDD2.n109 171.744
R2460 VDD2.n144 VDD2.n109 171.744
R2461 VDD2.n144 VDD2.n143 171.744
R2462 VDD2.n143 VDD2.n113 171.744
R2463 VDD2.n136 VDD2.n113 171.744
R2464 VDD2.n136 VDD2.n135 171.744
R2465 VDD2.n135 VDD2.n117 171.744
R2466 VDD2.n128 VDD2.n117 171.744
R2467 VDD2.n128 VDD2.n127 171.744
R2468 VDD2.n127 VDD2.n121 171.744
R2469 VDD2.n33 VDD2.n27 171.744
R2470 VDD2.n34 VDD2.n33 171.744
R2471 VDD2.n34 VDD2.n23 171.744
R2472 VDD2.n41 VDD2.n23 171.744
R2473 VDD2.n42 VDD2.n41 171.744
R2474 VDD2.n42 VDD2.n19 171.744
R2475 VDD2.n49 VDD2.n19 171.744
R2476 VDD2.n50 VDD2.n49 171.744
R2477 VDD2.n50 VDD2.n15 171.744
R2478 VDD2.n57 VDD2.n15 171.744
R2479 VDD2.n58 VDD2.n57 171.744
R2480 VDD2.n58 VDD2.n11 171.744
R2481 VDD2.n65 VDD2.n11 171.744
R2482 VDD2.n66 VDD2.n65 171.744
R2483 VDD2.n66 VDD2.n7 171.744
R2484 VDD2.n74 VDD2.n7 171.744
R2485 VDD2.n75 VDD2.n74 171.744
R2486 VDD2.n76 VDD2.n75 171.744
R2487 VDD2.n76 VDD2.n3 171.744
R2488 VDD2.n83 VDD2.n3 171.744
R2489 VDD2.n84 VDD2.n83 171.744
R2490 VDD2.t0 VDD2.n121 85.8723
R2491 VDD2.t1 VDD2.n27 85.8723
R2492 VDD2.n92 VDD2.n91 72.7658
R2493 VDD2 VDD2.n185 72.7629
R2494 VDD2.n184 VDD2.n183 71.3537
R2495 VDD2.n90 VDD2.n89 71.3535
R2496 VDD2.n90 VDD2.n88 52.3725
R2497 VDD2.n182 VDD2.n181 50.4157
R2498 VDD2.n182 VDD2.n92 46.9416
R2499 VDD2.n123 VDD2.n122 16.3895
R2500 VDD2.n29 VDD2.n28 16.3895
R2501 VDD2.n170 VDD2.n99 13.1884
R2502 VDD2.n77 VDD2.n6 13.1884
R2503 VDD2.n171 VDD2.n97 12.8005
R2504 VDD2.n166 VDD2.n101 12.8005
R2505 VDD2.n126 VDD2.n125 12.8005
R2506 VDD2.n32 VDD2.n31 12.8005
R2507 VDD2.n73 VDD2.n72 12.8005
R2508 VDD2.n78 VDD2.n4 12.8005
R2509 VDD2.n175 VDD2.n174 12.0247
R2510 VDD2.n165 VDD2.n102 12.0247
R2511 VDD2.n129 VDD2.n120 12.0247
R2512 VDD2.n35 VDD2.n26 12.0247
R2513 VDD2.n71 VDD2.n8 12.0247
R2514 VDD2.n82 VDD2.n81 12.0247
R2515 VDD2.n178 VDD2.n95 11.249
R2516 VDD2.n162 VDD2.n161 11.249
R2517 VDD2.n130 VDD2.n118 11.249
R2518 VDD2.n36 VDD2.n24 11.249
R2519 VDD2.n68 VDD2.n67 11.249
R2520 VDD2.n85 VDD2.n2 11.249
R2521 VDD2.n179 VDD2.n93 10.4732
R2522 VDD2.n158 VDD2.n104 10.4732
R2523 VDD2.n134 VDD2.n133 10.4732
R2524 VDD2.n40 VDD2.n39 10.4732
R2525 VDD2.n64 VDD2.n10 10.4732
R2526 VDD2.n86 VDD2.n0 10.4732
R2527 VDD2.n157 VDD2.n106 9.69747
R2528 VDD2.n137 VDD2.n116 9.69747
R2529 VDD2.n43 VDD2.n22 9.69747
R2530 VDD2.n63 VDD2.n12 9.69747
R2531 VDD2.n181 VDD2.n180 9.45567
R2532 VDD2.n88 VDD2.n87 9.45567
R2533 VDD2.n149 VDD2.n148 9.3005
R2534 VDD2.n108 VDD2.n107 9.3005
R2535 VDD2.n155 VDD2.n154 9.3005
R2536 VDD2.n157 VDD2.n156 9.3005
R2537 VDD2.n104 VDD2.n103 9.3005
R2538 VDD2.n163 VDD2.n162 9.3005
R2539 VDD2.n165 VDD2.n164 9.3005
R2540 VDD2.n101 VDD2.n98 9.3005
R2541 VDD2.n180 VDD2.n179 9.3005
R2542 VDD2.n95 VDD2.n94 9.3005
R2543 VDD2.n174 VDD2.n173 9.3005
R2544 VDD2.n172 VDD2.n171 9.3005
R2545 VDD2.n147 VDD2.n146 9.3005
R2546 VDD2.n112 VDD2.n111 9.3005
R2547 VDD2.n141 VDD2.n140 9.3005
R2548 VDD2.n139 VDD2.n138 9.3005
R2549 VDD2.n116 VDD2.n115 9.3005
R2550 VDD2.n133 VDD2.n132 9.3005
R2551 VDD2.n131 VDD2.n130 9.3005
R2552 VDD2.n120 VDD2.n119 9.3005
R2553 VDD2.n125 VDD2.n124 9.3005
R2554 VDD2.n87 VDD2.n86 9.3005
R2555 VDD2.n2 VDD2.n1 9.3005
R2556 VDD2.n81 VDD2.n80 9.3005
R2557 VDD2.n79 VDD2.n78 9.3005
R2558 VDD2.n18 VDD2.n17 9.3005
R2559 VDD2.n47 VDD2.n46 9.3005
R2560 VDD2.n45 VDD2.n44 9.3005
R2561 VDD2.n22 VDD2.n21 9.3005
R2562 VDD2.n39 VDD2.n38 9.3005
R2563 VDD2.n37 VDD2.n36 9.3005
R2564 VDD2.n26 VDD2.n25 9.3005
R2565 VDD2.n31 VDD2.n30 9.3005
R2566 VDD2.n53 VDD2.n52 9.3005
R2567 VDD2.n55 VDD2.n54 9.3005
R2568 VDD2.n14 VDD2.n13 9.3005
R2569 VDD2.n61 VDD2.n60 9.3005
R2570 VDD2.n63 VDD2.n62 9.3005
R2571 VDD2.n10 VDD2.n9 9.3005
R2572 VDD2.n69 VDD2.n68 9.3005
R2573 VDD2.n71 VDD2.n70 9.3005
R2574 VDD2.n72 VDD2.n5 9.3005
R2575 VDD2.n154 VDD2.n153 8.92171
R2576 VDD2.n138 VDD2.n114 8.92171
R2577 VDD2.n44 VDD2.n20 8.92171
R2578 VDD2.n60 VDD2.n59 8.92171
R2579 VDD2.n150 VDD2.n108 8.14595
R2580 VDD2.n142 VDD2.n141 8.14595
R2581 VDD2.n48 VDD2.n47 8.14595
R2582 VDD2.n56 VDD2.n14 8.14595
R2583 VDD2.n149 VDD2.n110 7.3702
R2584 VDD2.n145 VDD2.n112 7.3702
R2585 VDD2.n51 VDD2.n18 7.3702
R2586 VDD2.n55 VDD2.n16 7.3702
R2587 VDD2.n146 VDD2.n110 6.59444
R2588 VDD2.n146 VDD2.n145 6.59444
R2589 VDD2.n52 VDD2.n51 6.59444
R2590 VDD2.n52 VDD2.n16 6.59444
R2591 VDD2.n150 VDD2.n149 5.81868
R2592 VDD2.n142 VDD2.n112 5.81868
R2593 VDD2.n48 VDD2.n18 5.81868
R2594 VDD2.n56 VDD2.n55 5.81868
R2595 VDD2.n153 VDD2.n108 5.04292
R2596 VDD2.n141 VDD2.n114 5.04292
R2597 VDD2.n47 VDD2.n20 5.04292
R2598 VDD2.n59 VDD2.n14 5.04292
R2599 VDD2.n154 VDD2.n106 4.26717
R2600 VDD2.n138 VDD2.n137 4.26717
R2601 VDD2.n44 VDD2.n43 4.26717
R2602 VDD2.n60 VDD2.n12 4.26717
R2603 VDD2.n124 VDD2.n123 3.70982
R2604 VDD2.n30 VDD2.n29 3.70982
R2605 VDD2.n181 VDD2.n93 3.49141
R2606 VDD2.n158 VDD2.n157 3.49141
R2607 VDD2.n134 VDD2.n116 3.49141
R2608 VDD2.n40 VDD2.n22 3.49141
R2609 VDD2.n64 VDD2.n63 3.49141
R2610 VDD2.n88 VDD2.n0 3.49141
R2611 VDD2.n179 VDD2.n178 2.71565
R2612 VDD2.n161 VDD2.n104 2.71565
R2613 VDD2.n133 VDD2.n118 2.71565
R2614 VDD2.n39 VDD2.n24 2.71565
R2615 VDD2.n67 VDD2.n10 2.71565
R2616 VDD2.n86 VDD2.n85 2.71565
R2617 VDD2.n185 VDD2.t5 2.01195
R2618 VDD2.n185 VDD2.t6 2.01195
R2619 VDD2.n183 VDD2.t4 2.01195
R2620 VDD2.n183 VDD2.t9 2.01195
R2621 VDD2.n91 VDD2.t8 2.01195
R2622 VDD2.n91 VDD2.t3 2.01195
R2623 VDD2.n89 VDD2.t2 2.01195
R2624 VDD2.n89 VDD2.t7 2.01195
R2625 VDD2.n184 VDD2.n182 1.9574
R2626 VDD2.n175 VDD2.n95 1.93989
R2627 VDD2.n162 VDD2.n102 1.93989
R2628 VDD2.n130 VDD2.n129 1.93989
R2629 VDD2.n36 VDD2.n35 1.93989
R2630 VDD2.n68 VDD2.n8 1.93989
R2631 VDD2.n82 VDD2.n2 1.93989
R2632 VDD2.n174 VDD2.n97 1.16414
R2633 VDD2.n166 VDD2.n165 1.16414
R2634 VDD2.n126 VDD2.n120 1.16414
R2635 VDD2.n32 VDD2.n26 1.16414
R2636 VDD2.n73 VDD2.n71 1.16414
R2637 VDD2.n81 VDD2.n4 1.16414
R2638 VDD2 VDD2.n184 0.547914
R2639 VDD2.n92 VDD2.n90 0.434378
R2640 VDD2.n171 VDD2.n170 0.388379
R2641 VDD2.n101 VDD2.n99 0.388379
R2642 VDD2.n125 VDD2.n122 0.388379
R2643 VDD2.n31 VDD2.n28 0.388379
R2644 VDD2.n72 VDD2.n6 0.388379
R2645 VDD2.n78 VDD2.n77 0.388379
R2646 VDD2.n180 VDD2.n94 0.155672
R2647 VDD2.n173 VDD2.n94 0.155672
R2648 VDD2.n173 VDD2.n172 0.155672
R2649 VDD2.n172 VDD2.n98 0.155672
R2650 VDD2.n164 VDD2.n98 0.155672
R2651 VDD2.n164 VDD2.n163 0.155672
R2652 VDD2.n163 VDD2.n103 0.155672
R2653 VDD2.n156 VDD2.n103 0.155672
R2654 VDD2.n156 VDD2.n155 0.155672
R2655 VDD2.n155 VDD2.n107 0.155672
R2656 VDD2.n148 VDD2.n107 0.155672
R2657 VDD2.n148 VDD2.n147 0.155672
R2658 VDD2.n147 VDD2.n111 0.155672
R2659 VDD2.n140 VDD2.n111 0.155672
R2660 VDD2.n140 VDD2.n139 0.155672
R2661 VDD2.n139 VDD2.n115 0.155672
R2662 VDD2.n132 VDD2.n115 0.155672
R2663 VDD2.n132 VDD2.n131 0.155672
R2664 VDD2.n131 VDD2.n119 0.155672
R2665 VDD2.n124 VDD2.n119 0.155672
R2666 VDD2.n30 VDD2.n25 0.155672
R2667 VDD2.n37 VDD2.n25 0.155672
R2668 VDD2.n38 VDD2.n37 0.155672
R2669 VDD2.n38 VDD2.n21 0.155672
R2670 VDD2.n45 VDD2.n21 0.155672
R2671 VDD2.n46 VDD2.n45 0.155672
R2672 VDD2.n46 VDD2.n17 0.155672
R2673 VDD2.n53 VDD2.n17 0.155672
R2674 VDD2.n54 VDD2.n53 0.155672
R2675 VDD2.n54 VDD2.n13 0.155672
R2676 VDD2.n61 VDD2.n13 0.155672
R2677 VDD2.n62 VDD2.n61 0.155672
R2678 VDD2.n62 VDD2.n9 0.155672
R2679 VDD2.n69 VDD2.n9 0.155672
R2680 VDD2.n70 VDD2.n69 0.155672
R2681 VDD2.n70 VDD2.n5 0.155672
R2682 VDD2.n79 VDD2.n5 0.155672
R2683 VDD2.n80 VDD2.n79 0.155672
R2684 VDD2.n80 VDD2.n1 0.155672
R2685 VDD2.n87 VDD2.n1 0.155672
C0 VN VDD1 0.152137f
C1 w_n3694_n4200# VDD2 2.93932f
C2 VN VDD2 13.264501f
C3 VDD1 B 2.54224f
C4 VTAIL VDD1 12.709f
C5 VDD2 B 2.63445f
C6 VTAIL VDD2 12.753401f
C7 w_n3694_n4200# VP 8.24207f
C8 VN VP 8.188331f
C9 VDD1 VDD2 1.74536f
C10 VN w_n3694_n4200# 7.76316f
C11 B VP 1.96913f
C12 w_n3694_n4200# B 10.6034f
C13 VTAIL VP 13.4729f
C14 VN B 1.16747f
C15 VTAIL w_n3694_n4200# 3.72141f
C16 VN VTAIL 13.4585f
C17 VDD1 VP 13.607599f
C18 VTAIL B 4.32019f
C19 w_n3694_n4200# VDD1 2.82997f
C20 VDD2 VP 0.50012f
C21 VDD2 VSUBS 1.987389f
C22 VDD1 VSUBS 1.797193f
C23 VTAIL VSUBS 1.289803f
C24 VN VSUBS 6.7958f
C25 VP VSUBS 3.535051f
C26 B VSUBS 4.898168f
C27 w_n3694_n4200# VSUBS 0.190034p
C28 VDD2.n0 VSUBS 0.028914f
C29 VDD2.n1 VSUBS 0.026831f
C30 VDD2.n2 VSUBS 0.014418f
C31 VDD2.n3 VSUBS 0.034078f
C32 VDD2.n4 VSUBS 0.015266f
C33 VDD2.n5 VSUBS 0.026831f
C34 VDD2.n6 VSUBS 0.014842f
C35 VDD2.n7 VSUBS 0.034078f
C36 VDD2.n8 VSUBS 0.015266f
C37 VDD2.n9 VSUBS 0.026831f
C38 VDD2.n10 VSUBS 0.014418f
C39 VDD2.n11 VSUBS 0.034078f
C40 VDD2.n12 VSUBS 0.015266f
C41 VDD2.n13 VSUBS 0.026831f
C42 VDD2.n14 VSUBS 0.014418f
C43 VDD2.n15 VSUBS 0.034078f
C44 VDD2.n16 VSUBS 0.015266f
C45 VDD2.n17 VSUBS 0.026831f
C46 VDD2.n18 VSUBS 0.014418f
C47 VDD2.n19 VSUBS 0.034078f
C48 VDD2.n20 VSUBS 0.015266f
C49 VDD2.n21 VSUBS 0.026831f
C50 VDD2.n22 VSUBS 0.014418f
C51 VDD2.n23 VSUBS 0.034078f
C52 VDD2.n24 VSUBS 0.015266f
C53 VDD2.n25 VSUBS 0.026831f
C54 VDD2.n26 VSUBS 0.014418f
C55 VDD2.n27 VSUBS 0.025558f
C56 VDD2.n28 VSUBS 0.021679f
C57 VDD2.t1 VSUBS 0.073032f
C58 VDD2.n29 VSUBS 0.198313f
C59 VDD2.n30 VSUBS 1.85448f
C60 VDD2.n31 VSUBS 0.014418f
C61 VDD2.n32 VSUBS 0.015266f
C62 VDD2.n33 VSUBS 0.034078f
C63 VDD2.n34 VSUBS 0.034078f
C64 VDD2.n35 VSUBS 0.015266f
C65 VDD2.n36 VSUBS 0.014418f
C66 VDD2.n37 VSUBS 0.026831f
C67 VDD2.n38 VSUBS 0.026831f
C68 VDD2.n39 VSUBS 0.014418f
C69 VDD2.n40 VSUBS 0.015266f
C70 VDD2.n41 VSUBS 0.034078f
C71 VDD2.n42 VSUBS 0.034078f
C72 VDD2.n43 VSUBS 0.015266f
C73 VDD2.n44 VSUBS 0.014418f
C74 VDD2.n45 VSUBS 0.026831f
C75 VDD2.n46 VSUBS 0.026831f
C76 VDD2.n47 VSUBS 0.014418f
C77 VDD2.n48 VSUBS 0.015266f
C78 VDD2.n49 VSUBS 0.034078f
C79 VDD2.n50 VSUBS 0.034078f
C80 VDD2.n51 VSUBS 0.015266f
C81 VDD2.n52 VSUBS 0.014418f
C82 VDD2.n53 VSUBS 0.026831f
C83 VDD2.n54 VSUBS 0.026831f
C84 VDD2.n55 VSUBS 0.014418f
C85 VDD2.n56 VSUBS 0.015266f
C86 VDD2.n57 VSUBS 0.034078f
C87 VDD2.n58 VSUBS 0.034078f
C88 VDD2.n59 VSUBS 0.015266f
C89 VDD2.n60 VSUBS 0.014418f
C90 VDD2.n61 VSUBS 0.026831f
C91 VDD2.n62 VSUBS 0.026831f
C92 VDD2.n63 VSUBS 0.014418f
C93 VDD2.n64 VSUBS 0.015266f
C94 VDD2.n65 VSUBS 0.034078f
C95 VDD2.n66 VSUBS 0.034078f
C96 VDD2.n67 VSUBS 0.015266f
C97 VDD2.n68 VSUBS 0.014418f
C98 VDD2.n69 VSUBS 0.026831f
C99 VDD2.n70 VSUBS 0.026831f
C100 VDD2.n71 VSUBS 0.014418f
C101 VDD2.n72 VSUBS 0.014418f
C102 VDD2.n73 VSUBS 0.015266f
C103 VDD2.n74 VSUBS 0.034078f
C104 VDD2.n75 VSUBS 0.034078f
C105 VDD2.n76 VSUBS 0.034078f
C106 VDD2.n77 VSUBS 0.014842f
C107 VDD2.n78 VSUBS 0.014418f
C108 VDD2.n79 VSUBS 0.026831f
C109 VDD2.n80 VSUBS 0.026831f
C110 VDD2.n81 VSUBS 0.014418f
C111 VDD2.n82 VSUBS 0.015266f
C112 VDD2.n83 VSUBS 0.034078f
C113 VDD2.n84 VSUBS 0.080567f
C114 VDD2.n85 VSUBS 0.015266f
C115 VDD2.n86 VSUBS 0.014418f
C116 VDD2.n87 VSUBS 0.06495f
C117 VDD2.n88 VSUBS 0.067338f
C118 VDD2.t2 VSUBS 0.342631f
C119 VDD2.t7 VSUBS 0.342631f
C120 VDD2.n89 VSUBS 2.81429f
C121 VDD2.n90 VSUBS 0.936506f
C122 VDD2.t8 VSUBS 0.342631f
C123 VDD2.t3 VSUBS 0.342631f
C124 VDD2.n91 VSUBS 2.83014f
C125 VDD2.n92 VSUBS 3.31356f
C126 VDD2.n93 VSUBS 0.028914f
C127 VDD2.n94 VSUBS 0.026831f
C128 VDD2.n95 VSUBS 0.014418f
C129 VDD2.n96 VSUBS 0.034078f
C130 VDD2.n97 VSUBS 0.015266f
C131 VDD2.n98 VSUBS 0.026831f
C132 VDD2.n99 VSUBS 0.014842f
C133 VDD2.n100 VSUBS 0.034078f
C134 VDD2.n101 VSUBS 0.014418f
C135 VDD2.n102 VSUBS 0.015266f
C136 VDD2.n103 VSUBS 0.026831f
C137 VDD2.n104 VSUBS 0.014418f
C138 VDD2.n105 VSUBS 0.034078f
C139 VDD2.n106 VSUBS 0.015266f
C140 VDD2.n107 VSUBS 0.026831f
C141 VDD2.n108 VSUBS 0.014418f
C142 VDD2.n109 VSUBS 0.034078f
C143 VDD2.n110 VSUBS 0.015266f
C144 VDD2.n111 VSUBS 0.026831f
C145 VDD2.n112 VSUBS 0.014418f
C146 VDD2.n113 VSUBS 0.034078f
C147 VDD2.n114 VSUBS 0.015266f
C148 VDD2.n115 VSUBS 0.026831f
C149 VDD2.n116 VSUBS 0.014418f
C150 VDD2.n117 VSUBS 0.034078f
C151 VDD2.n118 VSUBS 0.015266f
C152 VDD2.n119 VSUBS 0.026831f
C153 VDD2.n120 VSUBS 0.014418f
C154 VDD2.n121 VSUBS 0.025558f
C155 VDD2.n122 VSUBS 0.021679f
C156 VDD2.t0 VSUBS 0.073032f
C157 VDD2.n123 VSUBS 0.198313f
C158 VDD2.n124 VSUBS 1.85448f
C159 VDD2.n125 VSUBS 0.014418f
C160 VDD2.n126 VSUBS 0.015266f
C161 VDD2.n127 VSUBS 0.034078f
C162 VDD2.n128 VSUBS 0.034078f
C163 VDD2.n129 VSUBS 0.015266f
C164 VDD2.n130 VSUBS 0.014418f
C165 VDD2.n131 VSUBS 0.026831f
C166 VDD2.n132 VSUBS 0.026831f
C167 VDD2.n133 VSUBS 0.014418f
C168 VDD2.n134 VSUBS 0.015266f
C169 VDD2.n135 VSUBS 0.034078f
C170 VDD2.n136 VSUBS 0.034078f
C171 VDD2.n137 VSUBS 0.015266f
C172 VDD2.n138 VSUBS 0.014418f
C173 VDD2.n139 VSUBS 0.026831f
C174 VDD2.n140 VSUBS 0.026831f
C175 VDD2.n141 VSUBS 0.014418f
C176 VDD2.n142 VSUBS 0.015266f
C177 VDD2.n143 VSUBS 0.034078f
C178 VDD2.n144 VSUBS 0.034078f
C179 VDD2.n145 VSUBS 0.015266f
C180 VDD2.n146 VSUBS 0.014418f
C181 VDD2.n147 VSUBS 0.026831f
C182 VDD2.n148 VSUBS 0.026831f
C183 VDD2.n149 VSUBS 0.014418f
C184 VDD2.n150 VSUBS 0.015266f
C185 VDD2.n151 VSUBS 0.034078f
C186 VDD2.n152 VSUBS 0.034078f
C187 VDD2.n153 VSUBS 0.015266f
C188 VDD2.n154 VSUBS 0.014418f
C189 VDD2.n155 VSUBS 0.026831f
C190 VDD2.n156 VSUBS 0.026831f
C191 VDD2.n157 VSUBS 0.014418f
C192 VDD2.n158 VSUBS 0.015266f
C193 VDD2.n159 VSUBS 0.034078f
C194 VDD2.n160 VSUBS 0.034078f
C195 VDD2.n161 VSUBS 0.015266f
C196 VDD2.n162 VSUBS 0.014418f
C197 VDD2.n163 VSUBS 0.026831f
C198 VDD2.n164 VSUBS 0.026831f
C199 VDD2.n165 VSUBS 0.014418f
C200 VDD2.n166 VSUBS 0.015266f
C201 VDD2.n167 VSUBS 0.034078f
C202 VDD2.n168 VSUBS 0.034078f
C203 VDD2.n169 VSUBS 0.034078f
C204 VDD2.n170 VSUBS 0.014842f
C205 VDD2.n171 VSUBS 0.014418f
C206 VDD2.n172 VSUBS 0.026831f
C207 VDD2.n173 VSUBS 0.026831f
C208 VDD2.n174 VSUBS 0.014418f
C209 VDD2.n175 VSUBS 0.015266f
C210 VDD2.n176 VSUBS 0.034078f
C211 VDD2.n177 VSUBS 0.080567f
C212 VDD2.n178 VSUBS 0.015266f
C213 VDD2.n179 VSUBS 0.014418f
C214 VDD2.n180 VSUBS 0.06495f
C215 VDD2.n181 VSUBS 0.059023f
C216 VDD2.n182 VSUBS 3.17096f
C217 VDD2.t4 VSUBS 0.342631f
C218 VDD2.t9 VSUBS 0.342631f
C219 VDD2.n183 VSUBS 2.8143f
C220 VDD2.n184 VSUBS 0.730666f
C221 VDD2.t5 VSUBS 0.342631f
C222 VDD2.t6 VSUBS 0.342631f
C223 VDD2.n185 VSUBS 2.83009f
C224 VN.n0 VSUBS 0.030824f
C225 VN.t6 VSUBS 2.65229f
C226 VN.n1 VSUBS 0.028634f
C227 VN.n2 VSUBS 0.030824f
C228 VN.t1 VSUBS 2.65229f
C229 VN.n3 VSUBS 0.054103f
C230 VN.n4 VSUBS 0.030824f
C231 VN.t2 VSUBS 2.65229f
C232 VN.n5 VSUBS 0.059785f
C233 VN.n6 VSUBS 0.030824f
C234 VN.t7 VSUBS 2.65229f
C235 VN.n7 VSUBS 1.00372f
C236 VN.t8 VSUBS 2.8048f
C237 VN.n8 VSUBS 1.00571f
C238 VN.n9 VSUBS 0.229729f
C239 VN.n10 VSUBS 0.04418f
C240 VN.n11 VSUBS 0.054103f
C241 VN.n12 VSUBS 0.032887f
C242 VN.n13 VSUBS 0.030824f
C243 VN.n14 VSUBS 0.030824f
C244 VN.n15 VSUBS 0.030824f
C245 VN.n16 VSUBS 0.959877f
C246 VN.n17 VSUBS 0.059785f
C247 VN.n18 VSUBS 0.032887f
C248 VN.n19 VSUBS 0.030824f
C249 VN.n20 VSUBS 0.030824f
C250 VN.n21 VSUBS 0.030824f
C251 VN.n22 VSUBS 0.04418f
C252 VN.n23 VSUBS 0.930935f
C253 VN.n24 VSUBS 0.041922f
C254 VN.n25 VSUBS 0.056589f
C255 VN.n26 VSUBS 0.030824f
C256 VN.n27 VSUBS 0.030824f
C257 VN.n28 VSUBS 0.030824f
C258 VN.n29 VSUBS 0.061552f
C259 VN.n30 VSUBS 0.031199f
C260 VN.n31 VSUBS 1.00482f
C261 VN.n32 VSUBS 0.034251f
C262 VN.n33 VSUBS 0.030824f
C263 VN.t9 VSUBS 2.65229f
C264 VN.n34 VSUBS 0.028634f
C265 VN.n35 VSUBS 0.030824f
C266 VN.t5 VSUBS 2.65229f
C267 VN.n36 VSUBS 0.054103f
C268 VN.n37 VSUBS 0.030824f
C269 VN.t0 VSUBS 2.65229f
C270 VN.n38 VSUBS 0.059785f
C271 VN.n39 VSUBS 0.030824f
C272 VN.t4 VSUBS 2.65229f
C273 VN.n40 VSUBS 1.00372f
C274 VN.t3 VSUBS 2.8048f
C275 VN.n41 VSUBS 1.00571f
C276 VN.n42 VSUBS 0.229729f
C277 VN.n43 VSUBS 0.04418f
C278 VN.n44 VSUBS 0.054103f
C279 VN.n45 VSUBS 0.032887f
C280 VN.n46 VSUBS 0.030824f
C281 VN.n47 VSUBS 0.030824f
C282 VN.n48 VSUBS 0.030824f
C283 VN.n49 VSUBS 0.959877f
C284 VN.n50 VSUBS 0.059785f
C285 VN.n51 VSUBS 0.032887f
C286 VN.n52 VSUBS 0.030824f
C287 VN.n53 VSUBS 0.030824f
C288 VN.n54 VSUBS 0.030824f
C289 VN.n55 VSUBS 0.04418f
C290 VN.n56 VSUBS 0.930935f
C291 VN.n57 VSUBS 0.041922f
C292 VN.n58 VSUBS 0.056589f
C293 VN.n59 VSUBS 0.030824f
C294 VN.n60 VSUBS 0.030824f
C295 VN.n61 VSUBS 0.030824f
C296 VN.n62 VSUBS 0.061552f
C297 VN.n63 VSUBS 0.031199f
C298 VN.n64 VSUBS 1.00482f
C299 VN.n65 VSUBS 1.83649f
C300 VDD1.n0 VSUBS 0.028824f
C301 VDD1.n1 VSUBS 0.026747f
C302 VDD1.n2 VSUBS 0.014373f
C303 VDD1.n3 VSUBS 0.033971f
C304 VDD1.n4 VSUBS 0.015218f
C305 VDD1.n5 VSUBS 0.026747f
C306 VDD1.n6 VSUBS 0.014795f
C307 VDD1.n7 VSUBS 0.033971f
C308 VDD1.n8 VSUBS 0.014373f
C309 VDD1.n9 VSUBS 0.015218f
C310 VDD1.n10 VSUBS 0.026747f
C311 VDD1.n11 VSUBS 0.014373f
C312 VDD1.n12 VSUBS 0.033971f
C313 VDD1.n13 VSUBS 0.015218f
C314 VDD1.n14 VSUBS 0.026747f
C315 VDD1.n15 VSUBS 0.014373f
C316 VDD1.n16 VSUBS 0.033971f
C317 VDD1.n17 VSUBS 0.015218f
C318 VDD1.n18 VSUBS 0.026747f
C319 VDD1.n19 VSUBS 0.014373f
C320 VDD1.n20 VSUBS 0.033971f
C321 VDD1.n21 VSUBS 0.015218f
C322 VDD1.n22 VSUBS 0.026747f
C323 VDD1.n23 VSUBS 0.014373f
C324 VDD1.n24 VSUBS 0.033971f
C325 VDD1.n25 VSUBS 0.015218f
C326 VDD1.n26 VSUBS 0.026747f
C327 VDD1.n27 VSUBS 0.014373f
C328 VDD1.n28 VSUBS 0.025479f
C329 VDD1.n29 VSUBS 0.021611f
C330 VDD1.t9 VSUBS 0.072803f
C331 VDD1.n30 VSUBS 0.197693f
C332 VDD1.n31 VSUBS 1.84869f
C333 VDD1.n32 VSUBS 0.014373f
C334 VDD1.n33 VSUBS 0.015218f
C335 VDD1.n34 VSUBS 0.033971f
C336 VDD1.n35 VSUBS 0.033971f
C337 VDD1.n36 VSUBS 0.015218f
C338 VDD1.n37 VSUBS 0.014373f
C339 VDD1.n38 VSUBS 0.026747f
C340 VDD1.n39 VSUBS 0.026747f
C341 VDD1.n40 VSUBS 0.014373f
C342 VDD1.n41 VSUBS 0.015218f
C343 VDD1.n42 VSUBS 0.033971f
C344 VDD1.n43 VSUBS 0.033971f
C345 VDD1.n44 VSUBS 0.015218f
C346 VDD1.n45 VSUBS 0.014373f
C347 VDD1.n46 VSUBS 0.026747f
C348 VDD1.n47 VSUBS 0.026747f
C349 VDD1.n48 VSUBS 0.014373f
C350 VDD1.n49 VSUBS 0.015218f
C351 VDD1.n50 VSUBS 0.033971f
C352 VDD1.n51 VSUBS 0.033971f
C353 VDD1.n52 VSUBS 0.015218f
C354 VDD1.n53 VSUBS 0.014373f
C355 VDD1.n54 VSUBS 0.026747f
C356 VDD1.n55 VSUBS 0.026747f
C357 VDD1.n56 VSUBS 0.014373f
C358 VDD1.n57 VSUBS 0.015218f
C359 VDD1.n58 VSUBS 0.033971f
C360 VDD1.n59 VSUBS 0.033971f
C361 VDD1.n60 VSUBS 0.015218f
C362 VDD1.n61 VSUBS 0.014373f
C363 VDD1.n62 VSUBS 0.026747f
C364 VDD1.n63 VSUBS 0.026747f
C365 VDD1.n64 VSUBS 0.014373f
C366 VDD1.n65 VSUBS 0.015218f
C367 VDD1.n66 VSUBS 0.033971f
C368 VDD1.n67 VSUBS 0.033971f
C369 VDD1.n68 VSUBS 0.015218f
C370 VDD1.n69 VSUBS 0.014373f
C371 VDD1.n70 VSUBS 0.026747f
C372 VDD1.n71 VSUBS 0.026747f
C373 VDD1.n72 VSUBS 0.014373f
C374 VDD1.n73 VSUBS 0.015218f
C375 VDD1.n74 VSUBS 0.033971f
C376 VDD1.n75 VSUBS 0.033971f
C377 VDD1.n76 VSUBS 0.033971f
C378 VDD1.n77 VSUBS 0.014795f
C379 VDD1.n78 VSUBS 0.014373f
C380 VDD1.n79 VSUBS 0.026747f
C381 VDD1.n80 VSUBS 0.026747f
C382 VDD1.n81 VSUBS 0.014373f
C383 VDD1.n82 VSUBS 0.015218f
C384 VDD1.n83 VSUBS 0.033971f
C385 VDD1.n84 VSUBS 0.080316f
C386 VDD1.n85 VSUBS 0.015218f
C387 VDD1.n86 VSUBS 0.014373f
C388 VDD1.n87 VSUBS 0.064747f
C389 VDD1.n88 VSUBS 0.067127f
C390 VDD1.t6 VSUBS 0.34156f
C391 VDD1.t5 VSUBS 0.34156f
C392 VDD1.n89 VSUBS 2.8055f
C393 VDD1.n90 VSUBS 0.941922f
C394 VDD1.n91 VSUBS 0.028824f
C395 VDD1.n92 VSUBS 0.026747f
C396 VDD1.n93 VSUBS 0.014373f
C397 VDD1.n94 VSUBS 0.033971f
C398 VDD1.n95 VSUBS 0.015218f
C399 VDD1.n96 VSUBS 0.026747f
C400 VDD1.n97 VSUBS 0.014795f
C401 VDD1.n98 VSUBS 0.033971f
C402 VDD1.n99 VSUBS 0.015218f
C403 VDD1.n100 VSUBS 0.026747f
C404 VDD1.n101 VSUBS 0.014373f
C405 VDD1.n102 VSUBS 0.033971f
C406 VDD1.n103 VSUBS 0.015218f
C407 VDD1.n104 VSUBS 0.026747f
C408 VDD1.n105 VSUBS 0.014373f
C409 VDD1.n106 VSUBS 0.033971f
C410 VDD1.n107 VSUBS 0.015218f
C411 VDD1.n108 VSUBS 0.026747f
C412 VDD1.n109 VSUBS 0.014373f
C413 VDD1.n110 VSUBS 0.033971f
C414 VDD1.n111 VSUBS 0.015218f
C415 VDD1.n112 VSUBS 0.026747f
C416 VDD1.n113 VSUBS 0.014373f
C417 VDD1.n114 VSUBS 0.033971f
C418 VDD1.n115 VSUBS 0.015218f
C419 VDD1.n116 VSUBS 0.026747f
C420 VDD1.n117 VSUBS 0.014373f
C421 VDD1.n118 VSUBS 0.025479f
C422 VDD1.n119 VSUBS 0.021611f
C423 VDD1.t1 VSUBS 0.072803f
C424 VDD1.n120 VSUBS 0.197693f
C425 VDD1.n121 VSUBS 1.84869f
C426 VDD1.n122 VSUBS 0.014373f
C427 VDD1.n123 VSUBS 0.015218f
C428 VDD1.n124 VSUBS 0.033971f
C429 VDD1.n125 VSUBS 0.033971f
C430 VDD1.n126 VSUBS 0.015218f
C431 VDD1.n127 VSUBS 0.014373f
C432 VDD1.n128 VSUBS 0.026747f
C433 VDD1.n129 VSUBS 0.026747f
C434 VDD1.n130 VSUBS 0.014373f
C435 VDD1.n131 VSUBS 0.015218f
C436 VDD1.n132 VSUBS 0.033971f
C437 VDD1.n133 VSUBS 0.033971f
C438 VDD1.n134 VSUBS 0.015218f
C439 VDD1.n135 VSUBS 0.014373f
C440 VDD1.n136 VSUBS 0.026747f
C441 VDD1.n137 VSUBS 0.026747f
C442 VDD1.n138 VSUBS 0.014373f
C443 VDD1.n139 VSUBS 0.015218f
C444 VDD1.n140 VSUBS 0.033971f
C445 VDD1.n141 VSUBS 0.033971f
C446 VDD1.n142 VSUBS 0.015218f
C447 VDD1.n143 VSUBS 0.014373f
C448 VDD1.n144 VSUBS 0.026747f
C449 VDD1.n145 VSUBS 0.026747f
C450 VDD1.n146 VSUBS 0.014373f
C451 VDD1.n147 VSUBS 0.015218f
C452 VDD1.n148 VSUBS 0.033971f
C453 VDD1.n149 VSUBS 0.033971f
C454 VDD1.n150 VSUBS 0.015218f
C455 VDD1.n151 VSUBS 0.014373f
C456 VDD1.n152 VSUBS 0.026747f
C457 VDD1.n153 VSUBS 0.026747f
C458 VDD1.n154 VSUBS 0.014373f
C459 VDD1.n155 VSUBS 0.015218f
C460 VDD1.n156 VSUBS 0.033971f
C461 VDD1.n157 VSUBS 0.033971f
C462 VDD1.n158 VSUBS 0.015218f
C463 VDD1.n159 VSUBS 0.014373f
C464 VDD1.n160 VSUBS 0.026747f
C465 VDD1.n161 VSUBS 0.026747f
C466 VDD1.n162 VSUBS 0.014373f
C467 VDD1.n163 VSUBS 0.014373f
C468 VDD1.n164 VSUBS 0.015218f
C469 VDD1.n165 VSUBS 0.033971f
C470 VDD1.n166 VSUBS 0.033971f
C471 VDD1.n167 VSUBS 0.033971f
C472 VDD1.n168 VSUBS 0.014795f
C473 VDD1.n169 VSUBS 0.014373f
C474 VDD1.n170 VSUBS 0.026747f
C475 VDD1.n171 VSUBS 0.026747f
C476 VDD1.n172 VSUBS 0.014373f
C477 VDD1.n173 VSUBS 0.015218f
C478 VDD1.n174 VSUBS 0.033971f
C479 VDD1.n175 VSUBS 0.080316f
C480 VDD1.n176 VSUBS 0.015218f
C481 VDD1.n177 VSUBS 0.014373f
C482 VDD1.n178 VSUBS 0.064747f
C483 VDD1.n179 VSUBS 0.067127f
C484 VDD1.t4 VSUBS 0.34156f
C485 VDD1.t8 VSUBS 0.34156f
C486 VDD1.n180 VSUBS 2.80549f
C487 VDD1.n181 VSUBS 0.933579f
C488 VDD1.t0 VSUBS 0.34156f
C489 VDD1.t3 VSUBS 0.34156f
C490 VDD1.n182 VSUBS 2.82129f
C491 VDD1.n183 VSUBS 3.42073f
C492 VDD1.t2 VSUBS 0.34156f
C493 VDD1.t7 VSUBS 0.34156f
C494 VDD1.n184 VSUBS 2.80549f
C495 VDD1.n185 VSUBS 3.73394f
C496 VTAIL.t19 VSUBS 0.350025f
C497 VTAIL.t5 VSUBS 0.350025f
C498 VTAIL.n0 VSUBS 2.71637f
C499 VTAIL.n1 VSUBS 0.909329f
C500 VTAIL.n2 VSUBS 0.029538f
C501 VTAIL.n3 VSUBS 0.02741f
C502 VTAIL.n4 VSUBS 0.014729f
C503 VTAIL.n5 VSUBS 0.034813f
C504 VTAIL.n6 VSUBS 0.015595f
C505 VTAIL.n7 VSUBS 0.02741f
C506 VTAIL.n8 VSUBS 0.015162f
C507 VTAIL.n9 VSUBS 0.034813f
C508 VTAIL.n10 VSUBS 0.015595f
C509 VTAIL.n11 VSUBS 0.02741f
C510 VTAIL.n12 VSUBS 0.014729f
C511 VTAIL.n13 VSUBS 0.034813f
C512 VTAIL.n14 VSUBS 0.015595f
C513 VTAIL.n15 VSUBS 0.02741f
C514 VTAIL.n16 VSUBS 0.014729f
C515 VTAIL.n17 VSUBS 0.034813f
C516 VTAIL.n18 VSUBS 0.015595f
C517 VTAIL.n19 VSUBS 0.02741f
C518 VTAIL.n20 VSUBS 0.014729f
C519 VTAIL.n21 VSUBS 0.034813f
C520 VTAIL.n22 VSUBS 0.015595f
C521 VTAIL.n23 VSUBS 0.02741f
C522 VTAIL.n24 VSUBS 0.014729f
C523 VTAIL.n25 VSUBS 0.034813f
C524 VTAIL.n26 VSUBS 0.015595f
C525 VTAIL.n27 VSUBS 0.02741f
C526 VTAIL.n28 VSUBS 0.014729f
C527 VTAIL.n29 VSUBS 0.02611f
C528 VTAIL.n30 VSUBS 0.022147f
C529 VTAIL.t11 VSUBS 0.074608f
C530 VTAIL.n31 VSUBS 0.202592f
C531 VTAIL.n32 VSUBS 1.8945f
C532 VTAIL.n33 VSUBS 0.014729f
C533 VTAIL.n34 VSUBS 0.015595f
C534 VTAIL.n35 VSUBS 0.034813f
C535 VTAIL.n36 VSUBS 0.034813f
C536 VTAIL.n37 VSUBS 0.015595f
C537 VTAIL.n38 VSUBS 0.014729f
C538 VTAIL.n39 VSUBS 0.02741f
C539 VTAIL.n40 VSUBS 0.02741f
C540 VTAIL.n41 VSUBS 0.014729f
C541 VTAIL.n42 VSUBS 0.015595f
C542 VTAIL.n43 VSUBS 0.034813f
C543 VTAIL.n44 VSUBS 0.034813f
C544 VTAIL.n45 VSUBS 0.015595f
C545 VTAIL.n46 VSUBS 0.014729f
C546 VTAIL.n47 VSUBS 0.02741f
C547 VTAIL.n48 VSUBS 0.02741f
C548 VTAIL.n49 VSUBS 0.014729f
C549 VTAIL.n50 VSUBS 0.015595f
C550 VTAIL.n51 VSUBS 0.034813f
C551 VTAIL.n52 VSUBS 0.034813f
C552 VTAIL.n53 VSUBS 0.015595f
C553 VTAIL.n54 VSUBS 0.014729f
C554 VTAIL.n55 VSUBS 0.02741f
C555 VTAIL.n56 VSUBS 0.02741f
C556 VTAIL.n57 VSUBS 0.014729f
C557 VTAIL.n58 VSUBS 0.015595f
C558 VTAIL.n59 VSUBS 0.034813f
C559 VTAIL.n60 VSUBS 0.034813f
C560 VTAIL.n61 VSUBS 0.015595f
C561 VTAIL.n62 VSUBS 0.014729f
C562 VTAIL.n63 VSUBS 0.02741f
C563 VTAIL.n64 VSUBS 0.02741f
C564 VTAIL.n65 VSUBS 0.014729f
C565 VTAIL.n66 VSUBS 0.015595f
C566 VTAIL.n67 VSUBS 0.034813f
C567 VTAIL.n68 VSUBS 0.034813f
C568 VTAIL.n69 VSUBS 0.015595f
C569 VTAIL.n70 VSUBS 0.014729f
C570 VTAIL.n71 VSUBS 0.02741f
C571 VTAIL.n72 VSUBS 0.02741f
C572 VTAIL.n73 VSUBS 0.014729f
C573 VTAIL.n74 VSUBS 0.014729f
C574 VTAIL.n75 VSUBS 0.015595f
C575 VTAIL.n76 VSUBS 0.034813f
C576 VTAIL.n77 VSUBS 0.034813f
C577 VTAIL.n78 VSUBS 0.034813f
C578 VTAIL.n79 VSUBS 0.015162f
C579 VTAIL.n80 VSUBS 0.014729f
C580 VTAIL.n81 VSUBS 0.02741f
C581 VTAIL.n82 VSUBS 0.02741f
C582 VTAIL.n83 VSUBS 0.014729f
C583 VTAIL.n84 VSUBS 0.015595f
C584 VTAIL.n85 VSUBS 0.034813f
C585 VTAIL.n86 VSUBS 0.082306f
C586 VTAIL.n87 VSUBS 0.015595f
C587 VTAIL.n88 VSUBS 0.014729f
C588 VTAIL.n89 VSUBS 0.066352f
C589 VTAIL.n90 VSUBS 0.041393f
C590 VTAIL.n91 VSUBS 0.325847f
C591 VTAIL.t17 VSUBS 0.350025f
C592 VTAIL.t16 VSUBS 0.350025f
C593 VTAIL.n92 VSUBS 2.71637f
C594 VTAIL.n93 VSUBS 0.992319f
C595 VTAIL.t14 VSUBS 0.350025f
C596 VTAIL.t10 VSUBS 0.350025f
C597 VTAIL.n94 VSUBS 2.71637f
C598 VTAIL.n95 VSUBS 2.76787f
C599 VTAIL.t2 VSUBS 0.350025f
C600 VTAIL.t1 VSUBS 0.350025f
C601 VTAIL.n96 VSUBS 2.71639f
C602 VTAIL.n97 VSUBS 2.76785f
C603 VTAIL.t3 VSUBS 0.350025f
C604 VTAIL.t4 VSUBS 0.350025f
C605 VTAIL.n98 VSUBS 2.71639f
C606 VTAIL.n99 VSUBS 0.992303f
C607 VTAIL.n100 VSUBS 0.029538f
C608 VTAIL.n101 VSUBS 0.02741f
C609 VTAIL.n102 VSUBS 0.014729f
C610 VTAIL.n103 VSUBS 0.034813f
C611 VTAIL.n104 VSUBS 0.015595f
C612 VTAIL.n105 VSUBS 0.02741f
C613 VTAIL.n106 VSUBS 0.015162f
C614 VTAIL.n107 VSUBS 0.034813f
C615 VTAIL.n108 VSUBS 0.014729f
C616 VTAIL.n109 VSUBS 0.015595f
C617 VTAIL.n110 VSUBS 0.02741f
C618 VTAIL.n111 VSUBS 0.014729f
C619 VTAIL.n112 VSUBS 0.034813f
C620 VTAIL.n113 VSUBS 0.015595f
C621 VTAIL.n114 VSUBS 0.02741f
C622 VTAIL.n115 VSUBS 0.014729f
C623 VTAIL.n116 VSUBS 0.034813f
C624 VTAIL.n117 VSUBS 0.015595f
C625 VTAIL.n118 VSUBS 0.02741f
C626 VTAIL.n119 VSUBS 0.014729f
C627 VTAIL.n120 VSUBS 0.034813f
C628 VTAIL.n121 VSUBS 0.015595f
C629 VTAIL.n122 VSUBS 0.02741f
C630 VTAIL.n123 VSUBS 0.014729f
C631 VTAIL.n124 VSUBS 0.034813f
C632 VTAIL.n125 VSUBS 0.015595f
C633 VTAIL.n126 VSUBS 0.02741f
C634 VTAIL.n127 VSUBS 0.014729f
C635 VTAIL.n128 VSUBS 0.02611f
C636 VTAIL.n129 VSUBS 0.022147f
C637 VTAIL.t0 VSUBS 0.074608f
C638 VTAIL.n130 VSUBS 0.202592f
C639 VTAIL.n131 VSUBS 1.8945f
C640 VTAIL.n132 VSUBS 0.014729f
C641 VTAIL.n133 VSUBS 0.015595f
C642 VTAIL.n134 VSUBS 0.034813f
C643 VTAIL.n135 VSUBS 0.034813f
C644 VTAIL.n136 VSUBS 0.015595f
C645 VTAIL.n137 VSUBS 0.014729f
C646 VTAIL.n138 VSUBS 0.02741f
C647 VTAIL.n139 VSUBS 0.02741f
C648 VTAIL.n140 VSUBS 0.014729f
C649 VTAIL.n141 VSUBS 0.015595f
C650 VTAIL.n142 VSUBS 0.034813f
C651 VTAIL.n143 VSUBS 0.034813f
C652 VTAIL.n144 VSUBS 0.015595f
C653 VTAIL.n145 VSUBS 0.014729f
C654 VTAIL.n146 VSUBS 0.02741f
C655 VTAIL.n147 VSUBS 0.02741f
C656 VTAIL.n148 VSUBS 0.014729f
C657 VTAIL.n149 VSUBS 0.015595f
C658 VTAIL.n150 VSUBS 0.034813f
C659 VTAIL.n151 VSUBS 0.034813f
C660 VTAIL.n152 VSUBS 0.015595f
C661 VTAIL.n153 VSUBS 0.014729f
C662 VTAIL.n154 VSUBS 0.02741f
C663 VTAIL.n155 VSUBS 0.02741f
C664 VTAIL.n156 VSUBS 0.014729f
C665 VTAIL.n157 VSUBS 0.015595f
C666 VTAIL.n158 VSUBS 0.034813f
C667 VTAIL.n159 VSUBS 0.034813f
C668 VTAIL.n160 VSUBS 0.015595f
C669 VTAIL.n161 VSUBS 0.014729f
C670 VTAIL.n162 VSUBS 0.02741f
C671 VTAIL.n163 VSUBS 0.02741f
C672 VTAIL.n164 VSUBS 0.014729f
C673 VTAIL.n165 VSUBS 0.015595f
C674 VTAIL.n166 VSUBS 0.034813f
C675 VTAIL.n167 VSUBS 0.034813f
C676 VTAIL.n168 VSUBS 0.015595f
C677 VTAIL.n169 VSUBS 0.014729f
C678 VTAIL.n170 VSUBS 0.02741f
C679 VTAIL.n171 VSUBS 0.02741f
C680 VTAIL.n172 VSUBS 0.014729f
C681 VTAIL.n173 VSUBS 0.015595f
C682 VTAIL.n174 VSUBS 0.034813f
C683 VTAIL.n175 VSUBS 0.034813f
C684 VTAIL.n176 VSUBS 0.034813f
C685 VTAIL.n177 VSUBS 0.015162f
C686 VTAIL.n178 VSUBS 0.014729f
C687 VTAIL.n179 VSUBS 0.02741f
C688 VTAIL.n180 VSUBS 0.02741f
C689 VTAIL.n181 VSUBS 0.014729f
C690 VTAIL.n182 VSUBS 0.015595f
C691 VTAIL.n183 VSUBS 0.034813f
C692 VTAIL.n184 VSUBS 0.082306f
C693 VTAIL.n185 VSUBS 0.015595f
C694 VTAIL.n186 VSUBS 0.014729f
C695 VTAIL.n187 VSUBS 0.066352f
C696 VTAIL.n188 VSUBS 0.041393f
C697 VTAIL.n189 VSUBS 0.325847f
C698 VTAIL.t18 VSUBS 0.350025f
C699 VTAIL.t9 VSUBS 0.350025f
C700 VTAIL.n190 VSUBS 2.71639f
C701 VTAIL.n191 VSUBS 0.947381f
C702 VTAIL.t13 VSUBS 0.350025f
C703 VTAIL.t15 VSUBS 0.350025f
C704 VTAIL.n192 VSUBS 2.71639f
C705 VTAIL.n193 VSUBS 0.992303f
C706 VTAIL.n194 VSUBS 0.029538f
C707 VTAIL.n195 VSUBS 0.02741f
C708 VTAIL.n196 VSUBS 0.014729f
C709 VTAIL.n197 VSUBS 0.034813f
C710 VTAIL.n198 VSUBS 0.015595f
C711 VTAIL.n199 VSUBS 0.02741f
C712 VTAIL.n200 VSUBS 0.015162f
C713 VTAIL.n201 VSUBS 0.034813f
C714 VTAIL.n202 VSUBS 0.014729f
C715 VTAIL.n203 VSUBS 0.015595f
C716 VTAIL.n204 VSUBS 0.02741f
C717 VTAIL.n205 VSUBS 0.014729f
C718 VTAIL.n206 VSUBS 0.034813f
C719 VTAIL.n207 VSUBS 0.015595f
C720 VTAIL.n208 VSUBS 0.02741f
C721 VTAIL.n209 VSUBS 0.014729f
C722 VTAIL.n210 VSUBS 0.034813f
C723 VTAIL.n211 VSUBS 0.015595f
C724 VTAIL.n212 VSUBS 0.02741f
C725 VTAIL.n213 VSUBS 0.014729f
C726 VTAIL.n214 VSUBS 0.034813f
C727 VTAIL.n215 VSUBS 0.015595f
C728 VTAIL.n216 VSUBS 0.02741f
C729 VTAIL.n217 VSUBS 0.014729f
C730 VTAIL.n218 VSUBS 0.034813f
C731 VTAIL.n219 VSUBS 0.015595f
C732 VTAIL.n220 VSUBS 0.02741f
C733 VTAIL.n221 VSUBS 0.014729f
C734 VTAIL.n222 VSUBS 0.02611f
C735 VTAIL.n223 VSUBS 0.022147f
C736 VTAIL.t12 VSUBS 0.074608f
C737 VTAIL.n224 VSUBS 0.202592f
C738 VTAIL.n225 VSUBS 1.8945f
C739 VTAIL.n226 VSUBS 0.014729f
C740 VTAIL.n227 VSUBS 0.015595f
C741 VTAIL.n228 VSUBS 0.034813f
C742 VTAIL.n229 VSUBS 0.034813f
C743 VTAIL.n230 VSUBS 0.015595f
C744 VTAIL.n231 VSUBS 0.014729f
C745 VTAIL.n232 VSUBS 0.02741f
C746 VTAIL.n233 VSUBS 0.02741f
C747 VTAIL.n234 VSUBS 0.014729f
C748 VTAIL.n235 VSUBS 0.015595f
C749 VTAIL.n236 VSUBS 0.034813f
C750 VTAIL.n237 VSUBS 0.034813f
C751 VTAIL.n238 VSUBS 0.015595f
C752 VTAIL.n239 VSUBS 0.014729f
C753 VTAIL.n240 VSUBS 0.02741f
C754 VTAIL.n241 VSUBS 0.02741f
C755 VTAIL.n242 VSUBS 0.014729f
C756 VTAIL.n243 VSUBS 0.015595f
C757 VTAIL.n244 VSUBS 0.034813f
C758 VTAIL.n245 VSUBS 0.034813f
C759 VTAIL.n246 VSUBS 0.015595f
C760 VTAIL.n247 VSUBS 0.014729f
C761 VTAIL.n248 VSUBS 0.02741f
C762 VTAIL.n249 VSUBS 0.02741f
C763 VTAIL.n250 VSUBS 0.014729f
C764 VTAIL.n251 VSUBS 0.015595f
C765 VTAIL.n252 VSUBS 0.034813f
C766 VTAIL.n253 VSUBS 0.034813f
C767 VTAIL.n254 VSUBS 0.015595f
C768 VTAIL.n255 VSUBS 0.014729f
C769 VTAIL.n256 VSUBS 0.02741f
C770 VTAIL.n257 VSUBS 0.02741f
C771 VTAIL.n258 VSUBS 0.014729f
C772 VTAIL.n259 VSUBS 0.015595f
C773 VTAIL.n260 VSUBS 0.034813f
C774 VTAIL.n261 VSUBS 0.034813f
C775 VTAIL.n262 VSUBS 0.015595f
C776 VTAIL.n263 VSUBS 0.014729f
C777 VTAIL.n264 VSUBS 0.02741f
C778 VTAIL.n265 VSUBS 0.02741f
C779 VTAIL.n266 VSUBS 0.014729f
C780 VTAIL.n267 VSUBS 0.015595f
C781 VTAIL.n268 VSUBS 0.034813f
C782 VTAIL.n269 VSUBS 0.034813f
C783 VTAIL.n270 VSUBS 0.034813f
C784 VTAIL.n271 VSUBS 0.015162f
C785 VTAIL.n272 VSUBS 0.014729f
C786 VTAIL.n273 VSUBS 0.02741f
C787 VTAIL.n274 VSUBS 0.02741f
C788 VTAIL.n275 VSUBS 0.014729f
C789 VTAIL.n276 VSUBS 0.015595f
C790 VTAIL.n277 VSUBS 0.034813f
C791 VTAIL.n278 VSUBS 0.082306f
C792 VTAIL.n279 VSUBS 0.015595f
C793 VTAIL.n280 VSUBS 0.014729f
C794 VTAIL.n281 VSUBS 0.066352f
C795 VTAIL.n282 VSUBS 0.041393f
C796 VTAIL.n283 VSUBS 1.97349f
C797 VTAIL.n284 VSUBS 0.029538f
C798 VTAIL.n285 VSUBS 0.02741f
C799 VTAIL.n286 VSUBS 0.014729f
C800 VTAIL.n287 VSUBS 0.034813f
C801 VTAIL.n288 VSUBS 0.015595f
C802 VTAIL.n289 VSUBS 0.02741f
C803 VTAIL.n290 VSUBS 0.015162f
C804 VTAIL.n291 VSUBS 0.034813f
C805 VTAIL.n292 VSUBS 0.015595f
C806 VTAIL.n293 VSUBS 0.02741f
C807 VTAIL.n294 VSUBS 0.014729f
C808 VTAIL.n295 VSUBS 0.034813f
C809 VTAIL.n296 VSUBS 0.015595f
C810 VTAIL.n297 VSUBS 0.02741f
C811 VTAIL.n298 VSUBS 0.014729f
C812 VTAIL.n299 VSUBS 0.034813f
C813 VTAIL.n300 VSUBS 0.015595f
C814 VTAIL.n301 VSUBS 0.02741f
C815 VTAIL.n302 VSUBS 0.014729f
C816 VTAIL.n303 VSUBS 0.034813f
C817 VTAIL.n304 VSUBS 0.015595f
C818 VTAIL.n305 VSUBS 0.02741f
C819 VTAIL.n306 VSUBS 0.014729f
C820 VTAIL.n307 VSUBS 0.034813f
C821 VTAIL.n308 VSUBS 0.015595f
C822 VTAIL.n309 VSUBS 0.02741f
C823 VTAIL.n310 VSUBS 0.014729f
C824 VTAIL.n311 VSUBS 0.02611f
C825 VTAIL.n312 VSUBS 0.022147f
C826 VTAIL.t8 VSUBS 0.074608f
C827 VTAIL.n313 VSUBS 0.202592f
C828 VTAIL.n314 VSUBS 1.8945f
C829 VTAIL.n315 VSUBS 0.014729f
C830 VTAIL.n316 VSUBS 0.015595f
C831 VTAIL.n317 VSUBS 0.034813f
C832 VTAIL.n318 VSUBS 0.034813f
C833 VTAIL.n319 VSUBS 0.015595f
C834 VTAIL.n320 VSUBS 0.014729f
C835 VTAIL.n321 VSUBS 0.02741f
C836 VTAIL.n322 VSUBS 0.02741f
C837 VTAIL.n323 VSUBS 0.014729f
C838 VTAIL.n324 VSUBS 0.015595f
C839 VTAIL.n325 VSUBS 0.034813f
C840 VTAIL.n326 VSUBS 0.034813f
C841 VTAIL.n327 VSUBS 0.015595f
C842 VTAIL.n328 VSUBS 0.014729f
C843 VTAIL.n329 VSUBS 0.02741f
C844 VTAIL.n330 VSUBS 0.02741f
C845 VTAIL.n331 VSUBS 0.014729f
C846 VTAIL.n332 VSUBS 0.015595f
C847 VTAIL.n333 VSUBS 0.034813f
C848 VTAIL.n334 VSUBS 0.034813f
C849 VTAIL.n335 VSUBS 0.015595f
C850 VTAIL.n336 VSUBS 0.014729f
C851 VTAIL.n337 VSUBS 0.02741f
C852 VTAIL.n338 VSUBS 0.02741f
C853 VTAIL.n339 VSUBS 0.014729f
C854 VTAIL.n340 VSUBS 0.015595f
C855 VTAIL.n341 VSUBS 0.034813f
C856 VTAIL.n342 VSUBS 0.034813f
C857 VTAIL.n343 VSUBS 0.015595f
C858 VTAIL.n344 VSUBS 0.014729f
C859 VTAIL.n345 VSUBS 0.02741f
C860 VTAIL.n346 VSUBS 0.02741f
C861 VTAIL.n347 VSUBS 0.014729f
C862 VTAIL.n348 VSUBS 0.015595f
C863 VTAIL.n349 VSUBS 0.034813f
C864 VTAIL.n350 VSUBS 0.034813f
C865 VTAIL.n351 VSUBS 0.015595f
C866 VTAIL.n352 VSUBS 0.014729f
C867 VTAIL.n353 VSUBS 0.02741f
C868 VTAIL.n354 VSUBS 0.02741f
C869 VTAIL.n355 VSUBS 0.014729f
C870 VTAIL.n356 VSUBS 0.014729f
C871 VTAIL.n357 VSUBS 0.015595f
C872 VTAIL.n358 VSUBS 0.034813f
C873 VTAIL.n359 VSUBS 0.034813f
C874 VTAIL.n360 VSUBS 0.034813f
C875 VTAIL.n361 VSUBS 0.015162f
C876 VTAIL.n362 VSUBS 0.014729f
C877 VTAIL.n363 VSUBS 0.02741f
C878 VTAIL.n364 VSUBS 0.02741f
C879 VTAIL.n365 VSUBS 0.014729f
C880 VTAIL.n366 VSUBS 0.015595f
C881 VTAIL.n367 VSUBS 0.034813f
C882 VTAIL.n368 VSUBS 0.082306f
C883 VTAIL.n369 VSUBS 0.015595f
C884 VTAIL.n370 VSUBS 0.014729f
C885 VTAIL.n371 VSUBS 0.066352f
C886 VTAIL.n372 VSUBS 0.041393f
C887 VTAIL.n373 VSUBS 1.97349f
C888 VTAIL.t7 VSUBS 0.350025f
C889 VTAIL.t6 VSUBS 0.350025f
C890 VTAIL.n374 VSUBS 2.71637f
C891 VTAIL.n375 VSUBS 0.857555f
C892 VP.n0 VSUBS 0.03136f
C893 VP.t6 VSUBS 2.6984f
C894 VP.n1 VSUBS 0.029132f
C895 VP.n2 VSUBS 0.03136f
C896 VP.t9 VSUBS 2.6984f
C897 VP.n3 VSUBS 0.055044f
C898 VP.n4 VSUBS 0.03136f
C899 VP.t1 VSUBS 2.6984f
C900 VP.n5 VSUBS 0.060824f
C901 VP.n6 VSUBS 0.03136f
C902 VP.t5 VSUBS 2.6984f
C903 VP.n7 VSUBS 0.94712f
C904 VP.n8 VSUBS 0.03136f
C905 VP.n9 VSUBS 0.062622f
C906 VP.n10 VSUBS 0.03136f
C907 VP.t2 VSUBS 2.6984f
C908 VP.n11 VSUBS 0.029132f
C909 VP.n12 VSUBS 0.03136f
C910 VP.t7 VSUBS 2.6984f
C911 VP.n13 VSUBS 0.055044f
C912 VP.n14 VSUBS 0.03136f
C913 VP.t4 VSUBS 2.6984f
C914 VP.n15 VSUBS 0.060824f
C915 VP.n16 VSUBS 0.03136f
C916 VP.t3 VSUBS 2.6984f
C917 VP.n17 VSUBS 1.02117f
C918 VP.t0 VSUBS 2.85357f
C919 VP.n18 VSUBS 1.02319f
C920 VP.n19 VSUBS 0.233723f
C921 VP.n20 VSUBS 0.044948f
C922 VP.n21 VSUBS 0.055044f
C923 VP.n22 VSUBS 0.033459f
C924 VP.n23 VSUBS 0.03136f
C925 VP.n24 VSUBS 0.03136f
C926 VP.n25 VSUBS 0.03136f
C927 VP.n26 VSUBS 0.976565f
C928 VP.n27 VSUBS 0.060824f
C929 VP.n28 VSUBS 0.033459f
C930 VP.n29 VSUBS 0.03136f
C931 VP.n30 VSUBS 0.03136f
C932 VP.n31 VSUBS 0.03136f
C933 VP.n32 VSUBS 0.044948f
C934 VP.n33 VSUBS 0.94712f
C935 VP.n34 VSUBS 0.042651f
C936 VP.n35 VSUBS 0.057573f
C937 VP.n36 VSUBS 0.03136f
C938 VP.n37 VSUBS 0.03136f
C939 VP.n38 VSUBS 0.03136f
C940 VP.n39 VSUBS 0.062622f
C941 VP.n40 VSUBS 0.031742f
C942 VP.n41 VSUBS 1.02229f
C943 VP.n42 VSUBS 1.84808f
C944 VP.n43 VSUBS 1.86958f
C945 VP.t8 VSUBS 2.6984f
C946 VP.n44 VSUBS 1.02229f
C947 VP.n45 VSUBS 0.031742f
C948 VP.n46 VSUBS 0.03136f
C949 VP.n47 VSUBS 0.03136f
C950 VP.n48 VSUBS 0.03136f
C951 VP.n49 VSUBS 0.029132f
C952 VP.n50 VSUBS 0.057573f
C953 VP.n51 VSUBS 0.042651f
C954 VP.n52 VSUBS 0.03136f
C955 VP.n53 VSUBS 0.03136f
C956 VP.n54 VSUBS 0.044948f
C957 VP.n55 VSUBS 0.055044f
C958 VP.n56 VSUBS 0.033459f
C959 VP.n57 VSUBS 0.03136f
C960 VP.n58 VSUBS 0.03136f
C961 VP.n59 VSUBS 0.03136f
C962 VP.n60 VSUBS 0.976565f
C963 VP.n61 VSUBS 0.060824f
C964 VP.n62 VSUBS 0.033459f
C965 VP.n63 VSUBS 0.03136f
C966 VP.n64 VSUBS 0.03136f
C967 VP.n65 VSUBS 0.03136f
C968 VP.n66 VSUBS 0.044948f
C969 VP.n67 VSUBS 0.94712f
C970 VP.n68 VSUBS 0.042651f
C971 VP.n69 VSUBS 0.057573f
C972 VP.n70 VSUBS 0.03136f
C973 VP.n71 VSUBS 0.03136f
C974 VP.n72 VSUBS 0.03136f
C975 VP.n73 VSUBS 0.062622f
C976 VP.n74 VSUBS 0.031742f
C977 VP.n75 VSUBS 1.02229f
C978 VP.n76 VSUBS 0.034846f
C979 B.n0 VSUBS 0.00507f
C980 B.n1 VSUBS 0.00507f
C981 B.n2 VSUBS 0.008018f
C982 B.n3 VSUBS 0.008018f
C983 B.n4 VSUBS 0.008018f
C984 B.n5 VSUBS 0.008018f
C985 B.n6 VSUBS 0.008018f
C986 B.n7 VSUBS 0.008018f
C987 B.n8 VSUBS 0.008018f
C988 B.n9 VSUBS 0.008018f
C989 B.n10 VSUBS 0.008018f
C990 B.n11 VSUBS 0.008018f
C991 B.n12 VSUBS 0.008018f
C992 B.n13 VSUBS 0.008018f
C993 B.n14 VSUBS 0.008018f
C994 B.n15 VSUBS 0.008018f
C995 B.n16 VSUBS 0.008018f
C996 B.n17 VSUBS 0.008018f
C997 B.n18 VSUBS 0.008018f
C998 B.n19 VSUBS 0.008018f
C999 B.n20 VSUBS 0.008018f
C1000 B.n21 VSUBS 0.008018f
C1001 B.n22 VSUBS 0.008018f
C1002 B.n23 VSUBS 0.008018f
C1003 B.n24 VSUBS 0.008018f
C1004 B.n25 VSUBS 0.008018f
C1005 B.n26 VSUBS 0.02036f
C1006 B.n27 VSUBS 0.008018f
C1007 B.n28 VSUBS 0.008018f
C1008 B.n29 VSUBS 0.008018f
C1009 B.n30 VSUBS 0.008018f
C1010 B.n31 VSUBS 0.008018f
C1011 B.n32 VSUBS 0.008018f
C1012 B.n33 VSUBS 0.008018f
C1013 B.n34 VSUBS 0.008018f
C1014 B.n35 VSUBS 0.008018f
C1015 B.n36 VSUBS 0.008018f
C1016 B.n37 VSUBS 0.008018f
C1017 B.n38 VSUBS 0.008018f
C1018 B.n39 VSUBS 0.008018f
C1019 B.n40 VSUBS 0.008018f
C1020 B.n41 VSUBS 0.008018f
C1021 B.n42 VSUBS 0.008018f
C1022 B.n43 VSUBS 0.008018f
C1023 B.n44 VSUBS 0.008018f
C1024 B.n45 VSUBS 0.008018f
C1025 B.n46 VSUBS 0.008018f
C1026 B.n47 VSUBS 0.008018f
C1027 B.n48 VSUBS 0.008018f
C1028 B.n49 VSUBS 0.008018f
C1029 B.n50 VSUBS 0.008018f
C1030 B.n51 VSUBS 0.008018f
C1031 B.n52 VSUBS 0.008018f
C1032 B.n53 VSUBS 0.008018f
C1033 B.t2 VSUBS 0.351633f
C1034 B.t1 VSUBS 0.381564f
C1035 B.t0 VSUBS 1.56953f
C1036 B.n54 VSUBS 0.56787f
C1037 B.n55 VSUBS 0.347703f
C1038 B.n56 VSUBS 0.008018f
C1039 B.n57 VSUBS 0.008018f
C1040 B.n58 VSUBS 0.008018f
C1041 B.n59 VSUBS 0.008018f
C1042 B.t8 VSUBS 0.351637f
C1043 B.t7 VSUBS 0.381568f
C1044 B.t6 VSUBS 1.56953f
C1045 B.n60 VSUBS 0.567867f
C1046 B.n61 VSUBS 0.347699f
C1047 B.n62 VSUBS 0.008018f
C1048 B.n63 VSUBS 0.008018f
C1049 B.n64 VSUBS 0.008018f
C1050 B.n65 VSUBS 0.008018f
C1051 B.n66 VSUBS 0.008018f
C1052 B.n67 VSUBS 0.008018f
C1053 B.n68 VSUBS 0.008018f
C1054 B.n69 VSUBS 0.008018f
C1055 B.n70 VSUBS 0.008018f
C1056 B.n71 VSUBS 0.008018f
C1057 B.n72 VSUBS 0.008018f
C1058 B.n73 VSUBS 0.008018f
C1059 B.n74 VSUBS 0.008018f
C1060 B.n75 VSUBS 0.008018f
C1061 B.n76 VSUBS 0.008018f
C1062 B.n77 VSUBS 0.008018f
C1063 B.n78 VSUBS 0.008018f
C1064 B.n79 VSUBS 0.008018f
C1065 B.n80 VSUBS 0.008018f
C1066 B.n81 VSUBS 0.008018f
C1067 B.n82 VSUBS 0.008018f
C1068 B.n83 VSUBS 0.008018f
C1069 B.n84 VSUBS 0.008018f
C1070 B.n85 VSUBS 0.008018f
C1071 B.n86 VSUBS 0.008018f
C1072 B.n87 VSUBS 0.008018f
C1073 B.n88 VSUBS 0.019495f
C1074 B.n89 VSUBS 0.008018f
C1075 B.n90 VSUBS 0.008018f
C1076 B.n91 VSUBS 0.008018f
C1077 B.n92 VSUBS 0.008018f
C1078 B.n93 VSUBS 0.008018f
C1079 B.n94 VSUBS 0.008018f
C1080 B.n95 VSUBS 0.008018f
C1081 B.n96 VSUBS 0.008018f
C1082 B.n97 VSUBS 0.008018f
C1083 B.n98 VSUBS 0.008018f
C1084 B.n99 VSUBS 0.008018f
C1085 B.n100 VSUBS 0.008018f
C1086 B.n101 VSUBS 0.008018f
C1087 B.n102 VSUBS 0.008018f
C1088 B.n103 VSUBS 0.008018f
C1089 B.n104 VSUBS 0.008018f
C1090 B.n105 VSUBS 0.008018f
C1091 B.n106 VSUBS 0.008018f
C1092 B.n107 VSUBS 0.008018f
C1093 B.n108 VSUBS 0.008018f
C1094 B.n109 VSUBS 0.008018f
C1095 B.n110 VSUBS 0.008018f
C1096 B.n111 VSUBS 0.008018f
C1097 B.n112 VSUBS 0.008018f
C1098 B.n113 VSUBS 0.008018f
C1099 B.n114 VSUBS 0.008018f
C1100 B.n115 VSUBS 0.008018f
C1101 B.n116 VSUBS 0.008018f
C1102 B.n117 VSUBS 0.008018f
C1103 B.n118 VSUBS 0.008018f
C1104 B.n119 VSUBS 0.008018f
C1105 B.n120 VSUBS 0.008018f
C1106 B.n121 VSUBS 0.008018f
C1107 B.n122 VSUBS 0.008018f
C1108 B.n123 VSUBS 0.008018f
C1109 B.n124 VSUBS 0.008018f
C1110 B.n125 VSUBS 0.008018f
C1111 B.n126 VSUBS 0.008018f
C1112 B.n127 VSUBS 0.008018f
C1113 B.n128 VSUBS 0.008018f
C1114 B.n129 VSUBS 0.008018f
C1115 B.n130 VSUBS 0.008018f
C1116 B.n131 VSUBS 0.008018f
C1117 B.n132 VSUBS 0.008018f
C1118 B.n133 VSUBS 0.008018f
C1119 B.n134 VSUBS 0.008018f
C1120 B.n135 VSUBS 0.008018f
C1121 B.n136 VSUBS 0.008018f
C1122 B.n137 VSUBS 0.02036f
C1123 B.n138 VSUBS 0.008018f
C1124 B.n139 VSUBS 0.008018f
C1125 B.n140 VSUBS 0.008018f
C1126 B.n141 VSUBS 0.008018f
C1127 B.n142 VSUBS 0.008018f
C1128 B.n143 VSUBS 0.008018f
C1129 B.n144 VSUBS 0.008018f
C1130 B.n145 VSUBS 0.008018f
C1131 B.n146 VSUBS 0.008018f
C1132 B.n147 VSUBS 0.008018f
C1133 B.n148 VSUBS 0.008018f
C1134 B.n149 VSUBS 0.008018f
C1135 B.n150 VSUBS 0.008018f
C1136 B.n151 VSUBS 0.008018f
C1137 B.n152 VSUBS 0.008018f
C1138 B.n153 VSUBS 0.008018f
C1139 B.n154 VSUBS 0.008018f
C1140 B.n155 VSUBS 0.008018f
C1141 B.n156 VSUBS 0.008018f
C1142 B.n157 VSUBS 0.008018f
C1143 B.n158 VSUBS 0.008018f
C1144 B.n159 VSUBS 0.008018f
C1145 B.n160 VSUBS 0.008018f
C1146 B.n161 VSUBS 0.008018f
C1147 B.n162 VSUBS 0.008018f
C1148 B.n163 VSUBS 0.008018f
C1149 B.t10 VSUBS 0.351637f
C1150 B.t11 VSUBS 0.381568f
C1151 B.t9 VSUBS 1.56953f
C1152 B.n164 VSUBS 0.567867f
C1153 B.n165 VSUBS 0.347699f
C1154 B.n166 VSUBS 0.018577f
C1155 B.n167 VSUBS 0.008018f
C1156 B.n168 VSUBS 0.008018f
C1157 B.n169 VSUBS 0.008018f
C1158 B.n170 VSUBS 0.008018f
C1159 B.n171 VSUBS 0.008018f
C1160 B.t4 VSUBS 0.351633f
C1161 B.t5 VSUBS 0.381564f
C1162 B.t3 VSUBS 1.56953f
C1163 B.n172 VSUBS 0.56787f
C1164 B.n173 VSUBS 0.347703f
C1165 B.n174 VSUBS 0.008018f
C1166 B.n175 VSUBS 0.008018f
C1167 B.n176 VSUBS 0.008018f
C1168 B.n177 VSUBS 0.008018f
C1169 B.n178 VSUBS 0.008018f
C1170 B.n179 VSUBS 0.008018f
C1171 B.n180 VSUBS 0.008018f
C1172 B.n181 VSUBS 0.008018f
C1173 B.n182 VSUBS 0.008018f
C1174 B.n183 VSUBS 0.008018f
C1175 B.n184 VSUBS 0.008018f
C1176 B.n185 VSUBS 0.008018f
C1177 B.n186 VSUBS 0.008018f
C1178 B.n187 VSUBS 0.008018f
C1179 B.n188 VSUBS 0.008018f
C1180 B.n189 VSUBS 0.008018f
C1181 B.n190 VSUBS 0.008018f
C1182 B.n191 VSUBS 0.008018f
C1183 B.n192 VSUBS 0.008018f
C1184 B.n193 VSUBS 0.008018f
C1185 B.n194 VSUBS 0.008018f
C1186 B.n195 VSUBS 0.008018f
C1187 B.n196 VSUBS 0.008018f
C1188 B.n197 VSUBS 0.008018f
C1189 B.n198 VSUBS 0.008018f
C1190 B.n199 VSUBS 0.008018f
C1191 B.n200 VSUBS 0.019495f
C1192 B.n201 VSUBS 0.008018f
C1193 B.n202 VSUBS 0.008018f
C1194 B.n203 VSUBS 0.008018f
C1195 B.n204 VSUBS 0.008018f
C1196 B.n205 VSUBS 0.008018f
C1197 B.n206 VSUBS 0.008018f
C1198 B.n207 VSUBS 0.008018f
C1199 B.n208 VSUBS 0.008018f
C1200 B.n209 VSUBS 0.008018f
C1201 B.n210 VSUBS 0.008018f
C1202 B.n211 VSUBS 0.008018f
C1203 B.n212 VSUBS 0.008018f
C1204 B.n213 VSUBS 0.008018f
C1205 B.n214 VSUBS 0.008018f
C1206 B.n215 VSUBS 0.008018f
C1207 B.n216 VSUBS 0.008018f
C1208 B.n217 VSUBS 0.008018f
C1209 B.n218 VSUBS 0.008018f
C1210 B.n219 VSUBS 0.008018f
C1211 B.n220 VSUBS 0.008018f
C1212 B.n221 VSUBS 0.008018f
C1213 B.n222 VSUBS 0.008018f
C1214 B.n223 VSUBS 0.008018f
C1215 B.n224 VSUBS 0.008018f
C1216 B.n225 VSUBS 0.008018f
C1217 B.n226 VSUBS 0.008018f
C1218 B.n227 VSUBS 0.008018f
C1219 B.n228 VSUBS 0.008018f
C1220 B.n229 VSUBS 0.008018f
C1221 B.n230 VSUBS 0.008018f
C1222 B.n231 VSUBS 0.008018f
C1223 B.n232 VSUBS 0.008018f
C1224 B.n233 VSUBS 0.008018f
C1225 B.n234 VSUBS 0.008018f
C1226 B.n235 VSUBS 0.008018f
C1227 B.n236 VSUBS 0.008018f
C1228 B.n237 VSUBS 0.008018f
C1229 B.n238 VSUBS 0.008018f
C1230 B.n239 VSUBS 0.008018f
C1231 B.n240 VSUBS 0.008018f
C1232 B.n241 VSUBS 0.008018f
C1233 B.n242 VSUBS 0.008018f
C1234 B.n243 VSUBS 0.008018f
C1235 B.n244 VSUBS 0.008018f
C1236 B.n245 VSUBS 0.008018f
C1237 B.n246 VSUBS 0.008018f
C1238 B.n247 VSUBS 0.008018f
C1239 B.n248 VSUBS 0.008018f
C1240 B.n249 VSUBS 0.008018f
C1241 B.n250 VSUBS 0.008018f
C1242 B.n251 VSUBS 0.008018f
C1243 B.n252 VSUBS 0.008018f
C1244 B.n253 VSUBS 0.008018f
C1245 B.n254 VSUBS 0.008018f
C1246 B.n255 VSUBS 0.008018f
C1247 B.n256 VSUBS 0.008018f
C1248 B.n257 VSUBS 0.008018f
C1249 B.n258 VSUBS 0.008018f
C1250 B.n259 VSUBS 0.008018f
C1251 B.n260 VSUBS 0.008018f
C1252 B.n261 VSUBS 0.008018f
C1253 B.n262 VSUBS 0.008018f
C1254 B.n263 VSUBS 0.008018f
C1255 B.n264 VSUBS 0.008018f
C1256 B.n265 VSUBS 0.008018f
C1257 B.n266 VSUBS 0.008018f
C1258 B.n267 VSUBS 0.008018f
C1259 B.n268 VSUBS 0.008018f
C1260 B.n269 VSUBS 0.008018f
C1261 B.n270 VSUBS 0.008018f
C1262 B.n271 VSUBS 0.008018f
C1263 B.n272 VSUBS 0.008018f
C1264 B.n273 VSUBS 0.008018f
C1265 B.n274 VSUBS 0.008018f
C1266 B.n275 VSUBS 0.008018f
C1267 B.n276 VSUBS 0.008018f
C1268 B.n277 VSUBS 0.008018f
C1269 B.n278 VSUBS 0.008018f
C1270 B.n279 VSUBS 0.008018f
C1271 B.n280 VSUBS 0.008018f
C1272 B.n281 VSUBS 0.008018f
C1273 B.n282 VSUBS 0.008018f
C1274 B.n283 VSUBS 0.008018f
C1275 B.n284 VSUBS 0.008018f
C1276 B.n285 VSUBS 0.008018f
C1277 B.n286 VSUBS 0.008018f
C1278 B.n287 VSUBS 0.008018f
C1279 B.n288 VSUBS 0.008018f
C1280 B.n289 VSUBS 0.008018f
C1281 B.n290 VSUBS 0.008018f
C1282 B.n291 VSUBS 0.008018f
C1283 B.n292 VSUBS 0.008018f
C1284 B.n293 VSUBS 0.019495f
C1285 B.n294 VSUBS 0.02036f
C1286 B.n295 VSUBS 0.02036f
C1287 B.n296 VSUBS 0.008018f
C1288 B.n297 VSUBS 0.008018f
C1289 B.n298 VSUBS 0.008018f
C1290 B.n299 VSUBS 0.008018f
C1291 B.n300 VSUBS 0.008018f
C1292 B.n301 VSUBS 0.008018f
C1293 B.n302 VSUBS 0.008018f
C1294 B.n303 VSUBS 0.008018f
C1295 B.n304 VSUBS 0.008018f
C1296 B.n305 VSUBS 0.008018f
C1297 B.n306 VSUBS 0.008018f
C1298 B.n307 VSUBS 0.008018f
C1299 B.n308 VSUBS 0.008018f
C1300 B.n309 VSUBS 0.008018f
C1301 B.n310 VSUBS 0.008018f
C1302 B.n311 VSUBS 0.008018f
C1303 B.n312 VSUBS 0.008018f
C1304 B.n313 VSUBS 0.008018f
C1305 B.n314 VSUBS 0.008018f
C1306 B.n315 VSUBS 0.008018f
C1307 B.n316 VSUBS 0.008018f
C1308 B.n317 VSUBS 0.008018f
C1309 B.n318 VSUBS 0.008018f
C1310 B.n319 VSUBS 0.008018f
C1311 B.n320 VSUBS 0.008018f
C1312 B.n321 VSUBS 0.008018f
C1313 B.n322 VSUBS 0.008018f
C1314 B.n323 VSUBS 0.008018f
C1315 B.n324 VSUBS 0.008018f
C1316 B.n325 VSUBS 0.008018f
C1317 B.n326 VSUBS 0.008018f
C1318 B.n327 VSUBS 0.008018f
C1319 B.n328 VSUBS 0.008018f
C1320 B.n329 VSUBS 0.008018f
C1321 B.n330 VSUBS 0.008018f
C1322 B.n331 VSUBS 0.008018f
C1323 B.n332 VSUBS 0.008018f
C1324 B.n333 VSUBS 0.008018f
C1325 B.n334 VSUBS 0.008018f
C1326 B.n335 VSUBS 0.008018f
C1327 B.n336 VSUBS 0.008018f
C1328 B.n337 VSUBS 0.008018f
C1329 B.n338 VSUBS 0.008018f
C1330 B.n339 VSUBS 0.008018f
C1331 B.n340 VSUBS 0.008018f
C1332 B.n341 VSUBS 0.008018f
C1333 B.n342 VSUBS 0.008018f
C1334 B.n343 VSUBS 0.008018f
C1335 B.n344 VSUBS 0.008018f
C1336 B.n345 VSUBS 0.008018f
C1337 B.n346 VSUBS 0.008018f
C1338 B.n347 VSUBS 0.008018f
C1339 B.n348 VSUBS 0.008018f
C1340 B.n349 VSUBS 0.008018f
C1341 B.n350 VSUBS 0.008018f
C1342 B.n351 VSUBS 0.008018f
C1343 B.n352 VSUBS 0.008018f
C1344 B.n353 VSUBS 0.008018f
C1345 B.n354 VSUBS 0.008018f
C1346 B.n355 VSUBS 0.008018f
C1347 B.n356 VSUBS 0.008018f
C1348 B.n357 VSUBS 0.008018f
C1349 B.n358 VSUBS 0.008018f
C1350 B.n359 VSUBS 0.008018f
C1351 B.n360 VSUBS 0.008018f
C1352 B.n361 VSUBS 0.008018f
C1353 B.n362 VSUBS 0.008018f
C1354 B.n363 VSUBS 0.008018f
C1355 B.n364 VSUBS 0.008018f
C1356 B.n365 VSUBS 0.008018f
C1357 B.n366 VSUBS 0.008018f
C1358 B.n367 VSUBS 0.008018f
C1359 B.n368 VSUBS 0.008018f
C1360 B.n369 VSUBS 0.008018f
C1361 B.n370 VSUBS 0.008018f
C1362 B.n371 VSUBS 0.008018f
C1363 B.n372 VSUBS 0.008018f
C1364 B.n373 VSUBS 0.008018f
C1365 B.n374 VSUBS 0.005542f
C1366 B.n375 VSUBS 0.018577f
C1367 B.n376 VSUBS 0.006485f
C1368 B.n377 VSUBS 0.008018f
C1369 B.n378 VSUBS 0.008018f
C1370 B.n379 VSUBS 0.008018f
C1371 B.n380 VSUBS 0.008018f
C1372 B.n381 VSUBS 0.008018f
C1373 B.n382 VSUBS 0.008018f
C1374 B.n383 VSUBS 0.008018f
C1375 B.n384 VSUBS 0.008018f
C1376 B.n385 VSUBS 0.008018f
C1377 B.n386 VSUBS 0.008018f
C1378 B.n387 VSUBS 0.008018f
C1379 B.n388 VSUBS 0.006485f
C1380 B.n389 VSUBS 0.008018f
C1381 B.n390 VSUBS 0.008018f
C1382 B.n391 VSUBS 0.005542f
C1383 B.n392 VSUBS 0.008018f
C1384 B.n393 VSUBS 0.008018f
C1385 B.n394 VSUBS 0.008018f
C1386 B.n395 VSUBS 0.008018f
C1387 B.n396 VSUBS 0.008018f
C1388 B.n397 VSUBS 0.008018f
C1389 B.n398 VSUBS 0.008018f
C1390 B.n399 VSUBS 0.008018f
C1391 B.n400 VSUBS 0.008018f
C1392 B.n401 VSUBS 0.008018f
C1393 B.n402 VSUBS 0.008018f
C1394 B.n403 VSUBS 0.008018f
C1395 B.n404 VSUBS 0.008018f
C1396 B.n405 VSUBS 0.008018f
C1397 B.n406 VSUBS 0.008018f
C1398 B.n407 VSUBS 0.008018f
C1399 B.n408 VSUBS 0.008018f
C1400 B.n409 VSUBS 0.008018f
C1401 B.n410 VSUBS 0.008018f
C1402 B.n411 VSUBS 0.008018f
C1403 B.n412 VSUBS 0.008018f
C1404 B.n413 VSUBS 0.008018f
C1405 B.n414 VSUBS 0.008018f
C1406 B.n415 VSUBS 0.008018f
C1407 B.n416 VSUBS 0.008018f
C1408 B.n417 VSUBS 0.008018f
C1409 B.n418 VSUBS 0.008018f
C1410 B.n419 VSUBS 0.008018f
C1411 B.n420 VSUBS 0.008018f
C1412 B.n421 VSUBS 0.008018f
C1413 B.n422 VSUBS 0.008018f
C1414 B.n423 VSUBS 0.008018f
C1415 B.n424 VSUBS 0.008018f
C1416 B.n425 VSUBS 0.008018f
C1417 B.n426 VSUBS 0.008018f
C1418 B.n427 VSUBS 0.008018f
C1419 B.n428 VSUBS 0.008018f
C1420 B.n429 VSUBS 0.008018f
C1421 B.n430 VSUBS 0.008018f
C1422 B.n431 VSUBS 0.008018f
C1423 B.n432 VSUBS 0.008018f
C1424 B.n433 VSUBS 0.008018f
C1425 B.n434 VSUBS 0.008018f
C1426 B.n435 VSUBS 0.008018f
C1427 B.n436 VSUBS 0.008018f
C1428 B.n437 VSUBS 0.008018f
C1429 B.n438 VSUBS 0.008018f
C1430 B.n439 VSUBS 0.008018f
C1431 B.n440 VSUBS 0.008018f
C1432 B.n441 VSUBS 0.008018f
C1433 B.n442 VSUBS 0.008018f
C1434 B.n443 VSUBS 0.008018f
C1435 B.n444 VSUBS 0.008018f
C1436 B.n445 VSUBS 0.008018f
C1437 B.n446 VSUBS 0.008018f
C1438 B.n447 VSUBS 0.008018f
C1439 B.n448 VSUBS 0.008018f
C1440 B.n449 VSUBS 0.008018f
C1441 B.n450 VSUBS 0.008018f
C1442 B.n451 VSUBS 0.008018f
C1443 B.n452 VSUBS 0.008018f
C1444 B.n453 VSUBS 0.008018f
C1445 B.n454 VSUBS 0.008018f
C1446 B.n455 VSUBS 0.008018f
C1447 B.n456 VSUBS 0.008018f
C1448 B.n457 VSUBS 0.008018f
C1449 B.n458 VSUBS 0.008018f
C1450 B.n459 VSUBS 0.008018f
C1451 B.n460 VSUBS 0.008018f
C1452 B.n461 VSUBS 0.008018f
C1453 B.n462 VSUBS 0.008018f
C1454 B.n463 VSUBS 0.008018f
C1455 B.n464 VSUBS 0.008018f
C1456 B.n465 VSUBS 0.008018f
C1457 B.n466 VSUBS 0.008018f
C1458 B.n467 VSUBS 0.008018f
C1459 B.n468 VSUBS 0.008018f
C1460 B.n469 VSUBS 0.008018f
C1461 B.n470 VSUBS 0.02036f
C1462 B.n471 VSUBS 0.019495f
C1463 B.n472 VSUBS 0.019495f
C1464 B.n473 VSUBS 0.008018f
C1465 B.n474 VSUBS 0.008018f
C1466 B.n475 VSUBS 0.008018f
C1467 B.n476 VSUBS 0.008018f
C1468 B.n477 VSUBS 0.008018f
C1469 B.n478 VSUBS 0.008018f
C1470 B.n479 VSUBS 0.008018f
C1471 B.n480 VSUBS 0.008018f
C1472 B.n481 VSUBS 0.008018f
C1473 B.n482 VSUBS 0.008018f
C1474 B.n483 VSUBS 0.008018f
C1475 B.n484 VSUBS 0.008018f
C1476 B.n485 VSUBS 0.008018f
C1477 B.n486 VSUBS 0.008018f
C1478 B.n487 VSUBS 0.008018f
C1479 B.n488 VSUBS 0.008018f
C1480 B.n489 VSUBS 0.008018f
C1481 B.n490 VSUBS 0.008018f
C1482 B.n491 VSUBS 0.008018f
C1483 B.n492 VSUBS 0.008018f
C1484 B.n493 VSUBS 0.008018f
C1485 B.n494 VSUBS 0.008018f
C1486 B.n495 VSUBS 0.008018f
C1487 B.n496 VSUBS 0.008018f
C1488 B.n497 VSUBS 0.008018f
C1489 B.n498 VSUBS 0.008018f
C1490 B.n499 VSUBS 0.008018f
C1491 B.n500 VSUBS 0.008018f
C1492 B.n501 VSUBS 0.008018f
C1493 B.n502 VSUBS 0.008018f
C1494 B.n503 VSUBS 0.008018f
C1495 B.n504 VSUBS 0.008018f
C1496 B.n505 VSUBS 0.008018f
C1497 B.n506 VSUBS 0.008018f
C1498 B.n507 VSUBS 0.008018f
C1499 B.n508 VSUBS 0.008018f
C1500 B.n509 VSUBS 0.008018f
C1501 B.n510 VSUBS 0.008018f
C1502 B.n511 VSUBS 0.008018f
C1503 B.n512 VSUBS 0.008018f
C1504 B.n513 VSUBS 0.008018f
C1505 B.n514 VSUBS 0.008018f
C1506 B.n515 VSUBS 0.008018f
C1507 B.n516 VSUBS 0.008018f
C1508 B.n517 VSUBS 0.008018f
C1509 B.n518 VSUBS 0.008018f
C1510 B.n519 VSUBS 0.008018f
C1511 B.n520 VSUBS 0.008018f
C1512 B.n521 VSUBS 0.008018f
C1513 B.n522 VSUBS 0.008018f
C1514 B.n523 VSUBS 0.008018f
C1515 B.n524 VSUBS 0.008018f
C1516 B.n525 VSUBS 0.008018f
C1517 B.n526 VSUBS 0.008018f
C1518 B.n527 VSUBS 0.008018f
C1519 B.n528 VSUBS 0.008018f
C1520 B.n529 VSUBS 0.008018f
C1521 B.n530 VSUBS 0.008018f
C1522 B.n531 VSUBS 0.008018f
C1523 B.n532 VSUBS 0.008018f
C1524 B.n533 VSUBS 0.008018f
C1525 B.n534 VSUBS 0.008018f
C1526 B.n535 VSUBS 0.008018f
C1527 B.n536 VSUBS 0.008018f
C1528 B.n537 VSUBS 0.008018f
C1529 B.n538 VSUBS 0.008018f
C1530 B.n539 VSUBS 0.008018f
C1531 B.n540 VSUBS 0.008018f
C1532 B.n541 VSUBS 0.008018f
C1533 B.n542 VSUBS 0.008018f
C1534 B.n543 VSUBS 0.008018f
C1535 B.n544 VSUBS 0.008018f
C1536 B.n545 VSUBS 0.008018f
C1537 B.n546 VSUBS 0.008018f
C1538 B.n547 VSUBS 0.008018f
C1539 B.n548 VSUBS 0.008018f
C1540 B.n549 VSUBS 0.008018f
C1541 B.n550 VSUBS 0.008018f
C1542 B.n551 VSUBS 0.008018f
C1543 B.n552 VSUBS 0.008018f
C1544 B.n553 VSUBS 0.008018f
C1545 B.n554 VSUBS 0.008018f
C1546 B.n555 VSUBS 0.008018f
C1547 B.n556 VSUBS 0.008018f
C1548 B.n557 VSUBS 0.008018f
C1549 B.n558 VSUBS 0.008018f
C1550 B.n559 VSUBS 0.008018f
C1551 B.n560 VSUBS 0.008018f
C1552 B.n561 VSUBS 0.008018f
C1553 B.n562 VSUBS 0.008018f
C1554 B.n563 VSUBS 0.008018f
C1555 B.n564 VSUBS 0.008018f
C1556 B.n565 VSUBS 0.008018f
C1557 B.n566 VSUBS 0.008018f
C1558 B.n567 VSUBS 0.008018f
C1559 B.n568 VSUBS 0.008018f
C1560 B.n569 VSUBS 0.008018f
C1561 B.n570 VSUBS 0.008018f
C1562 B.n571 VSUBS 0.008018f
C1563 B.n572 VSUBS 0.008018f
C1564 B.n573 VSUBS 0.008018f
C1565 B.n574 VSUBS 0.008018f
C1566 B.n575 VSUBS 0.008018f
C1567 B.n576 VSUBS 0.008018f
C1568 B.n577 VSUBS 0.008018f
C1569 B.n578 VSUBS 0.008018f
C1570 B.n579 VSUBS 0.008018f
C1571 B.n580 VSUBS 0.008018f
C1572 B.n581 VSUBS 0.008018f
C1573 B.n582 VSUBS 0.008018f
C1574 B.n583 VSUBS 0.008018f
C1575 B.n584 VSUBS 0.008018f
C1576 B.n585 VSUBS 0.008018f
C1577 B.n586 VSUBS 0.008018f
C1578 B.n587 VSUBS 0.008018f
C1579 B.n588 VSUBS 0.008018f
C1580 B.n589 VSUBS 0.008018f
C1581 B.n590 VSUBS 0.008018f
C1582 B.n591 VSUBS 0.008018f
C1583 B.n592 VSUBS 0.008018f
C1584 B.n593 VSUBS 0.008018f
C1585 B.n594 VSUBS 0.008018f
C1586 B.n595 VSUBS 0.008018f
C1587 B.n596 VSUBS 0.008018f
C1588 B.n597 VSUBS 0.008018f
C1589 B.n598 VSUBS 0.008018f
C1590 B.n599 VSUBS 0.008018f
C1591 B.n600 VSUBS 0.008018f
C1592 B.n601 VSUBS 0.008018f
C1593 B.n602 VSUBS 0.008018f
C1594 B.n603 VSUBS 0.008018f
C1595 B.n604 VSUBS 0.008018f
C1596 B.n605 VSUBS 0.008018f
C1597 B.n606 VSUBS 0.008018f
C1598 B.n607 VSUBS 0.008018f
C1599 B.n608 VSUBS 0.008018f
C1600 B.n609 VSUBS 0.008018f
C1601 B.n610 VSUBS 0.008018f
C1602 B.n611 VSUBS 0.008018f
C1603 B.n612 VSUBS 0.008018f
C1604 B.n613 VSUBS 0.008018f
C1605 B.n614 VSUBS 0.008018f
C1606 B.n615 VSUBS 0.02036f
C1607 B.n616 VSUBS 0.019495f
C1608 B.n617 VSUBS 0.02036f
C1609 B.n618 VSUBS 0.008018f
C1610 B.n619 VSUBS 0.008018f
C1611 B.n620 VSUBS 0.008018f
C1612 B.n621 VSUBS 0.008018f
C1613 B.n622 VSUBS 0.008018f
C1614 B.n623 VSUBS 0.008018f
C1615 B.n624 VSUBS 0.008018f
C1616 B.n625 VSUBS 0.008018f
C1617 B.n626 VSUBS 0.008018f
C1618 B.n627 VSUBS 0.008018f
C1619 B.n628 VSUBS 0.008018f
C1620 B.n629 VSUBS 0.008018f
C1621 B.n630 VSUBS 0.008018f
C1622 B.n631 VSUBS 0.008018f
C1623 B.n632 VSUBS 0.008018f
C1624 B.n633 VSUBS 0.008018f
C1625 B.n634 VSUBS 0.008018f
C1626 B.n635 VSUBS 0.008018f
C1627 B.n636 VSUBS 0.008018f
C1628 B.n637 VSUBS 0.008018f
C1629 B.n638 VSUBS 0.008018f
C1630 B.n639 VSUBS 0.008018f
C1631 B.n640 VSUBS 0.008018f
C1632 B.n641 VSUBS 0.008018f
C1633 B.n642 VSUBS 0.008018f
C1634 B.n643 VSUBS 0.008018f
C1635 B.n644 VSUBS 0.008018f
C1636 B.n645 VSUBS 0.008018f
C1637 B.n646 VSUBS 0.008018f
C1638 B.n647 VSUBS 0.008018f
C1639 B.n648 VSUBS 0.008018f
C1640 B.n649 VSUBS 0.008018f
C1641 B.n650 VSUBS 0.008018f
C1642 B.n651 VSUBS 0.008018f
C1643 B.n652 VSUBS 0.008018f
C1644 B.n653 VSUBS 0.008018f
C1645 B.n654 VSUBS 0.008018f
C1646 B.n655 VSUBS 0.008018f
C1647 B.n656 VSUBS 0.008018f
C1648 B.n657 VSUBS 0.008018f
C1649 B.n658 VSUBS 0.008018f
C1650 B.n659 VSUBS 0.008018f
C1651 B.n660 VSUBS 0.008018f
C1652 B.n661 VSUBS 0.008018f
C1653 B.n662 VSUBS 0.008018f
C1654 B.n663 VSUBS 0.008018f
C1655 B.n664 VSUBS 0.008018f
C1656 B.n665 VSUBS 0.008018f
C1657 B.n666 VSUBS 0.008018f
C1658 B.n667 VSUBS 0.008018f
C1659 B.n668 VSUBS 0.008018f
C1660 B.n669 VSUBS 0.008018f
C1661 B.n670 VSUBS 0.008018f
C1662 B.n671 VSUBS 0.008018f
C1663 B.n672 VSUBS 0.008018f
C1664 B.n673 VSUBS 0.008018f
C1665 B.n674 VSUBS 0.008018f
C1666 B.n675 VSUBS 0.008018f
C1667 B.n676 VSUBS 0.008018f
C1668 B.n677 VSUBS 0.008018f
C1669 B.n678 VSUBS 0.008018f
C1670 B.n679 VSUBS 0.008018f
C1671 B.n680 VSUBS 0.008018f
C1672 B.n681 VSUBS 0.008018f
C1673 B.n682 VSUBS 0.008018f
C1674 B.n683 VSUBS 0.008018f
C1675 B.n684 VSUBS 0.008018f
C1676 B.n685 VSUBS 0.008018f
C1677 B.n686 VSUBS 0.008018f
C1678 B.n687 VSUBS 0.008018f
C1679 B.n688 VSUBS 0.008018f
C1680 B.n689 VSUBS 0.008018f
C1681 B.n690 VSUBS 0.008018f
C1682 B.n691 VSUBS 0.008018f
C1683 B.n692 VSUBS 0.008018f
C1684 B.n693 VSUBS 0.008018f
C1685 B.n694 VSUBS 0.008018f
C1686 B.n695 VSUBS 0.008018f
C1687 B.n696 VSUBS 0.008018f
C1688 B.n697 VSUBS 0.005542f
C1689 B.n698 VSUBS 0.018577f
C1690 B.n699 VSUBS 0.006485f
C1691 B.n700 VSUBS 0.008018f
C1692 B.n701 VSUBS 0.008018f
C1693 B.n702 VSUBS 0.008018f
C1694 B.n703 VSUBS 0.008018f
C1695 B.n704 VSUBS 0.008018f
C1696 B.n705 VSUBS 0.008018f
C1697 B.n706 VSUBS 0.008018f
C1698 B.n707 VSUBS 0.008018f
C1699 B.n708 VSUBS 0.008018f
C1700 B.n709 VSUBS 0.008018f
C1701 B.n710 VSUBS 0.008018f
C1702 B.n711 VSUBS 0.006485f
C1703 B.n712 VSUBS 0.018577f
C1704 B.n713 VSUBS 0.005542f
C1705 B.n714 VSUBS 0.008018f
C1706 B.n715 VSUBS 0.008018f
C1707 B.n716 VSUBS 0.008018f
C1708 B.n717 VSUBS 0.008018f
C1709 B.n718 VSUBS 0.008018f
C1710 B.n719 VSUBS 0.008018f
C1711 B.n720 VSUBS 0.008018f
C1712 B.n721 VSUBS 0.008018f
C1713 B.n722 VSUBS 0.008018f
C1714 B.n723 VSUBS 0.008018f
C1715 B.n724 VSUBS 0.008018f
C1716 B.n725 VSUBS 0.008018f
C1717 B.n726 VSUBS 0.008018f
C1718 B.n727 VSUBS 0.008018f
C1719 B.n728 VSUBS 0.008018f
C1720 B.n729 VSUBS 0.008018f
C1721 B.n730 VSUBS 0.008018f
C1722 B.n731 VSUBS 0.008018f
C1723 B.n732 VSUBS 0.008018f
C1724 B.n733 VSUBS 0.008018f
C1725 B.n734 VSUBS 0.008018f
C1726 B.n735 VSUBS 0.008018f
C1727 B.n736 VSUBS 0.008018f
C1728 B.n737 VSUBS 0.008018f
C1729 B.n738 VSUBS 0.008018f
C1730 B.n739 VSUBS 0.008018f
C1731 B.n740 VSUBS 0.008018f
C1732 B.n741 VSUBS 0.008018f
C1733 B.n742 VSUBS 0.008018f
C1734 B.n743 VSUBS 0.008018f
C1735 B.n744 VSUBS 0.008018f
C1736 B.n745 VSUBS 0.008018f
C1737 B.n746 VSUBS 0.008018f
C1738 B.n747 VSUBS 0.008018f
C1739 B.n748 VSUBS 0.008018f
C1740 B.n749 VSUBS 0.008018f
C1741 B.n750 VSUBS 0.008018f
C1742 B.n751 VSUBS 0.008018f
C1743 B.n752 VSUBS 0.008018f
C1744 B.n753 VSUBS 0.008018f
C1745 B.n754 VSUBS 0.008018f
C1746 B.n755 VSUBS 0.008018f
C1747 B.n756 VSUBS 0.008018f
C1748 B.n757 VSUBS 0.008018f
C1749 B.n758 VSUBS 0.008018f
C1750 B.n759 VSUBS 0.008018f
C1751 B.n760 VSUBS 0.008018f
C1752 B.n761 VSUBS 0.008018f
C1753 B.n762 VSUBS 0.008018f
C1754 B.n763 VSUBS 0.008018f
C1755 B.n764 VSUBS 0.008018f
C1756 B.n765 VSUBS 0.008018f
C1757 B.n766 VSUBS 0.008018f
C1758 B.n767 VSUBS 0.008018f
C1759 B.n768 VSUBS 0.008018f
C1760 B.n769 VSUBS 0.008018f
C1761 B.n770 VSUBS 0.008018f
C1762 B.n771 VSUBS 0.008018f
C1763 B.n772 VSUBS 0.008018f
C1764 B.n773 VSUBS 0.008018f
C1765 B.n774 VSUBS 0.008018f
C1766 B.n775 VSUBS 0.008018f
C1767 B.n776 VSUBS 0.008018f
C1768 B.n777 VSUBS 0.008018f
C1769 B.n778 VSUBS 0.008018f
C1770 B.n779 VSUBS 0.008018f
C1771 B.n780 VSUBS 0.008018f
C1772 B.n781 VSUBS 0.008018f
C1773 B.n782 VSUBS 0.008018f
C1774 B.n783 VSUBS 0.008018f
C1775 B.n784 VSUBS 0.008018f
C1776 B.n785 VSUBS 0.008018f
C1777 B.n786 VSUBS 0.008018f
C1778 B.n787 VSUBS 0.008018f
C1779 B.n788 VSUBS 0.008018f
C1780 B.n789 VSUBS 0.008018f
C1781 B.n790 VSUBS 0.008018f
C1782 B.n791 VSUBS 0.008018f
C1783 B.n792 VSUBS 0.008018f
C1784 B.n793 VSUBS 0.02036f
C1785 B.n794 VSUBS 0.019495f
C1786 B.n795 VSUBS 0.019495f
C1787 B.n796 VSUBS 0.008018f
C1788 B.n797 VSUBS 0.008018f
C1789 B.n798 VSUBS 0.008018f
C1790 B.n799 VSUBS 0.008018f
C1791 B.n800 VSUBS 0.008018f
C1792 B.n801 VSUBS 0.008018f
C1793 B.n802 VSUBS 0.008018f
C1794 B.n803 VSUBS 0.008018f
C1795 B.n804 VSUBS 0.008018f
C1796 B.n805 VSUBS 0.008018f
C1797 B.n806 VSUBS 0.008018f
C1798 B.n807 VSUBS 0.008018f
C1799 B.n808 VSUBS 0.008018f
C1800 B.n809 VSUBS 0.008018f
C1801 B.n810 VSUBS 0.008018f
C1802 B.n811 VSUBS 0.008018f
C1803 B.n812 VSUBS 0.008018f
C1804 B.n813 VSUBS 0.008018f
C1805 B.n814 VSUBS 0.008018f
C1806 B.n815 VSUBS 0.008018f
C1807 B.n816 VSUBS 0.008018f
C1808 B.n817 VSUBS 0.008018f
C1809 B.n818 VSUBS 0.008018f
C1810 B.n819 VSUBS 0.008018f
C1811 B.n820 VSUBS 0.008018f
C1812 B.n821 VSUBS 0.008018f
C1813 B.n822 VSUBS 0.008018f
C1814 B.n823 VSUBS 0.008018f
C1815 B.n824 VSUBS 0.008018f
C1816 B.n825 VSUBS 0.008018f
C1817 B.n826 VSUBS 0.008018f
C1818 B.n827 VSUBS 0.008018f
C1819 B.n828 VSUBS 0.008018f
C1820 B.n829 VSUBS 0.008018f
C1821 B.n830 VSUBS 0.008018f
C1822 B.n831 VSUBS 0.008018f
C1823 B.n832 VSUBS 0.008018f
C1824 B.n833 VSUBS 0.008018f
C1825 B.n834 VSUBS 0.008018f
C1826 B.n835 VSUBS 0.008018f
C1827 B.n836 VSUBS 0.008018f
C1828 B.n837 VSUBS 0.008018f
C1829 B.n838 VSUBS 0.008018f
C1830 B.n839 VSUBS 0.008018f
C1831 B.n840 VSUBS 0.008018f
C1832 B.n841 VSUBS 0.008018f
C1833 B.n842 VSUBS 0.008018f
C1834 B.n843 VSUBS 0.008018f
C1835 B.n844 VSUBS 0.008018f
C1836 B.n845 VSUBS 0.008018f
C1837 B.n846 VSUBS 0.008018f
C1838 B.n847 VSUBS 0.008018f
C1839 B.n848 VSUBS 0.008018f
C1840 B.n849 VSUBS 0.008018f
C1841 B.n850 VSUBS 0.008018f
C1842 B.n851 VSUBS 0.008018f
C1843 B.n852 VSUBS 0.008018f
C1844 B.n853 VSUBS 0.008018f
C1845 B.n854 VSUBS 0.008018f
C1846 B.n855 VSUBS 0.008018f
C1847 B.n856 VSUBS 0.008018f
C1848 B.n857 VSUBS 0.008018f
C1849 B.n858 VSUBS 0.008018f
C1850 B.n859 VSUBS 0.008018f
C1851 B.n860 VSUBS 0.008018f
C1852 B.n861 VSUBS 0.008018f
C1853 B.n862 VSUBS 0.008018f
C1854 B.n863 VSUBS 0.008018f
C1855 B.n864 VSUBS 0.008018f
C1856 B.n865 VSUBS 0.008018f
C1857 B.n866 VSUBS 0.008018f
C1858 B.n867 VSUBS 0.018156f
.ends

