* NGSPICE file created from diff_pair_sample_1609.ext - technology: sky130A

.subckt diff_pair_sample_1609 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t1 w_n5130_n2414# sky130_fd_pr__pfet_01v8 ad=2.8197 pd=15.24 as=1.19295 ps=7.56 w=7.23 l=3.83
X1 VTAIL.t14 VP.t1 VDD1.t2 w_n5130_n2414# sky130_fd_pr__pfet_01v8 ad=1.19295 pd=7.56 as=1.19295 ps=7.56 w=7.23 l=3.83
X2 VTAIL.t3 VN.t0 VDD2.t7 w_n5130_n2414# sky130_fd_pr__pfet_01v8 ad=2.8197 pd=15.24 as=1.19295 ps=7.56 w=7.23 l=3.83
X3 VDD1.t6 VP.t2 VTAIL.t13 w_n5130_n2414# sky130_fd_pr__pfet_01v8 ad=1.19295 pd=7.56 as=1.19295 ps=7.56 w=7.23 l=3.83
X4 VDD2.t6 VN.t1 VTAIL.t0 w_n5130_n2414# sky130_fd_pr__pfet_01v8 ad=1.19295 pd=7.56 as=1.19295 ps=7.56 w=7.23 l=3.83
X5 B.t11 B.t9 B.t10 w_n5130_n2414# sky130_fd_pr__pfet_01v8 ad=2.8197 pd=15.24 as=0 ps=0 w=7.23 l=3.83
X6 VDD2.t5 VN.t2 VTAIL.t1 w_n5130_n2414# sky130_fd_pr__pfet_01v8 ad=1.19295 pd=7.56 as=1.19295 ps=7.56 w=7.23 l=3.83
X7 VDD1.t5 VP.t3 VTAIL.t12 w_n5130_n2414# sky130_fd_pr__pfet_01v8 ad=1.19295 pd=7.56 as=2.8197 ps=15.24 w=7.23 l=3.83
X8 VTAIL.t4 VN.t3 VDD2.t4 w_n5130_n2414# sky130_fd_pr__pfet_01v8 ad=2.8197 pd=15.24 as=1.19295 ps=7.56 w=7.23 l=3.83
X9 VDD2.t3 VN.t4 VTAIL.t5 w_n5130_n2414# sky130_fd_pr__pfet_01v8 ad=1.19295 pd=7.56 as=2.8197 ps=15.24 w=7.23 l=3.83
X10 VTAIL.t11 VP.t4 VDD1.t7 w_n5130_n2414# sky130_fd_pr__pfet_01v8 ad=2.8197 pd=15.24 as=1.19295 ps=7.56 w=7.23 l=3.83
X11 VTAIL.t10 VP.t5 VDD1.t0 w_n5130_n2414# sky130_fd_pr__pfet_01v8 ad=1.19295 pd=7.56 as=1.19295 ps=7.56 w=7.23 l=3.83
X12 VDD1.t3 VP.t6 VTAIL.t9 w_n5130_n2414# sky130_fd_pr__pfet_01v8 ad=1.19295 pd=7.56 as=2.8197 ps=15.24 w=7.23 l=3.83
X13 B.t8 B.t6 B.t7 w_n5130_n2414# sky130_fd_pr__pfet_01v8 ad=2.8197 pd=15.24 as=0 ps=0 w=7.23 l=3.83
X14 VDD1.t4 VP.t7 VTAIL.t8 w_n5130_n2414# sky130_fd_pr__pfet_01v8 ad=1.19295 pd=7.56 as=1.19295 ps=7.56 w=7.23 l=3.83
X15 VTAIL.t6 VN.t5 VDD2.t2 w_n5130_n2414# sky130_fd_pr__pfet_01v8 ad=1.19295 pd=7.56 as=1.19295 ps=7.56 w=7.23 l=3.83
X16 B.t5 B.t3 B.t4 w_n5130_n2414# sky130_fd_pr__pfet_01v8 ad=2.8197 pd=15.24 as=0 ps=0 w=7.23 l=3.83
X17 B.t2 B.t0 B.t1 w_n5130_n2414# sky130_fd_pr__pfet_01v8 ad=2.8197 pd=15.24 as=0 ps=0 w=7.23 l=3.83
X18 VTAIL.t7 VN.t6 VDD2.t1 w_n5130_n2414# sky130_fd_pr__pfet_01v8 ad=1.19295 pd=7.56 as=1.19295 ps=7.56 w=7.23 l=3.83
X19 VDD2.t0 VN.t7 VTAIL.t2 w_n5130_n2414# sky130_fd_pr__pfet_01v8 ad=1.19295 pd=7.56 as=2.8197 ps=15.24 w=7.23 l=3.83
R0 VP.n23 VP.n22 161.3
R1 VP.n24 VP.n19 161.3
R2 VP.n26 VP.n25 161.3
R3 VP.n27 VP.n18 161.3
R4 VP.n29 VP.n28 161.3
R5 VP.n30 VP.n17 161.3
R6 VP.n32 VP.n31 161.3
R7 VP.n33 VP.n16 161.3
R8 VP.n36 VP.n35 161.3
R9 VP.n37 VP.n15 161.3
R10 VP.n39 VP.n38 161.3
R11 VP.n40 VP.n14 161.3
R12 VP.n42 VP.n41 161.3
R13 VP.n43 VP.n13 161.3
R14 VP.n45 VP.n44 161.3
R15 VP.n46 VP.n12 161.3
R16 VP.n88 VP.n0 161.3
R17 VP.n87 VP.n86 161.3
R18 VP.n85 VP.n1 161.3
R19 VP.n84 VP.n83 161.3
R20 VP.n82 VP.n2 161.3
R21 VP.n81 VP.n80 161.3
R22 VP.n79 VP.n3 161.3
R23 VP.n78 VP.n77 161.3
R24 VP.n75 VP.n4 161.3
R25 VP.n74 VP.n73 161.3
R26 VP.n72 VP.n5 161.3
R27 VP.n71 VP.n70 161.3
R28 VP.n69 VP.n6 161.3
R29 VP.n68 VP.n67 161.3
R30 VP.n66 VP.n7 161.3
R31 VP.n65 VP.n64 161.3
R32 VP.n62 VP.n8 161.3
R33 VP.n61 VP.n60 161.3
R34 VP.n59 VP.n9 161.3
R35 VP.n58 VP.n57 161.3
R36 VP.n56 VP.n10 161.3
R37 VP.n55 VP.n54 161.3
R38 VP.n53 VP.n11 161.3
R39 VP.n52 VP.n51 161.3
R40 VP.n20 VP.t0 77.5753
R41 VP.n21 VP.n20 58.9368
R42 VP.n50 VP.n49 58.2041
R43 VP.n90 VP.n89 58.2041
R44 VP.n48 VP.n47 58.2041
R45 VP.n70 VP.n69 56.5193
R46 VP.n28 VP.n27 56.5193
R47 VP.n49 VP.n48 53.2994
R48 VP.n57 VP.n56 49.2348
R49 VP.n83 VP.n82 49.2348
R50 VP.n41 VP.n40 49.2348
R51 VP.n50 VP.t4 45.4948
R52 VP.n63 VP.t7 45.4948
R53 VP.n76 VP.t5 45.4948
R54 VP.n89 VP.t6 45.4948
R55 VP.n47 VP.t3 45.4948
R56 VP.n34 VP.t1 45.4948
R57 VP.n21 VP.t2 45.4948
R58 VP.n56 VP.n55 31.752
R59 VP.n83 VP.n1 31.752
R60 VP.n41 VP.n13 31.752
R61 VP.n51 VP.n11 24.4675
R62 VP.n55 VP.n11 24.4675
R63 VP.n57 VP.n9 24.4675
R64 VP.n61 VP.n9 24.4675
R65 VP.n62 VP.n61 24.4675
R66 VP.n64 VP.n7 24.4675
R67 VP.n68 VP.n7 24.4675
R68 VP.n69 VP.n68 24.4675
R69 VP.n70 VP.n5 24.4675
R70 VP.n74 VP.n5 24.4675
R71 VP.n75 VP.n74 24.4675
R72 VP.n77 VP.n3 24.4675
R73 VP.n81 VP.n3 24.4675
R74 VP.n82 VP.n81 24.4675
R75 VP.n87 VP.n1 24.4675
R76 VP.n88 VP.n87 24.4675
R77 VP.n45 VP.n13 24.4675
R78 VP.n46 VP.n45 24.4675
R79 VP.n28 VP.n17 24.4675
R80 VP.n32 VP.n17 24.4675
R81 VP.n33 VP.n32 24.4675
R82 VP.n35 VP.n15 24.4675
R83 VP.n39 VP.n15 24.4675
R84 VP.n40 VP.n39 24.4675
R85 VP.n22 VP.n19 24.4675
R86 VP.n26 VP.n19 24.4675
R87 VP.n27 VP.n26 24.4675
R88 VP.n51 VP.n50 23.9782
R89 VP.n89 VP.n88 23.9782
R90 VP.n47 VP.n46 23.9782
R91 VP.n64 VP.n63 16.1487
R92 VP.n76 VP.n75 16.1487
R93 VP.n34 VP.n33 16.1487
R94 VP.n22 VP.n21 16.1487
R95 VP.n63 VP.n62 8.31928
R96 VP.n77 VP.n76 8.31928
R97 VP.n35 VP.n34 8.31928
R98 VP.n23 VP.n20 2.5472
R99 VP.n48 VP.n12 0.417535
R100 VP.n52 VP.n49 0.417535
R101 VP.n90 VP.n0 0.417535
R102 VP VP.n90 0.394291
R103 VP.n24 VP.n23 0.189894
R104 VP.n25 VP.n24 0.189894
R105 VP.n25 VP.n18 0.189894
R106 VP.n29 VP.n18 0.189894
R107 VP.n30 VP.n29 0.189894
R108 VP.n31 VP.n30 0.189894
R109 VP.n31 VP.n16 0.189894
R110 VP.n36 VP.n16 0.189894
R111 VP.n37 VP.n36 0.189894
R112 VP.n38 VP.n37 0.189894
R113 VP.n38 VP.n14 0.189894
R114 VP.n42 VP.n14 0.189894
R115 VP.n43 VP.n42 0.189894
R116 VP.n44 VP.n43 0.189894
R117 VP.n44 VP.n12 0.189894
R118 VP.n53 VP.n52 0.189894
R119 VP.n54 VP.n53 0.189894
R120 VP.n54 VP.n10 0.189894
R121 VP.n58 VP.n10 0.189894
R122 VP.n59 VP.n58 0.189894
R123 VP.n60 VP.n59 0.189894
R124 VP.n60 VP.n8 0.189894
R125 VP.n65 VP.n8 0.189894
R126 VP.n66 VP.n65 0.189894
R127 VP.n67 VP.n66 0.189894
R128 VP.n67 VP.n6 0.189894
R129 VP.n71 VP.n6 0.189894
R130 VP.n72 VP.n71 0.189894
R131 VP.n73 VP.n72 0.189894
R132 VP.n73 VP.n4 0.189894
R133 VP.n78 VP.n4 0.189894
R134 VP.n79 VP.n78 0.189894
R135 VP.n80 VP.n79 0.189894
R136 VP.n80 VP.n2 0.189894
R137 VP.n84 VP.n2 0.189894
R138 VP.n85 VP.n84 0.189894
R139 VP.n86 VP.n85 0.189894
R140 VP.n86 VP.n0 0.189894
R141 VDD1 VDD1.n0 89.5992
R142 VDD1.n3 VDD1.n2 89.4856
R143 VDD1.n3 VDD1.n1 89.4856
R144 VDD1.n5 VDD1.n4 87.7478
R145 VDD1.n5 VDD1.n3 46.669
R146 VDD1.n4 VDD1.t2 4.49635
R147 VDD1.n4 VDD1.t5 4.49635
R148 VDD1.n0 VDD1.t1 4.49635
R149 VDD1.n0 VDD1.t6 4.49635
R150 VDD1.n2 VDD1.t0 4.49635
R151 VDD1.n2 VDD1.t3 4.49635
R152 VDD1.n1 VDD1.t7 4.49635
R153 VDD1.n1 VDD1.t4 4.49635
R154 VDD1 VDD1.n5 1.73541
R155 VTAIL.n273 VTAIL.n272 585
R156 VTAIL.n275 VTAIL.n274 585
R157 VTAIL.n268 VTAIL.n267 585
R158 VTAIL.n281 VTAIL.n280 585
R159 VTAIL.n283 VTAIL.n282 585
R160 VTAIL.n264 VTAIL.n263 585
R161 VTAIL.n289 VTAIL.n288 585
R162 VTAIL.n291 VTAIL.n290 585
R163 VTAIL.n15 VTAIL.n14 585
R164 VTAIL.n17 VTAIL.n16 585
R165 VTAIL.n10 VTAIL.n9 585
R166 VTAIL.n23 VTAIL.n22 585
R167 VTAIL.n25 VTAIL.n24 585
R168 VTAIL.n6 VTAIL.n5 585
R169 VTAIL.n31 VTAIL.n30 585
R170 VTAIL.n33 VTAIL.n32 585
R171 VTAIL.n51 VTAIL.n50 585
R172 VTAIL.n53 VTAIL.n52 585
R173 VTAIL.n46 VTAIL.n45 585
R174 VTAIL.n59 VTAIL.n58 585
R175 VTAIL.n61 VTAIL.n60 585
R176 VTAIL.n42 VTAIL.n41 585
R177 VTAIL.n67 VTAIL.n66 585
R178 VTAIL.n69 VTAIL.n68 585
R179 VTAIL.n89 VTAIL.n88 585
R180 VTAIL.n91 VTAIL.n90 585
R181 VTAIL.n84 VTAIL.n83 585
R182 VTAIL.n97 VTAIL.n96 585
R183 VTAIL.n99 VTAIL.n98 585
R184 VTAIL.n80 VTAIL.n79 585
R185 VTAIL.n105 VTAIL.n104 585
R186 VTAIL.n107 VTAIL.n106 585
R187 VTAIL.n255 VTAIL.n254 585
R188 VTAIL.n253 VTAIL.n252 585
R189 VTAIL.n228 VTAIL.n227 585
R190 VTAIL.n247 VTAIL.n246 585
R191 VTAIL.n245 VTAIL.n244 585
R192 VTAIL.n232 VTAIL.n231 585
R193 VTAIL.n239 VTAIL.n238 585
R194 VTAIL.n237 VTAIL.n236 585
R195 VTAIL.n217 VTAIL.n216 585
R196 VTAIL.n215 VTAIL.n214 585
R197 VTAIL.n190 VTAIL.n189 585
R198 VTAIL.n209 VTAIL.n208 585
R199 VTAIL.n207 VTAIL.n206 585
R200 VTAIL.n194 VTAIL.n193 585
R201 VTAIL.n201 VTAIL.n200 585
R202 VTAIL.n199 VTAIL.n198 585
R203 VTAIL.n181 VTAIL.n180 585
R204 VTAIL.n179 VTAIL.n178 585
R205 VTAIL.n154 VTAIL.n153 585
R206 VTAIL.n173 VTAIL.n172 585
R207 VTAIL.n171 VTAIL.n170 585
R208 VTAIL.n158 VTAIL.n157 585
R209 VTAIL.n165 VTAIL.n164 585
R210 VTAIL.n163 VTAIL.n162 585
R211 VTAIL.n143 VTAIL.n142 585
R212 VTAIL.n141 VTAIL.n140 585
R213 VTAIL.n116 VTAIL.n115 585
R214 VTAIL.n135 VTAIL.n134 585
R215 VTAIL.n133 VTAIL.n132 585
R216 VTAIL.n120 VTAIL.n119 585
R217 VTAIL.n127 VTAIL.n126 585
R218 VTAIL.n125 VTAIL.n124 585
R219 VTAIL.n290 VTAIL.n260 498.474
R220 VTAIL.n32 VTAIL.n2 498.474
R221 VTAIL.n68 VTAIL.n38 498.474
R222 VTAIL.n106 VTAIL.n76 498.474
R223 VTAIL.n254 VTAIL.n224 498.474
R224 VTAIL.n216 VTAIL.n186 498.474
R225 VTAIL.n180 VTAIL.n150 498.474
R226 VTAIL.n142 VTAIL.n112 498.474
R227 VTAIL.n271 VTAIL.t2 329.053
R228 VTAIL.n13 VTAIL.t4 329.053
R229 VTAIL.n49 VTAIL.t9 329.053
R230 VTAIL.n87 VTAIL.t11 329.053
R231 VTAIL.n235 VTAIL.t12 329.053
R232 VTAIL.n197 VTAIL.t15 329.053
R233 VTAIL.n161 VTAIL.t5 329.053
R234 VTAIL.n123 VTAIL.t3 329.053
R235 VTAIL.n274 VTAIL.n273 171.744
R236 VTAIL.n274 VTAIL.n267 171.744
R237 VTAIL.n281 VTAIL.n267 171.744
R238 VTAIL.n282 VTAIL.n281 171.744
R239 VTAIL.n282 VTAIL.n263 171.744
R240 VTAIL.n289 VTAIL.n263 171.744
R241 VTAIL.n290 VTAIL.n289 171.744
R242 VTAIL.n16 VTAIL.n15 171.744
R243 VTAIL.n16 VTAIL.n9 171.744
R244 VTAIL.n23 VTAIL.n9 171.744
R245 VTAIL.n24 VTAIL.n23 171.744
R246 VTAIL.n24 VTAIL.n5 171.744
R247 VTAIL.n31 VTAIL.n5 171.744
R248 VTAIL.n32 VTAIL.n31 171.744
R249 VTAIL.n52 VTAIL.n51 171.744
R250 VTAIL.n52 VTAIL.n45 171.744
R251 VTAIL.n59 VTAIL.n45 171.744
R252 VTAIL.n60 VTAIL.n59 171.744
R253 VTAIL.n60 VTAIL.n41 171.744
R254 VTAIL.n67 VTAIL.n41 171.744
R255 VTAIL.n68 VTAIL.n67 171.744
R256 VTAIL.n90 VTAIL.n89 171.744
R257 VTAIL.n90 VTAIL.n83 171.744
R258 VTAIL.n97 VTAIL.n83 171.744
R259 VTAIL.n98 VTAIL.n97 171.744
R260 VTAIL.n98 VTAIL.n79 171.744
R261 VTAIL.n105 VTAIL.n79 171.744
R262 VTAIL.n106 VTAIL.n105 171.744
R263 VTAIL.n254 VTAIL.n253 171.744
R264 VTAIL.n253 VTAIL.n227 171.744
R265 VTAIL.n246 VTAIL.n227 171.744
R266 VTAIL.n246 VTAIL.n245 171.744
R267 VTAIL.n245 VTAIL.n231 171.744
R268 VTAIL.n238 VTAIL.n231 171.744
R269 VTAIL.n238 VTAIL.n237 171.744
R270 VTAIL.n216 VTAIL.n215 171.744
R271 VTAIL.n215 VTAIL.n189 171.744
R272 VTAIL.n208 VTAIL.n189 171.744
R273 VTAIL.n208 VTAIL.n207 171.744
R274 VTAIL.n207 VTAIL.n193 171.744
R275 VTAIL.n200 VTAIL.n193 171.744
R276 VTAIL.n200 VTAIL.n199 171.744
R277 VTAIL.n180 VTAIL.n179 171.744
R278 VTAIL.n179 VTAIL.n153 171.744
R279 VTAIL.n172 VTAIL.n153 171.744
R280 VTAIL.n172 VTAIL.n171 171.744
R281 VTAIL.n171 VTAIL.n157 171.744
R282 VTAIL.n164 VTAIL.n157 171.744
R283 VTAIL.n164 VTAIL.n163 171.744
R284 VTAIL.n142 VTAIL.n141 171.744
R285 VTAIL.n141 VTAIL.n115 171.744
R286 VTAIL.n134 VTAIL.n115 171.744
R287 VTAIL.n134 VTAIL.n133 171.744
R288 VTAIL.n133 VTAIL.n119 171.744
R289 VTAIL.n126 VTAIL.n119 171.744
R290 VTAIL.n126 VTAIL.n125 171.744
R291 VTAIL.n273 VTAIL.t2 85.8723
R292 VTAIL.n15 VTAIL.t4 85.8723
R293 VTAIL.n51 VTAIL.t9 85.8723
R294 VTAIL.n89 VTAIL.t11 85.8723
R295 VTAIL.n237 VTAIL.t12 85.8723
R296 VTAIL.n199 VTAIL.t15 85.8723
R297 VTAIL.n163 VTAIL.t5 85.8723
R298 VTAIL.n125 VTAIL.t3 85.8723
R299 VTAIL.n223 VTAIL.n222 71.0691
R300 VTAIL.n149 VTAIL.n148 71.0691
R301 VTAIL.n1 VTAIL.n0 71.069
R302 VTAIL.n75 VTAIL.n74 71.069
R303 VTAIL.n295 VTAIL.n294 35.0944
R304 VTAIL.n37 VTAIL.n36 35.0944
R305 VTAIL.n73 VTAIL.n72 35.0944
R306 VTAIL.n111 VTAIL.n110 35.0944
R307 VTAIL.n259 VTAIL.n258 35.0944
R308 VTAIL.n221 VTAIL.n220 35.0944
R309 VTAIL.n185 VTAIL.n184 35.0944
R310 VTAIL.n147 VTAIL.n146 35.0944
R311 VTAIL.n295 VTAIL.n259 22.1858
R312 VTAIL.n147 VTAIL.n111 22.1858
R313 VTAIL.n292 VTAIL.n291 12.8005
R314 VTAIL.n34 VTAIL.n33 12.8005
R315 VTAIL.n70 VTAIL.n69 12.8005
R316 VTAIL.n108 VTAIL.n107 12.8005
R317 VTAIL.n256 VTAIL.n255 12.8005
R318 VTAIL.n218 VTAIL.n217 12.8005
R319 VTAIL.n182 VTAIL.n181 12.8005
R320 VTAIL.n144 VTAIL.n143 12.8005
R321 VTAIL.n288 VTAIL.n262 12.0247
R322 VTAIL.n30 VTAIL.n4 12.0247
R323 VTAIL.n66 VTAIL.n40 12.0247
R324 VTAIL.n104 VTAIL.n78 12.0247
R325 VTAIL.n252 VTAIL.n226 12.0247
R326 VTAIL.n214 VTAIL.n188 12.0247
R327 VTAIL.n178 VTAIL.n152 12.0247
R328 VTAIL.n140 VTAIL.n114 12.0247
R329 VTAIL.n287 VTAIL.n264 11.249
R330 VTAIL.n29 VTAIL.n6 11.249
R331 VTAIL.n65 VTAIL.n42 11.249
R332 VTAIL.n103 VTAIL.n80 11.249
R333 VTAIL.n251 VTAIL.n228 11.249
R334 VTAIL.n213 VTAIL.n190 11.249
R335 VTAIL.n177 VTAIL.n154 11.249
R336 VTAIL.n139 VTAIL.n116 11.249
R337 VTAIL.n272 VTAIL.n271 10.7237
R338 VTAIL.n14 VTAIL.n13 10.7237
R339 VTAIL.n50 VTAIL.n49 10.7237
R340 VTAIL.n88 VTAIL.n87 10.7237
R341 VTAIL.n236 VTAIL.n235 10.7237
R342 VTAIL.n198 VTAIL.n197 10.7237
R343 VTAIL.n162 VTAIL.n161 10.7237
R344 VTAIL.n124 VTAIL.n123 10.7237
R345 VTAIL.n284 VTAIL.n283 10.4732
R346 VTAIL.n26 VTAIL.n25 10.4732
R347 VTAIL.n62 VTAIL.n61 10.4732
R348 VTAIL.n100 VTAIL.n99 10.4732
R349 VTAIL.n248 VTAIL.n247 10.4732
R350 VTAIL.n210 VTAIL.n209 10.4732
R351 VTAIL.n174 VTAIL.n173 10.4732
R352 VTAIL.n136 VTAIL.n135 10.4732
R353 VTAIL.n280 VTAIL.n266 9.69747
R354 VTAIL.n22 VTAIL.n8 9.69747
R355 VTAIL.n58 VTAIL.n44 9.69747
R356 VTAIL.n96 VTAIL.n82 9.69747
R357 VTAIL.n244 VTAIL.n230 9.69747
R358 VTAIL.n206 VTAIL.n192 9.69747
R359 VTAIL.n170 VTAIL.n156 9.69747
R360 VTAIL.n132 VTAIL.n118 9.69747
R361 VTAIL.n294 VTAIL.n293 9.45567
R362 VTAIL.n36 VTAIL.n35 9.45567
R363 VTAIL.n72 VTAIL.n71 9.45567
R364 VTAIL.n110 VTAIL.n109 9.45567
R365 VTAIL.n258 VTAIL.n257 9.45567
R366 VTAIL.n220 VTAIL.n219 9.45567
R367 VTAIL.n184 VTAIL.n183 9.45567
R368 VTAIL.n146 VTAIL.n145 9.45567
R369 VTAIL.n270 VTAIL.n269 9.3005
R370 VTAIL.n277 VTAIL.n276 9.3005
R371 VTAIL.n279 VTAIL.n278 9.3005
R372 VTAIL.n266 VTAIL.n265 9.3005
R373 VTAIL.n285 VTAIL.n284 9.3005
R374 VTAIL.n287 VTAIL.n286 9.3005
R375 VTAIL.n262 VTAIL.n261 9.3005
R376 VTAIL.n293 VTAIL.n292 9.3005
R377 VTAIL.n12 VTAIL.n11 9.3005
R378 VTAIL.n19 VTAIL.n18 9.3005
R379 VTAIL.n21 VTAIL.n20 9.3005
R380 VTAIL.n8 VTAIL.n7 9.3005
R381 VTAIL.n27 VTAIL.n26 9.3005
R382 VTAIL.n29 VTAIL.n28 9.3005
R383 VTAIL.n4 VTAIL.n3 9.3005
R384 VTAIL.n35 VTAIL.n34 9.3005
R385 VTAIL.n48 VTAIL.n47 9.3005
R386 VTAIL.n55 VTAIL.n54 9.3005
R387 VTAIL.n57 VTAIL.n56 9.3005
R388 VTAIL.n44 VTAIL.n43 9.3005
R389 VTAIL.n63 VTAIL.n62 9.3005
R390 VTAIL.n65 VTAIL.n64 9.3005
R391 VTAIL.n40 VTAIL.n39 9.3005
R392 VTAIL.n71 VTAIL.n70 9.3005
R393 VTAIL.n86 VTAIL.n85 9.3005
R394 VTAIL.n93 VTAIL.n92 9.3005
R395 VTAIL.n95 VTAIL.n94 9.3005
R396 VTAIL.n82 VTAIL.n81 9.3005
R397 VTAIL.n101 VTAIL.n100 9.3005
R398 VTAIL.n103 VTAIL.n102 9.3005
R399 VTAIL.n78 VTAIL.n77 9.3005
R400 VTAIL.n109 VTAIL.n108 9.3005
R401 VTAIL.n234 VTAIL.n233 9.3005
R402 VTAIL.n241 VTAIL.n240 9.3005
R403 VTAIL.n243 VTAIL.n242 9.3005
R404 VTAIL.n230 VTAIL.n229 9.3005
R405 VTAIL.n249 VTAIL.n248 9.3005
R406 VTAIL.n251 VTAIL.n250 9.3005
R407 VTAIL.n226 VTAIL.n225 9.3005
R408 VTAIL.n257 VTAIL.n256 9.3005
R409 VTAIL.n196 VTAIL.n195 9.3005
R410 VTAIL.n203 VTAIL.n202 9.3005
R411 VTAIL.n205 VTAIL.n204 9.3005
R412 VTAIL.n192 VTAIL.n191 9.3005
R413 VTAIL.n211 VTAIL.n210 9.3005
R414 VTAIL.n213 VTAIL.n212 9.3005
R415 VTAIL.n188 VTAIL.n187 9.3005
R416 VTAIL.n219 VTAIL.n218 9.3005
R417 VTAIL.n160 VTAIL.n159 9.3005
R418 VTAIL.n167 VTAIL.n166 9.3005
R419 VTAIL.n169 VTAIL.n168 9.3005
R420 VTAIL.n156 VTAIL.n155 9.3005
R421 VTAIL.n175 VTAIL.n174 9.3005
R422 VTAIL.n177 VTAIL.n176 9.3005
R423 VTAIL.n152 VTAIL.n151 9.3005
R424 VTAIL.n183 VTAIL.n182 9.3005
R425 VTAIL.n122 VTAIL.n121 9.3005
R426 VTAIL.n129 VTAIL.n128 9.3005
R427 VTAIL.n131 VTAIL.n130 9.3005
R428 VTAIL.n118 VTAIL.n117 9.3005
R429 VTAIL.n137 VTAIL.n136 9.3005
R430 VTAIL.n139 VTAIL.n138 9.3005
R431 VTAIL.n114 VTAIL.n113 9.3005
R432 VTAIL.n145 VTAIL.n144 9.3005
R433 VTAIL.n279 VTAIL.n268 8.92171
R434 VTAIL.n21 VTAIL.n10 8.92171
R435 VTAIL.n57 VTAIL.n46 8.92171
R436 VTAIL.n95 VTAIL.n84 8.92171
R437 VTAIL.n243 VTAIL.n232 8.92171
R438 VTAIL.n205 VTAIL.n194 8.92171
R439 VTAIL.n169 VTAIL.n158 8.92171
R440 VTAIL.n131 VTAIL.n120 8.92171
R441 VTAIL.n276 VTAIL.n275 8.14595
R442 VTAIL.n18 VTAIL.n17 8.14595
R443 VTAIL.n54 VTAIL.n53 8.14595
R444 VTAIL.n92 VTAIL.n91 8.14595
R445 VTAIL.n240 VTAIL.n239 8.14595
R446 VTAIL.n202 VTAIL.n201 8.14595
R447 VTAIL.n166 VTAIL.n165 8.14595
R448 VTAIL.n128 VTAIL.n127 8.14595
R449 VTAIL.n294 VTAIL.n260 7.75445
R450 VTAIL.n36 VTAIL.n2 7.75445
R451 VTAIL.n72 VTAIL.n38 7.75445
R452 VTAIL.n110 VTAIL.n76 7.75445
R453 VTAIL.n258 VTAIL.n224 7.75445
R454 VTAIL.n220 VTAIL.n186 7.75445
R455 VTAIL.n184 VTAIL.n150 7.75445
R456 VTAIL.n146 VTAIL.n112 7.75445
R457 VTAIL.n272 VTAIL.n270 7.3702
R458 VTAIL.n14 VTAIL.n12 7.3702
R459 VTAIL.n50 VTAIL.n48 7.3702
R460 VTAIL.n88 VTAIL.n86 7.3702
R461 VTAIL.n236 VTAIL.n234 7.3702
R462 VTAIL.n198 VTAIL.n196 7.3702
R463 VTAIL.n162 VTAIL.n160 7.3702
R464 VTAIL.n124 VTAIL.n122 7.3702
R465 VTAIL.n292 VTAIL.n260 6.08283
R466 VTAIL.n34 VTAIL.n2 6.08283
R467 VTAIL.n70 VTAIL.n38 6.08283
R468 VTAIL.n108 VTAIL.n76 6.08283
R469 VTAIL.n256 VTAIL.n224 6.08283
R470 VTAIL.n218 VTAIL.n186 6.08283
R471 VTAIL.n182 VTAIL.n150 6.08283
R472 VTAIL.n144 VTAIL.n112 6.08283
R473 VTAIL.n275 VTAIL.n270 5.81868
R474 VTAIL.n17 VTAIL.n12 5.81868
R475 VTAIL.n53 VTAIL.n48 5.81868
R476 VTAIL.n91 VTAIL.n86 5.81868
R477 VTAIL.n239 VTAIL.n234 5.81868
R478 VTAIL.n201 VTAIL.n196 5.81868
R479 VTAIL.n165 VTAIL.n160 5.81868
R480 VTAIL.n127 VTAIL.n122 5.81868
R481 VTAIL.n276 VTAIL.n268 5.04292
R482 VTAIL.n18 VTAIL.n10 5.04292
R483 VTAIL.n54 VTAIL.n46 5.04292
R484 VTAIL.n92 VTAIL.n84 5.04292
R485 VTAIL.n240 VTAIL.n232 5.04292
R486 VTAIL.n202 VTAIL.n194 5.04292
R487 VTAIL.n166 VTAIL.n158 5.04292
R488 VTAIL.n128 VTAIL.n120 5.04292
R489 VTAIL.n0 VTAIL.t1 4.49635
R490 VTAIL.n0 VTAIL.t7 4.49635
R491 VTAIL.n74 VTAIL.t8 4.49635
R492 VTAIL.n74 VTAIL.t10 4.49635
R493 VTAIL.n222 VTAIL.t13 4.49635
R494 VTAIL.n222 VTAIL.t14 4.49635
R495 VTAIL.n148 VTAIL.t0 4.49635
R496 VTAIL.n148 VTAIL.t6 4.49635
R497 VTAIL.n280 VTAIL.n279 4.26717
R498 VTAIL.n22 VTAIL.n21 4.26717
R499 VTAIL.n58 VTAIL.n57 4.26717
R500 VTAIL.n96 VTAIL.n95 4.26717
R501 VTAIL.n244 VTAIL.n243 4.26717
R502 VTAIL.n206 VTAIL.n205 4.26717
R503 VTAIL.n170 VTAIL.n169 4.26717
R504 VTAIL.n132 VTAIL.n131 4.26717
R505 VTAIL.n149 VTAIL.n147 3.58671
R506 VTAIL.n185 VTAIL.n149 3.58671
R507 VTAIL.n223 VTAIL.n221 3.58671
R508 VTAIL.n259 VTAIL.n223 3.58671
R509 VTAIL.n111 VTAIL.n75 3.58671
R510 VTAIL.n75 VTAIL.n73 3.58671
R511 VTAIL.n37 VTAIL.n1 3.58671
R512 VTAIL VTAIL.n295 3.52852
R513 VTAIL.n283 VTAIL.n266 3.49141
R514 VTAIL.n25 VTAIL.n8 3.49141
R515 VTAIL.n61 VTAIL.n44 3.49141
R516 VTAIL.n99 VTAIL.n82 3.49141
R517 VTAIL.n247 VTAIL.n230 3.49141
R518 VTAIL.n209 VTAIL.n192 3.49141
R519 VTAIL.n173 VTAIL.n156 3.49141
R520 VTAIL.n135 VTAIL.n118 3.49141
R521 VTAIL.n284 VTAIL.n264 2.71565
R522 VTAIL.n26 VTAIL.n6 2.71565
R523 VTAIL.n62 VTAIL.n42 2.71565
R524 VTAIL.n100 VTAIL.n80 2.71565
R525 VTAIL.n248 VTAIL.n228 2.71565
R526 VTAIL.n210 VTAIL.n190 2.71565
R527 VTAIL.n174 VTAIL.n154 2.71565
R528 VTAIL.n136 VTAIL.n116 2.71565
R529 VTAIL.n271 VTAIL.n269 2.41305
R530 VTAIL.n13 VTAIL.n11 2.41305
R531 VTAIL.n49 VTAIL.n47 2.41305
R532 VTAIL.n87 VTAIL.n85 2.41305
R533 VTAIL.n235 VTAIL.n233 2.41305
R534 VTAIL.n197 VTAIL.n195 2.41305
R535 VTAIL.n161 VTAIL.n159 2.41305
R536 VTAIL.n123 VTAIL.n121 2.41305
R537 VTAIL.n288 VTAIL.n287 1.93989
R538 VTAIL.n30 VTAIL.n29 1.93989
R539 VTAIL.n66 VTAIL.n65 1.93989
R540 VTAIL.n104 VTAIL.n103 1.93989
R541 VTAIL.n252 VTAIL.n251 1.93989
R542 VTAIL.n214 VTAIL.n213 1.93989
R543 VTAIL.n178 VTAIL.n177 1.93989
R544 VTAIL.n140 VTAIL.n139 1.93989
R545 VTAIL.n291 VTAIL.n262 1.16414
R546 VTAIL.n33 VTAIL.n4 1.16414
R547 VTAIL.n69 VTAIL.n40 1.16414
R548 VTAIL.n107 VTAIL.n78 1.16414
R549 VTAIL.n255 VTAIL.n226 1.16414
R550 VTAIL.n217 VTAIL.n188 1.16414
R551 VTAIL.n181 VTAIL.n152 1.16414
R552 VTAIL.n143 VTAIL.n114 1.16414
R553 VTAIL.n221 VTAIL.n185 0.470328
R554 VTAIL.n73 VTAIL.n37 0.470328
R555 VTAIL.n277 VTAIL.n269 0.155672
R556 VTAIL.n278 VTAIL.n277 0.155672
R557 VTAIL.n278 VTAIL.n265 0.155672
R558 VTAIL.n285 VTAIL.n265 0.155672
R559 VTAIL.n286 VTAIL.n285 0.155672
R560 VTAIL.n286 VTAIL.n261 0.155672
R561 VTAIL.n293 VTAIL.n261 0.155672
R562 VTAIL.n19 VTAIL.n11 0.155672
R563 VTAIL.n20 VTAIL.n19 0.155672
R564 VTAIL.n20 VTAIL.n7 0.155672
R565 VTAIL.n27 VTAIL.n7 0.155672
R566 VTAIL.n28 VTAIL.n27 0.155672
R567 VTAIL.n28 VTAIL.n3 0.155672
R568 VTAIL.n35 VTAIL.n3 0.155672
R569 VTAIL.n55 VTAIL.n47 0.155672
R570 VTAIL.n56 VTAIL.n55 0.155672
R571 VTAIL.n56 VTAIL.n43 0.155672
R572 VTAIL.n63 VTAIL.n43 0.155672
R573 VTAIL.n64 VTAIL.n63 0.155672
R574 VTAIL.n64 VTAIL.n39 0.155672
R575 VTAIL.n71 VTAIL.n39 0.155672
R576 VTAIL.n93 VTAIL.n85 0.155672
R577 VTAIL.n94 VTAIL.n93 0.155672
R578 VTAIL.n94 VTAIL.n81 0.155672
R579 VTAIL.n101 VTAIL.n81 0.155672
R580 VTAIL.n102 VTAIL.n101 0.155672
R581 VTAIL.n102 VTAIL.n77 0.155672
R582 VTAIL.n109 VTAIL.n77 0.155672
R583 VTAIL.n257 VTAIL.n225 0.155672
R584 VTAIL.n250 VTAIL.n225 0.155672
R585 VTAIL.n250 VTAIL.n249 0.155672
R586 VTAIL.n249 VTAIL.n229 0.155672
R587 VTAIL.n242 VTAIL.n229 0.155672
R588 VTAIL.n242 VTAIL.n241 0.155672
R589 VTAIL.n241 VTAIL.n233 0.155672
R590 VTAIL.n219 VTAIL.n187 0.155672
R591 VTAIL.n212 VTAIL.n187 0.155672
R592 VTAIL.n212 VTAIL.n211 0.155672
R593 VTAIL.n211 VTAIL.n191 0.155672
R594 VTAIL.n204 VTAIL.n191 0.155672
R595 VTAIL.n204 VTAIL.n203 0.155672
R596 VTAIL.n203 VTAIL.n195 0.155672
R597 VTAIL.n183 VTAIL.n151 0.155672
R598 VTAIL.n176 VTAIL.n151 0.155672
R599 VTAIL.n176 VTAIL.n175 0.155672
R600 VTAIL.n175 VTAIL.n155 0.155672
R601 VTAIL.n168 VTAIL.n155 0.155672
R602 VTAIL.n168 VTAIL.n167 0.155672
R603 VTAIL.n167 VTAIL.n159 0.155672
R604 VTAIL.n145 VTAIL.n113 0.155672
R605 VTAIL.n138 VTAIL.n113 0.155672
R606 VTAIL.n138 VTAIL.n137 0.155672
R607 VTAIL.n137 VTAIL.n117 0.155672
R608 VTAIL.n130 VTAIL.n117 0.155672
R609 VTAIL.n130 VTAIL.n129 0.155672
R610 VTAIL.n129 VTAIL.n121 0.155672
R611 VTAIL VTAIL.n1 0.0586897
R612 VN.n71 VN.n37 161.3
R613 VN.n70 VN.n69 161.3
R614 VN.n68 VN.n38 161.3
R615 VN.n67 VN.n66 161.3
R616 VN.n65 VN.n39 161.3
R617 VN.n64 VN.n63 161.3
R618 VN.n62 VN.n40 161.3
R619 VN.n61 VN.n60 161.3
R620 VN.n58 VN.n41 161.3
R621 VN.n57 VN.n56 161.3
R622 VN.n55 VN.n42 161.3
R623 VN.n54 VN.n53 161.3
R624 VN.n52 VN.n43 161.3
R625 VN.n51 VN.n50 161.3
R626 VN.n49 VN.n44 161.3
R627 VN.n48 VN.n47 161.3
R628 VN.n34 VN.n0 161.3
R629 VN.n33 VN.n32 161.3
R630 VN.n31 VN.n1 161.3
R631 VN.n30 VN.n29 161.3
R632 VN.n28 VN.n2 161.3
R633 VN.n27 VN.n26 161.3
R634 VN.n25 VN.n3 161.3
R635 VN.n24 VN.n23 161.3
R636 VN.n21 VN.n4 161.3
R637 VN.n20 VN.n19 161.3
R638 VN.n18 VN.n5 161.3
R639 VN.n17 VN.n16 161.3
R640 VN.n15 VN.n6 161.3
R641 VN.n14 VN.n13 161.3
R642 VN.n12 VN.n7 161.3
R643 VN.n11 VN.n10 161.3
R644 VN.n8 VN.t3 77.5757
R645 VN.n45 VN.t4 77.5757
R646 VN.n9 VN.n8 58.9368
R647 VN.n46 VN.n45 58.9368
R648 VN.n36 VN.n35 58.2041
R649 VN.n73 VN.n72 58.2041
R650 VN.n16 VN.n15 56.5193
R651 VN.n53 VN.n52 56.5193
R652 VN VN.n73 53.3375
R653 VN.n29 VN.n28 49.2348
R654 VN.n66 VN.n65 49.2348
R655 VN.n9 VN.t2 45.4948
R656 VN.n22 VN.t6 45.4948
R657 VN.n35 VN.t7 45.4948
R658 VN.n46 VN.t5 45.4948
R659 VN.n59 VN.t1 45.4948
R660 VN.n72 VN.t0 45.4948
R661 VN.n29 VN.n1 31.752
R662 VN.n66 VN.n38 31.752
R663 VN.n10 VN.n7 24.4675
R664 VN.n14 VN.n7 24.4675
R665 VN.n15 VN.n14 24.4675
R666 VN.n16 VN.n5 24.4675
R667 VN.n20 VN.n5 24.4675
R668 VN.n21 VN.n20 24.4675
R669 VN.n23 VN.n3 24.4675
R670 VN.n27 VN.n3 24.4675
R671 VN.n28 VN.n27 24.4675
R672 VN.n33 VN.n1 24.4675
R673 VN.n34 VN.n33 24.4675
R674 VN.n52 VN.n51 24.4675
R675 VN.n51 VN.n44 24.4675
R676 VN.n47 VN.n44 24.4675
R677 VN.n65 VN.n64 24.4675
R678 VN.n64 VN.n40 24.4675
R679 VN.n60 VN.n40 24.4675
R680 VN.n58 VN.n57 24.4675
R681 VN.n57 VN.n42 24.4675
R682 VN.n53 VN.n42 24.4675
R683 VN.n71 VN.n70 24.4675
R684 VN.n70 VN.n38 24.4675
R685 VN.n35 VN.n34 23.9782
R686 VN.n72 VN.n71 23.9782
R687 VN.n10 VN.n9 16.1487
R688 VN.n22 VN.n21 16.1487
R689 VN.n47 VN.n46 16.1487
R690 VN.n59 VN.n58 16.1487
R691 VN.n23 VN.n22 8.31928
R692 VN.n60 VN.n59 8.31928
R693 VN.n48 VN.n45 2.54723
R694 VN.n11 VN.n8 2.54723
R695 VN.n73 VN.n37 0.417535
R696 VN.n36 VN.n0 0.417535
R697 VN VN.n36 0.394291
R698 VN.n69 VN.n37 0.189894
R699 VN.n69 VN.n68 0.189894
R700 VN.n68 VN.n67 0.189894
R701 VN.n67 VN.n39 0.189894
R702 VN.n63 VN.n39 0.189894
R703 VN.n63 VN.n62 0.189894
R704 VN.n62 VN.n61 0.189894
R705 VN.n61 VN.n41 0.189894
R706 VN.n56 VN.n41 0.189894
R707 VN.n56 VN.n55 0.189894
R708 VN.n55 VN.n54 0.189894
R709 VN.n54 VN.n43 0.189894
R710 VN.n50 VN.n43 0.189894
R711 VN.n50 VN.n49 0.189894
R712 VN.n49 VN.n48 0.189894
R713 VN.n12 VN.n11 0.189894
R714 VN.n13 VN.n12 0.189894
R715 VN.n13 VN.n6 0.189894
R716 VN.n17 VN.n6 0.189894
R717 VN.n18 VN.n17 0.189894
R718 VN.n19 VN.n18 0.189894
R719 VN.n19 VN.n4 0.189894
R720 VN.n24 VN.n4 0.189894
R721 VN.n25 VN.n24 0.189894
R722 VN.n26 VN.n25 0.189894
R723 VN.n26 VN.n2 0.189894
R724 VN.n30 VN.n2 0.189894
R725 VN.n31 VN.n30 0.189894
R726 VN.n32 VN.n31 0.189894
R727 VN.n32 VN.n0 0.189894
R728 VDD2.n2 VDD2.n1 89.4856
R729 VDD2.n2 VDD2.n0 89.4856
R730 VDD2 VDD2.n5 89.4827
R731 VDD2.n4 VDD2.n3 87.7479
R732 VDD2.n4 VDD2.n2 46.086
R733 VDD2.n5 VDD2.t2 4.49635
R734 VDD2.n5 VDD2.t3 4.49635
R735 VDD2.n3 VDD2.t7 4.49635
R736 VDD2.n3 VDD2.t6 4.49635
R737 VDD2.n1 VDD2.t1 4.49635
R738 VDD2.n1 VDD2.t0 4.49635
R739 VDD2.n0 VDD2.t4 4.49635
R740 VDD2.n0 VDD2.t5 4.49635
R741 VDD2 VDD2.n4 1.85179
R742 B.n625 B.n624 585
R743 B.n626 B.n73 585
R744 B.n628 B.n627 585
R745 B.n629 B.n72 585
R746 B.n631 B.n630 585
R747 B.n632 B.n71 585
R748 B.n634 B.n633 585
R749 B.n635 B.n70 585
R750 B.n637 B.n636 585
R751 B.n638 B.n69 585
R752 B.n640 B.n639 585
R753 B.n641 B.n68 585
R754 B.n643 B.n642 585
R755 B.n644 B.n67 585
R756 B.n646 B.n645 585
R757 B.n647 B.n66 585
R758 B.n649 B.n648 585
R759 B.n650 B.n65 585
R760 B.n652 B.n651 585
R761 B.n653 B.n64 585
R762 B.n655 B.n654 585
R763 B.n656 B.n63 585
R764 B.n658 B.n657 585
R765 B.n659 B.n62 585
R766 B.n661 B.n660 585
R767 B.n662 B.n61 585
R768 B.n664 B.n663 585
R769 B.n665 B.n58 585
R770 B.n668 B.n667 585
R771 B.n669 B.n57 585
R772 B.n671 B.n670 585
R773 B.n672 B.n56 585
R774 B.n674 B.n673 585
R775 B.n675 B.n55 585
R776 B.n677 B.n676 585
R777 B.n678 B.n51 585
R778 B.n680 B.n679 585
R779 B.n681 B.n50 585
R780 B.n683 B.n682 585
R781 B.n684 B.n49 585
R782 B.n686 B.n685 585
R783 B.n687 B.n48 585
R784 B.n689 B.n688 585
R785 B.n690 B.n47 585
R786 B.n692 B.n691 585
R787 B.n693 B.n46 585
R788 B.n695 B.n694 585
R789 B.n696 B.n45 585
R790 B.n698 B.n697 585
R791 B.n699 B.n44 585
R792 B.n701 B.n700 585
R793 B.n702 B.n43 585
R794 B.n704 B.n703 585
R795 B.n705 B.n42 585
R796 B.n707 B.n706 585
R797 B.n708 B.n41 585
R798 B.n710 B.n709 585
R799 B.n711 B.n40 585
R800 B.n713 B.n712 585
R801 B.n714 B.n39 585
R802 B.n716 B.n715 585
R803 B.n717 B.n38 585
R804 B.n719 B.n718 585
R805 B.n720 B.n37 585
R806 B.n722 B.n721 585
R807 B.n623 B.n74 585
R808 B.n622 B.n621 585
R809 B.n620 B.n75 585
R810 B.n619 B.n618 585
R811 B.n617 B.n76 585
R812 B.n616 B.n615 585
R813 B.n614 B.n77 585
R814 B.n613 B.n612 585
R815 B.n611 B.n78 585
R816 B.n610 B.n609 585
R817 B.n608 B.n79 585
R818 B.n607 B.n606 585
R819 B.n605 B.n80 585
R820 B.n604 B.n603 585
R821 B.n602 B.n81 585
R822 B.n601 B.n600 585
R823 B.n599 B.n82 585
R824 B.n598 B.n597 585
R825 B.n596 B.n83 585
R826 B.n595 B.n594 585
R827 B.n593 B.n84 585
R828 B.n592 B.n591 585
R829 B.n590 B.n85 585
R830 B.n589 B.n588 585
R831 B.n587 B.n86 585
R832 B.n586 B.n585 585
R833 B.n584 B.n87 585
R834 B.n583 B.n582 585
R835 B.n581 B.n88 585
R836 B.n580 B.n579 585
R837 B.n578 B.n89 585
R838 B.n577 B.n576 585
R839 B.n575 B.n90 585
R840 B.n574 B.n573 585
R841 B.n572 B.n91 585
R842 B.n571 B.n570 585
R843 B.n569 B.n92 585
R844 B.n568 B.n567 585
R845 B.n566 B.n93 585
R846 B.n565 B.n564 585
R847 B.n563 B.n94 585
R848 B.n562 B.n561 585
R849 B.n560 B.n95 585
R850 B.n559 B.n558 585
R851 B.n557 B.n96 585
R852 B.n556 B.n555 585
R853 B.n554 B.n97 585
R854 B.n553 B.n552 585
R855 B.n551 B.n98 585
R856 B.n550 B.n549 585
R857 B.n548 B.n99 585
R858 B.n547 B.n546 585
R859 B.n545 B.n100 585
R860 B.n544 B.n543 585
R861 B.n542 B.n101 585
R862 B.n541 B.n540 585
R863 B.n539 B.n102 585
R864 B.n538 B.n537 585
R865 B.n536 B.n103 585
R866 B.n535 B.n534 585
R867 B.n533 B.n104 585
R868 B.n532 B.n531 585
R869 B.n530 B.n105 585
R870 B.n529 B.n528 585
R871 B.n527 B.n106 585
R872 B.n526 B.n525 585
R873 B.n524 B.n107 585
R874 B.n523 B.n522 585
R875 B.n521 B.n108 585
R876 B.n520 B.n519 585
R877 B.n518 B.n109 585
R878 B.n517 B.n516 585
R879 B.n515 B.n110 585
R880 B.n514 B.n513 585
R881 B.n512 B.n111 585
R882 B.n511 B.n510 585
R883 B.n509 B.n112 585
R884 B.n508 B.n507 585
R885 B.n506 B.n113 585
R886 B.n505 B.n504 585
R887 B.n503 B.n114 585
R888 B.n502 B.n501 585
R889 B.n500 B.n115 585
R890 B.n499 B.n498 585
R891 B.n497 B.n116 585
R892 B.n496 B.n495 585
R893 B.n494 B.n117 585
R894 B.n493 B.n492 585
R895 B.n491 B.n118 585
R896 B.n490 B.n489 585
R897 B.n488 B.n119 585
R898 B.n487 B.n486 585
R899 B.n485 B.n120 585
R900 B.n484 B.n483 585
R901 B.n482 B.n121 585
R902 B.n481 B.n480 585
R903 B.n479 B.n122 585
R904 B.n478 B.n477 585
R905 B.n476 B.n123 585
R906 B.n475 B.n474 585
R907 B.n473 B.n124 585
R908 B.n472 B.n471 585
R909 B.n470 B.n125 585
R910 B.n469 B.n468 585
R911 B.n467 B.n126 585
R912 B.n466 B.n465 585
R913 B.n464 B.n127 585
R914 B.n463 B.n462 585
R915 B.n461 B.n128 585
R916 B.n460 B.n459 585
R917 B.n458 B.n129 585
R918 B.n457 B.n456 585
R919 B.n455 B.n130 585
R920 B.n454 B.n453 585
R921 B.n452 B.n131 585
R922 B.n451 B.n450 585
R923 B.n449 B.n132 585
R924 B.n448 B.n447 585
R925 B.n446 B.n133 585
R926 B.n445 B.n444 585
R927 B.n443 B.n134 585
R928 B.n442 B.n441 585
R929 B.n440 B.n135 585
R930 B.n439 B.n438 585
R931 B.n437 B.n136 585
R932 B.n436 B.n435 585
R933 B.n434 B.n137 585
R934 B.n433 B.n432 585
R935 B.n431 B.n138 585
R936 B.n430 B.n429 585
R937 B.n428 B.n139 585
R938 B.n427 B.n426 585
R939 B.n425 B.n140 585
R940 B.n424 B.n423 585
R941 B.n422 B.n141 585
R942 B.n421 B.n420 585
R943 B.n419 B.n142 585
R944 B.n418 B.n417 585
R945 B.n416 B.n143 585
R946 B.n315 B.n314 585
R947 B.n316 B.n177 585
R948 B.n318 B.n317 585
R949 B.n319 B.n176 585
R950 B.n321 B.n320 585
R951 B.n322 B.n175 585
R952 B.n324 B.n323 585
R953 B.n325 B.n174 585
R954 B.n327 B.n326 585
R955 B.n328 B.n173 585
R956 B.n330 B.n329 585
R957 B.n331 B.n172 585
R958 B.n333 B.n332 585
R959 B.n334 B.n171 585
R960 B.n336 B.n335 585
R961 B.n337 B.n170 585
R962 B.n339 B.n338 585
R963 B.n340 B.n169 585
R964 B.n342 B.n341 585
R965 B.n343 B.n168 585
R966 B.n345 B.n344 585
R967 B.n346 B.n167 585
R968 B.n348 B.n347 585
R969 B.n349 B.n166 585
R970 B.n351 B.n350 585
R971 B.n352 B.n165 585
R972 B.n354 B.n353 585
R973 B.n355 B.n162 585
R974 B.n358 B.n357 585
R975 B.n359 B.n161 585
R976 B.n361 B.n360 585
R977 B.n362 B.n160 585
R978 B.n364 B.n363 585
R979 B.n365 B.n159 585
R980 B.n367 B.n366 585
R981 B.n368 B.n158 585
R982 B.n373 B.n372 585
R983 B.n374 B.n157 585
R984 B.n376 B.n375 585
R985 B.n377 B.n156 585
R986 B.n379 B.n378 585
R987 B.n380 B.n155 585
R988 B.n382 B.n381 585
R989 B.n383 B.n154 585
R990 B.n385 B.n384 585
R991 B.n386 B.n153 585
R992 B.n388 B.n387 585
R993 B.n389 B.n152 585
R994 B.n391 B.n390 585
R995 B.n392 B.n151 585
R996 B.n394 B.n393 585
R997 B.n395 B.n150 585
R998 B.n397 B.n396 585
R999 B.n398 B.n149 585
R1000 B.n400 B.n399 585
R1001 B.n401 B.n148 585
R1002 B.n403 B.n402 585
R1003 B.n404 B.n147 585
R1004 B.n406 B.n405 585
R1005 B.n407 B.n146 585
R1006 B.n409 B.n408 585
R1007 B.n410 B.n145 585
R1008 B.n412 B.n411 585
R1009 B.n413 B.n144 585
R1010 B.n415 B.n414 585
R1011 B.n313 B.n178 585
R1012 B.n312 B.n311 585
R1013 B.n310 B.n179 585
R1014 B.n309 B.n308 585
R1015 B.n307 B.n180 585
R1016 B.n306 B.n305 585
R1017 B.n304 B.n181 585
R1018 B.n303 B.n302 585
R1019 B.n301 B.n182 585
R1020 B.n300 B.n299 585
R1021 B.n298 B.n183 585
R1022 B.n297 B.n296 585
R1023 B.n295 B.n184 585
R1024 B.n294 B.n293 585
R1025 B.n292 B.n185 585
R1026 B.n291 B.n290 585
R1027 B.n289 B.n186 585
R1028 B.n288 B.n287 585
R1029 B.n286 B.n187 585
R1030 B.n285 B.n284 585
R1031 B.n283 B.n188 585
R1032 B.n282 B.n281 585
R1033 B.n280 B.n189 585
R1034 B.n279 B.n278 585
R1035 B.n277 B.n190 585
R1036 B.n276 B.n275 585
R1037 B.n274 B.n191 585
R1038 B.n273 B.n272 585
R1039 B.n271 B.n192 585
R1040 B.n270 B.n269 585
R1041 B.n268 B.n193 585
R1042 B.n267 B.n266 585
R1043 B.n265 B.n194 585
R1044 B.n264 B.n263 585
R1045 B.n262 B.n195 585
R1046 B.n261 B.n260 585
R1047 B.n259 B.n196 585
R1048 B.n258 B.n257 585
R1049 B.n256 B.n197 585
R1050 B.n255 B.n254 585
R1051 B.n253 B.n198 585
R1052 B.n252 B.n251 585
R1053 B.n250 B.n199 585
R1054 B.n249 B.n248 585
R1055 B.n247 B.n200 585
R1056 B.n246 B.n245 585
R1057 B.n244 B.n201 585
R1058 B.n243 B.n242 585
R1059 B.n241 B.n202 585
R1060 B.n240 B.n239 585
R1061 B.n238 B.n203 585
R1062 B.n237 B.n236 585
R1063 B.n235 B.n204 585
R1064 B.n234 B.n233 585
R1065 B.n232 B.n205 585
R1066 B.n231 B.n230 585
R1067 B.n229 B.n206 585
R1068 B.n228 B.n227 585
R1069 B.n226 B.n207 585
R1070 B.n225 B.n224 585
R1071 B.n223 B.n208 585
R1072 B.n222 B.n221 585
R1073 B.n220 B.n209 585
R1074 B.n219 B.n218 585
R1075 B.n217 B.n210 585
R1076 B.n216 B.n215 585
R1077 B.n214 B.n211 585
R1078 B.n213 B.n212 585
R1079 B.n2 B.n0 585
R1080 B.n825 B.n1 585
R1081 B.n824 B.n823 585
R1082 B.n822 B.n3 585
R1083 B.n821 B.n820 585
R1084 B.n819 B.n4 585
R1085 B.n818 B.n817 585
R1086 B.n816 B.n5 585
R1087 B.n815 B.n814 585
R1088 B.n813 B.n6 585
R1089 B.n812 B.n811 585
R1090 B.n810 B.n7 585
R1091 B.n809 B.n808 585
R1092 B.n807 B.n8 585
R1093 B.n806 B.n805 585
R1094 B.n804 B.n9 585
R1095 B.n803 B.n802 585
R1096 B.n801 B.n10 585
R1097 B.n800 B.n799 585
R1098 B.n798 B.n11 585
R1099 B.n797 B.n796 585
R1100 B.n795 B.n12 585
R1101 B.n794 B.n793 585
R1102 B.n792 B.n13 585
R1103 B.n791 B.n790 585
R1104 B.n789 B.n14 585
R1105 B.n788 B.n787 585
R1106 B.n786 B.n15 585
R1107 B.n785 B.n784 585
R1108 B.n783 B.n16 585
R1109 B.n782 B.n781 585
R1110 B.n780 B.n17 585
R1111 B.n779 B.n778 585
R1112 B.n777 B.n18 585
R1113 B.n776 B.n775 585
R1114 B.n774 B.n19 585
R1115 B.n773 B.n772 585
R1116 B.n771 B.n20 585
R1117 B.n770 B.n769 585
R1118 B.n768 B.n21 585
R1119 B.n767 B.n766 585
R1120 B.n765 B.n22 585
R1121 B.n764 B.n763 585
R1122 B.n762 B.n23 585
R1123 B.n761 B.n760 585
R1124 B.n759 B.n24 585
R1125 B.n758 B.n757 585
R1126 B.n756 B.n25 585
R1127 B.n755 B.n754 585
R1128 B.n753 B.n26 585
R1129 B.n752 B.n751 585
R1130 B.n750 B.n27 585
R1131 B.n749 B.n748 585
R1132 B.n747 B.n28 585
R1133 B.n746 B.n745 585
R1134 B.n744 B.n29 585
R1135 B.n743 B.n742 585
R1136 B.n741 B.n30 585
R1137 B.n740 B.n739 585
R1138 B.n738 B.n31 585
R1139 B.n737 B.n736 585
R1140 B.n735 B.n32 585
R1141 B.n734 B.n733 585
R1142 B.n732 B.n33 585
R1143 B.n731 B.n730 585
R1144 B.n729 B.n34 585
R1145 B.n728 B.n727 585
R1146 B.n726 B.n35 585
R1147 B.n725 B.n724 585
R1148 B.n723 B.n36 585
R1149 B.n827 B.n826 585
R1150 B.n315 B.n178 526.135
R1151 B.n723 B.n722 526.135
R1152 B.n416 B.n415 526.135
R1153 B.n625 B.n74 526.135
R1154 B.n369 B.t11 370.454
R1155 B.n59 B.t1 370.454
R1156 B.n163 B.t8 370.452
R1157 B.n52 B.t4 370.452
R1158 B.n370 B.t10 289.774
R1159 B.n60 B.t2 289.774
R1160 B.n164 B.t7 289.774
R1161 B.n53 B.t5 289.774
R1162 B.n369 B.t9 254.862
R1163 B.n163 B.t6 254.862
R1164 B.n52 B.t3 254.862
R1165 B.n59 B.t0 254.862
R1166 B.n311 B.n178 163.367
R1167 B.n311 B.n310 163.367
R1168 B.n310 B.n309 163.367
R1169 B.n309 B.n180 163.367
R1170 B.n305 B.n180 163.367
R1171 B.n305 B.n304 163.367
R1172 B.n304 B.n303 163.367
R1173 B.n303 B.n182 163.367
R1174 B.n299 B.n182 163.367
R1175 B.n299 B.n298 163.367
R1176 B.n298 B.n297 163.367
R1177 B.n297 B.n184 163.367
R1178 B.n293 B.n184 163.367
R1179 B.n293 B.n292 163.367
R1180 B.n292 B.n291 163.367
R1181 B.n291 B.n186 163.367
R1182 B.n287 B.n186 163.367
R1183 B.n287 B.n286 163.367
R1184 B.n286 B.n285 163.367
R1185 B.n285 B.n188 163.367
R1186 B.n281 B.n188 163.367
R1187 B.n281 B.n280 163.367
R1188 B.n280 B.n279 163.367
R1189 B.n279 B.n190 163.367
R1190 B.n275 B.n190 163.367
R1191 B.n275 B.n274 163.367
R1192 B.n274 B.n273 163.367
R1193 B.n273 B.n192 163.367
R1194 B.n269 B.n192 163.367
R1195 B.n269 B.n268 163.367
R1196 B.n268 B.n267 163.367
R1197 B.n267 B.n194 163.367
R1198 B.n263 B.n194 163.367
R1199 B.n263 B.n262 163.367
R1200 B.n262 B.n261 163.367
R1201 B.n261 B.n196 163.367
R1202 B.n257 B.n196 163.367
R1203 B.n257 B.n256 163.367
R1204 B.n256 B.n255 163.367
R1205 B.n255 B.n198 163.367
R1206 B.n251 B.n198 163.367
R1207 B.n251 B.n250 163.367
R1208 B.n250 B.n249 163.367
R1209 B.n249 B.n200 163.367
R1210 B.n245 B.n200 163.367
R1211 B.n245 B.n244 163.367
R1212 B.n244 B.n243 163.367
R1213 B.n243 B.n202 163.367
R1214 B.n239 B.n202 163.367
R1215 B.n239 B.n238 163.367
R1216 B.n238 B.n237 163.367
R1217 B.n237 B.n204 163.367
R1218 B.n233 B.n204 163.367
R1219 B.n233 B.n232 163.367
R1220 B.n232 B.n231 163.367
R1221 B.n231 B.n206 163.367
R1222 B.n227 B.n206 163.367
R1223 B.n227 B.n226 163.367
R1224 B.n226 B.n225 163.367
R1225 B.n225 B.n208 163.367
R1226 B.n221 B.n208 163.367
R1227 B.n221 B.n220 163.367
R1228 B.n220 B.n219 163.367
R1229 B.n219 B.n210 163.367
R1230 B.n215 B.n210 163.367
R1231 B.n215 B.n214 163.367
R1232 B.n214 B.n213 163.367
R1233 B.n213 B.n2 163.367
R1234 B.n826 B.n2 163.367
R1235 B.n826 B.n825 163.367
R1236 B.n825 B.n824 163.367
R1237 B.n824 B.n3 163.367
R1238 B.n820 B.n3 163.367
R1239 B.n820 B.n819 163.367
R1240 B.n819 B.n818 163.367
R1241 B.n818 B.n5 163.367
R1242 B.n814 B.n5 163.367
R1243 B.n814 B.n813 163.367
R1244 B.n813 B.n812 163.367
R1245 B.n812 B.n7 163.367
R1246 B.n808 B.n7 163.367
R1247 B.n808 B.n807 163.367
R1248 B.n807 B.n806 163.367
R1249 B.n806 B.n9 163.367
R1250 B.n802 B.n9 163.367
R1251 B.n802 B.n801 163.367
R1252 B.n801 B.n800 163.367
R1253 B.n800 B.n11 163.367
R1254 B.n796 B.n11 163.367
R1255 B.n796 B.n795 163.367
R1256 B.n795 B.n794 163.367
R1257 B.n794 B.n13 163.367
R1258 B.n790 B.n13 163.367
R1259 B.n790 B.n789 163.367
R1260 B.n789 B.n788 163.367
R1261 B.n788 B.n15 163.367
R1262 B.n784 B.n15 163.367
R1263 B.n784 B.n783 163.367
R1264 B.n783 B.n782 163.367
R1265 B.n782 B.n17 163.367
R1266 B.n778 B.n17 163.367
R1267 B.n778 B.n777 163.367
R1268 B.n777 B.n776 163.367
R1269 B.n776 B.n19 163.367
R1270 B.n772 B.n19 163.367
R1271 B.n772 B.n771 163.367
R1272 B.n771 B.n770 163.367
R1273 B.n770 B.n21 163.367
R1274 B.n766 B.n21 163.367
R1275 B.n766 B.n765 163.367
R1276 B.n765 B.n764 163.367
R1277 B.n764 B.n23 163.367
R1278 B.n760 B.n23 163.367
R1279 B.n760 B.n759 163.367
R1280 B.n759 B.n758 163.367
R1281 B.n758 B.n25 163.367
R1282 B.n754 B.n25 163.367
R1283 B.n754 B.n753 163.367
R1284 B.n753 B.n752 163.367
R1285 B.n752 B.n27 163.367
R1286 B.n748 B.n27 163.367
R1287 B.n748 B.n747 163.367
R1288 B.n747 B.n746 163.367
R1289 B.n746 B.n29 163.367
R1290 B.n742 B.n29 163.367
R1291 B.n742 B.n741 163.367
R1292 B.n741 B.n740 163.367
R1293 B.n740 B.n31 163.367
R1294 B.n736 B.n31 163.367
R1295 B.n736 B.n735 163.367
R1296 B.n735 B.n734 163.367
R1297 B.n734 B.n33 163.367
R1298 B.n730 B.n33 163.367
R1299 B.n730 B.n729 163.367
R1300 B.n729 B.n728 163.367
R1301 B.n728 B.n35 163.367
R1302 B.n724 B.n35 163.367
R1303 B.n724 B.n723 163.367
R1304 B.n316 B.n315 163.367
R1305 B.n317 B.n316 163.367
R1306 B.n317 B.n176 163.367
R1307 B.n321 B.n176 163.367
R1308 B.n322 B.n321 163.367
R1309 B.n323 B.n322 163.367
R1310 B.n323 B.n174 163.367
R1311 B.n327 B.n174 163.367
R1312 B.n328 B.n327 163.367
R1313 B.n329 B.n328 163.367
R1314 B.n329 B.n172 163.367
R1315 B.n333 B.n172 163.367
R1316 B.n334 B.n333 163.367
R1317 B.n335 B.n334 163.367
R1318 B.n335 B.n170 163.367
R1319 B.n339 B.n170 163.367
R1320 B.n340 B.n339 163.367
R1321 B.n341 B.n340 163.367
R1322 B.n341 B.n168 163.367
R1323 B.n345 B.n168 163.367
R1324 B.n346 B.n345 163.367
R1325 B.n347 B.n346 163.367
R1326 B.n347 B.n166 163.367
R1327 B.n351 B.n166 163.367
R1328 B.n352 B.n351 163.367
R1329 B.n353 B.n352 163.367
R1330 B.n353 B.n162 163.367
R1331 B.n358 B.n162 163.367
R1332 B.n359 B.n358 163.367
R1333 B.n360 B.n359 163.367
R1334 B.n360 B.n160 163.367
R1335 B.n364 B.n160 163.367
R1336 B.n365 B.n364 163.367
R1337 B.n366 B.n365 163.367
R1338 B.n366 B.n158 163.367
R1339 B.n373 B.n158 163.367
R1340 B.n374 B.n373 163.367
R1341 B.n375 B.n374 163.367
R1342 B.n375 B.n156 163.367
R1343 B.n379 B.n156 163.367
R1344 B.n380 B.n379 163.367
R1345 B.n381 B.n380 163.367
R1346 B.n381 B.n154 163.367
R1347 B.n385 B.n154 163.367
R1348 B.n386 B.n385 163.367
R1349 B.n387 B.n386 163.367
R1350 B.n387 B.n152 163.367
R1351 B.n391 B.n152 163.367
R1352 B.n392 B.n391 163.367
R1353 B.n393 B.n392 163.367
R1354 B.n393 B.n150 163.367
R1355 B.n397 B.n150 163.367
R1356 B.n398 B.n397 163.367
R1357 B.n399 B.n398 163.367
R1358 B.n399 B.n148 163.367
R1359 B.n403 B.n148 163.367
R1360 B.n404 B.n403 163.367
R1361 B.n405 B.n404 163.367
R1362 B.n405 B.n146 163.367
R1363 B.n409 B.n146 163.367
R1364 B.n410 B.n409 163.367
R1365 B.n411 B.n410 163.367
R1366 B.n411 B.n144 163.367
R1367 B.n415 B.n144 163.367
R1368 B.n417 B.n416 163.367
R1369 B.n417 B.n142 163.367
R1370 B.n421 B.n142 163.367
R1371 B.n422 B.n421 163.367
R1372 B.n423 B.n422 163.367
R1373 B.n423 B.n140 163.367
R1374 B.n427 B.n140 163.367
R1375 B.n428 B.n427 163.367
R1376 B.n429 B.n428 163.367
R1377 B.n429 B.n138 163.367
R1378 B.n433 B.n138 163.367
R1379 B.n434 B.n433 163.367
R1380 B.n435 B.n434 163.367
R1381 B.n435 B.n136 163.367
R1382 B.n439 B.n136 163.367
R1383 B.n440 B.n439 163.367
R1384 B.n441 B.n440 163.367
R1385 B.n441 B.n134 163.367
R1386 B.n445 B.n134 163.367
R1387 B.n446 B.n445 163.367
R1388 B.n447 B.n446 163.367
R1389 B.n447 B.n132 163.367
R1390 B.n451 B.n132 163.367
R1391 B.n452 B.n451 163.367
R1392 B.n453 B.n452 163.367
R1393 B.n453 B.n130 163.367
R1394 B.n457 B.n130 163.367
R1395 B.n458 B.n457 163.367
R1396 B.n459 B.n458 163.367
R1397 B.n459 B.n128 163.367
R1398 B.n463 B.n128 163.367
R1399 B.n464 B.n463 163.367
R1400 B.n465 B.n464 163.367
R1401 B.n465 B.n126 163.367
R1402 B.n469 B.n126 163.367
R1403 B.n470 B.n469 163.367
R1404 B.n471 B.n470 163.367
R1405 B.n471 B.n124 163.367
R1406 B.n475 B.n124 163.367
R1407 B.n476 B.n475 163.367
R1408 B.n477 B.n476 163.367
R1409 B.n477 B.n122 163.367
R1410 B.n481 B.n122 163.367
R1411 B.n482 B.n481 163.367
R1412 B.n483 B.n482 163.367
R1413 B.n483 B.n120 163.367
R1414 B.n487 B.n120 163.367
R1415 B.n488 B.n487 163.367
R1416 B.n489 B.n488 163.367
R1417 B.n489 B.n118 163.367
R1418 B.n493 B.n118 163.367
R1419 B.n494 B.n493 163.367
R1420 B.n495 B.n494 163.367
R1421 B.n495 B.n116 163.367
R1422 B.n499 B.n116 163.367
R1423 B.n500 B.n499 163.367
R1424 B.n501 B.n500 163.367
R1425 B.n501 B.n114 163.367
R1426 B.n505 B.n114 163.367
R1427 B.n506 B.n505 163.367
R1428 B.n507 B.n506 163.367
R1429 B.n507 B.n112 163.367
R1430 B.n511 B.n112 163.367
R1431 B.n512 B.n511 163.367
R1432 B.n513 B.n512 163.367
R1433 B.n513 B.n110 163.367
R1434 B.n517 B.n110 163.367
R1435 B.n518 B.n517 163.367
R1436 B.n519 B.n518 163.367
R1437 B.n519 B.n108 163.367
R1438 B.n523 B.n108 163.367
R1439 B.n524 B.n523 163.367
R1440 B.n525 B.n524 163.367
R1441 B.n525 B.n106 163.367
R1442 B.n529 B.n106 163.367
R1443 B.n530 B.n529 163.367
R1444 B.n531 B.n530 163.367
R1445 B.n531 B.n104 163.367
R1446 B.n535 B.n104 163.367
R1447 B.n536 B.n535 163.367
R1448 B.n537 B.n536 163.367
R1449 B.n537 B.n102 163.367
R1450 B.n541 B.n102 163.367
R1451 B.n542 B.n541 163.367
R1452 B.n543 B.n542 163.367
R1453 B.n543 B.n100 163.367
R1454 B.n547 B.n100 163.367
R1455 B.n548 B.n547 163.367
R1456 B.n549 B.n548 163.367
R1457 B.n549 B.n98 163.367
R1458 B.n553 B.n98 163.367
R1459 B.n554 B.n553 163.367
R1460 B.n555 B.n554 163.367
R1461 B.n555 B.n96 163.367
R1462 B.n559 B.n96 163.367
R1463 B.n560 B.n559 163.367
R1464 B.n561 B.n560 163.367
R1465 B.n561 B.n94 163.367
R1466 B.n565 B.n94 163.367
R1467 B.n566 B.n565 163.367
R1468 B.n567 B.n566 163.367
R1469 B.n567 B.n92 163.367
R1470 B.n571 B.n92 163.367
R1471 B.n572 B.n571 163.367
R1472 B.n573 B.n572 163.367
R1473 B.n573 B.n90 163.367
R1474 B.n577 B.n90 163.367
R1475 B.n578 B.n577 163.367
R1476 B.n579 B.n578 163.367
R1477 B.n579 B.n88 163.367
R1478 B.n583 B.n88 163.367
R1479 B.n584 B.n583 163.367
R1480 B.n585 B.n584 163.367
R1481 B.n585 B.n86 163.367
R1482 B.n589 B.n86 163.367
R1483 B.n590 B.n589 163.367
R1484 B.n591 B.n590 163.367
R1485 B.n591 B.n84 163.367
R1486 B.n595 B.n84 163.367
R1487 B.n596 B.n595 163.367
R1488 B.n597 B.n596 163.367
R1489 B.n597 B.n82 163.367
R1490 B.n601 B.n82 163.367
R1491 B.n602 B.n601 163.367
R1492 B.n603 B.n602 163.367
R1493 B.n603 B.n80 163.367
R1494 B.n607 B.n80 163.367
R1495 B.n608 B.n607 163.367
R1496 B.n609 B.n608 163.367
R1497 B.n609 B.n78 163.367
R1498 B.n613 B.n78 163.367
R1499 B.n614 B.n613 163.367
R1500 B.n615 B.n614 163.367
R1501 B.n615 B.n76 163.367
R1502 B.n619 B.n76 163.367
R1503 B.n620 B.n619 163.367
R1504 B.n621 B.n620 163.367
R1505 B.n621 B.n74 163.367
R1506 B.n722 B.n37 163.367
R1507 B.n718 B.n37 163.367
R1508 B.n718 B.n717 163.367
R1509 B.n717 B.n716 163.367
R1510 B.n716 B.n39 163.367
R1511 B.n712 B.n39 163.367
R1512 B.n712 B.n711 163.367
R1513 B.n711 B.n710 163.367
R1514 B.n710 B.n41 163.367
R1515 B.n706 B.n41 163.367
R1516 B.n706 B.n705 163.367
R1517 B.n705 B.n704 163.367
R1518 B.n704 B.n43 163.367
R1519 B.n700 B.n43 163.367
R1520 B.n700 B.n699 163.367
R1521 B.n699 B.n698 163.367
R1522 B.n698 B.n45 163.367
R1523 B.n694 B.n45 163.367
R1524 B.n694 B.n693 163.367
R1525 B.n693 B.n692 163.367
R1526 B.n692 B.n47 163.367
R1527 B.n688 B.n47 163.367
R1528 B.n688 B.n687 163.367
R1529 B.n687 B.n686 163.367
R1530 B.n686 B.n49 163.367
R1531 B.n682 B.n49 163.367
R1532 B.n682 B.n681 163.367
R1533 B.n681 B.n680 163.367
R1534 B.n680 B.n51 163.367
R1535 B.n676 B.n51 163.367
R1536 B.n676 B.n675 163.367
R1537 B.n675 B.n674 163.367
R1538 B.n674 B.n56 163.367
R1539 B.n670 B.n56 163.367
R1540 B.n670 B.n669 163.367
R1541 B.n669 B.n668 163.367
R1542 B.n668 B.n58 163.367
R1543 B.n663 B.n58 163.367
R1544 B.n663 B.n662 163.367
R1545 B.n662 B.n661 163.367
R1546 B.n661 B.n62 163.367
R1547 B.n657 B.n62 163.367
R1548 B.n657 B.n656 163.367
R1549 B.n656 B.n655 163.367
R1550 B.n655 B.n64 163.367
R1551 B.n651 B.n64 163.367
R1552 B.n651 B.n650 163.367
R1553 B.n650 B.n649 163.367
R1554 B.n649 B.n66 163.367
R1555 B.n645 B.n66 163.367
R1556 B.n645 B.n644 163.367
R1557 B.n644 B.n643 163.367
R1558 B.n643 B.n68 163.367
R1559 B.n639 B.n68 163.367
R1560 B.n639 B.n638 163.367
R1561 B.n638 B.n637 163.367
R1562 B.n637 B.n70 163.367
R1563 B.n633 B.n70 163.367
R1564 B.n633 B.n632 163.367
R1565 B.n632 B.n631 163.367
R1566 B.n631 B.n72 163.367
R1567 B.n627 B.n72 163.367
R1568 B.n627 B.n626 163.367
R1569 B.n626 B.n625 163.367
R1570 B.n370 B.n369 80.6793
R1571 B.n164 B.n163 80.6793
R1572 B.n53 B.n52 80.6793
R1573 B.n60 B.n59 80.6793
R1574 B.n371 B.n370 59.5399
R1575 B.n356 B.n164 59.5399
R1576 B.n54 B.n53 59.5399
R1577 B.n666 B.n60 59.5399
R1578 B.n721 B.n36 34.1859
R1579 B.n624 B.n623 34.1859
R1580 B.n414 B.n143 34.1859
R1581 B.n314 B.n313 34.1859
R1582 B B.n827 18.0485
R1583 B.n721 B.n720 10.6151
R1584 B.n720 B.n719 10.6151
R1585 B.n719 B.n38 10.6151
R1586 B.n715 B.n38 10.6151
R1587 B.n715 B.n714 10.6151
R1588 B.n714 B.n713 10.6151
R1589 B.n713 B.n40 10.6151
R1590 B.n709 B.n40 10.6151
R1591 B.n709 B.n708 10.6151
R1592 B.n708 B.n707 10.6151
R1593 B.n707 B.n42 10.6151
R1594 B.n703 B.n42 10.6151
R1595 B.n703 B.n702 10.6151
R1596 B.n702 B.n701 10.6151
R1597 B.n701 B.n44 10.6151
R1598 B.n697 B.n44 10.6151
R1599 B.n697 B.n696 10.6151
R1600 B.n696 B.n695 10.6151
R1601 B.n695 B.n46 10.6151
R1602 B.n691 B.n46 10.6151
R1603 B.n691 B.n690 10.6151
R1604 B.n690 B.n689 10.6151
R1605 B.n689 B.n48 10.6151
R1606 B.n685 B.n48 10.6151
R1607 B.n685 B.n684 10.6151
R1608 B.n684 B.n683 10.6151
R1609 B.n683 B.n50 10.6151
R1610 B.n679 B.n678 10.6151
R1611 B.n678 B.n677 10.6151
R1612 B.n677 B.n55 10.6151
R1613 B.n673 B.n55 10.6151
R1614 B.n673 B.n672 10.6151
R1615 B.n672 B.n671 10.6151
R1616 B.n671 B.n57 10.6151
R1617 B.n667 B.n57 10.6151
R1618 B.n665 B.n664 10.6151
R1619 B.n664 B.n61 10.6151
R1620 B.n660 B.n61 10.6151
R1621 B.n660 B.n659 10.6151
R1622 B.n659 B.n658 10.6151
R1623 B.n658 B.n63 10.6151
R1624 B.n654 B.n63 10.6151
R1625 B.n654 B.n653 10.6151
R1626 B.n653 B.n652 10.6151
R1627 B.n652 B.n65 10.6151
R1628 B.n648 B.n65 10.6151
R1629 B.n648 B.n647 10.6151
R1630 B.n647 B.n646 10.6151
R1631 B.n646 B.n67 10.6151
R1632 B.n642 B.n67 10.6151
R1633 B.n642 B.n641 10.6151
R1634 B.n641 B.n640 10.6151
R1635 B.n640 B.n69 10.6151
R1636 B.n636 B.n69 10.6151
R1637 B.n636 B.n635 10.6151
R1638 B.n635 B.n634 10.6151
R1639 B.n634 B.n71 10.6151
R1640 B.n630 B.n71 10.6151
R1641 B.n630 B.n629 10.6151
R1642 B.n629 B.n628 10.6151
R1643 B.n628 B.n73 10.6151
R1644 B.n624 B.n73 10.6151
R1645 B.n418 B.n143 10.6151
R1646 B.n419 B.n418 10.6151
R1647 B.n420 B.n419 10.6151
R1648 B.n420 B.n141 10.6151
R1649 B.n424 B.n141 10.6151
R1650 B.n425 B.n424 10.6151
R1651 B.n426 B.n425 10.6151
R1652 B.n426 B.n139 10.6151
R1653 B.n430 B.n139 10.6151
R1654 B.n431 B.n430 10.6151
R1655 B.n432 B.n431 10.6151
R1656 B.n432 B.n137 10.6151
R1657 B.n436 B.n137 10.6151
R1658 B.n437 B.n436 10.6151
R1659 B.n438 B.n437 10.6151
R1660 B.n438 B.n135 10.6151
R1661 B.n442 B.n135 10.6151
R1662 B.n443 B.n442 10.6151
R1663 B.n444 B.n443 10.6151
R1664 B.n444 B.n133 10.6151
R1665 B.n448 B.n133 10.6151
R1666 B.n449 B.n448 10.6151
R1667 B.n450 B.n449 10.6151
R1668 B.n450 B.n131 10.6151
R1669 B.n454 B.n131 10.6151
R1670 B.n455 B.n454 10.6151
R1671 B.n456 B.n455 10.6151
R1672 B.n456 B.n129 10.6151
R1673 B.n460 B.n129 10.6151
R1674 B.n461 B.n460 10.6151
R1675 B.n462 B.n461 10.6151
R1676 B.n462 B.n127 10.6151
R1677 B.n466 B.n127 10.6151
R1678 B.n467 B.n466 10.6151
R1679 B.n468 B.n467 10.6151
R1680 B.n468 B.n125 10.6151
R1681 B.n472 B.n125 10.6151
R1682 B.n473 B.n472 10.6151
R1683 B.n474 B.n473 10.6151
R1684 B.n474 B.n123 10.6151
R1685 B.n478 B.n123 10.6151
R1686 B.n479 B.n478 10.6151
R1687 B.n480 B.n479 10.6151
R1688 B.n480 B.n121 10.6151
R1689 B.n484 B.n121 10.6151
R1690 B.n485 B.n484 10.6151
R1691 B.n486 B.n485 10.6151
R1692 B.n486 B.n119 10.6151
R1693 B.n490 B.n119 10.6151
R1694 B.n491 B.n490 10.6151
R1695 B.n492 B.n491 10.6151
R1696 B.n492 B.n117 10.6151
R1697 B.n496 B.n117 10.6151
R1698 B.n497 B.n496 10.6151
R1699 B.n498 B.n497 10.6151
R1700 B.n498 B.n115 10.6151
R1701 B.n502 B.n115 10.6151
R1702 B.n503 B.n502 10.6151
R1703 B.n504 B.n503 10.6151
R1704 B.n504 B.n113 10.6151
R1705 B.n508 B.n113 10.6151
R1706 B.n509 B.n508 10.6151
R1707 B.n510 B.n509 10.6151
R1708 B.n510 B.n111 10.6151
R1709 B.n514 B.n111 10.6151
R1710 B.n515 B.n514 10.6151
R1711 B.n516 B.n515 10.6151
R1712 B.n516 B.n109 10.6151
R1713 B.n520 B.n109 10.6151
R1714 B.n521 B.n520 10.6151
R1715 B.n522 B.n521 10.6151
R1716 B.n522 B.n107 10.6151
R1717 B.n526 B.n107 10.6151
R1718 B.n527 B.n526 10.6151
R1719 B.n528 B.n527 10.6151
R1720 B.n528 B.n105 10.6151
R1721 B.n532 B.n105 10.6151
R1722 B.n533 B.n532 10.6151
R1723 B.n534 B.n533 10.6151
R1724 B.n534 B.n103 10.6151
R1725 B.n538 B.n103 10.6151
R1726 B.n539 B.n538 10.6151
R1727 B.n540 B.n539 10.6151
R1728 B.n540 B.n101 10.6151
R1729 B.n544 B.n101 10.6151
R1730 B.n545 B.n544 10.6151
R1731 B.n546 B.n545 10.6151
R1732 B.n546 B.n99 10.6151
R1733 B.n550 B.n99 10.6151
R1734 B.n551 B.n550 10.6151
R1735 B.n552 B.n551 10.6151
R1736 B.n552 B.n97 10.6151
R1737 B.n556 B.n97 10.6151
R1738 B.n557 B.n556 10.6151
R1739 B.n558 B.n557 10.6151
R1740 B.n558 B.n95 10.6151
R1741 B.n562 B.n95 10.6151
R1742 B.n563 B.n562 10.6151
R1743 B.n564 B.n563 10.6151
R1744 B.n564 B.n93 10.6151
R1745 B.n568 B.n93 10.6151
R1746 B.n569 B.n568 10.6151
R1747 B.n570 B.n569 10.6151
R1748 B.n570 B.n91 10.6151
R1749 B.n574 B.n91 10.6151
R1750 B.n575 B.n574 10.6151
R1751 B.n576 B.n575 10.6151
R1752 B.n576 B.n89 10.6151
R1753 B.n580 B.n89 10.6151
R1754 B.n581 B.n580 10.6151
R1755 B.n582 B.n581 10.6151
R1756 B.n582 B.n87 10.6151
R1757 B.n586 B.n87 10.6151
R1758 B.n587 B.n586 10.6151
R1759 B.n588 B.n587 10.6151
R1760 B.n588 B.n85 10.6151
R1761 B.n592 B.n85 10.6151
R1762 B.n593 B.n592 10.6151
R1763 B.n594 B.n593 10.6151
R1764 B.n594 B.n83 10.6151
R1765 B.n598 B.n83 10.6151
R1766 B.n599 B.n598 10.6151
R1767 B.n600 B.n599 10.6151
R1768 B.n600 B.n81 10.6151
R1769 B.n604 B.n81 10.6151
R1770 B.n605 B.n604 10.6151
R1771 B.n606 B.n605 10.6151
R1772 B.n606 B.n79 10.6151
R1773 B.n610 B.n79 10.6151
R1774 B.n611 B.n610 10.6151
R1775 B.n612 B.n611 10.6151
R1776 B.n612 B.n77 10.6151
R1777 B.n616 B.n77 10.6151
R1778 B.n617 B.n616 10.6151
R1779 B.n618 B.n617 10.6151
R1780 B.n618 B.n75 10.6151
R1781 B.n622 B.n75 10.6151
R1782 B.n623 B.n622 10.6151
R1783 B.n314 B.n177 10.6151
R1784 B.n318 B.n177 10.6151
R1785 B.n319 B.n318 10.6151
R1786 B.n320 B.n319 10.6151
R1787 B.n320 B.n175 10.6151
R1788 B.n324 B.n175 10.6151
R1789 B.n325 B.n324 10.6151
R1790 B.n326 B.n325 10.6151
R1791 B.n326 B.n173 10.6151
R1792 B.n330 B.n173 10.6151
R1793 B.n331 B.n330 10.6151
R1794 B.n332 B.n331 10.6151
R1795 B.n332 B.n171 10.6151
R1796 B.n336 B.n171 10.6151
R1797 B.n337 B.n336 10.6151
R1798 B.n338 B.n337 10.6151
R1799 B.n338 B.n169 10.6151
R1800 B.n342 B.n169 10.6151
R1801 B.n343 B.n342 10.6151
R1802 B.n344 B.n343 10.6151
R1803 B.n344 B.n167 10.6151
R1804 B.n348 B.n167 10.6151
R1805 B.n349 B.n348 10.6151
R1806 B.n350 B.n349 10.6151
R1807 B.n350 B.n165 10.6151
R1808 B.n354 B.n165 10.6151
R1809 B.n355 B.n354 10.6151
R1810 B.n357 B.n161 10.6151
R1811 B.n361 B.n161 10.6151
R1812 B.n362 B.n361 10.6151
R1813 B.n363 B.n362 10.6151
R1814 B.n363 B.n159 10.6151
R1815 B.n367 B.n159 10.6151
R1816 B.n368 B.n367 10.6151
R1817 B.n372 B.n368 10.6151
R1818 B.n376 B.n157 10.6151
R1819 B.n377 B.n376 10.6151
R1820 B.n378 B.n377 10.6151
R1821 B.n378 B.n155 10.6151
R1822 B.n382 B.n155 10.6151
R1823 B.n383 B.n382 10.6151
R1824 B.n384 B.n383 10.6151
R1825 B.n384 B.n153 10.6151
R1826 B.n388 B.n153 10.6151
R1827 B.n389 B.n388 10.6151
R1828 B.n390 B.n389 10.6151
R1829 B.n390 B.n151 10.6151
R1830 B.n394 B.n151 10.6151
R1831 B.n395 B.n394 10.6151
R1832 B.n396 B.n395 10.6151
R1833 B.n396 B.n149 10.6151
R1834 B.n400 B.n149 10.6151
R1835 B.n401 B.n400 10.6151
R1836 B.n402 B.n401 10.6151
R1837 B.n402 B.n147 10.6151
R1838 B.n406 B.n147 10.6151
R1839 B.n407 B.n406 10.6151
R1840 B.n408 B.n407 10.6151
R1841 B.n408 B.n145 10.6151
R1842 B.n412 B.n145 10.6151
R1843 B.n413 B.n412 10.6151
R1844 B.n414 B.n413 10.6151
R1845 B.n313 B.n312 10.6151
R1846 B.n312 B.n179 10.6151
R1847 B.n308 B.n179 10.6151
R1848 B.n308 B.n307 10.6151
R1849 B.n307 B.n306 10.6151
R1850 B.n306 B.n181 10.6151
R1851 B.n302 B.n181 10.6151
R1852 B.n302 B.n301 10.6151
R1853 B.n301 B.n300 10.6151
R1854 B.n300 B.n183 10.6151
R1855 B.n296 B.n183 10.6151
R1856 B.n296 B.n295 10.6151
R1857 B.n295 B.n294 10.6151
R1858 B.n294 B.n185 10.6151
R1859 B.n290 B.n185 10.6151
R1860 B.n290 B.n289 10.6151
R1861 B.n289 B.n288 10.6151
R1862 B.n288 B.n187 10.6151
R1863 B.n284 B.n187 10.6151
R1864 B.n284 B.n283 10.6151
R1865 B.n283 B.n282 10.6151
R1866 B.n282 B.n189 10.6151
R1867 B.n278 B.n189 10.6151
R1868 B.n278 B.n277 10.6151
R1869 B.n277 B.n276 10.6151
R1870 B.n276 B.n191 10.6151
R1871 B.n272 B.n191 10.6151
R1872 B.n272 B.n271 10.6151
R1873 B.n271 B.n270 10.6151
R1874 B.n270 B.n193 10.6151
R1875 B.n266 B.n193 10.6151
R1876 B.n266 B.n265 10.6151
R1877 B.n265 B.n264 10.6151
R1878 B.n264 B.n195 10.6151
R1879 B.n260 B.n195 10.6151
R1880 B.n260 B.n259 10.6151
R1881 B.n259 B.n258 10.6151
R1882 B.n258 B.n197 10.6151
R1883 B.n254 B.n197 10.6151
R1884 B.n254 B.n253 10.6151
R1885 B.n253 B.n252 10.6151
R1886 B.n252 B.n199 10.6151
R1887 B.n248 B.n199 10.6151
R1888 B.n248 B.n247 10.6151
R1889 B.n247 B.n246 10.6151
R1890 B.n246 B.n201 10.6151
R1891 B.n242 B.n201 10.6151
R1892 B.n242 B.n241 10.6151
R1893 B.n241 B.n240 10.6151
R1894 B.n240 B.n203 10.6151
R1895 B.n236 B.n203 10.6151
R1896 B.n236 B.n235 10.6151
R1897 B.n235 B.n234 10.6151
R1898 B.n234 B.n205 10.6151
R1899 B.n230 B.n205 10.6151
R1900 B.n230 B.n229 10.6151
R1901 B.n229 B.n228 10.6151
R1902 B.n228 B.n207 10.6151
R1903 B.n224 B.n207 10.6151
R1904 B.n224 B.n223 10.6151
R1905 B.n223 B.n222 10.6151
R1906 B.n222 B.n209 10.6151
R1907 B.n218 B.n209 10.6151
R1908 B.n218 B.n217 10.6151
R1909 B.n217 B.n216 10.6151
R1910 B.n216 B.n211 10.6151
R1911 B.n212 B.n211 10.6151
R1912 B.n212 B.n0 10.6151
R1913 B.n823 B.n1 10.6151
R1914 B.n823 B.n822 10.6151
R1915 B.n822 B.n821 10.6151
R1916 B.n821 B.n4 10.6151
R1917 B.n817 B.n4 10.6151
R1918 B.n817 B.n816 10.6151
R1919 B.n816 B.n815 10.6151
R1920 B.n815 B.n6 10.6151
R1921 B.n811 B.n6 10.6151
R1922 B.n811 B.n810 10.6151
R1923 B.n810 B.n809 10.6151
R1924 B.n809 B.n8 10.6151
R1925 B.n805 B.n8 10.6151
R1926 B.n805 B.n804 10.6151
R1927 B.n804 B.n803 10.6151
R1928 B.n803 B.n10 10.6151
R1929 B.n799 B.n10 10.6151
R1930 B.n799 B.n798 10.6151
R1931 B.n798 B.n797 10.6151
R1932 B.n797 B.n12 10.6151
R1933 B.n793 B.n12 10.6151
R1934 B.n793 B.n792 10.6151
R1935 B.n792 B.n791 10.6151
R1936 B.n791 B.n14 10.6151
R1937 B.n787 B.n14 10.6151
R1938 B.n787 B.n786 10.6151
R1939 B.n786 B.n785 10.6151
R1940 B.n785 B.n16 10.6151
R1941 B.n781 B.n16 10.6151
R1942 B.n781 B.n780 10.6151
R1943 B.n780 B.n779 10.6151
R1944 B.n779 B.n18 10.6151
R1945 B.n775 B.n18 10.6151
R1946 B.n775 B.n774 10.6151
R1947 B.n774 B.n773 10.6151
R1948 B.n773 B.n20 10.6151
R1949 B.n769 B.n20 10.6151
R1950 B.n769 B.n768 10.6151
R1951 B.n768 B.n767 10.6151
R1952 B.n767 B.n22 10.6151
R1953 B.n763 B.n22 10.6151
R1954 B.n763 B.n762 10.6151
R1955 B.n762 B.n761 10.6151
R1956 B.n761 B.n24 10.6151
R1957 B.n757 B.n24 10.6151
R1958 B.n757 B.n756 10.6151
R1959 B.n756 B.n755 10.6151
R1960 B.n755 B.n26 10.6151
R1961 B.n751 B.n26 10.6151
R1962 B.n751 B.n750 10.6151
R1963 B.n750 B.n749 10.6151
R1964 B.n749 B.n28 10.6151
R1965 B.n745 B.n28 10.6151
R1966 B.n745 B.n744 10.6151
R1967 B.n744 B.n743 10.6151
R1968 B.n743 B.n30 10.6151
R1969 B.n739 B.n30 10.6151
R1970 B.n739 B.n738 10.6151
R1971 B.n738 B.n737 10.6151
R1972 B.n737 B.n32 10.6151
R1973 B.n733 B.n32 10.6151
R1974 B.n733 B.n732 10.6151
R1975 B.n732 B.n731 10.6151
R1976 B.n731 B.n34 10.6151
R1977 B.n727 B.n34 10.6151
R1978 B.n727 B.n726 10.6151
R1979 B.n726 B.n725 10.6151
R1980 B.n725 B.n36 10.6151
R1981 B.n679 B.n54 6.5566
R1982 B.n667 B.n666 6.5566
R1983 B.n357 B.n356 6.5566
R1984 B.n372 B.n371 6.5566
R1985 B.n54 B.n50 4.05904
R1986 B.n666 B.n665 4.05904
R1987 B.n356 B.n355 4.05904
R1988 B.n371 B.n157 4.05904
R1989 B.n827 B.n0 2.81026
R1990 B.n827 B.n1 2.81026
C0 VN VDD2 5.77426f
C1 B VDD2 2.03141f
C2 VDD2 VTAIL 7.36846f
C3 w_n5130_n2414# VDD2 2.38572f
C4 VDD1 VDD2 2.41499f
C5 VP VDD2 0.650422f
C6 VN B 1.45543f
C7 VN VTAIL 6.81044f
C8 w_n5130_n2414# VN 10.699f
C9 VDD1 VN 0.153818f
C10 B VTAIL 3.82758f
C11 w_n5130_n2414# B 10.662999f
C12 VDD1 B 1.89668f
C13 w_n5130_n2414# VTAIL 3.28826f
C14 VN VP 8.28644f
C15 VDD1 VTAIL 7.30579f
C16 w_n5130_n2414# VDD1 2.21941f
C17 VP B 2.58447f
C18 VP VTAIL 6.82455f
C19 w_n5130_n2414# VP 11.368599f
C20 VDD1 VP 6.26885f
C21 VDD2 VSUBS 2.489532f
C22 VDD1 VSUBS 3.19056f
C23 VTAIL VSUBS 1.375722f
C24 VN VSUBS 8.414491f
C25 VP VSUBS 4.703552f
C26 B VSUBS 5.972622f
C27 w_n5130_n2414# VSUBS 0.153962p
C28 B.n0 VSUBS 0.006048f
C29 B.n1 VSUBS 0.006048f
C30 B.n2 VSUBS 0.009564f
C31 B.n3 VSUBS 0.009564f
C32 B.n4 VSUBS 0.009564f
C33 B.n5 VSUBS 0.009564f
C34 B.n6 VSUBS 0.009564f
C35 B.n7 VSUBS 0.009564f
C36 B.n8 VSUBS 0.009564f
C37 B.n9 VSUBS 0.009564f
C38 B.n10 VSUBS 0.009564f
C39 B.n11 VSUBS 0.009564f
C40 B.n12 VSUBS 0.009564f
C41 B.n13 VSUBS 0.009564f
C42 B.n14 VSUBS 0.009564f
C43 B.n15 VSUBS 0.009564f
C44 B.n16 VSUBS 0.009564f
C45 B.n17 VSUBS 0.009564f
C46 B.n18 VSUBS 0.009564f
C47 B.n19 VSUBS 0.009564f
C48 B.n20 VSUBS 0.009564f
C49 B.n21 VSUBS 0.009564f
C50 B.n22 VSUBS 0.009564f
C51 B.n23 VSUBS 0.009564f
C52 B.n24 VSUBS 0.009564f
C53 B.n25 VSUBS 0.009564f
C54 B.n26 VSUBS 0.009564f
C55 B.n27 VSUBS 0.009564f
C56 B.n28 VSUBS 0.009564f
C57 B.n29 VSUBS 0.009564f
C58 B.n30 VSUBS 0.009564f
C59 B.n31 VSUBS 0.009564f
C60 B.n32 VSUBS 0.009564f
C61 B.n33 VSUBS 0.009564f
C62 B.n34 VSUBS 0.009564f
C63 B.n35 VSUBS 0.009564f
C64 B.n36 VSUBS 0.022184f
C65 B.n37 VSUBS 0.009564f
C66 B.n38 VSUBS 0.009564f
C67 B.n39 VSUBS 0.009564f
C68 B.n40 VSUBS 0.009564f
C69 B.n41 VSUBS 0.009564f
C70 B.n42 VSUBS 0.009564f
C71 B.n43 VSUBS 0.009564f
C72 B.n44 VSUBS 0.009564f
C73 B.n45 VSUBS 0.009564f
C74 B.n46 VSUBS 0.009564f
C75 B.n47 VSUBS 0.009564f
C76 B.n48 VSUBS 0.009564f
C77 B.n49 VSUBS 0.009564f
C78 B.n50 VSUBS 0.00661f
C79 B.n51 VSUBS 0.009564f
C80 B.t5 VSUBS 0.152521f
C81 B.t4 VSUBS 0.20426f
C82 B.t3 VSUBS 1.80674f
C83 B.n52 VSUBS 0.333512f
C84 B.n53 VSUBS 0.251215f
C85 B.n54 VSUBS 0.022159f
C86 B.n55 VSUBS 0.009564f
C87 B.n56 VSUBS 0.009564f
C88 B.n57 VSUBS 0.009564f
C89 B.n58 VSUBS 0.009564f
C90 B.t2 VSUBS 0.152524f
C91 B.t1 VSUBS 0.204263f
C92 B.t0 VSUBS 1.80674f
C93 B.n59 VSUBS 0.33351f
C94 B.n60 VSUBS 0.251212f
C95 B.n61 VSUBS 0.009564f
C96 B.n62 VSUBS 0.009564f
C97 B.n63 VSUBS 0.009564f
C98 B.n64 VSUBS 0.009564f
C99 B.n65 VSUBS 0.009564f
C100 B.n66 VSUBS 0.009564f
C101 B.n67 VSUBS 0.009564f
C102 B.n68 VSUBS 0.009564f
C103 B.n69 VSUBS 0.009564f
C104 B.n70 VSUBS 0.009564f
C105 B.n71 VSUBS 0.009564f
C106 B.n72 VSUBS 0.009564f
C107 B.n73 VSUBS 0.009564f
C108 B.n74 VSUBS 0.022184f
C109 B.n75 VSUBS 0.009564f
C110 B.n76 VSUBS 0.009564f
C111 B.n77 VSUBS 0.009564f
C112 B.n78 VSUBS 0.009564f
C113 B.n79 VSUBS 0.009564f
C114 B.n80 VSUBS 0.009564f
C115 B.n81 VSUBS 0.009564f
C116 B.n82 VSUBS 0.009564f
C117 B.n83 VSUBS 0.009564f
C118 B.n84 VSUBS 0.009564f
C119 B.n85 VSUBS 0.009564f
C120 B.n86 VSUBS 0.009564f
C121 B.n87 VSUBS 0.009564f
C122 B.n88 VSUBS 0.009564f
C123 B.n89 VSUBS 0.009564f
C124 B.n90 VSUBS 0.009564f
C125 B.n91 VSUBS 0.009564f
C126 B.n92 VSUBS 0.009564f
C127 B.n93 VSUBS 0.009564f
C128 B.n94 VSUBS 0.009564f
C129 B.n95 VSUBS 0.009564f
C130 B.n96 VSUBS 0.009564f
C131 B.n97 VSUBS 0.009564f
C132 B.n98 VSUBS 0.009564f
C133 B.n99 VSUBS 0.009564f
C134 B.n100 VSUBS 0.009564f
C135 B.n101 VSUBS 0.009564f
C136 B.n102 VSUBS 0.009564f
C137 B.n103 VSUBS 0.009564f
C138 B.n104 VSUBS 0.009564f
C139 B.n105 VSUBS 0.009564f
C140 B.n106 VSUBS 0.009564f
C141 B.n107 VSUBS 0.009564f
C142 B.n108 VSUBS 0.009564f
C143 B.n109 VSUBS 0.009564f
C144 B.n110 VSUBS 0.009564f
C145 B.n111 VSUBS 0.009564f
C146 B.n112 VSUBS 0.009564f
C147 B.n113 VSUBS 0.009564f
C148 B.n114 VSUBS 0.009564f
C149 B.n115 VSUBS 0.009564f
C150 B.n116 VSUBS 0.009564f
C151 B.n117 VSUBS 0.009564f
C152 B.n118 VSUBS 0.009564f
C153 B.n119 VSUBS 0.009564f
C154 B.n120 VSUBS 0.009564f
C155 B.n121 VSUBS 0.009564f
C156 B.n122 VSUBS 0.009564f
C157 B.n123 VSUBS 0.009564f
C158 B.n124 VSUBS 0.009564f
C159 B.n125 VSUBS 0.009564f
C160 B.n126 VSUBS 0.009564f
C161 B.n127 VSUBS 0.009564f
C162 B.n128 VSUBS 0.009564f
C163 B.n129 VSUBS 0.009564f
C164 B.n130 VSUBS 0.009564f
C165 B.n131 VSUBS 0.009564f
C166 B.n132 VSUBS 0.009564f
C167 B.n133 VSUBS 0.009564f
C168 B.n134 VSUBS 0.009564f
C169 B.n135 VSUBS 0.009564f
C170 B.n136 VSUBS 0.009564f
C171 B.n137 VSUBS 0.009564f
C172 B.n138 VSUBS 0.009564f
C173 B.n139 VSUBS 0.009564f
C174 B.n140 VSUBS 0.009564f
C175 B.n141 VSUBS 0.009564f
C176 B.n142 VSUBS 0.009564f
C177 B.n143 VSUBS 0.022184f
C178 B.n144 VSUBS 0.009564f
C179 B.n145 VSUBS 0.009564f
C180 B.n146 VSUBS 0.009564f
C181 B.n147 VSUBS 0.009564f
C182 B.n148 VSUBS 0.009564f
C183 B.n149 VSUBS 0.009564f
C184 B.n150 VSUBS 0.009564f
C185 B.n151 VSUBS 0.009564f
C186 B.n152 VSUBS 0.009564f
C187 B.n153 VSUBS 0.009564f
C188 B.n154 VSUBS 0.009564f
C189 B.n155 VSUBS 0.009564f
C190 B.n156 VSUBS 0.009564f
C191 B.n157 VSUBS 0.00661f
C192 B.n158 VSUBS 0.009564f
C193 B.n159 VSUBS 0.009564f
C194 B.n160 VSUBS 0.009564f
C195 B.n161 VSUBS 0.009564f
C196 B.n162 VSUBS 0.009564f
C197 B.t7 VSUBS 0.152521f
C198 B.t8 VSUBS 0.20426f
C199 B.t6 VSUBS 1.80674f
C200 B.n163 VSUBS 0.333512f
C201 B.n164 VSUBS 0.251215f
C202 B.n165 VSUBS 0.009564f
C203 B.n166 VSUBS 0.009564f
C204 B.n167 VSUBS 0.009564f
C205 B.n168 VSUBS 0.009564f
C206 B.n169 VSUBS 0.009564f
C207 B.n170 VSUBS 0.009564f
C208 B.n171 VSUBS 0.009564f
C209 B.n172 VSUBS 0.009564f
C210 B.n173 VSUBS 0.009564f
C211 B.n174 VSUBS 0.009564f
C212 B.n175 VSUBS 0.009564f
C213 B.n176 VSUBS 0.009564f
C214 B.n177 VSUBS 0.009564f
C215 B.n178 VSUBS 0.022184f
C216 B.n179 VSUBS 0.009564f
C217 B.n180 VSUBS 0.009564f
C218 B.n181 VSUBS 0.009564f
C219 B.n182 VSUBS 0.009564f
C220 B.n183 VSUBS 0.009564f
C221 B.n184 VSUBS 0.009564f
C222 B.n185 VSUBS 0.009564f
C223 B.n186 VSUBS 0.009564f
C224 B.n187 VSUBS 0.009564f
C225 B.n188 VSUBS 0.009564f
C226 B.n189 VSUBS 0.009564f
C227 B.n190 VSUBS 0.009564f
C228 B.n191 VSUBS 0.009564f
C229 B.n192 VSUBS 0.009564f
C230 B.n193 VSUBS 0.009564f
C231 B.n194 VSUBS 0.009564f
C232 B.n195 VSUBS 0.009564f
C233 B.n196 VSUBS 0.009564f
C234 B.n197 VSUBS 0.009564f
C235 B.n198 VSUBS 0.009564f
C236 B.n199 VSUBS 0.009564f
C237 B.n200 VSUBS 0.009564f
C238 B.n201 VSUBS 0.009564f
C239 B.n202 VSUBS 0.009564f
C240 B.n203 VSUBS 0.009564f
C241 B.n204 VSUBS 0.009564f
C242 B.n205 VSUBS 0.009564f
C243 B.n206 VSUBS 0.009564f
C244 B.n207 VSUBS 0.009564f
C245 B.n208 VSUBS 0.009564f
C246 B.n209 VSUBS 0.009564f
C247 B.n210 VSUBS 0.009564f
C248 B.n211 VSUBS 0.009564f
C249 B.n212 VSUBS 0.009564f
C250 B.n213 VSUBS 0.009564f
C251 B.n214 VSUBS 0.009564f
C252 B.n215 VSUBS 0.009564f
C253 B.n216 VSUBS 0.009564f
C254 B.n217 VSUBS 0.009564f
C255 B.n218 VSUBS 0.009564f
C256 B.n219 VSUBS 0.009564f
C257 B.n220 VSUBS 0.009564f
C258 B.n221 VSUBS 0.009564f
C259 B.n222 VSUBS 0.009564f
C260 B.n223 VSUBS 0.009564f
C261 B.n224 VSUBS 0.009564f
C262 B.n225 VSUBS 0.009564f
C263 B.n226 VSUBS 0.009564f
C264 B.n227 VSUBS 0.009564f
C265 B.n228 VSUBS 0.009564f
C266 B.n229 VSUBS 0.009564f
C267 B.n230 VSUBS 0.009564f
C268 B.n231 VSUBS 0.009564f
C269 B.n232 VSUBS 0.009564f
C270 B.n233 VSUBS 0.009564f
C271 B.n234 VSUBS 0.009564f
C272 B.n235 VSUBS 0.009564f
C273 B.n236 VSUBS 0.009564f
C274 B.n237 VSUBS 0.009564f
C275 B.n238 VSUBS 0.009564f
C276 B.n239 VSUBS 0.009564f
C277 B.n240 VSUBS 0.009564f
C278 B.n241 VSUBS 0.009564f
C279 B.n242 VSUBS 0.009564f
C280 B.n243 VSUBS 0.009564f
C281 B.n244 VSUBS 0.009564f
C282 B.n245 VSUBS 0.009564f
C283 B.n246 VSUBS 0.009564f
C284 B.n247 VSUBS 0.009564f
C285 B.n248 VSUBS 0.009564f
C286 B.n249 VSUBS 0.009564f
C287 B.n250 VSUBS 0.009564f
C288 B.n251 VSUBS 0.009564f
C289 B.n252 VSUBS 0.009564f
C290 B.n253 VSUBS 0.009564f
C291 B.n254 VSUBS 0.009564f
C292 B.n255 VSUBS 0.009564f
C293 B.n256 VSUBS 0.009564f
C294 B.n257 VSUBS 0.009564f
C295 B.n258 VSUBS 0.009564f
C296 B.n259 VSUBS 0.009564f
C297 B.n260 VSUBS 0.009564f
C298 B.n261 VSUBS 0.009564f
C299 B.n262 VSUBS 0.009564f
C300 B.n263 VSUBS 0.009564f
C301 B.n264 VSUBS 0.009564f
C302 B.n265 VSUBS 0.009564f
C303 B.n266 VSUBS 0.009564f
C304 B.n267 VSUBS 0.009564f
C305 B.n268 VSUBS 0.009564f
C306 B.n269 VSUBS 0.009564f
C307 B.n270 VSUBS 0.009564f
C308 B.n271 VSUBS 0.009564f
C309 B.n272 VSUBS 0.009564f
C310 B.n273 VSUBS 0.009564f
C311 B.n274 VSUBS 0.009564f
C312 B.n275 VSUBS 0.009564f
C313 B.n276 VSUBS 0.009564f
C314 B.n277 VSUBS 0.009564f
C315 B.n278 VSUBS 0.009564f
C316 B.n279 VSUBS 0.009564f
C317 B.n280 VSUBS 0.009564f
C318 B.n281 VSUBS 0.009564f
C319 B.n282 VSUBS 0.009564f
C320 B.n283 VSUBS 0.009564f
C321 B.n284 VSUBS 0.009564f
C322 B.n285 VSUBS 0.009564f
C323 B.n286 VSUBS 0.009564f
C324 B.n287 VSUBS 0.009564f
C325 B.n288 VSUBS 0.009564f
C326 B.n289 VSUBS 0.009564f
C327 B.n290 VSUBS 0.009564f
C328 B.n291 VSUBS 0.009564f
C329 B.n292 VSUBS 0.009564f
C330 B.n293 VSUBS 0.009564f
C331 B.n294 VSUBS 0.009564f
C332 B.n295 VSUBS 0.009564f
C333 B.n296 VSUBS 0.009564f
C334 B.n297 VSUBS 0.009564f
C335 B.n298 VSUBS 0.009564f
C336 B.n299 VSUBS 0.009564f
C337 B.n300 VSUBS 0.009564f
C338 B.n301 VSUBS 0.009564f
C339 B.n302 VSUBS 0.009564f
C340 B.n303 VSUBS 0.009564f
C341 B.n304 VSUBS 0.009564f
C342 B.n305 VSUBS 0.009564f
C343 B.n306 VSUBS 0.009564f
C344 B.n307 VSUBS 0.009564f
C345 B.n308 VSUBS 0.009564f
C346 B.n309 VSUBS 0.009564f
C347 B.n310 VSUBS 0.009564f
C348 B.n311 VSUBS 0.009564f
C349 B.n312 VSUBS 0.009564f
C350 B.n313 VSUBS 0.022184f
C351 B.n314 VSUBS 0.023948f
C352 B.n315 VSUBS 0.023948f
C353 B.n316 VSUBS 0.009564f
C354 B.n317 VSUBS 0.009564f
C355 B.n318 VSUBS 0.009564f
C356 B.n319 VSUBS 0.009564f
C357 B.n320 VSUBS 0.009564f
C358 B.n321 VSUBS 0.009564f
C359 B.n322 VSUBS 0.009564f
C360 B.n323 VSUBS 0.009564f
C361 B.n324 VSUBS 0.009564f
C362 B.n325 VSUBS 0.009564f
C363 B.n326 VSUBS 0.009564f
C364 B.n327 VSUBS 0.009564f
C365 B.n328 VSUBS 0.009564f
C366 B.n329 VSUBS 0.009564f
C367 B.n330 VSUBS 0.009564f
C368 B.n331 VSUBS 0.009564f
C369 B.n332 VSUBS 0.009564f
C370 B.n333 VSUBS 0.009564f
C371 B.n334 VSUBS 0.009564f
C372 B.n335 VSUBS 0.009564f
C373 B.n336 VSUBS 0.009564f
C374 B.n337 VSUBS 0.009564f
C375 B.n338 VSUBS 0.009564f
C376 B.n339 VSUBS 0.009564f
C377 B.n340 VSUBS 0.009564f
C378 B.n341 VSUBS 0.009564f
C379 B.n342 VSUBS 0.009564f
C380 B.n343 VSUBS 0.009564f
C381 B.n344 VSUBS 0.009564f
C382 B.n345 VSUBS 0.009564f
C383 B.n346 VSUBS 0.009564f
C384 B.n347 VSUBS 0.009564f
C385 B.n348 VSUBS 0.009564f
C386 B.n349 VSUBS 0.009564f
C387 B.n350 VSUBS 0.009564f
C388 B.n351 VSUBS 0.009564f
C389 B.n352 VSUBS 0.009564f
C390 B.n353 VSUBS 0.009564f
C391 B.n354 VSUBS 0.009564f
C392 B.n355 VSUBS 0.00661f
C393 B.n356 VSUBS 0.022159f
C394 B.n357 VSUBS 0.007736f
C395 B.n358 VSUBS 0.009564f
C396 B.n359 VSUBS 0.009564f
C397 B.n360 VSUBS 0.009564f
C398 B.n361 VSUBS 0.009564f
C399 B.n362 VSUBS 0.009564f
C400 B.n363 VSUBS 0.009564f
C401 B.n364 VSUBS 0.009564f
C402 B.n365 VSUBS 0.009564f
C403 B.n366 VSUBS 0.009564f
C404 B.n367 VSUBS 0.009564f
C405 B.n368 VSUBS 0.009564f
C406 B.t10 VSUBS 0.152524f
C407 B.t11 VSUBS 0.204263f
C408 B.t9 VSUBS 1.80674f
C409 B.n369 VSUBS 0.33351f
C410 B.n370 VSUBS 0.251212f
C411 B.n371 VSUBS 0.022159f
C412 B.n372 VSUBS 0.007736f
C413 B.n373 VSUBS 0.009564f
C414 B.n374 VSUBS 0.009564f
C415 B.n375 VSUBS 0.009564f
C416 B.n376 VSUBS 0.009564f
C417 B.n377 VSUBS 0.009564f
C418 B.n378 VSUBS 0.009564f
C419 B.n379 VSUBS 0.009564f
C420 B.n380 VSUBS 0.009564f
C421 B.n381 VSUBS 0.009564f
C422 B.n382 VSUBS 0.009564f
C423 B.n383 VSUBS 0.009564f
C424 B.n384 VSUBS 0.009564f
C425 B.n385 VSUBS 0.009564f
C426 B.n386 VSUBS 0.009564f
C427 B.n387 VSUBS 0.009564f
C428 B.n388 VSUBS 0.009564f
C429 B.n389 VSUBS 0.009564f
C430 B.n390 VSUBS 0.009564f
C431 B.n391 VSUBS 0.009564f
C432 B.n392 VSUBS 0.009564f
C433 B.n393 VSUBS 0.009564f
C434 B.n394 VSUBS 0.009564f
C435 B.n395 VSUBS 0.009564f
C436 B.n396 VSUBS 0.009564f
C437 B.n397 VSUBS 0.009564f
C438 B.n398 VSUBS 0.009564f
C439 B.n399 VSUBS 0.009564f
C440 B.n400 VSUBS 0.009564f
C441 B.n401 VSUBS 0.009564f
C442 B.n402 VSUBS 0.009564f
C443 B.n403 VSUBS 0.009564f
C444 B.n404 VSUBS 0.009564f
C445 B.n405 VSUBS 0.009564f
C446 B.n406 VSUBS 0.009564f
C447 B.n407 VSUBS 0.009564f
C448 B.n408 VSUBS 0.009564f
C449 B.n409 VSUBS 0.009564f
C450 B.n410 VSUBS 0.009564f
C451 B.n411 VSUBS 0.009564f
C452 B.n412 VSUBS 0.009564f
C453 B.n413 VSUBS 0.009564f
C454 B.n414 VSUBS 0.023948f
C455 B.n415 VSUBS 0.023948f
C456 B.n416 VSUBS 0.022184f
C457 B.n417 VSUBS 0.009564f
C458 B.n418 VSUBS 0.009564f
C459 B.n419 VSUBS 0.009564f
C460 B.n420 VSUBS 0.009564f
C461 B.n421 VSUBS 0.009564f
C462 B.n422 VSUBS 0.009564f
C463 B.n423 VSUBS 0.009564f
C464 B.n424 VSUBS 0.009564f
C465 B.n425 VSUBS 0.009564f
C466 B.n426 VSUBS 0.009564f
C467 B.n427 VSUBS 0.009564f
C468 B.n428 VSUBS 0.009564f
C469 B.n429 VSUBS 0.009564f
C470 B.n430 VSUBS 0.009564f
C471 B.n431 VSUBS 0.009564f
C472 B.n432 VSUBS 0.009564f
C473 B.n433 VSUBS 0.009564f
C474 B.n434 VSUBS 0.009564f
C475 B.n435 VSUBS 0.009564f
C476 B.n436 VSUBS 0.009564f
C477 B.n437 VSUBS 0.009564f
C478 B.n438 VSUBS 0.009564f
C479 B.n439 VSUBS 0.009564f
C480 B.n440 VSUBS 0.009564f
C481 B.n441 VSUBS 0.009564f
C482 B.n442 VSUBS 0.009564f
C483 B.n443 VSUBS 0.009564f
C484 B.n444 VSUBS 0.009564f
C485 B.n445 VSUBS 0.009564f
C486 B.n446 VSUBS 0.009564f
C487 B.n447 VSUBS 0.009564f
C488 B.n448 VSUBS 0.009564f
C489 B.n449 VSUBS 0.009564f
C490 B.n450 VSUBS 0.009564f
C491 B.n451 VSUBS 0.009564f
C492 B.n452 VSUBS 0.009564f
C493 B.n453 VSUBS 0.009564f
C494 B.n454 VSUBS 0.009564f
C495 B.n455 VSUBS 0.009564f
C496 B.n456 VSUBS 0.009564f
C497 B.n457 VSUBS 0.009564f
C498 B.n458 VSUBS 0.009564f
C499 B.n459 VSUBS 0.009564f
C500 B.n460 VSUBS 0.009564f
C501 B.n461 VSUBS 0.009564f
C502 B.n462 VSUBS 0.009564f
C503 B.n463 VSUBS 0.009564f
C504 B.n464 VSUBS 0.009564f
C505 B.n465 VSUBS 0.009564f
C506 B.n466 VSUBS 0.009564f
C507 B.n467 VSUBS 0.009564f
C508 B.n468 VSUBS 0.009564f
C509 B.n469 VSUBS 0.009564f
C510 B.n470 VSUBS 0.009564f
C511 B.n471 VSUBS 0.009564f
C512 B.n472 VSUBS 0.009564f
C513 B.n473 VSUBS 0.009564f
C514 B.n474 VSUBS 0.009564f
C515 B.n475 VSUBS 0.009564f
C516 B.n476 VSUBS 0.009564f
C517 B.n477 VSUBS 0.009564f
C518 B.n478 VSUBS 0.009564f
C519 B.n479 VSUBS 0.009564f
C520 B.n480 VSUBS 0.009564f
C521 B.n481 VSUBS 0.009564f
C522 B.n482 VSUBS 0.009564f
C523 B.n483 VSUBS 0.009564f
C524 B.n484 VSUBS 0.009564f
C525 B.n485 VSUBS 0.009564f
C526 B.n486 VSUBS 0.009564f
C527 B.n487 VSUBS 0.009564f
C528 B.n488 VSUBS 0.009564f
C529 B.n489 VSUBS 0.009564f
C530 B.n490 VSUBS 0.009564f
C531 B.n491 VSUBS 0.009564f
C532 B.n492 VSUBS 0.009564f
C533 B.n493 VSUBS 0.009564f
C534 B.n494 VSUBS 0.009564f
C535 B.n495 VSUBS 0.009564f
C536 B.n496 VSUBS 0.009564f
C537 B.n497 VSUBS 0.009564f
C538 B.n498 VSUBS 0.009564f
C539 B.n499 VSUBS 0.009564f
C540 B.n500 VSUBS 0.009564f
C541 B.n501 VSUBS 0.009564f
C542 B.n502 VSUBS 0.009564f
C543 B.n503 VSUBS 0.009564f
C544 B.n504 VSUBS 0.009564f
C545 B.n505 VSUBS 0.009564f
C546 B.n506 VSUBS 0.009564f
C547 B.n507 VSUBS 0.009564f
C548 B.n508 VSUBS 0.009564f
C549 B.n509 VSUBS 0.009564f
C550 B.n510 VSUBS 0.009564f
C551 B.n511 VSUBS 0.009564f
C552 B.n512 VSUBS 0.009564f
C553 B.n513 VSUBS 0.009564f
C554 B.n514 VSUBS 0.009564f
C555 B.n515 VSUBS 0.009564f
C556 B.n516 VSUBS 0.009564f
C557 B.n517 VSUBS 0.009564f
C558 B.n518 VSUBS 0.009564f
C559 B.n519 VSUBS 0.009564f
C560 B.n520 VSUBS 0.009564f
C561 B.n521 VSUBS 0.009564f
C562 B.n522 VSUBS 0.009564f
C563 B.n523 VSUBS 0.009564f
C564 B.n524 VSUBS 0.009564f
C565 B.n525 VSUBS 0.009564f
C566 B.n526 VSUBS 0.009564f
C567 B.n527 VSUBS 0.009564f
C568 B.n528 VSUBS 0.009564f
C569 B.n529 VSUBS 0.009564f
C570 B.n530 VSUBS 0.009564f
C571 B.n531 VSUBS 0.009564f
C572 B.n532 VSUBS 0.009564f
C573 B.n533 VSUBS 0.009564f
C574 B.n534 VSUBS 0.009564f
C575 B.n535 VSUBS 0.009564f
C576 B.n536 VSUBS 0.009564f
C577 B.n537 VSUBS 0.009564f
C578 B.n538 VSUBS 0.009564f
C579 B.n539 VSUBS 0.009564f
C580 B.n540 VSUBS 0.009564f
C581 B.n541 VSUBS 0.009564f
C582 B.n542 VSUBS 0.009564f
C583 B.n543 VSUBS 0.009564f
C584 B.n544 VSUBS 0.009564f
C585 B.n545 VSUBS 0.009564f
C586 B.n546 VSUBS 0.009564f
C587 B.n547 VSUBS 0.009564f
C588 B.n548 VSUBS 0.009564f
C589 B.n549 VSUBS 0.009564f
C590 B.n550 VSUBS 0.009564f
C591 B.n551 VSUBS 0.009564f
C592 B.n552 VSUBS 0.009564f
C593 B.n553 VSUBS 0.009564f
C594 B.n554 VSUBS 0.009564f
C595 B.n555 VSUBS 0.009564f
C596 B.n556 VSUBS 0.009564f
C597 B.n557 VSUBS 0.009564f
C598 B.n558 VSUBS 0.009564f
C599 B.n559 VSUBS 0.009564f
C600 B.n560 VSUBS 0.009564f
C601 B.n561 VSUBS 0.009564f
C602 B.n562 VSUBS 0.009564f
C603 B.n563 VSUBS 0.009564f
C604 B.n564 VSUBS 0.009564f
C605 B.n565 VSUBS 0.009564f
C606 B.n566 VSUBS 0.009564f
C607 B.n567 VSUBS 0.009564f
C608 B.n568 VSUBS 0.009564f
C609 B.n569 VSUBS 0.009564f
C610 B.n570 VSUBS 0.009564f
C611 B.n571 VSUBS 0.009564f
C612 B.n572 VSUBS 0.009564f
C613 B.n573 VSUBS 0.009564f
C614 B.n574 VSUBS 0.009564f
C615 B.n575 VSUBS 0.009564f
C616 B.n576 VSUBS 0.009564f
C617 B.n577 VSUBS 0.009564f
C618 B.n578 VSUBS 0.009564f
C619 B.n579 VSUBS 0.009564f
C620 B.n580 VSUBS 0.009564f
C621 B.n581 VSUBS 0.009564f
C622 B.n582 VSUBS 0.009564f
C623 B.n583 VSUBS 0.009564f
C624 B.n584 VSUBS 0.009564f
C625 B.n585 VSUBS 0.009564f
C626 B.n586 VSUBS 0.009564f
C627 B.n587 VSUBS 0.009564f
C628 B.n588 VSUBS 0.009564f
C629 B.n589 VSUBS 0.009564f
C630 B.n590 VSUBS 0.009564f
C631 B.n591 VSUBS 0.009564f
C632 B.n592 VSUBS 0.009564f
C633 B.n593 VSUBS 0.009564f
C634 B.n594 VSUBS 0.009564f
C635 B.n595 VSUBS 0.009564f
C636 B.n596 VSUBS 0.009564f
C637 B.n597 VSUBS 0.009564f
C638 B.n598 VSUBS 0.009564f
C639 B.n599 VSUBS 0.009564f
C640 B.n600 VSUBS 0.009564f
C641 B.n601 VSUBS 0.009564f
C642 B.n602 VSUBS 0.009564f
C643 B.n603 VSUBS 0.009564f
C644 B.n604 VSUBS 0.009564f
C645 B.n605 VSUBS 0.009564f
C646 B.n606 VSUBS 0.009564f
C647 B.n607 VSUBS 0.009564f
C648 B.n608 VSUBS 0.009564f
C649 B.n609 VSUBS 0.009564f
C650 B.n610 VSUBS 0.009564f
C651 B.n611 VSUBS 0.009564f
C652 B.n612 VSUBS 0.009564f
C653 B.n613 VSUBS 0.009564f
C654 B.n614 VSUBS 0.009564f
C655 B.n615 VSUBS 0.009564f
C656 B.n616 VSUBS 0.009564f
C657 B.n617 VSUBS 0.009564f
C658 B.n618 VSUBS 0.009564f
C659 B.n619 VSUBS 0.009564f
C660 B.n620 VSUBS 0.009564f
C661 B.n621 VSUBS 0.009564f
C662 B.n622 VSUBS 0.009564f
C663 B.n623 VSUBS 0.023264f
C664 B.n624 VSUBS 0.022869f
C665 B.n625 VSUBS 0.023948f
C666 B.n626 VSUBS 0.009564f
C667 B.n627 VSUBS 0.009564f
C668 B.n628 VSUBS 0.009564f
C669 B.n629 VSUBS 0.009564f
C670 B.n630 VSUBS 0.009564f
C671 B.n631 VSUBS 0.009564f
C672 B.n632 VSUBS 0.009564f
C673 B.n633 VSUBS 0.009564f
C674 B.n634 VSUBS 0.009564f
C675 B.n635 VSUBS 0.009564f
C676 B.n636 VSUBS 0.009564f
C677 B.n637 VSUBS 0.009564f
C678 B.n638 VSUBS 0.009564f
C679 B.n639 VSUBS 0.009564f
C680 B.n640 VSUBS 0.009564f
C681 B.n641 VSUBS 0.009564f
C682 B.n642 VSUBS 0.009564f
C683 B.n643 VSUBS 0.009564f
C684 B.n644 VSUBS 0.009564f
C685 B.n645 VSUBS 0.009564f
C686 B.n646 VSUBS 0.009564f
C687 B.n647 VSUBS 0.009564f
C688 B.n648 VSUBS 0.009564f
C689 B.n649 VSUBS 0.009564f
C690 B.n650 VSUBS 0.009564f
C691 B.n651 VSUBS 0.009564f
C692 B.n652 VSUBS 0.009564f
C693 B.n653 VSUBS 0.009564f
C694 B.n654 VSUBS 0.009564f
C695 B.n655 VSUBS 0.009564f
C696 B.n656 VSUBS 0.009564f
C697 B.n657 VSUBS 0.009564f
C698 B.n658 VSUBS 0.009564f
C699 B.n659 VSUBS 0.009564f
C700 B.n660 VSUBS 0.009564f
C701 B.n661 VSUBS 0.009564f
C702 B.n662 VSUBS 0.009564f
C703 B.n663 VSUBS 0.009564f
C704 B.n664 VSUBS 0.009564f
C705 B.n665 VSUBS 0.00661f
C706 B.n666 VSUBS 0.022159f
C707 B.n667 VSUBS 0.007736f
C708 B.n668 VSUBS 0.009564f
C709 B.n669 VSUBS 0.009564f
C710 B.n670 VSUBS 0.009564f
C711 B.n671 VSUBS 0.009564f
C712 B.n672 VSUBS 0.009564f
C713 B.n673 VSUBS 0.009564f
C714 B.n674 VSUBS 0.009564f
C715 B.n675 VSUBS 0.009564f
C716 B.n676 VSUBS 0.009564f
C717 B.n677 VSUBS 0.009564f
C718 B.n678 VSUBS 0.009564f
C719 B.n679 VSUBS 0.007736f
C720 B.n680 VSUBS 0.009564f
C721 B.n681 VSUBS 0.009564f
C722 B.n682 VSUBS 0.009564f
C723 B.n683 VSUBS 0.009564f
C724 B.n684 VSUBS 0.009564f
C725 B.n685 VSUBS 0.009564f
C726 B.n686 VSUBS 0.009564f
C727 B.n687 VSUBS 0.009564f
C728 B.n688 VSUBS 0.009564f
C729 B.n689 VSUBS 0.009564f
C730 B.n690 VSUBS 0.009564f
C731 B.n691 VSUBS 0.009564f
C732 B.n692 VSUBS 0.009564f
C733 B.n693 VSUBS 0.009564f
C734 B.n694 VSUBS 0.009564f
C735 B.n695 VSUBS 0.009564f
C736 B.n696 VSUBS 0.009564f
C737 B.n697 VSUBS 0.009564f
C738 B.n698 VSUBS 0.009564f
C739 B.n699 VSUBS 0.009564f
C740 B.n700 VSUBS 0.009564f
C741 B.n701 VSUBS 0.009564f
C742 B.n702 VSUBS 0.009564f
C743 B.n703 VSUBS 0.009564f
C744 B.n704 VSUBS 0.009564f
C745 B.n705 VSUBS 0.009564f
C746 B.n706 VSUBS 0.009564f
C747 B.n707 VSUBS 0.009564f
C748 B.n708 VSUBS 0.009564f
C749 B.n709 VSUBS 0.009564f
C750 B.n710 VSUBS 0.009564f
C751 B.n711 VSUBS 0.009564f
C752 B.n712 VSUBS 0.009564f
C753 B.n713 VSUBS 0.009564f
C754 B.n714 VSUBS 0.009564f
C755 B.n715 VSUBS 0.009564f
C756 B.n716 VSUBS 0.009564f
C757 B.n717 VSUBS 0.009564f
C758 B.n718 VSUBS 0.009564f
C759 B.n719 VSUBS 0.009564f
C760 B.n720 VSUBS 0.009564f
C761 B.n721 VSUBS 0.023948f
C762 B.n722 VSUBS 0.023948f
C763 B.n723 VSUBS 0.022184f
C764 B.n724 VSUBS 0.009564f
C765 B.n725 VSUBS 0.009564f
C766 B.n726 VSUBS 0.009564f
C767 B.n727 VSUBS 0.009564f
C768 B.n728 VSUBS 0.009564f
C769 B.n729 VSUBS 0.009564f
C770 B.n730 VSUBS 0.009564f
C771 B.n731 VSUBS 0.009564f
C772 B.n732 VSUBS 0.009564f
C773 B.n733 VSUBS 0.009564f
C774 B.n734 VSUBS 0.009564f
C775 B.n735 VSUBS 0.009564f
C776 B.n736 VSUBS 0.009564f
C777 B.n737 VSUBS 0.009564f
C778 B.n738 VSUBS 0.009564f
C779 B.n739 VSUBS 0.009564f
C780 B.n740 VSUBS 0.009564f
C781 B.n741 VSUBS 0.009564f
C782 B.n742 VSUBS 0.009564f
C783 B.n743 VSUBS 0.009564f
C784 B.n744 VSUBS 0.009564f
C785 B.n745 VSUBS 0.009564f
C786 B.n746 VSUBS 0.009564f
C787 B.n747 VSUBS 0.009564f
C788 B.n748 VSUBS 0.009564f
C789 B.n749 VSUBS 0.009564f
C790 B.n750 VSUBS 0.009564f
C791 B.n751 VSUBS 0.009564f
C792 B.n752 VSUBS 0.009564f
C793 B.n753 VSUBS 0.009564f
C794 B.n754 VSUBS 0.009564f
C795 B.n755 VSUBS 0.009564f
C796 B.n756 VSUBS 0.009564f
C797 B.n757 VSUBS 0.009564f
C798 B.n758 VSUBS 0.009564f
C799 B.n759 VSUBS 0.009564f
C800 B.n760 VSUBS 0.009564f
C801 B.n761 VSUBS 0.009564f
C802 B.n762 VSUBS 0.009564f
C803 B.n763 VSUBS 0.009564f
C804 B.n764 VSUBS 0.009564f
C805 B.n765 VSUBS 0.009564f
C806 B.n766 VSUBS 0.009564f
C807 B.n767 VSUBS 0.009564f
C808 B.n768 VSUBS 0.009564f
C809 B.n769 VSUBS 0.009564f
C810 B.n770 VSUBS 0.009564f
C811 B.n771 VSUBS 0.009564f
C812 B.n772 VSUBS 0.009564f
C813 B.n773 VSUBS 0.009564f
C814 B.n774 VSUBS 0.009564f
C815 B.n775 VSUBS 0.009564f
C816 B.n776 VSUBS 0.009564f
C817 B.n777 VSUBS 0.009564f
C818 B.n778 VSUBS 0.009564f
C819 B.n779 VSUBS 0.009564f
C820 B.n780 VSUBS 0.009564f
C821 B.n781 VSUBS 0.009564f
C822 B.n782 VSUBS 0.009564f
C823 B.n783 VSUBS 0.009564f
C824 B.n784 VSUBS 0.009564f
C825 B.n785 VSUBS 0.009564f
C826 B.n786 VSUBS 0.009564f
C827 B.n787 VSUBS 0.009564f
C828 B.n788 VSUBS 0.009564f
C829 B.n789 VSUBS 0.009564f
C830 B.n790 VSUBS 0.009564f
C831 B.n791 VSUBS 0.009564f
C832 B.n792 VSUBS 0.009564f
C833 B.n793 VSUBS 0.009564f
C834 B.n794 VSUBS 0.009564f
C835 B.n795 VSUBS 0.009564f
C836 B.n796 VSUBS 0.009564f
C837 B.n797 VSUBS 0.009564f
C838 B.n798 VSUBS 0.009564f
C839 B.n799 VSUBS 0.009564f
C840 B.n800 VSUBS 0.009564f
C841 B.n801 VSUBS 0.009564f
C842 B.n802 VSUBS 0.009564f
C843 B.n803 VSUBS 0.009564f
C844 B.n804 VSUBS 0.009564f
C845 B.n805 VSUBS 0.009564f
C846 B.n806 VSUBS 0.009564f
C847 B.n807 VSUBS 0.009564f
C848 B.n808 VSUBS 0.009564f
C849 B.n809 VSUBS 0.009564f
C850 B.n810 VSUBS 0.009564f
C851 B.n811 VSUBS 0.009564f
C852 B.n812 VSUBS 0.009564f
C853 B.n813 VSUBS 0.009564f
C854 B.n814 VSUBS 0.009564f
C855 B.n815 VSUBS 0.009564f
C856 B.n816 VSUBS 0.009564f
C857 B.n817 VSUBS 0.009564f
C858 B.n818 VSUBS 0.009564f
C859 B.n819 VSUBS 0.009564f
C860 B.n820 VSUBS 0.009564f
C861 B.n821 VSUBS 0.009564f
C862 B.n822 VSUBS 0.009564f
C863 B.n823 VSUBS 0.009564f
C864 B.n824 VSUBS 0.009564f
C865 B.n825 VSUBS 0.009564f
C866 B.n826 VSUBS 0.009564f
C867 B.n827 VSUBS 0.021657f
C868 VDD2.t4 VSUBS 0.208793f
C869 VDD2.t5 VSUBS 0.208793f
C870 VDD2.n0 VSUBS 1.50393f
C871 VDD2.t1 VSUBS 0.208793f
C872 VDD2.t0 VSUBS 0.208793f
C873 VDD2.n1 VSUBS 1.50393f
C874 VDD2.n2 VSUBS 5.99479f
C875 VDD2.t7 VSUBS 0.208793f
C876 VDD2.t6 VSUBS 0.208793f
C877 VDD2.n3 VSUBS 1.47981f
C878 VDD2.n4 VSUBS 4.70391f
C879 VDD2.t2 VSUBS 0.208793f
C880 VDD2.t3 VSUBS 0.208793f
C881 VDD2.n5 VSUBS 1.50387f
C882 VN.n0 VSUBS 0.054154f
C883 VN.t7 VSUBS 2.13118f
C884 VN.n1 VSUBS 0.05791f
C885 VN.n2 VSUBS 0.02879f
C886 VN.n3 VSUBS 0.053657f
C887 VN.n4 VSUBS 0.02879f
C888 VN.t6 VSUBS 2.13118f
C889 VN.n5 VSUBS 0.053657f
C890 VN.n6 VSUBS 0.02879f
C891 VN.n7 VSUBS 0.053657f
C892 VN.t3 VSUBS 2.54481f
C893 VN.n8 VSUBS 0.848786f
C894 VN.t2 VSUBS 2.13118f
C895 VN.n9 VSUBS 0.879276f
C896 VN.n10 VSUBS 0.04465f
C897 VN.n11 VSUBS 0.373587f
C898 VN.n12 VSUBS 0.02879f
C899 VN.n13 VSUBS 0.02879f
C900 VN.n14 VSUBS 0.053657f
C901 VN.n15 VSUBS 0.042028f
C902 VN.n16 VSUBS 0.042028f
C903 VN.n17 VSUBS 0.02879f
C904 VN.n18 VSUBS 0.02879f
C905 VN.n19 VSUBS 0.02879f
C906 VN.n20 VSUBS 0.053657f
C907 VN.n21 VSUBS 0.04465f
C908 VN.n22 VSUBS 0.771218f
C909 VN.n23 VSUBS 0.036173f
C910 VN.n24 VSUBS 0.02879f
C911 VN.n25 VSUBS 0.02879f
C912 VN.n26 VSUBS 0.02879f
C913 VN.n27 VSUBS 0.053657f
C914 VN.n28 VSUBS 0.053388f
C915 VN.n29 VSUBS 0.026415f
C916 VN.n30 VSUBS 0.02879f
C917 VN.n31 VSUBS 0.02879f
C918 VN.n32 VSUBS 0.02879f
C919 VN.n33 VSUBS 0.053657f
C920 VN.n34 VSUBS 0.053127f
C921 VN.n35 VSUBS 0.901865f
C922 VN.n36 VSUBS 0.083738f
C923 VN.n37 VSUBS 0.054154f
C924 VN.t0 VSUBS 2.13118f
C925 VN.n38 VSUBS 0.05791f
C926 VN.n39 VSUBS 0.02879f
C927 VN.n40 VSUBS 0.053657f
C928 VN.n41 VSUBS 0.02879f
C929 VN.t1 VSUBS 2.13118f
C930 VN.n42 VSUBS 0.053657f
C931 VN.n43 VSUBS 0.02879f
C932 VN.n44 VSUBS 0.053657f
C933 VN.t4 VSUBS 2.54481f
C934 VN.n45 VSUBS 0.848786f
C935 VN.t5 VSUBS 2.13118f
C936 VN.n46 VSUBS 0.879276f
C937 VN.n47 VSUBS 0.04465f
C938 VN.n48 VSUBS 0.373587f
C939 VN.n49 VSUBS 0.02879f
C940 VN.n50 VSUBS 0.02879f
C941 VN.n51 VSUBS 0.053657f
C942 VN.n52 VSUBS 0.042028f
C943 VN.n53 VSUBS 0.042028f
C944 VN.n54 VSUBS 0.02879f
C945 VN.n55 VSUBS 0.02879f
C946 VN.n56 VSUBS 0.02879f
C947 VN.n57 VSUBS 0.053657f
C948 VN.n58 VSUBS 0.04465f
C949 VN.n59 VSUBS 0.771218f
C950 VN.n60 VSUBS 0.036173f
C951 VN.n61 VSUBS 0.02879f
C952 VN.n62 VSUBS 0.02879f
C953 VN.n63 VSUBS 0.02879f
C954 VN.n64 VSUBS 0.053657f
C955 VN.n65 VSUBS 0.053388f
C956 VN.n66 VSUBS 0.026415f
C957 VN.n67 VSUBS 0.02879f
C958 VN.n68 VSUBS 0.02879f
C959 VN.n69 VSUBS 0.02879f
C960 VN.n70 VSUBS 0.053657f
C961 VN.n71 VSUBS 0.053127f
C962 VN.n72 VSUBS 0.901865f
C963 VN.n73 VSUBS 1.83098f
C964 VTAIL.t1 VSUBS 0.16732f
C965 VTAIL.t7 VSUBS 0.16732f
C966 VTAIL.n0 VSUBS 1.07435f
C967 VTAIL.n1 VSUBS 0.896336f
C968 VTAIL.n2 VSUBS 0.03152f
C969 VTAIL.n3 VSUBS 0.029286f
C970 VTAIL.n4 VSUBS 0.015737f
C971 VTAIL.n5 VSUBS 0.037196f
C972 VTAIL.n6 VSUBS 0.016662f
C973 VTAIL.n7 VSUBS 0.029286f
C974 VTAIL.n8 VSUBS 0.015737f
C975 VTAIL.n9 VSUBS 0.037196f
C976 VTAIL.n10 VSUBS 0.016662f
C977 VTAIL.n11 VSUBS 0.826415f
C978 VTAIL.n12 VSUBS 0.015737f
C979 VTAIL.t4 VSUBS 0.079902f
C980 VTAIL.n13 VSUBS 0.16766f
C981 VTAIL.n14 VSUBS 0.02798f
C982 VTAIL.n15 VSUBS 0.027897f
C983 VTAIL.n16 VSUBS 0.037196f
C984 VTAIL.n17 VSUBS 0.016662f
C985 VTAIL.n18 VSUBS 0.015737f
C986 VTAIL.n19 VSUBS 0.029286f
C987 VTAIL.n20 VSUBS 0.029286f
C988 VTAIL.n21 VSUBS 0.015737f
C989 VTAIL.n22 VSUBS 0.016662f
C990 VTAIL.n23 VSUBS 0.037196f
C991 VTAIL.n24 VSUBS 0.037196f
C992 VTAIL.n25 VSUBS 0.016662f
C993 VTAIL.n26 VSUBS 0.015737f
C994 VTAIL.n27 VSUBS 0.029286f
C995 VTAIL.n28 VSUBS 0.029286f
C996 VTAIL.n29 VSUBS 0.015737f
C997 VTAIL.n30 VSUBS 0.016662f
C998 VTAIL.n31 VSUBS 0.037196f
C999 VTAIL.n32 VSUBS 0.092342f
C1000 VTAIL.n33 VSUBS 0.016662f
C1001 VTAIL.n34 VSUBS 0.030903f
C1002 VTAIL.n35 VSUBS 0.073693f
C1003 VTAIL.n36 VSUBS 0.070705f
C1004 VTAIL.n37 VSUBS 0.411153f
C1005 VTAIL.n38 VSUBS 0.03152f
C1006 VTAIL.n39 VSUBS 0.029286f
C1007 VTAIL.n40 VSUBS 0.015737f
C1008 VTAIL.n41 VSUBS 0.037196f
C1009 VTAIL.n42 VSUBS 0.016662f
C1010 VTAIL.n43 VSUBS 0.029286f
C1011 VTAIL.n44 VSUBS 0.015737f
C1012 VTAIL.n45 VSUBS 0.037196f
C1013 VTAIL.n46 VSUBS 0.016662f
C1014 VTAIL.n47 VSUBS 0.826415f
C1015 VTAIL.n48 VSUBS 0.015737f
C1016 VTAIL.t9 VSUBS 0.079902f
C1017 VTAIL.n49 VSUBS 0.16766f
C1018 VTAIL.n50 VSUBS 0.02798f
C1019 VTAIL.n51 VSUBS 0.027897f
C1020 VTAIL.n52 VSUBS 0.037196f
C1021 VTAIL.n53 VSUBS 0.016662f
C1022 VTAIL.n54 VSUBS 0.015737f
C1023 VTAIL.n55 VSUBS 0.029286f
C1024 VTAIL.n56 VSUBS 0.029286f
C1025 VTAIL.n57 VSUBS 0.015737f
C1026 VTAIL.n58 VSUBS 0.016662f
C1027 VTAIL.n59 VSUBS 0.037196f
C1028 VTAIL.n60 VSUBS 0.037196f
C1029 VTAIL.n61 VSUBS 0.016662f
C1030 VTAIL.n62 VSUBS 0.015737f
C1031 VTAIL.n63 VSUBS 0.029286f
C1032 VTAIL.n64 VSUBS 0.029286f
C1033 VTAIL.n65 VSUBS 0.015737f
C1034 VTAIL.n66 VSUBS 0.016662f
C1035 VTAIL.n67 VSUBS 0.037196f
C1036 VTAIL.n68 VSUBS 0.092342f
C1037 VTAIL.n69 VSUBS 0.016662f
C1038 VTAIL.n70 VSUBS 0.030903f
C1039 VTAIL.n71 VSUBS 0.073693f
C1040 VTAIL.n72 VSUBS 0.070705f
C1041 VTAIL.n73 VSUBS 0.411153f
C1042 VTAIL.t8 VSUBS 0.16732f
C1043 VTAIL.t10 VSUBS 0.16732f
C1044 VTAIL.n74 VSUBS 1.07435f
C1045 VTAIL.n75 VSUBS 1.22926f
C1046 VTAIL.n76 VSUBS 0.03152f
C1047 VTAIL.n77 VSUBS 0.029286f
C1048 VTAIL.n78 VSUBS 0.015737f
C1049 VTAIL.n79 VSUBS 0.037196f
C1050 VTAIL.n80 VSUBS 0.016662f
C1051 VTAIL.n81 VSUBS 0.029286f
C1052 VTAIL.n82 VSUBS 0.015737f
C1053 VTAIL.n83 VSUBS 0.037196f
C1054 VTAIL.n84 VSUBS 0.016662f
C1055 VTAIL.n85 VSUBS 0.826415f
C1056 VTAIL.n86 VSUBS 0.015737f
C1057 VTAIL.t11 VSUBS 0.079902f
C1058 VTAIL.n87 VSUBS 0.16766f
C1059 VTAIL.n88 VSUBS 0.02798f
C1060 VTAIL.n89 VSUBS 0.027897f
C1061 VTAIL.n90 VSUBS 0.037196f
C1062 VTAIL.n91 VSUBS 0.016662f
C1063 VTAIL.n92 VSUBS 0.015737f
C1064 VTAIL.n93 VSUBS 0.029286f
C1065 VTAIL.n94 VSUBS 0.029286f
C1066 VTAIL.n95 VSUBS 0.015737f
C1067 VTAIL.n96 VSUBS 0.016662f
C1068 VTAIL.n97 VSUBS 0.037196f
C1069 VTAIL.n98 VSUBS 0.037196f
C1070 VTAIL.n99 VSUBS 0.016662f
C1071 VTAIL.n100 VSUBS 0.015737f
C1072 VTAIL.n101 VSUBS 0.029286f
C1073 VTAIL.n102 VSUBS 0.029286f
C1074 VTAIL.n103 VSUBS 0.015737f
C1075 VTAIL.n104 VSUBS 0.016662f
C1076 VTAIL.n105 VSUBS 0.037196f
C1077 VTAIL.n106 VSUBS 0.092342f
C1078 VTAIL.n107 VSUBS 0.016662f
C1079 VTAIL.n108 VSUBS 0.030903f
C1080 VTAIL.n109 VSUBS 0.073693f
C1081 VTAIL.n110 VSUBS 0.070705f
C1082 VTAIL.n111 VSUBS 1.69119f
C1083 VTAIL.n112 VSUBS 0.03152f
C1084 VTAIL.n113 VSUBS 0.029286f
C1085 VTAIL.n114 VSUBS 0.015737f
C1086 VTAIL.n115 VSUBS 0.037196f
C1087 VTAIL.n116 VSUBS 0.016662f
C1088 VTAIL.n117 VSUBS 0.029286f
C1089 VTAIL.n118 VSUBS 0.015737f
C1090 VTAIL.n119 VSUBS 0.037196f
C1091 VTAIL.n120 VSUBS 0.016662f
C1092 VTAIL.n121 VSUBS 0.826415f
C1093 VTAIL.n122 VSUBS 0.015737f
C1094 VTAIL.t3 VSUBS 0.079902f
C1095 VTAIL.n123 VSUBS 0.16766f
C1096 VTAIL.n124 VSUBS 0.02798f
C1097 VTAIL.n125 VSUBS 0.027897f
C1098 VTAIL.n126 VSUBS 0.037196f
C1099 VTAIL.n127 VSUBS 0.016662f
C1100 VTAIL.n128 VSUBS 0.015737f
C1101 VTAIL.n129 VSUBS 0.029286f
C1102 VTAIL.n130 VSUBS 0.029286f
C1103 VTAIL.n131 VSUBS 0.015737f
C1104 VTAIL.n132 VSUBS 0.016662f
C1105 VTAIL.n133 VSUBS 0.037196f
C1106 VTAIL.n134 VSUBS 0.037196f
C1107 VTAIL.n135 VSUBS 0.016662f
C1108 VTAIL.n136 VSUBS 0.015737f
C1109 VTAIL.n137 VSUBS 0.029286f
C1110 VTAIL.n138 VSUBS 0.029286f
C1111 VTAIL.n139 VSUBS 0.015737f
C1112 VTAIL.n140 VSUBS 0.016662f
C1113 VTAIL.n141 VSUBS 0.037196f
C1114 VTAIL.n142 VSUBS 0.092342f
C1115 VTAIL.n143 VSUBS 0.016662f
C1116 VTAIL.n144 VSUBS 0.030903f
C1117 VTAIL.n145 VSUBS 0.073693f
C1118 VTAIL.n146 VSUBS 0.070705f
C1119 VTAIL.n147 VSUBS 1.69119f
C1120 VTAIL.t0 VSUBS 0.16732f
C1121 VTAIL.t6 VSUBS 0.16732f
C1122 VTAIL.n148 VSUBS 1.07436f
C1123 VTAIL.n149 VSUBS 1.22925f
C1124 VTAIL.n150 VSUBS 0.03152f
C1125 VTAIL.n151 VSUBS 0.029286f
C1126 VTAIL.n152 VSUBS 0.015737f
C1127 VTAIL.n153 VSUBS 0.037196f
C1128 VTAIL.n154 VSUBS 0.016662f
C1129 VTAIL.n155 VSUBS 0.029286f
C1130 VTAIL.n156 VSUBS 0.015737f
C1131 VTAIL.n157 VSUBS 0.037196f
C1132 VTAIL.n158 VSUBS 0.016662f
C1133 VTAIL.n159 VSUBS 0.826415f
C1134 VTAIL.n160 VSUBS 0.015737f
C1135 VTAIL.t5 VSUBS 0.079902f
C1136 VTAIL.n161 VSUBS 0.16766f
C1137 VTAIL.n162 VSUBS 0.02798f
C1138 VTAIL.n163 VSUBS 0.027897f
C1139 VTAIL.n164 VSUBS 0.037196f
C1140 VTAIL.n165 VSUBS 0.016662f
C1141 VTAIL.n166 VSUBS 0.015737f
C1142 VTAIL.n167 VSUBS 0.029286f
C1143 VTAIL.n168 VSUBS 0.029286f
C1144 VTAIL.n169 VSUBS 0.015737f
C1145 VTAIL.n170 VSUBS 0.016662f
C1146 VTAIL.n171 VSUBS 0.037196f
C1147 VTAIL.n172 VSUBS 0.037196f
C1148 VTAIL.n173 VSUBS 0.016662f
C1149 VTAIL.n174 VSUBS 0.015737f
C1150 VTAIL.n175 VSUBS 0.029286f
C1151 VTAIL.n176 VSUBS 0.029286f
C1152 VTAIL.n177 VSUBS 0.015737f
C1153 VTAIL.n178 VSUBS 0.016662f
C1154 VTAIL.n179 VSUBS 0.037196f
C1155 VTAIL.n180 VSUBS 0.092342f
C1156 VTAIL.n181 VSUBS 0.016662f
C1157 VTAIL.n182 VSUBS 0.030903f
C1158 VTAIL.n183 VSUBS 0.073693f
C1159 VTAIL.n184 VSUBS 0.070705f
C1160 VTAIL.n185 VSUBS 0.411153f
C1161 VTAIL.n186 VSUBS 0.03152f
C1162 VTAIL.n187 VSUBS 0.029286f
C1163 VTAIL.n188 VSUBS 0.015737f
C1164 VTAIL.n189 VSUBS 0.037196f
C1165 VTAIL.n190 VSUBS 0.016662f
C1166 VTAIL.n191 VSUBS 0.029286f
C1167 VTAIL.n192 VSUBS 0.015737f
C1168 VTAIL.n193 VSUBS 0.037196f
C1169 VTAIL.n194 VSUBS 0.016662f
C1170 VTAIL.n195 VSUBS 0.826415f
C1171 VTAIL.n196 VSUBS 0.015737f
C1172 VTAIL.t15 VSUBS 0.079902f
C1173 VTAIL.n197 VSUBS 0.16766f
C1174 VTAIL.n198 VSUBS 0.02798f
C1175 VTAIL.n199 VSUBS 0.027897f
C1176 VTAIL.n200 VSUBS 0.037196f
C1177 VTAIL.n201 VSUBS 0.016662f
C1178 VTAIL.n202 VSUBS 0.015737f
C1179 VTAIL.n203 VSUBS 0.029286f
C1180 VTAIL.n204 VSUBS 0.029286f
C1181 VTAIL.n205 VSUBS 0.015737f
C1182 VTAIL.n206 VSUBS 0.016662f
C1183 VTAIL.n207 VSUBS 0.037196f
C1184 VTAIL.n208 VSUBS 0.037196f
C1185 VTAIL.n209 VSUBS 0.016662f
C1186 VTAIL.n210 VSUBS 0.015737f
C1187 VTAIL.n211 VSUBS 0.029286f
C1188 VTAIL.n212 VSUBS 0.029286f
C1189 VTAIL.n213 VSUBS 0.015737f
C1190 VTAIL.n214 VSUBS 0.016662f
C1191 VTAIL.n215 VSUBS 0.037196f
C1192 VTAIL.n216 VSUBS 0.092342f
C1193 VTAIL.n217 VSUBS 0.016662f
C1194 VTAIL.n218 VSUBS 0.030903f
C1195 VTAIL.n219 VSUBS 0.073693f
C1196 VTAIL.n220 VSUBS 0.070705f
C1197 VTAIL.n221 VSUBS 0.411153f
C1198 VTAIL.t13 VSUBS 0.16732f
C1199 VTAIL.t14 VSUBS 0.16732f
C1200 VTAIL.n222 VSUBS 1.07436f
C1201 VTAIL.n223 VSUBS 1.22925f
C1202 VTAIL.n224 VSUBS 0.03152f
C1203 VTAIL.n225 VSUBS 0.029286f
C1204 VTAIL.n226 VSUBS 0.015737f
C1205 VTAIL.n227 VSUBS 0.037196f
C1206 VTAIL.n228 VSUBS 0.016662f
C1207 VTAIL.n229 VSUBS 0.029286f
C1208 VTAIL.n230 VSUBS 0.015737f
C1209 VTAIL.n231 VSUBS 0.037196f
C1210 VTAIL.n232 VSUBS 0.016662f
C1211 VTAIL.n233 VSUBS 0.826415f
C1212 VTAIL.n234 VSUBS 0.015737f
C1213 VTAIL.t12 VSUBS 0.079902f
C1214 VTAIL.n235 VSUBS 0.16766f
C1215 VTAIL.n236 VSUBS 0.02798f
C1216 VTAIL.n237 VSUBS 0.027897f
C1217 VTAIL.n238 VSUBS 0.037196f
C1218 VTAIL.n239 VSUBS 0.016662f
C1219 VTAIL.n240 VSUBS 0.015737f
C1220 VTAIL.n241 VSUBS 0.029286f
C1221 VTAIL.n242 VSUBS 0.029286f
C1222 VTAIL.n243 VSUBS 0.015737f
C1223 VTAIL.n244 VSUBS 0.016662f
C1224 VTAIL.n245 VSUBS 0.037196f
C1225 VTAIL.n246 VSUBS 0.037196f
C1226 VTAIL.n247 VSUBS 0.016662f
C1227 VTAIL.n248 VSUBS 0.015737f
C1228 VTAIL.n249 VSUBS 0.029286f
C1229 VTAIL.n250 VSUBS 0.029286f
C1230 VTAIL.n251 VSUBS 0.015737f
C1231 VTAIL.n252 VSUBS 0.016662f
C1232 VTAIL.n253 VSUBS 0.037196f
C1233 VTAIL.n254 VSUBS 0.092342f
C1234 VTAIL.n255 VSUBS 0.016662f
C1235 VTAIL.n256 VSUBS 0.030903f
C1236 VTAIL.n257 VSUBS 0.073693f
C1237 VTAIL.n258 VSUBS 0.070705f
C1238 VTAIL.n259 VSUBS 1.69119f
C1239 VTAIL.n260 VSUBS 0.03152f
C1240 VTAIL.n261 VSUBS 0.029286f
C1241 VTAIL.n262 VSUBS 0.015737f
C1242 VTAIL.n263 VSUBS 0.037196f
C1243 VTAIL.n264 VSUBS 0.016662f
C1244 VTAIL.n265 VSUBS 0.029286f
C1245 VTAIL.n266 VSUBS 0.015737f
C1246 VTAIL.n267 VSUBS 0.037196f
C1247 VTAIL.n268 VSUBS 0.016662f
C1248 VTAIL.n269 VSUBS 0.826415f
C1249 VTAIL.n270 VSUBS 0.015737f
C1250 VTAIL.t2 VSUBS 0.079902f
C1251 VTAIL.n271 VSUBS 0.16766f
C1252 VTAIL.n272 VSUBS 0.02798f
C1253 VTAIL.n273 VSUBS 0.027897f
C1254 VTAIL.n274 VSUBS 0.037196f
C1255 VTAIL.n275 VSUBS 0.016662f
C1256 VTAIL.n276 VSUBS 0.015737f
C1257 VTAIL.n277 VSUBS 0.029286f
C1258 VTAIL.n278 VSUBS 0.029286f
C1259 VTAIL.n279 VSUBS 0.015737f
C1260 VTAIL.n280 VSUBS 0.016662f
C1261 VTAIL.n281 VSUBS 0.037196f
C1262 VTAIL.n282 VSUBS 0.037196f
C1263 VTAIL.n283 VSUBS 0.016662f
C1264 VTAIL.n284 VSUBS 0.015737f
C1265 VTAIL.n285 VSUBS 0.029286f
C1266 VTAIL.n286 VSUBS 0.029286f
C1267 VTAIL.n287 VSUBS 0.015737f
C1268 VTAIL.n288 VSUBS 0.016662f
C1269 VTAIL.n289 VSUBS 0.037196f
C1270 VTAIL.n290 VSUBS 0.092342f
C1271 VTAIL.n291 VSUBS 0.016662f
C1272 VTAIL.n292 VSUBS 0.030903f
C1273 VTAIL.n293 VSUBS 0.073693f
C1274 VTAIL.n294 VSUBS 0.070705f
C1275 VTAIL.n295 VSUBS 1.6857f
C1276 VDD1.t1 VSUBS 0.188728f
C1277 VDD1.t6 VSUBS 0.188728f
C1278 VDD1.n0 VSUBS 1.36104f
C1279 VDD1.t7 VSUBS 0.188728f
C1280 VDD1.t4 VSUBS 0.188728f
C1281 VDD1.n1 VSUBS 1.3594f
C1282 VDD1.t0 VSUBS 0.188728f
C1283 VDD1.t3 VSUBS 0.188728f
C1284 VDD1.n2 VSUBS 1.3594f
C1285 VDD1.n3 VSUBS 5.48683f
C1286 VDD1.t2 VSUBS 0.188728f
C1287 VDD1.t5 VSUBS 0.188728f
C1288 VDD1.n4 VSUBS 1.3376f
C1289 VDD1.n5 VSUBS 4.29334f
C1290 VP.n0 VSUBS 0.060744f
C1291 VP.t6 VSUBS 2.39052f
C1292 VP.n1 VSUBS 0.064957f
C1293 VP.n2 VSUBS 0.032293f
C1294 VP.n3 VSUBS 0.060187f
C1295 VP.n4 VSUBS 0.032293f
C1296 VP.t5 VSUBS 2.39052f
C1297 VP.n5 VSUBS 0.060187f
C1298 VP.n6 VSUBS 0.032293f
C1299 VP.n7 VSUBS 0.060187f
C1300 VP.n8 VSUBS 0.032293f
C1301 VP.t7 VSUBS 2.39052f
C1302 VP.n9 VSUBS 0.060187f
C1303 VP.n10 VSUBS 0.032293f
C1304 VP.n11 VSUBS 0.060187f
C1305 VP.n12 VSUBS 0.060744f
C1306 VP.t3 VSUBS 2.39052f
C1307 VP.n13 VSUBS 0.064957f
C1308 VP.n14 VSUBS 0.032293f
C1309 VP.n15 VSUBS 0.060187f
C1310 VP.n16 VSUBS 0.032293f
C1311 VP.t1 VSUBS 2.39052f
C1312 VP.n17 VSUBS 0.060187f
C1313 VP.n18 VSUBS 0.032293f
C1314 VP.n19 VSUBS 0.060187f
C1315 VP.t0 VSUBS 2.85448f
C1316 VP.n20 VSUBS 0.952078f
C1317 VP.t2 VSUBS 2.39052f
C1318 VP.n21 VSUBS 0.986275f
C1319 VP.n22 VSUBS 0.050084f
C1320 VP.n23 VSUBS 0.41905f
C1321 VP.n24 VSUBS 0.032293f
C1322 VP.n25 VSUBS 0.032293f
C1323 VP.n26 VSUBS 0.060187f
C1324 VP.n27 VSUBS 0.047143f
C1325 VP.n28 VSUBS 0.047143f
C1326 VP.n29 VSUBS 0.032293f
C1327 VP.n30 VSUBS 0.032293f
C1328 VP.n31 VSUBS 0.032293f
C1329 VP.n32 VSUBS 0.060187f
C1330 VP.n33 VSUBS 0.050084f
C1331 VP.n34 VSUBS 0.865067f
C1332 VP.n35 VSUBS 0.040575f
C1333 VP.n36 VSUBS 0.032293f
C1334 VP.n37 VSUBS 0.032293f
C1335 VP.n38 VSUBS 0.032293f
C1336 VP.n39 VSUBS 0.060187f
C1337 VP.n40 VSUBS 0.059885f
C1338 VP.n41 VSUBS 0.02963f
C1339 VP.n42 VSUBS 0.032293f
C1340 VP.n43 VSUBS 0.032293f
C1341 VP.n44 VSUBS 0.032293f
C1342 VP.n45 VSUBS 0.060187f
C1343 VP.n46 VSUBS 0.059592f
C1344 VP.n47 VSUBS 1.01161f
C1345 VP.n48 VSUBS 2.04574f
C1346 VP.n49 VSUBS 2.06752f
C1347 VP.t4 VSUBS 2.39052f
C1348 VP.n50 VSUBS 1.01161f
C1349 VP.n51 VSUBS 0.059592f
C1350 VP.n52 VSUBS 0.060744f
C1351 VP.n53 VSUBS 0.032293f
C1352 VP.n54 VSUBS 0.032293f
C1353 VP.n55 VSUBS 0.064957f
C1354 VP.n56 VSUBS 0.02963f
C1355 VP.n57 VSUBS 0.059885f
C1356 VP.n58 VSUBS 0.032293f
C1357 VP.n59 VSUBS 0.032293f
C1358 VP.n60 VSUBS 0.032293f
C1359 VP.n61 VSUBS 0.060187f
C1360 VP.n62 VSUBS 0.040575f
C1361 VP.n63 VSUBS 0.865067f
C1362 VP.n64 VSUBS 0.050084f
C1363 VP.n65 VSUBS 0.032293f
C1364 VP.n66 VSUBS 0.032293f
C1365 VP.n67 VSUBS 0.032293f
C1366 VP.n68 VSUBS 0.060187f
C1367 VP.n69 VSUBS 0.047143f
C1368 VP.n70 VSUBS 0.047143f
C1369 VP.n71 VSUBS 0.032293f
C1370 VP.n72 VSUBS 0.032293f
C1371 VP.n73 VSUBS 0.032293f
C1372 VP.n74 VSUBS 0.060187f
C1373 VP.n75 VSUBS 0.050084f
C1374 VP.n76 VSUBS 0.865067f
C1375 VP.n77 VSUBS 0.040575f
C1376 VP.n78 VSUBS 0.032293f
C1377 VP.n79 VSUBS 0.032293f
C1378 VP.n80 VSUBS 0.032293f
C1379 VP.n81 VSUBS 0.060187f
C1380 VP.n82 VSUBS 0.059885f
C1381 VP.n83 VSUBS 0.02963f
C1382 VP.n84 VSUBS 0.032293f
C1383 VP.n85 VSUBS 0.032293f
C1384 VP.n86 VSUBS 0.032293f
C1385 VP.n87 VSUBS 0.060187f
C1386 VP.n88 VSUBS 0.059592f
C1387 VP.n89 VSUBS 1.01161f
C1388 VP.n90 VSUBS 0.093927f
.ends

