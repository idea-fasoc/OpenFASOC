* NGSPICE file created from diff_pair_sample_0646.ext - technology: sky130A

.subckt diff_pair_sample_0646 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 w_n1530_n3732# sky130_fd_pr__pfet_01v8 ad=5.382 pd=28.38 as=5.382 ps=28.38 w=13.8 l=1.07
X1 B.t11 B.t9 B.t10 w_n1530_n3732# sky130_fd_pr__pfet_01v8 ad=5.382 pd=28.38 as=0 ps=0 w=13.8 l=1.07
X2 VDD1.t1 VP.t0 VTAIL.t0 w_n1530_n3732# sky130_fd_pr__pfet_01v8 ad=5.382 pd=28.38 as=5.382 ps=28.38 w=13.8 l=1.07
X3 B.t8 B.t6 B.t7 w_n1530_n3732# sky130_fd_pr__pfet_01v8 ad=5.382 pd=28.38 as=0 ps=0 w=13.8 l=1.07
X4 VDD1.t0 VP.t1 VTAIL.t1 w_n1530_n3732# sky130_fd_pr__pfet_01v8 ad=5.382 pd=28.38 as=5.382 ps=28.38 w=13.8 l=1.07
X5 B.t5 B.t3 B.t4 w_n1530_n3732# sky130_fd_pr__pfet_01v8 ad=5.382 pd=28.38 as=0 ps=0 w=13.8 l=1.07
X6 VDD2.t0 VN.t1 VTAIL.t2 w_n1530_n3732# sky130_fd_pr__pfet_01v8 ad=5.382 pd=28.38 as=5.382 ps=28.38 w=13.8 l=1.07
X7 B.t2 B.t0 B.t1 w_n1530_n3732# sky130_fd_pr__pfet_01v8 ad=5.382 pd=28.38 as=0 ps=0 w=13.8 l=1.07
R0 VN VN.t1 551.644
R1 VN VN.t0 509.337
R2 VTAIL.n2 VTAIL.t1 55.2965
R3 VTAIL.n1 VTAIL.t2 55.2965
R4 VTAIL.n3 VTAIL.t3 55.2964
R5 VTAIL.n0 VTAIL.t0 55.2964
R6 VTAIL.n1 VTAIL.n0 26.6945
R7 VTAIL.n3 VTAIL.n2 25.4876
R8 VTAIL.n2 VTAIL.n1 1.07378
R9 VTAIL VTAIL.n0 0.830241
R10 VTAIL VTAIL.n3 0.244034
R11 VDD2.n0 VDD2.t1 109.963
R12 VDD2.n0 VDD2.t0 71.9753
R13 VDD2 VDD2.n0 0.360414
R14 B.n327 B.n84 585
R15 B.n326 B.n325 585
R16 B.n324 B.n85 585
R17 B.n323 B.n322 585
R18 B.n321 B.n86 585
R19 B.n320 B.n319 585
R20 B.n318 B.n87 585
R21 B.n317 B.n316 585
R22 B.n315 B.n88 585
R23 B.n314 B.n313 585
R24 B.n312 B.n89 585
R25 B.n311 B.n310 585
R26 B.n309 B.n90 585
R27 B.n308 B.n307 585
R28 B.n306 B.n91 585
R29 B.n305 B.n304 585
R30 B.n303 B.n92 585
R31 B.n302 B.n301 585
R32 B.n300 B.n93 585
R33 B.n299 B.n298 585
R34 B.n297 B.n94 585
R35 B.n296 B.n295 585
R36 B.n294 B.n95 585
R37 B.n293 B.n292 585
R38 B.n291 B.n96 585
R39 B.n290 B.n289 585
R40 B.n288 B.n97 585
R41 B.n287 B.n286 585
R42 B.n285 B.n98 585
R43 B.n284 B.n283 585
R44 B.n282 B.n99 585
R45 B.n281 B.n280 585
R46 B.n279 B.n100 585
R47 B.n278 B.n277 585
R48 B.n276 B.n101 585
R49 B.n275 B.n274 585
R50 B.n273 B.n102 585
R51 B.n272 B.n271 585
R52 B.n270 B.n103 585
R53 B.n269 B.n268 585
R54 B.n267 B.n104 585
R55 B.n266 B.n265 585
R56 B.n264 B.n105 585
R57 B.n263 B.n262 585
R58 B.n261 B.n106 585
R59 B.n260 B.n259 585
R60 B.n258 B.n107 585
R61 B.n257 B.n256 585
R62 B.n252 B.n108 585
R63 B.n251 B.n250 585
R64 B.n249 B.n109 585
R65 B.n248 B.n247 585
R66 B.n246 B.n110 585
R67 B.n245 B.n244 585
R68 B.n243 B.n111 585
R69 B.n242 B.n241 585
R70 B.n240 B.n112 585
R71 B.n238 B.n237 585
R72 B.n236 B.n115 585
R73 B.n235 B.n234 585
R74 B.n233 B.n116 585
R75 B.n232 B.n231 585
R76 B.n230 B.n117 585
R77 B.n229 B.n228 585
R78 B.n227 B.n118 585
R79 B.n226 B.n225 585
R80 B.n224 B.n119 585
R81 B.n223 B.n222 585
R82 B.n221 B.n120 585
R83 B.n220 B.n219 585
R84 B.n218 B.n121 585
R85 B.n217 B.n216 585
R86 B.n215 B.n122 585
R87 B.n214 B.n213 585
R88 B.n212 B.n123 585
R89 B.n211 B.n210 585
R90 B.n209 B.n124 585
R91 B.n208 B.n207 585
R92 B.n206 B.n125 585
R93 B.n205 B.n204 585
R94 B.n203 B.n126 585
R95 B.n202 B.n201 585
R96 B.n200 B.n127 585
R97 B.n199 B.n198 585
R98 B.n197 B.n128 585
R99 B.n196 B.n195 585
R100 B.n194 B.n129 585
R101 B.n193 B.n192 585
R102 B.n191 B.n130 585
R103 B.n190 B.n189 585
R104 B.n188 B.n131 585
R105 B.n187 B.n186 585
R106 B.n185 B.n132 585
R107 B.n184 B.n183 585
R108 B.n182 B.n133 585
R109 B.n181 B.n180 585
R110 B.n179 B.n134 585
R111 B.n178 B.n177 585
R112 B.n176 B.n135 585
R113 B.n175 B.n174 585
R114 B.n173 B.n136 585
R115 B.n172 B.n171 585
R116 B.n170 B.n137 585
R117 B.n169 B.n168 585
R118 B.n329 B.n328 585
R119 B.n330 B.n83 585
R120 B.n332 B.n331 585
R121 B.n333 B.n82 585
R122 B.n335 B.n334 585
R123 B.n336 B.n81 585
R124 B.n338 B.n337 585
R125 B.n339 B.n80 585
R126 B.n341 B.n340 585
R127 B.n342 B.n79 585
R128 B.n344 B.n343 585
R129 B.n345 B.n78 585
R130 B.n347 B.n346 585
R131 B.n348 B.n77 585
R132 B.n350 B.n349 585
R133 B.n351 B.n76 585
R134 B.n353 B.n352 585
R135 B.n354 B.n75 585
R136 B.n356 B.n355 585
R137 B.n357 B.n74 585
R138 B.n359 B.n358 585
R139 B.n360 B.n73 585
R140 B.n362 B.n361 585
R141 B.n363 B.n72 585
R142 B.n365 B.n364 585
R143 B.n366 B.n71 585
R144 B.n368 B.n367 585
R145 B.n369 B.n70 585
R146 B.n371 B.n370 585
R147 B.n372 B.n69 585
R148 B.n374 B.n373 585
R149 B.n375 B.n68 585
R150 B.n377 B.n376 585
R151 B.n378 B.n67 585
R152 B.n535 B.n10 585
R153 B.n534 B.n533 585
R154 B.n532 B.n11 585
R155 B.n531 B.n530 585
R156 B.n529 B.n12 585
R157 B.n528 B.n527 585
R158 B.n526 B.n13 585
R159 B.n525 B.n524 585
R160 B.n523 B.n14 585
R161 B.n522 B.n521 585
R162 B.n520 B.n15 585
R163 B.n519 B.n518 585
R164 B.n517 B.n16 585
R165 B.n516 B.n515 585
R166 B.n514 B.n17 585
R167 B.n513 B.n512 585
R168 B.n511 B.n18 585
R169 B.n510 B.n509 585
R170 B.n508 B.n19 585
R171 B.n507 B.n506 585
R172 B.n505 B.n20 585
R173 B.n504 B.n503 585
R174 B.n502 B.n21 585
R175 B.n501 B.n500 585
R176 B.n499 B.n22 585
R177 B.n498 B.n497 585
R178 B.n496 B.n23 585
R179 B.n495 B.n494 585
R180 B.n493 B.n24 585
R181 B.n492 B.n491 585
R182 B.n490 B.n25 585
R183 B.n489 B.n488 585
R184 B.n487 B.n26 585
R185 B.n486 B.n485 585
R186 B.n484 B.n27 585
R187 B.n483 B.n482 585
R188 B.n481 B.n28 585
R189 B.n480 B.n479 585
R190 B.n478 B.n29 585
R191 B.n477 B.n476 585
R192 B.n475 B.n30 585
R193 B.n474 B.n473 585
R194 B.n472 B.n31 585
R195 B.n471 B.n470 585
R196 B.n469 B.n32 585
R197 B.n468 B.n467 585
R198 B.n466 B.n33 585
R199 B.n464 B.n463 585
R200 B.n462 B.n36 585
R201 B.n461 B.n460 585
R202 B.n459 B.n37 585
R203 B.n458 B.n457 585
R204 B.n456 B.n38 585
R205 B.n455 B.n454 585
R206 B.n453 B.n39 585
R207 B.n452 B.n451 585
R208 B.n450 B.n40 585
R209 B.n449 B.n448 585
R210 B.n447 B.n41 585
R211 B.n446 B.n445 585
R212 B.n444 B.n45 585
R213 B.n443 B.n442 585
R214 B.n441 B.n46 585
R215 B.n440 B.n439 585
R216 B.n438 B.n47 585
R217 B.n437 B.n436 585
R218 B.n435 B.n48 585
R219 B.n434 B.n433 585
R220 B.n432 B.n49 585
R221 B.n431 B.n430 585
R222 B.n429 B.n50 585
R223 B.n428 B.n427 585
R224 B.n426 B.n51 585
R225 B.n425 B.n424 585
R226 B.n423 B.n52 585
R227 B.n422 B.n421 585
R228 B.n420 B.n53 585
R229 B.n419 B.n418 585
R230 B.n417 B.n54 585
R231 B.n416 B.n415 585
R232 B.n414 B.n55 585
R233 B.n413 B.n412 585
R234 B.n411 B.n56 585
R235 B.n410 B.n409 585
R236 B.n408 B.n57 585
R237 B.n407 B.n406 585
R238 B.n405 B.n58 585
R239 B.n404 B.n403 585
R240 B.n402 B.n59 585
R241 B.n401 B.n400 585
R242 B.n399 B.n60 585
R243 B.n398 B.n397 585
R244 B.n396 B.n61 585
R245 B.n395 B.n394 585
R246 B.n393 B.n62 585
R247 B.n392 B.n391 585
R248 B.n390 B.n63 585
R249 B.n389 B.n388 585
R250 B.n387 B.n64 585
R251 B.n386 B.n385 585
R252 B.n384 B.n65 585
R253 B.n383 B.n382 585
R254 B.n381 B.n66 585
R255 B.n380 B.n379 585
R256 B.n537 B.n536 585
R257 B.n538 B.n9 585
R258 B.n540 B.n539 585
R259 B.n541 B.n8 585
R260 B.n543 B.n542 585
R261 B.n544 B.n7 585
R262 B.n546 B.n545 585
R263 B.n547 B.n6 585
R264 B.n549 B.n548 585
R265 B.n550 B.n5 585
R266 B.n552 B.n551 585
R267 B.n553 B.n4 585
R268 B.n555 B.n554 585
R269 B.n556 B.n3 585
R270 B.n558 B.n557 585
R271 B.n559 B.n0 585
R272 B.n2 B.n1 585
R273 B.n146 B.n145 585
R274 B.n148 B.n147 585
R275 B.n149 B.n144 585
R276 B.n151 B.n150 585
R277 B.n152 B.n143 585
R278 B.n154 B.n153 585
R279 B.n155 B.n142 585
R280 B.n157 B.n156 585
R281 B.n158 B.n141 585
R282 B.n160 B.n159 585
R283 B.n161 B.n140 585
R284 B.n163 B.n162 585
R285 B.n164 B.n139 585
R286 B.n166 B.n165 585
R287 B.n167 B.n138 585
R288 B.n113 B.t3 514.202
R289 B.n253 B.t9 514.202
R290 B.n42 B.t6 514.202
R291 B.n34 B.t0 514.202
R292 B.n169 B.n138 434.841
R293 B.n329 B.n84 434.841
R294 B.n379 B.n378 434.841
R295 B.n536 B.n535 434.841
R296 B.n561 B.n560 256.663
R297 B.n560 B.n559 235.042
R298 B.n560 B.n2 235.042
R299 B.n170 B.n169 163.367
R300 B.n171 B.n170 163.367
R301 B.n171 B.n136 163.367
R302 B.n175 B.n136 163.367
R303 B.n176 B.n175 163.367
R304 B.n177 B.n176 163.367
R305 B.n177 B.n134 163.367
R306 B.n181 B.n134 163.367
R307 B.n182 B.n181 163.367
R308 B.n183 B.n182 163.367
R309 B.n183 B.n132 163.367
R310 B.n187 B.n132 163.367
R311 B.n188 B.n187 163.367
R312 B.n189 B.n188 163.367
R313 B.n189 B.n130 163.367
R314 B.n193 B.n130 163.367
R315 B.n194 B.n193 163.367
R316 B.n195 B.n194 163.367
R317 B.n195 B.n128 163.367
R318 B.n199 B.n128 163.367
R319 B.n200 B.n199 163.367
R320 B.n201 B.n200 163.367
R321 B.n201 B.n126 163.367
R322 B.n205 B.n126 163.367
R323 B.n206 B.n205 163.367
R324 B.n207 B.n206 163.367
R325 B.n207 B.n124 163.367
R326 B.n211 B.n124 163.367
R327 B.n212 B.n211 163.367
R328 B.n213 B.n212 163.367
R329 B.n213 B.n122 163.367
R330 B.n217 B.n122 163.367
R331 B.n218 B.n217 163.367
R332 B.n219 B.n218 163.367
R333 B.n219 B.n120 163.367
R334 B.n223 B.n120 163.367
R335 B.n224 B.n223 163.367
R336 B.n225 B.n224 163.367
R337 B.n225 B.n118 163.367
R338 B.n229 B.n118 163.367
R339 B.n230 B.n229 163.367
R340 B.n231 B.n230 163.367
R341 B.n231 B.n116 163.367
R342 B.n235 B.n116 163.367
R343 B.n236 B.n235 163.367
R344 B.n237 B.n236 163.367
R345 B.n237 B.n112 163.367
R346 B.n242 B.n112 163.367
R347 B.n243 B.n242 163.367
R348 B.n244 B.n243 163.367
R349 B.n244 B.n110 163.367
R350 B.n248 B.n110 163.367
R351 B.n249 B.n248 163.367
R352 B.n250 B.n249 163.367
R353 B.n250 B.n108 163.367
R354 B.n257 B.n108 163.367
R355 B.n258 B.n257 163.367
R356 B.n259 B.n258 163.367
R357 B.n259 B.n106 163.367
R358 B.n263 B.n106 163.367
R359 B.n264 B.n263 163.367
R360 B.n265 B.n264 163.367
R361 B.n265 B.n104 163.367
R362 B.n269 B.n104 163.367
R363 B.n270 B.n269 163.367
R364 B.n271 B.n270 163.367
R365 B.n271 B.n102 163.367
R366 B.n275 B.n102 163.367
R367 B.n276 B.n275 163.367
R368 B.n277 B.n276 163.367
R369 B.n277 B.n100 163.367
R370 B.n281 B.n100 163.367
R371 B.n282 B.n281 163.367
R372 B.n283 B.n282 163.367
R373 B.n283 B.n98 163.367
R374 B.n287 B.n98 163.367
R375 B.n288 B.n287 163.367
R376 B.n289 B.n288 163.367
R377 B.n289 B.n96 163.367
R378 B.n293 B.n96 163.367
R379 B.n294 B.n293 163.367
R380 B.n295 B.n294 163.367
R381 B.n295 B.n94 163.367
R382 B.n299 B.n94 163.367
R383 B.n300 B.n299 163.367
R384 B.n301 B.n300 163.367
R385 B.n301 B.n92 163.367
R386 B.n305 B.n92 163.367
R387 B.n306 B.n305 163.367
R388 B.n307 B.n306 163.367
R389 B.n307 B.n90 163.367
R390 B.n311 B.n90 163.367
R391 B.n312 B.n311 163.367
R392 B.n313 B.n312 163.367
R393 B.n313 B.n88 163.367
R394 B.n317 B.n88 163.367
R395 B.n318 B.n317 163.367
R396 B.n319 B.n318 163.367
R397 B.n319 B.n86 163.367
R398 B.n323 B.n86 163.367
R399 B.n324 B.n323 163.367
R400 B.n325 B.n324 163.367
R401 B.n325 B.n84 163.367
R402 B.n378 B.n377 163.367
R403 B.n377 B.n68 163.367
R404 B.n373 B.n68 163.367
R405 B.n373 B.n372 163.367
R406 B.n372 B.n371 163.367
R407 B.n371 B.n70 163.367
R408 B.n367 B.n70 163.367
R409 B.n367 B.n366 163.367
R410 B.n366 B.n365 163.367
R411 B.n365 B.n72 163.367
R412 B.n361 B.n72 163.367
R413 B.n361 B.n360 163.367
R414 B.n360 B.n359 163.367
R415 B.n359 B.n74 163.367
R416 B.n355 B.n74 163.367
R417 B.n355 B.n354 163.367
R418 B.n354 B.n353 163.367
R419 B.n353 B.n76 163.367
R420 B.n349 B.n76 163.367
R421 B.n349 B.n348 163.367
R422 B.n348 B.n347 163.367
R423 B.n347 B.n78 163.367
R424 B.n343 B.n78 163.367
R425 B.n343 B.n342 163.367
R426 B.n342 B.n341 163.367
R427 B.n341 B.n80 163.367
R428 B.n337 B.n80 163.367
R429 B.n337 B.n336 163.367
R430 B.n336 B.n335 163.367
R431 B.n335 B.n82 163.367
R432 B.n331 B.n82 163.367
R433 B.n331 B.n330 163.367
R434 B.n330 B.n329 163.367
R435 B.n535 B.n534 163.367
R436 B.n534 B.n11 163.367
R437 B.n530 B.n11 163.367
R438 B.n530 B.n529 163.367
R439 B.n529 B.n528 163.367
R440 B.n528 B.n13 163.367
R441 B.n524 B.n13 163.367
R442 B.n524 B.n523 163.367
R443 B.n523 B.n522 163.367
R444 B.n522 B.n15 163.367
R445 B.n518 B.n15 163.367
R446 B.n518 B.n517 163.367
R447 B.n517 B.n516 163.367
R448 B.n516 B.n17 163.367
R449 B.n512 B.n17 163.367
R450 B.n512 B.n511 163.367
R451 B.n511 B.n510 163.367
R452 B.n510 B.n19 163.367
R453 B.n506 B.n19 163.367
R454 B.n506 B.n505 163.367
R455 B.n505 B.n504 163.367
R456 B.n504 B.n21 163.367
R457 B.n500 B.n21 163.367
R458 B.n500 B.n499 163.367
R459 B.n499 B.n498 163.367
R460 B.n498 B.n23 163.367
R461 B.n494 B.n23 163.367
R462 B.n494 B.n493 163.367
R463 B.n493 B.n492 163.367
R464 B.n492 B.n25 163.367
R465 B.n488 B.n25 163.367
R466 B.n488 B.n487 163.367
R467 B.n487 B.n486 163.367
R468 B.n486 B.n27 163.367
R469 B.n482 B.n27 163.367
R470 B.n482 B.n481 163.367
R471 B.n481 B.n480 163.367
R472 B.n480 B.n29 163.367
R473 B.n476 B.n29 163.367
R474 B.n476 B.n475 163.367
R475 B.n475 B.n474 163.367
R476 B.n474 B.n31 163.367
R477 B.n470 B.n31 163.367
R478 B.n470 B.n469 163.367
R479 B.n469 B.n468 163.367
R480 B.n468 B.n33 163.367
R481 B.n463 B.n33 163.367
R482 B.n463 B.n462 163.367
R483 B.n462 B.n461 163.367
R484 B.n461 B.n37 163.367
R485 B.n457 B.n37 163.367
R486 B.n457 B.n456 163.367
R487 B.n456 B.n455 163.367
R488 B.n455 B.n39 163.367
R489 B.n451 B.n39 163.367
R490 B.n451 B.n450 163.367
R491 B.n450 B.n449 163.367
R492 B.n449 B.n41 163.367
R493 B.n445 B.n41 163.367
R494 B.n445 B.n444 163.367
R495 B.n444 B.n443 163.367
R496 B.n443 B.n46 163.367
R497 B.n439 B.n46 163.367
R498 B.n439 B.n438 163.367
R499 B.n438 B.n437 163.367
R500 B.n437 B.n48 163.367
R501 B.n433 B.n48 163.367
R502 B.n433 B.n432 163.367
R503 B.n432 B.n431 163.367
R504 B.n431 B.n50 163.367
R505 B.n427 B.n50 163.367
R506 B.n427 B.n426 163.367
R507 B.n426 B.n425 163.367
R508 B.n425 B.n52 163.367
R509 B.n421 B.n52 163.367
R510 B.n421 B.n420 163.367
R511 B.n420 B.n419 163.367
R512 B.n419 B.n54 163.367
R513 B.n415 B.n54 163.367
R514 B.n415 B.n414 163.367
R515 B.n414 B.n413 163.367
R516 B.n413 B.n56 163.367
R517 B.n409 B.n56 163.367
R518 B.n409 B.n408 163.367
R519 B.n408 B.n407 163.367
R520 B.n407 B.n58 163.367
R521 B.n403 B.n58 163.367
R522 B.n403 B.n402 163.367
R523 B.n402 B.n401 163.367
R524 B.n401 B.n60 163.367
R525 B.n397 B.n60 163.367
R526 B.n397 B.n396 163.367
R527 B.n396 B.n395 163.367
R528 B.n395 B.n62 163.367
R529 B.n391 B.n62 163.367
R530 B.n391 B.n390 163.367
R531 B.n390 B.n389 163.367
R532 B.n389 B.n64 163.367
R533 B.n385 B.n64 163.367
R534 B.n385 B.n384 163.367
R535 B.n384 B.n383 163.367
R536 B.n383 B.n66 163.367
R537 B.n379 B.n66 163.367
R538 B.n536 B.n9 163.367
R539 B.n540 B.n9 163.367
R540 B.n541 B.n540 163.367
R541 B.n542 B.n541 163.367
R542 B.n542 B.n7 163.367
R543 B.n546 B.n7 163.367
R544 B.n547 B.n546 163.367
R545 B.n548 B.n547 163.367
R546 B.n548 B.n5 163.367
R547 B.n552 B.n5 163.367
R548 B.n553 B.n552 163.367
R549 B.n554 B.n553 163.367
R550 B.n554 B.n3 163.367
R551 B.n558 B.n3 163.367
R552 B.n559 B.n558 163.367
R553 B.n146 B.n2 163.367
R554 B.n147 B.n146 163.367
R555 B.n147 B.n144 163.367
R556 B.n151 B.n144 163.367
R557 B.n152 B.n151 163.367
R558 B.n153 B.n152 163.367
R559 B.n153 B.n142 163.367
R560 B.n157 B.n142 163.367
R561 B.n158 B.n157 163.367
R562 B.n159 B.n158 163.367
R563 B.n159 B.n140 163.367
R564 B.n163 B.n140 163.367
R565 B.n164 B.n163 163.367
R566 B.n165 B.n164 163.367
R567 B.n165 B.n138 163.367
R568 B.n253 B.t10 137.78
R569 B.n42 B.t8 137.78
R570 B.n113 B.t4 137.762
R571 B.n34 B.t2 137.762
R572 B.n254 B.t11 110.627
R573 B.n43 B.t7 110.627
R574 B.n114 B.t5 110.611
R575 B.n35 B.t1 110.611
R576 B.n239 B.n114 59.5399
R577 B.n255 B.n254 59.5399
R578 B.n44 B.n43 59.5399
R579 B.n465 B.n35 59.5399
R580 B.n328 B.n327 28.2542
R581 B.n537 B.n10 28.2542
R582 B.n380 B.n67 28.2542
R583 B.n168 B.n167 28.2542
R584 B.n114 B.n113 27.152
R585 B.n254 B.n253 27.152
R586 B.n43 B.n42 27.152
R587 B.n35 B.n34 27.152
R588 B B.n561 18.0485
R589 B.n538 B.n537 10.6151
R590 B.n539 B.n538 10.6151
R591 B.n539 B.n8 10.6151
R592 B.n543 B.n8 10.6151
R593 B.n544 B.n543 10.6151
R594 B.n545 B.n544 10.6151
R595 B.n545 B.n6 10.6151
R596 B.n549 B.n6 10.6151
R597 B.n550 B.n549 10.6151
R598 B.n551 B.n550 10.6151
R599 B.n551 B.n4 10.6151
R600 B.n555 B.n4 10.6151
R601 B.n556 B.n555 10.6151
R602 B.n557 B.n556 10.6151
R603 B.n557 B.n0 10.6151
R604 B.n533 B.n10 10.6151
R605 B.n533 B.n532 10.6151
R606 B.n532 B.n531 10.6151
R607 B.n531 B.n12 10.6151
R608 B.n527 B.n12 10.6151
R609 B.n527 B.n526 10.6151
R610 B.n526 B.n525 10.6151
R611 B.n525 B.n14 10.6151
R612 B.n521 B.n14 10.6151
R613 B.n521 B.n520 10.6151
R614 B.n520 B.n519 10.6151
R615 B.n519 B.n16 10.6151
R616 B.n515 B.n16 10.6151
R617 B.n515 B.n514 10.6151
R618 B.n514 B.n513 10.6151
R619 B.n513 B.n18 10.6151
R620 B.n509 B.n18 10.6151
R621 B.n509 B.n508 10.6151
R622 B.n508 B.n507 10.6151
R623 B.n507 B.n20 10.6151
R624 B.n503 B.n20 10.6151
R625 B.n503 B.n502 10.6151
R626 B.n502 B.n501 10.6151
R627 B.n501 B.n22 10.6151
R628 B.n497 B.n22 10.6151
R629 B.n497 B.n496 10.6151
R630 B.n496 B.n495 10.6151
R631 B.n495 B.n24 10.6151
R632 B.n491 B.n24 10.6151
R633 B.n491 B.n490 10.6151
R634 B.n490 B.n489 10.6151
R635 B.n489 B.n26 10.6151
R636 B.n485 B.n26 10.6151
R637 B.n485 B.n484 10.6151
R638 B.n484 B.n483 10.6151
R639 B.n483 B.n28 10.6151
R640 B.n479 B.n28 10.6151
R641 B.n479 B.n478 10.6151
R642 B.n478 B.n477 10.6151
R643 B.n477 B.n30 10.6151
R644 B.n473 B.n30 10.6151
R645 B.n473 B.n472 10.6151
R646 B.n472 B.n471 10.6151
R647 B.n471 B.n32 10.6151
R648 B.n467 B.n32 10.6151
R649 B.n467 B.n466 10.6151
R650 B.n464 B.n36 10.6151
R651 B.n460 B.n36 10.6151
R652 B.n460 B.n459 10.6151
R653 B.n459 B.n458 10.6151
R654 B.n458 B.n38 10.6151
R655 B.n454 B.n38 10.6151
R656 B.n454 B.n453 10.6151
R657 B.n453 B.n452 10.6151
R658 B.n452 B.n40 10.6151
R659 B.n448 B.n447 10.6151
R660 B.n447 B.n446 10.6151
R661 B.n446 B.n45 10.6151
R662 B.n442 B.n45 10.6151
R663 B.n442 B.n441 10.6151
R664 B.n441 B.n440 10.6151
R665 B.n440 B.n47 10.6151
R666 B.n436 B.n47 10.6151
R667 B.n436 B.n435 10.6151
R668 B.n435 B.n434 10.6151
R669 B.n434 B.n49 10.6151
R670 B.n430 B.n49 10.6151
R671 B.n430 B.n429 10.6151
R672 B.n429 B.n428 10.6151
R673 B.n428 B.n51 10.6151
R674 B.n424 B.n51 10.6151
R675 B.n424 B.n423 10.6151
R676 B.n423 B.n422 10.6151
R677 B.n422 B.n53 10.6151
R678 B.n418 B.n53 10.6151
R679 B.n418 B.n417 10.6151
R680 B.n417 B.n416 10.6151
R681 B.n416 B.n55 10.6151
R682 B.n412 B.n55 10.6151
R683 B.n412 B.n411 10.6151
R684 B.n411 B.n410 10.6151
R685 B.n410 B.n57 10.6151
R686 B.n406 B.n57 10.6151
R687 B.n406 B.n405 10.6151
R688 B.n405 B.n404 10.6151
R689 B.n404 B.n59 10.6151
R690 B.n400 B.n59 10.6151
R691 B.n400 B.n399 10.6151
R692 B.n399 B.n398 10.6151
R693 B.n398 B.n61 10.6151
R694 B.n394 B.n61 10.6151
R695 B.n394 B.n393 10.6151
R696 B.n393 B.n392 10.6151
R697 B.n392 B.n63 10.6151
R698 B.n388 B.n63 10.6151
R699 B.n388 B.n387 10.6151
R700 B.n387 B.n386 10.6151
R701 B.n386 B.n65 10.6151
R702 B.n382 B.n65 10.6151
R703 B.n382 B.n381 10.6151
R704 B.n381 B.n380 10.6151
R705 B.n376 B.n67 10.6151
R706 B.n376 B.n375 10.6151
R707 B.n375 B.n374 10.6151
R708 B.n374 B.n69 10.6151
R709 B.n370 B.n69 10.6151
R710 B.n370 B.n369 10.6151
R711 B.n369 B.n368 10.6151
R712 B.n368 B.n71 10.6151
R713 B.n364 B.n71 10.6151
R714 B.n364 B.n363 10.6151
R715 B.n363 B.n362 10.6151
R716 B.n362 B.n73 10.6151
R717 B.n358 B.n73 10.6151
R718 B.n358 B.n357 10.6151
R719 B.n357 B.n356 10.6151
R720 B.n356 B.n75 10.6151
R721 B.n352 B.n75 10.6151
R722 B.n352 B.n351 10.6151
R723 B.n351 B.n350 10.6151
R724 B.n350 B.n77 10.6151
R725 B.n346 B.n77 10.6151
R726 B.n346 B.n345 10.6151
R727 B.n345 B.n344 10.6151
R728 B.n344 B.n79 10.6151
R729 B.n340 B.n79 10.6151
R730 B.n340 B.n339 10.6151
R731 B.n339 B.n338 10.6151
R732 B.n338 B.n81 10.6151
R733 B.n334 B.n81 10.6151
R734 B.n334 B.n333 10.6151
R735 B.n333 B.n332 10.6151
R736 B.n332 B.n83 10.6151
R737 B.n328 B.n83 10.6151
R738 B.n145 B.n1 10.6151
R739 B.n148 B.n145 10.6151
R740 B.n149 B.n148 10.6151
R741 B.n150 B.n149 10.6151
R742 B.n150 B.n143 10.6151
R743 B.n154 B.n143 10.6151
R744 B.n155 B.n154 10.6151
R745 B.n156 B.n155 10.6151
R746 B.n156 B.n141 10.6151
R747 B.n160 B.n141 10.6151
R748 B.n161 B.n160 10.6151
R749 B.n162 B.n161 10.6151
R750 B.n162 B.n139 10.6151
R751 B.n166 B.n139 10.6151
R752 B.n167 B.n166 10.6151
R753 B.n168 B.n137 10.6151
R754 B.n172 B.n137 10.6151
R755 B.n173 B.n172 10.6151
R756 B.n174 B.n173 10.6151
R757 B.n174 B.n135 10.6151
R758 B.n178 B.n135 10.6151
R759 B.n179 B.n178 10.6151
R760 B.n180 B.n179 10.6151
R761 B.n180 B.n133 10.6151
R762 B.n184 B.n133 10.6151
R763 B.n185 B.n184 10.6151
R764 B.n186 B.n185 10.6151
R765 B.n186 B.n131 10.6151
R766 B.n190 B.n131 10.6151
R767 B.n191 B.n190 10.6151
R768 B.n192 B.n191 10.6151
R769 B.n192 B.n129 10.6151
R770 B.n196 B.n129 10.6151
R771 B.n197 B.n196 10.6151
R772 B.n198 B.n197 10.6151
R773 B.n198 B.n127 10.6151
R774 B.n202 B.n127 10.6151
R775 B.n203 B.n202 10.6151
R776 B.n204 B.n203 10.6151
R777 B.n204 B.n125 10.6151
R778 B.n208 B.n125 10.6151
R779 B.n209 B.n208 10.6151
R780 B.n210 B.n209 10.6151
R781 B.n210 B.n123 10.6151
R782 B.n214 B.n123 10.6151
R783 B.n215 B.n214 10.6151
R784 B.n216 B.n215 10.6151
R785 B.n216 B.n121 10.6151
R786 B.n220 B.n121 10.6151
R787 B.n221 B.n220 10.6151
R788 B.n222 B.n221 10.6151
R789 B.n222 B.n119 10.6151
R790 B.n226 B.n119 10.6151
R791 B.n227 B.n226 10.6151
R792 B.n228 B.n227 10.6151
R793 B.n228 B.n117 10.6151
R794 B.n232 B.n117 10.6151
R795 B.n233 B.n232 10.6151
R796 B.n234 B.n233 10.6151
R797 B.n234 B.n115 10.6151
R798 B.n238 B.n115 10.6151
R799 B.n241 B.n240 10.6151
R800 B.n241 B.n111 10.6151
R801 B.n245 B.n111 10.6151
R802 B.n246 B.n245 10.6151
R803 B.n247 B.n246 10.6151
R804 B.n247 B.n109 10.6151
R805 B.n251 B.n109 10.6151
R806 B.n252 B.n251 10.6151
R807 B.n256 B.n252 10.6151
R808 B.n260 B.n107 10.6151
R809 B.n261 B.n260 10.6151
R810 B.n262 B.n261 10.6151
R811 B.n262 B.n105 10.6151
R812 B.n266 B.n105 10.6151
R813 B.n267 B.n266 10.6151
R814 B.n268 B.n267 10.6151
R815 B.n268 B.n103 10.6151
R816 B.n272 B.n103 10.6151
R817 B.n273 B.n272 10.6151
R818 B.n274 B.n273 10.6151
R819 B.n274 B.n101 10.6151
R820 B.n278 B.n101 10.6151
R821 B.n279 B.n278 10.6151
R822 B.n280 B.n279 10.6151
R823 B.n280 B.n99 10.6151
R824 B.n284 B.n99 10.6151
R825 B.n285 B.n284 10.6151
R826 B.n286 B.n285 10.6151
R827 B.n286 B.n97 10.6151
R828 B.n290 B.n97 10.6151
R829 B.n291 B.n290 10.6151
R830 B.n292 B.n291 10.6151
R831 B.n292 B.n95 10.6151
R832 B.n296 B.n95 10.6151
R833 B.n297 B.n296 10.6151
R834 B.n298 B.n297 10.6151
R835 B.n298 B.n93 10.6151
R836 B.n302 B.n93 10.6151
R837 B.n303 B.n302 10.6151
R838 B.n304 B.n303 10.6151
R839 B.n304 B.n91 10.6151
R840 B.n308 B.n91 10.6151
R841 B.n309 B.n308 10.6151
R842 B.n310 B.n309 10.6151
R843 B.n310 B.n89 10.6151
R844 B.n314 B.n89 10.6151
R845 B.n315 B.n314 10.6151
R846 B.n316 B.n315 10.6151
R847 B.n316 B.n87 10.6151
R848 B.n320 B.n87 10.6151
R849 B.n321 B.n320 10.6151
R850 B.n322 B.n321 10.6151
R851 B.n322 B.n85 10.6151
R852 B.n326 B.n85 10.6151
R853 B.n327 B.n326 10.6151
R854 B.n466 B.n465 8.74196
R855 B.n448 B.n44 8.74196
R856 B.n239 B.n238 8.74196
R857 B.n255 B.n107 8.74196
R858 B.n561 B.n0 8.11757
R859 B.n561 B.n1 8.11757
R860 B.n465 B.n464 1.87367
R861 B.n44 B.n40 1.87367
R862 B.n240 B.n239 1.87367
R863 B.n256 B.n255 1.87367
R864 VP.n0 VP.t1 551.264
R865 VP.n0 VP.t0 509.286
R866 VP VP.n0 0.0516364
R867 VDD1 VDD1.t1 110.788
R868 VDD1 VDD1.t0 72.3352
C0 VDD1 VDD2 0.499821f
C1 VTAIL w_n1530_n3732# 3.14618f
C2 VTAIL VN 2.05795f
C3 B VP 1.1185f
C4 VDD1 VP 2.70658f
C5 B w_n1530_n3732# 7.66511f
C6 B VN 0.809647f
C7 VP VDD2 0.27029f
C8 VDD1 w_n1530_n3732# 1.74224f
C9 VDD1 VN 0.148424f
C10 w_n1530_n3732# VDD2 1.75061f
C11 VN VDD2 2.58905f
C12 B VTAIL 3.26569f
C13 VDD1 VTAIL 5.83414f
C14 VTAIL VDD2 5.87092f
C15 VP w_n1530_n3732# 2.1982f
C16 VN VP 5.0644f
C17 VN w_n1530_n3732# 2.0066f
C18 B VDD1 1.61423f
C19 VTAIL VP 2.07252f
C20 B VDD2 1.63139f
C21 VDD2 VSUBS 0.833122f
C22 VDD1 VSUBS 4.266845f
C23 VTAIL VSUBS 0.882527f
C24 VN VSUBS 7.90304f
C25 VP VSUBS 1.288925f
C26 B VSUBS 2.919746f
C27 w_n1530_n3732# VSUBS 70.1168f
C28 VDD1.t0 VSUBS 2.29135f
C29 VDD1.t1 VSUBS 2.87932f
C30 VP.t1 VSUBS 3.08875f
C31 VP.t0 VSUBS 2.84683f
C32 VP.n0 VSUBS 6.1296f
C33 B.n0 VSUBS 0.006055f
C34 B.n1 VSUBS 0.006055f
C35 B.n2 VSUBS 0.008954f
C36 B.n3 VSUBS 0.006862f
C37 B.n4 VSUBS 0.006862f
C38 B.n5 VSUBS 0.006862f
C39 B.n6 VSUBS 0.006862f
C40 B.n7 VSUBS 0.006862f
C41 B.n8 VSUBS 0.006862f
C42 B.n9 VSUBS 0.006862f
C43 B.n10 VSUBS 0.015146f
C44 B.n11 VSUBS 0.006862f
C45 B.n12 VSUBS 0.006862f
C46 B.n13 VSUBS 0.006862f
C47 B.n14 VSUBS 0.006862f
C48 B.n15 VSUBS 0.006862f
C49 B.n16 VSUBS 0.006862f
C50 B.n17 VSUBS 0.006862f
C51 B.n18 VSUBS 0.006862f
C52 B.n19 VSUBS 0.006862f
C53 B.n20 VSUBS 0.006862f
C54 B.n21 VSUBS 0.006862f
C55 B.n22 VSUBS 0.006862f
C56 B.n23 VSUBS 0.006862f
C57 B.n24 VSUBS 0.006862f
C58 B.n25 VSUBS 0.006862f
C59 B.n26 VSUBS 0.006862f
C60 B.n27 VSUBS 0.006862f
C61 B.n28 VSUBS 0.006862f
C62 B.n29 VSUBS 0.006862f
C63 B.n30 VSUBS 0.006862f
C64 B.n31 VSUBS 0.006862f
C65 B.n32 VSUBS 0.006862f
C66 B.n33 VSUBS 0.006862f
C67 B.t1 VSUBS 0.447042f
C68 B.t2 VSUBS 0.45778f
C69 B.t0 VSUBS 0.610572f
C70 B.n34 VSUBS 0.176761f
C71 B.n35 VSUBS 0.064271f
C72 B.n36 VSUBS 0.006862f
C73 B.n37 VSUBS 0.006862f
C74 B.n38 VSUBS 0.006862f
C75 B.n39 VSUBS 0.006862f
C76 B.n40 VSUBS 0.004036f
C77 B.n41 VSUBS 0.006862f
C78 B.t7 VSUBS 0.447031f
C79 B.t8 VSUBS 0.45777f
C80 B.t6 VSUBS 0.610572f
C81 B.n42 VSUBS 0.176771f
C82 B.n43 VSUBS 0.064282f
C83 B.n44 VSUBS 0.015898f
C84 B.n45 VSUBS 0.006862f
C85 B.n46 VSUBS 0.006862f
C86 B.n47 VSUBS 0.006862f
C87 B.n48 VSUBS 0.006862f
C88 B.n49 VSUBS 0.006862f
C89 B.n50 VSUBS 0.006862f
C90 B.n51 VSUBS 0.006862f
C91 B.n52 VSUBS 0.006862f
C92 B.n53 VSUBS 0.006862f
C93 B.n54 VSUBS 0.006862f
C94 B.n55 VSUBS 0.006862f
C95 B.n56 VSUBS 0.006862f
C96 B.n57 VSUBS 0.006862f
C97 B.n58 VSUBS 0.006862f
C98 B.n59 VSUBS 0.006862f
C99 B.n60 VSUBS 0.006862f
C100 B.n61 VSUBS 0.006862f
C101 B.n62 VSUBS 0.006862f
C102 B.n63 VSUBS 0.006862f
C103 B.n64 VSUBS 0.006862f
C104 B.n65 VSUBS 0.006862f
C105 B.n66 VSUBS 0.006862f
C106 B.n67 VSUBS 0.014118f
C107 B.n68 VSUBS 0.006862f
C108 B.n69 VSUBS 0.006862f
C109 B.n70 VSUBS 0.006862f
C110 B.n71 VSUBS 0.006862f
C111 B.n72 VSUBS 0.006862f
C112 B.n73 VSUBS 0.006862f
C113 B.n74 VSUBS 0.006862f
C114 B.n75 VSUBS 0.006862f
C115 B.n76 VSUBS 0.006862f
C116 B.n77 VSUBS 0.006862f
C117 B.n78 VSUBS 0.006862f
C118 B.n79 VSUBS 0.006862f
C119 B.n80 VSUBS 0.006862f
C120 B.n81 VSUBS 0.006862f
C121 B.n82 VSUBS 0.006862f
C122 B.n83 VSUBS 0.006862f
C123 B.n84 VSUBS 0.015146f
C124 B.n85 VSUBS 0.006862f
C125 B.n86 VSUBS 0.006862f
C126 B.n87 VSUBS 0.006862f
C127 B.n88 VSUBS 0.006862f
C128 B.n89 VSUBS 0.006862f
C129 B.n90 VSUBS 0.006862f
C130 B.n91 VSUBS 0.006862f
C131 B.n92 VSUBS 0.006862f
C132 B.n93 VSUBS 0.006862f
C133 B.n94 VSUBS 0.006862f
C134 B.n95 VSUBS 0.006862f
C135 B.n96 VSUBS 0.006862f
C136 B.n97 VSUBS 0.006862f
C137 B.n98 VSUBS 0.006862f
C138 B.n99 VSUBS 0.006862f
C139 B.n100 VSUBS 0.006862f
C140 B.n101 VSUBS 0.006862f
C141 B.n102 VSUBS 0.006862f
C142 B.n103 VSUBS 0.006862f
C143 B.n104 VSUBS 0.006862f
C144 B.n105 VSUBS 0.006862f
C145 B.n106 VSUBS 0.006862f
C146 B.n107 VSUBS 0.006256f
C147 B.n108 VSUBS 0.006862f
C148 B.n109 VSUBS 0.006862f
C149 B.n110 VSUBS 0.006862f
C150 B.n111 VSUBS 0.006862f
C151 B.n112 VSUBS 0.006862f
C152 B.t5 VSUBS 0.447042f
C153 B.t4 VSUBS 0.45778f
C154 B.t3 VSUBS 0.610572f
C155 B.n113 VSUBS 0.176761f
C156 B.n114 VSUBS 0.064271f
C157 B.n115 VSUBS 0.006862f
C158 B.n116 VSUBS 0.006862f
C159 B.n117 VSUBS 0.006862f
C160 B.n118 VSUBS 0.006862f
C161 B.n119 VSUBS 0.006862f
C162 B.n120 VSUBS 0.006862f
C163 B.n121 VSUBS 0.006862f
C164 B.n122 VSUBS 0.006862f
C165 B.n123 VSUBS 0.006862f
C166 B.n124 VSUBS 0.006862f
C167 B.n125 VSUBS 0.006862f
C168 B.n126 VSUBS 0.006862f
C169 B.n127 VSUBS 0.006862f
C170 B.n128 VSUBS 0.006862f
C171 B.n129 VSUBS 0.006862f
C172 B.n130 VSUBS 0.006862f
C173 B.n131 VSUBS 0.006862f
C174 B.n132 VSUBS 0.006862f
C175 B.n133 VSUBS 0.006862f
C176 B.n134 VSUBS 0.006862f
C177 B.n135 VSUBS 0.006862f
C178 B.n136 VSUBS 0.006862f
C179 B.n137 VSUBS 0.006862f
C180 B.n138 VSUBS 0.014118f
C181 B.n139 VSUBS 0.006862f
C182 B.n140 VSUBS 0.006862f
C183 B.n141 VSUBS 0.006862f
C184 B.n142 VSUBS 0.006862f
C185 B.n143 VSUBS 0.006862f
C186 B.n144 VSUBS 0.006862f
C187 B.n145 VSUBS 0.006862f
C188 B.n146 VSUBS 0.006862f
C189 B.n147 VSUBS 0.006862f
C190 B.n148 VSUBS 0.006862f
C191 B.n149 VSUBS 0.006862f
C192 B.n150 VSUBS 0.006862f
C193 B.n151 VSUBS 0.006862f
C194 B.n152 VSUBS 0.006862f
C195 B.n153 VSUBS 0.006862f
C196 B.n154 VSUBS 0.006862f
C197 B.n155 VSUBS 0.006862f
C198 B.n156 VSUBS 0.006862f
C199 B.n157 VSUBS 0.006862f
C200 B.n158 VSUBS 0.006862f
C201 B.n159 VSUBS 0.006862f
C202 B.n160 VSUBS 0.006862f
C203 B.n161 VSUBS 0.006862f
C204 B.n162 VSUBS 0.006862f
C205 B.n163 VSUBS 0.006862f
C206 B.n164 VSUBS 0.006862f
C207 B.n165 VSUBS 0.006862f
C208 B.n166 VSUBS 0.006862f
C209 B.n167 VSUBS 0.014118f
C210 B.n168 VSUBS 0.015146f
C211 B.n169 VSUBS 0.015146f
C212 B.n170 VSUBS 0.006862f
C213 B.n171 VSUBS 0.006862f
C214 B.n172 VSUBS 0.006862f
C215 B.n173 VSUBS 0.006862f
C216 B.n174 VSUBS 0.006862f
C217 B.n175 VSUBS 0.006862f
C218 B.n176 VSUBS 0.006862f
C219 B.n177 VSUBS 0.006862f
C220 B.n178 VSUBS 0.006862f
C221 B.n179 VSUBS 0.006862f
C222 B.n180 VSUBS 0.006862f
C223 B.n181 VSUBS 0.006862f
C224 B.n182 VSUBS 0.006862f
C225 B.n183 VSUBS 0.006862f
C226 B.n184 VSUBS 0.006862f
C227 B.n185 VSUBS 0.006862f
C228 B.n186 VSUBS 0.006862f
C229 B.n187 VSUBS 0.006862f
C230 B.n188 VSUBS 0.006862f
C231 B.n189 VSUBS 0.006862f
C232 B.n190 VSUBS 0.006862f
C233 B.n191 VSUBS 0.006862f
C234 B.n192 VSUBS 0.006862f
C235 B.n193 VSUBS 0.006862f
C236 B.n194 VSUBS 0.006862f
C237 B.n195 VSUBS 0.006862f
C238 B.n196 VSUBS 0.006862f
C239 B.n197 VSUBS 0.006862f
C240 B.n198 VSUBS 0.006862f
C241 B.n199 VSUBS 0.006862f
C242 B.n200 VSUBS 0.006862f
C243 B.n201 VSUBS 0.006862f
C244 B.n202 VSUBS 0.006862f
C245 B.n203 VSUBS 0.006862f
C246 B.n204 VSUBS 0.006862f
C247 B.n205 VSUBS 0.006862f
C248 B.n206 VSUBS 0.006862f
C249 B.n207 VSUBS 0.006862f
C250 B.n208 VSUBS 0.006862f
C251 B.n209 VSUBS 0.006862f
C252 B.n210 VSUBS 0.006862f
C253 B.n211 VSUBS 0.006862f
C254 B.n212 VSUBS 0.006862f
C255 B.n213 VSUBS 0.006862f
C256 B.n214 VSUBS 0.006862f
C257 B.n215 VSUBS 0.006862f
C258 B.n216 VSUBS 0.006862f
C259 B.n217 VSUBS 0.006862f
C260 B.n218 VSUBS 0.006862f
C261 B.n219 VSUBS 0.006862f
C262 B.n220 VSUBS 0.006862f
C263 B.n221 VSUBS 0.006862f
C264 B.n222 VSUBS 0.006862f
C265 B.n223 VSUBS 0.006862f
C266 B.n224 VSUBS 0.006862f
C267 B.n225 VSUBS 0.006862f
C268 B.n226 VSUBS 0.006862f
C269 B.n227 VSUBS 0.006862f
C270 B.n228 VSUBS 0.006862f
C271 B.n229 VSUBS 0.006862f
C272 B.n230 VSUBS 0.006862f
C273 B.n231 VSUBS 0.006862f
C274 B.n232 VSUBS 0.006862f
C275 B.n233 VSUBS 0.006862f
C276 B.n234 VSUBS 0.006862f
C277 B.n235 VSUBS 0.006862f
C278 B.n236 VSUBS 0.006862f
C279 B.n237 VSUBS 0.006862f
C280 B.n238 VSUBS 0.006256f
C281 B.n239 VSUBS 0.015898f
C282 B.n240 VSUBS 0.004036f
C283 B.n241 VSUBS 0.006862f
C284 B.n242 VSUBS 0.006862f
C285 B.n243 VSUBS 0.006862f
C286 B.n244 VSUBS 0.006862f
C287 B.n245 VSUBS 0.006862f
C288 B.n246 VSUBS 0.006862f
C289 B.n247 VSUBS 0.006862f
C290 B.n248 VSUBS 0.006862f
C291 B.n249 VSUBS 0.006862f
C292 B.n250 VSUBS 0.006862f
C293 B.n251 VSUBS 0.006862f
C294 B.n252 VSUBS 0.006862f
C295 B.t11 VSUBS 0.447031f
C296 B.t10 VSUBS 0.45777f
C297 B.t9 VSUBS 0.610572f
C298 B.n253 VSUBS 0.176771f
C299 B.n254 VSUBS 0.064282f
C300 B.n255 VSUBS 0.015898f
C301 B.n256 VSUBS 0.004036f
C302 B.n257 VSUBS 0.006862f
C303 B.n258 VSUBS 0.006862f
C304 B.n259 VSUBS 0.006862f
C305 B.n260 VSUBS 0.006862f
C306 B.n261 VSUBS 0.006862f
C307 B.n262 VSUBS 0.006862f
C308 B.n263 VSUBS 0.006862f
C309 B.n264 VSUBS 0.006862f
C310 B.n265 VSUBS 0.006862f
C311 B.n266 VSUBS 0.006862f
C312 B.n267 VSUBS 0.006862f
C313 B.n268 VSUBS 0.006862f
C314 B.n269 VSUBS 0.006862f
C315 B.n270 VSUBS 0.006862f
C316 B.n271 VSUBS 0.006862f
C317 B.n272 VSUBS 0.006862f
C318 B.n273 VSUBS 0.006862f
C319 B.n274 VSUBS 0.006862f
C320 B.n275 VSUBS 0.006862f
C321 B.n276 VSUBS 0.006862f
C322 B.n277 VSUBS 0.006862f
C323 B.n278 VSUBS 0.006862f
C324 B.n279 VSUBS 0.006862f
C325 B.n280 VSUBS 0.006862f
C326 B.n281 VSUBS 0.006862f
C327 B.n282 VSUBS 0.006862f
C328 B.n283 VSUBS 0.006862f
C329 B.n284 VSUBS 0.006862f
C330 B.n285 VSUBS 0.006862f
C331 B.n286 VSUBS 0.006862f
C332 B.n287 VSUBS 0.006862f
C333 B.n288 VSUBS 0.006862f
C334 B.n289 VSUBS 0.006862f
C335 B.n290 VSUBS 0.006862f
C336 B.n291 VSUBS 0.006862f
C337 B.n292 VSUBS 0.006862f
C338 B.n293 VSUBS 0.006862f
C339 B.n294 VSUBS 0.006862f
C340 B.n295 VSUBS 0.006862f
C341 B.n296 VSUBS 0.006862f
C342 B.n297 VSUBS 0.006862f
C343 B.n298 VSUBS 0.006862f
C344 B.n299 VSUBS 0.006862f
C345 B.n300 VSUBS 0.006862f
C346 B.n301 VSUBS 0.006862f
C347 B.n302 VSUBS 0.006862f
C348 B.n303 VSUBS 0.006862f
C349 B.n304 VSUBS 0.006862f
C350 B.n305 VSUBS 0.006862f
C351 B.n306 VSUBS 0.006862f
C352 B.n307 VSUBS 0.006862f
C353 B.n308 VSUBS 0.006862f
C354 B.n309 VSUBS 0.006862f
C355 B.n310 VSUBS 0.006862f
C356 B.n311 VSUBS 0.006862f
C357 B.n312 VSUBS 0.006862f
C358 B.n313 VSUBS 0.006862f
C359 B.n314 VSUBS 0.006862f
C360 B.n315 VSUBS 0.006862f
C361 B.n316 VSUBS 0.006862f
C362 B.n317 VSUBS 0.006862f
C363 B.n318 VSUBS 0.006862f
C364 B.n319 VSUBS 0.006862f
C365 B.n320 VSUBS 0.006862f
C366 B.n321 VSUBS 0.006862f
C367 B.n322 VSUBS 0.006862f
C368 B.n323 VSUBS 0.006862f
C369 B.n324 VSUBS 0.006862f
C370 B.n325 VSUBS 0.006862f
C371 B.n326 VSUBS 0.006862f
C372 B.n327 VSUBS 0.014209f
C373 B.n328 VSUBS 0.015055f
C374 B.n329 VSUBS 0.014118f
C375 B.n330 VSUBS 0.006862f
C376 B.n331 VSUBS 0.006862f
C377 B.n332 VSUBS 0.006862f
C378 B.n333 VSUBS 0.006862f
C379 B.n334 VSUBS 0.006862f
C380 B.n335 VSUBS 0.006862f
C381 B.n336 VSUBS 0.006862f
C382 B.n337 VSUBS 0.006862f
C383 B.n338 VSUBS 0.006862f
C384 B.n339 VSUBS 0.006862f
C385 B.n340 VSUBS 0.006862f
C386 B.n341 VSUBS 0.006862f
C387 B.n342 VSUBS 0.006862f
C388 B.n343 VSUBS 0.006862f
C389 B.n344 VSUBS 0.006862f
C390 B.n345 VSUBS 0.006862f
C391 B.n346 VSUBS 0.006862f
C392 B.n347 VSUBS 0.006862f
C393 B.n348 VSUBS 0.006862f
C394 B.n349 VSUBS 0.006862f
C395 B.n350 VSUBS 0.006862f
C396 B.n351 VSUBS 0.006862f
C397 B.n352 VSUBS 0.006862f
C398 B.n353 VSUBS 0.006862f
C399 B.n354 VSUBS 0.006862f
C400 B.n355 VSUBS 0.006862f
C401 B.n356 VSUBS 0.006862f
C402 B.n357 VSUBS 0.006862f
C403 B.n358 VSUBS 0.006862f
C404 B.n359 VSUBS 0.006862f
C405 B.n360 VSUBS 0.006862f
C406 B.n361 VSUBS 0.006862f
C407 B.n362 VSUBS 0.006862f
C408 B.n363 VSUBS 0.006862f
C409 B.n364 VSUBS 0.006862f
C410 B.n365 VSUBS 0.006862f
C411 B.n366 VSUBS 0.006862f
C412 B.n367 VSUBS 0.006862f
C413 B.n368 VSUBS 0.006862f
C414 B.n369 VSUBS 0.006862f
C415 B.n370 VSUBS 0.006862f
C416 B.n371 VSUBS 0.006862f
C417 B.n372 VSUBS 0.006862f
C418 B.n373 VSUBS 0.006862f
C419 B.n374 VSUBS 0.006862f
C420 B.n375 VSUBS 0.006862f
C421 B.n376 VSUBS 0.006862f
C422 B.n377 VSUBS 0.006862f
C423 B.n378 VSUBS 0.014118f
C424 B.n379 VSUBS 0.015146f
C425 B.n380 VSUBS 0.015146f
C426 B.n381 VSUBS 0.006862f
C427 B.n382 VSUBS 0.006862f
C428 B.n383 VSUBS 0.006862f
C429 B.n384 VSUBS 0.006862f
C430 B.n385 VSUBS 0.006862f
C431 B.n386 VSUBS 0.006862f
C432 B.n387 VSUBS 0.006862f
C433 B.n388 VSUBS 0.006862f
C434 B.n389 VSUBS 0.006862f
C435 B.n390 VSUBS 0.006862f
C436 B.n391 VSUBS 0.006862f
C437 B.n392 VSUBS 0.006862f
C438 B.n393 VSUBS 0.006862f
C439 B.n394 VSUBS 0.006862f
C440 B.n395 VSUBS 0.006862f
C441 B.n396 VSUBS 0.006862f
C442 B.n397 VSUBS 0.006862f
C443 B.n398 VSUBS 0.006862f
C444 B.n399 VSUBS 0.006862f
C445 B.n400 VSUBS 0.006862f
C446 B.n401 VSUBS 0.006862f
C447 B.n402 VSUBS 0.006862f
C448 B.n403 VSUBS 0.006862f
C449 B.n404 VSUBS 0.006862f
C450 B.n405 VSUBS 0.006862f
C451 B.n406 VSUBS 0.006862f
C452 B.n407 VSUBS 0.006862f
C453 B.n408 VSUBS 0.006862f
C454 B.n409 VSUBS 0.006862f
C455 B.n410 VSUBS 0.006862f
C456 B.n411 VSUBS 0.006862f
C457 B.n412 VSUBS 0.006862f
C458 B.n413 VSUBS 0.006862f
C459 B.n414 VSUBS 0.006862f
C460 B.n415 VSUBS 0.006862f
C461 B.n416 VSUBS 0.006862f
C462 B.n417 VSUBS 0.006862f
C463 B.n418 VSUBS 0.006862f
C464 B.n419 VSUBS 0.006862f
C465 B.n420 VSUBS 0.006862f
C466 B.n421 VSUBS 0.006862f
C467 B.n422 VSUBS 0.006862f
C468 B.n423 VSUBS 0.006862f
C469 B.n424 VSUBS 0.006862f
C470 B.n425 VSUBS 0.006862f
C471 B.n426 VSUBS 0.006862f
C472 B.n427 VSUBS 0.006862f
C473 B.n428 VSUBS 0.006862f
C474 B.n429 VSUBS 0.006862f
C475 B.n430 VSUBS 0.006862f
C476 B.n431 VSUBS 0.006862f
C477 B.n432 VSUBS 0.006862f
C478 B.n433 VSUBS 0.006862f
C479 B.n434 VSUBS 0.006862f
C480 B.n435 VSUBS 0.006862f
C481 B.n436 VSUBS 0.006862f
C482 B.n437 VSUBS 0.006862f
C483 B.n438 VSUBS 0.006862f
C484 B.n439 VSUBS 0.006862f
C485 B.n440 VSUBS 0.006862f
C486 B.n441 VSUBS 0.006862f
C487 B.n442 VSUBS 0.006862f
C488 B.n443 VSUBS 0.006862f
C489 B.n444 VSUBS 0.006862f
C490 B.n445 VSUBS 0.006862f
C491 B.n446 VSUBS 0.006862f
C492 B.n447 VSUBS 0.006862f
C493 B.n448 VSUBS 0.006256f
C494 B.n449 VSUBS 0.006862f
C495 B.n450 VSUBS 0.006862f
C496 B.n451 VSUBS 0.006862f
C497 B.n452 VSUBS 0.006862f
C498 B.n453 VSUBS 0.006862f
C499 B.n454 VSUBS 0.006862f
C500 B.n455 VSUBS 0.006862f
C501 B.n456 VSUBS 0.006862f
C502 B.n457 VSUBS 0.006862f
C503 B.n458 VSUBS 0.006862f
C504 B.n459 VSUBS 0.006862f
C505 B.n460 VSUBS 0.006862f
C506 B.n461 VSUBS 0.006862f
C507 B.n462 VSUBS 0.006862f
C508 B.n463 VSUBS 0.006862f
C509 B.n464 VSUBS 0.004036f
C510 B.n465 VSUBS 0.015898f
C511 B.n466 VSUBS 0.006256f
C512 B.n467 VSUBS 0.006862f
C513 B.n468 VSUBS 0.006862f
C514 B.n469 VSUBS 0.006862f
C515 B.n470 VSUBS 0.006862f
C516 B.n471 VSUBS 0.006862f
C517 B.n472 VSUBS 0.006862f
C518 B.n473 VSUBS 0.006862f
C519 B.n474 VSUBS 0.006862f
C520 B.n475 VSUBS 0.006862f
C521 B.n476 VSUBS 0.006862f
C522 B.n477 VSUBS 0.006862f
C523 B.n478 VSUBS 0.006862f
C524 B.n479 VSUBS 0.006862f
C525 B.n480 VSUBS 0.006862f
C526 B.n481 VSUBS 0.006862f
C527 B.n482 VSUBS 0.006862f
C528 B.n483 VSUBS 0.006862f
C529 B.n484 VSUBS 0.006862f
C530 B.n485 VSUBS 0.006862f
C531 B.n486 VSUBS 0.006862f
C532 B.n487 VSUBS 0.006862f
C533 B.n488 VSUBS 0.006862f
C534 B.n489 VSUBS 0.006862f
C535 B.n490 VSUBS 0.006862f
C536 B.n491 VSUBS 0.006862f
C537 B.n492 VSUBS 0.006862f
C538 B.n493 VSUBS 0.006862f
C539 B.n494 VSUBS 0.006862f
C540 B.n495 VSUBS 0.006862f
C541 B.n496 VSUBS 0.006862f
C542 B.n497 VSUBS 0.006862f
C543 B.n498 VSUBS 0.006862f
C544 B.n499 VSUBS 0.006862f
C545 B.n500 VSUBS 0.006862f
C546 B.n501 VSUBS 0.006862f
C547 B.n502 VSUBS 0.006862f
C548 B.n503 VSUBS 0.006862f
C549 B.n504 VSUBS 0.006862f
C550 B.n505 VSUBS 0.006862f
C551 B.n506 VSUBS 0.006862f
C552 B.n507 VSUBS 0.006862f
C553 B.n508 VSUBS 0.006862f
C554 B.n509 VSUBS 0.006862f
C555 B.n510 VSUBS 0.006862f
C556 B.n511 VSUBS 0.006862f
C557 B.n512 VSUBS 0.006862f
C558 B.n513 VSUBS 0.006862f
C559 B.n514 VSUBS 0.006862f
C560 B.n515 VSUBS 0.006862f
C561 B.n516 VSUBS 0.006862f
C562 B.n517 VSUBS 0.006862f
C563 B.n518 VSUBS 0.006862f
C564 B.n519 VSUBS 0.006862f
C565 B.n520 VSUBS 0.006862f
C566 B.n521 VSUBS 0.006862f
C567 B.n522 VSUBS 0.006862f
C568 B.n523 VSUBS 0.006862f
C569 B.n524 VSUBS 0.006862f
C570 B.n525 VSUBS 0.006862f
C571 B.n526 VSUBS 0.006862f
C572 B.n527 VSUBS 0.006862f
C573 B.n528 VSUBS 0.006862f
C574 B.n529 VSUBS 0.006862f
C575 B.n530 VSUBS 0.006862f
C576 B.n531 VSUBS 0.006862f
C577 B.n532 VSUBS 0.006862f
C578 B.n533 VSUBS 0.006862f
C579 B.n534 VSUBS 0.006862f
C580 B.n535 VSUBS 0.015146f
C581 B.n536 VSUBS 0.014118f
C582 B.n537 VSUBS 0.014118f
C583 B.n538 VSUBS 0.006862f
C584 B.n539 VSUBS 0.006862f
C585 B.n540 VSUBS 0.006862f
C586 B.n541 VSUBS 0.006862f
C587 B.n542 VSUBS 0.006862f
C588 B.n543 VSUBS 0.006862f
C589 B.n544 VSUBS 0.006862f
C590 B.n545 VSUBS 0.006862f
C591 B.n546 VSUBS 0.006862f
C592 B.n547 VSUBS 0.006862f
C593 B.n548 VSUBS 0.006862f
C594 B.n549 VSUBS 0.006862f
C595 B.n550 VSUBS 0.006862f
C596 B.n551 VSUBS 0.006862f
C597 B.n552 VSUBS 0.006862f
C598 B.n553 VSUBS 0.006862f
C599 B.n554 VSUBS 0.006862f
C600 B.n555 VSUBS 0.006862f
C601 B.n556 VSUBS 0.006862f
C602 B.n557 VSUBS 0.006862f
C603 B.n558 VSUBS 0.006862f
C604 B.n559 VSUBS 0.008954f
C605 B.n560 VSUBS 0.009539f
C606 B.n561 VSUBS 0.018969f
C607 VDD2.t1 VSUBS 2.87774f
C608 VDD2.t0 VSUBS 2.3092f
C609 VDD2.n0 VSUBS 3.24901f
C610 VTAIL.t0 VSUBS 3.01569f
C611 VTAIL.n0 VSUBS 2.5923f
C612 VTAIL.t2 VSUBS 3.01571f
C613 VTAIL.n1 VSUBS 2.61461f
C614 VTAIL.t1 VSUBS 3.01571f
C615 VTAIL.n2 VSUBS 2.50397f
C616 VTAIL.t3 VSUBS 3.01569f
C617 VTAIL.n3 VSUBS 2.42792f
C618 VN.t0 VSUBS 2.75697f
C619 VN.t1 VSUBS 2.9961f
.ends

