* NGSPICE file created from diff_pair_sample_0827.ext - technology: sky130A

.subckt diff_pair_sample_0827 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=1.54935 pd=9.72 as=1.54935 ps=9.72 w=9.39 l=2.88
X1 VTAIL.t1 VN.t0 VDD2.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=3.6621 pd=19.56 as=1.54935 ps=9.72 w=9.39 l=2.88
X2 VDD2.t6 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.54935 pd=9.72 as=1.54935 ps=9.72 w=9.39 l=2.88
X3 VTAIL.t8 VP.t1 VDD1.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=3.6621 pd=19.56 as=1.54935 ps=9.72 w=9.39 l=2.88
X4 VDD1.t5 VP.t2 VTAIL.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=1.54935 pd=9.72 as=3.6621 ps=19.56 w=9.39 l=2.88
X5 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=3.6621 pd=19.56 as=0 ps=0 w=9.39 l=2.88
X6 VTAIL.t0 VN.t2 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.54935 pd=9.72 as=1.54935 ps=9.72 w=9.39 l=2.88
X7 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=3.6621 pd=19.56 as=0 ps=0 w=9.39 l=2.88
X8 VTAIL.t10 VP.t3 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.54935 pd=9.72 as=1.54935 ps=9.72 w=9.39 l=2.88
X9 VDD1.t3 VP.t4 VTAIL.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=1.54935 pd=9.72 as=1.54935 ps=9.72 w=9.39 l=2.88
X10 VTAIL.t6 VN.t3 VDD2.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=3.6621 pd=19.56 as=1.54935 ps=9.72 w=9.39 l=2.88
X11 VDD1.t2 VP.t5 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=1.54935 pd=9.72 as=3.6621 ps=19.56 w=9.39 l=2.88
X12 VTAIL.t13 VP.t6 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.54935 pd=9.72 as=1.54935 ps=9.72 w=9.39 l=2.88
X13 VTAIL.t7 VP.t7 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=3.6621 pd=19.56 as=1.54935 ps=9.72 w=9.39 l=2.88
X14 VDD2.t3 VN.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.54935 pd=9.72 as=3.6621 ps=19.56 w=9.39 l=2.88
X15 VDD2.t2 VN.t5 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=1.54935 pd=9.72 as=3.6621 ps=19.56 w=9.39 l=2.88
X16 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=3.6621 pd=19.56 as=0 ps=0 w=9.39 l=2.88
X17 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.6621 pd=19.56 as=0 ps=0 w=9.39 l=2.88
X18 VTAIL.t2 VN.t6 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.54935 pd=9.72 as=1.54935 ps=9.72 w=9.39 l=2.88
X19 VDD2.t0 VN.t7 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.54935 pd=9.72 as=1.54935 ps=9.72 w=9.39 l=2.88
R0 VP.n19 VP.n16 161.3
R1 VP.n21 VP.n20 161.3
R2 VP.n22 VP.n15 161.3
R3 VP.n24 VP.n23 161.3
R4 VP.n25 VP.n14 161.3
R5 VP.n28 VP.n27 161.3
R6 VP.n29 VP.n13 161.3
R7 VP.n31 VP.n30 161.3
R8 VP.n32 VP.n12 161.3
R9 VP.n34 VP.n33 161.3
R10 VP.n35 VP.n11 161.3
R11 VP.n37 VP.n36 161.3
R12 VP.n38 VP.n10 161.3
R13 VP.n74 VP.n0 161.3
R14 VP.n73 VP.n72 161.3
R15 VP.n71 VP.n1 161.3
R16 VP.n70 VP.n69 161.3
R17 VP.n68 VP.n2 161.3
R18 VP.n67 VP.n66 161.3
R19 VP.n65 VP.n3 161.3
R20 VP.n64 VP.n63 161.3
R21 VP.n61 VP.n4 161.3
R22 VP.n60 VP.n59 161.3
R23 VP.n58 VP.n5 161.3
R24 VP.n57 VP.n56 161.3
R25 VP.n55 VP.n6 161.3
R26 VP.n53 VP.n52 161.3
R27 VP.n51 VP.n7 161.3
R28 VP.n50 VP.n49 161.3
R29 VP.n48 VP.n8 161.3
R30 VP.n47 VP.n46 161.3
R31 VP.n45 VP.n9 161.3
R32 VP.n44 VP.n43 161.3
R33 VP.n17 VP.t7 111.825
R34 VP.n42 VP.n41 107.576
R35 VP.n76 VP.n75 107.576
R36 VP.n40 VP.n39 107.576
R37 VP.n42 VP.t1 78.5765
R38 VP.n54 VP.t4 78.5765
R39 VP.n62 VP.t3 78.5765
R40 VP.n75 VP.t5 78.5765
R41 VP.n39 VP.t2 78.5765
R42 VP.n26 VP.t6 78.5765
R43 VP.n18 VP.t0 78.5765
R44 VP.n60 VP.n5 56.5193
R45 VP.n24 VP.n15 56.5193
R46 VP.n18 VP.n17 56.3164
R47 VP.n41 VP.n40 50.2117
R48 VP.n49 VP.n48 44.3785
R49 VP.n69 VP.n68 44.3785
R50 VP.n33 VP.n32 44.3785
R51 VP.n48 VP.n47 36.6083
R52 VP.n69 VP.n1 36.6083
R53 VP.n33 VP.n11 36.6083
R54 VP.n43 VP.n9 24.4675
R55 VP.n47 VP.n9 24.4675
R56 VP.n49 VP.n7 24.4675
R57 VP.n53 VP.n7 24.4675
R58 VP.n56 VP.n55 24.4675
R59 VP.n56 VP.n5 24.4675
R60 VP.n61 VP.n60 24.4675
R61 VP.n63 VP.n61 24.4675
R62 VP.n67 VP.n3 24.4675
R63 VP.n68 VP.n67 24.4675
R64 VP.n73 VP.n1 24.4675
R65 VP.n74 VP.n73 24.4675
R66 VP.n37 VP.n11 24.4675
R67 VP.n38 VP.n37 24.4675
R68 VP.n25 VP.n24 24.4675
R69 VP.n27 VP.n25 24.4675
R70 VP.n31 VP.n13 24.4675
R71 VP.n32 VP.n31 24.4675
R72 VP.n20 VP.n19 24.4675
R73 VP.n20 VP.n15 24.4675
R74 VP.n55 VP.n54 17.3721
R75 VP.n63 VP.n62 17.3721
R76 VP.n27 VP.n26 17.3721
R77 VP.n19 VP.n18 17.3721
R78 VP.n54 VP.n53 7.09593
R79 VP.n62 VP.n3 7.09593
R80 VP.n26 VP.n13 7.09593
R81 VP.n17 VP.n16 5.06027
R82 VP.n43 VP.n42 3.18121
R83 VP.n75 VP.n74 3.18121
R84 VP.n39 VP.n38 3.18121
R85 VP.n40 VP.n10 0.278367
R86 VP.n44 VP.n41 0.278367
R87 VP.n76 VP.n0 0.278367
R88 VP.n21 VP.n16 0.189894
R89 VP.n22 VP.n21 0.189894
R90 VP.n23 VP.n22 0.189894
R91 VP.n23 VP.n14 0.189894
R92 VP.n28 VP.n14 0.189894
R93 VP.n29 VP.n28 0.189894
R94 VP.n30 VP.n29 0.189894
R95 VP.n30 VP.n12 0.189894
R96 VP.n34 VP.n12 0.189894
R97 VP.n35 VP.n34 0.189894
R98 VP.n36 VP.n35 0.189894
R99 VP.n36 VP.n10 0.189894
R100 VP.n45 VP.n44 0.189894
R101 VP.n46 VP.n45 0.189894
R102 VP.n46 VP.n8 0.189894
R103 VP.n50 VP.n8 0.189894
R104 VP.n51 VP.n50 0.189894
R105 VP.n52 VP.n51 0.189894
R106 VP.n52 VP.n6 0.189894
R107 VP.n57 VP.n6 0.189894
R108 VP.n58 VP.n57 0.189894
R109 VP.n59 VP.n58 0.189894
R110 VP.n59 VP.n4 0.189894
R111 VP.n64 VP.n4 0.189894
R112 VP.n65 VP.n64 0.189894
R113 VP.n66 VP.n65 0.189894
R114 VP.n66 VP.n2 0.189894
R115 VP.n70 VP.n2 0.189894
R116 VP.n71 VP.n70 0.189894
R117 VP.n72 VP.n71 0.189894
R118 VP.n72 VP.n0 0.189894
R119 VP VP.n76 0.153454
R120 VTAIL.n402 VTAIL.n358 289.615
R121 VTAIL.n46 VTAIL.n2 289.615
R122 VTAIL.n96 VTAIL.n52 289.615
R123 VTAIL.n148 VTAIL.n104 289.615
R124 VTAIL.n352 VTAIL.n308 289.615
R125 VTAIL.n300 VTAIL.n256 289.615
R126 VTAIL.n250 VTAIL.n206 289.615
R127 VTAIL.n198 VTAIL.n154 289.615
R128 VTAIL.n375 VTAIL.n374 185
R129 VTAIL.n377 VTAIL.n376 185
R130 VTAIL.n370 VTAIL.n369 185
R131 VTAIL.n383 VTAIL.n382 185
R132 VTAIL.n385 VTAIL.n384 185
R133 VTAIL.n366 VTAIL.n365 185
R134 VTAIL.n392 VTAIL.n391 185
R135 VTAIL.n393 VTAIL.n364 185
R136 VTAIL.n395 VTAIL.n394 185
R137 VTAIL.n362 VTAIL.n361 185
R138 VTAIL.n401 VTAIL.n400 185
R139 VTAIL.n403 VTAIL.n402 185
R140 VTAIL.n19 VTAIL.n18 185
R141 VTAIL.n21 VTAIL.n20 185
R142 VTAIL.n14 VTAIL.n13 185
R143 VTAIL.n27 VTAIL.n26 185
R144 VTAIL.n29 VTAIL.n28 185
R145 VTAIL.n10 VTAIL.n9 185
R146 VTAIL.n36 VTAIL.n35 185
R147 VTAIL.n37 VTAIL.n8 185
R148 VTAIL.n39 VTAIL.n38 185
R149 VTAIL.n6 VTAIL.n5 185
R150 VTAIL.n45 VTAIL.n44 185
R151 VTAIL.n47 VTAIL.n46 185
R152 VTAIL.n69 VTAIL.n68 185
R153 VTAIL.n71 VTAIL.n70 185
R154 VTAIL.n64 VTAIL.n63 185
R155 VTAIL.n77 VTAIL.n76 185
R156 VTAIL.n79 VTAIL.n78 185
R157 VTAIL.n60 VTAIL.n59 185
R158 VTAIL.n86 VTAIL.n85 185
R159 VTAIL.n87 VTAIL.n58 185
R160 VTAIL.n89 VTAIL.n88 185
R161 VTAIL.n56 VTAIL.n55 185
R162 VTAIL.n95 VTAIL.n94 185
R163 VTAIL.n97 VTAIL.n96 185
R164 VTAIL.n121 VTAIL.n120 185
R165 VTAIL.n123 VTAIL.n122 185
R166 VTAIL.n116 VTAIL.n115 185
R167 VTAIL.n129 VTAIL.n128 185
R168 VTAIL.n131 VTAIL.n130 185
R169 VTAIL.n112 VTAIL.n111 185
R170 VTAIL.n138 VTAIL.n137 185
R171 VTAIL.n139 VTAIL.n110 185
R172 VTAIL.n141 VTAIL.n140 185
R173 VTAIL.n108 VTAIL.n107 185
R174 VTAIL.n147 VTAIL.n146 185
R175 VTAIL.n149 VTAIL.n148 185
R176 VTAIL.n353 VTAIL.n352 185
R177 VTAIL.n351 VTAIL.n350 185
R178 VTAIL.n312 VTAIL.n311 185
R179 VTAIL.n316 VTAIL.n314 185
R180 VTAIL.n345 VTAIL.n344 185
R181 VTAIL.n343 VTAIL.n342 185
R182 VTAIL.n318 VTAIL.n317 185
R183 VTAIL.n337 VTAIL.n336 185
R184 VTAIL.n335 VTAIL.n334 185
R185 VTAIL.n322 VTAIL.n321 185
R186 VTAIL.n329 VTAIL.n328 185
R187 VTAIL.n327 VTAIL.n326 185
R188 VTAIL.n301 VTAIL.n300 185
R189 VTAIL.n299 VTAIL.n298 185
R190 VTAIL.n260 VTAIL.n259 185
R191 VTAIL.n264 VTAIL.n262 185
R192 VTAIL.n293 VTAIL.n292 185
R193 VTAIL.n291 VTAIL.n290 185
R194 VTAIL.n266 VTAIL.n265 185
R195 VTAIL.n285 VTAIL.n284 185
R196 VTAIL.n283 VTAIL.n282 185
R197 VTAIL.n270 VTAIL.n269 185
R198 VTAIL.n277 VTAIL.n276 185
R199 VTAIL.n275 VTAIL.n274 185
R200 VTAIL.n251 VTAIL.n250 185
R201 VTAIL.n249 VTAIL.n248 185
R202 VTAIL.n210 VTAIL.n209 185
R203 VTAIL.n214 VTAIL.n212 185
R204 VTAIL.n243 VTAIL.n242 185
R205 VTAIL.n241 VTAIL.n240 185
R206 VTAIL.n216 VTAIL.n215 185
R207 VTAIL.n235 VTAIL.n234 185
R208 VTAIL.n233 VTAIL.n232 185
R209 VTAIL.n220 VTAIL.n219 185
R210 VTAIL.n227 VTAIL.n226 185
R211 VTAIL.n225 VTAIL.n224 185
R212 VTAIL.n199 VTAIL.n198 185
R213 VTAIL.n197 VTAIL.n196 185
R214 VTAIL.n158 VTAIL.n157 185
R215 VTAIL.n162 VTAIL.n160 185
R216 VTAIL.n191 VTAIL.n190 185
R217 VTAIL.n189 VTAIL.n188 185
R218 VTAIL.n164 VTAIL.n163 185
R219 VTAIL.n183 VTAIL.n182 185
R220 VTAIL.n181 VTAIL.n180 185
R221 VTAIL.n168 VTAIL.n167 185
R222 VTAIL.n175 VTAIL.n174 185
R223 VTAIL.n173 VTAIL.n172 185
R224 VTAIL.n373 VTAIL.t15 149.524
R225 VTAIL.n17 VTAIL.t1 149.524
R226 VTAIL.n67 VTAIL.t12 149.524
R227 VTAIL.n119 VTAIL.t8 149.524
R228 VTAIL.n325 VTAIL.t9 149.524
R229 VTAIL.n273 VTAIL.t7 149.524
R230 VTAIL.n223 VTAIL.t5 149.524
R231 VTAIL.n171 VTAIL.t6 149.524
R232 VTAIL.n376 VTAIL.n375 104.615
R233 VTAIL.n376 VTAIL.n369 104.615
R234 VTAIL.n383 VTAIL.n369 104.615
R235 VTAIL.n384 VTAIL.n383 104.615
R236 VTAIL.n384 VTAIL.n365 104.615
R237 VTAIL.n392 VTAIL.n365 104.615
R238 VTAIL.n393 VTAIL.n392 104.615
R239 VTAIL.n394 VTAIL.n393 104.615
R240 VTAIL.n394 VTAIL.n361 104.615
R241 VTAIL.n401 VTAIL.n361 104.615
R242 VTAIL.n402 VTAIL.n401 104.615
R243 VTAIL.n20 VTAIL.n19 104.615
R244 VTAIL.n20 VTAIL.n13 104.615
R245 VTAIL.n27 VTAIL.n13 104.615
R246 VTAIL.n28 VTAIL.n27 104.615
R247 VTAIL.n28 VTAIL.n9 104.615
R248 VTAIL.n36 VTAIL.n9 104.615
R249 VTAIL.n37 VTAIL.n36 104.615
R250 VTAIL.n38 VTAIL.n37 104.615
R251 VTAIL.n38 VTAIL.n5 104.615
R252 VTAIL.n45 VTAIL.n5 104.615
R253 VTAIL.n46 VTAIL.n45 104.615
R254 VTAIL.n70 VTAIL.n69 104.615
R255 VTAIL.n70 VTAIL.n63 104.615
R256 VTAIL.n77 VTAIL.n63 104.615
R257 VTAIL.n78 VTAIL.n77 104.615
R258 VTAIL.n78 VTAIL.n59 104.615
R259 VTAIL.n86 VTAIL.n59 104.615
R260 VTAIL.n87 VTAIL.n86 104.615
R261 VTAIL.n88 VTAIL.n87 104.615
R262 VTAIL.n88 VTAIL.n55 104.615
R263 VTAIL.n95 VTAIL.n55 104.615
R264 VTAIL.n96 VTAIL.n95 104.615
R265 VTAIL.n122 VTAIL.n121 104.615
R266 VTAIL.n122 VTAIL.n115 104.615
R267 VTAIL.n129 VTAIL.n115 104.615
R268 VTAIL.n130 VTAIL.n129 104.615
R269 VTAIL.n130 VTAIL.n111 104.615
R270 VTAIL.n138 VTAIL.n111 104.615
R271 VTAIL.n139 VTAIL.n138 104.615
R272 VTAIL.n140 VTAIL.n139 104.615
R273 VTAIL.n140 VTAIL.n107 104.615
R274 VTAIL.n147 VTAIL.n107 104.615
R275 VTAIL.n148 VTAIL.n147 104.615
R276 VTAIL.n352 VTAIL.n351 104.615
R277 VTAIL.n351 VTAIL.n311 104.615
R278 VTAIL.n316 VTAIL.n311 104.615
R279 VTAIL.n344 VTAIL.n316 104.615
R280 VTAIL.n344 VTAIL.n343 104.615
R281 VTAIL.n343 VTAIL.n317 104.615
R282 VTAIL.n336 VTAIL.n317 104.615
R283 VTAIL.n336 VTAIL.n335 104.615
R284 VTAIL.n335 VTAIL.n321 104.615
R285 VTAIL.n328 VTAIL.n321 104.615
R286 VTAIL.n328 VTAIL.n327 104.615
R287 VTAIL.n300 VTAIL.n299 104.615
R288 VTAIL.n299 VTAIL.n259 104.615
R289 VTAIL.n264 VTAIL.n259 104.615
R290 VTAIL.n292 VTAIL.n264 104.615
R291 VTAIL.n292 VTAIL.n291 104.615
R292 VTAIL.n291 VTAIL.n265 104.615
R293 VTAIL.n284 VTAIL.n265 104.615
R294 VTAIL.n284 VTAIL.n283 104.615
R295 VTAIL.n283 VTAIL.n269 104.615
R296 VTAIL.n276 VTAIL.n269 104.615
R297 VTAIL.n276 VTAIL.n275 104.615
R298 VTAIL.n250 VTAIL.n249 104.615
R299 VTAIL.n249 VTAIL.n209 104.615
R300 VTAIL.n214 VTAIL.n209 104.615
R301 VTAIL.n242 VTAIL.n214 104.615
R302 VTAIL.n242 VTAIL.n241 104.615
R303 VTAIL.n241 VTAIL.n215 104.615
R304 VTAIL.n234 VTAIL.n215 104.615
R305 VTAIL.n234 VTAIL.n233 104.615
R306 VTAIL.n233 VTAIL.n219 104.615
R307 VTAIL.n226 VTAIL.n219 104.615
R308 VTAIL.n226 VTAIL.n225 104.615
R309 VTAIL.n198 VTAIL.n197 104.615
R310 VTAIL.n197 VTAIL.n157 104.615
R311 VTAIL.n162 VTAIL.n157 104.615
R312 VTAIL.n190 VTAIL.n162 104.615
R313 VTAIL.n190 VTAIL.n189 104.615
R314 VTAIL.n189 VTAIL.n163 104.615
R315 VTAIL.n182 VTAIL.n163 104.615
R316 VTAIL.n182 VTAIL.n181 104.615
R317 VTAIL.n181 VTAIL.n167 104.615
R318 VTAIL.n174 VTAIL.n167 104.615
R319 VTAIL.n174 VTAIL.n173 104.615
R320 VTAIL.n375 VTAIL.t15 52.3082
R321 VTAIL.n19 VTAIL.t1 52.3082
R322 VTAIL.n69 VTAIL.t12 52.3082
R323 VTAIL.n121 VTAIL.t8 52.3082
R324 VTAIL.n327 VTAIL.t9 52.3082
R325 VTAIL.n275 VTAIL.t7 52.3082
R326 VTAIL.n225 VTAIL.t5 52.3082
R327 VTAIL.n173 VTAIL.t6 52.3082
R328 VTAIL.n307 VTAIL.n306 49.2323
R329 VTAIL.n205 VTAIL.n204 49.2323
R330 VTAIL.n1 VTAIL.n0 49.2322
R331 VTAIL.n103 VTAIL.n102 49.2322
R332 VTAIL.n407 VTAIL.n406 35.0944
R333 VTAIL.n51 VTAIL.n50 35.0944
R334 VTAIL.n101 VTAIL.n100 35.0944
R335 VTAIL.n153 VTAIL.n152 35.0944
R336 VTAIL.n357 VTAIL.n356 35.0944
R337 VTAIL.n305 VTAIL.n304 35.0944
R338 VTAIL.n255 VTAIL.n254 35.0944
R339 VTAIL.n203 VTAIL.n202 35.0944
R340 VTAIL.n407 VTAIL.n357 23.2289
R341 VTAIL.n203 VTAIL.n153 23.2289
R342 VTAIL.n395 VTAIL.n362 13.1884
R343 VTAIL.n39 VTAIL.n6 13.1884
R344 VTAIL.n89 VTAIL.n56 13.1884
R345 VTAIL.n141 VTAIL.n108 13.1884
R346 VTAIL.n314 VTAIL.n312 13.1884
R347 VTAIL.n262 VTAIL.n260 13.1884
R348 VTAIL.n212 VTAIL.n210 13.1884
R349 VTAIL.n160 VTAIL.n158 13.1884
R350 VTAIL.n396 VTAIL.n364 12.8005
R351 VTAIL.n400 VTAIL.n399 12.8005
R352 VTAIL.n40 VTAIL.n8 12.8005
R353 VTAIL.n44 VTAIL.n43 12.8005
R354 VTAIL.n90 VTAIL.n58 12.8005
R355 VTAIL.n94 VTAIL.n93 12.8005
R356 VTAIL.n142 VTAIL.n110 12.8005
R357 VTAIL.n146 VTAIL.n145 12.8005
R358 VTAIL.n350 VTAIL.n349 12.8005
R359 VTAIL.n346 VTAIL.n345 12.8005
R360 VTAIL.n298 VTAIL.n297 12.8005
R361 VTAIL.n294 VTAIL.n293 12.8005
R362 VTAIL.n248 VTAIL.n247 12.8005
R363 VTAIL.n244 VTAIL.n243 12.8005
R364 VTAIL.n196 VTAIL.n195 12.8005
R365 VTAIL.n192 VTAIL.n191 12.8005
R366 VTAIL.n391 VTAIL.n390 12.0247
R367 VTAIL.n403 VTAIL.n360 12.0247
R368 VTAIL.n35 VTAIL.n34 12.0247
R369 VTAIL.n47 VTAIL.n4 12.0247
R370 VTAIL.n85 VTAIL.n84 12.0247
R371 VTAIL.n97 VTAIL.n54 12.0247
R372 VTAIL.n137 VTAIL.n136 12.0247
R373 VTAIL.n149 VTAIL.n106 12.0247
R374 VTAIL.n353 VTAIL.n310 12.0247
R375 VTAIL.n342 VTAIL.n315 12.0247
R376 VTAIL.n301 VTAIL.n258 12.0247
R377 VTAIL.n290 VTAIL.n263 12.0247
R378 VTAIL.n251 VTAIL.n208 12.0247
R379 VTAIL.n240 VTAIL.n213 12.0247
R380 VTAIL.n199 VTAIL.n156 12.0247
R381 VTAIL.n188 VTAIL.n161 12.0247
R382 VTAIL.n389 VTAIL.n366 11.249
R383 VTAIL.n404 VTAIL.n358 11.249
R384 VTAIL.n33 VTAIL.n10 11.249
R385 VTAIL.n48 VTAIL.n2 11.249
R386 VTAIL.n83 VTAIL.n60 11.249
R387 VTAIL.n98 VTAIL.n52 11.249
R388 VTAIL.n135 VTAIL.n112 11.249
R389 VTAIL.n150 VTAIL.n104 11.249
R390 VTAIL.n354 VTAIL.n308 11.249
R391 VTAIL.n341 VTAIL.n318 11.249
R392 VTAIL.n302 VTAIL.n256 11.249
R393 VTAIL.n289 VTAIL.n266 11.249
R394 VTAIL.n252 VTAIL.n206 11.249
R395 VTAIL.n239 VTAIL.n216 11.249
R396 VTAIL.n200 VTAIL.n154 11.249
R397 VTAIL.n187 VTAIL.n164 11.249
R398 VTAIL.n386 VTAIL.n385 10.4732
R399 VTAIL.n30 VTAIL.n29 10.4732
R400 VTAIL.n80 VTAIL.n79 10.4732
R401 VTAIL.n132 VTAIL.n131 10.4732
R402 VTAIL.n338 VTAIL.n337 10.4732
R403 VTAIL.n286 VTAIL.n285 10.4732
R404 VTAIL.n236 VTAIL.n235 10.4732
R405 VTAIL.n184 VTAIL.n183 10.4732
R406 VTAIL.n374 VTAIL.n373 10.2747
R407 VTAIL.n18 VTAIL.n17 10.2747
R408 VTAIL.n68 VTAIL.n67 10.2747
R409 VTAIL.n120 VTAIL.n119 10.2747
R410 VTAIL.n326 VTAIL.n325 10.2747
R411 VTAIL.n274 VTAIL.n273 10.2747
R412 VTAIL.n224 VTAIL.n223 10.2747
R413 VTAIL.n172 VTAIL.n171 10.2747
R414 VTAIL.n382 VTAIL.n368 9.69747
R415 VTAIL.n26 VTAIL.n12 9.69747
R416 VTAIL.n76 VTAIL.n62 9.69747
R417 VTAIL.n128 VTAIL.n114 9.69747
R418 VTAIL.n334 VTAIL.n320 9.69747
R419 VTAIL.n282 VTAIL.n268 9.69747
R420 VTAIL.n232 VTAIL.n218 9.69747
R421 VTAIL.n180 VTAIL.n166 9.69747
R422 VTAIL.n406 VTAIL.n405 9.45567
R423 VTAIL.n50 VTAIL.n49 9.45567
R424 VTAIL.n100 VTAIL.n99 9.45567
R425 VTAIL.n152 VTAIL.n151 9.45567
R426 VTAIL.n356 VTAIL.n355 9.45567
R427 VTAIL.n304 VTAIL.n303 9.45567
R428 VTAIL.n254 VTAIL.n253 9.45567
R429 VTAIL.n202 VTAIL.n201 9.45567
R430 VTAIL.n405 VTAIL.n404 9.3005
R431 VTAIL.n360 VTAIL.n359 9.3005
R432 VTAIL.n399 VTAIL.n398 9.3005
R433 VTAIL.n372 VTAIL.n371 9.3005
R434 VTAIL.n379 VTAIL.n378 9.3005
R435 VTAIL.n381 VTAIL.n380 9.3005
R436 VTAIL.n368 VTAIL.n367 9.3005
R437 VTAIL.n387 VTAIL.n386 9.3005
R438 VTAIL.n389 VTAIL.n388 9.3005
R439 VTAIL.n390 VTAIL.n363 9.3005
R440 VTAIL.n397 VTAIL.n396 9.3005
R441 VTAIL.n49 VTAIL.n48 9.3005
R442 VTAIL.n4 VTAIL.n3 9.3005
R443 VTAIL.n43 VTAIL.n42 9.3005
R444 VTAIL.n16 VTAIL.n15 9.3005
R445 VTAIL.n23 VTAIL.n22 9.3005
R446 VTAIL.n25 VTAIL.n24 9.3005
R447 VTAIL.n12 VTAIL.n11 9.3005
R448 VTAIL.n31 VTAIL.n30 9.3005
R449 VTAIL.n33 VTAIL.n32 9.3005
R450 VTAIL.n34 VTAIL.n7 9.3005
R451 VTAIL.n41 VTAIL.n40 9.3005
R452 VTAIL.n99 VTAIL.n98 9.3005
R453 VTAIL.n54 VTAIL.n53 9.3005
R454 VTAIL.n93 VTAIL.n92 9.3005
R455 VTAIL.n66 VTAIL.n65 9.3005
R456 VTAIL.n73 VTAIL.n72 9.3005
R457 VTAIL.n75 VTAIL.n74 9.3005
R458 VTAIL.n62 VTAIL.n61 9.3005
R459 VTAIL.n81 VTAIL.n80 9.3005
R460 VTAIL.n83 VTAIL.n82 9.3005
R461 VTAIL.n84 VTAIL.n57 9.3005
R462 VTAIL.n91 VTAIL.n90 9.3005
R463 VTAIL.n151 VTAIL.n150 9.3005
R464 VTAIL.n106 VTAIL.n105 9.3005
R465 VTAIL.n145 VTAIL.n144 9.3005
R466 VTAIL.n118 VTAIL.n117 9.3005
R467 VTAIL.n125 VTAIL.n124 9.3005
R468 VTAIL.n127 VTAIL.n126 9.3005
R469 VTAIL.n114 VTAIL.n113 9.3005
R470 VTAIL.n133 VTAIL.n132 9.3005
R471 VTAIL.n135 VTAIL.n134 9.3005
R472 VTAIL.n136 VTAIL.n109 9.3005
R473 VTAIL.n143 VTAIL.n142 9.3005
R474 VTAIL.n324 VTAIL.n323 9.3005
R475 VTAIL.n331 VTAIL.n330 9.3005
R476 VTAIL.n333 VTAIL.n332 9.3005
R477 VTAIL.n320 VTAIL.n319 9.3005
R478 VTAIL.n339 VTAIL.n338 9.3005
R479 VTAIL.n341 VTAIL.n340 9.3005
R480 VTAIL.n315 VTAIL.n313 9.3005
R481 VTAIL.n347 VTAIL.n346 9.3005
R482 VTAIL.n355 VTAIL.n354 9.3005
R483 VTAIL.n310 VTAIL.n309 9.3005
R484 VTAIL.n349 VTAIL.n348 9.3005
R485 VTAIL.n272 VTAIL.n271 9.3005
R486 VTAIL.n279 VTAIL.n278 9.3005
R487 VTAIL.n281 VTAIL.n280 9.3005
R488 VTAIL.n268 VTAIL.n267 9.3005
R489 VTAIL.n287 VTAIL.n286 9.3005
R490 VTAIL.n289 VTAIL.n288 9.3005
R491 VTAIL.n263 VTAIL.n261 9.3005
R492 VTAIL.n295 VTAIL.n294 9.3005
R493 VTAIL.n303 VTAIL.n302 9.3005
R494 VTAIL.n258 VTAIL.n257 9.3005
R495 VTAIL.n297 VTAIL.n296 9.3005
R496 VTAIL.n222 VTAIL.n221 9.3005
R497 VTAIL.n229 VTAIL.n228 9.3005
R498 VTAIL.n231 VTAIL.n230 9.3005
R499 VTAIL.n218 VTAIL.n217 9.3005
R500 VTAIL.n237 VTAIL.n236 9.3005
R501 VTAIL.n239 VTAIL.n238 9.3005
R502 VTAIL.n213 VTAIL.n211 9.3005
R503 VTAIL.n245 VTAIL.n244 9.3005
R504 VTAIL.n253 VTAIL.n252 9.3005
R505 VTAIL.n208 VTAIL.n207 9.3005
R506 VTAIL.n247 VTAIL.n246 9.3005
R507 VTAIL.n170 VTAIL.n169 9.3005
R508 VTAIL.n177 VTAIL.n176 9.3005
R509 VTAIL.n179 VTAIL.n178 9.3005
R510 VTAIL.n166 VTAIL.n165 9.3005
R511 VTAIL.n185 VTAIL.n184 9.3005
R512 VTAIL.n187 VTAIL.n186 9.3005
R513 VTAIL.n161 VTAIL.n159 9.3005
R514 VTAIL.n193 VTAIL.n192 9.3005
R515 VTAIL.n201 VTAIL.n200 9.3005
R516 VTAIL.n156 VTAIL.n155 9.3005
R517 VTAIL.n195 VTAIL.n194 9.3005
R518 VTAIL.n381 VTAIL.n370 8.92171
R519 VTAIL.n25 VTAIL.n14 8.92171
R520 VTAIL.n75 VTAIL.n64 8.92171
R521 VTAIL.n127 VTAIL.n116 8.92171
R522 VTAIL.n333 VTAIL.n322 8.92171
R523 VTAIL.n281 VTAIL.n270 8.92171
R524 VTAIL.n231 VTAIL.n220 8.92171
R525 VTAIL.n179 VTAIL.n168 8.92171
R526 VTAIL.n378 VTAIL.n377 8.14595
R527 VTAIL.n22 VTAIL.n21 8.14595
R528 VTAIL.n72 VTAIL.n71 8.14595
R529 VTAIL.n124 VTAIL.n123 8.14595
R530 VTAIL.n330 VTAIL.n329 8.14595
R531 VTAIL.n278 VTAIL.n277 8.14595
R532 VTAIL.n228 VTAIL.n227 8.14595
R533 VTAIL.n176 VTAIL.n175 8.14595
R534 VTAIL.n374 VTAIL.n372 7.3702
R535 VTAIL.n18 VTAIL.n16 7.3702
R536 VTAIL.n68 VTAIL.n66 7.3702
R537 VTAIL.n120 VTAIL.n118 7.3702
R538 VTAIL.n326 VTAIL.n324 7.3702
R539 VTAIL.n274 VTAIL.n272 7.3702
R540 VTAIL.n224 VTAIL.n222 7.3702
R541 VTAIL.n172 VTAIL.n170 7.3702
R542 VTAIL.n377 VTAIL.n372 5.81868
R543 VTAIL.n21 VTAIL.n16 5.81868
R544 VTAIL.n71 VTAIL.n66 5.81868
R545 VTAIL.n123 VTAIL.n118 5.81868
R546 VTAIL.n329 VTAIL.n324 5.81868
R547 VTAIL.n277 VTAIL.n272 5.81868
R548 VTAIL.n227 VTAIL.n222 5.81868
R549 VTAIL.n175 VTAIL.n170 5.81868
R550 VTAIL.n378 VTAIL.n370 5.04292
R551 VTAIL.n22 VTAIL.n14 5.04292
R552 VTAIL.n72 VTAIL.n64 5.04292
R553 VTAIL.n124 VTAIL.n116 5.04292
R554 VTAIL.n330 VTAIL.n322 5.04292
R555 VTAIL.n278 VTAIL.n270 5.04292
R556 VTAIL.n228 VTAIL.n220 5.04292
R557 VTAIL.n176 VTAIL.n168 5.04292
R558 VTAIL.n382 VTAIL.n381 4.26717
R559 VTAIL.n26 VTAIL.n25 4.26717
R560 VTAIL.n76 VTAIL.n75 4.26717
R561 VTAIL.n128 VTAIL.n127 4.26717
R562 VTAIL.n334 VTAIL.n333 4.26717
R563 VTAIL.n282 VTAIL.n281 4.26717
R564 VTAIL.n232 VTAIL.n231 4.26717
R565 VTAIL.n180 VTAIL.n179 4.26717
R566 VTAIL.n385 VTAIL.n368 3.49141
R567 VTAIL.n29 VTAIL.n12 3.49141
R568 VTAIL.n79 VTAIL.n62 3.49141
R569 VTAIL.n131 VTAIL.n114 3.49141
R570 VTAIL.n337 VTAIL.n320 3.49141
R571 VTAIL.n285 VTAIL.n268 3.49141
R572 VTAIL.n235 VTAIL.n218 3.49141
R573 VTAIL.n183 VTAIL.n166 3.49141
R574 VTAIL.n373 VTAIL.n371 2.84303
R575 VTAIL.n17 VTAIL.n15 2.84303
R576 VTAIL.n67 VTAIL.n65 2.84303
R577 VTAIL.n119 VTAIL.n117 2.84303
R578 VTAIL.n325 VTAIL.n323 2.84303
R579 VTAIL.n273 VTAIL.n271 2.84303
R580 VTAIL.n223 VTAIL.n221 2.84303
R581 VTAIL.n171 VTAIL.n169 2.84303
R582 VTAIL.n205 VTAIL.n203 2.76774
R583 VTAIL.n255 VTAIL.n205 2.76774
R584 VTAIL.n307 VTAIL.n305 2.76774
R585 VTAIL.n357 VTAIL.n307 2.76774
R586 VTAIL.n153 VTAIL.n103 2.76774
R587 VTAIL.n103 VTAIL.n101 2.76774
R588 VTAIL.n51 VTAIL.n1 2.76774
R589 VTAIL.n386 VTAIL.n366 2.71565
R590 VTAIL.n406 VTAIL.n358 2.71565
R591 VTAIL.n30 VTAIL.n10 2.71565
R592 VTAIL.n50 VTAIL.n2 2.71565
R593 VTAIL.n80 VTAIL.n60 2.71565
R594 VTAIL.n100 VTAIL.n52 2.71565
R595 VTAIL.n132 VTAIL.n112 2.71565
R596 VTAIL.n152 VTAIL.n104 2.71565
R597 VTAIL.n356 VTAIL.n308 2.71565
R598 VTAIL.n338 VTAIL.n318 2.71565
R599 VTAIL.n304 VTAIL.n256 2.71565
R600 VTAIL.n286 VTAIL.n266 2.71565
R601 VTAIL.n254 VTAIL.n206 2.71565
R602 VTAIL.n236 VTAIL.n216 2.71565
R603 VTAIL.n202 VTAIL.n154 2.71565
R604 VTAIL.n184 VTAIL.n164 2.71565
R605 VTAIL VTAIL.n407 2.70955
R606 VTAIL.n0 VTAIL.t4 2.10913
R607 VTAIL.n0 VTAIL.t2 2.10913
R608 VTAIL.n102 VTAIL.t14 2.10913
R609 VTAIL.n102 VTAIL.t10 2.10913
R610 VTAIL.n306 VTAIL.t11 2.10913
R611 VTAIL.n306 VTAIL.t13 2.10913
R612 VTAIL.n204 VTAIL.t3 2.10913
R613 VTAIL.n204 VTAIL.t0 2.10913
R614 VTAIL.n391 VTAIL.n389 1.93989
R615 VTAIL.n404 VTAIL.n403 1.93989
R616 VTAIL.n35 VTAIL.n33 1.93989
R617 VTAIL.n48 VTAIL.n47 1.93989
R618 VTAIL.n85 VTAIL.n83 1.93989
R619 VTAIL.n98 VTAIL.n97 1.93989
R620 VTAIL.n137 VTAIL.n135 1.93989
R621 VTAIL.n150 VTAIL.n149 1.93989
R622 VTAIL.n354 VTAIL.n353 1.93989
R623 VTAIL.n342 VTAIL.n341 1.93989
R624 VTAIL.n302 VTAIL.n301 1.93989
R625 VTAIL.n290 VTAIL.n289 1.93989
R626 VTAIL.n252 VTAIL.n251 1.93989
R627 VTAIL.n240 VTAIL.n239 1.93989
R628 VTAIL.n200 VTAIL.n199 1.93989
R629 VTAIL.n188 VTAIL.n187 1.93989
R630 VTAIL.n390 VTAIL.n364 1.16414
R631 VTAIL.n400 VTAIL.n360 1.16414
R632 VTAIL.n34 VTAIL.n8 1.16414
R633 VTAIL.n44 VTAIL.n4 1.16414
R634 VTAIL.n84 VTAIL.n58 1.16414
R635 VTAIL.n94 VTAIL.n54 1.16414
R636 VTAIL.n136 VTAIL.n110 1.16414
R637 VTAIL.n146 VTAIL.n106 1.16414
R638 VTAIL.n350 VTAIL.n310 1.16414
R639 VTAIL.n345 VTAIL.n315 1.16414
R640 VTAIL.n298 VTAIL.n258 1.16414
R641 VTAIL.n293 VTAIL.n263 1.16414
R642 VTAIL.n248 VTAIL.n208 1.16414
R643 VTAIL.n243 VTAIL.n213 1.16414
R644 VTAIL.n196 VTAIL.n156 1.16414
R645 VTAIL.n191 VTAIL.n161 1.16414
R646 VTAIL.n305 VTAIL.n255 0.470328
R647 VTAIL.n101 VTAIL.n51 0.470328
R648 VTAIL.n396 VTAIL.n395 0.388379
R649 VTAIL.n399 VTAIL.n362 0.388379
R650 VTAIL.n40 VTAIL.n39 0.388379
R651 VTAIL.n43 VTAIL.n6 0.388379
R652 VTAIL.n90 VTAIL.n89 0.388379
R653 VTAIL.n93 VTAIL.n56 0.388379
R654 VTAIL.n142 VTAIL.n141 0.388379
R655 VTAIL.n145 VTAIL.n108 0.388379
R656 VTAIL.n349 VTAIL.n312 0.388379
R657 VTAIL.n346 VTAIL.n314 0.388379
R658 VTAIL.n297 VTAIL.n260 0.388379
R659 VTAIL.n294 VTAIL.n262 0.388379
R660 VTAIL.n247 VTAIL.n210 0.388379
R661 VTAIL.n244 VTAIL.n212 0.388379
R662 VTAIL.n195 VTAIL.n158 0.388379
R663 VTAIL.n192 VTAIL.n160 0.388379
R664 VTAIL.n379 VTAIL.n371 0.155672
R665 VTAIL.n380 VTAIL.n379 0.155672
R666 VTAIL.n380 VTAIL.n367 0.155672
R667 VTAIL.n387 VTAIL.n367 0.155672
R668 VTAIL.n388 VTAIL.n387 0.155672
R669 VTAIL.n388 VTAIL.n363 0.155672
R670 VTAIL.n397 VTAIL.n363 0.155672
R671 VTAIL.n398 VTAIL.n397 0.155672
R672 VTAIL.n398 VTAIL.n359 0.155672
R673 VTAIL.n405 VTAIL.n359 0.155672
R674 VTAIL.n23 VTAIL.n15 0.155672
R675 VTAIL.n24 VTAIL.n23 0.155672
R676 VTAIL.n24 VTAIL.n11 0.155672
R677 VTAIL.n31 VTAIL.n11 0.155672
R678 VTAIL.n32 VTAIL.n31 0.155672
R679 VTAIL.n32 VTAIL.n7 0.155672
R680 VTAIL.n41 VTAIL.n7 0.155672
R681 VTAIL.n42 VTAIL.n41 0.155672
R682 VTAIL.n42 VTAIL.n3 0.155672
R683 VTAIL.n49 VTAIL.n3 0.155672
R684 VTAIL.n73 VTAIL.n65 0.155672
R685 VTAIL.n74 VTAIL.n73 0.155672
R686 VTAIL.n74 VTAIL.n61 0.155672
R687 VTAIL.n81 VTAIL.n61 0.155672
R688 VTAIL.n82 VTAIL.n81 0.155672
R689 VTAIL.n82 VTAIL.n57 0.155672
R690 VTAIL.n91 VTAIL.n57 0.155672
R691 VTAIL.n92 VTAIL.n91 0.155672
R692 VTAIL.n92 VTAIL.n53 0.155672
R693 VTAIL.n99 VTAIL.n53 0.155672
R694 VTAIL.n125 VTAIL.n117 0.155672
R695 VTAIL.n126 VTAIL.n125 0.155672
R696 VTAIL.n126 VTAIL.n113 0.155672
R697 VTAIL.n133 VTAIL.n113 0.155672
R698 VTAIL.n134 VTAIL.n133 0.155672
R699 VTAIL.n134 VTAIL.n109 0.155672
R700 VTAIL.n143 VTAIL.n109 0.155672
R701 VTAIL.n144 VTAIL.n143 0.155672
R702 VTAIL.n144 VTAIL.n105 0.155672
R703 VTAIL.n151 VTAIL.n105 0.155672
R704 VTAIL.n355 VTAIL.n309 0.155672
R705 VTAIL.n348 VTAIL.n309 0.155672
R706 VTAIL.n348 VTAIL.n347 0.155672
R707 VTAIL.n347 VTAIL.n313 0.155672
R708 VTAIL.n340 VTAIL.n313 0.155672
R709 VTAIL.n340 VTAIL.n339 0.155672
R710 VTAIL.n339 VTAIL.n319 0.155672
R711 VTAIL.n332 VTAIL.n319 0.155672
R712 VTAIL.n332 VTAIL.n331 0.155672
R713 VTAIL.n331 VTAIL.n323 0.155672
R714 VTAIL.n303 VTAIL.n257 0.155672
R715 VTAIL.n296 VTAIL.n257 0.155672
R716 VTAIL.n296 VTAIL.n295 0.155672
R717 VTAIL.n295 VTAIL.n261 0.155672
R718 VTAIL.n288 VTAIL.n261 0.155672
R719 VTAIL.n288 VTAIL.n287 0.155672
R720 VTAIL.n287 VTAIL.n267 0.155672
R721 VTAIL.n280 VTAIL.n267 0.155672
R722 VTAIL.n280 VTAIL.n279 0.155672
R723 VTAIL.n279 VTAIL.n271 0.155672
R724 VTAIL.n253 VTAIL.n207 0.155672
R725 VTAIL.n246 VTAIL.n207 0.155672
R726 VTAIL.n246 VTAIL.n245 0.155672
R727 VTAIL.n245 VTAIL.n211 0.155672
R728 VTAIL.n238 VTAIL.n211 0.155672
R729 VTAIL.n238 VTAIL.n237 0.155672
R730 VTAIL.n237 VTAIL.n217 0.155672
R731 VTAIL.n230 VTAIL.n217 0.155672
R732 VTAIL.n230 VTAIL.n229 0.155672
R733 VTAIL.n229 VTAIL.n221 0.155672
R734 VTAIL.n201 VTAIL.n155 0.155672
R735 VTAIL.n194 VTAIL.n155 0.155672
R736 VTAIL.n194 VTAIL.n193 0.155672
R737 VTAIL.n193 VTAIL.n159 0.155672
R738 VTAIL.n186 VTAIL.n159 0.155672
R739 VTAIL.n186 VTAIL.n185 0.155672
R740 VTAIL.n185 VTAIL.n165 0.155672
R741 VTAIL.n178 VTAIL.n165 0.155672
R742 VTAIL.n178 VTAIL.n177 0.155672
R743 VTAIL.n177 VTAIL.n169 0.155672
R744 VTAIL VTAIL.n1 0.0586897
R745 VDD1 VDD1.n0 67.3529
R746 VDD1.n3 VDD1.n2 67.2392
R747 VDD1.n3 VDD1.n1 67.2392
R748 VDD1.n5 VDD1.n4 65.911
R749 VDD1.n5 VDD1.n3 44.8457
R750 VDD1.n4 VDD1.t1 2.10913
R751 VDD1.n4 VDD1.t5 2.10913
R752 VDD1.n0 VDD1.t0 2.10913
R753 VDD1.n0 VDD1.t7 2.10913
R754 VDD1.n2 VDD1.t4 2.10913
R755 VDD1.n2 VDD1.t2 2.10913
R756 VDD1.n1 VDD1.t6 2.10913
R757 VDD1.n1 VDD1.t3 2.10913
R758 VDD1 VDD1.n5 1.32593
R759 B.n839 B.n838 585
R760 B.n840 B.n839 585
R761 B.n295 B.n141 585
R762 B.n294 B.n293 585
R763 B.n292 B.n291 585
R764 B.n290 B.n289 585
R765 B.n288 B.n287 585
R766 B.n286 B.n285 585
R767 B.n284 B.n283 585
R768 B.n282 B.n281 585
R769 B.n280 B.n279 585
R770 B.n278 B.n277 585
R771 B.n276 B.n275 585
R772 B.n274 B.n273 585
R773 B.n272 B.n271 585
R774 B.n270 B.n269 585
R775 B.n268 B.n267 585
R776 B.n266 B.n265 585
R777 B.n264 B.n263 585
R778 B.n262 B.n261 585
R779 B.n260 B.n259 585
R780 B.n258 B.n257 585
R781 B.n256 B.n255 585
R782 B.n254 B.n253 585
R783 B.n252 B.n251 585
R784 B.n250 B.n249 585
R785 B.n248 B.n247 585
R786 B.n246 B.n245 585
R787 B.n244 B.n243 585
R788 B.n242 B.n241 585
R789 B.n240 B.n239 585
R790 B.n238 B.n237 585
R791 B.n236 B.n235 585
R792 B.n234 B.n233 585
R793 B.n232 B.n231 585
R794 B.n229 B.n228 585
R795 B.n227 B.n226 585
R796 B.n225 B.n224 585
R797 B.n223 B.n222 585
R798 B.n221 B.n220 585
R799 B.n219 B.n218 585
R800 B.n217 B.n216 585
R801 B.n215 B.n214 585
R802 B.n213 B.n212 585
R803 B.n211 B.n210 585
R804 B.n209 B.n208 585
R805 B.n207 B.n206 585
R806 B.n205 B.n204 585
R807 B.n203 B.n202 585
R808 B.n201 B.n200 585
R809 B.n199 B.n198 585
R810 B.n197 B.n196 585
R811 B.n195 B.n194 585
R812 B.n193 B.n192 585
R813 B.n191 B.n190 585
R814 B.n189 B.n188 585
R815 B.n187 B.n186 585
R816 B.n185 B.n184 585
R817 B.n183 B.n182 585
R818 B.n181 B.n180 585
R819 B.n179 B.n178 585
R820 B.n177 B.n176 585
R821 B.n175 B.n174 585
R822 B.n173 B.n172 585
R823 B.n171 B.n170 585
R824 B.n169 B.n168 585
R825 B.n167 B.n166 585
R826 B.n165 B.n164 585
R827 B.n163 B.n162 585
R828 B.n161 B.n160 585
R829 B.n159 B.n158 585
R830 B.n157 B.n156 585
R831 B.n155 B.n154 585
R832 B.n153 B.n152 585
R833 B.n151 B.n150 585
R834 B.n149 B.n148 585
R835 B.n103 B.n102 585
R836 B.n843 B.n842 585
R837 B.n837 B.n142 585
R838 B.n142 B.n100 585
R839 B.n836 B.n99 585
R840 B.n847 B.n99 585
R841 B.n835 B.n98 585
R842 B.n848 B.n98 585
R843 B.n834 B.n97 585
R844 B.n849 B.n97 585
R845 B.n833 B.n832 585
R846 B.n832 B.n93 585
R847 B.n831 B.n92 585
R848 B.n855 B.n92 585
R849 B.n830 B.n91 585
R850 B.n856 B.n91 585
R851 B.n829 B.n90 585
R852 B.n857 B.n90 585
R853 B.n828 B.n827 585
R854 B.n827 B.n89 585
R855 B.n826 B.n85 585
R856 B.n863 B.n85 585
R857 B.n825 B.n84 585
R858 B.n864 B.n84 585
R859 B.n824 B.n83 585
R860 B.n865 B.n83 585
R861 B.n823 B.n822 585
R862 B.n822 B.n79 585
R863 B.n821 B.n78 585
R864 B.n871 B.n78 585
R865 B.n820 B.n77 585
R866 B.n872 B.n77 585
R867 B.n819 B.n76 585
R868 B.n873 B.n76 585
R869 B.n818 B.n817 585
R870 B.n817 B.n72 585
R871 B.n816 B.n71 585
R872 B.n879 B.n71 585
R873 B.n815 B.n70 585
R874 B.n880 B.n70 585
R875 B.n814 B.n69 585
R876 B.n881 B.n69 585
R877 B.n813 B.n812 585
R878 B.n812 B.n68 585
R879 B.n811 B.n64 585
R880 B.n887 B.n64 585
R881 B.n810 B.n63 585
R882 B.n888 B.n63 585
R883 B.n809 B.n62 585
R884 B.n889 B.n62 585
R885 B.n808 B.n807 585
R886 B.n807 B.n58 585
R887 B.n806 B.n57 585
R888 B.n895 B.n57 585
R889 B.n805 B.n56 585
R890 B.n896 B.n56 585
R891 B.n804 B.n55 585
R892 B.n897 B.n55 585
R893 B.n803 B.n802 585
R894 B.n802 B.n51 585
R895 B.n801 B.n50 585
R896 B.n903 B.n50 585
R897 B.n800 B.n49 585
R898 B.n904 B.n49 585
R899 B.n799 B.n48 585
R900 B.n905 B.n48 585
R901 B.n798 B.n797 585
R902 B.n797 B.n44 585
R903 B.n796 B.n43 585
R904 B.n911 B.n43 585
R905 B.n795 B.n42 585
R906 B.n912 B.n42 585
R907 B.n794 B.n41 585
R908 B.n913 B.n41 585
R909 B.n793 B.n792 585
R910 B.n792 B.n37 585
R911 B.n791 B.n36 585
R912 B.n919 B.n36 585
R913 B.n790 B.n35 585
R914 B.n920 B.n35 585
R915 B.n789 B.n34 585
R916 B.n921 B.n34 585
R917 B.n788 B.n787 585
R918 B.n787 B.n30 585
R919 B.n786 B.n29 585
R920 B.n927 B.n29 585
R921 B.n785 B.n28 585
R922 B.n928 B.n28 585
R923 B.n784 B.n27 585
R924 B.n929 B.n27 585
R925 B.n783 B.n782 585
R926 B.n782 B.n23 585
R927 B.n781 B.n22 585
R928 B.n935 B.n22 585
R929 B.n780 B.n21 585
R930 B.n936 B.n21 585
R931 B.n779 B.n20 585
R932 B.n937 B.n20 585
R933 B.n778 B.n777 585
R934 B.n777 B.n16 585
R935 B.n776 B.n15 585
R936 B.n943 B.n15 585
R937 B.n775 B.n14 585
R938 B.n944 B.n14 585
R939 B.n774 B.n13 585
R940 B.n945 B.n13 585
R941 B.n773 B.n772 585
R942 B.n772 B.n12 585
R943 B.n771 B.n770 585
R944 B.n771 B.n8 585
R945 B.n769 B.n7 585
R946 B.n952 B.n7 585
R947 B.n768 B.n6 585
R948 B.n953 B.n6 585
R949 B.n767 B.n5 585
R950 B.n954 B.n5 585
R951 B.n766 B.n765 585
R952 B.n765 B.n4 585
R953 B.n764 B.n296 585
R954 B.n764 B.n763 585
R955 B.n754 B.n297 585
R956 B.n298 B.n297 585
R957 B.n756 B.n755 585
R958 B.n757 B.n756 585
R959 B.n753 B.n303 585
R960 B.n303 B.n302 585
R961 B.n752 B.n751 585
R962 B.n751 B.n750 585
R963 B.n305 B.n304 585
R964 B.n306 B.n305 585
R965 B.n743 B.n742 585
R966 B.n744 B.n743 585
R967 B.n741 B.n311 585
R968 B.n311 B.n310 585
R969 B.n740 B.n739 585
R970 B.n739 B.n738 585
R971 B.n313 B.n312 585
R972 B.n314 B.n313 585
R973 B.n731 B.n730 585
R974 B.n732 B.n731 585
R975 B.n729 B.n319 585
R976 B.n319 B.n318 585
R977 B.n728 B.n727 585
R978 B.n727 B.n726 585
R979 B.n321 B.n320 585
R980 B.n322 B.n321 585
R981 B.n719 B.n718 585
R982 B.n720 B.n719 585
R983 B.n717 B.n327 585
R984 B.n327 B.n326 585
R985 B.n716 B.n715 585
R986 B.n715 B.n714 585
R987 B.n329 B.n328 585
R988 B.n330 B.n329 585
R989 B.n707 B.n706 585
R990 B.n708 B.n707 585
R991 B.n705 B.n335 585
R992 B.n335 B.n334 585
R993 B.n704 B.n703 585
R994 B.n703 B.n702 585
R995 B.n337 B.n336 585
R996 B.n338 B.n337 585
R997 B.n695 B.n694 585
R998 B.n696 B.n695 585
R999 B.n693 B.n342 585
R1000 B.n346 B.n342 585
R1001 B.n692 B.n691 585
R1002 B.n691 B.n690 585
R1003 B.n344 B.n343 585
R1004 B.n345 B.n344 585
R1005 B.n683 B.n682 585
R1006 B.n684 B.n683 585
R1007 B.n681 B.n351 585
R1008 B.n351 B.n350 585
R1009 B.n680 B.n679 585
R1010 B.n679 B.n678 585
R1011 B.n353 B.n352 585
R1012 B.n354 B.n353 585
R1013 B.n671 B.n670 585
R1014 B.n672 B.n671 585
R1015 B.n669 B.n359 585
R1016 B.n359 B.n358 585
R1017 B.n668 B.n667 585
R1018 B.n667 B.n666 585
R1019 B.n361 B.n360 585
R1020 B.n659 B.n361 585
R1021 B.n658 B.n657 585
R1022 B.n660 B.n658 585
R1023 B.n656 B.n366 585
R1024 B.n366 B.n365 585
R1025 B.n655 B.n654 585
R1026 B.n654 B.n653 585
R1027 B.n368 B.n367 585
R1028 B.n369 B.n368 585
R1029 B.n646 B.n645 585
R1030 B.n647 B.n646 585
R1031 B.n644 B.n374 585
R1032 B.n374 B.n373 585
R1033 B.n643 B.n642 585
R1034 B.n642 B.n641 585
R1035 B.n376 B.n375 585
R1036 B.n377 B.n376 585
R1037 B.n634 B.n633 585
R1038 B.n635 B.n634 585
R1039 B.n632 B.n382 585
R1040 B.n382 B.n381 585
R1041 B.n631 B.n630 585
R1042 B.n630 B.n629 585
R1043 B.n384 B.n383 585
R1044 B.n622 B.n384 585
R1045 B.n621 B.n620 585
R1046 B.n623 B.n621 585
R1047 B.n619 B.n389 585
R1048 B.n389 B.n388 585
R1049 B.n618 B.n617 585
R1050 B.n617 B.n616 585
R1051 B.n391 B.n390 585
R1052 B.n392 B.n391 585
R1053 B.n609 B.n608 585
R1054 B.n610 B.n609 585
R1055 B.n607 B.n397 585
R1056 B.n397 B.n396 585
R1057 B.n606 B.n605 585
R1058 B.n605 B.n604 585
R1059 B.n399 B.n398 585
R1060 B.n400 B.n399 585
R1061 B.n600 B.n599 585
R1062 B.n403 B.n402 585
R1063 B.n596 B.n595 585
R1064 B.n597 B.n596 585
R1065 B.n594 B.n441 585
R1066 B.n593 B.n592 585
R1067 B.n591 B.n590 585
R1068 B.n589 B.n588 585
R1069 B.n587 B.n586 585
R1070 B.n585 B.n584 585
R1071 B.n583 B.n582 585
R1072 B.n581 B.n580 585
R1073 B.n579 B.n578 585
R1074 B.n577 B.n576 585
R1075 B.n575 B.n574 585
R1076 B.n573 B.n572 585
R1077 B.n571 B.n570 585
R1078 B.n569 B.n568 585
R1079 B.n567 B.n566 585
R1080 B.n565 B.n564 585
R1081 B.n563 B.n562 585
R1082 B.n561 B.n560 585
R1083 B.n559 B.n558 585
R1084 B.n557 B.n556 585
R1085 B.n555 B.n554 585
R1086 B.n553 B.n552 585
R1087 B.n551 B.n550 585
R1088 B.n549 B.n548 585
R1089 B.n547 B.n546 585
R1090 B.n545 B.n544 585
R1091 B.n543 B.n542 585
R1092 B.n541 B.n540 585
R1093 B.n539 B.n538 585
R1094 B.n537 B.n536 585
R1095 B.n535 B.n534 585
R1096 B.n532 B.n531 585
R1097 B.n530 B.n529 585
R1098 B.n528 B.n527 585
R1099 B.n526 B.n525 585
R1100 B.n524 B.n523 585
R1101 B.n522 B.n521 585
R1102 B.n520 B.n519 585
R1103 B.n518 B.n517 585
R1104 B.n516 B.n515 585
R1105 B.n514 B.n513 585
R1106 B.n512 B.n511 585
R1107 B.n510 B.n509 585
R1108 B.n508 B.n507 585
R1109 B.n506 B.n505 585
R1110 B.n504 B.n503 585
R1111 B.n502 B.n501 585
R1112 B.n500 B.n499 585
R1113 B.n498 B.n497 585
R1114 B.n496 B.n495 585
R1115 B.n494 B.n493 585
R1116 B.n492 B.n491 585
R1117 B.n490 B.n489 585
R1118 B.n488 B.n487 585
R1119 B.n486 B.n485 585
R1120 B.n484 B.n483 585
R1121 B.n482 B.n481 585
R1122 B.n480 B.n479 585
R1123 B.n478 B.n477 585
R1124 B.n476 B.n475 585
R1125 B.n474 B.n473 585
R1126 B.n472 B.n471 585
R1127 B.n470 B.n469 585
R1128 B.n468 B.n467 585
R1129 B.n466 B.n465 585
R1130 B.n464 B.n463 585
R1131 B.n462 B.n461 585
R1132 B.n460 B.n459 585
R1133 B.n458 B.n457 585
R1134 B.n456 B.n455 585
R1135 B.n454 B.n453 585
R1136 B.n452 B.n451 585
R1137 B.n450 B.n449 585
R1138 B.n448 B.n447 585
R1139 B.n601 B.n401 585
R1140 B.n401 B.n400 585
R1141 B.n603 B.n602 585
R1142 B.n604 B.n603 585
R1143 B.n395 B.n394 585
R1144 B.n396 B.n395 585
R1145 B.n612 B.n611 585
R1146 B.n611 B.n610 585
R1147 B.n613 B.n393 585
R1148 B.n393 B.n392 585
R1149 B.n615 B.n614 585
R1150 B.n616 B.n615 585
R1151 B.n387 B.n386 585
R1152 B.n388 B.n387 585
R1153 B.n625 B.n624 585
R1154 B.n624 B.n623 585
R1155 B.n626 B.n385 585
R1156 B.n622 B.n385 585
R1157 B.n628 B.n627 585
R1158 B.n629 B.n628 585
R1159 B.n380 B.n379 585
R1160 B.n381 B.n380 585
R1161 B.n637 B.n636 585
R1162 B.n636 B.n635 585
R1163 B.n638 B.n378 585
R1164 B.n378 B.n377 585
R1165 B.n640 B.n639 585
R1166 B.n641 B.n640 585
R1167 B.n372 B.n371 585
R1168 B.n373 B.n372 585
R1169 B.n649 B.n648 585
R1170 B.n648 B.n647 585
R1171 B.n650 B.n370 585
R1172 B.n370 B.n369 585
R1173 B.n652 B.n651 585
R1174 B.n653 B.n652 585
R1175 B.n364 B.n363 585
R1176 B.n365 B.n364 585
R1177 B.n662 B.n661 585
R1178 B.n661 B.n660 585
R1179 B.n663 B.n362 585
R1180 B.n659 B.n362 585
R1181 B.n665 B.n664 585
R1182 B.n666 B.n665 585
R1183 B.n357 B.n356 585
R1184 B.n358 B.n357 585
R1185 B.n674 B.n673 585
R1186 B.n673 B.n672 585
R1187 B.n675 B.n355 585
R1188 B.n355 B.n354 585
R1189 B.n677 B.n676 585
R1190 B.n678 B.n677 585
R1191 B.n349 B.n348 585
R1192 B.n350 B.n349 585
R1193 B.n686 B.n685 585
R1194 B.n685 B.n684 585
R1195 B.n687 B.n347 585
R1196 B.n347 B.n345 585
R1197 B.n689 B.n688 585
R1198 B.n690 B.n689 585
R1199 B.n341 B.n340 585
R1200 B.n346 B.n341 585
R1201 B.n698 B.n697 585
R1202 B.n697 B.n696 585
R1203 B.n699 B.n339 585
R1204 B.n339 B.n338 585
R1205 B.n701 B.n700 585
R1206 B.n702 B.n701 585
R1207 B.n333 B.n332 585
R1208 B.n334 B.n333 585
R1209 B.n710 B.n709 585
R1210 B.n709 B.n708 585
R1211 B.n711 B.n331 585
R1212 B.n331 B.n330 585
R1213 B.n713 B.n712 585
R1214 B.n714 B.n713 585
R1215 B.n325 B.n324 585
R1216 B.n326 B.n325 585
R1217 B.n722 B.n721 585
R1218 B.n721 B.n720 585
R1219 B.n723 B.n323 585
R1220 B.n323 B.n322 585
R1221 B.n725 B.n724 585
R1222 B.n726 B.n725 585
R1223 B.n317 B.n316 585
R1224 B.n318 B.n317 585
R1225 B.n734 B.n733 585
R1226 B.n733 B.n732 585
R1227 B.n735 B.n315 585
R1228 B.n315 B.n314 585
R1229 B.n737 B.n736 585
R1230 B.n738 B.n737 585
R1231 B.n309 B.n308 585
R1232 B.n310 B.n309 585
R1233 B.n746 B.n745 585
R1234 B.n745 B.n744 585
R1235 B.n747 B.n307 585
R1236 B.n307 B.n306 585
R1237 B.n749 B.n748 585
R1238 B.n750 B.n749 585
R1239 B.n301 B.n300 585
R1240 B.n302 B.n301 585
R1241 B.n759 B.n758 585
R1242 B.n758 B.n757 585
R1243 B.n760 B.n299 585
R1244 B.n299 B.n298 585
R1245 B.n762 B.n761 585
R1246 B.n763 B.n762 585
R1247 B.n3 B.n0 585
R1248 B.n4 B.n3 585
R1249 B.n951 B.n1 585
R1250 B.n952 B.n951 585
R1251 B.n950 B.n949 585
R1252 B.n950 B.n8 585
R1253 B.n948 B.n9 585
R1254 B.n12 B.n9 585
R1255 B.n947 B.n946 585
R1256 B.n946 B.n945 585
R1257 B.n11 B.n10 585
R1258 B.n944 B.n11 585
R1259 B.n942 B.n941 585
R1260 B.n943 B.n942 585
R1261 B.n940 B.n17 585
R1262 B.n17 B.n16 585
R1263 B.n939 B.n938 585
R1264 B.n938 B.n937 585
R1265 B.n19 B.n18 585
R1266 B.n936 B.n19 585
R1267 B.n934 B.n933 585
R1268 B.n935 B.n934 585
R1269 B.n932 B.n24 585
R1270 B.n24 B.n23 585
R1271 B.n931 B.n930 585
R1272 B.n930 B.n929 585
R1273 B.n26 B.n25 585
R1274 B.n928 B.n26 585
R1275 B.n926 B.n925 585
R1276 B.n927 B.n926 585
R1277 B.n924 B.n31 585
R1278 B.n31 B.n30 585
R1279 B.n923 B.n922 585
R1280 B.n922 B.n921 585
R1281 B.n33 B.n32 585
R1282 B.n920 B.n33 585
R1283 B.n918 B.n917 585
R1284 B.n919 B.n918 585
R1285 B.n916 B.n38 585
R1286 B.n38 B.n37 585
R1287 B.n915 B.n914 585
R1288 B.n914 B.n913 585
R1289 B.n40 B.n39 585
R1290 B.n912 B.n40 585
R1291 B.n910 B.n909 585
R1292 B.n911 B.n910 585
R1293 B.n908 B.n45 585
R1294 B.n45 B.n44 585
R1295 B.n907 B.n906 585
R1296 B.n906 B.n905 585
R1297 B.n47 B.n46 585
R1298 B.n904 B.n47 585
R1299 B.n902 B.n901 585
R1300 B.n903 B.n902 585
R1301 B.n900 B.n52 585
R1302 B.n52 B.n51 585
R1303 B.n899 B.n898 585
R1304 B.n898 B.n897 585
R1305 B.n54 B.n53 585
R1306 B.n896 B.n54 585
R1307 B.n894 B.n893 585
R1308 B.n895 B.n894 585
R1309 B.n892 B.n59 585
R1310 B.n59 B.n58 585
R1311 B.n891 B.n890 585
R1312 B.n890 B.n889 585
R1313 B.n61 B.n60 585
R1314 B.n888 B.n61 585
R1315 B.n886 B.n885 585
R1316 B.n887 B.n886 585
R1317 B.n884 B.n65 585
R1318 B.n68 B.n65 585
R1319 B.n883 B.n882 585
R1320 B.n882 B.n881 585
R1321 B.n67 B.n66 585
R1322 B.n880 B.n67 585
R1323 B.n878 B.n877 585
R1324 B.n879 B.n878 585
R1325 B.n876 B.n73 585
R1326 B.n73 B.n72 585
R1327 B.n875 B.n874 585
R1328 B.n874 B.n873 585
R1329 B.n75 B.n74 585
R1330 B.n872 B.n75 585
R1331 B.n870 B.n869 585
R1332 B.n871 B.n870 585
R1333 B.n868 B.n80 585
R1334 B.n80 B.n79 585
R1335 B.n867 B.n866 585
R1336 B.n866 B.n865 585
R1337 B.n82 B.n81 585
R1338 B.n864 B.n82 585
R1339 B.n862 B.n861 585
R1340 B.n863 B.n862 585
R1341 B.n860 B.n86 585
R1342 B.n89 B.n86 585
R1343 B.n859 B.n858 585
R1344 B.n858 B.n857 585
R1345 B.n88 B.n87 585
R1346 B.n856 B.n88 585
R1347 B.n854 B.n853 585
R1348 B.n855 B.n854 585
R1349 B.n852 B.n94 585
R1350 B.n94 B.n93 585
R1351 B.n851 B.n850 585
R1352 B.n850 B.n849 585
R1353 B.n96 B.n95 585
R1354 B.n848 B.n96 585
R1355 B.n846 B.n845 585
R1356 B.n847 B.n846 585
R1357 B.n844 B.n101 585
R1358 B.n101 B.n100 585
R1359 B.n955 B.n954 585
R1360 B.n953 B.n2 585
R1361 B.n842 B.n101 506.916
R1362 B.n839 B.n142 506.916
R1363 B.n447 B.n399 506.916
R1364 B.n599 B.n401 506.916
R1365 B.n143 B.t10 299.548
R1366 B.n444 B.t18 299.548
R1367 B.n145 B.t20 299.548
R1368 B.n442 B.t15 299.548
R1369 B.n145 B.t19 287.01
R1370 B.n143 B.t8 287.01
R1371 B.n444 B.t16 287.01
R1372 B.n442 B.t12 287.01
R1373 B.n840 B.n140 256.663
R1374 B.n840 B.n139 256.663
R1375 B.n840 B.n138 256.663
R1376 B.n840 B.n137 256.663
R1377 B.n840 B.n136 256.663
R1378 B.n840 B.n135 256.663
R1379 B.n840 B.n134 256.663
R1380 B.n840 B.n133 256.663
R1381 B.n840 B.n132 256.663
R1382 B.n840 B.n131 256.663
R1383 B.n840 B.n130 256.663
R1384 B.n840 B.n129 256.663
R1385 B.n840 B.n128 256.663
R1386 B.n840 B.n127 256.663
R1387 B.n840 B.n126 256.663
R1388 B.n840 B.n125 256.663
R1389 B.n840 B.n124 256.663
R1390 B.n840 B.n123 256.663
R1391 B.n840 B.n122 256.663
R1392 B.n840 B.n121 256.663
R1393 B.n840 B.n120 256.663
R1394 B.n840 B.n119 256.663
R1395 B.n840 B.n118 256.663
R1396 B.n840 B.n117 256.663
R1397 B.n840 B.n116 256.663
R1398 B.n840 B.n115 256.663
R1399 B.n840 B.n114 256.663
R1400 B.n840 B.n113 256.663
R1401 B.n840 B.n112 256.663
R1402 B.n840 B.n111 256.663
R1403 B.n840 B.n110 256.663
R1404 B.n840 B.n109 256.663
R1405 B.n840 B.n108 256.663
R1406 B.n840 B.n107 256.663
R1407 B.n840 B.n106 256.663
R1408 B.n840 B.n105 256.663
R1409 B.n840 B.n104 256.663
R1410 B.n841 B.n840 256.663
R1411 B.n598 B.n597 256.663
R1412 B.n597 B.n404 256.663
R1413 B.n597 B.n405 256.663
R1414 B.n597 B.n406 256.663
R1415 B.n597 B.n407 256.663
R1416 B.n597 B.n408 256.663
R1417 B.n597 B.n409 256.663
R1418 B.n597 B.n410 256.663
R1419 B.n597 B.n411 256.663
R1420 B.n597 B.n412 256.663
R1421 B.n597 B.n413 256.663
R1422 B.n597 B.n414 256.663
R1423 B.n597 B.n415 256.663
R1424 B.n597 B.n416 256.663
R1425 B.n597 B.n417 256.663
R1426 B.n597 B.n418 256.663
R1427 B.n597 B.n419 256.663
R1428 B.n597 B.n420 256.663
R1429 B.n597 B.n421 256.663
R1430 B.n597 B.n422 256.663
R1431 B.n597 B.n423 256.663
R1432 B.n597 B.n424 256.663
R1433 B.n597 B.n425 256.663
R1434 B.n597 B.n426 256.663
R1435 B.n597 B.n427 256.663
R1436 B.n597 B.n428 256.663
R1437 B.n597 B.n429 256.663
R1438 B.n597 B.n430 256.663
R1439 B.n597 B.n431 256.663
R1440 B.n597 B.n432 256.663
R1441 B.n597 B.n433 256.663
R1442 B.n597 B.n434 256.663
R1443 B.n597 B.n435 256.663
R1444 B.n597 B.n436 256.663
R1445 B.n597 B.n437 256.663
R1446 B.n597 B.n438 256.663
R1447 B.n597 B.n439 256.663
R1448 B.n597 B.n440 256.663
R1449 B.n957 B.n956 256.663
R1450 B.n144 B.t11 237.293
R1451 B.n445 B.t17 237.293
R1452 B.n146 B.t21 237.292
R1453 B.n443 B.t14 237.292
R1454 B.n148 B.n103 163.367
R1455 B.n152 B.n151 163.367
R1456 B.n156 B.n155 163.367
R1457 B.n160 B.n159 163.367
R1458 B.n164 B.n163 163.367
R1459 B.n168 B.n167 163.367
R1460 B.n172 B.n171 163.367
R1461 B.n176 B.n175 163.367
R1462 B.n180 B.n179 163.367
R1463 B.n184 B.n183 163.367
R1464 B.n188 B.n187 163.367
R1465 B.n192 B.n191 163.367
R1466 B.n196 B.n195 163.367
R1467 B.n200 B.n199 163.367
R1468 B.n204 B.n203 163.367
R1469 B.n208 B.n207 163.367
R1470 B.n212 B.n211 163.367
R1471 B.n216 B.n215 163.367
R1472 B.n220 B.n219 163.367
R1473 B.n224 B.n223 163.367
R1474 B.n228 B.n227 163.367
R1475 B.n233 B.n232 163.367
R1476 B.n237 B.n236 163.367
R1477 B.n241 B.n240 163.367
R1478 B.n245 B.n244 163.367
R1479 B.n249 B.n248 163.367
R1480 B.n253 B.n252 163.367
R1481 B.n257 B.n256 163.367
R1482 B.n261 B.n260 163.367
R1483 B.n265 B.n264 163.367
R1484 B.n269 B.n268 163.367
R1485 B.n273 B.n272 163.367
R1486 B.n277 B.n276 163.367
R1487 B.n281 B.n280 163.367
R1488 B.n285 B.n284 163.367
R1489 B.n289 B.n288 163.367
R1490 B.n293 B.n292 163.367
R1491 B.n839 B.n141 163.367
R1492 B.n605 B.n399 163.367
R1493 B.n605 B.n397 163.367
R1494 B.n609 B.n397 163.367
R1495 B.n609 B.n391 163.367
R1496 B.n617 B.n391 163.367
R1497 B.n617 B.n389 163.367
R1498 B.n621 B.n389 163.367
R1499 B.n621 B.n384 163.367
R1500 B.n630 B.n384 163.367
R1501 B.n630 B.n382 163.367
R1502 B.n634 B.n382 163.367
R1503 B.n634 B.n376 163.367
R1504 B.n642 B.n376 163.367
R1505 B.n642 B.n374 163.367
R1506 B.n646 B.n374 163.367
R1507 B.n646 B.n368 163.367
R1508 B.n654 B.n368 163.367
R1509 B.n654 B.n366 163.367
R1510 B.n658 B.n366 163.367
R1511 B.n658 B.n361 163.367
R1512 B.n667 B.n361 163.367
R1513 B.n667 B.n359 163.367
R1514 B.n671 B.n359 163.367
R1515 B.n671 B.n353 163.367
R1516 B.n679 B.n353 163.367
R1517 B.n679 B.n351 163.367
R1518 B.n683 B.n351 163.367
R1519 B.n683 B.n344 163.367
R1520 B.n691 B.n344 163.367
R1521 B.n691 B.n342 163.367
R1522 B.n695 B.n342 163.367
R1523 B.n695 B.n337 163.367
R1524 B.n703 B.n337 163.367
R1525 B.n703 B.n335 163.367
R1526 B.n707 B.n335 163.367
R1527 B.n707 B.n329 163.367
R1528 B.n715 B.n329 163.367
R1529 B.n715 B.n327 163.367
R1530 B.n719 B.n327 163.367
R1531 B.n719 B.n321 163.367
R1532 B.n727 B.n321 163.367
R1533 B.n727 B.n319 163.367
R1534 B.n731 B.n319 163.367
R1535 B.n731 B.n313 163.367
R1536 B.n739 B.n313 163.367
R1537 B.n739 B.n311 163.367
R1538 B.n743 B.n311 163.367
R1539 B.n743 B.n305 163.367
R1540 B.n751 B.n305 163.367
R1541 B.n751 B.n303 163.367
R1542 B.n756 B.n303 163.367
R1543 B.n756 B.n297 163.367
R1544 B.n764 B.n297 163.367
R1545 B.n765 B.n764 163.367
R1546 B.n765 B.n5 163.367
R1547 B.n6 B.n5 163.367
R1548 B.n7 B.n6 163.367
R1549 B.n771 B.n7 163.367
R1550 B.n772 B.n771 163.367
R1551 B.n772 B.n13 163.367
R1552 B.n14 B.n13 163.367
R1553 B.n15 B.n14 163.367
R1554 B.n777 B.n15 163.367
R1555 B.n777 B.n20 163.367
R1556 B.n21 B.n20 163.367
R1557 B.n22 B.n21 163.367
R1558 B.n782 B.n22 163.367
R1559 B.n782 B.n27 163.367
R1560 B.n28 B.n27 163.367
R1561 B.n29 B.n28 163.367
R1562 B.n787 B.n29 163.367
R1563 B.n787 B.n34 163.367
R1564 B.n35 B.n34 163.367
R1565 B.n36 B.n35 163.367
R1566 B.n792 B.n36 163.367
R1567 B.n792 B.n41 163.367
R1568 B.n42 B.n41 163.367
R1569 B.n43 B.n42 163.367
R1570 B.n797 B.n43 163.367
R1571 B.n797 B.n48 163.367
R1572 B.n49 B.n48 163.367
R1573 B.n50 B.n49 163.367
R1574 B.n802 B.n50 163.367
R1575 B.n802 B.n55 163.367
R1576 B.n56 B.n55 163.367
R1577 B.n57 B.n56 163.367
R1578 B.n807 B.n57 163.367
R1579 B.n807 B.n62 163.367
R1580 B.n63 B.n62 163.367
R1581 B.n64 B.n63 163.367
R1582 B.n812 B.n64 163.367
R1583 B.n812 B.n69 163.367
R1584 B.n70 B.n69 163.367
R1585 B.n71 B.n70 163.367
R1586 B.n817 B.n71 163.367
R1587 B.n817 B.n76 163.367
R1588 B.n77 B.n76 163.367
R1589 B.n78 B.n77 163.367
R1590 B.n822 B.n78 163.367
R1591 B.n822 B.n83 163.367
R1592 B.n84 B.n83 163.367
R1593 B.n85 B.n84 163.367
R1594 B.n827 B.n85 163.367
R1595 B.n827 B.n90 163.367
R1596 B.n91 B.n90 163.367
R1597 B.n92 B.n91 163.367
R1598 B.n832 B.n92 163.367
R1599 B.n832 B.n97 163.367
R1600 B.n98 B.n97 163.367
R1601 B.n99 B.n98 163.367
R1602 B.n142 B.n99 163.367
R1603 B.n596 B.n403 163.367
R1604 B.n596 B.n441 163.367
R1605 B.n592 B.n591 163.367
R1606 B.n588 B.n587 163.367
R1607 B.n584 B.n583 163.367
R1608 B.n580 B.n579 163.367
R1609 B.n576 B.n575 163.367
R1610 B.n572 B.n571 163.367
R1611 B.n568 B.n567 163.367
R1612 B.n564 B.n563 163.367
R1613 B.n560 B.n559 163.367
R1614 B.n556 B.n555 163.367
R1615 B.n552 B.n551 163.367
R1616 B.n548 B.n547 163.367
R1617 B.n544 B.n543 163.367
R1618 B.n540 B.n539 163.367
R1619 B.n536 B.n535 163.367
R1620 B.n531 B.n530 163.367
R1621 B.n527 B.n526 163.367
R1622 B.n523 B.n522 163.367
R1623 B.n519 B.n518 163.367
R1624 B.n515 B.n514 163.367
R1625 B.n511 B.n510 163.367
R1626 B.n507 B.n506 163.367
R1627 B.n503 B.n502 163.367
R1628 B.n499 B.n498 163.367
R1629 B.n495 B.n494 163.367
R1630 B.n491 B.n490 163.367
R1631 B.n487 B.n486 163.367
R1632 B.n483 B.n482 163.367
R1633 B.n479 B.n478 163.367
R1634 B.n475 B.n474 163.367
R1635 B.n471 B.n470 163.367
R1636 B.n467 B.n466 163.367
R1637 B.n463 B.n462 163.367
R1638 B.n459 B.n458 163.367
R1639 B.n455 B.n454 163.367
R1640 B.n451 B.n450 163.367
R1641 B.n603 B.n401 163.367
R1642 B.n603 B.n395 163.367
R1643 B.n611 B.n395 163.367
R1644 B.n611 B.n393 163.367
R1645 B.n615 B.n393 163.367
R1646 B.n615 B.n387 163.367
R1647 B.n624 B.n387 163.367
R1648 B.n624 B.n385 163.367
R1649 B.n628 B.n385 163.367
R1650 B.n628 B.n380 163.367
R1651 B.n636 B.n380 163.367
R1652 B.n636 B.n378 163.367
R1653 B.n640 B.n378 163.367
R1654 B.n640 B.n372 163.367
R1655 B.n648 B.n372 163.367
R1656 B.n648 B.n370 163.367
R1657 B.n652 B.n370 163.367
R1658 B.n652 B.n364 163.367
R1659 B.n661 B.n364 163.367
R1660 B.n661 B.n362 163.367
R1661 B.n665 B.n362 163.367
R1662 B.n665 B.n357 163.367
R1663 B.n673 B.n357 163.367
R1664 B.n673 B.n355 163.367
R1665 B.n677 B.n355 163.367
R1666 B.n677 B.n349 163.367
R1667 B.n685 B.n349 163.367
R1668 B.n685 B.n347 163.367
R1669 B.n689 B.n347 163.367
R1670 B.n689 B.n341 163.367
R1671 B.n697 B.n341 163.367
R1672 B.n697 B.n339 163.367
R1673 B.n701 B.n339 163.367
R1674 B.n701 B.n333 163.367
R1675 B.n709 B.n333 163.367
R1676 B.n709 B.n331 163.367
R1677 B.n713 B.n331 163.367
R1678 B.n713 B.n325 163.367
R1679 B.n721 B.n325 163.367
R1680 B.n721 B.n323 163.367
R1681 B.n725 B.n323 163.367
R1682 B.n725 B.n317 163.367
R1683 B.n733 B.n317 163.367
R1684 B.n733 B.n315 163.367
R1685 B.n737 B.n315 163.367
R1686 B.n737 B.n309 163.367
R1687 B.n745 B.n309 163.367
R1688 B.n745 B.n307 163.367
R1689 B.n749 B.n307 163.367
R1690 B.n749 B.n301 163.367
R1691 B.n758 B.n301 163.367
R1692 B.n758 B.n299 163.367
R1693 B.n762 B.n299 163.367
R1694 B.n762 B.n3 163.367
R1695 B.n955 B.n3 163.367
R1696 B.n951 B.n2 163.367
R1697 B.n951 B.n950 163.367
R1698 B.n950 B.n9 163.367
R1699 B.n946 B.n9 163.367
R1700 B.n946 B.n11 163.367
R1701 B.n942 B.n11 163.367
R1702 B.n942 B.n17 163.367
R1703 B.n938 B.n17 163.367
R1704 B.n938 B.n19 163.367
R1705 B.n934 B.n19 163.367
R1706 B.n934 B.n24 163.367
R1707 B.n930 B.n24 163.367
R1708 B.n930 B.n26 163.367
R1709 B.n926 B.n26 163.367
R1710 B.n926 B.n31 163.367
R1711 B.n922 B.n31 163.367
R1712 B.n922 B.n33 163.367
R1713 B.n918 B.n33 163.367
R1714 B.n918 B.n38 163.367
R1715 B.n914 B.n38 163.367
R1716 B.n914 B.n40 163.367
R1717 B.n910 B.n40 163.367
R1718 B.n910 B.n45 163.367
R1719 B.n906 B.n45 163.367
R1720 B.n906 B.n47 163.367
R1721 B.n902 B.n47 163.367
R1722 B.n902 B.n52 163.367
R1723 B.n898 B.n52 163.367
R1724 B.n898 B.n54 163.367
R1725 B.n894 B.n54 163.367
R1726 B.n894 B.n59 163.367
R1727 B.n890 B.n59 163.367
R1728 B.n890 B.n61 163.367
R1729 B.n886 B.n61 163.367
R1730 B.n886 B.n65 163.367
R1731 B.n882 B.n65 163.367
R1732 B.n882 B.n67 163.367
R1733 B.n878 B.n67 163.367
R1734 B.n878 B.n73 163.367
R1735 B.n874 B.n73 163.367
R1736 B.n874 B.n75 163.367
R1737 B.n870 B.n75 163.367
R1738 B.n870 B.n80 163.367
R1739 B.n866 B.n80 163.367
R1740 B.n866 B.n82 163.367
R1741 B.n862 B.n82 163.367
R1742 B.n862 B.n86 163.367
R1743 B.n858 B.n86 163.367
R1744 B.n858 B.n88 163.367
R1745 B.n854 B.n88 163.367
R1746 B.n854 B.n94 163.367
R1747 B.n850 B.n94 163.367
R1748 B.n850 B.n96 163.367
R1749 B.n846 B.n96 163.367
R1750 B.n846 B.n101 163.367
R1751 B.n597 B.n400 83.26
R1752 B.n840 B.n100 83.26
R1753 B.n842 B.n841 71.676
R1754 B.n148 B.n104 71.676
R1755 B.n152 B.n105 71.676
R1756 B.n156 B.n106 71.676
R1757 B.n160 B.n107 71.676
R1758 B.n164 B.n108 71.676
R1759 B.n168 B.n109 71.676
R1760 B.n172 B.n110 71.676
R1761 B.n176 B.n111 71.676
R1762 B.n180 B.n112 71.676
R1763 B.n184 B.n113 71.676
R1764 B.n188 B.n114 71.676
R1765 B.n192 B.n115 71.676
R1766 B.n196 B.n116 71.676
R1767 B.n200 B.n117 71.676
R1768 B.n204 B.n118 71.676
R1769 B.n208 B.n119 71.676
R1770 B.n212 B.n120 71.676
R1771 B.n216 B.n121 71.676
R1772 B.n220 B.n122 71.676
R1773 B.n224 B.n123 71.676
R1774 B.n228 B.n124 71.676
R1775 B.n233 B.n125 71.676
R1776 B.n237 B.n126 71.676
R1777 B.n241 B.n127 71.676
R1778 B.n245 B.n128 71.676
R1779 B.n249 B.n129 71.676
R1780 B.n253 B.n130 71.676
R1781 B.n257 B.n131 71.676
R1782 B.n261 B.n132 71.676
R1783 B.n265 B.n133 71.676
R1784 B.n269 B.n134 71.676
R1785 B.n273 B.n135 71.676
R1786 B.n277 B.n136 71.676
R1787 B.n281 B.n137 71.676
R1788 B.n285 B.n138 71.676
R1789 B.n289 B.n139 71.676
R1790 B.n293 B.n140 71.676
R1791 B.n141 B.n140 71.676
R1792 B.n292 B.n139 71.676
R1793 B.n288 B.n138 71.676
R1794 B.n284 B.n137 71.676
R1795 B.n280 B.n136 71.676
R1796 B.n276 B.n135 71.676
R1797 B.n272 B.n134 71.676
R1798 B.n268 B.n133 71.676
R1799 B.n264 B.n132 71.676
R1800 B.n260 B.n131 71.676
R1801 B.n256 B.n130 71.676
R1802 B.n252 B.n129 71.676
R1803 B.n248 B.n128 71.676
R1804 B.n244 B.n127 71.676
R1805 B.n240 B.n126 71.676
R1806 B.n236 B.n125 71.676
R1807 B.n232 B.n124 71.676
R1808 B.n227 B.n123 71.676
R1809 B.n223 B.n122 71.676
R1810 B.n219 B.n121 71.676
R1811 B.n215 B.n120 71.676
R1812 B.n211 B.n119 71.676
R1813 B.n207 B.n118 71.676
R1814 B.n203 B.n117 71.676
R1815 B.n199 B.n116 71.676
R1816 B.n195 B.n115 71.676
R1817 B.n191 B.n114 71.676
R1818 B.n187 B.n113 71.676
R1819 B.n183 B.n112 71.676
R1820 B.n179 B.n111 71.676
R1821 B.n175 B.n110 71.676
R1822 B.n171 B.n109 71.676
R1823 B.n167 B.n108 71.676
R1824 B.n163 B.n107 71.676
R1825 B.n159 B.n106 71.676
R1826 B.n155 B.n105 71.676
R1827 B.n151 B.n104 71.676
R1828 B.n841 B.n103 71.676
R1829 B.n599 B.n598 71.676
R1830 B.n441 B.n404 71.676
R1831 B.n591 B.n405 71.676
R1832 B.n587 B.n406 71.676
R1833 B.n583 B.n407 71.676
R1834 B.n579 B.n408 71.676
R1835 B.n575 B.n409 71.676
R1836 B.n571 B.n410 71.676
R1837 B.n567 B.n411 71.676
R1838 B.n563 B.n412 71.676
R1839 B.n559 B.n413 71.676
R1840 B.n555 B.n414 71.676
R1841 B.n551 B.n415 71.676
R1842 B.n547 B.n416 71.676
R1843 B.n543 B.n417 71.676
R1844 B.n539 B.n418 71.676
R1845 B.n535 B.n419 71.676
R1846 B.n530 B.n420 71.676
R1847 B.n526 B.n421 71.676
R1848 B.n522 B.n422 71.676
R1849 B.n518 B.n423 71.676
R1850 B.n514 B.n424 71.676
R1851 B.n510 B.n425 71.676
R1852 B.n506 B.n426 71.676
R1853 B.n502 B.n427 71.676
R1854 B.n498 B.n428 71.676
R1855 B.n494 B.n429 71.676
R1856 B.n490 B.n430 71.676
R1857 B.n486 B.n431 71.676
R1858 B.n482 B.n432 71.676
R1859 B.n478 B.n433 71.676
R1860 B.n474 B.n434 71.676
R1861 B.n470 B.n435 71.676
R1862 B.n466 B.n436 71.676
R1863 B.n462 B.n437 71.676
R1864 B.n458 B.n438 71.676
R1865 B.n454 B.n439 71.676
R1866 B.n450 B.n440 71.676
R1867 B.n598 B.n403 71.676
R1868 B.n592 B.n404 71.676
R1869 B.n588 B.n405 71.676
R1870 B.n584 B.n406 71.676
R1871 B.n580 B.n407 71.676
R1872 B.n576 B.n408 71.676
R1873 B.n572 B.n409 71.676
R1874 B.n568 B.n410 71.676
R1875 B.n564 B.n411 71.676
R1876 B.n560 B.n412 71.676
R1877 B.n556 B.n413 71.676
R1878 B.n552 B.n414 71.676
R1879 B.n548 B.n415 71.676
R1880 B.n544 B.n416 71.676
R1881 B.n540 B.n417 71.676
R1882 B.n536 B.n418 71.676
R1883 B.n531 B.n419 71.676
R1884 B.n527 B.n420 71.676
R1885 B.n523 B.n421 71.676
R1886 B.n519 B.n422 71.676
R1887 B.n515 B.n423 71.676
R1888 B.n511 B.n424 71.676
R1889 B.n507 B.n425 71.676
R1890 B.n503 B.n426 71.676
R1891 B.n499 B.n427 71.676
R1892 B.n495 B.n428 71.676
R1893 B.n491 B.n429 71.676
R1894 B.n487 B.n430 71.676
R1895 B.n483 B.n431 71.676
R1896 B.n479 B.n432 71.676
R1897 B.n475 B.n433 71.676
R1898 B.n471 B.n434 71.676
R1899 B.n467 B.n435 71.676
R1900 B.n463 B.n436 71.676
R1901 B.n459 B.n437 71.676
R1902 B.n455 B.n438 71.676
R1903 B.n451 B.n439 71.676
R1904 B.n447 B.n440 71.676
R1905 B.n956 B.n955 71.676
R1906 B.n956 B.n2 71.676
R1907 B.n146 B.n145 62.255
R1908 B.n144 B.n143 62.255
R1909 B.n445 B.n444 62.255
R1910 B.n443 B.n442 62.255
R1911 B.n147 B.n146 59.5399
R1912 B.n230 B.n144 59.5399
R1913 B.n446 B.n445 59.5399
R1914 B.n533 B.n443 59.5399
R1915 B.n604 B.n400 51.0063
R1916 B.n604 B.n396 51.0063
R1917 B.n610 B.n396 51.0063
R1918 B.n610 B.n392 51.0063
R1919 B.n616 B.n392 51.0063
R1920 B.n616 B.n388 51.0063
R1921 B.n623 B.n388 51.0063
R1922 B.n623 B.n622 51.0063
R1923 B.n629 B.n381 51.0063
R1924 B.n635 B.n381 51.0063
R1925 B.n635 B.n377 51.0063
R1926 B.n641 B.n377 51.0063
R1927 B.n641 B.n373 51.0063
R1928 B.n647 B.n373 51.0063
R1929 B.n647 B.n369 51.0063
R1930 B.n653 B.n369 51.0063
R1931 B.n653 B.n365 51.0063
R1932 B.n660 B.n365 51.0063
R1933 B.n660 B.n659 51.0063
R1934 B.n666 B.n358 51.0063
R1935 B.n672 B.n358 51.0063
R1936 B.n672 B.n354 51.0063
R1937 B.n678 B.n354 51.0063
R1938 B.n678 B.n350 51.0063
R1939 B.n684 B.n350 51.0063
R1940 B.n684 B.n345 51.0063
R1941 B.n690 B.n345 51.0063
R1942 B.n690 B.n346 51.0063
R1943 B.n696 B.n338 51.0063
R1944 B.n702 B.n338 51.0063
R1945 B.n702 B.n334 51.0063
R1946 B.n708 B.n334 51.0063
R1947 B.n708 B.n330 51.0063
R1948 B.n714 B.n330 51.0063
R1949 B.n714 B.n326 51.0063
R1950 B.n720 B.n326 51.0063
R1951 B.n726 B.n322 51.0063
R1952 B.n726 B.n318 51.0063
R1953 B.n732 B.n318 51.0063
R1954 B.n732 B.n314 51.0063
R1955 B.n738 B.n314 51.0063
R1956 B.n738 B.n310 51.0063
R1957 B.n744 B.n310 51.0063
R1958 B.n744 B.n306 51.0063
R1959 B.n750 B.n306 51.0063
R1960 B.n757 B.n302 51.0063
R1961 B.n757 B.n298 51.0063
R1962 B.n763 B.n298 51.0063
R1963 B.n763 B.n4 51.0063
R1964 B.n954 B.n4 51.0063
R1965 B.n954 B.n953 51.0063
R1966 B.n953 B.n952 51.0063
R1967 B.n952 B.n8 51.0063
R1968 B.n12 B.n8 51.0063
R1969 B.n945 B.n12 51.0063
R1970 B.n945 B.n944 51.0063
R1971 B.n943 B.n16 51.0063
R1972 B.n937 B.n16 51.0063
R1973 B.n937 B.n936 51.0063
R1974 B.n936 B.n935 51.0063
R1975 B.n935 B.n23 51.0063
R1976 B.n929 B.n23 51.0063
R1977 B.n929 B.n928 51.0063
R1978 B.n928 B.n927 51.0063
R1979 B.n927 B.n30 51.0063
R1980 B.n921 B.n920 51.0063
R1981 B.n920 B.n919 51.0063
R1982 B.n919 B.n37 51.0063
R1983 B.n913 B.n37 51.0063
R1984 B.n913 B.n912 51.0063
R1985 B.n912 B.n911 51.0063
R1986 B.n911 B.n44 51.0063
R1987 B.n905 B.n44 51.0063
R1988 B.n904 B.n903 51.0063
R1989 B.n903 B.n51 51.0063
R1990 B.n897 B.n51 51.0063
R1991 B.n897 B.n896 51.0063
R1992 B.n896 B.n895 51.0063
R1993 B.n895 B.n58 51.0063
R1994 B.n889 B.n58 51.0063
R1995 B.n889 B.n888 51.0063
R1996 B.n888 B.n887 51.0063
R1997 B.n881 B.n68 51.0063
R1998 B.n881 B.n880 51.0063
R1999 B.n880 B.n879 51.0063
R2000 B.n879 B.n72 51.0063
R2001 B.n873 B.n72 51.0063
R2002 B.n873 B.n872 51.0063
R2003 B.n872 B.n871 51.0063
R2004 B.n871 B.n79 51.0063
R2005 B.n865 B.n79 51.0063
R2006 B.n865 B.n864 51.0063
R2007 B.n864 B.n863 51.0063
R2008 B.n857 B.n89 51.0063
R2009 B.n857 B.n856 51.0063
R2010 B.n856 B.n855 51.0063
R2011 B.n855 B.n93 51.0063
R2012 B.n849 B.n93 51.0063
R2013 B.n849 B.n848 51.0063
R2014 B.n848 B.n847 51.0063
R2015 B.n847 B.n100 51.0063
R2016 B.n659 B.t6 43.5054
R2017 B.n68 B.t7 43.5054
R2018 B.t5 B.n302 42.0053
R2019 B.n944 B.t1 42.0053
R2020 B.n629 B.t13 40.5051
R2021 B.n863 B.t9 40.5051
R2022 B.n720 B.t0 37.5048
R2023 B.n921 B.t4 37.5048
R2024 B.n696 B.t3 36.0046
R2025 B.n905 B.t2 36.0046
R2026 B.n601 B.n600 32.9371
R2027 B.n448 B.n398 32.9371
R2028 B.n838 B.n837 32.9371
R2029 B.n844 B.n843 32.9371
R2030 B B.n957 18.0485
R2031 B.n346 B.t3 15.0022
R2032 B.t2 B.n904 15.0022
R2033 B.t0 B.n322 13.502
R2034 B.t4 B.n30 13.502
R2035 B.n602 B.n601 10.6151
R2036 B.n602 B.n394 10.6151
R2037 B.n612 B.n394 10.6151
R2038 B.n613 B.n612 10.6151
R2039 B.n614 B.n613 10.6151
R2040 B.n614 B.n386 10.6151
R2041 B.n625 B.n386 10.6151
R2042 B.n626 B.n625 10.6151
R2043 B.n627 B.n626 10.6151
R2044 B.n627 B.n379 10.6151
R2045 B.n637 B.n379 10.6151
R2046 B.n638 B.n637 10.6151
R2047 B.n639 B.n638 10.6151
R2048 B.n639 B.n371 10.6151
R2049 B.n649 B.n371 10.6151
R2050 B.n650 B.n649 10.6151
R2051 B.n651 B.n650 10.6151
R2052 B.n651 B.n363 10.6151
R2053 B.n662 B.n363 10.6151
R2054 B.n663 B.n662 10.6151
R2055 B.n664 B.n663 10.6151
R2056 B.n664 B.n356 10.6151
R2057 B.n674 B.n356 10.6151
R2058 B.n675 B.n674 10.6151
R2059 B.n676 B.n675 10.6151
R2060 B.n676 B.n348 10.6151
R2061 B.n686 B.n348 10.6151
R2062 B.n687 B.n686 10.6151
R2063 B.n688 B.n687 10.6151
R2064 B.n688 B.n340 10.6151
R2065 B.n698 B.n340 10.6151
R2066 B.n699 B.n698 10.6151
R2067 B.n700 B.n699 10.6151
R2068 B.n700 B.n332 10.6151
R2069 B.n710 B.n332 10.6151
R2070 B.n711 B.n710 10.6151
R2071 B.n712 B.n711 10.6151
R2072 B.n712 B.n324 10.6151
R2073 B.n722 B.n324 10.6151
R2074 B.n723 B.n722 10.6151
R2075 B.n724 B.n723 10.6151
R2076 B.n724 B.n316 10.6151
R2077 B.n734 B.n316 10.6151
R2078 B.n735 B.n734 10.6151
R2079 B.n736 B.n735 10.6151
R2080 B.n736 B.n308 10.6151
R2081 B.n746 B.n308 10.6151
R2082 B.n747 B.n746 10.6151
R2083 B.n748 B.n747 10.6151
R2084 B.n748 B.n300 10.6151
R2085 B.n759 B.n300 10.6151
R2086 B.n760 B.n759 10.6151
R2087 B.n761 B.n760 10.6151
R2088 B.n761 B.n0 10.6151
R2089 B.n600 B.n402 10.6151
R2090 B.n595 B.n402 10.6151
R2091 B.n595 B.n594 10.6151
R2092 B.n594 B.n593 10.6151
R2093 B.n593 B.n590 10.6151
R2094 B.n590 B.n589 10.6151
R2095 B.n589 B.n586 10.6151
R2096 B.n586 B.n585 10.6151
R2097 B.n585 B.n582 10.6151
R2098 B.n582 B.n581 10.6151
R2099 B.n581 B.n578 10.6151
R2100 B.n578 B.n577 10.6151
R2101 B.n577 B.n574 10.6151
R2102 B.n574 B.n573 10.6151
R2103 B.n573 B.n570 10.6151
R2104 B.n570 B.n569 10.6151
R2105 B.n569 B.n566 10.6151
R2106 B.n566 B.n565 10.6151
R2107 B.n565 B.n562 10.6151
R2108 B.n562 B.n561 10.6151
R2109 B.n561 B.n558 10.6151
R2110 B.n558 B.n557 10.6151
R2111 B.n557 B.n554 10.6151
R2112 B.n554 B.n553 10.6151
R2113 B.n553 B.n550 10.6151
R2114 B.n550 B.n549 10.6151
R2115 B.n549 B.n546 10.6151
R2116 B.n546 B.n545 10.6151
R2117 B.n545 B.n542 10.6151
R2118 B.n542 B.n541 10.6151
R2119 B.n541 B.n538 10.6151
R2120 B.n538 B.n537 10.6151
R2121 B.n537 B.n534 10.6151
R2122 B.n532 B.n529 10.6151
R2123 B.n529 B.n528 10.6151
R2124 B.n528 B.n525 10.6151
R2125 B.n525 B.n524 10.6151
R2126 B.n524 B.n521 10.6151
R2127 B.n521 B.n520 10.6151
R2128 B.n520 B.n517 10.6151
R2129 B.n517 B.n516 10.6151
R2130 B.n513 B.n512 10.6151
R2131 B.n512 B.n509 10.6151
R2132 B.n509 B.n508 10.6151
R2133 B.n508 B.n505 10.6151
R2134 B.n505 B.n504 10.6151
R2135 B.n504 B.n501 10.6151
R2136 B.n501 B.n500 10.6151
R2137 B.n500 B.n497 10.6151
R2138 B.n497 B.n496 10.6151
R2139 B.n496 B.n493 10.6151
R2140 B.n493 B.n492 10.6151
R2141 B.n492 B.n489 10.6151
R2142 B.n489 B.n488 10.6151
R2143 B.n488 B.n485 10.6151
R2144 B.n485 B.n484 10.6151
R2145 B.n484 B.n481 10.6151
R2146 B.n481 B.n480 10.6151
R2147 B.n480 B.n477 10.6151
R2148 B.n477 B.n476 10.6151
R2149 B.n476 B.n473 10.6151
R2150 B.n473 B.n472 10.6151
R2151 B.n472 B.n469 10.6151
R2152 B.n469 B.n468 10.6151
R2153 B.n468 B.n465 10.6151
R2154 B.n465 B.n464 10.6151
R2155 B.n464 B.n461 10.6151
R2156 B.n461 B.n460 10.6151
R2157 B.n460 B.n457 10.6151
R2158 B.n457 B.n456 10.6151
R2159 B.n456 B.n453 10.6151
R2160 B.n453 B.n452 10.6151
R2161 B.n452 B.n449 10.6151
R2162 B.n449 B.n448 10.6151
R2163 B.n606 B.n398 10.6151
R2164 B.n607 B.n606 10.6151
R2165 B.n608 B.n607 10.6151
R2166 B.n608 B.n390 10.6151
R2167 B.n618 B.n390 10.6151
R2168 B.n619 B.n618 10.6151
R2169 B.n620 B.n619 10.6151
R2170 B.n620 B.n383 10.6151
R2171 B.n631 B.n383 10.6151
R2172 B.n632 B.n631 10.6151
R2173 B.n633 B.n632 10.6151
R2174 B.n633 B.n375 10.6151
R2175 B.n643 B.n375 10.6151
R2176 B.n644 B.n643 10.6151
R2177 B.n645 B.n644 10.6151
R2178 B.n645 B.n367 10.6151
R2179 B.n655 B.n367 10.6151
R2180 B.n656 B.n655 10.6151
R2181 B.n657 B.n656 10.6151
R2182 B.n657 B.n360 10.6151
R2183 B.n668 B.n360 10.6151
R2184 B.n669 B.n668 10.6151
R2185 B.n670 B.n669 10.6151
R2186 B.n670 B.n352 10.6151
R2187 B.n680 B.n352 10.6151
R2188 B.n681 B.n680 10.6151
R2189 B.n682 B.n681 10.6151
R2190 B.n682 B.n343 10.6151
R2191 B.n692 B.n343 10.6151
R2192 B.n693 B.n692 10.6151
R2193 B.n694 B.n693 10.6151
R2194 B.n694 B.n336 10.6151
R2195 B.n704 B.n336 10.6151
R2196 B.n705 B.n704 10.6151
R2197 B.n706 B.n705 10.6151
R2198 B.n706 B.n328 10.6151
R2199 B.n716 B.n328 10.6151
R2200 B.n717 B.n716 10.6151
R2201 B.n718 B.n717 10.6151
R2202 B.n718 B.n320 10.6151
R2203 B.n728 B.n320 10.6151
R2204 B.n729 B.n728 10.6151
R2205 B.n730 B.n729 10.6151
R2206 B.n730 B.n312 10.6151
R2207 B.n740 B.n312 10.6151
R2208 B.n741 B.n740 10.6151
R2209 B.n742 B.n741 10.6151
R2210 B.n742 B.n304 10.6151
R2211 B.n752 B.n304 10.6151
R2212 B.n753 B.n752 10.6151
R2213 B.n755 B.n753 10.6151
R2214 B.n755 B.n754 10.6151
R2215 B.n754 B.n296 10.6151
R2216 B.n766 B.n296 10.6151
R2217 B.n767 B.n766 10.6151
R2218 B.n768 B.n767 10.6151
R2219 B.n769 B.n768 10.6151
R2220 B.n770 B.n769 10.6151
R2221 B.n773 B.n770 10.6151
R2222 B.n774 B.n773 10.6151
R2223 B.n775 B.n774 10.6151
R2224 B.n776 B.n775 10.6151
R2225 B.n778 B.n776 10.6151
R2226 B.n779 B.n778 10.6151
R2227 B.n780 B.n779 10.6151
R2228 B.n781 B.n780 10.6151
R2229 B.n783 B.n781 10.6151
R2230 B.n784 B.n783 10.6151
R2231 B.n785 B.n784 10.6151
R2232 B.n786 B.n785 10.6151
R2233 B.n788 B.n786 10.6151
R2234 B.n789 B.n788 10.6151
R2235 B.n790 B.n789 10.6151
R2236 B.n791 B.n790 10.6151
R2237 B.n793 B.n791 10.6151
R2238 B.n794 B.n793 10.6151
R2239 B.n795 B.n794 10.6151
R2240 B.n796 B.n795 10.6151
R2241 B.n798 B.n796 10.6151
R2242 B.n799 B.n798 10.6151
R2243 B.n800 B.n799 10.6151
R2244 B.n801 B.n800 10.6151
R2245 B.n803 B.n801 10.6151
R2246 B.n804 B.n803 10.6151
R2247 B.n805 B.n804 10.6151
R2248 B.n806 B.n805 10.6151
R2249 B.n808 B.n806 10.6151
R2250 B.n809 B.n808 10.6151
R2251 B.n810 B.n809 10.6151
R2252 B.n811 B.n810 10.6151
R2253 B.n813 B.n811 10.6151
R2254 B.n814 B.n813 10.6151
R2255 B.n815 B.n814 10.6151
R2256 B.n816 B.n815 10.6151
R2257 B.n818 B.n816 10.6151
R2258 B.n819 B.n818 10.6151
R2259 B.n820 B.n819 10.6151
R2260 B.n821 B.n820 10.6151
R2261 B.n823 B.n821 10.6151
R2262 B.n824 B.n823 10.6151
R2263 B.n825 B.n824 10.6151
R2264 B.n826 B.n825 10.6151
R2265 B.n828 B.n826 10.6151
R2266 B.n829 B.n828 10.6151
R2267 B.n830 B.n829 10.6151
R2268 B.n831 B.n830 10.6151
R2269 B.n833 B.n831 10.6151
R2270 B.n834 B.n833 10.6151
R2271 B.n835 B.n834 10.6151
R2272 B.n836 B.n835 10.6151
R2273 B.n837 B.n836 10.6151
R2274 B.n949 B.n1 10.6151
R2275 B.n949 B.n948 10.6151
R2276 B.n948 B.n947 10.6151
R2277 B.n947 B.n10 10.6151
R2278 B.n941 B.n10 10.6151
R2279 B.n941 B.n940 10.6151
R2280 B.n940 B.n939 10.6151
R2281 B.n939 B.n18 10.6151
R2282 B.n933 B.n18 10.6151
R2283 B.n933 B.n932 10.6151
R2284 B.n932 B.n931 10.6151
R2285 B.n931 B.n25 10.6151
R2286 B.n925 B.n25 10.6151
R2287 B.n925 B.n924 10.6151
R2288 B.n924 B.n923 10.6151
R2289 B.n923 B.n32 10.6151
R2290 B.n917 B.n32 10.6151
R2291 B.n917 B.n916 10.6151
R2292 B.n916 B.n915 10.6151
R2293 B.n915 B.n39 10.6151
R2294 B.n909 B.n39 10.6151
R2295 B.n909 B.n908 10.6151
R2296 B.n908 B.n907 10.6151
R2297 B.n907 B.n46 10.6151
R2298 B.n901 B.n46 10.6151
R2299 B.n901 B.n900 10.6151
R2300 B.n900 B.n899 10.6151
R2301 B.n899 B.n53 10.6151
R2302 B.n893 B.n53 10.6151
R2303 B.n893 B.n892 10.6151
R2304 B.n892 B.n891 10.6151
R2305 B.n891 B.n60 10.6151
R2306 B.n885 B.n60 10.6151
R2307 B.n885 B.n884 10.6151
R2308 B.n884 B.n883 10.6151
R2309 B.n883 B.n66 10.6151
R2310 B.n877 B.n66 10.6151
R2311 B.n877 B.n876 10.6151
R2312 B.n876 B.n875 10.6151
R2313 B.n875 B.n74 10.6151
R2314 B.n869 B.n74 10.6151
R2315 B.n869 B.n868 10.6151
R2316 B.n868 B.n867 10.6151
R2317 B.n867 B.n81 10.6151
R2318 B.n861 B.n81 10.6151
R2319 B.n861 B.n860 10.6151
R2320 B.n860 B.n859 10.6151
R2321 B.n859 B.n87 10.6151
R2322 B.n853 B.n87 10.6151
R2323 B.n853 B.n852 10.6151
R2324 B.n852 B.n851 10.6151
R2325 B.n851 B.n95 10.6151
R2326 B.n845 B.n95 10.6151
R2327 B.n845 B.n844 10.6151
R2328 B.n843 B.n102 10.6151
R2329 B.n149 B.n102 10.6151
R2330 B.n150 B.n149 10.6151
R2331 B.n153 B.n150 10.6151
R2332 B.n154 B.n153 10.6151
R2333 B.n157 B.n154 10.6151
R2334 B.n158 B.n157 10.6151
R2335 B.n161 B.n158 10.6151
R2336 B.n162 B.n161 10.6151
R2337 B.n165 B.n162 10.6151
R2338 B.n166 B.n165 10.6151
R2339 B.n169 B.n166 10.6151
R2340 B.n170 B.n169 10.6151
R2341 B.n173 B.n170 10.6151
R2342 B.n174 B.n173 10.6151
R2343 B.n177 B.n174 10.6151
R2344 B.n178 B.n177 10.6151
R2345 B.n181 B.n178 10.6151
R2346 B.n182 B.n181 10.6151
R2347 B.n185 B.n182 10.6151
R2348 B.n186 B.n185 10.6151
R2349 B.n189 B.n186 10.6151
R2350 B.n190 B.n189 10.6151
R2351 B.n193 B.n190 10.6151
R2352 B.n194 B.n193 10.6151
R2353 B.n197 B.n194 10.6151
R2354 B.n198 B.n197 10.6151
R2355 B.n201 B.n198 10.6151
R2356 B.n202 B.n201 10.6151
R2357 B.n205 B.n202 10.6151
R2358 B.n206 B.n205 10.6151
R2359 B.n209 B.n206 10.6151
R2360 B.n210 B.n209 10.6151
R2361 B.n214 B.n213 10.6151
R2362 B.n217 B.n214 10.6151
R2363 B.n218 B.n217 10.6151
R2364 B.n221 B.n218 10.6151
R2365 B.n222 B.n221 10.6151
R2366 B.n225 B.n222 10.6151
R2367 B.n226 B.n225 10.6151
R2368 B.n229 B.n226 10.6151
R2369 B.n234 B.n231 10.6151
R2370 B.n235 B.n234 10.6151
R2371 B.n238 B.n235 10.6151
R2372 B.n239 B.n238 10.6151
R2373 B.n242 B.n239 10.6151
R2374 B.n243 B.n242 10.6151
R2375 B.n246 B.n243 10.6151
R2376 B.n247 B.n246 10.6151
R2377 B.n250 B.n247 10.6151
R2378 B.n251 B.n250 10.6151
R2379 B.n254 B.n251 10.6151
R2380 B.n255 B.n254 10.6151
R2381 B.n258 B.n255 10.6151
R2382 B.n259 B.n258 10.6151
R2383 B.n262 B.n259 10.6151
R2384 B.n263 B.n262 10.6151
R2385 B.n266 B.n263 10.6151
R2386 B.n267 B.n266 10.6151
R2387 B.n270 B.n267 10.6151
R2388 B.n271 B.n270 10.6151
R2389 B.n274 B.n271 10.6151
R2390 B.n275 B.n274 10.6151
R2391 B.n278 B.n275 10.6151
R2392 B.n279 B.n278 10.6151
R2393 B.n282 B.n279 10.6151
R2394 B.n283 B.n282 10.6151
R2395 B.n286 B.n283 10.6151
R2396 B.n287 B.n286 10.6151
R2397 B.n290 B.n287 10.6151
R2398 B.n291 B.n290 10.6151
R2399 B.n294 B.n291 10.6151
R2400 B.n295 B.n294 10.6151
R2401 B.n838 B.n295 10.6151
R2402 B.n622 B.t13 10.5017
R2403 B.n89 B.t9 10.5017
R2404 B.n750 B.t5 9.00152
R2405 B.t1 B.n943 9.00152
R2406 B.n957 B.n0 8.11757
R2407 B.n957 B.n1 8.11757
R2408 B.n666 B.t6 7.50135
R2409 B.n887 B.t7 7.50135
R2410 B.n533 B.n532 6.5566
R2411 B.n516 B.n446 6.5566
R2412 B.n213 B.n147 6.5566
R2413 B.n230 B.n229 6.5566
R2414 B.n534 B.n533 4.05904
R2415 B.n513 B.n446 4.05904
R2416 B.n210 B.n147 4.05904
R2417 B.n231 B.n230 4.05904
R2418 VN.n59 VN.n31 161.3
R2419 VN.n58 VN.n57 161.3
R2420 VN.n56 VN.n32 161.3
R2421 VN.n55 VN.n54 161.3
R2422 VN.n53 VN.n33 161.3
R2423 VN.n52 VN.n51 161.3
R2424 VN.n50 VN.n34 161.3
R2425 VN.n49 VN.n48 161.3
R2426 VN.n47 VN.n35 161.3
R2427 VN.n46 VN.n45 161.3
R2428 VN.n44 VN.n37 161.3
R2429 VN.n43 VN.n42 161.3
R2430 VN.n41 VN.n38 161.3
R2431 VN.n28 VN.n0 161.3
R2432 VN.n27 VN.n26 161.3
R2433 VN.n25 VN.n1 161.3
R2434 VN.n24 VN.n23 161.3
R2435 VN.n22 VN.n2 161.3
R2436 VN.n21 VN.n20 161.3
R2437 VN.n19 VN.n3 161.3
R2438 VN.n18 VN.n17 161.3
R2439 VN.n15 VN.n4 161.3
R2440 VN.n14 VN.n13 161.3
R2441 VN.n12 VN.n5 161.3
R2442 VN.n11 VN.n10 161.3
R2443 VN.n9 VN.n6 161.3
R2444 VN.n7 VN.t0 111.825
R2445 VN.n39 VN.t4 111.825
R2446 VN.n30 VN.n29 107.576
R2447 VN.n61 VN.n60 107.576
R2448 VN.n8 VN.t7 78.5765
R2449 VN.n16 VN.t6 78.5765
R2450 VN.n29 VN.t5 78.5765
R2451 VN.n40 VN.t2 78.5765
R2452 VN.n36 VN.t1 78.5765
R2453 VN.n60 VN.t3 78.5765
R2454 VN.n14 VN.n5 56.5193
R2455 VN.n46 VN.n37 56.5193
R2456 VN.n8 VN.n7 56.3164
R2457 VN.n40 VN.n39 56.3164
R2458 VN VN.n61 50.4906
R2459 VN.n23 VN.n22 44.3785
R2460 VN.n54 VN.n53 44.3785
R2461 VN.n23 VN.n1 36.6083
R2462 VN.n54 VN.n32 36.6083
R2463 VN.n10 VN.n9 24.4675
R2464 VN.n10 VN.n5 24.4675
R2465 VN.n15 VN.n14 24.4675
R2466 VN.n17 VN.n15 24.4675
R2467 VN.n21 VN.n3 24.4675
R2468 VN.n22 VN.n21 24.4675
R2469 VN.n27 VN.n1 24.4675
R2470 VN.n28 VN.n27 24.4675
R2471 VN.n42 VN.n37 24.4675
R2472 VN.n42 VN.n41 24.4675
R2473 VN.n53 VN.n52 24.4675
R2474 VN.n52 VN.n34 24.4675
R2475 VN.n48 VN.n47 24.4675
R2476 VN.n47 VN.n46 24.4675
R2477 VN.n59 VN.n58 24.4675
R2478 VN.n58 VN.n32 24.4675
R2479 VN.n9 VN.n8 17.3721
R2480 VN.n17 VN.n16 17.3721
R2481 VN.n41 VN.n40 17.3721
R2482 VN.n48 VN.n36 17.3721
R2483 VN.n16 VN.n3 7.09593
R2484 VN.n36 VN.n34 7.09593
R2485 VN.n39 VN.n38 5.06027
R2486 VN.n7 VN.n6 5.06027
R2487 VN.n29 VN.n28 3.18121
R2488 VN.n60 VN.n59 3.18121
R2489 VN.n61 VN.n31 0.278367
R2490 VN.n30 VN.n0 0.278367
R2491 VN.n57 VN.n31 0.189894
R2492 VN.n57 VN.n56 0.189894
R2493 VN.n56 VN.n55 0.189894
R2494 VN.n55 VN.n33 0.189894
R2495 VN.n51 VN.n33 0.189894
R2496 VN.n51 VN.n50 0.189894
R2497 VN.n50 VN.n49 0.189894
R2498 VN.n49 VN.n35 0.189894
R2499 VN.n45 VN.n35 0.189894
R2500 VN.n45 VN.n44 0.189894
R2501 VN.n44 VN.n43 0.189894
R2502 VN.n43 VN.n38 0.189894
R2503 VN.n11 VN.n6 0.189894
R2504 VN.n12 VN.n11 0.189894
R2505 VN.n13 VN.n12 0.189894
R2506 VN.n13 VN.n4 0.189894
R2507 VN.n18 VN.n4 0.189894
R2508 VN.n19 VN.n18 0.189894
R2509 VN.n20 VN.n19 0.189894
R2510 VN.n20 VN.n2 0.189894
R2511 VN.n24 VN.n2 0.189894
R2512 VN.n25 VN.n24 0.189894
R2513 VN.n26 VN.n25 0.189894
R2514 VN.n26 VN.n0 0.189894
R2515 VN VN.n30 0.153454
R2516 VDD2.n2 VDD2.n1 67.2392
R2517 VDD2.n2 VDD2.n0 67.2392
R2518 VDD2 VDD2.n5 67.2364
R2519 VDD2.n4 VDD2.n3 65.9111
R2520 VDD2.n4 VDD2.n2 44.2627
R2521 VDD2.n5 VDD2.t5 2.10913
R2522 VDD2.n5 VDD2.t3 2.10913
R2523 VDD2.n3 VDD2.t4 2.10913
R2524 VDD2.n3 VDD2.t6 2.10913
R2525 VDD2.n1 VDD2.t1 2.10913
R2526 VDD2.n1 VDD2.t2 2.10913
R2527 VDD2.n0 VDD2.t7 2.10913
R2528 VDD2.n0 VDD2.t0 2.10913
R2529 VDD2 VDD2.n4 1.44231
C0 VDD2 VP 0.549121f
C1 VN VP 7.52067f
C2 VDD1 VP 7.43471f
C3 VTAIL VP 7.6528f
C4 VN VDD2 7.03901f
C5 VDD1 VDD2 1.92081f
C6 VTAIL VDD2 7.37552f
C7 VN VDD1 0.15189f
C8 VN VTAIL 7.6387f
C9 VTAIL VDD1 7.319231f
C10 VDD2 B 5.399974f
C11 VDD1 B 5.867634f
C12 VTAIL B 9.118374f
C13 VN B 16.362131f
C14 VP B 15.007509f
C15 VDD2.t7 B 0.17938f
C16 VDD2.t0 B 0.17938f
C17 VDD2.n0 B 1.58474f
C18 VDD2.t1 B 0.17938f
C19 VDD2.t2 B 0.17938f
C20 VDD2.n1 B 1.58474f
C21 VDD2.n2 B 3.16027f
C22 VDD2.t4 B 0.17938f
C23 VDD2.t6 B 0.17938f
C24 VDD2.n3 B 1.57441f
C25 VDD2.n4 B 2.74836f
C26 VDD2.t5 B 0.17938f
C27 VDD2.t3 B 0.17938f
C28 VDD2.n5 B 1.58471f
C29 VN.n0 B 0.028213f
C30 VN.t5 B 1.56421f
C31 VN.n1 B 0.043146f
C32 VN.n2 B 0.021399f
C33 VN.n3 B 0.025901f
C34 VN.n4 B 0.021399f
C35 VN.n5 B 0.031239f
C36 VN.n6 B 0.22652f
C37 VN.t7 B 1.56421f
C38 VN.t0 B 1.77401f
C39 VN.n7 B 0.601973f
C40 VN.n8 B 0.63105f
C41 VN.n9 B 0.034171f
C42 VN.n10 B 0.039882f
C43 VN.n11 B 0.021399f
C44 VN.n12 B 0.021399f
C45 VN.n13 B 0.021399f
C46 VN.n14 B 0.031239f
C47 VN.n15 B 0.039882f
C48 VN.t6 B 1.56421f
C49 VN.n16 B 0.560282f
C50 VN.n17 B 0.034171f
C51 VN.n18 B 0.021399f
C52 VN.n19 B 0.021399f
C53 VN.n20 B 0.021399f
C54 VN.n21 B 0.039882f
C55 VN.n22 B 0.041471f
C56 VN.n23 B 0.017743f
C57 VN.n24 B 0.021399f
C58 VN.n25 B 0.021399f
C59 VN.n26 B 0.021399f
C60 VN.n27 B 0.039882f
C61 VN.n28 B 0.022751f
C62 VN.n29 B 0.631984f
C63 VN.n30 B 0.040458f
C64 VN.n31 B 0.028213f
C65 VN.t3 B 1.56421f
C66 VN.n32 B 0.043146f
C67 VN.n33 B 0.021399f
C68 VN.n34 B 0.025901f
C69 VN.n35 B 0.021399f
C70 VN.t1 B 1.56421f
C71 VN.n36 B 0.560282f
C72 VN.n37 B 0.031239f
C73 VN.n38 B 0.22652f
C74 VN.t2 B 1.56421f
C75 VN.t4 B 1.77401f
C76 VN.n39 B 0.601973f
C77 VN.n40 B 0.63105f
C78 VN.n41 B 0.034171f
C79 VN.n42 B 0.039882f
C80 VN.n43 B 0.021399f
C81 VN.n44 B 0.021399f
C82 VN.n45 B 0.021399f
C83 VN.n46 B 0.031239f
C84 VN.n47 B 0.039882f
C85 VN.n48 B 0.034171f
C86 VN.n49 B 0.021399f
C87 VN.n50 B 0.021399f
C88 VN.n51 B 0.021399f
C89 VN.n52 B 0.039882f
C90 VN.n53 B 0.041471f
C91 VN.n54 B 0.017743f
C92 VN.n55 B 0.021399f
C93 VN.n56 B 0.021399f
C94 VN.n57 B 0.021399f
C95 VN.n58 B 0.039882f
C96 VN.n59 B 0.022751f
C97 VN.n60 B 0.631984f
C98 VN.n61 B 1.21537f
C99 VDD1.t0 B 0.181989f
C100 VDD1.t7 B 0.181989f
C101 VDD1.n0 B 1.60885f
C102 VDD1.t6 B 0.181989f
C103 VDD1.t3 B 0.181989f
C104 VDD1.n1 B 1.60779f
C105 VDD1.t4 B 0.181989f
C106 VDD1.t2 B 0.181989f
C107 VDD1.n2 B 1.60779f
C108 VDD1.n3 B 3.25725f
C109 VDD1.t1 B 0.181989f
C110 VDD1.t5 B 0.181989f
C111 VDD1.n4 B 1.5973f
C112 VDD1.n5 B 2.8187f
C113 VTAIL.t4 B 0.156128f
C114 VTAIL.t2 B 0.156128f
C115 VTAIL.n0 B 1.3145f
C116 VTAIL.n1 B 0.387583f
C117 VTAIL.n2 B 0.029433f
C118 VTAIL.n3 B 0.021041f
C119 VTAIL.n4 B 0.011306f
C120 VTAIL.n5 B 0.026724f
C121 VTAIL.n6 B 0.011639f
C122 VTAIL.n7 B 0.021041f
C123 VTAIL.n8 B 0.011972f
C124 VTAIL.n9 B 0.026724f
C125 VTAIL.n10 B 0.011972f
C126 VTAIL.n11 B 0.021041f
C127 VTAIL.n12 B 0.011306f
C128 VTAIL.n13 B 0.026724f
C129 VTAIL.n14 B 0.011972f
C130 VTAIL.n15 B 0.817201f
C131 VTAIL.n16 B 0.011306f
C132 VTAIL.t1 B 0.044844f
C133 VTAIL.n17 B 0.130626f
C134 VTAIL.n18 B 0.018892f
C135 VTAIL.n19 B 0.020043f
C136 VTAIL.n20 B 0.026724f
C137 VTAIL.n21 B 0.011972f
C138 VTAIL.n22 B 0.011306f
C139 VTAIL.n23 B 0.021041f
C140 VTAIL.n24 B 0.021041f
C141 VTAIL.n25 B 0.011306f
C142 VTAIL.n26 B 0.011972f
C143 VTAIL.n27 B 0.026724f
C144 VTAIL.n28 B 0.026724f
C145 VTAIL.n29 B 0.011972f
C146 VTAIL.n30 B 0.011306f
C147 VTAIL.n31 B 0.021041f
C148 VTAIL.n32 B 0.021041f
C149 VTAIL.n33 B 0.011306f
C150 VTAIL.n34 B 0.011306f
C151 VTAIL.n35 B 0.011972f
C152 VTAIL.n36 B 0.026724f
C153 VTAIL.n37 B 0.026724f
C154 VTAIL.n38 B 0.026724f
C155 VTAIL.n39 B 0.011639f
C156 VTAIL.n40 B 0.011306f
C157 VTAIL.n41 B 0.021041f
C158 VTAIL.n42 B 0.021041f
C159 VTAIL.n43 B 0.011306f
C160 VTAIL.n44 B 0.011972f
C161 VTAIL.n45 B 0.026724f
C162 VTAIL.n46 B 0.057603f
C163 VTAIL.n47 B 0.011972f
C164 VTAIL.n48 B 0.011306f
C165 VTAIL.n49 B 0.052946f
C166 VTAIL.n50 B 0.032333f
C167 VTAIL.n51 B 0.239876f
C168 VTAIL.n52 B 0.029433f
C169 VTAIL.n53 B 0.021041f
C170 VTAIL.n54 B 0.011306f
C171 VTAIL.n55 B 0.026724f
C172 VTAIL.n56 B 0.011639f
C173 VTAIL.n57 B 0.021041f
C174 VTAIL.n58 B 0.011972f
C175 VTAIL.n59 B 0.026724f
C176 VTAIL.n60 B 0.011972f
C177 VTAIL.n61 B 0.021041f
C178 VTAIL.n62 B 0.011306f
C179 VTAIL.n63 B 0.026724f
C180 VTAIL.n64 B 0.011972f
C181 VTAIL.n65 B 0.817201f
C182 VTAIL.n66 B 0.011306f
C183 VTAIL.t12 B 0.044844f
C184 VTAIL.n67 B 0.130626f
C185 VTAIL.n68 B 0.018892f
C186 VTAIL.n69 B 0.020043f
C187 VTAIL.n70 B 0.026724f
C188 VTAIL.n71 B 0.011972f
C189 VTAIL.n72 B 0.011306f
C190 VTAIL.n73 B 0.021041f
C191 VTAIL.n74 B 0.021041f
C192 VTAIL.n75 B 0.011306f
C193 VTAIL.n76 B 0.011972f
C194 VTAIL.n77 B 0.026724f
C195 VTAIL.n78 B 0.026724f
C196 VTAIL.n79 B 0.011972f
C197 VTAIL.n80 B 0.011306f
C198 VTAIL.n81 B 0.021041f
C199 VTAIL.n82 B 0.021041f
C200 VTAIL.n83 B 0.011306f
C201 VTAIL.n84 B 0.011306f
C202 VTAIL.n85 B 0.011972f
C203 VTAIL.n86 B 0.026724f
C204 VTAIL.n87 B 0.026724f
C205 VTAIL.n88 B 0.026724f
C206 VTAIL.n89 B 0.011639f
C207 VTAIL.n90 B 0.011306f
C208 VTAIL.n91 B 0.021041f
C209 VTAIL.n92 B 0.021041f
C210 VTAIL.n93 B 0.011306f
C211 VTAIL.n94 B 0.011972f
C212 VTAIL.n95 B 0.026724f
C213 VTAIL.n96 B 0.057603f
C214 VTAIL.n97 B 0.011972f
C215 VTAIL.n98 B 0.011306f
C216 VTAIL.n99 B 0.052946f
C217 VTAIL.n100 B 0.032333f
C218 VTAIL.n101 B 0.239876f
C219 VTAIL.t14 B 0.156128f
C220 VTAIL.t10 B 0.156128f
C221 VTAIL.n102 B 1.3145f
C222 VTAIL.n103 B 0.571252f
C223 VTAIL.n104 B 0.029433f
C224 VTAIL.n105 B 0.021041f
C225 VTAIL.n106 B 0.011306f
C226 VTAIL.n107 B 0.026724f
C227 VTAIL.n108 B 0.011639f
C228 VTAIL.n109 B 0.021041f
C229 VTAIL.n110 B 0.011972f
C230 VTAIL.n111 B 0.026724f
C231 VTAIL.n112 B 0.011972f
C232 VTAIL.n113 B 0.021041f
C233 VTAIL.n114 B 0.011306f
C234 VTAIL.n115 B 0.026724f
C235 VTAIL.n116 B 0.011972f
C236 VTAIL.n117 B 0.817201f
C237 VTAIL.n118 B 0.011306f
C238 VTAIL.t8 B 0.044844f
C239 VTAIL.n119 B 0.130626f
C240 VTAIL.n120 B 0.018892f
C241 VTAIL.n121 B 0.020043f
C242 VTAIL.n122 B 0.026724f
C243 VTAIL.n123 B 0.011972f
C244 VTAIL.n124 B 0.011306f
C245 VTAIL.n125 B 0.021041f
C246 VTAIL.n126 B 0.021041f
C247 VTAIL.n127 B 0.011306f
C248 VTAIL.n128 B 0.011972f
C249 VTAIL.n129 B 0.026724f
C250 VTAIL.n130 B 0.026724f
C251 VTAIL.n131 B 0.011972f
C252 VTAIL.n132 B 0.011306f
C253 VTAIL.n133 B 0.021041f
C254 VTAIL.n134 B 0.021041f
C255 VTAIL.n135 B 0.011306f
C256 VTAIL.n136 B 0.011306f
C257 VTAIL.n137 B 0.011972f
C258 VTAIL.n138 B 0.026724f
C259 VTAIL.n139 B 0.026724f
C260 VTAIL.n140 B 0.026724f
C261 VTAIL.n141 B 0.011639f
C262 VTAIL.n142 B 0.011306f
C263 VTAIL.n143 B 0.021041f
C264 VTAIL.n144 B 0.021041f
C265 VTAIL.n145 B 0.011306f
C266 VTAIL.n146 B 0.011972f
C267 VTAIL.n147 B 0.026724f
C268 VTAIL.n148 B 0.057603f
C269 VTAIL.n149 B 0.011972f
C270 VTAIL.n150 B 0.011306f
C271 VTAIL.n151 B 0.052946f
C272 VTAIL.n152 B 0.032333f
C273 VTAIL.n153 B 1.23027f
C274 VTAIL.n154 B 0.029433f
C275 VTAIL.n155 B 0.021041f
C276 VTAIL.n156 B 0.011306f
C277 VTAIL.n157 B 0.026724f
C278 VTAIL.n158 B 0.011639f
C279 VTAIL.n159 B 0.021041f
C280 VTAIL.n160 B 0.011639f
C281 VTAIL.n161 B 0.011306f
C282 VTAIL.n162 B 0.026724f
C283 VTAIL.n163 B 0.026724f
C284 VTAIL.n164 B 0.011972f
C285 VTAIL.n165 B 0.021041f
C286 VTAIL.n166 B 0.011306f
C287 VTAIL.n167 B 0.026724f
C288 VTAIL.n168 B 0.011972f
C289 VTAIL.n169 B 0.817201f
C290 VTAIL.n170 B 0.011306f
C291 VTAIL.t6 B 0.044844f
C292 VTAIL.n171 B 0.130626f
C293 VTAIL.n172 B 0.018892f
C294 VTAIL.n173 B 0.020043f
C295 VTAIL.n174 B 0.026724f
C296 VTAIL.n175 B 0.011972f
C297 VTAIL.n176 B 0.011306f
C298 VTAIL.n177 B 0.021041f
C299 VTAIL.n178 B 0.021041f
C300 VTAIL.n179 B 0.011306f
C301 VTAIL.n180 B 0.011972f
C302 VTAIL.n181 B 0.026724f
C303 VTAIL.n182 B 0.026724f
C304 VTAIL.n183 B 0.011972f
C305 VTAIL.n184 B 0.011306f
C306 VTAIL.n185 B 0.021041f
C307 VTAIL.n186 B 0.021041f
C308 VTAIL.n187 B 0.011306f
C309 VTAIL.n188 B 0.011972f
C310 VTAIL.n189 B 0.026724f
C311 VTAIL.n190 B 0.026724f
C312 VTAIL.n191 B 0.011972f
C313 VTAIL.n192 B 0.011306f
C314 VTAIL.n193 B 0.021041f
C315 VTAIL.n194 B 0.021041f
C316 VTAIL.n195 B 0.011306f
C317 VTAIL.n196 B 0.011972f
C318 VTAIL.n197 B 0.026724f
C319 VTAIL.n198 B 0.057603f
C320 VTAIL.n199 B 0.011972f
C321 VTAIL.n200 B 0.011306f
C322 VTAIL.n201 B 0.052946f
C323 VTAIL.n202 B 0.032333f
C324 VTAIL.n203 B 1.23027f
C325 VTAIL.t3 B 0.156128f
C326 VTAIL.t0 B 0.156128f
C327 VTAIL.n204 B 1.31451f
C328 VTAIL.n205 B 0.571244f
C329 VTAIL.n206 B 0.029433f
C330 VTAIL.n207 B 0.021041f
C331 VTAIL.n208 B 0.011306f
C332 VTAIL.n209 B 0.026724f
C333 VTAIL.n210 B 0.011639f
C334 VTAIL.n211 B 0.021041f
C335 VTAIL.n212 B 0.011639f
C336 VTAIL.n213 B 0.011306f
C337 VTAIL.n214 B 0.026724f
C338 VTAIL.n215 B 0.026724f
C339 VTAIL.n216 B 0.011972f
C340 VTAIL.n217 B 0.021041f
C341 VTAIL.n218 B 0.011306f
C342 VTAIL.n219 B 0.026724f
C343 VTAIL.n220 B 0.011972f
C344 VTAIL.n221 B 0.817201f
C345 VTAIL.n222 B 0.011306f
C346 VTAIL.t5 B 0.044844f
C347 VTAIL.n223 B 0.130626f
C348 VTAIL.n224 B 0.018892f
C349 VTAIL.n225 B 0.020043f
C350 VTAIL.n226 B 0.026724f
C351 VTAIL.n227 B 0.011972f
C352 VTAIL.n228 B 0.011306f
C353 VTAIL.n229 B 0.021041f
C354 VTAIL.n230 B 0.021041f
C355 VTAIL.n231 B 0.011306f
C356 VTAIL.n232 B 0.011972f
C357 VTAIL.n233 B 0.026724f
C358 VTAIL.n234 B 0.026724f
C359 VTAIL.n235 B 0.011972f
C360 VTAIL.n236 B 0.011306f
C361 VTAIL.n237 B 0.021041f
C362 VTAIL.n238 B 0.021041f
C363 VTAIL.n239 B 0.011306f
C364 VTAIL.n240 B 0.011972f
C365 VTAIL.n241 B 0.026724f
C366 VTAIL.n242 B 0.026724f
C367 VTAIL.n243 B 0.011972f
C368 VTAIL.n244 B 0.011306f
C369 VTAIL.n245 B 0.021041f
C370 VTAIL.n246 B 0.021041f
C371 VTAIL.n247 B 0.011306f
C372 VTAIL.n248 B 0.011972f
C373 VTAIL.n249 B 0.026724f
C374 VTAIL.n250 B 0.057603f
C375 VTAIL.n251 B 0.011972f
C376 VTAIL.n252 B 0.011306f
C377 VTAIL.n253 B 0.052946f
C378 VTAIL.n254 B 0.032333f
C379 VTAIL.n255 B 0.239876f
C380 VTAIL.n256 B 0.029433f
C381 VTAIL.n257 B 0.021041f
C382 VTAIL.n258 B 0.011306f
C383 VTAIL.n259 B 0.026724f
C384 VTAIL.n260 B 0.011639f
C385 VTAIL.n261 B 0.021041f
C386 VTAIL.n262 B 0.011639f
C387 VTAIL.n263 B 0.011306f
C388 VTAIL.n264 B 0.026724f
C389 VTAIL.n265 B 0.026724f
C390 VTAIL.n266 B 0.011972f
C391 VTAIL.n267 B 0.021041f
C392 VTAIL.n268 B 0.011306f
C393 VTAIL.n269 B 0.026724f
C394 VTAIL.n270 B 0.011972f
C395 VTAIL.n271 B 0.817201f
C396 VTAIL.n272 B 0.011306f
C397 VTAIL.t7 B 0.044844f
C398 VTAIL.n273 B 0.130626f
C399 VTAIL.n274 B 0.018892f
C400 VTAIL.n275 B 0.020043f
C401 VTAIL.n276 B 0.026724f
C402 VTAIL.n277 B 0.011972f
C403 VTAIL.n278 B 0.011306f
C404 VTAIL.n279 B 0.021041f
C405 VTAIL.n280 B 0.021041f
C406 VTAIL.n281 B 0.011306f
C407 VTAIL.n282 B 0.011972f
C408 VTAIL.n283 B 0.026724f
C409 VTAIL.n284 B 0.026724f
C410 VTAIL.n285 B 0.011972f
C411 VTAIL.n286 B 0.011306f
C412 VTAIL.n287 B 0.021041f
C413 VTAIL.n288 B 0.021041f
C414 VTAIL.n289 B 0.011306f
C415 VTAIL.n290 B 0.011972f
C416 VTAIL.n291 B 0.026724f
C417 VTAIL.n292 B 0.026724f
C418 VTAIL.n293 B 0.011972f
C419 VTAIL.n294 B 0.011306f
C420 VTAIL.n295 B 0.021041f
C421 VTAIL.n296 B 0.021041f
C422 VTAIL.n297 B 0.011306f
C423 VTAIL.n298 B 0.011972f
C424 VTAIL.n299 B 0.026724f
C425 VTAIL.n300 B 0.057603f
C426 VTAIL.n301 B 0.011972f
C427 VTAIL.n302 B 0.011306f
C428 VTAIL.n303 B 0.052946f
C429 VTAIL.n304 B 0.032333f
C430 VTAIL.n305 B 0.239876f
C431 VTAIL.t11 B 0.156128f
C432 VTAIL.t13 B 0.156128f
C433 VTAIL.n306 B 1.31451f
C434 VTAIL.n307 B 0.571244f
C435 VTAIL.n308 B 0.029433f
C436 VTAIL.n309 B 0.021041f
C437 VTAIL.n310 B 0.011306f
C438 VTAIL.n311 B 0.026724f
C439 VTAIL.n312 B 0.011639f
C440 VTAIL.n313 B 0.021041f
C441 VTAIL.n314 B 0.011639f
C442 VTAIL.n315 B 0.011306f
C443 VTAIL.n316 B 0.026724f
C444 VTAIL.n317 B 0.026724f
C445 VTAIL.n318 B 0.011972f
C446 VTAIL.n319 B 0.021041f
C447 VTAIL.n320 B 0.011306f
C448 VTAIL.n321 B 0.026724f
C449 VTAIL.n322 B 0.011972f
C450 VTAIL.n323 B 0.817201f
C451 VTAIL.n324 B 0.011306f
C452 VTAIL.t9 B 0.044844f
C453 VTAIL.n325 B 0.130626f
C454 VTAIL.n326 B 0.018892f
C455 VTAIL.n327 B 0.020043f
C456 VTAIL.n328 B 0.026724f
C457 VTAIL.n329 B 0.011972f
C458 VTAIL.n330 B 0.011306f
C459 VTAIL.n331 B 0.021041f
C460 VTAIL.n332 B 0.021041f
C461 VTAIL.n333 B 0.011306f
C462 VTAIL.n334 B 0.011972f
C463 VTAIL.n335 B 0.026724f
C464 VTAIL.n336 B 0.026724f
C465 VTAIL.n337 B 0.011972f
C466 VTAIL.n338 B 0.011306f
C467 VTAIL.n339 B 0.021041f
C468 VTAIL.n340 B 0.021041f
C469 VTAIL.n341 B 0.011306f
C470 VTAIL.n342 B 0.011972f
C471 VTAIL.n343 B 0.026724f
C472 VTAIL.n344 B 0.026724f
C473 VTAIL.n345 B 0.011972f
C474 VTAIL.n346 B 0.011306f
C475 VTAIL.n347 B 0.021041f
C476 VTAIL.n348 B 0.021041f
C477 VTAIL.n349 B 0.011306f
C478 VTAIL.n350 B 0.011972f
C479 VTAIL.n351 B 0.026724f
C480 VTAIL.n352 B 0.057603f
C481 VTAIL.n353 B 0.011972f
C482 VTAIL.n354 B 0.011306f
C483 VTAIL.n355 B 0.052946f
C484 VTAIL.n356 B 0.032333f
C485 VTAIL.n357 B 1.23027f
C486 VTAIL.n358 B 0.029433f
C487 VTAIL.n359 B 0.021041f
C488 VTAIL.n360 B 0.011306f
C489 VTAIL.n361 B 0.026724f
C490 VTAIL.n362 B 0.011639f
C491 VTAIL.n363 B 0.021041f
C492 VTAIL.n364 B 0.011972f
C493 VTAIL.n365 B 0.026724f
C494 VTAIL.n366 B 0.011972f
C495 VTAIL.n367 B 0.021041f
C496 VTAIL.n368 B 0.011306f
C497 VTAIL.n369 B 0.026724f
C498 VTAIL.n370 B 0.011972f
C499 VTAIL.n371 B 0.817201f
C500 VTAIL.n372 B 0.011306f
C501 VTAIL.t15 B 0.044844f
C502 VTAIL.n373 B 0.130626f
C503 VTAIL.n374 B 0.018892f
C504 VTAIL.n375 B 0.020043f
C505 VTAIL.n376 B 0.026724f
C506 VTAIL.n377 B 0.011972f
C507 VTAIL.n378 B 0.011306f
C508 VTAIL.n379 B 0.021041f
C509 VTAIL.n380 B 0.021041f
C510 VTAIL.n381 B 0.011306f
C511 VTAIL.n382 B 0.011972f
C512 VTAIL.n383 B 0.026724f
C513 VTAIL.n384 B 0.026724f
C514 VTAIL.n385 B 0.011972f
C515 VTAIL.n386 B 0.011306f
C516 VTAIL.n387 B 0.021041f
C517 VTAIL.n388 B 0.021041f
C518 VTAIL.n389 B 0.011306f
C519 VTAIL.n390 B 0.011306f
C520 VTAIL.n391 B 0.011972f
C521 VTAIL.n392 B 0.026724f
C522 VTAIL.n393 B 0.026724f
C523 VTAIL.n394 B 0.026724f
C524 VTAIL.n395 B 0.011639f
C525 VTAIL.n396 B 0.011306f
C526 VTAIL.n397 B 0.021041f
C527 VTAIL.n398 B 0.021041f
C528 VTAIL.n399 B 0.011306f
C529 VTAIL.n400 B 0.011972f
C530 VTAIL.n401 B 0.026724f
C531 VTAIL.n402 B 0.057603f
C532 VTAIL.n403 B 0.011972f
C533 VTAIL.n404 B 0.011306f
C534 VTAIL.n405 B 0.052946f
C535 VTAIL.n406 B 0.032333f
C536 VTAIL.n407 B 1.22632f
C537 VP.n0 B 0.02889f
C538 VP.t5 B 1.60178f
C539 VP.n1 B 0.044182f
C540 VP.n2 B 0.021913f
C541 VP.n3 B 0.026524f
C542 VP.n4 B 0.021913f
C543 VP.n5 B 0.031989f
C544 VP.n6 B 0.021913f
C545 VP.t4 B 1.60178f
C546 VP.n7 B 0.04084f
C547 VP.n8 B 0.021913f
C548 VP.n9 B 0.04084f
C549 VP.n10 B 0.02889f
C550 VP.t2 B 1.60178f
C551 VP.n11 B 0.044182f
C552 VP.n12 B 0.021913f
C553 VP.n13 B 0.026524f
C554 VP.n14 B 0.021913f
C555 VP.n15 B 0.031989f
C556 VP.n16 B 0.231961f
C557 VP.t0 B 1.60178f
C558 VP.t7 B 1.81662f
C559 VP.n17 B 0.616431f
C560 VP.n18 B 0.646207f
C561 VP.n19 B 0.034992f
C562 VP.n20 B 0.04084f
C563 VP.n21 B 0.021913f
C564 VP.n22 B 0.021913f
C565 VP.n23 B 0.021913f
C566 VP.n24 B 0.031989f
C567 VP.n25 B 0.04084f
C568 VP.t6 B 1.60178f
C569 VP.n26 B 0.573739f
C570 VP.n27 B 0.034992f
C571 VP.n28 B 0.021913f
C572 VP.n29 B 0.021913f
C573 VP.n30 B 0.021913f
C574 VP.n31 B 0.04084f
C575 VP.n32 B 0.042467f
C576 VP.n33 B 0.018169f
C577 VP.n34 B 0.021913f
C578 VP.n35 B 0.021913f
C579 VP.n36 B 0.021913f
C580 VP.n37 B 0.04084f
C581 VP.n38 B 0.023297f
C582 VP.n39 B 0.647163f
C583 VP.n40 B 1.2328f
C584 VP.n41 B 1.24848f
C585 VP.t1 B 1.60178f
C586 VP.n42 B 0.647163f
C587 VP.n43 B 0.023297f
C588 VP.n44 B 0.02889f
C589 VP.n45 B 0.021913f
C590 VP.n46 B 0.021913f
C591 VP.n47 B 0.044182f
C592 VP.n48 B 0.018169f
C593 VP.n49 B 0.042467f
C594 VP.n50 B 0.021913f
C595 VP.n51 B 0.021913f
C596 VP.n52 B 0.021913f
C597 VP.n53 B 0.026524f
C598 VP.n54 B 0.573739f
C599 VP.n55 B 0.034992f
C600 VP.n56 B 0.04084f
C601 VP.n57 B 0.021913f
C602 VP.n58 B 0.021913f
C603 VP.n59 B 0.021913f
C604 VP.n60 B 0.031989f
C605 VP.n61 B 0.04084f
C606 VP.t3 B 1.60178f
C607 VP.n62 B 0.573739f
C608 VP.n63 B 0.034992f
C609 VP.n64 B 0.021913f
C610 VP.n65 B 0.021913f
C611 VP.n66 B 0.021913f
C612 VP.n67 B 0.04084f
C613 VP.n68 B 0.042467f
C614 VP.n69 B 0.018169f
C615 VP.n70 B 0.021913f
C616 VP.n71 B 0.021913f
C617 VP.n72 B 0.021913f
C618 VP.n73 B 0.04084f
C619 VP.n74 B 0.023297f
C620 VP.n75 B 0.647163f
C621 VP.n76 B 0.04143f
.ends

