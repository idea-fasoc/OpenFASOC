* NGSPICE file created from diff_pair_sample_0732.ext - technology: sky130A

.subckt diff_pair_sample_0732 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8876 pd=10.46 as=0 ps=0 w=4.84 l=2.29
X1 VDD1.t1 VP.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8876 pd=10.46 as=1.8876 ps=10.46 w=4.84 l=2.29
X2 VDD1.t0 VP.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.8876 pd=10.46 as=1.8876 ps=10.46 w=4.84 l=2.29
X3 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.8876 pd=10.46 as=0 ps=0 w=4.84 l=2.29
X4 VDD2.t1 VN.t0 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8876 pd=10.46 as=1.8876 ps=10.46 w=4.84 l=2.29
X5 VDD2.t0 VN.t1 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.8876 pd=10.46 as=1.8876 ps=10.46 w=4.84 l=2.29
X6 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.8876 pd=10.46 as=0 ps=0 w=4.84 l=2.29
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8876 pd=10.46 as=0 ps=0 w=4.84 l=2.29
R0 B.n453 B.n452 585
R1 B.n454 B.n453 585
R2 B.n174 B.n72 585
R3 B.n173 B.n172 585
R4 B.n171 B.n170 585
R5 B.n169 B.n168 585
R6 B.n167 B.n166 585
R7 B.n165 B.n164 585
R8 B.n163 B.n162 585
R9 B.n161 B.n160 585
R10 B.n159 B.n158 585
R11 B.n157 B.n156 585
R12 B.n155 B.n154 585
R13 B.n153 B.n152 585
R14 B.n151 B.n150 585
R15 B.n149 B.n148 585
R16 B.n147 B.n146 585
R17 B.n145 B.n144 585
R18 B.n143 B.n142 585
R19 B.n141 B.n140 585
R20 B.n139 B.n138 585
R21 B.n137 B.n136 585
R22 B.n135 B.n134 585
R23 B.n133 B.n132 585
R24 B.n131 B.n130 585
R25 B.n129 B.n128 585
R26 B.n127 B.n126 585
R27 B.n125 B.n124 585
R28 B.n123 B.n122 585
R29 B.n121 B.n120 585
R30 B.n119 B.n118 585
R31 B.n116 B.n115 585
R32 B.n114 B.n113 585
R33 B.n112 B.n111 585
R34 B.n110 B.n109 585
R35 B.n108 B.n107 585
R36 B.n106 B.n105 585
R37 B.n104 B.n103 585
R38 B.n102 B.n101 585
R39 B.n100 B.n99 585
R40 B.n98 B.n97 585
R41 B.n96 B.n95 585
R42 B.n94 B.n93 585
R43 B.n92 B.n91 585
R44 B.n90 B.n89 585
R45 B.n88 B.n87 585
R46 B.n86 B.n85 585
R47 B.n84 B.n83 585
R48 B.n82 B.n81 585
R49 B.n80 B.n79 585
R50 B.n47 B.n46 585
R51 B.n457 B.n456 585
R52 B.n451 B.n73 585
R53 B.n73 B.n44 585
R54 B.n450 B.n43 585
R55 B.n461 B.n43 585
R56 B.n449 B.n42 585
R57 B.n462 B.n42 585
R58 B.n448 B.n41 585
R59 B.n463 B.n41 585
R60 B.n447 B.n446 585
R61 B.n446 B.n37 585
R62 B.n445 B.n36 585
R63 B.n469 B.n36 585
R64 B.n444 B.n35 585
R65 B.n470 B.n35 585
R66 B.n443 B.n34 585
R67 B.n471 B.n34 585
R68 B.n442 B.n441 585
R69 B.n441 B.n30 585
R70 B.n440 B.n29 585
R71 B.n477 B.n29 585
R72 B.n439 B.n28 585
R73 B.n478 B.n28 585
R74 B.n438 B.n27 585
R75 B.n479 B.n27 585
R76 B.n437 B.n436 585
R77 B.n436 B.n23 585
R78 B.n435 B.n22 585
R79 B.n485 B.n22 585
R80 B.n434 B.n21 585
R81 B.n486 B.n21 585
R82 B.n433 B.n20 585
R83 B.n487 B.n20 585
R84 B.n432 B.n431 585
R85 B.n431 B.n16 585
R86 B.n430 B.n15 585
R87 B.n493 B.n15 585
R88 B.n429 B.n14 585
R89 B.n494 B.n14 585
R90 B.n428 B.n13 585
R91 B.n495 B.n13 585
R92 B.n427 B.n426 585
R93 B.n426 B.n12 585
R94 B.n425 B.n424 585
R95 B.n425 B.n8 585
R96 B.n423 B.n7 585
R97 B.n502 B.n7 585
R98 B.n422 B.n6 585
R99 B.n503 B.n6 585
R100 B.n421 B.n5 585
R101 B.n504 B.n5 585
R102 B.n420 B.n419 585
R103 B.n419 B.n4 585
R104 B.n418 B.n175 585
R105 B.n418 B.n417 585
R106 B.n408 B.n176 585
R107 B.n177 B.n176 585
R108 B.n410 B.n409 585
R109 B.n411 B.n410 585
R110 B.n407 B.n181 585
R111 B.n185 B.n181 585
R112 B.n406 B.n405 585
R113 B.n405 B.n404 585
R114 B.n183 B.n182 585
R115 B.n184 B.n183 585
R116 B.n397 B.n396 585
R117 B.n398 B.n397 585
R118 B.n395 B.n190 585
R119 B.n190 B.n189 585
R120 B.n394 B.n393 585
R121 B.n393 B.n392 585
R122 B.n192 B.n191 585
R123 B.n193 B.n192 585
R124 B.n385 B.n384 585
R125 B.n386 B.n385 585
R126 B.n383 B.n198 585
R127 B.n198 B.n197 585
R128 B.n382 B.n381 585
R129 B.n381 B.n380 585
R130 B.n200 B.n199 585
R131 B.n201 B.n200 585
R132 B.n373 B.n372 585
R133 B.n374 B.n373 585
R134 B.n371 B.n206 585
R135 B.n206 B.n205 585
R136 B.n370 B.n369 585
R137 B.n369 B.n368 585
R138 B.n208 B.n207 585
R139 B.n209 B.n208 585
R140 B.n361 B.n360 585
R141 B.n362 B.n361 585
R142 B.n359 B.n214 585
R143 B.n214 B.n213 585
R144 B.n358 B.n357 585
R145 B.n357 B.n356 585
R146 B.n216 B.n215 585
R147 B.n217 B.n216 585
R148 B.n352 B.n351 585
R149 B.n220 B.n219 585
R150 B.n348 B.n347 585
R151 B.n349 B.n348 585
R152 B.n346 B.n245 585
R153 B.n345 B.n344 585
R154 B.n343 B.n342 585
R155 B.n341 B.n340 585
R156 B.n339 B.n338 585
R157 B.n337 B.n336 585
R158 B.n335 B.n334 585
R159 B.n333 B.n332 585
R160 B.n331 B.n330 585
R161 B.n329 B.n328 585
R162 B.n327 B.n326 585
R163 B.n325 B.n324 585
R164 B.n323 B.n322 585
R165 B.n321 B.n320 585
R166 B.n319 B.n318 585
R167 B.n317 B.n316 585
R168 B.n315 B.n314 585
R169 B.n313 B.n312 585
R170 B.n311 B.n310 585
R171 B.n309 B.n308 585
R172 B.n307 B.n306 585
R173 B.n305 B.n304 585
R174 B.n303 B.n302 585
R175 B.n301 B.n300 585
R176 B.n299 B.n298 585
R177 B.n297 B.n296 585
R178 B.n295 B.n294 585
R179 B.n292 B.n291 585
R180 B.n290 B.n289 585
R181 B.n288 B.n287 585
R182 B.n286 B.n285 585
R183 B.n284 B.n283 585
R184 B.n282 B.n281 585
R185 B.n280 B.n279 585
R186 B.n278 B.n277 585
R187 B.n276 B.n275 585
R188 B.n274 B.n273 585
R189 B.n272 B.n271 585
R190 B.n270 B.n269 585
R191 B.n268 B.n267 585
R192 B.n266 B.n265 585
R193 B.n264 B.n263 585
R194 B.n262 B.n261 585
R195 B.n260 B.n259 585
R196 B.n258 B.n257 585
R197 B.n256 B.n255 585
R198 B.n254 B.n253 585
R199 B.n252 B.n251 585
R200 B.n353 B.n218 585
R201 B.n218 B.n217 585
R202 B.n355 B.n354 585
R203 B.n356 B.n355 585
R204 B.n212 B.n211 585
R205 B.n213 B.n212 585
R206 B.n364 B.n363 585
R207 B.n363 B.n362 585
R208 B.n365 B.n210 585
R209 B.n210 B.n209 585
R210 B.n367 B.n366 585
R211 B.n368 B.n367 585
R212 B.n204 B.n203 585
R213 B.n205 B.n204 585
R214 B.n376 B.n375 585
R215 B.n375 B.n374 585
R216 B.n377 B.n202 585
R217 B.n202 B.n201 585
R218 B.n379 B.n378 585
R219 B.n380 B.n379 585
R220 B.n196 B.n195 585
R221 B.n197 B.n196 585
R222 B.n388 B.n387 585
R223 B.n387 B.n386 585
R224 B.n389 B.n194 585
R225 B.n194 B.n193 585
R226 B.n391 B.n390 585
R227 B.n392 B.n391 585
R228 B.n188 B.n187 585
R229 B.n189 B.n188 585
R230 B.n400 B.n399 585
R231 B.n399 B.n398 585
R232 B.n401 B.n186 585
R233 B.n186 B.n184 585
R234 B.n403 B.n402 585
R235 B.n404 B.n403 585
R236 B.n180 B.n179 585
R237 B.n185 B.n180 585
R238 B.n413 B.n412 585
R239 B.n412 B.n411 585
R240 B.n414 B.n178 585
R241 B.n178 B.n177 585
R242 B.n416 B.n415 585
R243 B.n417 B.n416 585
R244 B.n3 B.n0 585
R245 B.n4 B.n3 585
R246 B.n501 B.n1 585
R247 B.n502 B.n501 585
R248 B.n500 B.n499 585
R249 B.n500 B.n8 585
R250 B.n498 B.n9 585
R251 B.n12 B.n9 585
R252 B.n497 B.n496 585
R253 B.n496 B.n495 585
R254 B.n11 B.n10 585
R255 B.n494 B.n11 585
R256 B.n492 B.n491 585
R257 B.n493 B.n492 585
R258 B.n490 B.n17 585
R259 B.n17 B.n16 585
R260 B.n489 B.n488 585
R261 B.n488 B.n487 585
R262 B.n19 B.n18 585
R263 B.n486 B.n19 585
R264 B.n484 B.n483 585
R265 B.n485 B.n484 585
R266 B.n482 B.n24 585
R267 B.n24 B.n23 585
R268 B.n481 B.n480 585
R269 B.n480 B.n479 585
R270 B.n26 B.n25 585
R271 B.n478 B.n26 585
R272 B.n476 B.n475 585
R273 B.n477 B.n476 585
R274 B.n474 B.n31 585
R275 B.n31 B.n30 585
R276 B.n473 B.n472 585
R277 B.n472 B.n471 585
R278 B.n33 B.n32 585
R279 B.n470 B.n33 585
R280 B.n468 B.n467 585
R281 B.n469 B.n468 585
R282 B.n466 B.n38 585
R283 B.n38 B.n37 585
R284 B.n465 B.n464 585
R285 B.n464 B.n463 585
R286 B.n40 B.n39 585
R287 B.n462 B.n40 585
R288 B.n460 B.n459 585
R289 B.n461 B.n460 585
R290 B.n458 B.n45 585
R291 B.n45 B.n44 585
R292 B.n505 B.n504 585
R293 B.n503 B.n2 585
R294 B.n456 B.n45 478.086
R295 B.n453 B.n73 478.086
R296 B.n251 B.n216 478.086
R297 B.n351 B.n218 478.086
R298 B.n77 B.t6 258.462
R299 B.n74 B.t10 258.462
R300 B.n249 B.t13 258.462
R301 B.n246 B.t2 258.462
R302 B.n454 B.n71 256.663
R303 B.n454 B.n70 256.663
R304 B.n454 B.n69 256.663
R305 B.n454 B.n68 256.663
R306 B.n454 B.n67 256.663
R307 B.n454 B.n66 256.663
R308 B.n454 B.n65 256.663
R309 B.n454 B.n64 256.663
R310 B.n454 B.n63 256.663
R311 B.n454 B.n62 256.663
R312 B.n454 B.n61 256.663
R313 B.n454 B.n60 256.663
R314 B.n454 B.n59 256.663
R315 B.n454 B.n58 256.663
R316 B.n454 B.n57 256.663
R317 B.n454 B.n56 256.663
R318 B.n454 B.n55 256.663
R319 B.n454 B.n54 256.663
R320 B.n454 B.n53 256.663
R321 B.n454 B.n52 256.663
R322 B.n454 B.n51 256.663
R323 B.n454 B.n50 256.663
R324 B.n454 B.n49 256.663
R325 B.n454 B.n48 256.663
R326 B.n455 B.n454 256.663
R327 B.n350 B.n349 256.663
R328 B.n349 B.n221 256.663
R329 B.n349 B.n222 256.663
R330 B.n349 B.n223 256.663
R331 B.n349 B.n224 256.663
R332 B.n349 B.n225 256.663
R333 B.n349 B.n226 256.663
R334 B.n349 B.n227 256.663
R335 B.n349 B.n228 256.663
R336 B.n349 B.n229 256.663
R337 B.n349 B.n230 256.663
R338 B.n349 B.n231 256.663
R339 B.n349 B.n232 256.663
R340 B.n349 B.n233 256.663
R341 B.n349 B.n234 256.663
R342 B.n349 B.n235 256.663
R343 B.n349 B.n236 256.663
R344 B.n349 B.n237 256.663
R345 B.n349 B.n238 256.663
R346 B.n349 B.n239 256.663
R347 B.n349 B.n240 256.663
R348 B.n349 B.n241 256.663
R349 B.n349 B.n242 256.663
R350 B.n349 B.n243 256.663
R351 B.n349 B.n244 256.663
R352 B.n507 B.n506 256.663
R353 B.n79 B.n47 163.367
R354 B.n83 B.n82 163.367
R355 B.n87 B.n86 163.367
R356 B.n91 B.n90 163.367
R357 B.n95 B.n94 163.367
R358 B.n99 B.n98 163.367
R359 B.n103 B.n102 163.367
R360 B.n107 B.n106 163.367
R361 B.n111 B.n110 163.367
R362 B.n115 B.n114 163.367
R363 B.n120 B.n119 163.367
R364 B.n124 B.n123 163.367
R365 B.n128 B.n127 163.367
R366 B.n132 B.n131 163.367
R367 B.n136 B.n135 163.367
R368 B.n140 B.n139 163.367
R369 B.n144 B.n143 163.367
R370 B.n148 B.n147 163.367
R371 B.n152 B.n151 163.367
R372 B.n156 B.n155 163.367
R373 B.n160 B.n159 163.367
R374 B.n164 B.n163 163.367
R375 B.n168 B.n167 163.367
R376 B.n172 B.n171 163.367
R377 B.n453 B.n72 163.367
R378 B.n357 B.n216 163.367
R379 B.n357 B.n214 163.367
R380 B.n361 B.n214 163.367
R381 B.n361 B.n208 163.367
R382 B.n369 B.n208 163.367
R383 B.n369 B.n206 163.367
R384 B.n373 B.n206 163.367
R385 B.n373 B.n200 163.367
R386 B.n381 B.n200 163.367
R387 B.n381 B.n198 163.367
R388 B.n385 B.n198 163.367
R389 B.n385 B.n192 163.367
R390 B.n393 B.n192 163.367
R391 B.n393 B.n190 163.367
R392 B.n397 B.n190 163.367
R393 B.n397 B.n183 163.367
R394 B.n405 B.n183 163.367
R395 B.n405 B.n181 163.367
R396 B.n410 B.n181 163.367
R397 B.n410 B.n176 163.367
R398 B.n418 B.n176 163.367
R399 B.n419 B.n418 163.367
R400 B.n419 B.n5 163.367
R401 B.n6 B.n5 163.367
R402 B.n7 B.n6 163.367
R403 B.n425 B.n7 163.367
R404 B.n426 B.n425 163.367
R405 B.n426 B.n13 163.367
R406 B.n14 B.n13 163.367
R407 B.n15 B.n14 163.367
R408 B.n431 B.n15 163.367
R409 B.n431 B.n20 163.367
R410 B.n21 B.n20 163.367
R411 B.n22 B.n21 163.367
R412 B.n436 B.n22 163.367
R413 B.n436 B.n27 163.367
R414 B.n28 B.n27 163.367
R415 B.n29 B.n28 163.367
R416 B.n441 B.n29 163.367
R417 B.n441 B.n34 163.367
R418 B.n35 B.n34 163.367
R419 B.n36 B.n35 163.367
R420 B.n446 B.n36 163.367
R421 B.n446 B.n41 163.367
R422 B.n42 B.n41 163.367
R423 B.n43 B.n42 163.367
R424 B.n73 B.n43 163.367
R425 B.n348 B.n220 163.367
R426 B.n348 B.n245 163.367
R427 B.n344 B.n343 163.367
R428 B.n340 B.n339 163.367
R429 B.n336 B.n335 163.367
R430 B.n332 B.n331 163.367
R431 B.n328 B.n327 163.367
R432 B.n324 B.n323 163.367
R433 B.n320 B.n319 163.367
R434 B.n316 B.n315 163.367
R435 B.n312 B.n311 163.367
R436 B.n308 B.n307 163.367
R437 B.n304 B.n303 163.367
R438 B.n300 B.n299 163.367
R439 B.n296 B.n295 163.367
R440 B.n291 B.n290 163.367
R441 B.n287 B.n286 163.367
R442 B.n283 B.n282 163.367
R443 B.n279 B.n278 163.367
R444 B.n275 B.n274 163.367
R445 B.n271 B.n270 163.367
R446 B.n267 B.n266 163.367
R447 B.n263 B.n262 163.367
R448 B.n259 B.n258 163.367
R449 B.n255 B.n254 163.367
R450 B.n355 B.n218 163.367
R451 B.n355 B.n212 163.367
R452 B.n363 B.n212 163.367
R453 B.n363 B.n210 163.367
R454 B.n367 B.n210 163.367
R455 B.n367 B.n204 163.367
R456 B.n375 B.n204 163.367
R457 B.n375 B.n202 163.367
R458 B.n379 B.n202 163.367
R459 B.n379 B.n196 163.367
R460 B.n387 B.n196 163.367
R461 B.n387 B.n194 163.367
R462 B.n391 B.n194 163.367
R463 B.n391 B.n188 163.367
R464 B.n399 B.n188 163.367
R465 B.n399 B.n186 163.367
R466 B.n403 B.n186 163.367
R467 B.n403 B.n180 163.367
R468 B.n412 B.n180 163.367
R469 B.n412 B.n178 163.367
R470 B.n416 B.n178 163.367
R471 B.n416 B.n3 163.367
R472 B.n505 B.n3 163.367
R473 B.n501 B.n2 163.367
R474 B.n501 B.n500 163.367
R475 B.n500 B.n9 163.367
R476 B.n496 B.n9 163.367
R477 B.n496 B.n11 163.367
R478 B.n492 B.n11 163.367
R479 B.n492 B.n17 163.367
R480 B.n488 B.n17 163.367
R481 B.n488 B.n19 163.367
R482 B.n484 B.n19 163.367
R483 B.n484 B.n24 163.367
R484 B.n480 B.n24 163.367
R485 B.n480 B.n26 163.367
R486 B.n476 B.n26 163.367
R487 B.n476 B.n31 163.367
R488 B.n472 B.n31 163.367
R489 B.n472 B.n33 163.367
R490 B.n468 B.n33 163.367
R491 B.n468 B.n38 163.367
R492 B.n464 B.n38 163.367
R493 B.n464 B.n40 163.367
R494 B.n460 B.n40 163.367
R495 B.n460 B.n45 163.367
R496 B.n349 B.n217 135.938
R497 B.n454 B.n44 135.938
R498 B.n74 B.t11 122.683
R499 B.n249 B.t15 122.683
R500 B.n77 B.t8 122.677
R501 B.n246 B.t5 122.677
R502 B.n356 B.n217 73.9501
R503 B.n356 B.n213 73.9501
R504 B.n362 B.n213 73.9501
R505 B.n362 B.n209 73.9501
R506 B.n368 B.n209 73.9501
R507 B.n368 B.n205 73.9501
R508 B.n374 B.n205 73.9501
R509 B.n380 B.n201 73.9501
R510 B.n380 B.n197 73.9501
R511 B.n386 B.n197 73.9501
R512 B.n386 B.n193 73.9501
R513 B.n392 B.n193 73.9501
R514 B.n392 B.n189 73.9501
R515 B.n398 B.n189 73.9501
R516 B.n398 B.n184 73.9501
R517 B.n404 B.n184 73.9501
R518 B.n404 B.n185 73.9501
R519 B.n411 B.n177 73.9501
R520 B.n417 B.n177 73.9501
R521 B.n417 B.n4 73.9501
R522 B.n504 B.n4 73.9501
R523 B.n504 B.n503 73.9501
R524 B.n503 B.n502 73.9501
R525 B.n502 B.n8 73.9501
R526 B.n12 B.n8 73.9501
R527 B.n495 B.n12 73.9501
R528 B.n494 B.n493 73.9501
R529 B.n493 B.n16 73.9501
R530 B.n487 B.n16 73.9501
R531 B.n487 B.n486 73.9501
R532 B.n486 B.n485 73.9501
R533 B.n485 B.n23 73.9501
R534 B.n479 B.n23 73.9501
R535 B.n479 B.n478 73.9501
R536 B.n478 B.n477 73.9501
R537 B.n477 B.n30 73.9501
R538 B.n471 B.n470 73.9501
R539 B.n470 B.n469 73.9501
R540 B.n469 B.n37 73.9501
R541 B.n463 B.n37 73.9501
R542 B.n463 B.n462 73.9501
R543 B.n462 B.n461 73.9501
R544 B.n461 B.n44 73.9501
R545 B.n75 B.t12 71.8703
R546 B.n250 B.t14 71.8703
R547 B.n78 B.t9 71.8655
R548 B.n247 B.t4 71.8655
R549 B.n456 B.n455 71.676
R550 B.n79 B.n48 71.676
R551 B.n83 B.n49 71.676
R552 B.n87 B.n50 71.676
R553 B.n91 B.n51 71.676
R554 B.n95 B.n52 71.676
R555 B.n99 B.n53 71.676
R556 B.n103 B.n54 71.676
R557 B.n107 B.n55 71.676
R558 B.n111 B.n56 71.676
R559 B.n115 B.n57 71.676
R560 B.n120 B.n58 71.676
R561 B.n124 B.n59 71.676
R562 B.n128 B.n60 71.676
R563 B.n132 B.n61 71.676
R564 B.n136 B.n62 71.676
R565 B.n140 B.n63 71.676
R566 B.n144 B.n64 71.676
R567 B.n148 B.n65 71.676
R568 B.n152 B.n66 71.676
R569 B.n156 B.n67 71.676
R570 B.n160 B.n68 71.676
R571 B.n164 B.n69 71.676
R572 B.n168 B.n70 71.676
R573 B.n172 B.n71 71.676
R574 B.n72 B.n71 71.676
R575 B.n171 B.n70 71.676
R576 B.n167 B.n69 71.676
R577 B.n163 B.n68 71.676
R578 B.n159 B.n67 71.676
R579 B.n155 B.n66 71.676
R580 B.n151 B.n65 71.676
R581 B.n147 B.n64 71.676
R582 B.n143 B.n63 71.676
R583 B.n139 B.n62 71.676
R584 B.n135 B.n61 71.676
R585 B.n131 B.n60 71.676
R586 B.n127 B.n59 71.676
R587 B.n123 B.n58 71.676
R588 B.n119 B.n57 71.676
R589 B.n114 B.n56 71.676
R590 B.n110 B.n55 71.676
R591 B.n106 B.n54 71.676
R592 B.n102 B.n53 71.676
R593 B.n98 B.n52 71.676
R594 B.n94 B.n51 71.676
R595 B.n90 B.n50 71.676
R596 B.n86 B.n49 71.676
R597 B.n82 B.n48 71.676
R598 B.n455 B.n47 71.676
R599 B.n351 B.n350 71.676
R600 B.n245 B.n221 71.676
R601 B.n343 B.n222 71.676
R602 B.n339 B.n223 71.676
R603 B.n335 B.n224 71.676
R604 B.n331 B.n225 71.676
R605 B.n327 B.n226 71.676
R606 B.n323 B.n227 71.676
R607 B.n319 B.n228 71.676
R608 B.n315 B.n229 71.676
R609 B.n311 B.n230 71.676
R610 B.n307 B.n231 71.676
R611 B.n303 B.n232 71.676
R612 B.n299 B.n233 71.676
R613 B.n295 B.n234 71.676
R614 B.n290 B.n235 71.676
R615 B.n286 B.n236 71.676
R616 B.n282 B.n237 71.676
R617 B.n278 B.n238 71.676
R618 B.n274 B.n239 71.676
R619 B.n270 B.n240 71.676
R620 B.n266 B.n241 71.676
R621 B.n262 B.n242 71.676
R622 B.n258 B.n243 71.676
R623 B.n254 B.n244 71.676
R624 B.n350 B.n220 71.676
R625 B.n344 B.n221 71.676
R626 B.n340 B.n222 71.676
R627 B.n336 B.n223 71.676
R628 B.n332 B.n224 71.676
R629 B.n328 B.n225 71.676
R630 B.n324 B.n226 71.676
R631 B.n320 B.n227 71.676
R632 B.n316 B.n228 71.676
R633 B.n312 B.n229 71.676
R634 B.n308 B.n230 71.676
R635 B.n304 B.n231 71.676
R636 B.n300 B.n232 71.676
R637 B.n296 B.n233 71.676
R638 B.n291 B.n234 71.676
R639 B.n287 B.n235 71.676
R640 B.n283 B.n236 71.676
R641 B.n279 B.n237 71.676
R642 B.n275 B.n238 71.676
R643 B.n271 B.n239 71.676
R644 B.n267 B.n240 71.676
R645 B.n263 B.n241 71.676
R646 B.n259 B.n242 71.676
R647 B.n255 B.n243 71.676
R648 B.n251 B.n244 71.676
R649 B.n506 B.n505 71.676
R650 B.n506 B.n2 71.676
R651 B.n411 B.t1 70.6876
R652 B.n495 B.t0 70.6876
R653 B.t3 B.n201 64.1626
R654 B.t7 B.n30 64.1626
R655 B.n117 B.n78 59.5399
R656 B.n76 B.n75 59.5399
R657 B.n293 B.n250 59.5399
R658 B.n248 B.n247 59.5399
R659 B.n78 B.n77 50.8126
R660 B.n75 B.n74 50.8126
R661 B.n250 B.n249 50.8126
R662 B.n247 B.n246 50.8126
R663 B.n353 B.n352 31.0639
R664 B.n252 B.n215 31.0639
R665 B.n452 B.n451 31.0639
R666 B.n458 B.n457 31.0639
R667 B B.n507 18.0485
R668 B.n354 B.n353 10.6151
R669 B.n354 B.n211 10.6151
R670 B.n364 B.n211 10.6151
R671 B.n365 B.n364 10.6151
R672 B.n366 B.n365 10.6151
R673 B.n366 B.n203 10.6151
R674 B.n376 B.n203 10.6151
R675 B.n377 B.n376 10.6151
R676 B.n378 B.n377 10.6151
R677 B.n378 B.n195 10.6151
R678 B.n388 B.n195 10.6151
R679 B.n389 B.n388 10.6151
R680 B.n390 B.n389 10.6151
R681 B.n390 B.n187 10.6151
R682 B.n400 B.n187 10.6151
R683 B.n401 B.n400 10.6151
R684 B.n402 B.n401 10.6151
R685 B.n402 B.n179 10.6151
R686 B.n413 B.n179 10.6151
R687 B.n414 B.n413 10.6151
R688 B.n415 B.n414 10.6151
R689 B.n415 B.n0 10.6151
R690 B.n352 B.n219 10.6151
R691 B.n347 B.n219 10.6151
R692 B.n347 B.n346 10.6151
R693 B.n346 B.n345 10.6151
R694 B.n345 B.n342 10.6151
R695 B.n342 B.n341 10.6151
R696 B.n341 B.n338 10.6151
R697 B.n338 B.n337 10.6151
R698 B.n337 B.n334 10.6151
R699 B.n334 B.n333 10.6151
R700 B.n333 B.n330 10.6151
R701 B.n330 B.n329 10.6151
R702 B.n329 B.n326 10.6151
R703 B.n326 B.n325 10.6151
R704 B.n325 B.n322 10.6151
R705 B.n322 B.n321 10.6151
R706 B.n321 B.n318 10.6151
R707 B.n318 B.n317 10.6151
R708 B.n317 B.n314 10.6151
R709 B.n314 B.n313 10.6151
R710 B.n310 B.n309 10.6151
R711 B.n309 B.n306 10.6151
R712 B.n306 B.n305 10.6151
R713 B.n305 B.n302 10.6151
R714 B.n302 B.n301 10.6151
R715 B.n301 B.n298 10.6151
R716 B.n298 B.n297 10.6151
R717 B.n297 B.n294 10.6151
R718 B.n292 B.n289 10.6151
R719 B.n289 B.n288 10.6151
R720 B.n288 B.n285 10.6151
R721 B.n285 B.n284 10.6151
R722 B.n284 B.n281 10.6151
R723 B.n281 B.n280 10.6151
R724 B.n280 B.n277 10.6151
R725 B.n277 B.n276 10.6151
R726 B.n276 B.n273 10.6151
R727 B.n273 B.n272 10.6151
R728 B.n272 B.n269 10.6151
R729 B.n269 B.n268 10.6151
R730 B.n268 B.n265 10.6151
R731 B.n265 B.n264 10.6151
R732 B.n264 B.n261 10.6151
R733 B.n261 B.n260 10.6151
R734 B.n260 B.n257 10.6151
R735 B.n257 B.n256 10.6151
R736 B.n256 B.n253 10.6151
R737 B.n253 B.n252 10.6151
R738 B.n358 B.n215 10.6151
R739 B.n359 B.n358 10.6151
R740 B.n360 B.n359 10.6151
R741 B.n360 B.n207 10.6151
R742 B.n370 B.n207 10.6151
R743 B.n371 B.n370 10.6151
R744 B.n372 B.n371 10.6151
R745 B.n372 B.n199 10.6151
R746 B.n382 B.n199 10.6151
R747 B.n383 B.n382 10.6151
R748 B.n384 B.n383 10.6151
R749 B.n384 B.n191 10.6151
R750 B.n394 B.n191 10.6151
R751 B.n395 B.n394 10.6151
R752 B.n396 B.n395 10.6151
R753 B.n396 B.n182 10.6151
R754 B.n406 B.n182 10.6151
R755 B.n407 B.n406 10.6151
R756 B.n409 B.n407 10.6151
R757 B.n409 B.n408 10.6151
R758 B.n408 B.n175 10.6151
R759 B.n420 B.n175 10.6151
R760 B.n421 B.n420 10.6151
R761 B.n422 B.n421 10.6151
R762 B.n423 B.n422 10.6151
R763 B.n424 B.n423 10.6151
R764 B.n427 B.n424 10.6151
R765 B.n428 B.n427 10.6151
R766 B.n429 B.n428 10.6151
R767 B.n430 B.n429 10.6151
R768 B.n432 B.n430 10.6151
R769 B.n433 B.n432 10.6151
R770 B.n434 B.n433 10.6151
R771 B.n435 B.n434 10.6151
R772 B.n437 B.n435 10.6151
R773 B.n438 B.n437 10.6151
R774 B.n439 B.n438 10.6151
R775 B.n440 B.n439 10.6151
R776 B.n442 B.n440 10.6151
R777 B.n443 B.n442 10.6151
R778 B.n444 B.n443 10.6151
R779 B.n445 B.n444 10.6151
R780 B.n447 B.n445 10.6151
R781 B.n448 B.n447 10.6151
R782 B.n449 B.n448 10.6151
R783 B.n450 B.n449 10.6151
R784 B.n451 B.n450 10.6151
R785 B.n499 B.n1 10.6151
R786 B.n499 B.n498 10.6151
R787 B.n498 B.n497 10.6151
R788 B.n497 B.n10 10.6151
R789 B.n491 B.n10 10.6151
R790 B.n491 B.n490 10.6151
R791 B.n490 B.n489 10.6151
R792 B.n489 B.n18 10.6151
R793 B.n483 B.n18 10.6151
R794 B.n483 B.n482 10.6151
R795 B.n482 B.n481 10.6151
R796 B.n481 B.n25 10.6151
R797 B.n475 B.n25 10.6151
R798 B.n475 B.n474 10.6151
R799 B.n474 B.n473 10.6151
R800 B.n473 B.n32 10.6151
R801 B.n467 B.n32 10.6151
R802 B.n467 B.n466 10.6151
R803 B.n466 B.n465 10.6151
R804 B.n465 B.n39 10.6151
R805 B.n459 B.n39 10.6151
R806 B.n459 B.n458 10.6151
R807 B.n457 B.n46 10.6151
R808 B.n80 B.n46 10.6151
R809 B.n81 B.n80 10.6151
R810 B.n84 B.n81 10.6151
R811 B.n85 B.n84 10.6151
R812 B.n88 B.n85 10.6151
R813 B.n89 B.n88 10.6151
R814 B.n92 B.n89 10.6151
R815 B.n93 B.n92 10.6151
R816 B.n96 B.n93 10.6151
R817 B.n97 B.n96 10.6151
R818 B.n100 B.n97 10.6151
R819 B.n101 B.n100 10.6151
R820 B.n104 B.n101 10.6151
R821 B.n105 B.n104 10.6151
R822 B.n108 B.n105 10.6151
R823 B.n109 B.n108 10.6151
R824 B.n112 B.n109 10.6151
R825 B.n113 B.n112 10.6151
R826 B.n116 B.n113 10.6151
R827 B.n121 B.n118 10.6151
R828 B.n122 B.n121 10.6151
R829 B.n125 B.n122 10.6151
R830 B.n126 B.n125 10.6151
R831 B.n129 B.n126 10.6151
R832 B.n130 B.n129 10.6151
R833 B.n133 B.n130 10.6151
R834 B.n134 B.n133 10.6151
R835 B.n138 B.n137 10.6151
R836 B.n141 B.n138 10.6151
R837 B.n142 B.n141 10.6151
R838 B.n145 B.n142 10.6151
R839 B.n146 B.n145 10.6151
R840 B.n149 B.n146 10.6151
R841 B.n150 B.n149 10.6151
R842 B.n153 B.n150 10.6151
R843 B.n154 B.n153 10.6151
R844 B.n157 B.n154 10.6151
R845 B.n158 B.n157 10.6151
R846 B.n161 B.n158 10.6151
R847 B.n162 B.n161 10.6151
R848 B.n165 B.n162 10.6151
R849 B.n166 B.n165 10.6151
R850 B.n169 B.n166 10.6151
R851 B.n170 B.n169 10.6151
R852 B.n173 B.n170 10.6151
R853 B.n174 B.n173 10.6151
R854 B.n452 B.n174 10.6151
R855 B.n374 B.t3 9.78794
R856 B.n471 B.t7 9.78794
R857 B.n507 B.n0 8.11757
R858 B.n507 B.n1 8.11757
R859 B.n310 B.n248 6.5566
R860 B.n294 B.n293 6.5566
R861 B.n118 B.n117 6.5566
R862 B.n134 B.n76 6.5566
R863 B.n313 B.n248 4.05904
R864 B.n293 B.n292 4.05904
R865 B.n117 B.n116 4.05904
R866 B.n137 B.n76 4.05904
R867 B.n185 B.t1 3.26298
R868 B.t0 B.n494 3.26298
R869 VP.n0 VP.t1 138.561
R870 VP.n0 VP.t0 100.151
R871 VP VP.n0 0.336784
R872 VTAIL.n1 VTAIL.t0 55.4276
R873 VTAIL.n3 VTAIL.t1 55.4275
R874 VTAIL.n0 VTAIL.t2 55.4275
R875 VTAIL.n2 VTAIL.t3 55.4275
R876 VTAIL.n1 VTAIL.n0 21.0565
R877 VTAIL.n3 VTAIL.n2 18.7979
R878 VTAIL.n2 VTAIL.n1 1.59964
R879 VTAIL VTAIL.n0 1.09317
R880 VTAIL VTAIL.n3 0.506965
R881 VDD1 VDD1.t1 105.544
R882 VDD1 VDD1.t0 72.7292
R883 VN VN.t0 138.659
R884 VN VN.t1 100.489
R885 VDD2.n0 VDD2.t0 104.456
R886 VDD2.n0 VDD2.t1 72.1063
R887 VDD2 VDD2.n0 0.623345
C0 VP VTAIL 1.31397f
C1 VDD2 VDD1 0.636626f
C2 VN VDD1 0.152138f
C3 VDD2 VTAIL 3.14514f
C4 VN VTAIL 1.29978f
C5 VP VDD2 0.323902f
C6 VN VP 3.98284f
C7 VN VDD2 1.2495f
C8 VTAIL VDD1 3.09509f
C9 VP VDD1 1.4196f
C10 VDD2 B 2.994374f
C11 VDD1 B 4.79681f
C12 VTAIL B 4.120655f
C13 VN B 7.43062f
C14 VP B 5.403826f
C15 VDD2.t0 B 0.824059f
C16 VDD2.t1 B 0.586603f
C17 VDD2.n0 B 1.60463f
C18 VN.t1 B 0.865952f
C19 VN.t0 B 1.17514f
C20 VDD1.t0 B 0.57792f
C21 VDD1.t1 B 0.829366f
C22 VTAIL.t2 B 0.617859f
C23 VTAIL.n0 B 0.966285f
C24 VTAIL.t0 B 0.617863f
C25 VTAIL.n1 B 0.994045f
C26 VTAIL.t3 B 0.617859f
C27 VTAIL.n2 B 0.870233f
C28 VTAIL.t1 B 0.617859f
C29 VTAIL.n3 B 0.810333f
C30 VP.t1 B 1.18171f
C31 VP.t0 B 0.872061f
C32 VP.n0 B 1.8971f
.ends

