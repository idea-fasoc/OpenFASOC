* NGSPICE file created from diff_pair_sample_0570.ext - technology: sky130A

.subckt diff_pair_sample_0570 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.08735 pd=6.92 as=2.5701 ps=13.96 w=6.59 l=3.77
X1 VDD1.t3 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.08735 pd=6.92 as=2.5701 ps=13.96 w=6.59 l=3.77
X2 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=2.5701 pd=13.96 as=0 ps=0 w=6.59 l=3.77
X3 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=2.5701 pd=13.96 as=0 ps=0 w=6.59 l=3.77
X4 VTAIL.t2 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.5701 pd=13.96 as=1.08735 ps=6.92 w=6.59 l=3.77
X5 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5701 pd=13.96 as=0 ps=0 w=6.59 l=3.77
X6 VDD2.t2 VN.t1 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.08735 pd=6.92 as=2.5701 ps=13.96 w=6.59 l=3.77
X7 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5701 pd=13.96 as=0 ps=0 w=6.59 l=3.77
X8 VDD1.t1 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.08735 pd=6.92 as=2.5701 ps=13.96 w=6.59 l=3.77
X9 VTAIL.t4 VN.t2 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.5701 pd=13.96 as=1.08735 ps=6.92 w=6.59 l=3.77
X10 VTAIL.t1 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5701 pd=13.96 as=1.08735 ps=6.92 w=6.59 l=3.77
X11 VTAIL.t7 VN.t3 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5701 pd=13.96 as=1.08735 ps=6.92 w=6.59 l=3.77
R0 VN.n1 VN.t1 75.8784
R1 VN.n0 VN.t3 75.8784
R2 VN.n0 VN.t0 74.5357
R3 VN.n1 VN.t2 74.5357
R4 VN VN.n1 47.8771
R5 VN VN.n0 1.88085
R6 VTAIL.n270 VTAIL.n269 289.615
R7 VTAIL.n32 VTAIL.n31 289.615
R8 VTAIL.n66 VTAIL.n65 289.615
R9 VTAIL.n100 VTAIL.n99 289.615
R10 VTAIL.n236 VTAIL.n235 289.615
R11 VTAIL.n202 VTAIL.n201 289.615
R12 VTAIL.n168 VTAIL.n167 289.615
R13 VTAIL.n134 VTAIL.n133 289.615
R14 VTAIL.n248 VTAIL.n247 185
R15 VTAIL.n253 VTAIL.n252 185
R16 VTAIL.n255 VTAIL.n254 185
R17 VTAIL.n244 VTAIL.n243 185
R18 VTAIL.n261 VTAIL.n260 185
R19 VTAIL.n263 VTAIL.n262 185
R20 VTAIL.n240 VTAIL.n239 185
R21 VTAIL.n269 VTAIL.n268 185
R22 VTAIL.n10 VTAIL.n9 185
R23 VTAIL.n15 VTAIL.n14 185
R24 VTAIL.n17 VTAIL.n16 185
R25 VTAIL.n6 VTAIL.n5 185
R26 VTAIL.n23 VTAIL.n22 185
R27 VTAIL.n25 VTAIL.n24 185
R28 VTAIL.n2 VTAIL.n1 185
R29 VTAIL.n31 VTAIL.n30 185
R30 VTAIL.n44 VTAIL.n43 185
R31 VTAIL.n49 VTAIL.n48 185
R32 VTAIL.n51 VTAIL.n50 185
R33 VTAIL.n40 VTAIL.n39 185
R34 VTAIL.n57 VTAIL.n56 185
R35 VTAIL.n59 VTAIL.n58 185
R36 VTAIL.n36 VTAIL.n35 185
R37 VTAIL.n65 VTAIL.n64 185
R38 VTAIL.n78 VTAIL.n77 185
R39 VTAIL.n83 VTAIL.n82 185
R40 VTAIL.n85 VTAIL.n84 185
R41 VTAIL.n74 VTAIL.n73 185
R42 VTAIL.n91 VTAIL.n90 185
R43 VTAIL.n93 VTAIL.n92 185
R44 VTAIL.n70 VTAIL.n69 185
R45 VTAIL.n99 VTAIL.n98 185
R46 VTAIL.n235 VTAIL.n234 185
R47 VTAIL.n206 VTAIL.n205 185
R48 VTAIL.n229 VTAIL.n228 185
R49 VTAIL.n227 VTAIL.n226 185
R50 VTAIL.n210 VTAIL.n209 185
R51 VTAIL.n221 VTAIL.n220 185
R52 VTAIL.n219 VTAIL.n218 185
R53 VTAIL.n214 VTAIL.n213 185
R54 VTAIL.n201 VTAIL.n200 185
R55 VTAIL.n172 VTAIL.n171 185
R56 VTAIL.n195 VTAIL.n194 185
R57 VTAIL.n193 VTAIL.n192 185
R58 VTAIL.n176 VTAIL.n175 185
R59 VTAIL.n187 VTAIL.n186 185
R60 VTAIL.n185 VTAIL.n184 185
R61 VTAIL.n180 VTAIL.n179 185
R62 VTAIL.n167 VTAIL.n166 185
R63 VTAIL.n138 VTAIL.n137 185
R64 VTAIL.n161 VTAIL.n160 185
R65 VTAIL.n159 VTAIL.n158 185
R66 VTAIL.n142 VTAIL.n141 185
R67 VTAIL.n153 VTAIL.n152 185
R68 VTAIL.n151 VTAIL.n150 185
R69 VTAIL.n146 VTAIL.n145 185
R70 VTAIL.n133 VTAIL.n132 185
R71 VTAIL.n104 VTAIL.n103 185
R72 VTAIL.n127 VTAIL.n126 185
R73 VTAIL.n125 VTAIL.n124 185
R74 VTAIL.n108 VTAIL.n107 185
R75 VTAIL.n119 VTAIL.n118 185
R76 VTAIL.n117 VTAIL.n116 185
R77 VTAIL.n112 VTAIL.n111 185
R78 VTAIL.n181 VTAIL.t1 149.525
R79 VTAIL.n147 VTAIL.t6 149.525
R80 VTAIL.n113 VTAIL.t4 149.525
R81 VTAIL.n249 VTAIL.t5 149.525
R82 VTAIL.n11 VTAIL.t7 149.525
R83 VTAIL.n45 VTAIL.t3 149.525
R84 VTAIL.n79 VTAIL.t2 149.525
R85 VTAIL.n215 VTAIL.t0 149.525
R86 VTAIL.n253 VTAIL.n247 104.615
R87 VTAIL.n254 VTAIL.n253 104.615
R88 VTAIL.n254 VTAIL.n243 104.615
R89 VTAIL.n261 VTAIL.n243 104.615
R90 VTAIL.n262 VTAIL.n261 104.615
R91 VTAIL.n262 VTAIL.n239 104.615
R92 VTAIL.n269 VTAIL.n239 104.615
R93 VTAIL.n15 VTAIL.n9 104.615
R94 VTAIL.n16 VTAIL.n15 104.615
R95 VTAIL.n16 VTAIL.n5 104.615
R96 VTAIL.n23 VTAIL.n5 104.615
R97 VTAIL.n24 VTAIL.n23 104.615
R98 VTAIL.n24 VTAIL.n1 104.615
R99 VTAIL.n31 VTAIL.n1 104.615
R100 VTAIL.n49 VTAIL.n43 104.615
R101 VTAIL.n50 VTAIL.n49 104.615
R102 VTAIL.n50 VTAIL.n39 104.615
R103 VTAIL.n57 VTAIL.n39 104.615
R104 VTAIL.n58 VTAIL.n57 104.615
R105 VTAIL.n58 VTAIL.n35 104.615
R106 VTAIL.n65 VTAIL.n35 104.615
R107 VTAIL.n83 VTAIL.n77 104.615
R108 VTAIL.n84 VTAIL.n83 104.615
R109 VTAIL.n84 VTAIL.n73 104.615
R110 VTAIL.n91 VTAIL.n73 104.615
R111 VTAIL.n92 VTAIL.n91 104.615
R112 VTAIL.n92 VTAIL.n69 104.615
R113 VTAIL.n99 VTAIL.n69 104.615
R114 VTAIL.n235 VTAIL.n205 104.615
R115 VTAIL.n228 VTAIL.n205 104.615
R116 VTAIL.n228 VTAIL.n227 104.615
R117 VTAIL.n227 VTAIL.n209 104.615
R118 VTAIL.n220 VTAIL.n209 104.615
R119 VTAIL.n220 VTAIL.n219 104.615
R120 VTAIL.n219 VTAIL.n213 104.615
R121 VTAIL.n201 VTAIL.n171 104.615
R122 VTAIL.n194 VTAIL.n171 104.615
R123 VTAIL.n194 VTAIL.n193 104.615
R124 VTAIL.n193 VTAIL.n175 104.615
R125 VTAIL.n186 VTAIL.n175 104.615
R126 VTAIL.n186 VTAIL.n185 104.615
R127 VTAIL.n185 VTAIL.n179 104.615
R128 VTAIL.n167 VTAIL.n137 104.615
R129 VTAIL.n160 VTAIL.n137 104.615
R130 VTAIL.n160 VTAIL.n159 104.615
R131 VTAIL.n159 VTAIL.n141 104.615
R132 VTAIL.n152 VTAIL.n141 104.615
R133 VTAIL.n152 VTAIL.n151 104.615
R134 VTAIL.n151 VTAIL.n145 104.615
R135 VTAIL.n133 VTAIL.n103 104.615
R136 VTAIL.n126 VTAIL.n103 104.615
R137 VTAIL.n126 VTAIL.n125 104.615
R138 VTAIL.n125 VTAIL.n107 104.615
R139 VTAIL.n118 VTAIL.n107 104.615
R140 VTAIL.n118 VTAIL.n117 104.615
R141 VTAIL.n117 VTAIL.n111 104.615
R142 VTAIL.t5 VTAIL.n247 52.3082
R143 VTAIL.t7 VTAIL.n9 52.3082
R144 VTAIL.t3 VTAIL.n43 52.3082
R145 VTAIL.t2 VTAIL.n77 52.3082
R146 VTAIL.t0 VTAIL.n213 52.3082
R147 VTAIL.t1 VTAIL.n179 52.3082
R148 VTAIL.t6 VTAIL.n145 52.3082
R149 VTAIL.t4 VTAIL.n111 52.3082
R150 VTAIL.n271 VTAIL.n270 36.2581
R151 VTAIL.n33 VTAIL.n32 36.2581
R152 VTAIL.n67 VTAIL.n66 36.2581
R153 VTAIL.n101 VTAIL.n100 36.2581
R154 VTAIL.n237 VTAIL.n236 36.2581
R155 VTAIL.n203 VTAIL.n202 36.2581
R156 VTAIL.n169 VTAIL.n168 36.2581
R157 VTAIL.n135 VTAIL.n134 36.2581
R158 VTAIL.n271 VTAIL.n237 21.5824
R159 VTAIL.n135 VTAIL.n101 21.5824
R160 VTAIL.n268 VTAIL.n238 12.8005
R161 VTAIL.n30 VTAIL.n0 12.8005
R162 VTAIL.n64 VTAIL.n34 12.8005
R163 VTAIL.n98 VTAIL.n68 12.8005
R164 VTAIL.n234 VTAIL.n204 12.8005
R165 VTAIL.n200 VTAIL.n170 12.8005
R166 VTAIL.n166 VTAIL.n136 12.8005
R167 VTAIL.n132 VTAIL.n102 12.8005
R168 VTAIL.n267 VTAIL.n240 12.0247
R169 VTAIL.n29 VTAIL.n2 12.0247
R170 VTAIL.n63 VTAIL.n36 12.0247
R171 VTAIL.n97 VTAIL.n70 12.0247
R172 VTAIL.n233 VTAIL.n206 12.0247
R173 VTAIL.n199 VTAIL.n172 12.0247
R174 VTAIL.n165 VTAIL.n138 12.0247
R175 VTAIL.n131 VTAIL.n104 12.0247
R176 VTAIL.n264 VTAIL.n263 11.249
R177 VTAIL.n26 VTAIL.n25 11.249
R178 VTAIL.n60 VTAIL.n59 11.249
R179 VTAIL.n94 VTAIL.n93 11.249
R180 VTAIL.n230 VTAIL.n229 11.249
R181 VTAIL.n196 VTAIL.n195 11.249
R182 VTAIL.n162 VTAIL.n161 11.249
R183 VTAIL.n128 VTAIL.n127 11.249
R184 VTAIL.n260 VTAIL.n242 10.4732
R185 VTAIL.n22 VTAIL.n4 10.4732
R186 VTAIL.n56 VTAIL.n38 10.4732
R187 VTAIL.n90 VTAIL.n72 10.4732
R188 VTAIL.n226 VTAIL.n208 10.4732
R189 VTAIL.n192 VTAIL.n174 10.4732
R190 VTAIL.n158 VTAIL.n140 10.4732
R191 VTAIL.n124 VTAIL.n106 10.4732
R192 VTAIL.n249 VTAIL.n248 10.2746
R193 VTAIL.n11 VTAIL.n10 10.2746
R194 VTAIL.n45 VTAIL.n44 10.2746
R195 VTAIL.n79 VTAIL.n78 10.2746
R196 VTAIL.n215 VTAIL.n214 10.2746
R197 VTAIL.n181 VTAIL.n180 10.2746
R198 VTAIL.n147 VTAIL.n146 10.2746
R199 VTAIL.n113 VTAIL.n112 10.2746
R200 VTAIL.n259 VTAIL.n244 9.69747
R201 VTAIL.n21 VTAIL.n6 9.69747
R202 VTAIL.n55 VTAIL.n40 9.69747
R203 VTAIL.n89 VTAIL.n74 9.69747
R204 VTAIL.n225 VTAIL.n210 9.69747
R205 VTAIL.n191 VTAIL.n176 9.69747
R206 VTAIL.n157 VTAIL.n142 9.69747
R207 VTAIL.n123 VTAIL.n108 9.69747
R208 VTAIL.n266 VTAIL.n238 9.45567
R209 VTAIL.n28 VTAIL.n0 9.45567
R210 VTAIL.n62 VTAIL.n34 9.45567
R211 VTAIL.n96 VTAIL.n68 9.45567
R212 VTAIL.n232 VTAIL.n204 9.45567
R213 VTAIL.n198 VTAIL.n170 9.45567
R214 VTAIL.n164 VTAIL.n136 9.45567
R215 VTAIL.n130 VTAIL.n102 9.45567
R216 VTAIL.n251 VTAIL.n250 9.3005
R217 VTAIL.n246 VTAIL.n245 9.3005
R218 VTAIL.n257 VTAIL.n256 9.3005
R219 VTAIL.n259 VTAIL.n258 9.3005
R220 VTAIL.n242 VTAIL.n241 9.3005
R221 VTAIL.n265 VTAIL.n264 9.3005
R222 VTAIL.n267 VTAIL.n266 9.3005
R223 VTAIL.n13 VTAIL.n12 9.3005
R224 VTAIL.n8 VTAIL.n7 9.3005
R225 VTAIL.n19 VTAIL.n18 9.3005
R226 VTAIL.n21 VTAIL.n20 9.3005
R227 VTAIL.n4 VTAIL.n3 9.3005
R228 VTAIL.n27 VTAIL.n26 9.3005
R229 VTAIL.n29 VTAIL.n28 9.3005
R230 VTAIL.n47 VTAIL.n46 9.3005
R231 VTAIL.n42 VTAIL.n41 9.3005
R232 VTAIL.n53 VTAIL.n52 9.3005
R233 VTAIL.n55 VTAIL.n54 9.3005
R234 VTAIL.n38 VTAIL.n37 9.3005
R235 VTAIL.n61 VTAIL.n60 9.3005
R236 VTAIL.n63 VTAIL.n62 9.3005
R237 VTAIL.n81 VTAIL.n80 9.3005
R238 VTAIL.n76 VTAIL.n75 9.3005
R239 VTAIL.n87 VTAIL.n86 9.3005
R240 VTAIL.n89 VTAIL.n88 9.3005
R241 VTAIL.n72 VTAIL.n71 9.3005
R242 VTAIL.n95 VTAIL.n94 9.3005
R243 VTAIL.n97 VTAIL.n96 9.3005
R244 VTAIL.n233 VTAIL.n232 9.3005
R245 VTAIL.n231 VTAIL.n230 9.3005
R246 VTAIL.n208 VTAIL.n207 9.3005
R247 VTAIL.n225 VTAIL.n224 9.3005
R248 VTAIL.n223 VTAIL.n222 9.3005
R249 VTAIL.n212 VTAIL.n211 9.3005
R250 VTAIL.n217 VTAIL.n216 9.3005
R251 VTAIL.n178 VTAIL.n177 9.3005
R252 VTAIL.n189 VTAIL.n188 9.3005
R253 VTAIL.n191 VTAIL.n190 9.3005
R254 VTAIL.n174 VTAIL.n173 9.3005
R255 VTAIL.n197 VTAIL.n196 9.3005
R256 VTAIL.n199 VTAIL.n198 9.3005
R257 VTAIL.n183 VTAIL.n182 9.3005
R258 VTAIL.n144 VTAIL.n143 9.3005
R259 VTAIL.n155 VTAIL.n154 9.3005
R260 VTAIL.n157 VTAIL.n156 9.3005
R261 VTAIL.n140 VTAIL.n139 9.3005
R262 VTAIL.n163 VTAIL.n162 9.3005
R263 VTAIL.n165 VTAIL.n164 9.3005
R264 VTAIL.n149 VTAIL.n148 9.3005
R265 VTAIL.n110 VTAIL.n109 9.3005
R266 VTAIL.n121 VTAIL.n120 9.3005
R267 VTAIL.n123 VTAIL.n122 9.3005
R268 VTAIL.n106 VTAIL.n105 9.3005
R269 VTAIL.n129 VTAIL.n128 9.3005
R270 VTAIL.n131 VTAIL.n130 9.3005
R271 VTAIL.n115 VTAIL.n114 9.3005
R272 VTAIL.n256 VTAIL.n255 8.92171
R273 VTAIL.n18 VTAIL.n17 8.92171
R274 VTAIL.n52 VTAIL.n51 8.92171
R275 VTAIL.n86 VTAIL.n85 8.92171
R276 VTAIL.n222 VTAIL.n221 8.92171
R277 VTAIL.n188 VTAIL.n187 8.92171
R278 VTAIL.n154 VTAIL.n153 8.92171
R279 VTAIL.n120 VTAIL.n119 8.92171
R280 VTAIL.n252 VTAIL.n246 8.14595
R281 VTAIL.n14 VTAIL.n8 8.14595
R282 VTAIL.n48 VTAIL.n42 8.14595
R283 VTAIL.n82 VTAIL.n76 8.14595
R284 VTAIL.n218 VTAIL.n212 8.14595
R285 VTAIL.n184 VTAIL.n178 8.14595
R286 VTAIL.n150 VTAIL.n144 8.14595
R287 VTAIL.n116 VTAIL.n110 8.14595
R288 VTAIL.n251 VTAIL.n248 7.3702
R289 VTAIL.n13 VTAIL.n10 7.3702
R290 VTAIL.n47 VTAIL.n44 7.3702
R291 VTAIL.n81 VTAIL.n78 7.3702
R292 VTAIL.n217 VTAIL.n214 7.3702
R293 VTAIL.n183 VTAIL.n180 7.3702
R294 VTAIL.n149 VTAIL.n146 7.3702
R295 VTAIL.n115 VTAIL.n112 7.3702
R296 VTAIL.n252 VTAIL.n251 5.81868
R297 VTAIL.n14 VTAIL.n13 5.81868
R298 VTAIL.n48 VTAIL.n47 5.81868
R299 VTAIL.n82 VTAIL.n81 5.81868
R300 VTAIL.n218 VTAIL.n217 5.81868
R301 VTAIL.n184 VTAIL.n183 5.81868
R302 VTAIL.n150 VTAIL.n149 5.81868
R303 VTAIL.n116 VTAIL.n115 5.81868
R304 VTAIL.n255 VTAIL.n246 5.04292
R305 VTAIL.n17 VTAIL.n8 5.04292
R306 VTAIL.n51 VTAIL.n42 5.04292
R307 VTAIL.n85 VTAIL.n76 5.04292
R308 VTAIL.n221 VTAIL.n212 5.04292
R309 VTAIL.n187 VTAIL.n178 5.04292
R310 VTAIL.n153 VTAIL.n144 5.04292
R311 VTAIL.n119 VTAIL.n110 5.04292
R312 VTAIL.n256 VTAIL.n244 4.26717
R313 VTAIL.n18 VTAIL.n6 4.26717
R314 VTAIL.n52 VTAIL.n40 4.26717
R315 VTAIL.n86 VTAIL.n74 4.26717
R316 VTAIL.n222 VTAIL.n210 4.26717
R317 VTAIL.n188 VTAIL.n176 4.26717
R318 VTAIL.n154 VTAIL.n142 4.26717
R319 VTAIL.n120 VTAIL.n108 4.26717
R320 VTAIL.n169 VTAIL.n135 3.53498
R321 VTAIL.n237 VTAIL.n203 3.53498
R322 VTAIL.n101 VTAIL.n67 3.53498
R323 VTAIL.n260 VTAIL.n259 3.49141
R324 VTAIL.n22 VTAIL.n21 3.49141
R325 VTAIL.n56 VTAIL.n55 3.49141
R326 VTAIL.n90 VTAIL.n89 3.49141
R327 VTAIL.n226 VTAIL.n225 3.49141
R328 VTAIL.n192 VTAIL.n191 3.49141
R329 VTAIL.n158 VTAIL.n157 3.49141
R330 VTAIL.n124 VTAIL.n123 3.49141
R331 VTAIL.n182 VTAIL.n181 2.84308
R332 VTAIL.n148 VTAIL.n147 2.84308
R333 VTAIL.n114 VTAIL.n113 2.84308
R334 VTAIL.n250 VTAIL.n249 2.84308
R335 VTAIL.n12 VTAIL.n11 2.84308
R336 VTAIL.n46 VTAIL.n45 2.84308
R337 VTAIL.n80 VTAIL.n79 2.84308
R338 VTAIL.n216 VTAIL.n215 2.84308
R339 VTAIL.n263 VTAIL.n242 2.71565
R340 VTAIL.n25 VTAIL.n4 2.71565
R341 VTAIL.n59 VTAIL.n38 2.71565
R342 VTAIL.n93 VTAIL.n72 2.71565
R343 VTAIL.n229 VTAIL.n208 2.71565
R344 VTAIL.n195 VTAIL.n174 2.71565
R345 VTAIL.n161 VTAIL.n140 2.71565
R346 VTAIL.n127 VTAIL.n106 2.71565
R347 VTAIL.n264 VTAIL.n240 1.93989
R348 VTAIL.n26 VTAIL.n2 1.93989
R349 VTAIL.n60 VTAIL.n36 1.93989
R350 VTAIL.n94 VTAIL.n70 1.93989
R351 VTAIL.n230 VTAIL.n206 1.93989
R352 VTAIL.n196 VTAIL.n172 1.93989
R353 VTAIL.n162 VTAIL.n138 1.93989
R354 VTAIL.n128 VTAIL.n104 1.93989
R355 VTAIL VTAIL.n33 1.82593
R356 VTAIL VTAIL.n271 1.70955
R357 VTAIL.n268 VTAIL.n267 1.16414
R358 VTAIL.n30 VTAIL.n29 1.16414
R359 VTAIL.n64 VTAIL.n63 1.16414
R360 VTAIL.n98 VTAIL.n97 1.16414
R361 VTAIL.n234 VTAIL.n233 1.16414
R362 VTAIL.n200 VTAIL.n199 1.16414
R363 VTAIL.n166 VTAIL.n165 1.16414
R364 VTAIL.n132 VTAIL.n131 1.16414
R365 VTAIL.n203 VTAIL.n169 0.470328
R366 VTAIL.n67 VTAIL.n33 0.470328
R367 VTAIL.n270 VTAIL.n238 0.388379
R368 VTAIL.n32 VTAIL.n0 0.388379
R369 VTAIL.n66 VTAIL.n34 0.388379
R370 VTAIL.n100 VTAIL.n68 0.388379
R371 VTAIL.n236 VTAIL.n204 0.388379
R372 VTAIL.n202 VTAIL.n170 0.388379
R373 VTAIL.n168 VTAIL.n136 0.388379
R374 VTAIL.n134 VTAIL.n102 0.388379
R375 VTAIL.n250 VTAIL.n245 0.155672
R376 VTAIL.n257 VTAIL.n245 0.155672
R377 VTAIL.n258 VTAIL.n257 0.155672
R378 VTAIL.n258 VTAIL.n241 0.155672
R379 VTAIL.n265 VTAIL.n241 0.155672
R380 VTAIL.n266 VTAIL.n265 0.155672
R381 VTAIL.n12 VTAIL.n7 0.155672
R382 VTAIL.n19 VTAIL.n7 0.155672
R383 VTAIL.n20 VTAIL.n19 0.155672
R384 VTAIL.n20 VTAIL.n3 0.155672
R385 VTAIL.n27 VTAIL.n3 0.155672
R386 VTAIL.n28 VTAIL.n27 0.155672
R387 VTAIL.n46 VTAIL.n41 0.155672
R388 VTAIL.n53 VTAIL.n41 0.155672
R389 VTAIL.n54 VTAIL.n53 0.155672
R390 VTAIL.n54 VTAIL.n37 0.155672
R391 VTAIL.n61 VTAIL.n37 0.155672
R392 VTAIL.n62 VTAIL.n61 0.155672
R393 VTAIL.n80 VTAIL.n75 0.155672
R394 VTAIL.n87 VTAIL.n75 0.155672
R395 VTAIL.n88 VTAIL.n87 0.155672
R396 VTAIL.n88 VTAIL.n71 0.155672
R397 VTAIL.n95 VTAIL.n71 0.155672
R398 VTAIL.n96 VTAIL.n95 0.155672
R399 VTAIL.n232 VTAIL.n231 0.155672
R400 VTAIL.n231 VTAIL.n207 0.155672
R401 VTAIL.n224 VTAIL.n207 0.155672
R402 VTAIL.n224 VTAIL.n223 0.155672
R403 VTAIL.n223 VTAIL.n211 0.155672
R404 VTAIL.n216 VTAIL.n211 0.155672
R405 VTAIL.n198 VTAIL.n197 0.155672
R406 VTAIL.n197 VTAIL.n173 0.155672
R407 VTAIL.n190 VTAIL.n173 0.155672
R408 VTAIL.n190 VTAIL.n189 0.155672
R409 VTAIL.n189 VTAIL.n177 0.155672
R410 VTAIL.n182 VTAIL.n177 0.155672
R411 VTAIL.n164 VTAIL.n163 0.155672
R412 VTAIL.n163 VTAIL.n139 0.155672
R413 VTAIL.n156 VTAIL.n139 0.155672
R414 VTAIL.n156 VTAIL.n155 0.155672
R415 VTAIL.n155 VTAIL.n143 0.155672
R416 VTAIL.n148 VTAIL.n143 0.155672
R417 VTAIL.n130 VTAIL.n129 0.155672
R418 VTAIL.n129 VTAIL.n105 0.155672
R419 VTAIL.n122 VTAIL.n105 0.155672
R420 VTAIL.n122 VTAIL.n121 0.155672
R421 VTAIL.n121 VTAIL.n109 0.155672
R422 VTAIL.n114 VTAIL.n109 0.155672
R423 VDD2.n2 VDD2.n0 109.873
R424 VDD2.n2 VDD2.n1 69.8735
R425 VDD2.n1 VDD2.t1 3.00505
R426 VDD2.n1 VDD2.t2 3.00505
R427 VDD2.n0 VDD2.t0 3.00505
R428 VDD2.n0 VDD2.t3 3.00505
R429 VDD2 VDD2.n2 0.0586897
R430 B.n673 B.n672 585
R431 B.n674 B.n673 585
R432 B.n237 B.n114 585
R433 B.n236 B.n235 585
R434 B.n234 B.n233 585
R435 B.n232 B.n231 585
R436 B.n230 B.n229 585
R437 B.n228 B.n227 585
R438 B.n226 B.n225 585
R439 B.n224 B.n223 585
R440 B.n222 B.n221 585
R441 B.n220 B.n219 585
R442 B.n218 B.n217 585
R443 B.n216 B.n215 585
R444 B.n214 B.n213 585
R445 B.n212 B.n211 585
R446 B.n210 B.n209 585
R447 B.n208 B.n207 585
R448 B.n206 B.n205 585
R449 B.n204 B.n203 585
R450 B.n202 B.n201 585
R451 B.n200 B.n199 585
R452 B.n198 B.n197 585
R453 B.n196 B.n195 585
R454 B.n194 B.n193 585
R455 B.n192 B.n191 585
R456 B.n190 B.n189 585
R457 B.n187 B.n186 585
R458 B.n185 B.n184 585
R459 B.n183 B.n182 585
R460 B.n181 B.n180 585
R461 B.n179 B.n178 585
R462 B.n177 B.n176 585
R463 B.n175 B.n174 585
R464 B.n173 B.n172 585
R465 B.n171 B.n170 585
R466 B.n169 B.n168 585
R467 B.n167 B.n166 585
R468 B.n165 B.n164 585
R469 B.n163 B.n162 585
R470 B.n161 B.n160 585
R471 B.n159 B.n158 585
R472 B.n157 B.n156 585
R473 B.n155 B.n154 585
R474 B.n153 B.n152 585
R475 B.n151 B.n150 585
R476 B.n149 B.n148 585
R477 B.n147 B.n146 585
R478 B.n145 B.n144 585
R479 B.n143 B.n142 585
R480 B.n141 B.n140 585
R481 B.n139 B.n138 585
R482 B.n137 B.n136 585
R483 B.n135 B.n134 585
R484 B.n133 B.n132 585
R485 B.n131 B.n130 585
R486 B.n129 B.n128 585
R487 B.n127 B.n126 585
R488 B.n125 B.n124 585
R489 B.n123 B.n122 585
R490 B.n121 B.n120 585
R491 B.n82 B.n81 585
R492 B.n671 B.n83 585
R493 B.n675 B.n83 585
R494 B.n670 B.n669 585
R495 B.n669 B.n79 585
R496 B.n668 B.n78 585
R497 B.n681 B.n78 585
R498 B.n667 B.n77 585
R499 B.n682 B.n77 585
R500 B.n666 B.n76 585
R501 B.n683 B.n76 585
R502 B.n665 B.n664 585
R503 B.n664 B.n72 585
R504 B.n663 B.n71 585
R505 B.n689 B.n71 585
R506 B.n662 B.n70 585
R507 B.n690 B.n70 585
R508 B.n661 B.n69 585
R509 B.n691 B.n69 585
R510 B.n660 B.n659 585
R511 B.n659 B.n68 585
R512 B.n658 B.n64 585
R513 B.n697 B.n64 585
R514 B.n657 B.n63 585
R515 B.n698 B.n63 585
R516 B.n656 B.n62 585
R517 B.n699 B.n62 585
R518 B.n655 B.n654 585
R519 B.n654 B.n58 585
R520 B.n653 B.n57 585
R521 B.n705 B.n57 585
R522 B.n652 B.n56 585
R523 B.n706 B.n56 585
R524 B.n651 B.n55 585
R525 B.n707 B.n55 585
R526 B.n650 B.n649 585
R527 B.n649 B.n51 585
R528 B.n648 B.n50 585
R529 B.n713 B.n50 585
R530 B.n647 B.n49 585
R531 B.n714 B.n49 585
R532 B.n646 B.n48 585
R533 B.n715 B.n48 585
R534 B.n645 B.n644 585
R535 B.n644 B.n44 585
R536 B.n643 B.n43 585
R537 B.n721 B.n43 585
R538 B.n642 B.n42 585
R539 B.n722 B.n42 585
R540 B.n641 B.n41 585
R541 B.n723 B.n41 585
R542 B.n640 B.n639 585
R543 B.n639 B.n37 585
R544 B.n638 B.n36 585
R545 B.n729 B.n36 585
R546 B.n637 B.n35 585
R547 B.n730 B.n35 585
R548 B.n636 B.n34 585
R549 B.n731 B.n34 585
R550 B.n635 B.n634 585
R551 B.n634 B.n30 585
R552 B.n633 B.n29 585
R553 B.n737 B.n29 585
R554 B.n632 B.n28 585
R555 B.n738 B.n28 585
R556 B.n631 B.n27 585
R557 B.n739 B.n27 585
R558 B.n630 B.n629 585
R559 B.n629 B.n23 585
R560 B.n628 B.n22 585
R561 B.n745 B.n22 585
R562 B.n627 B.n21 585
R563 B.n746 B.n21 585
R564 B.n626 B.n20 585
R565 B.n747 B.n20 585
R566 B.n625 B.n624 585
R567 B.n624 B.n16 585
R568 B.n623 B.n15 585
R569 B.n753 B.n15 585
R570 B.n622 B.n14 585
R571 B.n754 B.n14 585
R572 B.n621 B.n13 585
R573 B.n755 B.n13 585
R574 B.n620 B.n619 585
R575 B.n619 B.n12 585
R576 B.n618 B.n617 585
R577 B.n618 B.n8 585
R578 B.n616 B.n7 585
R579 B.n762 B.n7 585
R580 B.n615 B.n6 585
R581 B.n763 B.n6 585
R582 B.n614 B.n5 585
R583 B.n764 B.n5 585
R584 B.n613 B.n612 585
R585 B.n612 B.n4 585
R586 B.n611 B.n238 585
R587 B.n611 B.n610 585
R588 B.n601 B.n239 585
R589 B.n240 B.n239 585
R590 B.n603 B.n602 585
R591 B.n604 B.n603 585
R592 B.n600 B.n245 585
R593 B.n245 B.n244 585
R594 B.n599 B.n598 585
R595 B.n598 B.n597 585
R596 B.n247 B.n246 585
R597 B.n248 B.n247 585
R598 B.n590 B.n589 585
R599 B.n591 B.n590 585
R600 B.n588 B.n253 585
R601 B.n253 B.n252 585
R602 B.n587 B.n586 585
R603 B.n586 B.n585 585
R604 B.n255 B.n254 585
R605 B.n256 B.n255 585
R606 B.n578 B.n577 585
R607 B.n579 B.n578 585
R608 B.n576 B.n261 585
R609 B.n261 B.n260 585
R610 B.n575 B.n574 585
R611 B.n574 B.n573 585
R612 B.n263 B.n262 585
R613 B.n264 B.n263 585
R614 B.n566 B.n565 585
R615 B.n567 B.n566 585
R616 B.n564 B.n269 585
R617 B.n269 B.n268 585
R618 B.n563 B.n562 585
R619 B.n562 B.n561 585
R620 B.n271 B.n270 585
R621 B.n272 B.n271 585
R622 B.n554 B.n553 585
R623 B.n555 B.n554 585
R624 B.n552 B.n277 585
R625 B.n277 B.n276 585
R626 B.n551 B.n550 585
R627 B.n550 B.n549 585
R628 B.n279 B.n278 585
R629 B.n280 B.n279 585
R630 B.n542 B.n541 585
R631 B.n543 B.n542 585
R632 B.n540 B.n285 585
R633 B.n285 B.n284 585
R634 B.n539 B.n538 585
R635 B.n538 B.n537 585
R636 B.n287 B.n286 585
R637 B.n288 B.n287 585
R638 B.n530 B.n529 585
R639 B.n531 B.n530 585
R640 B.n528 B.n293 585
R641 B.n293 B.n292 585
R642 B.n527 B.n526 585
R643 B.n526 B.n525 585
R644 B.n295 B.n294 585
R645 B.n296 B.n295 585
R646 B.n518 B.n517 585
R647 B.n519 B.n518 585
R648 B.n516 B.n301 585
R649 B.n301 B.n300 585
R650 B.n515 B.n514 585
R651 B.n514 B.n513 585
R652 B.n303 B.n302 585
R653 B.n506 B.n303 585
R654 B.n505 B.n504 585
R655 B.n507 B.n505 585
R656 B.n503 B.n308 585
R657 B.n308 B.n307 585
R658 B.n502 B.n501 585
R659 B.n501 B.n500 585
R660 B.n310 B.n309 585
R661 B.n311 B.n310 585
R662 B.n493 B.n492 585
R663 B.n494 B.n493 585
R664 B.n491 B.n316 585
R665 B.n316 B.n315 585
R666 B.n490 B.n489 585
R667 B.n489 B.n488 585
R668 B.n318 B.n317 585
R669 B.n319 B.n318 585
R670 B.n481 B.n480 585
R671 B.n482 B.n481 585
R672 B.n322 B.n321 585
R673 B.n359 B.n357 585
R674 B.n360 B.n356 585
R675 B.n360 B.n323 585
R676 B.n363 B.n362 585
R677 B.n364 B.n355 585
R678 B.n366 B.n365 585
R679 B.n368 B.n354 585
R680 B.n371 B.n370 585
R681 B.n372 B.n353 585
R682 B.n374 B.n373 585
R683 B.n376 B.n352 585
R684 B.n379 B.n378 585
R685 B.n380 B.n351 585
R686 B.n382 B.n381 585
R687 B.n384 B.n350 585
R688 B.n387 B.n386 585
R689 B.n388 B.n349 585
R690 B.n390 B.n389 585
R691 B.n392 B.n348 585
R692 B.n395 B.n394 585
R693 B.n396 B.n347 585
R694 B.n398 B.n397 585
R695 B.n400 B.n346 585
R696 B.n403 B.n402 585
R697 B.n404 B.n345 585
R698 B.n409 B.n408 585
R699 B.n411 B.n344 585
R700 B.n414 B.n413 585
R701 B.n415 B.n343 585
R702 B.n417 B.n416 585
R703 B.n419 B.n342 585
R704 B.n422 B.n421 585
R705 B.n423 B.n341 585
R706 B.n425 B.n424 585
R707 B.n427 B.n340 585
R708 B.n430 B.n429 585
R709 B.n431 B.n336 585
R710 B.n433 B.n432 585
R711 B.n435 B.n335 585
R712 B.n438 B.n437 585
R713 B.n439 B.n334 585
R714 B.n441 B.n440 585
R715 B.n443 B.n333 585
R716 B.n446 B.n445 585
R717 B.n447 B.n332 585
R718 B.n449 B.n448 585
R719 B.n451 B.n331 585
R720 B.n454 B.n453 585
R721 B.n455 B.n330 585
R722 B.n457 B.n456 585
R723 B.n459 B.n329 585
R724 B.n462 B.n461 585
R725 B.n463 B.n328 585
R726 B.n465 B.n464 585
R727 B.n467 B.n327 585
R728 B.n470 B.n469 585
R729 B.n471 B.n326 585
R730 B.n473 B.n472 585
R731 B.n475 B.n325 585
R732 B.n478 B.n477 585
R733 B.n479 B.n324 585
R734 B.n484 B.n483 585
R735 B.n483 B.n482 585
R736 B.n485 B.n320 585
R737 B.n320 B.n319 585
R738 B.n487 B.n486 585
R739 B.n488 B.n487 585
R740 B.n314 B.n313 585
R741 B.n315 B.n314 585
R742 B.n496 B.n495 585
R743 B.n495 B.n494 585
R744 B.n497 B.n312 585
R745 B.n312 B.n311 585
R746 B.n499 B.n498 585
R747 B.n500 B.n499 585
R748 B.n306 B.n305 585
R749 B.n307 B.n306 585
R750 B.n509 B.n508 585
R751 B.n508 B.n507 585
R752 B.n510 B.n304 585
R753 B.n506 B.n304 585
R754 B.n512 B.n511 585
R755 B.n513 B.n512 585
R756 B.n299 B.n298 585
R757 B.n300 B.n299 585
R758 B.n521 B.n520 585
R759 B.n520 B.n519 585
R760 B.n522 B.n297 585
R761 B.n297 B.n296 585
R762 B.n524 B.n523 585
R763 B.n525 B.n524 585
R764 B.n291 B.n290 585
R765 B.n292 B.n291 585
R766 B.n533 B.n532 585
R767 B.n532 B.n531 585
R768 B.n534 B.n289 585
R769 B.n289 B.n288 585
R770 B.n536 B.n535 585
R771 B.n537 B.n536 585
R772 B.n283 B.n282 585
R773 B.n284 B.n283 585
R774 B.n545 B.n544 585
R775 B.n544 B.n543 585
R776 B.n546 B.n281 585
R777 B.n281 B.n280 585
R778 B.n548 B.n547 585
R779 B.n549 B.n548 585
R780 B.n275 B.n274 585
R781 B.n276 B.n275 585
R782 B.n557 B.n556 585
R783 B.n556 B.n555 585
R784 B.n558 B.n273 585
R785 B.n273 B.n272 585
R786 B.n560 B.n559 585
R787 B.n561 B.n560 585
R788 B.n267 B.n266 585
R789 B.n268 B.n267 585
R790 B.n569 B.n568 585
R791 B.n568 B.n567 585
R792 B.n570 B.n265 585
R793 B.n265 B.n264 585
R794 B.n572 B.n571 585
R795 B.n573 B.n572 585
R796 B.n259 B.n258 585
R797 B.n260 B.n259 585
R798 B.n581 B.n580 585
R799 B.n580 B.n579 585
R800 B.n582 B.n257 585
R801 B.n257 B.n256 585
R802 B.n584 B.n583 585
R803 B.n585 B.n584 585
R804 B.n251 B.n250 585
R805 B.n252 B.n251 585
R806 B.n593 B.n592 585
R807 B.n592 B.n591 585
R808 B.n594 B.n249 585
R809 B.n249 B.n248 585
R810 B.n596 B.n595 585
R811 B.n597 B.n596 585
R812 B.n243 B.n242 585
R813 B.n244 B.n243 585
R814 B.n606 B.n605 585
R815 B.n605 B.n604 585
R816 B.n607 B.n241 585
R817 B.n241 B.n240 585
R818 B.n609 B.n608 585
R819 B.n610 B.n609 585
R820 B.n3 B.n0 585
R821 B.n4 B.n3 585
R822 B.n761 B.n1 585
R823 B.n762 B.n761 585
R824 B.n760 B.n759 585
R825 B.n760 B.n8 585
R826 B.n758 B.n9 585
R827 B.n12 B.n9 585
R828 B.n757 B.n756 585
R829 B.n756 B.n755 585
R830 B.n11 B.n10 585
R831 B.n754 B.n11 585
R832 B.n752 B.n751 585
R833 B.n753 B.n752 585
R834 B.n750 B.n17 585
R835 B.n17 B.n16 585
R836 B.n749 B.n748 585
R837 B.n748 B.n747 585
R838 B.n19 B.n18 585
R839 B.n746 B.n19 585
R840 B.n744 B.n743 585
R841 B.n745 B.n744 585
R842 B.n742 B.n24 585
R843 B.n24 B.n23 585
R844 B.n741 B.n740 585
R845 B.n740 B.n739 585
R846 B.n26 B.n25 585
R847 B.n738 B.n26 585
R848 B.n736 B.n735 585
R849 B.n737 B.n736 585
R850 B.n734 B.n31 585
R851 B.n31 B.n30 585
R852 B.n733 B.n732 585
R853 B.n732 B.n731 585
R854 B.n33 B.n32 585
R855 B.n730 B.n33 585
R856 B.n728 B.n727 585
R857 B.n729 B.n728 585
R858 B.n726 B.n38 585
R859 B.n38 B.n37 585
R860 B.n725 B.n724 585
R861 B.n724 B.n723 585
R862 B.n40 B.n39 585
R863 B.n722 B.n40 585
R864 B.n720 B.n719 585
R865 B.n721 B.n720 585
R866 B.n718 B.n45 585
R867 B.n45 B.n44 585
R868 B.n717 B.n716 585
R869 B.n716 B.n715 585
R870 B.n47 B.n46 585
R871 B.n714 B.n47 585
R872 B.n712 B.n711 585
R873 B.n713 B.n712 585
R874 B.n710 B.n52 585
R875 B.n52 B.n51 585
R876 B.n709 B.n708 585
R877 B.n708 B.n707 585
R878 B.n54 B.n53 585
R879 B.n706 B.n54 585
R880 B.n704 B.n703 585
R881 B.n705 B.n704 585
R882 B.n702 B.n59 585
R883 B.n59 B.n58 585
R884 B.n701 B.n700 585
R885 B.n700 B.n699 585
R886 B.n61 B.n60 585
R887 B.n698 B.n61 585
R888 B.n696 B.n695 585
R889 B.n697 B.n696 585
R890 B.n694 B.n65 585
R891 B.n68 B.n65 585
R892 B.n693 B.n692 585
R893 B.n692 B.n691 585
R894 B.n67 B.n66 585
R895 B.n690 B.n67 585
R896 B.n688 B.n687 585
R897 B.n689 B.n688 585
R898 B.n686 B.n73 585
R899 B.n73 B.n72 585
R900 B.n685 B.n684 585
R901 B.n684 B.n683 585
R902 B.n75 B.n74 585
R903 B.n682 B.n75 585
R904 B.n680 B.n679 585
R905 B.n681 B.n680 585
R906 B.n678 B.n80 585
R907 B.n80 B.n79 585
R908 B.n677 B.n676 585
R909 B.n676 B.n675 585
R910 B.n765 B.n764 585
R911 B.n763 B.n2 585
R912 B.n676 B.n82 463.671
R913 B.n673 B.n83 463.671
R914 B.n481 B.n324 463.671
R915 B.n483 B.n322 463.671
R916 B.n115 B.t6 268.435
R917 B.n337 B.t17 268.435
R918 B.n117 B.t9 268.435
R919 B.n405 B.t14 268.435
R920 B.n674 B.n113 256.663
R921 B.n674 B.n112 256.663
R922 B.n674 B.n111 256.663
R923 B.n674 B.n110 256.663
R924 B.n674 B.n109 256.663
R925 B.n674 B.n108 256.663
R926 B.n674 B.n107 256.663
R927 B.n674 B.n106 256.663
R928 B.n674 B.n105 256.663
R929 B.n674 B.n104 256.663
R930 B.n674 B.n103 256.663
R931 B.n674 B.n102 256.663
R932 B.n674 B.n101 256.663
R933 B.n674 B.n100 256.663
R934 B.n674 B.n99 256.663
R935 B.n674 B.n98 256.663
R936 B.n674 B.n97 256.663
R937 B.n674 B.n96 256.663
R938 B.n674 B.n95 256.663
R939 B.n674 B.n94 256.663
R940 B.n674 B.n93 256.663
R941 B.n674 B.n92 256.663
R942 B.n674 B.n91 256.663
R943 B.n674 B.n90 256.663
R944 B.n674 B.n89 256.663
R945 B.n674 B.n88 256.663
R946 B.n674 B.n87 256.663
R947 B.n674 B.n86 256.663
R948 B.n674 B.n85 256.663
R949 B.n674 B.n84 256.663
R950 B.n358 B.n323 256.663
R951 B.n361 B.n323 256.663
R952 B.n367 B.n323 256.663
R953 B.n369 B.n323 256.663
R954 B.n375 B.n323 256.663
R955 B.n377 B.n323 256.663
R956 B.n383 B.n323 256.663
R957 B.n385 B.n323 256.663
R958 B.n391 B.n323 256.663
R959 B.n393 B.n323 256.663
R960 B.n399 B.n323 256.663
R961 B.n401 B.n323 256.663
R962 B.n410 B.n323 256.663
R963 B.n412 B.n323 256.663
R964 B.n418 B.n323 256.663
R965 B.n420 B.n323 256.663
R966 B.n426 B.n323 256.663
R967 B.n428 B.n323 256.663
R968 B.n434 B.n323 256.663
R969 B.n436 B.n323 256.663
R970 B.n442 B.n323 256.663
R971 B.n444 B.n323 256.663
R972 B.n450 B.n323 256.663
R973 B.n452 B.n323 256.663
R974 B.n458 B.n323 256.663
R975 B.n460 B.n323 256.663
R976 B.n466 B.n323 256.663
R977 B.n468 B.n323 256.663
R978 B.n474 B.n323 256.663
R979 B.n476 B.n323 256.663
R980 B.n767 B.n766 256.663
R981 B.n117 B.t8 251.447
R982 B.n115 B.t4 251.447
R983 B.n337 B.t15 251.447
R984 B.n405 B.t11 251.447
R985 B.n116 B.t7 188.919
R986 B.n338 B.t16 188.919
R987 B.n118 B.t10 188.919
R988 B.n406 B.t13 188.919
R989 B.n122 B.n121 163.367
R990 B.n126 B.n125 163.367
R991 B.n130 B.n129 163.367
R992 B.n134 B.n133 163.367
R993 B.n138 B.n137 163.367
R994 B.n142 B.n141 163.367
R995 B.n146 B.n145 163.367
R996 B.n150 B.n149 163.367
R997 B.n154 B.n153 163.367
R998 B.n158 B.n157 163.367
R999 B.n162 B.n161 163.367
R1000 B.n166 B.n165 163.367
R1001 B.n170 B.n169 163.367
R1002 B.n174 B.n173 163.367
R1003 B.n178 B.n177 163.367
R1004 B.n182 B.n181 163.367
R1005 B.n186 B.n185 163.367
R1006 B.n191 B.n190 163.367
R1007 B.n195 B.n194 163.367
R1008 B.n199 B.n198 163.367
R1009 B.n203 B.n202 163.367
R1010 B.n207 B.n206 163.367
R1011 B.n211 B.n210 163.367
R1012 B.n215 B.n214 163.367
R1013 B.n219 B.n218 163.367
R1014 B.n223 B.n222 163.367
R1015 B.n227 B.n226 163.367
R1016 B.n231 B.n230 163.367
R1017 B.n235 B.n234 163.367
R1018 B.n673 B.n114 163.367
R1019 B.n481 B.n318 163.367
R1020 B.n489 B.n318 163.367
R1021 B.n489 B.n316 163.367
R1022 B.n493 B.n316 163.367
R1023 B.n493 B.n310 163.367
R1024 B.n501 B.n310 163.367
R1025 B.n501 B.n308 163.367
R1026 B.n505 B.n308 163.367
R1027 B.n505 B.n303 163.367
R1028 B.n514 B.n303 163.367
R1029 B.n514 B.n301 163.367
R1030 B.n518 B.n301 163.367
R1031 B.n518 B.n295 163.367
R1032 B.n526 B.n295 163.367
R1033 B.n526 B.n293 163.367
R1034 B.n530 B.n293 163.367
R1035 B.n530 B.n287 163.367
R1036 B.n538 B.n287 163.367
R1037 B.n538 B.n285 163.367
R1038 B.n542 B.n285 163.367
R1039 B.n542 B.n279 163.367
R1040 B.n550 B.n279 163.367
R1041 B.n550 B.n277 163.367
R1042 B.n554 B.n277 163.367
R1043 B.n554 B.n271 163.367
R1044 B.n562 B.n271 163.367
R1045 B.n562 B.n269 163.367
R1046 B.n566 B.n269 163.367
R1047 B.n566 B.n263 163.367
R1048 B.n574 B.n263 163.367
R1049 B.n574 B.n261 163.367
R1050 B.n578 B.n261 163.367
R1051 B.n578 B.n255 163.367
R1052 B.n586 B.n255 163.367
R1053 B.n586 B.n253 163.367
R1054 B.n590 B.n253 163.367
R1055 B.n590 B.n247 163.367
R1056 B.n598 B.n247 163.367
R1057 B.n598 B.n245 163.367
R1058 B.n603 B.n245 163.367
R1059 B.n603 B.n239 163.367
R1060 B.n611 B.n239 163.367
R1061 B.n612 B.n611 163.367
R1062 B.n612 B.n5 163.367
R1063 B.n6 B.n5 163.367
R1064 B.n7 B.n6 163.367
R1065 B.n618 B.n7 163.367
R1066 B.n619 B.n618 163.367
R1067 B.n619 B.n13 163.367
R1068 B.n14 B.n13 163.367
R1069 B.n15 B.n14 163.367
R1070 B.n624 B.n15 163.367
R1071 B.n624 B.n20 163.367
R1072 B.n21 B.n20 163.367
R1073 B.n22 B.n21 163.367
R1074 B.n629 B.n22 163.367
R1075 B.n629 B.n27 163.367
R1076 B.n28 B.n27 163.367
R1077 B.n29 B.n28 163.367
R1078 B.n634 B.n29 163.367
R1079 B.n634 B.n34 163.367
R1080 B.n35 B.n34 163.367
R1081 B.n36 B.n35 163.367
R1082 B.n639 B.n36 163.367
R1083 B.n639 B.n41 163.367
R1084 B.n42 B.n41 163.367
R1085 B.n43 B.n42 163.367
R1086 B.n644 B.n43 163.367
R1087 B.n644 B.n48 163.367
R1088 B.n49 B.n48 163.367
R1089 B.n50 B.n49 163.367
R1090 B.n649 B.n50 163.367
R1091 B.n649 B.n55 163.367
R1092 B.n56 B.n55 163.367
R1093 B.n57 B.n56 163.367
R1094 B.n654 B.n57 163.367
R1095 B.n654 B.n62 163.367
R1096 B.n63 B.n62 163.367
R1097 B.n64 B.n63 163.367
R1098 B.n659 B.n64 163.367
R1099 B.n659 B.n69 163.367
R1100 B.n70 B.n69 163.367
R1101 B.n71 B.n70 163.367
R1102 B.n664 B.n71 163.367
R1103 B.n664 B.n76 163.367
R1104 B.n77 B.n76 163.367
R1105 B.n78 B.n77 163.367
R1106 B.n669 B.n78 163.367
R1107 B.n669 B.n83 163.367
R1108 B.n360 B.n359 163.367
R1109 B.n362 B.n360 163.367
R1110 B.n366 B.n355 163.367
R1111 B.n370 B.n368 163.367
R1112 B.n374 B.n353 163.367
R1113 B.n378 B.n376 163.367
R1114 B.n382 B.n351 163.367
R1115 B.n386 B.n384 163.367
R1116 B.n390 B.n349 163.367
R1117 B.n394 B.n392 163.367
R1118 B.n398 B.n347 163.367
R1119 B.n402 B.n400 163.367
R1120 B.n409 B.n345 163.367
R1121 B.n413 B.n411 163.367
R1122 B.n417 B.n343 163.367
R1123 B.n421 B.n419 163.367
R1124 B.n425 B.n341 163.367
R1125 B.n429 B.n427 163.367
R1126 B.n433 B.n336 163.367
R1127 B.n437 B.n435 163.367
R1128 B.n441 B.n334 163.367
R1129 B.n445 B.n443 163.367
R1130 B.n449 B.n332 163.367
R1131 B.n453 B.n451 163.367
R1132 B.n457 B.n330 163.367
R1133 B.n461 B.n459 163.367
R1134 B.n465 B.n328 163.367
R1135 B.n469 B.n467 163.367
R1136 B.n473 B.n326 163.367
R1137 B.n477 B.n475 163.367
R1138 B.n483 B.n320 163.367
R1139 B.n487 B.n320 163.367
R1140 B.n487 B.n314 163.367
R1141 B.n495 B.n314 163.367
R1142 B.n495 B.n312 163.367
R1143 B.n499 B.n312 163.367
R1144 B.n499 B.n306 163.367
R1145 B.n508 B.n306 163.367
R1146 B.n508 B.n304 163.367
R1147 B.n512 B.n304 163.367
R1148 B.n512 B.n299 163.367
R1149 B.n520 B.n299 163.367
R1150 B.n520 B.n297 163.367
R1151 B.n524 B.n297 163.367
R1152 B.n524 B.n291 163.367
R1153 B.n532 B.n291 163.367
R1154 B.n532 B.n289 163.367
R1155 B.n536 B.n289 163.367
R1156 B.n536 B.n283 163.367
R1157 B.n544 B.n283 163.367
R1158 B.n544 B.n281 163.367
R1159 B.n548 B.n281 163.367
R1160 B.n548 B.n275 163.367
R1161 B.n556 B.n275 163.367
R1162 B.n556 B.n273 163.367
R1163 B.n560 B.n273 163.367
R1164 B.n560 B.n267 163.367
R1165 B.n568 B.n267 163.367
R1166 B.n568 B.n265 163.367
R1167 B.n572 B.n265 163.367
R1168 B.n572 B.n259 163.367
R1169 B.n580 B.n259 163.367
R1170 B.n580 B.n257 163.367
R1171 B.n584 B.n257 163.367
R1172 B.n584 B.n251 163.367
R1173 B.n592 B.n251 163.367
R1174 B.n592 B.n249 163.367
R1175 B.n596 B.n249 163.367
R1176 B.n596 B.n243 163.367
R1177 B.n605 B.n243 163.367
R1178 B.n605 B.n241 163.367
R1179 B.n609 B.n241 163.367
R1180 B.n609 B.n3 163.367
R1181 B.n765 B.n3 163.367
R1182 B.n761 B.n2 163.367
R1183 B.n761 B.n760 163.367
R1184 B.n760 B.n9 163.367
R1185 B.n756 B.n9 163.367
R1186 B.n756 B.n11 163.367
R1187 B.n752 B.n11 163.367
R1188 B.n752 B.n17 163.367
R1189 B.n748 B.n17 163.367
R1190 B.n748 B.n19 163.367
R1191 B.n744 B.n19 163.367
R1192 B.n744 B.n24 163.367
R1193 B.n740 B.n24 163.367
R1194 B.n740 B.n26 163.367
R1195 B.n736 B.n26 163.367
R1196 B.n736 B.n31 163.367
R1197 B.n732 B.n31 163.367
R1198 B.n732 B.n33 163.367
R1199 B.n728 B.n33 163.367
R1200 B.n728 B.n38 163.367
R1201 B.n724 B.n38 163.367
R1202 B.n724 B.n40 163.367
R1203 B.n720 B.n40 163.367
R1204 B.n720 B.n45 163.367
R1205 B.n716 B.n45 163.367
R1206 B.n716 B.n47 163.367
R1207 B.n712 B.n47 163.367
R1208 B.n712 B.n52 163.367
R1209 B.n708 B.n52 163.367
R1210 B.n708 B.n54 163.367
R1211 B.n704 B.n54 163.367
R1212 B.n704 B.n59 163.367
R1213 B.n700 B.n59 163.367
R1214 B.n700 B.n61 163.367
R1215 B.n696 B.n61 163.367
R1216 B.n696 B.n65 163.367
R1217 B.n692 B.n65 163.367
R1218 B.n692 B.n67 163.367
R1219 B.n688 B.n67 163.367
R1220 B.n688 B.n73 163.367
R1221 B.n684 B.n73 163.367
R1222 B.n684 B.n75 163.367
R1223 B.n680 B.n75 163.367
R1224 B.n680 B.n80 163.367
R1225 B.n676 B.n80 163.367
R1226 B.n482 B.n323 101.055
R1227 B.n675 B.n674 101.055
R1228 B.n118 B.n117 79.5157
R1229 B.n116 B.n115 79.5157
R1230 B.n338 B.n337 79.5157
R1231 B.n406 B.n405 79.5157
R1232 B.n84 B.n82 71.676
R1233 B.n122 B.n85 71.676
R1234 B.n126 B.n86 71.676
R1235 B.n130 B.n87 71.676
R1236 B.n134 B.n88 71.676
R1237 B.n138 B.n89 71.676
R1238 B.n142 B.n90 71.676
R1239 B.n146 B.n91 71.676
R1240 B.n150 B.n92 71.676
R1241 B.n154 B.n93 71.676
R1242 B.n158 B.n94 71.676
R1243 B.n162 B.n95 71.676
R1244 B.n166 B.n96 71.676
R1245 B.n170 B.n97 71.676
R1246 B.n174 B.n98 71.676
R1247 B.n178 B.n99 71.676
R1248 B.n182 B.n100 71.676
R1249 B.n186 B.n101 71.676
R1250 B.n191 B.n102 71.676
R1251 B.n195 B.n103 71.676
R1252 B.n199 B.n104 71.676
R1253 B.n203 B.n105 71.676
R1254 B.n207 B.n106 71.676
R1255 B.n211 B.n107 71.676
R1256 B.n215 B.n108 71.676
R1257 B.n219 B.n109 71.676
R1258 B.n223 B.n110 71.676
R1259 B.n227 B.n111 71.676
R1260 B.n231 B.n112 71.676
R1261 B.n235 B.n113 71.676
R1262 B.n114 B.n113 71.676
R1263 B.n234 B.n112 71.676
R1264 B.n230 B.n111 71.676
R1265 B.n226 B.n110 71.676
R1266 B.n222 B.n109 71.676
R1267 B.n218 B.n108 71.676
R1268 B.n214 B.n107 71.676
R1269 B.n210 B.n106 71.676
R1270 B.n206 B.n105 71.676
R1271 B.n202 B.n104 71.676
R1272 B.n198 B.n103 71.676
R1273 B.n194 B.n102 71.676
R1274 B.n190 B.n101 71.676
R1275 B.n185 B.n100 71.676
R1276 B.n181 B.n99 71.676
R1277 B.n177 B.n98 71.676
R1278 B.n173 B.n97 71.676
R1279 B.n169 B.n96 71.676
R1280 B.n165 B.n95 71.676
R1281 B.n161 B.n94 71.676
R1282 B.n157 B.n93 71.676
R1283 B.n153 B.n92 71.676
R1284 B.n149 B.n91 71.676
R1285 B.n145 B.n90 71.676
R1286 B.n141 B.n89 71.676
R1287 B.n137 B.n88 71.676
R1288 B.n133 B.n87 71.676
R1289 B.n129 B.n86 71.676
R1290 B.n125 B.n85 71.676
R1291 B.n121 B.n84 71.676
R1292 B.n358 B.n322 71.676
R1293 B.n362 B.n361 71.676
R1294 B.n367 B.n366 71.676
R1295 B.n370 B.n369 71.676
R1296 B.n375 B.n374 71.676
R1297 B.n378 B.n377 71.676
R1298 B.n383 B.n382 71.676
R1299 B.n386 B.n385 71.676
R1300 B.n391 B.n390 71.676
R1301 B.n394 B.n393 71.676
R1302 B.n399 B.n398 71.676
R1303 B.n402 B.n401 71.676
R1304 B.n410 B.n409 71.676
R1305 B.n413 B.n412 71.676
R1306 B.n418 B.n417 71.676
R1307 B.n421 B.n420 71.676
R1308 B.n426 B.n425 71.676
R1309 B.n429 B.n428 71.676
R1310 B.n434 B.n433 71.676
R1311 B.n437 B.n436 71.676
R1312 B.n442 B.n441 71.676
R1313 B.n445 B.n444 71.676
R1314 B.n450 B.n449 71.676
R1315 B.n453 B.n452 71.676
R1316 B.n458 B.n457 71.676
R1317 B.n461 B.n460 71.676
R1318 B.n466 B.n465 71.676
R1319 B.n469 B.n468 71.676
R1320 B.n474 B.n473 71.676
R1321 B.n477 B.n476 71.676
R1322 B.n359 B.n358 71.676
R1323 B.n361 B.n355 71.676
R1324 B.n368 B.n367 71.676
R1325 B.n369 B.n353 71.676
R1326 B.n376 B.n375 71.676
R1327 B.n377 B.n351 71.676
R1328 B.n384 B.n383 71.676
R1329 B.n385 B.n349 71.676
R1330 B.n392 B.n391 71.676
R1331 B.n393 B.n347 71.676
R1332 B.n400 B.n399 71.676
R1333 B.n401 B.n345 71.676
R1334 B.n411 B.n410 71.676
R1335 B.n412 B.n343 71.676
R1336 B.n419 B.n418 71.676
R1337 B.n420 B.n341 71.676
R1338 B.n427 B.n426 71.676
R1339 B.n428 B.n336 71.676
R1340 B.n435 B.n434 71.676
R1341 B.n436 B.n334 71.676
R1342 B.n443 B.n442 71.676
R1343 B.n444 B.n332 71.676
R1344 B.n451 B.n450 71.676
R1345 B.n452 B.n330 71.676
R1346 B.n459 B.n458 71.676
R1347 B.n460 B.n328 71.676
R1348 B.n467 B.n466 71.676
R1349 B.n468 B.n326 71.676
R1350 B.n475 B.n474 71.676
R1351 B.n476 B.n324 71.676
R1352 B.n766 B.n765 71.676
R1353 B.n766 B.n2 71.676
R1354 B.n482 B.n319 63.0431
R1355 B.n488 B.n319 63.0431
R1356 B.n488 B.n315 63.0431
R1357 B.n494 B.n315 63.0431
R1358 B.n494 B.n311 63.0431
R1359 B.n500 B.n311 63.0431
R1360 B.n500 B.n307 63.0431
R1361 B.n507 B.n307 63.0431
R1362 B.n507 B.n506 63.0431
R1363 B.n513 B.n300 63.0431
R1364 B.n519 B.n300 63.0431
R1365 B.n519 B.n296 63.0431
R1366 B.n525 B.n296 63.0431
R1367 B.n525 B.n292 63.0431
R1368 B.n531 B.n292 63.0431
R1369 B.n531 B.n288 63.0431
R1370 B.n537 B.n288 63.0431
R1371 B.n537 B.n284 63.0431
R1372 B.n543 B.n284 63.0431
R1373 B.n543 B.n280 63.0431
R1374 B.n549 B.n280 63.0431
R1375 B.n549 B.n276 63.0431
R1376 B.n555 B.n276 63.0431
R1377 B.n561 B.n272 63.0431
R1378 B.n561 B.n268 63.0431
R1379 B.n567 B.n268 63.0431
R1380 B.n567 B.n264 63.0431
R1381 B.n573 B.n264 63.0431
R1382 B.n573 B.n260 63.0431
R1383 B.n579 B.n260 63.0431
R1384 B.n579 B.n256 63.0431
R1385 B.n585 B.n256 63.0431
R1386 B.n585 B.n252 63.0431
R1387 B.n591 B.n252 63.0431
R1388 B.n597 B.n248 63.0431
R1389 B.n597 B.n244 63.0431
R1390 B.n604 B.n244 63.0431
R1391 B.n604 B.n240 63.0431
R1392 B.n610 B.n240 63.0431
R1393 B.n610 B.n4 63.0431
R1394 B.n764 B.n4 63.0431
R1395 B.n764 B.n763 63.0431
R1396 B.n763 B.n762 63.0431
R1397 B.n762 B.n8 63.0431
R1398 B.n12 B.n8 63.0431
R1399 B.n755 B.n12 63.0431
R1400 B.n755 B.n754 63.0431
R1401 B.n754 B.n753 63.0431
R1402 B.n753 B.n16 63.0431
R1403 B.n747 B.n746 63.0431
R1404 B.n746 B.n745 63.0431
R1405 B.n745 B.n23 63.0431
R1406 B.n739 B.n23 63.0431
R1407 B.n739 B.n738 63.0431
R1408 B.n738 B.n737 63.0431
R1409 B.n737 B.n30 63.0431
R1410 B.n731 B.n30 63.0431
R1411 B.n731 B.n730 63.0431
R1412 B.n730 B.n729 63.0431
R1413 B.n729 B.n37 63.0431
R1414 B.n723 B.n722 63.0431
R1415 B.n722 B.n721 63.0431
R1416 B.n721 B.n44 63.0431
R1417 B.n715 B.n44 63.0431
R1418 B.n715 B.n714 63.0431
R1419 B.n714 B.n713 63.0431
R1420 B.n713 B.n51 63.0431
R1421 B.n707 B.n51 63.0431
R1422 B.n707 B.n706 63.0431
R1423 B.n706 B.n705 63.0431
R1424 B.n705 B.n58 63.0431
R1425 B.n699 B.n58 63.0431
R1426 B.n699 B.n698 63.0431
R1427 B.n698 B.n697 63.0431
R1428 B.n691 B.n68 63.0431
R1429 B.n691 B.n690 63.0431
R1430 B.n690 B.n689 63.0431
R1431 B.n689 B.n72 63.0431
R1432 B.n683 B.n72 63.0431
R1433 B.n683 B.n682 63.0431
R1434 B.n682 B.n681 63.0431
R1435 B.n681 B.n79 63.0431
R1436 B.n675 B.n79 63.0431
R1437 B.n119 B.n118 59.5399
R1438 B.n188 B.n116 59.5399
R1439 B.n339 B.n338 59.5399
R1440 B.n407 B.n406 59.5399
R1441 B.n591 B.t3 54.6992
R1442 B.n747 B.t1 54.6992
R1443 B.n555 B.t2 50.9908
R1444 B.n723 B.t0 50.9908
R1445 B.n506 B.t12 34.3031
R1446 B.n68 B.t5 34.3031
R1447 B.n484 B.n321 30.1273
R1448 B.n480 B.n479 30.1273
R1449 B.n677 B.n81 30.1273
R1450 B.n672 B.n671 30.1273
R1451 B.n513 B.t12 28.7405
R1452 B.n697 B.t5 28.7405
R1453 B B.n767 18.0485
R1454 B.t2 B.n272 12.0528
R1455 B.t0 B.n37 12.0528
R1456 B.n485 B.n484 10.6151
R1457 B.n486 B.n485 10.6151
R1458 B.n486 B.n313 10.6151
R1459 B.n496 B.n313 10.6151
R1460 B.n497 B.n496 10.6151
R1461 B.n498 B.n497 10.6151
R1462 B.n498 B.n305 10.6151
R1463 B.n509 B.n305 10.6151
R1464 B.n510 B.n509 10.6151
R1465 B.n511 B.n510 10.6151
R1466 B.n511 B.n298 10.6151
R1467 B.n521 B.n298 10.6151
R1468 B.n522 B.n521 10.6151
R1469 B.n523 B.n522 10.6151
R1470 B.n523 B.n290 10.6151
R1471 B.n533 B.n290 10.6151
R1472 B.n534 B.n533 10.6151
R1473 B.n535 B.n534 10.6151
R1474 B.n535 B.n282 10.6151
R1475 B.n545 B.n282 10.6151
R1476 B.n546 B.n545 10.6151
R1477 B.n547 B.n546 10.6151
R1478 B.n547 B.n274 10.6151
R1479 B.n557 B.n274 10.6151
R1480 B.n558 B.n557 10.6151
R1481 B.n559 B.n558 10.6151
R1482 B.n559 B.n266 10.6151
R1483 B.n569 B.n266 10.6151
R1484 B.n570 B.n569 10.6151
R1485 B.n571 B.n570 10.6151
R1486 B.n571 B.n258 10.6151
R1487 B.n581 B.n258 10.6151
R1488 B.n582 B.n581 10.6151
R1489 B.n583 B.n582 10.6151
R1490 B.n583 B.n250 10.6151
R1491 B.n593 B.n250 10.6151
R1492 B.n594 B.n593 10.6151
R1493 B.n595 B.n594 10.6151
R1494 B.n595 B.n242 10.6151
R1495 B.n606 B.n242 10.6151
R1496 B.n607 B.n606 10.6151
R1497 B.n608 B.n607 10.6151
R1498 B.n608 B.n0 10.6151
R1499 B.n357 B.n321 10.6151
R1500 B.n357 B.n356 10.6151
R1501 B.n363 B.n356 10.6151
R1502 B.n364 B.n363 10.6151
R1503 B.n365 B.n364 10.6151
R1504 B.n365 B.n354 10.6151
R1505 B.n371 B.n354 10.6151
R1506 B.n372 B.n371 10.6151
R1507 B.n373 B.n372 10.6151
R1508 B.n373 B.n352 10.6151
R1509 B.n379 B.n352 10.6151
R1510 B.n380 B.n379 10.6151
R1511 B.n381 B.n380 10.6151
R1512 B.n381 B.n350 10.6151
R1513 B.n387 B.n350 10.6151
R1514 B.n388 B.n387 10.6151
R1515 B.n389 B.n388 10.6151
R1516 B.n389 B.n348 10.6151
R1517 B.n395 B.n348 10.6151
R1518 B.n396 B.n395 10.6151
R1519 B.n397 B.n396 10.6151
R1520 B.n397 B.n346 10.6151
R1521 B.n403 B.n346 10.6151
R1522 B.n404 B.n403 10.6151
R1523 B.n408 B.n404 10.6151
R1524 B.n414 B.n344 10.6151
R1525 B.n415 B.n414 10.6151
R1526 B.n416 B.n415 10.6151
R1527 B.n416 B.n342 10.6151
R1528 B.n422 B.n342 10.6151
R1529 B.n423 B.n422 10.6151
R1530 B.n424 B.n423 10.6151
R1531 B.n424 B.n340 10.6151
R1532 B.n431 B.n430 10.6151
R1533 B.n432 B.n431 10.6151
R1534 B.n432 B.n335 10.6151
R1535 B.n438 B.n335 10.6151
R1536 B.n439 B.n438 10.6151
R1537 B.n440 B.n439 10.6151
R1538 B.n440 B.n333 10.6151
R1539 B.n446 B.n333 10.6151
R1540 B.n447 B.n446 10.6151
R1541 B.n448 B.n447 10.6151
R1542 B.n448 B.n331 10.6151
R1543 B.n454 B.n331 10.6151
R1544 B.n455 B.n454 10.6151
R1545 B.n456 B.n455 10.6151
R1546 B.n456 B.n329 10.6151
R1547 B.n462 B.n329 10.6151
R1548 B.n463 B.n462 10.6151
R1549 B.n464 B.n463 10.6151
R1550 B.n464 B.n327 10.6151
R1551 B.n470 B.n327 10.6151
R1552 B.n471 B.n470 10.6151
R1553 B.n472 B.n471 10.6151
R1554 B.n472 B.n325 10.6151
R1555 B.n478 B.n325 10.6151
R1556 B.n479 B.n478 10.6151
R1557 B.n480 B.n317 10.6151
R1558 B.n490 B.n317 10.6151
R1559 B.n491 B.n490 10.6151
R1560 B.n492 B.n491 10.6151
R1561 B.n492 B.n309 10.6151
R1562 B.n502 B.n309 10.6151
R1563 B.n503 B.n502 10.6151
R1564 B.n504 B.n503 10.6151
R1565 B.n504 B.n302 10.6151
R1566 B.n515 B.n302 10.6151
R1567 B.n516 B.n515 10.6151
R1568 B.n517 B.n516 10.6151
R1569 B.n517 B.n294 10.6151
R1570 B.n527 B.n294 10.6151
R1571 B.n528 B.n527 10.6151
R1572 B.n529 B.n528 10.6151
R1573 B.n529 B.n286 10.6151
R1574 B.n539 B.n286 10.6151
R1575 B.n540 B.n539 10.6151
R1576 B.n541 B.n540 10.6151
R1577 B.n541 B.n278 10.6151
R1578 B.n551 B.n278 10.6151
R1579 B.n552 B.n551 10.6151
R1580 B.n553 B.n552 10.6151
R1581 B.n553 B.n270 10.6151
R1582 B.n563 B.n270 10.6151
R1583 B.n564 B.n563 10.6151
R1584 B.n565 B.n564 10.6151
R1585 B.n565 B.n262 10.6151
R1586 B.n575 B.n262 10.6151
R1587 B.n576 B.n575 10.6151
R1588 B.n577 B.n576 10.6151
R1589 B.n577 B.n254 10.6151
R1590 B.n587 B.n254 10.6151
R1591 B.n588 B.n587 10.6151
R1592 B.n589 B.n588 10.6151
R1593 B.n589 B.n246 10.6151
R1594 B.n599 B.n246 10.6151
R1595 B.n600 B.n599 10.6151
R1596 B.n602 B.n600 10.6151
R1597 B.n602 B.n601 10.6151
R1598 B.n601 B.n238 10.6151
R1599 B.n613 B.n238 10.6151
R1600 B.n614 B.n613 10.6151
R1601 B.n615 B.n614 10.6151
R1602 B.n616 B.n615 10.6151
R1603 B.n617 B.n616 10.6151
R1604 B.n620 B.n617 10.6151
R1605 B.n621 B.n620 10.6151
R1606 B.n622 B.n621 10.6151
R1607 B.n623 B.n622 10.6151
R1608 B.n625 B.n623 10.6151
R1609 B.n626 B.n625 10.6151
R1610 B.n627 B.n626 10.6151
R1611 B.n628 B.n627 10.6151
R1612 B.n630 B.n628 10.6151
R1613 B.n631 B.n630 10.6151
R1614 B.n632 B.n631 10.6151
R1615 B.n633 B.n632 10.6151
R1616 B.n635 B.n633 10.6151
R1617 B.n636 B.n635 10.6151
R1618 B.n637 B.n636 10.6151
R1619 B.n638 B.n637 10.6151
R1620 B.n640 B.n638 10.6151
R1621 B.n641 B.n640 10.6151
R1622 B.n642 B.n641 10.6151
R1623 B.n643 B.n642 10.6151
R1624 B.n645 B.n643 10.6151
R1625 B.n646 B.n645 10.6151
R1626 B.n647 B.n646 10.6151
R1627 B.n648 B.n647 10.6151
R1628 B.n650 B.n648 10.6151
R1629 B.n651 B.n650 10.6151
R1630 B.n652 B.n651 10.6151
R1631 B.n653 B.n652 10.6151
R1632 B.n655 B.n653 10.6151
R1633 B.n656 B.n655 10.6151
R1634 B.n657 B.n656 10.6151
R1635 B.n658 B.n657 10.6151
R1636 B.n660 B.n658 10.6151
R1637 B.n661 B.n660 10.6151
R1638 B.n662 B.n661 10.6151
R1639 B.n663 B.n662 10.6151
R1640 B.n665 B.n663 10.6151
R1641 B.n666 B.n665 10.6151
R1642 B.n667 B.n666 10.6151
R1643 B.n668 B.n667 10.6151
R1644 B.n670 B.n668 10.6151
R1645 B.n671 B.n670 10.6151
R1646 B.n759 B.n1 10.6151
R1647 B.n759 B.n758 10.6151
R1648 B.n758 B.n757 10.6151
R1649 B.n757 B.n10 10.6151
R1650 B.n751 B.n10 10.6151
R1651 B.n751 B.n750 10.6151
R1652 B.n750 B.n749 10.6151
R1653 B.n749 B.n18 10.6151
R1654 B.n743 B.n18 10.6151
R1655 B.n743 B.n742 10.6151
R1656 B.n742 B.n741 10.6151
R1657 B.n741 B.n25 10.6151
R1658 B.n735 B.n25 10.6151
R1659 B.n735 B.n734 10.6151
R1660 B.n734 B.n733 10.6151
R1661 B.n733 B.n32 10.6151
R1662 B.n727 B.n32 10.6151
R1663 B.n727 B.n726 10.6151
R1664 B.n726 B.n725 10.6151
R1665 B.n725 B.n39 10.6151
R1666 B.n719 B.n39 10.6151
R1667 B.n719 B.n718 10.6151
R1668 B.n718 B.n717 10.6151
R1669 B.n717 B.n46 10.6151
R1670 B.n711 B.n46 10.6151
R1671 B.n711 B.n710 10.6151
R1672 B.n710 B.n709 10.6151
R1673 B.n709 B.n53 10.6151
R1674 B.n703 B.n53 10.6151
R1675 B.n703 B.n702 10.6151
R1676 B.n702 B.n701 10.6151
R1677 B.n701 B.n60 10.6151
R1678 B.n695 B.n60 10.6151
R1679 B.n695 B.n694 10.6151
R1680 B.n694 B.n693 10.6151
R1681 B.n693 B.n66 10.6151
R1682 B.n687 B.n66 10.6151
R1683 B.n687 B.n686 10.6151
R1684 B.n686 B.n685 10.6151
R1685 B.n685 B.n74 10.6151
R1686 B.n679 B.n74 10.6151
R1687 B.n679 B.n678 10.6151
R1688 B.n678 B.n677 10.6151
R1689 B.n120 B.n81 10.6151
R1690 B.n123 B.n120 10.6151
R1691 B.n124 B.n123 10.6151
R1692 B.n127 B.n124 10.6151
R1693 B.n128 B.n127 10.6151
R1694 B.n131 B.n128 10.6151
R1695 B.n132 B.n131 10.6151
R1696 B.n135 B.n132 10.6151
R1697 B.n136 B.n135 10.6151
R1698 B.n139 B.n136 10.6151
R1699 B.n140 B.n139 10.6151
R1700 B.n143 B.n140 10.6151
R1701 B.n144 B.n143 10.6151
R1702 B.n147 B.n144 10.6151
R1703 B.n148 B.n147 10.6151
R1704 B.n151 B.n148 10.6151
R1705 B.n152 B.n151 10.6151
R1706 B.n155 B.n152 10.6151
R1707 B.n156 B.n155 10.6151
R1708 B.n159 B.n156 10.6151
R1709 B.n160 B.n159 10.6151
R1710 B.n163 B.n160 10.6151
R1711 B.n164 B.n163 10.6151
R1712 B.n167 B.n164 10.6151
R1713 B.n168 B.n167 10.6151
R1714 B.n172 B.n171 10.6151
R1715 B.n175 B.n172 10.6151
R1716 B.n176 B.n175 10.6151
R1717 B.n179 B.n176 10.6151
R1718 B.n180 B.n179 10.6151
R1719 B.n183 B.n180 10.6151
R1720 B.n184 B.n183 10.6151
R1721 B.n187 B.n184 10.6151
R1722 B.n192 B.n189 10.6151
R1723 B.n193 B.n192 10.6151
R1724 B.n196 B.n193 10.6151
R1725 B.n197 B.n196 10.6151
R1726 B.n200 B.n197 10.6151
R1727 B.n201 B.n200 10.6151
R1728 B.n204 B.n201 10.6151
R1729 B.n205 B.n204 10.6151
R1730 B.n208 B.n205 10.6151
R1731 B.n209 B.n208 10.6151
R1732 B.n212 B.n209 10.6151
R1733 B.n213 B.n212 10.6151
R1734 B.n216 B.n213 10.6151
R1735 B.n217 B.n216 10.6151
R1736 B.n220 B.n217 10.6151
R1737 B.n221 B.n220 10.6151
R1738 B.n224 B.n221 10.6151
R1739 B.n225 B.n224 10.6151
R1740 B.n228 B.n225 10.6151
R1741 B.n229 B.n228 10.6151
R1742 B.n232 B.n229 10.6151
R1743 B.n233 B.n232 10.6151
R1744 B.n236 B.n233 10.6151
R1745 B.n237 B.n236 10.6151
R1746 B.n672 B.n237 10.6151
R1747 B.t3 B.n248 8.34437
R1748 B.t1 B.n16 8.34437
R1749 B.n767 B.n0 8.11757
R1750 B.n767 B.n1 8.11757
R1751 B.n407 B.n344 6.5566
R1752 B.n340 B.n339 6.5566
R1753 B.n171 B.n119 6.5566
R1754 B.n188 B.n187 6.5566
R1755 B.n408 B.n407 4.05904
R1756 B.n430 B.n339 4.05904
R1757 B.n168 B.n119 4.05904
R1758 B.n189 B.n188 4.05904
R1759 VP.n21 VP.n20 161.3
R1760 VP.n19 VP.n1 161.3
R1761 VP.n18 VP.n17 161.3
R1762 VP.n16 VP.n2 161.3
R1763 VP.n15 VP.n14 161.3
R1764 VP.n13 VP.n3 161.3
R1765 VP.n12 VP.n11 161.3
R1766 VP.n10 VP.n4 161.3
R1767 VP.n9 VP.n8 161.3
R1768 VP.n7 VP.n6 87.6207
R1769 VP.n22 VP.n0 87.6207
R1770 VP.n5 VP.t3 75.8783
R1771 VP.n5 VP.t0 74.5357
R1772 VP.n6 VP.n5 47.7117
R1773 VP.n7 VP.t1 42.1276
R1774 VP.n0 VP.t2 42.1276
R1775 VP.n14 VP.n13 40.4934
R1776 VP.n14 VP.n2 40.4934
R1777 VP.n8 VP.n4 24.4675
R1778 VP.n12 VP.n4 24.4675
R1779 VP.n13 VP.n12 24.4675
R1780 VP.n18 VP.n2 24.4675
R1781 VP.n19 VP.n18 24.4675
R1782 VP.n20 VP.n19 24.4675
R1783 VP.n8 VP.n7 2.4472
R1784 VP.n20 VP.n0 2.4472
R1785 VP.n9 VP.n6 0.354971
R1786 VP.n22 VP.n21 0.354971
R1787 VP VP.n22 0.26696
R1788 VP.n10 VP.n9 0.189894
R1789 VP.n11 VP.n10 0.189894
R1790 VP.n11 VP.n3 0.189894
R1791 VP.n15 VP.n3 0.189894
R1792 VP.n16 VP.n15 0.189894
R1793 VP.n17 VP.n16 0.189894
R1794 VP.n17 VP.n1 0.189894
R1795 VP.n21 VP.n1 0.189894
R1796 VDD1 VDD1.n1 110.397
R1797 VDD1 VDD1.n0 69.9317
R1798 VDD1.n0 VDD1.t0 3.00505
R1799 VDD1.n0 VDD1.t3 3.00505
R1800 VDD1.n1 VDD1.t2 3.00505
R1801 VDD1.n1 VDD1.t1 3.00505
C0 VP VDD1 3.23434f
C1 VTAIL VP 3.41693f
C2 VP VN 6.03381f
C3 VDD2 VP 0.468609f
C4 VTAIL VDD1 4.60812f
C5 VDD1 VN 0.149912f
C6 VTAIL VN 3.40282f
C7 VDD2 VDD1 1.30985f
C8 VDD2 VTAIL 4.67017f
C9 VDD2 VN 2.91667f
C10 VDD2 B 4.012885f
C11 VDD1 B 8.11826f
C12 VTAIL B 7.099483f
C13 VN B 12.47928f
C14 VP B 10.892694f
C15 VDD1.t0 B 0.149375f
C16 VDD1.t3 B 0.149375f
C17 VDD1.n0 B 1.2723f
C18 VDD1.t2 B 0.149375f
C19 VDD1.t1 B 0.149375f
C20 VDD1.n1 B 1.83298f
C21 VP.t2 B 1.54794f
C22 VP.n0 B 0.651716f
C23 VP.n1 B 0.023417f
C24 VP.n2 B 0.046541f
C25 VP.n3 B 0.023417f
C26 VP.n4 B 0.043643f
C27 VP.t3 B 1.88491f
C28 VP.t0 B 1.87195f
C29 VP.n5 B 2.48429f
C30 VP.n6 B 1.2657f
C31 VP.t1 B 1.54794f
C32 VP.n7 B 0.651716f
C33 VP.n8 B 0.024251f
C34 VP.n9 B 0.037794f
C35 VP.n10 B 0.023417f
C36 VP.n11 B 0.023417f
C37 VP.n12 B 0.043643f
C38 VP.n13 B 0.046541f
C39 VP.n14 B 0.01893f
C40 VP.n15 B 0.023417f
C41 VP.n16 B 0.023417f
C42 VP.n17 B 0.023417f
C43 VP.n18 B 0.043643f
C44 VP.n19 B 0.043643f
C45 VP.n20 B 0.024251f
C46 VP.n21 B 0.037794f
C47 VP.n22 B 0.071844f
C48 VDD2.t0 B 0.147549f
C49 VDD2.t3 B 0.147549f
C50 VDD2.n0 B 1.7855f
C51 VDD2.t1 B 0.147549f
C52 VDD2.t2 B 0.147549f
C53 VDD2.n1 B 1.25629f
C54 VDD2.n2 B 3.63924f
C55 VTAIL.n0 B 0.011507f
C56 VTAIL.n1 B 0.025891f
C57 VTAIL.n2 B 0.011598f
C58 VTAIL.n3 B 0.020385f
C59 VTAIL.n4 B 0.010954f
C60 VTAIL.n5 B 0.025891f
C61 VTAIL.n6 B 0.011598f
C62 VTAIL.n7 B 0.020385f
C63 VTAIL.n8 B 0.010954f
C64 VTAIL.n9 B 0.019419f
C65 VTAIL.n10 B 0.018303f
C66 VTAIL.t7 B 0.043198f
C67 VTAIL.n11 B 0.104746f
C68 VTAIL.n12 B 0.537693f
C69 VTAIL.n13 B 0.010954f
C70 VTAIL.n14 B 0.011598f
C71 VTAIL.n15 B 0.025891f
C72 VTAIL.n16 B 0.025891f
C73 VTAIL.n17 B 0.011598f
C74 VTAIL.n18 B 0.010954f
C75 VTAIL.n19 B 0.020385f
C76 VTAIL.n20 B 0.020385f
C77 VTAIL.n21 B 0.010954f
C78 VTAIL.n22 B 0.011598f
C79 VTAIL.n23 B 0.025891f
C80 VTAIL.n24 B 0.025891f
C81 VTAIL.n25 B 0.011598f
C82 VTAIL.n26 B 0.010954f
C83 VTAIL.n27 B 0.020385f
C84 VTAIL.n28 B 0.053524f
C85 VTAIL.n29 B 0.010954f
C86 VTAIL.n30 B 0.011598f
C87 VTAIL.n31 B 0.053861f
C88 VTAIL.n32 B 0.045679f
C89 VTAIL.n33 B 0.171485f
C90 VTAIL.n34 B 0.011507f
C91 VTAIL.n35 B 0.025891f
C92 VTAIL.n36 B 0.011598f
C93 VTAIL.n37 B 0.020385f
C94 VTAIL.n38 B 0.010954f
C95 VTAIL.n39 B 0.025891f
C96 VTAIL.n40 B 0.011598f
C97 VTAIL.n41 B 0.020385f
C98 VTAIL.n42 B 0.010954f
C99 VTAIL.n43 B 0.019419f
C100 VTAIL.n44 B 0.018303f
C101 VTAIL.t3 B 0.043198f
C102 VTAIL.n45 B 0.104746f
C103 VTAIL.n46 B 0.537693f
C104 VTAIL.n47 B 0.010954f
C105 VTAIL.n48 B 0.011598f
C106 VTAIL.n49 B 0.025891f
C107 VTAIL.n50 B 0.025891f
C108 VTAIL.n51 B 0.011598f
C109 VTAIL.n52 B 0.010954f
C110 VTAIL.n53 B 0.020385f
C111 VTAIL.n54 B 0.020385f
C112 VTAIL.n55 B 0.010954f
C113 VTAIL.n56 B 0.011598f
C114 VTAIL.n57 B 0.025891f
C115 VTAIL.n58 B 0.025891f
C116 VTAIL.n59 B 0.011598f
C117 VTAIL.n60 B 0.010954f
C118 VTAIL.n61 B 0.020385f
C119 VTAIL.n62 B 0.053524f
C120 VTAIL.n63 B 0.010954f
C121 VTAIL.n64 B 0.011598f
C122 VTAIL.n65 B 0.053861f
C123 VTAIL.n66 B 0.045679f
C124 VTAIL.n67 B 0.283744f
C125 VTAIL.n68 B 0.011507f
C126 VTAIL.n69 B 0.025891f
C127 VTAIL.n70 B 0.011598f
C128 VTAIL.n71 B 0.020385f
C129 VTAIL.n72 B 0.010954f
C130 VTAIL.n73 B 0.025891f
C131 VTAIL.n74 B 0.011598f
C132 VTAIL.n75 B 0.020385f
C133 VTAIL.n76 B 0.010954f
C134 VTAIL.n77 B 0.019419f
C135 VTAIL.n78 B 0.018303f
C136 VTAIL.t2 B 0.043198f
C137 VTAIL.n79 B 0.104746f
C138 VTAIL.n80 B 0.537693f
C139 VTAIL.n81 B 0.010954f
C140 VTAIL.n82 B 0.011598f
C141 VTAIL.n83 B 0.025891f
C142 VTAIL.n84 B 0.025891f
C143 VTAIL.n85 B 0.011598f
C144 VTAIL.n86 B 0.010954f
C145 VTAIL.n87 B 0.020385f
C146 VTAIL.n88 B 0.020385f
C147 VTAIL.n89 B 0.010954f
C148 VTAIL.n90 B 0.011598f
C149 VTAIL.n91 B 0.025891f
C150 VTAIL.n92 B 0.025891f
C151 VTAIL.n93 B 0.011598f
C152 VTAIL.n94 B 0.010954f
C153 VTAIL.n95 B 0.020385f
C154 VTAIL.n96 B 0.053524f
C155 VTAIL.n97 B 0.010954f
C156 VTAIL.n98 B 0.011598f
C157 VTAIL.n99 B 0.053861f
C158 VTAIL.n100 B 0.045679f
C159 VTAIL.n101 B 1.13511f
C160 VTAIL.n102 B 0.011507f
C161 VTAIL.n103 B 0.025891f
C162 VTAIL.n104 B 0.011598f
C163 VTAIL.n105 B 0.020385f
C164 VTAIL.n106 B 0.010954f
C165 VTAIL.n107 B 0.025891f
C166 VTAIL.n108 B 0.011598f
C167 VTAIL.n109 B 0.020385f
C168 VTAIL.n110 B 0.010954f
C169 VTAIL.n111 B 0.019419f
C170 VTAIL.n112 B 0.018303f
C171 VTAIL.t4 B 0.043198f
C172 VTAIL.n113 B 0.104746f
C173 VTAIL.n114 B 0.537693f
C174 VTAIL.n115 B 0.010954f
C175 VTAIL.n116 B 0.011598f
C176 VTAIL.n117 B 0.025891f
C177 VTAIL.n118 B 0.025891f
C178 VTAIL.n119 B 0.011598f
C179 VTAIL.n120 B 0.010954f
C180 VTAIL.n121 B 0.020385f
C181 VTAIL.n122 B 0.020385f
C182 VTAIL.n123 B 0.010954f
C183 VTAIL.n124 B 0.011598f
C184 VTAIL.n125 B 0.025891f
C185 VTAIL.n126 B 0.025891f
C186 VTAIL.n127 B 0.011598f
C187 VTAIL.n128 B 0.010954f
C188 VTAIL.n129 B 0.020385f
C189 VTAIL.n130 B 0.053524f
C190 VTAIL.n131 B 0.010954f
C191 VTAIL.n132 B 0.011598f
C192 VTAIL.n133 B 0.053861f
C193 VTAIL.n134 B 0.045679f
C194 VTAIL.n135 B 1.13511f
C195 VTAIL.n136 B 0.011507f
C196 VTAIL.n137 B 0.025891f
C197 VTAIL.n138 B 0.011598f
C198 VTAIL.n139 B 0.020385f
C199 VTAIL.n140 B 0.010954f
C200 VTAIL.n141 B 0.025891f
C201 VTAIL.n142 B 0.011598f
C202 VTAIL.n143 B 0.020385f
C203 VTAIL.n144 B 0.010954f
C204 VTAIL.n145 B 0.019419f
C205 VTAIL.n146 B 0.018303f
C206 VTAIL.t6 B 0.043198f
C207 VTAIL.n147 B 0.104746f
C208 VTAIL.n148 B 0.537693f
C209 VTAIL.n149 B 0.010954f
C210 VTAIL.n150 B 0.011598f
C211 VTAIL.n151 B 0.025891f
C212 VTAIL.n152 B 0.025891f
C213 VTAIL.n153 B 0.011598f
C214 VTAIL.n154 B 0.010954f
C215 VTAIL.n155 B 0.020385f
C216 VTAIL.n156 B 0.020385f
C217 VTAIL.n157 B 0.010954f
C218 VTAIL.n158 B 0.011598f
C219 VTAIL.n159 B 0.025891f
C220 VTAIL.n160 B 0.025891f
C221 VTAIL.n161 B 0.011598f
C222 VTAIL.n162 B 0.010954f
C223 VTAIL.n163 B 0.020385f
C224 VTAIL.n164 B 0.053524f
C225 VTAIL.n165 B 0.010954f
C226 VTAIL.n166 B 0.011598f
C227 VTAIL.n167 B 0.053861f
C228 VTAIL.n168 B 0.045679f
C229 VTAIL.n169 B 0.283744f
C230 VTAIL.n170 B 0.011507f
C231 VTAIL.n171 B 0.025891f
C232 VTAIL.n172 B 0.011598f
C233 VTAIL.n173 B 0.020385f
C234 VTAIL.n174 B 0.010954f
C235 VTAIL.n175 B 0.025891f
C236 VTAIL.n176 B 0.011598f
C237 VTAIL.n177 B 0.020385f
C238 VTAIL.n178 B 0.010954f
C239 VTAIL.n179 B 0.019419f
C240 VTAIL.n180 B 0.018303f
C241 VTAIL.t1 B 0.043198f
C242 VTAIL.n181 B 0.104746f
C243 VTAIL.n182 B 0.537693f
C244 VTAIL.n183 B 0.010954f
C245 VTAIL.n184 B 0.011598f
C246 VTAIL.n185 B 0.025891f
C247 VTAIL.n186 B 0.025891f
C248 VTAIL.n187 B 0.011598f
C249 VTAIL.n188 B 0.010954f
C250 VTAIL.n189 B 0.020385f
C251 VTAIL.n190 B 0.020385f
C252 VTAIL.n191 B 0.010954f
C253 VTAIL.n192 B 0.011598f
C254 VTAIL.n193 B 0.025891f
C255 VTAIL.n194 B 0.025891f
C256 VTAIL.n195 B 0.011598f
C257 VTAIL.n196 B 0.010954f
C258 VTAIL.n197 B 0.020385f
C259 VTAIL.n198 B 0.053524f
C260 VTAIL.n199 B 0.010954f
C261 VTAIL.n200 B 0.011598f
C262 VTAIL.n201 B 0.053861f
C263 VTAIL.n202 B 0.045679f
C264 VTAIL.n203 B 0.283744f
C265 VTAIL.n204 B 0.011507f
C266 VTAIL.n205 B 0.025891f
C267 VTAIL.n206 B 0.011598f
C268 VTAIL.n207 B 0.020385f
C269 VTAIL.n208 B 0.010954f
C270 VTAIL.n209 B 0.025891f
C271 VTAIL.n210 B 0.011598f
C272 VTAIL.n211 B 0.020385f
C273 VTAIL.n212 B 0.010954f
C274 VTAIL.n213 B 0.019419f
C275 VTAIL.n214 B 0.018303f
C276 VTAIL.t0 B 0.043198f
C277 VTAIL.n215 B 0.104746f
C278 VTAIL.n216 B 0.537693f
C279 VTAIL.n217 B 0.010954f
C280 VTAIL.n218 B 0.011598f
C281 VTAIL.n219 B 0.025891f
C282 VTAIL.n220 B 0.025891f
C283 VTAIL.n221 B 0.011598f
C284 VTAIL.n222 B 0.010954f
C285 VTAIL.n223 B 0.020385f
C286 VTAIL.n224 B 0.020385f
C287 VTAIL.n225 B 0.010954f
C288 VTAIL.n226 B 0.011598f
C289 VTAIL.n227 B 0.025891f
C290 VTAIL.n228 B 0.025891f
C291 VTAIL.n229 B 0.011598f
C292 VTAIL.n230 B 0.010954f
C293 VTAIL.n231 B 0.020385f
C294 VTAIL.n232 B 0.053524f
C295 VTAIL.n233 B 0.010954f
C296 VTAIL.n234 B 0.011598f
C297 VTAIL.n235 B 0.053861f
C298 VTAIL.n236 B 0.045679f
C299 VTAIL.n237 B 1.13511f
C300 VTAIL.n238 B 0.011507f
C301 VTAIL.n239 B 0.025891f
C302 VTAIL.n240 B 0.011598f
C303 VTAIL.n241 B 0.020385f
C304 VTAIL.n242 B 0.010954f
C305 VTAIL.n243 B 0.025891f
C306 VTAIL.n244 B 0.011598f
C307 VTAIL.n245 B 0.020385f
C308 VTAIL.n246 B 0.010954f
C309 VTAIL.n247 B 0.019419f
C310 VTAIL.n248 B 0.018303f
C311 VTAIL.t5 B 0.043198f
C312 VTAIL.n249 B 0.104746f
C313 VTAIL.n250 B 0.537693f
C314 VTAIL.n251 B 0.010954f
C315 VTAIL.n252 B 0.011598f
C316 VTAIL.n253 B 0.025891f
C317 VTAIL.n254 B 0.025891f
C318 VTAIL.n255 B 0.011598f
C319 VTAIL.n256 B 0.010954f
C320 VTAIL.n257 B 0.020385f
C321 VTAIL.n258 B 0.020385f
C322 VTAIL.n259 B 0.010954f
C323 VTAIL.n260 B 0.011598f
C324 VTAIL.n261 B 0.025891f
C325 VTAIL.n262 B 0.025891f
C326 VTAIL.n263 B 0.011598f
C327 VTAIL.n264 B 0.010954f
C328 VTAIL.n265 B 0.020385f
C329 VTAIL.n266 B 0.053524f
C330 VTAIL.n267 B 0.010954f
C331 VTAIL.n268 B 0.011598f
C332 VTAIL.n269 B 0.053861f
C333 VTAIL.n270 B 0.045679f
C334 VTAIL.n271 B 1.01521f
C335 VN.t0 B 1.82261f
C336 VN.t3 B 1.83524f
C337 VN.n0 B 1.08364f
C338 VN.t2 B 1.82261f
C339 VN.t1 B 1.83524f
C340 VN.n1 B 2.42826f
.ends

