* NGSPICE file created from diff_pair_sample_0616.ext - technology: sky130A

.subckt diff_pair_sample_0616 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2358_n3650# sky130_fd_pr__pfet_01v8 ad=5.2299 pd=27.6 as=0 ps=0 w=13.41 l=3.14
X1 VDD1.t1 VP.t0 VTAIL.t2 w_n2358_n3650# sky130_fd_pr__pfet_01v8 ad=5.2299 pd=27.6 as=5.2299 ps=27.6 w=13.41 l=3.14
X2 B.t8 B.t6 B.t7 w_n2358_n3650# sky130_fd_pr__pfet_01v8 ad=5.2299 pd=27.6 as=0 ps=0 w=13.41 l=3.14
X3 VDD2.t1 VN.t0 VTAIL.t0 w_n2358_n3650# sky130_fd_pr__pfet_01v8 ad=5.2299 pd=27.6 as=5.2299 ps=27.6 w=13.41 l=3.14
X4 VDD1.t0 VP.t1 VTAIL.t3 w_n2358_n3650# sky130_fd_pr__pfet_01v8 ad=5.2299 pd=27.6 as=5.2299 ps=27.6 w=13.41 l=3.14
X5 B.t5 B.t3 B.t4 w_n2358_n3650# sky130_fd_pr__pfet_01v8 ad=5.2299 pd=27.6 as=0 ps=0 w=13.41 l=3.14
X6 B.t2 B.t0 B.t1 w_n2358_n3650# sky130_fd_pr__pfet_01v8 ad=5.2299 pd=27.6 as=0 ps=0 w=13.41 l=3.14
X7 VDD2.t0 VN.t1 VTAIL.t1 w_n2358_n3650# sky130_fd_pr__pfet_01v8 ad=5.2299 pd=27.6 as=5.2299 ps=27.6 w=13.41 l=3.14
R0 B.n361 B.n360 585
R1 B.n359 B.n100 585
R2 B.n358 B.n357 585
R3 B.n356 B.n101 585
R4 B.n355 B.n354 585
R5 B.n353 B.n102 585
R6 B.n352 B.n351 585
R7 B.n350 B.n103 585
R8 B.n349 B.n348 585
R9 B.n347 B.n104 585
R10 B.n346 B.n345 585
R11 B.n344 B.n105 585
R12 B.n343 B.n342 585
R13 B.n341 B.n106 585
R14 B.n340 B.n339 585
R15 B.n338 B.n107 585
R16 B.n337 B.n336 585
R17 B.n335 B.n108 585
R18 B.n334 B.n333 585
R19 B.n332 B.n109 585
R20 B.n331 B.n330 585
R21 B.n329 B.n110 585
R22 B.n328 B.n327 585
R23 B.n326 B.n111 585
R24 B.n325 B.n324 585
R25 B.n323 B.n112 585
R26 B.n322 B.n321 585
R27 B.n320 B.n113 585
R28 B.n319 B.n318 585
R29 B.n317 B.n114 585
R30 B.n316 B.n315 585
R31 B.n314 B.n115 585
R32 B.n313 B.n312 585
R33 B.n311 B.n116 585
R34 B.n310 B.n309 585
R35 B.n308 B.n117 585
R36 B.n307 B.n306 585
R37 B.n305 B.n118 585
R38 B.n304 B.n303 585
R39 B.n302 B.n119 585
R40 B.n301 B.n300 585
R41 B.n299 B.n120 585
R42 B.n298 B.n297 585
R43 B.n296 B.n121 585
R44 B.n295 B.n294 585
R45 B.n293 B.n122 585
R46 B.n292 B.n291 585
R47 B.n287 B.n123 585
R48 B.n286 B.n285 585
R49 B.n284 B.n124 585
R50 B.n283 B.n282 585
R51 B.n281 B.n125 585
R52 B.n280 B.n279 585
R53 B.n278 B.n126 585
R54 B.n277 B.n276 585
R55 B.n274 B.n127 585
R56 B.n273 B.n272 585
R57 B.n271 B.n130 585
R58 B.n270 B.n269 585
R59 B.n268 B.n131 585
R60 B.n267 B.n266 585
R61 B.n265 B.n132 585
R62 B.n264 B.n263 585
R63 B.n262 B.n133 585
R64 B.n261 B.n260 585
R65 B.n259 B.n134 585
R66 B.n258 B.n257 585
R67 B.n256 B.n135 585
R68 B.n255 B.n254 585
R69 B.n253 B.n136 585
R70 B.n252 B.n251 585
R71 B.n250 B.n137 585
R72 B.n249 B.n248 585
R73 B.n247 B.n138 585
R74 B.n246 B.n245 585
R75 B.n244 B.n139 585
R76 B.n243 B.n242 585
R77 B.n241 B.n140 585
R78 B.n240 B.n239 585
R79 B.n238 B.n141 585
R80 B.n237 B.n236 585
R81 B.n235 B.n142 585
R82 B.n234 B.n233 585
R83 B.n232 B.n143 585
R84 B.n231 B.n230 585
R85 B.n229 B.n144 585
R86 B.n228 B.n227 585
R87 B.n226 B.n145 585
R88 B.n225 B.n224 585
R89 B.n223 B.n146 585
R90 B.n222 B.n221 585
R91 B.n220 B.n147 585
R92 B.n219 B.n218 585
R93 B.n217 B.n148 585
R94 B.n216 B.n215 585
R95 B.n214 B.n149 585
R96 B.n213 B.n212 585
R97 B.n211 B.n150 585
R98 B.n210 B.n209 585
R99 B.n208 B.n151 585
R100 B.n207 B.n206 585
R101 B.n362 B.n99 585
R102 B.n364 B.n363 585
R103 B.n365 B.n98 585
R104 B.n367 B.n366 585
R105 B.n368 B.n97 585
R106 B.n370 B.n369 585
R107 B.n371 B.n96 585
R108 B.n373 B.n372 585
R109 B.n374 B.n95 585
R110 B.n376 B.n375 585
R111 B.n377 B.n94 585
R112 B.n379 B.n378 585
R113 B.n380 B.n93 585
R114 B.n382 B.n381 585
R115 B.n383 B.n92 585
R116 B.n385 B.n384 585
R117 B.n386 B.n91 585
R118 B.n388 B.n387 585
R119 B.n389 B.n90 585
R120 B.n391 B.n390 585
R121 B.n392 B.n89 585
R122 B.n394 B.n393 585
R123 B.n395 B.n88 585
R124 B.n397 B.n396 585
R125 B.n398 B.n87 585
R126 B.n400 B.n399 585
R127 B.n401 B.n86 585
R128 B.n403 B.n402 585
R129 B.n404 B.n85 585
R130 B.n406 B.n405 585
R131 B.n407 B.n84 585
R132 B.n409 B.n408 585
R133 B.n410 B.n83 585
R134 B.n412 B.n411 585
R135 B.n413 B.n82 585
R136 B.n415 B.n414 585
R137 B.n416 B.n81 585
R138 B.n418 B.n417 585
R139 B.n419 B.n80 585
R140 B.n421 B.n420 585
R141 B.n422 B.n79 585
R142 B.n424 B.n423 585
R143 B.n425 B.n78 585
R144 B.n427 B.n426 585
R145 B.n428 B.n77 585
R146 B.n430 B.n429 585
R147 B.n431 B.n76 585
R148 B.n433 B.n432 585
R149 B.n434 B.n75 585
R150 B.n436 B.n435 585
R151 B.n437 B.n74 585
R152 B.n439 B.n438 585
R153 B.n440 B.n73 585
R154 B.n442 B.n441 585
R155 B.n443 B.n72 585
R156 B.n445 B.n444 585
R157 B.n446 B.n71 585
R158 B.n448 B.n447 585
R159 B.n601 B.n16 585
R160 B.n600 B.n599 585
R161 B.n598 B.n17 585
R162 B.n597 B.n596 585
R163 B.n595 B.n18 585
R164 B.n594 B.n593 585
R165 B.n592 B.n19 585
R166 B.n591 B.n590 585
R167 B.n589 B.n20 585
R168 B.n588 B.n587 585
R169 B.n586 B.n21 585
R170 B.n585 B.n584 585
R171 B.n583 B.n22 585
R172 B.n582 B.n581 585
R173 B.n580 B.n23 585
R174 B.n579 B.n578 585
R175 B.n577 B.n24 585
R176 B.n576 B.n575 585
R177 B.n574 B.n25 585
R178 B.n573 B.n572 585
R179 B.n571 B.n26 585
R180 B.n570 B.n569 585
R181 B.n568 B.n27 585
R182 B.n567 B.n566 585
R183 B.n565 B.n28 585
R184 B.n564 B.n563 585
R185 B.n562 B.n29 585
R186 B.n561 B.n560 585
R187 B.n559 B.n30 585
R188 B.n558 B.n557 585
R189 B.n556 B.n31 585
R190 B.n555 B.n554 585
R191 B.n553 B.n32 585
R192 B.n552 B.n551 585
R193 B.n550 B.n33 585
R194 B.n549 B.n548 585
R195 B.n547 B.n34 585
R196 B.n546 B.n545 585
R197 B.n544 B.n35 585
R198 B.n543 B.n542 585
R199 B.n541 B.n36 585
R200 B.n540 B.n539 585
R201 B.n538 B.n37 585
R202 B.n537 B.n536 585
R203 B.n535 B.n38 585
R204 B.n534 B.n533 585
R205 B.n531 B.n39 585
R206 B.n530 B.n529 585
R207 B.n528 B.n42 585
R208 B.n527 B.n526 585
R209 B.n525 B.n43 585
R210 B.n524 B.n523 585
R211 B.n522 B.n44 585
R212 B.n521 B.n520 585
R213 B.n519 B.n45 585
R214 B.n517 B.n516 585
R215 B.n515 B.n48 585
R216 B.n514 B.n513 585
R217 B.n512 B.n49 585
R218 B.n511 B.n510 585
R219 B.n509 B.n50 585
R220 B.n508 B.n507 585
R221 B.n506 B.n51 585
R222 B.n505 B.n504 585
R223 B.n503 B.n52 585
R224 B.n502 B.n501 585
R225 B.n500 B.n53 585
R226 B.n499 B.n498 585
R227 B.n497 B.n54 585
R228 B.n496 B.n495 585
R229 B.n494 B.n55 585
R230 B.n493 B.n492 585
R231 B.n491 B.n56 585
R232 B.n490 B.n489 585
R233 B.n488 B.n57 585
R234 B.n487 B.n486 585
R235 B.n485 B.n58 585
R236 B.n484 B.n483 585
R237 B.n482 B.n59 585
R238 B.n481 B.n480 585
R239 B.n479 B.n60 585
R240 B.n478 B.n477 585
R241 B.n476 B.n61 585
R242 B.n475 B.n474 585
R243 B.n473 B.n62 585
R244 B.n472 B.n471 585
R245 B.n470 B.n63 585
R246 B.n469 B.n468 585
R247 B.n467 B.n64 585
R248 B.n466 B.n465 585
R249 B.n464 B.n65 585
R250 B.n463 B.n462 585
R251 B.n461 B.n66 585
R252 B.n460 B.n459 585
R253 B.n458 B.n67 585
R254 B.n457 B.n456 585
R255 B.n455 B.n68 585
R256 B.n454 B.n453 585
R257 B.n452 B.n69 585
R258 B.n451 B.n450 585
R259 B.n449 B.n70 585
R260 B.n603 B.n602 585
R261 B.n604 B.n15 585
R262 B.n606 B.n605 585
R263 B.n607 B.n14 585
R264 B.n609 B.n608 585
R265 B.n610 B.n13 585
R266 B.n612 B.n611 585
R267 B.n613 B.n12 585
R268 B.n615 B.n614 585
R269 B.n616 B.n11 585
R270 B.n618 B.n617 585
R271 B.n619 B.n10 585
R272 B.n621 B.n620 585
R273 B.n622 B.n9 585
R274 B.n624 B.n623 585
R275 B.n625 B.n8 585
R276 B.n627 B.n626 585
R277 B.n628 B.n7 585
R278 B.n630 B.n629 585
R279 B.n631 B.n6 585
R280 B.n633 B.n632 585
R281 B.n634 B.n5 585
R282 B.n636 B.n635 585
R283 B.n637 B.n4 585
R284 B.n639 B.n638 585
R285 B.n640 B.n3 585
R286 B.n642 B.n641 585
R287 B.n643 B.n0 585
R288 B.n2 B.n1 585
R289 B.n166 B.n165 585
R290 B.n168 B.n167 585
R291 B.n169 B.n164 585
R292 B.n171 B.n170 585
R293 B.n172 B.n163 585
R294 B.n174 B.n173 585
R295 B.n175 B.n162 585
R296 B.n177 B.n176 585
R297 B.n178 B.n161 585
R298 B.n180 B.n179 585
R299 B.n181 B.n160 585
R300 B.n183 B.n182 585
R301 B.n184 B.n159 585
R302 B.n186 B.n185 585
R303 B.n187 B.n158 585
R304 B.n189 B.n188 585
R305 B.n190 B.n157 585
R306 B.n192 B.n191 585
R307 B.n193 B.n156 585
R308 B.n195 B.n194 585
R309 B.n196 B.n155 585
R310 B.n198 B.n197 585
R311 B.n199 B.n154 585
R312 B.n201 B.n200 585
R313 B.n202 B.n153 585
R314 B.n204 B.n203 585
R315 B.n205 B.n152 585
R316 B.n206 B.n205 511.721
R317 B.n360 B.n99 511.721
R318 B.n449 B.n448 511.721
R319 B.n602 B.n601 511.721
R320 B.n288 B.t10 468.291
R321 B.n46 B.t8 468.291
R322 B.n128 B.t4 468.291
R323 B.n40 B.t2 468.291
R324 B.n289 B.t11 400.995
R325 B.n47 B.t7 400.995
R326 B.n129 B.t5 400.993
R327 B.n41 B.t1 400.993
R328 B.n128 B.t3 311.663
R329 B.n288 B.t9 311.663
R330 B.n46 B.t6 311.663
R331 B.n40 B.t0 311.663
R332 B.n645 B.n644 256.663
R333 B.n644 B.n643 235.042
R334 B.n644 B.n2 235.042
R335 B.n206 B.n151 163.367
R336 B.n210 B.n151 163.367
R337 B.n211 B.n210 163.367
R338 B.n212 B.n211 163.367
R339 B.n212 B.n149 163.367
R340 B.n216 B.n149 163.367
R341 B.n217 B.n216 163.367
R342 B.n218 B.n217 163.367
R343 B.n218 B.n147 163.367
R344 B.n222 B.n147 163.367
R345 B.n223 B.n222 163.367
R346 B.n224 B.n223 163.367
R347 B.n224 B.n145 163.367
R348 B.n228 B.n145 163.367
R349 B.n229 B.n228 163.367
R350 B.n230 B.n229 163.367
R351 B.n230 B.n143 163.367
R352 B.n234 B.n143 163.367
R353 B.n235 B.n234 163.367
R354 B.n236 B.n235 163.367
R355 B.n236 B.n141 163.367
R356 B.n240 B.n141 163.367
R357 B.n241 B.n240 163.367
R358 B.n242 B.n241 163.367
R359 B.n242 B.n139 163.367
R360 B.n246 B.n139 163.367
R361 B.n247 B.n246 163.367
R362 B.n248 B.n247 163.367
R363 B.n248 B.n137 163.367
R364 B.n252 B.n137 163.367
R365 B.n253 B.n252 163.367
R366 B.n254 B.n253 163.367
R367 B.n254 B.n135 163.367
R368 B.n258 B.n135 163.367
R369 B.n259 B.n258 163.367
R370 B.n260 B.n259 163.367
R371 B.n260 B.n133 163.367
R372 B.n264 B.n133 163.367
R373 B.n265 B.n264 163.367
R374 B.n266 B.n265 163.367
R375 B.n266 B.n131 163.367
R376 B.n270 B.n131 163.367
R377 B.n271 B.n270 163.367
R378 B.n272 B.n271 163.367
R379 B.n272 B.n127 163.367
R380 B.n277 B.n127 163.367
R381 B.n278 B.n277 163.367
R382 B.n279 B.n278 163.367
R383 B.n279 B.n125 163.367
R384 B.n283 B.n125 163.367
R385 B.n284 B.n283 163.367
R386 B.n285 B.n284 163.367
R387 B.n285 B.n123 163.367
R388 B.n292 B.n123 163.367
R389 B.n293 B.n292 163.367
R390 B.n294 B.n293 163.367
R391 B.n294 B.n121 163.367
R392 B.n298 B.n121 163.367
R393 B.n299 B.n298 163.367
R394 B.n300 B.n299 163.367
R395 B.n300 B.n119 163.367
R396 B.n304 B.n119 163.367
R397 B.n305 B.n304 163.367
R398 B.n306 B.n305 163.367
R399 B.n306 B.n117 163.367
R400 B.n310 B.n117 163.367
R401 B.n311 B.n310 163.367
R402 B.n312 B.n311 163.367
R403 B.n312 B.n115 163.367
R404 B.n316 B.n115 163.367
R405 B.n317 B.n316 163.367
R406 B.n318 B.n317 163.367
R407 B.n318 B.n113 163.367
R408 B.n322 B.n113 163.367
R409 B.n323 B.n322 163.367
R410 B.n324 B.n323 163.367
R411 B.n324 B.n111 163.367
R412 B.n328 B.n111 163.367
R413 B.n329 B.n328 163.367
R414 B.n330 B.n329 163.367
R415 B.n330 B.n109 163.367
R416 B.n334 B.n109 163.367
R417 B.n335 B.n334 163.367
R418 B.n336 B.n335 163.367
R419 B.n336 B.n107 163.367
R420 B.n340 B.n107 163.367
R421 B.n341 B.n340 163.367
R422 B.n342 B.n341 163.367
R423 B.n342 B.n105 163.367
R424 B.n346 B.n105 163.367
R425 B.n347 B.n346 163.367
R426 B.n348 B.n347 163.367
R427 B.n348 B.n103 163.367
R428 B.n352 B.n103 163.367
R429 B.n353 B.n352 163.367
R430 B.n354 B.n353 163.367
R431 B.n354 B.n101 163.367
R432 B.n358 B.n101 163.367
R433 B.n359 B.n358 163.367
R434 B.n360 B.n359 163.367
R435 B.n448 B.n71 163.367
R436 B.n444 B.n71 163.367
R437 B.n444 B.n443 163.367
R438 B.n443 B.n442 163.367
R439 B.n442 B.n73 163.367
R440 B.n438 B.n73 163.367
R441 B.n438 B.n437 163.367
R442 B.n437 B.n436 163.367
R443 B.n436 B.n75 163.367
R444 B.n432 B.n75 163.367
R445 B.n432 B.n431 163.367
R446 B.n431 B.n430 163.367
R447 B.n430 B.n77 163.367
R448 B.n426 B.n77 163.367
R449 B.n426 B.n425 163.367
R450 B.n425 B.n424 163.367
R451 B.n424 B.n79 163.367
R452 B.n420 B.n79 163.367
R453 B.n420 B.n419 163.367
R454 B.n419 B.n418 163.367
R455 B.n418 B.n81 163.367
R456 B.n414 B.n81 163.367
R457 B.n414 B.n413 163.367
R458 B.n413 B.n412 163.367
R459 B.n412 B.n83 163.367
R460 B.n408 B.n83 163.367
R461 B.n408 B.n407 163.367
R462 B.n407 B.n406 163.367
R463 B.n406 B.n85 163.367
R464 B.n402 B.n85 163.367
R465 B.n402 B.n401 163.367
R466 B.n401 B.n400 163.367
R467 B.n400 B.n87 163.367
R468 B.n396 B.n87 163.367
R469 B.n396 B.n395 163.367
R470 B.n395 B.n394 163.367
R471 B.n394 B.n89 163.367
R472 B.n390 B.n89 163.367
R473 B.n390 B.n389 163.367
R474 B.n389 B.n388 163.367
R475 B.n388 B.n91 163.367
R476 B.n384 B.n91 163.367
R477 B.n384 B.n383 163.367
R478 B.n383 B.n382 163.367
R479 B.n382 B.n93 163.367
R480 B.n378 B.n93 163.367
R481 B.n378 B.n377 163.367
R482 B.n377 B.n376 163.367
R483 B.n376 B.n95 163.367
R484 B.n372 B.n95 163.367
R485 B.n372 B.n371 163.367
R486 B.n371 B.n370 163.367
R487 B.n370 B.n97 163.367
R488 B.n366 B.n97 163.367
R489 B.n366 B.n365 163.367
R490 B.n365 B.n364 163.367
R491 B.n364 B.n99 163.367
R492 B.n601 B.n600 163.367
R493 B.n600 B.n17 163.367
R494 B.n596 B.n17 163.367
R495 B.n596 B.n595 163.367
R496 B.n595 B.n594 163.367
R497 B.n594 B.n19 163.367
R498 B.n590 B.n19 163.367
R499 B.n590 B.n589 163.367
R500 B.n589 B.n588 163.367
R501 B.n588 B.n21 163.367
R502 B.n584 B.n21 163.367
R503 B.n584 B.n583 163.367
R504 B.n583 B.n582 163.367
R505 B.n582 B.n23 163.367
R506 B.n578 B.n23 163.367
R507 B.n578 B.n577 163.367
R508 B.n577 B.n576 163.367
R509 B.n576 B.n25 163.367
R510 B.n572 B.n25 163.367
R511 B.n572 B.n571 163.367
R512 B.n571 B.n570 163.367
R513 B.n570 B.n27 163.367
R514 B.n566 B.n27 163.367
R515 B.n566 B.n565 163.367
R516 B.n565 B.n564 163.367
R517 B.n564 B.n29 163.367
R518 B.n560 B.n29 163.367
R519 B.n560 B.n559 163.367
R520 B.n559 B.n558 163.367
R521 B.n558 B.n31 163.367
R522 B.n554 B.n31 163.367
R523 B.n554 B.n553 163.367
R524 B.n553 B.n552 163.367
R525 B.n552 B.n33 163.367
R526 B.n548 B.n33 163.367
R527 B.n548 B.n547 163.367
R528 B.n547 B.n546 163.367
R529 B.n546 B.n35 163.367
R530 B.n542 B.n35 163.367
R531 B.n542 B.n541 163.367
R532 B.n541 B.n540 163.367
R533 B.n540 B.n37 163.367
R534 B.n536 B.n37 163.367
R535 B.n536 B.n535 163.367
R536 B.n535 B.n534 163.367
R537 B.n534 B.n39 163.367
R538 B.n529 B.n39 163.367
R539 B.n529 B.n528 163.367
R540 B.n528 B.n527 163.367
R541 B.n527 B.n43 163.367
R542 B.n523 B.n43 163.367
R543 B.n523 B.n522 163.367
R544 B.n522 B.n521 163.367
R545 B.n521 B.n45 163.367
R546 B.n516 B.n45 163.367
R547 B.n516 B.n515 163.367
R548 B.n515 B.n514 163.367
R549 B.n514 B.n49 163.367
R550 B.n510 B.n49 163.367
R551 B.n510 B.n509 163.367
R552 B.n509 B.n508 163.367
R553 B.n508 B.n51 163.367
R554 B.n504 B.n51 163.367
R555 B.n504 B.n503 163.367
R556 B.n503 B.n502 163.367
R557 B.n502 B.n53 163.367
R558 B.n498 B.n53 163.367
R559 B.n498 B.n497 163.367
R560 B.n497 B.n496 163.367
R561 B.n496 B.n55 163.367
R562 B.n492 B.n55 163.367
R563 B.n492 B.n491 163.367
R564 B.n491 B.n490 163.367
R565 B.n490 B.n57 163.367
R566 B.n486 B.n57 163.367
R567 B.n486 B.n485 163.367
R568 B.n485 B.n484 163.367
R569 B.n484 B.n59 163.367
R570 B.n480 B.n59 163.367
R571 B.n480 B.n479 163.367
R572 B.n479 B.n478 163.367
R573 B.n478 B.n61 163.367
R574 B.n474 B.n61 163.367
R575 B.n474 B.n473 163.367
R576 B.n473 B.n472 163.367
R577 B.n472 B.n63 163.367
R578 B.n468 B.n63 163.367
R579 B.n468 B.n467 163.367
R580 B.n467 B.n466 163.367
R581 B.n466 B.n65 163.367
R582 B.n462 B.n65 163.367
R583 B.n462 B.n461 163.367
R584 B.n461 B.n460 163.367
R585 B.n460 B.n67 163.367
R586 B.n456 B.n67 163.367
R587 B.n456 B.n455 163.367
R588 B.n455 B.n454 163.367
R589 B.n454 B.n69 163.367
R590 B.n450 B.n69 163.367
R591 B.n450 B.n449 163.367
R592 B.n602 B.n15 163.367
R593 B.n606 B.n15 163.367
R594 B.n607 B.n606 163.367
R595 B.n608 B.n607 163.367
R596 B.n608 B.n13 163.367
R597 B.n612 B.n13 163.367
R598 B.n613 B.n612 163.367
R599 B.n614 B.n613 163.367
R600 B.n614 B.n11 163.367
R601 B.n618 B.n11 163.367
R602 B.n619 B.n618 163.367
R603 B.n620 B.n619 163.367
R604 B.n620 B.n9 163.367
R605 B.n624 B.n9 163.367
R606 B.n625 B.n624 163.367
R607 B.n626 B.n625 163.367
R608 B.n626 B.n7 163.367
R609 B.n630 B.n7 163.367
R610 B.n631 B.n630 163.367
R611 B.n632 B.n631 163.367
R612 B.n632 B.n5 163.367
R613 B.n636 B.n5 163.367
R614 B.n637 B.n636 163.367
R615 B.n638 B.n637 163.367
R616 B.n638 B.n3 163.367
R617 B.n642 B.n3 163.367
R618 B.n643 B.n642 163.367
R619 B.n165 B.n2 163.367
R620 B.n168 B.n165 163.367
R621 B.n169 B.n168 163.367
R622 B.n170 B.n169 163.367
R623 B.n170 B.n163 163.367
R624 B.n174 B.n163 163.367
R625 B.n175 B.n174 163.367
R626 B.n176 B.n175 163.367
R627 B.n176 B.n161 163.367
R628 B.n180 B.n161 163.367
R629 B.n181 B.n180 163.367
R630 B.n182 B.n181 163.367
R631 B.n182 B.n159 163.367
R632 B.n186 B.n159 163.367
R633 B.n187 B.n186 163.367
R634 B.n188 B.n187 163.367
R635 B.n188 B.n157 163.367
R636 B.n192 B.n157 163.367
R637 B.n193 B.n192 163.367
R638 B.n194 B.n193 163.367
R639 B.n194 B.n155 163.367
R640 B.n198 B.n155 163.367
R641 B.n199 B.n198 163.367
R642 B.n200 B.n199 163.367
R643 B.n200 B.n153 163.367
R644 B.n204 B.n153 163.367
R645 B.n205 B.n204 163.367
R646 B.n129 B.n128 67.2975
R647 B.n289 B.n288 67.2975
R648 B.n47 B.n46 67.2975
R649 B.n41 B.n40 67.2975
R650 B.n275 B.n129 59.5399
R651 B.n290 B.n289 59.5399
R652 B.n518 B.n47 59.5399
R653 B.n532 B.n41 59.5399
R654 B.n603 B.n16 33.2493
R655 B.n447 B.n70 33.2493
R656 B.n362 B.n361 33.2493
R657 B.n207 B.n152 33.2493
R658 B B.n645 18.0485
R659 B.n604 B.n603 10.6151
R660 B.n605 B.n604 10.6151
R661 B.n605 B.n14 10.6151
R662 B.n609 B.n14 10.6151
R663 B.n610 B.n609 10.6151
R664 B.n611 B.n610 10.6151
R665 B.n611 B.n12 10.6151
R666 B.n615 B.n12 10.6151
R667 B.n616 B.n615 10.6151
R668 B.n617 B.n616 10.6151
R669 B.n617 B.n10 10.6151
R670 B.n621 B.n10 10.6151
R671 B.n622 B.n621 10.6151
R672 B.n623 B.n622 10.6151
R673 B.n623 B.n8 10.6151
R674 B.n627 B.n8 10.6151
R675 B.n628 B.n627 10.6151
R676 B.n629 B.n628 10.6151
R677 B.n629 B.n6 10.6151
R678 B.n633 B.n6 10.6151
R679 B.n634 B.n633 10.6151
R680 B.n635 B.n634 10.6151
R681 B.n635 B.n4 10.6151
R682 B.n639 B.n4 10.6151
R683 B.n640 B.n639 10.6151
R684 B.n641 B.n640 10.6151
R685 B.n641 B.n0 10.6151
R686 B.n599 B.n16 10.6151
R687 B.n599 B.n598 10.6151
R688 B.n598 B.n597 10.6151
R689 B.n597 B.n18 10.6151
R690 B.n593 B.n18 10.6151
R691 B.n593 B.n592 10.6151
R692 B.n592 B.n591 10.6151
R693 B.n591 B.n20 10.6151
R694 B.n587 B.n20 10.6151
R695 B.n587 B.n586 10.6151
R696 B.n586 B.n585 10.6151
R697 B.n585 B.n22 10.6151
R698 B.n581 B.n22 10.6151
R699 B.n581 B.n580 10.6151
R700 B.n580 B.n579 10.6151
R701 B.n579 B.n24 10.6151
R702 B.n575 B.n24 10.6151
R703 B.n575 B.n574 10.6151
R704 B.n574 B.n573 10.6151
R705 B.n573 B.n26 10.6151
R706 B.n569 B.n26 10.6151
R707 B.n569 B.n568 10.6151
R708 B.n568 B.n567 10.6151
R709 B.n567 B.n28 10.6151
R710 B.n563 B.n28 10.6151
R711 B.n563 B.n562 10.6151
R712 B.n562 B.n561 10.6151
R713 B.n561 B.n30 10.6151
R714 B.n557 B.n30 10.6151
R715 B.n557 B.n556 10.6151
R716 B.n556 B.n555 10.6151
R717 B.n555 B.n32 10.6151
R718 B.n551 B.n32 10.6151
R719 B.n551 B.n550 10.6151
R720 B.n550 B.n549 10.6151
R721 B.n549 B.n34 10.6151
R722 B.n545 B.n34 10.6151
R723 B.n545 B.n544 10.6151
R724 B.n544 B.n543 10.6151
R725 B.n543 B.n36 10.6151
R726 B.n539 B.n36 10.6151
R727 B.n539 B.n538 10.6151
R728 B.n538 B.n537 10.6151
R729 B.n537 B.n38 10.6151
R730 B.n533 B.n38 10.6151
R731 B.n531 B.n530 10.6151
R732 B.n530 B.n42 10.6151
R733 B.n526 B.n42 10.6151
R734 B.n526 B.n525 10.6151
R735 B.n525 B.n524 10.6151
R736 B.n524 B.n44 10.6151
R737 B.n520 B.n44 10.6151
R738 B.n520 B.n519 10.6151
R739 B.n517 B.n48 10.6151
R740 B.n513 B.n48 10.6151
R741 B.n513 B.n512 10.6151
R742 B.n512 B.n511 10.6151
R743 B.n511 B.n50 10.6151
R744 B.n507 B.n50 10.6151
R745 B.n507 B.n506 10.6151
R746 B.n506 B.n505 10.6151
R747 B.n505 B.n52 10.6151
R748 B.n501 B.n52 10.6151
R749 B.n501 B.n500 10.6151
R750 B.n500 B.n499 10.6151
R751 B.n499 B.n54 10.6151
R752 B.n495 B.n54 10.6151
R753 B.n495 B.n494 10.6151
R754 B.n494 B.n493 10.6151
R755 B.n493 B.n56 10.6151
R756 B.n489 B.n56 10.6151
R757 B.n489 B.n488 10.6151
R758 B.n488 B.n487 10.6151
R759 B.n487 B.n58 10.6151
R760 B.n483 B.n58 10.6151
R761 B.n483 B.n482 10.6151
R762 B.n482 B.n481 10.6151
R763 B.n481 B.n60 10.6151
R764 B.n477 B.n60 10.6151
R765 B.n477 B.n476 10.6151
R766 B.n476 B.n475 10.6151
R767 B.n475 B.n62 10.6151
R768 B.n471 B.n62 10.6151
R769 B.n471 B.n470 10.6151
R770 B.n470 B.n469 10.6151
R771 B.n469 B.n64 10.6151
R772 B.n465 B.n64 10.6151
R773 B.n465 B.n464 10.6151
R774 B.n464 B.n463 10.6151
R775 B.n463 B.n66 10.6151
R776 B.n459 B.n66 10.6151
R777 B.n459 B.n458 10.6151
R778 B.n458 B.n457 10.6151
R779 B.n457 B.n68 10.6151
R780 B.n453 B.n68 10.6151
R781 B.n453 B.n452 10.6151
R782 B.n452 B.n451 10.6151
R783 B.n451 B.n70 10.6151
R784 B.n447 B.n446 10.6151
R785 B.n446 B.n445 10.6151
R786 B.n445 B.n72 10.6151
R787 B.n441 B.n72 10.6151
R788 B.n441 B.n440 10.6151
R789 B.n440 B.n439 10.6151
R790 B.n439 B.n74 10.6151
R791 B.n435 B.n74 10.6151
R792 B.n435 B.n434 10.6151
R793 B.n434 B.n433 10.6151
R794 B.n433 B.n76 10.6151
R795 B.n429 B.n76 10.6151
R796 B.n429 B.n428 10.6151
R797 B.n428 B.n427 10.6151
R798 B.n427 B.n78 10.6151
R799 B.n423 B.n78 10.6151
R800 B.n423 B.n422 10.6151
R801 B.n422 B.n421 10.6151
R802 B.n421 B.n80 10.6151
R803 B.n417 B.n80 10.6151
R804 B.n417 B.n416 10.6151
R805 B.n416 B.n415 10.6151
R806 B.n415 B.n82 10.6151
R807 B.n411 B.n82 10.6151
R808 B.n411 B.n410 10.6151
R809 B.n410 B.n409 10.6151
R810 B.n409 B.n84 10.6151
R811 B.n405 B.n84 10.6151
R812 B.n405 B.n404 10.6151
R813 B.n404 B.n403 10.6151
R814 B.n403 B.n86 10.6151
R815 B.n399 B.n86 10.6151
R816 B.n399 B.n398 10.6151
R817 B.n398 B.n397 10.6151
R818 B.n397 B.n88 10.6151
R819 B.n393 B.n88 10.6151
R820 B.n393 B.n392 10.6151
R821 B.n392 B.n391 10.6151
R822 B.n391 B.n90 10.6151
R823 B.n387 B.n90 10.6151
R824 B.n387 B.n386 10.6151
R825 B.n386 B.n385 10.6151
R826 B.n385 B.n92 10.6151
R827 B.n381 B.n92 10.6151
R828 B.n381 B.n380 10.6151
R829 B.n380 B.n379 10.6151
R830 B.n379 B.n94 10.6151
R831 B.n375 B.n94 10.6151
R832 B.n375 B.n374 10.6151
R833 B.n374 B.n373 10.6151
R834 B.n373 B.n96 10.6151
R835 B.n369 B.n96 10.6151
R836 B.n369 B.n368 10.6151
R837 B.n368 B.n367 10.6151
R838 B.n367 B.n98 10.6151
R839 B.n363 B.n98 10.6151
R840 B.n363 B.n362 10.6151
R841 B.n166 B.n1 10.6151
R842 B.n167 B.n166 10.6151
R843 B.n167 B.n164 10.6151
R844 B.n171 B.n164 10.6151
R845 B.n172 B.n171 10.6151
R846 B.n173 B.n172 10.6151
R847 B.n173 B.n162 10.6151
R848 B.n177 B.n162 10.6151
R849 B.n178 B.n177 10.6151
R850 B.n179 B.n178 10.6151
R851 B.n179 B.n160 10.6151
R852 B.n183 B.n160 10.6151
R853 B.n184 B.n183 10.6151
R854 B.n185 B.n184 10.6151
R855 B.n185 B.n158 10.6151
R856 B.n189 B.n158 10.6151
R857 B.n190 B.n189 10.6151
R858 B.n191 B.n190 10.6151
R859 B.n191 B.n156 10.6151
R860 B.n195 B.n156 10.6151
R861 B.n196 B.n195 10.6151
R862 B.n197 B.n196 10.6151
R863 B.n197 B.n154 10.6151
R864 B.n201 B.n154 10.6151
R865 B.n202 B.n201 10.6151
R866 B.n203 B.n202 10.6151
R867 B.n203 B.n152 10.6151
R868 B.n208 B.n207 10.6151
R869 B.n209 B.n208 10.6151
R870 B.n209 B.n150 10.6151
R871 B.n213 B.n150 10.6151
R872 B.n214 B.n213 10.6151
R873 B.n215 B.n214 10.6151
R874 B.n215 B.n148 10.6151
R875 B.n219 B.n148 10.6151
R876 B.n220 B.n219 10.6151
R877 B.n221 B.n220 10.6151
R878 B.n221 B.n146 10.6151
R879 B.n225 B.n146 10.6151
R880 B.n226 B.n225 10.6151
R881 B.n227 B.n226 10.6151
R882 B.n227 B.n144 10.6151
R883 B.n231 B.n144 10.6151
R884 B.n232 B.n231 10.6151
R885 B.n233 B.n232 10.6151
R886 B.n233 B.n142 10.6151
R887 B.n237 B.n142 10.6151
R888 B.n238 B.n237 10.6151
R889 B.n239 B.n238 10.6151
R890 B.n239 B.n140 10.6151
R891 B.n243 B.n140 10.6151
R892 B.n244 B.n243 10.6151
R893 B.n245 B.n244 10.6151
R894 B.n245 B.n138 10.6151
R895 B.n249 B.n138 10.6151
R896 B.n250 B.n249 10.6151
R897 B.n251 B.n250 10.6151
R898 B.n251 B.n136 10.6151
R899 B.n255 B.n136 10.6151
R900 B.n256 B.n255 10.6151
R901 B.n257 B.n256 10.6151
R902 B.n257 B.n134 10.6151
R903 B.n261 B.n134 10.6151
R904 B.n262 B.n261 10.6151
R905 B.n263 B.n262 10.6151
R906 B.n263 B.n132 10.6151
R907 B.n267 B.n132 10.6151
R908 B.n268 B.n267 10.6151
R909 B.n269 B.n268 10.6151
R910 B.n269 B.n130 10.6151
R911 B.n273 B.n130 10.6151
R912 B.n274 B.n273 10.6151
R913 B.n276 B.n126 10.6151
R914 B.n280 B.n126 10.6151
R915 B.n281 B.n280 10.6151
R916 B.n282 B.n281 10.6151
R917 B.n282 B.n124 10.6151
R918 B.n286 B.n124 10.6151
R919 B.n287 B.n286 10.6151
R920 B.n291 B.n287 10.6151
R921 B.n295 B.n122 10.6151
R922 B.n296 B.n295 10.6151
R923 B.n297 B.n296 10.6151
R924 B.n297 B.n120 10.6151
R925 B.n301 B.n120 10.6151
R926 B.n302 B.n301 10.6151
R927 B.n303 B.n302 10.6151
R928 B.n303 B.n118 10.6151
R929 B.n307 B.n118 10.6151
R930 B.n308 B.n307 10.6151
R931 B.n309 B.n308 10.6151
R932 B.n309 B.n116 10.6151
R933 B.n313 B.n116 10.6151
R934 B.n314 B.n313 10.6151
R935 B.n315 B.n314 10.6151
R936 B.n315 B.n114 10.6151
R937 B.n319 B.n114 10.6151
R938 B.n320 B.n319 10.6151
R939 B.n321 B.n320 10.6151
R940 B.n321 B.n112 10.6151
R941 B.n325 B.n112 10.6151
R942 B.n326 B.n325 10.6151
R943 B.n327 B.n326 10.6151
R944 B.n327 B.n110 10.6151
R945 B.n331 B.n110 10.6151
R946 B.n332 B.n331 10.6151
R947 B.n333 B.n332 10.6151
R948 B.n333 B.n108 10.6151
R949 B.n337 B.n108 10.6151
R950 B.n338 B.n337 10.6151
R951 B.n339 B.n338 10.6151
R952 B.n339 B.n106 10.6151
R953 B.n343 B.n106 10.6151
R954 B.n344 B.n343 10.6151
R955 B.n345 B.n344 10.6151
R956 B.n345 B.n104 10.6151
R957 B.n349 B.n104 10.6151
R958 B.n350 B.n349 10.6151
R959 B.n351 B.n350 10.6151
R960 B.n351 B.n102 10.6151
R961 B.n355 B.n102 10.6151
R962 B.n356 B.n355 10.6151
R963 B.n357 B.n356 10.6151
R964 B.n357 B.n100 10.6151
R965 B.n361 B.n100 10.6151
R966 B.n645 B.n0 8.11757
R967 B.n645 B.n1 8.11757
R968 B.n532 B.n531 6.5566
R969 B.n519 B.n518 6.5566
R970 B.n276 B.n275 6.5566
R971 B.n291 B.n290 6.5566
R972 B.n533 B.n532 4.05904
R973 B.n518 B.n517 4.05904
R974 B.n275 B.n274 4.05904
R975 B.n290 B.n122 4.05904
R976 VP.n0 VP.t1 188.869
R977 VP.n0 VP.t0 141.713
R978 VP VP.n0 0.52637
R979 VTAIL.n241 VTAIL.n240 585
R980 VTAIL.n243 VTAIL.n242 585
R981 VTAIL.n236 VTAIL.n235 585
R982 VTAIL.n249 VTAIL.n248 585
R983 VTAIL.n251 VTAIL.n250 585
R984 VTAIL.n232 VTAIL.n231 585
R985 VTAIL.n257 VTAIL.n256 585
R986 VTAIL.n259 VTAIL.n258 585
R987 VTAIL.n228 VTAIL.n227 585
R988 VTAIL.n265 VTAIL.n264 585
R989 VTAIL.n267 VTAIL.n266 585
R990 VTAIL.n224 VTAIL.n223 585
R991 VTAIL.n273 VTAIL.n272 585
R992 VTAIL.n275 VTAIL.n274 585
R993 VTAIL.n220 VTAIL.n219 585
R994 VTAIL.n281 VTAIL.n280 585
R995 VTAIL.n283 VTAIL.n282 585
R996 VTAIL.n25 VTAIL.n24 585
R997 VTAIL.n27 VTAIL.n26 585
R998 VTAIL.n20 VTAIL.n19 585
R999 VTAIL.n33 VTAIL.n32 585
R1000 VTAIL.n35 VTAIL.n34 585
R1001 VTAIL.n16 VTAIL.n15 585
R1002 VTAIL.n41 VTAIL.n40 585
R1003 VTAIL.n43 VTAIL.n42 585
R1004 VTAIL.n12 VTAIL.n11 585
R1005 VTAIL.n49 VTAIL.n48 585
R1006 VTAIL.n51 VTAIL.n50 585
R1007 VTAIL.n8 VTAIL.n7 585
R1008 VTAIL.n57 VTAIL.n56 585
R1009 VTAIL.n59 VTAIL.n58 585
R1010 VTAIL.n4 VTAIL.n3 585
R1011 VTAIL.n65 VTAIL.n64 585
R1012 VTAIL.n67 VTAIL.n66 585
R1013 VTAIL.n211 VTAIL.n210 585
R1014 VTAIL.n209 VTAIL.n208 585
R1015 VTAIL.n148 VTAIL.n147 585
R1016 VTAIL.n203 VTAIL.n202 585
R1017 VTAIL.n201 VTAIL.n200 585
R1018 VTAIL.n152 VTAIL.n151 585
R1019 VTAIL.n195 VTAIL.n194 585
R1020 VTAIL.n193 VTAIL.n192 585
R1021 VTAIL.n156 VTAIL.n155 585
R1022 VTAIL.n187 VTAIL.n186 585
R1023 VTAIL.n185 VTAIL.n184 585
R1024 VTAIL.n160 VTAIL.n159 585
R1025 VTAIL.n179 VTAIL.n178 585
R1026 VTAIL.n177 VTAIL.n176 585
R1027 VTAIL.n164 VTAIL.n163 585
R1028 VTAIL.n171 VTAIL.n170 585
R1029 VTAIL.n169 VTAIL.n168 585
R1030 VTAIL.n139 VTAIL.n138 585
R1031 VTAIL.n137 VTAIL.n136 585
R1032 VTAIL.n76 VTAIL.n75 585
R1033 VTAIL.n131 VTAIL.n130 585
R1034 VTAIL.n129 VTAIL.n128 585
R1035 VTAIL.n80 VTAIL.n79 585
R1036 VTAIL.n123 VTAIL.n122 585
R1037 VTAIL.n121 VTAIL.n120 585
R1038 VTAIL.n84 VTAIL.n83 585
R1039 VTAIL.n115 VTAIL.n114 585
R1040 VTAIL.n113 VTAIL.n112 585
R1041 VTAIL.n88 VTAIL.n87 585
R1042 VTAIL.n107 VTAIL.n106 585
R1043 VTAIL.n105 VTAIL.n104 585
R1044 VTAIL.n92 VTAIL.n91 585
R1045 VTAIL.n99 VTAIL.n98 585
R1046 VTAIL.n97 VTAIL.n96 585
R1047 VTAIL.n282 VTAIL.n216 498.474
R1048 VTAIL.n66 VTAIL.n0 498.474
R1049 VTAIL.n210 VTAIL.n144 498.474
R1050 VTAIL.n138 VTAIL.n72 498.474
R1051 VTAIL.n239 VTAIL.t1 327.466
R1052 VTAIL.n23 VTAIL.t2 327.466
R1053 VTAIL.n167 VTAIL.t3 327.466
R1054 VTAIL.n95 VTAIL.t0 327.466
R1055 VTAIL.n242 VTAIL.n241 171.744
R1056 VTAIL.n242 VTAIL.n235 171.744
R1057 VTAIL.n249 VTAIL.n235 171.744
R1058 VTAIL.n250 VTAIL.n249 171.744
R1059 VTAIL.n250 VTAIL.n231 171.744
R1060 VTAIL.n257 VTAIL.n231 171.744
R1061 VTAIL.n258 VTAIL.n257 171.744
R1062 VTAIL.n258 VTAIL.n227 171.744
R1063 VTAIL.n265 VTAIL.n227 171.744
R1064 VTAIL.n266 VTAIL.n265 171.744
R1065 VTAIL.n266 VTAIL.n223 171.744
R1066 VTAIL.n273 VTAIL.n223 171.744
R1067 VTAIL.n274 VTAIL.n273 171.744
R1068 VTAIL.n274 VTAIL.n219 171.744
R1069 VTAIL.n281 VTAIL.n219 171.744
R1070 VTAIL.n282 VTAIL.n281 171.744
R1071 VTAIL.n26 VTAIL.n25 171.744
R1072 VTAIL.n26 VTAIL.n19 171.744
R1073 VTAIL.n33 VTAIL.n19 171.744
R1074 VTAIL.n34 VTAIL.n33 171.744
R1075 VTAIL.n34 VTAIL.n15 171.744
R1076 VTAIL.n41 VTAIL.n15 171.744
R1077 VTAIL.n42 VTAIL.n41 171.744
R1078 VTAIL.n42 VTAIL.n11 171.744
R1079 VTAIL.n49 VTAIL.n11 171.744
R1080 VTAIL.n50 VTAIL.n49 171.744
R1081 VTAIL.n50 VTAIL.n7 171.744
R1082 VTAIL.n57 VTAIL.n7 171.744
R1083 VTAIL.n58 VTAIL.n57 171.744
R1084 VTAIL.n58 VTAIL.n3 171.744
R1085 VTAIL.n65 VTAIL.n3 171.744
R1086 VTAIL.n66 VTAIL.n65 171.744
R1087 VTAIL.n210 VTAIL.n209 171.744
R1088 VTAIL.n209 VTAIL.n147 171.744
R1089 VTAIL.n202 VTAIL.n147 171.744
R1090 VTAIL.n202 VTAIL.n201 171.744
R1091 VTAIL.n201 VTAIL.n151 171.744
R1092 VTAIL.n194 VTAIL.n151 171.744
R1093 VTAIL.n194 VTAIL.n193 171.744
R1094 VTAIL.n193 VTAIL.n155 171.744
R1095 VTAIL.n186 VTAIL.n155 171.744
R1096 VTAIL.n186 VTAIL.n185 171.744
R1097 VTAIL.n185 VTAIL.n159 171.744
R1098 VTAIL.n178 VTAIL.n159 171.744
R1099 VTAIL.n178 VTAIL.n177 171.744
R1100 VTAIL.n177 VTAIL.n163 171.744
R1101 VTAIL.n170 VTAIL.n163 171.744
R1102 VTAIL.n170 VTAIL.n169 171.744
R1103 VTAIL.n138 VTAIL.n137 171.744
R1104 VTAIL.n137 VTAIL.n75 171.744
R1105 VTAIL.n130 VTAIL.n75 171.744
R1106 VTAIL.n130 VTAIL.n129 171.744
R1107 VTAIL.n129 VTAIL.n79 171.744
R1108 VTAIL.n122 VTAIL.n79 171.744
R1109 VTAIL.n122 VTAIL.n121 171.744
R1110 VTAIL.n121 VTAIL.n83 171.744
R1111 VTAIL.n114 VTAIL.n83 171.744
R1112 VTAIL.n114 VTAIL.n113 171.744
R1113 VTAIL.n113 VTAIL.n87 171.744
R1114 VTAIL.n106 VTAIL.n87 171.744
R1115 VTAIL.n106 VTAIL.n105 171.744
R1116 VTAIL.n105 VTAIL.n91 171.744
R1117 VTAIL.n98 VTAIL.n91 171.744
R1118 VTAIL.n98 VTAIL.n97 171.744
R1119 VTAIL.n241 VTAIL.t1 85.8723
R1120 VTAIL.n25 VTAIL.t2 85.8723
R1121 VTAIL.n169 VTAIL.t3 85.8723
R1122 VTAIL.n97 VTAIL.t0 85.8723
R1123 VTAIL.n287 VTAIL.n286 36.2581
R1124 VTAIL.n71 VTAIL.n70 36.2581
R1125 VTAIL.n215 VTAIL.n214 36.2581
R1126 VTAIL.n143 VTAIL.n142 36.2581
R1127 VTAIL.n143 VTAIL.n71 29.91
R1128 VTAIL.n287 VTAIL.n215 26.9186
R1129 VTAIL.n240 VTAIL.n239 16.3895
R1130 VTAIL.n24 VTAIL.n23 16.3895
R1131 VTAIL.n168 VTAIL.n167 16.3895
R1132 VTAIL.n96 VTAIL.n95 16.3895
R1133 VTAIL.n243 VTAIL.n238 12.8005
R1134 VTAIL.n284 VTAIL.n283 12.8005
R1135 VTAIL.n27 VTAIL.n22 12.8005
R1136 VTAIL.n68 VTAIL.n67 12.8005
R1137 VTAIL.n212 VTAIL.n211 12.8005
R1138 VTAIL.n171 VTAIL.n166 12.8005
R1139 VTAIL.n140 VTAIL.n139 12.8005
R1140 VTAIL.n99 VTAIL.n94 12.8005
R1141 VTAIL.n244 VTAIL.n236 12.0247
R1142 VTAIL.n280 VTAIL.n218 12.0247
R1143 VTAIL.n28 VTAIL.n20 12.0247
R1144 VTAIL.n64 VTAIL.n2 12.0247
R1145 VTAIL.n208 VTAIL.n146 12.0247
R1146 VTAIL.n172 VTAIL.n164 12.0247
R1147 VTAIL.n136 VTAIL.n74 12.0247
R1148 VTAIL.n100 VTAIL.n92 12.0247
R1149 VTAIL.n248 VTAIL.n247 11.249
R1150 VTAIL.n279 VTAIL.n220 11.249
R1151 VTAIL.n32 VTAIL.n31 11.249
R1152 VTAIL.n63 VTAIL.n4 11.249
R1153 VTAIL.n207 VTAIL.n148 11.249
R1154 VTAIL.n176 VTAIL.n175 11.249
R1155 VTAIL.n135 VTAIL.n76 11.249
R1156 VTAIL.n104 VTAIL.n103 11.249
R1157 VTAIL.n251 VTAIL.n234 10.4732
R1158 VTAIL.n276 VTAIL.n275 10.4732
R1159 VTAIL.n35 VTAIL.n18 10.4732
R1160 VTAIL.n60 VTAIL.n59 10.4732
R1161 VTAIL.n204 VTAIL.n203 10.4732
R1162 VTAIL.n179 VTAIL.n162 10.4732
R1163 VTAIL.n132 VTAIL.n131 10.4732
R1164 VTAIL.n107 VTAIL.n90 10.4732
R1165 VTAIL.n252 VTAIL.n232 9.69747
R1166 VTAIL.n272 VTAIL.n222 9.69747
R1167 VTAIL.n36 VTAIL.n16 9.69747
R1168 VTAIL.n56 VTAIL.n6 9.69747
R1169 VTAIL.n200 VTAIL.n150 9.69747
R1170 VTAIL.n180 VTAIL.n160 9.69747
R1171 VTAIL.n128 VTAIL.n78 9.69747
R1172 VTAIL.n108 VTAIL.n88 9.69747
R1173 VTAIL.n286 VTAIL.n285 9.45567
R1174 VTAIL.n70 VTAIL.n69 9.45567
R1175 VTAIL.n214 VTAIL.n213 9.45567
R1176 VTAIL.n142 VTAIL.n141 9.45567
R1177 VTAIL.n261 VTAIL.n260 9.3005
R1178 VTAIL.n230 VTAIL.n229 9.3005
R1179 VTAIL.n255 VTAIL.n254 9.3005
R1180 VTAIL.n253 VTAIL.n252 9.3005
R1181 VTAIL.n234 VTAIL.n233 9.3005
R1182 VTAIL.n247 VTAIL.n246 9.3005
R1183 VTAIL.n245 VTAIL.n244 9.3005
R1184 VTAIL.n238 VTAIL.n237 9.3005
R1185 VTAIL.n263 VTAIL.n262 9.3005
R1186 VTAIL.n226 VTAIL.n225 9.3005
R1187 VTAIL.n269 VTAIL.n268 9.3005
R1188 VTAIL.n271 VTAIL.n270 9.3005
R1189 VTAIL.n222 VTAIL.n221 9.3005
R1190 VTAIL.n277 VTAIL.n276 9.3005
R1191 VTAIL.n279 VTAIL.n278 9.3005
R1192 VTAIL.n218 VTAIL.n217 9.3005
R1193 VTAIL.n285 VTAIL.n284 9.3005
R1194 VTAIL.n45 VTAIL.n44 9.3005
R1195 VTAIL.n14 VTAIL.n13 9.3005
R1196 VTAIL.n39 VTAIL.n38 9.3005
R1197 VTAIL.n37 VTAIL.n36 9.3005
R1198 VTAIL.n18 VTAIL.n17 9.3005
R1199 VTAIL.n31 VTAIL.n30 9.3005
R1200 VTAIL.n29 VTAIL.n28 9.3005
R1201 VTAIL.n22 VTAIL.n21 9.3005
R1202 VTAIL.n47 VTAIL.n46 9.3005
R1203 VTAIL.n10 VTAIL.n9 9.3005
R1204 VTAIL.n53 VTAIL.n52 9.3005
R1205 VTAIL.n55 VTAIL.n54 9.3005
R1206 VTAIL.n6 VTAIL.n5 9.3005
R1207 VTAIL.n61 VTAIL.n60 9.3005
R1208 VTAIL.n63 VTAIL.n62 9.3005
R1209 VTAIL.n2 VTAIL.n1 9.3005
R1210 VTAIL.n69 VTAIL.n68 9.3005
R1211 VTAIL.n154 VTAIL.n153 9.3005
R1212 VTAIL.n197 VTAIL.n196 9.3005
R1213 VTAIL.n199 VTAIL.n198 9.3005
R1214 VTAIL.n150 VTAIL.n149 9.3005
R1215 VTAIL.n205 VTAIL.n204 9.3005
R1216 VTAIL.n207 VTAIL.n206 9.3005
R1217 VTAIL.n146 VTAIL.n145 9.3005
R1218 VTAIL.n213 VTAIL.n212 9.3005
R1219 VTAIL.n191 VTAIL.n190 9.3005
R1220 VTAIL.n189 VTAIL.n188 9.3005
R1221 VTAIL.n158 VTAIL.n157 9.3005
R1222 VTAIL.n183 VTAIL.n182 9.3005
R1223 VTAIL.n181 VTAIL.n180 9.3005
R1224 VTAIL.n162 VTAIL.n161 9.3005
R1225 VTAIL.n175 VTAIL.n174 9.3005
R1226 VTAIL.n173 VTAIL.n172 9.3005
R1227 VTAIL.n166 VTAIL.n165 9.3005
R1228 VTAIL.n82 VTAIL.n81 9.3005
R1229 VTAIL.n125 VTAIL.n124 9.3005
R1230 VTAIL.n127 VTAIL.n126 9.3005
R1231 VTAIL.n78 VTAIL.n77 9.3005
R1232 VTAIL.n133 VTAIL.n132 9.3005
R1233 VTAIL.n135 VTAIL.n134 9.3005
R1234 VTAIL.n74 VTAIL.n73 9.3005
R1235 VTAIL.n141 VTAIL.n140 9.3005
R1236 VTAIL.n119 VTAIL.n118 9.3005
R1237 VTAIL.n117 VTAIL.n116 9.3005
R1238 VTAIL.n86 VTAIL.n85 9.3005
R1239 VTAIL.n111 VTAIL.n110 9.3005
R1240 VTAIL.n109 VTAIL.n108 9.3005
R1241 VTAIL.n90 VTAIL.n89 9.3005
R1242 VTAIL.n103 VTAIL.n102 9.3005
R1243 VTAIL.n101 VTAIL.n100 9.3005
R1244 VTAIL.n94 VTAIL.n93 9.3005
R1245 VTAIL.n256 VTAIL.n255 8.92171
R1246 VTAIL.n271 VTAIL.n224 8.92171
R1247 VTAIL.n40 VTAIL.n39 8.92171
R1248 VTAIL.n55 VTAIL.n8 8.92171
R1249 VTAIL.n199 VTAIL.n152 8.92171
R1250 VTAIL.n184 VTAIL.n183 8.92171
R1251 VTAIL.n127 VTAIL.n80 8.92171
R1252 VTAIL.n112 VTAIL.n111 8.92171
R1253 VTAIL.n259 VTAIL.n230 8.14595
R1254 VTAIL.n268 VTAIL.n267 8.14595
R1255 VTAIL.n43 VTAIL.n14 8.14595
R1256 VTAIL.n52 VTAIL.n51 8.14595
R1257 VTAIL.n196 VTAIL.n195 8.14595
R1258 VTAIL.n187 VTAIL.n158 8.14595
R1259 VTAIL.n124 VTAIL.n123 8.14595
R1260 VTAIL.n115 VTAIL.n86 8.14595
R1261 VTAIL.n286 VTAIL.n216 7.75445
R1262 VTAIL.n70 VTAIL.n0 7.75445
R1263 VTAIL.n214 VTAIL.n144 7.75445
R1264 VTAIL.n142 VTAIL.n72 7.75445
R1265 VTAIL.n260 VTAIL.n228 7.3702
R1266 VTAIL.n264 VTAIL.n226 7.3702
R1267 VTAIL.n44 VTAIL.n12 7.3702
R1268 VTAIL.n48 VTAIL.n10 7.3702
R1269 VTAIL.n192 VTAIL.n154 7.3702
R1270 VTAIL.n188 VTAIL.n156 7.3702
R1271 VTAIL.n120 VTAIL.n82 7.3702
R1272 VTAIL.n116 VTAIL.n84 7.3702
R1273 VTAIL.n263 VTAIL.n228 6.59444
R1274 VTAIL.n264 VTAIL.n263 6.59444
R1275 VTAIL.n47 VTAIL.n12 6.59444
R1276 VTAIL.n48 VTAIL.n47 6.59444
R1277 VTAIL.n192 VTAIL.n191 6.59444
R1278 VTAIL.n191 VTAIL.n156 6.59444
R1279 VTAIL.n120 VTAIL.n119 6.59444
R1280 VTAIL.n119 VTAIL.n84 6.59444
R1281 VTAIL.n284 VTAIL.n216 6.08283
R1282 VTAIL.n68 VTAIL.n0 6.08283
R1283 VTAIL.n212 VTAIL.n144 6.08283
R1284 VTAIL.n140 VTAIL.n72 6.08283
R1285 VTAIL.n260 VTAIL.n259 5.81868
R1286 VTAIL.n267 VTAIL.n226 5.81868
R1287 VTAIL.n44 VTAIL.n43 5.81868
R1288 VTAIL.n51 VTAIL.n10 5.81868
R1289 VTAIL.n195 VTAIL.n154 5.81868
R1290 VTAIL.n188 VTAIL.n187 5.81868
R1291 VTAIL.n123 VTAIL.n82 5.81868
R1292 VTAIL.n116 VTAIL.n115 5.81868
R1293 VTAIL.n256 VTAIL.n230 5.04292
R1294 VTAIL.n268 VTAIL.n224 5.04292
R1295 VTAIL.n40 VTAIL.n14 5.04292
R1296 VTAIL.n52 VTAIL.n8 5.04292
R1297 VTAIL.n196 VTAIL.n152 5.04292
R1298 VTAIL.n184 VTAIL.n158 5.04292
R1299 VTAIL.n124 VTAIL.n80 5.04292
R1300 VTAIL.n112 VTAIL.n86 5.04292
R1301 VTAIL.n255 VTAIL.n232 4.26717
R1302 VTAIL.n272 VTAIL.n271 4.26717
R1303 VTAIL.n39 VTAIL.n16 4.26717
R1304 VTAIL.n56 VTAIL.n55 4.26717
R1305 VTAIL.n200 VTAIL.n199 4.26717
R1306 VTAIL.n183 VTAIL.n160 4.26717
R1307 VTAIL.n128 VTAIL.n127 4.26717
R1308 VTAIL.n111 VTAIL.n88 4.26717
R1309 VTAIL.n239 VTAIL.n237 3.70982
R1310 VTAIL.n23 VTAIL.n21 3.70982
R1311 VTAIL.n167 VTAIL.n165 3.70982
R1312 VTAIL.n95 VTAIL.n93 3.70982
R1313 VTAIL.n252 VTAIL.n251 3.49141
R1314 VTAIL.n275 VTAIL.n222 3.49141
R1315 VTAIL.n36 VTAIL.n35 3.49141
R1316 VTAIL.n59 VTAIL.n6 3.49141
R1317 VTAIL.n203 VTAIL.n150 3.49141
R1318 VTAIL.n180 VTAIL.n179 3.49141
R1319 VTAIL.n131 VTAIL.n78 3.49141
R1320 VTAIL.n108 VTAIL.n107 3.49141
R1321 VTAIL.n248 VTAIL.n234 2.71565
R1322 VTAIL.n276 VTAIL.n220 2.71565
R1323 VTAIL.n32 VTAIL.n18 2.71565
R1324 VTAIL.n60 VTAIL.n4 2.71565
R1325 VTAIL.n204 VTAIL.n148 2.71565
R1326 VTAIL.n176 VTAIL.n162 2.71565
R1327 VTAIL.n132 VTAIL.n76 2.71565
R1328 VTAIL.n104 VTAIL.n90 2.71565
R1329 VTAIL.n215 VTAIL.n143 1.96602
R1330 VTAIL.n247 VTAIL.n236 1.93989
R1331 VTAIL.n280 VTAIL.n279 1.93989
R1332 VTAIL.n31 VTAIL.n20 1.93989
R1333 VTAIL.n64 VTAIL.n63 1.93989
R1334 VTAIL.n208 VTAIL.n207 1.93989
R1335 VTAIL.n175 VTAIL.n164 1.93989
R1336 VTAIL.n136 VTAIL.n135 1.93989
R1337 VTAIL.n103 VTAIL.n92 1.93989
R1338 VTAIL VTAIL.n71 1.27636
R1339 VTAIL.n244 VTAIL.n243 1.16414
R1340 VTAIL.n283 VTAIL.n218 1.16414
R1341 VTAIL.n28 VTAIL.n27 1.16414
R1342 VTAIL.n67 VTAIL.n2 1.16414
R1343 VTAIL.n211 VTAIL.n146 1.16414
R1344 VTAIL.n172 VTAIL.n171 1.16414
R1345 VTAIL.n139 VTAIL.n74 1.16414
R1346 VTAIL.n100 VTAIL.n99 1.16414
R1347 VTAIL VTAIL.n287 0.690155
R1348 VTAIL.n240 VTAIL.n238 0.388379
R1349 VTAIL.n24 VTAIL.n22 0.388379
R1350 VTAIL.n168 VTAIL.n166 0.388379
R1351 VTAIL.n96 VTAIL.n94 0.388379
R1352 VTAIL.n245 VTAIL.n237 0.155672
R1353 VTAIL.n246 VTAIL.n245 0.155672
R1354 VTAIL.n246 VTAIL.n233 0.155672
R1355 VTAIL.n253 VTAIL.n233 0.155672
R1356 VTAIL.n254 VTAIL.n253 0.155672
R1357 VTAIL.n254 VTAIL.n229 0.155672
R1358 VTAIL.n261 VTAIL.n229 0.155672
R1359 VTAIL.n262 VTAIL.n261 0.155672
R1360 VTAIL.n262 VTAIL.n225 0.155672
R1361 VTAIL.n269 VTAIL.n225 0.155672
R1362 VTAIL.n270 VTAIL.n269 0.155672
R1363 VTAIL.n270 VTAIL.n221 0.155672
R1364 VTAIL.n277 VTAIL.n221 0.155672
R1365 VTAIL.n278 VTAIL.n277 0.155672
R1366 VTAIL.n278 VTAIL.n217 0.155672
R1367 VTAIL.n285 VTAIL.n217 0.155672
R1368 VTAIL.n29 VTAIL.n21 0.155672
R1369 VTAIL.n30 VTAIL.n29 0.155672
R1370 VTAIL.n30 VTAIL.n17 0.155672
R1371 VTAIL.n37 VTAIL.n17 0.155672
R1372 VTAIL.n38 VTAIL.n37 0.155672
R1373 VTAIL.n38 VTAIL.n13 0.155672
R1374 VTAIL.n45 VTAIL.n13 0.155672
R1375 VTAIL.n46 VTAIL.n45 0.155672
R1376 VTAIL.n46 VTAIL.n9 0.155672
R1377 VTAIL.n53 VTAIL.n9 0.155672
R1378 VTAIL.n54 VTAIL.n53 0.155672
R1379 VTAIL.n54 VTAIL.n5 0.155672
R1380 VTAIL.n61 VTAIL.n5 0.155672
R1381 VTAIL.n62 VTAIL.n61 0.155672
R1382 VTAIL.n62 VTAIL.n1 0.155672
R1383 VTAIL.n69 VTAIL.n1 0.155672
R1384 VTAIL.n213 VTAIL.n145 0.155672
R1385 VTAIL.n206 VTAIL.n145 0.155672
R1386 VTAIL.n206 VTAIL.n205 0.155672
R1387 VTAIL.n205 VTAIL.n149 0.155672
R1388 VTAIL.n198 VTAIL.n149 0.155672
R1389 VTAIL.n198 VTAIL.n197 0.155672
R1390 VTAIL.n197 VTAIL.n153 0.155672
R1391 VTAIL.n190 VTAIL.n153 0.155672
R1392 VTAIL.n190 VTAIL.n189 0.155672
R1393 VTAIL.n189 VTAIL.n157 0.155672
R1394 VTAIL.n182 VTAIL.n157 0.155672
R1395 VTAIL.n182 VTAIL.n181 0.155672
R1396 VTAIL.n181 VTAIL.n161 0.155672
R1397 VTAIL.n174 VTAIL.n161 0.155672
R1398 VTAIL.n174 VTAIL.n173 0.155672
R1399 VTAIL.n173 VTAIL.n165 0.155672
R1400 VTAIL.n141 VTAIL.n73 0.155672
R1401 VTAIL.n134 VTAIL.n73 0.155672
R1402 VTAIL.n134 VTAIL.n133 0.155672
R1403 VTAIL.n133 VTAIL.n77 0.155672
R1404 VTAIL.n126 VTAIL.n77 0.155672
R1405 VTAIL.n126 VTAIL.n125 0.155672
R1406 VTAIL.n125 VTAIL.n81 0.155672
R1407 VTAIL.n118 VTAIL.n81 0.155672
R1408 VTAIL.n118 VTAIL.n117 0.155672
R1409 VTAIL.n117 VTAIL.n85 0.155672
R1410 VTAIL.n110 VTAIL.n85 0.155672
R1411 VTAIL.n110 VTAIL.n109 0.155672
R1412 VTAIL.n109 VTAIL.n89 0.155672
R1413 VTAIL.n102 VTAIL.n89 0.155672
R1414 VTAIL.n102 VTAIL.n101 0.155672
R1415 VTAIL.n101 VTAIL.n93 0.155672
R1416 VDD1.n67 VDD1.n66 585
R1417 VDD1.n65 VDD1.n64 585
R1418 VDD1.n4 VDD1.n3 585
R1419 VDD1.n59 VDD1.n58 585
R1420 VDD1.n57 VDD1.n56 585
R1421 VDD1.n8 VDD1.n7 585
R1422 VDD1.n51 VDD1.n50 585
R1423 VDD1.n49 VDD1.n48 585
R1424 VDD1.n12 VDD1.n11 585
R1425 VDD1.n43 VDD1.n42 585
R1426 VDD1.n41 VDD1.n40 585
R1427 VDD1.n16 VDD1.n15 585
R1428 VDD1.n35 VDD1.n34 585
R1429 VDD1.n33 VDD1.n32 585
R1430 VDD1.n20 VDD1.n19 585
R1431 VDD1.n27 VDD1.n26 585
R1432 VDD1.n25 VDD1.n24 585
R1433 VDD1.n96 VDD1.n95 585
R1434 VDD1.n98 VDD1.n97 585
R1435 VDD1.n91 VDD1.n90 585
R1436 VDD1.n104 VDD1.n103 585
R1437 VDD1.n106 VDD1.n105 585
R1438 VDD1.n87 VDD1.n86 585
R1439 VDD1.n112 VDD1.n111 585
R1440 VDD1.n114 VDD1.n113 585
R1441 VDD1.n83 VDD1.n82 585
R1442 VDD1.n120 VDD1.n119 585
R1443 VDD1.n122 VDD1.n121 585
R1444 VDD1.n79 VDD1.n78 585
R1445 VDD1.n128 VDD1.n127 585
R1446 VDD1.n130 VDD1.n129 585
R1447 VDD1.n75 VDD1.n74 585
R1448 VDD1.n136 VDD1.n135 585
R1449 VDD1.n138 VDD1.n137 585
R1450 VDD1.n66 VDD1.n0 498.474
R1451 VDD1.n137 VDD1.n71 498.474
R1452 VDD1.n23 VDD1.t0 327.466
R1453 VDD1.n94 VDD1.t1 327.466
R1454 VDD1.n66 VDD1.n65 171.744
R1455 VDD1.n65 VDD1.n3 171.744
R1456 VDD1.n58 VDD1.n3 171.744
R1457 VDD1.n58 VDD1.n57 171.744
R1458 VDD1.n57 VDD1.n7 171.744
R1459 VDD1.n50 VDD1.n7 171.744
R1460 VDD1.n50 VDD1.n49 171.744
R1461 VDD1.n49 VDD1.n11 171.744
R1462 VDD1.n42 VDD1.n11 171.744
R1463 VDD1.n42 VDD1.n41 171.744
R1464 VDD1.n41 VDD1.n15 171.744
R1465 VDD1.n34 VDD1.n15 171.744
R1466 VDD1.n34 VDD1.n33 171.744
R1467 VDD1.n33 VDD1.n19 171.744
R1468 VDD1.n26 VDD1.n19 171.744
R1469 VDD1.n26 VDD1.n25 171.744
R1470 VDD1.n97 VDD1.n96 171.744
R1471 VDD1.n97 VDD1.n90 171.744
R1472 VDD1.n104 VDD1.n90 171.744
R1473 VDD1.n105 VDD1.n104 171.744
R1474 VDD1.n105 VDD1.n86 171.744
R1475 VDD1.n112 VDD1.n86 171.744
R1476 VDD1.n113 VDD1.n112 171.744
R1477 VDD1.n113 VDD1.n82 171.744
R1478 VDD1.n120 VDD1.n82 171.744
R1479 VDD1.n121 VDD1.n120 171.744
R1480 VDD1.n121 VDD1.n78 171.744
R1481 VDD1.n128 VDD1.n78 171.744
R1482 VDD1.n129 VDD1.n128 171.744
R1483 VDD1.n129 VDD1.n74 171.744
R1484 VDD1.n136 VDD1.n74 171.744
R1485 VDD1.n137 VDD1.n136 171.744
R1486 VDD1 VDD1.n141 95.4121
R1487 VDD1.n25 VDD1.t0 85.8723
R1488 VDD1.n96 VDD1.t1 85.8723
R1489 VDD1 VDD1.n70 53.7429
R1490 VDD1.n24 VDD1.n23 16.3895
R1491 VDD1.n95 VDD1.n94 16.3895
R1492 VDD1.n68 VDD1.n67 12.8005
R1493 VDD1.n27 VDD1.n22 12.8005
R1494 VDD1.n98 VDD1.n93 12.8005
R1495 VDD1.n139 VDD1.n138 12.8005
R1496 VDD1.n64 VDD1.n2 12.0247
R1497 VDD1.n28 VDD1.n20 12.0247
R1498 VDD1.n99 VDD1.n91 12.0247
R1499 VDD1.n135 VDD1.n73 12.0247
R1500 VDD1.n63 VDD1.n4 11.249
R1501 VDD1.n32 VDD1.n31 11.249
R1502 VDD1.n103 VDD1.n102 11.249
R1503 VDD1.n134 VDD1.n75 11.249
R1504 VDD1.n60 VDD1.n59 10.4732
R1505 VDD1.n35 VDD1.n18 10.4732
R1506 VDD1.n106 VDD1.n89 10.4732
R1507 VDD1.n131 VDD1.n130 10.4732
R1508 VDD1.n56 VDD1.n6 9.69747
R1509 VDD1.n36 VDD1.n16 9.69747
R1510 VDD1.n107 VDD1.n87 9.69747
R1511 VDD1.n127 VDD1.n77 9.69747
R1512 VDD1.n70 VDD1.n69 9.45567
R1513 VDD1.n141 VDD1.n140 9.45567
R1514 VDD1.n10 VDD1.n9 9.3005
R1515 VDD1.n53 VDD1.n52 9.3005
R1516 VDD1.n55 VDD1.n54 9.3005
R1517 VDD1.n6 VDD1.n5 9.3005
R1518 VDD1.n61 VDD1.n60 9.3005
R1519 VDD1.n63 VDD1.n62 9.3005
R1520 VDD1.n2 VDD1.n1 9.3005
R1521 VDD1.n69 VDD1.n68 9.3005
R1522 VDD1.n47 VDD1.n46 9.3005
R1523 VDD1.n45 VDD1.n44 9.3005
R1524 VDD1.n14 VDD1.n13 9.3005
R1525 VDD1.n39 VDD1.n38 9.3005
R1526 VDD1.n37 VDD1.n36 9.3005
R1527 VDD1.n18 VDD1.n17 9.3005
R1528 VDD1.n31 VDD1.n30 9.3005
R1529 VDD1.n29 VDD1.n28 9.3005
R1530 VDD1.n22 VDD1.n21 9.3005
R1531 VDD1.n116 VDD1.n115 9.3005
R1532 VDD1.n85 VDD1.n84 9.3005
R1533 VDD1.n110 VDD1.n109 9.3005
R1534 VDD1.n108 VDD1.n107 9.3005
R1535 VDD1.n89 VDD1.n88 9.3005
R1536 VDD1.n102 VDD1.n101 9.3005
R1537 VDD1.n100 VDD1.n99 9.3005
R1538 VDD1.n93 VDD1.n92 9.3005
R1539 VDD1.n118 VDD1.n117 9.3005
R1540 VDD1.n81 VDD1.n80 9.3005
R1541 VDD1.n124 VDD1.n123 9.3005
R1542 VDD1.n126 VDD1.n125 9.3005
R1543 VDD1.n77 VDD1.n76 9.3005
R1544 VDD1.n132 VDD1.n131 9.3005
R1545 VDD1.n134 VDD1.n133 9.3005
R1546 VDD1.n73 VDD1.n72 9.3005
R1547 VDD1.n140 VDD1.n139 9.3005
R1548 VDD1.n55 VDD1.n8 8.92171
R1549 VDD1.n40 VDD1.n39 8.92171
R1550 VDD1.n111 VDD1.n110 8.92171
R1551 VDD1.n126 VDD1.n79 8.92171
R1552 VDD1.n52 VDD1.n51 8.14595
R1553 VDD1.n43 VDD1.n14 8.14595
R1554 VDD1.n114 VDD1.n85 8.14595
R1555 VDD1.n123 VDD1.n122 8.14595
R1556 VDD1.n70 VDD1.n0 7.75445
R1557 VDD1.n141 VDD1.n71 7.75445
R1558 VDD1.n48 VDD1.n10 7.3702
R1559 VDD1.n44 VDD1.n12 7.3702
R1560 VDD1.n115 VDD1.n83 7.3702
R1561 VDD1.n119 VDD1.n81 7.3702
R1562 VDD1.n48 VDD1.n47 6.59444
R1563 VDD1.n47 VDD1.n12 6.59444
R1564 VDD1.n118 VDD1.n83 6.59444
R1565 VDD1.n119 VDD1.n118 6.59444
R1566 VDD1.n68 VDD1.n0 6.08283
R1567 VDD1.n139 VDD1.n71 6.08283
R1568 VDD1.n51 VDD1.n10 5.81868
R1569 VDD1.n44 VDD1.n43 5.81868
R1570 VDD1.n115 VDD1.n114 5.81868
R1571 VDD1.n122 VDD1.n81 5.81868
R1572 VDD1.n52 VDD1.n8 5.04292
R1573 VDD1.n40 VDD1.n14 5.04292
R1574 VDD1.n111 VDD1.n85 5.04292
R1575 VDD1.n123 VDD1.n79 5.04292
R1576 VDD1.n56 VDD1.n55 4.26717
R1577 VDD1.n39 VDD1.n16 4.26717
R1578 VDD1.n110 VDD1.n87 4.26717
R1579 VDD1.n127 VDD1.n126 4.26717
R1580 VDD1.n23 VDD1.n21 3.70982
R1581 VDD1.n94 VDD1.n92 3.70982
R1582 VDD1.n59 VDD1.n6 3.49141
R1583 VDD1.n36 VDD1.n35 3.49141
R1584 VDD1.n107 VDD1.n106 3.49141
R1585 VDD1.n130 VDD1.n77 3.49141
R1586 VDD1.n60 VDD1.n4 2.71565
R1587 VDD1.n32 VDD1.n18 2.71565
R1588 VDD1.n103 VDD1.n89 2.71565
R1589 VDD1.n131 VDD1.n75 2.71565
R1590 VDD1.n64 VDD1.n63 1.93989
R1591 VDD1.n31 VDD1.n20 1.93989
R1592 VDD1.n102 VDD1.n91 1.93989
R1593 VDD1.n135 VDD1.n134 1.93989
R1594 VDD1.n67 VDD1.n2 1.16414
R1595 VDD1.n28 VDD1.n27 1.16414
R1596 VDD1.n99 VDD1.n98 1.16414
R1597 VDD1.n138 VDD1.n73 1.16414
R1598 VDD1.n24 VDD1.n22 0.388379
R1599 VDD1.n95 VDD1.n93 0.388379
R1600 VDD1.n69 VDD1.n1 0.155672
R1601 VDD1.n62 VDD1.n1 0.155672
R1602 VDD1.n62 VDD1.n61 0.155672
R1603 VDD1.n61 VDD1.n5 0.155672
R1604 VDD1.n54 VDD1.n5 0.155672
R1605 VDD1.n54 VDD1.n53 0.155672
R1606 VDD1.n53 VDD1.n9 0.155672
R1607 VDD1.n46 VDD1.n9 0.155672
R1608 VDD1.n46 VDD1.n45 0.155672
R1609 VDD1.n45 VDD1.n13 0.155672
R1610 VDD1.n38 VDD1.n13 0.155672
R1611 VDD1.n38 VDD1.n37 0.155672
R1612 VDD1.n37 VDD1.n17 0.155672
R1613 VDD1.n30 VDD1.n17 0.155672
R1614 VDD1.n30 VDD1.n29 0.155672
R1615 VDD1.n29 VDD1.n21 0.155672
R1616 VDD1.n100 VDD1.n92 0.155672
R1617 VDD1.n101 VDD1.n100 0.155672
R1618 VDD1.n101 VDD1.n88 0.155672
R1619 VDD1.n108 VDD1.n88 0.155672
R1620 VDD1.n109 VDD1.n108 0.155672
R1621 VDD1.n109 VDD1.n84 0.155672
R1622 VDD1.n116 VDD1.n84 0.155672
R1623 VDD1.n117 VDD1.n116 0.155672
R1624 VDD1.n117 VDD1.n80 0.155672
R1625 VDD1.n124 VDD1.n80 0.155672
R1626 VDD1.n125 VDD1.n124 0.155672
R1627 VDD1.n125 VDD1.n76 0.155672
R1628 VDD1.n132 VDD1.n76 0.155672
R1629 VDD1.n133 VDD1.n132 0.155672
R1630 VDD1.n133 VDD1.n72 0.155672
R1631 VDD1.n140 VDD1.n72 0.155672
R1632 VN VN.t0 188.775
R1633 VN VN.t1 142.238
R1634 VDD2.n138 VDD2.n137 585
R1635 VDD2.n136 VDD2.n135 585
R1636 VDD2.n75 VDD2.n74 585
R1637 VDD2.n130 VDD2.n129 585
R1638 VDD2.n128 VDD2.n127 585
R1639 VDD2.n79 VDD2.n78 585
R1640 VDD2.n122 VDD2.n121 585
R1641 VDD2.n120 VDD2.n119 585
R1642 VDD2.n83 VDD2.n82 585
R1643 VDD2.n114 VDD2.n113 585
R1644 VDD2.n112 VDD2.n111 585
R1645 VDD2.n87 VDD2.n86 585
R1646 VDD2.n106 VDD2.n105 585
R1647 VDD2.n104 VDD2.n103 585
R1648 VDD2.n91 VDD2.n90 585
R1649 VDD2.n98 VDD2.n97 585
R1650 VDD2.n96 VDD2.n95 585
R1651 VDD2.n25 VDD2.n24 585
R1652 VDD2.n27 VDD2.n26 585
R1653 VDD2.n20 VDD2.n19 585
R1654 VDD2.n33 VDD2.n32 585
R1655 VDD2.n35 VDD2.n34 585
R1656 VDD2.n16 VDD2.n15 585
R1657 VDD2.n41 VDD2.n40 585
R1658 VDD2.n43 VDD2.n42 585
R1659 VDD2.n12 VDD2.n11 585
R1660 VDD2.n49 VDD2.n48 585
R1661 VDD2.n51 VDD2.n50 585
R1662 VDD2.n8 VDD2.n7 585
R1663 VDD2.n57 VDD2.n56 585
R1664 VDD2.n59 VDD2.n58 585
R1665 VDD2.n4 VDD2.n3 585
R1666 VDD2.n65 VDD2.n64 585
R1667 VDD2.n67 VDD2.n66 585
R1668 VDD2.n137 VDD2.n71 498.474
R1669 VDD2.n66 VDD2.n0 498.474
R1670 VDD2.n94 VDD2.t1 327.466
R1671 VDD2.n23 VDD2.t0 327.466
R1672 VDD2.n137 VDD2.n136 171.744
R1673 VDD2.n136 VDD2.n74 171.744
R1674 VDD2.n129 VDD2.n74 171.744
R1675 VDD2.n129 VDD2.n128 171.744
R1676 VDD2.n128 VDD2.n78 171.744
R1677 VDD2.n121 VDD2.n78 171.744
R1678 VDD2.n121 VDD2.n120 171.744
R1679 VDD2.n120 VDD2.n82 171.744
R1680 VDD2.n113 VDD2.n82 171.744
R1681 VDD2.n113 VDD2.n112 171.744
R1682 VDD2.n112 VDD2.n86 171.744
R1683 VDD2.n105 VDD2.n86 171.744
R1684 VDD2.n105 VDD2.n104 171.744
R1685 VDD2.n104 VDD2.n90 171.744
R1686 VDD2.n97 VDD2.n90 171.744
R1687 VDD2.n97 VDD2.n96 171.744
R1688 VDD2.n26 VDD2.n25 171.744
R1689 VDD2.n26 VDD2.n19 171.744
R1690 VDD2.n33 VDD2.n19 171.744
R1691 VDD2.n34 VDD2.n33 171.744
R1692 VDD2.n34 VDD2.n15 171.744
R1693 VDD2.n41 VDD2.n15 171.744
R1694 VDD2.n42 VDD2.n41 171.744
R1695 VDD2.n42 VDD2.n11 171.744
R1696 VDD2.n49 VDD2.n11 171.744
R1697 VDD2.n50 VDD2.n49 171.744
R1698 VDD2.n50 VDD2.n7 171.744
R1699 VDD2.n57 VDD2.n7 171.744
R1700 VDD2.n58 VDD2.n57 171.744
R1701 VDD2.n58 VDD2.n3 171.744
R1702 VDD2.n65 VDD2.n3 171.744
R1703 VDD2.n66 VDD2.n65 171.744
R1704 VDD2.n142 VDD2.n70 94.1394
R1705 VDD2.n96 VDD2.t1 85.8723
R1706 VDD2.n25 VDD2.t0 85.8723
R1707 VDD2.n142 VDD2.n141 52.9369
R1708 VDD2.n95 VDD2.n94 16.3895
R1709 VDD2.n24 VDD2.n23 16.3895
R1710 VDD2.n139 VDD2.n138 12.8005
R1711 VDD2.n98 VDD2.n93 12.8005
R1712 VDD2.n27 VDD2.n22 12.8005
R1713 VDD2.n68 VDD2.n67 12.8005
R1714 VDD2.n135 VDD2.n73 12.0247
R1715 VDD2.n99 VDD2.n91 12.0247
R1716 VDD2.n28 VDD2.n20 12.0247
R1717 VDD2.n64 VDD2.n2 12.0247
R1718 VDD2.n134 VDD2.n75 11.249
R1719 VDD2.n103 VDD2.n102 11.249
R1720 VDD2.n32 VDD2.n31 11.249
R1721 VDD2.n63 VDD2.n4 11.249
R1722 VDD2.n131 VDD2.n130 10.4732
R1723 VDD2.n106 VDD2.n89 10.4732
R1724 VDD2.n35 VDD2.n18 10.4732
R1725 VDD2.n60 VDD2.n59 10.4732
R1726 VDD2.n127 VDD2.n77 9.69747
R1727 VDD2.n107 VDD2.n87 9.69747
R1728 VDD2.n36 VDD2.n16 9.69747
R1729 VDD2.n56 VDD2.n6 9.69747
R1730 VDD2.n141 VDD2.n140 9.45567
R1731 VDD2.n70 VDD2.n69 9.45567
R1732 VDD2.n81 VDD2.n80 9.3005
R1733 VDD2.n124 VDD2.n123 9.3005
R1734 VDD2.n126 VDD2.n125 9.3005
R1735 VDD2.n77 VDD2.n76 9.3005
R1736 VDD2.n132 VDD2.n131 9.3005
R1737 VDD2.n134 VDD2.n133 9.3005
R1738 VDD2.n73 VDD2.n72 9.3005
R1739 VDD2.n140 VDD2.n139 9.3005
R1740 VDD2.n118 VDD2.n117 9.3005
R1741 VDD2.n116 VDD2.n115 9.3005
R1742 VDD2.n85 VDD2.n84 9.3005
R1743 VDD2.n110 VDD2.n109 9.3005
R1744 VDD2.n108 VDD2.n107 9.3005
R1745 VDD2.n89 VDD2.n88 9.3005
R1746 VDD2.n102 VDD2.n101 9.3005
R1747 VDD2.n100 VDD2.n99 9.3005
R1748 VDD2.n93 VDD2.n92 9.3005
R1749 VDD2.n45 VDD2.n44 9.3005
R1750 VDD2.n14 VDD2.n13 9.3005
R1751 VDD2.n39 VDD2.n38 9.3005
R1752 VDD2.n37 VDD2.n36 9.3005
R1753 VDD2.n18 VDD2.n17 9.3005
R1754 VDD2.n31 VDD2.n30 9.3005
R1755 VDD2.n29 VDD2.n28 9.3005
R1756 VDD2.n22 VDD2.n21 9.3005
R1757 VDD2.n47 VDD2.n46 9.3005
R1758 VDD2.n10 VDD2.n9 9.3005
R1759 VDD2.n53 VDD2.n52 9.3005
R1760 VDD2.n55 VDD2.n54 9.3005
R1761 VDD2.n6 VDD2.n5 9.3005
R1762 VDD2.n61 VDD2.n60 9.3005
R1763 VDD2.n63 VDD2.n62 9.3005
R1764 VDD2.n2 VDD2.n1 9.3005
R1765 VDD2.n69 VDD2.n68 9.3005
R1766 VDD2.n126 VDD2.n79 8.92171
R1767 VDD2.n111 VDD2.n110 8.92171
R1768 VDD2.n40 VDD2.n39 8.92171
R1769 VDD2.n55 VDD2.n8 8.92171
R1770 VDD2.n123 VDD2.n122 8.14595
R1771 VDD2.n114 VDD2.n85 8.14595
R1772 VDD2.n43 VDD2.n14 8.14595
R1773 VDD2.n52 VDD2.n51 8.14595
R1774 VDD2.n141 VDD2.n71 7.75445
R1775 VDD2.n70 VDD2.n0 7.75445
R1776 VDD2.n119 VDD2.n81 7.3702
R1777 VDD2.n115 VDD2.n83 7.3702
R1778 VDD2.n44 VDD2.n12 7.3702
R1779 VDD2.n48 VDD2.n10 7.3702
R1780 VDD2.n119 VDD2.n118 6.59444
R1781 VDD2.n118 VDD2.n83 6.59444
R1782 VDD2.n47 VDD2.n12 6.59444
R1783 VDD2.n48 VDD2.n47 6.59444
R1784 VDD2.n139 VDD2.n71 6.08283
R1785 VDD2.n68 VDD2.n0 6.08283
R1786 VDD2.n122 VDD2.n81 5.81868
R1787 VDD2.n115 VDD2.n114 5.81868
R1788 VDD2.n44 VDD2.n43 5.81868
R1789 VDD2.n51 VDD2.n10 5.81868
R1790 VDD2.n123 VDD2.n79 5.04292
R1791 VDD2.n111 VDD2.n85 5.04292
R1792 VDD2.n40 VDD2.n14 5.04292
R1793 VDD2.n52 VDD2.n8 5.04292
R1794 VDD2.n127 VDD2.n126 4.26717
R1795 VDD2.n110 VDD2.n87 4.26717
R1796 VDD2.n39 VDD2.n16 4.26717
R1797 VDD2.n56 VDD2.n55 4.26717
R1798 VDD2.n94 VDD2.n92 3.70982
R1799 VDD2.n23 VDD2.n21 3.70982
R1800 VDD2.n130 VDD2.n77 3.49141
R1801 VDD2.n107 VDD2.n106 3.49141
R1802 VDD2.n36 VDD2.n35 3.49141
R1803 VDD2.n59 VDD2.n6 3.49141
R1804 VDD2.n131 VDD2.n75 2.71565
R1805 VDD2.n103 VDD2.n89 2.71565
R1806 VDD2.n32 VDD2.n18 2.71565
R1807 VDD2.n60 VDD2.n4 2.71565
R1808 VDD2.n135 VDD2.n134 1.93989
R1809 VDD2.n102 VDD2.n91 1.93989
R1810 VDD2.n31 VDD2.n20 1.93989
R1811 VDD2.n64 VDD2.n63 1.93989
R1812 VDD2.n138 VDD2.n73 1.16414
R1813 VDD2.n99 VDD2.n98 1.16414
R1814 VDD2.n28 VDD2.n27 1.16414
R1815 VDD2.n67 VDD2.n2 1.16414
R1816 VDD2 VDD2.n142 0.806535
R1817 VDD2.n95 VDD2.n93 0.388379
R1818 VDD2.n24 VDD2.n22 0.388379
R1819 VDD2.n140 VDD2.n72 0.155672
R1820 VDD2.n133 VDD2.n72 0.155672
R1821 VDD2.n133 VDD2.n132 0.155672
R1822 VDD2.n132 VDD2.n76 0.155672
R1823 VDD2.n125 VDD2.n76 0.155672
R1824 VDD2.n125 VDD2.n124 0.155672
R1825 VDD2.n124 VDD2.n80 0.155672
R1826 VDD2.n117 VDD2.n80 0.155672
R1827 VDD2.n117 VDD2.n116 0.155672
R1828 VDD2.n116 VDD2.n84 0.155672
R1829 VDD2.n109 VDD2.n84 0.155672
R1830 VDD2.n109 VDD2.n108 0.155672
R1831 VDD2.n108 VDD2.n88 0.155672
R1832 VDD2.n101 VDD2.n88 0.155672
R1833 VDD2.n101 VDD2.n100 0.155672
R1834 VDD2.n100 VDD2.n92 0.155672
R1835 VDD2.n29 VDD2.n21 0.155672
R1836 VDD2.n30 VDD2.n29 0.155672
R1837 VDD2.n30 VDD2.n17 0.155672
R1838 VDD2.n37 VDD2.n17 0.155672
R1839 VDD2.n38 VDD2.n37 0.155672
R1840 VDD2.n38 VDD2.n13 0.155672
R1841 VDD2.n45 VDD2.n13 0.155672
R1842 VDD2.n46 VDD2.n45 0.155672
R1843 VDD2.n46 VDD2.n9 0.155672
R1844 VDD2.n53 VDD2.n9 0.155672
R1845 VDD2.n54 VDD2.n53 0.155672
R1846 VDD2.n54 VDD2.n5 0.155672
R1847 VDD2.n61 VDD2.n5 0.155672
R1848 VDD2.n62 VDD2.n61 0.155672
R1849 VDD2.n62 VDD2.n1 0.155672
R1850 VDD2.n69 VDD2.n1 0.155672
C0 w_n2358_n3650# VN 3.34787f
C1 w_n2358_n3650# VDD1 1.93898f
C2 w_n2358_n3650# VDD2 1.97151f
C3 VDD1 VN 0.14837f
C4 w_n2358_n3650# VP 3.6494f
C5 B w_n2358_n3650# 9.78749f
C6 VDD2 VN 3.1609f
C7 VP VN 5.97466f
C8 B VN 1.15726f
C9 VDD1 VDD2 0.740412f
C10 VDD1 VP 3.36587f
C11 B VDD1 1.89058f
C12 VP VDD2 0.355844f
C13 B VDD2 1.92546f
C14 B VP 1.65515f
C15 w_n2358_n3650# VTAIL 2.94693f
C16 VTAIL VN 2.80045f
C17 VDD1 VTAIL 5.52164f
C18 VTAIL VDD2 5.5761f
C19 VTAIL VP 2.81472f
C20 B VTAIL 4.19003f
C21 VDD2 VSUBS 0.975344f
C22 VDD1 VSUBS 4.02452f
C23 VTAIL VSUBS 1.118992f
C24 VN VSUBS 8.3255f
C25 VP VSUBS 1.902301f
C26 B VSUBS 4.423581f
C27 w_n2358_n3650# VSUBS 0.105742p
C28 VDD2.n0 VSUBS 0.022574f
C29 VDD2.n1 VSUBS 0.020385f
C30 VDD2.n2 VSUBS 0.010954f
C31 VDD2.n3 VSUBS 0.025891f
C32 VDD2.n4 VSUBS 0.011598f
C33 VDD2.n5 VSUBS 0.020385f
C34 VDD2.n6 VSUBS 0.010954f
C35 VDD2.n7 VSUBS 0.025891f
C36 VDD2.n8 VSUBS 0.011598f
C37 VDD2.n9 VSUBS 0.020385f
C38 VDD2.n10 VSUBS 0.010954f
C39 VDD2.n11 VSUBS 0.025891f
C40 VDD2.n12 VSUBS 0.011598f
C41 VDD2.n13 VSUBS 0.020385f
C42 VDD2.n14 VSUBS 0.010954f
C43 VDD2.n15 VSUBS 0.025891f
C44 VDD2.n16 VSUBS 0.011598f
C45 VDD2.n17 VSUBS 0.020385f
C46 VDD2.n18 VSUBS 0.010954f
C47 VDD2.n19 VSUBS 0.025891f
C48 VDD2.n20 VSUBS 0.011598f
C49 VDD2.n21 VSUBS 1.15446f
C50 VDD2.n22 VSUBS 0.010954f
C51 VDD2.t0 VSUBS 0.055348f
C52 VDD2.n23 VSUBS 0.134135f
C53 VDD2.n24 VSUBS 0.016471f
C54 VDD2.n25 VSUBS 0.019418f
C55 VDD2.n26 VSUBS 0.025891f
C56 VDD2.n27 VSUBS 0.011598f
C57 VDD2.n28 VSUBS 0.010954f
C58 VDD2.n29 VSUBS 0.020385f
C59 VDD2.n30 VSUBS 0.020385f
C60 VDD2.n31 VSUBS 0.010954f
C61 VDD2.n32 VSUBS 0.011598f
C62 VDD2.n33 VSUBS 0.025891f
C63 VDD2.n34 VSUBS 0.025891f
C64 VDD2.n35 VSUBS 0.011598f
C65 VDD2.n36 VSUBS 0.010954f
C66 VDD2.n37 VSUBS 0.020385f
C67 VDD2.n38 VSUBS 0.020385f
C68 VDD2.n39 VSUBS 0.010954f
C69 VDD2.n40 VSUBS 0.011598f
C70 VDD2.n41 VSUBS 0.025891f
C71 VDD2.n42 VSUBS 0.025891f
C72 VDD2.n43 VSUBS 0.011598f
C73 VDD2.n44 VSUBS 0.010954f
C74 VDD2.n45 VSUBS 0.020385f
C75 VDD2.n46 VSUBS 0.020385f
C76 VDD2.n47 VSUBS 0.010954f
C77 VDD2.n48 VSUBS 0.011598f
C78 VDD2.n49 VSUBS 0.025891f
C79 VDD2.n50 VSUBS 0.025891f
C80 VDD2.n51 VSUBS 0.011598f
C81 VDD2.n52 VSUBS 0.010954f
C82 VDD2.n53 VSUBS 0.020385f
C83 VDD2.n54 VSUBS 0.020385f
C84 VDD2.n55 VSUBS 0.010954f
C85 VDD2.n56 VSUBS 0.011598f
C86 VDD2.n57 VSUBS 0.025891f
C87 VDD2.n58 VSUBS 0.025891f
C88 VDD2.n59 VSUBS 0.011598f
C89 VDD2.n60 VSUBS 0.010954f
C90 VDD2.n61 VSUBS 0.020385f
C91 VDD2.n62 VSUBS 0.020385f
C92 VDD2.n63 VSUBS 0.010954f
C93 VDD2.n64 VSUBS 0.011598f
C94 VDD2.n65 VSUBS 0.025891f
C95 VDD2.n66 VSUBS 0.065434f
C96 VDD2.n67 VSUBS 0.011598f
C97 VDD2.n68 VSUBS 0.021511f
C98 VDD2.n69 VSUBS 0.052966f
C99 VDD2.n70 VSUBS 0.664077f
C100 VDD2.n71 VSUBS 0.022574f
C101 VDD2.n72 VSUBS 0.020385f
C102 VDD2.n73 VSUBS 0.010954f
C103 VDD2.n74 VSUBS 0.025891f
C104 VDD2.n75 VSUBS 0.011598f
C105 VDD2.n76 VSUBS 0.020385f
C106 VDD2.n77 VSUBS 0.010954f
C107 VDD2.n78 VSUBS 0.025891f
C108 VDD2.n79 VSUBS 0.011598f
C109 VDD2.n80 VSUBS 0.020385f
C110 VDD2.n81 VSUBS 0.010954f
C111 VDD2.n82 VSUBS 0.025891f
C112 VDD2.n83 VSUBS 0.011598f
C113 VDD2.n84 VSUBS 0.020385f
C114 VDD2.n85 VSUBS 0.010954f
C115 VDD2.n86 VSUBS 0.025891f
C116 VDD2.n87 VSUBS 0.011598f
C117 VDD2.n88 VSUBS 0.020385f
C118 VDD2.n89 VSUBS 0.010954f
C119 VDD2.n90 VSUBS 0.025891f
C120 VDD2.n91 VSUBS 0.011598f
C121 VDD2.n92 VSUBS 1.15446f
C122 VDD2.n93 VSUBS 0.010954f
C123 VDD2.t1 VSUBS 0.055348f
C124 VDD2.n94 VSUBS 0.134135f
C125 VDD2.n95 VSUBS 0.016471f
C126 VDD2.n96 VSUBS 0.019418f
C127 VDD2.n97 VSUBS 0.025891f
C128 VDD2.n98 VSUBS 0.011598f
C129 VDD2.n99 VSUBS 0.010954f
C130 VDD2.n100 VSUBS 0.020385f
C131 VDD2.n101 VSUBS 0.020385f
C132 VDD2.n102 VSUBS 0.010954f
C133 VDD2.n103 VSUBS 0.011598f
C134 VDD2.n104 VSUBS 0.025891f
C135 VDD2.n105 VSUBS 0.025891f
C136 VDD2.n106 VSUBS 0.011598f
C137 VDD2.n107 VSUBS 0.010954f
C138 VDD2.n108 VSUBS 0.020385f
C139 VDD2.n109 VSUBS 0.020385f
C140 VDD2.n110 VSUBS 0.010954f
C141 VDD2.n111 VSUBS 0.011598f
C142 VDD2.n112 VSUBS 0.025891f
C143 VDD2.n113 VSUBS 0.025891f
C144 VDD2.n114 VSUBS 0.011598f
C145 VDD2.n115 VSUBS 0.010954f
C146 VDD2.n116 VSUBS 0.020385f
C147 VDD2.n117 VSUBS 0.020385f
C148 VDD2.n118 VSUBS 0.010954f
C149 VDD2.n119 VSUBS 0.011598f
C150 VDD2.n120 VSUBS 0.025891f
C151 VDD2.n121 VSUBS 0.025891f
C152 VDD2.n122 VSUBS 0.011598f
C153 VDD2.n123 VSUBS 0.010954f
C154 VDD2.n124 VSUBS 0.020385f
C155 VDD2.n125 VSUBS 0.020385f
C156 VDD2.n126 VSUBS 0.010954f
C157 VDD2.n127 VSUBS 0.011598f
C158 VDD2.n128 VSUBS 0.025891f
C159 VDD2.n129 VSUBS 0.025891f
C160 VDD2.n130 VSUBS 0.011598f
C161 VDD2.n131 VSUBS 0.010954f
C162 VDD2.n132 VSUBS 0.020385f
C163 VDD2.n133 VSUBS 0.020385f
C164 VDD2.n134 VSUBS 0.010954f
C165 VDD2.n135 VSUBS 0.011598f
C166 VDD2.n136 VSUBS 0.025891f
C167 VDD2.n137 VSUBS 0.065434f
C168 VDD2.n138 VSUBS 0.011598f
C169 VDD2.n139 VSUBS 0.021511f
C170 VDD2.n140 VSUBS 0.052966f
C171 VDD2.n141 VSUBS 0.064756f
C172 VDD2.n142 VSUBS 2.72486f
C173 VN.t1 VSUBS 4.4495f
C174 VN.t0 VSUBS 5.2352f
C175 VDD1.n0 VSUBS 0.022637f
C176 VDD1.n1 VSUBS 0.020441f
C177 VDD1.n2 VSUBS 0.010984f
C178 VDD1.n3 VSUBS 0.025963f
C179 VDD1.n4 VSUBS 0.01163f
C180 VDD1.n5 VSUBS 0.020441f
C181 VDD1.n6 VSUBS 0.010984f
C182 VDD1.n7 VSUBS 0.025963f
C183 VDD1.n8 VSUBS 0.01163f
C184 VDD1.n9 VSUBS 0.020441f
C185 VDD1.n10 VSUBS 0.010984f
C186 VDD1.n11 VSUBS 0.025963f
C187 VDD1.n12 VSUBS 0.01163f
C188 VDD1.n13 VSUBS 0.020441f
C189 VDD1.n14 VSUBS 0.010984f
C190 VDD1.n15 VSUBS 0.025963f
C191 VDD1.n16 VSUBS 0.01163f
C192 VDD1.n17 VSUBS 0.020441f
C193 VDD1.n18 VSUBS 0.010984f
C194 VDD1.n19 VSUBS 0.025963f
C195 VDD1.n20 VSUBS 0.01163f
C196 VDD1.n21 VSUBS 1.15767f
C197 VDD1.n22 VSUBS 0.010984f
C198 VDD1.t0 VSUBS 0.055502f
C199 VDD1.n23 VSUBS 0.134508f
C200 VDD1.n24 VSUBS 0.016516f
C201 VDD1.n25 VSUBS 0.019472f
C202 VDD1.n26 VSUBS 0.025963f
C203 VDD1.n27 VSUBS 0.01163f
C204 VDD1.n28 VSUBS 0.010984f
C205 VDD1.n29 VSUBS 0.020441f
C206 VDD1.n30 VSUBS 0.020441f
C207 VDD1.n31 VSUBS 0.010984f
C208 VDD1.n32 VSUBS 0.01163f
C209 VDD1.n33 VSUBS 0.025963f
C210 VDD1.n34 VSUBS 0.025963f
C211 VDD1.n35 VSUBS 0.01163f
C212 VDD1.n36 VSUBS 0.010984f
C213 VDD1.n37 VSUBS 0.020441f
C214 VDD1.n38 VSUBS 0.020441f
C215 VDD1.n39 VSUBS 0.010984f
C216 VDD1.n40 VSUBS 0.01163f
C217 VDD1.n41 VSUBS 0.025963f
C218 VDD1.n42 VSUBS 0.025963f
C219 VDD1.n43 VSUBS 0.01163f
C220 VDD1.n44 VSUBS 0.010984f
C221 VDD1.n45 VSUBS 0.020441f
C222 VDD1.n46 VSUBS 0.020441f
C223 VDD1.n47 VSUBS 0.010984f
C224 VDD1.n48 VSUBS 0.01163f
C225 VDD1.n49 VSUBS 0.025963f
C226 VDD1.n50 VSUBS 0.025963f
C227 VDD1.n51 VSUBS 0.01163f
C228 VDD1.n52 VSUBS 0.010984f
C229 VDD1.n53 VSUBS 0.020441f
C230 VDD1.n54 VSUBS 0.020441f
C231 VDD1.n55 VSUBS 0.010984f
C232 VDD1.n56 VSUBS 0.01163f
C233 VDD1.n57 VSUBS 0.025963f
C234 VDD1.n58 VSUBS 0.025963f
C235 VDD1.n59 VSUBS 0.01163f
C236 VDD1.n60 VSUBS 0.010984f
C237 VDD1.n61 VSUBS 0.020441f
C238 VDD1.n62 VSUBS 0.020441f
C239 VDD1.n63 VSUBS 0.010984f
C240 VDD1.n64 VSUBS 0.01163f
C241 VDD1.n65 VSUBS 0.025963f
C242 VDD1.n66 VSUBS 0.065616f
C243 VDD1.n67 VSUBS 0.01163f
C244 VDD1.n68 VSUBS 0.021571f
C245 VDD1.n69 VSUBS 0.053113f
C246 VDD1.n70 VSUBS 0.066373f
C247 VDD1.n71 VSUBS 0.022637f
C248 VDD1.n72 VSUBS 0.020441f
C249 VDD1.n73 VSUBS 0.010984f
C250 VDD1.n74 VSUBS 0.025963f
C251 VDD1.n75 VSUBS 0.01163f
C252 VDD1.n76 VSUBS 0.020441f
C253 VDD1.n77 VSUBS 0.010984f
C254 VDD1.n78 VSUBS 0.025963f
C255 VDD1.n79 VSUBS 0.01163f
C256 VDD1.n80 VSUBS 0.020441f
C257 VDD1.n81 VSUBS 0.010984f
C258 VDD1.n82 VSUBS 0.025963f
C259 VDD1.n83 VSUBS 0.01163f
C260 VDD1.n84 VSUBS 0.020441f
C261 VDD1.n85 VSUBS 0.010984f
C262 VDD1.n86 VSUBS 0.025963f
C263 VDD1.n87 VSUBS 0.01163f
C264 VDD1.n88 VSUBS 0.020441f
C265 VDD1.n89 VSUBS 0.010984f
C266 VDD1.n90 VSUBS 0.025963f
C267 VDD1.n91 VSUBS 0.01163f
C268 VDD1.n92 VSUBS 1.15767f
C269 VDD1.n93 VSUBS 0.010984f
C270 VDD1.t1 VSUBS 0.055502f
C271 VDD1.n94 VSUBS 0.134508f
C272 VDD1.n95 VSUBS 0.016516f
C273 VDD1.n96 VSUBS 0.019472f
C274 VDD1.n97 VSUBS 0.025963f
C275 VDD1.n98 VSUBS 0.01163f
C276 VDD1.n99 VSUBS 0.010984f
C277 VDD1.n100 VSUBS 0.020441f
C278 VDD1.n101 VSUBS 0.020441f
C279 VDD1.n102 VSUBS 0.010984f
C280 VDD1.n103 VSUBS 0.01163f
C281 VDD1.n104 VSUBS 0.025963f
C282 VDD1.n105 VSUBS 0.025963f
C283 VDD1.n106 VSUBS 0.01163f
C284 VDD1.n107 VSUBS 0.010984f
C285 VDD1.n108 VSUBS 0.020441f
C286 VDD1.n109 VSUBS 0.020441f
C287 VDD1.n110 VSUBS 0.010984f
C288 VDD1.n111 VSUBS 0.01163f
C289 VDD1.n112 VSUBS 0.025963f
C290 VDD1.n113 VSUBS 0.025963f
C291 VDD1.n114 VSUBS 0.01163f
C292 VDD1.n115 VSUBS 0.010984f
C293 VDD1.n116 VSUBS 0.020441f
C294 VDD1.n117 VSUBS 0.020441f
C295 VDD1.n118 VSUBS 0.010984f
C296 VDD1.n119 VSUBS 0.01163f
C297 VDD1.n120 VSUBS 0.025963f
C298 VDD1.n121 VSUBS 0.025963f
C299 VDD1.n122 VSUBS 0.01163f
C300 VDD1.n123 VSUBS 0.010984f
C301 VDD1.n124 VSUBS 0.020441f
C302 VDD1.n125 VSUBS 0.020441f
C303 VDD1.n126 VSUBS 0.010984f
C304 VDD1.n127 VSUBS 0.01163f
C305 VDD1.n128 VSUBS 0.025963f
C306 VDD1.n129 VSUBS 0.025963f
C307 VDD1.n130 VSUBS 0.01163f
C308 VDD1.n131 VSUBS 0.010984f
C309 VDD1.n132 VSUBS 0.020441f
C310 VDD1.n133 VSUBS 0.020441f
C311 VDD1.n134 VSUBS 0.010984f
C312 VDD1.n135 VSUBS 0.01163f
C313 VDD1.n136 VSUBS 0.025963f
C314 VDD1.n137 VSUBS 0.065616f
C315 VDD1.n138 VSUBS 0.01163f
C316 VDD1.n139 VSUBS 0.021571f
C317 VDD1.n140 VSUBS 0.053113f
C318 VDD1.n141 VSUBS 0.709498f
C319 VTAIL.n0 VSUBS 0.032532f
C320 VTAIL.n1 VSUBS 0.029376f
C321 VTAIL.n2 VSUBS 0.015786f
C322 VTAIL.n3 VSUBS 0.037311f
C323 VTAIL.n4 VSUBS 0.016714f
C324 VTAIL.n5 VSUBS 0.029376f
C325 VTAIL.n6 VSUBS 0.015786f
C326 VTAIL.n7 VSUBS 0.037311f
C327 VTAIL.n8 VSUBS 0.016714f
C328 VTAIL.n9 VSUBS 0.029376f
C329 VTAIL.n10 VSUBS 0.015786f
C330 VTAIL.n11 VSUBS 0.037311f
C331 VTAIL.n12 VSUBS 0.016714f
C332 VTAIL.n13 VSUBS 0.029376f
C333 VTAIL.n14 VSUBS 0.015786f
C334 VTAIL.n15 VSUBS 0.037311f
C335 VTAIL.n16 VSUBS 0.016714f
C336 VTAIL.n17 VSUBS 0.029376f
C337 VTAIL.n18 VSUBS 0.015786f
C338 VTAIL.n19 VSUBS 0.037311f
C339 VTAIL.n20 VSUBS 0.016714f
C340 VTAIL.n21 VSUBS 1.66369f
C341 VTAIL.n22 VSUBS 0.015786f
C342 VTAIL.t2 VSUBS 0.079762f
C343 VTAIL.n23 VSUBS 0.193303f
C344 VTAIL.n24 VSUBS 0.023736f
C345 VTAIL.n25 VSUBS 0.027983f
C346 VTAIL.n26 VSUBS 0.037311f
C347 VTAIL.n27 VSUBS 0.016714f
C348 VTAIL.n28 VSUBS 0.015786f
C349 VTAIL.n29 VSUBS 0.029376f
C350 VTAIL.n30 VSUBS 0.029376f
C351 VTAIL.n31 VSUBS 0.015786f
C352 VTAIL.n32 VSUBS 0.016714f
C353 VTAIL.n33 VSUBS 0.037311f
C354 VTAIL.n34 VSUBS 0.037311f
C355 VTAIL.n35 VSUBS 0.016714f
C356 VTAIL.n36 VSUBS 0.015786f
C357 VTAIL.n37 VSUBS 0.029376f
C358 VTAIL.n38 VSUBS 0.029376f
C359 VTAIL.n39 VSUBS 0.015786f
C360 VTAIL.n40 VSUBS 0.016714f
C361 VTAIL.n41 VSUBS 0.037311f
C362 VTAIL.n42 VSUBS 0.037311f
C363 VTAIL.n43 VSUBS 0.016714f
C364 VTAIL.n44 VSUBS 0.015786f
C365 VTAIL.n45 VSUBS 0.029376f
C366 VTAIL.n46 VSUBS 0.029376f
C367 VTAIL.n47 VSUBS 0.015786f
C368 VTAIL.n48 VSUBS 0.016714f
C369 VTAIL.n49 VSUBS 0.037311f
C370 VTAIL.n50 VSUBS 0.037311f
C371 VTAIL.n51 VSUBS 0.016714f
C372 VTAIL.n52 VSUBS 0.015786f
C373 VTAIL.n53 VSUBS 0.029376f
C374 VTAIL.n54 VSUBS 0.029376f
C375 VTAIL.n55 VSUBS 0.015786f
C376 VTAIL.n56 VSUBS 0.016714f
C377 VTAIL.n57 VSUBS 0.037311f
C378 VTAIL.n58 VSUBS 0.037311f
C379 VTAIL.n59 VSUBS 0.016714f
C380 VTAIL.n60 VSUBS 0.015786f
C381 VTAIL.n61 VSUBS 0.029376f
C382 VTAIL.n62 VSUBS 0.029376f
C383 VTAIL.n63 VSUBS 0.015786f
C384 VTAIL.n64 VSUBS 0.016714f
C385 VTAIL.n65 VSUBS 0.037311f
C386 VTAIL.n66 VSUBS 0.094297f
C387 VTAIL.n67 VSUBS 0.016714f
C388 VTAIL.n68 VSUBS 0.030999f
C389 VTAIL.n69 VSUBS 0.07633f
C390 VTAIL.n70 VSUBS 0.073094f
C391 VTAIL.n71 VSUBS 2.21025f
C392 VTAIL.n72 VSUBS 0.032532f
C393 VTAIL.n73 VSUBS 0.029376f
C394 VTAIL.n74 VSUBS 0.015786f
C395 VTAIL.n75 VSUBS 0.037311f
C396 VTAIL.n76 VSUBS 0.016714f
C397 VTAIL.n77 VSUBS 0.029376f
C398 VTAIL.n78 VSUBS 0.015786f
C399 VTAIL.n79 VSUBS 0.037311f
C400 VTAIL.n80 VSUBS 0.016714f
C401 VTAIL.n81 VSUBS 0.029376f
C402 VTAIL.n82 VSUBS 0.015786f
C403 VTAIL.n83 VSUBS 0.037311f
C404 VTAIL.n84 VSUBS 0.016714f
C405 VTAIL.n85 VSUBS 0.029376f
C406 VTAIL.n86 VSUBS 0.015786f
C407 VTAIL.n87 VSUBS 0.037311f
C408 VTAIL.n88 VSUBS 0.016714f
C409 VTAIL.n89 VSUBS 0.029376f
C410 VTAIL.n90 VSUBS 0.015786f
C411 VTAIL.n91 VSUBS 0.037311f
C412 VTAIL.n92 VSUBS 0.016714f
C413 VTAIL.n93 VSUBS 1.66369f
C414 VTAIL.n94 VSUBS 0.015786f
C415 VTAIL.t0 VSUBS 0.079762f
C416 VTAIL.n95 VSUBS 0.193303f
C417 VTAIL.n96 VSUBS 0.023736f
C418 VTAIL.n97 VSUBS 0.027983f
C419 VTAIL.n98 VSUBS 0.037311f
C420 VTAIL.n99 VSUBS 0.016714f
C421 VTAIL.n100 VSUBS 0.015786f
C422 VTAIL.n101 VSUBS 0.029376f
C423 VTAIL.n102 VSUBS 0.029376f
C424 VTAIL.n103 VSUBS 0.015786f
C425 VTAIL.n104 VSUBS 0.016714f
C426 VTAIL.n105 VSUBS 0.037311f
C427 VTAIL.n106 VSUBS 0.037311f
C428 VTAIL.n107 VSUBS 0.016714f
C429 VTAIL.n108 VSUBS 0.015786f
C430 VTAIL.n109 VSUBS 0.029376f
C431 VTAIL.n110 VSUBS 0.029376f
C432 VTAIL.n111 VSUBS 0.015786f
C433 VTAIL.n112 VSUBS 0.016714f
C434 VTAIL.n113 VSUBS 0.037311f
C435 VTAIL.n114 VSUBS 0.037311f
C436 VTAIL.n115 VSUBS 0.016714f
C437 VTAIL.n116 VSUBS 0.015786f
C438 VTAIL.n117 VSUBS 0.029376f
C439 VTAIL.n118 VSUBS 0.029376f
C440 VTAIL.n119 VSUBS 0.015786f
C441 VTAIL.n120 VSUBS 0.016714f
C442 VTAIL.n121 VSUBS 0.037311f
C443 VTAIL.n122 VSUBS 0.037311f
C444 VTAIL.n123 VSUBS 0.016714f
C445 VTAIL.n124 VSUBS 0.015786f
C446 VTAIL.n125 VSUBS 0.029376f
C447 VTAIL.n126 VSUBS 0.029376f
C448 VTAIL.n127 VSUBS 0.015786f
C449 VTAIL.n128 VSUBS 0.016714f
C450 VTAIL.n129 VSUBS 0.037311f
C451 VTAIL.n130 VSUBS 0.037311f
C452 VTAIL.n131 VSUBS 0.016714f
C453 VTAIL.n132 VSUBS 0.015786f
C454 VTAIL.n133 VSUBS 0.029376f
C455 VTAIL.n134 VSUBS 0.029376f
C456 VTAIL.n135 VSUBS 0.015786f
C457 VTAIL.n136 VSUBS 0.016714f
C458 VTAIL.n137 VSUBS 0.037311f
C459 VTAIL.n138 VSUBS 0.094297f
C460 VTAIL.n139 VSUBS 0.016714f
C461 VTAIL.n140 VSUBS 0.030999f
C462 VTAIL.n141 VSUBS 0.07633f
C463 VTAIL.n142 VSUBS 0.073094f
C464 VTAIL.n143 VSUBS 2.27554f
C465 VTAIL.n144 VSUBS 0.032532f
C466 VTAIL.n145 VSUBS 0.029376f
C467 VTAIL.n146 VSUBS 0.015786f
C468 VTAIL.n147 VSUBS 0.037311f
C469 VTAIL.n148 VSUBS 0.016714f
C470 VTAIL.n149 VSUBS 0.029376f
C471 VTAIL.n150 VSUBS 0.015786f
C472 VTAIL.n151 VSUBS 0.037311f
C473 VTAIL.n152 VSUBS 0.016714f
C474 VTAIL.n153 VSUBS 0.029376f
C475 VTAIL.n154 VSUBS 0.015786f
C476 VTAIL.n155 VSUBS 0.037311f
C477 VTAIL.n156 VSUBS 0.016714f
C478 VTAIL.n157 VSUBS 0.029376f
C479 VTAIL.n158 VSUBS 0.015786f
C480 VTAIL.n159 VSUBS 0.037311f
C481 VTAIL.n160 VSUBS 0.016714f
C482 VTAIL.n161 VSUBS 0.029376f
C483 VTAIL.n162 VSUBS 0.015786f
C484 VTAIL.n163 VSUBS 0.037311f
C485 VTAIL.n164 VSUBS 0.016714f
C486 VTAIL.n165 VSUBS 1.66369f
C487 VTAIL.n166 VSUBS 0.015786f
C488 VTAIL.t3 VSUBS 0.079762f
C489 VTAIL.n167 VSUBS 0.193303f
C490 VTAIL.n168 VSUBS 0.023736f
C491 VTAIL.n169 VSUBS 0.027983f
C492 VTAIL.n170 VSUBS 0.037311f
C493 VTAIL.n171 VSUBS 0.016714f
C494 VTAIL.n172 VSUBS 0.015786f
C495 VTAIL.n173 VSUBS 0.029376f
C496 VTAIL.n174 VSUBS 0.029376f
C497 VTAIL.n175 VSUBS 0.015786f
C498 VTAIL.n176 VSUBS 0.016714f
C499 VTAIL.n177 VSUBS 0.037311f
C500 VTAIL.n178 VSUBS 0.037311f
C501 VTAIL.n179 VSUBS 0.016714f
C502 VTAIL.n180 VSUBS 0.015786f
C503 VTAIL.n181 VSUBS 0.029376f
C504 VTAIL.n182 VSUBS 0.029376f
C505 VTAIL.n183 VSUBS 0.015786f
C506 VTAIL.n184 VSUBS 0.016714f
C507 VTAIL.n185 VSUBS 0.037311f
C508 VTAIL.n186 VSUBS 0.037311f
C509 VTAIL.n187 VSUBS 0.016714f
C510 VTAIL.n188 VSUBS 0.015786f
C511 VTAIL.n189 VSUBS 0.029376f
C512 VTAIL.n190 VSUBS 0.029376f
C513 VTAIL.n191 VSUBS 0.015786f
C514 VTAIL.n192 VSUBS 0.016714f
C515 VTAIL.n193 VSUBS 0.037311f
C516 VTAIL.n194 VSUBS 0.037311f
C517 VTAIL.n195 VSUBS 0.016714f
C518 VTAIL.n196 VSUBS 0.015786f
C519 VTAIL.n197 VSUBS 0.029376f
C520 VTAIL.n198 VSUBS 0.029376f
C521 VTAIL.n199 VSUBS 0.015786f
C522 VTAIL.n200 VSUBS 0.016714f
C523 VTAIL.n201 VSUBS 0.037311f
C524 VTAIL.n202 VSUBS 0.037311f
C525 VTAIL.n203 VSUBS 0.016714f
C526 VTAIL.n204 VSUBS 0.015786f
C527 VTAIL.n205 VSUBS 0.029376f
C528 VTAIL.n206 VSUBS 0.029376f
C529 VTAIL.n207 VSUBS 0.015786f
C530 VTAIL.n208 VSUBS 0.016714f
C531 VTAIL.n209 VSUBS 0.037311f
C532 VTAIL.n210 VSUBS 0.094297f
C533 VTAIL.n211 VSUBS 0.016714f
C534 VTAIL.n212 VSUBS 0.030999f
C535 VTAIL.n213 VSUBS 0.07633f
C536 VTAIL.n214 VSUBS 0.073094f
C537 VTAIL.n215 VSUBS 1.99238f
C538 VTAIL.n216 VSUBS 0.032532f
C539 VTAIL.n217 VSUBS 0.029376f
C540 VTAIL.n218 VSUBS 0.015786f
C541 VTAIL.n219 VSUBS 0.037311f
C542 VTAIL.n220 VSUBS 0.016714f
C543 VTAIL.n221 VSUBS 0.029376f
C544 VTAIL.n222 VSUBS 0.015786f
C545 VTAIL.n223 VSUBS 0.037311f
C546 VTAIL.n224 VSUBS 0.016714f
C547 VTAIL.n225 VSUBS 0.029376f
C548 VTAIL.n226 VSUBS 0.015786f
C549 VTAIL.n227 VSUBS 0.037311f
C550 VTAIL.n228 VSUBS 0.016714f
C551 VTAIL.n229 VSUBS 0.029376f
C552 VTAIL.n230 VSUBS 0.015786f
C553 VTAIL.n231 VSUBS 0.037311f
C554 VTAIL.n232 VSUBS 0.016714f
C555 VTAIL.n233 VSUBS 0.029376f
C556 VTAIL.n234 VSUBS 0.015786f
C557 VTAIL.n235 VSUBS 0.037311f
C558 VTAIL.n236 VSUBS 0.016714f
C559 VTAIL.n237 VSUBS 1.66369f
C560 VTAIL.n238 VSUBS 0.015786f
C561 VTAIL.t1 VSUBS 0.079762f
C562 VTAIL.n239 VSUBS 0.193303f
C563 VTAIL.n240 VSUBS 0.023736f
C564 VTAIL.n241 VSUBS 0.027983f
C565 VTAIL.n242 VSUBS 0.037311f
C566 VTAIL.n243 VSUBS 0.016714f
C567 VTAIL.n244 VSUBS 0.015786f
C568 VTAIL.n245 VSUBS 0.029376f
C569 VTAIL.n246 VSUBS 0.029376f
C570 VTAIL.n247 VSUBS 0.015786f
C571 VTAIL.n248 VSUBS 0.016714f
C572 VTAIL.n249 VSUBS 0.037311f
C573 VTAIL.n250 VSUBS 0.037311f
C574 VTAIL.n251 VSUBS 0.016714f
C575 VTAIL.n252 VSUBS 0.015786f
C576 VTAIL.n253 VSUBS 0.029376f
C577 VTAIL.n254 VSUBS 0.029376f
C578 VTAIL.n255 VSUBS 0.015786f
C579 VTAIL.n256 VSUBS 0.016714f
C580 VTAIL.n257 VSUBS 0.037311f
C581 VTAIL.n258 VSUBS 0.037311f
C582 VTAIL.n259 VSUBS 0.016714f
C583 VTAIL.n260 VSUBS 0.015786f
C584 VTAIL.n261 VSUBS 0.029376f
C585 VTAIL.n262 VSUBS 0.029376f
C586 VTAIL.n263 VSUBS 0.015786f
C587 VTAIL.n264 VSUBS 0.016714f
C588 VTAIL.n265 VSUBS 0.037311f
C589 VTAIL.n266 VSUBS 0.037311f
C590 VTAIL.n267 VSUBS 0.016714f
C591 VTAIL.n268 VSUBS 0.015786f
C592 VTAIL.n269 VSUBS 0.029376f
C593 VTAIL.n270 VSUBS 0.029376f
C594 VTAIL.n271 VSUBS 0.015786f
C595 VTAIL.n272 VSUBS 0.016714f
C596 VTAIL.n273 VSUBS 0.037311f
C597 VTAIL.n274 VSUBS 0.037311f
C598 VTAIL.n275 VSUBS 0.016714f
C599 VTAIL.n276 VSUBS 0.015786f
C600 VTAIL.n277 VSUBS 0.029376f
C601 VTAIL.n278 VSUBS 0.029376f
C602 VTAIL.n279 VSUBS 0.015786f
C603 VTAIL.n280 VSUBS 0.016714f
C604 VTAIL.n281 VSUBS 0.037311f
C605 VTAIL.n282 VSUBS 0.094297f
C606 VTAIL.n283 VSUBS 0.016714f
C607 VTAIL.n284 VSUBS 0.030999f
C608 VTAIL.n285 VSUBS 0.07633f
C609 VTAIL.n286 VSUBS 0.073094f
C610 VTAIL.n287 VSUBS 1.87161f
C611 VP.t1 VSUBS 5.42366f
C612 VP.t0 VSUBS 4.60417f
C613 VP.n0 VSUBS 5.65317f
C614 B.n0 VSUBS 0.004983f
C615 B.n1 VSUBS 0.004983f
C616 B.n2 VSUBS 0.00737f
C617 B.n3 VSUBS 0.005648f
C618 B.n4 VSUBS 0.005648f
C619 B.n5 VSUBS 0.005648f
C620 B.n6 VSUBS 0.005648f
C621 B.n7 VSUBS 0.005648f
C622 B.n8 VSUBS 0.005648f
C623 B.n9 VSUBS 0.005648f
C624 B.n10 VSUBS 0.005648f
C625 B.n11 VSUBS 0.005648f
C626 B.n12 VSUBS 0.005648f
C627 B.n13 VSUBS 0.005648f
C628 B.n14 VSUBS 0.005648f
C629 B.n15 VSUBS 0.005648f
C630 B.n16 VSUBS 0.013668f
C631 B.n17 VSUBS 0.005648f
C632 B.n18 VSUBS 0.005648f
C633 B.n19 VSUBS 0.005648f
C634 B.n20 VSUBS 0.005648f
C635 B.n21 VSUBS 0.005648f
C636 B.n22 VSUBS 0.005648f
C637 B.n23 VSUBS 0.005648f
C638 B.n24 VSUBS 0.005648f
C639 B.n25 VSUBS 0.005648f
C640 B.n26 VSUBS 0.005648f
C641 B.n27 VSUBS 0.005648f
C642 B.n28 VSUBS 0.005648f
C643 B.n29 VSUBS 0.005648f
C644 B.n30 VSUBS 0.005648f
C645 B.n31 VSUBS 0.005648f
C646 B.n32 VSUBS 0.005648f
C647 B.n33 VSUBS 0.005648f
C648 B.n34 VSUBS 0.005648f
C649 B.n35 VSUBS 0.005648f
C650 B.n36 VSUBS 0.005648f
C651 B.n37 VSUBS 0.005648f
C652 B.n38 VSUBS 0.005648f
C653 B.n39 VSUBS 0.005648f
C654 B.t1 VSUBS 0.195898f
C655 B.t2 VSUBS 0.226426f
C656 B.t0 VSUBS 1.55638f
C657 B.n40 VSUBS 0.359118f
C658 B.n41 VSUBS 0.220486f
C659 B.n42 VSUBS 0.005648f
C660 B.n43 VSUBS 0.005648f
C661 B.n44 VSUBS 0.005648f
C662 B.n45 VSUBS 0.005648f
C663 B.t7 VSUBS 0.195901f
C664 B.t8 VSUBS 0.226428f
C665 B.t6 VSUBS 1.55638f
C666 B.n46 VSUBS 0.359116f
C667 B.n47 VSUBS 0.220483f
C668 B.n48 VSUBS 0.005648f
C669 B.n49 VSUBS 0.005648f
C670 B.n50 VSUBS 0.005648f
C671 B.n51 VSUBS 0.005648f
C672 B.n52 VSUBS 0.005648f
C673 B.n53 VSUBS 0.005648f
C674 B.n54 VSUBS 0.005648f
C675 B.n55 VSUBS 0.005648f
C676 B.n56 VSUBS 0.005648f
C677 B.n57 VSUBS 0.005648f
C678 B.n58 VSUBS 0.005648f
C679 B.n59 VSUBS 0.005648f
C680 B.n60 VSUBS 0.005648f
C681 B.n61 VSUBS 0.005648f
C682 B.n62 VSUBS 0.005648f
C683 B.n63 VSUBS 0.005648f
C684 B.n64 VSUBS 0.005648f
C685 B.n65 VSUBS 0.005648f
C686 B.n66 VSUBS 0.005648f
C687 B.n67 VSUBS 0.005648f
C688 B.n68 VSUBS 0.005648f
C689 B.n69 VSUBS 0.005648f
C690 B.n70 VSUBS 0.013668f
C691 B.n71 VSUBS 0.005648f
C692 B.n72 VSUBS 0.005648f
C693 B.n73 VSUBS 0.005648f
C694 B.n74 VSUBS 0.005648f
C695 B.n75 VSUBS 0.005648f
C696 B.n76 VSUBS 0.005648f
C697 B.n77 VSUBS 0.005648f
C698 B.n78 VSUBS 0.005648f
C699 B.n79 VSUBS 0.005648f
C700 B.n80 VSUBS 0.005648f
C701 B.n81 VSUBS 0.005648f
C702 B.n82 VSUBS 0.005648f
C703 B.n83 VSUBS 0.005648f
C704 B.n84 VSUBS 0.005648f
C705 B.n85 VSUBS 0.005648f
C706 B.n86 VSUBS 0.005648f
C707 B.n87 VSUBS 0.005648f
C708 B.n88 VSUBS 0.005648f
C709 B.n89 VSUBS 0.005648f
C710 B.n90 VSUBS 0.005648f
C711 B.n91 VSUBS 0.005648f
C712 B.n92 VSUBS 0.005648f
C713 B.n93 VSUBS 0.005648f
C714 B.n94 VSUBS 0.005648f
C715 B.n95 VSUBS 0.005648f
C716 B.n96 VSUBS 0.005648f
C717 B.n97 VSUBS 0.005648f
C718 B.n98 VSUBS 0.005648f
C719 B.n99 VSUBS 0.013076f
C720 B.n100 VSUBS 0.005648f
C721 B.n101 VSUBS 0.005648f
C722 B.n102 VSUBS 0.005648f
C723 B.n103 VSUBS 0.005648f
C724 B.n104 VSUBS 0.005648f
C725 B.n105 VSUBS 0.005648f
C726 B.n106 VSUBS 0.005648f
C727 B.n107 VSUBS 0.005648f
C728 B.n108 VSUBS 0.005648f
C729 B.n109 VSUBS 0.005648f
C730 B.n110 VSUBS 0.005648f
C731 B.n111 VSUBS 0.005648f
C732 B.n112 VSUBS 0.005648f
C733 B.n113 VSUBS 0.005648f
C734 B.n114 VSUBS 0.005648f
C735 B.n115 VSUBS 0.005648f
C736 B.n116 VSUBS 0.005648f
C737 B.n117 VSUBS 0.005648f
C738 B.n118 VSUBS 0.005648f
C739 B.n119 VSUBS 0.005648f
C740 B.n120 VSUBS 0.005648f
C741 B.n121 VSUBS 0.005648f
C742 B.n122 VSUBS 0.003904f
C743 B.n123 VSUBS 0.005648f
C744 B.n124 VSUBS 0.005648f
C745 B.n125 VSUBS 0.005648f
C746 B.n126 VSUBS 0.005648f
C747 B.n127 VSUBS 0.005648f
C748 B.t5 VSUBS 0.195898f
C749 B.t4 VSUBS 0.226426f
C750 B.t3 VSUBS 1.55638f
C751 B.n128 VSUBS 0.359118f
C752 B.n129 VSUBS 0.220486f
C753 B.n130 VSUBS 0.005648f
C754 B.n131 VSUBS 0.005648f
C755 B.n132 VSUBS 0.005648f
C756 B.n133 VSUBS 0.005648f
C757 B.n134 VSUBS 0.005648f
C758 B.n135 VSUBS 0.005648f
C759 B.n136 VSUBS 0.005648f
C760 B.n137 VSUBS 0.005648f
C761 B.n138 VSUBS 0.005648f
C762 B.n139 VSUBS 0.005648f
C763 B.n140 VSUBS 0.005648f
C764 B.n141 VSUBS 0.005648f
C765 B.n142 VSUBS 0.005648f
C766 B.n143 VSUBS 0.005648f
C767 B.n144 VSUBS 0.005648f
C768 B.n145 VSUBS 0.005648f
C769 B.n146 VSUBS 0.005648f
C770 B.n147 VSUBS 0.005648f
C771 B.n148 VSUBS 0.005648f
C772 B.n149 VSUBS 0.005648f
C773 B.n150 VSUBS 0.005648f
C774 B.n151 VSUBS 0.005648f
C775 B.n152 VSUBS 0.013076f
C776 B.n153 VSUBS 0.005648f
C777 B.n154 VSUBS 0.005648f
C778 B.n155 VSUBS 0.005648f
C779 B.n156 VSUBS 0.005648f
C780 B.n157 VSUBS 0.005648f
C781 B.n158 VSUBS 0.005648f
C782 B.n159 VSUBS 0.005648f
C783 B.n160 VSUBS 0.005648f
C784 B.n161 VSUBS 0.005648f
C785 B.n162 VSUBS 0.005648f
C786 B.n163 VSUBS 0.005648f
C787 B.n164 VSUBS 0.005648f
C788 B.n165 VSUBS 0.005648f
C789 B.n166 VSUBS 0.005648f
C790 B.n167 VSUBS 0.005648f
C791 B.n168 VSUBS 0.005648f
C792 B.n169 VSUBS 0.005648f
C793 B.n170 VSUBS 0.005648f
C794 B.n171 VSUBS 0.005648f
C795 B.n172 VSUBS 0.005648f
C796 B.n173 VSUBS 0.005648f
C797 B.n174 VSUBS 0.005648f
C798 B.n175 VSUBS 0.005648f
C799 B.n176 VSUBS 0.005648f
C800 B.n177 VSUBS 0.005648f
C801 B.n178 VSUBS 0.005648f
C802 B.n179 VSUBS 0.005648f
C803 B.n180 VSUBS 0.005648f
C804 B.n181 VSUBS 0.005648f
C805 B.n182 VSUBS 0.005648f
C806 B.n183 VSUBS 0.005648f
C807 B.n184 VSUBS 0.005648f
C808 B.n185 VSUBS 0.005648f
C809 B.n186 VSUBS 0.005648f
C810 B.n187 VSUBS 0.005648f
C811 B.n188 VSUBS 0.005648f
C812 B.n189 VSUBS 0.005648f
C813 B.n190 VSUBS 0.005648f
C814 B.n191 VSUBS 0.005648f
C815 B.n192 VSUBS 0.005648f
C816 B.n193 VSUBS 0.005648f
C817 B.n194 VSUBS 0.005648f
C818 B.n195 VSUBS 0.005648f
C819 B.n196 VSUBS 0.005648f
C820 B.n197 VSUBS 0.005648f
C821 B.n198 VSUBS 0.005648f
C822 B.n199 VSUBS 0.005648f
C823 B.n200 VSUBS 0.005648f
C824 B.n201 VSUBS 0.005648f
C825 B.n202 VSUBS 0.005648f
C826 B.n203 VSUBS 0.005648f
C827 B.n204 VSUBS 0.005648f
C828 B.n205 VSUBS 0.013076f
C829 B.n206 VSUBS 0.013668f
C830 B.n207 VSUBS 0.013668f
C831 B.n208 VSUBS 0.005648f
C832 B.n209 VSUBS 0.005648f
C833 B.n210 VSUBS 0.005648f
C834 B.n211 VSUBS 0.005648f
C835 B.n212 VSUBS 0.005648f
C836 B.n213 VSUBS 0.005648f
C837 B.n214 VSUBS 0.005648f
C838 B.n215 VSUBS 0.005648f
C839 B.n216 VSUBS 0.005648f
C840 B.n217 VSUBS 0.005648f
C841 B.n218 VSUBS 0.005648f
C842 B.n219 VSUBS 0.005648f
C843 B.n220 VSUBS 0.005648f
C844 B.n221 VSUBS 0.005648f
C845 B.n222 VSUBS 0.005648f
C846 B.n223 VSUBS 0.005648f
C847 B.n224 VSUBS 0.005648f
C848 B.n225 VSUBS 0.005648f
C849 B.n226 VSUBS 0.005648f
C850 B.n227 VSUBS 0.005648f
C851 B.n228 VSUBS 0.005648f
C852 B.n229 VSUBS 0.005648f
C853 B.n230 VSUBS 0.005648f
C854 B.n231 VSUBS 0.005648f
C855 B.n232 VSUBS 0.005648f
C856 B.n233 VSUBS 0.005648f
C857 B.n234 VSUBS 0.005648f
C858 B.n235 VSUBS 0.005648f
C859 B.n236 VSUBS 0.005648f
C860 B.n237 VSUBS 0.005648f
C861 B.n238 VSUBS 0.005648f
C862 B.n239 VSUBS 0.005648f
C863 B.n240 VSUBS 0.005648f
C864 B.n241 VSUBS 0.005648f
C865 B.n242 VSUBS 0.005648f
C866 B.n243 VSUBS 0.005648f
C867 B.n244 VSUBS 0.005648f
C868 B.n245 VSUBS 0.005648f
C869 B.n246 VSUBS 0.005648f
C870 B.n247 VSUBS 0.005648f
C871 B.n248 VSUBS 0.005648f
C872 B.n249 VSUBS 0.005648f
C873 B.n250 VSUBS 0.005648f
C874 B.n251 VSUBS 0.005648f
C875 B.n252 VSUBS 0.005648f
C876 B.n253 VSUBS 0.005648f
C877 B.n254 VSUBS 0.005648f
C878 B.n255 VSUBS 0.005648f
C879 B.n256 VSUBS 0.005648f
C880 B.n257 VSUBS 0.005648f
C881 B.n258 VSUBS 0.005648f
C882 B.n259 VSUBS 0.005648f
C883 B.n260 VSUBS 0.005648f
C884 B.n261 VSUBS 0.005648f
C885 B.n262 VSUBS 0.005648f
C886 B.n263 VSUBS 0.005648f
C887 B.n264 VSUBS 0.005648f
C888 B.n265 VSUBS 0.005648f
C889 B.n266 VSUBS 0.005648f
C890 B.n267 VSUBS 0.005648f
C891 B.n268 VSUBS 0.005648f
C892 B.n269 VSUBS 0.005648f
C893 B.n270 VSUBS 0.005648f
C894 B.n271 VSUBS 0.005648f
C895 B.n272 VSUBS 0.005648f
C896 B.n273 VSUBS 0.005648f
C897 B.n274 VSUBS 0.003904f
C898 B.n275 VSUBS 0.013085f
C899 B.n276 VSUBS 0.004568f
C900 B.n277 VSUBS 0.005648f
C901 B.n278 VSUBS 0.005648f
C902 B.n279 VSUBS 0.005648f
C903 B.n280 VSUBS 0.005648f
C904 B.n281 VSUBS 0.005648f
C905 B.n282 VSUBS 0.005648f
C906 B.n283 VSUBS 0.005648f
C907 B.n284 VSUBS 0.005648f
C908 B.n285 VSUBS 0.005648f
C909 B.n286 VSUBS 0.005648f
C910 B.n287 VSUBS 0.005648f
C911 B.t11 VSUBS 0.195901f
C912 B.t10 VSUBS 0.226428f
C913 B.t9 VSUBS 1.55638f
C914 B.n288 VSUBS 0.359116f
C915 B.n289 VSUBS 0.220483f
C916 B.n290 VSUBS 0.013085f
C917 B.n291 VSUBS 0.004568f
C918 B.n292 VSUBS 0.005648f
C919 B.n293 VSUBS 0.005648f
C920 B.n294 VSUBS 0.005648f
C921 B.n295 VSUBS 0.005648f
C922 B.n296 VSUBS 0.005648f
C923 B.n297 VSUBS 0.005648f
C924 B.n298 VSUBS 0.005648f
C925 B.n299 VSUBS 0.005648f
C926 B.n300 VSUBS 0.005648f
C927 B.n301 VSUBS 0.005648f
C928 B.n302 VSUBS 0.005648f
C929 B.n303 VSUBS 0.005648f
C930 B.n304 VSUBS 0.005648f
C931 B.n305 VSUBS 0.005648f
C932 B.n306 VSUBS 0.005648f
C933 B.n307 VSUBS 0.005648f
C934 B.n308 VSUBS 0.005648f
C935 B.n309 VSUBS 0.005648f
C936 B.n310 VSUBS 0.005648f
C937 B.n311 VSUBS 0.005648f
C938 B.n312 VSUBS 0.005648f
C939 B.n313 VSUBS 0.005648f
C940 B.n314 VSUBS 0.005648f
C941 B.n315 VSUBS 0.005648f
C942 B.n316 VSUBS 0.005648f
C943 B.n317 VSUBS 0.005648f
C944 B.n318 VSUBS 0.005648f
C945 B.n319 VSUBS 0.005648f
C946 B.n320 VSUBS 0.005648f
C947 B.n321 VSUBS 0.005648f
C948 B.n322 VSUBS 0.005648f
C949 B.n323 VSUBS 0.005648f
C950 B.n324 VSUBS 0.005648f
C951 B.n325 VSUBS 0.005648f
C952 B.n326 VSUBS 0.005648f
C953 B.n327 VSUBS 0.005648f
C954 B.n328 VSUBS 0.005648f
C955 B.n329 VSUBS 0.005648f
C956 B.n330 VSUBS 0.005648f
C957 B.n331 VSUBS 0.005648f
C958 B.n332 VSUBS 0.005648f
C959 B.n333 VSUBS 0.005648f
C960 B.n334 VSUBS 0.005648f
C961 B.n335 VSUBS 0.005648f
C962 B.n336 VSUBS 0.005648f
C963 B.n337 VSUBS 0.005648f
C964 B.n338 VSUBS 0.005648f
C965 B.n339 VSUBS 0.005648f
C966 B.n340 VSUBS 0.005648f
C967 B.n341 VSUBS 0.005648f
C968 B.n342 VSUBS 0.005648f
C969 B.n343 VSUBS 0.005648f
C970 B.n344 VSUBS 0.005648f
C971 B.n345 VSUBS 0.005648f
C972 B.n346 VSUBS 0.005648f
C973 B.n347 VSUBS 0.005648f
C974 B.n348 VSUBS 0.005648f
C975 B.n349 VSUBS 0.005648f
C976 B.n350 VSUBS 0.005648f
C977 B.n351 VSUBS 0.005648f
C978 B.n352 VSUBS 0.005648f
C979 B.n353 VSUBS 0.005648f
C980 B.n354 VSUBS 0.005648f
C981 B.n355 VSUBS 0.005648f
C982 B.n356 VSUBS 0.005648f
C983 B.n357 VSUBS 0.005648f
C984 B.n358 VSUBS 0.005648f
C985 B.n359 VSUBS 0.005648f
C986 B.n360 VSUBS 0.013668f
C987 B.n361 VSUBS 0.013012f
C988 B.n362 VSUBS 0.013732f
C989 B.n363 VSUBS 0.005648f
C990 B.n364 VSUBS 0.005648f
C991 B.n365 VSUBS 0.005648f
C992 B.n366 VSUBS 0.005648f
C993 B.n367 VSUBS 0.005648f
C994 B.n368 VSUBS 0.005648f
C995 B.n369 VSUBS 0.005648f
C996 B.n370 VSUBS 0.005648f
C997 B.n371 VSUBS 0.005648f
C998 B.n372 VSUBS 0.005648f
C999 B.n373 VSUBS 0.005648f
C1000 B.n374 VSUBS 0.005648f
C1001 B.n375 VSUBS 0.005648f
C1002 B.n376 VSUBS 0.005648f
C1003 B.n377 VSUBS 0.005648f
C1004 B.n378 VSUBS 0.005648f
C1005 B.n379 VSUBS 0.005648f
C1006 B.n380 VSUBS 0.005648f
C1007 B.n381 VSUBS 0.005648f
C1008 B.n382 VSUBS 0.005648f
C1009 B.n383 VSUBS 0.005648f
C1010 B.n384 VSUBS 0.005648f
C1011 B.n385 VSUBS 0.005648f
C1012 B.n386 VSUBS 0.005648f
C1013 B.n387 VSUBS 0.005648f
C1014 B.n388 VSUBS 0.005648f
C1015 B.n389 VSUBS 0.005648f
C1016 B.n390 VSUBS 0.005648f
C1017 B.n391 VSUBS 0.005648f
C1018 B.n392 VSUBS 0.005648f
C1019 B.n393 VSUBS 0.005648f
C1020 B.n394 VSUBS 0.005648f
C1021 B.n395 VSUBS 0.005648f
C1022 B.n396 VSUBS 0.005648f
C1023 B.n397 VSUBS 0.005648f
C1024 B.n398 VSUBS 0.005648f
C1025 B.n399 VSUBS 0.005648f
C1026 B.n400 VSUBS 0.005648f
C1027 B.n401 VSUBS 0.005648f
C1028 B.n402 VSUBS 0.005648f
C1029 B.n403 VSUBS 0.005648f
C1030 B.n404 VSUBS 0.005648f
C1031 B.n405 VSUBS 0.005648f
C1032 B.n406 VSUBS 0.005648f
C1033 B.n407 VSUBS 0.005648f
C1034 B.n408 VSUBS 0.005648f
C1035 B.n409 VSUBS 0.005648f
C1036 B.n410 VSUBS 0.005648f
C1037 B.n411 VSUBS 0.005648f
C1038 B.n412 VSUBS 0.005648f
C1039 B.n413 VSUBS 0.005648f
C1040 B.n414 VSUBS 0.005648f
C1041 B.n415 VSUBS 0.005648f
C1042 B.n416 VSUBS 0.005648f
C1043 B.n417 VSUBS 0.005648f
C1044 B.n418 VSUBS 0.005648f
C1045 B.n419 VSUBS 0.005648f
C1046 B.n420 VSUBS 0.005648f
C1047 B.n421 VSUBS 0.005648f
C1048 B.n422 VSUBS 0.005648f
C1049 B.n423 VSUBS 0.005648f
C1050 B.n424 VSUBS 0.005648f
C1051 B.n425 VSUBS 0.005648f
C1052 B.n426 VSUBS 0.005648f
C1053 B.n427 VSUBS 0.005648f
C1054 B.n428 VSUBS 0.005648f
C1055 B.n429 VSUBS 0.005648f
C1056 B.n430 VSUBS 0.005648f
C1057 B.n431 VSUBS 0.005648f
C1058 B.n432 VSUBS 0.005648f
C1059 B.n433 VSUBS 0.005648f
C1060 B.n434 VSUBS 0.005648f
C1061 B.n435 VSUBS 0.005648f
C1062 B.n436 VSUBS 0.005648f
C1063 B.n437 VSUBS 0.005648f
C1064 B.n438 VSUBS 0.005648f
C1065 B.n439 VSUBS 0.005648f
C1066 B.n440 VSUBS 0.005648f
C1067 B.n441 VSUBS 0.005648f
C1068 B.n442 VSUBS 0.005648f
C1069 B.n443 VSUBS 0.005648f
C1070 B.n444 VSUBS 0.005648f
C1071 B.n445 VSUBS 0.005648f
C1072 B.n446 VSUBS 0.005648f
C1073 B.n447 VSUBS 0.013076f
C1074 B.n448 VSUBS 0.013076f
C1075 B.n449 VSUBS 0.013668f
C1076 B.n450 VSUBS 0.005648f
C1077 B.n451 VSUBS 0.005648f
C1078 B.n452 VSUBS 0.005648f
C1079 B.n453 VSUBS 0.005648f
C1080 B.n454 VSUBS 0.005648f
C1081 B.n455 VSUBS 0.005648f
C1082 B.n456 VSUBS 0.005648f
C1083 B.n457 VSUBS 0.005648f
C1084 B.n458 VSUBS 0.005648f
C1085 B.n459 VSUBS 0.005648f
C1086 B.n460 VSUBS 0.005648f
C1087 B.n461 VSUBS 0.005648f
C1088 B.n462 VSUBS 0.005648f
C1089 B.n463 VSUBS 0.005648f
C1090 B.n464 VSUBS 0.005648f
C1091 B.n465 VSUBS 0.005648f
C1092 B.n466 VSUBS 0.005648f
C1093 B.n467 VSUBS 0.005648f
C1094 B.n468 VSUBS 0.005648f
C1095 B.n469 VSUBS 0.005648f
C1096 B.n470 VSUBS 0.005648f
C1097 B.n471 VSUBS 0.005648f
C1098 B.n472 VSUBS 0.005648f
C1099 B.n473 VSUBS 0.005648f
C1100 B.n474 VSUBS 0.005648f
C1101 B.n475 VSUBS 0.005648f
C1102 B.n476 VSUBS 0.005648f
C1103 B.n477 VSUBS 0.005648f
C1104 B.n478 VSUBS 0.005648f
C1105 B.n479 VSUBS 0.005648f
C1106 B.n480 VSUBS 0.005648f
C1107 B.n481 VSUBS 0.005648f
C1108 B.n482 VSUBS 0.005648f
C1109 B.n483 VSUBS 0.005648f
C1110 B.n484 VSUBS 0.005648f
C1111 B.n485 VSUBS 0.005648f
C1112 B.n486 VSUBS 0.005648f
C1113 B.n487 VSUBS 0.005648f
C1114 B.n488 VSUBS 0.005648f
C1115 B.n489 VSUBS 0.005648f
C1116 B.n490 VSUBS 0.005648f
C1117 B.n491 VSUBS 0.005648f
C1118 B.n492 VSUBS 0.005648f
C1119 B.n493 VSUBS 0.005648f
C1120 B.n494 VSUBS 0.005648f
C1121 B.n495 VSUBS 0.005648f
C1122 B.n496 VSUBS 0.005648f
C1123 B.n497 VSUBS 0.005648f
C1124 B.n498 VSUBS 0.005648f
C1125 B.n499 VSUBS 0.005648f
C1126 B.n500 VSUBS 0.005648f
C1127 B.n501 VSUBS 0.005648f
C1128 B.n502 VSUBS 0.005648f
C1129 B.n503 VSUBS 0.005648f
C1130 B.n504 VSUBS 0.005648f
C1131 B.n505 VSUBS 0.005648f
C1132 B.n506 VSUBS 0.005648f
C1133 B.n507 VSUBS 0.005648f
C1134 B.n508 VSUBS 0.005648f
C1135 B.n509 VSUBS 0.005648f
C1136 B.n510 VSUBS 0.005648f
C1137 B.n511 VSUBS 0.005648f
C1138 B.n512 VSUBS 0.005648f
C1139 B.n513 VSUBS 0.005648f
C1140 B.n514 VSUBS 0.005648f
C1141 B.n515 VSUBS 0.005648f
C1142 B.n516 VSUBS 0.005648f
C1143 B.n517 VSUBS 0.003904f
C1144 B.n518 VSUBS 0.013085f
C1145 B.n519 VSUBS 0.004568f
C1146 B.n520 VSUBS 0.005648f
C1147 B.n521 VSUBS 0.005648f
C1148 B.n522 VSUBS 0.005648f
C1149 B.n523 VSUBS 0.005648f
C1150 B.n524 VSUBS 0.005648f
C1151 B.n525 VSUBS 0.005648f
C1152 B.n526 VSUBS 0.005648f
C1153 B.n527 VSUBS 0.005648f
C1154 B.n528 VSUBS 0.005648f
C1155 B.n529 VSUBS 0.005648f
C1156 B.n530 VSUBS 0.005648f
C1157 B.n531 VSUBS 0.004568f
C1158 B.n532 VSUBS 0.013085f
C1159 B.n533 VSUBS 0.003904f
C1160 B.n534 VSUBS 0.005648f
C1161 B.n535 VSUBS 0.005648f
C1162 B.n536 VSUBS 0.005648f
C1163 B.n537 VSUBS 0.005648f
C1164 B.n538 VSUBS 0.005648f
C1165 B.n539 VSUBS 0.005648f
C1166 B.n540 VSUBS 0.005648f
C1167 B.n541 VSUBS 0.005648f
C1168 B.n542 VSUBS 0.005648f
C1169 B.n543 VSUBS 0.005648f
C1170 B.n544 VSUBS 0.005648f
C1171 B.n545 VSUBS 0.005648f
C1172 B.n546 VSUBS 0.005648f
C1173 B.n547 VSUBS 0.005648f
C1174 B.n548 VSUBS 0.005648f
C1175 B.n549 VSUBS 0.005648f
C1176 B.n550 VSUBS 0.005648f
C1177 B.n551 VSUBS 0.005648f
C1178 B.n552 VSUBS 0.005648f
C1179 B.n553 VSUBS 0.005648f
C1180 B.n554 VSUBS 0.005648f
C1181 B.n555 VSUBS 0.005648f
C1182 B.n556 VSUBS 0.005648f
C1183 B.n557 VSUBS 0.005648f
C1184 B.n558 VSUBS 0.005648f
C1185 B.n559 VSUBS 0.005648f
C1186 B.n560 VSUBS 0.005648f
C1187 B.n561 VSUBS 0.005648f
C1188 B.n562 VSUBS 0.005648f
C1189 B.n563 VSUBS 0.005648f
C1190 B.n564 VSUBS 0.005648f
C1191 B.n565 VSUBS 0.005648f
C1192 B.n566 VSUBS 0.005648f
C1193 B.n567 VSUBS 0.005648f
C1194 B.n568 VSUBS 0.005648f
C1195 B.n569 VSUBS 0.005648f
C1196 B.n570 VSUBS 0.005648f
C1197 B.n571 VSUBS 0.005648f
C1198 B.n572 VSUBS 0.005648f
C1199 B.n573 VSUBS 0.005648f
C1200 B.n574 VSUBS 0.005648f
C1201 B.n575 VSUBS 0.005648f
C1202 B.n576 VSUBS 0.005648f
C1203 B.n577 VSUBS 0.005648f
C1204 B.n578 VSUBS 0.005648f
C1205 B.n579 VSUBS 0.005648f
C1206 B.n580 VSUBS 0.005648f
C1207 B.n581 VSUBS 0.005648f
C1208 B.n582 VSUBS 0.005648f
C1209 B.n583 VSUBS 0.005648f
C1210 B.n584 VSUBS 0.005648f
C1211 B.n585 VSUBS 0.005648f
C1212 B.n586 VSUBS 0.005648f
C1213 B.n587 VSUBS 0.005648f
C1214 B.n588 VSUBS 0.005648f
C1215 B.n589 VSUBS 0.005648f
C1216 B.n590 VSUBS 0.005648f
C1217 B.n591 VSUBS 0.005648f
C1218 B.n592 VSUBS 0.005648f
C1219 B.n593 VSUBS 0.005648f
C1220 B.n594 VSUBS 0.005648f
C1221 B.n595 VSUBS 0.005648f
C1222 B.n596 VSUBS 0.005648f
C1223 B.n597 VSUBS 0.005648f
C1224 B.n598 VSUBS 0.005648f
C1225 B.n599 VSUBS 0.005648f
C1226 B.n600 VSUBS 0.005648f
C1227 B.n601 VSUBS 0.013668f
C1228 B.n602 VSUBS 0.013076f
C1229 B.n603 VSUBS 0.013076f
C1230 B.n604 VSUBS 0.005648f
C1231 B.n605 VSUBS 0.005648f
C1232 B.n606 VSUBS 0.005648f
C1233 B.n607 VSUBS 0.005648f
C1234 B.n608 VSUBS 0.005648f
C1235 B.n609 VSUBS 0.005648f
C1236 B.n610 VSUBS 0.005648f
C1237 B.n611 VSUBS 0.005648f
C1238 B.n612 VSUBS 0.005648f
C1239 B.n613 VSUBS 0.005648f
C1240 B.n614 VSUBS 0.005648f
C1241 B.n615 VSUBS 0.005648f
C1242 B.n616 VSUBS 0.005648f
C1243 B.n617 VSUBS 0.005648f
C1244 B.n618 VSUBS 0.005648f
C1245 B.n619 VSUBS 0.005648f
C1246 B.n620 VSUBS 0.005648f
C1247 B.n621 VSUBS 0.005648f
C1248 B.n622 VSUBS 0.005648f
C1249 B.n623 VSUBS 0.005648f
C1250 B.n624 VSUBS 0.005648f
C1251 B.n625 VSUBS 0.005648f
C1252 B.n626 VSUBS 0.005648f
C1253 B.n627 VSUBS 0.005648f
C1254 B.n628 VSUBS 0.005648f
C1255 B.n629 VSUBS 0.005648f
C1256 B.n630 VSUBS 0.005648f
C1257 B.n631 VSUBS 0.005648f
C1258 B.n632 VSUBS 0.005648f
C1259 B.n633 VSUBS 0.005648f
C1260 B.n634 VSUBS 0.005648f
C1261 B.n635 VSUBS 0.005648f
C1262 B.n636 VSUBS 0.005648f
C1263 B.n637 VSUBS 0.005648f
C1264 B.n638 VSUBS 0.005648f
C1265 B.n639 VSUBS 0.005648f
C1266 B.n640 VSUBS 0.005648f
C1267 B.n641 VSUBS 0.005648f
C1268 B.n642 VSUBS 0.005648f
C1269 B.n643 VSUBS 0.00737f
C1270 B.n644 VSUBS 0.007851f
C1271 B.n645 VSUBS 0.015612f
.ends

