| units: 500000 tech: sky130A format: MIT
x a_n579_n1047# a_n674_n997# a_n549_n997# a_n1366_n1488# s=30000,700 d=30000,700 l=30 w=600 x=-318 y=-996 sky130_fd_pr__nfet_01v8
x a_n579_201# a_n549_397# a_n674_n997# a_n1366_n1488# s=30000,700 d=30000,700 l=30 w=600 x=289 y=-996 sky130_fd_pr__nfet_01v8
x a_n1366_n1488# a_n1366_n1488# a_n1366_n1488# a_n1366_n1488# d=57000,1390 l=30 w=600 x=897 y=397 sky130_fd_pr__nfet_01v8
x a_n579_201# a_n674_n997# a_n549_397# a_n1366_n1488# s=57000,1390 d=30000,700 l=30 w=600 x=159 y=-996 sky130_fd_pr__nfet_01v8
x a_n579_n1047# a_n549_n997# a_n674_n997# a_n1366_n1488# s=30000,700 d=57000,1390 l=30 w=600 x=-188 y=-996 sky130_fd_pr__nfet_01v8
x a_n1366_n1488# a_n1366_n1488# a_n1366_n1488# a_n1366_n1488# d=57000,1390 l=30 w=600 x=-926 y=397 sky130_fd_pr__nfet_01v8
x a_n579_n1047# a_n549_n997# a_n674_n997# a_n1366_n1488# s=30000,700 d=30000,700 l=30 w=600 x=289 y=397 sky130_fd_pr__nfet_01v8
x a_n579_201# a_n549_397# a_n674_n997# a_n1366_n1488# s=30000,700 d=57000,1390 l=30 w=600 x=549 y=-996 sky130_fd_pr__nfet_01v8
x a_n579_n1047# a_n674_n997# a_n549_n997# a_n1366_n1488# s=57000,1390 d=30000,700 l=30 w=600 x=159 y=397 sky130_fd_pr__nfet_01v8
x a_n579_n1047# a_n549_n997# a_n674_n997# a_n1366_n1488# s=30000,700 d=57000,1390 l=30 w=600 x=549 y=397 sky130_fd_pr__nfet_01v8
x a_n579_201# a_n674_n997# a_n549_397# a_n1366_n1488# s=30000,700 d=30000,700 l=30 w=600 x=419 y=-996 sky130_fd_pr__nfet_01v8
x a_n579_201# a_n549_397# a_n674_n997# a_n1366_n1488# s=30000,700 d=57000,1390 l=30 w=600 x=-188 y=397 sky130_fd_pr__nfet_01v8
x a_n579_n1047# a_n674_n997# a_n549_n997# a_n1366_n1488# s=30000,700 d=30000,700 l=30 w=600 x=419 y=397 sky130_fd_pr__nfet_01v8
x a_n579_201# a_n674_n997# a_n549_397# a_n1366_n1488# s=57000,1390 d=30000,700 l=30 w=600 x=-578 y=397 sky130_fd_pr__nfet_01v8
x a_n579_n1047# a_n674_n997# a_n549_n997# a_n1366_n1488# s=57000,1390 d=30000,700 l=30 w=600 x=-578 y=-996 sky130_fd_pr__nfet_01v8
x a_n1366_n1488# a_n1366_n1488# a_n1366_n1488# a_n1366_n1488# d=57000,1390 l=30 w=600 x=-926 y=-996 sky130_fd_pr__nfet_01v8
x a_n1366_n1488# a_n1366_n1488# a_n1366_n1488# a_n1366_n1488# d=57000,1390 l=30 w=600 x=897 y=-996 sky130_fd_pr__nfet_01v8
x a_n579_201# a_n549_397# a_n674_n997# a_n1366_n1488# s=30000,700 d=30000,700 l=30 w=600 x=-448 y=397 sky130_fd_pr__nfet_01v8
x a_n579_201# a_n674_n997# a_n549_397# a_n1366_n1488# s=30000,700 d=30000,700 l=30 w=600 x=-318 y=397 sky130_fd_pr__nfet_01v8
x a_n579_n1047# a_n549_n997# a_n674_n997# a_n1366_n1488# s=30000,700 d=30000,700 l=30 w=600 x=-448 y=-996 sky130_fd_pr__nfet_01v8
C a_n549_397# a_n579_n1047# 0.2
C a_n579_201# a_n549_397# 0.9
C a_n579_201# a_n579_n1047# 3.2
C a_n549_n997# a_n674_n997# 5.6
C a_n549_397# a_n674_n997# 5.6
C a_n549_n997# a_n549_397# 0.6
C a_n674_n997# a_n579_n1047# 0.8
C a_n549_n997# a_n579_n1047# 0.8
C a_n579_201# a_n674_n997# 0.8
C a_n549_n997# a_n579_201# 0.3
C a_n549_n997#0 2.0
R a_n549_n997# 4368
C a_n549_397#0 2.2
R a_n549_397# 4368
C a_n674_n997#0 3.4
R a_n674_n997# 13714
C a_n579_n1047#0 4.2
R a_n579_n1047# 10536
C a_n579_201#0 4.1
R a_n579_201# 10535
R a_n1366_n1488# 42346
