* NGSPICE file created from diff_pair_sample_1424.ext - technology: sky130A

.subckt diff_pair_sample_1424 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.6871 pd=14.56 as=2.6871 ps=14.56 w=6.89 l=1.04
X1 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=2.6871 pd=14.56 as=0 ps=0 w=6.89 l=1.04
X2 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.6871 pd=14.56 as=2.6871 ps=14.56 w=6.89 l=1.04
X3 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=2.6871 pd=14.56 as=0 ps=0 w=6.89 l=1.04
X4 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.6871 pd=14.56 as=2.6871 ps=14.56 w=6.89 l=1.04
X5 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.6871 pd=14.56 as=0 ps=0 w=6.89 l=1.04
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.6871 pd=14.56 as=0 ps=0 w=6.89 l=1.04
X7 VDD2.t0 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.6871 pd=14.56 as=2.6871 ps=14.56 w=6.89 l=1.04
R0 VN VN.t0 396.01
R1 VN VN.t1 359.017
R2 VTAIL.n1 VTAIL.t2 54.5118
R3 VTAIL.n3 VTAIL.t3 54.5117
R4 VTAIL.n0 VTAIL.t0 54.5117
R5 VTAIL.n2 VTAIL.t1 54.5117
R6 VTAIL.n1 VTAIL.n0 20.6858
R7 VTAIL.n3 VTAIL.n2 19.5048
R8 VTAIL.n2 VTAIL.n1 1.06084
R9 VTAIL VTAIL.n0 0.823776
R10 VTAIL VTAIL.n3 0.237569
R11 VDD2.n0 VDD2.t0 103.168
R12 VDD2.n0 VDD2.t1 71.1905
R13 VDD2 VDD2.n0 0.353948
R14 B.n456 B.n455 585
R15 B.n457 B.n456 585
R16 B.n192 B.n65 585
R17 B.n191 B.n190 585
R18 B.n189 B.n188 585
R19 B.n187 B.n186 585
R20 B.n185 B.n184 585
R21 B.n183 B.n182 585
R22 B.n181 B.n180 585
R23 B.n179 B.n178 585
R24 B.n177 B.n176 585
R25 B.n175 B.n174 585
R26 B.n173 B.n172 585
R27 B.n171 B.n170 585
R28 B.n169 B.n168 585
R29 B.n167 B.n166 585
R30 B.n165 B.n164 585
R31 B.n163 B.n162 585
R32 B.n161 B.n160 585
R33 B.n159 B.n158 585
R34 B.n157 B.n156 585
R35 B.n155 B.n154 585
R36 B.n153 B.n152 585
R37 B.n151 B.n150 585
R38 B.n149 B.n148 585
R39 B.n147 B.n146 585
R40 B.n145 B.n144 585
R41 B.n143 B.n142 585
R42 B.n141 B.n140 585
R43 B.n139 B.n138 585
R44 B.n137 B.n136 585
R45 B.n135 B.n134 585
R46 B.n133 B.n132 585
R47 B.n131 B.n130 585
R48 B.n129 B.n128 585
R49 B.n127 B.n126 585
R50 B.n125 B.n124 585
R51 B.n122 B.n121 585
R52 B.n120 B.n119 585
R53 B.n118 B.n117 585
R54 B.n116 B.n115 585
R55 B.n114 B.n113 585
R56 B.n112 B.n111 585
R57 B.n110 B.n109 585
R58 B.n108 B.n107 585
R59 B.n106 B.n105 585
R60 B.n104 B.n103 585
R61 B.n102 B.n101 585
R62 B.n100 B.n99 585
R63 B.n98 B.n97 585
R64 B.n96 B.n95 585
R65 B.n94 B.n93 585
R66 B.n92 B.n91 585
R67 B.n90 B.n89 585
R68 B.n88 B.n87 585
R69 B.n86 B.n85 585
R70 B.n84 B.n83 585
R71 B.n82 B.n81 585
R72 B.n80 B.n79 585
R73 B.n78 B.n77 585
R74 B.n76 B.n75 585
R75 B.n74 B.n73 585
R76 B.n72 B.n71 585
R77 B.n32 B.n31 585
R78 B.n454 B.n33 585
R79 B.n458 B.n33 585
R80 B.n453 B.n452 585
R81 B.n452 B.n29 585
R82 B.n451 B.n28 585
R83 B.n464 B.n28 585
R84 B.n450 B.n27 585
R85 B.n465 B.n27 585
R86 B.n449 B.n26 585
R87 B.n466 B.n26 585
R88 B.n448 B.n447 585
R89 B.n447 B.n25 585
R90 B.n446 B.n21 585
R91 B.n472 B.n21 585
R92 B.n445 B.n20 585
R93 B.n473 B.n20 585
R94 B.n444 B.n19 585
R95 B.n474 B.n19 585
R96 B.n443 B.n442 585
R97 B.n442 B.n15 585
R98 B.n441 B.n14 585
R99 B.n480 B.n14 585
R100 B.n440 B.n13 585
R101 B.n481 B.n13 585
R102 B.n439 B.n12 585
R103 B.n482 B.n12 585
R104 B.n438 B.n437 585
R105 B.n437 B.n8 585
R106 B.n436 B.n7 585
R107 B.n488 B.n7 585
R108 B.n435 B.n6 585
R109 B.n489 B.n6 585
R110 B.n434 B.n5 585
R111 B.n490 B.n5 585
R112 B.n433 B.n432 585
R113 B.n432 B.n4 585
R114 B.n431 B.n193 585
R115 B.n431 B.n430 585
R116 B.n421 B.n194 585
R117 B.n195 B.n194 585
R118 B.n423 B.n422 585
R119 B.n424 B.n423 585
R120 B.n420 B.n200 585
R121 B.n200 B.n199 585
R122 B.n419 B.n418 585
R123 B.n418 B.n417 585
R124 B.n202 B.n201 585
R125 B.n203 B.n202 585
R126 B.n410 B.n409 585
R127 B.n411 B.n410 585
R128 B.n408 B.n208 585
R129 B.n208 B.n207 585
R130 B.n407 B.n406 585
R131 B.n406 B.n405 585
R132 B.n210 B.n209 585
R133 B.n398 B.n210 585
R134 B.n397 B.n396 585
R135 B.n399 B.n397 585
R136 B.n395 B.n215 585
R137 B.n215 B.n214 585
R138 B.n394 B.n393 585
R139 B.n393 B.n392 585
R140 B.n217 B.n216 585
R141 B.n218 B.n217 585
R142 B.n385 B.n384 585
R143 B.n386 B.n385 585
R144 B.n221 B.n220 585
R145 B.n258 B.n257 585
R146 B.n259 B.n255 585
R147 B.n255 B.n222 585
R148 B.n261 B.n260 585
R149 B.n263 B.n254 585
R150 B.n266 B.n265 585
R151 B.n267 B.n253 585
R152 B.n269 B.n268 585
R153 B.n271 B.n252 585
R154 B.n274 B.n273 585
R155 B.n275 B.n251 585
R156 B.n277 B.n276 585
R157 B.n279 B.n250 585
R158 B.n282 B.n281 585
R159 B.n283 B.n249 585
R160 B.n285 B.n284 585
R161 B.n287 B.n248 585
R162 B.n290 B.n289 585
R163 B.n291 B.n247 585
R164 B.n293 B.n292 585
R165 B.n295 B.n246 585
R166 B.n298 B.n297 585
R167 B.n299 B.n245 585
R168 B.n301 B.n300 585
R169 B.n303 B.n244 585
R170 B.n306 B.n305 585
R171 B.n307 B.n241 585
R172 B.n310 B.n309 585
R173 B.n312 B.n240 585
R174 B.n315 B.n314 585
R175 B.n316 B.n239 585
R176 B.n318 B.n317 585
R177 B.n320 B.n238 585
R178 B.n323 B.n322 585
R179 B.n324 B.n237 585
R180 B.n329 B.n328 585
R181 B.n331 B.n236 585
R182 B.n334 B.n333 585
R183 B.n335 B.n235 585
R184 B.n337 B.n336 585
R185 B.n339 B.n234 585
R186 B.n342 B.n341 585
R187 B.n343 B.n233 585
R188 B.n345 B.n344 585
R189 B.n347 B.n232 585
R190 B.n350 B.n349 585
R191 B.n351 B.n231 585
R192 B.n353 B.n352 585
R193 B.n355 B.n230 585
R194 B.n358 B.n357 585
R195 B.n359 B.n229 585
R196 B.n361 B.n360 585
R197 B.n363 B.n228 585
R198 B.n366 B.n365 585
R199 B.n367 B.n227 585
R200 B.n369 B.n368 585
R201 B.n371 B.n226 585
R202 B.n374 B.n373 585
R203 B.n375 B.n225 585
R204 B.n377 B.n376 585
R205 B.n379 B.n224 585
R206 B.n382 B.n381 585
R207 B.n383 B.n223 585
R208 B.n388 B.n387 585
R209 B.n387 B.n386 585
R210 B.n389 B.n219 585
R211 B.n219 B.n218 585
R212 B.n391 B.n390 585
R213 B.n392 B.n391 585
R214 B.n213 B.n212 585
R215 B.n214 B.n213 585
R216 B.n401 B.n400 585
R217 B.n400 B.n399 585
R218 B.n402 B.n211 585
R219 B.n398 B.n211 585
R220 B.n404 B.n403 585
R221 B.n405 B.n404 585
R222 B.n206 B.n205 585
R223 B.n207 B.n206 585
R224 B.n413 B.n412 585
R225 B.n412 B.n411 585
R226 B.n414 B.n204 585
R227 B.n204 B.n203 585
R228 B.n416 B.n415 585
R229 B.n417 B.n416 585
R230 B.n198 B.n197 585
R231 B.n199 B.n198 585
R232 B.n426 B.n425 585
R233 B.n425 B.n424 585
R234 B.n427 B.n196 585
R235 B.n196 B.n195 585
R236 B.n429 B.n428 585
R237 B.n430 B.n429 585
R238 B.n2 B.n0 585
R239 B.n4 B.n2 585
R240 B.n3 B.n1 585
R241 B.n489 B.n3 585
R242 B.n487 B.n486 585
R243 B.n488 B.n487 585
R244 B.n485 B.n9 585
R245 B.n9 B.n8 585
R246 B.n484 B.n483 585
R247 B.n483 B.n482 585
R248 B.n11 B.n10 585
R249 B.n481 B.n11 585
R250 B.n479 B.n478 585
R251 B.n480 B.n479 585
R252 B.n477 B.n16 585
R253 B.n16 B.n15 585
R254 B.n476 B.n475 585
R255 B.n475 B.n474 585
R256 B.n18 B.n17 585
R257 B.n473 B.n18 585
R258 B.n471 B.n470 585
R259 B.n472 B.n471 585
R260 B.n469 B.n22 585
R261 B.n25 B.n22 585
R262 B.n468 B.n467 585
R263 B.n467 B.n466 585
R264 B.n24 B.n23 585
R265 B.n465 B.n24 585
R266 B.n463 B.n462 585
R267 B.n464 B.n463 585
R268 B.n461 B.n30 585
R269 B.n30 B.n29 585
R270 B.n460 B.n459 585
R271 B.n459 B.n458 585
R272 B.n492 B.n491 585
R273 B.n491 B.n490 585
R274 B.n387 B.n221 516.524
R275 B.n459 B.n32 516.524
R276 B.n385 B.n223 516.524
R277 B.n456 B.n33 516.524
R278 B.n325 B.t9 362.853
R279 B.n242 B.t13 362.853
R280 B.n69 B.t6 362.853
R281 B.n66 B.t2 362.853
R282 B.n457 B.n64 256.663
R283 B.n457 B.n63 256.663
R284 B.n457 B.n62 256.663
R285 B.n457 B.n61 256.663
R286 B.n457 B.n60 256.663
R287 B.n457 B.n59 256.663
R288 B.n457 B.n58 256.663
R289 B.n457 B.n57 256.663
R290 B.n457 B.n56 256.663
R291 B.n457 B.n55 256.663
R292 B.n457 B.n54 256.663
R293 B.n457 B.n53 256.663
R294 B.n457 B.n52 256.663
R295 B.n457 B.n51 256.663
R296 B.n457 B.n50 256.663
R297 B.n457 B.n49 256.663
R298 B.n457 B.n48 256.663
R299 B.n457 B.n47 256.663
R300 B.n457 B.n46 256.663
R301 B.n457 B.n45 256.663
R302 B.n457 B.n44 256.663
R303 B.n457 B.n43 256.663
R304 B.n457 B.n42 256.663
R305 B.n457 B.n41 256.663
R306 B.n457 B.n40 256.663
R307 B.n457 B.n39 256.663
R308 B.n457 B.n38 256.663
R309 B.n457 B.n37 256.663
R310 B.n457 B.n36 256.663
R311 B.n457 B.n35 256.663
R312 B.n457 B.n34 256.663
R313 B.n256 B.n222 256.663
R314 B.n262 B.n222 256.663
R315 B.n264 B.n222 256.663
R316 B.n270 B.n222 256.663
R317 B.n272 B.n222 256.663
R318 B.n278 B.n222 256.663
R319 B.n280 B.n222 256.663
R320 B.n286 B.n222 256.663
R321 B.n288 B.n222 256.663
R322 B.n294 B.n222 256.663
R323 B.n296 B.n222 256.663
R324 B.n302 B.n222 256.663
R325 B.n304 B.n222 256.663
R326 B.n311 B.n222 256.663
R327 B.n313 B.n222 256.663
R328 B.n319 B.n222 256.663
R329 B.n321 B.n222 256.663
R330 B.n330 B.n222 256.663
R331 B.n332 B.n222 256.663
R332 B.n338 B.n222 256.663
R333 B.n340 B.n222 256.663
R334 B.n346 B.n222 256.663
R335 B.n348 B.n222 256.663
R336 B.n354 B.n222 256.663
R337 B.n356 B.n222 256.663
R338 B.n362 B.n222 256.663
R339 B.n364 B.n222 256.663
R340 B.n370 B.n222 256.663
R341 B.n372 B.n222 256.663
R342 B.n378 B.n222 256.663
R343 B.n380 B.n222 256.663
R344 B.n387 B.n219 163.367
R345 B.n391 B.n219 163.367
R346 B.n391 B.n213 163.367
R347 B.n400 B.n213 163.367
R348 B.n400 B.n211 163.367
R349 B.n404 B.n211 163.367
R350 B.n404 B.n206 163.367
R351 B.n412 B.n206 163.367
R352 B.n412 B.n204 163.367
R353 B.n416 B.n204 163.367
R354 B.n416 B.n198 163.367
R355 B.n425 B.n198 163.367
R356 B.n425 B.n196 163.367
R357 B.n429 B.n196 163.367
R358 B.n429 B.n2 163.367
R359 B.n491 B.n2 163.367
R360 B.n491 B.n3 163.367
R361 B.n487 B.n3 163.367
R362 B.n487 B.n9 163.367
R363 B.n483 B.n9 163.367
R364 B.n483 B.n11 163.367
R365 B.n479 B.n11 163.367
R366 B.n479 B.n16 163.367
R367 B.n475 B.n16 163.367
R368 B.n475 B.n18 163.367
R369 B.n471 B.n18 163.367
R370 B.n471 B.n22 163.367
R371 B.n467 B.n22 163.367
R372 B.n467 B.n24 163.367
R373 B.n463 B.n24 163.367
R374 B.n463 B.n30 163.367
R375 B.n459 B.n30 163.367
R376 B.n257 B.n255 163.367
R377 B.n261 B.n255 163.367
R378 B.n265 B.n263 163.367
R379 B.n269 B.n253 163.367
R380 B.n273 B.n271 163.367
R381 B.n277 B.n251 163.367
R382 B.n281 B.n279 163.367
R383 B.n285 B.n249 163.367
R384 B.n289 B.n287 163.367
R385 B.n293 B.n247 163.367
R386 B.n297 B.n295 163.367
R387 B.n301 B.n245 163.367
R388 B.n305 B.n303 163.367
R389 B.n310 B.n241 163.367
R390 B.n314 B.n312 163.367
R391 B.n318 B.n239 163.367
R392 B.n322 B.n320 163.367
R393 B.n329 B.n237 163.367
R394 B.n333 B.n331 163.367
R395 B.n337 B.n235 163.367
R396 B.n341 B.n339 163.367
R397 B.n345 B.n233 163.367
R398 B.n349 B.n347 163.367
R399 B.n353 B.n231 163.367
R400 B.n357 B.n355 163.367
R401 B.n361 B.n229 163.367
R402 B.n365 B.n363 163.367
R403 B.n369 B.n227 163.367
R404 B.n373 B.n371 163.367
R405 B.n377 B.n225 163.367
R406 B.n381 B.n379 163.367
R407 B.n385 B.n217 163.367
R408 B.n393 B.n217 163.367
R409 B.n393 B.n215 163.367
R410 B.n397 B.n215 163.367
R411 B.n397 B.n210 163.367
R412 B.n406 B.n210 163.367
R413 B.n406 B.n208 163.367
R414 B.n410 B.n208 163.367
R415 B.n410 B.n202 163.367
R416 B.n418 B.n202 163.367
R417 B.n418 B.n200 163.367
R418 B.n423 B.n200 163.367
R419 B.n423 B.n194 163.367
R420 B.n431 B.n194 163.367
R421 B.n432 B.n431 163.367
R422 B.n432 B.n5 163.367
R423 B.n6 B.n5 163.367
R424 B.n7 B.n6 163.367
R425 B.n437 B.n7 163.367
R426 B.n437 B.n12 163.367
R427 B.n13 B.n12 163.367
R428 B.n14 B.n13 163.367
R429 B.n442 B.n14 163.367
R430 B.n442 B.n19 163.367
R431 B.n20 B.n19 163.367
R432 B.n21 B.n20 163.367
R433 B.n447 B.n21 163.367
R434 B.n447 B.n26 163.367
R435 B.n27 B.n26 163.367
R436 B.n28 B.n27 163.367
R437 B.n452 B.n28 163.367
R438 B.n452 B.n33 163.367
R439 B.n73 B.n72 163.367
R440 B.n77 B.n76 163.367
R441 B.n81 B.n80 163.367
R442 B.n85 B.n84 163.367
R443 B.n89 B.n88 163.367
R444 B.n93 B.n92 163.367
R445 B.n97 B.n96 163.367
R446 B.n101 B.n100 163.367
R447 B.n105 B.n104 163.367
R448 B.n109 B.n108 163.367
R449 B.n113 B.n112 163.367
R450 B.n117 B.n116 163.367
R451 B.n121 B.n120 163.367
R452 B.n126 B.n125 163.367
R453 B.n130 B.n129 163.367
R454 B.n134 B.n133 163.367
R455 B.n138 B.n137 163.367
R456 B.n142 B.n141 163.367
R457 B.n146 B.n145 163.367
R458 B.n150 B.n149 163.367
R459 B.n154 B.n153 163.367
R460 B.n158 B.n157 163.367
R461 B.n162 B.n161 163.367
R462 B.n166 B.n165 163.367
R463 B.n170 B.n169 163.367
R464 B.n174 B.n173 163.367
R465 B.n178 B.n177 163.367
R466 B.n182 B.n181 163.367
R467 B.n186 B.n185 163.367
R468 B.n190 B.n189 163.367
R469 B.n456 B.n65 163.367
R470 B.n386 B.n222 121.871
R471 B.n458 B.n457 121.871
R472 B.n325 B.t12 97.3253
R473 B.n66 B.t4 97.3253
R474 B.n242 B.t15 97.3176
R475 B.n69 B.t7 97.3176
R476 B.n256 B.n221 71.676
R477 B.n262 B.n261 71.676
R478 B.n265 B.n264 71.676
R479 B.n270 B.n269 71.676
R480 B.n273 B.n272 71.676
R481 B.n278 B.n277 71.676
R482 B.n281 B.n280 71.676
R483 B.n286 B.n285 71.676
R484 B.n289 B.n288 71.676
R485 B.n294 B.n293 71.676
R486 B.n297 B.n296 71.676
R487 B.n302 B.n301 71.676
R488 B.n305 B.n304 71.676
R489 B.n311 B.n310 71.676
R490 B.n314 B.n313 71.676
R491 B.n319 B.n318 71.676
R492 B.n322 B.n321 71.676
R493 B.n330 B.n329 71.676
R494 B.n333 B.n332 71.676
R495 B.n338 B.n337 71.676
R496 B.n341 B.n340 71.676
R497 B.n346 B.n345 71.676
R498 B.n349 B.n348 71.676
R499 B.n354 B.n353 71.676
R500 B.n357 B.n356 71.676
R501 B.n362 B.n361 71.676
R502 B.n365 B.n364 71.676
R503 B.n370 B.n369 71.676
R504 B.n373 B.n372 71.676
R505 B.n378 B.n377 71.676
R506 B.n381 B.n380 71.676
R507 B.n34 B.n32 71.676
R508 B.n73 B.n35 71.676
R509 B.n77 B.n36 71.676
R510 B.n81 B.n37 71.676
R511 B.n85 B.n38 71.676
R512 B.n89 B.n39 71.676
R513 B.n93 B.n40 71.676
R514 B.n97 B.n41 71.676
R515 B.n101 B.n42 71.676
R516 B.n105 B.n43 71.676
R517 B.n109 B.n44 71.676
R518 B.n113 B.n45 71.676
R519 B.n117 B.n46 71.676
R520 B.n121 B.n47 71.676
R521 B.n126 B.n48 71.676
R522 B.n130 B.n49 71.676
R523 B.n134 B.n50 71.676
R524 B.n138 B.n51 71.676
R525 B.n142 B.n52 71.676
R526 B.n146 B.n53 71.676
R527 B.n150 B.n54 71.676
R528 B.n154 B.n55 71.676
R529 B.n158 B.n56 71.676
R530 B.n162 B.n57 71.676
R531 B.n166 B.n58 71.676
R532 B.n170 B.n59 71.676
R533 B.n174 B.n60 71.676
R534 B.n178 B.n61 71.676
R535 B.n182 B.n62 71.676
R536 B.n186 B.n63 71.676
R537 B.n190 B.n64 71.676
R538 B.n65 B.n64 71.676
R539 B.n189 B.n63 71.676
R540 B.n185 B.n62 71.676
R541 B.n181 B.n61 71.676
R542 B.n177 B.n60 71.676
R543 B.n173 B.n59 71.676
R544 B.n169 B.n58 71.676
R545 B.n165 B.n57 71.676
R546 B.n161 B.n56 71.676
R547 B.n157 B.n55 71.676
R548 B.n153 B.n54 71.676
R549 B.n149 B.n53 71.676
R550 B.n145 B.n52 71.676
R551 B.n141 B.n51 71.676
R552 B.n137 B.n50 71.676
R553 B.n133 B.n49 71.676
R554 B.n129 B.n48 71.676
R555 B.n125 B.n47 71.676
R556 B.n120 B.n46 71.676
R557 B.n116 B.n45 71.676
R558 B.n112 B.n44 71.676
R559 B.n108 B.n43 71.676
R560 B.n104 B.n42 71.676
R561 B.n100 B.n41 71.676
R562 B.n96 B.n40 71.676
R563 B.n92 B.n39 71.676
R564 B.n88 B.n38 71.676
R565 B.n84 B.n37 71.676
R566 B.n80 B.n36 71.676
R567 B.n76 B.n35 71.676
R568 B.n72 B.n34 71.676
R569 B.n257 B.n256 71.676
R570 B.n263 B.n262 71.676
R571 B.n264 B.n253 71.676
R572 B.n271 B.n270 71.676
R573 B.n272 B.n251 71.676
R574 B.n279 B.n278 71.676
R575 B.n280 B.n249 71.676
R576 B.n287 B.n286 71.676
R577 B.n288 B.n247 71.676
R578 B.n295 B.n294 71.676
R579 B.n296 B.n245 71.676
R580 B.n303 B.n302 71.676
R581 B.n304 B.n241 71.676
R582 B.n312 B.n311 71.676
R583 B.n313 B.n239 71.676
R584 B.n320 B.n319 71.676
R585 B.n321 B.n237 71.676
R586 B.n331 B.n330 71.676
R587 B.n332 B.n235 71.676
R588 B.n339 B.n338 71.676
R589 B.n340 B.n233 71.676
R590 B.n347 B.n346 71.676
R591 B.n348 B.n231 71.676
R592 B.n355 B.n354 71.676
R593 B.n356 B.n229 71.676
R594 B.n363 B.n362 71.676
R595 B.n364 B.n227 71.676
R596 B.n371 B.n370 71.676
R597 B.n372 B.n225 71.676
R598 B.n379 B.n378 71.676
R599 B.n380 B.n223 71.676
R600 B.n326 B.t11 70.7556
R601 B.n67 B.t5 70.7556
R602 B.n243 B.t14 70.7479
R603 B.n70 B.t8 70.7479
R604 B.n386 B.n218 61.3874
R605 B.n392 B.n218 61.3874
R606 B.n392 B.n214 61.3874
R607 B.n399 B.n214 61.3874
R608 B.n399 B.n398 61.3874
R609 B.n405 B.n207 61.3874
R610 B.n411 B.n207 61.3874
R611 B.n411 B.n203 61.3874
R612 B.n417 B.n203 61.3874
R613 B.n417 B.n199 61.3874
R614 B.n424 B.n199 61.3874
R615 B.n430 B.n195 61.3874
R616 B.n430 B.n4 61.3874
R617 B.n490 B.n4 61.3874
R618 B.n490 B.n489 61.3874
R619 B.n489 B.n488 61.3874
R620 B.n488 B.n8 61.3874
R621 B.n482 B.n481 61.3874
R622 B.n481 B.n480 61.3874
R623 B.n480 B.n15 61.3874
R624 B.n474 B.n15 61.3874
R625 B.n474 B.n473 61.3874
R626 B.n473 B.n472 61.3874
R627 B.n466 B.n25 61.3874
R628 B.n466 B.n465 61.3874
R629 B.n465 B.n464 61.3874
R630 B.n464 B.n29 61.3874
R631 B.n458 B.n29 61.3874
R632 B.n327 B.n326 59.5399
R633 B.n308 B.n243 59.5399
R634 B.n123 B.n70 59.5399
R635 B.n68 B.n67 59.5399
R636 B.n405 B.t10 52.36
R637 B.n472 B.t3 52.36
R638 B.t0 B.n195 37.916
R639 B.t1 B.n8 37.916
R640 B.n460 B.n31 33.5615
R641 B.n455 B.n454 33.5615
R642 B.n384 B.n383 33.5615
R643 B.n388 B.n220 33.5615
R644 B.n326 B.n325 26.5702
R645 B.n243 B.n242 26.5702
R646 B.n70 B.n69 26.5702
R647 B.n67 B.n66 26.5702
R648 B.n424 B.t0 23.472
R649 B.n482 B.t1 23.472
R650 B B.n492 18.0485
R651 B.n71 B.n31 10.6151
R652 B.n74 B.n71 10.6151
R653 B.n75 B.n74 10.6151
R654 B.n78 B.n75 10.6151
R655 B.n79 B.n78 10.6151
R656 B.n82 B.n79 10.6151
R657 B.n83 B.n82 10.6151
R658 B.n86 B.n83 10.6151
R659 B.n87 B.n86 10.6151
R660 B.n90 B.n87 10.6151
R661 B.n91 B.n90 10.6151
R662 B.n94 B.n91 10.6151
R663 B.n95 B.n94 10.6151
R664 B.n98 B.n95 10.6151
R665 B.n99 B.n98 10.6151
R666 B.n102 B.n99 10.6151
R667 B.n103 B.n102 10.6151
R668 B.n106 B.n103 10.6151
R669 B.n107 B.n106 10.6151
R670 B.n110 B.n107 10.6151
R671 B.n111 B.n110 10.6151
R672 B.n114 B.n111 10.6151
R673 B.n115 B.n114 10.6151
R674 B.n118 B.n115 10.6151
R675 B.n119 B.n118 10.6151
R676 B.n122 B.n119 10.6151
R677 B.n127 B.n124 10.6151
R678 B.n128 B.n127 10.6151
R679 B.n131 B.n128 10.6151
R680 B.n132 B.n131 10.6151
R681 B.n135 B.n132 10.6151
R682 B.n136 B.n135 10.6151
R683 B.n139 B.n136 10.6151
R684 B.n140 B.n139 10.6151
R685 B.n144 B.n143 10.6151
R686 B.n147 B.n144 10.6151
R687 B.n148 B.n147 10.6151
R688 B.n151 B.n148 10.6151
R689 B.n152 B.n151 10.6151
R690 B.n155 B.n152 10.6151
R691 B.n156 B.n155 10.6151
R692 B.n159 B.n156 10.6151
R693 B.n160 B.n159 10.6151
R694 B.n163 B.n160 10.6151
R695 B.n164 B.n163 10.6151
R696 B.n167 B.n164 10.6151
R697 B.n168 B.n167 10.6151
R698 B.n171 B.n168 10.6151
R699 B.n172 B.n171 10.6151
R700 B.n175 B.n172 10.6151
R701 B.n176 B.n175 10.6151
R702 B.n179 B.n176 10.6151
R703 B.n180 B.n179 10.6151
R704 B.n183 B.n180 10.6151
R705 B.n184 B.n183 10.6151
R706 B.n187 B.n184 10.6151
R707 B.n188 B.n187 10.6151
R708 B.n191 B.n188 10.6151
R709 B.n192 B.n191 10.6151
R710 B.n455 B.n192 10.6151
R711 B.n384 B.n216 10.6151
R712 B.n394 B.n216 10.6151
R713 B.n395 B.n394 10.6151
R714 B.n396 B.n395 10.6151
R715 B.n396 B.n209 10.6151
R716 B.n407 B.n209 10.6151
R717 B.n408 B.n407 10.6151
R718 B.n409 B.n408 10.6151
R719 B.n409 B.n201 10.6151
R720 B.n419 B.n201 10.6151
R721 B.n420 B.n419 10.6151
R722 B.n422 B.n420 10.6151
R723 B.n422 B.n421 10.6151
R724 B.n421 B.n193 10.6151
R725 B.n433 B.n193 10.6151
R726 B.n434 B.n433 10.6151
R727 B.n435 B.n434 10.6151
R728 B.n436 B.n435 10.6151
R729 B.n438 B.n436 10.6151
R730 B.n439 B.n438 10.6151
R731 B.n440 B.n439 10.6151
R732 B.n441 B.n440 10.6151
R733 B.n443 B.n441 10.6151
R734 B.n444 B.n443 10.6151
R735 B.n445 B.n444 10.6151
R736 B.n446 B.n445 10.6151
R737 B.n448 B.n446 10.6151
R738 B.n449 B.n448 10.6151
R739 B.n450 B.n449 10.6151
R740 B.n451 B.n450 10.6151
R741 B.n453 B.n451 10.6151
R742 B.n454 B.n453 10.6151
R743 B.n258 B.n220 10.6151
R744 B.n259 B.n258 10.6151
R745 B.n260 B.n259 10.6151
R746 B.n260 B.n254 10.6151
R747 B.n266 B.n254 10.6151
R748 B.n267 B.n266 10.6151
R749 B.n268 B.n267 10.6151
R750 B.n268 B.n252 10.6151
R751 B.n274 B.n252 10.6151
R752 B.n275 B.n274 10.6151
R753 B.n276 B.n275 10.6151
R754 B.n276 B.n250 10.6151
R755 B.n282 B.n250 10.6151
R756 B.n283 B.n282 10.6151
R757 B.n284 B.n283 10.6151
R758 B.n284 B.n248 10.6151
R759 B.n290 B.n248 10.6151
R760 B.n291 B.n290 10.6151
R761 B.n292 B.n291 10.6151
R762 B.n292 B.n246 10.6151
R763 B.n298 B.n246 10.6151
R764 B.n299 B.n298 10.6151
R765 B.n300 B.n299 10.6151
R766 B.n300 B.n244 10.6151
R767 B.n306 B.n244 10.6151
R768 B.n307 B.n306 10.6151
R769 B.n309 B.n240 10.6151
R770 B.n315 B.n240 10.6151
R771 B.n316 B.n315 10.6151
R772 B.n317 B.n316 10.6151
R773 B.n317 B.n238 10.6151
R774 B.n323 B.n238 10.6151
R775 B.n324 B.n323 10.6151
R776 B.n328 B.n324 10.6151
R777 B.n334 B.n236 10.6151
R778 B.n335 B.n334 10.6151
R779 B.n336 B.n335 10.6151
R780 B.n336 B.n234 10.6151
R781 B.n342 B.n234 10.6151
R782 B.n343 B.n342 10.6151
R783 B.n344 B.n343 10.6151
R784 B.n344 B.n232 10.6151
R785 B.n350 B.n232 10.6151
R786 B.n351 B.n350 10.6151
R787 B.n352 B.n351 10.6151
R788 B.n352 B.n230 10.6151
R789 B.n358 B.n230 10.6151
R790 B.n359 B.n358 10.6151
R791 B.n360 B.n359 10.6151
R792 B.n360 B.n228 10.6151
R793 B.n366 B.n228 10.6151
R794 B.n367 B.n366 10.6151
R795 B.n368 B.n367 10.6151
R796 B.n368 B.n226 10.6151
R797 B.n374 B.n226 10.6151
R798 B.n375 B.n374 10.6151
R799 B.n376 B.n375 10.6151
R800 B.n376 B.n224 10.6151
R801 B.n382 B.n224 10.6151
R802 B.n383 B.n382 10.6151
R803 B.n389 B.n388 10.6151
R804 B.n390 B.n389 10.6151
R805 B.n390 B.n212 10.6151
R806 B.n401 B.n212 10.6151
R807 B.n402 B.n401 10.6151
R808 B.n403 B.n402 10.6151
R809 B.n403 B.n205 10.6151
R810 B.n413 B.n205 10.6151
R811 B.n414 B.n413 10.6151
R812 B.n415 B.n414 10.6151
R813 B.n415 B.n197 10.6151
R814 B.n426 B.n197 10.6151
R815 B.n427 B.n426 10.6151
R816 B.n428 B.n427 10.6151
R817 B.n428 B.n0 10.6151
R818 B.n486 B.n1 10.6151
R819 B.n486 B.n485 10.6151
R820 B.n485 B.n484 10.6151
R821 B.n484 B.n10 10.6151
R822 B.n478 B.n10 10.6151
R823 B.n478 B.n477 10.6151
R824 B.n477 B.n476 10.6151
R825 B.n476 B.n17 10.6151
R826 B.n470 B.n17 10.6151
R827 B.n470 B.n469 10.6151
R828 B.n469 B.n468 10.6151
R829 B.n468 B.n23 10.6151
R830 B.n462 B.n23 10.6151
R831 B.n462 B.n461 10.6151
R832 B.n461 B.n460 10.6151
R833 B.n398 B.t10 9.02799
R834 B.n25 B.t3 9.02799
R835 B.n124 B.n123 7.18099
R836 B.n140 B.n68 7.18099
R837 B.n309 B.n308 7.18099
R838 B.n328 B.n327 7.18099
R839 B.n123 B.n122 3.43465
R840 B.n143 B.n68 3.43465
R841 B.n308 B.n307 3.43465
R842 B.n327 B.n236 3.43465
R843 B.n492 B.n0 2.81026
R844 B.n492 B.n1 2.81026
R845 VP.n0 VP.t1 395.63
R846 VP.n0 VP.t0 358.966
R847 VP VP.n0 0.0516364
R848 VDD1 VDD1.t1 103.989
R849 VDD1 VDD1.t0 71.5439
C0 VDD2 VTAIL 3.64005f
C1 VDD1 VN 0.148744f
C2 VP VTAIL 1.22618f
C3 VDD2 VDD1 0.495088f
C4 VDD2 VN 1.39956f
C5 VP VDD1 1.51696f
C6 VP VN 3.76898f
C7 VDD1 VTAIL 3.60038f
C8 VTAIL VN 1.21184f
C9 VDD2 VP 0.268456f
C10 VDD2 B 2.941929f
C11 VDD1 B 4.66763f
C12 VTAIL B 4.462699f
C13 VN B 6.33309f
C14 VP B 4.030796f
C15 VDD1.t0 B 0.863178f
C16 VDD1.t1 B 1.10765f
C17 VP.t1 B 0.851207f
C18 VP.t0 B 0.745616f
C19 VP.n0 B 2.18635f
C20 VDD2.t0 B 1.10823f
C21 VDD2.t1 B 0.875439f
C22 VDD2.n0 B 1.57089f
C23 VTAIL.t0 B 0.920393f
C24 VTAIL.n0 B 0.898287f
C25 VTAIL.t2 B 0.920401f
C26 VTAIL.n1 B 0.910808f
C27 VTAIL.t1 B 0.920393f
C28 VTAIL.n2 B 0.848398f
C29 VTAIL.t3 B 0.920393f
C30 VTAIL.n3 B 0.804888f
C31 VN.t1 B 0.737416f
C32 VN.t0 B 0.844647f
.ends

