* NGSPICE file created from diff_pair_sample_0060.ext - technology: sky130A

.subckt diff_pair_sample_0060 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=2.26545 pd=14.06 as=2.26545 ps=14.06 w=13.73 l=3.97
X1 VTAIL.t2 VP.t0 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.26545 pd=14.06 as=2.26545 ps=14.06 w=13.73 l=3.97
X2 VDD1.t4 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.3547 pd=28.24 as=2.26545 ps=14.06 w=13.73 l=3.97
X3 VDD2.t3 VN.t1 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=5.3547 pd=28.24 as=2.26545 ps=14.06 w=13.73 l=3.97
X4 VDD1.t3 VP.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.26545 pd=14.06 as=5.3547 ps=28.24 w=13.73 l=3.97
X5 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=5.3547 pd=28.24 as=0 ps=0 w=13.73 l=3.97
X6 VTAIL.t9 VN.t2 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.26545 pd=14.06 as=2.26545 ps=14.06 w=13.73 l=3.97
X7 VDD2.t5 VN.t3 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=2.26545 pd=14.06 as=5.3547 ps=28.24 w=13.73 l=3.97
X8 VDD2.t4 VN.t4 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=5.3547 pd=28.24 as=2.26545 ps=14.06 w=13.73 l=3.97
X9 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=5.3547 pd=28.24 as=0 ps=0 w=13.73 l=3.97
X10 VDD2.t1 VN.t5 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.26545 pd=14.06 as=5.3547 ps=28.24 w=13.73 l=3.97
X11 VDD1.t2 VP.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=5.3547 pd=28.24 as=2.26545 ps=14.06 w=13.73 l=3.97
X12 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.3547 pd=28.24 as=0 ps=0 w=13.73 l=3.97
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.3547 pd=28.24 as=0 ps=0 w=13.73 l=3.97
X14 VTAIL.t5 VP.t4 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=2.26545 pd=14.06 as=2.26545 ps=14.06 w=13.73 l=3.97
X15 VDD1.t0 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.26545 pd=14.06 as=5.3547 ps=28.24 w=13.73 l=3.97
R0 VN.n42 VN.n41 161.3
R1 VN.n40 VN.n23 161.3
R2 VN.n39 VN.n38 161.3
R3 VN.n37 VN.n24 161.3
R4 VN.n36 VN.n35 161.3
R5 VN.n34 VN.n25 161.3
R6 VN.n33 VN.n32 161.3
R7 VN.n31 VN.n26 161.3
R8 VN.n30 VN.n29 161.3
R9 VN.n20 VN.n19 161.3
R10 VN.n18 VN.n1 161.3
R11 VN.n17 VN.n16 161.3
R12 VN.n15 VN.n2 161.3
R13 VN.n14 VN.n13 161.3
R14 VN.n12 VN.n3 161.3
R15 VN.n11 VN.n10 161.3
R16 VN.n9 VN.n4 161.3
R17 VN.n8 VN.n7 161.3
R18 VN.n27 VN.t5 116.038
R19 VN.n5 VN.t4 116.038
R20 VN.n21 VN.n0 87.6207
R21 VN.n43 VN.n22 87.6207
R22 VN.n6 VN.t2 83.3489
R23 VN.n0 VN.t3 83.3489
R24 VN.n28 VN.t0 83.3489
R25 VN.n22 VN.t1 83.3489
R26 VN.n28 VN.n27 62.9379
R27 VN.n6 VN.n5 62.9379
R28 VN VN.n43 55.6117
R29 VN.n13 VN.n12 50.2061
R30 VN.n35 VN.n34 50.2061
R31 VN.n13 VN.n2 30.7807
R32 VN.n35 VN.n24 30.7807
R33 VN.n7 VN.n4 24.4675
R34 VN.n11 VN.n4 24.4675
R35 VN.n12 VN.n11 24.4675
R36 VN.n17 VN.n2 24.4675
R37 VN.n18 VN.n17 24.4675
R38 VN.n19 VN.n18 24.4675
R39 VN.n34 VN.n33 24.4675
R40 VN.n33 VN.n26 24.4675
R41 VN.n29 VN.n26 24.4675
R42 VN.n41 VN.n40 24.4675
R43 VN.n40 VN.n39 24.4675
R44 VN.n39 VN.n24 24.4675
R45 VN.n7 VN.n6 12.234
R46 VN.n29 VN.n28 12.234
R47 VN.n30 VN.n27 2.47757
R48 VN.n8 VN.n5 2.47757
R49 VN.n19 VN.n0 2.4472
R50 VN.n41 VN.n22 2.4472
R51 VN.n43 VN.n42 0.354971
R52 VN.n21 VN.n20 0.354971
R53 VN VN.n21 0.26696
R54 VN.n42 VN.n23 0.189894
R55 VN.n38 VN.n23 0.189894
R56 VN.n38 VN.n37 0.189894
R57 VN.n37 VN.n36 0.189894
R58 VN.n36 VN.n25 0.189894
R59 VN.n32 VN.n25 0.189894
R60 VN.n32 VN.n31 0.189894
R61 VN.n31 VN.n30 0.189894
R62 VN.n9 VN.n8 0.189894
R63 VN.n10 VN.n9 0.189894
R64 VN.n10 VN.n3 0.189894
R65 VN.n14 VN.n3 0.189894
R66 VN.n15 VN.n14 0.189894
R67 VN.n16 VN.n15 0.189894
R68 VN.n16 VN.n1 0.189894
R69 VN.n20 VN.n1 0.189894
R70 VDD2.n1 VDD2.t4 68.5308
R71 VDD2.n2 VDD2.t3 65.8062
R72 VDD2.n1 VDD2.n0 65.2353
R73 VDD2 VDD2.n3 65.2325
R74 VDD2.n2 VDD2.n1 47.5989
R75 VDD2 VDD2.n2 2.83886
R76 VDD2.n3 VDD2.t2 1.4426
R77 VDD2.n3 VDD2.t1 1.4426
R78 VDD2.n0 VDD2.t0 1.4426
R79 VDD2.n0 VDD2.t5 1.4426
R80 VTAIL.n7 VTAIL.t6 49.1274
R81 VTAIL.n11 VTAIL.t8 49.1272
R82 VTAIL.n2 VTAIL.t3 49.1272
R83 VTAIL.n10 VTAIL.t0 49.1272
R84 VTAIL.n9 VTAIL.n8 47.6853
R85 VTAIL.n6 VTAIL.n5 47.6853
R86 VTAIL.n1 VTAIL.n0 47.6851
R87 VTAIL.n4 VTAIL.n3 47.6851
R88 VTAIL.n6 VTAIL.n4 31.6169
R89 VTAIL.n11 VTAIL.n10 27.91
R90 VTAIL.n7 VTAIL.n6 3.7074
R91 VTAIL.n10 VTAIL.n9 3.7074
R92 VTAIL.n4 VTAIL.n2 3.7074
R93 VTAIL VTAIL.n11 2.72248
R94 VTAIL.n9 VTAIL.n7 2.32378
R95 VTAIL.n2 VTAIL.n1 2.32378
R96 VTAIL.n0 VTAIL.t7 1.4426
R97 VTAIL.n0 VTAIL.t9 1.4426
R98 VTAIL.n3 VTAIL.t4 1.4426
R99 VTAIL.n3 VTAIL.t5 1.4426
R100 VTAIL.n8 VTAIL.t1 1.4426
R101 VTAIL.n8 VTAIL.t2 1.4426
R102 VTAIL.n5 VTAIL.t10 1.4426
R103 VTAIL.n5 VTAIL.t11 1.4426
R104 VTAIL VTAIL.n1 0.985414
R105 B.n791 B.n790 585
R106 B.n791 B.n107 585
R107 B.n794 B.n793 585
R108 B.n795 B.n163 585
R109 B.n797 B.n796 585
R110 B.n799 B.n162 585
R111 B.n802 B.n801 585
R112 B.n803 B.n161 585
R113 B.n805 B.n804 585
R114 B.n807 B.n160 585
R115 B.n810 B.n809 585
R116 B.n811 B.n159 585
R117 B.n813 B.n812 585
R118 B.n815 B.n158 585
R119 B.n818 B.n817 585
R120 B.n819 B.n157 585
R121 B.n821 B.n820 585
R122 B.n823 B.n156 585
R123 B.n826 B.n825 585
R124 B.n827 B.n155 585
R125 B.n829 B.n828 585
R126 B.n831 B.n154 585
R127 B.n834 B.n833 585
R128 B.n835 B.n153 585
R129 B.n837 B.n836 585
R130 B.n839 B.n152 585
R131 B.n842 B.n841 585
R132 B.n843 B.n151 585
R133 B.n845 B.n844 585
R134 B.n847 B.n150 585
R135 B.n850 B.n849 585
R136 B.n851 B.n149 585
R137 B.n853 B.n852 585
R138 B.n855 B.n148 585
R139 B.n858 B.n857 585
R140 B.n859 B.n147 585
R141 B.n861 B.n860 585
R142 B.n863 B.n146 585
R143 B.n866 B.n865 585
R144 B.n867 B.n145 585
R145 B.n869 B.n868 585
R146 B.n871 B.n144 585
R147 B.n874 B.n873 585
R148 B.n875 B.n143 585
R149 B.n877 B.n876 585
R150 B.n879 B.n142 585
R151 B.n882 B.n881 585
R152 B.n883 B.n139 585
R153 B.n886 B.n885 585
R154 B.n888 B.n138 585
R155 B.n891 B.n890 585
R156 B.n892 B.n137 585
R157 B.n894 B.n893 585
R158 B.n896 B.n136 585
R159 B.n899 B.n898 585
R160 B.n900 B.n132 585
R161 B.n902 B.n901 585
R162 B.n904 B.n131 585
R163 B.n907 B.n906 585
R164 B.n908 B.n130 585
R165 B.n910 B.n909 585
R166 B.n912 B.n129 585
R167 B.n915 B.n914 585
R168 B.n916 B.n128 585
R169 B.n918 B.n917 585
R170 B.n920 B.n127 585
R171 B.n923 B.n922 585
R172 B.n924 B.n126 585
R173 B.n926 B.n925 585
R174 B.n928 B.n125 585
R175 B.n931 B.n930 585
R176 B.n932 B.n124 585
R177 B.n934 B.n933 585
R178 B.n936 B.n123 585
R179 B.n939 B.n938 585
R180 B.n940 B.n122 585
R181 B.n942 B.n941 585
R182 B.n944 B.n121 585
R183 B.n947 B.n946 585
R184 B.n948 B.n120 585
R185 B.n950 B.n949 585
R186 B.n952 B.n119 585
R187 B.n955 B.n954 585
R188 B.n956 B.n118 585
R189 B.n958 B.n957 585
R190 B.n960 B.n117 585
R191 B.n963 B.n962 585
R192 B.n964 B.n116 585
R193 B.n966 B.n965 585
R194 B.n968 B.n115 585
R195 B.n971 B.n970 585
R196 B.n972 B.n114 585
R197 B.n974 B.n973 585
R198 B.n976 B.n113 585
R199 B.n979 B.n978 585
R200 B.n980 B.n112 585
R201 B.n982 B.n981 585
R202 B.n984 B.n111 585
R203 B.n987 B.n986 585
R204 B.n988 B.n110 585
R205 B.n990 B.n989 585
R206 B.n992 B.n109 585
R207 B.n995 B.n994 585
R208 B.n996 B.n108 585
R209 B.n789 B.n106 585
R210 B.n999 B.n106 585
R211 B.n788 B.n105 585
R212 B.n1000 B.n105 585
R213 B.n787 B.n104 585
R214 B.n1001 B.n104 585
R215 B.n786 B.n785 585
R216 B.n785 B.n100 585
R217 B.n784 B.n99 585
R218 B.n1007 B.n99 585
R219 B.n783 B.n98 585
R220 B.n1008 B.n98 585
R221 B.n782 B.n97 585
R222 B.n1009 B.n97 585
R223 B.n781 B.n780 585
R224 B.n780 B.n93 585
R225 B.n779 B.n92 585
R226 B.n1015 B.n92 585
R227 B.n778 B.n91 585
R228 B.n1016 B.n91 585
R229 B.n777 B.n90 585
R230 B.n1017 B.n90 585
R231 B.n776 B.n775 585
R232 B.n775 B.n86 585
R233 B.n774 B.n85 585
R234 B.n1023 B.n85 585
R235 B.n773 B.n84 585
R236 B.n1024 B.n84 585
R237 B.n772 B.n83 585
R238 B.n1025 B.n83 585
R239 B.n771 B.n770 585
R240 B.n770 B.n79 585
R241 B.n769 B.n78 585
R242 B.n1031 B.n78 585
R243 B.n768 B.n77 585
R244 B.n1032 B.n77 585
R245 B.n767 B.n76 585
R246 B.n1033 B.n76 585
R247 B.n766 B.n765 585
R248 B.n765 B.n72 585
R249 B.n764 B.n71 585
R250 B.n1039 B.n71 585
R251 B.n763 B.n70 585
R252 B.n1040 B.n70 585
R253 B.n762 B.n69 585
R254 B.n1041 B.n69 585
R255 B.n761 B.n760 585
R256 B.n760 B.n65 585
R257 B.n759 B.n64 585
R258 B.n1047 B.n64 585
R259 B.n758 B.n63 585
R260 B.n1048 B.n63 585
R261 B.n757 B.n62 585
R262 B.n1049 B.n62 585
R263 B.n756 B.n755 585
R264 B.n755 B.n58 585
R265 B.n754 B.n57 585
R266 B.n1055 B.n57 585
R267 B.n753 B.n56 585
R268 B.n1056 B.n56 585
R269 B.n752 B.n55 585
R270 B.n1057 B.n55 585
R271 B.n751 B.n750 585
R272 B.n750 B.n51 585
R273 B.n749 B.n50 585
R274 B.n1063 B.n50 585
R275 B.n748 B.n49 585
R276 B.n1064 B.n49 585
R277 B.n747 B.n48 585
R278 B.n1065 B.n48 585
R279 B.n746 B.n745 585
R280 B.n745 B.n44 585
R281 B.n744 B.n43 585
R282 B.n1071 B.n43 585
R283 B.n743 B.n42 585
R284 B.n1072 B.n42 585
R285 B.n742 B.n41 585
R286 B.n1073 B.n41 585
R287 B.n741 B.n740 585
R288 B.n740 B.n37 585
R289 B.n739 B.n36 585
R290 B.n1079 B.n36 585
R291 B.n738 B.n35 585
R292 B.n1080 B.n35 585
R293 B.n737 B.n34 585
R294 B.n1081 B.n34 585
R295 B.n736 B.n735 585
R296 B.n735 B.n30 585
R297 B.n734 B.n29 585
R298 B.n1087 B.n29 585
R299 B.n733 B.n28 585
R300 B.n1088 B.n28 585
R301 B.n732 B.n27 585
R302 B.n1089 B.n27 585
R303 B.n731 B.n730 585
R304 B.n730 B.n23 585
R305 B.n729 B.n22 585
R306 B.n1095 B.n22 585
R307 B.n728 B.n21 585
R308 B.n1096 B.n21 585
R309 B.n727 B.n20 585
R310 B.n1097 B.n20 585
R311 B.n726 B.n725 585
R312 B.n725 B.n16 585
R313 B.n724 B.n15 585
R314 B.n1103 B.n15 585
R315 B.n723 B.n14 585
R316 B.n1104 B.n14 585
R317 B.n722 B.n13 585
R318 B.n1105 B.n13 585
R319 B.n721 B.n720 585
R320 B.n720 B.n12 585
R321 B.n719 B.n718 585
R322 B.n719 B.n8 585
R323 B.n717 B.n7 585
R324 B.n1112 B.n7 585
R325 B.n716 B.n6 585
R326 B.n1113 B.n6 585
R327 B.n715 B.n5 585
R328 B.n1114 B.n5 585
R329 B.n714 B.n713 585
R330 B.n713 B.n4 585
R331 B.n712 B.n164 585
R332 B.n712 B.n711 585
R333 B.n702 B.n165 585
R334 B.n166 B.n165 585
R335 B.n704 B.n703 585
R336 B.n705 B.n704 585
R337 B.n701 B.n171 585
R338 B.n171 B.n170 585
R339 B.n700 B.n699 585
R340 B.n699 B.n698 585
R341 B.n173 B.n172 585
R342 B.n174 B.n173 585
R343 B.n691 B.n690 585
R344 B.n692 B.n691 585
R345 B.n689 B.n179 585
R346 B.n179 B.n178 585
R347 B.n688 B.n687 585
R348 B.n687 B.n686 585
R349 B.n181 B.n180 585
R350 B.n182 B.n181 585
R351 B.n679 B.n678 585
R352 B.n680 B.n679 585
R353 B.n677 B.n187 585
R354 B.n187 B.n186 585
R355 B.n676 B.n675 585
R356 B.n675 B.n674 585
R357 B.n189 B.n188 585
R358 B.n190 B.n189 585
R359 B.n667 B.n666 585
R360 B.n668 B.n667 585
R361 B.n665 B.n195 585
R362 B.n195 B.n194 585
R363 B.n664 B.n663 585
R364 B.n663 B.n662 585
R365 B.n197 B.n196 585
R366 B.n198 B.n197 585
R367 B.n655 B.n654 585
R368 B.n656 B.n655 585
R369 B.n653 B.n202 585
R370 B.n206 B.n202 585
R371 B.n652 B.n651 585
R372 B.n651 B.n650 585
R373 B.n204 B.n203 585
R374 B.n205 B.n204 585
R375 B.n643 B.n642 585
R376 B.n644 B.n643 585
R377 B.n641 B.n211 585
R378 B.n211 B.n210 585
R379 B.n640 B.n639 585
R380 B.n639 B.n638 585
R381 B.n213 B.n212 585
R382 B.n214 B.n213 585
R383 B.n631 B.n630 585
R384 B.n632 B.n631 585
R385 B.n629 B.n219 585
R386 B.n219 B.n218 585
R387 B.n628 B.n627 585
R388 B.n627 B.n626 585
R389 B.n221 B.n220 585
R390 B.n222 B.n221 585
R391 B.n619 B.n618 585
R392 B.n620 B.n619 585
R393 B.n617 B.n226 585
R394 B.n230 B.n226 585
R395 B.n616 B.n615 585
R396 B.n615 B.n614 585
R397 B.n228 B.n227 585
R398 B.n229 B.n228 585
R399 B.n607 B.n606 585
R400 B.n608 B.n607 585
R401 B.n605 B.n235 585
R402 B.n235 B.n234 585
R403 B.n604 B.n603 585
R404 B.n603 B.n602 585
R405 B.n237 B.n236 585
R406 B.n238 B.n237 585
R407 B.n595 B.n594 585
R408 B.n596 B.n595 585
R409 B.n593 B.n243 585
R410 B.n243 B.n242 585
R411 B.n592 B.n591 585
R412 B.n591 B.n590 585
R413 B.n245 B.n244 585
R414 B.n246 B.n245 585
R415 B.n583 B.n582 585
R416 B.n584 B.n583 585
R417 B.n581 B.n251 585
R418 B.n251 B.n250 585
R419 B.n580 B.n579 585
R420 B.n579 B.n578 585
R421 B.n253 B.n252 585
R422 B.n254 B.n253 585
R423 B.n571 B.n570 585
R424 B.n572 B.n571 585
R425 B.n569 B.n258 585
R426 B.n262 B.n258 585
R427 B.n568 B.n567 585
R428 B.n567 B.n566 585
R429 B.n260 B.n259 585
R430 B.n261 B.n260 585
R431 B.n559 B.n558 585
R432 B.n560 B.n559 585
R433 B.n557 B.n267 585
R434 B.n267 B.n266 585
R435 B.n556 B.n555 585
R436 B.n555 B.n554 585
R437 B.n269 B.n268 585
R438 B.n270 B.n269 585
R439 B.n547 B.n546 585
R440 B.n548 B.n547 585
R441 B.n545 B.n275 585
R442 B.n275 B.n274 585
R443 B.n544 B.n543 585
R444 B.n543 B.n542 585
R445 B.n539 B.n279 585
R446 B.n538 B.n537 585
R447 B.n535 B.n280 585
R448 B.n535 B.n278 585
R449 B.n534 B.n533 585
R450 B.n532 B.n531 585
R451 B.n530 B.n282 585
R452 B.n528 B.n527 585
R453 B.n526 B.n283 585
R454 B.n525 B.n524 585
R455 B.n522 B.n284 585
R456 B.n520 B.n519 585
R457 B.n518 B.n285 585
R458 B.n517 B.n516 585
R459 B.n514 B.n286 585
R460 B.n512 B.n511 585
R461 B.n510 B.n287 585
R462 B.n509 B.n508 585
R463 B.n506 B.n288 585
R464 B.n504 B.n503 585
R465 B.n502 B.n289 585
R466 B.n501 B.n500 585
R467 B.n498 B.n290 585
R468 B.n496 B.n495 585
R469 B.n494 B.n291 585
R470 B.n493 B.n492 585
R471 B.n490 B.n292 585
R472 B.n488 B.n487 585
R473 B.n486 B.n293 585
R474 B.n485 B.n484 585
R475 B.n482 B.n294 585
R476 B.n480 B.n479 585
R477 B.n478 B.n295 585
R478 B.n477 B.n476 585
R479 B.n474 B.n296 585
R480 B.n472 B.n471 585
R481 B.n470 B.n297 585
R482 B.n469 B.n468 585
R483 B.n466 B.n298 585
R484 B.n464 B.n463 585
R485 B.n462 B.n299 585
R486 B.n461 B.n460 585
R487 B.n458 B.n300 585
R488 B.n456 B.n455 585
R489 B.n454 B.n301 585
R490 B.n453 B.n452 585
R491 B.n450 B.n302 585
R492 B.n448 B.n447 585
R493 B.n445 B.n303 585
R494 B.n444 B.n443 585
R495 B.n441 B.n306 585
R496 B.n439 B.n438 585
R497 B.n437 B.n307 585
R498 B.n436 B.n435 585
R499 B.n433 B.n308 585
R500 B.n431 B.n430 585
R501 B.n429 B.n309 585
R502 B.n427 B.n426 585
R503 B.n424 B.n312 585
R504 B.n422 B.n421 585
R505 B.n420 B.n313 585
R506 B.n419 B.n418 585
R507 B.n416 B.n314 585
R508 B.n414 B.n413 585
R509 B.n412 B.n315 585
R510 B.n411 B.n410 585
R511 B.n408 B.n316 585
R512 B.n406 B.n405 585
R513 B.n404 B.n317 585
R514 B.n403 B.n402 585
R515 B.n400 B.n318 585
R516 B.n398 B.n397 585
R517 B.n396 B.n319 585
R518 B.n395 B.n394 585
R519 B.n392 B.n320 585
R520 B.n390 B.n389 585
R521 B.n388 B.n321 585
R522 B.n387 B.n386 585
R523 B.n384 B.n322 585
R524 B.n382 B.n381 585
R525 B.n380 B.n323 585
R526 B.n379 B.n378 585
R527 B.n376 B.n324 585
R528 B.n374 B.n373 585
R529 B.n372 B.n325 585
R530 B.n371 B.n370 585
R531 B.n368 B.n326 585
R532 B.n366 B.n365 585
R533 B.n364 B.n327 585
R534 B.n363 B.n362 585
R535 B.n360 B.n328 585
R536 B.n358 B.n357 585
R537 B.n356 B.n329 585
R538 B.n355 B.n354 585
R539 B.n352 B.n330 585
R540 B.n350 B.n349 585
R541 B.n348 B.n331 585
R542 B.n347 B.n346 585
R543 B.n344 B.n332 585
R544 B.n342 B.n341 585
R545 B.n340 B.n333 585
R546 B.n339 B.n338 585
R547 B.n336 B.n334 585
R548 B.n277 B.n276 585
R549 B.n541 B.n540 585
R550 B.n542 B.n541 585
R551 B.n273 B.n272 585
R552 B.n274 B.n273 585
R553 B.n550 B.n549 585
R554 B.n549 B.n548 585
R555 B.n551 B.n271 585
R556 B.n271 B.n270 585
R557 B.n553 B.n552 585
R558 B.n554 B.n553 585
R559 B.n265 B.n264 585
R560 B.n266 B.n265 585
R561 B.n562 B.n561 585
R562 B.n561 B.n560 585
R563 B.n563 B.n263 585
R564 B.n263 B.n261 585
R565 B.n565 B.n564 585
R566 B.n566 B.n565 585
R567 B.n257 B.n256 585
R568 B.n262 B.n257 585
R569 B.n574 B.n573 585
R570 B.n573 B.n572 585
R571 B.n575 B.n255 585
R572 B.n255 B.n254 585
R573 B.n577 B.n576 585
R574 B.n578 B.n577 585
R575 B.n249 B.n248 585
R576 B.n250 B.n249 585
R577 B.n586 B.n585 585
R578 B.n585 B.n584 585
R579 B.n587 B.n247 585
R580 B.n247 B.n246 585
R581 B.n589 B.n588 585
R582 B.n590 B.n589 585
R583 B.n241 B.n240 585
R584 B.n242 B.n241 585
R585 B.n598 B.n597 585
R586 B.n597 B.n596 585
R587 B.n599 B.n239 585
R588 B.n239 B.n238 585
R589 B.n601 B.n600 585
R590 B.n602 B.n601 585
R591 B.n233 B.n232 585
R592 B.n234 B.n233 585
R593 B.n610 B.n609 585
R594 B.n609 B.n608 585
R595 B.n611 B.n231 585
R596 B.n231 B.n229 585
R597 B.n613 B.n612 585
R598 B.n614 B.n613 585
R599 B.n225 B.n224 585
R600 B.n230 B.n225 585
R601 B.n622 B.n621 585
R602 B.n621 B.n620 585
R603 B.n623 B.n223 585
R604 B.n223 B.n222 585
R605 B.n625 B.n624 585
R606 B.n626 B.n625 585
R607 B.n217 B.n216 585
R608 B.n218 B.n217 585
R609 B.n634 B.n633 585
R610 B.n633 B.n632 585
R611 B.n635 B.n215 585
R612 B.n215 B.n214 585
R613 B.n637 B.n636 585
R614 B.n638 B.n637 585
R615 B.n209 B.n208 585
R616 B.n210 B.n209 585
R617 B.n646 B.n645 585
R618 B.n645 B.n644 585
R619 B.n647 B.n207 585
R620 B.n207 B.n205 585
R621 B.n649 B.n648 585
R622 B.n650 B.n649 585
R623 B.n201 B.n200 585
R624 B.n206 B.n201 585
R625 B.n658 B.n657 585
R626 B.n657 B.n656 585
R627 B.n659 B.n199 585
R628 B.n199 B.n198 585
R629 B.n661 B.n660 585
R630 B.n662 B.n661 585
R631 B.n193 B.n192 585
R632 B.n194 B.n193 585
R633 B.n670 B.n669 585
R634 B.n669 B.n668 585
R635 B.n671 B.n191 585
R636 B.n191 B.n190 585
R637 B.n673 B.n672 585
R638 B.n674 B.n673 585
R639 B.n185 B.n184 585
R640 B.n186 B.n185 585
R641 B.n682 B.n681 585
R642 B.n681 B.n680 585
R643 B.n683 B.n183 585
R644 B.n183 B.n182 585
R645 B.n685 B.n684 585
R646 B.n686 B.n685 585
R647 B.n177 B.n176 585
R648 B.n178 B.n177 585
R649 B.n694 B.n693 585
R650 B.n693 B.n692 585
R651 B.n695 B.n175 585
R652 B.n175 B.n174 585
R653 B.n697 B.n696 585
R654 B.n698 B.n697 585
R655 B.n169 B.n168 585
R656 B.n170 B.n169 585
R657 B.n707 B.n706 585
R658 B.n706 B.n705 585
R659 B.n708 B.n167 585
R660 B.n167 B.n166 585
R661 B.n710 B.n709 585
R662 B.n711 B.n710 585
R663 B.n3 B.n0 585
R664 B.n4 B.n3 585
R665 B.n1111 B.n1 585
R666 B.n1112 B.n1111 585
R667 B.n1110 B.n1109 585
R668 B.n1110 B.n8 585
R669 B.n1108 B.n9 585
R670 B.n12 B.n9 585
R671 B.n1107 B.n1106 585
R672 B.n1106 B.n1105 585
R673 B.n11 B.n10 585
R674 B.n1104 B.n11 585
R675 B.n1102 B.n1101 585
R676 B.n1103 B.n1102 585
R677 B.n1100 B.n17 585
R678 B.n17 B.n16 585
R679 B.n1099 B.n1098 585
R680 B.n1098 B.n1097 585
R681 B.n19 B.n18 585
R682 B.n1096 B.n19 585
R683 B.n1094 B.n1093 585
R684 B.n1095 B.n1094 585
R685 B.n1092 B.n24 585
R686 B.n24 B.n23 585
R687 B.n1091 B.n1090 585
R688 B.n1090 B.n1089 585
R689 B.n26 B.n25 585
R690 B.n1088 B.n26 585
R691 B.n1086 B.n1085 585
R692 B.n1087 B.n1086 585
R693 B.n1084 B.n31 585
R694 B.n31 B.n30 585
R695 B.n1083 B.n1082 585
R696 B.n1082 B.n1081 585
R697 B.n33 B.n32 585
R698 B.n1080 B.n33 585
R699 B.n1078 B.n1077 585
R700 B.n1079 B.n1078 585
R701 B.n1076 B.n38 585
R702 B.n38 B.n37 585
R703 B.n1075 B.n1074 585
R704 B.n1074 B.n1073 585
R705 B.n40 B.n39 585
R706 B.n1072 B.n40 585
R707 B.n1070 B.n1069 585
R708 B.n1071 B.n1070 585
R709 B.n1068 B.n45 585
R710 B.n45 B.n44 585
R711 B.n1067 B.n1066 585
R712 B.n1066 B.n1065 585
R713 B.n47 B.n46 585
R714 B.n1064 B.n47 585
R715 B.n1062 B.n1061 585
R716 B.n1063 B.n1062 585
R717 B.n1060 B.n52 585
R718 B.n52 B.n51 585
R719 B.n1059 B.n1058 585
R720 B.n1058 B.n1057 585
R721 B.n54 B.n53 585
R722 B.n1056 B.n54 585
R723 B.n1054 B.n1053 585
R724 B.n1055 B.n1054 585
R725 B.n1052 B.n59 585
R726 B.n59 B.n58 585
R727 B.n1051 B.n1050 585
R728 B.n1050 B.n1049 585
R729 B.n61 B.n60 585
R730 B.n1048 B.n61 585
R731 B.n1046 B.n1045 585
R732 B.n1047 B.n1046 585
R733 B.n1044 B.n66 585
R734 B.n66 B.n65 585
R735 B.n1043 B.n1042 585
R736 B.n1042 B.n1041 585
R737 B.n68 B.n67 585
R738 B.n1040 B.n68 585
R739 B.n1038 B.n1037 585
R740 B.n1039 B.n1038 585
R741 B.n1036 B.n73 585
R742 B.n73 B.n72 585
R743 B.n1035 B.n1034 585
R744 B.n1034 B.n1033 585
R745 B.n75 B.n74 585
R746 B.n1032 B.n75 585
R747 B.n1030 B.n1029 585
R748 B.n1031 B.n1030 585
R749 B.n1028 B.n80 585
R750 B.n80 B.n79 585
R751 B.n1027 B.n1026 585
R752 B.n1026 B.n1025 585
R753 B.n82 B.n81 585
R754 B.n1024 B.n82 585
R755 B.n1022 B.n1021 585
R756 B.n1023 B.n1022 585
R757 B.n1020 B.n87 585
R758 B.n87 B.n86 585
R759 B.n1019 B.n1018 585
R760 B.n1018 B.n1017 585
R761 B.n89 B.n88 585
R762 B.n1016 B.n89 585
R763 B.n1014 B.n1013 585
R764 B.n1015 B.n1014 585
R765 B.n1012 B.n94 585
R766 B.n94 B.n93 585
R767 B.n1011 B.n1010 585
R768 B.n1010 B.n1009 585
R769 B.n96 B.n95 585
R770 B.n1008 B.n96 585
R771 B.n1006 B.n1005 585
R772 B.n1007 B.n1006 585
R773 B.n1004 B.n101 585
R774 B.n101 B.n100 585
R775 B.n1003 B.n1002 585
R776 B.n1002 B.n1001 585
R777 B.n103 B.n102 585
R778 B.n1000 B.n103 585
R779 B.n998 B.n997 585
R780 B.n999 B.n998 585
R781 B.n1115 B.n1114 585
R782 B.n1113 B.n2 585
R783 B.n998 B.n108 530.939
R784 B.n791 B.n106 530.939
R785 B.n543 B.n277 530.939
R786 B.n541 B.n279 530.939
R787 B.n133 B.t6 292.818
R788 B.n140 B.t17 292.818
R789 B.n310 B.t14 292.818
R790 B.n304 B.t10 292.818
R791 B.n792 B.n107 256.663
R792 B.n798 B.n107 256.663
R793 B.n800 B.n107 256.663
R794 B.n806 B.n107 256.663
R795 B.n808 B.n107 256.663
R796 B.n814 B.n107 256.663
R797 B.n816 B.n107 256.663
R798 B.n822 B.n107 256.663
R799 B.n824 B.n107 256.663
R800 B.n830 B.n107 256.663
R801 B.n832 B.n107 256.663
R802 B.n838 B.n107 256.663
R803 B.n840 B.n107 256.663
R804 B.n846 B.n107 256.663
R805 B.n848 B.n107 256.663
R806 B.n854 B.n107 256.663
R807 B.n856 B.n107 256.663
R808 B.n862 B.n107 256.663
R809 B.n864 B.n107 256.663
R810 B.n870 B.n107 256.663
R811 B.n872 B.n107 256.663
R812 B.n878 B.n107 256.663
R813 B.n880 B.n107 256.663
R814 B.n887 B.n107 256.663
R815 B.n889 B.n107 256.663
R816 B.n895 B.n107 256.663
R817 B.n897 B.n107 256.663
R818 B.n903 B.n107 256.663
R819 B.n905 B.n107 256.663
R820 B.n911 B.n107 256.663
R821 B.n913 B.n107 256.663
R822 B.n919 B.n107 256.663
R823 B.n921 B.n107 256.663
R824 B.n927 B.n107 256.663
R825 B.n929 B.n107 256.663
R826 B.n935 B.n107 256.663
R827 B.n937 B.n107 256.663
R828 B.n943 B.n107 256.663
R829 B.n945 B.n107 256.663
R830 B.n951 B.n107 256.663
R831 B.n953 B.n107 256.663
R832 B.n959 B.n107 256.663
R833 B.n961 B.n107 256.663
R834 B.n967 B.n107 256.663
R835 B.n969 B.n107 256.663
R836 B.n975 B.n107 256.663
R837 B.n977 B.n107 256.663
R838 B.n983 B.n107 256.663
R839 B.n985 B.n107 256.663
R840 B.n991 B.n107 256.663
R841 B.n993 B.n107 256.663
R842 B.n536 B.n278 256.663
R843 B.n281 B.n278 256.663
R844 B.n529 B.n278 256.663
R845 B.n523 B.n278 256.663
R846 B.n521 B.n278 256.663
R847 B.n515 B.n278 256.663
R848 B.n513 B.n278 256.663
R849 B.n507 B.n278 256.663
R850 B.n505 B.n278 256.663
R851 B.n499 B.n278 256.663
R852 B.n497 B.n278 256.663
R853 B.n491 B.n278 256.663
R854 B.n489 B.n278 256.663
R855 B.n483 B.n278 256.663
R856 B.n481 B.n278 256.663
R857 B.n475 B.n278 256.663
R858 B.n473 B.n278 256.663
R859 B.n467 B.n278 256.663
R860 B.n465 B.n278 256.663
R861 B.n459 B.n278 256.663
R862 B.n457 B.n278 256.663
R863 B.n451 B.n278 256.663
R864 B.n449 B.n278 256.663
R865 B.n442 B.n278 256.663
R866 B.n440 B.n278 256.663
R867 B.n434 B.n278 256.663
R868 B.n432 B.n278 256.663
R869 B.n425 B.n278 256.663
R870 B.n423 B.n278 256.663
R871 B.n417 B.n278 256.663
R872 B.n415 B.n278 256.663
R873 B.n409 B.n278 256.663
R874 B.n407 B.n278 256.663
R875 B.n401 B.n278 256.663
R876 B.n399 B.n278 256.663
R877 B.n393 B.n278 256.663
R878 B.n391 B.n278 256.663
R879 B.n385 B.n278 256.663
R880 B.n383 B.n278 256.663
R881 B.n377 B.n278 256.663
R882 B.n375 B.n278 256.663
R883 B.n369 B.n278 256.663
R884 B.n367 B.n278 256.663
R885 B.n361 B.n278 256.663
R886 B.n359 B.n278 256.663
R887 B.n353 B.n278 256.663
R888 B.n351 B.n278 256.663
R889 B.n345 B.n278 256.663
R890 B.n343 B.n278 256.663
R891 B.n337 B.n278 256.663
R892 B.n335 B.n278 256.663
R893 B.n1117 B.n1116 256.663
R894 B.n994 B.n992 163.367
R895 B.n990 B.n110 163.367
R896 B.n986 B.n984 163.367
R897 B.n982 B.n112 163.367
R898 B.n978 B.n976 163.367
R899 B.n974 B.n114 163.367
R900 B.n970 B.n968 163.367
R901 B.n966 B.n116 163.367
R902 B.n962 B.n960 163.367
R903 B.n958 B.n118 163.367
R904 B.n954 B.n952 163.367
R905 B.n950 B.n120 163.367
R906 B.n946 B.n944 163.367
R907 B.n942 B.n122 163.367
R908 B.n938 B.n936 163.367
R909 B.n934 B.n124 163.367
R910 B.n930 B.n928 163.367
R911 B.n926 B.n126 163.367
R912 B.n922 B.n920 163.367
R913 B.n918 B.n128 163.367
R914 B.n914 B.n912 163.367
R915 B.n910 B.n130 163.367
R916 B.n906 B.n904 163.367
R917 B.n902 B.n132 163.367
R918 B.n898 B.n896 163.367
R919 B.n894 B.n137 163.367
R920 B.n890 B.n888 163.367
R921 B.n886 B.n139 163.367
R922 B.n881 B.n879 163.367
R923 B.n877 B.n143 163.367
R924 B.n873 B.n871 163.367
R925 B.n869 B.n145 163.367
R926 B.n865 B.n863 163.367
R927 B.n861 B.n147 163.367
R928 B.n857 B.n855 163.367
R929 B.n853 B.n149 163.367
R930 B.n849 B.n847 163.367
R931 B.n845 B.n151 163.367
R932 B.n841 B.n839 163.367
R933 B.n837 B.n153 163.367
R934 B.n833 B.n831 163.367
R935 B.n829 B.n155 163.367
R936 B.n825 B.n823 163.367
R937 B.n821 B.n157 163.367
R938 B.n817 B.n815 163.367
R939 B.n813 B.n159 163.367
R940 B.n809 B.n807 163.367
R941 B.n805 B.n161 163.367
R942 B.n801 B.n799 163.367
R943 B.n797 B.n163 163.367
R944 B.n793 B.n791 163.367
R945 B.n543 B.n275 163.367
R946 B.n547 B.n275 163.367
R947 B.n547 B.n269 163.367
R948 B.n555 B.n269 163.367
R949 B.n555 B.n267 163.367
R950 B.n559 B.n267 163.367
R951 B.n559 B.n260 163.367
R952 B.n567 B.n260 163.367
R953 B.n567 B.n258 163.367
R954 B.n571 B.n258 163.367
R955 B.n571 B.n253 163.367
R956 B.n579 B.n253 163.367
R957 B.n579 B.n251 163.367
R958 B.n583 B.n251 163.367
R959 B.n583 B.n245 163.367
R960 B.n591 B.n245 163.367
R961 B.n591 B.n243 163.367
R962 B.n595 B.n243 163.367
R963 B.n595 B.n237 163.367
R964 B.n603 B.n237 163.367
R965 B.n603 B.n235 163.367
R966 B.n607 B.n235 163.367
R967 B.n607 B.n228 163.367
R968 B.n615 B.n228 163.367
R969 B.n615 B.n226 163.367
R970 B.n619 B.n226 163.367
R971 B.n619 B.n221 163.367
R972 B.n627 B.n221 163.367
R973 B.n627 B.n219 163.367
R974 B.n631 B.n219 163.367
R975 B.n631 B.n213 163.367
R976 B.n639 B.n213 163.367
R977 B.n639 B.n211 163.367
R978 B.n643 B.n211 163.367
R979 B.n643 B.n204 163.367
R980 B.n651 B.n204 163.367
R981 B.n651 B.n202 163.367
R982 B.n655 B.n202 163.367
R983 B.n655 B.n197 163.367
R984 B.n663 B.n197 163.367
R985 B.n663 B.n195 163.367
R986 B.n667 B.n195 163.367
R987 B.n667 B.n189 163.367
R988 B.n675 B.n189 163.367
R989 B.n675 B.n187 163.367
R990 B.n679 B.n187 163.367
R991 B.n679 B.n181 163.367
R992 B.n687 B.n181 163.367
R993 B.n687 B.n179 163.367
R994 B.n691 B.n179 163.367
R995 B.n691 B.n173 163.367
R996 B.n699 B.n173 163.367
R997 B.n699 B.n171 163.367
R998 B.n704 B.n171 163.367
R999 B.n704 B.n165 163.367
R1000 B.n712 B.n165 163.367
R1001 B.n713 B.n712 163.367
R1002 B.n713 B.n5 163.367
R1003 B.n6 B.n5 163.367
R1004 B.n7 B.n6 163.367
R1005 B.n719 B.n7 163.367
R1006 B.n720 B.n719 163.367
R1007 B.n720 B.n13 163.367
R1008 B.n14 B.n13 163.367
R1009 B.n15 B.n14 163.367
R1010 B.n725 B.n15 163.367
R1011 B.n725 B.n20 163.367
R1012 B.n21 B.n20 163.367
R1013 B.n22 B.n21 163.367
R1014 B.n730 B.n22 163.367
R1015 B.n730 B.n27 163.367
R1016 B.n28 B.n27 163.367
R1017 B.n29 B.n28 163.367
R1018 B.n735 B.n29 163.367
R1019 B.n735 B.n34 163.367
R1020 B.n35 B.n34 163.367
R1021 B.n36 B.n35 163.367
R1022 B.n740 B.n36 163.367
R1023 B.n740 B.n41 163.367
R1024 B.n42 B.n41 163.367
R1025 B.n43 B.n42 163.367
R1026 B.n745 B.n43 163.367
R1027 B.n745 B.n48 163.367
R1028 B.n49 B.n48 163.367
R1029 B.n50 B.n49 163.367
R1030 B.n750 B.n50 163.367
R1031 B.n750 B.n55 163.367
R1032 B.n56 B.n55 163.367
R1033 B.n57 B.n56 163.367
R1034 B.n755 B.n57 163.367
R1035 B.n755 B.n62 163.367
R1036 B.n63 B.n62 163.367
R1037 B.n64 B.n63 163.367
R1038 B.n760 B.n64 163.367
R1039 B.n760 B.n69 163.367
R1040 B.n70 B.n69 163.367
R1041 B.n71 B.n70 163.367
R1042 B.n765 B.n71 163.367
R1043 B.n765 B.n76 163.367
R1044 B.n77 B.n76 163.367
R1045 B.n78 B.n77 163.367
R1046 B.n770 B.n78 163.367
R1047 B.n770 B.n83 163.367
R1048 B.n84 B.n83 163.367
R1049 B.n85 B.n84 163.367
R1050 B.n775 B.n85 163.367
R1051 B.n775 B.n90 163.367
R1052 B.n91 B.n90 163.367
R1053 B.n92 B.n91 163.367
R1054 B.n780 B.n92 163.367
R1055 B.n780 B.n97 163.367
R1056 B.n98 B.n97 163.367
R1057 B.n99 B.n98 163.367
R1058 B.n785 B.n99 163.367
R1059 B.n785 B.n104 163.367
R1060 B.n105 B.n104 163.367
R1061 B.n106 B.n105 163.367
R1062 B.n537 B.n535 163.367
R1063 B.n535 B.n534 163.367
R1064 B.n531 B.n530 163.367
R1065 B.n528 B.n283 163.367
R1066 B.n524 B.n522 163.367
R1067 B.n520 B.n285 163.367
R1068 B.n516 B.n514 163.367
R1069 B.n512 B.n287 163.367
R1070 B.n508 B.n506 163.367
R1071 B.n504 B.n289 163.367
R1072 B.n500 B.n498 163.367
R1073 B.n496 B.n291 163.367
R1074 B.n492 B.n490 163.367
R1075 B.n488 B.n293 163.367
R1076 B.n484 B.n482 163.367
R1077 B.n480 B.n295 163.367
R1078 B.n476 B.n474 163.367
R1079 B.n472 B.n297 163.367
R1080 B.n468 B.n466 163.367
R1081 B.n464 B.n299 163.367
R1082 B.n460 B.n458 163.367
R1083 B.n456 B.n301 163.367
R1084 B.n452 B.n450 163.367
R1085 B.n448 B.n303 163.367
R1086 B.n443 B.n441 163.367
R1087 B.n439 B.n307 163.367
R1088 B.n435 B.n433 163.367
R1089 B.n431 B.n309 163.367
R1090 B.n426 B.n424 163.367
R1091 B.n422 B.n313 163.367
R1092 B.n418 B.n416 163.367
R1093 B.n414 B.n315 163.367
R1094 B.n410 B.n408 163.367
R1095 B.n406 B.n317 163.367
R1096 B.n402 B.n400 163.367
R1097 B.n398 B.n319 163.367
R1098 B.n394 B.n392 163.367
R1099 B.n390 B.n321 163.367
R1100 B.n386 B.n384 163.367
R1101 B.n382 B.n323 163.367
R1102 B.n378 B.n376 163.367
R1103 B.n374 B.n325 163.367
R1104 B.n370 B.n368 163.367
R1105 B.n366 B.n327 163.367
R1106 B.n362 B.n360 163.367
R1107 B.n358 B.n329 163.367
R1108 B.n354 B.n352 163.367
R1109 B.n350 B.n331 163.367
R1110 B.n346 B.n344 163.367
R1111 B.n342 B.n333 163.367
R1112 B.n338 B.n336 163.367
R1113 B.n541 B.n273 163.367
R1114 B.n549 B.n273 163.367
R1115 B.n549 B.n271 163.367
R1116 B.n553 B.n271 163.367
R1117 B.n553 B.n265 163.367
R1118 B.n561 B.n265 163.367
R1119 B.n561 B.n263 163.367
R1120 B.n565 B.n263 163.367
R1121 B.n565 B.n257 163.367
R1122 B.n573 B.n257 163.367
R1123 B.n573 B.n255 163.367
R1124 B.n577 B.n255 163.367
R1125 B.n577 B.n249 163.367
R1126 B.n585 B.n249 163.367
R1127 B.n585 B.n247 163.367
R1128 B.n589 B.n247 163.367
R1129 B.n589 B.n241 163.367
R1130 B.n597 B.n241 163.367
R1131 B.n597 B.n239 163.367
R1132 B.n601 B.n239 163.367
R1133 B.n601 B.n233 163.367
R1134 B.n609 B.n233 163.367
R1135 B.n609 B.n231 163.367
R1136 B.n613 B.n231 163.367
R1137 B.n613 B.n225 163.367
R1138 B.n621 B.n225 163.367
R1139 B.n621 B.n223 163.367
R1140 B.n625 B.n223 163.367
R1141 B.n625 B.n217 163.367
R1142 B.n633 B.n217 163.367
R1143 B.n633 B.n215 163.367
R1144 B.n637 B.n215 163.367
R1145 B.n637 B.n209 163.367
R1146 B.n645 B.n209 163.367
R1147 B.n645 B.n207 163.367
R1148 B.n649 B.n207 163.367
R1149 B.n649 B.n201 163.367
R1150 B.n657 B.n201 163.367
R1151 B.n657 B.n199 163.367
R1152 B.n661 B.n199 163.367
R1153 B.n661 B.n193 163.367
R1154 B.n669 B.n193 163.367
R1155 B.n669 B.n191 163.367
R1156 B.n673 B.n191 163.367
R1157 B.n673 B.n185 163.367
R1158 B.n681 B.n185 163.367
R1159 B.n681 B.n183 163.367
R1160 B.n685 B.n183 163.367
R1161 B.n685 B.n177 163.367
R1162 B.n693 B.n177 163.367
R1163 B.n693 B.n175 163.367
R1164 B.n697 B.n175 163.367
R1165 B.n697 B.n169 163.367
R1166 B.n706 B.n169 163.367
R1167 B.n706 B.n167 163.367
R1168 B.n710 B.n167 163.367
R1169 B.n710 B.n3 163.367
R1170 B.n1115 B.n3 163.367
R1171 B.n1111 B.n2 163.367
R1172 B.n1111 B.n1110 163.367
R1173 B.n1110 B.n9 163.367
R1174 B.n1106 B.n9 163.367
R1175 B.n1106 B.n11 163.367
R1176 B.n1102 B.n11 163.367
R1177 B.n1102 B.n17 163.367
R1178 B.n1098 B.n17 163.367
R1179 B.n1098 B.n19 163.367
R1180 B.n1094 B.n19 163.367
R1181 B.n1094 B.n24 163.367
R1182 B.n1090 B.n24 163.367
R1183 B.n1090 B.n26 163.367
R1184 B.n1086 B.n26 163.367
R1185 B.n1086 B.n31 163.367
R1186 B.n1082 B.n31 163.367
R1187 B.n1082 B.n33 163.367
R1188 B.n1078 B.n33 163.367
R1189 B.n1078 B.n38 163.367
R1190 B.n1074 B.n38 163.367
R1191 B.n1074 B.n40 163.367
R1192 B.n1070 B.n40 163.367
R1193 B.n1070 B.n45 163.367
R1194 B.n1066 B.n45 163.367
R1195 B.n1066 B.n47 163.367
R1196 B.n1062 B.n47 163.367
R1197 B.n1062 B.n52 163.367
R1198 B.n1058 B.n52 163.367
R1199 B.n1058 B.n54 163.367
R1200 B.n1054 B.n54 163.367
R1201 B.n1054 B.n59 163.367
R1202 B.n1050 B.n59 163.367
R1203 B.n1050 B.n61 163.367
R1204 B.n1046 B.n61 163.367
R1205 B.n1046 B.n66 163.367
R1206 B.n1042 B.n66 163.367
R1207 B.n1042 B.n68 163.367
R1208 B.n1038 B.n68 163.367
R1209 B.n1038 B.n73 163.367
R1210 B.n1034 B.n73 163.367
R1211 B.n1034 B.n75 163.367
R1212 B.n1030 B.n75 163.367
R1213 B.n1030 B.n80 163.367
R1214 B.n1026 B.n80 163.367
R1215 B.n1026 B.n82 163.367
R1216 B.n1022 B.n82 163.367
R1217 B.n1022 B.n87 163.367
R1218 B.n1018 B.n87 163.367
R1219 B.n1018 B.n89 163.367
R1220 B.n1014 B.n89 163.367
R1221 B.n1014 B.n94 163.367
R1222 B.n1010 B.n94 163.367
R1223 B.n1010 B.n96 163.367
R1224 B.n1006 B.n96 163.367
R1225 B.n1006 B.n101 163.367
R1226 B.n1002 B.n101 163.367
R1227 B.n1002 B.n103 163.367
R1228 B.n998 B.n103 163.367
R1229 B.n140 B.t18 153.5
R1230 B.n310 B.t16 153.5
R1231 B.n133 B.t8 153.482
R1232 B.n304 B.t13 153.482
R1233 B.n134 B.n133 83.3944
R1234 B.n141 B.n140 83.3944
R1235 B.n311 B.n310 83.3944
R1236 B.n305 B.n304 83.3944
R1237 B.n542 B.n278 79.2954
R1238 B.n999 B.n107 79.2954
R1239 B.n993 B.n108 71.676
R1240 B.n992 B.n991 71.676
R1241 B.n985 B.n110 71.676
R1242 B.n984 B.n983 71.676
R1243 B.n977 B.n112 71.676
R1244 B.n976 B.n975 71.676
R1245 B.n969 B.n114 71.676
R1246 B.n968 B.n967 71.676
R1247 B.n961 B.n116 71.676
R1248 B.n960 B.n959 71.676
R1249 B.n953 B.n118 71.676
R1250 B.n952 B.n951 71.676
R1251 B.n945 B.n120 71.676
R1252 B.n944 B.n943 71.676
R1253 B.n937 B.n122 71.676
R1254 B.n936 B.n935 71.676
R1255 B.n929 B.n124 71.676
R1256 B.n928 B.n927 71.676
R1257 B.n921 B.n126 71.676
R1258 B.n920 B.n919 71.676
R1259 B.n913 B.n128 71.676
R1260 B.n912 B.n911 71.676
R1261 B.n905 B.n130 71.676
R1262 B.n904 B.n903 71.676
R1263 B.n897 B.n132 71.676
R1264 B.n896 B.n895 71.676
R1265 B.n889 B.n137 71.676
R1266 B.n888 B.n887 71.676
R1267 B.n880 B.n139 71.676
R1268 B.n879 B.n878 71.676
R1269 B.n872 B.n143 71.676
R1270 B.n871 B.n870 71.676
R1271 B.n864 B.n145 71.676
R1272 B.n863 B.n862 71.676
R1273 B.n856 B.n147 71.676
R1274 B.n855 B.n854 71.676
R1275 B.n848 B.n149 71.676
R1276 B.n847 B.n846 71.676
R1277 B.n840 B.n151 71.676
R1278 B.n839 B.n838 71.676
R1279 B.n832 B.n153 71.676
R1280 B.n831 B.n830 71.676
R1281 B.n824 B.n155 71.676
R1282 B.n823 B.n822 71.676
R1283 B.n816 B.n157 71.676
R1284 B.n815 B.n814 71.676
R1285 B.n808 B.n159 71.676
R1286 B.n807 B.n806 71.676
R1287 B.n800 B.n161 71.676
R1288 B.n799 B.n798 71.676
R1289 B.n792 B.n163 71.676
R1290 B.n793 B.n792 71.676
R1291 B.n798 B.n797 71.676
R1292 B.n801 B.n800 71.676
R1293 B.n806 B.n805 71.676
R1294 B.n809 B.n808 71.676
R1295 B.n814 B.n813 71.676
R1296 B.n817 B.n816 71.676
R1297 B.n822 B.n821 71.676
R1298 B.n825 B.n824 71.676
R1299 B.n830 B.n829 71.676
R1300 B.n833 B.n832 71.676
R1301 B.n838 B.n837 71.676
R1302 B.n841 B.n840 71.676
R1303 B.n846 B.n845 71.676
R1304 B.n849 B.n848 71.676
R1305 B.n854 B.n853 71.676
R1306 B.n857 B.n856 71.676
R1307 B.n862 B.n861 71.676
R1308 B.n865 B.n864 71.676
R1309 B.n870 B.n869 71.676
R1310 B.n873 B.n872 71.676
R1311 B.n878 B.n877 71.676
R1312 B.n881 B.n880 71.676
R1313 B.n887 B.n886 71.676
R1314 B.n890 B.n889 71.676
R1315 B.n895 B.n894 71.676
R1316 B.n898 B.n897 71.676
R1317 B.n903 B.n902 71.676
R1318 B.n906 B.n905 71.676
R1319 B.n911 B.n910 71.676
R1320 B.n914 B.n913 71.676
R1321 B.n919 B.n918 71.676
R1322 B.n922 B.n921 71.676
R1323 B.n927 B.n926 71.676
R1324 B.n930 B.n929 71.676
R1325 B.n935 B.n934 71.676
R1326 B.n938 B.n937 71.676
R1327 B.n943 B.n942 71.676
R1328 B.n946 B.n945 71.676
R1329 B.n951 B.n950 71.676
R1330 B.n954 B.n953 71.676
R1331 B.n959 B.n958 71.676
R1332 B.n962 B.n961 71.676
R1333 B.n967 B.n966 71.676
R1334 B.n970 B.n969 71.676
R1335 B.n975 B.n974 71.676
R1336 B.n978 B.n977 71.676
R1337 B.n983 B.n982 71.676
R1338 B.n986 B.n985 71.676
R1339 B.n991 B.n990 71.676
R1340 B.n994 B.n993 71.676
R1341 B.n536 B.n279 71.676
R1342 B.n534 B.n281 71.676
R1343 B.n530 B.n529 71.676
R1344 B.n523 B.n283 71.676
R1345 B.n522 B.n521 71.676
R1346 B.n515 B.n285 71.676
R1347 B.n514 B.n513 71.676
R1348 B.n507 B.n287 71.676
R1349 B.n506 B.n505 71.676
R1350 B.n499 B.n289 71.676
R1351 B.n498 B.n497 71.676
R1352 B.n491 B.n291 71.676
R1353 B.n490 B.n489 71.676
R1354 B.n483 B.n293 71.676
R1355 B.n482 B.n481 71.676
R1356 B.n475 B.n295 71.676
R1357 B.n474 B.n473 71.676
R1358 B.n467 B.n297 71.676
R1359 B.n466 B.n465 71.676
R1360 B.n459 B.n299 71.676
R1361 B.n458 B.n457 71.676
R1362 B.n451 B.n301 71.676
R1363 B.n450 B.n449 71.676
R1364 B.n442 B.n303 71.676
R1365 B.n441 B.n440 71.676
R1366 B.n434 B.n307 71.676
R1367 B.n433 B.n432 71.676
R1368 B.n425 B.n309 71.676
R1369 B.n424 B.n423 71.676
R1370 B.n417 B.n313 71.676
R1371 B.n416 B.n415 71.676
R1372 B.n409 B.n315 71.676
R1373 B.n408 B.n407 71.676
R1374 B.n401 B.n317 71.676
R1375 B.n400 B.n399 71.676
R1376 B.n393 B.n319 71.676
R1377 B.n392 B.n391 71.676
R1378 B.n385 B.n321 71.676
R1379 B.n384 B.n383 71.676
R1380 B.n377 B.n323 71.676
R1381 B.n376 B.n375 71.676
R1382 B.n369 B.n325 71.676
R1383 B.n368 B.n367 71.676
R1384 B.n361 B.n327 71.676
R1385 B.n360 B.n359 71.676
R1386 B.n353 B.n329 71.676
R1387 B.n352 B.n351 71.676
R1388 B.n345 B.n331 71.676
R1389 B.n344 B.n343 71.676
R1390 B.n337 B.n333 71.676
R1391 B.n336 B.n335 71.676
R1392 B.n537 B.n536 71.676
R1393 B.n531 B.n281 71.676
R1394 B.n529 B.n528 71.676
R1395 B.n524 B.n523 71.676
R1396 B.n521 B.n520 71.676
R1397 B.n516 B.n515 71.676
R1398 B.n513 B.n512 71.676
R1399 B.n508 B.n507 71.676
R1400 B.n505 B.n504 71.676
R1401 B.n500 B.n499 71.676
R1402 B.n497 B.n496 71.676
R1403 B.n492 B.n491 71.676
R1404 B.n489 B.n488 71.676
R1405 B.n484 B.n483 71.676
R1406 B.n481 B.n480 71.676
R1407 B.n476 B.n475 71.676
R1408 B.n473 B.n472 71.676
R1409 B.n468 B.n467 71.676
R1410 B.n465 B.n464 71.676
R1411 B.n460 B.n459 71.676
R1412 B.n457 B.n456 71.676
R1413 B.n452 B.n451 71.676
R1414 B.n449 B.n448 71.676
R1415 B.n443 B.n442 71.676
R1416 B.n440 B.n439 71.676
R1417 B.n435 B.n434 71.676
R1418 B.n432 B.n431 71.676
R1419 B.n426 B.n425 71.676
R1420 B.n423 B.n422 71.676
R1421 B.n418 B.n417 71.676
R1422 B.n415 B.n414 71.676
R1423 B.n410 B.n409 71.676
R1424 B.n407 B.n406 71.676
R1425 B.n402 B.n401 71.676
R1426 B.n399 B.n398 71.676
R1427 B.n394 B.n393 71.676
R1428 B.n391 B.n390 71.676
R1429 B.n386 B.n385 71.676
R1430 B.n383 B.n382 71.676
R1431 B.n378 B.n377 71.676
R1432 B.n375 B.n374 71.676
R1433 B.n370 B.n369 71.676
R1434 B.n367 B.n366 71.676
R1435 B.n362 B.n361 71.676
R1436 B.n359 B.n358 71.676
R1437 B.n354 B.n353 71.676
R1438 B.n351 B.n350 71.676
R1439 B.n346 B.n345 71.676
R1440 B.n343 B.n342 71.676
R1441 B.n338 B.n337 71.676
R1442 B.n335 B.n277 71.676
R1443 B.n1116 B.n1115 71.676
R1444 B.n1116 B.n2 71.676
R1445 B.n141 B.t19 70.1057
R1446 B.n311 B.t15 70.1057
R1447 B.n134 B.t9 70.088
R1448 B.n305 B.t12 70.088
R1449 B.n135 B.n134 59.5399
R1450 B.n884 B.n141 59.5399
R1451 B.n428 B.n311 59.5399
R1452 B.n446 B.n305 59.5399
R1453 B.n542 B.n274 39.3586
R1454 B.n548 B.n274 39.3586
R1455 B.n548 B.n270 39.3586
R1456 B.n554 B.n270 39.3586
R1457 B.n554 B.n266 39.3586
R1458 B.n560 B.n266 39.3586
R1459 B.n560 B.n261 39.3586
R1460 B.n566 B.n261 39.3586
R1461 B.n566 B.n262 39.3586
R1462 B.n572 B.n254 39.3586
R1463 B.n578 B.n254 39.3586
R1464 B.n578 B.n250 39.3586
R1465 B.n584 B.n250 39.3586
R1466 B.n584 B.n246 39.3586
R1467 B.n590 B.n246 39.3586
R1468 B.n590 B.n242 39.3586
R1469 B.n596 B.n242 39.3586
R1470 B.n596 B.n238 39.3586
R1471 B.n602 B.n238 39.3586
R1472 B.n602 B.n234 39.3586
R1473 B.n608 B.n234 39.3586
R1474 B.n608 B.n229 39.3586
R1475 B.n614 B.n229 39.3586
R1476 B.n614 B.n230 39.3586
R1477 B.n620 B.n222 39.3586
R1478 B.n626 B.n222 39.3586
R1479 B.n626 B.n218 39.3586
R1480 B.n632 B.n218 39.3586
R1481 B.n632 B.n214 39.3586
R1482 B.n638 B.n214 39.3586
R1483 B.n638 B.n210 39.3586
R1484 B.n644 B.n210 39.3586
R1485 B.n644 B.n205 39.3586
R1486 B.n650 B.n205 39.3586
R1487 B.n650 B.n206 39.3586
R1488 B.n656 B.n198 39.3586
R1489 B.n662 B.n198 39.3586
R1490 B.n662 B.n194 39.3586
R1491 B.n668 B.n194 39.3586
R1492 B.n668 B.n190 39.3586
R1493 B.n674 B.n190 39.3586
R1494 B.n674 B.n186 39.3586
R1495 B.n680 B.n186 39.3586
R1496 B.n680 B.n182 39.3586
R1497 B.n686 B.n182 39.3586
R1498 B.n686 B.n178 39.3586
R1499 B.n692 B.n178 39.3586
R1500 B.n698 B.n174 39.3586
R1501 B.n698 B.n170 39.3586
R1502 B.n705 B.n170 39.3586
R1503 B.n705 B.n166 39.3586
R1504 B.n711 B.n166 39.3586
R1505 B.n711 B.n4 39.3586
R1506 B.n1114 B.n4 39.3586
R1507 B.n1114 B.n1113 39.3586
R1508 B.n1113 B.n1112 39.3586
R1509 B.n1112 B.n8 39.3586
R1510 B.n12 B.n8 39.3586
R1511 B.n1105 B.n12 39.3586
R1512 B.n1105 B.n1104 39.3586
R1513 B.n1104 B.n1103 39.3586
R1514 B.n1103 B.n16 39.3586
R1515 B.n1097 B.n1096 39.3586
R1516 B.n1096 B.n1095 39.3586
R1517 B.n1095 B.n23 39.3586
R1518 B.n1089 B.n23 39.3586
R1519 B.n1089 B.n1088 39.3586
R1520 B.n1088 B.n1087 39.3586
R1521 B.n1087 B.n30 39.3586
R1522 B.n1081 B.n30 39.3586
R1523 B.n1081 B.n1080 39.3586
R1524 B.n1080 B.n1079 39.3586
R1525 B.n1079 B.n37 39.3586
R1526 B.n1073 B.n37 39.3586
R1527 B.n1072 B.n1071 39.3586
R1528 B.n1071 B.n44 39.3586
R1529 B.n1065 B.n44 39.3586
R1530 B.n1065 B.n1064 39.3586
R1531 B.n1064 B.n1063 39.3586
R1532 B.n1063 B.n51 39.3586
R1533 B.n1057 B.n51 39.3586
R1534 B.n1057 B.n1056 39.3586
R1535 B.n1056 B.n1055 39.3586
R1536 B.n1055 B.n58 39.3586
R1537 B.n1049 B.n58 39.3586
R1538 B.n1048 B.n1047 39.3586
R1539 B.n1047 B.n65 39.3586
R1540 B.n1041 B.n65 39.3586
R1541 B.n1041 B.n1040 39.3586
R1542 B.n1040 B.n1039 39.3586
R1543 B.n1039 B.n72 39.3586
R1544 B.n1033 B.n72 39.3586
R1545 B.n1033 B.n1032 39.3586
R1546 B.n1032 B.n1031 39.3586
R1547 B.n1031 B.n79 39.3586
R1548 B.n1025 B.n79 39.3586
R1549 B.n1025 B.n1024 39.3586
R1550 B.n1024 B.n1023 39.3586
R1551 B.n1023 B.n86 39.3586
R1552 B.n1017 B.n86 39.3586
R1553 B.n1016 B.n1015 39.3586
R1554 B.n1015 B.n93 39.3586
R1555 B.n1009 B.n93 39.3586
R1556 B.n1009 B.n1008 39.3586
R1557 B.n1008 B.n1007 39.3586
R1558 B.n1007 B.n100 39.3586
R1559 B.n1001 B.n100 39.3586
R1560 B.n1001 B.n1000 39.3586
R1561 B.n1000 B.n999 39.3586
R1562 B.n206 B.t5 36.4646
R1563 B.t2 B.n1072 36.4646
R1564 B.n540 B.n539 34.4981
R1565 B.n544 B.n276 34.4981
R1566 B.n790 B.n789 34.4981
R1567 B.n997 B.n996 34.4981
R1568 B.n620 B.t4 28.3615
R1569 B.n1049 B.t0 28.3615
R1570 B.n572 B.t11 22.5735
R1571 B.n692 B.t3 22.5735
R1572 B.n1097 B.t1 22.5735
R1573 B.n1017 B.t7 22.5735
R1574 B B.n1117 18.0485
R1575 B.n262 B.t11 16.7856
R1576 B.t3 B.n174 16.7856
R1577 B.t1 B.n16 16.7856
R1578 B.t7 B.n1016 16.7856
R1579 B.n230 B.t4 10.9976
R1580 B.t0 B.n1048 10.9976
R1581 B.n540 B.n272 10.6151
R1582 B.n550 B.n272 10.6151
R1583 B.n551 B.n550 10.6151
R1584 B.n552 B.n551 10.6151
R1585 B.n552 B.n264 10.6151
R1586 B.n562 B.n264 10.6151
R1587 B.n563 B.n562 10.6151
R1588 B.n564 B.n563 10.6151
R1589 B.n564 B.n256 10.6151
R1590 B.n574 B.n256 10.6151
R1591 B.n575 B.n574 10.6151
R1592 B.n576 B.n575 10.6151
R1593 B.n576 B.n248 10.6151
R1594 B.n586 B.n248 10.6151
R1595 B.n587 B.n586 10.6151
R1596 B.n588 B.n587 10.6151
R1597 B.n588 B.n240 10.6151
R1598 B.n598 B.n240 10.6151
R1599 B.n599 B.n598 10.6151
R1600 B.n600 B.n599 10.6151
R1601 B.n600 B.n232 10.6151
R1602 B.n610 B.n232 10.6151
R1603 B.n611 B.n610 10.6151
R1604 B.n612 B.n611 10.6151
R1605 B.n612 B.n224 10.6151
R1606 B.n622 B.n224 10.6151
R1607 B.n623 B.n622 10.6151
R1608 B.n624 B.n623 10.6151
R1609 B.n624 B.n216 10.6151
R1610 B.n634 B.n216 10.6151
R1611 B.n635 B.n634 10.6151
R1612 B.n636 B.n635 10.6151
R1613 B.n636 B.n208 10.6151
R1614 B.n646 B.n208 10.6151
R1615 B.n647 B.n646 10.6151
R1616 B.n648 B.n647 10.6151
R1617 B.n648 B.n200 10.6151
R1618 B.n658 B.n200 10.6151
R1619 B.n659 B.n658 10.6151
R1620 B.n660 B.n659 10.6151
R1621 B.n660 B.n192 10.6151
R1622 B.n670 B.n192 10.6151
R1623 B.n671 B.n670 10.6151
R1624 B.n672 B.n671 10.6151
R1625 B.n672 B.n184 10.6151
R1626 B.n682 B.n184 10.6151
R1627 B.n683 B.n682 10.6151
R1628 B.n684 B.n683 10.6151
R1629 B.n684 B.n176 10.6151
R1630 B.n694 B.n176 10.6151
R1631 B.n695 B.n694 10.6151
R1632 B.n696 B.n695 10.6151
R1633 B.n696 B.n168 10.6151
R1634 B.n707 B.n168 10.6151
R1635 B.n708 B.n707 10.6151
R1636 B.n709 B.n708 10.6151
R1637 B.n709 B.n0 10.6151
R1638 B.n539 B.n538 10.6151
R1639 B.n538 B.n280 10.6151
R1640 B.n533 B.n280 10.6151
R1641 B.n533 B.n532 10.6151
R1642 B.n532 B.n282 10.6151
R1643 B.n527 B.n282 10.6151
R1644 B.n527 B.n526 10.6151
R1645 B.n526 B.n525 10.6151
R1646 B.n525 B.n284 10.6151
R1647 B.n519 B.n284 10.6151
R1648 B.n519 B.n518 10.6151
R1649 B.n518 B.n517 10.6151
R1650 B.n517 B.n286 10.6151
R1651 B.n511 B.n286 10.6151
R1652 B.n511 B.n510 10.6151
R1653 B.n510 B.n509 10.6151
R1654 B.n509 B.n288 10.6151
R1655 B.n503 B.n288 10.6151
R1656 B.n503 B.n502 10.6151
R1657 B.n502 B.n501 10.6151
R1658 B.n501 B.n290 10.6151
R1659 B.n495 B.n290 10.6151
R1660 B.n495 B.n494 10.6151
R1661 B.n494 B.n493 10.6151
R1662 B.n493 B.n292 10.6151
R1663 B.n487 B.n292 10.6151
R1664 B.n487 B.n486 10.6151
R1665 B.n486 B.n485 10.6151
R1666 B.n485 B.n294 10.6151
R1667 B.n479 B.n294 10.6151
R1668 B.n479 B.n478 10.6151
R1669 B.n478 B.n477 10.6151
R1670 B.n477 B.n296 10.6151
R1671 B.n471 B.n296 10.6151
R1672 B.n471 B.n470 10.6151
R1673 B.n470 B.n469 10.6151
R1674 B.n469 B.n298 10.6151
R1675 B.n463 B.n298 10.6151
R1676 B.n463 B.n462 10.6151
R1677 B.n462 B.n461 10.6151
R1678 B.n461 B.n300 10.6151
R1679 B.n455 B.n300 10.6151
R1680 B.n455 B.n454 10.6151
R1681 B.n454 B.n453 10.6151
R1682 B.n453 B.n302 10.6151
R1683 B.n447 B.n302 10.6151
R1684 B.n445 B.n444 10.6151
R1685 B.n444 B.n306 10.6151
R1686 B.n438 B.n306 10.6151
R1687 B.n438 B.n437 10.6151
R1688 B.n437 B.n436 10.6151
R1689 B.n436 B.n308 10.6151
R1690 B.n430 B.n308 10.6151
R1691 B.n430 B.n429 10.6151
R1692 B.n427 B.n312 10.6151
R1693 B.n421 B.n312 10.6151
R1694 B.n421 B.n420 10.6151
R1695 B.n420 B.n419 10.6151
R1696 B.n419 B.n314 10.6151
R1697 B.n413 B.n314 10.6151
R1698 B.n413 B.n412 10.6151
R1699 B.n412 B.n411 10.6151
R1700 B.n411 B.n316 10.6151
R1701 B.n405 B.n316 10.6151
R1702 B.n405 B.n404 10.6151
R1703 B.n404 B.n403 10.6151
R1704 B.n403 B.n318 10.6151
R1705 B.n397 B.n318 10.6151
R1706 B.n397 B.n396 10.6151
R1707 B.n396 B.n395 10.6151
R1708 B.n395 B.n320 10.6151
R1709 B.n389 B.n320 10.6151
R1710 B.n389 B.n388 10.6151
R1711 B.n388 B.n387 10.6151
R1712 B.n387 B.n322 10.6151
R1713 B.n381 B.n322 10.6151
R1714 B.n381 B.n380 10.6151
R1715 B.n380 B.n379 10.6151
R1716 B.n379 B.n324 10.6151
R1717 B.n373 B.n324 10.6151
R1718 B.n373 B.n372 10.6151
R1719 B.n372 B.n371 10.6151
R1720 B.n371 B.n326 10.6151
R1721 B.n365 B.n326 10.6151
R1722 B.n365 B.n364 10.6151
R1723 B.n364 B.n363 10.6151
R1724 B.n363 B.n328 10.6151
R1725 B.n357 B.n328 10.6151
R1726 B.n357 B.n356 10.6151
R1727 B.n356 B.n355 10.6151
R1728 B.n355 B.n330 10.6151
R1729 B.n349 B.n330 10.6151
R1730 B.n349 B.n348 10.6151
R1731 B.n348 B.n347 10.6151
R1732 B.n347 B.n332 10.6151
R1733 B.n341 B.n332 10.6151
R1734 B.n341 B.n340 10.6151
R1735 B.n340 B.n339 10.6151
R1736 B.n339 B.n334 10.6151
R1737 B.n334 B.n276 10.6151
R1738 B.n545 B.n544 10.6151
R1739 B.n546 B.n545 10.6151
R1740 B.n546 B.n268 10.6151
R1741 B.n556 B.n268 10.6151
R1742 B.n557 B.n556 10.6151
R1743 B.n558 B.n557 10.6151
R1744 B.n558 B.n259 10.6151
R1745 B.n568 B.n259 10.6151
R1746 B.n569 B.n568 10.6151
R1747 B.n570 B.n569 10.6151
R1748 B.n570 B.n252 10.6151
R1749 B.n580 B.n252 10.6151
R1750 B.n581 B.n580 10.6151
R1751 B.n582 B.n581 10.6151
R1752 B.n582 B.n244 10.6151
R1753 B.n592 B.n244 10.6151
R1754 B.n593 B.n592 10.6151
R1755 B.n594 B.n593 10.6151
R1756 B.n594 B.n236 10.6151
R1757 B.n604 B.n236 10.6151
R1758 B.n605 B.n604 10.6151
R1759 B.n606 B.n605 10.6151
R1760 B.n606 B.n227 10.6151
R1761 B.n616 B.n227 10.6151
R1762 B.n617 B.n616 10.6151
R1763 B.n618 B.n617 10.6151
R1764 B.n618 B.n220 10.6151
R1765 B.n628 B.n220 10.6151
R1766 B.n629 B.n628 10.6151
R1767 B.n630 B.n629 10.6151
R1768 B.n630 B.n212 10.6151
R1769 B.n640 B.n212 10.6151
R1770 B.n641 B.n640 10.6151
R1771 B.n642 B.n641 10.6151
R1772 B.n642 B.n203 10.6151
R1773 B.n652 B.n203 10.6151
R1774 B.n653 B.n652 10.6151
R1775 B.n654 B.n653 10.6151
R1776 B.n654 B.n196 10.6151
R1777 B.n664 B.n196 10.6151
R1778 B.n665 B.n664 10.6151
R1779 B.n666 B.n665 10.6151
R1780 B.n666 B.n188 10.6151
R1781 B.n676 B.n188 10.6151
R1782 B.n677 B.n676 10.6151
R1783 B.n678 B.n677 10.6151
R1784 B.n678 B.n180 10.6151
R1785 B.n688 B.n180 10.6151
R1786 B.n689 B.n688 10.6151
R1787 B.n690 B.n689 10.6151
R1788 B.n690 B.n172 10.6151
R1789 B.n700 B.n172 10.6151
R1790 B.n701 B.n700 10.6151
R1791 B.n703 B.n701 10.6151
R1792 B.n703 B.n702 10.6151
R1793 B.n702 B.n164 10.6151
R1794 B.n714 B.n164 10.6151
R1795 B.n715 B.n714 10.6151
R1796 B.n716 B.n715 10.6151
R1797 B.n717 B.n716 10.6151
R1798 B.n718 B.n717 10.6151
R1799 B.n721 B.n718 10.6151
R1800 B.n722 B.n721 10.6151
R1801 B.n723 B.n722 10.6151
R1802 B.n724 B.n723 10.6151
R1803 B.n726 B.n724 10.6151
R1804 B.n727 B.n726 10.6151
R1805 B.n728 B.n727 10.6151
R1806 B.n729 B.n728 10.6151
R1807 B.n731 B.n729 10.6151
R1808 B.n732 B.n731 10.6151
R1809 B.n733 B.n732 10.6151
R1810 B.n734 B.n733 10.6151
R1811 B.n736 B.n734 10.6151
R1812 B.n737 B.n736 10.6151
R1813 B.n738 B.n737 10.6151
R1814 B.n739 B.n738 10.6151
R1815 B.n741 B.n739 10.6151
R1816 B.n742 B.n741 10.6151
R1817 B.n743 B.n742 10.6151
R1818 B.n744 B.n743 10.6151
R1819 B.n746 B.n744 10.6151
R1820 B.n747 B.n746 10.6151
R1821 B.n748 B.n747 10.6151
R1822 B.n749 B.n748 10.6151
R1823 B.n751 B.n749 10.6151
R1824 B.n752 B.n751 10.6151
R1825 B.n753 B.n752 10.6151
R1826 B.n754 B.n753 10.6151
R1827 B.n756 B.n754 10.6151
R1828 B.n757 B.n756 10.6151
R1829 B.n758 B.n757 10.6151
R1830 B.n759 B.n758 10.6151
R1831 B.n761 B.n759 10.6151
R1832 B.n762 B.n761 10.6151
R1833 B.n763 B.n762 10.6151
R1834 B.n764 B.n763 10.6151
R1835 B.n766 B.n764 10.6151
R1836 B.n767 B.n766 10.6151
R1837 B.n768 B.n767 10.6151
R1838 B.n769 B.n768 10.6151
R1839 B.n771 B.n769 10.6151
R1840 B.n772 B.n771 10.6151
R1841 B.n773 B.n772 10.6151
R1842 B.n774 B.n773 10.6151
R1843 B.n776 B.n774 10.6151
R1844 B.n777 B.n776 10.6151
R1845 B.n778 B.n777 10.6151
R1846 B.n779 B.n778 10.6151
R1847 B.n781 B.n779 10.6151
R1848 B.n782 B.n781 10.6151
R1849 B.n783 B.n782 10.6151
R1850 B.n784 B.n783 10.6151
R1851 B.n786 B.n784 10.6151
R1852 B.n787 B.n786 10.6151
R1853 B.n788 B.n787 10.6151
R1854 B.n789 B.n788 10.6151
R1855 B.n1109 B.n1 10.6151
R1856 B.n1109 B.n1108 10.6151
R1857 B.n1108 B.n1107 10.6151
R1858 B.n1107 B.n10 10.6151
R1859 B.n1101 B.n10 10.6151
R1860 B.n1101 B.n1100 10.6151
R1861 B.n1100 B.n1099 10.6151
R1862 B.n1099 B.n18 10.6151
R1863 B.n1093 B.n18 10.6151
R1864 B.n1093 B.n1092 10.6151
R1865 B.n1092 B.n1091 10.6151
R1866 B.n1091 B.n25 10.6151
R1867 B.n1085 B.n25 10.6151
R1868 B.n1085 B.n1084 10.6151
R1869 B.n1084 B.n1083 10.6151
R1870 B.n1083 B.n32 10.6151
R1871 B.n1077 B.n32 10.6151
R1872 B.n1077 B.n1076 10.6151
R1873 B.n1076 B.n1075 10.6151
R1874 B.n1075 B.n39 10.6151
R1875 B.n1069 B.n39 10.6151
R1876 B.n1069 B.n1068 10.6151
R1877 B.n1068 B.n1067 10.6151
R1878 B.n1067 B.n46 10.6151
R1879 B.n1061 B.n46 10.6151
R1880 B.n1061 B.n1060 10.6151
R1881 B.n1060 B.n1059 10.6151
R1882 B.n1059 B.n53 10.6151
R1883 B.n1053 B.n53 10.6151
R1884 B.n1053 B.n1052 10.6151
R1885 B.n1052 B.n1051 10.6151
R1886 B.n1051 B.n60 10.6151
R1887 B.n1045 B.n60 10.6151
R1888 B.n1045 B.n1044 10.6151
R1889 B.n1044 B.n1043 10.6151
R1890 B.n1043 B.n67 10.6151
R1891 B.n1037 B.n67 10.6151
R1892 B.n1037 B.n1036 10.6151
R1893 B.n1036 B.n1035 10.6151
R1894 B.n1035 B.n74 10.6151
R1895 B.n1029 B.n74 10.6151
R1896 B.n1029 B.n1028 10.6151
R1897 B.n1028 B.n1027 10.6151
R1898 B.n1027 B.n81 10.6151
R1899 B.n1021 B.n81 10.6151
R1900 B.n1021 B.n1020 10.6151
R1901 B.n1020 B.n1019 10.6151
R1902 B.n1019 B.n88 10.6151
R1903 B.n1013 B.n88 10.6151
R1904 B.n1013 B.n1012 10.6151
R1905 B.n1012 B.n1011 10.6151
R1906 B.n1011 B.n95 10.6151
R1907 B.n1005 B.n95 10.6151
R1908 B.n1005 B.n1004 10.6151
R1909 B.n1004 B.n1003 10.6151
R1910 B.n1003 B.n102 10.6151
R1911 B.n997 B.n102 10.6151
R1912 B.n996 B.n995 10.6151
R1913 B.n995 B.n109 10.6151
R1914 B.n989 B.n109 10.6151
R1915 B.n989 B.n988 10.6151
R1916 B.n988 B.n987 10.6151
R1917 B.n987 B.n111 10.6151
R1918 B.n981 B.n111 10.6151
R1919 B.n981 B.n980 10.6151
R1920 B.n980 B.n979 10.6151
R1921 B.n979 B.n113 10.6151
R1922 B.n973 B.n113 10.6151
R1923 B.n973 B.n972 10.6151
R1924 B.n972 B.n971 10.6151
R1925 B.n971 B.n115 10.6151
R1926 B.n965 B.n115 10.6151
R1927 B.n965 B.n964 10.6151
R1928 B.n964 B.n963 10.6151
R1929 B.n963 B.n117 10.6151
R1930 B.n957 B.n117 10.6151
R1931 B.n957 B.n956 10.6151
R1932 B.n956 B.n955 10.6151
R1933 B.n955 B.n119 10.6151
R1934 B.n949 B.n119 10.6151
R1935 B.n949 B.n948 10.6151
R1936 B.n948 B.n947 10.6151
R1937 B.n947 B.n121 10.6151
R1938 B.n941 B.n121 10.6151
R1939 B.n941 B.n940 10.6151
R1940 B.n940 B.n939 10.6151
R1941 B.n939 B.n123 10.6151
R1942 B.n933 B.n123 10.6151
R1943 B.n933 B.n932 10.6151
R1944 B.n932 B.n931 10.6151
R1945 B.n931 B.n125 10.6151
R1946 B.n925 B.n125 10.6151
R1947 B.n925 B.n924 10.6151
R1948 B.n924 B.n923 10.6151
R1949 B.n923 B.n127 10.6151
R1950 B.n917 B.n127 10.6151
R1951 B.n917 B.n916 10.6151
R1952 B.n916 B.n915 10.6151
R1953 B.n915 B.n129 10.6151
R1954 B.n909 B.n129 10.6151
R1955 B.n909 B.n908 10.6151
R1956 B.n908 B.n907 10.6151
R1957 B.n907 B.n131 10.6151
R1958 B.n901 B.n900 10.6151
R1959 B.n900 B.n899 10.6151
R1960 B.n899 B.n136 10.6151
R1961 B.n893 B.n136 10.6151
R1962 B.n893 B.n892 10.6151
R1963 B.n892 B.n891 10.6151
R1964 B.n891 B.n138 10.6151
R1965 B.n885 B.n138 10.6151
R1966 B.n883 B.n882 10.6151
R1967 B.n882 B.n142 10.6151
R1968 B.n876 B.n142 10.6151
R1969 B.n876 B.n875 10.6151
R1970 B.n875 B.n874 10.6151
R1971 B.n874 B.n144 10.6151
R1972 B.n868 B.n144 10.6151
R1973 B.n868 B.n867 10.6151
R1974 B.n867 B.n866 10.6151
R1975 B.n866 B.n146 10.6151
R1976 B.n860 B.n146 10.6151
R1977 B.n860 B.n859 10.6151
R1978 B.n859 B.n858 10.6151
R1979 B.n858 B.n148 10.6151
R1980 B.n852 B.n148 10.6151
R1981 B.n852 B.n851 10.6151
R1982 B.n851 B.n850 10.6151
R1983 B.n850 B.n150 10.6151
R1984 B.n844 B.n150 10.6151
R1985 B.n844 B.n843 10.6151
R1986 B.n843 B.n842 10.6151
R1987 B.n842 B.n152 10.6151
R1988 B.n836 B.n152 10.6151
R1989 B.n836 B.n835 10.6151
R1990 B.n835 B.n834 10.6151
R1991 B.n834 B.n154 10.6151
R1992 B.n828 B.n154 10.6151
R1993 B.n828 B.n827 10.6151
R1994 B.n827 B.n826 10.6151
R1995 B.n826 B.n156 10.6151
R1996 B.n820 B.n156 10.6151
R1997 B.n820 B.n819 10.6151
R1998 B.n819 B.n818 10.6151
R1999 B.n818 B.n158 10.6151
R2000 B.n812 B.n158 10.6151
R2001 B.n812 B.n811 10.6151
R2002 B.n811 B.n810 10.6151
R2003 B.n810 B.n160 10.6151
R2004 B.n804 B.n160 10.6151
R2005 B.n804 B.n803 10.6151
R2006 B.n803 B.n802 10.6151
R2007 B.n802 B.n162 10.6151
R2008 B.n796 B.n162 10.6151
R2009 B.n796 B.n795 10.6151
R2010 B.n795 B.n794 10.6151
R2011 B.n794 B.n790 10.6151
R2012 B.n1117 B.n0 8.11757
R2013 B.n1117 B.n1 8.11757
R2014 B.n446 B.n445 6.5566
R2015 B.n429 B.n428 6.5566
R2016 B.n901 B.n135 6.5566
R2017 B.n885 B.n884 6.5566
R2018 B.n447 B.n446 4.05904
R2019 B.n428 B.n427 4.05904
R2020 B.n135 B.n131 4.05904
R2021 B.n884 B.n883 4.05904
R2022 B.n656 B.t5 2.89448
R2023 B.n1073 B.t2 2.89448
R2024 VP.n18 VP.n17 161.3
R2025 VP.n19 VP.n14 161.3
R2026 VP.n21 VP.n20 161.3
R2027 VP.n22 VP.n13 161.3
R2028 VP.n24 VP.n23 161.3
R2029 VP.n25 VP.n12 161.3
R2030 VP.n27 VP.n26 161.3
R2031 VP.n28 VP.n11 161.3
R2032 VP.n30 VP.n29 161.3
R2033 VP.n61 VP.n60 161.3
R2034 VP.n59 VP.n1 161.3
R2035 VP.n58 VP.n57 161.3
R2036 VP.n56 VP.n2 161.3
R2037 VP.n55 VP.n54 161.3
R2038 VP.n53 VP.n3 161.3
R2039 VP.n52 VP.n51 161.3
R2040 VP.n50 VP.n4 161.3
R2041 VP.n49 VP.n48 161.3
R2042 VP.n46 VP.n5 161.3
R2043 VP.n45 VP.n44 161.3
R2044 VP.n43 VP.n6 161.3
R2045 VP.n42 VP.n41 161.3
R2046 VP.n40 VP.n7 161.3
R2047 VP.n39 VP.n38 161.3
R2048 VP.n37 VP.n8 161.3
R2049 VP.n36 VP.n35 161.3
R2050 VP.n34 VP.n9 161.3
R2051 VP.n15 VP.t1 116.038
R2052 VP.n33 VP.n32 87.6207
R2053 VP.n62 VP.n0 87.6207
R2054 VP.n31 VP.n10 87.6207
R2055 VP.n33 VP.t3 83.3489
R2056 VP.n47 VP.t4 83.3489
R2057 VP.n0 VP.t5 83.3489
R2058 VP.n10 VP.t2 83.3489
R2059 VP.n16 VP.t0 83.3489
R2060 VP.n16 VP.n15 62.9379
R2061 VP.n32 VP.n31 55.4463
R2062 VP.n41 VP.n40 50.2061
R2063 VP.n54 VP.n53 50.2061
R2064 VP.n23 VP.n22 50.2061
R2065 VP.n40 VP.n39 30.7807
R2066 VP.n54 VP.n2 30.7807
R2067 VP.n23 VP.n12 30.7807
R2068 VP.n35 VP.n34 24.4675
R2069 VP.n35 VP.n8 24.4675
R2070 VP.n39 VP.n8 24.4675
R2071 VP.n41 VP.n6 24.4675
R2072 VP.n45 VP.n6 24.4675
R2073 VP.n46 VP.n45 24.4675
R2074 VP.n48 VP.n4 24.4675
R2075 VP.n52 VP.n4 24.4675
R2076 VP.n53 VP.n52 24.4675
R2077 VP.n58 VP.n2 24.4675
R2078 VP.n59 VP.n58 24.4675
R2079 VP.n60 VP.n59 24.4675
R2080 VP.n27 VP.n12 24.4675
R2081 VP.n28 VP.n27 24.4675
R2082 VP.n29 VP.n28 24.4675
R2083 VP.n17 VP.n14 24.4675
R2084 VP.n21 VP.n14 24.4675
R2085 VP.n22 VP.n21 24.4675
R2086 VP.n47 VP.n46 12.234
R2087 VP.n48 VP.n47 12.234
R2088 VP.n17 VP.n16 12.234
R2089 VP.n18 VP.n15 2.47756
R2090 VP.n34 VP.n33 2.4472
R2091 VP.n60 VP.n0 2.4472
R2092 VP.n29 VP.n10 2.4472
R2093 VP.n31 VP.n30 0.354971
R2094 VP.n32 VP.n9 0.354971
R2095 VP.n62 VP.n61 0.354971
R2096 VP VP.n62 0.26696
R2097 VP.n19 VP.n18 0.189894
R2098 VP.n20 VP.n19 0.189894
R2099 VP.n20 VP.n13 0.189894
R2100 VP.n24 VP.n13 0.189894
R2101 VP.n25 VP.n24 0.189894
R2102 VP.n26 VP.n25 0.189894
R2103 VP.n26 VP.n11 0.189894
R2104 VP.n30 VP.n11 0.189894
R2105 VP.n36 VP.n9 0.189894
R2106 VP.n37 VP.n36 0.189894
R2107 VP.n38 VP.n37 0.189894
R2108 VP.n38 VP.n7 0.189894
R2109 VP.n42 VP.n7 0.189894
R2110 VP.n43 VP.n42 0.189894
R2111 VP.n44 VP.n43 0.189894
R2112 VP.n44 VP.n5 0.189894
R2113 VP.n49 VP.n5 0.189894
R2114 VP.n50 VP.n49 0.189894
R2115 VP.n51 VP.n50 0.189894
R2116 VP.n51 VP.n3 0.189894
R2117 VP.n55 VP.n3 0.189894
R2118 VP.n56 VP.n55 0.189894
R2119 VP.n57 VP.n56 0.189894
R2120 VP.n57 VP.n1 0.189894
R2121 VP.n61 VP.n1 0.189894
R2122 VDD1 VDD1.t4 68.6446
R2123 VDD1.n1 VDD1.t2 68.5308
R2124 VDD1.n1 VDD1.n0 65.2353
R2125 VDD1.n3 VDD1.n2 64.3639
R2126 VDD1.n3 VDD1.n1 50.0354
R2127 VDD1.n2 VDD1.t5 1.4426
R2128 VDD1.n2 VDD1.t3 1.4426
R2129 VDD1.n0 VDD1.t1 1.4426
R2130 VDD1.n0 VDD1.t0 1.4426
R2131 VDD1 VDD1.n3 0.869035
C0 VDD2 VTAIL 8.852691f
C1 VP VN 8.57703f
C2 VDD1 VP 8.5857f
C3 VDD1 VN 0.15259f
C4 VP VTAIL 8.587941f
C5 VN VTAIL 8.57295f
C6 VDD2 VP 0.573835f
C7 VDD2 VN 8.16695f
C8 VDD1 VTAIL 8.79187f
C9 VDD2 VDD1 1.94166f
C10 VDD2 B 7.337388f
C11 VDD1 B 7.724684f
C12 VTAIL B 9.383815f
C13 VN B 17.051f
C14 VP B 15.767994f
C15 VDD1.t4 B 2.7199f
C16 VDD1.t2 B 2.7189f
C17 VDD1.t1 B 0.234849f
C18 VDD1.t0 B 0.234849f
C19 VDD1.n0 B 2.12339f
C20 VDD1.n1 B 3.24915f
C21 VDD1.t5 B 0.234849f
C22 VDD1.t3 B 0.234849f
C23 VDD1.n2 B 2.11669f
C24 VDD1.n3 B 2.85703f
C25 VP.t5 B 2.62899f
C26 VP.n0 B 0.982956f
C27 VP.n1 B 0.017638f
C28 VP.n2 B 0.035336f
C29 VP.n3 B 0.017638f
C30 VP.n4 B 0.032874f
C31 VP.n5 B 0.017638f
C32 VP.t4 B 2.62899f
C33 VP.n6 B 0.032874f
C34 VP.n7 B 0.017638f
C35 VP.n8 B 0.032874f
C36 VP.n9 B 0.028468f
C37 VP.t3 B 2.62899f
C38 VP.t2 B 2.62899f
C39 VP.n10 B 0.982956f
C40 VP.n11 B 0.017638f
C41 VP.n12 B 0.035336f
C42 VP.n13 B 0.017638f
C43 VP.n14 B 0.032874f
C44 VP.t1 B 2.92707f
C45 VP.n15 B 0.931088f
C46 VP.t0 B 2.62899f
C47 VP.n16 B 0.978718f
C48 VP.n17 B 0.024759f
C49 VP.n18 B 0.230723f
C50 VP.n19 B 0.017638f
C51 VP.n20 B 0.017638f
C52 VP.n21 B 0.032874f
C53 VP.n22 B 0.032373f
C54 VP.n23 B 0.016663f
C55 VP.n24 B 0.017638f
C56 VP.n25 B 0.017638f
C57 VP.n26 B 0.017638f
C58 VP.n27 B 0.032874f
C59 VP.n28 B 0.032874f
C60 VP.n29 B 0.018267f
C61 VP.n30 B 0.028468f
C62 VP.n31 B 1.17492f
C63 VP.n32 B 1.18636f
C64 VP.n33 B 0.982956f
C65 VP.n34 B 0.018267f
C66 VP.n35 B 0.032874f
C67 VP.n36 B 0.017638f
C68 VP.n37 B 0.017638f
C69 VP.n38 B 0.017638f
C70 VP.n39 B 0.035336f
C71 VP.n40 B 0.016663f
C72 VP.n41 B 0.032373f
C73 VP.n42 B 0.017638f
C74 VP.n43 B 0.017638f
C75 VP.n44 B 0.017638f
C76 VP.n45 B 0.032874f
C77 VP.n46 B 0.024759f
C78 VP.n47 B 0.914364f
C79 VP.n48 B 0.024759f
C80 VP.n49 B 0.017638f
C81 VP.n50 B 0.017638f
C82 VP.n51 B 0.017638f
C83 VP.n52 B 0.032874f
C84 VP.n53 B 0.032373f
C85 VP.n54 B 0.016663f
C86 VP.n55 B 0.017638f
C87 VP.n56 B 0.017638f
C88 VP.n57 B 0.017638f
C89 VP.n58 B 0.032874f
C90 VP.n59 B 0.032874f
C91 VP.n60 B 0.018267f
C92 VP.n61 B 0.028468f
C93 VP.n62 B 0.056098f
C94 VTAIL.t7 B 0.26212f
C95 VTAIL.t9 B 0.26212f
C96 VTAIL.n0 B 2.29655f
C97 VTAIL.n1 B 0.483722f
C98 VTAIL.t3 B 2.93072f
C99 VTAIL.n2 B 0.77632f
C100 VTAIL.t4 B 0.26212f
C101 VTAIL.t5 B 0.26212f
C102 VTAIL.n3 B 2.29655f
C103 VTAIL.n4 B 2.34145f
C104 VTAIL.t10 B 0.26212f
C105 VTAIL.t11 B 0.26212f
C106 VTAIL.n5 B 2.29656f
C107 VTAIL.n6 B 2.34145f
C108 VTAIL.t6 B 2.93072f
C109 VTAIL.n7 B 0.776317f
C110 VTAIL.t1 B 0.26212f
C111 VTAIL.t2 B 0.26212f
C112 VTAIL.n8 B 2.29656f
C113 VTAIL.n9 B 0.695612f
C114 VTAIL.t0 B 2.93072f
C115 VTAIL.n10 B 2.13359f
C116 VTAIL.t8 B 2.93072f
C117 VTAIL.n11 B 2.05692f
C118 VDD2.t4 B 2.68436f
C119 VDD2.t0 B 0.231865f
C120 VDD2.t5 B 0.231865f
C121 VDD2.n0 B 2.09642f
C122 VDD2.n1 B 3.06901f
C123 VDD2.t3 B 2.66759f
C124 VDD2.n2 B 2.81562f
C125 VDD2.t2 B 0.231865f
C126 VDD2.t1 B 0.231865f
C127 VDD2.n3 B 2.09638f
C128 VN.t3 B 2.58574f
C129 VN.n0 B 0.966787f
C130 VN.n1 B 0.017348f
C131 VN.n2 B 0.034755f
C132 VN.n3 B 0.017348f
C133 VN.n4 B 0.032333f
C134 VN.t4 B 2.87893f
C135 VN.n5 B 0.915772f
C136 VN.t2 B 2.58574f
C137 VN.n6 B 0.962619f
C138 VN.n7 B 0.024351f
C139 VN.n8 B 0.226927f
C140 VN.n9 B 0.017348f
C141 VN.n10 B 0.017348f
C142 VN.n11 B 0.032333f
C143 VN.n12 B 0.03184f
C144 VN.n13 B 0.016389f
C145 VN.n14 B 0.017348f
C146 VN.n15 B 0.017348f
C147 VN.n16 B 0.017348f
C148 VN.n17 B 0.032333f
C149 VN.n18 B 0.032333f
C150 VN.n19 B 0.017966f
C151 VN.n20 B 0.028f
C152 VN.n21 B 0.055175f
C153 VN.t1 B 2.58574f
C154 VN.n22 B 0.966787f
C155 VN.n23 B 0.017348f
C156 VN.n24 B 0.034755f
C157 VN.n25 B 0.017348f
C158 VN.n26 B 0.032333f
C159 VN.t5 B 2.87893f
C160 VN.n27 B 0.915772f
C161 VN.t0 B 2.58574f
C162 VN.n28 B 0.962619f
C163 VN.n29 B 0.024351f
C164 VN.n30 B 0.226927f
C165 VN.n31 B 0.017348f
C166 VN.n32 B 0.017348f
C167 VN.n33 B 0.032333f
C168 VN.n34 B 0.03184f
C169 VN.n35 B 0.016389f
C170 VN.n36 B 0.017348f
C171 VN.n37 B 0.017348f
C172 VN.n38 B 0.017348f
C173 VN.n39 B 0.032333f
C174 VN.n40 B 0.032333f
C175 VN.n41 B 0.017966f
C176 VN.n42 B 0.028f
C177 VN.n43 B 1.16245f
.ends

