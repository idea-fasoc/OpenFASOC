* NGSPICE file created from diff_pair_sample_0951.ext - technology: sky130A

.subckt diff_pair_sample_0951 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t12 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=6.1776 pd=32.46 as=2.6136 ps=16.17 w=15.84 l=2.72
X1 VDD2.t9 VN.t0 VTAIL.t5 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=6.1776 pd=32.46 as=2.6136 ps=16.17 w=15.84 l=2.72
X2 VDD2.t8 VN.t1 VTAIL.t9 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=2.6136 pd=16.17 as=6.1776 ps=32.46 w=15.84 l=2.72
X3 VDD2.t7 VN.t2 VTAIL.t3 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=6.1776 pd=32.46 as=2.6136 ps=16.17 w=15.84 l=2.72
X4 B.t11 B.t9 B.t10 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=6.1776 pd=32.46 as=0 ps=0 w=15.84 l=2.72
X5 VTAIL.t14 VP.t1 VDD1.t8 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=2.6136 pd=16.17 as=2.6136 ps=16.17 w=15.84 l=2.72
X6 VTAIL.t2 VN.t3 VDD2.t6 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=2.6136 pd=16.17 as=2.6136 ps=16.17 w=15.84 l=2.72
X7 VTAIL.t1 VN.t4 VDD2.t5 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=2.6136 pd=16.17 as=2.6136 ps=16.17 w=15.84 l=2.72
X8 VTAIL.t17 VP.t2 VDD1.t7 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=2.6136 pd=16.17 as=2.6136 ps=16.17 w=15.84 l=2.72
X9 VTAIL.t6 VN.t5 VDD2.t4 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=2.6136 pd=16.17 as=2.6136 ps=16.17 w=15.84 l=2.72
X10 B.t8 B.t6 B.t7 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=6.1776 pd=32.46 as=0 ps=0 w=15.84 l=2.72
X11 VDD2.t3 VN.t6 VTAIL.t4 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=2.6136 pd=16.17 as=6.1776 ps=32.46 w=15.84 l=2.72
X12 VDD2.t2 VN.t7 VTAIL.t7 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=2.6136 pd=16.17 as=2.6136 ps=16.17 w=15.84 l=2.72
X13 B.t5 B.t3 B.t4 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=6.1776 pd=32.46 as=0 ps=0 w=15.84 l=2.72
X14 VDD1.t6 VP.t3 VTAIL.t13 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=2.6136 pd=16.17 as=6.1776 ps=32.46 w=15.84 l=2.72
X15 VDD1.t5 VP.t4 VTAIL.t18 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=6.1776 pd=32.46 as=2.6136 ps=16.17 w=15.84 l=2.72
X16 B.t2 B.t0 B.t1 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=6.1776 pd=32.46 as=0 ps=0 w=15.84 l=2.72
X17 VDD1.t4 VP.t5 VTAIL.t11 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=2.6136 pd=16.17 as=2.6136 ps=16.17 w=15.84 l=2.72
X18 VTAIL.t16 VP.t6 VDD1.t3 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=2.6136 pd=16.17 as=2.6136 ps=16.17 w=15.84 l=2.72
X19 VDD1.t2 VP.t7 VTAIL.t19 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=2.6136 pd=16.17 as=2.6136 ps=16.17 w=15.84 l=2.72
X20 VDD2.t1 VN.t8 VTAIL.t8 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=2.6136 pd=16.17 as=2.6136 ps=16.17 w=15.84 l=2.72
X21 VTAIL.t10 VP.t8 VDD1.t1 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=2.6136 pd=16.17 as=2.6136 ps=16.17 w=15.84 l=2.72
X22 VDD1.t0 VP.t9 VTAIL.t15 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=2.6136 pd=16.17 as=6.1776 ps=32.46 w=15.84 l=2.72
X23 VTAIL.t0 VN.t9 VDD2.t0 w_n4630_n4136# sky130_fd_pr__pfet_01v8 ad=2.6136 pd=16.17 as=2.6136 ps=16.17 w=15.84 l=2.72
R0 VP.n24 VP.t4 172.297
R1 VP.n27 VP.n26 161.3
R2 VP.n28 VP.n23 161.3
R3 VP.n30 VP.n29 161.3
R4 VP.n31 VP.n22 161.3
R5 VP.n33 VP.n32 161.3
R6 VP.n34 VP.n21 161.3
R7 VP.n36 VP.n35 161.3
R8 VP.n37 VP.n20 161.3
R9 VP.n39 VP.n38 161.3
R10 VP.n40 VP.n19 161.3
R11 VP.n42 VP.n41 161.3
R12 VP.n43 VP.n18 161.3
R13 VP.n45 VP.n44 161.3
R14 VP.n47 VP.n46 161.3
R15 VP.n48 VP.n16 161.3
R16 VP.n50 VP.n49 161.3
R17 VP.n51 VP.n15 161.3
R18 VP.n53 VP.n52 161.3
R19 VP.n54 VP.n14 161.3
R20 VP.n96 VP.n0 161.3
R21 VP.n95 VP.n94 161.3
R22 VP.n93 VP.n1 161.3
R23 VP.n92 VP.n91 161.3
R24 VP.n90 VP.n2 161.3
R25 VP.n89 VP.n88 161.3
R26 VP.n87 VP.n86 161.3
R27 VP.n85 VP.n4 161.3
R28 VP.n84 VP.n83 161.3
R29 VP.n82 VP.n5 161.3
R30 VP.n81 VP.n80 161.3
R31 VP.n79 VP.n6 161.3
R32 VP.n78 VP.n77 161.3
R33 VP.n76 VP.n7 161.3
R34 VP.n75 VP.n74 161.3
R35 VP.n73 VP.n8 161.3
R36 VP.n72 VP.n71 161.3
R37 VP.n70 VP.n9 161.3
R38 VP.n69 VP.n68 161.3
R39 VP.n66 VP.n10 161.3
R40 VP.n65 VP.n64 161.3
R41 VP.n63 VP.n11 161.3
R42 VP.n62 VP.n61 161.3
R43 VP.n60 VP.n12 161.3
R44 VP.n59 VP.n58 161.3
R45 VP.n78 VP.t7 140.347
R46 VP.n13 VP.t0 140.347
R47 VP.n67 VP.t8 140.347
R48 VP.n3 VP.t6 140.347
R49 VP.n97 VP.t3 140.347
R50 VP.n36 VP.t5 140.347
R51 VP.n55 VP.t9 140.347
R52 VP.n17 VP.t1 140.347
R53 VP.n25 VP.t2 140.347
R54 VP.n57 VP.n13 105.99
R55 VP.n98 VP.n97 105.99
R56 VP.n56 VP.n55 105.99
R57 VP.n25 VP.n24 70.8607
R58 VP.n57 VP.n56 56.6474
R59 VP.n61 VP.n11 47.8428
R60 VP.n91 VP.n1 47.8428
R61 VP.n49 VP.n15 47.8428
R62 VP.n73 VP.n72 42.999
R63 VP.n84 VP.n5 42.999
R64 VP.n42 VP.n19 42.999
R65 VP.n31 VP.n30 42.999
R66 VP.n74 VP.n73 38.1551
R67 VP.n80 VP.n5 38.1551
R68 VP.n38 VP.n19 38.1551
R69 VP.n32 VP.n31 38.1551
R70 VP.n65 VP.n11 33.3113
R71 VP.n91 VP.n90 33.3113
R72 VP.n49 VP.n48 33.3113
R73 VP.n60 VP.n59 24.5923
R74 VP.n61 VP.n60 24.5923
R75 VP.n66 VP.n65 24.5923
R76 VP.n68 VP.n9 24.5923
R77 VP.n72 VP.n9 24.5923
R78 VP.n74 VP.n7 24.5923
R79 VP.n78 VP.n7 24.5923
R80 VP.n79 VP.n78 24.5923
R81 VP.n80 VP.n79 24.5923
R82 VP.n85 VP.n84 24.5923
R83 VP.n86 VP.n85 24.5923
R84 VP.n90 VP.n89 24.5923
R85 VP.n95 VP.n1 24.5923
R86 VP.n96 VP.n95 24.5923
R87 VP.n53 VP.n15 24.5923
R88 VP.n54 VP.n53 24.5923
R89 VP.n43 VP.n42 24.5923
R90 VP.n44 VP.n43 24.5923
R91 VP.n48 VP.n47 24.5923
R92 VP.n32 VP.n21 24.5923
R93 VP.n36 VP.n21 24.5923
R94 VP.n37 VP.n36 24.5923
R95 VP.n38 VP.n37 24.5923
R96 VP.n26 VP.n23 24.5923
R97 VP.n30 VP.n23 24.5923
R98 VP.n67 VP.n66 22.1332
R99 VP.n89 VP.n3 22.1332
R100 VP.n47 VP.n17 22.1332
R101 VP.n27 VP.n24 7.15857
R102 VP.n59 VP.n13 4.91887
R103 VP.n97 VP.n96 4.91887
R104 VP.n55 VP.n54 4.91887
R105 VP.n68 VP.n67 2.45968
R106 VP.n86 VP.n3 2.45968
R107 VP.n44 VP.n17 2.45968
R108 VP.n26 VP.n25 2.45968
R109 VP.n56 VP.n14 0.278335
R110 VP.n58 VP.n57 0.278335
R111 VP.n98 VP.n0 0.278335
R112 VP.n28 VP.n27 0.189894
R113 VP.n29 VP.n28 0.189894
R114 VP.n29 VP.n22 0.189894
R115 VP.n33 VP.n22 0.189894
R116 VP.n34 VP.n33 0.189894
R117 VP.n35 VP.n34 0.189894
R118 VP.n35 VP.n20 0.189894
R119 VP.n39 VP.n20 0.189894
R120 VP.n40 VP.n39 0.189894
R121 VP.n41 VP.n40 0.189894
R122 VP.n41 VP.n18 0.189894
R123 VP.n45 VP.n18 0.189894
R124 VP.n46 VP.n45 0.189894
R125 VP.n46 VP.n16 0.189894
R126 VP.n50 VP.n16 0.189894
R127 VP.n51 VP.n50 0.189894
R128 VP.n52 VP.n51 0.189894
R129 VP.n52 VP.n14 0.189894
R130 VP.n58 VP.n12 0.189894
R131 VP.n62 VP.n12 0.189894
R132 VP.n63 VP.n62 0.189894
R133 VP.n64 VP.n63 0.189894
R134 VP.n64 VP.n10 0.189894
R135 VP.n69 VP.n10 0.189894
R136 VP.n70 VP.n69 0.189894
R137 VP.n71 VP.n70 0.189894
R138 VP.n71 VP.n8 0.189894
R139 VP.n75 VP.n8 0.189894
R140 VP.n76 VP.n75 0.189894
R141 VP.n77 VP.n76 0.189894
R142 VP.n77 VP.n6 0.189894
R143 VP.n81 VP.n6 0.189894
R144 VP.n82 VP.n81 0.189894
R145 VP.n83 VP.n82 0.189894
R146 VP.n83 VP.n4 0.189894
R147 VP.n87 VP.n4 0.189894
R148 VP.n88 VP.n87 0.189894
R149 VP.n88 VP.n2 0.189894
R150 VP.n92 VP.n2 0.189894
R151 VP.n93 VP.n92 0.189894
R152 VP.n94 VP.n93 0.189894
R153 VP.n94 VP.n0 0.189894
R154 VP VP.n98 0.153485
R155 VTAIL.n11 VTAIL.t4 57.7243
R156 VTAIL.n16 VTAIL.t15 57.7242
R157 VTAIL.n17 VTAIL.t9 57.7241
R158 VTAIL.n2 VTAIL.t13 57.7241
R159 VTAIL.n15 VTAIL.n14 55.6723
R160 VTAIL.n13 VTAIL.n12 55.6723
R161 VTAIL.n10 VTAIL.n9 55.6723
R162 VTAIL.n8 VTAIL.n7 55.6723
R163 VTAIL.n19 VTAIL.n18 55.672
R164 VTAIL.n1 VTAIL.n0 55.672
R165 VTAIL.n4 VTAIL.n3 55.672
R166 VTAIL.n6 VTAIL.n5 55.672
R167 VTAIL.n8 VTAIL.n6 31.2807
R168 VTAIL.n17 VTAIL.n16 28.6514
R169 VTAIL.n10 VTAIL.n8 2.62981
R170 VTAIL.n11 VTAIL.n10 2.62981
R171 VTAIL.n15 VTAIL.n13 2.62981
R172 VTAIL.n16 VTAIL.n15 2.62981
R173 VTAIL.n6 VTAIL.n4 2.62981
R174 VTAIL.n4 VTAIL.n2 2.62981
R175 VTAIL.n19 VTAIL.n17 2.62981
R176 VTAIL.n18 VTAIL.t8 2.05258
R177 VTAIL.n18 VTAIL.t0 2.05258
R178 VTAIL.n0 VTAIL.t3 2.05258
R179 VTAIL.n0 VTAIL.t1 2.05258
R180 VTAIL.n3 VTAIL.t19 2.05258
R181 VTAIL.n3 VTAIL.t16 2.05258
R182 VTAIL.n5 VTAIL.t12 2.05258
R183 VTAIL.n5 VTAIL.t10 2.05258
R184 VTAIL.n14 VTAIL.t11 2.05258
R185 VTAIL.n14 VTAIL.t14 2.05258
R186 VTAIL.n12 VTAIL.t18 2.05258
R187 VTAIL.n12 VTAIL.t17 2.05258
R188 VTAIL.n9 VTAIL.t7 2.05258
R189 VTAIL.n9 VTAIL.t6 2.05258
R190 VTAIL.n7 VTAIL.t5 2.05258
R191 VTAIL.n7 VTAIL.t2 2.05258
R192 VTAIL VTAIL.n1 2.03067
R193 VTAIL.n13 VTAIL.n11 1.78498
R194 VTAIL.n2 VTAIL.n1 1.78498
R195 VTAIL VTAIL.n19 0.599638
R196 VDD1.n1 VDD1.t5 77.0324
R197 VDD1.n3 VDD1.t9 77.0323
R198 VDD1.n5 VDD1.n4 74.2674
R199 VDD1.n1 VDD1.n0 72.351
R200 VDD1.n7 VDD1.n6 72.3509
R201 VDD1.n3 VDD1.n2 72.3508
R202 VDD1.n7 VDD1.n5 51.7574
R203 VDD1.n6 VDD1.t8 2.05258
R204 VDD1.n6 VDD1.t0 2.05258
R205 VDD1.n0 VDD1.t7 2.05258
R206 VDD1.n0 VDD1.t4 2.05258
R207 VDD1.n4 VDD1.t3 2.05258
R208 VDD1.n4 VDD1.t6 2.05258
R209 VDD1.n2 VDD1.t1 2.05258
R210 VDD1.n2 VDD1.t2 2.05258
R211 VDD1 VDD1.n7 1.91429
R212 VDD1 VDD1.n1 0.716017
R213 VDD1.n5 VDD1.n3 0.602482
R214 VN.n10 VN.t2 172.297
R215 VN.n53 VN.t6 172.297
R216 VN.n83 VN.n43 161.3
R217 VN.n82 VN.n81 161.3
R218 VN.n80 VN.n44 161.3
R219 VN.n79 VN.n78 161.3
R220 VN.n77 VN.n45 161.3
R221 VN.n76 VN.n75 161.3
R222 VN.n74 VN.n73 161.3
R223 VN.n72 VN.n47 161.3
R224 VN.n71 VN.n70 161.3
R225 VN.n69 VN.n48 161.3
R226 VN.n68 VN.n67 161.3
R227 VN.n66 VN.n49 161.3
R228 VN.n65 VN.n64 161.3
R229 VN.n63 VN.n50 161.3
R230 VN.n62 VN.n61 161.3
R231 VN.n60 VN.n51 161.3
R232 VN.n59 VN.n58 161.3
R233 VN.n57 VN.n52 161.3
R234 VN.n56 VN.n55 161.3
R235 VN.n40 VN.n0 161.3
R236 VN.n39 VN.n38 161.3
R237 VN.n37 VN.n1 161.3
R238 VN.n36 VN.n35 161.3
R239 VN.n34 VN.n2 161.3
R240 VN.n33 VN.n32 161.3
R241 VN.n31 VN.n30 161.3
R242 VN.n29 VN.n4 161.3
R243 VN.n28 VN.n27 161.3
R244 VN.n26 VN.n5 161.3
R245 VN.n25 VN.n24 161.3
R246 VN.n23 VN.n6 161.3
R247 VN.n22 VN.n21 161.3
R248 VN.n20 VN.n7 161.3
R249 VN.n19 VN.n18 161.3
R250 VN.n17 VN.n8 161.3
R251 VN.n16 VN.n15 161.3
R252 VN.n14 VN.n9 161.3
R253 VN.n13 VN.n12 161.3
R254 VN.n22 VN.t8 140.347
R255 VN.n11 VN.t4 140.347
R256 VN.n3 VN.t9 140.347
R257 VN.n41 VN.t1 140.347
R258 VN.n65 VN.t7 140.347
R259 VN.n54 VN.t5 140.347
R260 VN.n46 VN.t3 140.347
R261 VN.n84 VN.t0 140.347
R262 VN.n42 VN.n41 105.99
R263 VN.n85 VN.n84 105.99
R264 VN.n11 VN.n10 70.8607
R265 VN.n54 VN.n53 70.8607
R266 VN VN.n85 56.9262
R267 VN.n35 VN.n1 47.8428
R268 VN.n78 VN.n44 47.8428
R269 VN.n17 VN.n16 42.999
R270 VN.n28 VN.n5 42.999
R271 VN.n60 VN.n59 42.999
R272 VN.n71 VN.n48 42.999
R273 VN.n18 VN.n17 38.1551
R274 VN.n24 VN.n5 38.1551
R275 VN.n61 VN.n60 38.1551
R276 VN.n67 VN.n48 38.1551
R277 VN.n35 VN.n34 33.3113
R278 VN.n78 VN.n77 33.3113
R279 VN.n12 VN.n9 24.5923
R280 VN.n16 VN.n9 24.5923
R281 VN.n18 VN.n7 24.5923
R282 VN.n22 VN.n7 24.5923
R283 VN.n23 VN.n22 24.5923
R284 VN.n24 VN.n23 24.5923
R285 VN.n29 VN.n28 24.5923
R286 VN.n30 VN.n29 24.5923
R287 VN.n34 VN.n33 24.5923
R288 VN.n39 VN.n1 24.5923
R289 VN.n40 VN.n39 24.5923
R290 VN.n59 VN.n52 24.5923
R291 VN.n55 VN.n52 24.5923
R292 VN.n67 VN.n66 24.5923
R293 VN.n66 VN.n65 24.5923
R294 VN.n65 VN.n50 24.5923
R295 VN.n61 VN.n50 24.5923
R296 VN.n77 VN.n76 24.5923
R297 VN.n73 VN.n72 24.5923
R298 VN.n72 VN.n71 24.5923
R299 VN.n83 VN.n82 24.5923
R300 VN.n82 VN.n44 24.5923
R301 VN.n33 VN.n3 22.1332
R302 VN.n76 VN.n46 22.1332
R303 VN.n56 VN.n53 7.15857
R304 VN.n13 VN.n10 7.15857
R305 VN.n41 VN.n40 4.91887
R306 VN.n84 VN.n83 4.91887
R307 VN.n12 VN.n11 2.45968
R308 VN.n30 VN.n3 2.45968
R309 VN.n55 VN.n54 2.45968
R310 VN.n73 VN.n46 2.45968
R311 VN.n85 VN.n43 0.278335
R312 VN.n42 VN.n0 0.278335
R313 VN.n81 VN.n43 0.189894
R314 VN.n81 VN.n80 0.189894
R315 VN.n80 VN.n79 0.189894
R316 VN.n79 VN.n45 0.189894
R317 VN.n75 VN.n45 0.189894
R318 VN.n75 VN.n74 0.189894
R319 VN.n74 VN.n47 0.189894
R320 VN.n70 VN.n47 0.189894
R321 VN.n70 VN.n69 0.189894
R322 VN.n69 VN.n68 0.189894
R323 VN.n68 VN.n49 0.189894
R324 VN.n64 VN.n49 0.189894
R325 VN.n64 VN.n63 0.189894
R326 VN.n63 VN.n62 0.189894
R327 VN.n62 VN.n51 0.189894
R328 VN.n58 VN.n51 0.189894
R329 VN.n58 VN.n57 0.189894
R330 VN.n57 VN.n56 0.189894
R331 VN.n14 VN.n13 0.189894
R332 VN.n15 VN.n14 0.189894
R333 VN.n15 VN.n8 0.189894
R334 VN.n19 VN.n8 0.189894
R335 VN.n20 VN.n19 0.189894
R336 VN.n21 VN.n20 0.189894
R337 VN.n21 VN.n6 0.189894
R338 VN.n25 VN.n6 0.189894
R339 VN.n26 VN.n25 0.189894
R340 VN.n27 VN.n26 0.189894
R341 VN.n27 VN.n4 0.189894
R342 VN.n31 VN.n4 0.189894
R343 VN.n32 VN.n31 0.189894
R344 VN.n32 VN.n2 0.189894
R345 VN.n36 VN.n2 0.189894
R346 VN.n37 VN.n36 0.189894
R347 VN.n38 VN.n37 0.189894
R348 VN.n38 VN.n0 0.189894
R349 VN VN.n42 0.153485
R350 VDD2.n1 VDD2.t7 77.0323
R351 VDD2.n4 VDD2.t9 74.4031
R352 VDD2.n3 VDD2.n2 74.2674
R353 VDD2 VDD2.n7 74.2646
R354 VDD2.n6 VDD2.n5 72.351
R355 VDD2.n1 VDD2.n0 72.3508
R356 VDD2.n4 VDD2.n3 49.8597
R357 VDD2.n6 VDD2.n4 2.62981
R358 VDD2.n7 VDD2.t4 2.05258
R359 VDD2.n7 VDD2.t3 2.05258
R360 VDD2.n5 VDD2.t6 2.05258
R361 VDD2.n5 VDD2.t2 2.05258
R362 VDD2.n2 VDD2.t0 2.05258
R363 VDD2.n2 VDD2.t8 2.05258
R364 VDD2.n0 VDD2.t5 2.05258
R365 VDD2.n0 VDD2.t1 2.05258
R366 VDD2 VDD2.n6 0.716017
R367 VDD2.n3 VDD2.n1 0.602482
R368 B.n704 B.n703 585
R369 B.n705 B.n94 585
R370 B.n707 B.n706 585
R371 B.n708 B.n93 585
R372 B.n710 B.n709 585
R373 B.n711 B.n92 585
R374 B.n713 B.n712 585
R375 B.n714 B.n91 585
R376 B.n716 B.n715 585
R377 B.n717 B.n90 585
R378 B.n719 B.n718 585
R379 B.n720 B.n89 585
R380 B.n722 B.n721 585
R381 B.n723 B.n88 585
R382 B.n725 B.n724 585
R383 B.n726 B.n87 585
R384 B.n728 B.n727 585
R385 B.n729 B.n86 585
R386 B.n731 B.n730 585
R387 B.n732 B.n85 585
R388 B.n734 B.n733 585
R389 B.n735 B.n84 585
R390 B.n737 B.n736 585
R391 B.n738 B.n83 585
R392 B.n740 B.n739 585
R393 B.n741 B.n82 585
R394 B.n743 B.n742 585
R395 B.n744 B.n81 585
R396 B.n746 B.n745 585
R397 B.n747 B.n80 585
R398 B.n749 B.n748 585
R399 B.n750 B.n79 585
R400 B.n752 B.n751 585
R401 B.n753 B.n78 585
R402 B.n755 B.n754 585
R403 B.n756 B.n77 585
R404 B.n758 B.n757 585
R405 B.n759 B.n76 585
R406 B.n761 B.n760 585
R407 B.n762 B.n75 585
R408 B.n764 B.n763 585
R409 B.n765 B.n74 585
R410 B.n767 B.n766 585
R411 B.n768 B.n73 585
R412 B.n770 B.n769 585
R413 B.n771 B.n72 585
R414 B.n773 B.n772 585
R415 B.n774 B.n71 585
R416 B.n776 B.n775 585
R417 B.n777 B.n70 585
R418 B.n779 B.n778 585
R419 B.n780 B.n69 585
R420 B.n782 B.n781 585
R421 B.n784 B.n783 585
R422 B.n785 B.n65 585
R423 B.n787 B.n786 585
R424 B.n788 B.n64 585
R425 B.n790 B.n789 585
R426 B.n791 B.n63 585
R427 B.n793 B.n792 585
R428 B.n794 B.n62 585
R429 B.n796 B.n795 585
R430 B.n798 B.n59 585
R431 B.n800 B.n799 585
R432 B.n801 B.n58 585
R433 B.n803 B.n802 585
R434 B.n804 B.n57 585
R435 B.n806 B.n805 585
R436 B.n807 B.n56 585
R437 B.n809 B.n808 585
R438 B.n810 B.n55 585
R439 B.n812 B.n811 585
R440 B.n813 B.n54 585
R441 B.n815 B.n814 585
R442 B.n816 B.n53 585
R443 B.n818 B.n817 585
R444 B.n819 B.n52 585
R445 B.n821 B.n820 585
R446 B.n822 B.n51 585
R447 B.n824 B.n823 585
R448 B.n825 B.n50 585
R449 B.n827 B.n826 585
R450 B.n828 B.n49 585
R451 B.n830 B.n829 585
R452 B.n831 B.n48 585
R453 B.n833 B.n832 585
R454 B.n834 B.n47 585
R455 B.n836 B.n835 585
R456 B.n837 B.n46 585
R457 B.n839 B.n838 585
R458 B.n840 B.n45 585
R459 B.n842 B.n841 585
R460 B.n843 B.n44 585
R461 B.n845 B.n844 585
R462 B.n846 B.n43 585
R463 B.n848 B.n847 585
R464 B.n849 B.n42 585
R465 B.n851 B.n850 585
R466 B.n852 B.n41 585
R467 B.n854 B.n853 585
R468 B.n855 B.n40 585
R469 B.n857 B.n856 585
R470 B.n858 B.n39 585
R471 B.n860 B.n859 585
R472 B.n861 B.n38 585
R473 B.n863 B.n862 585
R474 B.n864 B.n37 585
R475 B.n866 B.n865 585
R476 B.n867 B.n36 585
R477 B.n869 B.n868 585
R478 B.n870 B.n35 585
R479 B.n872 B.n871 585
R480 B.n873 B.n34 585
R481 B.n875 B.n874 585
R482 B.n876 B.n33 585
R483 B.n702 B.n95 585
R484 B.n701 B.n700 585
R485 B.n699 B.n96 585
R486 B.n698 B.n697 585
R487 B.n696 B.n97 585
R488 B.n695 B.n694 585
R489 B.n693 B.n98 585
R490 B.n692 B.n691 585
R491 B.n690 B.n99 585
R492 B.n689 B.n688 585
R493 B.n687 B.n100 585
R494 B.n686 B.n685 585
R495 B.n684 B.n101 585
R496 B.n683 B.n682 585
R497 B.n681 B.n102 585
R498 B.n680 B.n679 585
R499 B.n678 B.n103 585
R500 B.n677 B.n676 585
R501 B.n675 B.n104 585
R502 B.n674 B.n673 585
R503 B.n672 B.n105 585
R504 B.n671 B.n670 585
R505 B.n669 B.n106 585
R506 B.n668 B.n667 585
R507 B.n666 B.n107 585
R508 B.n665 B.n664 585
R509 B.n663 B.n108 585
R510 B.n662 B.n661 585
R511 B.n660 B.n109 585
R512 B.n659 B.n658 585
R513 B.n657 B.n110 585
R514 B.n656 B.n655 585
R515 B.n654 B.n111 585
R516 B.n653 B.n652 585
R517 B.n651 B.n112 585
R518 B.n650 B.n649 585
R519 B.n648 B.n113 585
R520 B.n647 B.n646 585
R521 B.n645 B.n114 585
R522 B.n644 B.n643 585
R523 B.n642 B.n115 585
R524 B.n641 B.n640 585
R525 B.n639 B.n116 585
R526 B.n638 B.n637 585
R527 B.n636 B.n117 585
R528 B.n635 B.n634 585
R529 B.n633 B.n118 585
R530 B.n632 B.n631 585
R531 B.n630 B.n119 585
R532 B.n629 B.n628 585
R533 B.n627 B.n120 585
R534 B.n626 B.n625 585
R535 B.n624 B.n121 585
R536 B.n623 B.n622 585
R537 B.n621 B.n122 585
R538 B.n620 B.n619 585
R539 B.n618 B.n123 585
R540 B.n617 B.n616 585
R541 B.n615 B.n124 585
R542 B.n614 B.n613 585
R543 B.n612 B.n125 585
R544 B.n611 B.n610 585
R545 B.n609 B.n126 585
R546 B.n608 B.n607 585
R547 B.n606 B.n127 585
R548 B.n605 B.n604 585
R549 B.n603 B.n128 585
R550 B.n602 B.n601 585
R551 B.n600 B.n129 585
R552 B.n599 B.n598 585
R553 B.n597 B.n130 585
R554 B.n596 B.n595 585
R555 B.n594 B.n131 585
R556 B.n593 B.n592 585
R557 B.n591 B.n132 585
R558 B.n590 B.n589 585
R559 B.n588 B.n133 585
R560 B.n587 B.n586 585
R561 B.n585 B.n134 585
R562 B.n584 B.n583 585
R563 B.n582 B.n135 585
R564 B.n581 B.n580 585
R565 B.n579 B.n136 585
R566 B.n578 B.n577 585
R567 B.n576 B.n137 585
R568 B.n575 B.n574 585
R569 B.n573 B.n138 585
R570 B.n572 B.n571 585
R571 B.n570 B.n139 585
R572 B.n569 B.n568 585
R573 B.n567 B.n140 585
R574 B.n566 B.n565 585
R575 B.n564 B.n141 585
R576 B.n563 B.n562 585
R577 B.n561 B.n142 585
R578 B.n560 B.n559 585
R579 B.n558 B.n143 585
R580 B.n557 B.n556 585
R581 B.n555 B.n144 585
R582 B.n554 B.n553 585
R583 B.n552 B.n145 585
R584 B.n551 B.n550 585
R585 B.n549 B.n146 585
R586 B.n548 B.n547 585
R587 B.n546 B.n147 585
R588 B.n545 B.n544 585
R589 B.n543 B.n148 585
R590 B.n542 B.n541 585
R591 B.n540 B.n149 585
R592 B.n539 B.n538 585
R593 B.n537 B.n150 585
R594 B.n536 B.n535 585
R595 B.n534 B.n151 585
R596 B.n533 B.n532 585
R597 B.n531 B.n152 585
R598 B.n530 B.n529 585
R599 B.n528 B.n153 585
R600 B.n527 B.n526 585
R601 B.n525 B.n154 585
R602 B.n524 B.n523 585
R603 B.n522 B.n155 585
R604 B.n521 B.n520 585
R605 B.n519 B.n156 585
R606 B.n518 B.n517 585
R607 B.n516 B.n157 585
R608 B.n342 B.n219 585
R609 B.n344 B.n343 585
R610 B.n345 B.n218 585
R611 B.n347 B.n346 585
R612 B.n348 B.n217 585
R613 B.n350 B.n349 585
R614 B.n351 B.n216 585
R615 B.n353 B.n352 585
R616 B.n354 B.n215 585
R617 B.n356 B.n355 585
R618 B.n357 B.n214 585
R619 B.n359 B.n358 585
R620 B.n360 B.n213 585
R621 B.n362 B.n361 585
R622 B.n363 B.n212 585
R623 B.n365 B.n364 585
R624 B.n366 B.n211 585
R625 B.n368 B.n367 585
R626 B.n369 B.n210 585
R627 B.n371 B.n370 585
R628 B.n372 B.n209 585
R629 B.n374 B.n373 585
R630 B.n375 B.n208 585
R631 B.n377 B.n376 585
R632 B.n378 B.n207 585
R633 B.n380 B.n379 585
R634 B.n381 B.n206 585
R635 B.n383 B.n382 585
R636 B.n384 B.n205 585
R637 B.n386 B.n385 585
R638 B.n387 B.n204 585
R639 B.n389 B.n388 585
R640 B.n390 B.n203 585
R641 B.n392 B.n391 585
R642 B.n393 B.n202 585
R643 B.n395 B.n394 585
R644 B.n396 B.n201 585
R645 B.n398 B.n397 585
R646 B.n399 B.n200 585
R647 B.n401 B.n400 585
R648 B.n402 B.n199 585
R649 B.n404 B.n403 585
R650 B.n405 B.n198 585
R651 B.n407 B.n406 585
R652 B.n408 B.n197 585
R653 B.n410 B.n409 585
R654 B.n411 B.n196 585
R655 B.n413 B.n412 585
R656 B.n414 B.n195 585
R657 B.n416 B.n415 585
R658 B.n417 B.n194 585
R659 B.n419 B.n418 585
R660 B.n420 B.n191 585
R661 B.n423 B.n422 585
R662 B.n424 B.n190 585
R663 B.n426 B.n425 585
R664 B.n427 B.n189 585
R665 B.n429 B.n428 585
R666 B.n430 B.n188 585
R667 B.n432 B.n431 585
R668 B.n433 B.n187 585
R669 B.n435 B.n434 585
R670 B.n437 B.n436 585
R671 B.n438 B.n183 585
R672 B.n440 B.n439 585
R673 B.n441 B.n182 585
R674 B.n443 B.n442 585
R675 B.n444 B.n181 585
R676 B.n446 B.n445 585
R677 B.n447 B.n180 585
R678 B.n449 B.n448 585
R679 B.n450 B.n179 585
R680 B.n452 B.n451 585
R681 B.n453 B.n178 585
R682 B.n455 B.n454 585
R683 B.n456 B.n177 585
R684 B.n458 B.n457 585
R685 B.n459 B.n176 585
R686 B.n461 B.n460 585
R687 B.n462 B.n175 585
R688 B.n464 B.n463 585
R689 B.n465 B.n174 585
R690 B.n467 B.n466 585
R691 B.n468 B.n173 585
R692 B.n470 B.n469 585
R693 B.n471 B.n172 585
R694 B.n473 B.n472 585
R695 B.n474 B.n171 585
R696 B.n476 B.n475 585
R697 B.n477 B.n170 585
R698 B.n479 B.n478 585
R699 B.n480 B.n169 585
R700 B.n482 B.n481 585
R701 B.n483 B.n168 585
R702 B.n485 B.n484 585
R703 B.n486 B.n167 585
R704 B.n488 B.n487 585
R705 B.n489 B.n166 585
R706 B.n491 B.n490 585
R707 B.n492 B.n165 585
R708 B.n494 B.n493 585
R709 B.n495 B.n164 585
R710 B.n497 B.n496 585
R711 B.n498 B.n163 585
R712 B.n500 B.n499 585
R713 B.n501 B.n162 585
R714 B.n503 B.n502 585
R715 B.n504 B.n161 585
R716 B.n506 B.n505 585
R717 B.n507 B.n160 585
R718 B.n509 B.n508 585
R719 B.n510 B.n159 585
R720 B.n512 B.n511 585
R721 B.n513 B.n158 585
R722 B.n515 B.n514 585
R723 B.n341 B.n340 585
R724 B.n339 B.n220 585
R725 B.n338 B.n337 585
R726 B.n336 B.n221 585
R727 B.n335 B.n334 585
R728 B.n333 B.n222 585
R729 B.n332 B.n331 585
R730 B.n330 B.n223 585
R731 B.n329 B.n328 585
R732 B.n327 B.n224 585
R733 B.n326 B.n325 585
R734 B.n324 B.n225 585
R735 B.n323 B.n322 585
R736 B.n321 B.n226 585
R737 B.n320 B.n319 585
R738 B.n318 B.n227 585
R739 B.n317 B.n316 585
R740 B.n315 B.n228 585
R741 B.n314 B.n313 585
R742 B.n312 B.n229 585
R743 B.n311 B.n310 585
R744 B.n309 B.n230 585
R745 B.n308 B.n307 585
R746 B.n306 B.n231 585
R747 B.n305 B.n304 585
R748 B.n303 B.n232 585
R749 B.n302 B.n301 585
R750 B.n300 B.n233 585
R751 B.n299 B.n298 585
R752 B.n297 B.n234 585
R753 B.n296 B.n295 585
R754 B.n294 B.n235 585
R755 B.n293 B.n292 585
R756 B.n291 B.n236 585
R757 B.n290 B.n289 585
R758 B.n288 B.n237 585
R759 B.n287 B.n286 585
R760 B.n285 B.n238 585
R761 B.n284 B.n283 585
R762 B.n282 B.n239 585
R763 B.n281 B.n280 585
R764 B.n279 B.n240 585
R765 B.n278 B.n277 585
R766 B.n276 B.n241 585
R767 B.n275 B.n274 585
R768 B.n273 B.n242 585
R769 B.n272 B.n271 585
R770 B.n270 B.n243 585
R771 B.n269 B.n268 585
R772 B.n267 B.n244 585
R773 B.n266 B.n265 585
R774 B.n264 B.n245 585
R775 B.n263 B.n262 585
R776 B.n261 B.n246 585
R777 B.n260 B.n259 585
R778 B.n258 B.n247 585
R779 B.n257 B.n256 585
R780 B.n255 B.n248 585
R781 B.n254 B.n253 585
R782 B.n252 B.n249 585
R783 B.n251 B.n250 585
R784 B.n2 B.n0 585
R785 B.n969 B.n1 585
R786 B.n968 B.n967 585
R787 B.n966 B.n3 585
R788 B.n965 B.n964 585
R789 B.n963 B.n4 585
R790 B.n962 B.n961 585
R791 B.n960 B.n5 585
R792 B.n959 B.n958 585
R793 B.n957 B.n6 585
R794 B.n956 B.n955 585
R795 B.n954 B.n7 585
R796 B.n953 B.n952 585
R797 B.n951 B.n8 585
R798 B.n950 B.n949 585
R799 B.n948 B.n9 585
R800 B.n947 B.n946 585
R801 B.n945 B.n10 585
R802 B.n944 B.n943 585
R803 B.n942 B.n11 585
R804 B.n941 B.n940 585
R805 B.n939 B.n12 585
R806 B.n938 B.n937 585
R807 B.n936 B.n13 585
R808 B.n935 B.n934 585
R809 B.n933 B.n14 585
R810 B.n932 B.n931 585
R811 B.n930 B.n15 585
R812 B.n929 B.n928 585
R813 B.n927 B.n16 585
R814 B.n926 B.n925 585
R815 B.n924 B.n17 585
R816 B.n923 B.n922 585
R817 B.n921 B.n18 585
R818 B.n920 B.n919 585
R819 B.n918 B.n19 585
R820 B.n917 B.n916 585
R821 B.n915 B.n20 585
R822 B.n914 B.n913 585
R823 B.n912 B.n21 585
R824 B.n911 B.n910 585
R825 B.n909 B.n22 585
R826 B.n908 B.n907 585
R827 B.n906 B.n23 585
R828 B.n905 B.n904 585
R829 B.n903 B.n24 585
R830 B.n902 B.n901 585
R831 B.n900 B.n25 585
R832 B.n899 B.n898 585
R833 B.n897 B.n26 585
R834 B.n896 B.n895 585
R835 B.n894 B.n27 585
R836 B.n893 B.n892 585
R837 B.n891 B.n28 585
R838 B.n890 B.n889 585
R839 B.n888 B.n29 585
R840 B.n887 B.n886 585
R841 B.n885 B.n30 585
R842 B.n884 B.n883 585
R843 B.n882 B.n31 585
R844 B.n881 B.n880 585
R845 B.n879 B.n32 585
R846 B.n878 B.n877 585
R847 B.n971 B.n970 585
R848 B.n340 B.n219 521.33
R849 B.n878 B.n33 521.33
R850 B.n514 B.n157 521.33
R851 B.n704 B.n95 521.33
R852 B.n184 B.t6 348.568
R853 B.n192 B.t0 348.568
R854 B.n60 B.t3 348.568
R855 B.n66 B.t9 348.568
R856 B.n184 B.t8 169.477
R857 B.n66 B.t10 169.477
R858 B.n192 B.t2 169.458
R859 B.n60 B.t4 169.458
R860 B.n340 B.n339 163.367
R861 B.n339 B.n338 163.367
R862 B.n338 B.n221 163.367
R863 B.n334 B.n221 163.367
R864 B.n334 B.n333 163.367
R865 B.n333 B.n332 163.367
R866 B.n332 B.n223 163.367
R867 B.n328 B.n223 163.367
R868 B.n328 B.n327 163.367
R869 B.n327 B.n326 163.367
R870 B.n326 B.n225 163.367
R871 B.n322 B.n225 163.367
R872 B.n322 B.n321 163.367
R873 B.n321 B.n320 163.367
R874 B.n320 B.n227 163.367
R875 B.n316 B.n227 163.367
R876 B.n316 B.n315 163.367
R877 B.n315 B.n314 163.367
R878 B.n314 B.n229 163.367
R879 B.n310 B.n229 163.367
R880 B.n310 B.n309 163.367
R881 B.n309 B.n308 163.367
R882 B.n308 B.n231 163.367
R883 B.n304 B.n231 163.367
R884 B.n304 B.n303 163.367
R885 B.n303 B.n302 163.367
R886 B.n302 B.n233 163.367
R887 B.n298 B.n233 163.367
R888 B.n298 B.n297 163.367
R889 B.n297 B.n296 163.367
R890 B.n296 B.n235 163.367
R891 B.n292 B.n235 163.367
R892 B.n292 B.n291 163.367
R893 B.n291 B.n290 163.367
R894 B.n290 B.n237 163.367
R895 B.n286 B.n237 163.367
R896 B.n286 B.n285 163.367
R897 B.n285 B.n284 163.367
R898 B.n284 B.n239 163.367
R899 B.n280 B.n239 163.367
R900 B.n280 B.n279 163.367
R901 B.n279 B.n278 163.367
R902 B.n278 B.n241 163.367
R903 B.n274 B.n241 163.367
R904 B.n274 B.n273 163.367
R905 B.n273 B.n272 163.367
R906 B.n272 B.n243 163.367
R907 B.n268 B.n243 163.367
R908 B.n268 B.n267 163.367
R909 B.n267 B.n266 163.367
R910 B.n266 B.n245 163.367
R911 B.n262 B.n245 163.367
R912 B.n262 B.n261 163.367
R913 B.n261 B.n260 163.367
R914 B.n260 B.n247 163.367
R915 B.n256 B.n247 163.367
R916 B.n256 B.n255 163.367
R917 B.n255 B.n254 163.367
R918 B.n254 B.n249 163.367
R919 B.n250 B.n249 163.367
R920 B.n250 B.n2 163.367
R921 B.n970 B.n2 163.367
R922 B.n970 B.n969 163.367
R923 B.n969 B.n968 163.367
R924 B.n968 B.n3 163.367
R925 B.n964 B.n3 163.367
R926 B.n964 B.n963 163.367
R927 B.n963 B.n962 163.367
R928 B.n962 B.n5 163.367
R929 B.n958 B.n5 163.367
R930 B.n958 B.n957 163.367
R931 B.n957 B.n956 163.367
R932 B.n956 B.n7 163.367
R933 B.n952 B.n7 163.367
R934 B.n952 B.n951 163.367
R935 B.n951 B.n950 163.367
R936 B.n950 B.n9 163.367
R937 B.n946 B.n9 163.367
R938 B.n946 B.n945 163.367
R939 B.n945 B.n944 163.367
R940 B.n944 B.n11 163.367
R941 B.n940 B.n11 163.367
R942 B.n940 B.n939 163.367
R943 B.n939 B.n938 163.367
R944 B.n938 B.n13 163.367
R945 B.n934 B.n13 163.367
R946 B.n934 B.n933 163.367
R947 B.n933 B.n932 163.367
R948 B.n932 B.n15 163.367
R949 B.n928 B.n15 163.367
R950 B.n928 B.n927 163.367
R951 B.n927 B.n926 163.367
R952 B.n926 B.n17 163.367
R953 B.n922 B.n17 163.367
R954 B.n922 B.n921 163.367
R955 B.n921 B.n920 163.367
R956 B.n920 B.n19 163.367
R957 B.n916 B.n19 163.367
R958 B.n916 B.n915 163.367
R959 B.n915 B.n914 163.367
R960 B.n914 B.n21 163.367
R961 B.n910 B.n21 163.367
R962 B.n910 B.n909 163.367
R963 B.n909 B.n908 163.367
R964 B.n908 B.n23 163.367
R965 B.n904 B.n23 163.367
R966 B.n904 B.n903 163.367
R967 B.n903 B.n902 163.367
R968 B.n902 B.n25 163.367
R969 B.n898 B.n25 163.367
R970 B.n898 B.n897 163.367
R971 B.n897 B.n896 163.367
R972 B.n896 B.n27 163.367
R973 B.n892 B.n27 163.367
R974 B.n892 B.n891 163.367
R975 B.n891 B.n890 163.367
R976 B.n890 B.n29 163.367
R977 B.n886 B.n29 163.367
R978 B.n886 B.n885 163.367
R979 B.n885 B.n884 163.367
R980 B.n884 B.n31 163.367
R981 B.n880 B.n31 163.367
R982 B.n880 B.n879 163.367
R983 B.n879 B.n878 163.367
R984 B.n344 B.n219 163.367
R985 B.n345 B.n344 163.367
R986 B.n346 B.n345 163.367
R987 B.n346 B.n217 163.367
R988 B.n350 B.n217 163.367
R989 B.n351 B.n350 163.367
R990 B.n352 B.n351 163.367
R991 B.n352 B.n215 163.367
R992 B.n356 B.n215 163.367
R993 B.n357 B.n356 163.367
R994 B.n358 B.n357 163.367
R995 B.n358 B.n213 163.367
R996 B.n362 B.n213 163.367
R997 B.n363 B.n362 163.367
R998 B.n364 B.n363 163.367
R999 B.n364 B.n211 163.367
R1000 B.n368 B.n211 163.367
R1001 B.n369 B.n368 163.367
R1002 B.n370 B.n369 163.367
R1003 B.n370 B.n209 163.367
R1004 B.n374 B.n209 163.367
R1005 B.n375 B.n374 163.367
R1006 B.n376 B.n375 163.367
R1007 B.n376 B.n207 163.367
R1008 B.n380 B.n207 163.367
R1009 B.n381 B.n380 163.367
R1010 B.n382 B.n381 163.367
R1011 B.n382 B.n205 163.367
R1012 B.n386 B.n205 163.367
R1013 B.n387 B.n386 163.367
R1014 B.n388 B.n387 163.367
R1015 B.n388 B.n203 163.367
R1016 B.n392 B.n203 163.367
R1017 B.n393 B.n392 163.367
R1018 B.n394 B.n393 163.367
R1019 B.n394 B.n201 163.367
R1020 B.n398 B.n201 163.367
R1021 B.n399 B.n398 163.367
R1022 B.n400 B.n399 163.367
R1023 B.n400 B.n199 163.367
R1024 B.n404 B.n199 163.367
R1025 B.n405 B.n404 163.367
R1026 B.n406 B.n405 163.367
R1027 B.n406 B.n197 163.367
R1028 B.n410 B.n197 163.367
R1029 B.n411 B.n410 163.367
R1030 B.n412 B.n411 163.367
R1031 B.n412 B.n195 163.367
R1032 B.n416 B.n195 163.367
R1033 B.n417 B.n416 163.367
R1034 B.n418 B.n417 163.367
R1035 B.n418 B.n191 163.367
R1036 B.n423 B.n191 163.367
R1037 B.n424 B.n423 163.367
R1038 B.n425 B.n424 163.367
R1039 B.n425 B.n189 163.367
R1040 B.n429 B.n189 163.367
R1041 B.n430 B.n429 163.367
R1042 B.n431 B.n430 163.367
R1043 B.n431 B.n187 163.367
R1044 B.n435 B.n187 163.367
R1045 B.n436 B.n435 163.367
R1046 B.n436 B.n183 163.367
R1047 B.n440 B.n183 163.367
R1048 B.n441 B.n440 163.367
R1049 B.n442 B.n441 163.367
R1050 B.n442 B.n181 163.367
R1051 B.n446 B.n181 163.367
R1052 B.n447 B.n446 163.367
R1053 B.n448 B.n447 163.367
R1054 B.n448 B.n179 163.367
R1055 B.n452 B.n179 163.367
R1056 B.n453 B.n452 163.367
R1057 B.n454 B.n453 163.367
R1058 B.n454 B.n177 163.367
R1059 B.n458 B.n177 163.367
R1060 B.n459 B.n458 163.367
R1061 B.n460 B.n459 163.367
R1062 B.n460 B.n175 163.367
R1063 B.n464 B.n175 163.367
R1064 B.n465 B.n464 163.367
R1065 B.n466 B.n465 163.367
R1066 B.n466 B.n173 163.367
R1067 B.n470 B.n173 163.367
R1068 B.n471 B.n470 163.367
R1069 B.n472 B.n471 163.367
R1070 B.n472 B.n171 163.367
R1071 B.n476 B.n171 163.367
R1072 B.n477 B.n476 163.367
R1073 B.n478 B.n477 163.367
R1074 B.n478 B.n169 163.367
R1075 B.n482 B.n169 163.367
R1076 B.n483 B.n482 163.367
R1077 B.n484 B.n483 163.367
R1078 B.n484 B.n167 163.367
R1079 B.n488 B.n167 163.367
R1080 B.n489 B.n488 163.367
R1081 B.n490 B.n489 163.367
R1082 B.n490 B.n165 163.367
R1083 B.n494 B.n165 163.367
R1084 B.n495 B.n494 163.367
R1085 B.n496 B.n495 163.367
R1086 B.n496 B.n163 163.367
R1087 B.n500 B.n163 163.367
R1088 B.n501 B.n500 163.367
R1089 B.n502 B.n501 163.367
R1090 B.n502 B.n161 163.367
R1091 B.n506 B.n161 163.367
R1092 B.n507 B.n506 163.367
R1093 B.n508 B.n507 163.367
R1094 B.n508 B.n159 163.367
R1095 B.n512 B.n159 163.367
R1096 B.n513 B.n512 163.367
R1097 B.n514 B.n513 163.367
R1098 B.n518 B.n157 163.367
R1099 B.n519 B.n518 163.367
R1100 B.n520 B.n519 163.367
R1101 B.n520 B.n155 163.367
R1102 B.n524 B.n155 163.367
R1103 B.n525 B.n524 163.367
R1104 B.n526 B.n525 163.367
R1105 B.n526 B.n153 163.367
R1106 B.n530 B.n153 163.367
R1107 B.n531 B.n530 163.367
R1108 B.n532 B.n531 163.367
R1109 B.n532 B.n151 163.367
R1110 B.n536 B.n151 163.367
R1111 B.n537 B.n536 163.367
R1112 B.n538 B.n537 163.367
R1113 B.n538 B.n149 163.367
R1114 B.n542 B.n149 163.367
R1115 B.n543 B.n542 163.367
R1116 B.n544 B.n543 163.367
R1117 B.n544 B.n147 163.367
R1118 B.n548 B.n147 163.367
R1119 B.n549 B.n548 163.367
R1120 B.n550 B.n549 163.367
R1121 B.n550 B.n145 163.367
R1122 B.n554 B.n145 163.367
R1123 B.n555 B.n554 163.367
R1124 B.n556 B.n555 163.367
R1125 B.n556 B.n143 163.367
R1126 B.n560 B.n143 163.367
R1127 B.n561 B.n560 163.367
R1128 B.n562 B.n561 163.367
R1129 B.n562 B.n141 163.367
R1130 B.n566 B.n141 163.367
R1131 B.n567 B.n566 163.367
R1132 B.n568 B.n567 163.367
R1133 B.n568 B.n139 163.367
R1134 B.n572 B.n139 163.367
R1135 B.n573 B.n572 163.367
R1136 B.n574 B.n573 163.367
R1137 B.n574 B.n137 163.367
R1138 B.n578 B.n137 163.367
R1139 B.n579 B.n578 163.367
R1140 B.n580 B.n579 163.367
R1141 B.n580 B.n135 163.367
R1142 B.n584 B.n135 163.367
R1143 B.n585 B.n584 163.367
R1144 B.n586 B.n585 163.367
R1145 B.n586 B.n133 163.367
R1146 B.n590 B.n133 163.367
R1147 B.n591 B.n590 163.367
R1148 B.n592 B.n591 163.367
R1149 B.n592 B.n131 163.367
R1150 B.n596 B.n131 163.367
R1151 B.n597 B.n596 163.367
R1152 B.n598 B.n597 163.367
R1153 B.n598 B.n129 163.367
R1154 B.n602 B.n129 163.367
R1155 B.n603 B.n602 163.367
R1156 B.n604 B.n603 163.367
R1157 B.n604 B.n127 163.367
R1158 B.n608 B.n127 163.367
R1159 B.n609 B.n608 163.367
R1160 B.n610 B.n609 163.367
R1161 B.n610 B.n125 163.367
R1162 B.n614 B.n125 163.367
R1163 B.n615 B.n614 163.367
R1164 B.n616 B.n615 163.367
R1165 B.n616 B.n123 163.367
R1166 B.n620 B.n123 163.367
R1167 B.n621 B.n620 163.367
R1168 B.n622 B.n621 163.367
R1169 B.n622 B.n121 163.367
R1170 B.n626 B.n121 163.367
R1171 B.n627 B.n626 163.367
R1172 B.n628 B.n627 163.367
R1173 B.n628 B.n119 163.367
R1174 B.n632 B.n119 163.367
R1175 B.n633 B.n632 163.367
R1176 B.n634 B.n633 163.367
R1177 B.n634 B.n117 163.367
R1178 B.n638 B.n117 163.367
R1179 B.n639 B.n638 163.367
R1180 B.n640 B.n639 163.367
R1181 B.n640 B.n115 163.367
R1182 B.n644 B.n115 163.367
R1183 B.n645 B.n644 163.367
R1184 B.n646 B.n645 163.367
R1185 B.n646 B.n113 163.367
R1186 B.n650 B.n113 163.367
R1187 B.n651 B.n650 163.367
R1188 B.n652 B.n651 163.367
R1189 B.n652 B.n111 163.367
R1190 B.n656 B.n111 163.367
R1191 B.n657 B.n656 163.367
R1192 B.n658 B.n657 163.367
R1193 B.n658 B.n109 163.367
R1194 B.n662 B.n109 163.367
R1195 B.n663 B.n662 163.367
R1196 B.n664 B.n663 163.367
R1197 B.n664 B.n107 163.367
R1198 B.n668 B.n107 163.367
R1199 B.n669 B.n668 163.367
R1200 B.n670 B.n669 163.367
R1201 B.n670 B.n105 163.367
R1202 B.n674 B.n105 163.367
R1203 B.n675 B.n674 163.367
R1204 B.n676 B.n675 163.367
R1205 B.n676 B.n103 163.367
R1206 B.n680 B.n103 163.367
R1207 B.n681 B.n680 163.367
R1208 B.n682 B.n681 163.367
R1209 B.n682 B.n101 163.367
R1210 B.n686 B.n101 163.367
R1211 B.n687 B.n686 163.367
R1212 B.n688 B.n687 163.367
R1213 B.n688 B.n99 163.367
R1214 B.n692 B.n99 163.367
R1215 B.n693 B.n692 163.367
R1216 B.n694 B.n693 163.367
R1217 B.n694 B.n97 163.367
R1218 B.n698 B.n97 163.367
R1219 B.n699 B.n698 163.367
R1220 B.n700 B.n699 163.367
R1221 B.n700 B.n95 163.367
R1222 B.n874 B.n33 163.367
R1223 B.n874 B.n873 163.367
R1224 B.n873 B.n872 163.367
R1225 B.n872 B.n35 163.367
R1226 B.n868 B.n35 163.367
R1227 B.n868 B.n867 163.367
R1228 B.n867 B.n866 163.367
R1229 B.n866 B.n37 163.367
R1230 B.n862 B.n37 163.367
R1231 B.n862 B.n861 163.367
R1232 B.n861 B.n860 163.367
R1233 B.n860 B.n39 163.367
R1234 B.n856 B.n39 163.367
R1235 B.n856 B.n855 163.367
R1236 B.n855 B.n854 163.367
R1237 B.n854 B.n41 163.367
R1238 B.n850 B.n41 163.367
R1239 B.n850 B.n849 163.367
R1240 B.n849 B.n848 163.367
R1241 B.n848 B.n43 163.367
R1242 B.n844 B.n43 163.367
R1243 B.n844 B.n843 163.367
R1244 B.n843 B.n842 163.367
R1245 B.n842 B.n45 163.367
R1246 B.n838 B.n45 163.367
R1247 B.n838 B.n837 163.367
R1248 B.n837 B.n836 163.367
R1249 B.n836 B.n47 163.367
R1250 B.n832 B.n47 163.367
R1251 B.n832 B.n831 163.367
R1252 B.n831 B.n830 163.367
R1253 B.n830 B.n49 163.367
R1254 B.n826 B.n49 163.367
R1255 B.n826 B.n825 163.367
R1256 B.n825 B.n824 163.367
R1257 B.n824 B.n51 163.367
R1258 B.n820 B.n51 163.367
R1259 B.n820 B.n819 163.367
R1260 B.n819 B.n818 163.367
R1261 B.n818 B.n53 163.367
R1262 B.n814 B.n53 163.367
R1263 B.n814 B.n813 163.367
R1264 B.n813 B.n812 163.367
R1265 B.n812 B.n55 163.367
R1266 B.n808 B.n55 163.367
R1267 B.n808 B.n807 163.367
R1268 B.n807 B.n806 163.367
R1269 B.n806 B.n57 163.367
R1270 B.n802 B.n57 163.367
R1271 B.n802 B.n801 163.367
R1272 B.n801 B.n800 163.367
R1273 B.n800 B.n59 163.367
R1274 B.n795 B.n59 163.367
R1275 B.n795 B.n794 163.367
R1276 B.n794 B.n793 163.367
R1277 B.n793 B.n63 163.367
R1278 B.n789 B.n63 163.367
R1279 B.n789 B.n788 163.367
R1280 B.n788 B.n787 163.367
R1281 B.n787 B.n65 163.367
R1282 B.n783 B.n65 163.367
R1283 B.n783 B.n782 163.367
R1284 B.n782 B.n69 163.367
R1285 B.n778 B.n69 163.367
R1286 B.n778 B.n777 163.367
R1287 B.n777 B.n776 163.367
R1288 B.n776 B.n71 163.367
R1289 B.n772 B.n71 163.367
R1290 B.n772 B.n771 163.367
R1291 B.n771 B.n770 163.367
R1292 B.n770 B.n73 163.367
R1293 B.n766 B.n73 163.367
R1294 B.n766 B.n765 163.367
R1295 B.n765 B.n764 163.367
R1296 B.n764 B.n75 163.367
R1297 B.n760 B.n75 163.367
R1298 B.n760 B.n759 163.367
R1299 B.n759 B.n758 163.367
R1300 B.n758 B.n77 163.367
R1301 B.n754 B.n77 163.367
R1302 B.n754 B.n753 163.367
R1303 B.n753 B.n752 163.367
R1304 B.n752 B.n79 163.367
R1305 B.n748 B.n79 163.367
R1306 B.n748 B.n747 163.367
R1307 B.n747 B.n746 163.367
R1308 B.n746 B.n81 163.367
R1309 B.n742 B.n81 163.367
R1310 B.n742 B.n741 163.367
R1311 B.n741 B.n740 163.367
R1312 B.n740 B.n83 163.367
R1313 B.n736 B.n83 163.367
R1314 B.n736 B.n735 163.367
R1315 B.n735 B.n734 163.367
R1316 B.n734 B.n85 163.367
R1317 B.n730 B.n85 163.367
R1318 B.n730 B.n729 163.367
R1319 B.n729 B.n728 163.367
R1320 B.n728 B.n87 163.367
R1321 B.n724 B.n87 163.367
R1322 B.n724 B.n723 163.367
R1323 B.n723 B.n722 163.367
R1324 B.n722 B.n89 163.367
R1325 B.n718 B.n89 163.367
R1326 B.n718 B.n717 163.367
R1327 B.n717 B.n716 163.367
R1328 B.n716 B.n91 163.367
R1329 B.n712 B.n91 163.367
R1330 B.n712 B.n711 163.367
R1331 B.n711 B.n710 163.367
R1332 B.n710 B.n93 163.367
R1333 B.n706 B.n93 163.367
R1334 B.n706 B.n705 163.367
R1335 B.n705 B.n704 163.367
R1336 B.n185 B.t7 110.326
R1337 B.n67 B.t11 110.326
R1338 B.n193 B.t1 110.306
R1339 B.n61 B.t5 110.306
R1340 B.n186 B.n185 59.5399
R1341 B.n421 B.n193 59.5399
R1342 B.n797 B.n61 59.5399
R1343 B.n68 B.n67 59.5399
R1344 B.n185 B.n184 59.152
R1345 B.n193 B.n192 59.152
R1346 B.n61 B.n60 59.152
R1347 B.n67 B.n66 59.152
R1348 B.n877 B.n876 33.8737
R1349 B.n703 B.n702 33.8737
R1350 B.n516 B.n515 33.8737
R1351 B.n342 B.n341 33.8737
R1352 B B.n971 18.0485
R1353 B.n876 B.n875 10.6151
R1354 B.n875 B.n34 10.6151
R1355 B.n871 B.n34 10.6151
R1356 B.n871 B.n870 10.6151
R1357 B.n870 B.n869 10.6151
R1358 B.n869 B.n36 10.6151
R1359 B.n865 B.n36 10.6151
R1360 B.n865 B.n864 10.6151
R1361 B.n864 B.n863 10.6151
R1362 B.n863 B.n38 10.6151
R1363 B.n859 B.n38 10.6151
R1364 B.n859 B.n858 10.6151
R1365 B.n858 B.n857 10.6151
R1366 B.n857 B.n40 10.6151
R1367 B.n853 B.n40 10.6151
R1368 B.n853 B.n852 10.6151
R1369 B.n852 B.n851 10.6151
R1370 B.n851 B.n42 10.6151
R1371 B.n847 B.n42 10.6151
R1372 B.n847 B.n846 10.6151
R1373 B.n846 B.n845 10.6151
R1374 B.n845 B.n44 10.6151
R1375 B.n841 B.n44 10.6151
R1376 B.n841 B.n840 10.6151
R1377 B.n840 B.n839 10.6151
R1378 B.n839 B.n46 10.6151
R1379 B.n835 B.n46 10.6151
R1380 B.n835 B.n834 10.6151
R1381 B.n834 B.n833 10.6151
R1382 B.n833 B.n48 10.6151
R1383 B.n829 B.n48 10.6151
R1384 B.n829 B.n828 10.6151
R1385 B.n828 B.n827 10.6151
R1386 B.n827 B.n50 10.6151
R1387 B.n823 B.n50 10.6151
R1388 B.n823 B.n822 10.6151
R1389 B.n822 B.n821 10.6151
R1390 B.n821 B.n52 10.6151
R1391 B.n817 B.n52 10.6151
R1392 B.n817 B.n816 10.6151
R1393 B.n816 B.n815 10.6151
R1394 B.n815 B.n54 10.6151
R1395 B.n811 B.n54 10.6151
R1396 B.n811 B.n810 10.6151
R1397 B.n810 B.n809 10.6151
R1398 B.n809 B.n56 10.6151
R1399 B.n805 B.n56 10.6151
R1400 B.n805 B.n804 10.6151
R1401 B.n804 B.n803 10.6151
R1402 B.n803 B.n58 10.6151
R1403 B.n799 B.n58 10.6151
R1404 B.n799 B.n798 10.6151
R1405 B.n796 B.n62 10.6151
R1406 B.n792 B.n62 10.6151
R1407 B.n792 B.n791 10.6151
R1408 B.n791 B.n790 10.6151
R1409 B.n790 B.n64 10.6151
R1410 B.n786 B.n64 10.6151
R1411 B.n786 B.n785 10.6151
R1412 B.n785 B.n784 10.6151
R1413 B.n781 B.n780 10.6151
R1414 B.n780 B.n779 10.6151
R1415 B.n779 B.n70 10.6151
R1416 B.n775 B.n70 10.6151
R1417 B.n775 B.n774 10.6151
R1418 B.n774 B.n773 10.6151
R1419 B.n773 B.n72 10.6151
R1420 B.n769 B.n72 10.6151
R1421 B.n769 B.n768 10.6151
R1422 B.n768 B.n767 10.6151
R1423 B.n767 B.n74 10.6151
R1424 B.n763 B.n74 10.6151
R1425 B.n763 B.n762 10.6151
R1426 B.n762 B.n761 10.6151
R1427 B.n761 B.n76 10.6151
R1428 B.n757 B.n76 10.6151
R1429 B.n757 B.n756 10.6151
R1430 B.n756 B.n755 10.6151
R1431 B.n755 B.n78 10.6151
R1432 B.n751 B.n78 10.6151
R1433 B.n751 B.n750 10.6151
R1434 B.n750 B.n749 10.6151
R1435 B.n749 B.n80 10.6151
R1436 B.n745 B.n80 10.6151
R1437 B.n745 B.n744 10.6151
R1438 B.n744 B.n743 10.6151
R1439 B.n743 B.n82 10.6151
R1440 B.n739 B.n82 10.6151
R1441 B.n739 B.n738 10.6151
R1442 B.n738 B.n737 10.6151
R1443 B.n737 B.n84 10.6151
R1444 B.n733 B.n84 10.6151
R1445 B.n733 B.n732 10.6151
R1446 B.n732 B.n731 10.6151
R1447 B.n731 B.n86 10.6151
R1448 B.n727 B.n86 10.6151
R1449 B.n727 B.n726 10.6151
R1450 B.n726 B.n725 10.6151
R1451 B.n725 B.n88 10.6151
R1452 B.n721 B.n88 10.6151
R1453 B.n721 B.n720 10.6151
R1454 B.n720 B.n719 10.6151
R1455 B.n719 B.n90 10.6151
R1456 B.n715 B.n90 10.6151
R1457 B.n715 B.n714 10.6151
R1458 B.n714 B.n713 10.6151
R1459 B.n713 B.n92 10.6151
R1460 B.n709 B.n92 10.6151
R1461 B.n709 B.n708 10.6151
R1462 B.n708 B.n707 10.6151
R1463 B.n707 B.n94 10.6151
R1464 B.n703 B.n94 10.6151
R1465 B.n517 B.n516 10.6151
R1466 B.n517 B.n156 10.6151
R1467 B.n521 B.n156 10.6151
R1468 B.n522 B.n521 10.6151
R1469 B.n523 B.n522 10.6151
R1470 B.n523 B.n154 10.6151
R1471 B.n527 B.n154 10.6151
R1472 B.n528 B.n527 10.6151
R1473 B.n529 B.n528 10.6151
R1474 B.n529 B.n152 10.6151
R1475 B.n533 B.n152 10.6151
R1476 B.n534 B.n533 10.6151
R1477 B.n535 B.n534 10.6151
R1478 B.n535 B.n150 10.6151
R1479 B.n539 B.n150 10.6151
R1480 B.n540 B.n539 10.6151
R1481 B.n541 B.n540 10.6151
R1482 B.n541 B.n148 10.6151
R1483 B.n545 B.n148 10.6151
R1484 B.n546 B.n545 10.6151
R1485 B.n547 B.n546 10.6151
R1486 B.n547 B.n146 10.6151
R1487 B.n551 B.n146 10.6151
R1488 B.n552 B.n551 10.6151
R1489 B.n553 B.n552 10.6151
R1490 B.n553 B.n144 10.6151
R1491 B.n557 B.n144 10.6151
R1492 B.n558 B.n557 10.6151
R1493 B.n559 B.n558 10.6151
R1494 B.n559 B.n142 10.6151
R1495 B.n563 B.n142 10.6151
R1496 B.n564 B.n563 10.6151
R1497 B.n565 B.n564 10.6151
R1498 B.n565 B.n140 10.6151
R1499 B.n569 B.n140 10.6151
R1500 B.n570 B.n569 10.6151
R1501 B.n571 B.n570 10.6151
R1502 B.n571 B.n138 10.6151
R1503 B.n575 B.n138 10.6151
R1504 B.n576 B.n575 10.6151
R1505 B.n577 B.n576 10.6151
R1506 B.n577 B.n136 10.6151
R1507 B.n581 B.n136 10.6151
R1508 B.n582 B.n581 10.6151
R1509 B.n583 B.n582 10.6151
R1510 B.n583 B.n134 10.6151
R1511 B.n587 B.n134 10.6151
R1512 B.n588 B.n587 10.6151
R1513 B.n589 B.n588 10.6151
R1514 B.n589 B.n132 10.6151
R1515 B.n593 B.n132 10.6151
R1516 B.n594 B.n593 10.6151
R1517 B.n595 B.n594 10.6151
R1518 B.n595 B.n130 10.6151
R1519 B.n599 B.n130 10.6151
R1520 B.n600 B.n599 10.6151
R1521 B.n601 B.n600 10.6151
R1522 B.n601 B.n128 10.6151
R1523 B.n605 B.n128 10.6151
R1524 B.n606 B.n605 10.6151
R1525 B.n607 B.n606 10.6151
R1526 B.n607 B.n126 10.6151
R1527 B.n611 B.n126 10.6151
R1528 B.n612 B.n611 10.6151
R1529 B.n613 B.n612 10.6151
R1530 B.n613 B.n124 10.6151
R1531 B.n617 B.n124 10.6151
R1532 B.n618 B.n617 10.6151
R1533 B.n619 B.n618 10.6151
R1534 B.n619 B.n122 10.6151
R1535 B.n623 B.n122 10.6151
R1536 B.n624 B.n623 10.6151
R1537 B.n625 B.n624 10.6151
R1538 B.n625 B.n120 10.6151
R1539 B.n629 B.n120 10.6151
R1540 B.n630 B.n629 10.6151
R1541 B.n631 B.n630 10.6151
R1542 B.n631 B.n118 10.6151
R1543 B.n635 B.n118 10.6151
R1544 B.n636 B.n635 10.6151
R1545 B.n637 B.n636 10.6151
R1546 B.n637 B.n116 10.6151
R1547 B.n641 B.n116 10.6151
R1548 B.n642 B.n641 10.6151
R1549 B.n643 B.n642 10.6151
R1550 B.n643 B.n114 10.6151
R1551 B.n647 B.n114 10.6151
R1552 B.n648 B.n647 10.6151
R1553 B.n649 B.n648 10.6151
R1554 B.n649 B.n112 10.6151
R1555 B.n653 B.n112 10.6151
R1556 B.n654 B.n653 10.6151
R1557 B.n655 B.n654 10.6151
R1558 B.n655 B.n110 10.6151
R1559 B.n659 B.n110 10.6151
R1560 B.n660 B.n659 10.6151
R1561 B.n661 B.n660 10.6151
R1562 B.n661 B.n108 10.6151
R1563 B.n665 B.n108 10.6151
R1564 B.n666 B.n665 10.6151
R1565 B.n667 B.n666 10.6151
R1566 B.n667 B.n106 10.6151
R1567 B.n671 B.n106 10.6151
R1568 B.n672 B.n671 10.6151
R1569 B.n673 B.n672 10.6151
R1570 B.n673 B.n104 10.6151
R1571 B.n677 B.n104 10.6151
R1572 B.n678 B.n677 10.6151
R1573 B.n679 B.n678 10.6151
R1574 B.n679 B.n102 10.6151
R1575 B.n683 B.n102 10.6151
R1576 B.n684 B.n683 10.6151
R1577 B.n685 B.n684 10.6151
R1578 B.n685 B.n100 10.6151
R1579 B.n689 B.n100 10.6151
R1580 B.n690 B.n689 10.6151
R1581 B.n691 B.n690 10.6151
R1582 B.n691 B.n98 10.6151
R1583 B.n695 B.n98 10.6151
R1584 B.n696 B.n695 10.6151
R1585 B.n697 B.n696 10.6151
R1586 B.n697 B.n96 10.6151
R1587 B.n701 B.n96 10.6151
R1588 B.n702 B.n701 10.6151
R1589 B.n343 B.n342 10.6151
R1590 B.n343 B.n218 10.6151
R1591 B.n347 B.n218 10.6151
R1592 B.n348 B.n347 10.6151
R1593 B.n349 B.n348 10.6151
R1594 B.n349 B.n216 10.6151
R1595 B.n353 B.n216 10.6151
R1596 B.n354 B.n353 10.6151
R1597 B.n355 B.n354 10.6151
R1598 B.n355 B.n214 10.6151
R1599 B.n359 B.n214 10.6151
R1600 B.n360 B.n359 10.6151
R1601 B.n361 B.n360 10.6151
R1602 B.n361 B.n212 10.6151
R1603 B.n365 B.n212 10.6151
R1604 B.n366 B.n365 10.6151
R1605 B.n367 B.n366 10.6151
R1606 B.n367 B.n210 10.6151
R1607 B.n371 B.n210 10.6151
R1608 B.n372 B.n371 10.6151
R1609 B.n373 B.n372 10.6151
R1610 B.n373 B.n208 10.6151
R1611 B.n377 B.n208 10.6151
R1612 B.n378 B.n377 10.6151
R1613 B.n379 B.n378 10.6151
R1614 B.n379 B.n206 10.6151
R1615 B.n383 B.n206 10.6151
R1616 B.n384 B.n383 10.6151
R1617 B.n385 B.n384 10.6151
R1618 B.n385 B.n204 10.6151
R1619 B.n389 B.n204 10.6151
R1620 B.n390 B.n389 10.6151
R1621 B.n391 B.n390 10.6151
R1622 B.n391 B.n202 10.6151
R1623 B.n395 B.n202 10.6151
R1624 B.n396 B.n395 10.6151
R1625 B.n397 B.n396 10.6151
R1626 B.n397 B.n200 10.6151
R1627 B.n401 B.n200 10.6151
R1628 B.n402 B.n401 10.6151
R1629 B.n403 B.n402 10.6151
R1630 B.n403 B.n198 10.6151
R1631 B.n407 B.n198 10.6151
R1632 B.n408 B.n407 10.6151
R1633 B.n409 B.n408 10.6151
R1634 B.n409 B.n196 10.6151
R1635 B.n413 B.n196 10.6151
R1636 B.n414 B.n413 10.6151
R1637 B.n415 B.n414 10.6151
R1638 B.n415 B.n194 10.6151
R1639 B.n419 B.n194 10.6151
R1640 B.n420 B.n419 10.6151
R1641 B.n422 B.n190 10.6151
R1642 B.n426 B.n190 10.6151
R1643 B.n427 B.n426 10.6151
R1644 B.n428 B.n427 10.6151
R1645 B.n428 B.n188 10.6151
R1646 B.n432 B.n188 10.6151
R1647 B.n433 B.n432 10.6151
R1648 B.n434 B.n433 10.6151
R1649 B.n438 B.n437 10.6151
R1650 B.n439 B.n438 10.6151
R1651 B.n439 B.n182 10.6151
R1652 B.n443 B.n182 10.6151
R1653 B.n444 B.n443 10.6151
R1654 B.n445 B.n444 10.6151
R1655 B.n445 B.n180 10.6151
R1656 B.n449 B.n180 10.6151
R1657 B.n450 B.n449 10.6151
R1658 B.n451 B.n450 10.6151
R1659 B.n451 B.n178 10.6151
R1660 B.n455 B.n178 10.6151
R1661 B.n456 B.n455 10.6151
R1662 B.n457 B.n456 10.6151
R1663 B.n457 B.n176 10.6151
R1664 B.n461 B.n176 10.6151
R1665 B.n462 B.n461 10.6151
R1666 B.n463 B.n462 10.6151
R1667 B.n463 B.n174 10.6151
R1668 B.n467 B.n174 10.6151
R1669 B.n468 B.n467 10.6151
R1670 B.n469 B.n468 10.6151
R1671 B.n469 B.n172 10.6151
R1672 B.n473 B.n172 10.6151
R1673 B.n474 B.n473 10.6151
R1674 B.n475 B.n474 10.6151
R1675 B.n475 B.n170 10.6151
R1676 B.n479 B.n170 10.6151
R1677 B.n480 B.n479 10.6151
R1678 B.n481 B.n480 10.6151
R1679 B.n481 B.n168 10.6151
R1680 B.n485 B.n168 10.6151
R1681 B.n486 B.n485 10.6151
R1682 B.n487 B.n486 10.6151
R1683 B.n487 B.n166 10.6151
R1684 B.n491 B.n166 10.6151
R1685 B.n492 B.n491 10.6151
R1686 B.n493 B.n492 10.6151
R1687 B.n493 B.n164 10.6151
R1688 B.n497 B.n164 10.6151
R1689 B.n498 B.n497 10.6151
R1690 B.n499 B.n498 10.6151
R1691 B.n499 B.n162 10.6151
R1692 B.n503 B.n162 10.6151
R1693 B.n504 B.n503 10.6151
R1694 B.n505 B.n504 10.6151
R1695 B.n505 B.n160 10.6151
R1696 B.n509 B.n160 10.6151
R1697 B.n510 B.n509 10.6151
R1698 B.n511 B.n510 10.6151
R1699 B.n511 B.n158 10.6151
R1700 B.n515 B.n158 10.6151
R1701 B.n341 B.n220 10.6151
R1702 B.n337 B.n220 10.6151
R1703 B.n337 B.n336 10.6151
R1704 B.n336 B.n335 10.6151
R1705 B.n335 B.n222 10.6151
R1706 B.n331 B.n222 10.6151
R1707 B.n331 B.n330 10.6151
R1708 B.n330 B.n329 10.6151
R1709 B.n329 B.n224 10.6151
R1710 B.n325 B.n224 10.6151
R1711 B.n325 B.n324 10.6151
R1712 B.n324 B.n323 10.6151
R1713 B.n323 B.n226 10.6151
R1714 B.n319 B.n226 10.6151
R1715 B.n319 B.n318 10.6151
R1716 B.n318 B.n317 10.6151
R1717 B.n317 B.n228 10.6151
R1718 B.n313 B.n228 10.6151
R1719 B.n313 B.n312 10.6151
R1720 B.n312 B.n311 10.6151
R1721 B.n311 B.n230 10.6151
R1722 B.n307 B.n230 10.6151
R1723 B.n307 B.n306 10.6151
R1724 B.n306 B.n305 10.6151
R1725 B.n305 B.n232 10.6151
R1726 B.n301 B.n232 10.6151
R1727 B.n301 B.n300 10.6151
R1728 B.n300 B.n299 10.6151
R1729 B.n299 B.n234 10.6151
R1730 B.n295 B.n234 10.6151
R1731 B.n295 B.n294 10.6151
R1732 B.n294 B.n293 10.6151
R1733 B.n293 B.n236 10.6151
R1734 B.n289 B.n236 10.6151
R1735 B.n289 B.n288 10.6151
R1736 B.n288 B.n287 10.6151
R1737 B.n287 B.n238 10.6151
R1738 B.n283 B.n238 10.6151
R1739 B.n283 B.n282 10.6151
R1740 B.n282 B.n281 10.6151
R1741 B.n281 B.n240 10.6151
R1742 B.n277 B.n240 10.6151
R1743 B.n277 B.n276 10.6151
R1744 B.n276 B.n275 10.6151
R1745 B.n275 B.n242 10.6151
R1746 B.n271 B.n242 10.6151
R1747 B.n271 B.n270 10.6151
R1748 B.n270 B.n269 10.6151
R1749 B.n269 B.n244 10.6151
R1750 B.n265 B.n244 10.6151
R1751 B.n265 B.n264 10.6151
R1752 B.n264 B.n263 10.6151
R1753 B.n263 B.n246 10.6151
R1754 B.n259 B.n246 10.6151
R1755 B.n259 B.n258 10.6151
R1756 B.n258 B.n257 10.6151
R1757 B.n257 B.n248 10.6151
R1758 B.n253 B.n248 10.6151
R1759 B.n253 B.n252 10.6151
R1760 B.n252 B.n251 10.6151
R1761 B.n251 B.n0 10.6151
R1762 B.n967 B.n1 10.6151
R1763 B.n967 B.n966 10.6151
R1764 B.n966 B.n965 10.6151
R1765 B.n965 B.n4 10.6151
R1766 B.n961 B.n4 10.6151
R1767 B.n961 B.n960 10.6151
R1768 B.n960 B.n959 10.6151
R1769 B.n959 B.n6 10.6151
R1770 B.n955 B.n6 10.6151
R1771 B.n955 B.n954 10.6151
R1772 B.n954 B.n953 10.6151
R1773 B.n953 B.n8 10.6151
R1774 B.n949 B.n8 10.6151
R1775 B.n949 B.n948 10.6151
R1776 B.n948 B.n947 10.6151
R1777 B.n947 B.n10 10.6151
R1778 B.n943 B.n10 10.6151
R1779 B.n943 B.n942 10.6151
R1780 B.n942 B.n941 10.6151
R1781 B.n941 B.n12 10.6151
R1782 B.n937 B.n12 10.6151
R1783 B.n937 B.n936 10.6151
R1784 B.n936 B.n935 10.6151
R1785 B.n935 B.n14 10.6151
R1786 B.n931 B.n14 10.6151
R1787 B.n931 B.n930 10.6151
R1788 B.n930 B.n929 10.6151
R1789 B.n929 B.n16 10.6151
R1790 B.n925 B.n16 10.6151
R1791 B.n925 B.n924 10.6151
R1792 B.n924 B.n923 10.6151
R1793 B.n923 B.n18 10.6151
R1794 B.n919 B.n18 10.6151
R1795 B.n919 B.n918 10.6151
R1796 B.n918 B.n917 10.6151
R1797 B.n917 B.n20 10.6151
R1798 B.n913 B.n20 10.6151
R1799 B.n913 B.n912 10.6151
R1800 B.n912 B.n911 10.6151
R1801 B.n911 B.n22 10.6151
R1802 B.n907 B.n22 10.6151
R1803 B.n907 B.n906 10.6151
R1804 B.n906 B.n905 10.6151
R1805 B.n905 B.n24 10.6151
R1806 B.n901 B.n24 10.6151
R1807 B.n901 B.n900 10.6151
R1808 B.n900 B.n899 10.6151
R1809 B.n899 B.n26 10.6151
R1810 B.n895 B.n26 10.6151
R1811 B.n895 B.n894 10.6151
R1812 B.n894 B.n893 10.6151
R1813 B.n893 B.n28 10.6151
R1814 B.n889 B.n28 10.6151
R1815 B.n889 B.n888 10.6151
R1816 B.n888 B.n887 10.6151
R1817 B.n887 B.n30 10.6151
R1818 B.n883 B.n30 10.6151
R1819 B.n883 B.n882 10.6151
R1820 B.n882 B.n881 10.6151
R1821 B.n881 B.n32 10.6151
R1822 B.n877 B.n32 10.6151
R1823 B.n797 B.n796 6.5566
R1824 B.n784 B.n68 6.5566
R1825 B.n422 B.n421 6.5566
R1826 B.n434 B.n186 6.5566
R1827 B.n798 B.n797 4.05904
R1828 B.n781 B.n68 4.05904
R1829 B.n421 B.n420 4.05904
R1830 B.n437 B.n186 4.05904
R1831 B.n971 B.n0 2.81026
R1832 B.n971 B.n1 2.81026
C0 VN VDD1 0.153704f
C1 VP B 2.37776f
C2 VN B 1.36283f
C3 w_n4630_n4136# VDD2 3.24606f
C4 VTAIL VDD2 12.2052f
C5 VDD1 w_n4630_n4136# 3.09628f
C6 VTAIL VDD1 12.154099f
C7 VP VN 9.279769f
C8 w_n4630_n4136# B 11.8255f
C9 VTAIL B 4.64766f
C10 VDD1 VDD2 2.25111f
C11 VP w_n4630_n4136# 10.607599f
C12 VP VTAIL 14.5799f
C13 VDD2 B 2.95421f
C14 VN w_n4630_n4136# 10.0044f
C15 VN VTAIL 14.5655f
C16 VDD1 B 2.83162f
C17 VP VDD2 0.599252f
C18 VTAIL w_n4630_n4136# 3.75198f
C19 VN VDD2 14.047501f
C20 VP VDD1 14.488501f
C21 VDD2 VSUBS 2.28681f
C22 VDD1 VSUBS 2.110595f
C23 VTAIL VSUBS 1.45408f
C24 VN VSUBS 8.00163f
C25 VP VSUBS 4.522943f
C26 B VSUBS 5.840923f
C27 w_n4630_n4136# VSUBS 0.23463p
C28 B.n0 VSUBS 0.005313f
C29 B.n1 VSUBS 0.005313f
C30 B.n2 VSUBS 0.008402f
C31 B.n3 VSUBS 0.008402f
C32 B.n4 VSUBS 0.008402f
C33 B.n5 VSUBS 0.008402f
C34 B.n6 VSUBS 0.008402f
C35 B.n7 VSUBS 0.008402f
C36 B.n8 VSUBS 0.008402f
C37 B.n9 VSUBS 0.008402f
C38 B.n10 VSUBS 0.008402f
C39 B.n11 VSUBS 0.008402f
C40 B.n12 VSUBS 0.008402f
C41 B.n13 VSUBS 0.008402f
C42 B.n14 VSUBS 0.008402f
C43 B.n15 VSUBS 0.008402f
C44 B.n16 VSUBS 0.008402f
C45 B.n17 VSUBS 0.008402f
C46 B.n18 VSUBS 0.008402f
C47 B.n19 VSUBS 0.008402f
C48 B.n20 VSUBS 0.008402f
C49 B.n21 VSUBS 0.008402f
C50 B.n22 VSUBS 0.008402f
C51 B.n23 VSUBS 0.008402f
C52 B.n24 VSUBS 0.008402f
C53 B.n25 VSUBS 0.008402f
C54 B.n26 VSUBS 0.008402f
C55 B.n27 VSUBS 0.008402f
C56 B.n28 VSUBS 0.008402f
C57 B.n29 VSUBS 0.008402f
C58 B.n30 VSUBS 0.008402f
C59 B.n31 VSUBS 0.008402f
C60 B.n32 VSUBS 0.008402f
C61 B.n33 VSUBS 0.020386f
C62 B.n34 VSUBS 0.008402f
C63 B.n35 VSUBS 0.008402f
C64 B.n36 VSUBS 0.008402f
C65 B.n37 VSUBS 0.008402f
C66 B.n38 VSUBS 0.008402f
C67 B.n39 VSUBS 0.008402f
C68 B.n40 VSUBS 0.008402f
C69 B.n41 VSUBS 0.008402f
C70 B.n42 VSUBS 0.008402f
C71 B.n43 VSUBS 0.008402f
C72 B.n44 VSUBS 0.008402f
C73 B.n45 VSUBS 0.008402f
C74 B.n46 VSUBS 0.008402f
C75 B.n47 VSUBS 0.008402f
C76 B.n48 VSUBS 0.008402f
C77 B.n49 VSUBS 0.008402f
C78 B.n50 VSUBS 0.008402f
C79 B.n51 VSUBS 0.008402f
C80 B.n52 VSUBS 0.008402f
C81 B.n53 VSUBS 0.008402f
C82 B.n54 VSUBS 0.008402f
C83 B.n55 VSUBS 0.008402f
C84 B.n56 VSUBS 0.008402f
C85 B.n57 VSUBS 0.008402f
C86 B.n58 VSUBS 0.008402f
C87 B.n59 VSUBS 0.008402f
C88 B.t5 VSUBS 0.635793f
C89 B.t4 VSUBS 0.661989f
C90 B.t3 VSUBS 2.32141f
C91 B.n60 VSUBS 0.361251f
C92 B.n61 VSUBS 0.087031f
C93 B.n62 VSUBS 0.008402f
C94 B.n63 VSUBS 0.008402f
C95 B.n64 VSUBS 0.008402f
C96 B.n65 VSUBS 0.008402f
C97 B.t11 VSUBS 0.635773f
C98 B.t10 VSUBS 0.661973f
C99 B.t9 VSUBS 2.32141f
C100 B.n66 VSUBS 0.361266f
C101 B.n67 VSUBS 0.08705f
C102 B.n68 VSUBS 0.019467f
C103 B.n69 VSUBS 0.008402f
C104 B.n70 VSUBS 0.008402f
C105 B.n71 VSUBS 0.008402f
C106 B.n72 VSUBS 0.008402f
C107 B.n73 VSUBS 0.008402f
C108 B.n74 VSUBS 0.008402f
C109 B.n75 VSUBS 0.008402f
C110 B.n76 VSUBS 0.008402f
C111 B.n77 VSUBS 0.008402f
C112 B.n78 VSUBS 0.008402f
C113 B.n79 VSUBS 0.008402f
C114 B.n80 VSUBS 0.008402f
C115 B.n81 VSUBS 0.008402f
C116 B.n82 VSUBS 0.008402f
C117 B.n83 VSUBS 0.008402f
C118 B.n84 VSUBS 0.008402f
C119 B.n85 VSUBS 0.008402f
C120 B.n86 VSUBS 0.008402f
C121 B.n87 VSUBS 0.008402f
C122 B.n88 VSUBS 0.008402f
C123 B.n89 VSUBS 0.008402f
C124 B.n90 VSUBS 0.008402f
C125 B.n91 VSUBS 0.008402f
C126 B.n92 VSUBS 0.008402f
C127 B.n93 VSUBS 0.008402f
C128 B.n94 VSUBS 0.008402f
C129 B.n95 VSUBS 0.019896f
C130 B.n96 VSUBS 0.008402f
C131 B.n97 VSUBS 0.008402f
C132 B.n98 VSUBS 0.008402f
C133 B.n99 VSUBS 0.008402f
C134 B.n100 VSUBS 0.008402f
C135 B.n101 VSUBS 0.008402f
C136 B.n102 VSUBS 0.008402f
C137 B.n103 VSUBS 0.008402f
C138 B.n104 VSUBS 0.008402f
C139 B.n105 VSUBS 0.008402f
C140 B.n106 VSUBS 0.008402f
C141 B.n107 VSUBS 0.008402f
C142 B.n108 VSUBS 0.008402f
C143 B.n109 VSUBS 0.008402f
C144 B.n110 VSUBS 0.008402f
C145 B.n111 VSUBS 0.008402f
C146 B.n112 VSUBS 0.008402f
C147 B.n113 VSUBS 0.008402f
C148 B.n114 VSUBS 0.008402f
C149 B.n115 VSUBS 0.008402f
C150 B.n116 VSUBS 0.008402f
C151 B.n117 VSUBS 0.008402f
C152 B.n118 VSUBS 0.008402f
C153 B.n119 VSUBS 0.008402f
C154 B.n120 VSUBS 0.008402f
C155 B.n121 VSUBS 0.008402f
C156 B.n122 VSUBS 0.008402f
C157 B.n123 VSUBS 0.008402f
C158 B.n124 VSUBS 0.008402f
C159 B.n125 VSUBS 0.008402f
C160 B.n126 VSUBS 0.008402f
C161 B.n127 VSUBS 0.008402f
C162 B.n128 VSUBS 0.008402f
C163 B.n129 VSUBS 0.008402f
C164 B.n130 VSUBS 0.008402f
C165 B.n131 VSUBS 0.008402f
C166 B.n132 VSUBS 0.008402f
C167 B.n133 VSUBS 0.008402f
C168 B.n134 VSUBS 0.008402f
C169 B.n135 VSUBS 0.008402f
C170 B.n136 VSUBS 0.008402f
C171 B.n137 VSUBS 0.008402f
C172 B.n138 VSUBS 0.008402f
C173 B.n139 VSUBS 0.008402f
C174 B.n140 VSUBS 0.008402f
C175 B.n141 VSUBS 0.008402f
C176 B.n142 VSUBS 0.008402f
C177 B.n143 VSUBS 0.008402f
C178 B.n144 VSUBS 0.008402f
C179 B.n145 VSUBS 0.008402f
C180 B.n146 VSUBS 0.008402f
C181 B.n147 VSUBS 0.008402f
C182 B.n148 VSUBS 0.008402f
C183 B.n149 VSUBS 0.008402f
C184 B.n150 VSUBS 0.008402f
C185 B.n151 VSUBS 0.008402f
C186 B.n152 VSUBS 0.008402f
C187 B.n153 VSUBS 0.008402f
C188 B.n154 VSUBS 0.008402f
C189 B.n155 VSUBS 0.008402f
C190 B.n156 VSUBS 0.008402f
C191 B.n157 VSUBS 0.019896f
C192 B.n158 VSUBS 0.008402f
C193 B.n159 VSUBS 0.008402f
C194 B.n160 VSUBS 0.008402f
C195 B.n161 VSUBS 0.008402f
C196 B.n162 VSUBS 0.008402f
C197 B.n163 VSUBS 0.008402f
C198 B.n164 VSUBS 0.008402f
C199 B.n165 VSUBS 0.008402f
C200 B.n166 VSUBS 0.008402f
C201 B.n167 VSUBS 0.008402f
C202 B.n168 VSUBS 0.008402f
C203 B.n169 VSUBS 0.008402f
C204 B.n170 VSUBS 0.008402f
C205 B.n171 VSUBS 0.008402f
C206 B.n172 VSUBS 0.008402f
C207 B.n173 VSUBS 0.008402f
C208 B.n174 VSUBS 0.008402f
C209 B.n175 VSUBS 0.008402f
C210 B.n176 VSUBS 0.008402f
C211 B.n177 VSUBS 0.008402f
C212 B.n178 VSUBS 0.008402f
C213 B.n179 VSUBS 0.008402f
C214 B.n180 VSUBS 0.008402f
C215 B.n181 VSUBS 0.008402f
C216 B.n182 VSUBS 0.008402f
C217 B.n183 VSUBS 0.008402f
C218 B.t7 VSUBS 0.635773f
C219 B.t8 VSUBS 0.661973f
C220 B.t6 VSUBS 2.32141f
C221 B.n184 VSUBS 0.361266f
C222 B.n185 VSUBS 0.08705f
C223 B.n186 VSUBS 0.019467f
C224 B.n187 VSUBS 0.008402f
C225 B.n188 VSUBS 0.008402f
C226 B.n189 VSUBS 0.008402f
C227 B.n190 VSUBS 0.008402f
C228 B.n191 VSUBS 0.008402f
C229 B.t1 VSUBS 0.635793f
C230 B.t2 VSUBS 0.661989f
C231 B.t0 VSUBS 2.32141f
C232 B.n192 VSUBS 0.361251f
C233 B.n193 VSUBS 0.087031f
C234 B.n194 VSUBS 0.008402f
C235 B.n195 VSUBS 0.008402f
C236 B.n196 VSUBS 0.008402f
C237 B.n197 VSUBS 0.008402f
C238 B.n198 VSUBS 0.008402f
C239 B.n199 VSUBS 0.008402f
C240 B.n200 VSUBS 0.008402f
C241 B.n201 VSUBS 0.008402f
C242 B.n202 VSUBS 0.008402f
C243 B.n203 VSUBS 0.008402f
C244 B.n204 VSUBS 0.008402f
C245 B.n205 VSUBS 0.008402f
C246 B.n206 VSUBS 0.008402f
C247 B.n207 VSUBS 0.008402f
C248 B.n208 VSUBS 0.008402f
C249 B.n209 VSUBS 0.008402f
C250 B.n210 VSUBS 0.008402f
C251 B.n211 VSUBS 0.008402f
C252 B.n212 VSUBS 0.008402f
C253 B.n213 VSUBS 0.008402f
C254 B.n214 VSUBS 0.008402f
C255 B.n215 VSUBS 0.008402f
C256 B.n216 VSUBS 0.008402f
C257 B.n217 VSUBS 0.008402f
C258 B.n218 VSUBS 0.008402f
C259 B.n219 VSUBS 0.020386f
C260 B.n220 VSUBS 0.008402f
C261 B.n221 VSUBS 0.008402f
C262 B.n222 VSUBS 0.008402f
C263 B.n223 VSUBS 0.008402f
C264 B.n224 VSUBS 0.008402f
C265 B.n225 VSUBS 0.008402f
C266 B.n226 VSUBS 0.008402f
C267 B.n227 VSUBS 0.008402f
C268 B.n228 VSUBS 0.008402f
C269 B.n229 VSUBS 0.008402f
C270 B.n230 VSUBS 0.008402f
C271 B.n231 VSUBS 0.008402f
C272 B.n232 VSUBS 0.008402f
C273 B.n233 VSUBS 0.008402f
C274 B.n234 VSUBS 0.008402f
C275 B.n235 VSUBS 0.008402f
C276 B.n236 VSUBS 0.008402f
C277 B.n237 VSUBS 0.008402f
C278 B.n238 VSUBS 0.008402f
C279 B.n239 VSUBS 0.008402f
C280 B.n240 VSUBS 0.008402f
C281 B.n241 VSUBS 0.008402f
C282 B.n242 VSUBS 0.008402f
C283 B.n243 VSUBS 0.008402f
C284 B.n244 VSUBS 0.008402f
C285 B.n245 VSUBS 0.008402f
C286 B.n246 VSUBS 0.008402f
C287 B.n247 VSUBS 0.008402f
C288 B.n248 VSUBS 0.008402f
C289 B.n249 VSUBS 0.008402f
C290 B.n250 VSUBS 0.008402f
C291 B.n251 VSUBS 0.008402f
C292 B.n252 VSUBS 0.008402f
C293 B.n253 VSUBS 0.008402f
C294 B.n254 VSUBS 0.008402f
C295 B.n255 VSUBS 0.008402f
C296 B.n256 VSUBS 0.008402f
C297 B.n257 VSUBS 0.008402f
C298 B.n258 VSUBS 0.008402f
C299 B.n259 VSUBS 0.008402f
C300 B.n260 VSUBS 0.008402f
C301 B.n261 VSUBS 0.008402f
C302 B.n262 VSUBS 0.008402f
C303 B.n263 VSUBS 0.008402f
C304 B.n264 VSUBS 0.008402f
C305 B.n265 VSUBS 0.008402f
C306 B.n266 VSUBS 0.008402f
C307 B.n267 VSUBS 0.008402f
C308 B.n268 VSUBS 0.008402f
C309 B.n269 VSUBS 0.008402f
C310 B.n270 VSUBS 0.008402f
C311 B.n271 VSUBS 0.008402f
C312 B.n272 VSUBS 0.008402f
C313 B.n273 VSUBS 0.008402f
C314 B.n274 VSUBS 0.008402f
C315 B.n275 VSUBS 0.008402f
C316 B.n276 VSUBS 0.008402f
C317 B.n277 VSUBS 0.008402f
C318 B.n278 VSUBS 0.008402f
C319 B.n279 VSUBS 0.008402f
C320 B.n280 VSUBS 0.008402f
C321 B.n281 VSUBS 0.008402f
C322 B.n282 VSUBS 0.008402f
C323 B.n283 VSUBS 0.008402f
C324 B.n284 VSUBS 0.008402f
C325 B.n285 VSUBS 0.008402f
C326 B.n286 VSUBS 0.008402f
C327 B.n287 VSUBS 0.008402f
C328 B.n288 VSUBS 0.008402f
C329 B.n289 VSUBS 0.008402f
C330 B.n290 VSUBS 0.008402f
C331 B.n291 VSUBS 0.008402f
C332 B.n292 VSUBS 0.008402f
C333 B.n293 VSUBS 0.008402f
C334 B.n294 VSUBS 0.008402f
C335 B.n295 VSUBS 0.008402f
C336 B.n296 VSUBS 0.008402f
C337 B.n297 VSUBS 0.008402f
C338 B.n298 VSUBS 0.008402f
C339 B.n299 VSUBS 0.008402f
C340 B.n300 VSUBS 0.008402f
C341 B.n301 VSUBS 0.008402f
C342 B.n302 VSUBS 0.008402f
C343 B.n303 VSUBS 0.008402f
C344 B.n304 VSUBS 0.008402f
C345 B.n305 VSUBS 0.008402f
C346 B.n306 VSUBS 0.008402f
C347 B.n307 VSUBS 0.008402f
C348 B.n308 VSUBS 0.008402f
C349 B.n309 VSUBS 0.008402f
C350 B.n310 VSUBS 0.008402f
C351 B.n311 VSUBS 0.008402f
C352 B.n312 VSUBS 0.008402f
C353 B.n313 VSUBS 0.008402f
C354 B.n314 VSUBS 0.008402f
C355 B.n315 VSUBS 0.008402f
C356 B.n316 VSUBS 0.008402f
C357 B.n317 VSUBS 0.008402f
C358 B.n318 VSUBS 0.008402f
C359 B.n319 VSUBS 0.008402f
C360 B.n320 VSUBS 0.008402f
C361 B.n321 VSUBS 0.008402f
C362 B.n322 VSUBS 0.008402f
C363 B.n323 VSUBS 0.008402f
C364 B.n324 VSUBS 0.008402f
C365 B.n325 VSUBS 0.008402f
C366 B.n326 VSUBS 0.008402f
C367 B.n327 VSUBS 0.008402f
C368 B.n328 VSUBS 0.008402f
C369 B.n329 VSUBS 0.008402f
C370 B.n330 VSUBS 0.008402f
C371 B.n331 VSUBS 0.008402f
C372 B.n332 VSUBS 0.008402f
C373 B.n333 VSUBS 0.008402f
C374 B.n334 VSUBS 0.008402f
C375 B.n335 VSUBS 0.008402f
C376 B.n336 VSUBS 0.008402f
C377 B.n337 VSUBS 0.008402f
C378 B.n338 VSUBS 0.008402f
C379 B.n339 VSUBS 0.008402f
C380 B.n340 VSUBS 0.019896f
C381 B.n341 VSUBS 0.019896f
C382 B.n342 VSUBS 0.020386f
C383 B.n343 VSUBS 0.008402f
C384 B.n344 VSUBS 0.008402f
C385 B.n345 VSUBS 0.008402f
C386 B.n346 VSUBS 0.008402f
C387 B.n347 VSUBS 0.008402f
C388 B.n348 VSUBS 0.008402f
C389 B.n349 VSUBS 0.008402f
C390 B.n350 VSUBS 0.008402f
C391 B.n351 VSUBS 0.008402f
C392 B.n352 VSUBS 0.008402f
C393 B.n353 VSUBS 0.008402f
C394 B.n354 VSUBS 0.008402f
C395 B.n355 VSUBS 0.008402f
C396 B.n356 VSUBS 0.008402f
C397 B.n357 VSUBS 0.008402f
C398 B.n358 VSUBS 0.008402f
C399 B.n359 VSUBS 0.008402f
C400 B.n360 VSUBS 0.008402f
C401 B.n361 VSUBS 0.008402f
C402 B.n362 VSUBS 0.008402f
C403 B.n363 VSUBS 0.008402f
C404 B.n364 VSUBS 0.008402f
C405 B.n365 VSUBS 0.008402f
C406 B.n366 VSUBS 0.008402f
C407 B.n367 VSUBS 0.008402f
C408 B.n368 VSUBS 0.008402f
C409 B.n369 VSUBS 0.008402f
C410 B.n370 VSUBS 0.008402f
C411 B.n371 VSUBS 0.008402f
C412 B.n372 VSUBS 0.008402f
C413 B.n373 VSUBS 0.008402f
C414 B.n374 VSUBS 0.008402f
C415 B.n375 VSUBS 0.008402f
C416 B.n376 VSUBS 0.008402f
C417 B.n377 VSUBS 0.008402f
C418 B.n378 VSUBS 0.008402f
C419 B.n379 VSUBS 0.008402f
C420 B.n380 VSUBS 0.008402f
C421 B.n381 VSUBS 0.008402f
C422 B.n382 VSUBS 0.008402f
C423 B.n383 VSUBS 0.008402f
C424 B.n384 VSUBS 0.008402f
C425 B.n385 VSUBS 0.008402f
C426 B.n386 VSUBS 0.008402f
C427 B.n387 VSUBS 0.008402f
C428 B.n388 VSUBS 0.008402f
C429 B.n389 VSUBS 0.008402f
C430 B.n390 VSUBS 0.008402f
C431 B.n391 VSUBS 0.008402f
C432 B.n392 VSUBS 0.008402f
C433 B.n393 VSUBS 0.008402f
C434 B.n394 VSUBS 0.008402f
C435 B.n395 VSUBS 0.008402f
C436 B.n396 VSUBS 0.008402f
C437 B.n397 VSUBS 0.008402f
C438 B.n398 VSUBS 0.008402f
C439 B.n399 VSUBS 0.008402f
C440 B.n400 VSUBS 0.008402f
C441 B.n401 VSUBS 0.008402f
C442 B.n402 VSUBS 0.008402f
C443 B.n403 VSUBS 0.008402f
C444 B.n404 VSUBS 0.008402f
C445 B.n405 VSUBS 0.008402f
C446 B.n406 VSUBS 0.008402f
C447 B.n407 VSUBS 0.008402f
C448 B.n408 VSUBS 0.008402f
C449 B.n409 VSUBS 0.008402f
C450 B.n410 VSUBS 0.008402f
C451 B.n411 VSUBS 0.008402f
C452 B.n412 VSUBS 0.008402f
C453 B.n413 VSUBS 0.008402f
C454 B.n414 VSUBS 0.008402f
C455 B.n415 VSUBS 0.008402f
C456 B.n416 VSUBS 0.008402f
C457 B.n417 VSUBS 0.008402f
C458 B.n418 VSUBS 0.008402f
C459 B.n419 VSUBS 0.008402f
C460 B.n420 VSUBS 0.005807f
C461 B.n421 VSUBS 0.019467f
C462 B.n422 VSUBS 0.006796f
C463 B.n423 VSUBS 0.008402f
C464 B.n424 VSUBS 0.008402f
C465 B.n425 VSUBS 0.008402f
C466 B.n426 VSUBS 0.008402f
C467 B.n427 VSUBS 0.008402f
C468 B.n428 VSUBS 0.008402f
C469 B.n429 VSUBS 0.008402f
C470 B.n430 VSUBS 0.008402f
C471 B.n431 VSUBS 0.008402f
C472 B.n432 VSUBS 0.008402f
C473 B.n433 VSUBS 0.008402f
C474 B.n434 VSUBS 0.006796f
C475 B.n435 VSUBS 0.008402f
C476 B.n436 VSUBS 0.008402f
C477 B.n437 VSUBS 0.005807f
C478 B.n438 VSUBS 0.008402f
C479 B.n439 VSUBS 0.008402f
C480 B.n440 VSUBS 0.008402f
C481 B.n441 VSUBS 0.008402f
C482 B.n442 VSUBS 0.008402f
C483 B.n443 VSUBS 0.008402f
C484 B.n444 VSUBS 0.008402f
C485 B.n445 VSUBS 0.008402f
C486 B.n446 VSUBS 0.008402f
C487 B.n447 VSUBS 0.008402f
C488 B.n448 VSUBS 0.008402f
C489 B.n449 VSUBS 0.008402f
C490 B.n450 VSUBS 0.008402f
C491 B.n451 VSUBS 0.008402f
C492 B.n452 VSUBS 0.008402f
C493 B.n453 VSUBS 0.008402f
C494 B.n454 VSUBS 0.008402f
C495 B.n455 VSUBS 0.008402f
C496 B.n456 VSUBS 0.008402f
C497 B.n457 VSUBS 0.008402f
C498 B.n458 VSUBS 0.008402f
C499 B.n459 VSUBS 0.008402f
C500 B.n460 VSUBS 0.008402f
C501 B.n461 VSUBS 0.008402f
C502 B.n462 VSUBS 0.008402f
C503 B.n463 VSUBS 0.008402f
C504 B.n464 VSUBS 0.008402f
C505 B.n465 VSUBS 0.008402f
C506 B.n466 VSUBS 0.008402f
C507 B.n467 VSUBS 0.008402f
C508 B.n468 VSUBS 0.008402f
C509 B.n469 VSUBS 0.008402f
C510 B.n470 VSUBS 0.008402f
C511 B.n471 VSUBS 0.008402f
C512 B.n472 VSUBS 0.008402f
C513 B.n473 VSUBS 0.008402f
C514 B.n474 VSUBS 0.008402f
C515 B.n475 VSUBS 0.008402f
C516 B.n476 VSUBS 0.008402f
C517 B.n477 VSUBS 0.008402f
C518 B.n478 VSUBS 0.008402f
C519 B.n479 VSUBS 0.008402f
C520 B.n480 VSUBS 0.008402f
C521 B.n481 VSUBS 0.008402f
C522 B.n482 VSUBS 0.008402f
C523 B.n483 VSUBS 0.008402f
C524 B.n484 VSUBS 0.008402f
C525 B.n485 VSUBS 0.008402f
C526 B.n486 VSUBS 0.008402f
C527 B.n487 VSUBS 0.008402f
C528 B.n488 VSUBS 0.008402f
C529 B.n489 VSUBS 0.008402f
C530 B.n490 VSUBS 0.008402f
C531 B.n491 VSUBS 0.008402f
C532 B.n492 VSUBS 0.008402f
C533 B.n493 VSUBS 0.008402f
C534 B.n494 VSUBS 0.008402f
C535 B.n495 VSUBS 0.008402f
C536 B.n496 VSUBS 0.008402f
C537 B.n497 VSUBS 0.008402f
C538 B.n498 VSUBS 0.008402f
C539 B.n499 VSUBS 0.008402f
C540 B.n500 VSUBS 0.008402f
C541 B.n501 VSUBS 0.008402f
C542 B.n502 VSUBS 0.008402f
C543 B.n503 VSUBS 0.008402f
C544 B.n504 VSUBS 0.008402f
C545 B.n505 VSUBS 0.008402f
C546 B.n506 VSUBS 0.008402f
C547 B.n507 VSUBS 0.008402f
C548 B.n508 VSUBS 0.008402f
C549 B.n509 VSUBS 0.008402f
C550 B.n510 VSUBS 0.008402f
C551 B.n511 VSUBS 0.008402f
C552 B.n512 VSUBS 0.008402f
C553 B.n513 VSUBS 0.008402f
C554 B.n514 VSUBS 0.020386f
C555 B.n515 VSUBS 0.020386f
C556 B.n516 VSUBS 0.019896f
C557 B.n517 VSUBS 0.008402f
C558 B.n518 VSUBS 0.008402f
C559 B.n519 VSUBS 0.008402f
C560 B.n520 VSUBS 0.008402f
C561 B.n521 VSUBS 0.008402f
C562 B.n522 VSUBS 0.008402f
C563 B.n523 VSUBS 0.008402f
C564 B.n524 VSUBS 0.008402f
C565 B.n525 VSUBS 0.008402f
C566 B.n526 VSUBS 0.008402f
C567 B.n527 VSUBS 0.008402f
C568 B.n528 VSUBS 0.008402f
C569 B.n529 VSUBS 0.008402f
C570 B.n530 VSUBS 0.008402f
C571 B.n531 VSUBS 0.008402f
C572 B.n532 VSUBS 0.008402f
C573 B.n533 VSUBS 0.008402f
C574 B.n534 VSUBS 0.008402f
C575 B.n535 VSUBS 0.008402f
C576 B.n536 VSUBS 0.008402f
C577 B.n537 VSUBS 0.008402f
C578 B.n538 VSUBS 0.008402f
C579 B.n539 VSUBS 0.008402f
C580 B.n540 VSUBS 0.008402f
C581 B.n541 VSUBS 0.008402f
C582 B.n542 VSUBS 0.008402f
C583 B.n543 VSUBS 0.008402f
C584 B.n544 VSUBS 0.008402f
C585 B.n545 VSUBS 0.008402f
C586 B.n546 VSUBS 0.008402f
C587 B.n547 VSUBS 0.008402f
C588 B.n548 VSUBS 0.008402f
C589 B.n549 VSUBS 0.008402f
C590 B.n550 VSUBS 0.008402f
C591 B.n551 VSUBS 0.008402f
C592 B.n552 VSUBS 0.008402f
C593 B.n553 VSUBS 0.008402f
C594 B.n554 VSUBS 0.008402f
C595 B.n555 VSUBS 0.008402f
C596 B.n556 VSUBS 0.008402f
C597 B.n557 VSUBS 0.008402f
C598 B.n558 VSUBS 0.008402f
C599 B.n559 VSUBS 0.008402f
C600 B.n560 VSUBS 0.008402f
C601 B.n561 VSUBS 0.008402f
C602 B.n562 VSUBS 0.008402f
C603 B.n563 VSUBS 0.008402f
C604 B.n564 VSUBS 0.008402f
C605 B.n565 VSUBS 0.008402f
C606 B.n566 VSUBS 0.008402f
C607 B.n567 VSUBS 0.008402f
C608 B.n568 VSUBS 0.008402f
C609 B.n569 VSUBS 0.008402f
C610 B.n570 VSUBS 0.008402f
C611 B.n571 VSUBS 0.008402f
C612 B.n572 VSUBS 0.008402f
C613 B.n573 VSUBS 0.008402f
C614 B.n574 VSUBS 0.008402f
C615 B.n575 VSUBS 0.008402f
C616 B.n576 VSUBS 0.008402f
C617 B.n577 VSUBS 0.008402f
C618 B.n578 VSUBS 0.008402f
C619 B.n579 VSUBS 0.008402f
C620 B.n580 VSUBS 0.008402f
C621 B.n581 VSUBS 0.008402f
C622 B.n582 VSUBS 0.008402f
C623 B.n583 VSUBS 0.008402f
C624 B.n584 VSUBS 0.008402f
C625 B.n585 VSUBS 0.008402f
C626 B.n586 VSUBS 0.008402f
C627 B.n587 VSUBS 0.008402f
C628 B.n588 VSUBS 0.008402f
C629 B.n589 VSUBS 0.008402f
C630 B.n590 VSUBS 0.008402f
C631 B.n591 VSUBS 0.008402f
C632 B.n592 VSUBS 0.008402f
C633 B.n593 VSUBS 0.008402f
C634 B.n594 VSUBS 0.008402f
C635 B.n595 VSUBS 0.008402f
C636 B.n596 VSUBS 0.008402f
C637 B.n597 VSUBS 0.008402f
C638 B.n598 VSUBS 0.008402f
C639 B.n599 VSUBS 0.008402f
C640 B.n600 VSUBS 0.008402f
C641 B.n601 VSUBS 0.008402f
C642 B.n602 VSUBS 0.008402f
C643 B.n603 VSUBS 0.008402f
C644 B.n604 VSUBS 0.008402f
C645 B.n605 VSUBS 0.008402f
C646 B.n606 VSUBS 0.008402f
C647 B.n607 VSUBS 0.008402f
C648 B.n608 VSUBS 0.008402f
C649 B.n609 VSUBS 0.008402f
C650 B.n610 VSUBS 0.008402f
C651 B.n611 VSUBS 0.008402f
C652 B.n612 VSUBS 0.008402f
C653 B.n613 VSUBS 0.008402f
C654 B.n614 VSUBS 0.008402f
C655 B.n615 VSUBS 0.008402f
C656 B.n616 VSUBS 0.008402f
C657 B.n617 VSUBS 0.008402f
C658 B.n618 VSUBS 0.008402f
C659 B.n619 VSUBS 0.008402f
C660 B.n620 VSUBS 0.008402f
C661 B.n621 VSUBS 0.008402f
C662 B.n622 VSUBS 0.008402f
C663 B.n623 VSUBS 0.008402f
C664 B.n624 VSUBS 0.008402f
C665 B.n625 VSUBS 0.008402f
C666 B.n626 VSUBS 0.008402f
C667 B.n627 VSUBS 0.008402f
C668 B.n628 VSUBS 0.008402f
C669 B.n629 VSUBS 0.008402f
C670 B.n630 VSUBS 0.008402f
C671 B.n631 VSUBS 0.008402f
C672 B.n632 VSUBS 0.008402f
C673 B.n633 VSUBS 0.008402f
C674 B.n634 VSUBS 0.008402f
C675 B.n635 VSUBS 0.008402f
C676 B.n636 VSUBS 0.008402f
C677 B.n637 VSUBS 0.008402f
C678 B.n638 VSUBS 0.008402f
C679 B.n639 VSUBS 0.008402f
C680 B.n640 VSUBS 0.008402f
C681 B.n641 VSUBS 0.008402f
C682 B.n642 VSUBS 0.008402f
C683 B.n643 VSUBS 0.008402f
C684 B.n644 VSUBS 0.008402f
C685 B.n645 VSUBS 0.008402f
C686 B.n646 VSUBS 0.008402f
C687 B.n647 VSUBS 0.008402f
C688 B.n648 VSUBS 0.008402f
C689 B.n649 VSUBS 0.008402f
C690 B.n650 VSUBS 0.008402f
C691 B.n651 VSUBS 0.008402f
C692 B.n652 VSUBS 0.008402f
C693 B.n653 VSUBS 0.008402f
C694 B.n654 VSUBS 0.008402f
C695 B.n655 VSUBS 0.008402f
C696 B.n656 VSUBS 0.008402f
C697 B.n657 VSUBS 0.008402f
C698 B.n658 VSUBS 0.008402f
C699 B.n659 VSUBS 0.008402f
C700 B.n660 VSUBS 0.008402f
C701 B.n661 VSUBS 0.008402f
C702 B.n662 VSUBS 0.008402f
C703 B.n663 VSUBS 0.008402f
C704 B.n664 VSUBS 0.008402f
C705 B.n665 VSUBS 0.008402f
C706 B.n666 VSUBS 0.008402f
C707 B.n667 VSUBS 0.008402f
C708 B.n668 VSUBS 0.008402f
C709 B.n669 VSUBS 0.008402f
C710 B.n670 VSUBS 0.008402f
C711 B.n671 VSUBS 0.008402f
C712 B.n672 VSUBS 0.008402f
C713 B.n673 VSUBS 0.008402f
C714 B.n674 VSUBS 0.008402f
C715 B.n675 VSUBS 0.008402f
C716 B.n676 VSUBS 0.008402f
C717 B.n677 VSUBS 0.008402f
C718 B.n678 VSUBS 0.008402f
C719 B.n679 VSUBS 0.008402f
C720 B.n680 VSUBS 0.008402f
C721 B.n681 VSUBS 0.008402f
C722 B.n682 VSUBS 0.008402f
C723 B.n683 VSUBS 0.008402f
C724 B.n684 VSUBS 0.008402f
C725 B.n685 VSUBS 0.008402f
C726 B.n686 VSUBS 0.008402f
C727 B.n687 VSUBS 0.008402f
C728 B.n688 VSUBS 0.008402f
C729 B.n689 VSUBS 0.008402f
C730 B.n690 VSUBS 0.008402f
C731 B.n691 VSUBS 0.008402f
C732 B.n692 VSUBS 0.008402f
C733 B.n693 VSUBS 0.008402f
C734 B.n694 VSUBS 0.008402f
C735 B.n695 VSUBS 0.008402f
C736 B.n696 VSUBS 0.008402f
C737 B.n697 VSUBS 0.008402f
C738 B.n698 VSUBS 0.008402f
C739 B.n699 VSUBS 0.008402f
C740 B.n700 VSUBS 0.008402f
C741 B.n701 VSUBS 0.008402f
C742 B.n702 VSUBS 0.020853f
C743 B.n703 VSUBS 0.019429f
C744 B.n704 VSUBS 0.020386f
C745 B.n705 VSUBS 0.008402f
C746 B.n706 VSUBS 0.008402f
C747 B.n707 VSUBS 0.008402f
C748 B.n708 VSUBS 0.008402f
C749 B.n709 VSUBS 0.008402f
C750 B.n710 VSUBS 0.008402f
C751 B.n711 VSUBS 0.008402f
C752 B.n712 VSUBS 0.008402f
C753 B.n713 VSUBS 0.008402f
C754 B.n714 VSUBS 0.008402f
C755 B.n715 VSUBS 0.008402f
C756 B.n716 VSUBS 0.008402f
C757 B.n717 VSUBS 0.008402f
C758 B.n718 VSUBS 0.008402f
C759 B.n719 VSUBS 0.008402f
C760 B.n720 VSUBS 0.008402f
C761 B.n721 VSUBS 0.008402f
C762 B.n722 VSUBS 0.008402f
C763 B.n723 VSUBS 0.008402f
C764 B.n724 VSUBS 0.008402f
C765 B.n725 VSUBS 0.008402f
C766 B.n726 VSUBS 0.008402f
C767 B.n727 VSUBS 0.008402f
C768 B.n728 VSUBS 0.008402f
C769 B.n729 VSUBS 0.008402f
C770 B.n730 VSUBS 0.008402f
C771 B.n731 VSUBS 0.008402f
C772 B.n732 VSUBS 0.008402f
C773 B.n733 VSUBS 0.008402f
C774 B.n734 VSUBS 0.008402f
C775 B.n735 VSUBS 0.008402f
C776 B.n736 VSUBS 0.008402f
C777 B.n737 VSUBS 0.008402f
C778 B.n738 VSUBS 0.008402f
C779 B.n739 VSUBS 0.008402f
C780 B.n740 VSUBS 0.008402f
C781 B.n741 VSUBS 0.008402f
C782 B.n742 VSUBS 0.008402f
C783 B.n743 VSUBS 0.008402f
C784 B.n744 VSUBS 0.008402f
C785 B.n745 VSUBS 0.008402f
C786 B.n746 VSUBS 0.008402f
C787 B.n747 VSUBS 0.008402f
C788 B.n748 VSUBS 0.008402f
C789 B.n749 VSUBS 0.008402f
C790 B.n750 VSUBS 0.008402f
C791 B.n751 VSUBS 0.008402f
C792 B.n752 VSUBS 0.008402f
C793 B.n753 VSUBS 0.008402f
C794 B.n754 VSUBS 0.008402f
C795 B.n755 VSUBS 0.008402f
C796 B.n756 VSUBS 0.008402f
C797 B.n757 VSUBS 0.008402f
C798 B.n758 VSUBS 0.008402f
C799 B.n759 VSUBS 0.008402f
C800 B.n760 VSUBS 0.008402f
C801 B.n761 VSUBS 0.008402f
C802 B.n762 VSUBS 0.008402f
C803 B.n763 VSUBS 0.008402f
C804 B.n764 VSUBS 0.008402f
C805 B.n765 VSUBS 0.008402f
C806 B.n766 VSUBS 0.008402f
C807 B.n767 VSUBS 0.008402f
C808 B.n768 VSUBS 0.008402f
C809 B.n769 VSUBS 0.008402f
C810 B.n770 VSUBS 0.008402f
C811 B.n771 VSUBS 0.008402f
C812 B.n772 VSUBS 0.008402f
C813 B.n773 VSUBS 0.008402f
C814 B.n774 VSUBS 0.008402f
C815 B.n775 VSUBS 0.008402f
C816 B.n776 VSUBS 0.008402f
C817 B.n777 VSUBS 0.008402f
C818 B.n778 VSUBS 0.008402f
C819 B.n779 VSUBS 0.008402f
C820 B.n780 VSUBS 0.008402f
C821 B.n781 VSUBS 0.005807f
C822 B.n782 VSUBS 0.008402f
C823 B.n783 VSUBS 0.008402f
C824 B.n784 VSUBS 0.006796f
C825 B.n785 VSUBS 0.008402f
C826 B.n786 VSUBS 0.008402f
C827 B.n787 VSUBS 0.008402f
C828 B.n788 VSUBS 0.008402f
C829 B.n789 VSUBS 0.008402f
C830 B.n790 VSUBS 0.008402f
C831 B.n791 VSUBS 0.008402f
C832 B.n792 VSUBS 0.008402f
C833 B.n793 VSUBS 0.008402f
C834 B.n794 VSUBS 0.008402f
C835 B.n795 VSUBS 0.008402f
C836 B.n796 VSUBS 0.006796f
C837 B.n797 VSUBS 0.019467f
C838 B.n798 VSUBS 0.005807f
C839 B.n799 VSUBS 0.008402f
C840 B.n800 VSUBS 0.008402f
C841 B.n801 VSUBS 0.008402f
C842 B.n802 VSUBS 0.008402f
C843 B.n803 VSUBS 0.008402f
C844 B.n804 VSUBS 0.008402f
C845 B.n805 VSUBS 0.008402f
C846 B.n806 VSUBS 0.008402f
C847 B.n807 VSUBS 0.008402f
C848 B.n808 VSUBS 0.008402f
C849 B.n809 VSUBS 0.008402f
C850 B.n810 VSUBS 0.008402f
C851 B.n811 VSUBS 0.008402f
C852 B.n812 VSUBS 0.008402f
C853 B.n813 VSUBS 0.008402f
C854 B.n814 VSUBS 0.008402f
C855 B.n815 VSUBS 0.008402f
C856 B.n816 VSUBS 0.008402f
C857 B.n817 VSUBS 0.008402f
C858 B.n818 VSUBS 0.008402f
C859 B.n819 VSUBS 0.008402f
C860 B.n820 VSUBS 0.008402f
C861 B.n821 VSUBS 0.008402f
C862 B.n822 VSUBS 0.008402f
C863 B.n823 VSUBS 0.008402f
C864 B.n824 VSUBS 0.008402f
C865 B.n825 VSUBS 0.008402f
C866 B.n826 VSUBS 0.008402f
C867 B.n827 VSUBS 0.008402f
C868 B.n828 VSUBS 0.008402f
C869 B.n829 VSUBS 0.008402f
C870 B.n830 VSUBS 0.008402f
C871 B.n831 VSUBS 0.008402f
C872 B.n832 VSUBS 0.008402f
C873 B.n833 VSUBS 0.008402f
C874 B.n834 VSUBS 0.008402f
C875 B.n835 VSUBS 0.008402f
C876 B.n836 VSUBS 0.008402f
C877 B.n837 VSUBS 0.008402f
C878 B.n838 VSUBS 0.008402f
C879 B.n839 VSUBS 0.008402f
C880 B.n840 VSUBS 0.008402f
C881 B.n841 VSUBS 0.008402f
C882 B.n842 VSUBS 0.008402f
C883 B.n843 VSUBS 0.008402f
C884 B.n844 VSUBS 0.008402f
C885 B.n845 VSUBS 0.008402f
C886 B.n846 VSUBS 0.008402f
C887 B.n847 VSUBS 0.008402f
C888 B.n848 VSUBS 0.008402f
C889 B.n849 VSUBS 0.008402f
C890 B.n850 VSUBS 0.008402f
C891 B.n851 VSUBS 0.008402f
C892 B.n852 VSUBS 0.008402f
C893 B.n853 VSUBS 0.008402f
C894 B.n854 VSUBS 0.008402f
C895 B.n855 VSUBS 0.008402f
C896 B.n856 VSUBS 0.008402f
C897 B.n857 VSUBS 0.008402f
C898 B.n858 VSUBS 0.008402f
C899 B.n859 VSUBS 0.008402f
C900 B.n860 VSUBS 0.008402f
C901 B.n861 VSUBS 0.008402f
C902 B.n862 VSUBS 0.008402f
C903 B.n863 VSUBS 0.008402f
C904 B.n864 VSUBS 0.008402f
C905 B.n865 VSUBS 0.008402f
C906 B.n866 VSUBS 0.008402f
C907 B.n867 VSUBS 0.008402f
C908 B.n868 VSUBS 0.008402f
C909 B.n869 VSUBS 0.008402f
C910 B.n870 VSUBS 0.008402f
C911 B.n871 VSUBS 0.008402f
C912 B.n872 VSUBS 0.008402f
C913 B.n873 VSUBS 0.008402f
C914 B.n874 VSUBS 0.008402f
C915 B.n875 VSUBS 0.008402f
C916 B.n876 VSUBS 0.020386f
C917 B.n877 VSUBS 0.019896f
C918 B.n878 VSUBS 0.019896f
C919 B.n879 VSUBS 0.008402f
C920 B.n880 VSUBS 0.008402f
C921 B.n881 VSUBS 0.008402f
C922 B.n882 VSUBS 0.008402f
C923 B.n883 VSUBS 0.008402f
C924 B.n884 VSUBS 0.008402f
C925 B.n885 VSUBS 0.008402f
C926 B.n886 VSUBS 0.008402f
C927 B.n887 VSUBS 0.008402f
C928 B.n888 VSUBS 0.008402f
C929 B.n889 VSUBS 0.008402f
C930 B.n890 VSUBS 0.008402f
C931 B.n891 VSUBS 0.008402f
C932 B.n892 VSUBS 0.008402f
C933 B.n893 VSUBS 0.008402f
C934 B.n894 VSUBS 0.008402f
C935 B.n895 VSUBS 0.008402f
C936 B.n896 VSUBS 0.008402f
C937 B.n897 VSUBS 0.008402f
C938 B.n898 VSUBS 0.008402f
C939 B.n899 VSUBS 0.008402f
C940 B.n900 VSUBS 0.008402f
C941 B.n901 VSUBS 0.008402f
C942 B.n902 VSUBS 0.008402f
C943 B.n903 VSUBS 0.008402f
C944 B.n904 VSUBS 0.008402f
C945 B.n905 VSUBS 0.008402f
C946 B.n906 VSUBS 0.008402f
C947 B.n907 VSUBS 0.008402f
C948 B.n908 VSUBS 0.008402f
C949 B.n909 VSUBS 0.008402f
C950 B.n910 VSUBS 0.008402f
C951 B.n911 VSUBS 0.008402f
C952 B.n912 VSUBS 0.008402f
C953 B.n913 VSUBS 0.008402f
C954 B.n914 VSUBS 0.008402f
C955 B.n915 VSUBS 0.008402f
C956 B.n916 VSUBS 0.008402f
C957 B.n917 VSUBS 0.008402f
C958 B.n918 VSUBS 0.008402f
C959 B.n919 VSUBS 0.008402f
C960 B.n920 VSUBS 0.008402f
C961 B.n921 VSUBS 0.008402f
C962 B.n922 VSUBS 0.008402f
C963 B.n923 VSUBS 0.008402f
C964 B.n924 VSUBS 0.008402f
C965 B.n925 VSUBS 0.008402f
C966 B.n926 VSUBS 0.008402f
C967 B.n927 VSUBS 0.008402f
C968 B.n928 VSUBS 0.008402f
C969 B.n929 VSUBS 0.008402f
C970 B.n930 VSUBS 0.008402f
C971 B.n931 VSUBS 0.008402f
C972 B.n932 VSUBS 0.008402f
C973 B.n933 VSUBS 0.008402f
C974 B.n934 VSUBS 0.008402f
C975 B.n935 VSUBS 0.008402f
C976 B.n936 VSUBS 0.008402f
C977 B.n937 VSUBS 0.008402f
C978 B.n938 VSUBS 0.008402f
C979 B.n939 VSUBS 0.008402f
C980 B.n940 VSUBS 0.008402f
C981 B.n941 VSUBS 0.008402f
C982 B.n942 VSUBS 0.008402f
C983 B.n943 VSUBS 0.008402f
C984 B.n944 VSUBS 0.008402f
C985 B.n945 VSUBS 0.008402f
C986 B.n946 VSUBS 0.008402f
C987 B.n947 VSUBS 0.008402f
C988 B.n948 VSUBS 0.008402f
C989 B.n949 VSUBS 0.008402f
C990 B.n950 VSUBS 0.008402f
C991 B.n951 VSUBS 0.008402f
C992 B.n952 VSUBS 0.008402f
C993 B.n953 VSUBS 0.008402f
C994 B.n954 VSUBS 0.008402f
C995 B.n955 VSUBS 0.008402f
C996 B.n956 VSUBS 0.008402f
C997 B.n957 VSUBS 0.008402f
C998 B.n958 VSUBS 0.008402f
C999 B.n959 VSUBS 0.008402f
C1000 B.n960 VSUBS 0.008402f
C1001 B.n961 VSUBS 0.008402f
C1002 B.n962 VSUBS 0.008402f
C1003 B.n963 VSUBS 0.008402f
C1004 B.n964 VSUBS 0.008402f
C1005 B.n965 VSUBS 0.008402f
C1006 B.n966 VSUBS 0.008402f
C1007 B.n967 VSUBS 0.008402f
C1008 B.n968 VSUBS 0.008402f
C1009 B.n969 VSUBS 0.008402f
C1010 B.n970 VSUBS 0.008402f
C1011 B.n971 VSUBS 0.019026f
C1012 VDD2.t7 VSUBS 3.8865f
C1013 VDD2.t5 VSUBS 0.36184f
C1014 VDD2.t1 VSUBS 0.36184f
C1015 VDD2.n0 VSUBS 2.9679f
C1016 VDD2.n1 VSUBS 1.72411f
C1017 VDD2.t0 VSUBS 0.36184f
C1018 VDD2.t8 VSUBS 0.36184f
C1019 VDD2.n2 VSUBS 2.9933f
C1020 VDD2.n3 VSUBS 4.01436f
C1021 VDD2.t9 VSUBS 3.85565f
C1022 VDD2.n4 VSUBS 4.33916f
C1023 VDD2.t6 VSUBS 0.36184f
C1024 VDD2.t2 VSUBS 0.36184f
C1025 VDD2.n5 VSUBS 2.96791f
C1026 VDD2.n6 VSUBS 0.860165f
C1027 VDD2.t4 VSUBS 0.36184f
C1028 VDD2.t3 VSUBS 0.36184f
C1029 VDD2.n7 VSUBS 2.99324f
C1030 VN.n0 VSUBS 0.033641f
C1031 VN.t1 VSUBS 3.01634f
C1032 VN.n1 VSUBS 0.047775f
C1033 VN.n2 VSUBS 0.025518f
C1034 VN.t9 VSUBS 3.01634f
C1035 VN.n3 VSUBS 1.05042f
C1036 VN.n4 VSUBS 0.025518f
C1037 VN.n5 VSUBS 0.020814f
C1038 VN.n6 VSUBS 0.025518f
C1039 VN.t8 VSUBS 3.01634f
C1040 VN.n7 VSUBS 0.047321f
C1041 VN.n8 VSUBS 0.025518f
C1042 VN.n9 VSUBS 0.047321f
C1043 VN.t2 VSUBS 3.24072f
C1044 VN.n10 VSUBS 1.0974f
C1045 VN.t4 VSUBS 3.01634f
C1046 VN.n11 VSUBS 1.11775f
C1047 VN.n12 VSUBS 0.026296f
C1048 VN.n13 VSUBS 0.249637f
C1049 VN.n14 VSUBS 0.025518f
C1050 VN.n15 VSUBS 0.025518f
C1051 VN.n16 VSUBS 0.049721f
C1052 VN.n17 VSUBS 0.020814f
C1053 VN.n18 VSUBS 0.050975f
C1054 VN.n19 VSUBS 0.025518f
C1055 VN.n20 VSUBS 0.025518f
C1056 VN.n21 VSUBS 0.025518f
C1057 VN.n22 VSUBS 1.07438f
C1058 VN.n23 VSUBS 0.047321f
C1059 VN.n24 VSUBS 0.050975f
C1060 VN.n25 VSUBS 0.025518f
C1061 VN.n26 VSUBS 0.025518f
C1062 VN.n27 VSUBS 0.025518f
C1063 VN.n28 VSUBS 0.049721f
C1064 VN.n29 VSUBS 0.047321f
C1065 VN.n30 VSUBS 0.026296f
C1066 VN.n31 VSUBS 0.025518f
C1067 VN.n32 VSUBS 0.025518f
C1068 VN.n33 VSUBS 0.044985f
C1069 VN.n34 VSUBS 0.051235f
C1070 VN.n35 VSUBS 0.022501f
C1071 VN.n36 VSUBS 0.025518f
C1072 VN.n37 VSUBS 0.025518f
C1073 VN.n38 VSUBS 0.025518f
C1074 VN.n39 VSUBS 0.047321f
C1075 VN.n40 VSUBS 0.028632f
C1076 VN.n41 VSUBS 1.13246f
C1077 VN.n42 VSUBS 0.045664f
C1078 VN.n43 VSUBS 0.033641f
C1079 VN.t0 VSUBS 3.01634f
C1080 VN.n44 VSUBS 0.047775f
C1081 VN.n45 VSUBS 0.025518f
C1082 VN.t3 VSUBS 3.01634f
C1083 VN.n46 VSUBS 1.05042f
C1084 VN.n47 VSUBS 0.025518f
C1085 VN.n48 VSUBS 0.020814f
C1086 VN.n49 VSUBS 0.025518f
C1087 VN.t7 VSUBS 3.01634f
C1088 VN.n50 VSUBS 0.047321f
C1089 VN.n51 VSUBS 0.025518f
C1090 VN.n52 VSUBS 0.047321f
C1091 VN.t6 VSUBS 3.24072f
C1092 VN.n53 VSUBS 1.0974f
C1093 VN.t5 VSUBS 3.01634f
C1094 VN.n54 VSUBS 1.11775f
C1095 VN.n55 VSUBS 0.026296f
C1096 VN.n56 VSUBS 0.249637f
C1097 VN.n57 VSUBS 0.025518f
C1098 VN.n58 VSUBS 0.025518f
C1099 VN.n59 VSUBS 0.049721f
C1100 VN.n60 VSUBS 0.020814f
C1101 VN.n61 VSUBS 0.050975f
C1102 VN.n62 VSUBS 0.025518f
C1103 VN.n63 VSUBS 0.025518f
C1104 VN.n64 VSUBS 0.025518f
C1105 VN.n65 VSUBS 1.07438f
C1106 VN.n66 VSUBS 0.047321f
C1107 VN.n67 VSUBS 0.050975f
C1108 VN.n68 VSUBS 0.025518f
C1109 VN.n69 VSUBS 0.025518f
C1110 VN.n70 VSUBS 0.025518f
C1111 VN.n71 VSUBS 0.049721f
C1112 VN.n72 VSUBS 0.047321f
C1113 VN.n73 VSUBS 0.026296f
C1114 VN.n74 VSUBS 0.025518f
C1115 VN.n75 VSUBS 0.025518f
C1116 VN.n76 VSUBS 0.044985f
C1117 VN.n77 VSUBS 0.051235f
C1118 VN.n78 VSUBS 0.022501f
C1119 VN.n79 VSUBS 0.025518f
C1120 VN.n80 VSUBS 0.025518f
C1121 VN.n81 VSUBS 0.025518f
C1122 VN.n82 VSUBS 0.047321f
C1123 VN.n83 VSUBS 0.028632f
C1124 VN.n84 VSUBS 1.13246f
C1125 VN.n85 VSUBS 1.71445f
C1126 VDD1.t5 VSUBS 3.89693f
C1127 VDD1.t7 VSUBS 0.362809f
C1128 VDD1.t4 VSUBS 0.362809f
C1129 VDD1.n0 VSUBS 2.97585f
C1130 VDD1.n1 VSUBS 1.73819f
C1131 VDD1.t9 VSUBS 3.89691f
C1132 VDD1.t1 VSUBS 0.362809f
C1133 VDD1.t2 VSUBS 0.362809f
C1134 VDD1.n2 VSUBS 2.97585f
C1135 VDD1.n3 VSUBS 1.72873f
C1136 VDD1.t3 VSUBS 0.362809f
C1137 VDD1.t6 VSUBS 0.362809f
C1138 VDD1.n4 VSUBS 3.00131f
C1139 VDD1.n5 VSUBS 4.17671f
C1140 VDD1.t8 VSUBS 0.362809f
C1141 VDD1.t0 VSUBS 0.362809f
C1142 VDD1.n6 VSUBS 2.97584f
C1143 VDD1.n7 VSUBS 4.38563f
C1144 VTAIL.t3 VSUBS 0.349578f
C1145 VTAIL.t1 VSUBS 0.349578f
C1146 VTAIL.n0 VSUBS 2.71013f
C1147 VTAIL.n1 VSUBS 0.992537f
C1148 VTAIL.t13 VSUBS 3.5457f
C1149 VTAIL.n2 VSUBS 1.16428f
C1150 VTAIL.t19 VSUBS 0.349578f
C1151 VTAIL.t16 VSUBS 0.349578f
C1152 VTAIL.n3 VSUBS 2.71013f
C1153 VTAIL.n4 VSUBS 1.12248f
C1154 VTAIL.t12 VSUBS 0.349578f
C1155 VTAIL.t10 VSUBS 0.349578f
C1156 VTAIL.n5 VSUBS 2.71013f
C1157 VTAIL.n6 VSUBS 2.96727f
C1158 VTAIL.t5 VSUBS 0.349578f
C1159 VTAIL.t2 VSUBS 0.349578f
C1160 VTAIL.n7 VSUBS 2.71014f
C1161 VTAIL.n8 VSUBS 2.96727f
C1162 VTAIL.t7 VSUBS 0.349578f
C1163 VTAIL.t6 VSUBS 0.349578f
C1164 VTAIL.n9 VSUBS 2.71014f
C1165 VTAIL.n10 VSUBS 1.12247f
C1166 VTAIL.t4 VSUBS 3.54573f
C1167 VTAIL.n11 VSUBS 1.16425f
C1168 VTAIL.t18 VSUBS 0.349578f
C1169 VTAIL.t17 VSUBS 0.349578f
C1170 VTAIL.n12 VSUBS 2.71014f
C1171 VTAIL.n13 VSUBS 1.04645f
C1172 VTAIL.t11 VSUBS 0.349578f
C1173 VTAIL.t14 VSUBS 0.349578f
C1174 VTAIL.n14 VSUBS 2.71014f
C1175 VTAIL.n15 VSUBS 1.12247f
C1176 VTAIL.t15 VSUBS 3.5457f
C1177 VTAIL.n16 VSUBS 2.84848f
C1178 VTAIL.t9 VSUBS 3.5457f
C1179 VTAIL.n17 VSUBS 2.84848f
C1180 VTAIL.t8 VSUBS 0.349578f
C1181 VTAIL.t0 VSUBS 0.349578f
C1182 VTAIL.n18 VSUBS 2.71013f
C1183 VTAIL.n19 VSUBS 0.939785f
C1184 VP.n0 VSUBS 0.036127f
C1185 VP.t3 VSUBS 3.23917f
C1186 VP.n1 VSUBS 0.051305f
C1187 VP.n2 VSUBS 0.027403f
C1188 VP.t6 VSUBS 3.23917f
C1189 VP.n3 VSUBS 1.12802f
C1190 VP.n4 VSUBS 0.027403f
C1191 VP.n5 VSUBS 0.022352f
C1192 VP.n6 VSUBS 0.027403f
C1193 VP.t7 VSUBS 3.23917f
C1194 VP.n7 VSUBS 0.050817f
C1195 VP.n8 VSUBS 0.027403f
C1196 VP.n9 VSUBS 0.050817f
C1197 VP.n10 VSUBS 0.027403f
C1198 VP.t8 VSUBS 3.23917f
C1199 VP.n11 VSUBS 0.024163f
C1200 VP.n12 VSUBS 0.027403f
C1201 VP.t0 VSUBS 3.23917f
C1202 VP.n13 VSUBS 1.21612f
C1203 VP.n14 VSUBS 0.036127f
C1204 VP.t9 VSUBS 3.23917f
C1205 VP.n15 VSUBS 0.051305f
C1206 VP.n16 VSUBS 0.027403f
C1207 VP.t1 VSUBS 3.23917f
C1208 VP.n17 VSUBS 1.12802f
C1209 VP.n18 VSUBS 0.027403f
C1210 VP.n19 VSUBS 0.022352f
C1211 VP.n20 VSUBS 0.027403f
C1212 VP.t5 VSUBS 3.23917f
C1213 VP.n21 VSUBS 0.050817f
C1214 VP.n22 VSUBS 0.027403f
C1215 VP.n23 VSUBS 0.050817f
C1216 VP.t4 VSUBS 3.48012f
C1217 VP.n24 VSUBS 1.17846f
C1218 VP.t2 VSUBS 3.23917f
C1219 VP.n25 VSUBS 1.20032f
C1220 VP.n26 VSUBS 0.028239f
C1221 VP.n27 VSUBS 0.268079f
C1222 VP.n28 VSUBS 0.027403f
C1223 VP.n29 VSUBS 0.027403f
C1224 VP.n30 VSUBS 0.053395f
C1225 VP.n31 VSUBS 0.022352f
C1226 VP.n32 VSUBS 0.054741f
C1227 VP.n33 VSUBS 0.027403f
C1228 VP.n34 VSUBS 0.027403f
C1229 VP.n35 VSUBS 0.027403f
C1230 VP.n36 VSUBS 1.15375f
C1231 VP.n37 VSUBS 0.050817f
C1232 VP.n38 VSUBS 0.054741f
C1233 VP.n39 VSUBS 0.027403f
C1234 VP.n40 VSUBS 0.027403f
C1235 VP.n41 VSUBS 0.027403f
C1236 VP.n42 VSUBS 0.053395f
C1237 VP.n43 VSUBS 0.050817f
C1238 VP.n44 VSUBS 0.028239f
C1239 VP.n45 VSUBS 0.027403f
C1240 VP.n46 VSUBS 0.027403f
C1241 VP.n47 VSUBS 0.048308f
C1242 VP.n48 VSUBS 0.05502f
C1243 VP.n49 VSUBS 0.024163f
C1244 VP.n50 VSUBS 0.027403f
C1245 VP.n51 VSUBS 0.027403f
C1246 VP.n52 VSUBS 0.027403f
C1247 VP.n53 VSUBS 0.050817f
C1248 VP.n54 VSUBS 0.030747f
C1249 VP.n55 VSUBS 1.21612f
C1250 VP.n56 VSUBS 1.82665f
C1251 VP.n57 VSUBS 1.84409f
C1252 VP.n58 VSUBS 0.036127f
C1253 VP.n59 VSUBS 0.030747f
C1254 VP.n60 VSUBS 0.050817f
C1255 VP.n61 VSUBS 0.051305f
C1256 VP.n62 VSUBS 0.027403f
C1257 VP.n63 VSUBS 0.027403f
C1258 VP.n64 VSUBS 0.027403f
C1259 VP.n65 VSUBS 0.05502f
C1260 VP.n66 VSUBS 0.048308f
C1261 VP.n67 VSUBS 1.12802f
C1262 VP.n68 VSUBS 0.028239f
C1263 VP.n69 VSUBS 0.027403f
C1264 VP.n70 VSUBS 0.027403f
C1265 VP.n71 VSUBS 0.027403f
C1266 VP.n72 VSUBS 0.053395f
C1267 VP.n73 VSUBS 0.022352f
C1268 VP.n74 VSUBS 0.054741f
C1269 VP.n75 VSUBS 0.027403f
C1270 VP.n76 VSUBS 0.027403f
C1271 VP.n77 VSUBS 0.027403f
C1272 VP.n78 VSUBS 1.15375f
C1273 VP.n79 VSUBS 0.050817f
C1274 VP.n80 VSUBS 0.054741f
C1275 VP.n81 VSUBS 0.027403f
C1276 VP.n82 VSUBS 0.027403f
C1277 VP.n83 VSUBS 0.027403f
C1278 VP.n84 VSUBS 0.053395f
C1279 VP.n85 VSUBS 0.050817f
C1280 VP.n86 VSUBS 0.028239f
C1281 VP.n87 VSUBS 0.027403f
C1282 VP.n88 VSUBS 0.027403f
C1283 VP.n89 VSUBS 0.048308f
C1284 VP.n90 VSUBS 0.05502f
C1285 VP.n91 VSUBS 0.024163f
C1286 VP.n92 VSUBS 0.027403f
C1287 VP.n93 VSUBS 0.027403f
C1288 VP.n94 VSUBS 0.027403f
C1289 VP.n95 VSUBS 0.050817f
C1290 VP.n96 VSUBS 0.030747f
C1291 VP.n97 VSUBS 1.21612f
C1292 VP.n98 VSUBS 0.049038f
.ends

