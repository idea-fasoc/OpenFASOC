* NGSPICE file created from diff_pair_sample_0748.ext - technology: sky130A

.subckt diff_pair_sample_0748 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 w_n1674_n4862# sky130_fd_pr__pfet_01v8 ad=7.5933 pd=39.72 as=7.5933 ps=39.72 w=19.47 l=1.43
X1 VDD1.t0 VP.t1 VTAIL.t3 w_n1674_n4862# sky130_fd_pr__pfet_01v8 ad=7.5933 pd=39.72 as=7.5933 ps=39.72 w=19.47 l=1.43
X2 B.t11 B.t9 B.t10 w_n1674_n4862# sky130_fd_pr__pfet_01v8 ad=7.5933 pd=39.72 as=0 ps=0 w=19.47 l=1.43
X3 VDD2.t1 VN.t0 VTAIL.t0 w_n1674_n4862# sky130_fd_pr__pfet_01v8 ad=7.5933 pd=39.72 as=7.5933 ps=39.72 w=19.47 l=1.43
X4 B.t8 B.t6 B.t7 w_n1674_n4862# sky130_fd_pr__pfet_01v8 ad=7.5933 pd=39.72 as=0 ps=0 w=19.47 l=1.43
X5 B.t5 B.t3 B.t4 w_n1674_n4862# sky130_fd_pr__pfet_01v8 ad=7.5933 pd=39.72 as=0 ps=0 w=19.47 l=1.43
X6 B.t2 B.t0 B.t1 w_n1674_n4862# sky130_fd_pr__pfet_01v8 ad=7.5933 pd=39.72 as=0 ps=0 w=19.47 l=1.43
X7 VDD2.t0 VN.t1 VTAIL.t1 w_n1674_n4862# sky130_fd_pr__pfet_01v8 ad=7.5933 pd=39.72 as=7.5933 ps=39.72 w=19.47 l=1.43
R0 VP.n0 VP.t0 483.587
R1 VP.n0 VP.t1 436.373
R2 VP VP.n0 0.146778
R3 VTAIL.n353 VTAIL.n352 585
R4 VTAIL.n350 VTAIL.n349 585
R5 VTAIL.n359 VTAIL.n358 585
R6 VTAIL.n361 VTAIL.n360 585
R7 VTAIL.n346 VTAIL.n345 585
R8 VTAIL.n367 VTAIL.n366 585
R9 VTAIL.n370 VTAIL.n369 585
R10 VTAIL.n368 VTAIL.n342 585
R11 VTAIL.n375 VTAIL.n341 585
R12 VTAIL.n377 VTAIL.n376 585
R13 VTAIL.n379 VTAIL.n378 585
R14 VTAIL.n338 VTAIL.n337 585
R15 VTAIL.n385 VTAIL.n384 585
R16 VTAIL.n387 VTAIL.n386 585
R17 VTAIL.n334 VTAIL.n333 585
R18 VTAIL.n393 VTAIL.n392 585
R19 VTAIL.n395 VTAIL.n394 585
R20 VTAIL.n330 VTAIL.n329 585
R21 VTAIL.n401 VTAIL.n400 585
R22 VTAIL.n403 VTAIL.n402 585
R23 VTAIL.n326 VTAIL.n325 585
R24 VTAIL.n409 VTAIL.n408 585
R25 VTAIL.n411 VTAIL.n410 585
R26 VTAIL.n322 VTAIL.n321 585
R27 VTAIL.n417 VTAIL.n416 585
R28 VTAIL.n419 VTAIL.n418 585
R29 VTAIL.n35 VTAIL.n34 585
R30 VTAIL.n32 VTAIL.n31 585
R31 VTAIL.n41 VTAIL.n40 585
R32 VTAIL.n43 VTAIL.n42 585
R33 VTAIL.n28 VTAIL.n27 585
R34 VTAIL.n49 VTAIL.n48 585
R35 VTAIL.n52 VTAIL.n51 585
R36 VTAIL.n50 VTAIL.n24 585
R37 VTAIL.n57 VTAIL.n23 585
R38 VTAIL.n59 VTAIL.n58 585
R39 VTAIL.n61 VTAIL.n60 585
R40 VTAIL.n20 VTAIL.n19 585
R41 VTAIL.n67 VTAIL.n66 585
R42 VTAIL.n69 VTAIL.n68 585
R43 VTAIL.n16 VTAIL.n15 585
R44 VTAIL.n75 VTAIL.n74 585
R45 VTAIL.n77 VTAIL.n76 585
R46 VTAIL.n12 VTAIL.n11 585
R47 VTAIL.n83 VTAIL.n82 585
R48 VTAIL.n85 VTAIL.n84 585
R49 VTAIL.n8 VTAIL.n7 585
R50 VTAIL.n91 VTAIL.n90 585
R51 VTAIL.n93 VTAIL.n92 585
R52 VTAIL.n4 VTAIL.n3 585
R53 VTAIL.n99 VTAIL.n98 585
R54 VTAIL.n101 VTAIL.n100 585
R55 VTAIL.n313 VTAIL.n312 585
R56 VTAIL.n311 VTAIL.n310 585
R57 VTAIL.n216 VTAIL.n215 585
R58 VTAIL.n305 VTAIL.n304 585
R59 VTAIL.n303 VTAIL.n302 585
R60 VTAIL.n220 VTAIL.n219 585
R61 VTAIL.n297 VTAIL.n296 585
R62 VTAIL.n295 VTAIL.n294 585
R63 VTAIL.n224 VTAIL.n223 585
R64 VTAIL.n289 VTAIL.n288 585
R65 VTAIL.n287 VTAIL.n286 585
R66 VTAIL.n228 VTAIL.n227 585
R67 VTAIL.n281 VTAIL.n280 585
R68 VTAIL.n279 VTAIL.n278 585
R69 VTAIL.n232 VTAIL.n231 585
R70 VTAIL.n273 VTAIL.n272 585
R71 VTAIL.n271 VTAIL.n270 585
R72 VTAIL.n269 VTAIL.n235 585
R73 VTAIL.n239 VTAIL.n236 585
R74 VTAIL.n264 VTAIL.n263 585
R75 VTAIL.n262 VTAIL.n261 585
R76 VTAIL.n241 VTAIL.n240 585
R77 VTAIL.n256 VTAIL.n255 585
R78 VTAIL.n254 VTAIL.n253 585
R79 VTAIL.n245 VTAIL.n244 585
R80 VTAIL.n248 VTAIL.n247 585
R81 VTAIL.n207 VTAIL.n206 585
R82 VTAIL.n205 VTAIL.n204 585
R83 VTAIL.n110 VTAIL.n109 585
R84 VTAIL.n199 VTAIL.n198 585
R85 VTAIL.n197 VTAIL.n196 585
R86 VTAIL.n114 VTAIL.n113 585
R87 VTAIL.n191 VTAIL.n190 585
R88 VTAIL.n189 VTAIL.n188 585
R89 VTAIL.n118 VTAIL.n117 585
R90 VTAIL.n183 VTAIL.n182 585
R91 VTAIL.n181 VTAIL.n180 585
R92 VTAIL.n122 VTAIL.n121 585
R93 VTAIL.n175 VTAIL.n174 585
R94 VTAIL.n173 VTAIL.n172 585
R95 VTAIL.n126 VTAIL.n125 585
R96 VTAIL.n167 VTAIL.n166 585
R97 VTAIL.n165 VTAIL.n164 585
R98 VTAIL.n163 VTAIL.n129 585
R99 VTAIL.n133 VTAIL.n130 585
R100 VTAIL.n158 VTAIL.n157 585
R101 VTAIL.n156 VTAIL.n155 585
R102 VTAIL.n135 VTAIL.n134 585
R103 VTAIL.n150 VTAIL.n149 585
R104 VTAIL.n148 VTAIL.n147 585
R105 VTAIL.n139 VTAIL.n138 585
R106 VTAIL.n142 VTAIL.n141 585
R107 VTAIL.n418 VTAIL.n318 498.474
R108 VTAIL.n100 VTAIL.n0 498.474
R109 VTAIL.n312 VTAIL.n212 498.474
R110 VTAIL.n206 VTAIL.n106 498.474
R111 VTAIL.t1 VTAIL.n351 329.036
R112 VTAIL.t3 VTAIL.n33 329.036
R113 VTAIL.t2 VTAIL.n246 329.036
R114 VTAIL.t0 VTAIL.n140 329.036
R115 VTAIL.n352 VTAIL.n349 171.744
R116 VTAIL.n359 VTAIL.n349 171.744
R117 VTAIL.n360 VTAIL.n359 171.744
R118 VTAIL.n360 VTAIL.n345 171.744
R119 VTAIL.n367 VTAIL.n345 171.744
R120 VTAIL.n369 VTAIL.n367 171.744
R121 VTAIL.n369 VTAIL.n368 171.744
R122 VTAIL.n368 VTAIL.n341 171.744
R123 VTAIL.n377 VTAIL.n341 171.744
R124 VTAIL.n378 VTAIL.n377 171.744
R125 VTAIL.n378 VTAIL.n337 171.744
R126 VTAIL.n385 VTAIL.n337 171.744
R127 VTAIL.n386 VTAIL.n385 171.744
R128 VTAIL.n386 VTAIL.n333 171.744
R129 VTAIL.n393 VTAIL.n333 171.744
R130 VTAIL.n394 VTAIL.n393 171.744
R131 VTAIL.n394 VTAIL.n329 171.744
R132 VTAIL.n401 VTAIL.n329 171.744
R133 VTAIL.n402 VTAIL.n401 171.744
R134 VTAIL.n402 VTAIL.n325 171.744
R135 VTAIL.n409 VTAIL.n325 171.744
R136 VTAIL.n410 VTAIL.n409 171.744
R137 VTAIL.n410 VTAIL.n321 171.744
R138 VTAIL.n417 VTAIL.n321 171.744
R139 VTAIL.n418 VTAIL.n417 171.744
R140 VTAIL.n34 VTAIL.n31 171.744
R141 VTAIL.n41 VTAIL.n31 171.744
R142 VTAIL.n42 VTAIL.n41 171.744
R143 VTAIL.n42 VTAIL.n27 171.744
R144 VTAIL.n49 VTAIL.n27 171.744
R145 VTAIL.n51 VTAIL.n49 171.744
R146 VTAIL.n51 VTAIL.n50 171.744
R147 VTAIL.n50 VTAIL.n23 171.744
R148 VTAIL.n59 VTAIL.n23 171.744
R149 VTAIL.n60 VTAIL.n59 171.744
R150 VTAIL.n60 VTAIL.n19 171.744
R151 VTAIL.n67 VTAIL.n19 171.744
R152 VTAIL.n68 VTAIL.n67 171.744
R153 VTAIL.n68 VTAIL.n15 171.744
R154 VTAIL.n75 VTAIL.n15 171.744
R155 VTAIL.n76 VTAIL.n75 171.744
R156 VTAIL.n76 VTAIL.n11 171.744
R157 VTAIL.n83 VTAIL.n11 171.744
R158 VTAIL.n84 VTAIL.n83 171.744
R159 VTAIL.n84 VTAIL.n7 171.744
R160 VTAIL.n91 VTAIL.n7 171.744
R161 VTAIL.n92 VTAIL.n91 171.744
R162 VTAIL.n92 VTAIL.n3 171.744
R163 VTAIL.n99 VTAIL.n3 171.744
R164 VTAIL.n100 VTAIL.n99 171.744
R165 VTAIL.n312 VTAIL.n311 171.744
R166 VTAIL.n311 VTAIL.n215 171.744
R167 VTAIL.n304 VTAIL.n215 171.744
R168 VTAIL.n304 VTAIL.n303 171.744
R169 VTAIL.n303 VTAIL.n219 171.744
R170 VTAIL.n296 VTAIL.n219 171.744
R171 VTAIL.n296 VTAIL.n295 171.744
R172 VTAIL.n295 VTAIL.n223 171.744
R173 VTAIL.n288 VTAIL.n223 171.744
R174 VTAIL.n288 VTAIL.n287 171.744
R175 VTAIL.n287 VTAIL.n227 171.744
R176 VTAIL.n280 VTAIL.n227 171.744
R177 VTAIL.n280 VTAIL.n279 171.744
R178 VTAIL.n279 VTAIL.n231 171.744
R179 VTAIL.n272 VTAIL.n231 171.744
R180 VTAIL.n272 VTAIL.n271 171.744
R181 VTAIL.n271 VTAIL.n235 171.744
R182 VTAIL.n239 VTAIL.n235 171.744
R183 VTAIL.n263 VTAIL.n239 171.744
R184 VTAIL.n263 VTAIL.n262 171.744
R185 VTAIL.n262 VTAIL.n240 171.744
R186 VTAIL.n255 VTAIL.n240 171.744
R187 VTAIL.n255 VTAIL.n254 171.744
R188 VTAIL.n254 VTAIL.n244 171.744
R189 VTAIL.n247 VTAIL.n244 171.744
R190 VTAIL.n206 VTAIL.n205 171.744
R191 VTAIL.n205 VTAIL.n109 171.744
R192 VTAIL.n198 VTAIL.n109 171.744
R193 VTAIL.n198 VTAIL.n197 171.744
R194 VTAIL.n197 VTAIL.n113 171.744
R195 VTAIL.n190 VTAIL.n113 171.744
R196 VTAIL.n190 VTAIL.n189 171.744
R197 VTAIL.n189 VTAIL.n117 171.744
R198 VTAIL.n182 VTAIL.n117 171.744
R199 VTAIL.n182 VTAIL.n181 171.744
R200 VTAIL.n181 VTAIL.n121 171.744
R201 VTAIL.n174 VTAIL.n121 171.744
R202 VTAIL.n174 VTAIL.n173 171.744
R203 VTAIL.n173 VTAIL.n125 171.744
R204 VTAIL.n166 VTAIL.n125 171.744
R205 VTAIL.n166 VTAIL.n165 171.744
R206 VTAIL.n165 VTAIL.n129 171.744
R207 VTAIL.n133 VTAIL.n129 171.744
R208 VTAIL.n157 VTAIL.n133 171.744
R209 VTAIL.n157 VTAIL.n156 171.744
R210 VTAIL.n156 VTAIL.n134 171.744
R211 VTAIL.n149 VTAIL.n134 171.744
R212 VTAIL.n149 VTAIL.n148 171.744
R213 VTAIL.n148 VTAIL.n138 171.744
R214 VTAIL.n141 VTAIL.n138 171.744
R215 VTAIL.n352 VTAIL.t1 85.8723
R216 VTAIL.n34 VTAIL.t3 85.8723
R217 VTAIL.n247 VTAIL.t2 85.8723
R218 VTAIL.n141 VTAIL.t0 85.8723
R219 VTAIL.n423 VTAIL.n422 35.0944
R220 VTAIL.n105 VTAIL.n104 35.0944
R221 VTAIL.n317 VTAIL.n316 35.0944
R222 VTAIL.n211 VTAIL.n210 35.0944
R223 VTAIL.n211 VTAIL.n105 32.1858
R224 VTAIL.n423 VTAIL.n317 30.6686
R225 VTAIL.n376 VTAIL.n375 13.1884
R226 VTAIL.n58 VTAIL.n57 13.1884
R227 VTAIL.n270 VTAIL.n269 13.1884
R228 VTAIL.n164 VTAIL.n163 13.1884
R229 VTAIL.n374 VTAIL.n342 12.8005
R230 VTAIL.n379 VTAIL.n340 12.8005
R231 VTAIL.n420 VTAIL.n419 12.8005
R232 VTAIL.n56 VTAIL.n24 12.8005
R233 VTAIL.n61 VTAIL.n22 12.8005
R234 VTAIL.n102 VTAIL.n101 12.8005
R235 VTAIL.n314 VTAIL.n313 12.8005
R236 VTAIL.n273 VTAIL.n234 12.8005
R237 VTAIL.n268 VTAIL.n236 12.8005
R238 VTAIL.n208 VTAIL.n207 12.8005
R239 VTAIL.n167 VTAIL.n128 12.8005
R240 VTAIL.n162 VTAIL.n130 12.8005
R241 VTAIL.n371 VTAIL.n370 12.0247
R242 VTAIL.n380 VTAIL.n338 12.0247
R243 VTAIL.n416 VTAIL.n320 12.0247
R244 VTAIL.n53 VTAIL.n52 12.0247
R245 VTAIL.n62 VTAIL.n20 12.0247
R246 VTAIL.n98 VTAIL.n2 12.0247
R247 VTAIL.n310 VTAIL.n214 12.0247
R248 VTAIL.n274 VTAIL.n232 12.0247
R249 VTAIL.n265 VTAIL.n264 12.0247
R250 VTAIL.n204 VTAIL.n108 12.0247
R251 VTAIL.n168 VTAIL.n126 12.0247
R252 VTAIL.n159 VTAIL.n158 12.0247
R253 VTAIL.n366 VTAIL.n344 11.249
R254 VTAIL.n384 VTAIL.n383 11.249
R255 VTAIL.n415 VTAIL.n322 11.249
R256 VTAIL.n48 VTAIL.n26 11.249
R257 VTAIL.n66 VTAIL.n65 11.249
R258 VTAIL.n97 VTAIL.n4 11.249
R259 VTAIL.n309 VTAIL.n216 11.249
R260 VTAIL.n278 VTAIL.n277 11.249
R261 VTAIL.n261 VTAIL.n238 11.249
R262 VTAIL.n203 VTAIL.n110 11.249
R263 VTAIL.n172 VTAIL.n171 11.249
R264 VTAIL.n155 VTAIL.n132 11.249
R265 VTAIL.n353 VTAIL.n351 10.7239
R266 VTAIL.n35 VTAIL.n33 10.7239
R267 VTAIL.n248 VTAIL.n246 10.7239
R268 VTAIL.n142 VTAIL.n140 10.7239
R269 VTAIL.n365 VTAIL.n346 10.4732
R270 VTAIL.n387 VTAIL.n336 10.4732
R271 VTAIL.n412 VTAIL.n411 10.4732
R272 VTAIL.n47 VTAIL.n28 10.4732
R273 VTAIL.n69 VTAIL.n18 10.4732
R274 VTAIL.n94 VTAIL.n93 10.4732
R275 VTAIL.n306 VTAIL.n305 10.4732
R276 VTAIL.n281 VTAIL.n230 10.4732
R277 VTAIL.n260 VTAIL.n241 10.4732
R278 VTAIL.n200 VTAIL.n199 10.4732
R279 VTAIL.n175 VTAIL.n124 10.4732
R280 VTAIL.n154 VTAIL.n135 10.4732
R281 VTAIL.n362 VTAIL.n361 9.69747
R282 VTAIL.n388 VTAIL.n334 9.69747
R283 VTAIL.n408 VTAIL.n324 9.69747
R284 VTAIL.n44 VTAIL.n43 9.69747
R285 VTAIL.n70 VTAIL.n16 9.69747
R286 VTAIL.n90 VTAIL.n6 9.69747
R287 VTAIL.n302 VTAIL.n218 9.69747
R288 VTAIL.n282 VTAIL.n228 9.69747
R289 VTAIL.n257 VTAIL.n256 9.69747
R290 VTAIL.n196 VTAIL.n112 9.69747
R291 VTAIL.n176 VTAIL.n122 9.69747
R292 VTAIL.n151 VTAIL.n150 9.69747
R293 VTAIL.n422 VTAIL.n421 9.45567
R294 VTAIL.n104 VTAIL.n103 9.45567
R295 VTAIL.n316 VTAIL.n315 9.45567
R296 VTAIL.n210 VTAIL.n209 9.45567
R297 VTAIL.n397 VTAIL.n396 9.3005
R298 VTAIL.n332 VTAIL.n331 9.3005
R299 VTAIL.n391 VTAIL.n390 9.3005
R300 VTAIL.n389 VTAIL.n388 9.3005
R301 VTAIL.n336 VTAIL.n335 9.3005
R302 VTAIL.n383 VTAIL.n382 9.3005
R303 VTAIL.n381 VTAIL.n380 9.3005
R304 VTAIL.n340 VTAIL.n339 9.3005
R305 VTAIL.n355 VTAIL.n354 9.3005
R306 VTAIL.n357 VTAIL.n356 9.3005
R307 VTAIL.n348 VTAIL.n347 9.3005
R308 VTAIL.n363 VTAIL.n362 9.3005
R309 VTAIL.n365 VTAIL.n364 9.3005
R310 VTAIL.n344 VTAIL.n343 9.3005
R311 VTAIL.n372 VTAIL.n371 9.3005
R312 VTAIL.n374 VTAIL.n373 9.3005
R313 VTAIL.n399 VTAIL.n398 9.3005
R314 VTAIL.n328 VTAIL.n327 9.3005
R315 VTAIL.n405 VTAIL.n404 9.3005
R316 VTAIL.n407 VTAIL.n406 9.3005
R317 VTAIL.n324 VTAIL.n323 9.3005
R318 VTAIL.n413 VTAIL.n412 9.3005
R319 VTAIL.n415 VTAIL.n414 9.3005
R320 VTAIL.n320 VTAIL.n319 9.3005
R321 VTAIL.n421 VTAIL.n420 9.3005
R322 VTAIL.n79 VTAIL.n78 9.3005
R323 VTAIL.n14 VTAIL.n13 9.3005
R324 VTAIL.n73 VTAIL.n72 9.3005
R325 VTAIL.n71 VTAIL.n70 9.3005
R326 VTAIL.n18 VTAIL.n17 9.3005
R327 VTAIL.n65 VTAIL.n64 9.3005
R328 VTAIL.n63 VTAIL.n62 9.3005
R329 VTAIL.n22 VTAIL.n21 9.3005
R330 VTAIL.n37 VTAIL.n36 9.3005
R331 VTAIL.n39 VTAIL.n38 9.3005
R332 VTAIL.n30 VTAIL.n29 9.3005
R333 VTAIL.n45 VTAIL.n44 9.3005
R334 VTAIL.n47 VTAIL.n46 9.3005
R335 VTAIL.n26 VTAIL.n25 9.3005
R336 VTAIL.n54 VTAIL.n53 9.3005
R337 VTAIL.n56 VTAIL.n55 9.3005
R338 VTAIL.n81 VTAIL.n80 9.3005
R339 VTAIL.n10 VTAIL.n9 9.3005
R340 VTAIL.n87 VTAIL.n86 9.3005
R341 VTAIL.n89 VTAIL.n88 9.3005
R342 VTAIL.n6 VTAIL.n5 9.3005
R343 VTAIL.n95 VTAIL.n94 9.3005
R344 VTAIL.n97 VTAIL.n96 9.3005
R345 VTAIL.n2 VTAIL.n1 9.3005
R346 VTAIL.n103 VTAIL.n102 9.3005
R347 VTAIL.n250 VTAIL.n249 9.3005
R348 VTAIL.n252 VTAIL.n251 9.3005
R349 VTAIL.n243 VTAIL.n242 9.3005
R350 VTAIL.n258 VTAIL.n257 9.3005
R351 VTAIL.n260 VTAIL.n259 9.3005
R352 VTAIL.n238 VTAIL.n237 9.3005
R353 VTAIL.n266 VTAIL.n265 9.3005
R354 VTAIL.n268 VTAIL.n267 9.3005
R355 VTAIL.n222 VTAIL.n221 9.3005
R356 VTAIL.n299 VTAIL.n298 9.3005
R357 VTAIL.n301 VTAIL.n300 9.3005
R358 VTAIL.n218 VTAIL.n217 9.3005
R359 VTAIL.n307 VTAIL.n306 9.3005
R360 VTAIL.n309 VTAIL.n308 9.3005
R361 VTAIL.n214 VTAIL.n213 9.3005
R362 VTAIL.n315 VTAIL.n314 9.3005
R363 VTAIL.n293 VTAIL.n292 9.3005
R364 VTAIL.n291 VTAIL.n290 9.3005
R365 VTAIL.n226 VTAIL.n225 9.3005
R366 VTAIL.n285 VTAIL.n284 9.3005
R367 VTAIL.n283 VTAIL.n282 9.3005
R368 VTAIL.n230 VTAIL.n229 9.3005
R369 VTAIL.n277 VTAIL.n276 9.3005
R370 VTAIL.n275 VTAIL.n274 9.3005
R371 VTAIL.n234 VTAIL.n233 9.3005
R372 VTAIL.n144 VTAIL.n143 9.3005
R373 VTAIL.n146 VTAIL.n145 9.3005
R374 VTAIL.n137 VTAIL.n136 9.3005
R375 VTAIL.n152 VTAIL.n151 9.3005
R376 VTAIL.n154 VTAIL.n153 9.3005
R377 VTAIL.n132 VTAIL.n131 9.3005
R378 VTAIL.n160 VTAIL.n159 9.3005
R379 VTAIL.n162 VTAIL.n161 9.3005
R380 VTAIL.n116 VTAIL.n115 9.3005
R381 VTAIL.n193 VTAIL.n192 9.3005
R382 VTAIL.n195 VTAIL.n194 9.3005
R383 VTAIL.n112 VTAIL.n111 9.3005
R384 VTAIL.n201 VTAIL.n200 9.3005
R385 VTAIL.n203 VTAIL.n202 9.3005
R386 VTAIL.n108 VTAIL.n107 9.3005
R387 VTAIL.n209 VTAIL.n208 9.3005
R388 VTAIL.n187 VTAIL.n186 9.3005
R389 VTAIL.n185 VTAIL.n184 9.3005
R390 VTAIL.n120 VTAIL.n119 9.3005
R391 VTAIL.n179 VTAIL.n178 9.3005
R392 VTAIL.n177 VTAIL.n176 9.3005
R393 VTAIL.n124 VTAIL.n123 9.3005
R394 VTAIL.n171 VTAIL.n170 9.3005
R395 VTAIL.n169 VTAIL.n168 9.3005
R396 VTAIL.n128 VTAIL.n127 9.3005
R397 VTAIL.n358 VTAIL.n348 8.92171
R398 VTAIL.n392 VTAIL.n391 8.92171
R399 VTAIL.n407 VTAIL.n326 8.92171
R400 VTAIL.n40 VTAIL.n30 8.92171
R401 VTAIL.n74 VTAIL.n73 8.92171
R402 VTAIL.n89 VTAIL.n8 8.92171
R403 VTAIL.n301 VTAIL.n220 8.92171
R404 VTAIL.n286 VTAIL.n285 8.92171
R405 VTAIL.n253 VTAIL.n243 8.92171
R406 VTAIL.n195 VTAIL.n114 8.92171
R407 VTAIL.n180 VTAIL.n179 8.92171
R408 VTAIL.n147 VTAIL.n137 8.92171
R409 VTAIL.n357 VTAIL.n350 8.14595
R410 VTAIL.n395 VTAIL.n332 8.14595
R411 VTAIL.n404 VTAIL.n403 8.14595
R412 VTAIL.n39 VTAIL.n32 8.14595
R413 VTAIL.n77 VTAIL.n14 8.14595
R414 VTAIL.n86 VTAIL.n85 8.14595
R415 VTAIL.n298 VTAIL.n297 8.14595
R416 VTAIL.n289 VTAIL.n226 8.14595
R417 VTAIL.n252 VTAIL.n245 8.14595
R418 VTAIL.n192 VTAIL.n191 8.14595
R419 VTAIL.n183 VTAIL.n120 8.14595
R420 VTAIL.n146 VTAIL.n139 8.14595
R421 VTAIL.n422 VTAIL.n318 7.75445
R422 VTAIL.n104 VTAIL.n0 7.75445
R423 VTAIL.n316 VTAIL.n212 7.75445
R424 VTAIL.n210 VTAIL.n106 7.75445
R425 VTAIL.n354 VTAIL.n353 7.3702
R426 VTAIL.n396 VTAIL.n330 7.3702
R427 VTAIL.n400 VTAIL.n328 7.3702
R428 VTAIL.n36 VTAIL.n35 7.3702
R429 VTAIL.n78 VTAIL.n12 7.3702
R430 VTAIL.n82 VTAIL.n10 7.3702
R431 VTAIL.n294 VTAIL.n222 7.3702
R432 VTAIL.n290 VTAIL.n224 7.3702
R433 VTAIL.n249 VTAIL.n248 7.3702
R434 VTAIL.n188 VTAIL.n116 7.3702
R435 VTAIL.n184 VTAIL.n118 7.3702
R436 VTAIL.n143 VTAIL.n142 7.3702
R437 VTAIL.n399 VTAIL.n330 6.59444
R438 VTAIL.n400 VTAIL.n399 6.59444
R439 VTAIL.n81 VTAIL.n12 6.59444
R440 VTAIL.n82 VTAIL.n81 6.59444
R441 VTAIL.n294 VTAIL.n293 6.59444
R442 VTAIL.n293 VTAIL.n224 6.59444
R443 VTAIL.n188 VTAIL.n187 6.59444
R444 VTAIL.n187 VTAIL.n118 6.59444
R445 VTAIL.n420 VTAIL.n318 6.08283
R446 VTAIL.n102 VTAIL.n0 6.08283
R447 VTAIL.n314 VTAIL.n212 6.08283
R448 VTAIL.n208 VTAIL.n106 6.08283
R449 VTAIL.n354 VTAIL.n350 5.81868
R450 VTAIL.n396 VTAIL.n395 5.81868
R451 VTAIL.n403 VTAIL.n328 5.81868
R452 VTAIL.n36 VTAIL.n32 5.81868
R453 VTAIL.n78 VTAIL.n77 5.81868
R454 VTAIL.n85 VTAIL.n10 5.81868
R455 VTAIL.n297 VTAIL.n222 5.81868
R456 VTAIL.n290 VTAIL.n289 5.81868
R457 VTAIL.n249 VTAIL.n245 5.81868
R458 VTAIL.n191 VTAIL.n116 5.81868
R459 VTAIL.n184 VTAIL.n183 5.81868
R460 VTAIL.n143 VTAIL.n139 5.81868
R461 VTAIL.n358 VTAIL.n357 5.04292
R462 VTAIL.n392 VTAIL.n332 5.04292
R463 VTAIL.n404 VTAIL.n326 5.04292
R464 VTAIL.n40 VTAIL.n39 5.04292
R465 VTAIL.n74 VTAIL.n14 5.04292
R466 VTAIL.n86 VTAIL.n8 5.04292
R467 VTAIL.n298 VTAIL.n220 5.04292
R468 VTAIL.n286 VTAIL.n226 5.04292
R469 VTAIL.n253 VTAIL.n252 5.04292
R470 VTAIL.n192 VTAIL.n114 5.04292
R471 VTAIL.n180 VTAIL.n120 5.04292
R472 VTAIL.n147 VTAIL.n146 5.04292
R473 VTAIL.n361 VTAIL.n348 4.26717
R474 VTAIL.n391 VTAIL.n334 4.26717
R475 VTAIL.n408 VTAIL.n407 4.26717
R476 VTAIL.n43 VTAIL.n30 4.26717
R477 VTAIL.n73 VTAIL.n16 4.26717
R478 VTAIL.n90 VTAIL.n89 4.26717
R479 VTAIL.n302 VTAIL.n301 4.26717
R480 VTAIL.n285 VTAIL.n228 4.26717
R481 VTAIL.n256 VTAIL.n243 4.26717
R482 VTAIL.n196 VTAIL.n195 4.26717
R483 VTAIL.n179 VTAIL.n122 4.26717
R484 VTAIL.n150 VTAIL.n137 4.26717
R485 VTAIL.n362 VTAIL.n346 3.49141
R486 VTAIL.n388 VTAIL.n387 3.49141
R487 VTAIL.n411 VTAIL.n324 3.49141
R488 VTAIL.n44 VTAIL.n28 3.49141
R489 VTAIL.n70 VTAIL.n69 3.49141
R490 VTAIL.n93 VTAIL.n6 3.49141
R491 VTAIL.n305 VTAIL.n218 3.49141
R492 VTAIL.n282 VTAIL.n281 3.49141
R493 VTAIL.n257 VTAIL.n241 3.49141
R494 VTAIL.n199 VTAIL.n112 3.49141
R495 VTAIL.n176 VTAIL.n175 3.49141
R496 VTAIL.n151 VTAIL.n135 3.49141
R497 VTAIL.n366 VTAIL.n365 2.71565
R498 VTAIL.n384 VTAIL.n336 2.71565
R499 VTAIL.n412 VTAIL.n322 2.71565
R500 VTAIL.n48 VTAIL.n47 2.71565
R501 VTAIL.n66 VTAIL.n18 2.71565
R502 VTAIL.n94 VTAIL.n4 2.71565
R503 VTAIL.n306 VTAIL.n216 2.71565
R504 VTAIL.n278 VTAIL.n230 2.71565
R505 VTAIL.n261 VTAIL.n260 2.71565
R506 VTAIL.n200 VTAIL.n110 2.71565
R507 VTAIL.n172 VTAIL.n124 2.71565
R508 VTAIL.n155 VTAIL.n154 2.71565
R509 VTAIL.n250 VTAIL.n246 2.41282
R510 VTAIL.n144 VTAIL.n140 2.41282
R511 VTAIL.n355 VTAIL.n351 2.41282
R512 VTAIL.n37 VTAIL.n33 2.41282
R513 VTAIL.n370 VTAIL.n344 1.93989
R514 VTAIL.n383 VTAIL.n338 1.93989
R515 VTAIL.n416 VTAIL.n415 1.93989
R516 VTAIL.n52 VTAIL.n26 1.93989
R517 VTAIL.n65 VTAIL.n20 1.93989
R518 VTAIL.n98 VTAIL.n97 1.93989
R519 VTAIL.n310 VTAIL.n309 1.93989
R520 VTAIL.n277 VTAIL.n232 1.93989
R521 VTAIL.n264 VTAIL.n238 1.93989
R522 VTAIL.n204 VTAIL.n203 1.93989
R523 VTAIL.n171 VTAIL.n126 1.93989
R524 VTAIL.n158 VTAIL.n132 1.93989
R525 VTAIL.n317 VTAIL.n211 1.22895
R526 VTAIL.n371 VTAIL.n342 1.16414
R527 VTAIL.n380 VTAIL.n379 1.16414
R528 VTAIL.n419 VTAIL.n320 1.16414
R529 VTAIL.n53 VTAIL.n24 1.16414
R530 VTAIL.n62 VTAIL.n61 1.16414
R531 VTAIL.n101 VTAIL.n2 1.16414
R532 VTAIL.n313 VTAIL.n214 1.16414
R533 VTAIL.n274 VTAIL.n273 1.16414
R534 VTAIL.n265 VTAIL.n236 1.16414
R535 VTAIL.n207 VTAIL.n108 1.16414
R536 VTAIL.n168 VTAIL.n167 1.16414
R537 VTAIL.n159 VTAIL.n130 1.16414
R538 VTAIL VTAIL.n105 0.907828
R539 VTAIL.n375 VTAIL.n374 0.388379
R540 VTAIL.n376 VTAIL.n340 0.388379
R541 VTAIL.n57 VTAIL.n56 0.388379
R542 VTAIL.n58 VTAIL.n22 0.388379
R543 VTAIL.n270 VTAIL.n234 0.388379
R544 VTAIL.n269 VTAIL.n268 0.388379
R545 VTAIL.n164 VTAIL.n128 0.388379
R546 VTAIL.n163 VTAIL.n162 0.388379
R547 VTAIL VTAIL.n423 0.321621
R548 VTAIL.n356 VTAIL.n355 0.155672
R549 VTAIL.n356 VTAIL.n347 0.155672
R550 VTAIL.n363 VTAIL.n347 0.155672
R551 VTAIL.n364 VTAIL.n363 0.155672
R552 VTAIL.n364 VTAIL.n343 0.155672
R553 VTAIL.n372 VTAIL.n343 0.155672
R554 VTAIL.n373 VTAIL.n372 0.155672
R555 VTAIL.n373 VTAIL.n339 0.155672
R556 VTAIL.n381 VTAIL.n339 0.155672
R557 VTAIL.n382 VTAIL.n381 0.155672
R558 VTAIL.n382 VTAIL.n335 0.155672
R559 VTAIL.n389 VTAIL.n335 0.155672
R560 VTAIL.n390 VTAIL.n389 0.155672
R561 VTAIL.n390 VTAIL.n331 0.155672
R562 VTAIL.n397 VTAIL.n331 0.155672
R563 VTAIL.n398 VTAIL.n397 0.155672
R564 VTAIL.n398 VTAIL.n327 0.155672
R565 VTAIL.n405 VTAIL.n327 0.155672
R566 VTAIL.n406 VTAIL.n405 0.155672
R567 VTAIL.n406 VTAIL.n323 0.155672
R568 VTAIL.n413 VTAIL.n323 0.155672
R569 VTAIL.n414 VTAIL.n413 0.155672
R570 VTAIL.n414 VTAIL.n319 0.155672
R571 VTAIL.n421 VTAIL.n319 0.155672
R572 VTAIL.n38 VTAIL.n37 0.155672
R573 VTAIL.n38 VTAIL.n29 0.155672
R574 VTAIL.n45 VTAIL.n29 0.155672
R575 VTAIL.n46 VTAIL.n45 0.155672
R576 VTAIL.n46 VTAIL.n25 0.155672
R577 VTAIL.n54 VTAIL.n25 0.155672
R578 VTAIL.n55 VTAIL.n54 0.155672
R579 VTAIL.n55 VTAIL.n21 0.155672
R580 VTAIL.n63 VTAIL.n21 0.155672
R581 VTAIL.n64 VTAIL.n63 0.155672
R582 VTAIL.n64 VTAIL.n17 0.155672
R583 VTAIL.n71 VTAIL.n17 0.155672
R584 VTAIL.n72 VTAIL.n71 0.155672
R585 VTAIL.n72 VTAIL.n13 0.155672
R586 VTAIL.n79 VTAIL.n13 0.155672
R587 VTAIL.n80 VTAIL.n79 0.155672
R588 VTAIL.n80 VTAIL.n9 0.155672
R589 VTAIL.n87 VTAIL.n9 0.155672
R590 VTAIL.n88 VTAIL.n87 0.155672
R591 VTAIL.n88 VTAIL.n5 0.155672
R592 VTAIL.n95 VTAIL.n5 0.155672
R593 VTAIL.n96 VTAIL.n95 0.155672
R594 VTAIL.n96 VTAIL.n1 0.155672
R595 VTAIL.n103 VTAIL.n1 0.155672
R596 VTAIL.n315 VTAIL.n213 0.155672
R597 VTAIL.n308 VTAIL.n213 0.155672
R598 VTAIL.n308 VTAIL.n307 0.155672
R599 VTAIL.n307 VTAIL.n217 0.155672
R600 VTAIL.n300 VTAIL.n217 0.155672
R601 VTAIL.n300 VTAIL.n299 0.155672
R602 VTAIL.n299 VTAIL.n221 0.155672
R603 VTAIL.n292 VTAIL.n221 0.155672
R604 VTAIL.n292 VTAIL.n291 0.155672
R605 VTAIL.n291 VTAIL.n225 0.155672
R606 VTAIL.n284 VTAIL.n225 0.155672
R607 VTAIL.n284 VTAIL.n283 0.155672
R608 VTAIL.n283 VTAIL.n229 0.155672
R609 VTAIL.n276 VTAIL.n229 0.155672
R610 VTAIL.n276 VTAIL.n275 0.155672
R611 VTAIL.n275 VTAIL.n233 0.155672
R612 VTAIL.n267 VTAIL.n233 0.155672
R613 VTAIL.n267 VTAIL.n266 0.155672
R614 VTAIL.n266 VTAIL.n237 0.155672
R615 VTAIL.n259 VTAIL.n237 0.155672
R616 VTAIL.n259 VTAIL.n258 0.155672
R617 VTAIL.n258 VTAIL.n242 0.155672
R618 VTAIL.n251 VTAIL.n242 0.155672
R619 VTAIL.n251 VTAIL.n250 0.155672
R620 VTAIL.n209 VTAIL.n107 0.155672
R621 VTAIL.n202 VTAIL.n107 0.155672
R622 VTAIL.n202 VTAIL.n201 0.155672
R623 VTAIL.n201 VTAIL.n111 0.155672
R624 VTAIL.n194 VTAIL.n111 0.155672
R625 VTAIL.n194 VTAIL.n193 0.155672
R626 VTAIL.n193 VTAIL.n115 0.155672
R627 VTAIL.n186 VTAIL.n115 0.155672
R628 VTAIL.n186 VTAIL.n185 0.155672
R629 VTAIL.n185 VTAIL.n119 0.155672
R630 VTAIL.n178 VTAIL.n119 0.155672
R631 VTAIL.n178 VTAIL.n177 0.155672
R632 VTAIL.n177 VTAIL.n123 0.155672
R633 VTAIL.n170 VTAIL.n123 0.155672
R634 VTAIL.n170 VTAIL.n169 0.155672
R635 VTAIL.n169 VTAIL.n127 0.155672
R636 VTAIL.n161 VTAIL.n127 0.155672
R637 VTAIL.n161 VTAIL.n160 0.155672
R638 VTAIL.n160 VTAIL.n131 0.155672
R639 VTAIL.n153 VTAIL.n131 0.155672
R640 VTAIL.n153 VTAIL.n152 0.155672
R641 VTAIL.n152 VTAIL.n136 0.155672
R642 VTAIL.n145 VTAIL.n136 0.155672
R643 VTAIL.n145 VTAIL.n144 0.155672
R644 VDD1.n101 VDD1.n100 585
R645 VDD1.n99 VDD1.n98 585
R646 VDD1.n4 VDD1.n3 585
R647 VDD1.n93 VDD1.n92 585
R648 VDD1.n91 VDD1.n90 585
R649 VDD1.n8 VDD1.n7 585
R650 VDD1.n85 VDD1.n84 585
R651 VDD1.n83 VDD1.n82 585
R652 VDD1.n12 VDD1.n11 585
R653 VDD1.n77 VDD1.n76 585
R654 VDD1.n75 VDD1.n74 585
R655 VDD1.n16 VDD1.n15 585
R656 VDD1.n69 VDD1.n68 585
R657 VDD1.n67 VDD1.n66 585
R658 VDD1.n20 VDD1.n19 585
R659 VDD1.n61 VDD1.n60 585
R660 VDD1.n59 VDD1.n58 585
R661 VDD1.n57 VDD1.n23 585
R662 VDD1.n27 VDD1.n24 585
R663 VDD1.n52 VDD1.n51 585
R664 VDD1.n50 VDD1.n49 585
R665 VDD1.n29 VDD1.n28 585
R666 VDD1.n44 VDD1.n43 585
R667 VDD1.n42 VDD1.n41 585
R668 VDD1.n33 VDD1.n32 585
R669 VDD1.n36 VDD1.n35 585
R670 VDD1.n140 VDD1.n139 585
R671 VDD1.n137 VDD1.n136 585
R672 VDD1.n146 VDD1.n145 585
R673 VDD1.n148 VDD1.n147 585
R674 VDD1.n133 VDD1.n132 585
R675 VDD1.n154 VDD1.n153 585
R676 VDD1.n157 VDD1.n156 585
R677 VDD1.n155 VDD1.n129 585
R678 VDD1.n162 VDD1.n128 585
R679 VDD1.n164 VDD1.n163 585
R680 VDD1.n166 VDD1.n165 585
R681 VDD1.n125 VDD1.n124 585
R682 VDD1.n172 VDD1.n171 585
R683 VDD1.n174 VDD1.n173 585
R684 VDD1.n121 VDD1.n120 585
R685 VDD1.n180 VDD1.n179 585
R686 VDD1.n182 VDD1.n181 585
R687 VDD1.n117 VDD1.n116 585
R688 VDD1.n188 VDD1.n187 585
R689 VDD1.n190 VDD1.n189 585
R690 VDD1.n113 VDD1.n112 585
R691 VDD1.n196 VDD1.n195 585
R692 VDD1.n198 VDD1.n197 585
R693 VDD1.n109 VDD1.n108 585
R694 VDD1.n204 VDD1.n203 585
R695 VDD1.n206 VDD1.n205 585
R696 VDD1.n100 VDD1.n0 498.474
R697 VDD1.n205 VDD1.n105 498.474
R698 VDD1.t1 VDD1.n34 329.036
R699 VDD1.t0 VDD1.n138 329.036
R700 VDD1.n100 VDD1.n99 171.744
R701 VDD1.n99 VDD1.n3 171.744
R702 VDD1.n92 VDD1.n3 171.744
R703 VDD1.n92 VDD1.n91 171.744
R704 VDD1.n91 VDD1.n7 171.744
R705 VDD1.n84 VDD1.n7 171.744
R706 VDD1.n84 VDD1.n83 171.744
R707 VDD1.n83 VDD1.n11 171.744
R708 VDD1.n76 VDD1.n11 171.744
R709 VDD1.n76 VDD1.n75 171.744
R710 VDD1.n75 VDD1.n15 171.744
R711 VDD1.n68 VDD1.n15 171.744
R712 VDD1.n68 VDD1.n67 171.744
R713 VDD1.n67 VDD1.n19 171.744
R714 VDD1.n60 VDD1.n19 171.744
R715 VDD1.n60 VDD1.n59 171.744
R716 VDD1.n59 VDD1.n23 171.744
R717 VDD1.n27 VDD1.n23 171.744
R718 VDD1.n51 VDD1.n27 171.744
R719 VDD1.n51 VDD1.n50 171.744
R720 VDD1.n50 VDD1.n28 171.744
R721 VDD1.n43 VDD1.n28 171.744
R722 VDD1.n43 VDD1.n42 171.744
R723 VDD1.n42 VDD1.n32 171.744
R724 VDD1.n35 VDD1.n32 171.744
R725 VDD1.n139 VDD1.n136 171.744
R726 VDD1.n146 VDD1.n136 171.744
R727 VDD1.n147 VDD1.n146 171.744
R728 VDD1.n147 VDD1.n132 171.744
R729 VDD1.n154 VDD1.n132 171.744
R730 VDD1.n156 VDD1.n154 171.744
R731 VDD1.n156 VDD1.n155 171.744
R732 VDD1.n155 VDD1.n128 171.744
R733 VDD1.n164 VDD1.n128 171.744
R734 VDD1.n165 VDD1.n164 171.744
R735 VDD1.n165 VDD1.n124 171.744
R736 VDD1.n172 VDD1.n124 171.744
R737 VDD1.n173 VDD1.n172 171.744
R738 VDD1.n173 VDD1.n120 171.744
R739 VDD1.n180 VDD1.n120 171.744
R740 VDD1.n181 VDD1.n180 171.744
R741 VDD1.n181 VDD1.n116 171.744
R742 VDD1.n188 VDD1.n116 171.744
R743 VDD1.n189 VDD1.n188 171.744
R744 VDD1.n189 VDD1.n112 171.744
R745 VDD1.n196 VDD1.n112 171.744
R746 VDD1.n197 VDD1.n196 171.744
R747 VDD1.n197 VDD1.n108 171.744
R748 VDD1.n204 VDD1.n108 171.744
R749 VDD1.n205 VDD1.n204 171.744
R750 VDD1 VDD1.n209 96.1558
R751 VDD1.n35 VDD1.t1 85.8723
R752 VDD1.n139 VDD1.t0 85.8723
R753 VDD1 VDD1.n104 52.2107
R754 VDD1.n58 VDD1.n57 13.1884
R755 VDD1.n163 VDD1.n162 13.1884
R756 VDD1.n102 VDD1.n101 12.8005
R757 VDD1.n61 VDD1.n22 12.8005
R758 VDD1.n56 VDD1.n24 12.8005
R759 VDD1.n161 VDD1.n129 12.8005
R760 VDD1.n166 VDD1.n127 12.8005
R761 VDD1.n207 VDD1.n206 12.8005
R762 VDD1.n98 VDD1.n2 12.0247
R763 VDD1.n62 VDD1.n20 12.0247
R764 VDD1.n53 VDD1.n52 12.0247
R765 VDD1.n158 VDD1.n157 12.0247
R766 VDD1.n167 VDD1.n125 12.0247
R767 VDD1.n203 VDD1.n107 12.0247
R768 VDD1.n97 VDD1.n4 11.249
R769 VDD1.n66 VDD1.n65 11.249
R770 VDD1.n49 VDD1.n26 11.249
R771 VDD1.n153 VDD1.n131 11.249
R772 VDD1.n171 VDD1.n170 11.249
R773 VDD1.n202 VDD1.n109 11.249
R774 VDD1.n36 VDD1.n34 10.7239
R775 VDD1.n140 VDD1.n138 10.7239
R776 VDD1.n94 VDD1.n93 10.4732
R777 VDD1.n69 VDD1.n18 10.4732
R778 VDD1.n48 VDD1.n29 10.4732
R779 VDD1.n152 VDD1.n133 10.4732
R780 VDD1.n174 VDD1.n123 10.4732
R781 VDD1.n199 VDD1.n198 10.4732
R782 VDD1.n90 VDD1.n6 9.69747
R783 VDD1.n70 VDD1.n16 9.69747
R784 VDD1.n45 VDD1.n44 9.69747
R785 VDD1.n149 VDD1.n148 9.69747
R786 VDD1.n175 VDD1.n121 9.69747
R787 VDD1.n195 VDD1.n111 9.69747
R788 VDD1.n104 VDD1.n103 9.45567
R789 VDD1.n209 VDD1.n208 9.45567
R790 VDD1.n38 VDD1.n37 9.3005
R791 VDD1.n40 VDD1.n39 9.3005
R792 VDD1.n31 VDD1.n30 9.3005
R793 VDD1.n46 VDD1.n45 9.3005
R794 VDD1.n48 VDD1.n47 9.3005
R795 VDD1.n26 VDD1.n25 9.3005
R796 VDD1.n54 VDD1.n53 9.3005
R797 VDD1.n56 VDD1.n55 9.3005
R798 VDD1.n10 VDD1.n9 9.3005
R799 VDD1.n87 VDD1.n86 9.3005
R800 VDD1.n89 VDD1.n88 9.3005
R801 VDD1.n6 VDD1.n5 9.3005
R802 VDD1.n95 VDD1.n94 9.3005
R803 VDD1.n97 VDD1.n96 9.3005
R804 VDD1.n2 VDD1.n1 9.3005
R805 VDD1.n103 VDD1.n102 9.3005
R806 VDD1.n81 VDD1.n80 9.3005
R807 VDD1.n79 VDD1.n78 9.3005
R808 VDD1.n14 VDD1.n13 9.3005
R809 VDD1.n73 VDD1.n72 9.3005
R810 VDD1.n71 VDD1.n70 9.3005
R811 VDD1.n18 VDD1.n17 9.3005
R812 VDD1.n65 VDD1.n64 9.3005
R813 VDD1.n63 VDD1.n62 9.3005
R814 VDD1.n22 VDD1.n21 9.3005
R815 VDD1.n184 VDD1.n183 9.3005
R816 VDD1.n119 VDD1.n118 9.3005
R817 VDD1.n178 VDD1.n177 9.3005
R818 VDD1.n176 VDD1.n175 9.3005
R819 VDD1.n123 VDD1.n122 9.3005
R820 VDD1.n170 VDD1.n169 9.3005
R821 VDD1.n168 VDD1.n167 9.3005
R822 VDD1.n127 VDD1.n126 9.3005
R823 VDD1.n142 VDD1.n141 9.3005
R824 VDD1.n144 VDD1.n143 9.3005
R825 VDD1.n135 VDD1.n134 9.3005
R826 VDD1.n150 VDD1.n149 9.3005
R827 VDD1.n152 VDD1.n151 9.3005
R828 VDD1.n131 VDD1.n130 9.3005
R829 VDD1.n159 VDD1.n158 9.3005
R830 VDD1.n161 VDD1.n160 9.3005
R831 VDD1.n186 VDD1.n185 9.3005
R832 VDD1.n115 VDD1.n114 9.3005
R833 VDD1.n192 VDD1.n191 9.3005
R834 VDD1.n194 VDD1.n193 9.3005
R835 VDD1.n111 VDD1.n110 9.3005
R836 VDD1.n200 VDD1.n199 9.3005
R837 VDD1.n202 VDD1.n201 9.3005
R838 VDD1.n107 VDD1.n106 9.3005
R839 VDD1.n208 VDD1.n207 9.3005
R840 VDD1.n89 VDD1.n8 8.92171
R841 VDD1.n74 VDD1.n73 8.92171
R842 VDD1.n41 VDD1.n31 8.92171
R843 VDD1.n145 VDD1.n135 8.92171
R844 VDD1.n179 VDD1.n178 8.92171
R845 VDD1.n194 VDD1.n113 8.92171
R846 VDD1.n86 VDD1.n85 8.14595
R847 VDD1.n77 VDD1.n14 8.14595
R848 VDD1.n40 VDD1.n33 8.14595
R849 VDD1.n144 VDD1.n137 8.14595
R850 VDD1.n182 VDD1.n119 8.14595
R851 VDD1.n191 VDD1.n190 8.14595
R852 VDD1.n104 VDD1.n0 7.75445
R853 VDD1.n209 VDD1.n105 7.75445
R854 VDD1.n82 VDD1.n10 7.3702
R855 VDD1.n78 VDD1.n12 7.3702
R856 VDD1.n37 VDD1.n36 7.3702
R857 VDD1.n141 VDD1.n140 7.3702
R858 VDD1.n183 VDD1.n117 7.3702
R859 VDD1.n187 VDD1.n115 7.3702
R860 VDD1.n82 VDD1.n81 6.59444
R861 VDD1.n81 VDD1.n12 6.59444
R862 VDD1.n186 VDD1.n117 6.59444
R863 VDD1.n187 VDD1.n186 6.59444
R864 VDD1.n102 VDD1.n0 6.08283
R865 VDD1.n207 VDD1.n105 6.08283
R866 VDD1.n85 VDD1.n10 5.81868
R867 VDD1.n78 VDD1.n77 5.81868
R868 VDD1.n37 VDD1.n33 5.81868
R869 VDD1.n141 VDD1.n137 5.81868
R870 VDD1.n183 VDD1.n182 5.81868
R871 VDD1.n190 VDD1.n115 5.81868
R872 VDD1.n86 VDD1.n8 5.04292
R873 VDD1.n74 VDD1.n14 5.04292
R874 VDD1.n41 VDD1.n40 5.04292
R875 VDD1.n145 VDD1.n144 5.04292
R876 VDD1.n179 VDD1.n119 5.04292
R877 VDD1.n191 VDD1.n113 5.04292
R878 VDD1.n90 VDD1.n89 4.26717
R879 VDD1.n73 VDD1.n16 4.26717
R880 VDD1.n44 VDD1.n31 4.26717
R881 VDD1.n148 VDD1.n135 4.26717
R882 VDD1.n178 VDD1.n121 4.26717
R883 VDD1.n195 VDD1.n194 4.26717
R884 VDD1.n93 VDD1.n6 3.49141
R885 VDD1.n70 VDD1.n69 3.49141
R886 VDD1.n45 VDD1.n29 3.49141
R887 VDD1.n149 VDD1.n133 3.49141
R888 VDD1.n175 VDD1.n174 3.49141
R889 VDD1.n198 VDD1.n111 3.49141
R890 VDD1.n94 VDD1.n4 2.71565
R891 VDD1.n66 VDD1.n18 2.71565
R892 VDD1.n49 VDD1.n48 2.71565
R893 VDD1.n153 VDD1.n152 2.71565
R894 VDD1.n171 VDD1.n123 2.71565
R895 VDD1.n199 VDD1.n109 2.71565
R896 VDD1.n38 VDD1.n34 2.41282
R897 VDD1.n142 VDD1.n138 2.41282
R898 VDD1.n98 VDD1.n97 1.93989
R899 VDD1.n65 VDD1.n20 1.93989
R900 VDD1.n52 VDD1.n26 1.93989
R901 VDD1.n157 VDD1.n131 1.93989
R902 VDD1.n170 VDD1.n125 1.93989
R903 VDD1.n203 VDD1.n202 1.93989
R904 VDD1.n101 VDD1.n2 1.16414
R905 VDD1.n62 VDD1.n61 1.16414
R906 VDD1.n53 VDD1.n24 1.16414
R907 VDD1.n158 VDD1.n129 1.16414
R908 VDD1.n167 VDD1.n166 1.16414
R909 VDD1.n206 VDD1.n107 1.16414
R910 VDD1.n58 VDD1.n22 0.388379
R911 VDD1.n57 VDD1.n56 0.388379
R912 VDD1.n162 VDD1.n161 0.388379
R913 VDD1.n163 VDD1.n127 0.388379
R914 VDD1.n103 VDD1.n1 0.155672
R915 VDD1.n96 VDD1.n1 0.155672
R916 VDD1.n96 VDD1.n95 0.155672
R917 VDD1.n95 VDD1.n5 0.155672
R918 VDD1.n88 VDD1.n5 0.155672
R919 VDD1.n88 VDD1.n87 0.155672
R920 VDD1.n87 VDD1.n9 0.155672
R921 VDD1.n80 VDD1.n9 0.155672
R922 VDD1.n80 VDD1.n79 0.155672
R923 VDD1.n79 VDD1.n13 0.155672
R924 VDD1.n72 VDD1.n13 0.155672
R925 VDD1.n72 VDD1.n71 0.155672
R926 VDD1.n71 VDD1.n17 0.155672
R927 VDD1.n64 VDD1.n17 0.155672
R928 VDD1.n64 VDD1.n63 0.155672
R929 VDD1.n63 VDD1.n21 0.155672
R930 VDD1.n55 VDD1.n21 0.155672
R931 VDD1.n55 VDD1.n54 0.155672
R932 VDD1.n54 VDD1.n25 0.155672
R933 VDD1.n47 VDD1.n25 0.155672
R934 VDD1.n47 VDD1.n46 0.155672
R935 VDD1.n46 VDD1.n30 0.155672
R936 VDD1.n39 VDD1.n30 0.155672
R937 VDD1.n39 VDD1.n38 0.155672
R938 VDD1.n143 VDD1.n142 0.155672
R939 VDD1.n143 VDD1.n134 0.155672
R940 VDD1.n150 VDD1.n134 0.155672
R941 VDD1.n151 VDD1.n150 0.155672
R942 VDD1.n151 VDD1.n130 0.155672
R943 VDD1.n159 VDD1.n130 0.155672
R944 VDD1.n160 VDD1.n159 0.155672
R945 VDD1.n160 VDD1.n126 0.155672
R946 VDD1.n168 VDD1.n126 0.155672
R947 VDD1.n169 VDD1.n168 0.155672
R948 VDD1.n169 VDD1.n122 0.155672
R949 VDD1.n176 VDD1.n122 0.155672
R950 VDD1.n177 VDD1.n176 0.155672
R951 VDD1.n177 VDD1.n118 0.155672
R952 VDD1.n184 VDD1.n118 0.155672
R953 VDD1.n185 VDD1.n184 0.155672
R954 VDD1.n185 VDD1.n114 0.155672
R955 VDD1.n192 VDD1.n114 0.155672
R956 VDD1.n193 VDD1.n192 0.155672
R957 VDD1.n193 VDD1.n110 0.155672
R958 VDD1.n200 VDD1.n110 0.155672
R959 VDD1.n201 VDD1.n200 0.155672
R960 VDD1.n201 VDD1.n106 0.155672
R961 VDD1.n208 VDD1.n106 0.155672
R962 B.n416 B.n415 585
R963 B.n414 B.n103 585
R964 B.n413 B.n412 585
R965 B.n411 B.n104 585
R966 B.n410 B.n409 585
R967 B.n408 B.n105 585
R968 B.n407 B.n406 585
R969 B.n405 B.n106 585
R970 B.n404 B.n403 585
R971 B.n402 B.n107 585
R972 B.n401 B.n400 585
R973 B.n399 B.n108 585
R974 B.n398 B.n397 585
R975 B.n396 B.n109 585
R976 B.n395 B.n394 585
R977 B.n393 B.n110 585
R978 B.n392 B.n391 585
R979 B.n390 B.n111 585
R980 B.n389 B.n388 585
R981 B.n387 B.n112 585
R982 B.n386 B.n385 585
R983 B.n384 B.n113 585
R984 B.n383 B.n382 585
R985 B.n381 B.n114 585
R986 B.n380 B.n379 585
R987 B.n378 B.n115 585
R988 B.n377 B.n376 585
R989 B.n375 B.n116 585
R990 B.n374 B.n373 585
R991 B.n372 B.n117 585
R992 B.n371 B.n370 585
R993 B.n369 B.n118 585
R994 B.n368 B.n367 585
R995 B.n366 B.n119 585
R996 B.n365 B.n364 585
R997 B.n363 B.n120 585
R998 B.n362 B.n361 585
R999 B.n360 B.n121 585
R1000 B.n359 B.n358 585
R1001 B.n357 B.n122 585
R1002 B.n356 B.n355 585
R1003 B.n354 B.n123 585
R1004 B.n353 B.n352 585
R1005 B.n351 B.n124 585
R1006 B.n350 B.n349 585
R1007 B.n348 B.n125 585
R1008 B.n347 B.n346 585
R1009 B.n345 B.n126 585
R1010 B.n344 B.n343 585
R1011 B.n342 B.n127 585
R1012 B.n341 B.n340 585
R1013 B.n339 B.n128 585
R1014 B.n338 B.n337 585
R1015 B.n336 B.n129 585
R1016 B.n335 B.n334 585
R1017 B.n333 B.n130 585
R1018 B.n332 B.n331 585
R1019 B.n330 B.n131 585
R1020 B.n329 B.n328 585
R1021 B.n327 B.n132 585
R1022 B.n326 B.n325 585
R1023 B.n324 B.n133 585
R1024 B.n323 B.n322 585
R1025 B.n321 B.n134 585
R1026 B.n320 B.n319 585
R1027 B.n315 B.n135 585
R1028 B.n314 B.n313 585
R1029 B.n312 B.n136 585
R1030 B.n311 B.n310 585
R1031 B.n309 B.n137 585
R1032 B.n308 B.n307 585
R1033 B.n306 B.n138 585
R1034 B.n305 B.n304 585
R1035 B.n302 B.n139 585
R1036 B.n301 B.n300 585
R1037 B.n299 B.n142 585
R1038 B.n298 B.n297 585
R1039 B.n296 B.n143 585
R1040 B.n295 B.n294 585
R1041 B.n293 B.n144 585
R1042 B.n292 B.n291 585
R1043 B.n290 B.n145 585
R1044 B.n289 B.n288 585
R1045 B.n287 B.n146 585
R1046 B.n286 B.n285 585
R1047 B.n284 B.n147 585
R1048 B.n283 B.n282 585
R1049 B.n281 B.n148 585
R1050 B.n280 B.n279 585
R1051 B.n278 B.n149 585
R1052 B.n277 B.n276 585
R1053 B.n275 B.n150 585
R1054 B.n274 B.n273 585
R1055 B.n272 B.n151 585
R1056 B.n271 B.n270 585
R1057 B.n269 B.n152 585
R1058 B.n268 B.n267 585
R1059 B.n266 B.n153 585
R1060 B.n265 B.n264 585
R1061 B.n263 B.n154 585
R1062 B.n262 B.n261 585
R1063 B.n260 B.n155 585
R1064 B.n259 B.n258 585
R1065 B.n257 B.n156 585
R1066 B.n256 B.n255 585
R1067 B.n254 B.n157 585
R1068 B.n253 B.n252 585
R1069 B.n251 B.n158 585
R1070 B.n250 B.n249 585
R1071 B.n248 B.n159 585
R1072 B.n247 B.n246 585
R1073 B.n245 B.n160 585
R1074 B.n244 B.n243 585
R1075 B.n242 B.n161 585
R1076 B.n241 B.n240 585
R1077 B.n239 B.n162 585
R1078 B.n238 B.n237 585
R1079 B.n236 B.n163 585
R1080 B.n235 B.n234 585
R1081 B.n233 B.n164 585
R1082 B.n232 B.n231 585
R1083 B.n230 B.n165 585
R1084 B.n229 B.n228 585
R1085 B.n227 B.n166 585
R1086 B.n226 B.n225 585
R1087 B.n224 B.n167 585
R1088 B.n223 B.n222 585
R1089 B.n221 B.n168 585
R1090 B.n220 B.n219 585
R1091 B.n218 B.n169 585
R1092 B.n217 B.n216 585
R1093 B.n215 B.n170 585
R1094 B.n214 B.n213 585
R1095 B.n212 B.n171 585
R1096 B.n211 B.n210 585
R1097 B.n209 B.n172 585
R1098 B.n208 B.n207 585
R1099 B.n417 B.n102 585
R1100 B.n419 B.n418 585
R1101 B.n420 B.n101 585
R1102 B.n422 B.n421 585
R1103 B.n423 B.n100 585
R1104 B.n425 B.n424 585
R1105 B.n426 B.n99 585
R1106 B.n428 B.n427 585
R1107 B.n429 B.n98 585
R1108 B.n431 B.n430 585
R1109 B.n432 B.n97 585
R1110 B.n434 B.n433 585
R1111 B.n435 B.n96 585
R1112 B.n437 B.n436 585
R1113 B.n438 B.n95 585
R1114 B.n440 B.n439 585
R1115 B.n441 B.n94 585
R1116 B.n443 B.n442 585
R1117 B.n444 B.n93 585
R1118 B.n446 B.n445 585
R1119 B.n447 B.n92 585
R1120 B.n449 B.n448 585
R1121 B.n450 B.n91 585
R1122 B.n452 B.n451 585
R1123 B.n453 B.n90 585
R1124 B.n455 B.n454 585
R1125 B.n456 B.n89 585
R1126 B.n458 B.n457 585
R1127 B.n459 B.n88 585
R1128 B.n461 B.n460 585
R1129 B.n462 B.n87 585
R1130 B.n464 B.n463 585
R1131 B.n465 B.n86 585
R1132 B.n467 B.n466 585
R1133 B.n468 B.n85 585
R1134 B.n470 B.n469 585
R1135 B.n471 B.n84 585
R1136 B.n473 B.n472 585
R1137 B.n680 B.n11 585
R1138 B.n679 B.n678 585
R1139 B.n677 B.n12 585
R1140 B.n676 B.n675 585
R1141 B.n674 B.n13 585
R1142 B.n673 B.n672 585
R1143 B.n671 B.n14 585
R1144 B.n670 B.n669 585
R1145 B.n668 B.n15 585
R1146 B.n667 B.n666 585
R1147 B.n665 B.n16 585
R1148 B.n664 B.n663 585
R1149 B.n662 B.n17 585
R1150 B.n661 B.n660 585
R1151 B.n659 B.n18 585
R1152 B.n658 B.n657 585
R1153 B.n656 B.n19 585
R1154 B.n655 B.n654 585
R1155 B.n653 B.n20 585
R1156 B.n652 B.n651 585
R1157 B.n650 B.n21 585
R1158 B.n649 B.n648 585
R1159 B.n647 B.n22 585
R1160 B.n646 B.n645 585
R1161 B.n644 B.n23 585
R1162 B.n643 B.n642 585
R1163 B.n641 B.n24 585
R1164 B.n640 B.n639 585
R1165 B.n638 B.n25 585
R1166 B.n637 B.n636 585
R1167 B.n635 B.n26 585
R1168 B.n634 B.n633 585
R1169 B.n632 B.n27 585
R1170 B.n631 B.n630 585
R1171 B.n629 B.n28 585
R1172 B.n628 B.n627 585
R1173 B.n626 B.n29 585
R1174 B.n625 B.n624 585
R1175 B.n623 B.n30 585
R1176 B.n622 B.n621 585
R1177 B.n620 B.n31 585
R1178 B.n619 B.n618 585
R1179 B.n617 B.n32 585
R1180 B.n616 B.n615 585
R1181 B.n614 B.n33 585
R1182 B.n613 B.n612 585
R1183 B.n611 B.n34 585
R1184 B.n610 B.n609 585
R1185 B.n608 B.n35 585
R1186 B.n607 B.n606 585
R1187 B.n605 B.n36 585
R1188 B.n604 B.n603 585
R1189 B.n602 B.n37 585
R1190 B.n601 B.n600 585
R1191 B.n599 B.n38 585
R1192 B.n598 B.n597 585
R1193 B.n596 B.n39 585
R1194 B.n595 B.n594 585
R1195 B.n593 B.n40 585
R1196 B.n592 B.n591 585
R1197 B.n590 B.n41 585
R1198 B.n589 B.n588 585
R1199 B.n587 B.n42 585
R1200 B.n586 B.n585 585
R1201 B.n583 B.n43 585
R1202 B.n582 B.n581 585
R1203 B.n580 B.n46 585
R1204 B.n579 B.n578 585
R1205 B.n577 B.n47 585
R1206 B.n576 B.n575 585
R1207 B.n574 B.n48 585
R1208 B.n573 B.n572 585
R1209 B.n571 B.n49 585
R1210 B.n569 B.n568 585
R1211 B.n567 B.n52 585
R1212 B.n566 B.n565 585
R1213 B.n564 B.n53 585
R1214 B.n563 B.n562 585
R1215 B.n561 B.n54 585
R1216 B.n560 B.n559 585
R1217 B.n558 B.n55 585
R1218 B.n557 B.n556 585
R1219 B.n555 B.n56 585
R1220 B.n554 B.n553 585
R1221 B.n552 B.n57 585
R1222 B.n551 B.n550 585
R1223 B.n549 B.n58 585
R1224 B.n548 B.n547 585
R1225 B.n546 B.n59 585
R1226 B.n545 B.n544 585
R1227 B.n543 B.n60 585
R1228 B.n542 B.n541 585
R1229 B.n540 B.n61 585
R1230 B.n539 B.n538 585
R1231 B.n537 B.n62 585
R1232 B.n536 B.n535 585
R1233 B.n534 B.n63 585
R1234 B.n533 B.n532 585
R1235 B.n531 B.n64 585
R1236 B.n530 B.n529 585
R1237 B.n528 B.n65 585
R1238 B.n527 B.n526 585
R1239 B.n525 B.n66 585
R1240 B.n524 B.n523 585
R1241 B.n522 B.n67 585
R1242 B.n521 B.n520 585
R1243 B.n519 B.n68 585
R1244 B.n518 B.n517 585
R1245 B.n516 B.n69 585
R1246 B.n515 B.n514 585
R1247 B.n513 B.n70 585
R1248 B.n512 B.n511 585
R1249 B.n510 B.n71 585
R1250 B.n509 B.n508 585
R1251 B.n507 B.n72 585
R1252 B.n506 B.n505 585
R1253 B.n504 B.n73 585
R1254 B.n503 B.n502 585
R1255 B.n501 B.n74 585
R1256 B.n500 B.n499 585
R1257 B.n498 B.n75 585
R1258 B.n497 B.n496 585
R1259 B.n495 B.n76 585
R1260 B.n494 B.n493 585
R1261 B.n492 B.n77 585
R1262 B.n491 B.n490 585
R1263 B.n489 B.n78 585
R1264 B.n488 B.n487 585
R1265 B.n486 B.n79 585
R1266 B.n485 B.n484 585
R1267 B.n483 B.n80 585
R1268 B.n482 B.n481 585
R1269 B.n480 B.n81 585
R1270 B.n479 B.n478 585
R1271 B.n477 B.n82 585
R1272 B.n476 B.n475 585
R1273 B.n474 B.n83 585
R1274 B.n682 B.n681 585
R1275 B.n683 B.n10 585
R1276 B.n685 B.n684 585
R1277 B.n686 B.n9 585
R1278 B.n688 B.n687 585
R1279 B.n689 B.n8 585
R1280 B.n691 B.n690 585
R1281 B.n692 B.n7 585
R1282 B.n694 B.n693 585
R1283 B.n695 B.n6 585
R1284 B.n697 B.n696 585
R1285 B.n698 B.n5 585
R1286 B.n700 B.n699 585
R1287 B.n701 B.n4 585
R1288 B.n703 B.n702 585
R1289 B.n704 B.n3 585
R1290 B.n706 B.n705 585
R1291 B.n707 B.n0 585
R1292 B.n2 B.n1 585
R1293 B.n182 B.n181 585
R1294 B.n184 B.n183 585
R1295 B.n185 B.n180 585
R1296 B.n187 B.n186 585
R1297 B.n188 B.n179 585
R1298 B.n190 B.n189 585
R1299 B.n191 B.n178 585
R1300 B.n193 B.n192 585
R1301 B.n194 B.n177 585
R1302 B.n196 B.n195 585
R1303 B.n197 B.n176 585
R1304 B.n199 B.n198 585
R1305 B.n200 B.n175 585
R1306 B.n202 B.n201 585
R1307 B.n203 B.n174 585
R1308 B.n205 B.n204 585
R1309 B.n206 B.n173 585
R1310 B.n316 B.t4 544.197
R1311 B.n50 B.t11 544.197
R1312 B.n140 B.t1 544.197
R1313 B.n44 B.t8 544.197
R1314 B.n140 B.t0 533.301
R1315 B.n316 B.t3 533.301
R1316 B.n50 B.t9 533.301
R1317 B.n44 B.t6 533.301
R1318 B.n317 B.t5 510.065
R1319 B.n51 B.t10 510.065
R1320 B.n141 B.t2 510.065
R1321 B.n45 B.t7 510.065
R1322 B.n208 B.n173 473.281
R1323 B.n417 B.n416 473.281
R1324 B.n472 B.n83 473.281
R1325 B.n682 B.n11 473.281
R1326 B.n709 B.n708 256.663
R1327 B.n708 B.n707 235.042
R1328 B.n708 B.n2 235.042
R1329 B.n209 B.n208 163.367
R1330 B.n210 B.n209 163.367
R1331 B.n210 B.n171 163.367
R1332 B.n214 B.n171 163.367
R1333 B.n215 B.n214 163.367
R1334 B.n216 B.n215 163.367
R1335 B.n216 B.n169 163.367
R1336 B.n220 B.n169 163.367
R1337 B.n221 B.n220 163.367
R1338 B.n222 B.n221 163.367
R1339 B.n222 B.n167 163.367
R1340 B.n226 B.n167 163.367
R1341 B.n227 B.n226 163.367
R1342 B.n228 B.n227 163.367
R1343 B.n228 B.n165 163.367
R1344 B.n232 B.n165 163.367
R1345 B.n233 B.n232 163.367
R1346 B.n234 B.n233 163.367
R1347 B.n234 B.n163 163.367
R1348 B.n238 B.n163 163.367
R1349 B.n239 B.n238 163.367
R1350 B.n240 B.n239 163.367
R1351 B.n240 B.n161 163.367
R1352 B.n244 B.n161 163.367
R1353 B.n245 B.n244 163.367
R1354 B.n246 B.n245 163.367
R1355 B.n246 B.n159 163.367
R1356 B.n250 B.n159 163.367
R1357 B.n251 B.n250 163.367
R1358 B.n252 B.n251 163.367
R1359 B.n252 B.n157 163.367
R1360 B.n256 B.n157 163.367
R1361 B.n257 B.n256 163.367
R1362 B.n258 B.n257 163.367
R1363 B.n258 B.n155 163.367
R1364 B.n262 B.n155 163.367
R1365 B.n263 B.n262 163.367
R1366 B.n264 B.n263 163.367
R1367 B.n264 B.n153 163.367
R1368 B.n268 B.n153 163.367
R1369 B.n269 B.n268 163.367
R1370 B.n270 B.n269 163.367
R1371 B.n270 B.n151 163.367
R1372 B.n274 B.n151 163.367
R1373 B.n275 B.n274 163.367
R1374 B.n276 B.n275 163.367
R1375 B.n276 B.n149 163.367
R1376 B.n280 B.n149 163.367
R1377 B.n281 B.n280 163.367
R1378 B.n282 B.n281 163.367
R1379 B.n282 B.n147 163.367
R1380 B.n286 B.n147 163.367
R1381 B.n287 B.n286 163.367
R1382 B.n288 B.n287 163.367
R1383 B.n288 B.n145 163.367
R1384 B.n292 B.n145 163.367
R1385 B.n293 B.n292 163.367
R1386 B.n294 B.n293 163.367
R1387 B.n294 B.n143 163.367
R1388 B.n298 B.n143 163.367
R1389 B.n299 B.n298 163.367
R1390 B.n300 B.n299 163.367
R1391 B.n300 B.n139 163.367
R1392 B.n305 B.n139 163.367
R1393 B.n306 B.n305 163.367
R1394 B.n307 B.n306 163.367
R1395 B.n307 B.n137 163.367
R1396 B.n311 B.n137 163.367
R1397 B.n312 B.n311 163.367
R1398 B.n313 B.n312 163.367
R1399 B.n313 B.n135 163.367
R1400 B.n320 B.n135 163.367
R1401 B.n321 B.n320 163.367
R1402 B.n322 B.n321 163.367
R1403 B.n322 B.n133 163.367
R1404 B.n326 B.n133 163.367
R1405 B.n327 B.n326 163.367
R1406 B.n328 B.n327 163.367
R1407 B.n328 B.n131 163.367
R1408 B.n332 B.n131 163.367
R1409 B.n333 B.n332 163.367
R1410 B.n334 B.n333 163.367
R1411 B.n334 B.n129 163.367
R1412 B.n338 B.n129 163.367
R1413 B.n339 B.n338 163.367
R1414 B.n340 B.n339 163.367
R1415 B.n340 B.n127 163.367
R1416 B.n344 B.n127 163.367
R1417 B.n345 B.n344 163.367
R1418 B.n346 B.n345 163.367
R1419 B.n346 B.n125 163.367
R1420 B.n350 B.n125 163.367
R1421 B.n351 B.n350 163.367
R1422 B.n352 B.n351 163.367
R1423 B.n352 B.n123 163.367
R1424 B.n356 B.n123 163.367
R1425 B.n357 B.n356 163.367
R1426 B.n358 B.n357 163.367
R1427 B.n358 B.n121 163.367
R1428 B.n362 B.n121 163.367
R1429 B.n363 B.n362 163.367
R1430 B.n364 B.n363 163.367
R1431 B.n364 B.n119 163.367
R1432 B.n368 B.n119 163.367
R1433 B.n369 B.n368 163.367
R1434 B.n370 B.n369 163.367
R1435 B.n370 B.n117 163.367
R1436 B.n374 B.n117 163.367
R1437 B.n375 B.n374 163.367
R1438 B.n376 B.n375 163.367
R1439 B.n376 B.n115 163.367
R1440 B.n380 B.n115 163.367
R1441 B.n381 B.n380 163.367
R1442 B.n382 B.n381 163.367
R1443 B.n382 B.n113 163.367
R1444 B.n386 B.n113 163.367
R1445 B.n387 B.n386 163.367
R1446 B.n388 B.n387 163.367
R1447 B.n388 B.n111 163.367
R1448 B.n392 B.n111 163.367
R1449 B.n393 B.n392 163.367
R1450 B.n394 B.n393 163.367
R1451 B.n394 B.n109 163.367
R1452 B.n398 B.n109 163.367
R1453 B.n399 B.n398 163.367
R1454 B.n400 B.n399 163.367
R1455 B.n400 B.n107 163.367
R1456 B.n404 B.n107 163.367
R1457 B.n405 B.n404 163.367
R1458 B.n406 B.n405 163.367
R1459 B.n406 B.n105 163.367
R1460 B.n410 B.n105 163.367
R1461 B.n411 B.n410 163.367
R1462 B.n412 B.n411 163.367
R1463 B.n412 B.n103 163.367
R1464 B.n416 B.n103 163.367
R1465 B.n472 B.n471 163.367
R1466 B.n471 B.n470 163.367
R1467 B.n470 B.n85 163.367
R1468 B.n466 B.n85 163.367
R1469 B.n466 B.n465 163.367
R1470 B.n465 B.n464 163.367
R1471 B.n464 B.n87 163.367
R1472 B.n460 B.n87 163.367
R1473 B.n460 B.n459 163.367
R1474 B.n459 B.n458 163.367
R1475 B.n458 B.n89 163.367
R1476 B.n454 B.n89 163.367
R1477 B.n454 B.n453 163.367
R1478 B.n453 B.n452 163.367
R1479 B.n452 B.n91 163.367
R1480 B.n448 B.n91 163.367
R1481 B.n448 B.n447 163.367
R1482 B.n447 B.n446 163.367
R1483 B.n446 B.n93 163.367
R1484 B.n442 B.n93 163.367
R1485 B.n442 B.n441 163.367
R1486 B.n441 B.n440 163.367
R1487 B.n440 B.n95 163.367
R1488 B.n436 B.n95 163.367
R1489 B.n436 B.n435 163.367
R1490 B.n435 B.n434 163.367
R1491 B.n434 B.n97 163.367
R1492 B.n430 B.n97 163.367
R1493 B.n430 B.n429 163.367
R1494 B.n429 B.n428 163.367
R1495 B.n428 B.n99 163.367
R1496 B.n424 B.n99 163.367
R1497 B.n424 B.n423 163.367
R1498 B.n423 B.n422 163.367
R1499 B.n422 B.n101 163.367
R1500 B.n418 B.n101 163.367
R1501 B.n418 B.n417 163.367
R1502 B.n678 B.n11 163.367
R1503 B.n678 B.n677 163.367
R1504 B.n677 B.n676 163.367
R1505 B.n676 B.n13 163.367
R1506 B.n672 B.n13 163.367
R1507 B.n672 B.n671 163.367
R1508 B.n671 B.n670 163.367
R1509 B.n670 B.n15 163.367
R1510 B.n666 B.n15 163.367
R1511 B.n666 B.n665 163.367
R1512 B.n665 B.n664 163.367
R1513 B.n664 B.n17 163.367
R1514 B.n660 B.n17 163.367
R1515 B.n660 B.n659 163.367
R1516 B.n659 B.n658 163.367
R1517 B.n658 B.n19 163.367
R1518 B.n654 B.n19 163.367
R1519 B.n654 B.n653 163.367
R1520 B.n653 B.n652 163.367
R1521 B.n652 B.n21 163.367
R1522 B.n648 B.n21 163.367
R1523 B.n648 B.n647 163.367
R1524 B.n647 B.n646 163.367
R1525 B.n646 B.n23 163.367
R1526 B.n642 B.n23 163.367
R1527 B.n642 B.n641 163.367
R1528 B.n641 B.n640 163.367
R1529 B.n640 B.n25 163.367
R1530 B.n636 B.n25 163.367
R1531 B.n636 B.n635 163.367
R1532 B.n635 B.n634 163.367
R1533 B.n634 B.n27 163.367
R1534 B.n630 B.n27 163.367
R1535 B.n630 B.n629 163.367
R1536 B.n629 B.n628 163.367
R1537 B.n628 B.n29 163.367
R1538 B.n624 B.n29 163.367
R1539 B.n624 B.n623 163.367
R1540 B.n623 B.n622 163.367
R1541 B.n622 B.n31 163.367
R1542 B.n618 B.n31 163.367
R1543 B.n618 B.n617 163.367
R1544 B.n617 B.n616 163.367
R1545 B.n616 B.n33 163.367
R1546 B.n612 B.n33 163.367
R1547 B.n612 B.n611 163.367
R1548 B.n611 B.n610 163.367
R1549 B.n610 B.n35 163.367
R1550 B.n606 B.n35 163.367
R1551 B.n606 B.n605 163.367
R1552 B.n605 B.n604 163.367
R1553 B.n604 B.n37 163.367
R1554 B.n600 B.n37 163.367
R1555 B.n600 B.n599 163.367
R1556 B.n599 B.n598 163.367
R1557 B.n598 B.n39 163.367
R1558 B.n594 B.n39 163.367
R1559 B.n594 B.n593 163.367
R1560 B.n593 B.n592 163.367
R1561 B.n592 B.n41 163.367
R1562 B.n588 B.n41 163.367
R1563 B.n588 B.n587 163.367
R1564 B.n587 B.n586 163.367
R1565 B.n586 B.n43 163.367
R1566 B.n581 B.n43 163.367
R1567 B.n581 B.n580 163.367
R1568 B.n580 B.n579 163.367
R1569 B.n579 B.n47 163.367
R1570 B.n575 B.n47 163.367
R1571 B.n575 B.n574 163.367
R1572 B.n574 B.n573 163.367
R1573 B.n573 B.n49 163.367
R1574 B.n568 B.n49 163.367
R1575 B.n568 B.n567 163.367
R1576 B.n567 B.n566 163.367
R1577 B.n566 B.n53 163.367
R1578 B.n562 B.n53 163.367
R1579 B.n562 B.n561 163.367
R1580 B.n561 B.n560 163.367
R1581 B.n560 B.n55 163.367
R1582 B.n556 B.n55 163.367
R1583 B.n556 B.n555 163.367
R1584 B.n555 B.n554 163.367
R1585 B.n554 B.n57 163.367
R1586 B.n550 B.n57 163.367
R1587 B.n550 B.n549 163.367
R1588 B.n549 B.n548 163.367
R1589 B.n548 B.n59 163.367
R1590 B.n544 B.n59 163.367
R1591 B.n544 B.n543 163.367
R1592 B.n543 B.n542 163.367
R1593 B.n542 B.n61 163.367
R1594 B.n538 B.n61 163.367
R1595 B.n538 B.n537 163.367
R1596 B.n537 B.n536 163.367
R1597 B.n536 B.n63 163.367
R1598 B.n532 B.n63 163.367
R1599 B.n532 B.n531 163.367
R1600 B.n531 B.n530 163.367
R1601 B.n530 B.n65 163.367
R1602 B.n526 B.n65 163.367
R1603 B.n526 B.n525 163.367
R1604 B.n525 B.n524 163.367
R1605 B.n524 B.n67 163.367
R1606 B.n520 B.n67 163.367
R1607 B.n520 B.n519 163.367
R1608 B.n519 B.n518 163.367
R1609 B.n518 B.n69 163.367
R1610 B.n514 B.n69 163.367
R1611 B.n514 B.n513 163.367
R1612 B.n513 B.n512 163.367
R1613 B.n512 B.n71 163.367
R1614 B.n508 B.n71 163.367
R1615 B.n508 B.n507 163.367
R1616 B.n507 B.n506 163.367
R1617 B.n506 B.n73 163.367
R1618 B.n502 B.n73 163.367
R1619 B.n502 B.n501 163.367
R1620 B.n501 B.n500 163.367
R1621 B.n500 B.n75 163.367
R1622 B.n496 B.n75 163.367
R1623 B.n496 B.n495 163.367
R1624 B.n495 B.n494 163.367
R1625 B.n494 B.n77 163.367
R1626 B.n490 B.n77 163.367
R1627 B.n490 B.n489 163.367
R1628 B.n489 B.n488 163.367
R1629 B.n488 B.n79 163.367
R1630 B.n484 B.n79 163.367
R1631 B.n484 B.n483 163.367
R1632 B.n483 B.n482 163.367
R1633 B.n482 B.n81 163.367
R1634 B.n478 B.n81 163.367
R1635 B.n478 B.n477 163.367
R1636 B.n477 B.n476 163.367
R1637 B.n476 B.n83 163.367
R1638 B.n683 B.n682 163.367
R1639 B.n684 B.n683 163.367
R1640 B.n684 B.n9 163.367
R1641 B.n688 B.n9 163.367
R1642 B.n689 B.n688 163.367
R1643 B.n690 B.n689 163.367
R1644 B.n690 B.n7 163.367
R1645 B.n694 B.n7 163.367
R1646 B.n695 B.n694 163.367
R1647 B.n696 B.n695 163.367
R1648 B.n696 B.n5 163.367
R1649 B.n700 B.n5 163.367
R1650 B.n701 B.n700 163.367
R1651 B.n702 B.n701 163.367
R1652 B.n702 B.n3 163.367
R1653 B.n706 B.n3 163.367
R1654 B.n707 B.n706 163.367
R1655 B.n181 B.n2 163.367
R1656 B.n184 B.n181 163.367
R1657 B.n185 B.n184 163.367
R1658 B.n186 B.n185 163.367
R1659 B.n186 B.n179 163.367
R1660 B.n190 B.n179 163.367
R1661 B.n191 B.n190 163.367
R1662 B.n192 B.n191 163.367
R1663 B.n192 B.n177 163.367
R1664 B.n196 B.n177 163.367
R1665 B.n197 B.n196 163.367
R1666 B.n198 B.n197 163.367
R1667 B.n198 B.n175 163.367
R1668 B.n202 B.n175 163.367
R1669 B.n203 B.n202 163.367
R1670 B.n204 B.n203 163.367
R1671 B.n204 B.n173 163.367
R1672 B.n303 B.n141 59.5399
R1673 B.n318 B.n317 59.5399
R1674 B.n570 B.n51 59.5399
R1675 B.n584 B.n45 59.5399
R1676 B.n141 B.n140 34.1338
R1677 B.n317 B.n316 34.1338
R1678 B.n51 B.n50 34.1338
R1679 B.n45 B.n44 34.1338
R1680 B.n681 B.n680 30.7517
R1681 B.n474 B.n473 30.7517
R1682 B.n415 B.n102 30.7517
R1683 B.n207 B.n206 30.7517
R1684 B B.n709 18.0485
R1685 B.n681 B.n10 10.6151
R1686 B.n685 B.n10 10.6151
R1687 B.n686 B.n685 10.6151
R1688 B.n687 B.n686 10.6151
R1689 B.n687 B.n8 10.6151
R1690 B.n691 B.n8 10.6151
R1691 B.n692 B.n691 10.6151
R1692 B.n693 B.n692 10.6151
R1693 B.n693 B.n6 10.6151
R1694 B.n697 B.n6 10.6151
R1695 B.n698 B.n697 10.6151
R1696 B.n699 B.n698 10.6151
R1697 B.n699 B.n4 10.6151
R1698 B.n703 B.n4 10.6151
R1699 B.n704 B.n703 10.6151
R1700 B.n705 B.n704 10.6151
R1701 B.n705 B.n0 10.6151
R1702 B.n680 B.n679 10.6151
R1703 B.n679 B.n12 10.6151
R1704 B.n675 B.n12 10.6151
R1705 B.n675 B.n674 10.6151
R1706 B.n674 B.n673 10.6151
R1707 B.n673 B.n14 10.6151
R1708 B.n669 B.n14 10.6151
R1709 B.n669 B.n668 10.6151
R1710 B.n668 B.n667 10.6151
R1711 B.n667 B.n16 10.6151
R1712 B.n663 B.n16 10.6151
R1713 B.n663 B.n662 10.6151
R1714 B.n662 B.n661 10.6151
R1715 B.n661 B.n18 10.6151
R1716 B.n657 B.n18 10.6151
R1717 B.n657 B.n656 10.6151
R1718 B.n656 B.n655 10.6151
R1719 B.n655 B.n20 10.6151
R1720 B.n651 B.n20 10.6151
R1721 B.n651 B.n650 10.6151
R1722 B.n650 B.n649 10.6151
R1723 B.n649 B.n22 10.6151
R1724 B.n645 B.n22 10.6151
R1725 B.n645 B.n644 10.6151
R1726 B.n644 B.n643 10.6151
R1727 B.n643 B.n24 10.6151
R1728 B.n639 B.n24 10.6151
R1729 B.n639 B.n638 10.6151
R1730 B.n638 B.n637 10.6151
R1731 B.n637 B.n26 10.6151
R1732 B.n633 B.n26 10.6151
R1733 B.n633 B.n632 10.6151
R1734 B.n632 B.n631 10.6151
R1735 B.n631 B.n28 10.6151
R1736 B.n627 B.n28 10.6151
R1737 B.n627 B.n626 10.6151
R1738 B.n626 B.n625 10.6151
R1739 B.n625 B.n30 10.6151
R1740 B.n621 B.n30 10.6151
R1741 B.n621 B.n620 10.6151
R1742 B.n620 B.n619 10.6151
R1743 B.n619 B.n32 10.6151
R1744 B.n615 B.n32 10.6151
R1745 B.n615 B.n614 10.6151
R1746 B.n614 B.n613 10.6151
R1747 B.n613 B.n34 10.6151
R1748 B.n609 B.n34 10.6151
R1749 B.n609 B.n608 10.6151
R1750 B.n608 B.n607 10.6151
R1751 B.n607 B.n36 10.6151
R1752 B.n603 B.n36 10.6151
R1753 B.n603 B.n602 10.6151
R1754 B.n602 B.n601 10.6151
R1755 B.n601 B.n38 10.6151
R1756 B.n597 B.n38 10.6151
R1757 B.n597 B.n596 10.6151
R1758 B.n596 B.n595 10.6151
R1759 B.n595 B.n40 10.6151
R1760 B.n591 B.n40 10.6151
R1761 B.n591 B.n590 10.6151
R1762 B.n590 B.n589 10.6151
R1763 B.n589 B.n42 10.6151
R1764 B.n585 B.n42 10.6151
R1765 B.n583 B.n582 10.6151
R1766 B.n582 B.n46 10.6151
R1767 B.n578 B.n46 10.6151
R1768 B.n578 B.n577 10.6151
R1769 B.n577 B.n576 10.6151
R1770 B.n576 B.n48 10.6151
R1771 B.n572 B.n48 10.6151
R1772 B.n572 B.n571 10.6151
R1773 B.n569 B.n52 10.6151
R1774 B.n565 B.n52 10.6151
R1775 B.n565 B.n564 10.6151
R1776 B.n564 B.n563 10.6151
R1777 B.n563 B.n54 10.6151
R1778 B.n559 B.n54 10.6151
R1779 B.n559 B.n558 10.6151
R1780 B.n558 B.n557 10.6151
R1781 B.n557 B.n56 10.6151
R1782 B.n553 B.n56 10.6151
R1783 B.n553 B.n552 10.6151
R1784 B.n552 B.n551 10.6151
R1785 B.n551 B.n58 10.6151
R1786 B.n547 B.n58 10.6151
R1787 B.n547 B.n546 10.6151
R1788 B.n546 B.n545 10.6151
R1789 B.n545 B.n60 10.6151
R1790 B.n541 B.n60 10.6151
R1791 B.n541 B.n540 10.6151
R1792 B.n540 B.n539 10.6151
R1793 B.n539 B.n62 10.6151
R1794 B.n535 B.n62 10.6151
R1795 B.n535 B.n534 10.6151
R1796 B.n534 B.n533 10.6151
R1797 B.n533 B.n64 10.6151
R1798 B.n529 B.n64 10.6151
R1799 B.n529 B.n528 10.6151
R1800 B.n528 B.n527 10.6151
R1801 B.n527 B.n66 10.6151
R1802 B.n523 B.n66 10.6151
R1803 B.n523 B.n522 10.6151
R1804 B.n522 B.n521 10.6151
R1805 B.n521 B.n68 10.6151
R1806 B.n517 B.n68 10.6151
R1807 B.n517 B.n516 10.6151
R1808 B.n516 B.n515 10.6151
R1809 B.n515 B.n70 10.6151
R1810 B.n511 B.n70 10.6151
R1811 B.n511 B.n510 10.6151
R1812 B.n510 B.n509 10.6151
R1813 B.n509 B.n72 10.6151
R1814 B.n505 B.n72 10.6151
R1815 B.n505 B.n504 10.6151
R1816 B.n504 B.n503 10.6151
R1817 B.n503 B.n74 10.6151
R1818 B.n499 B.n74 10.6151
R1819 B.n499 B.n498 10.6151
R1820 B.n498 B.n497 10.6151
R1821 B.n497 B.n76 10.6151
R1822 B.n493 B.n76 10.6151
R1823 B.n493 B.n492 10.6151
R1824 B.n492 B.n491 10.6151
R1825 B.n491 B.n78 10.6151
R1826 B.n487 B.n78 10.6151
R1827 B.n487 B.n486 10.6151
R1828 B.n486 B.n485 10.6151
R1829 B.n485 B.n80 10.6151
R1830 B.n481 B.n80 10.6151
R1831 B.n481 B.n480 10.6151
R1832 B.n480 B.n479 10.6151
R1833 B.n479 B.n82 10.6151
R1834 B.n475 B.n82 10.6151
R1835 B.n475 B.n474 10.6151
R1836 B.n473 B.n84 10.6151
R1837 B.n469 B.n84 10.6151
R1838 B.n469 B.n468 10.6151
R1839 B.n468 B.n467 10.6151
R1840 B.n467 B.n86 10.6151
R1841 B.n463 B.n86 10.6151
R1842 B.n463 B.n462 10.6151
R1843 B.n462 B.n461 10.6151
R1844 B.n461 B.n88 10.6151
R1845 B.n457 B.n88 10.6151
R1846 B.n457 B.n456 10.6151
R1847 B.n456 B.n455 10.6151
R1848 B.n455 B.n90 10.6151
R1849 B.n451 B.n90 10.6151
R1850 B.n451 B.n450 10.6151
R1851 B.n450 B.n449 10.6151
R1852 B.n449 B.n92 10.6151
R1853 B.n445 B.n92 10.6151
R1854 B.n445 B.n444 10.6151
R1855 B.n444 B.n443 10.6151
R1856 B.n443 B.n94 10.6151
R1857 B.n439 B.n94 10.6151
R1858 B.n439 B.n438 10.6151
R1859 B.n438 B.n437 10.6151
R1860 B.n437 B.n96 10.6151
R1861 B.n433 B.n96 10.6151
R1862 B.n433 B.n432 10.6151
R1863 B.n432 B.n431 10.6151
R1864 B.n431 B.n98 10.6151
R1865 B.n427 B.n98 10.6151
R1866 B.n427 B.n426 10.6151
R1867 B.n426 B.n425 10.6151
R1868 B.n425 B.n100 10.6151
R1869 B.n421 B.n100 10.6151
R1870 B.n421 B.n420 10.6151
R1871 B.n420 B.n419 10.6151
R1872 B.n419 B.n102 10.6151
R1873 B.n182 B.n1 10.6151
R1874 B.n183 B.n182 10.6151
R1875 B.n183 B.n180 10.6151
R1876 B.n187 B.n180 10.6151
R1877 B.n188 B.n187 10.6151
R1878 B.n189 B.n188 10.6151
R1879 B.n189 B.n178 10.6151
R1880 B.n193 B.n178 10.6151
R1881 B.n194 B.n193 10.6151
R1882 B.n195 B.n194 10.6151
R1883 B.n195 B.n176 10.6151
R1884 B.n199 B.n176 10.6151
R1885 B.n200 B.n199 10.6151
R1886 B.n201 B.n200 10.6151
R1887 B.n201 B.n174 10.6151
R1888 B.n205 B.n174 10.6151
R1889 B.n206 B.n205 10.6151
R1890 B.n207 B.n172 10.6151
R1891 B.n211 B.n172 10.6151
R1892 B.n212 B.n211 10.6151
R1893 B.n213 B.n212 10.6151
R1894 B.n213 B.n170 10.6151
R1895 B.n217 B.n170 10.6151
R1896 B.n218 B.n217 10.6151
R1897 B.n219 B.n218 10.6151
R1898 B.n219 B.n168 10.6151
R1899 B.n223 B.n168 10.6151
R1900 B.n224 B.n223 10.6151
R1901 B.n225 B.n224 10.6151
R1902 B.n225 B.n166 10.6151
R1903 B.n229 B.n166 10.6151
R1904 B.n230 B.n229 10.6151
R1905 B.n231 B.n230 10.6151
R1906 B.n231 B.n164 10.6151
R1907 B.n235 B.n164 10.6151
R1908 B.n236 B.n235 10.6151
R1909 B.n237 B.n236 10.6151
R1910 B.n237 B.n162 10.6151
R1911 B.n241 B.n162 10.6151
R1912 B.n242 B.n241 10.6151
R1913 B.n243 B.n242 10.6151
R1914 B.n243 B.n160 10.6151
R1915 B.n247 B.n160 10.6151
R1916 B.n248 B.n247 10.6151
R1917 B.n249 B.n248 10.6151
R1918 B.n249 B.n158 10.6151
R1919 B.n253 B.n158 10.6151
R1920 B.n254 B.n253 10.6151
R1921 B.n255 B.n254 10.6151
R1922 B.n255 B.n156 10.6151
R1923 B.n259 B.n156 10.6151
R1924 B.n260 B.n259 10.6151
R1925 B.n261 B.n260 10.6151
R1926 B.n261 B.n154 10.6151
R1927 B.n265 B.n154 10.6151
R1928 B.n266 B.n265 10.6151
R1929 B.n267 B.n266 10.6151
R1930 B.n267 B.n152 10.6151
R1931 B.n271 B.n152 10.6151
R1932 B.n272 B.n271 10.6151
R1933 B.n273 B.n272 10.6151
R1934 B.n273 B.n150 10.6151
R1935 B.n277 B.n150 10.6151
R1936 B.n278 B.n277 10.6151
R1937 B.n279 B.n278 10.6151
R1938 B.n279 B.n148 10.6151
R1939 B.n283 B.n148 10.6151
R1940 B.n284 B.n283 10.6151
R1941 B.n285 B.n284 10.6151
R1942 B.n285 B.n146 10.6151
R1943 B.n289 B.n146 10.6151
R1944 B.n290 B.n289 10.6151
R1945 B.n291 B.n290 10.6151
R1946 B.n291 B.n144 10.6151
R1947 B.n295 B.n144 10.6151
R1948 B.n296 B.n295 10.6151
R1949 B.n297 B.n296 10.6151
R1950 B.n297 B.n142 10.6151
R1951 B.n301 B.n142 10.6151
R1952 B.n302 B.n301 10.6151
R1953 B.n304 B.n138 10.6151
R1954 B.n308 B.n138 10.6151
R1955 B.n309 B.n308 10.6151
R1956 B.n310 B.n309 10.6151
R1957 B.n310 B.n136 10.6151
R1958 B.n314 B.n136 10.6151
R1959 B.n315 B.n314 10.6151
R1960 B.n319 B.n315 10.6151
R1961 B.n323 B.n134 10.6151
R1962 B.n324 B.n323 10.6151
R1963 B.n325 B.n324 10.6151
R1964 B.n325 B.n132 10.6151
R1965 B.n329 B.n132 10.6151
R1966 B.n330 B.n329 10.6151
R1967 B.n331 B.n330 10.6151
R1968 B.n331 B.n130 10.6151
R1969 B.n335 B.n130 10.6151
R1970 B.n336 B.n335 10.6151
R1971 B.n337 B.n336 10.6151
R1972 B.n337 B.n128 10.6151
R1973 B.n341 B.n128 10.6151
R1974 B.n342 B.n341 10.6151
R1975 B.n343 B.n342 10.6151
R1976 B.n343 B.n126 10.6151
R1977 B.n347 B.n126 10.6151
R1978 B.n348 B.n347 10.6151
R1979 B.n349 B.n348 10.6151
R1980 B.n349 B.n124 10.6151
R1981 B.n353 B.n124 10.6151
R1982 B.n354 B.n353 10.6151
R1983 B.n355 B.n354 10.6151
R1984 B.n355 B.n122 10.6151
R1985 B.n359 B.n122 10.6151
R1986 B.n360 B.n359 10.6151
R1987 B.n361 B.n360 10.6151
R1988 B.n361 B.n120 10.6151
R1989 B.n365 B.n120 10.6151
R1990 B.n366 B.n365 10.6151
R1991 B.n367 B.n366 10.6151
R1992 B.n367 B.n118 10.6151
R1993 B.n371 B.n118 10.6151
R1994 B.n372 B.n371 10.6151
R1995 B.n373 B.n372 10.6151
R1996 B.n373 B.n116 10.6151
R1997 B.n377 B.n116 10.6151
R1998 B.n378 B.n377 10.6151
R1999 B.n379 B.n378 10.6151
R2000 B.n379 B.n114 10.6151
R2001 B.n383 B.n114 10.6151
R2002 B.n384 B.n383 10.6151
R2003 B.n385 B.n384 10.6151
R2004 B.n385 B.n112 10.6151
R2005 B.n389 B.n112 10.6151
R2006 B.n390 B.n389 10.6151
R2007 B.n391 B.n390 10.6151
R2008 B.n391 B.n110 10.6151
R2009 B.n395 B.n110 10.6151
R2010 B.n396 B.n395 10.6151
R2011 B.n397 B.n396 10.6151
R2012 B.n397 B.n108 10.6151
R2013 B.n401 B.n108 10.6151
R2014 B.n402 B.n401 10.6151
R2015 B.n403 B.n402 10.6151
R2016 B.n403 B.n106 10.6151
R2017 B.n407 B.n106 10.6151
R2018 B.n408 B.n407 10.6151
R2019 B.n409 B.n408 10.6151
R2020 B.n409 B.n104 10.6151
R2021 B.n413 B.n104 10.6151
R2022 B.n414 B.n413 10.6151
R2023 B.n415 B.n414 10.6151
R2024 B.n709 B.n0 8.11757
R2025 B.n709 B.n1 8.11757
R2026 B.n584 B.n583 6.5566
R2027 B.n571 B.n570 6.5566
R2028 B.n304 B.n303 6.5566
R2029 B.n319 B.n318 6.5566
R2030 B.n585 B.n584 4.05904
R2031 B.n570 B.n569 4.05904
R2032 B.n303 B.n302 4.05904
R2033 B.n318 B.n134 4.05904
R2034 VN VN.t0 483.873
R2035 VN VN.t1 436.519
R2036 VDD2.n206 VDD2.n205 585
R2037 VDD2.n204 VDD2.n203 585
R2038 VDD2.n109 VDD2.n108 585
R2039 VDD2.n198 VDD2.n197 585
R2040 VDD2.n196 VDD2.n195 585
R2041 VDD2.n113 VDD2.n112 585
R2042 VDD2.n190 VDD2.n189 585
R2043 VDD2.n188 VDD2.n187 585
R2044 VDD2.n117 VDD2.n116 585
R2045 VDD2.n182 VDD2.n181 585
R2046 VDD2.n180 VDD2.n179 585
R2047 VDD2.n121 VDD2.n120 585
R2048 VDD2.n174 VDD2.n173 585
R2049 VDD2.n172 VDD2.n171 585
R2050 VDD2.n125 VDD2.n124 585
R2051 VDD2.n166 VDD2.n165 585
R2052 VDD2.n164 VDD2.n163 585
R2053 VDD2.n162 VDD2.n128 585
R2054 VDD2.n132 VDD2.n129 585
R2055 VDD2.n157 VDD2.n156 585
R2056 VDD2.n155 VDD2.n154 585
R2057 VDD2.n134 VDD2.n133 585
R2058 VDD2.n149 VDD2.n148 585
R2059 VDD2.n147 VDD2.n146 585
R2060 VDD2.n138 VDD2.n137 585
R2061 VDD2.n141 VDD2.n140 585
R2062 VDD2.n35 VDD2.n34 585
R2063 VDD2.n32 VDD2.n31 585
R2064 VDD2.n41 VDD2.n40 585
R2065 VDD2.n43 VDD2.n42 585
R2066 VDD2.n28 VDD2.n27 585
R2067 VDD2.n49 VDD2.n48 585
R2068 VDD2.n52 VDD2.n51 585
R2069 VDD2.n50 VDD2.n24 585
R2070 VDD2.n57 VDD2.n23 585
R2071 VDD2.n59 VDD2.n58 585
R2072 VDD2.n61 VDD2.n60 585
R2073 VDD2.n20 VDD2.n19 585
R2074 VDD2.n67 VDD2.n66 585
R2075 VDD2.n69 VDD2.n68 585
R2076 VDD2.n16 VDD2.n15 585
R2077 VDD2.n75 VDD2.n74 585
R2078 VDD2.n77 VDD2.n76 585
R2079 VDD2.n12 VDD2.n11 585
R2080 VDD2.n83 VDD2.n82 585
R2081 VDD2.n85 VDD2.n84 585
R2082 VDD2.n8 VDD2.n7 585
R2083 VDD2.n91 VDD2.n90 585
R2084 VDD2.n93 VDD2.n92 585
R2085 VDD2.n4 VDD2.n3 585
R2086 VDD2.n99 VDD2.n98 585
R2087 VDD2.n101 VDD2.n100 585
R2088 VDD2.n205 VDD2.n105 498.474
R2089 VDD2.n100 VDD2.n0 498.474
R2090 VDD2.t1 VDD2.n139 329.036
R2091 VDD2.t0 VDD2.n33 329.036
R2092 VDD2.n205 VDD2.n204 171.744
R2093 VDD2.n204 VDD2.n108 171.744
R2094 VDD2.n197 VDD2.n108 171.744
R2095 VDD2.n197 VDD2.n196 171.744
R2096 VDD2.n196 VDD2.n112 171.744
R2097 VDD2.n189 VDD2.n112 171.744
R2098 VDD2.n189 VDD2.n188 171.744
R2099 VDD2.n188 VDD2.n116 171.744
R2100 VDD2.n181 VDD2.n116 171.744
R2101 VDD2.n181 VDD2.n180 171.744
R2102 VDD2.n180 VDD2.n120 171.744
R2103 VDD2.n173 VDD2.n120 171.744
R2104 VDD2.n173 VDD2.n172 171.744
R2105 VDD2.n172 VDD2.n124 171.744
R2106 VDD2.n165 VDD2.n124 171.744
R2107 VDD2.n165 VDD2.n164 171.744
R2108 VDD2.n164 VDD2.n128 171.744
R2109 VDD2.n132 VDD2.n128 171.744
R2110 VDD2.n156 VDD2.n132 171.744
R2111 VDD2.n156 VDD2.n155 171.744
R2112 VDD2.n155 VDD2.n133 171.744
R2113 VDD2.n148 VDD2.n133 171.744
R2114 VDD2.n148 VDD2.n147 171.744
R2115 VDD2.n147 VDD2.n137 171.744
R2116 VDD2.n140 VDD2.n137 171.744
R2117 VDD2.n34 VDD2.n31 171.744
R2118 VDD2.n41 VDD2.n31 171.744
R2119 VDD2.n42 VDD2.n41 171.744
R2120 VDD2.n42 VDD2.n27 171.744
R2121 VDD2.n49 VDD2.n27 171.744
R2122 VDD2.n51 VDD2.n49 171.744
R2123 VDD2.n51 VDD2.n50 171.744
R2124 VDD2.n50 VDD2.n23 171.744
R2125 VDD2.n59 VDD2.n23 171.744
R2126 VDD2.n60 VDD2.n59 171.744
R2127 VDD2.n60 VDD2.n19 171.744
R2128 VDD2.n67 VDD2.n19 171.744
R2129 VDD2.n68 VDD2.n67 171.744
R2130 VDD2.n68 VDD2.n15 171.744
R2131 VDD2.n75 VDD2.n15 171.744
R2132 VDD2.n76 VDD2.n75 171.744
R2133 VDD2.n76 VDD2.n11 171.744
R2134 VDD2.n83 VDD2.n11 171.744
R2135 VDD2.n84 VDD2.n83 171.744
R2136 VDD2.n84 VDD2.n7 171.744
R2137 VDD2.n91 VDD2.n7 171.744
R2138 VDD2.n92 VDD2.n91 171.744
R2139 VDD2.n92 VDD2.n3 171.744
R2140 VDD2.n99 VDD2.n3 171.744
R2141 VDD2.n100 VDD2.n99 171.744
R2142 VDD2.n210 VDD2.n104 95.2516
R2143 VDD2.n140 VDD2.t1 85.8723
R2144 VDD2.n34 VDD2.t0 85.8723
R2145 VDD2.n210 VDD2.n209 51.7732
R2146 VDD2.n163 VDD2.n162 13.1884
R2147 VDD2.n58 VDD2.n57 13.1884
R2148 VDD2.n207 VDD2.n206 12.8005
R2149 VDD2.n166 VDD2.n127 12.8005
R2150 VDD2.n161 VDD2.n129 12.8005
R2151 VDD2.n56 VDD2.n24 12.8005
R2152 VDD2.n61 VDD2.n22 12.8005
R2153 VDD2.n102 VDD2.n101 12.8005
R2154 VDD2.n203 VDD2.n107 12.0247
R2155 VDD2.n167 VDD2.n125 12.0247
R2156 VDD2.n158 VDD2.n157 12.0247
R2157 VDD2.n53 VDD2.n52 12.0247
R2158 VDD2.n62 VDD2.n20 12.0247
R2159 VDD2.n98 VDD2.n2 12.0247
R2160 VDD2.n202 VDD2.n109 11.249
R2161 VDD2.n171 VDD2.n170 11.249
R2162 VDD2.n154 VDD2.n131 11.249
R2163 VDD2.n48 VDD2.n26 11.249
R2164 VDD2.n66 VDD2.n65 11.249
R2165 VDD2.n97 VDD2.n4 11.249
R2166 VDD2.n141 VDD2.n139 10.7239
R2167 VDD2.n35 VDD2.n33 10.7239
R2168 VDD2.n199 VDD2.n198 10.4732
R2169 VDD2.n174 VDD2.n123 10.4732
R2170 VDD2.n153 VDD2.n134 10.4732
R2171 VDD2.n47 VDD2.n28 10.4732
R2172 VDD2.n69 VDD2.n18 10.4732
R2173 VDD2.n94 VDD2.n93 10.4732
R2174 VDD2.n195 VDD2.n111 9.69747
R2175 VDD2.n175 VDD2.n121 9.69747
R2176 VDD2.n150 VDD2.n149 9.69747
R2177 VDD2.n44 VDD2.n43 9.69747
R2178 VDD2.n70 VDD2.n16 9.69747
R2179 VDD2.n90 VDD2.n6 9.69747
R2180 VDD2.n209 VDD2.n208 9.45567
R2181 VDD2.n104 VDD2.n103 9.45567
R2182 VDD2.n143 VDD2.n142 9.3005
R2183 VDD2.n145 VDD2.n144 9.3005
R2184 VDD2.n136 VDD2.n135 9.3005
R2185 VDD2.n151 VDD2.n150 9.3005
R2186 VDD2.n153 VDD2.n152 9.3005
R2187 VDD2.n131 VDD2.n130 9.3005
R2188 VDD2.n159 VDD2.n158 9.3005
R2189 VDD2.n161 VDD2.n160 9.3005
R2190 VDD2.n115 VDD2.n114 9.3005
R2191 VDD2.n192 VDD2.n191 9.3005
R2192 VDD2.n194 VDD2.n193 9.3005
R2193 VDD2.n111 VDD2.n110 9.3005
R2194 VDD2.n200 VDD2.n199 9.3005
R2195 VDD2.n202 VDD2.n201 9.3005
R2196 VDD2.n107 VDD2.n106 9.3005
R2197 VDD2.n208 VDD2.n207 9.3005
R2198 VDD2.n186 VDD2.n185 9.3005
R2199 VDD2.n184 VDD2.n183 9.3005
R2200 VDD2.n119 VDD2.n118 9.3005
R2201 VDD2.n178 VDD2.n177 9.3005
R2202 VDD2.n176 VDD2.n175 9.3005
R2203 VDD2.n123 VDD2.n122 9.3005
R2204 VDD2.n170 VDD2.n169 9.3005
R2205 VDD2.n168 VDD2.n167 9.3005
R2206 VDD2.n127 VDD2.n126 9.3005
R2207 VDD2.n79 VDD2.n78 9.3005
R2208 VDD2.n14 VDD2.n13 9.3005
R2209 VDD2.n73 VDD2.n72 9.3005
R2210 VDD2.n71 VDD2.n70 9.3005
R2211 VDD2.n18 VDD2.n17 9.3005
R2212 VDD2.n65 VDD2.n64 9.3005
R2213 VDD2.n63 VDD2.n62 9.3005
R2214 VDD2.n22 VDD2.n21 9.3005
R2215 VDD2.n37 VDD2.n36 9.3005
R2216 VDD2.n39 VDD2.n38 9.3005
R2217 VDD2.n30 VDD2.n29 9.3005
R2218 VDD2.n45 VDD2.n44 9.3005
R2219 VDD2.n47 VDD2.n46 9.3005
R2220 VDD2.n26 VDD2.n25 9.3005
R2221 VDD2.n54 VDD2.n53 9.3005
R2222 VDD2.n56 VDD2.n55 9.3005
R2223 VDD2.n81 VDD2.n80 9.3005
R2224 VDD2.n10 VDD2.n9 9.3005
R2225 VDD2.n87 VDD2.n86 9.3005
R2226 VDD2.n89 VDD2.n88 9.3005
R2227 VDD2.n6 VDD2.n5 9.3005
R2228 VDD2.n95 VDD2.n94 9.3005
R2229 VDD2.n97 VDD2.n96 9.3005
R2230 VDD2.n2 VDD2.n1 9.3005
R2231 VDD2.n103 VDD2.n102 9.3005
R2232 VDD2.n194 VDD2.n113 8.92171
R2233 VDD2.n179 VDD2.n178 8.92171
R2234 VDD2.n146 VDD2.n136 8.92171
R2235 VDD2.n40 VDD2.n30 8.92171
R2236 VDD2.n74 VDD2.n73 8.92171
R2237 VDD2.n89 VDD2.n8 8.92171
R2238 VDD2.n191 VDD2.n190 8.14595
R2239 VDD2.n182 VDD2.n119 8.14595
R2240 VDD2.n145 VDD2.n138 8.14595
R2241 VDD2.n39 VDD2.n32 8.14595
R2242 VDD2.n77 VDD2.n14 8.14595
R2243 VDD2.n86 VDD2.n85 8.14595
R2244 VDD2.n209 VDD2.n105 7.75445
R2245 VDD2.n104 VDD2.n0 7.75445
R2246 VDD2.n187 VDD2.n115 7.3702
R2247 VDD2.n183 VDD2.n117 7.3702
R2248 VDD2.n142 VDD2.n141 7.3702
R2249 VDD2.n36 VDD2.n35 7.3702
R2250 VDD2.n78 VDD2.n12 7.3702
R2251 VDD2.n82 VDD2.n10 7.3702
R2252 VDD2.n187 VDD2.n186 6.59444
R2253 VDD2.n186 VDD2.n117 6.59444
R2254 VDD2.n81 VDD2.n12 6.59444
R2255 VDD2.n82 VDD2.n81 6.59444
R2256 VDD2.n207 VDD2.n105 6.08283
R2257 VDD2.n102 VDD2.n0 6.08283
R2258 VDD2.n190 VDD2.n115 5.81868
R2259 VDD2.n183 VDD2.n182 5.81868
R2260 VDD2.n142 VDD2.n138 5.81868
R2261 VDD2.n36 VDD2.n32 5.81868
R2262 VDD2.n78 VDD2.n77 5.81868
R2263 VDD2.n85 VDD2.n10 5.81868
R2264 VDD2.n191 VDD2.n113 5.04292
R2265 VDD2.n179 VDD2.n119 5.04292
R2266 VDD2.n146 VDD2.n145 5.04292
R2267 VDD2.n40 VDD2.n39 5.04292
R2268 VDD2.n74 VDD2.n14 5.04292
R2269 VDD2.n86 VDD2.n8 5.04292
R2270 VDD2.n195 VDD2.n194 4.26717
R2271 VDD2.n178 VDD2.n121 4.26717
R2272 VDD2.n149 VDD2.n136 4.26717
R2273 VDD2.n43 VDD2.n30 4.26717
R2274 VDD2.n73 VDD2.n16 4.26717
R2275 VDD2.n90 VDD2.n89 4.26717
R2276 VDD2.n198 VDD2.n111 3.49141
R2277 VDD2.n175 VDD2.n174 3.49141
R2278 VDD2.n150 VDD2.n134 3.49141
R2279 VDD2.n44 VDD2.n28 3.49141
R2280 VDD2.n70 VDD2.n69 3.49141
R2281 VDD2.n93 VDD2.n6 3.49141
R2282 VDD2.n199 VDD2.n109 2.71565
R2283 VDD2.n171 VDD2.n123 2.71565
R2284 VDD2.n154 VDD2.n153 2.71565
R2285 VDD2.n48 VDD2.n47 2.71565
R2286 VDD2.n66 VDD2.n18 2.71565
R2287 VDD2.n94 VDD2.n4 2.71565
R2288 VDD2.n143 VDD2.n139 2.41282
R2289 VDD2.n37 VDD2.n33 2.41282
R2290 VDD2.n203 VDD2.n202 1.93989
R2291 VDD2.n170 VDD2.n125 1.93989
R2292 VDD2.n157 VDD2.n131 1.93989
R2293 VDD2.n52 VDD2.n26 1.93989
R2294 VDD2.n65 VDD2.n20 1.93989
R2295 VDD2.n98 VDD2.n97 1.93989
R2296 VDD2.n206 VDD2.n107 1.16414
R2297 VDD2.n167 VDD2.n166 1.16414
R2298 VDD2.n158 VDD2.n129 1.16414
R2299 VDD2.n53 VDD2.n24 1.16414
R2300 VDD2.n62 VDD2.n61 1.16414
R2301 VDD2.n101 VDD2.n2 1.16414
R2302 VDD2 VDD2.n210 0.438
R2303 VDD2.n163 VDD2.n127 0.388379
R2304 VDD2.n162 VDD2.n161 0.388379
R2305 VDD2.n57 VDD2.n56 0.388379
R2306 VDD2.n58 VDD2.n22 0.388379
R2307 VDD2.n208 VDD2.n106 0.155672
R2308 VDD2.n201 VDD2.n106 0.155672
R2309 VDD2.n201 VDD2.n200 0.155672
R2310 VDD2.n200 VDD2.n110 0.155672
R2311 VDD2.n193 VDD2.n110 0.155672
R2312 VDD2.n193 VDD2.n192 0.155672
R2313 VDD2.n192 VDD2.n114 0.155672
R2314 VDD2.n185 VDD2.n114 0.155672
R2315 VDD2.n185 VDD2.n184 0.155672
R2316 VDD2.n184 VDD2.n118 0.155672
R2317 VDD2.n177 VDD2.n118 0.155672
R2318 VDD2.n177 VDD2.n176 0.155672
R2319 VDD2.n176 VDD2.n122 0.155672
R2320 VDD2.n169 VDD2.n122 0.155672
R2321 VDD2.n169 VDD2.n168 0.155672
R2322 VDD2.n168 VDD2.n126 0.155672
R2323 VDD2.n160 VDD2.n126 0.155672
R2324 VDD2.n160 VDD2.n159 0.155672
R2325 VDD2.n159 VDD2.n130 0.155672
R2326 VDD2.n152 VDD2.n130 0.155672
R2327 VDD2.n152 VDD2.n151 0.155672
R2328 VDD2.n151 VDD2.n135 0.155672
R2329 VDD2.n144 VDD2.n135 0.155672
R2330 VDD2.n144 VDD2.n143 0.155672
R2331 VDD2.n38 VDD2.n37 0.155672
R2332 VDD2.n38 VDD2.n29 0.155672
R2333 VDD2.n45 VDD2.n29 0.155672
R2334 VDD2.n46 VDD2.n45 0.155672
R2335 VDD2.n46 VDD2.n25 0.155672
R2336 VDD2.n54 VDD2.n25 0.155672
R2337 VDD2.n55 VDD2.n54 0.155672
R2338 VDD2.n55 VDD2.n21 0.155672
R2339 VDD2.n63 VDD2.n21 0.155672
R2340 VDD2.n64 VDD2.n63 0.155672
R2341 VDD2.n64 VDD2.n17 0.155672
R2342 VDD2.n71 VDD2.n17 0.155672
R2343 VDD2.n72 VDD2.n71 0.155672
R2344 VDD2.n72 VDD2.n13 0.155672
R2345 VDD2.n79 VDD2.n13 0.155672
R2346 VDD2.n80 VDD2.n79 0.155672
R2347 VDD2.n80 VDD2.n9 0.155672
R2348 VDD2.n87 VDD2.n9 0.155672
R2349 VDD2.n88 VDD2.n87 0.155672
R2350 VDD2.n88 VDD2.n5 0.155672
R2351 VDD2.n95 VDD2.n5 0.155672
R2352 VDD2.n96 VDD2.n95 0.155672
R2353 VDD2.n96 VDD2.n1 0.155672
R2354 VDD2.n103 VDD2.n1 0.155672
C0 w_n1674_n4862# VTAIL 3.92723f
C1 VP VTAIL 3.14335f
C2 w_n1674_n4862# B 9.6382f
C3 B VP 1.28149f
C4 VN VTAIL 3.12872f
C5 B VN 0.939766f
C6 VDD2 w_n1674_n4862# 2.19734f
C7 VDD2 VP 0.284932f
C8 VDD2 VN 3.85728f
C9 VTAIL VDD1 7.32557f
C10 B VDD1 2.10523f
C11 w_n1674_n4862# VP 2.55608f
C12 B VTAIL 4.61661f
C13 VDD2 VDD1 0.539812f
C14 w_n1674_n4862# VN 2.34536f
C15 VP VN 6.288549f
C16 VDD2 VTAIL 7.36366f
C17 VDD2 B 2.1251f
C18 w_n1674_n4862# VDD1 2.18527f
C19 VP VDD1 3.9893f
C20 VN VDD1 0.147586f
C21 VDD2 VSUBS 1.070869f
C22 VDD1 VSUBS 5.3073f
C23 VTAIL VSUBS 1.151385f
C24 VN VSUBS 9.235399f
C25 VP VSUBS 1.609614f
C26 B VSUBS 3.662663f
C27 w_n1674_n4862# VSUBS 99.4155f
C28 VDD2.n0 VSUBS 0.029916f
C29 VDD2.n1 VSUBS 0.027795f
C30 VDD2.n2 VSUBS 0.014936f
C31 VDD2.n3 VSUBS 0.035303f
C32 VDD2.n4 VSUBS 0.015815f
C33 VDD2.n5 VSUBS 0.027795f
C34 VDD2.n6 VSUBS 0.014936f
C35 VDD2.n7 VSUBS 0.035303f
C36 VDD2.n8 VSUBS 0.015815f
C37 VDD2.n9 VSUBS 0.027795f
C38 VDD2.n10 VSUBS 0.014936f
C39 VDD2.n11 VSUBS 0.035303f
C40 VDD2.n12 VSUBS 0.015815f
C41 VDD2.n13 VSUBS 0.027795f
C42 VDD2.n14 VSUBS 0.014936f
C43 VDD2.n15 VSUBS 0.035303f
C44 VDD2.n16 VSUBS 0.015815f
C45 VDD2.n17 VSUBS 0.027795f
C46 VDD2.n18 VSUBS 0.014936f
C47 VDD2.n19 VSUBS 0.035303f
C48 VDD2.n20 VSUBS 0.015815f
C49 VDD2.n21 VSUBS 0.027795f
C50 VDD2.n22 VSUBS 0.014936f
C51 VDD2.n23 VSUBS 0.035303f
C52 VDD2.n24 VSUBS 0.015815f
C53 VDD2.n25 VSUBS 0.027795f
C54 VDD2.n26 VSUBS 0.014936f
C55 VDD2.n27 VSUBS 0.035303f
C56 VDD2.n28 VSUBS 0.015815f
C57 VDD2.n29 VSUBS 0.027795f
C58 VDD2.n30 VSUBS 0.014936f
C59 VDD2.n31 VSUBS 0.035303f
C60 VDD2.n32 VSUBS 0.015815f
C61 VDD2.n33 VSUBS 0.312788f
C62 VDD2.t0 VSUBS 0.076777f
C63 VDD2.n34 VSUBS 0.026478f
C64 VDD2.n35 VSUBS 0.026557f
C65 VDD2.n36 VSUBS 0.014936f
C66 VDD2.n37 VSUBS 2.27545f
C67 VDD2.n38 VSUBS 0.027795f
C68 VDD2.n39 VSUBS 0.014936f
C69 VDD2.n40 VSUBS 0.015815f
C70 VDD2.n41 VSUBS 0.035303f
C71 VDD2.n42 VSUBS 0.035303f
C72 VDD2.n43 VSUBS 0.015815f
C73 VDD2.n44 VSUBS 0.014936f
C74 VDD2.n45 VSUBS 0.027795f
C75 VDD2.n46 VSUBS 0.027795f
C76 VDD2.n47 VSUBS 0.014936f
C77 VDD2.n48 VSUBS 0.015815f
C78 VDD2.n49 VSUBS 0.035303f
C79 VDD2.n50 VSUBS 0.035303f
C80 VDD2.n51 VSUBS 0.035303f
C81 VDD2.n52 VSUBS 0.015815f
C82 VDD2.n53 VSUBS 0.014936f
C83 VDD2.n54 VSUBS 0.027795f
C84 VDD2.n55 VSUBS 0.027795f
C85 VDD2.n56 VSUBS 0.014936f
C86 VDD2.n57 VSUBS 0.015375f
C87 VDD2.n58 VSUBS 0.015375f
C88 VDD2.n59 VSUBS 0.035303f
C89 VDD2.n60 VSUBS 0.035303f
C90 VDD2.n61 VSUBS 0.015815f
C91 VDD2.n62 VSUBS 0.014936f
C92 VDD2.n63 VSUBS 0.027795f
C93 VDD2.n64 VSUBS 0.027795f
C94 VDD2.n65 VSUBS 0.014936f
C95 VDD2.n66 VSUBS 0.015815f
C96 VDD2.n67 VSUBS 0.035303f
C97 VDD2.n68 VSUBS 0.035303f
C98 VDD2.n69 VSUBS 0.015815f
C99 VDD2.n70 VSUBS 0.014936f
C100 VDD2.n71 VSUBS 0.027795f
C101 VDD2.n72 VSUBS 0.027795f
C102 VDD2.n73 VSUBS 0.014936f
C103 VDD2.n74 VSUBS 0.015815f
C104 VDD2.n75 VSUBS 0.035303f
C105 VDD2.n76 VSUBS 0.035303f
C106 VDD2.n77 VSUBS 0.015815f
C107 VDD2.n78 VSUBS 0.014936f
C108 VDD2.n79 VSUBS 0.027795f
C109 VDD2.n80 VSUBS 0.027795f
C110 VDD2.n81 VSUBS 0.014936f
C111 VDD2.n82 VSUBS 0.015815f
C112 VDD2.n83 VSUBS 0.035303f
C113 VDD2.n84 VSUBS 0.035303f
C114 VDD2.n85 VSUBS 0.015815f
C115 VDD2.n86 VSUBS 0.014936f
C116 VDD2.n87 VSUBS 0.027795f
C117 VDD2.n88 VSUBS 0.027795f
C118 VDD2.n89 VSUBS 0.014936f
C119 VDD2.n90 VSUBS 0.015815f
C120 VDD2.n91 VSUBS 0.035303f
C121 VDD2.n92 VSUBS 0.035303f
C122 VDD2.n93 VSUBS 0.015815f
C123 VDD2.n94 VSUBS 0.014936f
C124 VDD2.n95 VSUBS 0.027795f
C125 VDD2.n96 VSUBS 0.027795f
C126 VDD2.n97 VSUBS 0.014936f
C127 VDD2.n98 VSUBS 0.015815f
C128 VDD2.n99 VSUBS 0.035303f
C129 VDD2.n100 VSUBS 0.087644f
C130 VDD2.n101 VSUBS 0.015815f
C131 VDD2.n102 VSUBS 0.029331f
C132 VDD2.n103 VSUBS 0.069944f
C133 VDD2.n104 VSUBS 1.03365f
C134 VDD2.n105 VSUBS 0.029916f
C135 VDD2.n106 VSUBS 0.027795f
C136 VDD2.n107 VSUBS 0.014936f
C137 VDD2.n108 VSUBS 0.035303f
C138 VDD2.n109 VSUBS 0.015815f
C139 VDD2.n110 VSUBS 0.027795f
C140 VDD2.n111 VSUBS 0.014936f
C141 VDD2.n112 VSUBS 0.035303f
C142 VDD2.n113 VSUBS 0.015815f
C143 VDD2.n114 VSUBS 0.027795f
C144 VDD2.n115 VSUBS 0.014936f
C145 VDD2.n116 VSUBS 0.035303f
C146 VDD2.n117 VSUBS 0.015815f
C147 VDD2.n118 VSUBS 0.027795f
C148 VDD2.n119 VSUBS 0.014936f
C149 VDD2.n120 VSUBS 0.035303f
C150 VDD2.n121 VSUBS 0.015815f
C151 VDD2.n122 VSUBS 0.027795f
C152 VDD2.n123 VSUBS 0.014936f
C153 VDD2.n124 VSUBS 0.035303f
C154 VDD2.n125 VSUBS 0.015815f
C155 VDD2.n126 VSUBS 0.027795f
C156 VDD2.n127 VSUBS 0.014936f
C157 VDD2.n128 VSUBS 0.035303f
C158 VDD2.n129 VSUBS 0.015815f
C159 VDD2.n130 VSUBS 0.027795f
C160 VDD2.n131 VSUBS 0.014936f
C161 VDD2.n132 VSUBS 0.035303f
C162 VDD2.n133 VSUBS 0.035303f
C163 VDD2.n134 VSUBS 0.015815f
C164 VDD2.n135 VSUBS 0.027795f
C165 VDD2.n136 VSUBS 0.014936f
C166 VDD2.n137 VSUBS 0.035303f
C167 VDD2.n138 VSUBS 0.015815f
C168 VDD2.n139 VSUBS 0.312788f
C169 VDD2.t1 VSUBS 0.076777f
C170 VDD2.n140 VSUBS 0.026478f
C171 VDD2.n141 VSUBS 0.026557f
C172 VDD2.n142 VSUBS 0.014936f
C173 VDD2.n143 VSUBS 2.27545f
C174 VDD2.n144 VSUBS 0.027795f
C175 VDD2.n145 VSUBS 0.014936f
C176 VDD2.n146 VSUBS 0.015815f
C177 VDD2.n147 VSUBS 0.035303f
C178 VDD2.n148 VSUBS 0.035303f
C179 VDD2.n149 VSUBS 0.015815f
C180 VDD2.n150 VSUBS 0.014936f
C181 VDD2.n151 VSUBS 0.027795f
C182 VDD2.n152 VSUBS 0.027795f
C183 VDD2.n153 VSUBS 0.014936f
C184 VDD2.n154 VSUBS 0.015815f
C185 VDD2.n155 VSUBS 0.035303f
C186 VDD2.n156 VSUBS 0.035303f
C187 VDD2.n157 VSUBS 0.015815f
C188 VDD2.n158 VSUBS 0.014936f
C189 VDD2.n159 VSUBS 0.027795f
C190 VDD2.n160 VSUBS 0.027795f
C191 VDD2.n161 VSUBS 0.014936f
C192 VDD2.n162 VSUBS 0.015375f
C193 VDD2.n163 VSUBS 0.015375f
C194 VDD2.n164 VSUBS 0.035303f
C195 VDD2.n165 VSUBS 0.035303f
C196 VDD2.n166 VSUBS 0.015815f
C197 VDD2.n167 VSUBS 0.014936f
C198 VDD2.n168 VSUBS 0.027795f
C199 VDD2.n169 VSUBS 0.027795f
C200 VDD2.n170 VSUBS 0.014936f
C201 VDD2.n171 VSUBS 0.015815f
C202 VDD2.n172 VSUBS 0.035303f
C203 VDD2.n173 VSUBS 0.035303f
C204 VDD2.n174 VSUBS 0.015815f
C205 VDD2.n175 VSUBS 0.014936f
C206 VDD2.n176 VSUBS 0.027795f
C207 VDD2.n177 VSUBS 0.027795f
C208 VDD2.n178 VSUBS 0.014936f
C209 VDD2.n179 VSUBS 0.015815f
C210 VDD2.n180 VSUBS 0.035303f
C211 VDD2.n181 VSUBS 0.035303f
C212 VDD2.n182 VSUBS 0.015815f
C213 VDD2.n183 VSUBS 0.014936f
C214 VDD2.n184 VSUBS 0.027795f
C215 VDD2.n185 VSUBS 0.027795f
C216 VDD2.n186 VSUBS 0.014936f
C217 VDD2.n187 VSUBS 0.015815f
C218 VDD2.n188 VSUBS 0.035303f
C219 VDD2.n189 VSUBS 0.035303f
C220 VDD2.n190 VSUBS 0.015815f
C221 VDD2.n191 VSUBS 0.014936f
C222 VDD2.n192 VSUBS 0.027795f
C223 VDD2.n193 VSUBS 0.027795f
C224 VDD2.n194 VSUBS 0.014936f
C225 VDD2.n195 VSUBS 0.015815f
C226 VDD2.n196 VSUBS 0.035303f
C227 VDD2.n197 VSUBS 0.035303f
C228 VDD2.n198 VSUBS 0.015815f
C229 VDD2.n199 VSUBS 0.014936f
C230 VDD2.n200 VSUBS 0.027795f
C231 VDD2.n201 VSUBS 0.027795f
C232 VDD2.n202 VSUBS 0.014936f
C233 VDD2.n203 VSUBS 0.015815f
C234 VDD2.n204 VSUBS 0.035303f
C235 VDD2.n205 VSUBS 0.087644f
C236 VDD2.n206 VSUBS 0.015815f
C237 VDD2.n207 VSUBS 0.029331f
C238 VDD2.n208 VSUBS 0.069944f
C239 VDD2.n209 VSUBS 0.086258f
C240 VDD2.n210 VSUBS 4.02336f
C241 VN.t1 VSUBS 4.11181f
C242 VN.t0 VSUBS 4.47093f
C243 B.n0 VSUBS 0.006862f
C244 B.n1 VSUBS 0.006862f
C245 B.n2 VSUBS 0.010149f
C246 B.n3 VSUBS 0.007777f
C247 B.n4 VSUBS 0.007777f
C248 B.n5 VSUBS 0.007777f
C249 B.n6 VSUBS 0.007777f
C250 B.n7 VSUBS 0.007777f
C251 B.n8 VSUBS 0.007777f
C252 B.n9 VSUBS 0.007777f
C253 B.n10 VSUBS 0.007777f
C254 B.n11 VSUBS 0.018035f
C255 B.n12 VSUBS 0.007777f
C256 B.n13 VSUBS 0.007777f
C257 B.n14 VSUBS 0.007777f
C258 B.n15 VSUBS 0.007777f
C259 B.n16 VSUBS 0.007777f
C260 B.n17 VSUBS 0.007777f
C261 B.n18 VSUBS 0.007777f
C262 B.n19 VSUBS 0.007777f
C263 B.n20 VSUBS 0.007777f
C264 B.n21 VSUBS 0.007777f
C265 B.n22 VSUBS 0.007777f
C266 B.n23 VSUBS 0.007777f
C267 B.n24 VSUBS 0.007777f
C268 B.n25 VSUBS 0.007777f
C269 B.n26 VSUBS 0.007777f
C270 B.n27 VSUBS 0.007777f
C271 B.n28 VSUBS 0.007777f
C272 B.n29 VSUBS 0.007777f
C273 B.n30 VSUBS 0.007777f
C274 B.n31 VSUBS 0.007777f
C275 B.n32 VSUBS 0.007777f
C276 B.n33 VSUBS 0.007777f
C277 B.n34 VSUBS 0.007777f
C278 B.n35 VSUBS 0.007777f
C279 B.n36 VSUBS 0.007777f
C280 B.n37 VSUBS 0.007777f
C281 B.n38 VSUBS 0.007777f
C282 B.n39 VSUBS 0.007777f
C283 B.n40 VSUBS 0.007777f
C284 B.n41 VSUBS 0.007777f
C285 B.n42 VSUBS 0.007777f
C286 B.n43 VSUBS 0.007777f
C287 B.t7 VSUBS 0.429683f
C288 B.t8 VSUBS 0.452775f
C289 B.t6 VSUBS 1.30377f
C290 B.n44 VSUBS 0.616958f
C291 B.n45 VSUBS 0.379266f
C292 B.n46 VSUBS 0.007777f
C293 B.n47 VSUBS 0.007777f
C294 B.n48 VSUBS 0.007777f
C295 B.n49 VSUBS 0.007777f
C296 B.t10 VSUBS 0.429687f
C297 B.t11 VSUBS 0.452779f
C298 B.t9 VSUBS 1.30377f
C299 B.n50 VSUBS 0.616954f
C300 B.n51 VSUBS 0.379262f
C301 B.n52 VSUBS 0.007777f
C302 B.n53 VSUBS 0.007777f
C303 B.n54 VSUBS 0.007777f
C304 B.n55 VSUBS 0.007777f
C305 B.n56 VSUBS 0.007777f
C306 B.n57 VSUBS 0.007777f
C307 B.n58 VSUBS 0.007777f
C308 B.n59 VSUBS 0.007777f
C309 B.n60 VSUBS 0.007777f
C310 B.n61 VSUBS 0.007777f
C311 B.n62 VSUBS 0.007777f
C312 B.n63 VSUBS 0.007777f
C313 B.n64 VSUBS 0.007777f
C314 B.n65 VSUBS 0.007777f
C315 B.n66 VSUBS 0.007777f
C316 B.n67 VSUBS 0.007777f
C317 B.n68 VSUBS 0.007777f
C318 B.n69 VSUBS 0.007777f
C319 B.n70 VSUBS 0.007777f
C320 B.n71 VSUBS 0.007777f
C321 B.n72 VSUBS 0.007777f
C322 B.n73 VSUBS 0.007777f
C323 B.n74 VSUBS 0.007777f
C324 B.n75 VSUBS 0.007777f
C325 B.n76 VSUBS 0.007777f
C326 B.n77 VSUBS 0.007777f
C327 B.n78 VSUBS 0.007777f
C328 B.n79 VSUBS 0.007777f
C329 B.n80 VSUBS 0.007777f
C330 B.n81 VSUBS 0.007777f
C331 B.n82 VSUBS 0.007777f
C332 B.n83 VSUBS 0.018035f
C333 B.n84 VSUBS 0.007777f
C334 B.n85 VSUBS 0.007777f
C335 B.n86 VSUBS 0.007777f
C336 B.n87 VSUBS 0.007777f
C337 B.n88 VSUBS 0.007777f
C338 B.n89 VSUBS 0.007777f
C339 B.n90 VSUBS 0.007777f
C340 B.n91 VSUBS 0.007777f
C341 B.n92 VSUBS 0.007777f
C342 B.n93 VSUBS 0.007777f
C343 B.n94 VSUBS 0.007777f
C344 B.n95 VSUBS 0.007777f
C345 B.n96 VSUBS 0.007777f
C346 B.n97 VSUBS 0.007777f
C347 B.n98 VSUBS 0.007777f
C348 B.n99 VSUBS 0.007777f
C349 B.n100 VSUBS 0.007777f
C350 B.n101 VSUBS 0.007777f
C351 B.n102 VSUBS 0.01794f
C352 B.n103 VSUBS 0.007777f
C353 B.n104 VSUBS 0.007777f
C354 B.n105 VSUBS 0.007777f
C355 B.n106 VSUBS 0.007777f
C356 B.n107 VSUBS 0.007777f
C357 B.n108 VSUBS 0.007777f
C358 B.n109 VSUBS 0.007777f
C359 B.n110 VSUBS 0.007777f
C360 B.n111 VSUBS 0.007777f
C361 B.n112 VSUBS 0.007777f
C362 B.n113 VSUBS 0.007777f
C363 B.n114 VSUBS 0.007777f
C364 B.n115 VSUBS 0.007777f
C365 B.n116 VSUBS 0.007777f
C366 B.n117 VSUBS 0.007777f
C367 B.n118 VSUBS 0.007777f
C368 B.n119 VSUBS 0.007777f
C369 B.n120 VSUBS 0.007777f
C370 B.n121 VSUBS 0.007777f
C371 B.n122 VSUBS 0.007777f
C372 B.n123 VSUBS 0.007777f
C373 B.n124 VSUBS 0.007777f
C374 B.n125 VSUBS 0.007777f
C375 B.n126 VSUBS 0.007777f
C376 B.n127 VSUBS 0.007777f
C377 B.n128 VSUBS 0.007777f
C378 B.n129 VSUBS 0.007777f
C379 B.n130 VSUBS 0.007777f
C380 B.n131 VSUBS 0.007777f
C381 B.n132 VSUBS 0.007777f
C382 B.n133 VSUBS 0.007777f
C383 B.n134 VSUBS 0.005376f
C384 B.n135 VSUBS 0.007777f
C385 B.n136 VSUBS 0.007777f
C386 B.n137 VSUBS 0.007777f
C387 B.n138 VSUBS 0.007777f
C388 B.n139 VSUBS 0.007777f
C389 B.t2 VSUBS 0.429683f
C390 B.t1 VSUBS 0.452775f
C391 B.t0 VSUBS 1.30377f
C392 B.n140 VSUBS 0.616958f
C393 B.n141 VSUBS 0.379266f
C394 B.n142 VSUBS 0.007777f
C395 B.n143 VSUBS 0.007777f
C396 B.n144 VSUBS 0.007777f
C397 B.n145 VSUBS 0.007777f
C398 B.n146 VSUBS 0.007777f
C399 B.n147 VSUBS 0.007777f
C400 B.n148 VSUBS 0.007777f
C401 B.n149 VSUBS 0.007777f
C402 B.n150 VSUBS 0.007777f
C403 B.n151 VSUBS 0.007777f
C404 B.n152 VSUBS 0.007777f
C405 B.n153 VSUBS 0.007777f
C406 B.n154 VSUBS 0.007777f
C407 B.n155 VSUBS 0.007777f
C408 B.n156 VSUBS 0.007777f
C409 B.n157 VSUBS 0.007777f
C410 B.n158 VSUBS 0.007777f
C411 B.n159 VSUBS 0.007777f
C412 B.n160 VSUBS 0.007777f
C413 B.n161 VSUBS 0.007777f
C414 B.n162 VSUBS 0.007777f
C415 B.n163 VSUBS 0.007777f
C416 B.n164 VSUBS 0.007777f
C417 B.n165 VSUBS 0.007777f
C418 B.n166 VSUBS 0.007777f
C419 B.n167 VSUBS 0.007777f
C420 B.n168 VSUBS 0.007777f
C421 B.n169 VSUBS 0.007777f
C422 B.n170 VSUBS 0.007777f
C423 B.n171 VSUBS 0.007777f
C424 B.n172 VSUBS 0.007777f
C425 B.n173 VSUBS 0.016964f
C426 B.n174 VSUBS 0.007777f
C427 B.n175 VSUBS 0.007777f
C428 B.n176 VSUBS 0.007777f
C429 B.n177 VSUBS 0.007777f
C430 B.n178 VSUBS 0.007777f
C431 B.n179 VSUBS 0.007777f
C432 B.n180 VSUBS 0.007777f
C433 B.n181 VSUBS 0.007777f
C434 B.n182 VSUBS 0.007777f
C435 B.n183 VSUBS 0.007777f
C436 B.n184 VSUBS 0.007777f
C437 B.n185 VSUBS 0.007777f
C438 B.n186 VSUBS 0.007777f
C439 B.n187 VSUBS 0.007777f
C440 B.n188 VSUBS 0.007777f
C441 B.n189 VSUBS 0.007777f
C442 B.n190 VSUBS 0.007777f
C443 B.n191 VSUBS 0.007777f
C444 B.n192 VSUBS 0.007777f
C445 B.n193 VSUBS 0.007777f
C446 B.n194 VSUBS 0.007777f
C447 B.n195 VSUBS 0.007777f
C448 B.n196 VSUBS 0.007777f
C449 B.n197 VSUBS 0.007777f
C450 B.n198 VSUBS 0.007777f
C451 B.n199 VSUBS 0.007777f
C452 B.n200 VSUBS 0.007777f
C453 B.n201 VSUBS 0.007777f
C454 B.n202 VSUBS 0.007777f
C455 B.n203 VSUBS 0.007777f
C456 B.n204 VSUBS 0.007777f
C457 B.n205 VSUBS 0.007777f
C458 B.n206 VSUBS 0.016964f
C459 B.n207 VSUBS 0.018035f
C460 B.n208 VSUBS 0.018035f
C461 B.n209 VSUBS 0.007777f
C462 B.n210 VSUBS 0.007777f
C463 B.n211 VSUBS 0.007777f
C464 B.n212 VSUBS 0.007777f
C465 B.n213 VSUBS 0.007777f
C466 B.n214 VSUBS 0.007777f
C467 B.n215 VSUBS 0.007777f
C468 B.n216 VSUBS 0.007777f
C469 B.n217 VSUBS 0.007777f
C470 B.n218 VSUBS 0.007777f
C471 B.n219 VSUBS 0.007777f
C472 B.n220 VSUBS 0.007777f
C473 B.n221 VSUBS 0.007777f
C474 B.n222 VSUBS 0.007777f
C475 B.n223 VSUBS 0.007777f
C476 B.n224 VSUBS 0.007777f
C477 B.n225 VSUBS 0.007777f
C478 B.n226 VSUBS 0.007777f
C479 B.n227 VSUBS 0.007777f
C480 B.n228 VSUBS 0.007777f
C481 B.n229 VSUBS 0.007777f
C482 B.n230 VSUBS 0.007777f
C483 B.n231 VSUBS 0.007777f
C484 B.n232 VSUBS 0.007777f
C485 B.n233 VSUBS 0.007777f
C486 B.n234 VSUBS 0.007777f
C487 B.n235 VSUBS 0.007777f
C488 B.n236 VSUBS 0.007777f
C489 B.n237 VSUBS 0.007777f
C490 B.n238 VSUBS 0.007777f
C491 B.n239 VSUBS 0.007777f
C492 B.n240 VSUBS 0.007777f
C493 B.n241 VSUBS 0.007777f
C494 B.n242 VSUBS 0.007777f
C495 B.n243 VSUBS 0.007777f
C496 B.n244 VSUBS 0.007777f
C497 B.n245 VSUBS 0.007777f
C498 B.n246 VSUBS 0.007777f
C499 B.n247 VSUBS 0.007777f
C500 B.n248 VSUBS 0.007777f
C501 B.n249 VSUBS 0.007777f
C502 B.n250 VSUBS 0.007777f
C503 B.n251 VSUBS 0.007777f
C504 B.n252 VSUBS 0.007777f
C505 B.n253 VSUBS 0.007777f
C506 B.n254 VSUBS 0.007777f
C507 B.n255 VSUBS 0.007777f
C508 B.n256 VSUBS 0.007777f
C509 B.n257 VSUBS 0.007777f
C510 B.n258 VSUBS 0.007777f
C511 B.n259 VSUBS 0.007777f
C512 B.n260 VSUBS 0.007777f
C513 B.n261 VSUBS 0.007777f
C514 B.n262 VSUBS 0.007777f
C515 B.n263 VSUBS 0.007777f
C516 B.n264 VSUBS 0.007777f
C517 B.n265 VSUBS 0.007777f
C518 B.n266 VSUBS 0.007777f
C519 B.n267 VSUBS 0.007777f
C520 B.n268 VSUBS 0.007777f
C521 B.n269 VSUBS 0.007777f
C522 B.n270 VSUBS 0.007777f
C523 B.n271 VSUBS 0.007777f
C524 B.n272 VSUBS 0.007777f
C525 B.n273 VSUBS 0.007777f
C526 B.n274 VSUBS 0.007777f
C527 B.n275 VSUBS 0.007777f
C528 B.n276 VSUBS 0.007777f
C529 B.n277 VSUBS 0.007777f
C530 B.n278 VSUBS 0.007777f
C531 B.n279 VSUBS 0.007777f
C532 B.n280 VSUBS 0.007777f
C533 B.n281 VSUBS 0.007777f
C534 B.n282 VSUBS 0.007777f
C535 B.n283 VSUBS 0.007777f
C536 B.n284 VSUBS 0.007777f
C537 B.n285 VSUBS 0.007777f
C538 B.n286 VSUBS 0.007777f
C539 B.n287 VSUBS 0.007777f
C540 B.n288 VSUBS 0.007777f
C541 B.n289 VSUBS 0.007777f
C542 B.n290 VSUBS 0.007777f
C543 B.n291 VSUBS 0.007777f
C544 B.n292 VSUBS 0.007777f
C545 B.n293 VSUBS 0.007777f
C546 B.n294 VSUBS 0.007777f
C547 B.n295 VSUBS 0.007777f
C548 B.n296 VSUBS 0.007777f
C549 B.n297 VSUBS 0.007777f
C550 B.n298 VSUBS 0.007777f
C551 B.n299 VSUBS 0.007777f
C552 B.n300 VSUBS 0.007777f
C553 B.n301 VSUBS 0.007777f
C554 B.n302 VSUBS 0.005376f
C555 B.n303 VSUBS 0.018019f
C556 B.n304 VSUBS 0.006291f
C557 B.n305 VSUBS 0.007777f
C558 B.n306 VSUBS 0.007777f
C559 B.n307 VSUBS 0.007777f
C560 B.n308 VSUBS 0.007777f
C561 B.n309 VSUBS 0.007777f
C562 B.n310 VSUBS 0.007777f
C563 B.n311 VSUBS 0.007777f
C564 B.n312 VSUBS 0.007777f
C565 B.n313 VSUBS 0.007777f
C566 B.n314 VSUBS 0.007777f
C567 B.n315 VSUBS 0.007777f
C568 B.t5 VSUBS 0.429687f
C569 B.t4 VSUBS 0.452779f
C570 B.t3 VSUBS 1.30377f
C571 B.n316 VSUBS 0.616954f
C572 B.n317 VSUBS 0.379262f
C573 B.n318 VSUBS 0.018019f
C574 B.n319 VSUBS 0.006291f
C575 B.n320 VSUBS 0.007777f
C576 B.n321 VSUBS 0.007777f
C577 B.n322 VSUBS 0.007777f
C578 B.n323 VSUBS 0.007777f
C579 B.n324 VSUBS 0.007777f
C580 B.n325 VSUBS 0.007777f
C581 B.n326 VSUBS 0.007777f
C582 B.n327 VSUBS 0.007777f
C583 B.n328 VSUBS 0.007777f
C584 B.n329 VSUBS 0.007777f
C585 B.n330 VSUBS 0.007777f
C586 B.n331 VSUBS 0.007777f
C587 B.n332 VSUBS 0.007777f
C588 B.n333 VSUBS 0.007777f
C589 B.n334 VSUBS 0.007777f
C590 B.n335 VSUBS 0.007777f
C591 B.n336 VSUBS 0.007777f
C592 B.n337 VSUBS 0.007777f
C593 B.n338 VSUBS 0.007777f
C594 B.n339 VSUBS 0.007777f
C595 B.n340 VSUBS 0.007777f
C596 B.n341 VSUBS 0.007777f
C597 B.n342 VSUBS 0.007777f
C598 B.n343 VSUBS 0.007777f
C599 B.n344 VSUBS 0.007777f
C600 B.n345 VSUBS 0.007777f
C601 B.n346 VSUBS 0.007777f
C602 B.n347 VSUBS 0.007777f
C603 B.n348 VSUBS 0.007777f
C604 B.n349 VSUBS 0.007777f
C605 B.n350 VSUBS 0.007777f
C606 B.n351 VSUBS 0.007777f
C607 B.n352 VSUBS 0.007777f
C608 B.n353 VSUBS 0.007777f
C609 B.n354 VSUBS 0.007777f
C610 B.n355 VSUBS 0.007777f
C611 B.n356 VSUBS 0.007777f
C612 B.n357 VSUBS 0.007777f
C613 B.n358 VSUBS 0.007777f
C614 B.n359 VSUBS 0.007777f
C615 B.n360 VSUBS 0.007777f
C616 B.n361 VSUBS 0.007777f
C617 B.n362 VSUBS 0.007777f
C618 B.n363 VSUBS 0.007777f
C619 B.n364 VSUBS 0.007777f
C620 B.n365 VSUBS 0.007777f
C621 B.n366 VSUBS 0.007777f
C622 B.n367 VSUBS 0.007777f
C623 B.n368 VSUBS 0.007777f
C624 B.n369 VSUBS 0.007777f
C625 B.n370 VSUBS 0.007777f
C626 B.n371 VSUBS 0.007777f
C627 B.n372 VSUBS 0.007777f
C628 B.n373 VSUBS 0.007777f
C629 B.n374 VSUBS 0.007777f
C630 B.n375 VSUBS 0.007777f
C631 B.n376 VSUBS 0.007777f
C632 B.n377 VSUBS 0.007777f
C633 B.n378 VSUBS 0.007777f
C634 B.n379 VSUBS 0.007777f
C635 B.n380 VSUBS 0.007777f
C636 B.n381 VSUBS 0.007777f
C637 B.n382 VSUBS 0.007777f
C638 B.n383 VSUBS 0.007777f
C639 B.n384 VSUBS 0.007777f
C640 B.n385 VSUBS 0.007777f
C641 B.n386 VSUBS 0.007777f
C642 B.n387 VSUBS 0.007777f
C643 B.n388 VSUBS 0.007777f
C644 B.n389 VSUBS 0.007777f
C645 B.n390 VSUBS 0.007777f
C646 B.n391 VSUBS 0.007777f
C647 B.n392 VSUBS 0.007777f
C648 B.n393 VSUBS 0.007777f
C649 B.n394 VSUBS 0.007777f
C650 B.n395 VSUBS 0.007777f
C651 B.n396 VSUBS 0.007777f
C652 B.n397 VSUBS 0.007777f
C653 B.n398 VSUBS 0.007777f
C654 B.n399 VSUBS 0.007777f
C655 B.n400 VSUBS 0.007777f
C656 B.n401 VSUBS 0.007777f
C657 B.n402 VSUBS 0.007777f
C658 B.n403 VSUBS 0.007777f
C659 B.n404 VSUBS 0.007777f
C660 B.n405 VSUBS 0.007777f
C661 B.n406 VSUBS 0.007777f
C662 B.n407 VSUBS 0.007777f
C663 B.n408 VSUBS 0.007777f
C664 B.n409 VSUBS 0.007777f
C665 B.n410 VSUBS 0.007777f
C666 B.n411 VSUBS 0.007777f
C667 B.n412 VSUBS 0.007777f
C668 B.n413 VSUBS 0.007777f
C669 B.n414 VSUBS 0.007777f
C670 B.n415 VSUBS 0.017059f
C671 B.n416 VSUBS 0.018035f
C672 B.n417 VSUBS 0.016964f
C673 B.n418 VSUBS 0.007777f
C674 B.n419 VSUBS 0.007777f
C675 B.n420 VSUBS 0.007777f
C676 B.n421 VSUBS 0.007777f
C677 B.n422 VSUBS 0.007777f
C678 B.n423 VSUBS 0.007777f
C679 B.n424 VSUBS 0.007777f
C680 B.n425 VSUBS 0.007777f
C681 B.n426 VSUBS 0.007777f
C682 B.n427 VSUBS 0.007777f
C683 B.n428 VSUBS 0.007777f
C684 B.n429 VSUBS 0.007777f
C685 B.n430 VSUBS 0.007777f
C686 B.n431 VSUBS 0.007777f
C687 B.n432 VSUBS 0.007777f
C688 B.n433 VSUBS 0.007777f
C689 B.n434 VSUBS 0.007777f
C690 B.n435 VSUBS 0.007777f
C691 B.n436 VSUBS 0.007777f
C692 B.n437 VSUBS 0.007777f
C693 B.n438 VSUBS 0.007777f
C694 B.n439 VSUBS 0.007777f
C695 B.n440 VSUBS 0.007777f
C696 B.n441 VSUBS 0.007777f
C697 B.n442 VSUBS 0.007777f
C698 B.n443 VSUBS 0.007777f
C699 B.n444 VSUBS 0.007777f
C700 B.n445 VSUBS 0.007777f
C701 B.n446 VSUBS 0.007777f
C702 B.n447 VSUBS 0.007777f
C703 B.n448 VSUBS 0.007777f
C704 B.n449 VSUBS 0.007777f
C705 B.n450 VSUBS 0.007777f
C706 B.n451 VSUBS 0.007777f
C707 B.n452 VSUBS 0.007777f
C708 B.n453 VSUBS 0.007777f
C709 B.n454 VSUBS 0.007777f
C710 B.n455 VSUBS 0.007777f
C711 B.n456 VSUBS 0.007777f
C712 B.n457 VSUBS 0.007777f
C713 B.n458 VSUBS 0.007777f
C714 B.n459 VSUBS 0.007777f
C715 B.n460 VSUBS 0.007777f
C716 B.n461 VSUBS 0.007777f
C717 B.n462 VSUBS 0.007777f
C718 B.n463 VSUBS 0.007777f
C719 B.n464 VSUBS 0.007777f
C720 B.n465 VSUBS 0.007777f
C721 B.n466 VSUBS 0.007777f
C722 B.n467 VSUBS 0.007777f
C723 B.n468 VSUBS 0.007777f
C724 B.n469 VSUBS 0.007777f
C725 B.n470 VSUBS 0.007777f
C726 B.n471 VSUBS 0.007777f
C727 B.n472 VSUBS 0.016964f
C728 B.n473 VSUBS 0.016964f
C729 B.n474 VSUBS 0.018035f
C730 B.n475 VSUBS 0.007777f
C731 B.n476 VSUBS 0.007777f
C732 B.n477 VSUBS 0.007777f
C733 B.n478 VSUBS 0.007777f
C734 B.n479 VSUBS 0.007777f
C735 B.n480 VSUBS 0.007777f
C736 B.n481 VSUBS 0.007777f
C737 B.n482 VSUBS 0.007777f
C738 B.n483 VSUBS 0.007777f
C739 B.n484 VSUBS 0.007777f
C740 B.n485 VSUBS 0.007777f
C741 B.n486 VSUBS 0.007777f
C742 B.n487 VSUBS 0.007777f
C743 B.n488 VSUBS 0.007777f
C744 B.n489 VSUBS 0.007777f
C745 B.n490 VSUBS 0.007777f
C746 B.n491 VSUBS 0.007777f
C747 B.n492 VSUBS 0.007777f
C748 B.n493 VSUBS 0.007777f
C749 B.n494 VSUBS 0.007777f
C750 B.n495 VSUBS 0.007777f
C751 B.n496 VSUBS 0.007777f
C752 B.n497 VSUBS 0.007777f
C753 B.n498 VSUBS 0.007777f
C754 B.n499 VSUBS 0.007777f
C755 B.n500 VSUBS 0.007777f
C756 B.n501 VSUBS 0.007777f
C757 B.n502 VSUBS 0.007777f
C758 B.n503 VSUBS 0.007777f
C759 B.n504 VSUBS 0.007777f
C760 B.n505 VSUBS 0.007777f
C761 B.n506 VSUBS 0.007777f
C762 B.n507 VSUBS 0.007777f
C763 B.n508 VSUBS 0.007777f
C764 B.n509 VSUBS 0.007777f
C765 B.n510 VSUBS 0.007777f
C766 B.n511 VSUBS 0.007777f
C767 B.n512 VSUBS 0.007777f
C768 B.n513 VSUBS 0.007777f
C769 B.n514 VSUBS 0.007777f
C770 B.n515 VSUBS 0.007777f
C771 B.n516 VSUBS 0.007777f
C772 B.n517 VSUBS 0.007777f
C773 B.n518 VSUBS 0.007777f
C774 B.n519 VSUBS 0.007777f
C775 B.n520 VSUBS 0.007777f
C776 B.n521 VSUBS 0.007777f
C777 B.n522 VSUBS 0.007777f
C778 B.n523 VSUBS 0.007777f
C779 B.n524 VSUBS 0.007777f
C780 B.n525 VSUBS 0.007777f
C781 B.n526 VSUBS 0.007777f
C782 B.n527 VSUBS 0.007777f
C783 B.n528 VSUBS 0.007777f
C784 B.n529 VSUBS 0.007777f
C785 B.n530 VSUBS 0.007777f
C786 B.n531 VSUBS 0.007777f
C787 B.n532 VSUBS 0.007777f
C788 B.n533 VSUBS 0.007777f
C789 B.n534 VSUBS 0.007777f
C790 B.n535 VSUBS 0.007777f
C791 B.n536 VSUBS 0.007777f
C792 B.n537 VSUBS 0.007777f
C793 B.n538 VSUBS 0.007777f
C794 B.n539 VSUBS 0.007777f
C795 B.n540 VSUBS 0.007777f
C796 B.n541 VSUBS 0.007777f
C797 B.n542 VSUBS 0.007777f
C798 B.n543 VSUBS 0.007777f
C799 B.n544 VSUBS 0.007777f
C800 B.n545 VSUBS 0.007777f
C801 B.n546 VSUBS 0.007777f
C802 B.n547 VSUBS 0.007777f
C803 B.n548 VSUBS 0.007777f
C804 B.n549 VSUBS 0.007777f
C805 B.n550 VSUBS 0.007777f
C806 B.n551 VSUBS 0.007777f
C807 B.n552 VSUBS 0.007777f
C808 B.n553 VSUBS 0.007777f
C809 B.n554 VSUBS 0.007777f
C810 B.n555 VSUBS 0.007777f
C811 B.n556 VSUBS 0.007777f
C812 B.n557 VSUBS 0.007777f
C813 B.n558 VSUBS 0.007777f
C814 B.n559 VSUBS 0.007777f
C815 B.n560 VSUBS 0.007777f
C816 B.n561 VSUBS 0.007777f
C817 B.n562 VSUBS 0.007777f
C818 B.n563 VSUBS 0.007777f
C819 B.n564 VSUBS 0.007777f
C820 B.n565 VSUBS 0.007777f
C821 B.n566 VSUBS 0.007777f
C822 B.n567 VSUBS 0.007777f
C823 B.n568 VSUBS 0.007777f
C824 B.n569 VSUBS 0.005376f
C825 B.n570 VSUBS 0.018019f
C826 B.n571 VSUBS 0.006291f
C827 B.n572 VSUBS 0.007777f
C828 B.n573 VSUBS 0.007777f
C829 B.n574 VSUBS 0.007777f
C830 B.n575 VSUBS 0.007777f
C831 B.n576 VSUBS 0.007777f
C832 B.n577 VSUBS 0.007777f
C833 B.n578 VSUBS 0.007777f
C834 B.n579 VSUBS 0.007777f
C835 B.n580 VSUBS 0.007777f
C836 B.n581 VSUBS 0.007777f
C837 B.n582 VSUBS 0.007777f
C838 B.n583 VSUBS 0.006291f
C839 B.n584 VSUBS 0.018019f
C840 B.n585 VSUBS 0.005376f
C841 B.n586 VSUBS 0.007777f
C842 B.n587 VSUBS 0.007777f
C843 B.n588 VSUBS 0.007777f
C844 B.n589 VSUBS 0.007777f
C845 B.n590 VSUBS 0.007777f
C846 B.n591 VSUBS 0.007777f
C847 B.n592 VSUBS 0.007777f
C848 B.n593 VSUBS 0.007777f
C849 B.n594 VSUBS 0.007777f
C850 B.n595 VSUBS 0.007777f
C851 B.n596 VSUBS 0.007777f
C852 B.n597 VSUBS 0.007777f
C853 B.n598 VSUBS 0.007777f
C854 B.n599 VSUBS 0.007777f
C855 B.n600 VSUBS 0.007777f
C856 B.n601 VSUBS 0.007777f
C857 B.n602 VSUBS 0.007777f
C858 B.n603 VSUBS 0.007777f
C859 B.n604 VSUBS 0.007777f
C860 B.n605 VSUBS 0.007777f
C861 B.n606 VSUBS 0.007777f
C862 B.n607 VSUBS 0.007777f
C863 B.n608 VSUBS 0.007777f
C864 B.n609 VSUBS 0.007777f
C865 B.n610 VSUBS 0.007777f
C866 B.n611 VSUBS 0.007777f
C867 B.n612 VSUBS 0.007777f
C868 B.n613 VSUBS 0.007777f
C869 B.n614 VSUBS 0.007777f
C870 B.n615 VSUBS 0.007777f
C871 B.n616 VSUBS 0.007777f
C872 B.n617 VSUBS 0.007777f
C873 B.n618 VSUBS 0.007777f
C874 B.n619 VSUBS 0.007777f
C875 B.n620 VSUBS 0.007777f
C876 B.n621 VSUBS 0.007777f
C877 B.n622 VSUBS 0.007777f
C878 B.n623 VSUBS 0.007777f
C879 B.n624 VSUBS 0.007777f
C880 B.n625 VSUBS 0.007777f
C881 B.n626 VSUBS 0.007777f
C882 B.n627 VSUBS 0.007777f
C883 B.n628 VSUBS 0.007777f
C884 B.n629 VSUBS 0.007777f
C885 B.n630 VSUBS 0.007777f
C886 B.n631 VSUBS 0.007777f
C887 B.n632 VSUBS 0.007777f
C888 B.n633 VSUBS 0.007777f
C889 B.n634 VSUBS 0.007777f
C890 B.n635 VSUBS 0.007777f
C891 B.n636 VSUBS 0.007777f
C892 B.n637 VSUBS 0.007777f
C893 B.n638 VSUBS 0.007777f
C894 B.n639 VSUBS 0.007777f
C895 B.n640 VSUBS 0.007777f
C896 B.n641 VSUBS 0.007777f
C897 B.n642 VSUBS 0.007777f
C898 B.n643 VSUBS 0.007777f
C899 B.n644 VSUBS 0.007777f
C900 B.n645 VSUBS 0.007777f
C901 B.n646 VSUBS 0.007777f
C902 B.n647 VSUBS 0.007777f
C903 B.n648 VSUBS 0.007777f
C904 B.n649 VSUBS 0.007777f
C905 B.n650 VSUBS 0.007777f
C906 B.n651 VSUBS 0.007777f
C907 B.n652 VSUBS 0.007777f
C908 B.n653 VSUBS 0.007777f
C909 B.n654 VSUBS 0.007777f
C910 B.n655 VSUBS 0.007777f
C911 B.n656 VSUBS 0.007777f
C912 B.n657 VSUBS 0.007777f
C913 B.n658 VSUBS 0.007777f
C914 B.n659 VSUBS 0.007777f
C915 B.n660 VSUBS 0.007777f
C916 B.n661 VSUBS 0.007777f
C917 B.n662 VSUBS 0.007777f
C918 B.n663 VSUBS 0.007777f
C919 B.n664 VSUBS 0.007777f
C920 B.n665 VSUBS 0.007777f
C921 B.n666 VSUBS 0.007777f
C922 B.n667 VSUBS 0.007777f
C923 B.n668 VSUBS 0.007777f
C924 B.n669 VSUBS 0.007777f
C925 B.n670 VSUBS 0.007777f
C926 B.n671 VSUBS 0.007777f
C927 B.n672 VSUBS 0.007777f
C928 B.n673 VSUBS 0.007777f
C929 B.n674 VSUBS 0.007777f
C930 B.n675 VSUBS 0.007777f
C931 B.n676 VSUBS 0.007777f
C932 B.n677 VSUBS 0.007777f
C933 B.n678 VSUBS 0.007777f
C934 B.n679 VSUBS 0.007777f
C935 B.n680 VSUBS 0.018035f
C936 B.n681 VSUBS 0.016964f
C937 B.n682 VSUBS 0.016964f
C938 B.n683 VSUBS 0.007777f
C939 B.n684 VSUBS 0.007777f
C940 B.n685 VSUBS 0.007777f
C941 B.n686 VSUBS 0.007777f
C942 B.n687 VSUBS 0.007777f
C943 B.n688 VSUBS 0.007777f
C944 B.n689 VSUBS 0.007777f
C945 B.n690 VSUBS 0.007777f
C946 B.n691 VSUBS 0.007777f
C947 B.n692 VSUBS 0.007777f
C948 B.n693 VSUBS 0.007777f
C949 B.n694 VSUBS 0.007777f
C950 B.n695 VSUBS 0.007777f
C951 B.n696 VSUBS 0.007777f
C952 B.n697 VSUBS 0.007777f
C953 B.n698 VSUBS 0.007777f
C954 B.n699 VSUBS 0.007777f
C955 B.n700 VSUBS 0.007777f
C956 B.n701 VSUBS 0.007777f
C957 B.n702 VSUBS 0.007777f
C958 B.n703 VSUBS 0.007777f
C959 B.n704 VSUBS 0.007777f
C960 B.n705 VSUBS 0.007777f
C961 B.n706 VSUBS 0.007777f
C962 B.n707 VSUBS 0.010149f
C963 B.n708 VSUBS 0.010811f
C964 B.n709 VSUBS 0.021499f
C965 VDD1.n0 VSUBS 0.029721f
C966 VDD1.n1 VSUBS 0.027614f
C967 VDD1.n2 VSUBS 0.014838f
C968 VDD1.n3 VSUBS 0.035073f
C969 VDD1.n4 VSUBS 0.015711f
C970 VDD1.n5 VSUBS 0.027614f
C971 VDD1.n6 VSUBS 0.014838f
C972 VDD1.n7 VSUBS 0.035073f
C973 VDD1.n8 VSUBS 0.015711f
C974 VDD1.n9 VSUBS 0.027614f
C975 VDD1.n10 VSUBS 0.014838f
C976 VDD1.n11 VSUBS 0.035073f
C977 VDD1.n12 VSUBS 0.015711f
C978 VDD1.n13 VSUBS 0.027614f
C979 VDD1.n14 VSUBS 0.014838f
C980 VDD1.n15 VSUBS 0.035073f
C981 VDD1.n16 VSUBS 0.015711f
C982 VDD1.n17 VSUBS 0.027614f
C983 VDD1.n18 VSUBS 0.014838f
C984 VDD1.n19 VSUBS 0.035073f
C985 VDD1.n20 VSUBS 0.015711f
C986 VDD1.n21 VSUBS 0.027614f
C987 VDD1.n22 VSUBS 0.014838f
C988 VDD1.n23 VSUBS 0.035073f
C989 VDD1.n24 VSUBS 0.015711f
C990 VDD1.n25 VSUBS 0.027614f
C991 VDD1.n26 VSUBS 0.014838f
C992 VDD1.n27 VSUBS 0.035073f
C993 VDD1.n28 VSUBS 0.035073f
C994 VDD1.n29 VSUBS 0.015711f
C995 VDD1.n30 VSUBS 0.027614f
C996 VDD1.n31 VSUBS 0.014838f
C997 VDD1.n32 VSUBS 0.035073f
C998 VDD1.n33 VSUBS 0.015711f
C999 VDD1.n34 VSUBS 0.310743f
C1000 VDD1.t1 VSUBS 0.076275f
C1001 VDD1.n35 VSUBS 0.026305f
C1002 VDD1.n36 VSUBS 0.026384f
C1003 VDD1.n37 VSUBS 0.014838f
C1004 VDD1.n38 VSUBS 2.26057f
C1005 VDD1.n39 VSUBS 0.027614f
C1006 VDD1.n40 VSUBS 0.014838f
C1007 VDD1.n41 VSUBS 0.015711f
C1008 VDD1.n42 VSUBS 0.035073f
C1009 VDD1.n43 VSUBS 0.035073f
C1010 VDD1.n44 VSUBS 0.015711f
C1011 VDD1.n45 VSUBS 0.014838f
C1012 VDD1.n46 VSUBS 0.027614f
C1013 VDD1.n47 VSUBS 0.027614f
C1014 VDD1.n48 VSUBS 0.014838f
C1015 VDD1.n49 VSUBS 0.015711f
C1016 VDD1.n50 VSUBS 0.035073f
C1017 VDD1.n51 VSUBS 0.035073f
C1018 VDD1.n52 VSUBS 0.015711f
C1019 VDD1.n53 VSUBS 0.014838f
C1020 VDD1.n54 VSUBS 0.027614f
C1021 VDD1.n55 VSUBS 0.027614f
C1022 VDD1.n56 VSUBS 0.014838f
C1023 VDD1.n57 VSUBS 0.015275f
C1024 VDD1.n58 VSUBS 0.015275f
C1025 VDD1.n59 VSUBS 0.035073f
C1026 VDD1.n60 VSUBS 0.035073f
C1027 VDD1.n61 VSUBS 0.015711f
C1028 VDD1.n62 VSUBS 0.014838f
C1029 VDD1.n63 VSUBS 0.027614f
C1030 VDD1.n64 VSUBS 0.027614f
C1031 VDD1.n65 VSUBS 0.014838f
C1032 VDD1.n66 VSUBS 0.015711f
C1033 VDD1.n67 VSUBS 0.035073f
C1034 VDD1.n68 VSUBS 0.035073f
C1035 VDD1.n69 VSUBS 0.015711f
C1036 VDD1.n70 VSUBS 0.014838f
C1037 VDD1.n71 VSUBS 0.027614f
C1038 VDD1.n72 VSUBS 0.027614f
C1039 VDD1.n73 VSUBS 0.014838f
C1040 VDD1.n74 VSUBS 0.015711f
C1041 VDD1.n75 VSUBS 0.035073f
C1042 VDD1.n76 VSUBS 0.035073f
C1043 VDD1.n77 VSUBS 0.015711f
C1044 VDD1.n78 VSUBS 0.014838f
C1045 VDD1.n79 VSUBS 0.027614f
C1046 VDD1.n80 VSUBS 0.027614f
C1047 VDD1.n81 VSUBS 0.014838f
C1048 VDD1.n82 VSUBS 0.015711f
C1049 VDD1.n83 VSUBS 0.035073f
C1050 VDD1.n84 VSUBS 0.035073f
C1051 VDD1.n85 VSUBS 0.015711f
C1052 VDD1.n86 VSUBS 0.014838f
C1053 VDD1.n87 VSUBS 0.027614f
C1054 VDD1.n88 VSUBS 0.027614f
C1055 VDD1.n89 VSUBS 0.014838f
C1056 VDD1.n90 VSUBS 0.015711f
C1057 VDD1.n91 VSUBS 0.035073f
C1058 VDD1.n92 VSUBS 0.035073f
C1059 VDD1.n93 VSUBS 0.015711f
C1060 VDD1.n94 VSUBS 0.014838f
C1061 VDD1.n95 VSUBS 0.027614f
C1062 VDD1.n96 VSUBS 0.027614f
C1063 VDD1.n97 VSUBS 0.014838f
C1064 VDD1.n98 VSUBS 0.015711f
C1065 VDD1.n99 VSUBS 0.035073f
C1066 VDD1.n100 VSUBS 0.087071f
C1067 VDD1.n101 VSUBS 0.015711f
C1068 VDD1.n102 VSUBS 0.029139f
C1069 VDD1.n103 VSUBS 0.069486f
C1070 VDD1.n104 VSUBS 0.086493f
C1071 VDD1.n105 VSUBS 0.029721f
C1072 VDD1.n106 VSUBS 0.027614f
C1073 VDD1.n107 VSUBS 0.014838f
C1074 VDD1.n108 VSUBS 0.035073f
C1075 VDD1.n109 VSUBS 0.015711f
C1076 VDD1.n110 VSUBS 0.027614f
C1077 VDD1.n111 VSUBS 0.014838f
C1078 VDD1.n112 VSUBS 0.035073f
C1079 VDD1.n113 VSUBS 0.015711f
C1080 VDD1.n114 VSUBS 0.027614f
C1081 VDD1.n115 VSUBS 0.014838f
C1082 VDD1.n116 VSUBS 0.035073f
C1083 VDD1.n117 VSUBS 0.015711f
C1084 VDD1.n118 VSUBS 0.027614f
C1085 VDD1.n119 VSUBS 0.014838f
C1086 VDD1.n120 VSUBS 0.035073f
C1087 VDD1.n121 VSUBS 0.015711f
C1088 VDD1.n122 VSUBS 0.027614f
C1089 VDD1.n123 VSUBS 0.014838f
C1090 VDD1.n124 VSUBS 0.035073f
C1091 VDD1.n125 VSUBS 0.015711f
C1092 VDD1.n126 VSUBS 0.027614f
C1093 VDD1.n127 VSUBS 0.014838f
C1094 VDD1.n128 VSUBS 0.035073f
C1095 VDD1.n129 VSUBS 0.015711f
C1096 VDD1.n130 VSUBS 0.027614f
C1097 VDD1.n131 VSUBS 0.014838f
C1098 VDD1.n132 VSUBS 0.035073f
C1099 VDD1.n133 VSUBS 0.015711f
C1100 VDD1.n134 VSUBS 0.027614f
C1101 VDD1.n135 VSUBS 0.014838f
C1102 VDD1.n136 VSUBS 0.035073f
C1103 VDD1.n137 VSUBS 0.015711f
C1104 VDD1.n138 VSUBS 0.310743f
C1105 VDD1.t0 VSUBS 0.076275f
C1106 VDD1.n139 VSUBS 0.026305f
C1107 VDD1.n140 VSUBS 0.026384f
C1108 VDD1.n141 VSUBS 0.014838f
C1109 VDD1.n142 VSUBS 2.26057f
C1110 VDD1.n143 VSUBS 0.027614f
C1111 VDD1.n144 VSUBS 0.014838f
C1112 VDD1.n145 VSUBS 0.015711f
C1113 VDD1.n146 VSUBS 0.035073f
C1114 VDD1.n147 VSUBS 0.035073f
C1115 VDD1.n148 VSUBS 0.015711f
C1116 VDD1.n149 VSUBS 0.014838f
C1117 VDD1.n150 VSUBS 0.027614f
C1118 VDD1.n151 VSUBS 0.027614f
C1119 VDD1.n152 VSUBS 0.014838f
C1120 VDD1.n153 VSUBS 0.015711f
C1121 VDD1.n154 VSUBS 0.035073f
C1122 VDD1.n155 VSUBS 0.035073f
C1123 VDD1.n156 VSUBS 0.035073f
C1124 VDD1.n157 VSUBS 0.015711f
C1125 VDD1.n158 VSUBS 0.014838f
C1126 VDD1.n159 VSUBS 0.027614f
C1127 VDD1.n160 VSUBS 0.027614f
C1128 VDD1.n161 VSUBS 0.014838f
C1129 VDD1.n162 VSUBS 0.015275f
C1130 VDD1.n163 VSUBS 0.015275f
C1131 VDD1.n164 VSUBS 0.035073f
C1132 VDD1.n165 VSUBS 0.035073f
C1133 VDD1.n166 VSUBS 0.015711f
C1134 VDD1.n167 VSUBS 0.014838f
C1135 VDD1.n168 VSUBS 0.027614f
C1136 VDD1.n169 VSUBS 0.027614f
C1137 VDD1.n170 VSUBS 0.014838f
C1138 VDD1.n171 VSUBS 0.015711f
C1139 VDD1.n172 VSUBS 0.035073f
C1140 VDD1.n173 VSUBS 0.035073f
C1141 VDD1.n174 VSUBS 0.015711f
C1142 VDD1.n175 VSUBS 0.014838f
C1143 VDD1.n176 VSUBS 0.027614f
C1144 VDD1.n177 VSUBS 0.027614f
C1145 VDD1.n178 VSUBS 0.014838f
C1146 VDD1.n179 VSUBS 0.015711f
C1147 VDD1.n180 VSUBS 0.035073f
C1148 VDD1.n181 VSUBS 0.035073f
C1149 VDD1.n182 VSUBS 0.015711f
C1150 VDD1.n183 VSUBS 0.014838f
C1151 VDD1.n184 VSUBS 0.027614f
C1152 VDD1.n185 VSUBS 0.027614f
C1153 VDD1.n186 VSUBS 0.014838f
C1154 VDD1.n187 VSUBS 0.015711f
C1155 VDD1.n188 VSUBS 0.035073f
C1156 VDD1.n189 VSUBS 0.035073f
C1157 VDD1.n190 VSUBS 0.015711f
C1158 VDD1.n191 VSUBS 0.014838f
C1159 VDD1.n192 VSUBS 0.027614f
C1160 VDD1.n193 VSUBS 0.027614f
C1161 VDD1.n194 VSUBS 0.014838f
C1162 VDD1.n195 VSUBS 0.015711f
C1163 VDD1.n196 VSUBS 0.035073f
C1164 VDD1.n197 VSUBS 0.035073f
C1165 VDD1.n198 VSUBS 0.015711f
C1166 VDD1.n199 VSUBS 0.014838f
C1167 VDD1.n200 VSUBS 0.027614f
C1168 VDD1.n201 VSUBS 0.027614f
C1169 VDD1.n202 VSUBS 0.014838f
C1170 VDD1.n203 VSUBS 0.015711f
C1171 VDD1.n204 VSUBS 0.035073f
C1172 VDD1.n205 VSUBS 0.087071f
C1173 VDD1.n206 VSUBS 0.015711f
C1174 VDD1.n207 VSUBS 0.029139f
C1175 VDD1.n208 VSUBS 0.069486f
C1176 VDD1.n209 VSUBS 1.07401f
C1177 VTAIL.n0 VSUBS 0.029462f
C1178 VTAIL.n1 VSUBS 0.027374f
C1179 VTAIL.n2 VSUBS 0.01471f
C1180 VTAIL.n3 VSUBS 0.034768f
C1181 VTAIL.n4 VSUBS 0.015575f
C1182 VTAIL.n5 VSUBS 0.027374f
C1183 VTAIL.n6 VSUBS 0.01471f
C1184 VTAIL.n7 VSUBS 0.034768f
C1185 VTAIL.n8 VSUBS 0.015575f
C1186 VTAIL.n9 VSUBS 0.027374f
C1187 VTAIL.n10 VSUBS 0.01471f
C1188 VTAIL.n11 VSUBS 0.034768f
C1189 VTAIL.n12 VSUBS 0.015575f
C1190 VTAIL.n13 VSUBS 0.027374f
C1191 VTAIL.n14 VSUBS 0.01471f
C1192 VTAIL.n15 VSUBS 0.034768f
C1193 VTAIL.n16 VSUBS 0.015575f
C1194 VTAIL.n17 VSUBS 0.027374f
C1195 VTAIL.n18 VSUBS 0.01471f
C1196 VTAIL.n19 VSUBS 0.034768f
C1197 VTAIL.n20 VSUBS 0.015575f
C1198 VTAIL.n21 VSUBS 0.027374f
C1199 VTAIL.n22 VSUBS 0.01471f
C1200 VTAIL.n23 VSUBS 0.034768f
C1201 VTAIL.n24 VSUBS 0.015575f
C1202 VTAIL.n25 VSUBS 0.027374f
C1203 VTAIL.n26 VSUBS 0.01471f
C1204 VTAIL.n27 VSUBS 0.034768f
C1205 VTAIL.n28 VSUBS 0.015575f
C1206 VTAIL.n29 VSUBS 0.027374f
C1207 VTAIL.n30 VSUBS 0.01471f
C1208 VTAIL.n31 VSUBS 0.034768f
C1209 VTAIL.n32 VSUBS 0.015575f
C1210 VTAIL.n33 VSUBS 0.308045f
C1211 VTAIL.t3 VSUBS 0.075612f
C1212 VTAIL.n34 VSUBS 0.026076f
C1213 VTAIL.n35 VSUBS 0.026154f
C1214 VTAIL.n36 VSUBS 0.01471f
C1215 VTAIL.n37 VSUBS 2.24094f
C1216 VTAIL.n38 VSUBS 0.027374f
C1217 VTAIL.n39 VSUBS 0.01471f
C1218 VTAIL.n40 VSUBS 0.015575f
C1219 VTAIL.n41 VSUBS 0.034768f
C1220 VTAIL.n42 VSUBS 0.034768f
C1221 VTAIL.n43 VSUBS 0.015575f
C1222 VTAIL.n44 VSUBS 0.01471f
C1223 VTAIL.n45 VSUBS 0.027374f
C1224 VTAIL.n46 VSUBS 0.027374f
C1225 VTAIL.n47 VSUBS 0.01471f
C1226 VTAIL.n48 VSUBS 0.015575f
C1227 VTAIL.n49 VSUBS 0.034768f
C1228 VTAIL.n50 VSUBS 0.034768f
C1229 VTAIL.n51 VSUBS 0.034768f
C1230 VTAIL.n52 VSUBS 0.015575f
C1231 VTAIL.n53 VSUBS 0.01471f
C1232 VTAIL.n54 VSUBS 0.027374f
C1233 VTAIL.n55 VSUBS 0.027374f
C1234 VTAIL.n56 VSUBS 0.01471f
C1235 VTAIL.n57 VSUBS 0.015142f
C1236 VTAIL.n58 VSUBS 0.015142f
C1237 VTAIL.n59 VSUBS 0.034768f
C1238 VTAIL.n60 VSUBS 0.034768f
C1239 VTAIL.n61 VSUBS 0.015575f
C1240 VTAIL.n62 VSUBS 0.01471f
C1241 VTAIL.n63 VSUBS 0.027374f
C1242 VTAIL.n64 VSUBS 0.027374f
C1243 VTAIL.n65 VSUBS 0.01471f
C1244 VTAIL.n66 VSUBS 0.015575f
C1245 VTAIL.n67 VSUBS 0.034768f
C1246 VTAIL.n68 VSUBS 0.034768f
C1247 VTAIL.n69 VSUBS 0.015575f
C1248 VTAIL.n70 VSUBS 0.01471f
C1249 VTAIL.n71 VSUBS 0.027374f
C1250 VTAIL.n72 VSUBS 0.027374f
C1251 VTAIL.n73 VSUBS 0.01471f
C1252 VTAIL.n74 VSUBS 0.015575f
C1253 VTAIL.n75 VSUBS 0.034768f
C1254 VTAIL.n76 VSUBS 0.034768f
C1255 VTAIL.n77 VSUBS 0.015575f
C1256 VTAIL.n78 VSUBS 0.01471f
C1257 VTAIL.n79 VSUBS 0.027374f
C1258 VTAIL.n80 VSUBS 0.027374f
C1259 VTAIL.n81 VSUBS 0.01471f
C1260 VTAIL.n82 VSUBS 0.015575f
C1261 VTAIL.n83 VSUBS 0.034768f
C1262 VTAIL.n84 VSUBS 0.034768f
C1263 VTAIL.n85 VSUBS 0.015575f
C1264 VTAIL.n86 VSUBS 0.01471f
C1265 VTAIL.n87 VSUBS 0.027374f
C1266 VTAIL.n88 VSUBS 0.027374f
C1267 VTAIL.n89 VSUBS 0.01471f
C1268 VTAIL.n90 VSUBS 0.015575f
C1269 VTAIL.n91 VSUBS 0.034768f
C1270 VTAIL.n92 VSUBS 0.034768f
C1271 VTAIL.n93 VSUBS 0.015575f
C1272 VTAIL.n94 VSUBS 0.01471f
C1273 VTAIL.n95 VSUBS 0.027374f
C1274 VTAIL.n96 VSUBS 0.027374f
C1275 VTAIL.n97 VSUBS 0.01471f
C1276 VTAIL.n98 VSUBS 0.015575f
C1277 VTAIL.n99 VSUBS 0.034768f
C1278 VTAIL.n100 VSUBS 0.086314f
C1279 VTAIL.n101 VSUBS 0.015575f
C1280 VTAIL.n102 VSUBS 0.028886f
C1281 VTAIL.n103 VSUBS 0.068883f
C1282 VTAIL.n104 VSUBS 0.066089f
C1283 VTAIL.n105 VSUBS 2.22656f
C1284 VTAIL.n106 VSUBS 0.029462f
C1285 VTAIL.n107 VSUBS 0.027374f
C1286 VTAIL.n108 VSUBS 0.01471f
C1287 VTAIL.n109 VSUBS 0.034768f
C1288 VTAIL.n110 VSUBS 0.015575f
C1289 VTAIL.n111 VSUBS 0.027374f
C1290 VTAIL.n112 VSUBS 0.01471f
C1291 VTAIL.n113 VSUBS 0.034768f
C1292 VTAIL.n114 VSUBS 0.015575f
C1293 VTAIL.n115 VSUBS 0.027374f
C1294 VTAIL.n116 VSUBS 0.01471f
C1295 VTAIL.n117 VSUBS 0.034768f
C1296 VTAIL.n118 VSUBS 0.015575f
C1297 VTAIL.n119 VSUBS 0.027374f
C1298 VTAIL.n120 VSUBS 0.01471f
C1299 VTAIL.n121 VSUBS 0.034768f
C1300 VTAIL.n122 VSUBS 0.015575f
C1301 VTAIL.n123 VSUBS 0.027374f
C1302 VTAIL.n124 VSUBS 0.01471f
C1303 VTAIL.n125 VSUBS 0.034768f
C1304 VTAIL.n126 VSUBS 0.015575f
C1305 VTAIL.n127 VSUBS 0.027374f
C1306 VTAIL.n128 VSUBS 0.01471f
C1307 VTAIL.n129 VSUBS 0.034768f
C1308 VTAIL.n130 VSUBS 0.015575f
C1309 VTAIL.n131 VSUBS 0.027374f
C1310 VTAIL.n132 VSUBS 0.01471f
C1311 VTAIL.n133 VSUBS 0.034768f
C1312 VTAIL.n134 VSUBS 0.034768f
C1313 VTAIL.n135 VSUBS 0.015575f
C1314 VTAIL.n136 VSUBS 0.027374f
C1315 VTAIL.n137 VSUBS 0.01471f
C1316 VTAIL.n138 VSUBS 0.034768f
C1317 VTAIL.n139 VSUBS 0.015575f
C1318 VTAIL.n140 VSUBS 0.308044f
C1319 VTAIL.t0 VSUBS 0.075612f
C1320 VTAIL.n141 VSUBS 0.026076f
C1321 VTAIL.n142 VSUBS 0.026154f
C1322 VTAIL.n143 VSUBS 0.01471f
C1323 VTAIL.n144 VSUBS 2.24094f
C1324 VTAIL.n145 VSUBS 0.027374f
C1325 VTAIL.n146 VSUBS 0.01471f
C1326 VTAIL.n147 VSUBS 0.015575f
C1327 VTAIL.n148 VSUBS 0.034768f
C1328 VTAIL.n149 VSUBS 0.034768f
C1329 VTAIL.n150 VSUBS 0.015575f
C1330 VTAIL.n151 VSUBS 0.01471f
C1331 VTAIL.n152 VSUBS 0.027374f
C1332 VTAIL.n153 VSUBS 0.027374f
C1333 VTAIL.n154 VSUBS 0.01471f
C1334 VTAIL.n155 VSUBS 0.015575f
C1335 VTAIL.n156 VSUBS 0.034768f
C1336 VTAIL.n157 VSUBS 0.034768f
C1337 VTAIL.n158 VSUBS 0.015575f
C1338 VTAIL.n159 VSUBS 0.01471f
C1339 VTAIL.n160 VSUBS 0.027374f
C1340 VTAIL.n161 VSUBS 0.027374f
C1341 VTAIL.n162 VSUBS 0.01471f
C1342 VTAIL.n163 VSUBS 0.015142f
C1343 VTAIL.n164 VSUBS 0.015142f
C1344 VTAIL.n165 VSUBS 0.034768f
C1345 VTAIL.n166 VSUBS 0.034768f
C1346 VTAIL.n167 VSUBS 0.015575f
C1347 VTAIL.n168 VSUBS 0.01471f
C1348 VTAIL.n169 VSUBS 0.027374f
C1349 VTAIL.n170 VSUBS 0.027374f
C1350 VTAIL.n171 VSUBS 0.01471f
C1351 VTAIL.n172 VSUBS 0.015575f
C1352 VTAIL.n173 VSUBS 0.034768f
C1353 VTAIL.n174 VSUBS 0.034768f
C1354 VTAIL.n175 VSUBS 0.015575f
C1355 VTAIL.n176 VSUBS 0.01471f
C1356 VTAIL.n177 VSUBS 0.027374f
C1357 VTAIL.n178 VSUBS 0.027374f
C1358 VTAIL.n179 VSUBS 0.01471f
C1359 VTAIL.n180 VSUBS 0.015575f
C1360 VTAIL.n181 VSUBS 0.034768f
C1361 VTAIL.n182 VSUBS 0.034768f
C1362 VTAIL.n183 VSUBS 0.015575f
C1363 VTAIL.n184 VSUBS 0.01471f
C1364 VTAIL.n185 VSUBS 0.027374f
C1365 VTAIL.n186 VSUBS 0.027374f
C1366 VTAIL.n187 VSUBS 0.01471f
C1367 VTAIL.n188 VSUBS 0.015575f
C1368 VTAIL.n189 VSUBS 0.034768f
C1369 VTAIL.n190 VSUBS 0.034768f
C1370 VTAIL.n191 VSUBS 0.015575f
C1371 VTAIL.n192 VSUBS 0.01471f
C1372 VTAIL.n193 VSUBS 0.027374f
C1373 VTAIL.n194 VSUBS 0.027374f
C1374 VTAIL.n195 VSUBS 0.01471f
C1375 VTAIL.n196 VSUBS 0.015575f
C1376 VTAIL.n197 VSUBS 0.034768f
C1377 VTAIL.n198 VSUBS 0.034768f
C1378 VTAIL.n199 VSUBS 0.015575f
C1379 VTAIL.n200 VSUBS 0.01471f
C1380 VTAIL.n201 VSUBS 0.027374f
C1381 VTAIL.n202 VSUBS 0.027374f
C1382 VTAIL.n203 VSUBS 0.01471f
C1383 VTAIL.n204 VSUBS 0.015575f
C1384 VTAIL.n205 VSUBS 0.034768f
C1385 VTAIL.n206 VSUBS 0.086314f
C1386 VTAIL.n207 VSUBS 0.015575f
C1387 VTAIL.n208 VSUBS 0.028886f
C1388 VTAIL.n209 VSUBS 0.068883f
C1389 VTAIL.n210 VSUBS 0.066089f
C1390 VTAIL.n211 VSUBS 2.25488f
C1391 VTAIL.n212 VSUBS 0.029462f
C1392 VTAIL.n213 VSUBS 0.027374f
C1393 VTAIL.n214 VSUBS 0.01471f
C1394 VTAIL.n215 VSUBS 0.034768f
C1395 VTAIL.n216 VSUBS 0.015575f
C1396 VTAIL.n217 VSUBS 0.027374f
C1397 VTAIL.n218 VSUBS 0.01471f
C1398 VTAIL.n219 VSUBS 0.034768f
C1399 VTAIL.n220 VSUBS 0.015575f
C1400 VTAIL.n221 VSUBS 0.027374f
C1401 VTAIL.n222 VSUBS 0.01471f
C1402 VTAIL.n223 VSUBS 0.034768f
C1403 VTAIL.n224 VSUBS 0.015575f
C1404 VTAIL.n225 VSUBS 0.027374f
C1405 VTAIL.n226 VSUBS 0.01471f
C1406 VTAIL.n227 VSUBS 0.034768f
C1407 VTAIL.n228 VSUBS 0.015575f
C1408 VTAIL.n229 VSUBS 0.027374f
C1409 VTAIL.n230 VSUBS 0.01471f
C1410 VTAIL.n231 VSUBS 0.034768f
C1411 VTAIL.n232 VSUBS 0.015575f
C1412 VTAIL.n233 VSUBS 0.027374f
C1413 VTAIL.n234 VSUBS 0.01471f
C1414 VTAIL.n235 VSUBS 0.034768f
C1415 VTAIL.n236 VSUBS 0.015575f
C1416 VTAIL.n237 VSUBS 0.027374f
C1417 VTAIL.n238 VSUBS 0.01471f
C1418 VTAIL.n239 VSUBS 0.034768f
C1419 VTAIL.n240 VSUBS 0.034768f
C1420 VTAIL.n241 VSUBS 0.015575f
C1421 VTAIL.n242 VSUBS 0.027374f
C1422 VTAIL.n243 VSUBS 0.01471f
C1423 VTAIL.n244 VSUBS 0.034768f
C1424 VTAIL.n245 VSUBS 0.015575f
C1425 VTAIL.n246 VSUBS 0.308044f
C1426 VTAIL.t2 VSUBS 0.075612f
C1427 VTAIL.n247 VSUBS 0.026076f
C1428 VTAIL.n248 VSUBS 0.026154f
C1429 VTAIL.n249 VSUBS 0.01471f
C1430 VTAIL.n250 VSUBS 2.24094f
C1431 VTAIL.n251 VSUBS 0.027374f
C1432 VTAIL.n252 VSUBS 0.01471f
C1433 VTAIL.n253 VSUBS 0.015575f
C1434 VTAIL.n254 VSUBS 0.034768f
C1435 VTAIL.n255 VSUBS 0.034768f
C1436 VTAIL.n256 VSUBS 0.015575f
C1437 VTAIL.n257 VSUBS 0.01471f
C1438 VTAIL.n258 VSUBS 0.027374f
C1439 VTAIL.n259 VSUBS 0.027374f
C1440 VTAIL.n260 VSUBS 0.01471f
C1441 VTAIL.n261 VSUBS 0.015575f
C1442 VTAIL.n262 VSUBS 0.034768f
C1443 VTAIL.n263 VSUBS 0.034768f
C1444 VTAIL.n264 VSUBS 0.015575f
C1445 VTAIL.n265 VSUBS 0.01471f
C1446 VTAIL.n266 VSUBS 0.027374f
C1447 VTAIL.n267 VSUBS 0.027374f
C1448 VTAIL.n268 VSUBS 0.01471f
C1449 VTAIL.n269 VSUBS 0.015142f
C1450 VTAIL.n270 VSUBS 0.015142f
C1451 VTAIL.n271 VSUBS 0.034768f
C1452 VTAIL.n272 VSUBS 0.034768f
C1453 VTAIL.n273 VSUBS 0.015575f
C1454 VTAIL.n274 VSUBS 0.01471f
C1455 VTAIL.n275 VSUBS 0.027374f
C1456 VTAIL.n276 VSUBS 0.027374f
C1457 VTAIL.n277 VSUBS 0.01471f
C1458 VTAIL.n278 VSUBS 0.015575f
C1459 VTAIL.n279 VSUBS 0.034768f
C1460 VTAIL.n280 VSUBS 0.034768f
C1461 VTAIL.n281 VSUBS 0.015575f
C1462 VTAIL.n282 VSUBS 0.01471f
C1463 VTAIL.n283 VSUBS 0.027374f
C1464 VTAIL.n284 VSUBS 0.027374f
C1465 VTAIL.n285 VSUBS 0.01471f
C1466 VTAIL.n286 VSUBS 0.015575f
C1467 VTAIL.n287 VSUBS 0.034768f
C1468 VTAIL.n288 VSUBS 0.034768f
C1469 VTAIL.n289 VSUBS 0.015575f
C1470 VTAIL.n290 VSUBS 0.01471f
C1471 VTAIL.n291 VSUBS 0.027374f
C1472 VTAIL.n292 VSUBS 0.027374f
C1473 VTAIL.n293 VSUBS 0.01471f
C1474 VTAIL.n294 VSUBS 0.015575f
C1475 VTAIL.n295 VSUBS 0.034768f
C1476 VTAIL.n296 VSUBS 0.034768f
C1477 VTAIL.n297 VSUBS 0.015575f
C1478 VTAIL.n298 VSUBS 0.01471f
C1479 VTAIL.n299 VSUBS 0.027374f
C1480 VTAIL.n300 VSUBS 0.027374f
C1481 VTAIL.n301 VSUBS 0.01471f
C1482 VTAIL.n302 VSUBS 0.015575f
C1483 VTAIL.n303 VSUBS 0.034768f
C1484 VTAIL.n304 VSUBS 0.034768f
C1485 VTAIL.n305 VSUBS 0.015575f
C1486 VTAIL.n306 VSUBS 0.01471f
C1487 VTAIL.n307 VSUBS 0.027374f
C1488 VTAIL.n308 VSUBS 0.027374f
C1489 VTAIL.n309 VSUBS 0.01471f
C1490 VTAIL.n310 VSUBS 0.015575f
C1491 VTAIL.n311 VSUBS 0.034768f
C1492 VTAIL.n312 VSUBS 0.086314f
C1493 VTAIL.n313 VSUBS 0.015575f
C1494 VTAIL.n314 VSUBS 0.028886f
C1495 VTAIL.n315 VSUBS 0.068883f
C1496 VTAIL.n316 VSUBS 0.066089f
C1497 VTAIL.n317 VSUBS 2.12105f
C1498 VTAIL.n318 VSUBS 0.029462f
C1499 VTAIL.n319 VSUBS 0.027374f
C1500 VTAIL.n320 VSUBS 0.01471f
C1501 VTAIL.n321 VSUBS 0.034768f
C1502 VTAIL.n322 VSUBS 0.015575f
C1503 VTAIL.n323 VSUBS 0.027374f
C1504 VTAIL.n324 VSUBS 0.01471f
C1505 VTAIL.n325 VSUBS 0.034768f
C1506 VTAIL.n326 VSUBS 0.015575f
C1507 VTAIL.n327 VSUBS 0.027374f
C1508 VTAIL.n328 VSUBS 0.01471f
C1509 VTAIL.n329 VSUBS 0.034768f
C1510 VTAIL.n330 VSUBS 0.015575f
C1511 VTAIL.n331 VSUBS 0.027374f
C1512 VTAIL.n332 VSUBS 0.01471f
C1513 VTAIL.n333 VSUBS 0.034768f
C1514 VTAIL.n334 VSUBS 0.015575f
C1515 VTAIL.n335 VSUBS 0.027374f
C1516 VTAIL.n336 VSUBS 0.01471f
C1517 VTAIL.n337 VSUBS 0.034768f
C1518 VTAIL.n338 VSUBS 0.015575f
C1519 VTAIL.n339 VSUBS 0.027374f
C1520 VTAIL.n340 VSUBS 0.01471f
C1521 VTAIL.n341 VSUBS 0.034768f
C1522 VTAIL.n342 VSUBS 0.015575f
C1523 VTAIL.n343 VSUBS 0.027374f
C1524 VTAIL.n344 VSUBS 0.01471f
C1525 VTAIL.n345 VSUBS 0.034768f
C1526 VTAIL.n346 VSUBS 0.015575f
C1527 VTAIL.n347 VSUBS 0.027374f
C1528 VTAIL.n348 VSUBS 0.01471f
C1529 VTAIL.n349 VSUBS 0.034768f
C1530 VTAIL.n350 VSUBS 0.015575f
C1531 VTAIL.n351 VSUBS 0.308045f
C1532 VTAIL.t1 VSUBS 0.075612f
C1533 VTAIL.n352 VSUBS 0.026076f
C1534 VTAIL.n353 VSUBS 0.026154f
C1535 VTAIL.n354 VSUBS 0.01471f
C1536 VTAIL.n355 VSUBS 2.24094f
C1537 VTAIL.n356 VSUBS 0.027374f
C1538 VTAIL.n357 VSUBS 0.01471f
C1539 VTAIL.n358 VSUBS 0.015575f
C1540 VTAIL.n359 VSUBS 0.034768f
C1541 VTAIL.n360 VSUBS 0.034768f
C1542 VTAIL.n361 VSUBS 0.015575f
C1543 VTAIL.n362 VSUBS 0.01471f
C1544 VTAIL.n363 VSUBS 0.027374f
C1545 VTAIL.n364 VSUBS 0.027374f
C1546 VTAIL.n365 VSUBS 0.01471f
C1547 VTAIL.n366 VSUBS 0.015575f
C1548 VTAIL.n367 VSUBS 0.034768f
C1549 VTAIL.n368 VSUBS 0.034768f
C1550 VTAIL.n369 VSUBS 0.034768f
C1551 VTAIL.n370 VSUBS 0.015575f
C1552 VTAIL.n371 VSUBS 0.01471f
C1553 VTAIL.n372 VSUBS 0.027374f
C1554 VTAIL.n373 VSUBS 0.027374f
C1555 VTAIL.n374 VSUBS 0.01471f
C1556 VTAIL.n375 VSUBS 0.015142f
C1557 VTAIL.n376 VSUBS 0.015142f
C1558 VTAIL.n377 VSUBS 0.034768f
C1559 VTAIL.n378 VSUBS 0.034768f
C1560 VTAIL.n379 VSUBS 0.015575f
C1561 VTAIL.n380 VSUBS 0.01471f
C1562 VTAIL.n381 VSUBS 0.027374f
C1563 VTAIL.n382 VSUBS 0.027374f
C1564 VTAIL.n383 VSUBS 0.01471f
C1565 VTAIL.n384 VSUBS 0.015575f
C1566 VTAIL.n385 VSUBS 0.034768f
C1567 VTAIL.n386 VSUBS 0.034768f
C1568 VTAIL.n387 VSUBS 0.015575f
C1569 VTAIL.n388 VSUBS 0.01471f
C1570 VTAIL.n389 VSUBS 0.027374f
C1571 VTAIL.n390 VSUBS 0.027374f
C1572 VTAIL.n391 VSUBS 0.01471f
C1573 VTAIL.n392 VSUBS 0.015575f
C1574 VTAIL.n393 VSUBS 0.034768f
C1575 VTAIL.n394 VSUBS 0.034768f
C1576 VTAIL.n395 VSUBS 0.015575f
C1577 VTAIL.n396 VSUBS 0.01471f
C1578 VTAIL.n397 VSUBS 0.027374f
C1579 VTAIL.n398 VSUBS 0.027374f
C1580 VTAIL.n399 VSUBS 0.01471f
C1581 VTAIL.n400 VSUBS 0.015575f
C1582 VTAIL.n401 VSUBS 0.034768f
C1583 VTAIL.n402 VSUBS 0.034768f
C1584 VTAIL.n403 VSUBS 0.015575f
C1585 VTAIL.n404 VSUBS 0.01471f
C1586 VTAIL.n405 VSUBS 0.027374f
C1587 VTAIL.n406 VSUBS 0.027374f
C1588 VTAIL.n407 VSUBS 0.01471f
C1589 VTAIL.n408 VSUBS 0.015575f
C1590 VTAIL.n409 VSUBS 0.034768f
C1591 VTAIL.n410 VSUBS 0.034768f
C1592 VTAIL.n411 VSUBS 0.015575f
C1593 VTAIL.n412 VSUBS 0.01471f
C1594 VTAIL.n413 VSUBS 0.027374f
C1595 VTAIL.n414 VSUBS 0.027374f
C1596 VTAIL.n415 VSUBS 0.01471f
C1597 VTAIL.n416 VSUBS 0.015575f
C1598 VTAIL.n417 VSUBS 0.034768f
C1599 VTAIL.n418 VSUBS 0.086314f
C1600 VTAIL.n419 VSUBS 0.015575f
C1601 VTAIL.n420 VSUBS 0.028886f
C1602 VTAIL.n421 VSUBS 0.068883f
C1603 VTAIL.n422 VSUBS 0.066089f
C1604 VTAIL.n423 VSUBS 2.04102f
C1605 VP.t0 VSUBS 4.60111f
C1606 VP.t1 VSUBS 4.23544f
C1607 VP.n0 VSUBS 7.11348f
.ends

