* NGSPICE file created from diff_pair_sample_1579.ext - technology: sky130A

.subckt diff_pair_sample_1579 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t14 VN.t0 VDD2.t1 w_n3350_n1784# sky130_fd_pr__pfet_01v8 ad=1.5912 pd=8.94 as=0.6732 ps=4.41 w=4.08 l=2.05
X1 B.t11 B.t9 B.t10 w_n3350_n1784# sky130_fd_pr__pfet_01v8 ad=1.5912 pd=8.94 as=0 ps=0 w=4.08 l=2.05
X2 B.t8 B.t6 B.t7 w_n3350_n1784# sky130_fd_pr__pfet_01v8 ad=1.5912 pd=8.94 as=0 ps=0 w=4.08 l=2.05
X3 VDD1.t7 VP.t0 VTAIL.t3 w_n3350_n1784# sky130_fd_pr__pfet_01v8 ad=0.6732 pd=4.41 as=0.6732 ps=4.41 w=4.08 l=2.05
X4 VTAIL.t13 VN.t1 VDD2.t0 w_n3350_n1784# sky130_fd_pr__pfet_01v8 ad=1.5912 pd=8.94 as=0.6732 ps=4.41 w=4.08 l=2.05
X5 VDD1.t6 VP.t1 VTAIL.t15 w_n3350_n1784# sky130_fd_pr__pfet_01v8 ad=0.6732 pd=4.41 as=1.5912 ps=8.94 w=4.08 l=2.05
X6 VDD2.t5 VN.t2 VTAIL.t12 w_n3350_n1784# sky130_fd_pr__pfet_01v8 ad=0.6732 pd=4.41 as=1.5912 ps=8.94 w=4.08 l=2.05
X7 VTAIL.t5 VP.t2 VDD1.t5 w_n3350_n1784# sky130_fd_pr__pfet_01v8 ad=0.6732 pd=4.41 as=0.6732 ps=4.41 w=4.08 l=2.05
X8 VDD2.t6 VN.t3 VTAIL.t11 w_n3350_n1784# sky130_fd_pr__pfet_01v8 ad=0.6732 pd=4.41 as=0.6732 ps=4.41 w=4.08 l=2.05
X9 VDD1.t4 VP.t3 VTAIL.t2 w_n3350_n1784# sky130_fd_pr__pfet_01v8 ad=0.6732 pd=4.41 as=1.5912 ps=8.94 w=4.08 l=2.05
X10 VDD1.t3 VP.t4 VTAIL.t1 w_n3350_n1784# sky130_fd_pr__pfet_01v8 ad=0.6732 pd=4.41 as=0.6732 ps=4.41 w=4.08 l=2.05
X11 VTAIL.t10 VN.t4 VDD2.t4 w_n3350_n1784# sky130_fd_pr__pfet_01v8 ad=0.6732 pd=4.41 as=0.6732 ps=4.41 w=4.08 l=2.05
X12 VTAIL.t9 VN.t5 VDD2.t3 w_n3350_n1784# sky130_fd_pr__pfet_01v8 ad=0.6732 pd=4.41 as=0.6732 ps=4.41 w=4.08 l=2.05
X13 VTAIL.t0 VP.t5 VDD1.t2 w_n3350_n1784# sky130_fd_pr__pfet_01v8 ad=1.5912 pd=8.94 as=0.6732 ps=4.41 w=4.08 l=2.05
X14 B.t5 B.t3 B.t4 w_n3350_n1784# sky130_fd_pr__pfet_01v8 ad=1.5912 pd=8.94 as=0 ps=0 w=4.08 l=2.05
X15 VTAIL.t6 VP.t6 VDD1.t1 w_n3350_n1784# sky130_fd_pr__pfet_01v8 ad=0.6732 pd=4.41 as=0.6732 ps=4.41 w=4.08 l=2.05
X16 VTAIL.t4 VP.t7 VDD1.t0 w_n3350_n1784# sky130_fd_pr__pfet_01v8 ad=1.5912 pd=8.94 as=0.6732 ps=4.41 w=4.08 l=2.05
X17 VDD2.t2 VN.t6 VTAIL.t8 w_n3350_n1784# sky130_fd_pr__pfet_01v8 ad=0.6732 pd=4.41 as=1.5912 ps=8.94 w=4.08 l=2.05
X18 VDD2.t7 VN.t7 VTAIL.t7 w_n3350_n1784# sky130_fd_pr__pfet_01v8 ad=0.6732 pd=4.41 as=0.6732 ps=4.41 w=4.08 l=2.05
X19 B.t2 B.t0 B.t1 w_n3350_n1784# sky130_fd_pr__pfet_01v8 ad=1.5912 pd=8.94 as=0 ps=0 w=4.08 l=2.05
R0 VN.n43 VN.n23 161.3
R1 VN.n42 VN.n41 161.3
R2 VN.n40 VN.n24 161.3
R3 VN.n39 VN.n38 161.3
R4 VN.n37 VN.n25 161.3
R5 VN.n35 VN.n34 161.3
R6 VN.n33 VN.n26 161.3
R7 VN.n32 VN.n31 161.3
R8 VN.n30 VN.n27 161.3
R9 VN.n20 VN.n0 161.3
R10 VN.n19 VN.n18 161.3
R11 VN.n17 VN.n1 161.3
R12 VN.n16 VN.n15 161.3
R13 VN.n14 VN.n2 161.3
R14 VN.n12 VN.n11 161.3
R15 VN.n10 VN.n3 161.3
R16 VN.n9 VN.n8 161.3
R17 VN.n7 VN.n4 161.3
R18 VN.n22 VN.n21 95.1695
R19 VN.n45 VN.n44 95.1695
R20 VN.n5 VN.t0 81.2878
R21 VN.n28 VN.t2 81.2878
R22 VN.n8 VN.n3 56.5617
R23 VN.n31 VN.n26 56.5617
R24 VN.n19 VN.n1 53.171
R25 VN.n42 VN.n24 53.171
R26 VN.n6 VN.n5 49.1088
R27 VN.n29 VN.n28 49.1088
R28 VN.n6 VN.t3 47.9654
R29 VN.n13 VN.t4 47.9654
R30 VN.n21 VN.t6 47.9654
R31 VN.n29 VN.t5 47.9654
R32 VN.n36 VN.t7 47.9654
R33 VN.n44 VN.t1 47.9654
R34 VN VN.n45 42.5739
R35 VN.n15 VN.n1 27.983
R36 VN.n38 VN.n24 27.983
R37 VN.n8 VN.n7 24.5923
R38 VN.n12 VN.n3 24.5923
R39 VN.n15 VN.n14 24.5923
R40 VN.n20 VN.n19 24.5923
R41 VN.n31 VN.n30 24.5923
R42 VN.n38 VN.n37 24.5923
R43 VN.n35 VN.n26 24.5923
R44 VN.n43 VN.n42 24.5923
R45 VN.n7 VN.n6 21.6413
R46 VN.n13 VN.n12 21.6413
R47 VN.n30 VN.n29 21.6413
R48 VN.n36 VN.n35 21.6413
R49 VN.n21 VN.n20 15.7393
R50 VN.n44 VN.n43 15.7393
R51 VN.n28 VN.n27 9.35282
R52 VN.n5 VN.n4 9.35282
R53 VN.n14 VN.n13 2.95152
R54 VN.n37 VN.n36 2.95152
R55 VN.n45 VN.n23 0.278335
R56 VN.n22 VN.n0 0.278335
R57 VN.n41 VN.n23 0.189894
R58 VN.n41 VN.n40 0.189894
R59 VN.n40 VN.n39 0.189894
R60 VN.n39 VN.n25 0.189894
R61 VN.n34 VN.n25 0.189894
R62 VN.n34 VN.n33 0.189894
R63 VN.n33 VN.n32 0.189894
R64 VN.n32 VN.n27 0.189894
R65 VN.n9 VN.n4 0.189894
R66 VN.n10 VN.n9 0.189894
R67 VN.n11 VN.n10 0.189894
R68 VN.n11 VN.n2 0.189894
R69 VN.n16 VN.n2 0.189894
R70 VN.n17 VN.n16 0.189894
R71 VN.n18 VN.n17 0.189894
R72 VN.n18 VN.n0 0.189894
R73 VN VN.n22 0.153485
R74 VDD2.n2 VDD2.n1 107.029
R75 VDD2.n2 VDD2.n0 107.029
R76 VDD2 VDD2.n5 107.026
R77 VDD2.n4 VDD2.n3 106.059
R78 VDD2.n4 VDD2.n2 36.4653
R79 VDD2.n5 VDD2.t3 7.96741
R80 VDD2.n5 VDD2.t5 7.96741
R81 VDD2.n3 VDD2.t0 7.96741
R82 VDD2.n3 VDD2.t7 7.96741
R83 VDD2.n1 VDD2.t4 7.96741
R84 VDD2.n1 VDD2.t2 7.96741
R85 VDD2.n0 VDD2.t1 7.96741
R86 VDD2.n0 VDD2.t6 7.96741
R87 VDD2 VDD2.n4 1.08455
R88 VTAIL.n11 VTAIL.t4 97.3475
R89 VTAIL.n10 VTAIL.t12 97.3475
R90 VTAIL.n7 VTAIL.t13 97.3475
R91 VTAIL.n15 VTAIL.t8 97.3472
R92 VTAIL.n2 VTAIL.t14 97.3472
R93 VTAIL.n3 VTAIL.t15 97.3472
R94 VTAIL.n6 VTAIL.t0 97.3472
R95 VTAIL.n14 VTAIL.t2 97.3472
R96 VTAIL.n13 VTAIL.n12 89.3806
R97 VTAIL.n9 VTAIL.n8 89.3806
R98 VTAIL.n1 VTAIL.n0 89.3803
R99 VTAIL.n5 VTAIL.n4 89.3803
R100 VTAIL.n15 VTAIL.n14 17.9358
R101 VTAIL.n7 VTAIL.n6 17.9358
R102 VTAIL.n0 VTAIL.t11 7.96741
R103 VTAIL.n0 VTAIL.t10 7.96741
R104 VTAIL.n4 VTAIL.t1 7.96741
R105 VTAIL.n4 VTAIL.t6 7.96741
R106 VTAIL.n12 VTAIL.t3 7.96741
R107 VTAIL.n12 VTAIL.t5 7.96741
R108 VTAIL.n8 VTAIL.t7 7.96741
R109 VTAIL.n8 VTAIL.t9 7.96741
R110 VTAIL.n9 VTAIL.n7 2.05222
R111 VTAIL.n10 VTAIL.n9 2.05222
R112 VTAIL.n13 VTAIL.n11 2.05222
R113 VTAIL.n14 VTAIL.n13 2.05222
R114 VTAIL.n6 VTAIL.n5 2.05222
R115 VTAIL.n5 VTAIL.n3 2.05222
R116 VTAIL.n2 VTAIL.n1 2.05222
R117 VTAIL VTAIL.n15 1.99403
R118 VTAIL.n11 VTAIL.n10 0.470328
R119 VTAIL.n3 VTAIL.n2 0.470328
R120 VTAIL VTAIL.n1 0.0586897
R121 B.n408 B.n51 585
R122 B.n410 B.n409 585
R123 B.n411 B.n50 585
R124 B.n413 B.n412 585
R125 B.n414 B.n49 585
R126 B.n416 B.n415 585
R127 B.n417 B.n48 585
R128 B.n419 B.n418 585
R129 B.n420 B.n47 585
R130 B.n422 B.n421 585
R131 B.n423 B.n46 585
R132 B.n425 B.n424 585
R133 B.n426 B.n45 585
R134 B.n428 B.n427 585
R135 B.n429 B.n44 585
R136 B.n431 B.n430 585
R137 B.n432 B.n43 585
R138 B.n434 B.n433 585
R139 B.n436 B.n40 585
R140 B.n438 B.n437 585
R141 B.n439 B.n39 585
R142 B.n441 B.n440 585
R143 B.n442 B.n38 585
R144 B.n444 B.n443 585
R145 B.n445 B.n37 585
R146 B.n447 B.n446 585
R147 B.n448 B.n33 585
R148 B.n450 B.n449 585
R149 B.n451 B.n32 585
R150 B.n453 B.n452 585
R151 B.n454 B.n31 585
R152 B.n456 B.n455 585
R153 B.n457 B.n30 585
R154 B.n459 B.n458 585
R155 B.n460 B.n29 585
R156 B.n462 B.n461 585
R157 B.n463 B.n28 585
R158 B.n465 B.n464 585
R159 B.n466 B.n27 585
R160 B.n468 B.n467 585
R161 B.n469 B.n26 585
R162 B.n471 B.n470 585
R163 B.n472 B.n25 585
R164 B.n474 B.n473 585
R165 B.n475 B.n24 585
R166 B.n477 B.n476 585
R167 B.n407 B.n406 585
R168 B.n405 B.n52 585
R169 B.n404 B.n403 585
R170 B.n402 B.n53 585
R171 B.n401 B.n400 585
R172 B.n399 B.n54 585
R173 B.n398 B.n397 585
R174 B.n396 B.n55 585
R175 B.n395 B.n394 585
R176 B.n393 B.n56 585
R177 B.n392 B.n391 585
R178 B.n390 B.n57 585
R179 B.n389 B.n388 585
R180 B.n387 B.n58 585
R181 B.n386 B.n385 585
R182 B.n384 B.n59 585
R183 B.n383 B.n382 585
R184 B.n381 B.n60 585
R185 B.n380 B.n379 585
R186 B.n378 B.n61 585
R187 B.n377 B.n376 585
R188 B.n375 B.n62 585
R189 B.n374 B.n373 585
R190 B.n372 B.n63 585
R191 B.n371 B.n370 585
R192 B.n369 B.n64 585
R193 B.n368 B.n367 585
R194 B.n366 B.n65 585
R195 B.n365 B.n364 585
R196 B.n363 B.n66 585
R197 B.n362 B.n361 585
R198 B.n360 B.n67 585
R199 B.n359 B.n358 585
R200 B.n357 B.n68 585
R201 B.n356 B.n355 585
R202 B.n354 B.n69 585
R203 B.n353 B.n352 585
R204 B.n351 B.n70 585
R205 B.n350 B.n349 585
R206 B.n348 B.n71 585
R207 B.n347 B.n346 585
R208 B.n345 B.n72 585
R209 B.n344 B.n343 585
R210 B.n342 B.n73 585
R211 B.n341 B.n340 585
R212 B.n339 B.n74 585
R213 B.n338 B.n337 585
R214 B.n336 B.n75 585
R215 B.n335 B.n334 585
R216 B.n333 B.n76 585
R217 B.n332 B.n331 585
R218 B.n330 B.n77 585
R219 B.n329 B.n328 585
R220 B.n327 B.n78 585
R221 B.n326 B.n325 585
R222 B.n324 B.n79 585
R223 B.n323 B.n322 585
R224 B.n321 B.n80 585
R225 B.n320 B.n319 585
R226 B.n318 B.n81 585
R227 B.n317 B.n316 585
R228 B.n315 B.n82 585
R229 B.n314 B.n313 585
R230 B.n312 B.n83 585
R231 B.n311 B.n310 585
R232 B.n309 B.n84 585
R233 B.n308 B.n307 585
R234 B.n306 B.n85 585
R235 B.n305 B.n304 585
R236 B.n303 B.n86 585
R237 B.n302 B.n301 585
R238 B.n300 B.n87 585
R239 B.n299 B.n298 585
R240 B.n297 B.n88 585
R241 B.n296 B.n295 585
R242 B.n294 B.n89 585
R243 B.n293 B.n292 585
R244 B.n291 B.n90 585
R245 B.n290 B.n289 585
R246 B.n288 B.n91 585
R247 B.n287 B.n286 585
R248 B.n285 B.n92 585
R249 B.n284 B.n283 585
R250 B.n282 B.n93 585
R251 B.n281 B.n280 585
R252 B.n279 B.n94 585
R253 B.n278 B.n277 585
R254 B.n207 B.n122 585
R255 B.n209 B.n208 585
R256 B.n210 B.n121 585
R257 B.n212 B.n211 585
R258 B.n213 B.n120 585
R259 B.n215 B.n214 585
R260 B.n216 B.n119 585
R261 B.n218 B.n217 585
R262 B.n219 B.n118 585
R263 B.n221 B.n220 585
R264 B.n222 B.n117 585
R265 B.n224 B.n223 585
R266 B.n225 B.n116 585
R267 B.n227 B.n226 585
R268 B.n228 B.n115 585
R269 B.n230 B.n229 585
R270 B.n231 B.n114 585
R271 B.n233 B.n232 585
R272 B.n235 B.n234 585
R273 B.n236 B.n110 585
R274 B.n238 B.n237 585
R275 B.n239 B.n109 585
R276 B.n241 B.n240 585
R277 B.n242 B.n108 585
R278 B.n244 B.n243 585
R279 B.n245 B.n107 585
R280 B.n247 B.n246 585
R281 B.n248 B.n104 585
R282 B.n251 B.n250 585
R283 B.n252 B.n103 585
R284 B.n254 B.n253 585
R285 B.n255 B.n102 585
R286 B.n257 B.n256 585
R287 B.n258 B.n101 585
R288 B.n260 B.n259 585
R289 B.n261 B.n100 585
R290 B.n263 B.n262 585
R291 B.n264 B.n99 585
R292 B.n266 B.n265 585
R293 B.n267 B.n98 585
R294 B.n269 B.n268 585
R295 B.n270 B.n97 585
R296 B.n272 B.n271 585
R297 B.n273 B.n96 585
R298 B.n275 B.n274 585
R299 B.n276 B.n95 585
R300 B.n206 B.n205 585
R301 B.n204 B.n123 585
R302 B.n203 B.n202 585
R303 B.n201 B.n124 585
R304 B.n200 B.n199 585
R305 B.n198 B.n125 585
R306 B.n197 B.n196 585
R307 B.n195 B.n126 585
R308 B.n194 B.n193 585
R309 B.n192 B.n127 585
R310 B.n191 B.n190 585
R311 B.n189 B.n128 585
R312 B.n188 B.n187 585
R313 B.n186 B.n129 585
R314 B.n185 B.n184 585
R315 B.n183 B.n130 585
R316 B.n182 B.n181 585
R317 B.n180 B.n131 585
R318 B.n179 B.n178 585
R319 B.n177 B.n132 585
R320 B.n176 B.n175 585
R321 B.n174 B.n133 585
R322 B.n173 B.n172 585
R323 B.n171 B.n134 585
R324 B.n170 B.n169 585
R325 B.n168 B.n135 585
R326 B.n167 B.n166 585
R327 B.n165 B.n136 585
R328 B.n164 B.n163 585
R329 B.n162 B.n137 585
R330 B.n161 B.n160 585
R331 B.n159 B.n138 585
R332 B.n158 B.n157 585
R333 B.n156 B.n139 585
R334 B.n155 B.n154 585
R335 B.n153 B.n140 585
R336 B.n152 B.n151 585
R337 B.n150 B.n141 585
R338 B.n149 B.n148 585
R339 B.n147 B.n142 585
R340 B.n146 B.n145 585
R341 B.n144 B.n143 585
R342 B.n2 B.n0 585
R343 B.n541 B.n1 585
R344 B.n540 B.n539 585
R345 B.n538 B.n3 585
R346 B.n537 B.n536 585
R347 B.n535 B.n4 585
R348 B.n534 B.n533 585
R349 B.n532 B.n5 585
R350 B.n531 B.n530 585
R351 B.n529 B.n6 585
R352 B.n528 B.n527 585
R353 B.n526 B.n7 585
R354 B.n525 B.n524 585
R355 B.n523 B.n8 585
R356 B.n522 B.n521 585
R357 B.n520 B.n9 585
R358 B.n519 B.n518 585
R359 B.n517 B.n10 585
R360 B.n516 B.n515 585
R361 B.n514 B.n11 585
R362 B.n513 B.n512 585
R363 B.n511 B.n12 585
R364 B.n510 B.n509 585
R365 B.n508 B.n13 585
R366 B.n507 B.n506 585
R367 B.n505 B.n14 585
R368 B.n504 B.n503 585
R369 B.n502 B.n15 585
R370 B.n501 B.n500 585
R371 B.n499 B.n16 585
R372 B.n498 B.n497 585
R373 B.n496 B.n17 585
R374 B.n495 B.n494 585
R375 B.n493 B.n18 585
R376 B.n492 B.n491 585
R377 B.n490 B.n19 585
R378 B.n489 B.n488 585
R379 B.n487 B.n20 585
R380 B.n486 B.n485 585
R381 B.n484 B.n21 585
R382 B.n483 B.n482 585
R383 B.n481 B.n22 585
R384 B.n480 B.n479 585
R385 B.n478 B.n23 585
R386 B.n543 B.n542 585
R387 B.n205 B.n122 535.745
R388 B.n476 B.n23 535.745
R389 B.n277 B.n276 535.745
R390 B.n408 B.n407 535.745
R391 B.n105 B.t9 254.998
R392 B.n111 B.t3 254.998
R393 B.n34 B.t6 254.998
R394 B.n41 B.t0 254.998
R395 B.n105 B.t11 165.249
R396 B.n41 B.t1 165.249
R397 B.n111 B.t5 165.244
R398 B.n34 B.t7 165.244
R399 B.n205 B.n204 163.367
R400 B.n204 B.n203 163.367
R401 B.n203 B.n124 163.367
R402 B.n199 B.n124 163.367
R403 B.n199 B.n198 163.367
R404 B.n198 B.n197 163.367
R405 B.n197 B.n126 163.367
R406 B.n193 B.n126 163.367
R407 B.n193 B.n192 163.367
R408 B.n192 B.n191 163.367
R409 B.n191 B.n128 163.367
R410 B.n187 B.n128 163.367
R411 B.n187 B.n186 163.367
R412 B.n186 B.n185 163.367
R413 B.n185 B.n130 163.367
R414 B.n181 B.n130 163.367
R415 B.n181 B.n180 163.367
R416 B.n180 B.n179 163.367
R417 B.n179 B.n132 163.367
R418 B.n175 B.n132 163.367
R419 B.n175 B.n174 163.367
R420 B.n174 B.n173 163.367
R421 B.n173 B.n134 163.367
R422 B.n169 B.n134 163.367
R423 B.n169 B.n168 163.367
R424 B.n168 B.n167 163.367
R425 B.n167 B.n136 163.367
R426 B.n163 B.n136 163.367
R427 B.n163 B.n162 163.367
R428 B.n162 B.n161 163.367
R429 B.n161 B.n138 163.367
R430 B.n157 B.n138 163.367
R431 B.n157 B.n156 163.367
R432 B.n156 B.n155 163.367
R433 B.n155 B.n140 163.367
R434 B.n151 B.n140 163.367
R435 B.n151 B.n150 163.367
R436 B.n150 B.n149 163.367
R437 B.n149 B.n142 163.367
R438 B.n145 B.n142 163.367
R439 B.n145 B.n144 163.367
R440 B.n144 B.n2 163.367
R441 B.n542 B.n2 163.367
R442 B.n542 B.n541 163.367
R443 B.n541 B.n540 163.367
R444 B.n540 B.n3 163.367
R445 B.n536 B.n3 163.367
R446 B.n536 B.n535 163.367
R447 B.n535 B.n534 163.367
R448 B.n534 B.n5 163.367
R449 B.n530 B.n5 163.367
R450 B.n530 B.n529 163.367
R451 B.n529 B.n528 163.367
R452 B.n528 B.n7 163.367
R453 B.n524 B.n7 163.367
R454 B.n524 B.n523 163.367
R455 B.n523 B.n522 163.367
R456 B.n522 B.n9 163.367
R457 B.n518 B.n9 163.367
R458 B.n518 B.n517 163.367
R459 B.n517 B.n516 163.367
R460 B.n516 B.n11 163.367
R461 B.n512 B.n11 163.367
R462 B.n512 B.n511 163.367
R463 B.n511 B.n510 163.367
R464 B.n510 B.n13 163.367
R465 B.n506 B.n13 163.367
R466 B.n506 B.n505 163.367
R467 B.n505 B.n504 163.367
R468 B.n504 B.n15 163.367
R469 B.n500 B.n15 163.367
R470 B.n500 B.n499 163.367
R471 B.n499 B.n498 163.367
R472 B.n498 B.n17 163.367
R473 B.n494 B.n17 163.367
R474 B.n494 B.n493 163.367
R475 B.n493 B.n492 163.367
R476 B.n492 B.n19 163.367
R477 B.n488 B.n19 163.367
R478 B.n488 B.n487 163.367
R479 B.n487 B.n486 163.367
R480 B.n486 B.n21 163.367
R481 B.n482 B.n21 163.367
R482 B.n482 B.n481 163.367
R483 B.n481 B.n480 163.367
R484 B.n480 B.n23 163.367
R485 B.n209 B.n122 163.367
R486 B.n210 B.n209 163.367
R487 B.n211 B.n210 163.367
R488 B.n211 B.n120 163.367
R489 B.n215 B.n120 163.367
R490 B.n216 B.n215 163.367
R491 B.n217 B.n216 163.367
R492 B.n217 B.n118 163.367
R493 B.n221 B.n118 163.367
R494 B.n222 B.n221 163.367
R495 B.n223 B.n222 163.367
R496 B.n223 B.n116 163.367
R497 B.n227 B.n116 163.367
R498 B.n228 B.n227 163.367
R499 B.n229 B.n228 163.367
R500 B.n229 B.n114 163.367
R501 B.n233 B.n114 163.367
R502 B.n234 B.n233 163.367
R503 B.n234 B.n110 163.367
R504 B.n238 B.n110 163.367
R505 B.n239 B.n238 163.367
R506 B.n240 B.n239 163.367
R507 B.n240 B.n108 163.367
R508 B.n244 B.n108 163.367
R509 B.n245 B.n244 163.367
R510 B.n246 B.n245 163.367
R511 B.n246 B.n104 163.367
R512 B.n251 B.n104 163.367
R513 B.n252 B.n251 163.367
R514 B.n253 B.n252 163.367
R515 B.n253 B.n102 163.367
R516 B.n257 B.n102 163.367
R517 B.n258 B.n257 163.367
R518 B.n259 B.n258 163.367
R519 B.n259 B.n100 163.367
R520 B.n263 B.n100 163.367
R521 B.n264 B.n263 163.367
R522 B.n265 B.n264 163.367
R523 B.n265 B.n98 163.367
R524 B.n269 B.n98 163.367
R525 B.n270 B.n269 163.367
R526 B.n271 B.n270 163.367
R527 B.n271 B.n96 163.367
R528 B.n275 B.n96 163.367
R529 B.n276 B.n275 163.367
R530 B.n277 B.n94 163.367
R531 B.n281 B.n94 163.367
R532 B.n282 B.n281 163.367
R533 B.n283 B.n282 163.367
R534 B.n283 B.n92 163.367
R535 B.n287 B.n92 163.367
R536 B.n288 B.n287 163.367
R537 B.n289 B.n288 163.367
R538 B.n289 B.n90 163.367
R539 B.n293 B.n90 163.367
R540 B.n294 B.n293 163.367
R541 B.n295 B.n294 163.367
R542 B.n295 B.n88 163.367
R543 B.n299 B.n88 163.367
R544 B.n300 B.n299 163.367
R545 B.n301 B.n300 163.367
R546 B.n301 B.n86 163.367
R547 B.n305 B.n86 163.367
R548 B.n306 B.n305 163.367
R549 B.n307 B.n306 163.367
R550 B.n307 B.n84 163.367
R551 B.n311 B.n84 163.367
R552 B.n312 B.n311 163.367
R553 B.n313 B.n312 163.367
R554 B.n313 B.n82 163.367
R555 B.n317 B.n82 163.367
R556 B.n318 B.n317 163.367
R557 B.n319 B.n318 163.367
R558 B.n319 B.n80 163.367
R559 B.n323 B.n80 163.367
R560 B.n324 B.n323 163.367
R561 B.n325 B.n324 163.367
R562 B.n325 B.n78 163.367
R563 B.n329 B.n78 163.367
R564 B.n330 B.n329 163.367
R565 B.n331 B.n330 163.367
R566 B.n331 B.n76 163.367
R567 B.n335 B.n76 163.367
R568 B.n336 B.n335 163.367
R569 B.n337 B.n336 163.367
R570 B.n337 B.n74 163.367
R571 B.n341 B.n74 163.367
R572 B.n342 B.n341 163.367
R573 B.n343 B.n342 163.367
R574 B.n343 B.n72 163.367
R575 B.n347 B.n72 163.367
R576 B.n348 B.n347 163.367
R577 B.n349 B.n348 163.367
R578 B.n349 B.n70 163.367
R579 B.n353 B.n70 163.367
R580 B.n354 B.n353 163.367
R581 B.n355 B.n354 163.367
R582 B.n355 B.n68 163.367
R583 B.n359 B.n68 163.367
R584 B.n360 B.n359 163.367
R585 B.n361 B.n360 163.367
R586 B.n361 B.n66 163.367
R587 B.n365 B.n66 163.367
R588 B.n366 B.n365 163.367
R589 B.n367 B.n366 163.367
R590 B.n367 B.n64 163.367
R591 B.n371 B.n64 163.367
R592 B.n372 B.n371 163.367
R593 B.n373 B.n372 163.367
R594 B.n373 B.n62 163.367
R595 B.n377 B.n62 163.367
R596 B.n378 B.n377 163.367
R597 B.n379 B.n378 163.367
R598 B.n379 B.n60 163.367
R599 B.n383 B.n60 163.367
R600 B.n384 B.n383 163.367
R601 B.n385 B.n384 163.367
R602 B.n385 B.n58 163.367
R603 B.n389 B.n58 163.367
R604 B.n390 B.n389 163.367
R605 B.n391 B.n390 163.367
R606 B.n391 B.n56 163.367
R607 B.n395 B.n56 163.367
R608 B.n396 B.n395 163.367
R609 B.n397 B.n396 163.367
R610 B.n397 B.n54 163.367
R611 B.n401 B.n54 163.367
R612 B.n402 B.n401 163.367
R613 B.n403 B.n402 163.367
R614 B.n403 B.n52 163.367
R615 B.n407 B.n52 163.367
R616 B.n476 B.n475 163.367
R617 B.n475 B.n474 163.367
R618 B.n474 B.n25 163.367
R619 B.n470 B.n25 163.367
R620 B.n470 B.n469 163.367
R621 B.n469 B.n468 163.367
R622 B.n468 B.n27 163.367
R623 B.n464 B.n27 163.367
R624 B.n464 B.n463 163.367
R625 B.n463 B.n462 163.367
R626 B.n462 B.n29 163.367
R627 B.n458 B.n29 163.367
R628 B.n458 B.n457 163.367
R629 B.n457 B.n456 163.367
R630 B.n456 B.n31 163.367
R631 B.n452 B.n31 163.367
R632 B.n452 B.n451 163.367
R633 B.n451 B.n450 163.367
R634 B.n450 B.n33 163.367
R635 B.n446 B.n33 163.367
R636 B.n446 B.n445 163.367
R637 B.n445 B.n444 163.367
R638 B.n444 B.n38 163.367
R639 B.n440 B.n38 163.367
R640 B.n440 B.n439 163.367
R641 B.n439 B.n438 163.367
R642 B.n438 B.n40 163.367
R643 B.n433 B.n40 163.367
R644 B.n433 B.n432 163.367
R645 B.n432 B.n431 163.367
R646 B.n431 B.n44 163.367
R647 B.n427 B.n44 163.367
R648 B.n427 B.n426 163.367
R649 B.n426 B.n425 163.367
R650 B.n425 B.n46 163.367
R651 B.n421 B.n46 163.367
R652 B.n421 B.n420 163.367
R653 B.n420 B.n419 163.367
R654 B.n419 B.n48 163.367
R655 B.n415 B.n48 163.367
R656 B.n415 B.n414 163.367
R657 B.n414 B.n413 163.367
R658 B.n413 B.n50 163.367
R659 B.n409 B.n50 163.367
R660 B.n409 B.n408 163.367
R661 B.n106 B.t10 119.091
R662 B.n42 B.t2 119.091
R663 B.n112 B.t4 119.088
R664 B.n35 B.t8 119.088
R665 B.n249 B.n106 59.5399
R666 B.n113 B.n112 59.5399
R667 B.n36 B.n35 59.5399
R668 B.n435 B.n42 59.5399
R669 B.n106 B.n105 46.1581
R670 B.n112 B.n111 46.1581
R671 B.n35 B.n34 46.1581
R672 B.n42 B.n41 46.1581
R673 B.n478 B.n477 34.8103
R674 B.n406 B.n51 34.8103
R675 B.n278 B.n95 34.8103
R676 B.n207 B.n206 34.8103
R677 B B.n543 18.0485
R678 B.n477 B.n24 10.6151
R679 B.n473 B.n24 10.6151
R680 B.n473 B.n472 10.6151
R681 B.n472 B.n471 10.6151
R682 B.n471 B.n26 10.6151
R683 B.n467 B.n26 10.6151
R684 B.n467 B.n466 10.6151
R685 B.n466 B.n465 10.6151
R686 B.n465 B.n28 10.6151
R687 B.n461 B.n28 10.6151
R688 B.n461 B.n460 10.6151
R689 B.n460 B.n459 10.6151
R690 B.n459 B.n30 10.6151
R691 B.n455 B.n30 10.6151
R692 B.n455 B.n454 10.6151
R693 B.n454 B.n453 10.6151
R694 B.n453 B.n32 10.6151
R695 B.n449 B.n448 10.6151
R696 B.n448 B.n447 10.6151
R697 B.n447 B.n37 10.6151
R698 B.n443 B.n37 10.6151
R699 B.n443 B.n442 10.6151
R700 B.n442 B.n441 10.6151
R701 B.n441 B.n39 10.6151
R702 B.n437 B.n39 10.6151
R703 B.n437 B.n436 10.6151
R704 B.n434 B.n43 10.6151
R705 B.n430 B.n43 10.6151
R706 B.n430 B.n429 10.6151
R707 B.n429 B.n428 10.6151
R708 B.n428 B.n45 10.6151
R709 B.n424 B.n45 10.6151
R710 B.n424 B.n423 10.6151
R711 B.n423 B.n422 10.6151
R712 B.n422 B.n47 10.6151
R713 B.n418 B.n47 10.6151
R714 B.n418 B.n417 10.6151
R715 B.n417 B.n416 10.6151
R716 B.n416 B.n49 10.6151
R717 B.n412 B.n49 10.6151
R718 B.n412 B.n411 10.6151
R719 B.n411 B.n410 10.6151
R720 B.n410 B.n51 10.6151
R721 B.n279 B.n278 10.6151
R722 B.n280 B.n279 10.6151
R723 B.n280 B.n93 10.6151
R724 B.n284 B.n93 10.6151
R725 B.n285 B.n284 10.6151
R726 B.n286 B.n285 10.6151
R727 B.n286 B.n91 10.6151
R728 B.n290 B.n91 10.6151
R729 B.n291 B.n290 10.6151
R730 B.n292 B.n291 10.6151
R731 B.n292 B.n89 10.6151
R732 B.n296 B.n89 10.6151
R733 B.n297 B.n296 10.6151
R734 B.n298 B.n297 10.6151
R735 B.n298 B.n87 10.6151
R736 B.n302 B.n87 10.6151
R737 B.n303 B.n302 10.6151
R738 B.n304 B.n303 10.6151
R739 B.n304 B.n85 10.6151
R740 B.n308 B.n85 10.6151
R741 B.n309 B.n308 10.6151
R742 B.n310 B.n309 10.6151
R743 B.n310 B.n83 10.6151
R744 B.n314 B.n83 10.6151
R745 B.n315 B.n314 10.6151
R746 B.n316 B.n315 10.6151
R747 B.n316 B.n81 10.6151
R748 B.n320 B.n81 10.6151
R749 B.n321 B.n320 10.6151
R750 B.n322 B.n321 10.6151
R751 B.n322 B.n79 10.6151
R752 B.n326 B.n79 10.6151
R753 B.n327 B.n326 10.6151
R754 B.n328 B.n327 10.6151
R755 B.n328 B.n77 10.6151
R756 B.n332 B.n77 10.6151
R757 B.n333 B.n332 10.6151
R758 B.n334 B.n333 10.6151
R759 B.n334 B.n75 10.6151
R760 B.n338 B.n75 10.6151
R761 B.n339 B.n338 10.6151
R762 B.n340 B.n339 10.6151
R763 B.n340 B.n73 10.6151
R764 B.n344 B.n73 10.6151
R765 B.n345 B.n344 10.6151
R766 B.n346 B.n345 10.6151
R767 B.n346 B.n71 10.6151
R768 B.n350 B.n71 10.6151
R769 B.n351 B.n350 10.6151
R770 B.n352 B.n351 10.6151
R771 B.n352 B.n69 10.6151
R772 B.n356 B.n69 10.6151
R773 B.n357 B.n356 10.6151
R774 B.n358 B.n357 10.6151
R775 B.n358 B.n67 10.6151
R776 B.n362 B.n67 10.6151
R777 B.n363 B.n362 10.6151
R778 B.n364 B.n363 10.6151
R779 B.n364 B.n65 10.6151
R780 B.n368 B.n65 10.6151
R781 B.n369 B.n368 10.6151
R782 B.n370 B.n369 10.6151
R783 B.n370 B.n63 10.6151
R784 B.n374 B.n63 10.6151
R785 B.n375 B.n374 10.6151
R786 B.n376 B.n375 10.6151
R787 B.n376 B.n61 10.6151
R788 B.n380 B.n61 10.6151
R789 B.n381 B.n380 10.6151
R790 B.n382 B.n381 10.6151
R791 B.n382 B.n59 10.6151
R792 B.n386 B.n59 10.6151
R793 B.n387 B.n386 10.6151
R794 B.n388 B.n387 10.6151
R795 B.n388 B.n57 10.6151
R796 B.n392 B.n57 10.6151
R797 B.n393 B.n392 10.6151
R798 B.n394 B.n393 10.6151
R799 B.n394 B.n55 10.6151
R800 B.n398 B.n55 10.6151
R801 B.n399 B.n398 10.6151
R802 B.n400 B.n399 10.6151
R803 B.n400 B.n53 10.6151
R804 B.n404 B.n53 10.6151
R805 B.n405 B.n404 10.6151
R806 B.n406 B.n405 10.6151
R807 B.n208 B.n207 10.6151
R808 B.n208 B.n121 10.6151
R809 B.n212 B.n121 10.6151
R810 B.n213 B.n212 10.6151
R811 B.n214 B.n213 10.6151
R812 B.n214 B.n119 10.6151
R813 B.n218 B.n119 10.6151
R814 B.n219 B.n218 10.6151
R815 B.n220 B.n219 10.6151
R816 B.n220 B.n117 10.6151
R817 B.n224 B.n117 10.6151
R818 B.n225 B.n224 10.6151
R819 B.n226 B.n225 10.6151
R820 B.n226 B.n115 10.6151
R821 B.n230 B.n115 10.6151
R822 B.n231 B.n230 10.6151
R823 B.n232 B.n231 10.6151
R824 B.n236 B.n235 10.6151
R825 B.n237 B.n236 10.6151
R826 B.n237 B.n109 10.6151
R827 B.n241 B.n109 10.6151
R828 B.n242 B.n241 10.6151
R829 B.n243 B.n242 10.6151
R830 B.n243 B.n107 10.6151
R831 B.n247 B.n107 10.6151
R832 B.n248 B.n247 10.6151
R833 B.n250 B.n103 10.6151
R834 B.n254 B.n103 10.6151
R835 B.n255 B.n254 10.6151
R836 B.n256 B.n255 10.6151
R837 B.n256 B.n101 10.6151
R838 B.n260 B.n101 10.6151
R839 B.n261 B.n260 10.6151
R840 B.n262 B.n261 10.6151
R841 B.n262 B.n99 10.6151
R842 B.n266 B.n99 10.6151
R843 B.n267 B.n266 10.6151
R844 B.n268 B.n267 10.6151
R845 B.n268 B.n97 10.6151
R846 B.n272 B.n97 10.6151
R847 B.n273 B.n272 10.6151
R848 B.n274 B.n273 10.6151
R849 B.n274 B.n95 10.6151
R850 B.n206 B.n123 10.6151
R851 B.n202 B.n123 10.6151
R852 B.n202 B.n201 10.6151
R853 B.n201 B.n200 10.6151
R854 B.n200 B.n125 10.6151
R855 B.n196 B.n125 10.6151
R856 B.n196 B.n195 10.6151
R857 B.n195 B.n194 10.6151
R858 B.n194 B.n127 10.6151
R859 B.n190 B.n127 10.6151
R860 B.n190 B.n189 10.6151
R861 B.n189 B.n188 10.6151
R862 B.n188 B.n129 10.6151
R863 B.n184 B.n129 10.6151
R864 B.n184 B.n183 10.6151
R865 B.n183 B.n182 10.6151
R866 B.n182 B.n131 10.6151
R867 B.n178 B.n131 10.6151
R868 B.n178 B.n177 10.6151
R869 B.n177 B.n176 10.6151
R870 B.n176 B.n133 10.6151
R871 B.n172 B.n133 10.6151
R872 B.n172 B.n171 10.6151
R873 B.n171 B.n170 10.6151
R874 B.n170 B.n135 10.6151
R875 B.n166 B.n135 10.6151
R876 B.n166 B.n165 10.6151
R877 B.n165 B.n164 10.6151
R878 B.n164 B.n137 10.6151
R879 B.n160 B.n137 10.6151
R880 B.n160 B.n159 10.6151
R881 B.n159 B.n158 10.6151
R882 B.n158 B.n139 10.6151
R883 B.n154 B.n139 10.6151
R884 B.n154 B.n153 10.6151
R885 B.n153 B.n152 10.6151
R886 B.n152 B.n141 10.6151
R887 B.n148 B.n141 10.6151
R888 B.n148 B.n147 10.6151
R889 B.n147 B.n146 10.6151
R890 B.n146 B.n143 10.6151
R891 B.n143 B.n0 10.6151
R892 B.n539 B.n1 10.6151
R893 B.n539 B.n538 10.6151
R894 B.n538 B.n537 10.6151
R895 B.n537 B.n4 10.6151
R896 B.n533 B.n4 10.6151
R897 B.n533 B.n532 10.6151
R898 B.n532 B.n531 10.6151
R899 B.n531 B.n6 10.6151
R900 B.n527 B.n6 10.6151
R901 B.n527 B.n526 10.6151
R902 B.n526 B.n525 10.6151
R903 B.n525 B.n8 10.6151
R904 B.n521 B.n8 10.6151
R905 B.n521 B.n520 10.6151
R906 B.n520 B.n519 10.6151
R907 B.n519 B.n10 10.6151
R908 B.n515 B.n10 10.6151
R909 B.n515 B.n514 10.6151
R910 B.n514 B.n513 10.6151
R911 B.n513 B.n12 10.6151
R912 B.n509 B.n12 10.6151
R913 B.n509 B.n508 10.6151
R914 B.n508 B.n507 10.6151
R915 B.n507 B.n14 10.6151
R916 B.n503 B.n14 10.6151
R917 B.n503 B.n502 10.6151
R918 B.n502 B.n501 10.6151
R919 B.n501 B.n16 10.6151
R920 B.n497 B.n16 10.6151
R921 B.n497 B.n496 10.6151
R922 B.n496 B.n495 10.6151
R923 B.n495 B.n18 10.6151
R924 B.n491 B.n18 10.6151
R925 B.n491 B.n490 10.6151
R926 B.n490 B.n489 10.6151
R927 B.n489 B.n20 10.6151
R928 B.n485 B.n20 10.6151
R929 B.n485 B.n484 10.6151
R930 B.n484 B.n483 10.6151
R931 B.n483 B.n22 10.6151
R932 B.n479 B.n22 10.6151
R933 B.n479 B.n478 10.6151
R934 B.n36 B.n32 9.36635
R935 B.n435 B.n434 9.36635
R936 B.n232 B.n113 9.36635
R937 B.n250 B.n249 9.36635
R938 B.n543 B.n0 2.81026
R939 B.n543 B.n1 2.81026
R940 B.n449 B.n36 1.24928
R941 B.n436 B.n435 1.24928
R942 B.n235 B.n113 1.24928
R943 B.n249 B.n248 1.24928
R944 VP.n15 VP.n12 161.3
R945 VP.n17 VP.n16 161.3
R946 VP.n18 VP.n11 161.3
R947 VP.n20 VP.n19 161.3
R948 VP.n22 VP.n10 161.3
R949 VP.n24 VP.n23 161.3
R950 VP.n25 VP.n9 161.3
R951 VP.n27 VP.n26 161.3
R952 VP.n28 VP.n8 161.3
R953 VP.n54 VP.n0 161.3
R954 VP.n53 VP.n52 161.3
R955 VP.n51 VP.n1 161.3
R956 VP.n50 VP.n49 161.3
R957 VP.n48 VP.n2 161.3
R958 VP.n46 VP.n45 161.3
R959 VP.n44 VP.n3 161.3
R960 VP.n43 VP.n42 161.3
R961 VP.n41 VP.n4 161.3
R962 VP.n39 VP.n38 161.3
R963 VP.n37 VP.n5 161.3
R964 VP.n36 VP.n35 161.3
R965 VP.n34 VP.n6 161.3
R966 VP.n33 VP.n32 161.3
R967 VP.n31 VP.n7 95.1695
R968 VP.n56 VP.n55 95.1695
R969 VP.n30 VP.n29 95.1695
R970 VP.n13 VP.t7 81.2878
R971 VP.n42 VP.n3 56.5617
R972 VP.n16 VP.n11 56.5617
R973 VP.n35 VP.n34 53.171
R974 VP.n53 VP.n1 53.171
R975 VP.n27 VP.n9 53.171
R976 VP.n14 VP.n13 49.1088
R977 VP.n7 VP.t5 47.9654
R978 VP.n40 VP.t4 47.9654
R979 VP.n47 VP.t6 47.9654
R980 VP.n55 VP.t1 47.9654
R981 VP.n29 VP.t3 47.9654
R982 VP.n21 VP.t2 47.9654
R983 VP.n14 VP.t0 47.9654
R984 VP.n31 VP.n30 42.2951
R985 VP.n35 VP.n5 27.983
R986 VP.n49 VP.n1 27.983
R987 VP.n23 VP.n9 27.983
R988 VP.n34 VP.n33 24.5923
R989 VP.n39 VP.n5 24.5923
R990 VP.n42 VP.n41 24.5923
R991 VP.n46 VP.n3 24.5923
R992 VP.n49 VP.n48 24.5923
R993 VP.n54 VP.n53 24.5923
R994 VP.n28 VP.n27 24.5923
R995 VP.n20 VP.n11 24.5923
R996 VP.n23 VP.n22 24.5923
R997 VP.n16 VP.n15 24.5923
R998 VP.n41 VP.n40 21.6413
R999 VP.n47 VP.n46 21.6413
R1000 VP.n21 VP.n20 21.6413
R1001 VP.n15 VP.n14 21.6413
R1002 VP.n33 VP.n7 15.7393
R1003 VP.n55 VP.n54 15.7393
R1004 VP.n29 VP.n28 15.7393
R1005 VP.n13 VP.n12 9.35282
R1006 VP.n40 VP.n39 2.95152
R1007 VP.n48 VP.n47 2.95152
R1008 VP.n22 VP.n21 2.95152
R1009 VP.n30 VP.n8 0.278335
R1010 VP.n32 VP.n31 0.278335
R1011 VP.n56 VP.n0 0.278335
R1012 VP.n17 VP.n12 0.189894
R1013 VP.n18 VP.n17 0.189894
R1014 VP.n19 VP.n18 0.189894
R1015 VP.n19 VP.n10 0.189894
R1016 VP.n24 VP.n10 0.189894
R1017 VP.n25 VP.n24 0.189894
R1018 VP.n26 VP.n25 0.189894
R1019 VP.n26 VP.n8 0.189894
R1020 VP.n32 VP.n6 0.189894
R1021 VP.n36 VP.n6 0.189894
R1022 VP.n37 VP.n36 0.189894
R1023 VP.n38 VP.n37 0.189894
R1024 VP.n38 VP.n4 0.189894
R1025 VP.n43 VP.n4 0.189894
R1026 VP.n44 VP.n43 0.189894
R1027 VP.n45 VP.n44 0.189894
R1028 VP.n45 VP.n2 0.189894
R1029 VP.n50 VP.n2 0.189894
R1030 VP.n51 VP.n50 0.189894
R1031 VP.n52 VP.n51 0.189894
R1032 VP.n52 VP.n0 0.189894
R1033 VP VP.n56 0.153485
R1034 VDD1 VDD1.n0 107.144
R1035 VDD1.n3 VDD1.n2 107.029
R1036 VDD1.n3 VDD1.n1 107.029
R1037 VDD1.n5 VDD1.n4 106.059
R1038 VDD1.n5 VDD1.n3 37.0483
R1039 VDD1.n4 VDD1.t5 7.96741
R1040 VDD1.n4 VDD1.t4 7.96741
R1041 VDD1.n0 VDD1.t0 7.96741
R1042 VDD1.n0 VDD1.t7 7.96741
R1043 VDD1.n2 VDD1.t1 7.96741
R1044 VDD1.n2 VDD1.t6 7.96741
R1045 VDD1.n1 VDD1.t2 7.96741
R1046 VDD1.n1 VDD1.t3 7.96741
R1047 VDD1 VDD1.n5 0.968172
C0 VN VTAIL 3.81522f
C1 B VDD2 1.3478f
C2 VN VP 5.52742f
C3 VN VDD1 0.155265f
C4 w_n3350_n1784# VN 6.52089f
C5 VN VDD2 3.09499f
C6 VN B 1.02862f
C7 VTAIL VP 3.82933f
C8 VTAIL VDD1 5.0449f
C9 VP VDD1 3.40418f
C10 w_n3350_n1784# VTAIL 2.34338f
C11 w_n3350_n1784# VP 6.95337f
C12 w_n3350_n1784# VDD1 1.56125f
C13 VTAIL VDD2 5.09563f
C14 VP VDD2 0.466204f
C15 VDD2 VDD1 1.4908f
C16 VTAIL B 2.18061f
C17 B VP 1.75182f
C18 B VDD1 1.26895f
C19 w_n3350_n1784# VDD2 1.65253f
C20 w_n3350_n1784# B 7.06583f
C21 VDD2 VSUBS 1.344111f
C22 VDD1 VSUBS 1.896425f
C23 VTAIL VSUBS 0.589288f
C24 VN VSUBS 5.74435f
C25 VP VSUBS 2.514303f
C26 B VSUBS 3.50689f
C27 w_n3350_n1784# VSUBS 75.2142f
C28 VDD1.t0 VSUBS 0.079725f
C29 VDD1.t7 VSUBS 0.079725f
C30 VDD1.n0 VSUBS 0.474662f
C31 VDD1.t2 VSUBS 0.079725f
C32 VDD1.t3 VSUBS 0.079725f
C33 VDD1.n1 VSUBS 0.47394f
C34 VDD1.t1 VSUBS 0.079725f
C35 VDD1.t6 VSUBS 0.079725f
C36 VDD1.n2 VSUBS 0.47394f
C37 VDD1.n3 VSUBS 2.80412f
C38 VDD1.t5 VSUBS 0.079725f
C39 VDD1.t4 VSUBS 0.079725f
C40 VDD1.n4 VSUBS 0.468458f
C41 VDD1.n5 VSUBS 2.29693f
C42 VP.n0 VSUBS 0.062432f
C43 VP.t1 VSUBS 1.01936f
C44 VP.n1 VSUBS 0.049539f
C45 VP.n2 VSUBS 0.047357f
C46 VP.t6 VSUBS 1.01936f
C47 VP.n3 VSUBS 0.068841f
C48 VP.n4 VSUBS 0.047357f
C49 VP.t4 VSUBS 1.01936f
C50 VP.n5 VSUBS 0.092337f
C51 VP.n6 VSUBS 0.047357f
C52 VP.t5 VSUBS 1.01936f
C53 VP.n7 VSUBS 0.549932f
C54 VP.n8 VSUBS 0.062432f
C55 VP.t3 VSUBS 1.01936f
C56 VP.n9 VSUBS 0.049539f
C57 VP.n10 VSUBS 0.047357f
C58 VP.t2 VSUBS 1.01936f
C59 VP.n11 VSUBS 0.068841f
C60 VP.n12 VSUBS 0.396346f
C61 VP.t0 VSUBS 1.01936f
C62 VP.t7 VSUBS 1.28834f
C63 VP.n13 VSUBS 0.511327f
C64 VP.n14 VSUBS 0.546238f
C65 VP.n15 VSUBS 0.082617f
C66 VP.n16 VSUBS 0.068841f
C67 VP.n17 VSUBS 0.047357f
C68 VP.n18 VSUBS 0.047357f
C69 VP.n19 VSUBS 0.047357f
C70 VP.n20 VSUBS 0.082617f
C71 VP.n21 VSUBS 0.413369f
C72 VP.n22 VSUBS 0.049668f
C73 VP.n23 VSUBS 0.092337f
C74 VP.n24 VSUBS 0.047357f
C75 VP.n25 VSUBS 0.047357f
C76 VP.n26 VSUBS 0.047357f
C77 VP.n27 VSUBS 0.083625f
C78 VP.n28 VSUBS 0.072212f
C79 VP.n29 VSUBS 0.549932f
C80 VP.n30 VSUBS 2.02197f
C81 VP.n31 VSUBS 2.06234f
C82 VP.n32 VSUBS 0.062432f
C83 VP.n33 VSUBS 0.072212f
C84 VP.n34 VSUBS 0.083625f
C85 VP.n35 VSUBS 0.049539f
C86 VP.n36 VSUBS 0.047357f
C87 VP.n37 VSUBS 0.047357f
C88 VP.n38 VSUBS 0.047357f
C89 VP.n39 VSUBS 0.049668f
C90 VP.n40 VSUBS 0.413369f
C91 VP.n41 VSUBS 0.082617f
C92 VP.n42 VSUBS 0.068841f
C93 VP.n43 VSUBS 0.047357f
C94 VP.n44 VSUBS 0.047357f
C95 VP.n45 VSUBS 0.047357f
C96 VP.n46 VSUBS 0.082617f
C97 VP.n47 VSUBS 0.413369f
C98 VP.n48 VSUBS 0.049668f
C99 VP.n49 VSUBS 0.092337f
C100 VP.n50 VSUBS 0.047357f
C101 VP.n51 VSUBS 0.047357f
C102 VP.n52 VSUBS 0.047357f
C103 VP.n53 VSUBS 0.083625f
C104 VP.n54 VSUBS 0.072212f
C105 VP.n55 VSUBS 0.549932f
C106 VP.n56 VSUBS 0.063168f
C107 B.n0 VSUBS 0.005812f
C108 B.n1 VSUBS 0.005812f
C109 B.n2 VSUBS 0.00919f
C110 B.n3 VSUBS 0.00919f
C111 B.n4 VSUBS 0.00919f
C112 B.n5 VSUBS 0.00919f
C113 B.n6 VSUBS 0.00919f
C114 B.n7 VSUBS 0.00919f
C115 B.n8 VSUBS 0.00919f
C116 B.n9 VSUBS 0.00919f
C117 B.n10 VSUBS 0.00919f
C118 B.n11 VSUBS 0.00919f
C119 B.n12 VSUBS 0.00919f
C120 B.n13 VSUBS 0.00919f
C121 B.n14 VSUBS 0.00919f
C122 B.n15 VSUBS 0.00919f
C123 B.n16 VSUBS 0.00919f
C124 B.n17 VSUBS 0.00919f
C125 B.n18 VSUBS 0.00919f
C126 B.n19 VSUBS 0.00919f
C127 B.n20 VSUBS 0.00919f
C128 B.n21 VSUBS 0.00919f
C129 B.n22 VSUBS 0.00919f
C130 B.n23 VSUBS 0.021951f
C131 B.n24 VSUBS 0.00919f
C132 B.n25 VSUBS 0.00919f
C133 B.n26 VSUBS 0.00919f
C134 B.n27 VSUBS 0.00919f
C135 B.n28 VSUBS 0.00919f
C136 B.n29 VSUBS 0.00919f
C137 B.n30 VSUBS 0.00919f
C138 B.n31 VSUBS 0.00919f
C139 B.n32 VSUBS 0.00865f
C140 B.n33 VSUBS 0.00919f
C141 B.t8 VSUBS 0.141841f
C142 B.t7 VSUBS 0.162456f
C143 B.t6 VSUBS 0.522932f
C144 B.n34 VSUBS 0.114746f
C145 B.n35 VSUBS 0.086911f
C146 B.n36 VSUBS 0.021293f
C147 B.n37 VSUBS 0.00919f
C148 B.n38 VSUBS 0.00919f
C149 B.n39 VSUBS 0.00919f
C150 B.n40 VSUBS 0.00919f
C151 B.t2 VSUBS 0.141841f
C152 B.t1 VSUBS 0.162456f
C153 B.t0 VSUBS 0.522932f
C154 B.n41 VSUBS 0.114746f
C155 B.n42 VSUBS 0.086911f
C156 B.n43 VSUBS 0.00919f
C157 B.n44 VSUBS 0.00919f
C158 B.n45 VSUBS 0.00919f
C159 B.n46 VSUBS 0.00919f
C160 B.n47 VSUBS 0.00919f
C161 B.n48 VSUBS 0.00919f
C162 B.n49 VSUBS 0.00919f
C163 B.n50 VSUBS 0.00919f
C164 B.n51 VSUBS 0.021901f
C165 B.n52 VSUBS 0.00919f
C166 B.n53 VSUBS 0.00919f
C167 B.n54 VSUBS 0.00919f
C168 B.n55 VSUBS 0.00919f
C169 B.n56 VSUBS 0.00919f
C170 B.n57 VSUBS 0.00919f
C171 B.n58 VSUBS 0.00919f
C172 B.n59 VSUBS 0.00919f
C173 B.n60 VSUBS 0.00919f
C174 B.n61 VSUBS 0.00919f
C175 B.n62 VSUBS 0.00919f
C176 B.n63 VSUBS 0.00919f
C177 B.n64 VSUBS 0.00919f
C178 B.n65 VSUBS 0.00919f
C179 B.n66 VSUBS 0.00919f
C180 B.n67 VSUBS 0.00919f
C181 B.n68 VSUBS 0.00919f
C182 B.n69 VSUBS 0.00919f
C183 B.n70 VSUBS 0.00919f
C184 B.n71 VSUBS 0.00919f
C185 B.n72 VSUBS 0.00919f
C186 B.n73 VSUBS 0.00919f
C187 B.n74 VSUBS 0.00919f
C188 B.n75 VSUBS 0.00919f
C189 B.n76 VSUBS 0.00919f
C190 B.n77 VSUBS 0.00919f
C191 B.n78 VSUBS 0.00919f
C192 B.n79 VSUBS 0.00919f
C193 B.n80 VSUBS 0.00919f
C194 B.n81 VSUBS 0.00919f
C195 B.n82 VSUBS 0.00919f
C196 B.n83 VSUBS 0.00919f
C197 B.n84 VSUBS 0.00919f
C198 B.n85 VSUBS 0.00919f
C199 B.n86 VSUBS 0.00919f
C200 B.n87 VSUBS 0.00919f
C201 B.n88 VSUBS 0.00919f
C202 B.n89 VSUBS 0.00919f
C203 B.n90 VSUBS 0.00919f
C204 B.n91 VSUBS 0.00919f
C205 B.n92 VSUBS 0.00919f
C206 B.n93 VSUBS 0.00919f
C207 B.n94 VSUBS 0.00919f
C208 B.n95 VSUBS 0.02292f
C209 B.n96 VSUBS 0.00919f
C210 B.n97 VSUBS 0.00919f
C211 B.n98 VSUBS 0.00919f
C212 B.n99 VSUBS 0.00919f
C213 B.n100 VSUBS 0.00919f
C214 B.n101 VSUBS 0.00919f
C215 B.n102 VSUBS 0.00919f
C216 B.n103 VSUBS 0.00919f
C217 B.n104 VSUBS 0.00919f
C218 B.t10 VSUBS 0.141841f
C219 B.t11 VSUBS 0.162456f
C220 B.t9 VSUBS 0.522932f
C221 B.n105 VSUBS 0.114746f
C222 B.n106 VSUBS 0.086911f
C223 B.n107 VSUBS 0.00919f
C224 B.n108 VSUBS 0.00919f
C225 B.n109 VSUBS 0.00919f
C226 B.n110 VSUBS 0.00919f
C227 B.t4 VSUBS 0.141841f
C228 B.t5 VSUBS 0.162456f
C229 B.t3 VSUBS 0.522932f
C230 B.n111 VSUBS 0.114746f
C231 B.n112 VSUBS 0.086911f
C232 B.n113 VSUBS 0.021293f
C233 B.n114 VSUBS 0.00919f
C234 B.n115 VSUBS 0.00919f
C235 B.n116 VSUBS 0.00919f
C236 B.n117 VSUBS 0.00919f
C237 B.n118 VSUBS 0.00919f
C238 B.n119 VSUBS 0.00919f
C239 B.n120 VSUBS 0.00919f
C240 B.n121 VSUBS 0.00919f
C241 B.n122 VSUBS 0.02292f
C242 B.n123 VSUBS 0.00919f
C243 B.n124 VSUBS 0.00919f
C244 B.n125 VSUBS 0.00919f
C245 B.n126 VSUBS 0.00919f
C246 B.n127 VSUBS 0.00919f
C247 B.n128 VSUBS 0.00919f
C248 B.n129 VSUBS 0.00919f
C249 B.n130 VSUBS 0.00919f
C250 B.n131 VSUBS 0.00919f
C251 B.n132 VSUBS 0.00919f
C252 B.n133 VSUBS 0.00919f
C253 B.n134 VSUBS 0.00919f
C254 B.n135 VSUBS 0.00919f
C255 B.n136 VSUBS 0.00919f
C256 B.n137 VSUBS 0.00919f
C257 B.n138 VSUBS 0.00919f
C258 B.n139 VSUBS 0.00919f
C259 B.n140 VSUBS 0.00919f
C260 B.n141 VSUBS 0.00919f
C261 B.n142 VSUBS 0.00919f
C262 B.n143 VSUBS 0.00919f
C263 B.n144 VSUBS 0.00919f
C264 B.n145 VSUBS 0.00919f
C265 B.n146 VSUBS 0.00919f
C266 B.n147 VSUBS 0.00919f
C267 B.n148 VSUBS 0.00919f
C268 B.n149 VSUBS 0.00919f
C269 B.n150 VSUBS 0.00919f
C270 B.n151 VSUBS 0.00919f
C271 B.n152 VSUBS 0.00919f
C272 B.n153 VSUBS 0.00919f
C273 B.n154 VSUBS 0.00919f
C274 B.n155 VSUBS 0.00919f
C275 B.n156 VSUBS 0.00919f
C276 B.n157 VSUBS 0.00919f
C277 B.n158 VSUBS 0.00919f
C278 B.n159 VSUBS 0.00919f
C279 B.n160 VSUBS 0.00919f
C280 B.n161 VSUBS 0.00919f
C281 B.n162 VSUBS 0.00919f
C282 B.n163 VSUBS 0.00919f
C283 B.n164 VSUBS 0.00919f
C284 B.n165 VSUBS 0.00919f
C285 B.n166 VSUBS 0.00919f
C286 B.n167 VSUBS 0.00919f
C287 B.n168 VSUBS 0.00919f
C288 B.n169 VSUBS 0.00919f
C289 B.n170 VSUBS 0.00919f
C290 B.n171 VSUBS 0.00919f
C291 B.n172 VSUBS 0.00919f
C292 B.n173 VSUBS 0.00919f
C293 B.n174 VSUBS 0.00919f
C294 B.n175 VSUBS 0.00919f
C295 B.n176 VSUBS 0.00919f
C296 B.n177 VSUBS 0.00919f
C297 B.n178 VSUBS 0.00919f
C298 B.n179 VSUBS 0.00919f
C299 B.n180 VSUBS 0.00919f
C300 B.n181 VSUBS 0.00919f
C301 B.n182 VSUBS 0.00919f
C302 B.n183 VSUBS 0.00919f
C303 B.n184 VSUBS 0.00919f
C304 B.n185 VSUBS 0.00919f
C305 B.n186 VSUBS 0.00919f
C306 B.n187 VSUBS 0.00919f
C307 B.n188 VSUBS 0.00919f
C308 B.n189 VSUBS 0.00919f
C309 B.n190 VSUBS 0.00919f
C310 B.n191 VSUBS 0.00919f
C311 B.n192 VSUBS 0.00919f
C312 B.n193 VSUBS 0.00919f
C313 B.n194 VSUBS 0.00919f
C314 B.n195 VSUBS 0.00919f
C315 B.n196 VSUBS 0.00919f
C316 B.n197 VSUBS 0.00919f
C317 B.n198 VSUBS 0.00919f
C318 B.n199 VSUBS 0.00919f
C319 B.n200 VSUBS 0.00919f
C320 B.n201 VSUBS 0.00919f
C321 B.n202 VSUBS 0.00919f
C322 B.n203 VSUBS 0.00919f
C323 B.n204 VSUBS 0.00919f
C324 B.n205 VSUBS 0.021951f
C325 B.n206 VSUBS 0.021951f
C326 B.n207 VSUBS 0.02292f
C327 B.n208 VSUBS 0.00919f
C328 B.n209 VSUBS 0.00919f
C329 B.n210 VSUBS 0.00919f
C330 B.n211 VSUBS 0.00919f
C331 B.n212 VSUBS 0.00919f
C332 B.n213 VSUBS 0.00919f
C333 B.n214 VSUBS 0.00919f
C334 B.n215 VSUBS 0.00919f
C335 B.n216 VSUBS 0.00919f
C336 B.n217 VSUBS 0.00919f
C337 B.n218 VSUBS 0.00919f
C338 B.n219 VSUBS 0.00919f
C339 B.n220 VSUBS 0.00919f
C340 B.n221 VSUBS 0.00919f
C341 B.n222 VSUBS 0.00919f
C342 B.n223 VSUBS 0.00919f
C343 B.n224 VSUBS 0.00919f
C344 B.n225 VSUBS 0.00919f
C345 B.n226 VSUBS 0.00919f
C346 B.n227 VSUBS 0.00919f
C347 B.n228 VSUBS 0.00919f
C348 B.n229 VSUBS 0.00919f
C349 B.n230 VSUBS 0.00919f
C350 B.n231 VSUBS 0.00919f
C351 B.n232 VSUBS 0.00865f
C352 B.n233 VSUBS 0.00919f
C353 B.n234 VSUBS 0.00919f
C354 B.n235 VSUBS 0.005136f
C355 B.n236 VSUBS 0.00919f
C356 B.n237 VSUBS 0.00919f
C357 B.n238 VSUBS 0.00919f
C358 B.n239 VSUBS 0.00919f
C359 B.n240 VSUBS 0.00919f
C360 B.n241 VSUBS 0.00919f
C361 B.n242 VSUBS 0.00919f
C362 B.n243 VSUBS 0.00919f
C363 B.n244 VSUBS 0.00919f
C364 B.n245 VSUBS 0.00919f
C365 B.n246 VSUBS 0.00919f
C366 B.n247 VSUBS 0.00919f
C367 B.n248 VSUBS 0.005136f
C368 B.n249 VSUBS 0.021293f
C369 B.n250 VSUBS 0.00865f
C370 B.n251 VSUBS 0.00919f
C371 B.n252 VSUBS 0.00919f
C372 B.n253 VSUBS 0.00919f
C373 B.n254 VSUBS 0.00919f
C374 B.n255 VSUBS 0.00919f
C375 B.n256 VSUBS 0.00919f
C376 B.n257 VSUBS 0.00919f
C377 B.n258 VSUBS 0.00919f
C378 B.n259 VSUBS 0.00919f
C379 B.n260 VSUBS 0.00919f
C380 B.n261 VSUBS 0.00919f
C381 B.n262 VSUBS 0.00919f
C382 B.n263 VSUBS 0.00919f
C383 B.n264 VSUBS 0.00919f
C384 B.n265 VSUBS 0.00919f
C385 B.n266 VSUBS 0.00919f
C386 B.n267 VSUBS 0.00919f
C387 B.n268 VSUBS 0.00919f
C388 B.n269 VSUBS 0.00919f
C389 B.n270 VSUBS 0.00919f
C390 B.n271 VSUBS 0.00919f
C391 B.n272 VSUBS 0.00919f
C392 B.n273 VSUBS 0.00919f
C393 B.n274 VSUBS 0.00919f
C394 B.n275 VSUBS 0.00919f
C395 B.n276 VSUBS 0.02292f
C396 B.n277 VSUBS 0.021951f
C397 B.n278 VSUBS 0.021951f
C398 B.n279 VSUBS 0.00919f
C399 B.n280 VSUBS 0.00919f
C400 B.n281 VSUBS 0.00919f
C401 B.n282 VSUBS 0.00919f
C402 B.n283 VSUBS 0.00919f
C403 B.n284 VSUBS 0.00919f
C404 B.n285 VSUBS 0.00919f
C405 B.n286 VSUBS 0.00919f
C406 B.n287 VSUBS 0.00919f
C407 B.n288 VSUBS 0.00919f
C408 B.n289 VSUBS 0.00919f
C409 B.n290 VSUBS 0.00919f
C410 B.n291 VSUBS 0.00919f
C411 B.n292 VSUBS 0.00919f
C412 B.n293 VSUBS 0.00919f
C413 B.n294 VSUBS 0.00919f
C414 B.n295 VSUBS 0.00919f
C415 B.n296 VSUBS 0.00919f
C416 B.n297 VSUBS 0.00919f
C417 B.n298 VSUBS 0.00919f
C418 B.n299 VSUBS 0.00919f
C419 B.n300 VSUBS 0.00919f
C420 B.n301 VSUBS 0.00919f
C421 B.n302 VSUBS 0.00919f
C422 B.n303 VSUBS 0.00919f
C423 B.n304 VSUBS 0.00919f
C424 B.n305 VSUBS 0.00919f
C425 B.n306 VSUBS 0.00919f
C426 B.n307 VSUBS 0.00919f
C427 B.n308 VSUBS 0.00919f
C428 B.n309 VSUBS 0.00919f
C429 B.n310 VSUBS 0.00919f
C430 B.n311 VSUBS 0.00919f
C431 B.n312 VSUBS 0.00919f
C432 B.n313 VSUBS 0.00919f
C433 B.n314 VSUBS 0.00919f
C434 B.n315 VSUBS 0.00919f
C435 B.n316 VSUBS 0.00919f
C436 B.n317 VSUBS 0.00919f
C437 B.n318 VSUBS 0.00919f
C438 B.n319 VSUBS 0.00919f
C439 B.n320 VSUBS 0.00919f
C440 B.n321 VSUBS 0.00919f
C441 B.n322 VSUBS 0.00919f
C442 B.n323 VSUBS 0.00919f
C443 B.n324 VSUBS 0.00919f
C444 B.n325 VSUBS 0.00919f
C445 B.n326 VSUBS 0.00919f
C446 B.n327 VSUBS 0.00919f
C447 B.n328 VSUBS 0.00919f
C448 B.n329 VSUBS 0.00919f
C449 B.n330 VSUBS 0.00919f
C450 B.n331 VSUBS 0.00919f
C451 B.n332 VSUBS 0.00919f
C452 B.n333 VSUBS 0.00919f
C453 B.n334 VSUBS 0.00919f
C454 B.n335 VSUBS 0.00919f
C455 B.n336 VSUBS 0.00919f
C456 B.n337 VSUBS 0.00919f
C457 B.n338 VSUBS 0.00919f
C458 B.n339 VSUBS 0.00919f
C459 B.n340 VSUBS 0.00919f
C460 B.n341 VSUBS 0.00919f
C461 B.n342 VSUBS 0.00919f
C462 B.n343 VSUBS 0.00919f
C463 B.n344 VSUBS 0.00919f
C464 B.n345 VSUBS 0.00919f
C465 B.n346 VSUBS 0.00919f
C466 B.n347 VSUBS 0.00919f
C467 B.n348 VSUBS 0.00919f
C468 B.n349 VSUBS 0.00919f
C469 B.n350 VSUBS 0.00919f
C470 B.n351 VSUBS 0.00919f
C471 B.n352 VSUBS 0.00919f
C472 B.n353 VSUBS 0.00919f
C473 B.n354 VSUBS 0.00919f
C474 B.n355 VSUBS 0.00919f
C475 B.n356 VSUBS 0.00919f
C476 B.n357 VSUBS 0.00919f
C477 B.n358 VSUBS 0.00919f
C478 B.n359 VSUBS 0.00919f
C479 B.n360 VSUBS 0.00919f
C480 B.n361 VSUBS 0.00919f
C481 B.n362 VSUBS 0.00919f
C482 B.n363 VSUBS 0.00919f
C483 B.n364 VSUBS 0.00919f
C484 B.n365 VSUBS 0.00919f
C485 B.n366 VSUBS 0.00919f
C486 B.n367 VSUBS 0.00919f
C487 B.n368 VSUBS 0.00919f
C488 B.n369 VSUBS 0.00919f
C489 B.n370 VSUBS 0.00919f
C490 B.n371 VSUBS 0.00919f
C491 B.n372 VSUBS 0.00919f
C492 B.n373 VSUBS 0.00919f
C493 B.n374 VSUBS 0.00919f
C494 B.n375 VSUBS 0.00919f
C495 B.n376 VSUBS 0.00919f
C496 B.n377 VSUBS 0.00919f
C497 B.n378 VSUBS 0.00919f
C498 B.n379 VSUBS 0.00919f
C499 B.n380 VSUBS 0.00919f
C500 B.n381 VSUBS 0.00919f
C501 B.n382 VSUBS 0.00919f
C502 B.n383 VSUBS 0.00919f
C503 B.n384 VSUBS 0.00919f
C504 B.n385 VSUBS 0.00919f
C505 B.n386 VSUBS 0.00919f
C506 B.n387 VSUBS 0.00919f
C507 B.n388 VSUBS 0.00919f
C508 B.n389 VSUBS 0.00919f
C509 B.n390 VSUBS 0.00919f
C510 B.n391 VSUBS 0.00919f
C511 B.n392 VSUBS 0.00919f
C512 B.n393 VSUBS 0.00919f
C513 B.n394 VSUBS 0.00919f
C514 B.n395 VSUBS 0.00919f
C515 B.n396 VSUBS 0.00919f
C516 B.n397 VSUBS 0.00919f
C517 B.n398 VSUBS 0.00919f
C518 B.n399 VSUBS 0.00919f
C519 B.n400 VSUBS 0.00919f
C520 B.n401 VSUBS 0.00919f
C521 B.n402 VSUBS 0.00919f
C522 B.n403 VSUBS 0.00919f
C523 B.n404 VSUBS 0.00919f
C524 B.n405 VSUBS 0.00919f
C525 B.n406 VSUBS 0.02297f
C526 B.n407 VSUBS 0.021951f
C527 B.n408 VSUBS 0.02292f
C528 B.n409 VSUBS 0.00919f
C529 B.n410 VSUBS 0.00919f
C530 B.n411 VSUBS 0.00919f
C531 B.n412 VSUBS 0.00919f
C532 B.n413 VSUBS 0.00919f
C533 B.n414 VSUBS 0.00919f
C534 B.n415 VSUBS 0.00919f
C535 B.n416 VSUBS 0.00919f
C536 B.n417 VSUBS 0.00919f
C537 B.n418 VSUBS 0.00919f
C538 B.n419 VSUBS 0.00919f
C539 B.n420 VSUBS 0.00919f
C540 B.n421 VSUBS 0.00919f
C541 B.n422 VSUBS 0.00919f
C542 B.n423 VSUBS 0.00919f
C543 B.n424 VSUBS 0.00919f
C544 B.n425 VSUBS 0.00919f
C545 B.n426 VSUBS 0.00919f
C546 B.n427 VSUBS 0.00919f
C547 B.n428 VSUBS 0.00919f
C548 B.n429 VSUBS 0.00919f
C549 B.n430 VSUBS 0.00919f
C550 B.n431 VSUBS 0.00919f
C551 B.n432 VSUBS 0.00919f
C552 B.n433 VSUBS 0.00919f
C553 B.n434 VSUBS 0.00865f
C554 B.n435 VSUBS 0.021293f
C555 B.n436 VSUBS 0.005136f
C556 B.n437 VSUBS 0.00919f
C557 B.n438 VSUBS 0.00919f
C558 B.n439 VSUBS 0.00919f
C559 B.n440 VSUBS 0.00919f
C560 B.n441 VSUBS 0.00919f
C561 B.n442 VSUBS 0.00919f
C562 B.n443 VSUBS 0.00919f
C563 B.n444 VSUBS 0.00919f
C564 B.n445 VSUBS 0.00919f
C565 B.n446 VSUBS 0.00919f
C566 B.n447 VSUBS 0.00919f
C567 B.n448 VSUBS 0.00919f
C568 B.n449 VSUBS 0.005136f
C569 B.n450 VSUBS 0.00919f
C570 B.n451 VSUBS 0.00919f
C571 B.n452 VSUBS 0.00919f
C572 B.n453 VSUBS 0.00919f
C573 B.n454 VSUBS 0.00919f
C574 B.n455 VSUBS 0.00919f
C575 B.n456 VSUBS 0.00919f
C576 B.n457 VSUBS 0.00919f
C577 B.n458 VSUBS 0.00919f
C578 B.n459 VSUBS 0.00919f
C579 B.n460 VSUBS 0.00919f
C580 B.n461 VSUBS 0.00919f
C581 B.n462 VSUBS 0.00919f
C582 B.n463 VSUBS 0.00919f
C583 B.n464 VSUBS 0.00919f
C584 B.n465 VSUBS 0.00919f
C585 B.n466 VSUBS 0.00919f
C586 B.n467 VSUBS 0.00919f
C587 B.n468 VSUBS 0.00919f
C588 B.n469 VSUBS 0.00919f
C589 B.n470 VSUBS 0.00919f
C590 B.n471 VSUBS 0.00919f
C591 B.n472 VSUBS 0.00919f
C592 B.n473 VSUBS 0.00919f
C593 B.n474 VSUBS 0.00919f
C594 B.n475 VSUBS 0.00919f
C595 B.n476 VSUBS 0.02292f
C596 B.n477 VSUBS 0.02292f
C597 B.n478 VSUBS 0.021951f
C598 B.n479 VSUBS 0.00919f
C599 B.n480 VSUBS 0.00919f
C600 B.n481 VSUBS 0.00919f
C601 B.n482 VSUBS 0.00919f
C602 B.n483 VSUBS 0.00919f
C603 B.n484 VSUBS 0.00919f
C604 B.n485 VSUBS 0.00919f
C605 B.n486 VSUBS 0.00919f
C606 B.n487 VSUBS 0.00919f
C607 B.n488 VSUBS 0.00919f
C608 B.n489 VSUBS 0.00919f
C609 B.n490 VSUBS 0.00919f
C610 B.n491 VSUBS 0.00919f
C611 B.n492 VSUBS 0.00919f
C612 B.n493 VSUBS 0.00919f
C613 B.n494 VSUBS 0.00919f
C614 B.n495 VSUBS 0.00919f
C615 B.n496 VSUBS 0.00919f
C616 B.n497 VSUBS 0.00919f
C617 B.n498 VSUBS 0.00919f
C618 B.n499 VSUBS 0.00919f
C619 B.n500 VSUBS 0.00919f
C620 B.n501 VSUBS 0.00919f
C621 B.n502 VSUBS 0.00919f
C622 B.n503 VSUBS 0.00919f
C623 B.n504 VSUBS 0.00919f
C624 B.n505 VSUBS 0.00919f
C625 B.n506 VSUBS 0.00919f
C626 B.n507 VSUBS 0.00919f
C627 B.n508 VSUBS 0.00919f
C628 B.n509 VSUBS 0.00919f
C629 B.n510 VSUBS 0.00919f
C630 B.n511 VSUBS 0.00919f
C631 B.n512 VSUBS 0.00919f
C632 B.n513 VSUBS 0.00919f
C633 B.n514 VSUBS 0.00919f
C634 B.n515 VSUBS 0.00919f
C635 B.n516 VSUBS 0.00919f
C636 B.n517 VSUBS 0.00919f
C637 B.n518 VSUBS 0.00919f
C638 B.n519 VSUBS 0.00919f
C639 B.n520 VSUBS 0.00919f
C640 B.n521 VSUBS 0.00919f
C641 B.n522 VSUBS 0.00919f
C642 B.n523 VSUBS 0.00919f
C643 B.n524 VSUBS 0.00919f
C644 B.n525 VSUBS 0.00919f
C645 B.n526 VSUBS 0.00919f
C646 B.n527 VSUBS 0.00919f
C647 B.n528 VSUBS 0.00919f
C648 B.n529 VSUBS 0.00919f
C649 B.n530 VSUBS 0.00919f
C650 B.n531 VSUBS 0.00919f
C651 B.n532 VSUBS 0.00919f
C652 B.n533 VSUBS 0.00919f
C653 B.n534 VSUBS 0.00919f
C654 B.n535 VSUBS 0.00919f
C655 B.n536 VSUBS 0.00919f
C656 B.n537 VSUBS 0.00919f
C657 B.n538 VSUBS 0.00919f
C658 B.n539 VSUBS 0.00919f
C659 B.n540 VSUBS 0.00919f
C660 B.n541 VSUBS 0.00919f
C661 B.n542 VSUBS 0.00919f
C662 B.n543 VSUBS 0.02081f
C663 VTAIL.t11 VSUBS 0.099904f
C664 VTAIL.t10 VSUBS 0.099904f
C665 VTAIL.n0 VSUBS 0.50557f
C666 VTAIL.n1 VSUBS 0.692424f
C667 VTAIL.t14 VSUBS 0.722537f
C668 VTAIL.n2 VSUBS 0.789023f
C669 VTAIL.t15 VSUBS 0.722537f
C670 VTAIL.n3 VSUBS 0.789023f
C671 VTAIL.t1 VSUBS 0.099904f
C672 VTAIL.t6 VSUBS 0.099904f
C673 VTAIL.n4 VSUBS 0.50557f
C674 VTAIL.n5 VSUBS 0.891468f
C675 VTAIL.t0 VSUBS 0.722537f
C676 VTAIL.n6 VSUBS 1.71906f
C677 VTAIL.t13 VSUBS 0.72254f
C678 VTAIL.n7 VSUBS 1.71905f
C679 VTAIL.t7 VSUBS 0.099904f
C680 VTAIL.t9 VSUBS 0.099904f
C681 VTAIL.n8 VSUBS 0.505574f
C682 VTAIL.n9 VSUBS 0.891465f
C683 VTAIL.t12 VSUBS 0.72254f
C684 VTAIL.n10 VSUBS 0.78902f
C685 VTAIL.t4 VSUBS 0.72254f
C686 VTAIL.n11 VSUBS 0.78902f
C687 VTAIL.t3 VSUBS 0.099904f
C688 VTAIL.t5 VSUBS 0.099904f
C689 VTAIL.n12 VSUBS 0.505574f
C690 VTAIL.n13 VSUBS 0.891465f
C691 VTAIL.t2 VSUBS 0.722537f
C692 VTAIL.n14 VSUBS 1.71906f
C693 VTAIL.t8 VSUBS 0.722537f
C694 VTAIL.n15 VSUBS 1.71325f
C695 VDD2.t1 VSUBS 0.078683f
C696 VDD2.t6 VSUBS 0.078683f
C697 VDD2.n0 VSUBS 0.467741f
C698 VDD2.t4 VSUBS 0.078683f
C699 VDD2.t2 VSUBS 0.078683f
C700 VDD2.n1 VSUBS 0.467741f
C701 VDD2.n2 VSUBS 2.71608f
C702 VDD2.t0 VSUBS 0.078683f
C703 VDD2.t7 VSUBS 0.078683f
C704 VDD2.n3 VSUBS 0.462334f
C705 VDD2.n4 VSUBS 2.23727f
C706 VDD2.t3 VSUBS 0.078683f
C707 VDD2.t5 VSUBS 0.078683f
C708 VDD2.n5 VSUBS 0.467718f
C709 VN.n0 VSUBS 0.059695f
C710 VN.t6 VSUBS 0.974666f
C711 VN.n1 VSUBS 0.047367f
C712 VN.n2 VSUBS 0.045281f
C713 VN.t4 VSUBS 0.974666f
C714 VN.n3 VSUBS 0.065823f
C715 VN.n4 VSUBS 0.37897f
C716 VN.t3 VSUBS 0.974666f
C717 VN.t0 VSUBS 1.23185f
C718 VN.n5 VSUBS 0.48891f
C719 VN.n6 VSUBS 0.522291f
C720 VN.n7 VSUBS 0.078995f
C721 VN.n8 VSUBS 0.065823f
C722 VN.n9 VSUBS 0.045281f
C723 VN.n10 VSUBS 0.045281f
C724 VN.n11 VSUBS 0.045281f
C725 VN.n12 VSUBS 0.078995f
C726 VN.n13 VSUBS 0.395247f
C727 VN.n14 VSUBS 0.04749f
C728 VN.n15 VSUBS 0.088289f
C729 VN.n16 VSUBS 0.045281f
C730 VN.n17 VSUBS 0.045281f
C731 VN.n18 VSUBS 0.045281f
C732 VN.n19 VSUBS 0.079959f
C733 VN.n20 VSUBS 0.069046f
C734 VN.n21 VSUBS 0.525823f
C735 VN.n22 VSUBS 0.060399f
C736 VN.n23 VSUBS 0.059695f
C737 VN.t1 VSUBS 0.974666f
C738 VN.n24 VSUBS 0.047367f
C739 VN.n25 VSUBS 0.045281f
C740 VN.t7 VSUBS 0.974666f
C741 VN.n26 VSUBS 0.065823f
C742 VN.n27 VSUBS 0.37897f
C743 VN.t5 VSUBS 0.974666f
C744 VN.t2 VSUBS 1.23185f
C745 VN.n28 VSUBS 0.48891f
C746 VN.n29 VSUBS 0.522291f
C747 VN.n30 VSUBS 0.078995f
C748 VN.n31 VSUBS 0.065823f
C749 VN.n32 VSUBS 0.045281f
C750 VN.n33 VSUBS 0.045281f
C751 VN.n34 VSUBS 0.045281f
C752 VN.n35 VSUBS 0.078995f
C753 VN.n36 VSUBS 0.395247f
C754 VN.n37 VSUBS 0.04749f
C755 VN.n38 VSUBS 0.088289f
C756 VN.n39 VSUBS 0.045281f
C757 VN.n40 VSUBS 0.045281f
C758 VN.n41 VSUBS 0.045281f
C759 VN.n42 VSUBS 0.079959f
C760 VN.n43 VSUBS 0.069046f
C761 VN.n44 VSUBS 0.525823f
C762 VN.n45 VSUBS 1.95837f
.ends

