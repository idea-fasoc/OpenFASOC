* NGSPICE file created from diff_pair_sample_0310.ext - technology: sky130A

.subckt diff_pair_sample_0310 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.5148 pd=3.42 as=0.2178 ps=1.65 w=1.32 l=3.1
X1 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=0.5148 pd=3.42 as=0 ps=0 w=1.32 l=3.1
X2 VDD1.t1 VP.t1 VTAIL.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2178 pd=1.65 as=0.2178 ps=1.65 w=1.32 l=3.1
X3 VTAIL.t6 VN.t0 VDD2.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=0.2178 pd=1.65 as=0.2178 ps=1.65 w=1.32 l=3.1
X4 VDD1.t0 VP.t2 VTAIL.t13 B.t4 sky130_fd_pr__nfet_01v8 ad=0.2178 pd=1.65 as=0.5148 ps=3.42 w=1.32 l=3.1
X5 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=0.5148 pd=3.42 as=0 ps=0 w=1.32 l=3.1
X6 VTAIL.t12 VP.t3 VDD1.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5148 pd=3.42 as=0.2178 ps=1.65 w=1.32 l=3.1
X7 VTAIL.t5 VN.t1 VDD2.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5148 pd=3.42 as=0.2178 ps=1.65 w=1.32 l=3.1
X8 VDD1.t5 VP.t4 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2178 pd=1.65 as=0.5148 ps=3.42 w=1.32 l=3.1
X9 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=0.5148 pd=3.42 as=0 ps=0 w=1.32 l=3.1
X10 VTAIL.t10 VP.t5 VDD1.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=0.2178 pd=1.65 as=0.2178 ps=1.65 w=1.32 l=3.1
X11 VDD1.t6 VP.t6 VTAIL.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=0.2178 pd=1.65 as=0.2178 ps=1.65 w=1.32 l=3.1
X12 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.5148 pd=3.42 as=0 ps=0 w=1.32 l=3.1
X13 VTAIL.t2 VN.t2 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.2178 pd=1.65 as=0.2178 ps=1.65 w=1.32 l=3.1
X14 VDD2.t4 VN.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.2178 pd=1.65 as=0.5148 ps=3.42 w=1.32 l=3.1
X15 VDD2.t3 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2178 pd=1.65 as=0.2178 ps=1.65 w=1.32 l=3.1
X16 VDD2.t2 VN.t5 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.2178 pd=1.65 as=0.2178 ps=1.65 w=1.32 l=3.1
X17 VTAIL.t8 VP.t7 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.2178 pd=1.65 as=0.2178 ps=1.65 w=1.32 l=3.1
X18 VTAIL.t1 VN.t6 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.5148 pd=3.42 as=0.2178 ps=1.65 w=1.32 l=3.1
X19 VDD2.t0 VN.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2178 pd=1.65 as=0.5148 ps=3.42 w=1.32 l=3.1
R0 VP.n21 VP.n18 161.3
R1 VP.n23 VP.n22 161.3
R2 VP.n24 VP.n17 161.3
R3 VP.n26 VP.n25 161.3
R4 VP.n27 VP.n16 161.3
R5 VP.n29 VP.n28 161.3
R6 VP.n31 VP.n30 161.3
R7 VP.n32 VP.n14 161.3
R8 VP.n34 VP.n33 161.3
R9 VP.n35 VP.n13 161.3
R10 VP.n37 VP.n36 161.3
R11 VP.n38 VP.n12 161.3
R12 VP.n40 VP.n39 161.3
R13 VP.n75 VP.n74 161.3
R14 VP.n73 VP.n1 161.3
R15 VP.n72 VP.n71 161.3
R16 VP.n70 VP.n2 161.3
R17 VP.n69 VP.n68 161.3
R18 VP.n67 VP.n3 161.3
R19 VP.n66 VP.n65 161.3
R20 VP.n64 VP.n63 161.3
R21 VP.n62 VP.n5 161.3
R22 VP.n61 VP.n60 161.3
R23 VP.n59 VP.n6 161.3
R24 VP.n58 VP.n57 161.3
R25 VP.n56 VP.n7 161.3
R26 VP.n54 VP.n53 161.3
R27 VP.n52 VP.n8 161.3
R28 VP.n51 VP.n50 161.3
R29 VP.n49 VP.n9 161.3
R30 VP.n48 VP.n47 161.3
R31 VP.n46 VP.n10 161.3
R32 VP.n45 VP.n44 161.3
R33 VP.n43 VP.n42 70.818
R34 VP.n76 VP.n0 70.818
R35 VP.n41 VP.n11 70.818
R36 VP.n61 VP.n6 56.5617
R37 VP.n26 VP.n17 56.5617
R38 VP.n49 VP.n48 56.5617
R39 VP.n72 VP.n2 56.5617
R40 VP.n37 VP.n13 56.5617
R41 VP.n20 VP.n19 51.1977
R42 VP.n42 VP.n41 45.2799
R43 VP.n19 VP.t3 43.7243
R44 VP.n44 VP.n10 24.5923
R45 VP.n48 VP.n10 24.5923
R46 VP.n50 VP.n49 24.5923
R47 VP.n50 VP.n8 24.5923
R48 VP.n54 VP.n8 24.5923
R49 VP.n57 VP.n56 24.5923
R50 VP.n57 VP.n6 24.5923
R51 VP.n62 VP.n61 24.5923
R52 VP.n63 VP.n62 24.5923
R53 VP.n67 VP.n66 24.5923
R54 VP.n68 VP.n67 24.5923
R55 VP.n68 VP.n2 24.5923
R56 VP.n73 VP.n72 24.5923
R57 VP.n74 VP.n73 24.5923
R58 VP.n38 VP.n37 24.5923
R59 VP.n39 VP.n38 24.5923
R60 VP.n27 VP.n26 24.5923
R61 VP.n28 VP.n27 24.5923
R62 VP.n32 VP.n31 24.5923
R63 VP.n33 VP.n32 24.5923
R64 VP.n33 VP.n13 24.5923
R65 VP.n22 VP.n21 24.5923
R66 VP.n22 VP.n17 24.5923
R67 VP.n56 VP.n55 22.8709
R68 VP.n63 VP.n4 22.8709
R69 VP.n28 VP.n15 22.8709
R70 VP.n21 VP.n20 22.8709
R71 VP.n44 VP.n43 19.4281
R72 VP.n74 VP.n0 19.4281
R73 VP.n39 VP.n11 19.4281
R74 VP.n43 VP.t0 10.2624
R75 VP.n55 VP.t1 10.2624
R76 VP.n4 VP.t5 10.2624
R77 VP.n0 VP.t2 10.2624
R78 VP.n11 VP.t4 10.2624
R79 VP.n15 VP.t7 10.2624
R80 VP.n20 VP.t6 10.2624
R81 VP.n19 VP.n18 3.93217
R82 VP.n55 VP.n54 1.72193
R83 VP.n66 VP.n4 1.72193
R84 VP.n31 VP.n15 1.72193
R85 VP.n41 VP.n40 0.354861
R86 VP.n45 VP.n42 0.354861
R87 VP.n76 VP.n75 0.354861
R88 VP VP.n76 0.267071
R89 VP.n23 VP.n18 0.189894
R90 VP.n24 VP.n23 0.189894
R91 VP.n25 VP.n24 0.189894
R92 VP.n25 VP.n16 0.189894
R93 VP.n29 VP.n16 0.189894
R94 VP.n30 VP.n29 0.189894
R95 VP.n30 VP.n14 0.189894
R96 VP.n34 VP.n14 0.189894
R97 VP.n35 VP.n34 0.189894
R98 VP.n36 VP.n35 0.189894
R99 VP.n36 VP.n12 0.189894
R100 VP.n40 VP.n12 0.189894
R101 VP.n46 VP.n45 0.189894
R102 VP.n47 VP.n46 0.189894
R103 VP.n47 VP.n9 0.189894
R104 VP.n51 VP.n9 0.189894
R105 VP.n52 VP.n51 0.189894
R106 VP.n53 VP.n52 0.189894
R107 VP.n53 VP.n7 0.189894
R108 VP.n58 VP.n7 0.189894
R109 VP.n59 VP.n58 0.189894
R110 VP.n60 VP.n59 0.189894
R111 VP.n60 VP.n5 0.189894
R112 VP.n64 VP.n5 0.189894
R113 VP.n65 VP.n64 0.189894
R114 VP.n65 VP.n3 0.189894
R115 VP.n69 VP.n3 0.189894
R116 VP.n70 VP.n69 0.189894
R117 VP.n71 VP.n70 0.189894
R118 VP.n71 VP.n1 0.189894
R119 VP.n75 VP.n1 0.189894
R120 VDD1 VDD1.n0 148.74
R121 VDD1.n3 VDD1.n2 148.627
R122 VDD1.n3 VDD1.n1 148.627
R123 VDD1.n5 VDD1.n4 147.204
R124 VDD1.n5 VDD1.n3 38.7423
R125 VDD1.n4 VDD1.t4 15.0005
R126 VDD1.n4 VDD1.t5 15.0005
R127 VDD1.n0 VDD1.t2 15.0005
R128 VDD1.n0 VDD1.t6 15.0005
R129 VDD1.n2 VDD1.t7 15.0005
R130 VDD1.n2 VDD1.t0 15.0005
R131 VDD1.n1 VDD1.t3 15.0005
R132 VDD1.n1 VDD1.t1 15.0005
R133 VDD1 VDD1.n5 1.42076
R134 VTAIL.n15 VTAIL.t0 156.684
R135 VTAIL.n2 VTAIL.t5 156.684
R136 VTAIL.n3 VTAIL.t13 156.684
R137 VTAIL.n6 VTAIL.t15 156.684
R138 VTAIL.n14 VTAIL.t11 156.684
R139 VTAIL.n11 VTAIL.t12 156.684
R140 VTAIL.n10 VTAIL.t4 156.684
R141 VTAIL.n7 VTAIL.t1 156.684
R142 VTAIL.n1 VTAIL.n0 130.526
R143 VTAIL.n5 VTAIL.n4 130.526
R144 VTAIL.n13 VTAIL.n12 130.525
R145 VTAIL.n9 VTAIL.n8 130.525
R146 VTAIL.n15 VTAIL.n14 16.4617
R147 VTAIL.n7 VTAIL.n6 16.4617
R148 VTAIL.n0 VTAIL.t7 15.0005
R149 VTAIL.n0 VTAIL.t2 15.0005
R150 VTAIL.n4 VTAIL.t14 15.0005
R151 VTAIL.n4 VTAIL.t10 15.0005
R152 VTAIL.n12 VTAIL.t9 15.0005
R153 VTAIL.n12 VTAIL.t8 15.0005
R154 VTAIL.n8 VTAIL.t3 15.0005
R155 VTAIL.n8 VTAIL.t6 15.0005
R156 VTAIL.n9 VTAIL.n7 2.9574
R157 VTAIL.n10 VTAIL.n9 2.9574
R158 VTAIL.n13 VTAIL.n11 2.9574
R159 VTAIL.n14 VTAIL.n13 2.9574
R160 VTAIL.n6 VTAIL.n5 2.9574
R161 VTAIL.n5 VTAIL.n3 2.9574
R162 VTAIL.n2 VTAIL.n1 2.9574
R163 VTAIL VTAIL.n15 2.89921
R164 VTAIL.n11 VTAIL.n10 0.470328
R165 VTAIL.n3 VTAIL.n2 0.470328
R166 VTAIL VTAIL.n1 0.0586897
R167 B.n574 B.n573 585
R168 B.n575 B.n128 585
R169 B.n577 B.n576 585
R170 B.n579 B.n127 585
R171 B.n582 B.n581 585
R172 B.n583 B.n126 585
R173 B.n585 B.n584 585
R174 B.n587 B.n125 585
R175 B.n589 B.n588 585
R176 B.n591 B.n590 585
R177 B.n594 B.n593 585
R178 B.n595 B.n120 585
R179 B.n597 B.n596 585
R180 B.n599 B.n119 585
R181 B.n602 B.n601 585
R182 B.n603 B.n118 585
R183 B.n605 B.n604 585
R184 B.n607 B.n117 585
R185 B.n609 B.n608 585
R186 B.n611 B.n610 585
R187 B.n614 B.n613 585
R188 B.n615 B.n112 585
R189 B.n617 B.n616 585
R190 B.n619 B.n111 585
R191 B.n622 B.n621 585
R192 B.n623 B.n110 585
R193 B.n625 B.n624 585
R194 B.n627 B.n109 585
R195 B.n630 B.n629 585
R196 B.n631 B.n108 585
R197 B.n571 B.n106 585
R198 B.n634 B.n106 585
R199 B.n570 B.n105 585
R200 B.n635 B.n105 585
R201 B.n569 B.n104 585
R202 B.n636 B.n104 585
R203 B.n568 B.n567 585
R204 B.n567 B.n100 585
R205 B.n566 B.n99 585
R206 B.n642 B.n99 585
R207 B.n565 B.n98 585
R208 B.n643 B.n98 585
R209 B.n564 B.n97 585
R210 B.n644 B.n97 585
R211 B.n563 B.n562 585
R212 B.n562 B.n93 585
R213 B.n561 B.n92 585
R214 B.n650 B.n92 585
R215 B.n560 B.n91 585
R216 B.n651 B.n91 585
R217 B.n559 B.n90 585
R218 B.n652 B.n90 585
R219 B.n558 B.n557 585
R220 B.n557 B.n86 585
R221 B.n556 B.n85 585
R222 B.n658 B.n85 585
R223 B.n555 B.n84 585
R224 B.n659 B.n84 585
R225 B.n554 B.n83 585
R226 B.n660 B.n83 585
R227 B.n553 B.n552 585
R228 B.n552 B.n79 585
R229 B.n551 B.n78 585
R230 B.n666 B.n78 585
R231 B.n550 B.n77 585
R232 B.n667 B.n77 585
R233 B.n549 B.n76 585
R234 B.n668 B.n76 585
R235 B.n548 B.n547 585
R236 B.n547 B.n72 585
R237 B.n546 B.n71 585
R238 B.n674 B.n71 585
R239 B.n545 B.n70 585
R240 B.n675 B.n70 585
R241 B.n544 B.n69 585
R242 B.n676 B.n69 585
R243 B.n543 B.n542 585
R244 B.n542 B.n65 585
R245 B.n541 B.n64 585
R246 B.n682 B.n64 585
R247 B.n540 B.n63 585
R248 B.n683 B.n63 585
R249 B.n539 B.n62 585
R250 B.n684 B.n62 585
R251 B.n538 B.n537 585
R252 B.n537 B.n58 585
R253 B.n536 B.n57 585
R254 B.n690 B.n57 585
R255 B.n535 B.n56 585
R256 B.n691 B.n56 585
R257 B.n534 B.n55 585
R258 B.n692 B.n55 585
R259 B.n533 B.n532 585
R260 B.n532 B.n54 585
R261 B.n531 B.n50 585
R262 B.n698 B.n50 585
R263 B.n530 B.n49 585
R264 B.n699 B.n49 585
R265 B.n529 B.n48 585
R266 B.n700 B.n48 585
R267 B.n528 B.n527 585
R268 B.n527 B.n44 585
R269 B.n526 B.n43 585
R270 B.n706 B.n43 585
R271 B.n525 B.n42 585
R272 B.n707 B.n42 585
R273 B.n524 B.n41 585
R274 B.n708 B.n41 585
R275 B.n523 B.n522 585
R276 B.n522 B.n37 585
R277 B.n521 B.n36 585
R278 B.n714 B.n36 585
R279 B.n520 B.n35 585
R280 B.n715 B.n35 585
R281 B.n519 B.n34 585
R282 B.n716 B.n34 585
R283 B.n518 B.n517 585
R284 B.n517 B.n30 585
R285 B.n516 B.n29 585
R286 B.n722 B.n29 585
R287 B.n515 B.n28 585
R288 B.n723 B.n28 585
R289 B.n514 B.n27 585
R290 B.n724 B.n27 585
R291 B.n513 B.n512 585
R292 B.n512 B.n23 585
R293 B.n511 B.n22 585
R294 B.n730 B.n22 585
R295 B.n510 B.n21 585
R296 B.n731 B.n21 585
R297 B.n509 B.n20 585
R298 B.n732 B.n20 585
R299 B.n508 B.n507 585
R300 B.n507 B.n19 585
R301 B.n506 B.n15 585
R302 B.n738 B.n15 585
R303 B.n505 B.n14 585
R304 B.n739 B.n14 585
R305 B.n504 B.n13 585
R306 B.n740 B.n13 585
R307 B.n503 B.n502 585
R308 B.n502 B.n12 585
R309 B.n501 B.n500 585
R310 B.n501 B.n8 585
R311 B.n499 B.n7 585
R312 B.n747 B.n7 585
R313 B.n498 B.n6 585
R314 B.n748 B.n6 585
R315 B.n497 B.n5 585
R316 B.n749 B.n5 585
R317 B.n496 B.n495 585
R318 B.n495 B.n4 585
R319 B.n494 B.n129 585
R320 B.n494 B.n493 585
R321 B.n484 B.n130 585
R322 B.n131 B.n130 585
R323 B.n486 B.n485 585
R324 B.n487 B.n486 585
R325 B.n483 B.n136 585
R326 B.n136 B.n135 585
R327 B.n482 B.n481 585
R328 B.n481 B.n480 585
R329 B.n138 B.n137 585
R330 B.n473 B.n138 585
R331 B.n472 B.n471 585
R332 B.n474 B.n472 585
R333 B.n470 B.n143 585
R334 B.n143 B.n142 585
R335 B.n469 B.n468 585
R336 B.n468 B.n467 585
R337 B.n145 B.n144 585
R338 B.n146 B.n145 585
R339 B.n460 B.n459 585
R340 B.n461 B.n460 585
R341 B.n458 B.n151 585
R342 B.n151 B.n150 585
R343 B.n457 B.n456 585
R344 B.n456 B.n455 585
R345 B.n153 B.n152 585
R346 B.n154 B.n153 585
R347 B.n448 B.n447 585
R348 B.n449 B.n448 585
R349 B.n446 B.n158 585
R350 B.n162 B.n158 585
R351 B.n445 B.n444 585
R352 B.n444 B.n443 585
R353 B.n160 B.n159 585
R354 B.n161 B.n160 585
R355 B.n436 B.n435 585
R356 B.n437 B.n436 585
R357 B.n434 B.n167 585
R358 B.n167 B.n166 585
R359 B.n433 B.n432 585
R360 B.n432 B.n431 585
R361 B.n169 B.n168 585
R362 B.n170 B.n169 585
R363 B.n424 B.n423 585
R364 B.n425 B.n424 585
R365 B.n422 B.n175 585
R366 B.n175 B.n174 585
R367 B.n421 B.n420 585
R368 B.n420 B.n419 585
R369 B.n177 B.n176 585
R370 B.n412 B.n177 585
R371 B.n411 B.n410 585
R372 B.n413 B.n411 585
R373 B.n409 B.n182 585
R374 B.n182 B.n181 585
R375 B.n408 B.n407 585
R376 B.n407 B.n406 585
R377 B.n184 B.n183 585
R378 B.n185 B.n184 585
R379 B.n399 B.n398 585
R380 B.n400 B.n399 585
R381 B.n397 B.n190 585
R382 B.n190 B.n189 585
R383 B.n396 B.n395 585
R384 B.n395 B.n394 585
R385 B.n192 B.n191 585
R386 B.n193 B.n192 585
R387 B.n387 B.n386 585
R388 B.n388 B.n387 585
R389 B.n385 B.n197 585
R390 B.n201 B.n197 585
R391 B.n384 B.n383 585
R392 B.n383 B.n382 585
R393 B.n199 B.n198 585
R394 B.n200 B.n199 585
R395 B.n375 B.n374 585
R396 B.n376 B.n375 585
R397 B.n373 B.n206 585
R398 B.n206 B.n205 585
R399 B.n372 B.n371 585
R400 B.n371 B.n370 585
R401 B.n208 B.n207 585
R402 B.n209 B.n208 585
R403 B.n363 B.n362 585
R404 B.n364 B.n363 585
R405 B.n361 B.n214 585
R406 B.n214 B.n213 585
R407 B.n360 B.n359 585
R408 B.n359 B.n358 585
R409 B.n216 B.n215 585
R410 B.n217 B.n216 585
R411 B.n351 B.n350 585
R412 B.n352 B.n351 585
R413 B.n349 B.n222 585
R414 B.n222 B.n221 585
R415 B.n348 B.n347 585
R416 B.n347 B.n346 585
R417 B.n224 B.n223 585
R418 B.n225 B.n224 585
R419 B.n339 B.n338 585
R420 B.n340 B.n339 585
R421 B.n337 B.n230 585
R422 B.n230 B.n229 585
R423 B.n336 B.n335 585
R424 B.n335 B.n334 585
R425 B.n232 B.n231 585
R426 B.n233 B.n232 585
R427 B.n327 B.n326 585
R428 B.n328 B.n327 585
R429 B.n325 B.n238 585
R430 B.n238 B.n237 585
R431 B.n324 B.n323 585
R432 B.n323 B.n322 585
R433 B.n319 B.n242 585
R434 B.n318 B.n317 585
R435 B.n315 B.n243 585
R436 B.n315 B.n241 585
R437 B.n314 B.n313 585
R438 B.n312 B.n311 585
R439 B.n310 B.n245 585
R440 B.n308 B.n307 585
R441 B.n306 B.n246 585
R442 B.n305 B.n304 585
R443 B.n302 B.n247 585
R444 B.n300 B.n299 585
R445 B.n298 B.n248 585
R446 B.n297 B.n296 585
R447 B.n294 B.n252 585
R448 B.n292 B.n291 585
R449 B.n290 B.n253 585
R450 B.n289 B.n288 585
R451 B.n286 B.n254 585
R452 B.n284 B.n283 585
R453 B.n282 B.n255 585
R454 B.n280 B.n279 585
R455 B.n277 B.n258 585
R456 B.n275 B.n274 585
R457 B.n273 B.n259 585
R458 B.n272 B.n271 585
R459 B.n269 B.n260 585
R460 B.n267 B.n266 585
R461 B.n265 B.n261 585
R462 B.n264 B.n263 585
R463 B.n240 B.n239 585
R464 B.n241 B.n240 585
R465 B.n321 B.n320 585
R466 B.n322 B.n321 585
R467 B.n236 B.n235 585
R468 B.n237 B.n236 585
R469 B.n330 B.n329 585
R470 B.n329 B.n328 585
R471 B.n331 B.n234 585
R472 B.n234 B.n233 585
R473 B.n333 B.n332 585
R474 B.n334 B.n333 585
R475 B.n228 B.n227 585
R476 B.n229 B.n228 585
R477 B.n342 B.n341 585
R478 B.n341 B.n340 585
R479 B.n343 B.n226 585
R480 B.n226 B.n225 585
R481 B.n345 B.n344 585
R482 B.n346 B.n345 585
R483 B.n220 B.n219 585
R484 B.n221 B.n220 585
R485 B.n354 B.n353 585
R486 B.n353 B.n352 585
R487 B.n355 B.n218 585
R488 B.n218 B.n217 585
R489 B.n357 B.n356 585
R490 B.n358 B.n357 585
R491 B.n212 B.n211 585
R492 B.n213 B.n212 585
R493 B.n366 B.n365 585
R494 B.n365 B.n364 585
R495 B.n367 B.n210 585
R496 B.n210 B.n209 585
R497 B.n369 B.n368 585
R498 B.n370 B.n369 585
R499 B.n204 B.n203 585
R500 B.n205 B.n204 585
R501 B.n378 B.n377 585
R502 B.n377 B.n376 585
R503 B.n379 B.n202 585
R504 B.n202 B.n200 585
R505 B.n381 B.n380 585
R506 B.n382 B.n381 585
R507 B.n196 B.n195 585
R508 B.n201 B.n196 585
R509 B.n390 B.n389 585
R510 B.n389 B.n388 585
R511 B.n391 B.n194 585
R512 B.n194 B.n193 585
R513 B.n393 B.n392 585
R514 B.n394 B.n393 585
R515 B.n188 B.n187 585
R516 B.n189 B.n188 585
R517 B.n402 B.n401 585
R518 B.n401 B.n400 585
R519 B.n403 B.n186 585
R520 B.n186 B.n185 585
R521 B.n405 B.n404 585
R522 B.n406 B.n405 585
R523 B.n180 B.n179 585
R524 B.n181 B.n180 585
R525 B.n415 B.n414 585
R526 B.n414 B.n413 585
R527 B.n416 B.n178 585
R528 B.n412 B.n178 585
R529 B.n418 B.n417 585
R530 B.n419 B.n418 585
R531 B.n173 B.n172 585
R532 B.n174 B.n173 585
R533 B.n427 B.n426 585
R534 B.n426 B.n425 585
R535 B.n428 B.n171 585
R536 B.n171 B.n170 585
R537 B.n430 B.n429 585
R538 B.n431 B.n430 585
R539 B.n165 B.n164 585
R540 B.n166 B.n165 585
R541 B.n439 B.n438 585
R542 B.n438 B.n437 585
R543 B.n440 B.n163 585
R544 B.n163 B.n161 585
R545 B.n442 B.n441 585
R546 B.n443 B.n442 585
R547 B.n157 B.n156 585
R548 B.n162 B.n157 585
R549 B.n451 B.n450 585
R550 B.n450 B.n449 585
R551 B.n452 B.n155 585
R552 B.n155 B.n154 585
R553 B.n454 B.n453 585
R554 B.n455 B.n454 585
R555 B.n149 B.n148 585
R556 B.n150 B.n149 585
R557 B.n463 B.n462 585
R558 B.n462 B.n461 585
R559 B.n464 B.n147 585
R560 B.n147 B.n146 585
R561 B.n466 B.n465 585
R562 B.n467 B.n466 585
R563 B.n141 B.n140 585
R564 B.n142 B.n141 585
R565 B.n476 B.n475 585
R566 B.n475 B.n474 585
R567 B.n477 B.n139 585
R568 B.n473 B.n139 585
R569 B.n479 B.n478 585
R570 B.n480 B.n479 585
R571 B.n134 B.n133 585
R572 B.n135 B.n134 585
R573 B.n489 B.n488 585
R574 B.n488 B.n487 585
R575 B.n490 B.n132 585
R576 B.n132 B.n131 585
R577 B.n492 B.n491 585
R578 B.n493 B.n492 585
R579 B.n3 B.n0 585
R580 B.n4 B.n3 585
R581 B.n746 B.n1 585
R582 B.n747 B.n746 585
R583 B.n745 B.n744 585
R584 B.n745 B.n8 585
R585 B.n743 B.n9 585
R586 B.n12 B.n9 585
R587 B.n742 B.n741 585
R588 B.n741 B.n740 585
R589 B.n11 B.n10 585
R590 B.n739 B.n11 585
R591 B.n737 B.n736 585
R592 B.n738 B.n737 585
R593 B.n735 B.n16 585
R594 B.n19 B.n16 585
R595 B.n734 B.n733 585
R596 B.n733 B.n732 585
R597 B.n18 B.n17 585
R598 B.n731 B.n18 585
R599 B.n729 B.n728 585
R600 B.n730 B.n729 585
R601 B.n727 B.n24 585
R602 B.n24 B.n23 585
R603 B.n726 B.n725 585
R604 B.n725 B.n724 585
R605 B.n26 B.n25 585
R606 B.n723 B.n26 585
R607 B.n721 B.n720 585
R608 B.n722 B.n721 585
R609 B.n719 B.n31 585
R610 B.n31 B.n30 585
R611 B.n718 B.n717 585
R612 B.n717 B.n716 585
R613 B.n33 B.n32 585
R614 B.n715 B.n33 585
R615 B.n713 B.n712 585
R616 B.n714 B.n713 585
R617 B.n711 B.n38 585
R618 B.n38 B.n37 585
R619 B.n710 B.n709 585
R620 B.n709 B.n708 585
R621 B.n40 B.n39 585
R622 B.n707 B.n40 585
R623 B.n705 B.n704 585
R624 B.n706 B.n705 585
R625 B.n703 B.n45 585
R626 B.n45 B.n44 585
R627 B.n702 B.n701 585
R628 B.n701 B.n700 585
R629 B.n47 B.n46 585
R630 B.n699 B.n47 585
R631 B.n697 B.n696 585
R632 B.n698 B.n697 585
R633 B.n695 B.n51 585
R634 B.n54 B.n51 585
R635 B.n694 B.n693 585
R636 B.n693 B.n692 585
R637 B.n53 B.n52 585
R638 B.n691 B.n53 585
R639 B.n689 B.n688 585
R640 B.n690 B.n689 585
R641 B.n687 B.n59 585
R642 B.n59 B.n58 585
R643 B.n686 B.n685 585
R644 B.n685 B.n684 585
R645 B.n61 B.n60 585
R646 B.n683 B.n61 585
R647 B.n681 B.n680 585
R648 B.n682 B.n681 585
R649 B.n679 B.n66 585
R650 B.n66 B.n65 585
R651 B.n678 B.n677 585
R652 B.n677 B.n676 585
R653 B.n68 B.n67 585
R654 B.n675 B.n68 585
R655 B.n673 B.n672 585
R656 B.n674 B.n673 585
R657 B.n671 B.n73 585
R658 B.n73 B.n72 585
R659 B.n670 B.n669 585
R660 B.n669 B.n668 585
R661 B.n75 B.n74 585
R662 B.n667 B.n75 585
R663 B.n665 B.n664 585
R664 B.n666 B.n665 585
R665 B.n663 B.n80 585
R666 B.n80 B.n79 585
R667 B.n662 B.n661 585
R668 B.n661 B.n660 585
R669 B.n82 B.n81 585
R670 B.n659 B.n82 585
R671 B.n657 B.n656 585
R672 B.n658 B.n657 585
R673 B.n655 B.n87 585
R674 B.n87 B.n86 585
R675 B.n654 B.n653 585
R676 B.n653 B.n652 585
R677 B.n89 B.n88 585
R678 B.n651 B.n89 585
R679 B.n649 B.n648 585
R680 B.n650 B.n649 585
R681 B.n647 B.n94 585
R682 B.n94 B.n93 585
R683 B.n646 B.n645 585
R684 B.n645 B.n644 585
R685 B.n96 B.n95 585
R686 B.n643 B.n96 585
R687 B.n641 B.n640 585
R688 B.n642 B.n641 585
R689 B.n639 B.n101 585
R690 B.n101 B.n100 585
R691 B.n638 B.n637 585
R692 B.n637 B.n636 585
R693 B.n103 B.n102 585
R694 B.n635 B.n103 585
R695 B.n633 B.n632 585
R696 B.n634 B.n633 585
R697 B.n750 B.n749 585
R698 B.n748 B.n2 585
R699 B.n633 B.n108 506.916
R700 B.n573 B.n106 506.916
R701 B.n323 B.n240 506.916
R702 B.n321 B.n242 506.916
R703 B.n572 B.n107 256.663
R704 B.n578 B.n107 256.663
R705 B.n580 B.n107 256.663
R706 B.n586 B.n107 256.663
R707 B.n124 B.n107 256.663
R708 B.n592 B.n107 256.663
R709 B.n598 B.n107 256.663
R710 B.n600 B.n107 256.663
R711 B.n606 B.n107 256.663
R712 B.n116 B.n107 256.663
R713 B.n612 B.n107 256.663
R714 B.n618 B.n107 256.663
R715 B.n620 B.n107 256.663
R716 B.n626 B.n107 256.663
R717 B.n628 B.n107 256.663
R718 B.n316 B.n241 256.663
R719 B.n244 B.n241 256.663
R720 B.n309 B.n241 256.663
R721 B.n303 B.n241 256.663
R722 B.n301 B.n241 256.663
R723 B.n295 B.n241 256.663
R724 B.n293 B.n241 256.663
R725 B.n287 B.n241 256.663
R726 B.n285 B.n241 256.663
R727 B.n278 B.n241 256.663
R728 B.n276 B.n241 256.663
R729 B.n270 B.n241 256.663
R730 B.n268 B.n241 256.663
R731 B.n262 B.n241 256.663
R732 B.n752 B.n751 256.663
R733 B.n113 B.t20 217.088
R734 B.n249 B.t11 217.088
R735 B.n121 B.t14 217.088
R736 B.n256 B.t18 217.088
R737 B.n322 B.n241 211.827
R738 B.n634 B.n107 211.827
R739 B.n113 B.t19 209.304
R740 B.n121 B.t12 209.304
R741 B.n256 B.t16 209.304
R742 B.n249 B.t8 209.304
R743 B.n629 B.n627 163.367
R744 B.n625 B.n110 163.367
R745 B.n621 B.n619 163.367
R746 B.n617 B.n112 163.367
R747 B.n613 B.n611 163.367
R748 B.n608 B.n607 163.367
R749 B.n605 B.n118 163.367
R750 B.n601 B.n599 163.367
R751 B.n597 B.n120 163.367
R752 B.n593 B.n591 163.367
R753 B.n588 B.n587 163.367
R754 B.n585 B.n126 163.367
R755 B.n581 B.n579 163.367
R756 B.n577 B.n128 163.367
R757 B.n323 B.n238 163.367
R758 B.n327 B.n238 163.367
R759 B.n327 B.n232 163.367
R760 B.n335 B.n232 163.367
R761 B.n335 B.n230 163.367
R762 B.n339 B.n230 163.367
R763 B.n339 B.n224 163.367
R764 B.n347 B.n224 163.367
R765 B.n347 B.n222 163.367
R766 B.n351 B.n222 163.367
R767 B.n351 B.n216 163.367
R768 B.n359 B.n216 163.367
R769 B.n359 B.n214 163.367
R770 B.n363 B.n214 163.367
R771 B.n363 B.n208 163.367
R772 B.n371 B.n208 163.367
R773 B.n371 B.n206 163.367
R774 B.n375 B.n206 163.367
R775 B.n375 B.n199 163.367
R776 B.n383 B.n199 163.367
R777 B.n383 B.n197 163.367
R778 B.n387 B.n197 163.367
R779 B.n387 B.n192 163.367
R780 B.n395 B.n192 163.367
R781 B.n395 B.n190 163.367
R782 B.n399 B.n190 163.367
R783 B.n399 B.n184 163.367
R784 B.n407 B.n184 163.367
R785 B.n407 B.n182 163.367
R786 B.n411 B.n182 163.367
R787 B.n411 B.n177 163.367
R788 B.n420 B.n177 163.367
R789 B.n420 B.n175 163.367
R790 B.n424 B.n175 163.367
R791 B.n424 B.n169 163.367
R792 B.n432 B.n169 163.367
R793 B.n432 B.n167 163.367
R794 B.n436 B.n167 163.367
R795 B.n436 B.n160 163.367
R796 B.n444 B.n160 163.367
R797 B.n444 B.n158 163.367
R798 B.n448 B.n158 163.367
R799 B.n448 B.n153 163.367
R800 B.n456 B.n153 163.367
R801 B.n456 B.n151 163.367
R802 B.n460 B.n151 163.367
R803 B.n460 B.n145 163.367
R804 B.n468 B.n145 163.367
R805 B.n468 B.n143 163.367
R806 B.n472 B.n143 163.367
R807 B.n472 B.n138 163.367
R808 B.n481 B.n138 163.367
R809 B.n481 B.n136 163.367
R810 B.n486 B.n136 163.367
R811 B.n486 B.n130 163.367
R812 B.n494 B.n130 163.367
R813 B.n495 B.n494 163.367
R814 B.n495 B.n5 163.367
R815 B.n6 B.n5 163.367
R816 B.n7 B.n6 163.367
R817 B.n501 B.n7 163.367
R818 B.n502 B.n501 163.367
R819 B.n502 B.n13 163.367
R820 B.n14 B.n13 163.367
R821 B.n15 B.n14 163.367
R822 B.n507 B.n15 163.367
R823 B.n507 B.n20 163.367
R824 B.n21 B.n20 163.367
R825 B.n22 B.n21 163.367
R826 B.n512 B.n22 163.367
R827 B.n512 B.n27 163.367
R828 B.n28 B.n27 163.367
R829 B.n29 B.n28 163.367
R830 B.n517 B.n29 163.367
R831 B.n517 B.n34 163.367
R832 B.n35 B.n34 163.367
R833 B.n36 B.n35 163.367
R834 B.n522 B.n36 163.367
R835 B.n522 B.n41 163.367
R836 B.n42 B.n41 163.367
R837 B.n43 B.n42 163.367
R838 B.n527 B.n43 163.367
R839 B.n527 B.n48 163.367
R840 B.n49 B.n48 163.367
R841 B.n50 B.n49 163.367
R842 B.n532 B.n50 163.367
R843 B.n532 B.n55 163.367
R844 B.n56 B.n55 163.367
R845 B.n57 B.n56 163.367
R846 B.n537 B.n57 163.367
R847 B.n537 B.n62 163.367
R848 B.n63 B.n62 163.367
R849 B.n64 B.n63 163.367
R850 B.n542 B.n64 163.367
R851 B.n542 B.n69 163.367
R852 B.n70 B.n69 163.367
R853 B.n71 B.n70 163.367
R854 B.n547 B.n71 163.367
R855 B.n547 B.n76 163.367
R856 B.n77 B.n76 163.367
R857 B.n78 B.n77 163.367
R858 B.n552 B.n78 163.367
R859 B.n552 B.n83 163.367
R860 B.n84 B.n83 163.367
R861 B.n85 B.n84 163.367
R862 B.n557 B.n85 163.367
R863 B.n557 B.n90 163.367
R864 B.n91 B.n90 163.367
R865 B.n92 B.n91 163.367
R866 B.n562 B.n92 163.367
R867 B.n562 B.n97 163.367
R868 B.n98 B.n97 163.367
R869 B.n99 B.n98 163.367
R870 B.n567 B.n99 163.367
R871 B.n567 B.n104 163.367
R872 B.n105 B.n104 163.367
R873 B.n106 B.n105 163.367
R874 B.n317 B.n315 163.367
R875 B.n315 B.n314 163.367
R876 B.n311 B.n310 163.367
R877 B.n308 B.n246 163.367
R878 B.n304 B.n302 163.367
R879 B.n300 B.n248 163.367
R880 B.n296 B.n294 163.367
R881 B.n292 B.n253 163.367
R882 B.n288 B.n286 163.367
R883 B.n284 B.n255 163.367
R884 B.n279 B.n277 163.367
R885 B.n275 B.n259 163.367
R886 B.n271 B.n269 163.367
R887 B.n267 B.n261 163.367
R888 B.n263 B.n240 163.367
R889 B.n321 B.n236 163.367
R890 B.n329 B.n236 163.367
R891 B.n329 B.n234 163.367
R892 B.n333 B.n234 163.367
R893 B.n333 B.n228 163.367
R894 B.n341 B.n228 163.367
R895 B.n341 B.n226 163.367
R896 B.n345 B.n226 163.367
R897 B.n345 B.n220 163.367
R898 B.n353 B.n220 163.367
R899 B.n353 B.n218 163.367
R900 B.n357 B.n218 163.367
R901 B.n357 B.n212 163.367
R902 B.n365 B.n212 163.367
R903 B.n365 B.n210 163.367
R904 B.n369 B.n210 163.367
R905 B.n369 B.n204 163.367
R906 B.n377 B.n204 163.367
R907 B.n377 B.n202 163.367
R908 B.n381 B.n202 163.367
R909 B.n381 B.n196 163.367
R910 B.n389 B.n196 163.367
R911 B.n389 B.n194 163.367
R912 B.n393 B.n194 163.367
R913 B.n393 B.n188 163.367
R914 B.n401 B.n188 163.367
R915 B.n401 B.n186 163.367
R916 B.n405 B.n186 163.367
R917 B.n405 B.n180 163.367
R918 B.n414 B.n180 163.367
R919 B.n414 B.n178 163.367
R920 B.n418 B.n178 163.367
R921 B.n418 B.n173 163.367
R922 B.n426 B.n173 163.367
R923 B.n426 B.n171 163.367
R924 B.n430 B.n171 163.367
R925 B.n430 B.n165 163.367
R926 B.n438 B.n165 163.367
R927 B.n438 B.n163 163.367
R928 B.n442 B.n163 163.367
R929 B.n442 B.n157 163.367
R930 B.n450 B.n157 163.367
R931 B.n450 B.n155 163.367
R932 B.n454 B.n155 163.367
R933 B.n454 B.n149 163.367
R934 B.n462 B.n149 163.367
R935 B.n462 B.n147 163.367
R936 B.n466 B.n147 163.367
R937 B.n466 B.n141 163.367
R938 B.n475 B.n141 163.367
R939 B.n475 B.n139 163.367
R940 B.n479 B.n139 163.367
R941 B.n479 B.n134 163.367
R942 B.n488 B.n134 163.367
R943 B.n488 B.n132 163.367
R944 B.n492 B.n132 163.367
R945 B.n492 B.n3 163.367
R946 B.n750 B.n3 163.367
R947 B.n746 B.n2 163.367
R948 B.n746 B.n745 163.367
R949 B.n745 B.n9 163.367
R950 B.n741 B.n9 163.367
R951 B.n741 B.n11 163.367
R952 B.n737 B.n11 163.367
R953 B.n737 B.n16 163.367
R954 B.n733 B.n16 163.367
R955 B.n733 B.n18 163.367
R956 B.n729 B.n18 163.367
R957 B.n729 B.n24 163.367
R958 B.n725 B.n24 163.367
R959 B.n725 B.n26 163.367
R960 B.n721 B.n26 163.367
R961 B.n721 B.n31 163.367
R962 B.n717 B.n31 163.367
R963 B.n717 B.n33 163.367
R964 B.n713 B.n33 163.367
R965 B.n713 B.n38 163.367
R966 B.n709 B.n38 163.367
R967 B.n709 B.n40 163.367
R968 B.n705 B.n40 163.367
R969 B.n705 B.n45 163.367
R970 B.n701 B.n45 163.367
R971 B.n701 B.n47 163.367
R972 B.n697 B.n47 163.367
R973 B.n697 B.n51 163.367
R974 B.n693 B.n51 163.367
R975 B.n693 B.n53 163.367
R976 B.n689 B.n53 163.367
R977 B.n689 B.n59 163.367
R978 B.n685 B.n59 163.367
R979 B.n685 B.n61 163.367
R980 B.n681 B.n61 163.367
R981 B.n681 B.n66 163.367
R982 B.n677 B.n66 163.367
R983 B.n677 B.n68 163.367
R984 B.n673 B.n68 163.367
R985 B.n673 B.n73 163.367
R986 B.n669 B.n73 163.367
R987 B.n669 B.n75 163.367
R988 B.n665 B.n75 163.367
R989 B.n665 B.n80 163.367
R990 B.n661 B.n80 163.367
R991 B.n661 B.n82 163.367
R992 B.n657 B.n82 163.367
R993 B.n657 B.n87 163.367
R994 B.n653 B.n87 163.367
R995 B.n653 B.n89 163.367
R996 B.n649 B.n89 163.367
R997 B.n649 B.n94 163.367
R998 B.n645 B.n94 163.367
R999 B.n645 B.n96 163.367
R1000 B.n641 B.n96 163.367
R1001 B.n641 B.n101 163.367
R1002 B.n637 B.n101 163.367
R1003 B.n637 B.n103 163.367
R1004 B.n633 B.n103 163.367
R1005 B.n114 B.t21 150.566
R1006 B.n122 B.t15 150.566
R1007 B.n257 B.t17 150.566
R1008 B.n250 B.t10 150.566
R1009 B.n322 B.n237 113.419
R1010 B.n328 B.n237 113.419
R1011 B.n328 B.n233 113.419
R1012 B.n334 B.n233 113.419
R1013 B.n334 B.n229 113.419
R1014 B.n340 B.n229 113.419
R1015 B.n340 B.n225 113.419
R1016 B.n346 B.n225 113.419
R1017 B.n352 B.n221 113.419
R1018 B.n352 B.n217 113.419
R1019 B.n358 B.n217 113.419
R1020 B.n358 B.n213 113.419
R1021 B.n364 B.n213 113.419
R1022 B.n364 B.n209 113.419
R1023 B.n370 B.n209 113.419
R1024 B.n370 B.n205 113.419
R1025 B.n376 B.n205 113.419
R1026 B.n376 B.n200 113.419
R1027 B.n382 B.n200 113.419
R1028 B.n382 B.n201 113.419
R1029 B.n388 B.n193 113.419
R1030 B.n394 B.n193 113.419
R1031 B.n394 B.n189 113.419
R1032 B.n400 B.n189 113.419
R1033 B.n400 B.n185 113.419
R1034 B.n406 B.n185 113.419
R1035 B.n406 B.n181 113.419
R1036 B.n413 B.n181 113.419
R1037 B.n413 B.n412 113.419
R1038 B.n419 B.n174 113.419
R1039 B.n425 B.n174 113.419
R1040 B.n425 B.n170 113.419
R1041 B.n431 B.n170 113.419
R1042 B.n431 B.n166 113.419
R1043 B.n437 B.n166 113.419
R1044 B.n437 B.n161 113.419
R1045 B.n443 B.n161 113.419
R1046 B.n443 B.n162 113.419
R1047 B.n449 B.n154 113.419
R1048 B.n455 B.n154 113.419
R1049 B.n455 B.n150 113.419
R1050 B.n461 B.n150 113.419
R1051 B.n461 B.n146 113.419
R1052 B.n467 B.n146 113.419
R1053 B.n467 B.n142 113.419
R1054 B.n474 B.n142 113.419
R1055 B.n474 B.n473 113.419
R1056 B.n480 B.n135 113.419
R1057 B.n487 B.n135 113.419
R1058 B.n487 B.n131 113.419
R1059 B.n493 B.n131 113.419
R1060 B.n493 B.n4 113.419
R1061 B.n749 B.n4 113.419
R1062 B.n749 B.n748 113.419
R1063 B.n748 B.n747 113.419
R1064 B.n747 B.n8 113.419
R1065 B.n12 B.n8 113.419
R1066 B.n740 B.n12 113.419
R1067 B.n740 B.n739 113.419
R1068 B.n739 B.n738 113.419
R1069 B.n732 B.n19 113.419
R1070 B.n732 B.n731 113.419
R1071 B.n731 B.n730 113.419
R1072 B.n730 B.n23 113.419
R1073 B.n724 B.n23 113.419
R1074 B.n724 B.n723 113.419
R1075 B.n723 B.n722 113.419
R1076 B.n722 B.n30 113.419
R1077 B.n716 B.n30 113.419
R1078 B.n715 B.n714 113.419
R1079 B.n714 B.n37 113.419
R1080 B.n708 B.n37 113.419
R1081 B.n708 B.n707 113.419
R1082 B.n707 B.n706 113.419
R1083 B.n706 B.n44 113.419
R1084 B.n700 B.n44 113.419
R1085 B.n700 B.n699 113.419
R1086 B.n699 B.n698 113.419
R1087 B.n692 B.n54 113.419
R1088 B.n692 B.n691 113.419
R1089 B.n691 B.n690 113.419
R1090 B.n690 B.n58 113.419
R1091 B.n684 B.n58 113.419
R1092 B.n684 B.n683 113.419
R1093 B.n683 B.n682 113.419
R1094 B.n682 B.n65 113.419
R1095 B.n676 B.n65 113.419
R1096 B.n675 B.n674 113.419
R1097 B.n674 B.n72 113.419
R1098 B.n668 B.n72 113.419
R1099 B.n668 B.n667 113.419
R1100 B.n667 B.n666 113.419
R1101 B.n666 B.n79 113.419
R1102 B.n660 B.n79 113.419
R1103 B.n660 B.n659 113.419
R1104 B.n659 B.n658 113.419
R1105 B.n658 B.n86 113.419
R1106 B.n652 B.n86 113.419
R1107 B.n652 B.n651 113.419
R1108 B.n650 B.n93 113.419
R1109 B.n644 B.n93 113.419
R1110 B.n644 B.n643 113.419
R1111 B.n643 B.n642 113.419
R1112 B.n642 B.n100 113.419
R1113 B.n636 B.n100 113.419
R1114 B.n636 B.n635 113.419
R1115 B.n635 B.n634 113.419
R1116 B.n473 B.t4 96.7405
R1117 B.n19 B.t5 96.7405
R1118 B.n162 B.t6 86.7329
R1119 B.t7 B.n715 86.7329
R1120 B.t9 B.n221 80.0611
R1121 B.n651 B.t13 80.0611
R1122 B.n412 B.t3 76.7253
R1123 B.n54 B.t2 76.7253
R1124 B.n628 B.n108 71.676
R1125 B.n627 B.n626 71.676
R1126 B.n620 B.n110 71.676
R1127 B.n619 B.n618 71.676
R1128 B.n612 B.n112 71.676
R1129 B.n611 B.n116 71.676
R1130 B.n607 B.n606 71.676
R1131 B.n600 B.n118 71.676
R1132 B.n599 B.n598 71.676
R1133 B.n592 B.n120 71.676
R1134 B.n591 B.n124 71.676
R1135 B.n587 B.n586 71.676
R1136 B.n580 B.n126 71.676
R1137 B.n579 B.n578 71.676
R1138 B.n572 B.n128 71.676
R1139 B.n573 B.n572 71.676
R1140 B.n578 B.n577 71.676
R1141 B.n581 B.n580 71.676
R1142 B.n586 B.n585 71.676
R1143 B.n588 B.n124 71.676
R1144 B.n593 B.n592 71.676
R1145 B.n598 B.n597 71.676
R1146 B.n601 B.n600 71.676
R1147 B.n606 B.n605 71.676
R1148 B.n608 B.n116 71.676
R1149 B.n613 B.n612 71.676
R1150 B.n618 B.n617 71.676
R1151 B.n621 B.n620 71.676
R1152 B.n626 B.n625 71.676
R1153 B.n629 B.n628 71.676
R1154 B.n316 B.n242 71.676
R1155 B.n314 B.n244 71.676
R1156 B.n310 B.n309 71.676
R1157 B.n303 B.n246 71.676
R1158 B.n302 B.n301 71.676
R1159 B.n295 B.n248 71.676
R1160 B.n294 B.n293 71.676
R1161 B.n287 B.n253 71.676
R1162 B.n286 B.n285 71.676
R1163 B.n278 B.n255 71.676
R1164 B.n277 B.n276 71.676
R1165 B.n270 B.n259 71.676
R1166 B.n269 B.n268 71.676
R1167 B.n262 B.n261 71.676
R1168 B.n317 B.n316 71.676
R1169 B.n311 B.n244 71.676
R1170 B.n309 B.n308 71.676
R1171 B.n304 B.n303 71.676
R1172 B.n301 B.n300 71.676
R1173 B.n296 B.n295 71.676
R1174 B.n293 B.n292 71.676
R1175 B.n288 B.n287 71.676
R1176 B.n285 B.n284 71.676
R1177 B.n279 B.n278 71.676
R1178 B.n276 B.n275 71.676
R1179 B.n271 B.n270 71.676
R1180 B.n268 B.n267 71.676
R1181 B.n263 B.n262 71.676
R1182 B.n751 B.n750 71.676
R1183 B.n751 B.n2 71.676
R1184 B.n201 B.t1 66.7177
R1185 B.t0 B.n675 66.7177
R1186 B.n114 B.n113 66.5217
R1187 B.n122 B.n121 66.5217
R1188 B.n257 B.n256 66.5217
R1189 B.n250 B.n249 66.5217
R1190 B.n115 B.n114 59.5399
R1191 B.n123 B.n122 59.5399
R1192 B.n281 B.n257 59.5399
R1193 B.n251 B.n250 59.5399
R1194 B.n388 B.t1 46.7025
R1195 B.n676 B.t0 46.7025
R1196 B.n419 B.t3 36.695
R1197 B.n698 B.t2 36.695
R1198 B.n346 B.t9 33.3591
R1199 B.t13 B.n650 33.3591
R1200 B.n320 B.n319 32.9371
R1201 B.n324 B.n239 32.9371
R1202 B.n574 B.n571 32.9371
R1203 B.n632 B.n631 32.9371
R1204 B.n449 B.t6 26.6874
R1205 B.n716 B.t7 26.6874
R1206 B B.n752 18.0485
R1207 B.n480 B.t4 16.6798
R1208 B.n738 B.t5 16.6798
R1209 B.n320 B.n235 10.6151
R1210 B.n330 B.n235 10.6151
R1211 B.n331 B.n330 10.6151
R1212 B.n332 B.n331 10.6151
R1213 B.n332 B.n227 10.6151
R1214 B.n342 B.n227 10.6151
R1215 B.n343 B.n342 10.6151
R1216 B.n344 B.n343 10.6151
R1217 B.n344 B.n219 10.6151
R1218 B.n354 B.n219 10.6151
R1219 B.n355 B.n354 10.6151
R1220 B.n356 B.n355 10.6151
R1221 B.n356 B.n211 10.6151
R1222 B.n366 B.n211 10.6151
R1223 B.n367 B.n366 10.6151
R1224 B.n368 B.n367 10.6151
R1225 B.n368 B.n203 10.6151
R1226 B.n378 B.n203 10.6151
R1227 B.n379 B.n378 10.6151
R1228 B.n380 B.n379 10.6151
R1229 B.n380 B.n195 10.6151
R1230 B.n390 B.n195 10.6151
R1231 B.n391 B.n390 10.6151
R1232 B.n392 B.n391 10.6151
R1233 B.n392 B.n187 10.6151
R1234 B.n402 B.n187 10.6151
R1235 B.n403 B.n402 10.6151
R1236 B.n404 B.n403 10.6151
R1237 B.n404 B.n179 10.6151
R1238 B.n415 B.n179 10.6151
R1239 B.n416 B.n415 10.6151
R1240 B.n417 B.n416 10.6151
R1241 B.n417 B.n172 10.6151
R1242 B.n427 B.n172 10.6151
R1243 B.n428 B.n427 10.6151
R1244 B.n429 B.n428 10.6151
R1245 B.n429 B.n164 10.6151
R1246 B.n439 B.n164 10.6151
R1247 B.n440 B.n439 10.6151
R1248 B.n441 B.n440 10.6151
R1249 B.n441 B.n156 10.6151
R1250 B.n451 B.n156 10.6151
R1251 B.n452 B.n451 10.6151
R1252 B.n453 B.n452 10.6151
R1253 B.n453 B.n148 10.6151
R1254 B.n463 B.n148 10.6151
R1255 B.n464 B.n463 10.6151
R1256 B.n465 B.n464 10.6151
R1257 B.n465 B.n140 10.6151
R1258 B.n476 B.n140 10.6151
R1259 B.n477 B.n476 10.6151
R1260 B.n478 B.n477 10.6151
R1261 B.n478 B.n133 10.6151
R1262 B.n489 B.n133 10.6151
R1263 B.n490 B.n489 10.6151
R1264 B.n491 B.n490 10.6151
R1265 B.n491 B.n0 10.6151
R1266 B.n319 B.n318 10.6151
R1267 B.n318 B.n243 10.6151
R1268 B.n313 B.n243 10.6151
R1269 B.n313 B.n312 10.6151
R1270 B.n312 B.n245 10.6151
R1271 B.n307 B.n245 10.6151
R1272 B.n307 B.n306 10.6151
R1273 B.n306 B.n305 10.6151
R1274 B.n305 B.n247 10.6151
R1275 B.n299 B.n298 10.6151
R1276 B.n298 B.n297 10.6151
R1277 B.n297 B.n252 10.6151
R1278 B.n291 B.n252 10.6151
R1279 B.n291 B.n290 10.6151
R1280 B.n290 B.n289 10.6151
R1281 B.n289 B.n254 10.6151
R1282 B.n283 B.n254 10.6151
R1283 B.n283 B.n282 10.6151
R1284 B.n280 B.n258 10.6151
R1285 B.n274 B.n258 10.6151
R1286 B.n274 B.n273 10.6151
R1287 B.n273 B.n272 10.6151
R1288 B.n272 B.n260 10.6151
R1289 B.n266 B.n260 10.6151
R1290 B.n266 B.n265 10.6151
R1291 B.n265 B.n264 10.6151
R1292 B.n264 B.n239 10.6151
R1293 B.n325 B.n324 10.6151
R1294 B.n326 B.n325 10.6151
R1295 B.n326 B.n231 10.6151
R1296 B.n336 B.n231 10.6151
R1297 B.n337 B.n336 10.6151
R1298 B.n338 B.n337 10.6151
R1299 B.n338 B.n223 10.6151
R1300 B.n348 B.n223 10.6151
R1301 B.n349 B.n348 10.6151
R1302 B.n350 B.n349 10.6151
R1303 B.n350 B.n215 10.6151
R1304 B.n360 B.n215 10.6151
R1305 B.n361 B.n360 10.6151
R1306 B.n362 B.n361 10.6151
R1307 B.n362 B.n207 10.6151
R1308 B.n372 B.n207 10.6151
R1309 B.n373 B.n372 10.6151
R1310 B.n374 B.n373 10.6151
R1311 B.n374 B.n198 10.6151
R1312 B.n384 B.n198 10.6151
R1313 B.n385 B.n384 10.6151
R1314 B.n386 B.n385 10.6151
R1315 B.n386 B.n191 10.6151
R1316 B.n396 B.n191 10.6151
R1317 B.n397 B.n396 10.6151
R1318 B.n398 B.n397 10.6151
R1319 B.n398 B.n183 10.6151
R1320 B.n408 B.n183 10.6151
R1321 B.n409 B.n408 10.6151
R1322 B.n410 B.n409 10.6151
R1323 B.n410 B.n176 10.6151
R1324 B.n421 B.n176 10.6151
R1325 B.n422 B.n421 10.6151
R1326 B.n423 B.n422 10.6151
R1327 B.n423 B.n168 10.6151
R1328 B.n433 B.n168 10.6151
R1329 B.n434 B.n433 10.6151
R1330 B.n435 B.n434 10.6151
R1331 B.n435 B.n159 10.6151
R1332 B.n445 B.n159 10.6151
R1333 B.n446 B.n445 10.6151
R1334 B.n447 B.n446 10.6151
R1335 B.n447 B.n152 10.6151
R1336 B.n457 B.n152 10.6151
R1337 B.n458 B.n457 10.6151
R1338 B.n459 B.n458 10.6151
R1339 B.n459 B.n144 10.6151
R1340 B.n469 B.n144 10.6151
R1341 B.n470 B.n469 10.6151
R1342 B.n471 B.n470 10.6151
R1343 B.n471 B.n137 10.6151
R1344 B.n482 B.n137 10.6151
R1345 B.n483 B.n482 10.6151
R1346 B.n485 B.n483 10.6151
R1347 B.n485 B.n484 10.6151
R1348 B.n484 B.n129 10.6151
R1349 B.n496 B.n129 10.6151
R1350 B.n497 B.n496 10.6151
R1351 B.n498 B.n497 10.6151
R1352 B.n499 B.n498 10.6151
R1353 B.n500 B.n499 10.6151
R1354 B.n503 B.n500 10.6151
R1355 B.n504 B.n503 10.6151
R1356 B.n505 B.n504 10.6151
R1357 B.n506 B.n505 10.6151
R1358 B.n508 B.n506 10.6151
R1359 B.n509 B.n508 10.6151
R1360 B.n510 B.n509 10.6151
R1361 B.n511 B.n510 10.6151
R1362 B.n513 B.n511 10.6151
R1363 B.n514 B.n513 10.6151
R1364 B.n515 B.n514 10.6151
R1365 B.n516 B.n515 10.6151
R1366 B.n518 B.n516 10.6151
R1367 B.n519 B.n518 10.6151
R1368 B.n520 B.n519 10.6151
R1369 B.n521 B.n520 10.6151
R1370 B.n523 B.n521 10.6151
R1371 B.n524 B.n523 10.6151
R1372 B.n525 B.n524 10.6151
R1373 B.n526 B.n525 10.6151
R1374 B.n528 B.n526 10.6151
R1375 B.n529 B.n528 10.6151
R1376 B.n530 B.n529 10.6151
R1377 B.n531 B.n530 10.6151
R1378 B.n533 B.n531 10.6151
R1379 B.n534 B.n533 10.6151
R1380 B.n535 B.n534 10.6151
R1381 B.n536 B.n535 10.6151
R1382 B.n538 B.n536 10.6151
R1383 B.n539 B.n538 10.6151
R1384 B.n540 B.n539 10.6151
R1385 B.n541 B.n540 10.6151
R1386 B.n543 B.n541 10.6151
R1387 B.n544 B.n543 10.6151
R1388 B.n545 B.n544 10.6151
R1389 B.n546 B.n545 10.6151
R1390 B.n548 B.n546 10.6151
R1391 B.n549 B.n548 10.6151
R1392 B.n550 B.n549 10.6151
R1393 B.n551 B.n550 10.6151
R1394 B.n553 B.n551 10.6151
R1395 B.n554 B.n553 10.6151
R1396 B.n555 B.n554 10.6151
R1397 B.n556 B.n555 10.6151
R1398 B.n558 B.n556 10.6151
R1399 B.n559 B.n558 10.6151
R1400 B.n560 B.n559 10.6151
R1401 B.n561 B.n560 10.6151
R1402 B.n563 B.n561 10.6151
R1403 B.n564 B.n563 10.6151
R1404 B.n565 B.n564 10.6151
R1405 B.n566 B.n565 10.6151
R1406 B.n568 B.n566 10.6151
R1407 B.n569 B.n568 10.6151
R1408 B.n570 B.n569 10.6151
R1409 B.n571 B.n570 10.6151
R1410 B.n744 B.n1 10.6151
R1411 B.n744 B.n743 10.6151
R1412 B.n743 B.n742 10.6151
R1413 B.n742 B.n10 10.6151
R1414 B.n736 B.n10 10.6151
R1415 B.n736 B.n735 10.6151
R1416 B.n735 B.n734 10.6151
R1417 B.n734 B.n17 10.6151
R1418 B.n728 B.n17 10.6151
R1419 B.n728 B.n727 10.6151
R1420 B.n727 B.n726 10.6151
R1421 B.n726 B.n25 10.6151
R1422 B.n720 B.n25 10.6151
R1423 B.n720 B.n719 10.6151
R1424 B.n719 B.n718 10.6151
R1425 B.n718 B.n32 10.6151
R1426 B.n712 B.n32 10.6151
R1427 B.n712 B.n711 10.6151
R1428 B.n711 B.n710 10.6151
R1429 B.n710 B.n39 10.6151
R1430 B.n704 B.n39 10.6151
R1431 B.n704 B.n703 10.6151
R1432 B.n703 B.n702 10.6151
R1433 B.n702 B.n46 10.6151
R1434 B.n696 B.n46 10.6151
R1435 B.n696 B.n695 10.6151
R1436 B.n695 B.n694 10.6151
R1437 B.n694 B.n52 10.6151
R1438 B.n688 B.n52 10.6151
R1439 B.n688 B.n687 10.6151
R1440 B.n687 B.n686 10.6151
R1441 B.n686 B.n60 10.6151
R1442 B.n680 B.n60 10.6151
R1443 B.n680 B.n679 10.6151
R1444 B.n679 B.n678 10.6151
R1445 B.n678 B.n67 10.6151
R1446 B.n672 B.n67 10.6151
R1447 B.n672 B.n671 10.6151
R1448 B.n671 B.n670 10.6151
R1449 B.n670 B.n74 10.6151
R1450 B.n664 B.n74 10.6151
R1451 B.n664 B.n663 10.6151
R1452 B.n663 B.n662 10.6151
R1453 B.n662 B.n81 10.6151
R1454 B.n656 B.n81 10.6151
R1455 B.n656 B.n655 10.6151
R1456 B.n655 B.n654 10.6151
R1457 B.n654 B.n88 10.6151
R1458 B.n648 B.n88 10.6151
R1459 B.n648 B.n647 10.6151
R1460 B.n647 B.n646 10.6151
R1461 B.n646 B.n95 10.6151
R1462 B.n640 B.n95 10.6151
R1463 B.n640 B.n639 10.6151
R1464 B.n639 B.n638 10.6151
R1465 B.n638 B.n102 10.6151
R1466 B.n632 B.n102 10.6151
R1467 B.n631 B.n630 10.6151
R1468 B.n630 B.n109 10.6151
R1469 B.n624 B.n109 10.6151
R1470 B.n624 B.n623 10.6151
R1471 B.n623 B.n622 10.6151
R1472 B.n622 B.n111 10.6151
R1473 B.n616 B.n111 10.6151
R1474 B.n616 B.n615 10.6151
R1475 B.n615 B.n614 10.6151
R1476 B.n610 B.n609 10.6151
R1477 B.n609 B.n117 10.6151
R1478 B.n604 B.n117 10.6151
R1479 B.n604 B.n603 10.6151
R1480 B.n603 B.n602 10.6151
R1481 B.n602 B.n119 10.6151
R1482 B.n596 B.n119 10.6151
R1483 B.n596 B.n595 10.6151
R1484 B.n595 B.n594 10.6151
R1485 B.n590 B.n589 10.6151
R1486 B.n589 B.n125 10.6151
R1487 B.n584 B.n125 10.6151
R1488 B.n584 B.n583 10.6151
R1489 B.n583 B.n582 10.6151
R1490 B.n582 B.n127 10.6151
R1491 B.n576 B.n127 10.6151
R1492 B.n576 B.n575 10.6151
R1493 B.n575 B.n574 10.6151
R1494 B.n251 B.n247 9.36635
R1495 B.n281 B.n280 9.36635
R1496 B.n614 B.n115 9.36635
R1497 B.n590 B.n123 9.36635
R1498 B.n752 B.n0 8.11757
R1499 B.n752 B.n1 8.11757
R1500 B.n299 B.n251 1.24928
R1501 B.n282 B.n281 1.24928
R1502 B.n610 B.n115 1.24928
R1503 B.n594 B.n123 1.24928
R1504 VN.n60 VN.n59 161.3
R1505 VN.n58 VN.n32 161.3
R1506 VN.n57 VN.n56 161.3
R1507 VN.n55 VN.n33 161.3
R1508 VN.n54 VN.n53 161.3
R1509 VN.n52 VN.n34 161.3
R1510 VN.n51 VN.n50 161.3
R1511 VN.n49 VN.n48 161.3
R1512 VN.n47 VN.n36 161.3
R1513 VN.n46 VN.n45 161.3
R1514 VN.n44 VN.n37 161.3
R1515 VN.n43 VN.n42 161.3
R1516 VN.n41 VN.n38 161.3
R1517 VN.n29 VN.n28 161.3
R1518 VN.n27 VN.n1 161.3
R1519 VN.n26 VN.n25 161.3
R1520 VN.n24 VN.n2 161.3
R1521 VN.n23 VN.n22 161.3
R1522 VN.n21 VN.n3 161.3
R1523 VN.n20 VN.n19 161.3
R1524 VN.n18 VN.n17 161.3
R1525 VN.n16 VN.n5 161.3
R1526 VN.n15 VN.n14 161.3
R1527 VN.n13 VN.n6 161.3
R1528 VN.n12 VN.n11 161.3
R1529 VN.n10 VN.n7 161.3
R1530 VN.n30 VN.n0 70.818
R1531 VN.n61 VN.n31 70.818
R1532 VN.n15 VN.n6 56.5617
R1533 VN.n46 VN.n37 56.5617
R1534 VN.n26 VN.n2 56.5617
R1535 VN.n57 VN.n33 56.5617
R1536 VN.n9 VN.n8 51.1977
R1537 VN.n40 VN.n39 51.1977
R1538 VN VN.n61 45.4451
R1539 VN.n39 VN.t3 43.7245
R1540 VN.n8 VN.t1 43.7245
R1541 VN.n11 VN.n10 24.5923
R1542 VN.n11 VN.n6 24.5923
R1543 VN.n16 VN.n15 24.5923
R1544 VN.n17 VN.n16 24.5923
R1545 VN.n21 VN.n20 24.5923
R1546 VN.n22 VN.n21 24.5923
R1547 VN.n22 VN.n2 24.5923
R1548 VN.n27 VN.n26 24.5923
R1549 VN.n28 VN.n27 24.5923
R1550 VN.n42 VN.n37 24.5923
R1551 VN.n42 VN.n41 24.5923
R1552 VN.n53 VN.n33 24.5923
R1553 VN.n53 VN.n52 24.5923
R1554 VN.n52 VN.n51 24.5923
R1555 VN.n48 VN.n47 24.5923
R1556 VN.n47 VN.n46 24.5923
R1557 VN.n59 VN.n58 24.5923
R1558 VN.n58 VN.n57 24.5923
R1559 VN.n10 VN.n9 22.8709
R1560 VN.n17 VN.n4 22.8709
R1561 VN.n41 VN.n40 22.8709
R1562 VN.n48 VN.n35 22.8709
R1563 VN.n28 VN.n0 19.4281
R1564 VN.n59 VN.n31 19.4281
R1565 VN.n9 VN.t5 10.2624
R1566 VN.n4 VN.t2 10.2624
R1567 VN.n0 VN.t7 10.2624
R1568 VN.n40 VN.t0 10.2624
R1569 VN.n35 VN.t4 10.2624
R1570 VN.n31 VN.t6 10.2624
R1571 VN.n39 VN.n38 3.9322
R1572 VN.n8 VN.n7 3.9322
R1573 VN.n20 VN.n4 1.72193
R1574 VN.n51 VN.n35 1.72193
R1575 VN.n61 VN.n60 0.354861
R1576 VN.n30 VN.n29 0.354861
R1577 VN VN.n30 0.267071
R1578 VN.n60 VN.n32 0.189894
R1579 VN.n56 VN.n32 0.189894
R1580 VN.n56 VN.n55 0.189894
R1581 VN.n55 VN.n54 0.189894
R1582 VN.n54 VN.n34 0.189894
R1583 VN.n50 VN.n34 0.189894
R1584 VN.n50 VN.n49 0.189894
R1585 VN.n49 VN.n36 0.189894
R1586 VN.n45 VN.n36 0.189894
R1587 VN.n45 VN.n44 0.189894
R1588 VN.n44 VN.n43 0.189894
R1589 VN.n43 VN.n38 0.189894
R1590 VN.n12 VN.n7 0.189894
R1591 VN.n13 VN.n12 0.189894
R1592 VN.n14 VN.n13 0.189894
R1593 VN.n14 VN.n5 0.189894
R1594 VN.n18 VN.n5 0.189894
R1595 VN.n19 VN.n18 0.189894
R1596 VN.n19 VN.n3 0.189894
R1597 VN.n23 VN.n3 0.189894
R1598 VN.n24 VN.n23 0.189894
R1599 VN.n25 VN.n24 0.189894
R1600 VN.n25 VN.n1 0.189894
R1601 VN.n29 VN.n1 0.189894
R1602 VDD2.n2 VDD2.n1 148.627
R1603 VDD2.n2 VDD2.n0 148.627
R1604 VDD2 VDD2.n5 148.625
R1605 VDD2.n4 VDD2.n3 147.203
R1606 VDD2.n4 VDD2.n2 38.1593
R1607 VDD2.n5 VDD2.t7 15.0005
R1608 VDD2.n5 VDD2.t4 15.0005
R1609 VDD2.n3 VDD2.t1 15.0005
R1610 VDD2.n3 VDD2.t3 15.0005
R1611 VDD2.n1 VDD2.t5 15.0005
R1612 VDD2.n1 VDD2.t0 15.0005
R1613 VDD2.n0 VDD2.t6 15.0005
R1614 VDD2.n0 VDD2.t2 15.0005
R1615 VDD2 VDD2.n4 1.53714
C0 VP VDD2 0.581773f
C1 VN VDD1 0.159736f
C2 VTAIL VN 2.85749f
C3 VN VP 6.29938f
C4 VN VDD2 1.40396f
C5 VTAIL VDD1 4.95777f
C6 VP VDD1 1.82208f
C7 VDD1 VDD2 2.03873f
C8 VTAIL VP 2.8716f
C9 VTAIL VDD2 5.01554f
C10 VDD2 B 5.030758f
C11 VDD1 B 5.500801f
C12 VTAIL B 3.856455f
C13 VN B 16.51349f
C14 VP B 15.036797f
C15 VDD2.t6 B 0.02736f
C16 VDD2.t2 B 0.02736f
C17 VDD2.n0 B 0.142633f
C18 VDD2.t5 B 0.02736f
C19 VDD2.t0 B 0.02736f
C20 VDD2.n1 B 0.142633f
C21 VDD2.n2 B 3.02052f
C22 VDD2.t1 B 0.02736f
C23 VDD2.t3 B 0.02736f
C24 VDD2.n3 B 0.137165f
C25 VDD2.n4 B 2.3807f
C26 VDD2.t7 B 0.02736f
C27 VDD2.t4 B 0.02736f
C28 VDD2.n5 B 0.142616f
C29 VN.t7 B 0.233176f
C30 VN.n0 B 0.237554f
C31 VN.n1 B 0.027203f
C32 VN.n2 B 0.034275f
C33 VN.n3 B 0.027203f
C34 VN.t2 B 0.233176f
C35 VN.n4 B 0.128887f
C36 VN.n5 B 0.027203f
C37 VN.n6 B 0.039543f
C38 VN.n7 B 0.310476f
C39 VN.t5 B 0.233176f
C40 VN.t1 B 0.478398f
C41 VN.n8 B 0.233782f
C42 VN.n9 B 0.228071f
C43 VN.n10 B 0.048702f
C44 VN.n11 B 0.050445f
C45 VN.n12 B 0.027203f
C46 VN.n13 B 0.027203f
C47 VN.n14 B 0.027203f
C48 VN.n15 B 0.039543f
C49 VN.n16 B 0.050445f
C50 VN.n17 B 0.048702f
C51 VN.n18 B 0.027203f
C52 VN.n19 B 0.027203f
C53 VN.n20 B 0.027285f
C54 VN.n21 B 0.050445f
C55 VN.n22 B 0.050445f
C56 VN.n23 B 0.027203f
C57 VN.n24 B 0.027203f
C58 VN.n25 B 0.027203f
C59 VN.n26 B 0.044812f
C60 VN.n27 B 0.050445f
C61 VN.n28 B 0.045215f
C62 VN.n29 B 0.043898f
C63 VN.n30 B 0.058308f
C64 VN.t6 B 0.233176f
C65 VN.n31 B 0.237554f
C66 VN.n32 B 0.027203f
C67 VN.n33 B 0.034275f
C68 VN.n34 B 0.027203f
C69 VN.t4 B 0.233176f
C70 VN.n35 B 0.128887f
C71 VN.n36 B 0.027203f
C72 VN.n37 B 0.039543f
C73 VN.n38 B 0.310476f
C74 VN.t0 B 0.233176f
C75 VN.t3 B 0.478398f
C76 VN.n39 B 0.233782f
C77 VN.n40 B 0.228071f
C78 VN.n41 B 0.048702f
C79 VN.n42 B 0.050445f
C80 VN.n43 B 0.027203f
C81 VN.n44 B 0.027203f
C82 VN.n45 B 0.027203f
C83 VN.n46 B 0.039543f
C84 VN.n47 B 0.050445f
C85 VN.n48 B 0.048702f
C86 VN.n49 B 0.027203f
C87 VN.n50 B 0.027203f
C88 VN.n51 B 0.027285f
C89 VN.n52 B 0.050445f
C90 VN.n53 B 0.050445f
C91 VN.n54 B 0.027203f
C92 VN.n55 B 0.027203f
C93 VN.n56 B 0.027203f
C94 VN.n57 B 0.044812f
C95 VN.n58 B 0.050445f
C96 VN.n59 B 0.045215f
C97 VN.n60 B 0.043898f
C98 VN.n61 B 1.34145f
C99 VTAIL.t7 B 0.038324f
C100 VTAIL.t2 B 0.038324f
C101 VTAIL.n0 B 0.159038f
C102 VTAIL.n1 B 0.606115f
C103 VTAIL.t5 B 0.223464f
C104 VTAIL.n2 B 0.694941f
C105 VTAIL.t13 B 0.223464f
C106 VTAIL.n3 B 0.694941f
C107 VTAIL.t14 B 0.038324f
C108 VTAIL.t10 B 0.038324f
C109 VTAIL.n4 B 0.159038f
C110 VTAIL.n5 B 0.949281f
C111 VTAIL.t15 B 0.223464f
C112 VTAIL.n6 B 1.62316f
C113 VTAIL.t1 B 0.223464f
C114 VTAIL.n7 B 1.62316f
C115 VTAIL.t3 B 0.038324f
C116 VTAIL.t6 B 0.038324f
C117 VTAIL.n8 B 0.159037f
C118 VTAIL.n9 B 0.949281f
C119 VTAIL.t4 B 0.223464f
C120 VTAIL.n10 B 0.694941f
C121 VTAIL.t12 B 0.223464f
C122 VTAIL.n11 B 0.694941f
C123 VTAIL.t9 B 0.038324f
C124 VTAIL.t8 B 0.038324f
C125 VTAIL.n12 B 0.159037f
C126 VTAIL.n13 B 0.949281f
C127 VTAIL.t11 B 0.223464f
C128 VTAIL.n14 B 1.62316f
C129 VTAIL.t0 B 0.223464f
C130 VTAIL.n15 B 1.61628f
C131 VDD1.t2 B 0.026986f
C132 VDD1.t6 B 0.026986f
C133 VDD1.n0 B 0.141205f
C134 VDD1.t3 B 0.026986f
C135 VDD1.t1 B 0.026986f
C136 VDD1.n1 B 0.140686f
C137 VDD1.t7 B 0.026986f
C138 VDD1.t0 B 0.026986f
C139 VDD1.n2 B 0.140686f
C140 VDD1.n3 B 3.0331f
C141 VDD1.t4 B 0.026986f
C142 VDD1.t5 B 0.026986f
C143 VDD1.n4 B 0.135293f
C144 VDD1.n5 B 2.38024f
C145 VP.t2 B 0.234149f
C146 VP.n0 B 0.238545f
C147 VP.n1 B 0.027316f
C148 VP.n2 B 0.034418f
C149 VP.n3 B 0.027316f
C150 VP.t5 B 0.234149f
C151 VP.n4 B 0.129425f
C152 VP.n5 B 0.027316f
C153 VP.n6 B 0.039708f
C154 VP.n7 B 0.027316f
C155 VP.t1 B 0.234149f
C156 VP.n8 B 0.050655f
C157 VP.n9 B 0.027316f
C158 VP.n10 B 0.050655f
C159 VP.t4 B 0.234149f
C160 VP.n11 B 0.238545f
C161 VP.n12 B 0.027316f
C162 VP.n13 B 0.034418f
C163 VP.n14 B 0.027316f
C164 VP.t7 B 0.234149f
C165 VP.n15 B 0.129425f
C166 VP.n16 B 0.027316f
C167 VP.n17 B 0.039708f
C168 VP.n18 B 0.311773f
C169 VP.t6 B 0.234149f
C170 VP.t3 B 0.480394f
C171 VP.n19 B 0.234758f
C172 VP.n20 B 0.229023f
C173 VP.n21 B 0.048905f
C174 VP.n22 B 0.050655f
C175 VP.n23 B 0.027316f
C176 VP.n24 B 0.027316f
C177 VP.n25 B 0.027316f
C178 VP.n26 B 0.039708f
C179 VP.n27 B 0.050655f
C180 VP.n28 B 0.048905f
C181 VP.n29 B 0.027316f
C182 VP.n30 B 0.027316f
C183 VP.n31 B 0.027399f
C184 VP.n32 B 0.050655f
C185 VP.n33 B 0.050655f
C186 VP.n34 B 0.027316f
C187 VP.n35 B 0.027316f
C188 VP.n36 B 0.027316f
C189 VP.n37 B 0.044999f
C190 VP.n38 B 0.050655f
C191 VP.n39 B 0.045404f
C192 VP.n40 B 0.044081f
C193 VP.n41 B 1.33548f
C194 VP.n42 B 1.35723f
C195 VP.t0 B 0.234149f
C196 VP.n43 B 0.238545f
C197 VP.n44 B 0.045404f
C198 VP.n45 B 0.044081f
C199 VP.n46 B 0.027316f
C200 VP.n47 B 0.027316f
C201 VP.n48 B 0.044999f
C202 VP.n49 B 0.034418f
C203 VP.n50 B 0.050655f
C204 VP.n51 B 0.027316f
C205 VP.n52 B 0.027316f
C206 VP.n53 B 0.027316f
C207 VP.n54 B 0.027399f
C208 VP.n55 B 0.129425f
C209 VP.n56 B 0.048905f
C210 VP.n57 B 0.050655f
C211 VP.n58 B 0.027316f
C212 VP.n59 B 0.027316f
C213 VP.n60 B 0.027316f
C214 VP.n61 B 0.039708f
C215 VP.n62 B 0.050655f
C216 VP.n63 B 0.048905f
C217 VP.n64 B 0.027316f
C218 VP.n65 B 0.027316f
C219 VP.n66 B 0.027399f
C220 VP.n67 B 0.050655f
C221 VP.n68 B 0.050655f
C222 VP.n69 B 0.027316f
C223 VP.n70 B 0.027316f
C224 VP.n71 B 0.027316f
C225 VP.n72 B 0.044999f
C226 VP.n73 B 0.050655f
C227 VP.n74 B 0.045404f
C228 VP.n75 B 0.044081f
C229 VP.n76 B 0.058551f
.ends

