* NGSPICE file created from diff_pair_sample_1186.ext - technology: sky130A

.subckt diff_pair_sample_1186 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t6 VN.t0 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=2.8665 pd=15.48 as=1.21275 ps=7.68 w=7.35 l=3.05
X1 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=2.8665 pd=15.48 as=0 ps=0 w=7.35 l=3.05
X2 VDD1.t3 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.21275 pd=7.68 as=2.8665 ps=15.48 w=7.35 l=3.05
X3 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=2.8665 pd=15.48 as=0 ps=0 w=7.35 l=3.05
X4 VDD2.t1 VN.t1 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.21275 pd=7.68 as=2.8665 ps=15.48 w=7.35 l=3.05
X5 VTAIL.t4 VN.t2 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=2.8665 pd=15.48 as=1.21275 ps=7.68 w=7.35 l=3.05
X6 VTAIL.t7 VP.t1 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.8665 pd=15.48 as=1.21275 ps=7.68 w=7.35 l=3.05
X7 VDD1.t1 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.21275 pd=7.68 as=2.8665 ps=15.48 w=7.35 l=3.05
X8 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.8665 pd=15.48 as=0 ps=0 w=7.35 l=3.05
X9 VDD2.t2 VN.t3 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.21275 pd=7.68 as=2.8665 ps=15.48 w=7.35 l=3.05
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.8665 pd=15.48 as=0 ps=0 w=7.35 l=3.05
X11 VTAIL.t0 VP.t3 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.8665 pd=15.48 as=1.21275 ps=7.68 w=7.35 l=3.05
R0 VN.n1 VN.t3 92.5657
R1 VN.n0 VN.t0 92.5657
R2 VN.n0 VN.t1 91.5625
R3 VN.n1 VN.t2 91.5625
R4 VN VN.n1 47.3317
R5 VN VN.n0 2.91879
R6 VDD2.n2 VDD2.n0 102.248
R7 VDD2.n2 VDD2.n1 63.4549
R8 VDD2.n1 VDD2.t3 2.69438
R9 VDD2.n1 VDD2.t2 2.69438
R10 VDD2.n0 VDD2.t0 2.69438
R11 VDD2.n0 VDD2.t1 2.69438
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n314 VTAIL.n280 289.615
R14 VTAIL.n34 VTAIL.n0 289.615
R15 VTAIL.n74 VTAIL.n40 289.615
R16 VTAIL.n114 VTAIL.n80 289.615
R17 VTAIL.n274 VTAIL.n240 289.615
R18 VTAIL.n234 VTAIL.n200 289.615
R19 VTAIL.n194 VTAIL.n160 289.615
R20 VTAIL.n154 VTAIL.n120 289.615
R21 VTAIL.n292 VTAIL.n291 185
R22 VTAIL.n297 VTAIL.n296 185
R23 VTAIL.n299 VTAIL.n298 185
R24 VTAIL.n288 VTAIL.n287 185
R25 VTAIL.n305 VTAIL.n304 185
R26 VTAIL.n307 VTAIL.n306 185
R27 VTAIL.n284 VTAIL.n283 185
R28 VTAIL.n313 VTAIL.n312 185
R29 VTAIL.n315 VTAIL.n314 185
R30 VTAIL.n12 VTAIL.n11 185
R31 VTAIL.n17 VTAIL.n16 185
R32 VTAIL.n19 VTAIL.n18 185
R33 VTAIL.n8 VTAIL.n7 185
R34 VTAIL.n25 VTAIL.n24 185
R35 VTAIL.n27 VTAIL.n26 185
R36 VTAIL.n4 VTAIL.n3 185
R37 VTAIL.n33 VTAIL.n32 185
R38 VTAIL.n35 VTAIL.n34 185
R39 VTAIL.n52 VTAIL.n51 185
R40 VTAIL.n57 VTAIL.n56 185
R41 VTAIL.n59 VTAIL.n58 185
R42 VTAIL.n48 VTAIL.n47 185
R43 VTAIL.n65 VTAIL.n64 185
R44 VTAIL.n67 VTAIL.n66 185
R45 VTAIL.n44 VTAIL.n43 185
R46 VTAIL.n73 VTAIL.n72 185
R47 VTAIL.n75 VTAIL.n74 185
R48 VTAIL.n92 VTAIL.n91 185
R49 VTAIL.n97 VTAIL.n96 185
R50 VTAIL.n99 VTAIL.n98 185
R51 VTAIL.n88 VTAIL.n87 185
R52 VTAIL.n105 VTAIL.n104 185
R53 VTAIL.n107 VTAIL.n106 185
R54 VTAIL.n84 VTAIL.n83 185
R55 VTAIL.n113 VTAIL.n112 185
R56 VTAIL.n115 VTAIL.n114 185
R57 VTAIL.n275 VTAIL.n274 185
R58 VTAIL.n273 VTAIL.n272 185
R59 VTAIL.n244 VTAIL.n243 185
R60 VTAIL.n267 VTAIL.n266 185
R61 VTAIL.n265 VTAIL.n264 185
R62 VTAIL.n248 VTAIL.n247 185
R63 VTAIL.n259 VTAIL.n258 185
R64 VTAIL.n257 VTAIL.n256 185
R65 VTAIL.n252 VTAIL.n251 185
R66 VTAIL.n235 VTAIL.n234 185
R67 VTAIL.n233 VTAIL.n232 185
R68 VTAIL.n204 VTAIL.n203 185
R69 VTAIL.n227 VTAIL.n226 185
R70 VTAIL.n225 VTAIL.n224 185
R71 VTAIL.n208 VTAIL.n207 185
R72 VTAIL.n219 VTAIL.n218 185
R73 VTAIL.n217 VTAIL.n216 185
R74 VTAIL.n212 VTAIL.n211 185
R75 VTAIL.n195 VTAIL.n194 185
R76 VTAIL.n193 VTAIL.n192 185
R77 VTAIL.n164 VTAIL.n163 185
R78 VTAIL.n187 VTAIL.n186 185
R79 VTAIL.n185 VTAIL.n184 185
R80 VTAIL.n168 VTAIL.n167 185
R81 VTAIL.n179 VTAIL.n178 185
R82 VTAIL.n177 VTAIL.n176 185
R83 VTAIL.n172 VTAIL.n171 185
R84 VTAIL.n155 VTAIL.n154 185
R85 VTAIL.n153 VTAIL.n152 185
R86 VTAIL.n124 VTAIL.n123 185
R87 VTAIL.n147 VTAIL.n146 185
R88 VTAIL.n145 VTAIL.n144 185
R89 VTAIL.n128 VTAIL.n127 185
R90 VTAIL.n139 VTAIL.n138 185
R91 VTAIL.n137 VTAIL.n136 185
R92 VTAIL.n132 VTAIL.n131 185
R93 VTAIL.n293 VTAIL.t5 147.659
R94 VTAIL.n13 VTAIL.t6 147.659
R95 VTAIL.n53 VTAIL.t1 147.659
R96 VTAIL.n93 VTAIL.t0 147.659
R97 VTAIL.n253 VTAIL.t2 147.659
R98 VTAIL.n213 VTAIL.t7 147.659
R99 VTAIL.n173 VTAIL.t3 147.659
R100 VTAIL.n133 VTAIL.t4 147.659
R101 VTAIL.n297 VTAIL.n291 104.615
R102 VTAIL.n298 VTAIL.n297 104.615
R103 VTAIL.n298 VTAIL.n287 104.615
R104 VTAIL.n305 VTAIL.n287 104.615
R105 VTAIL.n306 VTAIL.n305 104.615
R106 VTAIL.n306 VTAIL.n283 104.615
R107 VTAIL.n313 VTAIL.n283 104.615
R108 VTAIL.n314 VTAIL.n313 104.615
R109 VTAIL.n17 VTAIL.n11 104.615
R110 VTAIL.n18 VTAIL.n17 104.615
R111 VTAIL.n18 VTAIL.n7 104.615
R112 VTAIL.n25 VTAIL.n7 104.615
R113 VTAIL.n26 VTAIL.n25 104.615
R114 VTAIL.n26 VTAIL.n3 104.615
R115 VTAIL.n33 VTAIL.n3 104.615
R116 VTAIL.n34 VTAIL.n33 104.615
R117 VTAIL.n57 VTAIL.n51 104.615
R118 VTAIL.n58 VTAIL.n57 104.615
R119 VTAIL.n58 VTAIL.n47 104.615
R120 VTAIL.n65 VTAIL.n47 104.615
R121 VTAIL.n66 VTAIL.n65 104.615
R122 VTAIL.n66 VTAIL.n43 104.615
R123 VTAIL.n73 VTAIL.n43 104.615
R124 VTAIL.n74 VTAIL.n73 104.615
R125 VTAIL.n97 VTAIL.n91 104.615
R126 VTAIL.n98 VTAIL.n97 104.615
R127 VTAIL.n98 VTAIL.n87 104.615
R128 VTAIL.n105 VTAIL.n87 104.615
R129 VTAIL.n106 VTAIL.n105 104.615
R130 VTAIL.n106 VTAIL.n83 104.615
R131 VTAIL.n113 VTAIL.n83 104.615
R132 VTAIL.n114 VTAIL.n113 104.615
R133 VTAIL.n274 VTAIL.n273 104.615
R134 VTAIL.n273 VTAIL.n243 104.615
R135 VTAIL.n266 VTAIL.n243 104.615
R136 VTAIL.n266 VTAIL.n265 104.615
R137 VTAIL.n265 VTAIL.n247 104.615
R138 VTAIL.n258 VTAIL.n247 104.615
R139 VTAIL.n258 VTAIL.n257 104.615
R140 VTAIL.n257 VTAIL.n251 104.615
R141 VTAIL.n234 VTAIL.n233 104.615
R142 VTAIL.n233 VTAIL.n203 104.615
R143 VTAIL.n226 VTAIL.n203 104.615
R144 VTAIL.n226 VTAIL.n225 104.615
R145 VTAIL.n225 VTAIL.n207 104.615
R146 VTAIL.n218 VTAIL.n207 104.615
R147 VTAIL.n218 VTAIL.n217 104.615
R148 VTAIL.n217 VTAIL.n211 104.615
R149 VTAIL.n194 VTAIL.n193 104.615
R150 VTAIL.n193 VTAIL.n163 104.615
R151 VTAIL.n186 VTAIL.n163 104.615
R152 VTAIL.n186 VTAIL.n185 104.615
R153 VTAIL.n185 VTAIL.n167 104.615
R154 VTAIL.n178 VTAIL.n167 104.615
R155 VTAIL.n178 VTAIL.n177 104.615
R156 VTAIL.n177 VTAIL.n171 104.615
R157 VTAIL.n154 VTAIL.n153 104.615
R158 VTAIL.n153 VTAIL.n123 104.615
R159 VTAIL.n146 VTAIL.n123 104.615
R160 VTAIL.n146 VTAIL.n145 104.615
R161 VTAIL.n145 VTAIL.n127 104.615
R162 VTAIL.n138 VTAIL.n127 104.615
R163 VTAIL.n138 VTAIL.n137 104.615
R164 VTAIL.n137 VTAIL.n131 104.615
R165 VTAIL.t5 VTAIL.n291 52.3082
R166 VTAIL.t6 VTAIL.n11 52.3082
R167 VTAIL.t1 VTAIL.n51 52.3082
R168 VTAIL.t0 VTAIL.n91 52.3082
R169 VTAIL.t2 VTAIL.n251 52.3082
R170 VTAIL.t7 VTAIL.n211 52.3082
R171 VTAIL.t3 VTAIL.n171 52.3082
R172 VTAIL.t4 VTAIL.n131 52.3082
R173 VTAIL.n319 VTAIL.n318 30.4399
R174 VTAIL.n39 VTAIL.n38 30.4399
R175 VTAIL.n79 VTAIL.n78 30.4399
R176 VTAIL.n119 VTAIL.n118 30.4399
R177 VTAIL.n279 VTAIL.n278 30.4399
R178 VTAIL.n239 VTAIL.n238 30.4399
R179 VTAIL.n199 VTAIL.n198 30.4399
R180 VTAIL.n159 VTAIL.n158 30.4399
R181 VTAIL.n319 VTAIL.n279 21.6169
R182 VTAIL.n159 VTAIL.n119 21.6169
R183 VTAIL.n293 VTAIL.n292 15.6677
R184 VTAIL.n13 VTAIL.n12 15.6677
R185 VTAIL.n53 VTAIL.n52 15.6677
R186 VTAIL.n93 VTAIL.n92 15.6677
R187 VTAIL.n253 VTAIL.n252 15.6677
R188 VTAIL.n213 VTAIL.n212 15.6677
R189 VTAIL.n173 VTAIL.n172 15.6677
R190 VTAIL.n133 VTAIL.n132 15.6677
R191 VTAIL.n296 VTAIL.n295 12.8005
R192 VTAIL.n16 VTAIL.n15 12.8005
R193 VTAIL.n56 VTAIL.n55 12.8005
R194 VTAIL.n96 VTAIL.n95 12.8005
R195 VTAIL.n256 VTAIL.n255 12.8005
R196 VTAIL.n216 VTAIL.n215 12.8005
R197 VTAIL.n176 VTAIL.n175 12.8005
R198 VTAIL.n136 VTAIL.n135 12.8005
R199 VTAIL.n299 VTAIL.n290 12.0247
R200 VTAIL.n19 VTAIL.n10 12.0247
R201 VTAIL.n59 VTAIL.n50 12.0247
R202 VTAIL.n99 VTAIL.n90 12.0247
R203 VTAIL.n259 VTAIL.n250 12.0247
R204 VTAIL.n219 VTAIL.n210 12.0247
R205 VTAIL.n179 VTAIL.n170 12.0247
R206 VTAIL.n139 VTAIL.n130 12.0247
R207 VTAIL.n300 VTAIL.n288 11.249
R208 VTAIL.n20 VTAIL.n8 11.249
R209 VTAIL.n60 VTAIL.n48 11.249
R210 VTAIL.n100 VTAIL.n88 11.249
R211 VTAIL.n260 VTAIL.n248 11.249
R212 VTAIL.n220 VTAIL.n208 11.249
R213 VTAIL.n180 VTAIL.n168 11.249
R214 VTAIL.n140 VTAIL.n128 11.249
R215 VTAIL.n304 VTAIL.n303 10.4732
R216 VTAIL.n24 VTAIL.n23 10.4732
R217 VTAIL.n64 VTAIL.n63 10.4732
R218 VTAIL.n104 VTAIL.n103 10.4732
R219 VTAIL.n264 VTAIL.n263 10.4732
R220 VTAIL.n224 VTAIL.n223 10.4732
R221 VTAIL.n184 VTAIL.n183 10.4732
R222 VTAIL.n144 VTAIL.n143 10.4732
R223 VTAIL.n307 VTAIL.n286 9.69747
R224 VTAIL.n27 VTAIL.n6 9.69747
R225 VTAIL.n67 VTAIL.n46 9.69747
R226 VTAIL.n107 VTAIL.n86 9.69747
R227 VTAIL.n267 VTAIL.n246 9.69747
R228 VTAIL.n227 VTAIL.n206 9.69747
R229 VTAIL.n187 VTAIL.n166 9.69747
R230 VTAIL.n147 VTAIL.n126 9.69747
R231 VTAIL.n318 VTAIL.n317 9.45567
R232 VTAIL.n38 VTAIL.n37 9.45567
R233 VTAIL.n78 VTAIL.n77 9.45567
R234 VTAIL.n118 VTAIL.n117 9.45567
R235 VTAIL.n278 VTAIL.n277 9.45567
R236 VTAIL.n238 VTAIL.n237 9.45567
R237 VTAIL.n198 VTAIL.n197 9.45567
R238 VTAIL.n158 VTAIL.n157 9.45567
R239 VTAIL.n317 VTAIL.n316 9.3005
R240 VTAIL.n311 VTAIL.n310 9.3005
R241 VTAIL.n309 VTAIL.n308 9.3005
R242 VTAIL.n286 VTAIL.n285 9.3005
R243 VTAIL.n303 VTAIL.n302 9.3005
R244 VTAIL.n301 VTAIL.n300 9.3005
R245 VTAIL.n290 VTAIL.n289 9.3005
R246 VTAIL.n295 VTAIL.n294 9.3005
R247 VTAIL.n282 VTAIL.n281 9.3005
R248 VTAIL.n37 VTAIL.n36 9.3005
R249 VTAIL.n31 VTAIL.n30 9.3005
R250 VTAIL.n29 VTAIL.n28 9.3005
R251 VTAIL.n6 VTAIL.n5 9.3005
R252 VTAIL.n23 VTAIL.n22 9.3005
R253 VTAIL.n21 VTAIL.n20 9.3005
R254 VTAIL.n10 VTAIL.n9 9.3005
R255 VTAIL.n15 VTAIL.n14 9.3005
R256 VTAIL.n2 VTAIL.n1 9.3005
R257 VTAIL.n77 VTAIL.n76 9.3005
R258 VTAIL.n71 VTAIL.n70 9.3005
R259 VTAIL.n69 VTAIL.n68 9.3005
R260 VTAIL.n46 VTAIL.n45 9.3005
R261 VTAIL.n63 VTAIL.n62 9.3005
R262 VTAIL.n61 VTAIL.n60 9.3005
R263 VTAIL.n50 VTAIL.n49 9.3005
R264 VTAIL.n55 VTAIL.n54 9.3005
R265 VTAIL.n42 VTAIL.n41 9.3005
R266 VTAIL.n117 VTAIL.n116 9.3005
R267 VTAIL.n111 VTAIL.n110 9.3005
R268 VTAIL.n109 VTAIL.n108 9.3005
R269 VTAIL.n86 VTAIL.n85 9.3005
R270 VTAIL.n103 VTAIL.n102 9.3005
R271 VTAIL.n101 VTAIL.n100 9.3005
R272 VTAIL.n90 VTAIL.n89 9.3005
R273 VTAIL.n95 VTAIL.n94 9.3005
R274 VTAIL.n82 VTAIL.n81 9.3005
R275 VTAIL.n277 VTAIL.n276 9.3005
R276 VTAIL.n242 VTAIL.n241 9.3005
R277 VTAIL.n271 VTAIL.n270 9.3005
R278 VTAIL.n269 VTAIL.n268 9.3005
R279 VTAIL.n246 VTAIL.n245 9.3005
R280 VTAIL.n263 VTAIL.n262 9.3005
R281 VTAIL.n261 VTAIL.n260 9.3005
R282 VTAIL.n250 VTAIL.n249 9.3005
R283 VTAIL.n255 VTAIL.n254 9.3005
R284 VTAIL.n237 VTAIL.n236 9.3005
R285 VTAIL.n202 VTAIL.n201 9.3005
R286 VTAIL.n231 VTAIL.n230 9.3005
R287 VTAIL.n229 VTAIL.n228 9.3005
R288 VTAIL.n206 VTAIL.n205 9.3005
R289 VTAIL.n223 VTAIL.n222 9.3005
R290 VTAIL.n221 VTAIL.n220 9.3005
R291 VTAIL.n210 VTAIL.n209 9.3005
R292 VTAIL.n215 VTAIL.n214 9.3005
R293 VTAIL.n197 VTAIL.n196 9.3005
R294 VTAIL.n162 VTAIL.n161 9.3005
R295 VTAIL.n191 VTAIL.n190 9.3005
R296 VTAIL.n189 VTAIL.n188 9.3005
R297 VTAIL.n166 VTAIL.n165 9.3005
R298 VTAIL.n183 VTAIL.n182 9.3005
R299 VTAIL.n181 VTAIL.n180 9.3005
R300 VTAIL.n170 VTAIL.n169 9.3005
R301 VTAIL.n175 VTAIL.n174 9.3005
R302 VTAIL.n157 VTAIL.n156 9.3005
R303 VTAIL.n122 VTAIL.n121 9.3005
R304 VTAIL.n151 VTAIL.n150 9.3005
R305 VTAIL.n149 VTAIL.n148 9.3005
R306 VTAIL.n126 VTAIL.n125 9.3005
R307 VTAIL.n143 VTAIL.n142 9.3005
R308 VTAIL.n141 VTAIL.n140 9.3005
R309 VTAIL.n130 VTAIL.n129 9.3005
R310 VTAIL.n135 VTAIL.n134 9.3005
R311 VTAIL.n308 VTAIL.n284 8.92171
R312 VTAIL.n28 VTAIL.n4 8.92171
R313 VTAIL.n68 VTAIL.n44 8.92171
R314 VTAIL.n108 VTAIL.n84 8.92171
R315 VTAIL.n268 VTAIL.n244 8.92171
R316 VTAIL.n228 VTAIL.n204 8.92171
R317 VTAIL.n188 VTAIL.n164 8.92171
R318 VTAIL.n148 VTAIL.n124 8.92171
R319 VTAIL.n312 VTAIL.n311 8.14595
R320 VTAIL.n32 VTAIL.n31 8.14595
R321 VTAIL.n72 VTAIL.n71 8.14595
R322 VTAIL.n112 VTAIL.n111 8.14595
R323 VTAIL.n272 VTAIL.n271 8.14595
R324 VTAIL.n232 VTAIL.n231 8.14595
R325 VTAIL.n192 VTAIL.n191 8.14595
R326 VTAIL.n152 VTAIL.n151 8.14595
R327 VTAIL.n315 VTAIL.n282 7.3702
R328 VTAIL.n318 VTAIL.n280 7.3702
R329 VTAIL.n35 VTAIL.n2 7.3702
R330 VTAIL.n38 VTAIL.n0 7.3702
R331 VTAIL.n75 VTAIL.n42 7.3702
R332 VTAIL.n78 VTAIL.n40 7.3702
R333 VTAIL.n115 VTAIL.n82 7.3702
R334 VTAIL.n118 VTAIL.n80 7.3702
R335 VTAIL.n278 VTAIL.n240 7.3702
R336 VTAIL.n275 VTAIL.n242 7.3702
R337 VTAIL.n238 VTAIL.n200 7.3702
R338 VTAIL.n235 VTAIL.n202 7.3702
R339 VTAIL.n198 VTAIL.n160 7.3702
R340 VTAIL.n195 VTAIL.n162 7.3702
R341 VTAIL.n158 VTAIL.n120 7.3702
R342 VTAIL.n155 VTAIL.n122 7.3702
R343 VTAIL.n316 VTAIL.n315 6.59444
R344 VTAIL.n316 VTAIL.n280 6.59444
R345 VTAIL.n36 VTAIL.n35 6.59444
R346 VTAIL.n36 VTAIL.n0 6.59444
R347 VTAIL.n76 VTAIL.n75 6.59444
R348 VTAIL.n76 VTAIL.n40 6.59444
R349 VTAIL.n116 VTAIL.n115 6.59444
R350 VTAIL.n116 VTAIL.n80 6.59444
R351 VTAIL.n276 VTAIL.n240 6.59444
R352 VTAIL.n276 VTAIL.n275 6.59444
R353 VTAIL.n236 VTAIL.n200 6.59444
R354 VTAIL.n236 VTAIL.n235 6.59444
R355 VTAIL.n196 VTAIL.n160 6.59444
R356 VTAIL.n196 VTAIL.n195 6.59444
R357 VTAIL.n156 VTAIL.n120 6.59444
R358 VTAIL.n156 VTAIL.n155 6.59444
R359 VTAIL.n312 VTAIL.n282 5.81868
R360 VTAIL.n32 VTAIL.n2 5.81868
R361 VTAIL.n72 VTAIL.n42 5.81868
R362 VTAIL.n112 VTAIL.n82 5.81868
R363 VTAIL.n272 VTAIL.n242 5.81868
R364 VTAIL.n232 VTAIL.n202 5.81868
R365 VTAIL.n192 VTAIL.n162 5.81868
R366 VTAIL.n152 VTAIL.n122 5.81868
R367 VTAIL.n311 VTAIL.n284 5.04292
R368 VTAIL.n31 VTAIL.n4 5.04292
R369 VTAIL.n71 VTAIL.n44 5.04292
R370 VTAIL.n111 VTAIL.n84 5.04292
R371 VTAIL.n271 VTAIL.n244 5.04292
R372 VTAIL.n231 VTAIL.n204 5.04292
R373 VTAIL.n191 VTAIL.n164 5.04292
R374 VTAIL.n151 VTAIL.n124 5.04292
R375 VTAIL.n254 VTAIL.n253 4.38565
R376 VTAIL.n214 VTAIL.n213 4.38565
R377 VTAIL.n174 VTAIL.n173 4.38565
R378 VTAIL.n134 VTAIL.n133 4.38565
R379 VTAIL.n294 VTAIL.n293 4.38565
R380 VTAIL.n14 VTAIL.n13 4.38565
R381 VTAIL.n54 VTAIL.n53 4.38565
R382 VTAIL.n94 VTAIL.n93 4.38565
R383 VTAIL.n308 VTAIL.n307 4.26717
R384 VTAIL.n28 VTAIL.n27 4.26717
R385 VTAIL.n68 VTAIL.n67 4.26717
R386 VTAIL.n108 VTAIL.n107 4.26717
R387 VTAIL.n268 VTAIL.n267 4.26717
R388 VTAIL.n228 VTAIL.n227 4.26717
R389 VTAIL.n188 VTAIL.n187 4.26717
R390 VTAIL.n148 VTAIL.n147 4.26717
R391 VTAIL.n304 VTAIL.n286 3.49141
R392 VTAIL.n24 VTAIL.n6 3.49141
R393 VTAIL.n64 VTAIL.n46 3.49141
R394 VTAIL.n104 VTAIL.n86 3.49141
R395 VTAIL.n264 VTAIL.n246 3.49141
R396 VTAIL.n224 VTAIL.n206 3.49141
R397 VTAIL.n184 VTAIL.n166 3.49141
R398 VTAIL.n144 VTAIL.n126 3.49141
R399 VTAIL.n199 VTAIL.n159 2.91429
R400 VTAIL.n279 VTAIL.n239 2.91429
R401 VTAIL.n119 VTAIL.n79 2.91429
R402 VTAIL.n303 VTAIL.n288 2.71565
R403 VTAIL.n23 VTAIL.n8 2.71565
R404 VTAIL.n63 VTAIL.n48 2.71565
R405 VTAIL.n103 VTAIL.n88 2.71565
R406 VTAIL.n263 VTAIL.n248 2.71565
R407 VTAIL.n223 VTAIL.n208 2.71565
R408 VTAIL.n183 VTAIL.n168 2.71565
R409 VTAIL.n143 VTAIL.n128 2.71565
R410 VTAIL.n300 VTAIL.n299 1.93989
R411 VTAIL.n20 VTAIL.n19 1.93989
R412 VTAIL.n60 VTAIL.n59 1.93989
R413 VTAIL.n100 VTAIL.n99 1.93989
R414 VTAIL.n260 VTAIL.n259 1.93989
R415 VTAIL.n220 VTAIL.n219 1.93989
R416 VTAIL.n180 VTAIL.n179 1.93989
R417 VTAIL.n140 VTAIL.n139 1.93989
R418 VTAIL VTAIL.n39 1.51559
R419 VTAIL VTAIL.n319 1.39921
R420 VTAIL.n296 VTAIL.n290 1.16414
R421 VTAIL.n16 VTAIL.n10 1.16414
R422 VTAIL.n56 VTAIL.n50 1.16414
R423 VTAIL.n96 VTAIL.n90 1.16414
R424 VTAIL.n256 VTAIL.n250 1.16414
R425 VTAIL.n216 VTAIL.n210 1.16414
R426 VTAIL.n176 VTAIL.n170 1.16414
R427 VTAIL.n136 VTAIL.n130 1.16414
R428 VTAIL.n239 VTAIL.n199 0.470328
R429 VTAIL.n79 VTAIL.n39 0.470328
R430 VTAIL.n295 VTAIL.n292 0.388379
R431 VTAIL.n15 VTAIL.n12 0.388379
R432 VTAIL.n55 VTAIL.n52 0.388379
R433 VTAIL.n95 VTAIL.n92 0.388379
R434 VTAIL.n255 VTAIL.n252 0.388379
R435 VTAIL.n215 VTAIL.n212 0.388379
R436 VTAIL.n175 VTAIL.n172 0.388379
R437 VTAIL.n135 VTAIL.n132 0.388379
R438 VTAIL.n294 VTAIL.n289 0.155672
R439 VTAIL.n301 VTAIL.n289 0.155672
R440 VTAIL.n302 VTAIL.n301 0.155672
R441 VTAIL.n302 VTAIL.n285 0.155672
R442 VTAIL.n309 VTAIL.n285 0.155672
R443 VTAIL.n310 VTAIL.n309 0.155672
R444 VTAIL.n310 VTAIL.n281 0.155672
R445 VTAIL.n317 VTAIL.n281 0.155672
R446 VTAIL.n14 VTAIL.n9 0.155672
R447 VTAIL.n21 VTAIL.n9 0.155672
R448 VTAIL.n22 VTAIL.n21 0.155672
R449 VTAIL.n22 VTAIL.n5 0.155672
R450 VTAIL.n29 VTAIL.n5 0.155672
R451 VTAIL.n30 VTAIL.n29 0.155672
R452 VTAIL.n30 VTAIL.n1 0.155672
R453 VTAIL.n37 VTAIL.n1 0.155672
R454 VTAIL.n54 VTAIL.n49 0.155672
R455 VTAIL.n61 VTAIL.n49 0.155672
R456 VTAIL.n62 VTAIL.n61 0.155672
R457 VTAIL.n62 VTAIL.n45 0.155672
R458 VTAIL.n69 VTAIL.n45 0.155672
R459 VTAIL.n70 VTAIL.n69 0.155672
R460 VTAIL.n70 VTAIL.n41 0.155672
R461 VTAIL.n77 VTAIL.n41 0.155672
R462 VTAIL.n94 VTAIL.n89 0.155672
R463 VTAIL.n101 VTAIL.n89 0.155672
R464 VTAIL.n102 VTAIL.n101 0.155672
R465 VTAIL.n102 VTAIL.n85 0.155672
R466 VTAIL.n109 VTAIL.n85 0.155672
R467 VTAIL.n110 VTAIL.n109 0.155672
R468 VTAIL.n110 VTAIL.n81 0.155672
R469 VTAIL.n117 VTAIL.n81 0.155672
R470 VTAIL.n277 VTAIL.n241 0.155672
R471 VTAIL.n270 VTAIL.n241 0.155672
R472 VTAIL.n270 VTAIL.n269 0.155672
R473 VTAIL.n269 VTAIL.n245 0.155672
R474 VTAIL.n262 VTAIL.n245 0.155672
R475 VTAIL.n262 VTAIL.n261 0.155672
R476 VTAIL.n261 VTAIL.n249 0.155672
R477 VTAIL.n254 VTAIL.n249 0.155672
R478 VTAIL.n237 VTAIL.n201 0.155672
R479 VTAIL.n230 VTAIL.n201 0.155672
R480 VTAIL.n230 VTAIL.n229 0.155672
R481 VTAIL.n229 VTAIL.n205 0.155672
R482 VTAIL.n222 VTAIL.n205 0.155672
R483 VTAIL.n222 VTAIL.n221 0.155672
R484 VTAIL.n221 VTAIL.n209 0.155672
R485 VTAIL.n214 VTAIL.n209 0.155672
R486 VTAIL.n197 VTAIL.n161 0.155672
R487 VTAIL.n190 VTAIL.n161 0.155672
R488 VTAIL.n190 VTAIL.n189 0.155672
R489 VTAIL.n189 VTAIL.n165 0.155672
R490 VTAIL.n182 VTAIL.n165 0.155672
R491 VTAIL.n182 VTAIL.n181 0.155672
R492 VTAIL.n181 VTAIL.n169 0.155672
R493 VTAIL.n174 VTAIL.n169 0.155672
R494 VTAIL.n157 VTAIL.n121 0.155672
R495 VTAIL.n150 VTAIL.n121 0.155672
R496 VTAIL.n150 VTAIL.n149 0.155672
R497 VTAIL.n149 VTAIL.n125 0.155672
R498 VTAIL.n142 VTAIL.n125 0.155672
R499 VTAIL.n142 VTAIL.n141 0.155672
R500 VTAIL.n141 VTAIL.n129 0.155672
R501 VTAIL.n134 VTAIL.n129 0.155672
R502 B.n513 B.n108 585
R503 B.n108 B.n71 585
R504 B.n515 B.n514 585
R505 B.n517 B.n107 585
R506 B.n520 B.n519 585
R507 B.n521 B.n106 585
R508 B.n523 B.n522 585
R509 B.n525 B.n105 585
R510 B.n528 B.n527 585
R511 B.n529 B.n104 585
R512 B.n531 B.n530 585
R513 B.n533 B.n103 585
R514 B.n536 B.n535 585
R515 B.n537 B.n102 585
R516 B.n539 B.n538 585
R517 B.n541 B.n101 585
R518 B.n544 B.n543 585
R519 B.n545 B.n100 585
R520 B.n547 B.n546 585
R521 B.n549 B.n99 585
R522 B.n552 B.n551 585
R523 B.n553 B.n98 585
R524 B.n555 B.n554 585
R525 B.n557 B.n97 585
R526 B.n560 B.n559 585
R527 B.n561 B.n96 585
R528 B.n563 B.n562 585
R529 B.n565 B.n95 585
R530 B.n568 B.n567 585
R531 B.n570 B.n92 585
R532 B.n572 B.n571 585
R533 B.n574 B.n91 585
R534 B.n577 B.n576 585
R535 B.n578 B.n90 585
R536 B.n580 B.n579 585
R537 B.n582 B.n89 585
R538 B.n585 B.n584 585
R539 B.n586 B.n86 585
R540 B.n589 B.n588 585
R541 B.n591 B.n85 585
R542 B.n594 B.n593 585
R543 B.n595 B.n84 585
R544 B.n597 B.n596 585
R545 B.n599 B.n83 585
R546 B.n602 B.n601 585
R547 B.n603 B.n82 585
R548 B.n605 B.n604 585
R549 B.n607 B.n81 585
R550 B.n610 B.n609 585
R551 B.n611 B.n80 585
R552 B.n613 B.n612 585
R553 B.n615 B.n79 585
R554 B.n618 B.n617 585
R555 B.n619 B.n78 585
R556 B.n621 B.n620 585
R557 B.n623 B.n77 585
R558 B.n626 B.n625 585
R559 B.n627 B.n76 585
R560 B.n629 B.n628 585
R561 B.n631 B.n75 585
R562 B.n634 B.n633 585
R563 B.n635 B.n74 585
R564 B.n637 B.n636 585
R565 B.n639 B.n73 585
R566 B.n642 B.n641 585
R567 B.n643 B.n72 585
R568 B.n512 B.n70 585
R569 B.n646 B.n70 585
R570 B.n511 B.n69 585
R571 B.n647 B.n69 585
R572 B.n510 B.n68 585
R573 B.n648 B.n68 585
R574 B.n509 B.n508 585
R575 B.n508 B.n64 585
R576 B.n507 B.n63 585
R577 B.n654 B.n63 585
R578 B.n506 B.n62 585
R579 B.n655 B.n62 585
R580 B.n505 B.n61 585
R581 B.n656 B.n61 585
R582 B.n504 B.n503 585
R583 B.n503 B.n57 585
R584 B.n502 B.n56 585
R585 B.n662 B.n56 585
R586 B.n501 B.n55 585
R587 B.n663 B.n55 585
R588 B.n500 B.n54 585
R589 B.n664 B.n54 585
R590 B.n499 B.n498 585
R591 B.n498 B.n50 585
R592 B.n497 B.n49 585
R593 B.n670 B.n49 585
R594 B.n496 B.n48 585
R595 B.n671 B.n48 585
R596 B.n495 B.n47 585
R597 B.n672 B.n47 585
R598 B.n494 B.n493 585
R599 B.n493 B.n43 585
R600 B.n492 B.n42 585
R601 B.n678 B.n42 585
R602 B.n491 B.n41 585
R603 B.n679 B.n41 585
R604 B.n490 B.n40 585
R605 B.n680 B.n40 585
R606 B.n489 B.n488 585
R607 B.n488 B.n36 585
R608 B.n487 B.n35 585
R609 B.n686 B.n35 585
R610 B.n486 B.n34 585
R611 B.n687 B.n34 585
R612 B.n485 B.n33 585
R613 B.n688 B.n33 585
R614 B.n484 B.n483 585
R615 B.n483 B.n29 585
R616 B.n482 B.n28 585
R617 B.n694 B.n28 585
R618 B.n481 B.n27 585
R619 B.n695 B.n27 585
R620 B.n480 B.n26 585
R621 B.n696 B.n26 585
R622 B.n479 B.n478 585
R623 B.n478 B.n22 585
R624 B.n477 B.n21 585
R625 B.n702 B.n21 585
R626 B.n476 B.n20 585
R627 B.n703 B.n20 585
R628 B.n475 B.n19 585
R629 B.n704 B.n19 585
R630 B.n474 B.n473 585
R631 B.n473 B.n18 585
R632 B.n472 B.n14 585
R633 B.n710 B.n14 585
R634 B.n471 B.n13 585
R635 B.n711 B.n13 585
R636 B.n470 B.n12 585
R637 B.n712 B.n12 585
R638 B.n469 B.n468 585
R639 B.n468 B.n8 585
R640 B.n467 B.n7 585
R641 B.n718 B.n7 585
R642 B.n466 B.n6 585
R643 B.n719 B.n6 585
R644 B.n465 B.n5 585
R645 B.n720 B.n5 585
R646 B.n464 B.n463 585
R647 B.n463 B.n4 585
R648 B.n462 B.n109 585
R649 B.n462 B.n461 585
R650 B.n452 B.n110 585
R651 B.n111 B.n110 585
R652 B.n454 B.n453 585
R653 B.n455 B.n454 585
R654 B.n451 B.n116 585
R655 B.n116 B.n115 585
R656 B.n450 B.n449 585
R657 B.n449 B.n448 585
R658 B.n118 B.n117 585
R659 B.n441 B.n118 585
R660 B.n440 B.n439 585
R661 B.n442 B.n440 585
R662 B.n438 B.n123 585
R663 B.n123 B.n122 585
R664 B.n437 B.n436 585
R665 B.n436 B.n435 585
R666 B.n125 B.n124 585
R667 B.n126 B.n125 585
R668 B.n428 B.n427 585
R669 B.n429 B.n428 585
R670 B.n426 B.n131 585
R671 B.n131 B.n130 585
R672 B.n425 B.n424 585
R673 B.n424 B.n423 585
R674 B.n133 B.n132 585
R675 B.n134 B.n133 585
R676 B.n416 B.n415 585
R677 B.n417 B.n416 585
R678 B.n414 B.n138 585
R679 B.n142 B.n138 585
R680 B.n413 B.n412 585
R681 B.n412 B.n411 585
R682 B.n140 B.n139 585
R683 B.n141 B.n140 585
R684 B.n404 B.n403 585
R685 B.n405 B.n404 585
R686 B.n402 B.n147 585
R687 B.n147 B.n146 585
R688 B.n401 B.n400 585
R689 B.n400 B.n399 585
R690 B.n149 B.n148 585
R691 B.n150 B.n149 585
R692 B.n392 B.n391 585
R693 B.n393 B.n392 585
R694 B.n390 B.n155 585
R695 B.n155 B.n154 585
R696 B.n389 B.n388 585
R697 B.n388 B.n387 585
R698 B.n157 B.n156 585
R699 B.n158 B.n157 585
R700 B.n380 B.n379 585
R701 B.n381 B.n380 585
R702 B.n378 B.n163 585
R703 B.n163 B.n162 585
R704 B.n377 B.n376 585
R705 B.n376 B.n375 585
R706 B.n165 B.n164 585
R707 B.n166 B.n165 585
R708 B.n368 B.n367 585
R709 B.n369 B.n368 585
R710 B.n366 B.n171 585
R711 B.n171 B.n170 585
R712 B.n365 B.n364 585
R713 B.n364 B.n363 585
R714 B.n173 B.n172 585
R715 B.n174 B.n173 585
R716 B.n356 B.n355 585
R717 B.n357 B.n356 585
R718 B.n354 B.n179 585
R719 B.n179 B.n178 585
R720 B.n353 B.n352 585
R721 B.n352 B.n351 585
R722 B.n348 B.n183 585
R723 B.n347 B.n346 585
R724 B.n344 B.n184 585
R725 B.n344 B.n182 585
R726 B.n343 B.n342 585
R727 B.n341 B.n340 585
R728 B.n339 B.n186 585
R729 B.n337 B.n336 585
R730 B.n335 B.n187 585
R731 B.n334 B.n333 585
R732 B.n331 B.n188 585
R733 B.n329 B.n328 585
R734 B.n327 B.n189 585
R735 B.n326 B.n325 585
R736 B.n323 B.n190 585
R737 B.n321 B.n320 585
R738 B.n319 B.n191 585
R739 B.n318 B.n317 585
R740 B.n315 B.n192 585
R741 B.n313 B.n312 585
R742 B.n311 B.n193 585
R743 B.n310 B.n309 585
R744 B.n307 B.n194 585
R745 B.n305 B.n304 585
R746 B.n303 B.n195 585
R747 B.n302 B.n301 585
R748 B.n299 B.n196 585
R749 B.n297 B.n296 585
R750 B.n295 B.n197 585
R751 B.n293 B.n292 585
R752 B.n290 B.n200 585
R753 B.n288 B.n287 585
R754 B.n286 B.n201 585
R755 B.n285 B.n284 585
R756 B.n282 B.n202 585
R757 B.n280 B.n279 585
R758 B.n278 B.n203 585
R759 B.n277 B.n276 585
R760 B.n274 B.n273 585
R761 B.n272 B.n271 585
R762 B.n270 B.n208 585
R763 B.n268 B.n267 585
R764 B.n266 B.n209 585
R765 B.n265 B.n264 585
R766 B.n262 B.n210 585
R767 B.n260 B.n259 585
R768 B.n258 B.n211 585
R769 B.n257 B.n256 585
R770 B.n254 B.n212 585
R771 B.n252 B.n251 585
R772 B.n250 B.n213 585
R773 B.n249 B.n248 585
R774 B.n246 B.n214 585
R775 B.n244 B.n243 585
R776 B.n242 B.n215 585
R777 B.n241 B.n240 585
R778 B.n238 B.n216 585
R779 B.n236 B.n235 585
R780 B.n234 B.n217 585
R781 B.n233 B.n232 585
R782 B.n230 B.n218 585
R783 B.n228 B.n227 585
R784 B.n226 B.n219 585
R785 B.n225 B.n224 585
R786 B.n222 B.n220 585
R787 B.n181 B.n180 585
R788 B.n350 B.n349 585
R789 B.n351 B.n350 585
R790 B.n177 B.n176 585
R791 B.n178 B.n177 585
R792 B.n359 B.n358 585
R793 B.n358 B.n357 585
R794 B.n360 B.n175 585
R795 B.n175 B.n174 585
R796 B.n362 B.n361 585
R797 B.n363 B.n362 585
R798 B.n169 B.n168 585
R799 B.n170 B.n169 585
R800 B.n371 B.n370 585
R801 B.n370 B.n369 585
R802 B.n372 B.n167 585
R803 B.n167 B.n166 585
R804 B.n374 B.n373 585
R805 B.n375 B.n374 585
R806 B.n161 B.n160 585
R807 B.n162 B.n161 585
R808 B.n383 B.n382 585
R809 B.n382 B.n381 585
R810 B.n384 B.n159 585
R811 B.n159 B.n158 585
R812 B.n386 B.n385 585
R813 B.n387 B.n386 585
R814 B.n153 B.n152 585
R815 B.n154 B.n153 585
R816 B.n395 B.n394 585
R817 B.n394 B.n393 585
R818 B.n396 B.n151 585
R819 B.n151 B.n150 585
R820 B.n398 B.n397 585
R821 B.n399 B.n398 585
R822 B.n145 B.n144 585
R823 B.n146 B.n145 585
R824 B.n407 B.n406 585
R825 B.n406 B.n405 585
R826 B.n408 B.n143 585
R827 B.n143 B.n141 585
R828 B.n410 B.n409 585
R829 B.n411 B.n410 585
R830 B.n137 B.n136 585
R831 B.n142 B.n137 585
R832 B.n419 B.n418 585
R833 B.n418 B.n417 585
R834 B.n420 B.n135 585
R835 B.n135 B.n134 585
R836 B.n422 B.n421 585
R837 B.n423 B.n422 585
R838 B.n129 B.n128 585
R839 B.n130 B.n129 585
R840 B.n431 B.n430 585
R841 B.n430 B.n429 585
R842 B.n432 B.n127 585
R843 B.n127 B.n126 585
R844 B.n434 B.n433 585
R845 B.n435 B.n434 585
R846 B.n121 B.n120 585
R847 B.n122 B.n121 585
R848 B.n444 B.n443 585
R849 B.n443 B.n442 585
R850 B.n445 B.n119 585
R851 B.n441 B.n119 585
R852 B.n447 B.n446 585
R853 B.n448 B.n447 585
R854 B.n114 B.n113 585
R855 B.n115 B.n114 585
R856 B.n457 B.n456 585
R857 B.n456 B.n455 585
R858 B.n458 B.n112 585
R859 B.n112 B.n111 585
R860 B.n460 B.n459 585
R861 B.n461 B.n460 585
R862 B.n2 B.n0 585
R863 B.n4 B.n2 585
R864 B.n3 B.n1 585
R865 B.n719 B.n3 585
R866 B.n717 B.n716 585
R867 B.n718 B.n717 585
R868 B.n715 B.n9 585
R869 B.n9 B.n8 585
R870 B.n714 B.n713 585
R871 B.n713 B.n712 585
R872 B.n11 B.n10 585
R873 B.n711 B.n11 585
R874 B.n709 B.n708 585
R875 B.n710 B.n709 585
R876 B.n707 B.n15 585
R877 B.n18 B.n15 585
R878 B.n706 B.n705 585
R879 B.n705 B.n704 585
R880 B.n17 B.n16 585
R881 B.n703 B.n17 585
R882 B.n701 B.n700 585
R883 B.n702 B.n701 585
R884 B.n699 B.n23 585
R885 B.n23 B.n22 585
R886 B.n698 B.n697 585
R887 B.n697 B.n696 585
R888 B.n25 B.n24 585
R889 B.n695 B.n25 585
R890 B.n693 B.n692 585
R891 B.n694 B.n693 585
R892 B.n691 B.n30 585
R893 B.n30 B.n29 585
R894 B.n690 B.n689 585
R895 B.n689 B.n688 585
R896 B.n32 B.n31 585
R897 B.n687 B.n32 585
R898 B.n685 B.n684 585
R899 B.n686 B.n685 585
R900 B.n683 B.n37 585
R901 B.n37 B.n36 585
R902 B.n682 B.n681 585
R903 B.n681 B.n680 585
R904 B.n39 B.n38 585
R905 B.n679 B.n39 585
R906 B.n677 B.n676 585
R907 B.n678 B.n677 585
R908 B.n675 B.n44 585
R909 B.n44 B.n43 585
R910 B.n674 B.n673 585
R911 B.n673 B.n672 585
R912 B.n46 B.n45 585
R913 B.n671 B.n46 585
R914 B.n669 B.n668 585
R915 B.n670 B.n669 585
R916 B.n667 B.n51 585
R917 B.n51 B.n50 585
R918 B.n666 B.n665 585
R919 B.n665 B.n664 585
R920 B.n53 B.n52 585
R921 B.n663 B.n53 585
R922 B.n661 B.n660 585
R923 B.n662 B.n661 585
R924 B.n659 B.n58 585
R925 B.n58 B.n57 585
R926 B.n658 B.n657 585
R927 B.n657 B.n656 585
R928 B.n60 B.n59 585
R929 B.n655 B.n60 585
R930 B.n653 B.n652 585
R931 B.n654 B.n653 585
R932 B.n651 B.n65 585
R933 B.n65 B.n64 585
R934 B.n650 B.n649 585
R935 B.n649 B.n648 585
R936 B.n67 B.n66 585
R937 B.n647 B.n67 585
R938 B.n645 B.n644 585
R939 B.n646 B.n645 585
R940 B.n722 B.n721 585
R941 B.n721 B.n720 585
R942 B.n350 B.n183 526.135
R943 B.n645 B.n72 526.135
R944 B.n352 B.n181 526.135
R945 B.n108 B.n70 526.135
R946 B.n204 B.t10 267.719
R947 B.n93 B.t13 267.719
R948 B.n198 B.t7 267.719
R949 B.n87 B.t16 267.719
R950 B.n204 B.t8 266.716
R951 B.n198 B.t4 266.716
R952 B.n87 B.t15 266.716
R953 B.n93 B.t11 266.716
R954 B.n516 B.n71 256.663
R955 B.n518 B.n71 256.663
R956 B.n524 B.n71 256.663
R957 B.n526 B.n71 256.663
R958 B.n532 B.n71 256.663
R959 B.n534 B.n71 256.663
R960 B.n540 B.n71 256.663
R961 B.n542 B.n71 256.663
R962 B.n548 B.n71 256.663
R963 B.n550 B.n71 256.663
R964 B.n556 B.n71 256.663
R965 B.n558 B.n71 256.663
R966 B.n564 B.n71 256.663
R967 B.n566 B.n71 256.663
R968 B.n573 B.n71 256.663
R969 B.n575 B.n71 256.663
R970 B.n581 B.n71 256.663
R971 B.n583 B.n71 256.663
R972 B.n590 B.n71 256.663
R973 B.n592 B.n71 256.663
R974 B.n598 B.n71 256.663
R975 B.n600 B.n71 256.663
R976 B.n606 B.n71 256.663
R977 B.n608 B.n71 256.663
R978 B.n614 B.n71 256.663
R979 B.n616 B.n71 256.663
R980 B.n622 B.n71 256.663
R981 B.n624 B.n71 256.663
R982 B.n630 B.n71 256.663
R983 B.n632 B.n71 256.663
R984 B.n638 B.n71 256.663
R985 B.n640 B.n71 256.663
R986 B.n345 B.n182 256.663
R987 B.n185 B.n182 256.663
R988 B.n338 B.n182 256.663
R989 B.n332 B.n182 256.663
R990 B.n330 B.n182 256.663
R991 B.n324 B.n182 256.663
R992 B.n322 B.n182 256.663
R993 B.n316 B.n182 256.663
R994 B.n314 B.n182 256.663
R995 B.n308 B.n182 256.663
R996 B.n306 B.n182 256.663
R997 B.n300 B.n182 256.663
R998 B.n298 B.n182 256.663
R999 B.n291 B.n182 256.663
R1000 B.n289 B.n182 256.663
R1001 B.n283 B.n182 256.663
R1002 B.n281 B.n182 256.663
R1003 B.n275 B.n182 256.663
R1004 B.n207 B.n182 256.663
R1005 B.n269 B.n182 256.663
R1006 B.n263 B.n182 256.663
R1007 B.n261 B.n182 256.663
R1008 B.n255 B.n182 256.663
R1009 B.n253 B.n182 256.663
R1010 B.n247 B.n182 256.663
R1011 B.n245 B.n182 256.663
R1012 B.n239 B.n182 256.663
R1013 B.n237 B.n182 256.663
R1014 B.n231 B.n182 256.663
R1015 B.n229 B.n182 256.663
R1016 B.n223 B.n182 256.663
R1017 B.n221 B.n182 256.663
R1018 B.n205 B.t9 202.167
R1019 B.n94 B.t14 202.167
R1020 B.n199 B.t6 202.167
R1021 B.n88 B.t17 202.167
R1022 B.n350 B.n177 163.367
R1023 B.n358 B.n177 163.367
R1024 B.n358 B.n175 163.367
R1025 B.n362 B.n175 163.367
R1026 B.n362 B.n169 163.367
R1027 B.n370 B.n169 163.367
R1028 B.n370 B.n167 163.367
R1029 B.n374 B.n167 163.367
R1030 B.n374 B.n161 163.367
R1031 B.n382 B.n161 163.367
R1032 B.n382 B.n159 163.367
R1033 B.n386 B.n159 163.367
R1034 B.n386 B.n153 163.367
R1035 B.n394 B.n153 163.367
R1036 B.n394 B.n151 163.367
R1037 B.n398 B.n151 163.367
R1038 B.n398 B.n145 163.367
R1039 B.n406 B.n145 163.367
R1040 B.n406 B.n143 163.367
R1041 B.n410 B.n143 163.367
R1042 B.n410 B.n137 163.367
R1043 B.n418 B.n137 163.367
R1044 B.n418 B.n135 163.367
R1045 B.n422 B.n135 163.367
R1046 B.n422 B.n129 163.367
R1047 B.n430 B.n129 163.367
R1048 B.n430 B.n127 163.367
R1049 B.n434 B.n127 163.367
R1050 B.n434 B.n121 163.367
R1051 B.n443 B.n121 163.367
R1052 B.n443 B.n119 163.367
R1053 B.n447 B.n119 163.367
R1054 B.n447 B.n114 163.367
R1055 B.n456 B.n114 163.367
R1056 B.n456 B.n112 163.367
R1057 B.n460 B.n112 163.367
R1058 B.n460 B.n2 163.367
R1059 B.n721 B.n2 163.367
R1060 B.n721 B.n3 163.367
R1061 B.n717 B.n3 163.367
R1062 B.n717 B.n9 163.367
R1063 B.n713 B.n9 163.367
R1064 B.n713 B.n11 163.367
R1065 B.n709 B.n11 163.367
R1066 B.n709 B.n15 163.367
R1067 B.n705 B.n15 163.367
R1068 B.n705 B.n17 163.367
R1069 B.n701 B.n17 163.367
R1070 B.n701 B.n23 163.367
R1071 B.n697 B.n23 163.367
R1072 B.n697 B.n25 163.367
R1073 B.n693 B.n25 163.367
R1074 B.n693 B.n30 163.367
R1075 B.n689 B.n30 163.367
R1076 B.n689 B.n32 163.367
R1077 B.n685 B.n32 163.367
R1078 B.n685 B.n37 163.367
R1079 B.n681 B.n37 163.367
R1080 B.n681 B.n39 163.367
R1081 B.n677 B.n39 163.367
R1082 B.n677 B.n44 163.367
R1083 B.n673 B.n44 163.367
R1084 B.n673 B.n46 163.367
R1085 B.n669 B.n46 163.367
R1086 B.n669 B.n51 163.367
R1087 B.n665 B.n51 163.367
R1088 B.n665 B.n53 163.367
R1089 B.n661 B.n53 163.367
R1090 B.n661 B.n58 163.367
R1091 B.n657 B.n58 163.367
R1092 B.n657 B.n60 163.367
R1093 B.n653 B.n60 163.367
R1094 B.n653 B.n65 163.367
R1095 B.n649 B.n65 163.367
R1096 B.n649 B.n67 163.367
R1097 B.n645 B.n67 163.367
R1098 B.n346 B.n344 163.367
R1099 B.n344 B.n343 163.367
R1100 B.n340 B.n339 163.367
R1101 B.n337 B.n187 163.367
R1102 B.n333 B.n331 163.367
R1103 B.n329 B.n189 163.367
R1104 B.n325 B.n323 163.367
R1105 B.n321 B.n191 163.367
R1106 B.n317 B.n315 163.367
R1107 B.n313 B.n193 163.367
R1108 B.n309 B.n307 163.367
R1109 B.n305 B.n195 163.367
R1110 B.n301 B.n299 163.367
R1111 B.n297 B.n197 163.367
R1112 B.n292 B.n290 163.367
R1113 B.n288 B.n201 163.367
R1114 B.n284 B.n282 163.367
R1115 B.n280 B.n203 163.367
R1116 B.n276 B.n274 163.367
R1117 B.n271 B.n270 163.367
R1118 B.n268 B.n209 163.367
R1119 B.n264 B.n262 163.367
R1120 B.n260 B.n211 163.367
R1121 B.n256 B.n254 163.367
R1122 B.n252 B.n213 163.367
R1123 B.n248 B.n246 163.367
R1124 B.n244 B.n215 163.367
R1125 B.n240 B.n238 163.367
R1126 B.n236 B.n217 163.367
R1127 B.n232 B.n230 163.367
R1128 B.n228 B.n219 163.367
R1129 B.n224 B.n222 163.367
R1130 B.n352 B.n179 163.367
R1131 B.n356 B.n179 163.367
R1132 B.n356 B.n173 163.367
R1133 B.n364 B.n173 163.367
R1134 B.n364 B.n171 163.367
R1135 B.n368 B.n171 163.367
R1136 B.n368 B.n165 163.367
R1137 B.n376 B.n165 163.367
R1138 B.n376 B.n163 163.367
R1139 B.n380 B.n163 163.367
R1140 B.n380 B.n157 163.367
R1141 B.n388 B.n157 163.367
R1142 B.n388 B.n155 163.367
R1143 B.n392 B.n155 163.367
R1144 B.n392 B.n149 163.367
R1145 B.n400 B.n149 163.367
R1146 B.n400 B.n147 163.367
R1147 B.n404 B.n147 163.367
R1148 B.n404 B.n140 163.367
R1149 B.n412 B.n140 163.367
R1150 B.n412 B.n138 163.367
R1151 B.n416 B.n138 163.367
R1152 B.n416 B.n133 163.367
R1153 B.n424 B.n133 163.367
R1154 B.n424 B.n131 163.367
R1155 B.n428 B.n131 163.367
R1156 B.n428 B.n125 163.367
R1157 B.n436 B.n125 163.367
R1158 B.n436 B.n123 163.367
R1159 B.n440 B.n123 163.367
R1160 B.n440 B.n118 163.367
R1161 B.n449 B.n118 163.367
R1162 B.n449 B.n116 163.367
R1163 B.n454 B.n116 163.367
R1164 B.n454 B.n110 163.367
R1165 B.n462 B.n110 163.367
R1166 B.n463 B.n462 163.367
R1167 B.n463 B.n5 163.367
R1168 B.n6 B.n5 163.367
R1169 B.n7 B.n6 163.367
R1170 B.n468 B.n7 163.367
R1171 B.n468 B.n12 163.367
R1172 B.n13 B.n12 163.367
R1173 B.n14 B.n13 163.367
R1174 B.n473 B.n14 163.367
R1175 B.n473 B.n19 163.367
R1176 B.n20 B.n19 163.367
R1177 B.n21 B.n20 163.367
R1178 B.n478 B.n21 163.367
R1179 B.n478 B.n26 163.367
R1180 B.n27 B.n26 163.367
R1181 B.n28 B.n27 163.367
R1182 B.n483 B.n28 163.367
R1183 B.n483 B.n33 163.367
R1184 B.n34 B.n33 163.367
R1185 B.n35 B.n34 163.367
R1186 B.n488 B.n35 163.367
R1187 B.n488 B.n40 163.367
R1188 B.n41 B.n40 163.367
R1189 B.n42 B.n41 163.367
R1190 B.n493 B.n42 163.367
R1191 B.n493 B.n47 163.367
R1192 B.n48 B.n47 163.367
R1193 B.n49 B.n48 163.367
R1194 B.n498 B.n49 163.367
R1195 B.n498 B.n54 163.367
R1196 B.n55 B.n54 163.367
R1197 B.n56 B.n55 163.367
R1198 B.n503 B.n56 163.367
R1199 B.n503 B.n61 163.367
R1200 B.n62 B.n61 163.367
R1201 B.n63 B.n62 163.367
R1202 B.n508 B.n63 163.367
R1203 B.n508 B.n68 163.367
R1204 B.n69 B.n68 163.367
R1205 B.n70 B.n69 163.367
R1206 B.n641 B.n639 163.367
R1207 B.n637 B.n74 163.367
R1208 B.n633 B.n631 163.367
R1209 B.n629 B.n76 163.367
R1210 B.n625 B.n623 163.367
R1211 B.n621 B.n78 163.367
R1212 B.n617 B.n615 163.367
R1213 B.n613 B.n80 163.367
R1214 B.n609 B.n607 163.367
R1215 B.n605 B.n82 163.367
R1216 B.n601 B.n599 163.367
R1217 B.n597 B.n84 163.367
R1218 B.n593 B.n591 163.367
R1219 B.n589 B.n86 163.367
R1220 B.n584 B.n582 163.367
R1221 B.n580 B.n90 163.367
R1222 B.n576 B.n574 163.367
R1223 B.n572 B.n92 163.367
R1224 B.n567 B.n565 163.367
R1225 B.n563 B.n96 163.367
R1226 B.n559 B.n557 163.367
R1227 B.n555 B.n98 163.367
R1228 B.n551 B.n549 163.367
R1229 B.n547 B.n100 163.367
R1230 B.n543 B.n541 163.367
R1231 B.n539 B.n102 163.367
R1232 B.n535 B.n533 163.367
R1233 B.n531 B.n104 163.367
R1234 B.n527 B.n525 163.367
R1235 B.n523 B.n106 163.367
R1236 B.n519 B.n517 163.367
R1237 B.n515 B.n108 163.367
R1238 B.n351 B.n182 103.683
R1239 B.n646 B.n71 103.683
R1240 B.n345 B.n183 71.676
R1241 B.n343 B.n185 71.676
R1242 B.n339 B.n338 71.676
R1243 B.n332 B.n187 71.676
R1244 B.n331 B.n330 71.676
R1245 B.n324 B.n189 71.676
R1246 B.n323 B.n322 71.676
R1247 B.n316 B.n191 71.676
R1248 B.n315 B.n314 71.676
R1249 B.n308 B.n193 71.676
R1250 B.n307 B.n306 71.676
R1251 B.n300 B.n195 71.676
R1252 B.n299 B.n298 71.676
R1253 B.n291 B.n197 71.676
R1254 B.n290 B.n289 71.676
R1255 B.n283 B.n201 71.676
R1256 B.n282 B.n281 71.676
R1257 B.n275 B.n203 71.676
R1258 B.n274 B.n207 71.676
R1259 B.n270 B.n269 71.676
R1260 B.n263 B.n209 71.676
R1261 B.n262 B.n261 71.676
R1262 B.n255 B.n211 71.676
R1263 B.n254 B.n253 71.676
R1264 B.n247 B.n213 71.676
R1265 B.n246 B.n245 71.676
R1266 B.n239 B.n215 71.676
R1267 B.n238 B.n237 71.676
R1268 B.n231 B.n217 71.676
R1269 B.n230 B.n229 71.676
R1270 B.n223 B.n219 71.676
R1271 B.n222 B.n221 71.676
R1272 B.n640 B.n72 71.676
R1273 B.n639 B.n638 71.676
R1274 B.n632 B.n74 71.676
R1275 B.n631 B.n630 71.676
R1276 B.n624 B.n76 71.676
R1277 B.n623 B.n622 71.676
R1278 B.n616 B.n78 71.676
R1279 B.n615 B.n614 71.676
R1280 B.n608 B.n80 71.676
R1281 B.n607 B.n606 71.676
R1282 B.n600 B.n82 71.676
R1283 B.n599 B.n598 71.676
R1284 B.n592 B.n84 71.676
R1285 B.n591 B.n590 71.676
R1286 B.n583 B.n86 71.676
R1287 B.n582 B.n581 71.676
R1288 B.n575 B.n90 71.676
R1289 B.n574 B.n573 71.676
R1290 B.n566 B.n92 71.676
R1291 B.n565 B.n564 71.676
R1292 B.n558 B.n96 71.676
R1293 B.n557 B.n556 71.676
R1294 B.n550 B.n98 71.676
R1295 B.n549 B.n548 71.676
R1296 B.n542 B.n100 71.676
R1297 B.n541 B.n540 71.676
R1298 B.n534 B.n102 71.676
R1299 B.n533 B.n532 71.676
R1300 B.n526 B.n104 71.676
R1301 B.n525 B.n524 71.676
R1302 B.n518 B.n106 71.676
R1303 B.n517 B.n516 71.676
R1304 B.n516 B.n515 71.676
R1305 B.n519 B.n518 71.676
R1306 B.n524 B.n523 71.676
R1307 B.n527 B.n526 71.676
R1308 B.n532 B.n531 71.676
R1309 B.n535 B.n534 71.676
R1310 B.n540 B.n539 71.676
R1311 B.n543 B.n542 71.676
R1312 B.n548 B.n547 71.676
R1313 B.n551 B.n550 71.676
R1314 B.n556 B.n555 71.676
R1315 B.n559 B.n558 71.676
R1316 B.n564 B.n563 71.676
R1317 B.n567 B.n566 71.676
R1318 B.n573 B.n572 71.676
R1319 B.n576 B.n575 71.676
R1320 B.n581 B.n580 71.676
R1321 B.n584 B.n583 71.676
R1322 B.n590 B.n589 71.676
R1323 B.n593 B.n592 71.676
R1324 B.n598 B.n597 71.676
R1325 B.n601 B.n600 71.676
R1326 B.n606 B.n605 71.676
R1327 B.n609 B.n608 71.676
R1328 B.n614 B.n613 71.676
R1329 B.n617 B.n616 71.676
R1330 B.n622 B.n621 71.676
R1331 B.n625 B.n624 71.676
R1332 B.n630 B.n629 71.676
R1333 B.n633 B.n632 71.676
R1334 B.n638 B.n637 71.676
R1335 B.n641 B.n640 71.676
R1336 B.n346 B.n345 71.676
R1337 B.n340 B.n185 71.676
R1338 B.n338 B.n337 71.676
R1339 B.n333 B.n332 71.676
R1340 B.n330 B.n329 71.676
R1341 B.n325 B.n324 71.676
R1342 B.n322 B.n321 71.676
R1343 B.n317 B.n316 71.676
R1344 B.n314 B.n313 71.676
R1345 B.n309 B.n308 71.676
R1346 B.n306 B.n305 71.676
R1347 B.n301 B.n300 71.676
R1348 B.n298 B.n297 71.676
R1349 B.n292 B.n291 71.676
R1350 B.n289 B.n288 71.676
R1351 B.n284 B.n283 71.676
R1352 B.n281 B.n280 71.676
R1353 B.n276 B.n275 71.676
R1354 B.n271 B.n207 71.676
R1355 B.n269 B.n268 71.676
R1356 B.n264 B.n263 71.676
R1357 B.n261 B.n260 71.676
R1358 B.n256 B.n255 71.676
R1359 B.n253 B.n252 71.676
R1360 B.n248 B.n247 71.676
R1361 B.n245 B.n244 71.676
R1362 B.n240 B.n239 71.676
R1363 B.n237 B.n236 71.676
R1364 B.n232 B.n231 71.676
R1365 B.n229 B.n228 71.676
R1366 B.n224 B.n223 71.676
R1367 B.n221 B.n181 71.676
R1368 B.n205 B.n204 65.552
R1369 B.n199 B.n198 65.552
R1370 B.n88 B.n87 65.552
R1371 B.n94 B.n93 65.552
R1372 B.n206 B.n205 59.5399
R1373 B.n294 B.n199 59.5399
R1374 B.n587 B.n88 59.5399
R1375 B.n569 B.n94 59.5399
R1376 B.n351 B.n178 59.248
R1377 B.n357 B.n178 59.248
R1378 B.n357 B.n174 59.248
R1379 B.n363 B.n174 59.248
R1380 B.n363 B.n170 59.248
R1381 B.n369 B.n170 59.248
R1382 B.n369 B.n166 59.248
R1383 B.n375 B.n166 59.248
R1384 B.n381 B.n162 59.248
R1385 B.n381 B.n158 59.248
R1386 B.n387 B.n158 59.248
R1387 B.n387 B.n154 59.248
R1388 B.n393 B.n154 59.248
R1389 B.n393 B.n150 59.248
R1390 B.n399 B.n150 59.248
R1391 B.n399 B.n146 59.248
R1392 B.n405 B.n146 59.248
R1393 B.n405 B.n141 59.248
R1394 B.n411 B.n141 59.248
R1395 B.n411 B.n142 59.248
R1396 B.n417 B.n134 59.248
R1397 B.n423 B.n134 59.248
R1398 B.n423 B.n130 59.248
R1399 B.n429 B.n130 59.248
R1400 B.n429 B.n126 59.248
R1401 B.n435 B.n126 59.248
R1402 B.n435 B.n122 59.248
R1403 B.n442 B.n122 59.248
R1404 B.n442 B.n441 59.248
R1405 B.n448 B.n115 59.248
R1406 B.n455 B.n115 59.248
R1407 B.n455 B.n111 59.248
R1408 B.n461 B.n111 59.248
R1409 B.n461 B.n4 59.248
R1410 B.n720 B.n4 59.248
R1411 B.n720 B.n719 59.248
R1412 B.n719 B.n718 59.248
R1413 B.n718 B.n8 59.248
R1414 B.n712 B.n8 59.248
R1415 B.n712 B.n711 59.248
R1416 B.n711 B.n710 59.248
R1417 B.n704 B.n18 59.248
R1418 B.n704 B.n703 59.248
R1419 B.n703 B.n702 59.248
R1420 B.n702 B.n22 59.248
R1421 B.n696 B.n22 59.248
R1422 B.n696 B.n695 59.248
R1423 B.n695 B.n694 59.248
R1424 B.n694 B.n29 59.248
R1425 B.n688 B.n29 59.248
R1426 B.n687 B.n686 59.248
R1427 B.n686 B.n36 59.248
R1428 B.n680 B.n36 59.248
R1429 B.n680 B.n679 59.248
R1430 B.n679 B.n678 59.248
R1431 B.n678 B.n43 59.248
R1432 B.n672 B.n43 59.248
R1433 B.n672 B.n671 59.248
R1434 B.n671 B.n670 59.248
R1435 B.n670 B.n50 59.248
R1436 B.n664 B.n50 59.248
R1437 B.n664 B.n663 59.248
R1438 B.n662 B.n57 59.248
R1439 B.n656 B.n57 59.248
R1440 B.n656 B.n655 59.248
R1441 B.n655 B.n654 59.248
R1442 B.n654 B.n64 59.248
R1443 B.n648 B.n64 59.248
R1444 B.n648 B.n647 59.248
R1445 B.n647 B.n646 59.248
R1446 B.t5 B.n162 39.2084
R1447 B.n663 B.t12 39.2084
R1448 B.n644 B.n643 34.1859
R1449 B.n513 B.n512 34.1859
R1450 B.n353 B.n180 34.1859
R1451 B.n349 B.n348 34.1859
R1452 B.n448 B.t1 33.9807
R1453 B.n710 B.t3 33.9807
R1454 B.n417 B.t0 30.4955
R1455 B.n688 B.t2 30.4955
R1456 B.n142 B.t0 28.753
R1457 B.t2 B.n687 28.753
R1458 B.n441 B.t1 25.2678
R1459 B.n18 B.t3 25.2678
R1460 B.n375 B.t5 20.0401
R1461 B.t12 B.n662 20.0401
R1462 B B.n722 18.0485
R1463 B.n643 B.n642 10.6151
R1464 B.n642 B.n73 10.6151
R1465 B.n636 B.n73 10.6151
R1466 B.n636 B.n635 10.6151
R1467 B.n635 B.n634 10.6151
R1468 B.n634 B.n75 10.6151
R1469 B.n628 B.n75 10.6151
R1470 B.n628 B.n627 10.6151
R1471 B.n627 B.n626 10.6151
R1472 B.n626 B.n77 10.6151
R1473 B.n620 B.n77 10.6151
R1474 B.n620 B.n619 10.6151
R1475 B.n619 B.n618 10.6151
R1476 B.n618 B.n79 10.6151
R1477 B.n612 B.n79 10.6151
R1478 B.n612 B.n611 10.6151
R1479 B.n611 B.n610 10.6151
R1480 B.n610 B.n81 10.6151
R1481 B.n604 B.n81 10.6151
R1482 B.n604 B.n603 10.6151
R1483 B.n603 B.n602 10.6151
R1484 B.n602 B.n83 10.6151
R1485 B.n596 B.n83 10.6151
R1486 B.n596 B.n595 10.6151
R1487 B.n595 B.n594 10.6151
R1488 B.n594 B.n85 10.6151
R1489 B.n588 B.n85 10.6151
R1490 B.n586 B.n585 10.6151
R1491 B.n585 B.n89 10.6151
R1492 B.n579 B.n89 10.6151
R1493 B.n579 B.n578 10.6151
R1494 B.n578 B.n577 10.6151
R1495 B.n577 B.n91 10.6151
R1496 B.n571 B.n91 10.6151
R1497 B.n571 B.n570 10.6151
R1498 B.n568 B.n95 10.6151
R1499 B.n562 B.n95 10.6151
R1500 B.n562 B.n561 10.6151
R1501 B.n561 B.n560 10.6151
R1502 B.n560 B.n97 10.6151
R1503 B.n554 B.n97 10.6151
R1504 B.n554 B.n553 10.6151
R1505 B.n553 B.n552 10.6151
R1506 B.n552 B.n99 10.6151
R1507 B.n546 B.n99 10.6151
R1508 B.n546 B.n545 10.6151
R1509 B.n545 B.n544 10.6151
R1510 B.n544 B.n101 10.6151
R1511 B.n538 B.n101 10.6151
R1512 B.n538 B.n537 10.6151
R1513 B.n537 B.n536 10.6151
R1514 B.n536 B.n103 10.6151
R1515 B.n530 B.n103 10.6151
R1516 B.n530 B.n529 10.6151
R1517 B.n529 B.n528 10.6151
R1518 B.n528 B.n105 10.6151
R1519 B.n522 B.n105 10.6151
R1520 B.n522 B.n521 10.6151
R1521 B.n521 B.n520 10.6151
R1522 B.n520 B.n107 10.6151
R1523 B.n514 B.n107 10.6151
R1524 B.n514 B.n513 10.6151
R1525 B.n354 B.n353 10.6151
R1526 B.n355 B.n354 10.6151
R1527 B.n355 B.n172 10.6151
R1528 B.n365 B.n172 10.6151
R1529 B.n366 B.n365 10.6151
R1530 B.n367 B.n366 10.6151
R1531 B.n367 B.n164 10.6151
R1532 B.n377 B.n164 10.6151
R1533 B.n378 B.n377 10.6151
R1534 B.n379 B.n378 10.6151
R1535 B.n379 B.n156 10.6151
R1536 B.n389 B.n156 10.6151
R1537 B.n390 B.n389 10.6151
R1538 B.n391 B.n390 10.6151
R1539 B.n391 B.n148 10.6151
R1540 B.n401 B.n148 10.6151
R1541 B.n402 B.n401 10.6151
R1542 B.n403 B.n402 10.6151
R1543 B.n403 B.n139 10.6151
R1544 B.n413 B.n139 10.6151
R1545 B.n414 B.n413 10.6151
R1546 B.n415 B.n414 10.6151
R1547 B.n415 B.n132 10.6151
R1548 B.n425 B.n132 10.6151
R1549 B.n426 B.n425 10.6151
R1550 B.n427 B.n426 10.6151
R1551 B.n427 B.n124 10.6151
R1552 B.n437 B.n124 10.6151
R1553 B.n438 B.n437 10.6151
R1554 B.n439 B.n438 10.6151
R1555 B.n439 B.n117 10.6151
R1556 B.n450 B.n117 10.6151
R1557 B.n451 B.n450 10.6151
R1558 B.n453 B.n451 10.6151
R1559 B.n453 B.n452 10.6151
R1560 B.n452 B.n109 10.6151
R1561 B.n464 B.n109 10.6151
R1562 B.n465 B.n464 10.6151
R1563 B.n466 B.n465 10.6151
R1564 B.n467 B.n466 10.6151
R1565 B.n469 B.n467 10.6151
R1566 B.n470 B.n469 10.6151
R1567 B.n471 B.n470 10.6151
R1568 B.n472 B.n471 10.6151
R1569 B.n474 B.n472 10.6151
R1570 B.n475 B.n474 10.6151
R1571 B.n476 B.n475 10.6151
R1572 B.n477 B.n476 10.6151
R1573 B.n479 B.n477 10.6151
R1574 B.n480 B.n479 10.6151
R1575 B.n481 B.n480 10.6151
R1576 B.n482 B.n481 10.6151
R1577 B.n484 B.n482 10.6151
R1578 B.n485 B.n484 10.6151
R1579 B.n486 B.n485 10.6151
R1580 B.n487 B.n486 10.6151
R1581 B.n489 B.n487 10.6151
R1582 B.n490 B.n489 10.6151
R1583 B.n491 B.n490 10.6151
R1584 B.n492 B.n491 10.6151
R1585 B.n494 B.n492 10.6151
R1586 B.n495 B.n494 10.6151
R1587 B.n496 B.n495 10.6151
R1588 B.n497 B.n496 10.6151
R1589 B.n499 B.n497 10.6151
R1590 B.n500 B.n499 10.6151
R1591 B.n501 B.n500 10.6151
R1592 B.n502 B.n501 10.6151
R1593 B.n504 B.n502 10.6151
R1594 B.n505 B.n504 10.6151
R1595 B.n506 B.n505 10.6151
R1596 B.n507 B.n506 10.6151
R1597 B.n509 B.n507 10.6151
R1598 B.n510 B.n509 10.6151
R1599 B.n511 B.n510 10.6151
R1600 B.n512 B.n511 10.6151
R1601 B.n348 B.n347 10.6151
R1602 B.n347 B.n184 10.6151
R1603 B.n342 B.n184 10.6151
R1604 B.n342 B.n341 10.6151
R1605 B.n341 B.n186 10.6151
R1606 B.n336 B.n186 10.6151
R1607 B.n336 B.n335 10.6151
R1608 B.n335 B.n334 10.6151
R1609 B.n334 B.n188 10.6151
R1610 B.n328 B.n188 10.6151
R1611 B.n328 B.n327 10.6151
R1612 B.n327 B.n326 10.6151
R1613 B.n326 B.n190 10.6151
R1614 B.n320 B.n190 10.6151
R1615 B.n320 B.n319 10.6151
R1616 B.n319 B.n318 10.6151
R1617 B.n318 B.n192 10.6151
R1618 B.n312 B.n192 10.6151
R1619 B.n312 B.n311 10.6151
R1620 B.n311 B.n310 10.6151
R1621 B.n310 B.n194 10.6151
R1622 B.n304 B.n194 10.6151
R1623 B.n304 B.n303 10.6151
R1624 B.n303 B.n302 10.6151
R1625 B.n302 B.n196 10.6151
R1626 B.n296 B.n196 10.6151
R1627 B.n296 B.n295 10.6151
R1628 B.n293 B.n200 10.6151
R1629 B.n287 B.n200 10.6151
R1630 B.n287 B.n286 10.6151
R1631 B.n286 B.n285 10.6151
R1632 B.n285 B.n202 10.6151
R1633 B.n279 B.n202 10.6151
R1634 B.n279 B.n278 10.6151
R1635 B.n278 B.n277 10.6151
R1636 B.n273 B.n272 10.6151
R1637 B.n272 B.n208 10.6151
R1638 B.n267 B.n208 10.6151
R1639 B.n267 B.n266 10.6151
R1640 B.n266 B.n265 10.6151
R1641 B.n265 B.n210 10.6151
R1642 B.n259 B.n210 10.6151
R1643 B.n259 B.n258 10.6151
R1644 B.n258 B.n257 10.6151
R1645 B.n257 B.n212 10.6151
R1646 B.n251 B.n212 10.6151
R1647 B.n251 B.n250 10.6151
R1648 B.n250 B.n249 10.6151
R1649 B.n249 B.n214 10.6151
R1650 B.n243 B.n214 10.6151
R1651 B.n243 B.n242 10.6151
R1652 B.n242 B.n241 10.6151
R1653 B.n241 B.n216 10.6151
R1654 B.n235 B.n216 10.6151
R1655 B.n235 B.n234 10.6151
R1656 B.n234 B.n233 10.6151
R1657 B.n233 B.n218 10.6151
R1658 B.n227 B.n218 10.6151
R1659 B.n227 B.n226 10.6151
R1660 B.n226 B.n225 10.6151
R1661 B.n225 B.n220 10.6151
R1662 B.n220 B.n180 10.6151
R1663 B.n349 B.n176 10.6151
R1664 B.n359 B.n176 10.6151
R1665 B.n360 B.n359 10.6151
R1666 B.n361 B.n360 10.6151
R1667 B.n361 B.n168 10.6151
R1668 B.n371 B.n168 10.6151
R1669 B.n372 B.n371 10.6151
R1670 B.n373 B.n372 10.6151
R1671 B.n373 B.n160 10.6151
R1672 B.n383 B.n160 10.6151
R1673 B.n384 B.n383 10.6151
R1674 B.n385 B.n384 10.6151
R1675 B.n385 B.n152 10.6151
R1676 B.n395 B.n152 10.6151
R1677 B.n396 B.n395 10.6151
R1678 B.n397 B.n396 10.6151
R1679 B.n397 B.n144 10.6151
R1680 B.n407 B.n144 10.6151
R1681 B.n408 B.n407 10.6151
R1682 B.n409 B.n408 10.6151
R1683 B.n409 B.n136 10.6151
R1684 B.n419 B.n136 10.6151
R1685 B.n420 B.n419 10.6151
R1686 B.n421 B.n420 10.6151
R1687 B.n421 B.n128 10.6151
R1688 B.n431 B.n128 10.6151
R1689 B.n432 B.n431 10.6151
R1690 B.n433 B.n432 10.6151
R1691 B.n433 B.n120 10.6151
R1692 B.n444 B.n120 10.6151
R1693 B.n445 B.n444 10.6151
R1694 B.n446 B.n445 10.6151
R1695 B.n446 B.n113 10.6151
R1696 B.n457 B.n113 10.6151
R1697 B.n458 B.n457 10.6151
R1698 B.n459 B.n458 10.6151
R1699 B.n459 B.n0 10.6151
R1700 B.n716 B.n1 10.6151
R1701 B.n716 B.n715 10.6151
R1702 B.n715 B.n714 10.6151
R1703 B.n714 B.n10 10.6151
R1704 B.n708 B.n10 10.6151
R1705 B.n708 B.n707 10.6151
R1706 B.n707 B.n706 10.6151
R1707 B.n706 B.n16 10.6151
R1708 B.n700 B.n16 10.6151
R1709 B.n700 B.n699 10.6151
R1710 B.n699 B.n698 10.6151
R1711 B.n698 B.n24 10.6151
R1712 B.n692 B.n24 10.6151
R1713 B.n692 B.n691 10.6151
R1714 B.n691 B.n690 10.6151
R1715 B.n690 B.n31 10.6151
R1716 B.n684 B.n31 10.6151
R1717 B.n684 B.n683 10.6151
R1718 B.n683 B.n682 10.6151
R1719 B.n682 B.n38 10.6151
R1720 B.n676 B.n38 10.6151
R1721 B.n676 B.n675 10.6151
R1722 B.n675 B.n674 10.6151
R1723 B.n674 B.n45 10.6151
R1724 B.n668 B.n45 10.6151
R1725 B.n668 B.n667 10.6151
R1726 B.n667 B.n666 10.6151
R1727 B.n666 B.n52 10.6151
R1728 B.n660 B.n52 10.6151
R1729 B.n660 B.n659 10.6151
R1730 B.n659 B.n658 10.6151
R1731 B.n658 B.n59 10.6151
R1732 B.n652 B.n59 10.6151
R1733 B.n652 B.n651 10.6151
R1734 B.n651 B.n650 10.6151
R1735 B.n650 B.n66 10.6151
R1736 B.n644 B.n66 10.6151
R1737 B.n587 B.n586 6.5566
R1738 B.n570 B.n569 6.5566
R1739 B.n294 B.n293 6.5566
R1740 B.n277 B.n206 6.5566
R1741 B.n588 B.n587 4.05904
R1742 B.n569 B.n568 4.05904
R1743 B.n295 B.n294 4.05904
R1744 B.n273 B.n206 4.05904
R1745 B.n722 B.n0 2.81026
R1746 B.n722 B.n1 2.81026
R1747 VP.n15 VP.n14 161.3
R1748 VP.n13 VP.n1 161.3
R1749 VP.n12 VP.n11 161.3
R1750 VP.n10 VP.n2 161.3
R1751 VP.n9 VP.n8 161.3
R1752 VP.n7 VP.n3 161.3
R1753 VP.n4 VP.t1 92.5654
R1754 VP.n4 VP.t0 91.5625
R1755 VP.n6 VP.n5 68.5364
R1756 VP.n16 VP.n0 68.5364
R1757 VP.n6 VP.t3 58.0775
R1758 VP.n0 VP.t2 58.0775
R1759 VP.n12 VP.n2 56.5193
R1760 VP.n5 VP.n4 47.1663
R1761 VP.n8 VP.n7 24.4675
R1762 VP.n8 VP.n2 24.4675
R1763 VP.n13 VP.n12 24.4675
R1764 VP.n14 VP.n13 24.4675
R1765 VP.n7 VP.n6 21.5315
R1766 VP.n14 VP.n0 21.5315
R1767 VP.n5 VP.n3 0.354971
R1768 VP.n16 VP.n15 0.354971
R1769 VP VP.n16 0.26696
R1770 VP.n9 VP.n3 0.189894
R1771 VP.n10 VP.n9 0.189894
R1772 VP.n11 VP.n10 0.189894
R1773 VP.n11 VP.n1 0.189894
R1774 VP.n15 VP.n1 0.189894
R1775 VDD1 VDD1.n1 102.772
R1776 VDD1 VDD1.n0 63.5131
R1777 VDD1.n0 VDD1.t2 2.69438
R1778 VDD1.n0 VDD1.t3 2.69438
R1779 VDD1.n1 VDD1.t0 2.69438
R1780 VDD1.n1 VDD1.t1 2.69438
C0 VDD1 VP 3.38124f
C1 VDD1 VN 0.149549f
C2 VTAIL VP 3.31632f
C3 VDD1 VDD2 1.13624f
C4 VTAIL VN 3.30221f
C5 VN VP 5.65435f
C6 VTAIL VDD2 4.51827f
C7 VP VDD2 0.423082f
C8 VTAIL VDD1 4.46104f
C9 VN VDD2 3.10856f
C10 VDD2 B 3.667217f
C11 VDD1 B 7.56926f
C12 VTAIL B 7.525908f
C13 VN B 11.226151f
C14 VP B 9.592009f
C15 VDD1.t2 B 0.163885f
C16 VDD1.t3 B 0.163885f
C17 VDD1.n0 B 1.39711f
C18 VDD1.t0 B 0.163885f
C19 VDD1.t1 B 0.163885f
C20 VDD1.n1 B 1.97965f
C21 VP.t2 B 1.54079f
C22 VP.n0 B 0.667424f
C23 VP.n1 B 0.025691f
C24 VP.n2 B 0.037503f
C25 VP.n3 B 0.041464f
C26 VP.t3 B 1.54079f
C27 VP.t1 B 1.81982f
C28 VP.t0 B 1.81197f
C29 VP.n4 B 2.47455f
C30 VP.n5 B 1.3252f
C31 VP.n6 B 0.667424f
C32 VP.n7 B 0.045044f
C33 VP.n8 B 0.047881f
C34 VP.n9 B 0.025691f
C35 VP.n10 B 0.025691f
C36 VP.n11 B 0.025691f
C37 VP.n12 B 0.037503f
C38 VP.n13 B 0.047881f
C39 VP.n14 B 0.045044f
C40 VP.n15 B 0.041464f
C41 VP.n16 B 0.05201f
C42 VTAIL.n0 B 0.026195f
C43 VTAIL.n1 B 0.018726f
C44 VTAIL.n2 B 0.010063f
C45 VTAIL.n3 B 0.023784f
C46 VTAIL.n4 B 0.010655f
C47 VTAIL.n5 B 0.018726f
C48 VTAIL.n6 B 0.010063f
C49 VTAIL.n7 B 0.023784f
C50 VTAIL.n8 B 0.010655f
C51 VTAIL.n9 B 0.018726f
C52 VTAIL.n10 B 0.010063f
C53 VTAIL.n11 B 0.017838f
C54 VTAIL.n12 B 0.01405f
C55 VTAIL.t6 B 0.038756f
C56 VTAIL.n13 B 0.086282f
C57 VTAIL.n14 B 0.561718f
C58 VTAIL.n15 B 0.010063f
C59 VTAIL.n16 B 0.010655f
C60 VTAIL.n17 B 0.023784f
C61 VTAIL.n18 B 0.023784f
C62 VTAIL.n19 B 0.010655f
C63 VTAIL.n20 B 0.010063f
C64 VTAIL.n21 B 0.018726f
C65 VTAIL.n22 B 0.018726f
C66 VTAIL.n23 B 0.010063f
C67 VTAIL.n24 B 0.010655f
C68 VTAIL.n25 B 0.023784f
C69 VTAIL.n26 B 0.023784f
C70 VTAIL.n27 B 0.010655f
C71 VTAIL.n28 B 0.010063f
C72 VTAIL.n29 B 0.018726f
C73 VTAIL.n30 B 0.018726f
C74 VTAIL.n31 B 0.010063f
C75 VTAIL.n32 B 0.010655f
C76 VTAIL.n33 B 0.023784f
C77 VTAIL.n34 B 0.051266f
C78 VTAIL.n35 B 0.010655f
C79 VTAIL.n36 B 0.010063f
C80 VTAIL.n37 B 0.040982f
C81 VTAIL.n38 B 0.02859f
C82 VTAIL.n39 B 0.134466f
C83 VTAIL.n40 B 0.026195f
C84 VTAIL.n41 B 0.018726f
C85 VTAIL.n42 B 0.010063f
C86 VTAIL.n43 B 0.023784f
C87 VTAIL.n44 B 0.010655f
C88 VTAIL.n45 B 0.018726f
C89 VTAIL.n46 B 0.010063f
C90 VTAIL.n47 B 0.023784f
C91 VTAIL.n48 B 0.010655f
C92 VTAIL.n49 B 0.018726f
C93 VTAIL.n50 B 0.010063f
C94 VTAIL.n51 B 0.017838f
C95 VTAIL.n52 B 0.01405f
C96 VTAIL.t1 B 0.038756f
C97 VTAIL.n53 B 0.086282f
C98 VTAIL.n54 B 0.561718f
C99 VTAIL.n55 B 0.010063f
C100 VTAIL.n56 B 0.010655f
C101 VTAIL.n57 B 0.023784f
C102 VTAIL.n58 B 0.023784f
C103 VTAIL.n59 B 0.010655f
C104 VTAIL.n60 B 0.010063f
C105 VTAIL.n61 B 0.018726f
C106 VTAIL.n62 B 0.018726f
C107 VTAIL.n63 B 0.010063f
C108 VTAIL.n64 B 0.010655f
C109 VTAIL.n65 B 0.023784f
C110 VTAIL.n66 B 0.023784f
C111 VTAIL.n67 B 0.010655f
C112 VTAIL.n68 B 0.010063f
C113 VTAIL.n69 B 0.018726f
C114 VTAIL.n70 B 0.018726f
C115 VTAIL.n71 B 0.010063f
C116 VTAIL.n72 B 0.010655f
C117 VTAIL.n73 B 0.023784f
C118 VTAIL.n74 B 0.051266f
C119 VTAIL.n75 B 0.010655f
C120 VTAIL.n76 B 0.010063f
C121 VTAIL.n77 B 0.040982f
C122 VTAIL.n78 B 0.02859f
C123 VTAIL.n79 B 0.218863f
C124 VTAIL.n80 B 0.026195f
C125 VTAIL.n81 B 0.018726f
C126 VTAIL.n82 B 0.010063f
C127 VTAIL.n83 B 0.023784f
C128 VTAIL.n84 B 0.010655f
C129 VTAIL.n85 B 0.018726f
C130 VTAIL.n86 B 0.010063f
C131 VTAIL.n87 B 0.023784f
C132 VTAIL.n88 B 0.010655f
C133 VTAIL.n89 B 0.018726f
C134 VTAIL.n90 B 0.010063f
C135 VTAIL.n91 B 0.017838f
C136 VTAIL.n92 B 0.01405f
C137 VTAIL.t0 B 0.038756f
C138 VTAIL.n93 B 0.086282f
C139 VTAIL.n94 B 0.561718f
C140 VTAIL.n95 B 0.010063f
C141 VTAIL.n96 B 0.010655f
C142 VTAIL.n97 B 0.023784f
C143 VTAIL.n98 B 0.023784f
C144 VTAIL.n99 B 0.010655f
C145 VTAIL.n100 B 0.010063f
C146 VTAIL.n101 B 0.018726f
C147 VTAIL.n102 B 0.018726f
C148 VTAIL.n103 B 0.010063f
C149 VTAIL.n104 B 0.010655f
C150 VTAIL.n105 B 0.023784f
C151 VTAIL.n106 B 0.023784f
C152 VTAIL.n107 B 0.010655f
C153 VTAIL.n108 B 0.010063f
C154 VTAIL.n109 B 0.018726f
C155 VTAIL.n110 B 0.018726f
C156 VTAIL.n111 B 0.010063f
C157 VTAIL.n112 B 0.010655f
C158 VTAIL.n113 B 0.023784f
C159 VTAIL.n114 B 0.051266f
C160 VTAIL.n115 B 0.010655f
C161 VTAIL.n116 B 0.010063f
C162 VTAIL.n117 B 0.040982f
C163 VTAIL.n118 B 0.02859f
C164 VTAIL.n119 B 1.00303f
C165 VTAIL.n120 B 0.026195f
C166 VTAIL.n121 B 0.018726f
C167 VTAIL.n122 B 0.010063f
C168 VTAIL.n123 B 0.023784f
C169 VTAIL.n124 B 0.010655f
C170 VTAIL.n125 B 0.018726f
C171 VTAIL.n126 B 0.010063f
C172 VTAIL.n127 B 0.023784f
C173 VTAIL.n128 B 0.010655f
C174 VTAIL.n129 B 0.018726f
C175 VTAIL.n130 B 0.010063f
C176 VTAIL.n131 B 0.017838f
C177 VTAIL.n132 B 0.01405f
C178 VTAIL.t4 B 0.038756f
C179 VTAIL.n133 B 0.086282f
C180 VTAIL.n134 B 0.561718f
C181 VTAIL.n135 B 0.010063f
C182 VTAIL.n136 B 0.010655f
C183 VTAIL.n137 B 0.023784f
C184 VTAIL.n138 B 0.023784f
C185 VTAIL.n139 B 0.010655f
C186 VTAIL.n140 B 0.010063f
C187 VTAIL.n141 B 0.018726f
C188 VTAIL.n142 B 0.018726f
C189 VTAIL.n143 B 0.010063f
C190 VTAIL.n144 B 0.010655f
C191 VTAIL.n145 B 0.023784f
C192 VTAIL.n146 B 0.023784f
C193 VTAIL.n147 B 0.010655f
C194 VTAIL.n148 B 0.010063f
C195 VTAIL.n149 B 0.018726f
C196 VTAIL.n150 B 0.018726f
C197 VTAIL.n151 B 0.010063f
C198 VTAIL.n152 B 0.010655f
C199 VTAIL.n153 B 0.023784f
C200 VTAIL.n154 B 0.051266f
C201 VTAIL.n155 B 0.010655f
C202 VTAIL.n156 B 0.010063f
C203 VTAIL.n157 B 0.040982f
C204 VTAIL.n158 B 0.02859f
C205 VTAIL.n159 B 1.00303f
C206 VTAIL.n160 B 0.026195f
C207 VTAIL.n161 B 0.018726f
C208 VTAIL.n162 B 0.010063f
C209 VTAIL.n163 B 0.023784f
C210 VTAIL.n164 B 0.010655f
C211 VTAIL.n165 B 0.018726f
C212 VTAIL.n166 B 0.010063f
C213 VTAIL.n167 B 0.023784f
C214 VTAIL.n168 B 0.010655f
C215 VTAIL.n169 B 0.018726f
C216 VTAIL.n170 B 0.010063f
C217 VTAIL.n171 B 0.017838f
C218 VTAIL.n172 B 0.01405f
C219 VTAIL.t3 B 0.038756f
C220 VTAIL.n173 B 0.086282f
C221 VTAIL.n174 B 0.561718f
C222 VTAIL.n175 B 0.010063f
C223 VTAIL.n176 B 0.010655f
C224 VTAIL.n177 B 0.023784f
C225 VTAIL.n178 B 0.023784f
C226 VTAIL.n179 B 0.010655f
C227 VTAIL.n180 B 0.010063f
C228 VTAIL.n181 B 0.018726f
C229 VTAIL.n182 B 0.018726f
C230 VTAIL.n183 B 0.010063f
C231 VTAIL.n184 B 0.010655f
C232 VTAIL.n185 B 0.023784f
C233 VTAIL.n186 B 0.023784f
C234 VTAIL.n187 B 0.010655f
C235 VTAIL.n188 B 0.010063f
C236 VTAIL.n189 B 0.018726f
C237 VTAIL.n190 B 0.018726f
C238 VTAIL.n191 B 0.010063f
C239 VTAIL.n192 B 0.010655f
C240 VTAIL.n193 B 0.023784f
C241 VTAIL.n194 B 0.051266f
C242 VTAIL.n195 B 0.010655f
C243 VTAIL.n196 B 0.010063f
C244 VTAIL.n197 B 0.040982f
C245 VTAIL.n198 B 0.02859f
C246 VTAIL.n199 B 0.218863f
C247 VTAIL.n200 B 0.026195f
C248 VTAIL.n201 B 0.018726f
C249 VTAIL.n202 B 0.010063f
C250 VTAIL.n203 B 0.023784f
C251 VTAIL.n204 B 0.010655f
C252 VTAIL.n205 B 0.018726f
C253 VTAIL.n206 B 0.010063f
C254 VTAIL.n207 B 0.023784f
C255 VTAIL.n208 B 0.010655f
C256 VTAIL.n209 B 0.018726f
C257 VTAIL.n210 B 0.010063f
C258 VTAIL.n211 B 0.017838f
C259 VTAIL.n212 B 0.01405f
C260 VTAIL.t7 B 0.038756f
C261 VTAIL.n213 B 0.086282f
C262 VTAIL.n214 B 0.561718f
C263 VTAIL.n215 B 0.010063f
C264 VTAIL.n216 B 0.010655f
C265 VTAIL.n217 B 0.023784f
C266 VTAIL.n218 B 0.023784f
C267 VTAIL.n219 B 0.010655f
C268 VTAIL.n220 B 0.010063f
C269 VTAIL.n221 B 0.018726f
C270 VTAIL.n222 B 0.018726f
C271 VTAIL.n223 B 0.010063f
C272 VTAIL.n224 B 0.010655f
C273 VTAIL.n225 B 0.023784f
C274 VTAIL.n226 B 0.023784f
C275 VTAIL.n227 B 0.010655f
C276 VTAIL.n228 B 0.010063f
C277 VTAIL.n229 B 0.018726f
C278 VTAIL.n230 B 0.018726f
C279 VTAIL.n231 B 0.010063f
C280 VTAIL.n232 B 0.010655f
C281 VTAIL.n233 B 0.023784f
C282 VTAIL.n234 B 0.051266f
C283 VTAIL.n235 B 0.010655f
C284 VTAIL.n236 B 0.010063f
C285 VTAIL.n237 B 0.040982f
C286 VTAIL.n238 B 0.02859f
C287 VTAIL.n239 B 0.218863f
C288 VTAIL.n240 B 0.026195f
C289 VTAIL.n241 B 0.018726f
C290 VTAIL.n242 B 0.010063f
C291 VTAIL.n243 B 0.023784f
C292 VTAIL.n244 B 0.010655f
C293 VTAIL.n245 B 0.018726f
C294 VTAIL.n246 B 0.010063f
C295 VTAIL.n247 B 0.023784f
C296 VTAIL.n248 B 0.010655f
C297 VTAIL.n249 B 0.018726f
C298 VTAIL.n250 B 0.010063f
C299 VTAIL.n251 B 0.017838f
C300 VTAIL.n252 B 0.01405f
C301 VTAIL.t2 B 0.038756f
C302 VTAIL.n253 B 0.086282f
C303 VTAIL.n254 B 0.561718f
C304 VTAIL.n255 B 0.010063f
C305 VTAIL.n256 B 0.010655f
C306 VTAIL.n257 B 0.023784f
C307 VTAIL.n258 B 0.023784f
C308 VTAIL.n259 B 0.010655f
C309 VTAIL.n260 B 0.010063f
C310 VTAIL.n261 B 0.018726f
C311 VTAIL.n262 B 0.018726f
C312 VTAIL.n263 B 0.010063f
C313 VTAIL.n264 B 0.010655f
C314 VTAIL.n265 B 0.023784f
C315 VTAIL.n266 B 0.023784f
C316 VTAIL.n267 B 0.010655f
C317 VTAIL.n268 B 0.010063f
C318 VTAIL.n269 B 0.018726f
C319 VTAIL.n270 B 0.018726f
C320 VTAIL.n271 B 0.010063f
C321 VTAIL.n272 B 0.010655f
C322 VTAIL.n273 B 0.023784f
C323 VTAIL.n274 B 0.051266f
C324 VTAIL.n275 B 0.010655f
C325 VTAIL.n276 B 0.010063f
C326 VTAIL.n277 B 0.040982f
C327 VTAIL.n278 B 0.02859f
C328 VTAIL.n279 B 1.00303f
C329 VTAIL.n280 B 0.026195f
C330 VTAIL.n281 B 0.018726f
C331 VTAIL.n282 B 0.010063f
C332 VTAIL.n283 B 0.023784f
C333 VTAIL.n284 B 0.010655f
C334 VTAIL.n285 B 0.018726f
C335 VTAIL.n286 B 0.010063f
C336 VTAIL.n287 B 0.023784f
C337 VTAIL.n288 B 0.010655f
C338 VTAIL.n289 B 0.018726f
C339 VTAIL.n290 B 0.010063f
C340 VTAIL.n291 B 0.017838f
C341 VTAIL.n292 B 0.01405f
C342 VTAIL.t5 B 0.038756f
C343 VTAIL.n293 B 0.086282f
C344 VTAIL.n294 B 0.561718f
C345 VTAIL.n295 B 0.010063f
C346 VTAIL.n296 B 0.010655f
C347 VTAIL.n297 B 0.023784f
C348 VTAIL.n298 B 0.023784f
C349 VTAIL.n299 B 0.010655f
C350 VTAIL.n300 B 0.010063f
C351 VTAIL.n301 B 0.018726f
C352 VTAIL.n302 B 0.018726f
C353 VTAIL.n303 B 0.010063f
C354 VTAIL.n304 B 0.010655f
C355 VTAIL.n305 B 0.023784f
C356 VTAIL.n306 B 0.023784f
C357 VTAIL.n307 B 0.010655f
C358 VTAIL.n308 B 0.010063f
C359 VTAIL.n309 B 0.018726f
C360 VTAIL.n310 B 0.018726f
C361 VTAIL.n311 B 0.010063f
C362 VTAIL.n312 B 0.010655f
C363 VTAIL.n313 B 0.023784f
C364 VTAIL.n314 B 0.051266f
C365 VTAIL.n315 B 0.010655f
C366 VTAIL.n316 B 0.010063f
C367 VTAIL.n317 B 0.040982f
C368 VTAIL.n318 B 0.02859f
C369 VTAIL.n319 B 0.911612f
C370 VDD2.t0 B 0.159769f
C371 VDD2.t1 B 0.159769f
C372 VDD2.n0 B 1.90437f
C373 VDD2.t3 B 0.159769f
C374 VDD2.t2 B 0.159769f
C375 VDD2.n1 B 1.36156f
C376 VDD2.n2 B 3.43081f
C377 VN.t1 B 1.763f
C378 VN.t0 B 1.77063f
C379 VN.n0 B 1.07506f
C380 VN.t3 B 1.77063f
C381 VN.t2 B 1.763f
C382 VN.n1 B 2.41801f
.ends

