* NGSPICE file created from diff_pair_sample_1481.ext - technology: sky130A

.subckt diff_pair_sample_1481 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t6 VN.t0 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6107 pd=9.04 as=0.68145 ps=4.46 w=4.13 l=0.99
X1 VDD1.t3 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.68145 pd=4.46 as=1.6107 ps=9.04 w=4.13 l=0.99
X2 VDD1.t2 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.68145 pd=4.46 as=1.6107 ps=9.04 w=4.13 l=0.99
X3 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=1.6107 pd=9.04 as=0 ps=0 w=4.13 l=0.99
X4 VDD2.t3 VN.t1 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=0.68145 pd=4.46 as=1.6107 ps=9.04 w=4.13 l=0.99
X5 VTAIL.t4 VN.t2 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6107 pd=9.04 as=0.68145 ps=4.46 w=4.13 l=0.99
X6 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=1.6107 pd=9.04 as=0 ps=0 w=4.13 l=0.99
X7 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6107 pd=9.04 as=0 ps=0 w=4.13 l=0.99
X8 VTAIL.t7 VP.t2 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6107 pd=9.04 as=0.68145 ps=4.46 w=4.13 l=0.99
X9 VDD2.t2 VN.t3 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.68145 pd=4.46 as=1.6107 ps=9.04 w=4.13 l=0.99
X10 VTAIL.t2 VP.t3 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6107 pd=9.04 as=0.68145 ps=4.46 w=4.13 l=0.99
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6107 pd=9.04 as=0 ps=0 w=4.13 l=0.99
R0 VN.n0 VN.t0 159.07
R1 VN.n1 VN.t3 159.07
R2 VN.n1 VN.t2 158.982
R3 VN.n0 VN.t1 158.982
R4 VN VN.n1 66.9478
R5 VN VN.n0 31.2622
R6 VDD2.n2 VDD2.n0 101.249
R7 VDD2.n2 VDD2.n1 70.5607
R8 VDD2.n1 VDD2.t1 4.79469
R9 VDD2.n1 VDD2.t2 4.79469
R10 VDD2.n0 VDD2.t0 4.79469
R11 VDD2.n0 VDD2.t3 4.79469
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t7 58.6763
R14 VTAIL.n4 VTAIL.t3 58.6763
R15 VTAIL.n3 VTAIL.t4 58.6763
R16 VTAIL.n6 VTAIL.t0 58.676
R17 VTAIL.n7 VTAIL.t5 58.676
R18 VTAIL.n0 VTAIL.t6 58.676
R19 VTAIL.n1 VTAIL.t1 58.676
R20 VTAIL.n2 VTAIL.t2 58.676
R21 VTAIL.n7 VTAIL.n6 17.0652
R22 VTAIL.n3 VTAIL.n2 17.0652
R23 VTAIL.n4 VTAIL.n3 1.13843
R24 VTAIL.n6 VTAIL.n5 1.13843
R25 VTAIL.n2 VTAIL.n1 1.13843
R26 VTAIL VTAIL.n0 0.627655
R27 VTAIL VTAIL.n7 0.511276
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 B.n401 B.n400 585
R31 B.n402 B.n401 585
R32 B.n156 B.n62 585
R33 B.n155 B.n154 585
R34 B.n153 B.n152 585
R35 B.n151 B.n150 585
R36 B.n149 B.n148 585
R37 B.n147 B.n146 585
R38 B.n145 B.n144 585
R39 B.n143 B.n142 585
R40 B.n141 B.n140 585
R41 B.n139 B.n138 585
R42 B.n137 B.n136 585
R43 B.n135 B.n134 585
R44 B.n133 B.n132 585
R45 B.n131 B.n130 585
R46 B.n129 B.n128 585
R47 B.n127 B.n126 585
R48 B.n125 B.n124 585
R49 B.n123 B.n122 585
R50 B.n121 B.n120 585
R51 B.n119 B.n118 585
R52 B.n117 B.n116 585
R53 B.n115 B.n114 585
R54 B.n113 B.n112 585
R55 B.n111 B.n110 585
R56 B.n109 B.n108 585
R57 B.n107 B.n106 585
R58 B.n105 B.n104 585
R59 B.n102 B.n101 585
R60 B.n100 B.n99 585
R61 B.n98 B.n97 585
R62 B.n96 B.n95 585
R63 B.n94 B.n93 585
R64 B.n92 B.n91 585
R65 B.n90 B.n89 585
R66 B.n88 B.n87 585
R67 B.n86 B.n85 585
R68 B.n84 B.n83 585
R69 B.n82 B.n81 585
R70 B.n80 B.n79 585
R71 B.n78 B.n77 585
R72 B.n76 B.n75 585
R73 B.n74 B.n73 585
R74 B.n72 B.n71 585
R75 B.n70 B.n69 585
R76 B.n39 B.n38 585
R77 B.n405 B.n404 585
R78 B.n399 B.n63 585
R79 B.n63 B.n36 585
R80 B.n398 B.n35 585
R81 B.n409 B.n35 585
R82 B.n397 B.n34 585
R83 B.n410 B.n34 585
R84 B.n396 B.n33 585
R85 B.n411 B.n33 585
R86 B.n395 B.n394 585
R87 B.n394 B.n32 585
R88 B.n393 B.n28 585
R89 B.n417 B.n28 585
R90 B.n392 B.n27 585
R91 B.n418 B.n27 585
R92 B.n391 B.n26 585
R93 B.n419 B.n26 585
R94 B.n390 B.n389 585
R95 B.n389 B.n22 585
R96 B.n388 B.n21 585
R97 B.n425 B.n21 585
R98 B.n387 B.n20 585
R99 B.n426 B.n20 585
R100 B.n386 B.n19 585
R101 B.n427 B.n19 585
R102 B.n385 B.n384 585
R103 B.n384 B.n18 585
R104 B.n383 B.n14 585
R105 B.n433 B.n14 585
R106 B.n382 B.n13 585
R107 B.n434 B.n13 585
R108 B.n381 B.n12 585
R109 B.n435 B.n12 585
R110 B.n380 B.n379 585
R111 B.n379 B.n378 585
R112 B.n377 B.n376 585
R113 B.n377 B.n8 585
R114 B.n375 B.n7 585
R115 B.n442 B.n7 585
R116 B.n374 B.n6 585
R117 B.n443 B.n6 585
R118 B.n373 B.n5 585
R119 B.n444 B.n5 585
R120 B.n372 B.n371 585
R121 B.n371 B.n4 585
R122 B.n370 B.n157 585
R123 B.n370 B.n369 585
R124 B.n360 B.n158 585
R125 B.n159 B.n158 585
R126 B.n362 B.n361 585
R127 B.n363 B.n362 585
R128 B.n359 B.n164 585
R129 B.n164 B.n163 585
R130 B.n358 B.n357 585
R131 B.n357 B.n356 585
R132 B.n166 B.n165 585
R133 B.n349 B.n166 585
R134 B.n348 B.n347 585
R135 B.n350 B.n348 585
R136 B.n346 B.n171 585
R137 B.n171 B.n170 585
R138 B.n345 B.n344 585
R139 B.n344 B.n343 585
R140 B.n173 B.n172 585
R141 B.n174 B.n173 585
R142 B.n336 B.n335 585
R143 B.n337 B.n336 585
R144 B.n334 B.n179 585
R145 B.n179 B.n178 585
R146 B.n333 B.n332 585
R147 B.n332 B.n331 585
R148 B.n181 B.n180 585
R149 B.n324 B.n181 585
R150 B.n323 B.n322 585
R151 B.n325 B.n323 585
R152 B.n321 B.n186 585
R153 B.n186 B.n185 585
R154 B.n320 B.n319 585
R155 B.n319 B.n318 585
R156 B.n188 B.n187 585
R157 B.n189 B.n188 585
R158 B.n314 B.n313 585
R159 B.n192 B.n191 585
R160 B.n310 B.n309 585
R161 B.n311 B.n310 585
R162 B.n308 B.n215 585
R163 B.n307 B.n306 585
R164 B.n305 B.n304 585
R165 B.n303 B.n302 585
R166 B.n301 B.n300 585
R167 B.n299 B.n298 585
R168 B.n297 B.n296 585
R169 B.n295 B.n294 585
R170 B.n293 B.n292 585
R171 B.n291 B.n290 585
R172 B.n289 B.n288 585
R173 B.n287 B.n286 585
R174 B.n285 B.n284 585
R175 B.n283 B.n282 585
R176 B.n281 B.n280 585
R177 B.n279 B.n278 585
R178 B.n277 B.n276 585
R179 B.n275 B.n274 585
R180 B.n273 B.n272 585
R181 B.n271 B.n270 585
R182 B.n269 B.n268 585
R183 B.n267 B.n266 585
R184 B.n265 B.n264 585
R185 B.n263 B.n262 585
R186 B.n261 B.n260 585
R187 B.n258 B.n257 585
R188 B.n256 B.n255 585
R189 B.n254 B.n253 585
R190 B.n252 B.n251 585
R191 B.n250 B.n249 585
R192 B.n248 B.n247 585
R193 B.n246 B.n245 585
R194 B.n244 B.n243 585
R195 B.n242 B.n241 585
R196 B.n240 B.n239 585
R197 B.n238 B.n237 585
R198 B.n236 B.n235 585
R199 B.n234 B.n233 585
R200 B.n232 B.n231 585
R201 B.n230 B.n229 585
R202 B.n228 B.n227 585
R203 B.n226 B.n225 585
R204 B.n224 B.n223 585
R205 B.n222 B.n221 585
R206 B.n315 B.n190 585
R207 B.n190 B.n189 585
R208 B.n317 B.n316 585
R209 B.n318 B.n317 585
R210 B.n184 B.n183 585
R211 B.n185 B.n184 585
R212 B.n327 B.n326 585
R213 B.n326 B.n325 585
R214 B.n328 B.n182 585
R215 B.n324 B.n182 585
R216 B.n330 B.n329 585
R217 B.n331 B.n330 585
R218 B.n177 B.n176 585
R219 B.n178 B.n177 585
R220 B.n339 B.n338 585
R221 B.n338 B.n337 585
R222 B.n340 B.n175 585
R223 B.n175 B.n174 585
R224 B.n342 B.n341 585
R225 B.n343 B.n342 585
R226 B.n169 B.n168 585
R227 B.n170 B.n169 585
R228 B.n352 B.n351 585
R229 B.n351 B.n350 585
R230 B.n353 B.n167 585
R231 B.n349 B.n167 585
R232 B.n355 B.n354 585
R233 B.n356 B.n355 585
R234 B.n162 B.n161 585
R235 B.n163 B.n162 585
R236 B.n365 B.n364 585
R237 B.n364 B.n363 585
R238 B.n366 B.n160 585
R239 B.n160 B.n159 585
R240 B.n368 B.n367 585
R241 B.n369 B.n368 585
R242 B.n3 B.n0 585
R243 B.n4 B.n3 585
R244 B.n441 B.n1 585
R245 B.n442 B.n441 585
R246 B.n440 B.n439 585
R247 B.n440 B.n8 585
R248 B.n438 B.n9 585
R249 B.n378 B.n9 585
R250 B.n437 B.n436 585
R251 B.n436 B.n435 585
R252 B.n11 B.n10 585
R253 B.n434 B.n11 585
R254 B.n432 B.n431 585
R255 B.n433 B.n432 585
R256 B.n430 B.n15 585
R257 B.n18 B.n15 585
R258 B.n429 B.n428 585
R259 B.n428 B.n427 585
R260 B.n17 B.n16 585
R261 B.n426 B.n17 585
R262 B.n424 B.n423 585
R263 B.n425 B.n424 585
R264 B.n422 B.n23 585
R265 B.n23 B.n22 585
R266 B.n421 B.n420 585
R267 B.n420 B.n419 585
R268 B.n25 B.n24 585
R269 B.n418 B.n25 585
R270 B.n416 B.n415 585
R271 B.n417 B.n416 585
R272 B.n414 B.n29 585
R273 B.n32 B.n29 585
R274 B.n413 B.n412 585
R275 B.n412 B.n411 585
R276 B.n31 B.n30 585
R277 B.n410 B.n31 585
R278 B.n408 B.n407 585
R279 B.n409 B.n408 585
R280 B.n406 B.n37 585
R281 B.n37 B.n36 585
R282 B.n445 B.n444 585
R283 B.n443 B.n2 585
R284 B.n404 B.n37 502.111
R285 B.n401 B.n63 502.111
R286 B.n221 B.n188 502.111
R287 B.n313 B.n190 502.111
R288 B.n67 B.t15 303.397
R289 B.n64 B.t11 303.397
R290 B.n219 B.t4 303.397
R291 B.n216 B.t8 303.397
R292 B.n402 B.n61 256.663
R293 B.n402 B.n60 256.663
R294 B.n402 B.n59 256.663
R295 B.n402 B.n58 256.663
R296 B.n402 B.n57 256.663
R297 B.n402 B.n56 256.663
R298 B.n402 B.n55 256.663
R299 B.n402 B.n54 256.663
R300 B.n402 B.n53 256.663
R301 B.n402 B.n52 256.663
R302 B.n402 B.n51 256.663
R303 B.n402 B.n50 256.663
R304 B.n402 B.n49 256.663
R305 B.n402 B.n48 256.663
R306 B.n402 B.n47 256.663
R307 B.n402 B.n46 256.663
R308 B.n402 B.n45 256.663
R309 B.n402 B.n44 256.663
R310 B.n402 B.n43 256.663
R311 B.n402 B.n42 256.663
R312 B.n402 B.n41 256.663
R313 B.n402 B.n40 256.663
R314 B.n403 B.n402 256.663
R315 B.n312 B.n311 256.663
R316 B.n311 B.n193 256.663
R317 B.n311 B.n194 256.663
R318 B.n311 B.n195 256.663
R319 B.n311 B.n196 256.663
R320 B.n311 B.n197 256.663
R321 B.n311 B.n198 256.663
R322 B.n311 B.n199 256.663
R323 B.n311 B.n200 256.663
R324 B.n311 B.n201 256.663
R325 B.n311 B.n202 256.663
R326 B.n311 B.n203 256.663
R327 B.n311 B.n204 256.663
R328 B.n311 B.n205 256.663
R329 B.n311 B.n206 256.663
R330 B.n311 B.n207 256.663
R331 B.n311 B.n208 256.663
R332 B.n311 B.n209 256.663
R333 B.n311 B.n210 256.663
R334 B.n311 B.n211 256.663
R335 B.n311 B.n212 256.663
R336 B.n311 B.n213 256.663
R337 B.n311 B.n214 256.663
R338 B.n447 B.n446 256.663
R339 B.n311 B.n189 164.912
R340 B.n402 B.n36 164.912
R341 B.n69 B.n39 163.367
R342 B.n73 B.n72 163.367
R343 B.n77 B.n76 163.367
R344 B.n81 B.n80 163.367
R345 B.n85 B.n84 163.367
R346 B.n89 B.n88 163.367
R347 B.n93 B.n92 163.367
R348 B.n97 B.n96 163.367
R349 B.n101 B.n100 163.367
R350 B.n106 B.n105 163.367
R351 B.n110 B.n109 163.367
R352 B.n114 B.n113 163.367
R353 B.n118 B.n117 163.367
R354 B.n122 B.n121 163.367
R355 B.n126 B.n125 163.367
R356 B.n130 B.n129 163.367
R357 B.n134 B.n133 163.367
R358 B.n138 B.n137 163.367
R359 B.n142 B.n141 163.367
R360 B.n146 B.n145 163.367
R361 B.n150 B.n149 163.367
R362 B.n154 B.n153 163.367
R363 B.n401 B.n62 163.367
R364 B.n319 B.n188 163.367
R365 B.n319 B.n186 163.367
R366 B.n323 B.n186 163.367
R367 B.n323 B.n181 163.367
R368 B.n332 B.n181 163.367
R369 B.n332 B.n179 163.367
R370 B.n336 B.n179 163.367
R371 B.n336 B.n173 163.367
R372 B.n344 B.n173 163.367
R373 B.n344 B.n171 163.367
R374 B.n348 B.n171 163.367
R375 B.n348 B.n166 163.367
R376 B.n357 B.n166 163.367
R377 B.n357 B.n164 163.367
R378 B.n362 B.n164 163.367
R379 B.n362 B.n158 163.367
R380 B.n370 B.n158 163.367
R381 B.n371 B.n370 163.367
R382 B.n371 B.n5 163.367
R383 B.n6 B.n5 163.367
R384 B.n7 B.n6 163.367
R385 B.n377 B.n7 163.367
R386 B.n379 B.n377 163.367
R387 B.n379 B.n12 163.367
R388 B.n13 B.n12 163.367
R389 B.n14 B.n13 163.367
R390 B.n384 B.n14 163.367
R391 B.n384 B.n19 163.367
R392 B.n20 B.n19 163.367
R393 B.n21 B.n20 163.367
R394 B.n389 B.n21 163.367
R395 B.n389 B.n26 163.367
R396 B.n27 B.n26 163.367
R397 B.n28 B.n27 163.367
R398 B.n394 B.n28 163.367
R399 B.n394 B.n33 163.367
R400 B.n34 B.n33 163.367
R401 B.n35 B.n34 163.367
R402 B.n63 B.n35 163.367
R403 B.n310 B.n192 163.367
R404 B.n310 B.n215 163.367
R405 B.n306 B.n305 163.367
R406 B.n302 B.n301 163.367
R407 B.n298 B.n297 163.367
R408 B.n294 B.n293 163.367
R409 B.n290 B.n289 163.367
R410 B.n286 B.n285 163.367
R411 B.n282 B.n281 163.367
R412 B.n278 B.n277 163.367
R413 B.n274 B.n273 163.367
R414 B.n270 B.n269 163.367
R415 B.n266 B.n265 163.367
R416 B.n262 B.n261 163.367
R417 B.n257 B.n256 163.367
R418 B.n253 B.n252 163.367
R419 B.n249 B.n248 163.367
R420 B.n245 B.n244 163.367
R421 B.n241 B.n240 163.367
R422 B.n237 B.n236 163.367
R423 B.n233 B.n232 163.367
R424 B.n229 B.n228 163.367
R425 B.n225 B.n224 163.367
R426 B.n317 B.n190 163.367
R427 B.n317 B.n184 163.367
R428 B.n326 B.n184 163.367
R429 B.n326 B.n182 163.367
R430 B.n330 B.n182 163.367
R431 B.n330 B.n177 163.367
R432 B.n338 B.n177 163.367
R433 B.n338 B.n175 163.367
R434 B.n342 B.n175 163.367
R435 B.n342 B.n169 163.367
R436 B.n351 B.n169 163.367
R437 B.n351 B.n167 163.367
R438 B.n355 B.n167 163.367
R439 B.n355 B.n162 163.367
R440 B.n364 B.n162 163.367
R441 B.n364 B.n160 163.367
R442 B.n368 B.n160 163.367
R443 B.n368 B.n3 163.367
R444 B.n445 B.n3 163.367
R445 B.n441 B.n2 163.367
R446 B.n441 B.n440 163.367
R447 B.n440 B.n9 163.367
R448 B.n436 B.n9 163.367
R449 B.n436 B.n11 163.367
R450 B.n432 B.n11 163.367
R451 B.n432 B.n15 163.367
R452 B.n428 B.n15 163.367
R453 B.n428 B.n17 163.367
R454 B.n424 B.n17 163.367
R455 B.n424 B.n23 163.367
R456 B.n420 B.n23 163.367
R457 B.n420 B.n25 163.367
R458 B.n416 B.n25 163.367
R459 B.n416 B.n29 163.367
R460 B.n412 B.n29 163.367
R461 B.n412 B.n31 163.367
R462 B.n408 B.n31 163.367
R463 B.n408 B.n37 163.367
R464 B.n64 B.t13 97.7784
R465 B.n219 B.t7 97.7784
R466 B.n67 B.t16 97.7745
R467 B.n216 B.t10 97.7745
R468 B.n318 B.n189 79.5327
R469 B.n318 B.n185 79.5327
R470 B.n325 B.n185 79.5327
R471 B.n325 B.n324 79.5327
R472 B.n331 B.n178 79.5327
R473 B.n337 B.n178 79.5327
R474 B.n337 B.n174 79.5327
R475 B.n343 B.n174 79.5327
R476 B.n343 B.n170 79.5327
R477 B.n350 B.n170 79.5327
R478 B.n350 B.n349 79.5327
R479 B.n356 B.n163 79.5327
R480 B.n363 B.n163 79.5327
R481 B.n369 B.n159 79.5327
R482 B.n369 B.n4 79.5327
R483 B.n444 B.n4 79.5327
R484 B.n444 B.n443 79.5327
R485 B.n443 B.n442 79.5327
R486 B.n442 B.n8 79.5327
R487 B.n378 B.n8 79.5327
R488 B.n435 B.n434 79.5327
R489 B.n434 B.n433 79.5327
R490 B.n427 B.n18 79.5327
R491 B.n427 B.n426 79.5327
R492 B.n426 B.n425 79.5327
R493 B.n425 B.n22 79.5327
R494 B.n419 B.n22 79.5327
R495 B.n419 B.n418 79.5327
R496 B.n418 B.n417 79.5327
R497 B.n411 B.n32 79.5327
R498 B.n411 B.n410 79.5327
R499 B.n410 B.n409 79.5327
R500 B.n409 B.n36 79.5327
R501 B.n324 B.t5 78.3631
R502 B.n32 B.t12 78.3631
R503 B.n363 B.t1 76.0239
R504 B.n435 B.t3 76.0239
R505 B.n356 B.t2 73.6847
R506 B.n433 B.t0 73.6847
R507 B.n65 B.t14 72.1784
R508 B.n220 B.t6 72.1784
R509 B.n68 B.t17 72.1745
R510 B.n217 B.t9 72.1745
R511 B.n404 B.n403 71.676
R512 B.n69 B.n40 71.676
R513 B.n73 B.n41 71.676
R514 B.n77 B.n42 71.676
R515 B.n81 B.n43 71.676
R516 B.n85 B.n44 71.676
R517 B.n89 B.n45 71.676
R518 B.n93 B.n46 71.676
R519 B.n97 B.n47 71.676
R520 B.n101 B.n48 71.676
R521 B.n106 B.n49 71.676
R522 B.n110 B.n50 71.676
R523 B.n114 B.n51 71.676
R524 B.n118 B.n52 71.676
R525 B.n122 B.n53 71.676
R526 B.n126 B.n54 71.676
R527 B.n130 B.n55 71.676
R528 B.n134 B.n56 71.676
R529 B.n138 B.n57 71.676
R530 B.n142 B.n58 71.676
R531 B.n146 B.n59 71.676
R532 B.n150 B.n60 71.676
R533 B.n154 B.n61 71.676
R534 B.n62 B.n61 71.676
R535 B.n153 B.n60 71.676
R536 B.n149 B.n59 71.676
R537 B.n145 B.n58 71.676
R538 B.n141 B.n57 71.676
R539 B.n137 B.n56 71.676
R540 B.n133 B.n55 71.676
R541 B.n129 B.n54 71.676
R542 B.n125 B.n53 71.676
R543 B.n121 B.n52 71.676
R544 B.n117 B.n51 71.676
R545 B.n113 B.n50 71.676
R546 B.n109 B.n49 71.676
R547 B.n105 B.n48 71.676
R548 B.n100 B.n47 71.676
R549 B.n96 B.n46 71.676
R550 B.n92 B.n45 71.676
R551 B.n88 B.n44 71.676
R552 B.n84 B.n43 71.676
R553 B.n80 B.n42 71.676
R554 B.n76 B.n41 71.676
R555 B.n72 B.n40 71.676
R556 B.n403 B.n39 71.676
R557 B.n313 B.n312 71.676
R558 B.n215 B.n193 71.676
R559 B.n305 B.n194 71.676
R560 B.n301 B.n195 71.676
R561 B.n297 B.n196 71.676
R562 B.n293 B.n197 71.676
R563 B.n289 B.n198 71.676
R564 B.n285 B.n199 71.676
R565 B.n281 B.n200 71.676
R566 B.n277 B.n201 71.676
R567 B.n273 B.n202 71.676
R568 B.n269 B.n203 71.676
R569 B.n265 B.n204 71.676
R570 B.n261 B.n205 71.676
R571 B.n256 B.n206 71.676
R572 B.n252 B.n207 71.676
R573 B.n248 B.n208 71.676
R574 B.n244 B.n209 71.676
R575 B.n240 B.n210 71.676
R576 B.n236 B.n211 71.676
R577 B.n232 B.n212 71.676
R578 B.n228 B.n213 71.676
R579 B.n224 B.n214 71.676
R580 B.n312 B.n192 71.676
R581 B.n306 B.n193 71.676
R582 B.n302 B.n194 71.676
R583 B.n298 B.n195 71.676
R584 B.n294 B.n196 71.676
R585 B.n290 B.n197 71.676
R586 B.n286 B.n198 71.676
R587 B.n282 B.n199 71.676
R588 B.n278 B.n200 71.676
R589 B.n274 B.n201 71.676
R590 B.n270 B.n202 71.676
R591 B.n266 B.n203 71.676
R592 B.n262 B.n204 71.676
R593 B.n257 B.n205 71.676
R594 B.n253 B.n206 71.676
R595 B.n249 B.n207 71.676
R596 B.n245 B.n208 71.676
R597 B.n241 B.n209 71.676
R598 B.n237 B.n210 71.676
R599 B.n233 B.n211 71.676
R600 B.n229 B.n212 71.676
R601 B.n225 B.n213 71.676
R602 B.n221 B.n214 71.676
R603 B.n446 B.n445 71.676
R604 B.n446 B.n2 71.676
R605 B.n103 B.n68 59.5399
R606 B.n66 B.n65 59.5399
R607 B.n259 B.n220 59.5399
R608 B.n218 B.n217 59.5399
R609 B.n315 B.n314 32.6249
R610 B.n222 B.n187 32.6249
R611 B.n400 B.n399 32.6249
R612 B.n406 B.n405 32.6249
R613 B.n68 B.n67 25.6005
R614 B.n65 B.n64 25.6005
R615 B.n220 B.n219 25.6005
R616 B.n217 B.n216 25.6005
R617 B B.n447 18.0485
R618 B.n316 B.n315 10.6151
R619 B.n316 B.n183 10.6151
R620 B.n327 B.n183 10.6151
R621 B.n328 B.n327 10.6151
R622 B.n329 B.n328 10.6151
R623 B.n329 B.n176 10.6151
R624 B.n339 B.n176 10.6151
R625 B.n340 B.n339 10.6151
R626 B.n341 B.n340 10.6151
R627 B.n341 B.n168 10.6151
R628 B.n352 B.n168 10.6151
R629 B.n353 B.n352 10.6151
R630 B.n354 B.n353 10.6151
R631 B.n354 B.n161 10.6151
R632 B.n365 B.n161 10.6151
R633 B.n366 B.n365 10.6151
R634 B.n367 B.n366 10.6151
R635 B.n367 B.n0 10.6151
R636 B.n314 B.n191 10.6151
R637 B.n309 B.n191 10.6151
R638 B.n309 B.n308 10.6151
R639 B.n308 B.n307 10.6151
R640 B.n307 B.n304 10.6151
R641 B.n304 B.n303 10.6151
R642 B.n303 B.n300 10.6151
R643 B.n300 B.n299 10.6151
R644 B.n299 B.n296 10.6151
R645 B.n296 B.n295 10.6151
R646 B.n295 B.n292 10.6151
R647 B.n292 B.n291 10.6151
R648 B.n291 B.n288 10.6151
R649 B.n288 B.n287 10.6151
R650 B.n287 B.n284 10.6151
R651 B.n284 B.n283 10.6151
R652 B.n283 B.n280 10.6151
R653 B.n280 B.n279 10.6151
R654 B.n276 B.n275 10.6151
R655 B.n275 B.n272 10.6151
R656 B.n272 B.n271 10.6151
R657 B.n271 B.n268 10.6151
R658 B.n268 B.n267 10.6151
R659 B.n267 B.n264 10.6151
R660 B.n264 B.n263 10.6151
R661 B.n263 B.n260 10.6151
R662 B.n258 B.n255 10.6151
R663 B.n255 B.n254 10.6151
R664 B.n254 B.n251 10.6151
R665 B.n251 B.n250 10.6151
R666 B.n250 B.n247 10.6151
R667 B.n247 B.n246 10.6151
R668 B.n246 B.n243 10.6151
R669 B.n243 B.n242 10.6151
R670 B.n242 B.n239 10.6151
R671 B.n239 B.n238 10.6151
R672 B.n238 B.n235 10.6151
R673 B.n235 B.n234 10.6151
R674 B.n234 B.n231 10.6151
R675 B.n231 B.n230 10.6151
R676 B.n230 B.n227 10.6151
R677 B.n227 B.n226 10.6151
R678 B.n226 B.n223 10.6151
R679 B.n223 B.n222 10.6151
R680 B.n320 B.n187 10.6151
R681 B.n321 B.n320 10.6151
R682 B.n322 B.n321 10.6151
R683 B.n322 B.n180 10.6151
R684 B.n333 B.n180 10.6151
R685 B.n334 B.n333 10.6151
R686 B.n335 B.n334 10.6151
R687 B.n335 B.n172 10.6151
R688 B.n345 B.n172 10.6151
R689 B.n346 B.n345 10.6151
R690 B.n347 B.n346 10.6151
R691 B.n347 B.n165 10.6151
R692 B.n358 B.n165 10.6151
R693 B.n359 B.n358 10.6151
R694 B.n361 B.n359 10.6151
R695 B.n361 B.n360 10.6151
R696 B.n360 B.n157 10.6151
R697 B.n372 B.n157 10.6151
R698 B.n373 B.n372 10.6151
R699 B.n374 B.n373 10.6151
R700 B.n375 B.n374 10.6151
R701 B.n376 B.n375 10.6151
R702 B.n380 B.n376 10.6151
R703 B.n381 B.n380 10.6151
R704 B.n382 B.n381 10.6151
R705 B.n383 B.n382 10.6151
R706 B.n385 B.n383 10.6151
R707 B.n386 B.n385 10.6151
R708 B.n387 B.n386 10.6151
R709 B.n388 B.n387 10.6151
R710 B.n390 B.n388 10.6151
R711 B.n391 B.n390 10.6151
R712 B.n392 B.n391 10.6151
R713 B.n393 B.n392 10.6151
R714 B.n395 B.n393 10.6151
R715 B.n396 B.n395 10.6151
R716 B.n397 B.n396 10.6151
R717 B.n398 B.n397 10.6151
R718 B.n399 B.n398 10.6151
R719 B.n439 B.n1 10.6151
R720 B.n439 B.n438 10.6151
R721 B.n438 B.n437 10.6151
R722 B.n437 B.n10 10.6151
R723 B.n431 B.n10 10.6151
R724 B.n431 B.n430 10.6151
R725 B.n430 B.n429 10.6151
R726 B.n429 B.n16 10.6151
R727 B.n423 B.n16 10.6151
R728 B.n423 B.n422 10.6151
R729 B.n422 B.n421 10.6151
R730 B.n421 B.n24 10.6151
R731 B.n415 B.n24 10.6151
R732 B.n415 B.n414 10.6151
R733 B.n414 B.n413 10.6151
R734 B.n413 B.n30 10.6151
R735 B.n407 B.n30 10.6151
R736 B.n407 B.n406 10.6151
R737 B.n405 B.n38 10.6151
R738 B.n70 B.n38 10.6151
R739 B.n71 B.n70 10.6151
R740 B.n74 B.n71 10.6151
R741 B.n75 B.n74 10.6151
R742 B.n78 B.n75 10.6151
R743 B.n79 B.n78 10.6151
R744 B.n82 B.n79 10.6151
R745 B.n83 B.n82 10.6151
R746 B.n86 B.n83 10.6151
R747 B.n87 B.n86 10.6151
R748 B.n90 B.n87 10.6151
R749 B.n91 B.n90 10.6151
R750 B.n94 B.n91 10.6151
R751 B.n95 B.n94 10.6151
R752 B.n98 B.n95 10.6151
R753 B.n99 B.n98 10.6151
R754 B.n102 B.n99 10.6151
R755 B.n107 B.n104 10.6151
R756 B.n108 B.n107 10.6151
R757 B.n111 B.n108 10.6151
R758 B.n112 B.n111 10.6151
R759 B.n115 B.n112 10.6151
R760 B.n116 B.n115 10.6151
R761 B.n119 B.n116 10.6151
R762 B.n120 B.n119 10.6151
R763 B.n124 B.n123 10.6151
R764 B.n127 B.n124 10.6151
R765 B.n128 B.n127 10.6151
R766 B.n131 B.n128 10.6151
R767 B.n132 B.n131 10.6151
R768 B.n135 B.n132 10.6151
R769 B.n136 B.n135 10.6151
R770 B.n139 B.n136 10.6151
R771 B.n140 B.n139 10.6151
R772 B.n143 B.n140 10.6151
R773 B.n144 B.n143 10.6151
R774 B.n147 B.n144 10.6151
R775 B.n148 B.n147 10.6151
R776 B.n151 B.n148 10.6151
R777 B.n152 B.n151 10.6151
R778 B.n155 B.n152 10.6151
R779 B.n156 B.n155 10.6151
R780 B.n400 B.n156 10.6151
R781 B.n447 B.n0 8.11757
R782 B.n447 B.n1 8.11757
R783 B.n276 B.n218 6.5566
R784 B.n260 B.n259 6.5566
R785 B.n104 B.n103 6.5566
R786 B.n120 B.n66 6.5566
R787 B.n349 B.t2 5.84845
R788 B.n18 B.t0 5.84845
R789 B.n279 B.n218 4.05904
R790 B.n259 B.n258 4.05904
R791 B.n103 B.n102 4.05904
R792 B.n123 B.n66 4.05904
R793 B.t1 B.n159 3.50927
R794 B.n378 B.t3 3.50927
R795 B.n331 B.t5 1.17009
R796 B.n417 B.t12 1.17009
R797 VP.n0 VP.t2 159.07
R798 VP.n0 VP.t1 158.982
R799 VP.n2 VP.t3 140.463
R800 VP.n3 VP.t0 140.463
R801 VP.n4 VP.n3 80.6037
R802 VP.n2 VP.n1 80.6037
R803 VP.n1 VP.n0 66.6623
R804 VP.n3 VP.n2 48.2005
R805 VP.n4 VP.n1 0.380177
R806 VP VP.n4 0.146778
R807 VDD1 VDD1.n1 101.775
R808 VDD1 VDD1.n0 70.6189
R809 VDD1.n0 VDD1.t1 4.79469
R810 VDD1.n0 VDD1.t2 4.79469
R811 VDD1.n1 VDD1.t0 4.79469
R812 VDD1.n1 VDD1.t3 4.79469
C0 VN VP 3.57991f
C1 VP VTAIL 1.51655f
C2 VDD2 VP 0.296508f
C3 VN VDD1 0.151841f
C4 VDD1 VTAIL 3.15625f
C5 VDD2 VDD1 0.636212f
C6 VN VTAIL 1.50245f
C7 VDD2 VN 1.44595f
C8 VDD2 VTAIL 3.19967f
C9 VDD1 VP 1.58992f
C10 VDD2 B 2.210995f
C11 VDD1 B 4.1125f
C12 VTAIL B 4.32142f
C13 VN B 6.26268f
C14 VP B 4.868329f
C15 VDD1.t1 B 0.059719f
C16 VDD1.t2 B 0.059719f
C17 VDD1.n0 B 0.472575f
C18 VDD1.t0 B 0.059719f
C19 VDD1.t3 B 0.059719f
C20 VDD1.n1 B 0.703919f
C21 VP.t1 B 0.325743f
C22 VP.t2 B 0.32585f
C23 VP.n0 B 0.735921f
C24 VP.n1 B 1.22585f
C25 VP.t3 B 0.307332f
C26 VP.n2 B 0.158047f
C27 VP.t0 B 0.307332f
C28 VP.n3 B 0.158047f
C29 VP.n4 B 0.032413f
C30 VTAIL.t6 B 0.400355f
C31 VTAIL.n0 B 0.196055f
C32 VTAIL.t1 B 0.400355f
C33 VTAIL.n1 B 0.218026f
C34 VTAIL.t2 B 0.400355f
C35 VTAIL.n2 B 0.581263f
C36 VTAIL.t4 B 0.400357f
C37 VTAIL.n3 B 0.581261f
C38 VTAIL.t3 B 0.400357f
C39 VTAIL.n4 B 0.218025f
C40 VTAIL.t7 B 0.400357f
C41 VTAIL.n5 B 0.218025f
C42 VTAIL.t0 B 0.400355f
C43 VTAIL.n6 B 0.581263f
C44 VTAIL.t5 B 0.400355f
C45 VTAIL.n7 B 0.554285f
C46 VDD2.t0 B 0.061008f
C47 VDD2.t3 B 0.061008f
C48 VDD2.n0 B 0.70469f
C49 VDD2.t1 B 0.061008f
C50 VDD2.t2 B 0.061008f
C51 VDD2.n1 B 0.482586f
C52 VDD2.n2 B 1.69613f
C53 VN.t0 B 0.322637f
C54 VN.t1 B 0.32253f
C55 VN.n0 B 0.277079f
C56 VN.t3 B 0.322637f
C57 VN.t2 B 0.32253f
C58 VN.n1 B 0.738178f
.ends

