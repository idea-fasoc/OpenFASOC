* NGSPICE file created from diff_pair_sample_1503.ext - technology: sky130A

.subckt diff_pair_sample_1503 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9141 pd=5.87 as=2.1606 ps=11.86 w=5.54 l=0.22
X1 VDD1.t3 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9141 pd=5.87 as=2.1606 ps=11.86 w=5.54 l=0.22
X2 VTAIL.t7 VN.t1 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.1606 pd=11.86 as=0.9141 ps=5.87 w=5.54 l=0.22
X3 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=2.1606 pd=11.86 as=0 ps=0 w=5.54 l=0.22
X4 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=2.1606 pd=11.86 as=0 ps=0 w=5.54 l=0.22
X5 VTAIL.t6 VN.t2 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1606 pd=11.86 as=0.9141 ps=5.87 w=5.54 l=0.22
X6 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.1606 pd=11.86 as=0 ps=0 w=5.54 l=0.22
X7 VTAIL.t3 VP.t1 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.1606 pd=11.86 as=0.9141 ps=5.87 w=5.54 l=0.22
X8 VTAIL.t2 VP.t2 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1606 pd=11.86 as=0.9141 ps=5.87 w=5.54 l=0.22
X9 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.1606 pd=11.86 as=0 ps=0 w=5.54 l=0.22
X10 VDD2.t0 VN.t3 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9141 pd=5.87 as=2.1606 ps=11.86 w=5.54 l=0.22
X11 VDD1.t0 VP.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9141 pd=5.87 as=2.1606 ps=11.86 w=5.54 l=0.22
R0 VN.n0 VN.t3 789.458
R1 VN.n0 VN.t1 789.458
R2 VN.n1 VN.t2 789.458
R3 VN.n1 VN.t0 789.458
R4 VN VN.n1 195.773
R5 VN VN.n0 161.351
R6 VTAIL.n5 VTAIL.t3 52.8258
R7 VTAIL.n4 VTAIL.t5 52.8258
R8 VTAIL.n3 VTAIL.t6 52.8258
R9 VTAIL.n7 VTAIL.t4 52.8256
R10 VTAIL.n0 VTAIL.t7 52.8256
R11 VTAIL.n1 VTAIL.t1 52.8256
R12 VTAIL.n2 VTAIL.t2 52.8256
R13 VTAIL.n6 VTAIL.t0 52.8256
R14 VTAIL.n7 VTAIL.n6 17.6341
R15 VTAIL.n3 VTAIL.n2 17.6341
R16 VTAIL.n4 VTAIL.n3 0.474638
R17 VTAIL.n6 VTAIL.n5 0.474638
R18 VTAIL.n2 VTAIL.n1 0.474638
R19 VTAIL.n5 VTAIL.n4 0.470328
R20 VTAIL.n1 VTAIL.n0 0.470328
R21 VTAIL VTAIL.n0 0.295759
R22 VTAIL VTAIL.n7 0.179379
R23 VDD2.n2 VDD2.n0 95.8607
R24 VDD2.n2 VDD2.n1 65.9305
R25 VDD2.n1 VDD2.t1 3.57451
R26 VDD2.n1 VDD2.t3 3.57451
R27 VDD2.n0 VDD2.t2 3.57451
R28 VDD2.n0 VDD2.t0 3.57451
R29 VDD2 VDD2.n2 0.0586897
R30 B.n224 B.t15 837.755
R31 B.n221 B.t8 837.755
R32 B.n59 B.t12 837.755
R33 B.n56 B.t4 837.755
R34 B.n393 B.n392 585
R35 B.n394 B.n393 585
R36 B.n168 B.n55 585
R37 B.n167 B.n166 585
R38 B.n165 B.n164 585
R39 B.n163 B.n162 585
R40 B.n161 B.n160 585
R41 B.n159 B.n158 585
R42 B.n157 B.n156 585
R43 B.n155 B.n154 585
R44 B.n153 B.n152 585
R45 B.n151 B.n150 585
R46 B.n149 B.n148 585
R47 B.n147 B.n146 585
R48 B.n145 B.n144 585
R49 B.n143 B.n142 585
R50 B.n141 B.n140 585
R51 B.n139 B.n138 585
R52 B.n137 B.n136 585
R53 B.n135 B.n134 585
R54 B.n133 B.n132 585
R55 B.n131 B.n130 585
R56 B.n129 B.n128 585
R57 B.n127 B.n126 585
R58 B.n125 B.n124 585
R59 B.n123 B.n122 585
R60 B.n121 B.n120 585
R61 B.n119 B.n118 585
R62 B.n117 B.n116 585
R63 B.n115 B.n114 585
R64 B.n113 B.n112 585
R65 B.n111 B.n110 585
R66 B.n109 B.n108 585
R67 B.n106 B.n105 585
R68 B.n104 B.n103 585
R69 B.n102 B.n101 585
R70 B.n100 B.n99 585
R71 B.n98 B.n97 585
R72 B.n96 B.n95 585
R73 B.n94 B.n93 585
R74 B.n92 B.n91 585
R75 B.n90 B.n89 585
R76 B.n88 B.n87 585
R77 B.n86 B.n85 585
R78 B.n84 B.n83 585
R79 B.n82 B.n81 585
R80 B.n80 B.n79 585
R81 B.n78 B.n77 585
R82 B.n76 B.n75 585
R83 B.n74 B.n73 585
R84 B.n72 B.n71 585
R85 B.n70 B.n69 585
R86 B.n68 B.n67 585
R87 B.n66 B.n65 585
R88 B.n64 B.n63 585
R89 B.n62 B.n61 585
R90 B.n391 B.n27 585
R91 B.n395 B.n27 585
R92 B.n390 B.n26 585
R93 B.n396 B.n26 585
R94 B.n389 B.n388 585
R95 B.n388 B.n22 585
R96 B.n387 B.n21 585
R97 B.n402 B.n21 585
R98 B.n386 B.n20 585
R99 B.n403 B.n20 585
R100 B.n385 B.n19 585
R101 B.n404 B.n19 585
R102 B.n384 B.n383 585
R103 B.n383 B.n15 585
R104 B.n382 B.n14 585
R105 B.n410 B.n14 585
R106 B.n381 B.n13 585
R107 B.n411 B.n13 585
R108 B.n380 B.n12 585
R109 B.n412 B.n12 585
R110 B.n379 B.n378 585
R111 B.n378 B.n11 585
R112 B.n377 B.n7 585
R113 B.n418 B.n7 585
R114 B.n376 B.n6 585
R115 B.n419 B.n6 585
R116 B.n375 B.n5 585
R117 B.n420 B.n5 585
R118 B.n374 B.n373 585
R119 B.n373 B.n4 585
R120 B.n372 B.n169 585
R121 B.n372 B.n371 585
R122 B.n361 B.n170 585
R123 B.n364 B.n170 585
R124 B.n363 B.n362 585
R125 B.n365 B.n363 585
R126 B.n360 B.n174 585
R127 B.n178 B.n174 585
R128 B.n359 B.n358 585
R129 B.n358 B.n357 585
R130 B.n176 B.n175 585
R131 B.n177 B.n176 585
R132 B.n350 B.n349 585
R133 B.n351 B.n350 585
R134 B.n348 B.n182 585
R135 B.n186 B.n182 585
R136 B.n347 B.n346 585
R137 B.n346 B.n345 585
R138 B.n184 B.n183 585
R139 B.n185 B.n184 585
R140 B.n338 B.n337 585
R141 B.n339 B.n338 585
R142 B.n336 B.n191 585
R143 B.n191 B.n190 585
R144 B.n330 B.n329 585
R145 B.n328 B.n220 585
R146 B.n327 B.n219 585
R147 B.n332 B.n219 585
R148 B.n326 B.n325 585
R149 B.n324 B.n323 585
R150 B.n322 B.n321 585
R151 B.n320 B.n319 585
R152 B.n318 B.n317 585
R153 B.n316 B.n315 585
R154 B.n314 B.n313 585
R155 B.n312 B.n311 585
R156 B.n310 B.n309 585
R157 B.n308 B.n307 585
R158 B.n306 B.n305 585
R159 B.n304 B.n303 585
R160 B.n302 B.n301 585
R161 B.n300 B.n299 585
R162 B.n298 B.n297 585
R163 B.n296 B.n295 585
R164 B.n294 B.n293 585
R165 B.n292 B.n291 585
R166 B.n290 B.n289 585
R167 B.n288 B.n287 585
R168 B.n286 B.n285 585
R169 B.n284 B.n283 585
R170 B.n282 B.n281 585
R171 B.n280 B.n279 585
R172 B.n278 B.n277 585
R173 B.n276 B.n275 585
R174 B.n274 B.n273 585
R175 B.n272 B.n271 585
R176 B.n270 B.n269 585
R177 B.n267 B.n266 585
R178 B.n265 B.n264 585
R179 B.n263 B.n262 585
R180 B.n261 B.n260 585
R181 B.n259 B.n258 585
R182 B.n257 B.n256 585
R183 B.n255 B.n254 585
R184 B.n253 B.n252 585
R185 B.n251 B.n250 585
R186 B.n249 B.n248 585
R187 B.n247 B.n246 585
R188 B.n245 B.n244 585
R189 B.n243 B.n242 585
R190 B.n241 B.n240 585
R191 B.n239 B.n238 585
R192 B.n237 B.n236 585
R193 B.n235 B.n234 585
R194 B.n233 B.n232 585
R195 B.n231 B.n230 585
R196 B.n229 B.n228 585
R197 B.n227 B.n226 585
R198 B.n193 B.n192 585
R199 B.n335 B.n334 585
R200 B.n189 B.n188 585
R201 B.n190 B.n189 585
R202 B.n341 B.n340 585
R203 B.n340 B.n339 585
R204 B.n342 B.n187 585
R205 B.n187 B.n185 585
R206 B.n344 B.n343 585
R207 B.n345 B.n344 585
R208 B.n181 B.n180 585
R209 B.n186 B.n181 585
R210 B.n353 B.n352 585
R211 B.n352 B.n351 585
R212 B.n354 B.n179 585
R213 B.n179 B.n177 585
R214 B.n356 B.n355 585
R215 B.n357 B.n356 585
R216 B.n173 B.n172 585
R217 B.n178 B.n173 585
R218 B.n367 B.n366 585
R219 B.n366 B.n365 585
R220 B.n368 B.n171 585
R221 B.n364 B.n171 585
R222 B.n370 B.n369 585
R223 B.n371 B.n370 585
R224 B.n2 B.n0 585
R225 B.n4 B.n2 585
R226 B.n3 B.n1 585
R227 B.n419 B.n3 585
R228 B.n417 B.n416 585
R229 B.n418 B.n417 585
R230 B.n415 B.n8 585
R231 B.n11 B.n8 585
R232 B.n414 B.n413 585
R233 B.n413 B.n412 585
R234 B.n10 B.n9 585
R235 B.n411 B.n10 585
R236 B.n409 B.n408 585
R237 B.n410 B.n409 585
R238 B.n407 B.n16 585
R239 B.n16 B.n15 585
R240 B.n406 B.n405 585
R241 B.n405 B.n404 585
R242 B.n18 B.n17 585
R243 B.n403 B.n18 585
R244 B.n401 B.n400 585
R245 B.n402 B.n401 585
R246 B.n399 B.n23 585
R247 B.n23 B.n22 585
R248 B.n398 B.n397 585
R249 B.n397 B.n396 585
R250 B.n25 B.n24 585
R251 B.n395 B.n25 585
R252 B.n422 B.n421 585
R253 B.n421 B.n420 585
R254 B.n330 B.n189 487.695
R255 B.n61 B.n25 487.695
R256 B.n334 B.n191 487.695
R257 B.n393 B.n27 487.695
R258 B.n394 B.n54 256.663
R259 B.n394 B.n53 256.663
R260 B.n394 B.n52 256.663
R261 B.n394 B.n51 256.663
R262 B.n394 B.n50 256.663
R263 B.n394 B.n49 256.663
R264 B.n394 B.n48 256.663
R265 B.n394 B.n47 256.663
R266 B.n394 B.n46 256.663
R267 B.n394 B.n45 256.663
R268 B.n394 B.n44 256.663
R269 B.n394 B.n43 256.663
R270 B.n394 B.n42 256.663
R271 B.n394 B.n41 256.663
R272 B.n394 B.n40 256.663
R273 B.n394 B.n39 256.663
R274 B.n394 B.n38 256.663
R275 B.n394 B.n37 256.663
R276 B.n394 B.n36 256.663
R277 B.n394 B.n35 256.663
R278 B.n394 B.n34 256.663
R279 B.n394 B.n33 256.663
R280 B.n394 B.n32 256.663
R281 B.n394 B.n31 256.663
R282 B.n394 B.n30 256.663
R283 B.n394 B.n29 256.663
R284 B.n394 B.n28 256.663
R285 B.n332 B.n331 256.663
R286 B.n332 B.n194 256.663
R287 B.n332 B.n195 256.663
R288 B.n332 B.n196 256.663
R289 B.n332 B.n197 256.663
R290 B.n332 B.n198 256.663
R291 B.n332 B.n199 256.663
R292 B.n332 B.n200 256.663
R293 B.n332 B.n201 256.663
R294 B.n332 B.n202 256.663
R295 B.n332 B.n203 256.663
R296 B.n332 B.n204 256.663
R297 B.n332 B.n205 256.663
R298 B.n332 B.n206 256.663
R299 B.n332 B.n207 256.663
R300 B.n332 B.n208 256.663
R301 B.n332 B.n209 256.663
R302 B.n332 B.n210 256.663
R303 B.n332 B.n211 256.663
R304 B.n332 B.n212 256.663
R305 B.n332 B.n213 256.663
R306 B.n332 B.n214 256.663
R307 B.n332 B.n215 256.663
R308 B.n332 B.n216 256.663
R309 B.n332 B.n217 256.663
R310 B.n332 B.n218 256.663
R311 B.n333 B.n332 256.663
R312 B.n340 B.n189 163.367
R313 B.n340 B.n187 163.367
R314 B.n344 B.n187 163.367
R315 B.n344 B.n181 163.367
R316 B.n352 B.n181 163.367
R317 B.n352 B.n179 163.367
R318 B.n356 B.n179 163.367
R319 B.n356 B.n173 163.367
R320 B.n366 B.n173 163.367
R321 B.n366 B.n171 163.367
R322 B.n370 B.n171 163.367
R323 B.n370 B.n2 163.367
R324 B.n421 B.n2 163.367
R325 B.n421 B.n3 163.367
R326 B.n417 B.n3 163.367
R327 B.n417 B.n8 163.367
R328 B.n413 B.n8 163.367
R329 B.n413 B.n10 163.367
R330 B.n409 B.n10 163.367
R331 B.n409 B.n16 163.367
R332 B.n405 B.n16 163.367
R333 B.n405 B.n18 163.367
R334 B.n401 B.n18 163.367
R335 B.n401 B.n23 163.367
R336 B.n397 B.n23 163.367
R337 B.n397 B.n25 163.367
R338 B.n220 B.n219 163.367
R339 B.n325 B.n219 163.367
R340 B.n323 B.n322 163.367
R341 B.n319 B.n318 163.367
R342 B.n315 B.n314 163.367
R343 B.n311 B.n310 163.367
R344 B.n307 B.n306 163.367
R345 B.n303 B.n302 163.367
R346 B.n299 B.n298 163.367
R347 B.n295 B.n294 163.367
R348 B.n291 B.n290 163.367
R349 B.n287 B.n286 163.367
R350 B.n283 B.n282 163.367
R351 B.n279 B.n278 163.367
R352 B.n275 B.n274 163.367
R353 B.n271 B.n270 163.367
R354 B.n266 B.n265 163.367
R355 B.n262 B.n261 163.367
R356 B.n258 B.n257 163.367
R357 B.n254 B.n253 163.367
R358 B.n250 B.n249 163.367
R359 B.n246 B.n245 163.367
R360 B.n242 B.n241 163.367
R361 B.n238 B.n237 163.367
R362 B.n234 B.n233 163.367
R363 B.n230 B.n229 163.367
R364 B.n226 B.n193 163.367
R365 B.n338 B.n191 163.367
R366 B.n338 B.n184 163.367
R367 B.n346 B.n184 163.367
R368 B.n346 B.n182 163.367
R369 B.n350 B.n182 163.367
R370 B.n350 B.n176 163.367
R371 B.n358 B.n176 163.367
R372 B.n358 B.n174 163.367
R373 B.n363 B.n174 163.367
R374 B.n363 B.n170 163.367
R375 B.n372 B.n170 163.367
R376 B.n373 B.n372 163.367
R377 B.n373 B.n5 163.367
R378 B.n6 B.n5 163.367
R379 B.n7 B.n6 163.367
R380 B.n378 B.n7 163.367
R381 B.n378 B.n12 163.367
R382 B.n13 B.n12 163.367
R383 B.n14 B.n13 163.367
R384 B.n383 B.n14 163.367
R385 B.n383 B.n19 163.367
R386 B.n20 B.n19 163.367
R387 B.n21 B.n20 163.367
R388 B.n388 B.n21 163.367
R389 B.n388 B.n26 163.367
R390 B.n27 B.n26 163.367
R391 B.n65 B.n64 163.367
R392 B.n69 B.n68 163.367
R393 B.n73 B.n72 163.367
R394 B.n77 B.n76 163.367
R395 B.n81 B.n80 163.367
R396 B.n85 B.n84 163.367
R397 B.n89 B.n88 163.367
R398 B.n93 B.n92 163.367
R399 B.n97 B.n96 163.367
R400 B.n101 B.n100 163.367
R401 B.n105 B.n104 163.367
R402 B.n110 B.n109 163.367
R403 B.n114 B.n113 163.367
R404 B.n118 B.n117 163.367
R405 B.n122 B.n121 163.367
R406 B.n126 B.n125 163.367
R407 B.n130 B.n129 163.367
R408 B.n134 B.n133 163.367
R409 B.n138 B.n137 163.367
R410 B.n142 B.n141 163.367
R411 B.n146 B.n145 163.367
R412 B.n150 B.n149 163.367
R413 B.n154 B.n153 163.367
R414 B.n158 B.n157 163.367
R415 B.n162 B.n161 163.367
R416 B.n166 B.n165 163.367
R417 B.n393 B.n55 163.367
R418 B.n332 B.n190 122.844
R419 B.n395 B.n394 122.844
R420 B.n224 B.t17 82.3444
R421 B.n56 B.t6 82.3444
R422 B.n221 B.t11 82.3386
R423 B.n59 B.t13 82.3386
R424 B.n225 B.t16 71.6778
R425 B.n57 B.t7 71.6778
R426 B.n331 B.n330 71.676
R427 B.n325 B.n194 71.676
R428 B.n322 B.n195 71.676
R429 B.n318 B.n196 71.676
R430 B.n314 B.n197 71.676
R431 B.n310 B.n198 71.676
R432 B.n306 B.n199 71.676
R433 B.n302 B.n200 71.676
R434 B.n298 B.n201 71.676
R435 B.n294 B.n202 71.676
R436 B.n290 B.n203 71.676
R437 B.n286 B.n204 71.676
R438 B.n282 B.n205 71.676
R439 B.n278 B.n206 71.676
R440 B.n274 B.n207 71.676
R441 B.n270 B.n208 71.676
R442 B.n265 B.n209 71.676
R443 B.n261 B.n210 71.676
R444 B.n257 B.n211 71.676
R445 B.n253 B.n212 71.676
R446 B.n249 B.n213 71.676
R447 B.n245 B.n214 71.676
R448 B.n241 B.n215 71.676
R449 B.n237 B.n216 71.676
R450 B.n233 B.n217 71.676
R451 B.n229 B.n218 71.676
R452 B.n333 B.n193 71.676
R453 B.n61 B.n28 71.676
R454 B.n65 B.n29 71.676
R455 B.n69 B.n30 71.676
R456 B.n73 B.n31 71.676
R457 B.n77 B.n32 71.676
R458 B.n81 B.n33 71.676
R459 B.n85 B.n34 71.676
R460 B.n89 B.n35 71.676
R461 B.n93 B.n36 71.676
R462 B.n97 B.n37 71.676
R463 B.n101 B.n38 71.676
R464 B.n105 B.n39 71.676
R465 B.n110 B.n40 71.676
R466 B.n114 B.n41 71.676
R467 B.n118 B.n42 71.676
R468 B.n122 B.n43 71.676
R469 B.n126 B.n44 71.676
R470 B.n130 B.n45 71.676
R471 B.n134 B.n46 71.676
R472 B.n138 B.n47 71.676
R473 B.n142 B.n48 71.676
R474 B.n146 B.n49 71.676
R475 B.n150 B.n50 71.676
R476 B.n154 B.n51 71.676
R477 B.n158 B.n52 71.676
R478 B.n162 B.n53 71.676
R479 B.n166 B.n54 71.676
R480 B.n55 B.n54 71.676
R481 B.n165 B.n53 71.676
R482 B.n161 B.n52 71.676
R483 B.n157 B.n51 71.676
R484 B.n153 B.n50 71.676
R485 B.n149 B.n49 71.676
R486 B.n145 B.n48 71.676
R487 B.n141 B.n47 71.676
R488 B.n137 B.n46 71.676
R489 B.n133 B.n45 71.676
R490 B.n129 B.n44 71.676
R491 B.n125 B.n43 71.676
R492 B.n121 B.n42 71.676
R493 B.n117 B.n41 71.676
R494 B.n113 B.n40 71.676
R495 B.n109 B.n39 71.676
R496 B.n104 B.n38 71.676
R497 B.n100 B.n37 71.676
R498 B.n96 B.n36 71.676
R499 B.n92 B.n35 71.676
R500 B.n88 B.n34 71.676
R501 B.n84 B.n33 71.676
R502 B.n80 B.n32 71.676
R503 B.n76 B.n31 71.676
R504 B.n72 B.n30 71.676
R505 B.n68 B.n29 71.676
R506 B.n64 B.n28 71.676
R507 B.n331 B.n220 71.676
R508 B.n323 B.n194 71.676
R509 B.n319 B.n195 71.676
R510 B.n315 B.n196 71.676
R511 B.n311 B.n197 71.676
R512 B.n307 B.n198 71.676
R513 B.n303 B.n199 71.676
R514 B.n299 B.n200 71.676
R515 B.n295 B.n201 71.676
R516 B.n291 B.n202 71.676
R517 B.n287 B.n203 71.676
R518 B.n283 B.n204 71.676
R519 B.n279 B.n205 71.676
R520 B.n275 B.n206 71.676
R521 B.n271 B.n207 71.676
R522 B.n266 B.n208 71.676
R523 B.n262 B.n209 71.676
R524 B.n258 B.n210 71.676
R525 B.n254 B.n211 71.676
R526 B.n250 B.n212 71.676
R527 B.n246 B.n213 71.676
R528 B.n242 B.n214 71.676
R529 B.n238 B.n215 71.676
R530 B.n234 B.n216 71.676
R531 B.n230 B.n217 71.676
R532 B.n226 B.n218 71.676
R533 B.n334 B.n333 71.676
R534 B.n222 B.t10 71.672
R535 B.n60 B.t14 71.672
R536 B.n339 B.n190 69.036
R537 B.n339 B.n185 69.036
R538 B.n345 B.n185 69.036
R539 B.n345 B.n186 69.036
R540 B.n351 B.n177 69.036
R541 B.n357 B.n177 69.036
R542 B.n357 B.n178 69.036
R543 B.n365 B.n364 69.036
R544 B.n371 B.n4 69.036
R545 B.n420 B.n4 69.036
R546 B.n420 B.n419 69.036
R547 B.n419 B.n418 69.036
R548 B.n412 B.n11 69.036
R549 B.n411 B.n410 69.036
R550 B.n410 B.n15 69.036
R551 B.n404 B.n15 69.036
R552 B.n403 B.n402 69.036
R553 B.n402 B.n22 69.036
R554 B.n396 B.n22 69.036
R555 B.n396 B.n395 69.036
R556 B.n178 B.t2 67.0056
R557 B.t0 B.n411 67.0056
R558 B.n268 B.n225 59.5399
R559 B.n223 B.n222 59.5399
R560 B.n107 B.n60 59.5399
R561 B.n58 B.n57 59.5399
R562 B.n351 B.t9 58.8838
R563 B.n404 B.t5 58.8838
R564 B.n364 B.t1 40.6096
R565 B.n11 B.t3 40.6096
R566 B.n62 B.n24 31.6883
R567 B.n392 B.n391 31.6883
R568 B.n336 B.n335 31.6883
R569 B.n329 B.n188 31.6883
R570 B.n371 B.t1 28.4269
R571 B.n418 B.t3 28.4269
R572 B B.n422 18.0485
R573 B.n225 B.n224 10.6672
R574 B.n222 B.n221 10.6672
R575 B.n60 B.n59 10.6672
R576 B.n57 B.n56 10.6672
R577 B.n63 B.n62 10.6151
R578 B.n66 B.n63 10.6151
R579 B.n67 B.n66 10.6151
R580 B.n70 B.n67 10.6151
R581 B.n71 B.n70 10.6151
R582 B.n74 B.n71 10.6151
R583 B.n75 B.n74 10.6151
R584 B.n78 B.n75 10.6151
R585 B.n79 B.n78 10.6151
R586 B.n82 B.n79 10.6151
R587 B.n83 B.n82 10.6151
R588 B.n86 B.n83 10.6151
R589 B.n87 B.n86 10.6151
R590 B.n90 B.n87 10.6151
R591 B.n91 B.n90 10.6151
R592 B.n94 B.n91 10.6151
R593 B.n95 B.n94 10.6151
R594 B.n98 B.n95 10.6151
R595 B.n99 B.n98 10.6151
R596 B.n102 B.n99 10.6151
R597 B.n103 B.n102 10.6151
R598 B.n106 B.n103 10.6151
R599 B.n111 B.n108 10.6151
R600 B.n112 B.n111 10.6151
R601 B.n115 B.n112 10.6151
R602 B.n116 B.n115 10.6151
R603 B.n119 B.n116 10.6151
R604 B.n120 B.n119 10.6151
R605 B.n123 B.n120 10.6151
R606 B.n124 B.n123 10.6151
R607 B.n128 B.n127 10.6151
R608 B.n131 B.n128 10.6151
R609 B.n132 B.n131 10.6151
R610 B.n135 B.n132 10.6151
R611 B.n136 B.n135 10.6151
R612 B.n139 B.n136 10.6151
R613 B.n140 B.n139 10.6151
R614 B.n143 B.n140 10.6151
R615 B.n144 B.n143 10.6151
R616 B.n147 B.n144 10.6151
R617 B.n148 B.n147 10.6151
R618 B.n151 B.n148 10.6151
R619 B.n152 B.n151 10.6151
R620 B.n155 B.n152 10.6151
R621 B.n156 B.n155 10.6151
R622 B.n159 B.n156 10.6151
R623 B.n160 B.n159 10.6151
R624 B.n163 B.n160 10.6151
R625 B.n164 B.n163 10.6151
R626 B.n167 B.n164 10.6151
R627 B.n168 B.n167 10.6151
R628 B.n392 B.n168 10.6151
R629 B.n337 B.n336 10.6151
R630 B.n337 B.n183 10.6151
R631 B.n347 B.n183 10.6151
R632 B.n348 B.n347 10.6151
R633 B.n349 B.n348 10.6151
R634 B.n349 B.n175 10.6151
R635 B.n359 B.n175 10.6151
R636 B.n360 B.n359 10.6151
R637 B.n362 B.n360 10.6151
R638 B.n362 B.n361 10.6151
R639 B.n361 B.n169 10.6151
R640 B.n374 B.n169 10.6151
R641 B.n375 B.n374 10.6151
R642 B.n376 B.n375 10.6151
R643 B.n377 B.n376 10.6151
R644 B.n379 B.n377 10.6151
R645 B.n380 B.n379 10.6151
R646 B.n381 B.n380 10.6151
R647 B.n382 B.n381 10.6151
R648 B.n384 B.n382 10.6151
R649 B.n385 B.n384 10.6151
R650 B.n386 B.n385 10.6151
R651 B.n387 B.n386 10.6151
R652 B.n389 B.n387 10.6151
R653 B.n390 B.n389 10.6151
R654 B.n391 B.n390 10.6151
R655 B.n329 B.n328 10.6151
R656 B.n328 B.n327 10.6151
R657 B.n327 B.n326 10.6151
R658 B.n326 B.n324 10.6151
R659 B.n324 B.n321 10.6151
R660 B.n321 B.n320 10.6151
R661 B.n320 B.n317 10.6151
R662 B.n317 B.n316 10.6151
R663 B.n316 B.n313 10.6151
R664 B.n313 B.n312 10.6151
R665 B.n312 B.n309 10.6151
R666 B.n309 B.n308 10.6151
R667 B.n308 B.n305 10.6151
R668 B.n305 B.n304 10.6151
R669 B.n304 B.n301 10.6151
R670 B.n301 B.n300 10.6151
R671 B.n300 B.n297 10.6151
R672 B.n297 B.n296 10.6151
R673 B.n296 B.n293 10.6151
R674 B.n293 B.n292 10.6151
R675 B.n292 B.n289 10.6151
R676 B.n289 B.n288 10.6151
R677 B.n285 B.n284 10.6151
R678 B.n284 B.n281 10.6151
R679 B.n281 B.n280 10.6151
R680 B.n280 B.n277 10.6151
R681 B.n277 B.n276 10.6151
R682 B.n276 B.n273 10.6151
R683 B.n273 B.n272 10.6151
R684 B.n272 B.n269 10.6151
R685 B.n267 B.n264 10.6151
R686 B.n264 B.n263 10.6151
R687 B.n263 B.n260 10.6151
R688 B.n260 B.n259 10.6151
R689 B.n259 B.n256 10.6151
R690 B.n256 B.n255 10.6151
R691 B.n255 B.n252 10.6151
R692 B.n252 B.n251 10.6151
R693 B.n251 B.n248 10.6151
R694 B.n248 B.n247 10.6151
R695 B.n247 B.n244 10.6151
R696 B.n244 B.n243 10.6151
R697 B.n243 B.n240 10.6151
R698 B.n240 B.n239 10.6151
R699 B.n239 B.n236 10.6151
R700 B.n236 B.n235 10.6151
R701 B.n235 B.n232 10.6151
R702 B.n232 B.n231 10.6151
R703 B.n231 B.n228 10.6151
R704 B.n228 B.n227 10.6151
R705 B.n227 B.n192 10.6151
R706 B.n335 B.n192 10.6151
R707 B.n341 B.n188 10.6151
R708 B.n342 B.n341 10.6151
R709 B.n343 B.n342 10.6151
R710 B.n343 B.n180 10.6151
R711 B.n353 B.n180 10.6151
R712 B.n354 B.n353 10.6151
R713 B.n355 B.n354 10.6151
R714 B.n355 B.n172 10.6151
R715 B.n367 B.n172 10.6151
R716 B.n368 B.n367 10.6151
R717 B.n369 B.n368 10.6151
R718 B.n369 B.n0 10.6151
R719 B.n416 B.n1 10.6151
R720 B.n416 B.n415 10.6151
R721 B.n415 B.n414 10.6151
R722 B.n414 B.n9 10.6151
R723 B.n408 B.n9 10.6151
R724 B.n408 B.n407 10.6151
R725 B.n407 B.n406 10.6151
R726 B.n406 B.n17 10.6151
R727 B.n400 B.n17 10.6151
R728 B.n400 B.n399 10.6151
R729 B.n399 B.n398 10.6151
R730 B.n398 B.n24 10.6151
R731 B.n186 B.t9 10.1528
R732 B.t5 B.n403 10.1528
R733 B.n108 B.n107 7.18099
R734 B.n124 B.n58 7.18099
R735 B.n285 B.n223 7.18099
R736 B.n269 B.n268 7.18099
R737 B.n107 B.n106 3.43465
R738 B.n127 B.n58 3.43465
R739 B.n288 B.n223 3.43465
R740 B.n268 B.n267 3.43465
R741 B.n422 B.n0 2.81026
R742 B.n422 B.n1 2.81026
R743 B.n365 B.t2 2.03096
R744 B.n412 B.t0 2.03096
R745 VP.n1 VP.t3 789.458
R746 VP.n1 VP.t2 789.458
R747 VP.n0 VP.t1 789.458
R748 VP.n0 VP.t0 789.458
R749 VP.n2 VP.n0 195.392
R750 VP.n2 VP.n1 161.3
R751 VP VP.n2 0.0516364
R752 VDD1 VDD1.n1 96.3855
R753 VDD1 VDD1.n0 65.9887
R754 VDD1.n0 VDD1.t2 3.57451
R755 VDD1.n0 VDD1.t3 3.57451
R756 VDD1.n1 VDD1.t1 3.57451
R757 VDD1.n1 VDD1.t0 3.57451
C0 VDD2 VTAIL 5.60235f
C1 VN VTAIL 0.741227f
C2 VP VDD2 0.244334f
C3 VP VN 3.2749f
C4 VDD2 VN 0.970097f
C5 VDD1 VTAIL 5.5641f
C6 VP VDD1 1.06598f
C7 VDD2 VDD1 0.462207f
C8 VDD1 VN 0.148321f
C9 VP VTAIL 0.755333f
C10 VDD2 B 1.91215f
C11 VDD1 B 4.66318f
C12 VTAIL B 4.513675f
C13 VN B 5.68573f
C14 VP B 3.393206f
C15 VDD1.t2 B 0.123949f
C16 VDD1.t3 B 0.123949f
C17 VDD1.n0 B 1.02304f
C18 VDD1.t1 B 0.123949f
C19 VDD1.t0 B 0.123949f
C20 VDD1.n1 B 1.40969f
C21 VP.t1 B 0.148f
C22 VP.t0 B 0.148f
C23 VP.n0 B 0.356117f
C24 VP.t2 B 0.148f
C25 VP.t3 B 0.148f
C26 VP.n1 B 0.149907f
C27 VP.n2 B 2.18572f
C28 VDD2.t2 B 0.126308f
C29 VDD2.t0 B 0.126308f
C30 VDD2.n0 B 1.41321f
C31 VDD2.t1 B 0.126308f
C32 VDD2.t3 B 0.126308f
C33 VDD2.n1 B 1.04225f
C34 VDD2.n2 B 2.58902f
C35 VTAIL.t7 B 0.824763f
C36 VTAIL.n0 B 0.283071f
C37 VTAIL.t1 B 0.824763f
C38 VTAIL.n1 B 0.294225f
C39 VTAIL.t2 B 0.824763f
C40 VTAIL.n2 B 0.856249f
C41 VTAIL.t6 B 0.824767f
C42 VTAIL.n3 B 0.856245f
C43 VTAIL.t5 B 0.824767f
C44 VTAIL.n4 B 0.294221f
C45 VTAIL.t3 B 0.824767f
C46 VTAIL.n5 B 0.294221f
C47 VTAIL.t0 B 0.824763f
C48 VTAIL.n6 B 0.856249f
C49 VTAIL.t4 B 0.824763f
C50 VTAIL.n7 B 0.837838f
C51 VN.t1 B 0.145428f
C52 VN.t3 B 0.145428f
C53 VN.n0 B 0.147314f
C54 VN.t2 B 0.145428f
C55 VN.t0 B 0.145428f
C56 VN.n1 B 0.356577f
.ends

