* NGSPICE file created from diff_pair_sample_1084.ext - technology: sky130A

.subckt diff_pair_sample_1084 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=6.6885 pd=35.08 as=0 ps=0 w=17.15 l=2.44
X1 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=6.6885 pd=35.08 as=0 ps=0 w=17.15 l=2.44
X2 VDD2.t3 VN.t0 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=2.82975 pd=17.48 as=6.6885 ps=35.08 w=17.15 l=2.44
X3 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=6.6885 pd=35.08 as=0 ps=0 w=17.15 l=2.44
X4 VTAIL.t5 VN.t1 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=6.6885 pd=35.08 as=2.82975 ps=17.48 w=17.15 l=2.44
X5 VTAIL.t4 VN.t2 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=6.6885 pd=35.08 as=2.82975 ps=17.48 w=17.15 l=2.44
X6 VDD2.t0 VN.t3 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.82975 pd=17.48 as=6.6885 ps=35.08 w=17.15 l=2.44
X7 VDD1.t3 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.82975 pd=17.48 as=6.6885 ps=35.08 w=17.15 l=2.44
X8 VDD1.t2 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.82975 pd=17.48 as=6.6885 ps=35.08 w=17.15 l=2.44
X9 VTAIL.t1 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.6885 pd=35.08 as=2.82975 ps=17.48 w=17.15 l=2.44
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.6885 pd=35.08 as=0 ps=0 w=17.15 l=2.44
X11 VTAIL.t2 VP.t3 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=6.6885 pd=35.08 as=2.82975 ps=17.48 w=17.15 l=2.44
R0 B.n887 B.n886 585
R1 B.n888 B.n887 585
R2 B.n371 B.n124 585
R3 B.n370 B.n369 585
R4 B.n368 B.n367 585
R5 B.n366 B.n365 585
R6 B.n364 B.n363 585
R7 B.n362 B.n361 585
R8 B.n360 B.n359 585
R9 B.n358 B.n357 585
R10 B.n356 B.n355 585
R11 B.n354 B.n353 585
R12 B.n352 B.n351 585
R13 B.n350 B.n349 585
R14 B.n348 B.n347 585
R15 B.n346 B.n345 585
R16 B.n344 B.n343 585
R17 B.n342 B.n341 585
R18 B.n340 B.n339 585
R19 B.n338 B.n337 585
R20 B.n336 B.n335 585
R21 B.n334 B.n333 585
R22 B.n332 B.n331 585
R23 B.n330 B.n329 585
R24 B.n328 B.n327 585
R25 B.n326 B.n325 585
R26 B.n324 B.n323 585
R27 B.n322 B.n321 585
R28 B.n320 B.n319 585
R29 B.n318 B.n317 585
R30 B.n316 B.n315 585
R31 B.n314 B.n313 585
R32 B.n312 B.n311 585
R33 B.n310 B.n309 585
R34 B.n308 B.n307 585
R35 B.n306 B.n305 585
R36 B.n304 B.n303 585
R37 B.n302 B.n301 585
R38 B.n300 B.n299 585
R39 B.n298 B.n297 585
R40 B.n296 B.n295 585
R41 B.n294 B.n293 585
R42 B.n292 B.n291 585
R43 B.n290 B.n289 585
R44 B.n288 B.n287 585
R45 B.n286 B.n285 585
R46 B.n284 B.n283 585
R47 B.n282 B.n281 585
R48 B.n280 B.n279 585
R49 B.n278 B.n277 585
R50 B.n276 B.n275 585
R51 B.n274 B.n273 585
R52 B.n272 B.n271 585
R53 B.n270 B.n269 585
R54 B.n268 B.n267 585
R55 B.n266 B.n265 585
R56 B.n264 B.n263 585
R57 B.n262 B.n261 585
R58 B.n260 B.n259 585
R59 B.n258 B.n257 585
R60 B.n256 B.n255 585
R61 B.n254 B.n253 585
R62 B.n252 B.n251 585
R63 B.n250 B.n249 585
R64 B.n248 B.n247 585
R65 B.n246 B.n245 585
R66 B.n244 B.n243 585
R67 B.n241 B.n240 585
R68 B.n239 B.n238 585
R69 B.n237 B.n236 585
R70 B.n235 B.n234 585
R71 B.n233 B.n232 585
R72 B.n231 B.n230 585
R73 B.n229 B.n228 585
R74 B.n227 B.n226 585
R75 B.n225 B.n224 585
R76 B.n223 B.n222 585
R77 B.n221 B.n220 585
R78 B.n219 B.n218 585
R79 B.n217 B.n216 585
R80 B.n215 B.n214 585
R81 B.n213 B.n212 585
R82 B.n211 B.n210 585
R83 B.n209 B.n208 585
R84 B.n207 B.n206 585
R85 B.n205 B.n204 585
R86 B.n203 B.n202 585
R87 B.n201 B.n200 585
R88 B.n199 B.n198 585
R89 B.n197 B.n196 585
R90 B.n195 B.n194 585
R91 B.n193 B.n192 585
R92 B.n191 B.n190 585
R93 B.n189 B.n188 585
R94 B.n187 B.n186 585
R95 B.n185 B.n184 585
R96 B.n183 B.n182 585
R97 B.n181 B.n180 585
R98 B.n179 B.n178 585
R99 B.n177 B.n176 585
R100 B.n175 B.n174 585
R101 B.n173 B.n172 585
R102 B.n171 B.n170 585
R103 B.n169 B.n168 585
R104 B.n167 B.n166 585
R105 B.n165 B.n164 585
R106 B.n163 B.n162 585
R107 B.n161 B.n160 585
R108 B.n159 B.n158 585
R109 B.n157 B.n156 585
R110 B.n155 B.n154 585
R111 B.n153 B.n152 585
R112 B.n151 B.n150 585
R113 B.n149 B.n148 585
R114 B.n147 B.n146 585
R115 B.n145 B.n144 585
R116 B.n143 B.n142 585
R117 B.n141 B.n140 585
R118 B.n139 B.n138 585
R119 B.n137 B.n136 585
R120 B.n135 B.n134 585
R121 B.n133 B.n132 585
R122 B.n131 B.n130 585
R123 B.n61 B.n60 585
R124 B.n885 B.n62 585
R125 B.n889 B.n62 585
R126 B.n884 B.n883 585
R127 B.n883 B.n58 585
R128 B.n882 B.n57 585
R129 B.n895 B.n57 585
R130 B.n881 B.n56 585
R131 B.n896 B.n56 585
R132 B.n880 B.n55 585
R133 B.n897 B.n55 585
R134 B.n879 B.n878 585
R135 B.n878 B.n51 585
R136 B.n877 B.n50 585
R137 B.n903 B.n50 585
R138 B.n876 B.n49 585
R139 B.n904 B.n49 585
R140 B.n875 B.n48 585
R141 B.n905 B.n48 585
R142 B.n874 B.n873 585
R143 B.n873 B.n44 585
R144 B.n872 B.n43 585
R145 B.n911 B.n43 585
R146 B.n871 B.n42 585
R147 B.n912 B.n42 585
R148 B.n870 B.n41 585
R149 B.n913 B.n41 585
R150 B.n869 B.n868 585
R151 B.n868 B.n37 585
R152 B.n867 B.n36 585
R153 B.n919 B.n36 585
R154 B.n866 B.n35 585
R155 B.n920 B.n35 585
R156 B.n865 B.n34 585
R157 B.n921 B.n34 585
R158 B.n864 B.n863 585
R159 B.n863 B.n30 585
R160 B.n862 B.n29 585
R161 B.n927 B.n29 585
R162 B.n861 B.n28 585
R163 B.n928 B.n28 585
R164 B.n860 B.n27 585
R165 B.n929 B.n27 585
R166 B.n859 B.n858 585
R167 B.n858 B.n23 585
R168 B.n857 B.n22 585
R169 B.n935 B.n22 585
R170 B.n856 B.n21 585
R171 B.n936 B.n21 585
R172 B.n855 B.n20 585
R173 B.n937 B.n20 585
R174 B.n854 B.n853 585
R175 B.n853 B.n16 585
R176 B.n852 B.n15 585
R177 B.n943 B.n15 585
R178 B.n851 B.n14 585
R179 B.n944 B.n14 585
R180 B.n850 B.n13 585
R181 B.n945 B.n13 585
R182 B.n849 B.n848 585
R183 B.n848 B.n12 585
R184 B.n847 B.n846 585
R185 B.n847 B.n8 585
R186 B.n845 B.n7 585
R187 B.n952 B.n7 585
R188 B.n844 B.n6 585
R189 B.n953 B.n6 585
R190 B.n843 B.n5 585
R191 B.n954 B.n5 585
R192 B.n842 B.n841 585
R193 B.n841 B.n4 585
R194 B.n840 B.n372 585
R195 B.n840 B.n839 585
R196 B.n830 B.n373 585
R197 B.n374 B.n373 585
R198 B.n832 B.n831 585
R199 B.n833 B.n832 585
R200 B.n829 B.n379 585
R201 B.n379 B.n378 585
R202 B.n828 B.n827 585
R203 B.n827 B.n826 585
R204 B.n381 B.n380 585
R205 B.n382 B.n381 585
R206 B.n819 B.n818 585
R207 B.n820 B.n819 585
R208 B.n817 B.n387 585
R209 B.n387 B.n386 585
R210 B.n816 B.n815 585
R211 B.n815 B.n814 585
R212 B.n389 B.n388 585
R213 B.n390 B.n389 585
R214 B.n807 B.n806 585
R215 B.n808 B.n807 585
R216 B.n805 B.n395 585
R217 B.n395 B.n394 585
R218 B.n804 B.n803 585
R219 B.n803 B.n802 585
R220 B.n397 B.n396 585
R221 B.n398 B.n397 585
R222 B.n795 B.n794 585
R223 B.n796 B.n795 585
R224 B.n793 B.n403 585
R225 B.n403 B.n402 585
R226 B.n792 B.n791 585
R227 B.n791 B.n790 585
R228 B.n405 B.n404 585
R229 B.n406 B.n405 585
R230 B.n783 B.n782 585
R231 B.n784 B.n783 585
R232 B.n781 B.n411 585
R233 B.n411 B.n410 585
R234 B.n780 B.n779 585
R235 B.n779 B.n778 585
R236 B.n413 B.n412 585
R237 B.n414 B.n413 585
R238 B.n771 B.n770 585
R239 B.n772 B.n771 585
R240 B.n769 B.n418 585
R241 B.n422 B.n418 585
R242 B.n768 B.n767 585
R243 B.n767 B.n766 585
R244 B.n420 B.n419 585
R245 B.n421 B.n420 585
R246 B.n759 B.n758 585
R247 B.n760 B.n759 585
R248 B.n757 B.n427 585
R249 B.n427 B.n426 585
R250 B.n756 B.n755 585
R251 B.n755 B.n754 585
R252 B.n429 B.n428 585
R253 B.n430 B.n429 585
R254 B.n747 B.n746 585
R255 B.n748 B.n747 585
R256 B.n433 B.n432 585
R257 B.n503 B.n502 585
R258 B.n504 B.n500 585
R259 B.n500 B.n434 585
R260 B.n506 B.n505 585
R261 B.n508 B.n499 585
R262 B.n511 B.n510 585
R263 B.n512 B.n498 585
R264 B.n514 B.n513 585
R265 B.n516 B.n497 585
R266 B.n519 B.n518 585
R267 B.n520 B.n496 585
R268 B.n522 B.n521 585
R269 B.n524 B.n495 585
R270 B.n527 B.n526 585
R271 B.n528 B.n494 585
R272 B.n530 B.n529 585
R273 B.n532 B.n493 585
R274 B.n535 B.n534 585
R275 B.n536 B.n492 585
R276 B.n538 B.n537 585
R277 B.n540 B.n491 585
R278 B.n543 B.n542 585
R279 B.n544 B.n490 585
R280 B.n546 B.n545 585
R281 B.n548 B.n489 585
R282 B.n551 B.n550 585
R283 B.n552 B.n488 585
R284 B.n554 B.n553 585
R285 B.n556 B.n487 585
R286 B.n559 B.n558 585
R287 B.n560 B.n486 585
R288 B.n562 B.n561 585
R289 B.n564 B.n485 585
R290 B.n567 B.n566 585
R291 B.n568 B.n484 585
R292 B.n570 B.n569 585
R293 B.n572 B.n483 585
R294 B.n575 B.n574 585
R295 B.n576 B.n482 585
R296 B.n578 B.n577 585
R297 B.n580 B.n481 585
R298 B.n583 B.n582 585
R299 B.n584 B.n480 585
R300 B.n586 B.n585 585
R301 B.n588 B.n479 585
R302 B.n591 B.n590 585
R303 B.n592 B.n478 585
R304 B.n594 B.n593 585
R305 B.n596 B.n477 585
R306 B.n599 B.n598 585
R307 B.n600 B.n476 585
R308 B.n602 B.n601 585
R309 B.n604 B.n475 585
R310 B.n607 B.n606 585
R311 B.n608 B.n474 585
R312 B.n610 B.n609 585
R313 B.n612 B.n473 585
R314 B.n615 B.n614 585
R315 B.n616 B.n469 585
R316 B.n618 B.n617 585
R317 B.n620 B.n468 585
R318 B.n623 B.n622 585
R319 B.n624 B.n467 585
R320 B.n626 B.n625 585
R321 B.n628 B.n466 585
R322 B.n631 B.n630 585
R323 B.n633 B.n463 585
R324 B.n635 B.n634 585
R325 B.n637 B.n462 585
R326 B.n640 B.n639 585
R327 B.n641 B.n461 585
R328 B.n643 B.n642 585
R329 B.n645 B.n460 585
R330 B.n648 B.n647 585
R331 B.n649 B.n459 585
R332 B.n651 B.n650 585
R333 B.n653 B.n458 585
R334 B.n656 B.n655 585
R335 B.n657 B.n457 585
R336 B.n659 B.n658 585
R337 B.n661 B.n456 585
R338 B.n664 B.n663 585
R339 B.n665 B.n455 585
R340 B.n667 B.n666 585
R341 B.n669 B.n454 585
R342 B.n672 B.n671 585
R343 B.n673 B.n453 585
R344 B.n675 B.n674 585
R345 B.n677 B.n452 585
R346 B.n680 B.n679 585
R347 B.n681 B.n451 585
R348 B.n683 B.n682 585
R349 B.n685 B.n450 585
R350 B.n688 B.n687 585
R351 B.n689 B.n449 585
R352 B.n691 B.n690 585
R353 B.n693 B.n448 585
R354 B.n696 B.n695 585
R355 B.n697 B.n447 585
R356 B.n699 B.n698 585
R357 B.n701 B.n446 585
R358 B.n704 B.n703 585
R359 B.n705 B.n445 585
R360 B.n707 B.n706 585
R361 B.n709 B.n444 585
R362 B.n712 B.n711 585
R363 B.n713 B.n443 585
R364 B.n715 B.n714 585
R365 B.n717 B.n442 585
R366 B.n720 B.n719 585
R367 B.n721 B.n441 585
R368 B.n723 B.n722 585
R369 B.n725 B.n440 585
R370 B.n728 B.n727 585
R371 B.n729 B.n439 585
R372 B.n731 B.n730 585
R373 B.n733 B.n438 585
R374 B.n736 B.n735 585
R375 B.n737 B.n437 585
R376 B.n739 B.n738 585
R377 B.n741 B.n436 585
R378 B.n744 B.n743 585
R379 B.n745 B.n435 585
R380 B.n750 B.n749 585
R381 B.n749 B.n748 585
R382 B.n751 B.n431 585
R383 B.n431 B.n430 585
R384 B.n753 B.n752 585
R385 B.n754 B.n753 585
R386 B.n425 B.n424 585
R387 B.n426 B.n425 585
R388 B.n762 B.n761 585
R389 B.n761 B.n760 585
R390 B.n763 B.n423 585
R391 B.n423 B.n421 585
R392 B.n765 B.n764 585
R393 B.n766 B.n765 585
R394 B.n417 B.n416 585
R395 B.n422 B.n417 585
R396 B.n774 B.n773 585
R397 B.n773 B.n772 585
R398 B.n775 B.n415 585
R399 B.n415 B.n414 585
R400 B.n777 B.n776 585
R401 B.n778 B.n777 585
R402 B.n409 B.n408 585
R403 B.n410 B.n409 585
R404 B.n786 B.n785 585
R405 B.n785 B.n784 585
R406 B.n787 B.n407 585
R407 B.n407 B.n406 585
R408 B.n789 B.n788 585
R409 B.n790 B.n789 585
R410 B.n401 B.n400 585
R411 B.n402 B.n401 585
R412 B.n798 B.n797 585
R413 B.n797 B.n796 585
R414 B.n799 B.n399 585
R415 B.n399 B.n398 585
R416 B.n801 B.n800 585
R417 B.n802 B.n801 585
R418 B.n393 B.n392 585
R419 B.n394 B.n393 585
R420 B.n810 B.n809 585
R421 B.n809 B.n808 585
R422 B.n811 B.n391 585
R423 B.n391 B.n390 585
R424 B.n813 B.n812 585
R425 B.n814 B.n813 585
R426 B.n385 B.n384 585
R427 B.n386 B.n385 585
R428 B.n822 B.n821 585
R429 B.n821 B.n820 585
R430 B.n823 B.n383 585
R431 B.n383 B.n382 585
R432 B.n825 B.n824 585
R433 B.n826 B.n825 585
R434 B.n377 B.n376 585
R435 B.n378 B.n377 585
R436 B.n835 B.n834 585
R437 B.n834 B.n833 585
R438 B.n836 B.n375 585
R439 B.n375 B.n374 585
R440 B.n838 B.n837 585
R441 B.n839 B.n838 585
R442 B.n3 B.n0 585
R443 B.n4 B.n3 585
R444 B.n951 B.n1 585
R445 B.n952 B.n951 585
R446 B.n950 B.n949 585
R447 B.n950 B.n8 585
R448 B.n948 B.n9 585
R449 B.n12 B.n9 585
R450 B.n947 B.n946 585
R451 B.n946 B.n945 585
R452 B.n11 B.n10 585
R453 B.n944 B.n11 585
R454 B.n942 B.n941 585
R455 B.n943 B.n942 585
R456 B.n940 B.n17 585
R457 B.n17 B.n16 585
R458 B.n939 B.n938 585
R459 B.n938 B.n937 585
R460 B.n19 B.n18 585
R461 B.n936 B.n19 585
R462 B.n934 B.n933 585
R463 B.n935 B.n934 585
R464 B.n932 B.n24 585
R465 B.n24 B.n23 585
R466 B.n931 B.n930 585
R467 B.n930 B.n929 585
R468 B.n26 B.n25 585
R469 B.n928 B.n26 585
R470 B.n926 B.n925 585
R471 B.n927 B.n926 585
R472 B.n924 B.n31 585
R473 B.n31 B.n30 585
R474 B.n923 B.n922 585
R475 B.n922 B.n921 585
R476 B.n33 B.n32 585
R477 B.n920 B.n33 585
R478 B.n918 B.n917 585
R479 B.n919 B.n918 585
R480 B.n916 B.n38 585
R481 B.n38 B.n37 585
R482 B.n915 B.n914 585
R483 B.n914 B.n913 585
R484 B.n40 B.n39 585
R485 B.n912 B.n40 585
R486 B.n910 B.n909 585
R487 B.n911 B.n910 585
R488 B.n908 B.n45 585
R489 B.n45 B.n44 585
R490 B.n907 B.n906 585
R491 B.n906 B.n905 585
R492 B.n47 B.n46 585
R493 B.n904 B.n47 585
R494 B.n902 B.n901 585
R495 B.n903 B.n902 585
R496 B.n900 B.n52 585
R497 B.n52 B.n51 585
R498 B.n899 B.n898 585
R499 B.n898 B.n897 585
R500 B.n54 B.n53 585
R501 B.n896 B.n54 585
R502 B.n894 B.n893 585
R503 B.n895 B.n894 585
R504 B.n892 B.n59 585
R505 B.n59 B.n58 585
R506 B.n891 B.n890 585
R507 B.n890 B.n889 585
R508 B.n955 B.n954 585
R509 B.n953 B.n2 585
R510 B.n890 B.n61 516.524
R511 B.n887 B.n62 516.524
R512 B.n747 B.n435 516.524
R513 B.n749 B.n433 516.524
R514 B.n128 B.t8 377.183
R515 B.n125 B.t4 377.183
R516 B.n464 B.t15 377.183
R517 B.n470 B.t11 377.183
R518 B.n888 B.n123 256.663
R519 B.n888 B.n122 256.663
R520 B.n888 B.n121 256.663
R521 B.n888 B.n120 256.663
R522 B.n888 B.n119 256.663
R523 B.n888 B.n118 256.663
R524 B.n888 B.n117 256.663
R525 B.n888 B.n116 256.663
R526 B.n888 B.n115 256.663
R527 B.n888 B.n114 256.663
R528 B.n888 B.n113 256.663
R529 B.n888 B.n112 256.663
R530 B.n888 B.n111 256.663
R531 B.n888 B.n110 256.663
R532 B.n888 B.n109 256.663
R533 B.n888 B.n108 256.663
R534 B.n888 B.n107 256.663
R535 B.n888 B.n106 256.663
R536 B.n888 B.n105 256.663
R537 B.n888 B.n104 256.663
R538 B.n888 B.n103 256.663
R539 B.n888 B.n102 256.663
R540 B.n888 B.n101 256.663
R541 B.n888 B.n100 256.663
R542 B.n888 B.n99 256.663
R543 B.n888 B.n98 256.663
R544 B.n888 B.n97 256.663
R545 B.n888 B.n96 256.663
R546 B.n888 B.n95 256.663
R547 B.n888 B.n94 256.663
R548 B.n888 B.n93 256.663
R549 B.n888 B.n92 256.663
R550 B.n888 B.n91 256.663
R551 B.n888 B.n90 256.663
R552 B.n888 B.n89 256.663
R553 B.n888 B.n88 256.663
R554 B.n888 B.n87 256.663
R555 B.n888 B.n86 256.663
R556 B.n888 B.n85 256.663
R557 B.n888 B.n84 256.663
R558 B.n888 B.n83 256.663
R559 B.n888 B.n82 256.663
R560 B.n888 B.n81 256.663
R561 B.n888 B.n80 256.663
R562 B.n888 B.n79 256.663
R563 B.n888 B.n78 256.663
R564 B.n888 B.n77 256.663
R565 B.n888 B.n76 256.663
R566 B.n888 B.n75 256.663
R567 B.n888 B.n74 256.663
R568 B.n888 B.n73 256.663
R569 B.n888 B.n72 256.663
R570 B.n888 B.n71 256.663
R571 B.n888 B.n70 256.663
R572 B.n888 B.n69 256.663
R573 B.n888 B.n68 256.663
R574 B.n888 B.n67 256.663
R575 B.n888 B.n66 256.663
R576 B.n888 B.n65 256.663
R577 B.n888 B.n64 256.663
R578 B.n888 B.n63 256.663
R579 B.n501 B.n434 256.663
R580 B.n507 B.n434 256.663
R581 B.n509 B.n434 256.663
R582 B.n515 B.n434 256.663
R583 B.n517 B.n434 256.663
R584 B.n523 B.n434 256.663
R585 B.n525 B.n434 256.663
R586 B.n531 B.n434 256.663
R587 B.n533 B.n434 256.663
R588 B.n539 B.n434 256.663
R589 B.n541 B.n434 256.663
R590 B.n547 B.n434 256.663
R591 B.n549 B.n434 256.663
R592 B.n555 B.n434 256.663
R593 B.n557 B.n434 256.663
R594 B.n563 B.n434 256.663
R595 B.n565 B.n434 256.663
R596 B.n571 B.n434 256.663
R597 B.n573 B.n434 256.663
R598 B.n579 B.n434 256.663
R599 B.n581 B.n434 256.663
R600 B.n587 B.n434 256.663
R601 B.n589 B.n434 256.663
R602 B.n595 B.n434 256.663
R603 B.n597 B.n434 256.663
R604 B.n603 B.n434 256.663
R605 B.n605 B.n434 256.663
R606 B.n611 B.n434 256.663
R607 B.n613 B.n434 256.663
R608 B.n619 B.n434 256.663
R609 B.n621 B.n434 256.663
R610 B.n627 B.n434 256.663
R611 B.n629 B.n434 256.663
R612 B.n636 B.n434 256.663
R613 B.n638 B.n434 256.663
R614 B.n644 B.n434 256.663
R615 B.n646 B.n434 256.663
R616 B.n652 B.n434 256.663
R617 B.n654 B.n434 256.663
R618 B.n660 B.n434 256.663
R619 B.n662 B.n434 256.663
R620 B.n668 B.n434 256.663
R621 B.n670 B.n434 256.663
R622 B.n676 B.n434 256.663
R623 B.n678 B.n434 256.663
R624 B.n684 B.n434 256.663
R625 B.n686 B.n434 256.663
R626 B.n692 B.n434 256.663
R627 B.n694 B.n434 256.663
R628 B.n700 B.n434 256.663
R629 B.n702 B.n434 256.663
R630 B.n708 B.n434 256.663
R631 B.n710 B.n434 256.663
R632 B.n716 B.n434 256.663
R633 B.n718 B.n434 256.663
R634 B.n724 B.n434 256.663
R635 B.n726 B.n434 256.663
R636 B.n732 B.n434 256.663
R637 B.n734 B.n434 256.663
R638 B.n740 B.n434 256.663
R639 B.n742 B.n434 256.663
R640 B.n957 B.n956 256.663
R641 B.n132 B.n131 163.367
R642 B.n136 B.n135 163.367
R643 B.n140 B.n139 163.367
R644 B.n144 B.n143 163.367
R645 B.n148 B.n147 163.367
R646 B.n152 B.n151 163.367
R647 B.n156 B.n155 163.367
R648 B.n160 B.n159 163.367
R649 B.n164 B.n163 163.367
R650 B.n168 B.n167 163.367
R651 B.n172 B.n171 163.367
R652 B.n176 B.n175 163.367
R653 B.n180 B.n179 163.367
R654 B.n184 B.n183 163.367
R655 B.n188 B.n187 163.367
R656 B.n192 B.n191 163.367
R657 B.n196 B.n195 163.367
R658 B.n200 B.n199 163.367
R659 B.n204 B.n203 163.367
R660 B.n208 B.n207 163.367
R661 B.n212 B.n211 163.367
R662 B.n216 B.n215 163.367
R663 B.n220 B.n219 163.367
R664 B.n224 B.n223 163.367
R665 B.n228 B.n227 163.367
R666 B.n232 B.n231 163.367
R667 B.n236 B.n235 163.367
R668 B.n240 B.n239 163.367
R669 B.n245 B.n244 163.367
R670 B.n249 B.n248 163.367
R671 B.n253 B.n252 163.367
R672 B.n257 B.n256 163.367
R673 B.n261 B.n260 163.367
R674 B.n265 B.n264 163.367
R675 B.n269 B.n268 163.367
R676 B.n273 B.n272 163.367
R677 B.n277 B.n276 163.367
R678 B.n281 B.n280 163.367
R679 B.n285 B.n284 163.367
R680 B.n289 B.n288 163.367
R681 B.n293 B.n292 163.367
R682 B.n297 B.n296 163.367
R683 B.n301 B.n300 163.367
R684 B.n305 B.n304 163.367
R685 B.n309 B.n308 163.367
R686 B.n313 B.n312 163.367
R687 B.n317 B.n316 163.367
R688 B.n321 B.n320 163.367
R689 B.n325 B.n324 163.367
R690 B.n329 B.n328 163.367
R691 B.n333 B.n332 163.367
R692 B.n337 B.n336 163.367
R693 B.n341 B.n340 163.367
R694 B.n345 B.n344 163.367
R695 B.n349 B.n348 163.367
R696 B.n353 B.n352 163.367
R697 B.n357 B.n356 163.367
R698 B.n361 B.n360 163.367
R699 B.n365 B.n364 163.367
R700 B.n369 B.n368 163.367
R701 B.n887 B.n124 163.367
R702 B.n747 B.n429 163.367
R703 B.n755 B.n429 163.367
R704 B.n755 B.n427 163.367
R705 B.n759 B.n427 163.367
R706 B.n759 B.n420 163.367
R707 B.n767 B.n420 163.367
R708 B.n767 B.n418 163.367
R709 B.n771 B.n418 163.367
R710 B.n771 B.n413 163.367
R711 B.n779 B.n413 163.367
R712 B.n779 B.n411 163.367
R713 B.n783 B.n411 163.367
R714 B.n783 B.n405 163.367
R715 B.n791 B.n405 163.367
R716 B.n791 B.n403 163.367
R717 B.n795 B.n403 163.367
R718 B.n795 B.n397 163.367
R719 B.n803 B.n397 163.367
R720 B.n803 B.n395 163.367
R721 B.n807 B.n395 163.367
R722 B.n807 B.n389 163.367
R723 B.n815 B.n389 163.367
R724 B.n815 B.n387 163.367
R725 B.n819 B.n387 163.367
R726 B.n819 B.n381 163.367
R727 B.n827 B.n381 163.367
R728 B.n827 B.n379 163.367
R729 B.n832 B.n379 163.367
R730 B.n832 B.n373 163.367
R731 B.n840 B.n373 163.367
R732 B.n841 B.n840 163.367
R733 B.n841 B.n5 163.367
R734 B.n6 B.n5 163.367
R735 B.n7 B.n6 163.367
R736 B.n847 B.n7 163.367
R737 B.n848 B.n847 163.367
R738 B.n848 B.n13 163.367
R739 B.n14 B.n13 163.367
R740 B.n15 B.n14 163.367
R741 B.n853 B.n15 163.367
R742 B.n853 B.n20 163.367
R743 B.n21 B.n20 163.367
R744 B.n22 B.n21 163.367
R745 B.n858 B.n22 163.367
R746 B.n858 B.n27 163.367
R747 B.n28 B.n27 163.367
R748 B.n29 B.n28 163.367
R749 B.n863 B.n29 163.367
R750 B.n863 B.n34 163.367
R751 B.n35 B.n34 163.367
R752 B.n36 B.n35 163.367
R753 B.n868 B.n36 163.367
R754 B.n868 B.n41 163.367
R755 B.n42 B.n41 163.367
R756 B.n43 B.n42 163.367
R757 B.n873 B.n43 163.367
R758 B.n873 B.n48 163.367
R759 B.n49 B.n48 163.367
R760 B.n50 B.n49 163.367
R761 B.n878 B.n50 163.367
R762 B.n878 B.n55 163.367
R763 B.n56 B.n55 163.367
R764 B.n57 B.n56 163.367
R765 B.n883 B.n57 163.367
R766 B.n883 B.n62 163.367
R767 B.n502 B.n500 163.367
R768 B.n506 B.n500 163.367
R769 B.n510 B.n508 163.367
R770 B.n514 B.n498 163.367
R771 B.n518 B.n516 163.367
R772 B.n522 B.n496 163.367
R773 B.n526 B.n524 163.367
R774 B.n530 B.n494 163.367
R775 B.n534 B.n532 163.367
R776 B.n538 B.n492 163.367
R777 B.n542 B.n540 163.367
R778 B.n546 B.n490 163.367
R779 B.n550 B.n548 163.367
R780 B.n554 B.n488 163.367
R781 B.n558 B.n556 163.367
R782 B.n562 B.n486 163.367
R783 B.n566 B.n564 163.367
R784 B.n570 B.n484 163.367
R785 B.n574 B.n572 163.367
R786 B.n578 B.n482 163.367
R787 B.n582 B.n580 163.367
R788 B.n586 B.n480 163.367
R789 B.n590 B.n588 163.367
R790 B.n594 B.n478 163.367
R791 B.n598 B.n596 163.367
R792 B.n602 B.n476 163.367
R793 B.n606 B.n604 163.367
R794 B.n610 B.n474 163.367
R795 B.n614 B.n612 163.367
R796 B.n618 B.n469 163.367
R797 B.n622 B.n620 163.367
R798 B.n626 B.n467 163.367
R799 B.n630 B.n628 163.367
R800 B.n635 B.n463 163.367
R801 B.n639 B.n637 163.367
R802 B.n643 B.n461 163.367
R803 B.n647 B.n645 163.367
R804 B.n651 B.n459 163.367
R805 B.n655 B.n653 163.367
R806 B.n659 B.n457 163.367
R807 B.n663 B.n661 163.367
R808 B.n667 B.n455 163.367
R809 B.n671 B.n669 163.367
R810 B.n675 B.n453 163.367
R811 B.n679 B.n677 163.367
R812 B.n683 B.n451 163.367
R813 B.n687 B.n685 163.367
R814 B.n691 B.n449 163.367
R815 B.n695 B.n693 163.367
R816 B.n699 B.n447 163.367
R817 B.n703 B.n701 163.367
R818 B.n707 B.n445 163.367
R819 B.n711 B.n709 163.367
R820 B.n715 B.n443 163.367
R821 B.n719 B.n717 163.367
R822 B.n723 B.n441 163.367
R823 B.n727 B.n725 163.367
R824 B.n731 B.n439 163.367
R825 B.n735 B.n733 163.367
R826 B.n739 B.n437 163.367
R827 B.n743 B.n741 163.367
R828 B.n749 B.n431 163.367
R829 B.n753 B.n431 163.367
R830 B.n753 B.n425 163.367
R831 B.n761 B.n425 163.367
R832 B.n761 B.n423 163.367
R833 B.n765 B.n423 163.367
R834 B.n765 B.n417 163.367
R835 B.n773 B.n417 163.367
R836 B.n773 B.n415 163.367
R837 B.n777 B.n415 163.367
R838 B.n777 B.n409 163.367
R839 B.n785 B.n409 163.367
R840 B.n785 B.n407 163.367
R841 B.n789 B.n407 163.367
R842 B.n789 B.n401 163.367
R843 B.n797 B.n401 163.367
R844 B.n797 B.n399 163.367
R845 B.n801 B.n399 163.367
R846 B.n801 B.n393 163.367
R847 B.n809 B.n393 163.367
R848 B.n809 B.n391 163.367
R849 B.n813 B.n391 163.367
R850 B.n813 B.n385 163.367
R851 B.n821 B.n385 163.367
R852 B.n821 B.n383 163.367
R853 B.n825 B.n383 163.367
R854 B.n825 B.n377 163.367
R855 B.n834 B.n377 163.367
R856 B.n834 B.n375 163.367
R857 B.n838 B.n375 163.367
R858 B.n838 B.n3 163.367
R859 B.n955 B.n3 163.367
R860 B.n951 B.n2 163.367
R861 B.n951 B.n950 163.367
R862 B.n950 B.n9 163.367
R863 B.n946 B.n9 163.367
R864 B.n946 B.n11 163.367
R865 B.n942 B.n11 163.367
R866 B.n942 B.n17 163.367
R867 B.n938 B.n17 163.367
R868 B.n938 B.n19 163.367
R869 B.n934 B.n19 163.367
R870 B.n934 B.n24 163.367
R871 B.n930 B.n24 163.367
R872 B.n930 B.n26 163.367
R873 B.n926 B.n26 163.367
R874 B.n926 B.n31 163.367
R875 B.n922 B.n31 163.367
R876 B.n922 B.n33 163.367
R877 B.n918 B.n33 163.367
R878 B.n918 B.n38 163.367
R879 B.n914 B.n38 163.367
R880 B.n914 B.n40 163.367
R881 B.n910 B.n40 163.367
R882 B.n910 B.n45 163.367
R883 B.n906 B.n45 163.367
R884 B.n906 B.n47 163.367
R885 B.n902 B.n47 163.367
R886 B.n902 B.n52 163.367
R887 B.n898 B.n52 163.367
R888 B.n898 B.n54 163.367
R889 B.n894 B.n54 163.367
R890 B.n894 B.n59 163.367
R891 B.n890 B.n59 163.367
R892 B.n125 B.t6 123.933
R893 B.n464 B.t17 123.933
R894 B.n128 B.t9 123.909
R895 B.n470 B.t14 123.909
R896 B.n63 B.n61 71.676
R897 B.n132 B.n64 71.676
R898 B.n136 B.n65 71.676
R899 B.n140 B.n66 71.676
R900 B.n144 B.n67 71.676
R901 B.n148 B.n68 71.676
R902 B.n152 B.n69 71.676
R903 B.n156 B.n70 71.676
R904 B.n160 B.n71 71.676
R905 B.n164 B.n72 71.676
R906 B.n168 B.n73 71.676
R907 B.n172 B.n74 71.676
R908 B.n176 B.n75 71.676
R909 B.n180 B.n76 71.676
R910 B.n184 B.n77 71.676
R911 B.n188 B.n78 71.676
R912 B.n192 B.n79 71.676
R913 B.n196 B.n80 71.676
R914 B.n200 B.n81 71.676
R915 B.n204 B.n82 71.676
R916 B.n208 B.n83 71.676
R917 B.n212 B.n84 71.676
R918 B.n216 B.n85 71.676
R919 B.n220 B.n86 71.676
R920 B.n224 B.n87 71.676
R921 B.n228 B.n88 71.676
R922 B.n232 B.n89 71.676
R923 B.n236 B.n90 71.676
R924 B.n240 B.n91 71.676
R925 B.n245 B.n92 71.676
R926 B.n249 B.n93 71.676
R927 B.n253 B.n94 71.676
R928 B.n257 B.n95 71.676
R929 B.n261 B.n96 71.676
R930 B.n265 B.n97 71.676
R931 B.n269 B.n98 71.676
R932 B.n273 B.n99 71.676
R933 B.n277 B.n100 71.676
R934 B.n281 B.n101 71.676
R935 B.n285 B.n102 71.676
R936 B.n289 B.n103 71.676
R937 B.n293 B.n104 71.676
R938 B.n297 B.n105 71.676
R939 B.n301 B.n106 71.676
R940 B.n305 B.n107 71.676
R941 B.n309 B.n108 71.676
R942 B.n313 B.n109 71.676
R943 B.n317 B.n110 71.676
R944 B.n321 B.n111 71.676
R945 B.n325 B.n112 71.676
R946 B.n329 B.n113 71.676
R947 B.n333 B.n114 71.676
R948 B.n337 B.n115 71.676
R949 B.n341 B.n116 71.676
R950 B.n345 B.n117 71.676
R951 B.n349 B.n118 71.676
R952 B.n353 B.n119 71.676
R953 B.n357 B.n120 71.676
R954 B.n361 B.n121 71.676
R955 B.n365 B.n122 71.676
R956 B.n369 B.n123 71.676
R957 B.n124 B.n123 71.676
R958 B.n368 B.n122 71.676
R959 B.n364 B.n121 71.676
R960 B.n360 B.n120 71.676
R961 B.n356 B.n119 71.676
R962 B.n352 B.n118 71.676
R963 B.n348 B.n117 71.676
R964 B.n344 B.n116 71.676
R965 B.n340 B.n115 71.676
R966 B.n336 B.n114 71.676
R967 B.n332 B.n113 71.676
R968 B.n328 B.n112 71.676
R969 B.n324 B.n111 71.676
R970 B.n320 B.n110 71.676
R971 B.n316 B.n109 71.676
R972 B.n312 B.n108 71.676
R973 B.n308 B.n107 71.676
R974 B.n304 B.n106 71.676
R975 B.n300 B.n105 71.676
R976 B.n296 B.n104 71.676
R977 B.n292 B.n103 71.676
R978 B.n288 B.n102 71.676
R979 B.n284 B.n101 71.676
R980 B.n280 B.n100 71.676
R981 B.n276 B.n99 71.676
R982 B.n272 B.n98 71.676
R983 B.n268 B.n97 71.676
R984 B.n264 B.n96 71.676
R985 B.n260 B.n95 71.676
R986 B.n256 B.n94 71.676
R987 B.n252 B.n93 71.676
R988 B.n248 B.n92 71.676
R989 B.n244 B.n91 71.676
R990 B.n239 B.n90 71.676
R991 B.n235 B.n89 71.676
R992 B.n231 B.n88 71.676
R993 B.n227 B.n87 71.676
R994 B.n223 B.n86 71.676
R995 B.n219 B.n85 71.676
R996 B.n215 B.n84 71.676
R997 B.n211 B.n83 71.676
R998 B.n207 B.n82 71.676
R999 B.n203 B.n81 71.676
R1000 B.n199 B.n80 71.676
R1001 B.n195 B.n79 71.676
R1002 B.n191 B.n78 71.676
R1003 B.n187 B.n77 71.676
R1004 B.n183 B.n76 71.676
R1005 B.n179 B.n75 71.676
R1006 B.n175 B.n74 71.676
R1007 B.n171 B.n73 71.676
R1008 B.n167 B.n72 71.676
R1009 B.n163 B.n71 71.676
R1010 B.n159 B.n70 71.676
R1011 B.n155 B.n69 71.676
R1012 B.n151 B.n68 71.676
R1013 B.n147 B.n67 71.676
R1014 B.n143 B.n66 71.676
R1015 B.n139 B.n65 71.676
R1016 B.n135 B.n64 71.676
R1017 B.n131 B.n63 71.676
R1018 B.n501 B.n433 71.676
R1019 B.n507 B.n506 71.676
R1020 B.n510 B.n509 71.676
R1021 B.n515 B.n514 71.676
R1022 B.n518 B.n517 71.676
R1023 B.n523 B.n522 71.676
R1024 B.n526 B.n525 71.676
R1025 B.n531 B.n530 71.676
R1026 B.n534 B.n533 71.676
R1027 B.n539 B.n538 71.676
R1028 B.n542 B.n541 71.676
R1029 B.n547 B.n546 71.676
R1030 B.n550 B.n549 71.676
R1031 B.n555 B.n554 71.676
R1032 B.n558 B.n557 71.676
R1033 B.n563 B.n562 71.676
R1034 B.n566 B.n565 71.676
R1035 B.n571 B.n570 71.676
R1036 B.n574 B.n573 71.676
R1037 B.n579 B.n578 71.676
R1038 B.n582 B.n581 71.676
R1039 B.n587 B.n586 71.676
R1040 B.n590 B.n589 71.676
R1041 B.n595 B.n594 71.676
R1042 B.n598 B.n597 71.676
R1043 B.n603 B.n602 71.676
R1044 B.n606 B.n605 71.676
R1045 B.n611 B.n610 71.676
R1046 B.n614 B.n613 71.676
R1047 B.n619 B.n618 71.676
R1048 B.n622 B.n621 71.676
R1049 B.n627 B.n626 71.676
R1050 B.n630 B.n629 71.676
R1051 B.n636 B.n635 71.676
R1052 B.n639 B.n638 71.676
R1053 B.n644 B.n643 71.676
R1054 B.n647 B.n646 71.676
R1055 B.n652 B.n651 71.676
R1056 B.n655 B.n654 71.676
R1057 B.n660 B.n659 71.676
R1058 B.n663 B.n662 71.676
R1059 B.n668 B.n667 71.676
R1060 B.n671 B.n670 71.676
R1061 B.n676 B.n675 71.676
R1062 B.n679 B.n678 71.676
R1063 B.n684 B.n683 71.676
R1064 B.n687 B.n686 71.676
R1065 B.n692 B.n691 71.676
R1066 B.n695 B.n694 71.676
R1067 B.n700 B.n699 71.676
R1068 B.n703 B.n702 71.676
R1069 B.n708 B.n707 71.676
R1070 B.n711 B.n710 71.676
R1071 B.n716 B.n715 71.676
R1072 B.n719 B.n718 71.676
R1073 B.n724 B.n723 71.676
R1074 B.n727 B.n726 71.676
R1075 B.n732 B.n731 71.676
R1076 B.n735 B.n734 71.676
R1077 B.n740 B.n739 71.676
R1078 B.n743 B.n742 71.676
R1079 B.n502 B.n501 71.676
R1080 B.n508 B.n507 71.676
R1081 B.n509 B.n498 71.676
R1082 B.n516 B.n515 71.676
R1083 B.n517 B.n496 71.676
R1084 B.n524 B.n523 71.676
R1085 B.n525 B.n494 71.676
R1086 B.n532 B.n531 71.676
R1087 B.n533 B.n492 71.676
R1088 B.n540 B.n539 71.676
R1089 B.n541 B.n490 71.676
R1090 B.n548 B.n547 71.676
R1091 B.n549 B.n488 71.676
R1092 B.n556 B.n555 71.676
R1093 B.n557 B.n486 71.676
R1094 B.n564 B.n563 71.676
R1095 B.n565 B.n484 71.676
R1096 B.n572 B.n571 71.676
R1097 B.n573 B.n482 71.676
R1098 B.n580 B.n579 71.676
R1099 B.n581 B.n480 71.676
R1100 B.n588 B.n587 71.676
R1101 B.n589 B.n478 71.676
R1102 B.n596 B.n595 71.676
R1103 B.n597 B.n476 71.676
R1104 B.n604 B.n603 71.676
R1105 B.n605 B.n474 71.676
R1106 B.n612 B.n611 71.676
R1107 B.n613 B.n469 71.676
R1108 B.n620 B.n619 71.676
R1109 B.n621 B.n467 71.676
R1110 B.n628 B.n627 71.676
R1111 B.n629 B.n463 71.676
R1112 B.n637 B.n636 71.676
R1113 B.n638 B.n461 71.676
R1114 B.n645 B.n644 71.676
R1115 B.n646 B.n459 71.676
R1116 B.n653 B.n652 71.676
R1117 B.n654 B.n457 71.676
R1118 B.n661 B.n660 71.676
R1119 B.n662 B.n455 71.676
R1120 B.n669 B.n668 71.676
R1121 B.n670 B.n453 71.676
R1122 B.n677 B.n676 71.676
R1123 B.n678 B.n451 71.676
R1124 B.n685 B.n684 71.676
R1125 B.n686 B.n449 71.676
R1126 B.n693 B.n692 71.676
R1127 B.n694 B.n447 71.676
R1128 B.n701 B.n700 71.676
R1129 B.n702 B.n445 71.676
R1130 B.n709 B.n708 71.676
R1131 B.n710 B.n443 71.676
R1132 B.n717 B.n716 71.676
R1133 B.n718 B.n441 71.676
R1134 B.n725 B.n724 71.676
R1135 B.n726 B.n439 71.676
R1136 B.n733 B.n732 71.676
R1137 B.n734 B.n437 71.676
R1138 B.n741 B.n740 71.676
R1139 B.n742 B.n435 71.676
R1140 B.n956 B.n955 71.676
R1141 B.n956 B.n2 71.676
R1142 B.n126 B.t7 70.211
R1143 B.n465 B.t16 70.211
R1144 B.n129 B.t10 70.1883
R1145 B.n471 B.t13 70.1883
R1146 B.n748 B.n434 62.297
R1147 B.n889 B.n888 62.297
R1148 B.n242 B.n129 59.5399
R1149 B.n127 B.n126 59.5399
R1150 B.n632 B.n465 59.5399
R1151 B.n472 B.n471 59.5399
R1152 B.n129 B.n128 53.7217
R1153 B.n126 B.n125 53.7217
R1154 B.n465 B.n464 53.7217
R1155 B.n471 B.n470 53.7217
R1156 B.n750 B.n432 33.5615
R1157 B.n746 B.n745 33.5615
R1158 B.n886 B.n885 33.5615
R1159 B.n891 B.n60 33.5615
R1160 B.n748 B.n430 33.3561
R1161 B.n754 B.n430 33.3561
R1162 B.n754 B.n426 33.3561
R1163 B.n760 B.n426 33.3561
R1164 B.n760 B.n421 33.3561
R1165 B.n766 B.n421 33.3561
R1166 B.n766 B.n422 33.3561
R1167 B.n772 B.n414 33.3561
R1168 B.n778 B.n414 33.3561
R1169 B.n778 B.n410 33.3561
R1170 B.n784 B.n410 33.3561
R1171 B.n784 B.n406 33.3561
R1172 B.n790 B.n406 33.3561
R1173 B.n790 B.n402 33.3561
R1174 B.n796 B.n402 33.3561
R1175 B.n796 B.n398 33.3561
R1176 B.n802 B.n398 33.3561
R1177 B.n808 B.n394 33.3561
R1178 B.n808 B.n390 33.3561
R1179 B.n814 B.n390 33.3561
R1180 B.n814 B.n386 33.3561
R1181 B.n820 B.n386 33.3561
R1182 B.n820 B.n382 33.3561
R1183 B.n826 B.n382 33.3561
R1184 B.n833 B.n378 33.3561
R1185 B.n833 B.n374 33.3561
R1186 B.n839 B.n374 33.3561
R1187 B.n839 B.n4 33.3561
R1188 B.n954 B.n4 33.3561
R1189 B.n954 B.n953 33.3561
R1190 B.n953 B.n952 33.3561
R1191 B.n952 B.n8 33.3561
R1192 B.n12 B.n8 33.3561
R1193 B.n945 B.n12 33.3561
R1194 B.n945 B.n944 33.3561
R1195 B.n943 B.n16 33.3561
R1196 B.n937 B.n16 33.3561
R1197 B.n937 B.n936 33.3561
R1198 B.n936 B.n935 33.3561
R1199 B.n935 B.n23 33.3561
R1200 B.n929 B.n23 33.3561
R1201 B.n929 B.n928 33.3561
R1202 B.n927 B.n30 33.3561
R1203 B.n921 B.n30 33.3561
R1204 B.n921 B.n920 33.3561
R1205 B.n920 B.n919 33.3561
R1206 B.n919 B.n37 33.3561
R1207 B.n913 B.n37 33.3561
R1208 B.n913 B.n912 33.3561
R1209 B.n912 B.n911 33.3561
R1210 B.n911 B.n44 33.3561
R1211 B.n905 B.n44 33.3561
R1212 B.n904 B.n903 33.3561
R1213 B.n903 B.n51 33.3561
R1214 B.n897 B.n51 33.3561
R1215 B.n897 B.n896 33.3561
R1216 B.n896 B.n895 33.3561
R1217 B.n895 B.n58 33.3561
R1218 B.n889 B.n58 33.3561
R1219 B.n826 B.t3 27.4698
R1220 B.t2 B.n943 27.4698
R1221 B.n772 B.t12 22.5646
R1222 B.n802 B.t1 22.5646
R1223 B.t0 B.n927 22.5646
R1224 B.n905 B.t5 22.5646
R1225 B B.n957 18.0485
R1226 B.n422 B.t12 10.792
R1227 B.t1 B.n394 10.792
R1228 B.n928 B.t0 10.792
R1229 B.t5 B.n904 10.792
R1230 B.n751 B.n750 10.6151
R1231 B.n752 B.n751 10.6151
R1232 B.n752 B.n424 10.6151
R1233 B.n762 B.n424 10.6151
R1234 B.n763 B.n762 10.6151
R1235 B.n764 B.n763 10.6151
R1236 B.n764 B.n416 10.6151
R1237 B.n774 B.n416 10.6151
R1238 B.n775 B.n774 10.6151
R1239 B.n776 B.n775 10.6151
R1240 B.n776 B.n408 10.6151
R1241 B.n786 B.n408 10.6151
R1242 B.n787 B.n786 10.6151
R1243 B.n788 B.n787 10.6151
R1244 B.n788 B.n400 10.6151
R1245 B.n798 B.n400 10.6151
R1246 B.n799 B.n798 10.6151
R1247 B.n800 B.n799 10.6151
R1248 B.n800 B.n392 10.6151
R1249 B.n810 B.n392 10.6151
R1250 B.n811 B.n810 10.6151
R1251 B.n812 B.n811 10.6151
R1252 B.n812 B.n384 10.6151
R1253 B.n822 B.n384 10.6151
R1254 B.n823 B.n822 10.6151
R1255 B.n824 B.n823 10.6151
R1256 B.n824 B.n376 10.6151
R1257 B.n835 B.n376 10.6151
R1258 B.n836 B.n835 10.6151
R1259 B.n837 B.n836 10.6151
R1260 B.n837 B.n0 10.6151
R1261 B.n503 B.n432 10.6151
R1262 B.n504 B.n503 10.6151
R1263 B.n505 B.n504 10.6151
R1264 B.n505 B.n499 10.6151
R1265 B.n511 B.n499 10.6151
R1266 B.n512 B.n511 10.6151
R1267 B.n513 B.n512 10.6151
R1268 B.n513 B.n497 10.6151
R1269 B.n519 B.n497 10.6151
R1270 B.n520 B.n519 10.6151
R1271 B.n521 B.n520 10.6151
R1272 B.n521 B.n495 10.6151
R1273 B.n527 B.n495 10.6151
R1274 B.n528 B.n527 10.6151
R1275 B.n529 B.n528 10.6151
R1276 B.n529 B.n493 10.6151
R1277 B.n535 B.n493 10.6151
R1278 B.n536 B.n535 10.6151
R1279 B.n537 B.n536 10.6151
R1280 B.n537 B.n491 10.6151
R1281 B.n543 B.n491 10.6151
R1282 B.n544 B.n543 10.6151
R1283 B.n545 B.n544 10.6151
R1284 B.n545 B.n489 10.6151
R1285 B.n551 B.n489 10.6151
R1286 B.n552 B.n551 10.6151
R1287 B.n553 B.n552 10.6151
R1288 B.n553 B.n487 10.6151
R1289 B.n559 B.n487 10.6151
R1290 B.n560 B.n559 10.6151
R1291 B.n561 B.n560 10.6151
R1292 B.n561 B.n485 10.6151
R1293 B.n567 B.n485 10.6151
R1294 B.n568 B.n567 10.6151
R1295 B.n569 B.n568 10.6151
R1296 B.n569 B.n483 10.6151
R1297 B.n575 B.n483 10.6151
R1298 B.n576 B.n575 10.6151
R1299 B.n577 B.n576 10.6151
R1300 B.n577 B.n481 10.6151
R1301 B.n583 B.n481 10.6151
R1302 B.n584 B.n583 10.6151
R1303 B.n585 B.n584 10.6151
R1304 B.n585 B.n479 10.6151
R1305 B.n591 B.n479 10.6151
R1306 B.n592 B.n591 10.6151
R1307 B.n593 B.n592 10.6151
R1308 B.n593 B.n477 10.6151
R1309 B.n599 B.n477 10.6151
R1310 B.n600 B.n599 10.6151
R1311 B.n601 B.n600 10.6151
R1312 B.n601 B.n475 10.6151
R1313 B.n607 B.n475 10.6151
R1314 B.n608 B.n607 10.6151
R1315 B.n609 B.n608 10.6151
R1316 B.n609 B.n473 10.6151
R1317 B.n616 B.n615 10.6151
R1318 B.n617 B.n616 10.6151
R1319 B.n617 B.n468 10.6151
R1320 B.n623 B.n468 10.6151
R1321 B.n624 B.n623 10.6151
R1322 B.n625 B.n624 10.6151
R1323 B.n625 B.n466 10.6151
R1324 B.n631 B.n466 10.6151
R1325 B.n634 B.n633 10.6151
R1326 B.n634 B.n462 10.6151
R1327 B.n640 B.n462 10.6151
R1328 B.n641 B.n640 10.6151
R1329 B.n642 B.n641 10.6151
R1330 B.n642 B.n460 10.6151
R1331 B.n648 B.n460 10.6151
R1332 B.n649 B.n648 10.6151
R1333 B.n650 B.n649 10.6151
R1334 B.n650 B.n458 10.6151
R1335 B.n656 B.n458 10.6151
R1336 B.n657 B.n656 10.6151
R1337 B.n658 B.n657 10.6151
R1338 B.n658 B.n456 10.6151
R1339 B.n664 B.n456 10.6151
R1340 B.n665 B.n664 10.6151
R1341 B.n666 B.n665 10.6151
R1342 B.n666 B.n454 10.6151
R1343 B.n672 B.n454 10.6151
R1344 B.n673 B.n672 10.6151
R1345 B.n674 B.n673 10.6151
R1346 B.n674 B.n452 10.6151
R1347 B.n680 B.n452 10.6151
R1348 B.n681 B.n680 10.6151
R1349 B.n682 B.n681 10.6151
R1350 B.n682 B.n450 10.6151
R1351 B.n688 B.n450 10.6151
R1352 B.n689 B.n688 10.6151
R1353 B.n690 B.n689 10.6151
R1354 B.n690 B.n448 10.6151
R1355 B.n696 B.n448 10.6151
R1356 B.n697 B.n696 10.6151
R1357 B.n698 B.n697 10.6151
R1358 B.n698 B.n446 10.6151
R1359 B.n704 B.n446 10.6151
R1360 B.n705 B.n704 10.6151
R1361 B.n706 B.n705 10.6151
R1362 B.n706 B.n444 10.6151
R1363 B.n712 B.n444 10.6151
R1364 B.n713 B.n712 10.6151
R1365 B.n714 B.n713 10.6151
R1366 B.n714 B.n442 10.6151
R1367 B.n720 B.n442 10.6151
R1368 B.n721 B.n720 10.6151
R1369 B.n722 B.n721 10.6151
R1370 B.n722 B.n440 10.6151
R1371 B.n728 B.n440 10.6151
R1372 B.n729 B.n728 10.6151
R1373 B.n730 B.n729 10.6151
R1374 B.n730 B.n438 10.6151
R1375 B.n736 B.n438 10.6151
R1376 B.n737 B.n736 10.6151
R1377 B.n738 B.n737 10.6151
R1378 B.n738 B.n436 10.6151
R1379 B.n744 B.n436 10.6151
R1380 B.n745 B.n744 10.6151
R1381 B.n746 B.n428 10.6151
R1382 B.n756 B.n428 10.6151
R1383 B.n757 B.n756 10.6151
R1384 B.n758 B.n757 10.6151
R1385 B.n758 B.n419 10.6151
R1386 B.n768 B.n419 10.6151
R1387 B.n769 B.n768 10.6151
R1388 B.n770 B.n769 10.6151
R1389 B.n770 B.n412 10.6151
R1390 B.n780 B.n412 10.6151
R1391 B.n781 B.n780 10.6151
R1392 B.n782 B.n781 10.6151
R1393 B.n782 B.n404 10.6151
R1394 B.n792 B.n404 10.6151
R1395 B.n793 B.n792 10.6151
R1396 B.n794 B.n793 10.6151
R1397 B.n794 B.n396 10.6151
R1398 B.n804 B.n396 10.6151
R1399 B.n805 B.n804 10.6151
R1400 B.n806 B.n805 10.6151
R1401 B.n806 B.n388 10.6151
R1402 B.n816 B.n388 10.6151
R1403 B.n817 B.n816 10.6151
R1404 B.n818 B.n817 10.6151
R1405 B.n818 B.n380 10.6151
R1406 B.n828 B.n380 10.6151
R1407 B.n829 B.n828 10.6151
R1408 B.n831 B.n829 10.6151
R1409 B.n831 B.n830 10.6151
R1410 B.n830 B.n372 10.6151
R1411 B.n842 B.n372 10.6151
R1412 B.n843 B.n842 10.6151
R1413 B.n844 B.n843 10.6151
R1414 B.n845 B.n844 10.6151
R1415 B.n846 B.n845 10.6151
R1416 B.n849 B.n846 10.6151
R1417 B.n850 B.n849 10.6151
R1418 B.n851 B.n850 10.6151
R1419 B.n852 B.n851 10.6151
R1420 B.n854 B.n852 10.6151
R1421 B.n855 B.n854 10.6151
R1422 B.n856 B.n855 10.6151
R1423 B.n857 B.n856 10.6151
R1424 B.n859 B.n857 10.6151
R1425 B.n860 B.n859 10.6151
R1426 B.n861 B.n860 10.6151
R1427 B.n862 B.n861 10.6151
R1428 B.n864 B.n862 10.6151
R1429 B.n865 B.n864 10.6151
R1430 B.n866 B.n865 10.6151
R1431 B.n867 B.n866 10.6151
R1432 B.n869 B.n867 10.6151
R1433 B.n870 B.n869 10.6151
R1434 B.n871 B.n870 10.6151
R1435 B.n872 B.n871 10.6151
R1436 B.n874 B.n872 10.6151
R1437 B.n875 B.n874 10.6151
R1438 B.n876 B.n875 10.6151
R1439 B.n877 B.n876 10.6151
R1440 B.n879 B.n877 10.6151
R1441 B.n880 B.n879 10.6151
R1442 B.n881 B.n880 10.6151
R1443 B.n882 B.n881 10.6151
R1444 B.n884 B.n882 10.6151
R1445 B.n885 B.n884 10.6151
R1446 B.n949 B.n1 10.6151
R1447 B.n949 B.n948 10.6151
R1448 B.n948 B.n947 10.6151
R1449 B.n947 B.n10 10.6151
R1450 B.n941 B.n10 10.6151
R1451 B.n941 B.n940 10.6151
R1452 B.n940 B.n939 10.6151
R1453 B.n939 B.n18 10.6151
R1454 B.n933 B.n18 10.6151
R1455 B.n933 B.n932 10.6151
R1456 B.n932 B.n931 10.6151
R1457 B.n931 B.n25 10.6151
R1458 B.n925 B.n25 10.6151
R1459 B.n925 B.n924 10.6151
R1460 B.n924 B.n923 10.6151
R1461 B.n923 B.n32 10.6151
R1462 B.n917 B.n32 10.6151
R1463 B.n917 B.n916 10.6151
R1464 B.n916 B.n915 10.6151
R1465 B.n915 B.n39 10.6151
R1466 B.n909 B.n39 10.6151
R1467 B.n909 B.n908 10.6151
R1468 B.n908 B.n907 10.6151
R1469 B.n907 B.n46 10.6151
R1470 B.n901 B.n46 10.6151
R1471 B.n901 B.n900 10.6151
R1472 B.n900 B.n899 10.6151
R1473 B.n899 B.n53 10.6151
R1474 B.n893 B.n53 10.6151
R1475 B.n893 B.n892 10.6151
R1476 B.n892 B.n891 10.6151
R1477 B.n130 B.n60 10.6151
R1478 B.n133 B.n130 10.6151
R1479 B.n134 B.n133 10.6151
R1480 B.n137 B.n134 10.6151
R1481 B.n138 B.n137 10.6151
R1482 B.n141 B.n138 10.6151
R1483 B.n142 B.n141 10.6151
R1484 B.n145 B.n142 10.6151
R1485 B.n146 B.n145 10.6151
R1486 B.n149 B.n146 10.6151
R1487 B.n150 B.n149 10.6151
R1488 B.n153 B.n150 10.6151
R1489 B.n154 B.n153 10.6151
R1490 B.n157 B.n154 10.6151
R1491 B.n158 B.n157 10.6151
R1492 B.n161 B.n158 10.6151
R1493 B.n162 B.n161 10.6151
R1494 B.n165 B.n162 10.6151
R1495 B.n166 B.n165 10.6151
R1496 B.n169 B.n166 10.6151
R1497 B.n170 B.n169 10.6151
R1498 B.n173 B.n170 10.6151
R1499 B.n174 B.n173 10.6151
R1500 B.n177 B.n174 10.6151
R1501 B.n178 B.n177 10.6151
R1502 B.n181 B.n178 10.6151
R1503 B.n182 B.n181 10.6151
R1504 B.n185 B.n182 10.6151
R1505 B.n186 B.n185 10.6151
R1506 B.n189 B.n186 10.6151
R1507 B.n190 B.n189 10.6151
R1508 B.n193 B.n190 10.6151
R1509 B.n194 B.n193 10.6151
R1510 B.n197 B.n194 10.6151
R1511 B.n198 B.n197 10.6151
R1512 B.n201 B.n198 10.6151
R1513 B.n202 B.n201 10.6151
R1514 B.n205 B.n202 10.6151
R1515 B.n206 B.n205 10.6151
R1516 B.n209 B.n206 10.6151
R1517 B.n210 B.n209 10.6151
R1518 B.n213 B.n210 10.6151
R1519 B.n214 B.n213 10.6151
R1520 B.n217 B.n214 10.6151
R1521 B.n218 B.n217 10.6151
R1522 B.n221 B.n218 10.6151
R1523 B.n222 B.n221 10.6151
R1524 B.n225 B.n222 10.6151
R1525 B.n226 B.n225 10.6151
R1526 B.n229 B.n226 10.6151
R1527 B.n230 B.n229 10.6151
R1528 B.n233 B.n230 10.6151
R1529 B.n234 B.n233 10.6151
R1530 B.n237 B.n234 10.6151
R1531 B.n238 B.n237 10.6151
R1532 B.n241 B.n238 10.6151
R1533 B.n246 B.n243 10.6151
R1534 B.n247 B.n246 10.6151
R1535 B.n250 B.n247 10.6151
R1536 B.n251 B.n250 10.6151
R1537 B.n254 B.n251 10.6151
R1538 B.n255 B.n254 10.6151
R1539 B.n258 B.n255 10.6151
R1540 B.n259 B.n258 10.6151
R1541 B.n263 B.n262 10.6151
R1542 B.n266 B.n263 10.6151
R1543 B.n267 B.n266 10.6151
R1544 B.n270 B.n267 10.6151
R1545 B.n271 B.n270 10.6151
R1546 B.n274 B.n271 10.6151
R1547 B.n275 B.n274 10.6151
R1548 B.n278 B.n275 10.6151
R1549 B.n279 B.n278 10.6151
R1550 B.n282 B.n279 10.6151
R1551 B.n283 B.n282 10.6151
R1552 B.n286 B.n283 10.6151
R1553 B.n287 B.n286 10.6151
R1554 B.n290 B.n287 10.6151
R1555 B.n291 B.n290 10.6151
R1556 B.n294 B.n291 10.6151
R1557 B.n295 B.n294 10.6151
R1558 B.n298 B.n295 10.6151
R1559 B.n299 B.n298 10.6151
R1560 B.n302 B.n299 10.6151
R1561 B.n303 B.n302 10.6151
R1562 B.n306 B.n303 10.6151
R1563 B.n307 B.n306 10.6151
R1564 B.n310 B.n307 10.6151
R1565 B.n311 B.n310 10.6151
R1566 B.n314 B.n311 10.6151
R1567 B.n315 B.n314 10.6151
R1568 B.n318 B.n315 10.6151
R1569 B.n319 B.n318 10.6151
R1570 B.n322 B.n319 10.6151
R1571 B.n323 B.n322 10.6151
R1572 B.n326 B.n323 10.6151
R1573 B.n327 B.n326 10.6151
R1574 B.n330 B.n327 10.6151
R1575 B.n331 B.n330 10.6151
R1576 B.n334 B.n331 10.6151
R1577 B.n335 B.n334 10.6151
R1578 B.n338 B.n335 10.6151
R1579 B.n339 B.n338 10.6151
R1580 B.n342 B.n339 10.6151
R1581 B.n343 B.n342 10.6151
R1582 B.n346 B.n343 10.6151
R1583 B.n347 B.n346 10.6151
R1584 B.n350 B.n347 10.6151
R1585 B.n351 B.n350 10.6151
R1586 B.n354 B.n351 10.6151
R1587 B.n355 B.n354 10.6151
R1588 B.n358 B.n355 10.6151
R1589 B.n359 B.n358 10.6151
R1590 B.n362 B.n359 10.6151
R1591 B.n363 B.n362 10.6151
R1592 B.n366 B.n363 10.6151
R1593 B.n367 B.n366 10.6151
R1594 B.n370 B.n367 10.6151
R1595 B.n371 B.n370 10.6151
R1596 B.n886 B.n371 10.6151
R1597 B.n957 B.n0 8.11757
R1598 B.n957 B.n1 8.11757
R1599 B.n615 B.n472 6.5566
R1600 B.n632 B.n631 6.5566
R1601 B.n243 B.n242 6.5566
R1602 B.n259 B.n127 6.5566
R1603 B.t3 B.n378 5.88679
R1604 B.n944 B.t2 5.88679
R1605 B.n473 B.n472 4.05904
R1606 B.n633 B.n632 4.05904
R1607 B.n242 B.n241 4.05904
R1608 B.n262 B.n127 4.05904
R1609 VN.n0 VN.t2 204.322
R1610 VN.n1 VN.t3 204.322
R1611 VN.n0 VN.t0 203.576
R1612 VN.n1 VN.t1 203.576
R1613 VN VN.n1 54.5548
R1614 VN VN.n0 4.64949
R1615 VTAIL.n5 VTAIL.t2 44.9838
R1616 VTAIL.n4 VTAIL.t6 44.9838
R1617 VTAIL.n3 VTAIL.t5 44.9838
R1618 VTAIL.n7 VTAIL.t7 44.9837
R1619 VTAIL.n0 VTAIL.t4 44.9837
R1620 VTAIL.n1 VTAIL.t3 44.9837
R1621 VTAIL.n2 VTAIL.t1 44.9837
R1622 VTAIL.n6 VTAIL.t0 44.9837
R1623 VTAIL.n7 VTAIL.n6 29.5393
R1624 VTAIL.n3 VTAIL.n2 29.5393
R1625 VTAIL.n4 VTAIL.n3 2.38843
R1626 VTAIL.n6 VTAIL.n5 2.38843
R1627 VTAIL.n2 VTAIL.n1 2.38843
R1628 VTAIL VTAIL.n0 1.25266
R1629 VTAIL VTAIL.n7 1.13628
R1630 VTAIL.n5 VTAIL.n4 0.470328
R1631 VTAIL.n1 VTAIL.n0 0.470328
R1632 VDD2.n2 VDD2.n0 106.171
R1633 VDD2.n2 VDD2.n1 60.5079
R1634 VDD2.n1 VDD2.t2 1.15502
R1635 VDD2.n1 VDD2.t0 1.15502
R1636 VDD2.n0 VDD2.t1 1.15502
R1637 VDD2.n0 VDD2.t3 1.15502
R1638 VDD2 VDD2.n2 0.0586897
R1639 VP.n4 VP.t3 204.322
R1640 VP.n4 VP.t1 203.576
R1641 VP.n3 VP.t2 169.392
R1642 VP.n15 VP.t0 169.392
R1643 VP.n14 VP.n0 161.3
R1644 VP.n13 VP.n12 161.3
R1645 VP.n11 VP.n1 161.3
R1646 VP.n10 VP.n9 161.3
R1647 VP.n8 VP.n2 161.3
R1648 VP.n7 VP.n6 161.3
R1649 VP.n5 VP.n3 104.15
R1650 VP.n16 VP.n15 104.15
R1651 VP.n9 VP.n1 56.5193
R1652 VP.n5 VP.n4 54.2759
R1653 VP.n8 VP.n7 24.4675
R1654 VP.n9 VP.n8 24.4675
R1655 VP.n13 VP.n1 24.4675
R1656 VP.n14 VP.n13 24.4675
R1657 VP.n7 VP.n3 6.60659
R1658 VP.n15 VP.n14 6.60659
R1659 VP.n6 VP.n5 0.278367
R1660 VP.n16 VP.n0 0.278367
R1661 VP.n6 VP.n2 0.189894
R1662 VP.n10 VP.n2 0.189894
R1663 VP.n11 VP.n10 0.189894
R1664 VP.n12 VP.n11 0.189894
R1665 VP.n12 VP.n0 0.189894
R1666 VP VP.n16 0.153454
R1667 VDD1 VDD1.n1 106.695
R1668 VDD1 VDD1.n0 60.5661
R1669 VDD1.n0 VDD1.t0 1.15502
R1670 VDD1.n0 VDD1.t2 1.15502
R1671 VDD1.n1 VDD1.t1 1.15502
R1672 VDD1.n1 VDD1.t3 1.15502
C0 VP VTAIL 6.25101f
C1 VDD2 VTAIL 6.69478f
C2 VN VTAIL 6.23691f
C3 VDD1 VP 6.80712f
C4 VDD1 VDD2 0.99445f
C5 VDD1 VN 0.148988f
C6 VP VDD2 0.384257f
C7 VP VN 7.03286f
C8 VDD2 VN 6.57255f
C9 VDD1 VTAIL 6.64165f
C10 VDD2 B 4.072531f
C11 VDD1 B 8.655139f
C12 VTAIL B 13.071259f
C13 VN B 10.843639f
C14 VP B 8.947468f
C15 VDD1.t0 B 0.360104f
C16 VDD1.t2 B 0.360104f
C17 VDD1.n0 B 3.27405f
C18 VDD1.t1 B 0.360104f
C19 VDD1.t3 B 0.360104f
C20 VDD1.n1 B 4.15894f
C21 VP.n0 B 0.03398f
C22 VP.t0 B 2.96377f
C23 VP.n1 B 0.037625f
C24 VP.n2 B 0.025774f
C25 VP.t2 B 2.96377f
C26 VP.n3 B 1.10743f
C27 VP.t1 B 3.16272f
C28 VP.t3 B 3.16703f
C29 VP.n4 B 3.5744f
C30 VP.n5 B 1.57955f
C31 VP.n6 B 0.03398f
C32 VP.n7 B 0.030722f
C33 VP.n8 B 0.048035f
C34 VP.n9 B 0.037625f
C35 VP.n10 B 0.025774f
C36 VP.n11 B 0.025774f
C37 VP.n12 B 0.025774f
C38 VP.n13 B 0.048035f
C39 VP.n14 B 0.030722f
C40 VP.n15 B 1.10743f
C41 VP.n16 B 0.042574f
C42 VDD2.t1 B 0.360053f
C43 VDD2.t3 B 0.360053f
C44 VDD2.n0 B 4.13009f
C45 VDD2.t2 B 0.360053f
C46 VDD2.t0 B 0.360053f
C47 VDD2.n1 B 3.27317f
C48 VDD2.n2 B 4.24638f
C49 VTAIL.t4 B 2.3556f
C50 VTAIL.n0 B 0.295661f
C51 VTAIL.t3 B 2.3556f
C52 VTAIL.n1 B 0.351861f
C53 VTAIL.t1 B 2.3556f
C54 VTAIL.n2 B 1.38693f
C55 VTAIL.t5 B 2.35562f
C56 VTAIL.n3 B 1.38692f
C57 VTAIL.t6 B 2.35562f
C58 VTAIL.n4 B 0.351846f
C59 VTAIL.t2 B 2.35562f
C60 VTAIL.n5 B 0.351846f
C61 VTAIL.t0 B 2.3556f
C62 VTAIL.n6 B 1.38693f
C63 VTAIL.t7 B 2.3556f
C64 VTAIL.n7 B 1.32497f
C65 VN.t2 B 3.11415f
C66 VN.t0 B 3.10991f
C67 VN.n0 B 2.0367f
C68 VN.t3 B 3.11415f
C69 VN.t1 B 3.10991f
C70 VN.n1 B 3.5279f
.ends

