* NGSPICE file created from diff_pair_sample_1265.ext - technology: sky130A

.subckt diff_pair_sample_1265 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t11 w_n4570_n3366# sky130_fd_pr__pfet_01v8 ad=1.97835 pd=12.32 as=4.6761 ps=24.76 w=11.99 l=3.27
X1 VDD2.t7 VN.t0 VTAIL.t1 w_n4570_n3366# sky130_fd_pr__pfet_01v8 ad=1.97835 pd=12.32 as=4.6761 ps=24.76 w=11.99 l=3.27
X2 VDD2.t6 VN.t1 VTAIL.t2 w_n4570_n3366# sky130_fd_pr__pfet_01v8 ad=1.97835 pd=12.32 as=1.97835 ps=12.32 w=11.99 l=3.27
X3 VTAIL.t3 VN.t2 VDD2.t5 w_n4570_n3366# sky130_fd_pr__pfet_01v8 ad=1.97835 pd=12.32 as=1.97835 ps=12.32 w=11.99 l=3.27
X4 VTAIL.t4 VN.t3 VDD2.t4 w_n4570_n3366# sky130_fd_pr__pfet_01v8 ad=4.6761 pd=24.76 as=1.97835 ps=12.32 w=11.99 l=3.27
X5 B.t11 B.t9 B.t10 w_n4570_n3366# sky130_fd_pr__pfet_01v8 ad=4.6761 pd=24.76 as=0 ps=0 w=11.99 l=3.27
X6 B.t8 B.t6 B.t7 w_n4570_n3366# sky130_fd_pr__pfet_01v8 ad=4.6761 pd=24.76 as=0 ps=0 w=11.99 l=3.27
X7 VDD2.t3 VN.t4 VTAIL.t0 w_n4570_n3366# sky130_fd_pr__pfet_01v8 ad=1.97835 pd=12.32 as=4.6761 ps=24.76 w=11.99 l=3.27
X8 VDD2.t2 VN.t5 VTAIL.t6 w_n4570_n3366# sky130_fd_pr__pfet_01v8 ad=1.97835 pd=12.32 as=1.97835 ps=12.32 w=11.99 l=3.27
X9 VDD1.t6 VP.t1 VTAIL.t8 w_n4570_n3366# sky130_fd_pr__pfet_01v8 ad=1.97835 pd=12.32 as=1.97835 ps=12.32 w=11.99 l=3.27
X10 VDD1.t5 VP.t2 VTAIL.t12 w_n4570_n3366# sky130_fd_pr__pfet_01v8 ad=1.97835 pd=12.32 as=1.97835 ps=12.32 w=11.99 l=3.27
X11 VTAIL.t10 VP.t3 VDD1.t4 w_n4570_n3366# sky130_fd_pr__pfet_01v8 ad=1.97835 pd=12.32 as=1.97835 ps=12.32 w=11.99 l=3.27
X12 VTAIL.t9 VP.t4 VDD1.t3 w_n4570_n3366# sky130_fd_pr__pfet_01v8 ad=4.6761 pd=24.76 as=1.97835 ps=12.32 w=11.99 l=3.27
X13 VTAIL.t5 VN.t6 VDD2.t1 w_n4570_n3366# sky130_fd_pr__pfet_01v8 ad=4.6761 pd=24.76 as=1.97835 ps=12.32 w=11.99 l=3.27
X14 B.t5 B.t3 B.t4 w_n4570_n3366# sky130_fd_pr__pfet_01v8 ad=4.6761 pd=24.76 as=0 ps=0 w=11.99 l=3.27
X15 VTAIL.t7 VN.t7 VDD2.t0 w_n4570_n3366# sky130_fd_pr__pfet_01v8 ad=1.97835 pd=12.32 as=1.97835 ps=12.32 w=11.99 l=3.27
X16 B.t2 B.t0 B.t1 w_n4570_n3366# sky130_fd_pr__pfet_01v8 ad=4.6761 pd=24.76 as=0 ps=0 w=11.99 l=3.27
X17 VTAIL.t13 VP.t5 VDD1.t2 w_n4570_n3366# sky130_fd_pr__pfet_01v8 ad=1.97835 pd=12.32 as=1.97835 ps=12.32 w=11.99 l=3.27
X18 VTAIL.t15 VP.t6 VDD1.t1 w_n4570_n3366# sky130_fd_pr__pfet_01v8 ad=4.6761 pd=24.76 as=1.97835 ps=12.32 w=11.99 l=3.27
X19 VDD1.t0 VP.t7 VTAIL.t14 w_n4570_n3366# sky130_fd_pr__pfet_01v8 ad=1.97835 pd=12.32 as=4.6761 ps=24.76 w=11.99 l=3.27
R0 VP.n24 VP.n23 161.3
R1 VP.n25 VP.n20 161.3
R2 VP.n27 VP.n26 161.3
R3 VP.n28 VP.n19 161.3
R4 VP.n30 VP.n29 161.3
R5 VP.n31 VP.n18 161.3
R6 VP.n33 VP.n32 161.3
R7 VP.n35 VP.n34 161.3
R8 VP.n36 VP.n16 161.3
R9 VP.n38 VP.n37 161.3
R10 VP.n39 VP.n15 161.3
R11 VP.n41 VP.n40 161.3
R12 VP.n42 VP.n14 161.3
R13 VP.n44 VP.n43 161.3
R14 VP.n79 VP.n78 161.3
R15 VP.n77 VP.n1 161.3
R16 VP.n76 VP.n75 161.3
R17 VP.n74 VP.n2 161.3
R18 VP.n73 VP.n72 161.3
R19 VP.n71 VP.n3 161.3
R20 VP.n70 VP.n69 161.3
R21 VP.n68 VP.n67 161.3
R22 VP.n66 VP.n5 161.3
R23 VP.n65 VP.n64 161.3
R24 VP.n63 VP.n6 161.3
R25 VP.n62 VP.n61 161.3
R26 VP.n60 VP.n7 161.3
R27 VP.n59 VP.n58 161.3
R28 VP.n57 VP.n56 161.3
R29 VP.n55 VP.n9 161.3
R30 VP.n54 VP.n53 161.3
R31 VP.n52 VP.n10 161.3
R32 VP.n51 VP.n50 161.3
R33 VP.n49 VP.n11 161.3
R34 VP.n48 VP.n47 161.3
R35 VP.n22 VP.t6 121.709
R36 VP.n12 VP.t4 88.3672
R37 VP.n8 VP.t2 88.3672
R38 VP.n4 VP.t5 88.3672
R39 VP.n0 VP.t7 88.3672
R40 VP.n13 VP.t0 88.3672
R41 VP.n17 VP.t3 88.3672
R42 VP.n21 VP.t1 88.3672
R43 VP.n46 VP.n12 70.4938
R44 VP.n80 VP.n0 70.4938
R45 VP.n45 VP.n13 70.4938
R46 VP.n22 VP.n21 59.4932
R47 VP.n46 VP.n45 54.2039
R48 VP.n50 VP.n10 50.2061
R49 VP.n76 VP.n2 50.2061
R50 VP.n41 VP.n15 50.2061
R51 VP.n61 VP.n6 40.4934
R52 VP.n65 VP.n6 40.4934
R53 VP.n30 VP.n19 40.4934
R54 VP.n26 VP.n19 40.4934
R55 VP.n54 VP.n10 30.7807
R56 VP.n72 VP.n2 30.7807
R57 VP.n37 VP.n15 30.7807
R58 VP.n49 VP.n48 24.4675
R59 VP.n50 VP.n49 24.4675
R60 VP.n55 VP.n54 24.4675
R61 VP.n56 VP.n55 24.4675
R62 VP.n60 VP.n59 24.4675
R63 VP.n61 VP.n60 24.4675
R64 VP.n66 VP.n65 24.4675
R65 VP.n67 VP.n66 24.4675
R66 VP.n71 VP.n70 24.4675
R67 VP.n72 VP.n71 24.4675
R68 VP.n77 VP.n76 24.4675
R69 VP.n78 VP.n77 24.4675
R70 VP.n42 VP.n41 24.4675
R71 VP.n43 VP.n42 24.4675
R72 VP.n31 VP.n30 24.4675
R73 VP.n32 VP.n31 24.4675
R74 VP.n36 VP.n35 24.4675
R75 VP.n37 VP.n36 24.4675
R76 VP.n25 VP.n24 24.4675
R77 VP.n26 VP.n25 24.4675
R78 VP.n48 VP.n12 19.5741
R79 VP.n78 VP.n0 19.5741
R80 VP.n43 VP.n13 19.5741
R81 VP.n59 VP.n8 14.6807
R82 VP.n67 VP.n4 14.6807
R83 VP.n32 VP.n17 14.6807
R84 VP.n24 VP.n21 14.6807
R85 VP.n56 VP.n8 9.7873
R86 VP.n70 VP.n4 9.7873
R87 VP.n35 VP.n17 9.7873
R88 VP.n23 VP.n22 3.92585
R89 VP.n45 VP.n44 0.354971
R90 VP.n47 VP.n46 0.354971
R91 VP.n80 VP.n79 0.354971
R92 VP VP.n80 0.26696
R93 VP.n23 VP.n20 0.189894
R94 VP.n27 VP.n20 0.189894
R95 VP.n28 VP.n27 0.189894
R96 VP.n29 VP.n28 0.189894
R97 VP.n29 VP.n18 0.189894
R98 VP.n33 VP.n18 0.189894
R99 VP.n34 VP.n33 0.189894
R100 VP.n34 VP.n16 0.189894
R101 VP.n38 VP.n16 0.189894
R102 VP.n39 VP.n38 0.189894
R103 VP.n40 VP.n39 0.189894
R104 VP.n40 VP.n14 0.189894
R105 VP.n44 VP.n14 0.189894
R106 VP.n47 VP.n11 0.189894
R107 VP.n51 VP.n11 0.189894
R108 VP.n52 VP.n51 0.189894
R109 VP.n53 VP.n52 0.189894
R110 VP.n53 VP.n9 0.189894
R111 VP.n57 VP.n9 0.189894
R112 VP.n58 VP.n57 0.189894
R113 VP.n58 VP.n7 0.189894
R114 VP.n62 VP.n7 0.189894
R115 VP.n63 VP.n62 0.189894
R116 VP.n64 VP.n63 0.189894
R117 VP.n64 VP.n5 0.189894
R118 VP.n68 VP.n5 0.189894
R119 VP.n69 VP.n68 0.189894
R120 VP.n69 VP.n3 0.189894
R121 VP.n73 VP.n3 0.189894
R122 VP.n74 VP.n73 0.189894
R123 VP.n75 VP.n74 0.189894
R124 VP.n75 VP.n1 0.189894
R125 VP.n79 VP.n1 0.189894
R126 VTAIL.n534 VTAIL.n533 756.745
R127 VTAIL.n66 VTAIL.n65 756.745
R128 VTAIL.n132 VTAIL.n131 756.745
R129 VTAIL.n200 VTAIL.n199 756.745
R130 VTAIL.n468 VTAIL.n467 756.745
R131 VTAIL.n400 VTAIL.n399 756.745
R132 VTAIL.n334 VTAIL.n333 756.745
R133 VTAIL.n266 VTAIL.n265 756.745
R134 VTAIL.n493 VTAIL.n492 585
R135 VTAIL.n495 VTAIL.n494 585
R136 VTAIL.n488 VTAIL.n487 585
R137 VTAIL.n501 VTAIL.n500 585
R138 VTAIL.n503 VTAIL.n502 585
R139 VTAIL.n484 VTAIL.n483 585
R140 VTAIL.n509 VTAIL.n508 585
R141 VTAIL.n511 VTAIL.n510 585
R142 VTAIL.n480 VTAIL.n479 585
R143 VTAIL.n517 VTAIL.n516 585
R144 VTAIL.n519 VTAIL.n518 585
R145 VTAIL.n476 VTAIL.n475 585
R146 VTAIL.n525 VTAIL.n524 585
R147 VTAIL.n527 VTAIL.n526 585
R148 VTAIL.n472 VTAIL.n471 585
R149 VTAIL.n533 VTAIL.n532 585
R150 VTAIL.n25 VTAIL.n24 585
R151 VTAIL.n27 VTAIL.n26 585
R152 VTAIL.n20 VTAIL.n19 585
R153 VTAIL.n33 VTAIL.n32 585
R154 VTAIL.n35 VTAIL.n34 585
R155 VTAIL.n16 VTAIL.n15 585
R156 VTAIL.n41 VTAIL.n40 585
R157 VTAIL.n43 VTAIL.n42 585
R158 VTAIL.n12 VTAIL.n11 585
R159 VTAIL.n49 VTAIL.n48 585
R160 VTAIL.n51 VTAIL.n50 585
R161 VTAIL.n8 VTAIL.n7 585
R162 VTAIL.n57 VTAIL.n56 585
R163 VTAIL.n59 VTAIL.n58 585
R164 VTAIL.n4 VTAIL.n3 585
R165 VTAIL.n65 VTAIL.n64 585
R166 VTAIL.n91 VTAIL.n90 585
R167 VTAIL.n93 VTAIL.n92 585
R168 VTAIL.n86 VTAIL.n85 585
R169 VTAIL.n99 VTAIL.n98 585
R170 VTAIL.n101 VTAIL.n100 585
R171 VTAIL.n82 VTAIL.n81 585
R172 VTAIL.n107 VTAIL.n106 585
R173 VTAIL.n109 VTAIL.n108 585
R174 VTAIL.n78 VTAIL.n77 585
R175 VTAIL.n115 VTAIL.n114 585
R176 VTAIL.n117 VTAIL.n116 585
R177 VTAIL.n74 VTAIL.n73 585
R178 VTAIL.n123 VTAIL.n122 585
R179 VTAIL.n125 VTAIL.n124 585
R180 VTAIL.n70 VTAIL.n69 585
R181 VTAIL.n131 VTAIL.n130 585
R182 VTAIL.n159 VTAIL.n158 585
R183 VTAIL.n161 VTAIL.n160 585
R184 VTAIL.n154 VTAIL.n153 585
R185 VTAIL.n167 VTAIL.n166 585
R186 VTAIL.n169 VTAIL.n168 585
R187 VTAIL.n150 VTAIL.n149 585
R188 VTAIL.n175 VTAIL.n174 585
R189 VTAIL.n177 VTAIL.n176 585
R190 VTAIL.n146 VTAIL.n145 585
R191 VTAIL.n183 VTAIL.n182 585
R192 VTAIL.n185 VTAIL.n184 585
R193 VTAIL.n142 VTAIL.n141 585
R194 VTAIL.n191 VTAIL.n190 585
R195 VTAIL.n193 VTAIL.n192 585
R196 VTAIL.n138 VTAIL.n137 585
R197 VTAIL.n199 VTAIL.n198 585
R198 VTAIL.n467 VTAIL.n466 585
R199 VTAIL.n406 VTAIL.n405 585
R200 VTAIL.n461 VTAIL.n460 585
R201 VTAIL.n459 VTAIL.n458 585
R202 VTAIL.n410 VTAIL.n409 585
R203 VTAIL.n453 VTAIL.n452 585
R204 VTAIL.n451 VTAIL.n450 585
R205 VTAIL.n414 VTAIL.n413 585
R206 VTAIL.n445 VTAIL.n444 585
R207 VTAIL.n443 VTAIL.n442 585
R208 VTAIL.n418 VTAIL.n417 585
R209 VTAIL.n437 VTAIL.n436 585
R210 VTAIL.n435 VTAIL.n434 585
R211 VTAIL.n422 VTAIL.n421 585
R212 VTAIL.n429 VTAIL.n428 585
R213 VTAIL.n427 VTAIL.n426 585
R214 VTAIL.n399 VTAIL.n398 585
R215 VTAIL.n338 VTAIL.n337 585
R216 VTAIL.n393 VTAIL.n392 585
R217 VTAIL.n391 VTAIL.n390 585
R218 VTAIL.n342 VTAIL.n341 585
R219 VTAIL.n385 VTAIL.n384 585
R220 VTAIL.n383 VTAIL.n382 585
R221 VTAIL.n346 VTAIL.n345 585
R222 VTAIL.n377 VTAIL.n376 585
R223 VTAIL.n375 VTAIL.n374 585
R224 VTAIL.n350 VTAIL.n349 585
R225 VTAIL.n369 VTAIL.n368 585
R226 VTAIL.n367 VTAIL.n366 585
R227 VTAIL.n354 VTAIL.n353 585
R228 VTAIL.n361 VTAIL.n360 585
R229 VTAIL.n359 VTAIL.n358 585
R230 VTAIL.n333 VTAIL.n332 585
R231 VTAIL.n272 VTAIL.n271 585
R232 VTAIL.n327 VTAIL.n326 585
R233 VTAIL.n325 VTAIL.n324 585
R234 VTAIL.n276 VTAIL.n275 585
R235 VTAIL.n319 VTAIL.n318 585
R236 VTAIL.n317 VTAIL.n316 585
R237 VTAIL.n280 VTAIL.n279 585
R238 VTAIL.n311 VTAIL.n310 585
R239 VTAIL.n309 VTAIL.n308 585
R240 VTAIL.n284 VTAIL.n283 585
R241 VTAIL.n303 VTAIL.n302 585
R242 VTAIL.n301 VTAIL.n300 585
R243 VTAIL.n288 VTAIL.n287 585
R244 VTAIL.n295 VTAIL.n294 585
R245 VTAIL.n293 VTAIL.n292 585
R246 VTAIL.n265 VTAIL.n264 585
R247 VTAIL.n204 VTAIL.n203 585
R248 VTAIL.n259 VTAIL.n258 585
R249 VTAIL.n257 VTAIL.n256 585
R250 VTAIL.n208 VTAIL.n207 585
R251 VTAIL.n251 VTAIL.n250 585
R252 VTAIL.n249 VTAIL.n248 585
R253 VTAIL.n212 VTAIL.n211 585
R254 VTAIL.n243 VTAIL.n242 585
R255 VTAIL.n241 VTAIL.n240 585
R256 VTAIL.n216 VTAIL.n215 585
R257 VTAIL.n235 VTAIL.n234 585
R258 VTAIL.n233 VTAIL.n232 585
R259 VTAIL.n220 VTAIL.n219 585
R260 VTAIL.n227 VTAIL.n226 585
R261 VTAIL.n225 VTAIL.n224 585
R262 VTAIL.n425 VTAIL.t11 327.466
R263 VTAIL.n357 VTAIL.t15 327.466
R264 VTAIL.n291 VTAIL.t0 327.466
R265 VTAIL.n223 VTAIL.t5 327.466
R266 VTAIL.n491 VTAIL.t1 327.466
R267 VTAIL.n23 VTAIL.t4 327.466
R268 VTAIL.n89 VTAIL.t14 327.466
R269 VTAIL.n157 VTAIL.t9 327.466
R270 VTAIL.n494 VTAIL.n493 171.744
R271 VTAIL.n494 VTAIL.n487 171.744
R272 VTAIL.n501 VTAIL.n487 171.744
R273 VTAIL.n502 VTAIL.n501 171.744
R274 VTAIL.n502 VTAIL.n483 171.744
R275 VTAIL.n509 VTAIL.n483 171.744
R276 VTAIL.n510 VTAIL.n509 171.744
R277 VTAIL.n510 VTAIL.n479 171.744
R278 VTAIL.n517 VTAIL.n479 171.744
R279 VTAIL.n518 VTAIL.n517 171.744
R280 VTAIL.n518 VTAIL.n475 171.744
R281 VTAIL.n525 VTAIL.n475 171.744
R282 VTAIL.n526 VTAIL.n525 171.744
R283 VTAIL.n526 VTAIL.n471 171.744
R284 VTAIL.n533 VTAIL.n471 171.744
R285 VTAIL.n26 VTAIL.n25 171.744
R286 VTAIL.n26 VTAIL.n19 171.744
R287 VTAIL.n33 VTAIL.n19 171.744
R288 VTAIL.n34 VTAIL.n33 171.744
R289 VTAIL.n34 VTAIL.n15 171.744
R290 VTAIL.n41 VTAIL.n15 171.744
R291 VTAIL.n42 VTAIL.n41 171.744
R292 VTAIL.n42 VTAIL.n11 171.744
R293 VTAIL.n49 VTAIL.n11 171.744
R294 VTAIL.n50 VTAIL.n49 171.744
R295 VTAIL.n50 VTAIL.n7 171.744
R296 VTAIL.n57 VTAIL.n7 171.744
R297 VTAIL.n58 VTAIL.n57 171.744
R298 VTAIL.n58 VTAIL.n3 171.744
R299 VTAIL.n65 VTAIL.n3 171.744
R300 VTAIL.n92 VTAIL.n91 171.744
R301 VTAIL.n92 VTAIL.n85 171.744
R302 VTAIL.n99 VTAIL.n85 171.744
R303 VTAIL.n100 VTAIL.n99 171.744
R304 VTAIL.n100 VTAIL.n81 171.744
R305 VTAIL.n107 VTAIL.n81 171.744
R306 VTAIL.n108 VTAIL.n107 171.744
R307 VTAIL.n108 VTAIL.n77 171.744
R308 VTAIL.n115 VTAIL.n77 171.744
R309 VTAIL.n116 VTAIL.n115 171.744
R310 VTAIL.n116 VTAIL.n73 171.744
R311 VTAIL.n123 VTAIL.n73 171.744
R312 VTAIL.n124 VTAIL.n123 171.744
R313 VTAIL.n124 VTAIL.n69 171.744
R314 VTAIL.n131 VTAIL.n69 171.744
R315 VTAIL.n160 VTAIL.n159 171.744
R316 VTAIL.n160 VTAIL.n153 171.744
R317 VTAIL.n167 VTAIL.n153 171.744
R318 VTAIL.n168 VTAIL.n167 171.744
R319 VTAIL.n168 VTAIL.n149 171.744
R320 VTAIL.n175 VTAIL.n149 171.744
R321 VTAIL.n176 VTAIL.n175 171.744
R322 VTAIL.n176 VTAIL.n145 171.744
R323 VTAIL.n183 VTAIL.n145 171.744
R324 VTAIL.n184 VTAIL.n183 171.744
R325 VTAIL.n184 VTAIL.n141 171.744
R326 VTAIL.n191 VTAIL.n141 171.744
R327 VTAIL.n192 VTAIL.n191 171.744
R328 VTAIL.n192 VTAIL.n137 171.744
R329 VTAIL.n199 VTAIL.n137 171.744
R330 VTAIL.n467 VTAIL.n405 171.744
R331 VTAIL.n460 VTAIL.n405 171.744
R332 VTAIL.n460 VTAIL.n459 171.744
R333 VTAIL.n459 VTAIL.n409 171.744
R334 VTAIL.n452 VTAIL.n409 171.744
R335 VTAIL.n452 VTAIL.n451 171.744
R336 VTAIL.n451 VTAIL.n413 171.744
R337 VTAIL.n444 VTAIL.n413 171.744
R338 VTAIL.n444 VTAIL.n443 171.744
R339 VTAIL.n443 VTAIL.n417 171.744
R340 VTAIL.n436 VTAIL.n417 171.744
R341 VTAIL.n436 VTAIL.n435 171.744
R342 VTAIL.n435 VTAIL.n421 171.744
R343 VTAIL.n428 VTAIL.n421 171.744
R344 VTAIL.n428 VTAIL.n427 171.744
R345 VTAIL.n399 VTAIL.n337 171.744
R346 VTAIL.n392 VTAIL.n337 171.744
R347 VTAIL.n392 VTAIL.n391 171.744
R348 VTAIL.n391 VTAIL.n341 171.744
R349 VTAIL.n384 VTAIL.n341 171.744
R350 VTAIL.n384 VTAIL.n383 171.744
R351 VTAIL.n383 VTAIL.n345 171.744
R352 VTAIL.n376 VTAIL.n345 171.744
R353 VTAIL.n376 VTAIL.n375 171.744
R354 VTAIL.n375 VTAIL.n349 171.744
R355 VTAIL.n368 VTAIL.n349 171.744
R356 VTAIL.n368 VTAIL.n367 171.744
R357 VTAIL.n367 VTAIL.n353 171.744
R358 VTAIL.n360 VTAIL.n353 171.744
R359 VTAIL.n360 VTAIL.n359 171.744
R360 VTAIL.n333 VTAIL.n271 171.744
R361 VTAIL.n326 VTAIL.n271 171.744
R362 VTAIL.n326 VTAIL.n325 171.744
R363 VTAIL.n325 VTAIL.n275 171.744
R364 VTAIL.n318 VTAIL.n275 171.744
R365 VTAIL.n318 VTAIL.n317 171.744
R366 VTAIL.n317 VTAIL.n279 171.744
R367 VTAIL.n310 VTAIL.n279 171.744
R368 VTAIL.n310 VTAIL.n309 171.744
R369 VTAIL.n309 VTAIL.n283 171.744
R370 VTAIL.n302 VTAIL.n283 171.744
R371 VTAIL.n302 VTAIL.n301 171.744
R372 VTAIL.n301 VTAIL.n287 171.744
R373 VTAIL.n294 VTAIL.n287 171.744
R374 VTAIL.n294 VTAIL.n293 171.744
R375 VTAIL.n265 VTAIL.n203 171.744
R376 VTAIL.n258 VTAIL.n203 171.744
R377 VTAIL.n258 VTAIL.n257 171.744
R378 VTAIL.n257 VTAIL.n207 171.744
R379 VTAIL.n250 VTAIL.n207 171.744
R380 VTAIL.n250 VTAIL.n249 171.744
R381 VTAIL.n249 VTAIL.n211 171.744
R382 VTAIL.n242 VTAIL.n211 171.744
R383 VTAIL.n242 VTAIL.n241 171.744
R384 VTAIL.n241 VTAIL.n215 171.744
R385 VTAIL.n234 VTAIL.n215 171.744
R386 VTAIL.n234 VTAIL.n233 171.744
R387 VTAIL.n233 VTAIL.n219 171.744
R388 VTAIL.n226 VTAIL.n219 171.744
R389 VTAIL.n226 VTAIL.n225 171.744
R390 VTAIL.n493 VTAIL.t1 85.8723
R391 VTAIL.n25 VTAIL.t4 85.8723
R392 VTAIL.n91 VTAIL.t14 85.8723
R393 VTAIL.n159 VTAIL.t9 85.8723
R394 VTAIL.n427 VTAIL.t11 85.8723
R395 VTAIL.n359 VTAIL.t15 85.8723
R396 VTAIL.n293 VTAIL.t0 85.8723
R397 VTAIL.n225 VTAIL.t5 85.8723
R398 VTAIL.n403 VTAIL.n402 61.1977
R399 VTAIL.n269 VTAIL.n268 61.1977
R400 VTAIL.n1 VTAIL.n0 61.1976
R401 VTAIL.n135 VTAIL.n134 61.1976
R402 VTAIL.n535 VTAIL.n534 35.4823
R403 VTAIL.n67 VTAIL.n66 35.4823
R404 VTAIL.n133 VTAIL.n132 35.4823
R405 VTAIL.n201 VTAIL.n200 35.4823
R406 VTAIL.n469 VTAIL.n468 35.4823
R407 VTAIL.n401 VTAIL.n400 35.4823
R408 VTAIL.n335 VTAIL.n334 35.4823
R409 VTAIL.n267 VTAIL.n266 35.4823
R410 VTAIL.n535 VTAIL.n469 25.8065
R411 VTAIL.n267 VTAIL.n201 25.8065
R412 VTAIL.n492 VTAIL.n491 16.3895
R413 VTAIL.n24 VTAIL.n23 16.3895
R414 VTAIL.n90 VTAIL.n89 16.3895
R415 VTAIL.n158 VTAIL.n157 16.3895
R416 VTAIL.n426 VTAIL.n425 16.3895
R417 VTAIL.n358 VTAIL.n357 16.3895
R418 VTAIL.n292 VTAIL.n291 16.3895
R419 VTAIL.n224 VTAIL.n223 16.3895
R420 VTAIL.n495 VTAIL.n490 12.8005
R421 VTAIL.n27 VTAIL.n22 12.8005
R422 VTAIL.n93 VTAIL.n88 12.8005
R423 VTAIL.n161 VTAIL.n156 12.8005
R424 VTAIL.n429 VTAIL.n424 12.8005
R425 VTAIL.n361 VTAIL.n356 12.8005
R426 VTAIL.n295 VTAIL.n290 12.8005
R427 VTAIL.n227 VTAIL.n222 12.8005
R428 VTAIL.n496 VTAIL.n488 12.0247
R429 VTAIL.n532 VTAIL.n470 12.0247
R430 VTAIL.n28 VTAIL.n20 12.0247
R431 VTAIL.n64 VTAIL.n2 12.0247
R432 VTAIL.n94 VTAIL.n86 12.0247
R433 VTAIL.n130 VTAIL.n68 12.0247
R434 VTAIL.n162 VTAIL.n154 12.0247
R435 VTAIL.n198 VTAIL.n136 12.0247
R436 VTAIL.n466 VTAIL.n404 12.0247
R437 VTAIL.n430 VTAIL.n422 12.0247
R438 VTAIL.n398 VTAIL.n336 12.0247
R439 VTAIL.n362 VTAIL.n354 12.0247
R440 VTAIL.n332 VTAIL.n270 12.0247
R441 VTAIL.n296 VTAIL.n288 12.0247
R442 VTAIL.n264 VTAIL.n202 12.0247
R443 VTAIL.n228 VTAIL.n220 12.0247
R444 VTAIL.n500 VTAIL.n499 11.249
R445 VTAIL.n531 VTAIL.n472 11.249
R446 VTAIL.n32 VTAIL.n31 11.249
R447 VTAIL.n63 VTAIL.n4 11.249
R448 VTAIL.n98 VTAIL.n97 11.249
R449 VTAIL.n129 VTAIL.n70 11.249
R450 VTAIL.n166 VTAIL.n165 11.249
R451 VTAIL.n197 VTAIL.n138 11.249
R452 VTAIL.n465 VTAIL.n406 11.249
R453 VTAIL.n434 VTAIL.n433 11.249
R454 VTAIL.n397 VTAIL.n338 11.249
R455 VTAIL.n366 VTAIL.n365 11.249
R456 VTAIL.n331 VTAIL.n272 11.249
R457 VTAIL.n300 VTAIL.n299 11.249
R458 VTAIL.n263 VTAIL.n204 11.249
R459 VTAIL.n232 VTAIL.n231 11.249
R460 VTAIL.n503 VTAIL.n486 10.4732
R461 VTAIL.n528 VTAIL.n527 10.4732
R462 VTAIL.n35 VTAIL.n18 10.4732
R463 VTAIL.n60 VTAIL.n59 10.4732
R464 VTAIL.n101 VTAIL.n84 10.4732
R465 VTAIL.n126 VTAIL.n125 10.4732
R466 VTAIL.n169 VTAIL.n152 10.4732
R467 VTAIL.n194 VTAIL.n193 10.4732
R468 VTAIL.n462 VTAIL.n461 10.4732
R469 VTAIL.n437 VTAIL.n420 10.4732
R470 VTAIL.n394 VTAIL.n393 10.4732
R471 VTAIL.n369 VTAIL.n352 10.4732
R472 VTAIL.n328 VTAIL.n327 10.4732
R473 VTAIL.n303 VTAIL.n286 10.4732
R474 VTAIL.n260 VTAIL.n259 10.4732
R475 VTAIL.n235 VTAIL.n218 10.4732
R476 VTAIL.n504 VTAIL.n484 9.69747
R477 VTAIL.n524 VTAIL.n474 9.69747
R478 VTAIL.n36 VTAIL.n16 9.69747
R479 VTAIL.n56 VTAIL.n6 9.69747
R480 VTAIL.n102 VTAIL.n82 9.69747
R481 VTAIL.n122 VTAIL.n72 9.69747
R482 VTAIL.n170 VTAIL.n150 9.69747
R483 VTAIL.n190 VTAIL.n140 9.69747
R484 VTAIL.n458 VTAIL.n408 9.69747
R485 VTAIL.n438 VTAIL.n418 9.69747
R486 VTAIL.n390 VTAIL.n340 9.69747
R487 VTAIL.n370 VTAIL.n350 9.69747
R488 VTAIL.n324 VTAIL.n274 9.69747
R489 VTAIL.n304 VTAIL.n284 9.69747
R490 VTAIL.n256 VTAIL.n206 9.69747
R491 VTAIL.n236 VTAIL.n216 9.69747
R492 VTAIL.n530 VTAIL.n470 9.45567
R493 VTAIL.n62 VTAIL.n2 9.45567
R494 VTAIL.n128 VTAIL.n68 9.45567
R495 VTAIL.n196 VTAIL.n136 9.45567
R496 VTAIL.n464 VTAIL.n404 9.45567
R497 VTAIL.n396 VTAIL.n336 9.45567
R498 VTAIL.n330 VTAIL.n270 9.45567
R499 VTAIL.n262 VTAIL.n202 9.45567
R500 VTAIL.n515 VTAIL.n514 9.3005
R501 VTAIL.n478 VTAIL.n477 9.3005
R502 VTAIL.n521 VTAIL.n520 9.3005
R503 VTAIL.n523 VTAIL.n522 9.3005
R504 VTAIL.n474 VTAIL.n473 9.3005
R505 VTAIL.n529 VTAIL.n528 9.3005
R506 VTAIL.n531 VTAIL.n530 9.3005
R507 VTAIL.n482 VTAIL.n481 9.3005
R508 VTAIL.n507 VTAIL.n506 9.3005
R509 VTAIL.n505 VTAIL.n504 9.3005
R510 VTAIL.n486 VTAIL.n485 9.3005
R511 VTAIL.n499 VTAIL.n498 9.3005
R512 VTAIL.n497 VTAIL.n496 9.3005
R513 VTAIL.n490 VTAIL.n489 9.3005
R514 VTAIL.n513 VTAIL.n512 9.3005
R515 VTAIL.n47 VTAIL.n46 9.3005
R516 VTAIL.n10 VTAIL.n9 9.3005
R517 VTAIL.n53 VTAIL.n52 9.3005
R518 VTAIL.n55 VTAIL.n54 9.3005
R519 VTAIL.n6 VTAIL.n5 9.3005
R520 VTAIL.n61 VTAIL.n60 9.3005
R521 VTAIL.n63 VTAIL.n62 9.3005
R522 VTAIL.n14 VTAIL.n13 9.3005
R523 VTAIL.n39 VTAIL.n38 9.3005
R524 VTAIL.n37 VTAIL.n36 9.3005
R525 VTAIL.n18 VTAIL.n17 9.3005
R526 VTAIL.n31 VTAIL.n30 9.3005
R527 VTAIL.n29 VTAIL.n28 9.3005
R528 VTAIL.n22 VTAIL.n21 9.3005
R529 VTAIL.n45 VTAIL.n44 9.3005
R530 VTAIL.n113 VTAIL.n112 9.3005
R531 VTAIL.n76 VTAIL.n75 9.3005
R532 VTAIL.n119 VTAIL.n118 9.3005
R533 VTAIL.n121 VTAIL.n120 9.3005
R534 VTAIL.n72 VTAIL.n71 9.3005
R535 VTAIL.n127 VTAIL.n126 9.3005
R536 VTAIL.n129 VTAIL.n128 9.3005
R537 VTAIL.n80 VTAIL.n79 9.3005
R538 VTAIL.n105 VTAIL.n104 9.3005
R539 VTAIL.n103 VTAIL.n102 9.3005
R540 VTAIL.n84 VTAIL.n83 9.3005
R541 VTAIL.n97 VTAIL.n96 9.3005
R542 VTAIL.n95 VTAIL.n94 9.3005
R543 VTAIL.n88 VTAIL.n87 9.3005
R544 VTAIL.n111 VTAIL.n110 9.3005
R545 VTAIL.n181 VTAIL.n180 9.3005
R546 VTAIL.n144 VTAIL.n143 9.3005
R547 VTAIL.n187 VTAIL.n186 9.3005
R548 VTAIL.n189 VTAIL.n188 9.3005
R549 VTAIL.n140 VTAIL.n139 9.3005
R550 VTAIL.n195 VTAIL.n194 9.3005
R551 VTAIL.n197 VTAIL.n196 9.3005
R552 VTAIL.n148 VTAIL.n147 9.3005
R553 VTAIL.n173 VTAIL.n172 9.3005
R554 VTAIL.n171 VTAIL.n170 9.3005
R555 VTAIL.n152 VTAIL.n151 9.3005
R556 VTAIL.n165 VTAIL.n164 9.3005
R557 VTAIL.n163 VTAIL.n162 9.3005
R558 VTAIL.n156 VTAIL.n155 9.3005
R559 VTAIL.n179 VTAIL.n178 9.3005
R560 VTAIL.n465 VTAIL.n464 9.3005
R561 VTAIL.n463 VTAIL.n462 9.3005
R562 VTAIL.n408 VTAIL.n407 9.3005
R563 VTAIL.n457 VTAIL.n456 9.3005
R564 VTAIL.n455 VTAIL.n454 9.3005
R565 VTAIL.n412 VTAIL.n411 9.3005
R566 VTAIL.n449 VTAIL.n448 9.3005
R567 VTAIL.n447 VTAIL.n446 9.3005
R568 VTAIL.n416 VTAIL.n415 9.3005
R569 VTAIL.n441 VTAIL.n440 9.3005
R570 VTAIL.n439 VTAIL.n438 9.3005
R571 VTAIL.n420 VTAIL.n419 9.3005
R572 VTAIL.n433 VTAIL.n432 9.3005
R573 VTAIL.n431 VTAIL.n430 9.3005
R574 VTAIL.n424 VTAIL.n423 9.3005
R575 VTAIL.n344 VTAIL.n343 9.3005
R576 VTAIL.n387 VTAIL.n386 9.3005
R577 VTAIL.n389 VTAIL.n388 9.3005
R578 VTAIL.n340 VTAIL.n339 9.3005
R579 VTAIL.n395 VTAIL.n394 9.3005
R580 VTAIL.n397 VTAIL.n396 9.3005
R581 VTAIL.n381 VTAIL.n380 9.3005
R582 VTAIL.n379 VTAIL.n378 9.3005
R583 VTAIL.n348 VTAIL.n347 9.3005
R584 VTAIL.n373 VTAIL.n372 9.3005
R585 VTAIL.n371 VTAIL.n370 9.3005
R586 VTAIL.n352 VTAIL.n351 9.3005
R587 VTAIL.n365 VTAIL.n364 9.3005
R588 VTAIL.n363 VTAIL.n362 9.3005
R589 VTAIL.n356 VTAIL.n355 9.3005
R590 VTAIL.n278 VTAIL.n277 9.3005
R591 VTAIL.n321 VTAIL.n320 9.3005
R592 VTAIL.n323 VTAIL.n322 9.3005
R593 VTAIL.n274 VTAIL.n273 9.3005
R594 VTAIL.n329 VTAIL.n328 9.3005
R595 VTAIL.n331 VTAIL.n330 9.3005
R596 VTAIL.n315 VTAIL.n314 9.3005
R597 VTAIL.n313 VTAIL.n312 9.3005
R598 VTAIL.n282 VTAIL.n281 9.3005
R599 VTAIL.n307 VTAIL.n306 9.3005
R600 VTAIL.n305 VTAIL.n304 9.3005
R601 VTAIL.n286 VTAIL.n285 9.3005
R602 VTAIL.n299 VTAIL.n298 9.3005
R603 VTAIL.n297 VTAIL.n296 9.3005
R604 VTAIL.n290 VTAIL.n289 9.3005
R605 VTAIL.n210 VTAIL.n209 9.3005
R606 VTAIL.n253 VTAIL.n252 9.3005
R607 VTAIL.n255 VTAIL.n254 9.3005
R608 VTAIL.n206 VTAIL.n205 9.3005
R609 VTAIL.n261 VTAIL.n260 9.3005
R610 VTAIL.n263 VTAIL.n262 9.3005
R611 VTAIL.n247 VTAIL.n246 9.3005
R612 VTAIL.n245 VTAIL.n244 9.3005
R613 VTAIL.n214 VTAIL.n213 9.3005
R614 VTAIL.n239 VTAIL.n238 9.3005
R615 VTAIL.n237 VTAIL.n236 9.3005
R616 VTAIL.n218 VTAIL.n217 9.3005
R617 VTAIL.n231 VTAIL.n230 9.3005
R618 VTAIL.n229 VTAIL.n228 9.3005
R619 VTAIL.n222 VTAIL.n221 9.3005
R620 VTAIL.n508 VTAIL.n507 8.92171
R621 VTAIL.n523 VTAIL.n476 8.92171
R622 VTAIL.n40 VTAIL.n39 8.92171
R623 VTAIL.n55 VTAIL.n8 8.92171
R624 VTAIL.n106 VTAIL.n105 8.92171
R625 VTAIL.n121 VTAIL.n74 8.92171
R626 VTAIL.n174 VTAIL.n173 8.92171
R627 VTAIL.n189 VTAIL.n142 8.92171
R628 VTAIL.n457 VTAIL.n410 8.92171
R629 VTAIL.n442 VTAIL.n441 8.92171
R630 VTAIL.n389 VTAIL.n342 8.92171
R631 VTAIL.n374 VTAIL.n373 8.92171
R632 VTAIL.n323 VTAIL.n276 8.92171
R633 VTAIL.n308 VTAIL.n307 8.92171
R634 VTAIL.n255 VTAIL.n208 8.92171
R635 VTAIL.n240 VTAIL.n239 8.92171
R636 VTAIL.n511 VTAIL.n482 8.14595
R637 VTAIL.n520 VTAIL.n519 8.14595
R638 VTAIL.n43 VTAIL.n14 8.14595
R639 VTAIL.n52 VTAIL.n51 8.14595
R640 VTAIL.n109 VTAIL.n80 8.14595
R641 VTAIL.n118 VTAIL.n117 8.14595
R642 VTAIL.n177 VTAIL.n148 8.14595
R643 VTAIL.n186 VTAIL.n185 8.14595
R644 VTAIL.n454 VTAIL.n453 8.14595
R645 VTAIL.n445 VTAIL.n416 8.14595
R646 VTAIL.n386 VTAIL.n385 8.14595
R647 VTAIL.n377 VTAIL.n348 8.14595
R648 VTAIL.n320 VTAIL.n319 8.14595
R649 VTAIL.n311 VTAIL.n282 8.14595
R650 VTAIL.n252 VTAIL.n251 8.14595
R651 VTAIL.n243 VTAIL.n214 8.14595
R652 VTAIL.n512 VTAIL.n480 7.3702
R653 VTAIL.n516 VTAIL.n478 7.3702
R654 VTAIL.n44 VTAIL.n12 7.3702
R655 VTAIL.n48 VTAIL.n10 7.3702
R656 VTAIL.n110 VTAIL.n78 7.3702
R657 VTAIL.n114 VTAIL.n76 7.3702
R658 VTAIL.n178 VTAIL.n146 7.3702
R659 VTAIL.n182 VTAIL.n144 7.3702
R660 VTAIL.n450 VTAIL.n412 7.3702
R661 VTAIL.n446 VTAIL.n414 7.3702
R662 VTAIL.n382 VTAIL.n344 7.3702
R663 VTAIL.n378 VTAIL.n346 7.3702
R664 VTAIL.n316 VTAIL.n278 7.3702
R665 VTAIL.n312 VTAIL.n280 7.3702
R666 VTAIL.n248 VTAIL.n210 7.3702
R667 VTAIL.n244 VTAIL.n212 7.3702
R668 VTAIL.n515 VTAIL.n480 6.59444
R669 VTAIL.n516 VTAIL.n515 6.59444
R670 VTAIL.n47 VTAIL.n12 6.59444
R671 VTAIL.n48 VTAIL.n47 6.59444
R672 VTAIL.n113 VTAIL.n78 6.59444
R673 VTAIL.n114 VTAIL.n113 6.59444
R674 VTAIL.n181 VTAIL.n146 6.59444
R675 VTAIL.n182 VTAIL.n181 6.59444
R676 VTAIL.n450 VTAIL.n449 6.59444
R677 VTAIL.n449 VTAIL.n414 6.59444
R678 VTAIL.n382 VTAIL.n381 6.59444
R679 VTAIL.n381 VTAIL.n346 6.59444
R680 VTAIL.n316 VTAIL.n315 6.59444
R681 VTAIL.n315 VTAIL.n280 6.59444
R682 VTAIL.n248 VTAIL.n247 6.59444
R683 VTAIL.n247 VTAIL.n212 6.59444
R684 VTAIL.n512 VTAIL.n511 5.81868
R685 VTAIL.n519 VTAIL.n478 5.81868
R686 VTAIL.n44 VTAIL.n43 5.81868
R687 VTAIL.n51 VTAIL.n10 5.81868
R688 VTAIL.n110 VTAIL.n109 5.81868
R689 VTAIL.n117 VTAIL.n76 5.81868
R690 VTAIL.n178 VTAIL.n177 5.81868
R691 VTAIL.n185 VTAIL.n144 5.81868
R692 VTAIL.n453 VTAIL.n412 5.81868
R693 VTAIL.n446 VTAIL.n445 5.81868
R694 VTAIL.n385 VTAIL.n344 5.81868
R695 VTAIL.n378 VTAIL.n377 5.81868
R696 VTAIL.n319 VTAIL.n278 5.81868
R697 VTAIL.n312 VTAIL.n311 5.81868
R698 VTAIL.n251 VTAIL.n210 5.81868
R699 VTAIL.n244 VTAIL.n243 5.81868
R700 VTAIL.n508 VTAIL.n482 5.04292
R701 VTAIL.n520 VTAIL.n476 5.04292
R702 VTAIL.n40 VTAIL.n14 5.04292
R703 VTAIL.n52 VTAIL.n8 5.04292
R704 VTAIL.n106 VTAIL.n80 5.04292
R705 VTAIL.n118 VTAIL.n74 5.04292
R706 VTAIL.n174 VTAIL.n148 5.04292
R707 VTAIL.n186 VTAIL.n142 5.04292
R708 VTAIL.n454 VTAIL.n410 5.04292
R709 VTAIL.n442 VTAIL.n416 5.04292
R710 VTAIL.n386 VTAIL.n342 5.04292
R711 VTAIL.n374 VTAIL.n348 5.04292
R712 VTAIL.n320 VTAIL.n276 5.04292
R713 VTAIL.n308 VTAIL.n282 5.04292
R714 VTAIL.n252 VTAIL.n208 5.04292
R715 VTAIL.n240 VTAIL.n214 5.04292
R716 VTAIL.n507 VTAIL.n484 4.26717
R717 VTAIL.n524 VTAIL.n523 4.26717
R718 VTAIL.n39 VTAIL.n16 4.26717
R719 VTAIL.n56 VTAIL.n55 4.26717
R720 VTAIL.n105 VTAIL.n82 4.26717
R721 VTAIL.n122 VTAIL.n121 4.26717
R722 VTAIL.n173 VTAIL.n150 4.26717
R723 VTAIL.n190 VTAIL.n189 4.26717
R724 VTAIL.n458 VTAIL.n457 4.26717
R725 VTAIL.n441 VTAIL.n418 4.26717
R726 VTAIL.n390 VTAIL.n389 4.26717
R727 VTAIL.n373 VTAIL.n350 4.26717
R728 VTAIL.n324 VTAIL.n323 4.26717
R729 VTAIL.n307 VTAIL.n284 4.26717
R730 VTAIL.n256 VTAIL.n255 4.26717
R731 VTAIL.n239 VTAIL.n216 4.26717
R732 VTAIL.n425 VTAIL.n423 3.70982
R733 VTAIL.n357 VTAIL.n355 3.70982
R734 VTAIL.n291 VTAIL.n289 3.70982
R735 VTAIL.n223 VTAIL.n221 3.70982
R736 VTAIL.n491 VTAIL.n489 3.70982
R737 VTAIL.n23 VTAIL.n21 3.70982
R738 VTAIL.n89 VTAIL.n87 3.70982
R739 VTAIL.n157 VTAIL.n155 3.70982
R740 VTAIL.n504 VTAIL.n503 3.49141
R741 VTAIL.n527 VTAIL.n474 3.49141
R742 VTAIL.n36 VTAIL.n35 3.49141
R743 VTAIL.n59 VTAIL.n6 3.49141
R744 VTAIL.n102 VTAIL.n101 3.49141
R745 VTAIL.n125 VTAIL.n72 3.49141
R746 VTAIL.n170 VTAIL.n169 3.49141
R747 VTAIL.n193 VTAIL.n140 3.49141
R748 VTAIL.n461 VTAIL.n408 3.49141
R749 VTAIL.n438 VTAIL.n437 3.49141
R750 VTAIL.n393 VTAIL.n340 3.49141
R751 VTAIL.n370 VTAIL.n369 3.49141
R752 VTAIL.n327 VTAIL.n274 3.49141
R753 VTAIL.n304 VTAIL.n303 3.49141
R754 VTAIL.n259 VTAIL.n206 3.49141
R755 VTAIL.n236 VTAIL.n235 3.49141
R756 VTAIL.n269 VTAIL.n267 3.10395
R757 VTAIL.n335 VTAIL.n269 3.10395
R758 VTAIL.n403 VTAIL.n401 3.10395
R759 VTAIL.n469 VTAIL.n403 3.10395
R760 VTAIL.n201 VTAIL.n135 3.10395
R761 VTAIL.n135 VTAIL.n133 3.10395
R762 VTAIL.n67 VTAIL.n1 3.10395
R763 VTAIL VTAIL.n535 3.04576
R764 VTAIL.n500 VTAIL.n486 2.71565
R765 VTAIL.n528 VTAIL.n472 2.71565
R766 VTAIL.n32 VTAIL.n18 2.71565
R767 VTAIL.n60 VTAIL.n4 2.71565
R768 VTAIL.n98 VTAIL.n84 2.71565
R769 VTAIL.n126 VTAIL.n70 2.71565
R770 VTAIL.n166 VTAIL.n152 2.71565
R771 VTAIL.n194 VTAIL.n138 2.71565
R772 VTAIL.n462 VTAIL.n406 2.71565
R773 VTAIL.n434 VTAIL.n420 2.71565
R774 VTAIL.n394 VTAIL.n338 2.71565
R775 VTAIL.n366 VTAIL.n352 2.71565
R776 VTAIL.n328 VTAIL.n272 2.71565
R777 VTAIL.n300 VTAIL.n286 2.71565
R778 VTAIL.n260 VTAIL.n204 2.71565
R779 VTAIL.n232 VTAIL.n218 2.71565
R780 VTAIL.n0 VTAIL.t6 2.71151
R781 VTAIL.n0 VTAIL.t3 2.71151
R782 VTAIL.n134 VTAIL.t12 2.71151
R783 VTAIL.n134 VTAIL.t13 2.71151
R784 VTAIL.n402 VTAIL.t8 2.71151
R785 VTAIL.n402 VTAIL.t10 2.71151
R786 VTAIL.n268 VTAIL.t2 2.71151
R787 VTAIL.n268 VTAIL.t7 2.71151
R788 VTAIL.n499 VTAIL.n488 1.93989
R789 VTAIL.n532 VTAIL.n531 1.93989
R790 VTAIL.n31 VTAIL.n20 1.93989
R791 VTAIL.n64 VTAIL.n63 1.93989
R792 VTAIL.n97 VTAIL.n86 1.93989
R793 VTAIL.n130 VTAIL.n129 1.93989
R794 VTAIL.n165 VTAIL.n154 1.93989
R795 VTAIL.n198 VTAIL.n197 1.93989
R796 VTAIL.n466 VTAIL.n465 1.93989
R797 VTAIL.n433 VTAIL.n422 1.93989
R798 VTAIL.n398 VTAIL.n397 1.93989
R799 VTAIL.n365 VTAIL.n354 1.93989
R800 VTAIL.n332 VTAIL.n331 1.93989
R801 VTAIL.n299 VTAIL.n288 1.93989
R802 VTAIL.n264 VTAIL.n263 1.93989
R803 VTAIL.n231 VTAIL.n220 1.93989
R804 VTAIL.n496 VTAIL.n495 1.16414
R805 VTAIL.n534 VTAIL.n470 1.16414
R806 VTAIL.n28 VTAIL.n27 1.16414
R807 VTAIL.n66 VTAIL.n2 1.16414
R808 VTAIL.n94 VTAIL.n93 1.16414
R809 VTAIL.n132 VTAIL.n68 1.16414
R810 VTAIL.n162 VTAIL.n161 1.16414
R811 VTAIL.n200 VTAIL.n136 1.16414
R812 VTAIL.n468 VTAIL.n404 1.16414
R813 VTAIL.n430 VTAIL.n429 1.16414
R814 VTAIL.n400 VTAIL.n336 1.16414
R815 VTAIL.n362 VTAIL.n361 1.16414
R816 VTAIL.n334 VTAIL.n270 1.16414
R817 VTAIL.n296 VTAIL.n295 1.16414
R818 VTAIL.n266 VTAIL.n202 1.16414
R819 VTAIL.n228 VTAIL.n227 1.16414
R820 VTAIL.n401 VTAIL.n335 0.470328
R821 VTAIL.n133 VTAIL.n67 0.470328
R822 VTAIL.n492 VTAIL.n490 0.388379
R823 VTAIL.n24 VTAIL.n22 0.388379
R824 VTAIL.n90 VTAIL.n88 0.388379
R825 VTAIL.n158 VTAIL.n156 0.388379
R826 VTAIL.n426 VTAIL.n424 0.388379
R827 VTAIL.n358 VTAIL.n356 0.388379
R828 VTAIL.n292 VTAIL.n290 0.388379
R829 VTAIL.n224 VTAIL.n222 0.388379
R830 VTAIL.n497 VTAIL.n489 0.155672
R831 VTAIL.n498 VTAIL.n497 0.155672
R832 VTAIL.n498 VTAIL.n485 0.155672
R833 VTAIL.n505 VTAIL.n485 0.155672
R834 VTAIL.n506 VTAIL.n505 0.155672
R835 VTAIL.n506 VTAIL.n481 0.155672
R836 VTAIL.n513 VTAIL.n481 0.155672
R837 VTAIL.n514 VTAIL.n513 0.155672
R838 VTAIL.n514 VTAIL.n477 0.155672
R839 VTAIL.n521 VTAIL.n477 0.155672
R840 VTAIL.n522 VTAIL.n521 0.155672
R841 VTAIL.n522 VTAIL.n473 0.155672
R842 VTAIL.n529 VTAIL.n473 0.155672
R843 VTAIL.n530 VTAIL.n529 0.155672
R844 VTAIL.n29 VTAIL.n21 0.155672
R845 VTAIL.n30 VTAIL.n29 0.155672
R846 VTAIL.n30 VTAIL.n17 0.155672
R847 VTAIL.n37 VTAIL.n17 0.155672
R848 VTAIL.n38 VTAIL.n37 0.155672
R849 VTAIL.n38 VTAIL.n13 0.155672
R850 VTAIL.n45 VTAIL.n13 0.155672
R851 VTAIL.n46 VTAIL.n45 0.155672
R852 VTAIL.n46 VTAIL.n9 0.155672
R853 VTAIL.n53 VTAIL.n9 0.155672
R854 VTAIL.n54 VTAIL.n53 0.155672
R855 VTAIL.n54 VTAIL.n5 0.155672
R856 VTAIL.n61 VTAIL.n5 0.155672
R857 VTAIL.n62 VTAIL.n61 0.155672
R858 VTAIL.n95 VTAIL.n87 0.155672
R859 VTAIL.n96 VTAIL.n95 0.155672
R860 VTAIL.n96 VTAIL.n83 0.155672
R861 VTAIL.n103 VTAIL.n83 0.155672
R862 VTAIL.n104 VTAIL.n103 0.155672
R863 VTAIL.n104 VTAIL.n79 0.155672
R864 VTAIL.n111 VTAIL.n79 0.155672
R865 VTAIL.n112 VTAIL.n111 0.155672
R866 VTAIL.n112 VTAIL.n75 0.155672
R867 VTAIL.n119 VTAIL.n75 0.155672
R868 VTAIL.n120 VTAIL.n119 0.155672
R869 VTAIL.n120 VTAIL.n71 0.155672
R870 VTAIL.n127 VTAIL.n71 0.155672
R871 VTAIL.n128 VTAIL.n127 0.155672
R872 VTAIL.n163 VTAIL.n155 0.155672
R873 VTAIL.n164 VTAIL.n163 0.155672
R874 VTAIL.n164 VTAIL.n151 0.155672
R875 VTAIL.n171 VTAIL.n151 0.155672
R876 VTAIL.n172 VTAIL.n171 0.155672
R877 VTAIL.n172 VTAIL.n147 0.155672
R878 VTAIL.n179 VTAIL.n147 0.155672
R879 VTAIL.n180 VTAIL.n179 0.155672
R880 VTAIL.n180 VTAIL.n143 0.155672
R881 VTAIL.n187 VTAIL.n143 0.155672
R882 VTAIL.n188 VTAIL.n187 0.155672
R883 VTAIL.n188 VTAIL.n139 0.155672
R884 VTAIL.n195 VTAIL.n139 0.155672
R885 VTAIL.n196 VTAIL.n195 0.155672
R886 VTAIL.n464 VTAIL.n463 0.155672
R887 VTAIL.n463 VTAIL.n407 0.155672
R888 VTAIL.n456 VTAIL.n407 0.155672
R889 VTAIL.n456 VTAIL.n455 0.155672
R890 VTAIL.n455 VTAIL.n411 0.155672
R891 VTAIL.n448 VTAIL.n411 0.155672
R892 VTAIL.n448 VTAIL.n447 0.155672
R893 VTAIL.n447 VTAIL.n415 0.155672
R894 VTAIL.n440 VTAIL.n415 0.155672
R895 VTAIL.n440 VTAIL.n439 0.155672
R896 VTAIL.n439 VTAIL.n419 0.155672
R897 VTAIL.n432 VTAIL.n419 0.155672
R898 VTAIL.n432 VTAIL.n431 0.155672
R899 VTAIL.n431 VTAIL.n423 0.155672
R900 VTAIL.n396 VTAIL.n395 0.155672
R901 VTAIL.n395 VTAIL.n339 0.155672
R902 VTAIL.n388 VTAIL.n339 0.155672
R903 VTAIL.n388 VTAIL.n387 0.155672
R904 VTAIL.n387 VTAIL.n343 0.155672
R905 VTAIL.n380 VTAIL.n343 0.155672
R906 VTAIL.n380 VTAIL.n379 0.155672
R907 VTAIL.n379 VTAIL.n347 0.155672
R908 VTAIL.n372 VTAIL.n347 0.155672
R909 VTAIL.n372 VTAIL.n371 0.155672
R910 VTAIL.n371 VTAIL.n351 0.155672
R911 VTAIL.n364 VTAIL.n351 0.155672
R912 VTAIL.n364 VTAIL.n363 0.155672
R913 VTAIL.n363 VTAIL.n355 0.155672
R914 VTAIL.n330 VTAIL.n329 0.155672
R915 VTAIL.n329 VTAIL.n273 0.155672
R916 VTAIL.n322 VTAIL.n273 0.155672
R917 VTAIL.n322 VTAIL.n321 0.155672
R918 VTAIL.n321 VTAIL.n277 0.155672
R919 VTAIL.n314 VTAIL.n277 0.155672
R920 VTAIL.n314 VTAIL.n313 0.155672
R921 VTAIL.n313 VTAIL.n281 0.155672
R922 VTAIL.n306 VTAIL.n281 0.155672
R923 VTAIL.n306 VTAIL.n305 0.155672
R924 VTAIL.n305 VTAIL.n285 0.155672
R925 VTAIL.n298 VTAIL.n285 0.155672
R926 VTAIL.n298 VTAIL.n297 0.155672
R927 VTAIL.n297 VTAIL.n289 0.155672
R928 VTAIL.n262 VTAIL.n261 0.155672
R929 VTAIL.n261 VTAIL.n205 0.155672
R930 VTAIL.n254 VTAIL.n205 0.155672
R931 VTAIL.n254 VTAIL.n253 0.155672
R932 VTAIL.n253 VTAIL.n209 0.155672
R933 VTAIL.n246 VTAIL.n209 0.155672
R934 VTAIL.n246 VTAIL.n245 0.155672
R935 VTAIL.n245 VTAIL.n213 0.155672
R936 VTAIL.n238 VTAIL.n213 0.155672
R937 VTAIL.n238 VTAIL.n237 0.155672
R938 VTAIL.n237 VTAIL.n217 0.155672
R939 VTAIL.n230 VTAIL.n217 0.155672
R940 VTAIL.n230 VTAIL.n229 0.155672
R941 VTAIL.n229 VTAIL.n221 0.155672
R942 VTAIL VTAIL.n1 0.0586897
R943 VDD1 VDD1.n0 79.4864
R944 VDD1.n3 VDD1.n2 79.3727
R945 VDD1.n3 VDD1.n1 79.3727
R946 VDD1.n5 VDD1.n4 77.8754
R947 VDD1.n5 VDD1.n3 48.6
R948 VDD1.n4 VDD1.t4 2.71151
R949 VDD1.n4 VDD1.t7 2.71151
R950 VDD1.n0 VDD1.t1 2.71151
R951 VDD1.n0 VDD1.t6 2.71151
R952 VDD1.n2 VDD1.t2 2.71151
R953 VDD1.n2 VDD1.t0 2.71151
R954 VDD1.n1 VDD1.t3 2.71151
R955 VDD1.n1 VDD1.t5 2.71151
R956 VDD1 VDD1.n5 1.49403
R957 VN.n64 VN.n63 161.3
R958 VN.n62 VN.n34 161.3
R959 VN.n61 VN.n60 161.3
R960 VN.n59 VN.n35 161.3
R961 VN.n58 VN.n57 161.3
R962 VN.n56 VN.n36 161.3
R963 VN.n55 VN.n54 161.3
R964 VN.n53 VN.n52 161.3
R965 VN.n51 VN.n38 161.3
R966 VN.n50 VN.n49 161.3
R967 VN.n48 VN.n39 161.3
R968 VN.n47 VN.n46 161.3
R969 VN.n45 VN.n40 161.3
R970 VN.n44 VN.n43 161.3
R971 VN.n31 VN.n30 161.3
R972 VN.n29 VN.n1 161.3
R973 VN.n28 VN.n27 161.3
R974 VN.n26 VN.n2 161.3
R975 VN.n25 VN.n24 161.3
R976 VN.n23 VN.n3 161.3
R977 VN.n22 VN.n21 161.3
R978 VN.n20 VN.n19 161.3
R979 VN.n18 VN.n5 161.3
R980 VN.n17 VN.n16 161.3
R981 VN.n15 VN.n6 161.3
R982 VN.n14 VN.n13 161.3
R983 VN.n12 VN.n7 161.3
R984 VN.n11 VN.n10 161.3
R985 VN.n42 VN.t4 121.709
R986 VN.n9 VN.t3 121.709
R987 VN.n8 VN.t5 88.3672
R988 VN.n4 VN.t2 88.3672
R989 VN.n0 VN.t0 88.3672
R990 VN.n41 VN.t7 88.3672
R991 VN.n37 VN.t1 88.3672
R992 VN.n33 VN.t6 88.3672
R993 VN.n32 VN.n0 70.4938
R994 VN.n65 VN.n33 70.4938
R995 VN.n9 VN.n8 59.4932
R996 VN.n42 VN.n41 59.4932
R997 VN VN.n65 54.3692
R998 VN.n28 VN.n2 50.2061
R999 VN.n61 VN.n35 50.2061
R1000 VN.n13 VN.n6 40.4934
R1001 VN.n17 VN.n6 40.4934
R1002 VN.n46 VN.n39 40.4934
R1003 VN.n50 VN.n39 40.4934
R1004 VN.n24 VN.n2 30.7807
R1005 VN.n57 VN.n35 30.7807
R1006 VN.n12 VN.n11 24.4675
R1007 VN.n13 VN.n12 24.4675
R1008 VN.n18 VN.n17 24.4675
R1009 VN.n19 VN.n18 24.4675
R1010 VN.n23 VN.n22 24.4675
R1011 VN.n24 VN.n23 24.4675
R1012 VN.n29 VN.n28 24.4675
R1013 VN.n30 VN.n29 24.4675
R1014 VN.n46 VN.n45 24.4675
R1015 VN.n45 VN.n44 24.4675
R1016 VN.n57 VN.n56 24.4675
R1017 VN.n56 VN.n55 24.4675
R1018 VN.n52 VN.n51 24.4675
R1019 VN.n51 VN.n50 24.4675
R1020 VN.n63 VN.n62 24.4675
R1021 VN.n62 VN.n61 24.4675
R1022 VN.n30 VN.n0 19.5741
R1023 VN.n63 VN.n33 19.5741
R1024 VN.n11 VN.n8 14.6807
R1025 VN.n19 VN.n4 14.6807
R1026 VN.n44 VN.n41 14.6807
R1027 VN.n52 VN.n37 14.6807
R1028 VN.n22 VN.n4 9.7873
R1029 VN.n55 VN.n37 9.7873
R1030 VN.n10 VN.n9 3.92587
R1031 VN.n43 VN.n42 3.92587
R1032 VN.n65 VN.n64 0.354971
R1033 VN.n32 VN.n31 0.354971
R1034 VN VN.n32 0.26696
R1035 VN.n64 VN.n34 0.189894
R1036 VN.n60 VN.n34 0.189894
R1037 VN.n60 VN.n59 0.189894
R1038 VN.n59 VN.n58 0.189894
R1039 VN.n58 VN.n36 0.189894
R1040 VN.n54 VN.n36 0.189894
R1041 VN.n54 VN.n53 0.189894
R1042 VN.n53 VN.n38 0.189894
R1043 VN.n49 VN.n38 0.189894
R1044 VN.n49 VN.n48 0.189894
R1045 VN.n48 VN.n47 0.189894
R1046 VN.n47 VN.n40 0.189894
R1047 VN.n43 VN.n40 0.189894
R1048 VN.n10 VN.n7 0.189894
R1049 VN.n14 VN.n7 0.189894
R1050 VN.n15 VN.n14 0.189894
R1051 VN.n16 VN.n15 0.189894
R1052 VN.n16 VN.n5 0.189894
R1053 VN.n20 VN.n5 0.189894
R1054 VN.n21 VN.n20 0.189894
R1055 VN.n21 VN.n3 0.189894
R1056 VN.n25 VN.n3 0.189894
R1057 VN.n26 VN.n25 0.189894
R1058 VN.n27 VN.n26 0.189894
R1059 VN.n27 VN.n1 0.189894
R1060 VN.n31 VN.n1 0.189894
R1061 VDD2.n2 VDD2.n1 79.3727
R1062 VDD2.n2 VDD2.n0 79.3727
R1063 VDD2 VDD2.n5 79.369
R1064 VDD2.n4 VDD2.n3 77.8765
R1065 VDD2.n4 VDD2.n2 48.017
R1066 VDD2.n5 VDD2.t0 2.71151
R1067 VDD2.n5 VDD2.t3 2.71151
R1068 VDD2.n3 VDD2.t1 2.71151
R1069 VDD2.n3 VDD2.t6 2.71151
R1070 VDD2.n1 VDD2.t5 2.71151
R1071 VDD2.n1 VDD2.t7 2.71151
R1072 VDD2.n0 VDD2.t4 2.71151
R1073 VDD2.n0 VDD2.t2 2.71151
R1074 VDD2 VDD2.n4 1.61041
R1075 B.n642 B.n83 585
R1076 B.n644 B.n643 585
R1077 B.n645 B.n82 585
R1078 B.n647 B.n646 585
R1079 B.n648 B.n81 585
R1080 B.n650 B.n649 585
R1081 B.n651 B.n80 585
R1082 B.n653 B.n652 585
R1083 B.n654 B.n79 585
R1084 B.n656 B.n655 585
R1085 B.n657 B.n78 585
R1086 B.n659 B.n658 585
R1087 B.n660 B.n77 585
R1088 B.n662 B.n661 585
R1089 B.n663 B.n76 585
R1090 B.n665 B.n664 585
R1091 B.n666 B.n75 585
R1092 B.n668 B.n667 585
R1093 B.n669 B.n74 585
R1094 B.n671 B.n670 585
R1095 B.n672 B.n73 585
R1096 B.n674 B.n673 585
R1097 B.n675 B.n72 585
R1098 B.n677 B.n676 585
R1099 B.n678 B.n71 585
R1100 B.n680 B.n679 585
R1101 B.n681 B.n70 585
R1102 B.n683 B.n682 585
R1103 B.n684 B.n69 585
R1104 B.n686 B.n685 585
R1105 B.n687 B.n68 585
R1106 B.n689 B.n688 585
R1107 B.n690 B.n67 585
R1108 B.n692 B.n691 585
R1109 B.n693 B.n66 585
R1110 B.n695 B.n694 585
R1111 B.n696 B.n65 585
R1112 B.n698 B.n697 585
R1113 B.n699 B.n64 585
R1114 B.n701 B.n700 585
R1115 B.n702 B.n63 585
R1116 B.n704 B.n703 585
R1117 B.n706 B.n705 585
R1118 B.n707 B.n59 585
R1119 B.n709 B.n708 585
R1120 B.n710 B.n58 585
R1121 B.n712 B.n711 585
R1122 B.n713 B.n57 585
R1123 B.n715 B.n714 585
R1124 B.n716 B.n56 585
R1125 B.n718 B.n717 585
R1126 B.n720 B.n53 585
R1127 B.n722 B.n721 585
R1128 B.n723 B.n52 585
R1129 B.n725 B.n724 585
R1130 B.n726 B.n51 585
R1131 B.n728 B.n727 585
R1132 B.n729 B.n50 585
R1133 B.n731 B.n730 585
R1134 B.n732 B.n49 585
R1135 B.n734 B.n733 585
R1136 B.n735 B.n48 585
R1137 B.n737 B.n736 585
R1138 B.n738 B.n47 585
R1139 B.n740 B.n739 585
R1140 B.n741 B.n46 585
R1141 B.n743 B.n742 585
R1142 B.n744 B.n45 585
R1143 B.n746 B.n745 585
R1144 B.n747 B.n44 585
R1145 B.n749 B.n748 585
R1146 B.n750 B.n43 585
R1147 B.n752 B.n751 585
R1148 B.n753 B.n42 585
R1149 B.n755 B.n754 585
R1150 B.n756 B.n41 585
R1151 B.n758 B.n757 585
R1152 B.n759 B.n40 585
R1153 B.n761 B.n760 585
R1154 B.n762 B.n39 585
R1155 B.n764 B.n763 585
R1156 B.n765 B.n38 585
R1157 B.n767 B.n766 585
R1158 B.n768 B.n37 585
R1159 B.n770 B.n769 585
R1160 B.n771 B.n36 585
R1161 B.n773 B.n772 585
R1162 B.n774 B.n35 585
R1163 B.n776 B.n775 585
R1164 B.n777 B.n34 585
R1165 B.n779 B.n778 585
R1166 B.n780 B.n33 585
R1167 B.n782 B.n781 585
R1168 B.n641 B.n640 585
R1169 B.n639 B.n84 585
R1170 B.n638 B.n637 585
R1171 B.n636 B.n85 585
R1172 B.n635 B.n634 585
R1173 B.n633 B.n86 585
R1174 B.n632 B.n631 585
R1175 B.n630 B.n87 585
R1176 B.n629 B.n628 585
R1177 B.n627 B.n88 585
R1178 B.n626 B.n625 585
R1179 B.n624 B.n89 585
R1180 B.n623 B.n622 585
R1181 B.n621 B.n90 585
R1182 B.n620 B.n619 585
R1183 B.n618 B.n91 585
R1184 B.n617 B.n616 585
R1185 B.n615 B.n92 585
R1186 B.n614 B.n613 585
R1187 B.n612 B.n93 585
R1188 B.n611 B.n610 585
R1189 B.n609 B.n94 585
R1190 B.n608 B.n607 585
R1191 B.n606 B.n95 585
R1192 B.n605 B.n604 585
R1193 B.n603 B.n96 585
R1194 B.n602 B.n601 585
R1195 B.n600 B.n97 585
R1196 B.n599 B.n598 585
R1197 B.n597 B.n98 585
R1198 B.n596 B.n595 585
R1199 B.n594 B.n99 585
R1200 B.n593 B.n592 585
R1201 B.n591 B.n100 585
R1202 B.n590 B.n589 585
R1203 B.n588 B.n101 585
R1204 B.n587 B.n586 585
R1205 B.n585 B.n102 585
R1206 B.n584 B.n583 585
R1207 B.n582 B.n103 585
R1208 B.n581 B.n580 585
R1209 B.n579 B.n104 585
R1210 B.n578 B.n577 585
R1211 B.n576 B.n105 585
R1212 B.n575 B.n574 585
R1213 B.n573 B.n106 585
R1214 B.n572 B.n571 585
R1215 B.n570 B.n107 585
R1216 B.n569 B.n568 585
R1217 B.n567 B.n108 585
R1218 B.n566 B.n565 585
R1219 B.n564 B.n109 585
R1220 B.n563 B.n562 585
R1221 B.n561 B.n110 585
R1222 B.n560 B.n559 585
R1223 B.n558 B.n111 585
R1224 B.n557 B.n556 585
R1225 B.n555 B.n112 585
R1226 B.n554 B.n553 585
R1227 B.n552 B.n113 585
R1228 B.n551 B.n550 585
R1229 B.n549 B.n114 585
R1230 B.n548 B.n547 585
R1231 B.n546 B.n115 585
R1232 B.n545 B.n544 585
R1233 B.n543 B.n116 585
R1234 B.n542 B.n541 585
R1235 B.n540 B.n117 585
R1236 B.n539 B.n538 585
R1237 B.n537 B.n118 585
R1238 B.n536 B.n535 585
R1239 B.n534 B.n119 585
R1240 B.n533 B.n532 585
R1241 B.n531 B.n120 585
R1242 B.n530 B.n529 585
R1243 B.n528 B.n121 585
R1244 B.n527 B.n526 585
R1245 B.n525 B.n122 585
R1246 B.n524 B.n523 585
R1247 B.n522 B.n123 585
R1248 B.n521 B.n520 585
R1249 B.n519 B.n124 585
R1250 B.n518 B.n517 585
R1251 B.n516 B.n125 585
R1252 B.n515 B.n514 585
R1253 B.n513 B.n126 585
R1254 B.n512 B.n511 585
R1255 B.n510 B.n127 585
R1256 B.n509 B.n508 585
R1257 B.n507 B.n128 585
R1258 B.n506 B.n505 585
R1259 B.n504 B.n129 585
R1260 B.n503 B.n502 585
R1261 B.n501 B.n130 585
R1262 B.n500 B.n499 585
R1263 B.n498 B.n131 585
R1264 B.n497 B.n496 585
R1265 B.n495 B.n132 585
R1266 B.n494 B.n493 585
R1267 B.n492 B.n133 585
R1268 B.n491 B.n490 585
R1269 B.n489 B.n134 585
R1270 B.n488 B.n487 585
R1271 B.n486 B.n135 585
R1272 B.n485 B.n484 585
R1273 B.n483 B.n136 585
R1274 B.n482 B.n481 585
R1275 B.n480 B.n137 585
R1276 B.n479 B.n478 585
R1277 B.n477 B.n138 585
R1278 B.n476 B.n475 585
R1279 B.n474 B.n139 585
R1280 B.n473 B.n472 585
R1281 B.n471 B.n140 585
R1282 B.n470 B.n469 585
R1283 B.n468 B.n141 585
R1284 B.n467 B.n466 585
R1285 B.n465 B.n142 585
R1286 B.n464 B.n463 585
R1287 B.n462 B.n143 585
R1288 B.n461 B.n460 585
R1289 B.n459 B.n144 585
R1290 B.n458 B.n457 585
R1291 B.n317 B.n316 585
R1292 B.n318 B.n195 585
R1293 B.n320 B.n319 585
R1294 B.n321 B.n194 585
R1295 B.n323 B.n322 585
R1296 B.n324 B.n193 585
R1297 B.n326 B.n325 585
R1298 B.n327 B.n192 585
R1299 B.n329 B.n328 585
R1300 B.n330 B.n191 585
R1301 B.n332 B.n331 585
R1302 B.n333 B.n190 585
R1303 B.n335 B.n334 585
R1304 B.n336 B.n189 585
R1305 B.n338 B.n337 585
R1306 B.n339 B.n188 585
R1307 B.n341 B.n340 585
R1308 B.n342 B.n187 585
R1309 B.n344 B.n343 585
R1310 B.n345 B.n186 585
R1311 B.n347 B.n346 585
R1312 B.n348 B.n185 585
R1313 B.n350 B.n349 585
R1314 B.n351 B.n184 585
R1315 B.n353 B.n352 585
R1316 B.n354 B.n183 585
R1317 B.n356 B.n355 585
R1318 B.n357 B.n182 585
R1319 B.n359 B.n358 585
R1320 B.n360 B.n181 585
R1321 B.n362 B.n361 585
R1322 B.n363 B.n180 585
R1323 B.n365 B.n364 585
R1324 B.n366 B.n179 585
R1325 B.n368 B.n367 585
R1326 B.n369 B.n178 585
R1327 B.n371 B.n370 585
R1328 B.n372 B.n177 585
R1329 B.n374 B.n373 585
R1330 B.n375 B.n176 585
R1331 B.n377 B.n376 585
R1332 B.n378 B.n173 585
R1333 B.n381 B.n380 585
R1334 B.n382 B.n172 585
R1335 B.n384 B.n383 585
R1336 B.n385 B.n171 585
R1337 B.n387 B.n386 585
R1338 B.n388 B.n170 585
R1339 B.n390 B.n389 585
R1340 B.n391 B.n169 585
R1341 B.n393 B.n392 585
R1342 B.n395 B.n394 585
R1343 B.n396 B.n165 585
R1344 B.n398 B.n397 585
R1345 B.n399 B.n164 585
R1346 B.n401 B.n400 585
R1347 B.n402 B.n163 585
R1348 B.n404 B.n403 585
R1349 B.n405 B.n162 585
R1350 B.n407 B.n406 585
R1351 B.n408 B.n161 585
R1352 B.n410 B.n409 585
R1353 B.n411 B.n160 585
R1354 B.n413 B.n412 585
R1355 B.n414 B.n159 585
R1356 B.n416 B.n415 585
R1357 B.n417 B.n158 585
R1358 B.n419 B.n418 585
R1359 B.n420 B.n157 585
R1360 B.n422 B.n421 585
R1361 B.n423 B.n156 585
R1362 B.n425 B.n424 585
R1363 B.n426 B.n155 585
R1364 B.n428 B.n427 585
R1365 B.n429 B.n154 585
R1366 B.n431 B.n430 585
R1367 B.n432 B.n153 585
R1368 B.n434 B.n433 585
R1369 B.n435 B.n152 585
R1370 B.n437 B.n436 585
R1371 B.n438 B.n151 585
R1372 B.n440 B.n439 585
R1373 B.n441 B.n150 585
R1374 B.n443 B.n442 585
R1375 B.n444 B.n149 585
R1376 B.n446 B.n445 585
R1377 B.n447 B.n148 585
R1378 B.n449 B.n448 585
R1379 B.n450 B.n147 585
R1380 B.n452 B.n451 585
R1381 B.n453 B.n146 585
R1382 B.n455 B.n454 585
R1383 B.n456 B.n145 585
R1384 B.n315 B.n196 585
R1385 B.n314 B.n313 585
R1386 B.n312 B.n197 585
R1387 B.n311 B.n310 585
R1388 B.n309 B.n198 585
R1389 B.n308 B.n307 585
R1390 B.n306 B.n199 585
R1391 B.n305 B.n304 585
R1392 B.n303 B.n200 585
R1393 B.n302 B.n301 585
R1394 B.n300 B.n201 585
R1395 B.n299 B.n298 585
R1396 B.n297 B.n202 585
R1397 B.n296 B.n295 585
R1398 B.n294 B.n203 585
R1399 B.n293 B.n292 585
R1400 B.n291 B.n204 585
R1401 B.n290 B.n289 585
R1402 B.n288 B.n205 585
R1403 B.n287 B.n286 585
R1404 B.n285 B.n206 585
R1405 B.n284 B.n283 585
R1406 B.n282 B.n207 585
R1407 B.n281 B.n280 585
R1408 B.n279 B.n208 585
R1409 B.n278 B.n277 585
R1410 B.n276 B.n209 585
R1411 B.n275 B.n274 585
R1412 B.n273 B.n210 585
R1413 B.n272 B.n271 585
R1414 B.n270 B.n211 585
R1415 B.n269 B.n268 585
R1416 B.n267 B.n212 585
R1417 B.n266 B.n265 585
R1418 B.n264 B.n213 585
R1419 B.n263 B.n262 585
R1420 B.n261 B.n214 585
R1421 B.n260 B.n259 585
R1422 B.n258 B.n215 585
R1423 B.n257 B.n256 585
R1424 B.n255 B.n216 585
R1425 B.n254 B.n253 585
R1426 B.n252 B.n217 585
R1427 B.n251 B.n250 585
R1428 B.n249 B.n218 585
R1429 B.n248 B.n247 585
R1430 B.n246 B.n219 585
R1431 B.n245 B.n244 585
R1432 B.n243 B.n220 585
R1433 B.n242 B.n241 585
R1434 B.n240 B.n221 585
R1435 B.n239 B.n238 585
R1436 B.n237 B.n222 585
R1437 B.n236 B.n235 585
R1438 B.n234 B.n223 585
R1439 B.n233 B.n232 585
R1440 B.n231 B.n224 585
R1441 B.n230 B.n229 585
R1442 B.n228 B.n225 585
R1443 B.n227 B.n226 585
R1444 B.n2 B.n0 585
R1445 B.n873 B.n1 585
R1446 B.n872 B.n871 585
R1447 B.n870 B.n3 585
R1448 B.n869 B.n868 585
R1449 B.n867 B.n4 585
R1450 B.n866 B.n865 585
R1451 B.n864 B.n5 585
R1452 B.n863 B.n862 585
R1453 B.n861 B.n6 585
R1454 B.n860 B.n859 585
R1455 B.n858 B.n7 585
R1456 B.n857 B.n856 585
R1457 B.n855 B.n8 585
R1458 B.n854 B.n853 585
R1459 B.n852 B.n9 585
R1460 B.n851 B.n850 585
R1461 B.n849 B.n10 585
R1462 B.n848 B.n847 585
R1463 B.n846 B.n11 585
R1464 B.n845 B.n844 585
R1465 B.n843 B.n12 585
R1466 B.n842 B.n841 585
R1467 B.n840 B.n13 585
R1468 B.n839 B.n838 585
R1469 B.n837 B.n14 585
R1470 B.n836 B.n835 585
R1471 B.n834 B.n15 585
R1472 B.n833 B.n832 585
R1473 B.n831 B.n16 585
R1474 B.n830 B.n829 585
R1475 B.n828 B.n17 585
R1476 B.n827 B.n826 585
R1477 B.n825 B.n18 585
R1478 B.n824 B.n823 585
R1479 B.n822 B.n19 585
R1480 B.n821 B.n820 585
R1481 B.n819 B.n20 585
R1482 B.n818 B.n817 585
R1483 B.n816 B.n21 585
R1484 B.n815 B.n814 585
R1485 B.n813 B.n22 585
R1486 B.n812 B.n811 585
R1487 B.n810 B.n23 585
R1488 B.n809 B.n808 585
R1489 B.n807 B.n24 585
R1490 B.n806 B.n805 585
R1491 B.n804 B.n25 585
R1492 B.n803 B.n802 585
R1493 B.n801 B.n26 585
R1494 B.n800 B.n799 585
R1495 B.n798 B.n27 585
R1496 B.n797 B.n796 585
R1497 B.n795 B.n28 585
R1498 B.n794 B.n793 585
R1499 B.n792 B.n29 585
R1500 B.n791 B.n790 585
R1501 B.n789 B.n30 585
R1502 B.n788 B.n787 585
R1503 B.n786 B.n31 585
R1504 B.n785 B.n784 585
R1505 B.n783 B.n32 585
R1506 B.n875 B.n874 585
R1507 B.n316 B.n315 487.695
R1508 B.n783 B.n782 487.695
R1509 B.n458 B.n145 487.695
R1510 B.n640 B.n83 487.695
R1511 B.n166 B.t11 445.154
R1512 B.n60 B.t1 445.154
R1513 B.n174 B.t8 445.154
R1514 B.n54 B.t4 445.154
R1515 B.n167 B.t10 375.337
R1516 B.n61 B.t2 375.337
R1517 B.n175 B.t7 375.337
R1518 B.n55 B.t5 375.337
R1519 B.n166 B.t9 297.241
R1520 B.n174 B.t6 297.241
R1521 B.n54 B.t3 297.241
R1522 B.n60 B.t0 297.241
R1523 B.n315 B.n314 163.367
R1524 B.n314 B.n197 163.367
R1525 B.n310 B.n197 163.367
R1526 B.n310 B.n309 163.367
R1527 B.n309 B.n308 163.367
R1528 B.n308 B.n199 163.367
R1529 B.n304 B.n199 163.367
R1530 B.n304 B.n303 163.367
R1531 B.n303 B.n302 163.367
R1532 B.n302 B.n201 163.367
R1533 B.n298 B.n201 163.367
R1534 B.n298 B.n297 163.367
R1535 B.n297 B.n296 163.367
R1536 B.n296 B.n203 163.367
R1537 B.n292 B.n203 163.367
R1538 B.n292 B.n291 163.367
R1539 B.n291 B.n290 163.367
R1540 B.n290 B.n205 163.367
R1541 B.n286 B.n205 163.367
R1542 B.n286 B.n285 163.367
R1543 B.n285 B.n284 163.367
R1544 B.n284 B.n207 163.367
R1545 B.n280 B.n207 163.367
R1546 B.n280 B.n279 163.367
R1547 B.n279 B.n278 163.367
R1548 B.n278 B.n209 163.367
R1549 B.n274 B.n209 163.367
R1550 B.n274 B.n273 163.367
R1551 B.n273 B.n272 163.367
R1552 B.n272 B.n211 163.367
R1553 B.n268 B.n211 163.367
R1554 B.n268 B.n267 163.367
R1555 B.n267 B.n266 163.367
R1556 B.n266 B.n213 163.367
R1557 B.n262 B.n213 163.367
R1558 B.n262 B.n261 163.367
R1559 B.n261 B.n260 163.367
R1560 B.n260 B.n215 163.367
R1561 B.n256 B.n215 163.367
R1562 B.n256 B.n255 163.367
R1563 B.n255 B.n254 163.367
R1564 B.n254 B.n217 163.367
R1565 B.n250 B.n217 163.367
R1566 B.n250 B.n249 163.367
R1567 B.n249 B.n248 163.367
R1568 B.n248 B.n219 163.367
R1569 B.n244 B.n219 163.367
R1570 B.n244 B.n243 163.367
R1571 B.n243 B.n242 163.367
R1572 B.n242 B.n221 163.367
R1573 B.n238 B.n221 163.367
R1574 B.n238 B.n237 163.367
R1575 B.n237 B.n236 163.367
R1576 B.n236 B.n223 163.367
R1577 B.n232 B.n223 163.367
R1578 B.n232 B.n231 163.367
R1579 B.n231 B.n230 163.367
R1580 B.n230 B.n225 163.367
R1581 B.n226 B.n225 163.367
R1582 B.n226 B.n2 163.367
R1583 B.n874 B.n2 163.367
R1584 B.n874 B.n873 163.367
R1585 B.n873 B.n872 163.367
R1586 B.n872 B.n3 163.367
R1587 B.n868 B.n3 163.367
R1588 B.n868 B.n867 163.367
R1589 B.n867 B.n866 163.367
R1590 B.n866 B.n5 163.367
R1591 B.n862 B.n5 163.367
R1592 B.n862 B.n861 163.367
R1593 B.n861 B.n860 163.367
R1594 B.n860 B.n7 163.367
R1595 B.n856 B.n7 163.367
R1596 B.n856 B.n855 163.367
R1597 B.n855 B.n854 163.367
R1598 B.n854 B.n9 163.367
R1599 B.n850 B.n9 163.367
R1600 B.n850 B.n849 163.367
R1601 B.n849 B.n848 163.367
R1602 B.n848 B.n11 163.367
R1603 B.n844 B.n11 163.367
R1604 B.n844 B.n843 163.367
R1605 B.n843 B.n842 163.367
R1606 B.n842 B.n13 163.367
R1607 B.n838 B.n13 163.367
R1608 B.n838 B.n837 163.367
R1609 B.n837 B.n836 163.367
R1610 B.n836 B.n15 163.367
R1611 B.n832 B.n15 163.367
R1612 B.n832 B.n831 163.367
R1613 B.n831 B.n830 163.367
R1614 B.n830 B.n17 163.367
R1615 B.n826 B.n17 163.367
R1616 B.n826 B.n825 163.367
R1617 B.n825 B.n824 163.367
R1618 B.n824 B.n19 163.367
R1619 B.n820 B.n19 163.367
R1620 B.n820 B.n819 163.367
R1621 B.n819 B.n818 163.367
R1622 B.n818 B.n21 163.367
R1623 B.n814 B.n21 163.367
R1624 B.n814 B.n813 163.367
R1625 B.n813 B.n812 163.367
R1626 B.n812 B.n23 163.367
R1627 B.n808 B.n23 163.367
R1628 B.n808 B.n807 163.367
R1629 B.n807 B.n806 163.367
R1630 B.n806 B.n25 163.367
R1631 B.n802 B.n25 163.367
R1632 B.n802 B.n801 163.367
R1633 B.n801 B.n800 163.367
R1634 B.n800 B.n27 163.367
R1635 B.n796 B.n27 163.367
R1636 B.n796 B.n795 163.367
R1637 B.n795 B.n794 163.367
R1638 B.n794 B.n29 163.367
R1639 B.n790 B.n29 163.367
R1640 B.n790 B.n789 163.367
R1641 B.n789 B.n788 163.367
R1642 B.n788 B.n31 163.367
R1643 B.n784 B.n31 163.367
R1644 B.n784 B.n783 163.367
R1645 B.n316 B.n195 163.367
R1646 B.n320 B.n195 163.367
R1647 B.n321 B.n320 163.367
R1648 B.n322 B.n321 163.367
R1649 B.n322 B.n193 163.367
R1650 B.n326 B.n193 163.367
R1651 B.n327 B.n326 163.367
R1652 B.n328 B.n327 163.367
R1653 B.n328 B.n191 163.367
R1654 B.n332 B.n191 163.367
R1655 B.n333 B.n332 163.367
R1656 B.n334 B.n333 163.367
R1657 B.n334 B.n189 163.367
R1658 B.n338 B.n189 163.367
R1659 B.n339 B.n338 163.367
R1660 B.n340 B.n339 163.367
R1661 B.n340 B.n187 163.367
R1662 B.n344 B.n187 163.367
R1663 B.n345 B.n344 163.367
R1664 B.n346 B.n345 163.367
R1665 B.n346 B.n185 163.367
R1666 B.n350 B.n185 163.367
R1667 B.n351 B.n350 163.367
R1668 B.n352 B.n351 163.367
R1669 B.n352 B.n183 163.367
R1670 B.n356 B.n183 163.367
R1671 B.n357 B.n356 163.367
R1672 B.n358 B.n357 163.367
R1673 B.n358 B.n181 163.367
R1674 B.n362 B.n181 163.367
R1675 B.n363 B.n362 163.367
R1676 B.n364 B.n363 163.367
R1677 B.n364 B.n179 163.367
R1678 B.n368 B.n179 163.367
R1679 B.n369 B.n368 163.367
R1680 B.n370 B.n369 163.367
R1681 B.n370 B.n177 163.367
R1682 B.n374 B.n177 163.367
R1683 B.n375 B.n374 163.367
R1684 B.n376 B.n375 163.367
R1685 B.n376 B.n173 163.367
R1686 B.n381 B.n173 163.367
R1687 B.n382 B.n381 163.367
R1688 B.n383 B.n382 163.367
R1689 B.n383 B.n171 163.367
R1690 B.n387 B.n171 163.367
R1691 B.n388 B.n387 163.367
R1692 B.n389 B.n388 163.367
R1693 B.n389 B.n169 163.367
R1694 B.n393 B.n169 163.367
R1695 B.n394 B.n393 163.367
R1696 B.n394 B.n165 163.367
R1697 B.n398 B.n165 163.367
R1698 B.n399 B.n398 163.367
R1699 B.n400 B.n399 163.367
R1700 B.n400 B.n163 163.367
R1701 B.n404 B.n163 163.367
R1702 B.n405 B.n404 163.367
R1703 B.n406 B.n405 163.367
R1704 B.n406 B.n161 163.367
R1705 B.n410 B.n161 163.367
R1706 B.n411 B.n410 163.367
R1707 B.n412 B.n411 163.367
R1708 B.n412 B.n159 163.367
R1709 B.n416 B.n159 163.367
R1710 B.n417 B.n416 163.367
R1711 B.n418 B.n417 163.367
R1712 B.n418 B.n157 163.367
R1713 B.n422 B.n157 163.367
R1714 B.n423 B.n422 163.367
R1715 B.n424 B.n423 163.367
R1716 B.n424 B.n155 163.367
R1717 B.n428 B.n155 163.367
R1718 B.n429 B.n428 163.367
R1719 B.n430 B.n429 163.367
R1720 B.n430 B.n153 163.367
R1721 B.n434 B.n153 163.367
R1722 B.n435 B.n434 163.367
R1723 B.n436 B.n435 163.367
R1724 B.n436 B.n151 163.367
R1725 B.n440 B.n151 163.367
R1726 B.n441 B.n440 163.367
R1727 B.n442 B.n441 163.367
R1728 B.n442 B.n149 163.367
R1729 B.n446 B.n149 163.367
R1730 B.n447 B.n446 163.367
R1731 B.n448 B.n447 163.367
R1732 B.n448 B.n147 163.367
R1733 B.n452 B.n147 163.367
R1734 B.n453 B.n452 163.367
R1735 B.n454 B.n453 163.367
R1736 B.n454 B.n145 163.367
R1737 B.n459 B.n458 163.367
R1738 B.n460 B.n459 163.367
R1739 B.n460 B.n143 163.367
R1740 B.n464 B.n143 163.367
R1741 B.n465 B.n464 163.367
R1742 B.n466 B.n465 163.367
R1743 B.n466 B.n141 163.367
R1744 B.n470 B.n141 163.367
R1745 B.n471 B.n470 163.367
R1746 B.n472 B.n471 163.367
R1747 B.n472 B.n139 163.367
R1748 B.n476 B.n139 163.367
R1749 B.n477 B.n476 163.367
R1750 B.n478 B.n477 163.367
R1751 B.n478 B.n137 163.367
R1752 B.n482 B.n137 163.367
R1753 B.n483 B.n482 163.367
R1754 B.n484 B.n483 163.367
R1755 B.n484 B.n135 163.367
R1756 B.n488 B.n135 163.367
R1757 B.n489 B.n488 163.367
R1758 B.n490 B.n489 163.367
R1759 B.n490 B.n133 163.367
R1760 B.n494 B.n133 163.367
R1761 B.n495 B.n494 163.367
R1762 B.n496 B.n495 163.367
R1763 B.n496 B.n131 163.367
R1764 B.n500 B.n131 163.367
R1765 B.n501 B.n500 163.367
R1766 B.n502 B.n501 163.367
R1767 B.n502 B.n129 163.367
R1768 B.n506 B.n129 163.367
R1769 B.n507 B.n506 163.367
R1770 B.n508 B.n507 163.367
R1771 B.n508 B.n127 163.367
R1772 B.n512 B.n127 163.367
R1773 B.n513 B.n512 163.367
R1774 B.n514 B.n513 163.367
R1775 B.n514 B.n125 163.367
R1776 B.n518 B.n125 163.367
R1777 B.n519 B.n518 163.367
R1778 B.n520 B.n519 163.367
R1779 B.n520 B.n123 163.367
R1780 B.n524 B.n123 163.367
R1781 B.n525 B.n524 163.367
R1782 B.n526 B.n525 163.367
R1783 B.n526 B.n121 163.367
R1784 B.n530 B.n121 163.367
R1785 B.n531 B.n530 163.367
R1786 B.n532 B.n531 163.367
R1787 B.n532 B.n119 163.367
R1788 B.n536 B.n119 163.367
R1789 B.n537 B.n536 163.367
R1790 B.n538 B.n537 163.367
R1791 B.n538 B.n117 163.367
R1792 B.n542 B.n117 163.367
R1793 B.n543 B.n542 163.367
R1794 B.n544 B.n543 163.367
R1795 B.n544 B.n115 163.367
R1796 B.n548 B.n115 163.367
R1797 B.n549 B.n548 163.367
R1798 B.n550 B.n549 163.367
R1799 B.n550 B.n113 163.367
R1800 B.n554 B.n113 163.367
R1801 B.n555 B.n554 163.367
R1802 B.n556 B.n555 163.367
R1803 B.n556 B.n111 163.367
R1804 B.n560 B.n111 163.367
R1805 B.n561 B.n560 163.367
R1806 B.n562 B.n561 163.367
R1807 B.n562 B.n109 163.367
R1808 B.n566 B.n109 163.367
R1809 B.n567 B.n566 163.367
R1810 B.n568 B.n567 163.367
R1811 B.n568 B.n107 163.367
R1812 B.n572 B.n107 163.367
R1813 B.n573 B.n572 163.367
R1814 B.n574 B.n573 163.367
R1815 B.n574 B.n105 163.367
R1816 B.n578 B.n105 163.367
R1817 B.n579 B.n578 163.367
R1818 B.n580 B.n579 163.367
R1819 B.n580 B.n103 163.367
R1820 B.n584 B.n103 163.367
R1821 B.n585 B.n584 163.367
R1822 B.n586 B.n585 163.367
R1823 B.n586 B.n101 163.367
R1824 B.n590 B.n101 163.367
R1825 B.n591 B.n590 163.367
R1826 B.n592 B.n591 163.367
R1827 B.n592 B.n99 163.367
R1828 B.n596 B.n99 163.367
R1829 B.n597 B.n596 163.367
R1830 B.n598 B.n597 163.367
R1831 B.n598 B.n97 163.367
R1832 B.n602 B.n97 163.367
R1833 B.n603 B.n602 163.367
R1834 B.n604 B.n603 163.367
R1835 B.n604 B.n95 163.367
R1836 B.n608 B.n95 163.367
R1837 B.n609 B.n608 163.367
R1838 B.n610 B.n609 163.367
R1839 B.n610 B.n93 163.367
R1840 B.n614 B.n93 163.367
R1841 B.n615 B.n614 163.367
R1842 B.n616 B.n615 163.367
R1843 B.n616 B.n91 163.367
R1844 B.n620 B.n91 163.367
R1845 B.n621 B.n620 163.367
R1846 B.n622 B.n621 163.367
R1847 B.n622 B.n89 163.367
R1848 B.n626 B.n89 163.367
R1849 B.n627 B.n626 163.367
R1850 B.n628 B.n627 163.367
R1851 B.n628 B.n87 163.367
R1852 B.n632 B.n87 163.367
R1853 B.n633 B.n632 163.367
R1854 B.n634 B.n633 163.367
R1855 B.n634 B.n85 163.367
R1856 B.n638 B.n85 163.367
R1857 B.n639 B.n638 163.367
R1858 B.n640 B.n639 163.367
R1859 B.n782 B.n33 163.367
R1860 B.n778 B.n33 163.367
R1861 B.n778 B.n777 163.367
R1862 B.n777 B.n776 163.367
R1863 B.n776 B.n35 163.367
R1864 B.n772 B.n35 163.367
R1865 B.n772 B.n771 163.367
R1866 B.n771 B.n770 163.367
R1867 B.n770 B.n37 163.367
R1868 B.n766 B.n37 163.367
R1869 B.n766 B.n765 163.367
R1870 B.n765 B.n764 163.367
R1871 B.n764 B.n39 163.367
R1872 B.n760 B.n39 163.367
R1873 B.n760 B.n759 163.367
R1874 B.n759 B.n758 163.367
R1875 B.n758 B.n41 163.367
R1876 B.n754 B.n41 163.367
R1877 B.n754 B.n753 163.367
R1878 B.n753 B.n752 163.367
R1879 B.n752 B.n43 163.367
R1880 B.n748 B.n43 163.367
R1881 B.n748 B.n747 163.367
R1882 B.n747 B.n746 163.367
R1883 B.n746 B.n45 163.367
R1884 B.n742 B.n45 163.367
R1885 B.n742 B.n741 163.367
R1886 B.n741 B.n740 163.367
R1887 B.n740 B.n47 163.367
R1888 B.n736 B.n47 163.367
R1889 B.n736 B.n735 163.367
R1890 B.n735 B.n734 163.367
R1891 B.n734 B.n49 163.367
R1892 B.n730 B.n49 163.367
R1893 B.n730 B.n729 163.367
R1894 B.n729 B.n728 163.367
R1895 B.n728 B.n51 163.367
R1896 B.n724 B.n51 163.367
R1897 B.n724 B.n723 163.367
R1898 B.n723 B.n722 163.367
R1899 B.n722 B.n53 163.367
R1900 B.n717 B.n53 163.367
R1901 B.n717 B.n716 163.367
R1902 B.n716 B.n715 163.367
R1903 B.n715 B.n57 163.367
R1904 B.n711 B.n57 163.367
R1905 B.n711 B.n710 163.367
R1906 B.n710 B.n709 163.367
R1907 B.n709 B.n59 163.367
R1908 B.n705 B.n59 163.367
R1909 B.n705 B.n704 163.367
R1910 B.n704 B.n63 163.367
R1911 B.n700 B.n63 163.367
R1912 B.n700 B.n699 163.367
R1913 B.n699 B.n698 163.367
R1914 B.n698 B.n65 163.367
R1915 B.n694 B.n65 163.367
R1916 B.n694 B.n693 163.367
R1917 B.n693 B.n692 163.367
R1918 B.n692 B.n67 163.367
R1919 B.n688 B.n67 163.367
R1920 B.n688 B.n687 163.367
R1921 B.n687 B.n686 163.367
R1922 B.n686 B.n69 163.367
R1923 B.n682 B.n69 163.367
R1924 B.n682 B.n681 163.367
R1925 B.n681 B.n680 163.367
R1926 B.n680 B.n71 163.367
R1927 B.n676 B.n71 163.367
R1928 B.n676 B.n675 163.367
R1929 B.n675 B.n674 163.367
R1930 B.n674 B.n73 163.367
R1931 B.n670 B.n73 163.367
R1932 B.n670 B.n669 163.367
R1933 B.n669 B.n668 163.367
R1934 B.n668 B.n75 163.367
R1935 B.n664 B.n75 163.367
R1936 B.n664 B.n663 163.367
R1937 B.n663 B.n662 163.367
R1938 B.n662 B.n77 163.367
R1939 B.n658 B.n77 163.367
R1940 B.n658 B.n657 163.367
R1941 B.n657 B.n656 163.367
R1942 B.n656 B.n79 163.367
R1943 B.n652 B.n79 163.367
R1944 B.n652 B.n651 163.367
R1945 B.n651 B.n650 163.367
R1946 B.n650 B.n81 163.367
R1947 B.n646 B.n81 163.367
R1948 B.n646 B.n645 163.367
R1949 B.n645 B.n644 163.367
R1950 B.n644 B.n83 163.367
R1951 B.n167 B.n166 69.8187
R1952 B.n175 B.n174 69.8187
R1953 B.n55 B.n54 69.8187
R1954 B.n61 B.n60 69.8187
R1955 B.n168 B.n167 59.5399
R1956 B.n379 B.n175 59.5399
R1957 B.n719 B.n55 59.5399
R1958 B.n62 B.n61 59.5399
R1959 B.n781 B.n32 31.6883
R1960 B.n642 B.n641 31.6883
R1961 B.n457 B.n456 31.6883
R1962 B.n317 B.n196 31.6883
R1963 B B.n875 18.0485
R1964 B.n781 B.n780 10.6151
R1965 B.n780 B.n779 10.6151
R1966 B.n779 B.n34 10.6151
R1967 B.n775 B.n34 10.6151
R1968 B.n775 B.n774 10.6151
R1969 B.n774 B.n773 10.6151
R1970 B.n773 B.n36 10.6151
R1971 B.n769 B.n36 10.6151
R1972 B.n769 B.n768 10.6151
R1973 B.n768 B.n767 10.6151
R1974 B.n767 B.n38 10.6151
R1975 B.n763 B.n38 10.6151
R1976 B.n763 B.n762 10.6151
R1977 B.n762 B.n761 10.6151
R1978 B.n761 B.n40 10.6151
R1979 B.n757 B.n40 10.6151
R1980 B.n757 B.n756 10.6151
R1981 B.n756 B.n755 10.6151
R1982 B.n755 B.n42 10.6151
R1983 B.n751 B.n42 10.6151
R1984 B.n751 B.n750 10.6151
R1985 B.n750 B.n749 10.6151
R1986 B.n749 B.n44 10.6151
R1987 B.n745 B.n44 10.6151
R1988 B.n745 B.n744 10.6151
R1989 B.n744 B.n743 10.6151
R1990 B.n743 B.n46 10.6151
R1991 B.n739 B.n46 10.6151
R1992 B.n739 B.n738 10.6151
R1993 B.n738 B.n737 10.6151
R1994 B.n737 B.n48 10.6151
R1995 B.n733 B.n48 10.6151
R1996 B.n733 B.n732 10.6151
R1997 B.n732 B.n731 10.6151
R1998 B.n731 B.n50 10.6151
R1999 B.n727 B.n50 10.6151
R2000 B.n727 B.n726 10.6151
R2001 B.n726 B.n725 10.6151
R2002 B.n725 B.n52 10.6151
R2003 B.n721 B.n52 10.6151
R2004 B.n721 B.n720 10.6151
R2005 B.n718 B.n56 10.6151
R2006 B.n714 B.n56 10.6151
R2007 B.n714 B.n713 10.6151
R2008 B.n713 B.n712 10.6151
R2009 B.n712 B.n58 10.6151
R2010 B.n708 B.n58 10.6151
R2011 B.n708 B.n707 10.6151
R2012 B.n707 B.n706 10.6151
R2013 B.n703 B.n702 10.6151
R2014 B.n702 B.n701 10.6151
R2015 B.n701 B.n64 10.6151
R2016 B.n697 B.n64 10.6151
R2017 B.n697 B.n696 10.6151
R2018 B.n696 B.n695 10.6151
R2019 B.n695 B.n66 10.6151
R2020 B.n691 B.n66 10.6151
R2021 B.n691 B.n690 10.6151
R2022 B.n690 B.n689 10.6151
R2023 B.n689 B.n68 10.6151
R2024 B.n685 B.n68 10.6151
R2025 B.n685 B.n684 10.6151
R2026 B.n684 B.n683 10.6151
R2027 B.n683 B.n70 10.6151
R2028 B.n679 B.n70 10.6151
R2029 B.n679 B.n678 10.6151
R2030 B.n678 B.n677 10.6151
R2031 B.n677 B.n72 10.6151
R2032 B.n673 B.n72 10.6151
R2033 B.n673 B.n672 10.6151
R2034 B.n672 B.n671 10.6151
R2035 B.n671 B.n74 10.6151
R2036 B.n667 B.n74 10.6151
R2037 B.n667 B.n666 10.6151
R2038 B.n666 B.n665 10.6151
R2039 B.n665 B.n76 10.6151
R2040 B.n661 B.n76 10.6151
R2041 B.n661 B.n660 10.6151
R2042 B.n660 B.n659 10.6151
R2043 B.n659 B.n78 10.6151
R2044 B.n655 B.n78 10.6151
R2045 B.n655 B.n654 10.6151
R2046 B.n654 B.n653 10.6151
R2047 B.n653 B.n80 10.6151
R2048 B.n649 B.n80 10.6151
R2049 B.n649 B.n648 10.6151
R2050 B.n648 B.n647 10.6151
R2051 B.n647 B.n82 10.6151
R2052 B.n643 B.n82 10.6151
R2053 B.n643 B.n642 10.6151
R2054 B.n457 B.n144 10.6151
R2055 B.n461 B.n144 10.6151
R2056 B.n462 B.n461 10.6151
R2057 B.n463 B.n462 10.6151
R2058 B.n463 B.n142 10.6151
R2059 B.n467 B.n142 10.6151
R2060 B.n468 B.n467 10.6151
R2061 B.n469 B.n468 10.6151
R2062 B.n469 B.n140 10.6151
R2063 B.n473 B.n140 10.6151
R2064 B.n474 B.n473 10.6151
R2065 B.n475 B.n474 10.6151
R2066 B.n475 B.n138 10.6151
R2067 B.n479 B.n138 10.6151
R2068 B.n480 B.n479 10.6151
R2069 B.n481 B.n480 10.6151
R2070 B.n481 B.n136 10.6151
R2071 B.n485 B.n136 10.6151
R2072 B.n486 B.n485 10.6151
R2073 B.n487 B.n486 10.6151
R2074 B.n487 B.n134 10.6151
R2075 B.n491 B.n134 10.6151
R2076 B.n492 B.n491 10.6151
R2077 B.n493 B.n492 10.6151
R2078 B.n493 B.n132 10.6151
R2079 B.n497 B.n132 10.6151
R2080 B.n498 B.n497 10.6151
R2081 B.n499 B.n498 10.6151
R2082 B.n499 B.n130 10.6151
R2083 B.n503 B.n130 10.6151
R2084 B.n504 B.n503 10.6151
R2085 B.n505 B.n504 10.6151
R2086 B.n505 B.n128 10.6151
R2087 B.n509 B.n128 10.6151
R2088 B.n510 B.n509 10.6151
R2089 B.n511 B.n510 10.6151
R2090 B.n511 B.n126 10.6151
R2091 B.n515 B.n126 10.6151
R2092 B.n516 B.n515 10.6151
R2093 B.n517 B.n516 10.6151
R2094 B.n517 B.n124 10.6151
R2095 B.n521 B.n124 10.6151
R2096 B.n522 B.n521 10.6151
R2097 B.n523 B.n522 10.6151
R2098 B.n523 B.n122 10.6151
R2099 B.n527 B.n122 10.6151
R2100 B.n528 B.n527 10.6151
R2101 B.n529 B.n528 10.6151
R2102 B.n529 B.n120 10.6151
R2103 B.n533 B.n120 10.6151
R2104 B.n534 B.n533 10.6151
R2105 B.n535 B.n534 10.6151
R2106 B.n535 B.n118 10.6151
R2107 B.n539 B.n118 10.6151
R2108 B.n540 B.n539 10.6151
R2109 B.n541 B.n540 10.6151
R2110 B.n541 B.n116 10.6151
R2111 B.n545 B.n116 10.6151
R2112 B.n546 B.n545 10.6151
R2113 B.n547 B.n546 10.6151
R2114 B.n547 B.n114 10.6151
R2115 B.n551 B.n114 10.6151
R2116 B.n552 B.n551 10.6151
R2117 B.n553 B.n552 10.6151
R2118 B.n553 B.n112 10.6151
R2119 B.n557 B.n112 10.6151
R2120 B.n558 B.n557 10.6151
R2121 B.n559 B.n558 10.6151
R2122 B.n559 B.n110 10.6151
R2123 B.n563 B.n110 10.6151
R2124 B.n564 B.n563 10.6151
R2125 B.n565 B.n564 10.6151
R2126 B.n565 B.n108 10.6151
R2127 B.n569 B.n108 10.6151
R2128 B.n570 B.n569 10.6151
R2129 B.n571 B.n570 10.6151
R2130 B.n571 B.n106 10.6151
R2131 B.n575 B.n106 10.6151
R2132 B.n576 B.n575 10.6151
R2133 B.n577 B.n576 10.6151
R2134 B.n577 B.n104 10.6151
R2135 B.n581 B.n104 10.6151
R2136 B.n582 B.n581 10.6151
R2137 B.n583 B.n582 10.6151
R2138 B.n583 B.n102 10.6151
R2139 B.n587 B.n102 10.6151
R2140 B.n588 B.n587 10.6151
R2141 B.n589 B.n588 10.6151
R2142 B.n589 B.n100 10.6151
R2143 B.n593 B.n100 10.6151
R2144 B.n594 B.n593 10.6151
R2145 B.n595 B.n594 10.6151
R2146 B.n595 B.n98 10.6151
R2147 B.n599 B.n98 10.6151
R2148 B.n600 B.n599 10.6151
R2149 B.n601 B.n600 10.6151
R2150 B.n601 B.n96 10.6151
R2151 B.n605 B.n96 10.6151
R2152 B.n606 B.n605 10.6151
R2153 B.n607 B.n606 10.6151
R2154 B.n607 B.n94 10.6151
R2155 B.n611 B.n94 10.6151
R2156 B.n612 B.n611 10.6151
R2157 B.n613 B.n612 10.6151
R2158 B.n613 B.n92 10.6151
R2159 B.n617 B.n92 10.6151
R2160 B.n618 B.n617 10.6151
R2161 B.n619 B.n618 10.6151
R2162 B.n619 B.n90 10.6151
R2163 B.n623 B.n90 10.6151
R2164 B.n624 B.n623 10.6151
R2165 B.n625 B.n624 10.6151
R2166 B.n625 B.n88 10.6151
R2167 B.n629 B.n88 10.6151
R2168 B.n630 B.n629 10.6151
R2169 B.n631 B.n630 10.6151
R2170 B.n631 B.n86 10.6151
R2171 B.n635 B.n86 10.6151
R2172 B.n636 B.n635 10.6151
R2173 B.n637 B.n636 10.6151
R2174 B.n637 B.n84 10.6151
R2175 B.n641 B.n84 10.6151
R2176 B.n318 B.n317 10.6151
R2177 B.n319 B.n318 10.6151
R2178 B.n319 B.n194 10.6151
R2179 B.n323 B.n194 10.6151
R2180 B.n324 B.n323 10.6151
R2181 B.n325 B.n324 10.6151
R2182 B.n325 B.n192 10.6151
R2183 B.n329 B.n192 10.6151
R2184 B.n330 B.n329 10.6151
R2185 B.n331 B.n330 10.6151
R2186 B.n331 B.n190 10.6151
R2187 B.n335 B.n190 10.6151
R2188 B.n336 B.n335 10.6151
R2189 B.n337 B.n336 10.6151
R2190 B.n337 B.n188 10.6151
R2191 B.n341 B.n188 10.6151
R2192 B.n342 B.n341 10.6151
R2193 B.n343 B.n342 10.6151
R2194 B.n343 B.n186 10.6151
R2195 B.n347 B.n186 10.6151
R2196 B.n348 B.n347 10.6151
R2197 B.n349 B.n348 10.6151
R2198 B.n349 B.n184 10.6151
R2199 B.n353 B.n184 10.6151
R2200 B.n354 B.n353 10.6151
R2201 B.n355 B.n354 10.6151
R2202 B.n355 B.n182 10.6151
R2203 B.n359 B.n182 10.6151
R2204 B.n360 B.n359 10.6151
R2205 B.n361 B.n360 10.6151
R2206 B.n361 B.n180 10.6151
R2207 B.n365 B.n180 10.6151
R2208 B.n366 B.n365 10.6151
R2209 B.n367 B.n366 10.6151
R2210 B.n367 B.n178 10.6151
R2211 B.n371 B.n178 10.6151
R2212 B.n372 B.n371 10.6151
R2213 B.n373 B.n372 10.6151
R2214 B.n373 B.n176 10.6151
R2215 B.n377 B.n176 10.6151
R2216 B.n378 B.n377 10.6151
R2217 B.n380 B.n172 10.6151
R2218 B.n384 B.n172 10.6151
R2219 B.n385 B.n384 10.6151
R2220 B.n386 B.n385 10.6151
R2221 B.n386 B.n170 10.6151
R2222 B.n390 B.n170 10.6151
R2223 B.n391 B.n390 10.6151
R2224 B.n392 B.n391 10.6151
R2225 B.n396 B.n395 10.6151
R2226 B.n397 B.n396 10.6151
R2227 B.n397 B.n164 10.6151
R2228 B.n401 B.n164 10.6151
R2229 B.n402 B.n401 10.6151
R2230 B.n403 B.n402 10.6151
R2231 B.n403 B.n162 10.6151
R2232 B.n407 B.n162 10.6151
R2233 B.n408 B.n407 10.6151
R2234 B.n409 B.n408 10.6151
R2235 B.n409 B.n160 10.6151
R2236 B.n413 B.n160 10.6151
R2237 B.n414 B.n413 10.6151
R2238 B.n415 B.n414 10.6151
R2239 B.n415 B.n158 10.6151
R2240 B.n419 B.n158 10.6151
R2241 B.n420 B.n419 10.6151
R2242 B.n421 B.n420 10.6151
R2243 B.n421 B.n156 10.6151
R2244 B.n425 B.n156 10.6151
R2245 B.n426 B.n425 10.6151
R2246 B.n427 B.n426 10.6151
R2247 B.n427 B.n154 10.6151
R2248 B.n431 B.n154 10.6151
R2249 B.n432 B.n431 10.6151
R2250 B.n433 B.n432 10.6151
R2251 B.n433 B.n152 10.6151
R2252 B.n437 B.n152 10.6151
R2253 B.n438 B.n437 10.6151
R2254 B.n439 B.n438 10.6151
R2255 B.n439 B.n150 10.6151
R2256 B.n443 B.n150 10.6151
R2257 B.n444 B.n443 10.6151
R2258 B.n445 B.n444 10.6151
R2259 B.n445 B.n148 10.6151
R2260 B.n449 B.n148 10.6151
R2261 B.n450 B.n449 10.6151
R2262 B.n451 B.n450 10.6151
R2263 B.n451 B.n146 10.6151
R2264 B.n455 B.n146 10.6151
R2265 B.n456 B.n455 10.6151
R2266 B.n313 B.n196 10.6151
R2267 B.n313 B.n312 10.6151
R2268 B.n312 B.n311 10.6151
R2269 B.n311 B.n198 10.6151
R2270 B.n307 B.n198 10.6151
R2271 B.n307 B.n306 10.6151
R2272 B.n306 B.n305 10.6151
R2273 B.n305 B.n200 10.6151
R2274 B.n301 B.n200 10.6151
R2275 B.n301 B.n300 10.6151
R2276 B.n300 B.n299 10.6151
R2277 B.n299 B.n202 10.6151
R2278 B.n295 B.n202 10.6151
R2279 B.n295 B.n294 10.6151
R2280 B.n294 B.n293 10.6151
R2281 B.n293 B.n204 10.6151
R2282 B.n289 B.n204 10.6151
R2283 B.n289 B.n288 10.6151
R2284 B.n288 B.n287 10.6151
R2285 B.n287 B.n206 10.6151
R2286 B.n283 B.n206 10.6151
R2287 B.n283 B.n282 10.6151
R2288 B.n282 B.n281 10.6151
R2289 B.n281 B.n208 10.6151
R2290 B.n277 B.n208 10.6151
R2291 B.n277 B.n276 10.6151
R2292 B.n276 B.n275 10.6151
R2293 B.n275 B.n210 10.6151
R2294 B.n271 B.n210 10.6151
R2295 B.n271 B.n270 10.6151
R2296 B.n270 B.n269 10.6151
R2297 B.n269 B.n212 10.6151
R2298 B.n265 B.n212 10.6151
R2299 B.n265 B.n264 10.6151
R2300 B.n264 B.n263 10.6151
R2301 B.n263 B.n214 10.6151
R2302 B.n259 B.n214 10.6151
R2303 B.n259 B.n258 10.6151
R2304 B.n258 B.n257 10.6151
R2305 B.n257 B.n216 10.6151
R2306 B.n253 B.n216 10.6151
R2307 B.n253 B.n252 10.6151
R2308 B.n252 B.n251 10.6151
R2309 B.n251 B.n218 10.6151
R2310 B.n247 B.n218 10.6151
R2311 B.n247 B.n246 10.6151
R2312 B.n246 B.n245 10.6151
R2313 B.n245 B.n220 10.6151
R2314 B.n241 B.n220 10.6151
R2315 B.n241 B.n240 10.6151
R2316 B.n240 B.n239 10.6151
R2317 B.n239 B.n222 10.6151
R2318 B.n235 B.n222 10.6151
R2319 B.n235 B.n234 10.6151
R2320 B.n234 B.n233 10.6151
R2321 B.n233 B.n224 10.6151
R2322 B.n229 B.n224 10.6151
R2323 B.n229 B.n228 10.6151
R2324 B.n228 B.n227 10.6151
R2325 B.n227 B.n0 10.6151
R2326 B.n871 B.n1 10.6151
R2327 B.n871 B.n870 10.6151
R2328 B.n870 B.n869 10.6151
R2329 B.n869 B.n4 10.6151
R2330 B.n865 B.n4 10.6151
R2331 B.n865 B.n864 10.6151
R2332 B.n864 B.n863 10.6151
R2333 B.n863 B.n6 10.6151
R2334 B.n859 B.n6 10.6151
R2335 B.n859 B.n858 10.6151
R2336 B.n858 B.n857 10.6151
R2337 B.n857 B.n8 10.6151
R2338 B.n853 B.n8 10.6151
R2339 B.n853 B.n852 10.6151
R2340 B.n852 B.n851 10.6151
R2341 B.n851 B.n10 10.6151
R2342 B.n847 B.n10 10.6151
R2343 B.n847 B.n846 10.6151
R2344 B.n846 B.n845 10.6151
R2345 B.n845 B.n12 10.6151
R2346 B.n841 B.n12 10.6151
R2347 B.n841 B.n840 10.6151
R2348 B.n840 B.n839 10.6151
R2349 B.n839 B.n14 10.6151
R2350 B.n835 B.n14 10.6151
R2351 B.n835 B.n834 10.6151
R2352 B.n834 B.n833 10.6151
R2353 B.n833 B.n16 10.6151
R2354 B.n829 B.n16 10.6151
R2355 B.n829 B.n828 10.6151
R2356 B.n828 B.n827 10.6151
R2357 B.n827 B.n18 10.6151
R2358 B.n823 B.n18 10.6151
R2359 B.n823 B.n822 10.6151
R2360 B.n822 B.n821 10.6151
R2361 B.n821 B.n20 10.6151
R2362 B.n817 B.n20 10.6151
R2363 B.n817 B.n816 10.6151
R2364 B.n816 B.n815 10.6151
R2365 B.n815 B.n22 10.6151
R2366 B.n811 B.n22 10.6151
R2367 B.n811 B.n810 10.6151
R2368 B.n810 B.n809 10.6151
R2369 B.n809 B.n24 10.6151
R2370 B.n805 B.n24 10.6151
R2371 B.n805 B.n804 10.6151
R2372 B.n804 B.n803 10.6151
R2373 B.n803 B.n26 10.6151
R2374 B.n799 B.n26 10.6151
R2375 B.n799 B.n798 10.6151
R2376 B.n798 B.n797 10.6151
R2377 B.n797 B.n28 10.6151
R2378 B.n793 B.n28 10.6151
R2379 B.n793 B.n792 10.6151
R2380 B.n792 B.n791 10.6151
R2381 B.n791 B.n30 10.6151
R2382 B.n787 B.n30 10.6151
R2383 B.n787 B.n786 10.6151
R2384 B.n786 B.n785 10.6151
R2385 B.n785 B.n32 10.6151
R2386 B.n719 B.n718 6.5566
R2387 B.n706 B.n62 6.5566
R2388 B.n380 B.n379 6.5566
R2389 B.n392 B.n168 6.5566
R2390 B.n720 B.n719 4.05904
R2391 B.n703 B.n62 4.05904
R2392 B.n379 B.n378 4.05904
R2393 B.n395 B.n168 4.05904
R2394 B.n875 B.n0 2.81026
R2395 B.n875 B.n1 2.81026
C0 VP VTAIL 9.686069f
C1 B w_n4570_n3366# 11.138201f
C2 B VN 1.38108f
C3 w_n4570_n3366# VDD2 2.31174f
C4 VP VDD1 9.483871f
C5 VN VDD2 9.04758f
C6 B VP 2.38251f
C7 VP VDD2 0.590847f
C8 VTAIL VDD1 8.30755f
C9 B VTAIL 5.26606f
C10 VTAIL VDD2 8.366461f
C11 B VDD1 1.8533f
C12 VDD1 VDD2 2.12564f
C13 B VDD2 1.9704f
C14 w_n4570_n3366# VN 9.48423f
C15 VP w_n4570_n3366# 10.0795f
C16 VP VN 8.478379f
C17 w_n4570_n3366# VTAIL 4.2603f
C18 VN VTAIL 9.671969f
C19 w_n4570_n3366# VDD1 2.16893f
C20 VN VDD1 0.152821f
C21 VDD2 VSUBS 2.183754f
C22 VDD1 VSUBS 2.95358f
C23 VTAIL VSUBS 1.457169f
C24 VN VSUBS 7.6412f
C25 VP VSUBS 4.282788f
C26 B VSUBS 5.749957f
C27 w_n4570_n3366# VSUBS 0.189363p
C28 B.n0 VSUBS 0.004635f
C29 B.n1 VSUBS 0.004635f
C30 B.n2 VSUBS 0.007329f
C31 B.n3 VSUBS 0.007329f
C32 B.n4 VSUBS 0.007329f
C33 B.n5 VSUBS 0.007329f
C34 B.n6 VSUBS 0.007329f
C35 B.n7 VSUBS 0.007329f
C36 B.n8 VSUBS 0.007329f
C37 B.n9 VSUBS 0.007329f
C38 B.n10 VSUBS 0.007329f
C39 B.n11 VSUBS 0.007329f
C40 B.n12 VSUBS 0.007329f
C41 B.n13 VSUBS 0.007329f
C42 B.n14 VSUBS 0.007329f
C43 B.n15 VSUBS 0.007329f
C44 B.n16 VSUBS 0.007329f
C45 B.n17 VSUBS 0.007329f
C46 B.n18 VSUBS 0.007329f
C47 B.n19 VSUBS 0.007329f
C48 B.n20 VSUBS 0.007329f
C49 B.n21 VSUBS 0.007329f
C50 B.n22 VSUBS 0.007329f
C51 B.n23 VSUBS 0.007329f
C52 B.n24 VSUBS 0.007329f
C53 B.n25 VSUBS 0.007329f
C54 B.n26 VSUBS 0.007329f
C55 B.n27 VSUBS 0.007329f
C56 B.n28 VSUBS 0.007329f
C57 B.n29 VSUBS 0.007329f
C58 B.n30 VSUBS 0.007329f
C59 B.n31 VSUBS 0.007329f
C60 B.n32 VSUBS 0.01626f
C61 B.n33 VSUBS 0.007329f
C62 B.n34 VSUBS 0.007329f
C63 B.n35 VSUBS 0.007329f
C64 B.n36 VSUBS 0.007329f
C65 B.n37 VSUBS 0.007329f
C66 B.n38 VSUBS 0.007329f
C67 B.n39 VSUBS 0.007329f
C68 B.n40 VSUBS 0.007329f
C69 B.n41 VSUBS 0.007329f
C70 B.n42 VSUBS 0.007329f
C71 B.n43 VSUBS 0.007329f
C72 B.n44 VSUBS 0.007329f
C73 B.n45 VSUBS 0.007329f
C74 B.n46 VSUBS 0.007329f
C75 B.n47 VSUBS 0.007329f
C76 B.n48 VSUBS 0.007329f
C77 B.n49 VSUBS 0.007329f
C78 B.n50 VSUBS 0.007329f
C79 B.n51 VSUBS 0.007329f
C80 B.n52 VSUBS 0.007329f
C81 B.n53 VSUBS 0.007329f
C82 B.t5 VSUBS 0.220581f
C83 B.t4 VSUBS 0.260753f
C84 B.t3 VSUBS 1.89781f
C85 B.n54 VSUBS 0.416564f
C86 B.n55 VSUBS 0.266588f
C87 B.n56 VSUBS 0.007329f
C88 B.n57 VSUBS 0.007329f
C89 B.n58 VSUBS 0.007329f
C90 B.n59 VSUBS 0.007329f
C91 B.t2 VSUBS 0.220584f
C92 B.t1 VSUBS 0.260756f
C93 B.t0 VSUBS 1.89781f
C94 B.n60 VSUBS 0.416561f
C95 B.n61 VSUBS 0.266585f
C96 B.n62 VSUBS 0.016981f
C97 B.n63 VSUBS 0.007329f
C98 B.n64 VSUBS 0.007329f
C99 B.n65 VSUBS 0.007329f
C100 B.n66 VSUBS 0.007329f
C101 B.n67 VSUBS 0.007329f
C102 B.n68 VSUBS 0.007329f
C103 B.n69 VSUBS 0.007329f
C104 B.n70 VSUBS 0.007329f
C105 B.n71 VSUBS 0.007329f
C106 B.n72 VSUBS 0.007329f
C107 B.n73 VSUBS 0.007329f
C108 B.n74 VSUBS 0.007329f
C109 B.n75 VSUBS 0.007329f
C110 B.n76 VSUBS 0.007329f
C111 B.n77 VSUBS 0.007329f
C112 B.n78 VSUBS 0.007329f
C113 B.n79 VSUBS 0.007329f
C114 B.n80 VSUBS 0.007329f
C115 B.n81 VSUBS 0.007329f
C116 B.n82 VSUBS 0.007329f
C117 B.n83 VSUBS 0.01737f
C118 B.n84 VSUBS 0.007329f
C119 B.n85 VSUBS 0.007329f
C120 B.n86 VSUBS 0.007329f
C121 B.n87 VSUBS 0.007329f
C122 B.n88 VSUBS 0.007329f
C123 B.n89 VSUBS 0.007329f
C124 B.n90 VSUBS 0.007329f
C125 B.n91 VSUBS 0.007329f
C126 B.n92 VSUBS 0.007329f
C127 B.n93 VSUBS 0.007329f
C128 B.n94 VSUBS 0.007329f
C129 B.n95 VSUBS 0.007329f
C130 B.n96 VSUBS 0.007329f
C131 B.n97 VSUBS 0.007329f
C132 B.n98 VSUBS 0.007329f
C133 B.n99 VSUBS 0.007329f
C134 B.n100 VSUBS 0.007329f
C135 B.n101 VSUBS 0.007329f
C136 B.n102 VSUBS 0.007329f
C137 B.n103 VSUBS 0.007329f
C138 B.n104 VSUBS 0.007329f
C139 B.n105 VSUBS 0.007329f
C140 B.n106 VSUBS 0.007329f
C141 B.n107 VSUBS 0.007329f
C142 B.n108 VSUBS 0.007329f
C143 B.n109 VSUBS 0.007329f
C144 B.n110 VSUBS 0.007329f
C145 B.n111 VSUBS 0.007329f
C146 B.n112 VSUBS 0.007329f
C147 B.n113 VSUBS 0.007329f
C148 B.n114 VSUBS 0.007329f
C149 B.n115 VSUBS 0.007329f
C150 B.n116 VSUBS 0.007329f
C151 B.n117 VSUBS 0.007329f
C152 B.n118 VSUBS 0.007329f
C153 B.n119 VSUBS 0.007329f
C154 B.n120 VSUBS 0.007329f
C155 B.n121 VSUBS 0.007329f
C156 B.n122 VSUBS 0.007329f
C157 B.n123 VSUBS 0.007329f
C158 B.n124 VSUBS 0.007329f
C159 B.n125 VSUBS 0.007329f
C160 B.n126 VSUBS 0.007329f
C161 B.n127 VSUBS 0.007329f
C162 B.n128 VSUBS 0.007329f
C163 B.n129 VSUBS 0.007329f
C164 B.n130 VSUBS 0.007329f
C165 B.n131 VSUBS 0.007329f
C166 B.n132 VSUBS 0.007329f
C167 B.n133 VSUBS 0.007329f
C168 B.n134 VSUBS 0.007329f
C169 B.n135 VSUBS 0.007329f
C170 B.n136 VSUBS 0.007329f
C171 B.n137 VSUBS 0.007329f
C172 B.n138 VSUBS 0.007329f
C173 B.n139 VSUBS 0.007329f
C174 B.n140 VSUBS 0.007329f
C175 B.n141 VSUBS 0.007329f
C176 B.n142 VSUBS 0.007329f
C177 B.n143 VSUBS 0.007329f
C178 B.n144 VSUBS 0.007329f
C179 B.n145 VSUBS 0.01737f
C180 B.n146 VSUBS 0.007329f
C181 B.n147 VSUBS 0.007329f
C182 B.n148 VSUBS 0.007329f
C183 B.n149 VSUBS 0.007329f
C184 B.n150 VSUBS 0.007329f
C185 B.n151 VSUBS 0.007329f
C186 B.n152 VSUBS 0.007329f
C187 B.n153 VSUBS 0.007329f
C188 B.n154 VSUBS 0.007329f
C189 B.n155 VSUBS 0.007329f
C190 B.n156 VSUBS 0.007329f
C191 B.n157 VSUBS 0.007329f
C192 B.n158 VSUBS 0.007329f
C193 B.n159 VSUBS 0.007329f
C194 B.n160 VSUBS 0.007329f
C195 B.n161 VSUBS 0.007329f
C196 B.n162 VSUBS 0.007329f
C197 B.n163 VSUBS 0.007329f
C198 B.n164 VSUBS 0.007329f
C199 B.n165 VSUBS 0.007329f
C200 B.t10 VSUBS 0.220584f
C201 B.t11 VSUBS 0.260756f
C202 B.t9 VSUBS 1.89781f
C203 B.n166 VSUBS 0.416561f
C204 B.n167 VSUBS 0.266585f
C205 B.n168 VSUBS 0.016981f
C206 B.n169 VSUBS 0.007329f
C207 B.n170 VSUBS 0.007329f
C208 B.n171 VSUBS 0.007329f
C209 B.n172 VSUBS 0.007329f
C210 B.n173 VSUBS 0.007329f
C211 B.t7 VSUBS 0.220581f
C212 B.t8 VSUBS 0.260753f
C213 B.t6 VSUBS 1.89781f
C214 B.n174 VSUBS 0.416564f
C215 B.n175 VSUBS 0.266588f
C216 B.n176 VSUBS 0.007329f
C217 B.n177 VSUBS 0.007329f
C218 B.n178 VSUBS 0.007329f
C219 B.n179 VSUBS 0.007329f
C220 B.n180 VSUBS 0.007329f
C221 B.n181 VSUBS 0.007329f
C222 B.n182 VSUBS 0.007329f
C223 B.n183 VSUBS 0.007329f
C224 B.n184 VSUBS 0.007329f
C225 B.n185 VSUBS 0.007329f
C226 B.n186 VSUBS 0.007329f
C227 B.n187 VSUBS 0.007329f
C228 B.n188 VSUBS 0.007329f
C229 B.n189 VSUBS 0.007329f
C230 B.n190 VSUBS 0.007329f
C231 B.n191 VSUBS 0.007329f
C232 B.n192 VSUBS 0.007329f
C233 B.n193 VSUBS 0.007329f
C234 B.n194 VSUBS 0.007329f
C235 B.n195 VSUBS 0.007329f
C236 B.n196 VSUBS 0.01626f
C237 B.n197 VSUBS 0.007329f
C238 B.n198 VSUBS 0.007329f
C239 B.n199 VSUBS 0.007329f
C240 B.n200 VSUBS 0.007329f
C241 B.n201 VSUBS 0.007329f
C242 B.n202 VSUBS 0.007329f
C243 B.n203 VSUBS 0.007329f
C244 B.n204 VSUBS 0.007329f
C245 B.n205 VSUBS 0.007329f
C246 B.n206 VSUBS 0.007329f
C247 B.n207 VSUBS 0.007329f
C248 B.n208 VSUBS 0.007329f
C249 B.n209 VSUBS 0.007329f
C250 B.n210 VSUBS 0.007329f
C251 B.n211 VSUBS 0.007329f
C252 B.n212 VSUBS 0.007329f
C253 B.n213 VSUBS 0.007329f
C254 B.n214 VSUBS 0.007329f
C255 B.n215 VSUBS 0.007329f
C256 B.n216 VSUBS 0.007329f
C257 B.n217 VSUBS 0.007329f
C258 B.n218 VSUBS 0.007329f
C259 B.n219 VSUBS 0.007329f
C260 B.n220 VSUBS 0.007329f
C261 B.n221 VSUBS 0.007329f
C262 B.n222 VSUBS 0.007329f
C263 B.n223 VSUBS 0.007329f
C264 B.n224 VSUBS 0.007329f
C265 B.n225 VSUBS 0.007329f
C266 B.n226 VSUBS 0.007329f
C267 B.n227 VSUBS 0.007329f
C268 B.n228 VSUBS 0.007329f
C269 B.n229 VSUBS 0.007329f
C270 B.n230 VSUBS 0.007329f
C271 B.n231 VSUBS 0.007329f
C272 B.n232 VSUBS 0.007329f
C273 B.n233 VSUBS 0.007329f
C274 B.n234 VSUBS 0.007329f
C275 B.n235 VSUBS 0.007329f
C276 B.n236 VSUBS 0.007329f
C277 B.n237 VSUBS 0.007329f
C278 B.n238 VSUBS 0.007329f
C279 B.n239 VSUBS 0.007329f
C280 B.n240 VSUBS 0.007329f
C281 B.n241 VSUBS 0.007329f
C282 B.n242 VSUBS 0.007329f
C283 B.n243 VSUBS 0.007329f
C284 B.n244 VSUBS 0.007329f
C285 B.n245 VSUBS 0.007329f
C286 B.n246 VSUBS 0.007329f
C287 B.n247 VSUBS 0.007329f
C288 B.n248 VSUBS 0.007329f
C289 B.n249 VSUBS 0.007329f
C290 B.n250 VSUBS 0.007329f
C291 B.n251 VSUBS 0.007329f
C292 B.n252 VSUBS 0.007329f
C293 B.n253 VSUBS 0.007329f
C294 B.n254 VSUBS 0.007329f
C295 B.n255 VSUBS 0.007329f
C296 B.n256 VSUBS 0.007329f
C297 B.n257 VSUBS 0.007329f
C298 B.n258 VSUBS 0.007329f
C299 B.n259 VSUBS 0.007329f
C300 B.n260 VSUBS 0.007329f
C301 B.n261 VSUBS 0.007329f
C302 B.n262 VSUBS 0.007329f
C303 B.n263 VSUBS 0.007329f
C304 B.n264 VSUBS 0.007329f
C305 B.n265 VSUBS 0.007329f
C306 B.n266 VSUBS 0.007329f
C307 B.n267 VSUBS 0.007329f
C308 B.n268 VSUBS 0.007329f
C309 B.n269 VSUBS 0.007329f
C310 B.n270 VSUBS 0.007329f
C311 B.n271 VSUBS 0.007329f
C312 B.n272 VSUBS 0.007329f
C313 B.n273 VSUBS 0.007329f
C314 B.n274 VSUBS 0.007329f
C315 B.n275 VSUBS 0.007329f
C316 B.n276 VSUBS 0.007329f
C317 B.n277 VSUBS 0.007329f
C318 B.n278 VSUBS 0.007329f
C319 B.n279 VSUBS 0.007329f
C320 B.n280 VSUBS 0.007329f
C321 B.n281 VSUBS 0.007329f
C322 B.n282 VSUBS 0.007329f
C323 B.n283 VSUBS 0.007329f
C324 B.n284 VSUBS 0.007329f
C325 B.n285 VSUBS 0.007329f
C326 B.n286 VSUBS 0.007329f
C327 B.n287 VSUBS 0.007329f
C328 B.n288 VSUBS 0.007329f
C329 B.n289 VSUBS 0.007329f
C330 B.n290 VSUBS 0.007329f
C331 B.n291 VSUBS 0.007329f
C332 B.n292 VSUBS 0.007329f
C333 B.n293 VSUBS 0.007329f
C334 B.n294 VSUBS 0.007329f
C335 B.n295 VSUBS 0.007329f
C336 B.n296 VSUBS 0.007329f
C337 B.n297 VSUBS 0.007329f
C338 B.n298 VSUBS 0.007329f
C339 B.n299 VSUBS 0.007329f
C340 B.n300 VSUBS 0.007329f
C341 B.n301 VSUBS 0.007329f
C342 B.n302 VSUBS 0.007329f
C343 B.n303 VSUBS 0.007329f
C344 B.n304 VSUBS 0.007329f
C345 B.n305 VSUBS 0.007329f
C346 B.n306 VSUBS 0.007329f
C347 B.n307 VSUBS 0.007329f
C348 B.n308 VSUBS 0.007329f
C349 B.n309 VSUBS 0.007329f
C350 B.n310 VSUBS 0.007329f
C351 B.n311 VSUBS 0.007329f
C352 B.n312 VSUBS 0.007329f
C353 B.n313 VSUBS 0.007329f
C354 B.n314 VSUBS 0.007329f
C355 B.n315 VSUBS 0.01626f
C356 B.n316 VSUBS 0.01737f
C357 B.n317 VSUBS 0.01737f
C358 B.n318 VSUBS 0.007329f
C359 B.n319 VSUBS 0.007329f
C360 B.n320 VSUBS 0.007329f
C361 B.n321 VSUBS 0.007329f
C362 B.n322 VSUBS 0.007329f
C363 B.n323 VSUBS 0.007329f
C364 B.n324 VSUBS 0.007329f
C365 B.n325 VSUBS 0.007329f
C366 B.n326 VSUBS 0.007329f
C367 B.n327 VSUBS 0.007329f
C368 B.n328 VSUBS 0.007329f
C369 B.n329 VSUBS 0.007329f
C370 B.n330 VSUBS 0.007329f
C371 B.n331 VSUBS 0.007329f
C372 B.n332 VSUBS 0.007329f
C373 B.n333 VSUBS 0.007329f
C374 B.n334 VSUBS 0.007329f
C375 B.n335 VSUBS 0.007329f
C376 B.n336 VSUBS 0.007329f
C377 B.n337 VSUBS 0.007329f
C378 B.n338 VSUBS 0.007329f
C379 B.n339 VSUBS 0.007329f
C380 B.n340 VSUBS 0.007329f
C381 B.n341 VSUBS 0.007329f
C382 B.n342 VSUBS 0.007329f
C383 B.n343 VSUBS 0.007329f
C384 B.n344 VSUBS 0.007329f
C385 B.n345 VSUBS 0.007329f
C386 B.n346 VSUBS 0.007329f
C387 B.n347 VSUBS 0.007329f
C388 B.n348 VSUBS 0.007329f
C389 B.n349 VSUBS 0.007329f
C390 B.n350 VSUBS 0.007329f
C391 B.n351 VSUBS 0.007329f
C392 B.n352 VSUBS 0.007329f
C393 B.n353 VSUBS 0.007329f
C394 B.n354 VSUBS 0.007329f
C395 B.n355 VSUBS 0.007329f
C396 B.n356 VSUBS 0.007329f
C397 B.n357 VSUBS 0.007329f
C398 B.n358 VSUBS 0.007329f
C399 B.n359 VSUBS 0.007329f
C400 B.n360 VSUBS 0.007329f
C401 B.n361 VSUBS 0.007329f
C402 B.n362 VSUBS 0.007329f
C403 B.n363 VSUBS 0.007329f
C404 B.n364 VSUBS 0.007329f
C405 B.n365 VSUBS 0.007329f
C406 B.n366 VSUBS 0.007329f
C407 B.n367 VSUBS 0.007329f
C408 B.n368 VSUBS 0.007329f
C409 B.n369 VSUBS 0.007329f
C410 B.n370 VSUBS 0.007329f
C411 B.n371 VSUBS 0.007329f
C412 B.n372 VSUBS 0.007329f
C413 B.n373 VSUBS 0.007329f
C414 B.n374 VSUBS 0.007329f
C415 B.n375 VSUBS 0.007329f
C416 B.n376 VSUBS 0.007329f
C417 B.n377 VSUBS 0.007329f
C418 B.n378 VSUBS 0.005066f
C419 B.n379 VSUBS 0.016981f
C420 B.n380 VSUBS 0.005928f
C421 B.n381 VSUBS 0.007329f
C422 B.n382 VSUBS 0.007329f
C423 B.n383 VSUBS 0.007329f
C424 B.n384 VSUBS 0.007329f
C425 B.n385 VSUBS 0.007329f
C426 B.n386 VSUBS 0.007329f
C427 B.n387 VSUBS 0.007329f
C428 B.n388 VSUBS 0.007329f
C429 B.n389 VSUBS 0.007329f
C430 B.n390 VSUBS 0.007329f
C431 B.n391 VSUBS 0.007329f
C432 B.n392 VSUBS 0.005928f
C433 B.n393 VSUBS 0.007329f
C434 B.n394 VSUBS 0.007329f
C435 B.n395 VSUBS 0.005066f
C436 B.n396 VSUBS 0.007329f
C437 B.n397 VSUBS 0.007329f
C438 B.n398 VSUBS 0.007329f
C439 B.n399 VSUBS 0.007329f
C440 B.n400 VSUBS 0.007329f
C441 B.n401 VSUBS 0.007329f
C442 B.n402 VSUBS 0.007329f
C443 B.n403 VSUBS 0.007329f
C444 B.n404 VSUBS 0.007329f
C445 B.n405 VSUBS 0.007329f
C446 B.n406 VSUBS 0.007329f
C447 B.n407 VSUBS 0.007329f
C448 B.n408 VSUBS 0.007329f
C449 B.n409 VSUBS 0.007329f
C450 B.n410 VSUBS 0.007329f
C451 B.n411 VSUBS 0.007329f
C452 B.n412 VSUBS 0.007329f
C453 B.n413 VSUBS 0.007329f
C454 B.n414 VSUBS 0.007329f
C455 B.n415 VSUBS 0.007329f
C456 B.n416 VSUBS 0.007329f
C457 B.n417 VSUBS 0.007329f
C458 B.n418 VSUBS 0.007329f
C459 B.n419 VSUBS 0.007329f
C460 B.n420 VSUBS 0.007329f
C461 B.n421 VSUBS 0.007329f
C462 B.n422 VSUBS 0.007329f
C463 B.n423 VSUBS 0.007329f
C464 B.n424 VSUBS 0.007329f
C465 B.n425 VSUBS 0.007329f
C466 B.n426 VSUBS 0.007329f
C467 B.n427 VSUBS 0.007329f
C468 B.n428 VSUBS 0.007329f
C469 B.n429 VSUBS 0.007329f
C470 B.n430 VSUBS 0.007329f
C471 B.n431 VSUBS 0.007329f
C472 B.n432 VSUBS 0.007329f
C473 B.n433 VSUBS 0.007329f
C474 B.n434 VSUBS 0.007329f
C475 B.n435 VSUBS 0.007329f
C476 B.n436 VSUBS 0.007329f
C477 B.n437 VSUBS 0.007329f
C478 B.n438 VSUBS 0.007329f
C479 B.n439 VSUBS 0.007329f
C480 B.n440 VSUBS 0.007329f
C481 B.n441 VSUBS 0.007329f
C482 B.n442 VSUBS 0.007329f
C483 B.n443 VSUBS 0.007329f
C484 B.n444 VSUBS 0.007329f
C485 B.n445 VSUBS 0.007329f
C486 B.n446 VSUBS 0.007329f
C487 B.n447 VSUBS 0.007329f
C488 B.n448 VSUBS 0.007329f
C489 B.n449 VSUBS 0.007329f
C490 B.n450 VSUBS 0.007329f
C491 B.n451 VSUBS 0.007329f
C492 B.n452 VSUBS 0.007329f
C493 B.n453 VSUBS 0.007329f
C494 B.n454 VSUBS 0.007329f
C495 B.n455 VSUBS 0.007329f
C496 B.n456 VSUBS 0.01737f
C497 B.n457 VSUBS 0.01626f
C498 B.n458 VSUBS 0.01626f
C499 B.n459 VSUBS 0.007329f
C500 B.n460 VSUBS 0.007329f
C501 B.n461 VSUBS 0.007329f
C502 B.n462 VSUBS 0.007329f
C503 B.n463 VSUBS 0.007329f
C504 B.n464 VSUBS 0.007329f
C505 B.n465 VSUBS 0.007329f
C506 B.n466 VSUBS 0.007329f
C507 B.n467 VSUBS 0.007329f
C508 B.n468 VSUBS 0.007329f
C509 B.n469 VSUBS 0.007329f
C510 B.n470 VSUBS 0.007329f
C511 B.n471 VSUBS 0.007329f
C512 B.n472 VSUBS 0.007329f
C513 B.n473 VSUBS 0.007329f
C514 B.n474 VSUBS 0.007329f
C515 B.n475 VSUBS 0.007329f
C516 B.n476 VSUBS 0.007329f
C517 B.n477 VSUBS 0.007329f
C518 B.n478 VSUBS 0.007329f
C519 B.n479 VSUBS 0.007329f
C520 B.n480 VSUBS 0.007329f
C521 B.n481 VSUBS 0.007329f
C522 B.n482 VSUBS 0.007329f
C523 B.n483 VSUBS 0.007329f
C524 B.n484 VSUBS 0.007329f
C525 B.n485 VSUBS 0.007329f
C526 B.n486 VSUBS 0.007329f
C527 B.n487 VSUBS 0.007329f
C528 B.n488 VSUBS 0.007329f
C529 B.n489 VSUBS 0.007329f
C530 B.n490 VSUBS 0.007329f
C531 B.n491 VSUBS 0.007329f
C532 B.n492 VSUBS 0.007329f
C533 B.n493 VSUBS 0.007329f
C534 B.n494 VSUBS 0.007329f
C535 B.n495 VSUBS 0.007329f
C536 B.n496 VSUBS 0.007329f
C537 B.n497 VSUBS 0.007329f
C538 B.n498 VSUBS 0.007329f
C539 B.n499 VSUBS 0.007329f
C540 B.n500 VSUBS 0.007329f
C541 B.n501 VSUBS 0.007329f
C542 B.n502 VSUBS 0.007329f
C543 B.n503 VSUBS 0.007329f
C544 B.n504 VSUBS 0.007329f
C545 B.n505 VSUBS 0.007329f
C546 B.n506 VSUBS 0.007329f
C547 B.n507 VSUBS 0.007329f
C548 B.n508 VSUBS 0.007329f
C549 B.n509 VSUBS 0.007329f
C550 B.n510 VSUBS 0.007329f
C551 B.n511 VSUBS 0.007329f
C552 B.n512 VSUBS 0.007329f
C553 B.n513 VSUBS 0.007329f
C554 B.n514 VSUBS 0.007329f
C555 B.n515 VSUBS 0.007329f
C556 B.n516 VSUBS 0.007329f
C557 B.n517 VSUBS 0.007329f
C558 B.n518 VSUBS 0.007329f
C559 B.n519 VSUBS 0.007329f
C560 B.n520 VSUBS 0.007329f
C561 B.n521 VSUBS 0.007329f
C562 B.n522 VSUBS 0.007329f
C563 B.n523 VSUBS 0.007329f
C564 B.n524 VSUBS 0.007329f
C565 B.n525 VSUBS 0.007329f
C566 B.n526 VSUBS 0.007329f
C567 B.n527 VSUBS 0.007329f
C568 B.n528 VSUBS 0.007329f
C569 B.n529 VSUBS 0.007329f
C570 B.n530 VSUBS 0.007329f
C571 B.n531 VSUBS 0.007329f
C572 B.n532 VSUBS 0.007329f
C573 B.n533 VSUBS 0.007329f
C574 B.n534 VSUBS 0.007329f
C575 B.n535 VSUBS 0.007329f
C576 B.n536 VSUBS 0.007329f
C577 B.n537 VSUBS 0.007329f
C578 B.n538 VSUBS 0.007329f
C579 B.n539 VSUBS 0.007329f
C580 B.n540 VSUBS 0.007329f
C581 B.n541 VSUBS 0.007329f
C582 B.n542 VSUBS 0.007329f
C583 B.n543 VSUBS 0.007329f
C584 B.n544 VSUBS 0.007329f
C585 B.n545 VSUBS 0.007329f
C586 B.n546 VSUBS 0.007329f
C587 B.n547 VSUBS 0.007329f
C588 B.n548 VSUBS 0.007329f
C589 B.n549 VSUBS 0.007329f
C590 B.n550 VSUBS 0.007329f
C591 B.n551 VSUBS 0.007329f
C592 B.n552 VSUBS 0.007329f
C593 B.n553 VSUBS 0.007329f
C594 B.n554 VSUBS 0.007329f
C595 B.n555 VSUBS 0.007329f
C596 B.n556 VSUBS 0.007329f
C597 B.n557 VSUBS 0.007329f
C598 B.n558 VSUBS 0.007329f
C599 B.n559 VSUBS 0.007329f
C600 B.n560 VSUBS 0.007329f
C601 B.n561 VSUBS 0.007329f
C602 B.n562 VSUBS 0.007329f
C603 B.n563 VSUBS 0.007329f
C604 B.n564 VSUBS 0.007329f
C605 B.n565 VSUBS 0.007329f
C606 B.n566 VSUBS 0.007329f
C607 B.n567 VSUBS 0.007329f
C608 B.n568 VSUBS 0.007329f
C609 B.n569 VSUBS 0.007329f
C610 B.n570 VSUBS 0.007329f
C611 B.n571 VSUBS 0.007329f
C612 B.n572 VSUBS 0.007329f
C613 B.n573 VSUBS 0.007329f
C614 B.n574 VSUBS 0.007329f
C615 B.n575 VSUBS 0.007329f
C616 B.n576 VSUBS 0.007329f
C617 B.n577 VSUBS 0.007329f
C618 B.n578 VSUBS 0.007329f
C619 B.n579 VSUBS 0.007329f
C620 B.n580 VSUBS 0.007329f
C621 B.n581 VSUBS 0.007329f
C622 B.n582 VSUBS 0.007329f
C623 B.n583 VSUBS 0.007329f
C624 B.n584 VSUBS 0.007329f
C625 B.n585 VSUBS 0.007329f
C626 B.n586 VSUBS 0.007329f
C627 B.n587 VSUBS 0.007329f
C628 B.n588 VSUBS 0.007329f
C629 B.n589 VSUBS 0.007329f
C630 B.n590 VSUBS 0.007329f
C631 B.n591 VSUBS 0.007329f
C632 B.n592 VSUBS 0.007329f
C633 B.n593 VSUBS 0.007329f
C634 B.n594 VSUBS 0.007329f
C635 B.n595 VSUBS 0.007329f
C636 B.n596 VSUBS 0.007329f
C637 B.n597 VSUBS 0.007329f
C638 B.n598 VSUBS 0.007329f
C639 B.n599 VSUBS 0.007329f
C640 B.n600 VSUBS 0.007329f
C641 B.n601 VSUBS 0.007329f
C642 B.n602 VSUBS 0.007329f
C643 B.n603 VSUBS 0.007329f
C644 B.n604 VSUBS 0.007329f
C645 B.n605 VSUBS 0.007329f
C646 B.n606 VSUBS 0.007329f
C647 B.n607 VSUBS 0.007329f
C648 B.n608 VSUBS 0.007329f
C649 B.n609 VSUBS 0.007329f
C650 B.n610 VSUBS 0.007329f
C651 B.n611 VSUBS 0.007329f
C652 B.n612 VSUBS 0.007329f
C653 B.n613 VSUBS 0.007329f
C654 B.n614 VSUBS 0.007329f
C655 B.n615 VSUBS 0.007329f
C656 B.n616 VSUBS 0.007329f
C657 B.n617 VSUBS 0.007329f
C658 B.n618 VSUBS 0.007329f
C659 B.n619 VSUBS 0.007329f
C660 B.n620 VSUBS 0.007329f
C661 B.n621 VSUBS 0.007329f
C662 B.n622 VSUBS 0.007329f
C663 B.n623 VSUBS 0.007329f
C664 B.n624 VSUBS 0.007329f
C665 B.n625 VSUBS 0.007329f
C666 B.n626 VSUBS 0.007329f
C667 B.n627 VSUBS 0.007329f
C668 B.n628 VSUBS 0.007329f
C669 B.n629 VSUBS 0.007329f
C670 B.n630 VSUBS 0.007329f
C671 B.n631 VSUBS 0.007329f
C672 B.n632 VSUBS 0.007329f
C673 B.n633 VSUBS 0.007329f
C674 B.n634 VSUBS 0.007329f
C675 B.n635 VSUBS 0.007329f
C676 B.n636 VSUBS 0.007329f
C677 B.n637 VSUBS 0.007329f
C678 B.n638 VSUBS 0.007329f
C679 B.n639 VSUBS 0.007329f
C680 B.n640 VSUBS 0.01626f
C681 B.n641 VSUBS 0.017152f
C682 B.n642 VSUBS 0.016477f
C683 B.n643 VSUBS 0.007329f
C684 B.n644 VSUBS 0.007329f
C685 B.n645 VSUBS 0.007329f
C686 B.n646 VSUBS 0.007329f
C687 B.n647 VSUBS 0.007329f
C688 B.n648 VSUBS 0.007329f
C689 B.n649 VSUBS 0.007329f
C690 B.n650 VSUBS 0.007329f
C691 B.n651 VSUBS 0.007329f
C692 B.n652 VSUBS 0.007329f
C693 B.n653 VSUBS 0.007329f
C694 B.n654 VSUBS 0.007329f
C695 B.n655 VSUBS 0.007329f
C696 B.n656 VSUBS 0.007329f
C697 B.n657 VSUBS 0.007329f
C698 B.n658 VSUBS 0.007329f
C699 B.n659 VSUBS 0.007329f
C700 B.n660 VSUBS 0.007329f
C701 B.n661 VSUBS 0.007329f
C702 B.n662 VSUBS 0.007329f
C703 B.n663 VSUBS 0.007329f
C704 B.n664 VSUBS 0.007329f
C705 B.n665 VSUBS 0.007329f
C706 B.n666 VSUBS 0.007329f
C707 B.n667 VSUBS 0.007329f
C708 B.n668 VSUBS 0.007329f
C709 B.n669 VSUBS 0.007329f
C710 B.n670 VSUBS 0.007329f
C711 B.n671 VSUBS 0.007329f
C712 B.n672 VSUBS 0.007329f
C713 B.n673 VSUBS 0.007329f
C714 B.n674 VSUBS 0.007329f
C715 B.n675 VSUBS 0.007329f
C716 B.n676 VSUBS 0.007329f
C717 B.n677 VSUBS 0.007329f
C718 B.n678 VSUBS 0.007329f
C719 B.n679 VSUBS 0.007329f
C720 B.n680 VSUBS 0.007329f
C721 B.n681 VSUBS 0.007329f
C722 B.n682 VSUBS 0.007329f
C723 B.n683 VSUBS 0.007329f
C724 B.n684 VSUBS 0.007329f
C725 B.n685 VSUBS 0.007329f
C726 B.n686 VSUBS 0.007329f
C727 B.n687 VSUBS 0.007329f
C728 B.n688 VSUBS 0.007329f
C729 B.n689 VSUBS 0.007329f
C730 B.n690 VSUBS 0.007329f
C731 B.n691 VSUBS 0.007329f
C732 B.n692 VSUBS 0.007329f
C733 B.n693 VSUBS 0.007329f
C734 B.n694 VSUBS 0.007329f
C735 B.n695 VSUBS 0.007329f
C736 B.n696 VSUBS 0.007329f
C737 B.n697 VSUBS 0.007329f
C738 B.n698 VSUBS 0.007329f
C739 B.n699 VSUBS 0.007329f
C740 B.n700 VSUBS 0.007329f
C741 B.n701 VSUBS 0.007329f
C742 B.n702 VSUBS 0.007329f
C743 B.n703 VSUBS 0.005066f
C744 B.n704 VSUBS 0.007329f
C745 B.n705 VSUBS 0.007329f
C746 B.n706 VSUBS 0.005928f
C747 B.n707 VSUBS 0.007329f
C748 B.n708 VSUBS 0.007329f
C749 B.n709 VSUBS 0.007329f
C750 B.n710 VSUBS 0.007329f
C751 B.n711 VSUBS 0.007329f
C752 B.n712 VSUBS 0.007329f
C753 B.n713 VSUBS 0.007329f
C754 B.n714 VSUBS 0.007329f
C755 B.n715 VSUBS 0.007329f
C756 B.n716 VSUBS 0.007329f
C757 B.n717 VSUBS 0.007329f
C758 B.n718 VSUBS 0.005928f
C759 B.n719 VSUBS 0.016981f
C760 B.n720 VSUBS 0.005066f
C761 B.n721 VSUBS 0.007329f
C762 B.n722 VSUBS 0.007329f
C763 B.n723 VSUBS 0.007329f
C764 B.n724 VSUBS 0.007329f
C765 B.n725 VSUBS 0.007329f
C766 B.n726 VSUBS 0.007329f
C767 B.n727 VSUBS 0.007329f
C768 B.n728 VSUBS 0.007329f
C769 B.n729 VSUBS 0.007329f
C770 B.n730 VSUBS 0.007329f
C771 B.n731 VSUBS 0.007329f
C772 B.n732 VSUBS 0.007329f
C773 B.n733 VSUBS 0.007329f
C774 B.n734 VSUBS 0.007329f
C775 B.n735 VSUBS 0.007329f
C776 B.n736 VSUBS 0.007329f
C777 B.n737 VSUBS 0.007329f
C778 B.n738 VSUBS 0.007329f
C779 B.n739 VSUBS 0.007329f
C780 B.n740 VSUBS 0.007329f
C781 B.n741 VSUBS 0.007329f
C782 B.n742 VSUBS 0.007329f
C783 B.n743 VSUBS 0.007329f
C784 B.n744 VSUBS 0.007329f
C785 B.n745 VSUBS 0.007329f
C786 B.n746 VSUBS 0.007329f
C787 B.n747 VSUBS 0.007329f
C788 B.n748 VSUBS 0.007329f
C789 B.n749 VSUBS 0.007329f
C790 B.n750 VSUBS 0.007329f
C791 B.n751 VSUBS 0.007329f
C792 B.n752 VSUBS 0.007329f
C793 B.n753 VSUBS 0.007329f
C794 B.n754 VSUBS 0.007329f
C795 B.n755 VSUBS 0.007329f
C796 B.n756 VSUBS 0.007329f
C797 B.n757 VSUBS 0.007329f
C798 B.n758 VSUBS 0.007329f
C799 B.n759 VSUBS 0.007329f
C800 B.n760 VSUBS 0.007329f
C801 B.n761 VSUBS 0.007329f
C802 B.n762 VSUBS 0.007329f
C803 B.n763 VSUBS 0.007329f
C804 B.n764 VSUBS 0.007329f
C805 B.n765 VSUBS 0.007329f
C806 B.n766 VSUBS 0.007329f
C807 B.n767 VSUBS 0.007329f
C808 B.n768 VSUBS 0.007329f
C809 B.n769 VSUBS 0.007329f
C810 B.n770 VSUBS 0.007329f
C811 B.n771 VSUBS 0.007329f
C812 B.n772 VSUBS 0.007329f
C813 B.n773 VSUBS 0.007329f
C814 B.n774 VSUBS 0.007329f
C815 B.n775 VSUBS 0.007329f
C816 B.n776 VSUBS 0.007329f
C817 B.n777 VSUBS 0.007329f
C818 B.n778 VSUBS 0.007329f
C819 B.n779 VSUBS 0.007329f
C820 B.n780 VSUBS 0.007329f
C821 B.n781 VSUBS 0.01737f
C822 B.n782 VSUBS 0.01737f
C823 B.n783 VSUBS 0.01626f
C824 B.n784 VSUBS 0.007329f
C825 B.n785 VSUBS 0.007329f
C826 B.n786 VSUBS 0.007329f
C827 B.n787 VSUBS 0.007329f
C828 B.n788 VSUBS 0.007329f
C829 B.n789 VSUBS 0.007329f
C830 B.n790 VSUBS 0.007329f
C831 B.n791 VSUBS 0.007329f
C832 B.n792 VSUBS 0.007329f
C833 B.n793 VSUBS 0.007329f
C834 B.n794 VSUBS 0.007329f
C835 B.n795 VSUBS 0.007329f
C836 B.n796 VSUBS 0.007329f
C837 B.n797 VSUBS 0.007329f
C838 B.n798 VSUBS 0.007329f
C839 B.n799 VSUBS 0.007329f
C840 B.n800 VSUBS 0.007329f
C841 B.n801 VSUBS 0.007329f
C842 B.n802 VSUBS 0.007329f
C843 B.n803 VSUBS 0.007329f
C844 B.n804 VSUBS 0.007329f
C845 B.n805 VSUBS 0.007329f
C846 B.n806 VSUBS 0.007329f
C847 B.n807 VSUBS 0.007329f
C848 B.n808 VSUBS 0.007329f
C849 B.n809 VSUBS 0.007329f
C850 B.n810 VSUBS 0.007329f
C851 B.n811 VSUBS 0.007329f
C852 B.n812 VSUBS 0.007329f
C853 B.n813 VSUBS 0.007329f
C854 B.n814 VSUBS 0.007329f
C855 B.n815 VSUBS 0.007329f
C856 B.n816 VSUBS 0.007329f
C857 B.n817 VSUBS 0.007329f
C858 B.n818 VSUBS 0.007329f
C859 B.n819 VSUBS 0.007329f
C860 B.n820 VSUBS 0.007329f
C861 B.n821 VSUBS 0.007329f
C862 B.n822 VSUBS 0.007329f
C863 B.n823 VSUBS 0.007329f
C864 B.n824 VSUBS 0.007329f
C865 B.n825 VSUBS 0.007329f
C866 B.n826 VSUBS 0.007329f
C867 B.n827 VSUBS 0.007329f
C868 B.n828 VSUBS 0.007329f
C869 B.n829 VSUBS 0.007329f
C870 B.n830 VSUBS 0.007329f
C871 B.n831 VSUBS 0.007329f
C872 B.n832 VSUBS 0.007329f
C873 B.n833 VSUBS 0.007329f
C874 B.n834 VSUBS 0.007329f
C875 B.n835 VSUBS 0.007329f
C876 B.n836 VSUBS 0.007329f
C877 B.n837 VSUBS 0.007329f
C878 B.n838 VSUBS 0.007329f
C879 B.n839 VSUBS 0.007329f
C880 B.n840 VSUBS 0.007329f
C881 B.n841 VSUBS 0.007329f
C882 B.n842 VSUBS 0.007329f
C883 B.n843 VSUBS 0.007329f
C884 B.n844 VSUBS 0.007329f
C885 B.n845 VSUBS 0.007329f
C886 B.n846 VSUBS 0.007329f
C887 B.n847 VSUBS 0.007329f
C888 B.n848 VSUBS 0.007329f
C889 B.n849 VSUBS 0.007329f
C890 B.n850 VSUBS 0.007329f
C891 B.n851 VSUBS 0.007329f
C892 B.n852 VSUBS 0.007329f
C893 B.n853 VSUBS 0.007329f
C894 B.n854 VSUBS 0.007329f
C895 B.n855 VSUBS 0.007329f
C896 B.n856 VSUBS 0.007329f
C897 B.n857 VSUBS 0.007329f
C898 B.n858 VSUBS 0.007329f
C899 B.n859 VSUBS 0.007329f
C900 B.n860 VSUBS 0.007329f
C901 B.n861 VSUBS 0.007329f
C902 B.n862 VSUBS 0.007329f
C903 B.n863 VSUBS 0.007329f
C904 B.n864 VSUBS 0.007329f
C905 B.n865 VSUBS 0.007329f
C906 B.n866 VSUBS 0.007329f
C907 B.n867 VSUBS 0.007329f
C908 B.n868 VSUBS 0.007329f
C909 B.n869 VSUBS 0.007329f
C910 B.n870 VSUBS 0.007329f
C911 B.n871 VSUBS 0.007329f
C912 B.n872 VSUBS 0.007329f
C913 B.n873 VSUBS 0.007329f
C914 B.n874 VSUBS 0.007329f
C915 B.n875 VSUBS 0.016596f
C916 VDD2.t4 VSUBS 0.286049f
C917 VDD2.t2 VSUBS 0.286049f
C918 VDD2.n0 VSUBS 2.28054f
C919 VDD2.t5 VSUBS 0.286049f
C920 VDD2.t7 VSUBS 0.286049f
C921 VDD2.n1 VSUBS 2.28054f
C922 VDD2.n2 VSUBS 4.99802f
C923 VDD2.t1 VSUBS 0.286049f
C924 VDD2.t6 VSUBS 0.286049f
C925 VDD2.n3 VSUBS 2.26176f
C926 VDD2.n4 VSUBS 4.13088f
C927 VDD2.t0 VSUBS 0.286049f
C928 VDD2.t3 VSUBS 0.286049f
C929 VDD2.n5 VSUBS 2.28049f
C930 VN.t0 VSUBS 2.7542f
C931 VN.n0 VSUBS 1.07721f
C932 VN.n1 VSUBS 0.025783f
C933 VN.n2 VSUBS 0.024357f
C934 VN.n3 VSUBS 0.025783f
C935 VN.t2 VSUBS 2.7542f
C936 VN.n4 VSUBS 0.968043f
C937 VN.n5 VSUBS 0.025783f
C938 VN.n6 VSUBS 0.020843f
C939 VN.n7 VSUBS 0.025783f
C940 VN.t5 VSUBS 2.7542f
C941 VN.n8 VSUBS 1.05593f
C942 VN.t3 VSUBS 3.07118f
C943 VN.n9 VSUBS 1.00536f
C944 VN.n10 VSUBS 0.299271f
C945 VN.n11 VSUBS 0.038563f
C946 VN.n12 VSUBS 0.048053f
C947 VN.n13 VSUBS 0.051243f
C948 VN.n14 VSUBS 0.025783f
C949 VN.n15 VSUBS 0.025783f
C950 VN.n16 VSUBS 0.025783f
C951 VN.n17 VSUBS 0.051243f
C952 VN.n18 VSUBS 0.048053f
C953 VN.n19 VSUBS 0.038563f
C954 VN.n20 VSUBS 0.025783f
C955 VN.n21 VSUBS 0.025783f
C956 VN.n22 VSUBS 0.033819f
C957 VN.n23 VSUBS 0.048053f
C958 VN.n24 VSUBS 0.051652f
C959 VN.n25 VSUBS 0.025783f
C960 VN.n26 VSUBS 0.025783f
C961 VN.n27 VSUBS 0.025783f
C962 VN.n28 VSUBS 0.047321f
C963 VN.n29 VSUBS 0.048053f
C964 VN.n30 VSUBS 0.043308f
C965 VN.n31 VSUBS 0.041613f
C966 VN.n32 VSUBS 0.056488f
C967 VN.t6 VSUBS 2.7542f
C968 VN.n33 VSUBS 1.07721f
C969 VN.n34 VSUBS 0.025783f
C970 VN.n35 VSUBS 0.024357f
C971 VN.n36 VSUBS 0.025783f
C972 VN.t1 VSUBS 2.7542f
C973 VN.n37 VSUBS 0.968043f
C974 VN.n38 VSUBS 0.025783f
C975 VN.n39 VSUBS 0.020843f
C976 VN.n40 VSUBS 0.025783f
C977 VN.t7 VSUBS 2.7542f
C978 VN.n41 VSUBS 1.05593f
C979 VN.t4 VSUBS 3.07118f
C980 VN.n42 VSUBS 1.00536f
C981 VN.n43 VSUBS 0.299271f
C982 VN.n44 VSUBS 0.038563f
C983 VN.n45 VSUBS 0.048053f
C984 VN.n46 VSUBS 0.051243f
C985 VN.n47 VSUBS 0.025783f
C986 VN.n48 VSUBS 0.025783f
C987 VN.n49 VSUBS 0.025783f
C988 VN.n50 VSUBS 0.051243f
C989 VN.n51 VSUBS 0.048053f
C990 VN.n52 VSUBS 0.038563f
C991 VN.n53 VSUBS 0.025783f
C992 VN.n54 VSUBS 0.025783f
C993 VN.n55 VSUBS 0.033819f
C994 VN.n56 VSUBS 0.048053f
C995 VN.n57 VSUBS 0.051652f
C996 VN.n58 VSUBS 0.025783f
C997 VN.n59 VSUBS 0.025783f
C998 VN.n60 VSUBS 0.025783f
C999 VN.n61 VSUBS 0.047321f
C1000 VN.n62 VSUBS 0.048053f
C1001 VN.n63 VSUBS 0.043308f
C1002 VN.n64 VSUBS 0.041613f
C1003 VN.n65 VSUBS 1.64985f
C1004 VDD1.t1 VSUBS 0.288509f
C1005 VDD1.t6 VSUBS 0.288509f
C1006 VDD1.n0 VSUBS 2.30179f
C1007 VDD1.t3 VSUBS 0.288509f
C1008 VDD1.t5 VSUBS 0.288509f
C1009 VDD1.n1 VSUBS 2.30016f
C1010 VDD1.t2 VSUBS 0.288509f
C1011 VDD1.t0 VSUBS 0.288509f
C1012 VDD1.n2 VSUBS 2.30016f
C1013 VDD1.n3 VSUBS 5.104f
C1014 VDD1.t4 VSUBS 0.288509f
C1015 VDD1.t7 VSUBS 0.288509f
C1016 VDD1.n4 VSUBS 2.2812f
C1017 VDD1.n5 VSUBS 4.20448f
C1018 VTAIL.t6 VSUBS 0.244327f
C1019 VTAIL.t3 VSUBS 0.244327f
C1020 VTAIL.n0 VSUBS 1.80822f
C1021 VTAIL.n1 VSUBS 0.80986f
C1022 VTAIL.n2 VSUBS 0.014556f
C1023 VTAIL.n3 VSUBS 0.032752f
C1024 VTAIL.n4 VSUBS 0.014672f
C1025 VTAIL.n5 VSUBS 0.025787f
C1026 VTAIL.n6 VSUBS 0.013857f
C1027 VTAIL.n7 VSUBS 0.032752f
C1028 VTAIL.n8 VSUBS 0.014672f
C1029 VTAIL.n9 VSUBS 0.025787f
C1030 VTAIL.n10 VSUBS 0.013857f
C1031 VTAIL.n11 VSUBS 0.032752f
C1032 VTAIL.n12 VSUBS 0.014672f
C1033 VTAIL.n13 VSUBS 0.025787f
C1034 VTAIL.n14 VSUBS 0.013857f
C1035 VTAIL.n15 VSUBS 0.032752f
C1036 VTAIL.n16 VSUBS 0.014672f
C1037 VTAIL.n17 VSUBS 0.025787f
C1038 VTAIL.n18 VSUBS 0.013857f
C1039 VTAIL.n19 VSUBS 0.032752f
C1040 VTAIL.n20 VSUBS 0.014672f
C1041 VTAIL.n21 VSUBS 1.29417f
C1042 VTAIL.n22 VSUBS 0.013857f
C1043 VTAIL.t4 VSUBS 0.069928f
C1044 VTAIL.n23 VSUBS 0.158886f
C1045 VTAIL.n24 VSUBS 0.020836f
C1046 VTAIL.n25 VSUBS 0.024564f
C1047 VTAIL.n26 VSUBS 0.032752f
C1048 VTAIL.n27 VSUBS 0.014672f
C1049 VTAIL.n28 VSUBS 0.013857f
C1050 VTAIL.n29 VSUBS 0.025787f
C1051 VTAIL.n30 VSUBS 0.025787f
C1052 VTAIL.n31 VSUBS 0.013857f
C1053 VTAIL.n32 VSUBS 0.014672f
C1054 VTAIL.n33 VSUBS 0.032752f
C1055 VTAIL.n34 VSUBS 0.032752f
C1056 VTAIL.n35 VSUBS 0.014672f
C1057 VTAIL.n36 VSUBS 0.013857f
C1058 VTAIL.n37 VSUBS 0.025787f
C1059 VTAIL.n38 VSUBS 0.025787f
C1060 VTAIL.n39 VSUBS 0.013857f
C1061 VTAIL.n40 VSUBS 0.014672f
C1062 VTAIL.n41 VSUBS 0.032752f
C1063 VTAIL.n42 VSUBS 0.032752f
C1064 VTAIL.n43 VSUBS 0.014672f
C1065 VTAIL.n44 VSUBS 0.013857f
C1066 VTAIL.n45 VSUBS 0.025787f
C1067 VTAIL.n46 VSUBS 0.025787f
C1068 VTAIL.n47 VSUBS 0.013857f
C1069 VTAIL.n48 VSUBS 0.014672f
C1070 VTAIL.n49 VSUBS 0.032752f
C1071 VTAIL.n50 VSUBS 0.032752f
C1072 VTAIL.n51 VSUBS 0.014672f
C1073 VTAIL.n52 VSUBS 0.013857f
C1074 VTAIL.n53 VSUBS 0.025787f
C1075 VTAIL.n54 VSUBS 0.025787f
C1076 VTAIL.n55 VSUBS 0.013857f
C1077 VTAIL.n56 VSUBS 0.014672f
C1078 VTAIL.n57 VSUBS 0.032752f
C1079 VTAIL.n58 VSUBS 0.032752f
C1080 VTAIL.n59 VSUBS 0.014672f
C1081 VTAIL.n60 VSUBS 0.013857f
C1082 VTAIL.n61 VSUBS 0.025787f
C1083 VTAIL.n62 VSUBS 0.067708f
C1084 VTAIL.n63 VSUBS 0.013857f
C1085 VTAIL.n64 VSUBS 0.014672f
C1086 VTAIL.n65 VSUBS 0.074082f
C1087 VTAIL.n66 VSUBS 0.049892f
C1088 VTAIL.n67 VSUBS 0.322319f
C1089 VTAIL.n68 VSUBS 0.014556f
C1090 VTAIL.n69 VSUBS 0.032752f
C1091 VTAIL.n70 VSUBS 0.014672f
C1092 VTAIL.n71 VSUBS 0.025787f
C1093 VTAIL.n72 VSUBS 0.013857f
C1094 VTAIL.n73 VSUBS 0.032752f
C1095 VTAIL.n74 VSUBS 0.014672f
C1096 VTAIL.n75 VSUBS 0.025787f
C1097 VTAIL.n76 VSUBS 0.013857f
C1098 VTAIL.n77 VSUBS 0.032752f
C1099 VTAIL.n78 VSUBS 0.014672f
C1100 VTAIL.n79 VSUBS 0.025787f
C1101 VTAIL.n80 VSUBS 0.013857f
C1102 VTAIL.n81 VSUBS 0.032752f
C1103 VTAIL.n82 VSUBS 0.014672f
C1104 VTAIL.n83 VSUBS 0.025787f
C1105 VTAIL.n84 VSUBS 0.013857f
C1106 VTAIL.n85 VSUBS 0.032752f
C1107 VTAIL.n86 VSUBS 0.014672f
C1108 VTAIL.n87 VSUBS 1.29417f
C1109 VTAIL.n88 VSUBS 0.013857f
C1110 VTAIL.t14 VSUBS 0.069928f
C1111 VTAIL.n89 VSUBS 0.158886f
C1112 VTAIL.n90 VSUBS 0.020836f
C1113 VTAIL.n91 VSUBS 0.024564f
C1114 VTAIL.n92 VSUBS 0.032752f
C1115 VTAIL.n93 VSUBS 0.014672f
C1116 VTAIL.n94 VSUBS 0.013857f
C1117 VTAIL.n95 VSUBS 0.025787f
C1118 VTAIL.n96 VSUBS 0.025787f
C1119 VTAIL.n97 VSUBS 0.013857f
C1120 VTAIL.n98 VSUBS 0.014672f
C1121 VTAIL.n99 VSUBS 0.032752f
C1122 VTAIL.n100 VSUBS 0.032752f
C1123 VTAIL.n101 VSUBS 0.014672f
C1124 VTAIL.n102 VSUBS 0.013857f
C1125 VTAIL.n103 VSUBS 0.025787f
C1126 VTAIL.n104 VSUBS 0.025787f
C1127 VTAIL.n105 VSUBS 0.013857f
C1128 VTAIL.n106 VSUBS 0.014672f
C1129 VTAIL.n107 VSUBS 0.032752f
C1130 VTAIL.n108 VSUBS 0.032752f
C1131 VTAIL.n109 VSUBS 0.014672f
C1132 VTAIL.n110 VSUBS 0.013857f
C1133 VTAIL.n111 VSUBS 0.025787f
C1134 VTAIL.n112 VSUBS 0.025787f
C1135 VTAIL.n113 VSUBS 0.013857f
C1136 VTAIL.n114 VSUBS 0.014672f
C1137 VTAIL.n115 VSUBS 0.032752f
C1138 VTAIL.n116 VSUBS 0.032752f
C1139 VTAIL.n117 VSUBS 0.014672f
C1140 VTAIL.n118 VSUBS 0.013857f
C1141 VTAIL.n119 VSUBS 0.025787f
C1142 VTAIL.n120 VSUBS 0.025787f
C1143 VTAIL.n121 VSUBS 0.013857f
C1144 VTAIL.n122 VSUBS 0.014672f
C1145 VTAIL.n123 VSUBS 0.032752f
C1146 VTAIL.n124 VSUBS 0.032752f
C1147 VTAIL.n125 VSUBS 0.014672f
C1148 VTAIL.n126 VSUBS 0.013857f
C1149 VTAIL.n127 VSUBS 0.025787f
C1150 VTAIL.n128 VSUBS 0.067708f
C1151 VTAIL.n129 VSUBS 0.013857f
C1152 VTAIL.n130 VSUBS 0.014672f
C1153 VTAIL.n131 VSUBS 0.074082f
C1154 VTAIL.n132 VSUBS 0.049892f
C1155 VTAIL.n133 VSUBS 0.322319f
C1156 VTAIL.t12 VSUBS 0.244327f
C1157 VTAIL.t13 VSUBS 0.244327f
C1158 VTAIL.n134 VSUBS 1.80822f
C1159 VTAIL.n135 VSUBS 1.06289f
C1160 VTAIL.n136 VSUBS 0.014556f
C1161 VTAIL.n137 VSUBS 0.032752f
C1162 VTAIL.n138 VSUBS 0.014672f
C1163 VTAIL.n139 VSUBS 0.025787f
C1164 VTAIL.n140 VSUBS 0.013857f
C1165 VTAIL.n141 VSUBS 0.032752f
C1166 VTAIL.n142 VSUBS 0.014672f
C1167 VTAIL.n143 VSUBS 0.025787f
C1168 VTAIL.n144 VSUBS 0.013857f
C1169 VTAIL.n145 VSUBS 0.032752f
C1170 VTAIL.n146 VSUBS 0.014672f
C1171 VTAIL.n147 VSUBS 0.025787f
C1172 VTAIL.n148 VSUBS 0.013857f
C1173 VTAIL.n149 VSUBS 0.032752f
C1174 VTAIL.n150 VSUBS 0.014672f
C1175 VTAIL.n151 VSUBS 0.025787f
C1176 VTAIL.n152 VSUBS 0.013857f
C1177 VTAIL.n153 VSUBS 0.032752f
C1178 VTAIL.n154 VSUBS 0.014672f
C1179 VTAIL.n155 VSUBS 1.29417f
C1180 VTAIL.n156 VSUBS 0.013857f
C1181 VTAIL.t9 VSUBS 0.069928f
C1182 VTAIL.n157 VSUBS 0.158886f
C1183 VTAIL.n158 VSUBS 0.020836f
C1184 VTAIL.n159 VSUBS 0.024564f
C1185 VTAIL.n160 VSUBS 0.032752f
C1186 VTAIL.n161 VSUBS 0.014672f
C1187 VTAIL.n162 VSUBS 0.013857f
C1188 VTAIL.n163 VSUBS 0.025787f
C1189 VTAIL.n164 VSUBS 0.025787f
C1190 VTAIL.n165 VSUBS 0.013857f
C1191 VTAIL.n166 VSUBS 0.014672f
C1192 VTAIL.n167 VSUBS 0.032752f
C1193 VTAIL.n168 VSUBS 0.032752f
C1194 VTAIL.n169 VSUBS 0.014672f
C1195 VTAIL.n170 VSUBS 0.013857f
C1196 VTAIL.n171 VSUBS 0.025787f
C1197 VTAIL.n172 VSUBS 0.025787f
C1198 VTAIL.n173 VSUBS 0.013857f
C1199 VTAIL.n174 VSUBS 0.014672f
C1200 VTAIL.n175 VSUBS 0.032752f
C1201 VTAIL.n176 VSUBS 0.032752f
C1202 VTAIL.n177 VSUBS 0.014672f
C1203 VTAIL.n178 VSUBS 0.013857f
C1204 VTAIL.n179 VSUBS 0.025787f
C1205 VTAIL.n180 VSUBS 0.025787f
C1206 VTAIL.n181 VSUBS 0.013857f
C1207 VTAIL.n182 VSUBS 0.014672f
C1208 VTAIL.n183 VSUBS 0.032752f
C1209 VTAIL.n184 VSUBS 0.032752f
C1210 VTAIL.n185 VSUBS 0.014672f
C1211 VTAIL.n186 VSUBS 0.013857f
C1212 VTAIL.n187 VSUBS 0.025787f
C1213 VTAIL.n188 VSUBS 0.025787f
C1214 VTAIL.n189 VSUBS 0.013857f
C1215 VTAIL.n190 VSUBS 0.014672f
C1216 VTAIL.n191 VSUBS 0.032752f
C1217 VTAIL.n192 VSUBS 0.032752f
C1218 VTAIL.n193 VSUBS 0.014672f
C1219 VTAIL.n194 VSUBS 0.013857f
C1220 VTAIL.n195 VSUBS 0.025787f
C1221 VTAIL.n196 VSUBS 0.067708f
C1222 VTAIL.n197 VSUBS 0.013857f
C1223 VTAIL.n198 VSUBS 0.014672f
C1224 VTAIL.n199 VSUBS 0.074082f
C1225 VTAIL.n200 VSUBS 0.049892f
C1226 VTAIL.n201 VSUBS 1.75028f
C1227 VTAIL.n202 VSUBS 0.014556f
C1228 VTAIL.n203 VSUBS 0.032752f
C1229 VTAIL.n204 VSUBS 0.014672f
C1230 VTAIL.n205 VSUBS 0.025787f
C1231 VTAIL.n206 VSUBS 0.013857f
C1232 VTAIL.n207 VSUBS 0.032752f
C1233 VTAIL.n208 VSUBS 0.014672f
C1234 VTAIL.n209 VSUBS 0.025787f
C1235 VTAIL.n210 VSUBS 0.013857f
C1236 VTAIL.n211 VSUBS 0.032752f
C1237 VTAIL.n212 VSUBS 0.014672f
C1238 VTAIL.n213 VSUBS 0.025787f
C1239 VTAIL.n214 VSUBS 0.013857f
C1240 VTAIL.n215 VSUBS 0.032752f
C1241 VTAIL.n216 VSUBS 0.014672f
C1242 VTAIL.n217 VSUBS 0.025787f
C1243 VTAIL.n218 VSUBS 0.013857f
C1244 VTAIL.n219 VSUBS 0.032752f
C1245 VTAIL.n220 VSUBS 0.014672f
C1246 VTAIL.n221 VSUBS 1.29417f
C1247 VTAIL.n222 VSUBS 0.013857f
C1248 VTAIL.t5 VSUBS 0.069928f
C1249 VTAIL.n223 VSUBS 0.158886f
C1250 VTAIL.n224 VSUBS 0.020836f
C1251 VTAIL.n225 VSUBS 0.024564f
C1252 VTAIL.n226 VSUBS 0.032752f
C1253 VTAIL.n227 VSUBS 0.014672f
C1254 VTAIL.n228 VSUBS 0.013857f
C1255 VTAIL.n229 VSUBS 0.025787f
C1256 VTAIL.n230 VSUBS 0.025787f
C1257 VTAIL.n231 VSUBS 0.013857f
C1258 VTAIL.n232 VSUBS 0.014672f
C1259 VTAIL.n233 VSUBS 0.032752f
C1260 VTAIL.n234 VSUBS 0.032752f
C1261 VTAIL.n235 VSUBS 0.014672f
C1262 VTAIL.n236 VSUBS 0.013857f
C1263 VTAIL.n237 VSUBS 0.025787f
C1264 VTAIL.n238 VSUBS 0.025787f
C1265 VTAIL.n239 VSUBS 0.013857f
C1266 VTAIL.n240 VSUBS 0.014672f
C1267 VTAIL.n241 VSUBS 0.032752f
C1268 VTAIL.n242 VSUBS 0.032752f
C1269 VTAIL.n243 VSUBS 0.014672f
C1270 VTAIL.n244 VSUBS 0.013857f
C1271 VTAIL.n245 VSUBS 0.025787f
C1272 VTAIL.n246 VSUBS 0.025787f
C1273 VTAIL.n247 VSUBS 0.013857f
C1274 VTAIL.n248 VSUBS 0.014672f
C1275 VTAIL.n249 VSUBS 0.032752f
C1276 VTAIL.n250 VSUBS 0.032752f
C1277 VTAIL.n251 VSUBS 0.014672f
C1278 VTAIL.n252 VSUBS 0.013857f
C1279 VTAIL.n253 VSUBS 0.025787f
C1280 VTAIL.n254 VSUBS 0.025787f
C1281 VTAIL.n255 VSUBS 0.013857f
C1282 VTAIL.n256 VSUBS 0.014672f
C1283 VTAIL.n257 VSUBS 0.032752f
C1284 VTAIL.n258 VSUBS 0.032752f
C1285 VTAIL.n259 VSUBS 0.014672f
C1286 VTAIL.n260 VSUBS 0.013857f
C1287 VTAIL.n261 VSUBS 0.025787f
C1288 VTAIL.n262 VSUBS 0.067708f
C1289 VTAIL.n263 VSUBS 0.013857f
C1290 VTAIL.n264 VSUBS 0.014672f
C1291 VTAIL.n265 VSUBS 0.074082f
C1292 VTAIL.n266 VSUBS 0.049892f
C1293 VTAIL.n267 VSUBS 1.75028f
C1294 VTAIL.t2 VSUBS 0.244327f
C1295 VTAIL.t7 VSUBS 0.244327f
C1296 VTAIL.n268 VSUBS 1.80823f
C1297 VTAIL.n269 VSUBS 1.06289f
C1298 VTAIL.n270 VSUBS 0.014556f
C1299 VTAIL.n271 VSUBS 0.032752f
C1300 VTAIL.n272 VSUBS 0.014672f
C1301 VTAIL.n273 VSUBS 0.025787f
C1302 VTAIL.n274 VSUBS 0.013857f
C1303 VTAIL.n275 VSUBS 0.032752f
C1304 VTAIL.n276 VSUBS 0.014672f
C1305 VTAIL.n277 VSUBS 0.025787f
C1306 VTAIL.n278 VSUBS 0.013857f
C1307 VTAIL.n279 VSUBS 0.032752f
C1308 VTAIL.n280 VSUBS 0.014672f
C1309 VTAIL.n281 VSUBS 0.025787f
C1310 VTAIL.n282 VSUBS 0.013857f
C1311 VTAIL.n283 VSUBS 0.032752f
C1312 VTAIL.n284 VSUBS 0.014672f
C1313 VTAIL.n285 VSUBS 0.025787f
C1314 VTAIL.n286 VSUBS 0.013857f
C1315 VTAIL.n287 VSUBS 0.032752f
C1316 VTAIL.n288 VSUBS 0.014672f
C1317 VTAIL.n289 VSUBS 1.29417f
C1318 VTAIL.n290 VSUBS 0.013857f
C1319 VTAIL.t0 VSUBS 0.069928f
C1320 VTAIL.n291 VSUBS 0.158886f
C1321 VTAIL.n292 VSUBS 0.020836f
C1322 VTAIL.n293 VSUBS 0.024564f
C1323 VTAIL.n294 VSUBS 0.032752f
C1324 VTAIL.n295 VSUBS 0.014672f
C1325 VTAIL.n296 VSUBS 0.013857f
C1326 VTAIL.n297 VSUBS 0.025787f
C1327 VTAIL.n298 VSUBS 0.025787f
C1328 VTAIL.n299 VSUBS 0.013857f
C1329 VTAIL.n300 VSUBS 0.014672f
C1330 VTAIL.n301 VSUBS 0.032752f
C1331 VTAIL.n302 VSUBS 0.032752f
C1332 VTAIL.n303 VSUBS 0.014672f
C1333 VTAIL.n304 VSUBS 0.013857f
C1334 VTAIL.n305 VSUBS 0.025787f
C1335 VTAIL.n306 VSUBS 0.025787f
C1336 VTAIL.n307 VSUBS 0.013857f
C1337 VTAIL.n308 VSUBS 0.014672f
C1338 VTAIL.n309 VSUBS 0.032752f
C1339 VTAIL.n310 VSUBS 0.032752f
C1340 VTAIL.n311 VSUBS 0.014672f
C1341 VTAIL.n312 VSUBS 0.013857f
C1342 VTAIL.n313 VSUBS 0.025787f
C1343 VTAIL.n314 VSUBS 0.025787f
C1344 VTAIL.n315 VSUBS 0.013857f
C1345 VTAIL.n316 VSUBS 0.014672f
C1346 VTAIL.n317 VSUBS 0.032752f
C1347 VTAIL.n318 VSUBS 0.032752f
C1348 VTAIL.n319 VSUBS 0.014672f
C1349 VTAIL.n320 VSUBS 0.013857f
C1350 VTAIL.n321 VSUBS 0.025787f
C1351 VTAIL.n322 VSUBS 0.025787f
C1352 VTAIL.n323 VSUBS 0.013857f
C1353 VTAIL.n324 VSUBS 0.014672f
C1354 VTAIL.n325 VSUBS 0.032752f
C1355 VTAIL.n326 VSUBS 0.032752f
C1356 VTAIL.n327 VSUBS 0.014672f
C1357 VTAIL.n328 VSUBS 0.013857f
C1358 VTAIL.n329 VSUBS 0.025787f
C1359 VTAIL.n330 VSUBS 0.067708f
C1360 VTAIL.n331 VSUBS 0.013857f
C1361 VTAIL.n332 VSUBS 0.014672f
C1362 VTAIL.n333 VSUBS 0.074082f
C1363 VTAIL.n334 VSUBS 0.049892f
C1364 VTAIL.n335 VSUBS 0.322319f
C1365 VTAIL.n336 VSUBS 0.014556f
C1366 VTAIL.n337 VSUBS 0.032752f
C1367 VTAIL.n338 VSUBS 0.014672f
C1368 VTAIL.n339 VSUBS 0.025787f
C1369 VTAIL.n340 VSUBS 0.013857f
C1370 VTAIL.n341 VSUBS 0.032752f
C1371 VTAIL.n342 VSUBS 0.014672f
C1372 VTAIL.n343 VSUBS 0.025787f
C1373 VTAIL.n344 VSUBS 0.013857f
C1374 VTAIL.n345 VSUBS 0.032752f
C1375 VTAIL.n346 VSUBS 0.014672f
C1376 VTAIL.n347 VSUBS 0.025787f
C1377 VTAIL.n348 VSUBS 0.013857f
C1378 VTAIL.n349 VSUBS 0.032752f
C1379 VTAIL.n350 VSUBS 0.014672f
C1380 VTAIL.n351 VSUBS 0.025787f
C1381 VTAIL.n352 VSUBS 0.013857f
C1382 VTAIL.n353 VSUBS 0.032752f
C1383 VTAIL.n354 VSUBS 0.014672f
C1384 VTAIL.n355 VSUBS 1.29417f
C1385 VTAIL.n356 VSUBS 0.013857f
C1386 VTAIL.t15 VSUBS 0.069928f
C1387 VTAIL.n357 VSUBS 0.158886f
C1388 VTAIL.n358 VSUBS 0.020836f
C1389 VTAIL.n359 VSUBS 0.024564f
C1390 VTAIL.n360 VSUBS 0.032752f
C1391 VTAIL.n361 VSUBS 0.014672f
C1392 VTAIL.n362 VSUBS 0.013857f
C1393 VTAIL.n363 VSUBS 0.025787f
C1394 VTAIL.n364 VSUBS 0.025787f
C1395 VTAIL.n365 VSUBS 0.013857f
C1396 VTAIL.n366 VSUBS 0.014672f
C1397 VTAIL.n367 VSUBS 0.032752f
C1398 VTAIL.n368 VSUBS 0.032752f
C1399 VTAIL.n369 VSUBS 0.014672f
C1400 VTAIL.n370 VSUBS 0.013857f
C1401 VTAIL.n371 VSUBS 0.025787f
C1402 VTAIL.n372 VSUBS 0.025787f
C1403 VTAIL.n373 VSUBS 0.013857f
C1404 VTAIL.n374 VSUBS 0.014672f
C1405 VTAIL.n375 VSUBS 0.032752f
C1406 VTAIL.n376 VSUBS 0.032752f
C1407 VTAIL.n377 VSUBS 0.014672f
C1408 VTAIL.n378 VSUBS 0.013857f
C1409 VTAIL.n379 VSUBS 0.025787f
C1410 VTAIL.n380 VSUBS 0.025787f
C1411 VTAIL.n381 VSUBS 0.013857f
C1412 VTAIL.n382 VSUBS 0.014672f
C1413 VTAIL.n383 VSUBS 0.032752f
C1414 VTAIL.n384 VSUBS 0.032752f
C1415 VTAIL.n385 VSUBS 0.014672f
C1416 VTAIL.n386 VSUBS 0.013857f
C1417 VTAIL.n387 VSUBS 0.025787f
C1418 VTAIL.n388 VSUBS 0.025787f
C1419 VTAIL.n389 VSUBS 0.013857f
C1420 VTAIL.n390 VSUBS 0.014672f
C1421 VTAIL.n391 VSUBS 0.032752f
C1422 VTAIL.n392 VSUBS 0.032752f
C1423 VTAIL.n393 VSUBS 0.014672f
C1424 VTAIL.n394 VSUBS 0.013857f
C1425 VTAIL.n395 VSUBS 0.025787f
C1426 VTAIL.n396 VSUBS 0.067708f
C1427 VTAIL.n397 VSUBS 0.013857f
C1428 VTAIL.n398 VSUBS 0.014672f
C1429 VTAIL.n399 VSUBS 0.074082f
C1430 VTAIL.n400 VSUBS 0.049892f
C1431 VTAIL.n401 VSUBS 0.322319f
C1432 VTAIL.t8 VSUBS 0.244327f
C1433 VTAIL.t10 VSUBS 0.244327f
C1434 VTAIL.n402 VSUBS 1.80823f
C1435 VTAIL.n403 VSUBS 1.06289f
C1436 VTAIL.n404 VSUBS 0.014556f
C1437 VTAIL.n405 VSUBS 0.032752f
C1438 VTAIL.n406 VSUBS 0.014672f
C1439 VTAIL.n407 VSUBS 0.025787f
C1440 VTAIL.n408 VSUBS 0.013857f
C1441 VTAIL.n409 VSUBS 0.032752f
C1442 VTAIL.n410 VSUBS 0.014672f
C1443 VTAIL.n411 VSUBS 0.025787f
C1444 VTAIL.n412 VSUBS 0.013857f
C1445 VTAIL.n413 VSUBS 0.032752f
C1446 VTAIL.n414 VSUBS 0.014672f
C1447 VTAIL.n415 VSUBS 0.025787f
C1448 VTAIL.n416 VSUBS 0.013857f
C1449 VTAIL.n417 VSUBS 0.032752f
C1450 VTAIL.n418 VSUBS 0.014672f
C1451 VTAIL.n419 VSUBS 0.025787f
C1452 VTAIL.n420 VSUBS 0.013857f
C1453 VTAIL.n421 VSUBS 0.032752f
C1454 VTAIL.n422 VSUBS 0.014672f
C1455 VTAIL.n423 VSUBS 1.29417f
C1456 VTAIL.n424 VSUBS 0.013857f
C1457 VTAIL.t11 VSUBS 0.069928f
C1458 VTAIL.n425 VSUBS 0.158886f
C1459 VTAIL.n426 VSUBS 0.020836f
C1460 VTAIL.n427 VSUBS 0.024564f
C1461 VTAIL.n428 VSUBS 0.032752f
C1462 VTAIL.n429 VSUBS 0.014672f
C1463 VTAIL.n430 VSUBS 0.013857f
C1464 VTAIL.n431 VSUBS 0.025787f
C1465 VTAIL.n432 VSUBS 0.025787f
C1466 VTAIL.n433 VSUBS 0.013857f
C1467 VTAIL.n434 VSUBS 0.014672f
C1468 VTAIL.n435 VSUBS 0.032752f
C1469 VTAIL.n436 VSUBS 0.032752f
C1470 VTAIL.n437 VSUBS 0.014672f
C1471 VTAIL.n438 VSUBS 0.013857f
C1472 VTAIL.n439 VSUBS 0.025787f
C1473 VTAIL.n440 VSUBS 0.025787f
C1474 VTAIL.n441 VSUBS 0.013857f
C1475 VTAIL.n442 VSUBS 0.014672f
C1476 VTAIL.n443 VSUBS 0.032752f
C1477 VTAIL.n444 VSUBS 0.032752f
C1478 VTAIL.n445 VSUBS 0.014672f
C1479 VTAIL.n446 VSUBS 0.013857f
C1480 VTAIL.n447 VSUBS 0.025787f
C1481 VTAIL.n448 VSUBS 0.025787f
C1482 VTAIL.n449 VSUBS 0.013857f
C1483 VTAIL.n450 VSUBS 0.014672f
C1484 VTAIL.n451 VSUBS 0.032752f
C1485 VTAIL.n452 VSUBS 0.032752f
C1486 VTAIL.n453 VSUBS 0.014672f
C1487 VTAIL.n454 VSUBS 0.013857f
C1488 VTAIL.n455 VSUBS 0.025787f
C1489 VTAIL.n456 VSUBS 0.025787f
C1490 VTAIL.n457 VSUBS 0.013857f
C1491 VTAIL.n458 VSUBS 0.014672f
C1492 VTAIL.n459 VSUBS 0.032752f
C1493 VTAIL.n460 VSUBS 0.032752f
C1494 VTAIL.n461 VSUBS 0.014672f
C1495 VTAIL.n462 VSUBS 0.013857f
C1496 VTAIL.n463 VSUBS 0.025787f
C1497 VTAIL.n464 VSUBS 0.067708f
C1498 VTAIL.n465 VSUBS 0.013857f
C1499 VTAIL.n466 VSUBS 0.014672f
C1500 VTAIL.n467 VSUBS 0.074082f
C1501 VTAIL.n468 VSUBS 0.049892f
C1502 VTAIL.n469 VSUBS 1.75028f
C1503 VTAIL.n470 VSUBS 0.014556f
C1504 VTAIL.n471 VSUBS 0.032752f
C1505 VTAIL.n472 VSUBS 0.014672f
C1506 VTAIL.n473 VSUBS 0.025787f
C1507 VTAIL.n474 VSUBS 0.013857f
C1508 VTAIL.n475 VSUBS 0.032752f
C1509 VTAIL.n476 VSUBS 0.014672f
C1510 VTAIL.n477 VSUBS 0.025787f
C1511 VTAIL.n478 VSUBS 0.013857f
C1512 VTAIL.n479 VSUBS 0.032752f
C1513 VTAIL.n480 VSUBS 0.014672f
C1514 VTAIL.n481 VSUBS 0.025787f
C1515 VTAIL.n482 VSUBS 0.013857f
C1516 VTAIL.n483 VSUBS 0.032752f
C1517 VTAIL.n484 VSUBS 0.014672f
C1518 VTAIL.n485 VSUBS 0.025787f
C1519 VTAIL.n486 VSUBS 0.013857f
C1520 VTAIL.n487 VSUBS 0.032752f
C1521 VTAIL.n488 VSUBS 0.014672f
C1522 VTAIL.n489 VSUBS 1.29417f
C1523 VTAIL.n490 VSUBS 0.013857f
C1524 VTAIL.t1 VSUBS 0.069928f
C1525 VTAIL.n491 VSUBS 0.158886f
C1526 VTAIL.n492 VSUBS 0.020836f
C1527 VTAIL.n493 VSUBS 0.024564f
C1528 VTAIL.n494 VSUBS 0.032752f
C1529 VTAIL.n495 VSUBS 0.014672f
C1530 VTAIL.n496 VSUBS 0.013857f
C1531 VTAIL.n497 VSUBS 0.025787f
C1532 VTAIL.n498 VSUBS 0.025787f
C1533 VTAIL.n499 VSUBS 0.013857f
C1534 VTAIL.n500 VSUBS 0.014672f
C1535 VTAIL.n501 VSUBS 0.032752f
C1536 VTAIL.n502 VSUBS 0.032752f
C1537 VTAIL.n503 VSUBS 0.014672f
C1538 VTAIL.n504 VSUBS 0.013857f
C1539 VTAIL.n505 VSUBS 0.025787f
C1540 VTAIL.n506 VSUBS 0.025787f
C1541 VTAIL.n507 VSUBS 0.013857f
C1542 VTAIL.n508 VSUBS 0.014672f
C1543 VTAIL.n509 VSUBS 0.032752f
C1544 VTAIL.n510 VSUBS 0.032752f
C1545 VTAIL.n511 VSUBS 0.014672f
C1546 VTAIL.n512 VSUBS 0.013857f
C1547 VTAIL.n513 VSUBS 0.025787f
C1548 VTAIL.n514 VSUBS 0.025787f
C1549 VTAIL.n515 VSUBS 0.013857f
C1550 VTAIL.n516 VSUBS 0.014672f
C1551 VTAIL.n517 VSUBS 0.032752f
C1552 VTAIL.n518 VSUBS 0.032752f
C1553 VTAIL.n519 VSUBS 0.014672f
C1554 VTAIL.n520 VSUBS 0.013857f
C1555 VTAIL.n521 VSUBS 0.025787f
C1556 VTAIL.n522 VSUBS 0.025787f
C1557 VTAIL.n523 VSUBS 0.013857f
C1558 VTAIL.n524 VSUBS 0.014672f
C1559 VTAIL.n525 VSUBS 0.032752f
C1560 VTAIL.n526 VSUBS 0.032752f
C1561 VTAIL.n527 VSUBS 0.014672f
C1562 VTAIL.n528 VSUBS 0.013857f
C1563 VTAIL.n529 VSUBS 0.025787f
C1564 VTAIL.n530 VSUBS 0.067708f
C1565 VTAIL.n531 VSUBS 0.013857f
C1566 VTAIL.n532 VSUBS 0.014672f
C1567 VTAIL.n533 VSUBS 0.074082f
C1568 VTAIL.n534 VSUBS 0.049892f
C1569 VTAIL.n535 VSUBS 1.74545f
C1570 VP.t7 VSUBS 3.01984f
C1571 VP.n0 VSUBS 1.18111f
C1572 VP.n1 VSUBS 0.02827f
C1573 VP.n2 VSUBS 0.026706f
C1574 VP.n3 VSUBS 0.02827f
C1575 VP.t5 VSUBS 3.01984f
C1576 VP.n4 VSUBS 1.06141f
C1577 VP.n5 VSUBS 0.02827f
C1578 VP.n6 VSUBS 0.022853f
C1579 VP.n7 VSUBS 0.02827f
C1580 VP.t2 VSUBS 3.01984f
C1581 VP.n8 VSUBS 1.06141f
C1582 VP.n9 VSUBS 0.02827f
C1583 VP.n10 VSUBS 0.026706f
C1584 VP.n11 VSUBS 0.02827f
C1585 VP.t4 VSUBS 3.01984f
C1586 VP.n12 VSUBS 1.18111f
C1587 VP.t0 VSUBS 3.01984f
C1588 VP.n13 VSUBS 1.18111f
C1589 VP.n14 VSUBS 0.02827f
C1590 VP.n15 VSUBS 0.026706f
C1591 VP.n16 VSUBS 0.02827f
C1592 VP.t3 VSUBS 3.01984f
C1593 VP.n17 VSUBS 1.06141f
C1594 VP.n18 VSUBS 0.02827f
C1595 VP.n19 VSUBS 0.022853f
C1596 VP.n20 VSUBS 0.02827f
C1597 VP.t1 VSUBS 3.01984f
C1598 VP.n21 VSUBS 1.15778f
C1599 VP.t6 VSUBS 3.3674f
C1600 VP.n22 VSUBS 1.10233f
C1601 VP.n23 VSUBS 0.328137f
C1602 VP.n24 VSUBS 0.042283f
C1603 VP.n25 VSUBS 0.052688f
C1604 VP.n26 VSUBS 0.056186f
C1605 VP.n27 VSUBS 0.02827f
C1606 VP.n28 VSUBS 0.02827f
C1607 VP.n29 VSUBS 0.02827f
C1608 VP.n30 VSUBS 0.056186f
C1609 VP.n31 VSUBS 0.052688f
C1610 VP.n32 VSUBS 0.042283f
C1611 VP.n33 VSUBS 0.02827f
C1612 VP.n34 VSUBS 0.02827f
C1613 VP.n35 VSUBS 0.03708f
C1614 VP.n36 VSUBS 0.052688f
C1615 VP.n37 VSUBS 0.056634f
C1616 VP.n38 VSUBS 0.02827f
C1617 VP.n39 VSUBS 0.02827f
C1618 VP.n40 VSUBS 0.02827f
C1619 VP.n41 VSUBS 0.051885f
C1620 VP.n42 VSUBS 0.052688f
C1621 VP.n43 VSUBS 0.047485f
C1622 VP.n44 VSUBS 0.045627f
C1623 VP.n45 VSUBS 1.79773f
C1624 VP.n46 VSUBS 1.81648f
C1625 VP.n47 VSUBS 0.045627f
C1626 VP.n48 VSUBS 0.047485f
C1627 VP.n49 VSUBS 0.052688f
C1628 VP.n50 VSUBS 0.051885f
C1629 VP.n51 VSUBS 0.02827f
C1630 VP.n52 VSUBS 0.02827f
C1631 VP.n53 VSUBS 0.02827f
C1632 VP.n54 VSUBS 0.056634f
C1633 VP.n55 VSUBS 0.052688f
C1634 VP.n56 VSUBS 0.03708f
C1635 VP.n57 VSUBS 0.02827f
C1636 VP.n58 VSUBS 0.02827f
C1637 VP.n59 VSUBS 0.042283f
C1638 VP.n60 VSUBS 0.052688f
C1639 VP.n61 VSUBS 0.056186f
C1640 VP.n62 VSUBS 0.02827f
C1641 VP.n63 VSUBS 0.02827f
C1642 VP.n64 VSUBS 0.02827f
C1643 VP.n65 VSUBS 0.056186f
C1644 VP.n66 VSUBS 0.052688f
C1645 VP.n67 VSUBS 0.042283f
C1646 VP.n68 VSUBS 0.02827f
C1647 VP.n69 VSUBS 0.02827f
C1648 VP.n70 VSUBS 0.03708f
C1649 VP.n71 VSUBS 0.052688f
C1650 VP.n72 VSUBS 0.056634f
C1651 VP.n73 VSUBS 0.02827f
C1652 VP.n74 VSUBS 0.02827f
C1653 VP.n75 VSUBS 0.02827f
C1654 VP.n76 VSUBS 0.051885f
C1655 VP.n77 VSUBS 0.052688f
C1656 VP.n78 VSUBS 0.047485f
C1657 VP.n79 VSUBS 0.045627f
C1658 VP.n80 VSUBS 0.061936f
.ends

