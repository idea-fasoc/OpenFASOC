* NGSPICE file created from diff_pair_sample_1335.ext - technology: sky130A

.subckt diff_pair_sample_1335 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8541 pd=5.16 as=0.8541 ps=5.16 w=2.19 l=3.52
X1 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=0.8541 pd=5.16 as=0 ps=0 w=2.19 l=3.52
X2 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8541 pd=5.16 as=0.8541 ps=5.16 w=2.19 l=3.52
X3 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=0.8541 pd=5.16 as=0 ps=0 w=2.19 l=3.52
X4 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.8541 pd=5.16 as=0.8541 ps=5.16 w=2.19 l=3.52
X5 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.8541 pd=5.16 as=0 ps=0 w=2.19 l=3.52
X6 VDD1.t0 VP.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.8541 pd=5.16 as=0.8541 ps=5.16 w=2.19 l=3.52
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.8541 pd=5.16 as=0 ps=0 w=2.19 l=3.52
R0 VP.n0 VP.t0 93.4464
R1 VP.n0 VP.t1 53.7823
R2 VP VP.n0 0.52637
R3 VTAIL.n2 VTAIL.t2 86.0239
R4 VTAIL.n3 VTAIL.t1 86.0238
R5 VTAIL.n0 VTAIL.t3 86.0238
R6 VTAIL.n1 VTAIL.t0 86.0237
R7 VTAIL.n1 VTAIL.n0 20.8927
R8 VTAIL.n3 VTAIL.n2 17.5738
R9 VTAIL.n2 VTAIL.n1 2.12981
R10 VTAIL VTAIL.n0 1.35826
R11 VTAIL VTAIL.n3 0.772052
R12 VDD1 VDD1.t0 136.243
R13 VDD1 VDD1.t1 103.591
R14 B.n363 B.n81 585
R15 B.n81 B.n58 585
R16 B.n365 B.n364 585
R17 B.n367 B.n80 585
R18 B.n370 B.n369 585
R19 B.n371 B.n79 585
R20 B.n373 B.n372 585
R21 B.n375 B.n78 585
R22 B.n378 B.n377 585
R23 B.n379 B.n77 585
R24 B.n381 B.n380 585
R25 B.n383 B.n76 585
R26 B.n385 B.n384 585
R27 B.n387 B.n386 585
R28 B.n390 B.n389 585
R29 B.n391 B.n71 585
R30 B.n393 B.n392 585
R31 B.n395 B.n70 585
R32 B.n398 B.n397 585
R33 B.n399 B.n69 585
R34 B.n401 B.n400 585
R35 B.n403 B.n68 585
R36 B.n406 B.n405 585
R37 B.n408 B.n65 585
R38 B.n410 B.n409 585
R39 B.n412 B.n64 585
R40 B.n415 B.n414 585
R41 B.n416 B.n63 585
R42 B.n418 B.n417 585
R43 B.n420 B.n62 585
R44 B.n423 B.n422 585
R45 B.n424 B.n61 585
R46 B.n426 B.n425 585
R47 B.n428 B.n60 585
R48 B.n431 B.n430 585
R49 B.n432 B.n59 585
R50 B.n362 B.n57 585
R51 B.n435 B.n57 585
R52 B.n361 B.n56 585
R53 B.n436 B.n56 585
R54 B.n360 B.n55 585
R55 B.n437 B.n55 585
R56 B.n359 B.n358 585
R57 B.n358 B.n51 585
R58 B.n357 B.n50 585
R59 B.n443 B.n50 585
R60 B.n356 B.n49 585
R61 B.n444 B.n49 585
R62 B.n355 B.n48 585
R63 B.n445 B.n48 585
R64 B.n354 B.n353 585
R65 B.n353 B.n44 585
R66 B.n352 B.n43 585
R67 B.n451 B.n43 585
R68 B.n351 B.n42 585
R69 B.n452 B.n42 585
R70 B.n350 B.n41 585
R71 B.n453 B.n41 585
R72 B.n349 B.n348 585
R73 B.n348 B.n37 585
R74 B.n347 B.n36 585
R75 B.n459 B.n36 585
R76 B.n346 B.n35 585
R77 B.n460 B.n35 585
R78 B.n345 B.n34 585
R79 B.n461 B.n34 585
R80 B.n344 B.n343 585
R81 B.n343 B.n30 585
R82 B.n342 B.n29 585
R83 B.n467 B.n29 585
R84 B.n341 B.n28 585
R85 B.n468 B.n28 585
R86 B.n340 B.n27 585
R87 B.n469 B.n27 585
R88 B.n339 B.n338 585
R89 B.n338 B.n23 585
R90 B.n337 B.n22 585
R91 B.n475 B.n22 585
R92 B.n336 B.n21 585
R93 B.n476 B.n21 585
R94 B.n335 B.n20 585
R95 B.n477 B.n20 585
R96 B.n334 B.n333 585
R97 B.n333 B.n19 585
R98 B.n332 B.n15 585
R99 B.n483 B.n15 585
R100 B.n331 B.n14 585
R101 B.n484 B.n14 585
R102 B.n330 B.n13 585
R103 B.n485 B.n13 585
R104 B.n329 B.n328 585
R105 B.n328 B.n12 585
R106 B.n327 B.n326 585
R107 B.n327 B.n8 585
R108 B.n325 B.n7 585
R109 B.n492 B.n7 585
R110 B.n324 B.n6 585
R111 B.n493 B.n6 585
R112 B.n323 B.n5 585
R113 B.n494 B.n5 585
R114 B.n322 B.n321 585
R115 B.n321 B.n4 585
R116 B.n320 B.n82 585
R117 B.n320 B.n319 585
R118 B.n310 B.n83 585
R119 B.n84 B.n83 585
R120 B.n312 B.n311 585
R121 B.n313 B.n312 585
R122 B.n309 B.n89 585
R123 B.n89 B.n88 585
R124 B.n308 B.n307 585
R125 B.n307 B.n306 585
R126 B.n91 B.n90 585
R127 B.n299 B.n91 585
R128 B.n298 B.n297 585
R129 B.n300 B.n298 585
R130 B.n296 B.n96 585
R131 B.n96 B.n95 585
R132 B.n295 B.n294 585
R133 B.n294 B.n293 585
R134 B.n98 B.n97 585
R135 B.n99 B.n98 585
R136 B.n286 B.n285 585
R137 B.n287 B.n286 585
R138 B.n284 B.n104 585
R139 B.n104 B.n103 585
R140 B.n283 B.n282 585
R141 B.n282 B.n281 585
R142 B.n106 B.n105 585
R143 B.n107 B.n106 585
R144 B.n274 B.n273 585
R145 B.n275 B.n274 585
R146 B.n272 B.n112 585
R147 B.n112 B.n111 585
R148 B.n271 B.n270 585
R149 B.n270 B.n269 585
R150 B.n114 B.n113 585
R151 B.n115 B.n114 585
R152 B.n262 B.n261 585
R153 B.n263 B.n262 585
R154 B.n260 B.n120 585
R155 B.n120 B.n119 585
R156 B.n259 B.n258 585
R157 B.n258 B.n257 585
R158 B.n122 B.n121 585
R159 B.n123 B.n122 585
R160 B.n250 B.n249 585
R161 B.n251 B.n250 585
R162 B.n248 B.n128 585
R163 B.n128 B.n127 585
R164 B.n247 B.n246 585
R165 B.n246 B.n245 585
R166 B.n130 B.n129 585
R167 B.n131 B.n130 585
R168 B.n238 B.n237 585
R169 B.n239 B.n238 585
R170 B.n236 B.n136 585
R171 B.n136 B.n135 585
R172 B.n235 B.n234 585
R173 B.n234 B.n233 585
R174 B.n230 B.n140 585
R175 B.n229 B.n228 585
R176 B.n226 B.n141 585
R177 B.n226 B.n139 585
R178 B.n225 B.n224 585
R179 B.n223 B.n222 585
R180 B.n221 B.n143 585
R181 B.n219 B.n218 585
R182 B.n217 B.n144 585
R183 B.n216 B.n215 585
R184 B.n213 B.n145 585
R185 B.n211 B.n210 585
R186 B.n209 B.n146 585
R187 B.n208 B.n207 585
R188 B.n205 B.n204 585
R189 B.n203 B.n202 585
R190 B.n201 B.n151 585
R191 B.n199 B.n198 585
R192 B.n197 B.n152 585
R193 B.n196 B.n195 585
R194 B.n193 B.n153 585
R195 B.n191 B.n190 585
R196 B.n189 B.n154 585
R197 B.n187 B.n186 585
R198 B.n184 B.n157 585
R199 B.n182 B.n181 585
R200 B.n180 B.n158 585
R201 B.n179 B.n178 585
R202 B.n176 B.n159 585
R203 B.n174 B.n173 585
R204 B.n172 B.n160 585
R205 B.n171 B.n170 585
R206 B.n168 B.n161 585
R207 B.n166 B.n165 585
R208 B.n164 B.n163 585
R209 B.n138 B.n137 585
R210 B.n232 B.n231 585
R211 B.n233 B.n232 585
R212 B.n134 B.n133 585
R213 B.n135 B.n134 585
R214 B.n241 B.n240 585
R215 B.n240 B.n239 585
R216 B.n242 B.n132 585
R217 B.n132 B.n131 585
R218 B.n244 B.n243 585
R219 B.n245 B.n244 585
R220 B.n126 B.n125 585
R221 B.n127 B.n126 585
R222 B.n253 B.n252 585
R223 B.n252 B.n251 585
R224 B.n254 B.n124 585
R225 B.n124 B.n123 585
R226 B.n256 B.n255 585
R227 B.n257 B.n256 585
R228 B.n118 B.n117 585
R229 B.n119 B.n118 585
R230 B.n265 B.n264 585
R231 B.n264 B.n263 585
R232 B.n266 B.n116 585
R233 B.n116 B.n115 585
R234 B.n268 B.n267 585
R235 B.n269 B.n268 585
R236 B.n110 B.n109 585
R237 B.n111 B.n110 585
R238 B.n277 B.n276 585
R239 B.n276 B.n275 585
R240 B.n278 B.n108 585
R241 B.n108 B.n107 585
R242 B.n280 B.n279 585
R243 B.n281 B.n280 585
R244 B.n102 B.n101 585
R245 B.n103 B.n102 585
R246 B.n289 B.n288 585
R247 B.n288 B.n287 585
R248 B.n290 B.n100 585
R249 B.n100 B.n99 585
R250 B.n292 B.n291 585
R251 B.n293 B.n292 585
R252 B.n94 B.n93 585
R253 B.n95 B.n94 585
R254 B.n302 B.n301 585
R255 B.n301 B.n300 585
R256 B.n303 B.n92 585
R257 B.n299 B.n92 585
R258 B.n305 B.n304 585
R259 B.n306 B.n305 585
R260 B.n87 B.n86 585
R261 B.n88 B.n87 585
R262 B.n315 B.n314 585
R263 B.n314 B.n313 585
R264 B.n316 B.n85 585
R265 B.n85 B.n84 585
R266 B.n318 B.n317 585
R267 B.n319 B.n318 585
R268 B.n3 B.n0 585
R269 B.n4 B.n3 585
R270 B.n491 B.n1 585
R271 B.n492 B.n491 585
R272 B.n490 B.n489 585
R273 B.n490 B.n8 585
R274 B.n488 B.n9 585
R275 B.n12 B.n9 585
R276 B.n487 B.n486 585
R277 B.n486 B.n485 585
R278 B.n11 B.n10 585
R279 B.n484 B.n11 585
R280 B.n482 B.n481 585
R281 B.n483 B.n482 585
R282 B.n480 B.n16 585
R283 B.n19 B.n16 585
R284 B.n479 B.n478 585
R285 B.n478 B.n477 585
R286 B.n18 B.n17 585
R287 B.n476 B.n18 585
R288 B.n474 B.n473 585
R289 B.n475 B.n474 585
R290 B.n472 B.n24 585
R291 B.n24 B.n23 585
R292 B.n471 B.n470 585
R293 B.n470 B.n469 585
R294 B.n26 B.n25 585
R295 B.n468 B.n26 585
R296 B.n466 B.n465 585
R297 B.n467 B.n466 585
R298 B.n464 B.n31 585
R299 B.n31 B.n30 585
R300 B.n463 B.n462 585
R301 B.n462 B.n461 585
R302 B.n33 B.n32 585
R303 B.n460 B.n33 585
R304 B.n458 B.n457 585
R305 B.n459 B.n458 585
R306 B.n456 B.n38 585
R307 B.n38 B.n37 585
R308 B.n455 B.n454 585
R309 B.n454 B.n453 585
R310 B.n40 B.n39 585
R311 B.n452 B.n40 585
R312 B.n450 B.n449 585
R313 B.n451 B.n450 585
R314 B.n448 B.n45 585
R315 B.n45 B.n44 585
R316 B.n447 B.n446 585
R317 B.n446 B.n445 585
R318 B.n47 B.n46 585
R319 B.n444 B.n47 585
R320 B.n442 B.n441 585
R321 B.n443 B.n442 585
R322 B.n440 B.n52 585
R323 B.n52 B.n51 585
R324 B.n439 B.n438 585
R325 B.n438 B.n437 585
R326 B.n54 B.n53 585
R327 B.n436 B.n54 585
R328 B.n434 B.n433 585
R329 B.n435 B.n434 585
R330 B.n495 B.n494 585
R331 B.n493 B.n2 585
R332 B.n434 B.n59 550.159
R333 B.n81 B.n57 550.159
R334 B.n234 B.n138 550.159
R335 B.n232 B.n140 550.159
R336 B.n366 B.n58 256.663
R337 B.n368 B.n58 256.663
R338 B.n374 B.n58 256.663
R339 B.n376 B.n58 256.663
R340 B.n382 B.n58 256.663
R341 B.n75 B.n58 256.663
R342 B.n388 B.n58 256.663
R343 B.n394 B.n58 256.663
R344 B.n396 B.n58 256.663
R345 B.n402 B.n58 256.663
R346 B.n404 B.n58 256.663
R347 B.n411 B.n58 256.663
R348 B.n413 B.n58 256.663
R349 B.n419 B.n58 256.663
R350 B.n421 B.n58 256.663
R351 B.n427 B.n58 256.663
R352 B.n429 B.n58 256.663
R353 B.n227 B.n139 256.663
R354 B.n142 B.n139 256.663
R355 B.n220 B.n139 256.663
R356 B.n214 B.n139 256.663
R357 B.n212 B.n139 256.663
R358 B.n206 B.n139 256.663
R359 B.n150 B.n139 256.663
R360 B.n200 B.n139 256.663
R361 B.n194 B.n139 256.663
R362 B.n192 B.n139 256.663
R363 B.n185 B.n139 256.663
R364 B.n183 B.n139 256.663
R365 B.n177 B.n139 256.663
R366 B.n175 B.n139 256.663
R367 B.n169 B.n139 256.663
R368 B.n167 B.n139 256.663
R369 B.n162 B.n139 256.663
R370 B.n497 B.n496 256.663
R371 B.n66 B.t2 224.106
R372 B.n72 B.t6 224.106
R373 B.n155 B.t13 224.106
R374 B.n147 B.t9 224.106
R375 B.n233 B.n139 207.77
R376 B.n435 B.n58 207.77
R377 B.n430 B.n428 163.367
R378 B.n426 B.n61 163.367
R379 B.n422 B.n420 163.367
R380 B.n418 B.n63 163.367
R381 B.n414 B.n412 163.367
R382 B.n410 B.n65 163.367
R383 B.n405 B.n403 163.367
R384 B.n401 B.n69 163.367
R385 B.n397 B.n395 163.367
R386 B.n393 B.n71 163.367
R387 B.n389 B.n387 163.367
R388 B.n384 B.n383 163.367
R389 B.n381 B.n77 163.367
R390 B.n377 B.n375 163.367
R391 B.n373 B.n79 163.367
R392 B.n369 B.n367 163.367
R393 B.n365 B.n81 163.367
R394 B.n234 B.n136 163.367
R395 B.n238 B.n136 163.367
R396 B.n238 B.n130 163.367
R397 B.n246 B.n130 163.367
R398 B.n246 B.n128 163.367
R399 B.n250 B.n128 163.367
R400 B.n250 B.n122 163.367
R401 B.n258 B.n122 163.367
R402 B.n258 B.n120 163.367
R403 B.n262 B.n120 163.367
R404 B.n262 B.n114 163.367
R405 B.n270 B.n114 163.367
R406 B.n270 B.n112 163.367
R407 B.n274 B.n112 163.367
R408 B.n274 B.n106 163.367
R409 B.n282 B.n106 163.367
R410 B.n282 B.n104 163.367
R411 B.n286 B.n104 163.367
R412 B.n286 B.n98 163.367
R413 B.n294 B.n98 163.367
R414 B.n294 B.n96 163.367
R415 B.n298 B.n96 163.367
R416 B.n298 B.n91 163.367
R417 B.n307 B.n91 163.367
R418 B.n307 B.n89 163.367
R419 B.n312 B.n89 163.367
R420 B.n312 B.n83 163.367
R421 B.n320 B.n83 163.367
R422 B.n321 B.n320 163.367
R423 B.n321 B.n5 163.367
R424 B.n6 B.n5 163.367
R425 B.n7 B.n6 163.367
R426 B.n327 B.n7 163.367
R427 B.n328 B.n327 163.367
R428 B.n328 B.n13 163.367
R429 B.n14 B.n13 163.367
R430 B.n15 B.n14 163.367
R431 B.n333 B.n15 163.367
R432 B.n333 B.n20 163.367
R433 B.n21 B.n20 163.367
R434 B.n22 B.n21 163.367
R435 B.n338 B.n22 163.367
R436 B.n338 B.n27 163.367
R437 B.n28 B.n27 163.367
R438 B.n29 B.n28 163.367
R439 B.n343 B.n29 163.367
R440 B.n343 B.n34 163.367
R441 B.n35 B.n34 163.367
R442 B.n36 B.n35 163.367
R443 B.n348 B.n36 163.367
R444 B.n348 B.n41 163.367
R445 B.n42 B.n41 163.367
R446 B.n43 B.n42 163.367
R447 B.n353 B.n43 163.367
R448 B.n353 B.n48 163.367
R449 B.n49 B.n48 163.367
R450 B.n50 B.n49 163.367
R451 B.n358 B.n50 163.367
R452 B.n358 B.n55 163.367
R453 B.n56 B.n55 163.367
R454 B.n57 B.n56 163.367
R455 B.n228 B.n226 163.367
R456 B.n226 B.n225 163.367
R457 B.n222 B.n221 163.367
R458 B.n219 B.n144 163.367
R459 B.n215 B.n213 163.367
R460 B.n211 B.n146 163.367
R461 B.n207 B.n205 163.367
R462 B.n202 B.n201 163.367
R463 B.n199 B.n152 163.367
R464 B.n195 B.n193 163.367
R465 B.n191 B.n154 163.367
R466 B.n186 B.n184 163.367
R467 B.n182 B.n158 163.367
R468 B.n178 B.n176 163.367
R469 B.n174 B.n160 163.367
R470 B.n170 B.n168 163.367
R471 B.n166 B.n163 163.367
R472 B.n232 B.n134 163.367
R473 B.n240 B.n134 163.367
R474 B.n240 B.n132 163.367
R475 B.n244 B.n132 163.367
R476 B.n244 B.n126 163.367
R477 B.n252 B.n126 163.367
R478 B.n252 B.n124 163.367
R479 B.n256 B.n124 163.367
R480 B.n256 B.n118 163.367
R481 B.n264 B.n118 163.367
R482 B.n264 B.n116 163.367
R483 B.n268 B.n116 163.367
R484 B.n268 B.n110 163.367
R485 B.n276 B.n110 163.367
R486 B.n276 B.n108 163.367
R487 B.n280 B.n108 163.367
R488 B.n280 B.n102 163.367
R489 B.n288 B.n102 163.367
R490 B.n288 B.n100 163.367
R491 B.n292 B.n100 163.367
R492 B.n292 B.n94 163.367
R493 B.n301 B.n94 163.367
R494 B.n301 B.n92 163.367
R495 B.n305 B.n92 163.367
R496 B.n305 B.n87 163.367
R497 B.n314 B.n87 163.367
R498 B.n314 B.n85 163.367
R499 B.n318 B.n85 163.367
R500 B.n318 B.n3 163.367
R501 B.n495 B.n3 163.367
R502 B.n491 B.n2 163.367
R503 B.n491 B.n490 163.367
R504 B.n490 B.n9 163.367
R505 B.n486 B.n9 163.367
R506 B.n486 B.n11 163.367
R507 B.n482 B.n11 163.367
R508 B.n482 B.n16 163.367
R509 B.n478 B.n16 163.367
R510 B.n478 B.n18 163.367
R511 B.n474 B.n18 163.367
R512 B.n474 B.n24 163.367
R513 B.n470 B.n24 163.367
R514 B.n470 B.n26 163.367
R515 B.n466 B.n26 163.367
R516 B.n466 B.n31 163.367
R517 B.n462 B.n31 163.367
R518 B.n462 B.n33 163.367
R519 B.n458 B.n33 163.367
R520 B.n458 B.n38 163.367
R521 B.n454 B.n38 163.367
R522 B.n454 B.n40 163.367
R523 B.n450 B.n40 163.367
R524 B.n450 B.n45 163.367
R525 B.n446 B.n45 163.367
R526 B.n446 B.n47 163.367
R527 B.n442 B.n47 163.367
R528 B.n442 B.n52 163.367
R529 B.n438 B.n52 163.367
R530 B.n438 B.n54 163.367
R531 B.n434 B.n54 163.367
R532 B.n72 B.t7 160.221
R533 B.n155 B.t15 160.221
R534 B.n66 B.t4 160.221
R535 B.n147 B.t12 160.221
R536 B.n233 B.n135 100.201
R537 B.n239 B.n135 100.201
R538 B.n239 B.n131 100.201
R539 B.n245 B.n131 100.201
R540 B.n245 B.n127 100.201
R541 B.n251 B.n127 100.201
R542 B.n251 B.n123 100.201
R543 B.n257 B.n123 100.201
R544 B.n263 B.n119 100.201
R545 B.n263 B.n115 100.201
R546 B.n269 B.n115 100.201
R547 B.n269 B.n111 100.201
R548 B.n275 B.n111 100.201
R549 B.n275 B.n107 100.201
R550 B.n281 B.n107 100.201
R551 B.n281 B.n103 100.201
R552 B.n287 B.n103 100.201
R553 B.n287 B.n99 100.201
R554 B.n293 B.n99 100.201
R555 B.n293 B.n95 100.201
R556 B.n300 B.n95 100.201
R557 B.n300 B.n299 100.201
R558 B.n306 B.n88 100.201
R559 B.n313 B.n88 100.201
R560 B.n313 B.n84 100.201
R561 B.n319 B.n84 100.201
R562 B.n319 B.n4 100.201
R563 B.n494 B.n4 100.201
R564 B.n494 B.n493 100.201
R565 B.n493 B.n492 100.201
R566 B.n492 B.n8 100.201
R567 B.n12 B.n8 100.201
R568 B.n485 B.n12 100.201
R569 B.n485 B.n484 100.201
R570 B.n484 B.n483 100.201
R571 B.n477 B.n19 100.201
R572 B.n477 B.n476 100.201
R573 B.n476 B.n475 100.201
R574 B.n475 B.n23 100.201
R575 B.n469 B.n23 100.201
R576 B.n469 B.n468 100.201
R577 B.n468 B.n467 100.201
R578 B.n467 B.n30 100.201
R579 B.n461 B.n30 100.201
R580 B.n461 B.n460 100.201
R581 B.n460 B.n459 100.201
R582 B.n459 B.n37 100.201
R583 B.n453 B.n37 100.201
R584 B.n453 B.n452 100.201
R585 B.n451 B.n44 100.201
R586 B.n445 B.n44 100.201
R587 B.n445 B.n444 100.201
R588 B.n444 B.n443 100.201
R589 B.n443 B.n51 100.201
R590 B.n437 B.n51 100.201
R591 B.n437 B.n436 100.201
R592 B.n436 B.n435 100.201
R593 B.n73 B.t8 85.5549
R594 B.n156 B.t14 85.5549
R595 B.n67 B.t5 85.5546
R596 B.n148 B.t11 85.5546
R597 B.n306 B.t0 76.6248
R598 B.n483 B.t1 76.6248
R599 B.n67 B.n66 74.6672
R600 B.n73 B.n72 74.6672
R601 B.n156 B.n155 74.6672
R602 B.n148 B.n147 74.6672
R603 B.n429 B.n59 71.676
R604 B.n428 B.n427 71.676
R605 B.n421 B.n61 71.676
R606 B.n420 B.n419 71.676
R607 B.n413 B.n63 71.676
R608 B.n412 B.n411 71.676
R609 B.n404 B.n65 71.676
R610 B.n403 B.n402 71.676
R611 B.n396 B.n69 71.676
R612 B.n395 B.n394 71.676
R613 B.n388 B.n71 71.676
R614 B.n387 B.n75 71.676
R615 B.n383 B.n382 71.676
R616 B.n376 B.n77 71.676
R617 B.n375 B.n374 71.676
R618 B.n368 B.n79 71.676
R619 B.n367 B.n366 71.676
R620 B.n366 B.n365 71.676
R621 B.n369 B.n368 71.676
R622 B.n374 B.n373 71.676
R623 B.n377 B.n376 71.676
R624 B.n382 B.n381 71.676
R625 B.n384 B.n75 71.676
R626 B.n389 B.n388 71.676
R627 B.n394 B.n393 71.676
R628 B.n397 B.n396 71.676
R629 B.n402 B.n401 71.676
R630 B.n405 B.n404 71.676
R631 B.n411 B.n410 71.676
R632 B.n414 B.n413 71.676
R633 B.n419 B.n418 71.676
R634 B.n422 B.n421 71.676
R635 B.n427 B.n426 71.676
R636 B.n430 B.n429 71.676
R637 B.n227 B.n140 71.676
R638 B.n225 B.n142 71.676
R639 B.n221 B.n220 71.676
R640 B.n214 B.n144 71.676
R641 B.n213 B.n212 71.676
R642 B.n206 B.n146 71.676
R643 B.n205 B.n150 71.676
R644 B.n201 B.n200 71.676
R645 B.n194 B.n152 71.676
R646 B.n193 B.n192 71.676
R647 B.n185 B.n154 71.676
R648 B.n184 B.n183 71.676
R649 B.n177 B.n158 71.676
R650 B.n176 B.n175 71.676
R651 B.n169 B.n160 71.676
R652 B.n168 B.n167 71.676
R653 B.n163 B.n162 71.676
R654 B.n228 B.n227 71.676
R655 B.n222 B.n142 71.676
R656 B.n220 B.n219 71.676
R657 B.n215 B.n214 71.676
R658 B.n212 B.n211 71.676
R659 B.n207 B.n206 71.676
R660 B.n202 B.n150 71.676
R661 B.n200 B.n199 71.676
R662 B.n195 B.n194 71.676
R663 B.n192 B.n191 71.676
R664 B.n186 B.n185 71.676
R665 B.n183 B.n182 71.676
R666 B.n178 B.n177 71.676
R667 B.n175 B.n174 71.676
R668 B.n170 B.n169 71.676
R669 B.n167 B.n166 71.676
R670 B.n162 B.n138 71.676
R671 B.n496 B.n495 71.676
R672 B.n496 B.n2 71.676
R673 B.n257 B.t10 70.7306
R674 B.t3 B.n451 70.7306
R675 B.n407 B.n67 59.5399
R676 B.n74 B.n73 59.5399
R677 B.n188 B.n156 59.5399
R678 B.n149 B.n148 59.5399
R679 B.n363 B.n362 35.7468
R680 B.n231 B.n230 35.7468
R681 B.n235 B.n137 35.7468
R682 B.n433 B.n432 35.7468
R683 B.t10 B.n119 29.4714
R684 B.n452 B.t3 29.4714
R685 B.n299 B.t0 23.5772
R686 B.n19 B.t1 23.5772
R687 B B.n497 18.0485
R688 B.n231 B.n133 10.6151
R689 B.n241 B.n133 10.6151
R690 B.n242 B.n241 10.6151
R691 B.n243 B.n242 10.6151
R692 B.n243 B.n125 10.6151
R693 B.n253 B.n125 10.6151
R694 B.n254 B.n253 10.6151
R695 B.n255 B.n254 10.6151
R696 B.n255 B.n117 10.6151
R697 B.n265 B.n117 10.6151
R698 B.n266 B.n265 10.6151
R699 B.n267 B.n266 10.6151
R700 B.n267 B.n109 10.6151
R701 B.n277 B.n109 10.6151
R702 B.n278 B.n277 10.6151
R703 B.n279 B.n278 10.6151
R704 B.n279 B.n101 10.6151
R705 B.n289 B.n101 10.6151
R706 B.n290 B.n289 10.6151
R707 B.n291 B.n290 10.6151
R708 B.n291 B.n93 10.6151
R709 B.n302 B.n93 10.6151
R710 B.n303 B.n302 10.6151
R711 B.n304 B.n303 10.6151
R712 B.n304 B.n86 10.6151
R713 B.n315 B.n86 10.6151
R714 B.n316 B.n315 10.6151
R715 B.n317 B.n316 10.6151
R716 B.n317 B.n0 10.6151
R717 B.n230 B.n229 10.6151
R718 B.n229 B.n141 10.6151
R719 B.n224 B.n141 10.6151
R720 B.n224 B.n223 10.6151
R721 B.n223 B.n143 10.6151
R722 B.n218 B.n143 10.6151
R723 B.n218 B.n217 10.6151
R724 B.n217 B.n216 10.6151
R725 B.n216 B.n145 10.6151
R726 B.n210 B.n145 10.6151
R727 B.n210 B.n209 10.6151
R728 B.n209 B.n208 10.6151
R729 B.n204 B.n203 10.6151
R730 B.n203 B.n151 10.6151
R731 B.n198 B.n151 10.6151
R732 B.n198 B.n197 10.6151
R733 B.n197 B.n196 10.6151
R734 B.n196 B.n153 10.6151
R735 B.n190 B.n153 10.6151
R736 B.n190 B.n189 10.6151
R737 B.n187 B.n157 10.6151
R738 B.n181 B.n157 10.6151
R739 B.n181 B.n180 10.6151
R740 B.n180 B.n179 10.6151
R741 B.n179 B.n159 10.6151
R742 B.n173 B.n159 10.6151
R743 B.n173 B.n172 10.6151
R744 B.n172 B.n171 10.6151
R745 B.n171 B.n161 10.6151
R746 B.n165 B.n161 10.6151
R747 B.n165 B.n164 10.6151
R748 B.n164 B.n137 10.6151
R749 B.n236 B.n235 10.6151
R750 B.n237 B.n236 10.6151
R751 B.n237 B.n129 10.6151
R752 B.n247 B.n129 10.6151
R753 B.n248 B.n247 10.6151
R754 B.n249 B.n248 10.6151
R755 B.n249 B.n121 10.6151
R756 B.n259 B.n121 10.6151
R757 B.n260 B.n259 10.6151
R758 B.n261 B.n260 10.6151
R759 B.n261 B.n113 10.6151
R760 B.n271 B.n113 10.6151
R761 B.n272 B.n271 10.6151
R762 B.n273 B.n272 10.6151
R763 B.n273 B.n105 10.6151
R764 B.n283 B.n105 10.6151
R765 B.n284 B.n283 10.6151
R766 B.n285 B.n284 10.6151
R767 B.n285 B.n97 10.6151
R768 B.n295 B.n97 10.6151
R769 B.n296 B.n295 10.6151
R770 B.n297 B.n296 10.6151
R771 B.n297 B.n90 10.6151
R772 B.n308 B.n90 10.6151
R773 B.n309 B.n308 10.6151
R774 B.n311 B.n309 10.6151
R775 B.n311 B.n310 10.6151
R776 B.n310 B.n82 10.6151
R777 B.n322 B.n82 10.6151
R778 B.n323 B.n322 10.6151
R779 B.n324 B.n323 10.6151
R780 B.n325 B.n324 10.6151
R781 B.n326 B.n325 10.6151
R782 B.n329 B.n326 10.6151
R783 B.n330 B.n329 10.6151
R784 B.n331 B.n330 10.6151
R785 B.n332 B.n331 10.6151
R786 B.n334 B.n332 10.6151
R787 B.n335 B.n334 10.6151
R788 B.n336 B.n335 10.6151
R789 B.n337 B.n336 10.6151
R790 B.n339 B.n337 10.6151
R791 B.n340 B.n339 10.6151
R792 B.n341 B.n340 10.6151
R793 B.n342 B.n341 10.6151
R794 B.n344 B.n342 10.6151
R795 B.n345 B.n344 10.6151
R796 B.n346 B.n345 10.6151
R797 B.n347 B.n346 10.6151
R798 B.n349 B.n347 10.6151
R799 B.n350 B.n349 10.6151
R800 B.n351 B.n350 10.6151
R801 B.n352 B.n351 10.6151
R802 B.n354 B.n352 10.6151
R803 B.n355 B.n354 10.6151
R804 B.n356 B.n355 10.6151
R805 B.n357 B.n356 10.6151
R806 B.n359 B.n357 10.6151
R807 B.n360 B.n359 10.6151
R808 B.n361 B.n360 10.6151
R809 B.n362 B.n361 10.6151
R810 B.n489 B.n1 10.6151
R811 B.n489 B.n488 10.6151
R812 B.n488 B.n487 10.6151
R813 B.n487 B.n10 10.6151
R814 B.n481 B.n10 10.6151
R815 B.n481 B.n480 10.6151
R816 B.n480 B.n479 10.6151
R817 B.n479 B.n17 10.6151
R818 B.n473 B.n17 10.6151
R819 B.n473 B.n472 10.6151
R820 B.n472 B.n471 10.6151
R821 B.n471 B.n25 10.6151
R822 B.n465 B.n25 10.6151
R823 B.n465 B.n464 10.6151
R824 B.n464 B.n463 10.6151
R825 B.n463 B.n32 10.6151
R826 B.n457 B.n32 10.6151
R827 B.n457 B.n456 10.6151
R828 B.n456 B.n455 10.6151
R829 B.n455 B.n39 10.6151
R830 B.n449 B.n39 10.6151
R831 B.n449 B.n448 10.6151
R832 B.n448 B.n447 10.6151
R833 B.n447 B.n46 10.6151
R834 B.n441 B.n46 10.6151
R835 B.n441 B.n440 10.6151
R836 B.n440 B.n439 10.6151
R837 B.n439 B.n53 10.6151
R838 B.n433 B.n53 10.6151
R839 B.n432 B.n431 10.6151
R840 B.n431 B.n60 10.6151
R841 B.n425 B.n60 10.6151
R842 B.n425 B.n424 10.6151
R843 B.n424 B.n423 10.6151
R844 B.n423 B.n62 10.6151
R845 B.n417 B.n62 10.6151
R846 B.n417 B.n416 10.6151
R847 B.n416 B.n415 10.6151
R848 B.n415 B.n64 10.6151
R849 B.n409 B.n64 10.6151
R850 B.n409 B.n408 10.6151
R851 B.n406 B.n68 10.6151
R852 B.n400 B.n68 10.6151
R853 B.n400 B.n399 10.6151
R854 B.n399 B.n398 10.6151
R855 B.n398 B.n70 10.6151
R856 B.n392 B.n70 10.6151
R857 B.n392 B.n391 10.6151
R858 B.n391 B.n390 10.6151
R859 B.n386 B.n385 10.6151
R860 B.n385 B.n76 10.6151
R861 B.n380 B.n76 10.6151
R862 B.n380 B.n379 10.6151
R863 B.n379 B.n378 10.6151
R864 B.n378 B.n78 10.6151
R865 B.n372 B.n78 10.6151
R866 B.n372 B.n371 10.6151
R867 B.n371 B.n370 10.6151
R868 B.n370 B.n80 10.6151
R869 B.n364 B.n80 10.6151
R870 B.n364 B.n363 10.6151
R871 B.n497 B.n0 8.11757
R872 B.n497 B.n1 8.11757
R873 B.n204 B.n149 6.5566
R874 B.n189 B.n188 6.5566
R875 B.n407 B.n406 6.5566
R876 B.n390 B.n74 6.5566
R877 B.n208 B.n149 4.05904
R878 B.n188 B.n187 4.05904
R879 B.n408 B.n407 4.05904
R880 B.n386 B.n74 4.05904
R881 VN VN.t1 93.3536
R882 VN VN.t0 54.3081
R883 VDD2.n0 VDD2.t1 134.887
R884 VDD2.n0 VDD2.t0 102.703
R885 VDD2 VDD2.n0 0.888431
C0 VP VDD1 0.963648f
C1 VP VDD2 0.377891f
C2 VP VTAIL 1.1438f
C3 VDD1 VDD2 0.774293f
C4 VDD1 VTAIL 2.77442f
C5 VTAIL VDD2 2.83364f
C6 VN VP 4.07631f
C7 VN VDD1 0.154582f
C8 VN VDD2 0.742014f
C9 VN VTAIL 1.12968f
C10 VDD2 B 2.970265f
C11 VDD1 B 5.09606f
C12 VTAIL B 3.36985f
C13 VN B 8.74273f
C14 VP B 6.63784f
C15 VDD2.t1 B 0.479588f
C16 VDD2.t0 B 0.270959f
C17 VDD2.n0 B 1.90259f
C18 VN.t0 B 0.761205f
C19 VN.t1 B 1.29538f
C20 VDD1.t1 B 0.266494f
C21 VDD1.t0 B 0.490186f
C22 VTAIL.t3 B 0.292691f
C23 VTAIL.n0 B 1.16899f
C24 VTAIL.t0 B 0.292693f
C25 VTAIL.n1 B 1.22258f
C26 VTAIL.t2 B 0.292691f
C27 VTAIL.n2 B 0.992035f
C28 VTAIL.t1 B 0.292691f
C29 VTAIL.n3 B 0.89772f
C30 VP.t0 B 1.30554f
C31 VP.t1 B 0.765018f
C32 VP.n0 B 1.93346f
.ends

