* NGSPICE file created from diff_pair_sample_0560.ext - technology: sky130A

.subckt diff_pair_sample_0560 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t17 VN.t0 VDD2.t8 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=1.50645 pd=9.46 as=1.50645 ps=9.46 w=9.13 l=0.29
X1 VDD1.t9 VP.t0 VTAIL.t4 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=1.50645 pd=9.46 as=3.5607 ps=19.04 w=9.13 l=0.29
X2 VDD2.t7 VN.t1 VTAIL.t16 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=1.50645 pd=9.46 as=1.50645 ps=9.46 w=9.13 l=0.29
X3 VTAIL.t15 VN.t2 VDD2.t6 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=1.50645 pd=9.46 as=1.50645 ps=9.46 w=9.13 l=0.29
X4 VDD1.t8 VP.t1 VTAIL.t5 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=1.50645 pd=9.46 as=1.50645 ps=9.46 w=9.13 l=0.29
X5 VDD2.t0 VN.t3 VTAIL.t14 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=1.50645 pd=9.46 as=1.50645 ps=9.46 w=9.13 l=0.29
X6 VTAIL.t18 VP.t2 VDD1.t7 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=1.50645 pd=9.46 as=1.50645 ps=9.46 w=9.13 l=0.29
X7 VDD1.t6 VP.t3 VTAIL.t7 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=1.50645 pd=9.46 as=3.5607 ps=19.04 w=9.13 l=0.29
X8 VDD2.t9 VN.t4 VTAIL.t13 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=3.5607 pd=19.04 as=1.50645 ps=9.46 w=9.13 l=0.29
X9 VTAIL.t12 VN.t5 VDD2.t2 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=1.50645 pd=9.46 as=1.50645 ps=9.46 w=9.13 l=0.29
X10 VTAIL.t1 VP.t4 VDD1.t5 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=1.50645 pd=9.46 as=1.50645 ps=9.46 w=9.13 l=0.29
X11 VTAIL.t11 VN.t6 VDD2.t3 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=1.50645 pd=9.46 as=1.50645 ps=9.46 w=9.13 l=0.29
X12 VDD2.t4 VN.t7 VTAIL.t10 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=1.50645 pd=9.46 as=3.5607 ps=19.04 w=9.13 l=0.29
X13 VDD2.t1 VN.t8 VTAIL.t9 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=1.50645 pd=9.46 as=3.5607 ps=19.04 w=9.13 l=0.29
X14 VDD1.t4 VP.t5 VTAIL.t19 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=1.50645 pd=9.46 as=1.50645 ps=9.46 w=9.13 l=0.29
X15 VDD1.t3 VP.t6 VTAIL.t6 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=3.5607 pd=19.04 as=1.50645 ps=9.46 w=9.13 l=0.29
X16 VTAIL.t0 VP.t7 VDD1.t2 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=1.50645 pd=9.46 as=1.50645 ps=9.46 w=9.13 l=0.29
X17 B.t11 B.t9 B.t10 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=3.5607 pd=19.04 as=0 ps=0 w=9.13 l=0.29
X18 VDD2.t5 VN.t9 VTAIL.t8 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=3.5607 pd=19.04 as=1.50645 ps=9.46 w=9.13 l=0.29
X19 VTAIL.t2 VP.t8 VDD1.t1 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=1.50645 pd=9.46 as=1.50645 ps=9.46 w=9.13 l=0.29
X20 B.t8 B.t6 B.t7 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=3.5607 pd=19.04 as=0 ps=0 w=9.13 l=0.29
X21 B.t5 B.t3 B.t4 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=3.5607 pd=19.04 as=0 ps=0 w=9.13 l=0.29
X22 B.t2 B.t0 B.t1 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=3.5607 pd=19.04 as=0 ps=0 w=9.13 l=0.29
X23 VDD1.t0 VP.t9 VTAIL.t3 w_n1714_n2794# sky130_fd_pr__pfet_01v8 ad=3.5607 pd=19.04 as=1.50645 ps=9.46 w=9.13 l=0.29
R0 VN.n9 VN.t8 902.655
R1 VN.n3 VN.t9 902.655
R2 VN.n20 VN.t4 902.655
R3 VN.n14 VN.t7 902.655
R4 VN.n6 VN.t3 867.601
R5 VN.n8 VN.t2 867.601
R6 VN.n2 VN.t0 867.601
R7 VN.n17 VN.t1 867.601
R8 VN.n19 VN.t6 867.601
R9 VN.n13 VN.t5 867.601
R10 VN.n15 VN.n14 161.489
R11 VN.n4 VN.n3 161.489
R12 VN.n10 VN.n9 161.3
R13 VN.n21 VN.n20 161.3
R14 VN.n18 VN.n11 161.3
R15 VN.n17 VN.n16 161.3
R16 VN.n15 VN.n12 161.3
R17 VN.n7 VN.n0 161.3
R18 VN.n6 VN.n5 161.3
R19 VN.n4 VN.n1 161.3
R20 VN.n6 VN.n1 73.0308
R21 VN.n7 VN.n6 73.0308
R22 VN.n18 VN.n17 73.0308
R23 VN.n17 VN.n12 73.0308
R24 VN.n3 VN.n2 55.5035
R25 VN.n9 VN.n8 55.5035
R26 VN.n20 VN.n19 55.5035
R27 VN.n14 VN.n13 55.5035
R28 VN VN.n21 38.7978
R29 VN.n2 VN.n1 17.5278
R30 VN.n8 VN.n7 17.5278
R31 VN.n19 VN.n18 17.5278
R32 VN.n13 VN.n12 17.5278
R33 VN.n21 VN.n11 0.189894
R34 VN.n16 VN.n11 0.189894
R35 VN.n16 VN.n15 0.189894
R36 VN.n5 VN.n4 0.189894
R37 VN.n5 VN.n0 0.189894
R38 VN.n10 VN.n0 0.189894
R39 VN VN.n10 0.0516364
R40 VDD2.n1 VDD2.t5 81.7584
R41 VDD2.n4 VDD2.t9 81.2241
R42 VDD2.n3 VDD2.n2 78.0092
R43 VDD2 VDD2.n7 78.0065
R44 VDD2.n6 VDD2.n5 77.6639
R45 VDD2.n1 VDD2.n0 77.6636
R46 VDD2.n4 VDD2.n3 34.1248
R47 VDD2.n7 VDD2.t2 3.56074
R48 VDD2.n7 VDD2.t4 3.56074
R49 VDD2.n5 VDD2.t3 3.56074
R50 VDD2.n5 VDD2.t7 3.56074
R51 VDD2.n2 VDD2.t6 3.56074
R52 VDD2.n2 VDD2.t1 3.56074
R53 VDD2.n0 VDD2.t8 3.56074
R54 VDD2.n0 VDD2.t0 3.56074
R55 VDD2.n6 VDD2.n4 0.534983
R56 VDD2 VDD2.n6 0.19231
R57 VDD2.n3 VDD2.n1 0.0787747
R58 VTAIL.n16 VTAIL.t7 64.5453
R59 VTAIL.n11 VTAIL.t10 64.5453
R60 VTAIL.n17 VTAIL.t9 64.5451
R61 VTAIL.n2 VTAIL.t4 64.5451
R62 VTAIL.n15 VTAIL.n14 60.9851
R63 VTAIL.n13 VTAIL.n12 60.9851
R64 VTAIL.n10 VTAIL.n9 60.9851
R65 VTAIL.n8 VTAIL.n7 60.9851
R66 VTAIL.n19 VTAIL.n18 60.9849
R67 VTAIL.n1 VTAIL.n0 60.9849
R68 VTAIL.n4 VTAIL.n3 60.9849
R69 VTAIL.n6 VTAIL.n5 60.9849
R70 VTAIL.n8 VTAIL.n6 21.3065
R71 VTAIL.n17 VTAIL.n16 20.7721
R72 VTAIL.n18 VTAIL.t14 3.56074
R73 VTAIL.n18 VTAIL.t15 3.56074
R74 VTAIL.n0 VTAIL.t8 3.56074
R75 VTAIL.n0 VTAIL.t17 3.56074
R76 VTAIL.n3 VTAIL.t5 3.56074
R77 VTAIL.n3 VTAIL.t18 3.56074
R78 VTAIL.n5 VTAIL.t3 3.56074
R79 VTAIL.n5 VTAIL.t2 3.56074
R80 VTAIL.n14 VTAIL.t19 3.56074
R81 VTAIL.n14 VTAIL.t1 3.56074
R82 VTAIL.n12 VTAIL.t6 3.56074
R83 VTAIL.n12 VTAIL.t0 3.56074
R84 VTAIL.n9 VTAIL.t16 3.56074
R85 VTAIL.n9 VTAIL.t12 3.56074
R86 VTAIL.n7 VTAIL.t13 3.56074
R87 VTAIL.n7 VTAIL.t11 3.56074
R88 VTAIL.n13 VTAIL.n11 0.737569
R89 VTAIL.n2 VTAIL.n1 0.737569
R90 VTAIL.n10 VTAIL.n8 0.534983
R91 VTAIL.n11 VTAIL.n10 0.534983
R92 VTAIL.n15 VTAIL.n13 0.534983
R93 VTAIL.n16 VTAIL.n15 0.534983
R94 VTAIL.n6 VTAIL.n4 0.534983
R95 VTAIL.n4 VTAIL.n2 0.534983
R96 VTAIL.n19 VTAIL.n17 0.534983
R97 VTAIL VTAIL.n1 0.459552
R98 VTAIL VTAIL.n19 0.075931
R99 VP.n21 VP.t0 902.655
R100 VP.n14 VP.t9 902.655
R101 VP.n5 VP.t6 902.655
R102 VP.n11 VP.t3 902.655
R103 VP.n18 VP.t1 867.601
R104 VP.n20 VP.t2 867.601
R105 VP.n13 VP.t8 867.601
R106 VP.n8 VP.t5 867.601
R107 VP.n4 VP.t7 867.601
R108 VP.n10 VP.t4 867.601
R109 VP.n6 VP.n5 161.489
R110 VP.n22 VP.n21 161.3
R111 VP.n6 VP.n3 161.3
R112 VP.n8 VP.n7 161.3
R113 VP.n9 VP.n2 161.3
R114 VP.n12 VP.n11 161.3
R115 VP.n19 VP.n0 161.3
R116 VP.n18 VP.n17 161.3
R117 VP.n16 VP.n1 161.3
R118 VP.n15 VP.n14 161.3
R119 VP.n18 VP.n1 73.0308
R120 VP.n19 VP.n18 73.0308
R121 VP.n8 VP.n3 73.0308
R122 VP.n9 VP.n8 73.0308
R123 VP.n14 VP.n13 55.5035
R124 VP.n21 VP.n20 55.5035
R125 VP.n5 VP.n4 55.5035
R126 VP.n11 VP.n10 55.5035
R127 VP.n15 VP.n12 38.4172
R128 VP.n13 VP.n1 17.5278
R129 VP.n20 VP.n19 17.5278
R130 VP.n4 VP.n3 17.5278
R131 VP.n10 VP.n9 17.5278
R132 VP.n7 VP.n6 0.189894
R133 VP.n7 VP.n2 0.189894
R134 VP.n12 VP.n2 0.189894
R135 VP.n16 VP.n15 0.189894
R136 VP.n17 VP.n16 0.189894
R137 VP.n17 VP.n0 0.189894
R138 VP.n22 VP.n0 0.189894
R139 VP VP.n22 0.0516364
R140 VDD1.n1 VDD1.t3 81.7586
R141 VDD1.n3 VDD1.t0 81.7584
R142 VDD1.n5 VDD1.n4 78.0092
R143 VDD1.n7 VDD1.n6 77.6639
R144 VDD1.n1 VDD1.n0 77.6639
R145 VDD1.n3 VDD1.n2 77.6636
R146 VDD1.n7 VDD1.n5 34.975
R147 VDD1.n6 VDD1.t5 3.56074
R148 VDD1.n6 VDD1.t6 3.56074
R149 VDD1.n0 VDD1.t2 3.56074
R150 VDD1.n0 VDD1.t4 3.56074
R151 VDD1.n4 VDD1.t7 3.56074
R152 VDD1.n4 VDD1.t9 3.56074
R153 VDD1.n2 VDD1.t1 3.56074
R154 VDD1.n2 VDD1.t8 3.56074
R155 VDD1 VDD1.n7 0.343172
R156 VDD1 VDD1.n1 0.19231
R157 VDD1.n5 VDD1.n3 0.0787747
R158 B.n90 B.t0 976.386
R159 B.n98 B.t9 976.386
R160 B.n28 B.t6 976.386
R161 B.n36 B.t3 976.386
R162 B.n327 B.n326 585
R163 B.n328 B.n53 585
R164 B.n330 B.n329 585
R165 B.n331 B.n52 585
R166 B.n333 B.n332 585
R167 B.n334 B.n51 585
R168 B.n336 B.n335 585
R169 B.n337 B.n50 585
R170 B.n339 B.n338 585
R171 B.n340 B.n49 585
R172 B.n342 B.n341 585
R173 B.n343 B.n48 585
R174 B.n345 B.n344 585
R175 B.n346 B.n47 585
R176 B.n348 B.n347 585
R177 B.n349 B.n46 585
R178 B.n351 B.n350 585
R179 B.n352 B.n45 585
R180 B.n354 B.n353 585
R181 B.n355 B.n44 585
R182 B.n357 B.n356 585
R183 B.n358 B.n43 585
R184 B.n360 B.n359 585
R185 B.n361 B.n42 585
R186 B.n363 B.n362 585
R187 B.n364 B.n41 585
R188 B.n366 B.n365 585
R189 B.n367 B.n40 585
R190 B.n369 B.n368 585
R191 B.n370 B.n39 585
R192 B.n372 B.n371 585
R193 B.n373 B.n38 585
R194 B.n375 B.n374 585
R195 B.n377 B.n35 585
R196 B.n379 B.n378 585
R197 B.n380 B.n34 585
R198 B.n382 B.n381 585
R199 B.n383 B.n33 585
R200 B.n385 B.n384 585
R201 B.n386 B.n32 585
R202 B.n388 B.n387 585
R203 B.n389 B.n31 585
R204 B.n391 B.n390 585
R205 B.n393 B.n392 585
R206 B.n394 B.n27 585
R207 B.n396 B.n395 585
R208 B.n397 B.n26 585
R209 B.n399 B.n398 585
R210 B.n400 B.n25 585
R211 B.n402 B.n401 585
R212 B.n403 B.n24 585
R213 B.n405 B.n404 585
R214 B.n406 B.n23 585
R215 B.n408 B.n407 585
R216 B.n409 B.n22 585
R217 B.n411 B.n410 585
R218 B.n412 B.n21 585
R219 B.n414 B.n413 585
R220 B.n415 B.n20 585
R221 B.n417 B.n416 585
R222 B.n418 B.n19 585
R223 B.n420 B.n419 585
R224 B.n421 B.n18 585
R225 B.n423 B.n422 585
R226 B.n424 B.n17 585
R227 B.n426 B.n425 585
R228 B.n427 B.n16 585
R229 B.n429 B.n428 585
R230 B.n430 B.n15 585
R231 B.n432 B.n431 585
R232 B.n433 B.n14 585
R233 B.n435 B.n434 585
R234 B.n436 B.n13 585
R235 B.n438 B.n437 585
R236 B.n439 B.n12 585
R237 B.n441 B.n440 585
R238 B.n325 B.n54 585
R239 B.n324 B.n323 585
R240 B.n322 B.n55 585
R241 B.n321 B.n320 585
R242 B.n319 B.n56 585
R243 B.n318 B.n317 585
R244 B.n316 B.n57 585
R245 B.n315 B.n314 585
R246 B.n313 B.n58 585
R247 B.n312 B.n311 585
R248 B.n310 B.n59 585
R249 B.n309 B.n308 585
R250 B.n307 B.n60 585
R251 B.n306 B.n305 585
R252 B.n304 B.n61 585
R253 B.n303 B.n302 585
R254 B.n301 B.n62 585
R255 B.n300 B.n299 585
R256 B.n298 B.n63 585
R257 B.n297 B.n296 585
R258 B.n295 B.n64 585
R259 B.n294 B.n293 585
R260 B.n292 B.n65 585
R261 B.n291 B.n290 585
R262 B.n289 B.n66 585
R263 B.n288 B.n287 585
R264 B.n286 B.n67 585
R265 B.n285 B.n284 585
R266 B.n283 B.n68 585
R267 B.n282 B.n281 585
R268 B.n280 B.n69 585
R269 B.n279 B.n278 585
R270 B.n277 B.n70 585
R271 B.n276 B.n275 585
R272 B.n274 B.n71 585
R273 B.n273 B.n272 585
R274 B.n271 B.n72 585
R275 B.n270 B.n269 585
R276 B.n268 B.n73 585
R277 B.n153 B.n152 585
R278 B.n154 B.n115 585
R279 B.n156 B.n155 585
R280 B.n157 B.n114 585
R281 B.n159 B.n158 585
R282 B.n160 B.n113 585
R283 B.n162 B.n161 585
R284 B.n163 B.n112 585
R285 B.n165 B.n164 585
R286 B.n166 B.n111 585
R287 B.n168 B.n167 585
R288 B.n169 B.n110 585
R289 B.n171 B.n170 585
R290 B.n172 B.n109 585
R291 B.n174 B.n173 585
R292 B.n175 B.n108 585
R293 B.n177 B.n176 585
R294 B.n178 B.n107 585
R295 B.n180 B.n179 585
R296 B.n181 B.n106 585
R297 B.n183 B.n182 585
R298 B.n184 B.n105 585
R299 B.n186 B.n185 585
R300 B.n187 B.n104 585
R301 B.n189 B.n188 585
R302 B.n190 B.n103 585
R303 B.n192 B.n191 585
R304 B.n193 B.n102 585
R305 B.n195 B.n194 585
R306 B.n196 B.n101 585
R307 B.n198 B.n197 585
R308 B.n199 B.n100 585
R309 B.n201 B.n200 585
R310 B.n203 B.n97 585
R311 B.n205 B.n204 585
R312 B.n206 B.n96 585
R313 B.n208 B.n207 585
R314 B.n209 B.n95 585
R315 B.n211 B.n210 585
R316 B.n212 B.n94 585
R317 B.n214 B.n213 585
R318 B.n215 B.n93 585
R319 B.n217 B.n216 585
R320 B.n219 B.n218 585
R321 B.n220 B.n89 585
R322 B.n222 B.n221 585
R323 B.n223 B.n88 585
R324 B.n225 B.n224 585
R325 B.n226 B.n87 585
R326 B.n228 B.n227 585
R327 B.n229 B.n86 585
R328 B.n231 B.n230 585
R329 B.n232 B.n85 585
R330 B.n234 B.n233 585
R331 B.n235 B.n84 585
R332 B.n237 B.n236 585
R333 B.n238 B.n83 585
R334 B.n240 B.n239 585
R335 B.n241 B.n82 585
R336 B.n243 B.n242 585
R337 B.n244 B.n81 585
R338 B.n246 B.n245 585
R339 B.n247 B.n80 585
R340 B.n249 B.n248 585
R341 B.n250 B.n79 585
R342 B.n252 B.n251 585
R343 B.n253 B.n78 585
R344 B.n255 B.n254 585
R345 B.n256 B.n77 585
R346 B.n258 B.n257 585
R347 B.n259 B.n76 585
R348 B.n261 B.n260 585
R349 B.n262 B.n75 585
R350 B.n264 B.n263 585
R351 B.n265 B.n74 585
R352 B.n267 B.n266 585
R353 B.n151 B.n116 585
R354 B.n150 B.n149 585
R355 B.n148 B.n117 585
R356 B.n147 B.n146 585
R357 B.n145 B.n118 585
R358 B.n144 B.n143 585
R359 B.n142 B.n119 585
R360 B.n141 B.n140 585
R361 B.n139 B.n120 585
R362 B.n138 B.n137 585
R363 B.n136 B.n121 585
R364 B.n135 B.n134 585
R365 B.n133 B.n122 585
R366 B.n132 B.n131 585
R367 B.n130 B.n123 585
R368 B.n129 B.n128 585
R369 B.n127 B.n124 585
R370 B.n126 B.n125 585
R371 B.n2 B.n0 585
R372 B.n469 B.n1 585
R373 B.n468 B.n467 585
R374 B.n466 B.n3 585
R375 B.n465 B.n464 585
R376 B.n463 B.n4 585
R377 B.n462 B.n461 585
R378 B.n460 B.n5 585
R379 B.n459 B.n458 585
R380 B.n457 B.n6 585
R381 B.n456 B.n455 585
R382 B.n454 B.n7 585
R383 B.n453 B.n452 585
R384 B.n451 B.n8 585
R385 B.n450 B.n449 585
R386 B.n448 B.n9 585
R387 B.n447 B.n446 585
R388 B.n445 B.n10 585
R389 B.n444 B.n443 585
R390 B.n442 B.n11 585
R391 B.n471 B.n470 585
R392 B.n152 B.n151 502.111
R393 B.n440 B.n11 502.111
R394 B.n266 B.n73 502.111
R395 B.n326 B.n325 502.111
R396 B.n151 B.n150 163.367
R397 B.n150 B.n117 163.367
R398 B.n146 B.n117 163.367
R399 B.n146 B.n145 163.367
R400 B.n145 B.n144 163.367
R401 B.n144 B.n119 163.367
R402 B.n140 B.n119 163.367
R403 B.n140 B.n139 163.367
R404 B.n139 B.n138 163.367
R405 B.n138 B.n121 163.367
R406 B.n134 B.n121 163.367
R407 B.n134 B.n133 163.367
R408 B.n133 B.n132 163.367
R409 B.n132 B.n123 163.367
R410 B.n128 B.n123 163.367
R411 B.n128 B.n127 163.367
R412 B.n127 B.n126 163.367
R413 B.n126 B.n2 163.367
R414 B.n470 B.n2 163.367
R415 B.n470 B.n469 163.367
R416 B.n469 B.n468 163.367
R417 B.n468 B.n3 163.367
R418 B.n464 B.n3 163.367
R419 B.n464 B.n463 163.367
R420 B.n463 B.n462 163.367
R421 B.n462 B.n5 163.367
R422 B.n458 B.n5 163.367
R423 B.n458 B.n457 163.367
R424 B.n457 B.n456 163.367
R425 B.n456 B.n7 163.367
R426 B.n452 B.n7 163.367
R427 B.n452 B.n451 163.367
R428 B.n451 B.n450 163.367
R429 B.n450 B.n9 163.367
R430 B.n446 B.n9 163.367
R431 B.n446 B.n445 163.367
R432 B.n445 B.n444 163.367
R433 B.n444 B.n11 163.367
R434 B.n152 B.n115 163.367
R435 B.n156 B.n115 163.367
R436 B.n157 B.n156 163.367
R437 B.n158 B.n157 163.367
R438 B.n158 B.n113 163.367
R439 B.n162 B.n113 163.367
R440 B.n163 B.n162 163.367
R441 B.n164 B.n163 163.367
R442 B.n164 B.n111 163.367
R443 B.n168 B.n111 163.367
R444 B.n169 B.n168 163.367
R445 B.n170 B.n169 163.367
R446 B.n170 B.n109 163.367
R447 B.n174 B.n109 163.367
R448 B.n175 B.n174 163.367
R449 B.n176 B.n175 163.367
R450 B.n176 B.n107 163.367
R451 B.n180 B.n107 163.367
R452 B.n181 B.n180 163.367
R453 B.n182 B.n181 163.367
R454 B.n182 B.n105 163.367
R455 B.n186 B.n105 163.367
R456 B.n187 B.n186 163.367
R457 B.n188 B.n187 163.367
R458 B.n188 B.n103 163.367
R459 B.n192 B.n103 163.367
R460 B.n193 B.n192 163.367
R461 B.n194 B.n193 163.367
R462 B.n194 B.n101 163.367
R463 B.n198 B.n101 163.367
R464 B.n199 B.n198 163.367
R465 B.n200 B.n199 163.367
R466 B.n200 B.n97 163.367
R467 B.n205 B.n97 163.367
R468 B.n206 B.n205 163.367
R469 B.n207 B.n206 163.367
R470 B.n207 B.n95 163.367
R471 B.n211 B.n95 163.367
R472 B.n212 B.n211 163.367
R473 B.n213 B.n212 163.367
R474 B.n213 B.n93 163.367
R475 B.n217 B.n93 163.367
R476 B.n218 B.n217 163.367
R477 B.n218 B.n89 163.367
R478 B.n222 B.n89 163.367
R479 B.n223 B.n222 163.367
R480 B.n224 B.n223 163.367
R481 B.n224 B.n87 163.367
R482 B.n228 B.n87 163.367
R483 B.n229 B.n228 163.367
R484 B.n230 B.n229 163.367
R485 B.n230 B.n85 163.367
R486 B.n234 B.n85 163.367
R487 B.n235 B.n234 163.367
R488 B.n236 B.n235 163.367
R489 B.n236 B.n83 163.367
R490 B.n240 B.n83 163.367
R491 B.n241 B.n240 163.367
R492 B.n242 B.n241 163.367
R493 B.n242 B.n81 163.367
R494 B.n246 B.n81 163.367
R495 B.n247 B.n246 163.367
R496 B.n248 B.n247 163.367
R497 B.n248 B.n79 163.367
R498 B.n252 B.n79 163.367
R499 B.n253 B.n252 163.367
R500 B.n254 B.n253 163.367
R501 B.n254 B.n77 163.367
R502 B.n258 B.n77 163.367
R503 B.n259 B.n258 163.367
R504 B.n260 B.n259 163.367
R505 B.n260 B.n75 163.367
R506 B.n264 B.n75 163.367
R507 B.n265 B.n264 163.367
R508 B.n266 B.n265 163.367
R509 B.n270 B.n73 163.367
R510 B.n271 B.n270 163.367
R511 B.n272 B.n271 163.367
R512 B.n272 B.n71 163.367
R513 B.n276 B.n71 163.367
R514 B.n277 B.n276 163.367
R515 B.n278 B.n277 163.367
R516 B.n278 B.n69 163.367
R517 B.n282 B.n69 163.367
R518 B.n283 B.n282 163.367
R519 B.n284 B.n283 163.367
R520 B.n284 B.n67 163.367
R521 B.n288 B.n67 163.367
R522 B.n289 B.n288 163.367
R523 B.n290 B.n289 163.367
R524 B.n290 B.n65 163.367
R525 B.n294 B.n65 163.367
R526 B.n295 B.n294 163.367
R527 B.n296 B.n295 163.367
R528 B.n296 B.n63 163.367
R529 B.n300 B.n63 163.367
R530 B.n301 B.n300 163.367
R531 B.n302 B.n301 163.367
R532 B.n302 B.n61 163.367
R533 B.n306 B.n61 163.367
R534 B.n307 B.n306 163.367
R535 B.n308 B.n307 163.367
R536 B.n308 B.n59 163.367
R537 B.n312 B.n59 163.367
R538 B.n313 B.n312 163.367
R539 B.n314 B.n313 163.367
R540 B.n314 B.n57 163.367
R541 B.n318 B.n57 163.367
R542 B.n319 B.n318 163.367
R543 B.n320 B.n319 163.367
R544 B.n320 B.n55 163.367
R545 B.n324 B.n55 163.367
R546 B.n325 B.n324 163.367
R547 B.n440 B.n439 163.367
R548 B.n439 B.n438 163.367
R549 B.n438 B.n13 163.367
R550 B.n434 B.n13 163.367
R551 B.n434 B.n433 163.367
R552 B.n433 B.n432 163.367
R553 B.n432 B.n15 163.367
R554 B.n428 B.n15 163.367
R555 B.n428 B.n427 163.367
R556 B.n427 B.n426 163.367
R557 B.n426 B.n17 163.367
R558 B.n422 B.n17 163.367
R559 B.n422 B.n421 163.367
R560 B.n421 B.n420 163.367
R561 B.n420 B.n19 163.367
R562 B.n416 B.n19 163.367
R563 B.n416 B.n415 163.367
R564 B.n415 B.n414 163.367
R565 B.n414 B.n21 163.367
R566 B.n410 B.n21 163.367
R567 B.n410 B.n409 163.367
R568 B.n409 B.n408 163.367
R569 B.n408 B.n23 163.367
R570 B.n404 B.n23 163.367
R571 B.n404 B.n403 163.367
R572 B.n403 B.n402 163.367
R573 B.n402 B.n25 163.367
R574 B.n398 B.n25 163.367
R575 B.n398 B.n397 163.367
R576 B.n397 B.n396 163.367
R577 B.n396 B.n27 163.367
R578 B.n392 B.n27 163.367
R579 B.n392 B.n391 163.367
R580 B.n391 B.n31 163.367
R581 B.n387 B.n31 163.367
R582 B.n387 B.n386 163.367
R583 B.n386 B.n385 163.367
R584 B.n385 B.n33 163.367
R585 B.n381 B.n33 163.367
R586 B.n381 B.n380 163.367
R587 B.n380 B.n379 163.367
R588 B.n379 B.n35 163.367
R589 B.n374 B.n35 163.367
R590 B.n374 B.n373 163.367
R591 B.n373 B.n372 163.367
R592 B.n372 B.n39 163.367
R593 B.n368 B.n39 163.367
R594 B.n368 B.n367 163.367
R595 B.n367 B.n366 163.367
R596 B.n366 B.n41 163.367
R597 B.n362 B.n41 163.367
R598 B.n362 B.n361 163.367
R599 B.n361 B.n360 163.367
R600 B.n360 B.n43 163.367
R601 B.n356 B.n43 163.367
R602 B.n356 B.n355 163.367
R603 B.n355 B.n354 163.367
R604 B.n354 B.n45 163.367
R605 B.n350 B.n45 163.367
R606 B.n350 B.n349 163.367
R607 B.n349 B.n348 163.367
R608 B.n348 B.n47 163.367
R609 B.n344 B.n47 163.367
R610 B.n344 B.n343 163.367
R611 B.n343 B.n342 163.367
R612 B.n342 B.n49 163.367
R613 B.n338 B.n49 163.367
R614 B.n338 B.n337 163.367
R615 B.n337 B.n336 163.367
R616 B.n336 B.n51 163.367
R617 B.n332 B.n51 163.367
R618 B.n332 B.n331 163.367
R619 B.n331 B.n330 163.367
R620 B.n330 B.n53 163.367
R621 B.n326 B.n53 163.367
R622 B.n90 B.t2 125.692
R623 B.n36 B.t4 125.692
R624 B.n98 B.t11 125.681
R625 B.n28 B.t7 125.681
R626 B.n91 B.t1 113.666
R627 B.n37 B.t5 113.666
R628 B.n99 B.t10 113.656
R629 B.n29 B.t8 113.656
R630 B.n92 B.n91 59.5399
R631 B.n202 B.n99 59.5399
R632 B.n30 B.n29 59.5399
R633 B.n376 B.n37 59.5399
R634 B.n442 B.n441 32.6249
R635 B.n327 B.n54 32.6249
R636 B.n268 B.n267 32.6249
R637 B.n153 B.n116 32.6249
R638 B B.n471 18.0485
R639 B.n91 B.n90 12.0247
R640 B.n99 B.n98 12.0247
R641 B.n29 B.n28 12.0247
R642 B.n37 B.n36 12.0247
R643 B.n441 B.n12 10.6151
R644 B.n437 B.n12 10.6151
R645 B.n437 B.n436 10.6151
R646 B.n436 B.n435 10.6151
R647 B.n435 B.n14 10.6151
R648 B.n431 B.n14 10.6151
R649 B.n431 B.n430 10.6151
R650 B.n430 B.n429 10.6151
R651 B.n429 B.n16 10.6151
R652 B.n425 B.n16 10.6151
R653 B.n425 B.n424 10.6151
R654 B.n424 B.n423 10.6151
R655 B.n423 B.n18 10.6151
R656 B.n419 B.n18 10.6151
R657 B.n419 B.n418 10.6151
R658 B.n418 B.n417 10.6151
R659 B.n417 B.n20 10.6151
R660 B.n413 B.n20 10.6151
R661 B.n413 B.n412 10.6151
R662 B.n412 B.n411 10.6151
R663 B.n411 B.n22 10.6151
R664 B.n407 B.n22 10.6151
R665 B.n407 B.n406 10.6151
R666 B.n406 B.n405 10.6151
R667 B.n405 B.n24 10.6151
R668 B.n401 B.n24 10.6151
R669 B.n401 B.n400 10.6151
R670 B.n400 B.n399 10.6151
R671 B.n399 B.n26 10.6151
R672 B.n395 B.n26 10.6151
R673 B.n395 B.n394 10.6151
R674 B.n394 B.n393 10.6151
R675 B.n390 B.n389 10.6151
R676 B.n389 B.n388 10.6151
R677 B.n388 B.n32 10.6151
R678 B.n384 B.n32 10.6151
R679 B.n384 B.n383 10.6151
R680 B.n383 B.n382 10.6151
R681 B.n382 B.n34 10.6151
R682 B.n378 B.n34 10.6151
R683 B.n378 B.n377 10.6151
R684 B.n375 B.n38 10.6151
R685 B.n371 B.n38 10.6151
R686 B.n371 B.n370 10.6151
R687 B.n370 B.n369 10.6151
R688 B.n369 B.n40 10.6151
R689 B.n365 B.n40 10.6151
R690 B.n365 B.n364 10.6151
R691 B.n364 B.n363 10.6151
R692 B.n363 B.n42 10.6151
R693 B.n359 B.n42 10.6151
R694 B.n359 B.n358 10.6151
R695 B.n358 B.n357 10.6151
R696 B.n357 B.n44 10.6151
R697 B.n353 B.n44 10.6151
R698 B.n353 B.n352 10.6151
R699 B.n352 B.n351 10.6151
R700 B.n351 B.n46 10.6151
R701 B.n347 B.n46 10.6151
R702 B.n347 B.n346 10.6151
R703 B.n346 B.n345 10.6151
R704 B.n345 B.n48 10.6151
R705 B.n341 B.n48 10.6151
R706 B.n341 B.n340 10.6151
R707 B.n340 B.n339 10.6151
R708 B.n339 B.n50 10.6151
R709 B.n335 B.n50 10.6151
R710 B.n335 B.n334 10.6151
R711 B.n334 B.n333 10.6151
R712 B.n333 B.n52 10.6151
R713 B.n329 B.n52 10.6151
R714 B.n329 B.n328 10.6151
R715 B.n328 B.n327 10.6151
R716 B.n269 B.n268 10.6151
R717 B.n269 B.n72 10.6151
R718 B.n273 B.n72 10.6151
R719 B.n274 B.n273 10.6151
R720 B.n275 B.n274 10.6151
R721 B.n275 B.n70 10.6151
R722 B.n279 B.n70 10.6151
R723 B.n280 B.n279 10.6151
R724 B.n281 B.n280 10.6151
R725 B.n281 B.n68 10.6151
R726 B.n285 B.n68 10.6151
R727 B.n286 B.n285 10.6151
R728 B.n287 B.n286 10.6151
R729 B.n287 B.n66 10.6151
R730 B.n291 B.n66 10.6151
R731 B.n292 B.n291 10.6151
R732 B.n293 B.n292 10.6151
R733 B.n293 B.n64 10.6151
R734 B.n297 B.n64 10.6151
R735 B.n298 B.n297 10.6151
R736 B.n299 B.n298 10.6151
R737 B.n299 B.n62 10.6151
R738 B.n303 B.n62 10.6151
R739 B.n304 B.n303 10.6151
R740 B.n305 B.n304 10.6151
R741 B.n305 B.n60 10.6151
R742 B.n309 B.n60 10.6151
R743 B.n310 B.n309 10.6151
R744 B.n311 B.n310 10.6151
R745 B.n311 B.n58 10.6151
R746 B.n315 B.n58 10.6151
R747 B.n316 B.n315 10.6151
R748 B.n317 B.n316 10.6151
R749 B.n317 B.n56 10.6151
R750 B.n321 B.n56 10.6151
R751 B.n322 B.n321 10.6151
R752 B.n323 B.n322 10.6151
R753 B.n323 B.n54 10.6151
R754 B.n154 B.n153 10.6151
R755 B.n155 B.n154 10.6151
R756 B.n155 B.n114 10.6151
R757 B.n159 B.n114 10.6151
R758 B.n160 B.n159 10.6151
R759 B.n161 B.n160 10.6151
R760 B.n161 B.n112 10.6151
R761 B.n165 B.n112 10.6151
R762 B.n166 B.n165 10.6151
R763 B.n167 B.n166 10.6151
R764 B.n167 B.n110 10.6151
R765 B.n171 B.n110 10.6151
R766 B.n172 B.n171 10.6151
R767 B.n173 B.n172 10.6151
R768 B.n173 B.n108 10.6151
R769 B.n177 B.n108 10.6151
R770 B.n178 B.n177 10.6151
R771 B.n179 B.n178 10.6151
R772 B.n179 B.n106 10.6151
R773 B.n183 B.n106 10.6151
R774 B.n184 B.n183 10.6151
R775 B.n185 B.n184 10.6151
R776 B.n185 B.n104 10.6151
R777 B.n189 B.n104 10.6151
R778 B.n190 B.n189 10.6151
R779 B.n191 B.n190 10.6151
R780 B.n191 B.n102 10.6151
R781 B.n195 B.n102 10.6151
R782 B.n196 B.n195 10.6151
R783 B.n197 B.n196 10.6151
R784 B.n197 B.n100 10.6151
R785 B.n201 B.n100 10.6151
R786 B.n204 B.n203 10.6151
R787 B.n204 B.n96 10.6151
R788 B.n208 B.n96 10.6151
R789 B.n209 B.n208 10.6151
R790 B.n210 B.n209 10.6151
R791 B.n210 B.n94 10.6151
R792 B.n214 B.n94 10.6151
R793 B.n215 B.n214 10.6151
R794 B.n216 B.n215 10.6151
R795 B.n220 B.n219 10.6151
R796 B.n221 B.n220 10.6151
R797 B.n221 B.n88 10.6151
R798 B.n225 B.n88 10.6151
R799 B.n226 B.n225 10.6151
R800 B.n227 B.n226 10.6151
R801 B.n227 B.n86 10.6151
R802 B.n231 B.n86 10.6151
R803 B.n232 B.n231 10.6151
R804 B.n233 B.n232 10.6151
R805 B.n233 B.n84 10.6151
R806 B.n237 B.n84 10.6151
R807 B.n238 B.n237 10.6151
R808 B.n239 B.n238 10.6151
R809 B.n239 B.n82 10.6151
R810 B.n243 B.n82 10.6151
R811 B.n244 B.n243 10.6151
R812 B.n245 B.n244 10.6151
R813 B.n245 B.n80 10.6151
R814 B.n249 B.n80 10.6151
R815 B.n250 B.n249 10.6151
R816 B.n251 B.n250 10.6151
R817 B.n251 B.n78 10.6151
R818 B.n255 B.n78 10.6151
R819 B.n256 B.n255 10.6151
R820 B.n257 B.n256 10.6151
R821 B.n257 B.n76 10.6151
R822 B.n261 B.n76 10.6151
R823 B.n262 B.n261 10.6151
R824 B.n263 B.n262 10.6151
R825 B.n263 B.n74 10.6151
R826 B.n267 B.n74 10.6151
R827 B.n149 B.n116 10.6151
R828 B.n149 B.n148 10.6151
R829 B.n148 B.n147 10.6151
R830 B.n147 B.n118 10.6151
R831 B.n143 B.n118 10.6151
R832 B.n143 B.n142 10.6151
R833 B.n142 B.n141 10.6151
R834 B.n141 B.n120 10.6151
R835 B.n137 B.n120 10.6151
R836 B.n137 B.n136 10.6151
R837 B.n136 B.n135 10.6151
R838 B.n135 B.n122 10.6151
R839 B.n131 B.n122 10.6151
R840 B.n131 B.n130 10.6151
R841 B.n130 B.n129 10.6151
R842 B.n129 B.n124 10.6151
R843 B.n125 B.n124 10.6151
R844 B.n125 B.n0 10.6151
R845 B.n467 B.n1 10.6151
R846 B.n467 B.n466 10.6151
R847 B.n466 B.n465 10.6151
R848 B.n465 B.n4 10.6151
R849 B.n461 B.n4 10.6151
R850 B.n461 B.n460 10.6151
R851 B.n460 B.n459 10.6151
R852 B.n459 B.n6 10.6151
R853 B.n455 B.n6 10.6151
R854 B.n455 B.n454 10.6151
R855 B.n454 B.n453 10.6151
R856 B.n453 B.n8 10.6151
R857 B.n449 B.n8 10.6151
R858 B.n449 B.n448 10.6151
R859 B.n448 B.n447 10.6151
R860 B.n447 B.n10 10.6151
R861 B.n443 B.n10 10.6151
R862 B.n443 B.n442 10.6151
R863 B.n393 B.n30 9.36635
R864 B.n376 B.n375 9.36635
R865 B.n202 B.n201 9.36635
R866 B.n219 B.n92 9.36635
R867 B.n471 B.n0 2.81026
R868 B.n471 B.n1 2.81026
R869 B.n390 B.n30 1.24928
R870 B.n377 B.n376 1.24928
R871 B.n203 B.n202 1.24928
R872 B.n216 B.n92 1.24928
C0 VDD1 VTAIL 16.6386f
C1 VDD2 VP 0.288937f
C2 B VTAIL 1.97081f
C3 VDD1 VN 0.148026f
C4 B VN 0.657883f
C5 VP VDD1 3.18964f
C6 B VP 1.0084f
C7 w_n1714_n2794# VTAIL 2.57526f
C8 w_n1714_n2794# VN 2.91129f
C9 VDD2 VDD1 0.718743f
C10 B VDD2 1.34759f
C11 VP w_n1714_n2794# 3.12732f
C12 B VDD1 1.31898f
C13 VN VTAIL 2.77389f
C14 VDD2 w_n1714_n2794# 1.65814f
C15 VP VTAIL 2.7885f
C16 VP VN 4.4627f
C17 w_n1714_n2794# VDD1 1.63451f
C18 B w_n1714_n2794# 5.88195f
C19 VDD2 VTAIL 16.6702f
C20 VDD2 VN 3.05272f
C21 VDD2 VSUBS 1.319863f
C22 VDD1 VSUBS 0.920679f
C23 VTAIL VSUBS 0.508422f
C24 VN VSUBS 4.36482f
C25 VP VSUBS 1.201595f
C26 B VSUBS 2.2501f
C27 w_n1714_n2794# VSUBS 59.256397f
C28 B.n0 VSUBS 0.003861f
C29 B.n1 VSUBS 0.003861f
C30 B.n2 VSUBS 0.006106f
C31 B.n3 VSUBS 0.006106f
C32 B.n4 VSUBS 0.006106f
C33 B.n5 VSUBS 0.006106f
C34 B.n6 VSUBS 0.006106f
C35 B.n7 VSUBS 0.006106f
C36 B.n8 VSUBS 0.006106f
C37 B.n9 VSUBS 0.006106f
C38 B.n10 VSUBS 0.006106f
C39 B.n11 VSUBS 0.013881f
C40 B.n12 VSUBS 0.006106f
C41 B.n13 VSUBS 0.006106f
C42 B.n14 VSUBS 0.006106f
C43 B.n15 VSUBS 0.006106f
C44 B.n16 VSUBS 0.006106f
C45 B.n17 VSUBS 0.006106f
C46 B.n18 VSUBS 0.006106f
C47 B.n19 VSUBS 0.006106f
C48 B.n20 VSUBS 0.006106f
C49 B.n21 VSUBS 0.006106f
C50 B.n22 VSUBS 0.006106f
C51 B.n23 VSUBS 0.006106f
C52 B.n24 VSUBS 0.006106f
C53 B.n25 VSUBS 0.006106f
C54 B.n26 VSUBS 0.006106f
C55 B.n27 VSUBS 0.006106f
C56 B.t8 VSUBS 0.250796f
C57 B.t7 VSUBS 0.255137f
C58 B.t6 VSUBS 0.091681f
C59 B.n28 VSUBS 0.074585f
C60 B.n29 VSUBS 0.054091f
C61 B.n30 VSUBS 0.014147f
C62 B.n31 VSUBS 0.006106f
C63 B.n32 VSUBS 0.006106f
C64 B.n33 VSUBS 0.006106f
C65 B.n34 VSUBS 0.006106f
C66 B.n35 VSUBS 0.006106f
C67 B.t5 VSUBS 0.250793f
C68 B.t4 VSUBS 0.255135f
C69 B.t3 VSUBS 0.091681f
C70 B.n36 VSUBS 0.074588f
C71 B.n37 VSUBS 0.054093f
C72 B.n38 VSUBS 0.006106f
C73 B.n39 VSUBS 0.006106f
C74 B.n40 VSUBS 0.006106f
C75 B.n41 VSUBS 0.006106f
C76 B.n42 VSUBS 0.006106f
C77 B.n43 VSUBS 0.006106f
C78 B.n44 VSUBS 0.006106f
C79 B.n45 VSUBS 0.006106f
C80 B.n46 VSUBS 0.006106f
C81 B.n47 VSUBS 0.006106f
C82 B.n48 VSUBS 0.006106f
C83 B.n49 VSUBS 0.006106f
C84 B.n50 VSUBS 0.006106f
C85 B.n51 VSUBS 0.006106f
C86 B.n52 VSUBS 0.006106f
C87 B.n53 VSUBS 0.006106f
C88 B.n54 VSUBS 0.014603f
C89 B.n55 VSUBS 0.006106f
C90 B.n56 VSUBS 0.006106f
C91 B.n57 VSUBS 0.006106f
C92 B.n58 VSUBS 0.006106f
C93 B.n59 VSUBS 0.006106f
C94 B.n60 VSUBS 0.006106f
C95 B.n61 VSUBS 0.006106f
C96 B.n62 VSUBS 0.006106f
C97 B.n63 VSUBS 0.006106f
C98 B.n64 VSUBS 0.006106f
C99 B.n65 VSUBS 0.006106f
C100 B.n66 VSUBS 0.006106f
C101 B.n67 VSUBS 0.006106f
C102 B.n68 VSUBS 0.006106f
C103 B.n69 VSUBS 0.006106f
C104 B.n70 VSUBS 0.006106f
C105 B.n71 VSUBS 0.006106f
C106 B.n72 VSUBS 0.006106f
C107 B.n73 VSUBS 0.013881f
C108 B.n74 VSUBS 0.006106f
C109 B.n75 VSUBS 0.006106f
C110 B.n76 VSUBS 0.006106f
C111 B.n77 VSUBS 0.006106f
C112 B.n78 VSUBS 0.006106f
C113 B.n79 VSUBS 0.006106f
C114 B.n80 VSUBS 0.006106f
C115 B.n81 VSUBS 0.006106f
C116 B.n82 VSUBS 0.006106f
C117 B.n83 VSUBS 0.006106f
C118 B.n84 VSUBS 0.006106f
C119 B.n85 VSUBS 0.006106f
C120 B.n86 VSUBS 0.006106f
C121 B.n87 VSUBS 0.006106f
C122 B.n88 VSUBS 0.006106f
C123 B.n89 VSUBS 0.006106f
C124 B.t1 VSUBS 0.250793f
C125 B.t2 VSUBS 0.255135f
C126 B.t0 VSUBS 0.091681f
C127 B.n90 VSUBS 0.074588f
C128 B.n91 VSUBS 0.054093f
C129 B.n92 VSUBS 0.014147f
C130 B.n93 VSUBS 0.006106f
C131 B.n94 VSUBS 0.006106f
C132 B.n95 VSUBS 0.006106f
C133 B.n96 VSUBS 0.006106f
C134 B.n97 VSUBS 0.006106f
C135 B.t10 VSUBS 0.250796f
C136 B.t11 VSUBS 0.255137f
C137 B.t9 VSUBS 0.091681f
C138 B.n98 VSUBS 0.074585f
C139 B.n99 VSUBS 0.054091f
C140 B.n100 VSUBS 0.006106f
C141 B.n101 VSUBS 0.006106f
C142 B.n102 VSUBS 0.006106f
C143 B.n103 VSUBS 0.006106f
C144 B.n104 VSUBS 0.006106f
C145 B.n105 VSUBS 0.006106f
C146 B.n106 VSUBS 0.006106f
C147 B.n107 VSUBS 0.006106f
C148 B.n108 VSUBS 0.006106f
C149 B.n109 VSUBS 0.006106f
C150 B.n110 VSUBS 0.006106f
C151 B.n111 VSUBS 0.006106f
C152 B.n112 VSUBS 0.006106f
C153 B.n113 VSUBS 0.006106f
C154 B.n114 VSUBS 0.006106f
C155 B.n115 VSUBS 0.006106f
C156 B.n116 VSUBS 0.013881f
C157 B.n117 VSUBS 0.006106f
C158 B.n118 VSUBS 0.006106f
C159 B.n119 VSUBS 0.006106f
C160 B.n120 VSUBS 0.006106f
C161 B.n121 VSUBS 0.006106f
C162 B.n122 VSUBS 0.006106f
C163 B.n123 VSUBS 0.006106f
C164 B.n124 VSUBS 0.006106f
C165 B.n125 VSUBS 0.006106f
C166 B.n126 VSUBS 0.006106f
C167 B.n127 VSUBS 0.006106f
C168 B.n128 VSUBS 0.006106f
C169 B.n129 VSUBS 0.006106f
C170 B.n130 VSUBS 0.006106f
C171 B.n131 VSUBS 0.006106f
C172 B.n132 VSUBS 0.006106f
C173 B.n133 VSUBS 0.006106f
C174 B.n134 VSUBS 0.006106f
C175 B.n135 VSUBS 0.006106f
C176 B.n136 VSUBS 0.006106f
C177 B.n137 VSUBS 0.006106f
C178 B.n138 VSUBS 0.006106f
C179 B.n139 VSUBS 0.006106f
C180 B.n140 VSUBS 0.006106f
C181 B.n141 VSUBS 0.006106f
C182 B.n142 VSUBS 0.006106f
C183 B.n143 VSUBS 0.006106f
C184 B.n144 VSUBS 0.006106f
C185 B.n145 VSUBS 0.006106f
C186 B.n146 VSUBS 0.006106f
C187 B.n147 VSUBS 0.006106f
C188 B.n148 VSUBS 0.006106f
C189 B.n149 VSUBS 0.006106f
C190 B.n150 VSUBS 0.006106f
C191 B.n151 VSUBS 0.013881f
C192 B.n152 VSUBS 0.014674f
C193 B.n153 VSUBS 0.014674f
C194 B.n154 VSUBS 0.006106f
C195 B.n155 VSUBS 0.006106f
C196 B.n156 VSUBS 0.006106f
C197 B.n157 VSUBS 0.006106f
C198 B.n158 VSUBS 0.006106f
C199 B.n159 VSUBS 0.006106f
C200 B.n160 VSUBS 0.006106f
C201 B.n161 VSUBS 0.006106f
C202 B.n162 VSUBS 0.006106f
C203 B.n163 VSUBS 0.006106f
C204 B.n164 VSUBS 0.006106f
C205 B.n165 VSUBS 0.006106f
C206 B.n166 VSUBS 0.006106f
C207 B.n167 VSUBS 0.006106f
C208 B.n168 VSUBS 0.006106f
C209 B.n169 VSUBS 0.006106f
C210 B.n170 VSUBS 0.006106f
C211 B.n171 VSUBS 0.006106f
C212 B.n172 VSUBS 0.006106f
C213 B.n173 VSUBS 0.006106f
C214 B.n174 VSUBS 0.006106f
C215 B.n175 VSUBS 0.006106f
C216 B.n176 VSUBS 0.006106f
C217 B.n177 VSUBS 0.006106f
C218 B.n178 VSUBS 0.006106f
C219 B.n179 VSUBS 0.006106f
C220 B.n180 VSUBS 0.006106f
C221 B.n181 VSUBS 0.006106f
C222 B.n182 VSUBS 0.006106f
C223 B.n183 VSUBS 0.006106f
C224 B.n184 VSUBS 0.006106f
C225 B.n185 VSUBS 0.006106f
C226 B.n186 VSUBS 0.006106f
C227 B.n187 VSUBS 0.006106f
C228 B.n188 VSUBS 0.006106f
C229 B.n189 VSUBS 0.006106f
C230 B.n190 VSUBS 0.006106f
C231 B.n191 VSUBS 0.006106f
C232 B.n192 VSUBS 0.006106f
C233 B.n193 VSUBS 0.006106f
C234 B.n194 VSUBS 0.006106f
C235 B.n195 VSUBS 0.006106f
C236 B.n196 VSUBS 0.006106f
C237 B.n197 VSUBS 0.006106f
C238 B.n198 VSUBS 0.006106f
C239 B.n199 VSUBS 0.006106f
C240 B.n200 VSUBS 0.006106f
C241 B.n201 VSUBS 0.005747f
C242 B.n202 VSUBS 0.014147f
C243 B.n203 VSUBS 0.003412f
C244 B.n204 VSUBS 0.006106f
C245 B.n205 VSUBS 0.006106f
C246 B.n206 VSUBS 0.006106f
C247 B.n207 VSUBS 0.006106f
C248 B.n208 VSUBS 0.006106f
C249 B.n209 VSUBS 0.006106f
C250 B.n210 VSUBS 0.006106f
C251 B.n211 VSUBS 0.006106f
C252 B.n212 VSUBS 0.006106f
C253 B.n213 VSUBS 0.006106f
C254 B.n214 VSUBS 0.006106f
C255 B.n215 VSUBS 0.006106f
C256 B.n216 VSUBS 0.003412f
C257 B.n217 VSUBS 0.006106f
C258 B.n218 VSUBS 0.006106f
C259 B.n219 VSUBS 0.005747f
C260 B.n220 VSUBS 0.006106f
C261 B.n221 VSUBS 0.006106f
C262 B.n222 VSUBS 0.006106f
C263 B.n223 VSUBS 0.006106f
C264 B.n224 VSUBS 0.006106f
C265 B.n225 VSUBS 0.006106f
C266 B.n226 VSUBS 0.006106f
C267 B.n227 VSUBS 0.006106f
C268 B.n228 VSUBS 0.006106f
C269 B.n229 VSUBS 0.006106f
C270 B.n230 VSUBS 0.006106f
C271 B.n231 VSUBS 0.006106f
C272 B.n232 VSUBS 0.006106f
C273 B.n233 VSUBS 0.006106f
C274 B.n234 VSUBS 0.006106f
C275 B.n235 VSUBS 0.006106f
C276 B.n236 VSUBS 0.006106f
C277 B.n237 VSUBS 0.006106f
C278 B.n238 VSUBS 0.006106f
C279 B.n239 VSUBS 0.006106f
C280 B.n240 VSUBS 0.006106f
C281 B.n241 VSUBS 0.006106f
C282 B.n242 VSUBS 0.006106f
C283 B.n243 VSUBS 0.006106f
C284 B.n244 VSUBS 0.006106f
C285 B.n245 VSUBS 0.006106f
C286 B.n246 VSUBS 0.006106f
C287 B.n247 VSUBS 0.006106f
C288 B.n248 VSUBS 0.006106f
C289 B.n249 VSUBS 0.006106f
C290 B.n250 VSUBS 0.006106f
C291 B.n251 VSUBS 0.006106f
C292 B.n252 VSUBS 0.006106f
C293 B.n253 VSUBS 0.006106f
C294 B.n254 VSUBS 0.006106f
C295 B.n255 VSUBS 0.006106f
C296 B.n256 VSUBS 0.006106f
C297 B.n257 VSUBS 0.006106f
C298 B.n258 VSUBS 0.006106f
C299 B.n259 VSUBS 0.006106f
C300 B.n260 VSUBS 0.006106f
C301 B.n261 VSUBS 0.006106f
C302 B.n262 VSUBS 0.006106f
C303 B.n263 VSUBS 0.006106f
C304 B.n264 VSUBS 0.006106f
C305 B.n265 VSUBS 0.006106f
C306 B.n266 VSUBS 0.014674f
C307 B.n267 VSUBS 0.014674f
C308 B.n268 VSUBS 0.013881f
C309 B.n269 VSUBS 0.006106f
C310 B.n270 VSUBS 0.006106f
C311 B.n271 VSUBS 0.006106f
C312 B.n272 VSUBS 0.006106f
C313 B.n273 VSUBS 0.006106f
C314 B.n274 VSUBS 0.006106f
C315 B.n275 VSUBS 0.006106f
C316 B.n276 VSUBS 0.006106f
C317 B.n277 VSUBS 0.006106f
C318 B.n278 VSUBS 0.006106f
C319 B.n279 VSUBS 0.006106f
C320 B.n280 VSUBS 0.006106f
C321 B.n281 VSUBS 0.006106f
C322 B.n282 VSUBS 0.006106f
C323 B.n283 VSUBS 0.006106f
C324 B.n284 VSUBS 0.006106f
C325 B.n285 VSUBS 0.006106f
C326 B.n286 VSUBS 0.006106f
C327 B.n287 VSUBS 0.006106f
C328 B.n288 VSUBS 0.006106f
C329 B.n289 VSUBS 0.006106f
C330 B.n290 VSUBS 0.006106f
C331 B.n291 VSUBS 0.006106f
C332 B.n292 VSUBS 0.006106f
C333 B.n293 VSUBS 0.006106f
C334 B.n294 VSUBS 0.006106f
C335 B.n295 VSUBS 0.006106f
C336 B.n296 VSUBS 0.006106f
C337 B.n297 VSUBS 0.006106f
C338 B.n298 VSUBS 0.006106f
C339 B.n299 VSUBS 0.006106f
C340 B.n300 VSUBS 0.006106f
C341 B.n301 VSUBS 0.006106f
C342 B.n302 VSUBS 0.006106f
C343 B.n303 VSUBS 0.006106f
C344 B.n304 VSUBS 0.006106f
C345 B.n305 VSUBS 0.006106f
C346 B.n306 VSUBS 0.006106f
C347 B.n307 VSUBS 0.006106f
C348 B.n308 VSUBS 0.006106f
C349 B.n309 VSUBS 0.006106f
C350 B.n310 VSUBS 0.006106f
C351 B.n311 VSUBS 0.006106f
C352 B.n312 VSUBS 0.006106f
C353 B.n313 VSUBS 0.006106f
C354 B.n314 VSUBS 0.006106f
C355 B.n315 VSUBS 0.006106f
C356 B.n316 VSUBS 0.006106f
C357 B.n317 VSUBS 0.006106f
C358 B.n318 VSUBS 0.006106f
C359 B.n319 VSUBS 0.006106f
C360 B.n320 VSUBS 0.006106f
C361 B.n321 VSUBS 0.006106f
C362 B.n322 VSUBS 0.006106f
C363 B.n323 VSUBS 0.006106f
C364 B.n324 VSUBS 0.006106f
C365 B.n325 VSUBS 0.013881f
C366 B.n326 VSUBS 0.014674f
C367 B.n327 VSUBS 0.013951f
C368 B.n328 VSUBS 0.006106f
C369 B.n329 VSUBS 0.006106f
C370 B.n330 VSUBS 0.006106f
C371 B.n331 VSUBS 0.006106f
C372 B.n332 VSUBS 0.006106f
C373 B.n333 VSUBS 0.006106f
C374 B.n334 VSUBS 0.006106f
C375 B.n335 VSUBS 0.006106f
C376 B.n336 VSUBS 0.006106f
C377 B.n337 VSUBS 0.006106f
C378 B.n338 VSUBS 0.006106f
C379 B.n339 VSUBS 0.006106f
C380 B.n340 VSUBS 0.006106f
C381 B.n341 VSUBS 0.006106f
C382 B.n342 VSUBS 0.006106f
C383 B.n343 VSUBS 0.006106f
C384 B.n344 VSUBS 0.006106f
C385 B.n345 VSUBS 0.006106f
C386 B.n346 VSUBS 0.006106f
C387 B.n347 VSUBS 0.006106f
C388 B.n348 VSUBS 0.006106f
C389 B.n349 VSUBS 0.006106f
C390 B.n350 VSUBS 0.006106f
C391 B.n351 VSUBS 0.006106f
C392 B.n352 VSUBS 0.006106f
C393 B.n353 VSUBS 0.006106f
C394 B.n354 VSUBS 0.006106f
C395 B.n355 VSUBS 0.006106f
C396 B.n356 VSUBS 0.006106f
C397 B.n357 VSUBS 0.006106f
C398 B.n358 VSUBS 0.006106f
C399 B.n359 VSUBS 0.006106f
C400 B.n360 VSUBS 0.006106f
C401 B.n361 VSUBS 0.006106f
C402 B.n362 VSUBS 0.006106f
C403 B.n363 VSUBS 0.006106f
C404 B.n364 VSUBS 0.006106f
C405 B.n365 VSUBS 0.006106f
C406 B.n366 VSUBS 0.006106f
C407 B.n367 VSUBS 0.006106f
C408 B.n368 VSUBS 0.006106f
C409 B.n369 VSUBS 0.006106f
C410 B.n370 VSUBS 0.006106f
C411 B.n371 VSUBS 0.006106f
C412 B.n372 VSUBS 0.006106f
C413 B.n373 VSUBS 0.006106f
C414 B.n374 VSUBS 0.006106f
C415 B.n375 VSUBS 0.005747f
C416 B.n376 VSUBS 0.014147f
C417 B.n377 VSUBS 0.003412f
C418 B.n378 VSUBS 0.006106f
C419 B.n379 VSUBS 0.006106f
C420 B.n380 VSUBS 0.006106f
C421 B.n381 VSUBS 0.006106f
C422 B.n382 VSUBS 0.006106f
C423 B.n383 VSUBS 0.006106f
C424 B.n384 VSUBS 0.006106f
C425 B.n385 VSUBS 0.006106f
C426 B.n386 VSUBS 0.006106f
C427 B.n387 VSUBS 0.006106f
C428 B.n388 VSUBS 0.006106f
C429 B.n389 VSUBS 0.006106f
C430 B.n390 VSUBS 0.003412f
C431 B.n391 VSUBS 0.006106f
C432 B.n392 VSUBS 0.006106f
C433 B.n393 VSUBS 0.005747f
C434 B.n394 VSUBS 0.006106f
C435 B.n395 VSUBS 0.006106f
C436 B.n396 VSUBS 0.006106f
C437 B.n397 VSUBS 0.006106f
C438 B.n398 VSUBS 0.006106f
C439 B.n399 VSUBS 0.006106f
C440 B.n400 VSUBS 0.006106f
C441 B.n401 VSUBS 0.006106f
C442 B.n402 VSUBS 0.006106f
C443 B.n403 VSUBS 0.006106f
C444 B.n404 VSUBS 0.006106f
C445 B.n405 VSUBS 0.006106f
C446 B.n406 VSUBS 0.006106f
C447 B.n407 VSUBS 0.006106f
C448 B.n408 VSUBS 0.006106f
C449 B.n409 VSUBS 0.006106f
C450 B.n410 VSUBS 0.006106f
C451 B.n411 VSUBS 0.006106f
C452 B.n412 VSUBS 0.006106f
C453 B.n413 VSUBS 0.006106f
C454 B.n414 VSUBS 0.006106f
C455 B.n415 VSUBS 0.006106f
C456 B.n416 VSUBS 0.006106f
C457 B.n417 VSUBS 0.006106f
C458 B.n418 VSUBS 0.006106f
C459 B.n419 VSUBS 0.006106f
C460 B.n420 VSUBS 0.006106f
C461 B.n421 VSUBS 0.006106f
C462 B.n422 VSUBS 0.006106f
C463 B.n423 VSUBS 0.006106f
C464 B.n424 VSUBS 0.006106f
C465 B.n425 VSUBS 0.006106f
C466 B.n426 VSUBS 0.006106f
C467 B.n427 VSUBS 0.006106f
C468 B.n428 VSUBS 0.006106f
C469 B.n429 VSUBS 0.006106f
C470 B.n430 VSUBS 0.006106f
C471 B.n431 VSUBS 0.006106f
C472 B.n432 VSUBS 0.006106f
C473 B.n433 VSUBS 0.006106f
C474 B.n434 VSUBS 0.006106f
C475 B.n435 VSUBS 0.006106f
C476 B.n436 VSUBS 0.006106f
C477 B.n437 VSUBS 0.006106f
C478 B.n438 VSUBS 0.006106f
C479 B.n439 VSUBS 0.006106f
C480 B.n440 VSUBS 0.014674f
C481 B.n441 VSUBS 0.014674f
C482 B.n442 VSUBS 0.013881f
C483 B.n443 VSUBS 0.006106f
C484 B.n444 VSUBS 0.006106f
C485 B.n445 VSUBS 0.006106f
C486 B.n446 VSUBS 0.006106f
C487 B.n447 VSUBS 0.006106f
C488 B.n448 VSUBS 0.006106f
C489 B.n449 VSUBS 0.006106f
C490 B.n450 VSUBS 0.006106f
C491 B.n451 VSUBS 0.006106f
C492 B.n452 VSUBS 0.006106f
C493 B.n453 VSUBS 0.006106f
C494 B.n454 VSUBS 0.006106f
C495 B.n455 VSUBS 0.006106f
C496 B.n456 VSUBS 0.006106f
C497 B.n457 VSUBS 0.006106f
C498 B.n458 VSUBS 0.006106f
C499 B.n459 VSUBS 0.006106f
C500 B.n460 VSUBS 0.006106f
C501 B.n461 VSUBS 0.006106f
C502 B.n462 VSUBS 0.006106f
C503 B.n463 VSUBS 0.006106f
C504 B.n464 VSUBS 0.006106f
C505 B.n465 VSUBS 0.006106f
C506 B.n466 VSUBS 0.006106f
C507 B.n467 VSUBS 0.006106f
C508 B.n468 VSUBS 0.006106f
C509 B.n469 VSUBS 0.006106f
C510 B.n470 VSUBS 0.006106f
C511 B.n471 VSUBS 0.013826f
C512 VDD1.t3 VSUBS 2.08863f
C513 VDD1.t2 VSUBS 0.216078f
C514 VDD1.t4 VSUBS 0.216078f
C515 VDD1.n0 VSUBS 1.58037f
C516 VDD1.n1 VSUBS 1.31848f
C517 VDD1.t0 VSUBS 2.08862f
C518 VDD1.t1 VSUBS 0.216078f
C519 VDD1.t8 VSUBS 0.216078f
C520 VDD1.n2 VSUBS 1.58037f
C521 VDD1.n3 VSUBS 1.31641f
C522 VDD1.t7 VSUBS 0.216078f
C523 VDD1.t9 VSUBS 0.216078f
C524 VDD1.n4 VSUBS 1.58325f
C525 VDD1.n5 VSUBS 2.19245f
C526 VDD1.t5 VSUBS 0.216078f
C527 VDD1.t6 VSUBS 0.216078f
C528 VDD1.n6 VSUBS 1.58037f
C529 VDD1.n7 VSUBS 2.69083f
C530 VP.n0 VSUBS 0.071403f
C531 VP.t2 VSUBS 0.535813f
C532 VP.t1 VSUBS 0.535813f
C533 VP.n1 VSUBS 0.02897f
C534 VP.n2 VSUBS 0.071403f
C535 VP.t4 VSUBS 0.535813f
C536 VP.t5 VSUBS 0.535813f
C537 VP.n3 VSUBS 0.02897f
C538 VP.t6 VSUBS 0.544561f
C539 VP.t7 VSUBS 0.535813f
C540 VP.n4 VSUBS 0.223957f
C541 VP.n5 VSUBS 0.245596f
C542 VP.n6 VSUBS 0.154594f
C543 VP.n7 VSUBS 0.071403f
C544 VP.n8 VSUBS 0.247644f
C545 VP.n9 VSUBS 0.02897f
C546 VP.n10 VSUBS 0.223957f
C547 VP.t3 VSUBS 0.544561f
C548 VP.n11 VSUBS 0.245498f
C549 VP.n12 VSUBS 2.52804f
C550 VP.t9 VSUBS 0.544561f
C551 VP.t8 VSUBS 0.535813f
C552 VP.n13 VSUBS 0.223957f
C553 VP.n14 VSUBS 0.245498f
C554 VP.n15 VSUBS 2.59485f
C555 VP.n16 VSUBS 0.071403f
C556 VP.n17 VSUBS 0.071403f
C557 VP.n18 VSUBS 0.247644f
C558 VP.n19 VSUBS 0.02897f
C559 VP.n20 VSUBS 0.223957f
C560 VP.t0 VSUBS 0.544561f
C561 VP.n21 VSUBS 0.245498f
C562 VP.n22 VSUBS 0.055334f
C563 VTAIL.t8 VSUBS 0.242375f
C564 VTAIL.t17 VSUBS 0.242375f
C565 VTAIL.n0 VSUBS 1.60515f
C566 VTAIL.n1 VSUBS 0.870383f
C567 VTAIL.t4 VSUBS 2.15454f
C568 VTAIL.n2 VSUBS 0.990181f
C569 VTAIL.t5 VSUBS 0.242375f
C570 VTAIL.t18 VSUBS 0.242375f
C571 VTAIL.n3 VSUBS 1.60515f
C572 VTAIL.n4 VSUBS 0.856619f
C573 VTAIL.t3 VSUBS 0.242375f
C574 VTAIL.t2 VSUBS 0.242375f
C575 VTAIL.n5 VSUBS 1.60515f
C576 VTAIL.n6 VSUBS 2.2228f
C577 VTAIL.t13 VSUBS 0.242375f
C578 VTAIL.t11 VSUBS 0.242375f
C579 VTAIL.n7 VSUBS 1.60516f
C580 VTAIL.n8 VSUBS 2.22279f
C581 VTAIL.t16 VSUBS 0.242375f
C582 VTAIL.t12 VSUBS 0.242375f
C583 VTAIL.n9 VSUBS 1.60516f
C584 VTAIL.n10 VSUBS 0.856608f
C585 VTAIL.t10 VSUBS 2.15455f
C586 VTAIL.n11 VSUBS 0.990168f
C587 VTAIL.t6 VSUBS 0.242375f
C588 VTAIL.t0 VSUBS 0.242375f
C589 VTAIL.n12 VSUBS 1.60516f
C590 VTAIL.n13 VSUBS 0.878538f
C591 VTAIL.t19 VSUBS 0.242375f
C592 VTAIL.t1 VSUBS 0.242375f
C593 VTAIL.n14 VSUBS 1.60516f
C594 VTAIL.n15 VSUBS 0.856608f
C595 VTAIL.t7 VSUBS 2.15455f
C596 VTAIL.n16 VSUBS 2.27656f
C597 VTAIL.t9 VSUBS 2.15454f
C598 VTAIL.n17 VSUBS 2.27657f
C599 VTAIL.t14 VSUBS 0.242375f
C600 VTAIL.t15 VSUBS 0.242375f
C601 VTAIL.n18 VSUBS 1.60515f
C602 VTAIL.n19 VSUBS 0.806927f
C603 VDD2.t5 VSUBS 2.10036f
C604 VDD2.t8 VSUBS 0.217292f
C605 VDD2.t0 VSUBS 0.217292f
C606 VDD2.n0 VSUBS 1.58925f
C607 VDD2.n1 VSUBS 1.32381f
C608 VDD2.t6 VSUBS 0.217292f
C609 VDD2.t1 VSUBS 0.217292f
C610 VDD2.n2 VSUBS 1.59215f
C611 VDD2.n3 VSUBS 2.12407f
C612 VDD2.t9 VSUBS 2.09576f
C613 VDD2.n4 VSUBS 2.72826f
C614 VDD2.t3 VSUBS 0.217292f
C615 VDD2.t7 VSUBS 0.217292f
C616 VDD2.n5 VSUBS 1.58925f
C617 VDD2.n6 VSUBS 0.625435f
C618 VDD2.t2 VSUBS 0.217292f
C619 VDD2.t4 VSUBS 0.217292f
C620 VDD2.n7 VSUBS 1.59212f
C621 VN.n0 VSUBS 0.069316f
C622 VN.t2 VSUBS 0.520154f
C623 VN.t3 VSUBS 0.520154f
C624 VN.n1 VSUBS 0.028123f
C625 VN.t9 VSUBS 0.528647f
C626 VN.t0 VSUBS 0.520154f
C627 VN.n2 VSUBS 0.217412f
C628 VN.n3 VSUBS 0.238419f
C629 VN.n4 VSUBS 0.150077f
C630 VN.n5 VSUBS 0.069316f
C631 VN.n6 VSUBS 0.240406f
C632 VN.n7 VSUBS 0.028123f
C633 VN.n8 VSUBS 0.217412f
C634 VN.t8 VSUBS 0.528647f
C635 VN.n9 VSUBS 0.238324f
C636 VN.n10 VSUBS 0.053717f
C637 VN.n11 VSUBS 0.069316f
C638 VN.t4 VSUBS 0.528647f
C639 VN.t6 VSUBS 0.520154f
C640 VN.t1 VSUBS 0.520154f
C641 VN.n12 VSUBS 0.028123f
C642 VN.t5 VSUBS 0.520154f
C643 VN.n13 VSUBS 0.217412f
C644 VN.t7 VSUBS 0.528647f
C645 VN.n14 VSUBS 0.238419f
C646 VN.n15 VSUBS 0.150077f
C647 VN.n16 VSUBS 0.069316f
C648 VN.n17 VSUBS 0.240406f
C649 VN.n18 VSUBS 0.028123f
C650 VN.n19 VSUBS 0.217412f
C651 VN.n20 VSUBS 0.238324f
C652 VN.n21 VSUBS 2.49993f
.ends

