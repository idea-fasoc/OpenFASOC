* NGSPICE file created from diff_pair_sample_1384.ext - technology: sky130A

.subckt diff_pair_sample_1384 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t13 w_n3100_n4792# sky130_fd_pr__pfet_01v8 ad=3.1548 pd=19.45 as=7.4568 ps=39.02 w=19.12 l=1.8
X1 VDD2.t7 VN.t0 VTAIL.t5 w_n3100_n4792# sky130_fd_pr__pfet_01v8 ad=3.1548 pd=19.45 as=3.1548 ps=19.45 w=19.12 l=1.8
X2 VTAIL.t15 VP.t1 VDD1.t6 w_n3100_n4792# sky130_fd_pr__pfet_01v8 ad=7.4568 pd=39.02 as=3.1548 ps=19.45 w=19.12 l=1.8
X3 VTAIL.t1 VN.t1 VDD2.t6 w_n3100_n4792# sky130_fd_pr__pfet_01v8 ad=7.4568 pd=39.02 as=3.1548 ps=19.45 w=19.12 l=1.8
X4 B.t11 B.t9 B.t10 w_n3100_n4792# sky130_fd_pr__pfet_01v8 ad=7.4568 pd=39.02 as=0 ps=0 w=19.12 l=1.8
X5 B.t8 B.t6 B.t7 w_n3100_n4792# sky130_fd_pr__pfet_01v8 ad=7.4568 pd=39.02 as=0 ps=0 w=19.12 l=1.8
X6 VDD1.t5 VP.t2 VTAIL.t8 w_n3100_n4792# sky130_fd_pr__pfet_01v8 ad=3.1548 pd=19.45 as=7.4568 ps=39.02 w=19.12 l=1.8
X7 VDD2.t5 VN.t2 VTAIL.t0 w_n3100_n4792# sky130_fd_pr__pfet_01v8 ad=3.1548 pd=19.45 as=7.4568 ps=39.02 w=19.12 l=1.8
X8 B.t5 B.t3 B.t4 w_n3100_n4792# sky130_fd_pr__pfet_01v8 ad=7.4568 pd=39.02 as=0 ps=0 w=19.12 l=1.8
X9 VDD1.t4 VP.t3 VTAIL.t10 w_n3100_n4792# sky130_fd_pr__pfet_01v8 ad=3.1548 pd=19.45 as=3.1548 ps=19.45 w=19.12 l=1.8
X10 VDD2.t4 VN.t3 VTAIL.t4 w_n3100_n4792# sky130_fd_pr__pfet_01v8 ad=3.1548 pd=19.45 as=3.1548 ps=19.45 w=19.12 l=1.8
X11 VTAIL.t7 VN.t4 VDD2.t3 w_n3100_n4792# sky130_fd_pr__pfet_01v8 ad=3.1548 pd=19.45 as=3.1548 ps=19.45 w=19.12 l=1.8
X12 VTAIL.t9 VP.t4 VDD1.t3 w_n3100_n4792# sky130_fd_pr__pfet_01v8 ad=3.1548 pd=19.45 as=3.1548 ps=19.45 w=19.12 l=1.8
X13 VDD1.t2 VP.t5 VTAIL.t11 w_n3100_n4792# sky130_fd_pr__pfet_01v8 ad=3.1548 pd=19.45 as=3.1548 ps=19.45 w=19.12 l=1.8
X14 VTAIL.t12 VP.t6 VDD1.t1 w_n3100_n4792# sky130_fd_pr__pfet_01v8 ad=3.1548 pd=19.45 as=3.1548 ps=19.45 w=19.12 l=1.8
X15 VTAIL.t2 VN.t5 VDD2.t2 w_n3100_n4792# sky130_fd_pr__pfet_01v8 ad=3.1548 pd=19.45 as=3.1548 ps=19.45 w=19.12 l=1.8
X16 VTAIL.t6 VN.t6 VDD2.t1 w_n3100_n4792# sky130_fd_pr__pfet_01v8 ad=7.4568 pd=39.02 as=3.1548 ps=19.45 w=19.12 l=1.8
X17 VDD2.t0 VN.t7 VTAIL.t3 w_n3100_n4792# sky130_fd_pr__pfet_01v8 ad=3.1548 pd=19.45 as=7.4568 ps=39.02 w=19.12 l=1.8
X18 VTAIL.t14 VP.t7 VDD1.t0 w_n3100_n4792# sky130_fd_pr__pfet_01v8 ad=7.4568 pd=39.02 as=3.1548 ps=19.45 w=19.12 l=1.8
X19 B.t2 B.t0 B.t1 w_n3100_n4792# sky130_fd_pr__pfet_01v8 ad=7.4568 pd=39.02 as=0 ps=0 w=19.12 l=1.8
R0 VP.n10 VP.t1 287.122
R1 VP.n28 VP.t7 255.996
R2 VP.n35 VP.t5 255.996
R3 VP.n42 VP.t4 255.996
R4 VP.n49 VP.t2 255.996
R5 VP.n25 VP.t0 255.996
R6 VP.n18 VP.t6 255.996
R7 VP.n11 VP.t3 255.996
R8 VP.n13 VP.n12 161.3
R9 VP.n14 VP.n9 161.3
R10 VP.n16 VP.n15 161.3
R11 VP.n17 VP.n8 161.3
R12 VP.n20 VP.n19 161.3
R13 VP.n21 VP.n7 161.3
R14 VP.n23 VP.n22 161.3
R15 VP.n24 VP.n6 161.3
R16 VP.n48 VP.n0 161.3
R17 VP.n47 VP.n46 161.3
R18 VP.n45 VP.n1 161.3
R19 VP.n44 VP.n43 161.3
R20 VP.n41 VP.n2 161.3
R21 VP.n40 VP.n39 161.3
R22 VP.n38 VP.n3 161.3
R23 VP.n37 VP.n36 161.3
R24 VP.n34 VP.n4 161.3
R25 VP.n33 VP.n32 161.3
R26 VP.n31 VP.n5 161.3
R27 VP.n30 VP.n29 161.3
R28 VP.n28 VP.n27 89.0215
R29 VP.n50 VP.n49 89.0215
R30 VP.n26 VP.n25 89.0215
R31 VP.n40 VP.n3 56.5617
R32 VP.n16 VP.n9 56.5617
R33 VP.n11 VP.n10 54.4655
R34 VP.n27 VP.n26 52.5527
R35 VP.n33 VP.n5 52.2023
R36 VP.n47 VP.n1 52.2023
R37 VP.n23 VP.n7 52.2023
R38 VP.n29 VP.n5 28.9518
R39 VP.n48 VP.n47 28.9518
R40 VP.n24 VP.n23 28.9518
R41 VP.n34 VP.n33 24.5923
R42 VP.n36 VP.n3 24.5923
R43 VP.n41 VP.n40 24.5923
R44 VP.n43 VP.n1 24.5923
R45 VP.n17 VP.n16 24.5923
R46 VP.n19 VP.n7 24.5923
R47 VP.n12 VP.n9 24.5923
R48 VP.n29 VP.n28 21.8872
R49 VP.n49 VP.n48 21.8872
R50 VP.n25 VP.n24 21.8872
R51 VP.n36 VP.n35 15.4934
R52 VP.n42 VP.n41 15.4934
R53 VP.n18 VP.n17 15.4934
R54 VP.n12 VP.n11 15.4934
R55 VP.n13 VP.n10 12.9786
R56 VP.n35 VP.n34 9.09948
R57 VP.n43 VP.n42 9.09948
R58 VP.n19 VP.n18 9.09948
R59 VP.n26 VP.n6 0.278335
R60 VP.n30 VP.n27 0.278335
R61 VP.n50 VP.n0 0.278335
R62 VP.n14 VP.n13 0.189894
R63 VP.n15 VP.n14 0.189894
R64 VP.n15 VP.n8 0.189894
R65 VP.n20 VP.n8 0.189894
R66 VP.n21 VP.n20 0.189894
R67 VP.n22 VP.n21 0.189894
R68 VP.n22 VP.n6 0.189894
R69 VP.n31 VP.n30 0.189894
R70 VP.n32 VP.n31 0.189894
R71 VP.n32 VP.n4 0.189894
R72 VP.n37 VP.n4 0.189894
R73 VP.n38 VP.n37 0.189894
R74 VP.n39 VP.n38 0.189894
R75 VP.n39 VP.n2 0.189894
R76 VP.n44 VP.n2 0.189894
R77 VP.n45 VP.n44 0.189894
R78 VP.n46 VP.n45 0.189894
R79 VP.n46 VP.n0 0.189894
R80 VP VP.n50 0.153485
R81 VTAIL.n11 VTAIL.t15 56.0942
R82 VTAIL.n10 VTAIL.t0 56.0942
R83 VTAIL.n7 VTAIL.t6 56.0942
R84 VTAIL.n15 VTAIL.t3 56.0941
R85 VTAIL.n2 VTAIL.t1 56.0941
R86 VTAIL.n3 VTAIL.t8 56.0941
R87 VTAIL.n6 VTAIL.t14 56.0941
R88 VTAIL.n14 VTAIL.t13 56.0941
R89 VTAIL.n13 VTAIL.n12 54.3942
R90 VTAIL.n9 VTAIL.n8 54.3942
R91 VTAIL.n1 VTAIL.n0 54.393
R92 VTAIL.n5 VTAIL.n4 54.393
R93 VTAIL.n15 VTAIL.n14 30.6858
R94 VTAIL.n7 VTAIL.n6 30.6858
R95 VTAIL.n9 VTAIL.n7 1.83671
R96 VTAIL.n10 VTAIL.n9 1.83671
R97 VTAIL.n13 VTAIL.n11 1.83671
R98 VTAIL.n14 VTAIL.n13 1.83671
R99 VTAIL.n6 VTAIL.n5 1.83671
R100 VTAIL.n5 VTAIL.n3 1.83671
R101 VTAIL.n2 VTAIL.n1 1.83671
R102 VTAIL VTAIL.n15 1.77852
R103 VTAIL.n0 VTAIL.t4 1.70055
R104 VTAIL.n0 VTAIL.t7 1.70055
R105 VTAIL.n4 VTAIL.t11 1.70055
R106 VTAIL.n4 VTAIL.t9 1.70055
R107 VTAIL.n12 VTAIL.t10 1.70055
R108 VTAIL.n12 VTAIL.t12 1.70055
R109 VTAIL.n8 VTAIL.t5 1.70055
R110 VTAIL.n8 VTAIL.t2 1.70055
R111 VTAIL.n11 VTAIL.n10 0.470328
R112 VTAIL.n3 VTAIL.n2 0.470328
R113 VTAIL VTAIL.n1 0.0586897
R114 VDD1 VDD1.n0 72.0493
R115 VDD1.n3 VDD1.n2 71.9345
R116 VDD1.n3 VDD1.n1 71.9345
R117 VDD1.n5 VDD1.n4 71.0728
R118 VDD1.n5 VDD1.n3 49.044
R119 VDD1.n4 VDD1.t1 1.70055
R120 VDD1.n4 VDD1.t7 1.70055
R121 VDD1.n0 VDD1.t6 1.70055
R122 VDD1.n0 VDD1.t4 1.70055
R123 VDD1.n2 VDD1.t3 1.70055
R124 VDD1.n2 VDD1.t5 1.70055
R125 VDD1.n1 VDD1.t0 1.70055
R126 VDD1.n1 VDD1.t2 1.70055
R127 VDD1 VDD1.n5 0.860414
R128 VN.n4 VN.t1 287.122
R129 VN.n25 VN.t2 287.122
R130 VN.n5 VN.t3 255.996
R131 VN.n12 VN.t4 255.996
R132 VN.n19 VN.t7 255.996
R133 VN.n26 VN.t5 255.996
R134 VN.n33 VN.t0 255.996
R135 VN.n40 VN.t6 255.996
R136 VN.n39 VN.n21 161.3
R137 VN.n38 VN.n37 161.3
R138 VN.n36 VN.n22 161.3
R139 VN.n35 VN.n34 161.3
R140 VN.n32 VN.n23 161.3
R141 VN.n31 VN.n30 161.3
R142 VN.n29 VN.n24 161.3
R143 VN.n28 VN.n27 161.3
R144 VN.n18 VN.n0 161.3
R145 VN.n17 VN.n16 161.3
R146 VN.n15 VN.n1 161.3
R147 VN.n14 VN.n13 161.3
R148 VN.n11 VN.n2 161.3
R149 VN.n10 VN.n9 161.3
R150 VN.n8 VN.n3 161.3
R151 VN.n7 VN.n6 161.3
R152 VN.n20 VN.n19 89.0215
R153 VN.n41 VN.n40 89.0215
R154 VN.n10 VN.n3 56.5617
R155 VN.n31 VN.n24 56.5617
R156 VN.n5 VN.n4 54.4655
R157 VN.n26 VN.n25 54.4655
R158 VN VN.n41 52.8315
R159 VN.n17 VN.n1 52.2023
R160 VN.n38 VN.n22 52.2023
R161 VN.n18 VN.n17 28.9518
R162 VN.n39 VN.n38 28.9518
R163 VN.n6 VN.n3 24.5923
R164 VN.n11 VN.n10 24.5923
R165 VN.n13 VN.n1 24.5923
R166 VN.n27 VN.n24 24.5923
R167 VN.n34 VN.n22 24.5923
R168 VN.n32 VN.n31 24.5923
R169 VN.n19 VN.n18 21.8872
R170 VN.n40 VN.n39 21.8872
R171 VN.n6 VN.n5 15.4934
R172 VN.n12 VN.n11 15.4934
R173 VN.n27 VN.n26 15.4934
R174 VN.n33 VN.n32 15.4934
R175 VN.n28 VN.n25 12.9786
R176 VN.n7 VN.n4 12.9786
R177 VN.n13 VN.n12 9.09948
R178 VN.n34 VN.n33 9.09948
R179 VN.n41 VN.n21 0.278335
R180 VN.n20 VN.n0 0.278335
R181 VN.n37 VN.n21 0.189894
R182 VN.n37 VN.n36 0.189894
R183 VN.n36 VN.n35 0.189894
R184 VN.n35 VN.n23 0.189894
R185 VN.n30 VN.n23 0.189894
R186 VN.n30 VN.n29 0.189894
R187 VN.n29 VN.n28 0.189894
R188 VN.n8 VN.n7 0.189894
R189 VN.n9 VN.n8 0.189894
R190 VN.n9 VN.n2 0.189894
R191 VN.n14 VN.n2 0.189894
R192 VN.n15 VN.n14 0.189894
R193 VN.n16 VN.n15 0.189894
R194 VN.n16 VN.n0 0.189894
R195 VN VN.n20 0.153485
R196 VDD2.n2 VDD2.n1 71.9345
R197 VDD2.n2 VDD2.n0 71.9345
R198 VDD2 VDD2.n5 71.9327
R199 VDD2.n4 VDD2.n3 71.073
R200 VDD2.n4 VDD2.n2 48.461
R201 VDD2.n5 VDD2.t2 1.70055
R202 VDD2.n5 VDD2.t5 1.70055
R203 VDD2.n3 VDD2.t1 1.70055
R204 VDD2.n3 VDD2.t7 1.70055
R205 VDD2.n1 VDD2.t3 1.70055
R206 VDD2.n1 VDD2.t0 1.70055
R207 VDD2.n0 VDD2.t6 1.70055
R208 VDD2.n0 VDD2.t4 1.70055
R209 VDD2 VDD2.n4 0.976793
R210 B.n484 B.n133 585
R211 B.n483 B.n482 585
R212 B.n481 B.n134 585
R213 B.n480 B.n479 585
R214 B.n478 B.n135 585
R215 B.n477 B.n476 585
R216 B.n475 B.n136 585
R217 B.n474 B.n473 585
R218 B.n472 B.n137 585
R219 B.n471 B.n470 585
R220 B.n469 B.n138 585
R221 B.n468 B.n467 585
R222 B.n466 B.n139 585
R223 B.n465 B.n464 585
R224 B.n463 B.n140 585
R225 B.n462 B.n461 585
R226 B.n460 B.n141 585
R227 B.n459 B.n458 585
R228 B.n457 B.n142 585
R229 B.n456 B.n455 585
R230 B.n454 B.n143 585
R231 B.n453 B.n452 585
R232 B.n451 B.n144 585
R233 B.n450 B.n449 585
R234 B.n448 B.n145 585
R235 B.n447 B.n446 585
R236 B.n445 B.n146 585
R237 B.n444 B.n443 585
R238 B.n442 B.n147 585
R239 B.n441 B.n440 585
R240 B.n439 B.n148 585
R241 B.n438 B.n437 585
R242 B.n436 B.n149 585
R243 B.n435 B.n434 585
R244 B.n433 B.n150 585
R245 B.n432 B.n431 585
R246 B.n430 B.n151 585
R247 B.n429 B.n428 585
R248 B.n427 B.n152 585
R249 B.n426 B.n425 585
R250 B.n424 B.n153 585
R251 B.n423 B.n422 585
R252 B.n421 B.n154 585
R253 B.n420 B.n419 585
R254 B.n418 B.n155 585
R255 B.n417 B.n416 585
R256 B.n415 B.n156 585
R257 B.n414 B.n413 585
R258 B.n412 B.n157 585
R259 B.n411 B.n410 585
R260 B.n409 B.n158 585
R261 B.n408 B.n407 585
R262 B.n406 B.n159 585
R263 B.n405 B.n404 585
R264 B.n403 B.n160 585
R265 B.n402 B.n401 585
R266 B.n400 B.n161 585
R267 B.n399 B.n398 585
R268 B.n397 B.n162 585
R269 B.n396 B.n395 585
R270 B.n394 B.n163 585
R271 B.n393 B.n392 585
R272 B.n391 B.n164 585
R273 B.n390 B.n389 585
R274 B.n385 B.n165 585
R275 B.n384 B.n383 585
R276 B.n382 B.n166 585
R277 B.n381 B.n380 585
R278 B.n379 B.n167 585
R279 B.n378 B.n377 585
R280 B.n376 B.n168 585
R281 B.n375 B.n374 585
R282 B.n372 B.n169 585
R283 B.n371 B.n370 585
R284 B.n369 B.n172 585
R285 B.n368 B.n367 585
R286 B.n366 B.n173 585
R287 B.n365 B.n364 585
R288 B.n363 B.n174 585
R289 B.n362 B.n361 585
R290 B.n360 B.n175 585
R291 B.n359 B.n358 585
R292 B.n357 B.n176 585
R293 B.n356 B.n355 585
R294 B.n354 B.n177 585
R295 B.n353 B.n352 585
R296 B.n351 B.n178 585
R297 B.n350 B.n349 585
R298 B.n348 B.n179 585
R299 B.n347 B.n346 585
R300 B.n345 B.n180 585
R301 B.n344 B.n343 585
R302 B.n342 B.n181 585
R303 B.n341 B.n340 585
R304 B.n339 B.n182 585
R305 B.n338 B.n337 585
R306 B.n336 B.n183 585
R307 B.n335 B.n334 585
R308 B.n333 B.n184 585
R309 B.n332 B.n331 585
R310 B.n330 B.n185 585
R311 B.n329 B.n328 585
R312 B.n327 B.n186 585
R313 B.n326 B.n325 585
R314 B.n324 B.n187 585
R315 B.n323 B.n322 585
R316 B.n321 B.n188 585
R317 B.n320 B.n319 585
R318 B.n318 B.n189 585
R319 B.n317 B.n316 585
R320 B.n315 B.n190 585
R321 B.n314 B.n313 585
R322 B.n312 B.n191 585
R323 B.n311 B.n310 585
R324 B.n309 B.n192 585
R325 B.n308 B.n307 585
R326 B.n306 B.n193 585
R327 B.n305 B.n304 585
R328 B.n303 B.n194 585
R329 B.n302 B.n301 585
R330 B.n300 B.n195 585
R331 B.n299 B.n298 585
R332 B.n297 B.n196 585
R333 B.n296 B.n295 585
R334 B.n294 B.n197 585
R335 B.n293 B.n292 585
R336 B.n291 B.n198 585
R337 B.n290 B.n289 585
R338 B.n288 B.n199 585
R339 B.n287 B.n286 585
R340 B.n285 B.n200 585
R341 B.n284 B.n283 585
R342 B.n282 B.n201 585
R343 B.n281 B.n280 585
R344 B.n279 B.n202 585
R345 B.n486 B.n485 585
R346 B.n487 B.n132 585
R347 B.n489 B.n488 585
R348 B.n490 B.n131 585
R349 B.n492 B.n491 585
R350 B.n493 B.n130 585
R351 B.n495 B.n494 585
R352 B.n496 B.n129 585
R353 B.n498 B.n497 585
R354 B.n499 B.n128 585
R355 B.n501 B.n500 585
R356 B.n502 B.n127 585
R357 B.n504 B.n503 585
R358 B.n505 B.n126 585
R359 B.n507 B.n506 585
R360 B.n508 B.n125 585
R361 B.n510 B.n509 585
R362 B.n511 B.n124 585
R363 B.n513 B.n512 585
R364 B.n514 B.n123 585
R365 B.n516 B.n515 585
R366 B.n517 B.n122 585
R367 B.n519 B.n518 585
R368 B.n520 B.n121 585
R369 B.n522 B.n521 585
R370 B.n523 B.n120 585
R371 B.n525 B.n524 585
R372 B.n526 B.n119 585
R373 B.n528 B.n527 585
R374 B.n529 B.n118 585
R375 B.n531 B.n530 585
R376 B.n532 B.n117 585
R377 B.n534 B.n533 585
R378 B.n535 B.n116 585
R379 B.n537 B.n536 585
R380 B.n538 B.n115 585
R381 B.n540 B.n539 585
R382 B.n541 B.n114 585
R383 B.n543 B.n542 585
R384 B.n544 B.n113 585
R385 B.n546 B.n545 585
R386 B.n547 B.n112 585
R387 B.n549 B.n548 585
R388 B.n550 B.n111 585
R389 B.n552 B.n551 585
R390 B.n553 B.n110 585
R391 B.n555 B.n554 585
R392 B.n556 B.n109 585
R393 B.n558 B.n557 585
R394 B.n559 B.n108 585
R395 B.n561 B.n560 585
R396 B.n562 B.n107 585
R397 B.n564 B.n563 585
R398 B.n565 B.n106 585
R399 B.n567 B.n566 585
R400 B.n568 B.n105 585
R401 B.n570 B.n569 585
R402 B.n571 B.n104 585
R403 B.n573 B.n572 585
R404 B.n574 B.n103 585
R405 B.n576 B.n575 585
R406 B.n577 B.n102 585
R407 B.n579 B.n578 585
R408 B.n580 B.n101 585
R409 B.n582 B.n581 585
R410 B.n583 B.n100 585
R411 B.n585 B.n584 585
R412 B.n586 B.n99 585
R413 B.n588 B.n587 585
R414 B.n589 B.n98 585
R415 B.n591 B.n590 585
R416 B.n592 B.n97 585
R417 B.n594 B.n593 585
R418 B.n595 B.n96 585
R419 B.n597 B.n596 585
R420 B.n598 B.n95 585
R421 B.n600 B.n599 585
R422 B.n601 B.n94 585
R423 B.n603 B.n602 585
R424 B.n604 B.n93 585
R425 B.n809 B.n808 585
R426 B.n807 B.n22 585
R427 B.n806 B.n805 585
R428 B.n804 B.n23 585
R429 B.n803 B.n802 585
R430 B.n801 B.n24 585
R431 B.n800 B.n799 585
R432 B.n798 B.n25 585
R433 B.n797 B.n796 585
R434 B.n795 B.n26 585
R435 B.n794 B.n793 585
R436 B.n792 B.n27 585
R437 B.n791 B.n790 585
R438 B.n789 B.n28 585
R439 B.n788 B.n787 585
R440 B.n786 B.n29 585
R441 B.n785 B.n784 585
R442 B.n783 B.n30 585
R443 B.n782 B.n781 585
R444 B.n780 B.n31 585
R445 B.n779 B.n778 585
R446 B.n777 B.n32 585
R447 B.n776 B.n775 585
R448 B.n774 B.n33 585
R449 B.n773 B.n772 585
R450 B.n771 B.n34 585
R451 B.n770 B.n769 585
R452 B.n768 B.n35 585
R453 B.n767 B.n766 585
R454 B.n765 B.n36 585
R455 B.n764 B.n763 585
R456 B.n762 B.n37 585
R457 B.n761 B.n760 585
R458 B.n759 B.n38 585
R459 B.n758 B.n757 585
R460 B.n756 B.n39 585
R461 B.n755 B.n754 585
R462 B.n753 B.n40 585
R463 B.n752 B.n751 585
R464 B.n750 B.n41 585
R465 B.n749 B.n748 585
R466 B.n747 B.n42 585
R467 B.n746 B.n745 585
R468 B.n744 B.n43 585
R469 B.n743 B.n742 585
R470 B.n741 B.n44 585
R471 B.n740 B.n739 585
R472 B.n738 B.n45 585
R473 B.n737 B.n736 585
R474 B.n735 B.n46 585
R475 B.n734 B.n733 585
R476 B.n732 B.n47 585
R477 B.n731 B.n730 585
R478 B.n729 B.n48 585
R479 B.n728 B.n727 585
R480 B.n726 B.n49 585
R481 B.n725 B.n724 585
R482 B.n723 B.n50 585
R483 B.n722 B.n721 585
R484 B.n720 B.n51 585
R485 B.n719 B.n718 585
R486 B.n717 B.n52 585
R487 B.n716 B.n715 585
R488 B.n713 B.n53 585
R489 B.n712 B.n711 585
R490 B.n710 B.n56 585
R491 B.n709 B.n708 585
R492 B.n707 B.n57 585
R493 B.n706 B.n705 585
R494 B.n704 B.n58 585
R495 B.n703 B.n702 585
R496 B.n701 B.n59 585
R497 B.n699 B.n698 585
R498 B.n697 B.n62 585
R499 B.n696 B.n695 585
R500 B.n694 B.n63 585
R501 B.n693 B.n692 585
R502 B.n691 B.n64 585
R503 B.n690 B.n689 585
R504 B.n688 B.n65 585
R505 B.n687 B.n686 585
R506 B.n685 B.n66 585
R507 B.n684 B.n683 585
R508 B.n682 B.n67 585
R509 B.n681 B.n680 585
R510 B.n679 B.n68 585
R511 B.n678 B.n677 585
R512 B.n676 B.n69 585
R513 B.n675 B.n674 585
R514 B.n673 B.n70 585
R515 B.n672 B.n671 585
R516 B.n670 B.n71 585
R517 B.n669 B.n668 585
R518 B.n667 B.n72 585
R519 B.n666 B.n665 585
R520 B.n664 B.n73 585
R521 B.n663 B.n662 585
R522 B.n661 B.n74 585
R523 B.n660 B.n659 585
R524 B.n658 B.n75 585
R525 B.n657 B.n656 585
R526 B.n655 B.n76 585
R527 B.n654 B.n653 585
R528 B.n652 B.n77 585
R529 B.n651 B.n650 585
R530 B.n649 B.n78 585
R531 B.n648 B.n647 585
R532 B.n646 B.n79 585
R533 B.n645 B.n644 585
R534 B.n643 B.n80 585
R535 B.n642 B.n641 585
R536 B.n640 B.n81 585
R537 B.n639 B.n638 585
R538 B.n637 B.n82 585
R539 B.n636 B.n635 585
R540 B.n634 B.n83 585
R541 B.n633 B.n632 585
R542 B.n631 B.n84 585
R543 B.n630 B.n629 585
R544 B.n628 B.n85 585
R545 B.n627 B.n626 585
R546 B.n625 B.n86 585
R547 B.n624 B.n623 585
R548 B.n622 B.n87 585
R549 B.n621 B.n620 585
R550 B.n619 B.n88 585
R551 B.n618 B.n617 585
R552 B.n616 B.n89 585
R553 B.n615 B.n614 585
R554 B.n613 B.n90 585
R555 B.n612 B.n611 585
R556 B.n610 B.n91 585
R557 B.n609 B.n608 585
R558 B.n607 B.n92 585
R559 B.n606 B.n605 585
R560 B.n810 B.n21 585
R561 B.n812 B.n811 585
R562 B.n813 B.n20 585
R563 B.n815 B.n814 585
R564 B.n816 B.n19 585
R565 B.n818 B.n817 585
R566 B.n819 B.n18 585
R567 B.n821 B.n820 585
R568 B.n822 B.n17 585
R569 B.n824 B.n823 585
R570 B.n825 B.n16 585
R571 B.n827 B.n826 585
R572 B.n828 B.n15 585
R573 B.n830 B.n829 585
R574 B.n831 B.n14 585
R575 B.n833 B.n832 585
R576 B.n834 B.n13 585
R577 B.n836 B.n835 585
R578 B.n837 B.n12 585
R579 B.n839 B.n838 585
R580 B.n840 B.n11 585
R581 B.n842 B.n841 585
R582 B.n843 B.n10 585
R583 B.n845 B.n844 585
R584 B.n846 B.n9 585
R585 B.n848 B.n847 585
R586 B.n849 B.n8 585
R587 B.n851 B.n850 585
R588 B.n852 B.n7 585
R589 B.n854 B.n853 585
R590 B.n855 B.n6 585
R591 B.n857 B.n856 585
R592 B.n858 B.n5 585
R593 B.n860 B.n859 585
R594 B.n861 B.n4 585
R595 B.n863 B.n862 585
R596 B.n864 B.n3 585
R597 B.n866 B.n865 585
R598 B.n867 B.n0 585
R599 B.n2 B.n1 585
R600 B.n222 B.n221 585
R601 B.n224 B.n223 585
R602 B.n225 B.n220 585
R603 B.n227 B.n226 585
R604 B.n228 B.n219 585
R605 B.n230 B.n229 585
R606 B.n231 B.n218 585
R607 B.n233 B.n232 585
R608 B.n234 B.n217 585
R609 B.n236 B.n235 585
R610 B.n237 B.n216 585
R611 B.n239 B.n238 585
R612 B.n240 B.n215 585
R613 B.n242 B.n241 585
R614 B.n243 B.n214 585
R615 B.n245 B.n244 585
R616 B.n246 B.n213 585
R617 B.n248 B.n247 585
R618 B.n249 B.n212 585
R619 B.n251 B.n250 585
R620 B.n252 B.n211 585
R621 B.n254 B.n253 585
R622 B.n255 B.n210 585
R623 B.n257 B.n256 585
R624 B.n258 B.n209 585
R625 B.n260 B.n259 585
R626 B.n261 B.n208 585
R627 B.n263 B.n262 585
R628 B.n264 B.n207 585
R629 B.n266 B.n265 585
R630 B.n267 B.n206 585
R631 B.n269 B.n268 585
R632 B.n270 B.n205 585
R633 B.n272 B.n271 585
R634 B.n273 B.n204 585
R635 B.n275 B.n274 585
R636 B.n276 B.n203 585
R637 B.n278 B.n277 585
R638 B.n279 B.n278 463.671
R639 B.n486 B.n133 463.671
R640 B.n606 B.n93 463.671
R641 B.n808 B.n21 463.671
R642 B.n170 B.t0 462.401
R643 B.n386 B.t6 462.401
R644 B.n60 B.t9 462.401
R645 B.n54 B.t3 462.401
R646 B.n869 B.n868 256.663
R647 B.n868 B.n867 235.042
R648 B.n868 B.n2 235.042
R649 B.n280 B.n279 163.367
R650 B.n280 B.n201 163.367
R651 B.n284 B.n201 163.367
R652 B.n285 B.n284 163.367
R653 B.n286 B.n285 163.367
R654 B.n286 B.n199 163.367
R655 B.n290 B.n199 163.367
R656 B.n291 B.n290 163.367
R657 B.n292 B.n291 163.367
R658 B.n292 B.n197 163.367
R659 B.n296 B.n197 163.367
R660 B.n297 B.n296 163.367
R661 B.n298 B.n297 163.367
R662 B.n298 B.n195 163.367
R663 B.n302 B.n195 163.367
R664 B.n303 B.n302 163.367
R665 B.n304 B.n303 163.367
R666 B.n304 B.n193 163.367
R667 B.n308 B.n193 163.367
R668 B.n309 B.n308 163.367
R669 B.n310 B.n309 163.367
R670 B.n310 B.n191 163.367
R671 B.n314 B.n191 163.367
R672 B.n315 B.n314 163.367
R673 B.n316 B.n315 163.367
R674 B.n316 B.n189 163.367
R675 B.n320 B.n189 163.367
R676 B.n321 B.n320 163.367
R677 B.n322 B.n321 163.367
R678 B.n322 B.n187 163.367
R679 B.n326 B.n187 163.367
R680 B.n327 B.n326 163.367
R681 B.n328 B.n327 163.367
R682 B.n328 B.n185 163.367
R683 B.n332 B.n185 163.367
R684 B.n333 B.n332 163.367
R685 B.n334 B.n333 163.367
R686 B.n334 B.n183 163.367
R687 B.n338 B.n183 163.367
R688 B.n339 B.n338 163.367
R689 B.n340 B.n339 163.367
R690 B.n340 B.n181 163.367
R691 B.n344 B.n181 163.367
R692 B.n345 B.n344 163.367
R693 B.n346 B.n345 163.367
R694 B.n346 B.n179 163.367
R695 B.n350 B.n179 163.367
R696 B.n351 B.n350 163.367
R697 B.n352 B.n351 163.367
R698 B.n352 B.n177 163.367
R699 B.n356 B.n177 163.367
R700 B.n357 B.n356 163.367
R701 B.n358 B.n357 163.367
R702 B.n358 B.n175 163.367
R703 B.n362 B.n175 163.367
R704 B.n363 B.n362 163.367
R705 B.n364 B.n363 163.367
R706 B.n364 B.n173 163.367
R707 B.n368 B.n173 163.367
R708 B.n369 B.n368 163.367
R709 B.n370 B.n369 163.367
R710 B.n370 B.n169 163.367
R711 B.n375 B.n169 163.367
R712 B.n376 B.n375 163.367
R713 B.n377 B.n376 163.367
R714 B.n377 B.n167 163.367
R715 B.n381 B.n167 163.367
R716 B.n382 B.n381 163.367
R717 B.n383 B.n382 163.367
R718 B.n383 B.n165 163.367
R719 B.n390 B.n165 163.367
R720 B.n391 B.n390 163.367
R721 B.n392 B.n391 163.367
R722 B.n392 B.n163 163.367
R723 B.n396 B.n163 163.367
R724 B.n397 B.n396 163.367
R725 B.n398 B.n397 163.367
R726 B.n398 B.n161 163.367
R727 B.n402 B.n161 163.367
R728 B.n403 B.n402 163.367
R729 B.n404 B.n403 163.367
R730 B.n404 B.n159 163.367
R731 B.n408 B.n159 163.367
R732 B.n409 B.n408 163.367
R733 B.n410 B.n409 163.367
R734 B.n410 B.n157 163.367
R735 B.n414 B.n157 163.367
R736 B.n415 B.n414 163.367
R737 B.n416 B.n415 163.367
R738 B.n416 B.n155 163.367
R739 B.n420 B.n155 163.367
R740 B.n421 B.n420 163.367
R741 B.n422 B.n421 163.367
R742 B.n422 B.n153 163.367
R743 B.n426 B.n153 163.367
R744 B.n427 B.n426 163.367
R745 B.n428 B.n427 163.367
R746 B.n428 B.n151 163.367
R747 B.n432 B.n151 163.367
R748 B.n433 B.n432 163.367
R749 B.n434 B.n433 163.367
R750 B.n434 B.n149 163.367
R751 B.n438 B.n149 163.367
R752 B.n439 B.n438 163.367
R753 B.n440 B.n439 163.367
R754 B.n440 B.n147 163.367
R755 B.n444 B.n147 163.367
R756 B.n445 B.n444 163.367
R757 B.n446 B.n445 163.367
R758 B.n446 B.n145 163.367
R759 B.n450 B.n145 163.367
R760 B.n451 B.n450 163.367
R761 B.n452 B.n451 163.367
R762 B.n452 B.n143 163.367
R763 B.n456 B.n143 163.367
R764 B.n457 B.n456 163.367
R765 B.n458 B.n457 163.367
R766 B.n458 B.n141 163.367
R767 B.n462 B.n141 163.367
R768 B.n463 B.n462 163.367
R769 B.n464 B.n463 163.367
R770 B.n464 B.n139 163.367
R771 B.n468 B.n139 163.367
R772 B.n469 B.n468 163.367
R773 B.n470 B.n469 163.367
R774 B.n470 B.n137 163.367
R775 B.n474 B.n137 163.367
R776 B.n475 B.n474 163.367
R777 B.n476 B.n475 163.367
R778 B.n476 B.n135 163.367
R779 B.n480 B.n135 163.367
R780 B.n481 B.n480 163.367
R781 B.n482 B.n481 163.367
R782 B.n482 B.n133 163.367
R783 B.n602 B.n93 163.367
R784 B.n602 B.n601 163.367
R785 B.n601 B.n600 163.367
R786 B.n600 B.n95 163.367
R787 B.n596 B.n95 163.367
R788 B.n596 B.n595 163.367
R789 B.n595 B.n594 163.367
R790 B.n594 B.n97 163.367
R791 B.n590 B.n97 163.367
R792 B.n590 B.n589 163.367
R793 B.n589 B.n588 163.367
R794 B.n588 B.n99 163.367
R795 B.n584 B.n99 163.367
R796 B.n584 B.n583 163.367
R797 B.n583 B.n582 163.367
R798 B.n582 B.n101 163.367
R799 B.n578 B.n101 163.367
R800 B.n578 B.n577 163.367
R801 B.n577 B.n576 163.367
R802 B.n576 B.n103 163.367
R803 B.n572 B.n103 163.367
R804 B.n572 B.n571 163.367
R805 B.n571 B.n570 163.367
R806 B.n570 B.n105 163.367
R807 B.n566 B.n105 163.367
R808 B.n566 B.n565 163.367
R809 B.n565 B.n564 163.367
R810 B.n564 B.n107 163.367
R811 B.n560 B.n107 163.367
R812 B.n560 B.n559 163.367
R813 B.n559 B.n558 163.367
R814 B.n558 B.n109 163.367
R815 B.n554 B.n109 163.367
R816 B.n554 B.n553 163.367
R817 B.n553 B.n552 163.367
R818 B.n552 B.n111 163.367
R819 B.n548 B.n111 163.367
R820 B.n548 B.n547 163.367
R821 B.n547 B.n546 163.367
R822 B.n546 B.n113 163.367
R823 B.n542 B.n113 163.367
R824 B.n542 B.n541 163.367
R825 B.n541 B.n540 163.367
R826 B.n540 B.n115 163.367
R827 B.n536 B.n115 163.367
R828 B.n536 B.n535 163.367
R829 B.n535 B.n534 163.367
R830 B.n534 B.n117 163.367
R831 B.n530 B.n117 163.367
R832 B.n530 B.n529 163.367
R833 B.n529 B.n528 163.367
R834 B.n528 B.n119 163.367
R835 B.n524 B.n119 163.367
R836 B.n524 B.n523 163.367
R837 B.n523 B.n522 163.367
R838 B.n522 B.n121 163.367
R839 B.n518 B.n121 163.367
R840 B.n518 B.n517 163.367
R841 B.n517 B.n516 163.367
R842 B.n516 B.n123 163.367
R843 B.n512 B.n123 163.367
R844 B.n512 B.n511 163.367
R845 B.n511 B.n510 163.367
R846 B.n510 B.n125 163.367
R847 B.n506 B.n125 163.367
R848 B.n506 B.n505 163.367
R849 B.n505 B.n504 163.367
R850 B.n504 B.n127 163.367
R851 B.n500 B.n127 163.367
R852 B.n500 B.n499 163.367
R853 B.n499 B.n498 163.367
R854 B.n498 B.n129 163.367
R855 B.n494 B.n129 163.367
R856 B.n494 B.n493 163.367
R857 B.n493 B.n492 163.367
R858 B.n492 B.n131 163.367
R859 B.n488 B.n131 163.367
R860 B.n488 B.n487 163.367
R861 B.n487 B.n486 163.367
R862 B.n808 B.n807 163.367
R863 B.n807 B.n806 163.367
R864 B.n806 B.n23 163.367
R865 B.n802 B.n23 163.367
R866 B.n802 B.n801 163.367
R867 B.n801 B.n800 163.367
R868 B.n800 B.n25 163.367
R869 B.n796 B.n25 163.367
R870 B.n796 B.n795 163.367
R871 B.n795 B.n794 163.367
R872 B.n794 B.n27 163.367
R873 B.n790 B.n27 163.367
R874 B.n790 B.n789 163.367
R875 B.n789 B.n788 163.367
R876 B.n788 B.n29 163.367
R877 B.n784 B.n29 163.367
R878 B.n784 B.n783 163.367
R879 B.n783 B.n782 163.367
R880 B.n782 B.n31 163.367
R881 B.n778 B.n31 163.367
R882 B.n778 B.n777 163.367
R883 B.n777 B.n776 163.367
R884 B.n776 B.n33 163.367
R885 B.n772 B.n33 163.367
R886 B.n772 B.n771 163.367
R887 B.n771 B.n770 163.367
R888 B.n770 B.n35 163.367
R889 B.n766 B.n35 163.367
R890 B.n766 B.n765 163.367
R891 B.n765 B.n764 163.367
R892 B.n764 B.n37 163.367
R893 B.n760 B.n37 163.367
R894 B.n760 B.n759 163.367
R895 B.n759 B.n758 163.367
R896 B.n758 B.n39 163.367
R897 B.n754 B.n39 163.367
R898 B.n754 B.n753 163.367
R899 B.n753 B.n752 163.367
R900 B.n752 B.n41 163.367
R901 B.n748 B.n41 163.367
R902 B.n748 B.n747 163.367
R903 B.n747 B.n746 163.367
R904 B.n746 B.n43 163.367
R905 B.n742 B.n43 163.367
R906 B.n742 B.n741 163.367
R907 B.n741 B.n740 163.367
R908 B.n740 B.n45 163.367
R909 B.n736 B.n45 163.367
R910 B.n736 B.n735 163.367
R911 B.n735 B.n734 163.367
R912 B.n734 B.n47 163.367
R913 B.n730 B.n47 163.367
R914 B.n730 B.n729 163.367
R915 B.n729 B.n728 163.367
R916 B.n728 B.n49 163.367
R917 B.n724 B.n49 163.367
R918 B.n724 B.n723 163.367
R919 B.n723 B.n722 163.367
R920 B.n722 B.n51 163.367
R921 B.n718 B.n51 163.367
R922 B.n718 B.n717 163.367
R923 B.n717 B.n716 163.367
R924 B.n716 B.n53 163.367
R925 B.n711 B.n53 163.367
R926 B.n711 B.n710 163.367
R927 B.n710 B.n709 163.367
R928 B.n709 B.n57 163.367
R929 B.n705 B.n57 163.367
R930 B.n705 B.n704 163.367
R931 B.n704 B.n703 163.367
R932 B.n703 B.n59 163.367
R933 B.n698 B.n59 163.367
R934 B.n698 B.n697 163.367
R935 B.n697 B.n696 163.367
R936 B.n696 B.n63 163.367
R937 B.n692 B.n63 163.367
R938 B.n692 B.n691 163.367
R939 B.n691 B.n690 163.367
R940 B.n690 B.n65 163.367
R941 B.n686 B.n65 163.367
R942 B.n686 B.n685 163.367
R943 B.n685 B.n684 163.367
R944 B.n684 B.n67 163.367
R945 B.n680 B.n67 163.367
R946 B.n680 B.n679 163.367
R947 B.n679 B.n678 163.367
R948 B.n678 B.n69 163.367
R949 B.n674 B.n69 163.367
R950 B.n674 B.n673 163.367
R951 B.n673 B.n672 163.367
R952 B.n672 B.n71 163.367
R953 B.n668 B.n71 163.367
R954 B.n668 B.n667 163.367
R955 B.n667 B.n666 163.367
R956 B.n666 B.n73 163.367
R957 B.n662 B.n73 163.367
R958 B.n662 B.n661 163.367
R959 B.n661 B.n660 163.367
R960 B.n660 B.n75 163.367
R961 B.n656 B.n75 163.367
R962 B.n656 B.n655 163.367
R963 B.n655 B.n654 163.367
R964 B.n654 B.n77 163.367
R965 B.n650 B.n77 163.367
R966 B.n650 B.n649 163.367
R967 B.n649 B.n648 163.367
R968 B.n648 B.n79 163.367
R969 B.n644 B.n79 163.367
R970 B.n644 B.n643 163.367
R971 B.n643 B.n642 163.367
R972 B.n642 B.n81 163.367
R973 B.n638 B.n81 163.367
R974 B.n638 B.n637 163.367
R975 B.n637 B.n636 163.367
R976 B.n636 B.n83 163.367
R977 B.n632 B.n83 163.367
R978 B.n632 B.n631 163.367
R979 B.n631 B.n630 163.367
R980 B.n630 B.n85 163.367
R981 B.n626 B.n85 163.367
R982 B.n626 B.n625 163.367
R983 B.n625 B.n624 163.367
R984 B.n624 B.n87 163.367
R985 B.n620 B.n87 163.367
R986 B.n620 B.n619 163.367
R987 B.n619 B.n618 163.367
R988 B.n618 B.n89 163.367
R989 B.n614 B.n89 163.367
R990 B.n614 B.n613 163.367
R991 B.n613 B.n612 163.367
R992 B.n612 B.n91 163.367
R993 B.n608 B.n91 163.367
R994 B.n608 B.n607 163.367
R995 B.n607 B.n606 163.367
R996 B.n812 B.n21 163.367
R997 B.n813 B.n812 163.367
R998 B.n814 B.n813 163.367
R999 B.n814 B.n19 163.367
R1000 B.n818 B.n19 163.367
R1001 B.n819 B.n818 163.367
R1002 B.n820 B.n819 163.367
R1003 B.n820 B.n17 163.367
R1004 B.n824 B.n17 163.367
R1005 B.n825 B.n824 163.367
R1006 B.n826 B.n825 163.367
R1007 B.n826 B.n15 163.367
R1008 B.n830 B.n15 163.367
R1009 B.n831 B.n830 163.367
R1010 B.n832 B.n831 163.367
R1011 B.n832 B.n13 163.367
R1012 B.n836 B.n13 163.367
R1013 B.n837 B.n836 163.367
R1014 B.n838 B.n837 163.367
R1015 B.n838 B.n11 163.367
R1016 B.n842 B.n11 163.367
R1017 B.n843 B.n842 163.367
R1018 B.n844 B.n843 163.367
R1019 B.n844 B.n9 163.367
R1020 B.n848 B.n9 163.367
R1021 B.n849 B.n848 163.367
R1022 B.n850 B.n849 163.367
R1023 B.n850 B.n7 163.367
R1024 B.n854 B.n7 163.367
R1025 B.n855 B.n854 163.367
R1026 B.n856 B.n855 163.367
R1027 B.n856 B.n5 163.367
R1028 B.n860 B.n5 163.367
R1029 B.n861 B.n860 163.367
R1030 B.n862 B.n861 163.367
R1031 B.n862 B.n3 163.367
R1032 B.n866 B.n3 163.367
R1033 B.n867 B.n866 163.367
R1034 B.n221 B.n2 163.367
R1035 B.n224 B.n221 163.367
R1036 B.n225 B.n224 163.367
R1037 B.n226 B.n225 163.367
R1038 B.n226 B.n219 163.367
R1039 B.n230 B.n219 163.367
R1040 B.n231 B.n230 163.367
R1041 B.n232 B.n231 163.367
R1042 B.n232 B.n217 163.367
R1043 B.n236 B.n217 163.367
R1044 B.n237 B.n236 163.367
R1045 B.n238 B.n237 163.367
R1046 B.n238 B.n215 163.367
R1047 B.n242 B.n215 163.367
R1048 B.n243 B.n242 163.367
R1049 B.n244 B.n243 163.367
R1050 B.n244 B.n213 163.367
R1051 B.n248 B.n213 163.367
R1052 B.n249 B.n248 163.367
R1053 B.n250 B.n249 163.367
R1054 B.n250 B.n211 163.367
R1055 B.n254 B.n211 163.367
R1056 B.n255 B.n254 163.367
R1057 B.n256 B.n255 163.367
R1058 B.n256 B.n209 163.367
R1059 B.n260 B.n209 163.367
R1060 B.n261 B.n260 163.367
R1061 B.n262 B.n261 163.367
R1062 B.n262 B.n207 163.367
R1063 B.n266 B.n207 163.367
R1064 B.n267 B.n266 163.367
R1065 B.n268 B.n267 163.367
R1066 B.n268 B.n205 163.367
R1067 B.n272 B.n205 163.367
R1068 B.n273 B.n272 163.367
R1069 B.n274 B.n273 163.367
R1070 B.n274 B.n203 163.367
R1071 B.n278 B.n203 163.367
R1072 B.n386 B.t7 148.96
R1073 B.n60 B.t11 148.96
R1074 B.n170 B.t1 148.935
R1075 B.n54 B.t5 148.935
R1076 B.n387 B.t8 107.651
R1077 B.n61 B.t10 107.651
R1078 B.n171 B.t2 107.626
R1079 B.n55 B.t4 107.626
R1080 B.n373 B.n171 59.5399
R1081 B.n388 B.n387 59.5399
R1082 B.n700 B.n61 59.5399
R1083 B.n714 B.n55 59.5399
R1084 B.n171 B.n170 41.3096
R1085 B.n387 B.n386 41.3096
R1086 B.n61 B.n60 41.3096
R1087 B.n55 B.n54 41.3096
R1088 B.n810 B.n809 30.1273
R1089 B.n605 B.n604 30.1273
R1090 B.n485 B.n484 30.1273
R1091 B.n277 B.n202 30.1273
R1092 B B.n869 18.0485
R1093 B.n811 B.n810 10.6151
R1094 B.n811 B.n20 10.6151
R1095 B.n815 B.n20 10.6151
R1096 B.n816 B.n815 10.6151
R1097 B.n817 B.n816 10.6151
R1098 B.n817 B.n18 10.6151
R1099 B.n821 B.n18 10.6151
R1100 B.n822 B.n821 10.6151
R1101 B.n823 B.n822 10.6151
R1102 B.n823 B.n16 10.6151
R1103 B.n827 B.n16 10.6151
R1104 B.n828 B.n827 10.6151
R1105 B.n829 B.n828 10.6151
R1106 B.n829 B.n14 10.6151
R1107 B.n833 B.n14 10.6151
R1108 B.n834 B.n833 10.6151
R1109 B.n835 B.n834 10.6151
R1110 B.n835 B.n12 10.6151
R1111 B.n839 B.n12 10.6151
R1112 B.n840 B.n839 10.6151
R1113 B.n841 B.n840 10.6151
R1114 B.n841 B.n10 10.6151
R1115 B.n845 B.n10 10.6151
R1116 B.n846 B.n845 10.6151
R1117 B.n847 B.n846 10.6151
R1118 B.n847 B.n8 10.6151
R1119 B.n851 B.n8 10.6151
R1120 B.n852 B.n851 10.6151
R1121 B.n853 B.n852 10.6151
R1122 B.n853 B.n6 10.6151
R1123 B.n857 B.n6 10.6151
R1124 B.n858 B.n857 10.6151
R1125 B.n859 B.n858 10.6151
R1126 B.n859 B.n4 10.6151
R1127 B.n863 B.n4 10.6151
R1128 B.n864 B.n863 10.6151
R1129 B.n865 B.n864 10.6151
R1130 B.n865 B.n0 10.6151
R1131 B.n809 B.n22 10.6151
R1132 B.n805 B.n22 10.6151
R1133 B.n805 B.n804 10.6151
R1134 B.n804 B.n803 10.6151
R1135 B.n803 B.n24 10.6151
R1136 B.n799 B.n24 10.6151
R1137 B.n799 B.n798 10.6151
R1138 B.n798 B.n797 10.6151
R1139 B.n797 B.n26 10.6151
R1140 B.n793 B.n26 10.6151
R1141 B.n793 B.n792 10.6151
R1142 B.n792 B.n791 10.6151
R1143 B.n791 B.n28 10.6151
R1144 B.n787 B.n28 10.6151
R1145 B.n787 B.n786 10.6151
R1146 B.n786 B.n785 10.6151
R1147 B.n785 B.n30 10.6151
R1148 B.n781 B.n30 10.6151
R1149 B.n781 B.n780 10.6151
R1150 B.n780 B.n779 10.6151
R1151 B.n779 B.n32 10.6151
R1152 B.n775 B.n32 10.6151
R1153 B.n775 B.n774 10.6151
R1154 B.n774 B.n773 10.6151
R1155 B.n773 B.n34 10.6151
R1156 B.n769 B.n34 10.6151
R1157 B.n769 B.n768 10.6151
R1158 B.n768 B.n767 10.6151
R1159 B.n767 B.n36 10.6151
R1160 B.n763 B.n36 10.6151
R1161 B.n763 B.n762 10.6151
R1162 B.n762 B.n761 10.6151
R1163 B.n761 B.n38 10.6151
R1164 B.n757 B.n38 10.6151
R1165 B.n757 B.n756 10.6151
R1166 B.n756 B.n755 10.6151
R1167 B.n755 B.n40 10.6151
R1168 B.n751 B.n40 10.6151
R1169 B.n751 B.n750 10.6151
R1170 B.n750 B.n749 10.6151
R1171 B.n749 B.n42 10.6151
R1172 B.n745 B.n42 10.6151
R1173 B.n745 B.n744 10.6151
R1174 B.n744 B.n743 10.6151
R1175 B.n743 B.n44 10.6151
R1176 B.n739 B.n44 10.6151
R1177 B.n739 B.n738 10.6151
R1178 B.n738 B.n737 10.6151
R1179 B.n737 B.n46 10.6151
R1180 B.n733 B.n46 10.6151
R1181 B.n733 B.n732 10.6151
R1182 B.n732 B.n731 10.6151
R1183 B.n731 B.n48 10.6151
R1184 B.n727 B.n48 10.6151
R1185 B.n727 B.n726 10.6151
R1186 B.n726 B.n725 10.6151
R1187 B.n725 B.n50 10.6151
R1188 B.n721 B.n50 10.6151
R1189 B.n721 B.n720 10.6151
R1190 B.n720 B.n719 10.6151
R1191 B.n719 B.n52 10.6151
R1192 B.n715 B.n52 10.6151
R1193 B.n713 B.n712 10.6151
R1194 B.n712 B.n56 10.6151
R1195 B.n708 B.n56 10.6151
R1196 B.n708 B.n707 10.6151
R1197 B.n707 B.n706 10.6151
R1198 B.n706 B.n58 10.6151
R1199 B.n702 B.n58 10.6151
R1200 B.n702 B.n701 10.6151
R1201 B.n699 B.n62 10.6151
R1202 B.n695 B.n62 10.6151
R1203 B.n695 B.n694 10.6151
R1204 B.n694 B.n693 10.6151
R1205 B.n693 B.n64 10.6151
R1206 B.n689 B.n64 10.6151
R1207 B.n689 B.n688 10.6151
R1208 B.n688 B.n687 10.6151
R1209 B.n687 B.n66 10.6151
R1210 B.n683 B.n66 10.6151
R1211 B.n683 B.n682 10.6151
R1212 B.n682 B.n681 10.6151
R1213 B.n681 B.n68 10.6151
R1214 B.n677 B.n68 10.6151
R1215 B.n677 B.n676 10.6151
R1216 B.n676 B.n675 10.6151
R1217 B.n675 B.n70 10.6151
R1218 B.n671 B.n70 10.6151
R1219 B.n671 B.n670 10.6151
R1220 B.n670 B.n669 10.6151
R1221 B.n669 B.n72 10.6151
R1222 B.n665 B.n72 10.6151
R1223 B.n665 B.n664 10.6151
R1224 B.n664 B.n663 10.6151
R1225 B.n663 B.n74 10.6151
R1226 B.n659 B.n74 10.6151
R1227 B.n659 B.n658 10.6151
R1228 B.n658 B.n657 10.6151
R1229 B.n657 B.n76 10.6151
R1230 B.n653 B.n76 10.6151
R1231 B.n653 B.n652 10.6151
R1232 B.n652 B.n651 10.6151
R1233 B.n651 B.n78 10.6151
R1234 B.n647 B.n78 10.6151
R1235 B.n647 B.n646 10.6151
R1236 B.n646 B.n645 10.6151
R1237 B.n645 B.n80 10.6151
R1238 B.n641 B.n80 10.6151
R1239 B.n641 B.n640 10.6151
R1240 B.n640 B.n639 10.6151
R1241 B.n639 B.n82 10.6151
R1242 B.n635 B.n82 10.6151
R1243 B.n635 B.n634 10.6151
R1244 B.n634 B.n633 10.6151
R1245 B.n633 B.n84 10.6151
R1246 B.n629 B.n84 10.6151
R1247 B.n629 B.n628 10.6151
R1248 B.n628 B.n627 10.6151
R1249 B.n627 B.n86 10.6151
R1250 B.n623 B.n86 10.6151
R1251 B.n623 B.n622 10.6151
R1252 B.n622 B.n621 10.6151
R1253 B.n621 B.n88 10.6151
R1254 B.n617 B.n88 10.6151
R1255 B.n617 B.n616 10.6151
R1256 B.n616 B.n615 10.6151
R1257 B.n615 B.n90 10.6151
R1258 B.n611 B.n90 10.6151
R1259 B.n611 B.n610 10.6151
R1260 B.n610 B.n609 10.6151
R1261 B.n609 B.n92 10.6151
R1262 B.n605 B.n92 10.6151
R1263 B.n604 B.n603 10.6151
R1264 B.n603 B.n94 10.6151
R1265 B.n599 B.n94 10.6151
R1266 B.n599 B.n598 10.6151
R1267 B.n598 B.n597 10.6151
R1268 B.n597 B.n96 10.6151
R1269 B.n593 B.n96 10.6151
R1270 B.n593 B.n592 10.6151
R1271 B.n592 B.n591 10.6151
R1272 B.n591 B.n98 10.6151
R1273 B.n587 B.n98 10.6151
R1274 B.n587 B.n586 10.6151
R1275 B.n586 B.n585 10.6151
R1276 B.n585 B.n100 10.6151
R1277 B.n581 B.n100 10.6151
R1278 B.n581 B.n580 10.6151
R1279 B.n580 B.n579 10.6151
R1280 B.n579 B.n102 10.6151
R1281 B.n575 B.n102 10.6151
R1282 B.n575 B.n574 10.6151
R1283 B.n574 B.n573 10.6151
R1284 B.n573 B.n104 10.6151
R1285 B.n569 B.n104 10.6151
R1286 B.n569 B.n568 10.6151
R1287 B.n568 B.n567 10.6151
R1288 B.n567 B.n106 10.6151
R1289 B.n563 B.n106 10.6151
R1290 B.n563 B.n562 10.6151
R1291 B.n562 B.n561 10.6151
R1292 B.n561 B.n108 10.6151
R1293 B.n557 B.n108 10.6151
R1294 B.n557 B.n556 10.6151
R1295 B.n556 B.n555 10.6151
R1296 B.n555 B.n110 10.6151
R1297 B.n551 B.n110 10.6151
R1298 B.n551 B.n550 10.6151
R1299 B.n550 B.n549 10.6151
R1300 B.n549 B.n112 10.6151
R1301 B.n545 B.n112 10.6151
R1302 B.n545 B.n544 10.6151
R1303 B.n544 B.n543 10.6151
R1304 B.n543 B.n114 10.6151
R1305 B.n539 B.n114 10.6151
R1306 B.n539 B.n538 10.6151
R1307 B.n538 B.n537 10.6151
R1308 B.n537 B.n116 10.6151
R1309 B.n533 B.n116 10.6151
R1310 B.n533 B.n532 10.6151
R1311 B.n532 B.n531 10.6151
R1312 B.n531 B.n118 10.6151
R1313 B.n527 B.n118 10.6151
R1314 B.n527 B.n526 10.6151
R1315 B.n526 B.n525 10.6151
R1316 B.n525 B.n120 10.6151
R1317 B.n521 B.n120 10.6151
R1318 B.n521 B.n520 10.6151
R1319 B.n520 B.n519 10.6151
R1320 B.n519 B.n122 10.6151
R1321 B.n515 B.n122 10.6151
R1322 B.n515 B.n514 10.6151
R1323 B.n514 B.n513 10.6151
R1324 B.n513 B.n124 10.6151
R1325 B.n509 B.n124 10.6151
R1326 B.n509 B.n508 10.6151
R1327 B.n508 B.n507 10.6151
R1328 B.n507 B.n126 10.6151
R1329 B.n503 B.n126 10.6151
R1330 B.n503 B.n502 10.6151
R1331 B.n502 B.n501 10.6151
R1332 B.n501 B.n128 10.6151
R1333 B.n497 B.n128 10.6151
R1334 B.n497 B.n496 10.6151
R1335 B.n496 B.n495 10.6151
R1336 B.n495 B.n130 10.6151
R1337 B.n491 B.n130 10.6151
R1338 B.n491 B.n490 10.6151
R1339 B.n490 B.n489 10.6151
R1340 B.n489 B.n132 10.6151
R1341 B.n485 B.n132 10.6151
R1342 B.n222 B.n1 10.6151
R1343 B.n223 B.n222 10.6151
R1344 B.n223 B.n220 10.6151
R1345 B.n227 B.n220 10.6151
R1346 B.n228 B.n227 10.6151
R1347 B.n229 B.n228 10.6151
R1348 B.n229 B.n218 10.6151
R1349 B.n233 B.n218 10.6151
R1350 B.n234 B.n233 10.6151
R1351 B.n235 B.n234 10.6151
R1352 B.n235 B.n216 10.6151
R1353 B.n239 B.n216 10.6151
R1354 B.n240 B.n239 10.6151
R1355 B.n241 B.n240 10.6151
R1356 B.n241 B.n214 10.6151
R1357 B.n245 B.n214 10.6151
R1358 B.n246 B.n245 10.6151
R1359 B.n247 B.n246 10.6151
R1360 B.n247 B.n212 10.6151
R1361 B.n251 B.n212 10.6151
R1362 B.n252 B.n251 10.6151
R1363 B.n253 B.n252 10.6151
R1364 B.n253 B.n210 10.6151
R1365 B.n257 B.n210 10.6151
R1366 B.n258 B.n257 10.6151
R1367 B.n259 B.n258 10.6151
R1368 B.n259 B.n208 10.6151
R1369 B.n263 B.n208 10.6151
R1370 B.n264 B.n263 10.6151
R1371 B.n265 B.n264 10.6151
R1372 B.n265 B.n206 10.6151
R1373 B.n269 B.n206 10.6151
R1374 B.n270 B.n269 10.6151
R1375 B.n271 B.n270 10.6151
R1376 B.n271 B.n204 10.6151
R1377 B.n275 B.n204 10.6151
R1378 B.n276 B.n275 10.6151
R1379 B.n277 B.n276 10.6151
R1380 B.n281 B.n202 10.6151
R1381 B.n282 B.n281 10.6151
R1382 B.n283 B.n282 10.6151
R1383 B.n283 B.n200 10.6151
R1384 B.n287 B.n200 10.6151
R1385 B.n288 B.n287 10.6151
R1386 B.n289 B.n288 10.6151
R1387 B.n289 B.n198 10.6151
R1388 B.n293 B.n198 10.6151
R1389 B.n294 B.n293 10.6151
R1390 B.n295 B.n294 10.6151
R1391 B.n295 B.n196 10.6151
R1392 B.n299 B.n196 10.6151
R1393 B.n300 B.n299 10.6151
R1394 B.n301 B.n300 10.6151
R1395 B.n301 B.n194 10.6151
R1396 B.n305 B.n194 10.6151
R1397 B.n306 B.n305 10.6151
R1398 B.n307 B.n306 10.6151
R1399 B.n307 B.n192 10.6151
R1400 B.n311 B.n192 10.6151
R1401 B.n312 B.n311 10.6151
R1402 B.n313 B.n312 10.6151
R1403 B.n313 B.n190 10.6151
R1404 B.n317 B.n190 10.6151
R1405 B.n318 B.n317 10.6151
R1406 B.n319 B.n318 10.6151
R1407 B.n319 B.n188 10.6151
R1408 B.n323 B.n188 10.6151
R1409 B.n324 B.n323 10.6151
R1410 B.n325 B.n324 10.6151
R1411 B.n325 B.n186 10.6151
R1412 B.n329 B.n186 10.6151
R1413 B.n330 B.n329 10.6151
R1414 B.n331 B.n330 10.6151
R1415 B.n331 B.n184 10.6151
R1416 B.n335 B.n184 10.6151
R1417 B.n336 B.n335 10.6151
R1418 B.n337 B.n336 10.6151
R1419 B.n337 B.n182 10.6151
R1420 B.n341 B.n182 10.6151
R1421 B.n342 B.n341 10.6151
R1422 B.n343 B.n342 10.6151
R1423 B.n343 B.n180 10.6151
R1424 B.n347 B.n180 10.6151
R1425 B.n348 B.n347 10.6151
R1426 B.n349 B.n348 10.6151
R1427 B.n349 B.n178 10.6151
R1428 B.n353 B.n178 10.6151
R1429 B.n354 B.n353 10.6151
R1430 B.n355 B.n354 10.6151
R1431 B.n355 B.n176 10.6151
R1432 B.n359 B.n176 10.6151
R1433 B.n360 B.n359 10.6151
R1434 B.n361 B.n360 10.6151
R1435 B.n361 B.n174 10.6151
R1436 B.n365 B.n174 10.6151
R1437 B.n366 B.n365 10.6151
R1438 B.n367 B.n366 10.6151
R1439 B.n367 B.n172 10.6151
R1440 B.n371 B.n172 10.6151
R1441 B.n372 B.n371 10.6151
R1442 B.n374 B.n168 10.6151
R1443 B.n378 B.n168 10.6151
R1444 B.n379 B.n378 10.6151
R1445 B.n380 B.n379 10.6151
R1446 B.n380 B.n166 10.6151
R1447 B.n384 B.n166 10.6151
R1448 B.n385 B.n384 10.6151
R1449 B.n389 B.n385 10.6151
R1450 B.n393 B.n164 10.6151
R1451 B.n394 B.n393 10.6151
R1452 B.n395 B.n394 10.6151
R1453 B.n395 B.n162 10.6151
R1454 B.n399 B.n162 10.6151
R1455 B.n400 B.n399 10.6151
R1456 B.n401 B.n400 10.6151
R1457 B.n401 B.n160 10.6151
R1458 B.n405 B.n160 10.6151
R1459 B.n406 B.n405 10.6151
R1460 B.n407 B.n406 10.6151
R1461 B.n407 B.n158 10.6151
R1462 B.n411 B.n158 10.6151
R1463 B.n412 B.n411 10.6151
R1464 B.n413 B.n412 10.6151
R1465 B.n413 B.n156 10.6151
R1466 B.n417 B.n156 10.6151
R1467 B.n418 B.n417 10.6151
R1468 B.n419 B.n418 10.6151
R1469 B.n419 B.n154 10.6151
R1470 B.n423 B.n154 10.6151
R1471 B.n424 B.n423 10.6151
R1472 B.n425 B.n424 10.6151
R1473 B.n425 B.n152 10.6151
R1474 B.n429 B.n152 10.6151
R1475 B.n430 B.n429 10.6151
R1476 B.n431 B.n430 10.6151
R1477 B.n431 B.n150 10.6151
R1478 B.n435 B.n150 10.6151
R1479 B.n436 B.n435 10.6151
R1480 B.n437 B.n436 10.6151
R1481 B.n437 B.n148 10.6151
R1482 B.n441 B.n148 10.6151
R1483 B.n442 B.n441 10.6151
R1484 B.n443 B.n442 10.6151
R1485 B.n443 B.n146 10.6151
R1486 B.n447 B.n146 10.6151
R1487 B.n448 B.n447 10.6151
R1488 B.n449 B.n448 10.6151
R1489 B.n449 B.n144 10.6151
R1490 B.n453 B.n144 10.6151
R1491 B.n454 B.n453 10.6151
R1492 B.n455 B.n454 10.6151
R1493 B.n455 B.n142 10.6151
R1494 B.n459 B.n142 10.6151
R1495 B.n460 B.n459 10.6151
R1496 B.n461 B.n460 10.6151
R1497 B.n461 B.n140 10.6151
R1498 B.n465 B.n140 10.6151
R1499 B.n466 B.n465 10.6151
R1500 B.n467 B.n466 10.6151
R1501 B.n467 B.n138 10.6151
R1502 B.n471 B.n138 10.6151
R1503 B.n472 B.n471 10.6151
R1504 B.n473 B.n472 10.6151
R1505 B.n473 B.n136 10.6151
R1506 B.n477 B.n136 10.6151
R1507 B.n478 B.n477 10.6151
R1508 B.n479 B.n478 10.6151
R1509 B.n479 B.n134 10.6151
R1510 B.n483 B.n134 10.6151
R1511 B.n484 B.n483 10.6151
R1512 B.n869 B.n0 8.11757
R1513 B.n869 B.n1 8.11757
R1514 B.n714 B.n713 6.5566
R1515 B.n701 B.n700 6.5566
R1516 B.n374 B.n373 6.5566
R1517 B.n389 B.n388 6.5566
R1518 B.n715 B.n714 4.05904
R1519 B.n700 B.n699 4.05904
R1520 B.n373 B.n372 4.05904
R1521 B.n388 B.n164 4.05904
C0 VP VN 8.001471f
C1 w_n3100_n4792# VDD1 1.88271f
C2 B VTAIL 6.78474f
C3 VN VDD1 0.150516f
C4 VDD2 VTAIL 11.1993f
C5 VP VDD1 12.747299f
C6 w_n3100_n4792# B 10.886701f
C7 VN B 1.12571f
C8 w_n3100_n4792# VDD2 1.96386f
C9 VP B 1.79213f
C10 VN VDD2 12.464f
C11 VP VDD2 0.434777f
C12 B VDD1 1.59802f
C13 VDD2 VDD1 1.36049f
C14 w_n3100_n4792# VTAIL 5.82093f
C15 VN VTAIL 12.3076f
C16 VP VTAIL 12.3217f
C17 B VDD2 1.66887f
C18 VDD1 VTAIL 11.1503f
C19 w_n3100_n4792# VN 6.21828f
C20 VP w_n3100_n4792# 6.61836f
C21 VDD2 VSUBS 1.763768f
C22 VDD1 VSUBS 2.265364f
C23 VTAIL VSUBS 1.52858f
C24 VN VSUBS 6.12851f
C25 VP VSUBS 3.036208f
C26 B VSUBS 4.710509f
C27 w_n3100_n4792# VSUBS 0.181499p
C28 B.n0 VSUBS 0.005778f
C29 B.n1 VSUBS 0.005778f
C30 B.n2 VSUBS 0.008545f
C31 B.n3 VSUBS 0.006548f
C32 B.n4 VSUBS 0.006548f
C33 B.n5 VSUBS 0.006548f
C34 B.n6 VSUBS 0.006548f
C35 B.n7 VSUBS 0.006548f
C36 B.n8 VSUBS 0.006548f
C37 B.n9 VSUBS 0.006548f
C38 B.n10 VSUBS 0.006548f
C39 B.n11 VSUBS 0.006548f
C40 B.n12 VSUBS 0.006548f
C41 B.n13 VSUBS 0.006548f
C42 B.n14 VSUBS 0.006548f
C43 B.n15 VSUBS 0.006548f
C44 B.n16 VSUBS 0.006548f
C45 B.n17 VSUBS 0.006548f
C46 B.n18 VSUBS 0.006548f
C47 B.n19 VSUBS 0.006548f
C48 B.n20 VSUBS 0.006548f
C49 B.n21 VSUBS 0.014081f
C50 B.n22 VSUBS 0.006548f
C51 B.n23 VSUBS 0.006548f
C52 B.n24 VSUBS 0.006548f
C53 B.n25 VSUBS 0.006548f
C54 B.n26 VSUBS 0.006548f
C55 B.n27 VSUBS 0.006548f
C56 B.n28 VSUBS 0.006548f
C57 B.n29 VSUBS 0.006548f
C58 B.n30 VSUBS 0.006548f
C59 B.n31 VSUBS 0.006548f
C60 B.n32 VSUBS 0.006548f
C61 B.n33 VSUBS 0.006548f
C62 B.n34 VSUBS 0.006548f
C63 B.n35 VSUBS 0.006548f
C64 B.n36 VSUBS 0.006548f
C65 B.n37 VSUBS 0.006548f
C66 B.n38 VSUBS 0.006548f
C67 B.n39 VSUBS 0.006548f
C68 B.n40 VSUBS 0.006548f
C69 B.n41 VSUBS 0.006548f
C70 B.n42 VSUBS 0.006548f
C71 B.n43 VSUBS 0.006548f
C72 B.n44 VSUBS 0.006548f
C73 B.n45 VSUBS 0.006548f
C74 B.n46 VSUBS 0.006548f
C75 B.n47 VSUBS 0.006548f
C76 B.n48 VSUBS 0.006548f
C77 B.n49 VSUBS 0.006548f
C78 B.n50 VSUBS 0.006548f
C79 B.n51 VSUBS 0.006548f
C80 B.n52 VSUBS 0.006548f
C81 B.n53 VSUBS 0.006548f
C82 B.t4 VSUBS 0.606278f
C83 B.t5 VSUBS 0.621554f
C84 B.t3 VSUBS 1.38273f
C85 B.n54 VSUBS 0.29536f
C86 B.n55 VSUBS 0.064414f
C87 B.n56 VSUBS 0.006548f
C88 B.n57 VSUBS 0.006548f
C89 B.n58 VSUBS 0.006548f
C90 B.n59 VSUBS 0.006548f
C91 B.t10 VSUBS 0.606253f
C92 B.t11 VSUBS 0.621533f
C93 B.t9 VSUBS 1.38273f
C94 B.n60 VSUBS 0.29538f
C95 B.n61 VSUBS 0.064439f
C96 B.n62 VSUBS 0.006548f
C97 B.n63 VSUBS 0.006548f
C98 B.n64 VSUBS 0.006548f
C99 B.n65 VSUBS 0.006548f
C100 B.n66 VSUBS 0.006548f
C101 B.n67 VSUBS 0.006548f
C102 B.n68 VSUBS 0.006548f
C103 B.n69 VSUBS 0.006548f
C104 B.n70 VSUBS 0.006548f
C105 B.n71 VSUBS 0.006548f
C106 B.n72 VSUBS 0.006548f
C107 B.n73 VSUBS 0.006548f
C108 B.n74 VSUBS 0.006548f
C109 B.n75 VSUBS 0.006548f
C110 B.n76 VSUBS 0.006548f
C111 B.n77 VSUBS 0.006548f
C112 B.n78 VSUBS 0.006548f
C113 B.n79 VSUBS 0.006548f
C114 B.n80 VSUBS 0.006548f
C115 B.n81 VSUBS 0.006548f
C116 B.n82 VSUBS 0.006548f
C117 B.n83 VSUBS 0.006548f
C118 B.n84 VSUBS 0.006548f
C119 B.n85 VSUBS 0.006548f
C120 B.n86 VSUBS 0.006548f
C121 B.n87 VSUBS 0.006548f
C122 B.n88 VSUBS 0.006548f
C123 B.n89 VSUBS 0.006548f
C124 B.n90 VSUBS 0.006548f
C125 B.n91 VSUBS 0.006548f
C126 B.n92 VSUBS 0.006548f
C127 B.n93 VSUBS 0.014081f
C128 B.n94 VSUBS 0.006548f
C129 B.n95 VSUBS 0.006548f
C130 B.n96 VSUBS 0.006548f
C131 B.n97 VSUBS 0.006548f
C132 B.n98 VSUBS 0.006548f
C133 B.n99 VSUBS 0.006548f
C134 B.n100 VSUBS 0.006548f
C135 B.n101 VSUBS 0.006548f
C136 B.n102 VSUBS 0.006548f
C137 B.n103 VSUBS 0.006548f
C138 B.n104 VSUBS 0.006548f
C139 B.n105 VSUBS 0.006548f
C140 B.n106 VSUBS 0.006548f
C141 B.n107 VSUBS 0.006548f
C142 B.n108 VSUBS 0.006548f
C143 B.n109 VSUBS 0.006548f
C144 B.n110 VSUBS 0.006548f
C145 B.n111 VSUBS 0.006548f
C146 B.n112 VSUBS 0.006548f
C147 B.n113 VSUBS 0.006548f
C148 B.n114 VSUBS 0.006548f
C149 B.n115 VSUBS 0.006548f
C150 B.n116 VSUBS 0.006548f
C151 B.n117 VSUBS 0.006548f
C152 B.n118 VSUBS 0.006548f
C153 B.n119 VSUBS 0.006548f
C154 B.n120 VSUBS 0.006548f
C155 B.n121 VSUBS 0.006548f
C156 B.n122 VSUBS 0.006548f
C157 B.n123 VSUBS 0.006548f
C158 B.n124 VSUBS 0.006548f
C159 B.n125 VSUBS 0.006548f
C160 B.n126 VSUBS 0.006548f
C161 B.n127 VSUBS 0.006548f
C162 B.n128 VSUBS 0.006548f
C163 B.n129 VSUBS 0.006548f
C164 B.n130 VSUBS 0.006548f
C165 B.n131 VSUBS 0.006548f
C166 B.n132 VSUBS 0.006548f
C167 B.n133 VSUBS 0.015001f
C168 B.n134 VSUBS 0.006548f
C169 B.n135 VSUBS 0.006548f
C170 B.n136 VSUBS 0.006548f
C171 B.n137 VSUBS 0.006548f
C172 B.n138 VSUBS 0.006548f
C173 B.n139 VSUBS 0.006548f
C174 B.n140 VSUBS 0.006548f
C175 B.n141 VSUBS 0.006548f
C176 B.n142 VSUBS 0.006548f
C177 B.n143 VSUBS 0.006548f
C178 B.n144 VSUBS 0.006548f
C179 B.n145 VSUBS 0.006548f
C180 B.n146 VSUBS 0.006548f
C181 B.n147 VSUBS 0.006548f
C182 B.n148 VSUBS 0.006548f
C183 B.n149 VSUBS 0.006548f
C184 B.n150 VSUBS 0.006548f
C185 B.n151 VSUBS 0.006548f
C186 B.n152 VSUBS 0.006548f
C187 B.n153 VSUBS 0.006548f
C188 B.n154 VSUBS 0.006548f
C189 B.n155 VSUBS 0.006548f
C190 B.n156 VSUBS 0.006548f
C191 B.n157 VSUBS 0.006548f
C192 B.n158 VSUBS 0.006548f
C193 B.n159 VSUBS 0.006548f
C194 B.n160 VSUBS 0.006548f
C195 B.n161 VSUBS 0.006548f
C196 B.n162 VSUBS 0.006548f
C197 B.n163 VSUBS 0.006548f
C198 B.n164 VSUBS 0.004526f
C199 B.n165 VSUBS 0.006548f
C200 B.n166 VSUBS 0.006548f
C201 B.n167 VSUBS 0.006548f
C202 B.n168 VSUBS 0.006548f
C203 B.n169 VSUBS 0.006548f
C204 B.t2 VSUBS 0.606278f
C205 B.t1 VSUBS 0.621554f
C206 B.t0 VSUBS 1.38273f
C207 B.n170 VSUBS 0.29536f
C208 B.n171 VSUBS 0.064414f
C209 B.n172 VSUBS 0.006548f
C210 B.n173 VSUBS 0.006548f
C211 B.n174 VSUBS 0.006548f
C212 B.n175 VSUBS 0.006548f
C213 B.n176 VSUBS 0.006548f
C214 B.n177 VSUBS 0.006548f
C215 B.n178 VSUBS 0.006548f
C216 B.n179 VSUBS 0.006548f
C217 B.n180 VSUBS 0.006548f
C218 B.n181 VSUBS 0.006548f
C219 B.n182 VSUBS 0.006548f
C220 B.n183 VSUBS 0.006548f
C221 B.n184 VSUBS 0.006548f
C222 B.n185 VSUBS 0.006548f
C223 B.n186 VSUBS 0.006548f
C224 B.n187 VSUBS 0.006548f
C225 B.n188 VSUBS 0.006548f
C226 B.n189 VSUBS 0.006548f
C227 B.n190 VSUBS 0.006548f
C228 B.n191 VSUBS 0.006548f
C229 B.n192 VSUBS 0.006548f
C230 B.n193 VSUBS 0.006548f
C231 B.n194 VSUBS 0.006548f
C232 B.n195 VSUBS 0.006548f
C233 B.n196 VSUBS 0.006548f
C234 B.n197 VSUBS 0.006548f
C235 B.n198 VSUBS 0.006548f
C236 B.n199 VSUBS 0.006548f
C237 B.n200 VSUBS 0.006548f
C238 B.n201 VSUBS 0.006548f
C239 B.n202 VSUBS 0.015001f
C240 B.n203 VSUBS 0.006548f
C241 B.n204 VSUBS 0.006548f
C242 B.n205 VSUBS 0.006548f
C243 B.n206 VSUBS 0.006548f
C244 B.n207 VSUBS 0.006548f
C245 B.n208 VSUBS 0.006548f
C246 B.n209 VSUBS 0.006548f
C247 B.n210 VSUBS 0.006548f
C248 B.n211 VSUBS 0.006548f
C249 B.n212 VSUBS 0.006548f
C250 B.n213 VSUBS 0.006548f
C251 B.n214 VSUBS 0.006548f
C252 B.n215 VSUBS 0.006548f
C253 B.n216 VSUBS 0.006548f
C254 B.n217 VSUBS 0.006548f
C255 B.n218 VSUBS 0.006548f
C256 B.n219 VSUBS 0.006548f
C257 B.n220 VSUBS 0.006548f
C258 B.n221 VSUBS 0.006548f
C259 B.n222 VSUBS 0.006548f
C260 B.n223 VSUBS 0.006548f
C261 B.n224 VSUBS 0.006548f
C262 B.n225 VSUBS 0.006548f
C263 B.n226 VSUBS 0.006548f
C264 B.n227 VSUBS 0.006548f
C265 B.n228 VSUBS 0.006548f
C266 B.n229 VSUBS 0.006548f
C267 B.n230 VSUBS 0.006548f
C268 B.n231 VSUBS 0.006548f
C269 B.n232 VSUBS 0.006548f
C270 B.n233 VSUBS 0.006548f
C271 B.n234 VSUBS 0.006548f
C272 B.n235 VSUBS 0.006548f
C273 B.n236 VSUBS 0.006548f
C274 B.n237 VSUBS 0.006548f
C275 B.n238 VSUBS 0.006548f
C276 B.n239 VSUBS 0.006548f
C277 B.n240 VSUBS 0.006548f
C278 B.n241 VSUBS 0.006548f
C279 B.n242 VSUBS 0.006548f
C280 B.n243 VSUBS 0.006548f
C281 B.n244 VSUBS 0.006548f
C282 B.n245 VSUBS 0.006548f
C283 B.n246 VSUBS 0.006548f
C284 B.n247 VSUBS 0.006548f
C285 B.n248 VSUBS 0.006548f
C286 B.n249 VSUBS 0.006548f
C287 B.n250 VSUBS 0.006548f
C288 B.n251 VSUBS 0.006548f
C289 B.n252 VSUBS 0.006548f
C290 B.n253 VSUBS 0.006548f
C291 B.n254 VSUBS 0.006548f
C292 B.n255 VSUBS 0.006548f
C293 B.n256 VSUBS 0.006548f
C294 B.n257 VSUBS 0.006548f
C295 B.n258 VSUBS 0.006548f
C296 B.n259 VSUBS 0.006548f
C297 B.n260 VSUBS 0.006548f
C298 B.n261 VSUBS 0.006548f
C299 B.n262 VSUBS 0.006548f
C300 B.n263 VSUBS 0.006548f
C301 B.n264 VSUBS 0.006548f
C302 B.n265 VSUBS 0.006548f
C303 B.n266 VSUBS 0.006548f
C304 B.n267 VSUBS 0.006548f
C305 B.n268 VSUBS 0.006548f
C306 B.n269 VSUBS 0.006548f
C307 B.n270 VSUBS 0.006548f
C308 B.n271 VSUBS 0.006548f
C309 B.n272 VSUBS 0.006548f
C310 B.n273 VSUBS 0.006548f
C311 B.n274 VSUBS 0.006548f
C312 B.n275 VSUBS 0.006548f
C313 B.n276 VSUBS 0.006548f
C314 B.n277 VSUBS 0.014081f
C315 B.n278 VSUBS 0.014081f
C316 B.n279 VSUBS 0.015001f
C317 B.n280 VSUBS 0.006548f
C318 B.n281 VSUBS 0.006548f
C319 B.n282 VSUBS 0.006548f
C320 B.n283 VSUBS 0.006548f
C321 B.n284 VSUBS 0.006548f
C322 B.n285 VSUBS 0.006548f
C323 B.n286 VSUBS 0.006548f
C324 B.n287 VSUBS 0.006548f
C325 B.n288 VSUBS 0.006548f
C326 B.n289 VSUBS 0.006548f
C327 B.n290 VSUBS 0.006548f
C328 B.n291 VSUBS 0.006548f
C329 B.n292 VSUBS 0.006548f
C330 B.n293 VSUBS 0.006548f
C331 B.n294 VSUBS 0.006548f
C332 B.n295 VSUBS 0.006548f
C333 B.n296 VSUBS 0.006548f
C334 B.n297 VSUBS 0.006548f
C335 B.n298 VSUBS 0.006548f
C336 B.n299 VSUBS 0.006548f
C337 B.n300 VSUBS 0.006548f
C338 B.n301 VSUBS 0.006548f
C339 B.n302 VSUBS 0.006548f
C340 B.n303 VSUBS 0.006548f
C341 B.n304 VSUBS 0.006548f
C342 B.n305 VSUBS 0.006548f
C343 B.n306 VSUBS 0.006548f
C344 B.n307 VSUBS 0.006548f
C345 B.n308 VSUBS 0.006548f
C346 B.n309 VSUBS 0.006548f
C347 B.n310 VSUBS 0.006548f
C348 B.n311 VSUBS 0.006548f
C349 B.n312 VSUBS 0.006548f
C350 B.n313 VSUBS 0.006548f
C351 B.n314 VSUBS 0.006548f
C352 B.n315 VSUBS 0.006548f
C353 B.n316 VSUBS 0.006548f
C354 B.n317 VSUBS 0.006548f
C355 B.n318 VSUBS 0.006548f
C356 B.n319 VSUBS 0.006548f
C357 B.n320 VSUBS 0.006548f
C358 B.n321 VSUBS 0.006548f
C359 B.n322 VSUBS 0.006548f
C360 B.n323 VSUBS 0.006548f
C361 B.n324 VSUBS 0.006548f
C362 B.n325 VSUBS 0.006548f
C363 B.n326 VSUBS 0.006548f
C364 B.n327 VSUBS 0.006548f
C365 B.n328 VSUBS 0.006548f
C366 B.n329 VSUBS 0.006548f
C367 B.n330 VSUBS 0.006548f
C368 B.n331 VSUBS 0.006548f
C369 B.n332 VSUBS 0.006548f
C370 B.n333 VSUBS 0.006548f
C371 B.n334 VSUBS 0.006548f
C372 B.n335 VSUBS 0.006548f
C373 B.n336 VSUBS 0.006548f
C374 B.n337 VSUBS 0.006548f
C375 B.n338 VSUBS 0.006548f
C376 B.n339 VSUBS 0.006548f
C377 B.n340 VSUBS 0.006548f
C378 B.n341 VSUBS 0.006548f
C379 B.n342 VSUBS 0.006548f
C380 B.n343 VSUBS 0.006548f
C381 B.n344 VSUBS 0.006548f
C382 B.n345 VSUBS 0.006548f
C383 B.n346 VSUBS 0.006548f
C384 B.n347 VSUBS 0.006548f
C385 B.n348 VSUBS 0.006548f
C386 B.n349 VSUBS 0.006548f
C387 B.n350 VSUBS 0.006548f
C388 B.n351 VSUBS 0.006548f
C389 B.n352 VSUBS 0.006548f
C390 B.n353 VSUBS 0.006548f
C391 B.n354 VSUBS 0.006548f
C392 B.n355 VSUBS 0.006548f
C393 B.n356 VSUBS 0.006548f
C394 B.n357 VSUBS 0.006548f
C395 B.n358 VSUBS 0.006548f
C396 B.n359 VSUBS 0.006548f
C397 B.n360 VSUBS 0.006548f
C398 B.n361 VSUBS 0.006548f
C399 B.n362 VSUBS 0.006548f
C400 B.n363 VSUBS 0.006548f
C401 B.n364 VSUBS 0.006548f
C402 B.n365 VSUBS 0.006548f
C403 B.n366 VSUBS 0.006548f
C404 B.n367 VSUBS 0.006548f
C405 B.n368 VSUBS 0.006548f
C406 B.n369 VSUBS 0.006548f
C407 B.n370 VSUBS 0.006548f
C408 B.n371 VSUBS 0.006548f
C409 B.n372 VSUBS 0.004526f
C410 B.n373 VSUBS 0.015171f
C411 B.n374 VSUBS 0.005296f
C412 B.n375 VSUBS 0.006548f
C413 B.n376 VSUBS 0.006548f
C414 B.n377 VSUBS 0.006548f
C415 B.n378 VSUBS 0.006548f
C416 B.n379 VSUBS 0.006548f
C417 B.n380 VSUBS 0.006548f
C418 B.n381 VSUBS 0.006548f
C419 B.n382 VSUBS 0.006548f
C420 B.n383 VSUBS 0.006548f
C421 B.n384 VSUBS 0.006548f
C422 B.n385 VSUBS 0.006548f
C423 B.t8 VSUBS 0.606253f
C424 B.t7 VSUBS 0.621533f
C425 B.t6 VSUBS 1.38273f
C426 B.n386 VSUBS 0.29538f
C427 B.n387 VSUBS 0.064439f
C428 B.n388 VSUBS 0.015171f
C429 B.n389 VSUBS 0.005296f
C430 B.n390 VSUBS 0.006548f
C431 B.n391 VSUBS 0.006548f
C432 B.n392 VSUBS 0.006548f
C433 B.n393 VSUBS 0.006548f
C434 B.n394 VSUBS 0.006548f
C435 B.n395 VSUBS 0.006548f
C436 B.n396 VSUBS 0.006548f
C437 B.n397 VSUBS 0.006548f
C438 B.n398 VSUBS 0.006548f
C439 B.n399 VSUBS 0.006548f
C440 B.n400 VSUBS 0.006548f
C441 B.n401 VSUBS 0.006548f
C442 B.n402 VSUBS 0.006548f
C443 B.n403 VSUBS 0.006548f
C444 B.n404 VSUBS 0.006548f
C445 B.n405 VSUBS 0.006548f
C446 B.n406 VSUBS 0.006548f
C447 B.n407 VSUBS 0.006548f
C448 B.n408 VSUBS 0.006548f
C449 B.n409 VSUBS 0.006548f
C450 B.n410 VSUBS 0.006548f
C451 B.n411 VSUBS 0.006548f
C452 B.n412 VSUBS 0.006548f
C453 B.n413 VSUBS 0.006548f
C454 B.n414 VSUBS 0.006548f
C455 B.n415 VSUBS 0.006548f
C456 B.n416 VSUBS 0.006548f
C457 B.n417 VSUBS 0.006548f
C458 B.n418 VSUBS 0.006548f
C459 B.n419 VSUBS 0.006548f
C460 B.n420 VSUBS 0.006548f
C461 B.n421 VSUBS 0.006548f
C462 B.n422 VSUBS 0.006548f
C463 B.n423 VSUBS 0.006548f
C464 B.n424 VSUBS 0.006548f
C465 B.n425 VSUBS 0.006548f
C466 B.n426 VSUBS 0.006548f
C467 B.n427 VSUBS 0.006548f
C468 B.n428 VSUBS 0.006548f
C469 B.n429 VSUBS 0.006548f
C470 B.n430 VSUBS 0.006548f
C471 B.n431 VSUBS 0.006548f
C472 B.n432 VSUBS 0.006548f
C473 B.n433 VSUBS 0.006548f
C474 B.n434 VSUBS 0.006548f
C475 B.n435 VSUBS 0.006548f
C476 B.n436 VSUBS 0.006548f
C477 B.n437 VSUBS 0.006548f
C478 B.n438 VSUBS 0.006548f
C479 B.n439 VSUBS 0.006548f
C480 B.n440 VSUBS 0.006548f
C481 B.n441 VSUBS 0.006548f
C482 B.n442 VSUBS 0.006548f
C483 B.n443 VSUBS 0.006548f
C484 B.n444 VSUBS 0.006548f
C485 B.n445 VSUBS 0.006548f
C486 B.n446 VSUBS 0.006548f
C487 B.n447 VSUBS 0.006548f
C488 B.n448 VSUBS 0.006548f
C489 B.n449 VSUBS 0.006548f
C490 B.n450 VSUBS 0.006548f
C491 B.n451 VSUBS 0.006548f
C492 B.n452 VSUBS 0.006548f
C493 B.n453 VSUBS 0.006548f
C494 B.n454 VSUBS 0.006548f
C495 B.n455 VSUBS 0.006548f
C496 B.n456 VSUBS 0.006548f
C497 B.n457 VSUBS 0.006548f
C498 B.n458 VSUBS 0.006548f
C499 B.n459 VSUBS 0.006548f
C500 B.n460 VSUBS 0.006548f
C501 B.n461 VSUBS 0.006548f
C502 B.n462 VSUBS 0.006548f
C503 B.n463 VSUBS 0.006548f
C504 B.n464 VSUBS 0.006548f
C505 B.n465 VSUBS 0.006548f
C506 B.n466 VSUBS 0.006548f
C507 B.n467 VSUBS 0.006548f
C508 B.n468 VSUBS 0.006548f
C509 B.n469 VSUBS 0.006548f
C510 B.n470 VSUBS 0.006548f
C511 B.n471 VSUBS 0.006548f
C512 B.n472 VSUBS 0.006548f
C513 B.n473 VSUBS 0.006548f
C514 B.n474 VSUBS 0.006548f
C515 B.n475 VSUBS 0.006548f
C516 B.n476 VSUBS 0.006548f
C517 B.n477 VSUBS 0.006548f
C518 B.n478 VSUBS 0.006548f
C519 B.n479 VSUBS 0.006548f
C520 B.n480 VSUBS 0.006548f
C521 B.n481 VSUBS 0.006548f
C522 B.n482 VSUBS 0.006548f
C523 B.n483 VSUBS 0.006548f
C524 B.n484 VSUBS 0.014162f
C525 B.n485 VSUBS 0.014919f
C526 B.n486 VSUBS 0.014081f
C527 B.n487 VSUBS 0.006548f
C528 B.n488 VSUBS 0.006548f
C529 B.n489 VSUBS 0.006548f
C530 B.n490 VSUBS 0.006548f
C531 B.n491 VSUBS 0.006548f
C532 B.n492 VSUBS 0.006548f
C533 B.n493 VSUBS 0.006548f
C534 B.n494 VSUBS 0.006548f
C535 B.n495 VSUBS 0.006548f
C536 B.n496 VSUBS 0.006548f
C537 B.n497 VSUBS 0.006548f
C538 B.n498 VSUBS 0.006548f
C539 B.n499 VSUBS 0.006548f
C540 B.n500 VSUBS 0.006548f
C541 B.n501 VSUBS 0.006548f
C542 B.n502 VSUBS 0.006548f
C543 B.n503 VSUBS 0.006548f
C544 B.n504 VSUBS 0.006548f
C545 B.n505 VSUBS 0.006548f
C546 B.n506 VSUBS 0.006548f
C547 B.n507 VSUBS 0.006548f
C548 B.n508 VSUBS 0.006548f
C549 B.n509 VSUBS 0.006548f
C550 B.n510 VSUBS 0.006548f
C551 B.n511 VSUBS 0.006548f
C552 B.n512 VSUBS 0.006548f
C553 B.n513 VSUBS 0.006548f
C554 B.n514 VSUBS 0.006548f
C555 B.n515 VSUBS 0.006548f
C556 B.n516 VSUBS 0.006548f
C557 B.n517 VSUBS 0.006548f
C558 B.n518 VSUBS 0.006548f
C559 B.n519 VSUBS 0.006548f
C560 B.n520 VSUBS 0.006548f
C561 B.n521 VSUBS 0.006548f
C562 B.n522 VSUBS 0.006548f
C563 B.n523 VSUBS 0.006548f
C564 B.n524 VSUBS 0.006548f
C565 B.n525 VSUBS 0.006548f
C566 B.n526 VSUBS 0.006548f
C567 B.n527 VSUBS 0.006548f
C568 B.n528 VSUBS 0.006548f
C569 B.n529 VSUBS 0.006548f
C570 B.n530 VSUBS 0.006548f
C571 B.n531 VSUBS 0.006548f
C572 B.n532 VSUBS 0.006548f
C573 B.n533 VSUBS 0.006548f
C574 B.n534 VSUBS 0.006548f
C575 B.n535 VSUBS 0.006548f
C576 B.n536 VSUBS 0.006548f
C577 B.n537 VSUBS 0.006548f
C578 B.n538 VSUBS 0.006548f
C579 B.n539 VSUBS 0.006548f
C580 B.n540 VSUBS 0.006548f
C581 B.n541 VSUBS 0.006548f
C582 B.n542 VSUBS 0.006548f
C583 B.n543 VSUBS 0.006548f
C584 B.n544 VSUBS 0.006548f
C585 B.n545 VSUBS 0.006548f
C586 B.n546 VSUBS 0.006548f
C587 B.n547 VSUBS 0.006548f
C588 B.n548 VSUBS 0.006548f
C589 B.n549 VSUBS 0.006548f
C590 B.n550 VSUBS 0.006548f
C591 B.n551 VSUBS 0.006548f
C592 B.n552 VSUBS 0.006548f
C593 B.n553 VSUBS 0.006548f
C594 B.n554 VSUBS 0.006548f
C595 B.n555 VSUBS 0.006548f
C596 B.n556 VSUBS 0.006548f
C597 B.n557 VSUBS 0.006548f
C598 B.n558 VSUBS 0.006548f
C599 B.n559 VSUBS 0.006548f
C600 B.n560 VSUBS 0.006548f
C601 B.n561 VSUBS 0.006548f
C602 B.n562 VSUBS 0.006548f
C603 B.n563 VSUBS 0.006548f
C604 B.n564 VSUBS 0.006548f
C605 B.n565 VSUBS 0.006548f
C606 B.n566 VSUBS 0.006548f
C607 B.n567 VSUBS 0.006548f
C608 B.n568 VSUBS 0.006548f
C609 B.n569 VSUBS 0.006548f
C610 B.n570 VSUBS 0.006548f
C611 B.n571 VSUBS 0.006548f
C612 B.n572 VSUBS 0.006548f
C613 B.n573 VSUBS 0.006548f
C614 B.n574 VSUBS 0.006548f
C615 B.n575 VSUBS 0.006548f
C616 B.n576 VSUBS 0.006548f
C617 B.n577 VSUBS 0.006548f
C618 B.n578 VSUBS 0.006548f
C619 B.n579 VSUBS 0.006548f
C620 B.n580 VSUBS 0.006548f
C621 B.n581 VSUBS 0.006548f
C622 B.n582 VSUBS 0.006548f
C623 B.n583 VSUBS 0.006548f
C624 B.n584 VSUBS 0.006548f
C625 B.n585 VSUBS 0.006548f
C626 B.n586 VSUBS 0.006548f
C627 B.n587 VSUBS 0.006548f
C628 B.n588 VSUBS 0.006548f
C629 B.n589 VSUBS 0.006548f
C630 B.n590 VSUBS 0.006548f
C631 B.n591 VSUBS 0.006548f
C632 B.n592 VSUBS 0.006548f
C633 B.n593 VSUBS 0.006548f
C634 B.n594 VSUBS 0.006548f
C635 B.n595 VSUBS 0.006548f
C636 B.n596 VSUBS 0.006548f
C637 B.n597 VSUBS 0.006548f
C638 B.n598 VSUBS 0.006548f
C639 B.n599 VSUBS 0.006548f
C640 B.n600 VSUBS 0.006548f
C641 B.n601 VSUBS 0.006548f
C642 B.n602 VSUBS 0.006548f
C643 B.n603 VSUBS 0.006548f
C644 B.n604 VSUBS 0.014081f
C645 B.n605 VSUBS 0.015001f
C646 B.n606 VSUBS 0.015001f
C647 B.n607 VSUBS 0.006548f
C648 B.n608 VSUBS 0.006548f
C649 B.n609 VSUBS 0.006548f
C650 B.n610 VSUBS 0.006548f
C651 B.n611 VSUBS 0.006548f
C652 B.n612 VSUBS 0.006548f
C653 B.n613 VSUBS 0.006548f
C654 B.n614 VSUBS 0.006548f
C655 B.n615 VSUBS 0.006548f
C656 B.n616 VSUBS 0.006548f
C657 B.n617 VSUBS 0.006548f
C658 B.n618 VSUBS 0.006548f
C659 B.n619 VSUBS 0.006548f
C660 B.n620 VSUBS 0.006548f
C661 B.n621 VSUBS 0.006548f
C662 B.n622 VSUBS 0.006548f
C663 B.n623 VSUBS 0.006548f
C664 B.n624 VSUBS 0.006548f
C665 B.n625 VSUBS 0.006548f
C666 B.n626 VSUBS 0.006548f
C667 B.n627 VSUBS 0.006548f
C668 B.n628 VSUBS 0.006548f
C669 B.n629 VSUBS 0.006548f
C670 B.n630 VSUBS 0.006548f
C671 B.n631 VSUBS 0.006548f
C672 B.n632 VSUBS 0.006548f
C673 B.n633 VSUBS 0.006548f
C674 B.n634 VSUBS 0.006548f
C675 B.n635 VSUBS 0.006548f
C676 B.n636 VSUBS 0.006548f
C677 B.n637 VSUBS 0.006548f
C678 B.n638 VSUBS 0.006548f
C679 B.n639 VSUBS 0.006548f
C680 B.n640 VSUBS 0.006548f
C681 B.n641 VSUBS 0.006548f
C682 B.n642 VSUBS 0.006548f
C683 B.n643 VSUBS 0.006548f
C684 B.n644 VSUBS 0.006548f
C685 B.n645 VSUBS 0.006548f
C686 B.n646 VSUBS 0.006548f
C687 B.n647 VSUBS 0.006548f
C688 B.n648 VSUBS 0.006548f
C689 B.n649 VSUBS 0.006548f
C690 B.n650 VSUBS 0.006548f
C691 B.n651 VSUBS 0.006548f
C692 B.n652 VSUBS 0.006548f
C693 B.n653 VSUBS 0.006548f
C694 B.n654 VSUBS 0.006548f
C695 B.n655 VSUBS 0.006548f
C696 B.n656 VSUBS 0.006548f
C697 B.n657 VSUBS 0.006548f
C698 B.n658 VSUBS 0.006548f
C699 B.n659 VSUBS 0.006548f
C700 B.n660 VSUBS 0.006548f
C701 B.n661 VSUBS 0.006548f
C702 B.n662 VSUBS 0.006548f
C703 B.n663 VSUBS 0.006548f
C704 B.n664 VSUBS 0.006548f
C705 B.n665 VSUBS 0.006548f
C706 B.n666 VSUBS 0.006548f
C707 B.n667 VSUBS 0.006548f
C708 B.n668 VSUBS 0.006548f
C709 B.n669 VSUBS 0.006548f
C710 B.n670 VSUBS 0.006548f
C711 B.n671 VSUBS 0.006548f
C712 B.n672 VSUBS 0.006548f
C713 B.n673 VSUBS 0.006548f
C714 B.n674 VSUBS 0.006548f
C715 B.n675 VSUBS 0.006548f
C716 B.n676 VSUBS 0.006548f
C717 B.n677 VSUBS 0.006548f
C718 B.n678 VSUBS 0.006548f
C719 B.n679 VSUBS 0.006548f
C720 B.n680 VSUBS 0.006548f
C721 B.n681 VSUBS 0.006548f
C722 B.n682 VSUBS 0.006548f
C723 B.n683 VSUBS 0.006548f
C724 B.n684 VSUBS 0.006548f
C725 B.n685 VSUBS 0.006548f
C726 B.n686 VSUBS 0.006548f
C727 B.n687 VSUBS 0.006548f
C728 B.n688 VSUBS 0.006548f
C729 B.n689 VSUBS 0.006548f
C730 B.n690 VSUBS 0.006548f
C731 B.n691 VSUBS 0.006548f
C732 B.n692 VSUBS 0.006548f
C733 B.n693 VSUBS 0.006548f
C734 B.n694 VSUBS 0.006548f
C735 B.n695 VSUBS 0.006548f
C736 B.n696 VSUBS 0.006548f
C737 B.n697 VSUBS 0.006548f
C738 B.n698 VSUBS 0.006548f
C739 B.n699 VSUBS 0.004526f
C740 B.n700 VSUBS 0.015171f
C741 B.n701 VSUBS 0.005296f
C742 B.n702 VSUBS 0.006548f
C743 B.n703 VSUBS 0.006548f
C744 B.n704 VSUBS 0.006548f
C745 B.n705 VSUBS 0.006548f
C746 B.n706 VSUBS 0.006548f
C747 B.n707 VSUBS 0.006548f
C748 B.n708 VSUBS 0.006548f
C749 B.n709 VSUBS 0.006548f
C750 B.n710 VSUBS 0.006548f
C751 B.n711 VSUBS 0.006548f
C752 B.n712 VSUBS 0.006548f
C753 B.n713 VSUBS 0.005296f
C754 B.n714 VSUBS 0.015171f
C755 B.n715 VSUBS 0.004526f
C756 B.n716 VSUBS 0.006548f
C757 B.n717 VSUBS 0.006548f
C758 B.n718 VSUBS 0.006548f
C759 B.n719 VSUBS 0.006548f
C760 B.n720 VSUBS 0.006548f
C761 B.n721 VSUBS 0.006548f
C762 B.n722 VSUBS 0.006548f
C763 B.n723 VSUBS 0.006548f
C764 B.n724 VSUBS 0.006548f
C765 B.n725 VSUBS 0.006548f
C766 B.n726 VSUBS 0.006548f
C767 B.n727 VSUBS 0.006548f
C768 B.n728 VSUBS 0.006548f
C769 B.n729 VSUBS 0.006548f
C770 B.n730 VSUBS 0.006548f
C771 B.n731 VSUBS 0.006548f
C772 B.n732 VSUBS 0.006548f
C773 B.n733 VSUBS 0.006548f
C774 B.n734 VSUBS 0.006548f
C775 B.n735 VSUBS 0.006548f
C776 B.n736 VSUBS 0.006548f
C777 B.n737 VSUBS 0.006548f
C778 B.n738 VSUBS 0.006548f
C779 B.n739 VSUBS 0.006548f
C780 B.n740 VSUBS 0.006548f
C781 B.n741 VSUBS 0.006548f
C782 B.n742 VSUBS 0.006548f
C783 B.n743 VSUBS 0.006548f
C784 B.n744 VSUBS 0.006548f
C785 B.n745 VSUBS 0.006548f
C786 B.n746 VSUBS 0.006548f
C787 B.n747 VSUBS 0.006548f
C788 B.n748 VSUBS 0.006548f
C789 B.n749 VSUBS 0.006548f
C790 B.n750 VSUBS 0.006548f
C791 B.n751 VSUBS 0.006548f
C792 B.n752 VSUBS 0.006548f
C793 B.n753 VSUBS 0.006548f
C794 B.n754 VSUBS 0.006548f
C795 B.n755 VSUBS 0.006548f
C796 B.n756 VSUBS 0.006548f
C797 B.n757 VSUBS 0.006548f
C798 B.n758 VSUBS 0.006548f
C799 B.n759 VSUBS 0.006548f
C800 B.n760 VSUBS 0.006548f
C801 B.n761 VSUBS 0.006548f
C802 B.n762 VSUBS 0.006548f
C803 B.n763 VSUBS 0.006548f
C804 B.n764 VSUBS 0.006548f
C805 B.n765 VSUBS 0.006548f
C806 B.n766 VSUBS 0.006548f
C807 B.n767 VSUBS 0.006548f
C808 B.n768 VSUBS 0.006548f
C809 B.n769 VSUBS 0.006548f
C810 B.n770 VSUBS 0.006548f
C811 B.n771 VSUBS 0.006548f
C812 B.n772 VSUBS 0.006548f
C813 B.n773 VSUBS 0.006548f
C814 B.n774 VSUBS 0.006548f
C815 B.n775 VSUBS 0.006548f
C816 B.n776 VSUBS 0.006548f
C817 B.n777 VSUBS 0.006548f
C818 B.n778 VSUBS 0.006548f
C819 B.n779 VSUBS 0.006548f
C820 B.n780 VSUBS 0.006548f
C821 B.n781 VSUBS 0.006548f
C822 B.n782 VSUBS 0.006548f
C823 B.n783 VSUBS 0.006548f
C824 B.n784 VSUBS 0.006548f
C825 B.n785 VSUBS 0.006548f
C826 B.n786 VSUBS 0.006548f
C827 B.n787 VSUBS 0.006548f
C828 B.n788 VSUBS 0.006548f
C829 B.n789 VSUBS 0.006548f
C830 B.n790 VSUBS 0.006548f
C831 B.n791 VSUBS 0.006548f
C832 B.n792 VSUBS 0.006548f
C833 B.n793 VSUBS 0.006548f
C834 B.n794 VSUBS 0.006548f
C835 B.n795 VSUBS 0.006548f
C836 B.n796 VSUBS 0.006548f
C837 B.n797 VSUBS 0.006548f
C838 B.n798 VSUBS 0.006548f
C839 B.n799 VSUBS 0.006548f
C840 B.n800 VSUBS 0.006548f
C841 B.n801 VSUBS 0.006548f
C842 B.n802 VSUBS 0.006548f
C843 B.n803 VSUBS 0.006548f
C844 B.n804 VSUBS 0.006548f
C845 B.n805 VSUBS 0.006548f
C846 B.n806 VSUBS 0.006548f
C847 B.n807 VSUBS 0.006548f
C848 B.n808 VSUBS 0.015001f
C849 B.n809 VSUBS 0.015001f
C850 B.n810 VSUBS 0.014081f
C851 B.n811 VSUBS 0.006548f
C852 B.n812 VSUBS 0.006548f
C853 B.n813 VSUBS 0.006548f
C854 B.n814 VSUBS 0.006548f
C855 B.n815 VSUBS 0.006548f
C856 B.n816 VSUBS 0.006548f
C857 B.n817 VSUBS 0.006548f
C858 B.n818 VSUBS 0.006548f
C859 B.n819 VSUBS 0.006548f
C860 B.n820 VSUBS 0.006548f
C861 B.n821 VSUBS 0.006548f
C862 B.n822 VSUBS 0.006548f
C863 B.n823 VSUBS 0.006548f
C864 B.n824 VSUBS 0.006548f
C865 B.n825 VSUBS 0.006548f
C866 B.n826 VSUBS 0.006548f
C867 B.n827 VSUBS 0.006548f
C868 B.n828 VSUBS 0.006548f
C869 B.n829 VSUBS 0.006548f
C870 B.n830 VSUBS 0.006548f
C871 B.n831 VSUBS 0.006548f
C872 B.n832 VSUBS 0.006548f
C873 B.n833 VSUBS 0.006548f
C874 B.n834 VSUBS 0.006548f
C875 B.n835 VSUBS 0.006548f
C876 B.n836 VSUBS 0.006548f
C877 B.n837 VSUBS 0.006548f
C878 B.n838 VSUBS 0.006548f
C879 B.n839 VSUBS 0.006548f
C880 B.n840 VSUBS 0.006548f
C881 B.n841 VSUBS 0.006548f
C882 B.n842 VSUBS 0.006548f
C883 B.n843 VSUBS 0.006548f
C884 B.n844 VSUBS 0.006548f
C885 B.n845 VSUBS 0.006548f
C886 B.n846 VSUBS 0.006548f
C887 B.n847 VSUBS 0.006548f
C888 B.n848 VSUBS 0.006548f
C889 B.n849 VSUBS 0.006548f
C890 B.n850 VSUBS 0.006548f
C891 B.n851 VSUBS 0.006548f
C892 B.n852 VSUBS 0.006548f
C893 B.n853 VSUBS 0.006548f
C894 B.n854 VSUBS 0.006548f
C895 B.n855 VSUBS 0.006548f
C896 B.n856 VSUBS 0.006548f
C897 B.n857 VSUBS 0.006548f
C898 B.n858 VSUBS 0.006548f
C899 B.n859 VSUBS 0.006548f
C900 B.n860 VSUBS 0.006548f
C901 B.n861 VSUBS 0.006548f
C902 B.n862 VSUBS 0.006548f
C903 B.n863 VSUBS 0.006548f
C904 B.n864 VSUBS 0.006548f
C905 B.n865 VSUBS 0.006548f
C906 B.n866 VSUBS 0.006548f
C907 B.n867 VSUBS 0.008545f
C908 B.n868 VSUBS 0.009103f
C909 B.n869 VSUBS 0.018101f
C910 VDD2.t6 VSUBS 0.374614f
C911 VDD2.t4 VSUBS 0.374614f
C912 VDD2.n0 VSUBS 3.16392f
C913 VDD2.t3 VSUBS 0.374614f
C914 VDD2.t0 VSUBS 0.374614f
C915 VDD2.n1 VSUBS 3.16392f
C916 VDD2.n2 VSUBS 3.76565f
C917 VDD2.t1 VSUBS 0.374614f
C918 VDD2.t7 VSUBS 0.374614f
C919 VDD2.n3 VSUBS 3.15556f
C920 VDD2.n4 VSUBS 3.45436f
C921 VDD2.t2 VSUBS 0.374614f
C922 VDD2.t5 VSUBS 0.374614f
C923 VDD2.n5 VSUBS 3.16387f
C924 VN.n0 VSUBS 0.042143f
C925 VN.t7 VSUBS 3.02946f
C926 VN.n1 VSUBS 0.057113f
C927 VN.n2 VSUBS 0.031967f
C928 VN.t4 VSUBS 3.02946f
C929 VN.n3 VSUBS 0.046469f
C930 VN.t1 VSUBS 3.15982f
C931 VN.n4 VSUBS 1.13964f
C932 VN.t3 VSUBS 3.02946f
C933 VN.n5 VSUBS 1.13136f
C934 VN.n6 VSUBS 0.048452f
C935 VN.n7 VSUBS 0.233633f
C936 VN.n8 VSUBS 0.031967f
C937 VN.n9 VSUBS 0.031967f
C938 VN.n10 VSUBS 0.046469f
C939 VN.n11 VSUBS 0.048452f
C940 VN.n12 VSUBS 1.057f
C941 VN.n13 VSUBS 0.040843f
C942 VN.n14 VSUBS 0.031967f
C943 VN.n15 VSUBS 0.031967f
C944 VN.n16 VSUBS 0.031967f
C945 VN.n17 VSUBS 0.032212f
C946 VN.n18 VSUBS 0.059674f
C947 VN.n19 VSUBS 1.14846f
C948 VN.n20 VSUBS 0.036051f
C949 VN.n21 VSUBS 0.042143f
C950 VN.t6 VSUBS 3.02946f
C951 VN.n22 VSUBS 0.057113f
C952 VN.n23 VSUBS 0.031967f
C953 VN.t0 VSUBS 3.02946f
C954 VN.n24 VSUBS 0.046469f
C955 VN.t2 VSUBS 3.15982f
C956 VN.n25 VSUBS 1.13964f
C957 VN.t5 VSUBS 3.02946f
C958 VN.n26 VSUBS 1.13136f
C959 VN.n27 VSUBS 0.048452f
C960 VN.n28 VSUBS 0.233633f
C961 VN.n29 VSUBS 0.031967f
C962 VN.n30 VSUBS 0.031967f
C963 VN.n31 VSUBS 0.046469f
C964 VN.n32 VSUBS 0.048452f
C965 VN.n33 VSUBS 1.057f
C966 VN.n34 VSUBS 0.040843f
C967 VN.n35 VSUBS 0.031967f
C968 VN.n36 VSUBS 0.031967f
C969 VN.n37 VSUBS 0.031967f
C970 VN.n38 VSUBS 0.032212f
C971 VN.n39 VSUBS 0.059674f
C972 VN.n40 VSUBS 1.14846f
C973 VN.n41 VSUBS 1.91171f
C974 VDD1.t6 VSUBS 0.376321f
C975 VDD1.t4 VSUBS 0.376321f
C976 VDD1.n0 VSUBS 3.17956f
C977 VDD1.t0 VSUBS 0.376321f
C978 VDD1.t2 VSUBS 0.376321f
C979 VDD1.n1 VSUBS 3.17834f
C980 VDD1.t3 VSUBS 0.376321f
C981 VDD1.t5 VSUBS 0.376321f
C982 VDD1.n2 VSUBS 3.17834f
C983 VDD1.n3 VSUBS 3.83482f
C984 VDD1.t1 VSUBS 0.376321f
C985 VDD1.t7 VSUBS 0.376321f
C986 VDD1.n4 VSUBS 3.16992f
C987 VDD1.n5 VSUBS 3.50076f
C988 VTAIL.t4 VSUBS 0.348883f
C989 VTAIL.t7 VSUBS 0.348883f
C990 VTAIL.n0 VSUBS 2.80535f
C991 VTAIL.n1 VSUBS 0.682649f
C992 VTAIL.t1 VSUBS 3.65355f
C993 VTAIL.n2 VSUBS 0.816575f
C994 VTAIL.t8 VSUBS 3.65355f
C995 VTAIL.n3 VSUBS 0.816575f
C996 VTAIL.t11 VSUBS 0.348883f
C997 VTAIL.t9 VSUBS 0.348883f
C998 VTAIL.n4 VSUBS 2.80535f
C999 VTAIL.n5 VSUBS 0.81494f
C1000 VTAIL.t14 VSUBS 3.65355f
C1001 VTAIL.n6 VSUBS 2.45828f
C1002 VTAIL.t6 VSUBS 3.65358f
C1003 VTAIL.n7 VSUBS 2.45824f
C1004 VTAIL.t5 VSUBS 0.348883f
C1005 VTAIL.t2 VSUBS 0.348883f
C1006 VTAIL.n8 VSUBS 2.80536f
C1007 VTAIL.n9 VSUBS 0.814923f
C1008 VTAIL.t0 VSUBS 3.65358f
C1009 VTAIL.n10 VSUBS 0.816541f
C1010 VTAIL.t15 VSUBS 3.65358f
C1011 VTAIL.n11 VSUBS 0.816541f
C1012 VTAIL.t10 VSUBS 0.348883f
C1013 VTAIL.t12 VSUBS 0.348883f
C1014 VTAIL.n12 VSUBS 2.80536f
C1015 VTAIL.n13 VSUBS 0.814923f
C1016 VTAIL.t13 VSUBS 3.65355f
C1017 VTAIL.n14 VSUBS 2.45828f
C1018 VTAIL.t3 VSUBS 3.65355f
C1019 VTAIL.n15 VSUBS 2.45395f
C1020 VP.n0 VSUBS 0.04284f
C1021 VP.t2 VSUBS 3.07961f
C1022 VP.n1 VSUBS 0.058058f
C1023 VP.n2 VSUBS 0.032496f
C1024 VP.t4 VSUBS 3.07961f
C1025 VP.n3 VSUBS 0.047238f
C1026 VP.n4 VSUBS 0.032496f
C1027 VP.t5 VSUBS 3.07961f
C1028 VP.n5 VSUBS 0.032745f
C1029 VP.n6 VSUBS 0.04284f
C1030 VP.t0 VSUBS 3.07961f
C1031 VP.n7 VSUBS 0.058058f
C1032 VP.n8 VSUBS 0.032496f
C1033 VP.t6 VSUBS 3.07961f
C1034 VP.n9 VSUBS 0.047238f
C1035 VP.t1 VSUBS 3.21213f
C1036 VP.n10 VSUBS 1.15851f
C1037 VP.t3 VSUBS 3.07961f
C1038 VP.n11 VSUBS 1.15009f
C1039 VP.n12 VSUBS 0.049254f
C1040 VP.n13 VSUBS 0.237501f
C1041 VP.n14 VSUBS 0.032496f
C1042 VP.n15 VSUBS 0.032496f
C1043 VP.n16 VSUBS 0.047238f
C1044 VP.n17 VSUBS 0.049254f
C1045 VP.n18 VSUBS 1.0745f
C1046 VP.n19 VSUBS 0.041519f
C1047 VP.n20 VSUBS 0.032496f
C1048 VP.n21 VSUBS 0.032496f
C1049 VP.n22 VSUBS 0.032496f
C1050 VP.n23 VSUBS 0.032745f
C1051 VP.n24 VSUBS 0.060662f
C1052 VP.n25 VSUBS 1.16747f
C1053 VP.n26 VSUBS 1.92603f
C1054 VP.n27 VSUBS 1.94832f
C1055 VP.t7 VSUBS 3.07961f
C1056 VP.n28 VSUBS 1.16747f
C1057 VP.n29 VSUBS 0.060662f
C1058 VP.n30 VSUBS 0.04284f
C1059 VP.n31 VSUBS 0.032496f
C1060 VP.n32 VSUBS 0.032496f
C1061 VP.n33 VSUBS 0.058058f
C1062 VP.n34 VSUBS 0.041519f
C1063 VP.n35 VSUBS 1.0745f
C1064 VP.n36 VSUBS 0.049254f
C1065 VP.n37 VSUBS 0.032496f
C1066 VP.n38 VSUBS 0.032496f
C1067 VP.n39 VSUBS 0.032496f
C1068 VP.n40 VSUBS 0.047238f
C1069 VP.n41 VSUBS 0.049254f
C1070 VP.n42 VSUBS 1.0745f
C1071 VP.n43 VSUBS 0.041519f
C1072 VP.n44 VSUBS 0.032496f
C1073 VP.n45 VSUBS 0.032496f
C1074 VP.n46 VSUBS 0.032496f
C1075 VP.n47 VSUBS 0.032745f
C1076 VP.n48 VSUBS 0.060662f
C1077 VP.n49 VSUBS 1.16747f
C1078 VP.n50 VSUBS 0.036648f
.ends

