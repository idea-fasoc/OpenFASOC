* NGSPICE file created from diff_pair_sample_0353.ext - technology: sky130A

.subckt diff_pair_sample_0353 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t6 w_n2584_n3996# sky130_fd_pr__pfet_01v8 ad=2.4981 pd=15.47 as=5.9046 ps=31.06 w=15.14 l=2.36
X1 VDD1.t2 VP.t1 VTAIL.t5 w_n2584_n3996# sky130_fd_pr__pfet_01v8 ad=2.4981 pd=15.47 as=5.9046 ps=31.06 w=15.14 l=2.36
X2 VDD2.t3 VN.t0 VTAIL.t7 w_n2584_n3996# sky130_fd_pr__pfet_01v8 ad=2.4981 pd=15.47 as=5.9046 ps=31.06 w=15.14 l=2.36
X3 VTAIL.t4 VP.t2 VDD1.t1 w_n2584_n3996# sky130_fd_pr__pfet_01v8 ad=5.9046 pd=31.06 as=2.4981 ps=15.47 w=15.14 l=2.36
X4 VDD2.t2 VN.t1 VTAIL.t0 w_n2584_n3996# sky130_fd_pr__pfet_01v8 ad=2.4981 pd=15.47 as=5.9046 ps=31.06 w=15.14 l=2.36
X5 VTAIL.t2 VN.t2 VDD2.t1 w_n2584_n3996# sky130_fd_pr__pfet_01v8 ad=5.9046 pd=31.06 as=2.4981 ps=15.47 w=15.14 l=2.36
X6 B.t11 B.t9 B.t10 w_n2584_n3996# sky130_fd_pr__pfet_01v8 ad=5.9046 pd=31.06 as=0 ps=0 w=15.14 l=2.36
X7 B.t8 B.t6 B.t7 w_n2584_n3996# sky130_fd_pr__pfet_01v8 ad=5.9046 pd=31.06 as=0 ps=0 w=15.14 l=2.36
X8 B.t5 B.t3 B.t4 w_n2584_n3996# sky130_fd_pr__pfet_01v8 ad=5.9046 pd=31.06 as=0 ps=0 w=15.14 l=2.36
X9 B.t2 B.t0 B.t1 w_n2584_n3996# sky130_fd_pr__pfet_01v8 ad=5.9046 pd=31.06 as=0 ps=0 w=15.14 l=2.36
X10 VTAIL.t3 VP.t3 VDD1.t0 w_n2584_n3996# sky130_fd_pr__pfet_01v8 ad=5.9046 pd=31.06 as=2.4981 ps=15.47 w=15.14 l=2.36
X11 VTAIL.t1 VN.t3 VDD2.t0 w_n2584_n3996# sky130_fd_pr__pfet_01v8 ad=5.9046 pd=31.06 as=2.4981 ps=15.47 w=15.14 l=2.36
R0 VP.n3 VP.t3 191.392
R1 VP.n3 VP.t0 190.726
R2 VP.n12 VP.n0 161.3
R3 VP.n11 VP.n10 161.3
R4 VP.n9 VP.n1 161.3
R5 VP.n8 VP.n7 161.3
R6 VP.n6 VP.n2 161.3
R7 VP.n5 VP.t2 154.608
R8 VP.n13 VP.t1 154.608
R9 VP.n5 VP.n4 93.9399
R10 VP.n14 VP.n13 93.9399
R11 VP.n4 VP.n3 53.382
R12 VP.n7 VP.n1 40.577
R13 VP.n11 VP.n1 40.577
R14 VP.n7 VP.n6 24.5923
R15 VP.n12 VP.n11 24.5923
R16 VP.n6 VP.n5 16.9689
R17 VP.n13 VP.n12 16.9689
R18 VP.n4 VP.n2 0.278335
R19 VP.n14 VP.n0 0.278335
R20 VP.n8 VP.n2 0.189894
R21 VP.n9 VP.n8 0.189894
R22 VP.n10 VP.n9 0.189894
R23 VP.n10 VP.n0 0.189894
R24 VP VP.n14 0.153485
R25 VTAIL.n5 VTAIL.t3 58.6885
R26 VTAIL.n4 VTAIL.t0 58.6885
R27 VTAIL.n3 VTAIL.t2 58.6885
R28 VTAIL.n7 VTAIL.t7 58.6882
R29 VTAIL.n0 VTAIL.t1 58.6882
R30 VTAIL.n1 VTAIL.t5 58.6882
R31 VTAIL.n2 VTAIL.t4 58.6882
R32 VTAIL.n6 VTAIL.t6 58.6882
R33 VTAIL.n7 VTAIL.n6 27.7376
R34 VTAIL.n3 VTAIL.n2 27.7376
R35 VTAIL.n4 VTAIL.n3 2.31947
R36 VTAIL.n6 VTAIL.n5 2.31947
R37 VTAIL.n2 VTAIL.n1 2.31947
R38 VTAIL VTAIL.n0 1.21817
R39 VTAIL VTAIL.n7 1.10179
R40 VTAIL.n5 VTAIL.n4 0.470328
R41 VTAIL.n1 VTAIL.n0 0.470328
R42 VDD1 VDD1.n1 117.469
R43 VDD1 VDD1.n0 73.2783
R44 VDD1.n0 VDD1.t0 2.14746
R45 VDD1.n0 VDD1.t3 2.14746
R46 VDD1.n1 VDD1.t1 2.14746
R47 VDD1.n1 VDD1.t2 2.14746
R48 VN.n0 VN.t3 191.392
R49 VN.n1 VN.t1 191.392
R50 VN.n0 VN.t0 190.726
R51 VN.n1 VN.t2 190.726
R52 VN VN.n1 53.6608
R53 VN VN.n0 5.39185
R54 VDD2.n2 VDD2.n0 116.944
R55 VDD2.n2 VDD2.n1 73.2201
R56 VDD2.n1 VDD2.t1 2.14746
R57 VDD2.n1 VDD2.t2 2.14746
R58 VDD2.n0 VDD2.t0 2.14746
R59 VDD2.n0 VDD2.t3 2.14746
R60 VDD2 VDD2.n2 0.0586897
R61 B.n499 B.n498 585
R62 B.n500 B.n77 585
R63 B.n502 B.n501 585
R64 B.n503 B.n76 585
R65 B.n505 B.n504 585
R66 B.n506 B.n75 585
R67 B.n508 B.n507 585
R68 B.n509 B.n74 585
R69 B.n511 B.n510 585
R70 B.n512 B.n73 585
R71 B.n514 B.n513 585
R72 B.n515 B.n72 585
R73 B.n517 B.n516 585
R74 B.n518 B.n71 585
R75 B.n520 B.n519 585
R76 B.n521 B.n70 585
R77 B.n523 B.n522 585
R78 B.n524 B.n69 585
R79 B.n526 B.n525 585
R80 B.n527 B.n68 585
R81 B.n529 B.n528 585
R82 B.n530 B.n67 585
R83 B.n532 B.n531 585
R84 B.n533 B.n66 585
R85 B.n535 B.n534 585
R86 B.n536 B.n65 585
R87 B.n538 B.n537 585
R88 B.n539 B.n64 585
R89 B.n541 B.n540 585
R90 B.n542 B.n63 585
R91 B.n544 B.n543 585
R92 B.n545 B.n62 585
R93 B.n547 B.n546 585
R94 B.n548 B.n61 585
R95 B.n550 B.n549 585
R96 B.n551 B.n60 585
R97 B.n553 B.n552 585
R98 B.n554 B.n59 585
R99 B.n556 B.n555 585
R100 B.n557 B.n58 585
R101 B.n559 B.n558 585
R102 B.n560 B.n57 585
R103 B.n562 B.n561 585
R104 B.n563 B.n56 585
R105 B.n565 B.n564 585
R106 B.n566 B.n55 585
R107 B.n568 B.n567 585
R108 B.n569 B.n54 585
R109 B.n571 B.n570 585
R110 B.n572 B.n53 585
R111 B.n574 B.n573 585
R112 B.n576 B.n575 585
R113 B.n577 B.n49 585
R114 B.n579 B.n578 585
R115 B.n580 B.n48 585
R116 B.n582 B.n581 585
R117 B.n583 B.n47 585
R118 B.n585 B.n584 585
R119 B.n586 B.n46 585
R120 B.n588 B.n587 585
R121 B.n590 B.n43 585
R122 B.n592 B.n591 585
R123 B.n593 B.n42 585
R124 B.n595 B.n594 585
R125 B.n596 B.n41 585
R126 B.n598 B.n597 585
R127 B.n599 B.n40 585
R128 B.n601 B.n600 585
R129 B.n602 B.n39 585
R130 B.n604 B.n603 585
R131 B.n605 B.n38 585
R132 B.n607 B.n606 585
R133 B.n608 B.n37 585
R134 B.n610 B.n609 585
R135 B.n611 B.n36 585
R136 B.n613 B.n612 585
R137 B.n614 B.n35 585
R138 B.n616 B.n615 585
R139 B.n617 B.n34 585
R140 B.n619 B.n618 585
R141 B.n620 B.n33 585
R142 B.n622 B.n621 585
R143 B.n623 B.n32 585
R144 B.n625 B.n624 585
R145 B.n626 B.n31 585
R146 B.n628 B.n627 585
R147 B.n629 B.n30 585
R148 B.n631 B.n630 585
R149 B.n632 B.n29 585
R150 B.n634 B.n633 585
R151 B.n635 B.n28 585
R152 B.n637 B.n636 585
R153 B.n638 B.n27 585
R154 B.n640 B.n639 585
R155 B.n641 B.n26 585
R156 B.n643 B.n642 585
R157 B.n644 B.n25 585
R158 B.n646 B.n645 585
R159 B.n647 B.n24 585
R160 B.n649 B.n648 585
R161 B.n650 B.n23 585
R162 B.n652 B.n651 585
R163 B.n653 B.n22 585
R164 B.n655 B.n654 585
R165 B.n656 B.n21 585
R166 B.n658 B.n657 585
R167 B.n659 B.n20 585
R168 B.n661 B.n660 585
R169 B.n662 B.n19 585
R170 B.n664 B.n663 585
R171 B.n665 B.n18 585
R172 B.n497 B.n78 585
R173 B.n496 B.n495 585
R174 B.n494 B.n79 585
R175 B.n493 B.n492 585
R176 B.n491 B.n80 585
R177 B.n490 B.n489 585
R178 B.n488 B.n81 585
R179 B.n487 B.n486 585
R180 B.n485 B.n82 585
R181 B.n484 B.n483 585
R182 B.n482 B.n83 585
R183 B.n481 B.n480 585
R184 B.n479 B.n84 585
R185 B.n478 B.n477 585
R186 B.n476 B.n85 585
R187 B.n475 B.n474 585
R188 B.n473 B.n86 585
R189 B.n472 B.n471 585
R190 B.n470 B.n87 585
R191 B.n469 B.n468 585
R192 B.n467 B.n88 585
R193 B.n466 B.n465 585
R194 B.n464 B.n89 585
R195 B.n463 B.n462 585
R196 B.n461 B.n90 585
R197 B.n460 B.n459 585
R198 B.n458 B.n91 585
R199 B.n457 B.n456 585
R200 B.n455 B.n92 585
R201 B.n454 B.n453 585
R202 B.n452 B.n93 585
R203 B.n451 B.n450 585
R204 B.n449 B.n94 585
R205 B.n448 B.n447 585
R206 B.n446 B.n95 585
R207 B.n445 B.n444 585
R208 B.n443 B.n96 585
R209 B.n442 B.n441 585
R210 B.n440 B.n97 585
R211 B.n439 B.n438 585
R212 B.n437 B.n98 585
R213 B.n436 B.n435 585
R214 B.n434 B.n99 585
R215 B.n433 B.n432 585
R216 B.n431 B.n100 585
R217 B.n430 B.n429 585
R218 B.n428 B.n101 585
R219 B.n427 B.n426 585
R220 B.n425 B.n102 585
R221 B.n424 B.n423 585
R222 B.n422 B.n103 585
R223 B.n421 B.n420 585
R224 B.n419 B.n104 585
R225 B.n418 B.n417 585
R226 B.n416 B.n105 585
R227 B.n415 B.n414 585
R228 B.n413 B.n106 585
R229 B.n412 B.n411 585
R230 B.n410 B.n107 585
R231 B.n409 B.n408 585
R232 B.n407 B.n108 585
R233 B.n406 B.n405 585
R234 B.n404 B.n109 585
R235 B.n403 B.n402 585
R236 B.n401 B.n110 585
R237 B.n233 B.n170 585
R238 B.n235 B.n234 585
R239 B.n236 B.n169 585
R240 B.n238 B.n237 585
R241 B.n239 B.n168 585
R242 B.n241 B.n240 585
R243 B.n242 B.n167 585
R244 B.n244 B.n243 585
R245 B.n245 B.n166 585
R246 B.n247 B.n246 585
R247 B.n248 B.n165 585
R248 B.n250 B.n249 585
R249 B.n251 B.n164 585
R250 B.n253 B.n252 585
R251 B.n254 B.n163 585
R252 B.n256 B.n255 585
R253 B.n257 B.n162 585
R254 B.n259 B.n258 585
R255 B.n260 B.n161 585
R256 B.n262 B.n261 585
R257 B.n263 B.n160 585
R258 B.n265 B.n264 585
R259 B.n266 B.n159 585
R260 B.n268 B.n267 585
R261 B.n269 B.n158 585
R262 B.n271 B.n270 585
R263 B.n272 B.n157 585
R264 B.n274 B.n273 585
R265 B.n275 B.n156 585
R266 B.n277 B.n276 585
R267 B.n278 B.n155 585
R268 B.n280 B.n279 585
R269 B.n281 B.n154 585
R270 B.n283 B.n282 585
R271 B.n284 B.n153 585
R272 B.n286 B.n285 585
R273 B.n287 B.n152 585
R274 B.n289 B.n288 585
R275 B.n290 B.n151 585
R276 B.n292 B.n291 585
R277 B.n293 B.n150 585
R278 B.n295 B.n294 585
R279 B.n296 B.n149 585
R280 B.n298 B.n297 585
R281 B.n299 B.n148 585
R282 B.n301 B.n300 585
R283 B.n302 B.n147 585
R284 B.n304 B.n303 585
R285 B.n305 B.n146 585
R286 B.n307 B.n306 585
R287 B.n308 B.n143 585
R288 B.n311 B.n310 585
R289 B.n312 B.n142 585
R290 B.n314 B.n313 585
R291 B.n315 B.n141 585
R292 B.n317 B.n316 585
R293 B.n318 B.n140 585
R294 B.n320 B.n319 585
R295 B.n321 B.n139 585
R296 B.n323 B.n322 585
R297 B.n325 B.n324 585
R298 B.n326 B.n135 585
R299 B.n328 B.n327 585
R300 B.n329 B.n134 585
R301 B.n331 B.n330 585
R302 B.n332 B.n133 585
R303 B.n334 B.n333 585
R304 B.n335 B.n132 585
R305 B.n337 B.n336 585
R306 B.n338 B.n131 585
R307 B.n340 B.n339 585
R308 B.n341 B.n130 585
R309 B.n343 B.n342 585
R310 B.n344 B.n129 585
R311 B.n346 B.n345 585
R312 B.n347 B.n128 585
R313 B.n349 B.n348 585
R314 B.n350 B.n127 585
R315 B.n352 B.n351 585
R316 B.n353 B.n126 585
R317 B.n355 B.n354 585
R318 B.n356 B.n125 585
R319 B.n358 B.n357 585
R320 B.n359 B.n124 585
R321 B.n361 B.n360 585
R322 B.n362 B.n123 585
R323 B.n364 B.n363 585
R324 B.n365 B.n122 585
R325 B.n367 B.n366 585
R326 B.n368 B.n121 585
R327 B.n370 B.n369 585
R328 B.n371 B.n120 585
R329 B.n373 B.n372 585
R330 B.n374 B.n119 585
R331 B.n376 B.n375 585
R332 B.n377 B.n118 585
R333 B.n379 B.n378 585
R334 B.n380 B.n117 585
R335 B.n382 B.n381 585
R336 B.n383 B.n116 585
R337 B.n385 B.n384 585
R338 B.n386 B.n115 585
R339 B.n388 B.n387 585
R340 B.n389 B.n114 585
R341 B.n391 B.n390 585
R342 B.n392 B.n113 585
R343 B.n394 B.n393 585
R344 B.n395 B.n112 585
R345 B.n397 B.n396 585
R346 B.n398 B.n111 585
R347 B.n400 B.n399 585
R348 B.n232 B.n231 585
R349 B.n230 B.n171 585
R350 B.n229 B.n228 585
R351 B.n227 B.n172 585
R352 B.n226 B.n225 585
R353 B.n224 B.n173 585
R354 B.n223 B.n222 585
R355 B.n221 B.n174 585
R356 B.n220 B.n219 585
R357 B.n218 B.n175 585
R358 B.n217 B.n216 585
R359 B.n215 B.n176 585
R360 B.n214 B.n213 585
R361 B.n212 B.n177 585
R362 B.n211 B.n210 585
R363 B.n209 B.n178 585
R364 B.n208 B.n207 585
R365 B.n206 B.n179 585
R366 B.n205 B.n204 585
R367 B.n203 B.n180 585
R368 B.n202 B.n201 585
R369 B.n200 B.n181 585
R370 B.n199 B.n198 585
R371 B.n197 B.n182 585
R372 B.n196 B.n195 585
R373 B.n194 B.n183 585
R374 B.n193 B.n192 585
R375 B.n191 B.n184 585
R376 B.n190 B.n189 585
R377 B.n188 B.n185 585
R378 B.n187 B.n186 585
R379 B.n2 B.n0 585
R380 B.n713 B.n1 585
R381 B.n712 B.n711 585
R382 B.n710 B.n3 585
R383 B.n709 B.n708 585
R384 B.n707 B.n4 585
R385 B.n706 B.n705 585
R386 B.n704 B.n5 585
R387 B.n703 B.n702 585
R388 B.n701 B.n6 585
R389 B.n700 B.n699 585
R390 B.n698 B.n7 585
R391 B.n697 B.n696 585
R392 B.n695 B.n8 585
R393 B.n694 B.n693 585
R394 B.n692 B.n9 585
R395 B.n691 B.n690 585
R396 B.n689 B.n10 585
R397 B.n688 B.n687 585
R398 B.n686 B.n11 585
R399 B.n685 B.n684 585
R400 B.n683 B.n12 585
R401 B.n682 B.n681 585
R402 B.n680 B.n13 585
R403 B.n679 B.n678 585
R404 B.n677 B.n14 585
R405 B.n676 B.n675 585
R406 B.n674 B.n15 585
R407 B.n673 B.n672 585
R408 B.n671 B.n16 585
R409 B.n670 B.n669 585
R410 B.n668 B.n17 585
R411 B.n667 B.n666 585
R412 B.n715 B.n714 585
R413 B.n233 B.n232 497.305
R414 B.n666 B.n665 497.305
R415 B.n401 B.n400 497.305
R416 B.n498 B.n497 497.305
R417 B.n136 B.t6 362.262
R418 B.n144 B.t9 362.262
R419 B.n44 B.t0 362.262
R420 B.n50 B.t3 362.262
R421 B.n232 B.n171 163.367
R422 B.n228 B.n171 163.367
R423 B.n228 B.n227 163.367
R424 B.n227 B.n226 163.367
R425 B.n226 B.n173 163.367
R426 B.n222 B.n173 163.367
R427 B.n222 B.n221 163.367
R428 B.n221 B.n220 163.367
R429 B.n220 B.n175 163.367
R430 B.n216 B.n175 163.367
R431 B.n216 B.n215 163.367
R432 B.n215 B.n214 163.367
R433 B.n214 B.n177 163.367
R434 B.n210 B.n177 163.367
R435 B.n210 B.n209 163.367
R436 B.n209 B.n208 163.367
R437 B.n208 B.n179 163.367
R438 B.n204 B.n179 163.367
R439 B.n204 B.n203 163.367
R440 B.n203 B.n202 163.367
R441 B.n202 B.n181 163.367
R442 B.n198 B.n181 163.367
R443 B.n198 B.n197 163.367
R444 B.n197 B.n196 163.367
R445 B.n196 B.n183 163.367
R446 B.n192 B.n183 163.367
R447 B.n192 B.n191 163.367
R448 B.n191 B.n190 163.367
R449 B.n190 B.n185 163.367
R450 B.n186 B.n185 163.367
R451 B.n186 B.n2 163.367
R452 B.n714 B.n2 163.367
R453 B.n714 B.n713 163.367
R454 B.n713 B.n712 163.367
R455 B.n712 B.n3 163.367
R456 B.n708 B.n3 163.367
R457 B.n708 B.n707 163.367
R458 B.n707 B.n706 163.367
R459 B.n706 B.n5 163.367
R460 B.n702 B.n5 163.367
R461 B.n702 B.n701 163.367
R462 B.n701 B.n700 163.367
R463 B.n700 B.n7 163.367
R464 B.n696 B.n7 163.367
R465 B.n696 B.n695 163.367
R466 B.n695 B.n694 163.367
R467 B.n694 B.n9 163.367
R468 B.n690 B.n9 163.367
R469 B.n690 B.n689 163.367
R470 B.n689 B.n688 163.367
R471 B.n688 B.n11 163.367
R472 B.n684 B.n11 163.367
R473 B.n684 B.n683 163.367
R474 B.n683 B.n682 163.367
R475 B.n682 B.n13 163.367
R476 B.n678 B.n13 163.367
R477 B.n678 B.n677 163.367
R478 B.n677 B.n676 163.367
R479 B.n676 B.n15 163.367
R480 B.n672 B.n15 163.367
R481 B.n672 B.n671 163.367
R482 B.n671 B.n670 163.367
R483 B.n670 B.n17 163.367
R484 B.n666 B.n17 163.367
R485 B.n234 B.n233 163.367
R486 B.n234 B.n169 163.367
R487 B.n238 B.n169 163.367
R488 B.n239 B.n238 163.367
R489 B.n240 B.n239 163.367
R490 B.n240 B.n167 163.367
R491 B.n244 B.n167 163.367
R492 B.n245 B.n244 163.367
R493 B.n246 B.n245 163.367
R494 B.n246 B.n165 163.367
R495 B.n250 B.n165 163.367
R496 B.n251 B.n250 163.367
R497 B.n252 B.n251 163.367
R498 B.n252 B.n163 163.367
R499 B.n256 B.n163 163.367
R500 B.n257 B.n256 163.367
R501 B.n258 B.n257 163.367
R502 B.n258 B.n161 163.367
R503 B.n262 B.n161 163.367
R504 B.n263 B.n262 163.367
R505 B.n264 B.n263 163.367
R506 B.n264 B.n159 163.367
R507 B.n268 B.n159 163.367
R508 B.n269 B.n268 163.367
R509 B.n270 B.n269 163.367
R510 B.n270 B.n157 163.367
R511 B.n274 B.n157 163.367
R512 B.n275 B.n274 163.367
R513 B.n276 B.n275 163.367
R514 B.n276 B.n155 163.367
R515 B.n280 B.n155 163.367
R516 B.n281 B.n280 163.367
R517 B.n282 B.n281 163.367
R518 B.n282 B.n153 163.367
R519 B.n286 B.n153 163.367
R520 B.n287 B.n286 163.367
R521 B.n288 B.n287 163.367
R522 B.n288 B.n151 163.367
R523 B.n292 B.n151 163.367
R524 B.n293 B.n292 163.367
R525 B.n294 B.n293 163.367
R526 B.n294 B.n149 163.367
R527 B.n298 B.n149 163.367
R528 B.n299 B.n298 163.367
R529 B.n300 B.n299 163.367
R530 B.n300 B.n147 163.367
R531 B.n304 B.n147 163.367
R532 B.n305 B.n304 163.367
R533 B.n306 B.n305 163.367
R534 B.n306 B.n143 163.367
R535 B.n311 B.n143 163.367
R536 B.n312 B.n311 163.367
R537 B.n313 B.n312 163.367
R538 B.n313 B.n141 163.367
R539 B.n317 B.n141 163.367
R540 B.n318 B.n317 163.367
R541 B.n319 B.n318 163.367
R542 B.n319 B.n139 163.367
R543 B.n323 B.n139 163.367
R544 B.n324 B.n323 163.367
R545 B.n324 B.n135 163.367
R546 B.n328 B.n135 163.367
R547 B.n329 B.n328 163.367
R548 B.n330 B.n329 163.367
R549 B.n330 B.n133 163.367
R550 B.n334 B.n133 163.367
R551 B.n335 B.n334 163.367
R552 B.n336 B.n335 163.367
R553 B.n336 B.n131 163.367
R554 B.n340 B.n131 163.367
R555 B.n341 B.n340 163.367
R556 B.n342 B.n341 163.367
R557 B.n342 B.n129 163.367
R558 B.n346 B.n129 163.367
R559 B.n347 B.n346 163.367
R560 B.n348 B.n347 163.367
R561 B.n348 B.n127 163.367
R562 B.n352 B.n127 163.367
R563 B.n353 B.n352 163.367
R564 B.n354 B.n353 163.367
R565 B.n354 B.n125 163.367
R566 B.n358 B.n125 163.367
R567 B.n359 B.n358 163.367
R568 B.n360 B.n359 163.367
R569 B.n360 B.n123 163.367
R570 B.n364 B.n123 163.367
R571 B.n365 B.n364 163.367
R572 B.n366 B.n365 163.367
R573 B.n366 B.n121 163.367
R574 B.n370 B.n121 163.367
R575 B.n371 B.n370 163.367
R576 B.n372 B.n371 163.367
R577 B.n372 B.n119 163.367
R578 B.n376 B.n119 163.367
R579 B.n377 B.n376 163.367
R580 B.n378 B.n377 163.367
R581 B.n378 B.n117 163.367
R582 B.n382 B.n117 163.367
R583 B.n383 B.n382 163.367
R584 B.n384 B.n383 163.367
R585 B.n384 B.n115 163.367
R586 B.n388 B.n115 163.367
R587 B.n389 B.n388 163.367
R588 B.n390 B.n389 163.367
R589 B.n390 B.n113 163.367
R590 B.n394 B.n113 163.367
R591 B.n395 B.n394 163.367
R592 B.n396 B.n395 163.367
R593 B.n396 B.n111 163.367
R594 B.n400 B.n111 163.367
R595 B.n402 B.n401 163.367
R596 B.n402 B.n109 163.367
R597 B.n406 B.n109 163.367
R598 B.n407 B.n406 163.367
R599 B.n408 B.n407 163.367
R600 B.n408 B.n107 163.367
R601 B.n412 B.n107 163.367
R602 B.n413 B.n412 163.367
R603 B.n414 B.n413 163.367
R604 B.n414 B.n105 163.367
R605 B.n418 B.n105 163.367
R606 B.n419 B.n418 163.367
R607 B.n420 B.n419 163.367
R608 B.n420 B.n103 163.367
R609 B.n424 B.n103 163.367
R610 B.n425 B.n424 163.367
R611 B.n426 B.n425 163.367
R612 B.n426 B.n101 163.367
R613 B.n430 B.n101 163.367
R614 B.n431 B.n430 163.367
R615 B.n432 B.n431 163.367
R616 B.n432 B.n99 163.367
R617 B.n436 B.n99 163.367
R618 B.n437 B.n436 163.367
R619 B.n438 B.n437 163.367
R620 B.n438 B.n97 163.367
R621 B.n442 B.n97 163.367
R622 B.n443 B.n442 163.367
R623 B.n444 B.n443 163.367
R624 B.n444 B.n95 163.367
R625 B.n448 B.n95 163.367
R626 B.n449 B.n448 163.367
R627 B.n450 B.n449 163.367
R628 B.n450 B.n93 163.367
R629 B.n454 B.n93 163.367
R630 B.n455 B.n454 163.367
R631 B.n456 B.n455 163.367
R632 B.n456 B.n91 163.367
R633 B.n460 B.n91 163.367
R634 B.n461 B.n460 163.367
R635 B.n462 B.n461 163.367
R636 B.n462 B.n89 163.367
R637 B.n466 B.n89 163.367
R638 B.n467 B.n466 163.367
R639 B.n468 B.n467 163.367
R640 B.n468 B.n87 163.367
R641 B.n472 B.n87 163.367
R642 B.n473 B.n472 163.367
R643 B.n474 B.n473 163.367
R644 B.n474 B.n85 163.367
R645 B.n478 B.n85 163.367
R646 B.n479 B.n478 163.367
R647 B.n480 B.n479 163.367
R648 B.n480 B.n83 163.367
R649 B.n484 B.n83 163.367
R650 B.n485 B.n484 163.367
R651 B.n486 B.n485 163.367
R652 B.n486 B.n81 163.367
R653 B.n490 B.n81 163.367
R654 B.n491 B.n490 163.367
R655 B.n492 B.n491 163.367
R656 B.n492 B.n79 163.367
R657 B.n496 B.n79 163.367
R658 B.n497 B.n496 163.367
R659 B.n665 B.n664 163.367
R660 B.n664 B.n19 163.367
R661 B.n660 B.n19 163.367
R662 B.n660 B.n659 163.367
R663 B.n659 B.n658 163.367
R664 B.n658 B.n21 163.367
R665 B.n654 B.n21 163.367
R666 B.n654 B.n653 163.367
R667 B.n653 B.n652 163.367
R668 B.n652 B.n23 163.367
R669 B.n648 B.n23 163.367
R670 B.n648 B.n647 163.367
R671 B.n647 B.n646 163.367
R672 B.n646 B.n25 163.367
R673 B.n642 B.n25 163.367
R674 B.n642 B.n641 163.367
R675 B.n641 B.n640 163.367
R676 B.n640 B.n27 163.367
R677 B.n636 B.n27 163.367
R678 B.n636 B.n635 163.367
R679 B.n635 B.n634 163.367
R680 B.n634 B.n29 163.367
R681 B.n630 B.n29 163.367
R682 B.n630 B.n629 163.367
R683 B.n629 B.n628 163.367
R684 B.n628 B.n31 163.367
R685 B.n624 B.n31 163.367
R686 B.n624 B.n623 163.367
R687 B.n623 B.n622 163.367
R688 B.n622 B.n33 163.367
R689 B.n618 B.n33 163.367
R690 B.n618 B.n617 163.367
R691 B.n617 B.n616 163.367
R692 B.n616 B.n35 163.367
R693 B.n612 B.n35 163.367
R694 B.n612 B.n611 163.367
R695 B.n611 B.n610 163.367
R696 B.n610 B.n37 163.367
R697 B.n606 B.n37 163.367
R698 B.n606 B.n605 163.367
R699 B.n605 B.n604 163.367
R700 B.n604 B.n39 163.367
R701 B.n600 B.n39 163.367
R702 B.n600 B.n599 163.367
R703 B.n599 B.n598 163.367
R704 B.n598 B.n41 163.367
R705 B.n594 B.n41 163.367
R706 B.n594 B.n593 163.367
R707 B.n593 B.n592 163.367
R708 B.n592 B.n43 163.367
R709 B.n587 B.n43 163.367
R710 B.n587 B.n586 163.367
R711 B.n586 B.n585 163.367
R712 B.n585 B.n47 163.367
R713 B.n581 B.n47 163.367
R714 B.n581 B.n580 163.367
R715 B.n580 B.n579 163.367
R716 B.n579 B.n49 163.367
R717 B.n575 B.n49 163.367
R718 B.n575 B.n574 163.367
R719 B.n574 B.n53 163.367
R720 B.n570 B.n53 163.367
R721 B.n570 B.n569 163.367
R722 B.n569 B.n568 163.367
R723 B.n568 B.n55 163.367
R724 B.n564 B.n55 163.367
R725 B.n564 B.n563 163.367
R726 B.n563 B.n562 163.367
R727 B.n562 B.n57 163.367
R728 B.n558 B.n57 163.367
R729 B.n558 B.n557 163.367
R730 B.n557 B.n556 163.367
R731 B.n556 B.n59 163.367
R732 B.n552 B.n59 163.367
R733 B.n552 B.n551 163.367
R734 B.n551 B.n550 163.367
R735 B.n550 B.n61 163.367
R736 B.n546 B.n61 163.367
R737 B.n546 B.n545 163.367
R738 B.n545 B.n544 163.367
R739 B.n544 B.n63 163.367
R740 B.n540 B.n63 163.367
R741 B.n540 B.n539 163.367
R742 B.n539 B.n538 163.367
R743 B.n538 B.n65 163.367
R744 B.n534 B.n65 163.367
R745 B.n534 B.n533 163.367
R746 B.n533 B.n532 163.367
R747 B.n532 B.n67 163.367
R748 B.n528 B.n67 163.367
R749 B.n528 B.n527 163.367
R750 B.n527 B.n526 163.367
R751 B.n526 B.n69 163.367
R752 B.n522 B.n69 163.367
R753 B.n522 B.n521 163.367
R754 B.n521 B.n520 163.367
R755 B.n520 B.n71 163.367
R756 B.n516 B.n71 163.367
R757 B.n516 B.n515 163.367
R758 B.n515 B.n514 163.367
R759 B.n514 B.n73 163.367
R760 B.n510 B.n73 163.367
R761 B.n510 B.n509 163.367
R762 B.n509 B.n508 163.367
R763 B.n508 B.n75 163.367
R764 B.n504 B.n75 163.367
R765 B.n504 B.n503 163.367
R766 B.n503 B.n502 163.367
R767 B.n502 B.n77 163.367
R768 B.n498 B.n77 163.367
R769 B.n136 B.t8 162.202
R770 B.n50 B.t4 162.202
R771 B.n144 B.t11 162.183
R772 B.n44 B.t1 162.183
R773 B.n137 B.t7 110.032
R774 B.n51 B.t5 110.032
R775 B.n145 B.t10 110.013
R776 B.n45 B.t2 110.013
R777 B.n138 B.n137 59.5399
R778 B.n309 B.n145 59.5399
R779 B.n589 B.n45 59.5399
R780 B.n52 B.n51 59.5399
R781 B.n137 B.n136 52.1702
R782 B.n145 B.n144 52.1702
R783 B.n45 B.n44 52.1702
R784 B.n51 B.n50 52.1702
R785 B.n667 B.n18 32.3127
R786 B.n499 B.n78 32.3127
R787 B.n399 B.n110 32.3127
R788 B.n231 B.n170 32.3127
R789 B B.n715 18.0485
R790 B.n663 B.n18 10.6151
R791 B.n663 B.n662 10.6151
R792 B.n662 B.n661 10.6151
R793 B.n661 B.n20 10.6151
R794 B.n657 B.n20 10.6151
R795 B.n657 B.n656 10.6151
R796 B.n656 B.n655 10.6151
R797 B.n655 B.n22 10.6151
R798 B.n651 B.n22 10.6151
R799 B.n651 B.n650 10.6151
R800 B.n650 B.n649 10.6151
R801 B.n649 B.n24 10.6151
R802 B.n645 B.n24 10.6151
R803 B.n645 B.n644 10.6151
R804 B.n644 B.n643 10.6151
R805 B.n643 B.n26 10.6151
R806 B.n639 B.n26 10.6151
R807 B.n639 B.n638 10.6151
R808 B.n638 B.n637 10.6151
R809 B.n637 B.n28 10.6151
R810 B.n633 B.n28 10.6151
R811 B.n633 B.n632 10.6151
R812 B.n632 B.n631 10.6151
R813 B.n631 B.n30 10.6151
R814 B.n627 B.n30 10.6151
R815 B.n627 B.n626 10.6151
R816 B.n626 B.n625 10.6151
R817 B.n625 B.n32 10.6151
R818 B.n621 B.n32 10.6151
R819 B.n621 B.n620 10.6151
R820 B.n620 B.n619 10.6151
R821 B.n619 B.n34 10.6151
R822 B.n615 B.n34 10.6151
R823 B.n615 B.n614 10.6151
R824 B.n614 B.n613 10.6151
R825 B.n613 B.n36 10.6151
R826 B.n609 B.n36 10.6151
R827 B.n609 B.n608 10.6151
R828 B.n608 B.n607 10.6151
R829 B.n607 B.n38 10.6151
R830 B.n603 B.n38 10.6151
R831 B.n603 B.n602 10.6151
R832 B.n602 B.n601 10.6151
R833 B.n601 B.n40 10.6151
R834 B.n597 B.n40 10.6151
R835 B.n597 B.n596 10.6151
R836 B.n596 B.n595 10.6151
R837 B.n595 B.n42 10.6151
R838 B.n591 B.n42 10.6151
R839 B.n591 B.n590 10.6151
R840 B.n588 B.n46 10.6151
R841 B.n584 B.n46 10.6151
R842 B.n584 B.n583 10.6151
R843 B.n583 B.n582 10.6151
R844 B.n582 B.n48 10.6151
R845 B.n578 B.n48 10.6151
R846 B.n578 B.n577 10.6151
R847 B.n577 B.n576 10.6151
R848 B.n573 B.n572 10.6151
R849 B.n572 B.n571 10.6151
R850 B.n571 B.n54 10.6151
R851 B.n567 B.n54 10.6151
R852 B.n567 B.n566 10.6151
R853 B.n566 B.n565 10.6151
R854 B.n565 B.n56 10.6151
R855 B.n561 B.n56 10.6151
R856 B.n561 B.n560 10.6151
R857 B.n560 B.n559 10.6151
R858 B.n559 B.n58 10.6151
R859 B.n555 B.n58 10.6151
R860 B.n555 B.n554 10.6151
R861 B.n554 B.n553 10.6151
R862 B.n553 B.n60 10.6151
R863 B.n549 B.n60 10.6151
R864 B.n549 B.n548 10.6151
R865 B.n548 B.n547 10.6151
R866 B.n547 B.n62 10.6151
R867 B.n543 B.n62 10.6151
R868 B.n543 B.n542 10.6151
R869 B.n542 B.n541 10.6151
R870 B.n541 B.n64 10.6151
R871 B.n537 B.n64 10.6151
R872 B.n537 B.n536 10.6151
R873 B.n536 B.n535 10.6151
R874 B.n535 B.n66 10.6151
R875 B.n531 B.n66 10.6151
R876 B.n531 B.n530 10.6151
R877 B.n530 B.n529 10.6151
R878 B.n529 B.n68 10.6151
R879 B.n525 B.n68 10.6151
R880 B.n525 B.n524 10.6151
R881 B.n524 B.n523 10.6151
R882 B.n523 B.n70 10.6151
R883 B.n519 B.n70 10.6151
R884 B.n519 B.n518 10.6151
R885 B.n518 B.n517 10.6151
R886 B.n517 B.n72 10.6151
R887 B.n513 B.n72 10.6151
R888 B.n513 B.n512 10.6151
R889 B.n512 B.n511 10.6151
R890 B.n511 B.n74 10.6151
R891 B.n507 B.n74 10.6151
R892 B.n507 B.n506 10.6151
R893 B.n506 B.n505 10.6151
R894 B.n505 B.n76 10.6151
R895 B.n501 B.n76 10.6151
R896 B.n501 B.n500 10.6151
R897 B.n500 B.n499 10.6151
R898 B.n403 B.n110 10.6151
R899 B.n404 B.n403 10.6151
R900 B.n405 B.n404 10.6151
R901 B.n405 B.n108 10.6151
R902 B.n409 B.n108 10.6151
R903 B.n410 B.n409 10.6151
R904 B.n411 B.n410 10.6151
R905 B.n411 B.n106 10.6151
R906 B.n415 B.n106 10.6151
R907 B.n416 B.n415 10.6151
R908 B.n417 B.n416 10.6151
R909 B.n417 B.n104 10.6151
R910 B.n421 B.n104 10.6151
R911 B.n422 B.n421 10.6151
R912 B.n423 B.n422 10.6151
R913 B.n423 B.n102 10.6151
R914 B.n427 B.n102 10.6151
R915 B.n428 B.n427 10.6151
R916 B.n429 B.n428 10.6151
R917 B.n429 B.n100 10.6151
R918 B.n433 B.n100 10.6151
R919 B.n434 B.n433 10.6151
R920 B.n435 B.n434 10.6151
R921 B.n435 B.n98 10.6151
R922 B.n439 B.n98 10.6151
R923 B.n440 B.n439 10.6151
R924 B.n441 B.n440 10.6151
R925 B.n441 B.n96 10.6151
R926 B.n445 B.n96 10.6151
R927 B.n446 B.n445 10.6151
R928 B.n447 B.n446 10.6151
R929 B.n447 B.n94 10.6151
R930 B.n451 B.n94 10.6151
R931 B.n452 B.n451 10.6151
R932 B.n453 B.n452 10.6151
R933 B.n453 B.n92 10.6151
R934 B.n457 B.n92 10.6151
R935 B.n458 B.n457 10.6151
R936 B.n459 B.n458 10.6151
R937 B.n459 B.n90 10.6151
R938 B.n463 B.n90 10.6151
R939 B.n464 B.n463 10.6151
R940 B.n465 B.n464 10.6151
R941 B.n465 B.n88 10.6151
R942 B.n469 B.n88 10.6151
R943 B.n470 B.n469 10.6151
R944 B.n471 B.n470 10.6151
R945 B.n471 B.n86 10.6151
R946 B.n475 B.n86 10.6151
R947 B.n476 B.n475 10.6151
R948 B.n477 B.n476 10.6151
R949 B.n477 B.n84 10.6151
R950 B.n481 B.n84 10.6151
R951 B.n482 B.n481 10.6151
R952 B.n483 B.n482 10.6151
R953 B.n483 B.n82 10.6151
R954 B.n487 B.n82 10.6151
R955 B.n488 B.n487 10.6151
R956 B.n489 B.n488 10.6151
R957 B.n489 B.n80 10.6151
R958 B.n493 B.n80 10.6151
R959 B.n494 B.n493 10.6151
R960 B.n495 B.n494 10.6151
R961 B.n495 B.n78 10.6151
R962 B.n235 B.n170 10.6151
R963 B.n236 B.n235 10.6151
R964 B.n237 B.n236 10.6151
R965 B.n237 B.n168 10.6151
R966 B.n241 B.n168 10.6151
R967 B.n242 B.n241 10.6151
R968 B.n243 B.n242 10.6151
R969 B.n243 B.n166 10.6151
R970 B.n247 B.n166 10.6151
R971 B.n248 B.n247 10.6151
R972 B.n249 B.n248 10.6151
R973 B.n249 B.n164 10.6151
R974 B.n253 B.n164 10.6151
R975 B.n254 B.n253 10.6151
R976 B.n255 B.n254 10.6151
R977 B.n255 B.n162 10.6151
R978 B.n259 B.n162 10.6151
R979 B.n260 B.n259 10.6151
R980 B.n261 B.n260 10.6151
R981 B.n261 B.n160 10.6151
R982 B.n265 B.n160 10.6151
R983 B.n266 B.n265 10.6151
R984 B.n267 B.n266 10.6151
R985 B.n267 B.n158 10.6151
R986 B.n271 B.n158 10.6151
R987 B.n272 B.n271 10.6151
R988 B.n273 B.n272 10.6151
R989 B.n273 B.n156 10.6151
R990 B.n277 B.n156 10.6151
R991 B.n278 B.n277 10.6151
R992 B.n279 B.n278 10.6151
R993 B.n279 B.n154 10.6151
R994 B.n283 B.n154 10.6151
R995 B.n284 B.n283 10.6151
R996 B.n285 B.n284 10.6151
R997 B.n285 B.n152 10.6151
R998 B.n289 B.n152 10.6151
R999 B.n290 B.n289 10.6151
R1000 B.n291 B.n290 10.6151
R1001 B.n291 B.n150 10.6151
R1002 B.n295 B.n150 10.6151
R1003 B.n296 B.n295 10.6151
R1004 B.n297 B.n296 10.6151
R1005 B.n297 B.n148 10.6151
R1006 B.n301 B.n148 10.6151
R1007 B.n302 B.n301 10.6151
R1008 B.n303 B.n302 10.6151
R1009 B.n303 B.n146 10.6151
R1010 B.n307 B.n146 10.6151
R1011 B.n308 B.n307 10.6151
R1012 B.n310 B.n142 10.6151
R1013 B.n314 B.n142 10.6151
R1014 B.n315 B.n314 10.6151
R1015 B.n316 B.n315 10.6151
R1016 B.n316 B.n140 10.6151
R1017 B.n320 B.n140 10.6151
R1018 B.n321 B.n320 10.6151
R1019 B.n322 B.n321 10.6151
R1020 B.n326 B.n325 10.6151
R1021 B.n327 B.n326 10.6151
R1022 B.n327 B.n134 10.6151
R1023 B.n331 B.n134 10.6151
R1024 B.n332 B.n331 10.6151
R1025 B.n333 B.n332 10.6151
R1026 B.n333 B.n132 10.6151
R1027 B.n337 B.n132 10.6151
R1028 B.n338 B.n337 10.6151
R1029 B.n339 B.n338 10.6151
R1030 B.n339 B.n130 10.6151
R1031 B.n343 B.n130 10.6151
R1032 B.n344 B.n343 10.6151
R1033 B.n345 B.n344 10.6151
R1034 B.n345 B.n128 10.6151
R1035 B.n349 B.n128 10.6151
R1036 B.n350 B.n349 10.6151
R1037 B.n351 B.n350 10.6151
R1038 B.n351 B.n126 10.6151
R1039 B.n355 B.n126 10.6151
R1040 B.n356 B.n355 10.6151
R1041 B.n357 B.n356 10.6151
R1042 B.n357 B.n124 10.6151
R1043 B.n361 B.n124 10.6151
R1044 B.n362 B.n361 10.6151
R1045 B.n363 B.n362 10.6151
R1046 B.n363 B.n122 10.6151
R1047 B.n367 B.n122 10.6151
R1048 B.n368 B.n367 10.6151
R1049 B.n369 B.n368 10.6151
R1050 B.n369 B.n120 10.6151
R1051 B.n373 B.n120 10.6151
R1052 B.n374 B.n373 10.6151
R1053 B.n375 B.n374 10.6151
R1054 B.n375 B.n118 10.6151
R1055 B.n379 B.n118 10.6151
R1056 B.n380 B.n379 10.6151
R1057 B.n381 B.n380 10.6151
R1058 B.n381 B.n116 10.6151
R1059 B.n385 B.n116 10.6151
R1060 B.n386 B.n385 10.6151
R1061 B.n387 B.n386 10.6151
R1062 B.n387 B.n114 10.6151
R1063 B.n391 B.n114 10.6151
R1064 B.n392 B.n391 10.6151
R1065 B.n393 B.n392 10.6151
R1066 B.n393 B.n112 10.6151
R1067 B.n397 B.n112 10.6151
R1068 B.n398 B.n397 10.6151
R1069 B.n399 B.n398 10.6151
R1070 B.n231 B.n230 10.6151
R1071 B.n230 B.n229 10.6151
R1072 B.n229 B.n172 10.6151
R1073 B.n225 B.n172 10.6151
R1074 B.n225 B.n224 10.6151
R1075 B.n224 B.n223 10.6151
R1076 B.n223 B.n174 10.6151
R1077 B.n219 B.n174 10.6151
R1078 B.n219 B.n218 10.6151
R1079 B.n218 B.n217 10.6151
R1080 B.n217 B.n176 10.6151
R1081 B.n213 B.n176 10.6151
R1082 B.n213 B.n212 10.6151
R1083 B.n212 B.n211 10.6151
R1084 B.n211 B.n178 10.6151
R1085 B.n207 B.n178 10.6151
R1086 B.n207 B.n206 10.6151
R1087 B.n206 B.n205 10.6151
R1088 B.n205 B.n180 10.6151
R1089 B.n201 B.n180 10.6151
R1090 B.n201 B.n200 10.6151
R1091 B.n200 B.n199 10.6151
R1092 B.n199 B.n182 10.6151
R1093 B.n195 B.n182 10.6151
R1094 B.n195 B.n194 10.6151
R1095 B.n194 B.n193 10.6151
R1096 B.n193 B.n184 10.6151
R1097 B.n189 B.n184 10.6151
R1098 B.n189 B.n188 10.6151
R1099 B.n188 B.n187 10.6151
R1100 B.n187 B.n0 10.6151
R1101 B.n711 B.n1 10.6151
R1102 B.n711 B.n710 10.6151
R1103 B.n710 B.n709 10.6151
R1104 B.n709 B.n4 10.6151
R1105 B.n705 B.n4 10.6151
R1106 B.n705 B.n704 10.6151
R1107 B.n704 B.n703 10.6151
R1108 B.n703 B.n6 10.6151
R1109 B.n699 B.n6 10.6151
R1110 B.n699 B.n698 10.6151
R1111 B.n698 B.n697 10.6151
R1112 B.n697 B.n8 10.6151
R1113 B.n693 B.n8 10.6151
R1114 B.n693 B.n692 10.6151
R1115 B.n692 B.n691 10.6151
R1116 B.n691 B.n10 10.6151
R1117 B.n687 B.n10 10.6151
R1118 B.n687 B.n686 10.6151
R1119 B.n686 B.n685 10.6151
R1120 B.n685 B.n12 10.6151
R1121 B.n681 B.n12 10.6151
R1122 B.n681 B.n680 10.6151
R1123 B.n680 B.n679 10.6151
R1124 B.n679 B.n14 10.6151
R1125 B.n675 B.n14 10.6151
R1126 B.n675 B.n674 10.6151
R1127 B.n674 B.n673 10.6151
R1128 B.n673 B.n16 10.6151
R1129 B.n669 B.n16 10.6151
R1130 B.n669 B.n668 10.6151
R1131 B.n668 B.n667 10.6151
R1132 B.n589 B.n588 6.5566
R1133 B.n576 B.n52 6.5566
R1134 B.n310 B.n309 6.5566
R1135 B.n322 B.n138 6.5566
R1136 B.n590 B.n589 4.05904
R1137 B.n573 B.n52 4.05904
R1138 B.n309 B.n308 4.05904
R1139 B.n325 B.n138 4.05904
R1140 B.n715 B.n0 2.81026
R1141 B.n715 B.n1 2.81026
C0 VDD1 w_n2584_n3996# 1.48846f
C1 VDD1 VP 6.03782f
C2 VTAIL w_n2584_n3996# 4.68374f
C3 VDD1 VN 0.148948f
C4 VTAIL VP 5.5576f
C5 VDD1 B 1.30542f
C6 VN VTAIL 5.54349f
C7 VTAIL B 5.85076f
C8 VDD2 w_n2584_n3996# 1.53924f
C9 VDD2 VP 0.379199f
C10 VN VDD2 5.80825f
C11 VDD2 B 1.35361f
C12 VDD1 VTAIL 6.15459f
C13 VP w_n2584_n3996# 4.71398f
C14 VDD1 VDD2 0.972164f
C15 VN w_n2584_n3996# 4.3824f
C16 w_n2584_n3996# B 9.83154f
C17 VN VP 6.59352f
C18 VP B 1.65271f
C19 VDD2 VTAIL 6.20719f
C20 VN B 1.10359f
C21 VDD2 VSUBS 0.9724f
C22 VDD1 VSUBS 5.98867f
C23 VTAIL VSUBS 1.335473f
C24 VN VSUBS 5.45717f
C25 VP VSUBS 2.277239f
C26 B VSUBS 4.328898f
C27 w_n2584_n3996# VSUBS 0.126606p
C28 B.n0 VSUBS 0.00409f
C29 B.n1 VSUBS 0.00409f
C30 B.n2 VSUBS 0.006468f
C31 B.n3 VSUBS 0.006468f
C32 B.n4 VSUBS 0.006468f
C33 B.n5 VSUBS 0.006468f
C34 B.n6 VSUBS 0.006468f
C35 B.n7 VSUBS 0.006468f
C36 B.n8 VSUBS 0.006468f
C37 B.n9 VSUBS 0.006468f
C38 B.n10 VSUBS 0.006468f
C39 B.n11 VSUBS 0.006468f
C40 B.n12 VSUBS 0.006468f
C41 B.n13 VSUBS 0.006468f
C42 B.n14 VSUBS 0.006468f
C43 B.n15 VSUBS 0.006468f
C44 B.n16 VSUBS 0.006468f
C45 B.n17 VSUBS 0.006468f
C46 B.n18 VSUBS 0.015208f
C47 B.n19 VSUBS 0.006468f
C48 B.n20 VSUBS 0.006468f
C49 B.n21 VSUBS 0.006468f
C50 B.n22 VSUBS 0.006468f
C51 B.n23 VSUBS 0.006468f
C52 B.n24 VSUBS 0.006468f
C53 B.n25 VSUBS 0.006468f
C54 B.n26 VSUBS 0.006468f
C55 B.n27 VSUBS 0.006468f
C56 B.n28 VSUBS 0.006468f
C57 B.n29 VSUBS 0.006468f
C58 B.n30 VSUBS 0.006468f
C59 B.n31 VSUBS 0.006468f
C60 B.n32 VSUBS 0.006468f
C61 B.n33 VSUBS 0.006468f
C62 B.n34 VSUBS 0.006468f
C63 B.n35 VSUBS 0.006468f
C64 B.n36 VSUBS 0.006468f
C65 B.n37 VSUBS 0.006468f
C66 B.n38 VSUBS 0.006468f
C67 B.n39 VSUBS 0.006468f
C68 B.n40 VSUBS 0.006468f
C69 B.n41 VSUBS 0.006468f
C70 B.n42 VSUBS 0.006468f
C71 B.n43 VSUBS 0.006468f
C72 B.t2 VSUBS 0.46609f
C73 B.t1 VSUBS 0.484221f
C74 B.t0 VSUBS 1.47117f
C75 B.n44 VSUBS 0.250624f
C76 B.n45 VSUBS 0.065591f
C77 B.n46 VSUBS 0.006468f
C78 B.n47 VSUBS 0.006468f
C79 B.n48 VSUBS 0.006468f
C80 B.n49 VSUBS 0.006468f
C81 B.t5 VSUBS 0.466077f
C82 B.t4 VSUBS 0.48421f
C83 B.t3 VSUBS 1.47117f
C84 B.n50 VSUBS 0.250636f
C85 B.n51 VSUBS 0.065604f
C86 B.n52 VSUBS 0.014986f
C87 B.n53 VSUBS 0.006468f
C88 B.n54 VSUBS 0.006468f
C89 B.n55 VSUBS 0.006468f
C90 B.n56 VSUBS 0.006468f
C91 B.n57 VSUBS 0.006468f
C92 B.n58 VSUBS 0.006468f
C93 B.n59 VSUBS 0.006468f
C94 B.n60 VSUBS 0.006468f
C95 B.n61 VSUBS 0.006468f
C96 B.n62 VSUBS 0.006468f
C97 B.n63 VSUBS 0.006468f
C98 B.n64 VSUBS 0.006468f
C99 B.n65 VSUBS 0.006468f
C100 B.n66 VSUBS 0.006468f
C101 B.n67 VSUBS 0.006468f
C102 B.n68 VSUBS 0.006468f
C103 B.n69 VSUBS 0.006468f
C104 B.n70 VSUBS 0.006468f
C105 B.n71 VSUBS 0.006468f
C106 B.n72 VSUBS 0.006468f
C107 B.n73 VSUBS 0.006468f
C108 B.n74 VSUBS 0.006468f
C109 B.n75 VSUBS 0.006468f
C110 B.n76 VSUBS 0.006468f
C111 B.n77 VSUBS 0.006468f
C112 B.n78 VSUBS 0.015623f
C113 B.n79 VSUBS 0.006468f
C114 B.n80 VSUBS 0.006468f
C115 B.n81 VSUBS 0.006468f
C116 B.n82 VSUBS 0.006468f
C117 B.n83 VSUBS 0.006468f
C118 B.n84 VSUBS 0.006468f
C119 B.n85 VSUBS 0.006468f
C120 B.n86 VSUBS 0.006468f
C121 B.n87 VSUBS 0.006468f
C122 B.n88 VSUBS 0.006468f
C123 B.n89 VSUBS 0.006468f
C124 B.n90 VSUBS 0.006468f
C125 B.n91 VSUBS 0.006468f
C126 B.n92 VSUBS 0.006468f
C127 B.n93 VSUBS 0.006468f
C128 B.n94 VSUBS 0.006468f
C129 B.n95 VSUBS 0.006468f
C130 B.n96 VSUBS 0.006468f
C131 B.n97 VSUBS 0.006468f
C132 B.n98 VSUBS 0.006468f
C133 B.n99 VSUBS 0.006468f
C134 B.n100 VSUBS 0.006468f
C135 B.n101 VSUBS 0.006468f
C136 B.n102 VSUBS 0.006468f
C137 B.n103 VSUBS 0.006468f
C138 B.n104 VSUBS 0.006468f
C139 B.n105 VSUBS 0.006468f
C140 B.n106 VSUBS 0.006468f
C141 B.n107 VSUBS 0.006468f
C142 B.n108 VSUBS 0.006468f
C143 B.n109 VSUBS 0.006468f
C144 B.n110 VSUBS 0.01485f
C145 B.n111 VSUBS 0.006468f
C146 B.n112 VSUBS 0.006468f
C147 B.n113 VSUBS 0.006468f
C148 B.n114 VSUBS 0.006468f
C149 B.n115 VSUBS 0.006468f
C150 B.n116 VSUBS 0.006468f
C151 B.n117 VSUBS 0.006468f
C152 B.n118 VSUBS 0.006468f
C153 B.n119 VSUBS 0.006468f
C154 B.n120 VSUBS 0.006468f
C155 B.n121 VSUBS 0.006468f
C156 B.n122 VSUBS 0.006468f
C157 B.n123 VSUBS 0.006468f
C158 B.n124 VSUBS 0.006468f
C159 B.n125 VSUBS 0.006468f
C160 B.n126 VSUBS 0.006468f
C161 B.n127 VSUBS 0.006468f
C162 B.n128 VSUBS 0.006468f
C163 B.n129 VSUBS 0.006468f
C164 B.n130 VSUBS 0.006468f
C165 B.n131 VSUBS 0.006468f
C166 B.n132 VSUBS 0.006468f
C167 B.n133 VSUBS 0.006468f
C168 B.n134 VSUBS 0.006468f
C169 B.n135 VSUBS 0.006468f
C170 B.t7 VSUBS 0.466077f
C171 B.t8 VSUBS 0.48421f
C172 B.t6 VSUBS 1.47117f
C173 B.n136 VSUBS 0.250636f
C174 B.n137 VSUBS 0.065604f
C175 B.n138 VSUBS 0.014986f
C176 B.n139 VSUBS 0.006468f
C177 B.n140 VSUBS 0.006468f
C178 B.n141 VSUBS 0.006468f
C179 B.n142 VSUBS 0.006468f
C180 B.n143 VSUBS 0.006468f
C181 B.t10 VSUBS 0.46609f
C182 B.t11 VSUBS 0.484221f
C183 B.t9 VSUBS 1.47117f
C184 B.n144 VSUBS 0.250624f
C185 B.n145 VSUBS 0.065591f
C186 B.n146 VSUBS 0.006468f
C187 B.n147 VSUBS 0.006468f
C188 B.n148 VSUBS 0.006468f
C189 B.n149 VSUBS 0.006468f
C190 B.n150 VSUBS 0.006468f
C191 B.n151 VSUBS 0.006468f
C192 B.n152 VSUBS 0.006468f
C193 B.n153 VSUBS 0.006468f
C194 B.n154 VSUBS 0.006468f
C195 B.n155 VSUBS 0.006468f
C196 B.n156 VSUBS 0.006468f
C197 B.n157 VSUBS 0.006468f
C198 B.n158 VSUBS 0.006468f
C199 B.n159 VSUBS 0.006468f
C200 B.n160 VSUBS 0.006468f
C201 B.n161 VSUBS 0.006468f
C202 B.n162 VSUBS 0.006468f
C203 B.n163 VSUBS 0.006468f
C204 B.n164 VSUBS 0.006468f
C205 B.n165 VSUBS 0.006468f
C206 B.n166 VSUBS 0.006468f
C207 B.n167 VSUBS 0.006468f
C208 B.n168 VSUBS 0.006468f
C209 B.n169 VSUBS 0.006468f
C210 B.n170 VSUBS 0.015208f
C211 B.n171 VSUBS 0.006468f
C212 B.n172 VSUBS 0.006468f
C213 B.n173 VSUBS 0.006468f
C214 B.n174 VSUBS 0.006468f
C215 B.n175 VSUBS 0.006468f
C216 B.n176 VSUBS 0.006468f
C217 B.n177 VSUBS 0.006468f
C218 B.n178 VSUBS 0.006468f
C219 B.n179 VSUBS 0.006468f
C220 B.n180 VSUBS 0.006468f
C221 B.n181 VSUBS 0.006468f
C222 B.n182 VSUBS 0.006468f
C223 B.n183 VSUBS 0.006468f
C224 B.n184 VSUBS 0.006468f
C225 B.n185 VSUBS 0.006468f
C226 B.n186 VSUBS 0.006468f
C227 B.n187 VSUBS 0.006468f
C228 B.n188 VSUBS 0.006468f
C229 B.n189 VSUBS 0.006468f
C230 B.n190 VSUBS 0.006468f
C231 B.n191 VSUBS 0.006468f
C232 B.n192 VSUBS 0.006468f
C233 B.n193 VSUBS 0.006468f
C234 B.n194 VSUBS 0.006468f
C235 B.n195 VSUBS 0.006468f
C236 B.n196 VSUBS 0.006468f
C237 B.n197 VSUBS 0.006468f
C238 B.n198 VSUBS 0.006468f
C239 B.n199 VSUBS 0.006468f
C240 B.n200 VSUBS 0.006468f
C241 B.n201 VSUBS 0.006468f
C242 B.n202 VSUBS 0.006468f
C243 B.n203 VSUBS 0.006468f
C244 B.n204 VSUBS 0.006468f
C245 B.n205 VSUBS 0.006468f
C246 B.n206 VSUBS 0.006468f
C247 B.n207 VSUBS 0.006468f
C248 B.n208 VSUBS 0.006468f
C249 B.n209 VSUBS 0.006468f
C250 B.n210 VSUBS 0.006468f
C251 B.n211 VSUBS 0.006468f
C252 B.n212 VSUBS 0.006468f
C253 B.n213 VSUBS 0.006468f
C254 B.n214 VSUBS 0.006468f
C255 B.n215 VSUBS 0.006468f
C256 B.n216 VSUBS 0.006468f
C257 B.n217 VSUBS 0.006468f
C258 B.n218 VSUBS 0.006468f
C259 B.n219 VSUBS 0.006468f
C260 B.n220 VSUBS 0.006468f
C261 B.n221 VSUBS 0.006468f
C262 B.n222 VSUBS 0.006468f
C263 B.n223 VSUBS 0.006468f
C264 B.n224 VSUBS 0.006468f
C265 B.n225 VSUBS 0.006468f
C266 B.n226 VSUBS 0.006468f
C267 B.n227 VSUBS 0.006468f
C268 B.n228 VSUBS 0.006468f
C269 B.n229 VSUBS 0.006468f
C270 B.n230 VSUBS 0.006468f
C271 B.n231 VSUBS 0.01485f
C272 B.n232 VSUBS 0.01485f
C273 B.n233 VSUBS 0.015208f
C274 B.n234 VSUBS 0.006468f
C275 B.n235 VSUBS 0.006468f
C276 B.n236 VSUBS 0.006468f
C277 B.n237 VSUBS 0.006468f
C278 B.n238 VSUBS 0.006468f
C279 B.n239 VSUBS 0.006468f
C280 B.n240 VSUBS 0.006468f
C281 B.n241 VSUBS 0.006468f
C282 B.n242 VSUBS 0.006468f
C283 B.n243 VSUBS 0.006468f
C284 B.n244 VSUBS 0.006468f
C285 B.n245 VSUBS 0.006468f
C286 B.n246 VSUBS 0.006468f
C287 B.n247 VSUBS 0.006468f
C288 B.n248 VSUBS 0.006468f
C289 B.n249 VSUBS 0.006468f
C290 B.n250 VSUBS 0.006468f
C291 B.n251 VSUBS 0.006468f
C292 B.n252 VSUBS 0.006468f
C293 B.n253 VSUBS 0.006468f
C294 B.n254 VSUBS 0.006468f
C295 B.n255 VSUBS 0.006468f
C296 B.n256 VSUBS 0.006468f
C297 B.n257 VSUBS 0.006468f
C298 B.n258 VSUBS 0.006468f
C299 B.n259 VSUBS 0.006468f
C300 B.n260 VSUBS 0.006468f
C301 B.n261 VSUBS 0.006468f
C302 B.n262 VSUBS 0.006468f
C303 B.n263 VSUBS 0.006468f
C304 B.n264 VSUBS 0.006468f
C305 B.n265 VSUBS 0.006468f
C306 B.n266 VSUBS 0.006468f
C307 B.n267 VSUBS 0.006468f
C308 B.n268 VSUBS 0.006468f
C309 B.n269 VSUBS 0.006468f
C310 B.n270 VSUBS 0.006468f
C311 B.n271 VSUBS 0.006468f
C312 B.n272 VSUBS 0.006468f
C313 B.n273 VSUBS 0.006468f
C314 B.n274 VSUBS 0.006468f
C315 B.n275 VSUBS 0.006468f
C316 B.n276 VSUBS 0.006468f
C317 B.n277 VSUBS 0.006468f
C318 B.n278 VSUBS 0.006468f
C319 B.n279 VSUBS 0.006468f
C320 B.n280 VSUBS 0.006468f
C321 B.n281 VSUBS 0.006468f
C322 B.n282 VSUBS 0.006468f
C323 B.n283 VSUBS 0.006468f
C324 B.n284 VSUBS 0.006468f
C325 B.n285 VSUBS 0.006468f
C326 B.n286 VSUBS 0.006468f
C327 B.n287 VSUBS 0.006468f
C328 B.n288 VSUBS 0.006468f
C329 B.n289 VSUBS 0.006468f
C330 B.n290 VSUBS 0.006468f
C331 B.n291 VSUBS 0.006468f
C332 B.n292 VSUBS 0.006468f
C333 B.n293 VSUBS 0.006468f
C334 B.n294 VSUBS 0.006468f
C335 B.n295 VSUBS 0.006468f
C336 B.n296 VSUBS 0.006468f
C337 B.n297 VSUBS 0.006468f
C338 B.n298 VSUBS 0.006468f
C339 B.n299 VSUBS 0.006468f
C340 B.n300 VSUBS 0.006468f
C341 B.n301 VSUBS 0.006468f
C342 B.n302 VSUBS 0.006468f
C343 B.n303 VSUBS 0.006468f
C344 B.n304 VSUBS 0.006468f
C345 B.n305 VSUBS 0.006468f
C346 B.n306 VSUBS 0.006468f
C347 B.n307 VSUBS 0.006468f
C348 B.n308 VSUBS 0.004471f
C349 B.n309 VSUBS 0.014986f
C350 B.n310 VSUBS 0.005232f
C351 B.n311 VSUBS 0.006468f
C352 B.n312 VSUBS 0.006468f
C353 B.n313 VSUBS 0.006468f
C354 B.n314 VSUBS 0.006468f
C355 B.n315 VSUBS 0.006468f
C356 B.n316 VSUBS 0.006468f
C357 B.n317 VSUBS 0.006468f
C358 B.n318 VSUBS 0.006468f
C359 B.n319 VSUBS 0.006468f
C360 B.n320 VSUBS 0.006468f
C361 B.n321 VSUBS 0.006468f
C362 B.n322 VSUBS 0.005232f
C363 B.n323 VSUBS 0.006468f
C364 B.n324 VSUBS 0.006468f
C365 B.n325 VSUBS 0.004471f
C366 B.n326 VSUBS 0.006468f
C367 B.n327 VSUBS 0.006468f
C368 B.n328 VSUBS 0.006468f
C369 B.n329 VSUBS 0.006468f
C370 B.n330 VSUBS 0.006468f
C371 B.n331 VSUBS 0.006468f
C372 B.n332 VSUBS 0.006468f
C373 B.n333 VSUBS 0.006468f
C374 B.n334 VSUBS 0.006468f
C375 B.n335 VSUBS 0.006468f
C376 B.n336 VSUBS 0.006468f
C377 B.n337 VSUBS 0.006468f
C378 B.n338 VSUBS 0.006468f
C379 B.n339 VSUBS 0.006468f
C380 B.n340 VSUBS 0.006468f
C381 B.n341 VSUBS 0.006468f
C382 B.n342 VSUBS 0.006468f
C383 B.n343 VSUBS 0.006468f
C384 B.n344 VSUBS 0.006468f
C385 B.n345 VSUBS 0.006468f
C386 B.n346 VSUBS 0.006468f
C387 B.n347 VSUBS 0.006468f
C388 B.n348 VSUBS 0.006468f
C389 B.n349 VSUBS 0.006468f
C390 B.n350 VSUBS 0.006468f
C391 B.n351 VSUBS 0.006468f
C392 B.n352 VSUBS 0.006468f
C393 B.n353 VSUBS 0.006468f
C394 B.n354 VSUBS 0.006468f
C395 B.n355 VSUBS 0.006468f
C396 B.n356 VSUBS 0.006468f
C397 B.n357 VSUBS 0.006468f
C398 B.n358 VSUBS 0.006468f
C399 B.n359 VSUBS 0.006468f
C400 B.n360 VSUBS 0.006468f
C401 B.n361 VSUBS 0.006468f
C402 B.n362 VSUBS 0.006468f
C403 B.n363 VSUBS 0.006468f
C404 B.n364 VSUBS 0.006468f
C405 B.n365 VSUBS 0.006468f
C406 B.n366 VSUBS 0.006468f
C407 B.n367 VSUBS 0.006468f
C408 B.n368 VSUBS 0.006468f
C409 B.n369 VSUBS 0.006468f
C410 B.n370 VSUBS 0.006468f
C411 B.n371 VSUBS 0.006468f
C412 B.n372 VSUBS 0.006468f
C413 B.n373 VSUBS 0.006468f
C414 B.n374 VSUBS 0.006468f
C415 B.n375 VSUBS 0.006468f
C416 B.n376 VSUBS 0.006468f
C417 B.n377 VSUBS 0.006468f
C418 B.n378 VSUBS 0.006468f
C419 B.n379 VSUBS 0.006468f
C420 B.n380 VSUBS 0.006468f
C421 B.n381 VSUBS 0.006468f
C422 B.n382 VSUBS 0.006468f
C423 B.n383 VSUBS 0.006468f
C424 B.n384 VSUBS 0.006468f
C425 B.n385 VSUBS 0.006468f
C426 B.n386 VSUBS 0.006468f
C427 B.n387 VSUBS 0.006468f
C428 B.n388 VSUBS 0.006468f
C429 B.n389 VSUBS 0.006468f
C430 B.n390 VSUBS 0.006468f
C431 B.n391 VSUBS 0.006468f
C432 B.n392 VSUBS 0.006468f
C433 B.n393 VSUBS 0.006468f
C434 B.n394 VSUBS 0.006468f
C435 B.n395 VSUBS 0.006468f
C436 B.n396 VSUBS 0.006468f
C437 B.n397 VSUBS 0.006468f
C438 B.n398 VSUBS 0.006468f
C439 B.n399 VSUBS 0.015208f
C440 B.n400 VSUBS 0.015208f
C441 B.n401 VSUBS 0.01485f
C442 B.n402 VSUBS 0.006468f
C443 B.n403 VSUBS 0.006468f
C444 B.n404 VSUBS 0.006468f
C445 B.n405 VSUBS 0.006468f
C446 B.n406 VSUBS 0.006468f
C447 B.n407 VSUBS 0.006468f
C448 B.n408 VSUBS 0.006468f
C449 B.n409 VSUBS 0.006468f
C450 B.n410 VSUBS 0.006468f
C451 B.n411 VSUBS 0.006468f
C452 B.n412 VSUBS 0.006468f
C453 B.n413 VSUBS 0.006468f
C454 B.n414 VSUBS 0.006468f
C455 B.n415 VSUBS 0.006468f
C456 B.n416 VSUBS 0.006468f
C457 B.n417 VSUBS 0.006468f
C458 B.n418 VSUBS 0.006468f
C459 B.n419 VSUBS 0.006468f
C460 B.n420 VSUBS 0.006468f
C461 B.n421 VSUBS 0.006468f
C462 B.n422 VSUBS 0.006468f
C463 B.n423 VSUBS 0.006468f
C464 B.n424 VSUBS 0.006468f
C465 B.n425 VSUBS 0.006468f
C466 B.n426 VSUBS 0.006468f
C467 B.n427 VSUBS 0.006468f
C468 B.n428 VSUBS 0.006468f
C469 B.n429 VSUBS 0.006468f
C470 B.n430 VSUBS 0.006468f
C471 B.n431 VSUBS 0.006468f
C472 B.n432 VSUBS 0.006468f
C473 B.n433 VSUBS 0.006468f
C474 B.n434 VSUBS 0.006468f
C475 B.n435 VSUBS 0.006468f
C476 B.n436 VSUBS 0.006468f
C477 B.n437 VSUBS 0.006468f
C478 B.n438 VSUBS 0.006468f
C479 B.n439 VSUBS 0.006468f
C480 B.n440 VSUBS 0.006468f
C481 B.n441 VSUBS 0.006468f
C482 B.n442 VSUBS 0.006468f
C483 B.n443 VSUBS 0.006468f
C484 B.n444 VSUBS 0.006468f
C485 B.n445 VSUBS 0.006468f
C486 B.n446 VSUBS 0.006468f
C487 B.n447 VSUBS 0.006468f
C488 B.n448 VSUBS 0.006468f
C489 B.n449 VSUBS 0.006468f
C490 B.n450 VSUBS 0.006468f
C491 B.n451 VSUBS 0.006468f
C492 B.n452 VSUBS 0.006468f
C493 B.n453 VSUBS 0.006468f
C494 B.n454 VSUBS 0.006468f
C495 B.n455 VSUBS 0.006468f
C496 B.n456 VSUBS 0.006468f
C497 B.n457 VSUBS 0.006468f
C498 B.n458 VSUBS 0.006468f
C499 B.n459 VSUBS 0.006468f
C500 B.n460 VSUBS 0.006468f
C501 B.n461 VSUBS 0.006468f
C502 B.n462 VSUBS 0.006468f
C503 B.n463 VSUBS 0.006468f
C504 B.n464 VSUBS 0.006468f
C505 B.n465 VSUBS 0.006468f
C506 B.n466 VSUBS 0.006468f
C507 B.n467 VSUBS 0.006468f
C508 B.n468 VSUBS 0.006468f
C509 B.n469 VSUBS 0.006468f
C510 B.n470 VSUBS 0.006468f
C511 B.n471 VSUBS 0.006468f
C512 B.n472 VSUBS 0.006468f
C513 B.n473 VSUBS 0.006468f
C514 B.n474 VSUBS 0.006468f
C515 B.n475 VSUBS 0.006468f
C516 B.n476 VSUBS 0.006468f
C517 B.n477 VSUBS 0.006468f
C518 B.n478 VSUBS 0.006468f
C519 B.n479 VSUBS 0.006468f
C520 B.n480 VSUBS 0.006468f
C521 B.n481 VSUBS 0.006468f
C522 B.n482 VSUBS 0.006468f
C523 B.n483 VSUBS 0.006468f
C524 B.n484 VSUBS 0.006468f
C525 B.n485 VSUBS 0.006468f
C526 B.n486 VSUBS 0.006468f
C527 B.n487 VSUBS 0.006468f
C528 B.n488 VSUBS 0.006468f
C529 B.n489 VSUBS 0.006468f
C530 B.n490 VSUBS 0.006468f
C531 B.n491 VSUBS 0.006468f
C532 B.n492 VSUBS 0.006468f
C533 B.n493 VSUBS 0.006468f
C534 B.n494 VSUBS 0.006468f
C535 B.n495 VSUBS 0.006468f
C536 B.n496 VSUBS 0.006468f
C537 B.n497 VSUBS 0.01485f
C538 B.n498 VSUBS 0.015208f
C539 B.n499 VSUBS 0.014436f
C540 B.n500 VSUBS 0.006468f
C541 B.n501 VSUBS 0.006468f
C542 B.n502 VSUBS 0.006468f
C543 B.n503 VSUBS 0.006468f
C544 B.n504 VSUBS 0.006468f
C545 B.n505 VSUBS 0.006468f
C546 B.n506 VSUBS 0.006468f
C547 B.n507 VSUBS 0.006468f
C548 B.n508 VSUBS 0.006468f
C549 B.n509 VSUBS 0.006468f
C550 B.n510 VSUBS 0.006468f
C551 B.n511 VSUBS 0.006468f
C552 B.n512 VSUBS 0.006468f
C553 B.n513 VSUBS 0.006468f
C554 B.n514 VSUBS 0.006468f
C555 B.n515 VSUBS 0.006468f
C556 B.n516 VSUBS 0.006468f
C557 B.n517 VSUBS 0.006468f
C558 B.n518 VSUBS 0.006468f
C559 B.n519 VSUBS 0.006468f
C560 B.n520 VSUBS 0.006468f
C561 B.n521 VSUBS 0.006468f
C562 B.n522 VSUBS 0.006468f
C563 B.n523 VSUBS 0.006468f
C564 B.n524 VSUBS 0.006468f
C565 B.n525 VSUBS 0.006468f
C566 B.n526 VSUBS 0.006468f
C567 B.n527 VSUBS 0.006468f
C568 B.n528 VSUBS 0.006468f
C569 B.n529 VSUBS 0.006468f
C570 B.n530 VSUBS 0.006468f
C571 B.n531 VSUBS 0.006468f
C572 B.n532 VSUBS 0.006468f
C573 B.n533 VSUBS 0.006468f
C574 B.n534 VSUBS 0.006468f
C575 B.n535 VSUBS 0.006468f
C576 B.n536 VSUBS 0.006468f
C577 B.n537 VSUBS 0.006468f
C578 B.n538 VSUBS 0.006468f
C579 B.n539 VSUBS 0.006468f
C580 B.n540 VSUBS 0.006468f
C581 B.n541 VSUBS 0.006468f
C582 B.n542 VSUBS 0.006468f
C583 B.n543 VSUBS 0.006468f
C584 B.n544 VSUBS 0.006468f
C585 B.n545 VSUBS 0.006468f
C586 B.n546 VSUBS 0.006468f
C587 B.n547 VSUBS 0.006468f
C588 B.n548 VSUBS 0.006468f
C589 B.n549 VSUBS 0.006468f
C590 B.n550 VSUBS 0.006468f
C591 B.n551 VSUBS 0.006468f
C592 B.n552 VSUBS 0.006468f
C593 B.n553 VSUBS 0.006468f
C594 B.n554 VSUBS 0.006468f
C595 B.n555 VSUBS 0.006468f
C596 B.n556 VSUBS 0.006468f
C597 B.n557 VSUBS 0.006468f
C598 B.n558 VSUBS 0.006468f
C599 B.n559 VSUBS 0.006468f
C600 B.n560 VSUBS 0.006468f
C601 B.n561 VSUBS 0.006468f
C602 B.n562 VSUBS 0.006468f
C603 B.n563 VSUBS 0.006468f
C604 B.n564 VSUBS 0.006468f
C605 B.n565 VSUBS 0.006468f
C606 B.n566 VSUBS 0.006468f
C607 B.n567 VSUBS 0.006468f
C608 B.n568 VSUBS 0.006468f
C609 B.n569 VSUBS 0.006468f
C610 B.n570 VSUBS 0.006468f
C611 B.n571 VSUBS 0.006468f
C612 B.n572 VSUBS 0.006468f
C613 B.n573 VSUBS 0.004471f
C614 B.n574 VSUBS 0.006468f
C615 B.n575 VSUBS 0.006468f
C616 B.n576 VSUBS 0.005232f
C617 B.n577 VSUBS 0.006468f
C618 B.n578 VSUBS 0.006468f
C619 B.n579 VSUBS 0.006468f
C620 B.n580 VSUBS 0.006468f
C621 B.n581 VSUBS 0.006468f
C622 B.n582 VSUBS 0.006468f
C623 B.n583 VSUBS 0.006468f
C624 B.n584 VSUBS 0.006468f
C625 B.n585 VSUBS 0.006468f
C626 B.n586 VSUBS 0.006468f
C627 B.n587 VSUBS 0.006468f
C628 B.n588 VSUBS 0.005232f
C629 B.n589 VSUBS 0.014986f
C630 B.n590 VSUBS 0.004471f
C631 B.n591 VSUBS 0.006468f
C632 B.n592 VSUBS 0.006468f
C633 B.n593 VSUBS 0.006468f
C634 B.n594 VSUBS 0.006468f
C635 B.n595 VSUBS 0.006468f
C636 B.n596 VSUBS 0.006468f
C637 B.n597 VSUBS 0.006468f
C638 B.n598 VSUBS 0.006468f
C639 B.n599 VSUBS 0.006468f
C640 B.n600 VSUBS 0.006468f
C641 B.n601 VSUBS 0.006468f
C642 B.n602 VSUBS 0.006468f
C643 B.n603 VSUBS 0.006468f
C644 B.n604 VSUBS 0.006468f
C645 B.n605 VSUBS 0.006468f
C646 B.n606 VSUBS 0.006468f
C647 B.n607 VSUBS 0.006468f
C648 B.n608 VSUBS 0.006468f
C649 B.n609 VSUBS 0.006468f
C650 B.n610 VSUBS 0.006468f
C651 B.n611 VSUBS 0.006468f
C652 B.n612 VSUBS 0.006468f
C653 B.n613 VSUBS 0.006468f
C654 B.n614 VSUBS 0.006468f
C655 B.n615 VSUBS 0.006468f
C656 B.n616 VSUBS 0.006468f
C657 B.n617 VSUBS 0.006468f
C658 B.n618 VSUBS 0.006468f
C659 B.n619 VSUBS 0.006468f
C660 B.n620 VSUBS 0.006468f
C661 B.n621 VSUBS 0.006468f
C662 B.n622 VSUBS 0.006468f
C663 B.n623 VSUBS 0.006468f
C664 B.n624 VSUBS 0.006468f
C665 B.n625 VSUBS 0.006468f
C666 B.n626 VSUBS 0.006468f
C667 B.n627 VSUBS 0.006468f
C668 B.n628 VSUBS 0.006468f
C669 B.n629 VSUBS 0.006468f
C670 B.n630 VSUBS 0.006468f
C671 B.n631 VSUBS 0.006468f
C672 B.n632 VSUBS 0.006468f
C673 B.n633 VSUBS 0.006468f
C674 B.n634 VSUBS 0.006468f
C675 B.n635 VSUBS 0.006468f
C676 B.n636 VSUBS 0.006468f
C677 B.n637 VSUBS 0.006468f
C678 B.n638 VSUBS 0.006468f
C679 B.n639 VSUBS 0.006468f
C680 B.n640 VSUBS 0.006468f
C681 B.n641 VSUBS 0.006468f
C682 B.n642 VSUBS 0.006468f
C683 B.n643 VSUBS 0.006468f
C684 B.n644 VSUBS 0.006468f
C685 B.n645 VSUBS 0.006468f
C686 B.n646 VSUBS 0.006468f
C687 B.n647 VSUBS 0.006468f
C688 B.n648 VSUBS 0.006468f
C689 B.n649 VSUBS 0.006468f
C690 B.n650 VSUBS 0.006468f
C691 B.n651 VSUBS 0.006468f
C692 B.n652 VSUBS 0.006468f
C693 B.n653 VSUBS 0.006468f
C694 B.n654 VSUBS 0.006468f
C695 B.n655 VSUBS 0.006468f
C696 B.n656 VSUBS 0.006468f
C697 B.n657 VSUBS 0.006468f
C698 B.n658 VSUBS 0.006468f
C699 B.n659 VSUBS 0.006468f
C700 B.n660 VSUBS 0.006468f
C701 B.n661 VSUBS 0.006468f
C702 B.n662 VSUBS 0.006468f
C703 B.n663 VSUBS 0.006468f
C704 B.n664 VSUBS 0.006468f
C705 B.n665 VSUBS 0.015208f
C706 B.n666 VSUBS 0.01485f
C707 B.n667 VSUBS 0.01485f
C708 B.n668 VSUBS 0.006468f
C709 B.n669 VSUBS 0.006468f
C710 B.n670 VSUBS 0.006468f
C711 B.n671 VSUBS 0.006468f
C712 B.n672 VSUBS 0.006468f
C713 B.n673 VSUBS 0.006468f
C714 B.n674 VSUBS 0.006468f
C715 B.n675 VSUBS 0.006468f
C716 B.n676 VSUBS 0.006468f
C717 B.n677 VSUBS 0.006468f
C718 B.n678 VSUBS 0.006468f
C719 B.n679 VSUBS 0.006468f
C720 B.n680 VSUBS 0.006468f
C721 B.n681 VSUBS 0.006468f
C722 B.n682 VSUBS 0.006468f
C723 B.n683 VSUBS 0.006468f
C724 B.n684 VSUBS 0.006468f
C725 B.n685 VSUBS 0.006468f
C726 B.n686 VSUBS 0.006468f
C727 B.n687 VSUBS 0.006468f
C728 B.n688 VSUBS 0.006468f
C729 B.n689 VSUBS 0.006468f
C730 B.n690 VSUBS 0.006468f
C731 B.n691 VSUBS 0.006468f
C732 B.n692 VSUBS 0.006468f
C733 B.n693 VSUBS 0.006468f
C734 B.n694 VSUBS 0.006468f
C735 B.n695 VSUBS 0.006468f
C736 B.n696 VSUBS 0.006468f
C737 B.n697 VSUBS 0.006468f
C738 B.n698 VSUBS 0.006468f
C739 B.n699 VSUBS 0.006468f
C740 B.n700 VSUBS 0.006468f
C741 B.n701 VSUBS 0.006468f
C742 B.n702 VSUBS 0.006468f
C743 B.n703 VSUBS 0.006468f
C744 B.n704 VSUBS 0.006468f
C745 B.n705 VSUBS 0.006468f
C746 B.n706 VSUBS 0.006468f
C747 B.n707 VSUBS 0.006468f
C748 B.n708 VSUBS 0.006468f
C749 B.n709 VSUBS 0.006468f
C750 B.n710 VSUBS 0.006468f
C751 B.n711 VSUBS 0.006468f
C752 B.n712 VSUBS 0.006468f
C753 B.n713 VSUBS 0.006468f
C754 B.n714 VSUBS 0.006468f
C755 B.n715 VSUBS 0.014646f
C756 VDD2.t0 VSUBS 0.317803f
C757 VDD2.t3 VSUBS 0.317803f
C758 VDD2.n0 VSUBS 3.38892f
C759 VDD2.t1 VSUBS 0.317803f
C760 VDD2.t2 VSUBS 0.317803f
C761 VDD2.n1 VSUBS 2.59263f
C762 VDD2.n2 VSUBS 4.54303f
C763 VN.t3 VSUBS 3.45633f
C764 VN.t0 VSUBS 3.45185f
C765 VN.n0 VSUBS 2.24432f
C766 VN.t1 VSUBS 3.45633f
C767 VN.t2 VSUBS 3.45185f
C768 VN.n1 VSUBS 4.03015f
C769 VDD1.t0 VSUBS 0.320479f
C770 VDD1.t3 VSUBS 0.320479f
C771 VDD1.n0 VSUBS 2.61503f
C772 VDD1.t1 VSUBS 0.320479f
C773 VDD1.t2 VSUBS 0.320479f
C774 VDD1.n1 VSUBS 3.44347f
C775 VTAIL.t1 VSUBS 2.74303f
C776 VTAIL.n0 VSUBS 0.73839f
C777 VTAIL.t5 VSUBS 2.74303f
C778 VTAIL.n1 VSUBS 0.819088f
C779 VTAIL.t4 VSUBS 2.74303f
C780 VTAIL.n2 VSUBS 2.21986f
C781 VTAIL.t2 VSUBS 2.74303f
C782 VTAIL.n3 VSUBS 2.21986f
C783 VTAIL.t0 VSUBS 2.74303f
C784 VTAIL.n4 VSUBS 0.819083f
C785 VTAIL.t3 VSUBS 2.74303f
C786 VTAIL.n5 VSUBS 0.819083f
C787 VTAIL.t6 VSUBS 2.74303f
C788 VTAIL.n6 VSUBS 2.21986f
C789 VTAIL.t7 VSUBS 2.74303f
C790 VTAIL.n7 VSUBS 2.13063f
C791 VP.n0 VSUBS 0.044367f
C792 VP.t1 VSUBS 3.29569f
C793 VP.n1 VSUBS 0.027181f
C794 VP.n2 VSUBS 0.044367f
C795 VP.t2 VSUBS 3.29569f
C796 VP.t0 VSUBS 3.55204f
C797 VP.t3 VSUBS 3.55666f
C798 VP.n3 VSUBS 4.12968f
C799 VP.n4 VSUBS 1.98633f
C800 VP.n5 VSUBS 1.26869f
C801 VP.n6 VSUBS 0.052857f
C802 VP.n7 VSUBS 0.066535f
C803 VP.n8 VSUBS 0.033654f
C804 VP.n9 VSUBS 0.033654f
C805 VP.n10 VSUBS 0.033654f
C806 VP.n11 VSUBS 0.066535f
C807 VP.n12 VSUBS 0.052857f
C808 VP.n13 VSUBS 1.26869f
C809 VP.n14 VSUBS 0.046037f
.ends

