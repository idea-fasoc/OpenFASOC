* NGSPICE file created from diff_pair_sample_0126.ext - technology: sky130A

.subckt diff_pair_sample_0126 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 w_n1318_n2868# sky130_fd_pr__pfet_01v8 ad=3.6972 pd=19.74 as=3.6972 ps=19.74 w=9.48 l=0.54
X1 B.t11 B.t9 B.t10 w_n1318_n2868# sky130_fd_pr__pfet_01v8 ad=3.6972 pd=19.74 as=0 ps=0 w=9.48 l=0.54
X2 VDD1.t1 VP.t0 VTAIL.t1 w_n1318_n2868# sky130_fd_pr__pfet_01v8 ad=3.6972 pd=19.74 as=3.6972 ps=19.74 w=9.48 l=0.54
X3 B.t8 B.t6 B.t7 w_n1318_n2868# sky130_fd_pr__pfet_01v8 ad=3.6972 pd=19.74 as=0 ps=0 w=9.48 l=0.54
X4 B.t5 B.t3 B.t4 w_n1318_n2868# sky130_fd_pr__pfet_01v8 ad=3.6972 pd=19.74 as=0 ps=0 w=9.48 l=0.54
X5 B.t2 B.t0 B.t1 w_n1318_n2868# sky130_fd_pr__pfet_01v8 ad=3.6972 pd=19.74 as=0 ps=0 w=9.48 l=0.54
X6 VDD1.t0 VP.t1 VTAIL.t0 w_n1318_n2868# sky130_fd_pr__pfet_01v8 ad=3.6972 pd=19.74 as=3.6972 ps=19.74 w=9.48 l=0.54
X7 VDD2.t0 VN.t1 VTAIL.t3 w_n1318_n2868# sky130_fd_pr__pfet_01v8 ad=3.6972 pd=19.74 as=3.6972 ps=19.74 w=9.48 l=0.54
R0 VN VN.t1 695.708
R1 VN VN.t0 658.08
R2 VTAIL.n202 VTAIL.n156 756.745
R3 VTAIL.n46 VTAIL.n0 756.745
R4 VTAIL.n150 VTAIL.n104 756.745
R5 VTAIL.n98 VTAIL.n52 756.745
R6 VTAIL.n172 VTAIL.n171 585
R7 VTAIL.n177 VTAIL.n176 585
R8 VTAIL.n179 VTAIL.n178 585
R9 VTAIL.n168 VTAIL.n167 585
R10 VTAIL.n185 VTAIL.n184 585
R11 VTAIL.n187 VTAIL.n186 585
R12 VTAIL.n164 VTAIL.n163 585
R13 VTAIL.n193 VTAIL.n192 585
R14 VTAIL.n195 VTAIL.n194 585
R15 VTAIL.n160 VTAIL.n159 585
R16 VTAIL.n201 VTAIL.n200 585
R17 VTAIL.n203 VTAIL.n202 585
R18 VTAIL.n16 VTAIL.n15 585
R19 VTAIL.n21 VTAIL.n20 585
R20 VTAIL.n23 VTAIL.n22 585
R21 VTAIL.n12 VTAIL.n11 585
R22 VTAIL.n29 VTAIL.n28 585
R23 VTAIL.n31 VTAIL.n30 585
R24 VTAIL.n8 VTAIL.n7 585
R25 VTAIL.n37 VTAIL.n36 585
R26 VTAIL.n39 VTAIL.n38 585
R27 VTAIL.n4 VTAIL.n3 585
R28 VTAIL.n45 VTAIL.n44 585
R29 VTAIL.n47 VTAIL.n46 585
R30 VTAIL.n151 VTAIL.n150 585
R31 VTAIL.n149 VTAIL.n148 585
R32 VTAIL.n108 VTAIL.n107 585
R33 VTAIL.n143 VTAIL.n142 585
R34 VTAIL.n141 VTAIL.n140 585
R35 VTAIL.n112 VTAIL.n111 585
R36 VTAIL.n135 VTAIL.n134 585
R37 VTAIL.n133 VTAIL.n132 585
R38 VTAIL.n116 VTAIL.n115 585
R39 VTAIL.n127 VTAIL.n126 585
R40 VTAIL.n125 VTAIL.n124 585
R41 VTAIL.n120 VTAIL.n119 585
R42 VTAIL.n99 VTAIL.n98 585
R43 VTAIL.n97 VTAIL.n96 585
R44 VTAIL.n56 VTAIL.n55 585
R45 VTAIL.n91 VTAIL.n90 585
R46 VTAIL.n89 VTAIL.n88 585
R47 VTAIL.n60 VTAIL.n59 585
R48 VTAIL.n83 VTAIL.n82 585
R49 VTAIL.n81 VTAIL.n80 585
R50 VTAIL.n64 VTAIL.n63 585
R51 VTAIL.n75 VTAIL.n74 585
R52 VTAIL.n73 VTAIL.n72 585
R53 VTAIL.n68 VTAIL.n67 585
R54 VTAIL.n173 VTAIL.t2 327.467
R55 VTAIL.n17 VTAIL.t1 327.467
R56 VTAIL.n69 VTAIL.t3 327.467
R57 VTAIL.n121 VTAIL.t0 327.467
R58 VTAIL.n177 VTAIL.n171 171.744
R59 VTAIL.n178 VTAIL.n177 171.744
R60 VTAIL.n178 VTAIL.n167 171.744
R61 VTAIL.n185 VTAIL.n167 171.744
R62 VTAIL.n186 VTAIL.n185 171.744
R63 VTAIL.n186 VTAIL.n163 171.744
R64 VTAIL.n193 VTAIL.n163 171.744
R65 VTAIL.n194 VTAIL.n193 171.744
R66 VTAIL.n194 VTAIL.n159 171.744
R67 VTAIL.n201 VTAIL.n159 171.744
R68 VTAIL.n202 VTAIL.n201 171.744
R69 VTAIL.n21 VTAIL.n15 171.744
R70 VTAIL.n22 VTAIL.n21 171.744
R71 VTAIL.n22 VTAIL.n11 171.744
R72 VTAIL.n29 VTAIL.n11 171.744
R73 VTAIL.n30 VTAIL.n29 171.744
R74 VTAIL.n30 VTAIL.n7 171.744
R75 VTAIL.n37 VTAIL.n7 171.744
R76 VTAIL.n38 VTAIL.n37 171.744
R77 VTAIL.n38 VTAIL.n3 171.744
R78 VTAIL.n45 VTAIL.n3 171.744
R79 VTAIL.n46 VTAIL.n45 171.744
R80 VTAIL.n150 VTAIL.n149 171.744
R81 VTAIL.n149 VTAIL.n107 171.744
R82 VTAIL.n142 VTAIL.n107 171.744
R83 VTAIL.n142 VTAIL.n141 171.744
R84 VTAIL.n141 VTAIL.n111 171.744
R85 VTAIL.n134 VTAIL.n111 171.744
R86 VTAIL.n134 VTAIL.n133 171.744
R87 VTAIL.n133 VTAIL.n115 171.744
R88 VTAIL.n126 VTAIL.n115 171.744
R89 VTAIL.n126 VTAIL.n125 171.744
R90 VTAIL.n125 VTAIL.n119 171.744
R91 VTAIL.n98 VTAIL.n97 171.744
R92 VTAIL.n97 VTAIL.n55 171.744
R93 VTAIL.n90 VTAIL.n55 171.744
R94 VTAIL.n90 VTAIL.n89 171.744
R95 VTAIL.n89 VTAIL.n59 171.744
R96 VTAIL.n82 VTAIL.n59 171.744
R97 VTAIL.n82 VTAIL.n81 171.744
R98 VTAIL.n81 VTAIL.n63 171.744
R99 VTAIL.n74 VTAIL.n63 171.744
R100 VTAIL.n74 VTAIL.n73 171.744
R101 VTAIL.n73 VTAIL.n67 171.744
R102 VTAIL.t2 VTAIL.n171 85.8723
R103 VTAIL.t1 VTAIL.n15 85.8723
R104 VTAIL.t0 VTAIL.n119 85.8723
R105 VTAIL.t3 VTAIL.n67 85.8723
R106 VTAIL.n207 VTAIL.n206 29.8581
R107 VTAIL.n51 VTAIL.n50 29.8581
R108 VTAIL.n155 VTAIL.n154 29.8581
R109 VTAIL.n103 VTAIL.n102 29.8581
R110 VTAIL.n103 VTAIL.n51 22.0565
R111 VTAIL.n207 VTAIL.n155 21.3065
R112 VTAIL.n173 VTAIL.n172 16.3895
R113 VTAIL.n17 VTAIL.n16 16.3895
R114 VTAIL.n121 VTAIL.n120 16.3895
R115 VTAIL.n69 VTAIL.n68 16.3895
R116 VTAIL.n176 VTAIL.n175 12.8005
R117 VTAIL.n20 VTAIL.n19 12.8005
R118 VTAIL.n124 VTAIL.n123 12.8005
R119 VTAIL.n72 VTAIL.n71 12.8005
R120 VTAIL.n179 VTAIL.n170 12.0247
R121 VTAIL.n23 VTAIL.n14 12.0247
R122 VTAIL.n127 VTAIL.n118 12.0247
R123 VTAIL.n75 VTAIL.n66 12.0247
R124 VTAIL.n180 VTAIL.n168 11.249
R125 VTAIL.n24 VTAIL.n12 11.249
R126 VTAIL.n128 VTAIL.n116 11.249
R127 VTAIL.n76 VTAIL.n64 11.249
R128 VTAIL.n184 VTAIL.n183 10.4732
R129 VTAIL.n28 VTAIL.n27 10.4732
R130 VTAIL.n132 VTAIL.n131 10.4732
R131 VTAIL.n80 VTAIL.n79 10.4732
R132 VTAIL.n187 VTAIL.n166 9.69747
R133 VTAIL.n206 VTAIL.n156 9.69747
R134 VTAIL.n31 VTAIL.n10 9.69747
R135 VTAIL.n50 VTAIL.n0 9.69747
R136 VTAIL.n154 VTAIL.n104 9.69747
R137 VTAIL.n135 VTAIL.n114 9.69747
R138 VTAIL.n102 VTAIL.n52 9.69747
R139 VTAIL.n83 VTAIL.n62 9.69747
R140 VTAIL.n206 VTAIL.n205 9.45567
R141 VTAIL.n50 VTAIL.n49 9.45567
R142 VTAIL.n154 VTAIL.n153 9.45567
R143 VTAIL.n102 VTAIL.n101 9.45567
R144 VTAIL.n197 VTAIL.n196 9.3005
R145 VTAIL.n199 VTAIL.n198 9.3005
R146 VTAIL.n158 VTAIL.n157 9.3005
R147 VTAIL.n205 VTAIL.n204 9.3005
R148 VTAIL.n191 VTAIL.n190 9.3005
R149 VTAIL.n189 VTAIL.n188 9.3005
R150 VTAIL.n166 VTAIL.n165 9.3005
R151 VTAIL.n183 VTAIL.n182 9.3005
R152 VTAIL.n181 VTAIL.n180 9.3005
R153 VTAIL.n170 VTAIL.n169 9.3005
R154 VTAIL.n175 VTAIL.n174 9.3005
R155 VTAIL.n162 VTAIL.n161 9.3005
R156 VTAIL.n41 VTAIL.n40 9.3005
R157 VTAIL.n43 VTAIL.n42 9.3005
R158 VTAIL.n2 VTAIL.n1 9.3005
R159 VTAIL.n49 VTAIL.n48 9.3005
R160 VTAIL.n35 VTAIL.n34 9.3005
R161 VTAIL.n33 VTAIL.n32 9.3005
R162 VTAIL.n10 VTAIL.n9 9.3005
R163 VTAIL.n27 VTAIL.n26 9.3005
R164 VTAIL.n25 VTAIL.n24 9.3005
R165 VTAIL.n14 VTAIL.n13 9.3005
R166 VTAIL.n19 VTAIL.n18 9.3005
R167 VTAIL.n6 VTAIL.n5 9.3005
R168 VTAIL.n106 VTAIL.n105 9.3005
R169 VTAIL.n147 VTAIL.n146 9.3005
R170 VTAIL.n145 VTAIL.n144 9.3005
R171 VTAIL.n110 VTAIL.n109 9.3005
R172 VTAIL.n139 VTAIL.n138 9.3005
R173 VTAIL.n137 VTAIL.n136 9.3005
R174 VTAIL.n114 VTAIL.n113 9.3005
R175 VTAIL.n131 VTAIL.n130 9.3005
R176 VTAIL.n129 VTAIL.n128 9.3005
R177 VTAIL.n118 VTAIL.n117 9.3005
R178 VTAIL.n123 VTAIL.n122 9.3005
R179 VTAIL.n153 VTAIL.n152 9.3005
R180 VTAIL.n95 VTAIL.n94 9.3005
R181 VTAIL.n54 VTAIL.n53 9.3005
R182 VTAIL.n101 VTAIL.n100 9.3005
R183 VTAIL.n93 VTAIL.n92 9.3005
R184 VTAIL.n58 VTAIL.n57 9.3005
R185 VTAIL.n87 VTAIL.n86 9.3005
R186 VTAIL.n85 VTAIL.n84 9.3005
R187 VTAIL.n62 VTAIL.n61 9.3005
R188 VTAIL.n79 VTAIL.n78 9.3005
R189 VTAIL.n77 VTAIL.n76 9.3005
R190 VTAIL.n66 VTAIL.n65 9.3005
R191 VTAIL.n71 VTAIL.n70 9.3005
R192 VTAIL.n188 VTAIL.n164 8.92171
R193 VTAIL.n204 VTAIL.n203 8.92171
R194 VTAIL.n32 VTAIL.n8 8.92171
R195 VTAIL.n48 VTAIL.n47 8.92171
R196 VTAIL.n152 VTAIL.n151 8.92171
R197 VTAIL.n136 VTAIL.n112 8.92171
R198 VTAIL.n100 VTAIL.n99 8.92171
R199 VTAIL.n84 VTAIL.n60 8.92171
R200 VTAIL.n192 VTAIL.n191 8.14595
R201 VTAIL.n200 VTAIL.n158 8.14595
R202 VTAIL.n36 VTAIL.n35 8.14595
R203 VTAIL.n44 VTAIL.n2 8.14595
R204 VTAIL.n148 VTAIL.n106 8.14595
R205 VTAIL.n140 VTAIL.n139 8.14595
R206 VTAIL.n96 VTAIL.n54 8.14595
R207 VTAIL.n88 VTAIL.n87 8.14595
R208 VTAIL.n195 VTAIL.n162 7.3702
R209 VTAIL.n199 VTAIL.n160 7.3702
R210 VTAIL.n39 VTAIL.n6 7.3702
R211 VTAIL.n43 VTAIL.n4 7.3702
R212 VTAIL.n147 VTAIL.n108 7.3702
R213 VTAIL.n143 VTAIL.n110 7.3702
R214 VTAIL.n95 VTAIL.n56 7.3702
R215 VTAIL.n91 VTAIL.n58 7.3702
R216 VTAIL.n196 VTAIL.n195 6.59444
R217 VTAIL.n196 VTAIL.n160 6.59444
R218 VTAIL.n40 VTAIL.n39 6.59444
R219 VTAIL.n40 VTAIL.n4 6.59444
R220 VTAIL.n144 VTAIL.n108 6.59444
R221 VTAIL.n144 VTAIL.n143 6.59444
R222 VTAIL.n92 VTAIL.n56 6.59444
R223 VTAIL.n92 VTAIL.n91 6.59444
R224 VTAIL.n192 VTAIL.n162 5.81868
R225 VTAIL.n200 VTAIL.n199 5.81868
R226 VTAIL.n36 VTAIL.n6 5.81868
R227 VTAIL.n44 VTAIL.n43 5.81868
R228 VTAIL.n148 VTAIL.n147 5.81868
R229 VTAIL.n140 VTAIL.n110 5.81868
R230 VTAIL.n96 VTAIL.n95 5.81868
R231 VTAIL.n88 VTAIL.n58 5.81868
R232 VTAIL.n191 VTAIL.n164 5.04292
R233 VTAIL.n203 VTAIL.n158 5.04292
R234 VTAIL.n35 VTAIL.n8 5.04292
R235 VTAIL.n47 VTAIL.n2 5.04292
R236 VTAIL.n151 VTAIL.n106 5.04292
R237 VTAIL.n139 VTAIL.n112 5.04292
R238 VTAIL.n99 VTAIL.n54 5.04292
R239 VTAIL.n87 VTAIL.n60 5.04292
R240 VTAIL.n188 VTAIL.n187 4.26717
R241 VTAIL.n204 VTAIL.n156 4.26717
R242 VTAIL.n32 VTAIL.n31 4.26717
R243 VTAIL.n48 VTAIL.n0 4.26717
R244 VTAIL.n152 VTAIL.n104 4.26717
R245 VTAIL.n136 VTAIL.n135 4.26717
R246 VTAIL.n100 VTAIL.n52 4.26717
R247 VTAIL.n84 VTAIL.n83 4.26717
R248 VTAIL.n174 VTAIL.n173 3.70984
R249 VTAIL.n18 VTAIL.n17 3.70984
R250 VTAIL.n70 VTAIL.n69 3.70984
R251 VTAIL.n122 VTAIL.n121 3.70984
R252 VTAIL.n184 VTAIL.n166 3.49141
R253 VTAIL.n28 VTAIL.n10 3.49141
R254 VTAIL.n132 VTAIL.n114 3.49141
R255 VTAIL.n80 VTAIL.n62 3.49141
R256 VTAIL.n183 VTAIL.n168 2.71565
R257 VTAIL.n27 VTAIL.n12 2.71565
R258 VTAIL.n131 VTAIL.n116 2.71565
R259 VTAIL.n79 VTAIL.n64 2.71565
R260 VTAIL.n180 VTAIL.n179 1.93989
R261 VTAIL.n24 VTAIL.n23 1.93989
R262 VTAIL.n128 VTAIL.n127 1.93989
R263 VTAIL.n76 VTAIL.n75 1.93989
R264 VTAIL.n176 VTAIL.n170 1.16414
R265 VTAIL.n20 VTAIL.n14 1.16414
R266 VTAIL.n124 VTAIL.n118 1.16414
R267 VTAIL.n72 VTAIL.n66 1.16414
R268 VTAIL.n155 VTAIL.n103 0.845328
R269 VTAIL VTAIL.n51 0.716017
R270 VTAIL.n175 VTAIL.n172 0.388379
R271 VTAIL.n19 VTAIL.n16 0.388379
R272 VTAIL.n123 VTAIL.n120 0.388379
R273 VTAIL.n71 VTAIL.n68 0.388379
R274 VTAIL.n174 VTAIL.n169 0.155672
R275 VTAIL.n181 VTAIL.n169 0.155672
R276 VTAIL.n182 VTAIL.n181 0.155672
R277 VTAIL.n182 VTAIL.n165 0.155672
R278 VTAIL.n189 VTAIL.n165 0.155672
R279 VTAIL.n190 VTAIL.n189 0.155672
R280 VTAIL.n190 VTAIL.n161 0.155672
R281 VTAIL.n197 VTAIL.n161 0.155672
R282 VTAIL.n198 VTAIL.n197 0.155672
R283 VTAIL.n198 VTAIL.n157 0.155672
R284 VTAIL.n205 VTAIL.n157 0.155672
R285 VTAIL.n18 VTAIL.n13 0.155672
R286 VTAIL.n25 VTAIL.n13 0.155672
R287 VTAIL.n26 VTAIL.n25 0.155672
R288 VTAIL.n26 VTAIL.n9 0.155672
R289 VTAIL.n33 VTAIL.n9 0.155672
R290 VTAIL.n34 VTAIL.n33 0.155672
R291 VTAIL.n34 VTAIL.n5 0.155672
R292 VTAIL.n41 VTAIL.n5 0.155672
R293 VTAIL.n42 VTAIL.n41 0.155672
R294 VTAIL.n42 VTAIL.n1 0.155672
R295 VTAIL.n49 VTAIL.n1 0.155672
R296 VTAIL.n153 VTAIL.n105 0.155672
R297 VTAIL.n146 VTAIL.n105 0.155672
R298 VTAIL.n146 VTAIL.n145 0.155672
R299 VTAIL.n145 VTAIL.n109 0.155672
R300 VTAIL.n138 VTAIL.n109 0.155672
R301 VTAIL.n138 VTAIL.n137 0.155672
R302 VTAIL.n137 VTAIL.n113 0.155672
R303 VTAIL.n130 VTAIL.n113 0.155672
R304 VTAIL.n130 VTAIL.n129 0.155672
R305 VTAIL.n129 VTAIL.n117 0.155672
R306 VTAIL.n122 VTAIL.n117 0.155672
R307 VTAIL.n101 VTAIL.n53 0.155672
R308 VTAIL.n94 VTAIL.n53 0.155672
R309 VTAIL.n94 VTAIL.n93 0.155672
R310 VTAIL.n93 VTAIL.n57 0.155672
R311 VTAIL.n86 VTAIL.n57 0.155672
R312 VTAIL.n86 VTAIL.n85 0.155672
R313 VTAIL.n85 VTAIL.n61 0.155672
R314 VTAIL.n78 VTAIL.n61 0.155672
R315 VTAIL.n78 VTAIL.n77 0.155672
R316 VTAIL.n77 VTAIL.n65 0.155672
R317 VTAIL.n70 VTAIL.n65 0.155672
R318 VTAIL VTAIL.n207 0.12981
R319 VDD2.n97 VDD2.n51 756.745
R320 VDD2.n46 VDD2.n0 756.745
R321 VDD2.n98 VDD2.n97 585
R322 VDD2.n96 VDD2.n95 585
R323 VDD2.n55 VDD2.n54 585
R324 VDD2.n90 VDD2.n89 585
R325 VDD2.n88 VDD2.n87 585
R326 VDD2.n59 VDD2.n58 585
R327 VDD2.n82 VDD2.n81 585
R328 VDD2.n80 VDD2.n79 585
R329 VDD2.n63 VDD2.n62 585
R330 VDD2.n74 VDD2.n73 585
R331 VDD2.n72 VDD2.n71 585
R332 VDD2.n67 VDD2.n66 585
R333 VDD2.n16 VDD2.n15 585
R334 VDD2.n21 VDD2.n20 585
R335 VDD2.n23 VDD2.n22 585
R336 VDD2.n12 VDD2.n11 585
R337 VDD2.n29 VDD2.n28 585
R338 VDD2.n31 VDD2.n30 585
R339 VDD2.n8 VDD2.n7 585
R340 VDD2.n37 VDD2.n36 585
R341 VDD2.n39 VDD2.n38 585
R342 VDD2.n4 VDD2.n3 585
R343 VDD2.n45 VDD2.n44 585
R344 VDD2.n47 VDD2.n46 585
R345 VDD2.n17 VDD2.t1 327.467
R346 VDD2.n68 VDD2.t0 327.467
R347 VDD2.n97 VDD2.n96 171.744
R348 VDD2.n96 VDD2.n54 171.744
R349 VDD2.n89 VDD2.n54 171.744
R350 VDD2.n89 VDD2.n88 171.744
R351 VDD2.n88 VDD2.n58 171.744
R352 VDD2.n81 VDD2.n58 171.744
R353 VDD2.n81 VDD2.n80 171.744
R354 VDD2.n80 VDD2.n62 171.744
R355 VDD2.n73 VDD2.n62 171.744
R356 VDD2.n73 VDD2.n72 171.744
R357 VDD2.n72 VDD2.n66 171.744
R358 VDD2.n21 VDD2.n15 171.744
R359 VDD2.n22 VDD2.n21 171.744
R360 VDD2.n22 VDD2.n11 171.744
R361 VDD2.n29 VDD2.n11 171.744
R362 VDD2.n30 VDD2.n29 171.744
R363 VDD2.n30 VDD2.n7 171.744
R364 VDD2.n37 VDD2.n7 171.744
R365 VDD2.n38 VDD2.n37 171.744
R366 VDD2.n38 VDD2.n3 171.744
R367 VDD2.n45 VDD2.n3 171.744
R368 VDD2.n46 VDD2.n45 171.744
R369 VDD2.t0 VDD2.n66 85.8723
R370 VDD2.t1 VDD2.n15 85.8723
R371 VDD2.n102 VDD2.n50 79.886
R372 VDD2.n102 VDD2.n101 46.5369
R373 VDD2.n68 VDD2.n67 16.3895
R374 VDD2.n17 VDD2.n16 16.3895
R375 VDD2.n71 VDD2.n70 12.8005
R376 VDD2.n20 VDD2.n19 12.8005
R377 VDD2.n74 VDD2.n65 12.0247
R378 VDD2.n23 VDD2.n14 12.0247
R379 VDD2.n75 VDD2.n63 11.249
R380 VDD2.n24 VDD2.n12 11.249
R381 VDD2.n79 VDD2.n78 10.4732
R382 VDD2.n28 VDD2.n27 10.4732
R383 VDD2.n101 VDD2.n51 9.69747
R384 VDD2.n82 VDD2.n61 9.69747
R385 VDD2.n31 VDD2.n10 9.69747
R386 VDD2.n50 VDD2.n0 9.69747
R387 VDD2.n101 VDD2.n100 9.45567
R388 VDD2.n50 VDD2.n49 9.45567
R389 VDD2.n53 VDD2.n52 9.3005
R390 VDD2.n94 VDD2.n93 9.3005
R391 VDD2.n92 VDD2.n91 9.3005
R392 VDD2.n57 VDD2.n56 9.3005
R393 VDD2.n86 VDD2.n85 9.3005
R394 VDD2.n84 VDD2.n83 9.3005
R395 VDD2.n61 VDD2.n60 9.3005
R396 VDD2.n78 VDD2.n77 9.3005
R397 VDD2.n76 VDD2.n75 9.3005
R398 VDD2.n65 VDD2.n64 9.3005
R399 VDD2.n70 VDD2.n69 9.3005
R400 VDD2.n100 VDD2.n99 9.3005
R401 VDD2.n41 VDD2.n40 9.3005
R402 VDD2.n43 VDD2.n42 9.3005
R403 VDD2.n2 VDD2.n1 9.3005
R404 VDD2.n49 VDD2.n48 9.3005
R405 VDD2.n35 VDD2.n34 9.3005
R406 VDD2.n33 VDD2.n32 9.3005
R407 VDD2.n10 VDD2.n9 9.3005
R408 VDD2.n27 VDD2.n26 9.3005
R409 VDD2.n25 VDD2.n24 9.3005
R410 VDD2.n14 VDD2.n13 9.3005
R411 VDD2.n19 VDD2.n18 9.3005
R412 VDD2.n6 VDD2.n5 9.3005
R413 VDD2.n99 VDD2.n98 8.92171
R414 VDD2.n83 VDD2.n59 8.92171
R415 VDD2.n32 VDD2.n8 8.92171
R416 VDD2.n48 VDD2.n47 8.92171
R417 VDD2.n95 VDD2.n53 8.14595
R418 VDD2.n87 VDD2.n86 8.14595
R419 VDD2.n36 VDD2.n35 8.14595
R420 VDD2.n44 VDD2.n2 8.14595
R421 VDD2.n94 VDD2.n55 7.3702
R422 VDD2.n90 VDD2.n57 7.3702
R423 VDD2.n39 VDD2.n6 7.3702
R424 VDD2.n43 VDD2.n4 7.3702
R425 VDD2.n91 VDD2.n55 6.59444
R426 VDD2.n91 VDD2.n90 6.59444
R427 VDD2.n40 VDD2.n39 6.59444
R428 VDD2.n40 VDD2.n4 6.59444
R429 VDD2.n95 VDD2.n94 5.81868
R430 VDD2.n87 VDD2.n57 5.81868
R431 VDD2.n36 VDD2.n6 5.81868
R432 VDD2.n44 VDD2.n43 5.81868
R433 VDD2.n98 VDD2.n53 5.04292
R434 VDD2.n86 VDD2.n59 5.04292
R435 VDD2.n35 VDD2.n8 5.04292
R436 VDD2.n47 VDD2.n2 5.04292
R437 VDD2.n99 VDD2.n51 4.26717
R438 VDD2.n83 VDD2.n82 4.26717
R439 VDD2.n32 VDD2.n31 4.26717
R440 VDD2.n48 VDD2.n0 4.26717
R441 VDD2.n18 VDD2.n17 3.70984
R442 VDD2.n69 VDD2.n68 3.70984
R443 VDD2.n79 VDD2.n61 3.49141
R444 VDD2.n28 VDD2.n10 3.49141
R445 VDD2.n78 VDD2.n63 2.71565
R446 VDD2.n27 VDD2.n12 2.71565
R447 VDD2.n75 VDD2.n74 1.93989
R448 VDD2.n24 VDD2.n23 1.93989
R449 VDD2.n71 VDD2.n65 1.16414
R450 VDD2.n20 VDD2.n14 1.16414
R451 VDD2.n70 VDD2.n67 0.388379
R452 VDD2.n19 VDD2.n16 0.388379
R453 VDD2 VDD2.n102 0.24619
R454 VDD2.n100 VDD2.n52 0.155672
R455 VDD2.n93 VDD2.n52 0.155672
R456 VDD2.n93 VDD2.n92 0.155672
R457 VDD2.n92 VDD2.n56 0.155672
R458 VDD2.n85 VDD2.n56 0.155672
R459 VDD2.n85 VDD2.n84 0.155672
R460 VDD2.n84 VDD2.n60 0.155672
R461 VDD2.n77 VDD2.n60 0.155672
R462 VDD2.n77 VDD2.n76 0.155672
R463 VDD2.n76 VDD2.n64 0.155672
R464 VDD2.n69 VDD2.n64 0.155672
R465 VDD2.n18 VDD2.n13 0.155672
R466 VDD2.n25 VDD2.n13 0.155672
R467 VDD2.n26 VDD2.n25 0.155672
R468 VDD2.n26 VDD2.n9 0.155672
R469 VDD2.n33 VDD2.n9 0.155672
R470 VDD2.n34 VDD2.n33 0.155672
R471 VDD2.n34 VDD2.n5 0.155672
R472 VDD2.n41 VDD2.n5 0.155672
R473 VDD2.n42 VDD2.n41 0.155672
R474 VDD2.n42 VDD2.n1 0.155672
R475 VDD2.n49 VDD2.n1 0.155672
R476 B.n83 B.t0 628.605
R477 B.n91 B.t3 628.605
R478 B.n26 B.t6 628.605
R479 B.n34 B.t9 628.605
R480 B.n293 B.n52 585
R481 B.n295 B.n294 585
R482 B.n296 B.n51 585
R483 B.n298 B.n297 585
R484 B.n299 B.n50 585
R485 B.n301 B.n300 585
R486 B.n302 B.n49 585
R487 B.n304 B.n303 585
R488 B.n305 B.n48 585
R489 B.n307 B.n306 585
R490 B.n308 B.n47 585
R491 B.n310 B.n309 585
R492 B.n311 B.n46 585
R493 B.n313 B.n312 585
R494 B.n314 B.n45 585
R495 B.n316 B.n315 585
R496 B.n317 B.n44 585
R497 B.n319 B.n318 585
R498 B.n320 B.n43 585
R499 B.n322 B.n321 585
R500 B.n323 B.n42 585
R501 B.n325 B.n324 585
R502 B.n326 B.n41 585
R503 B.n328 B.n327 585
R504 B.n329 B.n40 585
R505 B.n331 B.n330 585
R506 B.n332 B.n39 585
R507 B.n334 B.n333 585
R508 B.n335 B.n38 585
R509 B.n337 B.n336 585
R510 B.n338 B.n37 585
R511 B.n340 B.n339 585
R512 B.n341 B.n33 585
R513 B.n343 B.n342 585
R514 B.n344 B.n32 585
R515 B.n346 B.n345 585
R516 B.n347 B.n31 585
R517 B.n349 B.n348 585
R518 B.n350 B.n30 585
R519 B.n352 B.n351 585
R520 B.n353 B.n29 585
R521 B.n355 B.n354 585
R522 B.n356 B.n28 585
R523 B.n358 B.n357 585
R524 B.n360 B.n25 585
R525 B.n362 B.n361 585
R526 B.n363 B.n24 585
R527 B.n365 B.n364 585
R528 B.n366 B.n23 585
R529 B.n368 B.n367 585
R530 B.n369 B.n22 585
R531 B.n371 B.n370 585
R532 B.n372 B.n21 585
R533 B.n374 B.n373 585
R534 B.n375 B.n20 585
R535 B.n377 B.n376 585
R536 B.n378 B.n19 585
R537 B.n380 B.n379 585
R538 B.n381 B.n18 585
R539 B.n383 B.n382 585
R540 B.n384 B.n17 585
R541 B.n386 B.n385 585
R542 B.n387 B.n16 585
R543 B.n389 B.n388 585
R544 B.n390 B.n15 585
R545 B.n392 B.n391 585
R546 B.n393 B.n14 585
R547 B.n395 B.n394 585
R548 B.n396 B.n13 585
R549 B.n398 B.n397 585
R550 B.n399 B.n12 585
R551 B.n401 B.n400 585
R552 B.n402 B.n11 585
R553 B.n404 B.n403 585
R554 B.n405 B.n10 585
R555 B.n407 B.n406 585
R556 B.n408 B.n9 585
R557 B.n410 B.n409 585
R558 B.n292 B.n291 585
R559 B.n290 B.n53 585
R560 B.n289 B.n288 585
R561 B.n287 B.n54 585
R562 B.n286 B.n285 585
R563 B.n284 B.n55 585
R564 B.n283 B.n282 585
R565 B.n281 B.n56 585
R566 B.n280 B.n279 585
R567 B.n278 B.n57 585
R568 B.n277 B.n276 585
R569 B.n275 B.n58 585
R570 B.n274 B.n273 585
R571 B.n272 B.n59 585
R572 B.n271 B.n270 585
R573 B.n269 B.n60 585
R574 B.n268 B.n267 585
R575 B.n266 B.n61 585
R576 B.n265 B.n264 585
R577 B.n263 B.n62 585
R578 B.n262 B.n261 585
R579 B.n260 B.n63 585
R580 B.n259 B.n258 585
R581 B.n257 B.n64 585
R582 B.n256 B.n255 585
R583 B.n254 B.n65 585
R584 B.n253 B.n252 585
R585 B.n134 B.n109 585
R586 B.n136 B.n135 585
R587 B.n137 B.n108 585
R588 B.n139 B.n138 585
R589 B.n140 B.n107 585
R590 B.n142 B.n141 585
R591 B.n143 B.n106 585
R592 B.n145 B.n144 585
R593 B.n146 B.n105 585
R594 B.n148 B.n147 585
R595 B.n149 B.n104 585
R596 B.n151 B.n150 585
R597 B.n152 B.n103 585
R598 B.n154 B.n153 585
R599 B.n155 B.n102 585
R600 B.n157 B.n156 585
R601 B.n158 B.n101 585
R602 B.n160 B.n159 585
R603 B.n161 B.n100 585
R604 B.n163 B.n162 585
R605 B.n164 B.n99 585
R606 B.n166 B.n165 585
R607 B.n167 B.n98 585
R608 B.n169 B.n168 585
R609 B.n170 B.n97 585
R610 B.n172 B.n171 585
R611 B.n173 B.n96 585
R612 B.n175 B.n174 585
R613 B.n176 B.n95 585
R614 B.n178 B.n177 585
R615 B.n179 B.n94 585
R616 B.n181 B.n180 585
R617 B.n182 B.n93 585
R618 B.n184 B.n183 585
R619 B.n186 B.n90 585
R620 B.n188 B.n187 585
R621 B.n189 B.n89 585
R622 B.n191 B.n190 585
R623 B.n192 B.n88 585
R624 B.n194 B.n193 585
R625 B.n195 B.n87 585
R626 B.n197 B.n196 585
R627 B.n198 B.n86 585
R628 B.n200 B.n199 585
R629 B.n202 B.n201 585
R630 B.n203 B.n82 585
R631 B.n205 B.n204 585
R632 B.n206 B.n81 585
R633 B.n208 B.n207 585
R634 B.n209 B.n80 585
R635 B.n211 B.n210 585
R636 B.n212 B.n79 585
R637 B.n214 B.n213 585
R638 B.n215 B.n78 585
R639 B.n217 B.n216 585
R640 B.n218 B.n77 585
R641 B.n220 B.n219 585
R642 B.n221 B.n76 585
R643 B.n223 B.n222 585
R644 B.n224 B.n75 585
R645 B.n226 B.n225 585
R646 B.n227 B.n74 585
R647 B.n229 B.n228 585
R648 B.n230 B.n73 585
R649 B.n232 B.n231 585
R650 B.n233 B.n72 585
R651 B.n235 B.n234 585
R652 B.n236 B.n71 585
R653 B.n238 B.n237 585
R654 B.n239 B.n70 585
R655 B.n241 B.n240 585
R656 B.n242 B.n69 585
R657 B.n244 B.n243 585
R658 B.n245 B.n68 585
R659 B.n247 B.n246 585
R660 B.n248 B.n67 585
R661 B.n250 B.n249 585
R662 B.n251 B.n66 585
R663 B.n133 B.n132 585
R664 B.n131 B.n110 585
R665 B.n130 B.n129 585
R666 B.n128 B.n111 585
R667 B.n127 B.n126 585
R668 B.n125 B.n112 585
R669 B.n124 B.n123 585
R670 B.n122 B.n113 585
R671 B.n121 B.n120 585
R672 B.n119 B.n114 585
R673 B.n118 B.n117 585
R674 B.n116 B.n115 585
R675 B.n2 B.n0 585
R676 B.n429 B.n1 585
R677 B.n428 B.n427 585
R678 B.n426 B.n3 585
R679 B.n425 B.n424 585
R680 B.n423 B.n4 585
R681 B.n422 B.n421 585
R682 B.n420 B.n5 585
R683 B.n419 B.n418 585
R684 B.n417 B.n6 585
R685 B.n416 B.n415 585
R686 B.n414 B.n7 585
R687 B.n413 B.n412 585
R688 B.n411 B.n8 585
R689 B.n431 B.n430 585
R690 B.n134 B.n133 545.355
R691 B.n411 B.n410 545.355
R692 B.n253 B.n66 545.355
R693 B.n291 B.n52 545.355
R694 B.n83 B.t2 347.317
R695 B.n34 B.t10 347.317
R696 B.n91 B.t5 347.317
R697 B.n26 B.t7 347.317
R698 B.n84 B.t1 330.445
R699 B.n35 B.t11 330.445
R700 B.n92 B.t4 330.445
R701 B.n27 B.t8 330.445
R702 B.n133 B.n110 163.367
R703 B.n129 B.n110 163.367
R704 B.n129 B.n128 163.367
R705 B.n128 B.n127 163.367
R706 B.n127 B.n112 163.367
R707 B.n123 B.n112 163.367
R708 B.n123 B.n122 163.367
R709 B.n122 B.n121 163.367
R710 B.n121 B.n114 163.367
R711 B.n117 B.n114 163.367
R712 B.n117 B.n116 163.367
R713 B.n116 B.n2 163.367
R714 B.n430 B.n2 163.367
R715 B.n430 B.n429 163.367
R716 B.n429 B.n428 163.367
R717 B.n428 B.n3 163.367
R718 B.n424 B.n3 163.367
R719 B.n424 B.n423 163.367
R720 B.n423 B.n422 163.367
R721 B.n422 B.n5 163.367
R722 B.n418 B.n5 163.367
R723 B.n418 B.n417 163.367
R724 B.n417 B.n416 163.367
R725 B.n416 B.n7 163.367
R726 B.n412 B.n7 163.367
R727 B.n412 B.n411 163.367
R728 B.n135 B.n134 163.367
R729 B.n135 B.n108 163.367
R730 B.n139 B.n108 163.367
R731 B.n140 B.n139 163.367
R732 B.n141 B.n140 163.367
R733 B.n141 B.n106 163.367
R734 B.n145 B.n106 163.367
R735 B.n146 B.n145 163.367
R736 B.n147 B.n146 163.367
R737 B.n147 B.n104 163.367
R738 B.n151 B.n104 163.367
R739 B.n152 B.n151 163.367
R740 B.n153 B.n152 163.367
R741 B.n153 B.n102 163.367
R742 B.n157 B.n102 163.367
R743 B.n158 B.n157 163.367
R744 B.n159 B.n158 163.367
R745 B.n159 B.n100 163.367
R746 B.n163 B.n100 163.367
R747 B.n164 B.n163 163.367
R748 B.n165 B.n164 163.367
R749 B.n165 B.n98 163.367
R750 B.n169 B.n98 163.367
R751 B.n170 B.n169 163.367
R752 B.n171 B.n170 163.367
R753 B.n171 B.n96 163.367
R754 B.n175 B.n96 163.367
R755 B.n176 B.n175 163.367
R756 B.n177 B.n176 163.367
R757 B.n177 B.n94 163.367
R758 B.n181 B.n94 163.367
R759 B.n182 B.n181 163.367
R760 B.n183 B.n182 163.367
R761 B.n183 B.n90 163.367
R762 B.n188 B.n90 163.367
R763 B.n189 B.n188 163.367
R764 B.n190 B.n189 163.367
R765 B.n190 B.n88 163.367
R766 B.n194 B.n88 163.367
R767 B.n195 B.n194 163.367
R768 B.n196 B.n195 163.367
R769 B.n196 B.n86 163.367
R770 B.n200 B.n86 163.367
R771 B.n201 B.n200 163.367
R772 B.n201 B.n82 163.367
R773 B.n205 B.n82 163.367
R774 B.n206 B.n205 163.367
R775 B.n207 B.n206 163.367
R776 B.n207 B.n80 163.367
R777 B.n211 B.n80 163.367
R778 B.n212 B.n211 163.367
R779 B.n213 B.n212 163.367
R780 B.n213 B.n78 163.367
R781 B.n217 B.n78 163.367
R782 B.n218 B.n217 163.367
R783 B.n219 B.n218 163.367
R784 B.n219 B.n76 163.367
R785 B.n223 B.n76 163.367
R786 B.n224 B.n223 163.367
R787 B.n225 B.n224 163.367
R788 B.n225 B.n74 163.367
R789 B.n229 B.n74 163.367
R790 B.n230 B.n229 163.367
R791 B.n231 B.n230 163.367
R792 B.n231 B.n72 163.367
R793 B.n235 B.n72 163.367
R794 B.n236 B.n235 163.367
R795 B.n237 B.n236 163.367
R796 B.n237 B.n70 163.367
R797 B.n241 B.n70 163.367
R798 B.n242 B.n241 163.367
R799 B.n243 B.n242 163.367
R800 B.n243 B.n68 163.367
R801 B.n247 B.n68 163.367
R802 B.n248 B.n247 163.367
R803 B.n249 B.n248 163.367
R804 B.n249 B.n66 163.367
R805 B.n254 B.n253 163.367
R806 B.n255 B.n254 163.367
R807 B.n255 B.n64 163.367
R808 B.n259 B.n64 163.367
R809 B.n260 B.n259 163.367
R810 B.n261 B.n260 163.367
R811 B.n261 B.n62 163.367
R812 B.n265 B.n62 163.367
R813 B.n266 B.n265 163.367
R814 B.n267 B.n266 163.367
R815 B.n267 B.n60 163.367
R816 B.n271 B.n60 163.367
R817 B.n272 B.n271 163.367
R818 B.n273 B.n272 163.367
R819 B.n273 B.n58 163.367
R820 B.n277 B.n58 163.367
R821 B.n278 B.n277 163.367
R822 B.n279 B.n278 163.367
R823 B.n279 B.n56 163.367
R824 B.n283 B.n56 163.367
R825 B.n284 B.n283 163.367
R826 B.n285 B.n284 163.367
R827 B.n285 B.n54 163.367
R828 B.n289 B.n54 163.367
R829 B.n290 B.n289 163.367
R830 B.n291 B.n290 163.367
R831 B.n410 B.n9 163.367
R832 B.n406 B.n9 163.367
R833 B.n406 B.n405 163.367
R834 B.n405 B.n404 163.367
R835 B.n404 B.n11 163.367
R836 B.n400 B.n11 163.367
R837 B.n400 B.n399 163.367
R838 B.n399 B.n398 163.367
R839 B.n398 B.n13 163.367
R840 B.n394 B.n13 163.367
R841 B.n394 B.n393 163.367
R842 B.n393 B.n392 163.367
R843 B.n392 B.n15 163.367
R844 B.n388 B.n15 163.367
R845 B.n388 B.n387 163.367
R846 B.n387 B.n386 163.367
R847 B.n386 B.n17 163.367
R848 B.n382 B.n17 163.367
R849 B.n382 B.n381 163.367
R850 B.n381 B.n380 163.367
R851 B.n380 B.n19 163.367
R852 B.n376 B.n19 163.367
R853 B.n376 B.n375 163.367
R854 B.n375 B.n374 163.367
R855 B.n374 B.n21 163.367
R856 B.n370 B.n21 163.367
R857 B.n370 B.n369 163.367
R858 B.n369 B.n368 163.367
R859 B.n368 B.n23 163.367
R860 B.n364 B.n23 163.367
R861 B.n364 B.n363 163.367
R862 B.n363 B.n362 163.367
R863 B.n362 B.n25 163.367
R864 B.n357 B.n25 163.367
R865 B.n357 B.n356 163.367
R866 B.n356 B.n355 163.367
R867 B.n355 B.n29 163.367
R868 B.n351 B.n29 163.367
R869 B.n351 B.n350 163.367
R870 B.n350 B.n349 163.367
R871 B.n349 B.n31 163.367
R872 B.n345 B.n31 163.367
R873 B.n345 B.n344 163.367
R874 B.n344 B.n343 163.367
R875 B.n343 B.n33 163.367
R876 B.n339 B.n33 163.367
R877 B.n339 B.n338 163.367
R878 B.n338 B.n337 163.367
R879 B.n337 B.n38 163.367
R880 B.n333 B.n38 163.367
R881 B.n333 B.n332 163.367
R882 B.n332 B.n331 163.367
R883 B.n331 B.n40 163.367
R884 B.n327 B.n40 163.367
R885 B.n327 B.n326 163.367
R886 B.n326 B.n325 163.367
R887 B.n325 B.n42 163.367
R888 B.n321 B.n42 163.367
R889 B.n321 B.n320 163.367
R890 B.n320 B.n319 163.367
R891 B.n319 B.n44 163.367
R892 B.n315 B.n44 163.367
R893 B.n315 B.n314 163.367
R894 B.n314 B.n313 163.367
R895 B.n313 B.n46 163.367
R896 B.n309 B.n46 163.367
R897 B.n309 B.n308 163.367
R898 B.n308 B.n307 163.367
R899 B.n307 B.n48 163.367
R900 B.n303 B.n48 163.367
R901 B.n303 B.n302 163.367
R902 B.n302 B.n301 163.367
R903 B.n301 B.n50 163.367
R904 B.n297 B.n50 163.367
R905 B.n297 B.n296 163.367
R906 B.n296 B.n295 163.367
R907 B.n295 B.n52 163.367
R908 B.n85 B.n84 59.5399
R909 B.n185 B.n92 59.5399
R910 B.n359 B.n27 59.5399
R911 B.n36 B.n35 59.5399
R912 B.n293 B.n292 35.4346
R913 B.n409 B.n8 35.4346
R914 B.n252 B.n251 35.4346
R915 B.n132 B.n109 35.4346
R916 B B.n431 18.0485
R917 B.n84 B.n83 16.8732
R918 B.n92 B.n91 16.8732
R919 B.n27 B.n26 16.8732
R920 B.n35 B.n34 16.8732
R921 B.n409 B.n408 10.6151
R922 B.n408 B.n407 10.6151
R923 B.n407 B.n10 10.6151
R924 B.n403 B.n10 10.6151
R925 B.n403 B.n402 10.6151
R926 B.n402 B.n401 10.6151
R927 B.n401 B.n12 10.6151
R928 B.n397 B.n12 10.6151
R929 B.n397 B.n396 10.6151
R930 B.n396 B.n395 10.6151
R931 B.n395 B.n14 10.6151
R932 B.n391 B.n14 10.6151
R933 B.n391 B.n390 10.6151
R934 B.n390 B.n389 10.6151
R935 B.n389 B.n16 10.6151
R936 B.n385 B.n16 10.6151
R937 B.n385 B.n384 10.6151
R938 B.n384 B.n383 10.6151
R939 B.n383 B.n18 10.6151
R940 B.n379 B.n18 10.6151
R941 B.n379 B.n378 10.6151
R942 B.n378 B.n377 10.6151
R943 B.n377 B.n20 10.6151
R944 B.n373 B.n20 10.6151
R945 B.n373 B.n372 10.6151
R946 B.n372 B.n371 10.6151
R947 B.n371 B.n22 10.6151
R948 B.n367 B.n22 10.6151
R949 B.n367 B.n366 10.6151
R950 B.n366 B.n365 10.6151
R951 B.n365 B.n24 10.6151
R952 B.n361 B.n24 10.6151
R953 B.n361 B.n360 10.6151
R954 B.n358 B.n28 10.6151
R955 B.n354 B.n28 10.6151
R956 B.n354 B.n353 10.6151
R957 B.n353 B.n352 10.6151
R958 B.n352 B.n30 10.6151
R959 B.n348 B.n30 10.6151
R960 B.n348 B.n347 10.6151
R961 B.n347 B.n346 10.6151
R962 B.n346 B.n32 10.6151
R963 B.n342 B.n341 10.6151
R964 B.n341 B.n340 10.6151
R965 B.n340 B.n37 10.6151
R966 B.n336 B.n37 10.6151
R967 B.n336 B.n335 10.6151
R968 B.n335 B.n334 10.6151
R969 B.n334 B.n39 10.6151
R970 B.n330 B.n39 10.6151
R971 B.n330 B.n329 10.6151
R972 B.n329 B.n328 10.6151
R973 B.n328 B.n41 10.6151
R974 B.n324 B.n41 10.6151
R975 B.n324 B.n323 10.6151
R976 B.n323 B.n322 10.6151
R977 B.n322 B.n43 10.6151
R978 B.n318 B.n43 10.6151
R979 B.n318 B.n317 10.6151
R980 B.n317 B.n316 10.6151
R981 B.n316 B.n45 10.6151
R982 B.n312 B.n45 10.6151
R983 B.n312 B.n311 10.6151
R984 B.n311 B.n310 10.6151
R985 B.n310 B.n47 10.6151
R986 B.n306 B.n47 10.6151
R987 B.n306 B.n305 10.6151
R988 B.n305 B.n304 10.6151
R989 B.n304 B.n49 10.6151
R990 B.n300 B.n49 10.6151
R991 B.n300 B.n299 10.6151
R992 B.n299 B.n298 10.6151
R993 B.n298 B.n51 10.6151
R994 B.n294 B.n51 10.6151
R995 B.n294 B.n293 10.6151
R996 B.n252 B.n65 10.6151
R997 B.n256 B.n65 10.6151
R998 B.n257 B.n256 10.6151
R999 B.n258 B.n257 10.6151
R1000 B.n258 B.n63 10.6151
R1001 B.n262 B.n63 10.6151
R1002 B.n263 B.n262 10.6151
R1003 B.n264 B.n263 10.6151
R1004 B.n264 B.n61 10.6151
R1005 B.n268 B.n61 10.6151
R1006 B.n269 B.n268 10.6151
R1007 B.n270 B.n269 10.6151
R1008 B.n270 B.n59 10.6151
R1009 B.n274 B.n59 10.6151
R1010 B.n275 B.n274 10.6151
R1011 B.n276 B.n275 10.6151
R1012 B.n276 B.n57 10.6151
R1013 B.n280 B.n57 10.6151
R1014 B.n281 B.n280 10.6151
R1015 B.n282 B.n281 10.6151
R1016 B.n282 B.n55 10.6151
R1017 B.n286 B.n55 10.6151
R1018 B.n287 B.n286 10.6151
R1019 B.n288 B.n287 10.6151
R1020 B.n288 B.n53 10.6151
R1021 B.n292 B.n53 10.6151
R1022 B.n136 B.n109 10.6151
R1023 B.n137 B.n136 10.6151
R1024 B.n138 B.n137 10.6151
R1025 B.n138 B.n107 10.6151
R1026 B.n142 B.n107 10.6151
R1027 B.n143 B.n142 10.6151
R1028 B.n144 B.n143 10.6151
R1029 B.n144 B.n105 10.6151
R1030 B.n148 B.n105 10.6151
R1031 B.n149 B.n148 10.6151
R1032 B.n150 B.n149 10.6151
R1033 B.n150 B.n103 10.6151
R1034 B.n154 B.n103 10.6151
R1035 B.n155 B.n154 10.6151
R1036 B.n156 B.n155 10.6151
R1037 B.n156 B.n101 10.6151
R1038 B.n160 B.n101 10.6151
R1039 B.n161 B.n160 10.6151
R1040 B.n162 B.n161 10.6151
R1041 B.n162 B.n99 10.6151
R1042 B.n166 B.n99 10.6151
R1043 B.n167 B.n166 10.6151
R1044 B.n168 B.n167 10.6151
R1045 B.n168 B.n97 10.6151
R1046 B.n172 B.n97 10.6151
R1047 B.n173 B.n172 10.6151
R1048 B.n174 B.n173 10.6151
R1049 B.n174 B.n95 10.6151
R1050 B.n178 B.n95 10.6151
R1051 B.n179 B.n178 10.6151
R1052 B.n180 B.n179 10.6151
R1053 B.n180 B.n93 10.6151
R1054 B.n184 B.n93 10.6151
R1055 B.n187 B.n186 10.6151
R1056 B.n187 B.n89 10.6151
R1057 B.n191 B.n89 10.6151
R1058 B.n192 B.n191 10.6151
R1059 B.n193 B.n192 10.6151
R1060 B.n193 B.n87 10.6151
R1061 B.n197 B.n87 10.6151
R1062 B.n198 B.n197 10.6151
R1063 B.n199 B.n198 10.6151
R1064 B.n203 B.n202 10.6151
R1065 B.n204 B.n203 10.6151
R1066 B.n204 B.n81 10.6151
R1067 B.n208 B.n81 10.6151
R1068 B.n209 B.n208 10.6151
R1069 B.n210 B.n209 10.6151
R1070 B.n210 B.n79 10.6151
R1071 B.n214 B.n79 10.6151
R1072 B.n215 B.n214 10.6151
R1073 B.n216 B.n215 10.6151
R1074 B.n216 B.n77 10.6151
R1075 B.n220 B.n77 10.6151
R1076 B.n221 B.n220 10.6151
R1077 B.n222 B.n221 10.6151
R1078 B.n222 B.n75 10.6151
R1079 B.n226 B.n75 10.6151
R1080 B.n227 B.n226 10.6151
R1081 B.n228 B.n227 10.6151
R1082 B.n228 B.n73 10.6151
R1083 B.n232 B.n73 10.6151
R1084 B.n233 B.n232 10.6151
R1085 B.n234 B.n233 10.6151
R1086 B.n234 B.n71 10.6151
R1087 B.n238 B.n71 10.6151
R1088 B.n239 B.n238 10.6151
R1089 B.n240 B.n239 10.6151
R1090 B.n240 B.n69 10.6151
R1091 B.n244 B.n69 10.6151
R1092 B.n245 B.n244 10.6151
R1093 B.n246 B.n245 10.6151
R1094 B.n246 B.n67 10.6151
R1095 B.n250 B.n67 10.6151
R1096 B.n251 B.n250 10.6151
R1097 B.n132 B.n131 10.6151
R1098 B.n131 B.n130 10.6151
R1099 B.n130 B.n111 10.6151
R1100 B.n126 B.n111 10.6151
R1101 B.n126 B.n125 10.6151
R1102 B.n125 B.n124 10.6151
R1103 B.n124 B.n113 10.6151
R1104 B.n120 B.n113 10.6151
R1105 B.n120 B.n119 10.6151
R1106 B.n119 B.n118 10.6151
R1107 B.n118 B.n115 10.6151
R1108 B.n115 B.n0 10.6151
R1109 B.n427 B.n1 10.6151
R1110 B.n427 B.n426 10.6151
R1111 B.n426 B.n425 10.6151
R1112 B.n425 B.n4 10.6151
R1113 B.n421 B.n4 10.6151
R1114 B.n421 B.n420 10.6151
R1115 B.n420 B.n419 10.6151
R1116 B.n419 B.n6 10.6151
R1117 B.n415 B.n6 10.6151
R1118 B.n415 B.n414 10.6151
R1119 B.n414 B.n413 10.6151
R1120 B.n413 B.n8 10.6151
R1121 B.n360 B.n359 8.74196
R1122 B.n342 B.n36 8.74196
R1123 B.n185 B.n184 8.74196
R1124 B.n202 B.n85 8.74196
R1125 B.n431 B.n0 2.81026
R1126 B.n431 B.n1 2.81026
R1127 B.n359 B.n358 1.87367
R1128 B.n36 B.n32 1.87367
R1129 B.n186 B.n185 1.87367
R1130 B.n199 B.n85 1.87367
R1131 VP.n0 VP.t1 695.327
R1132 VP.n0 VP.t0 658.029
R1133 VP VP.n0 0.0516364
R1134 VDD1.n46 VDD1.n0 756.745
R1135 VDD1.n97 VDD1.n51 756.745
R1136 VDD1.n47 VDD1.n46 585
R1137 VDD1.n45 VDD1.n44 585
R1138 VDD1.n4 VDD1.n3 585
R1139 VDD1.n39 VDD1.n38 585
R1140 VDD1.n37 VDD1.n36 585
R1141 VDD1.n8 VDD1.n7 585
R1142 VDD1.n31 VDD1.n30 585
R1143 VDD1.n29 VDD1.n28 585
R1144 VDD1.n12 VDD1.n11 585
R1145 VDD1.n23 VDD1.n22 585
R1146 VDD1.n21 VDD1.n20 585
R1147 VDD1.n16 VDD1.n15 585
R1148 VDD1.n67 VDD1.n66 585
R1149 VDD1.n72 VDD1.n71 585
R1150 VDD1.n74 VDD1.n73 585
R1151 VDD1.n63 VDD1.n62 585
R1152 VDD1.n80 VDD1.n79 585
R1153 VDD1.n82 VDD1.n81 585
R1154 VDD1.n59 VDD1.n58 585
R1155 VDD1.n88 VDD1.n87 585
R1156 VDD1.n90 VDD1.n89 585
R1157 VDD1.n55 VDD1.n54 585
R1158 VDD1.n96 VDD1.n95 585
R1159 VDD1.n98 VDD1.n97 585
R1160 VDD1.n68 VDD1.t1 327.467
R1161 VDD1.n17 VDD1.t0 327.467
R1162 VDD1.n46 VDD1.n45 171.744
R1163 VDD1.n45 VDD1.n3 171.744
R1164 VDD1.n38 VDD1.n3 171.744
R1165 VDD1.n38 VDD1.n37 171.744
R1166 VDD1.n37 VDD1.n7 171.744
R1167 VDD1.n30 VDD1.n7 171.744
R1168 VDD1.n30 VDD1.n29 171.744
R1169 VDD1.n29 VDD1.n11 171.744
R1170 VDD1.n22 VDD1.n11 171.744
R1171 VDD1.n22 VDD1.n21 171.744
R1172 VDD1.n21 VDD1.n15 171.744
R1173 VDD1.n72 VDD1.n66 171.744
R1174 VDD1.n73 VDD1.n72 171.744
R1175 VDD1.n73 VDD1.n62 171.744
R1176 VDD1.n80 VDD1.n62 171.744
R1177 VDD1.n81 VDD1.n80 171.744
R1178 VDD1.n81 VDD1.n58 171.744
R1179 VDD1.n88 VDD1.n58 171.744
R1180 VDD1.n89 VDD1.n88 171.744
R1181 VDD1.n89 VDD1.n54 171.744
R1182 VDD1.n96 VDD1.n54 171.744
R1183 VDD1.n97 VDD1.n96 171.744
R1184 VDD1.t0 VDD1.n15 85.8723
R1185 VDD1.t1 VDD1.n66 85.8723
R1186 VDD1 VDD1.n101 80.5983
R1187 VDD1 VDD1.n50 46.7826
R1188 VDD1.n17 VDD1.n16 16.3895
R1189 VDD1.n68 VDD1.n67 16.3895
R1190 VDD1.n20 VDD1.n19 12.8005
R1191 VDD1.n71 VDD1.n70 12.8005
R1192 VDD1.n23 VDD1.n14 12.0247
R1193 VDD1.n74 VDD1.n65 12.0247
R1194 VDD1.n24 VDD1.n12 11.249
R1195 VDD1.n75 VDD1.n63 11.249
R1196 VDD1.n28 VDD1.n27 10.4732
R1197 VDD1.n79 VDD1.n78 10.4732
R1198 VDD1.n50 VDD1.n0 9.69747
R1199 VDD1.n31 VDD1.n10 9.69747
R1200 VDD1.n82 VDD1.n61 9.69747
R1201 VDD1.n101 VDD1.n51 9.69747
R1202 VDD1.n50 VDD1.n49 9.45567
R1203 VDD1.n101 VDD1.n100 9.45567
R1204 VDD1.n2 VDD1.n1 9.3005
R1205 VDD1.n43 VDD1.n42 9.3005
R1206 VDD1.n41 VDD1.n40 9.3005
R1207 VDD1.n6 VDD1.n5 9.3005
R1208 VDD1.n35 VDD1.n34 9.3005
R1209 VDD1.n33 VDD1.n32 9.3005
R1210 VDD1.n10 VDD1.n9 9.3005
R1211 VDD1.n27 VDD1.n26 9.3005
R1212 VDD1.n25 VDD1.n24 9.3005
R1213 VDD1.n14 VDD1.n13 9.3005
R1214 VDD1.n19 VDD1.n18 9.3005
R1215 VDD1.n49 VDD1.n48 9.3005
R1216 VDD1.n92 VDD1.n91 9.3005
R1217 VDD1.n94 VDD1.n93 9.3005
R1218 VDD1.n53 VDD1.n52 9.3005
R1219 VDD1.n100 VDD1.n99 9.3005
R1220 VDD1.n86 VDD1.n85 9.3005
R1221 VDD1.n84 VDD1.n83 9.3005
R1222 VDD1.n61 VDD1.n60 9.3005
R1223 VDD1.n78 VDD1.n77 9.3005
R1224 VDD1.n76 VDD1.n75 9.3005
R1225 VDD1.n65 VDD1.n64 9.3005
R1226 VDD1.n70 VDD1.n69 9.3005
R1227 VDD1.n57 VDD1.n56 9.3005
R1228 VDD1.n48 VDD1.n47 8.92171
R1229 VDD1.n32 VDD1.n8 8.92171
R1230 VDD1.n83 VDD1.n59 8.92171
R1231 VDD1.n99 VDD1.n98 8.92171
R1232 VDD1.n44 VDD1.n2 8.14595
R1233 VDD1.n36 VDD1.n35 8.14595
R1234 VDD1.n87 VDD1.n86 8.14595
R1235 VDD1.n95 VDD1.n53 8.14595
R1236 VDD1.n43 VDD1.n4 7.3702
R1237 VDD1.n39 VDD1.n6 7.3702
R1238 VDD1.n90 VDD1.n57 7.3702
R1239 VDD1.n94 VDD1.n55 7.3702
R1240 VDD1.n40 VDD1.n4 6.59444
R1241 VDD1.n40 VDD1.n39 6.59444
R1242 VDD1.n91 VDD1.n90 6.59444
R1243 VDD1.n91 VDD1.n55 6.59444
R1244 VDD1.n44 VDD1.n43 5.81868
R1245 VDD1.n36 VDD1.n6 5.81868
R1246 VDD1.n87 VDD1.n57 5.81868
R1247 VDD1.n95 VDD1.n94 5.81868
R1248 VDD1.n47 VDD1.n2 5.04292
R1249 VDD1.n35 VDD1.n8 5.04292
R1250 VDD1.n86 VDD1.n59 5.04292
R1251 VDD1.n98 VDD1.n53 5.04292
R1252 VDD1.n48 VDD1.n0 4.26717
R1253 VDD1.n32 VDD1.n31 4.26717
R1254 VDD1.n83 VDD1.n82 4.26717
R1255 VDD1.n99 VDD1.n51 4.26717
R1256 VDD1.n69 VDD1.n68 3.70984
R1257 VDD1.n18 VDD1.n17 3.70984
R1258 VDD1.n28 VDD1.n10 3.49141
R1259 VDD1.n79 VDD1.n61 3.49141
R1260 VDD1.n27 VDD1.n12 2.71565
R1261 VDD1.n78 VDD1.n63 2.71565
R1262 VDD1.n24 VDD1.n23 1.93989
R1263 VDD1.n75 VDD1.n74 1.93989
R1264 VDD1.n20 VDD1.n14 1.16414
R1265 VDD1.n71 VDD1.n65 1.16414
R1266 VDD1.n19 VDD1.n16 0.388379
R1267 VDD1.n70 VDD1.n67 0.388379
R1268 VDD1.n49 VDD1.n1 0.155672
R1269 VDD1.n42 VDD1.n1 0.155672
R1270 VDD1.n42 VDD1.n41 0.155672
R1271 VDD1.n41 VDD1.n5 0.155672
R1272 VDD1.n34 VDD1.n5 0.155672
R1273 VDD1.n34 VDD1.n33 0.155672
R1274 VDD1.n33 VDD1.n9 0.155672
R1275 VDD1.n26 VDD1.n9 0.155672
R1276 VDD1.n26 VDD1.n25 0.155672
R1277 VDD1.n25 VDD1.n13 0.155672
R1278 VDD1.n18 VDD1.n13 0.155672
R1279 VDD1.n69 VDD1.n64 0.155672
R1280 VDD1.n76 VDD1.n64 0.155672
R1281 VDD1.n77 VDD1.n76 0.155672
R1282 VDD1.n77 VDD1.n60 0.155672
R1283 VDD1.n84 VDD1.n60 0.155672
R1284 VDD1.n85 VDD1.n84 0.155672
R1285 VDD1.n85 VDD1.n56 0.155672
R1286 VDD1.n92 VDD1.n56 0.155672
R1287 VDD1.n93 VDD1.n92 0.155672
R1288 VDD1.n93 VDD1.n52 0.155672
R1289 VDD1.n100 VDD1.n52 0.155672
C0 VP VDD1 1.56888f
C1 w_n1318_n2868# VTAIL 2.5315f
C2 VTAIL VN 1.05348f
C3 w_n1318_n2868# VP 1.76794f
C4 VN VP 4.02476f
C5 VDD2 VTAIL 5.01563f
C6 w_n1318_n2868# VDD1 1.36776f
C7 VDD2 VP 0.247619f
C8 VN VDD1 0.148182f
C9 VDD2 VDD1 0.446474f
C10 B VTAIL 2.19142f
C11 B VP 0.928511f
C12 w_n1318_n2868# VN 1.60449f
C13 B VDD1 1.20491f
C14 VDD2 w_n1318_n2868# 1.3708f
C15 VDD2 VN 1.47313f
C16 B w_n1318_n2868# 5.88008f
C17 B VN 0.668062f
C18 B VDD2 1.21833f
C19 VTAIL VP 1.06803f
C20 VTAIL VDD1 4.982f
C21 VDD2 VSUBS 0.644279f
C22 VDD1 VSUBS 2.375414f
C23 VTAIL VSUBS 0.253581f
C24 VN VSUBS 4.23541f
C25 VP VSUBS 0.966114f
C26 B VSUBS 2.166998f
C27 w_n1318_n2868# VSUBS 46.7363f
C28 VDD1.n0 VSUBS 0.018493f
C29 VDD1.n1 VSUBS 0.016386f
C30 VDD1.n2 VSUBS 0.008805f
C31 VDD1.n3 VSUBS 0.020813f
C32 VDD1.n4 VSUBS 0.009323f
C33 VDD1.n5 VSUBS 0.016386f
C34 VDD1.n6 VSUBS 0.008805f
C35 VDD1.n7 VSUBS 0.020813f
C36 VDD1.n8 VSUBS 0.009323f
C37 VDD1.n9 VSUBS 0.016386f
C38 VDD1.n10 VSUBS 0.008805f
C39 VDD1.n11 VSUBS 0.020813f
C40 VDD1.n12 VSUBS 0.009323f
C41 VDD1.n13 VSUBS 0.016386f
C42 VDD1.n14 VSUBS 0.008805f
C43 VDD1.n15 VSUBS 0.01561f
C44 VDD1.n16 VSUBS 0.01324f
C45 VDD1.t0 VSUBS 0.04437f
C46 VDD1.n17 VSUBS 0.088869f
C47 VDD1.n18 VSUBS 0.6356f
C48 VDD1.n19 VSUBS 0.008805f
C49 VDD1.n20 VSUBS 0.009323f
C50 VDD1.n21 VSUBS 0.020813f
C51 VDD1.n22 VSUBS 0.020813f
C52 VDD1.n23 VSUBS 0.009323f
C53 VDD1.n24 VSUBS 0.008805f
C54 VDD1.n25 VSUBS 0.016386f
C55 VDD1.n26 VSUBS 0.016386f
C56 VDD1.n27 VSUBS 0.008805f
C57 VDD1.n28 VSUBS 0.009323f
C58 VDD1.n29 VSUBS 0.020813f
C59 VDD1.n30 VSUBS 0.020813f
C60 VDD1.n31 VSUBS 0.009323f
C61 VDD1.n32 VSUBS 0.008805f
C62 VDD1.n33 VSUBS 0.016386f
C63 VDD1.n34 VSUBS 0.016386f
C64 VDD1.n35 VSUBS 0.008805f
C65 VDD1.n36 VSUBS 0.009323f
C66 VDD1.n37 VSUBS 0.020813f
C67 VDD1.n38 VSUBS 0.020813f
C68 VDD1.n39 VSUBS 0.009323f
C69 VDD1.n40 VSUBS 0.008805f
C70 VDD1.n41 VSUBS 0.016386f
C71 VDD1.n42 VSUBS 0.016386f
C72 VDD1.n43 VSUBS 0.008805f
C73 VDD1.n44 VSUBS 0.009323f
C74 VDD1.n45 VSUBS 0.020813f
C75 VDD1.n46 VSUBS 0.052045f
C76 VDD1.n47 VSUBS 0.009323f
C77 VDD1.n48 VSUBS 0.008805f
C78 VDD1.n49 VSUBS 0.03519f
C79 VDD1.n50 VSUBS 0.037725f
C80 VDD1.n51 VSUBS 0.018493f
C81 VDD1.n52 VSUBS 0.016386f
C82 VDD1.n53 VSUBS 0.008805f
C83 VDD1.n54 VSUBS 0.020813f
C84 VDD1.n55 VSUBS 0.009323f
C85 VDD1.n56 VSUBS 0.016386f
C86 VDD1.n57 VSUBS 0.008805f
C87 VDD1.n58 VSUBS 0.020813f
C88 VDD1.n59 VSUBS 0.009323f
C89 VDD1.n60 VSUBS 0.016386f
C90 VDD1.n61 VSUBS 0.008805f
C91 VDD1.n62 VSUBS 0.020813f
C92 VDD1.n63 VSUBS 0.009323f
C93 VDD1.n64 VSUBS 0.016386f
C94 VDD1.n65 VSUBS 0.008805f
C95 VDD1.n66 VSUBS 0.01561f
C96 VDD1.n67 VSUBS 0.01324f
C97 VDD1.t1 VSUBS 0.04437f
C98 VDD1.n68 VSUBS 0.088869f
C99 VDD1.n69 VSUBS 0.6356f
C100 VDD1.n70 VSUBS 0.008805f
C101 VDD1.n71 VSUBS 0.009323f
C102 VDD1.n72 VSUBS 0.020813f
C103 VDD1.n73 VSUBS 0.020813f
C104 VDD1.n74 VSUBS 0.009323f
C105 VDD1.n75 VSUBS 0.008805f
C106 VDD1.n76 VSUBS 0.016386f
C107 VDD1.n77 VSUBS 0.016386f
C108 VDD1.n78 VSUBS 0.008805f
C109 VDD1.n79 VSUBS 0.009323f
C110 VDD1.n80 VSUBS 0.020813f
C111 VDD1.n81 VSUBS 0.020813f
C112 VDD1.n82 VSUBS 0.009323f
C113 VDD1.n83 VSUBS 0.008805f
C114 VDD1.n84 VSUBS 0.016386f
C115 VDD1.n85 VSUBS 0.016386f
C116 VDD1.n86 VSUBS 0.008805f
C117 VDD1.n87 VSUBS 0.009323f
C118 VDD1.n88 VSUBS 0.020813f
C119 VDD1.n89 VSUBS 0.020813f
C120 VDD1.n90 VSUBS 0.009323f
C121 VDD1.n91 VSUBS 0.008805f
C122 VDD1.n92 VSUBS 0.016386f
C123 VDD1.n93 VSUBS 0.016386f
C124 VDD1.n94 VSUBS 0.008805f
C125 VDD1.n95 VSUBS 0.009323f
C126 VDD1.n96 VSUBS 0.020813f
C127 VDD1.n97 VSUBS 0.052045f
C128 VDD1.n98 VSUBS 0.009323f
C129 VDD1.n99 VSUBS 0.008805f
C130 VDD1.n100 VSUBS 0.03519f
C131 VDD1.n101 VSUBS 0.372797f
C132 VP.t1 VSUBS 0.664485f
C133 VP.t0 VSUBS 0.589791f
C134 VP.n0 VSUBS 2.7366f
C135 B.n0 VSUBS 0.005041f
C136 B.n1 VSUBS 0.005041f
C137 B.n2 VSUBS 0.007971f
C138 B.n3 VSUBS 0.007971f
C139 B.n4 VSUBS 0.007971f
C140 B.n5 VSUBS 0.007971f
C141 B.n6 VSUBS 0.007971f
C142 B.n7 VSUBS 0.007971f
C143 B.n8 VSUBS 0.019154f
C144 B.n9 VSUBS 0.007971f
C145 B.n10 VSUBS 0.007971f
C146 B.n11 VSUBS 0.007971f
C147 B.n12 VSUBS 0.007971f
C148 B.n13 VSUBS 0.007971f
C149 B.n14 VSUBS 0.007971f
C150 B.n15 VSUBS 0.007971f
C151 B.n16 VSUBS 0.007971f
C152 B.n17 VSUBS 0.007971f
C153 B.n18 VSUBS 0.007971f
C154 B.n19 VSUBS 0.007971f
C155 B.n20 VSUBS 0.007971f
C156 B.n21 VSUBS 0.007971f
C157 B.n22 VSUBS 0.007971f
C158 B.n23 VSUBS 0.007971f
C159 B.n24 VSUBS 0.007971f
C160 B.n25 VSUBS 0.007971f
C161 B.t8 VSUBS 0.178607f
C162 B.t7 VSUBS 0.189472f
C163 B.t6 VSUBS 0.239712f
C164 B.n26 VSUBS 0.28024f
C165 B.n27 VSUBS 0.235015f
C166 B.n28 VSUBS 0.007971f
C167 B.n29 VSUBS 0.007971f
C168 B.n30 VSUBS 0.007971f
C169 B.n31 VSUBS 0.007971f
C170 B.n32 VSUBS 0.004689f
C171 B.n33 VSUBS 0.007971f
C172 B.t11 VSUBS 0.17861f
C173 B.t10 VSUBS 0.189475f
C174 B.t9 VSUBS 0.239712f
C175 B.n34 VSUBS 0.280237f
C176 B.n35 VSUBS 0.235012f
C177 B.n36 VSUBS 0.018469f
C178 B.n37 VSUBS 0.007971f
C179 B.n38 VSUBS 0.007971f
C180 B.n39 VSUBS 0.007971f
C181 B.n40 VSUBS 0.007971f
C182 B.n41 VSUBS 0.007971f
C183 B.n42 VSUBS 0.007971f
C184 B.n43 VSUBS 0.007971f
C185 B.n44 VSUBS 0.007971f
C186 B.n45 VSUBS 0.007971f
C187 B.n46 VSUBS 0.007971f
C188 B.n47 VSUBS 0.007971f
C189 B.n48 VSUBS 0.007971f
C190 B.n49 VSUBS 0.007971f
C191 B.n50 VSUBS 0.007971f
C192 B.n51 VSUBS 0.007971f
C193 B.n52 VSUBS 0.020234f
C194 B.n53 VSUBS 0.007971f
C195 B.n54 VSUBS 0.007971f
C196 B.n55 VSUBS 0.007971f
C197 B.n56 VSUBS 0.007971f
C198 B.n57 VSUBS 0.007971f
C199 B.n58 VSUBS 0.007971f
C200 B.n59 VSUBS 0.007971f
C201 B.n60 VSUBS 0.007971f
C202 B.n61 VSUBS 0.007971f
C203 B.n62 VSUBS 0.007971f
C204 B.n63 VSUBS 0.007971f
C205 B.n64 VSUBS 0.007971f
C206 B.n65 VSUBS 0.007971f
C207 B.n66 VSUBS 0.020234f
C208 B.n67 VSUBS 0.007971f
C209 B.n68 VSUBS 0.007971f
C210 B.n69 VSUBS 0.007971f
C211 B.n70 VSUBS 0.007971f
C212 B.n71 VSUBS 0.007971f
C213 B.n72 VSUBS 0.007971f
C214 B.n73 VSUBS 0.007971f
C215 B.n74 VSUBS 0.007971f
C216 B.n75 VSUBS 0.007971f
C217 B.n76 VSUBS 0.007971f
C218 B.n77 VSUBS 0.007971f
C219 B.n78 VSUBS 0.007971f
C220 B.n79 VSUBS 0.007971f
C221 B.n80 VSUBS 0.007971f
C222 B.n81 VSUBS 0.007971f
C223 B.n82 VSUBS 0.007971f
C224 B.t1 VSUBS 0.17861f
C225 B.t2 VSUBS 0.189475f
C226 B.t0 VSUBS 0.239712f
C227 B.n83 VSUBS 0.280237f
C228 B.n84 VSUBS 0.235012f
C229 B.n85 VSUBS 0.018469f
C230 B.n86 VSUBS 0.007971f
C231 B.n87 VSUBS 0.007971f
C232 B.n88 VSUBS 0.007971f
C233 B.n89 VSUBS 0.007971f
C234 B.n90 VSUBS 0.007971f
C235 B.t4 VSUBS 0.178607f
C236 B.t5 VSUBS 0.189472f
C237 B.t3 VSUBS 0.239712f
C238 B.n91 VSUBS 0.28024f
C239 B.n92 VSUBS 0.235015f
C240 B.n93 VSUBS 0.007971f
C241 B.n94 VSUBS 0.007971f
C242 B.n95 VSUBS 0.007971f
C243 B.n96 VSUBS 0.007971f
C244 B.n97 VSUBS 0.007971f
C245 B.n98 VSUBS 0.007971f
C246 B.n99 VSUBS 0.007971f
C247 B.n100 VSUBS 0.007971f
C248 B.n101 VSUBS 0.007971f
C249 B.n102 VSUBS 0.007971f
C250 B.n103 VSUBS 0.007971f
C251 B.n104 VSUBS 0.007971f
C252 B.n105 VSUBS 0.007971f
C253 B.n106 VSUBS 0.007971f
C254 B.n107 VSUBS 0.007971f
C255 B.n108 VSUBS 0.007971f
C256 B.n109 VSUBS 0.020234f
C257 B.n110 VSUBS 0.007971f
C258 B.n111 VSUBS 0.007971f
C259 B.n112 VSUBS 0.007971f
C260 B.n113 VSUBS 0.007971f
C261 B.n114 VSUBS 0.007971f
C262 B.n115 VSUBS 0.007971f
C263 B.n116 VSUBS 0.007971f
C264 B.n117 VSUBS 0.007971f
C265 B.n118 VSUBS 0.007971f
C266 B.n119 VSUBS 0.007971f
C267 B.n120 VSUBS 0.007971f
C268 B.n121 VSUBS 0.007971f
C269 B.n122 VSUBS 0.007971f
C270 B.n123 VSUBS 0.007971f
C271 B.n124 VSUBS 0.007971f
C272 B.n125 VSUBS 0.007971f
C273 B.n126 VSUBS 0.007971f
C274 B.n127 VSUBS 0.007971f
C275 B.n128 VSUBS 0.007971f
C276 B.n129 VSUBS 0.007971f
C277 B.n130 VSUBS 0.007971f
C278 B.n131 VSUBS 0.007971f
C279 B.n132 VSUBS 0.019154f
C280 B.n133 VSUBS 0.019154f
C281 B.n134 VSUBS 0.020234f
C282 B.n135 VSUBS 0.007971f
C283 B.n136 VSUBS 0.007971f
C284 B.n137 VSUBS 0.007971f
C285 B.n138 VSUBS 0.007971f
C286 B.n139 VSUBS 0.007971f
C287 B.n140 VSUBS 0.007971f
C288 B.n141 VSUBS 0.007971f
C289 B.n142 VSUBS 0.007971f
C290 B.n143 VSUBS 0.007971f
C291 B.n144 VSUBS 0.007971f
C292 B.n145 VSUBS 0.007971f
C293 B.n146 VSUBS 0.007971f
C294 B.n147 VSUBS 0.007971f
C295 B.n148 VSUBS 0.007971f
C296 B.n149 VSUBS 0.007971f
C297 B.n150 VSUBS 0.007971f
C298 B.n151 VSUBS 0.007971f
C299 B.n152 VSUBS 0.007971f
C300 B.n153 VSUBS 0.007971f
C301 B.n154 VSUBS 0.007971f
C302 B.n155 VSUBS 0.007971f
C303 B.n156 VSUBS 0.007971f
C304 B.n157 VSUBS 0.007971f
C305 B.n158 VSUBS 0.007971f
C306 B.n159 VSUBS 0.007971f
C307 B.n160 VSUBS 0.007971f
C308 B.n161 VSUBS 0.007971f
C309 B.n162 VSUBS 0.007971f
C310 B.n163 VSUBS 0.007971f
C311 B.n164 VSUBS 0.007971f
C312 B.n165 VSUBS 0.007971f
C313 B.n166 VSUBS 0.007971f
C314 B.n167 VSUBS 0.007971f
C315 B.n168 VSUBS 0.007971f
C316 B.n169 VSUBS 0.007971f
C317 B.n170 VSUBS 0.007971f
C318 B.n171 VSUBS 0.007971f
C319 B.n172 VSUBS 0.007971f
C320 B.n173 VSUBS 0.007971f
C321 B.n174 VSUBS 0.007971f
C322 B.n175 VSUBS 0.007971f
C323 B.n176 VSUBS 0.007971f
C324 B.n177 VSUBS 0.007971f
C325 B.n178 VSUBS 0.007971f
C326 B.n179 VSUBS 0.007971f
C327 B.n180 VSUBS 0.007971f
C328 B.n181 VSUBS 0.007971f
C329 B.n182 VSUBS 0.007971f
C330 B.n183 VSUBS 0.007971f
C331 B.n184 VSUBS 0.007268f
C332 B.n185 VSUBS 0.018469f
C333 B.n186 VSUBS 0.004689f
C334 B.n187 VSUBS 0.007971f
C335 B.n188 VSUBS 0.007971f
C336 B.n189 VSUBS 0.007971f
C337 B.n190 VSUBS 0.007971f
C338 B.n191 VSUBS 0.007971f
C339 B.n192 VSUBS 0.007971f
C340 B.n193 VSUBS 0.007971f
C341 B.n194 VSUBS 0.007971f
C342 B.n195 VSUBS 0.007971f
C343 B.n196 VSUBS 0.007971f
C344 B.n197 VSUBS 0.007971f
C345 B.n198 VSUBS 0.007971f
C346 B.n199 VSUBS 0.004689f
C347 B.n200 VSUBS 0.007971f
C348 B.n201 VSUBS 0.007971f
C349 B.n202 VSUBS 0.007268f
C350 B.n203 VSUBS 0.007971f
C351 B.n204 VSUBS 0.007971f
C352 B.n205 VSUBS 0.007971f
C353 B.n206 VSUBS 0.007971f
C354 B.n207 VSUBS 0.007971f
C355 B.n208 VSUBS 0.007971f
C356 B.n209 VSUBS 0.007971f
C357 B.n210 VSUBS 0.007971f
C358 B.n211 VSUBS 0.007971f
C359 B.n212 VSUBS 0.007971f
C360 B.n213 VSUBS 0.007971f
C361 B.n214 VSUBS 0.007971f
C362 B.n215 VSUBS 0.007971f
C363 B.n216 VSUBS 0.007971f
C364 B.n217 VSUBS 0.007971f
C365 B.n218 VSUBS 0.007971f
C366 B.n219 VSUBS 0.007971f
C367 B.n220 VSUBS 0.007971f
C368 B.n221 VSUBS 0.007971f
C369 B.n222 VSUBS 0.007971f
C370 B.n223 VSUBS 0.007971f
C371 B.n224 VSUBS 0.007971f
C372 B.n225 VSUBS 0.007971f
C373 B.n226 VSUBS 0.007971f
C374 B.n227 VSUBS 0.007971f
C375 B.n228 VSUBS 0.007971f
C376 B.n229 VSUBS 0.007971f
C377 B.n230 VSUBS 0.007971f
C378 B.n231 VSUBS 0.007971f
C379 B.n232 VSUBS 0.007971f
C380 B.n233 VSUBS 0.007971f
C381 B.n234 VSUBS 0.007971f
C382 B.n235 VSUBS 0.007971f
C383 B.n236 VSUBS 0.007971f
C384 B.n237 VSUBS 0.007971f
C385 B.n238 VSUBS 0.007971f
C386 B.n239 VSUBS 0.007971f
C387 B.n240 VSUBS 0.007971f
C388 B.n241 VSUBS 0.007971f
C389 B.n242 VSUBS 0.007971f
C390 B.n243 VSUBS 0.007971f
C391 B.n244 VSUBS 0.007971f
C392 B.n245 VSUBS 0.007971f
C393 B.n246 VSUBS 0.007971f
C394 B.n247 VSUBS 0.007971f
C395 B.n248 VSUBS 0.007971f
C396 B.n249 VSUBS 0.007971f
C397 B.n250 VSUBS 0.007971f
C398 B.n251 VSUBS 0.020234f
C399 B.n252 VSUBS 0.019154f
C400 B.n253 VSUBS 0.019154f
C401 B.n254 VSUBS 0.007971f
C402 B.n255 VSUBS 0.007971f
C403 B.n256 VSUBS 0.007971f
C404 B.n257 VSUBS 0.007971f
C405 B.n258 VSUBS 0.007971f
C406 B.n259 VSUBS 0.007971f
C407 B.n260 VSUBS 0.007971f
C408 B.n261 VSUBS 0.007971f
C409 B.n262 VSUBS 0.007971f
C410 B.n263 VSUBS 0.007971f
C411 B.n264 VSUBS 0.007971f
C412 B.n265 VSUBS 0.007971f
C413 B.n266 VSUBS 0.007971f
C414 B.n267 VSUBS 0.007971f
C415 B.n268 VSUBS 0.007971f
C416 B.n269 VSUBS 0.007971f
C417 B.n270 VSUBS 0.007971f
C418 B.n271 VSUBS 0.007971f
C419 B.n272 VSUBS 0.007971f
C420 B.n273 VSUBS 0.007971f
C421 B.n274 VSUBS 0.007971f
C422 B.n275 VSUBS 0.007971f
C423 B.n276 VSUBS 0.007971f
C424 B.n277 VSUBS 0.007971f
C425 B.n278 VSUBS 0.007971f
C426 B.n279 VSUBS 0.007971f
C427 B.n280 VSUBS 0.007971f
C428 B.n281 VSUBS 0.007971f
C429 B.n282 VSUBS 0.007971f
C430 B.n283 VSUBS 0.007971f
C431 B.n284 VSUBS 0.007971f
C432 B.n285 VSUBS 0.007971f
C433 B.n286 VSUBS 0.007971f
C434 B.n287 VSUBS 0.007971f
C435 B.n288 VSUBS 0.007971f
C436 B.n289 VSUBS 0.007971f
C437 B.n290 VSUBS 0.007971f
C438 B.n291 VSUBS 0.019154f
C439 B.n292 VSUBS 0.020022f
C440 B.n293 VSUBS 0.019366f
C441 B.n294 VSUBS 0.007971f
C442 B.n295 VSUBS 0.007971f
C443 B.n296 VSUBS 0.007971f
C444 B.n297 VSUBS 0.007971f
C445 B.n298 VSUBS 0.007971f
C446 B.n299 VSUBS 0.007971f
C447 B.n300 VSUBS 0.007971f
C448 B.n301 VSUBS 0.007971f
C449 B.n302 VSUBS 0.007971f
C450 B.n303 VSUBS 0.007971f
C451 B.n304 VSUBS 0.007971f
C452 B.n305 VSUBS 0.007971f
C453 B.n306 VSUBS 0.007971f
C454 B.n307 VSUBS 0.007971f
C455 B.n308 VSUBS 0.007971f
C456 B.n309 VSUBS 0.007971f
C457 B.n310 VSUBS 0.007971f
C458 B.n311 VSUBS 0.007971f
C459 B.n312 VSUBS 0.007971f
C460 B.n313 VSUBS 0.007971f
C461 B.n314 VSUBS 0.007971f
C462 B.n315 VSUBS 0.007971f
C463 B.n316 VSUBS 0.007971f
C464 B.n317 VSUBS 0.007971f
C465 B.n318 VSUBS 0.007971f
C466 B.n319 VSUBS 0.007971f
C467 B.n320 VSUBS 0.007971f
C468 B.n321 VSUBS 0.007971f
C469 B.n322 VSUBS 0.007971f
C470 B.n323 VSUBS 0.007971f
C471 B.n324 VSUBS 0.007971f
C472 B.n325 VSUBS 0.007971f
C473 B.n326 VSUBS 0.007971f
C474 B.n327 VSUBS 0.007971f
C475 B.n328 VSUBS 0.007971f
C476 B.n329 VSUBS 0.007971f
C477 B.n330 VSUBS 0.007971f
C478 B.n331 VSUBS 0.007971f
C479 B.n332 VSUBS 0.007971f
C480 B.n333 VSUBS 0.007971f
C481 B.n334 VSUBS 0.007971f
C482 B.n335 VSUBS 0.007971f
C483 B.n336 VSUBS 0.007971f
C484 B.n337 VSUBS 0.007971f
C485 B.n338 VSUBS 0.007971f
C486 B.n339 VSUBS 0.007971f
C487 B.n340 VSUBS 0.007971f
C488 B.n341 VSUBS 0.007971f
C489 B.n342 VSUBS 0.007268f
C490 B.n343 VSUBS 0.007971f
C491 B.n344 VSUBS 0.007971f
C492 B.n345 VSUBS 0.007971f
C493 B.n346 VSUBS 0.007971f
C494 B.n347 VSUBS 0.007971f
C495 B.n348 VSUBS 0.007971f
C496 B.n349 VSUBS 0.007971f
C497 B.n350 VSUBS 0.007971f
C498 B.n351 VSUBS 0.007971f
C499 B.n352 VSUBS 0.007971f
C500 B.n353 VSUBS 0.007971f
C501 B.n354 VSUBS 0.007971f
C502 B.n355 VSUBS 0.007971f
C503 B.n356 VSUBS 0.007971f
C504 B.n357 VSUBS 0.007971f
C505 B.n358 VSUBS 0.004689f
C506 B.n359 VSUBS 0.018469f
C507 B.n360 VSUBS 0.007268f
C508 B.n361 VSUBS 0.007971f
C509 B.n362 VSUBS 0.007971f
C510 B.n363 VSUBS 0.007971f
C511 B.n364 VSUBS 0.007971f
C512 B.n365 VSUBS 0.007971f
C513 B.n366 VSUBS 0.007971f
C514 B.n367 VSUBS 0.007971f
C515 B.n368 VSUBS 0.007971f
C516 B.n369 VSUBS 0.007971f
C517 B.n370 VSUBS 0.007971f
C518 B.n371 VSUBS 0.007971f
C519 B.n372 VSUBS 0.007971f
C520 B.n373 VSUBS 0.007971f
C521 B.n374 VSUBS 0.007971f
C522 B.n375 VSUBS 0.007971f
C523 B.n376 VSUBS 0.007971f
C524 B.n377 VSUBS 0.007971f
C525 B.n378 VSUBS 0.007971f
C526 B.n379 VSUBS 0.007971f
C527 B.n380 VSUBS 0.007971f
C528 B.n381 VSUBS 0.007971f
C529 B.n382 VSUBS 0.007971f
C530 B.n383 VSUBS 0.007971f
C531 B.n384 VSUBS 0.007971f
C532 B.n385 VSUBS 0.007971f
C533 B.n386 VSUBS 0.007971f
C534 B.n387 VSUBS 0.007971f
C535 B.n388 VSUBS 0.007971f
C536 B.n389 VSUBS 0.007971f
C537 B.n390 VSUBS 0.007971f
C538 B.n391 VSUBS 0.007971f
C539 B.n392 VSUBS 0.007971f
C540 B.n393 VSUBS 0.007971f
C541 B.n394 VSUBS 0.007971f
C542 B.n395 VSUBS 0.007971f
C543 B.n396 VSUBS 0.007971f
C544 B.n397 VSUBS 0.007971f
C545 B.n398 VSUBS 0.007971f
C546 B.n399 VSUBS 0.007971f
C547 B.n400 VSUBS 0.007971f
C548 B.n401 VSUBS 0.007971f
C549 B.n402 VSUBS 0.007971f
C550 B.n403 VSUBS 0.007971f
C551 B.n404 VSUBS 0.007971f
C552 B.n405 VSUBS 0.007971f
C553 B.n406 VSUBS 0.007971f
C554 B.n407 VSUBS 0.007971f
C555 B.n408 VSUBS 0.007971f
C556 B.n409 VSUBS 0.020234f
C557 B.n410 VSUBS 0.020234f
C558 B.n411 VSUBS 0.019154f
C559 B.n412 VSUBS 0.007971f
C560 B.n413 VSUBS 0.007971f
C561 B.n414 VSUBS 0.007971f
C562 B.n415 VSUBS 0.007971f
C563 B.n416 VSUBS 0.007971f
C564 B.n417 VSUBS 0.007971f
C565 B.n418 VSUBS 0.007971f
C566 B.n419 VSUBS 0.007971f
C567 B.n420 VSUBS 0.007971f
C568 B.n421 VSUBS 0.007971f
C569 B.n422 VSUBS 0.007971f
C570 B.n423 VSUBS 0.007971f
C571 B.n424 VSUBS 0.007971f
C572 B.n425 VSUBS 0.007971f
C573 B.n426 VSUBS 0.007971f
C574 B.n427 VSUBS 0.007971f
C575 B.n428 VSUBS 0.007971f
C576 B.n429 VSUBS 0.007971f
C577 B.n430 VSUBS 0.007971f
C578 B.n431 VSUBS 0.01805f
C579 VDD2.n0 VSUBS 0.018719f
C580 VDD2.n1 VSUBS 0.016587f
C581 VDD2.n2 VSUBS 0.008913f
C582 VDD2.n3 VSUBS 0.021068f
C583 VDD2.n4 VSUBS 0.009438f
C584 VDD2.n5 VSUBS 0.016587f
C585 VDD2.n6 VSUBS 0.008913f
C586 VDD2.n7 VSUBS 0.021068f
C587 VDD2.n8 VSUBS 0.009438f
C588 VDD2.n9 VSUBS 0.016587f
C589 VDD2.n10 VSUBS 0.008913f
C590 VDD2.n11 VSUBS 0.021068f
C591 VDD2.n12 VSUBS 0.009438f
C592 VDD2.n13 VSUBS 0.016587f
C593 VDD2.n14 VSUBS 0.008913f
C594 VDD2.n15 VSUBS 0.015801f
C595 VDD2.n16 VSUBS 0.013402f
C596 VDD2.t1 VSUBS 0.044914f
C597 VDD2.n17 VSUBS 0.089958f
C598 VDD2.n18 VSUBS 0.643388f
C599 VDD2.n19 VSUBS 0.008913f
C600 VDD2.n20 VSUBS 0.009438f
C601 VDD2.n21 VSUBS 0.021068f
C602 VDD2.n22 VSUBS 0.021068f
C603 VDD2.n23 VSUBS 0.009438f
C604 VDD2.n24 VSUBS 0.008913f
C605 VDD2.n25 VSUBS 0.016587f
C606 VDD2.n26 VSUBS 0.016587f
C607 VDD2.n27 VSUBS 0.008913f
C608 VDD2.n28 VSUBS 0.009438f
C609 VDD2.n29 VSUBS 0.021068f
C610 VDD2.n30 VSUBS 0.021068f
C611 VDD2.n31 VSUBS 0.009438f
C612 VDD2.n32 VSUBS 0.008913f
C613 VDD2.n33 VSUBS 0.016587f
C614 VDD2.n34 VSUBS 0.016587f
C615 VDD2.n35 VSUBS 0.008913f
C616 VDD2.n36 VSUBS 0.009438f
C617 VDD2.n37 VSUBS 0.021068f
C618 VDD2.n38 VSUBS 0.021068f
C619 VDD2.n39 VSUBS 0.009438f
C620 VDD2.n40 VSUBS 0.008913f
C621 VDD2.n41 VSUBS 0.016587f
C622 VDD2.n42 VSUBS 0.016587f
C623 VDD2.n43 VSUBS 0.008913f
C624 VDD2.n44 VSUBS 0.009438f
C625 VDD2.n45 VSUBS 0.021068f
C626 VDD2.n46 VSUBS 0.052683f
C627 VDD2.n47 VSUBS 0.009438f
C628 VDD2.n48 VSUBS 0.008913f
C629 VDD2.n49 VSUBS 0.035622f
C630 VDD2.n50 VSUBS 0.356499f
C631 VDD2.n51 VSUBS 0.018719f
C632 VDD2.n52 VSUBS 0.016587f
C633 VDD2.n53 VSUBS 0.008913f
C634 VDD2.n54 VSUBS 0.021068f
C635 VDD2.n55 VSUBS 0.009438f
C636 VDD2.n56 VSUBS 0.016587f
C637 VDD2.n57 VSUBS 0.008913f
C638 VDD2.n58 VSUBS 0.021068f
C639 VDD2.n59 VSUBS 0.009438f
C640 VDD2.n60 VSUBS 0.016587f
C641 VDD2.n61 VSUBS 0.008913f
C642 VDD2.n62 VSUBS 0.021068f
C643 VDD2.n63 VSUBS 0.009438f
C644 VDD2.n64 VSUBS 0.016587f
C645 VDD2.n65 VSUBS 0.008913f
C646 VDD2.n66 VSUBS 0.015801f
C647 VDD2.n67 VSUBS 0.013402f
C648 VDD2.t0 VSUBS 0.044914f
C649 VDD2.n68 VSUBS 0.089958f
C650 VDD2.n69 VSUBS 0.643388f
C651 VDD2.n70 VSUBS 0.008913f
C652 VDD2.n71 VSUBS 0.009438f
C653 VDD2.n72 VSUBS 0.021068f
C654 VDD2.n73 VSUBS 0.021068f
C655 VDD2.n74 VSUBS 0.009438f
C656 VDD2.n75 VSUBS 0.008913f
C657 VDD2.n76 VSUBS 0.016587f
C658 VDD2.n77 VSUBS 0.016587f
C659 VDD2.n78 VSUBS 0.008913f
C660 VDD2.n79 VSUBS 0.009438f
C661 VDD2.n80 VSUBS 0.021068f
C662 VDD2.n81 VSUBS 0.021068f
C663 VDD2.n82 VSUBS 0.009438f
C664 VDD2.n83 VSUBS 0.008913f
C665 VDD2.n84 VSUBS 0.016587f
C666 VDD2.n85 VSUBS 0.016587f
C667 VDD2.n86 VSUBS 0.008913f
C668 VDD2.n87 VSUBS 0.009438f
C669 VDD2.n88 VSUBS 0.021068f
C670 VDD2.n89 VSUBS 0.021068f
C671 VDD2.n90 VSUBS 0.009438f
C672 VDD2.n91 VSUBS 0.008913f
C673 VDD2.n92 VSUBS 0.016587f
C674 VDD2.n93 VSUBS 0.016587f
C675 VDD2.n94 VSUBS 0.008913f
C676 VDD2.n95 VSUBS 0.009438f
C677 VDD2.n96 VSUBS 0.021068f
C678 VDD2.n97 VSUBS 0.052683f
C679 VDD2.n98 VSUBS 0.009438f
C680 VDD2.n99 VSUBS 0.008913f
C681 VDD2.n100 VSUBS 0.035622f
C682 VDD2.n101 VSUBS 0.037959f
C683 VDD2.n102 VSUBS 1.56829f
C684 VTAIL.n0 VSUBS 0.02979f
C685 VTAIL.n1 VSUBS 0.026397f
C686 VTAIL.n2 VSUBS 0.014185f
C687 VTAIL.n3 VSUBS 0.033528f
C688 VTAIL.n4 VSUBS 0.015019f
C689 VTAIL.n5 VSUBS 0.026397f
C690 VTAIL.n6 VSUBS 0.014185f
C691 VTAIL.n7 VSUBS 0.033528f
C692 VTAIL.n8 VSUBS 0.015019f
C693 VTAIL.n9 VSUBS 0.026397f
C694 VTAIL.n10 VSUBS 0.014185f
C695 VTAIL.n11 VSUBS 0.033528f
C696 VTAIL.n12 VSUBS 0.015019f
C697 VTAIL.n13 VSUBS 0.026397f
C698 VTAIL.n14 VSUBS 0.014185f
C699 VTAIL.n15 VSUBS 0.025146f
C700 VTAIL.n16 VSUBS 0.021329f
C701 VTAIL.t1 VSUBS 0.071477f
C702 VTAIL.n17 VSUBS 0.143162f
C703 VTAIL.n18 VSUBS 1.0239f
C704 VTAIL.n19 VSUBS 0.014185f
C705 VTAIL.n20 VSUBS 0.015019f
C706 VTAIL.n21 VSUBS 0.033528f
C707 VTAIL.n22 VSUBS 0.033528f
C708 VTAIL.n23 VSUBS 0.015019f
C709 VTAIL.n24 VSUBS 0.014185f
C710 VTAIL.n25 VSUBS 0.026397f
C711 VTAIL.n26 VSUBS 0.026397f
C712 VTAIL.n27 VSUBS 0.014185f
C713 VTAIL.n28 VSUBS 0.015019f
C714 VTAIL.n29 VSUBS 0.033528f
C715 VTAIL.n30 VSUBS 0.033528f
C716 VTAIL.n31 VSUBS 0.015019f
C717 VTAIL.n32 VSUBS 0.014185f
C718 VTAIL.n33 VSUBS 0.026397f
C719 VTAIL.n34 VSUBS 0.026397f
C720 VTAIL.n35 VSUBS 0.014185f
C721 VTAIL.n36 VSUBS 0.015019f
C722 VTAIL.n37 VSUBS 0.033528f
C723 VTAIL.n38 VSUBS 0.033528f
C724 VTAIL.n39 VSUBS 0.015019f
C725 VTAIL.n40 VSUBS 0.014185f
C726 VTAIL.n41 VSUBS 0.026397f
C727 VTAIL.n42 VSUBS 0.026397f
C728 VTAIL.n43 VSUBS 0.014185f
C729 VTAIL.n44 VSUBS 0.015019f
C730 VTAIL.n45 VSUBS 0.033528f
C731 VTAIL.n46 VSUBS 0.08384f
C732 VTAIL.n47 VSUBS 0.015019f
C733 VTAIL.n48 VSUBS 0.014185f
C734 VTAIL.n49 VSUBS 0.056689f
C735 VTAIL.n50 VSUBS 0.042144f
C736 VTAIL.n51 VSUBS 1.26373f
C737 VTAIL.n52 VSUBS 0.02979f
C738 VTAIL.n53 VSUBS 0.026397f
C739 VTAIL.n54 VSUBS 0.014185f
C740 VTAIL.n55 VSUBS 0.033528f
C741 VTAIL.n56 VSUBS 0.015019f
C742 VTAIL.n57 VSUBS 0.026397f
C743 VTAIL.n58 VSUBS 0.014185f
C744 VTAIL.n59 VSUBS 0.033528f
C745 VTAIL.n60 VSUBS 0.015019f
C746 VTAIL.n61 VSUBS 0.026397f
C747 VTAIL.n62 VSUBS 0.014185f
C748 VTAIL.n63 VSUBS 0.033528f
C749 VTAIL.n64 VSUBS 0.015019f
C750 VTAIL.n65 VSUBS 0.026397f
C751 VTAIL.n66 VSUBS 0.014185f
C752 VTAIL.n67 VSUBS 0.025146f
C753 VTAIL.n68 VSUBS 0.021329f
C754 VTAIL.t3 VSUBS 0.071477f
C755 VTAIL.n69 VSUBS 0.143162f
C756 VTAIL.n70 VSUBS 1.0239f
C757 VTAIL.n71 VSUBS 0.014185f
C758 VTAIL.n72 VSUBS 0.015019f
C759 VTAIL.n73 VSUBS 0.033528f
C760 VTAIL.n74 VSUBS 0.033528f
C761 VTAIL.n75 VSUBS 0.015019f
C762 VTAIL.n76 VSUBS 0.014185f
C763 VTAIL.n77 VSUBS 0.026397f
C764 VTAIL.n78 VSUBS 0.026397f
C765 VTAIL.n79 VSUBS 0.014185f
C766 VTAIL.n80 VSUBS 0.015019f
C767 VTAIL.n81 VSUBS 0.033528f
C768 VTAIL.n82 VSUBS 0.033528f
C769 VTAIL.n83 VSUBS 0.015019f
C770 VTAIL.n84 VSUBS 0.014185f
C771 VTAIL.n85 VSUBS 0.026397f
C772 VTAIL.n86 VSUBS 0.026397f
C773 VTAIL.n87 VSUBS 0.014185f
C774 VTAIL.n88 VSUBS 0.015019f
C775 VTAIL.n89 VSUBS 0.033528f
C776 VTAIL.n90 VSUBS 0.033528f
C777 VTAIL.n91 VSUBS 0.015019f
C778 VTAIL.n92 VSUBS 0.014185f
C779 VTAIL.n93 VSUBS 0.026397f
C780 VTAIL.n94 VSUBS 0.026397f
C781 VTAIL.n95 VSUBS 0.014185f
C782 VTAIL.n96 VSUBS 0.015019f
C783 VTAIL.n97 VSUBS 0.033528f
C784 VTAIL.n98 VSUBS 0.08384f
C785 VTAIL.n99 VSUBS 0.015019f
C786 VTAIL.n100 VSUBS 0.014185f
C787 VTAIL.n101 VSUBS 0.056689f
C788 VTAIL.n102 VSUBS 0.042144f
C789 VTAIL.n103 VSUBS 1.27473f
C790 VTAIL.n104 VSUBS 0.02979f
C791 VTAIL.n105 VSUBS 0.026397f
C792 VTAIL.n106 VSUBS 0.014185f
C793 VTAIL.n107 VSUBS 0.033528f
C794 VTAIL.n108 VSUBS 0.015019f
C795 VTAIL.n109 VSUBS 0.026397f
C796 VTAIL.n110 VSUBS 0.014185f
C797 VTAIL.n111 VSUBS 0.033528f
C798 VTAIL.n112 VSUBS 0.015019f
C799 VTAIL.n113 VSUBS 0.026397f
C800 VTAIL.n114 VSUBS 0.014185f
C801 VTAIL.n115 VSUBS 0.033528f
C802 VTAIL.n116 VSUBS 0.015019f
C803 VTAIL.n117 VSUBS 0.026397f
C804 VTAIL.n118 VSUBS 0.014185f
C805 VTAIL.n119 VSUBS 0.025146f
C806 VTAIL.n120 VSUBS 0.021329f
C807 VTAIL.t0 VSUBS 0.071477f
C808 VTAIL.n121 VSUBS 0.143162f
C809 VTAIL.n122 VSUBS 1.0239f
C810 VTAIL.n123 VSUBS 0.014185f
C811 VTAIL.n124 VSUBS 0.015019f
C812 VTAIL.n125 VSUBS 0.033528f
C813 VTAIL.n126 VSUBS 0.033528f
C814 VTAIL.n127 VSUBS 0.015019f
C815 VTAIL.n128 VSUBS 0.014185f
C816 VTAIL.n129 VSUBS 0.026397f
C817 VTAIL.n130 VSUBS 0.026397f
C818 VTAIL.n131 VSUBS 0.014185f
C819 VTAIL.n132 VSUBS 0.015019f
C820 VTAIL.n133 VSUBS 0.033528f
C821 VTAIL.n134 VSUBS 0.033528f
C822 VTAIL.n135 VSUBS 0.015019f
C823 VTAIL.n136 VSUBS 0.014185f
C824 VTAIL.n137 VSUBS 0.026397f
C825 VTAIL.n138 VSUBS 0.026397f
C826 VTAIL.n139 VSUBS 0.014185f
C827 VTAIL.n140 VSUBS 0.015019f
C828 VTAIL.n141 VSUBS 0.033528f
C829 VTAIL.n142 VSUBS 0.033528f
C830 VTAIL.n143 VSUBS 0.015019f
C831 VTAIL.n144 VSUBS 0.014185f
C832 VTAIL.n145 VSUBS 0.026397f
C833 VTAIL.n146 VSUBS 0.026397f
C834 VTAIL.n147 VSUBS 0.014185f
C835 VTAIL.n148 VSUBS 0.015019f
C836 VTAIL.n149 VSUBS 0.033528f
C837 VTAIL.n150 VSUBS 0.08384f
C838 VTAIL.n151 VSUBS 0.015019f
C839 VTAIL.n152 VSUBS 0.014185f
C840 VTAIL.n153 VSUBS 0.056689f
C841 VTAIL.n154 VSUBS 0.042144f
C842 VTAIL.n155 VSUBS 1.21094f
C843 VTAIL.n156 VSUBS 0.02979f
C844 VTAIL.n157 VSUBS 0.026397f
C845 VTAIL.n158 VSUBS 0.014185f
C846 VTAIL.n159 VSUBS 0.033528f
C847 VTAIL.n160 VSUBS 0.015019f
C848 VTAIL.n161 VSUBS 0.026397f
C849 VTAIL.n162 VSUBS 0.014185f
C850 VTAIL.n163 VSUBS 0.033528f
C851 VTAIL.n164 VSUBS 0.015019f
C852 VTAIL.n165 VSUBS 0.026397f
C853 VTAIL.n166 VSUBS 0.014185f
C854 VTAIL.n167 VSUBS 0.033528f
C855 VTAIL.n168 VSUBS 0.015019f
C856 VTAIL.n169 VSUBS 0.026397f
C857 VTAIL.n170 VSUBS 0.014185f
C858 VTAIL.n171 VSUBS 0.025146f
C859 VTAIL.n172 VSUBS 0.021329f
C860 VTAIL.t2 VSUBS 0.071477f
C861 VTAIL.n173 VSUBS 0.143162f
C862 VTAIL.n174 VSUBS 1.0239f
C863 VTAIL.n175 VSUBS 0.014185f
C864 VTAIL.n176 VSUBS 0.015019f
C865 VTAIL.n177 VSUBS 0.033528f
C866 VTAIL.n178 VSUBS 0.033528f
C867 VTAIL.n179 VSUBS 0.015019f
C868 VTAIL.n180 VSUBS 0.014185f
C869 VTAIL.n181 VSUBS 0.026397f
C870 VTAIL.n182 VSUBS 0.026397f
C871 VTAIL.n183 VSUBS 0.014185f
C872 VTAIL.n184 VSUBS 0.015019f
C873 VTAIL.n185 VSUBS 0.033528f
C874 VTAIL.n186 VSUBS 0.033528f
C875 VTAIL.n187 VSUBS 0.015019f
C876 VTAIL.n188 VSUBS 0.014185f
C877 VTAIL.n189 VSUBS 0.026397f
C878 VTAIL.n190 VSUBS 0.026397f
C879 VTAIL.n191 VSUBS 0.014185f
C880 VTAIL.n192 VSUBS 0.015019f
C881 VTAIL.n193 VSUBS 0.033528f
C882 VTAIL.n194 VSUBS 0.033528f
C883 VTAIL.n195 VSUBS 0.015019f
C884 VTAIL.n196 VSUBS 0.014185f
C885 VTAIL.n197 VSUBS 0.026397f
C886 VTAIL.n198 VSUBS 0.026397f
C887 VTAIL.n199 VSUBS 0.014185f
C888 VTAIL.n200 VSUBS 0.015019f
C889 VTAIL.n201 VSUBS 0.033528f
C890 VTAIL.n202 VSUBS 0.08384f
C891 VTAIL.n203 VSUBS 0.015019f
C892 VTAIL.n204 VSUBS 0.014185f
C893 VTAIL.n205 VSUBS 0.056689f
C894 VTAIL.n206 VSUBS 0.042144f
C895 VTAIL.n207 VSUBS 1.15008f
C896 VN.t0 VSUBS 0.582327f
C897 VN.t1 VSUBS 0.658064f
.ends

