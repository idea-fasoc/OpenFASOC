* NGSPICE file created from diff_pair_sample_0346.ext - technology: sky130A

.subckt diff_pair_sample_0346 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=2.9211 pd=15.76 as=0 ps=0 w=7.49 l=2.32
X1 VDD2.t3 VN.t0 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.23585 pd=7.82 as=2.9211 ps=15.76 w=7.49 l=2.32
X2 VTAIL.t6 VN.t1 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9211 pd=15.76 as=1.23585 ps=7.82 w=7.49 l=2.32
X3 VDD1.t3 VP.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.23585 pd=7.82 as=2.9211 ps=15.76 w=7.49 l=2.32
X4 VTAIL.t7 VN.t2 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.9211 pd=15.76 as=1.23585 ps=7.82 w=7.49 l=2.32
X5 VDD2.t0 VN.t3 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.23585 pd=7.82 as=2.9211 ps=15.76 w=7.49 l=2.32
X6 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=2.9211 pd=15.76 as=0 ps=0 w=7.49 l=2.32
X7 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.9211 pd=15.76 as=0 ps=0 w=7.49 l=2.32
X8 VTAIL.t3 VP.t1 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9211 pd=15.76 as=1.23585 ps=7.82 w=7.49 l=2.32
X9 VTAIL.t0 VP.t2 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.9211 pd=15.76 as=1.23585 ps=7.82 w=7.49 l=2.32
X10 VDD1.t0 VP.t3 VTAIL.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.23585 pd=7.82 as=2.9211 ps=15.76 w=7.49 l=2.32
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.9211 pd=15.76 as=0 ps=0 w=7.49 l=2.32
R0 B.n590 B.n589 585
R1 B.n225 B.n93 585
R2 B.n224 B.n223 585
R3 B.n222 B.n221 585
R4 B.n220 B.n219 585
R5 B.n218 B.n217 585
R6 B.n216 B.n215 585
R7 B.n214 B.n213 585
R8 B.n212 B.n211 585
R9 B.n210 B.n209 585
R10 B.n208 B.n207 585
R11 B.n206 B.n205 585
R12 B.n204 B.n203 585
R13 B.n202 B.n201 585
R14 B.n200 B.n199 585
R15 B.n198 B.n197 585
R16 B.n196 B.n195 585
R17 B.n194 B.n193 585
R18 B.n192 B.n191 585
R19 B.n190 B.n189 585
R20 B.n188 B.n187 585
R21 B.n186 B.n185 585
R22 B.n184 B.n183 585
R23 B.n182 B.n181 585
R24 B.n180 B.n179 585
R25 B.n178 B.n177 585
R26 B.n176 B.n175 585
R27 B.n174 B.n173 585
R28 B.n172 B.n171 585
R29 B.n170 B.n169 585
R30 B.n168 B.n167 585
R31 B.n166 B.n165 585
R32 B.n164 B.n163 585
R33 B.n162 B.n161 585
R34 B.n160 B.n159 585
R35 B.n158 B.n157 585
R36 B.n156 B.n155 585
R37 B.n154 B.n153 585
R38 B.n152 B.n151 585
R39 B.n150 B.n149 585
R40 B.n148 B.n147 585
R41 B.n146 B.n145 585
R42 B.n144 B.n143 585
R43 B.n142 B.n141 585
R44 B.n140 B.n139 585
R45 B.n138 B.n137 585
R46 B.n136 B.n135 585
R47 B.n134 B.n133 585
R48 B.n132 B.n131 585
R49 B.n130 B.n129 585
R50 B.n128 B.n127 585
R51 B.n126 B.n125 585
R52 B.n124 B.n123 585
R53 B.n122 B.n121 585
R54 B.n120 B.n119 585
R55 B.n118 B.n117 585
R56 B.n116 B.n115 585
R57 B.n114 B.n113 585
R58 B.n112 B.n111 585
R59 B.n110 B.n109 585
R60 B.n108 B.n107 585
R61 B.n106 B.n105 585
R62 B.n104 B.n103 585
R63 B.n102 B.n101 585
R64 B.n61 B.n60 585
R65 B.n595 B.n594 585
R66 B.n588 B.n94 585
R67 B.n94 B.n58 585
R68 B.n587 B.n57 585
R69 B.n599 B.n57 585
R70 B.n586 B.n56 585
R71 B.n600 B.n56 585
R72 B.n585 B.n55 585
R73 B.n601 B.n55 585
R74 B.n584 B.n583 585
R75 B.n583 B.n51 585
R76 B.n582 B.n50 585
R77 B.n607 B.n50 585
R78 B.n581 B.n49 585
R79 B.n608 B.n49 585
R80 B.n580 B.n48 585
R81 B.n609 B.n48 585
R82 B.n579 B.n578 585
R83 B.n578 B.n44 585
R84 B.n577 B.n43 585
R85 B.n615 B.n43 585
R86 B.n576 B.n42 585
R87 B.n616 B.n42 585
R88 B.n575 B.n41 585
R89 B.n617 B.n41 585
R90 B.n574 B.n573 585
R91 B.n573 B.n37 585
R92 B.n572 B.n36 585
R93 B.n623 B.n36 585
R94 B.n571 B.n35 585
R95 B.n624 B.n35 585
R96 B.n570 B.n34 585
R97 B.n625 B.n34 585
R98 B.n569 B.n568 585
R99 B.n568 B.n30 585
R100 B.n567 B.n29 585
R101 B.n631 B.n29 585
R102 B.n566 B.n28 585
R103 B.n632 B.n28 585
R104 B.n565 B.n27 585
R105 B.n633 B.n27 585
R106 B.n564 B.n563 585
R107 B.n563 B.n23 585
R108 B.n562 B.n22 585
R109 B.n639 B.n22 585
R110 B.n561 B.n21 585
R111 B.n640 B.n21 585
R112 B.n560 B.n20 585
R113 B.n641 B.n20 585
R114 B.n559 B.n558 585
R115 B.n558 B.n16 585
R116 B.n557 B.n15 585
R117 B.n647 B.n15 585
R118 B.n556 B.n14 585
R119 B.t2 B.n14 585
R120 B.n555 B.n13 585
R121 B.n648 B.n13 585
R122 B.n554 B.n553 585
R123 B.n553 B.n12 585
R124 B.n552 B.n551 585
R125 B.n552 B.n8 585
R126 B.n550 B.n7 585
R127 B.n655 B.n7 585
R128 B.n549 B.n6 585
R129 B.n656 B.n6 585
R130 B.n548 B.n5 585
R131 B.n657 B.n5 585
R132 B.n547 B.n546 585
R133 B.n546 B.n4 585
R134 B.n545 B.n226 585
R135 B.n545 B.n544 585
R136 B.n535 B.n227 585
R137 B.n228 B.n227 585
R138 B.n537 B.n536 585
R139 B.n538 B.n537 585
R140 B.n534 B.n232 585
R141 B.n232 B.t3 585
R142 B.n533 B.n532 585
R143 B.n532 B.n531 585
R144 B.n234 B.n233 585
R145 B.n235 B.n234 585
R146 B.n524 B.n523 585
R147 B.n525 B.n524 585
R148 B.n522 B.n240 585
R149 B.n240 B.n239 585
R150 B.n521 B.n520 585
R151 B.n520 B.n519 585
R152 B.n242 B.n241 585
R153 B.n243 B.n242 585
R154 B.n512 B.n511 585
R155 B.n513 B.n512 585
R156 B.n510 B.n247 585
R157 B.n251 B.n247 585
R158 B.n509 B.n508 585
R159 B.n508 B.n507 585
R160 B.n249 B.n248 585
R161 B.n250 B.n249 585
R162 B.n500 B.n499 585
R163 B.n501 B.n500 585
R164 B.n498 B.n256 585
R165 B.n256 B.n255 585
R166 B.n497 B.n496 585
R167 B.n496 B.n495 585
R168 B.n258 B.n257 585
R169 B.n259 B.n258 585
R170 B.n488 B.n487 585
R171 B.n489 B.n488 585
R172 B.n486 B.n264 585
R173 B.n264 B.n263 585
R174 B.n485 B.n484 585
R175 B.n484 B.n483 585
R176 B.n266 B.n265 585
R177 B.n267 B.n266 585
R178 B.n476 B.n475 585
R179 B.n477 B.n476 585
R180 B.n474 B.n272 585
R181 B.n272 B.n271 585
R182 B.n473 B.n472 585
R183 B.n472 B.n471 585
R184 B.n274 B.n273 585
R185 B.n275 B.n274 585
R186 B.n464 B.n463 585
R187 B.n465 B.n464 585
R188 B.n462 B.n280 585
R189 B.n280 B.n279 585
R190 B.n461 B.n460 585
R191 B.n460 B.n459 585
R192 B.n282 B.n281 585
R193 B.n283 B.n282 585
R194 B.n455 B.n454 585
R195 B.n286 B.n285 585
R196 B.n451 B.n450 585
R197 B.n452 B.n451 585
R198 B.n449 B.n319 585
R199 B.n448 B.n447 585
R200 B.n446 B.n445 585
R201 B.n444 B.n443 585
R202 B.n442 B.n441 585
R203 B.n440 B.n439 585
R204 B.n438 B.n437 585
R205 B.n436 B.n435 585
R206 B.n434 B.n433 585
R207 B.n432 B.n431 585
R208 B.n430 B.n429 585
R209 B.n428 B.n427 585
R210 B.n426 B.n425 585
R211 B.n424 B.n423 585
R212 B.n422 B.n421 585
R213 B.n420 B.n419 585
R214 B.n418 B.n417 585
R215 B.n416 B.n415 585
R216 B.n414 B.n413 585
R217 B.n412 B.n411 585
R218 B.n410 B.n409 585
R219 B.n408 B.n407 585
R220 B.n406 B.n405 585
R221 B.n404 B.n403 585
R222 B.n402 B.n401 585
R223 B.n399 B.n398 585
R224 B.n397 B.n396 585
R225 B.n395 B.n394 585
R226 B.n393 B.n392 585
R227 B.n391 B.n390 585
R228 B.n389 B.n388 585
R229 B.n387 B.n386 585
R230 B.n385 B.n384 585
R231 B.n383 B.n382 585
R232 B.n381 B.n380 585
R233 B.n378 B.n377 585
R234 B.n376 B.n375 585
R235 B.n374 B.n373 585
R236 B.n372 B.n371 585
R237 B.n370 B.n369 585
R238 B.n368 B.n367 585
R239 B.n366 B.n365 585
R240 B.n364 B.n363 585
R241 B.n362 B.n361 585
R242 B.n360 B.n359 585
R243 B.n358 B.n357 585
R244 B.n356 B.n355 585
R245 B.n354 B.n353 585
R246 B.n352 B.n351 585
R247 B.n350 B.n349 585
R248 B.n348 B.n347 585
R249 B.n346 B.n345 585
R250 B.n344 B.n343 585
R251 B.n342 B.n341 585
R252 B.n340 B.n339 585
R253 B.n338 B.n337 585
R254 B.n336 B.n335 585
R255 B.n334 B.n333 585
R256 B.n332 B.n331 585
R257 B.n330 B.n329 585
R258 B.n328 B.n327 585
R259 B.n326 B.n325 585
R260 B.n324 B.n318 585
R261 B.n452 B.n318 585
R262 B.n456 B.n284 585
R263 B.n284 B.n283 585
R264 B.n458 B.n457 585
R265 B.n459 B.n458 585
R266 B.n278 B.n277 585
R267 B.n279 B.n278 585
R268 B.n467 B.n466 585
R269 B.n466 B.n465 585
R270 B.n468 B.n276 585
R271 B.n276 B.n275 585
R272 B.n470 B.n469 585
R273 B.n471 B.n470 585
R274 B.n270 B.n269 585
R275 B.n271 B.n270 585
R276 B.n479 B.n478 585
R277 B.n478 B.n477 585
R278 B.n480 B.n268 585
R279 B.n268 B.n267 585
R280 B.n482 B.n481 585
R281 B.n483 B.n482 585
R282 B.n262 B.n261 585
R283 B.n263 B.n262 585
R284 B.n491 B.n490 585
R285 B.n490 B.n489 585
R286 B.n492 B.n260 585
R287 B.n260 B.n259 585
R288 B.n494 B.n493 585
R289 B.n495 B.n494 585
R290 B.n254 B.n253 585
R291 B.n255 B.n254 585
R292 B.n503 B.n502 585
R293 B.n502 B.n501 585
R294 B.n504 B.n252 585
R295 B.n252 B.n250 585
R296 B.n506 B.n505 585
R297 B.n507 B.n506 585
R298 B.n246 B.n245 585
R299 B.n251 B.n246 585
R300 B.n515 B.n514 585
R301 B.n514 B.n513 585
R302 B.n516 B.n244 585
R303 B.n244 B.n243 585
R304 B.n518 B.n517 585
R305 B.n519 B.n518 585
R306 B.n238 B.n237 585
R307 B.n239 B.n238 585
R308 B.n527 B.n526 585
R309 B.n526 B.n525 585
R310 B.n528 B.n236 585
R311 B.n236 B.n235 585
R312 B.n530 B.n529 585
R313 B.n531 B.n530 585
R314 B.n231 B.n230 585
R315 B.t3 B.n231 585
R316 B.n540 B.n539 585
R317 B.n539 B.n538 585
R318 B.n541 B.n229 585
R319 B.n229 B.n228 585
R320 B.n543 B.n542 585
R321 B.n544 B.n543 585
R322 B.n3 B.n0 585
R323 B.n4 B.n3 585
R324 B.n654 B.n1 585
R325 B.n655 B.n654 585
R326 B.n653 B.n652 585
R327 B.n653 B.n8 585
R328 B.n651 B.n9 585
R329 B.n12 B.n9 585
R330 B.n650 B.n649 585
R331 B.n649 B.n648 585
R332 B.n11 B.n10 585
R333 B.t2 B.n11 585
R334 B.n646 B.n645 585
R335 B.n647 B.n646 585
R336 B.n644 B.n17 585
R337 B.n17 B.n16 585
R338 B.n643 B.n642 585
R339 B.n642 B.n641 585
R340 B.n19 B.n18 585
R341 B.n640 B.n19 585
R342 B.n638 B.n637 585
R343 B.n639 B.n638 585
R344 B.n636 B.n24 585
R345 B.n24 B.n23 585
R346 B.n635 B.n634 585
R347 B.n634 B.n633 585
R348 B.n26 B.n25 585
R349 B.n632 B.n26 585
R350 B.n630 B.n629 585
R351 B.n631 B.n630 585
R352 B.n628 B.n31 585
R353 B.n31 B.n30 585
R354 B.n627 B.n626 585
R355 B.n626 B.n625 585
R356 B.n33 B.n32 585
R357 B.n624 B.n33 585
R358 B.n622 B.n621 585
R359 B.n623 B.n622 585
R360 B.n620 B.n38 585
R361 B.n38 B.n37 585
R362 B.n619 B.n618 585
R363 B.n618 B.n617 585
R364 B.n40 B.n39 585
R365 B.n616 B.n40 585
R366 B.n614 B.n613 585
R367 B.n615 B.n614 585
R368 B.n612 B.n45 585
R369 B.n45 B.n44 585
R370 B.n611 B.n610 585
R371 B.n610 B.n609 585
R372 B.n47 B.n46 585
R373 B.n608 B.n47 585
R374 B.n606 B.n605 585
R375 B.n607 B.n606 585
R376 B.n604 B.n52 585
R377 B.n52 B.n51 585
R378 B.n603 B.n602 585
R379 B.n602 B.n601 585
R380 B.n54 B.n53 585
R381 B.n600 B.n54 585
R382 B.n598 B.n597 585
R383 B.n599 B.n598 585
R384 B.n596 B.n59 585
R385 B.n59 B.n58 585
R386 B.n658 B.n657 585
R387 B.n656 B.n2 585
R388 B.n594 B.n59 521.33
R389 B.n590 B.n94 521.33
R390 B.n318 B.n282 521.33
R391 B.n454 B.n284 521.33
R392 B.n98 B.t8 285.387
R393 B.n95 B.t15 285.387
R394 B.n322 B.t12 285.387
R395 B.n320 B.t4 285.387
R396 B.n592 B.n591 256.663
R397 B.n592 B.n92 256.663
R398 B.n592 B.n91 256.663
R399 B.n592 B.n90 256.663
R400 B.n592 B.n89 256.663
R401 B.n592 B.n88 256.663
R402 B.n592 B.n87 256.663
R403 B.n592 B.n86 256.663
R404 B.n592 B.n85 256.663
R405 B.n592 B.n84 256.663
R406 B.n592 B.n83 256.663
R407 B.n592 B.n82 256.663
R408 B.n592 B.n81 256.663
R409 B.n592 B.n80 256.663
R410 B.n592 B.n79 256.663
R411 B.n592 B.n78 256.663
R412 B.n592 B.n77 256.663
R413 B.n592 B.n76 256.663
R414 B.n592 B.n75 256.663
R415 B.n592 B.n74 256.663
R416 B.n592 B.n73 256.663
R417 B.n592 B.n72 256.663
R418 B.n592 B.n71 256.663
R419 B.n592 B.n70 256.663
R420 B.n592 B.n69 256.663
R421 B.n592 B.n68 256.663
R422 B.n592 B.n67 256.663
R423 B.n592 B.n66 256.663
R424 B.n592 B.n65 256.663
R425 B.n592 B.n64 256.663
R426 B.n592 B.n63 256.663
R427 B.n592 B.n62 256.663
R428 B.n593 B.n592 256.663
R429 B.n453 B.n452 256.663
R430 B.n452 B.n287 256.663
R431 B.n452 B.n288 256.663
R432 B.n452 B.n289 256.663
R433 B.n452 B.n290 256.663
R434 B.n452 B.n291 256.663
R435 B.n452 B.n292 256.663
R436 B.n452 B.n293 256.663
R437 B.n452 B.n294 256.663
R438 B.n452 B.n295 256.663
R439 B.n452 B.n296 256.663
R440 B.n452 B.n297 256.663
R441 B.n452 B.n298 256.663
R442 B.n452 B.n299 256.663
R443 B.n452 B.n300 256.663
R444 B.n452 B.n301 256.663
R445 B.n452 B.n302 256.663
R446 B.n452 B.n303 256.663
R447 B.n452 B.n304 256.663
R448 B.n452 B.n305 256.663
R449 B.n452 B.n306 256.663
R450 B.n452 B.n307 256.663
R451 B.n452 B.n308 256.663
R452 B.n452 B.n309 256.663
R453 B.n452 B.n310 256.663
R454 B.n452 B.n311 256.663
R455 B.n452 B.n312 256.663
R456 B.n452 B.n313 256.663
R457 B.n452 B.n314 256.663
R458 B.n452 B.n315 256.663
R459 B.n452 B.n316 256.663
R460 B.n452 B.n317 256.663
R461 B.n660 B.n659 256.663
R462 B.n101 B.n61 163.367
R463 B.n105 B.n104 163.367
R464 B.n109 B.n108 163.367
R465 B.n113 B.n112 163.367
R466 B.n117 B.n116 163.367
R467 B.n121 B.n120 163.367
R468 B.n125 B.n124 163.367
R469 B.n129 B.n128 163.367
R470 B.n133 B.n132 163.367
R471 B.n137 B.n136 163.367
R472 B.n141 B.n140 163.367
R473 B.n145 B.n144 163.367
R474 B.n149 B.n148 163.367
R475 B.n153 B.n152 163.367
R476 B.n157 B.n156 163.367
R477 B.n161 B.n160 163.367
R478 B.n165 B.n164 163.367
R479 B.n169 B.n168 163.367
R480 B.n173 B.n172 163.367
R481 B.n177 B.n176 163.367
R482 B.n181 B.n180 163.367
R483 B.n185 B.n184 163.367
R484 B.n189 B.n188 163.367
R485 B.n193 B.n192 163.367
R486 B.n197 B.n196 163.367
R487 B.n201 B.n200 163.367
R488 B.n205 B.n204 163.367
R489 B.n209 B.n208 163.367
R490 B.n213 B.n212 163.367
R491 B.n217 B.n216 163.367
R492 B.n221 B.n220 163.367
R493 B.n223 B.n93 163.367
R494 B.n460 B.n282 163.367
R495 B.n460 B.n280 163.367
R496 B.n464 B.n280 163.367
R497 B.n464 B.n274 163.367
R498 B.n472 B.n274 163.367
R499 B.n472 B.n272 163.367
R500 B.n476 B.n272 163.367
R501 B.n476 B.n266 163.367
R502 B.n484 B.n266 163.367
R503 B.n484 B.n264 163.367
R504 B.n488 B.n264 163.367
R505 B.n488 B.n258 163.367
R506 B.n496 B.n258 163.367
R507 B.n496 B.n256 163.367
R508 B.n500 B.n256 163.367
R509 B.n500 B.n249 163.367
R510 B.n508 B.n249 163.367
R511 B.n508 B.n247 163.367
R512 B.n512 B.n247 163.367
R513 B.n512 B.n242 163.367
R514 B.n520 B.n242 163.367
R515 B.n520 B.n240 163.367
R516 B.n524 B.n240 163.367
R517 B.n524 B.n234 163.367
R518 B.n532 B.n234 163.367
R519 B.n532 B.n232 163.367
R520 B.n537 B.n232 163.367
R521 B.n537 B.n227 163.367
R522 B.n545 B.n227 163.367
R523 B.n546 B.n545 163.367
R524 B.n546 B.n5 163.367
R525 B.n6 B.n5 163.367
R526 B.n7 B.n6 163.367
R527 B.n552 B.n7 163.367
R528 B.n553 B.n552 163.367
R529 B.n553 B.n13 163.367
R530 B.n14 B.n13 163.367
R531 B.n15 B.n14 163.367
R532 B.n558 B.n15 163.367
R533 B.n558 B.n20 163.367
R534 B.n21 B.n20 163.367
R535 B.n22 B.n21 163.367
R536 B.n563 B.n22 163.367
R537 B.n563 B.n27 163.367
R538 B.n28 B.n27 163.367
R539 B.n29 B.n28 163.367
R540 B.n568 B.n29 163.367
R541 B.n568 B.n34 163.367
R542 B.n35 B.n34 163.367
R543 B.n36 B.n35 163.367
R544 B.n573 B.n36 163.367
R545 B.n573 B.n41 163.367
R546 B.n42 B.n41 163.367
R547 B.n43 B.n42 163.367
R548 B.n578 B.n43 163.367
R549 B.n578 B.n48 163.367
R550 B.n49 B.n48 163.367
R551 B.n50 B.n49 163.367
R552 B.n583 B.n50 163.367
R553 B.n583 B.n55 163.367
R554 B.n56 B.n55 163.367
R555 B.n57 B.n56 163.367
R556 B.n94 B.n57 163.367
R557 B.n451 B.n286 163.367
R558 B.n451 B.n319 163.367
R559 B.n447 B.n446 163.367
R560 B.n443 B.n442 163.367
R561 B.n439 B.n438 163.367
R562 B.n435 B.n434 163.367
R563 B.n431 B.n430 163.367
R564 B.n427 B.n426 163.367
R565 B.n423 B.n422 163.367
R566 B.n419 B.n418 163.367
R567 B.n415 B.n414 163.367
R568 B.n411 B.n410 163.367
R569 B.n407 B.n406 163.367
R570 B.n403 B.n402 163.367
R571 B.n398 B.n397 163.367
R572 B.n394 B.n393 163.367
R573 B.n390 B.n389 163.367
R574 B.n386 B.n385 163.367
R575 B.n382 B.n381 163.367
R576 B.n377 B.n376 163.367
R577 B.n373 B.n372 163.367
R578 B.n369 B.n368 163.367
R579 B.n365 B.n364 163.367
R580 B.n361 B.n360 163.367
R581 B.n357 B.n356 163.367
R582 B.n353 B.n352 163.367
R583 B.n349 B.n348 163.367
R584 B.n345 B.n344 163.367
R585 B.n341 B.n340 163.367
R586 B.n337 B.n336 163.367
R587 B.n333 B.n332 163.367
R588 B.n329 B.n328 163.367
R589 B.n325 B.n318 163.367
R590 B.n458 B.n284 163.367
R591 B.n458 B.n278 163.367
R592 B.n466 B.n278 163.367
R593 B.n466 B.n276 163.367
R594 B.n470 B.n276 163.367
R595 B.n470 B.n270 163.367
R596 B.n478 B.n270 163.367
R597 B.n478 B.n268 163.367
R598 B.n482 B.n268 163.367
R599 B.n482 B.n262 163.367
R600 B.n490 B.n262 163.367
R601 B.n490 B.n260 163.367
R602 B.n494 B.n260 163.367
R603 B.n494 B.n254 163.367
R604 B.n502 B.n254 163.367
R605 B.n502 B.n252 163.367
R606 B.n506 B.n252 163.367
R607 B.n506 B.n246 163.367
R608 B.n514 B.n246 163.367
R609 B.n514 B.n244 163.367
R610 B.n518 B.n244 163.367
R611 B.n518 B.n238 163.367
R612 B.n526 B.n238 163.367
R613 B.n526 B.n236 163.367
R614 B.n530 B.n236 163.367
R615 B.n530 B.n231 163.367
R616 B.n539 B.n231 163.367
R617 B.n539 B.n229 163.367
R618 B.n543 B.n229 163.367
R619 B.n543 B.n3 163.367
R620 B.n658 B.n3 163.367
R621 B.n654 B.n2 163.367
R622 B.n654 B.n653 163.367
R623 B.n653 B.n9 163.367
R624 B.n649 B.n9 163.367
R625 B.n649 B.n11 163.367
R626 B.n646 B.n11 163.367
R627 B.n646 B.n17 163.367
R628 B.n642 B.n17 163.367
R629 B.n642 B.n19 163.367
R630 B.n638 B.n19 163.367
R631 B.n638 B.n24 163.367
R632 B.n634 B.n24 163.367
R633 B.n634 B.n26 163.367
R634 B.n630 B.n26 163.367
R635 B.n630 B.n31 163.367
R636 B.n626 B.n31 163.367
R637 B.n626 B.n33 163.367
R638 B.n622 B.n33 163.367
R639 B.n622 B.n38 163.367
R640 B.n618 B.n38 163.367
R641 B.n618 B.n40 163.367
R642 B.n614 B.n40 163.367
R643 B.n614 B.n45 163.367
R644 B.n610 B.n45 163.367
R645 B.n610 B.n47 163.367
R646 B.n606 B.n47 163.367
R647 B.n606 B.n52 163.367
R648 B.n602 B.n52 163.367
R649 B.n602 B.n54 163.367
R650 B.n598 B.n54 163.367
R651 B.n598 B.n59 163.367
R652 B.n95 B.t16 120.367
R653 B.n322 B.t14 120.367
R654 B.n98 B.t10 120.358
R655 B.n320 B.t7 120.358
R656 B.n452 B.n283 105.993
R657 B.n592 B.n58 105.993
R658 B.n594 B.n593 71.676
R659 B.n101 B.n62 71.676
R660 B.n105 B.n63 71.676
R661 B.n109 B.n64 71.676
R662 B.n113 B.n65 71.676
R663 B.n117 B.n66 71.676
R664 B.n121 B.n67 71.676
R665 B.n125 B.n68 71.676
R666 B.n129 B.n69 71.676
R667 B.n133 B.n70 71.676
R668 B.n137 B.n71 71.676
R669 B.n141 B.n72 71.676
R670 B.n145 B.n73 71.676
R671 B.n149 B.n74 71.676
R672 B.n153 B.n75 71.676
R673 B.n157 B.n76 71.676
R674 B.n161 B.n77 71.676
R675 B.n165 B.n78 71.676
R676 B.n169 B.n79 71.676
R677 B.n173 B.n80 71.676
R678 B.n177 B.n81 71.676
R679 B.n181 B.n82 71.676
R680 B.n185 B.n83 71.676
R681 B.n189 B.n84 71.676
R682 B.n193 B.n85 71.676
R683 B.n197 B.n86 71.676
R684 B.n201 B.n87 71.676
R685 B.n205 B.n88 71.676
R686 B.n209 B.n89 71.676
R687 B.n213 B.n90 71.676
R688 B.n217 B.n91 71.676
R689 B.n221 B.n92 71.676
R690 B.n591 B.n93 71.676
R691 B.n591 B.n590 71.676
R692 B.n223 B.n92 71.676
R693 B.n220 B.n91 71.676
R694 B.n216 B.n90 71.676
R695 B.n212 B.n89 71.676
R696 B.n208 B.n88 71.676
R697 B.n204 B.n87 71.676
R698 B.n200 B.n86 71.676
R699 B.n196 B.n85 71.676
R700 B.n192 B.n84 71.676
R701 B.n188 B.n83 71.676
R702 B.n184 B.n82 71.676
R703 B.n180 B.n81 71.676
R704 B.n176 B.n80 71.676
R705 B.n172 B.n79 71.676
R706 B.n168 B.n78 71.676
R707 B.n164 B.n77 71.676
R708 B.n160 B.n76 71.676
R709 B.n156 B.n75 71.676
R710 B.n152 B.n74 71.676
R711 B.n148 B.n73 71.676
R712 B.n144 B.n72 71.676
R713 B.n140 B.n71 71.676
R714 B.n136 B.n70 71.676
R715 B.n132 B.n69 71.676
R716 B.n128 B.n68 71.676
R717 B.n124 B.n67 71.676
R718 B.n120 B.n66 71.676
R719 B.n116 B.n65 71.676
R720 B.n112 B.n64 71.676
R721 B.n108 B.n63 71.676
R722 B.n104 B.n62 71.676
R723 B.n593 B.n61 71.676
R724 B.n454 B.n453 71.676
R725 B.n319 B.n287 71.676
R726 B.n446 B.n288 71.676
R727 B.n442 B.n289 71.676
R728 B.n438 B.n290 71.676
R729 B.n434 B.n291 71.676
R730 B.n430 B.n292 71.676
R731 B.n426 B.n293 71.676
R732 B.n422 B.n294 71.676
R733 B.n418 B.n295 71.676
R734 B.n414 B.n296 71.676
R735 B.n410 B.n297 71.676
R736 B.n406 B.n298 71.676
R737 B.n402 B.n299 71.676
R738 B.n397 B.n300 71.676
R739 B.n393 B.n301 71.676
R740 B.n389 B.n302 71.676
R741 B.n385 B.n303 71.676
R742 B.n381 B.n304 71.676
R743 B.n376 B.n305 71.676
R744 B.n372 B.n306 71.676
R745 B.n368 B.n307 71.676
R746 B.n364 B.n308 71.676
R747 B.n360 B.n309 71.676
R748 B.n356 B.n310 71.676
R749 B.n352 B.n311 71.676
R750 B.n348 B.n312 71.676
R751 B.n344 B.n313 71.676
R752 B.n340 B.n314 71.676
R753 B.n336 B.n315 71.676
R754 B.n332 B.n316 71.676
R755 B.n328 B.n317 71.676
R756 B.n453 B.n286 71.676
R757 B.n447 B.n287 71.676
R758 B.n443 B.n288 71.676
R759 B.n439 B.n289 71.676
R760 B.n435 B.n290 71.676
R761 B.n431 B.n291 71.676
R762 B.n427 B.n292 71.676
R763 B.n423 B.n293 71.676
R764 B.n419 B.n294 71.676
R765 B.n415 B.n295 71.676
R766 B.n411 B.n296 71.676
R767 B.n407 B.n297 71.676
R768 B.n403 B.n298 71.676
R769 B.n398 B.n299 71.676
R770 B.n394 B.n300 71.676
R771 B.n390 B.n301 71.676
R772 B.n386 B.n302 71.676
R773 B.n382 B.n303 71.676
R774 B.n377 B.n304 71.676
R775 B.n373 B.n305 71.676
R776 B.n369 B.n306 71.676
R777 B.n365 B.n307 71.676
R778 B.n361 B.n308 71.676
R779 B.n357 B.n309 71.676
R780 B.n353 B.n310 71.676
R781 B.n349 B.n311 71.676
R782 B.n345 B.n312 71.676
R783 B.n341 B.n313 71.676
R784 B.n337 B.n314 71.676
R785 B.n333 B.n315 71.676
R786 B.n329 B.n316 71.676
R787 B.n325 B.n317 71.676
R788 B.n659 B.n658 71.676
R789 B.n659 B.n2 71.676
R790 B.n96 B.t17 68.9723
R791 B.n323 B.t13 68.9723
R792 B.n99 B.t11 68.9635
R793 B.n321 B.t6 68.9635
R794 B.n100 B.n99 59.5399
R795 B.n97 B.n96 59.5399
R796 B.n379 B.n323 59.5399
R797 B.n400 B.n321 59.5399
R798 B.n459 B.n283 58.5982
R799 B.n459 B.n279 58.5982
R800 B.n465 B.n279 58.5982
R801 B.n465 B.n275 58.5982
R802 B.n471 B.n275 58.5982
R803 B.n471 B.n271 58.5982
R804 B.n477 B.n271 58.5982
R805 B.n483 B.n267 58.5982
R806 B.n483 B.n263 58.5982
R807 B.n489 B.n263 58.5982
R808 B.n489 B.n259 58.5982
R809 B.n495 B.n259 58.5982
R810 B.n495 B.n255 58.5982
R811 B.n501 B.n255 58.5982
R812 B.n501 B.n250 58.5982
R813 B.n507 B.n250 58.5982
R814 B.n507 B.n251 58.5982
R815 B.n513 B.n243 58.5982
R816 B.n519 B.n243 58.5982
R817 B.n519 B.n239 58.5982
R818 B.n525 B.n239 58.5982
R819 B.n525 B.n235 58.5982
R820 B.n531 B.n235 58.5982
R821 B.n531 B.t3 58.5982
R822 B.n538 B.t3 58.5982
R823 B.n538 B.n228 58.5982
R824 B.n544 B.n228 58.5982
R825 B.n544 B.n4 58.5982
R826 B.n657 B.n4 58.5982
R827 B.n657 B.n656 58.5982
R828 B.n656 B.n655 58.5982
R829 B.n655 B.n8 58.5982
R830 B.n12 B.n8 58.5982
R831 B.n648 B.n12 58.5982
R832 B.n648 B.t2 58.5982
R833 B.t2 B.n647 58.5982
R834 B.n647 B.n16 58.5982
R835 B.n641 B.n16 58.5982
R836 B.n641 B.n640 58.5982
R837 B.n640 B.n639 58.5982
R838 B.n639 B.n23 58.5982
R839 B.n633 B.n23 58.5982
R840 B.n632 B.n631 58.5982
R841 B.n631 B.n30 58.5982
R842 B.n625 B.n30 58.5982
R843 B.n625 B.n624 58.5982
R844 B.n624 B.n623 58.5982
R845 B.n623 B.n37 58.5982
R846 B.n617 B.n37 58.5982
R847 B.n617 B.n616 58.5982
R848 B.n616 B.n615 58.5982
R849 B.n615 B.n44 58.5982
R850 B.n609 B.n608 58.5982
R851 B.n608 B.n607 58.5982
R852 B.n607 B.n51 58.5982
R853 B.n601 B.n51 58.5982
R854 B.n601 B.n600 58.5982
R855 B.n600 B.n599 58.5982
R856 B.n599 B.n58 58.5982
R857 B.n99 B.n98 51.3944
R858 B.n96 B.n95 51.3944
R859 B.n323 B.n322 51.3944
R860 B.n321 B.n320 51.3944
R861 B.t5 B.n267 46.534
R862 B.n513 B.t1 46.534
R863 B.n633 B.t0 46.534
R864 B.t9 B.n44 46.534
R865 B.n456 B.n455 33.8737
R866 B.n324 B.n281 33.8737
R867 B.n589 B.n588 33.8737
R868 B.n596 B.n595 33.8737
R869 B B.n660 18.0485
R870 B.n477 B.t5 12.0647
R871 B.n251 B.t1 12.0647
R872 B.t0 B.n632 12.0647
R873 B.n609 B.t9 12.0647
R874 B.n457 B.n456 10.6151
R875 B.n457 B.n277 10.6151
R876 B.n467 B.n277 10.6151
R877 B.n468 B.n467 10.6151
R878 B.n469 B.n468 10.6151
R879 B.n469 B.n269 10.6151
R880 B.n479 B.n269 10.6151
R881 B.n480 B.n479 10.6151
R882 B.n481 B.n480 10.6151
R883 B.n481 B.n261 10.6151
R884 B.n491 B.n261 10.6151
R885 B.n492 B.n491 10.6151
R886 B.n493 B.n492 10.6151
R887 B.n493 B.n253 10.6151
R888 B.n503 B.n253 10.6151
R889 B.n504 B.n503 10.6151
R890 B.n505 B.n504 10.6151
R891 B.n505 B.n245 10.6151
R892 B.n515 B.n245 10.6151
R893 B.n516 B.n515 10.6151
R894 B.n517 B.n516 10.6151
R895 B.n517 B.n237 10.6151
R896 B.n527 B.n237 10.6151
R897 B.n528 B.n527 10.6151
R898 B.n529 B.n528 10.6151
R899 B.n529 B.n230 10.6151
R900 B.n540 B.n230 10.6151
R901 B.n541 B.n540 10.6151
R902 B.n542 B.n541 10.6151
R903 B.n542 B.n0 10.6151
R904 B.n455 B.n285 10.6151
R905 B.n450 B.n285 10.6151
R906 B.n450 B.n449 10.6151
R907 B.n449 B.n448 10.6151
R908 B.n448 B.n445 10.6151
R909 B.n445 B.n444 10.6151
R910 B.n444 B.n441 10.6151
R911 B.n441 B.n440 10.6151
R912 B.n440 B.n437 10.6151
R913 B.n437 B.n436 10.6151
R914 B.n436 B.n433 10.6151
R915 B.n433 B.n432 10.6151
R916 B.n432 B.n429 10.6151
R917 B.n429 B.n428 10.6151
R918 B.n428 B.n425 10.6151
R919 B.n425 B.n424 10.6151
R920 B.n424 B.n421 10.6151
R921 B.n421 B.n420 10.6151
R922 B.n420 B.n417 10.6151
R923 B.n417 B.n416 10.6151
R924 B.n416 B.n413 10.6151
R925 B.n413 B.n412 10.6151
R926 B.n412 B.n409 10.6151
R927 B.n409 B.n408 10.6151
R928 B.n408 B.n405 10.6151
R929 B.n405 B.n404 10.6151
R930 B.n404 B.n401 10.6151
R931 B.n399 B.n396 10.6151
R932 B.n396 B.n395 10.6151
R933 B.n395 B.n392 10.6151
R934 B.n392 B.n391 10.6151
R935 B.n391 B.n388 10.6151
R936 B.n388 B.n387 10.6151
R937 B.n387 B.n384 10.6151
R938 B.n384 B.n383 10.6151
R939 B.n383 B.n380 10.6151
R940 B.n378 B.n375 10.6151
R941 B.n375 B.n374 10.6151
R942 B.n374 B.n371 10.6151
R943 B.n371 B.n370 10.6151
R944 B.n370 B.n367 10.6151
R945 B.n367 B.n366 10.6151
R946 B.n366 B.n363 10.6151
R947 B.n363 B.n362 10.6151
R948 B.n362 B.n359 10.6151
R949 B.n359 B.n358 10.6151
R950 B.n358 B.n355 10.6151
R951 B.n355 B.n354 10.6151
R952 B.n354 B.n351 10.6151
R953 B.n351 B.n350 10.6151
R954 B.n350 B.n347 10.6151
R955 B.n347 B.n346 10.6151
R956 B.n346 B.n343 10.6151
R957 B.n343 B.n342 10.6151
R958 B.n342 B.n339 10.6151
R959 B.n339 B.n338 10.6151
R960 B.n338 B.n335 10.6151
R961 B.n335 B.n334 10.6151
R962 B.n334 B.n331 10.6151
R963 B.n331 B.n330 10.6151
R964 B.n330 B.n327 10.6151
R965 B.n327 B.n326 10.6151
R966 B.n326 B.n324 10.6151
R967 B.n461 B.n281 10.6151
R968 B.n462 B.n461 10.6151
R969 B.n463 B.n462 10.6151
R970 B.n463 B.n273 10.6151
R971 B.n473 B.n273 10.6151
R972 B.n474 B.n473 10.6151
R973 B.n475 B.n474 10.6151
R974 B.n475 B.n265 10.6151
R975 B.n485 B.n265 10.6151
R976 B.n486 B.n485 10.6151
R977 B.n487 B.n486 10.6151
R978 B.n487 B.n257 10.6151
R979 B.n497 B.n257 10.6151
R980 B.n498 B.n497 10.6151
R981 B.n499 B.n498 10.6151
R982 B.n499 B.n248 10.6151
R983 B.n509 B.n248 10.6151
R984 B.n510 B.n509 10.6151
R985 B.n511 B.n510 10.6151
R986 B.n511 B.n241 10.6151
R987 B.n521 B.n241 10.6151
R988 B.n522 B.n521 10.6151
R989 B.n523 B.n522 10.6151
R990 B.n523 B.n233 10.6151
R991 B.n533 B.n233 10.6151
R992 B.n534 B.n533 10.6151
R993 B.n536 B.n534 10.6151
R994 B.n536 B.n535 10.6151
R995 B.n535 B.n226 10.6151
R996 B.n547 B.n226 10.6151
R997 B.n548 B.n547 10.6151
R998 B.n549 B.n548 10.6151
R999 B.n550 B.n549 10.6151
R1000 B.n551 B.n550 10.6151
R1001 B.n554 B.n551 10.6151
R1002 B.n555 B.n554 10.6151
R1003 B.n556 B.n555 10.6151
R1004 B.n557 B.n556 10.6151
R1005 B.n559 B.n557 10.6151
R1006 B.n560 B.n559 10.6151
R1007 B.n561 B.n560 10.6151
R1008 B.n562 B.n561 10.6151
R1009 B.n564 B.n562 10.6151
R1010 B.n565 B.n564 10.6151
R1011 B.n566 B.n565 10.6151
R1012 B.n567 B.n566 10.6151
R1013 B.n569 B.n567 10.6151
R1014 B.n570 B.n569 10.6151
R1015 B.n571 B.n570 10.6151
R1016 B.n572 B.n571 10.6151
R1017 B.n574 B.n572 10.6151
R1018 B.n575 B.n574 10.6151
R1019 B.n576 B.n575 10.6151
R1020 B.n577 B.n576 10.6151
R1021 B.n579 B.n577 10.6151
R1022 B.n580 B.n579 10.6151
R1023 B.n581 B.n580 10.6151
R1024 B.n582 B.n581 10.6151
R1025 B.n584 B.n582 10.6151
R1026 B.n585 B.n584 10.6151
R1027 B.n586 B.n585 10.6151
R1028 B.n587 B.n586 10.6151
R1029 B.n588 B.n587 10.6151
R1030 B.n652 B.n1 10.6151
R1031 B.n652 B.n651 10.6151
R1032 B.n651 B.n650 10.6151
R1033 B.n650 B.n10 10.6151
R1034 B.n645 B.n10 10.6151
R1035 B.n645 B.n644 10.6151
R1036 B.n644 B.n643 10.6151
R1037 B.n643 B.n18 10.6151
R1038 B.n637 B.n18 10.6151
R1039 B.n637 B.n636 10.6151
R1040 B.n636 B.n635 10.6151
R1041 B.n635 B.n25 10.6151
R1042 B.n629 B.n25 10.6151
R1043 B.n629 B.n628 10.6151
R1044 B.n628 B.n627 10.6151
R1045 B.n627 B.n32 10.6151
R1046 B.n621 B.n32 10.6151
R1047 B.n621 B.n620 10.6151
R1048 B.n620 B.n619 10.6151
R1049 B.n619 B.n39 10.6151
R1050 B.n613 B.n39 10.6151
R1051 B.n613 B.n612 10.6151
R1052 B.n612 B.n611 10.6151
R1053 B.n611 B.n46 10.6151
R1054 B.n605 B.n46 10.6151
R1055 B.n605 B.n604 10.6151
R1056 B.n604 B.n603 10.6151
R1057 B.n603 B.n53 10.6151
R1058 B.n597 B.n53 10.6151
R1059 B.n597 B.n596 10.6151
R1060 B.n595 B.n60 10.6151
R1061 B.n102 B.n60 10.6151
R1062 B.n103 B.n102 10.6151
R1063 B.n106 B.n103 10.6151
R1064 B.n107 B.n106 10.6151
R1065 B.n110 B.n107 10.6151
R1066 B.n111 B.n110 10.6151
R1067 B.n114 B.n111 10.6151
R1068 B.n115 B.n114 10.6151
R1069 B.n118 B.n115 10.6151
R1070 B.n119 B.n118 10.6151
R1071 B.n122 B.n119 10.6151
R1072 B.n123 B.n122 10.6151
R1073 B.n126 B.n123 10.6151
R1074 B.n127 B.n126 10.6151
R1075 B.n130 B.n127 10.6151
R1076 B.n131 B.n130 10.6151
R1077 B.n134 B.n131 10.6151
R1078 B.n135 B.n134 10.6151
R1079 B.n138 B.n135 10.6151
R1080 B.n139 B.n138 10.6151
R1081 B.n142 B.n139 10.6151
R1082 B.n143 B.n142 10.6151
R1083 B.n146 B.n143 10.6151
R1084 B.n147 B.n146 10.6151
R1085 B.n150 B.n147 10.6151
R1086 B.n151 B.n150 10.6151
R1087 B.n155 B.n154 10.6151
R1088 B.n158 B.n155 10.6151
R1089 B.n159 B.n158 10.6151
R1090 B.n162 B.n159 10.6151
R1091 B.n163 B.n162 10.6151
R1092 B.n166 B.n163 10.6151
R1093 B.n167 B.n166 10.6151
R1094 B.n170 B.n167 10.6151
R1095 B.n171 B.n170 10.6151
R1096 B.n175 B.n174 10.6151
R1097 B.n178 B.n175 10.6151
R1098 B.n179 B.n178 10.6151
R1099 B.n182 B.n179 10.6151
R1100 B.n183 B.n182 10.6151
R1101 B.n186 B.n183 10.6151
R1102 B.n187 B.n186 10.6151
R1103 B.n190 B.n187 10.6151
R1104 B.n191 B.n190 10.6151
R1105 B.n194 B.n191 10.6151
R1106 B.n195 B.n194 10.6151
R1107 B.n198 B.n195 10.6151
R1108 B.n199 B.n198 10.6151
R1109 B.n202 B.n199 10.6151
R1110 B.n203 B.n202 10.6151
R1111 B.n206 B.n203 10.6151
R1112 B.n207 B.n206 10.6151
R1113 B.n210 B.n207 10.6151
R1114 B.n211 B.n210 10.6151
R1115 B.n214 B.n211 10.6151
R1116 B.n215 B.n214 10.6151
R1117 B.n218 B.n215 10.6151
R1118 B.n219 B.n218 10.6151
R1119 B.n222 B.n219 10.6151
R1120 B.n224 B.n222 10.6151
R1121 B.n225 B.n224 10.6151
R1122 B.n589 B.n225 10.6151
R1123 B.n401 B.n400 9.36635
R1124 B.n379 B.n378 9.36635
R1125 B.n151 B.n100 9.36635
R1126 B.n174 B.n97 9.36635
R1127 B.n660 B.n0 8.11757
R1128 B.n660 B.n1 8.11757
R1129 B.n400 B.n399 1.24928
R1130 B.n380 B.n379 1.24928
R1131 B.n154 B.n100 1.24928
R1132 B.n171 B.n97 1.24928
R1133 VN.n0 VN.t2 114.272
R1134 VN.n1 VN.t3 114.272
R1135 VN.n0 VN.t0 113.615
R1136 VN.n1 VN.t1 113.615
R1137 VN VN.n1 47.8362
R1138 VN VN.n0 5.51418
R1139 VTAIL.n5 VTAIL.t0 51.2257
R1140 VTAIL.n4 VTAIL.t5 51.2257
R1141 VTAIL.n3 VTAIL.t6 51.2257
R1142 VTAIL.n7 VTAIL.t4 51.2255
R1143 VTAIL.n0 VTAIL.t7 51.2255
R1144 VTAIL.n1 VTAIL.t1 51.2255
R1145 VTAIL.n2 VTAIL.t3 51.2255
R1146 VTAIL.n6 VTAIL.t2 51.2255
R1147 VTAIL.n7 VTAIL.n6 21.1083
R1148 VTAIL.n3 VTAIL.n2 21.1083
R1149 VTAIL.n4 VTAIL.n3 2.28498
R1150 VTAIL.n6 VTAIL.n5 2.28498
R1151 VTAIL.n2 VTAIL.n1 2.28498
R1152 VTAIL VTAIL.n0 1.20093
R1153 VTAIL VTAIL.n7 1.08455
R1154 VTAIL.n5 VTAIL.n4 0.470328
R1155 VTAIL.n1 VTAIL.n0 0.470328
R1156 VDD2.n2 VDD2.n0 102.285
R1157 VDD2.n2 VDD2.n1 65.2608
R1158 VDD2.n1 VDD2.t2 2.64402
R1159 VDD2.n1 VDD2.t0 2.64402
R1160 VDD2.n0 VDD2.t1 2.64402
R1161 VDD2.n0 VDD2.t3 2.64402
R1162 VDD2 VDD2.n2 0.0586897
R1163 VP.n12 VP.n0 161.3
R1164 VP.n11 VP.n10 161.3
R1165 VP.n9 VP.n1 161.3
R1166 VP.n8 VP.n7 161.3
R1167 VP.n6 VP.n2 161.3
R1168 VP.n3 VP.t2 114.272
R1169 VP.n3 VP.t0 113.615
R1170 VP.n5 VP.n4 94.8529
R1171 VP.n14 VP.n13 94.8529
R1172 VP.n5 VP.t1 77.8061
R1173 VP.n13 VP.t3 77.8061
R1174 VP.n4 VP.n3 47.5573
R1175 VP.n7 VP.n1 40.4934
R1176 VP.n11 VP.n1 40.4934
R1177 VP.n7 VP.n6 24.4675
R1178 VP.n12 VP.n11 24.4675
R1179 VP.n6 VP.n5 15.9041
R1180 VP.n13 VP.n12 15.9041
R1181 VP.n4 VP.n2 0.278367
R1182 VP.n14 VP.n0 0.278367
R1183 VP.n8 VP.n2 0.189894
R1184 VP.n9 VP.n8 0.189894
R1185 VP.n10 VP.n9 0.189894
R1186 VP.n10 VP.n0 0.189894
R1187 VP VP.n14 0.153454
R1188 VDD1 VDD1.n1 102.811
R1189 VDD1 VDD1.n0 65.319
R1190 VDD1.n0 VDD1.t1 2.64402
R1191 VDD1.n0 VDD1.t3 2.64402
R1192 VDD1.n1 VDD1.t2 2.64402
R1193 VDD1.n1 VDD1.t0 2.64402
C0 VDD2 VDD1 0.962074f
C1 VTAIL VDD2 4.30657f
C2 VP VDD1 3.24949f
C3 VTAIL VP 3.09858f
C4 VDD2 VN 3.02242f
C5 VTAIL VDD1 4.254241f
C6 VP VN 5.15314f
C7 VN VDD1 0.148577f
C8 VP VDD2 0.376318f
C9 VTAIL VN 3.08447f
C10 VDD2 B 3.249892f
C11 VDD1 B 6.83238f
C12 VTAIL B 7.223039f
C13 VN B 9.81551f
C14 VP B 8.038644f
C15 VDD1.t1 B 0.162505f
C16 VDD1.t3 B 0.162505f
C17 VDD1.n0 B 1.39929f
C18 VDD1.t2 B 0.162505f
C19 VDD1.t0 B 0.162505f
C20 VDD1.n1 B 1.92279f
C21 VP.n0 B 0.039237f
C22 VP.t3 B 1.3848f
C23 VP.n1 B 0.024059f
C24 VP.n2 B 0.039237f
C25 VP.t1 B 1.3848f
C26 VP.t0 B 1.60058f
C27 VP.t2 B 1.60444f
C28 VP.n3 B 2.36286f
C29 VP.n4 B 1.4637f
C30 VP.n5 B 0.608895f
C31 VP.n6 B 0.045881f
C32 VP.n7 B 0.05915f
C33 VP.n8 B 0.029761f
C34 VP.n9 B 0.029761f
C35 VP.n10 B 0.029761f
C36 VP.n11 B 0.05915f
C37 VP.n12 B 0.045881f
C38 VP.n13 B 0.608895f
C39 VP.n14 B 0.041338f
C40 VDD2.t1 B 0.160339f
C41 VDD2.t3 B 0.160339f
C42 VDD2.n0 B 1.87282f
C43 VDD2.t2 B 0.160339f
C44 VDD2.t0 B 0.160339f
C45 VDD2.n1 B 1.38026f
C46 VDD2.n2 B 3.20032f
C47 VTAIL.t7 B 1.1071f
C48 VTAIL.n0 B 0.317324f
C49 VTAIL.t1 B 1.1071f
C50 VTAIL.n1 B 0.380284f
C51 VTAIL.t3 B 1.1071f
C52 VTAIL.n2 B 1.10552f
C53 VTAIL.t6 B 1.1071f
C54 VTAIL.n3 B 1.10552f
C55 VTAIL.t5 B 1.1071f
C56 VTAIL.n4 B 0.380282f
C57 VTAIL.t0 B 1.1071f
C58 VTAIL.n5 B 0.380282f
C59 VTAIL.t2 B 1.1071f
C60 VTAIL.n6 B 1.10552f
C61 VTAIL.t4 B 1.1071f
C62 VTAIL.n7 B 1.0358f
C63 VN.t2 B 1.57083f
C64 VN.t0 B 1.56705f
C65 VN.n0 B 1.0151f
C66 VN.t3 B 1.57083f
C67 VN.t1 B 1.56705f
C68 VN.n1 B 2.32863f
.ends

