* NGSPICE file created from diff_pair_sample_0882.ext - technology: sky130A

.subckt diff_pair_sample_0882 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=1.5717 pd=8.84 as=0 ps=0 w=4.03 l=3.9
X1 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=1.5717 pd=8.84 as=0 ps=0 w=4.03 l=3.9
X2 VTAIL.t18 VP.t0 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.66495 pd=4.36 as=0.66495 ps=4.36 w=4.03 l=3.9
X3 VTAIL.t17 VP.t1 VDD1.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=0.66495 pd=4.36 as=0.66495 ps=4.36 w=4.03 l=3.9
X4 VDD2.t9 VN.t0 VTAIL.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=0.66495 pd=4.36 as=0.66495 ps=4.36 w=4.03 l=3.9
X5 VDD2.t8 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.5717 pd=8.84 as=0.66495 ps=4.36 w=4.03 l=3.9
X6 VTAIL.t8 VN.t2 VDD2.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=0.66495 pd=4.36 as=0.66495 ps=4.36 w=4.03 l=3.9
X7 VTAIL.t7 VN.t3 VDD2.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=0.66495 pd=4.36 as=0.66495 ps=4.36 w=4.03 l=3.9
X8 VTAIL.t16 VP.t2 VDD1.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=0.66495 pd=4.36 as=0.66495 ps=4.36 w=4.03 l=3.9
X9 VTAIL.t19 VN.t4 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.66495 pd=4.36 as=0.66495 ps=4.36 w=4.03 l=3.9
X10 VTAIL.t2 VN.t5 VDD2.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.66495 pd=4.36 as=0.66495 ps=4.36 w=4.03 l=3.9
X11 VDD1.t6 VP.t3 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=1.5717 pd=8.84 as=0.66495 ps=4.36 w=4.03 l=3.9
X12 VDD2.t3 VN.t6 VTAIL.t4 B.t8 sky130_fd_pr__nfet_01v8 ad=0.66495 pd=4.36 as=1.5717 ps=8.84 w=4.03 l=3.9
X13 VDD1.t5 VP.t4 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=1.5717 pd=8.84 as=0.66495 ps=4.36 w=4.03 l=3.9
X14 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=1.5717 pd=8.84 as=0 ps=0 w=4.03 l=3.9
X15 VDD2.t2 VN.t7 VTAIL.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=0.66495 pd=4.36 as=1.5717 ps=8.84 w=4.03 l=3.9
X16 VDD1.t1 VP.t5 VTAIL.t13 B.t6 sky130_fd_pr__nfet_01v8 ad=0.66495 pd=4.36 as=0.66495 ps=4.36 w=4.03 l=3.9
X17 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.5717 pd=8.84 as=0 ps=0 w=4.03 l=3.9
X18 VDD1.t7 VP.t6 VTAIL.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=0.66495 pd=4.36 as=0.66495 ps=4.36 w=4.03 l=3.9
X19 VDD1.t2 VP.t7 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=0.66495 pd=4.36 as=1.5717 ps=8.84 w=4.03 l=3.9
X20 VDD2.t1 VN.t8 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.66495 pd=4.36 as=0.66495 ps=4.36 w=4.03 l=3.9
X21 VDD1.t4 VP.t8 VTAIL.t10 B.t8 sky130_fd_pr__nfet_01v8 ad=0.66495 pd=4.36 as=1.5717 ps=8.84 w=4.03 l=3.9
X22 VDD2.t0 VN.t9 VTAIL.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=1.5717 pd=8.84 as=0.66495 ps=4.36 w=4.03 l=3.9
X23 VTAIL.t9 VP.t9 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.66495 pd=4.36 as=0.66495 ps=4.36 w=4.03 l=3.9
R0 B.n814 B.n813 585
R1 B.n815 B.n178 585
R2 B.n817 B.n816 585
R3 B.n819 B.n177 585
R4 B.n822 B.n821 585
R5 B.n823 B.n176 585
R6 B.n825 B.n824 585
R7 B.n827 B.n175 585
R8 B.n830 B.n829 585
R9 B.n831 B.n174 585
R10 B.n833 B.n832 585
R11 B.n835 B.n173 585
R12 B.n838 B.n837 585
R13 B.n839 B.n172 585
R14 B.n841 B.n840 585
R15 B.n843 B.n171 585
R16 B.n845 B.n844 585
R17 B.n847 B.n846 585
R18 B.n850 B.n849 585
R19 B.n851 B.n166 585
R20 B.n853 B.n852 585
R21 B.n855 B.n165 585
R22 B.n858 B.n857 585
R23 B.n859 B.n164 585
R24 B.n861 B.n860 585
R25 B.n863 B.n163 585
R26 B.n865 B.n864 585
R27 B.n867 B.n866 585
R28 B.n870 B.n869 585
R29 B.n871 B.n158 585
R30 B.n873 B.n872 585
R31 B.n875 B.n157 585
R32 B.n878 B.n877 585
R33 B.n879 B.n156 585
R34 B.n881 B.n880 585
R35 B.n883 B.n155 585
R36 B.n886 B.n885 585
R37 B.n887 B.n154 585
R38 B.n889 B.n888 585
R39 B.n891 B.n153 585
R40 B.n894 B.n893 585
R41 B.n895 B.n152 585
R42 B.n897 B.n896 585
R43 B.n899 B.n151 585
R44 B.n902 B.n901 585
R45 B.n903 B.n150 585
R46 B.n811 B.n148 585
R47 B.n906 B.n148 585
R48 B.n810 B.n147 585
R49 B.n907 B.n147 585
R50 B.n809 B.n146 585
R51 B.n908 B.n146 585
R52 B.n808 B.n807 585
R53 B.n807 B.n142 585
R54 B.n806 B.n141 585
R55 B.n914 B.n141 585
R56 B.n805 B.n140 585
R57 B.n915 B.n140 585
R58 B.n804 B.n139 585
R59 B.n916 B.n139 585
R60 B.n803 B.n802 585
R61 B.n802 B.n135 585
R62 B.n801 B.n134 585
R63 B.n922 B.n134 585
R64 B.n800 B.n133 585
R65 B.n923 B.n133 585
R66 B.n799 B.n132 585
R67 B.n924 B.n132 585
R68 B.n798 B.n797 585
R69 B.n797 B.n128 585
R70 B.n796 B.n127 585
R71 B.n930 B.n127 585
R72 B.n795 B.n126 585
R73 B.n931 B.n126 585
R74 B.n794 B.n125 585
R75 B.n932 B.n125 585
R76 B.n793 B.n792 585
R77 B.n792 B.n121 585
R78 B.n791 B.n120 585
R79 B.n938 B.n120 585
R80 B.n790 B.n119 585
R81 B.n939 B.n119 585
R82 B.n789 B.n118 585
R83 B.n940 B.n118 585
R84 B.n788 B.n787 585
R85 B.n787 B.n114 585
R86 B.n786 B.n113 585
R87 B.n946 B.n113 585
R88 B.n785 B.n112 585
R89 B.n947 B.n112 585
R90 B.n784 B.n111 585
R91 B.n948 B.n111 585
R92 B.n783 B.n782 585
R93 B.n782 B.n107 585
R94 B.n781 B.n106 585
R95 B.n954 B.n106 585
R96 B.n780 B.n105 585
R97 B.n955 B.n105 585
R98 B.n779 B.n104 585
R99 B.n956 B.n104 585
R100 B.n778 B.n777 585
R101 B.n777 B.n100 585
R102 B.n776 B.n99 585
R103 B.n962 B.n99 585
R104 B.n775 B.n98 585
R105 B.n963 B.n98 585
R106 B.n774 B.n97 585
R107 B.n964 B.n97 585
R108 B.n773 B.n772 585
R109 B.n772 B.n93 585
R110 B.n771 B.n92 585
R111 B.n970 B.n92 585
R112 B.n770 B.n91 585
R113 B.n971 B.n91 585
R114 B.n769 B.n90 585
R115 B.n972 B.n90 585
R116 B.n768 B.n767 585
R117 B.n767 B.n86 585
R118 B.n766 B.n85 585
R119 B.n978 B.n85 585
R120 B.n765 B.n84 585
R121 B.n979 B.n84 585
R122 B.n764 B.n83 585
R123 B.n980 B.n83 585
R124 B.n763 B.n762 585
R125 B.n762 B.n79 585
R126 B.n761 B.n78 585
R127 B.n986 B.n78 585
R128 B.n760 B.n77 585
R129 B.n987 B.n77 585
R130 B.n759 B.n76 585
R131 B.n988 B.n76 585
R132 B.n758 B.n757 585
R133 B.n757 B.n72 585
R134 B.n756 B.n71 585
R135 B.n994 B.n71 585
R136 B.n755 B.n70 585
R137 B.n995 B.n70 585
R138 B.n754 B.n69 585
R139 B.n996 B.n69 585
R140 B.n753 B.n752 585
R141 B.n752 B.n65 585
R142 B.n751 B.n64 585
R143 B.n1002 B.n64 585
R144 B.n750 B.n63 585
R145 B.n1003 B.n63 585
R146 B.n749 B.n62 585
R147 B.n1004 B.n62 585
R148 B.n748 B.n747 585
R149 B.n747 B.n58 585
R150 B.n746 B.n57 585
R151 B.n1010 B.n57 585
R152 B.n745 B.n56 585
R153 B.n1011 B.n56 585
R154 B.n744 B.n55 585
R155 B.n1012 B.n55 585
R156 B.n743 B.n742 585
R157 B.n742 B.n51 585
R158 B.n741 B.n50 585
R159 B.n1018 B.n50 585
R160 B.n740 B.n49 585
R161 B.n1019 B.n49 585
R162 B.n739 B.n48 585
R163 B.n1020 B.n48 585
R164 B.n738 B.n737 585
R165 B.n737 B.n44 585
R166 B.n736 B.n43 585
R167 B.n1026 B.n43 585
R168 B.n735 B.n42 585
R169 B.n1027 B.n42 585
R170 B.n734 B.n41 585
R171 B.n1028 B.n41 585
R172 B.n733 B.n732 585
R173 B.n732 B.n37 585
R174 B.n731 B.n36 585
R175 B.n1034 B.n36 585
R176 B.n730 B.n35 585
R177 B.n1035 B.n35 585
R178 B.n729 B.n34 585
R179 B.n1036 B.n34 585
R180 B.n728 B.n727 585
R181 B.n727 B.n30 585
R182 B.n726 B.n29 585
R183 B.n1042 B.n29 585
R184 B.n725 B.n28 585
R185 B.n1043 B.n28 585
R186 B.n724 B.n27 585
R187 B.n1044 B.n27 585
R188 B.n723 B.n722 585
R189 B.n722 B.n23 585
R190 B.n721 B.n22 585
R191 B.n1050 B.n22 585
R192 B.n720 B.n21 585
R193 B.n1051 B.n21 585
R194 B.n719 B.n20 585
R195 B.n1052 B.n20 585
R196 B.n718 B.n717 585
R197 B.n717 B.n16 585
R198 B.n716 B.n15 585
R199 B.n1058 B.n15 585
R200 B.n715 B.n14 585
R201 B.n1059 B.n14 585
R202 B.n714 B.n13 585
R203 B.n1060 B.n13 585
R204 B.n713 B.n712 585
R205 B.n712 B.n12 585
R206 B.n711 B.n710 585
R207 B.n711 B.n8 585
R208 B.n709 B.n7 585
R209 B.n1067 B.n7 585
R210 B.n708 B.n6 585
R211 B.n1068 B.n6 585
R212 B.n707 B.n5 585
R213 B.n1069 B.n5 585
R214 B.n706 B.n705 585
R215 B.n705 B.n4 585
R216 B.n704 B.n179 585
R217 B.n704 B.n703 585
R218 B.n694 B.n180 585
R219 B.n181 B.n180 585
R220 B.n696 B.n695 585
R221 B.n697 B.n696 585
R222 B.n693 B.n186 585
R223 B.n186 B.n185 585
R224 B.n692 B.n691 585
R225 B.n691 B.n690 585
R226 B.n188 B.n187 585
R227 B.n189 B.n188 585
R228 B.n683 B.n682 585
R229 B.n684 B.n683 585
R230 B.n681 B.n194 585
R231 B.n194 B.n193 585
R232 B.n680 B.n679 585
R233 B.n679 B.n678 585
R234 B.n196 B.n195 585
R235 B.n197 B.n196 585
R236 B.n671 B.n670 585
R237 B.n672 B.n671 585
R238 B.n669 B.n202 585
R239 B.n202 B.n201 585
R240 B.n668 B.n667 585
R241 B.n667 B.n666 585
R242 B.n204 B.n203 585
R243 B.n205 B.n204 585
R244 B.n659 B.n658 585
R245 B.n660 B.n659 585
R246 B.n657 B.n210 585
R247 B.n210 B.n209 585
R248 B.n656 B.n655 585
R249 B.n655 B.n654 585
R250 B.n212 B.n211 585
R251 B.n213 B.n212 585
R252 B.n647 B.n646 585
R253 B.n648 B.n647 585
R254 B.n645 B.n218 585
R255 B.n218 B.n217 585
R256 B.n644 B.n643 585
R257 B.n643 B.n642 585
R258 B.n220 B.n219 585
R259 B.n221 B.n220 585
R260 B.n635 B.n634 585
R261 B.n636 B.n635 585
R262 B.n633 B.n226 585
R263 B.n226 B.n225 585
R264 B.n632 B.n631 585
R265 B.n631 B.n630 585
R266 B.n228 B.n227 585
R267 B.n229 B.n228 585
R268 B.n623 B.n622 585
R269 B.n624 B.n623 585
R270 B.n621 B.n234 585
R271 B.n234 B.n233 585
R272 B.n620 B.n619 585
R273 B.n619 B.n618 585
R274 B.n236 B.n235 585
R275 B.n237 B.n236 585
R276 B.n611 B.n610 585
R277 B.n612 B.n611 585
R278 B.n609 B.n241 585
R279 B.n245 B.n241 585
R280 B.n608 B.n607 585
R281 B.n607 B.n606 585
R282 B.n243 B.n242 585
R283 B.n244 B.n243 585
R284 B.n599 B.n598 585
R285 B.n600 B.n599 585
R286 B.n597 B.n250 585
R287 B.n250 B.n249 585
R288 B.n596 B.n595 585
R289 B.n595 B.n594 585
R290 B.n252 B.n251 585
R291 B.n253 B.n252 585
R292 B.n587 B.n586 585
R293 B.n588 B.n587 585
R294 B.n585 B.n258 585
R295 B.n258 B.n257 585
R296 B.n584 B.n583 585
R297 B.n583 B.n582 585
R298 B.n260 B.n259 585
R299 B.n261 B.n260 585
R300 B.n575 B.n574 585
R301 B.n576 B.n575 585
R302 B.n573 B.n265 585
R303 B.n269 B.n265 585
R304 B.n572 B.n571 585
R305 B.n571 B.n570 585
R306 B.n267 B.n266 585
R307 B.n268 B.n267 585
R308 B.n563 B.n562 585
R309 B.n564 B.n563 585
R310 B.n561 B.n274 585
R311 B.n274 B.n273 585
R312 B.n560 B.n559 585
R313 B.n559 B.n558 585
R314 B.n276 B.n275 585
R315 B.n277 B.n276 585
R316 B.n551 B.n550 585
R317 B.n552 B.n551 585
R318 B.n549 B.n282 585
R319 B.n282 B.n281 585
R320 B.n548 B.n547 585
R321 B.n547 B.n546 585
R322 B.n284 B.n283 585
R323 B.n285 B.n284 585
R324 B.n539 B.n538 585
R325 B.n540 B.n539 585
R326 B.n537 B.n290 585
R327 B.n290 B.n289 585
R328 B.n536 B.n535 585
R329 B.n535 B.n534 585
R330 B.n292 B.n291 585
R331 B.n293 B.n292 585
R332 B.n527 B.n526 585
R333 B.n528 B.n527 585
R334 B.n525 B.n298 585
R335 B.n298 B.n297 585
R336 B.n524 B.n523 585
R337 B.n523 B.n522 585
R338 B.n300 B.n299 585
R339 B.n301 B.n300 585
R340 B.n515 B.n514 585
R341 B.n516 B.n515 585
R342 B.n513 B.n306 585
R343 B.n306 B.n305 585
R344 B.n512 B.n511 585
R345 B.n511 B.n510 585
R346 B.n308 B.n307 585
R347 B.n309 B.n308 585
R348 B.n503 B.n502 585
R349 B.n504 B.n503 585
R350 B.n501 B.n314 585
R351 B.n314 B.n313 585
R352 B.n500 B.n499 585
R353 B.n499 B.n498 585
R354 B.n316 B.n315 585
R355 B.n317 B.n316 585
R356 B.n491 B.n490 585
R357 B.n492 B.n491 585
R358 B.n489 B.n321 585
R359 B.n325 B.n321 585
R360 B.n488 B.n487 585
R361 B.n487 B.n486 585
R362 B.n323 B.n322 585
R363 B.n324 B.n323 585
R364 B.n479 B.n478 585
R365 B.n480 B.n479 585
R366 B.n477 B.n330 585
R367 B.n330 B.n329 585
R368 B.n476 B.n475 585
R369 B.n475 B.n474 585
R370 B.n332 B.n331 585
R371 B.n333 B.n332 585
R372 B.n467 B.n466 585
R373 B.n468 B.n467 585
R374 B.n465 B.n338 585
R375 B.n338 B.n337 585
R376 B.n464 B.n463 585
R377 B.n463 B.n462 585
R378 B.n459 B.n342 585
R379 B.n458 B.n457 585
R380 B.n455 B.n343 585
R381 B.n455 B.n341 585
R382 B.n454 B.n453 585
R383 B.n452 B.n451 585
R384 B.n450 B.n345 585
R385 B.n448 B.n447 585
R386 B.n446 B.n346 585
R387 B.n445 B.n444 585
R388 B.n442 B.n347 585
R389 B.n440 B.n439 585
R390 B.n438 B.n348 585
R391 B.n437 B.n436 585
R392 B.n434 B.n349 585
R393 B.n432 B.n431 585
R394 B.n430 B.n350 585
R395 B.n429 B.n428 585
R396 B.n426 B.n351 585
R397 B.n424 B.n423 585
R398 B.n422 B.n352 585
R399 B.n421 B.n420 585
R400 B.n418 B.n356 585
R401 B.n416 B.n415 585
R402 B.n414 B.n357 585
R403 B.n413 B.n412 585
R404 B.n410 B.n358 585
R405 B.n408 B.n407 585
R406 B.n406 B.n359 585
R407 B.n404 B.n403 585
R408 B.n401 B.n362 585
R409 B.n399 B.n398 585
R410 B.n397 B.n363 585
R411 B.n396 B.n395 585
R412 B.n393 B.n364 585
R413 B.n391 B.n390 585
R414 B.n389 B.n365 585
R415 B.n388 B.n387 585
R416 B.n385 B.n366 585
R417 B.n383 B.n382 585
R418 B.n381 B.n367 585
R419 B.n380 B.n379 585
R420 B.n377 B.n368 585
R421 B.n375 B.n374 585
R422 B.n373 B.n369 585
R423 B.n372 B.n371 585
R424 B.n340 B.n339 585
R425 B.n341 B.n340 585
R426 B.n461 B.n460 585
R427 B.n462 B.n461 585
R428 B.n336 B.n335 585
R429 B.n337 B.n336 585
R430 B.n470 B.n469 585
R431 B.n469 B.n468 585
R432 B.n471 B.n334 585
R433 B.n334 B.n333 585
R434 B.n473 B.n472 585
R435 B.n474 B.n473 585
R436 B.n328 B.n327 585
R437 B.n329 B.n328 585
R438 B.n482 B.n481 585
R439 B.n481 B.n480 585
R440 B.n483 B.n326 585
R441 B.n326 B.n324 585
R442 B.n485 B.n484 585
R443 B.n486 B.n485 585
R444 B.n320 B.n319 585
R445 B.n325 B.n320 585
R446 B.n494 B.n493 585
R447 B.n493 B.n492 585
R448 B.n495 B.n318 585
R449 B.n318 B.n317 585
R450 B.n497 B.n496 585
R451 B.n498 B.n497 585
R452 B.n312 B.n311 585
R453 B.n313 B.n312 585
R454 B.n506 B.n505 585
R455 B.n505 B.n504 585
R456 B.n507 B.n310 585
R457 B.n310 B.n309 585
R458 B.n509 B.n508 585
R459 B.n510 B.n509 585
R460 B.n304 B.n303 585
R461 B.n305 B.n304 585
R462 B.n518 B.n517 585
R463 B.n517 B.n516 585
R464 B.n519 B.n302 585
R465 B.n302 B.n301 585
R466 B.n521 B.n520 585
R467 B.n522 B.n521 585
R468 B.n296 B.n295 585
R469 B.n297 B.n296 585
R470 B.n530 B.n529 585
R471 B.n529 B.n528 585
R472 B.n531 B.n294 585
R473 B.n294 B.n293 585
R474 B.n533 B.n532 585
R475 B.n534 B.n533 585
R476 B.n288 B.n287 585
R477 B.n289 B.n288 585
R478 B.n542 B.n541 585
R479 B.n541 B.n540 585
R480 B.n543 B.n286 585
R481 B.n286 B.n285 585
R482 B.n545 B.n544 585
R483 B.n546 B.n545 585
R484 B.n280 B.n279 585
R485 B.n281 B.n280 585
R486 B.n554 B.n553 585
R487 B.n553 B.n552 585
R488 B.n555 B.n278 585
R489 B.n278 B.n277 585
R490 B.n557 B.n556 585
R491 B.n558 B.n557 585
R492 B.n272 B.n271 585
R493 B.n273 B.n272 585
R494 B.n566 B.n565 585
R495 B.n565 B.n564 585
R496 B.n567 B.n270 585
R497 B.n270 B.n268 585
R498 B.n569 B.n568 585
R499 B.n570 B.n569 585
R500 B.n264 B.n263 585
R501 B.n269 B.n264 585
R502 B.n578 B.n577 585
R503 B.n577 B.n576 585
R504 B.n579 B.n262 585
R505 B.n262 B.n261 585
R506 B.n581 B.n580 585
R507 B.n582 B.n581 585
R508 B.n256 B.n255 585
R509 B.n257 B.n256 585
R510 B.n590 B.n589 585
R511 B.n589 B.n588 585
R512 B.n591 B.n254 585
R513 B.n254 B.n253 585
R514 B.n593 B.n592 585
R515 B.n594 B.n593 585
R516 B.n248 B.n247 585
R517 B.n249 B.n248 585
R518 B.n602 B.n601 585
R519 B.n601 B.n600 585
R520 B.n603 B.n246 585
R521 B.n246 B.n244 585
R522 B.n605 B.n604 585
R523 B.n606 B.n605 585
R524 B.n240 B.n239 585
R525 B.n245 B.n240 585
R526 B.n614 B.n613 585
R527 B.n613 B.n612 585
R528 B.n615 B.n238 585
R529 B.n238 B.n237 585
R530 B.n617 B.n616 585
R531 B.n618 B.n617 585
R532 B.n232 B.n231 585
R533 B.n233 B.n232 585
R534 B.n626 B.n625 585
R535 B.n625 B.n624 585
R536 B.n627 B.n230 585
R537 B.n230 B.n229 585
R538 B.n629 B.n628 585
R539 B.n630 B.n629 585
R540 B.n224 B.n223 585
R541 B.n225 B.n224 585
R542 B.n638 B.n637 585
R543 B.n637 B.n636 585
R544 B.n639 B.n222 585
R545 B.n222 B.n221 585
R546 B.n641 B.n640 585
R547 B.n642 B.n641 585
R548 B.n216 B.n215 585
R549 B.n217 B.n216 585
R550 B.n650 B.n649 585
R551 B.n649 B.n648 585
R552 B.n651 B.n214 585
R553 B.n214 B.n213 585
R554 B.n653 B.n652 585
R555 B.n654 B.n653 585
R556 B.n208 B.n207 585
R557 B.n209 B.n208 585
R558 B.n662 B.n661 585
R559 B.n661 B.n660 585
R560 B.n663 B.n206 585
R561 B.n206 B.n205 585
R562 B.n665 B.n664 585
R563 B.n666 B.n665 585
R564 B.n200 B.n199 585
R565 B.n201 B.n200 585
R566 B.n674 B.n673 585
R567 B.n673 B.n672 585
R568 B.n675 B.n198 585
R569 B.n198 B.n197 585
R570 B.n677 B.n676 585
R571 B.n678 B.n677 585
R572 B.n192 B.n191 585
R573 B.n193 B.n192 585
R574 B.n686 B.n685 585
R575 B.n685 B.n684 585
R576 B.n687 B.n190 585
R577 B.n190 B.n189 585
R578 B.n689 B.n688 585
R579 B.n690 B.n689 585
R580 B.n184 B.n183 585
R581 B.n185 B.n184 585
R582 B.n699 B.n698 585
R583 B.n698 B.n697 585
R584 B.n700 B.n182 585
R585 B.n182 B.n181 585
R586 B.n702 B.n701 585
R587 B.n703 B.n702 585
R588 B.n3 B.n0 585
R589 B.n4 B.n3 585
R590 B.n1066 B.n1 585
R591 B.n1067 B.n1066 585
R592 B.n1065 B.n1064 585
R593 B.n1065 B.n8 585
R594 B.n1063 B.n9 585
R595 B.n12 B.n9 585
R596 B.n1062 B.n1061 585
R597 B.n1061 B.n1060 585
R598 B.n11 B.n10 585
R599 B.n1059 B.n11 585
R600 B.n1057 B.n1056 585
R601 B.n1058 B.n1057 585
R602 B.n1055 B.n17 585
R603 B.n17 B.n16 585
R604 B.n1054 B.n1053 585
R605 B.n1053 B.n1052 585
R606 B.n19 B.n18 585
R607 B.n1051 B.n19 585
R608 B.n1049 B.n1048 585
R609 B.n1050 B.n1049 585
R610 B.n1047 B.n24 585
R611 B.n24 B.n23 585
R612 B.n1046 B.n1045 585
R613 B.n1045 B.n1044 585
R614 B.n26 B.n25 585
R615 B.n1043 B.n26 585
R616 B.n1041 B.n1040 585
R617 B.n1042 B.n1041 585
R618 B.n1039 B.n31 585
R619 B.n31 B.n30 585
R620 B.n1038 B.n1037 585
R621 B.n1037 B.n1036 585
R622 B.n33 B.n32 585
R623 B.n1035 B.n33 585
R624 B.n1033 B.n1032 585
R625 B.n1034 B.n1033 585
R626 B.n1031 B.n38 585
R627 B.n38 B.n37 585
R628 B.n1030 B.n1029 585
R629 B.n1029 B.n1028 585
R630 B.n40 B.n39 585
R631 B.n1027 B.n40 585
R632 B.n1025 B.n1024 585
R633 B.n1026 B.n1025 585
R634 B.n1023 B.n45 585
R635 B.n45 B.n44 585
R636 B.n1022 B.n1021 585
R637 B.n1021 B.n1020 585
R638 B.n47 B.n46 585
R639 B.n1019 B.n47 585
R640 B.n1017 B.n1016 585
R641 B.n1018 B.n1017 585
R642 B.n1015 B.n52 585
R643 B.n52 B.n51 585
R644 B.n1014 B.n1013 585
R645 B.n1013 B.n1012 585
R646 B.n54 B.n53 585
R647 B.n1011 B.n54 585
R648 B.n1009 B.n1008 585
R649 B.n1010 B.n1009 585
R650 B.n1007 B.n59 585
R651 B.n59 B.n58 585
R652 B.n1006 B.n1005 585
R653 B.n1005 B.n1004 585
R654 B.n61 B.n60 585
R655 B.n1003 B.n61 585
R656 B.n1001 B.n1000 585
R657 B.n1002 B.n1001 585
R658 B.n999 B.n66 585
R659 B.n66 B.n65 585
R660 B.n998 B.n997 585
R661 B.n997 B.n996 585
R662 B.n68 B.n67 585
R663 B.n995 B.n68 585
R664 B.n993 B.n992 585
R665 B.n994 B.n993 585
R666 B.n991 B.n73 585
R667 B.n73 B.n72 585
R668 B.n990 B.n989 585
R669 B.n989 B.n988 585
R670 B.n75 B.n74 585
R671 B.n987 B.n75 585
R672 B.n985 B.n984 585
R673 B.n986 B.n985 585
R674 B.n983 B.n80 585
R675 B.n80 B.n79 585
R676 B.n982 B.n981 585
R677 B.n981 B.n980 585
R678 B.n82 B.n81 585
R679 B.n979 B.n82 585
R680 B.n977 B.n976 585
R681 B.n978 B.n977 585
R682 B.n975 B.n87 585
R683 B.n87 B.n86 585
R684 B.n974 B.n973 585
R685 B.n973 B.n972 585
R686 B.n89 B.n88 585
R687 B.n971 B.n89 585
R688 B.n969 B.n968 585
R689 B.n970 B.n969 585
R690 B.n967 B.n94 585
R691 B.n94 B.n93 585
R692 B.n966 B.n965 585
R693 B.n965 B.n964 585
R694 B.n96 B.n95 585
R695 B.n963 B.n96 585
R696 B.n961 B.n960 585
R697 B.n962 B.n961 585
R698 B.n959 B.n101 585
R699 B.n101 B.n100 585
R700 B.n958 B.n957 585
R701 B.n957 B.n956 585
R702 B.n103 B.n102 585
R703 B.n955 B.n103 585
R704 B.n953 B.n952 585
R705 B.n954 B.n953 585
R706 B.n951 B.n108 585
R707 B.n108 B.n107 585
R708 B.n950 B.n949 585
R709 B.n949 B.n948 585
R710 B.n110 B.n109 585
R711 B.n947 B.n110 585
R712 B.n945 B.n944 585
R713 B.n946 B.n945 585
R714 B.n943 B.n115 585
R715 B.n115 B.n114 585
R716 B.n942 B.n941 585
R717 B.n941 B.n940 585
R718 B.n117 B.n116 585
R719 B.n939 B.n117 585
R720 B.n937 B.n936 585
R721 B.n938 B.n937 585
R722 B.n935 B.n122 585
R723 B.n122 B.n121 585
R724 B.n934 B.n933 585
R725 B.n933 B.n932 585
R726 B.n124 B.n123 585
R727 B.n931 B.n124 585
R728 B.n929 B.n928 585
R729 B.n930 B.n929 585
R730 B.n927 B.n129 585
R731 B.n129 B.n128 585
R732 B.n926 B.n925 585
R733 B.n925 B.n924 585
R734 B.n131 B.n130 585
R735 B.n923 B.n131 585
R736 B.n921 B.n920 585
R737 B.n922 B.n921 585
R738 B.n919 B.n136 585
R739 B.n136 B.n135 585
R740 B.n918 B.n917 585
R741 B.n917 B.n916 585
R742 B.n138 B.n137 585
R743 B.n915 B.n138 585
R744 B.n913 B.n912 585
R745 B.n914 B.n913 585
R746 B.n911 B.n143 585
R747 B.n143 B.n142 585
R748 B.n910 B.n909 585
R749 B.n909 B.n908 585
R750 B.n145 B.n144 585
R751 B.n907 B.n145 585
R752 B.n905 B.n904 585
R753 B.n906 B.n905 585
R754 B.n1070 B.n1069 585
R755 B.n1068 B.n2 585
R756 B.n905 B.n150 535.745
R757 B.n813 B.n148 535.745
R758 B.n463 B.n340 535.745
R759 B.n461 B.n342 535.745
R760 B.n812 B.n149 256.663
R761 B.n818 B.n149 256.663
R762 B.n820 B.n149 256.663
R763 B.n826 B.n149 256.663
R764 B.n828 B.n149 256.663
R765 B.n834 B.n149 256.663
R766 B.n836 B.n149 256.663
R767 B.n842 B.n149 256.663
R768 B.n170 B.n149 256.663
R769 B.n848 B.n149 256.663
R770 B.n854 B.n149 256.663
R771 B.n856 B.n149 256.663
R772 B.n862 B.n149 256.663
R773 B.n162 B.n149 256.663
R774 B.n868 B.n149 256.663
R775 B.n874 B.n149 256.663
R776 B.n876 B.n149 256.663
R777 B.n882 B.n149 256.663
R778 B.n884 B.n149 256.663
R779 B.n890 B.n149 256.663
R780 B.n892 B.n149 256.663
R781 B.n898 B.n149 256.663
R782 B.n900 B.n149 256.663
R783 B.n456 B.n341 256.663
R784 B.n344 B.n341 256.663
R785 B.n449 B.n341 256.663
R786 B.n443 B.n341 256.663
R787 B.n441 B.n341 256.663
R788 B.n435 B.n341 256.663
R789 B.n433 B.n341 256.663
R790 B.n427 B.n341 256.663
R791 B.n425 B.n341 256.663
R792 B.n419 B.n341 256.663
R793 B.n417 B.n341 256.663
R794 B.n411 B.n341 256.663
R795 B.n409 B.n341 256.663
R796 B.n402 B.n341 256.663
R797 B.n400 B.n341 256.663
R798 B.n394 B.n341 256.663
R799 B.n392 B.n341 256.663
R800 B.n386 B.n341 256.663
R801 B.n384 B.n341 256.663
R802 B.n378 B.n341 256.663
R803 B.n376 B.n341 256.663
R804 B.n370 B.n341 256.663
R805 B.n1072 B.n1071 256.663
R806 B.n159 B.t10 234.322
R807 B.n167 B.t21 234.322
R808 B.n360 B.t14 234.322
R809 B.n353 B.t18 234.322
R810 B.n167 B.t22 227.879
R811 B.n360 B.t17 227.879
R812 B.n159 B.t12 227.879
R813 B.n353 B.t20 227.879
R814 B.n462 B.n341 166.685
R815 B.n906 B.n149 166.685
R816 B.n901 B.n899 163.367
R817 B.n897 B.n152 163.367
R818 B.n893 B.n891 163.367
R819 B.n889 B.n154 163.367
R820 B.n885 B.n883 163.367
R821 B.n881 B.n156 163.367
R822 B.n877 B.n875 163.367
R823 B.n873 B.n158 163.367
R824 B.n869 B.n867 163.367
R825 B.n864 B.n863 163.367
R826 B.n861 B.n164 163.367
R827 B.n857 B.n855 163.367
R828 B.n853 B.n166 163.367
R829 B.n849 B.n847 163.367
R830 B.n844 B.n843 163.367
R831 B.n841 B.n172 163.367
R832 B.n837 B.n835 163.367
R833 B.n833 B.n174 163.367
R834 B.n829 B.n827 163.367
R835 B.n825 B.n176 163.367
R836 B.n821 B.n819 163.367
R837 B.n817 B.n178 163.367
R838 B.n463 B.n338 163.367
R839 B.n467 B.n338 163.367
R840 B.n467 B.n332 163.367
R841 B.n475 B.n332 163.367
R842 B.n475 B.n330 163.367
R843 B.n479 B.n330 163.367
R844 B.n479 B.n323 163.367
R845 B.n487 B.n323 163.367
R846 B.n487 B.n321 163.367
R847 B.n491 B.n321 163.367
R848 B.n491 B.n316 163.367
R849 B.n499 B.n316 163.367
R850 B.n499 B.n314 163.367
R851 B.n503 B.n314 163.367
R852 B.n503 B.n308 163.367
R853 B.n511 B.n308 163.367
R854 B.n511 B.n306 163.367
R855 B.n515 B.n306 163.367
R856 B.n515 B.n300 163.367
R857 B.n523 B.n300 163.367
R858 B.n523 B.n298 163.367
R859 B.n527 B.n298 163.367
R860 B.n527 B.n292 163.367
R861 B.n535 B.n292 163.367
R862 B.n535 B.n290 163.367
R863 B.n539 B.n290 163.367
R864 B.n539 B.n284 163.367
R865 B.n547 B.n284 163.367
R866 B.n547 B.n282 163.367
R867 B.n551 B.n282 163.367
R868 B.n551 B.n276 163.367
R869 B.n559 B.n276 163.367
R870 B.n559 B.n274 163.367
R871 B.n563 B.n274 163.367
R872 B.n563 B.n267 163.367
R873 B.n571 B.n267 163.367
R874 B.n571 B.n265 163.367
R875 B.n575 B.n265 163.367
R876 B.n575 B.n260 163.367
R877 B.n583 B.n260 163.367
R878 B.n583 B.n258 163.367
R879 B.n587 B.n258 163.367
R880 B.n587 B.n252 163.367
R881 B.n595 B.n252 163.367
R882 B.n595 B.n250 163.367
R883 B.n599 B.n250 163.367
R884 B.n599 B.n243 163.367
R885 B.n607 B.n243 163.367
R886 B.n607 B.n241 163.367
R887 B.n611 B.n241 163.367
R888 B.n611 B.n236 163.367
R889 B.n619 B.n236 163.367
R890 B.n619 B.n234 163.367
R891 B.n623 B.n234 163.367
R892 B.n623 B.n228 163.367
R893 B.n631 B.n228 163.367
R894 B.n631 B.n226 163.367
R895 B.n635 B.n226 163.367
R896 B.n635 B.n220 163.367
R897 B.n643 B.n220 163.367
R898 B.n643 B.n218 163.367
R899 B.n647 B.n218 163.367
R900 B.n647 B.n212 163.367
R901 B.n655 B.n212 163.367
R902 B.n655 B.n210 163.367
R903 B.n659 B.n210 163.367
R904 B.n659 B.n204 163.367
R905 B.n667 B.n204 163.367
R906 B.n667 B.n202 163.367
R907 B.n671 B.n202 163.367
R908 B.n671 B.n196 163.367
R909 B.n679 B.n196 163.367
R910 B.n679 B.n194 163.367
R911 B.n683 B.n194 163.367
R912 B.n683 B.n188 163.367
R913 B.n691 B.n188 163.367
R914 B.n691 B.n186 163.367
R915 B.n696 B.n186 163.367
R916 B.n696 B.n180 163.367
R917 B.n704 B.n180 163.367
R918 B.n705 B.n704 163.367
R919 B.n705 B.n5 163.367
R920 B.n6 B.n5 163.367
R921 B.n7 B.n6 163.367
R922 B.n711 B.n7 163.367
R923 B.n712 B.n711 163.367
R924 B.n712 B.n13 163.367
R925 B.n14 B.n13 163.367
R926 B.n15 B.n14 163.367
R927 B.n717 B.n15 163.367
R928 B.n717 B.n20 163.367
R929 B.n21 B.n20 163.367
R930 B.n22 B.n21 163.367
R931 B.n722 B.n22 163.367
R932 B.n722 B.n27 163.367
R933 B.n28 B.n27 163.367
R934 B.n29 B.n28 163.367
R935 B.n727 B.n29 163.367
R936 B.n727 B.n34 163.367
R937 B.n35 B.n34 163.367
R938 B.n36 B.n35 163.367
R939 B.n732 B.n36 163.367
R940 B.n732 B.n41 163.367
R941 B.n42 B.n41 163.367
R942 B.n43 B.n42 163.367
R943 B.n737 B.n43 163.367
R944 B.n737 B.n48 163.367
R945 B.n49 B.n48 163.367
R946 B.n50 B.n49 163.367
R947 B.n742 B.n50 163.367
R948 B.n742 B.n55 163.367
R949 B.n56 B.n55 163.367
R950 B.n57 B.n56 163.367
R951 B.n747 B.n57 163.367
R952 B.n747 B.n62 163.367
R953 B.n63 B.n62 163.367
R954 B.n64 B.n63 163.367
R955 B.n752 B.n64 163.367
R956 B.n752 B.n69 163.367
R957 B.n70 B.n69 163.367
R958 B.n71 B.n70 163.367
R959 B.n757 B.n71 163.367
R960 B.n757 B.n76 163.367
R961 B.n77 B.n76 163.367
R962 B.n78 B.n77 163.367
R963 B.n762 B.n78 163.367
R964 B.n762 B.n83 163.367
R965 B.n84 B.n83 163.367
R966 B.n85 B.n84 163.367
R967 B.n767 B.n85 163.367
R968 B.n767 B.n90 163.367
R969 B.n91 B.n90 163.367
R970 B.n92 B.n91 163.367
R971 B.n772 B.n92 163.367
R972 B.n772 B.n97 163.367
R973 B.n98 B.n97 163.367
R974 B.n99 B.n98 163.367
R975 B.n777 B.n99 163.367
R976 B.n777 B.n104 163.367
R977 B.n105 B.n104 163.367
R978 B.n106 B.n105 163.367
R979 B.n782 B.n106 163.367
R980 B.n782 B.n111 163.367
R981 B.n112 B.n111 163.367
R982 B.n113 B.n112 163.367
R983 B.n787 B.n113 163.367
R984 B.n787 B.n118 163.367
R985 B.n119 B.n118 163.367
R986 B.n120 B.n119 163.367
R987 B.n792 B.n120 163.367
R988 B.n792 B.n125 163.367
R989 B.n126 B.n125 163.367
R990 B.n127 B.n126 163.367
R991 B.n797 B.n127 163.367
R992 B.n797 B.n132 163.367
R993 B.n133 B.n132 163.367
R994 B.n134 B.n133 163.367
R995 B.n802 B.n134 163.367
R996 B.n802 B.n139 163.367
R997 B.n140 B.n139 163.367
R998 B.n141 B.n140 163.367
R999 B.n807 B.n141 163.367
R1000 B.n807 B.n146 163.367
R1001 B.n147 B.n146 163.367
R1002 B.n148 B.n147 163.367
R1003 B.n457 B.n455 163.367
R1004 B.n455 B.n454 163.367
R1005 B.n451 B.n450 163.367
R1006 B.n448 B.n346 163.367
R1007 B.n444 B.n442 163.367
R1008 B.n440 B.n348 163.367
R1009 B.n436 B.n434 163.367
R1010 B.n432 B.n350 163.367
R1011 B.n428 B.n426 163.367
R1012 B.n424 B.n352 163.367
R1013 B.n420 B.n418 163.367
R1014 B.n416 B.n357 163.367
R1015 B.n412 B.n410 163.367
R1016 B.n408 B.n359 163.367
R1017 B.n403 B.n401 163.367
R1018 B.n399 B.n363 163.367
R1019 B.n395 B.n393 163.367
R1020 B.n391 B.n365 163.367
R1021 B.n387 B.n385 163.367
R1022 B.n383 B.n367 163.367
R1023 B.n379 B.n377 163.367
R1024 B.n375 B.n369 163.367
R1025 B.n371 B.n340 163.367
R1026 B.n461 B.n336 163.367
R1027 B.n469 B.n336 163.367
R1028 B.n469 B.n334 163.367
R1029 B.n473 B.n334 163.367
R1030 B.n473 B.n328 163.367
R1031 B.n481 B.n328 163.367
R1032 B.n481 B.n326 163.367
R1033 B.n485 B.n326 163.367
R1034 B.n485 B.n320 163.367
R1035 B.n493 B.n320 163.367
R1036 B.n493 B.n318 163.367
R1037 B.n497 B.n318 163.367
R1038 B.n497 B.n312 163.367
R1039 B.n505 B.n312 163.367
R1040 B.n505 B.n310 163.367
R1041 B.n509 B.n310 163.367
R1042 B.n509 B.n304 163.367
R1043 B.n517 B.n304 163.367
R1044 B.n517 B.n302 163.367
R1045 B.n521 B.n302 163.367
R1046 B.n521 B.n296 163.367
R1047 B.n529 B.n296 163.367
R1048 B.n529 B.n294 163.367
R1049 B.n533 B.n294 163.367
R1050 B.n533 B.n288 163.367
R1051 B.n541 B.n288 163.367
R1052 B.n541 B.n286 163.367
R1053 B.n545 B.n286 163.367
R1054 B.n545 B.n280 163.367
R1055 B.n553 B.n280 163.367
R1056 B.n553 B.n278 163.367
R1057 B.n557 B.n278 163.367
R1058 B.n557 B.n272 163.367
R1059 B.n565 B.n272 163.367
R1060 B.n565 B.n270 163.367
R1061 B.n569 B.n270 163.367
R1062 B.n569 B.n264 163.367
R1063 B.n577 B.n264 163.367
R1064 B.n577 B.n262 163.367
R1065 B.n581 B.n262 163.367
R1066 B.n581 B.n256 163.367
R1067 B.n589 B.n256 163.367
R1068 B.n589 B.n254 163.367
R1069 B.n593 B.n254 163.367
R1070 B.n593 B.n248 163.367
R1071 B.n601 B.n248 163.367
R1072 B.n601 B.n246 163.367
R1073 B.n605 B.n246 163.367
R1074 B.n605 B.n240 163.367
R1075 B.n613 B.n240 163.367
R1076 B.n613 B.n238 163.367
R1077 B.n617 B.n238 163.367
R1078 B.n617 B.n232 163.367
R1079 B.n625 B.n232 163.367
R1080 B.n625 B.n230 163.367
R1081 B.n629 B.n230 163.367
R1082 B.n629 B.n224 163.367
R1083 B.n637 B.n224 163.367
R1084 B.n637 B.n222 163.367
R1085 B.n641 B.n222 163.367
R1086 B.n641 B.n216 163.367
R1087 B.n649 B.n216 163.367
R1088 B.n649 B.n214 163.367
R1089 B.n653 B.n214 163.367
R1090 B.n653 B.n208 163.367
R1091 B.n661 B.n208 163.367
R1092 B.n661 B.n206 163.367
R1093 B.n665 B.n206 163.367
R1094 B.n665 B.n200 163.367
R1095 B.n673 B.n200 163.367
R1096 B.n673 B.n198 163.367
R1097 B.n677 B.n198 163.367
R1098 B.n677 B.n192 163.367
R1099 B.n685 B.n192 163.367
R1100 B.n685 B.n190 163.367
R1101 B.n689 B.n190 163.367
R1102 B.n689 B.n184 163.367
R1103 B.n698 B.n184 163.367
R1104 B.n698 B.n182 163.367
R1105 B.n702 B.n182 163.367
R1106 B.n702 B.n3 163.367
R1107 B.n1070 B.n3 163.367
R1108 B.n1066 B.n2 163.367
R1109 B.n1066 B.n1065 163.367
R1110 B.n1065 B.n9 163.367
R1111 B.n1061 B.n9 163.367
R1112 B.n1061 B.n11 163.367
R1113 B.n1057 B.n11 163.367
R1114 B.n1057 B.n17 163.367
R1115 B.n1053 B.n17 163.367
R1116 B.n1053 B.n19 163.367
R1117 B.n1049 B.n19 163.367
R1118 B.n1049 B.n24 163.367
R1119 B.n1045 B.n24 163.367
R1120 B.n1045 B.n26 163.367
R1121 B.n1041 B.n26 163.367
R1122 B.n1041 B.n31 163.367
R1123 B.n1037 B.n31 163.367
R1124 B.n1037 B.n33 163.367
R1125 B.n1033 B.n33 163.367
R1126 B.n1033 B.n38 163.367
R1127 B.n1029 B.n38 163.367
R1128 B.n1029 B.n40 163.367
R1129 B.n1025 B.n40 163.367
R1130 B.n1025 B.n45 163.367
R1131 B.n1021 B.n45 163.367
R1132 B.n1021 B.n47 163.367
R1133 B.n1017 B.n47 163.367
R1134 B.n1017 B.n52 163.367
R1135 B.n1013 B.n52 163.367
R1136 B.n1013 B.n54 163.367
R1137 B.n1009 B.n54 163.367
R1138 B.n1009 B.n59 163.367
R1139 B.n1005 B.n59 163.367
R1140 B.n1005 B.n61 163.367
R1141 B.n1001 B.n61 163.367
R1142 B.n1001 B.n66 163.367
R1143 B.n997 B.n66 163.367
R1144 B.n997 B.n68 163.367
R1145 B.n993 B.n68 163.367
R1146 B.n993 B.n73 163.367
R1147 B.n989 B.n73 163.367
R1148 B.n989 B.n75 163.367
R1149 B.n985 B.n75 163.367
R1150 B.n985 B.n80 163.367
R1151 B.n981 B.n80 163.367
R1152 B.n981 B.n82 163.367
R1153 B.n977 B.n82 163.367
R1154 B.n977 B.n87 163.367
R1155 B.n973 B.n87 163.367
R1156 B.n973 B.n89 163.367
R1157 B.n969 B.n89 163.367
R1158 B.n969 B.n94 163.367
R1159 B.n965 B.n94 163.367
R1160 B.n965 B.n96 163.367
R1161 B.n961 B.n96 163.367
R1162 B.n961 B.n101 163.367
R1163 B.n957 B.n101 163.367
R1164 B.n957 B.n103 163.367
R1165 B.n953 B.n103 163.367
R1166 B.n953 B.n108 163.367
R1167 B.n949 B.n108 163.367
R1168 B.n949 B.n110 163.367
R1169 B.n945 B.n110 163.367
R1170 B.n945 B.n115 163.367
R1171 B.n941 B.n115 163.367
R1172 B.n941 B.n117 163.367
R1173 B.n937 B.n117 163.367
R1174 B.n937 B.n122 163.367
R1175 B.n933 B.n122 163.367
R1176 B.n933 B.n124 163.367
R1177 B.n929 B.n124 163.367
R1178 B.n929 B.n129 163.367
R1179 B.n925 B.n129 163.367
R1180 B.n925 B.n131 163.367
R1181 B.n921 B.n131 163.367
R1182 B.n921 B.n136 163.367
R1183 B.n917 B.n136 163.367
R1184 B.n917 B.n138 163.367
R1185 B.n913 B.n138 163.367
R1186 B.n913 B.n143 163.367
R1187 B.n909 B.n143 163.367
R1188 B.n909 B.n145 163.367
R1189 B.n905 B.n145 163.367
R1190 B.n168 B.t23 145.843
R1191 B.n361 B.t16 145.843
R1192 B.n160 B.t13 145.841
R1193 B.n354 B.t19 145.841
R1194 B.n160 B.n159 82.0369
R1195 B.n168 B.n167 82.0369
R1196 B.n361 B.n360 82.0369
R1197 B.n354 B.n353 82.0369
R1198 B.n462 B.n337 80.3874
R1199 B.n468 B.n337 80.3874
R1200 B.n468 B.n333 80.3874
R1201 B.n474 B.n333 80.3874
R1202 B.n474 B.n329 80.3874
R1203 B.n480 B.n329 80.3874
R1204 B.n480 B.n324 80.3874
R1205 B.n486 B.n324 80.3874
R1206 B.n486 B.n325 80.3874
R1207 B.n492 B.n317 80.3874
R1208 B.n498 B.n317 80.3874
R1209 B.n498 B.n313 80.3874
R1210 B.n504 B.n313 80.3874
R1211 B.n504 B.n309 80.3874
R1212 B.n510 B.n309 80.3874
R1213 B.n510 B.n305 80.3874
R1214 B.n516 B.n305 80.3874
R1215 B.n516 B.n301 80.3874
R1216 B.n522 B.n301 80.3874
R1217 B.n522 B.n297 80.3874
R1218 B.n528 B.n297 80.3874
R1219 B.n528 B.n293 80.3874
R1220 B.n534 B.n293 80.3874
R1221 B.n540 B.n289 80.3874
R1222 B.n540 B.n285 80.3874
R1223 B.n546 B.n285 80.3874
R1224 B.n546 B.n281 80.3874
R1225 B.n552 B.n281 80.3874
R1226 B.n552 B.n277 80.3874
R1227 B.n558 B.n277 80.3874
R1228 B.n558 B.n273 80.3874
R1229 B.n564 B.n273 80.3874
R1230 B.n564 B.n268 80.3874
R1231 B.n570 B.n268 80.3874
R1232 B.n570 B.n269 80.3874
R1233 B.n576 B.n261 80.3874
R1234 B.n582 B.n261 80.3874
R1235 B.n582 B.n257 80.3874
R1236 B.n588 B.n257 80.3874
R1237 B.n588 B.n253 80.3874
R1238 B.n594 B.n253 80.3874
R1239 B.n594 B.n249 80.3874
R1240 B.n600 B.n249 80.3874
R1241 B.n600 B.n244 80.3874
R1242 B.n606 B.n244 80.3874
R1243 B.n606 B.n245 80.3874
R1244 B.n612 B.n237 80.3874
R1245 B.n618 B.n237 80.3874
R1246 B.n618 B.n233 80.3874
R1247 B.n624 B.n233 80.3874
R1248 B.n624 B.n229 80.3874
R1249 B.n630 B.n229 80.3874
R1250 B.n630 B.n225 80.3874
R1251 B.n636 B.n225 80.3874
R1252 B.n636 B.n221 80.3874
R1253 B.n642 B.n221 80.3874
R1254 B.n642 B.n217 80.3874
R1255 B.n648 B.n217 80.3874
R1256 B.n654 B.n213 80.3874
R1257 B.n654 B.n209 80.3874
R1258 B.n660 B.n209 80.3874
R1259 B.n660 B.n205 80.3874
R1260 B.n666 B.n205 80.3874
R1261 B.n666 B.n201 80.3874
R1262 B.n672 B.n201 80.3874
R1263 B.n672 B.n197 80.3874
R1264 B.n678 B.n197 80.3874
R1265 B.n678 B.n193 80.3874
R1266 B.n684 B.n193 80.3874
R1267 B.n690 B.n189 80.3874
R1268 B.n690 B.n185 80.3874
R1269 B.n697 B.n185 80.3874
R1270 B.n697 B.n181 80.3874
R1271 B.n703 B.n181 80.3874
R1272 B.n703 B.n4 80.3874
R1273 B.n1069 B.n4 80.3874
R1274 B.n1069 B.n1068 80.3874
R1275 B.n1068 B.n1067 80.3874
R1276 B.n1067 B.n8 80.3874
R1277 B.n12 B.n8 80.3874
R1278 B.n1060 B.n12 80.3874
R1279 B.n1060 B.n1059 80.3874
R1280 B.n1059 B.n1058 80.3874
R1281 B.n1058 B.n16 80.3874
R1282 B.n1052 B.n1051 80.3874
R1283 B.n1051 B.n1050 80.3874
R1284 B.n1050 B.n23 80.3874
R1285 B.n1044 B.n23 80.3874
R1286 B.n1044 B.n1043 80.3874
R1287 B.n1043 B.n1042 80.3874
R1288 B.n1042 B.n30 80.3874
R1289 B.n1036 B.n30 80.3874
R1290 B.n1036 B.n1035 80.3874
R1291 B.n1035 B.n1034 80.3874
R1292 B.n1034 B.n37 80.3874
R1293 B.n1028 B.n1027 80.3874
R1294 B.n1027 B.n1026 80.3874
R1295 B.n1026 B.n44 80.3874
R1296 B.n1020 B.n44 80.3874
R1297 B.n1020 B.n1019 80.3874
R1298 B.n1019 B.n1018 80.3874
R1299 B.n1018 B.n51 80.3874
R1300 B.n1012 B.n51 80.3874
R1301 B.n1012 B.n1011 80.3874
R1302 B.n1011 B.n1010 80.3874
R1303 B.n1010 B.n58 80.3874
R1304 B.n1004 B.n58 80.3874
R1305 B.n1003 B.n1002 80.3874
R1306 B.n1002 B.n65 80.3874
R1307 B.n996 B.n65 80.3874
R1308 B.n996 B.n995 80.3874
R1309 B.n995 B.n994 80.3874
R1310 B.n994 B.n72 80.3874
R1311 B.n988 B.n72 80.3874
R1312 B.n988 B.n987 80.3874
R1313 B.n987 B.n986 80.3874
R1314 B.n986 B.n79 80.3874
R1315 B.n980 B.n79 80.3874
R1316 B.n979 B.n978 80.3874
R1317 B.n978 B.n86 80.3874
R1318 B.n972 B.n86 80.3874
R1319 B.n972 B.n971 80.3874
R1320 B.n971 B.n970 80.3874
R1321 B.n970 B.n93 80.3874
R1322 B.n964 B.n93 80.3874
R1323 B.n964 B.n963 80.3874
R1324 B.n963 B.n962 80.3874
R1325 B.n962 B.n100 80.3874
R1326 B.n956 B.n100 80.3874
R1327 B.n956 B.n955 80.3874
R1328 B.n954 B.n107 80.3874
R1329 B.n948 B.n107 80.3874
R1330 B.n948 B.n947 80.3874
R1331 B.n947 B.n946 80.3874
R1332 B.n946 B.n114 80.3874
R1333 B.n940 B.n114 80.3874
R1334 B.n940 B.n939 80.3874
R1335 B.n939 B.n938 80.3874
R1336 B.n938 B.n121 80.3874
R1337 B.n932 B.n121 80.3874
R1338 B.n932 B.n931 80.3874
R1339 B.n931 B.n930 80.3874
R1340 B.n930 B.n128 80.3874
R1341 B.n924 B.n128 80.3874
R1342 B.n923 B.n922 80.3874
R1343 B.n922 B.n135 80.3874
R1344 B.n916 B.n135 80.3874
R1345 B.n916 B.n915 80.3874
R1346 B.n915 B.n914 80.3874
R1347 B.n914 B.n142 80.3874
R1348 B.n908 B.n142 80.3874
R1349 B.n908 B.n907 80.3874
R1350 B.n907 B.n906 80.3874
R1351 B.n534 B.t0 73.2944
R1352 B.t5 B.n954 73.2944
R1353 B.n900 B.n150 71.676
R1354 B.n899 B.n898 71.676
R1355 B.n892 B.n152 71.676
R1356 B.n891 B.n890 71.676
R1357 B.n884 B.n154 71.676
R1358 B.n883 B.n882 71.676
R1359 B.n876 B.n156 71.676
R1360 B.n875 B.n874 71.676
R1361 B.n868 B.n158 71.676
R1362 B.n867 B.n162 71.676
R1363 B.n863 B.n862 71.676
R1364 B.n856 B.n164 71.676
R1365 B.n855 B.n854 71.676
R1366 B.n848 B.n166 71.676
R1367 B.n847 B.n170 71.676
R1368 B.n843 B.n842 71.676
R1369 B.n836 B.n172 71.676
R1370 B.n835 B.n834 71.676
R1371 B.n828 B.n174 71.676
R1372 B.n827 B.n826 71.676
R1373 B.n820 B.n176 71.676
R1374 B.n819 B.n818 71.676
R1375 B.n812 B.n178 71.676
R1376 B.n813 B.n812 71.676
R1377 B.n818 B.n817 71.676
R1378 B.n821 B.n820 71.676
R1379 B.n826 B.n825 71.676
R1380 B.n829 B.n828 71.676
R1381 B.n834 B.n833 71.676
R1382 B.n837 B.n836 71.676
R1383 B.n842 B.n841 71.676
R1384 B.n844 B.n170 71.676
R1385 B.n849 B.n848 71.676
R1386 B.n854 B.n853 71.676
R1387 B.n857 B.n856 71.676
R1388 B.n862 B.n861 71.676
R1389 B.n864 B.n162 71.676
R1390 B.n869 B.n868 71.676
R1391 B.n874 B.n873 71.676
R1392 B.n877 B.n876 71.676
R1393 B.n882 B.n881 71.676
R1394 B.n885 B.n884 71.676
R1395 B.n890 B.n889 71.676
R1396 B.n893 B.n892 71.676
R1397 B.n898 B.n897 71.676
R1398 B.n901 B.n900 71.676
R1399 B.n456 B.n342 71.676
R1400 B.n454 B.n344 71.676
R1401 B.n450 B.n449 71.676
R1402 B.n443 B.n346 71.676
R1403 B.n442 B.n441 71.676
R1404 B.n435 B.n348 71.676
R1405 B.n434 B.n433 71.676
R1406 B.n427 B.n350 71.676
R1407 B.n426 B.n425 71.676
R1408 B.n419 B.n352 71.676
R1409 B.n418 B.n417 71.676
R1410 B.n411 B.n357 71.676
R1411 B.n410 B.n409 71.676
R1412 B.n402 B.n359 71.676
R1413 B.n401 B.n400 71.676
R1414 B.n394 B.n363 71.676
R1415 B.n393 B.n392 71.676
R1416 B.n386 B.n365 71.676
R1417 B.n385 B.n384 71.676
R1418 B.n378 B.n367 71.676
R1419 B.n377 B.n376 71.676
R1420 B.n370 B.n369 71.676
R1421 B.n457 B.n456 71.676
R1422 B.n451 B.n344 71.676
R1423 B.n449 B.n448 71.676
R1424 B.n444 B.n443 71.676
R1425 B.n441 B.n440 71.676
R1426 B.n436 B.n435 71.676
R1427 B.n433 B.n432 71.676
R1428 B.n428 B.n427 71.676
R1429 B.n425 B.n424 71.676
R1430 B.n420 B.n419 71.676
R1431 B.n417 B.n416 71.676
R1432 B.n412 B.n411 71.676
R1433 B.n409 B.n408 71.676
R1434 B.n403 B.n402 71.676
R1435 B.n400 B.n399 71.676
R1436 B.n395 B.n394 71.676
R1437 B.n392 B.n391 71.676
R1438 B.n387 B.n386 71.676
R1439 B.n384 B.n383 71.676
R1440 B.n379 B.n378 71.676
R1441 B.n376 B.n375 71.676
R1442 B.n371 B.n370 71.676
R1443 B.n1071 B.n1070 71.676
R1444 B.n1071 B.n2 71.676
R1445 B.n245 B.t6 63.8371
R1446 B.t1 B.n1003 63.8371
R1447 B.t9 B.n213 61.4728
R1448 B.t2 B.n37 61.4728
R1449 B.n161 B.n160 59.5399
R1450 B.n169 B.n168 59.5399
R1451 B.n405 B.n361 59.5399
R1452 B.n355 B.n354 59.5399
R1453 B.n492 B.t15 59.1085
R1454 B.n924 B.t11 59.1085
R1455 B.n684 B.t8 54.3799
R1456 B.n1052 B.t7 54.3799
R1457 B.n576 B.t3 52.0155
R1458 B.n980 B.t4 52.0155
R1459 B.n460 B.n459 34.8103
R1460 B.n464 B.n339 34.8103
R1461 B.n814 B.n811 34.8103
R1462 B.n904 B.n903 34.8103
R1463 B.n269 B.t3 28.3723
R1464 B.t4 B.n979 28.3723
R1465 B.t8 B.n189 26.008
R1466 B.t7 B.n16 26.008
R1467 B.n325 B.t15 21.2794
R1468 B.t11 B.n923 21.2794
R1469 B.n648 B.t9 18.9151
R1470 B.n1028 B.t2 18.9151
R1471 B B.n1072 18.0485
R1472 B.n612 B.t6 16.5507
R1473 B.n1004 B.t1 16.5507
R1474 B.n460 B.n335 10.6151
R1475 B.n470 B.n335 10.6151
R1476 B.n471 B.n470 10.6151
R1477 B.n472 B.n471 10.6151
R1478 B.n472 B.n327 10.6151
R1479 B.n482 B.n327 10.6151
R1480 B.n483 B.n482 10.6151
R1481 B.n484 B.n483 10.6151
R1482 B.n484 B.n319 10.6151
R1483 B.n494 B.n319 10.6151
R1484 B.n495 B.n494 10.6151
R1485 B.n496 B.n495 10.6151
R1486 B.n496 B.n311 10.6151
R1487 B.n506 B.n311 10.6151
R1488 B.n507 B.n506 10.6151
R1489 B.n508 B.n507 10.6151
R1490 B.n508 B.n303 10.6151
R1491 B.n518 B.n303 10.6151
R1492 B.n519 B.n518 10.6151
R1493 B.n520 B.n519 10.6151
R1494 B.n520 B.n295 10.6151
R1495 B.n530 B.n295 10.6151
R1496 B.n531 B.n530 10.6151
R1497 B.n532 B.n531 10.6151
R1498 B.n532 B.n287 10.6151
R1499 B.n542 B.n287 10.6151
R1500 B.n543 B.n542 10.6151
R1501 B.n544 B.n543 10.6151
R1502 B.n544 B.n279 10.6151
R1503 B.n554 B.n279 10.6151
R1504 B.n555 B.n554 10.6151
R1505 B.n556 B.n555 10.6151
R1506 B.n556 B.n271 10.6151
R1507 B.n566 B.n271 10.6151
R1508 B.n567 B.n566 10.6151
R1509 B.n568 B.n567 10.6151
R1510 B.n568 B.n263 10.6151
R1511 B.n578 B.n263 10.6151
R1512 B.n579 B.n578 10.6151
R1513 B.n580 B.n579 10.6151
R1514 B.n580 B.n255 10.6151
R1515 B.n590 B.n255 10.6151
R1516 B.n591 B.n590 10.6151
R1517 B.n592 B.n591 10.6151
R1518 B.n592 B.n247 10.6151
R1519 B.n602 B.n247 10.6151
R1520 B.n603 B.n602 10.6151
R1521 B.n604 B.n603 10.6151
R1522 B.n604 B.n239 10.6151
R1523 B.n614 B.n239 10.6151
R1524 B.n615 B.n614 10.6151
R1525 B.n616 B.n615 10.6151
R1526 B.n616 B.n231 10.6151
R1527 B.n626 B.n231 10.6151
R1528 B.n627 B.n626 10.6151
R1529 B.n628 B.n627 10.6151
R1530 B.n628 B.n223 10.6151
R1531 B.n638 B.n223 10.6151
R1532 B.n639 B.n638 10.6151
R1533 B.n640 B.n639 10.6151
R1534 B.n640 B.n215 10.6151
R1535 B.n650 B.n215 10.6151
R1536 B.n651 B.n650 10.6151
R1537 B.n652 B.n651 10.6151
R1538 B.n652 B.n207 10.6151
R1539 B.n662 B.n207 10.6151
R1540 B.n663 B.n662 10.6151
R1541 B.n664 B.n663 10.6151
R1542 B.n664 B.n199 10.6151
R1543 B.n674 B.n199 10.6151
R1544 B.n675 B.n674 10.6151
R1545 B.n676 B.n675 10.6151
R1546 B.n676 B.n191 10.6151
R1547 B.n686 B.n191 10.6151
R1548 B.n687 B.n686 10.6151
R1549 B.n688 B.n687 10.6151
R1550 B.n688 B.n183 10.6151
R1551 B.n699 B.n183 10.6151
R1552 B.n700 B.n699 10.6151
R1553 B.n701 B.n700 10.6151
R1554 B.n701 B.n0 10.6151
R1555 B.n459 B.n458 10.6151
R1556 B.n458 B.n343 10.6151
R1557 B.n453 B.n343 10.6151
R1558 B.n453 B.n452 10.6151
R1559 B.n452 B.n345 10.6151
R1560 B.n447 B.n345 10.6151
R1561 B.n447 B.n446 10.6151
R1562 B.n446 B.n445 10.6151
R1563 B.n445 B.n347 10.6151
R1564 B.n439 B.n347 10.6151
R1565 B.n439 B.n438 10.6151
R1566 B.n438 B.n437 10.6151
R1567 B.n437 B.n349 10.6151
R1568 B.n431 B.n349 10.6151
R1569 B.n431 B.n430 10.6151
R1570 B.n430 B.n429 10.6151
R1571 B.n429 B.n351 10.6151
R1572 B.n423 B.n422 10.6151
R1573 B.n422 B.n421 10.6151
R1574 B.n421 B.n356 10.6151
R1575 B.n415 B.n356 10.6151
R1576 B.n415 B.n414 10.6151
R1577 B.n414 B.n413 10.6151
R1578 B.n413 B.n358 10.6151
R1579 B.n407 B.n358 10.6151
R1580 B.n407 B.n406 10.6151
R1581 B.n404 B.n362 10.6151
R1582 B.n398 B.n362 10.6151
R1583 B.n398 B.n397 10.6151
R1584 B.n397 B.n396 10.6151
R1585 B.n396 B.n364 10.6151
R1586 B.n390 B.n364 10.6151
R1587 B.n390 B.n389 10.6151
R1588 B.n389 B.n388 10.6151
R1589 B.n388 B.n366 10.6151
R1590 B.n382 B.n366 10.6151
R1591 B.n382 B.n381 10.6151
R1592 B.n381 B.n380 10.6151
R1593 B.n380 B.n368 10.6151
R1594 B.n374 B.n368 10.6151
R1595 B.n374 B.n373 10.6151
R1596 B.n373 B.n372 10.6151
R1597 B.n372 B.n339 10.6151
R1598 B.n465 B.n464 10.6151
R1599 B.n466 B.n465 10.6151
R1600 B.n466 B.n331 10.6151
R1601 B.n476 B.n331 10.6151
R1602 B.n477 B.n476 10.6151
R1603 B.n478 B.n477 10.6151
R1604 B.n478 B.n322 10.6151
R1605 B.n488 B.n322 10.6151
R1606 B.n489 B.n488 10.6151
R1607 B.n490 B.n489 10.6151
R1608 B.n490 B.n315 10.6151
R1609 B.n500 B.n315 10.6151
R1610 B.n501 B.n500 10.6151
R1611 B.n502 B.n501 10.6151
R1612 B.n502 B.n307 10.6151
R1613 B.n512 B.n307 10.6151
R1614 B.n513 B.n512 10.6151
R1615 B.n514 B.n513 10.6151
R1616 B.n514 B.n299 10.6151
R1617 B.n524 B.n299 10.6151
R1618 B.n525 B.n524 10.6151
R1619 B.n526 B.n525 10.6151
R1620 B.n526 B.n291 10.6151
R1621 B.n536 B.n291 10.6151
R1622 B.n537 B.n536 10.6151
R1623 B.n538 B.n537 10.6151
R1624 B.n538 B.n283 10.6151
R1625 B.n548 B.n283 10.6151
R1626 B.n549 B.n548 10.6151
R1627 B.n550 B.n549 10.6151
R1628 B.n550 B.n275 10.6151
R1629 B.n560 B.n275 10.6151
R1630 B.n561 B.n560 10.6151
R1631 B.n562 B.n561 10.6151
R1632 B.n562 B.n266 10.6151
R1633 B.n572 B.n266 10.6151
R1634 B.n573 B.n572 10.6151
R1635 B.n574 B.n573 10.6151
R1636 B.n574 B.n259 10.6151
R1637 B.n584 B.n259 10.6151
R1638 B.n585 B.n584 10.6151
R1639 B.n586 B.n585 10.6151
R1640 B.n586 B.n251 10.6151
R1641 B.n596 B.n251 10.6151
R1642 B.n597 B.n596 10.6151
R1643 B.n598 B.n597 10.6151
R1644 B.n598 B.n242 10.6151
R1645 B.n608 B.n242 10.6151
R1646 B.n609 B.n608 10.6151
R1647 B.n610 B.n609 10.6151
R1648 B.n610 B.n235 10.6151
R1649 B.n620 B.n235 10.6151
R1650 B.n621 B.n620 10.6151
R1651 B.n622 B.n621 10.6151
R1652 B.n622 B.n227 10.6151
R1653 B.n632 B.n227 10.6151
R1654 B.n633 B.n632 10.6151
R1655 B.n634 B.n633 10.6151
R1656 B.n634 B.n219 10.6151
R1657 B.n644 B.n219 10.6151
R1658 B.n645 B.n644 10.6151
R1659 B.n646 B.n645 10.6151
R1660 B.n646 B.n211 10.6151
R1661 B.n656 B.n211 10.6151
R1662 B.n657 B.n656 10.6151
R1663 B.n658 B.n657 10.6151
R1664 B.n658 B.n203 10.6151
R1665 B.n668 B.n203 10.6151
R1666 B.n669 B.n668 10.6151
R1667 B.n670 B.n669 10.6151
R1668 B.n670 B.n195 10.6151
R1669 B.n680 B.n195 10.6151
R1670 B.n681 B.n680 10.6151
R1671 B.n682 B.n681 10.6151
R1672 B.n682 B.n187 10.6151
R1673 B.n692 B.n187 10.6151
R1674 B.n693 B.n692 10.6151
R1675 B.n695 B.n693 10.6151
R1676 B.n695 B.n694 10.6151
R1677 B.n694 B.n179 10.6151
R1678 B.n706 B.n179 10.6151
R1679 B.n707 B.n706 10.6151
R1680 B.n708 B.n707 10.6151
R1681 B.n709 B.n708 10.6151
R1682 B.n710 B.n709 10.6151
R1683 B.n713 B.n710 10.6151
R1684 B.n714 B.n713 10.6151
R1685 B.n715 B.n714 10.6151
R1686 B.n716 B.n715 10.6151
R1687 B.n718 B.n716 10.6151
R1688 B.n719 B.n718 10.6151
R1689 B.n720 B.n719 10.6151
R1690 B.n721 B.n720 10.6151
R1691 B.n723 B.n721 10.6151
R1692 B.n724 B.n723 10.6151
R1693 B.n725 B.n724 10.6151
R1694 B.n726 B.n725 10.6151
R1695 B.n728 B.n726 10.6151
R1696 B.n729 B.n728 10.6151
R1697 B.n730 B.n729 10.6151
R1698 B.n731 B.n730 10.6151
R1699 B.n733 B.n731 10.6151
R1700 B.n734 B.n733 10.6151
R1701 B.n735 B.n734 10.6151
R1702 B.n736 B.n735 10.6151
R1703 B.n738 B.n736 10.6151
R1704 B.n739 B.n738 10.6151
R1705 B.n740 B.n739 10.6151
R1706 B.n741 B.n740 10.6151
R1707 B.n743 B.n741 10.6151
R1708 B.n744 B.n743 10.6151
R1709 B.n745 B.n744 10.6151
R1710 B.n746 B.n745 10.6151
R1711 B.n748 B.n746 10.6151
R1712 B.n749 B.n748 10.6151
R1713 B.n750 B.n749 10.6151
R1714 B.n751 B.n750 10.6151
R1715 B.n753 B.n751 10.6151
R1716 B.n754 B.n753 10.6151
R1717 B.n755 B.n754 10.6151
R1718 B.n756 B.n755 10.6151
R1719 B.n758 B.n756 10.6151
R1720 B.n759 B.n758 10.6151
R1721 B.n760 B.n759 10.6151
R1722 B.n761 B.n760 10.6151
R1723 B.n763 B.n761 10.6151
R1724 B.n764 B.n763 10.6151
R1725 B.n765 B.n764 10.6151
R1726 B.n766 B.n765 10.6151
R1727 B.n768 B.n766 10.6151
R1728 B.n769 B.n768 10.6151
R1729 B.n770 B.n769 10.6151
R1730 B.n771 B.n770 10.6151
R1731 B.n773 B.n771 10.6151
R1732 B.n774 B.n773 10.6151
R1733 B.n775 B.n774 10.6151
R1734 B.n776 B.n775 10.6151
R1735 B.n778 B.n776 10.6151
R1736 B.n779 B.n778 10.6151
R1737 B.n780 B.n779 10.6151
R1738 B.n781 B.n780 10.6151
R1739 B.n783 B.n781 10.6151
R1740 B.n784 B.n783 10.6151
R1741 B.n785 B.n784 10.6151
R1742 B.n786 B.n785 10.6151
R1743 B.n788 B.n786 10.6151
R1744 B.n789 B.n788 10.6151
R1745 B.n790 B.n789 10.6151
R1746 B.n791 B.n790 10.6151
R1747 B.n793 B.n791 10.6151
R1748 B.n794 B.n793 10.6151
R1749 B.n795 B.n794 10.6151
R1750 B.n796 B.n795 10.6151
R1751 B.n798 B.n796 10.6151
R1752 B.n799 B.n798 10.6151
R1753 B.n800 B.n799 10.6151
R1754 B.n801 B.n800 10.6151
R1755 B.n803 B.n801 10.6151
R1756 B.n804 B.n803 10.6151
R1757 B.n805 B.n804 10.6151
R1758 B.n806 B.n805 10.6151
R1759 B.n808 B.n806 10.6151
R1760 B.n809 B.n808 10.6151
R1761 B.n810 B.n809 10.6151
R1762 B.n811 B.n810 10.6151
R1763 B.n1064 B.n1 10.6151
R1764 B.n1064 B.n1063 10.6151
R1765 B.n1063 B.n1062 10.6151
R1766 B.n1062 B.n10 10.6151
R1767 B.n1056 B.n10 10.6151
R1768 B.n1056 B.n1055 10.6151
R1769 B.n1055 B.n1054 10.6151
R1770 B.n1054 B.n18 10.6151
R1771 B.n1048 B.n18 10.6151
R1772 B.n1048 B.n1047 10.6151
R1773 B.n1047 B.n1046 10.6151
R1774 B.n1046 B.n25 10.6151
R1775 B.n1040 B.n25 10.6151
R1776 B.n1040 B.n1039 10.6151
R1777 B.n1039 B.n1038 10.6151
R1778 B.n1038 B.n32 10.6151
R1779 B.n1032 B.n32 10.6151
R1780 B.n1032 B.n1031 10.6151
R1781 B.n1031 B.n1030 10.6151
R1782 B.n1030 B.n39 10.6151
R1783 B.n1024 B.n39 10.6151
R1784 B.n1024 B.n1023 10.6151
R1785 B.n1023 B.n1022 10.6151
R1786 B.n1022 B.n46 10.6151
R1787 B.n1016 B.n46 10.6151
R1788 B.n1016 B.n1015 10.6151
R1789 B.n1015 B.n1014 10.6151
R1790 B.n1014 B.n53 10.6151
R1791 B.n1008 B.n53 10.6151
R1792 B.n1008 B.n1007 10.6151
R1793 B.n1007 B.n1006 10.6151
R1794 B.n1006 B.n60 10.6151
R1795 B.n1000 B.n60 10.6151
R1796 B.n1000 B.n999 10.6151
R1797 B.n999 B.n998 10.6151
R1798 B.n998 B.n67 10.6151
R1799 B.n992 B.n67 10.6151
R1800 B.n992 B.n991 10.6151
R1801 B.n991 B.n990 10.6151
R1802 B.n990 B.n74 10.6151
R1803 B.n984 B.n74 10.6151
R1804 B.n984 B.n983 10.6151
R1805 B.n983 B.n982 10.6151
R1806 B.n982 B.n81 10.6151
R1807 B.n976 B.n81 10.6151
R1808 B.n976 B.n975 10.6151
R1809 B.n975 B.n974 10.6151
R1810 B.n974 B.n88 10.6151
R1811 B.n968 B.n88 10.6151
R1812 B.n968 B.n967 10.6151
R1813 B.n967 B.n966 10.6151
R1814 B.n966 B.n95 10.6151
R1815 B.n960 B.n95 10.6151
R1816 B.n960 B.n959 10.6151
R1817 B.n959 B.n958 10.6151
R1818 B.n958 B.n102 10.6151
R1819 B.n952 B.n102 10.6151
R1820 B.n952 B.n951 10.6151
R1821 B.n951 B.n950 10.6151
R1822 B.n950 B.n109 10.6151
R1823 B.n944 B.n109 10.6151
R1824 B.n944 B.n943 10.6151
R1825 B.n943 B.n942 10.6151
R1826 B.n942 B.n116 10.6151
R1827 B.n936 B.n116 10.6151
R1828 B.n936 B.n935 10.6151
R1829 B.n935 B.n934 10.6151
R1830 B.n934 B.n123 10.6151
R1831 B.n928 B.n123 10.6151
R1832 B.n928 B.n927 10.6151
R1833 B.n927 B.n926 10.6151
R1834 B.n926 B.n130 10.6151
R1835 B.n920 B.n130 10.6151
R1836 B.n920 B.n919 10.6151
R1837 B.n919 B.n918 10.6151
R1838 B.n918 B.n137 10.6151
R1839 B.n912 B.n137 10.6151
R1840 B.n912 B.n911 10.6151
R1841 B.n911 B.n910 10.6151
R1842 B.n910 B.n144 10.6151
R1843 B.n904 B.n144 10.6151
R1844 B.n903 B.n902 10.6151
R1845 B.n902 B.n151 10.6151
R1846 B.n896 B.n151 10.6151
R1847 B.n896 B.n895 10.6151
R1848 B.n895 B.n894 10.6151
R1849 B.n894 B.n153 10.6151
R1850 B.n888 B.n153 10.6151
R1851 B.n888 B.n887 10.6151
R1852 B.n887 B.n886 10.6151
R1853 B.n886 B.n155 10.6151
R1854 B.n880 B.n155 10.6151
R1855 B.n880 B.n879 10.6151
R1856 B.n879 B.n878 10.6151
R1857 B.n878 B.n157 10.6151
R1858 B.n872 B.n157 10.6151
R1859 B.n872 B.n871 10.6151
R1860 B.n871 B.n870 10.6151
R1861 B.n866 B.n865 10.6151
R1862 B.n865 B.n163 10.6151
R1863 B.n860 B.n163 10.6151
R1864 B.n860 B.n859 10.6151
R1865 B.n859 B.n858 10.6151
R1866 B.n858 B.n165 10.6151
R1867 B.n852 B.n165 10.6151
R1868 B.n852 B.n851 10.6151
R1869 B.n851 B.n850 10.6151
R1870 B.n846 B.n845 10.6151
R1871 B.n845 B.n171 10.6151
R1872 B.n840 B.n171 10.6151
R1873 B.n840 B.n839 10.6151
R1874 B.n839 B.n838 10.6151
R1875 B.n838 B.n173 10.6151
R1876 B.n832 B.n173 10.6151
R1877 B.n832 B.n831 10.6151
R1878 B.n831 B.n830 10.6151
R1879 B.n830 B.n175 10.6151
R1880 B.n824 B.n175 10.6151
R1881 B.n824 B.n823 10.6151
R1882 B.n823 B.n822 10.6151
R1883 B.n822 B.n177 10.6151
R1884 B.n816 B.n177 10.6151
R1885 B.n816 B.n815 10.6151
R1886 B.n815 B.n814 10.6151
R1887 B.n355 B.n351 9.36635
R1888 B.n405 B.n404 9.36635
R1889 B.n870 B.n161 9.36635
R1890 B.n846 B.n169 9.36635
R1891 B.n1072 B.n0 8.11757
R1892 B.n1072 B.n1 8.11757
R1893 B.t0 B.n289 7.09346
R1894 B.n955 B.t5 7.09346
R1895 B.n423 B.n355 1.24928
R1896 B.n406 B.n405 1.24928
R1897 B.n866 B.n161 1.24928
R1898 B.n850 B.n169 1.24928
R1899 VP.n32 VP.n29 161.3
R1900 VP.n34 VP.n33 161.3
R1901 VP.n35 VP.n28 161.3
R1902 VP.n37 VP.n36 161.3
R1903 VP.n38 VP.n27 161.3
R1904 VP.n40 VP.n39 161.3
R1905 VP.n41 VP.n26 161.3
R1906 VP.n43 VP.n42 161.3
R1907 VP.n44 VP.n25 161.3
R1908 VP.n46 VP.n45 161.3
R1909 VP.n47 VP.n24 161.3
R1910 VP.n49 VP.n48 161.3
R1911 VP.n50 VP.n23 161.3
R1912 VP.n52 VP.n51 161.3
R1913 VP.n53 VP.n22 161.3
R1914 VP.n55 VP.n54 161.3
R1915 VP.n56 VP.n21 161.3
R1916 VP.n59 VP.n58 161.3
R1917 VP.n60 VP.n20 161.3
R1918 VP.n62 VP.n61 161.3
R1919 VP.n63 VP.n19 161.3
R1920 VP.n65 VP.n64 161.3
R1921 VP.n66 VP.n18 161.3
R1922 VP.n68 VP.n67 161.3
R1923 VP.n69 VP.n17 161.3
R1924 VP.n124 VP.n0 161.3
R1925 VP.n123 VP.n122 161.3
R1926 VP.n121 VP.n1 161.3
R1927 VP.n120 VP.n119 161.3
R1928 VP.n118 VP.n2 161.3
R1929 VP.n117 VP.n116 161.3
R1930 VP.n115 VP.n3 161.3
R1931 VP.n114 VP.n113 161.3
R1932 VP.n111 VP.n4 161.3
R1933 VP.n110 VP.n109 161.3
R1934 VP.n108 VP.n5 161.3
R1935 VP.n107 VP.n106 161.3
R1936 VP.n105 VP.n6 161.3
R1937 VP.n104 VP.n103 161.3
R1938 VP.n102 VP.n7 161.3
R1939 VP.n101 VP.n100 161.3
R1940 VP.n99 VP.n8 161.3
R1941 VP.n98 VP.n97 161.3
R1942 VP.n96 VP.n9 161.3
R1943 VP.n95 VP.n94 161.3
R1944 VP.n93 VP.n10 161.3
R1945 VP.n92 VP.n91 161.3
R1946 VP.n90 VP.n11 161.3
R1947 VP.n89 VP.n88 161.3
R1948 VP.n87 VP.n12 161.3
R1949 VP.n85 VP.n84 161.3
R1950 VP.n83 VP.n13 161.3
R1951 VP.n82 VP.n81 161.3
R1952 VP.n80 VP.n14 161.3
R1953 VP.n79 VP.n78 161.3
R1954 VP.n77 VP.n15 161.3
R1955 VP.n76 VP.n75 161.3
R1956 VP.n74 VP.n16 161.3
R1957 VP.n31 VP.n30 63.8768
R1958 VP.n73 VP.n72 59.6721
R1959 VP.n126 VP.n125 59.6721
R1960 VP.n71 VP.n70 59.6721
R1961 VP.n30 VP.t3 57.043
R1962 VP.n80 VP.n79 55.548
R1963 VP.n119 VP.n118 55.548
R1964 VP.n64 VP.n63 55.548
R1965 VP.n72 VP.n71 54.4017
R1966 VP.n93 VP.n92 51.663
R1967 VP.n106 VP.n105 51.663
R1968 VP.n51 VP.n50 51.663
R1969 VP.n38 VP.n37 51.663
R1970 VP.n94 VP.n93 29.3238
R1971 VP.n105 VP.n104 29.3238
R1972 VP.n50 VP.n49 29.3238
R1973 VP.n39 VP.n38 29.3238
R1974 VP.n79 VP.n15 25.4388
R1975 VP.n119 VP.n1 25.4388
R1976 VP.n64 VP.n18 25.4388
R1977 VP.n99 VP.t5 24.9038
R1978 VP.n73 VP.t4 24.9038
R1979 VP.n86 VP.t9 24.9038
R1980 VP.n112 VP.t2 24.9038
R1981 VP.n125 VP.t8 24.9038
R1982 VP.n44 VP.t6 24.9038
R1983 VP.n70 VP.t7 24.9038
R1984 VP.n57 VP.t1 24.9038
R1985 VP.n31 VP.t0 24.9038
R1986 VP.n75 VP.n74 24.4675
R1987 VP.n75 VP.n15 24.4675
R1988 VP.n81 VP.n80 24.4675
R1989 VP.n81 VP.n13 24.4675
R1990 VP.n85 VP.n13 24.4675
R1991 VP.n88 VP.n87 24.4675
R1992 VP.n88 VP.n11 24.4675
R1993 VP.n92 VP.n11 24.4675
R1994 VP.n94 VP.n9 24.4675
R1995 VP.n98 VP.n9 24.4675
R1996 VP.n99 VP.n98 24.4675
R1997 VP.n100 VP.n99 24.4675
R1998 VP.n100 VP.n7 24.4675
R1999 VP.n104 VP.n7 24.4675
R2000 VP.n106 VP.n5 24.4675
R2001 VP.n110 VP.n5 24.4675
R2002 VP.n111 VP.n110 24.4675
R2003 VP.n113 VP.n3 24.4675
R2004 VP.n117 VP.n3 24.4675
R2005 VP.n118 VP.n117 24.4675
R2006 VP.n123 VP.n1 24.4675
R2007 VP.n124 VP.n123 24.4675
R2008 VP.n68 VP.n18 24.4675
R2009 VP.n69 VP.n68 24.4675
R2010 VP.n51 VP.n22 24.4675
R2011 VP.n55 VP.n22 24.4675
R2012 VP.n56 VP.n55 24.4675
R2013 VP.n58 VP.n20 24.4675
R2014 VP.n62 VP.n20 24.4675
R2015 VP.n63 VP.n62 24.4675
R2016 VP.n39 VP.n26 24.4675
R2017 VP.n43 VP.n26 24.4675
R2018 VP.n44 VP.n43 24.4675
R2019 VP.n45 VP.n44 24.4675
R2020 VP.n45 VP.n24 24.4675
R2021 VP.n49 VP.n24 24.4675
R2022 VP.n33 VP.n32 24.4675
R2023 VP.n33 VP.n28 24.4675
R2024 VP.n37 VP.n28 24.4675
R2025 VP.n74 VP.n73 22.5101
R2026 VP.n125 VP.n124 22.5101
R2027 VP.n70 VP.n69 22.5101
R2028 VP.n86 VP.n85 13.2127
R2029 VP.n113 VP.n112 13.2127
R2030 VP.n58 VP.n57 13.2127
R2031 VP.n87 VP.n86 11.2553
R2032 VP.n112 VP.n111 11.2553
R2033 VP.n57 VP.n56 11.2553
R2034 VP.n32 VP.n31 11.2553
R2035 VP.n30 VP.n29 2.60578
R2036 VP.n71 VP.n17 0.417535
R2037 VP.n72 VP.n16 0.417535
R2038 VP.n126 VP.n0 0.417535
R2039 VP VP.n126 0.394291
R2040 VP.n34 VP.n29 0.189894
R2041 VP.n35 VP.n34 0.189894
R2042 VP.n36 VP.n35 0.189894
R2043 VP.n36 VP.n27 0.189894
R2044 VP.n40 VP.n27 0.189894
R2045 VP.n41 VP.n40 0.189894
R2046 VP.n42 VP.n41 0.189894
R2047 VP.n42 VP.n25 0.189894
R2048 VP.n46 VP.n25 0.189894
R2049 VP.n47 VP.n46 0.189894
R2050 VP.n48 VP.n47 0.189894
R2051 VP.n48 VP.n23 0.189894
R2052 VP.n52 VP.n23 0.189894
R2053 VP.n53 VP.n52 0.189894
R2054 VP.n54 VP.n53 0.189894
R2055 VP.n54 VP.n21 0.189894
R2056 VP.n59 VP.n21 0.189894
R2057 VP.n60 VP.n59 0.189894
R2058 VP.n61 VP.n60 0.189894
R2059 VP.n61 VP.n19 0.189894
R2060 VP.n65 VP.n19 0.189894
R2061 VP.n66 VP.n65 0.189894
R2062 VP.n67 VP.n66 0.189894
R2063 VP.n67 VP.n17 0.189894
R2064 VP.n76 VP.n16 0.189894
R2065 VP.n77 VP.n76 0.189894
R2066 VP.n78 VP.n77 0.189894
R2067 VP.n78 VP.n14 0.189894
R2068 VP.n82 VP.n14 0.189894
R2069 VP.n83 VP.n82 0.189894
R2070 VP.n84 VP.n83 0.189894
R2071 VP.n84 VP.n12 0.189894
R2072 VP.n89 VP.n12 0.189894
R2073 VP.n90 VP.n89 0.189894
R2074 VP.n91 VP.n90 0.189894
R2075 VP.n91 VP.n10 0.189894
R2076 VP.n95 VP.n10 0.189894
R2077 VP.n96 VP.n95 0.189894
R2078 VP.n97 VP.n96 0.189894
R2079 VP.n97 VP.n8 0.189894
R2080 VP.n101 VP.n8 0.189894
R2081 VP.n102 VP.n101 0.189894
R2082 VP.n103 VP.n102 0.189894
R2083 VP.n103 VP.n6 0.189894
R2084 VP.n107 VP.n6 0.189894
R2085 VP.n108 VP.n107 0.189894
R2086 VP.n109 VP.n108 0.189894
R2087 VP.n109 VP.n4 0.189894
R2088 VP.n114 VP.n4 0.189894
R2089 VP.n115 VP.n114 0.189894
R2090 VP.n116 VP.n115 0.189894
R2091 VP.n116 VP.n2 0.189894
R2092 VP.n120 VP.n2 0.189894
R2093 VP.n121 VP.n120 0.189894
R2094 VP.n122 VP.n121 0.189894
R2095 VP.n122 VP.n0 0.189894
R2096 VDD1.n14 VDD1.n0 289.615
R2097 VDD1.n35 VDD1.n21 289.615
R2098 VDD1.n15 VDD1.n14 185
R2099 VDD1.n13 VDD1.n12 185
R2100 VDD1.n4 VDD1.n3 185
R2101 VDD1.n7 VDD1.n6 185
R2102 VDD1.n28 VDD1.n27 185
R2103 VDD1.n25 VDD1.n24 185
R2104 VDD1.n34 VDD1.n33 185
R2105 VDD1.n36 VDD1.n35 185
R2106 VDD1.t6 VDD1.n5 147.888
R2107 VDD1.t5 VDD1.n26 147.888
R2108 VDD1.n14 VDD1.n13 104.615
R2109 VDD1.n13 VDD1.n3 104.615
R2110 VDD1.n6 VDD1.n3 104.615
R2111 VDD1.n27 VDD1.n24 104.615
R2112 VDD1.n34 VDD1.n24 104.615
R2113 VDD1.n35 VDD1.n34 104.615
R2114 VDD1.n43 VDD1.n42 79.8284
R2115 VDD1.n20 VDD1.n19 77.149
R2116 VDD1.n45 VDD1.n44 77.1488
R2117 VDD1.n41 VDD1.n40 77.1488
R2118 VDD1.n20 VDD1.n18 56.1955
R2119 VDD1.n41 VDD1.n39 56.1955
R2120 VDD1.n6 VDD1.t6 52.3082
R2121 VDD1.n27 VDD1.t5 52.3082
R2122 VDD1.n45 VDD1.n43 46.9168
R2123 VDD1.n7 VDD1.n5 15.6496
R2124 VDD1.n28 VDD1.n26 15.6496
R2125 VDD1.n8 VDD1.n4 12.8005
R2126 VDD1.n29 VDD1.n25 12.8005
R2127 VDD1.n12 VDD1.n11 12.0247
R2128 VDD1.n33 VDD1.n32 12.0247
R2129 VDD1.n15 VDD1.n2 11.249
R2130 VDD1.n36 VDD1.n23 11.249
R2131 VDD1.n16 VDD1.n0 10.4732
R2132 VDD1.n37 VDD1.n21 10.4732
R2133 VDD1.n18 VDD1.n17 9.45567
R2134 VDD1.n39 VDD1.n38 9.45567
R2135 VDD1.n17 VDD1.n16 9.3005
R2136 VDD1.n2 VDD1.n1 9.3005
R2137 VDD1.n11 VDD1.n10 9.3005
R2138 VDD1.n9 VDD1.n8 9.3005
R2139 VDD1.n38 VDD1.n37 9.3005
R2140 VDD1.n23 VDD1.n22 9.3005
R2141 VDD1.n32 VDD1.n31 9.3005
R2142 VDD1.n30 VDD1.n29 9.3005
R2143 VDD1.n44 VDD1.t8 4.91365
R2144 VDD1.n44 VDD1.t2 4.91365
R2145 VDD1.n19 VDD1.t0 4.91365
R2146 VDD1.n19 VDD1.t7 4.91365
R2147 VDD1.n42 VDD1.t9 4.91365
R2148 VDD1.n42 VDD1.t4 4.91365
R2149 VDD1.n40 VDD1.t3 4.91365
R2150 VDD1.n40 VDD1.t1 4.91365
R2151 VDD1.n9 VDD1.n5 4.40546
R2152 VDD1.n30 VDD1.n26 4.40546
R2153 VDD1.n18 VDD1.n0 3.49141
R2154 VDD1.n39 VDD1.n21 3.49141
R2155 VDD1.n16 VDD1.n15 2.71565
R2156 VDD1.n37 VDD1.n36 2.71565
R2157 VDD1 VDD1.n45 2.67722
R2158 VDD1.n12 VDD1.n2 1.93989
R2159 VDD1.n33 VDD1.n23 1.93989
R2160 VDD1.n11 VDD1.n4 1.16414
R2161 VDD1.n32 VDD1.n25 1.16414
R2162 VDD1 VDD1.n20 0.970328
R2163 VDD1.n43 VDD1.n41 0.856792
R2164 VDD1.n8 VDD1.n7 0.388379
R2165 VDD1.n29 VDD1.n28 0.388379
R2166 VDD1.n17 VDD1.n1 0.155672
R2167 VDD1.n10 VDD1.n1 0.155672
R2168 VDD1.n10 VDD1.n9 0.155672
R2169 VDD1.n31 VDD1.n30 0.155672
R2170 VDD1.n31 VDD1.n22 0.155672
R2171 VDD1.n38 VDD1.n22 0.155672
R2172 VTAIL.n88 VTAIL.n74 289.615
R2173 VTAIL.n16 VTAIL.n2 289.615
R2174 VTAIL.n68 VTAIL.n54 289.615
R2175 VTAIL.n44 VTAIL.n30 289.615
R2176 VTAIL.n81 VTAIL.n80 185
R2177 VTAIL.n78 VTAIL.n77 185
R2178 VTAIL.n87 VTAIL.n86 185
R2179 VTAIL.n89 VTAIL.n88 185
R2180 VTAIL.n9 VTAIL.n8 185
R2181 VTAIL.n6 VTAIL.n5 185
R2182 VTAIL.n15 VTAIL.n14 185
R2183 VTAIL.n17 VTAIL.n16 185
R2184 VTAIL.n69 VTAIL.n68 185
R2185 VTAIL.n67 VTAIL.n66 185
R2186 VTAIL.n58 VTAIL.n57 185
R2187 VTAIL.n61 VTAIL.n60 185
R2188 VTAIL.n45 VTAIL.n44 185
R2189 VTAIL.n43 VTAIL.n42 185
R2190 VTAIL.n34 VTAIL.n33 185
R2191 VTAIL.n37 VTAIL.n36 185
R2192 VTAIL.t1 VTAIL.n79 147.888
R2193 VTAIL.t10 VTAIL.n7 147.888
R2194 VTAIL.t11 VTAIL.n59 147.888
R2195 VTAIL.t4 VTAIL.n35 147.888
R2196 VTAIL.n80 VTAIL.n77 104.615
R2197 VTAIL.n87 VTAIL.n77 104.615
R2198 VTAIL.n88 VTAIL.n87 104.615
R2199 VTAIL.n8 VTAIL.n5 104.615
R2200 VTAIL.n15 VTAIL.n5 104.615
R2201 VTAIL.n16 VTAIL.n15 104.615
R2202 VTAIL.n68 VTAIL.n67 104.615
R2203 VTAIL.n67 VTAIL.n57 104.615
R2204 VTAIL.n60 VTAIL.n57 104.615
R2205 VTAIL.n44 VTAIL.n43 104.615
R2206 VTAIL.n43 VTAIL.n33 104.615
R2207 VTAIL.n36 VTAIL.n33 104.615
R2208 VTAIL.n53 VTAIL.n52 60.4702
R2209 VTAIL.n51 VTAIL.n50 60.4702
R2210 VTAIL.n29 VTAIL.n28 60.4702
R2211 VTAIL.n27 VTAIL.n26 60.4702
R2212 VTAIL.n95 VTAIL.n94 60.47
R2213 VTAIL.n1 VTAIL.n0 60.47
R2214 VTAIL.n23 VTAIL.n22 60.47
R2215 VTAIL.n25 VTAIL.n24 60.47
R2216 VTAIL.n80 VTAIL.t1 52.3082
R2217 VTAIL.n8 VTAIL.t10 52.3082
R2218 VTAIL.n60 VTAIL.t11 52.3082
R2219 VTAIL.n36 VTAIL.t4 52.3082
R2220 VTAIL.n93 VTAIL.n92 35.8702
R2221 VTAIL.n21 VTAIL.n20 35.8702
R2222 VTAIL.n73 VTAIL.n72 35.8702
R2223 VTAIL.n49 VTAIL.n48 35.8702
R2224 VTAIL.n27 VTAIL.n25 23.1341
R2225 VTAIL.n93 VTAIL.n73 19.4876
R2226 VTAIL.n81 VTAIL.n79 15.6496
R2227 VTAIL.n9 VTAIL.n7 15.6496
R2228 VTAIL.n61 VTAIL.n59 15.6496
R2229 VTAIL.n37 VTAIL.n35 15.6496
R2230 VTAIL.n82 VTAIL.n78 12.8005
R2231 VTAIL.n10 VTAIL.n6 12.8005
R2232 VTAIL.n62 VTAIL.n58 12.8005
R2233 VTAIL.n38 VTAIL.n34 12.8005
R2234 VTAIL.n86 VTAIL.n85 12.0247
R2235 VTAIL.n14 VTAIL.n13 12.0247
R2236 VTAIL.n66 VTAIL.n65 12.0247
R2237 VTAIL.n42 VTAIL.n41 12.0247
R2238 VTAIL.n89 VTAIL.n76 11.249
R2239 VTAIL.n17 VTAIL.n4 11.249
R2240 VTAIL.n69 VTAIL.n56 11.249
R2241 VTAIL.n45 VTAIL.n32 11.249
R2242 VTAIL.n90 VTAIL.n74 10.4732
R2243 VTAIL.n18 VTAIL.n2 10.4732
R2244 VTAIL.n70 VTAIL.n54 10.4732
R2245 VTAIL.n46 VTAIL.n30 10.4732
R2246 VTAIL.n92 VTAIL.n91 9.45567
R2247 VTAIL.n20 VTAIL.n19 9.45567
R2248 VTAIL.n72 VTAIL.n71 9.45567
R2249 VTAIL.n48 VTAIL.n47 9.45567
R2250 VTAIL.n91 VTAIL.n90 9.3005
R2251 VTAIL.n76 VTAIL.n75 9.3005
R2252 VTAIL.n85 VTAIL.n84 9.3005
R2253 VTAIL.n83 VTAIL.n82 9.3005
R2254 VTAIL.n19 VTAIL.n18 9.3005
R2255 VTAIL.n4 VTAIL.n3 9.3005
R2256 VTAIL.n13 VTAIL.n12 9.3005
R2257 VTAIL.n11 VTAIL.n10 9.3005
R2258 VTAIL.n71 VTAIL.n70 9.3005
R2259 VTAIL.n56 VTAIL.n55 9.3005
R2260 VTAIL.n65 VTAIL.n64 9.3005
R2261 VTAIL.n63 VTAIL.n62 9.3005
R2262 VTAIL.n47 VTAIL.n46 9.3005
R2263 VTAIL.n32 VTAIL.n31 9.3005
R2264 VTAIL.n41 VTAIL.n40 9.3005
R2265 VTAIL.n39 VTAIL.n38 9.3005
R2266 VTAIL.n94 VTAIL.t6 4.91365
R2267 VTAIL.n94 VTAIL.t8 4.91365
R2268 VTAIL.n0 VTAIL.t5 4.91365
R2269 VTAIL.n0 VTAIL.t19 4.91365
R2270 VTAIL.n22 VTAIL.t13 4.91365
R2271 VTAIL.n22 VTAIL.t16 4.91365
R2272 VTAIL.n24 VTAIL.t14 4.91365
R2273 VTAIL.n24 VTAIL.t9 4.91365
R2274 VTAIL.n52 VTAIL.t12 4.91365
R2275 VTAIL.n52 VTAIL.t17 4.91365
R2276 VTAIL.n50 VTAIL.t15 4.91365
R2277 VTAIL.n50 VTAIL.t18 4.91365
R2278 VTAIL.n28 VTAIL.t3 4.91365
R2279 VTAIL.n28 VTAIL.t7 4.91365
R2280 VTAIL.n26 VTAIL.t0 4.91365
R2281 VTAIL.n26 VTAIL.t2 4.91365
R2282 VTAIL.n83 VTAIL.n79 4.40546
R2283 VTAIL.n11 VTAIL.n7 4.40546
R2284 VTAIL.n63 VTAIL.n59 4.40546
R2285 VTAIL.n39 VTAIL.n35 4.40546
R2286 VTAIL.n29 VTAIL.n27 3.64705
R2287 VTAIL.n49 VTAIL.n29 3.64705
R2288 VTAIL.n53 VTAIL.n51 3.64705
R2289 VTAIL.n73 VTAIL.n53 3.64705
R2290 VTAIL.n25 VTAIL.n23 3.64705
R2291 VTAIL.n23 VTAIL.n21 3.64705
R2292 VTAIL.n95 VTAIL.n93 3.64705
R2293 VTAIL.n92 VTAIL.n74 3.49141
R2294 VTAIL.n20 VTAIL.n2 3.49141
R2295 VTAIL.n72 VTAIL.n54 3.49141
R2296 VTAIL.n48 VTAIL.n30 3.49141
R2297 VTAIL VTAIL.n1 2.7936
R2298 VTAIL.n90 VTAIL.n89 2.71565
R2299 VTAIL.n18 VTAIL.n17 2.71565
R2300 VTAIL.n70 VTAIL.n69 2.71565
R2301 VTAIL.n46 VTAIL.n45 2.71565
R2302 VTAIL.n51 VTAIL.n49 2.2936
R2303 VTAIL.n21 VTAIL.n1 2.2936
R2304 VTAIL.n86 VTAIL.n76 1.93989
R2305 VTAIL.n14 VTAIL.n4 1.93989
R2306 VTAIL.n66 VTAIL.n56 1.93989
R2307 VTAIL.n42 VTAIL.n32 1.93989
R2308 VTAIL.n85 VTAIL.n78 1.16414
R2309 VTAIL.n13 VTAIL.n6 1.16414
R2310 VTAIL.n65 VTAIL.n58 1.16414
R2311 VTAIL.n41 VTAIL.n34 1.16414
R2312 VTAIL VTAIL.n95 0.853948
R2313 VTAIL.n82 VTAIL.n81 0.388379
R2314 VTAIL.n10 VTAIL.n9 0.388379
R2315 VTAIL.n62 VTAIL.n61 0.388379
R2316 VTAIL.n38 VTAIL.n37 0.388379
R2317 VTAIL.n84 VTAIL.n83 0.155672
R2318 VTAIL.n84 VTAIL.n75 0.155672
R2319 VTAIL.n91 VTAIL.n75 0.155672
R2320 VTAIL.n12 VTAIL.n11 0.155672
R2321 VTAIL.n12 VTAIL.n3 0.155672
R2322 VTAIL.n19 VTAIL.n3 0.155672
R2323 VTAIL.n71 VTAIL.n55 0.155672
R2324 VTAIL.n64 VTAIL.n55 0.155672
R2325 VTAIL.n64 VTAIL.n63 0.155672
R2326 VTAIL.n47 VTAIL.n31 0.155672
R2327 VTAIL.n40 VTAIL.n31 0.155672
R2328 VTAIL.n40 VTAIL.n39 0.155672
R2329 VN.n107 VN.n55 161.3
R2330 VN.n106 VN.n105 161.3
R2331 VN.n104 VN.n56 161.3
R2332 VN.n103 VN.n102 161.3
R2333 VN.n101 VN.n57 161.3
R2334 VN.n100 VN.n99 161.3
R2335 VN.n98 VN.n58 161.3
R2336 VN.n97 VN.n96 161.3
R2337 VN.n94 VN.n59 161.3
R2338 VN.n93 VN.n92 161.3
R2339 VN.n91 VN.n60 161.3
R2340 VN.n90 VN.n89 161.3
R2341 VN.n88 VN.n61 161.3
R2342 VN.n87 VN.n86 161.3
R2343 VN.n85 VN.n62 161.3
R2344 VN.n84 VN.n83 161.3
R2345 VN.n82 VN.n63 161.3
R2346 VN.n81 VN.n80 161.3
R2347 VN.n79 VN.n64 161.3
R2348 VN.n78 VN.n77 161.3
R2349 VN.n76 VN.n65 161.3
R2350 VN.n75 VN.n74 161.3
R2351 VN.n73 VN.n66 161.3
R2352 VN.n72 VN.n71 161.3
R2353 VN.n70 VN.n67 161.3
R2354 VN.n52 VN.n0 161.3
R2355 VN.n51 VN.n50 161.3
R2356 VN.n49 VN.n1 161.3
R2357 VN.n48 VN.n47 161.3
R2358 VN.n46 VN.n2 161.3
R2359 VN.n45 VN.n44 161.3
R2360 VN.n43 VN.n3 161.3
R2361 VN.n42 VN.n41 161.3
R2362 VN.n39 VN.n4 161.3
R2363 VN.n38 VN.n37 161.3
R2364 VN.n36 VN.n5 161.3
R2365 VN.n35 VN.n34 161.3
R2366 VN.n33 VN.n6 161.3
R2367 VN.n32 VN.n31 161.3
R2368 VN.n30 VN.n7 161.3
R2369 VN.n29 VN.n28 161.3
R2370 VN.n27 VN.n8 161.3
R2371 VN.n26 VN.n25 161.3
R2372 VN.n24 VN.n9 161.3
R2373 VN.n23 VN.n22 161.3
R2374 VN.n21 VN.n10 161.3
R2375 VN.n20 VN.n19 161.3
R2376 VN.n18 VN.n11 161.3
R2377 VN.n17 VN.n16 161.3
R2378 VN.n15 VN.n12 161.3
R2379 VN.n14 VN.n13 63.8768
R2380 VN.n69 VN.n68 63.8768
R2381 VN.n54 VN.n53 59.6721
R2382 VN.n109 VN.n108 59.6721
R2383 VN.n13 VN.t9 57.0435
R2384 VN.n68 VN.t6 57.0435
R2385 VN.n47 VN.n46 55.548
R2386 VN.n102 VN.n101 55.548
R2387 VN VN.n109 54.4397
R2388 VN.n21 VN.n20 51.663
R2389 VN.n34 VN.n33 51.663
R2390 VN.n76 VN.n75 51.663
R2391 VN.n89 VN.n88 51.663
R2392 VN.n22 VN.n21 29.3238
R2393 VN.n33 VN.n32 29.3238
R2394 VN.n77 VN.n76 29.3238
R2395 VN.n88 VN.n87 29.3238
R2396 VN.n47 VN.n1 25.4388
R2397 VN.n102 VN.n56 25.4388
R2398 VN.n27 VN.t8 24.9038
R2399 VN.n14 VN.t4 24.9038
R2400 VN.n40 VN.t2 24.9038
R2401 VN.n53 VN.t7 24.9038
R2402 VN.n82 VN.t0 24.9038
R2403 VN.n69 VN.t3 24.9038
R2404 VN.n95 VN.t5 24.9038
R2405 VN.n108 VN.t1 24.9038
R2406 VN.n16 VN.n15 24.4675
R2407 VN.n16 VN.n11 24.4675
R2408 VN.n20 VN.n11 24.4675
R2409 VN.n22 VN.n9 24.4675
R2410 VN.n26 VN.n9 24.4675
R2411 VN.n27 VN.n26 24.4675
R2412 VN.n28 VN.n27 24.4675
R2413 VN.n28 VN.n7 24.4675
R2414 VN.n32 VN.n7 24.4675
R2415 VN.n34 VN.n5 24.4675
R2416 VN.n38 VN.n5 24.4675
R2417 VN.n39 VN.n38 24.4675
R2418 VN.n41 VN.n3 24.4675
R2419 VN.n45 VN.n3 24.4675
R2420 VN.n46 VN.n45 24.4675
R2421 VN.n51 VN.n1 24.4675
R2422 VN.n52 VN.n51 24.4675
R2423 VN.n75 VN.n66 24.4675
R2424 VN.n71 VN.n66 24.4675
R2425 VN.n71 VN.n70 24.4675
R2426 VN.n87 VN.n62 24.4675
R2427 VN.n83 VN.n62 24.4675
R2428 VN.n83 VN.n82 24.4675
R2429 VN.n82 VN.n81 24.4675
R2430 VN.n81 VN.n64 24.4675
R2431 VN.n77 VN.n64 24.4675
R2432 VN.n101 VN.n100 24.4675
R2433 VN.n100 VN.n58 24.4675
R2434 VN.n96 VN.n58 24.4675
R2435 VN.n94 VN.n93 24.4675
R2436 VN.n93 VN.n60 24.4675
R2437 VN.n89 VN.n60 24.4675
R2438 VN.n107 VN.n106 24.4675
R2439 VN.n106 VN.n56 24.4675
R2440 VN.n53 VN.n52 22.5101
R2441 VN.n108 VN.n107 22.5101
R2442 VN.n41 VN.n40 13.2127
R2443 VN.n96 VN.n95 13.2127
R2444 VN.n15 VN.n14 11.2553
R2445 VN.n40 VN.n39 11.2553
R2446 VN.n70 VN.n69 11.2553
R2447 VN.n95 VN.n94 11.2553
R2448 VN.n68 VN.n67 2.6058
R2449 VN.n13 VN.n12 2.6058
R2450 VN.n109 VN.n55 0.417535
R2451 VN.n54 VN.n0 0.417535
R2452 VN VN.n54 0.394291
R2453 VN.n105 VN.n55 0.189894
R2454 VN.n105 VN.n104 0.189894
R2455 VN.n104 VN.n103 0.189894
R2456 VN.n103 VN.n57 0.189894
R2457 VN.n99 VN.n57 0.189894
R2458 VN.n99 VN.n98 0.189894
R2459 VN.n98 VN.n97 0.189894
R2460 VN.n97 VN.n59 0.189894
R2461 VN.n92 VN.n59 0.189894
R2462 VN.n92 VN.n91 0.189894
R2463 VN.n91 VN.n90 0.189894
R2464 VN.n90 VN.n61 0.189894
R2465 VN.n86 VN.n61 0.189894
R2466 VN.n86 VN.n85 0.189894
R2467 VN.n85 VN.n84 0.189894
R2468 VN.n84 VN.n63 0.189894
R2469 VN.n80 VN.n63 0.189894
R2470 VN.n80 VN.n79 0.189894
R2471 VN.n79 VN.n78 0.189894
R2472 VN.n78 VN.n65 0.189894
R2473 VN.n74 VN.n65 0.189894
R2474 VN.n74 VN.n73 0.189894
R2475 VN.n73 VN.n72 0.189894
R2476 VN.n72 VN.n67 0.189894
R2477 VN.n17 VN.n12 0.189894
R2478 VN.n18 VN.n17 0.189894
R2479 VN.n19 VN.n18 0.189894
R2480 VN.n19 VN.n10 0.189894
R2481 VN.n23 VN.n10 0.189894
R2482 VN.n24 VN.n23 0.189894
R2483 VN.n25 VN.n24 0.189894
R2484 VN.n25 VN.n8 0.189894
R2485 VN.n29 VN.n8 0.189894
R2486 VN.n30 VN.n29 0.189894
R2487 VN.n31 VN.n30 0.189894
R2488 VN.n31 VN.n6 0.189894
R2489 VN.n35 VN.n6 0.189894
R2490 VN.n36 VN.n35 0.189894
R2491 VN.n37 VN.n36 0.189894
R2492 VN.n37 VN.n4 0.189894
R2493 VN.n42 VN.n4 0.189894
R2494 VN.n43 VN.n42 0.189894
R2495 VN.n44 VN.n43 0.189894
R2496 VN.n44 VN.n2 0.189894
R2497 VN.n48 VN.n2 0.189894
R2498 VN.n49 VN.n48 0.189894
R2499 VN.n50 VN.n49 0.189894
R2500 VN.n50 VN.n0 0.189894
R2501 VDD2.n37 VDD2.n23 289.615
R2502 VDD2.n14 VDD2.n0 289.615
R2503 VDD2.n38 VDD2.n37 185
R2504 VDD2.n36 VDD2.n35 185
R2505 VDD2.n27 VDD2.n26 185
R2506 VDD2.n30 VDD2.n29 185
R2507 VDD2.n7 VDD2.n6 185
R2508 VDD2.n4 VDD2.n3 185
R2509 VDD2.n13 VDD2.n12 185
R2510 VDD2.n15 VDD2.n14 185
R2511 VDD2.t8 VDD2.n28 147.888
R2512 VDD2.t0 VDD2.n5 147.888
R2513 VDD2.n37 VDD2.n36 104.615
R2514 VDD2.n36 VDD2.n26 104.615
R2515 VDD2.n29 VDD2.n26 104.615
R2516 VDD2.n6 VDD2.n3 104.615
R2517 VDD2.n13 VDD2.n3 104.615
R2518 VDD2.n14 VDD2.n13 104.615
R2519 VDD2.n22 VDD2.n21 79.8284
R2520 VDD2 VDD2.n45 79.8256
R2521 VDD2.n44 VDD2.n43 77.149
R2522 VDD2.n20 VDD2.n19 77.1488
R2523 VDD2.n20 VDD2.n18 56.1955
R2524 VDD2.n42 VDD2.n41 52.549
R2525 VDD2.n29 VDD2.t8 52.3082
R2526 VDD2.n6 VDD2.t0 52.3082
R2527 VDD2.n42 VDD2.n22 44.5106
R2528 VDD2.n30 VDD2.n28 15.6496
R2529 VDD2.n7 VDD2.n5 15.6496
R2530 VDD2.n31 VDD2.n27 12.8005
R2531 VDD2.n8 VDD2.n4 12.8005
R2532 VDD2.n35 VDD2.n34 12.0247
R2533 VDD2.n12 VDD2.n11 12.0247
R2534 VDD2.n38 VDD2.n25 11.249
R2535 VDD2.n15 VDD2.n2 11.249
R2536 VDD2.n39 VDD2.n23 10.4732
R2537 VDD2.n16 VDD2.n0 10.4732
R2538 VDD2.n41 VDD2.n40 9.45567
R2539 VDD2.n18 VDD2.n17 9.45567
R2540 VDD2.n40 VDD2.n39 9.3005
R2541 VDD2.n25 VDD2.n24 9.3005
R2542 VDD2.n34 VDD2.n33 9.3005
R2543 VDD2.n32 VDD2.n31 9.3005
R2544 VDD2.n17 VDD2.n16 9.3005
R2545 VDD2.n2 VDD2.n1 9.3005
R2546 VDD2.n11 VDD2.n10 9.3005
R2547 VDD2.n9 VDD2.n8 9.3005
R2548 VDD2.n45 VDD2.t6 4.91365
R2549 VDD2.n45 VDD2.t3 4.91365
R2550 VDD2.n43 VDD2.t4 4.91365
R2551 VDD2.n43 VDD2.t9 4.91365
R2552 VDD2.n21 VDD2.t7 4.91365
R2553 VDD2.n21 VDD2.t2 4.91365
R2554 VDD2.n19 VDD2.t5 4.91365
R2555 VDD2.n19 VDD2.t1 4.91365
R2556 VDD2.n32 VDD2.n28 4.40546
R2557 VDD2.n9 VDD2.n5 4.40546
R2558 VDD2.n44 VDD2.n42 3.64705
R2559 VDD2.n41 VDD2.n23 3.49141
R2560 VDD2.n18 VDD2.n0 3.49141
R2561 VDD2.n39 VDD2.n38 2.71565
R2562 VDD2.n16 VDD2.n15 2.71565
R2563 VDD2.n35 VDD2.n25 1.93989
R2564 VDD2.n12 VDD2.n2 1.93989
R2565 VDD2.n34 VDD2.n27 1.16414
R2566 VDD2.n11 VDD2.n4 1.16414
R2567 VDD2 VDD2.n44 0.970328
R2568 VDD2.n22 VDD2.n20 0.856792
R2569 VDD2.n31 VDD2.n30 0.388379
R2570 VDD2.n8 VDD2.n7 0.388379
R2571 VDD2.n40 VDD2.n24 0.155672
R2572 VDD2.n33 VDD2.n24 0.155672
R2573 VDD2.n33 VDD2.n32 0.155672
R2574 VDD2.n10 VDD2.n9 0.155672
R2575 VDD2.n10 VDD2.n1 0.155672
R2576 VDD2.n17 VDD2.n1 0.155672
C0 VDD1 VDD2 3.02125f
C1 VP VN 8.84749f
C2 VN VTAIL 6.12713f
C3 VP VTAIL 6.1415f
C4 VN VDD1 0.16069f
C5 VP VDD1 4.79283f
C6 VN VDD2 4.20345f
C7 VP VDD2 0.753993f
C8 VTAIL VDD1 8.03283f
C9 VTAIL VDD2 8.09471f
C10 VDD2 B 7.44563f
C11 VDD1 B 7.331359f
C12 VTAIL B 5.293057f
C13 VN B 23.61945f
C14 VP B 22.071432f
C15 VDD2.n0 B 0.041139f
C16 VDD2.n1 B 0.028316f
C17 VDD2.n2 B 0.015216f
C18 VDD2.n3 B 0.035965f
C19 VDD2.n4 B 0.016111f
C20 VDD2.n5 B 0.109957f
C21 VDD2.t0 B 0.059969f
C22 VDD2.n6 B 0.026974f
C23 VDD2.n7 B 0.021168f
C24 VDD2.n8 B 0.015216f
C25 VDD2.n9 B 0.413872f
C26 VDD2.n10 B 0.028316f
C27 VDD2.n11 B 0.015216f
C28 VDD2.n12 B 0.016111f
C29 VDD2.n13 B 0.035965f
C30 VDD2.n14 B 0.080224f
C31 VDD2.n15 B 0.016111f
C32 VDD2.n16 B 0.015216f
C33 VDD2.n17 B 0.072802f
C34 VDD2.n18 B 0.090249f
C35 VDD2.t5 B 0.090177f
C36 VDD2.t1 B 0.090177f
C37 VDD2.n19 B 0.708681f
C38 VDD2.n20 B 0.999091f
C39 VDD2.t7 B 0.090177f
C40 VDD2.t2 B 0.090177f
C41 VDD2.n21 B 0.735879f
C42 VDD2.n22 B 3.49686f
C43 VDD2.n23 B 0.041139f
C44 VDD2.n24 B 0.028316f
C45 VDD2.n25 B 0.015216f
C46 VDD2.n26 B 0.035965f
C47 VDD2.n27 B 0.016111f
C48 VDD2.n28 B 0.109957f
C49 VDD2.t8 B 0.059969f
C50 VDD2.n29 B 0.026974f
C51 VDD2.n30 B 0.021168f
C52 VDD2.n31 B 0.015216f
C53 VDD2.n32 B 0.413872f
C54 VDD2.n33 B 0.028316f
C55 VDD2.n34 B 0.015216f
C56 VDD2.n35 B 0.016111f
C57 VDD2.n36 B 0.035965f
C58 VDD2.n37 B 0.080224f
C59 VDD2.n38 B 0.016111f
C60 VDD2.n39 B 0.015216f
C61 VDD2.n40 B 0.072802f
C62 VDD2.n41 B 0.064847f
C63 VDD2.n42 B 3.15275f
C64 VDD2.t4 B 0.090177f
C65 VDD2.t9 B 0.090177f
C66 VDD2.n43 B 0.708684f
C67 VDD2.n44 B 0.642628f
C68 VDD2.t6 B 0.090177f
C69 VDD2.t3 B 0.090177f
C70 VDD2.n45 B 0.735834f
C71 VN.n0 B 0.03979f
C72 VN.t7 B 0.854667f
C73 VN.n1 B 0.040138f
C74 VN.n2 B 0.021153f
C75 VN.n3 B 0.039425f
C76 VN.n4 B 0.021153f
C77 VN.t2 B 0.854667f
C78 VN.n5 B 0.039425f
C79 VN.n6 B 0.021153f
C80 VN.n7 B 0.039425f
C81 VN.n8 B 0.021153f
C82 VN.t8 B 0.854667f
C83 VN.n9 B 0.039425f
C84 VN.n10 B 0.021153f
C85 VN.n11 B 0.039425f
C86 VN.n12 B 0.278112f
C87 VN.t4 B 0.854667f
C88 VN.t9 B 1.13517f
C89 VN.n13 B 0.414721f
C90 VN.n14 B 0.405971f
C91 VN.n15 B 0.028914f
C92 VN.n16 B 0.039425f
C93 VN.n17 B 0.021153f
C94 VN.n18 B 0.021153f
C95 VN.n19 B 0.021153f
C96 VN.n20 B 0.038195f
C97 VN.n21 B 0.02099f
C98 VN.n22 B 0.042004f
C99 VN.n23 B 0.021153f
C100 VN.n24 B 0.021153f
C101 VN.n25 B 0.021153f
C102 VN.n26 B 0.039425f
C103 VN.n27 B 0.350002f
C104 VN.n28 B 0.039425f
C105 VN.n29 B 0.021153f
C106 VN.n30 B 0.021153f
C107 VN.n31 B 0.021153f
C108 VN.n32 B 0.042004f
C109 VN.n33 B 0.02099f
C110 VN.n34 B 0.038195f
C111 VN.n35 B 0.021153f
C112 VN.n36 B 0.021153f
C113 VN.n37 B 0.021153f
C114 VN.n38 B 0.039425f
C115 VN.n39 B 0.028914f
C116 VN.n40 B 0.330042f
C117 VN.n41 B 0.030471f
C118 VN.n42 B 0.021153f
C119 VN.n43 B 0.021153f
C120 VN.n44 B 0.021153f
C121 VN.n45 B 0.039425f
C122 VN.n46 B 0.036375f
C123 VN.n47 B 0.024676f
C124 VN.n48 B 0.021153f
C125 VN.n49 B 0.021153f
C126 VN.n50 B 0.021153f
C127 VN.n51 B 0.039425f
C128 VN.n52 B 0.037868f
C129 VN.n53 B 0.424989f
C130 VN.n54 B 0.064016f
C131 VN.n55 B 0.03979f
C132 VN.t1 B 0.854667f
C133 VN.n56 B 0.040138f
C134 VN.n57 B 0.021153f
C135 VN.n58 B 0.039425f
C136 VN.n59 B 0.021153f
C137 VN.t5 B 0.854667f
C138 VN.n60 B 0.039425f
C139 VN.n61 B 0.021153f
C140 VN.n62 B 0.039425f
C141 VN.n63 B 0.021153f
C142 VN.t0 B 0.854667f
C143 VN.n64 B 0.039425f
C144 VN.n65 B 0.021153f
C145 VN.n66 B 0.039425f
C146 VN.n67 B 0.278112f
C147 VN.t3 B 0.854667f
C148 VN.t6 B 1.13517f
C149 VN.n68 B 0.414721f
C150 VN.n69 B 0.405971f
C151 VN.n70 B 0.028914f
C152 VN.n71 B 0.039425f
C153 VN.n72 B 0.021153f
C154 VN.n73 B 0.021153f
C155 VN.n74 B 0.021153f
C156 VN.n75 B 0.038195f
C157 VN.n76 B 0.02099f
C158 VN.n77 B 0.042004f
C159 VN.n78 B 0.021153f
C160 VN.n79 B 0.021153f
C161 VN.n80 B 0.021153f
C162 VN.n81 B 0.039425f
C163 VN.n82 B 0.350002f
C164 VN.n83 B 0.039425f
C165 VN.n84 B 0.021153f
C166 VN.n85 B 0.021153f
C167 VN.n86 B 0.021153f
C168 VN.n87 B 0.042004f
C169 VN.n88 B 0.02099f
C170 VN.n89 B 0.038195f
C171 VN.n90 B 0.021153f
C172 VN.n91 B 0.021153f
C173 VN.n92 B 0.021153f
C174 VN.n93 B 0.039425f
C175 VN.n94 B 0.028914f
C176 VN.n95 B 0.330042f
C177 VN.n96 B 0.030471f
C178 VN.n97 B 0.021153f
C179 VN.n98 B 0.021153f
C180 VN.n99 B 0.021153f
C181 VN.n100 B 0.039425f
C182 VN.n101 B 0.036375f
C183 VN.n102 B 0.024676f
C184 VN.n103 B 0.021153f
C185 VN.n104 B 0.021153f
C186 VN.n105 B 0.021153f
C187 VN.n106 B 0.039425f
C188 VN.n107 B 0.037868f
C189 VN.n108 B 0.424989f
C190 VN.n109 B 1.38594f
C191 VTAIL.t5 B 0.10594f
C192 VTAIL.t19 B 0.10594f
C193 VTAIL.n0 B 0.762555f
C194 VTAIL.n1 B 0.83011f
C195 VTAIL.n2 B 0.04833f
C196 VTAIL.n3 B 0.033266f
C197 VTAIL.n4 B 0.017876f
C198 VTAIL.n5 B 0.042252f
C199 VTAIL.n6 B 0.018927f
C200 VTAIL.n7 B 0.129178f
C201 VTAIL.t10 B 0.070452f
C202 VTAIL.n8 B 0.031689f
C203 VTAIL.n9 B 0.024868f
C204 VTAIL.n10 B 0.017876f
C205 VTAIL.n11 B 0.486216f
C206 VTAIL.n12 B 0.033266f
C207 VTAIL.n13 B 0.017876f
C208 VTAIL.n14 B 0.018927f
C209 VTAIL.n15 B 0.042252f
C210 VTAIL.n16 B 0.094246f
C211 VTAIL.n17 B 0.018927f
C212 VTAIL.n18 B 0.017876f
C213 VTAIL.n19 B 0.085528f
C214 VTAIL.n20 B 0.053273f
C215 VTAIL.n21 B 0.669975f
C216 VTAIL.t13 B 0.10594f
C217 VTAIL.t16 B 0.10594f
C218 VTAIL.n22 B 0.762555f
C219 VTAIL.n23 B 1.06667f
C220 VTAIL.t14 B 0.10594f
C221 VTAIL.t9 B 0.10594f
C222 VTAIL.n24 B 0.762555f
C223 VTAIL.n25 B 2.28182f
C224 VTAIL.t0 B 0.10594f
C225 VTAIL.t2 B 0.10594f
C226 VTAIL.n26 B 0.76256f
C227 VTAIL.n27 B 2.28182f
C228 VTAIL.t3 B 0.10594f
C229 VTAIL.t7 B 0.10594f
C230 VTAIL.n28 B 0.76256f
C231 VTAIL.n29 B 1.06666f
C232 VTAIL.n30 B 0.04833f
C233 VTAIL.n31 B 0.033266f
C234 VTAIL.n32 B 0.017876f
C235 VTAIL.n33 B 0.042252f
C236 VTAIL.n34 B 0.018927f
C237 VTAIL.n35 B 0.129178f
C238 VTAIL.t4 B 0.070452f
C239 VTAIL.n36 B 0.031689f
C240 VTAIL.n37 B 0.024868f
C241 VTAIL.n38 B 0.017876f
C242 VTAIL.n39 B 0.486216f
C243 VTAIL.n40 B 0.033266f
C244 VTAIL.n41 B 0.017876f
C245 VTAIL.n42 B 0.018927f
C246 VTAIL.n43 B 0.042252f
C247 VTAIL.n44 B 0.094246f
C248 VTAIL.n45 B 0.018927f
C249 VTAIL.n46 B 0.017876f
C250 VTAIL.n47 B 0.085528f
C251 VTAIL.n48 B 0.053273f
C252 VTAIL.n49 B 0.669975f
C253 VTAIL.t15 B 0.10594f
C254 VTAIL.t18 B 0.10594f
C255 VTAIL.n50 B 0.76256f
C256 VTAIL.n51 B 0.921587f
C257 VTAIL.t12 B 0.10594f
C258 VTAIL.t17 B 0.10594f
C259 VTAIL.n52 B 0.76256f
C260 VTAIL.n53 B 1.06666f
C261 VTAIL.n54 B 0.04833f
C262 VTAIL.n55 B 0.033266f
C263 VTAIL.n56 B 0.017876f
C264 VTAIL.n57 B 0.042252f
C265 VTAIL.n58 B 0.018927f
C266 VTAIL.n59 B 0.129178f
C267 VTAIL.t11 B 0.070452f
C268 VTAIL.n60 B 0.031689f
C269 VTAIL.n61 B 0.024868f
C270 VTAIL.n62 B 0.017876f
C271 VTAIL.n63 B 0.486216f
C272 VTAIL.n64 B 0.033266f
C273 VTAIL.n65 B 0.017876f
C274 VTAIL.n66 B 0.018927f
C275 VTAIL.n67 B 0.042252f
C276 VTAIL.n68 B 0.094246f
C277 VTAIL.n69 B 0.018927f
C278 VTAIL.n70 B 0.017876f
C279 VTAIL.n71 B 0.085528f
C280 VTAIL.n72 B 0.053273f
C281 VTAIL.n73 B 1.63933f
C282 VTAIL.n74 B 0.04833f
C283 VTAIL.n75 B 0.033266f
C284 VTAIL.n76 B 0.017876f
C285 VTAIL.n77 B 0.042252f
C286 VTAIL.n78 B 0.018927f
C287 VTAIL.n79 B 0.129178f
C288 VTAIL.t1 B 0.070452f
C289 VTAIL.n80 B 0.031689f
C290 VTAIL.n81 B 0.024868f
C291 VTAIL.n82 B 0.017876f
C292 VTAIL.n83 B 0.486216f
C293 VTAIL.n84 B 0.033266f
C294 VTAIL.n85 B 0.017876f
C295 VTAIL.n86 B 0.018927f
C296 VTAIL.n87 B 0.042252f
C297 VTAIL.n88 B 0.094246f
C298 VTAIL.n89 B 0.018927f
C299 VTAIL.n90 B 0.017876f
C300 VTAIL.n91 B 0.085528f
C301 VTAIL.n92 B 0.053273f
C302 VTAIL.n93 B 1.63933f
C303 VTAIL.t6 B 0.10594f
C304 VTAIL.t8 B 0.10594f
C305 VTAIL.n94 B 0.762555f
C306 VTAIL.n95 B 0.767274f
C307 VDD1.n0 B 0.042195f
C308 VDD1.n1 B 0.029043f
C309 VDD1.n2 B 0.015607f
C310 VDD1.n3 B 0.036888f
C311 VDD1.n4 B 0.016525f
C312 VDD1.n5 B 0.11278f
C313 VDD1.t6 B 0.061509f
C314 VDD1.n6 B 0.027666f
C315 VDD1.n7 B 0.021711f
C316 VDD1.n8 B 0.015607f
C317 VDD1.n9 B 0.424496f
C318 VDD1.n10 B 0.029043f
C319 VDD1.n11 B 0.015607f
C320 VDD1.n12 B 0.016525f
C321 VDD1.n13 B 0.036888f
C322 VDD1.n14 B 0.082283f
C323 VDD1.n15 B 0.016525f
C324 VDD1.n16 B 0.015607f
C325 VDD1.n17 B 0.074671f
C326 VDD1.n18 B 0.092566f
C327 VDD1.t0 B 0.092492f
C328 VDD1.t7 B 0.092492f
C329 VDD1.n19 B 0.726875f
C330 VDD1.n20 B 1.03457f
C331 VDD1.n21 B 0.042195f
C332 VDD1.n22 B 0.029043f
C333 VDD1.n23 B 0.015607f
C334 VDD1.n24 B 0.036888f
C335 VDD1.n25 B 0.016525f
C336 VDD1.n26 B 0.11278f
C337 VDD1.t5 B 0.061509f
C338 VDD1.n27 B 0.027666f
C339 VDD1.n28 B 0.021711f
C340 VDD1.n29 B 0.015607f
C341 VDD1.n30 B 0.424496f
C342 VDD1.n31 B 0.029043f
C343 VDD1.n32 B 0.015607f
C344 VDD1.n33 B 0.016525f
C345 VDD1.n34 B 0.036888f
C346 VDD1.n35 B 0.082283f
C347 VDD1.n36 B 0.016525f
C348 VDD1.n37 B 0.015607f
C349 VDD1.n38 B 0.074671f
C350 VDD1.n39 B 0.092566f
C351 VDD1.t3 B 0.092492f
C352 VDD1.t1 B 0.092492f
C353 VDD1.n40 B 0.726871f
C354 VDD1.n41 B 1.02474f
C355 VDD1.t9 B 0.092492f
C356 VDD1.t4 B 0.092492f
C357 VDD1.n42 B 0.754768f
C358 VDD1.n43 B 3.76456f
C359 VDD1.t8 B 0.092492f
C360 VDD1.t2 B 0.092492f
C361 VDD1.n44 B 0.726871f
C362 VDD1.n45 B 3.59207f
C363 VP.n0 B 0.041104f
C364 VP.t8 B 0.882889f
C365 VP.n1 B 0.041464f
C366 VP.n2 B 0.021852f
C367 VP.n3 B 0.040727f
C368 VP.n4 B 0.021852f
C369 VP.t2 B 0.882889f
C370 VP.n5 B 0.040727f
C371 VP.n6 B 0.021852f
C372 VP.n7 B 0.040727f
C373 VP.n8 B 0.021852f
C374 VP.t5 B 0.882889f
C375 VP.n9 B 0.040727f
C376 VP.n10 B 0.021852f
C377 VP.n11 B 0.040727f
C378 VP.n12 B 0.021852f
C379 VP.t9 B 0.882889f
C380 VP.n13 B 0.040727f
C381 VP.n14 B 0.021852f
C382 VP.n15 B 0.041464f
C383 VP.n16 B 0.041104f
C384 VP.t4 B 0.882889f
C385 VP.n17 B 0.041104f
C386 VP.t7 B 0.882889f
C387 VP.n18 B 0.041464f
C388 VP.n19 B 0.021852f
C389 VP.n20 B 0.040727f
C390 VP.n21 B 0.021852f
C391 VP.t1 B 0.882889f
C392 VP.n22 B 0.040727f
C393 VP.n23 B 0.021852f
C394 VP.n24 B 0.040727f
C395 VP.n25 B 0.021852f
C396 VP.t6 B 0.882889f
C397 VP.n26 B 0.040727f
C398 VP.n27 B 0.021852f
C399 VP.n28 B 0.040727f
C400 VP.n29 B 0.287296f
C401 VP.t0 B 0.882889f
C402 VP.t3 B 1.17265f
C403 VP.n30 B 0.428418f
C404 VP.n31 B 0.419377f
C405 VP.n32 B 0.029869f
C406 VP.n33 B 0.040727f
C407 VP.n34 B 0.021852f
C408 VP.n35 B 0.021852f
C409 VP.n36 B 0.021852f
C410 VP.n37 B 0.039457f
C411 VP.n38 B 0.021684f
C412 VP.n39 B 0.043391f
C413 VP.n40 B 0.021852f
C414 VP.n41 B 0.021852f
C415 VP.n42 B 0.021852f
C416 VP.n43 B 0.040727f
C417 VP.n44 B 0.36156f
C418 VP.n45 B 0.040727f
C419 VP.n46 B 0.021852f
C420 VP.n47 B 0.021852f
C421 VP.n48 B 0.021852f
C422 VP.n49 B 0.043391f
C423 VP.n50 B 0.021684f
C424 VP.n51 B 0.039457f
C425 VP.n52 B 0.021852f
C426 VP.n53 B 0.021852f
C427 VP.n54 B 0.021852f
C428 VP.n55 B 0.040727f
C429 VP.n56 B 0.029869f
C430 VP.n57 B 0.340941f
C431 VP.n58 B 0.031477f
C432 VP.n59 B 0.021852f
C433 VP.n60 B 0.021852f
C434 VP.n61 B 0.021852f
C435 VP.n62 B 0.040727f
C436 VP.n63 B 0.037577f
C437 VP.n64 B 0.02549f
C438 VP.n65 B 0.021852f
C439 VP.n66 B 0.021852f
C440 VP.n67 B 0.021852f
C441 VP.n68 B 0.040727f
C442 VP.n69 B 0.039118f
C443 VP.n70 B 0.439022f
C444 VP.n71 B 1.42634f
C445 VP.n72 B 1.44078f
C446 VP.n73 B 0.439022f
C447 VP.n74 B 0.039118f
C448 VP.n75 B 0.040727f
C449 VP.n76 B 0.021852f
C450 VP.n77 B 0.021852f
C451 VP.n78 B 0.021852f
C452 VP.n79 B 0.02549f
C453 VP.n80 B 0.037577f
C454 VP.n81 B 0.040727f
C455 VP.n82 B 0.021852f
C456 VP.n83 B 0.021852f
C457 VP.n84 B 0.021852f
C458 VP.n85 B 0.031477f
C459 VP.n86 B 0.340941f
C460 VP.n87 B 0.029869f
C461 VP.n88 B 0.040727f
C462 VP.n89 B 0.021852f
C463 VP.n90 B 0.021852f
C464 VP.n91 B 0.021852f
C465 VP.n92 B 0.039457f
C466 VP.n93 B 0.021684f
C467 VP.n94 B 0.043391f
C468 VP.n95 B 0.021852f
C469 VP.n96 B 0.021852f
C470 VP.n97 B 0.021852f
C471 VP.n98 B 0.040727f
C472 VP.n99 B 0.36156f
C473 VP.n100 B 0.040727f
C474 VP.n101 B 0.021852f
C475 VP.n102 B 0.021852f
C476 VP.n103 B 0.021852f
C477 VP.n104 B 0.043391f
C478 VP.n105 B 0.021684f
C479 VP.n106 B 0.039457f
C480 VP.n107 B 0.021852f
C481 VP.n108 B 0.021852f
C482 VP.n109 B 0.021852f
C483 VP.n110 B 0.040727f
C484 VP.n111 B 0.029869f
C485 VP.n112 B 0.340941f
C486 VP.n113 B 0.031477f
C487 VP.n114 B 0.021852f
C488 VP.n115 B 0.021852f
C489 VP.n116 B 0.021852f
C490 VP.n117 B 0.040727f
C491 VP.n118 B 0.037577f
C492 VP.n119 B 0.02549f
C493 VP.n120 B 0.021852f
C494 VP.n121 B 0.021852f
C495 VP.n122 B 0.021852f
C496 VP.n123 B 0.040727f
C497 VP.n124 B 0.039118f
C498 VP.n125 B 0.439022f
C499 VP.n126 B 0.066131f
.ends

