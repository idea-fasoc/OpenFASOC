* NGSPICE file created from diff_pair_sample_0240.ext - technology: sky130A

.subckt diff_pair_sample_0240 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=6.7509 pd=35.4 as=2.85615 ps=17.64 w=17.31 l=0.89
X1 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=6.7509 pd=35.4 as=0 ps=0 w=17.31 l=0.89
X2 VTAIL.t1 VP.t0 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.85615 pd=17.64 as=2.85615 ps=17.64 w=17.31 l=0.89
X3 VDD1.t4 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.7509 pd=35.4 as=2.85615 ps=17.64 w=17.31 l=0.89
X4 VTAIL.t3 VP.t2 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.85615 pd=17.64 as=2.85615 ps=17.64 w=17.31 l=0.89
X5 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=6.7509 pd=35.4 as=0 ps=0 w=17.31 l=0.89
X6 VDD2.t4 VN.t1 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=2.85615 pd=17.64 as=6.7509 ps=35.4 w=17.31 l=0.89
X7 VTAIL.t8 VN.t2 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.85615 pd=17.64 as=2.85615 ps=17.64 w=17.31 l=0.89
X8 VDD1.t2 VP.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.85615 pd=17.64 as=6.7509 ps=35.4 w=17.31 l=0.89
X9 VDD1.t1 VP.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.85615 pd=17.64 as=6.7509 ps=35.4 w=17.31 l=0.89
X10 VDD2.t2 VN.t3 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=2.85615 pd=17.64 as=6.7509 ps=35.4 w=17.31 l=0.89
X11 VTAIL.t11 VN.t4 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.85615 pd=17.64 as=2.85615 ps=17.64 w=17.31 l=0.89
X12 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.7509 pd=35.4 as=0 ps=0 w=17.31 l=0.89
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.7509 pd=35.4 as=0 ps=0 w=17.31 l=0.89
X14 VDD1.t0 VP.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.7509 pd=35.4 as=2.85615 ps=17.64 w=17.31 l=0.89
X15 VDD2.t0 VN.t5 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=6.7509 pd=35.4 as=2.85615 ps=17.64 w=17.31 l=0.89
R0 VN.n2 VN.t5 529.992
R1 VN.n10 VN.t3 529.992
R2 VN.n6 VN.t1 513.14
R3 VN.n14 VN.t0 513.14
R4 VN.n1 VN.t2 468.731
R5 VN.n9 VN.t4 468.731
R6 VN.n7 VN.n6 161.3
R7 VN.n15 VN.n14 161.3
R8 VN.n13 VN.n8 161.3
R9 VN.n12 VN.n11 161.3
R10 VN.n5 VN.n0 161.3
R11 VN.n4 VN.n3 161.3
R12 VN.n5 VN.n4 54.0911
R13 VN.n13 VN.n12 54.0911
R14 VN VN.n15 46.3509
R15 VN.n11 VN.n10 43.6035
R16 VN.n3 VN.n2 43.6035
R17 VN.n2 VN.n1 42.5728
R18 VN.n10 VN.n9 42.5728
R19 VN.n4 VN.n1 12.234
R20 VN.n12 VN.n9 12.234
R21 VN.n6 VN.n5 3.65202
R22 VN.n14 VN.n13 3.65202
R23 VN.n15 VN.n8 0.189894
R24 VN.n11 VN.n8 0.189894
R25 VN.n3 VN.n0 0.189894
R26 VN.n7 VN.n0 0.189894
R27 VN VN.n7 0.0516364
R28 VTAIL.n7 VTAIL.t9 48.0762
R29 VTAIL.n11 VTAIL.t10 48.076
R30 VTAIL.n2 VTAIL.t4 48.076
R31 VTAIL.n10 VTAIL.t5 48.076
R32 VTAIL.n9 VTAIL.n8 46.9324
R33 VTAIL.n6 VTAIL.n5 46.9324
R34 VTAIL.n1 VTAIL.n0 46.9321
R35 VTAIL.n4 VTAIL.n3 46.9321
R36 VTAIL.n6 VTAIL.n4 29.3927
R37 VTAIL.n11 VTAIL.n10 28.341
R38 VTAIL.n0 VTAIL.t7 1.14435
R39 VTAIL.n0 VTAIL.t8 1.14435
R40 VTAIL.n3 VTAIL.t2 1.14435
R41 VTAIL.n3 VTAIL.t1 1.14435
R42 VTAIL.n8 VTAIL.t0 1.14435
R43 VTAIL.n8 VTAIL.t3 1.14435
R44 VTAIL.n5 VTAIL.t6 1.14435
R45 VTAIL.n5 VTAIL.t11 1.14435
R46 VTAIL.n7 VTAIL.n6 1.05222
R47 VTAIL.n10 VTAIL.n9 1.05222
R48 VTAIL.n4 VTAIL.n2 1.05222
R49 VTAIL.n9 VTAIL.n7 0.99619
R50 VTAIL.n2 VTAIL.n1 0.99619
R51 VTAIL VTAIL.n11 0.731103
R52 VTAIL VTAIL.n1 0.321621
R53 VDD2.n1 VDD2.t0 65.4883
R54 VDD2.n2 VDD2.t5 64.7549
R55 VDD2.n1 VDD2.n0 63.8185
R56 VDD2 VDD2.n3 63.8157
R57 VDD2.n2 VDD2.n1 42.0558
R58 VDD2.n3 VDD2.t1 1.14435
R59 VDD2.n3 VDD2.t2 1.14435
R60 VDD2.n0 VDD2.t3 1.14435
R61 VDD2.n0 VDD2.t4 1.14435
R62 VDD2 VDD2.n2 0.847483
R63 B.n74 B.t17 670.85
R64 B.n82 B.t6 670.85
R65 B.n189 B.t14 670.85
R66 B.n181 B.t10 670.85
R67 B.n566 B.n565 585
R68 B.n568 B.n111 585
R69 B.n571 B.n570 585
R70 B.n572 B.n110 585
R71 B.n574 B.n573 585
R72 B.n576 B.n109 585
R73 B.n579 B.n578 585
R74 B.n580 B.n108 585
R75 B.n582 B.n581 585
R76 B.n584 B.n107 585
R77 B.n587 B.n586 585
R78 B.n588 B.n106 585
R79 B.n590 B.n589 585
R80 B.n592 B.n105 585
R81 B.n595 B.n594 585
R82 B.n596 B.n104 585
R83 B.n598 B.n597 585
R84 B.n600 B.n103 585
R85 B.n603 B.n602 585
R86 B.n604 B.n102 585
R87 B.n606 B.n605 585
R88 B.n608 B.n101 585
R89 B.n611 B.n610 585
R90 B.n612 B.n100 585
R91 B.n614 B.n613 585
R92 B.n616 B.n99 585
R93 B.n619 B.n618 585
R94 B.n620 B.n98 585
R95 B.n622 B.n621 585
R96 B.n624 B.n97 585
R97 B.n627 B.n626 585
R98 B.n628 B.n96 585
R99 B.n630 B.n629 585
R100 B.n632 B.n95 585
R101 B.n635 B.n634 585
R102 B.n636 B.n94 585
R103 B.n638 B.n637 585
R104 B.n640 B.n93 585
R105 B.n643 B.n642 585
R106 B.n644 B.n92 585
R107 B.n646 B.n645 585
R108 B.n648 B.n91 585
R109 B.n651 B.n650 585
R110 B.n652 B.n90 585
R111 B.n654 B.n653 585
R112 B.n656 B.n89 585
R113 B.n659 B.n658 585
R114 B.n660 B.n88 585
R115 B.n662 B.n661 585
R116 B.n664 B.n87 585
R117 B.n667 B.n666 585
R118 B.n668 B.n86 585
R119 B.n670 B.n669 585
R120 B.n672 B.n85 585
R121 B.n675 B.n674 585
R122 B.n676 B.n81 585
R123 B.n678 B.n677 585
R124 B.n680 B.n80 585
R125 B.n683 B.n682 585
R126 B.n684 B.n79 585
R127 B.n686 B.n685 585
R128 B.n688 B.n78 585
R129 B.n691 B.n690 585
R130 B.n692 B.n77 585
R131 B.n694 B.n693 585
R132 B.n696 B.n76 585
R133 B.n699 B.n698 585
R134 B.n701 B.n73 585
R135 B.n703 B.n702 585
R136 B.n705 B.n72 585
R137 B.n708 B.n707 585
R138 B.n709 B.n71 585
R139 B.n711 B.n710 585
R140 B.n713 B.n70 585
R141 B.n716 B.n715 585
R142 B.n717 B.n69 585
R143 B.n719 B.n718 585
R144 B.n721 B.n68 585
R145 B.n724 B.n723 585
R146 B.n725 B.n67 585
R147 B.n727 B.n726 585
R148 B.n729 B.n66 585
R149 B.n732 B.n731 585
R150 B.n733 B.n65 585
R151 B.n735 B.n734 585
R152 B.n737 B.n64 585
R153 B.n740 B.n739 585
R154 B.n741 B.n63 585
R155 B.n743 B.n742 585
R156 B.n745 B.n62 585
R157 B.n748 B.n747 585
R158 B.n749 B.n61 585
R159 B.n751 B.n750 585
R160 B.n753 B.n60 585
R161 B.n756 B.n755 585
R162 B.n757 B.n59 585
R163 B.n759 B.n758 585
R164 B.n761 B.n58 585
R165 B.n764 B.n763 585
R166 B.n765 B.n57 585
R167 B.n767 B.n766 585
R168 B.n769 B.n56 585
R169 B.n772 B.n771 585
R170 B.n773 B.n55 585
R171 B.n775 B.n774 585
R172 B.n777 B.n54 585
R173 B.n780 B.n779 585
R174 B.n781 B.n53 585
R175 B.n783 B.n782 585
R176 B.n785 B.n52 585
R177 B.n788 B.n787 585
R178 B.n789 B.n51 585
R179 B.n791 B.n790 585
R180 B.n793 B.n50 585
R181 B.n796 B.n795 585
R182 B.n797 B.n49 585
R183 B.n799 B.n798 585
R184 B.n801 B.n48 585
R185 B.n804 B.n803 585
R186 B.n805 B.n47 585
R187 B.n807 B.n806 585
R188 B.n809 B.n46 585
R189 B.n812 B.n811 585
R190 B.n813 B.n45 585
R191 B.n564 B.n43 585
R192 B.n816 B.n43 585
R193 B.n563 B.n42 585
R194 B.n817 B.n42 585
R195 B.n562 B.n41 585
R196 B.n818 B.n41 585
R197 B.n561 B.n560 585
R198 B.n560 B.n37 585
R199 B.n559 B.n36 585
R200 B.n824 B.n36 585
R201 B.n558 B.n35 585
R202 B.n825 B.n35 585
R203 B.n557 B.n34 585
R204 B.n826 B.n34 585
R205 B.n556 B.n555 585
R206 B.n555 B.n30 585
R207 B.n554 B.n29 585
R208 B.n832 B.n29 585
R209 B.n553 B.n28 585
R210 B.n833 B.n28 585
R211 B.n552 B.n27 585
R212 B.n834 B.n27 585
R213 B.n551 B.n550 585
R214 B.n550 B.n26 585
R215 B.n549 B.n22 585
R216 B.n840 B.n22 585
R217 B.n548 B.n21 585
R218 B.n841 B.n21 585
R219 B.n547 B.n20 585
R220 B.n842 B.n20 585
R221 B.n546 B.n545 585
R222 B.n545 B.n19 585
R223 B.n544 B.n15 585
R224 B.n848 B.n15 585
R225 B.n543 B.n14 585
R226 B.n849 B.n14 585
R227 B.n542 B.n13 585
R228 B.n850 B.n13 585
R229 B.n541 B.n540 585
R230 B.n540 B.n12 585
R231 B.n539 B.n538 585
R232 B.n539 B.n8 585
R233 B.n537 B.n7 585
R234 B.n857 B.n7 585
R235 B.n536 B.n6 585
R236 B.n858 B.n6 585
R237 B.n535 B.n5 585
R238 B.n859 B.n5 585
R239 B.n534 B.n533 585
R240 B.n533 B.n4 585
R241 B.n532 B.n112 585
R242 B.n532 B.n531 585
R243 B.n521 B.n113 585
R244 B.n524 B.n113 585
R245 B.n523 B.n522 585
R246 B.n525 B.n523 585
R247 B.n520 B.n118 585
R248 B.n118 B.n117 585
R249 B.n519 B.n518 585
R250 B.n518 B.n517 585
R251 B.n120 B.n119 585
R252 B.n510 B.n120 585
R253 B.n509 B.n508 585
R254 B.n511 B.n509 585
R255 B.n507 B.n125 585
R256 B.n125 B.n124 585
R257 B.n506 B.n505 585
R258 B.n505 B.n504 585
R259 B.n127 B.n126 585
R260 B.n497 B.n127 585
R261 B.n496 B.n495 585
R262 B.n498 B.n496 585
R263 B.n494 B.n132 585
R264 B.n132 B.n131 585
R265 B.n493 B.n492 585
R266 B.n492 B.n491 585
R267 B.n134 B.n133 585
R268 B.n135 B.n134 585
R269 B.n484 B.n483 585
R270 B.n485 B.n484 585
R271 B.n482 B.n139 585
R272 B.n143 B.n139 585
R273 B.n481 B.n480 585
R274 B.n480 B.n479 585
R275 B.n141 B.n140 585
R276 B.n142 B.n141 585
R277 B.n472 B.n471 585
R278 B.n473 B.n472 585
R279 B.n470 B.n148 585
R280 B.n148 B.n147 585
R281 B.n469 B.n468 585
R282 B.n468 B.n467 585
R283 B.n464 B.n152 585
R284 B.n463 B.n462 585
R285 B.n460 B.n153 585
R286 B.n460 B.n151 585
R287 B.n459 B.n458 585
R288 B.n457 B.n456 585
R289 B.n455 B.n155 585
R290 B.n453 B.n452 585
R291 B.n451 B.n156 585
R292 B.n450 B.n449 585
R293 B.n447 B.n157 585
R294 B.n445 B.n444 585
R295 B.n443 B.n158 585
R296 B.n442 B.n441 585
R297 B.n439 B.n159 585
R298 B.n437 B.n436 585
R299 B.n435 B.n160 585
R300 B.n434 B.n433 585
R301 B.n431 B.n161 585
R302 B.n429 B.n428 585
R303 B.n427 B.n162 585
R304 B.n426 B.n425 585
R305 B.n423 B.n163 585
R306 B.n421 B.n420 585
R307 B.n419 B.n164 585
R308 B.n418 B.n417 585
R309 B.n415 B.n165 585
R310 B.n413 B.n412 585
R311 B.n411 B.n166 585
R312 B.n410 B.n409 585
R313 B.n407 B.n167 585
R314 B.n405 B.n404 585
R315 B.n403 B.n168 585
R316 B.n402 B.n401 585
R317 B.n399 B.n169 585
R318 B.n397 B.n396 585
R319 B.n395 B.n170 585
R320 B.n394 B.n393 585
R321 B.n391 B.n171 585
R322 B.n389 B.n388 585
R323 B.n387 B.n172 585
R324 B.n386 B.n385 585
R325 B.n383 B.n173 585
R326 B.n381 B.n380 585
R327 B.n379 B.n174 585
R328 B.n378 B.n377 585
R329 B.n375 B.n175 585
R330 B.n373 B.n372 585
R331 B.n371 B.n176 585
R332 B.n370 B.n369 585
R333 B.n367 B.n177 585
R334 B.n365 B.n364 585
R335 B.n363 B.n178 585
R336 B.n362 B.n361 585
R337 B.n359 B.n179 585
R338 B.n357 B.n356 585
R339 B.n355 B.n180 585
R340 B.n354 B.n353 585
R341 B.n351 B.n350 585
R342 B.n349 B.n348 585
R343 B.n347 B.n185 585
R344 B.n345 B.n344 585
R345 B.n343 B.n186 585
R346 B.n342 B.n341 585
R347 B.n339 B.n187 585
R348 B.n337 B.n336 585
R349 B.n335 B.n188 585
R350 B.n334 B.n333 585
R351 B.n331 B.n330 585
R352 B.n329 B.n328 585
R353 B.n327 B.n193 585
R354 B.n325 B.n324 585
R355 B.n323 B.n194 585
R356 B.n322 B.n321 585
R357 B.n319 B.n195 585
R358 B.n317 B.n316 585
R359 B.n315 B.n196 585
R360 B.n314 B.n313 585
R361 B.n311 B.n197 585
R362 B.n309 B.n308 585
R363 B.n307 B.n198 585
R364 B.n306 B.n305 585
R365 B.n303 B.n199 585
R366 B.n301 B.n300 585
R367 B.n299 B.n200 585
R368 B.n298 B.n297 585
R369 B.n295 B.n201 585
R370 B.n293 B.n292 585
R371 B.n291 B.n202 585
R372 B.n290 B.n289 585
R373 B.n287 B.n203 585
R374 B.n285 B.n284 585
R375 B.n283 B.n204 585
R376 B.n282 B.n281 585
R377 B.n279 B.n205 585
R378 B.n277 B.n276 585
R379 B.n275 B.n206 585
R380 B.n274 B.n273 585
R381 B.n271 B.n207 585
R382 B.n269 B.n268 585
R383 B.n267 B.n208 585
R384 B.n266 B.n265 585
R385 B.n263 B.n209 585
R386 B.n261 B.n260 585
R387 B.n259 B.n210 585
R388 B.n258 B.n257 585
R389 B.n255 B.n211 585
R390 B.n253 B.n252 585
R391 B.n251 B.n212 585
R392 B.n250 B.n249 585
R393 B.n247 B.n213 585
R394 B.n245 B.n244 585
R395 B.n243 B.n214 585
R396 B.n242 B.n241 585
R397 B.n239 B.n215 585
R398 B.n237 B.n236 585
R399 B.n235 B.n216 585
R400 B.n234 B.n233 585
R401 B.n231 B.n217 585
R402 B.n229 B.n228 585
R403 B.n227 B.n218 585
R404 B.n226 B.n225 585
R405 B.n223 B.n219 585
R406 B.n221 B.n220 585
R407 B.n150 B.n149 585
R408 B.n151 B.n150 585
R409 B.n466 B.n465 585
R410 B.n467 B.n466 585
R411 B.n146 B.n145 585
R412 B.n147 B.n146 585
R413 B.n475 B.n474 585
R414 B.n474 B.n473 585
R415 B.n476 B.n144 585
R416 B.n144 B.n142 585
R417 B.n478 B.n477 585
R418 B.n479 B.n478 585
R419 B.n138 B.n137 585
R420 B.n143 B.n138 585
R421 B.n487 B.n486 585
R422 B.n486 B.n485 585
R423 B.n488 B.n136 585
R424 B.n136 B.n135 585
R425 B.n490 B.n489 585
R426 B.n491 B.n490 585
R427 B.n130 B.n129 585
R428 B.n131 B.n130 585
R429 B.n500 B.n499 585
R430 B.n499 B.n498 585
R431 B.n501 B.n128 585
R432 B.n497 B.n128 585
R433 B.n503 B.n502 585
R434 B.n504 B.n503 585
R435 B.n123 B.n122 585
R436 B.n124 B.n123 585
R437 B.n513 B.n512 585
R438 B.n512 B.n511 585
R439 B.n514 B.n121 585
R440 B.n510 B.n121 585
R441 B.n516 B.n515 585
R442 B.n517 B.n516 585
R443 B.n116 B.n115 585
R444 B.n117 B.n116 585
R445 B.n527 B.n526 585
R446 B.n526 B.n525 585
R447 B.n528 B.n114 585
R448 B.n524 B.n114 585
R449 B.n530 B.n529 585
R450 B.n531 B.n530 585
R451 B.n3 B.n0 585
R452 B.n4 B.n3 585
R453 B.n856 B.n1 585
R454 B.n857 B.n856 585
R455 B.n855 B.n854 585
R456 B.n855 B.n8 585
R457 B.n853 B.n9 585
R458 B.n12 B.n9 585
R459 B.n852 B.n851 585
R460 B.n851 B.n850 585
R461 B.n11 B.n10 585
R462 B.n849 B.n11 585
R463 B.n847 B.n846 585
R464 B.n848 B.n847 585
R465 B.n845 B.n16 585
R466 B.n19 B.n16 585
R467 B.n844 B.n843 585
R468 B.n843 B.n842 585
R469 B.n18 B.n17 585
R470 B.n841 B.n18 585
R471 B.n839 B.n838 585
R472 B.n840 B.n839 585
R473 B.n837 B.n23 585
R474 B.n26 B.n23 585
R475 B.n836 B.n835 585
R476 B.n835 B.n834 585
R477 B.n25 B.n24 585
R478 B.n833 B.n25 585
R479 B.n831 B.n830 585
R480 B.n832 B.n831 585
R481 B.n829 B.n31 585
R482 B.n31 B.n30 585
R483 B.n828 B.n827 585
R484 B.n827 B.n826 585
R485 B.n33 B.n32 585
R486 B.n825 B.n33 585
R487 B.n823 B.n822 585
R488 B.n824 B.n823 585
R489 B.n821 B.n38 585
R490 B.n38 B.n37 585
R491 B.n820 B.n819 585
R492 B.n819 B.n818 585
R493 B.n40 B.n39 585
R494 B.n817 B.n40 585
R495 B.n815 B.n814 585
R496 B.n816 B.n815 585
R497 B.n860 B.n859 585
R498 B.n858 B.n2 585
R499 B.n815 B.n45 497.305
R500 B.n566 B.n43 497.305
R501 B.n468 B.n150 497.305
R502 B.n466 B.n152 497.305
R503 B.n567 B.n44 256.663
R504 B.n569 B.n44 256.663
R505 B.n575 B.n44 256.663
R506 B.n577 B.n44 256.663
R507 B.n583 B.n44 256.663
R508 B.n585 B.n44 256.663
R509 B.n591 B.n44 256.663
R510 B.n593 B.n44 256.663
R511 B.n599 B.n44 256.663
R512 B.n601 B.n44 256.663
R513 B.n607 B.n44 256.663
R514 B.n609 B.n44 256.663
R515 B.n615 B.n44 256.663
R516 B.n617 B.n44 256.663
R517 B.n623 B.n44 256.663
R518 B.n625 B.n44 256.663
R519 B.n631 B.n44 256.663
R520 B.n633 B.n44 256.663
R521 B.n639 B.n44 256.663
R522 B.n641 B.n44 256.663
R523 B.n647 B.n44 256.663
R524 B.n649 B.n44 256.663
R525 B.n655 B.n44 256.663
R526 B.n657 B.n44 256.663
R527 B.n663 B.n44 256.663
R528 B.n665 B.n44 256.663
R529 B.n671 B.n44 256.663
R530 B.n673 B.n44 256.663
R531 B.n679 B.n44 256.663
R532 B.n681 B.n44 256.663
R533 B.n687 B.n44 256.663
R534 B.n689 B.n44 256.663
R535 B.n695 B.n44 256.663
R536 B.n697 B.n44 256.663
R537 B.n704 B.n44 256.663
R538 B.n706 B.n44 256.663
R539 B.n712 B.n44 256.663
R540 B.n714 B.n44 256.663
R541 B.n720 B.n44 256.663
R542 B.n722 B.n44 256.663
R543 B.n728 B.n44 256.663
R544 B.n730 B.n44 256.663
R545 B.n736 B.n44 256.663
R546 B.n738 B.n44 256.663
R547 B.n744 B.n44 256.663
R548 B.n746 B.n44 256.663
R549 B.n752 B.n44 256.663
R550 B.n754 B.n44 256.663
R551 B.n760 B.n44 256.663
R552 B.n762 B.n44 256.663
R553 B.n768 B.n44 256.663
R554 B.n770 B.n44 256.663
R555 B.n776 B.n44 256.663
R556 B.n778 B.n44 256.663
R557 B.n784 B.n44 256.663
R558 B.n786 B.n44 256.663
R559 B.n792 B.n44 256.663
R560 B.n794 B.n44 256.663
R561 B.n800 B.n44 256.663
R562 B.n802 B.n44 256.663
R563 B.n808 B.n44 256.663
R564 B.n810 B.n44 256.663
R565 B.n461 B.n151 256.663
R566 B.n154 B.n151 256.663
R567 B.n454 B.n151 256.663
R568 B.n448 B.n151 256.663
R569 B.n446 B.n151 256.663
R570 B.n440 B.n151 256.663
R571 B.n438 B.n151 256.663
R572 B.n432 B.n151 256.663
R573 B.n430 B.n151 256.663
R574 B.n424 B.n151 256.663
R575 B.n422 B.n151 256.663
R576 B.n416 B.n151 256.663
R577 B.n414 B.n151 256.663
R578 B.n408 B.n151 256.663
R579 B.n406 B.n151 256.663
R580 B.n400 B.n151 256.663
R581 B.n398 B.n151 256.663
R582 B.n392 B.n151 256.663
R583 B.n390 B.n151 256.663
R584 B.n384 B.n151 256.663
R585 B.n382 B.n151 256.663
R586 B.n376 B.n151 256.663
R587 B.n374 B.n151 256.663
R588 B.n368 B.n151 256.663
R589 B.n366 B.n151 256.663
R590 B.n360 B.n151 256.663
R591 B.n358 B.n151 256.663
R592 B.n352 B.n151 256.663
R593 B.n184 B.n151 256.663
R594 B.n346 B.n151 256.663
R595 B.n340 B.n151 256.663
R596 B.n338 B.n151 256.663
R597 B.n332 B.n151 256.663
R598 B.n192 B.n151 256.663
R599 B.n326 B.n151 256.663
R600 B.n320 B.n151 256.663
R601 B.n318 B.n151 256.663
R602 B.n312 B.n151 256.663
R603 B.n310 B.n151 256.663
R604 B.n304 B.n151 256.663
R605 B.n302 B.n151 256.663
R606 B.n296 B.n151 256.663
R607 B.n294 B.n151 256.663
R608 B.n288 B.n151 256.663
R609 B.n286 B.n151 256.663
R610 B.n280 B.n151 256.663
R611 B.n278 B.n151 256.663
R612 B.n272 B.n151 256.663
R613 B.n270 B.n151 256.663
R614 B.n264 B.n151 256.663
R615 B.n262 B.n151 256.663
R616 B.n256 B.n151 256.663
R617 B.n254 B.n151 256.663
R618 B.n248 B.n151 256.663
R619 B.n246 B.n151 256.663
R620 B.n240 B.n151 256.663
R621 B.n238 B.n151 256.663
R622 B.n232 B.n151 256.663
R623 B.n230 B.n151 256.663
R624 B.n224 B.n151 256.663
R625 B.n222 B.n151 256.663
R626 B.n862 B.n861 256.663
R627 B.n811 B.n809 163.367
R628 B.n807 B.n47 163.367
R629 B.n803 B.n801 163.367
R630 B.n799 B.n49 163.367
R631 B.n795 B.n793 163.367
R632 B.n791 B.n51 163.367
R633 B.n787 B.n785 163.367
R634 B.n783 B.n53 163.367
R635 B.n779 B.n777 163.367
R636 B.n775 B.n55 163.367
R637 B.n771 B.n769 163.367
R638 B.n767 B.n57 163.367
R639 B.n763 B.n761 163.367
R640 B.n759 B.n59 163.367
R641 B.n755 B.n753 163.367
R642 B.n751 B.n61 163.367
R643 B.n747 B.n745 163.367
R644 B.n743 B.n63 163.367
R645 B.n739 B.n737 163.367
R646 B.n735 B.n65 163.367
R647 B.n731 B.n729 163.367
R648 B.n727 B.n67 163.367
R649 B.n723 B.n721 163.367
R650 B.n719 B.n69 163.367
R651 B.n715 B.n713 163.367
R652 B.n711 B.n71 163.367
R653 B.n707 B.n705 163.367
R654 B.n703 B.n73 163.367
R655 B.n698 B.n696 163.367
R656 B.n694 B.n77 163.367
R657 B.n690 B.n688 163.367
R658 B.n686 B.n79 163.367
R659 B.n682 B.n680 163.367
R660 B.n678 B.n81 163.367
R661 B.n674 B.n672 163.367
R662 B.n670 B.n86 163.367
R663 B.n666 B.n664 163.367
R664 B.n662 B.n88 163.367
R665 B.n658 B.n656 163.367
R666 B.n654 B.n90 163.367
R667 B.n650 B.n648 163.367
R668 B.n646 B.n92 163.367
R669 B.n642 B.n640 163.367
R670 B.n638 B.n94 163.367
R671 B.n634 B.n632 163.367
R672 B.n630 B.n96 163.367
R673 B.n626 B.n624 163.367
R674 B.n622 B.n98 163.367
R675 B.n618 B.n616 163.367
R676 B.n614 B.n100 163.367
R677 B.n610 B.n608 163.367
R678 B.n606 B.n102 163.367
R679 B.n602 B.n600 163.367
R680 B.n598 B.n104 163.367
R681 B.n594 B.n592 163.367
R682 B.n590 B.n106 163.367
R683 B.n586 B.n584 163.367
R684 B.n582 B.n108 163.367
R685 B.n578 B.n576 163.367
R686 B.n574 B.n110 163.367
R687 B.n570 B.n568 163.367
R688 B.n468 B.n148 163.367
R689 B.n472 B.n148 163.367
R690 B.n472 B.n141 163.367
R691 B.n480 B.n141 163.367
R692 B.n480 B.n139 163.367
R693 B.n484 B.n139 163.367
R694 B.n484 B.n134 163.367
R695 B.n492 B.n134 163.367
R696 B.n492 B.n132 163.367
R697 B.n496 B.n132 163.367
R698 B.n496 B.n127 163.367
R699 B.n505 B.n127 163.367
R700 B.n505 B.n125 163.367
R701 B.n509 B.n125 163.367
R702 B.n509 B.n120 163.367
R703 B.n518 B.n120 163.367
R704 B.n518 B.n118 163.367
R705 B.n523 B.n118 163.367
R706 B.n523 B.n113 163.367
R707 B.n532 B.n113 163.367
R708 B.n533 B.n532 163.367
R709 B.n533 B.n5 163.367
R710 B.n6 B.n5 163.367
R711 B.n7 B.n6 163.367
R712 B.n539 B.n7 163.367
R713 B.n540 B.n539 163.367
R714 B.n540 B.n13 163.367
R715 B.n14 B.n13 163.367
R716 B.n15 B.n14 163.367
R717 B.n545 B.n15 163.367
R718 B.n545 B.n20 163.367
R719 B.n21 B.n20 163.367
R720 B.n22 B.n21 163.367
R721 B.n550 B.n22 163.367
R722 B.n550 B.n27 163.367
R723 B.n28 B.n27 163.367
R724 B.n29 B.n28 163.367
R725 B.n555 B.n29 163.367
R726 B.n555 B.n34 163.367
R727 B.n35 B.n34 163.367
R728 B.n36 B.n35 163.367
R729 B.n560 B.n36 163.367
R730 B.n560 B.n41 163.367
R731 B.n42 B.n41 163.367
R732 B.n43 B.n42 163.367
R733 B.n462 B.n460 163.367
R734 B.n460 B.n459 163.367
R735 B.n456 B.n455 163.367
R736 B.n453 B.n156 163.367
R737 B.n449 B.n447 163.367
R738 B.n445 B.n158 163.367
R739 B.n441 B.n439 163.367
R740 B.n437 B.n160 163.367
R741 B.n433 B.n431 163.367
R742 B.n429 B.n162 163.367
R743 B.n425 B.n423 163.367
R744 B.n421 B.n164 163.367
R745 B.n417 B.n415 163.367
R746 B.n413 B.n166 163.367
R747 B.n409 B.n407 163.367
R748 B.n405 B.n168 163.367
R749 B.n401 B.n399 163.367
R750 B.n397 B.n170 163.367
R751 B.n393 B.n391 163.367
R752 B.n389 B.n172 163.367
R753 B.n385 B.n383 163.367
R754 B.n381 B.n174 163.367
R755 B.n377 B.n375 163.367
R756 B.n373 B.n176 163.367
R757 B.n369 B.n367 163.367
R758 B.n365 B.n178 163.367
R759 B.n361 B.n359 163.367
R760 B.n357 B.n180 163.367
R761 B.n353 B.n351 163.367
R762 B.n348 B.n347 163.367
R763 B.n345 B.n186 163.367
R764 B.n341 B.n339 163.367
R765 B.n337 B.n188 163.367
R766 B.n333 B.n331 163.367
R767 B.n328 B.n327 163.367
R768 B.n325 B.n194 163.367
R769 B.n321 B.n319 163.367
R770 B.n317 B.n196 163.367
R771 B.n313 B.n311 163.367
R772 B.n309 B.n198 163.367
R773 B.n305 B.n303 163.367
R774 B.n301 B.n200 163.367
R775 B.n297 B.n295 163.367
R776 B.n293 B.n202 163.367
R777 B.n289 B.n287 163.367
R778 B.n285 B.n204 163.367
R779 B.n281 B.n279 163.367
R780 B.n277 B.n206 163.367
R781 B.n273 B.n271 163.367
R782 B.n269 B.n208 163.367
R783 B.n265 B.n263 163.367
R784 B.n261 B.n210 163.367
R785 B.n257 B.n255 163.367
R786 B.n253 B.n212 163.367
R787 B.n249 B.n247 163.367
R788 B.n245 B.n214 163.367
R789 B.n241 B.n239 163.367
R790 B.n237 B.n216 163.367
R791 B.n233 B.n231 163.367
R792 B.n229 B.n218 163.367
R793 B.n225 B.n223 163.367
R794 B.n221 B.n150 163.367
R795 B.n466 B.n146 163.367
R796 B.n474 B.n146 163.367
R797 B.n474 B.n144 163.367
R798 B.n478 B.n144 163.367
R799 B.n478 B.n138 163.367
R800 B.n486 B.n138 163.367
R801 B.n486 B.n136 163.367
R802 B.n490 B.n136 163.367
R803 B.n490 B.n130 163.367
R804 B.n499 B.n130 163.367
R805 B.n499 B.n128 163.367
R806 B.n503 B.n128 163.367
R807 B.n503 B.n123 163.367
R808 B.n512 B.n123 163.367
R809 B.n512 B.n121 163.367
R810 B.n516 B.n121 163.367
R811 B.n516 B.n116 163.367
R812 B.n526 B.n116 163.367
R813 B.n526 B.n114 163.367
R814 B.n530 B.n114 163.367
R815 B.n530 B.n3 163.367
R816 B.n860 B.n3 163.367
R817 B.n856 B.n2 163.367
R818 B.n856 B.n855 163.367
R819 B.n855 B.n9 163.367
R820 B.n851 B.n9 163.367
R821 B.n851 B.n11 163.367
R822 B.n847 B.n11 163.367
R823 B.n847 B.n16 163.367
R824 B.n843 B.n16 163.367
R825 B.n843 B.n18 163.367
R826 B.n839 B.n18 163.367
R827 B.n839 B.n23 163.367
R828 B.n835 B.n23 163.367
R829 B.n835 B.n25 163.367
R830 B.n831 B.n25 163.367
R831 B.n831 B.n31 163.367
R832 B.n827 B.n31 163.367
R833 B.n827 B.n33 163.367
R834 B.n823 B.n33 163.367
R835 B.n823 B.n38 163.367
R836 B.n819 B.n38 163.367
R837 B.n819 B.n40 163.367
R838 B.n815 B.n40 163.367
R839 B.n82 B.t8 96.964
R840 B.n189 B.t16 96.964
R841 B.n74 B.t18 96.9412
R842 B.n181 B.t13 96.9412
R843 B.n83 B.t9 73.3033
R844 B.n190 B.t15 73.3033
R845 B.n75 B.t19 73.2806
R846 B.n182 B.t12 73.2806
R847 B.n810 B.n45 71.676
R848 B.n809 B.n808 71.676
R849 B.n802 B.n47 71.676
R850 B.n801 B.n800 71.676
R851 B.n794 B.n49 71.676
R852 B.n793 B.n792 71.676
R853 B.n786 B.n51 71.676
R854 B.n785 B.n784 71.676
R855 B.n778 B.n53 71.676
R856 B.n777 B.n776 71.676
R857 B.n770 B.n55 71.676
R858 B.n769 B.n768 71.676
R859 B.n762 B.n57 71.676
R860 B.n761 B.n760 71.676
R861 B.n754 B.n59 71.676
R862 B.n753 B.n752 71.676
R863 B.n746 B.n61 71.676
R864 B.n745 B.n744 71.676
R865 B.n738 B.n63 71.676
R866 B.n737 B.n736 71.676
R867 B.n730 B.n65 71.676
R868 B.n729 B.n728 71.676
R869 B.n722 B.n67 71.676
R870 B.n721 B.n720 71.676
R871 B.n714 B.n69 71.676
R872 B.n713 B.n712 71.676
R873 B.n706 B.n71 71.676
R874 B.n705 B.n704 71.676
R875 B.n697 B.n73 71.676
R876 B.n696 B.n695 71.676
R877 B.n689 B.n77 71.676
R878 B.n688 B.n687 71.676
R879 B.n681 B.n79 71.676
R880 B.n680 B.n679 71.676
R881 B.n673 B.n81 71.676
R882 B.n672 B.n671 71.676
R883 B.n665 B.n86 71.676
R884 B.n664 B.n663 71.676
R885 B.n657 B.n88 71.676
R886 B.n656 B.n655 71.676
R887 B.n649 B.n90 71.676
R888 B.n648 B.n647 71.676
R889 B.n641 B.n92 71.676
R890 B.n640 B.n639 71.676
R891 B.n633 B.n94 71.676
R892 B.n632 B.n631 71.676
R893 B.n625 B.n96 71.676
R894 B.n624 B.n623 71.676
R895 B.n617 B.n98 71.676
R896 B.n616 B.n615 71.676
R897 B.n609 B.n100 71.676
R898 B.n608 B.n607 71.676
R899 B.n601 B.n102 71.676
R900 B.n600 B.n599 71.676
R901 B.n593 B.n104 71.676
R902 B.n592 B.n591 71.676
R903 B.n585 B.n106 71.676
R904 B.n584 B.n583 71.676
R905 B.n577 B.n108 71.676
R906 B.n576 B.n575 71.676
R907 B.n569 B.n110 71.676
R908 B.n568 B.n567 71.676
R909 B.n567 B.n566 71.676
R910 B.n570 B.n569 71.676
R911 B.n575 B.n574 71.676
R912 B.n578 B.n577 71.676
R913 B.n583 B.n582 71.676
R914 B.n586 B.n585 71.676
R915 B.n591 B.n590 71.676
R916 B.n594 B.n593 71.676
R917 B.n599 B.n598 71.676
R918 B.n602 B.n601 71.676
R919 B.n607 B.n606 71.676
R920 B.n610 B.n609 71.676
R921 B.n615 B.n614 71.676
R922 B.n618 B.n617 71.676
R923 B.n623 B.n622 71.676
R924 B.n626 B.n625 71.676
R925 B.n631 B.n630 71.676
R926 B.n634 B.n633 71.676
R927 B.n639 B.n638 71.676
R928 B.n642 B.n641 71.676
R929 B.n647 B.n646 71.676
R930 B.n650 B.n649 71.676
R931 B.n655 B.n654 71.676
R932 B.n658 B.n657 71.676
R933 B.n663 B.n662 71.676
R934 B.n666 B.n665 71.676
R935 B.n671 B.n670 71.676
R936 B.n674 B.n673 71.676
R937 B.n679 B.n678 71.676
R938 B.n682 B.n681 71.676
R939 B.n687 B.n686 71.676
R940 B.n690 B.n689 71.676
R941 B.n695 B.n694 71.676
R942 B.n698 B.n697 71.676
R943 B.n704 B.n703 71.676
R944 B.n707 B.n706 71.676
R945 B.n712 B.n711 71.676
R946 B.n715 B.n714 71.676
R947 B.n720 B.n719 71.676
R948 B.n723 B.n722 71.676
R949 B.n728 B.n727 71.676
R950 B.n731 B.n730 71.676
R951 B.n736 B.n735 71.676
R952 B.n739 B.n738 71.676
R953 B.n744 B.n743 71.676
R954 B.n747 B.n746 71.676
R955 B.n752 B.n751 71.676
R956 B.n755 B.n754 71.676
R957 B.n760 B.n759 71.676
R958 B.n763 B.n762 71.676
R959 B.n768 B.n767 71.676
R960 B.n771 B.n770 71.676
R961 B.n776 B.n775 71.676
R962 B.n779 B.n778 71.676
R963 B.n784 B.n783 71.676
R964 B.n787 B.n786 71.676
R965 B.n792 B.n791 71.676
R966 B.n795 B.n794 71.676
R967 B.n800 B.n799 71.676
R968 B.n803 B.n802 71.676
R969 B.n808 B.n807 71.676
R970 B.n811 B.n810 71.676
R971 B.n461 B.n152 71.676
R972 B.n459 B.n154 71.676
R973 B.n455 B.n454 71.676
R974 B.n448 B.n156 71.676
R975 B.n447 B.n446 71.676
R976 B.n440 B.n158 71.676
R977 B.n439 B.n438 71.676
R978 B.n432 B.n160 71.676
R979 B.n431 B.n430 71.676
R980 B.n424 B.n162 71.676
R981 B.n423 B.n422 71.676
R982 B.n416 B.n164 71.676
R983 B.n415 B.n414 71.676
R984 B.n408 B.n166 71.676
R985 B.n407 B.n406 71.676
R986 B.n400 B.n168 71.676
R987 B.n399 B.n398 71.676
R988 B.n392 B.n170 71.676
R989 B.n391 B.n390 71.676
R990 B.n384 B.n172 71.676
R991 B.n383 B.n382 71.676
R992 B.n376 B.n174 71.676
R993 B.n375 B.n374 71.676
R994 B.n368 B.n176 71.676
R995 B.n367 B.n366 71.676
R996 B.n360 B.n178 71.676
R997 B.n359 B.n358 71.676
R998 B.n352 B.n180 71.676
R999 B.n351 B.n184 71.676
R1000 B.n347 B.n346 71.676
R1001 B.n340 B.n186 71.676
R1002 B.n339 B.n338 71.676
R1003 B.n332 B.n188 71.676
R1004 B.n331 B.n192 71.676
R1005 B.n327 B.n326 71.676
R1006 B.n320 B.n194 71.676
R1007 B.n319 B.n318 71.676
R1008 B.n312 B.n196 71.676
R1009 B.n311 B.n310 71.676
R1010 B.n304 B.n198 71.676
R1011 B.n303 B.n302 71.676
R1012 B.n296 B.n200 71.676
R1013 B.n295 B.n294 71.676
R1014 B.n288 B.n202 71.676
R1015 B.n287 B.n286 71.676
R1016 B.n280 B.n204 71.676
R1017 B.n279 B.n278 71.676
R1018 B.n272 B.n206 71.676
R1019 B.n271 B.n270 71.676
R1020 B.n264 B.n208 71.676
R1021 B.n263 B.n262 71.676
R1022 B.n256 B.n210 71.676
R1023 B.n255 B.n254 71.676
R1024 B.n248 B.n212 71.676
R1025 B.n247 B.n246 71.676
R1026 B.n240 B.n214 71.676
R1027 B.n239 B.n238 71.676
R1028 B.n232 B.n216 71.676
R1029 B.n231 B.n230 71.676
R1030 B.n224 B.n218 71.676
R1031 B.n223 B.n222 71.676
R1032 B.n462 B.n461 71.676
R1033 B.n456 B.n154 71.676
R1034 B.n454 B.n453 71.676
R1035 B.n449 B.n448 71.676
R1036 B.n446 B.n445 71.676
R1037 B.n441 B.n440 71.676
R1038 B.n438 B.n437 71.676
R1039 B.n433 B.n432 71.676
R1040 B.n430 B.n429 71.676
R1041 B.n425 B.n424 71.676
R1042 B.n422 B.n421 71.676
R1043 B.n417 B.n416 71.676
R1044 B.n414 B.n413 71.676
R1045 B.n409 B.n408 71.676
R1046 B.n406 B.n405 71.676
R1047 B.n401 B.n400 71.676
R1048 B.n398 B.n397 71.676
R1049 B.n393 B.n392 71.676
R1050 B.n390 B.n389 71.676
R1051 B.n385 B.n384 71.676
R1052 B.n382 B.n381 71.676
R1053 B.n377 B.n376 71.676
R1054 B.n374 B.n373 71.676
R1055 B.n369 B.n368 71.676
R1056 B.n366 B.n365 71.676
R1057 B.n361 B.n360 71.676
R1058 B.n358 B.n357 71.676
R1059 B.n353 B.n352 71.676
R1060 B.n348 B.n184 71.676
R1061 B.n346 B.n345 71.676
R1062 B.n341 B.n340 71.676
R1063 B.n338 B.n337 71.676
R1064 B.n333 B.n332 71.676
R1065 B.n328 B.n192 71.676
R1066 B.n326 B.n325 71.676
R1067 B.n321 B.n320 71.676
R1068 B.n318 B.n317 71.676
R1069 B.n313 B.n312 71.676
R1070 B.n310 B.n309 71.676
R1071 B.n305 B.n304 71.676
R1072 B.n302 B.n301 71.676
R1073 B.n297 B.n296 71.676
R1074 B.n294 B.n293 71.676
R1075 B.n289 B.n288 71.676
R1076 B.n286 B.n285 71.676
R1077 B.n281 B.n280 71.676
R1078 B.n278 B.n277 71.676
R1079 B.n273 B.n272 71.676
R1080 B.n270 B.n269 71.676
R1081 B.n265 B.n264 71.676
R1082 B.n262 B.n261 71.676
R1083 B.n257 B.n256 71.676
R1084 B.n254 B.n253 71.676
R1085 B.n249 B.n248 71.676
R1086 B.n246 B.n245 71.676
R1087 B.n241 B.n240 71.676
R1088 B.n238 B.n237 71.676
R1089 B.n233 B.n232 71.676
R1090 B.n230 B.n229 71.676
R1091 B.n225 B.n224 71.676
R1092 B.n222 B.n221 71.676
R1093 B.n861 B.n860 71.676
R1094 B.n861 B.n2 71.676
R1095 B.n700 B.n75 59.5399
R1096 B.n84 B.n83 59.5399
R1097 B.n191 B.n190 59.5399
R1098 B.n183 B.n182 59.5399
R1099 B.n467 B.n151 58.9334
R1100 B.n816 B.n44 58.9334
R1101 B.n467 B.n147 33.1198
R1102 B.n473 B.n147 33.1198
R1103 B.n473 B.n142 33.1198
R1104 B.n479 B.n142 33.1198
R1105 B.n479 B.n143 33.1198
R1106 B.n485 B.n135 33.1198
R1107 B.n491 B.n135 33.1198
R1108 B.n491 B.n131 33.1198
R1109 B.n498 B.n131 33.1198
R1110 B.n498 B.n497 33.1198
R1111 B.n504 B.n124 33.1198
R1112 B.n511 B.n124 33.1198
R1113 B.n511 B.n510 33.1198
R1114 B.n517 B.n117 33.1198
R1115 B.n525 B.n117 33.1198
R1116 B.n525 B.n524 33.1198
R1117 B.n531 B.n4 33.1198
R1118 B.n859 B.n4 33.1198
R1119 B.n859 B.n858 33.1198
R1120 B.n858 B.n857 33.1198
R1121 B.n857 B.n8 33.1198
R1122 B.n850 B.n12 33.1198
R1123 B.n850 B.n849 33.1198
R1124 B.n849 B.n848 33.1198
R1125 B.n842 B.n19 33.1198
R1126 B.n842 B.n841 33.1198
R1127 B.n841 B.n840 33.1198
R1128 B.n834 B.n26 33.1198
R1129 B.n834 B.n833 33.1198
R1130 B.n833 B.n832 33.1198
R1131 B.n832 B.n30 33.1198
R1132 B.n826 B.n30 33.1198
R1133 B.n825 B.n824 33.1198
R1134 B.n824 B.n37 33.1198
R1135 B.n818 B.n37 33.1198
R1136 B.n818 B.n817 33.1198
R1137 B.n817 B.n816 33.1198
R1138 B.n465 B.n464 32.3127
R1139 B.n469 B.n149 32.3127
R1140 B.n565 B.n564 32.3127
R1141 B.n814 B.n813 32.3127
R1142 B.n497 B.t2 30.6846
R1143 B.n26 B.t5 30.6846
R1144 B.n531 B.t4 29.7105
R1145 B.t0 B.n8 29.7105
R1146 B.n485 B.t11 28.7364
R1147 B.n826 B.t7 28.7364
R1148 B.n75 B.n74 23.6611
R1149 B.n83 B.n82 23.6611
R1150 B.n190 B.n189 23.6611
R1151 B.n182 B.n181 23.6611
R1152 B B.n862 18.0485
R1153 B.n510 B.t1 17.0472
R1154 B.n19 B.t3 17.0472
R1155 B.n517 B.t1 16.0731
R1156 B.n848 B.t3 16.0731
R1157 B.n465 B.n145 10.6151
R1158 B.n475 B.n145 10.6151
R1159 B.n476 B.n475 10.6151
R1160 B.n477 B.n476 10.6151
R1161 B.n477 B.n137 10.6151
R1162 B.n487 B.n137 10.6151
R1163 B.n488 B.n487 10.6151
R1164 B.n489 B.n488 10.6151
R1165 B.n489 B.n129 10.6151
R1166 B.n500 B.n129 10.6151
R1167 B.n501 B.n500 10.6151
R1168 B.n502 B.n501 10.6151
R1169 B.n502 B.n122 10.6151
R1170 B.n513 B.n122 10.6151
R1171 B.n514 B.n513 10.6151
R1172 B.n515 B.n514 10.6151
R1173 B.n515 B.n115 10.6151
R1174 B.n527 B.n115 10.6151
R1175 B.n528 B.n527 10.6151
R1176 B.n529 B.n528 10.6151
R1177 B.n529 B.n0 10.6151
R1178 B.n464 B.n463 10.6151
R1179 B.n463 B.n153 10.6151
R1180 B.n458 B.n153 10.6151
R1181 B.n458 B.n457 10.6151
R1182 B.n457 B.n155 10.6151
R1183 B.n452 B.n155 10.6151
R1184 B.n452 B.n451 10.6151
R1185 B.n451 B.n450 10.6151
R1186 B.n450 B.n157 10.6151
R1187 B.n444 B.n157 10.6151
R1188 B.n444 B.n443 10.6151
R1189 B.n443 B.n442 10.6151
R1190 B.n442 B.n159 10.6151
R1191 B.n436 B.n159 10.6151
R1192 B.n436 B.n435 10.6151
R1193 B.n435 B.n434 10.6151
R1194 B.n434 B.n161 10.6151
R1195 B.n428 B.n161 10.6151
R1196 B.n428 B.n427 10.6151
R1197 B.n427 B.n426 10.6151
R1198 B.n426 B.n163 10.6151
R1199 B.n420 B.n163 10.6151
R1200 B.n420 B.n419 10.6151
R1201 B.n419 B.n418 10.6151
R1202 B.n418 B.n165 10.6151
R1203 B.n412 B.n165 10.6151
R1204 B.n412 B.n411 10.6151
R1205 B.n411 B.n410 10.6151
R1206 B.n410 B.n167 10.6151
R1207 B.n404 B.n167 10.6151
R1208 B.n404 B.n403 10.6151
R1209 B.n403 B.n402 10.6151
R1210 B.n402 B.n169 10.6151
R1211 B.n396 B.n169 10.6151
R1212 B.n396 B.n395 10.6151
R1213 B.n395 B.n394 10.6151
R1214 B.n394 B.n171 10.6151
R1215 B.n388 B.n171 10.6151
R1216 B.n388 B.n387 10.6151
R1217 B.n387 B.n386 10.6151
R1218 B.n386 B.n173 10.6151
R1219 B.n380 B.n173 10.6151
R1220 B.n380 B.n379 10.6151
R1221 B.n379 B.n378 10.6151
R1222 B.n378 B.n175 10.6151
R1223 B.n372 B.n175 10.6151
R1224 B.n372 B.n371 10.6151
R1225 B.n371 B.n370 10.6151
R1226 B.n370 B.n177 10.6151
R1227 B.n364 B.n177 10.6151
R1228 B.n364 B.n363 10.6151
R1229 B.n363 B.n362 10.6151
R1230 B.n362 B.n179 10.6151
R1231 B.n356 B.n179 10.6151
R1232 B.n356 B.n355 10.6151
R1233 B.n355 B.n354 10.6151
R1234 B.n350 B.n349 10.6151
R1235 B.n349 B.n185 10.6151
R1236 B.n344 B.n185 10.6151
R1237 B.n344 B.n343 10.6151
R1238 B.n343 B.n342 10.6151
R1239 B.n342 B.n187 10.6151
R1240 B.n336 B.n187 10.6151
R1241 B.n336 B.n335 10.6151
R1242 B.n335 B.n334 10.6151
R1243 B.n330 B.n329 10.6151
R1244 B.n329 B.n193 10.6151
R1245 B.n324 B.n193 10.6151
R1246 B.n324 B.n323 10.6151
R1247 B.n323 B.n322 10.6151
R1248 B.n322 B.n195 10.6151
R1249 B.n316 B.n195 10.6151
R1250 B.n316 B.n315 10.6151
R1251 B.n315 B.n314 10.6151
R1252 B.n314 B.n197 10.6151
R1253 B.n308 B.n197 10.6151
R1254 B.n308 B.n307 10.6151
R1255 B.n307 B.n306 10.6151
R1256 B.n306 B.n199 10.6151
R1257 B.n300 B.n199 10.6151
R1258 B.n300 B.n299 10.6151
R1259 B.n299 B.n298 10.6151
R1260 B.n298 B.n201 10.6151
R1261 B.n292 B.n201 10.6151
R1262 B.n292 B.n291 10.6151
R1263 B.n291 B.n290 10.6151
R1264 B.n290 B.n203 10.6151
R1265 B.n284 B.n203 10.6151
R1266 B.n284 B.n283 10.6151
R1267 B.n283 B.n282 10.6151
R1268 B.n282 B.n205 10.6151
R1269 B.n276 B.n205 10.6151
R1270 B.n276 B.n275 10.6151
R1271 B.n275 B.n274 10.6151
R1272 B.n274 B.n207 10.6151
R1273 B.n268 B.n207 10.6151
R1274 B.n268 B.n267 10.6151
R1275 B.n267 B.n266 10.6151
R1276 B.n266 B.n209 10.6151
R1277 B.n260 B.n209 10.6151
R1278 B.n260 B.n259 10.6151
R1279 B.n259 B.n258 10.6151
R1280 B.n258 B.n211 10.6151
R1281 B.n252 B.n211 10.6151
R1282 B.n252 B.n251 10.6151
R1283 B.n251 B.n250 10.6151
R1284 B.n250 B.n213 10.6151
R1285 B.n244 B.n213 10.6151
R1286 B.n244 B.n243 10.6151
R1287 B.n243 B.n242 10.6151
R1288 B.n242 B.n215 10.6151
R1289 B.n236 B.n215 10.6151
R1290 B.n236 B.n235 10.6151
R1291 B.n235 B.n234 10.6151
R1292 B.n234 B.n217 10.6151
R1293 B.n228 B.n217 10.6151
R1294 B.n228 B.n227 10.6151
R1295 B.n227 B.n226 10.6151
R1296 B.n226 B.n219 10.6151
R1297 B.n220 B.n219 10.6151
R1298 B.n220 B.n149 10.6151
R1299 B.n470 B.n469 10.6151
R1300 B.n471 B.n470 10.6151
R1301 B.n471 B.n140 10.6151
R1302 B.n481 B.n140 10.6151
R1303 B.n482 B.n481 10.6151
R1304 B.n483 B.n482 10.6151
R1305 B.n483 B.n133 10.6151
R1306 B.n493 B.n133 10.6151
R1307 B.n494 B.n493 10.6151
R1308 B.n495 B.n494 10.6151
R1309 B.n495 B.n126 10.6151
R1310 B.n506 B.n126 10.6151
R1311 B.n507 B.n506 10.6151
R1312 B.n508 B.n507 10.6151
R1313 B.n508 B.n119 10.6151
R1314 B.n519 B.n119 10.6151
R1315 B.n520 B.n519 10.6151
R1316 B.n522 B.n520 10.6151
R1317 B.n522 B.n521 10.6151
R1318 B.n521 B.n112 10.6151
R1319 B.n534 B.n112 10.6151
R1320 B.n535 B.n534 10.6151
R1321 B.n536 B.n535 10.6151
R1322 B.n537 B.n536 10.6151
R1323 B.n538 B.n537 10.6151
R1324 B.n541 B.n538 10.6151
R1325 B.n542 B.n541 10.6151
R1326 B.n543 B.n542 10.6151
R1327 B.n544 B.n543 10.6151
R1328 B.n546 B.n544 10.6151
R1329 B.n547 B.n546 10.6151
R1330 B.n548 B.n547 10.6151
R1331 B.n549 B.n548 10.6151
R1332 B.n551 B.n549 10.6151
R1333 B.n552 B.n551 10.6151
R1334 B.n553 B.n552 10.6151
R1335 B.n554 B.n553 10.6151
R1336 B.n556 B.n554 10.6151
R1337 B.n557 B.n556 10.6151
R1338 B.n558 B.n557 10.6151
R1339 B.n559 B.n558 10.6151
R1340 B.n561 B.n559 10.6151
R1341 B.n562 B.n561 10.6151
R1342 B.n563 B.n562 10.6151
R1343 B.n564 B.n563 10.6151
R1344 B.n854 B.n1 10.6151
R1345 B.n854 B.n853 10.6151
R1346 B.n853 B.n852 10.6151
R1347 B.n852 B.n10 10.6151
R1348 B.n846 B.n10 10.6151
R1349 B.n846 B.n845 10.6151
R1350 B.n845 B.n844 10.6151
R1351 B.n844 B.n17 10.6151
R1352 B.n838 B.n17 10.6151
R1353 B.n838 B.n837 10.6151
R1354 B.n837 B.n836 10.6151
R1355 B.n836 B.n24 10.6151
R1356 B.n830 B.n24 10.6151
R1357 B.n830 B.n829 10.6151
R1358 B.n829 B.n828 10.6151
R1359 B.n828 B.n32 10.6151
R1360 B.n822 B.n32 10.6151
R1361 B.n822 B.n821 10.6151
R1362 B.n821 B.n820 10.6151
R1363 B.n820 B.n39 10.6151
R1364 B.n814 B.n39 10.6151
R1365 B.n813 B.n812 10.6151
R1366 B.n812 B.n46 10.6151
R1367 B.n806 B.n46 10.6151
R1368 B.n806 B.n805 10.6151
R1369 B.n805 B.n804 10.6151
R1370 B.n804 B.n48 10.6151
R1371 B.n798 B.n48 10.6151
R1372 B.n798 B.n797 10.6151
R1373 B.n797 B.n796 10.6151
R1374 B.n796 B.n50 10.6151
R1375 B.n790 B.n50 10.6151
R1376 B.n790 B.n789 10.6151
R1377 B.n789 B.n788 10.6151
R1378 B.n788 B.n52 10.6151
R1379 B.n782 B.n52 10.6151
R1380 B.n782 B.n781 10.6151
R1381 B.n781 B.n780 10.6151
R1382 B.n780 B.n54 10.6151
R1383 B.n774 B.n54 10.6151
R1384 B.n774 B.n773 10.6151
R1385 B.n773 B.n772 10.6151
R1386 B.n772 B.n56 10.6151
R1387 B.n766 B.n56 10.6151
R1388 B.n766 B.n765 10.6151
R1389 B.n765 B.n764 10.6151
R1390 B.n764 B.n58 10.6151
R1391 B.n758 B.n58 10.6151
R1392 B.n758 B.n757 10.6151
R1393 B.n757 B.n756 10.6151
R1394 B.n756 B.n60 10.6151
R1395 B.n750 B.n60 10.6151
R1396 B.n750 B.n749 10.6151
R1397 B.n749 B.n748 10.6151
R1398 B.n748 B.n62 10.6151
R1399 B.n742 B.n62 10.6151
R1400 B.n742 B.n741 10.6151
R1401 B.n741 B.n740 10.6151
R1402 B.n740 B.n64 10.6151
R1403 B.n734 B.n64 10.6151
R1404 B.n734 B.n733 10.6151
R1405 B.n733 B.n732 10.6151
R1406 B.n732 B.n66 10.6151
R1407 B.n726 B.n66 10.6151
R1408 B.n726 B.n725 10.6151
R1409 B.n725 B.n724 10.6151
R1410 B.n724 B.n68 10.6151
R1411 B.n718 B.n68 10.6151
R1412 B.n718 B.n717 10.6151
R1413 B.n717 B.n716 10.6151
R1414 B.n716 B.n70 10.6151
R1415 B.n710 B.n70 10.6151
R1416 B.n710 B.n709 10.6151
R1417 B.n709 B.n708 10.6151
R1418 B.n708 B.n72 10.6151
R1419 B.n702 B.n72 10.6151
R1420 B.n702 B.n701 10.6151
R1421 B.n699 B.n76 10.6151
R1422 B.n693 B.n76 10.6151
R1423 B.n693 B.n692 10.6151
R1424 B.n692 B.n691 10.6151
R1425 B.n691 B.n78 10.6151
R1426 B.n685 B.n78 10.6151
R1427 B.n685 B.n684 10.6151
R1428 B.n684 B.n683 10.6151
R1429 B.n683 B.n80 10.6151
R1430 B.n677 B.n676 10.6151
R1431 B.n676 B.n675 10.6151
R1432 B.n675 B.n85 10.6151
R1433 B.n669 B.n85 10.6151
R1434 B.n669 B.n668 10.6151
R1435 B.n668 B.n667 10.6151
R1436 B.n667 B.n87 10.6151
R1437 B.n661 B.n87 10.6151
R1438 B.n661 B.n660 10.6151
R1439 B.n660 B.n659 10.6151
R1440 B.n659 B.n89 10.6151
R1441 B.n653 B.n89 10.6151
R1442 B.n653 B.n652 10.6151
R1443 B.n652 B.n651 10.6151
R1444 B.n651 B.n91 10.6151
R1445 B.n645 B.n91 10.6151
R1446 B.n645 B.n644 10.6151
R1447 B.n644 B.n643 10.6151
R1448 B.n643 B.n93 10.6151
R1449 B.n637 B.n93 10.6151
R1450 B.n637 B.n636 10.6151
R1451 B.n636 B.n635 10.6151
R1452 B.n635 B.n95 10.6151
R1453 B.n629 B.n95 10.6151
R1454 B.n629 B.n628 10.6151
R1455 B.n628 B.n627 10.6151
R1456 B.n627 B.n97 10.6151
R1457 B.n621 B.n97 10.6151
R1458 B.n621 B.n620 10.6151
R1459 B.n620 B.n619 10.6151
R1460 B.n619 B.n99 10.6151
R1461 B.n613 B.n99 10.6151
R1462 B.n613 B.n612 10.6151
R1463 B.n612 B.n611 10.6151
R1464 B.n611 B.n101 10.6151
R1465 B.n605 B.n101 10.6151
R1466 B.n605 B.n604 10.6151
R1467 B.n604 B.n603 10.6151
R1468 B.n603 B.n103 10.6151
R1469 B.n597 B.n103 10.6151
R1470 B.n597 B.n596 10.6151
R1471 B.n596 B.n595 10.6151
R1472 B.n595 B.n105 10.6151
R1473 B.n589 B.n105 10.6151
R1474 B.n589 B.n588 10.6151
R1475 B.n588 B.n587 10.6151
R1476 B.n587 B.n107 10.6151
R1477 B.n581 B.n107 10.6151
R1478 B.n581 B.n580 10.6151
R1479 B.n580 B.n579 10.6151
R1480 B.n579 B.n109 10.6151
R1481 B.n573 B.n109 10.6151
R1482 B.n573 B.n572 10.6151
R1483 B.n572 B.n571 10.6151
R1484 B.n571 B.n111 10.6151
R1485 B.n565 B.n111 10.6151
R1486 B.n354 B.n183 9.36635
R1487 B.n330 B.n191 9.36635
R1488 B.n701 B.n700 9.36635
R1489 B.n677 B.n84 9.36635
R1490 B.n862 B.n0 8.11757
R1491 B.n862 B.n1 8.11757
R1492 B.n143 B.t11 4.38394
R1493 B.t7 B.n825 4.38394
R1494 B.n524 B.t4 3.40984
R1495 B.n12 B.t0 3.40984
R1496 B.n504 B.t2 2.43574
R1497 B.n840 B.t5 2.43574
R1498 B.n350 B.n183 1.24928
R1499 B.n334 B.n191 1.24928
R1500 B.n700 B.n699 1.24928
R1501 B.n84 B.n80 1.24928
R1502 VP.n5 VP.t1 529.992
R1503 VP.n12 VP.t5 513.14
R1504 VP.n19 VP.t3 513.14
R1505 VP.n9 VP.t4 513.14
R1506 VP.n1 VP.t0 468.731
R1507 VP.n4 VP.t2 468.731
R1508 VP.n20 VP.n19 161.3
R1509 VP.n7 VP.n6 161.3
R1510 VP.n8 VP.n3 161.3
R1511 VP.n10 VP.n9 161.3
R1512 VP.n18 VP.n0 161.3
R1513 VP.n17 VP.n16 161.3
R1514 VP.n15 VP.n14 161.3
R1515 VP.n13 VP.n2 161.3
R1516 VP.n12 VP.n11 161.3
R1517 VP.n14 VP.n13 54.0911
R1518 VP.n18 VP.n17 54.0911
R1519 VP.n8 VP.n7 54.0911
R1520 VP.n11 VP.n10 45.9702
R1521 VP.n6 VP.n5 43.6035
R1522 VP.n5 VP.n4 42.5728
R1523 VP.n14 VP.n1 12.234
R1524 VP.n17 VP.n1 12.234
R1525 VP.n7 VP.n4 12.234
R1526 VP.n13 VP.n12 3.65202
R1527 VP.n19 VP.n18 3.65202
R1528 VP.n9 VP.n8 3.65202
R1529 VP.n6 VP.n3 0.189894
R1530 VP.n10 VP.n3 0.189894
R1531 VP.n11 VP.n2 0.189894
R1532 VP.n15 VP.n2 0.189894
R1533 VP.n16 VP.n15 0.189894
R1534 VP.n16 VP.n0 0.189894
R1535 VP.n20 VP.n0 0.189894
R1536 VP VP.n20 0.0516364
R1537 VDD1 VDD1.t4 65.6019
R1538 VDD1.n1 VDD1.t0 65.4883
R1539 VDD1.n1 VDD1.n0 63.8185
R1540 VDD1.n3 VDD1.n2 63.611
R1541 VDD1.n3 VDD1.n1 43.1647
R1542 VDD1.n2 VDD1.t3 1.14435
R1543 VDD1.n2 VDD1.t1 1.14435
R1544 VDD1.n0 VDD1.t5 1.14435
R1545 VDD1.n0 VDD1.t2 1.14435
R1546 VDD1 VDD1.n3 0.205241
C0 VN VP 6.24896f
C1 VDD1 VP 7.00046f
C2 VTAIL VDD2 12.3151f
C3 VN VDD2 6.84044f
C4 VTAIL VN 6.36537f
C5 VDD1 VDD2 0.7813f
C6 VDD2 VP 0.314407f
C7 VDD1 VTAIL 12.2817f
C8 VTAIL VP 6.38012f
C9 VDD1 VN 0.148408f
C10 VDD2 B 5.588265f
C11 VDD1 B 5.831073f
C12 VTAIL B 8.539495f
C13 VN B 8.795229f
C14 VP B 6.695338f
C15 VDD1.t4 B 3.6144f
C16 VDD1.t0 B 3.61376f
C17 VDD1.t5 B 0.310141f
C18 VDD1.t2 B 0.310141f
C19 VDD1.n0 B 2.82476f
C20 VDD1.n1 B 2.33432f
C21 VDD1.t3 B 0.310141f
C22 VDD1.t1 B 0.310141f
C23 VDD1.n2 B 2.82381f
C24 VDD1.n3 B 2.46036f
C25 VP.n0 B 0.041817f
C26 VP.t0 B 1.77065f
C27 VP.n1 B 0.640283f
C28 VP.n2 B 0.041817f
C29 VP.n3 B 0.041817f
C30 VP.t4 B 1.82767f
C31 VP.t2 B 1.77065f
C32 VP.n4 B 0.679118f
C33 VP.t1 B 1.84978f
C34 VP.n5 B 0.690889f
C35 VP.n6 B 0.174917f
C36 VP.n7 B 0.054058f
C37 VP.n8 B 0.013523f
C38 VP.n9 B 0.683394f
C39 VP.n10 B 1.99784f
C40 VP.n11 B 2.03054f
C41 VP.t5 B 1.82767f
C42 VP.n12 B 0.683394f
C43 VP.n13 B 0.013523f
C44 VP.n14 B 0.054058f
C45 VP.n15 B 0.041817f
C46 VP.n16 B 0.041817f
C47 VP.n17 B 0.054058f
C48 VP.n18 B 0.013523f
C49 VP.t3 B 1.82767f
C50 VP.n19 B 0.683394f
C51 VP.n20 B 0.032406f
C52 VDD2.t0 B 3.59189f
C53 VDD2.t3 B 0.308265f
C54 VDD2.t4 B 0.308265f
C55 VDD2.n0 B 2.80767f
C56 VDD2.n1 B 2.24514f
C57 VDD2.t5 B 3.58848f
C58 VDD2.n2 B 2.46653f
C59 VDD2.t1 B 0.308265f
C60 VDD2.t2 B 0.308265f
C61 VDD2.n3 B 2.80764f
C62 VTAIL.t7 B 0.316512f
C63 VTAIL.t8 B 0.316512f
C64 VTAIL.n0 B 2.81633f
C65 VTAIL.n1 B 0.320938f
C66 VTAIL.t4 B 3.59952f
C67 VTAIL.n2 B 0.455434f
C68 VTAIL.t2 B 0.316512f
C69 VTAIL.t1 B 0.316512f
C70 VTAIL.n3 B 2.81633f
C71 VTAIL.n4 B 1.8849f
C72 VTAIL.t6 B 0.316512f
C73 VTAIL.t11 B 0.316512f
C74 VTAIL.n5 B 2.81633f
C75 VTAIL.n6 B 1.8849f
C76 VTAIL.t9 B 3.59954f
C77 VTAIL.n7 B 0.455414f
C78 VTAIL.t0 B 0.316512f
C79 VTAIL.t3 B 0.316512f
C80 VTAIL.n8 B 2.81633f
C81 VTAIL.n9 B 0.375407f
C82 VTAIL.t5 B 3.59952f
C83 VTAIL.n10 B 1.88651f
C84 VTAIL.t10 B 3.59952f
C85 VTAIL.n11 B 1.86257f
C86 VN.n0 B 0.041266f
C87 VN.t2 B 1.74734f
C88 VN.n1 B 0.670178f
C89 VN.t5 B 1.82543f
C90 VN.n2 B 0.681795f
C91 VN.n3 B 0.172615f
C92 VN.n4 B 0.053346f
C93 VN.n5 B 0.013345f
C94 VN.t1 B 1.80361f
C95 VN.n6 B 0.674398f
C96 VN.n7 B 0.03198f
C97 VN.n8 B 0.041266f
C98 VN.t4 B 1.74734f
C99 VN.n9 B 0.670178f
C100 VN.t3 B 1.82543f
C101 VN.n10 B 0.681795f
C102 VN.n11 B 0.172615f
C103 VN.n12 B 0.053346f
C104 VN.n13 B 0.013345f
C105 VN.t0 B 1.80361f
C106 VN.n14 B 0.674398f
C107 VN.n15 B 1.99849f
.ends

