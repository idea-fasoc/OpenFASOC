* NGSPICE file created from diff_pair_sample_0897.ext - technology: sky130A

.subckt diff_pair_sample_0897 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t1 w_n2200_n3844# sky130_fd_pr__pfet_01v8 ad=5.6082 pd=29.54 as=2.3727 ps=14.71 w=14.38 l=1.72
X1 B.t11 B.t9 B.t10 w_n2200_n3844# sky130_fd_pr__pfet_01v8 ad=5.6082 pd=29.54 as=0 ps=0 w=14.38 l=1.72
X2 VTAIL.t1 VN.t0 VDD2.t3 w_n2200_n3844# sky130_fd_pr__pfet_01v8 ad=5.6082 pd=29.54 as=2.3727 ps=14.71 w=14.38 l=1.72
X3 B.t8 B.t6 B.t7 w_n2200_n3844# sky130_fd_pr__pfet_01v8 ad=5.6082 pd=29.54 as=0 ps=0 w=14.38 l=1.72
X4 VDD2.t2 VN.t1 VTAIL.t3 w_n2200_n3844# sky130_fd_pr__pfet_01v8 ad=2.3727 pd=14.71 as=5.6082 ps=29.54 w=14.38 l=1.72
X5 VDD1.t0 VP.t1 VTAIL.t6 w_n2200_n3844# sky130_fd_pr__pfet_01v8 ad=2.3727 pd=14.71 as=5.6082 ps=29.54 w=14.38 l=1.72
X6 VDD1.t3 VP.t2 VTAIL.t5 w_n2200_n3844# sky130_fd_pr__pfet_01v8 ad=2.3727 pd=14.71 as=5.6082 ps=29.54 w=14.38 l=1.72
X7 VDD2.t1 VN.t2 VTAIL.t2 w_n2200_n3844# sky130_fd_pr__pfet_01v8 ad=2.3727 pd=14.71 as=5.6082 ps=29.54 w=14.38 l=1.72
X8 VTAIL.t4 VP.t3 VDD1.t2 w_n2200_n3844# sky130_fd_pr__pfet_01v8 ad=5.6082 pd=29.54 as=2.3727 ps=14.71 w=14.38 l=1.72
X9 B.t5 B.t3 B.t4 w_n2200_n3844# sky130_fd_pr__pfet_01v8 ad=5.6082 pd=29.54 as=0 ps=0 w=14.38 l=1.72
X10 B.t2 B.t0 B.t1 w_n2200_n3844# sky130_fd_pr__pfet_01v8 ad=5.6082 pd=29.54 as=0 ps=0 w=14.38 l=1.72
X11 VTAIL.t0 VN.t3 VDD2.t0 w_n2200_n3844# sky130_fd_pr__pfet_01v8 ad=5.6082 pd=29.54 as=2.3727 ps=14.71 w=14.38 l=1.72
R0 VP.n3 VP.t0 236.756
R1 VP.n3 VP.t2 236.333
R2 VP.n5 VP.t3 201.488
R3 VP.n13 VP.t1 201.488
R4 VP.n5 VP.n4 184.427
R5 VP.n14 VP.n13 184.427
R6 VP.n12 VP.n0 161.3
R7 VP.n11 VP.n10 161.3
R8 VP.n9 VP.n1 161.3
R9 VP.n8 VP.n7 161.3
R10 VP.n6 VP.n2 161.3
R11 VP.n4 VP.n3 54.8003
R12 VP.n7 VP.n1 40.4106
R13 VP.n11 VP.n1 40.4106
R14 VP.n7 VP.n6 24.3439
R15 VP.n12 VP.n11 24.3439
R16 VP.n6 VP.n5 1.21767
R17 VP.n13 VP.n12 1.21767
R18 VP.n4 VP.n2 0.189894
R19 VP.n8 VP.n2 0.189894
R20 VP.n9 VP.n8 0.189894
R21 VP.n10 VP.n9 0.189894
R22 VP.n10 VP.n0 0.189894
R23 VP.n14 VP.n0 0.189894
R24 VP VP.n14 0.0516364
R25 VDD1 VDD1.n1 114.919
R26 VDD1 VDD1.n0 73.04
R27 VDD1.n0 VDD1.t1 2.26093
R28 VDD1.n0 VDD1.t3 2.26093
R29 VDD1.n1 VDD1.t2 2.26093
R30 VDD1.n1 VDD1.t0 2.26093
R31 VTAIL.n5 VTAIL.t7 58.5636
R32 VTAIL.n4 VTAIL.t3 58.5636
R33 VTAIL.n3 VTAIL.t0 58.5636
R34 VTAIL.n7 VTAIL.t2 58.5634
R35 VTAIL.n0 VTAIL.t1 58.5634
R36 VTAIL.n1 VTAIL.t6 58.5634
R37 VTAIL.n2 VTAIL.t4 58.5634
R38 VTAIL.n6 VTAIL.t5 58.5634
R39 VTAIL.n7 VTAIL.n6 26.5307
R40 VTAIL.n3 VTAIL.n2 26.5307
R41 VTAIL.n4 VTAIL.n3 1.76774
R42 VTAIL.n6 VTAIL.n5 1.76774
R43 VTAIL.n2 VTAIL.n1 1.76774
R44 VTAIL VTAIL.n0 0.94231
R45 VTAIL VTAIL.n7 0.825931
R46 VTAIL.n5 VTAIL.n4 0.470328
R47 VTAIL.n1 VTAIL.n0 0.470328
R48 B.n450 B.n449 585
R49 B.n451 B.n72 585
R50 B.n453 B.n452 585
R51 B.n454 B.n71 585
R52 B.n456 B.n455 585
R53 B.n457 B.n70 585
R54 B.n459 B.n458 585
R55 B.n460 B.n69 585
R56 B.n462 B.n461 585
R57 B.n463 B.n68 585
R58 B.n465 B.n464 585
R59 B.n466 B.n67 585
R60 B.n468 B.n467 585
R61 B.n469 B.n66 585
R62 B.n471 B.n470 585
R63 B.n472 B.n65 585
R64 B.n474 B.n473 585
R65 B.n475 B.n64 585
R66 B.n477 B.n476 585
R67 B.n478 B.n63 585
R68 B.n480 B.n479 585
R69 B.n481 B.n62 585
R70 B.n483 B.n482 585
R71 B.n484 B.n61 585
R72 B.n486 B.n485 585
R73 B.n487 B.n60 585
R74 B.n489 B.n488 585
R75 B.n490 B.n59 585
R76 B.n492 B.n491 585
R77 B.n493 B.n58 585
R78 B.n495 B.n494 585
R79 B.n496 B.n57 585
R80 B.n498 B.n497 585
R81 B.n499 B.n56 585
R82 B.n501 B.n500 585
R83 B.n502 B.n55 585
R84 B.n504 B.n503 585
R85 B.n505 B.n54 585
R86 B.n507 B.n506 585
R87 B.n508 B.n53 585
R88 B.n510 B.n509 585
R89 B.n511 B.n52 585
R90 B.n513 B.n512 585
R91 B.n514 B.n51 585
R92 B.n516 B.n515 585
R93 B.n517 B.n50 585
R94 B.n519 B.n518 585
R95 B.n520 B.n49 585
R96 B.n522 B.n521 585
R97 B.n524 B.n523 585
R98 B.n525 B.n45 585
R99 B.n527 B.n526 585
R100 B.n528 B.n44 585
R101 B.n530 B.n529 585
R102 B.n531 B.n43 585
R103 B.n533 B.n532 585
R104 B.n534 B.n42 585
R105 B.n536 B.n535 585
R106 B.n538 B.n39 585
R107 B.n540 B.n539 585
R108 B.n541 B.n38 585
R109 B.n543 B.n542 585
R110 B.n544 B.n37 585
R111 B.n546 B.n545 585
R112 B.n547 B.n36 585
R113 B.n549 B.n548 585
R114 B.n550 B.n35 585
R115 B.n552 B.n551 585
R116 B.n553 B.n34 585
R117 B.n555 B.n554 585
R118 B.n556 B.n33 585
R119 B.n558 B.n557 585
R120 B.n559 B.n32 585
R121 B.n561 B.n560 585
R122 B.n562 B.n31 585
R123 B.n564 B.n563 585
R124 B.n565 B.n30 585
R125 B.n567 B.n566 585
R126 B.n568 B.n29 585
R127 B.n570 B.n569 585
R128 B.n571 B.n28 585
R129 B.n573 B.n572 585
R130 B.n574 B.n27 585
R131 B.n576 B.n575 585
R132 B.n577 B.n26 585
R133 B.n579 B.n578 585
R134 B.n580 B.n25 585
R135 B.n582 B.n581 585
R136 B.n583 B.n24 585
R137 B.n585 B.n584 585
R138 B.n586 B.n23 585
R139 B.n588 B.n587 585
R140 B.n589 B.n22 585
R141 B.n591 B.n590 585
R142 B.n592 B.n21 585
R143 B.n594 B.n593 585
R144 B.n595 B.n20 585
R145 B.n597 B.n596 585
R146 B.n598 B.n19 585
R147 B.n600 B.n599 585
R148 B.n601 B.n18 585
R149 B.n603 B.n602 585
R150 B.n604 B.n17 585
R151 B.n606 B.n605 585
R152 B.n607 B.n16 585
R153 B.n609 B.n608 585
R154 B.n610 B.n15 585
R155 B.n448 B.n73 585
R156 B.n447 B.n446 585
R157 B.n445 B.n74 585
R158 B.n444 B.n443 585
R159 B.n442 B.n75 585
R160 B.n441 B.n440 585
R161 B.n439 B.n76 585
R162 B.n438 B.n437 585
R163 B.n436 B.n77 585
R164 B.n435 B.n434 585
R165 B.n433 B.n78 585
R166 B.n432 B.n431 585
R167 B.n430 B.n79 585
R168 B.n429 B.n428 585
R169 B.n427 B.n80 585
R170 B.n426 B.n425 585
R171 B.n424 B.n81 585
R172 B.n423 B.n422 585
R173 B.n421 B.n82 585
R174 B.n420 B.n419 585
R175 B.n418 B.n83 585
R176 B.n417 B.n416 585
R177 B.n415 B.n84 585
R178 B.n414 B.n413 585
R179 B.n412 B.n85 585
R180 B.n411 B.n410 585
R181 B.n409 B.n86 585
R182 B.n408 B.n407 585
R183 B.n406 B.n87 585
R184 B.n405 B.n404 585
R185 B.n403 B.n88 585
R186 B.n402 B.n401 585
R187 B.n400 B.n89 585
R188 B.n399 B.n398 585
R189 B.n397 B.n90 585
R190 B.n396 B.n395 585
R191 B.n394 B.n91 585
R192 B.n393 B.n392 585
R193 B.n391 B.n92 585
R194 B.n390 B.n389 585
R195 B.n388 B.n93 585
R196 B.n387 B.n386 585
R197 B.n385 B.n94 585
R198 B.n384 B.n383 585
R199 B.n382 B.n95 585
R200 B.n381 B.n380 585
R201 B.n379 B.n96 585
R202 B.n378 B.n377 585
R203 B.n376 B.n97 585
R204 B.n375 B.n374 585
R205 B.n373 B.n98 585
R206 B.n372 B.n371 585
R207 B.n370 B.n99 585
R208 B.n208 B.n157 585
R209 B.n210 B.n209 585
R210 B.n211 B.n156 585
R211 B.n213 B.n212 585
R212 B.n214 B.n155 585
R213 B.n216 B.n215 585
R214 B.n217 B.n154 585
R215 B.n219 B.n218 585
R216 B.n220 B.n153 585
R217 B.n222 B.n221 585
R218 B.n223 B.n152 585
R219 B.n225 B.n224 585
R220 B.n226 B.n151 585
R221 B.n228 B.n227 585
R222 B.n229 B.n150 585
R223 B.n231 B.n230 585
R224 B.n232 B.n149 585
R225 B.n234 B.n233 585
R226 B.n235 B.n148 585
R227 B.n237 B.n236 585
R228 B.n238 B.n147 585
R229 B.n240 B.n239 585
R230 B.n241 B.n146 585
R231 B.n243 B.n242 585
R232 B.n244 B.n145 585
R233 B.n246 B.n245 585
R234 B.n247 B.n144 585
R235 B.n249 B.n248 585
R236 B.n250 B.n143 585
R237 B.n252 B.n251 585
R238 B.n253 B.n142 585
R239 B.n255 B.n254 585
R240 B.n256 B.n141 585
R241 B.n258 B.n257 585
R242 B.n259 B.n140 585
R243 B.n261 B.n260 585
R244 B.n262 B.n139 585
R245 B.n264 B.n263 585
R246 B.n265 B.n138 585
R247 B.n267 B.n266 585
R248 B.n268 B.n137 585
R249 B.n270 B.n269 585
R250 B.n271 B.n136 585
R251 B.n273 B.n272 585
R252 B.n274 B.n135 585
R253 B.n276 B.n275 585
R254 B.n277 B.n134 585
R255 B.n279 B.n278 585
R256 B.n280 B.n131 585
R257 B.n283 B.n282 585
R258 B.n284 B.n130 585
R259 B.n286 B.n285 585
R260 B.n287 B.n129 585
R261 B.n289 B.n288 585
R262 B.n290 B.n128 585
R263 B.n292 B.n291 585
R264 B.n293 B.n127 585
R265 B.n295 B.n294 585
R266 B.n297 B.n296 585
R267 B.n298 B.n123 585
R268 B.n300 B.n299 585
R269 B.n301 B.n122 585
R270 B.n303 B.n302 585
R271 B.n304 B.n121 585
R272 B.n306 B.n305 585
R273 B.n307 B.n120 585
R274 B.n309 B.n308 585
R275 B.n310 B.n119 585
R276 B.n312 B.n311 585
R277 B.n313 B.n118 585
R278 B.n315 B.n314 585
R279 B.n316 B.n117 585
R280 B.n318 B.n317 585
R281 B.n319 B.n116 585
R282 B.n321 B.n320 585
R283 B.n322 B.n115 585
R284 B.n324 B.n323 585
R285 B.n325 B.n114 585
R286 B.n327 B.n326 585
R287 B.n328 B.n113 585
R288 B.n330 B.n329 585
R289 B.n331 B.n112 585
R290 B.n333 B.n332 585
R291 B.n334 B.n111 585
R292 B.n336 B.n335 585
R293 B.n337 B.n110 585
R294 B.n339 B.n338 585
R295 B.n340 B.n109 585
R296 B.n342 B.n341 585
R297 B.n343 B.n108 585
R298 B.n345 B.n344 585
R299 B.n346 B.n107 585
R300 B.n348 B.n347 585
R301 B.n349 B.n106 585
R302 B.n351 B.n350 585
R303 B.n352 B.n105 585
R304 B.n354 B.n353 585
R305 B.n355 B.n104 585
R306 B.n357 B.n356 585
R307 B.n358 B.n103 585
R308 B.n360 B.n359 585
R309 B.n361 B.n102 585
R310 B.n363 B.n362 585
R311 B.n364 B.n101 585
R312 B.n366 B.n365 585
R313 B.n367 B.n100 585
R314 B.n369 B.n368 585
R315 B.n207 B.n206 585
R316 B.n205 B.n158 585
R317 B.n204 B.n203 585
R318 B.n202 B.n159 585
R319 B.n201 B.n200 585
R320 B.n199 B.n160 585
R321 B.n198 B.n197 585
R322 B.n196 B.n161 585
R323 B.n195 B.n194 585
R324 B.n193 B.n162 585
R325 B.n192 B.n191 585
R326 B.n190 B.n163 585
R327 B.n189 B.n188 585
R328 B.n187 B.n164 585
R329 B.n186 B.n185 585
R330 B.n184 B.n165 585
R331 B.n183 B.n182 585
R332 B.n181 B.n166 585
R333 B.n180 B.n179 585
R334 B.n178 B.n167 585
R335 B.n177 B.n176 585
R336 B.n175 B.n168 585
R337 B.n174 B.n173 585
R338 B.n172 B.n169 585
R339 B.n171 B.n170 585
R340 B.n2 B.n0 585
R341 B.n649 B.n1 585
R342 B.n648 B.n647 585
R343 B.n646 B.n3 585
R344 B.n645 B.n644 585
R345 B.n643 B.n4 585
R346 B.n642 B.n641 585
R347 B.n640 B.n5 585
R348 B.n639 B.n638 585
R349 B.n637 B.n6 585
R350 B.n636 B.n635 585
R351 B.n634 B.n7 585
R352 B.n633 B.n632 585
R353 B.n631 B.n8 585
R354 B.n630 B.n629 585
R355 B.n628 B.n9 585
R356 B.n627 B.n626 585
R357 B.n625 B.n10 585
R358 B.n624 B.n623 585
R359 B.n622 B.n11 585
R360 B.n621 B.n620 585
R361 B.n619 B.n12 585
R362 B.n618 B.n617 585
R363 B.n616 B.n13 585
R364 B.n615 B.n614 585
R365 B.n613 B.n14 585
R366 B.n612 B.n611 585
R367 B.n651 B.n650 585
R368 B.n206 B.n157 516.524
R369 B.n612 B.n15 516.524
R370 B.n368 B.n99 516.524
R371 B.n450 B.n73 516.524
R372 B.n124 B.t0 407.663
R373 B.n132 B.t9 407.663
R374 B.n40 B.t3 407.663
R375 B.n46 B.t6 407.663
R376 B.n206 B.n205 163.367
R377 B.n205 B.n204 163.367
R378 B.n204 B.n159 163.367
R379 B.n200 B.n159 163.367
R380 B.n200 B.n199 163.367
R381 B.n199 B.n198 163.367
R382 B.n198 B.n161 163.367
R383 B.n194 B.n161 163.367
R384 B.n194 B.n193 163.367
R385 B.n193 B.n192 163.367
R386 B.n192 B.n163 163.367
R387 B.n188 B.n163 163.367
R388 B.n188 B.n187 163.367
R389 B.n187 B.n186 163.367
R390 B.n186 B.n165 163.367
R391 B.n182 B.n165 163.367
R392 B.n182 B.n181 163.367
R393 B.n181 B.n180 163.367
R394 B.n180 B.n167 163.367
R395 B.n176 B.n167 163.367
R396 B.n176 B.n175 163.367
R397 B.n175 B.n174 163.367
R398 B.n174 B.n169 163.367
R399 B.n170 B.n169 163.367
R400 B.n170 B.n2 163.367
R401 B.n650 B.n2 163.367
R402 B.n650 B.n649 163.367
R403 B.n649 B.n648 163.367
R404 B.n648 B.n3 163.367
R405 B.n644 B.n3 163.367
R406 B.n644 B.n643 163.367
R407 B.n643 B.n642 163.367
R408 B.n642 B.n5 163.367
R409 B.n638 B.n5 163.367
R410 B.n638 B.n637 163.367
R411 B.n637 B.n636 163.367
R412 B.n636 B.n7 163.367
R413 B.n632 B.n7 163.367
R414 B.n632 B.n631 163.367
R415 B.n631 B.n630 163.367
R416 B.n630 B.n9 163.367
R417 B.n626 B.n9 163.367
R418 B.n626 B.n625 163.367
R419 B.n625 B.n624 163.367
R420 B.n624 B.n11 163.367
R421 B.n620 B.n11 163.367
R422 B.n620 B.n619 163.367
R423 B.n619 B.n618 163.367
R424 B.n618 B.n13 163.367
R425 B.n614 B.n13 163.367
R426 B.n614 B.n613 163.367
R427 B.n613 B.n612 163.367
R428 B.n210 B.n157 163.367
R429 B.n211 B.n210 163.367
R430 B.n212 B.n211 163.367
R431 B.n212 B.n155 163.367
R432 B.n216 B.n155 163.367
R433 B.n217 B.n216 163.367
R434 B.n218 B.n217 163.367
R435 B.n218 B.n153 163.367
R436 B.n222 B.n153 163.367
R437 B.n223 B.n222 163.367
R438 B.n224 B.n223 163.367
R439 B.n224 B.n151 163.367
R440 B.n228 B.n151 163.367
R441 B.n229 B.n228 163.367
R442 B.n230 B.n229 163.367
R443 B.n230 B.n149 163.367
R444 B.n234 B.n149 163.367
R445 B.n235 B.n234 163.367
R446 B.n236 B.n235 163.367
R447 B.n236 B.n147 163.367
R448 B.n240 B.n147 163.367
R449 B.n241 B.n240 163.367
R450 B.n242 B.n241 163.367
R451 B.n242 B.n145 163.367
R452 B.n246 B.n145 163.367
R453 B.n247 B.n246 163.367
R454 B.n248 B.n247 163.367
R455 B.n248 B.n143 163.367
R456 B.n252 B.n143 163.367
R457 B.n253 B.n252 163.367
R458 B.n254 B.n253 163.367
R459 B.n254 B.n141 163.367
R460 B.n258 B.n141 163.367
R461 B.n259 B.n258 163.367
R462 B.n260 B.n259 163.367
R463 B.n260 B.n139 163.367
R464 B.n264 B.n139 163.367
R465 B.n265 B.n264 163.367
R466 B.n266 B.n265 163.367
R467 B.n266 B.n137 163.367
R468 B.n270 B.n137 163.367
R469 B.n271 B.n270 163.367
R470 B.n272 B.n271 163.367
R471 B.n272 B.n135 163.367
R472 B.n276 B.n135 163.367
R473 B.n277 B.n276 163.367
R474 B.n278 B.n277 163.367
R475 B.n278 B.n131 163.367
R476 B.n283 B.n131 163.367
R477 B.n284 B.n283 163.367
R478 B.n285 B.n284 163.367
R479 B.n285 B.n129 163.367
R480 B.n289 B.n129 163.367
R481 B.n290 B.n289 163.367
R482 B.n291 B.n290 163.367
R483 B.n291 B.n127 163.367
R484 B.n295 B.n127 163.367
R485 B.n296 B.n295 163.367
R486 B.n296 B.n123 163.367
R487 B.n300 B.n123 163.367
R488 B.n301 B.n300 163.367
R489 B.n302 B.n301 163.367
R490 B.n302 B.n121 163.367
R491 B.n306 B.n121 163.367
R492 B.n307 B.n306 163.367
R493 B.n308 B.n307 163.367
R494 B.n308 B.n119 163.367
R495 B.n312 B.n119 163.367
R496 B.n313 B.n312 163.367
R497 B.n314 B.n313 163.367
R498 B.n314 B.n117 163.367
R499 B.n318 B.n117 163.367
R500 B.n319 B.n318 163.367
R501 B.n320 B.n319 163.367
R502 B.n320 B.n115 163.367
R503 B.n324 B.n115 163.367
R504 B.n325 B.n324 163.367
R505 B.n326 B.n325 163.367
R506 B.n326 B.n113 163.367
R507 B.n330 B.n113 163.367
R508 B.n331 B.n330 163.367
R509 B.n332 B.n331 163.367
R510 B.n332 B.n111 163.367
R511 B.n336 B.n111 163.367
R512 B.n337 B.n336 163.367
R513 B.n338 B.n337 163.367
R514 B.n338 B.n109 163.367
R515 B.n342 B.n109 163.367
R516 B.n343 B.n342 163.367
R517 B.n344 B.n343 163.367
R518 B.n344 B.n107 163.367
R519 B.n348 B.n107 163.367
R520 B.n349 B.n348 163.367
R521 B.n350 B.n349 163.367
R522 B.n350 B.n105 163.367
R523 B.n354 B.n105 163.367
R524 B.n355 B.n354 163.367
R525 B.n356 B.n355 163.367
R526 B.n356 B.n103 163.367
R527 B.n360 B.n103 163.367
R528 B.n361 B.n360 163.367
R529 B.n362 B.n361 163.367
R530 B.n362 B.n101 163.367
R531 B.n366 B.n101 163.367
R532 B.n367 B.n366 163.367
R533 B.n368 B.n367 163.367
R534 B.n372 B.n99 163.367
R535 B.n373 B.n372 163.367
R536 B.n374 B.n373 163.367
R537 B.n374 B.n97 163.367
R538 B.n378 B.n97 163.367
R539 B.n379 B.n378 163.367
R540 B.n380 B.n379 163.367
R541 B.n380 B.n95 163.367
R542 B.n384 B.n95 163.367
R543 B.n385 B.n384 163.367
R544 B.n386 B.n385 163.367
R545 B.n386 B.n93 163.367
R546 B.n390 B.n93 163.367
R547 B.n391 B.n390 163.367
R548 B.n392 B.n391 163.367
R549 B.n392 B.n91 163.367
R550 B.n396 B.n91 163.367
R551 B.n397 B.n396 163.367
R552 B.n398 B.n397 163.367
R553 B.n398 B.n89 163.367
R554 B.n402 B.n89 163.367
R555 B.n403 B.n402 163.367
R556 B.n404 B.n403 163.367
R557 B.n404 B.n87 163.367
R558 B.n408 B.n87 163.367
R559 B.n409 B.n408 163.367
R560 B.n410 B.n409 163.367
R561 B.n410 B.n85 163.367
R562 B.n414 B.n85 163.367
R563 B.n415 B.n414 163.367
R564 B.n416 B.n415 163.367
R565 B.n416 B.n83 163.367
R566 B.n420 B.n83 163.367
R567 B.n421 B.n420 163.367
R568 B.n422 B.n421 163.367
R569 B.n422 B.n81 163.367
R570 B.n426 B.n81 163.367
R571 B.n427 B.n426 163.367
R572 B.n428 B.n427 163.367
R573 B.n428 B.n79 163.367
R574 B.n432 B.n79 163.367
R575 B.n433 B.n432 163.367
R576 B.n434 B.n433 163.367
R577 B.n434 B.n77 163.367
R578 B.n438 B.n77 163.367
R579 B.n439 B.n438 163.367
R580 B.n440 B.n439 163.367
R581 B.n440 B.n75 163.367
R582 B.n444 B.n75 163.367
R583 B.n445 B.n444 163.367
R584 B.n446 B.n445 163.367
R585 B.n446 B.n73 163.367
R586 B.n608 B.n15 163.367
R587 B.n608 B.n607 163.367
R588 B.n607 B.n606 163.367
R589 B.n606 B.n17 163.367
R590 B.n602 B.n17 163.367
R591 B.n602 B.n601 163.367
R592 B.n601 B.n600 163.367
R593 B.n600 B.n19 163.367
R594 B.n596 B.n19 163.367
R595 B.n596 B.n595 163.367
R596 B.n595 B.n594 163.367
R597 B.n594 B.n21 163.367
R598 B.n590 B.n21 163.367
R599 B.n590 B.n589 163.367
R600 B.n589 B.n588 163.367
R601 B.n588 B.n23 163.367
R602 B.n584 B.n23 163.367
R603 B.n584 B.n583 163.367
R604 B.n583 B.n582 163.367
R605 B.n582 B.n25 163.367
R606 B.n578 B.n25 163.367
R607 B.n578 B.n577 163.367
R608 B.n577 B.n576 163.367
R609 B.n576 B.n27 163.367
R610 B.n572 B.n27 163.367
R611 B.n572 B.n571 163.367
R612 B.n571 B.n570 163.367
R613 B.n570 B.n29 163.367
R614 B.n566 B.n29 163.367
R615 B.n566 B.n565 163.367
R616 B.n565 B.n564 163.367
R617 B.n564 B.n31 163.367
R618 B.n560 B.n31 163.367
R619 B.n560 B.n559 163.367
R620 B.n559 B.n558 163.367
R621 B.n558 B.n33 163.367
R622 B.n554 B.n33 163.367
R623 B.n554 B.n553 163.367
R624 B.n553 B.n552 163.367
R625 B.n552 B.n35 163.367
R626 B.n548 B.n35 163.367
R627 B.n548 B.n547 163.367
R628 B.n547 B.n546 163.367
R629 B.n546 B.n37 163.367
R630 B.n542 B.n37 163.367
R631 B.n542 B.n541 163.367
R632 B.n541 B.n540 163.367
R633 B.n540 B.n39 163.367
R634 B.n535 B.n39 163.367
R635 B.n535 B.n534 163.367
R636 B.n534 B.n533 163.367
R637 B.n533 B.n43 163.367
R638 B.n529 B.n43 163.367
R639 B.n529 B.n528 163.367
R640 B.n528 B.n527 163.367
R641 B.n527 B.n45 163.367
R642 B.n523 B.n45 163.367
R643 B.n523 B.n522 163.367
R644 B.n522 B.n49 163.367
R645 B.n518 B.n49 163.367
R646 B.n518 B.n517 163.367
R647 B.n517 B.n516 163.367
R648 B.n516 B.n51 163.367
R649 B.n512 B.n51 163.367
R650 B.n512 B.n511 163.367
R651 B.n511 B.n510 163.367
R652 B.n510 B.n53 163.367
R653 B.n506 B.n53 163.367
R654 B.n506 B.n505 163.367
R655 B.n505 B.n504 163.367
R656 B.n504 B.n55 163.367
R657 B.n500 B.n55 163.367
R658 B.n500 B.n499 163.367
R659 B.n499 B.n498 163.367
R660 B.n498 B.n57 163.367
R661 B.n494 B.n57 163.367
R662 B.n494 B.n493 163.367
R663 B.n493 B.n492 163.367
R664 B.n492 B.n59 163.367
R665 B.n488 B.n59 163.367
R666 B.n488 B.n487 163.367
R667 B.n487 B.n486 163.367
R668 B.n486 B.n61 163.367
R669 B.n482 B.n61 163.367
R670 B.n482 B.n481 163.367
R671 B.n481 B.n480 163.367
R672 B.n480 B.n63 163.367
R673 B.n476 B.n63 163.367
R674 B.n476 B.n475 163.367
R675 B.n475 B.n474 163.367
R676 B.n474 B.n65 163.367
R677 B.n470 B.n65 163.367
R678 B.n470 B.n469 163.367
R679 B.n469 B.n468 163.367
R680 B.n468 B.n67 163.367
R681 B.n464 B.n67 163.367
R682 B.n464 B.n463 163.367
R683 B.n463 B.n462 163.367
R684 B.n462 B.n69 163.367
R685 B.n458 B.n69 163.367
R686 B.n458 B.n457 163.367
R687 B.n457 B.n456 163.367
R688 B.n456 B.n71 163.367
R689 B.n452 B.n71 163.367
R690 B.n452 B.n451 163.367
R691 B.n451 B.n450 163.367
R692 B.n124 B.t2 148.351
R693 B.n46 B.t7 148.351
R694 B.n132 B.t11 148.333
R695 B.n40 B.t4 148.333
R696 B.n125 B.t1 108.594
R697 B.n47 B.t8 108.594
R698 B.n133 B.t10 108.576
R699 B.n41 B.t5 108.576
R700 B.n126 B.n125 59.5399
R701 B.n281 B.n133 59.5399
R702 B.n537 B.n41 59.5399
R703 B.n48 B.n47 59.5399
R704 B.n125 B.n124 39.7581
R705 B.n133 B.n132 39.7581
R706 B.n41 B.n40 39.7581
R707 B.n47 B.n46 39.7581
R708 B.n611 B.n610 33.5615
R709 B.n449 B.n448 33.5615
R710 B.n370 B.n369 33.5615
R711 B.n208 B.n207 33.5615
R712 B B.n651 18.0485
R713 B.n610 B.n609 10.6151
R714 B.n609 B.n16 10.6151
R715 B.n605 B.n16 10.6151
R716 B.n605 B.n604 10.6151
R717 B.n604 B.n603 10.6151
R718 B.n603 B.n18 10.6151
R719 B.n599 B.n18 10.6151
R720 B.n599 B.n598 10.6151
R721 B.n598 B.n597 10.6151
R722 B.n597 B.n20 10.6151
R723 B.n593 B.n20 10.6151
R724 B.n593 B.n592 10.6151
R725 B.n592 B.n591 10.6151
R726 B.n591 B.n22 10.6151
R727 B.n587 B.n22 10.6151
R728 B.n587 B.n586 10.6151
R729 B.n586 B.n585 10.6151
R730 B.n585 B.n24 10.6151
R731 B.n581 B.n24 10.6151
R732 B.n581 B.n580 10.6151
R733 B.n580 B.n579 10.6151
R734 B.n579 B.n26 10.6151
R735 B.n575 B.n26 10.6151
R736 B.n575 B.n574 10.6151
R737 B.n574 B.n573 10.6151
R738 B.n573 B.n28 10.6151
R739 B.n569 B.n28 10.6151
R740 B.n569 B.n568 10.6151
R741 B.n568 B.n567 10.6151
R742 B.n567 B.n30 10.6151
R743 B.n563 B.n30 10.6151
R744 B.n563 B.n562 10.6151
R745 B.n562 B.n561 10.6151
R746 B.n561 B.n32 10.6151
R747 B.n557 B.n32 10.6151
R748 B.n557 B.n556 10.6151
R749 B.n556 B.n555 10.6151
R750 B.n555 B.n34 10.6151
R751 B.n551 B.n34 10.6151
R752 B.n551 B.n550 10.6151
R753 B.n550 B.n549 10.6151
R754 B.n549 B.n36 10.6151
R755 B.n545 B.n36 10.6151
R756 B.n545 B.n544 10.6151
R757 B.n544 B.n543 10.6151
R758 B.n543 B.n38 10.6151
R759 B.n539 B.n38 10.6151
R760 B.n539 B.n538 10.6151
R761 B.n536 B.n42 10.6151
R762 B.n532 B.n42 10.6151
R763 B.n532 B.n531 10.6151
R764 B.n531 B.n530 10.6151
R765 B.n530 B.n44 10.6151
R766 B.n526 B.n44 10.6151
R767 B.n526 B.n525 10.6151
R768 B.n525 B.n524 10.6151
R769 B.n521 B.n520 10.6151
R770 B.n520 B.n519 10.6151
R771 B.n519 B.n50 10.6151
R772 B.n515 B.n50 10.6151
R773 B.n515 B.n514 10.6151
R774 B.n514 B.n513 10.6151
R775 B.n513 B.n52 10.6151
R776 B.n509 B.n52 10.6151
R777 B.n509 B.n508 10.6151
R778 B.n508 B.n507 10.6151
R779 B.n507 B.n54 10.6151
R780 B.n503 B.n54 10.6151
R781 B.n503 B.n502 10.6151
R782 B.n502 B.n501 10.6151
R783 B.n501 B.n56 10.6151
R784 B.n497 B.n56 10.6151
R785 B.n497 B.n496 10.6151
R786 B.n496 B.n495 10.6151
R787 B.n495 B.n58 10.6151
R788 B.n491 B.n58 10.6151
R789 B.n491 B.n490 10.6151
R790 B.n490 B.n489 10.6151
R791 B.n489 B.n60 10.6151
R792 B.n485 B.n60 10.6151
R793 B.n485 B.n484 10.6151
R794 B.n484 B.n483 10.6151
R795 B.n483 B.n62 10.6151
R796 B.n479 B.n62 10.6151
R797 B.n479 B.n478 10.6151
R798 B.n478 B.n477 10.6151
R799 B.n477 B.n64 10.6151
R800 B.n473 B.n64 10.6151
R801 B.n473 B.n472 10.6151
R802 B.n472 B.n471 10.6151
R803 B.n471 B.n66 10.6151
R804 B.n467 B.n66 10.6151
R805 B.n467 B.n466 10.6151
R806 B.n466 B.n465 10.6151
R807 B.n465 B.n68 10.6151
R808 B.n461 B.n68 10.6151
R809 B.n461 B.n460 10.6151
R810 B.n460 B.n459 10.6151
R811 B.n459 B.n70 10.6151
R812 B.n455 B.n70 10.6151
R813 B.n455 B.n454 10.6151
R814 B.n454 B.n453 10.6151
R815 B.n453 B.n72 10.6151
R816 B.n449 B.n72 10.6151
R817 B.n371 B.n370 10.6151
R818 B.n371 B.n98 10.6151
R819 B.n375 B.n98 10.6151
R820 B.n376 B.n375 10.6151
R821 B.n377 B.n376 10.6151
R822 B.n377 B.n96 10.6151
R823 B.n381 B.n96 10.6151
R824 B.n382 B.n381 10.6151
R825 B.n383 B.n382 10.6151
R826 B.n383 B.n94 10.6151
R827 B.n387 B.n94 10.6151
R828 B.n388 B.n387 10.6151
R829 B.n389 B.n388 10.6151
R830 B.n389 B.n92 10.6151
R831 B.n393 B.n92 10.6151
R832 B.n394 B.n393 10.6151
R833 B.n395 B.n394 10.6151
R834 B.n395 B.n90 10.6151
R835 B.n399 B.n90 10.6151
R836 B.n400 B.n399 10.6151
R837 B.n401 B.n400 10.6151
R838 B.n401 B.n88 10.6151
R839 B.n405 B.n88 10.6151
R840 B.n406 B.n405 10.6151
R841 B.n407 B.n406 10.6151
R842 B.n407 B.n86 10.6151
R843 B.n411 B.n86 10.6151
R844 B.n412 B.n411 10.6151
R845 B.n413 B.n412 10.6151
R846 B.n413 B.n84 10.6151
R847 B.n417 B.n84 10.6151
R848 B.n418 B.n417 10.6151
R849 B.n419 B.n418 10.6151
R850 B.n419 B.n82 10.6151
R851 B.n423 B.n82 10.6151
R852 B.n424 B.n423 10.6151
R853 B.n425 B.n424 10.6151
R854 B.n425 B.n80 10.6151
R855 B.n429 B.n80 10.6151
R856 B.n430 B.n429 10.6151
R857 B.n431 B.n430 10.6151
R858 B.n431 B.n78 10.6151
R859 B.n435 B.n78 10.6151
R860 B.n436 B.n435 10.6151
R861 B.n437 B.n436 10.6151
R862 B.n437 B.n76 10.6151
R863 B.n441 B.n76 10.6151
R864 B.n442 B.n441 10.6151
R865 B.n443 B.n442 10.6151
R866 B.n443 B.n74 10.6151
R867 B.n447 B.n74 10.6151
R868 B.n448 B.n447 10.6151
R869 B.n209 B.n208 10.6151
R870 B.n209 B.n156 10.6151
R871 B.n213 B.n156 10.6151
R872 B.n214 B.n213 10.6151
R873 B.n215 B.n214 10.6151
R874 B.n215 B.n154 10.6151
R875 B.n219 B.n154 10.6151
R876 B.n220 B.n219 10.6151
R877 B.n221 B.n220 10.6151
R878 B.n221 B.n152 10.6151
R879 B.n225 B.n152 10.6151
R880 B.n226 B.n225 10.6151
R881 B.n227 B.n226 10.6151
R882 B.n227 B.n150 10.6151
R883 B.n231 B.n150 10.6151
R884 B.n232 B.n231 10.6151
R885 B.n233 B.n232 10.6151
R886 B.n233 B.n148 10.6151
R887 B.n237 B.n148 10.6151
R888 B.n238 B.n237 10.6151
R889 B.n239 B.n238 10.6151
R890 B.n239 B.n146 10.6151
R891 B.n243 B.n146 10.6151
R892 B.n244 B.n243 10.6151
R893 B.n245 B.n244 10.6151
R894 B.n245 B.n144 10.6151
R895 B.n249 B.n144 10.6151
R896 B.n250 B.n249 10.6151
R897 B.n251 B.n250 10.6151
R898 B.n251 B.n142 10.6151
R899 B.n255 B.n142 10.6151
R900 B.n256 B.n255 10.6151
R901 B.n257 B.n256 10.6151
R902 B.n257 B.n140 10.6151
R903 B.n261 B.n140 10.6151
R904 B.n262 B.n261 10.6151
R905 B.n263 B.n262 10.6151
R906 B.n263 B.n138 10.6151
R907 B.n267 B.n138 10.6151
R908 B.n268 B.n267 10.6151
R909 B.n269 B.n268 10.6151
R910 B.n269 B.n136 10.6151
R911 B.n273 B.n136 10.6151
R912 B.n274 B.n273 10.6151
R913 B.n275 B.n274 10.6151
R914 B.n275 B.n134 10.6151
R915 B.n279 B.n134 10.6151
R916 B.n280 B.n279 10.6151
R917 B.n282 B.n130 10.6151
R918 B.n286 B.n130 10.6151
R919 B.n287 B.n286 10.6151
R920 B.n288 B.n287 10.6151
R921 B.n288 B.n128 10.6151
R922 B.n292 B.n128 10.6151
R923 B.n293 B.n292 10.6151
R924 B.n294 B.n293 10.6151
R925 B.n298 B.n297 10.6151
R926 B.n299 B.n298 10.6151
R927 B.n299 B.n122 10.6151
R928 B.n303 B.n122 10.6151
R929 B.n304 B.n303 10.6151
R930 B.n305 B.n304 10.6151
R931 B.n305 B.n120 10.6151
R932 B.n309 B.n120 10.6151
R933 B.n310 B.n309 10.6151
R934 B.n311 B.n310 10.6151
R935 B.n311 B.n118 10.6151
R936 B.n315 B.n118 10.6151
R937 B.n316 B.n315 10.6151
R938 B.n317 B.n316 10.6151
R939 B.n317 B.n116 10.6151
R940 B.n321 B.n116 10.6151
R941 B.n322 B.n321 10.6151
R942 B.n323 B.n322 10.6151
R943 B.n323 B.n114 10.6151
R944 B.n327 B.n114 10.6151
R945 B.n328 B.n327 10.6151
R946 B.n329 B.n328 10.6151
R947 B.n329 B.n112 10.6151
R948 B.n333 B.n112 10.6151
R949 B.n334 B.n333 10.6151
R950 B.n335 B.n334 10.6151
R951 B.n335 B.n110 10.6151
R952 B.n339 B.n110 10.6151
R953 B.n340 B.n339 10.6151
R954 B.n341 B.n340 10.6151
R955 B.n341 B.n108 10.6151
R956 B.n345 B.n108 10.6151
R957 B.n346 B.n345 10.6151
R958 B.n347 B.n346 10.6151
R959 B.n347 B.n106 10.6151
R960 B.n351 B.n106 10.6151
R961 B.n352 B.n351 10.6151
R962 B.n353 B.n352 10.6151
R963 B.n353 B.n104 10.6151
R964 B.n357 B.n104 10.6151
R965 B.n358 B.n357 10.6151
R966 B.n359 B.n358 10.6151
R967 B.n359 B.n102 10.6151
R968 B.n363 B.n102 10.6151
R969 B.n364 B.n363 10.6151
R970 B.n365 B.n364 10.6151
R971 B.n365 B.n100 10.6151
R972 B.n369 B.n100 10.6151
R973 B.n207 B.n158 10.6151
R974 B.n203 B.n158 10.6151
R975 B.n203 B.n202 10.6151
R976 B.n202 B.n201 10.6151
R977 B.n201 B.n160 10.6151
R978 B.n197 B.n160 10.6151
R979 B.n197 B.n196 10.6151
R980 B.n196 B.n195 10.6151
R981 B.n195 B.n162 10.6151
R982 B.n191 B.n162 10.6151
R983 B.n191 B.n190 10.6151
R984 B.n190 B.n189 10.6151
R985 B.n189 B.n164 10.6151
R986 B.n185 B.n164 10.6151
R987 B.n185 B.n184 10.6151
R988 B.n184 B.n183 10.6151
R989 B.n183 B.n166 10.6151
R990 B.n179 B.n166 10.6151
R991 B.n179 B.n178 10.6151
R992 B.n178 B.n177 10.6151
R993 B.n177 B.n168 10.6151
R994 B.n173 B.n168 10.6151
R995 B.n173 B.n172 10.6151
R996 B.n172 B.n171 10.6151
R997 B.n171 B.n0 10.6151
R998 B.n647 B.n1 10.6151
R999 B.n647 B.n646 10.6151
R1000 B.n646 B.n645 10.6151
R1001 B.n645 B.n4 10.6151
R1002 B.n641 B.n4 10.6151
R1003 B.n641 B.n640 10.6151
R1004 B.n640 B.n639 10.6151
R1005 B.n639 B.n6 10.6151
R1006 B.n635 B.n6 10.6151
R1007 B.n635 B.n634 10.6151
R1008 B.n634 B.n633 10.6151
R1009 B.n633 B.n8 10.6151
R1010 B.n629 B.n8 10.6151
R1011 B.n629 B.n628 10.6151
R1012 B.n628 B.n627 10.6151
R1013 B.n627 B.n10 10.6151
R1014 B.n623 B.n10 10.6151
R1015 B.n623 B.n622 10.6151
R1016 B.n622 B.n621 10.6151
R1017 B.n621 B.n12 10.6151
R1018 B.n617 B.n12 10.6151
R1019 B.n617 B.n616 10.6151
R1020 B.n616 B.n615 10.6151
R1021 B.n615 B.n14 10.6151
R1022 B.n611 B.n14 10.6151
R1023 B.n537 B.n536 6.5566
R1024 B.n524 B.n48 6.5566
R1025 B.n282 B.n281 6.5566
R1026 B.n294 B.n126 6.5566
R1027 B.n538 B.n537 4.05904
R1028 B.n521 B.n48 4.05904
R1029 B.n281 B.n280 4.05904
R1030 B.n297 B.n126 4.05904
R1031 B.n651 B.n0 2.81026
R1032 B.n651 B.n1 2.81026
R1033 VN.n0 VN.t0 236.756
R1034 VN.n1 VN.t1 236.756
R1035 VN.n0 VN.t2 236.333
R1036 VN.n1 VN.t3 236.333
R1037 VN VN.n1 55.181
R1038 VN VN.n0 9.5333
R1039 VDD2.n2 VDD2.n0 114.394
R1040 VDD2.n2 VDD2.n1 72.9818
R1041 VDD2.n1 VDD2.t0 2.26093
R1042 VDD2.n1 VDD2.t2 2.26093
R1043 VDD2.n0 VDD2.t3 2.26093
R1044 VDD2.n0 VDD2.t1 2.26093
R1045 VDD2 VDD2.n2 0.0586897
C0 B w_n2200_n3844# 8.82995f
C1 VTAIL w_n2200_n3844# 4.53388f
C2 VDD1 VDD2 0.811921f
C3 VN w_n2200_n3844# 3.61954f
C4 VP w_n2200_n3844# 3.90013f
C5 w_n2200_n3844# VDD1 1.34135f
C6 B VTAIL 5.23516f
C7 B VN 0.966661f
C8 VP B 1.4282f
C9 VN VTAIL 4.83442f
C10 VP VTAIL 4.84852f
C11 VP VN 6.00299f
C12 B VDD1 1.17127f
C13 w_n2200_n3844# VDD2 1.37778f
C14 VTAIL VDD1 6.11122f
C15 VN VDD1 0.147691f
C16 VP VDD1 5.33916f
C17 B VDD2 1.20904f
C18 VTAIL VDD2 6.15952f
C19 VN VDD2 5.14957f
C20 VP VDD2 0.337796f
C21 VDD2 VSUBS 0.86698f
C22 VDD1 VSUBS 5.54735f
C23 VTAIL VSUBS 1.191577f
C24 VN VSUBS 5.25066f
C25 VP VSUBS 1.893234f
C26 B VSUBS 3.715142f
C27 w_n2200_n3844# VSUBS 0.103778p
C28 VDD2.t3 VSUBS 0.302269f
C29 VDD2.t1 VSUBS 0.302269f
C30 VDD2.n0 VSUBS 3.18314f
C31 VDD2.t0 VSUBS 0.302269f
C32 VDD2.t2 VSUBS 0.302269f
C33 VDD2.n1 VSUBS 2.44545f
C34 VDD2.n2 VSUBS 4.30514f
C35 VN.t0 VSUBS 2.81996f
C36 VN.t2 VSUBS 2.81793f
C37 VN.n0 VSUBS 1.98415f
C38 VN.t1 VSUBS 2.81996f
C39 VN.t3 VSUBS 2.81793f
C40 VN.n1 VSUBS 3.73177f
C41 B.n0 VSUBS 0.004402f
C42 B.n1 VSUBS 0.004402f
C43 B.n2 VSUBS 0.006961f
C44 B.n3 VSUBS 0.006961f
C45 B.n4 VSUBS 0.006961f
C46 B.n5 VSUBS 0.006961f
C47 B.n6 VSUBS 0.006961f
C48 B.n7 VSUBS 0.006961f
C49 B.n8 VSUBS 0.006961f
C50 B.n9 VSUBS 0.006961f
C51 B.n10 VSUBS 0.006961f
C52 B.n11 VSUBS 0.006961f
C53 B.n12 VSUBS 0.006961f
C54 B.n13 VSUBS 0.006961f
C55 B.n14 VSUBS 0.006961f
C56 B.n15 VSUBS 0.01716f
C57 B.n16 VSUBS 0.006961f
C58 B.n17 VSUBS 0.006961f
C59 B.n18 VSUBS 0.006961f
C60 B.n19 VSUBS 0.006961f
C61 B.n20 VSUBS 0.006961f
C62 B.n21 VSUBS 0.006961f
C63 B.n22 VSUBS 0.006961f
C64 B.n23 VSUBS 0.006961f
C65 B.n24 VSUBS 0.006961f
C66 B.n25 VSUBS 0.006961f
C67 B.n26 VSUBS 0.006961f
C68 B.n27 VSUBS 0.006961f
C69 B.n28 VSUBS 0.006961f
C70 B.n29 VSUBS 0.006961f
C71 B.n30 VSUBS 0.006961f
C72 B.n31 VSUBS 0.006961f
C73 B.n32 VSUBS 0.006961f
C74 B.n33 VSUBS 0.006961f
C75 B.n34 VSUBS 0.006961f
C76 B.n35 VSUBS 0.006961f
C77 B.n36 VSUBS 0.006961f
C78 B.n37 VSUBS 0.006961f
C79 B.n38 VSUBS 0.006961f
C80 B.n39 VSUBS 0.006961f
C81 B.t5 VSUBS 0.474303f
C82 B.t4 VSUBS 0.489849f
C83 B.t3 VSUBS 1.07372f
C84 B.n40 VSUBS 0.226162f
C85 B.n41 VSUBS 0.067929f
C86 B.n42 VSUBS 0.006961f
C87 B.n43 VSUBS 0.006961f
C88 B.n44 VSUBS 0.006961f
C89 B.n45 VSUBS 0.006961f
C90 B.t8 VSUBS 0.474291f
C91 B.t7 VSUBS 0.489838f
C92 B.t6 VSUBS 1.07372f
C93 B.n46 VSUBS 0.226173f
C94 B.n47 VSUBS 0.067941f
C95 B.n48 VSUBS 0.016128f
C96 B.n49 VSUBS 0.006961f
C97 B.n50 VSUBS 0.006961f
C98 B.n51 VSUBS 0.006961f
C99 B.n52 VSUBS 0.006961f
C100 B.n53 VSUBS 0.006961f
C101 B.n54 VSUBS 0.006961f
C102 B.n55 VSUBS 0.006961f
C103 B.n56 VSUBS 0.006961f
C104 B.n57 VSUBS 0.006961f
C105 B.n58 VSUBS 0.006961f
C106 B.n59 VSUBS 0.006961f
C107 B.n60 VSUBS 0.006961f
C108 B.n61 VSUBS 0.006961f
C109 B.n62 VSUBS 0.006961f
C110 B.n63 VSUBS 0.006961f
C111 B.n64 VSUBS 0.006961f
C112 B.n65 VSUBS 0.006961f
C113 B.n66 VSUBS 0.006961f
C114 B.n67 VSUBS 0.006961f
C115 B.n68 VSUBS 0.006961f
C116 B.n69 VSUBS 0.006961f
C117 B.n70 VSUBS 0.006961f
C118 B.n71 VSUBS 0.006961f
C119 B.n72 VSUBS 0.006961f
C120 B.n73 VSUBS 0.016008f
C121 B.n74 VSUBS 0.006961f
C122 B.n75 VSUBS 0.006961f
C123 B.n76 VSUBS 0.006961f
C124 B.n77 VSUBS 0.006961f
C125 B.n78 VSUBS 0.006961f
C126 B.n79 VSUBS 0.006961f
C127 B.n80 VSUBS 0.006961f
C128 B.n81 VSUBS 0.006961f
C129 B.n82 VSUBS 0.006961f
C130 B.n83 VSUBS 0.006961f
C131 B.n84 VSUBS 0.006961f
C132 B.n85 VSUBS 0.006961f
C133 B.n86 VSUBS 0.006961f
C134 B.n87 VSUBS 0.006961f
C135 B.n88 VSUBS 0.006961f
C136 B.n89 VSUBS 0.006961f
C137 B.n90 VSUBS 0.006961f
C138 B.n91 VSUBS 0.006961f
C139 B.n92 VSUBS 0.006961f
C140 B.n93 VSUBS 0.006961f
C141 B.n94 VSUBS 0.006961f
C142 B.n95 VSUBS 0.006961f
C143 B.n96 VSUBS 0.006961f
C144 B.n97 VSUBS 0.006961f
C145 B.n98 VSUBS 0.006961f
C146 B.n99 VSUBS 0.016008f
C147 B.n100 VSUBS 0.006961f
C148 B.n101 VSUBS 0.006961f
C149 B.n102 VSUBS 0.006961f
C150 B.n103 VSUBS 0.006961f
C151 B.n104 VSUBS 0.006961f
C152 B.n105 VSUBS 0.006961f
C153 B.n106 VSUBS 0.006961f
C154 B.n107 VSUBS 0.006961f
C155 B.n108 VSUBS 0.006961f
C156 B.n109 VSUBS 0.006961f
C157 B.n110 VSUBS 0.006961f
C158 B.n111 VSUBS 0.006961f
C159 B.n112 VSUBS 0.006961f
C160 B.n113 VSUBS 0.006961f
C161 B.n114 VSUBS 0.006961f
C162 B.n115 VSUBS 0.006961f
C163 B.n116 VSUBS 0.006961f
C164 B.n117 VSUBS 0.006961f
C165 B.n118 VSUBS 0.006961f
C166 B.n119 VSUBS 0.006961f
C167 B.n120 VSUBS 0.006961f
C168 B.n121 VSUBS 0.006961f
C169 B.n122 VSUBS 0.006961f
C170 B.n123 VSUBS 0.006961f
C171 B.t1 VSUBS 0.474291f
C172 B.t2 VSUBS 0.489838f
C173 B.t0 VSUBS 1.07372f
C174 B.n124 VSUBS 0.226173f
C175 B.n125 VSUBS 0.067941f
C176 B.n126 VSUBS 0.016128f
C177 B.n127 VSUBS 0.006961f
C178 B.n128 VSUBS 0.006961f
C179 B.n129 VSUBS 0.006961f
C180 B.n130 VSUBS 0.006961f
C181 B.n131 VSUBS 0.006961f
C182 B.t10 VSUBS 0.474303f
C183 B.t11 VSUBS 0.489849f
C184 B.t9 VSUBS 1.07372f
C185 B.n132 VSUBS 0.226162f
C186 B.n133 VSUBS 0.067929f
C187 B.n134 VSUBS 0.006961f
C188 B.n135 VSUBS 0.006961f
C189 B.n136 VSUBS 0.006961f
C190 B.n137 VSUBS 0.006961f
C191 B.n138 VSUBS 0.006961f
C192 B.n139 VSUBS 0.006961f
C193 B.n140 VSUBS 0.006961f
C194 B.n141 VSUBS 0.006961f
C195 B.n142 VSUBS 0.006961f
C196 B.n143 VSUBS 0.006961f
C197 B.n144 VSUBS 0.006961f
C198 B.n145 VSUBS 0.006961f
C199 B.n146 VSUBS 0.006961f
C200 B.n147 VSUBS 0.006961f
C201 B.n148 VSUBS 0.006961f
C202 B.n149 VSUBS 0.006961f
C203 B.n150 VSUBS 0.006961f
C204 B.n151 VSUBS 0.006961f
C205 B.n152 VSUBS 0.006961f
C206 B.n153 VSUBS 0.006961f
C207 B.n154 VSUBS 0.006961f
C208 B.n155 VSUBS 0.006961f
C209 B.n156 VSUBS 0.006961f
C210 B.n157 VSUBS 0.01716f
C211 B.n158 VSUBS 0.006961f
C212 B.n159 VSUBS 0.006961f
C213 B.n160 VSUBS 0.006961f
C214 B.n161 VSUBS 0.006961f
C215 B.n162 VSUBS 0.006961f
C216 B.n163 VSUBS 0.006961f
C217 B.n164 VSUBS 0.006961f
C218 B.n165 VSUBS 0.006961f
C219 B.n166 VSUBS 0.006961f
C220 B.n167 VSUBS 0.006961f
C221 B.n168 VSUBS 0.006961f
C222 B.n169 VSUBS 0.006961f
C223 B.n170 VSUBS 0.006961f
C224 B.n171 VSUBS 0.006961f
C225 B.n172 VSUBS 0.006961f
C226 B.n173 VSUBS 0.006961f
C227 B.n174 VSUBS 0.006961f
C228 B.n175 VSUBS 0.006961f
C229 B.n176 VSUBS 0.006961f
C230 B.n177 VSUBS 0.006961f
C231 B.n178 VSUBS 0.006961f
C232 B.n179 VSUBS 0.006961f
C233 B.n180 VSUBS 0.006961f
C234 B.n181 VSUBS 0.006961f
C235 B.n182 VSUBS 0.006961f
C236 B.n183 VSUBS 0.006961f
C237 B.n184 VSUBS 0.006961f
C238 B.n185 VSUBS 0.006961f
C239 B.n186 VSUBS 0.006961f
C240 B.n187 VSUBS 0.006961f
C241 B.n188 VSUBS 0.006961f
C242 B.n189 VSUBS 0.006961f
C243 B.n190 VSUBS 0.006961f
C244 B.n191 VSUBS 0.006961f
C245 B.n192 VSUBS 0.006961f
C246 B.n193 VSUBS 0.006961f
C247 B.n194 VSUBS 0.006961f
C248 B.n195 VSUBS 0.006961f
C249 B.n196 VSUBS 0.006961f
C250 B.n197 VSUBS 0.006961f
C251 B.n198 VSUBS 0.006961f
C252 B.n199 VSUBS 0.006961f
C253 B.n200 VSUBS 0.006961f
C254 B.n201 VSUBS 0.006961f
C255 B.n202 VSUBS 0.006961f
C256 B.n203 VSUBS 0.006961f
C257 B.n204 VSUBS 0.006961f
C258 B.n205 VSUBS 0.006961f
C259 B.n206 VSUBS 0.016008f
C260 B.n207 VSUBS 0.016008f
C261 B.n208 VSUBS 0.01716f
C262 B.n209 VSUBS 0.006961f
C263 B.n210 VSUBS 0.006961f
C264 B.n211 VSUBS 0.006961f
C265 B.n212 VSUBS 0.006961f
C266 B.n213 VSUBS 0.006961f
C267 B.n214 VSUBS 0.006961f
C268 B.n215 VSUBS 0.006961f
C269 B.n216 VSUBS 0.006961f
C270 B.n217 VSUBS 0.006961f
C271 B.n218 VSUBS 0.006961f
C272 B.n219 VSUBS 0.006961f
C273 B.n220 VSUBS 0.006961f
C274 B.n221 VSUBS 0.006961f
C275 B.n222 VSUBS 0.006961f
C276 B.n223 VSUBS 0.006961f
C277 B.n224 VSUBS 0.006961f
C278 B.n225 VSUBS 0.006961f
C279 B.n226 VSUBS 0.006961f
C280 B.n227 VSUBS 0.006961f
C281 B.n228 VSUBS 0.006961f
C282 B.n229 VSUBS 0.006961f
C283 B.n230 VSUBS 0.006961f
C284 B.n231 VSUBS 0.006961f
C285 B.n232 VSUBS 0.006961f
C286 B.n233 VSUBS 0.006961f
C287 B.n234 VSUBS 0.006961f
C288 B.n235 VSUBS 0.006961f
C289 B.n236 VSUBS 0.006961f
C290 B.n237 VSUBS 0.006961f
C291 B.n238 VSUBS 0.006961f
C292 B.n239 VSUBS 0.006961f
C293 B.n240 VSUBS 0.006961f
C294 B.n241 VSUBS 0.006961f
C295 B.n242 VSUBS 0.006961f
C296 B.n243 VSUBS 0.006961f
C297 B.n244 VSUBS 0.006961f
C298 B.n245 VSUBS 0.006961f
C299 B.n246 VSUBS 0.006961f
C300 B.n247 VSUBS 0.006961f
C301 B.n248 VSUBS 0.006961f
C302 B.n249 VSUBS 0.006961f
C303 B.n250 VSUBS 0.006961f
C304 B.n251 VSUBS 0.006961f
C305 B.n252 VSUBS 0.006961f
C306 B.n253 VSUBS 0.006961f
C307 B.n254 VSUBS 0.006961f
C308 B.n255 VSUBS 0.006961f
C309 B.n256 VSUBS 0.006961f
C310 B.n257 VSUBS 0.006961f
C311 B.n258 VSUBS 0.006961f
C312 B.n259 VSUBS 0.006961f
C313 B.n260 VSUBS 0.006961f
C314 B.n261 VSUBS 0.006961f
C315 B.n262 VSUBS 0.006961f
C316 B.n263 VSUBS 0.006961f
C317 B.n264 VSUBS 0.006961f
C318 B.n265 VSUBS 0.006961f
C319 B.n266 VSUBS 0.006961f
C320 B.n267 VSUBS 0.006961f
C321 B.n268 VSUBS 0.006961f
C322 B.n269 VSUBS 0.006961f
C323 B.n270 VSUBS 0.006961f
C324 B.n271 VSUBS 0.006961f
C325 B.n272 VSUBS 0.006961f
C326 B.n273 VSUBS 0.006961f
C327 B.n274 VSUBS 0.006961f
C328 B.n275 VSUBS 0.006961f
C329 B.n276 VSUBS 0.006961f
C330 B.n277 VSUBS 0.006961f
C331 B.n278 VSUBS 0.006961f
C332 B.n279 VSUBS 0.006961f
C333 B.n280 VSUBS 0.004811f
C334 B.n281 VSUBS 0.016128f
C335 B.n282 VSUBS 0.00563f
C336 B.n283 VSUBS 0.006961f
C337 B.n284 VSUBS 0.006961f
C338 B.n285 VSUBS 0.006961f
C339 B.n286 VSUBS 0.006961f
C340 B.n287 VSUBS 0.006961f
C341 B.n288 VSUBS 0.006961f
C342 B.n289 VSUBS 0.006961f
C343 B.n290 VSUBS 0.006961f
C344 B.n291 VSUBS 0.006961f
C345 B.n292 VSUBS 0.006961f
C346 B.n293 VSUBS 0.006961f
C347 B.n294 VSUBS 0.00563f
C348 B.n295 VSUBS 0.006961f
C349 B.n296 VSUBS 0.006961f
C350 B.n297 VSUBS 0.004811f
C351 B.n298 VSUBS 0.006961f
C352 B.n299 VSUBS 0.006961f
C353 B.n300 VSUBS 0.006961f
C354 B.n301 VSUBS 0.006961f
C355 B.n302 VSUBS 0.006961f
C356 B.n303 VSUBS 0.006961f
C357 B.n304 VSUBS 0.006961f
C358 B.n305 VSUBS 0.006961f
C359 B.n306 VSUBS 0.006961f
C360 B.n307 VSUBS 0.006961f
C361 B.n308 VSUBS 0.006961f
C362 B.n309 VSUBS 0.006961f
C363 B.n310 VSUBS 0.006961f
C364 B.n311 VSUBS 0.006961f
C365 B.n312 VSUBS 0.006961f
C366 B.n313 VSUBS 0.006961f
C367 B.n314 VSUBS 0.006961f
C368 B.n315 VSUBS 0.006961f
C369 B.n316 VSUBS 0.006961f
C370 B.n317 VSUBS 0.006961f
C371 B.n318 VSUBS 0.006961f
C372 B.n319 VSUBS 0.006961f
C373 B.n320 VSUBS 0.006961f
C374 B.n321 VSUBS 0.006961f
C375 B.n322 VSUBS 0.006961f
C376 B.n323 VSUBS 0.006961f
C377 B.n324 VSUBS 0.006961f
C378 B.n325 VSUBS 0.006961f
C379 B.n326 VSUBS 0.006961f
C380 B.n327 VSUBS 0.006961f
C381 B.n328 VSUBS 0.006961f
C382 B.n329 VSUBS 0.006961f
C383 B.n330 VSUBS 0.006961f
C384 B.n331 VSUBS 0.006961f
C385 B.n332 VSUBS 0.006961f
C386 B.n333 VSUBS 0.006961f
C387 B.n334 VSUBS 0.006961f
C388 B.n335 VSUBS 0.006961f
C389 B.n336 VSUBS 0.006961f
C390 B.n337 VSUBS 0.006961f
C391 B.n338 VSUBS 0.006961f
C392 B.n339 VSUBS 0.006961f
C393 B.n340 VSUBS 0.006961f
C394 B.n341 VSUBS 0.006961f
C395 B.n342 VSUBS 0.006961f
C396 B.n343 VSUBS 0.006961f
C397 B.n344 VSUBS 0.006961f
C398 B.n345 VSUBS 0.006961f
C399 B.n346 VSUBS 0.006961f
C400 B.n347 VSUBS 0.006961f
C401 B.n348 VSUBS 0.006961f
C402 B.n349 VSUBS 0.006961f
C403 B.n350 VSUBS 0.006961f
C404 B.n351 VSUBS 0.006961f
C405 B.n352 VSUBS 0.006961f
C406 B.n353 VSUBS 0.006961f
C407 B.n354 VSUBS 0.006961f
C408 B.n355 VSUBS 0.006961f
C409 B.n356 VSUBS 0.006961f
C410 B.n357 VSUBS 0.006961f
C411 B.n358 VSUBS 0.006961f
C412 B.n359 VSUBS 0.006961f
C413 B.n360 VSUBS 0.006961f
C414 B.n361 VSUBS 0.006961f
C415 B.n362 VSUBS 0.006961f
C416 B.n363 VSUBS 0.006961f
C417 B.n364 VSUBS 0.006961f
C418 B.n365 VSUBS 0.006961f
C419 B.n366 VSUBS 0.006961f
C420 B.n367 VSUBS 0.006961f
C421 B.n368 VSUBS 0.01716f
C422 B.n369 VSUBS 0.01716f
C423 B.n370 VSUBS 0.016008f
C424 B.n371 VSUBS 0.006961f
C425 B.n372 VSUBS 0.006961f
C426 B.n373 VSUBS 0.006961f
C427 B.n374 VSUBS 0.006961f
C428 B.n375 VSUBS 0.006961f
C429 B.n376 VSUBS 0.006961f
C430 B.n377 VSUBS 0.006961f
C431 B.n378 VSUBS 0.006961f
C432 B.n379 VSUBS 0.006961f
C433 B.n380 VSUBS 0.006961f
C434 B.n381 VSUBS 0.006961f
C435 B.n382 VSUBS 0.006961f
C436 B.n383 VSUBS 0.006961f
C437 B.n384 VSUBS 0.006961f
C438 B.n385 VSUBS 0.006961f
C439 B.n386 VSUBS 0.006961f
C440 B.n387 VSUBS 0.006961f
C441 B.n388 VSUBS 0.006961f
C442 B.n389 VSUBS 0.006961f
C443 B.n390 VSUBS 0.006961f
C444 B.n391 VSUBS 0.006961f
C445 B.n392 VSUBS 0.006961f
C446 B.n393 VSUBS 0.006961f
C447 B.n394 VSUBS 0.006961f
C448 B.n395 VSUBS 0.006961f
C449 B.n396 VSUBS 0.006961f
C450 B.n397 VSUBS 0.006961f
C451 B.n398 VSUBS 0.006961f
C452 B.n399 VSUBS 0.006961f
C453 B.n400 VSUBS 0.006961f
C454 B.n401 VSUBS 0.006961f
C455 B.n402 VSUBS 0.006961f
C456 B.n403 VSUBS 0.006961f
C457 B.n404 VSUBS 0.006961f
C458 B.n405 VSUBS 0.006961f
C459 B.n406 VSUBS 0.006961f
C460 B.n407 VSUBS 0.006961f
C461 B.n408 VSUBS 0.006961f
C462 B.n409 VSUBS 0.006961f
C463 B.n410 VSUBS 0.006961f
C464 B.n411 VSUBS 0.006961f
C465 B.n412 VSUBS 0.006961f
C466 B.n413 VSUBS 0.006961f
C467 B.n414 VSUBS 0.006961f
C468 B.n415 VSUBS 0.006961f
C469 B.n416 VSUBS 0.006961f
C470 B.n417 VSUBS 0.006961f
C471 B.n418 VSUBS 0.006961f
C472 B.n419 VSUBS 0.006961f
C473 B.n420 VSUBS 0.006961f
C474 B.n421 VSUBS 0.006961f
C475 B.n422 VSUBS 0.006961f
C476 B.n423 VSUBS 0.006961f
C477 B.n424 VSUBS 0.006961f
C478 B.n425 VSUBS 0.006961f
C479 B.n426 VSUBS 0.006961f
C480 B.n427 VSUBS 0.006961f
C481 B.n428 VSUBS 0.006961f
C482 B.n429 VSUBS 0.006961f
C483 B.n430 VSUBS 0.006961f
C484 B.n431 VSUBS 0.006961f
C485 B.n432 VSUBS 0.006961f
C486 B.n433 VSUBS 0.006961f
C487 B.n434 VSUBS 0.006961f
C488 B.n435 VSUBS 0.006961f
C489 B.n436 VSUBS 0.006961f
C490 B.n437 VSUBS 0.006961f
C491 B.n438 VSUBS 0.006961f
C492 B.n439 VSUBS 0.006961f
C493 B.n440 VSUBS 0.006961f
C494 B.n441 VSUBS 0.006961f
C495 B.n442 VSUBS 0.006961f
C496 B.n443 VSUBS 0.006961f
C497 B.n444 VSUBS 0.006961f
C498 B.n445 VSUBS 0.006961f
C499 B.n446 VSUBS 0.006961f
C500 B.n447 VSUBS 0.006961f
C501 B.n448 VSUBS 0.016808f
C502 B.n449 VSUBS 0.016359f
C503 B.n450 VSUBS 0.01716f
C504 B.n451 VSUBS 0.006961f
C505 B.n452 VSUBS 0.006961f
C506 B.n453 VSUBS 0.006961f
C507 B.n454 VSUBS 0.006961f
C508 B.n455 VSUBS 0.006961f
C509 B.n456 VSUBS 0.006961f
C510 B.n457 VSUBS 0.006961f
C511 B.n458 VSUBS 0.006961f
C512 B.n459 VSUBS 0.006961f
C513 B.n460 VSUBS 0.006961f
C514 B.n461 VSUBS 0.006961f
C515 B.n462 VSUBS 0.006961f
C516 B.n463 VSUBS 0.006961f
C517 B.n464 VSUBS 0.006961f
C518 B.n465 VSUBS 0.006961f
C519 B.n466 VSUBS 0.006961f
C520 B.n467 VSUBS 0.006961f
C521 B.n468 VSUBS 0.006961f
C522 B.n469 VSUBS 0.006961f
C523 B.n470 VSUBS 0.006961f
C524 B.n471 VSUBS 0.006961f
C525 B.n472 VSUBS 0.006961f
C526 B.n473 VSUBS 0.006961f
C527 B.n474 VSUBS 0.006961f
C528 B.n475 VSUBS 0.006961f
C529 B.n476 VSUBS 0.006961f
C530 B.n477 VSUBS 0.006961f
C531 B.n478 VSUBS 0.006961f
C532 B.n479 VSUBS 0.006961f
C533 B.n480 VSUBS 0.006961f
C534 B.n481 VSUBS 0.006961f
C535 B.n482 VSUBS 0.006961f
C536 B.n483 VSUBS 0.006961f
C537 B.n484 VSUBS 0.006961f
C538 B.n485 VSUBS 0.006961f
C539 B.n486 VSUBS 0.006961f
C540 B.n487 VSUBS 0.006961f
C541 B.n488 VSUBS 0.006961f
C542 B.n489 VSUBS 0.006961f
C543 B.n490 VSUBS 0.006961f
C544 B.n491 VSUBS 0.006961f
C545 B.n492 VSUBS 0.006961f
C546 B.n493 VSUBS 0.006961f
C547 B.n494 VSUBS 0.006961f
C548 B.n495 VSUBS 0.006961f
C549 B.n496 VSUBS 0.006961f
C550 B.n497 VSUBS 0.006961f
C551 B.n498 VSUBS 0.006961f
C552 B.n499 VSUBS 0.006961f
C553 B.n500 VSUBS 0.006961f
C554 B.n501 VSUBS 0.006961f
C555 B.n502 VSUBS 0.006961f
C556 B.n503 VSUBS 0.006961f
C557 B.n504 VSUBS 0.006961f
C558 B.n505 VSUBS 0.006961f
C559 B.n506 VSUBS 0.006961f
C560 B.n507 VSUBS 0.006961f
C561 B.n508 VSUBS 0.006961f
C562 B.n509 VSUBS 0.006961f
C563 B.n510 VSUBS 0.006961f
C564 B.n511 VSUBS 0.006961f
C565 B.n512 VSUBS 0.006961f
C566 B.n513 VSUBS 0.006961f
C567 B.n514 VSUBS 0.006961f
C568 B.n515 VSUBS 0.006961f
C569 B.n516 VSUBS 0.006961f
C570 B.n517 VSUBS 0.006961f
C571 B.n518 VSUBS 0.006961f
C572 B.n519 VSUBS 0.006961f
C573 B.n520 VSUBS 0.006961f
C574 B.n521 VSUBS 0.004811f
C575 B.n522 VSUBS 0.006961f
C576 B.n523 VSUBS 0.006961f
C577 B.n524 VSUBS 0.00563f
C578 B.n525 VSUBS 0.006961f
C579 B.n526 VSUBS 0.006961f
C580 B.n527 VSUBS 0.006961f
C581 B.n528 VSUBS 0.006961f
C582 B.n529 VSUBS 0.006961f
C583 B.n530 VSUBS 0.006961f
C584 B.n531 VSUBS 0.006961f
C585 B.n532 VSUBS 0.006961f
C586 B.n533 VSUBS 0.006961f
C587 B.n534 VSUBS 0.006961f
C588 B.n535 VSUBS 0.006961f
C589 B.n536 VSUBS 0.00563f
C590 B.n537 VSUBS 0.016128f
C591 B.n538 VSUBS 0.004811f
C592 B.n539 VSUBS 0.006961f
C593 B.n540 VSUBS 0.006961f
C594 B.n541 VSUBS 0.006961f
C595 B.n542 VSUBS 0.006961f
C596 B.n543 VSUBS 0.006961f
C597 B.n544 VSUBS 0.006961f
C598 B.n545 VSUBS 0.006961f
C599 B.n546 VSUBS 0.006961f
C600 B.n547 VSUBS 0.006961f
C601 B.n548 VSUBS 0.006961f
C602 B.n549 VSUBS 0.006961f
C603 B.n550 VSUBS 0.006961f
C604 B.n551 VSUBS 0.006961f
C605 B.n552 VSUBS 0.006961f
C606 B.n553 VSUBS 0.006961f
C607 B.n554 VSUBS 0.006961f
C608 B.n555 VSUBS 0.006961f
C609 B.n556 VSUBS 0.006961f
C610 B.n557 VSUBS 0.006961f
C611 B.n558 VSUBS 0.006961f
C612 B.n559 VSUBS 0.006961f
C613 B.n560 VSUBS 0.006961f
C614 B.n561 VSUBS 0.006961f
C615 B.n562 VSUBS 0.006961f
C616 B.n563 VSUBS 0.006961f
C617 B.n564 VSUBS 0.006961f
C618 B.n565 VSUBS 0.006961f
C619 B.n566 VSUBS 0.006961f
C620 B.n567 VSUBS 0.006961f
C621 B.n568 VSUBS 0.006961f
C622 B.n569 VSUBS 0.006961f
C623 B.n570 VSUBS 0.006961f
C624 B.n571 VSUBS 0.006961f
C625 B.n572 VSUBS 0.006961f
C626 B.n573 VSUBS 0.006961f
C627 B.n574 VSUBS 0.006961f
C628 B.n575 VSUBS 0.006961f
C629 B.n576 VSUBS 0.006961f
C630 B.n577 VSUBS 0.006961f
C631 B.n578 VSUBS 0.006961f
C632 B.n579 VSUBS 0.006961f
C633 B.n580 VSUBS 0.006961f
C634 B.n581 VSUBS 0.006961f
C635 B.n582 VSUBS 0.006961f
C636 B.n583 VSUBS 0.006961f
C637 B.n584 VSUBS 0.006961f
C638 B.n585 VSUBS 0.006961f
C639 B.n586 VSUBS 0.006961f
C640 B.n587 VSUBS 0.006961f
C641 B.n588 VSUBS 0.006961f
C642 B.n589 VSUBS 0.006961f
C643 B.n590 VSUBS 0.006961f
C644 B.n591 VSUBS 0.006961f
C645 B.n592 VSUBS 0.006961f
C646 B.n593 VSUBS 0.006961f
C647 B.n594 VSUBS 0.006961f
C648 B.n595 VSUBS 0.006961f
C649 B.n596 VSUBS 0.006961f
C650 B.n597 VSUBS 0.006961f
C651 B.n598 VSUBS 0.006961f
C652 B.n599 VSUBS 0.006961f
C653 B.n600 VSUBS 0.006961f
C654 B.n601 VSUBS 0.006961f
C655 B.n602 VSUBS 0.006961f
C656 B.n603 VSUBS 0.006961f
C657 B.n604 VSUBS 0.006961f
C658 B.n605 VSUBS 0.006961f
C659 B.n606 VSUBS 0.006961f
C660 B.n607 VSUBS 0.006961f
C661 B.n608 VSUBS 0.006961f
C662 B.n609 VSUBS 0.006961f
C663 B.n610 VSUBS 0.01716f
C664 B.n611 VSUBS 0.016008f
C665 B.n612 VSUBS 0.016008f
C666 B.n613 VSUBS 0.006961f
C667 B.n614 VSUBS 0.006961f
C668 B.n615 VSUBS 0.006961f
C669 B.n616 VSUBS 0.006961f
C670 B.n617 VSUBS 0.006961f
C671 B.n618 VSUBS 0.006961f
C672 B.n619 VSUBS 0.006961f
C673 B.n620 VSUBS 0.006961f
C674 B.n621 VSUBS 0.006961f
C675 B.n622 VSUBS 0.006961f
C676 B.n623 VSUBS 0.006961f
C677 B.n624 VSUBS 0.006961f
C678 B.n625 VSUBS 0.006961f
C679 B.n626 VSUBS 0.006961f
C680 B.n627 VSUBS 0.006961f
C681 B.n628 VSUBS 0.006961f
C682 B.n629 VSUBS 0.006961f
C683 B.n630 VSUBS 0.006961f
C684 B.n631 VSUBS 0.006961f
C685 B.n632 VSUBS 0.006961f
C686 B.n633 VSUBS 0.006961f
C687 B.n634 VSUBS 0.006961f
C688 B.n635 VSUBS 0.006961f
C689 B.n636 VSUBS 0.006961f
C690 B.n637 VSUBS 0.006961f
C691 B.n638 VSUBS 0.006961f
C692 B.n639 VSUBS 0.006961f
C693 B.n640 VSUBS 0.006961f
C694 B.n641 VSUBS 0.006961f
C695 B.n642 VSUBS 0.006961f
C696 B.n643 VSUBS 0.006961f
C697 B.n644 VSUBS 0.006961f
C698 B.n645 VSUBS 0.006961f
C699 B.n646 VSUBS 0.006961f
C700 B.n647 VSUBS 0.006961f
C701 B.n648 VSUBS 0.006961f
C702 B.n649 VSUBS 0.006961f
C703 B.n650 VSUBS 0.006961f
C704 B.n651 VSUBS 0.015762f
C705 VTAIL.t1 VSUBS 2.53839f
C706 VTAIL.n0 VSUBS 0.705793f
C707 VTAIL.t6 VSUBS 2.53839f
C708 VTAIL.n1 VSUBS 0.765362f
C709 VTAIL.t4 VSUBS 2.53839f
C710 VTAIL.n2 VSUBS 2.05785f
C711 VTAIL.t0 VSUBS 2.53841f
C712 VTAIL.n3 VSUBS 2.05783f
C713 VTAIL.t3 VSUBS 2.53841f
C714 VTAIL.n4 VSUBS 0.765342f
C715 VTAIL.t7 VSUBS 2.53841f
C716 VTAIL.n5 VSUBS 0.765342f
C717 VTAIL.t5 VSUBS 2.53839f
C718 VTAIL.n6 VSUBS 2.05785f
C719 VTAIL.t2 VSUBS 2.53839f
C720 VTAIL.n7 VSUBS 1.98988f
C721 VDD1.t1 VSUBS 0.302316f
C722 VDD1.t3 VSUBS 0.302316f
C723 VDD1.n0 VSUBS 2.44635f
C724 VDD1.t2 VSUBS 0.302316f
C725 VDD1.t0 VSUBS 0.302316f
C726 VDD1.n1 VSUBS 3.20895f
C727 VP.n0 VSUBS 0.040291f
C728 VP.t1 VSUBS 2.72802f
C729 VP.n1 VSUBS 0.032604f
C730 VP.n2 VSUBS 0.040291f
C731 VP.t3 VSUBS 2.72802f
C732 VP.t0 VSUBS 2.90046f
C733 VP.t2 VSUBS 2.89836f
C734 VP.n3 VSUBS 3.81393f
C735 VP.n4 VSUBS 2.29696f
C736 VP.n5 VSUBS 1.05015f
C737 VP.n6 VSUBS 0.04007f
C738 VP.n7 VSUBS 0.080505f
C739 VP.n8 VSUBS 0.040291f
C740 VP.n9 VSUBS 0.040291f
C741 VP.n10 VSUBS 0.040291f
C742 VP.n11 VSUBS 0.080505f
C743 VP.n12 VSUBS 0.04007f
C744 VP.n13 VSUBS 1.05015f
C745 VP.n14 VSUBS 0.042977f
.ends

