* NGSPICE file created from diff_pair_sample_1292.ext - technology: sky130A

.subckt diff_pair_sample_1292 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t12 w_n3290_n1970# sky130_fd_pr__pfet_01v8 ad=0.82665 pd=5.34 as=1.9539 ps=10.8 w=5.01 l=1.99
X1 VTAIL.t2 VN.t0 VDD2.t7 w_n3290_n1970# sky130_fd_pr__pfet_01v8 ad=1.9539 pd=10.8 as=0.82665 ps=5.34 w=5.01 l=1.99
X2 VDD2.t6 VN.t1 VTAIL.t1 w_n3290_n1970# sky130_fd_pr__pfet_01v8 ad=0.82665 pd=5.34 as=1.9539 ps=10.8 w=5.01 l=1.99
X3 VTAIL.t4 VN.t2 VDD2.t5 w_n3290_n1970# sky130_fd_pr__pfet_01v8 ad=0.82665 pd=5.34 as=0.82665 ps=5.34 w=5.01 l=1.99
X4 B.t11 B.t9 B.t10 w_n3290_n1970# sky130_fd_pr__pfet_01v8 ad=1.9539 pd=10.8 as=0 ps=0 w=5.01 l=1.99
X5 VDD2.t4 VN.t3 VTAIL.t7 w_n3290_n1970# sky130_fd_pr__pfet_01v8 ad=0.82665 pd=5.34 as=0.82665 ps=5.34 w=5.01 l=1.99
X6 VDD2.t3 VN.t4 VTAIL.t3 w_n3290_n1970# sky130_fd_pr__pfet_01v8 ad=0.82665 pd=5.34 as=1.9539 ps=10.8 w=5.01 l=1.99
X7 VDD1.t6 VP.t1 VTAIL.t10 w_n3290_n1970# sky130_fd_pr__pfet_01v8 ad=0.82665 pd=5.34 as=0.82665 ps=5.34 w=5.01 l=1.99
X8 VDD1.t5 VP.t2 VTAIL.t9 w_n3290_n1970# sky130_fd_pr__pfet_01v8 ad=0.82665 pd=5.34 as=1.9539 ps=10.8 w=5.01 l=1.99
X9 B.t8 B.t6 B.t7 w_n3290_n1970# sky130_fd_pr__pfet_01v8 ad=1.9539 pd=10.8 as=0 ps=0 w=5.01 l=1.99
X10 B.t5 B.t3 B.t4 w_n3290_n1970# sky130_fd_pr__pfet_01v8 ad=1.9539 pd=10.8 as=0 ps=0 w=5.01 l=1.99
X11 VTAIL.t0 VN.t5 VDD2.t2 w_n3290_n1970# sky130_fd_pr__pfet_01v8 ad=0.82665 pd=5.34 as=0.82665 ps=5.34 w=5.01 l=1.99
X12 VDD2.t1 VN.t6 VTAIL.t6 w_n3290_n1970# sky130_fd_pr__pfet_01v8 ad=0.82665 pd=5.34 as=0.82665 ps=5.34 w=5.01 l=1.99
X13 VTAIL.t8 VP.t3 VDD1.t4 w_n3290_n1970# sky130_fd_pr__pfet_01v8 ad=1.9539 pd=10.8 as=0.82665 ps=5.34 w=5.01 l=1.99
X14 VTAIL.t13 VP.t4 VDD1.t3 w_n3290_n1970# sky130_fd_pr__pfet_01v8 ad=1.9539 pd=10.8 as=0.82665 ps=5.34 w=5.01 l=1.99
X15 VTAIL.t11 VP.t5 VDD1.t2 w_n3290_n1970# sky130_fd_pr__pfet_01v8 ad=0.82665 pd=5.34 as=0.82665 ps=5.34 w=5.01 l=1.99
X16 VDD1.t1 VP.t6 VTAIL.t15 w_n3290_n1970# sky130_fd_pr__pfet_01v8 ad=0.82665 pd=5.34 as=0.82665 ps=5.34 w=5.01 l=1.99
X17 VTAIL.t5 VN.t7 VDD2.t0 w_n3290_n1970# sky130_fd_pr__pfet_01v8 ad=1.9539 pd=10.8 as=0.82665 ps=5.34 w=5.01 l=1.99
X18 VTAIL.t14 VP.t7 VDD1.t0 w_n3290_n1970# sky130_fd_pr__pfet_01v8 ad=0.82665 pd=5.34 as=0.82665 ps=5.34 w=5.01 l=1.99
X19 B.t2 B.t0 B.t1 w_n3290_n1970# sky130_fd_pr__pfet_01v8 ad=1.9539 pd=10.8 as=0 ps=0 w=5.01 l=1.99
R0 VP.n14 VP.n11 161.3
R1 VP.n16 VP.n15 161.3
R2 VP.n17 VP.n10 161.3
R3 VP.n19 VP.n18 161.3
R4 VP.n20 VP.n9 161.3
R5 VP.n23 VP.n22 161.3
R6 VP.n24 VP.n8 161.3
R7 VP.n26 VP.n25 161.3
R8 VP.n27 VP.n7 161.3
R9 VP.n52 VP.n0 161.3
R10 VP.n51 VP.n50 161.3
R11 VP.n49 VP.n1 161.3
R12 VP.n48 VP.n47 161.3
R13 VP.n45 VP.n2 161.3
R14 VP.n44 VP.n43 161.3
R15 VP.n42 VP.n3 161.3
R16 VP.n41 VP.n40 161.3
R17 VP.n39 VP.n4 161.3
R18 VP.n37 VP.n36 161.3
R19 VP.n35 VP.n5 161.3
R20 VP.n34 VP.n33 161.3
R21 VP.n32 VP.n6 161.3
R22 VP.n12 VP.t3 91.6439
R23 VP.n31 VP.n30 87.2681
R24 VP.n54 VP.n53 87.2681
R25 VP.n29 VP.n28 87.2681
R26 VP.n13 VP.n12 62.4703
R27 VP.n31 VP.t4 60.6744
R28 VP.n38 VP.t1 60.6744
R29 VP.n46 VP.t7 60.6744
R30 VP.n53 VP.t2 60.6744
R31 VP.n28 VP.t0 60.6744
R32 VP.n21 VP.t5 60.6744
R33 VP.n13 VP.t6 60.6744
R34 VP.n33 VP.n5 56.5193
R35 VP.n26 VP.n8 56.5193
R36 VP.n51 VP.n1 56.5193
R37 VP.n30 VP.n29 42.8253
R38 VP.n40 VP.n3 40.4934
R39 VP.n44 VP.n3 40.4934
R40 VP.n19 VP.n10 40.4934
R41 VP.n15 VP.n10 40.4934
R42 VP.n33 VP.n32 24.4675
R43 VP.n37 VP.n5 24.4675
R44 VP.n40 VP.n39 24.4675
R45 VP.n45 VP.n44 24.4675
R46 VP.n47 VP.n1 24.4675
R47 VP.n52 VP.n51 24.4675
R48 VP.n27 VP.n26 24.4675
R49 VP.n20 VP.n19 24.4675
R50 VP.n22 VP.n8 24.4675
R51 VP.n15 VP.n14 24.4675
R52 VP.n32 VP.n31 23.4888
R53 VP.n53 VP.n52 23.4888
R54 VP.n28 VP.n27 23.4888
R55 VP.n38 VP.n37 16.6381
R56 VP.n47 VP.n46 16.6381
R57 VP.n22 VP.n21 16.6381
R58 VP.n12 VP.n11 12.8111
R59 VP.n39 VP.n38 7.82994
R60 VP.n46 VP.n45 7.82994
R61 VP.n21 VP.n20 7.82994
R62 VP.n14 VP.n13 7.82994
R63 VP.n29 VP.n7 0.278367
R64 VP.n30 VP.n6 0.278367
R65 VP.n54 VP.n0 0.278367
R66 VP.n16 VP.n11 0.189894
R67 VP.n17 VP.n16 0.189894
R68 VP.n18 VP.n17 0.189894
R69 VP.n18 VP.n9 0.189894
R70 VP.n23 VP.n9 0.189894
R71 VP.n24 VP.n23 0.189894
R72 VP.n25 VP.n24 0.189894
R73 VP.n25 VP.n7 0.189894
R74 VP.n34 VP.n6 0.189894
R75 VP.n35 VP.n34 0.189894
R76 VP.n36 VP.n35 0.189894
R77 VP.n36 VP.n4 0.189894
R78 VP.n41 VP.n4 0.189894
R79 VP.n42 VP.n41 0.189894
R80 VP.n43 VP.n42 0.189894
R81 VP.n43 VP.n2 0.189894
R82 VP.n48 VP.n2 0.189894
R83 VP.n49 VP.n48 0.189894
R84 VP.n50 VP.n49 0.189894
R85 VP.n50 VP.n0 0.189894
R86 VP VP.n54 0.153454
R87 VTAIL.n11 VTAIL.t8 91.9954
R88 VTAIL.n10 VTAIL.t1 91.9954
R89 VTAIL.n7 VTAIL.t5 91.9954
R90 VTAIL.n15 VTAIL.t3 91.9953
R91 VTAIL.n2 VTAIL.t2 91.9953
R92 VTAIL.n3 VTAIL.t9 91.9953
R93 VTAIL.n6 VTAIL.t13 91.9953
R94 VTAIL.n14 VTAIL.t12 91.9953
R95 VTAIL.n13 VTAIL.n12 85.5075
R96 VTAIL.n9 VTAIL.n8 85.5075
R97 VTAIL.n1 VTAIL.n0 85.5072
R98 VTAIL.n5 VTAIL.n4 85.5072
R99 VTAIL.n15 VTAIL.n14 18.6858
R100 VTAIL.n7 VTAIL.n6 18.6858
R101 VTAIL.n0 VTAIL.t7 6.48852
R102 VTAIL.n0 VTAIL.t4 6.48852
R103 VTAIL.n4 VTAIL.t10 6.48852
R104 VTAIL.n4 VTAIL.t14 6.48852
R105 VTAIL.n12 VTAIL.t15 6.48852
R106 VTAIL.n12 VTAIL.t11 6.48852
R107 VTAIL.n8 VTAIL.t6 6.48852
R108 VTAIL.n8 VTAIL.t0 6.48852
R109 VTAIL.n9 VTAIL.n7 2.0005
R110 VTAIL.n10 VTAIL.n9 2.0005
R111 VTAIL.n13 VTAIL.n11 2.0005
R112 VTAIL.n14 VTAIL.n13 2.0005
R113 VTAIL.n6 VTAIL.n5 2.0005
R114 VTAIL.n5 VTAIL.n3 2.0005
R115 VTAIL.n2 VTAIL.n1 2.0005
R116 VTAIL VTAIL.n15 1.94231
R117 VTAIL.n11 VTAIL.n10 0.470328
R118 VTAIL.n3 VTAIL.n2 0.470328
R119 VTAIL VTAIL.n1 0.0586897
R120 VDD1 VDD1.n0 103.245
R121 VDD1.n3 VDD1.n2 103.13
R122 VDD1.n3 VDD1.n1 103.13
R123 VDD1.n5 VDD1.n4 102.186
R124 VDD1.n5 VDD1.n3 37.6173
R125 VDD1.n4 VDD1.t2 6.48852
R126 VDD1.n4 VDD1.t7 6.48852
R127 VDD1.n0 VDD1.t4 6.48852
R128 VDD1.n0 VDD1.t1 6.48852
R129 VDD1.n2 VDD1.t0 6.48852
R130 VDD1.n2 VDD1.t5 6.48852
R131 VDD1.n1 VDD1.t3 6.48852
R132 VDD1.n1 VDD1.t6 6.48852
R133 VDD1 VDD1.n5 0.94231
R134 VN.n43 VN.n23 161.3
R135 VN.n42 VN.n41 161.3
R136 VN.n40 VN.n24 161.3
R137 VN.n39 VN.n38 161.3
R138 VN.n36 VN.n25 161.3
R139 VN.n35 VN.n34 161.3
R140 VN.n33 VN.n26 161.3
R141 VN.n32 VN.n31 161.3
R142 VN.n30 VN.n27 161.3
R143 VN.n20 VN.n0 161.3
R144 VN.n19 VN.n18 161.3
R145 VN.n17 VN.n1 161.3
R146 VN.n16 VN.n15 161.3
R147 VN.n13 VN.n2 161.3
R148 VN.n12 VN.n11 161.3
R149 VN.n10 VN.n3 161.3
R150 VN.n9 VN.n8 161.3
R151 VN.n7 VN.n4 161.3
R152 VN.n5 VN.t0 91.6439
R153 VN.n28 VN.t1 91.6439
R154 VN.n22 VN.n21 87.2681
R155 VN.n45 VN.n44 87.2681
R156 VN.n6 VN.n5 62.4703
R157 VN.n29 VN.n28 62.4703
R158 VN.n6 VN.t3 60.6744
R159 VN.n14 VN.t2 60.6744
R160 VN.n21 VN.t4 60.6744
R161 VN.n29 VN.t5 60.6744
R162 VN.n37 VN.t6 60.6744
R163 VN.n44 VN.t7 60.6744
R164 VN.n19 VN.n1 56.5193
R165 VN.n42 VN.n24 56.5193
R166 VN VN.n45 43.1042
R167 VN.n8 VN.n3 40.4934
R168 VN.n12 VN.n3 40.4934
R169 VN.n31 VN.n26 40.4934
R170 VN.n35 VN.n26 40.4934
R171 VN.n8 VN.n7 24.4675
R172 VN.n13 VN.n12 24.4675
R173 VN.n15 VN.n1 24.4675
R174 VN.n20 VN.n19 24.4675
R175 VN.n31 VN.n30 24.4675
R176 VN.n38 VN.n24 24.4675
R177 VN.n36 VN.n35 24.4675
R178 VN.n43 VN.n42 24.4675
R179 VN.n21 VN.n20 23.4888
R180 VN.n44 VN.n43 23.4888
R181 VN.n15 VN.n14 16.6381
R182 VN.n38 VN.n37 16.6381
R183 VN.n28 VN.n27 12.8111
R184 VN.n5 VN.n4 12.8111
R185 VN.n7 VN.n6 7.82994
R186 VN.n14 VN.n13 7.82994
R187 VN.n30 VN.n29 7.82994
R188 VN.n37 VN.n36 7.82994
R189 VN.n45 VN.n23 0.278367
R190 VN.n22 VN.n0 0.278367
R191 VN.n41 VN.n23 0.189894
R192 VN.n41 VN.n40 0.189894
R193 VN.n40 VN.n39 0.189894
R194 VN.n39 VN.n25 0.189894
R195 VN.n34 VN.n25 0.189894
R196 VN.n34 VN.n33 0.189894
R197 VN.n33 VN.n32 0.189894
R198 VN.n32 VN.n27 0.189894
R199 VN.n9 VN.n4 0.189894
R200 VN.n10 VN.n9 0.189894
R201 VN.n11 VN.n10 0.189894
R202 VN.n11 VN.n2 0.189894
R203 VN.n16 VN.n2 0.189894
R204 VN.n17 VN.n16 0.189894
R205 VN.n18 VN.n17 0.189894
R206 VN.n18 VN.n0 0.189894
R207 VN VN.n22 0.153454
R208 VDD2.n2 VDD2.n1 103.13
R209 VDD2.n2 VDD2.n0 103.13
R210 VDD2 VDD2.n5 103.127
R211 VDD2.n4 VDD2.n3 102.186
R212 VDD2.n4 VDD2.n2 37.0343
R213 VDD2.n5 VDD2.t2 6.48852
R214 VDD2.n5 VDD2.t6 6.48852
R215 VDD2.n3 VDD2.t0 6.48852
R216 VDD2.n3 VDD2.t1 6.48852
R217 VDD2.n1 VDD2.t5 6.48852
R218 VDD2.n1 VDD2.t3 6.48852
R219 VDD2.n0 VDD2.t7 6.48852
R220 VDD2.n0 VDD2.t4 6.48852
R221 VDD2 VDD2.n4 1.05869
R222 B.n417 B.n416 585
R223 B.n418 B.n53 585
R224 B.n420 B.n419 585
R225 B.n421 B.n52 585
R226 B.n423 B.n422 585
R227 B.n424 B.n51 585
R228 B.n426 B.n425 585
R229 B.n427 B.n50 585
R230 B.n429 B.n428 585
R231 B.n430 B.n49 585
R232 B.n432 B.n431 585
R233 B.n433 B.n48 585
R234 B.n435 B.n434 585
R235 B.n436 B.n47 585
R236 B.n438 B.n437 585
R237 B.n439 B.n46 585
R238 B.n441 B.n440 585
R239 B.n442 B.n45 585
R240 B.n444 B.n443 585
R241 B.n445 B.n41 585
R242 B.n447 B.n446 585
R243 B.n448 B.n40 585
R244 B.n450 B.n449 585
R245 B.n451 B.n39 585
R246 B.n453 B.n452 585
R247 B.n454 B.n38 585
R248 B.n456 B.n455 585
R249 B.n457 B.n37 585
R250 B.n459 B.n458 585
R251 B.n460 B.n36 585
R252 B.n462 B.n461 585
R253 B.n464 B.n33 585
R254 B.n466 B.n465 585
R255 B.n467 B.n32 585
R256 B.n469 B.n468 585
R257 B.n470 B.n31 585
R258 B.n472 B.n471 585
R259 B.n473 B.n30 585
R260 B.n475 B.n474 585
R261 B.n476 B.n29 585
R262 B.n478 B.n477 585
R263 B.n479 B.n28 585
R264 B.n481 B.n480 585
R265 B.n482 B.n27 585
R266 B.n484 B.n483 585
R267 B.n485 B.n26 585
R268 B.n487 B.n486 585
R269 B.n488 B.n25 585
R270 B.n490 B.n489 585
R271 B.n491 B.n24 585
R272 B.n493 B.n492 585
R273 B.n494 B.n23 585
R274 B.n415 B.n54 585
R275 B.n414 B.n413 585
R276 B.n412 B.n55 585
R277 B.n411 B.n410 585
R278 B.n409 B.n56 585
R279 B.n408 B.n407 585
R280 B.n406 B.n57 585
R281 B.n405 B.n404 585
R282 B.n403 B.n58 585
R283 B.n402 B.n401 585
R284 B.n400 B.n59 585
R285 B.n399 B.n398 585
R286 B.n397 B.n60 585
R287 B.n396 B.n395 585
R288 B.n394 B.n61 585
R289 B.n393 B.n392 585
R290 B.n391 B.n62 585
R291 B.n390 B.n389 585
R292 B.n388 B.n63 585
R293 B.n387 B.n386 585
R294 B.n385 B.n64 585
R295 B.n384 B.n383 585
R296 B.n382 B.n65 585
R297 B.n381 B.n380 585
R298 B.n379 B.n66 585
R299 B.n378 B.n377 585
R300 B.n376 B.n67 585
R301 B.n375 B.n374 585
R302 B.n373 B.n68 585
R303 B.n372 B.n371 585
R304 B.n370 B.n69 585
R305 B.n369 B.n368 585
R306 B.n367 B.n70 585
R307 B.n366 B.n365 585
R308 B.n364 B.n71 585
R309 B.n363 B.n362 585
R310 B.n361 B.n72 585
R311 B.n360 B.n359 585
R312 B.n358 B.n73 585
R313 B.n357 B.n356 585
R314 B.n355 B.n74 585
R315 B.n354 B.n353 585
R316 B.n352 B.n75 585
R317 B.n351 B.n350 585
R318 B.n349 B.n76 585
R319 B.n348 B.n347 585
R320 B.n346 B.n77 585
R321 B.n345 B.n344 585
R322 B.n343 B.n78 585
R323 B.n342 B.n341 585
R324 B.n340 B.n79 585
R325 B.n339 B.n338 585
R326 B.n337 B.n80 585
R327 B.n336 B.n335 585
R328 B.n334 B.n81 585
R329 B.n333 B.n332 585
R330 B.n331 B.n82 585
R331 B.n330 B.n329 585
R332 B.n328 B.n83 585
R333 B.n327 B.n326 585
R334 B.n325 B.n84 585
R335 B.n324 B.n323 585
R336 B.n322 B.n85 585
R337 B.n321 B.n320 585
R338 B.n319 B.n86 585
R339 B.n318 B.n317 585
R340 B.n316 B.n87 585
R341 B.n315 B.n314 585
R342 B.n313 B.n88 585
R343 B.n312 B.n311 585
R344 B.n310 B.n89 585
R345 B.n309 B.n308 585
R346 B.n307 B.n90 585
R347 B.n306 B.n305 585
R348 B.n304 B.n91 585
R349 B.n303 B.n302 585
R350 B.n301 B.n92 585
R351 B.n300 B.n299 585
R352 B.n298 B.n93 585
R353 B.n297 B.n296 585
R354 B.n295 B.n94 585
R355 B.n294 B.n293 585
R356 B.n292 B.n95 585
R357 B.n291 B.n290 585
R358 B.n289 B.n96 585
R359 B.n210 B.n209 585
R360 B.n211 B.n126 585
R361 B.n213 B.n212 585
R362 B.n214 B.n125 585
R363 B.n216 B.n215 585
R364 B.n217 B.n124 585
R365 B.n219 B.n218 585
R366 B.n220 B.n123 585
R367 B.n222 B.n221 585
R368 B.n223 B.n122 585
R369 B.n225 B.n224 585
R370 B.n226 B.n121 585
R371 B.n228 B.n227 585
R372 B.n229 B.n120 585
R373 B.n231 B.n230 585
R374 B.n232 B.n119 585
R375 B.n234 B.n233 585
R376 B.n235 B.n118 585
R377 B.n237 B.n236 585
R378 B.n238 B.n117 585
R379 B.n240 B.n239 585
R380 B.n242 B.n114 585
R381 B.n244 B.n243 585
R382 B.n245 B.n113 585
R383 B.n247 B.n246 585
R384 B.n248 B.n112 585
R385 B.n250 B.n249 585
R386 B.n251 B.n111 585
R387 B.n253 B.n252 585
R388 B.n254 B.n110 585
R389 B.n256 B.n255 585
R390 B.n258 B.n257 585
R391 B.n259 B.n106 585
R392 B.n261 B.n260 585
R393 B.n262 B.n105 585
R394 B.n264 B.n263 585
R395 B.n265 B.n104 585
R396 B.n267 B.n266 585
R397 B.n268 B.n103 585
R398 B.n270 B.n269 585
R399 B.n271 B.n102 585
R400 B.n273 B.n272 585
R401 B.n274 B.n101 585
R402 B.n276 B.n275 585
R403 B.n277 B.n100 585
R404 B.n279 B.n278 585
R405 B.n280 B.n99 585
R406 B.n282 B.n281 585
R407 B.n283 B.n98 585
R408 B.n285 B.n284 585
R409 B.n286 B.n97 585
R410 B.n288 B.n287 585
R411 B.n208 B.n127 585
R412 B.n207 B.n206 585
R413 B.n205 B.n128 585
R414 B.n204 B.n203 585
R415 B.n202 B.n129 585
R416 B.n201 B.n200 585
R417 B.n199 B.n130 585
R418 B.n198 B.n197 585
R419 B.n196 B.n131 585
R420 B.n195 B.n194 585
R421 B.n193 B.n132 585
R422 B.n192 B.n191 585
R423 B.n190 B.n133 585
R424 B.n189 B.n188 585
R425 B.n187 B.n134 585
R426 B.n186 B.n185 585
R427 B.n184 B.n135 585
R428 B.n183 B.n182 585
R429 B.n181 B.n136 585
R430 B.n180 B.n179 585
R431 B.n178 B.n137 585
R432 B.n177 B.n176 585
R433 B.n175 B.n138 585
R434 B.n174 B.n173 585
R435 B.n172 B.n139 585
R436 B.n171 B.n170 585
R437 B.n169 B.n140 585
R438 B.n168 B.n167 585
R439 B.n166 B.n141 585
R440 B.n165 B.n164 585
R441 B.n163 B.n142 585
R442 B.n162 B.n161 585
R443 B.n160 B.n143 585
R444 B.n159 B.n158 585
R445 B.n157 B.n144 585
R446 B.n156 B.n155 585
R447 B.n154 B.n145 585
R448 B.n153 B.n152 585
R449 B.n151 B.n146 585
R450 B.n150 B.n149 585
R451 B.n148 B.n147 585
R452 B.n2 B.n0 585
R453 B.n557 B.n1 585
R454 B.n556 B.n555 585
R455 B.n554 B.n3 585
R456 B.n553 B.n552 585
R457 B.n551 B.n4 585
R458 B.n550 B.n549 585
R459 B.n548 B.n5 585
R460 B.n547 B.n546 585
R461 B.n545 B.n6 585
R462 B.n544 B.n543 585
R463 B.n542 B.n7 585
R464 B.n541 B.n540 585
R465 B.n539 B.n8 585
R466 B.n538 B.n537 585
R467 B.n536 B.n9 585
R468 B.n535 B.n534 585
R469 B.n533 B.n10 585
R470 B.n532 B.n531 585
R471 B.n530 B.n11 585
R472 B.n529 B.n528 585
R473 B.n527 B.n12 585
R474 B.n526 B.n525 585
R475 B.n524 B.n13 585
R476 B.n523 B.n522 585
R477 B.n521 B.n14 585
R478 B.n520 B.n519 585
R479 B.n518 B.n15 585
R480 B.n517 B.n516 585
R481 B.n515 B.n16 585
R482 B.n514 B.n513 585
R483 B.n512 B.n17 585
R484 B.n511 B.n510 585
R485 B.n509 B.n18 585
R486 B.n508 B.n507 585
R487 B.n506 B.n19 585
R488 B.n505 B.n504 585
R489 B.n503 B.n20 585
R490 B.n502 B.n501 585
R491 B.n500 B.n21 585
R492 B.n499 B.n498 585
R493 B.n497 B.n22 585
R494 B.n496 B.n495 585
R495 B.n559 B.n558 585
R496 B.n209 B.n208 511.721
R497 B.n496 B.n23 511.721
R498 B.n287 B.n96 511.721
R499 B.n417 B.n54 511.721
R500 B.n107 B.t0 267.568
R501 B.n115 B.t9 267.568
R502 B.n34 B.t6 267.568
R503 B.n42 B.t3 267.568
R504 B.n107 B.t2 164.349
R505 B.n42 B.t4 164.349
R506 B.n115 B.t11 164.345
R507 B.n34 B.t7 164.345
R508 B.n208 B.n207 163.367
R509 B.n207 B.n128 163.367
R510 B.n203 B.n128 163.367
R511 B.n203 B.n202 163.367
R512 B.n202 B.n201 163.367
R513 B.n201 B.n130 163.367
R514 B.n197 B.n130 163.367
R515 B.n197 B.n196 163.367
R516 B.n196 B.n195 163.367
R517 B.n195 B.n132 163.367
R518 B.n191 B.n132 163.367
R519 B.n191 B.n190 163.367
R520 B.n190 B.n189 163.367
R521 B.n189 B.n134 163.367
R522 B.n185 B.n134 163.367
R523 B.n185 B.n184 163.367
R524 B.n184 B.n183 163.367
R525 B.n183 B.n136 163.367
R526 B.n179 B.n136 163.367
R527 B.n179 B.n178 163.367
R528 B.n178 B.n177 163.367
R529 B.n177 B.n138 163.367
R530 B.n173 B.n138 163.367
R531 B.n173 B.n172 163.367
R532 B.n172 B.n171 163.367
R533 B.n171 B.n140 163.367
R534 B.n167 B.n140 163.367
R535 B.n167 B.n166 163.367
R536 B.n166 B.n165 163.367
R537 B.n165 B.n142 163.367
R538 B.n161 B.n142 163.367
R539 B.n161 B.n160 163.367
R540 B.n160 B.n159 163.367
R541 B.n159 B.n144 163.367
R542 B.n155 B.n144 163.367
R543 B.n155 B.n154 163.367
R544 B.n154 B.n153 163.367
R545 B.n153 B.n146 163.367
R546 B.n149 B.n146 163.367
R547 B.n149 B.n148 163.367
R548 B.n148 B.n2 163.367
R549 B.n558 B.n2 163.367
R550 B.n558 B.n557 163.367
R551 B.n557 B.n556 163.367
R552 B.n556 B.n3 163.367
R553 B.n552 B.n3 163.367
R554 B.n552 B.n551 163.367
R555 B.n551 B.n550 163.367
R556 B.n550 B.n5 163.367
R557 B.n546 B.n5 163.367
R558 B.n546 B.n545 163.367
R559 B.n545 B.n544 163.367
R560 B.n544 B.n7 163.367
R561 B.n540 B.n7 163.367
R562 B.n540 B.n539 163.367
R563 B.n539 B.n538 163.367
R564 B.n538 B.n9 163.367
R565 B.n534 B.n9 163.367
R566 B.n534 B.n533 163.367
R567 B.n533 B.n532 163.367
R568 B.n532 B.n11 163.367
R569 B.n528 B.n11 163.367
R570 B.n528 B.n527 163.367
R571 B.n527 B.n526 163.367
R572 B.n526 B.n13 163.367
R573 B.n522 B.n13 163.367
R574 B.n522 B.n521 163.367
R575 B.n521 B.n520 163.367
R576 B.n520 B.n15 163.367
R577 B.n516 B.n15 163.367
R578 B.n516 B.n515 163.367
R579 B.n515 B.n514 163.367
R580 B.n514 B.n17 163.367
R581 B.n510 B.n17 163.367
R582 B.n510 B.n509 163.367
R583 B.n509 B.n508 163.367
R584 B.n508 B.n19 163.367
R585 B.n504 B.n19 163.367
R586 B.n504 B.n503 163.367
R587 B.n503 B.n502 163.367
R588 B.n502 B.n21 163.367
R589 B.n498 B.n21 163.367
R590 B.n498 B.n497 163.367
R591 B.n497 B.n496 163.367
R592 B.n209 B.n126 163.367
R593 B.n213 B.n126 163.367
R594 B.n214 B.n213 163.367
R595 B.n215 B.n214 163.367
R596 B.n215 B.n124 163.367
R597 B.n219 B.n124 163.367
R598 B.n220 B.n219 163.367
R599 B.n221 B.n220 163.367
R600 B.n221 B.n122 163.367
R601 B.n225 B.n122 163.367
R602 B.n226 B.n225 163.367
R603 B.n227 B.n226 163.367
R604 B.n227 B.n120 163.367
R605 B.n231 B.n120 163.367
R606 B.n232 B.n231 163.367
R607 B.n233 B.n232 163.367
R608 B.n233 B.n118 163.367
R609 B.n237 B.n118 163.367
R610 B.n238 B.n237 163.367
R611 B.n239 B.n238 163.367
R612 B.n239 B.n114 163.367
R613 B.n244 B.n114 163.367
R614 B.n245 B.n244 163.367
R615 B.n246 B.n245 163.367
R616 B.n246 B.n112 163.367
R617 B.n250 B.n112 163.367
R618 B.n251 B.n250 163.367
R619 B.n252 B.n251 163.367
R620 B.n252 B.n110 163.367
R621 B.n256 B.n110 163.367
R622 B.n257 B.n256 163.367
R623 B.n257 B.n106 163.367
R624 B.n261 B.n106 163.367
R625 B.n262 B.n261 163.367
R626 B.n263 B.n262 163.367
R627 B.n263 B.n104 163.367
R628 B.n267 B.n104 163.367
R629 B.n268 B.n267 163.367
R630 B.n269 B.n268 163.367
R631 B.n269 B.n102 163.367
R632 B.n273 B.n102 163.367
R633 B.n274 B.n273 163.367
R634 B.n275 B.n274 163.367
R635 B.n275 B.n100 163.367
R636 B.n279 B.n100 163.367
R637 B.n280 B.n279 163.367
R638 B.n281 B.n280 163.367
R639 B.n281 B.n98 163.367
R640 B.n285 B.n98 163.367
R641 B.n286 B.n285 163.367
R642 B.n287 B.n286 163.367
R643 B.n291 B.n96 163.367
R644 B.n292 B.n291 163.367
R645 B.n293 B.n292 163.367
R646 B.n293 B.n94 163.367
R647 B.n297 B.n94 163.367
R648 B.n298 B.n297 163.367
R649 B.n299 B.n298 163.367
R650 B.n299 B.n92 163.367
R651 B.n303 B.n92 163.367
R652 B.n304 B.n303 163.367
R653 B.n305 B.n304 163.367
R654 B.n305 B.n90 163.367
R655 B.n309 B.n90 163.367
R656 B.n310 B.n309 163.367
R657 B.n311 B.n310 163.367
R658 B.n311 B.n88 163.367
R659 B.n315 B.n88 163.367
R660 B.n316 B.n315 163.367
R661 B.n317 B.n316 163.367
R662 B.n317 B.n86 163.367
R663 B.n321 B.n86 163.367
R664 B.n322 B.n321 163.367
R665 B.n323 B.n322 163.367
R666 B.n323 B.n84 163.367
R667 B.n327 B.n84 163.367
R668 B.n328 B.n327 163.367
R669 B.n329 B.n328 163.367
R670 B.n329 B.n82 163.367
R671 B.n333 B.n82 163.367
R672 B.n334 B.n333 163.367
R673 B.n335 B.n334 163.367
R674 B.n335 B.n80 163.367
R675 B.n339 B.n80 163.367
R676 B.n340 B.n339 163.367
R677 B.n341 B.n340 163.367
R678 B.n341 B.n78 163.367
R679 B.n345 B.n78 163.367
R680 B.n346 B.n345 163.367
R681 B.n347 B.n346 163.367
R682 B.n347 B.n76 163.367
R683 B.n351 B.n76 163.367
R684 B.n352 B.n351 163.367
R685 B.n353 B.n352 163.367
R686 B.n353 B.n74 163.367
R687 B.n357 B.n74 163.367
R688 B.n358 B.n357 163.367
R689 B.n359 B.n358 163.367
R690 B.n359 B.n72 163.367
R691 B.n363 B.n72 163.367
R692 B.n364 B.n363 163.367
R693 B.n365 B.n364 163.367
R694 B.n365 B.n70 163.367
R695 B.n369 B.n70 163.367
R696 B.n370 B.n369 163.367
R697 B.n371 B.n370 163.367
R698 B.n371 B.n68 163.367
R699 B.n375 B.n68 163.367
R700 B.n376 B.n375 163.367
R701 B.n377 B.n376 163.367
R702 B.n377 B.n66 163.367
R703 B.n381 B.n66 163.367
R704 B.n382 B.n381 163.367
R705 B.n383 B.n382 163.367
R706 B.n383 B.n64 163.367
R707 B.n387 B.n64 163.367
R708 B.n388 B.n387 163.367
R709 B.n389 B.n388 163.367
R710 B.n389 B.n62 163.367
R711 B.n393 B.n62 163.367
R712 B.n394 B.n393 163.367
R713 B.n395 B.n394 163.367
R714 B.n395 B.n60 163.367
R715 B.n399 B.n60 163.367
R716 B.n400 B.n399 163.367
R717 B.n401 B.n400 163.367
R718 B.n401 B.n58 163.367
R719 B.n405 B.n58 163.367
R720 B.n406 B.n405 163.367
R721 B.n407 B.n406 163.367
R722 B.n407 B.n56 163.367
R723 B.n411 B.n56 163.367
R724 B.n412 B.n411 163.367
R725 B.n413 B.n412 163.367
R726 B.n413 B.n54 163.367
R727 B.n492 B.n23 163.367
R728 B.n492 B.n491 163.367
R729 B.n491 B.n490 163.367
R730 B.n490 B.n25 163.367
R731 B.n486 B.n25 163.367
R732 B.n486 B.n485 163.367
R733 B.n485 B.n484 163.367
R734 B.n484 B.n27 163.367
R735 B.n480 B.n27 163.367
R736 B.n480 B.n479 163.367
R737 B.n479 B.n478 163.367
R738 B.n478 B.n29 163.367
R739 B.n474 B.n29 163.367
R740 B.n474 B.n473 163.367
R741 B.n473 B.n472 163.367
R742 B.n472 B.n31 163.367
R743 B.n468 B.n31 163.367
R744 B.n468 B.n467 163.367
R745 B.n467 B.n466 163.367
R746 B.n466 B.n33 163.367
R747 B.n461 B.n33 163.367
R748 B.n461 B.n460 163.367
R749 B.n460 B.n459 163.367
R750 B.n459 B.n37 163.367
R751 B.n455 B.n37 163.367
R752 B.n455 B.n454 163.367
R753 B.n454 B.n453 163.367
R754 B.n453 B.n39 163.367
R755 B.n449 B.n39 163.367
R756 B.n449 B.n448 163.367
R757 B.n448 B.n447 163.367
R758 B.n447 B.n41 163.367
R759 B.n443 B.n41 163.367
R760 B.n443 B.n442 163.367
R761 B.n442 B.n441 163.367
R762 B.n441 B.n46 163.367
R763 B.n437 B.n46 163.367
R764 B.n437 B.n436 163.367
R765 B.n436 B.n435 163.367
R766 B.n435 B.n48 163.367
R767 B.n431 B.n48 163.367
R768 B.n431 B.n430 163.367
R769 B.n430 B.n429 163.367
R770 B.n429 B.n50 163.367
R771 B.n425 B.n50 163.367
R772 B.n425 B.n424 163.367
R773 B.n424 B.n423 163.367
R774 B.n423 B.n52 163.367
R775 B.n419 B.n52 163.367
R776 B.n419 B.n418 163.367
R777 B.n418 B.n417 163.367
R778 B.n108 B.t1 119.356
R779 B.n43 B.t5 119.356
R780 B.n116 B.t10 119.35
R781 B.n35 B.t8 119.35
R782 B.n109 B.n108 59.5399
R783 B.n241 B.n116 59.5399
R784 B.n463 B.n35 59.5399
R785 B.n44 B.n43 59.5399
R786 B.n108 B.n107 44.9944
R787 B.n116 B.n115 44.9944
R788 B.n35 B.n34 44.9944
R789 B.n43 B.n42 44.9944
R790 B.n495 B.n494 33.2493
R791 B.n416 B.n415 33.2493
R792 B.n289 B.n288 33.2493
R793 B.n210 B.n127 33.2493
R794 B B.n559 18.0485
R795 B.n494 B.n493 10.6151
R796 B.n493 B.n24 10.6151
R797 B.n489 B.n24 10.6151
R798 B.n489 B.n488 10.6151
R799 B.n488 B.n487 10.6151
R800 B.n487 B.n26 10.6151
R801 B.n483 B.n26 10.6151
R802 B.n483 B.n482 10.6151
R803 B.n482 B.n481 10.6151
R804 B.n481 B.n28 10.6151
R805 B.n477 B.n28 10.6151
R806 B.n477 B.n476 10.6151
R807 B.n476 B.n475 10.6151
R808 B.n475 B.n30 10.6151
R809 B.n471 B.n30 10.6151
R810 B.n471 B.n470 10.6151
R811 B.n470 B.n469 10.6151
R812 B.n469 B.n32 10.6151
R813 B.n465 B.n32 10.6151
R814 B.n465 B.n464 10.6151
R815 B.n462 B.n36 10.6151
R816 B.n458 B.n36 10.6151
R817 B.n458 B.n457 10.6151
R818 B.n457 B.n456 10.6151
R819 B.n456 B.n38 10.6151
R820 B.n452 B.n38 10.6151
R821 B.n452 B.n451 10.6151
R822 B.n451 B.n450 10.6151
R823 B.n450 B.n40 10.6151
R824 B.n446 B.n445 10.6151
R825 B.n445 B.n444 10.6151
R826 B.n444 B.n45 10.6151
R827 B.n440 B.n45 10.6151
R828 B.n440 B.n439 10.6151
R829 B.n439 B.n438 10.6151
R830 B.n438 B.n47 10.6151
R831 B.n434 B.n47 10.6151
R832 B.n434 B.n433 10.6151
R833 B.n433 B.n432 10.6151
R834 B.n432 B.n49 10.6151
R835 B.n428 B.n49 10.6151
R836 B.n428 B.n427 10.6151
R837 B.n427 B.n426 10.6151
R838 B.n426 B.n51 10.6151
R839 B.n422 B.n51 10.6151
R840 B.n422 B.n421 10.6151
R841 B.n421 B.n420 10.6151
R842 B.n420 B.n53 10.6151
R843 B.n416 B.n53 10.6151
R844 B.n290 B.n289 10.6151
R845 B.n290 B.n95 10.6151
R846 B.n294 B.n95 10.6151
R847 B.n295 B.n294 10.6151
R848 B.n296 B.n295 10.6151
R849 B.n296 B.n93 10.6151
R850 B.n300 B.n93 10.6151
R851 B.n301 B.n300 10.6151
R852 B.n302 B.n301 10.6151
R853 B.n302 B.n91 10.6151
R854 B.n306 B.n91 10.6151
R855 B.n307 B.n306 10.6151
R856 B.n308 B.n307 10.6151
R857 B.n308 B.n89 10.6151
R858 B.n312 B.n89 10.6151
R859 B.n313 B.n312 10.6151
R860 B.n314 B.n313 10.6151
R861 B.n314 B.n87 10.6151
R862 B.n318 B.n87 10.6151
R863 B.n319 B.n318 10.6151
R864 B.n320 B.n319 10.6151
R865 B.n320 B.n85 10.6151
R866 B.n324 B.n85 10.6151
R867 B.n325 B.n324 10.6151
R868 B.n326 B.n325 10.6151
R869 B.n326 B.n83 10.6151
R870 B.n330 B.n83 10.6151
R871 B.n331 B.n330 10.6151
R872 B.n332 B.n331 10.6151
R873 B.n332 B.n81 10.6151
R874 B.n336 B.n81 10.6151
R875 B.n337 B.n336 10.6151
R876 B.n338 B.n337 10.6151
R877 B.n338 B.n79 10.6151
R878 B.n342 B.n79 10.6151
R879 B.n343 B.n342 10.6151
R880 B.n344 B.n343 10.6151
R881 B.n344 B.n77 10.6151
R882 B.n348 B.n77 10.6151
R883 B.n349 B.n348 10.6151
R884 B.n350 B.n349 10.6151
R885 B.n350 B.n75 10.6151
R886 B.n354 B.n75 10.6151
R887 B.n355 B.n354 10.6151
R888 B.n356 B.n355 10.6151
R889 B.n356 B.n73 10.6151
R890 B.n360 B.n73 10.6151
R891 B.n361 B.n360 10.6151
R892 B.n362 B.n361 10.6151
R893 B.n362 B.n71 10.6151
R894 B.n366 B.n71 10.6151
R895 B.n367 B.n366 10.6151
R896 B.n368 B.n367 10.6151
R897 B.n368 B.n69 10.6151
R898 B.n372 B.n69 10.6151
R899 B.n373 B.n372 10.6151
R900 B.n374 B.n373 10.6151
R901 B.n374 B.n67 10.6151
R902 B.n378 B.n67 10.6151
R903 B.n379 B.n378 10.6151
R904 B.n380 B.n379 10.6151
R905 B.n380 B.n65 10.6151
R906 B.n384 B.n65 10.6151
R907 B.n385 B.n384 10.6151
R908 B.n386 B.n385 10.6151
R909 B.n386 B.n63 10.6151
R910 B.n390 B.n63 10.6151
R911 B.n391 B.n390 10.6151
R912 B.n392 B.n391 10.6151
R913 B.n392 B.n61 10.6151
R914 B.n396 B.n61 10.6151
R915 B.n397 B.n396 10.6151
R916 B.n398 B.n397 10.6151
R917 B.n398 B.n59 10.6151
R918 B.n402 B.n59 10.6151
R919 B.n403 B.n402 10.6151
R920 B.n404 B.n403 10.6151
R921 B.n404 B.n57 10.6151
R922 B.n408 B.n57 10.6151
R923 B.n409 B.n408 10.6151
R924 B.n410 B.n409 10.6151
R925 B.n410 B.n55 10.6151
R926 B.n414 B.n55 10.6151
R927 B.n415 B.n414 10.6151
R928 B.n211 B.n210 10.6151
R929 B.n212 B.n211 10.6151
R930 B.n212 B.n125 10.6151
R931 B.n216 B.n125 10.6151
R932 B.n217 B.n216 10.6151
R933 B.n218 B.n217 10.6151
R934 B.n218 B.n123 10.6151
R935 B.n222 B.n123 10.6151
R936 B.n223 B.n222 10.6151
R937 B.n224 B.n223 10.6151
R938 B.n224 B.n121 10.6151
R939 B.n228 B.n121 10.6151
R940 B.n229 B.n228 10.6151
R941 B.n230 B.n229 10.6151
R942 B.n230 B.n119 10.6151
R943 B.n234 B.n119 10.6151
R944 B.n235 B.n234 10.6151
R945 B.n236 B.n235 10.6151
R946 B.n236 B.n117 10.6151
R947 B.n240 B.n117 10.6151
R948 B.n243 B.n242 10.6151
R949 B.n243 B.n113 10.6151
R950 B.n247 B.n113 10.6151
R951 B.n248 B.n247 10.6151
R952 B.n249 B.n248 10.6151
R953 B.n249 B.n111 10.6151
R954 B.n253 B.n111 10.6151
R955 B.n254 B.n253 10.6151
R956 B.n255 B.n254 10.6151
R957 B.n259 B.n258 10.6151
R958 B.n260 B.n259 10.6151
R959 B.n260 B.n105 10.6151
R960 B.n264 B.n105 10.6151
R961 B.n265 B.n264 10.6151
R962 B.n266 B.n265 10.6151
R963 B.n266 B.n103 10.6151
R964 B.n270 B.n103 10.6151
R965 B.n271 B.n270 10.6151
R966 B.n272 B.n271 10.6151
R967 B.n272 B.n101 10.6151
R968 B.n276 B.n101 10.6151
R969 B.n277 B.n276 10.6151
R970 B.n278 B.n277 10.6151
R971 B.n278 B.n99 10.6151
R972 B.n282 B.n99 10.6151
R973 B.n283 B.n282 10.6151
R974 B.n284 B.n283 10.6151
R975 B.n284 B.n97 10.6151
R976 B.n288 B.n97 10.6151
R977 B.n206 B.n127 10.6151
R978 B.n206 B.n205 10.6151
R979 B.n205 B.n204 10.6151
R980 B.n204 B.n129 10.6151
R981 B.n200 B.n129 10.6151
R982 B.n200 B.n199 10.6151
R983 B.n199 B.n198 10.6151
R984 B.n198 B.n131 10.6151
R985 B.n194 B.n131 10.6151
R986 B.n194 B.n193 10.6151
R987 B.n193 B.n192 10.6151
R988 B.n192 B.n133 10.6151
R989 B.n188 B.n133 10.6151
R990 B.n188 B.n187 10.6151
R991 B.n187 B.n186 10.6151
R992 B.n186 B.n135 10.6151
R993 B.n182 B.n135 10.6151
R994 B.n182 B.n181 10.6151
R995 B.n181 B.n180 10.6151
R996 B.n180 B.n137 10.6151
R997 B.n176 B.n137 10.6151
R998 B.n176 B.n175 10.6151
R999 B.n175 B.n174 10.6151
R1000 B.n174 B.n139 10.6151
R1001 B.n170 B.n139 10.6151
R1002 B.n170 B.n169 10.6151
R1003 B.n169 B.n168 10.6151
R1004 B.n168 B.n141 10.6151
R1005 B.n164 B.n141 10.6151
R1006 B.n164 B.n163 10.6151
R1007 B.n163 B.n162 10.6151
R1008 B.n162 B.n143 10.6151
R1009 B.n158 B.n143 10.6151
R1010 B.n158 B.n157 10.6151
R1011 B.n157 B.n156 10.6151
R1012 B.n156 B.n145 10.6151
R1013 B.n152 B.n145 10.6151
R1014 B.n152 B.n151 10.6151
R1015 B.n151 B.n150 10.6151
R1016 B.n150 B.n147 10.6151
R1017 B.n147 B.n0 10.6151
R1018 B.n555 B.n1 10.6151
R1019 B.n555 B.n554 10.6151
R1020 B.n554 B.n553 10.6151
R1021 B.n553 B.n4 10.6151
R1022 B.n549 B.n4 10.6151
R1023 B.n549 B.n548 10.6151
R1024 B.n548 B.n547 10.6151
R1025 B.n547 B.n6 10.6151
R1026 B.n543 B.n6 10.6151
R1027 B.n543 B.n542 10.6151
R1028 B.n542 B.n541 10.6151
R1029 B.n541 B.n8 10.6151
R1030 B.n537 B.n8 10.6151
R1031 B.n537 B.n536 10.6151
R1032 B.n536 B.n535 10.6151
R1033 B.n535 B.n10 10.6151
R1034 B.n531 B.n10 10.6151
R1035 B.n531 B.n530 10.6151
R1036 B.n530 B.n529 10.6151
R1037 B.n529 B.n12 10.6151
R1038 B.n525 B.n12 10.6151
R1039 B.n525 B.n524 10.6151
R1040 B.n524 B.n523 10.6151
R1041 B.n523 B.n14 10.6151
R1042 B.n519 B.n14 10.6151
R1043 B.n519 B.n518 10.6151
R1044 B.n518 B.n517 10.6151
R1045 B.n517 B.n16 10.6151
R1046 B.n513 B.n16 10.6151
R1047 B.n513 B.n512 10.6151
R1048 B.n512 B.n511 10.6151
R1049 B.n511 B.n18 10.6151
R1050 B.n507 B.n18 10.6151
R1051 B.n507 B.n506 10.6151
R1052 B.n506 B.n505 10.6151
R1053 B.n505 B.n20 10.6151
R1054 B.n501 B.n20 10.6151
R1055 B.n501 B.n500 10.6151
R1056 B.n500 B.n499 10.6151
R1057 B.n499 B.n22 10.6151
R1058 B.n495 B.n22 10.6151
R1059 B.n464 B.n463 9.36635
R1060 B.n446 B.n44 9.36635
R1061 B.n241 B.n240 9.36635
R1062 B.n258 B.n109 9.36635
R1063 B.n559 B.n0 2.81026
R1064 B.n559 B.n1 2.81026
R1065 B.n463 B.n462 1.24928
R1066 B.n44 B.n40 1.24928
R1067 B.n242 B.n241 1.24928
R1068 B.n255 B.n109 1.24928
C0 VDD1 VTAIL 5.37456f
C1 B VDD2 1.35289f
C2 B VN 1.02529f
C3 w_n3290_n1970# VP 6.82409f
C4 VDD2 VTAIL 5.42489f
C5 w_n3290_n1970# VDD1 1.56972f
C6 VN VTAIL 4.32228f
C7 w_n3290_n1970# VDD2 1.65857f
C8 w_n3290_n1970# VN 6.39886f
C9 VP VDD1 3.97329f
C10 B VTAIL 2.46593f
C11 VDD2 VP 0.459046f
C12 VN VP 5.62148f
C13 w_n3290_n1970# B 7.230411f
C14 VDD2 VDD1 1.46057f
C15 VN VDD1 0.15071f
C16 w_n3290_n1970# VTAIL 2.54738f
C17 B VP 1.73495f
C18 VDD2 VN 3.67035f
C19 B VDD1 1.27597f
C20 VP VTAIL 4.33638f
C21 VDD2 VSUBS 1.375559f
C22 VDD1 VSUBS 1.929234f
C23 VTAIL VSUBS 0.618964f
C24 VN VSUBS 5.65257f
C25 VP VSUBS 2.518093f
C26 B VSUBS 3.527682f
C27 w_n3290_n1970# VSUBS 81.210396f
C28 B.n0 VSUBS 0.005523f
C29 B.n1 VSUBS 0.005523f
C30 B.n2 VSUBS 0.008733f
C31 B.n3 VSUBS 0.008733f
C32 B.n4 VSUBS 0.008733f
C33 B.n5 VSUBS 0.008733f
C34 B.n6 VSUBS 0.008733f
C35 B.n7 VSUBS 0.008733f
C36 B.n8 VSUBS 0.008733f
C37 B.n9 VSUBS 0.008733f
C38 B.n10 VSUBS 0.008733f
C39 B.n11 VSUBS 0.008733f
C40 B.n12 VSUBS 0.008733f
C41 B.n13 VSUBS 0.008733f
C42 B.n14 VSUBS 0.008733f
C43 B.n15 VSUBS 0.008733f
C44 B.n16 VSUBS 0.008733f
C45 B.n17 VSUBS 0.008733f
C46 B.n18 VSUBS 0.008733f
C47 B.n19 VSUBS 0.008733f
C48 B.n20 VSUBS 0.008733f
C49 B.n21 VSUBS 0.008733f
C50 B.n22 VSUBS 0.008733f
C51 B.n23 VSUBS 0.021481f
C52 B.n24 VSUBS 0.008733f
C53 B.n25 VSUBS 0.008733f
C54 B.n26 VSUBS 0.008733f
C55 B.n27 VSUBS 0.008733f
C56 B.n28 VSUBS 0.008733f
C57 B.n29 VSUBS 0.008733f
C58 B.n30 VSUBS 0.008733f
C59 B.n31 VSUBS 0.008733f
C60 B.n32 VSUBS 0.008733f
C61 B.n33 VSUBS 0.008733f
C62 B.t8 VSUBS 0.174482f
C63 B.t7 VSUBS 0.194215f
C64 B.t6 VSUBS 0.585583f
C65 B.n34 VSUBS 0.122169f
C66 B.n35 VSUBS 0.084532f
C67 B.n36 VSUBS 0.008733f
C68 B.n37 VSUBS 0.008733f
C69 B.n38 VSUBS 0.008733f
C70 B.n39 VSUBS 0.008733f
C71 B.n40 VSUBS 0.00488f
C72 B.n41 VSUBS 0.008733f
C73 B.t5 VSUBS 0.174482f
C74 B.t4 VSUBS 0.194215f
C75 B.t3 VSUBS 0.585583f
C76 B.n42 VSUBS 0.12217f
C77 B.n43 VSUBS 0.084532f
C78 B.n44 VSUBS 0.020234f
C79 B.n45 VSUBS 0.008733f
C80 B.n46 VSUBS 0.008733f
C81 B.n47 VSUBS 0.008733f
C82 B.n48 VSUBS 0.008733f
C83 B.n49 VSUBS 0.008733f
C84 B.n50 VSUBS 0.008733f
C85 B.n51 VSUBS 0.008733f
C86 B.n52 VSUBS 0.008733f
C87 B.n53 VSUBS 0.008733f
C88 B.n54 VSUBS 0.019874f
C89 B.n55 VSUBS 0.008733f
C90 B.n56 VSUBS 0.008733f
C91 B.n57 VSUBS 0.008733f
C92 B.n58 VSUBS 0.008733f
C93 B.n59 VSUBS 0.008733f
C94 B.n60 VSUBS 0.008733f
C95 B.n61 VSUBS 0.008733f
C96 B.n62 VSUBS 0.008733f
C97 B.n63 VSUBS 0.008733f
C98 B.n64 VSUBS 0.008733f
C99 B.n65 VSUBS 0.008733f
C100 B.n66 VSUBS 0.008733f
C101 B.n67 VSUBS 0.008733f
C102 B.n68 VSUBS 0.008733f
C103 B.n69 VSUBS 0.008733f
C104 B.n70 VSUBS 0.008733f
C105 B.n71 VSUBS 0.008733f
C106 B.n72 VSUBS 0.008733f
C107 B.n73 VSUBS 0.008733f
C108 B.n74 VSUBS 0.008733f
C109 B.n75 VSUBS 0.008733f
C110 B.n76 VSUBS 0.008733f
C111 B.n77 VSUBS 0.008733f
C112 B.n78 VSUBS 0.008733f
C113 B.n79 VSUBS 0.008733f
C114 B.n80 VSUBS 0.008733f
C115 B.n81 VSUBS 0.008733f
C116 B.n82 VSUBS 0.008733f
C117 B.n83 VSUBS 0.008733f
C118 B.n84 VSUBS 0.008733f
C119 B.n85 VSUBS 0.008733f
C120 B.n86 VSUBS 0.008733f
C121 B.n87 VSUBS 0.008733f
C122 B.n88 VSUBS 0.008733f
C123 B.n89 VSUBS 0.008733f
C124 B.n90 VSUBS 0.008733f
C125 B.n91 VSUBS 0.008733f
C126 B.n92 VSUBS 0.008733f
C127 B.n93 VSUBS 0.008733f
C128 B.n94 VSUBS 0.008733f
C129 B.n95 VSUBS 0.008733f
C130 B.n96 VSUBS 0.019874f
C131 B.n97 VSUBS 0.008733f
C132 B.n98 VSUBS 0.008733f
C133 B.n99 VSUBS 0.008733f
C134 B.n100 VSUBS 0.008733f
C135 B.n101 VSUBS 0.008733f
C136 B.n102 VSUBS 0.008733f
C137 B.n103 VSUBS 0.008733f
C138 B.n104 VSUBS 0.008733f
C139 B.n105 VSUBS 0.008733f
C140 B.n106 VSUBS 0.008733f
C141 B.t1 VSUBS 0.174482f
C142 B.t2 VSUBS 0.194215f
C143 B.t0 VSUBS 0.585583f
C144 B.n107 VSUBS 0.12217f
C145 B.n108 VSUBS 0.084532f
C146 B.n109 VSUBS 0.020234f
C147 B.n110 VSUBS 0.008733f
C148 B.n111 VSUBS 0.008733f
C149 B.n112 VSUBS 0.008733f
C150 B.n113 VSUBS 0.008733f
C151 B.n114 VSUBS 0.008733f
C152 B.t10 VSUBS 0.174482f
C153 B.t11 VSUBS 0.194215f
C154 B.t9 VSUBS 0.585583f
C155 B.n115 VSUBS 0.122169f
C156 B.n116 VSUBS 0.084532f
C157 B.n117 VSUBS 0.008733f
C158 B.n118 VSUBS 0.008733f
C159 B.n119 VSUBS 0.008733f
C160 B.n120 VSUBS 0.008733f
C161 B.n121 VSUBS 0.008733f
C162 B.n122 VSUBS 0.008733f
C163 B.n123 VSUBS 0.008733f
C164 B.n124 VSUBS 0.008733f
C165 B.n125 VSUBS 0.008733f
C166 B.n126 VSUBS 0.008733f
C167 B.n127 VSUBS 0.019874f
C168 B.n128 VSUBS 0.008733f
C169 B.n129 VSUBS 0.008733f
C170 B.n130 VSUBS 0.008733f
C171 B.n131 VSUBS 0.008733f
C172 B.n132 VSUBS 0.008733f
C173 B.n133 VSUBS 0.008733f
C174 B.n134 VSUBS 0.008733f
C175 B.n135 VSUBS 0.008733f
C176 B.n136 VSUBS 0.008733f
C177 B.n137 VSUBS 0.008733f
C178 B.n138 VSUBS 0.008733f
C179 B.n139 VSUBS 0.008733f
C180 B.n140 VSUBS 0.008733f
C181 B.n141 VSUBS 0.008733f
C182 B.n142 VSUBS 0.008733f
C183 B.n143 VSUBS 0.008733f
C184 B.n144 VSUBS 0.008733f
C185 B.n145 VSUBS 0.008733f
C186 B.n146 VSUBS 0.008733f
C187 B.n147 VSUBS 0.008733f
C188 B.n148 VSUBS 0.008733f
C189 B.n149 VSUBS 0.008733f
C190 B.n150 VSUBS 0.008733f
C191 B.n151 VSUBS 0.008733f
C192 B.n152 VSUBS 0.008733f
C193 B.n153 VSUBS 0.008733f
C194 B.n154 VSUBS 0.008733f
C195 B.n155 VSUBS 0.008733f
C196 B.n156 VSUBS 0.008733f
C197 B.n157 VSUBS 0.008733f
C198 B.n158 VSUBS 0.008733f
C199 B.n159 VSUBS 0.008733f
C200 B.n160 VSUBS 0.008733f
C201 B.n161 VSUBS 0.008733f
C202 B.n162 VSUBS 0.008733f
C203 B.n163 VSUBS 0.008733f
C204 B.n164 VSUBS 0.008733f
C205 B.n165 VSUBS 0.008733f
C206 B.n166 VSUBS 0.008733f
C207 B.n167 VSUBS 0.008733f
C208 B.n168 VSUBS 0.008733f
C209 B.n169 VSUBS 0.008733f
C210 B.n170 VSUBS 0.008733f
C211 B.n171 VSUBS 0.008733f
C212 B.n172 VSUBS 0.008733f
C213 B.n173 VSUBS 0.008733f
C214 B.n174 VSUBS 0.008733f
C215 B.n175 VSUBS 0.008733f
C216 B.n176 VSUBS 0.008733f
C217 B.n177 VSUBS 0.008733f
C218 B.n178 VSUBS 0.008733f
C219 B.n179 VSUBS 0.008733f
C220 B.n180 VSUBS 0.008733f
C221 B.n181 VSUBS 0.008733f
C222 B.n182 VSUBS 0.008733f
C223 B.n183 VSUBS 0.008733f
C224 B.n184 VSUBS 0.008733f
C225 B.n185 VSUBS 0.008733f
C226 B.n186 VSUBS 0.008733f
C227 B.n187 VSUBS 0.008733f
C228 B.n188 VSUBS 0.008733f
C229 B.n189 VSUBS 0.008733f
C230 B.n190 VSUBS 0.008733f
C231 B.n191 VSUBS 0.008733f
C232 B.n192 VSUBS 0.008733f
C233 B.n193 VSUBS 0.008733f
C234 B.n194 VSUBS 0.008733f
C235 B.n195 VSUBS 0.008733f
C236 B.n196 VSUBS 0.008733f
C237 B.n197 VSUBS 0.008733f
C238 B.n198 VSUBS 0.008733f
C239 B.n199 VSUBS 0.008733f
C240 B.n200 VSUBS 0.008733f
C241 B.n201 VSUBS 0.008733f
C242 B.n202 VSUBS 0.008733f
C243 B.n203 VSUBS 0.008733f
C244 B.n204 VSUBS 0.008733f
C245 B.n205 VSUBS 0.008733f
C246 B.n206 VSUBS 0.008733f
C247 B.n207 VSUBS 0.008733f
C248 B.n208 VSUBS 0.019874f
C249 B.n209 VSUBS 0.021481f
C250 B.n210 VSUBS 0.021481f
C251 B.n211 VSUBS 0.008733f
C252 B.n212 VSUBS 0.008733f
C253 B.n213 VSUBS 0.008733f
C254 B.n214 VSUBS 0.008733f
C255 B.n215 VSUBS 0.008733f
C256 B.n216 VSUBS 0.008733f
C257 B.n217 VSUBS 0.008733f
C258 B.n218 VSUBS 0.008733f
C259 B.n219 VSUBS 0.008733f
C260 B.n220 VSUBS 0.008733f
C261 B.n221 VSUBS 0.008733f
C262 B.n222 VSUBS 0.008733f
C263 B.n223 VSUBS 0.008733f
C264 B.n224 VSUBS 0.008733f
C265 B.n225 VSUBS 0.008733f
C266 B.n226 VSUBS 0.008733f
C267 B.n227 VSUBS 0.008733f
C268 B.n228 VSUBS 0.008733f
C269 B.n229 VSUBS 0.008733f
C270 B.n230 VSUBS 0.008733f
C271 B.n231 VSUBS 0.008733f
C272 B.n232 VSUBS 0.008733f
C273 B.n233 VSUBS 0.008733f
C274 B.n234 VSUBS 0.008733f
C275 B.n235 VSUBS 0.008733f
C276 B.n236 VSUBS 0.008733f
C277 B.n237 VSUBS 0.008733f
C278 B.n238 VSUBS 0.008733f
C279 B.n239 VSUBS 0.008733f
C280 B.n240 VSUBS 0.00822f
C281 B.n241 VSUBS 0.020234f
C282 B.n242 VSUBS 0.00488f
C283 B.n243 VSUBS 0.008733f
C284 B.n244 VSUBS 0.008733f
C285 B.n245 VSUBS 0.008733f
C286 B.n246 VSUBS 0.008733f
C287 B.n247 VSUBS 0.008733f
C288 B.n248 VSUBS 0.008733f
C289 B.n249 VSUBS 0.008733f
C290 B.n250 VSUBS 0.008733f
C291 B.n251 VSUBS 0.008733f
C292 B.n252 VSUBS 0.008733f
C293 B.n253 VSUBS 0.008733f
C294 B.n254 VSUBS 0.008733f
C295 B.n255 VSUBS 0.00488f
C296 B.n256 VSUBS 0.008733f
C297 B.n257 VSUBS 0.008733f
C298 B.n258 VSUBS 0.00822f
C299 B.n259 VSUBS 0.008733f
C300 B.n260 VSUBS 0.008733f
C301 B.n261 VSUBS 0.008733f
C302 B.n262 VSUBS 0.008733f
C303 B.n263 VSUBS 0.008733f
C304 B.n264 VSUBS 0.008733f
C305 B.n265 VSUBS 0.008733f
C306 B.n266 VSUBS 0.008733f
C307 B.n267 VSUBS 0.008733f
C308 B.n268 VSUBS 0.008733f
C309 B.n269 VSUBS 0.008733f
C310 B.n270 VSUBS 0.008733f
C311 B.n271 VSUBS 0.008733f
C312 B.n272 VSUBS 0.008733f
C313 B.n273 VSUBS 0.008733f
C314 B.n274 VSUBS 0.008733f
C315 B.n275 VSUBS 0.008733f
C316 B.n276 VSUBS 0.008733f
C317 B.n277 VSUBS 0.008733f
C318 B.n278 VSUBS 0.008733f
C319 B.n279 VSUBS 0.008733f
C320 B.n280 VSUBS 0.008733f
C321 B.n281 VSUBS 0.008733f
C322 B.n282 VSUBS 0.008733f
C323 B.n283 VSUBS 0.008733f
C324 B.n284 VSUBS 0.008733f
C325 B.n285 VSUBS 0.008733f
C326 B.n286 VSUBS 0.008733f
C327 B.n287 VSUBS 0.021481f
C328 B.n288 VSUBS 0.021481f
C329 B.n289 VSUBS 0.019874f
C330 B.n290 VSUBS 0.008733f
C331 B.n291 VSUBS 0.008733f
C332 B.n292 VSUBS 0.008733f
C333 B.n293 VSUBS 0.008733f
C334 B.n294 VSUBS 0.008733f
C335 B.n295 VSUBS 0.008733f
C336 B.n296 VSUBS 0.008733f
C337 B.n297 VSUBS 0.008733f
C338 B.n298 VSUBS 0.008733f
C339 B.n299 VSUBS 0.008733f
C340 B.n300 VSUBS 0.008733f
C341 B.n301 VSUBS 0.008733f
C342 B.n302 VSUBS 0.008733f
C343 B.n303 VSUBS 0.008733f
C344 B.n304 VSUBS 0.008733f
C345 B.n305 VSUBS 0.008733f
C346 B.n306 VSUBS 0.008733f
C347 B.n307 VSUBS 0.008733f
C348 B.n308 VSUBS 0.008733f
C349 B.n309 VSUBS 0.008733f
C350 B.n310 VSUBS 0.008733f
C351 B.n311 VSUBS 0.008733f
C352 B.n312 VSUBS 0.008733f
C353 B.n313 VSUBS 0.008733f
C354 B.n314 VSUBS 0.008733f
C355 B.n315 VSUBS 0.008733f
C356 B.n316 VSUBS 0.008733f
C357 B.n317 VSUBS 0.008733f
C358 B.n318 VSUBS 0.008733f
C359 B.n319 VSUBS 0.008733f
C360 B.n320 VSUBS 0.008733f
C361 B.n321 VSUBS 0.008733f
C362 B.n322 VSUBS 0.008733f
C363 B.n323 VSUBS 0.008733f
C364 B.n324 VSUBS 0.008733f
C365 B.n325 VSUBS 0.008733f
C366 B.n326 VSUBS 0.008733f
C367 B.n327 VSUBS 0.008733f
C368 B.n328 VSUBS 0.008733f
C369 B.n329 VSUBS 0.008733f
C370 B.n330 VSUBS 0.008733f
C371 B.n331 VSUBS 0.008733f
C372 B.n332 VSUBS 0.008733f
C373 B.n333 VSUBS 0.008733f
C374 B.n334 VSUBS 0.008733f
C375 B.n335 VSUBS 0.008733f
C376 B.n336 VSUBS 0.008733f
C377 B.n337 VSUBS 0.008733f
C378 B.n338 VSUBS 0.008733f
C379 B.n339 VSUBS 0.008733f
C380 B.n340 VSUBS 0.008733f
C381 B.n341 VSUBS 0.008733f
C382 B.n342 VSUBS 0.008733f
C383 B.n343 VSUBS 0.008733f
C384 B.n344 VSUBS 0.008733f
C385 B.n345 VSUBS 0.008733f
C386 B.n346 VSUBS 0.008733f
C387 B.n347 VSUBS 0.008733f
C388 B.n348 VSUBS 0.008733f
C389 B.n349 VSUBS 0.008733f
C390 B.n350 VSUBS 0.008733f
C391 B.n351 VSUBS 0.008733f
C392 B.n352 VSUBS 0.008733f
C393 B.n353 VSUBS 0.008733f
C394 B.n354 VSUBS 0.008733f
C395 B.n355 VSUBS 0.008733f
C396 B.n356 VSUBS 0.008733f
C397 B.n357 VSUBS 0.008733f
C398 B.n358 VSUBS 0.008733f
C399 B.n359 VSUBS 0.008733f
C400 B.n360 VSUBS 0.008733f
C401 B.n361 VSUBS 0.008733f
C402 B.n362 VSUBS 0.008733f
C403 B.n363 VSUBS 0.008733f
C404 B.n364 VSUBS 0.008733f
C405 B.n365 VSUBS 0.008733f
C406 B.n366 VSUBS 0.008733f
C407 B.n367 VSUBS 0.008733f
C408 B.n368 VSUBS 0.008733f
C409 B.n369 VSUBS 0.008733f
C410 B.n370 VSUBS 0.008733f
C411 B.n371 VSUBS 0.008733f
C412 B.n372 VSUBS 0.008733f
C413 B.n373 VSUBS 0.008733f
C414 B.n374 VSUBS 0.008733f
C415 B.n375 VSUBS 0.008733f
C416 B.n376 VSUBS 0.008733f
C417 B.n377 VSUBS 0.008733f
C418 B.n378 VSUBS 0.008733f
C419 B.n379 VSUBS 0.008733f
C420 B.n380 VSUBS 0.008733f
C421 B.n381 VSUBS 0.008733f
C422 B.n382 VSUBS 0.008733f
C423 B.n383 VSUBS 0.008733f
C424 B.n384 VSUBS 0.008733f
C425 B.n385 VSUBS 0.008733f
C426 B.n386 VSUBS 0.008733f
C427 B.n387 VSUBS 0.008733f
C428 B.n388 VSUBS 0.008733f
C429 B.n389 VSUBS 0.008733f
C430 B.n390 VSUBS 0.008733f
C431 B.n391 VSUBS 0.008733f
C432 B.n392 VSUBS 0.008733f
C433 B.n393 VSUBS 0.008733f
C434 B.n394 VSUBS 0.008733f
C435 B.n395 VSUBS 0.008733f
C436 B.n396 VSUBS 0.008733f
C437 B.n397 VSUBS 0.008733f
C438 B.n398 VSUBS 0.008733f
C439 B.n399 VSUBS 0.008733f
C440 B.n400 VSUBS 0.008733f
C441 B.n401 VSUBS 0.008733f
C442 B.n402 VSUBS 0.008733f
C443 B.n403 VSUBS 0.008733f
C444 B.n404 VSUBS 0.008733f
C445 B.n405 VSUBS 0.008733f
C446 B.n406 VSUBS 0.008733f
C447 B.n407 VSUBS 0.008733f
C448 B.n408 VSUBS 0.008733f
C449 B.n409 VSUBS 0.008733f
C450 B.n410 VSUBS 0.008733f
C451 B.n411 VSUBS 0.008733f
C452 B.n412 VSUBS 0.008733f
C453 B.n413 VSUBS 0.008733f
C454 B.n414 VSUBS 0.008733f
C455 B.n415 VSUBS 0.020887f
C456 B.n416 VSUBS 0.020467f
C457 B.n417 VSUBS 0.021481f
C458 B.n418 VSUBS 0.008733f
C459 B.n419 VSUBS 0.008733f
C460 B.n420 VSUBS 0.008733f
C461 B.n421 VSUBS 0.008733f
C462 B.n422 VSUBS 0.008733f
C463 B.n423 VSUBS 0.008733f
C464 B.n424 VSUBS 0.008733f
C465 B.n425 VSUBS 0.008733f
C466 B.n426 VSUBS 0.008733f
C467 B.n427 VSUBS 0.008733f
C468 B.n428 VSUBS 0.008733f
C469 B.n429 VSUBS 0.008733f
C470 B.n430 VSUBS 0.008733f
C471 B.n431 VSUBS 0.008733f
C472 B.n432 VSUBS 0.008733f
C473 B.n433 VSUBS 0.008733f
C474 B.n434 VSUBS 0.008733f
C475 B.n435 VSUBS 0.008733f
C476 B.n436 VSUBS 0.008733f
C477 B.n437 VSUBS 0.008733f
C478 B.n438 VSUBS 0.008733f
C479 B.n439 VSUBS 0.008733f
C480 B.n440 VSUBS 0.008733f
C481 B.n441 VSUBS 0.008733f
C482 B.n442 VSUBS 0.008733f
C483 B.n443 VSUBS 0.008733f
C484 B.n444 VSUBS 0.008733f
C485 B.n445 VSUBS 0.008733f
C486 B.n446 VSUBS 0.00822f
C487 B.n447 VSUBS 0.008733f
C488 B.n448 VSUBS 0.008733f
C489 B.n449 VSUBS 0.008733f
C490 B.n450 VSUBS 0.008733f
C491 B.n451 VSUBS 0.008733f
C492 B.n452 VSUBS 0.008733f
C493 B.n453 VSUBS 0.008733f
C494 B.n454 VSUBS 0.008733f
C495 B.n455 VSUBS 0.008733f
C496 B.n456 VSUBS 0.008733f
C497 B.n457 VSUBS 0.008733f
C498 B.n458 VSUBS 0.008733f
C499 B.n459 VSUBS 0.008733f
C500 B.n460 VSUBS 0.008733f
C501 B.n461 VSUBS 0.008733f
C502 B.n462 VSUBS 0.00488f
C503 B.n463 VSUBS 0.020234f
C504 B.n464 VSUBS 0.00822f
C505 B.n465 VSUBS 0.008733f
C506 B.n466 VSUBS 0.008733f
C507 B.n467 VSUBS 0.008733f
C508 B.n468 VSUBS 0.008733f
C509 B.n469 VSUBS 0.008733f
C510 B.n470 VSUBS 0.008733f
C511 B.n471 VSUBS 0.008733f
C512 B.n472 VSUBS 0.008733f
C513 B.n473 VSUBS 0.008733f
C514 B.n474 VSUBS 0.008733f
C515 B.n475 VSUBS 0.008733f
C516 B.n476 VSUBS 0.008733f
C517 B.n477 VSUBS 0.008733f
C518 B.n478 VSUBS 0.008733f
C519 B.n479 VSUBS 0.008733f
C520 B.n480 VSUBS 0.008733f
C521 B.n481 VSUBS 0.008733f
C522 B.n482 VSUBS 0.008733f
C523 B.n483 VSUBS 0.008733f
C524 B.n484 VSUBS 0.008733f
C525 B.n485 VSUBS 0.008733f
C526 B.n486 VSUBS 0.008733f
C527 B.n487 VSUBS 0.008733f
C528 B.n488 VSUBS 0.008733f
C529 B.n489 VSUBS 0.008733f
C530 B.n490 VSUBS 0.008733f
C531 B.n491 VSUBS 0.008733f
C532 B.n492 VSUBS 0.008733f
C533 B.n493 VSUBS 0.008733f
C534 B.n494 VSUBS 0.021481f
C535 B.n495 VSUBS 0.019874f
C536 B.n496 VSUBS 0.019874f
C537 B.n497 VSUBS 0.008733f
C538 B.n498 VSUBS 0.008733f
C539 B.n499 VSUBS 0.008733f
C540 B.n500 VSUBS 0.008733f
C541 B.n501 VSUBS 0.008733f
C542 B.n502 VSUBS 0.008733f
C543 B.n503 VSUBS 0.008733f
C544 B.n504 VSUBS 0.008733f
C545 B.n505 VSUBS 0.008733f
C546 B.n506 VSUBS 0.008733f
C547 B.n507 VSUBS 0.008733f
C548 B.n508 VSUBS 0.008733f
C549 B.n509 VSUBS 0.008733f
C550 B.n510 VSUBS 0.008733f
C551 B.n511 VSUBS 0.008733f
C552 B.n512 VSUBS 0.008733f
C553 B.n513 VSUBS 0.008733f
C554 B.n514 VSUBS 0.008733f
C555 B.n515 VSUBS 0.008733f
C556 B.n516 VSUBS 0.008733f
C557 B.n517 VSUBS 0.008733f
C558 B.n518 VSUBS 0.008733f
C559 B.n519 VSUBS 0.008733f
C560 B.n520 VSUBS 0.008733f
C561 B.n521 VSUBS 0.008733f
C562 B.n522 VSUBS 0.008733f
C563 B.n523 VSUBS 0.008733f
C564 B.n524 VSUBS 0.008733f
C565 B.n525 VSUBS 0.008733f
C566 B.n526 VSUBS 0.008733f
C567 B.n527 VSUBS 0.008733f
C568 B.n528 VSUBS 0.008733f
C569 B.n529 VSUBS 0.008733f
C570 B.n530 VSUBS 0.008733f
C571 B.n531 VSUBS 0.008733f
C572 B.n532 VSUBS 0.008733f
C573 B.n533 VSUBS 0.008733f
C574 B.n534 VSUBS 0.008733f
C575 B.n535 VSUBS 0.008733f
C576 B.n536 VSUBS 0.008733f
C577 B.n537 VSUBS 0.008733f
C578 B.n538 VSUBS 0.008733f
C579 B.n539 VSUBS 0.008733f
C580 B.n540 VSUBS 0.008733f
C581 B.n541 VSUBS 0.008733f
C582 B.n542 VSUBS 0.008733f
C583 B.n543 VSUBS 0.008733f
C584 B.n544 VSUBS 0.008733f
C585 B.n545 VSUBS 0.008733f
C586 B.n546 VSUBS 0.008733f
C587 B.n547 VSUBS 0.008733f
C588 B.n548 VSUBS 0.008733f
C589 B.n549 VSUBS 0.008733f
C590 B.n550 VSUBS 0.008733f
C591 B.n551 VSUBS 0.008733f
C592 B.n552 VSUBS 0.008733f
C593 B.n553 VSUBS 0.008733f
C594 B.n554 VSUBS 0.008733f
C595 B.n555 VSUBS 0.008733f
C596 B.n556 VSUBS 0.008733f
C597 B.n557 VSUBS 0.008733f
C598 B.n558 VSUBS 0.008733f
C599 B.n559 VSUBS 0.019775f
C600 VDD2.t7 VSUBS 0.096755f
C601 VDD2.t4 VSUBS 0.096755f
C602 VDD2.n0 VSUBS 0.614874f
C603 VDD2.t5 VSUBS 0.096755f
C604 VDD2.t3 VSUBS 0.096755f
C605 VDD2.n1 VSUBS 0.614874f
C606 VDD2.n2 VSUBS 2.78855f
C607 VDD2.t0 VSUBS 0.096755f
C608 VDD2.t1 VSUBS 0.096755f
C609 VDD2.n3 VSUBS 0.609235f
C610 VDD2.n4 VSUBS 2.31661f
C611 VDD2.t2 VSUBS 0.096755f
C612 VDD2.t6 VSUBS 0.096755f
C613 VDD2.n5 VSUBS 0.614849f
C614 VN.n0 VSUBS 0.05678f
C615 VN.t4 VSUBS 1.12326f
C616 VN.n1 VSUBS 0.071272f
C617 VN.n2 VSUBS 0.043068f
C618 VN.t2 VSUBS 1.12326f
C619 VN.n3 VSUBS 0.034816f
C620 VN.n4 VSUBS 0.321769f
C621 VN.t3 VSUBS 1.12326f
C622 VN.t0 VSUBS 1.34514f
C623 VN.n5 VSUBS 0.544426f
C624 VN.n6 VSUBS 0.536992f
C625 VN.n7 VSUBS 0.05332f
C626 VN.n8 VSUBS 0.085597f
C627 VN.n9 VSUBS 0.043068f
C628 VN.n10 VSUBS 0.043068f
C629 VN.n11 VSUBS 0.043068f
C630 VN.n12 VSUBS 0.085597f
C631 VN.n13 VSUBS 0.05332f
C632 VN.n14 VSUBS 0.440737f
C633 VN.n15 VSUBS 0.067586f
C634 VN.n16 VSUBS 0.043068f
C635 VN.n17 VSUBS 0.043068f
C636 VN.n18 VSUBS 0.043068f
C637 VN.n19 VSUBS 0.05447f
C638 VN.n20 VSUBS 0.078682f
C639 VN.n21 VSUBS 0.582022f
C640 VN.n22 VSUBS 0.047221f
C641 VN.n23 VSUBS 0.05678f
C642 VN.t7 VSUBS 1.12326f
C643 VN.n24 VSUBS 0.071272f
C644 VN.n25 VSUBS 0.043068f
C645 VN.t6 VSUBS 1.12326f
C646 VN.n26 VSUBS 0.034816f
C647 VN.n27 VSUBS 0.321769f
C648 VN.t5 VSUBS 1.12326f
C649 VN.t1 VSUBS 1.34514f
C650 VN.n28 VSUBS 0.544426f
C651 VN.n29 VSUBS 0.536992f
C652 VN.n30 VSUBS 0.05332f
C653 VN.n31 VSUBS 0.085597f
C654 VN.n32 VSUBS 0.043068f
C655 VN.n33 VSUBS 0.043068f
C656 VN.n34 VSUBS 0.043068f
C657 VN.n35 VSUBS 0.085597f
C658 VN.n36 VSUBS 0.05332f
C659 VN.n37 VSUBS 0.440737f
C660 VN.n38 VSUBS 0.067586f
C661 VN.n39 VSUBS 0.043068f
C662 VN.n40 VSUBS 0.043068f
C663 VN.n41 VSUBS 0.043068f
C664 VN.n42 VSUBS 0.05447f
C665 VN.n43 VSUBS 0.078682f
C666 VN.n44 VSUBS 0.582022f
C667 VN.n45 VSUBS 1.89162f
C668 VDD1.t4 VSUBS 0.098963f
C669 VDD1.t1 VSUBS 0.098963f
C670 VDD1.n0 VSUBS 0.629683f
C671 VDD1.t3 VSUBS 0.098963f
C672 VDD1.t6 VSUBS 0.098963f
C673 VDD1.n1 VSUBS 0.628906f
C674 VDD1.t0 VSUBS 0.098963f
C675 VDD1.t5 VSUBS 0.098963f
C676 VDD1.n2 VSUBS 0.628906f
C677 VDD1.n3 VSUBS 2.90483f
C678 VDD1.t2 VSUBS 0.098963f
C679 VDD1.t7 VSUBS 0.098963f
C680 VDD1.n4 VSUBS 0.623135f
C681 VDD1.n5 VSUBS 2.39979f
C682 VTAIL.t7 VSUBS 0.116488f
C683 VTAIL.t4 VSUBS 0.116488f
C684 VTAIL.n0 VSUBS 0.646849f
C685 VTAIL.n1 VSUBS 0.691568f
C686 VTAIL.t2 VSUBS 0.904734f
C687 VTAIL.n2 VSUBS 0.790405f
C688 VTAIL.t9 VSUBS 0.904734f
C689 VTAIL.n3 VSUBS 0.790405f
C690 VTAIL.t10 VSUBS 0.116488f
C691 VTAIL.t14 VSUBS 0.116488f
C692 VTAIL.n4 VSUBS 0.646849f
C693 VTAIL.n5 VSUBS 0.875668f
C694 VTAIL.t13 VSUBS 0.904734f
C695 VTAIL.n6 VSUBS 1.74463f
C696 VTAIL.t5 VSUBS 0.904739f
C697 VTAIL.n7 VSUBS 1.74463f
C698 VTAIL.t6 VSUBS 0.116488f
C699 VTAIL.t0 VSUBS 0.116488f
C700 VTAIL.n8 VSUBS 0.646852f
C701 VTAIL.n9 VSUBS 0.875664f
C702 VTAIL.t1 VSUBS 0.904739f
C703 VTAIL.n10 VSUBS 0.7904f
C704 VTAIL.t8 VSUBS 0.904739f
C705 VTAIL.n11 VSUBS 0.7904f
C706 VTAIL.t15 VSUBS 0.116488f
C707 VTAIL.t11 VSUBS 0.116488f
C708 VTAIL.n12 VSUBS 0.646852f
C709 VTAIL.n13 VSUBS 0.875664f
C710 VTAIL.t12 VSUBS 0.904734f
C711 VTAIL.n14 VSUBS 1.74463f
C712 VTAIL.t3 VSUBS 0.904734f
C713 VTAIL.n15 VSUBS 1.73912f
C714 VP.n0 VSUBS 0.058946f
C715 VP.t2 VSUBS 1.16611f
C716 VP.n1 VSUBS 0.07399f
C717 VP.n2 VSUBS 0.04471f
C718 VP.t7 VSUBS 1.16611f
C719 VP.n3 VSUBS 0.036144f
C720 VP.n4 VSUBS 0.04471f
C721 VP.t1 VSUBS 1.16611f
C722 VP.n5 VSUBS 0.07399f
C723 VP.n6 VSUBS 0.058946f
C724 VP.t4 VSUBS 1.16611f
C725 VP.n7 VSUBS 0.058946f
C726 VP.t0 VSUBS 1.16611f
C727 VP.n8 VSUBS 0.07399f
C728 VP.n9 VSUBS 0.04471f
C729 VP.t5 VSUBS 1.16611f
C730 VP.n10 VSUBS 0.036144f
C731 VP.n11 VSUBS 0.334043f
C732 VP.t6 VSUBS 1.16611f
C733 VP.t3 VSUBS 1.39645f
C734 VP.n12 VSUBS 0.565191f
C735 VP.n13 VSUBS 0.557474f
C736 VP.n14 VSUBS 0.055354f
C737 VP.n15 VSUBS 0.088862f
C738 VP.n16 VSUBS 0.04471f
C739 VP.n17 VSUBS 0.04471f
C740 VP.n18 VSUBS 0.04471f
C741 VP.n19 VSUBS 0.088862f
C742 VP.n20 VSUBS 0.055354f
C743 VP.n21 VSUBS 0.457548f
C744 VP.n22 VSUBS 0.070164f
C745 VP.n23 VSUBS 0.04471f
C746 VP.n24 VSUBS 0.04471f
C747 VP.n25 VSUBS 0.04471f
C748 VP.n26 VSUBS 0.056548f
C749 VP.n27 VSUBS 0.081683f
C750 VP.n28 VSUBS 0.604222f
C751 VP.n29 VSUBS 1.93911f
C752 VP.n30 VSUBS 1.97664f
C753 VP.n31 VSUBS 0.604222f
C754 VP.n32 VSUBS 0.081683f
C755 VP.n33 VSUBS 0.056548f
C756 VP.n34 VSUBS 0.04471f
C757 VP.n35 VSUBS 0.04471f
C758 VP.n36 VSUBS 0.04471f
C759 VP.n37 VSUBS 0.070164f
C760 VP.n38 VSUBS 0.457548f
C761 VP.n39 VSUBS 0.055354f
C762 VP.n40 VSUBS 0.088862f
C763 VP.n41 VSUBS 0.04471f
C764 VP.n42 VSUBS 0.04471f
C765 VP.n43 VSUBS 0.04471f
C766 VP.n44 VSUBS 0.088862f
C767 VP.n45 VSUBS 0.055354f
C768 VP.n46 VSUBS 0.457548f
C769 VP.n47 VSUBS 0.070164f
C770 VP.n48 VSUBS 0.04471f
C771 VP.n49 VSUBS 0.04471f
C772 VP.n50 VSUBS 0.04471f
C773 VP.n51 VSUBS 0.056548f
C774 VP.n52 VSUBS 0.081683f
C775 VP.n53 VSUBS 0.604222f
C776 VP.n54 VSUBS 0.049022f
.ends

