* NGSPICE file created from diff_pair_sample_1357.ext - technology: sky130A

.subckt diff_pair_sample_1357 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=4.5123 pd=23.92 as=0 ps=0 w=11.57 l=3.14
X1 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=4.5123 pd=23.92 as=4.5123 ps=23.92 w=11.57 l=3.14
X2 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=4.5123 pd=23.92 as=0 ps=0 w=11.57 l=3.14
X3 VDD1.t1 VP.t0 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=4.5123 pd=23.92 as=4.5123 ps=23.92 w=11.57 l=3.14
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.5123 pd=23.92 as=0 ps=0 w=11.57 l=3.14
X5 VDD1.t0 VP.t1 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=4.5123 pd=23.92 as=4.5123 ps=23.92 w=11.57 l=3.14
X6 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=4.5123 pd=23.92 as=4.5123 ps=23.92 w=11.57 l=3.14
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.5123 pd=23.92 as=0 ps=0 w=11.57 l=3.14
R0 B.n689 B.n688 585
R1 B.n281 B.n100 585
R2 B.n280 B.n279 585
R3 B.n278 B.n277 585
R4 B.n276 B.n275 585
R5 B.n274 B.n273 585
R6 B.n272 B.n271 585
R7 B.n270 B.n269 585
R8 B.n268 B.n267 585
R9 B.n266 B.n265 585
R10 B.n264 B.n263 585
R11 B.n262 B.n261 585
R12 B.n260 B.n259 585
R13 B.n258 B.n257 585
R14 B.n256 B.n255 585
R15 B.n254 B.n253 585
R16 B.n252 B.n251 585
R17 B.n250 B.n249 585
R18 B.n248 B.n247 585
R19 B.n246 B.n245 585
R20 B.n244 B.n243 585
R21 B.n242 B.n241 585
R22 B.n240 B.n239 585
R23 B.n238 B.n237 585
R24 B.n236 B.n235 585
R25 B.n234 B.n233 585
R26 B.n232 B.n231 585
R27 B.n230 B.n229 585
R28 B.n228 B.n227 585
R29 B.n226 B.n225 585
R30 B.n224 B.n223 585
R31 B.n222 B.n221 585
R32 B.n220 B.n219 585
R33 B.n218 B.n217 585
R34 B.n216 B.n215 585
R35 B.n214 B.n213 585
R36 B.n212 B.n211 585
R37 B.n210 B.n209 585
R38 B.n208 B.n207 585
R39 B.n206 B.n205 585
R40 B.n204 B.n203 585
R41 B.n202 B.n201 585
R42 B.n200 B.n199 585
R43 B.n198 B.n197 585
R44 B.n196 B.n195 585
R45 B.n194 B.n193 585
R46 B.n192 B.n191 585
R47 B.n190 B.n189 585
R48 B.n188 B.n187 585
R49 B.n186 B.n185 585
R50 B.n184 B.n183 585
R51 B.n182 B.n181 585
R52 B.n180 B.n179 585
R53 B.n178 B.n177 585
R54 B.n176 B.n175 585
R55 B.n174 B.n173 585
R56 B.n172 B.n171 585
R57 B.n170 B.n169 585
R58 B.n168 B.n167 585
R59 B.n166 B.n165 585
R60 B.n164 B.n163 585
R61 B.n162 B.n161 585
R62 B.n160 B.n159 585
R63 B.n158 B.n157 585
R64 B.n156 B.n155 585
R65 B.n154 B.n153 585
R66 B.n152 B.n151 585
R67 B.n150 B.n149 585
R68 B.n148 B.n147 585
R69 B.n146 B.n145 585
R70 B.n144 B.n143 585
R71 B.n142 B.n141 585
R72 B.n140 B.n139 585
R73 B.n138 B.n137 585
R74 B.n136 B.n135 585
R75 B.n134 B.n133 585
R76 B.n132 B.n131 585
R77 B.n130 B.n129 585
R78 B.n128 B.n127 585
R79 B.n126 B.n125 585
R80 B.n124 B.n123 585
R81 B.n122 B.n121 585
R82 B.n120 B.n119 585
R83 B.n118 B.n117 585
R84 B.n116 B.n115 585
R85 B.n114 B.n113 585
R86 B.n112 B.n111 585
R87 B.n110 B.n109 585
R88 B.n108 B.n107 585
R89 B.n54 B.n53 585
R90 B.n687 B.n55 585
R91 B.n692 B.n55 585
R92 B.n686 B.n685 585
R93 B.n685 B.n51 585
R94 B.n684 B.n50 585
R95 B.n698 B.n50 585
R96 B.n683 B.n49 585
R97 B.n699 B.n49 585
R98 B.n682 B.n48 585
R99 B.n700 B.n48 585
R100 B.n681 B.n680 585
R101 B.n680 B.n44 585
R102 B.n679 B.n43 585
R103 B.n706 B.n43 585
R104 B.n678 B.n42 585
R105 B.n707 B.n42 585
R106 B.n677 B.n41 585
R107 B.n708 B.n41 585
R108 B.n676 B.n675 585
R109 B.n675 B.n37 585
R110 B.n674 B.n36 585
R111 B.n714 B.n36 585
R112 B.n673 B.n35 585
R113 B.n715 B.n35 585
R114 B.n672 B.n34 585
R115 B.n716 B.n34 585
R116 B.n671 B.n670 585
R117 B.n670 B.n30 585
R118 B.n669 B.n29 585
R119 B.n722 B.n29 585
R120 B.n668 B.n28 585
R121 B.n723 B.n28 585
R122 B.n667 B.n27 585
R123 B.n724 B.n27 585
R124 B.n666 B.n665 585
R125 B.n665 B.n23 585
R126 B.n664 B.n22 585
R127 B.n730 B.n22 585
R128 B.n663 B.n21 585
R129 B.n731 B.n21 585
R130 B.n662 B.n20 585
R131 B.n732 B.n20 585
R132 B.n661 B.n660 585
R133 B.n660 B.n19 585
R134 B.n659 B.n15 585
R135 B.n738 B.n15 585
R136 B.n658 B.n14 585
R137 B.n739 B.n14 585
R138 B.n657 B.n13 585
R139 B.n740 B.n13 585
R140 B.n656 B.n655 585
R141 B.n655 B.n12 585
R142 B.n654 B.n653 585
R143 B.n654 B.n8 585
R144 B.n652 B.n7 585
R145 B.n747 B.n7 585
R146 B.n651 B.n6 585
R147 B.n748 B.n6 585
R148 B.n650 B.n5 585
R149 B.n749 B.n5 585
R150 B.n649 B.n648 585
R151 B.n648 B.n4 585
R152 B.n647 B.n282 585
R153 B.n647 B.n646 585
R154 B.n637 B.n283 585
R155 B.n284 B.n283 585
R156 B.n639 B.n638 585
R157 B.n640 B.n639 585
R158 B.n636 B.n289 585
R159 B.n289 B.n288 585
R160 B.n635 B.n634 585
R161 B.n634 B.n633 585
R162 B.n291 B.n290 585
R163 B.n626 B.n291 585
R164 B.n625 B.n624 585
R165 B.n627 B.n625 585
R166 B.n623 B.n296 585
R167 B.n296 B.n295 585
R168 B.n622 B.n621 585
R169 B.n621 B.n620 585
R170 B.n298 B.n297 585
R171 B.n299 B.n298 585
R172 B.n613 B.n612 585
R173 B.n614 B.n613 585
R174 B.n611 B.n304 585
R175 B.n304 B.n303 585
R176 B.n610 B.n609 585
R177 B.n609 B.n608 585
R178 B.n306 B.n305 585
R179 B.n307 B.n306 585
R180 B.n601 B.n600 585
R181 B.n602 B.n601 585
R182 B.n599 B.n312 585
R183 B.n312 B.n311 585
R184 B.n598 B.n597 585
R185 B.n597 B.n596 585
R186 B.n314 B.n313 585
R187 B.n315 B.n314 585
R188 B.n589 B.n588 585
R189 B.n590 B.n589 585
R190 B.n587 B.n320 585
R191 B.n320 B.n319 585
R192 B.n586 B.n585 585
R193 B.n585 B.n584 585
R194 B.n322 B.n321 585
R195 B.n323 B.n322 585
R196 B.n577 B.n576 585
R197 B.n578 B.n577 585
R198 B.n575 B.n328 585
R199 B.n328 B.n327 585
R200 B.n574 B.n573 585
R201 B.n573 B.n572 585
R202 B.n330 B.n329 585
R203 B.n331 B.n330 585
R204 B.n565 B.n564 585
R205 B.n566 B.n565 585
R206 B.n334 B.n333 585
R207 B.n385 B.n383 585
R208 B.n386 B.n382 585
R209 B.n386 B.n335 585
R210 B.n389 B.n388 585
R211 B.n390 B.n381 585
R212 B.n392 B.n391 585
R213 B.n394 B.n380 585
R214 B.n397 B.n396 585
R215 B.n398 B.n379 585
R216 B.n400 B.n399 585
R217 B.n402 B.n378 585
R218 B.n405 B.n404 585
R219 B.n406 B.n377 585
R220 B.n408 B.n407 585
R221 B.n410 B.n376 585
R222 B.n413 B.n412 585
R223 B.n414 B.n375 585
R224 B.n416 B.n415 585
R225 B.n418 B.n374 585
R226 B.n421 B.n420 585
R227 B.n422 B.n373 585
R228 B.n424 B.n423 585
R229 B.n426 B.n372 585
R230 B.n429 B.n428 585
R231 B.n430 B.n371 585
R232 B.n432 B.n431 585
R233 B.n434 B.n370 585
R234 B.n437 B.n436 585
R235 B.n438 B.n369 585
R236 B.n440 B.n439 585
R237 B.n442 B.n368 585
R238 B.n445 B.n444 585
R239 B.n446 B.n367 585
R240 B.n448 B.n447 585
R241 B.n450 B.n366 585
R242 B.n453 B.n452 585
R243 B.n454 B.n365 585
R244 B.n456 B.n455 585
R245 B.n458 B.n364 585
R246 B.n461 B.n460 585
R247 B.n463 B.n361 585
R248 B.n465 B.n464 585
R249 B.n467 B.n360 585
R250 B.n470 B.n469 585
R251 B.n471 B.n359 585
R252 B.n473 B.n472 585
R253 B.n475 B.n358 585
R254 B.n478 B.n477 585
R255 B.n479 B.n357 585
R256 B.n484 B.n483 585
R257 B.n486 B.n356 585
R258 B.n489 B.n488 585
R259 B.n490 B.n355 585
R260 B.n492 B.n491 585
R261 B.n494 B.n354 585
R262 B.n497 B.n496 585
R263 B.n498 B.n353 585
R264 B.n500 B.n499 585
R265 B.n502 B.n352 585
R266 B.n505 B.n504 585
R267 B.n506 B.n351 585
R268 B.n508 B.n507 585
R269 B.n510 B.n350 585
R270 B.n513 B.n512 585
R271 B.n514 B.n349 585
R272 B.n516 B.n515 585
R273 B.n518 B.n348 585
R274 B.n521 B.n520 585
R275 B.n522 B.n347 585
R276 B.n524 B.n523 585
R277 B.n526 B.n346 585
R278 B.n529 B.n528 585
R279 B.n530 B.n345 585
R280 B.n532 B.n531 585
R281 B.n534 B.n344 585
R282 B.n537 B.n536 585
R283 B.n538 B.n343 585
R284 B.n540 B.n539 585
R285 B.n542 B.n342 585
R286 B.n545 B.n544 585
R287 B.n546 B.n341 585
R288 B.n548 B.n547 585
R289 B.n550 B.n340 585
R290 B.n553 B.n552 585
R291 B.n554 B.n339 585
R292 B.n556 B.n555 585
R293 B.n558 B.n338 585
R294 B.n559 B.n337 585
R295 B.n562 B.n561 585
R296 B.n563 B.n336 585
R297 B.n336 B.n335 585
R298 B.n568 B.n567 585
R299 B.n567 B.n566 585
R300 B.n569 B.n332 585
R301 B.n332 B.n331 585
R302 B.n571 B.n570 585
R303 B.n572 B.n571 585
R304 B.n326 B.n325 585
R305 B.n327 B.n326 585
R306 B.n580 B.n579 585
R307 B.n579 B.n578 585
R308 B.n581 B.n324 585
R309 B.n324 B.n323 585
R310 B.n583 B.n582 585
R311 B.n584 B.n583 585
R312 B.n318 B.n317 585
R313 B.n319 B.n318 585
R314 B.n592 B.n591 585
R315 B.n591 B.n590 585
R316 B.n593 B.n316 585
R317 B.n316 B.n315 585
R318 B.n595 B.n594 585
R319 B.n596 B.n595 585
R320 B.n310 B.n309 585
R321 B.n311 B.n310 585
R322 B.n604 B.n603 585
R323 B.n603 B.n602 585
R324 B.n605 B.n308 585
R325 B.n308 B.n307 585
R326 B.n607 B.n606 585
R327 B.n608 B.n607 585
R328 B.n302 B.n301 585
R329 B.n303 B.n302 585
R330 B.n616 B.n615 585
R331 B.n615 B.n614 585
R332 B.n617 B.n300 585
R333 B.n300 B.n299 585
R334 B.n619 B.n618 585
R335 B.n620 B.n619 585
R336 B.n294 B.n293 585
R337 B.n295 B.n294 585
R338 B.n629 B.n628 585
R339 B.n628 B.n627 585
R340 B.n630 B.n292 585
R341 B.n626 B.n292 585
R342 B.n632 B.n631 585
R343 B.n633 B.n632 585
R344 B.n287 B.n286 585
R345 B.n288 B.n287 585
R346 B.n642 B.n641 585
R347 B.n641 B.n640 585
R348 B.n643 B.n285 585
R349 B.n285 B.n284 585
R350 B.n645 B.n644 585
R351 B.n646 B.n645 585
R352 B.n3 B.n0 585
R353 B.n4 B.n3 585
R354 B.n746 B.n1 585
R355 B.n747 B.n746 585
R356 B.n745 B.n744 585
R357 B.n745 B.n8 585
R358 B.n743 B.n9 585
R359 B.n12 B.n9 585
R360 B.n742 B.n741 585
R361 B.n741 B.n740 585
R362 B.n11 B.n10 585
R363 B.n739 B.n11 585
R364 B.n737 B.n736 585
R365 B.n738 B.n737 585
R366 B.n735 B.n16 585
R367 B.n19 B.n16 585
R368 B.n734 B.n733 585
R369 B.n733 B.n732 585
R370 B.n18 B.n17 585
R371 B.n731 B.n18 585
R372 B.n729 B.n728 585
R373 B.n730 B.n729 585
R374 B.n727 B.n24 585
R375 B.n24 B.n23 585
R376 B.n726 B.n725 585
R377 B.n725 B.n724 585
R378 B.n26 B.n25 585
R379 B.n723 B.n26 585
R380 B.n721 B.n720 585
R381 B.n722 B.n721 585
R382 B.n719 B.n31 585
R383 B.n31 B.n30 585
R384 B.n718 B.n717 585
R385 B.n717 B.n716 585
R386 B.n33 B.n32 585
R387 B.n715 B.n33 585
R388 B.n713 B.n712 585
R389 B.n714 B.n713 585
R390 B.n711 B.n38 585
R391 B.n38 B.n37 585
R392 B.n710 B.n709 585
R393 B.n709 B.n708 585
R394 B.n40 B.n39 585
R395 B.n707 B.n40 585
R396 B.n705 B.n704 585
R397 B.n706 B.n705 585
R398 B.n703 B.n45 585
R399 B.n45 B.n44 585
R400 B.n702 B.n701 585
R401 B.n701 B.n700 585
R402 B.n47 B.n46 585
R403 B.n699 B.n47 585
R404 B.n697 B.n696 585
R405 B.n698 B.n697 585
R406 B.n695 B.n52 585
R407 B.n52 B.n51 585
R408 B.n694 B.n693 585
R409 B.n693 B.n692 585
R410 B.n750 B.n749 585
R411 B.n748 B.n2 585
R412 B.n693 B.n54 526.135
R413 B.n689 B.n55 526.135
R414 B.n565 B.n336 526.135
R415 B.n567 B.n334 526.135
R416 B.n104 B.t2 297.541
R417 B.n101 B.t10 297.541
R418 B.n480 B.t6 297.541
R419 B.n362 B.t13 297.541
R420 B.n691 B.n690 256.663
R421 B.n691 B.n99 256.663
R422 B.n691 B.n98 256.663
R423 B.n691 B.n97 256.663
R424 B.n691 B.n96 256.663
R425 B.n691 B.n95 256.663
R426 B.n691 B.n94 256.663
R427 B.n691 B.n93 256.663
R428 B.n691 B.n92 256.663
R429 B.n691 B.n91 256.663
R430 B.n691 B.n90 256.663
R431 B.n691 B.n89 256.663
R432 B.n691 B.n88 256.663
R433 B.n691 B.n87 256.663
R434 B.n691 B.n86 256.663
R435 B.n691 B.n85 256.663
R436 B.n691 B.n84 256.663
R437 B.n691 B.n83 256.663
R438 B.n691 B.n82 256.663
R439 B.n691 B.n81 256.663
R440 B.n691 B.n80 256.663
R441 B.n691 B.n79 256.663
R442 B.n691 B.n78 256.663
R443 B.n691 B.n77 256.663
R444 B.n691 B.n76 256.663
R445 B.n691 B.n75 256.663
R446 B.n691 B.n74 256.663
R447 B.n691 B.n73 256.663
R448 B.n691 B.n72 256.663
R449 B.n691 B.n71 256.663
R450 B.n691 B.n70 256.663
R451 B.n691 B.n69 256.663
R452 B.n691 B.n68 256.663
R453 B.n691 B.n67 256.663
R454 B.n691 B.n66 256.663
R455 B.n691 B.n65 256.663
R456 B.n691 B.n64 256.663
R457 B.n691 B.n63 256.663
R458 B.n691 B.n62 256.663
R459 B.n691 B.n61 256.663
R460 B.n691 B.n60 256.663
R461 B.n691 B.n59 256.663
R462 B.n691 B.n58 256.663
R463 B.n691 B.n57 256.663
R464 B.n691 B.n56 256.663
R465 B.n384 B.n335 256.663
R466 B.n387 B.n335 256.663
R467 B.n393 B.n335 256.663
R468 B.n395 B.n335 256.663
R469 B.n401 B.n335 256.663
R470 B.n403 B.n335 256.663
R471 B.n409 B.n335 256.663
R472 B.n411 B.n335 256.663
R473 B.n417 B.n335 256.663
R474 B.n419 B.n335 256.663
R475 B.n425 B.n335 256.663
R476 B.n427 B.n335 256.663
R477 B.n433 B.n335 256.663
R478 B.n435 B.n335 256.663
R479 B.n441 B.n335 256.663
R480 B.n443 B.n335 256.663
R481 B.n449 B.n335 256.663
R482 B.n451 B.n335 256.663
R483 B.n457 B.n335 256.663
R484 B.n459 B.n335 256.663
R485 B.n466 B.n335 256.663
R486 B.n468 B.n335 256.663
R487 B.n474 B.n335 256.663
R488 B.n476 B.n335 256.663
R489 B.n485 B.n335 256.663
R490 B.n487 B.n335 256.663
R491 B.n493 B.n335 256.663
R492 B.n495 B.n335 256.663
R493 B.n501 B.n335 256.663
R494 B.n503 B.n335 256.663
R495 B.n509 B.n335 256.663
R496 B.n511 B.n335 256.663
R497 B.n517 B.n335 256.663
R498 B.n519 B.n335 256.663
R499 B.n525 B.n335 256.663
R500 B.n527 B.n335 256.663
R501 B.n533 B.n335 256.663
R502 B.n535 B.n335 256.663
R503 B.n541 B.n335 256.663
R504 B.n543 B.n335 256.663
R505 B.n549 B.n335 256.663
R506 B.n551 B.n335 256.663
R507 B.n557 B.n335 256.663
R508 B.n560 B.n335 256.663
R509 B.n752 B.n751 256.663
R510 B.n109 B.n108 163.367
R511 B.n113 B.n112 163.367
R512 B.n117 B.n116 163.367
R513 B.n121 B.n120 163.367
R514 B.n125 B.n124 163.367
R515 B.n129 B.n128 163.367
R516 B.n133 B.n132 163.367
R517 B.n137 B.n136 163.367
R518 B.n141 B.n140 163.367
R519 B.n145 B.n144 163.367
R520 B.n149 B.n148 163.367
R521 B.n153 B.n152 163.367
R522 B.n157 B.n156 163.367
R523 B.n161 B.n160 163.367
R524 B.n165 B.n164 163.367
R525 B.n169 B.n168 163.367
R526 B.n173 B.n172 163.367
R527 B.n177 B.n176 163.367
R528 B.n181 B.n180 163.367
R529 B.n185 B.n184 163.367
R530 B.n189 B.n188 163.367
R531 B.n193 B.n192 163.367
R532 B.n197 B.n196 163.367
R533 B.n201 B.n200 163.367
R534 B.n205 B.n204 163.367
R535 B.n209 B.n208 163.367
R536 B.n213 B.n212 163.367
R537 B.n217 B.n216 163.367
R538 B.n221 B.n220 163.367
R539 B.n225 B.n224 163.367
R540 B.n229 B.n228 163.367
R541 B.n233 B.n232 163.367
R542 B.n237 B.n236 163.367
R543 B.n241 B.n240 163.367
R544 B.n245 B.n244 163.367
R545 B.n249 B.n248 163.367
R546 B.n253 B.n252 163.367
R547 B.n257 B.n256 163.367
R548 B.n261 B.n260 163.367
R549 B.n265 B.n264 163.367
R550 B.n269 B.n268 163.367
R551 B.n273 B.n272 163.367
R552 B.n277 B.n276 163.367
R553 B.n279 B.n100 163.367
R554 B.n565 B.n330 163.367
R555 B.n573 B.n330 163.367
R556 B.n573 B.n328 163.367
R557 B.n577 B.n328 163.367
R558 B.n577 B.n322 163.367
R559 B.n585 B.n322 163.367
R560 B.n585 B.n320 163.367
R561 B.n589 B.n320 163.367
R562 B.n589 B.n314 163.367
R563 B.n597 B.n314 163.367
R564 B.n597 B.n312 163.367
R565 B.n601 B.n312 163.367
R566 B.n601 B.n306 163.367
R567 B.n609 B.n306 163.367
R568 B.n609 B.n304 163.367
R569 B.n613 B.n304 163.367
R570 B.n613 B.n298 163.367
R571 B.n621 B.n298 163.367
R572 B.n621 B.n296 163.367
R573 B.n625 B.n296 163.367
R574 B.n625 B.n291 163.367
R575 B.n634 B.n291 163.367
R576 B.n634 B.n289 163.367
R577 B.n639 B.n289 163.367
R578 B.n639 B.n283 163.367
R579 B.n647 B.n283 163.367
R580 B.n648 B.n647 163.367
R581 B.n648 B.n5 163.367
R582 B.n6 B.n5 163.367
R583 B.n7 B.n6 163.367
R584 B.n654 B.n7 163.367
R585 B.n655 B.n654 163.367
R586 B.n655 B.n13 163.367
R587 B.n14 B.n13 163.367
R588 B.n15 B.n14 163.367
R589 B.n660 B.n15 163.367
R590 B.n660 B.n20 163.367
R591 B.n21 B.n20 163.367
R592 B.n22 B.n21 163.367
R593 B.n665 B.n22 163.367
R594 B.n665 B.n27 163.367
R595 B.n28 B.n27 163.367
R596 B.n29 B.n28 163.367
R597 B.n670 B.n29 163.367
R598 B.n670 B.n34 163.367
R599 B.n35 B.n34 163.367
R600 B.n36 B.n35 163.367
R601 B.n675 B.n36 163.367
R602 B.n675 B.n41 163.367
R603 B.n42 B.n41 163.367
R604 B.n43 B.n42 163.367
R605 B.n680 B.n43 163.367
R606 B.n680 B.n48 163.367
R607 B.n49 B.n48 163.367
R608 B.n50 B.n49 163.367
R609 B.n685 B.n50 163.367
R610 B.n685 B.n55 163.367
R611 B.n386 B.n385 163.367
R612 B.n388 B.n386 163.367
R613 B.n392 B.n381 163.367
R614 B.n396 B.n394 163.367
R615 B.n400 B.n379 163.367
R616 B.n404 B.n402 163.367
R617 B.n408 B.n377 163.367
R618 B.n412 B.n410 163.367
R619 B.n416 B.n375 163.367
R620 B.n420 B.n418 163.367
R621 B.n424 B.n373 163.367
R622 B.n428 B.n426 163.367
R623 B.n432 B.n371 163.367
R624 B.n436 B.n434 163.367
R625 B.n440 B.n369 163.367
R626 B.n444 B.n442 163.367
R627 B.n448 B.n367 163.367
R628 B.n452 B.n450 163.367
R629 B.n456 B.n365 163.367
R630 B.n460 B.n458 163.367
R631 B.n465 B.n361 163.367
R632 B.n469 B.n467 163.367
R633 B.n473 B.n359 163.367
R634 B.n477 B.n475 163.367
R635 B.n484 B.n357 163.367
R636 B.n488 B.n486 163.367
R637 B.n492 B.n355 163.367
R638 B.n496 B.n494 163.367
R639 B.n500 B.n353 163.367
R640 B.n504 B.n502 163.367
R641 B.n508 B.n351 163.367
R642 B.n512 B.n510 163.367
R643 B.n516 B.n349 163.367
R644 B.n520 B.n518 163.367
R645 B.n524 B.n347 163.367
R646 B.n528 B.n526 163.367
R647 B.n532 B.n345 163.367
R648 B.n536 B.n534 163.367
R649 B.n540 B.n343 163.367
R650 B.n544 B.n542 163.367
R651 B.n548 B.n341 163.367
R652 B.n552 B.n550 163.367
R653 B.n556 B.n339 163.367
R654 B.n559 B.n558 163.367
R655 B.n561 B.n336 163.367
R656 B.n567 B.n332 163.367
R657 B.n571 B.n332 163.367
R658 B.n571 B.n326 163.367
R659 B.n579 B.n326 163.367
R660 B.n579 B.n324 163.367
R661 B.n583 B.n324 163.367
R662 B.n583 B.n318 163.367
R663 B.n591 B.n318 163.367
R664 B.n591 B.n316 163.367
R665 B.n595 B.n316 163.367
R666 B.n595 B.n310 163.367
R667 B.n603 B.n310 163.367
R668 B.n603 B.n308 163.367
R669 B.n607 B.n308 163.367
R670 B.n607 B.n302 163.367
R671 B.n615 B.n302 163.367
R672 B.n615 B.n300 163.367
R673 B.n619 B.n300 163.367
R674 B.n619 B.n294 163.367
R675 B.n628 B.n294 163.367
R676 B.n628 B.n292 163.367
R677 B.n632 B.n292 163.367
R678 B.n632 B.n287 163.367
R679 B.n641 B.n287 163.367
R680 B.n641 B.n285 163.367
R681 B.n645 B.n285 163.367
R682 B.n645 B.n3 163.367
R683 B.n750 B.n3 163.367
R684 B.n746 B.n2 163.367
R685 B.n746 B.n745 163.367
R686 B.n745 B.n9 163.367
R687 B.n741 B.n9 163.367
R688 B.n741 B.n11 163.367
R689 B.n737 B.n11 163.367
R690 B.n737 B.n16 163.367
R691 B.n733 B.n16 163.367
R692 B.n733 B.n18 163.367
R693 B.n729 B.n18 163.367
R694 B.n729 B.n24 163.367
R695 B.n725 B.n24 163.367
R696 B.n725 B.n26 163.367
R697 B.n721 B.n26 163.367
R698 B.n721 B.n31 163.367
R699 B.n717 B.n31 163.367
R700 B.n717 B.n33 163.367
R701 B.n713 B.n33 163.367
R702 B.n713 B.n38 163.367
R703 B.n709 B.n38 163.367
R704 B.n709 B.n40 163.367
R705 B.n705 B.n40 163.367
R706 B.n705 B.n45 163.367
R707 B.n701 B.n45 163.367
R708 B.n701 B.n47 163.367
R709 B.n697 B.n47 163.367
R710 B.n697 B.n52 163.367
R711 B.n693 B.n52 163.367
R712 B.n101 B.t11 135.341
R713 B.n480 B.t9 135.341
R714 B.n104 B.t4 135.327
R715 B.n362 B.t15 135.327
R716 B.n566 B.n335 81.6271
R717 B.n692 B.n691 81.6271
R718 B.n56 B.n54 71.676
R719 B.n109 B.n57 71.676
R720 B.n113 B.n58 71.676
R721 B.n117 B.n59 71.676
R722 B.n121 B.n60 71.676
R723 B.n125 B.n61 71.676
R724 B.n129 B.n62 71.676
R725 B.n133 B.n63 71.676
R726 B.n137 B.n64 71.676
R727 B.n141 B.n65 71.676
R728 B.n145 B.n66 71.676
R729 B.n149 B.n67 71.676
R730 B.n153 B.n68 71.676
R731 B.n157 B.n69 71.676
R732 B.n161 B.n70 71.676
R733 B.n165 B.n71 71.676
R734 B.n169 B.n72 71.676
R735 B.n173 B.n73 71.676
R736 B.n177 B.n74 71.676
R737 B.n181 B.n75 71.676
R738 B.n185 B.n76 71.676
R739 B.n189 B.n77 71.676
R740 B.n193 B.n78 71.676
R741 B.n197 B.n79 71.676
R742 B.n201 B.n80 71.676
R743 B.n205 B.n81 71.676
R744 B.n209 B.n82 71.676
R745 B.n213 B.n83 71.676
R746 B.n217 B.n84 71.676
R747 B.n221 B.n85 71.676
R748 B.n225 B.n86 71.676
R749 B.n229 B.n87 71.676
R750 B.n233 B.n88 71.676
R751 B.n237 B.n89 71.676
R752 B.n241 B.n90 71.676
R753 B.n245 B.n91 71.676
R754 B.n249 B.n92 71.676
R755 B.n253 B.n93 71.676
R756 B.n257 B.n94 71.676
R757 B.n261 B.n95 71.676
R758 B.n265 B.n96 71.676
R759 B.n269 B.n97 71.676
R760 B.n273 B.n98 71.676
R761 B.n277 B.n99 71.676
R762 B.n690 B.n100 71.676
R763 B.n690 B.n689 71.676
R764 B.n279 B.n99 71.676
R765 B.n276 B.n98 71.676
R766 B.n272 B.n97 71.676
R767 B.n268 B.n96 71.676
R768 B.n264 B.n95 71.676
R769 B.n260 B.n94 71.676
R770 B.n256 B.n93 71.676
R771 B.n252 B.n92 71.676
R772 B.n248 B.n91 71.676
R773 B.n244 B.n90 71.676
R774 B.n240 B.n89 71.676
R775 B.n236 B.n88 71.676
R776 B.n232 B.n87 71.676
R777 B.n228 B.n86 71.676
R778 B.n224 B.n85 71.676
R779 B.n220 B.n84 71.676
R780 B.n216 B.n83 71.676
R781 B.n212 B.n82 71.676
R782 B.n208 B.n81 71.676
R783 B.n204 B.n80 71.676
R784 B.n200 B.n79 71.676
R785 B.n196 B.n78 71.676
R786 B.n192 B.n77 71.676
R787 B.n188 B.n76 71.676
R788 B.n184 B.n75 71.676
R789 B.n180 B.n74 71.676
R790 B.n176 B.n73 71.676
R791 B.n172 B.n72 71.676
R792 B.n168 B.n71 71.676
R793 B.n164 B.n70 71.676
R794 B.n160 B.n69 71.676
R795 B.n156 B.n68 71.676
R796 B.n152 B.n67 71.676
R797 B.n148 B.n66 71.676
R798 B.n144 B.n65 71.676
R799 B.n140 B.n64 71.676
R800 B.n136 B.n63 71.676
R801 B.n132 B.n62 71.676
R802 B.n128 B.n61 71.676
R803 B.n124 B.n60 71.676
R804 B.n120 B.n59 71.676
R805 B.n116 B.n58 71.676
R806 B.n112 B.n57 71.676
R807 B.n108 B.n56 71.676
R808 B.n384 B.n334 71.676
R809 B.n388 B.n387 71.676
R810 B.n393 B.n392 71.676
R811 B.n396 B.n395 71.676
R812 B.n401 B.n400 71.676
R813 B.n404 B.n403 71.676
R814 B.n409 B.n408 71.676
R815 B.n412 B.n411 71.676
R816 B.n417 B.n416 71.676
R817 B.n420 B.n419 71.676
R818 B.n425 B.n424 71.676
R819 B.n428 B.n427 71.676
R820 B.n433 B.n432 71.676
R821 B.n436 B.n435 71.676
R822 B.n441 B.n440 71.676
R823 B.n444 B.n443 71.676
R824 B.n449 B.n448 71.676
R825 B.n452 B.n451 71.676
R826 B.n457 B.n456 71.676
R827 B.n460 B.n459 71.676
R828 B.n466 B.n465 71.676
R829 B.n469 B.n468 71.676
R830 B.n474 B.n473 71.676
R831 B.n477 B.n476 71.676
R832 B.n485 B.n484 71.676
R833 B.n488 B.n487 71.676
R834 B.n493 B.n492 71.676
R835 B.n496 B.n495 71.676
R836 B.n501 B.n500 71.676
R837 B.n504 B.n503 71.676
R838 B.n509 B.n508 71.676
R839 B.n512 B.n511 71.676
R840 B.n517 B.n516 71.676
R841 B.n520 B.n519 71.676
R842 B.n525 B.n524 71.676
R843 B.n528 B.n527 71.676
R844 B.n533 B.n532 71.676
R845 B.n536 B.n535 71.676
R846 B.n541 B.n540 71.676
R847 B.n544 B.n543 71.676
R848 B.n549 B.n548 71.676
R849 B.n552 B.n551 71.676
R850 B.n557 B.n556 71.676
R851 B.n560 B.n559 71.676
R852 B.n385 B.n384 71.676
R853 B.n387 B.n381 71.676
R854 B.n394 B.n393 71.676
R855 B.n395 B.n379 71.676
R856 B.n402 B.n401 71.676
R857 B.n403 B.n377 71.676
R858 B.n410 B.n409 71.676
R859 B.n411 B.n375 71.676
R860 B.n418 B.n417 71.676
R861 B.n419 B.n373 71.676
R862 B.n426 B.n425 71.676
R863 B.n427 B.n371 71.676
R864 B.n434 B.n433 71.676
R865 B.n435 B.n369 71.676
R866 B.n442 B.n441 71.676
R867 B.n443 B.n367 71.676
R868 B.n450 B.n449 71.676
R869 B.n451 B.n365 71.676
R870 B.n458 B.n457 71.676
R871 B.n459 B.n361 71.676
R872 B.n467 B.n466 71.676
R873 B.n468 B.n359 71.676
R874 B.n475 B.n474 71.676
R875 B.n476 B.n357 71.676
R876 B.n486 B.n485 71.676
R877 B.n487 B.n355 71.676
R878 B.n494 B.n493 71.676
R879 B.n495 B.n353 71.676
R880 B.n502 B.n501 71.676
R881 B.n503 B.n351 71.676
R882 B.n510 B.n509 71.676
R883 B.n511 B.n349 71.676
R884 B.n518 B.n517 71.676
R885 B.n519 B.n347 71.676
R886 B.n526 B.n525 71.676
R887 B.n527 B.n345 71.676
R888 B.n534 B.n533 71.676
R889 B.n535 B.n343 71.676
R890 B.n542 B.n541 71.676
R891 B.n543 B.n341 71.676
R892 B.n550 B.n549 71.676
R893 B.n551 B.n339 71.676
R894 B.n558 B.n557 71.676
R895 B.n561 B.n560 71.676
R896 B.n751 B.n750 71.676
R897 B.n751 B.n2 71.676
R898 B.n102 B.t12 68.0447
R899 B.n481 B.t8 68.0447
R900 B.n105 B.t5 68.0299
R901 B.n363 B.t14 68.0299
R902 B.n105 B.n104 67.2975
R903 B.n102 B.n101 67.2975
R904 B.n481 B.n480 67.2975
R905 B.n363 B.n362 67.2975
R906 B.n106 B.n105 59.5399
R907 B.n103 B.n102 59.5399
R908 B.n482 B.n481 59.5399
R909 B.n462 B.n363 59.5399
R910 B.n566 B.n331 44.4054
R911 B.n572 B.n331 44.4054
R912 B.n572 B.n327 44.4054
R913 B.n578 B.n327 44.4054
R914 B.n578 B.n323 44.4054
R915 B.n584 B.n323 44.4054
R916 B.n584 B.n319 44.4054
R917 B.n590 B.n319 44.4054
R918 B.n596 B.n315 44.4054
R919 B.n596 B.n311 44.4054
R920 B.n602 B.n311 44.4054
R921 B.n602 B.n307 44.4054
R922 B.n608 B.n307 44.4054
R923 B.n608 B.n303 44.4054
R924 B.n614 B.n303 44.4054
R925 B.n614 B.n299 44.4054
R926 B.n620 B.n299 44.4054
R927 B.n620 B.n295 44.4054
R928 B.n627 B.n295 44.4054
R929 B.n627 B.n626 44.4054
R930 B.n633 B.n288 44.4054
R931 B.n640 B.n288 44.4054
R932 B.n640 B.n284 44.4054
R933 B.n646 B.n284 44.4054
R934 B.n646 B.n4 44.4054
R935 B.n749 B.n4 44.4054
R936 B.n749 B.n748 44.4054
R937 B.n748 B.n747 44.4054
R938 B.n747 B.n8 44.4054
R939 B.n12 B.n8 44.4054
R940 B.n740 B.n12 44.4054
R941 B.n740 B.n739 44.4054
R942 B.n739 B.n738 44.4054
R943 B.n732 B.n19 44.4054
R944 B.n732 B.n731 44.4054
R945 B.n731 B.n730 44.4054
R946 B.n730 B.n23 44.4054
R947 B.n724 B.n23 44.4054
R948 B.n724 B.n723 44.4054
R949 B.n723 B.n722 44.4054
R950 B.n722 B.n30 44.4054
R951 B.n716 B.n30 44.4054
R952 B.n716 B.n715 44.4054
R953 B.n715 B.n714 44.4054
R954 B.n714 B.n37 44.4054
R955 B.n708 B.n707 44.4054
R956 B.n707 B.n706 44.4054
R957 B.n706 B.n44 44.4054
R958 B.n700 B.n44 44.4054
R959 B.n700 B.n699 44.4054
R960 B.n699 B.n698 44.4054
R961 B.n698 B.n51 44.4054
R962 B.n692 B.n51 44.4054
R963 B.n626 B.t0 35.2632
R964 B.n19 B.t1 35.2632
R965 B.n568 B.n333 34.1859
R966 B.n564 B.n563 34.1859
R967 B.n688 B.n687 34.1859
R968 B.n694 B.n53 34.1859
R969 B.t7 B.n315 27.427
R970 B.t3 B.n37 27.427
R971 B B.n752 18.0485
R972 B.n590 B.t7 16.9788
R973 B.n708 B.t3 16.9788
R974 B.n569 B.n568 10.6151
R975 B.n570 B.n569 10.6151
R976 B.n570 B.n325 10.6151
R977 B.n580 B.n325 10.6151
R978 B.n581 B.n580 10.6151
R979 B.n582 B.n581 10.6151
R980 B.n582 B.n317 10.6151
R981 B.n592 B.n317 10.6151
R982 B.n593 B.n592 10.6151
R983 B.n594 B.n593 10.6151
R984 B.n594 B.n309 10.6151
R985 B.n604 B.n309 10.6151
R986 B.n605 B.n604 10.6151
R987 B.n606 B.n605 10.6151
R988 B.n606 B.n301 10.6151
R989 B.n616 B.n301 10.6151
R990 B.n617 B.n616 10.6151
R991 B.n618 B.n617 10.6151
R992 B.n618 B.n293 10.6151
R993 B.n629 B.n293 10.6151
R994 B.n630 B.n629 10.6151
R995 B.n631 B.n630 10.6151
R996 B.n631 B.n286 10.6151
R997 B.n642 B.n286 10.6151
R998 B.n643 B.n642 10.6151
R999 B.n644 B.n643 10.6151
R1000 B.n644 B.n0 10.6151
R1001 B.n383 B.n333 10.6151
R1002 B.n383 B.n382 10.6151
R1003 B.n389 B.n382 10.6151
R1004 B.n390 B.n389 10.6151
R1005 B.n391 B.n390 10.6151
R1006 B.n391 B.n380 10.6151
R1007 B.n397 B.n380 10.6151
R1008 B.n398 B.n397 10.6151
R1009 B.n399 B.n398 10.6151
R1010 B.n399 B.n378 10.6151
R1011 B.n405 B.n378 10.6151
R1012 B.n406 B.n405 10.6151
R1013 B.n407 B.n406 10.6151
R1014 B.n407 B.n376 10.6151
R1015 B.n413 B.n376 10.6151
R1016 B.n414 B.n413 10.6151
R1017 B.n415 B.n414 10.6151
R1018 B.n415 B.n374 10.6151
R1019 B.n421 B.n374 10.6151
R1020 B.n422 B.n421 10.6151
R1021 B.n423 B.n422 10.6151
R1022 B.n423 B.n372 10.6151
R1023 B.n429 B.n372 10.6151
R1024 B.n430 B.n429 10.6151
R1025 B.n431 B.n430 10.6151
R1026 B.n431 B.n370 10.6151
R1027 B.n437 B.n370 10.6151
R1028 B.n438 B.n437 10.6151
R1029 B.n439 B.n438 10.6151
R1030 B.n439 B.n368 10.6151
R1031 B.n445 B.n368 10.6151
R1032 B.n446 B.n445 10.6151
R1033 B.n447 B.n446 10.6151
R1034 B.n447 B.n366 10.6151
R1035 B.n453 B.n366 10.6151
R1036 B.n454 B.n453 10.6151
R1037 B.n455 B.n454 10.6151
R1038 B.n455 B.n364 10.6151
R1039 B.n461 B.n364 10.6151
R1040 B.n464 B.n463 10.6151
R1041 B.n464 B.n360 10.6151
R1042 B.n470 B.n360 10.6151
R1043 B.n471 B.n470 10.6151
R1044 B.n472 B.n471 10.6151
R1045 B.n472 B.n358 10.6151
R1046 B.n478 B.n358 10.6151
R1047 B.n479 B.n478 10.6151
R1048 B.n483 B.n479 10.6151
R1049 B.n489 B.n356 10.6151
R1050 B.n490 B.n489 10.6151
R1051 B.n491 B.n490 10.6151
R1052 B.n491 B.n354 10.6151
R1053 B.n497 B.n354 10.6151
R1054 B.n498 B.n497 10.6151
R1055 B.n499 B.n498 10.6151
R1056 B.n499 B.n352 10.6151
R1057 B.n505 B.n352 10.6151
R1058 B.n506 B.n505 10.6151
R1059 B.n507 B.n506 10.6151
R1060 B.n507 B.n350 10.6151
R1061 B.n513 B.n350 10.6151
R1062 B.n514 B.n513 10.6151
R1063 B.n515 B.n514 10.6151
R1064 B.n515 B.n348 10.6151
R1065 B.n521 B.n348 10.6151
R1066 B.n522 B.n521 10.6151
R1067 B.n523 B.n522 10.6151
R1068 B.n523 B.n346 10.6151
R1069 B.n529 B.n346 10.6151
R1070 B.n530 B.n529 10.6151
R1071 B.n531 B.n530 10.6151
R1072 B.n531 B.n344 10.6151
R1073 B.n537 B.n344 10.6151
R1074 B.n538 B.n537 10.6151
R1075 B.n539 B.n538 10.6151
R1076 B.n539 B.n342 10.6151
R1077 B.n545 B.n342 10.6151
R1078 B.n546 B.n545 10.6151
R1079 B.n547 B.n546 10.6151
R1080 B.n547 B.n340 10.6151
R1081 B.n553 B.n340 10.6151
R1082 B.n554 B.n553 10.6151
R1083 B.n555 B.n554 10.6151
R1084 B.n555 B.n338 10.6151
R1085 B.n338 B.n337 10.6151
R1086 B.n562 B.n337 10.6151
R1087 B.n563 B.n562 10.6151
R1088 B.n564 B.n329 10.6151
R1089 B.n574 B.n329 10.6151
R1090 B.n575 B.n574 10.6151
R1091 B.n576 B.n575 10.6151
R1092 B.n576 B.n321 10.6151
R1093 B.n586 B.n321 10.6151
R1094 B.n587 B.n586 10.6151
R1095 B.n588 B.n587 10.6151
R1096 B.n588 B.n313 10.6151
R1097 B.n598 B.n313 10.6151
R1098 B.n599 B.n598 10.6151
R1099 B.n600 B.n599 10.6151
R1100 B.n600 B.n305 10.6151
R1101 B.n610 B.n305 10.6151
R1102 B.n611 B.n610 10.6151
R1103 B.n612 B.n611 10.6151
R1104 B.n612 B.n297 10.6151
R1105 B.n622 B.n297 10.6151
R1106 B.n623 B.n622 10.6151
R1107 B.n624 B.n623 10.6151
R1108 B.n624 B.n290 10.6151
R1109 B.n635 B.n290 10.6151
R1110 B.n636 B.n635 10.6151
R1111 B.n638 B.n636 10.6151
R1112 B.n638 B.n637 10.6151
R1113 B.n637 B.n282 10.6151
R1114 B.n649 B.n282 10.6151
R1115 B.n650 B.n649 10.6151
R1116 B.n651 B.n650 10.6151
R1117 B.n652 B.n651 10.6151
R1118 B.n653 B.n652 10.6151
R1119 B.n656 B.n653 10.6151
R1120 B.n657 B.n656 10.6151
R1121 B.n658 B.n657 10.6151
R1122 B.n659 B.n658 10.6151
R1123 B.n661 B.n659 10.6151
R1124 B.n662 B.n661 10.6151
R1125 B.n663 B.n662 10.6151
R1126 B.n664 B.n663 10.6151
R1127 B.n666 B.n664 10.6151
R1128 B.n667 B.n666 10.6151
R1129 B.n668 B.n667 10.6151
R1130 B.n669 B.n668 10.6151
R1131 B.n671 B.n669 10.6151
R1132 B.n672 B.n671 10.6151
R1133 B.n673 B.n672 10.6151
R1134 B.n674 B.n673 10.6151
R1135 B.n676 B.n674 10.6151
R1136 B.n677 B.n676 10.6151
R1137 B.n678 B.n677 10.6151
R1138 B.n679 B.n678 10.6151
R1139 B.n681 B.n679 10.6151
R1140 B.n682 B.n681 10.6151
R1141 B.n683 B.n682 10.6151
R1142 B.n684 B.n683 10.6151
R1143 B.n686 B.n684 10.6151
R1144 B.n687 B.n686 10.6151
R1145 B.n744 B.n1 10.6151
R1146 B.n744 B.n743 10.6151
R1147 B.n743 B.n742 10.6151
R1148 B.n742 B.n10 10.6151
R1149 B.n736 B.n10 10.6151
R1150 B.n736 B.n735 10.6151
R1151 B.n735 B.n734 10.6151
R1152 B.n734 B.n17 10.6151
R1153 B.n728 B.n17 10.6151
R1154 B.n728 B.n727 10.6151
R1155 B.n727 B.n726 10.6151
R1156 B.n726 B.n25 10.6151
R1157 B.n720 B.n25 10.6151
R1158 B.n720 B.n719 10.6151
R1159 B.n719 B.n718 10.6151
R1160 B.n718 B.n32 10.6151
R1161 B.n712 B.n32 10.6151
R1162 B.n712 B.n711 10.6151
R1163 B.n711 B.n710 10.6151
R1164 B.n710 B.n39 10.6151
R1165 B.n704 B.n39 10.6151
R1166 B.n704 B.n703 10.6151
R1167 B.n703 B.n702 10.6151
R1168 B.n702 B.n46 10.6151
R1169 B.n696 B.n46 10.6151
R1170 B.n696 B.n695 10.6151
R1171 B.n695 B.n694 10.6151
R1172 B.n107 B.n53 10.6151
R1173 B.n110 B.n107 10.6151
R1174 B.n111 B.n110 10.6151
R1175 B.n114 B.n111 10.6151
R1176 B.n115 B.n114 10.6151
R1177 B.n118 B.n115 10.6151
R1178 B.n119 B.n118 10.6151
R1179 B.n122 B.n119 10.6151
R1180 B.n123 B.n122 10.6151
R1181 B.n126 B.n123 10.6151
R1182 B.n127 B.n126 10.6151
R1183 B.n130 B.n127 10.6151
R1184 B.n131 B.n130 10.6151
R1185 B.n134 B.n131 10.6151
R1186 B.n135 B.n134 10.6151
R1187 B.n138 B.n135 10.6151
R1188 B.n139 B.n138 10.6151
R1189 B.n142 B.n139 10.6151
R1190 B.n143 B.n142 10.6151
R1191 B.n146 B.n143 10.6151
R1192 B.n147 B.n146 10.6151
R1193 B.n150 B.n147 10.6151
R1194 B.n151 B.n150 10.6151
R1195 B.n154 B.n151 10.6151
R1196 B.n155 B.n154 10.6151
R1197 B.n158 B.n155 10.6151
R1198 B.n159 B.n158 10.6151
R1199 B.n162 B.n159 10.6151
R1200 B.n163 B.n162 10.6151
R1201 B.n166 B.n163 10.6151
R1202 B.n167 B.n166 10.6151
R1203 B.n170 B.n167 10.6151
R1204 B.n171 B.n170 10.6151
R1205 B.n174 B.n171 10.6151
R1206 B.n175 B.n174 10.6151
R1207 B.n178 B.n175 10.6151
R1208 B.n179 B.n178 10.6151
R1209 B.n182 B.n179 10.6151
R1210 B.n183 B.n182 10.6151
R1211 B.n187 B.n186 10.6151
R1212 B.n190 B.n187 10.6151
R1213 B.n191 B.n190 10.6151
R1214 B.n194 B.n191 10.6151
R1215 B.n195 B.n194 10.6151
R1216 B.n198 B.n195 10.6151
R1217 B.n199 B.n198 10.6151
R1218 B.n202 B.n199 10.6151
R1219 B.n203 B.n202 10.6151
R1220 B.n207 B.n206 10.6151
R1221 B.n210 B.n207 10.6151
R1222 B.n211 B.n210 10.6151
R1223 B.n214 B.n211 10.6151
R1224 B.n215 B.n214 10.6151
R1225 B.n218 B.n215 10.6151
R1226 B.n219 B.n218 10.6151
R1227 B.n222 B.n219 10.6151
R1228 B.n223 B.n222 10.6151
R1229 B.n226 B.n223 10.6151
R1230 B.n227 B.n226 10.6151
R1231 B.n230 B.n227 10.6151
R1232 B.n231 B.n230 10.6151
R1233 B.n234 B.n231 10.6151
R1234 B.n235 B.n234 10.6151
R1235 B.n238 B.n235 10.6151
R1236 B.n239 B.n238 10.6151
R1237 B.n242 B.n239 10.6151
R1238 B.n243 B.n242 10.6151
R1239 B.n246 B.n243 10.6151
R1240 B.n247 B.n246 10.6151
R1241 B.n250 B.n247 10.6151
R1242 B.n251 B.n250 10.6151
R1243 B.n254 B.n251 10.6151
R1244 B.n255 B.n254 10.6151
R1245 B.n258 B.n255 10.6151
R1246 B.n259 B.n258 10.6151
R1247 B.n262 B.n259 10.6151
R1248 B.n263 B.n262 10.6151
R1249 B.n266 B.n263 10.6151
R1250 B.n267 B.n266 10.6151
R1251 B.n270 B.n267 10.6151
R1252 B.n271 B.n270 10.6151
R1253 B.n274 B.n271 10.6151
R1254 B.n275 B.n274 10.6151
R1255 B.n278 B.n275 10.6151
R1256 B.n280 B.n278 10.6151
R1257 B.n281 B.n280 10.6151
R1258 B.n688 B.n281 10.6151
R1259 B.n462 B.n461 9.36635
R1260 B.n482 B.n356 9.36635
R1261 B.n183 B.n106 9.36635
R1262 B.n206 B.n103 9.36635
R1263 B.n633 B.t0 9.14268
R1264 B.n738 B.t1 9.14268
R1265 B.n752 B.n0 8.11757
R1266 B.n752 B.n1 8.11757
R1267 B.n463 B.n462 1.24928
R1268 B.n483 B.n482 1.24928
R1269 B.n186 B.n106 1.24928
R1270 B.n203 B.n103 1.24928
R1271 VN VN.t1 173.26
R1272 VN VN.t0 128.115
R1273 VTAIL.n1 VTAIL.t2 49.6605
R1274 VTAIL.n3 VTAIL.t3 49.6596
R1275 VTAIL.n0 VTAIL.t1 49.6596
R1276 VTAIL.n2 VTAIL.t0 49.6594
R1277 VTAIL.n1 VTAIL.n0 28.3238
R1278 VTAIL.n3 VTAIL.n2 25.3324
R1279 VTAIL.n2 VTAIL.n1 1.96602
R1280 VTAIL VTAIL.n0 1.27636
R1281 VTAIL VTAIL.n3 0.690155
R1282 VDD2.n0 VDD2.t1 105.954
R1283 VDD2.n0 VDD2.t0 66.3382
R1284 VDD2 VDD2.n0 0.806535
R1285 VP.n0 VP.t1 173.352
R1286 VP.n0 VP.t0 127.59
R1287 VP VP.n0 0.52637
R1288 VDD1 VDD1.t1 107.228
R1289 VDD1 VDD1.t0 67.1442
C0 VDD2 VP 0.355717f
C1 VDD2 VTAIL 5.10548f
C2 VDD1 VDD2 0.740235f
C3 VDD2 VN 2.76166f
C4 VTAIL VP 2.50011f
C5 VDD1 VP 2.96677f
C6 VP VN 5.63392f
C7 VDD1 VTAIL 5.05066f
C8 VTAIL VN 2.48587f
C9 VDD1 VN 0.14837f
C10 VDD2 B 4.54265f
C11 VDD1 B 7.7816f
C12 VTAIL B 7.449738f
C13 VN B 11.181231f
C14 VP B 7.056954f
C15 VDD1.t0 B 2.168f
C16 VDD1.t1 B 2.75903f
C17 VP.t1 B 3.79098f
C18 VP.t0 B 3.16405f
C19 VP.n0 B 4.05119f
C20 VDD2.t1 B 2.67752f
C21 VDD2.t0 B 2.13143f
C22 VDD2.n0 B 2.93864f
C23 VTAIL.t1 B 2.13007f
C24 VTAIL.n0 B 1.72488f
C25 VTAIL.t2 B 2.13007f
C26 VTAIL.n1 B 1.77189f
C27 VTAIL.t0 B 2.13006f
C28 VTAIL.n2 B 1.56799f
C29 VTAIL.t3 B 2.13007f
C30 VTAIL.n3 B 1.48101f
C31 VN.t0 B 3.09999f
C32 VN.t1 B 3.70943f
.ends

