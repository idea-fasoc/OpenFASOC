* NGSPICE file created from diff_pair_sample_0131.ext - technology: sky130A

.subckt diff_pair_sample_0131 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t9 w_n3914_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=7.0083 ps=36.72 w=17.97 l=3.35
X1 VTAIL.t6 VP.t1 VDD1.t4 w_n3914_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=2.96505 ps=18.3 w=17.97 l=3.35
X2 VDD2.t5 VN.t0 VTAIL.t1 w_n3914_n4562# sky130_fd_pr__pfet_01v8 ad=7.0083 pd=36.72 as=2.96505 ps=18.3 w=17.97 l=3.35
X3 VTAIL.t3 VN.t1 VDD2.t4 w_n3914_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=2.96505 ps=18.3 w=17.97 l=3.35
X4 B.t11 B.t9 B.t10 w_n3914_n4562# sky130_fd_pr__pfet_01v8 ad=7.0083 pd=36.72 as=0 ps=0 w=17.97 l=3.35
X5 VDD2.t3 VN.t2 VTAIL.t5 w_n3914_n4562# sky130_fd_pr__pfet_01v8 ad=7.0083 pd=36.72 as=2.96505 ps=18.3 w=17.97 l=3.35
X6 VDD2.t2 VN.t3 VTAIL.t0 w_n3914_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=7.0083 ps=36.72 w=17.97 l=3.35
X7 VDD1.t3 VP.t2 VTAIL.t10 w_n3914_n4562# sky130_fd_pr__pfet_01v8 ad=7.0083 pd=36.72 as=2.96505 ps=18.3 w=17.97 l=3.35
X8 VTAIL.t2 VN.t4 VDD2.t1 w_n3914_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=2.96505 ps=18.3 w=17.97 l=3.35
X9 B.t8 B.t6 B.t7 w_n3914_n4562# sky130_fd_pr__pfet_01v8 ad=7.0083 pd=36.72 as=0 ps=0 w=17.97 l=3.35
X10 B.t5 B.t3 B.t4 w_n3914_n4562# sky130_fd_pr__pfet_01v8 ad=7.0083 pd=36.72 as=0 ps=0 w=17.97 l=3.35
X11 VDD2.t0 VN.t5 VTAIL.t4 w_n3914_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=7.0083 ps=36.72 w=17.97 l=3.35
X12 B.t2 B.t0 B.t1 w_n3914_n4562# sky130_fd_pr__pfet_01v8 ad=7.0083 pd=36.72 as=0 ps=0 w=17.97 l=3.35
X13 VTAIL.t8 VP.t3 VDD1.t2 w_n3914_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=2.96505 ps=18.3 w=17.97 l=3.35
X14 VDD1.t1 VP.t4 VTAIL.t11 w_n3914_n4562# sky130_fd_pr__pfet_01v8 ad=7.0083 pd=36.72 as=2.96505 ps=18.3 w=17.97 l=3.35
X15 VDD1.t0 VP.t5 VTAIL.t7 w_n3914_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=7.0083 ps=36.72 w=17.97 l=3.35
R0 VP.n14 VP.t4 162.486
R1 VP.n16 VP.n15 161.3
R2 VP.n17 VP.n12 161.3
R3 VP.n19 VP.n18 161.3
R4 VP.n20 VP.n11 161.3
R5 VP.n22 VP.n21 161.3
R6 VP.n23 VP.n10 161.3
R7 VP.n25 VP.n24 161.3
R8 VP.n50 VP.n49 161.3
R9 VP.n48 VP.n1 161.3
R10 VP.n47 VP.n46 161.3
R11 VP.n45 VP.n2 161.3
R12 VP.n44 VP.n43 161.3
R13 VP.n42 VP.n3 161.3
R14 VP.n41 VP.n40 161.3
R15 VP.n39 VP.n4 161.3
R16 VP.n38 VP.n37 161.3
R17 VP.n36 VP.n5 161.3
R18 VP.n35 VP.n34 161.3
R19 VP.n33 VP.n6 161.3
R20 VP.n32 VP.n31 161.3
R21 VP.n30 VP.n7 161.3
R22 VP.n29 VP.n28 161.3
R23 VP.n4 VP.t3 129.278
R24 VP.n8 VP.t2 129.278
R25 VP.n0 VP.t5 129.278
R26 VP.n13 VP.t1 129.278
R27 VP.n9 VP.t0 129.278
R28 VP.n27 VP.n8 81.2593
R29 VP.n51 VP.n0 81.2593
R30 VP.n26 VP.n9 81.2593
R31 VP.n27 VP.n26 56.1736
R32 VP.n35 VP.n6 56.0336
R33 VP.n43 VP.n2 56.0336
R34 VP.n18 VP.n11 56.0336
R35 VP.n14 VP.n13 50.0921
R36 VP.n31 VP.n6 24.9531
R37 VP.n47 VP.n2 24.9531
R38 VP.n22 VP.n11 24.9531
R39 VP.n30 VP.n29 24.4675
R40 VP.n31 VP.n30 24.4675
R41 VP.n36 VP.n35 24.4675
R42 VP.n37 VP.n36 24.4675
R43 VP.n37 VP.n4 24.4675
R44 VP.n41 VP.n4 24.4675
R45 VP.n42 VP.n41 24.4675
R46 VP.n43 VP.n42 24.4675
R47 VP.n48 VP.n47 24.4675
R48 VP.n49 VP.n48 24.4675
R49 VP.n23 VP.n22 24.4675
R50 VP.n24 VP.n23 24.4675
R51 VP.n16 VP.n13 24.4675
R52 VP.n17 VP.n16 24.4675
R53 VP.n18 VP.n17 24.4675
R54 VP.n29 VP.n8 8.80862
R55 VP.n49 VP.n0 8.80862
R56 VP.n24 VP.n9 8.80862
R57 VP.n15 VP.n14 3.19478
R58 VP.n26 VP.n25 0.354971
R59 VP.n28 VP.n27 0.354971
R60 VP.n51 VP.n50 0.354971
R61 VP VP.n51 0.26696
R62 VP.n15 VP.n12 0.189894
R63 VP.n19 VP.n12 0.189894
R64 VP.n20 VP.n19 0.189894
R65 VP.n21 VP.n20 0.189894
R66 VP.n21 VP.n10 0.189894
R67 VP.n25 VP.n10 0.189894
R68 VP.n28 VP.n7 0.189894
R69 VP.n32 VP.n7 0.189894
R70 VP.n33 VP.n32 0.189894
R71 VP.n34 VP.n33 0.189894
R72 VP.n34 VP.n5 0.189894
R73 VP.n38 VP.n5 0.189894
R74 VP.n39 VP.n38 0.189894
R75 VP.n40 VP.n39 0.189894
R76 VP.n40 VP.n3 0.189894
R77 VP.n44 VP.n3 0.189894
R78 VP.n45 VP.n44 0.189894
R79 VP.n46 VP.n45 0.189894
R80 VP.n46 VP.n1 0.189894
R81 VP.n50 VP.n1 0.189894
R82 VTAIL.n7 VTAIL.t0 55.7262
R83 VTAIL.n11 VTAIL.t4 55.726
R84 VTAIL.n2 VTAIL.t7 55.726
R85 VTAIL.n10 VTAIL.t9 55.726
R86 VTAIL.n9 VTAIL.n8 53.9174
R87 VTAIL.n6 VTAIL.n5 53.9174
R88 VTAIL.n1 VTAIL.n0 53.9171
R89 VTAIL.n4 VTAIL.n3 53.9171
R90 VTAIL.n6 VTAIL.n4 34.2031
R91 VTAIL.n11 VTAIL.n10 31.0307
R92 VTAIL.n7 VTAIL.n6 3.17291
R93 VTAIL.n10 VTAIL.n9 3.17291
R94 VTAIL.n4 VTAIL.n2 3.17291
R95 VTAIL VTAIL.n11 2.32162
R96 VTAIL.n9 VTAIL.n7 2.05653
R97 VTAIL.n2 VTAIL.n1 2.05653
R98 VTAIL.n0 VTAIL.t5 1.80935
R99 VTAIL.n0 VTAIL.t3 1.80935
R100 VTAIL.n3 VTAIL.t10 1.80935
R101 VTAIL.n3 VTAIL.t8 1.80935
R102 VTAIL.n8 VTAIL.t11 1.80935
R103 VTAIL.n8 VTAIL.t6 1.80935
R104 VTAIL.n5 VTAIL.t1 1.80935
R105 VTAIL.n5 VTAIL.t2 1.80935
R106 VTAIL VTAIL.n1 0.851793
R107 VDD1 VDD1.t1 74.8425
R108 VDD1.n1 VDD1.t3 74.7287
R109 VDD1.n1 VDD1.n0 71.3336
R110 VDD1.n3 VDD1.n2 70.596
R111 VDD1.n3 VDD1.n1 51.6862
R112 VDD1.n2 VDD1.t4 1.80935
R113 VDD1.n2 VDD1.t5 1.80935
R114 VDD1.n0 VDD1.t2 1.80935
R115 VDD1.n0 VDD1.t0 1.80935
R116 VDD1 VDD1.n3 0.735414
R117 VN.n23 VN.t3 162.486
R118 VN.n5 VN.t2 162.486
R119 VN.n34 VN.n33 161.3
R120 VN.n32 VN.n19 161.3
R121 VN.n31 VN.n30 161.3
R122 VN.n29 VN.n20 161.3
R123 VN.n28 VN.n27 161.3
R124 VN.n26 VN.n21 161.3
R125 VN.n25 VN.n24 161.3
R126 VN.n16 VN.n15 161.3
R127 VN.n14 VN.n1 161.3
R128 VN.n13 VN.n12 161.3
R129 VN.n11 VN.n2 161.3
R130 VN.n10 VN.n9 161.3
R131 VN.n8 VN.n3 161.3
R132 VN.n7 VN.n6 161.3
R133 VN.n4 VN.t1 129.278
R134 VN.n0 VN.t5 129.278
R135 VN.n22 VN.t4 129.278
R136 VN.n18 VN.t0 129.278
R137 VN.n17 VN.n0 81.2593
R138 VN.n35 VN.n18 81.2593
R139 VN VN.n35 56.3389
R140 VN.n9 VN.n2 56.0336
R141 VN.n27 VN.n20 56.0336
R142 VN.n5 VN.n4 50.0921
R143 VN.n23 VN.n22 50.0921
R144 VN.n13 VN.n2 24.9531
R145 VN.n31 VN.n20 24.9531
R146 VN.n7 VN.n4 24.4675
R147 VN.n8 VN.n7 24.4675
R148 VN.n9 VN.n8 24.4675
R149 VN.n14 VN.n13 24.4675
R150 VN.n15 VN.n14 24.4675
R151 VN.n27 VN.n26 24.4675
R152 VN.n26 VN.n25 24.4675
R153 VN.n25 VN.n22 24.4675
R154 VN.n33 VN.n32 24.4675
R155 VN.n32 VN.n31 24.4675
R156 VN.n15 VN.n0 8.80862
R157 VN.n33 VN.n18 8.80862
R158 VN.n24 VN.n23 3.1948
R159 VN.n6 VN.n5 3.1948
R160 VN.n35 VN.n34 0.354971
R161 VN.n17 VN.n16 0.354971
R162 VN VN.n17 0.26696
R163 VN.n34 VN.n19 0.189894
R164 VN.n30 VN.n19 0.189894
R165 VN.n30 VN.n29 0.189894
R166 VN.n29 VN.n28 0.189894
R167 VN.n28 VN.n21 0.189894
R168 VN.n24 VN.n21 0.189894
R169 VN.n6 VN.n3 0.189894
R170 VN.n10 VN.n3 0.189894
R171 VN.n11 VN.n10 0.189894
R172 VN.n12 VN.n11 0.189894
R173 VN.n12 VN.n1 0.189894
R174 VN.n16 VN.n1 0.189894
R175 VDD2.n1 VDD2.t3 74.7287
R176 VDD2.n2 VDD2.t5 72.405
R177 VDD2.n1 VDD2.n0 71.3336
R178 VDD2 VDD2.n3 71.3309
R179 VDD2.n2 VDD2.n1 49.517
R180 VDD2 VDD2.n2 2.438
R181 VDD2.n3 VDD2.t1 1.80935
R182 VDD2.n3 VDD2.t2 1.80935
R183 VDD2.n0 VDD2.t4 1.80935
R184 VDD2.n0 VDD2.t0 1.80935
R185 B.n509 B.n148 585
R186 B.n508 B.n507 585
R187 B.n506 B.n149 585
R188 B.n505 B.n504 585
R189 B.n503 B.n150 585
R190 B.n502 B.n501 585
R191 B.n500 B.n151 585
R192 B.n499 B.n498 585
R193 B.n497 B.n152 585
R194 B.n496 B.n495 585
R195 B.n494 B.n153 585
R196 B.n493 B.n492 585
R197 B.n491 B.n154 585
R198 B.n490 B.n489 585
R199 B.n488 B.n155 585
R200 B.n487 B.n486 585
R201 B.n485 B.n156 585
R202 B.n484 B.n483 585
R203 B.n482 B.n157 585
R204 B.n481 B.n480 585
R205 B.n479 B.n158 585
R206 B.n478 B.n477 585
R207 B.n476 B.n159 585
R208 B.n475 B.n474 585
R209 B.n473 B.n160 585
R210 B.n472 B.n471 585
R211 B.n470 B.n161 585
R212 B.n469 B.n468 585
R213 B.n467 B.n162 585
R214 B.n466 B.n465 585
R215 B.n464 B.n163 585
R216 B.n463 B.n462 585
R217 B.n461 B.n164 585
R218 B.n460 B.n459 585
R219 B.n458 B.n165 585
R220 B.n457 B.n456 585
R221 B.n455 B.n166 585
R222 B.n454 B.n453 585
R223 B.n452 B.n167 585
R224 B.n451 B.n450 585
R225 B.n449 B.n168 585
R226 B.n448 B.n447 585
R227 B.n446 B.n169 585
R228 B.n445 B.n444 585
R229 B.n443 B.n170 585
R230 B.n442 B.n441 585
R231 B.n440 B.n171 585
R232 B.n439 B.n438 585
R233 B.n437 B.n172 585
R234 B.n436 B.n435 585
R235 B.n434 B.n173 585
R236 B.n433 B.n432 585
R237 B.n431 B.n174 585
R238 B.n430 B.n429 585
R239 B.n428 B.n175 585
R240 B.n427 B.n426 585
R241 B.n425 B.n176 585
R242 B.n424 B.n423 585
R243 B.n422 B.n177 585
R244 B.n420 B.n419 585
R245 B.n418 B.n180 585
R246 B.n417 B.n416 585
R247 B.n415 B.n181 585
R248 B.n414 B.n413 585
R249 B.n412 B.n182 585
R250 B.n411 B.n410 585
R251 B.n409 B.n183 585
R252 B.n408 B.n407 585
R253 B.n406 B.n184 585
R254 B.n405 B.n404 585
R255 B.n400 B.n185 585
R256 B.n399 B.n398 585
R257 B.n397 B.n186 585
R258 B.n396 B.n395 585
R259 B.n394 B.n187 585
R260 B.n393 B.n392 585
R261 B.n391 B.n188 585
R262 B.n390 B.n389 585
R263 B.n388 B.n189 585
R264 B.n387 B.n386 585
R265 B.n385 B.n190 585
R266 B.n384 B.n383 585
R267 B.n382 B.n191 585
R268 B.n381 B.n380 585
R269 B.n379 B.n192 585
R270 B.n378 B.n377 585
R271 B.n376 B.n193 585
R272 B.n375 B.n374 585
R273 B.n373 B.n194 585
R274 B.n372 B.n371 585
R275 B.n370 B.n195 585
R276 B.n369 B.n368 585
R277 B.n367 B.n196 585
R278 B.n366 B.n365 585
R279 B.n364 B.n197 585
R280 B.n363 B.n362 585
R281 B.n361 B.n198 585
R282 B.n360 B.n359 585
R283 B.n358 B.n199 585
R284 B.n357 B.n356 585
R285 B.n355 B.n200 585
R286 B.n354 B.n353 585
R287 B.n352 B.n201 585
R288 B.n351 B.n350 585
R289 B.n349 B.n202 585
R290 B.n348 B.n347 585
R291 B.n346 B.n203 585
R292 B.n345 B.n344 585
R293 B.n343 B.n204 585
R294 B.n342 B.n341 585
R295 B.n340 B.n205 585
R296 B.n339 B.n338 585
R297 B.n337 B.n206 585
R298 B.n336 B.n335 585
R299 B.n334 B.n207 585
R300 B.n333 B.n332 585
R301 B.n331 B.n208 585
R302 B.n330 B.n329 585
R303 B.n328 B.n209 585
R304 B.n327 B.n326 585
R305 B.n325 B.n210 585
R306 B.n324 B.n323 585
R307 B.n322 B.n211 585
R308 B.n321 B.n320 585
R309 B.n319 B.n212 585
R310 B.n318 B.n317 585
R311 B.n316 B.n213 585
R312 B.n315 B.n314 585
R313 B.n511 B.n510 585
R314 B.n512 B.n147 585
R315 B.n514 B.n513 585
R316 B.n515 B.n146 585
R317 B.n517 B.n516 585
R318 B.n518 B.n145 585
R319 B.n520 B.n519 585
R320 B.n521 B.n144 585
R321 B.n523 B.n522 585
R322 B.n524 B.n143 585
R323 B.n526 B.n525 585
R324 B.n527 B.n142 585
R325 B.n529 B.n528 585
R326 B.n530 B.n141 585
R327 B.n532 B.n531 585
R328 B.n533 B.n140 585
R329 B.n535 B.n534 585
R330 B.n536 B.n139 585
R331 B.n538 B.n537 585
R332 B.n539 B.n138 585
R333 B.n541 B.n540 585
R334 B.n542 B.n137 585
R335 B.n544 B.n543 585
R336 B.n545 B.n136 585
R337 B.n547 B.n546 585
R338 B.n548 B.n135 585
R339 B.n550 B.n549 585
R340 B.n551 B.n134 585
R341 B.n553 B.n552 585
R342 B.n554 B.n133 585
R343 B.n556 B.n555 585
R344 B.n557 B.n132 585
R345 B.n559 B.n558 585
R346 B.n560 B.n131 585
R347 B.n562 B.n561 585
R348 B.n563 B.n130 585
R349 B.n565 B.n564 585
R350 B.n566 B.n129 585
R351 B.n568 B.n567 585
R352 B.n569 B.n128 585
R353 B.n571 B.n570 585
R354 B.n572 B.n127 585
R355 B.n574 B.n573 585
R356 B.n575 B.n126 585
R357 B.n577 B.n576 585
R358 B.n578 B.n125 585
R359 B.n580 B.n579 585
R360 B.n581 B.n124 585
R361 B.n583 B.n582 585
R362 B.n584 B.n123 585
R363 B.n586 B.n585 585
R364 B.n587 B.n122 585
R365 B.n589 B.n588 585
R366 B.n590 B.n121 585
R367 B.n592 B.n591 585
R368 B.n593 B.n120 585
R369 B.n595 B.n594 585
R370 B.n596 B.n119 585
R371 B.n598 B.n597 585
R372 B.n599 B.n118 585
R373 B.n601 B.n600 585
R374 B.n602 B.n117 585
R375 B.n604 B.n603 585
R376 B.n605 B.n116 585
R377 B.n607 B.n606 585
R378 B.n608 B.n115 585
R379 B.n610 B.n609 585
R380 B.n611 B.n114 585
R381 B.n613 B.n612 585
R382 B.n614 B.n113 585
R383 B.n616 B.n615 585
R384 B.n617 B.n112 585
R385 B.n619 B.n618 585
R386 B.n620 B.n111 585
R387 B.n622 B.n621 585
R388 B.n623 B.n110 585
R389 B.n625 B.n624 585
R390 B.n626 B.n109 585
R391 B.n628 B.n627 585
R392 B.n629 B.n108 585
R393 B.n631 B.n630 585
R394 B.n632 B.n107 585
R395 B.n634 B.n633 585
R396 B.n635 B.n106 585
R397 B.n637 B.n636 585
R398 B.n638 B.n105 585
R399 B.n640 B.n639 585
R400 B.n641 B.n104 585
R401 B.n643 B.n642 585
R402 B.n644 B.n103 585
R403 B.n646 B.n645 585
R404 B.n647 B.n102 585
R405 B.n649 B.n648 585
R406 B.n650 B.n101 585
R407 B.n652 B.n651 585
R408 B.n653 B.n100 585
R409 B.n655 B.n654 585
R410 B.n656 B.n99 585
R411 B.n658 B.n657 585
R412 B.n659 B.n98 585
R413 B.n661 B.n660 585
R414 B.n662 B.n97 585
R415 B.n664 B.n663 585
R416 B.n665 B.n96 585
R417 B.n859 B.n858 585
R418 B.n857 B.n28 585
R419 B.n856 B.n855 585
R420 B.n854 B.n29 585
R421 B.n853 B.n852 585
R422 B.n851 B.n30 585
R423 B.n850 B.n849 585
R424 B.n848 B.n31 585
R425 B.n847 B.n846 585
R426 B.n845 B.n32 585
R427 B.n844 B.n843 585
R428 B.n842 B.n33 585
R429 B.n841 B.n840 585
R430 B.n839 B.n34 585
R431 B.n838 B.n837 585
R432 B.n836 B.n35 585
R433 B.n835 B.n834 585
R434 B.n833 B.n36 585
R435 B.n832 B.n831 585
R436 B.n830 B.n37 585
R437 B.n829 B.n828 585
R438 B.n827 B.n38 585
R439 B.n826 B.n825 585
R440 B.n824 B.n39 585
R441 B.n823 B.n822 585
R442 B.n821 B.n40 585
R443 B.n820 B.n819 585
R444 B.n818 B.n41 585
R445 B.n817 B.n816 585
R446 B.n815 B.n42 585
R447 B.n814 B.n813 585
R448 B.n812 B.n43 585
R449 B.n811 B.n810 585
R450 B.n809 B.n44 585
R451 B.n808 B.n807 585
R452 B.n806 B.n45 585
R453 B.n805 B.n804 585
R454 B.n803 B.n46 585
R455 B.n802 B.n801 585
R456 B.n800 B.n47 585
R457 B.n799 B.n798 585
R458 B.n797 B.n48 585
R459 B.n796 B.n795 585
R460 B.n794 B.n49 585
R461 B.n793 B.n792 585
R462 B.n791 B.n50 585
R463 B.n790 B.n789 585
R464 B.n788 B.n51 585
R465 B.n787 B.n786 585
R466 B.n785 B.n52 585
R467 B.n784 B.n783 585
R468 B.n782 B.n53 585
R469 B.n781 B.n780 585
R470 B.n779 B.n54 585
R471 B.n778 B.n777 585
R472 B.n776 B.n55 585
R473 B.n775 B.n774 585
R474 B.n773 B.n56 585
R475 B.n772 B.n771 585
R476 B.n769 B.n57 585
R477 B.n768 B.n767 585
R478 B.n766 B.n60 585
R479 B.n765 B.n764 585
R480 B.n763 B.n61 585
R481 B.n762 B.n761 585
R482 B.n760 B.n62 585
R483 B.n759 B.n758 585
R484 B.n757 B.n63 585
R485 B.n756 B.n755 585
R486 B.n754 B.n753 585
R487 B.n752 B.n67 585
R488 B.n751 B.n750 585
R489 B.n749 B.n68 585
R490 B.n748 B.n747 585
R491 B.n746 B.n69 585
R492 B.n745 B.n744 585
R493 B.n743 B.n70 585
R494 B.n742 B.n741 585
R495 B.n740 B.n71 585
R496 B.n739 B.n738 585
R497 B.n737 B.n72 585
R498 B.n736 B.n735 585
R499 B.n734 B.n73 585
R500 B.n733 B.n732 585
R501 B.n731 B.n74 585
R502 B.n730 B.n729 585
R503 B.n728 B.n75 585
R504 B.n727 B.n726 585
R505 B.n725 B.n76 585
R506 B.n724 B.n723 585
R507 B.n722 B.n77 585
R508 B.n721 B.n720 585
R509 B.n719 B.n78 585
R510 B.n718 B.n717 585
R511 B.n716 B.n79 585
R512 B.n715 B.n714 585
R513 B.n713 B.n80 585
R514 B.n712 B.n711 585
R515 B.n710 B.n81 585
R516 B.n709 B.n708 585
R517 B.n707 B.n82 585
R518 B.n706 B.n705 585
R519 B.n704 B.n83 585
R520 B.n703 B.n702 585
R521 B.n701 B.n84 585
R522 B.n700 B.n699 585
R523 B.n698 B.n85 585
R524 B.n697 B.n696 585
R525 B.n695 B.n86 585
R526 B.n694 B.n693 585
R527 B.n692 B.n87 585
R528 B.n691 B.n690 585
R529 B.n689 B.n88 585
R530 B.n688 B.n687 585
R531 B.n686 B.n89 585
R532 B.n685 B.n684 585
R533 B.n683 B.n90 585
R534 B.n682 B.n681 585
R535 B.n680 B.n91 585
R536 B.n679 B.n678 585
R537 B.n677 B.n92 585
R538 B.n676 B.n675 585
R539 B.n674 B.n93 585
R540 B.n673 B.n672 585
R541 B.n671 B.n94 585
R542 B.n670 B.n669 585
R543 B.n668 B.n95 585
R544 B.n667 B.n666 585
R545 B.n860 B.n27 585
R546 B.n862 B.n861 585
R547 B.n863 B.n26 585
R548 B.n865 B.n864 585
R549 B.n866 B.n25 585
R550 B.n868 B.n867 585
R551 B.n869 B.n24 585
R552 B.n871 B.n870 585
R553 B.n872 B.n23 585
R554 B.n874 B.n873 585
R555 B.n875 B.n22 585
R556 B.n877 B.n876 585
R557 B.n878 B.n21 585
R558 B.n880 B.n879 585
R559 B.n881 B.n20 585
R560 B.n883 B.n882 585
R561 B.n884 B.n19 585
R562 B.n886 B.n885 585
R563 B.n887 B.n18 585
R564 B.n889 B.n888 585
R565 B.n890 B.n17 585
R566 B.n892 B.n891 585
R567 B.n893 B.n16 585
R568 B.n895 B.n894 585
R569 B.n896 B.n15 585
R570 B.n898 B.n897 585
R571 B.n899 B.n14 585
R572 B.n901 B.n900 585
R573 B.n902 B.n13 585
R574 B.n904 B.n903 585
R575 B.n905 B.n12 585
R576 B.n907 B.n906 585
R577 B.n908 B.n11 585
R578 B.n910 B.n909 585
R579 B.n911 B.n10 585
R580 B.n913 B.n912 585
R581 B.n914 B.n9 585
R582 B.n916 B.n915 585
R583 B.n917 B.n8 585
R584 B.n919 B.n918 585
R585 B.n920 B.n7 585
R586 B.n922 B.n921 585
R587 B.n923 B.n6 585
R588 B.n925 B.n924 585
R589 B.n926 B.n5 585
R590 B.n928 B.n927 585
R591 B.n929 B.n4 585
R592 B.n931 B.n930 585
R593 B.n932 B.n3 585
R594 B.n934 B.n933 585
R595 B.n935 B.n0 585
R596 B.n2 B.n1 585
R597 B.n240 B.n239 585
R598 B.n241 B.n238 585
R599 B.n243 B.n242 585
R600 B.n244 B.n237 585
R601 B.n246 B.n245 585
R602 B.n247 B.n236 585
R603 B.n249 B.n248 585
R604 B.n250 B.n235 585
R605 B.n252 B.n251 585
R606 B.n253 B.n234 585
R607 B.n255 B.n254 585
R608 B.n256 B.n233 585
R609 B.n258 B.n257 585
R610 B.n259 B.n232 585
R611 B.n261 B.n260 585
R612 B.n262 B.n231 585
R613 B.n264 B.n263 585
R614 B.n265 B.n230 585
R615 B.n267 B.n266 585
R616 B.n268 B.n229 585
R617 B.n270 B.n269 585
R618 B.n271 B.n228 585
R619 B.n273 B.n272 585
R620 B.n274 B.n227 585
R621 B.n276 B.n275 585
R622 B.n277 B.n226 585
R623 B.n279 B.n278 585
R624 B.n280 B.n225 585
R625 B.n282 B.n281 585
R626 B.n283 B.n224 585
R627 B.n285 B.n284 585
R628 B.n286 B.n223 585
R629 B.n288 B.n287 585
R630 B.n289 B.n222 585
R631 B.n291 B.n290 585
R632 B.n292 B.n221 585
R633 B.n294 B.n293 585
R634 B.n295 B.n220 585
R635 B.n297 B.n296 585
R636 B.n298 B.n219 585
R637 B.n300 B.n299 585
R638 B.n301 B.n218 585
R639 B.n303 B.n302 585
R640 B.n304 B.n217 585
R641 B.n306 B.n305 585
R642 B.n307 B.n216 585
R643 B.n309 B.n308 585
R644 B.n310 B.n215 585
R645 B.n312 B.n311 585
R646 B.n313 B.n214 585
R647 B.n314 B.n313 478.086
R648 B.n510 B.n509 478.086
R649 B.n666 B.n665 478.086
R650 B.n858 B.n27 478.086
R651 B.n401 B.t0 338.231
R652 B.n178 B.t3 338.231
R653 B.n64 B.t9 338.231
R654 B.n58 B.t6 338.231
R655 B.n937 B.n936 256.663
R656 B.n936 B.n935 235.042
R657 B.n936 B.n2 235.042
R658 B.n178 B.t4 183.201
R659 B.n64 B.t11 183.201
R660 B.n401 B.t1 183.178
R661 B.n58 B.t8 183.178
R662 B.n314 B.n213 163.367
R663 B.n318 B.n213 163.367
R664 B.n319 B.n318 163.367
R665 B.n320 B.n319 163.367
R666 B.n320 B.n211 163.367
R667 B.n324 B.n211 163.367
R668 B.n325 B.n324 163.367
R669 B.n326 B.n325 163.367
R670 B.n326 B.n209 163.367
R671 B.n330 B.n209 163.367
R672 B.n331 B.n330 163.367
R673 B.n332 B.n331 163.367
R674 B.n332 B.n207 163.367
R675 B.n336 B.n207 163.367
R676 B.n337 B.n336 163.367
R677 B.n338 B.n337 163.367
R678 B.n338 B.n205 163.367
R679 B.n342 B.n205 163.367
R680 B.n343 B.n342 163.367
R681 B.n344 B.n343 163.367
R682 B.n344 B.n203 163.367
R683 B.n348 B.n203 163.367
R684 B.n349 B.n348 163.367
R685 B.n350 B.n349 163.367
R686 B.n350 B.n201 163.367
R687 B.n354 B.n201 163.367
R688 B.n355 B.n354 163.367
R689 B.n356 B.n355 163.367
R690 B.n356 B.n199 163.367
R691 B.n360 B.n199 163.367
R692 B.n361 B.n360 163.367
R693 B.n362 B.n361 163.367
R694 B.n362 B.n197 163.367
R695 B.n366 B.n197 163.367
R696 B.n367 B.n366 163.367
R697 B.n368 B.n367 163.367
R698 B.n368 B.n195 163.367
R699 B.n372 B.n195 163.367
R700 B.n373 B.n372 163.367
R701 B.n374 B.n373 163.367
R702 B.n374 B.n193 163.367
R703 B.n378 B.n193 163.367
R704 B.n379 B.n378 163.367
R705 B.n380 B.n379 163.367
R706 B.n380 B.n191 163.367
R707 B.n384 B.n191 163.367
R708 B.n385 B.n384 163.367
R709 B.n386 B.n385 163.367
R710 B.n386 B.n189 163.367
R711 B.n390 B.n189 163.367
R712 B.n391 B.n390 163.367
R713 B.n392 B.n391 163.367
R714 B.n392 B.n187 163.367
R715 B.n396 B.n187 163.367
R716 B.n397 B.n396 163.367
R717 B.n398 B.n397 163.367
R718 B.n398 B.n185 163.367
R719 B.n405 B.n185 163.367
R720 B.n406 B.n405 163.367
R721 B.n407 B.n406 163.367
R722 B.n407 B.n183 163.367
R723 B.n411 B.n183 163.367
R724 B.n412 B.n411 163.367
R725 B.n413 B.n412 163.367
R726 B.n413 B.n181 163.367
R727 B.n417 B.n181 163.367
R728 B.n418 B.n417 163.367
R729 B.n419 B.n418 163.367
R730 B.n419 B.n177 163.367
R731 B.n424 B.n177 163.367
R732 B.n425 B.n424 163.367
R733 B.n426 B.n425 163.367
R734 B.n426 B.n175 163.367
R735 B.n430 B.n175 163.367
R736 B.n431 B.n430 163.367
R737 B.n432 B.n431 163.367
R738 B.n432 B.n173 163.367
R739 B.n436 B.n173 163.367
R740 B.n437 B.n436 163.367
R741 B.n438 B.n437 163.367
R742 B.n438 B.n171 163.367
R743 B.n442 B.n171 163.367
R744 B.n443 B.n442 163.367
R745 B.n444 B.n443 163.367
R746 B.n444 B.n169 163.367
R747 B.n448 B.n169 163.367
R748 B.n449 B.n448 163.367
R749 B.n450 B.n449 163.367
R750 B.n450 B.n167 163.367
R751 B.n454 B.n167 163.367
R752 B.n455 B.n454 163.367
R753 B.n456 B.n455 163.367
R754 B.n456 B.n165 163.367
R755 B.n460 B.n165 163.367
R756 B.n461 B.n460 163.367
R757 B.n462 B.n461 163.367
R758 B.n462 B.n163 163.367
R759 B.n466 B.n163 163.367
R760 B.n467 B.n466 163.367
R761 B.n468 B.n467 163.367
R762 B.n468 B.n161 163.367
R763 B.n472 B.n161 163.367
R764 B.n473 B.n472 163.367
R765 B.n474 B.n473 163.367
R766 B.n474 B.n159 163.367
R767 B.n478 B.n159 163.367
R768 B.n479 B.n478 163.367
R769 B.n480 B.n479 163.367
R770 B.n480 B.n157 163.367
R771 B.n484 B.n157 163.367
R772 B.n485 B.n484 163.367
R773 B.n486 B.n485 163.367
R774 B.n486 B.n155 163.367
R775 B.n490 B.n155 163.367
R776 B.n491 B.n490 163.367
R777 B.n492 B.n491 163.367
R778 B.n492 B.n153 163.367
R779 B.n496 B.n153 163.367
R780 B.n497 B.n496 163.367
R781 B.n498 B.n497 163.367
R782 B.n498 B.n151 163.367
R783 B.n502 B.n151 163.367
R784 B.n503 B.n502 163.367
R785 B.n504 B.n503 163.367
R786 B.n504 B.n149 163.367
R787 B.n508 B.n149 163.367
R788 B.n509 B.n508 163.367
R789 B.n665 B.n664 163.367
R790 B.n664 B.n97 163.367
R791 B.n660 B.n97 163.367
R792 B.n660 B.n659 163.367
R793 B.n659 B.n658 163.367
R794 B.n658 B.n99 163.367
R795 B.n654 B.n99 163.367
R796 B.n654 B.n653 163.367
R797 B.n653 B.n652 163.367
R798 B.n652 B.n101 163.367
R799 B.n648 B.n101 163.367
R800 B.n648 B.n647 163.367
R801 B.n647 B.n646 163.367
R802 B.n646 B.n103 163.367
R803 B.n642 B.n103 163.367
R804 B.n642 B.n641 163.367
R805 B.n641 B.n640 163.367
R806 B.n640 B.n105 163.367
R807 B.n636 B.n105 163.367
R808 B.n636 B.n635 163.367
R809 B.n635 B.n634 163.367
R810 B.n634 B.n107 163.367
R811 B.n630 B.n107 163.367
R812 B.n630 B.n629 163.367
R813 B.n629 B.n628 163.367
R814 B.n628 B.n109 163.367
R815 B.n624 B.n109 163.367
R816 B.n624 B.n623 163.367
R817 B.n623 B.n622 163.367
R818 B.n622 B.n111 163.367
R819 B.n618 B.n111 163.367
R820 B.n618 B.n617 163.367
R821 B.n617 B.n616 163.367
R822 B.n616 B.n113 163.367
R823 B.n612 B.n113 163.367
R824 B.n612 B.n611 163.367
R825 B.n611 B.n610 163.367
R826 B.n610 B.n115 163.367
R827 B.n606 B.n115 163.367
R828 B.n606 B.n605 163.367
R829 B.n605 B.n604 163.367
R830 B.n604 B.n117 163.367
R831 B.n600 B.n117 163.367
R832 B.n600 B.n599 163.367
R833 B.n599 B.n598 163.367
R834 B.n598 B.n119 163.367
R835 B.n594 B.n119 163.367
R836 B.n594 B.n593 163.367
R837 B.n593 B.n592 163.367
R838 B.n592 B.n121 163.367
R839 B.n588 B.n121 163.367
R840 B.n588 B.n587 163.367
R841 B.n587 B.n586 163.367
R842 B.n586 B.n123 163.367
R843 B.n582 B.n123 163.367
R844 B.n582 B.n581 163.367
R845 B.n581 B.n580 163.367
R846 B.n580 B.n125 163.367
R847 B.n576 B.n125 163.367
R848 B.n576 B.n575 163.367
R849 B.n575 B.n574 163.367
R850 B.n574 B.n127 163.367
R851 B.n570 B.n127 163.367
R852 B.n570 B.n569 163.367
R853 B.n569 B.n568 163.367
R854 B.n568 B.n129 163.367
R855 B.n564 B.n129 163.367
R856 B.n564 B.n563 163.367
R857 B.n563 B.n562 163.367
R858 B.n562 B.n131 163.367
R859 B.n558 B.n131 163.367
R860 B.n558 B.n557 163.367
R861 B.n557 B.n556 163.367
R862 B.n556 B.n133 163.367
R863 B.n552 B.n133 163.367
R864 B.n552 B.n551 163.367
R865 B.n551 B.n550 163.367
R866 B.n550 B.n135 163.367
R867 B.n546 B.n135 163.367
R868 B.n546 B.n545 163.367
R869 B.n545 B.n544 163.367
R870 B.n544 B.n137 163.367
R871 B.n540 B.n137 163.367
R872 B.n540 B.n539 163.367
R873 B.n539 B.n538 163.367
R874 B.n538 B.n139 163.367
R875 B.n534 B.n139 163.367
R876 B.n534 B.n533 163.367
R877 B.n533 B.n532 163.367
R878 B.n532 B.n141 163.367
R879 B.n528 B.n141 163.367
R880 B.n528 B.n527 163.367
R881 B.n527 B.n526 163.367
R882 B.n526 B.n143 163.367
R883 B.n522 B.n143 163.367
R884 B.n522 B.n521 163.367
R885 B.n521 B.n520 163.367
R886 B.n520 B.n145 163.367
R887 B.n516 B.n145 163.367
R888 B.n516 B.n515 163.367
R889 B.n515 B.n514 163.367
R890 B.n514 B.n147 163.367
R891 B.n510 B.n147 163.367
R892 B.n858 B.n857 163.367
R893 B.n857 B.n856 163.367
R894 B.n856 B.n29 163.367
R895 B.n852 B.n29 163.367
R896 B.n852 B.n851 163.367
R897 B.n851 B.n850 163.367
R898 B.n850 B.n31 163.367
R899 B.n846 B.n31 163.367
R900 B.n846 B.n845 163.367
R901 B.n845 B.n844 163.367
R902 B.n844 B.n33 163.367
R903 B.n840 B.n33 163.367
R904 B.n840 B.n839 163.367
R905 B.n839 B.n838 163.367
R906 B.n838 B.n35 163.367
R907 B.n834 B.n35 163.367
R908 B.n834 B.n833 163.367
R909 B.n833 B.n832 163.367
R910 B.n832 B.n37 163.367
R911 B.n828 B.n37 163.367
R912 B.n828 B.n827 163.367
R913 B.n827 B.n826 163.367
R914 B.n826 B.n39 163.367
R915 B.n822 B.n39 163.367
R916 B.n822 B.n821 163.367
R917 B.n821 B.n820 163.367
R918 B.n820 B.n41 163.367
R919 B.n816 B.n41 163.367
R920 B.n816 B.n815 163.367
R921 B.n815 B.n814 163.367
R922 B.n814 B.n43 163.367
R923 B.n810 B.n43 163.367
R924 B.n810 B.n809 163.367
R925 B.n809 B.n808 163.367
R926 B.n808 B.n45 163.367
R927 B.n804 B.n45 163.367
R928 B.n804 B.n803 163.367
R929 B.n803 B.n802 163.367
R930 B.n802 B.n47 163.367
R931 B.n798 B.n47 163.367
R932 B.n798 B.n797 163.367
R933 B.n797 B.n796 163.367
R934 B.n796 B.n49 163.367
R935 B.n792 B.n49 163.367
R936 B.n792 B.n791 163.367
R937 B.n791 B.n790 163.367
R938 B.n790 B.n51 163.367
R939 B.n786 B.n51 163.367
R940 B.n786 B.n785 163.367
R941 B.n785 B.n784 163.367
R942 B.n784 B.n53 163.367
R943 B.n780 B.n53 163.367
R944 B.n780 B.n779 163.367
R945 B.n779 B.n778 163.367
R946 B.n778 B.n55 163.367
R947 B.n774 B.n55 163.367
R948 B.n774 B.n773 163.367
R949 B.n773 B.n772 163.367
R950 B.n772 B.n57 163.367
R951 B.n767 B.n57 163.367
R952 B.n767 B.n766 163.367
R953 B.n766 B.n765 163.367
R954 B.n765 B.n61 163.367
R955 B.n761 B.n61 163.367
R956 B.n761 B.n760 163.367
R957 B.n760 B.n759 163.367
R958 B.n759 B.n63 163.367
R959 B.n755 B.n63 163.367
R960 B.n755 B.n754 163.367
R961 B.n754 B.n67 163.367
R962 B.n750 B.n67 163.367
R963 B.n750 B.n749 163.367
R964 B.n749 B.n748 163.367
R965 B.n748 B.n69 163.367
R966 B.n744 B.n69 163.367
R967 B.n744 B.n743 163.367
R968 B.n743 B.n742 163.367
R969 B.n742 B.n71 163.367
R970 B.n738 B.n71 163.367
R971 B.n738 B.n737 163.367
R972 B.n737 B.n736 163.367
R973 B.n736 B.n73 163.367
R974 B.n732 B.n73 163.367
R975 B.n732 B.n731 163.367
R976 B.n731 B.n730 163.367
R977 B.n730 B.n75 163.367
R978 B.n726 B.n75 163.367
R979 B.n726 B.n725 163.367
R980 B.n725 B.n724 163.367
R981 B.n724 B.n77 163.367
R982 B.n720 B.n77 163.367
R983 B.n720 B.n719 163.367
R984 B.n719 B.n718 163.367
R985 B.n718 B.n79 163.367
R986 B.n714 B.n79 163.367
R987 B.n714 B.n713 163.367
R988 B.n713 B.n712 163.367
R989 B.n712 B.n81 163.367
R990 B.n708 B.n81 163.367
R991 B.n708 B.n707 163.367
R992 B.n707 B.n706 163.367
R993 B.n706 B.n83 163.367
R994 B.n702 B.n83 163.367
R995 B.n702 B.n701 163.367
R996 B.n701 B.n700 163.367
R997 B.n700 B.n85 163.367
R998 B.n696 B.n85 163.367
R999 B.n696 B.n695 163.367
R1000 B.n695 B.n694 163.367
R1001 B.n694 B.n87 163.367
R1002 B.n690 B.n87 163.367
R1003 B.n690 B.n689 163.367
R1004 B.n689 B.n688 163.367
R1005 B.n688 B.n89 163.367
R1006 B.n684 B.n89 163.367
R1007 B.n684 B.n683 163.367
R1008 B.n683 B.n682 163.367
R1009 B.n682 B.n91 163.367
R1010 B.n678 B.n91 163.367
R1011 B.n678 B.n677 163.367
R1012 B.n677 B.n676 163.367
R1013 B.n676 B.n93 163.367
R1014 B.n672 B.n93 163.367
R1015 B.n672 B.n671 163.367
R1016 B.n671 B.n670 163.367
R1017 B.n670 B.n95 163.367
R1018 B.n666 B.n95 163.367
R1019 B.n862 B.n27 163.367
R1020 B.n863 B.n862 163.367
R1021 B.n864 B.n863 163.367
R1022 B.n864 B.n25 163.367
R1023 B.n868 B.n25 163.367
R1024 B.n869 B.n868 163.367
R1025 B.n870 B.n869 163.367
R1026 B.n870 B.n23 163.367
R1027 B.n874 B.n23 163.367
R1028 B.n875 B.n874 163.367
R1029 B.n876 B.n875 163.367
R1030 B.n876 B.n21 163.367
R1031 B.n880 B.n21 163.367
R1032 B.n881 B.n880 163.367
R1033 B.n882 B.n881 163.367
R1034 B.n882 B.n19 163.367
R1035 B.n886 B.n19 163.367
R1036 B.n887 B.n886 163.367
R1037 B.n888 B.n887 163.367
R1038 B.n888 B.n17 163.367
R1039 B.n892 B.n17 163.367
R1040 B.n893 B.n892 163.367
R1041 B.n894 B.n893 163.367
R1042 B.n894 B.n15 163.367
R1043 B.n898 B.n15 163.367
R1044 B.n899 B.n898 163.367
R1045 B.n900 B.n899 163.367
R1046 B.n900 B.n13 163.367
R1047 B.n904 B.n13 163.367
R1048 B.n905 B.n904 163.367
R1049 B.n906 B.n905 163.367
R1050 B.n906 B.n11 163.367
R1051 B.n910 B.n11 163.367
R1052 B.n911 B.n910 163.367
R1053 B.n912 B.n911 163.367
R1054 B.n912 B.n9 163.367
R1055 B.n916 B.n9 163.367
R1056 B.n917 B.n916 163.367
R1057 B.n918 B.n917 163.367
R1058 B.n918 B.n7 163.367
R1059 B.n922 B.n7 163.367
R1060 B.n923 B.n922 163.367
R1061 B.n924 B.n923 163.367
R1062 B.n924 B.n5 163.367
R1063 B.n928 B.n5 163.367
R1064 B.n929 B.n928 163.367
R1065 B.n930 B.n929 163.367
R1066 B.n930 B.n3 163.367
R1067 B.n934 B.n3 163.367
R1068 B.n935 B.n934 163.367
R1069 B.n240 B.n2 163.367
R1070 B.n241 B.n240 163.367
R1071 B.n242 B.n241 163.367
R1072 B.n242 B.n237 163.367
R1073 B.n246 B.n237 163.367
R1074 B.n247 B.n246 163.367
R1075 B.n248 B.n247 163.367
R1076 B.n248 B.n235 163.367
R1077 B.n252 B.n235 163.367
R1078 B.n253 B.n252 163.367
R1079 B.n254 B.n253 163.367
R1080 B.n254 B.n233 163.367
R1081 B.n258 B.n233 163.367
R1082 B.n259 B.n258 163.367
R1083 B.n260 B.n259 163.367
R1084 B.n260 B.n231 163.367
R1085 B.n264 B.n231 163.367
R1086 B.n265 B.n264 163.367
R1087 B.n266 B.n265 163.367
R1088 B.n266 B.n229 163.367
R1089 B.n270 B.n229 163.367
R1090 B.n271 B.n270 163.367
R1091 B.n272 B.n271 163.367
R1092 B.n272 B.n227 163.367
R1093 B.n276 B.n227 163.367
R1094 B.n277 B.n276 163.367
R1095 B.n278 B.n277 163.367
R1096 B.n278 B.n225 163.367
R1097 B.n282 B.n225 163.367
R1098 B.n283 B.n282 163.367
R1099 B.n284 B.n283 163.367
R1100 B.n284 B.n223 163.367
R1101 B.n288 B.n223 163.367
R1102 B.n289 B.n288 163.367
R1103 B.n290 B.n289 163.367
R1104 B.n290 B.n221 163.367
R1105 B.n294 B.n221 163.367
R1106 B.n295 B.n294 163.367
R1107 B.n296 B.n295 163.367
R1108 B.n296 B.n219 163.367
R1109 B.n300 B.n219 163.367
R1110 B.n301 B.n300 163.367
R1111 B.n302 B.n301 163.367
R1112 B.n302 B.n217 163.367
R1113 B.n306 B.n217 163.367
R1114 B.n307 B.n306 163.367
R1115 B.n308 B.n307 163.367
R1116 B.n308 B.n215 163.367
R1117 B.n312 B.n215 163.367
R1118 B.n313 B.n312 163.367
R1119 B.n179 B.t5 111.832
R1120 B.n65 B.t10 111.832
R1121 B.n402 B.t2 111.808
R1122 B.n59 B.t7 111.808
R1123 B.n402 B.n401 71.3702
R1124 B.n179 B.n178 71.3702
R1125 B.n65 B.n64 71.3702
R1126 B.n59 B.n58 71.3702
R1127 B.n403 B.n402 59.5399
R1128 B.n421 B.n179 59.5399
R1129 B.n66 B.n65 59.5399
R1130 B.n770 B.n59 59.5399
R1131 B.n860 B.n859 31.0639
R1132 B.n667 B.n96 31.0639
R1133 B.n511 B.n148 31.0639
R1134 B.n315 B.n214 31.0639
R1135 B B.n937 18.0485
R1136 B.n861 B.n860 10.6151
R1137 B.n861 B.n26 10.6151
R1138 B.n865 B.n26 10.6151
R1139 B.n866 B.n865 10.6151
R1140 B.n867 B.n866 10.6151
R1141 B.n867 B.n24 10.6151
R1142 B.n871 B.n24 10.6151
R1143 B.n872 B.n871 10.6151
R1144 B.n873 B.n872 10.6151
R1145 B.n873 B.n22 10.6151
R1146 B.n877 B.n22 10.6151
R1147 B.n878 B.n877 10.6151
R1148 B.n879 B.n878 10.6151
R1149 B.n879 B.n20 10.6151
R1150 B.n883 B.n20 10.6151
R1151 B.n884 B.n883 10.6151
R1152 B.n885 B.n884 10.6151
R1153 B.n885 B.n18 10.6151
R1154 B.n889 B.n18 10.6151
R1155 B.n890 B.n889 10.6151
R1156 B.n891 B.n890 10.6151
R1157 B.n891 B.n16 10.6151
R1158 B.n895 B.n16 10.6151
R1159 B.n896 B.n895 10.6151
R1160 B.n897 B.n896 10.6151
R1161 B.n897 B.n14 10.6151
R1162 B.n901 B.n14 10.6151
R1163 B.n902 B.n901 10.6151
R1164 B.n903 B.n902 10.6151
R1165 B.n903 B.n12 10.6151
R1166 B.n907 B.n12 10.6151
R1167 B.n908 B.n907 10.6151
R1168 B.n909 B.n908 10.6151
R1169 B.n909 B.n10 10.6151
R1170 B.n913 B.n10 10.6151
R1171 B.n914 B.n913 10.6151
R1172 B.n915 B.n914 10.6151
R1173 B.n915 B.n8 10.6151
R1174 B.n919 B.n8 10.6151
R1175 B.n920 B.n919 10.6151
R1176 B.n921 B.n920 10.6151
R1177 B.n921 B.n6 10.6151
R1178 B.n925 B.n6 10.6151
R1179 B.n926 B.n925 10.6151
R1180 B.n927 B.n926 10.6151
R1181 B.n927 B.n4 10.6151
R1182 B.n931 B.n4 10.6151
R1183 B.n932 B.n931 10.6151
R1184 B.n933 B.n932 10.6151
R1185 B.n933 B.n0 10.6151
R1186 B.n859 B.n28 10.6151
R1187 B.n855 B.n28 10.6151
R1188 B.n855 B.n854 10.6151
R1189 B.n854 B.n853 10.6151
R1190 B.n853 B.n30 10.6151
R1191 B.n849 B.n30 10.6151
R1192 B.n849 B.n848 10.6151
R1193 B.n848 B.n847 10.6151
R1194 B.n847 B.n32 10.6151
R1195 B.n843 B.n32 10.6151
R1196 B.n843 B.n842 10.6151
R1197 B.n842 B.n841 10.6151
R1198 B.n841 B.n34 10.6151
R1199 B.n837 B.n34 10.6151
R1200 B.n837 B.n836 10.6151
R1201 B.n836 B.n835 10.6151
R1202 B.n835 B.n36 10.6151
R1203 B.n831 B.n36 10.6151
R1204 B.n831 B.n830 10.6151
R1205 B.n830 B.n829 10.6151
R1206 B.n829 B.n38 10.6151
R1207 B.n825 B.n38 10.6151
R1208 B.n825 B.n824 10.6151
R1209 B.n824 B.n823 10.6151
R1210 B.n823 B.n40 10.6151
R1211 B.n819 B.n40 10.6151
R1212 B.n819 B.n818 10.6151
R1213 B.n818 B.n817 10.6151
R1214 B.n817 B.n42 10.6151
R1215 B.n813 B.n42 10.6151
R1216 B.n813 B.n812 10.6151
R1217 B.n812 B.n811 10.6151
R1218 B.n811 B.n44 10.6151
R1219 B.n807 B.n44 10.6151
R1220 B.n807 B.n806 10.6151
R1221 B.n806 B.n805 10.6151
R1222 B.n805 B.n46 10.6151
R1223 B.n801 B.n46 10.6151
R1224 B.n801 B.n800 10.6151
R1225 B.n800 B.n799 10.6151
R1226 B.n799 B.n48 10.6151
R1227 B.n795 B.n48 10.6151
R1228 B.n795 B.n794 10.6151
R1229 B.n794 B.n793 10.6151
R1230 B.n793 B.n50 10.6151
R1231 B.n789 B.n50 10.6151
R1232 B.n789 B.n788 10.6151
R1233 B.n788 B.n787 10.6151
R1234 B.n787 B.n52 10.6151
R1235 B.n783 B.n52 10.6151
R1236 B.n783 B.n782 10.6151
R1237 B.n782 B.n781 10.6151
R1238 B.n781 B.n54 10.6151
R1239 B.n777 B.n54 10.6151
R1240 B.n777 B.n776 10.6151
R1241 B.n776 B.n775 10.6151
R1242 B.n775 B.n56 10.6151
R1243 B.n771 B.n56 10.6151
R1244 B.n769 B.n768 10.6151
R1245 B.n768 B.n60 10.6151
R1246 B.n764 B.n60 10.6151
R1247 B.n764 B.n763 10.6151
R1248 B.n763 B.n762 10.6151
R1249 B.n762 B.n62 10.6151
R1250 B.n758 B.n62 10.6151
R1251 B.n758 B.n757 10.6151
R1252 B.n757 B.n756 10.6151
R1253 B.n753 B.n752 10.6151
R1254 B.n752 B.n751 10.6151
R1255 B.n751 B.n68 10.6151
R1256 B.n747 B.n68 10.6151
R1257 B.n747 B.n746 10.6151
R1258 B.n746 B.n745 10.6151
R1259 B.n745 B.n70 10.6151
R1260 B.n741 B.n70 10.6151
R1261 B.n741 B.n740 10.6151
R1262 B.n740 B.n739 10.6151
R1263 B.n739 B.n72 10.6151
R1264 B.n735 B.n72 10.6151
R1265 B.n735 B.n734 10.6151
R1266 B.n734 B.n733 10.6151
R1267 B.n733 B.n74 10.6151
R1268 B.n729 B.n74 10.6151
R1269 B.n729 B.n728 10.6151
R1270 B.n728 B.n727 10.6151
R1271 B.n727 B.n76 10.6151
R1272 B.n723 B.n76 10.6151
R1273 B.n723 B.n722 10.6151
R1274 B.n722 B.n721 10.6151
R1275 B.n721 B.n78 10.6151
R1276 B.n717 B.n78 10.6151
R1277 B.n717 B.n716 10.6151
R1278 B.n716 B.n715 10.6151
R1279 B.n715 B.n80 10.6151
R1280 B.n711 B.n80 10.6151
R1281 B.n711 B.n710 10.6151
R1282 B.n710 B.n709 10.6151
R1283 B.n709 B.n82 10.6151
R1284 B.n705 B.n82 10.6151
R1285 B.n705 B.n704 10.6151
R1286 B.n704 B.n703 10.6151
R1287 B.n703 B.n84 10.6151
R1288 B.n699 B.n84 10.6151
R1289 B.n699 B.n698 10.6151
R1290 B.n698 B.n697 10.6151
R1291 B.n697 B.n86 10.6151
R1292 B.n693 B.n86 10.6151
R1293 B.n693 B.n692 10.6151
R1294 B.n692 B.n691 10.6151
R1295 B.n691 B.n88 10.6151
R1296 B.n687 B.n88 10.6151
R1297 B.n687 B.n686 10.6151
R1298 B.n686 B.n685 10.6151
R1299 B.n685 B.n90 10.6151
R1300 B.n681 B.n90 10.6151
R1301 B.n681 B.n680 10.6151
R1302 B.n680 B.n679 10.6151
R1303 B.n679 B.n92 10.6151
R1304 B.n675 B.n92 10.6151
R1305 B.n675 B.n674 10.6151
R1306 B.n674 B.n673 10.6151
R1307 B.n673 B.n94 10.6151
R1308 B.n669 B.n94 10.6151
R1309 B.n669 B.n668 10.6151
R1310 B.n668 B.n667 10.6151
R1311 B.n663 B.n96 10.6151
R1312 B.n663 B.n662 10.6151
R1313 B.n662 B.n661 10.6151
R1314 B.n661 B.n98 10.6151
R1315 B.n657 B.n98 10.6151
R1316 B.n657 B.n656 10.6151
R1317 B.n656 B.n655 10.6151
R1318 B.n655 B.n100 10.6151
R1319 B.n651 B.n100 10.6151
R1320 B.n651 B.n650 10.6151
R1321 B.n650 B.n649 10.6151
R1322 B.n649 B.n102 10.6151
R1323 B.n645 B.n102 10.6151
R1324 B.n645 B.n644 10.6151
R1325 B.n644 B.n643 10.6151
R1326 B.n643 B.n104 10.6151
R1327 B.n639 B.n104 10.6151
R1328 B.n639 B.n638 10.6151
R1329 B.n638 B.n637 10.6151
R1330 B.n637 B.n106 10.6151
R1331 B.n633 B.n106 10.6151
R1332 B.n633 B.n632 10.6151
R1333 B.n632 B.n631 10.6151
R1334 B.n631 B.n108 10.6151
R1335 B.n627 B.n108 10.6151
R1336 B.n627 B.n626 10.6151
R1337 B.n626 B.n625 10.6151
R1338 B.n625 B.n110 10.6151
R1339 B.n621 B.n110 10.6151
R1340 B.n621 B.n620 10.6151
R1341 B.n620 B.n619 10.6151
R1342 B.n619 B.n112 10.6151
R1343 B.n615 B.n112 10.6151
R1344 B.n615 B.n614 10.6151
R1345 B.n614 B.n613 10.6151
R1346 B.n613 B.n114 10.6151
R1347 B.n609 B.n114 10.6151
R1348 B.n609 B.n608 10.6151
R1349 B.n608 B.n607 10.6151
R1350 B.n607 B.n116 10.6151
R1351 B.n603 B.n116 10.6151
R1352 B.n603 B.n602 10.6151
R1353 B.n602 B.n601 10.6151
R1354 B.n601 B.n118 10.6151
R1355 B.n597 B.n118 10.6151
R1356 B.n597 B.n596 10.6151
R1357 B.n596 B.n595 10.6151
R1358 B.n595 B.n120 10.6151
R1359 B.n591 B.n120 10.6151
R1360 B.n591 B.n590 10.6151
R1361 B.n590 B.n589 10.6151
R1362 B.n589 B.n122 10.6151
R1363 B.n585 B.n122 10.6151
R1364 B.n585 B.n584 10.6151
R1365 B.n584 B.n583 10.6151
R1366 B.n583 B.n124 10.6151
R1367 B.n579 B.n124 10.6151
R1368 B.n579 B.n578 10.6151
R1369 B.n578 B.n577 10.6151
R1370 B.n577 B.n126 10.6151
R1371 B.n573 B.n126 10.6151
R1372 B.n573 B.n572 10.6151
R1373 B.n572 B.n571 10.6151
R1374 B.n571 B.n128 10.6151
R1375 B.n567 B.n128 10.6151
R1376 B.n567 B.n566 10.6151
R1377 B.n566 B.n565 10.6151
R1378 B.n565 B.n130 10.6151
R1379 B.n561 B.n130 10.6151
R1380 B.n561 B.n560 10.6151
R1381 B.n560 B.n559 10.6151
R1382 B.n559 B.n132 10.6151
R1383 B.n555 B.n132 10.6151
R1384 B.n555 B.n554 10.6151
R1385 B.n554 B.n553 10.6151
R1386 B.n553 B.n134 10.6151
R1387 B.n549 B.n134 10.6151
R1388 B.n549 B.n548 10.6151
R1389 B.n548 B.n547 10.6151
R1390 B.n547 B.n136 10.6151
R1391 B.n543 B.n136 10.6151
R1392 B.n543 B.n542 10.6151
R1393 B.n542 B.n541 10.6151
R1394 B.n541 B.n138 10.6151
R1395 B.n537 B.n138 10.6151
R1396 B.n537 B.n536 10.6151
R1397 B.n536 B.n535 10.6151
R1398 B.n535 B.n140 10.6151
R1399 B.n531 B.n140 10.6151
R1400 B.n531 B.n530 10.6151
R1401 B.n530 B.n529 10.6151
R1402 B.n529 B.n142 10.6151
R1403 B.n525 B.n142 10.6151
R1404 B.n525 B.n524 10.6151
R1405 B.n524 B.n523 10.6151
R1406 B.n523 B.n144 10.6151
R1407 B.n519 B.n144 10.6151
R1408 B.n519 B.n518 10.6151
R1409 B.n518 B.n517 10.6151
R1410 B.n517 B.n146 10.6151
R1411 B.n513 B.n146 10.6151
R1412 B.n513 B.n512 10.6151
R1413 B.n512 B.n511 10.6151
R1414 B.n239 B.n1 10.6151
R1415 B.n239 B.n238 10.6151
R1416 B.n243 B.n238 10.6151
R1417 B.n244 B.n243 10.6151
R1418 B.n245 B.n244 10.6151
R1419 B.n245 B.n236 10.6151
R1420 B.n249 B.n236 10.6151
R1421 B.n250 B.n249 10.6151
R1422 B.n251 B.n250 10.6151
R1423 B.n251 B.n234 10.6151
R1424 B.n255 B.n234 10.6151
R1425 B.n256 B.n255 10.6151
R1426 B.n257 B.n256 10.6151
R1427 B.n257 B.n232 10.6151
R1428 B.n261 B.n232 10.6151
R1429 B.n262 B.n261 10.6151
R1430 B.n263 B.n262 10.6151
R1431 B.n263 B.n230 10.6151
R1432 B.n267 B.n230 10.6151
R1433 B.n268 B.n267 10.6151
R1434 B.n269 B.n268 10.6151
R1435 B.n269 B.n228 10.6151
R1436 B.n273 B.n228 10.6151
R1437 B.n274 B.n273 10.6151
R1438 B.n275 B.n274 10.6151
R1439 B.n275 B.n226 10.6151
R1440 B.n279 B.n226 10.6151
R1441 B.n280 B.n279 10.6151
R1442 B.n281 B.n280 10.6151
R1443 B.n281 B.n224 10.6151
R1444 B.n285 B.n224 10.6151
R1445 B.n286 B.n285 10.6151
R1446 B.n287 B.n286 10.6151
R1447 B.n287 B.n222 10.6151
R1448 B.n291 B.n222 10.6151
R1449 B.n292 B.n291 10.6151
R1450 B.n293 B.n292 10.6151
R1451 B.n293 B.n220 10.6151
R1452 B.n297 B.n220 10.6151
R1453 B.n298 B.n297 10.6151
R1454 B.n299 B.n298 10.6151
R1455 B.n299 B.n218 10.6151
R1456 B.n303 B.n218 10.6151
R1457 B.n304 B.n303 10.6151
R1458 B.n305 B.n304 10.6151
R1459 B.n305 B.n216 10.6151
R1460 B.n309 B.n216 10.6151
R1461 B.n310 B.n309 10.6151
R1462 B.n311 B.n310 10.6151
R1463 B.n311 B.n214 10.6151
R1464 B.n316 B.n315 10.6151
R1465 B.n317 B.n316 10.6151
R1466 B.n317 B.n212 10.6151
R1467 B.n321 B.n212 10.6151
R1468 B.n322 B.n321 10.6151
R1469 B.n323 B.n322 10.6151
R1470 B.n323 B.n210 10.6151
R1471 B.n327 B.n210 10.6151
R1472 B.n328 B.n327 10.6151
R1473 B.n329 B.n328 10.6151
R1474 B.n329 B.n208 10.6151
R1475 B.n333 B.n208 10.6151
R1476 B.n334 B.n333 10.6151
R1477 B.n335 B.n334 10.6151
R1478 B.n335 B.n206 10.6151
R1479 B.n339 B.n206 10.6151
R1480 B.n340 B.n339 10.6151
R1481 B.n341 B.n340 10.6151
R1482 B.n341 B.n204 10.6151
R1483 B.n345 B.n204 10.6151
R1484 B.n346 B.n345 10.6151
R1485 B.n347 B.n346 10.6151
R1486 B.n347 B.n202 10.6151
R1487 B.n351 B.n202 10.6151
R1488 B.n352 B.n351 10.6151
R1489 B.n353 B.n352 10.6151
R1490 B.n353 B.n200 10.6151
R1491 B.n357 B.n200 10.6151
R1492 B.n358 B.n357 10.6151
R1493 B.n359 B.n358 10.6151
R1494 B.n359 B.n198 10.6151
R1495 B.n363 B.n198 10.6151
R1496 B.n364 B.n363 10.6151
R1497 B.n365 B.n364 10.6151
R1498 B.n365 B.n196 10.6151
R1499 B.n369 B.n196 10.6151
R1500 B.n370 B.n369 10.6151
R1501 B.n371 B.n370 10.6151
R1502 B.n371 B.n194 10.6151
R1503 B.n375 B.n194 10.6151
R1504 B.n376 B.n375 10.6151
R1505 B.n377 B.n376 10.6151
R1506 B.n377 B.n192 10.6151
R1507 B.n381 B.n192 10.6151
R1508 B.n382 B.n381 10.6151
R1509 B.n383 B.n382 10.6151
R1510 B.n383 B.n190 10.6151
R1511 B.n387 B.n190 10.6151
R1512 B.n388 B.n387 10.6151
R1513 B.n389 B.n388 10.6151
R1514 B.n389 B.n188 10.6151
R1515 B.n393 B.n188 10.6151
R1516 B.n394 B.n393 10.6151
R1517 B.n395 B.n394 10.6151
R1518 B.n395 B.n186 10.6151
R1519 B.n399 B.n186 10.6151
R1520 B.n400 B.n399 10.6151
R1521 B.n404 B.n400 10.6151
R1522 B.n408 B.n184 10.6151
R1523 B.n409 B.n408 10.6151
R1524 B.n410 B.n409 10.6151
R1525 B.n410 B.n182 10.6151
R1526 B.n414 B.n182 10.6151
R1527 B.n415 B.n414 10.6151
R1528 B.n416 B.n415 10.6151
R1529 B.n416 B.n180 10.6151
R1530 B.n420 B.n180 10.6151
R1531 B.n423 B.n422 10.6151
R1532 B.n423 B.n176 10.6151
R1533 B.n427 B.n176 10.6151
R1534 B.n428 B.n427 10.6151
R1535 B.n429 B.n428 10.6151
R1536 B.n429 B.n174 10.6151
R1537 B.n433 B.n174 10.6151
R1538 B.n434 B.n433 10.6151
R1539 B.n435 B.n434 10.6151
R1540 B.n435 B.n172 10.6151
R1541 B.n439 B.n172 10.6151
R1542 B.n440 B.n439 10.6151
R1543 B.n441 B.n440 10.6151
R1544 B.n441 B.n170 10.6151
R1545 B.n445 B.n170 10.6151
R1546 B.n446 B.n445 10.6151
R1547 B.n447 B.n446 10.6151
R1548 B.n447 B.n168 10.6151
R1549 B.n451 B.n168 10.6151
R1550 B.n452 B.n451 10.6151
R1551 B.n453 B.n452 10.6151
R1552 B.n453 B.n166 10.6151
R1553 B.n457 B.n166 10.6151
R1554 B.n458 B.n457 10.6151
R1555 B.n459 B.n458 10.6151
R1556 B.n459 B.n164 10.6151
R1557 B.n463 B.n164 10.6151
R1558 B.n464 B.n463 10.6151
R1559 B.n465 B.n464 10.6151
R1560 B.n465 B.n162 10.6151
R1561 B.n469 B.n162 10.6151
R1562 B.n470 B.n469 10.6151
R1563 B.n471 B.n470 10.6151
R1564 B.n471 B.n160 10.6151
R1565 B.n475 B.n160 10.6151
R1566 B.n476 B.n475 10.6151
R1567 B.n477 B.n476 10.6151
R1568 B.n477 B.n158 10.6151
R1569 B.n481 B.n158 10.6151
R1570 B.n482 B.n481 10.6151
R1571 B.n483 B.n482 10.6151
R1572 B.n483 B.n156 10.6151
R1573 B.n487 B.n156 10.6151
R1574 B.n488 B.n487 10.6151
R1575 B.n489 B.n488 10.6151
R1576 B.n489 B.n154 10.6151
R1577 B.n493 B.n154 10.6151
R1578 B.n494 B.n493 10.6151
R1579 B.n495 B.n494 10.6151
R1580 B.n495 B.n152 10.6151
R1581 B.n499 B.n152 10.6151
R1582 B.n500 B.n499 10.6151
R1583 B.n501 B.n500 10.6151
R1584 B.n501 B.n150 10.6151
R1585 B.n505 B.n150 10.6151
R1586 B.n506 B.n505 10.6151
R1587 B.n507 B.n506 10.6151
R1588 B.n507 B.n148 10.6151
R1589 B.n771 B.n770 9.36635
R1590 B.n753 B.n66 9.36635
R1591 B.n404 B.n403 9.36635
R1592 B.n422 B.n421 9.36635
R1593 B.n937 B.n0 8.11757
R1594 B.n937 B.n1 8.11757
R1595 B.n770 B.n769 1.24928
R1596 B.n756 B.n66 1.24928
R1597 B.n403 B.n184 1.24928
R1598 B.n421 B.n420 1.24928
C0 B VDD2 2.85981f
C1 VDD1 B 2.76773f
C2 VTAIL VP 10.3894f
C3 VTAIL VDD2 9.9906f
C4 VTAIL VDD1 9.93514f
C5 VTAIL B 5.37815f
C6 VN w_n3914_n4562# 7.715089f
C7 VP w_n3914_n4562# 8.22321f
C8 VDD2 w_n3914_n4562# 2.9933f
C9 VDD1 w_n3914_n4562# 2.88426f
C10 VN VP 8.7653f
C11 B w_n3914_n4562# 12.3857f
C12 VN VDD2 10.3141f
C13 VN VDD1 0.151839f
C14 VTAIL w_n3914_n4562# 3.85567f
C15 VN B 1.39557f
C16 VP VDD2 0.522379f
C17 VDD1 VP 10.6807f
C18 B VP 2.2477f
C19 VN VTAIL 10.3751f
C20 VDD1 VDD2 1.70061f
C21 VDD2 VSUBS 2.25718f
C22 VDD1 VSUBS 2.81423f
C23 VTAIL VSUBS 1.550598f
C24 VN VSUBS 6.78622f
C25 VP VSUBS 3.736527f
C26 B VSUBS 5.882811f
C27 w_n3914_n4562# VSUBS 0.218354p
C28 B.n0 VSUBS 0.006519f
C29 B.n1 VSUBS 0.006519f
C30 B.n2 VSUBS 0.009641f
C31 B.n3 VSUBS 0.007388f
C32 B.n4 VSUBS 0.007388f
C33 B.n5 VSUBS 0.007388f
C34 B.n6 VSUBS 0.007388f
C35 B.n7 VSUBS 0.007388f
C36 B.n8 VSUBS 0.007388f
C37 B.n9 VSUBS 0.007388f
C38 B.n10 VSUBS 0.007388f
C39 B.n11 VSUBS 0.007388f
C40 B.n12 VSUBS 0.007388f
C41 B.n13 VSUBS 0.007388f
C42 B.n14 VSUBS 0.007388f
C43 B.n15 VSUBS 0.007388f
C44 B.n16 VSUBS 0.007388f
C45 B.n17 VSUBS 0.007388f
C46 B.n18 VSUBS 0.007388f
C47 B.n19 VSUBS 0.007388f
C48 B.n20 VSUBS 0.007388f
C49 B.n21 VSUBS 0.007388f
C50 B.n22 VSUBS 0.007388f
C51 B.n23 VSUBS 0.007388f
C52 B.n24 VSUBS 0.007388f
C53 B.n25 VSUBS 0.007388f
C54 B.n26 VSUBS 0.007388f
C55 B.n27 VSUBS 0.016339f
C56 B.n28 VSUBS 0.007388f
C57 B.n29 VSUBS 0.007388f
C58 B.n30 VSUBS 0.007388f
C59 B.n31 VSUBS 0.007388f
C60 B.n32 VSUBS 0.007388f
C61 B.n33 VSUBS 0.007388f
C62 B.n34 VSUBS 0.007388f
C63 B.n35 VSUBS 0.007388f
C64 B.n36 VSUBS 0.007388f
C65 B.n37 VSUBS 0.007388f
C66 B.n38 VSUBS 0.007388f
C67 B.n39 VSUBS 0.007388f
C68 B.n40 VSUBS 0.007388f
C69 B.n41 VSUBS 0.007388f
C70 B.n42 VSUBS 0.007388f
C71 B.n43 VSUBS 0.007388f
C72 B.n44 VSUBS 0.007388f
C73 B.n45 VSUBS 0.007388f
C74 B.n46 VSUBS 0.007388f
C75 B.n47 VSUBS 0.007388f
C76 B.n48 VSUBS 0.007388f
C77 B.n49 VSUBS 0.007388f
C78 B.n50 VSUBS 0.007388f
C79 B.n51 VSUBS 0.007388f
C80 B.n52 VSUBS 0.007388f
C81 B.n53 VSUBS 0.007388f
C82 B.n54 VSUBS 0.007388f
C83 B.n55 VSUBS 0.007388f
C84 B.n56 VSUBS 0.007388f
C85 B.n57 VSUBS 0.007388f
C86 B.t7 VSUBS 0.640214f
C87 B.t8 VSUBS 0.66703f
C88 B.t6 VSUBS 2.87062f
C89 B.n58 VSUBS 0.399712f
C90 B.n59 VSUBS 0.079362f
C91 B.n60 VSUBS 0.007388f
C92 B.n61 VSUBS 0.007388f
C93 B.n62 VSUBS 0.007388f
C94 B.n63 VSUBS 0.007388f
C95 B.t10 VSUBS 0.640191f
C96 B.t11 VSUBS 0.667013f
C97 B.t9 VSUBS 2.87062f
C98 B.n64 VSUBS 0.39973f
C99 B.n65 VSUBS 0.079385f
C100 B.n66 VSUBS 0.017117f
C101 B.n67 VSUBS 0.007388f
C102 B.n68 VSUBS 0.007388f
C103 B.n69 VSUBS 0.007388f
C104 B.n70 VSUBS 0.007388f
C105 B.n71 VSUBS 0.007388f
C106 B.n72 VSUBS 0.007388f
C107 B.n73 VSUBS 0.007388f
C108 B.n74 VSUBS 0.007388f
C109 B.n75 VSUBS 0.007388f
C110 B.n76 VSUBS 0.007388f
C111 B.n77 VSUBS 0.007388f
C112 B.n78 VSUBS 0.007388f
C113 B.n79 VSUBS 0.007388f
C114 B.n80 VSUBS 0.007388f
C115 B.n81 VSUBS 0.007388f
C116 B.n82 VSUBS 0.007388f
C117 B.n83 VSUBS 0.007388f
C118 B.n84 VSUBS 0.007388f
C119 B.n85 VSUBS 0.007388f
C120 B.n86 VSUBS 0.007388f
C121 B.n87 VSUBS 0.007388f
C122 B.n88 VSUBS 0.007388f
C123 B.n89 VSUBS 0.007388f
C124 B.n90 VSUBS 0.007388f
C125 B.n91 VSUBS 0.007388f
C126 B.n92 VSUBS 0.007388f
C127 B.n93 VSUBS 0.007388f
C128 B.n94 VSUBS 0.007388f
C129 B.n95 VSUBS 0.007388f
C130 B.n96 VSUBS 0.016339f
C131 B.n97 VSUBS 0.007388f
C132 B.n98 VSUBS 0.007388f
C133 B.n99 VSUBS 0.007388f
C134 B.n100 VSUBS 0.007388f
C135 B.n101 VSUBS 0.007388f
C136 B.n102 VSUBS 0.007388f
C137 B.n103 VSUBS 0.007388f
C138 B.n104 VSUBS 0.007388f
C139 B.n105 VSUBS 0.007388f
C140 B.n106 VSUBS 0.007388f
C141 B.n107 VSUBS 0.007388f
C142 B.n108 VSUBS 0.007388f
C143 B.n109 VSUBS 0.007388f
C144 B.n110 VSUBS 0.007388f
C145 B.n111 VSUBS 0.007388f
C146 B.n112 VSUBS 0.007388f
C147 B.n113 VSUBS 0.007388f
C148 B.n114 VSUBS 0.007388f
C149 B.n115 VSUBS 0.007388f
C150 B.n116 VSUBS 0.007388f
C151 B.n117 VSUBS 0.007388f
C152 B.n118 VSUBS 0.007388f
C153 B.n119 VSUBS 0.007388f
C154 B.n120 VSUBS 0.007388f
C155 B.n121 VSUBS 0.007388f
C156 B.n122 VSUBS 0.007388f
C157 B.n123 VSUBS 0.007388f
C158 B.n124 VSUBS 0.007388f
C159 B.n125 VSUBS 0.007388f
C160 B.n126 VSUBS 0.007388f
C161 B.n127 VSUBS 0.007388f
C162 B.n128 VSUBS 0.007388f
C163 B.n129 VSUBS 0.007388f
C164 B.n130 VSUBS 0.007388f
C165 B.n131 VSUBS 0.007388f
C166 B.n132 VSUBS 0.007388f
C167 B.n133 VSUBS 0.007388f
C168 B.n134 VSUBS 0.007388f
C169 B.n135 VSUBS 0.007388f
C170 B.n136 VSUBS 0.007388f
C171 B.n137 VSUBS 0.007388f
C172 B.n138 VSUBS 0.007388f
C173 B.n139 VSUBS 0.007388f
C174 B.n140 VSUBS 0.007388f
C175 B.n141 VSUBS 0.007388f
C176 B.n142 VSUBS 0.007388f
C177 B.n143 VSUBS 0.007388f
C178 B.n144 VSUBS 0.007388f
C179 B.n145 VSUBS 0.007388f
C180 B.n146 VSUBS 0.007388f
C181 B.n147 VSUBS 0.007388f
C182 B.n148 VSUBS 0.016205f
C183 B.n149 VSUBS 0.007388f
C184 B.n150 VSUBS 0.007388f
C185 B.n151 VSUBS 0.007388f
C186 B.n152 VSUBS 0.007388f
C187 B.n153 VSUBS 0.007388f
C188 B.n154 VSUBS 0.007388f
C189 B.n155 VSUBS 0.007388f
C190 B.n156 VSUBS 0.007388f
C191 B.n157 VSUBS 0.007388f
C192 B.n158 VSUBS 0.007388f
C193 B.n159 VSUBS 0.007388f
C194 B.n160 VSUBS 0.007388f
C195 B.n161 VSUBS 0.007388f
C196 B.n162 VSUBS 0.007388f
C197 B.n163 VSUBS 0.007388f
C198 B.n164 VSUBS 0.007388f
C199 B.n165 VSUBS 0.007388f
C200 B.n166 VSUBS 0.007388f
C201 B.n167 VSUBS 0.007388f
C202 B.n168 VSUBS 0.007388f
C203 B.n169 VSUBS 0.007388f
C204 B.n170 VSUBS 0.007388f
C205 B.n171 VSUBS 0.007388f
C206 B.n172 VSUBS 0.007388f
C207 B.n173 VSUBS 0.007388f
C208 B.n174 VSUBS 0.007388f
C209 B.n175 VSUBS 0.007388f
C210 B.n176 VSUBS 0.007388f
C211 B.n177 VSUBS 0.007388f
C212 B.t5 VSUBS 0.640191f
C213 B.t4 VSUBS 0.667013f
C214 B.t3 VSUBS 2.87062f
C215 B.n178 VSUBS 0.39973f
C216 B.n179 VSUBS 0.079385f
C217 B.n180 VSUBS 0.007388f
C218 B.n181 VSUBS 0.007388f
C219 B.n182 VSUBS 0.007388f
C220 B.n183 VSUBS 0.007388f
C221 B.n184 VSUBS 0.004128f
C222 B.n185 VSUBS 0.007388f
C223 B.n186 VSUBS 0.007388f
C224 B.n187 VSUBS 0.007388f
C225 B.n188 VSUBS 0.007388f
C226 B.n189 VSUBS 0.007388f
C227 B.n190 VSUBS 0.007388f
C228 B.n191 VSUBS 0.007388f
C229 B.n192 VSUBS 0.007388f
C230 B.n193 VSUBS 0.007388f
C231 B.n194 VSUBS 0.007388f
C232 B.n195 VSUBS 0.007388f
C233 B.n196 VSUBS 0.007388f
C234 B.n197 VSUBS 0.007388f
C235 B.n198 VSUBS 0.007388f
C236 B.n199 VSUBS 0.007388f
C237 B.n200 VSUBS 0.007388f
C238 B.n201 VSUBS 0.007388f
C239 B.n202 VSUBS 0.007388f
C240 B.n203 VSUBS 0.007388f
C241 B.n204 VSUBS 0.007388f
C242 B.n205 VSUBS 0.007388f
C243 B.n206 VSUBS 0.007388f
C244 B.n207 VSUBS 0.007388f
C245 B.n208 VSUBS 0.007388f
C246 B.n209 VSUBS 0.007388f
C247 B.n210 VSUBS 0.007388f
C248 B.n211 VSUBS 0.007388f
C249 B.n212 VSUBS 0.007388f
C250 B.n213 VSUBS 0.007388f
C251 B.n214 VSUBS 0.016339f
C252 B.n215 VSUBS 0.007388f
C253 B.n216 VSUBS 0.007388f
C254 B.n217 VSUBS 0.007388f
C255 B.n218 VSUBS 0.007388f
C256 B.n219 VSUBS 0.007388f
C257 B.n220 VSUBS 0.007388f
C258 B.n221 VSUBS 0.007388f
C259 B.n222 VSUBS 0.007388f
C260 B.n223 VSUBS 0.007388f
C261 B.n224 VSUBS 0.007388f
C262 B.n225 VSUBS 0.007388f
C263 B.n226 VSUBS 0.007388f
C264 B.n227 VSUBS 0.007388f
C265 B.n228 VSUBS 0.007388f
C266 B.n229 VSUBS 0.007388f
C267 B.n230 VSUBS 0.007388f
C268 B.n231 VSUBS 0.007388f
C269 B.n232 VSUBS 0.007388f
C270 B.n233 VSUBS 0.007388f
C271 B.n234 VSUBS 0.007388f
C272 B.n235 VSUBS 0.007388f
C273 B.n236 VSUBS 0.007388f
C274 B.n237 VSUBS 0.007388f
C275 B.n238 VSUBS 0.007388f
C276 B.n239 VSUBS 0.007388f
C277 B.n240 VSUBS 0.007388f
C278 B.n241 VSUBS 0.007388f
C279 B.n242 VSUBS 0.007388f
C280 B.n243 VSUBS 0.007388f
C281 B.n244 VSUBS 0.007388f
C282 B.n245 VSUBS 0.007388f
C283 B.n246 VSUBS 0.007388f
C284 B.n247 VSUBS 0.007388f
C285 B.n248 VSUBS 0.007388f
C286 B.n249 VSUBS 0.007388f
C287 B.n250 VSUBS 0.007388f
C288 B.n251 VSUBS 0.007388f
C289 B.n252 VSUBS 0.007388f
C290 B.n253 VSUBS 0.007388f
C291 B.n254 VSUBS 0.007388f
C292 B.n255 VSUBS 0.007388f
C293 B.n256 VSUBS 0.007388f
C294 B.n257 VSUBS 0.007388f
C295 B.n258 VSUBS 0.007388f
C296 B.n259 VSUBS 0.007388f
C297 B.n260 VSUBS 0.007388f
C298 B.n261 VSUBS 0.007388f
C299 B.n262 VSUBS 0.007388f
C300 B.n263 VSUBS 0.007388f
C301 B.n264 VSUBS 0.007388f
C302 B.n265 VSUBS 0.007388f
C303 B.n266 VSUBS 0.007388f
C304 B.n267 VSUBS 0.007388f
C305 B.n268 VSUBS 0.007388f
C306 B.n269 VSUBS 0.007388f
C307 B.n270 VSUBS 0.007388f
C308 B.n271 VSUBS 0.007388f
C309 B.n272 VSUBS 0.007388f
C310 B.n273 VSUBS 0.007388f
C311 B.n274 VSUBS 0.007388f
C312 B.n275 VSUBS 0.007388f
C313 B.n276 VSUBS 0.007388f
C314 B.n277 VSUBS 0.007388f
C315 B.n278 VSUBS 0.007388f
C316 B.n279 VSUBS 0.007388f
C317 B.n280 VSUBS 0.007388f
C318 B.n281 VSUBS 0.007388f
C319 B.n282 VSUBS 0.007388f
C320 B.n283 VSUBS 0.007388f
C321 B.n284 VSUBS 0.007388f
C322 B.n285 VSUBS 0.007388f
C323 B.n286 VSUBS 0.007388f
C324 B.n287 VSUBS 0.007388f
C325 B.n288 VSUBS 0.007388f
C326 B.n289 VSUBS 0.007388f
C327 B.n290 VSUBS 0.007388f
C328 B.n291 VSUBS 0.007388f
C329 B.n292 VSUBS 0.007388f
C330 B.n293 VSUBS 0.007388f
C331 B.n294 VSUBS 0.007388f
C332 B.n295 VSUBS 0.007388f
C333 B.n296 VSUBS 0.007388f
C334 B.n297 VSUBS 0.007388f
C335 B.n298 VSUBS 0.007388f
C336 B.n299 VSUBS 0.007388f
C337 B.n300 VSUBS 0.007388f
C338 B.n301 VSUBS 0.007388f
C339 B.n302 VSUBS 0.007388f
C340 B.n303 VSUBS 0.007388f
C341 B.n304 VSUBS 0.007388f
C342 B.n305 VSUBS 0.007388f
C343 B.n306 VSUBS 0.007388f
C344 B.n307 VSUBS 0.007388f
C345 B.n308 VSUBS 0.007388f
C346 B.n309 VSUBS 0.007388f
C347 B.n310 VSUBS 0.007388f
C348 B.n311 VSUBS 0.007388f
C349 B.n312 VSUBS 0.007388f
C350 B.n313 VSUBS 0.016339f
C351 B.n314 VSUBS 0.017123f
C352 B.n315 VSUBS 0.017123f
C353 B.n316 VSUBS 0.007388f
C354 B.n317 VSUBS 0.007388f
C355 B.n318 VSUBS 0.007388f
C356 B.n319 VSUBS 0.007388f
C357 B.n320 VSUBS 0.007388f
C358 B.n321 VSUBS 0.007388f
C359 B.n322 VSUBS 0.007388f
C360 B.n323 VSUBS 0.007388f
C361 B.n324 VSUBS 0.007388f
C362 B.n325 VSUBS 0.007388f
C363 B.n326 VSUBS 0.007388f
C364 B.n327 VSUBS 0.007388f
C365 B.n328 VSUBS 0.007388f
C366 B.n329 VSUBS 0.007388f
C367 B.n330 VSUBS 0.007388f
C368 B.n331 VSUBS 0.007388f
C369 B.n332 VSUBS 0.007388f
C370 B.n333 VSUBS 0.007388f
C371 B.n334 VSUBS 0.007388f
C372 B.n335 VSUBS 0.007388f
C373 B.n336 VSUBS 0.007388f
C374 B.n337 VSUBS 0.007388f
C375 B.n338 VSUBS 0.007388f
C376 B.n339 VSUBS 0.007388f
C377 B.n340 VSUBS 0.007388f
C378 B.n341 VSUBS 0.007388f
C379 B.n342 VSUBS 0.007388f
C380 B.n343 VSUBS 0.007388f
C381 B.n344 VSUBS 0.007388f
C382 B.n345 VSUBS 0.007388f
C383 B.n346 VSUBS 0.007388f
C384 B.n347 VSUBS 0.007388f
C385 B.n348 VSUBS 0.007388f
C386 B.n349 VSUBS 0.007388f
C387 B.n350 VSUBS 0.007388f
C388 B.n351 VSUBS 0.007388f
C389 B.n352 VSUBS 0.007388f
C390 B.n353 VSUBS 0.007388f
C391 B.n354 VSUBS 0.007388f
C392 B.n355 VSUBS 0.007388f
C393 B.n356 VSUBS 0.007388f
C394 B.n357 VSUBS 0.007388f
C395 B.n358 VSUBS 0.007388f
C396 B.n359 VSUBS 0.007388f
C397 B.n360 VSUBS 0.007388f
C398 B.n361 VSUBS 0.007388f
C399 B.n362 VSUBS 0.007388f
C400 B.n363 VSUBS 0.007388f
C401 B.n364 VSUBS 0.007388f
C402 B.n365 VSUBS 0.007388f
C403 B.n366 VSUBS 0.007388f
C404 B.n367 VSUBS 0.007388f
C405 B.n368 VSUBS 0.007388f
C406 B.n369 VSUBS 0.007388f
C407 B.n370 VSUBS 0.007388f
C408 B.n371 VSUBS 0.007388f
C409 B.n372 VSUBS 0.007388f
C410 B.n373 VSUBS 0.007388f
C411 B.n374 VSUBS 0.007388f
C412 B.n375 VSUBS 0.007388f
C413 B.n376 VSUBS 0.007388f
C414 B.n377 VSUBS 0.007388f
C415 B.n378 VSUBS 0.007388f
C416 B.n379 VSUBS 0.007388f
C417 B.n380 VSUBS 0.007388f
C418 B.n381 VSUBS 0.007388f
C419 B.n382 VSUBS 0.007388f
C420 B.n383 VSUBS 0.007388f
C421 B.n384 VSUBS 0.007388f
C422 B.n385 VSUBS 0.007388f
C423 B.n386 VSUBS 0.007388f
C424 B.n387 VSUBS 0.007388f
C425 B.n388 VSUBS 0.007388f
C426 B.n389 VSUBS 0.007388f
C427 B.n390 VSUBS 0.007388f
C428 B.n391 VSUBS 0.007388f
C429 B.n392 VSUBS 0.007388f
C430 B.n393 VSUBS 0.007388f
C431 B.n394 VSUBS 0.007388f
C432 B.n395 VSUBS 0.007388f
C433 B.n396 VSUBS 0.007388f
C434 B.n397 VSUBS 0.007388f
C435 B.n398 VSUBS 0.007388f
C436 B.n399 VSUBS 0.007388f
C437 B.n400 VSUBS 0.007388f
C438 B.t2 VSUBS 0.640214f
C439 B.t1 VSUBS 0.66703f
C440 B.t0 VSUBS 2.87062f
C441 B.n401 VSUBS 0.399712f
C442 B.n402 VSUBS 0.079362f
C443 B.n403 VSUBS 0.017117f
C444 B.n404 VSUBS 0.006953f
C445 B.n405 VSUBS 0.007388f
C446 B.n406 VSUBS 0.007388f
C447 B.n407 VSUBS 0.007388f
C448 B.n408 VSUBS 0.007388f
C449 B.n409 VSUBS 0.007388f
C450 B.n410 VSUBS 0.007388f
C451 B.n411 VSUBS 0.007388f
C452 B.n412 VSUBS 0.007388f
C453 B.n413 VSUBS 0.007388f
C454 B.n414 VSUBS 0.007388f
C455 B.n415 VSUBS 0.007388f
C456 B.n416 VSUBS 0.007388f
C457 B.n417 VSUBS 0.007388f
C458 B.n418 VSUBS 0.007388f
C459 B.n419 VSUBS 0.007388f
C460 B.n420 VSUBS 0.004128f
C461 B.n421 VSUBS 0.017117f
C462 B.n422 VSUBS 0.006953f
C463 B.n423 VSUBS 0.007388f
C464 B.n424 VSUBS 0.007388f
C465 B.n425 VSUBS 0.007388f
C466 B.n426 VSUBS 0.007388f
C467 B.n427 VSUBS 0.007388f
C468 B.n428 VSUBS 0.007388f
C469 B.n429 VSUBS 0.007388f
C470 B.n430 VSUBS 0.007388f
C471 B.n431 VSUBS 0.007388f
C472 B.n432 VSUBS 0.007388f
C473 B.n433 VSUBS 0.007388f
C474 B.n434 VSUBS 0.007388f
C475 B.n435 VSUBS 0.007388f
C476 B.n436 VSUBS 0.007388f
C477 B.n437 VSUBS 0.007388f
C478 B.n438 VSUBS 0.007388f
C479 B.n439 VSUBS 0.007388f
C480 B.n440 VSUBS 0.007388f
C481 B.n441 VSUBS 0.007388f
C482 B.n442 VSUBS 0.007388f
C483 B.n443 VSUBS 0.007388f
C484 B.n444 VSUBS 0.007388f
C485 B.n445 VSUBS 0.007388f
C486 B.n446 VSUBS 0.007388f
C487 B.n447 VSUBS 0.007388f
C488 B.n448 VSUBS 0.007388f
C489 B.n449 VSUBS 0.007388f
C490 B.n450 VSUBS 0.007388f
C491 B.n451 VSUBS 0.007388f
C492 B.n452 VSUBS 0.007388f
C493 B.n453 VSUBS 0.007388f
C494 B.n454 VSUBS 0.007388f
C495 B.n455 VSUBS 0.007388f
C496 B.n456 VSUBS 0.007388f
C497 B.n457 VSUBS 0.007388f
C498 B.n458 VSUBS 0.007388f
C499 B.n459 VSUBS 0.007388f
C500 B.n460 VSUBS 0.007388f
C501 B.n461 VSUBS 0.007388f
C502 B.n462 VSUBS 0.007388f
C503 B.n463 VSUBS 0.007388f
C504 B.n464 VSUBS 0.007388f
C505 B.n465 VSUBS 0.007388f
C506 B.n466 VSUBS 0.007388f
C507 B.n467 VSUBS 0.007388f
C508 B.n468 VSUBS 0.007388f
C509 B.n469 VSUBS 0.007388f
C510 B.n470 VSUBS 0.007388f
C511 B.n471 VSUBS 0.007388f
C512 B.n472 VSUBS 0.007388f
C513 B.n473 VSUBS 0.007388f
C514 B.n474 VSUBS 0.007388f
C515 B.n475 VSUBS 0.007388f
C516 B.n476 VSUBS 0.007388f
C517 B.n477 VSUBS 0.007388f
C518 B.n478 VSUBS 0.007388f
C519 B.n479 VSUBS 0.007388f
C520 B.n480 VSUBS 0.007388f
C521 B.n481 VSUBS 0.007388f
C522 B.n482 VSUBS 0.007388f
C523 B.n483 VSUBS 0.007388f
C524 B.n484 VSUBS 0.007388f
C525 B.n485 VSUBS 0.007388f
C526 B.n486 VSUBS 0.007388f
C527 B.n487 VSUBS 0.007388f
C528 B.n488 VSUBS 0.007388f
C529 B.n489 VSUBS 0.007388f
C530 B.n490 VSUBS 0.007388f
C531 B.n491 VSUBS 0.007388f
C532 B.n492 VSUBS 0.007388f
C533 B.n493 VSUBS 0.007388f
C534 B.n494 VSUBS 0.007388f
C535 B.n495 VSUBS 0.007388f
C536 B.n496 VSUBS 0.007388f
C537 B.n497 VSUBS 0.007388f
C538 B.n498 VSUBS 0.007388f
C539 B.n499 VSUBS 0.007388f
C540 B.n500 VSUBS 0.007388f
C541 B.n501 VSUBS 0.007388f
C542 B.n502 VSUBS 0.007388f
C543 B.n503 VSUBS 0.007388f
C544 B.n504 VSUBS 0.007388f
C545 B.n505 VSUBS 0.007388f
C546 B.n506 VSUBS 0.007388f
C547 B.n507 VSUBS 0.007388f
C548 B.n508 VSUBS 0.007388f
C549 B.n509 VSUBS 0.017123f
C550 B.n510 VSUBS 0.016339f
C551 B.n511 VSUBS 0.017257f
C552 B.n512 VSUBS 0.007388f
C553 B.n513 VSUBS 0.007388f
C554 B.n514 VSUBS 0.007388f
C555 B.n515 VSUBS 0.007388f
C556 B.n516 VSUBS 0.007388f
C557 B.n517 VSUBS 0.007388f
C558 B.n518 VSUBS 0.007388f
C559 B.n519 VSUBS 0.007388f
C560 B.n520 VSUBS 0.007388f
C561 B.n521 VSUBS 0.007388f
C562 B.n522 VSUBS 0.007388f
C563 B.n523 VSUBS 0.007388f
C564 B.n524 VSUBS 0.007388f
C565 B.n525 VSUBS 0.007388f
C566 B.n526 VSUBS 0.007388f
C567 B.n527 VSUBS 0.007388f
C568 B.n528 VSUBS 0.007388f
C569 B.n529 VSUBS 0.007388f
C570 B.n530 VSUBS 0.007388f
C571 B.n531 VSUBS 0.007388f
C572 B.n532 VSUBS 0.007388f
C573 B.n533 VSUBS 0.007388f
C574 B.n534 VSUBS 0.007388f
C575 B.n535 VSUBS 0.007388f
C576 B.n536 VSUBS 0.007388f
C577 B.n537 VSUBS 0.007388f
C578 B.n538 VSUBS 0.007388f
C579 B.n539 VSUBS 0.007388f
C580 B.n540 VSUBS 0.007388f
C581 B.n541 VSUBS 0.007388f
C582 B.n542 VSUBS 0.007388f
C583 B.n543 VSUBS 0.007388f
C584 B.n544 VSUBS 0.007388f
C585 B.n545 VSUBS 0.007388f
C586 B.n546 VSUBS 0.007388f
C587 B.n547 VSUBS 0.007388f
C588 B.n548 VSUBS 0.007388f
C589 B.n549 VSUBS 0.007388f
C590 B.n550 VSUBS 0.007388f
C591 B.n551 VSUBS 0.007388f
C592 B.n552 VSUBS 0.007388f
C593 B.n553 VSUBS 0.007388f
C594 B.n554 VSUBS 0.007388f
C595 B.n555 VSUBS 0.007388f
C596 B.n556 VSUBS 0.007388f
C597 B.n557 VSUBS 0.007388f
C598 B.n558 VSUBS 0.007388f
C599 B.n559 VSUBS 0.007388f
C600 B.n560 VSUBS 0.007388f
C601 B.n561 VSUBS 0.007388f
C602 B.n562 VSUBS 0.007388f
C603 B.n563 VSUBS 0.007388f
C604 B.n564 VSUBS 0.007388f
C605 B.n565 VSUBS 0.007388f
C606 B.n566 VSUBS 0.007388f
C607 B.n567 VSUBS 0.007388f
C608 B.n568 VSUBS 0.007388f
C609 B.n569 VSUBS 0.007388f
C610 B.n570 VSUBS 0.007388f
C611 B.n571 VSUBS 0.007388f
C612 B.n572 VSUBS 0.007388f
C613 B.n573 VSUBS 0.007388f
C614 B.n574 VSUBS 0.007388f
C615 B.n575 VSUBS 0.007388f
C616 B.n576 VSUBS 0.007388f
C617 B.n577 VSUBS 0.007388f
C618 B.n578 VSUBS 0.007388f
C619 B.n579 VSUBS 0.007388f
C620 B.n580 VSUBS 0.007388f
C621 B.n581 VSUBS 0.007388f
C622 B.n582 VSUBS 0.007388f
C623 B.n583 VSUBS 0.007388f
C624 B.n584 VSUBS 0.007388f
C625 B.n585 VSUBS 0.007388f
C626 B.n586 VSUBS 0.007388f
C627 B.n587 VSUBS 0.007388f
C628 B.n588 VSUBS 0.007388f
C629 B.n589 VSUBS 0.007388f
C630 B.n590 VSUBS 0.007388f
C631 B.n591 VSUBS 0.007388f
C632 B.n592 VSUBS 0.007388f
C633 B.n593 VSUBS 0.007388f
C634 B.n594 VSUBS 0.007388f
C635 B.n595 VSUBS 0.007388f
C636 B.n596 VSUBS 0.007388f
C637 B.n597 VSUBS 0.007388f
C638 B.n598 VSUBS 0.007388f
C639 B.n599 VSUBS 0.007388f
C640 B.n600 VSUBS 0.007388f
C641 B.n601 VSUBS 0.007388f
C642 B.n602 VSUBS 0.007388f
C643 B.n603 VSUBS 0.007388f
C644 B.n604 VSUBS 0.007388f
C645 B.n605 VSUBS 0.007388f
C646 B.n606 VSUBS 0.007388f
C647 B.n607 VSUBS 0.007388f
C648 B.n608 VSUBS 0.007388f
C649 B.n609 VSUBS 0.007388f
C650 B.n610 VSUBS 0.007388f
C651 B.n611 VSUBS 0.007388f
C652 B.n612 VSUBS 0.007388f
C653 B.n613 VSUBS 0.007388f
C654 B.n614 VSUBS 0.007388f
C655 B.n615 VSUBS 0.007388f
C656 B.n616 VSUBS 0.007388f
C657 B.n617 VSUBS 0.007388f
C658 B.n618 VSUBS 0.007388f
C659 B.n619 VSUBS 0.007388f
C660 B.n620 VSUBS 0.007388f
C661 B.n621 VSUBS 0.007388f
C662 B.n622 VSUBS 0.007388f
C663 B.n623 VSUBS 0.007388f
C664 B.n624 VSUBS 0.007388f
C665 B.n625 VSUBS 0.007388f
C666 B.n626 VSUBS 0.007388f
C667 B.n627 VSUBS 0.007388f
C668 B.n628 VSUBS 0.007388f
C669 B.n629 VSUBS 0.007388f
C670 B.n630 VSUBS 0.007388f
C671 B.n631 VSUBS 0.007388f
C672 B.n632 VSUBS 0.007388f
C673 B.n633 VSUBS 0.007388f
C674 B.n634 VSUBS 0.007388f
C675 B.n635 VSUBS 0.007388f
C676 B.n636 VSUBS 0.007388f
C677 B.n637 VSUBS 0.007388f
C678 B.n638 VSUBS 0.007388f
C679 B.n639 VSUBS 0.007388f
C680 B.n640 VSUBS 0.007388f
C681 B.n641 VSUBS 0.007388f
C682 B.n642 VSUBS 0.007388f
C683 B.n643 VSUBS 0.007388f
C684 B.n644 VSUBS 0.007388f
C685 B.n645 VSUBS 0.007388f
C686 B.n646 VSUBS 0.007388f
C687 B.n647 VSUBS 0.007388f
C688 B.n648 VSUBS 0.007388f
C689 B.n649 VSUBS 0.007388f
C690 B.n650 VSUBS 0.007388f
C691 B.n651 VSUBS 0.007388f
C692 B.n652 VSUBS 0.007388f
C693 B.n653 VSUBS 0.007388f
C694 B.n654 VSUBS 0.007388f
C695 B.n655 VSUBS 0.007388f
C696 B.n656 VSUBS 0.007388f
C697 B.n657 VSUBS 0.007388f
C698 B.n658 VSUBS 0.007388f
C699 B.n659 VSUBS 0.007388f
C700 B.n660 VSUBS 0.007388f
C701 B.n661 VSUBS 0.007388f
C702 B.n662 VSUBS 0.007388f
C703 B.n663 VSUBS 0.007388f
C704 B.n664 VSUBS 0.007388f
C705 B.n665 VSUBS 0.016339f
C706 B.n666 VSUBS 0.017123f
C707 B.n667 VSUBS 0.017123f
C708 B.n668 VSUBS 0.007388f
C709 B.n669 VSUBS 0.007388f
C710 B.n670 VSUBS 0.007388f
C711 B.n671 VSUBS 0.007388f
C712 B.n672 VSUBS 0.007388f
C713 B.n673 VSUBS 0.007388f
C714 B.n674 VSUBS 0.007388f
C715 B.n675 VSUBS 0.007388f
C716 B.n676 VSUBS 0.007388f
C717 B.n677 VSUBS 0.007388f
C718 B.n678 VSUBS 0.007388f
C719 B.n679 VSUBS 0.007388f
C720 B.n680 VSUBS 0.007388f
C721 B.n681 VSUBS 0.007388f
C722 B.n682 VSUBS 0.007388f
C723 B.n683 VSUBS 0.007388f
C724 B.n684 VSUBS 0.007388f
C725 B.n685 VSUBS 0.007388f
C726 B.n686 VSUBS 0.007388f
C727 B.n687 VSUBS 0.007388f
C728 B.n688 VSUBS 0.007388f
C729 B.n689 VSUBS 0.007388f
C730 B.n690 VSUBS 0.007388f
C731 B.n691 VSUBS 0.007388f
C732 B.n692 VSUBS 0.007388f
C733 B.n693 VSUBS 0.007388f
C734 B.n694 VSUBS 0.007388f
C735 B.n695 VSUBS 0.007388f
C736 B.n696 VSUBS 0.007388f
C737 B.n697 VSUBS 0.007388f
C738 B.n698 VSUBS 0.007388f
C739 B.n699 VSUBS 0.007388f
C740 B.n700 VSUBS 0.007388f
C741 B.n701 VSUBS 0.007388f
C742 B.n702 VSUBS 0.007388f
C743 B.n703 VSUBS 0.007388f
C744 B.n704 VSUBS 0.007388f
C745 B.n705 VSUBS 0.007388f
C746 B.n706 VSUBS 0.007388f
C747 B.n707 VSUBS 0.007388f
C748 B.n708 VSUBS 0.007388f
C749 B.n709 VSUBS 0.007388f
C750 B.n710 VSUBS 0.007388f
C751 B.n711 VSUBS 0.007388f
C752 B.n712 VSUBS 0.007388f
C753 B.n713 VSUBS 0.007388f
C754 B.n714 VSUBS 0.007388f
C755 B.n715 VSUBS 0.007388f
C756 B.n716 VSUBS 0.007388f
C757 B.n717 VSUBS 0.007388f
C758 B.n718 VSUBS 0.007388f
C759 B.n719 VSUBS 0.007388f
C760 B.n720 VSUBS 0.007388f
C761 B.n721 VSUBS 0.007388f
C762 B.n722 VSUBS 0.007388f
C763 B.n723 VSUBS 0.007388f
C764 B.n724 VSUBS 0.007388f
C765 B.n725 VSUBS 0.007388f
C766 B.n726 VSUBS 0.007388f
C767 B.n727 VSUBS 0.007388f
C768 B.n728 VSUBS 0.007388f
C769 B.n729 VSUBS 0.007388f
C770 B.n730 VSUBS 0.007388f
C771 B.n731 VSUBS 0.007388f
C772 B.n732 VSUBS 0.007388f
C773 B.n733 VSUBS 0.007388f
C774 B.n734 VSUBS 0.007388f
C775 B.n735 VSUBS 0.007388f
C776 B.n736 VSUBS 0.007388f
C777 B.n737 VSUBS 0.007388f
C778 B.n738 VSUBS 0.007388f
C779 B.n739 VSUBS 0.007388f
C780 B.n740 VSUBS 0.007388f
C781 B.n741 VSUBS 0.007388f
C782 B.n742 VSUBS 0.007388f
C783 B.n743 VSUBS 0.007388f
C784 B.n744 VSUBS 0.007388f
C785 B.n745 VSUBS 0.007388f
C786 B.n746 VSUBS 0.007388f
C787 B.n747 VSUBS 0.007388f
C788 B.n748 VSUBS 0.007388f
C789 B.n749 VSUBS 0.007388f
C790 B.n750 VSUBS 0.007388f
C791 B.n751 VSUBS 0.007388f
C792 B.n752 VSUBS 0.007388f
C793 B.n753 VSUBS 0.006953f
C794 B.n754 VSUBS 0.007388f
C795 B.n755 VSUBS 0.007388f
C796 B.n756 VSUBS 0.004128f
C797 B.n757 VSUBS 0.007388f
C798 B.n758 VSUBS 0.007388f
C799 B.n759 VSUBS 0.007388f
C800 B.n760 VSUBS 0.007388f
C801 B.n761 VSUBS 0.007388f
C802 B.n762 VSUBS 0.007388f
C803 B.n763 VSUBS 0.007388f
C804 B.n764 VSUBS 0.007388f
C805 B.n765 VSUBS 0.007388f
C806 B.n766 VSUBS 0.007388f
C807 B.n767 VSUBS 0.007388f
C808 B.n768 VSUBS 0.007388f
C809 B.n769 VSUBS 0.004128f
C810 B.n770 VSUBS 0.017117f
C811 B.n771 VSUBS 0.006953f
C812 B.n772 VSUBS 0.007388f
C813 B.n773 VSUBS 0.007388f
C814 B.n774 VSUBS 0.007388f
C815 B.n775 VSUBS 0.007388f
C816 B.n776 VSUBS 0.007388f
C817 B.n777 VSUBS 0.007388f
C818 B.n778 VSUBS 0.007388f
C819 B.n779 VSUBS 0.007388f
C820 B.n780 VSUBS 0.007388f
C821 B.n781 VSUBS 0.007388f
C822 B.n782 VSUBS 0.007388f
C823 B.n783 VSUBS 0.007388f
C824 B.n784 VSUBS 0.007388f
C825 B.n785 VSUBS 0.007388f
C826 B.n786 VSUBS 0.007388f
C827 B.n787 VSUBS 0.007388f
C828 B.n788 VSUBS 0.007388f
C829 B.n789 VSUBS 0.007388f
C830 B.n790 VSUBS 0.007388f
C831 B.n791 VSUBS 0.007388f
C832 B.n792 VSUBS 0.007388f
C833 B.n793 VSUBS 0.007388f
C834 B.n794 VSUBS 0.007388f
C835 B.n795 VSUBS 0.007388f
C836 B.n796 VSUBS 0.007388f
C837 B.n797 VSUBS 0.007388f
C838 B.n798 VSUBS 0.007388f
C839 B.n799 VSUBS 0.007388f
C840 B.n800 VSUBS 0.007388f
C841 B.n801 VSUBS 0.007388f
C842 B.n802 VSUBS 0.007388f
C843 B.n803 VSUBS 0.007388f
C844 B.n804 VSUBS 0.007388f
C845 B.n805 VSUBS 0.007388f
C846 B.n806 VSUBS 0.007388f
C847 B.n807 VSUBS 0.007388f
C848 B.n808 VSUBS 0.007388f
C849 B.n809 VSUBS 0.007388f
C850 B.n810 VSUBS 0.007388f
C851 B.n811 VSUBS 0.007388f
C852 B.n812 VSUBS 0.007388f
C853 B.n813 VSUBS 0.007388f
C854 B.n814 VSUBS 0.007388f
C855 B.n815 VSUBS 0.007388f
C856 B.n816 VSUBS 0.007388f
C857 B.n817 VSUBS 0.007388f
C858 B.n818 VSUBS 0.007388f
C859 B.n819 VSUBS 0.007388f
C860 B.n820 VSUBS 0.007388f
C861 B.n821 VSUBS 0.007388f
C862 B.n822 VSUBS 0.007388f
C863 B.n823 VSUBS 0.007388f
C864 B.n824 VSUBS 0.007388f
C865 B.n825 VSUBS 0.007388f
C866 B.n826 VSUBS 0.007388f
C867 B.n827 VSUBS 0.007388f
C868 B.n828 VSUBS 0.007388f
C869 B.n829 VSUBS 0.007388f
C870 B.n830 VSUBS 0.007388f
C871 B.n831 VSUBS 0.007388f
C872 B.n832 VSUBS 0.007388f
C873 B.n833 VSUBS 0.007388f
C874 B.n834 VSUBS 0.007388f
C875 B.n835 VSUBS 0.007388f
C876 B.n836 VSUBS 0.007388f
C877 B.n837 VSUBS 0.007388f
C878 B.n838 VSUBS 0.007388f
C879 B.n839 VSUBS 0.007388f
C880 B.n840 VSUBS 0.007388f
C881 B.n841 VSUBS 0.007388f
C882 B.n842 VSUBS 0.007388f
C883 B.n843 VSUBS 0.007388f
C884 B.n844 VSUBS 0.007388f
C885 B.n845 VSUBS 0.007388f
C886 B.n846 VSUBS 0.007388f
C887 B.n847 VSUBS 0.007388f
C888 B.n848 VSUBS 0.007388f
C889 B.n849 VSUBS 0.007388f
C890 B.n850 VSUBS 0.007388f
C891 B.n851 VSUBS 0.007388f
C892 B.n852 VSUBS 0.007388f
C893 B.n853 VSUBS 0.007388f
C894 B.n854 VSUBS 0.007388f
C895 B.n855 VSUBS 0.007388f
C896 B.n856 VSUBS 0.007388f
C897 B.n857 VSUBS 0.007388f
C898 B.n858 VSUBS 0.017123f
C899 B.n859 VSUBS 0.017123f
C900 B.n860 VSUBS 0.016339f
C901 B.n861 VSUBS 0.007388f
C902 B.n862 VSUBS 0.007388f
C903 B.n863 VSUBS 0.007388f
C904 B.n864 VSUBS 0.007388f
C905 B.n865 VSUBS 0.007388f
C906 B.n866 VSUBS 0.007388f
C907 B.n867 VSUBS 0.007388f
C908 B.n868 VSUBS 0.007388f
C909 B.n869 VSUBS 0.007388f
C910 B.n870 VSUBS 0.007388f
C911 B.n871 VSUBS 0.007388f
C912 B.n872 VSUBS 0.007388f
C913 B.n873 VSUBS 0.007388f
C914 B.n874 VSUBS 0.007388f
C915 B.n875 VSUBS 0.007388f
C916 B.n876 VSUBS 0.007388f
C917 B.n877 VSUBS 0.007388f
C918 B.n878 VSUBS 0.007388f
C919 B.n879 VSUBS 0.007388f
C920 B.n880 VSUBS 0.007388f
C921 B.n881 VSUBS 0.007388f
C922 B.n882 VSUBS 0.007388f
C923 B.n883 VSUBS 0.007388f
C924 B.n884 VSUBS 0.007388f
C925 B.n885 VSUBS 0.007388f
C926 B.n886 VSUBS 0.007388f
C927 B.n887 VSUBS 0.007388f
C928 B.n888 VSUBS 0.007388f
C929 B.n889 VSUBS 0.007388f
C930 B.n890 VSUBS 0.007388f
C931 B.n891 VSUBS 0.007388f
C932 B.n892 VSUBS 0.007388f
C933 B.n893 VSUBS 0.007388f
C934 B.n894 VSUBS 0.007388f
C935 B.n895 VSUBS 0.007388f
C936 B.n896 VSUBS 0.007388f
C937 B.n897 VSUBS 0.007388f
C938 B.n898 VSUBS 0.007388f
C939 B.n899 VSUBS 0.007388f
C940 B.n900 VSUBS 0.007388f
C941 B.n901 VSUBS 0.007388f
C942 B.n902 VSUBS 0.007388f
C943 B.n903 VSUBS 0.007388f
C944 B.n904 VSUBS 0.007388f
C945 B.n905 VSUBS 0.007388f
C946 B.n906 VSUBS 0.007388f
C947 B.n907 VSUBS 0.007388f
C948 B.n908 VSUBS 0.007388f
C949 B.n909 VSUBS 0.007388f
C950 B.n910 VSUBS 0.007388f
C951 B.n911 VSUBS 0.007388f
C952 B.n912 VSUBS 0.007388f
C953 B.n913 VSUBS 0.007388f
C954 B.n914 VSUBS 0.007388f
C955 B.n915 VSUBS 0.007388f
C956 B.n916 VSUBS 0.007388f
C957 B.n917 VSUBS 0.007388f
C958 B.n918 VSUBS 0.007388f
C959 B.n919 VSUBS 0.007388f
C960 B.n920 VSUBS 0.007388f
C961 B.n921 VSUBS 0.007388f
C962 B.n922 VSUBS 0.007388f
C963 B.n923 VSUBS 0.007388f
C964 B.n924 VSUBS 0.007388f
C965 B.n925 VSUBS 0.007388f
C966 B.n926 VSUBS 0.007388f
C967 B.n927 VSUBS 0.007388f
C968 B.n928 VSUBS 0.007388f
C969 B.n929 VSUBS 0.007388f
C970 B.n930 VSUBS 0.007388f
C971 B.n931 VSUBS 0.007388f
C972 B.n932 VSUBS 0.007388f
C973 B.n933 VSUBS 0.007388f
C974 B.n934 VSUBS 0.007388f
C975 B.n935 VSUBS 0.009641f
C976 B.n936 VSUBS 0.01027f
C977 B.n937 VSUBS 0.020422f
C978 VDD2.t3 VSUBS 4.20623f
C979 VDD2.t4 VSUBS 0.386987f
C980 VDD2.t0 VSUBS 0.386987f
C981 VDD2.n0 VSUBS 3.23096f
C982 VDD2.n1 VSUBS 4.554f
C983 VDD2.t5 VSUBS 4.18004f
C984 VDD2.n2 VSUBS 4.09658f
C985 VDD2.t1 VSUBS 0.386987f
C986 VDD2.t2 VSUBS 0.386987f
C987 VDD2.n3 VSUBS 3.2309f
C988 VN.t5 VSUBS 3.90512f
C989 VN.n0 VSUBS 1.43382f
C990 VN.n1 VSUBS 0.023585f
C991 VN.n2 VSUBS 0.02816f
C992 VN.n3 VSUBS 0.023585f
C993 VN.t1 VSUBS 3.90512f
C994 VN.n4 VSUBS 1.44063f
C995 VN.t2 VSUBS 4.2157f
C996 VN.n5 VSUBS 1.37343f
C997 VN.n6 VSUBS 0.287631f
C998 VN.n7 VSUBS 0.043956f
C999 VN.n8 VSUBS 0.043956f
C1000 VN.n9 VSUBS 0.040287f
C1001 VN.n10 VSUBS 0.023585f
C1002 VN.n11 VSUBS 0.023585f
C1003 VN.n12 VSUBS 0.023585f
C1004 VN.n13 VSUBS 0.044369f
C1005 VN.n14 VSUBS 0.043956f
C1006 VN.n15 VSUBS 0.030067f
C1007 VN.n16 VSUBS 0.038065f
C1008 VN.n17 VSUBS 0.06259f
C1009 VN.t0 VSUBS 3.90512f
C1010 VN.n18 VSUBS 1.43382f
C1011 VN.n19 VSUBS 0.023585f
C1012 VN.n20 VSUBS 0.02816f
C1013 VN.n21 VSUBS 0.023585f
C1014 VN.t4 VSUBS 3.90512f
C1015 VN.n22 VSUBS 1.44063f
C1016 VN.t3 VSUBS 4.2157f
C1017 VN.n23 VSUBS 1.37343f
C1018 VN.n24 VSUBS 0.287631f
C1019 VN.n25 VSUBS 0.043956f
C1020 VN.n26 VSUBS 0.043956f
C1021 VN.n27 VSUBS 0.040287f
C1022 VN.n28 VSUBS 0.023585f
C1023 VN.n29 VSUBS 0.023585f
C1024 VN.n30 VSUBS 0.023585f
C1025 VN.n31 VSUBS 0.044369f
C1026 VN.n32 VSUBS 0.043956f
C1027 VN.n33 VSUBS 0.030067f
C1028 VN.n34 VSUBS 0.038065f
C1029 VN.n35 VSUBS 1.59297f
C1030 VDD1.t1 VSUBS 4.20768f
C1031 VDD1.t3 VSUBS 4.20613f
C1032 VDD1.t2 VSUBS 0.386978f
C1033 VDD1.t0 VSUBS 0.386978f
C1034 VDD1.n0 VSUBS 3.23088f
C1035 VDD1.n1 VSUBS 4.71584f
C1036 VDD1.t4 VSUBS 0.386978f
C1037 VDD1.t5 VSUBS 0.386978f
C1038 VDD1.n2 VSUBS 3.22171f
C1039 VDD1.n3 VSUBS 4.06707f
C1040 VTAIL.t5 VSUBS 0.398314f
C1041 VTAIL.t3 VSUBS 0.398314f
C1042 VTAIL.n0 VSUBS 3.14907f
C1043 VTAIL.n1 VSUBS 0.936963f
C1044 VTAIL.t7 VSUBS 4.11083f
C1045 VTAIL.n2 VSUBS 1.2713f
C1046 VTAIL.t10 VSUBS 0.398314f
C1047 VTAIL.t8 VSUBS 0.398314f
C1048 VTAIL.n3 VSUBS 3.14907f
C1049 VTAIL.n4 VSUBS 3.31553f
C1050 VTAIL.t1 VSUBS 0.398314f
C1051 VTAIL.t2 VSUBS 0.398314f
C1052 VTAIL.n5 VSUBS 3.14908f
C1053 VTAIL.n6 VSUBS 3.31552f
C1054 VTAIL.t0 VSUBS 4.11084f
C1055 VTAIL.n7 VSUBS 1.27129f
C1056 VTAIL.t11 VSUBS 0.398314f
C1057 VTAIL.t6 VSUBS 0.398314f
C1058 VTAIL.n8 VSUBS 3.14908f
C1059 VTAIL.n9 VSUBS 1.14674f
C1060 VTAIL.t9 VSUBS 4.11083f
C1061 VTAIL.n10 VSUBS 3.15335f
C1062 VTAIL.t4 VSUBS 4.11083f
C1063 VTAIL.n11 VSUBS 3.07641f
C1064 VP.t5 VSUBS 4.23432f
C1065 VP.n0 VSUBS 1.55469f
C1066 VP.n1 VSUBS 0.025573f
C1067 VP.n2 VSUBS 0.030534f
C1068 VP.n3 VSUBS 0.025573f
C1069 VP.t3 VSUBS 4.23432f
C1070 VP.n4 VSUBS 1.48578f
C1071 VP.n5 VSUBS 0.025573f
C1072 VP.n6 VSUBS 0.030534f
C1073 VP.n7 VSUBS 0.025573f
C1074 VP.t2 VSUBS 4.23432f
C1075 VP.n8 VSUBS 1.55469f
C1076 VP.t0 VSUBS 4.23432f
C1077 VP.n9 VSUBS 1.55469f
C1078 VP.n10 VSUBS 0.025573f
C1079 VP.n11 VSUBS 0.030534f
C1080 VP.n12 VSUBS 0.025573f
C1081 VP.t1 VSUBS 4.23432f
C1082 VP.n13 VSUBS 1.56208f
C1083 VP.t4 VSUBS 4.57108f
C1084 VP.n14 VSUBS 1.48921f
C1085 VP.n15 VSUBS 0.311879f
C1086 VP.n16 VSUBS 0.047662f
C1087 VP.n17 VSUBS 0.047662f
C1088 VP.n18 VSUBS 0.043683f
C1089 VP.n19 VSUBS 0.025573f
C1090 VP.n20 VSUBS 0.025573f
C1091 VP.n21 VSUBS 0.025573f
C1092 VP.n22 VSUBS 0.048109f
C1093 VP.n23 VSUBS 0.047662f
C1094 VP.n24 VSUBS 0.032602f
C1095 VP.n25 VSUBS 0.041274f
C1096 VP.n26 VSUBS 1.71718f
C1097 VP.n27 VSUBS 1.73354f
C1098 VP.n28 VSUBS 0.041274f
C1099 VP.n29 VSUBS 0.032602f
C1100 VP.n30 VSUBS 0.047662f
C1101 VP.n31 VSUBS 0.048109f
C1102 VP.n32 VSUBS 0.025573f
C1103 VP.n33 VSUBS 0.025573f
C1104 VP.n34 VSUBS 0.025573f
C1105 VP.n35 VSUBS 0.043683f
C1106 VP.n36 VSUBS 0.047662f
C1107 VP.n37 VSUBS 0.047662f
C1108 VP.n38 VSUBS 0.025573f
C1109 VP.n39 VSUBS 0.025573f
C1110 VP.n40 VSUBS 0.025573f
C1111 VP.n41 VSUBS 0.047662f
C1112 VP.n42 VSUBS 0.047662f
C1113 VP.n43 VSUBS 0.043683f
C1114 VP.n44 VSUBS 0.025573f
C1115 VP.n45 VSUBS 0.025573f
C1116 VP.n46 VSUBS 0.025573f
C1117 VP.n47 VSUBS 0.048109f
C1118 VP.n48 VSUBS 0.047662f
C1119 VP.n49 VSUBS 0.032602f
C1120 VP.n50 VSUBS 0.041274f
C1121 VP.n51 VSUBS 0.067867f
.ends

