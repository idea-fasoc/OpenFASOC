* NGSPICE file created from diff_pair_sample_0520.ext - technology: sky130A

.subckt diff_pair_sample_0520 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t9 w_n3660_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=3.2076 ps=19.77 w=19.44 l=2.36
X1 B.t11 B.t9 B.t10 w_n3660_n4856# sky130_fd_pr__pfet_01v8 ad=7.5816 pd=39.66 as=0 ps=0 w=19.44 l=2.36
X2 VDD2.t7 VN.t0 VTAIL.t2 w_n3660_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=3.2076 ps=19.77 w=19.44 l=2.36
X3 VTAIL.t12 VP.t1 VDD1.t6 w_n3660_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=3.2076 ps=19.77 w=19.44 l=2.36
X4 VTAIL.t1 VN.t1 VDD2.t6 w_n3660_n4856# sky130_fd_pr__pfet_01v8 ad=7.5816 pd=39.66 as=3.2076 ps=19.77 w=19.44 l=2.36
X5 VDD1.t5 VP.t2 VTAIL.t10 w_n3660_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=7.5816 ps=39.66 w=19.44 l=2.36
X6 VTAIL.t5 VN.t2 VDD2.t5 w_n3660_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=3.2076 ps=19.77 w=19.44 l=2.36
X7 VDD2.t4 VN.t3 VTAIL.t0 w_n3660_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=7.5816 ps=39.66 w=19.44 l=2.36
X8 VDD1.t4 VP.t3 VTAIL.t13 w_n3660_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=3.2076 ps=19.77 w=19.44 l=2.36
X9 VTAIL.t3 VN.t4 VDD2.t3 w_n3660_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=3.2076 ps=19.77 w=19.44 l=2.36
X10 VTAIL.t14 VP.t4 VDD1.t3 w_n3660_n4856# sky130_fd_pr__pfet_01v8 ad=7.5816 pd=39.66 as=3.2076 ps=19.77 w=19.44 l=2.36
X11 VDD2.t2 VN.t5 VTAIL.t4 w_n3660_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=7.5816 ps=39.66 w=19.44 l=2.36
X12 VTAIL.t7 VN.t6 VDD2.t1 w_n3660_n4856# sky130_fd_pr__pfet_01v8 ad=7.5816 pd=39.66 as=3.2076 ps=19.77 w=19.44 l=2.36
X13 VDD1.t2 VP.t5 VTAIL.t11 w_n3660_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=7.5816 ps=39.66 w=19.44 l=2.36
X14 B.t8 B.t6 B.t7 w_n3660_n4856# sky130_fd_pr__pfet_01v8 ad=7.5816 pd=39.66 as=0 ps=0 w=19.44 l=2.36
X15 B.t5 B.t3 B.t4 w_n3660_n4856# sky130_fd_pr__pfet_01v8 ad=7.5816 pd=39.66 as=0 ps=0 w=19.44 l=2.36
X16 VDD2.t0 VN.t7 VTAIL.t6 w_n3660_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=3.2076 ps=19.77 w=19.44 l=2.36
X17 B.t2 B.t0 B.t1 w_n3660_n4856# sky130_fd_pr__pfet_01v8 ad=7.5816 pd=39.66 as=0 ps=0 w=19.44 l=2.36
X18 VTAIL.t8 VP.t6 VDD1.t1 w_n3660_n4856# sky130_fd_pr__pfet_01v8 ad=7.5816 pd=39.66 as=3.2076 ps=19.77 w=19.44 l=2.36
X19 VTAIL.t15 VP.t7 VDD1.t0 w_n3660_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=3.2076 ps=19.77 w=19.44 l=2.36
R0 VP.n15 VP.t6 230.635
R1 VP.n36 VP.t4 198.519
R2 VP.n43 VP.t3 198.519
R3 VP.n55 VP.t7 198.519
R4 VP.n63 VP.t5 198.519
R5 VP.n33 VP.t2 198.519
R6 VP.n25 VP.t1 198.519
R7 VP.n14 VP.t0 198.519
R8 VP.n16 VP.n13 161.3
R9 VP.n18 VP.n17 161.3
R10 VP.n19 VP.n12 161.3
R11 VP.n21 VP.n20 161.3
R12 VP.n22 VP.n11 161.3
R13 VP.n24 VP.n23 161.3
R14 VP.n26 VP.n10 161.3
R15 VP.n28 VP.n27 161.3
R16 VP.n29 VP.n9 161.3
R17 VP.n31 VP.n30 161.3
R18 VP.n32 VP.n8 161.3
R19 VP.n62 VP.n0 161.3
R20 VP.n61 VP.n60 161.3
R21 VP.n59 VP.n1 161.3
R22 VP.n58 VP.n57 161.3
R23 VP.n56 VP.n2 161.3
R24 VP.n54 VP.n53 161.3
R25 VP.n52 VP.n3 161.3
R26 VP.n51 VP.n50 161.3
R27 VP.n49 VP.n4 161.3
R28 VP.n48 VP.n47 161.3
R29 VP.n46 VP.n5 161.3
R30 VP.n45 VP.n44 161.3
R31 VP.n42 VP.n6 161.3
R32 VP.n41 VP.n40 161.3
R33 VP.n39 VP.n7 161.3
R34 VP.n38 VP.n37 161.3
R35 VP.n36 VP.n35 96.7304
R36 VP.n64 VP.n63 96.7304
R37 VP.n34 VP.n33 96.7304
R38 VP.n15 VP.n14 67.322
R39 VP.n50 VP.n49 56.4773
R40 VP.n20 VP.n19 56.4773
R41 VP.n35 VP.n34 55.4313
R42 VP.n42 VP.n41 46.253
R43 VP.n57 VP.n1 46.253
R44 VP.n27 VP.n9 46.253
R45 VP.n41 VP.n7 34.5682
R46 VP.n61 VP.n1 34.5682
R47 VP.n31 VP.n9 34.5682
R48 VP.n37 VP.n7 24.3439
R49 VP.n44 VP.n42 24.3439
R50 VP.n48 VP.n5 24.3439
R51 VP.n49 VP.n48 24.3439
R52 VP.n50 VP.n3 24.3439
R53 VP.n54 VP.n3 24.3439
R54 VP.n57 VP.n56 24.3439
R55 VP.n62 VP.n61 24.3439
R56 VP.n32 VP.n31 24.3439
R57 VP.n20 VP.n11 24.3439
R58 VP.n24 VP.n11 24.3439
R59 VP.n27 VP.n26 24.3439
R60 VP.n18 VP.n13 24.3439
R61 VP.n19 VP.n18 24.3439
R62 VP.n44 VP.n43 19.7187
R63 VP.n56 VP.n55 19.7187
R64 VP.n26 VP.n25 19.7187
R65 VP.n37 VP.n36 13.8763
R66 VP.n63 VP.n62 13.8763
R67 VP.n33 VP.n32 13.8763
R68 VP.n16 VP.n15 9.62344
R69 VP.n43 VP.n5 4.62575
R70 VP.n55 VP.n54 4.62575
R71 VP.n25 VP.n24 4.62575
R72 VP.n14 VP.n13 4.62575
R73 VP.n34 VP.n8 0.278398
R74 VP.n38 VP.n35 0.278398
R75 VP.n64 VP.n0 0.278398
R76 VP.n17 VP.n16 0.189894
R77 VP.n17 VP.n12 0.189894
R78 VP.n21 VP.n12 0.189894
R79 VP.n22 VP.n21 0.189894
R80 VP.n23 VP.n22 0.189894
R81 VP.n23 VP.n10 0.189894
R82 VP.n28 VP.n10 0.189894
R83 VP.n29 VP.n28 0.189894
R84 VP.n30 VP.n29 0.189894
R85 VP.n30 VP.n8 0.189894
R86 VP.n39 VP.n38 0.189894
R87 VP.n40 VP.n39 0.189894
R88 VP.n40 VP.n6 0.189894
R89 VP.n45 VP.n6 0.189894
R90 VP.n46 VP.n45 0.189894
R91 VP.n47 VP.n46 0.189894
R92 VP.n47 VP.n4 0.189894
R93 VP.n51 VP.n4 0.189894
R94 VP.n52 VP.n51 0.189894
R95 VP.n53 VP.n52 0.189894
R96 VP.n53 VP.n2 0.189894
R97 VP.n58 VP.n2 0.189894
R98 VP.n59 VP.n58 0.189894
R99 VP.n60 VP.n59 0.189894
R100 VP.n60 VP.n0 0.189894
R101 VP VP.n64 0.153422
R102 VTAIL.n785 VTAIL.n784 585
R103 VTAIL.n782 VTAIL.n781 585
R104 VTAIL.n791 VTAIL.n790 585
R105 VTAIL.n793 VTAIL.n792 585
R106 VTAIL.n778 VTAIL.n777 585
R107 VTAIL.n799 VTAIL.n798 585
R108 VTAIL.n802 VTAIL.n801 585
R109 VTAIL.n800 VTAIL.n774 585
R110 VTAIL.n807 VTAIL.n773 585
R111 VTAIL.n809 VTAIL.n808 585
R112 VTAIL.n811 VTAIL.n810 585
R113 VTAIL.n770 VTAIL.n769 585
R114 VTAIL.n817 VTAIL.n816 585
R115 VTAIL.n819 VTAIL.n818 585
R116 VTAIL.n766 VTAIL.n765 585
R117 VTAIL.n825 VTAIL.n824 585
R118 VTAIL.n827 VTAIL.n826 585
R119 VTAIL.n762 VTAIL.n761 585
R120 VTAIL.n833 VTAIL.n832 585
R121 VTAIL.n835 VTAIL.n834 585
R122 VTAIL.n758 VTAIL.n757 585
R123 VTAIL.n841 VTAIL.n840 585
R124 VTAIL.n843 VTAIL.n842 585
R125 VTAIL.n754 VTAIL.n753 585
R126 VTAIL.n849 VTAIL.n848 585
R127 VTAIL.n851 VTAIL.n850 585
R128 VTAIL.n37 VTAIL.n36 585
R129 VTAIL.n34 VTAIL.n33 585
R130 VTAIL.n43 VTAIL.n42 585
R131 VTAIL.n45 VTAIL.n44 585
R132 VTAIL.n30 VTAIL.n29 585
R133 VTAIL.n51 VTAIL.n50 585
R134 VTAIL.n54 VTAIL.n53 585
R135 VTAIL.n52 VTAIL.n26 585
R136 VTAIL.n59 VTAIL.n25 585
R137 VTAIL.n61 VTAIL.n60 585
R138 VTAIL.n63 VTAIL.n62 585
R139 VTAIL.n22 VTAIL.n21 585
R140 VTAIL.n69 VTAIL.n68 585
R141 VTAIL.n71 VTAIL.n70 585
R142 VTAIL.n18 VTAIL.n17 585
R143 VTAIL.n77 VTAIL.n76 585
R144 VTAIL.n79 VTAIL.n78 585
R145 VTAIL.n14 VTAIL.n13 585
R146 VTAIL.n85 VTAIL.n84 585
R147 VTAIL.n87 VTAIL.n86 585
R148 VTAIL.n10 VTAIL.n9 585
R149 VTAIL.n93 VTAIL.n92 585
R150 VTAIL.n95 VTAIL.n94 585
R151 VTAIL.n6 VTAIL.n5 585
R152 VTAIL.n101 VTAIL.n100 585
R153 VTAIL.n103 VTAIL.n102 585
R154 VTAIL.n143 VTAIL.n142 585
R155 VTAIL.n140 VTAIL.n139 585
R156 VTAIL.n149 VTAIL.n148 585
R157 VTAIL.n151 VTAIL.n150 585
R158 VTAIL.n136 VTAIL.n135 585
R159 VTAIL.n157 VTAIL.n156 585
R160 VTAIL.n160 VTAIL.n159 585
R161 VTAIL.n158 VTAIL.n132 585
R162 VTAIL.n165 VTAIL.n131 585
R163 VTAIL.n167 VTAIL.n166 585
R164 VTAIL.n169 VTAIL.n168 585
R165 VTAIL.n128 VTAIL.n127 585
R166 VTAIL.n175 VTAIL.n174 585
R167 VTAIL.n177 VTAIL.n176 585
R168 VTAIL.n124 VTAIL.n123 585
R169 VTAIL.n183 VTAIL.n182 585
R170 VTAIL.n185 VTAIL.n184 585
R171 VTAIL.n120 VTAIL.n119 585
R172 VTAIL.n191 VTAIL.n190 585
R173 VTAIL.n193 VTAIL.n192 585
R174 VTAIL.n116 VTAIL.n115 585
R175 VTAIL.n199 VTAIL.n198 585
R176 VTAIL.n201 VTAIL.n200 585
R177 VTAIL.n112 VTAIL.n111 585
R178 VTAIL.n207 VTAIL.n206 585
R179 VTAIL.n209 VTAIL.n208 585
R180 VTAIL.n251 VTAIL.n250 585
R181 VTAIL.n248 VTAIL.n247 585
R182 VTAIL.n257 VTAIL.n256 585
R183 VTAIL.n259 VTAIL.n258 585
R184 VTAIL.n244 VTAIL.n243 585
R185 VTAIL.n265 VTAIL.n264 585
R186 VTAIL.n268 VTAIL.n267 585
R187 VTAIL.n266 VTAIL.n240 585
R188 VTAIL.n273 VTAIL.n239 585
R189 VTAIL.n275 VTAIL.n274 585
R190 VTAIL.n277 VTAIL.n276 585
R191 VTAIL.n236 VTAIL.n235 585
R192 VTAIL.n283 VTAIL.n282 585
R193 VTAIL.n285 VTAIL.n284 585
R194 VTAIL.n232 VTAIL.n231 585
R195 VTAIL.n291 VTAIL.n290 585
R196 VTAIL.n293 VTAIL.n292 585
R197 VTAIL.n228 VTAIL.n227 585
R198 VTAIL.n299 VTAIL.n298 585
R199 VTAIL.n301 VTAIL.n300 585
R200 VTAIL.n224 VTAIL.n223 585
R201 VTAIL.n307 VTAIL.n306 585
R202 VTAIL.n309 VTAIL.n308 585
R203 VTAIL.n220 VTAIL.n219 585
R204 VTAIL.n315 VTAIL.n314 585
R205 VTAIL.n317 VTAIL.n316 585
R206 VTAIL.n745 VTAIL.n744 585
R207 VTAIL.n743 VTAIL.n742 585
R208 VTAIL.n648 VTAIL.n647 585
R209 VTAIL.n737 VTAIL.n736 585
R210 VTAIL.n735 VTAIL.n734 585
R211 VTAIL.n652 VTAIL.n651 585
R212 VTAIL.n729 VTAIL.n728 585
R213 VTAIL.n727 VTAIL.n726 585
R214 VTAIL.n656 VTAIL.n655 585
R215 VTAIL.n721 VTAIL.n720 585
R216 VTAIL.n719 VTAIL.n718 585
R217 VTAIL.n660 VTAIL.n659 585
R218 VTAIL.n713 VTAIL.n712 585
R219 VTAIL.n711 VTAIL.n710 585
R220 VTAIL.n664 VTAIL.n663 585
R221 VTAIL.n705 VTAIL.n704 585
R222 VTAIL.n703 VTAIL.n702 585
R223 VTAIL.n701 VTAIL.n667 585
R224 VTAIL.n671 VTAIL.n668 585
R225 VTAIL.n696 VTAIL.n695 585
R226 VTAIL.n694 VTAIL.n693 585
R227 VTAIL.n673 VTAIL.n672 585
R228 VTAIL.n688 VTAIL.n687 585
R229 VTAIL.n686 VTAIL.n685 585
R230 VTAIL.n677 VTAIL.n676 585
R231 VTAIL.n680 VTAIL.n679 585
R232 VTAIL.n637 VTAIL.n636 585
R233 VTAIL.n635 VTAIL.n634 585
R234 VTAIL.n540 VTAIL.n539 585
R235 VTAIL.n629 VTAIL.n628 585
R236 VTAIL.n627 VTAIL.n626 585
R237 VTAIL.n544 VTAIL.n543 585
R238 VTAIL.n621 VTAIL.n620 585
R239 VTAIL.n619 VTAIL.n618 585
R240 VTAIL.n548 VTAIL.n547 585
R241 VTAIL.n613 VTAIL.n612 585
R242 VTAIL.n611 VTAIL.n610 585
R243 VTAIL.n552 VTAIL.n551 585
R244 VTAIL.n605 VTAIL.n604 585
R245 VTAIL.n603 VTAIL.n602 585
R246 VTAIL.n556 VTAIL.n555 585
R247 VTAIL.n597 VTAIL.n596 585
R248 VTAIL.n595 VTAIL.n594 585
R249 VTAIL.n593 VTAIL.n559 585
R250 VTAIL.n563 VTAIL.n560 585
R251 VTAIL.n588 VTAIL.n587 585
R252 VTAIL.n586 VTAIL.n585 585
R253 VTAIL.n565 VTAIL.n564 585
R254 VTAIL.n580 VTAIL.n579 585
R255 VTAIL.n578 VTAIL.n577 585
R256 VTAIL.n569 VTAIL.n568 585
R257 VTAIL.n572 VTAIL.n571 585
R258 VTAIL.n531 VTAIL.n530 585
R259 VTAIL.n529 VTAIL.n528 585
R260 VTAIL.n434 VTAIL.n433 585
R261 VTAIL.n523 VTAIL.n522 585
R262 VTAIL.n521 VTAIL.n520 585
R263 VTAIL.n438 VTAIL.n437 585
R264 VTAIL.n515 VTAIL.n514 585
R265 VTAIL.n513 VTAIL.n512 585
R266 VTAIL.n442 VTAIL.n441 585
R267 VTAIL.n507 VTAIL.n506 585
R268 VTAIL.n505 VTAIL.n504 585
R269 VTAIL.n446 VTAIL.n445 585
R270 VTAIL.n499 VTAIL.n498 585
R271 VTAIL.n497 VTAIL.n496 585
R272 VTAIL.n450 VTAIL.n449 585
R273 VTAIL.n491 VTAIL.n490 585
R274 VTAIL.n489 VTAIL.n488 585
R275 VTAIL.n487 VTAIL.n453 585
R276 VTAIL.n457 VTAIL.n454 585
R277 VTAIL.n482 VTAIL.n481 585
R278 VTAIL.n480 VTAIL.n479 585
R279 VTAIL.n459 VTAIL.n458 585
R280 VTAIL.n474 VTAIL.n473 585
R281 VTAIL.n472 VTAIL.n471 585
R282 VTAIL.n463 VTAIL.n462 585
R283 VTAIL.n466 VTAIL.n465 585
R284 VTAIL.n423 VTAIL.n422 585
R285 VTAIL.n421 VTAIL.n420 585
R286 VTAIL.n326 VTAIL.n325 585
R287 VTAIL.n415 VTAIL.n414 585
R288 VTAIL.n413 VTAIL.n412 585
R289 VTAIL.n330 VTAIL.n329 585
R290 VTAIL.n407 VTAIL.n406 585
R291 VTAIL.n405 VTAIL.n404 585
R292 VTAIL.n334 VTAIL.n333 585
R293 VTAIL.n399 VTAIL.n398 585
R294 VTAIL.n397 VTAIL.n396 585
R295 VTAIL.n338 VTAIL.n337 585
R296 VTAIL.n391 VTAIL.n390 585
R297 VTAIL.n389 VTAIL.n388 585
R298 VTAIL.n342 VTAIL.n341 585
R299 VTAIL.n383 VTAIL.n382 585
R300 VTAIL.n381 VTAIL.n380 585
R301 VTAIL.n379 VTAIL.n345 585
R302 VTAIL.n349 VTAIL.n346 585
R303 VTAIL.n374 VTAIL.n373 585
R304 VTAIL.n372 VTAIL.n371 585
R305 VTAIL.n351 VTAIL.n350 585
R306 VTAIL.n366 VTAIL.n365 585
R307 VTAIL.n364 VTAIL.n363 585
R308 VTAIL.n355 VTAIL.n354 585
R309 VTAIL.n358 VTAIL.n357 585
R310 VTAIL.n850 VTAIL.n750 498.474
R311 VTAIL.n102 VTAIL.n2 498.474
R312 VTAIL.n208 VTAIL.n108 498.474
R313 VTAIL.n316 VTAIL.n216 498.474
R314 VTAIL.n744 VTAIL.n644 498.474
R315 VTAIL.n636 VTAIL.n536 498.474
R316 VTAIL.n530 VTAIL.n430 498.474
R317 VTAIL.n422 VTAIL.n322 498.474
R318 VTAIL.t4 VTAIL.n783 329.036
R319 VTAIL.t7 VTAIL.n35 329.036
R320 VTAIL.t11 VTAIL.n141 329.036
R321 VTAIL.t14 VTAIL.n249 329.036
R322 VTAIL.t10 VTAIL.n678 329.036
R323 VTAIL.t8 VTAIL.n570 329.036
R324 VTAIL.t0 VTAIL.n464 329.036
R325 VTAIL.t1 VTAIL.n356 329.036
R326 VTAIL.n784 VTAIL.n781 171.744
R327 VTAIL.n791 VTAIL.n781 171.744
R328 VTAIL.n792 VTAIL.n791 171.744
R329 VTAIL.n792 VTAIL.n777 171.744
R330 VTAIL.n799 VTAIL.n777 171.744
R331 VTAIL.n801 VTAIL.n799 171.744
R332 VTAIL.n801 VTAIL.n800 171.744
R333 VTAIL.n800 VTAIL.n773 171.744
R334 VTAIL.n809 VTAIL.n773 171.744
R335 VTAIL.n810 VTAIL.n809 171.744
R336 VTAIL.n810 VTAIL.n769 171.744
R337 VTAIL.n817 VTAIL.n769 171.744
R338 VTAIL.n818 VTAIL.n817 171.744
R339 VTAIL.n818 VTAIL.n765 171.744
R340 VTAIL.n825 VTAIL.n765 171.744
R341 VTAIL.n826 VTAIL.n825 171.744
R342 VTAIL.n826 VTAIL.n761 171.744
R343 VTAIL.n833 VTAIL.n761 171.744
R344 VTAIL.n834 VTAIL.n833 171.744
R345 VTAIL.n834 VTAIL.n757 171.744
R346 VTAIL.n841 VTAIL.n757 171.744
R347 VTAIL.n842 VTAIL.n841 171.744
R348 VTAIL.n842 VTAIL.n753 171.744
R349 VTAIL.n849 VTAIL.n753 171.744
R350 VTAIL.n850 VTAIL.n849 171.744
R351 VTAIL.n36 VTAIL.n33 171.744
R352 VTAIL.n43 VTAIL.n33 171.744
R353 VTAIL.n44 VTAIL.n43 171.744
R354 VTAIL.n44 VTAIL.n29 171.744
R355 VTAIL.n51 VTAIL.n29 171.744
R356 VTAIL.n53 VTAIL.n51 171.744
R357 VTAIL.n53 VTAIL.n52 171.744
R358 VTAIL.n52 VTAIL.n25 171.744
R359 VTAIL.n61 VTAIL.n25 171.744
R360 VTAIL.n62 VTAIL.n61 171.744
R361 VTAIL.n62 VTAIL.n21 171.744
R362 VTAIL.n69 VTAIL.n21 171.744
R363 VTAIL.n70 VTAIL.n69 171.744
R364 VTAIL.n70 VTAIL.n17 171.744
R365 VTAIL.n77 VTAIL.n17 171.744
R366 VTAIL.n78 VTAIL.n77 171.744
R367 VTAIL.n78 VTAIL.n13 171.744
R368 VTAIL.n85 VTAIL.n13 171.744
R369 VTAIL.n86 VTAIL.n85 171.744
R370 VTAIL.n86 VTAIL.n9 171.744
R371 VTAIL.n93 VTAIL.n9 171.744
R372 VTAIL.n94 VTAIL.n93 171.744
R373 VTAIL.n94 VTAIL.n5 171.744
R374 VTAIL.n101 VTAIL.n5 171.744
R375 VTAIL.n102 VTAIL.n101 171.744
R376 VTAIL.n142 VTAIL.n139 171.744
R377 VTAIL.n149 VTAIL.n139 171.744
R378 VTAIL.n150 VTAIL.n149 171.744
R379 VTAIL.n150 VTAIL.n135 171.744
R380 VTAIL.n157 VTAIL.n135 171.744
R381 VTAIL.n159 VTAIL.n157 171.744
R382 VTAIL.n159 VTAIL.n158 171.744
R383 VTAIL.n158 VTAIL.n131 171.744
R384 VTAIL.n167 VTAIL.n131 171.744
R385 VTAIL.n168 VTAIL.n167 171.744
R386 VTAIL.n168 VTAIL.n127 171.744
R387 VTAIL.n175 VTAIL.n127 171.744
R388 VTAIL.n176 VTAIL.n175 171.744
R389 VTAIL.n176 VTAIL.n123 171.744
R390 VTAIL.n183 VTAIL.n123 171.744
R391 VTAIL.n184 VTAIL.n183 171.744
R392 VTAIL.n184 VTAIL.n119 171.744
R393 VTAIL.n191 VTAIL.n119 171.744
R394 VTAIL.n192 VTAIL.n191 171.744
R395 VTAIL.n192 VTAIL.n115 171.744
R396 VTAIL.n199 VTAIL.n115 171.744
R397 VTAIL.n200 VTAIL.n199 171.744
R398 VTAIL.n200 VTAIL.n111 171.744
R399 VTAIL.n207 VTAIL.n111 171.744
R400 VTAIL.n208 VTAIL.n207 171.744
R401 VTAIL.n250 VTAIL.n247 171.744
R402 VTAIL.n257 VTAIL.n247 171.744
R403 VTAIL.n258 VTAIL.n257 171.744
R404 VTAIL.n258 VTAIL.n243 171.744
R405 VTAIL.n265 VTAIL.n243 171.744
R406 VTAIL.n267 VTAIL.n265 171.744
R407 VTAIL.n267 VTAIL.n266 171.744
R408 VTAIL.n266 VTAIL.n239 171.744
R409 VTAIL.n275 VTAIL.n239 171.744
R410 VTAIL.n276 VTAIL.n275 171.744
R411 VTAIL.n276 VTAIL.n235 171.744
R412 VTAIL.n283 VTAIL.n235 171.744
R413 VTAIL.n284 VTAIL.n283 171.744
R414 VTAIL.n284 VTAIL.n231 171.744
R415 VTAIL.n291 VTAIL.n231 171.744
R416 VTAIL.n292 VTAIL.n291 171.744
R417 VTAIL.n292 VTAIL.n227 171.744
R418 VTAIL.n299 VTAIL.n227 171.744
R419 VTAIL.n300 VTAIL.n299 171.744
R420 VTAIL.n300 VTAIL.n223 171.744
R421 VTAIL.n307 VTAIL.n223 171.744
R422 VTAIL.n308 VTAIL.n307 171.744
R423 VTAIL.n308 VTAIL.n219 171.744
R424 VTAIL.n315 VTAIL.n219 171.744
R425 VTAIL.n316 VTAIL.n315 171.744
R426 VTAIL.n744 VTAIL.n743 171.744
R427 VTAIL.n743 VTAIL.n647 171.744
R428 VTAIL.n736 VTAIL.n647 171.744
R429 VTAIL.n736 VTAIL.n735 171.744
R430 VTAIL.n735 VTAIL.n651 171.744
R431 VTAIL.n728 VTAIL.n651 171.744
R432 VTAIL.n728 VTAIL.n727 171.744
R433 VTAIL.n727 VTAIL.n655 171.744
R434 VTAIL.n720 VTAIL.n655 171.744
R435 VTAIL.n720 VTAIL.n719 171.744
R436 VTAIL.n719 VTAIL.n659 171.744
R437 VTAIL.n712 VTAIL.n659 171.744
R438 VTAIL.n712 VTAIL.n711 171.744
R439 VTAIL.n711 VTAIL.n663 171.744
R440 VTAIL.n704 VTAIL.n663 171.744
R441 VTAIL.n704 VTAIL.n703 171.744
R442 VTAIL.n703 VTAIL.n667 171.744
R443 VTAIL.n671 VTAIL.n667 171.744
R444 VTAIL.n695 VTAIL.n671 171.744
R445 VTAIL.n695 VTAIL.n694 171.744
R446 VTAIL.n694 VTAIL.n672 171.744
R447 VTAIL.n687 VTAIL.n672 171.744
R448 VTAIL.n687 VTAIL.n686 171.744
R449 VTAIL.n686 VTAIL.n676 171.744
R450 VTAIL.n679 VTAIL.n676 171.744
R451 VTAIL.n636 VTAIL.n635 171.744
R452 VTAIL.n635 VTAIL.n539 171.744
R453 VTAIL.n628 VTAIL.n539 171.744
R454 VTAIL.n628 VTAIL.n627 171.744
R455 VTAIL.n627 VTAIL.n543 171.744
R456 VTAIL.n620 VTAIL.n543 171.744
R457 VTAIL.n620 VTAIL.n619 171.744
R458 VTAIL.n619 VTAIL.n547 171.744
R459 VTAIL.n612 VTAIL.n547 171.744
R460 VTAIL.n612 VTAIL.n611 171.744
R461 VTAIL.n611 VTAIL.n551 171.744
R462 VTAIL.n604 VTAIL.n551 171.744
R463 VTAIL.n604 VTAIL.n603 171.744
R464 VTAIL.n603 VTAIL.n555 171.744
R465 VTAIL.n596 VTAIL.n555 171.744
R466 VTAIL.n596 VTAIL.n595 171.744
R467 VTAIL.n595 VTAIL.n559 171.744
R468 VTAIL.n563 VTAIL.n559 171.744
R469 VTAIL.n587 VTAIL.n563 171.744
R470 VTAIL.n587 VTAIL.n586 171.744
R471 VTAIL.n586 VTAIL.n564 171.744
R472 VTAIL.n579 VTAIL.n564 171.744
R473 VTAIL.n579 VTAIL.n578 171.744
R474 VTAIL.n578 VTAIL.n568 171.744
R475 VTAIL.n571 VTAIL.n568 171.744
R476 VTAIL.n530 VTAIL.n529 171.744
R477 VTAIL.n529 VTAIL.n433 171.744
R478 VTAIL.n522 VTAIL.n433 171.744
R479 VTAIL.n522 VTAIL.n521 171.744
R480 VTAIL.n521 VTAIL.n437 171.744
R481 VTAIL.n514 VTAIL.n437 171.744
R482 VTAIL.n514 VTAIL.n513 171.744
R483 VTAIL.n513 VTAIL.n441 171.744
R484 VTAIL.n506 VTAIL.n441 171.744
R485 VTAIL.n506 VTAIL.n505 171.744
R486 VTAIL.n505 VTAIL.n445 171.744
R487 VTAIL.n498 VTAIL.n445 171.744
R488 VTAIL.n498 VTAIL.n497 171.744
R489 VTAIL.n497 VTAIL.n449 171.744
R490 VTAIL.n490 VTAIL.n449 171.744
R491 VTAIL.n490 VTAIL.n489 171.744
R492 VTAIL.n489 VTAIL.n453 171.744
R493 VTAIL.n457 VTAIL.n453 171.744
R494 VTAIL.n481 VTAIL.n457 171.744
R495 VTAIL.n481 VTAIL.n480 171.744
R496 VTAIL.n480 VTAIL.n458 171.744
R497 VTAIL.n473 VTAIL.n458 171.744
R498 VTAIL.n473 VTAIL.n472 171.744
R499 VTAIL.n472 VTAIL.n462 171.744
R500 VTAIL.n465 VTAIL.n462 171.744
R501 VTAIL.n422 VTAIL.n421 171.744
R502 VTAIL.n421 VTAIL.n325 171.744
R503 VTAIL.n414 VTAIL.n325 171.744
R504 VTAIL.n414 VTAIL.n413 171.744
R505 VTAIL.n413 VTAIL.n329 171.744
R506 VTAIL.n406 VTAIL.n329 171.744
R507 VTAIL.n406 VTAIL.n405 171.744
R508 VTAIL.n405 VTAIL.n333 171.744
R509 VTAIL.n398 VTAIL.n333 171.744
R510 VTAIL.n398 VTAIL.n397 171.744
R511 VTAIL.n397 VTAIL.n337 171.744
R512 VTAIL.n390 VTAIL.n337 171.744
R513 VTAIL.n390 VTAIL.n389 171.744
R514 VTAIL.n389 VTAIL.n341 171.744
R515 VTAIL.n382 VTAIL.n341 171.744
R516 VTAIL.n382 VTAIL.n381 171.744
R517 VTAIL.n381 VTAIL.n345 171.744
R518 VTAIL.n349 VTAIL.n345 171.744
R519 VTAIL.n373 VTAIL.n349 171.744
R520 VTAIL.n373 VTAIL.n372 171.744
R521 VTAIL.n372 VTAIL.n350 171.744
R522 VTAIL.n365 VTAIL.n350 171.744
R523 VTAIL.n365 VTAIL.n364 171.744
R524 VTAIL.n364 VTAIL.n354 171.744
R525 VTAIL.n357 VTAIL.n354 171.744
R526 VTAIL.n784 VTAIL.t4 85.8723
R527 VTAIL.n36 VTAIL.t7 85.8723
R528 VTAIL.n142 VTAIL.t11 85.8723
R529 VTAIL.n250 VTAIL.t14 85.8723
R530 VTAIL.n679 VTAIL.t10 85.8723
R531 VTAIL.n571 VTAIL.t8 85.8723
R532 VTAIL.n465 VTAIL.t0 85.8723
R533 VTAIL.n357 VTAIL.t1 85.8723
R534 VTAIL.n643 VTAIL.n642 53.4917
R535 VTAIL.n429 VTAIL.n428 53.4917
R536 VTAIL.n1 VTAIL.n0 53.4916
R537 VTAIL.n215 VTAIL.n214 53.4916
R538 VTAIL.n855 VTAIL.n854 34.5126
R539 VTAIL.n107 VTAIL.n106 34.5126
R540 VTAIL.n213 VTAIL.n212 34.5126
R541 VTAIL.n321 VTAIL.n320 34.5126
R542 VTAIL.n749 VTAIL.n748 34.5126
R543 VTAIL.n641 VTAIL.n640 34.5126
R544 VTAIL.n535 VTAIL.n534 34.5126
R545 VTAIL.n427 VTAIL.n426 34.5126
R546 VTAIL.n855 VTAIL.n749 31.4445
R547 VTAIL.n427 VTAIL.n321 31.4445
R548 VTAIL.n808 VTAIL.n807 13.1884
R549 VTAIL.n60 VTAIL.n59 13.1884
R550 VTAIL.n166 VTAIL.n165 13.1884
R551 VTAIL.n274 VTAIL.n273 13.1884
R552 VTAIL.n702 VTAIL.n701 13.1884
R553 VTAIL.n594 VTAIL.n593 13.1884
R554 VTAIL.n488 VTAIL.n487 13.1884
R555 VTAIL.n380 VTAIL.n379 13.1884
R556 VTAIL.n806 VTAIL.n774 12.8005
R557 VTAIL.n811 VTAIL.n772 12.8005
R558 VTAIL.n852 VTAIL.n851 12.8005
R559 VTAIL.n58 VTAIL.n26 12.8005
R560 VTAIL.n63 VTAIL.n24 12.8005
R561 VTAIL.n104 VTAIL.n103 12.8005
R562 VTAIL.n164 VTAIL.n132 12.8005
R563 VTAIL.n169 VTAIL.n130 12.8005
R564 VTAIL.n210 VTAIL.n209 12.8005
R565 VTAIL.n272 VTAIL.n240 12.8005
R566 VTAIL.n277 VTAIL.n238 12.8005
R567 VTAIL.n318 VTAIL.n317 12.8005
R568 VTAIL.n746 VTAIL.n745 12.8005
R569 VTAIL.n705 VTAIL.n666 12.8005
R570 VTAIL.n700 VTAIL.n668 12.8005
R571 VTAIL.n638 VTAIL.n637 12.8005
R572 VTAIL.n597 VTAIL.n558 12.8005
R573 VTAIL.n592 VTAIL.n560 12.8005
R574 VTAIL.n532 VTAIL.n531 12.8005
R575 VTAIL.n491 VTAIL.n452 12.8005
R576 VTAIL.n486 VTAIL.n454 12.8005
R577 VTAIL.n424 VTAIL.n423 12.8005
R578 VTAIL.n383 VTAIL.n344 12.8005
R579 VTAIL.n378 VTAIL.n346 12.8005
R580 VTAIL.n803 VTAIL.n802 12.0247
R581 VTAIL.n812 VTAIL.n770 12.0247
R582 VTAIL.n848 VTAIL.n752 12.0247
R583 VTAIL.n55 VTAIL.n54 12.0247
R584 VTAIL.n64 VTAIL.n22 12.0247
R585 VTAIL.n100 VTAIL.n4 12.0247
R586 VTAIL.n161 VTAIL.n160 12.0247
R587 VTAIL.n170 VTAIL.n128 12.0247
R588 VTAIL.n206 VTAIL.n110 12.0247
R589 VTAIL.n269 VTAIL.n268 12.0247
R590 VTAIL.n278 VTAIL.n236 12.0247
R591 VTAIL.n314 VTAIL.n218 12.0247
R592 VTAIL.n742 VTAIL.n646 12.0247
R593 VTAIL.n706 VTAIL.n664 12.0247
R594 VTAIL.n697 VTAIL.n696 12.0247
R595 VTAIL.n634 VTAIL.n538 12.0247
R596 VTAIL.n598 VTAIL.n556 12.0247
R597 VTAIL.n589 VTAIL.n588 12.0247
R598 VTAIL.n528 VTAIL.n432 12.0247
R599 VTAIL.n492 VTAIL.n450 12.0247
R600 VTAIL.n483 VTAIL.n482 12.0247
R601 VTAIL.n420 VTAIL.n324 12.0247
R602 VTAIL.n384 VTAIL.n342 12.0247
R603 VTAIL.n375 VTAIL.n374 12.0247
R604 VTAIL.n798 VTAIL.n776 11.249
R605 VTAIL.n816 VTAIL.n815 11.249
R606 VTAIL.n847 VTAIL.n754 11.249
R607 VTAIL.n50 VTAIL.n28 11.249
R608 VTAIL.n68 VTAIL.n67 11.249
R609 VTAIL.n99 VTAIL.n6 11.249
R610 VTAIL.n156 VTAIL.n134 11.249
R611 VTAIL.n174 VTAIL.n173 11.249
R612 VTAIL.n205 VTAIL.n112 11.249
R613 VTAIL.n264 VTAIL.n242 11.249
R614 VTAIL.n282 VTAIL.n281 11.249
R615 VTAIL.n313 VTAIL.n220 11.249
R616 VTAIL.n741 VTAIL.n648 11.249
R617 VTAIL.n710 VTAIL.n709 11.249
R618 VTAIL.n693 VTAIL.n670 11.249
R619 VTAIL.n633 VTAIL.n540 11.249
R620 VTAIL.n602 VTAIL.n601 11.249
R621 VTAIL.n585 VTAIL.n562 11.249
R622 VTAIL.n527 VTAIL.n434 11.249
R623 VTAIL.n496 VTAIL.n495 11.249
R624 VTAIL.n479 VTAIL.n456 11.249
R625 VTAIL.n419 VTAIL.n326 11.249
R626 VTAIL.n388 VTAIL.n387 11.249
R627 VTAIL.n371 VTAIL.n348 11.249
R628 VTAIL.n785 VTAIL.n783 10.7239
R629 VTAIL.n37 VTAIL.n35 10.7239
R630 VTAIL.n143 VTAIL.n141 10.7239
R631 VTAIL.n251 VTAIL.n249 10.7239
R632 VTAIL.n680 VTAIL.n678 10.7239
R633 VTAIL.n572 VTAIL.n570 10.7239
R634 VTAIL.n466 VTAIL.n464 10.7239
R635 VTAIL.n358 VTAIL.n356 10.7239
R636 VTAIL.n797 VTAIL.n778 10.4732
R637 VTAIL.n819 VTAIL.n768 10.4732
R638 VTAIL.n844 VTAIL.n843 10.4732
R639 VTAIL.n49 VTAIL.n30 10.4732
R640 VTAIL.n71 VTAIL.n20 10.4732
R641 VTAIL.n96 VTAIL.n95 10.4732
R642 VTAIL.n155 VTAIL.n136 10.4732
R643 VTAIL.n177 VTAIL.n126 10.4732
R644 VTAIL.n202 VTAIL.n201 10.4732
R645 VTAIL.n263 VTAIL.n244 10.4732
R646 VTAIL.n285 VTAIL.n234 10.4732
R647 VTAIL.n310 VTAIL.n309 10.4732
R648 VTAIL.n738 VTAIL.n737 10.4732
R649 VTAIL.n713 VTAIL.n662 10.4732
R650 VTAIL.n692 VTAIL.n673 10.4732
R651 VTAIL.n630 VTAIL.n629 10.4732
R652 VTAIL.n605 VTAIL.n554 10.4732
R653 VTAIL.n584 VTAIL.n565 10.4732
R654 VTAIL.n524 VTAIL.n523 10.4732
R655 VTAIL.n499 VTAIL.n448 10.4732
R656 VTAIL.n478 VTAIL.n459 10.4732
R657 VTAIL.n416 VTAIL.n415 10.4732
R658 VTAIL.n391 VTAIL.n340 10.4732
R659 VTAIL.n370 VTAIL.n351 10.4732
R660 VTAIL.n794 VTAIL.n793 9.69747
R661 VTAIL.n820 VTAIL.n766 9.69747
R662 VTAIL.n840 VTAIL.n756 9.69747
R663 VTAIL.n46 VTAIL.n45 9.69747
R664 VTAIL.n72 VTAIL.n18 9.69747
R665 VTAIL.n92 VTAIL.n8 9.69747
R666 VTAIL.n152 VTAIL.n151 9.69747
R667 VTAIL.n178 VTAIL.n124 9.69747
R668 VTAIL.n198 VTAIL.n114 9.69747
R669 VTAIL.n260 VTAIL.n259 9.69747
R670 VTAIL.n286 VTAIL.n232 9.69747
R671 VTAIL.n306 VTAIL.n222 9.69747
R672 VTAIL.n734 VTAIL.n650 9.69747
R673 VTAIL.n714 VTAIL.n660 9.69747
R674 VTAIL.n689 VTAIL.n688 9.69747
R675 VTAIL.n626 VTAIL.n542 9.69747
R676 VTAIL.n606 VTAIL.n552 9.69747
R677 VTAIL.n581 VTAIL.n580 9.69747
R678 VTAIL.n520 VTAIL.n436 9.69747
R679 VTAIL.n500 VTAIL.n446 9.69747
R680 VTAIL.n475 VTAIL.n474 9.69747
R681 VTAIL.n412 VTAIL.n328 9.69747
R682 VTAIL.n392 VTAIL.n338 9.69747
R683 VTAIL.n367 VTAIL.n366 9.69747
R684 VTAIL.n854 VTAIL.n853 9.45567
R685 VTAIL.n106 VTAIL.n105 9.45567
R686 VTAIL.n212 VTAIL.n211 9.45567
R687 VTAIL.n320 VTAIL.n319 9.45567
R688 VTAIL.n748 VTAIL.n747 9.45567
R689 VTAIL.n640 VTAIL.n639 9.45567
R690 VTAIL.n534 VTAIL.n533 9.45567
R691 VTAIL.n426 VTAIL.n425 9.45567
R692 VTAIL.n829 VTAIL.n828 9.3005
R693 VTAIL.n764 VTAIL.n763 9.3005
R694 VTAIL.n823 VTAIL.n822 9.3005
R695 VTAIL.n821 VTAIL.n820 9.3005
R696 VTAIL.n768 VTAIL.n767 9.3005
R697 VTAIL.n815 VTAIL.n814 9.3005
R698 VTAIL.n813 VTAIL.n812 9.3005
R699 VTAIL.n772 VTAIL.n771 9.3005
R700 VTAIL.n787 VTAIL.n786 9.3005
R701 VTAIL.n789 VTAIL.n788 9.3005
R702 VTAIL.n780 VTAIL.n779 9.3005
R703 VTAIL.n795 VTAIL.n794 9.3005
R704 VTAIL.n797 VTAIL.n796 9.3005
R705 VTAIL.n776 VTAIL.n775 9.3005
R706 VTAIL.n804 VTAIL.n803 9.3005
R707 VTAIL.n806 VTAIL.n805 9.3005
R708 VTAIL.n831 VTAIL.n830 9.3005
R709 VTAIL.n760 VTAIL.n759 9.3005
R710 VTAIL.n837 VTAIL.n836 9.3005
R711 VTAIL.n839 VTAIL.n838 9.3005
R712 VTAIL.n756 VTAIL.n755 9.3005
R713 VTAIL.n845 VTAIL.n844 9.3005
R714 VTAIL.n847 VTAIL.n846 9.3005
R715 VTAIL.n752 VTAIL.n751 9.3005
R716 VTAIL.n853 VTAIL.n852 9.3005
R717 VTAIL.n81 VTAIL.n80 9.3005
R718 VTAIL.n16 VTAIL.n15 9.3005
R719 VTAIL.n75 VTAIL.n74 9.3005
R720 VTAIL.n73 VTAIL.n72 9.3005
R721 VTAIL.n20 VTAIL.n19 9.3005
R722 VTAIL.n67 VTAIL.n66 9.3005
R723 VTAIL.n65 VTAIL.n64 9.3005
R724 VTAIL.n24 VTAIL.n23 9.3005
R725 VTAIL.n39 VTAIL.n38 9.3005
R726 VTAIL.n41 VTAIL.n40 9.3005
R727 VTAIL.n32 VTAIL.n31 9.3005
R728 VTAIL.n47 VTAIL.n46 9.3005
R729 VTAIL.n49 VTAIL.n48 9.3005
R730 VTAIL.n28 VTAIL.n27 9.3005
R731 VTAIL.n56 VTAIL.n55 9.3005
R732 VTAIL.n58 VTAIL.n57 9.3005
R733 VTAIL.n83 VTAIL.n82 9.3005
R734 VTAIL.n12 VTAIL.n11 9.3005
R735 VTAIL.n89 VTAIL.n88 9.3005
R736 VTAIL.n91 VTAIL.n90 9.3005
R737 VTAIL.n8 VTAIL.n7 9.3005
R738 VTAIL.n97 VTAIL.n96 9.3005
R739 VTAIL.n99 VTAIL.n98 9.3005
R740 VTAIL.n4 VTAIL.n3 9.3005
R741 VTAIL.n105 VTAIL.n104 9.3005
R742 VTAIL.n187 VTAIL.n186 9.3005
R743 VTAIL.n122 VTAIL.n121 9.3005
R744 VTAIL.n181 VTAIL.n180 9.3005
R745 VTAIL.n179 VTAIL.n178 9.3005
R746 VTAIL.n126 VTAIL.n125 9.3005
R747 VTAIL.n173 VTAIL.n172 9.3005
R748 VTAIL.n171 VTAIL.n170 9.3005
R749 VTAIL.n130 VTAIL.n129 9.3005
R750 VTAIL.n145 VTAIL.n144 9.3005
R751 VTAIL.n147 VTAIL.n146 9.3005
R752 VTAIL.n138 VTAIL.n137 9.3005
R753 VTAIL.n153 VTAIL.n152 9.3005
R754 VTAIL.n155 VTAIL.n154 9.3005
R755 VTAIL.n134 VTAIL.n133 9.3005
R756 VTAIL.n162 VTAIL.n161 9.3005
R757 VTAIL.n164 VTAIL.n163 9.3005
R758 VTAIL.n189 VTAIL.n188 9.3005
R759 VTAIL.n118 VTAIL.n117 9.3005
R760 VTAIL.n195 VTAIL.n194 9.3005
R761 VTAIL.n197 VTAIL.n196 9.3005
R762 VTAIL.n114 VTAIL.n113 9.3005
R763 VTAIL.n203 VTAIL.n202 9.3005
R764 VTAIL.n205 VTAIL.n204 9.3005
R765 VTAIL.n110 VTAIL.n109 9.3005
R766 VTAIL.n211 VTAIL.n210 9.3005
R767 VTAIL.n295 VTAIL.n294 9.3005
R768 VTAIL.n230 VTAIL.n229 9.3005
R769 VTAIL.n289 VTAIL.n288 9.3005
R770 VTAIL.n287 VTAIL.n286 9.3005
R771 VTAIL.n234 VTAIL.n233 9.3005
R772 VTAIL.n281 VTAIL.n280 9.3005
R773 VTAIL.n279 VTAIL.n278 9.3005
R774 VTAIL.n238 VTAIL.n237 9.3005
R775 VTAIL.n253 VTAIL.n252 9.3005
R776 VTAIL.n255 VTAIL.n254 9.3005
R777 VTAIL.n246 VTAIL.n245 9.3005
R778 VTAIL.n261 VTAIL.n260 9.3005
R779 VTAIL.n263 VTAIL.n262 9.3005
R780 VTAIL.n242 VTAIL.n241 9.3005
R781 VTAIL.n270 VTAIL.n269 9.3005
R782 VTAIL.n272 VTAIL.n271 9.3005
R783 VTAIL.n297 VTAIL.n296 9.3005
R784 VTAIL.n226 VTAIL.n225 9.3005
R785 VTAIL.n303 VTAIL.n302 9.3005
R786 VTAIL.n305 VTAIL.n304 9.3005
R787 VTAIL.n222 VTAIL.n221 9.3005
R788 VTAIL.n311 VTAIL.n310 9.3005
R789 VTAIL.n313 VTAIL.n312 9.3005
R790 VTAIL.n218 VTAIL.n217 9.3005
R791 VTAIL.n319 VTAIL.n318 9.3005
R792 VTAIL.n682 VTAIL.n681 9.3005
R793 VTAIL.n684 VTAIL.n683 9.3005
R794 VTAIL.n675 VTAIL.n674 9.3005
R795 VTAIL.n690 VTAIL.n689 9.3005
R796 VTAIL.n692 VTAIL.n691 9.3005
R797 VTAIL.n670 VTAIL.n669 9.3005
R798 VTAIL.n698 VTAIL.n697 9.3005
R799 VTAIL.n700 VTAIL.n699 9.3005
R800 VTAIL.n654 VTAIL.n653 9.3005
R801 VTAIL.n731 VTAIL.n730 9.3005
R802 VTAIL.n733 VTAIL.n732 9.3005
R803 VTAIL.n650 VTAIL.n649 9.3005
R804 VTAIL.n739 VTAIL.n738 9.3005
R805 VTAIL.n741 VTAIL.n740 9.3005
R806 VTAIL.n646 VTAIL.n645 9.3005
R807 VTAIL.n747 VTAIL.n746 9.3005
R808 VTAIL.n725 VTAIL.n724 9.3005
R809 VTAIL.n723 VTAIL.n722 9.3005
R810 VTAIL.n658 VTAIL.n657 9.3005
R811 VTAIL.n717 VTAIL.n716 9.3005
R812 VTAIL.n715 VTAIL.n714 9.3005
R813 VTAIL.n662 VTAIL.n661 9.3005
R814 VTAIL.n709 VTAIL.n708 9.3005
R815 VTAIL.n707 VTAIL.n706 9.3005
R816 VTAIL.n666 VTAIL.n665 9.3005
R817 VTAIL.n574 VTAIL.n573 9.3005
R818 VTAIL.n576 VTAIL.n575 9.3005
R819 VTAIL.n567 VTAIL.n566 9.3005
R820 VTAIL.n582 VTAIL.n581 9.3005
R821 VTAIL.n584 VTAIL.n583 9.3005
R822 VTAIL.n562 VTAIL.n561 9.3005
R823 VTAIL.n590 VTAIL.n589 9.3005
R824 VTAIL.n592 VTAIL.n591 9.3005
R825 VTAIL.n546 VTAIL.n545 9.3005
R826 VTAIL.n623 VTAIL.n622 9.3005
R827 VTAIL.n625 VTAIL.n624 9.3005
R828 VTAIL.n542 VTAIL.n541 9.3005
R829 VTAIL.n631 VTAIL.n630 9.3005
R830 VTAIL.n633 VTAIL.n632 9.3005
R831 VTAIL.n538 VTAIL.n537 9.3005
R832 VTAIL.n639 VTAIL.n638 9.3005
R833 VTAIL.n617 VTAIL.n616 9.3005
R834 VTAIL.n615 VTAIL.n614 9.3005
R835 VTAIL.n550 VTAIL.n549 9.3005
R836 VTAIL.n609 VTAIL.n608 9.3005
R837 VTAIL.n607 VTAIL.n606 9.3005
R838 VTAIL.n554 VTAIL.n553 9.3005
R839 VTAIL.n601 VTAIL.n600 9.3005
R840 VTAIL.n599 VTAIL.n598 9.3005
R841 VTAIL.n558 VTAIL.n557 9.3005
R842 VTAIL.n468 VTAIL.n467 9.3005
R843 VTAIL.n470 VTAIL.n469 9.3005
R844 VTAIL.n461 VTAIL.n460 9.3005
R845 VTAIL.n476 VTAIL.n475 9.3005
R846 VTAIL.n478 VTAIL.n477 9.3005
R847 VTAIL.n456 VTAIL.n455 9.3005
R848 VTAIL.n484 VTAIL.n483 9.3005
R849 VTAIL.n486 VTAIL.n485 9.3005
R850 VTAIL.n440 VTAIL.n439 9.3005
R851 VTAIL.n517 VTAIL.n516 9.3005
R852 VTAIL.n519 VTAIL.n518 9.3005
R853 VTAIL.n436 VTAIL.n435 9.3005
R854 VTAIL.n525 VTAIL.n524 9.3005
R855 VTAIL.n527 VTAIL.n526 9.3005
R856 VTAIL.n432 VTAIL.n431 9.3005
R857 VTAIL.n533 VTAIL.n532 9.3005
R858 VTAIL.n511 VTAIL.n510 9.3005
R859 VTAIL.n509 VTAIL.n508 9.3005
R860 VTAIL.n444 VTAIL.n443 9.3005
R861 VTAIL.n503 VTAIL.n502 9.3005
R862 VTAIL.n501 VTAIL.n500 9.3005
R863 VTAIL.n448 VTAIL.n447 9.3005
R864 VTAIL.n495 VTAIL.n494 9.3005
R865 VTAIL.n493 VTAIL.n492 9.3005
R866 VTAIL.n452 VTAIL.n451 9.3005
R867 VTAIL.n360 VTAIL.n359 9.3005
R868 VTAIL.n362 VTAIL.n361 9.3005
R869 VTAIL.n353 VTAIL.n352 9.3005
R870 VTAIL.n368 VTAIL.n367 9.3005
R871 VTAIL.n370 VTAIL.n369 9.3005
R872 VTAIL.n348 VTAIL.n347 9.3005
R873 VTAIL.n376 VTAIL.n375 9.3005
R874 VTAIL.n378 VTAIL.n377 9.3005
R875 VTAIL.n332 VTAIL.n331 9.3005
R876 VTAIL.n409 VTAIL.n408 9.3005
R877 VTAIL.n411 VTAIL.n410 9.3005
R878 VTAIL.n328 VTAIL.n327 9.3005
R879 VTAIL.n417 VTAIL.n416 9.3005
R880 VTAIL.n419 VTAIL.n418 9.3005
R881 VTAIL.n324 VTAIL.n323 9.3005
R882 VTAIL.n425 VTAIL.n424 9.3005
R883 VTAIL.n403 VTAIL.n402 9.3005
R884 VTAIL.n401 VTAIL.n400 9.3005
R885 VTAIL.n336 VTAIL.n335 9.3005
R886 VTAIL.n395 VTAIL.n394 9.3005
R887 VTAIL.n393 VTAIL.n392 9.3005
R888 VTAIL.n340 VTAIL.n339 9.3005
R889 VTAIL.n387 VTAIL.n386 9.3005
R890 VTAIL.n385 VTAIL.n384 9.3005
R891 VTAIL.n344 VTAIL.n343 9.3005
R892 VTAIL.n790 VTAIL.n780 8.92171
R893 VTAIL.n824 VTAIL.n823 8.92171
R894 VTAIL.n839 VTAIL.n758 8.92171
R895 VTAIL.n42 VTAIL.n32 8.92171
R896 VTAIL.n76 VTAIL.n75 8.92171
R897 VTAIL.n91 VTAIL.n10 8.92171
R898 VTAIL.n148 VTAIL.n138 8.92171
R899 VTAIL.n182 VTAIL.n181 8.92171
R900 VTAIL.n197 VTAIL.n116 8.92171
R901 VTAIL.n256 VTAIL.n246 8.92171
R902 VTAIL.n290 VTAIL.n289 8.92171
R903 VTAIL.n305 VTAIL.n224 8.92171
R904 VTAIL.n733 VTAIL.n652 8.92171
R905 VTAIL.n718 VTAIL.n717 8.92171
R906 VTAIL.n685 VTAIL.n675 8.92171
R907 VTAIL.n625 VTAIL.n544 8.92171
R908 VTAIL.n610 VTAIL.n609 8.92171
R909 VTAIL.n577 VTAIL.n567 8.92171
R910 VTAIL.n519 VTAIL.n438 8.92171
R911 VTAIL.n504 VTAIL.n503 8.92171
R912 VTAIL.n471 VTAIL.n461 8.92171
R913 VTAIL.n411 VTAIL.n330 8.92171
R914 VTAIL.n396 VTAIL.n395 8.92171
R915 VTAIL.n363 VTAIL.n353 8.92171
R916 VTAIL.n789 VTAIL.n782 8.14595
R917 VTAIL.n827 VTAIL.n764 8.14595
R918 VTAIL.n836 VTAIL.n835 8.14595
R919 VTAIL.n41 VTAIL.n34 8.14595
R920 VTAIL.n79 VTAIL.n16 8.14595
R921 VTAIL.n88 VTAIL.n87 8.14595
R922 VTAIL.n147 VTAIL.n140 8.14595
R923 VTAIL.n185 VTAIL.n122 8.14595
R924 VTAIL.n194 VTAIL.n193 8.14595
R925 VTAIL.n255 VTAIL.n248 8.14595
R926 VTAIL.n293 VTAIL.n230 8.14595
R927 VTAIL.n302 VTAIL.n301 8.14595
R928 VTAIL.n730 VTAIL.n729 8.14595
R929 VTAIL.n721 VTAIL.n658 8.14595
R930 VTAIL.n684 VTAIL.n677 8.14595
R931 VTAIL.n622 VTAIL.n621 8.14595
R932 VTAIL.n613 VTAIL.n550 8.14595
R933 VTAIL.n576 VTAIL.n569 8.14595
R934 VTAIL.n516 VTAIL.n515 8.14595
R935 VTAIL.n507 VTAIL.n444 8.14595
R936 VTAIL.n470 VTAIL.n463 8.14595
R937 VTAIL.n408 VTAIL.n407 8.14595
R938 VTAIL.n399 VTAIL.n336 8.14595
R939 VTAIL.n362 VTAIL.n355 8.14595
R940 VTAIL.n854 VTAIL.n750 7.75445
R941 VTAIL.n106 VTAIL.n2 7.75445
R942 VTAIL.n212 VTAIL.n108 7.75445
R943 VTAIL.n320 VTAIL.n216 7.75445
R944 VTAIL.n748 VTAIL.n644 7.75445
R945 VTAIL.n640 VTAIL.n536 7.75445
R946 VTAIL.n534 VTAIL.n430 7.75445
R947 VTAIL.n426 VTAIL.n322 7.75445
R948 VTAIL.n786 VTAIL.n785 7.3702
R949 VTAIL.n828 VTAIL.n762 7.3702
R950 VTAIL.n832 VTAIL.n760 7.3702
R951 VTAIL.n38 VTAIL.n37 7.3702
R952 VTAIL.n80 VTAIL.n14 7.3702
R953 VTAIL.n84 VTAIL.n12 7.3702
R954 VTAIL.n144 VTAIL.n143 7.3702
R955 VTAIL.n186 VTAIL.n120 7.3702
R956 VTAIL.n190 VTAIL.n118 7.3702
R957 VTAIL.n252 VTAIL.n251 7.3702
R958 VTAIL.n294 VTAIL.n228 7.3702
R959 VTAIL.n298 VTAIL.n226 7.3702
R960 VTAIL.n726 VTAIL.n654 7.3702
R961 VTAIL.n722 VTAIL.n656 7.3702
R962 VTAIL.n681 VTAIL.n680 7.3702
R963 VTAIL.n618 VTAIL.n546 7.3702
R964 VTAIL.n614 VTAIL.n548 7.3702
R965 VTAIL.n573 VTAIL.n572 7.3702
R966 VTAIL.n512 VTAIL.n440 7.3702
R967 VTAIL.n508 VTAIL.n442 7.3702
R968 VTAIL.n467 VTAIL.n466 7.3702
R969 VTAIL.n404 VTAIL.n332 7.3702
R970 VTAIL.n400 VTAIL.n334 7.3702
R971 VTAIL.n359 VTAIL.n358 7.3702
R972 VTAIL.n831 VTAIL.n762 6.59444
R973 VTAIL.n832 VTAIL.n831 6.59444
R974 VTAIL.n83 VTAIL.n14 6.59444
R975 VTAIL.n84 VTAIL.n83 6.59444
R976 VTAIL.n189 VTAIL.n120 6.59444
R977 VTAIL.n190 VTAIL.n189 6.59444
R978 VTAIL.n297 VTAIL.n228 6.59444
R979 VTAIL.n298 VTAIL.n297 6.59444
R980 VTAIL.n726 VTAIL.n725 6.59444
R981 VTAIL.n725 VTAIL.n656 6.59444
R982 VTAIL.n618 VTAIL.n617 6.59444
R983 VTAIL.n617 VTAIL.n548 6.59444
R984 VTAIL.n512 VTAIL.n511 6.59444
R985 VTAIL.n511 VTAIL.n442 6.59444
R986 VTAIL.n404 VTAIL.n403 6.59444
R987 VTAIL.n403 VTAIL.n334 6.59444
R988 VTAIL.n852 VTAIL.n750 6.08283
R989 VTAIL.n104 VTAIL.n2 6.08283
R990 VTAIL.n210 VTAIL.n108 6.08283
R991 VTAIL.n318 VTAIL.n216 6.08283
R992 VTAIL.n746 VTAIL.n644 6.08283
R993 VTAIL.n638 VTAIL.n536 6.08283
R994 VTAIL.n532 VTAIL.n430 6.08283
R995 VTAIL.n424 VTAIL.n322 6.08283
R996 VTAIL.n786 VTAIL.n782 5.81868
R997 VTAIL.n828 VTAIL.n827 5.81868
R998 VTAIL.n835 VTAIL.n760 5.81868
R999 VTAIL.n38 VTAIL.n34 5.81868
R1000 VTAIL.n80 VTAIL.n79 5.81868
R1001 VTAIL.n87 VTAIL.n12 5.81868
R1002 VTAIL.n144 VTAIL.n140 5.81868
R1003 VTAIL.n186 VTAIL.n185 5.81868
R1004 VTAIL.n193 VTAIL.n118 5.81868
R1005 VTAIL.n252 VTAIL.n248 5.81868
R1006 VTAIL.n294 VTAIL.n293 5.81868
R1007 VTAIL.n301 VTAIL.n226 5.81868
R1008 VTAIL.n729 VTAIL.n654 5.81868
R1009 VTAIL.n722 VTAIL.n721 5.81868
R1010 VTAIL.n681 VTAIL.n677 5.81868
R1011 VTAIL.n621 VTAIL.n546 5.81868
R1012 VTAIL.n614 VTAIL.n613 5.81868
R1013 VTAIL.n573 VTAIL.n569 5.81868
R1014 VTAIL.n515 VTAIL.n440 5.81868
R1015 VTAIL.n508 VTAIL.n507 5.81868
R1016 VTAIL.n467 VTAIL.n463 5.81868
R1017 VTAIL.n407 VTAIL.n332 5.81868
R1018 VTAIL.n400 VTAIL.n399 5.81868
R1019 VTAIL.n359 VTAIL.n355 5.81868
R1020 VTAIL.n790 VTAIL.n789 5.04292
R1021 VTAIL.n824 VTAIL.n764 5.04292
R1022 VTAIL.n836 VTAIL.n758 5.04292
R1023 VTAIL.n42 VTAIL.n41 5.04292
R1024 VTAIL.n76 VTAIL.n16 5.04292
R1025 VTAIL.n88 VTAIL.n10 5.04292
R1026 VTAIL.n148 VTAIL.n147 5.04292
R1027 VTAIL.n182 VTAIL.n122 5.04292
R1028 VTAIL.n194 VTAIL.n116 5.04292
R1029 VTAIL.n256 VTAIL.n255 5.04292
R1030 VTAIL.n290 VTAIL.n230 5.04292
R1031 VTAIL.n302 VTAIL.n224 5.04292
R1032 VTAIL.n730 VTAIL.n652 5.04292
R1033 VTAIL.n718 VTAIL.n658 5.04292
R1034 VTAIL.n685 VTAIL.n684 5.04292
R1035 VTAIL.n622 VTAIL.n544 5.04292
R1036 VTAIL.n610 VTAIL.n550 5.04292
R1037 VTAIL.n577 VTAIL.n576 5.04292
R1038 VTAIL.n516 VTAIL.n438 5.04292
R1039 VTAIL.n504 VTAIL.n444 5.04292
R1040 VTAIL.n471 VTAIL.n470 5.04292
R1041 VTAIL.n408 VTAIL.n330 5.04292
R1042 VTAIL.n396 VTAIL.n336 5.04292
R1043 VTAIL.n363 VTAIL.n362 5.04292
R1044 VTAIL.n793 VTAIL.n780 4.26717
R1045 VTAIL.n823 VTAIL.n766 4.26717
R1046 VTAIL.n840 VTAIL.n839 4.26717
R1047 VTAIL.n45 VTAIL.n32 4.26717
R1048 VTAIL.n75 VTAIL.n18 4.26717
R1049 VTAIL.n92 VTAIL.n91 4.26717
R1050 VTAIL.n151 VTAIL.n138 4.26717
R1051 VTAIL.n181 VTAIL.n124 4.26717
R1052 VTAIL.n198 VTAIL.n197 4.26717
R1053 VTAIL.n259 VTAIL.n246 4.26717
R1054 VTAIL.n289 VTAIL.n232 4.26717
R1055 VTAIL.n306 VTAIL.n305 4.26717
R1056 VTAIL.n734 VTAIL.n733 4.26717
R1057 VTAIL.n717 VTAIL.n660 4.26717
R1058 VTAIL.n688 VTAIL.n675 4.26717
R1059 VTAIL.n626 VTAIL.n625 4.26717
R1060 VTAIL.n609 VTAIL.n552 4.26717
R1061 VTAIL.n580 VTAIL.n567 4.26717
R1062 VTAIL.n520 VTAIL.n519 4.26717
R1063 VTAIL.n503 VTAIL.n446 4.26717
R1064 VTAIL.n474 VTAIL.n461 4.26717
R1065 VTAIL.n412 VTAIL.n411 4.26717
R1066 VTAIL.n395 VTAIL.n338 4.26717
R1067 VTAIL.n366 VTAIL.n353 4.26717
R1068 VTAIL.n794 VTAIL.n778 3.49141
R1069 VTAIL.n820 VTAIL.n819 3.49141
R1070 VTAIL.n843 VTAIL.n756 3.49141
R1071 VTAIL.n46 VTAIL.n30 3.49141
R1072 VTAIL.n72 VTAIL.n71 3.49141
R1073 VTAIL.n95 VTAIL.n8 3.49141
R1074 VTAIL.n152 VTAIL.n136 3.49141
R1075 VTAIL.n178 VTAIL.n177 3.49141
R1076 VTAIL.n201 VTAIL.n114 3.49141
R1077 VTAIL.n260 VTAIL.n244 3.49141
R1078 VTAIL.n286 VTAIL.n285 3.49141
R1079 VTAIL.n309 VTAIL.n222 3.49141
R1080 VTAIL.n737 VTAIL.n650 3.49141
R1081 VTAIL.n714 VTAIL.n713 3.49141
R1082 VTAIL.n689 VTAIL.n673 3.49141
R1083 VTAIL.n629 VTAIL.n542 3.49141
R1084 VTAIL.n606 VTAIL.n605 3.49141
R1085 VTAIL.n581 VTAIL.n565 3.49141
R1086 VTAIL.n523 VTAIL.n436 3.49141
R1087 VTAIL.n500 VTAIL.n499 3.49141
R1088 VTAIL.n475 VTAIL.n459 3.49141
R1089 VTAIL.n415 VTAIL.n328 3.49141
R1090 VTAIL.n392 VTAIL.n391 3.49141
R1091 VTAIL.n367 VTAIL.n351 3.49141
R1092 VTAIL.n798 VTAIL.n797 2.71565
R1093 VTAIL.n816 VTAIL.n768 2.71565
R1094 VTAIL.n844 VTAIL.n754 2.71565
R1095 VTAIL.n50 VTAIL.n49 2.71565
R1096 VTAIL.n68 VTAIL.n20 2.71565
R1097 VTAIL.n96 VTAIL.n6 2.71565
R1098 VTAIL.n156 VTAIL.n155 2.71565
R1099 VTAIL.n174 VTAIL.n126 2.71565
R1100 VTAIL.n202 VTAIL.n112 2.71565
R1101 VTAIL.n264 VTAIL.n263 2.71565
R1102 VTAIL.n282 VTAIL.n234 2.71565
R1103 VTAIL.n310 VTAIL.n220 2.71565
R1104 VTAIL.n738 VTAIL.n648 2.71565
R1105 VTAIL.n710 VTAIL.n662 2.71565
R1106 VTAIL.n693 VTAIL.n692 2.71565
R1107 VTAIL.n630 VTAIL.n540 2.71565
R1108 VTAIL.n602 VTAIL.n554 2.71565
R1109 VTAIL.n585 VTAIL.n584 2.71565
R1110 VTAIL.n524 VTAIL.n434 2.71565
R1111 VTAIL.n496 VTAIL.n448 2.71565
R1112 VTAIL.n479 VTAIL.n478 2.71565
R1113 VTAIL.n416 VTAIL.n326 2.71565
R1114 VTAIL.n388 VTAIL.n340 2.71565
R1115 VTAIL.n371 VTAIL.n370 2.71565
R1116 VTAIL.n682 VTAIL.n678 2.41282
R1117 VTAIL.n574 VTAIL.n570 2.41282
R1118 VTAIL.n468 VTAIL.n464 2.41282
R1119 VTAIL.n360 VTAIL.n356 2.41282
R1120 VTAIL.n787 VTAIL.n783 2.41282
R1121 VTAIL.n39 VTAIL.n35 2.41282
R1122 VTAIL.n145 VTAIL.n141 2.41282
R1123 VTAIL.n253 VTAIL.n249 2.41282
R1124 VTAIL.n429 VTAIL.n427 2.31947
R1125 VTAIL.n535 VTAIL.n429 2.31947
R1126 VTAIL.n643 VTAIL.n641 2.31947
R1127 VTAIL.n749 VTAIL.n643 2.31947
R1128 VTAIL.n321 VTAIL.n215 2.31947
R1129 VTAIL.n215 VTAIL.n213 2.31947
R1130 VTAIL.n107 VTAIL.n1 2.31947
R1131 VTAIL VTAIL.n855 2.26128
R1132 VTAIL.n802 VTAIL.n776 1.93989
R1133 VTAIL.n815 VTAIL.n770 1.93989
R1134 VTAIL.n848 VTAIL.n847 1.93989
R1135 VTAIL.n54 VTAIL.n28 1.93989
R1136 VTAIL.n67 VTAIL.n22 1.93989
R1137 VTAIL.n100 VTAIL.n99 1.93989
R1138 VTAIL.n160 VTAIL.n134 1.93989
R1139 VTAIL.n173 VTAIL.n128 1.93989
R1140 VTAIL.n206 VTAIL.n205 1.93989
R1141 VTAIL.n268 VTAIL.n242 1.93989
R1142 VTAIL.n281 VTAIL.n236 1.93989
R1143 VTAIL.n314 VTAIL.n313 1.93989
R1144 VTAIL.n742 VTAIL.n741 1.93989
R1145 VTAIL.n709 VTAIL.n664 1.93989
R1146 VTAIL.n696 VTAIL.n670 1.93989
R1147 VTAIL.n634 VTAIL.n633 1.93989
R1148 VTAIL.n601 VTAIL.n556 1.93989
R1149 VTAIL.n588 VTAIL.n562 1.93989
R1150 VTAIL.n528 VTAIL.n527 1.93989
R1151 VTAIL.n495 VTAIL.n450 1.93989
R1152 VTAIL.n482 VTAIL.n456 1.93989
R1153 VTAIL.n420 VTAIL.n419 1.93989
R1154 VTAIL.n387 VTAIL.n342 1.93989
R1155 VTAIL.n374 VTAIL.n348 1.93989
R1156 VTAIL.n0 VTAIL.t6 1.67257
R1157 VTAIL.n0 VTAIL.t5 1.67257
R1158 VTAIL.n214 VTAIL.t13 1.67257
R1159 VTAIL.n214 VTAIL.t15 1.67257
R1160 VTAIL.n642 VTAIL.t9 1.67257
R1161 VTAIL.n642 VTAIL.t12 1.67257
R1162 VTAIL.n428 VTAIL.t2 1.67257
R1163 VTAIL.n428 VTAIL.t3 1.67257
R1164 VTAIL.n803 VTAIL.n774 1.16414
R1165 VTAIL.n812 VTAIL.n811 1.16414
R1166 VTAIL.n851 VTAIL.n752 1.16414
R1167 VTAIL.n55 VTAIL.n26 1.16414
R1168 VTAIL.n64 VTAIL.n63 1.16414
R1169 VTAIL.n103 VTAIL.n4 1.16414
R1170 VTAIL.n161 VTAIL.n132 1.16414
R1171 VTAIL.n170 VTAIL.n169 1.16414
R1172 VTAIL.n209 VTAIL.n110 1.16414
R1173 VTAIL.n269 VTAIL.n240 1.16414
R1174 VTAIL.n278 VTAIL.n277 1.16414
R1175 VTAIL.n317 VTAIL.n218 1.16414
R1176 VTAIL.n745 VTAIL.n646 1.16414
R1177 VTAIL.n706 VTAIL.n705 1.16414
R1178 VTAIL.n697 VTAIL.n668 1.16414
R1179 VTAIL.n637 VTAIL.n538 1.16414
R1180 VTAIL.n598 VTAIL.n597 1.16414
R1181 VTAIL.n589 VTAIL.n560 1.16414
R1182 VTAIL.n531 VTAIL.n432 1.16414
R1183 VTAIL.n492 VTAIL.n491 1.16414
R1184 VTAIL.n483 VTAIL.n454 1.16414
R1185 VTAIL.n423 VTAIL.n324 1.16414
R1186 VTAIL.n384 VTAIL.n383 1.16414
R1187 VTAIL.n375 VTAIL.n346 1.16414
R1188 VTAIL.n641 VTAIL.n535 0.470328
R1189 VTAIL.n213 VTAIL.n107 0.470328
R1190 VTAIL.n807 VTAIL.n806 0.388379
R1191 VTAIL.n808 VTAIL.n772 0.388379
R1192 VTAIL.n59 VTAIL.n58 0.388379
R1193 VTAIL.n60 VTAIL.n24 0.388379
R1194 VTAIL.n165 VTAIL.n164 0.388379
R1195 VTAIL.n166 VTAIL.n130 0.388379
R1196 VTAIL.n273 VTAIL.n272 0.388379
R1197 VTAIL.n274 VTAIL.n238 0.388379
R1198 VTAIL.n702 VTAIL.n666 0.388379
R1199 VTAIL.n701 VTAIL.n700 0.388379
R1200 VTAIL.n594 VTAIL.n558 0.388379
R1201 VTAIL.n593 VTAIL.n592 0.388379
R1202 VTAIL.n488 VTAIL.n452 0.388379
R1203 VTAIL.n487 VTAIL.n486 0.388379
R1204 VTAIL.n380 VTAIL.n344 0.388379
R1205 VTAIL.n379 VTAIL.n378 0.388379
R1206 VTAIL.n788 VTAIL.n787 0.155672
R1207 VTAIL.n788 VTAIL.n779 0.155672
R1208 VTAIL.n795 VTAIL.n779 0.155672
R1209 VTAIL.n796 VTAIL.n795 0.155672
R1210 VTAIL.n796 VTAIL.n775 0.155672
R1211 VTAIL.n804 VTAIL.n775 0.155672
R1212 VTAIL.n805 VTAIL.n804 0.155672
R1213 VTAIL.n805 VTAIL.n771 0.155672
R1214 VTAIL.n813 VTAIL.n771 0.155672
R1215 VTAIL.n814 VTAIL.n813 0.155672
R1216 VTAIL.n814 VTAIL.n767 0.155672
R1217 VTAIL.n821 VTAIL.n767 0.155672
R1218 VTAIL.n822 VTAIL.n821 0.155672
R1219 VTAIL.n822 VTAIL.n763 0.155672
R1220 VTAIL.n829 VTAIL.n763 0.155672
R1221 VTAIL.n830 VTAIL.n829 0.155672
R1222 VTAIL.n830 VTAIL.n759 0.155672
R1223 VTAIL.n837 VTAIL.n759 0.155672
R1224 VTAIL.n838 VTAIL.n837 0.155672
R1225 VTAIL.n838 VTAIL.n755 0.155672
R1226 VTAIL.n845 VTAIL.n755 0.155672
R1227 VTAIL.n846 VTAIL.n845 0.155672
R1228 VTAIL.n846 VTAIL.n751 0.155672
R1229 VTAIL.n853 VTAIL.n751 0.155672
R1230 VTAIL.n40 VTAIL.n39 0.155672
R1231 VTAIL.n40 VTAIL.n31 0.155672
R1232 VTAIL.n47 VTAIL.n31 0.155672
R1233 VTAIL.n48 VTAIL.n47 0.155672
R1234 VTAIL.n48 VTAIL.n27 0.155672
R1235 VTAIL.n56 VTAIL.n27 0.155672
R1236 VTAIL.n57 VTAIL.n56 0.155672
R1237 VTAIL.n57 VTAIL.n23 0.155672
R1238 VTAIL.n65 VTAIL.n23 0.155672
R1239 VTAIL.n66 VTAIL.n65 0.155672
R1240 VTAIL.n66 VTAIL.n19 0.155672
R1241 VTAIL.n73 VTAIL.n19 0.155672
R1242 VTAIL.n74 VTAIL.n73 0.155672
R1243 VTAIL.n74 VTAIL.n15 0.155672
R1244 VTAIL.n81 VTAIL.n15 0.155672
R1245 VTAIL.n82 VTAIL.n81 0.155672
R1246 VTAIL.n82 VTAIL.n11 0.155672
R1247 VTAIL.n89 VTAIL.n11 0.155672
R1248 VTAIL.n90 VTAIL.n89 0.155672
R1249 VTAIL.n90 VTAIL.n7 0.155672
R1250 VTAIL.n97 VTAIL.n7 0.155672
R1251 VTAIL.n98 VTAIL.n97 0.155672
R1252 VTAIL.n98 VTAIL.n3 0.155672
R1253 VTAIL.n105 VTAIL.n3 0.155672
R1254 VTAIL.n146 VTAIL.n145 0.155672
R1255 VTAIL.n146 VTAIL.n137 0.155672
R1256 VTAIL.n153 VTAIL.n137 0.155672
R1257 VTAIL.n154 VTAIL.n153 0.155672
R1258 VTAIL.n154 VTAIL.n133 0.155672
R1259 VTAIL.n162 VTAIL.n133 0.155672
R1260 VTAIL.n163 VTAIL.n162 0.155672
R1261 VTAIL.n163 VTAIL.n129 0.155672
R1262 VTAIL.n171 VTAIL.n129 0.155672
R1263 VTAIL.n172 VTAIL.n171 0.155672
R1264 VTAIL.n172 VTAIL.n125 0.155672
R1265 VTAIL.n179 VTAIL.n125 0.155672
R1266 VTAIL.n180 VTAIL.n179 0.155672
R1267 VTAIL.n180 VTAIL.n121 0.155672
R1268 VTAIL.n187 VTAIL.n121 0.155672
R1269 VTAIL.n188 VTAIL.n187 0.155672
R1270 VTAIL.n188 VTAIL.n117 0.155672
R1271 VTAIL.n195 VTAIL.n117 0.155672
R1272 VTAIL.n196 VTAIL.n195 0.155672
R1273 VTAIL.n196 VTAIL.n113 0.155672
R1274 VTAIL.n203 VTAIL.n113 0.155672
R1275 VTAIL.n204 VTAIL.n203 0.155672
R1276 VTAIL.n204 VTAIL.n109 0.155672
R1277 VTAIL.n211 VTAIL.n109 0.155672
R1278 VTAIL.n254 VTAIL.n253 0.155672
R1279 VTAIL.n254 VTAIL.n245 0.155672
R1280 VTAIL.n261 VTAIL.n245 0.155672
R1281 VTAIL.n262 VTAIL.n261 0.155672
R1282 VTAIL.n262 VTAIL.n241 0.155672
R1283 VTAIL.n270 VTAIL.n241 0.155672
R1284 VTAIL.n271 VTAIL.n270 0.155672
R1285 VTAIL.n271 VTAIL.n237 0.155672
R1286 VTAIL.n279 VTAIL.n237 0.155672
R1287 VTAIL.n280 VTAIL.n279 0.155672
R1288 VTAIL.n280 VTAIL.n233 0.155672
R1289 VTAIL.n287 VTAIL.n233 0.155672
R1290 VTAIL.n288 VTAIL.n287 0.155672
R1291 VTAIL.n288 VTAIL.n229 0.155672
R1292 VTAIL.n295 VTAIL.n229 0.155672
R1293 VTAIL.n296 VTAIL.n295 0.155672
R1294 VTAIL.n296 VTAIL.n225 0.155672
R1295 VTAIL.n303 VTAIL.n225 0.155672
R1296 VTAIL.n304 VTAIL.n303 0.155672
R1297 VTAIL.n304 VTAIL.n221 0.155672
R1298 VTAIL.n311 VTAIL.n221 0.155672
R1299 VTAIL.n312 VTAIL.n311 0.155672
R1300 VTAIL.n312 VTAIL.n217 0.155672
R1301 VTAIL.n319 VTAIL.n217 0.155672
R1302 VTAIL.n747 VTAIL.n645 0.155672
R1303 VTAIL.n740 VTAIL.n645 0.155672
R1304 VTAIL.n740 VTAIL.n739 0.155672
R1305 VTAIL.n739 VTAIL.n649 0.155672
R1306 VTAIL.n732 VTAIL.n649 0.155672
R1307 VTAIL.n732 VTAIL.n731 0.155672
R1308 VTAIL.n731 VTAIL.n653 0.155672
R1309 VTAIL.n724 VTAIL.n653 0.155672
R1310 VTAIL.n724 VTAIL.n723 0.155672
R1311 VTAIL.n723 VTAIL.n657 0.155672
R1312 VTAIL.n716 VTAIL.n657 0.155672
R1313 VTAIL.n716 VTAIL.n715 0.155672
R1314 VTAIL.n715 VTAIL.n661 0.155672
R1315 VTAIL.n708 VTAIL.n661 0.155672
R1316 VTAIL.n708 VTAIL.n707 0.155672
R1317 VTAIL.n707 VTAIL.n665 0.155672
R1318 VTAIL.n699 VTAIL.n665 0.155672
R1319 VTAIL.n699 VTAIL.n698 0.155672
R1320 VTAIL.n698 VTAIL.n669 0.155672
R1321 VTAIL.n691 VTAIL.n669 0.155672
R1322 VTAIL.n691 VTAIL.n690 0.155672
R1323 VTAIL.n690 VTAIL.n674 0.155672
R1324 VTAIL.n683 VTAIL.n674 0.155672
R1325 VTAIL.n683 VTAIL.n682 0.155672
R1326 VTAIL.n639 VTAIL.n537 0.155672
R1327 VTAIL.n632 VTAIL.n537 0.155672
R1328 VTAIL.n632 VTAIL.n631 0.155672
R1329 VTAIL.n631 VTAIL.n541 0.155672
R1330 VTAIL.n624 VTAIL.n541 0.155672
R1331 VTAIL.n624 VTAIL.n623 0.155672
R1332 VTAIL.n623 VTAIL.n545 0.155672
R1333 VTAIL.n616 VTAIL.n545 0.155672
R1334 VTAIL.n616 VTAIL.n615 0.155672
R1335 VTAIL.n615 VTAIL.n549 0.155672
R1336 VTAIL.n608 VTAIL.n549 0.155672
R1337 VTAIL.n608 VTAIL.n607 0.155672
R1338 VTAIL.n607 VTAIL.n553 0.155672
R1339 VTAIL.n600 VTAIL.n553 0.155672
R1340 VTAIL.n600 VTAIL.n599 0.155672
R1341 VTAIL.n599 VTAIL.n557 0.155672
R1342 VTAIL.n591 VTAIL.n557 0.155672
R1343 VTAIL.n591 VTAIL.n590 0.155672
R1344 VTAIL.n590 VTAIL.n561 0.155672
R1345 VTAIL.n583 VTAIL.n561 0.155672
R1346 VTAIL.n583 VTAIL.n582 0.155672
R1347 VTAIL.n582 VTAIL.n566 0.155672
R1348 VTAIL.n575 VTAIL.n566 0.155672
R1349 VTAIL.n575 VTAIL.n574 0.155672
R1350 VTAIL.n533 VTAIL.n431 0.155672
R1351 VTAIL.n526 VTAIL.n431 0.155672
R1352 VTAIL.n526 VTAIL.n525 0.155672
R1353 VTAIL.n525 VTAIL.n435 0.155672
R1354 VTAIL.n518 VTAIL.n435 0.155672
R1355 VTAIL.n518 VTAIL.n517 0.155672
R1356 VTAIL.n517 VTAIL.n439 0.155672
R1357 VTAIL.n510 VTAIL.n439 0.155672
R1358 VTAIL.n510 VTAIL.n509 0.155672
R1359 VTAIL.n509 VTAIL.n443 0.155672
R1360 VTAIL.n502 VTAIL.n443 0.155672
R1361 VTAIL.n502 VTAIL.n501 0.155672
R1362 VTAIL.n501 VTAIL.n447 0.155672
R1363 VTAIL.n494 VTAIL.n447 0.155672
R1364 VTAIL.n494 VTAIL.n493 0.155672
R1365 VTAIL.n493 VTAIL.n451 0.155672
R1366 VTAIL.n485 VTAIL.n451 0.155672
R1367 VTAIL.n485 VTAIL.n484 0.155672
R1368 VTAIL.n484 VTAIL.n455 0.155672
R1369 VTAIL.n477 VTAIL.n455 0.155672
R1370 VTAIL.n477 VTAIL.n476 0.155672
R1371 VTAIL.n476 VTAIL.n460 0.155672
R1372 VTAIL.n469 VTAIL.n460 0.155672
R1373 VTAIL.n469 VTAIL.n468 0.155672
R1374 VTAIL.n425 VTAIL.n323 0.155672
R1375 VTAIL.n418 VTAIL.n323 0.155672
R1376 VTAIL.n418 VTAIL.n417 0.155672
R1377 VTAIL.n417 VTAIL.n327 0.155672
R1378 VTAIL.n410 VTAIL.n327 0.155672
R1379 VTAIL.n410 VTAIL.n409 0.155672
R1380 VTAIL.n409 VTAIL.n331 0.155672
R1381 VTAIL.n402 VTAIL.n331 0.155672
R1382 VTAIL.n402 VTAIL.n401 0.155672
R1383 VTAIL.n401 VTAIL.n335 0.155672
R1384 VTAIL.n394 VTAIL.n335 0.155672
R1385 VTAIL.n394 VTAIL.n393 0.155672
R1386 VTAIL.n393 VTAIL.n339 0.155672
R1387 VTAIL.n386 VTAIL.n339 0.155672
R1388 VTAIL.n386 VTAIL.n385 0.155672
R1389 VTAIL.n385 VTAIL.n343 0.155672
R1390 VTAIL.n377 VTAIL.n343 0.155672
R1391 VTAIL.n377 VTAIL.n376 0.155672
R1392 VTAIL.n376 VTAIL.n347 0.155672
R1393 VTAIL.n369 VTAIL.n347 0.155672
R1394 VTAIL.n369 VTAIL.n368 0.155672
R1395 VTAIL.n368 VTAIL.n352 0.155672
R1396 VTAIL.n361 VTAIL.n352 0.155672
R1397 VTAIL.n361 VTAIL.n360 0.155672
R1398 VTAIL VTAIL.n1 0.0586897
R1399 VDD1 VDD1.n0 71.3882
R1400 VDD1.n3 VDD1.n2 71.2745
R1401 VDD1.n3 VDD1.n1 71.2745
R1402 VDD1.n5 VDD1.n4 70.1704
R1403 VDD1.n5 VDD1.n3 51.4923
R1404 VDD1.n4 VDD1.t6 1.67257
R1405 VDD1.n4 VDD1.t5 1.67257
R1406 VDD1.n0 VDD1.t1 1.67257
R1407 VDD1.n0 VDD1.t7 1.67257
R1408 VDD1.n2 VDD1.t0 1.67257
R1409 VDD1.n2 VDD1.t2 1.67257
R1410 VDD1.n1 VDD1.t3 1.67257
R1411 VDD1.n1 VDD1.t4 1.67257
R1412 VDD1 VDD1.n5 1.10179
R1413 B.n518 B.n517 585
R1414 B.n516 B.n147 585
R1415 B.n515 B.n514 585
R1416 B.n513 B.n148 585
R1417 B.n512 B.n511 585
R1418 B.n510 B.n149 585
R1419 B.n509 B.n508 585
R1420 B.n507 B.n150 585
R1421 B.n506 B.n505 585
R1422 B.n504 B.n151 585
R1423 B.n503 B.n502 585
R1424 B.n501 B.n152 585
R1425 B.n500 B.n499 585
R1426 B.n498 B.n153 585
R1427 B.n497 B.n496 585
R1428 B.n495 B.n154 585
R1429 B.n494 B.n493 585
R1430 B.n492 B.n155 585
R1431 B.n491 B.n490 585
R1432 B.n489 B.n156 585
R1433 B.n488 B.n487 585
R1434 B.n486 B.n157 585
R1435 B.n485 B.n484 585
R1436 B.n483 B.n158 585
R1437 B.n482 B.n481 585
R1438 B.n480 B.n159 585
R1439 B.n479 B.n478 585
R1440 B.n477 B.n160 585
R1441 B.n476 B.n475 585
R1442 B.n474 B.n161 585
R1443 B.n473 B.n472 585
R1444 B.n471 B.n162 585
R1445 B.n470 B.n469 585
R1446 B.n468 B.n163 585
R1447 B.n467 B.n466 585
R1448 B.n465 B.n164 585
R1449 B.n464 B.n463 585
R1450 B.n462 B.n165 585
R1451 B.n461 B.n460 585
R1452 B.n459 B.n166 585
R1453 B.n458 B.n457 585
R1454 B.n456 B.n167 585
R1455 B.n455 B.n454 585
R1456 B.n453 B.n168 585
R1457 B.n452 B.n451 585
R1458 B.n450 B.n169 585
R1459 B.n449 B.n448 585
R1460 B.n447 B.n170 585
R1461 B.n446 B.n445 585
R1462 B.n444 B.n171 585
R1463 B.n443 B.n442 585
R1464 B.n441 B.n172 585
R1465 B.n440 B.n439 585
R1466 B.n438 B.n173 585
R1467 B.n437 B.n436 585
R1468 B.n435 B.n174 585
R1469 B.n434 B.n433 585
R1470 B.n432 B.n175 585
R1471 B.n431 B.n430 585
R1472 B.n429 B.n176 585
R1473 B.n428 B.n427 585
R1474 B.n426 B.n177 585
R1475 B.n425 B.n424 585
R1476 B.n423 B.n178 585
R1477 B.n422 B.n421 585
R1478 B.n417 B.n179 585
R1479 B.n416 B.n415 585
R1480 B.n414 B.n180 585
R1481 B.n413 B.n412 585
R1482 B.n411 B.n181 585
R1483 B.n410 B.n409 585
R1484 B.n408 B.n182 585
R1485 B.n407 B.n406 585
R1486 B.n404 B.n183 585
R1487 B.n403 B.n402 585
R1488 B.n401 B.n186 585
R1489 B.n400 B.n399 585
R1490 B.n398 B.n187 585
R1491 B.n397 B.n396 585
R1492 B.n395 B.n188 585
R1493 B.n394 B.n393 585
R1494 B.n392 B.n189 585
R1495 B.n391 B.n390 585
R1496 B.n389 B.n190 585
R1497 B.n388 B.n387 585
R1498 B.n386 B.n191 585
R1499 B.n385 B.n384 585
R1500 B.n383 B.n192 585
R1501 B.n382 B.n381 585
R1502 B.n380 B.n193 585
R1503 B.n379 B.n378 585
R1504 B.n377 B.n194 585
R1505 B.n376 B.n375 585
R1506 B.n374 B.n195 585
R1507 B.n373 B.n372 585
R1508 B.n371 B.n196 585
R1509 B.n370 B.n369 585
R1510 B.n368 B.n197 585
R1511 B.n367 B.n366 585
R1512 B.n365 B.n198 585
R1513 B.n364 B.n363 585
R1514 B.n362 B.n199 585
R1515 B.n361 B.n360 585
R1516 B.n359 B.n200 585
R1517 B.n358 B.n357 585
R1518 B.n356 B.n201 585
R1519 B.n355 B.n354 585
R1520 B.n353 B.n202 585
R1521 B.n352 B.n351 585
R1522 B.n350 B.n203 585
R1523 B.n349 B.n348 585
R1524 B.n347 B.n204 585
R1525 B.n346 B.n345 585
R1526 B.n344 B.n205 585
R1527 B.n343 B.n342 585
R1528 B.n341 B.n206 585
R1529 B.n340 B.n339 585
R1530 B.n338 B.n207 585
R1531 B.n337 B.n336 585
R1532 B.n335 B.n208 585
R1533 B.n334 B.n333 585
R1534 B.n332 B.n209 585
R1535 B.n331 B.n330 585
R1536 B.n329 B.n210 585
R1537 B.n328 B.n327 585
R1538 B.n326 B.n211 585
R1539 B.n325 B.n324 585
R1540 B.n323 B.n212 585
R1541 B.n322 B.n321 585
R1542 B.n320 B.n213 585
R1543 B.n319 B.n318 585
R1544 B.n317 B.n214 585
R1545 B.n316 B.n315 585
R1546 B.n314 B.n215 585
R1547 B.n313 B.n312 585
R1548 B.n311 B.n216 585
R1549 B.n310 B.n309 585
R1550 B.n519 B.n146 585
R1551 B.n521 B.n520 585
R1552 B.n522 B.n145 585
R1553 B.n524 B.n523 585
R1554 B.n525 B.n144 585
R1555 B.n527 B.n526 585
R1556 B.n528 B.n143 585
R1557 B.n530 B.n529 585
R1558 B.n531 B.n142 585
R1559 B.n533 B.n532 585
R1560 B.n534 B.n141 585
R1561 B.n536 B.n535 585
R1562 B.n537 B.n140 585
R1563 B.n539 B.n538 585
R1564 B.n540 B.n139 585
R1565 B.n542 B.n541 585
R1566 B.n543 B.n138 585
R1567 B.n545 B.n544 585
R1568 B.n546 B.n137 585
R1569 B.n548 B.n547 585
R1570 B.n549 B.n136 585
R1571 B.n551 B.n550 585
R1572 B.n552 B.n135 585
R1573 B.n554 B.n553 585
R1574 B.n555 B.n134 585
R1575 B.n557 B.n556 585
R1576 B.n558 B.n133 585
R1577 B.n560 B.n559 585
R1578 B.n561 B.n132 585
R1579 B.n563 B.n562 585
R1580 B.n564 B.n131 585
R1581 B.n566 B.n565 585
R1582 B.n567 B.n130 585
R1583 B.n569 B.n568 585
R1584 B.n570 B.n129 585
R1585 B.n572 B.n571 585
R1586 B.n573 B.n128 585
R1587 B.n575 B.n574 585
R1588 B.n576 B.n127 585
R1589 B.n578 B.n577 585
R1590 B.n579 B.n126 585
R1591 B.n581 B.n580 585
R1592 B.n582 B.n125 585
R1593 B.n584 B.n583 585
R1594 B.n585 B.n124 585
R1595 B.n587 B.n586 585
R1596 B.n588 B.n123 585
R1597 B.n590 B.n589 585
R1598 B.n591 B.n122 585
R1599 B.n593 B.n592 585
R1600 B.n594 B.n121 585
R1601 B.n596 B.n595 585
R1602 B.n597 B.n120 585
R1603 B.n599 B.n598 585
R1604 B.n600 B.n119 585
R1605 B.n602 B.n601 585
R1606 B.n603 B.n118 585
R1607 B.n605 B.n604 585
R1608 B.n606 B.n117 585
R1609 B.n608 B.n607 585
R1610 B.n609 B.n116 585
R1611 B.n611 B.n610 585
R1612 B.n612 B.n115 585
R1613 B.n614 B.n613 585
R1614 B.n615 B.n114 585
R1615 B.n617 B.n616 585
R1616 B.n618 B.n113 585
R1617 B.n620 B.n619 585
R1618 B.n621 B.n112 585
R1619 B.n623 B.n622 585
R1620 B.n624 B.n111 585
R1621 B.n626 B.n625 585
R1622 B.n627 B.n110 585
R1623 B.n629 B.n628 585
R1624 B.n630 B.n109 585
R1625 B.n632 B.n631 585
R1626 B.n633 B.n108 585
R1627 B.n635 B.n634 585
R1628 B.n636 B.n107 585
R1629 B.n638 B.n637 585
R1630 B.n639 B.n106 585
R1631 B.n641 B.n640 585
R1632 B.n642 B.n105 585
R1633 B.n644 B.n643 585
R1634 B.n645 B.n104 585
R1635 B.n647 B.n646 585
R1636 B.n648 B.n103 585
R1637 B.n650 B.n649 585
R1638 B.n651 B.n102 585
R1639 B.n653 B.n652 585
R1640 B.n654 B.n101 585
R1641 B.n656 B.n655 585
R1642 B.n657 B.n100 585
R1643 B.n659 B.n658 585
R1644 B.n660 B.n99 585
R1645 B.n662 B.n661 585
R1646 B.n869 B.n868 585
R1647 B.n867 B.n26 585
R1648 B.n866 B.n865 585
R1649 B.n864 B.n27 585
R1650 B.n863 B.n862 585
R1651 B.n861 B.n28 585
R1652 B.n860 B.n859 585
R1653 B.n858 B.n29 585
R1654 B.n857 B.n856 585
R1655 B.n855 B.n30 585
R1656 B.n854 B.n853 585
R1657 B.n852 B.n31 585
R1658 B.n851 B.n850 585
R1659 B.n849 B.n32 585
R1660 B.n848 B.n847 585
R1661 B.n846 B.n33 585
R1662 B.n845 B.n844 585
R1663 B.n843 B.n34 585
R1664 B.n842 B.n841 585
R1665 B.n840 B.n35 585
R1666 B.n839 B.n838 585
R1667 B.n837 B.n36 585
R1668 B.n836 B.n835 585
R1669 B.n834 B.n37 585
R1670 B.n833 B.n832 585
R1671 B.n831 B.n38 585
R1672 B.n830 B.n829 585
R1673 B.n828 B.n39 585
R1674 B.n827 B.n826 585
R1675 B.n825 B.n40 585
R1676 B.n824 B.n823 585
R1677 B.n822 B.n41 585
R1678 B.n821 B.n820 585
R1679 B.n819 B.n42 585
R1680 B.n818 B.n817 585
R1681 B.n816 B.n43 585
R1682 B.n815 B.n814 585
R1683 B.n813 B.n44 585
R1684 B.n812 B.n811 585
R1685 B.n810 B.n45 585
R1686 B.n809 B.n808 585
R1687 B.n807 B.n46 585
R1688 B.n806 B.n805 585
R1689 B.n804 B.n47 585
R1690 B.n803 B.n802 585
R1691 B.n801 B.n48 585
R1692 B.n800 B.n799 585
R1693 B.n798 B.n49 585
R1694 B.n797 B.n796 585
R1695 B.n795 B.n50 585
R1696 B.n794 B.n793 585
R1697 B.n792 B.n51 585
R1698 B.n791 B.n790 585
R1699 B.n789 B.n52 585
R1700 B.n788 B.n787 585
R1701 B.n786 B.n53 585
R1702 B.n785 B.n784 585
R1703 B.n783 B.n54 585
R1704 B.n782 B.n781 585
R1705 B.n780 B.n55 585
R1706 B.n779 B.n778 585
R1707 B.n777 B.n56 585
R1708 B.n776 B.n775 585
R1709 B.n774 B.n57 585
R1710 B.n772 B.n771 585
R1711 B.n770 B.n60 585
R1712 B.n769 B.n768 585
R1713 B.n767 B.n61 585
R1714 B.n766 B.n765 585
R1715 B.n764 B.n62 585
R1716 B.n763 B.n762 585
R1717 B.n761 B.n63 585
R1718 B.n760 B.n759 585
R1719 B.n758 B.n757 585
R1720 B.n756 B.n67 585
R1721 B.n755 B.n754 585
R1722 B.n753 B.n68 585
R1723 B.n752 B.n751 585
R1724 B.n750 B.n69 585
R1725 B.n749 B.n748 585
R1726 B.n747 B.n70 585
R1727 B.n746 B.n745 585
R1728 B.n744 B.n71 585
R1729 B.n743 B.n742 585
R1730 B.n741 B.n72 585
R1731 B.n740 B.n739 585
R1732 B.n738 B.n73 585
R1733 B.n737 B.n736 585
R1734 B.n735 B.n74 585
R1735 B.n734 B.n733 585
R1736 B.n732 B.n75 585
R1737 B.n731 B.n730 585
R1738 B.n729 B.n76 585
R1739 B.n728 B.n727 585
R1740 B.n726 B.n77 585
R1741 B.n725 B.n724 585
R1742 B.n723 B.n78 585
R1743 B.n722 B.n721 585
R1744 B.n720 B.n79 585
R1745 B.n719 B.n718 585
R1746 B.n717 B.n80 585
R1747 B.n716 B.n715 585
R1748 B.n714 B.n81 585
R1749 B.n713 B.n712 585
R1750 B.n711 B.n82 585
R1751 B.n710 B.n709 585
R1752 B.n708 B.n83 585
R1753 B.n707 B.n706 585
R1754 B.n705 B.n84 585
R1755 B.n704 B.n703 585
R1756 B.n702 B.n85 585
R1757 B.n701 B.n700 585
R1758 B.n699 B.n86 585
R1759 B.n698 B.n697 585
R1760 B.n696 B.n87 585
R1761 B.n695 B.n694 585
R1762 B.n693 B.n88 585
R1763 B.n692 B.n691 585
R1764 B.n690 B.n89 585
R1765 B.n689 B.n688 585
R1766 B.n687 B.n90 585
R1767 B.n686 B.n685 585
R1768 B.n684 B.n91 585
R1769 B.n683 B.n682 585
R1770 B.n681 B.n92 585
R1771 B.n680 B.n679 585
R1772 B.n678 B.n93 585
R1773 B.n677 B.n676 585
R1774 B.n675 B.n94 585
R1775 B.n674 B.n673 585
R1776 B.n672 B.n95 585
R1777 B.n671 B.n670 585
R1778 B.n669 B.n96 585
R1779 B.n668 B.n667 585
R1780 B.n666 B.n97 585
R1781 B.n665 B.n664 585
R1782 B.n663 B.n98 585
R1783 B.n870 B.n25 585
R1784 B.n872 B.n871 585
R1785 B.n873 B.n24 585
R1786 B.n875 B.n874 585
R1787 B.n876 B.n23 585
R1788 B.n878 B.n877 585
R1789 B.n879 B.n22 585
R1790 B.n881 B.n880 585
R1791 B.n882 B.n21 585
R1792 B.n884 B.n883 585
R1793 B.n885 B.n20 585
R1794 B.n887 B.n886 585
R1795 B.n888 B.n19 585
R1796 B.n890 B.n889 585
R1797 B.n891 B.n18 585
R1798 B.n893 B.n892 585
R1799 B.n894 B.n17 585
R1800 B.n896 B.n895 585
R1801 B.n897 B.n16 585
R1802 B.n899 B.n898 585
R1803 B.n900 B.n15 585
R1804 B.n902 B.n901 585
R1805 B.n903 B.n14 585
R1806 B.n905 B.n904 585
R1807 B.n906 B.n13 585
R1808 B.n908 B.n907 585
R1809 B.n909 B.n12 585
R1810 B.n911 B.n910 585
R1811 B.n912 B.n11 585
R1812 B.n914 B.n913 585
R1813 B.n915 B.n10 585
R1814 B.n917 B.n916 585
R1815 B.n918 B.n9 585
R1816 B.n920 B.n919 585
R1817 B.n921 B.n8 585
R1818 B.n923 B.n922 585
R1819 B.n924 B.n7 585
R1820 B.n926 B.n925 585
R1821 B.n927 B.n6 585
R1822 B.n929 B.n928 585
R1823 B.n930 B.n5 585
R1824 B.n932 B.n931 585
R1825 B.n933 B.n4 585
R1826 B.n935 B.n934 585
R1827 B.n936 B.n3 585
R1828 B.n938 B.n937 585
R1829 B.n939 B.n0 585
R1830 B.n2 B.n1 585
R1831 B.n241 B.n240 585
R1832 B.n242 B.n239 585
R1833 B.n244 B.n243 585
R1834 B.n245 B.n238 585
R1835 B.n247 B.n246 585
R1836 B.n248 B.n237 585
R1837 B.n250 B.n249 585
R1838 B.n251 B.n236 585
R1839 B.n253 B.n252 585
R1840 B.n254 B.n235 585
R1841 B.n256 B.n255 585
R1842 B.n257 B.n234 585
R1843 B.n259 B.n258 585
R1844 B.n260 B.n233 585
R1845 B.n262 B.n261 585
R1846 B.n263 B.n232 585
R1847 B.n265 B.n264 585
R1848 B.n266 B.n231 585
R1849 B.n268 B.n267 585
R1850 B.n269 B.n230 585
R1851 B.n271 B.n270 585
R1852 B.n272 B.n229 585
R1853 B.n274 B.n273 585
R1854 B.n275 B.n228 585
R1855 B.n277 B.n276 585
R1856 B.n278 B.n227 585
R1857 B.n280 B.n279 585
R1858 B.n281 B.n226 585
R1859 B.n283 B.n282 585
R1860 B.n284 B.n225 585
R1861 B.n286 B.n285 585
R1862 B.n287 B.n224 585
R1863 B.n289 B.n288 585
R1864 B.n290 B.n223 585
R1865 B.n292 B.n291 585
R1866 B.n293 B.n222 585
R1867 B.n295 B.n294 585
R1868 B.n296 B.n221 585
R1869 B.n298 B.n297 585
R1870 B.n299 B.n220 585
R1871 B.n301 B.n300 585
R1872 B.n302 B.n219 585
R1873 B.n304 B.n303 585
R1874 B.n305 B.n218 585
R1875 B.n307 B.n306 585
R1876 B.n308 B.n217 585
R1877 B.n418 B.t7 561.653
R1878 B.n64 B.t11 561.653
R1879 B.n184 B.t1 561.653
R1880 B.n58 B.t5 561.653
R1881 B.n419 B.t8 509.483
R1882 B.n65 B.t10 509.483
R1883 B.n185 B.t2 509.483
R1884 B.n59 B.t4 509.483
R1885 B.n310 B.n217 492.5
R1886 B.n519 B.n518 492.5
R1887 B.n663 B.n662 492.5
R1888 B.n868 B.n25 492.5
R1889 B.n184 B.t0 406.173
R1890 B.n418 B.t6 406.173
R1891 B.n64 B.t9 406.173
R1892 B.n58 B.t3 406.173
R1893 B.n941 B.n940 256.663
R1894 B.n940 B.n939 235.042
R1895 B.n940 B.n2 235.042
R1896 B.n311 B.n310 163.367
R1897 B.n312 B.n311 163.367
R1898 B.n312 B.n215 163.367
R1899 B.n316 B.n215 163.367
R1900 B.n317 B.n316 163.367
R1901 B.n318 B.n317 163.367
R1902 B.n318 B.n213 163.367
R1903 B.n322 B.n213 163.367
R1904 B.n323 B.n322 163.367
R1905 B.n324 B.n323 163.367
R1906 B.n324 B.n211 163.367
R1907 B.n328 B.n211 163.367
R1908 B.n329 B.n328 163.367
R1909 B.n330 B.n329 163.367
R1910 B.n330 B.n209 163.367
R1911 B.n334 B.n209 163.367
R1912 B.n335 B.n334 163.367
R1913 B.n336 B.n335 163.367
R1914 B.n336 B.n207 163.367
R1915 B.n340 B.n207 163.367
R1916 B.n341 B.n340 163.367
R1917 B.n342 B.n341 163.367
R1918 B.n342 B.n205 163.367
R1919 B.n346 B.n205 163.367
R1920 B.n347 B.n346 163.367
R1921 B.n348 B.n347 163.367
R1922 B.n348 B.n203 163.367
R1923 B.n352 B.n203 163.367
R1924 B.n353 B.n352 163.367
R1925 B.n354 B.n353 163.367
R1926 B.n354 B.n201 163.367
R1927 B.n358 B.n201 163.367
R1928 B.n359 B.n358 163.367
R1929 B.n360 B.n359 163.367
R1930 B.n360 B.n199 163.367
R1931 B.n364 B.n199 163.367
R1932 B.n365 B.n364 163.367
R1933 B.n366 B.n365 163.367
R1934 B.n366 B.n197 163.367
R1935 B.n370 B.n197 163.367
R1936 B.n371 B.n370 163.367
R1937 B.n372 B.n371 163.367
R1938 B.n372 B.n195 163.367
R1939 B.n376 B.n195 163.367
R1940 B.n377 B.n376 163.367
R1941 B.n378 B.n377 163.367
R1942 B.n378 B.n193 163.367
R1943 B.n382 B.n193 163.367
R1944 B.n383 B.n382 163.367
R1945 B.n384 B.n383 163.367
R1946 B.n384 B.n191 163.367
R1947 B.n388 B.n191 163.367
R1948 B.n389 B.n388 163.367
R1949 B.n390 B.n389 163.367
R1950 B.n390 B.n189 163.367
R1951 B.n394 B.n189 163.367
R1952 B.n395 B.n394 163.367
R1953 B.n396 B.n395 163.367
R1954 B.n396 B.n187 163.367
R1955 B.n400 B.n187 163.367
R1956 B.n401 B.n400 163.367
R1957 B.n402 B.n401 163.367
R1958 B.n402 B.n183 163.367
R1959 B.n407 B.n183 163.367
R1960 B.n408 B.n407 163.367
R1961 B.n409 B.n408 163.367
R1962 B.n409 B.n181 163.367
R1963 B.n413 B.n181 163.367
R1964 B.n414 B.n413 163.367
R1965 B.n415 B.n414 163.367
R1966 B.n415 B.n179 163.367
R1967 B.n422 B.n179 163.367
R1968 B.n423 B.n422 163.367
R1969 B.n424 B.n423 163.367
R1970 B.n424 B.n177 163.367
R1971 B.n428 B.n177 163.367
R1972 B.n429 B.n428 163.367
R1973 B.n430 B.n429 163.367
R1974 B.n430 B.n175 163.367
R1975 B.n434 B.n175 163.367
R1976 B.n435 B.n434 163.367
R1977 B.n436 B.n435 163.367
R1978 B.n436 B.n173 163.367
R1979 B.n440 B.n173 163.367
R1980 B.n441 B.n440 163.367
R1981 B.n442 B.n441 163.367
R1982 B.n442 B.n171 163.367
R1983 B.n446 B.n171 163.367
R1984 B.n447 B.n446 163.367
R1985 B.n448 B.n447 163.367
R1986 B.n448 B.n169 163.367
R1987 B.n452 B.n169 163.367
R1988 B.n453 B.n452 163.367
R1989 B.n454 B.n453 163.367
R1990 B.n454 B.n167 163.367
R1991 B.n458 B.n167 163.367
R1992 B.n459 B.n458 163.367
R1993 B.n460 B.n459 163.367
R1994 B.n460 B.n165 163.367
R1995 B.n464 B.n165 163.367
R1996 B.n465 B.n464 163.367
R1997 B.n466 B.n465 163.367
R1998 B.n466 B.n163 163.367
R1999 B.n470 B.n163 163.367
R2000 B.n471 B.n470 163.367
R2001 B.n472 B.n471 163.367
R2002 B.n472 B.n161 163.367
R2003 B.n476 B.n161 163.367
R2004 B.n477 B.n476 163.367
R2005 B.n478 B.n477 163.367
R2006 B.n478 B.n159 163.367
R2007 B.n482 B.n159 163.367
R2008 B.n483 B.n482 163.367
R2009 B.n484 B.n483 163.367
R2010 B.n484 B.n157 163.367
R2011 B.n488 B.n157 163.367
R2012 B.n489 B.n488 163.367
R2013 B.n490 B.n489 163.367
R2014 B.n490 B.n155 163.367
R2015 B.n494 B.n155 163.367
R2016 B.n495 B.n494 163.367
R2017 B.n496 B.n495 163.367
R2018 B.n496 B.n153 163.367
R2019 B.n500 B.n153 163.367
R2020 B.n501 B.n500 163.367
R2021 B.n502 B.n501 163.367
R2022 B.n502 B.n151 163.367
R2023 B.n506 B.n151 163.367
R2024 B.n507 B.n506 163.367
R2025 B.n508 B.n507 163.367
R2026 B.n508 B.n149 163.367
R2027 B.n512 B.n149 163.367
R2028 B.n513 B.n512 163.367
R2029 B.n514 B.n513 163.367
R2030 B.n514 B.n147 163.367
R2031 B.n518 B.n147 163.367
R2032 B.n662 B.n99 163.367
R2033 B.n658 B.n99 163.367
R2034 B.n658 B.n657 163.367
R2035 B.n657 B.n656 163.367
R2036 B.n656 B.n101 163.367
R2037 B.n652 B.n101 163.367
R2038 B.n652 B.n651 163.367
R2039 B.n651 B.n650 163.367
R2040 B.n650 B.n103 163.367
R2041 B.n646 B.n103 163.367
R2042 B.n646 B.n645 163.367
R2043 B.n645 B.n644 163.367
R2044 B.n644 B.n105 163.367
R2045 B.n640 B.n105 163.367
R2046 B.n640 B.n639 163.367
R2047 B.n639 B.n638 163.367
R2048 B.n638 B.n107 163.367
R2049 B.n634 B.n107 163.367
R2050 B.n634 B.n633 163.367
R2051 B.n633 B.n632 163.367
R2052 B.n632 B.n109 163.367
R2053 B.n628 B.n109 163.367
R2054 B.n628 B.n627 163.367
R2055 B.n627 B.n626 163.367
R2056 B.n626 B.n111 163.367
R2057 B.n622 B.n111 163.367
R2058 B.n622 B.n621 163.367
R2059 B.n621 B.n620 163.367
R2060 B.n620 B.n113 163.367
R2061 B.n616 B.n113 163.367
R2062 B.n616 B.n615 163.367
R2063 B.n615 B.n614 163.367
R2064 B.n614 B.n115 163.367
R2065 B.n610 B.n115 163.367
R2066 B.n610 B.n609 163.367
R2067 B.n609 B.n608 163.367
R2068 B.n608 B.n117 163.367
R2069 B.n604 B.n117 163.367
R2070 B.n604 B.n603 163.367
R2071 B.n603 B.n602 163.367
R2072 B.n602 B.n119 163.367
R2073 B.n598 B.n119 163.367
R2074 B.n598 B.n597 163.367
R2075 B.n597 B.n596 163.367
R2076 B.n596 B.n121 163.367
R2077 B.n592 B.n121 163.367
R2078 B.n592 B.n591 163.367
R2079 B.n591 B.n590 163.367
R2080 B.n590 B.n123 163.367
R2081 B.n586 B.n123 163.367
R2082 B.n586 B.n585 163.367
R2083 B.n585 B.n584 163.367
R2084 B.n584 B.n125 163.367
R2085 B.n580 B.n125 163.367
R2086 B.n580 B.n579 163.367
R2087 B.n579 B.n578 163.367
R2088 B.n578 B.n127 163.367
R2089 B.n574 B.n127 163.367
R2090 B.n574 B.n573 163.367
R2091 B.n573 B.n572 163.367
R2092 B.n572 B.n129 163.367
R2093 B.n568 B.n129 163.367
R2094 B.n568 B.n567 163.367
R2095 B.n567 B.n566 163.367
R2096 B.n566 B.n131 163.367
R2097 B.n562 B.n131 163.367
R2098 B.n562 B.n561 163.367
R2099 B.n561 B.n560 163.367
R2100 B.n560 B.n133 163.367
R2101 B.n556 B.n133 163.367
R2102 B.n556 B.n555 163.367
R2103 B.n555 B.n554 163.367
R2104 B.n554 B.n135 163.367
R2105 B.n550 B.n135 163.367
R2106 B.n550 B.n549 163.367
R2107 B.n549 B.n548 163.367
R2108 B.n548 B.n137 163.367
R2109 B.n544 B.n137 163.367
R2110 B.n544 B.n543 163.367
R2111 B.n543 B.n542 163.367
R2112 B.n542 B.n139 163.367
R2113 B.n538 B.n139 163.367
R2114 B.n538 B.n537 163.367
R2115 B.n537 B.n536 163.367
R2116 B.n536 B.n141 163.367
R2117 B.n532 B.n141 163.367
R2118 B.n532 B.n531 163.367
R2119 B.n531 B.n530 163.367
R2120 B.n530 B.n143 163.367
R2121 B.n526 B.n143 163.367
R2122 B.n526 B.n525 163.367
R2123 B.n525 B.n524 163.367
R2124 B.n524 B.n145 163.367
R2125 B.n520 B.n145 163.367
R2126 B.n520 B.n519 163.367
R2127 B.n868 B.n867 163.367
R2128 B.n867 B.n866 163.367
R2129 B.n866 B.n27 163.367
R2130 B.n862 B.n27 163.367
R2131 B.n862 B.n861 163.367
R2132 B.n861 B.n860 163.367
R2133 B.n860 B.n29 163.367
R2134 B.n856 B.n29 163.367
R2135 B.n856 B.n855 163.367
R2136 B.n855 B.n854 163.367
R2137 B.n854 B.n31 163.367
R2138 B.n850 B.n31 163.367
R2139 B.n850 B.n849 163.367
R2140 B.n849 B.n848 163.367
R2141 B.n848 B.n33 163.367
R2142 B.n844 B.n33 163.367
R2143 B.n844 B.n843 163.367
R2144 B.n843 B.n842 163.367
R2145 B.n842 B.n35 163.367
R2146 B.n838 B.n35 163.367
R2147 B.n838 B.n837 163.367
R2148 B.n837 B.n836 163.367
R2149 B.n836 B.n37 163.367
R2150 B.n832 B.n37 163.367
R2151 B.n832 B.n831 163.367
R2152 B.n831 B.n830 163.367
R2153 B.n830 B.n39 163.367
R2154 B.n826 B.n39 163.367
R2155 B.n826 B.n825 163.367
R2156 B.n825 B.n824 163.367
R2157 B.n824 B.n41 163.367
R2158 B.n820 B.n41 163.367
R2159 B.n820 B.n819 163.367
R2160 B.n819 B.n818 163.367
R2161 B.n818 B.n43 163.367
R2162 B.n814 B.n43 163.367
R2163 B.n814 B.n813 163.367
R2164 B.n813 B.n812 163.367
R2165 B.n812 B.n45 163.367
R2166 B.n808 B.n45 163.367
R2167 B.n808 B.n807 163.367
R2168 B.n807 B.n806 163.367
R2169 B.n806 B.n47 163.367
R2170 B.n802 B.n47 163.367
R2171 B.n802 B.n801 163.367
R2172 B.n801 B.n800 163.367
R2173 B.n800 B.n49 163.367
R2174 B.n796 B.n49 163.367
R2175 B.n796 B.n795 163.367
R2176 B.n795 B.n794 163.367
R2177 B.n794 B.n51 163.367
R2178 B.n790 B.n51 163.367
R2179 B.n790 B.n789 163.367
R2180 B.n789 B.n788 163.367
R2181 B.n788 B.n53 163.367
R2182 B.n784 B.n53 163.367
R2183 B.n784 B.n783 163.367
R2184 B.n783 B.n782 163.367
R2185 B.n782 B.n55 163.367
R2186 B.n778 B.n55 163.367
R2187 B.n778 B.n777 163.367
R2188 B.n777 B.n776 163.367
R2189 B.n776 B.n57 163.367
R2190 B.n771 B.n57 163.367
R2191 B.n771 B.n770 163.367
R2192 B.n770 B.n769 163.367
R2193 B.n769 B.n61 163.367
R2194 B.n765 B.n61 163.367
R2195 B.n765 B.n764 163.367
R2196 B.n764 B.n763 163.367
R2197 B.n763 B.n63 163.367
R2198 B.n759 B.n63 163.367
R2199 B.n759 B.n758 163.367
R2200 B.n758 B.n67 163.367
R2201 B.n754 B.n67 163.367
R2202 B.n754 B.n753 163.367
R2203 B.n753 B.n752 163.367
R2204 B.n752 B.n69 163.367
R2205 B.n748 B.n69 163.367
R2206 B.n748 B.n747 163.367
R2207 B.n747 B.n746 163.367
R2208 B.n746 B.n71 163.367
R2209 B.n742 B.n71 163.367
R2210 B.n742 B.n741 163.367
R2211 B.n741 B.n740 163.367
R2212 B.n740 B.n73 163.367
R2213 B.n736 B.n73 163.367
R2214 B.n736 B.n735 163.367
R2215 B.n735 B.n734 163.367
R2216 B.n734 B.n75 163.367
R2217 B.n730 B.n75 163.367
R2218 B.n730 B.n729 163.367
R2219 B.n729 B.n728 163.367
R2220 B.n728 B.n77 163.367
R2221 B.n724 B.n77 163.367
R2222 B.n724 B.n723 163.367
R2223 B.n723 B.n722 163.367
R2224 B.n722 B.n79 163.367
R2225 B.n718 B.n79 163.367
R2226 B.n718 B.n717 163.367
R2227 B.n717 B.n716 163.367
R2228 B.n716 B.n81 163.367
R2229 B.n712 B.n81 163.367
R2230 B.n712 B.n711 163.367
R2231 B.n711 B.n710 163.367
R2232 B.n710 B.n83 163.367
R2233 B.n706 B.n83 163.367
R2234 B.n706 B.n705 163.367
R2235 B.n705 B.n704 163.367
R2236 B.n704 B.n85 163.367
R2237 B.n700 B.n85 163.367
R2238 B.n700 B.n699 163.367
R2239 B.n699 B.n698 163.367
R2240 B.n698 B.n87 163.367
R2241 B.n694 B.n87 163.367
R2242 B.n694 B.n693 163.367
R2243 B.n693 B.n692 163.367
R2244 B.n692 B.n89 163.367
R2245 B.n688 B.n89 163.367
R2246 B.n688 B.n687 163.367
R2247 B.n687 B.n686 163.367
R2248 B.n686 B.n91 163.367
R2249 B.n682 B.n91 163.367
R2250 B.n682 B.n681 163.367
R2251 B.n681 B.n680 163.367
R2252 B.n680 B.n93 163.367
R2253 B.n676 B.n93 163.367
R2254 B.n676 B.n675 163.367
R2255 B.n675 B.n674 163.367
R2256 B.n674 B.n95 163.367
R2257 B.n670 B.n95 163.367
R2258 B.n670 B.n669 163.367
R2259 B.n669 B.n668 163.367
R2260 B.n668 B.n97 163.367
R2261 B.n664 B.n97 163.367
R2262 B.n664 B.n663 163.367
R2263 B.n872 B.n25 163.367
R2264 B.n873 B.n872 163.367
R2265 B.n874 B.n873 163.367
R2266 B.n874 B.n23 163.367
R2267 B.n878 B.n23 163.367
R2268 B.n879 B.n878 163.367
R2269 B.n880 B.n879 163.367
R2270 B.n880 B.n21 163.367
R2271 B.n884 B.n21 163.367
R2272 B.n885 B.n884 163.367
R2273 B.n886 B.n885 163.367
R2274 B.n886 B.n19 163.367
R2275 B.n890 B.n19 163.367
R2276 B.n891 B.n890 163.367
R2277 B.n892 B.n891 163.367
R2278 B.n892 B.n17 163.367
R2279 B.n896 B.n17 163.367
R2280 B.n897 B.n896 163.367
R2281 B.n898 B.n897 163.367
R2282 B.n898 B.n15 163.367
R2283 B.n902 B.n15 163.367
R2284 B.n903 B.n902 163.367
R2285 B.n904 B.n903 163.367
R2286 B.n904 B.n13 163.367
R2287 B.n908 B.n13 163.367
R2288 B.n909 B.n908 163.367
R2289 B.n910 B.n909 163.367
R2290 B.n910 B.n11 163.367
R2291 B.n914 B.n11 163.367
R2292 B.n915 B.n914 163.367
R2293 B.n916 B.n915 163.367
R2294 B.n916 B.n9 163.367
R2295 B.n920 B.n9 163.367
R2296 B.n921 B.n920 163.367
R2297 B.n922 B.n921 163.367
R2298 B.n922 B.n7 163.367
R2299 B.n926 B.n7 163.367
R2300 B.n927 B.n926 163.367
R2301 B.n928 B.n927 163.367
R2302 B.n928 B.n5 163.367
R2303 B.n932 B.n5 163.367
R2304 B.n933 B.n932 163.367
R2305 B.n934 B.n933 163.367
R2306 B.n934 B.n3 163.367
R2307 B.n938 B.n3 163.367
R2308 B.n939 B.n938 163.367
R2309 B.n240 B.n2 163.367
R2310 B.n240 B.n239 163.367
R2311 B.n244 B.n239 163.367
R2312 B.n245 B.n244 163.367
R2313 B.n246 B.n245 163.367
R2314 B.n246 B.n237 163.367
R2315 B.n250 B.n237 163.367
R2316 B.n251 B.n250 163.367
R2317 B.n252 B.n251 163.367
R2318 B.n252 B.n235 163.367
R2319 B.n256 B.n235 163.367
R2320 B.n257 B.n256 163.367
R2321 B.n258 B.n257 163.367
R2322 B.n258 B.n233 163.367
R2323 B.n262 B.n233 163.367
R2324 B.n263 B.n262 163.367
R2325 B.n264 B.n263 163.367
R2326 B.n264 B.n231 163.367
R2327 B.n268 B.n231 163.367
R2328 B.n269 B.n268 163.367
R2329 B.n270 B.n269 163.367
R2330 B.n270 B.n229 163.367
R2331 B.n274 B.n229 163.367
R2332 B.n275 B.n274 163.367
R2333 B.n276 B.n275 163.367
R2334 B.n276 B.n227 163.367
R2335 B.n280 B.n227 163.367
R2336 B.n281 B.n280 163.367
R2337 B.n282 B.n281 163.367
R2338 B.n282 B.n225 163.367
R2339 B.n286 B.n225 163.367
R2340 B.n287 B.n286 163.367
R2341 B.n288 B.n287 163.367
R2342 B.n288 B.n223 163.367
R2343 B.n292 B.n223 163.367
R2344 B.n293 B.n292 163.367
R2345 B.n294 B.n293 163.367
R2346 B.n294 B.n221 163.367
R2347 B.n298 B.n221 163.367
R2348 B.n299 B.n298 163.367
R2349 B.n300 B.n299 163.367
R2350 B.n300 B.n219 163.367
R2351 B.n304 B.n219 163.367
R2352 B.n305 B.n304 163.367
R2353 B.n306 B.n305 163.367
R2354 B.n306 B.n217 163.367
R2355 B.n405 B.n185 59.5399
R2356 B.n420 B.n419 59.5399
R2357 B.n66 B.n65 59.5399
R2358 B.n773 B.n59 59.5399
R2359 B.n185 B.n184 52.1702
R2360 B.n419 B.n418 52.1702
R2361 B.n65 B.n64 52.1702
R2362 B.n59 B.n58 52.1702
R2363 B.n870 B.n869 32.0005
R2364 B.n661 B.n98 32.0005
R2365 B.n517 B.n146 32.0005
R2366 B.n309 B.n308 32.0005
R2367 B B.n941 18.0485
R2368 B.n871 B.n870 10.6151
R2369 B.n871 B.n24 10.6151
R2370 B.n875 B.n24 10.6151
R2371 B.n876 B.n875 10.6151
R2372 B.n877 B.n876 10.6151
R2373 B.n877 B.n22 10.6151
R2374 B.n881 B.n22 10.6151
R2375 B.n882 B.n881 10.6151
R2376 B.n883 B.n882 10.6151
R2377 B.n883 B.n20 10.6151
R2378 B.n887 B.n20 10.6151
R2379 B.n888 B.n887 10.6151
R2380 B.n889 B.n888 10.6151
R2381 B.n889 B.n18 10.6151
R2382 B.n893 B.n18 10.6151
R2383 B.n894 B.n893 10.6151
R2384 B.n895 B.n894 10.6151
R2385 B.n895 B.n16 10.6151
R2386 B.n899 B.n16 10.6151
R2387 B.n900 B.n899 10.6151
R2388 B.n901 B.n900 10.6151
R2389 B.n901 B.n14 10.6151
R2390 B.n905 B.n14 10.6151
R2391 B.n906 B.n905 10.6151
R2392 B.n907 B.n906 10.6151
R2393 B.n907 B.n12 10.6151
R2394 B.n911 B.n12 10.6151
R2395 B.n912 B.n911 10.6151
R2396 B.n913 B.n912 10.6151
R2397 B.n913 B.n10 10.6151
R2398 B.n917 B.n10 10.6151
R2399 B.n918 B.n917 10.6151
R2400 B.n919 B.n918 10.6151
R2401 B.n919 B.n8 10.6151
R2402 B.n923 B.n8 10.6151
R2403 B.n924 B.n923 10.6151
R2404 B.n925 B.n924 10.6151
R2405 B.n925 B.n6 10.6151
R2406 B.n929 B.n6 10.6151
R2407 B.n930 B.n929 10.6151
R2408 B.n931 B.n930 10.6151
R2409 B.n931 B.n4 10.6151
R2410 B.n935 B.n4 10.6151
R2411 B.n936 B.n935 10.6151
R2412 B.n937 B.n936 10.6151
R2413 B.n937 B.n0 10.6151
R2414 B.n869 B.n26 10.6151
R2415 B.n865 B.n26 10.6151
R2416 B.n865 B.n864 10.6151
R2417 B.n864 B.n863 10.6151
R2418 B.n863 B.n28 10.6151
R2419 B.n859 B.n28 10.6151
R2420 B.n859 B.n858 10.6151
R2421 B.n858 B.n857 10.6151
R2422 B.n857 B.n30 10.6151
R2423 B.n853 B.n30 10.6151
R2424 B.n853 B.n852 10.6151
R2425 B.n852 B.n851 10.6151
R2426 B.n851 B.n32 10.6151
R2427 B.n847 B.n32 10.6151
R2428 B.n847 B.n846 10.6151
R2429 B.n846 B.n845 10.6151
R2430 B.n845 B.n34 10.6151
R2431 B.n841 B.n34 10.6151
R2432 B.n841 B.n840 10.6151
R2433 B.n840 B.n839 10.6151
R2434 B.n839 B.n36 10.6151
R2435 B.n835 B.n36 10.6151
R2436 B.n835 B.n834 10.6151
R2437 B.n834 B.n833 10.6151
R2438 B.n833 B.n38 10.6151
R2439 B.n829 B.n38 10.6151
R2440 B.n829 B.n828 10.6151
R2441 B.n828 B.n827 10.6151
R2442 B.n827 B.n40 10.6151
R2443 B.n823 B.n40 10.6151
R2444 B.n823 B.n822 10.6151
R2445 B.n822 B.n821 10.6151
R2446 B.n821 B.n42 10.6151
R2447 B.n817 B.n42 10.6151
R2448 B.n817 B.n816 10.6151
R2449 B.n816 B.n815 10.6151
R2450 B.n815 B.n44 10.6151
R2451 B.n811 B.n44 10.6151
R2452 B.n811 B.n810 10.6151
R2453 B.n810 B.n809 10.6151
R2454 B.n809 B.n46 10.6151
R2455 B.n805 B.n46 10.6151
R2456 B.n805 B.n804 10.6151
R2457 B.n804 B.n803 10.6151
R2458 B.n803 B.n48 10.6151
R2459 B.n799 B.n48 10.6151
R2460 B.n799 B.n798 10.6151
R2461 B.n798 B.n797 10.6151
R2462 B.n797 B.n50 10.6151
R2463 B.n793 B.n50 10.6151
R2464 B.n793 B.n792 10.6151
R2465 B.n792 B.n791 10.6151
R2466 B.n791 B.n52 10.6151
R2467 B.n787 B.n52 10.6151
R2468 B.n787 B.n786 10.6151
R2469 B.n786 B.n785 10.6151
R2470 B.n785 B.n54 10.6151
R2471 B.n781 B.n54 10.6151
R2472 B.n781 B.n780 10.6151
R2473 B.n780 B.n779 10.6151
R2474 B.n779 B.n56 10.6151
R2475 B.n775 B.n56 10.6151
R2476 B.n775 B.n774 10.6151
R2477 B.n772 B.n60 10.6151
R2478 B.n768 B.n60 10.6151
R2479 B.n768 B.n767 10.6151
R2480 B.n767 B.n766 10.6151
R2481 B.n766 B.n62 10.6151
R2482 B.n762 B.n62 10.6151
R2483 B.n762 B.n761 10.6151
R2484 B.n761 B.n760 10.6151
R2485 B.n757 B.n756 10.6151
R2486 B.n756 B.n755 10.6151
R2487 B.n755 B.n68 10.6151
R2488 B.n751 B.n68 10.6151
R2489 B.n751 B.n750 10.6151
R2490 B.n750 B.n749 10.6151
R2491 B.n749 B.n70 10.6151
R2492 B.n745 B.n70 10.6151
R2493 B.n745 B.n744 10.6151
R2494 B.n744 B.n743 10.6151
R2495 B.n743 B.n72 10.6151
R2496 B.n739 B.n72 10.6151
R2497 B.n739 B.n738 10.6151
R2498 B.n738 B.n737 10.6151
R2499 B.n737 B.n74 10.6151
R2500 B.n733 B.n74 10.6151
R2501 B.n733 B.n732 10.6151
R2502 B.n732 B.n731 10.6151
R2503 B.n731 B.n76 10.6151
R2504 B.n727 B.n76 10.6151
R2505 B.n727 B.n726 10.6151
R2506 B.n726 B.n725 10.6151
R2507 B.n725 B.n78 10.6151
R2508 B.n721 B.n78 10.6151
R2509 B.n721 B.n720 10.6151
R2510 B.n720 B.n719 10.6151
R2511 B.n719 B.n80 10.6151
R2512 B.n715 B.n80 10.6151
R2513 B.n715 B.n714 10.6151
R2514 B.n714 B.n713 10.6151
R2515 B.n713 B.n82 10.6151
R2516 B.n709 B.n82 10.6151
R2517 B.n709 B.n708 10.6151
R2518 B.n708 B.n707 10.6151
R2519 B.n707 B.n84 10.6151
R2520 B.n703 B.n84 10.6151
R2521 B.n703 B.n702 10.6151
R2522 B.n702 B.n701 10.6151
R2523 B.n701 B.n86 10.6151
R2524 B.n697 B.n86 10.6151
R2525 B.n697 B.n696 10.6151
R2526 B.n696 B.n695 10.6151
R2527 B.n695 B.n88 10.6151
R2528 B.n691 B.n88 10.6151
R2529 B.n691 B.n690 10.6151
R2530 B.n690 B.n689 10.6151
R2531 B.n689 B.n90 10.6151
R2532 B.n685 B.n90 10.6151
R2533 B.n685 B.n684 10.6151
R2534 B.n684 B.n683 10.6151
R2535 B.n683 B.n92 10.6151
R2536 B.n679 B.n92 10.6151
R2537 B.n679 B.n678 10.6151
R2538 B.n678 B.n677 10.6151
R2539 B.n677 B.n94 10.6151
R2540 B.n673 B.n94 10.6151
R2541 B.n673 B.n672 10.6151
R2542 B.n672 B.n671 10.6151
R2543 B.n671 B.n96 10.6151
R2544 B.n667 B.n96 10.6151
R2545 B.n667 B.n666 10.6151
R2546 B.n666 B.n665 10.6151
R2547 B.n665 B.n98 10.6151
R2548 B.n661 B.n660 10.6151
R2549 B.n660 B.n659 10.6151
R2550 B.n659 B.n100 10.6151
R2551 B.n655 B.n100 10.6151
R2552 B.n655 B.n654 10.6151
R2553 B.n654 B.n653 10.6151
R2554 B.n653 B.n102 10.6151
R2555 B.n649 B.n102 10.6151
R2556 B.n649 B.n648 10.6151
R2557 B.n648 B.n647 10.6151
R2558 B.n647 B.n104 10.6151
R2559 B.n643 B.n104 10.6151
R2560 B.n643 B.n642 10.6151
R2561 B.n642 B.n641 10.6151
R2562 B.n641 B.n106 10.6151
R2563 B.n637 B.n106 10.6151
R2564 B.n637 B.n636 10.6151
R2565 B.n636 B.n635 10.6151
R2566 B.n635 B.n108 10.6151
R2567 B.n631 B.n108 10.6151
R2568 B.n631 B.n630 10.6151
R2569 B.n630 B.n629 10.6151
R2570 B.n629 B.n110 10.6151
R2571 B.n625 B.n110 10.6151
R2572 B.n625 B.n624 10.6151
R2573 B.n624 B.n623 10.6151
R2574 B.n623 B.n112 10.6151
R2575 B.n619 B.n112 10.6151
R2576 B.n619 B.n618 10.6151
R2577 B.n618 B.n617 10.6151
R2578 B.n617 B.n114 10.6151
R2579 B.n613 B.n114 10.6151
R2580 B.n613 B.n612 10.6151
R2581 B.n612 B.n611 10.6151
R2582 B.n611 B.n116 10.6151
R2583 B.n607 B.n116 10.6151
R2584 B.n607 B.n606 10.6151
R2585 B.n606 B.n605 10.6151
R2586 B.n605 B.n118 10.6151
R2587 B.n601 B.n118 10.6151
R2588 B.n601 B.n600 10.6151
R2589 B.n600 B.n599 10.6151
R2590 B.n599 B.n120 10.6151
R2591 B.n595 B.n120 10.6151
R2592 B.n595 B.n594 10.6151
R2593 B.n594 B.n593 10.6151
R2594 B.n593 B.n122 10.6151
R2595 B.n589 B.n122 10.6151
R2596 B.n589 B.n588 10.6151
R2597 B.n588 B.n587 10.6151
R2598 B.n587 B.n124 10.6151
R2599 B.n583 B.n124 10.6151
R2600 B.n583 B.n582 10.6151
R2601 B.n582 B.n581 10.6151
R2602 B.n581 B.n126 10.6151
R2603 B.n577 B.n126 10.6151
R2604 B.n577 B.n576 10.6151
R2605 B.n576 B.n575 10.6151
R2606 B.n575 B.n128 10.6151
R2607 B.n571 B.n128 10.6151
R2608 B.n571 B.n570 10.6151
R2609 B.n570 B.n569 10.6151
R2610 B.n569 B.n130 10.6151
R2611 B.n565 B.n130 10.6151
R2612 B.n565 B.n564 10.6151
R2613 B.n564 B.n563 10.6151
R2614 B.n563 B.n132 10.6151
R2615 B.n559 B.n132 10.6151
R2616 B.n559 B.n558 10.6151
R2617 B.n558 B.n557 10.6151
R2618 B.n557 B.n134 10.6151
R2619 B.n553 B.n134 10.6151
R2620 B.n553 B.n552 10.6151
R2621 B.n552 B.n551 10.6151
R2622 B.n551 B.n136 10.6151
R2623 B.n547 B.n136 10.6151
R2624 B.n547 B.n546 10.6151
R2625 B.n546 B.n545 10.6151
R2626 B.n545 B.n138 10.6151
R2627 B.n541 B.n138 10.6151
R2628 B.n541 B.n540 10.6151
R2629 B.n540 B.n539 10.6151
R2630 B.n539 B.n140 10.6151
R2631 B.n535 B.n140 10.6151
R2632 B.n535 B.n534 10.6151
R2633 B.n534 B.n533 10.6151
R2634 B.n533 B.n142 10.6151
R2635 B.n529 B.n142 10.6151
R2636 B.n529 B.n528 10.6151
R2637 B.n528 B.n527 10.6151
R2638 B.n527 B.n144 10.6151
R2639 B.n523 B.n144 10.6151
R2640 B.n523 B.n522 10.6151
R2641 B.n522 B.n521 10.6151
R2642 B.n521 B.n146 10.6151
R2643 B.n241 B.n1 10.6151
R2644 B.n242 B.n241 10.6151
R2645 B.n243 B.n242 10.6151
R2646 B.n243 B.n238 10.6151
R2647 B.n247 B.n238 10.6151
R2648 B.n248 B.n247 10.6151
R2649 B.n249 B.n248 10.6151
R2650 B.n249 B.n236 10.6151
R2651 B.n253 B.n236 10.6151
R2652 B.n254 B.n253 10.6151
R2653 B.n255 B.n254 10.6151
R2654 B.n255 B.n234 10.6151
R2655 B.n259 B.n234 10.6151
R2656 B.n260 B.n259 10.6151
R2657 B.n261 B.n260 10.6151
R2658 B.n261 B.n232 10.6151
R2659 B.n265 B.n232 10.6151
R2660 B.n266 B.n265 10.6151
R2661 B.n267 B.n266 10.6151
R2662 B.n267 B.n230 10.6151
R2663 B.n271 B.n230 10.6151
R2664 B.n272 B.n271 10.6151
R2665 B.n273 B.n272 10.6151
R2666 B.n273 B.n228 10.6151
R2667 B.n277 B.n228 10.6151
R2668 B.n278 B.n277 10.6151
R2669 B.n279 B.n278 10.6151
R2670 B.n279 B.n226 10.6151
R2671 B.n283 B.n226 10.6151
R2672 B.n284 B.n283 10.6151
R2673 B.n285 B.n284 10.6151
R2674 B.n285 B.n224 10.6151
R2675 B.n289 B.n224 10.6151
R2676 B.n290 B.n289 10.6151
R2677 B.n291 B.n290 10.6151
R2678 B.n291 B.n222 10.6151
R2679 B.n295 B.n222 10.6151
R2680 B.n296 B.n295 10.6151
R2681 B.n297 B.n296 10.6151
R2682 B.n297 B.n220 10.6151
R2683 B.n301 B.n220 10.6151
R2684 B.n302 B.n301 10.6151
R2685 B.n303 B.n302 10.6151
R2686 B.n303 B.n218 10.6151
R2687 B.n307 B.n218 10.6151
R2688 B.n308 B.n307 10.6151
R2689 B.n309 B.n216 10.6151
R2690 B.n313 B.n216 10.6151
R2691 B.n314 B.n313 10.6151
R2692 B.n315 B.n314 10.6151
R2693 B.n315 B.n214 10.6151
R2694 B.n319 B.n214 10.6151
R2695 B.n320 B.n319 10.6151
R2696 B.n321 B.n320 10.6151
R2697 B.n321 B.n212 10.6151
R2698 B.n325 B.n212 10.6151
R2699 B.n326 B.n325 10.6151
R2700 B.n327 B.n326 10.6151
R2701 B.n327 B.n210 10.6151
R2702 B.n331 B.n210 10.6151
R2703 B.n332 B.n331 10.6151
R2704 B.n333 B.n332 10.6151
R2705 B.n333 B.n208 10.6151
R2706 B.n337 B.n208 10.6151
R2707 B.n338 B.n337 10.6151
R2708 B.n339 B.n338 10.6151
R2709 B.n339 B.n206 10.6151
R2710 B.n343 B.n206 10.6151
R2711 B.n344 B.n343 10.6151
R2712 B.n345 B.n344 10.6151
R2713 B.n345 B.n204 10.6151
R2714 B.n349 B.n204 10.6151
R2715 B.n350 B.n349 10.6151
R2716 B.n351 B.n350 10.6151
R2717 B.n351 B.n202 10.6151
R2718 B.n355 B.n202 10.6151
R2719 B.n356 B.n355 10.6151
R2720 B.n357 B.n356 10.6151
R2721 B.n357 B.n200 10.6151
R2722 B.n361 B.n200 10.6151
R2723 B.n362 B.n361 10.6151
R2724 B.n363 B.n362 10.6151
R2725 B.n363 B.n198 10.6151
R2726 B.n367 B.n198 10.6151
R2727 B.n368 B.n367 10.6151
R2728 B.n369 B.n368 10.6151
R2729 B.n369 B.n196 10.6151
R2730 B.n373 B.n196 10.6151
R2731 B.n374 B.n373 10.6151
R2732 B.n375 B.n374 10.6151
R2733 B.n375 B.n194 10.6151
R2734 B.n379 B.n194 10.6151
R2735 B.n380 B.n379 10.6151
R2736 B.n381 B.n380 10.6151
R2737 B.n381 B.n192 10.6151
R2738 B.n385 B.n192 10.6151
R2739 B.n386 B.n385 10.6151
R2740 B.n387 B.n386 10.6151
R2741 B.n387 B.n190 10.6151
R2742 B.n391 B.n190 10.6151
R2743 B.n392 B.n391 10.6151
R2744 B.n393 B.n392 10.6151
R2745 B.n393 B.n188 10.6151
R2746 B.n397 B.n188 10.6151
R2747 B.n398 B.n397 10.6151
R2748 B.n399 B.n398 10.6151
R2749 B.n399 B.n186 10.6151
R2750 B.n403 B.n186 10.6151
R2751 B.n404 B.n403 10.6151
R2752 B.n406 B.n182 10.6151
R2753 B.n410 B.n182 10.6151
R2754 B.n411 B.n410 10.6151
R2755 B.n412 B.n411 10.6151
R2756 B.n412 B.n180 10.6151
R2757 B.n416 B.n180 10.6151
R2758 B.n417 B.n416 10.6151
R2759 B.n421 B.n417 10.6151
R2760 B.n425 B.n178 10.6151
R2761 B.n426 B.n425 10.6151
R2762 B.n427 B.n426 10.6151
R2763 B.n427 B.n176 10.6151
R2764 B.n431 B.n176 10.6151
R2765 B.n432 B.n431 10.6151
R2766 B.n433 B.n432 10.6151
R2767 B.n433 B.n174 10.6151
R2768 B.n437 B.n174 10.6151
R2769 B.n438 B.n437 10.6151
R2770 B.n439 B.n438 10.6151
R2771 B.n439 B.n172 10.6151
R2772 B.n443 B.n172 10.6151
R2773 B.n444 B.n443 10.6151
R2774 B.n445 B.n444 10.6151
R2775 B.n445 B.n170 10.6151
R2776 B.n449 B.n170 10.6151
R2777 B.n450 B.n449 10.6151
R2778 B.n451 B.n450 10.6151
R2779 B.n451 B.n168 10.6151
R2780 B.n455 B.n168 10.6151
R2781 B.n456 B.n455 10.6151
R2782 B.n457 B.n456 10.6151
R2783 B.n457 B.n166 10.6151
R2784 B.n461 B.n166 10.6151
R2785 B.n462 B.n461 10.6151
R2786 B.n463 B.n462 10.6151
R2787 B.n463 B.n164 10.6151
R2788 B.n467 B.n164 10.6151
R2789 B.n468 B.n467 10.6151
R2790 B.n469 B.n468 10.6151
R2791 B.n469 B.n162 10.6151
R2792 B.n473 B.n162 10.6151
R2793 B.n474 B.n473 10.6151
R2794 B.n475 B.n474 10.6151
R2795 B.n475 B.n160 10.6151
R2796 B.n479 B.n160 10.6151
R2797 B.n480 B.n479 10.6151
R2798 B.n481 B.n480 10.6151
R2799 B.n481 B.n158 10.6151
R2800 B.n485 B.n158 10.6151
R2801 B.n486 B.n485 10.6151
R2802 B.n487 B.n486 10.6151
R2803 B.n487 B.n156 10.6151
R2804 B.n491 B.n156 10.6151
R2805 B.n492 B.n491 10.6151
R2806 B.n493 B.n492 10.6151
R2807 B.n493 B.n154 10.6151
R2808 B.n497 B.n154 10.6151
R2809 B.n498 B.n497 10.6151
R2810 B.n499 B.n498 10.6151
R2811 B.n499 B.n152 10.6151
R2812 B.n503 B.n152 10.6151
R2813 B.n504 B.n503 10.6151
R2814 B.n505 B.n504 10.6151
R2815 B.n505 B.n150 10.6151
R2816 B.n509 B.n150 10.6151
R2817 B.n510 B.n509 10.6151
R2818 B.n511 B.n510 10.6151
R2819 B.n511 B.n148 10.6151
R2820 B.n515 B.n148 10.6151
R2821 B.n516 B.n515 10.6151
R2822 B.n517 B.n516 10.6151
R2823 B.n941 B.n0 8.11757
R2824 B.n941 B.n1 8.11757
R2825 B.n773 B.n772 6.5566
R2826 B.n760 B.n66 6.5566
R2827 B.n406 B.n405 6.5566
R2828 B.n421 B.n420 6.5566
R2829 B.n774 B.n773 4.05904
R2830 B.n757 B.n66 4.05904
R2831 B.n405 B.n404 4.05904
R2832 B.n420 B.n178 4.05904
R2833 VN.n7 VN.t6 230.635
R2834 VN.n34 VN.t3 230.635
R2835 VN.n6 VN.t7 198.519
R2836 VN.n17 VN.t2 198.519
R2837 VN.n25 VN.t5 198.519
R2838 VN.n33 VN.t4 198.519
R2839 VN.n44 VN.t0 198.519
R2840 VN.n52 VN.t1 198.519
R2841 VN.n51 VN.n27 161.3
R2842 VN.n50 VN.n49 161.3
R2843 VN.n48 VN.n28 161.3
R2844 VN.n47 VN.n46 161.3
R2845 VN.n45 VN.n29 161.3
R2846 VN.n43 VN.n42 161.3
R2847 VN.n41 VN.n30 161.3
R2848 VN.n40 VN.n39 161.3
R2849 VN.n38 VN.n31 161.3
R2850 VN.n37 VN.n36 161.3
R2851 VN.n35 VN.n32 161.3
R2852 VN.n24 VN.n0 161.3
R2853 VN.n23 VN.n22 161.3
R2854 VN.n21 VN.n1 161.3
R2855 VN.n20 VN.n19 161.3
R2856 VN.n18 VN.n2 161.3
R2857 VN.n16 VN.n15 161.3
R2858 VN.n14 VN.n3 161.3
R2859 VN.n13 VN.n12 161.3
R2860 VN.n11 VN.n4 161.3
R2861 VN.n10 VN.n9 161.3
R2862 VN.n8 VN.n5 161.3
R2863 VN.n26 VN.n25 96.7304
R2864 VN.n53 VN.n52 96.7304
R2865 VN.n7 VN.n6 67.322
R2866 VN.n34 VN.n33 67.322
R2867 VN.n12 VN.n11 56.4773
R2868 VN.n39 VN.n38 56.4773
R2869 VN VN.n53 55.7102
R2870 VN.n19 VN.n1 46.253
R2871 VN.n46 VN.n28 46.253
R2872 VN.n23 VN.n1 34.5682
R2873 VN.n50 VN.n28 34.5682
R2874 VN.n10 VN.n5 24.3439
R2875 VN.n11 VN.n10 24.3439
R2876 VN.n12 VN.n3 24.3439
R2877 VN.n16 VN.n3 24.3439
R2878 VN.n19 VN.n18 24.3439
R2879 VN.n24 VN.n23 24.3439
R2880 VN.n38 VN.n37 24.3439
R2881 VN.n37 VN.n32 24.3439
R2882 VN.n46 VN.n45 24.3439
R2883 VN.n43 VN.n30 24.3439
R2884 VN.n39 VN.n30 24.3439
R2885 VN.n51 VN.n50 24.3439
R2886 VN.n18 VN.n17 19.7187
R2887 VN.n45 VN.n44 19.7187
R2888 VN.n25 VN.n24 13.8763
R2889 VN.n52 VN.n51 13.8763
R2890 VN.n35 VN.n34 9.62344
R2891 VN.n8 VN.n7 9.62344
R2892 VN.n6 VN.n5 4.62575
R2893 VN.n17 VN.n16 4.62575
R2894 VN.n33 VN.n32 4.62575
R2895 VN.n44 VN.n43 4.62575
R2896 VN.n53 VN.n27 0.278398
R2897 VN.n26 VN.n0 0.278398
R2898 VN.n49 VN.n27 0.189894
R2899 VN.n49 VN.n48 0.189894
R2900 VN.n48 VN.n47 0.189894
R2901 VN.n47 VN.n29 0.189894
R2902 VN.n42 VN.n29 0.189894
R2903 VN.n42 VN.n41 0.189894
R2904 VN.n41 VN.n40 0.189894
R2905 VN.n40 VN.n31 0.189894
R2906 VN.n36 VN.n31 0.189894
R2907 VN.n36 VN.n35 0.189894
R2908 VN.n9 VN.n8 0.189894
R2909 VN.n9 VN.n4 0.189894
R2910 VN.n13 VN.n4 0.189894
R2911 VN.n14 VN.n13 0.189894
R2912 VN.n15 VN.n14 0.189894
R2913 VN.n15 VN.n2 0.189894
R2914 VN.n20 VN.n2 0.189894
R2915 VN.n21 VN.n20 0.189894
R2916 VN.n22 VN.n21 0.189894
R2917 VN.n22 VN.n0 0.189894
R2918 VN VN.n26 0.153422
R2919 VDD2.n2 VDD2.n1 71.2745
R2920 VDD2.n2 VDD2.n0 71.2745
R2921 VDD2 VDD2.n5 71.2716
R2922 VDD2.n4 VDD2.n3 70.1705
R2923 VDD2.n4 VDD2.n2 50.9093
R2924 VDD2.n5 VDD2.t3 1.67257
R2925 VDD2.n5 VDD2.t4 1.67257
R2926 VDD2.n3 VDD2.t6 1.67257
R2927 VDD2.n3 VDD2.t7 1.67257
R2928 VDD2.n1 VDD2.t5 1.67257
R2929 VDD2.n1 VDD2.t2 1.67257
R2930 VDD2.n0 VDD2.t1 1.67257
R2931 VDD2.n0 VDD2.t0 1.67257
R2932 VDD2 VDD2.n4 1.21817
C0 VDD1 VP 13.879701f
C1 VDD2 B 1.86635f
C2 VDD2 VP 0.493507f
C3 VN VTAIL 13.5238f
C4 w_n3660_n4856# B 11.8343f
C5 w_n3660_n4856# VP 8.00451f
C6 VDD1 VDD2 1.65046f
C7 VDD1 w_n3660_n4856# 2.07241f
C8 VN B 1.25318f
C9 VDD2 w_n3660_n4856# 2.17705f
C10 VTAIL B 7.2762f
C11 VN VP 8.75241f
C12 VTAIL VP 13.537901f
C13 VDD1 VN 0.150669f
C14 VDD1 VTAIL 10.691401f
C15 VDD2 VN 13.538099f
C16 VDD2 VTAIL 10.744201f
C17 VN w_n3660_n4856# 7.53008f
C18 B VP 2.04722f
C19 VTAIL w_n3660_n4856# 5.88347f
C20 VDD1 B 1.77788f
C21 VDD2 VSUBS 1.987937f
C22 VDD1 VSUBS 2.59261f
C23 VTAIL VSUBS 1.63845f
C24 VN VSUBS 6.7663f
C25 VP VSUBS 3.614202f
C26 B VSUBS 5.36046f
C27 w_n3660_n4856# VSUBS 0.217097p
C28 VDD2.t1 VSUBS 0.407925f
C29 VDD2.t0 VSUBS 0.407925f
C30 VDD2.n0 VSUBS 3.45136f
C31 VDD2.t5 VSUBS 0.407925f
C32 VDD2.t2 VSUBS 0.407925f
C33 VDD2.n1 VSUBS 3.45136f
C34 VDD2.n2 VSUBS 4.41012f
C35 VDD2.t6 VSUBS 0.407925f
C36 VDD2.t7 VSUBS 0.407925f
C37 VDD2.n3 VSUBS 3.43876f
C38 VDD2.n4 VSUBS 3.93421f
C39 VDD2.t3 VSUBS 0.407925f
C40 VDD2.t4 VSUBS 0.407925f
C41 VDD2.n5 VSUBS 3.45131f
C42 VN.n0 VSUBS 0.035828f
C43 VN.t5 VSUBS 3.43393f
C44 VN.n1 VSUBS 0.023283f
C45 VN.n2 VSUBS 0.027174f
C46 VN.t2 VSUBS 3.43393f
C47 VN.n3 VSUBS 0.050899f
C48 VN.n4 VSUBS 0.027174f
C49 VN.n5 VSUBS 0.030543f
C50 VN.t6 VSUBS 3.62103f
C51 VN.t7 VSUBS 3.43393f
C52 VN.n6 VSUBS 1.25682f
C53 VN.n7 VSUBS 1.25035f
C54 VN.n8 VSUBS 0.235707f
C55 VN.n9 VSUBS 0.027174f
C56 VN.n10 VSUBS 0.050899f
C57 VN.n11 VSUBS 0.039842f
C58 VN.n12 VSUBS 0.039842f
C59 VN.n13 VSUBS 0.027174f
C60 VN.n14 VSUBS 0.027174f
C61 VN.n15 VSUBS 0.027174f
C62 VN.n16 VSUBS 0.030543f
C63 VN.n17 VSUBS 1.18974f
C64 VN.n18 VSUBS 0.046124f
C65 VN.n19 VSUBS 0.05209f
C66 VN.n20 VSUBS 0.027174f
C67 VN.n21 VSUBS 0.027174f
C68 VN.n22 VSUBS 0.027174f
C69 VN.n23 VSUBS 0.055211f
C70 VN.n24 VSUBS 0.040093f
C71 VN.n25 VSUBS 1.27855f
C72 VN.n26 VSUBS 0.039517f
C73 VN.n27 VSUBS 0.035828f
C74 VN.t1 VSUBS 3.43393f
C75 VN.n28 VSUBS 0.023283f
C76 VN.n29 VSUBS 0.027174f
C77 VN.t0 VSUBS 3.43393f
C78 VN.n30 VSUBS 0.050899f
C79 VN.n31 VSUBS 0.027174f
C80 VN.n32 VSUBS 0.030543f
C81 VN.t3 VSUBS 3.62103f
C82 VN.t4 VSUBS 3.43393f
C83 VN.n33 VSUBS 1.25682f
C84 VN.n34 VSUBS 1.25035f
C85 VN.n35 VSUBS 0.235707f
C86 VN.n36 VSUBS 0.027174f
C87 VN.n37 VSUBS 0.050899f
C88 VN.n38 VSUBS 0.039842f
C89 VN.n39 VSUBS 0.039842f
C90 VN.n40 VSUBS 0.027174f
C91 VN.n41 VSUBS 0.027174f
C92 VN.n42 VSUBS 0.027174f
C93 VN.n43 VSUBS 0.030543f
C94 VN.n44 VSUBS 1.18974f
C95 VN.n45 VSUBS 0.046124f
C96 VN.n46 VSUBS 0.05209f
C97 VN.n47 VSUBS 0.027174f
C98 VN.n48 VSUBS 0.027174f
C99 VN.n49 VSUBS 0.027174f
C100 VN.n50 VSUBS 0.055211f
C101 VN.n51 VSUBS 0.040093f
C102 VN.n52 VSUBS 1.27855f
C103 VN.n53 VSUBS 1.76275f
C104 B.n0 VSUBS 0.00596f
C105 B.n1 VSUBS 0.00596f
C106 B.n2 VSUBS 0.008814f
C107 B.n3 VSUBS 0.006754f
C108 B.n4 VSUBS 0.006754f
C109 B.n5 VSUBS 0.006754f
C110 B.n6 VSUBS 0.006754f
C111 B.n7 VSUBS 0.006754f
C112 B.n8 VSUBS 0.006754f
C113 B.n9 VSUBS 0.006754f
C114 B.n10 VSUBS 0.006754f
C115 B.n11 VSUBS 0.006754f
C116 B.n12 VSUBS 0.006754f
C117 B.n13 VSUBS 0.006754f
C118 B.n14 VSUBS 0.006754f
C119 B.n15 VSUBS 0.006754f
C120 B.n16 VSUBS 0.006754f
C121 B.n17 VSUBS 0.006754f
C122 B.n18 VSUBS 0.006754f
C123 B.n19 VSUBS 0.006754f
C124 B.n20 VSUBS 0.006754f
C125 B.n21 VSUBS 0.006754f
C126 B.n22 VSUBS 0.006754f
C127 B.n23 VSUBS 0.006754f
C128 B.n24 VSUBS 0.006754f
C129 B.n25 VSUBS 0.014949f
C130 B.n26 VSUBS 0.006754f
C131 B.n27 VSUBS 0.006754f
C132 B.n28 VSUBS 0.006754f
C133 B.n29 VSUBS 0.006754f
C134 B.n30 VSUBS 0.006754f
C135 B.n31 VSUBS 0.006754f
C136 B.n32 VSUBS 0.006754f
C137 B.n33 VSUBS 0.006754f
C138 B.n34 VSUBS 0.006754f
C139 B.n35 VSUBS 0.006754f
C140 B.n36 VSUBS 0.006754f
C141 B.n37 VSUBS 0.006754f
C142 B.n38 VSUBS 0.006754f
C143 B.n39 VSUBS 0.006754f
C144 B.n40 VSUBS 0.006754f
C145 B.n41 VSUBS 0.006754f
C146 B.n42 VSUBS 0.006754f
C147 B.n43 VSUBS 0.006754f
C148 B.n44 VSUBS 0.006754f
C149 B.n45 VSUBS 0.006754f
C150 B.n46 VSUBS 0.006754f
C151 B.n47 VSUBS 0.006754f
C152 B.n48 VSUBS 0.006754f
C153 B.n49 VSUBS 0.006754f
C154 B.n50 VSUBS 0.006754f
C155 B.n51 VSUBS 0.006754f
C156 B.n52 VSUBS 0.006754f
C157 B.n53 VSUBS 0.006754f
C158 B.n54 VSUBS 0.006754f
C159 B.n55 VSUBS 0.006754f
C160 B.n56 VSUBS 0.006754f
C161 B.n57 VSUBS 0.006754f
C162 B.t4 VSUBS 0.372417f
C163 B.t5 VSUBS 0.402434f
C164 B.t3 VSUBS 1.93909f
C165 B.n58 VSUBS 0.603818f
C166 B.n59 VSUBS 0.332801f
C167 B.n60 VSUBS 0.006754f
C168 B.n61 VSUBS 0.006754f
C169 B.n62 VSUBS 0.006754f
C170 B.n63 VSUBS 0.006754f
C171 B.t10 VSUBS 0.37242f
C172 B.t11 VSUBS 0.402437f
C173 B.t9 VSUBS 1.93909f
C174 B.n64 VSUBS 0.603815f
C175 B.n65 VSUBS 0.332797f
C176 B.n66 VSUBS 0.015649f
C177 B.n67 VSUBS 0.006754f
C178 B.n68 VSUBS 0.006754f
C179 B.n69 VSUBS 0.006754f
C180 B.n70 VSUBS 0.006754f
C181 B.n71 VSUBS 0.006754f
C182 B.n72 VSUBS 0.006754f
C183 B.n73 VSUBS 0.006754f
C184 B.n74 VSUBS 0.006754f
C185 B.n75 VSUBS 0.006754f
C186 B.n76 VSUBS 0.006754f
C187 B.n77 VSUBS 0.006754f
C188 B.n78 VSUBS 0.006754f
C189 B.n79 VSUBS 0.006754f
C190 B.n80 VSUBS 0.006754f
C191 B.n81 VSUBS 0.006754f
C192 B.n82 VSUBS 0.006754f
C193 B.n83 VSUBS 0.006754f
C194 B.n84 VSUBS 0.006754f
C195 B.n85 VSUBS 0.006754f
C196 B.n86 VSUBS 0.006754f
C197 B.n87 VSUBS 0.006754f
C198 B.n88 VSUBS 0.006754f
C199 B.n89 VSUBS 0.006754f
C200 B.n90 VSUBS 0.006754f
C201 B.n91 VSUBS 0.006754f
C202 B.n92 VSUBS 0.006754f
C203 B.n93 VSUBS 0.006754f
C204 B.n94 VSUBS 0.006754f
C205 B.n95 VSUBS 0.006754f
C206 B.n96 VSUBS 0.006754f
C207 B.n97 VSUBS 0.006754f
C208 B.n98 VSUBS 0.01624f
C209 B.n99 VSUBS 0.006754f
C210 B.n100 VSUBS 0.006754f
C211 B.n101 VSUBS 0.006754f
C212 B.n102 VSUBS 0.006754f
C213 B.n103 VSUBS 0.006754f
C214 B.n104 VSUBS 0.006754f
C215 B.n105 VSUBS 0.006754f
C216 B.n106 VSUBS 0.006754f
C217 B.n107 VSUBS 0.006754f
C218 B.n108 VSUBS 0.006754f
C219 B.n109 VSUBS 0.006754f
C220 B.n110 VSUBS 0.006754f
C221 B.n111 VSUBS 0.006754f
C222 B.n112 VSUBS 0.006754f
C223 B.n113 VSUBS 0.006754f
C224 B.n114 VSUBS 0.006754f
C225 B.n115 VSUBS 0.006754f
C226 B.n116 VSUBS 0.006754f
C227 B.n117 VSUBS 0.006754f
C228 B.n118 VSUBS 0.006754f
C229 B.n119 VSUBS 0.006754f
C230 B.n120 VSUBS 0.006754f
C231 B.n121 VSUBS 0.006754f
C232 B.n122 VSUBS 0.006754f
C233 B.n123 VSUBS 0.006754f
C234 B.n124 VSUBS 0.006754f
C235 B.n125 VSUBS 0.006754f
C236 B.n126 VSUBS 0.006754f
C237 B.n127 VSUBS 0.006754f
C238 B.n128 VSUBS 0.006754f
C239 B.n129 VSUBS 0.006754f
C240 B.n130 VSUBS 0.006754f
C241 B.n131 VSUBS 0.006754f
C242 B.n132 VSUBS 0.006754f
C243 B.n133 VSUBS 0.006754f
C244 B.n134 VSUBS 0.006754f
C245 B.n135 VSUBS 0.006754f
C246 B.n136 VSUBS 0.006754f
C247 B.n137 VSUBS 0.006754f
C248 B.n138 VSUBS 0.006754f
C249 B.n139 VSUBS 0.006754f
C250 B.n140 VSUBS 0.006754f
C251 B.n141 VSUBS 0.006754f
C252 B.n142 VSUBS 0.006754f
C253 B.n143 VSUBS 0.006754f
C254 B.n144 VSUBS 0.006754f
C255 B.n145 VSUBS 0.006754f
C256 B.n146 VSUBS 0.015764f
C257 B.n147 VSUBS 0.006754f
C258 B.n148 VSUBS 0.006754f
C259 B.n149 VSUBS 0.006754f
C260 B.n150 VSUBS 0.006754f
C261 B.n151 VSUBS 0.006754f
C262 B.n152 VSUBS 0.006754f
C263 B.n153 VSUBS 0.006754f
C264 B.n154 VSUBS 0.006754f
C265 B.n155 VSUBS 0.006754f
C266 B.n156 VSUBS 0.006754f
C267 B.n157 VSUBS 0.006754f
C268 B.n158 VSUBS 0.006754f
C269 B.n159 VSUBS 0.006754f
C270 B.n160 VSUBS 0.006754f
C271 B.n161 VSUBS 0.006754f
C272 B.n162 VSUBS 0.006754f
C273 B.n163 VSUBS 0.006754f
C274 B.n164 VSUBS 0.006754f
C275 B.n165 VSUBS 0.006754f
C276 B.n166 VSUBS 0.006754f
C277 B.n167 VSUBS 0.006754f
C278 B.n168 VSUBS 0.006754f
C279 B.n169 VSUBS 0.006754f
C280 B.n170 VSUBS 0.006754f
C281 B.n171 VSUBS 0.006754f
C282 B.n172 VSUBS 0.006754f
C283 B.n173 VSUBS 0.006754f
C284 B.n174 VSUBS 0.006754f
C285 B.n175 VSUBS 0.006754f
C286 B.n176 VSUBS 0.006754f
C287 B.n177 VSUBS 0.006754f
C288 B.n178 VSUBS 0.004668f
C289 B.n179 VSUBS 0.006754f
C290 B.n180 VSUBS 0.006754f
C291 B.n181 VSUBS 0.006754f
C292 B.n182 VSUBS 0.006754f
C293 B.n183 VSUBS 0.006754f
C294 B.t2 VSUBS 0.372417f
C295 B.t1 VSUBS 0.402434f
C296 B.t0 VSUBS 1.93909f
C297 B.n184 VSUBS 0.603818f
C298 B.n185 VSUBS 0.332801f
C299 B.n186 VSUBS 0.006754f
C300 B.n187 VSUBS 0.006754f
C301 B.n188 VSUBS 0.006754f
C302 B.n189 VSUBS 0.006754f
C303 B.n190 VSUBS 0.006754f
C304 B.n191 VSUBS 0.006754f
C305 B.n192 VSUBS 0.006754f
C306 B.n193 VSUBS 0.006754f
C307 B.n194 VSUBS 0.006754f
C308 B.n195 VSUBS 0.006754f
C309 B.n196 VSUBS 0.006754f
C310 B.n197 VSUBS 0.006754f
C311 B.n198 VSUBS 0.006754f
C312 B.n199 VSUBS 0.006754f
C313 B.n200 VSUBS 0.006754f
C314 B.n201 VSUBS 0.006754f
C315 B.n202 VSUBS 0.006754f
C316 B.n203 VSUBS 0.006754f
C317 B.n204 VSUBS 0.006754f
C318 B.n205 VSUBS 0.006754f
C319 B.n206 VSUBS 0.006754f
C320 B.n207 VSUBS 0.006754f
C321 B.n208 VSUBS 0.006754f
C322 B.n209 VSUBS 0.006754f
C323 B.n210 VSUBS 0.006754f
C324 B.n211 VSUBS 0.006754f
C325 B.n212 VSUBS 0.006754f
C326 B.n213 VSUBS 0.006754f
C327 B.n214 VSUBS 0.006754f
C328 B.n215 VSUBS 0.006754f
C329 B.n216 VSUBS 0.006754f
C330 B.n217 VSUBS 0.014949f
C331 B.n218 VSUBS 0.006754f
C332 B.n219 VSUBS 0.006754f
C333 B.n220 VSUBS 0.006754f
C334 B.n221 VSUBS 0.006754f
C335 B.n222 VSUBS 0.006754f
C336 B.n223 VSUBS 0.006754f
C337 B.n224 VSUBS 0.006754f
C338 B.n225 VSUBS 0.006754f
C339 B.n226 VSUBS 0.006754f
C340 B.n227 VSUBS 0.006754f
C341 B.n228 VSUBS 0.006754f
C342 B.n229 VSUBS 0.006754f
C343 B.n230 VSUBS 0.006754f
C344 B.n231 VSUBS 0.006754f
C345 B.n232 VSUBS 0.006754f
C346 B.n233 VSUBS 0.006754f
C347 B.n234 VSUBS 0.006754f
C348 B.n235 VSUBS 0.006754f
C349 B.n236 VSUBS 0.006754f
C350 B.n237 VSUBS 0.006754f
C351 B.n238 VSUBS 0.006754f
C352 B.n239 VSUBS 0.006754f
C353 B.n240 VSUBS 0.006754f
C354 B.n241 VSUBS 0.006754f
C355 B.n242 VSUBS 0.006754f
C356 B.n243 VSUBS 0.006754f
C357 B.n244 VSUBS 0.006754f
C358 B.n245 VSUBS 0.006754f
C359 B.n246 VSUBS 0.006754f
C360 B.n247 VSUBS 0.006754f
C361 B.n248 VSUBS 0.006754f
C362 B.n249 VSUBS 0.006754f
C363 B.n250 VSUBS 0.006754f
C364 B.n251 VSUBS 0.006754f
C365 B.n252 VSUBS 0.006754f
C366 B.n253 VSUBS 0.006754f
C367 B.n254 VSUBS 0.006754f
C368 B.n255 VSUBS 0.006754f
C369 B.n256 VSUBS 0.006754f
C370 B.n257 VSUBS 0.006754f
C371 B.n258 VSUBS 0.006754f
C372 B.n259 VSUBS 0.006754f
C373 B.n260 VSUBS 0.006754f
C374 B.n261 VSUBS 0.006754f
C375 B.n262 VSUBS 0.006754f
C376 B.n263 VSUBS 0.006754f
C377 B.n264 VSUBS 0.006754f
C378 B.n265 VSUBS 0.006754f
C379 B.n266 VSUBS 0.006754f
C380 B.n267 VSUBS 0.006754f
C381 B.n268 VSUBS 0.006754f
C382 B.n269 VSUBS 0.006754f
C383 B.n270 VSUBS 0.006754f
C384 B.n271 VSUBS 0.006754f
C385 B.n272 VSUBS 0.006754f
C386 B.n273 VSUBS 0.006754f
C387 B.n274 VSUBS 0.006754f
C388 B.n275 VSUBS 0.006754f
C389 B.n276 VSUBS 0.006754f
C390 B.n277 VSUBS 0.006754f
C391 B.n278 VSUBS 0.006754f
C392 B.n279 VSUBS 0.006754f
C393 B.n280 VSUBS 0.006754f
C394 B.n281 VSUBS 0.006754f
C395 B.n282 VSUBS 0.006754f
C396 B.n283 VSUBS 0.006754f
C397 B.n284 VSUBS 0.006754f
C398 B.n285 VSUBS 0.006754f
C399 B.n286 VSUBS 0.006754f
C400 B.n287 VSUBS 0.006754f
C401 B.n288 VSUBS 0.006754f
C402 B.n289 VSUBS 0.006754f
C403 B.n290 VSUBS 0.006754f
C404 B.n291 VSUBS 0.006754f
C405 B.n292 VSUBS 0.006754f
C406 B.n293 VSUBS 0.006754f
C407 B.n294 VSUBS 0.006754f
C408 B.n295 VSUBS 0.006754f
C409 B.n296 VSUBS 0.006754f
C410 B.n297 VSUBS 0.006754f
C411 B.n298 VSUBS 0.006754f
C412 B.n299 VSUBS 0.006754f
C413 B.n300 VSUBS 0.006754f
C414 B.n301 VSUBS 0.006754f
C415 B.n302 VSUBS 0.006754f
C416 B.n303 VSUBS 0.006754f
C417 B.n304 VSUBS 0.006754f
C418 B.n305 VSUBS 0.006754f
C419 B.n306 VSUBS 0.006754f
C420 B.n307 VSUBS 0.006754f
C421 B.n308 VSUBS 0.014949f
C422 B.n309 VSUBS 0.01624f
C423 B.n310 VSUBS 0.01624f
C424 B.n311 VSUBS 0.006754f
C425 B.n312 VSUBS 0.006754f
C426 B.n313 VSUBS 0.006754f
C427 B.n314 VSUBS 0.006754f
C428 B.n315 VSUBS 0.006754f
C429 B.n316 VSUBS 0.006754f
C430 B.n317 VSUBS 0.006754f
C431 B.n318 VSUBS 0.006754f
C432 B.n319 VSUBS 0.006754f
C433 B.n320 VSUBS 0.006754f
C434 B.n321 VSUBS 0.006754f
C435 B.n322 VSUBS 0.006754f
C436 B.n323 VSUBS 0.006754f
C437 B.n324 VSUBS 0.006754f
C438 B.n325 VSUBS 0.006754f
C439 B.n326 VSUBS 0.006754f
C440 B.n327 VSUBS 0.006754f
C441 B.n328 VSUBS 0.006754f
C442 B.n329 VSUBS 0.006754f
C443 B.n330 VSUBS 0.006754f
C444 B.n331 VSUBS 0.006754f
C445 B.n332 VSUBS 0.006754f
C446 B.n333 VSUBS 0.006754f
C447 B.n334 VSUBS 0.006754f
C448 B.n335 VSUBS 0.006754f
C449 B.n336 VSUBS 0.006754f
C450 B.n337 VSUBS 0.006754f
C451 B.n338 VSUBS 0.006754f
C452 B.n339 VSUBS 0.006754f
C453 B.n340 VSUBS 0.006754f
C454 B.n341 VSUBS 0.006754f
C455 B.n342 VSUBS 0.006754f
C456 B.n343 VSUBS 0.006754f
C457 B.n344 VSUBS 0.006754f
C458 B.n345 VSUBS 0.006754f
C459 B.n346 VSUBS 0.006754f
C460 B.n347 VSUBS 0.006754f
C461 B.n348 VSUBS 0.006754f
C462 B.n349 VSUBS 0.006754f
C463 B.n350 VSUBS 0.006754f
C464 B.n351 VSUBS 0.006754f
C465 B.n352 VSUBS 0.006754f
C466 B.n353 VSUBS 0.006754f
C467 B.n354 VSUBS 0.006754f
C468 B.n355 VSUBS 0.006754f
C469 B.n356 VSUBS 0.006754f
C470 B.n357 VSUBS 0.006754f
C471 B.n358 VSUBS 0.006754f
C472 B.n359 VSUBS 0.006754f
C473 B.n360 VSUBS 0.006754f
C474 B.n361 VSUBS 0.006754f
C475 B.n362 VSUBS 0.006754f
C476 B.n363 VSUBS 0.006754f
C477 B.n364 VSUBS 0.006754f
C478 B.n365 VSUBS 0.006754f
C479 B.n366 VSUBS 0.006754f
C480 B.n367 VSUBS 0.006754f
C481 B.n368 VSUBS 0.006754f
C482 B.n369 VSUBS 0.006754f
C483 B.n370 VSUBS 0.006754f
C484 B.n371 VSUBS 0.006754f
C485 B.n372 VSUBS 0.006754f
C486 B.n373 VSUBS 0.006754f
C487 B.n374 VSUBS 0.006754f
C488 B.n375 VSUBS 0.006754f
C489 B.n376 VSUBS 0.006754f
C490 B.n377 VSUBS 0.006754f
C491 B.n378 VSUBS 0.006754f
C492 B.n379 VSUBS 0.006754f
C493 B.n380 VSUBS 0.006754f
C494 B.n381 VSUBS 0.006754f
C495 B.n382 VSUBS 0.006754f
C496 B.n383 VSUBS 0.006754f
C497 B.n384 VSUBS 0.006754f
C498 B.n385 VSUBS 0.006754f
C499 B.n386 VSUBS 0.006754f
C500 B.n387 VSUBS 0.006754f
C501 B.n388 VSUBS 0.006754f
C502 B.n389 VSUBS 0.006754f
C503 B.n390 VSUBS 0.006754f
C504 B.n391 VSUBS 0.006754f
C505 B.n392 VSUBS 0.006754f
C506 B.n393 VSUBS 0.006754f
C507 B.n394 VSUBS 0.006754f
C508 B.n395 VSUBS 0.006754f
C509 B.n396 VSUBS 0.006754f
C510 B.n397 VSUBS 0.006754f
C511 B.n398 VSUBS 0.006754f
C512 B.n399 VSUBS 0.006754f
C513 B.n400 VSUBS 0.006754f
C514 B.n401 VSUBS 0.006754f
C515 B.n402 VSUBS 0.006754f
C516 B.n403 VSUBS 0.006754f
C517 B.n404 VSUBS 0.004668f
C518 B.n405 VSUBS 0.015649f
C519 B.n406 VSUBS 0.005463f
C520 B.n407 VSUBS 0.006754f
C521 B.n408 VSUBS 0.006754f
C522 B.n409 VSUBS 0.006754f
C523 B.n410 VSUBS 0.006754f
C524 B.n411 VSUBS 0.006754f
C525 B.n412 VSUBS 0.006754f
C526 B.n413 VSUBS 0.006754f
C527 B.n414 VSUBS 0.006754f
C528 B.n415 VSUBS 0.006754f
C529 B.n416 VSUBS 0.006754f
C530 B.n417 VSUBS 0.006754f
C531 B.t8 VSUBS 0.37242f
C532 B.t7 VSUBS 0.402437f
C533 B.t6 VSUBS 1.93909f
C534 B.n418 VSUBS 0.603815f
C535 B.n419 VSUBS 0.332797f
C536 B.n420 VSUBS 0.015649f
C537 B.n421 VSUBS 0.005463f
C538 B.n422 VSUBS 0.006754f
C539 B.n423 VSUBS 0.006754f
C540 B.n424 VSUBS 0.006754f
C541 B.n425 VSUBS 0.006754f
C542 B.n426 VSUBS 0.006754f
C543 B.n427 VSUBS 0.006754f
C544 B.n428 VSUBS 0.006754f
C545 B.n429 VSUBS 0.006754f
C546 B.n430 VSUBS 0.006754f
C547 B.n431 VSUBS 0.006754f
C548 B.n432 VSUBS 0.006754f
C549 B.n433 VSUBS 0.006754f
C550 B.n434 VSUBS 0.006754f
C551 B.n435 VSUBS 0.006754f
C552 B.n436 VSUBS 0.006754f
C553 B.n437 VSUBS 0.006754f
C554 B.n438 VSUBS 0.006754f
C555 B.n439 VSUBS 0.006754f
C556 B.n440 VSUBS 0.006754f
C557 B.n441 VSUBS 0.006754f
C558 B.n442 VSUBS 0.006754f
C559 B.n443 VSUBS 0.006754f
C560 B.n444 VSUBS 0.006754f
C561 B.n445 VSUBS 0.006754f
C562 B.n446 VSUBS 0.006754f
C563 B.n447 VSUBS 0.006754f
C564 B.n448 VSUBS 0.006754f
C565 B.n449 VSUBS 0.006754f
C566 B.n450 VSUBS 0.006754f
C567 B.n451 VSUBS 0.006754f
C568 B.n452 VSUBS 0.006754f
C569 B.n453 VSUBS 0.006754f
C570 B.n454 VSUBS 0.006754f
C571 B.n455 VSUBS 0.006754f
C572 B.n456 VSUBS 0.006754f
C573 B.n457 VSUBS 0.006754f
C574 B.n458 VSUBS 0.006754f
C575 B.n459 VSUBS 0.006754f
C576 B.n460 VSUBS 0.006754f
C577 B.n461 VSUBS 0.006754f
C578 B.n462 VSUBS 0.006754f
C579 B.n463 VSUBS 0.006754f
C580 B.n464 VSUBS 0.006754f
C581 B.n465 VSUBS 0.006754f
C582 B.n466 VSUBS 0.006754f
C583 B.n467 VSUBS 0.006754f
C584 B.n468 VSUBS 0.006754f
C585 B.n469 VSUBS 0.006754f
C586 B.n470 VSUBS 0.006754f
C587 B.n471 VSUBS 0.006754f
C588 B.n472 VSUBS 0.006754f
C589 B.n473 VSUBS 0.006754f
C590 B.n474 VSUBS 0.006754f
C591 B.n475 VSUBS 0.006754f
C592 B.n476 VSUBS 0.006754f
C593 B.n477 VSUBS 0.006754f
C594 B.n478 VSUBS 0.006754f
C595 B.n479 VSUBS 0.006754f
C596 B.n480 VSUBS 0.006754f
C597 B.n481 VSUBS 0.006754f
C598 B.n482 VSUBS 0.006754f
C599 B.n483 VSUBS 0.006754f
C600 B.n484 VSUBS 0.006754f
C601 B.n485 VSUBS 0.006754f
C602 B.n486 VSUBS 0.006754f
C603 B.n487 VSUBS 0.006754f
C604 B.n488 VSUBS 0.006754f
C605 B.n489 VSUBS 0.006754f
C606 B.n490 VSUBS 0.006754f
C607 B.n491 VSUBS 0.006754f
C608 B.n492 VSUBS 0.006754f
C609 B.n493 VSUBS 0.006754f
C610 B.n494 VSUBS 0.006754f
C611 B.n495 VSUBS 0.006754f
C612 B.n496 VSUBS 0.006754f
C613 B.n497 VSUBS 0.006754f
C614 B.n498 VSUBS 0.006754f
C615 B.n499 VSUBS 0.006754f
C616 B.n500 VSUBS 0.006754f
C617 B.n501 VSUBS 0.006754f
C618 B.n502 VSUBS 0.006754f
C619 B.n503 VSUBS 0.006754f
C620 B.n504 VSUBS 0.006754f
C621 B.n505 VSUBS 0.006754f
C622 B.n506 VSUBS 0.006754f
C623 B.n507 VSUBS 0.006754f
C624 B.n508 VSUBS 0.006754f
C625 B.n509 VSUBS 0.006754f
C626 B.n510 VSUBS 0.006754f
C627 B.n511 VSUBS 0.006754f
C628 B.n512 VSUBS 0.006754f
C629 B.n513 VSUBS 0.006754f
C630 B.n514 VSUBS 0.006754f
C631 B.n515 VSUBS 0.006754f
C632 B.n516 VSUBS 0.006754f
C633 B.n517 VSUBS 0.015426f
C634 B.n518 VSUBS 0.01624f
C635 B.n519 VSUBS 0.014949f
C636 B.n520 VSUBS 0.006754f
C637 B.n521 VSUBS 0.006754f
C638 B.n522 VSUBS 0.006754f
C639 B.n523 VSUBS 0.006754f
C640 B.n524 VSUBS 0.006754f
C641 B.n525 VSUBS 0.006754f
C642 B.n526 VSUBS 0.006754f
C643 B.n527 VSUBS 0.006754f
C644 B.n528 VSUBS 0.006754f
C645 B.n529 VSUBS 0.006754f
C646 B.n530 VSUBS 0.006754f
C647 B.n531 VSUBS 0.006754f
C648 B.n532 VSUBS 0.006754f
C649 B.n533 VSUBS 0.006754f
C650 B.n534 VSUBS 0.006754f
C651 B.n535 VSUBS 0.006754f
C652 B.n536 VSUBS 0.006754f
C653 B.n537 VSUBS 0.006754f
C654 B.n538 VSUBS 0.006754f
C655 B.n539 VSUBS 0.006754f
C656 B.n540 VSUBS 0.006754f
C657 B.n541 VSUBS 0.006754f
C658 B.n542 VSUBS 0.006754f
C659 B.n543 VSUBS 0.006754f
C660 B.n544 VSUBS 0.006754f
C661 B.n545 VSUBS 0.006754f
C662 B.n546 VSUBS 0.006754f
C663 B.n547 VSUBS 0.006754f
C664 B.n548 VSUBS 0.006754f
C665 B.n549 VSUBS 0.006754f
C666 B.n550 VSUBS 0.006754f
C667 B.n551 VSUBS 0.006754f
C668 B.n552 VSUBS 0.006754f
C669 B.n553 VSUBS 0.006754f
C670 B.n554 VSUBS 0.006754f
C671 B.n555 VSUBS 0.006754f
C672 B.n556 VSUBS 0.006754f
C673 B.n557 VSUBS 0.006754f
C674 B.n558 VSUBS 0.006754f
C675 B.n559 VSUBS 0.006754f
C676 B.n560 VSUBS 0.006754f
C677 B.n561 VSUBS 0.006754f
C678 B.n562 VSUBS 0.006754f
C679 B.n563 VSUBS 0.006754f
C680 B.n564 VSUBS 0.006754f
C681 B.n565 VSUBS 0.006754f
C682 B.n566 VSUBS 0.006754f
C683 B.n567 VSUBS 0.006754f
C684 B.n568 VSUBS 0.006754f
C685 B.n569 VSUBS 0.006754f
C686 B.n570 VSUBS 0.006754f
C687 B.n571 VSUBS 0.006754f
C688 B.n572 VSUBS 0.006754f
C689 B.n573 VSUBS 0.006754f
C690 B.n574 VSUBS 0.006754f
C691 B.n575 VSUBS 0.006754f
C692 B.n576 VSUBS 0.006754f
C693 B.n577 VSUBS 0.006754f
C694 B.n578 VSUBS 0.006754f
C695 B.n579 VSUBS 0.006754f
C696 B.n580 VSUBS 0.006754f
C697 B.n581 VSUBS 0.006754f
C698 B.n582 VSUBS 0.006754f
C699 B.n583 VSUBS 0.006754f
C700 B.n584 VSUBS 0.006754f
C701 B.n585 VSUBS 0.006754f
C702 B.n586 VSUBS 0.006754f
C703 B.n587 VSUBS 0.006754f
C704 B.n588 VSUBS 0.006754f
C705 B.n589 VSUBS 0.006754f
C706 B.n590 VSUBS 0.006754f
C707 B.n591 VSUBS 0.006754f
C708 B.n592 VSUBS 0.006754f
C709 B.n593 VSUBS 0.006754f
C710 B.n594 VSUBS 0.006754f
C711 B.n595 VSUBS 0.006754f
C712 B.n596 VSUBS 0.006754f
C713 B.n597 VSUBS 0.006754f
C714 B.n598 VSUBS 0.006754f
C715 B.n599 VSUBS 0.006754f
C716 B.n600 VSUBS 0.006754f
C717 B.n601 VSUBS 0.006754f
C718 B.n602 VSUBS 0.006754f
C719 B.n603 VSUBS 0.006754f
C720 B.n604 VSUBS 0.006754f
C721 B.n605 VSUBS 0.006754f
C722 B.n606 VSUBS 0.006754f
C723 B.n607 VSUBS 0.006754f
C724 B.n608 VSUBS 0.006754f
C725 B.n609 VSUBS 0.006754f
C726 B.n610 VSUBS 0.006754f
C727 B.n611 VSUBS 0.006754f
C728 B.n612 VSUBS 0.006754f
C729 B.n613 VSUBS 0.006754f
C730 B.n614 VSUBS 0.006754f
C731 B.n615 VSUBS 0.006754f
C732 B.n616 VSUBS 0.006754f
C733 B.n617 VSUBS 0.006754f
C734 B.n618 VSUBS 0.006754f
C735 B.n619 VSUBS 0.006754f
C736 B.n620 VSUBS 0.006754f
C737 B.n621 VSUBS 0.006754f
C738 B.n622 VSUBS 0.006754f
C739 B.n623 VSUBS 0.006754f
C740 B.n624 VSUBS 0.006754f
C741 B.n625 VSUBS 0.006754f
C742 B.n626 VSUBS 0.006754f
C743 B.n627 VSUBS 0.006754f
C744 B.n628 VSUBS 0.006754f
C745 B.n629 VSUBS 0.006754f
C746 B.n630 VSUBS 0.006754f
C747 B.n631 VSUBS 0.006754f
C748 B.n632 VSUBS 0.006754f
C749 B.n633 VSUBS 0.006754f
C750 B.n634 VSUBS 0.006754f
C751 B.n635 VSUBS 0.006754f
C752 B.n636 VSUBS 0.006754f
C753 B.n637 VSUBS 0.006754f
C754 B.n638 VSUBS 0.006754f
C755 B.n639 VSUBS 0.006754f
C756 B.n640 VSUBS 0.006754f
C757 B.n641 VSUBS 0.006754f
C758 B.n642 VSUBS 0.006754f
C759 B.n643 VSUBS 0.006754f
C760 B.n644 VSUBS 0.006754f
C761 B.n645 VSUBS 0.006754f
C762 B.n646 VSUBS 0.006754f
C763 B.n647 VSUBS 0.006754f
C764 B.n648 VSUBS 0.006754f
C765 B.n649 VSUBS 0.006754f
C766 B.n650 VSUBS 0.006754f
C767 B.n651 VSUBS 0.006754f
C768 B.n652 VSUBS 0.006754f
C769 B.n653 VSUBS 0.006754f
C770 B.n654 VSUBS 0.006754f
C771 B.n655 VSUBS 0.006754f
C772 B.n656 VSUBS 0.006754f
C773 B.n657 VSUBS 0.006754f
C774 B.n658 VSUBS 0.006754f
C775 B.n659 VSUBS 0.006754f
C776 B.n660 VSUBS 0.006754f
C777 B.n661 VSUBS 0.014949f
C778 B.n662 VSUBS 0.014949f
C779 B.n663 VSUBS 0.01624f
C780 B.n664 VSUBS 0.006754f
C781 B.n665 VSUBS 0.006754f
C782 B.n666 VSUBS 0.006754f
C783 B.n667 VSUBS 0.006754f
C784 B.n668 VSUBS 0.006754f
C785 B.n669 VSUBS 0.006754f
C786 B.n670 VSUBS 0.006754f
C787 B.n671 VSUBS 0.006754f
C788 B.n672 VSUBS 0.006754f
C789 B.n673 VSUBS 0.006754f
C790 B.n674 VSUBS 0.006754f
C791 B.n675 VSUBS 0.006754f
C792 B.n676 VSUBS 0.006754f
C793 B.n677 VSUBS 0.006754f
C794 B.n678 VSUBS 0.006754f
C795 B.n679 VSUBS 0.006754f
C796 B.n680 VSUBS 0.006754f
C797 B.n681 VSUBS 0.006754f
C798 B.n682 VSUBS 0.006754f
C799 B.n683 VSUBS 0.006754f
C800 B.n684 VSUBS 0.006754f
C801 B.n685 VSUBS 0.006754f
C802 B.n686 VSUBS 0.006754f
C803 B.n687 VSUBS 0.006754f
C804 B.n688 VSUBS 0.006754f
C805 B.n689 VSUBS 0.006754f
C806 B.n690 VSUBS 0.006754f
C807 B.n691 VSUBS 0.006754f
C808 B.n692 VSUBS 0.006754f
C809 B.n693 VSUBS 0.006754f
C810 B.n694 VSUBS 0.006754f
C811 B.n695 VSUBS 0.006754f
C812 B.n696 VSUBS 0.006754f
C813 B.n697 VSUBS 0.006754f
C814 B.n698 VSUBS 0.006754f
C815 B.n699 VSUBS 0.006754f
C816 B.n700 VSUBS 0.006754f
C817 B.n701 VSUBS 0.006754f
C818 B.n702 VSUBS 0.006754f
C819 B.n703 VSUBS 0.006754f
C820 B.n704 VSUBS 0.006754f
C821 B.n705 VSUBS 0.006754f
C822 B.n706 VSUBS 0.006754f
C823 B.n707 VSUBS 0.006754f
C824 B.n708 VSUBS 0.006754f
C825 B.n709 VSUBS 0.006754f
C826 B.n710 VSUBS 0.006754f
C827 B.n711 VSUBS 0.006754f
C828 B.n712 VSUBS 0.006754f
C829 B.n713 VSUBS 0.006754f
C830 B.n714 VSUBS 0.006754f
C831 B.n715 VSUBS 0.006754f
C832 B.n716 VSUBS 0.006754f
C833 B.n717 VSUBS 0.006754f
C834 B.n718 VSUBS 0.006754f
C835 B.n719 VSUBS 0.006754f
C836 B.n720 VSUBS 0.006754f
C837 B.n721 VSUBS 0.006754f
C838 B.n722 VSUBS 0.006754f
C839 B.n723 VSUBS 0.006754f
C840 B.n724 VSUBS 0.006754f
C841 B.n725 VSUBS 0.006754f
C842 B.n726 VSUBS 0.006754f
C843 B.n727 VSUBS 0.006754f
C844 B.n728 VSUBS 0.006754f
C845 B.n729 VSUBS 0.006754f
C846 B.n730 VSUBS 0.006754f
C847 B.n731 VSUBS 0.006754f
C848 B.n732 VSUBS 0.006754f
C849 B.n733 VSUBS 0.006754f
C850 B.n734 VSUBS 0.006754f
C851 B.n735 VSUBS 0.006754f
C852 B.n736 VSUBS 0.006754f
C853 B.n737 VSUBS 0.006754f
C854 B.n738 VSUBS 0.006754f
C855 B.n739 VSUBS 0.006754f
C856 B.n740 VSUBS 0.006754f
C857 B.n741 VSUBS 0.006754f
C858 B.n742 VSUBS 0.006754f
C859 B.n743 VSUBS 0.006754f
C860 B.n744 VSUBS 0.006754f
C861 B.n745 VSUBS 0.006754f
C862 B.n746 VSUBS 0.006754f
C863 B.n747 VSUBS 0.006754f
C864 B.n748 VSUBS 0.006754f
C865 B.n749 VSUBS 0.006754f
C866 B.n750 VSUBS 0.006754f
C867 B.n751 VSUBS 0.006754f
C868 B.n752 VSUBS 0.006754f
C869 B.n753 VSUBS 0.006754f
C870 B.n754 VSUBS 0.006754f
C871 B.n755 VSUBS 0.006754f
C872 B.n756 VSUBS 0.006754f
C873 B.n757 VSUBS 0.004668f
C874 B.n758 VSUBS 0.006754f
C875 B.n759 VSUBS 0.006754f
C876 B.n760 VSUBS 0.005463f
C877 B.n761 VSUBS 0.006754f
C878 B.n762 VSUBS 0.006754f
C879 B.n763 VSUBS 0.006754f
C880 B.n764 VSUBS 0.006754f
C881 B.n765 VSUBS 0.006754f
C882 B.n766 VSUBS 0.006754f
C883 B.n767 VSUBS 0.006754f
C884 B.n768 VSUBS 0.006754f
C885 B.n769 VSUBS 0.006754f
C886 B.n770 VSUBS 0.006754f
C887 B.n771 VSUBS 0.006754f
C888 B.n772 VSUBS 0.005463f
C889 B.n773 VSUBS 0.015649f
C890 B.n774 VSUBS 0.004668f
C891 B.n775 VSUBS 0.006754f
C892 B.n776 VSUBS 0.006754f
C893 B.n777 VSUBS 0.006754f
C894 B.n778 VSUBS 0.006754f
C895 B.n779 VSUBS 0.006754f
C896 B.n780 VSUBS 0.006754f
C897 B.n781 VSUBS 0.006754f
C898 B.n782 VSUBS 0.006754f
C899 B.n783 VSUBS 0.006754f
C900 B.n784 VSUBS 0.006754f
C901 B.n785 VSUBS 0.006754f
C902 B.n786 VSUBS 0.006754f
C903 B.n787 VSUBS 0.006754f
C904 B.n788 VSUBS 0.006754f
C905 B.n789 VSUBS 0.006754f
C906 B.n790 VSUBS 0.006754f
C907 B.n791 VSUBS 0.006754f
C908 B.n792 VSUBS 0.006754f
C909 B.n793 VSUBS 0.006754f
C910 B.n794 VSUBS 0.006754f
C911 B.n795 VSUBS 0.006754f
C912 B.n796 VSUBS 0.006754f
C913 B.n797 VSUBS 0.006754f
C914 B.n798 VSUBS 0.006754f
C915 B.n799 VSUBS 0.006754f
C916 B.n800 VSUBS 0.006754f
C917 B.n801 VSUBS 0.006754f
C918 B.n802 VSUBS 0.006754f
C919 B.n803 VSUBS 0.006754f
C920 B.n804 VSUBS 0.006754f
C921 B.n805 VSUBS 0.006754f
C922 B.n806 VSUBS 0.006754f
C923 B.n807 VSUBS 0.006754f
C924 B.n808 VSUBS 0.006754f
C925 B.n809 VSUBS 0.006754f
C926 B.n810 VSUBS 0.006754f
C927 B.n811 VSUBS 0.006754f
C928 B.n812 VSUBS 0.006754f
C929 B.n813 VSUBS 0.006754f
C930 B.n814 VSUBS 0.006754f
C931 B.n815 VSUBS 0.006754f
C932 B.n816 VSUBS 0.006754f
C933 B.n817 VSUBS 0.006754f
C934 B.n818 VSUBS 0.006754f
C935 B.n819 VSUBS 0.006754f
C936 B.n820 VSUBS 0.006754f
C937 B.n821 VSUBS 0.006754f
C938 B.n822 VSUBS 0.006754f
C939 B.n823 VSUBS 0.006754f
C940 B.n824 VSUBS 0.006754f
C941 B.n825 VSUBS 0.006754f
C942 B.n826 VSUBS 0.006754f
C943 B.n827 VSUBS 0.006754f
C944 B.n828 VSUBS 0.006754f
C945 B.n829 VSUBS 0.006754f
C946 B.n830 VSUBS 0.006754f
C947 B.n831 VSUBS 0.006754f
C948 B.n832 VSUBS 0.006754f
C949 B.n833 VSUBS 0.006754f
C950 B.n834 VSUBS 0.006754f
C951 B.n835 VSUBS 0.006754f
C952 B.n836 VSUBS 0.006754f
C953 B.n837 VSUBS 0.006754f
C954 B.n838 VSUBS 0.006754f
C955 B.n839 VSUBS 0.006754f
C956 B.n840 VSUBS 0.006754f
C957 B.n841 VSUBS 0.006754f
C958 B.n842 VSUBS 0.006754f
C959 B.n843 VSUBS 0.006754f
C960 B.n844 VSUBS 0.006754f
C961 B.n845 VSUBS 0.006754f
C962 B.n846 VSUBS 0.006754f
C963 B.n847 VSUBS 0.006754f
C964 B.n848 VSUBS 0.006754f
C965 B.n849 VSUBS 0.006754f
C966 B.n850 VSUBS 0.006754f
C967 B.n851 VSUBS 0.006754f
C968 B.n852 VSUBS 0.006754f
C969 B.n853 VSUBS 0.006754f
C970 B.n854 VSUBS 0.006754f
C971 B.n855 VSUBS 0.006754f
C972 B.n856 VSUBS 0.006754f
C973 B.n857 VSUBS 0.006754f
C974 B.n858 VSUBS 0.006754f
C975 B.n859 VSUBS 0.006754f
C976 B.n860 VSUBS 0.006754f
C977 B.n861 VSUBS 0.006754f
C978 B.n862 VSUBS 0.006754f
C979 B.n863 VSUBS 0.006754f
C980 B.n864 VSUBS 0.006754f
C981 B.n865 VSUBS 0.006754f
C982 B.n866 VSUBS 0.006754f
C983 B.n867 VSUBS 0.006754f
C984 B.n868 VSUBS 0.01624f
C985 B.n869 VSUBS 0.01624f
C986 B.n870 VSUBS 0.014949f
C987 B.n871 VSUBS 0.006754f
C988 B.n872 VSUBS 0.006754f
C989 B.n873 VSUBS 0.006754f
C990 B.n874 VSUBS 0.006754f
C991 B.n875 VSUBS 0.006754f
C992 B.n876 VSUBS 0.006754f
C993 B.n877 VSUBS 0.006754f
C994 B.n878 VSUBS 0.006754f
C995 B.n879 VSUBS 0.006754f
C996 B.n880 VSUBS 0.006754f
C997 B.n881 VSUBS 0.006754f
C998 B.n882 VSUBS 0.006754f
C999 B.n883 VSUBS 0.006754f
C1000 B.n884 VSUBS 0.006754f
C1001 B.n885 VSUBS 0.006754f
C1002 B.n886 VSUBS 0.006754f
C1003 B.n887 VSUBS 0.006754f
C1004 B.n888 VSUBS 0.006754f
C1005 B.n889 VSUBS 0.006754f
C1006 B.n890 VSUBS 0.006754f
C1007 B.n891 VSUBS 0.006754f
C1008 B.n892 VSUBS 0.006754f
C1009 B.n893 VSUBS 0.006754f
C1010 B.n894 VSUBS 0.006754f
C1011 B.n895 VSUBS 0.006754f
C1012 B.n896 VSUBS 0.006754f
C1013 B.n897 VSUBS 0.006754f
C1014 B.n898 VSUBS 0.006754f
C1015 B.n899 VSUBS 0.006754f
C1016 B.n900 VSUBS 0.006754f
C1017 B.n901 VSUBS 0.006754f
C1018 B.n902 VSUBS 0.006754f
C1019 B.n903 VSUBS 0.006754f
C1020 B.n904 VSUBS 0.006754f
C1021 B.n905 VSUBS 0.006754f
C1022 B.n906 VSUBS 0.006754f
C1023 B.n907 VSUBS 0.006754f
C1024 B.n908 VSUBS 0.006754f
C1025 B.n909 VSUBS 0.006754f
C1026 B.n910 VSUBS 0.006754f
C1027 B.n911 VSUBS 0.006754f
C1028 B.n912 VSUBS 0.006754f
C1029 B.n913 VSUBS 0.006754f
C1030 B.n914 VSUBS 0.006754f
C1031 B.n915 VSUBS 0.006754f
C1032 B.n916 VSUBS 0.006754f
C1033 B.n917 VSUBS 0.006754f
C1034 B.n918 VSUBS 0.006754f
C1035 B.n919 VSUBS 0.006754f
C1036 B.n920 VSUBS 0.006754f
C1037 B.n921 VSUBS 0.006754f
C1038 B.n922 VSUBS 0.006754f
C1039 B.n923 VSUBS 0.006754f
C1040 B.n924 VSUBS 0.006754f
C1041 B.n925 VSUBS 0.006754f
C1042 B.n926 VSUBS 0.006754f
C1043 B.n927 VSUBS 0.006754f
C1044 B.n928 VSUBS 0.006754f
C1045 B.n929 VSUBS 0.006754f
C1046 B.n930 VSUBS 0.006754f
C1047 B.n931 VSUBS 0.006754f
C1048 B.n932 VSUBS 0.006754f
C1049 B.n933 VSUBS 0.006754f
C1050 B.n934 VSUBS 0.006754f
C1051 B.n935 VSUBS 0.006754f
C1052 B.n936 VSUBS 0.006754f
C1053 B.n937 VSUBS 0.006754f
C1054 B.n938 VSUBS 0.006754f
C1055 B.n939 VSUBS 0.008814f
C1056 B.n940 VSUBS 0.009389f
C1057 B.n941 VSUBS 0.018672f
C1058 VDD1.t1 VSUBS 0.411033f
C1059 VDD1.t7 VSUBS 0.411033f
C1060 VDD1.n0 VSUBS 3.47911f
C1061 VDD1.t3 VSUBS 0.411033f
C1062 VDD1.t4 VSUBS 0.411033f
C1063 VDD1.n1 VSUBS 3.47766f
C1064 VDD1.t0 VSUBS 0.411033f
C1065 VDD1.t2 VSUBS 0.411033f
C1066 VDD1.n2 VSUBS 3.47766f
C1067 VDD1.n3 VSUBS 4.49925f
C1068 VDD1.t6 VSUBS 0.411033f
C1069 VDD1.t5 VSUBS 0.411033f
C1070 VDD1.n4 VSUBS 3.46494f
C1071 VDD1.n5 VSUBS 3.99747f
C1072 VTAIL.t6 VSUBS 0.3568f
C1073 VTAIL.t5 VSUBS 0.3568f
C1074 VTAIL.n0 VSUBS 2.86997f
C1075 VTAIL.n1 VSUBS 0.730467f
C1076 VTAIL.n2 VSUBS 0.024637f
C1077 VTAIL.n3 VSUBS 0.023226f
C1078 VTAIL.n4 VSUBS 0.012481f
C1079 VTAIL.n5 VSUBS 0.0295f
C1080 VTAIL.n6 VSUBS 0.013215f
C1081 VTAIL.n7 VSUBS 0.023226f
C1082 VTAIL.n8 VSUBS 0.012481f
C1083 VTAIL.n9 VSUBS 0.0295f
C1084 VTAIL.n10 VSUBS 0.013215f
C1085 VTAIL.n11 VSUBS 0.023226f
C1086 VTAIL.n12 VSUBS 0.012481f
C1087 VTAIL.n13 VSUBS 0.0295f
C1088 VTAIL.n14 VSUBS 0.013215f
C1089 VTAIL.n15 VSUBS 0.023226f
C1090 VTAIL.n16 VSUBS 0.012481f
C1091 VTAIL.n17 VSUBS 0.0295f
C1092 VTAIL.n18 VSUBS 0.013215f
C1093 VTAIL.n19 VSUBS 0.023226f
C1094 VTAIL.n20 VSUBS 0.012481f
C1095 VTAIL.n21 VSUBS 0.0295f
C1096 VTAIL.n22 VSUBS 0.013215f
C1097 VTAIL.n23 VSUBS 0.023226f
C1098 VTAIL.n24 VSUBS 0.012481f
C1099 VTAIL.n25 VSUBS 0.0295f
C1100 VTAIL.n26 VSUBS 0.013215f
C1101 VTAIL.n27 VSUBS 0.023226f
C1102 VTAIL.n28 VSUBS 0.012481f
C1103 VTAIL.n29 VSUBS 0.0295f
C1104 VTAIL.n30 VSUBS 0.013215f
C1105 VTAIL.n31 VSUBS 0.023226f
C1106 VTAIL.n32 VSUBS 0.012481f
C1107 VTAIL.n33 VSUBS 0.0295f
C1108 VTAIL.n34 VSUBS 0.013215f
C1109 VTAIL.n35 VSUBS 0.261052f
C1110 VTAIL.t7 VSUBS 0.064153f
C1111 VTAIL.n36 VSUBS 0.022125f
C1112 VTAIL.n37 VSUBS 0.022191f
C1113 VTAIL.n38 VSUBS 0.012481f
C1114 VTAIL.n39 VSUBS 1.89832f
C1115 VTAIL.n40 VSUBS 0.023226f
C1116 VTAIL.n41 VSUBS 0.012481f
C1117 VTAIL.n42 VSUBS 0.013215f
C1118 VTAIL.n43 VSUBS 0.0295f
C1119 VTAIL.n44 VSUBS 0.0295f
C1120 VTAIL.n45 VSUBS 0.013215f
C1121 VTAIL.n46 VSUBS 0.012481f
C1122 VTAIL.n47 VSUBS 0.023226f
C1123 VTAIL.n48 VSUBS 0.023226f
C1124 VTAIL.n49 VSUBS 0.012481f
C1125 VTAIL.n50 VSUBS 0.013215f
C1126 VTAIL.n51 VSUBS 0.0295f
C1127 VTAIL.n52 VSUBS 0.0295f
C1128 VTAIL.n53 VSUBS 0.0295f
C1129 VTAIL.n54 VSUBS 0.013215f
C1130 VTAIL.n55 VSUBS 0.012481f
C1131 VTAIL.n56 VSUBS 0.023226f
C1132 VTAIL.n57 VSUBS 0.023226f
C1133 VTAIL.n58 VSUBS 0.012481f
C1134 VTAIL.n59 VSUBS 0.012848f
C1135 VTAIL.n60 VSUBS 0.012848f
C1136 VTAIL.n61 VSUBS 0.0295f
C1137 VTAIL.n62 VSUBS 0.0295f
C1138 VTAIL.n63 VSUBS 0.013215f
C1139 VTAIL.n64 VSUBS 0.012481f
C1140 VTAIL.n65 VSUBS 0.023226f
C1141 VTAIL.n66 VSUBS 0.023226f
C1142 VTAIL.n67 VSUBS 0.012481f
C1143 VTAIL.n68 VSUBS 0.013215f
C1144 VTAIL.n69 VSUBS 0.0295f
C1145 VTAIL.n70 VSUBS 0.0295f
C1146 VTAIL.n71 VSUBS 0.013215f
C1147 VTAIL.n72 VSUBS 0.012481f
C1148 VTAIL.n73 VSUBS 0.023226f
C1149 VTAIL.n74 VSUBS 0.023226f
C1150 VTAIL.n75 VSUBS 0.012481f
C1151 VTAIL.n76 VSUBS 0.013215f
C1152 VTAIL.n77 VSUBS 0.0295f
C1153 VTAIL.n78 VSUBS 0.0295f
C1154 VTAIL.n79 VSUBS 0.013215f
C1155 VTAIL.n80 VSUBS 0.012481f
C1156 VTAIL.n81 VSUBS 0.023226f
C1157 VTAIL.n82 VSUBS 0.023226f
C1158 VTAIL.n83 VSUBS 0.012481f
C1159 VTAIL.n84 VSUBS 0.013215f
C1160 VTAIL.n85 VSUBS 0.0295f
C1161 VTAIL.n86 VSUBS 0.0295f
C1162 VTAIL.n87 VSUBS 0.013215f
C1163 VTAIL.n88 VSUBS 0.012481f
C1164 VTAIL.n89 VSUBS 0.023226f
C1165 VTAIL.n90 VSUBS 0.023226f
C1166 VTAIL.n91 VSUBS 0.012481f
C1167 VTAIL.n92 VSUBS 0.013215f
C1168 VTAIL.n93 VSUBS 0.0295f
C1169 VTAIL.n94 VSUBS 0.0295f
C1170 VTAIL.n95 VSUBS 0.013215f
C1171 VTAIL.n96 VSUBS 0.012481f
C1172 VTAIL.n97 VSUBS 0.023226f
C1173 VTAIL.n98 VSUBS 0.023226f
C1174 VTAIL.n99 VSUBS 0.012481f
C1175 VTAIL.n100 VSUBS 0.013215f
C1176 VTAIL.n101 VSUBS 0.0295f
C1177 VTAIL.n102 VSUBS 0.072576f
C1178 VTAIL.n103 VSUBS 0.013215f
C1179 VTAIL.n104 VSUBS 0.024509f
C1180 VTAIL.n105 VSUBS 0.057493f
C1181 VTAIL.n106 VSUBS 0.055216f
C1182 VTAIL.n107 VSUBS 0.230701f
C1183 VTAIL.n108 VSUBS 0.024637f
C1184 VTAIL.n109 VSUBS 0.023226f
C1185 VTAIL.n110 VSUBS 0.012481f
C1186 VTAIL.n111 VSUBS 0.0295f
C1187 VTAIL.n112 VSUBS 0.013215f
C1188 VTAIL.n113 VSUBS 0.023226f
C1189 VTAIL.n114 VSUBS 0.012481f
C1190 VTAIL.n115 VSUBS 0.0295f
C1191 VTAIL.n116 VSUBS 0.013215f
C1192 VTAIL.n117 VSUBS 0.023226f
C1193 VTAIL.n118 VSUBS 0.012481f
C1194 VTAIL.n119 VSUBS 0.0295f
C1195 VTAIL.n120 VSUBS 0.013215f
C1196 VTAIL.n121 VSUBS 0.023226f
C1197 VTAIL.n122 VSUBS 0.012481f
C1198 VTAIL.n123 VSUBS 0.0295f
C1199 VTAIL.n124 VSUBS 0.013215f
C1200 VTAIL.n125 VSUBS 0.023226f
C1201 VTAIL.n126 VSUBS 0.012481f
C1202 VTAIL.n127 VSUBS 0.0295f
C1203 VTAIL.n128 VSUBS 0.013215f
C1204 VTAIL.n129 VSUBS 0.023226f
C1205 VTAIL.n130 VSUBS 0.012481f
C1206 VTAIL.n131 VSUBS 0.0295f
C1207 VTAIL.n132 VSUBS 0.013215f
C1208 VTAIL.n133 VSUBS 0.023226f
C1209 VTAIL.n134 VSUBS 0.012481f
C1210 VTAIL.n135 VSUBS 0.0295f
C1211 VTAIL.n136 VSUBS 0.013215f
C1212 VTAIL.n137 VSUBS 0.023226f
C1213 VTAIL.n138 VSUBS 0.012481f
C1214 VTAIL.n139 VSUBS 0.0295f
C1215 VTAIL.n140 VSUBS 0.013215f
C1216 VTAIL.n141 VSUBS 0.261052f
C1217 VTAIL.t11 VSUBS 0.064153f
C1218 VTAIL.n142 VSUBS 0.022125f
C1219 VTAIL.n143 VSUBS 0.022191f
C1220 VTAIL.n144 VSUBS 0.012481f
C1221 VTAIL.n145 VSUBS 1.89832f
C1222 VTAIL.n146 VSUBS 0.023226f
C1223 VTAIL.n147 VSUBS 0.012481f
C1224 VTAIL.n148 VSUBS 0.013215f
C1225 VTAIL.n149 VSUBS 0.0295f
C1226 VTAIL.n150 VSUBS 0.0295f
C1227 VTAIL.n151 VSUBS 0.013215f
C1228 VTAIL.n152 VSUBS 0.012481f
C1229 VTAIL.n153 VSUBS 0.023226f
C1230 VTAIL.n154 VSUBS 0.023226f
C1231 VTAIL.n155 VSUBS 0.012481f
C1232 VTAIL.n156 VSUBS 0.013215f
C1233 VTAIL.n157 VSUBS 0.0295f
C1234 VTAIL.n158 VSUBS 0.0295f
C1235 VTAIL.n159 VSUBS 0.0295f
C1236 VTAIL.n160 VSUBS 0.013215f
C1237 VTAIL.n161 VSUBS 0.012481f
C1238 VTAIL.n162 VSUBS 0.023226f
C1239 VTAIL.n163 VSUBS 0.023226f
C1240 VTAIL.n164 VSUBS 0.012481f
C1241 VTAIL.n165 VSUBS 0.012848f
C1242 VTAIL.n166 VSUBS 0.012848f
C1243 VTAIL.n167 VSUBS 0.0295f
C1244 VTAIL.n168 VSUBS 0.0295f
C1245 VTAIL.n169 VSUBS 0.013215f
C1246 VTAIL.n170 VSUBS 0.012481f
C1247 VTAIL.n171 VSUBS 0.023226f
C1248 VTAIL.n172 VSUBS 0.023226f
C1249 VTAIL.n173 VSUBS 0.012481f
C1250 VTAIL.n174 VSUBS 0.013215f
C1251 VTAIL.n175 VSUBS 0.0295f
C1252 VTAIL.n176 VSUBS 0.0295f
C1253 VTAIL.n177 VSUBS 0.013215f
C1254 VTAIL.n178 VSUBS 0.012481f
C1255 VTAIL.n179 VSUBS 0.023226f
C1256 VTAIL.n180 VSUBS 0.023226f
C1257 VTAIL.n181 VSUBS 0.012481f
C1258 VTAIL.n182 VSUBS 0.013215f
C1259 VTAIL.n183 VSUBS 0.0295f
C1260 VTAIL.n184 VSUBS 0.0295f
C1261 VTAIL.n185 VSUBS 0.013215f
C1262 VTAIL.n186 VSUBS 0.012481f
C1263 VTAIL.n187 VSUBS 0.023226f
C1264 VTAIL.n188 VSUBS 0.023226f
C1265 VTAIL.n189 VSUBS 0.012481f
C1266 VTAIL.n190 VSUBS 0.013215f
C1267 VTAIL.n191 VSUBS 0.0295f
C1268 VTAIL.n192 VSUBS 0.0295f
C1269 VTAIL.n193 VSUBS 0.013215f
C1270 VTAIL.n194 VSUBS 0.012481f
C1271 VTAIL.n195 VSUBS 0.023226f
C1272 VTAIL.n196 VSUBS 0.023226f
C1273 VTAIL.n197 VSUBS 0.012481f
C1274 VTAIL.n198 VSUBS 0.013215f
C1275 VTAIL.n199 VSUBS 0.0295f
C1276 VTAIL.n200 VSUBS 0.0295f
C1277 VTAIL.n201 VSUBS 0.013215f
C1278 VTAIL.n202 VSUBS 0.012481f
C1279 VTAIL.n203 VSUBS 0.023226f
C1280 VTAIL.n204 VSUBS 0.023226f
C1281 VTAIL.n205 VSUBS 0.012481f
C1282 VTAIL.n206 VSUBS 0.013215f
C1283 VTAIL.n207 VSUBS 0.0295f
C1284 VTAIL.n208 VSUBS 0.072576f
C1285 VTAIL.n209 VSUBS 0.013215f
C1286 VTAIL.n210 VSUBS 0.024509f
C1287 VTAIL.n211 VSUBS 0.057493f
C1288 VTAIL.n212 VSUBS 0.055216f
C1289 VTAIL.n213 VSUBS 0.230701f
C1290 VTAIL.t13 VSUBS 0.3568f
C1291 VTAIL.t15 VSUBS 0.3568f
C1292 VTAIL.n214 VSUBS 2.86997f
C1293 VTAIL.n215 VSUBS 0.899662f
C1294 VTAIL.n216 VSUBS 0.024637f
C1295 VTAIL.n217 VSUBS 0.023226f
C1296 VTAIL.n218 VSUBS 0.012481f
C1297 VTAIL.n219 VSUBS 0.0295f
C1298 VTAIL.n220 VSUBS 0.013215f
C1299 VTAIL.n221 VSUBS 0.023226f
C1300 VTAIL.n222 VSUBS 0.012481f
C1301 VTAIL.n223 VSUBS 0.0295f
C1302 VTAIL.n224 VSUBS 0.013215f
C1303 VTAIL.n225 VSUBS 0.023226f
C1304 VTAIL.n226 VSUBS 0.012481f
C1305 VTAIL.n227 VSUBS 0.0295f
C1306 VTAIL.n228 VSUBS 0.013215f
C1307 VTAIL.n229 VSUBS 0.023226f
C1308 VTAIL.n230 VSUBS 0.012481f
C1309 VTAIL.n231 VSUBS 0.0295f
C1310 VTAIL.n232 VSUBS 0.013215f
C1311 VTAIL.n233 VSUBS 0.023226f
C1312 VTAIL.n234 VSUBS 0.012481f
C1313 VTAIL.n235 VSUBS 0.0295f
C1314 VTAIL.n236 VSUBS 0.013215f
C1315 VTAIL.n237 VSUBS 0.023226f
C1316 VTAIL.n238 VSUBS 0.012481f
C1317 VTAIL.n239 VSUBS 0.0295f
C1318 VTAIL.n240 VSUBS 0.013215f
C1319 VTAIL.n241 VSUBS 0.023226f
C1320 VTAIL.n242 VSUBS 0.012481f
C1321 VTAIL.n243 VSUBS 0.0295f
C1322 VTAIL.n244 VSUBS 0.013215f
C1323 VTAIL.n245 VSUBS 0.023226f
C1324 VTAIL.n246 VSUBS 0.012481f
C1325 VTAIL.n247 VSUBS 0.0295f
C1326 VTAIL.n248 VSUBS 0.013215f
C1327 VTAIL.n249 VSUBS 0.261052f
C1328 VTAIL.t14 VSUBS 0.064153f
C1329 VTAIL.n250 VSUBS 0.022125f
C1330 VTAIL.n251 VSUBS 0.022191f
C1331 VTAIL.n252 VSUBS 0.012481f
C1332 VTAIL.n253 VSUBS 1.89832f
C1333 VTAIL.n254 VSUBS 0.023226f
C1334 VTAIL.n255 VSUBS 0.012481f
C1335 VTAIL.n256 VSUBS 0.013215f
C1336 VTAIL.n257 VSUBS 0.0295f
C1337 VTAIL.n258 VSUBS 0.0295f
C1338 VTAIL.n259 VSUBS 0.013215f
C1339 VTAIL.n260 VSUBS 0.012481f
C1340 VTAIL.n261 VSUBS 0.023226f
C1341 VTAIL.n262 VSUBS 0.023226f
C1342 VTAIL.n263 VSUBS 0.012481f
C1343 VTAIL.n264 VSUBS 0.013215f
C1344 VTAIL.n265 VSUBS 0.0295f
C1345 VTAIL.n266 VSUBS 0.0295f
C1346 VTAIL.n267 VSUBS 0.0295f
C1347 VTAIL.n268 VSUBS 0.013215f
C1348 VTAIL.n269 VSUBS 0.012481f
C1349 VTAIL.n270 VSUBS 0.023226f
C1350 VTAIL.n271 VSUBS 0.023226f
C1351 VTAIL.n272 VSUBS 0.012481f
C1352 VTAIL.n273 VSUBS 0.012848f
C1353 VTAIL.n274 VSUBS 0.012848f
C1354 VTAIL.n275 VSUBS 0.0295f
C1355 VTAIL.n276 VSUBS 0.0295f
C1356 VTAIL.n277 VSUBS 0.013215f
C1357 VTAIL.n278 VSUBS 0.012481f
C1358 VTAIL.n279 VSUBS 0.023226f
C1359 VTAIL.n280 VSUBS 0.023226f
C1360 VTAIL.n281 VSUBS 0.012481f
C1361 VTAIL.n282 VSUBS 0.013215f
C1362 VTAIL.n283 VSUBS 0.0295f
C1363 VTAIL.n284 VSUBS 0.0295f
C1364 VTAIL.n285 VSUBS 0.013215f
C1365 VTAIL.n286 VSUBS 0.012481f
C1366 VTAIL.n287 VSUBS 0.023226f
C1367 VTAIL.n288 VSUBS 0.023226f
C1368 VTAIL.n289 VSUBS 0.012481f
C1369 VTAIL.n290 VSUBS 0.013215f
C1370 VTAIL.n291 VSUBS 0.0295f
C1371 VTAIL.n292 VSUBS 0.0295f
C1372 VTAIL.n293 VSUBS 0.013215f
C1373 VTAIL.n294 VSUBS 0.012481f
C1374 VTAIL.n295 VSUBS 0.023226f
C1375 VTAIL.n296 VSUBS 0.023226f
C1376 VTAIL.n297 VSUBS 0.012481f
C1377 VTAIL.n298 VSUBS 0.013215f
C1378 VTAIL.n299 VSUBS 0.0295f
C1379 VTAIL.n300 VSUBS 0.0295f
C1380 VTAIL.n301 VSUBS 0.013215f
C1381 VTAIL.n302 VSUBS 0.012481f
C1382 VTAIL.n303 VSUBS 0.023226f
C1383 VTAIL.n304 VSUBS 0.023226f
C1384 VTAIL.n305 VSUBS 0.012481f
C1385 VTAIL.n306 VSUBS 0.013215f
C1386 VTAIL.n307 VSUBS 0.0295f
C1387 VTAIL.n308 VSUBS 0.0295f
C1388 VTAIL.n309 VSUBS 0.013215f
C1389 VTAIL.n310 VSUBS 0.012481f
C1390 VTAIL.n311 VSUBS 0.023226f
C1391 VTAIL.n312 VSUBS 0.023226f
C1392 VTAIL.n313 VSUBS 0.012481f
C1393 VTAIL.n314 VSUBS 0.013215f
C1394 VTAIL.n315 VSUBS 0.0295f
C1395 VTAIL.n316 VSUBS 0.072576f
C1396 VTAIL.n317 VSUBS 0.013215f
C1397 VTAIL.n318 VSUBS 0.024509f
C1398 VTAIL.n319 VSUBS 0.057493f
C1399 VTAIL.n320 VSUBS 0.055216f
C1400 VTAIL.n321 VSUBS 1.93879f
C1401 VTAIL.n322 VSUBS 0.024637f
C1402 VTAIL.n323 VSUBS 0.023226f
C1403 VTAIL.n324 VSUBS 0.012481f
C1404 VTAIL.n325 VSUBS 0.0295f
C1405 VTAIL.n326 VSUBS 0.013215f
C1406 VTAIL.n327 VSUBS 0.023226f
C1407 VTAIL.n328 VSUBS 0.012481f
C1408 VTAIL.n329 VSUBS 0.0295f
C1409 VTAIL.n330 VSUBS 0.013215f
C1410 VTAIL.n331 VSUBS 0.023226f
C1411 VTAIL.n332 VSUBS 0.012481f
C1412 VTAIL.n333 VSUBS 0.0295f
C1413 VTAIL.n334 VSUBS 0.013215f
C1414 VTAIL.n335 VSUBS 0.023226f
C1415 VTAIL.n336 VSUBS 0.012481f
C1416 VTAIL.n337 VSUBS 0.0295f
C1417 VTAIL.n338 VSUBS 0.013215f
C1418 VTAIL.n339 VSUBS 0.023226f
C1419 VTAIL.n340 VSUBS 0.012481f
C1420 VTAIL.n341 VSUBS 0.0295f
C1421 VTAIL.n342 VSUBS 0.013215f
C1422 VTAIL.n343 VSUBS 0.023226f
C1423 VTAIL.n344 VSUBS 0.012481f
C1424 VTAIL.n345 VSUBS 0.0295f
C1425 VTAIL.n346 VSUBS 0.013215f
C1426 VTAIL.n347 VSUBS 0.023226f
C1427 VTAIL.n348 VSUBS 0.012481f
C1428 VTAIL.n349 VSUBS 0.0295f
C1429 VTAIL.n350 VSUBS 0.0295f
C1430 VTAIL.n351 VSUBS 0.013215f
C1431 VTAIL.n352 VSUBS 0.023226f
C1432 VTAIL.n353 VSUBS 0.012481f
C1433 VTAIL.n354 VSUBS 0.0295f
C1434 VTAIL.n355 VSUBS 0.013215f
C1435 VTAIL.n356 VSUBS 0.261052f
C1436 VTAIL.t1 VSUBS 0.064153f
C1437 VTAIL.n357 VSUBS 0.022125f
C1438 VTAIL.n358 VSUBS 0.022191f
C1439 VTAIL.n359 VSUBS 0.012481f
C1440 VTAIL.n360 VSUBS 1.89832f
C1441 VTAIL.n361 VSUBS 0.023226f
C1442 VTAIL.n362 VSUBS 0.012481f
C1443 VTAIL.n363 VSUBS 0.013215f
C1444 VTAIL.n364 VSUBS 0.0295f
C1445 VTAIL.n365 VSUBS 0.0295f
C1446 VTAIL.n366 VSUBS 0.013215f
C1447 VTAIL.n367 VSUBS 0.012481f
C1448 VTAIL.n368 VSUBS 0.023226f
C1449 VTAIL.n369 VSUBS 0.023226f
C1450 VTAIL.n370 VSUBS 0.012481f
C1451 VTAIL.n371 VSUBS 0.013215f
C1452 VTAIL.n372 VSUBS 0.0295f
C1453 VTAIL.n373 VSUBS 0.0295f
C1454 VTAIL.n374 VSUBS 0.013215f
C1455 VTAIL.n375 VSUBS 0.012481f
C1456 VTAIL.n376 VSUBS 0.023226f
C1457 VTAIL.n377 VSUBS 0.023226f
C1458 VTAIL.n378 VSUBS 0.012481f
C1459 VTAIL.n379 VSUBS 0.012848f
C1460 VTAIL.n380 VSUBS 0.012848f
C1461 VTAIL.n381 VSUBS 0.0295f
C1462 VTAIL.n382 VSUBS 0.0295f
C1463 VTAIL.n383 VSUBS 0.013215f
C1464 VTAIL.n384 VSUBS 0.012481f
C1465 VTAIL.n385 VSUBS 0.023226f
C1466 VTAIL.n386 VSUBS 0.023226f
C1467 VTAIL.n387 VSUBS 0.012481f
C1468 VTAIL.n388 VSUBS 0.013215f
C1469 VTAIL.n389 VSUBS 0.0295f
C1470 VTAIL.n390 VSUBS 0.0295f
C1471 VTAIL.n391 VSUBS 0.013215f
C1472 VTAIL.n392 VSUBS 0.012481f
C1473 VTAIL.n393 VSUBS 0.023226f
C1474 VTAIL.n394 VSUBS 0.023226f
C1475 VTAIL.n395 VSUBS 0.012481f
C1476 VTAIL.n396 VSUBS 0.013215f
C1477 VTAIL.n397 VSUBS 0.0295f
C1478 VTAIL.n398 VSUBS 0.0295f
C1479 VTAIL.n399 VSUBS 0.013215f
C1480 VTAIL.n400 VSUBS 0.012481f
C1481 VTAIL.n401 VSUBS 0.023226f
C1482 VTAIL.n402 VSUBS 0.023226f
C1483 VTAIL.n403 VSUBS 0.012481f
C1484 VTAIL.n404 VSUBS 0.013215f
C1485 VTAIL.n405 VSUBS 0.0295f
C1486 VTAIL.n406 VSUBS 0.0295f
C1487 VTAIL.n407 VSUBS 0.013215f
C1488 VTAIL.n408 VSUBS 0.012481f
C1489 VTAIL.n409 VSUBS 0.023226f
C1490 VTAIL.n410 VSUBS 0.023226f
C1491 VTAIL.n411 VSUBS 0.012481f
C1492 VTAIL.n412 VSUBS 0.013215f
C1493 VTAIL.n413 VSUBS 0.0295f
C1494 VTAIL.n414 VSUBS 0.0295f
C1495 VTAIL.n415 VSUBS 0.013215f
C1496 VTAIL.n416 VSUBS 0.012481f
C1497 VTAIL.n417 VSUBS 0.023226f
C1498 VTAIL.n418 VSUBS 0.023226f
C1499 VTAIL.n419 VSUBS 0.012481f
C1500 VTAIL.n420 VSUBS 0.013215f
C1501 VTAIL.n421 VSUBS 0.0295f
C1502 VTAIL.n422 VSUBS 0.072576f
C1503 VTAIL.n423 VSUBS 0.013215f
C1504 VTAIL.n424 VSUBS 0.024509f
C1505 VTAIL.n425 VSUBS 0.057493f
C1506 VTAIL.n426 VSUBS 0.055216f
C1507 VTAIL.n427 VSUBS 1.93879f
C1508 VTAIL.t2 VSUBS 0.3568f
C1509 VTAIL.t3 VSUBS 0.3568f
C1510 VTAIL.n428 VSUBS 2.86999f
C1511 VTAIL.n429 VSUBS 0.899645f
C1512 VTAIL.n430 VSUBS 0.024637f
C1513 VTAIL.n431 VSUBS 0.023226f
C1514 VTAIL.n432 VSUBS 0.012481f
C1515 VTAIL.n433 VSUBS 0.0295f
C1516 VTAIL.n434 VSUBS 0.013215f
C1517 VTAIL.n435 VSUBS 0.023226f
C1518 VTAIL.n436 VSUBS 0.012481f
C1519 VTAIL.n437 VSUBS 0.0295f
C1520 VTAIL.n438 VSUBS 0.013215f
C1521 VTAIL.n439 VSUBS 0.023226f
C1522 VTAIL.n440 VSUBS 0.012481f
C1523 VTAIL.n441 VSUBS 0.0295f
C1524 VTAIL.n442 VSUBS 0.013215f
C1525 VTAIL.n443 VSUBS 0.023226f
C1526 VTAIL.n444 VSUBS 0.012481f
C1527 VTAIL.n445 VSUBS 0.0295f
C1528 VTAIL.n446 VSUBS 0.013215f
C1529 VTAIL.n447 VSUBS 0.023226f
C1530 VTAIL.n448 VSUBS 0.012481f
C1531 VTAIL.n449 VSUBS 0.0295f
C1532 VTAIL.n450 VSUBS 0.013215f
C1533 VTAIL.n451 VSUBS 0.023226f
C1534 VTAIL.n452 VSUBS 0.012481f
C1535 VTAIL.n453 VSUBS 0.0295f
C1536 VTAIL.n454 VSUBS 0.013215f
C1537 VTAIL.n455 VSUBS 0.023226f
C1538 VTAIL.n456 VSUBS 0.012481f
C1539 VTAIL.n457 VSUBS 0.0295f
C1540 VTAIL.n458 VSUBS 0.0295f
C1541 VTAIL.n459 VSUBS 0.013215f
C1542 VTAIL.n460 VSUBS 0.023226f
C1543 VTAIL.n461 VSUBS 0.012481f
C1544 VTAIL.n462 VSUBS 0.0295f
C1545 VTAIL.n463 VSUBS 0.013215f
C1546 VTAIL.n464 VSUBS 0.261052f
C1547 VTAIL.t0 VSUBS 0.064153f
C1548 VTAIL.n465 VSUBS 0.022125f
C1549 VTAIL.n466 VSUBS 0.022191f
C1550 VTAIL.n467 VSUBS 0.012481f
C1551 VTAIL.n468 VSUBS 1.89832f
C1552 VTAIL.n469 VSUBS 0.023226f
C1553 VTAIL.n470 VSUBS 0.012481f
C1554 VTAIL.n471 VSUBS 0.013215f
C1555 VTAIL.n472 VSUBS 0.0295f
C1556 VTAIL.n473 VSUBS 0.0295f
C1557 VTAIL.n474 VSUBS 0.013215f
C1558 VTAIL.n475 VSUBS 0.012481f
C1559 VTAIL.n476 VSUBS 0.023226f
C1560 VTAIL.n477 VSUBS 0.023226f
C1561 VTAIL.n478 VSUBS 0.012481f
C1562 VTAIL.n479 VSUBS 0.013215f
C1563 VTAIL.n480 VSUBS 0.0295f
C1564 VTAIL.n481 VSUBS 0.0295f
C1565 VTAIL.n482 VSUBS 0.013215f
C1566 VTAIL.n483 VSUBS 0.012481f
C1567 VTAIL.n484 VSUBS 0.023226f
C1568 VTAIL.n485 VSUBS 0.023226f
C1569 VTAIL.n486 VSUBS 0.012481f
C1570 VTAIL.n487 VSUBS 0.012848f
C1571 VTAIL.n488 VSUBS 0.012848f
C1572 VTAIL.n489 VSUBS 0.0295f
C1573 VTAIL.n490 VSUBS 0.0295f
C1574 VTAIL.n491 VSUBS 0.013215f
C1575 VTAIL.n492 VSUBS 0.012481f
C1576 VTAIL.n493 VSUBS 0.023226f
C1577 VTAIL.n494 VSUBS 0.023226f
C1578 VTAIL.n495 VSUBS 0.012481f
C1579 VTAIL.n496 VSUBS 0.013215f
C1580 VTAIL.n497 VSUBS 0.0295f
C1581 VTAIL.n498 VSUBS 0.0295f
C1582 VTAIL.n499 VSUBS 0.013215f
C1583 VTAIL.n500 VSUBS 0.012481f
C1584 VTAIL.n501 VSUBS 0.023226f
C1585 VTAIL.n502 VSUBS 0.023226f
C1586 VTAIL.n503 VSUBS 0.012481f
C1587 VTAIL.n504 VSUBS 0.013215f
C1588 VTAIL.n505 VSUBS 0.0295f
C1589 VTAIL.n506 VSUBS 0.0295f
C1590 VTAIL.n507 VSUBS 0.013215f
C1591 VTAIL.n508 VSUBS 0.012481f
C1592 VTAIL.n509 VSUBS 0.023226f
C1593 VTAIL.n510 VSUBS 0.023226f
C1594 VTAIL.n511 VSUBS 0.012481f
C1595 VTAIL.n512 VSUBS 0.013215f
C1596 VTAIL.n513 VSUBS 0.0295f
C1597 VTAIL.n514 VSUBS 0.0295f
C1598 VTAIL.n515 VSUBS 0.013215f
C1599 VTAIL.n516 VSUBS 0.012481f
C1600 VTAIL.n517 VSUBS 0.023226f
C1601 VTAIL.n518 VSUBS 0.023226f
C1602 VTAIL.n519 VSUBS 0.012481f
C1603 VTAIL.n520 VSUBS 0.013215f
C1604 VTAIL.n521 VSUBS 0.0295f
C1605 VTAIL.n522 VSUBS 0.0295f
C1606 VTAIL.n523 VSUBS 0.013215f
C1607 VTAIL.n524 VSUBS 0.012481f
C1608 VTAIL.n525 VSUBS 0.023226f
C1609 VTAIL.n526 VSUBS 0.023226f
C1610 VTAIL.n527 VSUBS 0.012481f
C1611 VTAIL.n528 VSUBS 0.013215f
C1612 VTAIL.n529 VSUBS 0.0295f
C1613 VTAIL.n530 VSUBS 0.072576f
C1614 VTAIL.n531 VSUBS 0.013215f
C1615 VTAIL.n532 VSUBS 0.024509f
C1616 VTAIL.n533 VSUBS 0.057493f
C1617 VTAIL.n534 VSUBS 0.055216f
C1618 VTAIL.n535 VSUBS 0.230701f
C1619 VTAIL.n536 VSUBS 0.024637f
C1620 VTAIL.n537 VSUBS 0.023226f
C1621 VTAIL.n538 VSUBS 0.012481f
C1622 VTAIL.n539 VSUBS 0.0295f
C1623 VTAIL.n540 VSUBS 0.013215f
C1624 VTAIL.n541 VSUBS 0.023226f
C1625 VTAIL.n542 VSUBS 0.012481f
C1626 VTAIL.n543 VSUBS 0.0295f
C1627 VTAIL.n544 VSUBS 0.013215f
C1628 VTAIL.n545 VSUBS 0.023226f
C1629 VTAIL.n546 VSUBS 0.012481f
C1630 VTAIL.n547 VSUBS 0.0295f
C1631 VTAIL.n548 VSUBS 0.013215f
C1632 VTAIL.n549 VSUBS 0.023226f
C1633 VTAIL.n550 VSUBS 0.012481f
C1634 VTAIL.n551 VSUBS 0.0295f
C1635 VTAIL.n552 VSUBS 0.013215f
C1636 VTAIL.n553 VSUBS 0.023226f
C1637 VTAIL.n554 VSUBS 0.012481f
C1638 VTAIL.n555 VSUBS 0.0295f
C1639 VTAIL.n556 VSUBS 0.013215f
C1640 VTAIL.n557 VSUBS 0.023226f
C1641 VTAIL.n558 VSUBS 0.012481f
C1642 VTAIL.n559 VSUBS 0.0295f
C1643 VTAIL.n560 VSUBS 0.013215f
C1644 VTAIL.n561 VSUBS 0.023226f
C1645 VTAIL.n562 VSUBS 0.012481f
C1646 VTAIL.n563 VSUBS 0.0295f
C1647 VTAIL.n564 VSUBS 0.0295f
C1648 VTAIL.n565 VSUBS 0.013215f
C1649 VTAIL.n566 VSUBS 0.023226f
C1650 VTAIL.n567 VSUBS 0.012481f
C1651 VTAIL.n568 VSUBS 0.0295f
C1652 VTAIL.n569 VSUBS 0.013215f
C1653 VTAIL.n570 VSUBS 0.261052f
C1654 VTAIL.t8 VSUBS 0.064153f
C1655 VTAIL.n571 VSUBS 0.022125f
C1656 VTAIL.n572 VSUBS 0.022191f
C1657 VTAIL.n573 VSUBS 0.012481f
C1658 VTAIL.n574 VSUBS 1.89832f
C1659 VTAIL.n575 VSUBS 0.023226f
C1660 VTAIL.n576 VSUBS 0.012481f
C1661 VTAIL.n577 VSUBS 0.013215f
C1662 VTAIL.n578 VSUBS 0.0295f
C1663 VTAIL.n579 VSUBS 0.0295f
C1664 VTAIL.n580 VSUBS 0.013215f
C1665 VTAIL.n581 VSUBS 0.012481f
C1666 VTAIL.n582 VSUBS 0.023226f
C1667 VTAIL.n583 VSUBS 0.023226f
C1668 VTAIL.n584 VSUBS 0.012481f
C1669 VTAIL.n585 VSUBS 0.013215f
C1670 VTAIL.n586 VSUBS 0.0295f
C1671 VTAIL.n587 VSUBS 0.0295f
C1672 VTAIL.n588 VSUBS 0.013215f
C1673 VTAIL.n589 VSUBS 0.012481f
C1674 VTAIL.n590 VSUBS 0.023226f
C1675 VTAIL.n591 VSUBS 0.023226f
C1676 VTAIL.n592 VSUBS 0.012481f
C1677 VTAIL.n593 VSUBS 0.012848f
C1678 VTAIL.n594 VSUBS 0.012848f
C1679 VTAIL.n595 VSUBS 0.0295f
C1680 VTAIL.n596 VSUBS 0.0295f
C1681 VTAIL.n597 VSUBS 0.013215f
C1682 VTAIL.n598 VSUBS 0.012481f
C1683 VTAIL.n599 VSUBS 0.023226f
C1684 VTAIL.n600 VSUBS 0.023226f
C1685 VTAIL.n601 VSUBS 0.012481f
C1686 VTAIL.n602 VSUBS 0.013215f
C1687 VTAIL.n603 VSUBS 0.0295f
C1688 VTAIL.n604 VSUBS 0.0295f
C1689 VTAIL.n605 VSUBS 0.013215f
C1690 VTAIL.n606 VSUBS 0.012481f
C1691 VTAIL.n607 VSUBS 0.023226f
C1692 VTAIL.n608 VSUBS 0.023226f
C1693 VTAIL.n609 VSUBS 0.012481f
C1694 VTAIL.n610 VSUBS 0.013215f
C1695 VTAIL.n611 VSUBS 0.0295f
C1696 VTAIL.n612 VSUBS 0.0295f
C1697 VTAIL.n613 VSUBS 0.013215f
C1698 VTAIL.n614 VSUBS 0.012481f
C1699 VTAIL.n615 VSUBS 0.023226f
C1700 VTAIL.n616 VSUBS 0.023226f
C1701 VTAIL.n617 VSUBS 0.012481f
C1702 VTAIL.n618 VSUBS 0.013215f
C1703 VTAIL.n619 VSUBS 0.0295f
C1704 VTAIL.n620 VSUBS 0.0295f
C1705 VTAIL.n621 VSUBS 0.013215f
C1706 VTAIL.n622 VSUBS 0.012481f
C1707 VTAIL.n623 VSUBS 0.023226f
C1708 VTAIL.n624 VSUBS 0.023226f
C1709 VTAIL.n625 VSUBS 0.012481f
C1710 VTAIL.n626 VSUBS 0.013215f
C1711 VTAIL.n627 VSUBS 0.0295f
C1712 VTAIL.n628 VSUBS 0.0295f
C1713 VTAIL.n629 VSUBS 0.013215f
C1714 VTAIL.n630 VSUBS 0.012481f
C1715 VTAIL.n631 VSUBS 0.023226f
C1716 VTAIL.n632 VSUBS 0.023226f
C1717 VTAIL.n633 VSUBS 0.012481f
C1718 VTAIL.n634 VSUBS 0.013215f
C1719 VTAIL.n635 VSUBS 0.0295f
C1720 VTAIL.n636 VSUBS 0.072576f
C1721 VTAIL.n637 VSUBS 0.013215f
C1722 VTAIL.n638 VSUBS 0.024509f
C1723 VTAIL.n639 VSUBS 0.057493f
C1724 VTAIL.n640 VSUBS 0.055216f
C1725 VTAIL.n641 VSUBS 0.230701f
C1726 VTAIL.t9 VSUBS 0.3568f
C1727 VTAIL.t12 VSUBS 0.3568f
C1728 VTAIL.n642 VSUBS 2.86999f
C1729 VTAIL.n643 VSUBS 0.899645f
C1730 VTAIL.n644 VSUBS 0.024637f
C1731 VTAIL.n645 VSUBS 0.023226f
C1732 VTAIL.n646 VSUBS 0.012481f
C1733 VTAIL.n647 VSUBS 0.0295f
C1734 VTAIL.n648 VSUBS 0.013215f
C1735 VTAIL.n649 VSUBS 0.023226f
C1736 VTAIL.n650 VSUBS 0.012481f
C1737 VTAIL.n651 VSUBS 0.0295f
C1738 VTAIL.n652 VSUBS 0.013215f
C1739 VTAIL.n653 VSUBS 0.023226f
C1740 VTAIL.n654 VSUBS 0.012481f
C1741 VTAIL.n655 VSUBS 0.0295f
C1742 VTAIL.n656 VSUBS 0.013215f
C1743 VTAIL.n657 VSUBS 0.023226f
C1744 VTAIL.n658 VSUBS 0.012481f
C1745 VTAIL.n659 VSUBS 0.0295f
C1746 VTAIL.n660 VSUBS 0.013215f
C1747 VTAIL.n661 VSUBS 0.023226f
C1748 VTAIL.n662 VSUBS 0.012481f
C1749 VTAIL.n663 VSUBS 0.0295f
C1750 VTAIL.n664 VSUBS 0.013215f
C1751 VTAIL.n665 VSUBS 0.023226f
C1752 VTAIL.n666 VSUBS 0.012481f
C1753 VTAIL.n667 VSUBS 0.0295f
C1754 VTAIL.n668 VSUBS 0.013215f
C1755 VTAIL.n669 VSUBS 0.023226f
C1756 VTAIL.n670 VSUBS 0.012481f
C1757 VTAIL.n671 VSUBS 0.0295f
C1758 VTAIL.n672 VSUBS 0.0295f
C1759 VTAIL.n673 VSUBS 0.013215f
C1760 VTAIL.n674 VSUBS 0.023226f
C1761 VTAIL.n675 VSUBS 0.012481f
C1762 VTAIL.n676 VSUBS 0.0295f
C1763 VTAIL.n677 VSUBS 0.013215f
C1764 VTAIL.n678 VSUBS 0.261052f
C1765 VTAIL.t10 VSUBS 0.064153f
C1766 VTAIL.n679 VSUBS 0.022125f
C1767 VTAIL.n680 VSUBS 0.022191f
C1768 VTAIL.n681 VSUBS 0.012481f
C1769 VTAIL.n682 VSUBS 1.89832f
C1770 VTAIL.n683 VSUBS 0.023226f
C1771 VTAIL.n684 VSUBS 0.012481f
C1772 VTAIL.n685 VSUBS 0.013215f
C1773 VTAIL.n686 VSUBS 0.0295f
C1774 VTAIL.n687 VSUBS 0.0295f
C1775 VTAIL.n688 VSUBS 0.013215f
C1776 VTAIL.n689 VSUBS 0.012481f
C1777 VTAIL.n690 VSUBS 0.023226f
C1778 VTAIL.n691 VSUBS 0.023226f
C1779 VTAIL.n692 VSUBS 0.012481f
C1780 VTAIL.n693 VSUBS 0.013215f
C1781 VTAIL.n694 VSUBS 0.0295f
C1782 VTAIL.n695 VSUBS 0.0295f
C1783 VTAIL.n696 VSUBS 0.013215f
C1784 VTAIL.n697 VSUBS 0.012481f
C1785 VTAIL.n698 VSUBS 0.023226f
C1786 VTAIL.n699 VSUBS 0.023226f
C1787 VTAIL.n700 VSUBS 0.012481f
C1788 VTAIL.n701 VSUBS 0.012848f
C1789 VTAIL.n702 VSUBS 0.012848f
C1790 VTAIL.n703 VSUBS 0.0295f
C1791 VTAIL.n704 VSUBS 0.0295f
C1792 VTAIL.n705 VSUBS 0.013215f
C1793 VTAIL.n706 VSUBS 0.012481f
C1794 VTAIL.n707 VSUBS 0.023226f
C1795 VTAIL.n708 VSUBS 0.023226f
C1796 VTAIL.n709 VSUBS 0.012481f
C1797 VTAIL.n710 VSUBS 0.013215f
C1798 VTAIL.n711 VSUBS 0.0295f
C1799 VTAIL.n712 VSUBS 0.0295f
C1800 VTAIL.n713 VSUBS 0.013215f
C1801 VTAIL.n714 VSUBS 0.012481f
C1802 VTAIL.n715 VSUBS 0.023226f
C1803 VTAIL.n716 VSUBS 0.023226f
C1804 VTAIL.n717 VSUBS 0.012481f
C1805 VTAIL.n718 VSUBS 0.013215f
C1806 VTAIL.n719 VSUBS 0.0295f
C1807 VTAIL.n720 VSUBS 0.0295f
C1808 VTAIL.n721 VSUBS 0.013215f
C1809 VTAIL.n722 VSUBS 0.012481f
C1810 VTAIL.n723 VSUBS 0.023226f
C1811 VTAIL.n724 VSUBS 0.023226f
C1812 VTAIL.n725 VSUBS 0.012481f
C1813 VTAIL.n726 VSUBS 0.013215f
C1814 VTAIL.n727 VSUBS 0.0295f
C1815 VTAIL.n728 VSUBS 0.0295f
C1816 VTAIL.n729 VSUBS 0.013215f
C1817 VTAIL.n730 VSUBS 0.012481f
C1818 VTAIL.n731 VSUBS 0.023226f
C1819 VTAIL.n732 VSUBS 0.023226f
C1820 VTAIL.n733 VSUBS 0.012481f
C1821 VTAIL.n734 VSUBS 0.013215f
C1822 VTAIL.n735 VSUBS 0.0295f
C1823 VTAIL.n736 VSUBS 0.0295f
C1824 VTAIL.n737 VSUBS 0.013215f
C1825 VTAIL.n738 VSUBS 0.012481f
C1826 VTAIL.n739 VSUBS 0.023226f
C1827 VTAIL.n740 VSUBS 0.023226f
C1828 VTAIL.n741 VSUBS 0.012481f
C1829 VTAIL.n742 VSUBS 0.013215f
C1830 VTAIL.n743 VSUBS 0.0295f
C1831 VTAIL.n744 VSUBS 0.072576f
C1832 VTAIL.n745 VSUBS 0.013215f
C1833 VTAIL.n746 VSUBS 0.024509f
C1834 VTAIL.n747 VSUBS 0.057493f
C1835 VTAIL.n748 VSUBS 0.055216f
C1836 VTAIL.n749 VSUBS 1.93879f
C1837 VTAIL.n750 VSUBS 0.024637f
C1838 VTAIL.n751 VSUBS 0.023226f
C1839 VTAIL.n752 VSUBS 0.012481f
C1840 VTAIL.n753 VSUBS 0.0295f
C1841 VTAIL.n754 VSUBS 0.013215f
C1842 VTAIL.n755 VSUBS 0.023226f
C1843 VTAIL.n756 VSUBS 0.012481f
C1844 VTAIL.n757 VSUBS 0.0295f
C1845 VTAIL.n758 VSUBS 0.013215f
C1846 VTAIL.n759 VSUBS 0.023226f
C1847 VTAIL.n760 VSUBS 0.012481f
C1848 VTAIL.n761 VSUBS 0.0295f
C1849 VTAIL.n762 VSUBS 0.013215f
C1850 VTAIL.n763 VSUBS 0.023226f
C1851 VTAIL.n764 VSUBS 0.012481f
C1852 VTAIL.n765 VSUBS 0.0295f
C1853 VTAIL.n766 VSUBS 0.013215f
C1854 VTAIL.n767 VSUBS 0.023226f
C1855 VTAIL.n768 VSUBS 0.012481f
C1856 VTAIL.n769 VSUBS 0.0295f
C1857 VTAIL.n770 VSUBS 0.013215f
C1858 VTAIL.n771 VSUBS 0.023226f
C1859 VTAIL.n772 VSUBS 0.012481f
C1860 VTAIL.n773 VSUBS 0.0295f
C1861 VTAIL.n774 VSUBS 0.013215f
C1862 VTAIL.n775 VSUBS 0.023226f
C1863 VTAIL.n776 VSUBS 0.012481f
C1864 VTAIL.n777 VSUBS 0.0295f
C1865 VTAIL.n778 VSUBS 0.013215f
C1866 VTAIL.n779 VSUBS 0.023226f
C1867 VTAIL.n780 VSUBS 0.012481f
C1868 VTAIL.n781 VSUBS 0.0295f
C1869 VTAIL.n782 VSUBS 0.013215f
C1870 VTAIL.n783 VSUBS 0.261052f
C1871 VTAIL.t4 VSUBS 0.064153f
C1872 VTAIL.n784 VSUBS 0.022125f
C1873 VTAIL.n785 VSUBS 0.022191f
C1874 VTAIL.n786 VSUBS 0.012481f
C1875 VTAIL.n787 VSUBS 1.89832f
C1876 VTAIL.n788 VSUBS 0.023226f
C1877 VTAIL.n789 VSUBS 0.012481f
C1878 VTAIL.n790 VSUBS 0.013215f
C1879 VTAIL.n791 VSUBS 0.0295f
C1880 VTAIL.n792 VSUBS 0.0295f
C1881 VTAIL.n793 VSUBS 0.013215f
C1882 VTAIL.n794 VSUBS 0.012481f
C1883 VTAIL.n795 VSUBS 0.023226f
C1884 VTAIL.n796 VSUBS 0.023226f
C1885 VTAIL.n797 VSUBS 0.012481f
C1886 VTAIL.n798 VSUBS 0.013215f
C1887 VTAIL.n799 VSUBS 0.0295f
C1888 VTAIL.n800 VSUBS 0.0295f
C1889 VTAIL.n801 VSUBS 0.0295f
C1890 VTAIL.n802 VSUBS 0.013215f
C1891 VTAIL.n803 VSUBS 0.012481f
C1892 VTAIL.n804 VSUBS 0.023226f
C1893 VTAIL.n805 VSUBS 0.023226f
C1894 VTAIL.n806 VSUBS 0.012481f
C1895 VTAIL.n807 VSUBS 0.012848f
C1896 VTAIL.n808 VSUBS 0.012848f
C1897 VTAIL.n809 VSUBS 0.0295f
C1898 VTAIL.n810 VSUBS 0.0295f
C1899 VTAIL.n811 VSUBS 0.013215f
C1900 VTAIL.n812 VSUBS 0.012481f
C1901 VTAIL.n813 VSUBS 0.023226f
C1902 VTAIL.n814 VSUBS 0.023226f
C1903 VTAIL.n815 VSUBS 0.012481f
C1904 VTAIL.n816 VSUBS 0.013215f
C1905 VTAIL.n817 VSUBS 0.0295f
C1906 VTAIL.n818 VSUBS 0.0295f
C1907 VTAIL.n819 VSUBS 0.013215f
C1908 VTAIL.n820 VSUBS 0.012481f
C1909 VTAIL.n821 VSUBS 0.023226f
C1910 VTAIL.n822 VSUBS 0.023226f
C1911 VTAIL.n823 VSUBS 0.012481f
C1912 VTAIL.n824 VSUBS 0.013215f
C1913 VTAIL.n825 VSUBS 0.0295f
C1914 VTAIL.n826 VSUBS 0.0295f
C1915 VTAIL.n827 VSUBS 0.013215f
C1916 VTAIL.n828 VSUBS 0.012481f
C1917 VTAIL.n829 VSUBS 0.023226f
C1918 VTAIL.n830 VSUBS 0.023226f
C1919 VTAIL.n831 VSUBS 0.012481f
C1920 VTAIL.n832 VSUBS 0.013215f
C1921 VTAIL.n833 VSUBS 0.0295f
C1922 VTAIL.n834 VSUBS 0.0295f
C1923 VTAIL.n835 VSUBS 0.013215f
C1924 VTAIL.n836 VSUBS 0.012481f
C1925 VTAIL.n837 VSUBS 0.023226f
C1926 VTAIL.n838 VSUBS 0.023226f
C1927 VTAIL.n839 VSUBS 0.012481f
C1928 VTAIL.n840 VSUBS 0.013215f
C1929 VTAIL.n841 VSUBS 0.0295f
C1930 VTAIL.n842 VSUBS 0.0295f
C1931 VTAIL.n843 VSUBS 0.013215f
C1932 VTAIL.n844 VSUBS 0.012481f
C1933 VTAIL.n845 VSUBS 0.023226f
C1934 VTAIL.n846 VSUBS 0.023226f
C1935 VTAIL.n847 VSUBS 0.012481f
C1936 VTAIL.n848 VSUBS 0.013215f
C1937 VTAIL.n849 VSUBS 0.0295f
C1938 VTAIL.n850 VSUBS 0.072576f
C1939 VTAIL.n851 VSUBS 0.013215f
C1940 VTAIL.n852 VSUBS 0.024509f
C1941 VTAIL.n853 VSUBS 0.057493f
C1942 VTAIL.n854 VSUBS 0.055216f
C1943 VTAIL.n855 VSUBS 1.93444f
C1944 VP.n0 VSUBS 0.038262f
C1945 VP.t5 VSUBS 3.66715f
C1946 VP.n1 VSUBS 0.024864f
C1947 VP.n2 VSUBS 0.02902f
C1948 VP.t7 VSUBS 3.66715f
C1949 VP.n3 VSUBS 0.054356f
C1950 VP.n4 VSUBS 0.02902f
C1951 VP.n5 VSUBS 0.032618f
C1952 VP.n6 VSUBS 0.02902f
C1953 VP.n7 VSUBS 0.05896f
C1954 VP.n8 VSUBS 0.038262f
C1955 VP.t2 VSUBS 3.66715f
C1956 VP.n9 VSUBS 0.024864f
C1957 VP.n10 VSUBS 0.02902f
C1958 VP.t1 VSUBS 3.66715f
C1959 VP.n11 VSUBS 0.054356f
C1960 VP.n12 VSUBS 0.02902f
C1961 VP.n13 VSUBS 0.032618f
C1962 VP.t6 VSUBS 3.86696f
C1963 VP.t0 VSUBS 3.66715f
C1964 VP.n14 VSUBS 1.34217f
C1965 VP.n15 VSUBS 1.33526f
C1966 VP.n16 VSUBS 0.251715f
C1967 VP.n17 VSUBS 0.02902f
C1968 VP.n18 VSUBS 0.054356f
C1969 VP.n19 VSUBS 0.042548f
C1970 VP.n20 VSUBS 0.042548f
C1971 VP.n21 VSUBS 0.02902f
C1972 VP.n22 VSUBS 0.02902f
C1973 VP.n23 VSUBS 0.02902f
C1974 VP.n24 VSUBS 0.032618f
C1975 VP.n25 VSUBS 1.27055f
C1976 VP.n26 VSUBS 0.049257f
C1977 VP.n27 VSUBS 0.055628f
C1978 VP.n28 VSUBS 0.02902f
C1979 VP.n29 VSUBS 0.02902f
C1980 VP.n30 VSUBS 0.02902f
C1981 VP.n31 VSUBS 0.05896f
C1982 VP.n32 VSUBS 0.042816f
C1983 VP.n33 VSUBS 1.36538f
C1984 VP.n34 VSUBS 1.86712f
C1985 VP.n35 VSUBS 1.88589f
C1986 VP.t4 VSUBS 3.66715f
C1987 VP.n36 VSUBS 1.36538f
C1988 VP.n37 VSUBS 0.042816f
C1989 VP.n38 VSUBS 0.038262f
C1990 VP.n39 VSUBS 0.02902f
C1991 VP.n40 VSUBS 0.02902f
C1992 VP.n41 VSUBS 0.024864f
C1993 VP.n42 VSUBS 0.055628f
C1994 VP.t3 VSUBS 3.66715f
C1995 VP.n43 VSUBS 1.27055f
C1996 VP.n44 VSUBS 0.049257f
C1997 VP.n45 VSUBS 0.02902f
C1998 VP.n46 VSUBS 0.02902f
C1999 VP.n47 VSUBS 0.02902f
C2000 VP.n48 VSUBS 0.054356f
C2001 VP.n49 VSUBS 0.042548f
C2002 VP.n50 VSUBS 0.042548f
C2003 VP.n51 VSUBS 0.02902f
C2004 VP.n52 VSUBS 0.02902f
C2005 VP.n53 VSUBS 0.02902f
C2006 VP.n54 VSUBS 0.032618f
C2007 VP.n55 VSUBS 1.27055f
C2008 VP.n56 VSUBS 0.049257f
C2009 VP.n57 VSUBS 0.055628f
C2010 VP.n58 VSUBS 0.02902f
C2011 VP.n59 VSUBS 0.02902f
C2012 VP.n60 VSUBS 0.02902f
C2013 VP.n61 VSUBS 0.05896f
C2014 VP.n62 VSUBS 0.042816f
C2015 VP.n63 VSUBS 1.36538f
C2016 VP.n64 VSUBS 0.042201f
.ends

