* NGSPICE file created from diff_pair_sample_1289.ext - technology: sky130A

.subckt diff_pair_sample_1289 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1498_n3422# sky130_fd_pr__pfet_01v8 ad=5.82825 pd=25.49 as=0 ps=0 w=12.27 l=0.16
X1 VDD1.t5 VP.t0 VTAIL.t5 w_n1498_n3422# sky130_fd_pr__pfet_01v8 ad=3.0675 pd=12.77 as=5.82825 ps=25.49 w=12.27 l=0.16
X2 VDD2.t5 VN.t0 VTAIL.t11 w_n1498_n3422# sky130_fd_pr__pfet_01v8 ad=5.82825 pd=25.49 as=3.0675 ps=12.77 w=12.27 l=0.16
X3 B.t8 B.t6 B.t7 w_n1498_n3422# sky130_fd_pr__pfet_01v8 ad=5.82825 pd=25.49 as=0 ps=0 w=12.27 l=0.16
X4 VTAIL.t7 VP.t1 VDD1.t4 w_n1498_n3422# sky130_fd_pr__pfet_01v8 ad=3.0675 pd=12.77 as=3.0675 ps=12.77 w=12.27 l=0.16
X5 VDD2.t4 VN.t1 VTAIL.t2 w_n1498_n3422# sky130_fd_pr__pfet_01v8 ad=3.0675 pd=12.77 as=5.82825 ps=25.49 w=12.27 l=0.16
X6 VDD2.t3 VN.t2 VTAIL.t1 w_n1498_n3422# sky130_fd_pr__pfet_01v8 ad=3.0675 pd=12.77 as=5.82825 ps=25.49 w=12.27 l=0.16
X7 VDD1.t3 VP.t2 VTAIL.t6 w_n1498_n3422# sky130_fd_pr__pfet_01v8 ad=5.82825 pd=25.49 as=3.0675 ps=12.77 w=12.27 l=0.16
X8 VTAIL.t10 VP.t3 VDD1.t2 w_n1498_n3422# sky130_fd_pr__pfet_01v8 ad=3.0675 pd=12.77 as=3.0675 ps=12.77 w=12.27 l=0.16
X9 VTAIL.t4 VN.t3 VDD2.t2 w_n1498_n3422# sky130_fd_pr__pfet_01v8 ad=3.0675 pd=12.77 as=3.0675 ps=12.77 w=12.27 l=0.16
X10 VDD1.t1 VP.t4 VTAIL.t9 w_n1498_n3422# sky130_fd_pr__pfet_01v8 ad=3.0675 pd=12.77 as=5.82825 ps=25.49 w=12.27 l=0.16
X11 B.t5 B.t3 B.t4 w_n1498_n3422# sky130_fd_pr__pfet_01v8 ad=5.82825 pd=25.49 as=0 ps=0 w=12.27 l=0.16
X12 VDD1.t0 VP.t5 VTAIL.t8 w_n1498_n3422# sky130_fd_pr__pfet_01v8 ad=5.82825 pd=25.49 as=3.0675 ps=12.77 w=12.27 l=0.16
X13 VTAIL.t3 VN.t4 VDD2.t1 w_n1498_n3422# sky130_fd_pr__pfet_01v8 ad=3.0675 pd=12.77 as=3.0675 ps=12.77 w=12.27 l=0.16
X14 VDD2.t0 VN.t5 VTAIL.t0 w_n1498_n3422# sky130_fd_pr__pfet_01v8 ad=5.82825 pd=25.49 as=3.0675 ps=12.77 w=12.27 l=0.16
X15 B.t2 B.t0 B.t1 w_n1498_n3422# sky130_fd_pr__pfet_01v8 ad=5.82825 pd=25.49 as=0 ps=0 w=12.27 l=0.16
R0 B.n100 B.t0 2099.58
R1 B.n106 B.t9 2099.58
R2 B.n32 B.t3 2099.58
R3 B.n38 B.t6 2099.58
R4 B.n352 B.n61 585
R5 B.n354 B.n353 585
R6 B.n355 B.n60 585
R7 B.n357 B.n356 585
R8 B.n358 B.n59 585
R9 B.n360 B.n359 585
R10 B.n361 B.n58 585
R11 B.n363 B.n362 585
R12 B.n364 B.n57 585
R13 B.n366 B.n365 585
R14 B.n367 B.n56 585
R15 B.n369 B.n368 585
R16 B.n370 B.n55 585
R17 B.n372 B.n371 585
R18 B.n373 B.n54 585
R19 B.n375 B.n374 585
R20 B.n376 B.n53 585
R21 B.n378 B.n377 585
R22 B.n379 B.n52 585
R23 B.n381 B.n380 585
R24 B.n382 B.n51 585
R25 B.n384 B.n383 585
R26 B.n385 B.n50 585
R27 B.n387 B.n386 585
R28 B.n388 B.n49 585
R29 B.n390 B.n389 585
R30 B.n391 B.n48 585
R31 B.n393 B.n392 585
R32 B.n394 B.n47 585
R33 B.n396 B.n395 585
R34 B.n397 B.n46 585
R35 B.n399 B.n398 585
R36 B.n400 B.n45 585
R37 B.n402 B.n401 585
R38 B.n403 B.n44 585
R39 B.n405 B.n404 585
R40 B.n406 B.n43 585
R41 B.n408 B.n407 585
R42 B.n409 B.n42 585
R43 B.n411 B.n410 585
R44 B.n412 B.n41 585
R45 B.n414 B.n413 585
R46 B.n416 B.n415 585
R47 B.n417 B.n37 585
R48 B.n419 B.n418 585
R49 B.n420 B.n36 585
R50 B.n422 B.n421 585
R51 B.n423 B.n35 585
R52 B.n425 B.n424 585
R53 B.n426 B.n34 585
R54 B.n428 B.n427 585
R55 B.n429 B.n31 585
R56 B.n432 B.n431 585
R57 B.n433 B.n30 585
R58 B.n435 B.n434 585
R59 B.n436 B.n29 585
R60 B.n438 B.n437 585
R61 B.n439 B.n28 585
R62 B.n441 B.n440 585
R63 B.n442 B.n27 585
R64 B.n444 B.n443 585
R65 B.n445 B.n26 585
R66 B.n447 B.n446 585
R67 B.n448 B.n25 585
R68 B.n450 B.n449 585
R69 B.n451 B.n24 585
R70 B.n453 B.n452 585
R71 B.n454 B.n23 585
R72 B.n456 B.n455 585
R73 B.n457 B.n22 585
R74 B.n459 B.n458 585
R75 B.n460 B.n21 585
R76 B.n462 B.n461 585
R77 B.n463 B.n20 585
R78 B.n465 B.n464 585
R79 B.n466 B.n19 585
R80 B.n468 B.n467 585
R81 B.n469 B.n18 585
R82 B.n471 B.n470 585
R83 B.n472 B.n17 585
R84 B.n474 B.n473 585
R85 B.n475 B.n16 585
R86 B.n477 B.n476 585
R87 B.n478 B.n15 585
R88 B.n480 B.n479 585
R89 B.n481 B.n14 585
R90 B.n483 B.n482 585
R91 B.n484 B.n13 585
R92 B.n486 B.n485 585
R93 B.n487 B.n12 585
R94 B.n489 B.n488 585
R95 B.n490 B.n11 585
R96 B.n492 B.n491 585
R97 B.n493 B.n10 585
R98 B.n351 B.n350 585
R99 B.n349 B.n62 585
R100 B.n348 B.n347 585
R101 B.n346 B.n63 585
R102 B.n345 B.n344 585
R103 B.n343 B.n64 585
R104 B.n342 B.n341 585
R105 B.n340 B.n65 585
R106 B.n339 B.n338 585
R107 B.n337 B.n66 585
R108 B.n336 B.n335 585
R109 B.n334 B.n67 585
R110 B.n333 B.n332 585
R111 B.n331 B.n68 585
R112 B.n330 B.n329 585
R113 B.n328 B.n69 585
R114 B.n327 B.n326 585
R115 B.n325 B.n70 585
R116 B.n324 B.n323 585
R117 B.n322 B.n71 585
R118 B.n321 B.n320 585
R119 B.n319 B.n72 585
R120 B.n318 B.n317 585
R121 B.n316 B.n73 585
R122 B.n315 B.n314 585
R123 B.n313 B.n74 585
R124 B.n312 B.n311 585
R125 B.n310 B.n75 585
R126 B.n309 B.n308 585
R127 B.n307 B.n76 585
R128 B.n306 B.n305 585
R129 B.n304 B.n77 585
R130 B.n303 B.n302 585
R131 B.n160 B.n129 585
R132 B.n162 B.n161 585
R133 B.n163 B.n128 585
R134 B.n165 B.n164 585
R135 B.n166 B.n127 585
R136 B.n168 B.n167 585
R137 B.n169 B.n126 585
R138 B.n171 B.n170 585
R139 B.n172 B.n125 585
R140 B.n174 B.n173 585
R141 B.n175 B.n124 585
R142 B.n177 B.n176 585
R143 B.n178 B.n123 585
R144 B.n180 B.n179 585
R145 B.n181 B.n122 585
R146 B.n183 B.n182 585
R147 B.n184 B.n121 585
R148 B.n186 B.n185 585
R149 B.n187 B.n120 585
R150 B.n189 B.n188 585
R151 B.n190 B.n119 585
R152 B.n192 B.n191 585
R153 B.n193 B.n118 585
R154 B.n195 B.n194 585
R155 B.n196 B.n117 585
R156 B.n198 B.n197 585
R157 B.n199 B.n116 585
R158 B.n201 B.n200 585
R159 B.n202 B.n115 585
R160 B.n204 B.n203 585
R161 B.n205 B.n114 585
R162 B.n207 B.n206 585
R163 B.n208 B.n113 585
R164 B.n210 B.n209 585
R165 B.n211 B.n112 585
R166 B.n213 B.n212 585
R167 B.n214 B.n111 585
R168 B.n216 B.n215 585
R169 B.n217 B.n110 585
R170 B.n219 B.n218 585
R171 B.n220 B.n109 585
R172 B.n222 B.n221 585
R173 B.n224 B.n223 585
R174 B.n225 B.n105 585
R175 B.n227 B.n226 585
R176 B.n228 B.n104 585
R177 B.n230 B.n229 585
R178 B.n231 B.n103 585
R179 B.n233 B.n232 585
R180 B.n234 B.n102 585
R181 B.n236 B.n235 585
R182 B.n237 B.n99 585
R183 B.n240 B.n239 585
R184 B.n241 B.n98 585
R185 B.n243 B.n242 585
R186 B.n244 B.n97 585
R187 B.n246 B.n245 585
R188 B.n247 B.n96 585
R189 B.n249 B.n248 585
R190 B.n250 B.n95 585
R191 B.n252 B.n251 585
R192 B.n253 B.n94 585
R193 B.n255 B.n254 585
R194 B.n256 B.n93 585
R195 B.n258 B.n257 585
R196 B.n259 B.n92 585
R197 B.n261 B.n260 585
R198 B.n262 B.n91 585
R199 B.n264 B.n263 585
R200 B.n265 B.n90 585
R201 B.n267 B.n266 585
R202 B.n268 B.n89 585
R203 B.n270 B.n269 585
R204 B.n271 B.n88 585
R205 B.n273 B.n272 585
R206 B.n274 B.n87 585
R207 B.n276 B.n275 585
R208 B.n277 B.n86 585
R209 B.n279 B.n278 585
R210 B.n280 B.n85 585
R211 B.n282 B.n281 585
R212 B.n283 B.n84 585
R213 B.n285 B.n284 585
R214 B.n286 B.n83 585
R215 B.n288 B.n287 585
R216 B.n289 B.n82 585
R217 B.n291 B.n290 585
R218 B.n292 B.n81 585
R219 B.n294 B.n293 585
R220 B.n295 B.n80 585
R221 B.n297 B.n296 585
R222 B.n298 B.n79 585
R223 B.n300 B.n299 585
R224 B.n301 B.n78 585
R225 B.n159 B.n158 585
R226 B.n157 B.n130 585
R227 B.n156 B.n155 585
R228 B.n154 B.n131 585
R229 B.n153 B.n152 585
R230 B.n151 B.n132 585
R231 B.n150 B.n149 585
R232 B.n148 B.n133 585
R233 B.n147 B.n146 585
R234 B.n145 B.n134 585
R235 B.n144 B.n143 585
R236 B.n142 B.n135 585
R237 B.n141 B.n140 585
R238 B.n139 B.n136 585
R239 B.n138 B.n137 585
R240 B.n2 B.n0 585
R241 B.n517 B.n1 585
R242 B.n516 B.n515 585
R243 B.n514 B.n3 585
R244 B.n513 B.n512 585
R245 B.n511 B.n4 585
R246 B.n510 B.n509 585
R247 B.n508 B.n5 585
R248 B.n507 B.n506 585
R249 B.n505 B.n6 585
R250 B.n504 B.n503 585
R251 B.n502 B.n7 585
R252 B.n501 B.n500 585
R253 B.n499 B.n8 585
R254 B.n498 B.n497 585
R255 B.n496 B.n9 585
R256 B.n495 B.n494 585
R257 B.n519 B.n518 585
R258 B.n158 B.n129 511.721
R259 B.n494 B.n493 511.721
R260 B.n302 B.n301 511.721
R261 B.n350 B.n61 511.721
R262 B.n158 B.n157 163.367
R263 B.n157 B.n156 163.367
R264 B.n156 B.n131 163.367
R265 B.n152 B.n131 163.367
R266 B.n152 B.n151 163.367
R267 B.n151 B.n150 163.367
R268 B.n150 B.n133 163.367
R269 B.n146 B.n133 163.367
R270 B.n146 B.n145 163.367
R271 B.n145 B.n144 163.367
R272 B.n144 B.n135 163.367
R273 B.n140 B.n135 163.367
R274 B.n140 B.n139 163.367
R275 B.n139 B.n138 163.367
R276 B.n138 B.n2 163.367
R277 B.n518 B.n2 163.367
R278 B.n518 B.n517 163.367
R279 B.n517 B.n516 163.367
R280 B.n516 B.n3 163.367
R281 B.n512 B.n3 163.367
R282 B.n512 B.n511 163.367
R283 B.n511 B.n510 163.367
R284 B.n510 B.n5 163.367
R285 B.n506 B.n5 163.367
R286 B.n506 B.n505 163.367
R287 B.n505 B.n504 163.367
R288 B.n504 B.n7 163.367
R289 B.n500 B.n7 163.367
R290 B.n500 B.n499 163.367
R291 B.n499 B.n498 163.367
R292 B.n498 B.n9 163.367
R293 B.n494 B.n9 163.367
R294 B.n162 B.n129 163.367
R295 B.n163 B.n162 163.367
R296 B.n164 B.n163 163.367
R297 B.n164 B.n127 163.367
R298 B.n168 B.n127 163.367
R299 B.n169 B.n168 163.367
R300 B.n170 B.n169 163.367
R301 B.n170 B.n125 163.367
R302 B.n174 B.n125 163.367
R303 B.n175 B.n174 163.367
R304 B.n176 B.n175 163.367
R305 B.n176 B.n123 163.367
R306 B.n180 B.n123 163.367
R307 B.n181 B.n180 163.367
R308 B.n182 B.n181 163.367
R309 B.n182 B.n121 163.367
R310 B.n186 B.n121 163.367
R311 B.n187 B.n186 163.367
R312 B.n188 B.n187 163.367
R313 B.n188 B.n119 163.367
R314 B.n192 B.n119 163.367
R315 B.n193 B.n192 163.367
R316 B.n194 B.n193 163.367
R317 B.n194 B.n117 163.367
R318 B.n198 B.n117 163.367
R319 B.n199 B.n198 163.367
R320 B.n200 B.n199 163.367
R321 B.n200 B.n115 163.367
R322 B.n204 B.n115 163.367
R323 B.n205 B.n204 163.367
R324 B.n206 B.n205 163.367
R325 B.n206 B.n113 163.367
R326 B.n210 B.n113 163.367
R327 B.n211 B.n210 163.367
R328 B.n212 B.n211 163.367
R329 B.n212 B.n111 163.367
R330 B.n216 B.n111 163.367
R331 B.n217 B.n216 163.367
R332 B.n218 B.n217 163.367
R333 B.n218 B.n109 163.367
R334 B.n222 B.n109 163.367
R335 B.n223 B.n222 163.367
R336 B.n223 B.n105 163.367
R337 B.n227 B.n105 163.367
R338 B.n228 B.n227 163.367
R339 B.n229 B.n228 163.367
R340 B.n229 B.n103 163.367
R341 B.n233 B.n103 163.367
R342 B.n234 B.n233 163.367
R343 B.n235 B.n234 163.367
R344 B.n235 B.n99 163.367
R345 B.n240 B.n99 163.367
R346 B.n241 B.n240 163.367
R347 B.n242 B.n241 163.367
R348 B.n242 B.n97 163.367
R349 B.n246 B.n97 163.367
R350 B.n247 B.n246 163.367
R351 B.n248 B.n247 163.367
R352 B.n248 B.n95 163.367
R353 B.n252 B.n95 163.367
R354 B.n253 B.n252 163.367
R355 B.n254 B.n253 163.367
R356 B.n254 B.n93 163.367
R357 B.n258 B.n93 163.367
R358 B.n259 B.n258 163.367
R359 B.n260 B.n259 163.367
R360 B.n260 B.n91 163.367
R361 B.n264 B.n91 163.367
R362 B.n265 B.n264 163.367
R363 B.n266 B.n265 163.367
R364 B.n266 B.n89 163.367
R365 B.n270 B.n89 163.367
R366 B.n271 B.n270 163.367
R367 B.n272 B.n271 163.367
R368 B.n272 B.n87 163.367
R369 B.n276 B.n87 163.367
R370 B.n277 B.n276 163.367
R371 B.n278 B.n277 163.367
R372 B.n278 B.n85 163.367
R373 B.n282 B.n85 163.367
R374 B.n283 B.n282 163.367
R375 B.n284 B.n283 163.367
R376 B.n284 B.n83 163.367
R377 B.n288 B.n83 163.367
R378 B.n289 B.n288 163.367
R379 B.n290 B.n289 163.367
R380 B.n290 B.n81 163.367
R381 B.n294 B.n81 163.367
R382 B.n295 B.n294 163.367
R383 B.n296 B.n295 163.367
R384 B.n296 B.n79 163.367
R385 B.n300 B.n79 163.367
R386 B.n301 B.n300 163.367
R387 B.n302 B.n77 163.367
R388 B.n306 B.n77 163.367
R389 B.n307 B.n306 163.367
R390 B.n308 B.n307 163.367
R391 B.n308 B.n75 163.367
R392 B.n312 B.n75 163.367
R393 B.n313 B.n312 163.367
R394 B.n314 B.n313 163.367
R395 B.n314 B.n73 163.367
R396 B.n318 B.n73 163.367
R397 B.n319 B.n318 163.367
R398 B.n320 B.n319 163.367
R399 B.n320 B.n71 163.367
R400 B.n324 B.n71 163.367
R401 B.n325 B.n324 163.367
R402 B.n326 B.n325 163.367
R403 B.n326 B.n69 163.367
R404 B.n330 B.n69 163.367
R405 B.n331 B.n330 163.367
R406 B.n332 B.n331 163.367
R407 B.n332 B.n67 163.367
R408 B.n336 B.n67 163.367
R409 B.n337 B.n336 163.367
R410 B.n338 B.n337 163.367
R411 B.n338 B.n65 163.367
R412 B.n342 B.n65 163.367
R413 B.n343 B.n342 163.367
R414 B.n344 B.n343 163.367
R415 B.n344 B.n63 163.367
R416 B.n348 B.n63 163.367
R417 B.n349 B.n348 163.367
R418 B.n350 B.n349 163.367
R419 B.n493 B.n492 163.367
R420 B.n492 B.n11 163.367
R421 B.n488 B.n11 163.367
R422 B.n488 B.n487 163.367
R423 B.n487 B.n486 163.367
R424 B.n486 B.n13 163.367
R425 B.n482 B.n13 163.367
R426 B.n482 B.n481 163.367
R427 B.n481 B.n480 163.367
R428 B.n480 B.n15 163.367
R429 B.n476 B.n15 163.367
R430 B.n476 B.n475 163.367
R431 B.n475 B.n474 163.367
R432 B.n474 B.n17 163.367
R433 B.n470 B.n17 163.367
R434 B.n470 B.n469 163.367
R435 B.n469 B.n468 163.367
R436 B.n468 B.n19 163.367
R437 B.n464 B.n19 163.367
R438 B.n464 B.n463 163.367
R439 B.n463 B.n462 163.367
R440 B.n462 B.n21 163.367
R441 B.n458 B.n21 163.367
R442 B.n458 B.n457 163.367
R443 B.n457 B.n456 163.367
R444 B.n456 B.n23 163.367
R445 B.n452 B.n23 163.367
R446 B.n452 B.n451 163.367
R447 B.n451 B.n450 163.367
R448 B.n450 B.n25 163.367
R449 B.n446 B.n25 163.367
R450 B.n446 B.n445 163.367
R451 B.n445 B.n444 163.367
R452 B.n444 B.n27 163.367
R453 B.n440 B.n27 163.367
R454 B.n440 B.n439 163.367
R455 B.n439 B.n438 163.367
R456 B.n438 B.n29 163.367
R457 B.n434 B.n29 163.367
R458 B.n434 B.n433 163.367
R459 B.n433 B.n432 163.367
R460 B.n432 B.n31 163.367
R461 B.n427 B.n31 163.367
R462 B.n427 B.n426 163.367
R463 B.n426 B.n425 163.367
R464 B.n425 B.n35 163.367
R465 B.n421 B.n35 163.367
R466 B.n421 B.n420 163.367
R467 B.n420 B.n419 163.367
R468 B.n419 B.n37 163.367
R469 B.n415 B.n37 163.367
R470 B.n415 B.n414 163.367
R471 B.n414 B.n41 163.367
R472 B.n410 B.n41 163.367
R473 B.n410 B.n409 163.367
R474 B.n409 B.n408 163.367
R475 B.n408 B.n43 163.367
R476 B.n404 B.n43 163.367
R477 B.n404 B.n403 163.367
R478 B.n403 B.n402 163.367
R479 B.n402 B.n45 163.367
R480 B.n398 B.n45 163.367
R481 B.n398 B.n397 163.367
R482 B.n397 B.n396 163.367
R483 B.n396 B.n47 163.367
R484 B.n392 B.n47 163.367
R485 B.n392 B.n391 163.367
R486 B.n391 B.n390 163.367
R487 B.n390 B.n49 163.367
R488 B.n386 B.n49 163.367
R489 B.n386 B.n385 163.367
R490 B.n385 B.n384 163.367
R491 B.n384 B.n51 163.367
R492 B.n380 B.n51 163.367
R493 B.n380 B.n379 163.367
R494 B.n379 B.n378 163.367
R495 B.n378 B.n53 163.367
R496 B.n374 B.n53 163.367
R497 B.n374 B.n373 163.367
R498 B.n373 B.n372 163.367
R499 B.n372 B.n55 163.367
R500 B.n368 B.n55 163.367
R501 B.n368 B.n367 163.367
R502 B.n367 B.n366 163.367
R503 B.n366 B.n57 163.367
R504 B.n362 B.n57 163.367
R505 B.n362 B.n361 163.367
R506 B.n361 B.n360 163.367
R507 B.n360 B.n59 163.367
R508 B.n356 B.n59 163.367
R509 B.n356 B.n355 163.367
R510 B.n355 B.n354 163.367
R511 B.n354 B.n61 163.367
R512 B.n100 B.t2 121.79
R513 B.n38 B.t7 121.79
R514 B.n106 B.t11 121.775
R515 B.n32 B.t4 121.775
R516 B.n101 B.t1 108.99
R517 B.n39 B.t8 108.99
R518 B.n107 B.t10 108.975
R519 B.n33 B.t5 108.975
R520 B.n238 B.n101 59.5399
R521 B.n108 B.n107 59.5399
R522 B.n430 B.n33 59.5399
R523 B.n40 B.n39 59.5399
R524 B.n495 B.n10 33.2493
R525 B.n352 B.n351 33.2493
R526 B.n303 B.n78 33.2493
R527 B.n160 B.n159 33.2493
R528 B B.n519 18.0485
R529 B.n101 B.n100 12.8005
R530 B.n107 B.n106 12.8005
R531 B.n33 B.n32 12.8005
R532 B.n39 B.n38 12.8005
R533 B.n491 B.n10 10.6151
R534 B.n491 B.n490 10.6151
R535 B.n490 B.n489 10.6151
R536 B.n489 B.n12 10.6151
R537 B.n485 B.n12 10.6151
R538 B.n485 B.n484 10.6151
R539 B.n484 B.n483 10.6151
R540 B.n483 B.n14 10.6151
R541 B.n479 B.n14 10.6151
R542 B.n479 B.n478 10.6151
R543 B.n478 B.n477 10.6151
R544 B.n477 B.n16 10.6151
R545 B.n473 B.n16 10.6151
R546 B.n473 B.n472 10.6151
R547 B.n472 B.n471 10.6151
R548 B.n471 B.n18 10.6151
R549 B.n467 B.n18 10.6151
R550 B.n467 B.n466 10.6151
R551 B.n466 B.n465 10.6151
R552 B.n465 B.n20 10.6151
R553 B.n461 B.n20 10.6151
R554 B.n461 B.n460 10.6151
R555 B.n460 B.n459 10.6151
R556 B.n459 B.n22 10.6151
R557 B.n455 B.n22 10.6151
R558 B.n455 B.n454 10.6151
R559 B.n454 B.n453 10.6151
R560 B.n453 B.n24 10.6151
R561 B.n449 B.n24 10.6151
R562 B.n449 B.n448 10.6151
R563 B.n448 B.n447 10.6151
R564 B.n447 B.n26 10.6151
R565 B.n443 B.n26 10.6151
R566 B.n443 B.n442 10.6151
R567 B.n442 B.n441 10.6151
R568 B.n441 B.n28 10.6151
R569 B.n437 B.n28 10.6151
R570 B.n437 B.n436 10.6151
R571 B.n436 B.n435 10.6151
R572 B.n435 B.n30 10.6151
R573 B.n431 B.n30 10.6151
R574 B.n429 B.n428 10.6151
R575 B.n428 B.n34 10.6151
R576 B.n424 B.n34 10.6151
R577 B.n424 B.n423 10.6151
R578 B.n423 B.n422 10.6151
R579 B.n422 B.n36 10.6151
R580 B.n418 B.n36 10.6151
R581 B.n418 B.n417 10.6151
R582 B.n417 B.n416 10.6151
R583 B.n413 B.n412 10.6151
R584 B.n412 B.n411 10.6151
R585 B.n411 B.n42 10.6151
R586 B.n407 B.n42 10.6151
R587 B.n407 B.n406 10.6151
R588 B.n406 B.n405 10.6151
R589 B.n405 B.n44 10.6151
R590 B.n401 B.n44 10.6151
R591 B.n401 B.n400 10.6151
R592 B.n400 B.n399 10.6151
R593 B.n399 B.n46 10.6151
R594 B.n395 B.n46 10.6151
R595 B.n395 B.n394 10.6151
R596 B.n394 B.n393 10.6151
R597 B.n393 B.n48 10.6151
R598 B.n389 B.n48 10.6151
R599 B.n389 B.n388 10.6151
R600 B.n388 B.n387 10.6151
R601 B.n387 B.n50 10.6151
R602 B.n383 B.n50 10.6151
R603 B.n383 B.n382 10.6151
R604 B.n382 B.n381 10.6151
R605 B.n381 B.n52 10.6151
R606 B.n377 B.n52 10.6151
R607 B.n377 B.n376 10.6151
R608 B.n376 B.n375 10.6151
R609 B.n375 B.n54 10.6151
R610 B.n371 B.n54 10.6151
R611 B.n371 B.n370 10.6151
R612 B.n370 B.n369 10.6151
R613 B.n369 B.n56 10.6151
R614 B.n365 B.n56 10.6151
R615 B.n365 B.n364 10.6151
R616 B.n364 B.n363 10.6151
R617 B.n363 B.n58 10.6151
R618 B.n359 B.n58 10.6151
R619 B.n359 B.n358 10.6151
R620 B.n358 B.n357 10.6151
R621 B.n357 B.n60 10.6151
R622 B.n353 B.n60 10.6151
R623 B.n353 B.n352 10.6151
R624 B.n304 B.n303 10.6151
R625 B.n305 B.n304 10.6151
R626 B.n305 B.n76 10.6151
R627 B.n309 B.n76 10.6151
R628 B.n310 B.n309 10.6151
R629 B.n311 B.n310 10.6151
R630 B.n311 B.n74 10.6151
R631 B.n315 B.n74 10.6151
R632 B.n316 B.n315 10.6151
R633 B.n317 B.n316 10.6151
R634 B.n317 B.n72 10.6151
R635 B.n321 B.n72 10.6151
R636 B.n322 B.n321 10.6151
R637 B.n323 B.n322 10.6151
R638 B.n323 B.n70 10.6151
R639 B.n327 B.n70 10.6151
R640 B.n328 B.n327 10.6151
R641 B.n329 B.n328 10.6151
R642 B.n329 B.n68 10.6151
R643 B.n333 B.n68 10.6151
R644 B.n334 B.n333 10.6151
R645 B.n335 B.n334 10.6151
R646 B.n335 B.n66 10.6151
R647 B.n339 B.n66 10.6151
R648 B.n340 B.n339 10.6151
R649 B.n341 B.n340 10.6151
R650 B.n341 B.n64 10.6151
R651 B.n345 B.n64 10.6151
R652 B.n346 B.n345 10.6151
R653 B.n347 B.n346 10.6151
R654 B.n347 B.n62 10.6151
R655 B.n351 B.n62 10.6151
R656 B.n161 B.n160 10.6151
R657 B.n161 B.n128 10.6151
R658 B.n165 B.n128 10.6151
R659 B.n166 B.n165 10.6151
R660 B.n167 B.n166 10.6151
R661 B.n167 B.n126 10.6151
R662 B.n171 B.n126 10.6151
R663 B.n172 B.n171 10.6151
R664 B.n173 B.n172 10.6151
R665 B.n173 B.n124 10.6151
R666 B.n177 B.n124 10.6151
R667 B.n178 B.n177 10.6151
R668 B.n179 B.n178 10.6151
R669 B.n179 B.n122 10.6151
R670 B.n183 B.n122 10.6151
R671 B.n184 B.n183 10.6151
R672 B.n185 B.n184 10.6151
R673 B.n185 B.n120 10.6151
R674 B.n189 B.n120 10.6151
R675 B.n190 B.n189 10.6151
R676 B.n191 B.n190 10.6151
R677 B.n191 B.n118 10.6151
R678 B.n195 B.n118 10.6151
R679 B.n196 B.n195 10.6151
R680 B.n197 B.n196 10.6151
R681 B.n197 B.n116 10.6151
R682 B.n201 B.n116 10.6151
R683 B.n202 B.n201 10.6151
R684 B.n203 B.n202 10.6151
R685 B.n203 B.n114 10.6151
R686 B.n207 B.n114 10.6151
R687 B.n208 B.n207 10.6151
R688 B.n209 B.n208 10.6151
R689 B.n209 B.n112 10.6151
R690 B.n213 B.n112 10.6151
R691 B.n214 B.n213 10.6151
R692 B.n215 B.n214 10.6151
R693 B.n215 B.n110 10.6151
R694 B.n219 B.n110 10.6151
R695 B.n220 B.n219 10.6151
R696 B.n221 B.n220 10.6151
R697 B.n225 B.n224 10.6151
R698 B.n226 B.n225 10.6151
R699 B.n226 B.n104 10.6151
R700 B.n230 B.n104 10.6151
R701 B.n231 B.n230 10.6151
R702 B.n232 B.n231 10.6151
R703 B.n232 B.n102 10.6151
R704 B.n236 B.n102 10.6151
R705 B.n237 B.n236 10.6151
R706 B.n239 B.n98 10.6151
R707 B.n243 B.n98 10.6151
R708 B.n244 B.n243 10.6151
R709 B.n245 B.n244 10.6151
R710 B.n245 B.n96 10.6151
R711 B.n249 B.n96 10.6151
R712 B.n250 B.n249 10.6151
R713 B.n251 B.n250 10.6151
R714 B.n251 B.n94 10.6151
R715 B.n255 B.n94 10.6151
R716 B.n256 B.n255 10.6151
R717 B.n257 B.n256 10.6151
R718 B.n257 B.n92 10.6151
R719 B.n261 B.n92 10.6151
R720 B.n262 B.n261 10.6151
R721 B.n263 B.n262 10.6151
R722 B.n263 B.n90 10.6151
R723 B.n267 B.n90 10.6151
R724 B.n268 B.n267 10.6151
R725 B.n269 B.n268 10.6151
R726 B.n269 B.n88 10.6151
R727 B.n273 B.n88 10.6151
R728 B.n274 B.n273 10.6151
R729 B.n275 B.n274 10.6151
R730 B.n275 B.n86 10.6151
R731 B.n279 B.n86 10.6151
R732 B.n280 B.n279 10.6151
R733 B.n281 B.n280 10.6151
R734 B.n281 B.n84 10.6151
R735 B.n285 B.n84 10.6151
R736 B.n286 B.n285 10.6151
R737 B.n287 B.n286 10.6151
R738 B.n287 B.n82 10.6151
R739 B.n291 B.n82 10.6151
R740 B.n292 B.n291 10.6151
R741 B.n293 B.n292 10.6151
R742 B.n293 B.n80 10.6151
R743 B.n297 B.n80 10.6151
R744 B.n298 B.n297 10.6151
R745 B.n299 B.n298 10.6151
R746 B.n299 B.n78 10.6151
R747 B.n159 B.n130 10.6151
R748 B.n155 B.n130 10.6151
R749 B.n155 B.n154 10.6151
R750 B.n154 B.n153 10.6151
R751 B.n153 B.n132 10.6151
R752 B.n149 B.n132 10.6151
R753 B.n149 B.n148 10.6151
R754 B.n148 B.n147 10.6151
R755 B.n147 B.n134 10.6151
R756 B.n143 B.n134 10.6151
R757 B.n143 B.n142 10.6151
R758 B.n142 B.n141 10.6151
R759 B.n141 B.n136 10.6151
R760 B.n137 B.n136 10.6151
R761 B.n137 B.n0 10.6151
R762 B.n515 B.n1 10.6151
R763 B.n515 B.n514 10.6151
R764 B.n514 B.n513 10.6151
R765 B.n513 B.n4 10.6151
R766 B.n509 B.n4 10.6151
R767 B.n509 B.n508 10.6151
R768 B.n508 B.n507 10.6151
R769 B.n507 B.n6 10.6151
R770 B.n503 B.n6 10.6151
R771 B.n503 B.n502 10.6151
R772 B.n502 B.n501 10.6151
R773 B.n501 B.n8 10.6151
R774 B.n497 B.n8 10.6151
R775 B.n497 B.n496 10.6151
R776 B.n496 B.n495 10.6151
R777 B.n431 B.n430 9.36635
R778 B.n413 B.n40 9.36635
R779 B.n221 B.n108 9.36635
R780 B.n239 B.n238 9.36635
R781 B.n519 B.n0 2.81026
R782 B.n519 B.n1 2.81026
R783 B.n430 B.n429 1.24928
R784 B.n416 B.n40 1.24928
R785 B.n224 B.n108 1.24928
R786 B.n238 B.n237 1.24928
R787 VP.n7 VP.t0 2105.37
R788 VP.n5 VP.t2 2105.37
R789 VP.n0 VP.t5 2105.37
R790 VP.n2 VP.t4 2105.37
R791 VP.n6 VP.t3 2045.49
R792 VP.n1 VP.t1 2045.49
R793 VP.n3 VP.n0 161.489
R794 VP.n8 VP.n7 161.3
R795 VP.n3 VP.n2 161.3
R796 VP.n5 VP.n4 161.3
R797 VP.n4 VP.n3 40.152
R798 VP.n6 VP.n5 36.5157
R799 VP.n7 VP.n6 36.5157
R800 VP.n1 VP.n0 36.5157
R801 VP.n2 VP.n1 36.5157
R802 VP.n8 VP.n4 0.189894
R803 VP VP.n8 0.0516364
R804 VTAIL.n7 VTAIL.t2 63.2675
R805 VTAIL.n11 VTAIL.t1 63.2665
R806 VTAIL.n2 VTAIL.t5 63.2665
R807 VTAIL.n10 VTAIL.t9 63.2663
R808 VTAIL.n9 VTAIL.n8 59.2537
R809 VTAIL.n6 VTAIL.n5 59.2537
R810 VTAIL.n1 VTAIL.n0 59.2535
R811 VTAIL.n4 VTAIL.n3 59.2535
R812 VTAIL.n6 VTAIL.n4 24.0824
R813 VTAIL.n11 VTAIL.n10 23.5134
R814 VTAIL.n0 VTAIL.t0 4.01435
R815 VTAIL.n0 VTAIL.t3 4.01435
R816 VTAIL.n3 VTAIL.t6 4.01435
R817 VTAIL.n3 VTAIL.t10 4.01435
R818 VTAIL.n8 VTAIL.t8 4.01435
R819 VTAIL.n8 VTAIL.t7 4.01435
R820 VTAIL.n5 VTAIL.t11 4.01435
R821 VTAIL.n5 VTAIL.t4 4.01435
R822 VTAIL.n9 VTAIL.n7 0.75481
R823 VTAIL.n2 VTAIL.n1 0.75481
R824 VTAIL.n7 VTAIL.n6 0.569465
R825 VTAIL.n10 VTAIL.n9 0.569465
R826 VTAIL.n4 VTAIL.n2 0.569465
R827 VTAIL VTAIL.n11 0.369034
R828 VTAIL VTAIL.n1 0.200931
R829 VDD1 VDD1.t0 80.4312
R830 VDD1.n1 VDD1.t3 80.3167
R831 VDD1.n1 VDD1.n0 76.0191
R832 VDD1.n3 VDD1.n2 75.9313
R833 VDD1.n3 VDD1.n1 37.0095
R834 VDD1.n2 VDD1.t4 4.01435
R835 VDD1.n2 VDD1.t1 4.01435
R836 VDD1.n0 VDD1.t2 4.01435
R837 VDD1.n0 VDD1.t5 4.01435
R838 VDD1 VDD1.n3 0.0845517
R839 VN.n2 VN.t2 2105.37
R840 VN.n0 VN.t5 2105.37
R841 VN.n6 VN.t0 2105.37
R842 VN.n4 VN.t1 2105.37
R843 VN.n1 VN.t4 2045.49
R844 VN.n5 VN.t3 2045.49
R845 VN.n7 VN.n4 161.489
R846 VN.n3 VN.n0 161.489
R847 VN.n3 VN.n2 161.3
R848 VN.n7 VN.n6 161.3
R849 VN VN.n7 40.5327
R850 VN.n1 VN.n0 36.5157
R851 VN.n2 VN.n1 36.5157
R852 VN.n6 VN.n5 36.5157
R853 VN.n5 VN.n4 36.5157
R854 VN VN.n3 0.0516364
R855 VDD2.n1 VDD2.t0 80.3167
R856 VDD2.n2 VDD2.t5 79.9463
R857 VDD2.n1 VDD2.n0 76.0191
R858 VDD2 VDD2.n3 76.0153
R859 VDD2.n2 VDD2.n1 36.142
R860 VDD2.n3 VDD2.t2 4.01435
R861 VDD2.n3 VDD2.t4 4.01435
R862 VDD2.n0 VDD2.t1 4.01435
R863 VDD2.n0 VDD2.t3 4.01435
R864 VDD2 VDD2.n2 0.485414
C0 B VDD1 1.46231f
C1 w_n1498_n3422# VDD1 1.72885f
C2 B VTAIL 2.4675f
C3 w_n1498_n3422# VTAIL 3.07109f
C4 B VP 0.971784f
C5 VP w_n1498_n3422# 2.398f
C6 VDD2 VDD1 0.580075f
C7 VDD2 VTAIL 14.331499f
C8 VN B 0.670468f
C9 VN w_n1498_n3422# 2.21066f
C10 VDD2 VP 0.266091f
C11 VTAIL VDD1 14.301701f
C12 VDD2 VN 1.91139f
C13 VP VDD1 2.02516f
C14 VP VTAIL 1.35719f
C15 VN VDD1 0.147253f
C16 VN VTAIL 1.34243f
C17 B w_n1498_n3422# 6.61617f
C18 VN VP 4.75389f
C19 VDD2 B 1.48309f
C20 VDD2 w_n1498_n3422# 1.74179f
C21 VDD2 VSUBS 1.188623f
C22 VDD1 VSUBS 1.543664f
C23 VTAIL VSUBS 0.597237f
C24 VN VSUBS 3.73754f
C25 VP VSUBS 1.088609f
C26 B VSUBS 2.324109f
C27 w_n1498_n3422# VSUBS 63.077797f
C28 VDD2.t0 VSUBS 2.30983f
C29 VDD2.t1 VSUBS 0.313185f
C30 VDD2.t3 VSUBS 0.313185f
C31 VDD2.n0 VSUBS 1.84959f
C32 VDD2.n1 VSUBS 2.12061f
C33 VDD2.t5 VSUBS 2.3074f
C34 VDD2.n2 VSUBS 2.13327f
C35 VDD2.t2 VSUBS 0.313185f
C36 VDD2.t4 VSUBS 0.313185f
C37 VDD2.n3 VSUBS 1.84957f
C38 VN.t5 VSUBS 0.300998f
C39 VN.n0 VSUBS 0.147144f
C40 VN.t4 VSUBS 0.297368f
C41 VN.n1 VSUBS 0.125312f
C42 VN.t2 VSUBS 0.300998f
C43 VN.n2 VSUBS 0.147062f
C44 VN.n3 VSUBS 0.110914f
C45 VN.t1 VSUBS 0.300998f
C46 VN.n4 VSUBS 0.147144f
C47 VN.t0 VSUBS 0.300998f
C48 VN.t3 VSUBS 0.297368f
C49 VN.n5 VSUBS 0.125312f
C50 VN.n6 VSUBS 0.147062f
C51 VN.n7 VSUBS 2.15474f
C52 VDD1.t0 VSUBS 2.61935f
C53 VDD1.t3 VSUBS 2.61847f
C54 VDD1.t2 VSUBS 0.355033f
C55 VDD1.t5 VSUBS 0.355033f
C56 VDD1.n0 VSUBS 2.09673f
C57 VDD1.n1 VSUBS 2.47039f
C58 VDD1.t4 VSUBS 0.355033f
C59 VDD1.t1 VSUBS 0.355033f
C60 VDD1.n2 VSUBS 2.09615f
C61 VDD1.n3 VSUBS 2.33475f
C62 VTAIL.t0 VSUBS 0.393498f
C63 VTAIL.t3 VSUBS 0.393498f
C64 VTAIL.n0 VSUBS 2.18855f
C65 VTAIL.n1 VSUBS 0.66434f
C66 VTAIL.t5 VSUBS 2.73803f
C67 VTAIL.n2 VSUBS 0.854964f
C68 VTAIL.t6 VSUBS 0.393498f
C69 VTAIL.t10 VSUBS 0.393498f
C70 VTAIL.n3 VSUBS 2.18855f
C71 VTAIL.n4 VSUBS 2.00601f
C72 VTAIL.t11 VSUBS 0.393498f
C73 VTAIL.t4 VSUBS 0.393498f
C74 VTAIL.n5 VSUBS 2.18856f
C75 VTAIL.n6 VSUBS 2.006f
C76 VTAIL.t2 VSUBS 2.73803f
C77 VTAIL.n7 VSUBS 0.85496f
C78 VTAIL.t8 VSUBS 0.393498f
C79 VTAIL.t7 VSUBS 0.393498f
C80 VTAIL.n8 VSUBS 2.18856f
C81 VTAIL.n9 VSUBS 0.696139f
C82 VTAIL.t9 VSUBS 2.73802f
C83 VTAIL.n10 VSUBS 2.11573f
C84 VTAIL.t1 VSUBS 2.73803f
C85 VTAIL.n11 VSUBS 2.09842f
C86 VP.t5 VSUBS 0.399902f
C87 VP.n0 VSUBS 0.195493f
C88 VP.t1 VSUBS 0.395079f
C89 VP.n1 VSUBS 0.166488f
C90 VP.t4 VSUBS 0.399902f
C91 VP.n2 VSUBS 0.195385f
C92 VP.n3 VSUBS 2.81588f
C93 VP.n4 VSUBS 2.78745f
C94 VP.t3 VSUBS 0.395079f
C95 VP.t2 VSUBS 0.399902f
C96 VP.n5 VSUBS 0.195385f
C97 VP.n6 VSUBS 0.166488f
C98 VP.t0 VSUBS 0.399902f
C99 VP.n7 VSUBS 0.195385f
C100 VP.n8 VSUBS 0.055184f
C101 B.n0 VSUBS 0.004856f
C102 B.n1 VSUBS 0.004856f
C103 B.n2 VSUBS 0.007679f
C104 B.n3 VSUBS 0.007679f
C105 B.n4 VSUBS 0.007679f
C106 B.n5 VSUBS 0.007679f
C107 B.n6 VSUBS 0.007679f
C108 B.n7 VSUBS 0.007679f
C109 B.n8 VSUBS 0.007679f
C110 B.n9 VSUBS 0.007679f
C111 B.n10 VSUBS 0.018366f
C112 B.n11 VSUBS 0.007679f
C113 B.n12 VSUBS 0.007679f
C114 B.n13 VSUBS 0.007679f
C115 B.n14 VSUBS 0.007679f
C116 B.n15 VSUBS 0.007679f
C117 B.n16 VSUBS 0.007679f
C118 B.n17 VSUBS 0.007679f
C119 B.n18 VSUBS 0.007679f
C120 B.n19 VSUBS 0.007679f
C121 B.n20 VSUBS 0.007679f
C122 B.n21 VSUBS 0.007679f
C123 B.n22 VSUBS 0.007679f
C124 B.n23 VSUBS 0.007679f
C125 B.n24 VSUBS 0.007679f
C126 B.n25 VSUBS 0.007679f
C127 B.n26 VSUBS 0.007679f
C128 B.n27 VSUBS 0.007679f
C129 B.n28 VSUBS 0.007679f
C130 B.n29 VSUBS 0.007679f
C131 B.n30 VSUBS 0.007679f
C132 B.n31 VSUBS 0.007679f
C133 B.t5 VSUBS 0.491242f
C134 B.t4 VSUBS 0.497906f
C135 B.t3 VSUBS 0.082818f
C136 B.n32 VSUBS 0.094059f
C137 B.n33 VSUBS 0.074352f
C138 B.n34 VSUBS 0.007679f
C139 B.n35 VSUBS 0.007679f
C140 B.n36 VSUBS 0.007679f
C141 B.n37 VSUBS 0.007679f
C142 B.t8 VSUBS 0.491233f
C143 B.t7 VSUBS 0.497897f
C144 B.t6 VSUBS 0.082818f
C145 B.n38 VSUBS 0.094068f
C146 B.n39 VSUBS 0.07436f
C147 B.n40 VSUBS 0.017791f
C148 B.n41 VSUBS 0.007679f
C149 B.n42 VSUBS 0.007679f
C150 B.n43 VSUBS 0.007679f
C151 B.n44 VSUBS 0.007679f
C152 B.n45 VSUBS 0.007679f
C153 B.n46 VSUBS 0.007679f
C154 B.n47 VSUBS 0.007679f
C155 B.n48 VSUBS 0.007679f
C156 B.n49 VSUBS 0.007679f
C157 B.n50 VSUBS 0.007679f
C158 B.n51 VSUBS 0.007679f
C159 B.n52 VSUBS 0.007679f
C160 B.n53 VSUBS 0.007679f
C161 B.n54 VSUBS 0.007679f
C162 B.n55 VSUBS 0.007679f
C163 B.n56 VSUBS 0.007679f
C164 B.n57 VSUBS 0.007679f
C165 B.n58 VSUBS 0.007679f
C166 B.n59 VSUBS 0.007679f
C167 B.n60 VSUBS 0.007679f
C168 B.n61 VSUBS 0.018366f
C169 B.n62 VSUBS 0.007679f
C170 B.n63 VSUBS 0.007679f
C171 B.n64 VSUBS 0.007679f
C172 B.n65 VSUBS 0.007679f
C173 B.n66 VSUBS 0.007679f
C174 B.n67 VSUBS 0.007679f
C175 B.n68 VSUBS 0.007679f
C176 B.n69 VSUBS 0.007679f
C177 B.n70 VSUBS 0.007679f
C178 B.n71 VSUBS 0.007679f
C179 B.n72 VSUBS 0.007679f
C180 B.n73 VSUBS 0.007679f
C181 B.n74 VSUBS 0.007679f
C182 B.n75 VSUBS 0.007679f
C183 B.n76 VSUBS 0.007679f
C184 B.n77 VSUBS 0.007679f
C185 B.n78 VSUBS 0.018366f
C186 B.n79 VSUBS 0.007679f
C187 B.n80 VSUBS 0.007679f
C188 B.n81 VSUBS 0.007679f
C189 B.n82 VSUBS 0.007679f
C190 B.n83 VSUBS 0.007679f
C191 B.n84 VSUBS 0.007679f
C192 B.n85 VSUBS 0.007679f
C193 B.n86 VSUBS 0.007679f
C194 B.n87 VSUBS 0.007679f
C195 B.n88 VSUBS 0.007679f
C196 B.n89 VSUBS 0.007679f
C197 B.n90 VSUBS 0.007679f
C198 B.n91 VSUBS 0.007679f
C199 B.n92 VSUBS 0.007679f
C200 B.n93 VSUBS 0.007679f
C201 B.n94 VSUBS 0.007679f
C202 B.n95 VSUBS 0.007679f
C203 B.n96 VSUBS 0.007679f
C204 B.n97 VSUBS 0.007679f
C205 B.n98 VSUBS 0.007679f
C206 B.n99 VSUBS 0.007679f
C207 B.t1 VSUBS 0.491233f
C208 B.t2 VSUBS 0.497897f
C209 B.t0 VSUBS 0.082818f
C210 B.n100 VSUBS 0.094068f
C211 B.n101 VSUBS 0.07436f
C212 B.n102 VSUBS 0.007679f
C213 B.n103 VSUBS 0.007679f
C214 B.n104 VSUBS 0.007679f
C215 B.n105 VSUBS 0.007679f
C216 B.t10 VSUBS 0.491242f
C217 B.t11 VSUBS 0.497906f
C218 B.t9 VSUBS 0.082818f
C219 B.n106 VSUBS 0.094059f
C220 B.n107 VSUBS 0.074352f
C221 B.n108 VSUBS 0.017791f
C222 B.n109 VSUBS 0.007679f
C223 B.n110 VSUBS 0.007679f
C224 B.n111 VSUBS 0.007679f
C225 B.n112 VSUBS 0.007679f
C226 B.n113 VSUBS 0.007679f
C227 B.n114 VSUBS 0.007679f
C228 B.n115 VSUBS 0.007679f
C229 B.n116 VSUBS 0.007679f
C230 B.n117 VSUBS 0.007679f
C231 B.n118 VSUBS 0.007679f
C232 B.n119 VSUBS 0.007679f
C233 B.n120 VSUBS 0.007679f
C234 B.n121 VSUBS 0.007679f
C235 B.n122 VSUBS 0.007679f
C236 B.n123 VSUBS 0.007679f
C237 B.n124 VSUBS 0.007679f
C238 B.n125 VSUBS 0.007679f
C239 B.n126 VSUBS 0.007679f
C240 B.n127 VSUBS 0.007679f
C241 B.n128 VSUBS 0.007679f
C242 B.n129 VSUBS 0.018366f
C243 B.n130 VSUBS 0.007679f
C244 B.n131 VSUBS 0.007679f
C245 B.n132 VSUBS 0.007679f
C246 B.n133 VSUBS 0.007679f
C247 B.n134 VSUBS 0.007679f
C248 B.n135 VSUBS 0.007679f
C249 B.n136 VSUBS 0.007679f
C250 B.n137 VSUBS 0.007679f
C251 B.n138 VSUBS 0.007679f
C252 B.n139 VSUBS 0.007679f
C253 B.n140 VSUBS 0.007679f
C254 B.n141 VSUBS 0.007679f
C255 B.n142 VSUBS 0.007679f
C256 B.n143 VSUBS 0.007679f
C257 B.n144 VSUBS 0.007679f
C258 B.n145 VSUBS 0.007679f
C259 B.n146 VSUBS 0.007679f
C260 B.n147 VSUBS 0.007679f
C261 B.n148 VSUBS 0.007679f
C262 B.n149 VSUBS 0.007679f
C263 B.n150 VSUBS 0.007679f
C264 B.n151 VSUBS 0.007679f
C265 B.n152 VSUBS 0.007679f
C266 B.n153 VSUBS 0.007679f
C267 B.n154 VSUBS 0.007679f
C268 B.n155 VSUBS 0.007679f
C269 B.n156 VSUBS 0.007679f
C270 B.n157 VSUBS 0.007679f
C271 B.n158 VSUBS 0.017996f
C272 B.n159 VSUBS 0.017996f
C273 B.n160 VSUBS 0.018366f
C274 B.n161 VSUBS 0.007679f
C275 B.n162 VSUBS 0.007679f
C276 B.n163 VSUBS 0.007679f
C277 B.n164 VSUBS 0.007679f
C278 B.n165 VSUBS 0.007679f
C279 B.n166 VSUBS 0.007679f
C280 B.n167 VSUBS 0.007679f
C281 B.n168 VSUBS 0.007679f
C282 B.n169 VSUBS 0.007679f
C283 B.n170 VSUBS 0.007679f
C284 B.n171 VSUBS 0.007679f
C285 B.n172 VSUBS 0.007679f
C286 B.n173 VSUBS 0.007679f
C287 B.n174 VSUBS 0.007679f
C288 B.n175 VSUBS 0.007679f
C289 B.n176 VSUBS 0.007679f
C290 B.n177 VSUBS 0.007679f
C291 B.n178 VSUBS 0.007679f
C292 B.n179 VSUBS 0.007679f
C293 B.n180 VSUBS 0.007679f
C294 B.n181 VSUBS 0.007679f
C295 B.n182 VSUBS 0.007679f
C296 B.n183 VSUBS 0.007679f
C297 B.n184 VSUBS 0.007679f
C298 B.n185 VSUBS 0.007679f
C299 B.n186 VSUBS 0.007679f
C300 B.n187 VSUBS 0.007679f
C301 B.n188 VSUBS 0.007679f
C302 B.n189 VSUBS 0.007679f
C303 B.n190 VSUBS 0.007679f
C304 B.n191 VSUBS 0.007679f
C305 B.n192 VSUBS 0.007679f
C306 B.n193 VSUBS 0.007679f
C307 B.n194 VSUBS 0.007679f
C308 B.n195 VSUBS 0.007679f
C309 B.n196 VSUBS 0.007679f
C310 B.n197 VSUBS 0.007679f
C311 B.n198 VSUBS 0.007679f
C312 B.n199 VSUBS 0.007679f
C313 B.n200 VSUBS 0.007679f
C314 B.n201 VSUBS 0.007679f
C315 B.n202 VSUBS 0.007679f
C316 B.n203 VSUBS 0.007679f
C317 B.n204 VSUBS 0.007679f
C318 B.n205 VSUBS 0.007679f
C319 B.n206 VSUBS 0.007679f
C320 B.n207 VSUBS 0.007679f
C321 B.n208 VSUBS 0.007679f
C322 B.n209 VSUBS 0.007679f
C323 B.n210 VSUBS 0.007679f
C324 B.n211 VSUBS 0.007679f
C325 B.n212 VSUBS 0.007679f
C326 B.n213 VSUBS 0.007679f
C327 B.n214 VSUBS 0.007679f
C328 B.n215 VSUBS 0.007679f
C329 B.n216 VSUBS 0.007679f
C330 B.n217 VSUBS 0.007679f
C331 B.n218 VSUBS 0.007679f
C332 B.n219 VSUBS 0.007679f
C333 B.n220 VSUBS 0.007679f
C334 B.n221 VSUBS 0.007227f
C335 B.n222 VSUBS 0.007679f
C336 B.n223 VSUBS 0.007679f
C337 B.n224 VSUBS 0.004291f
C338 B.n225 VSUBS 0.007679f
C339 B.n226 VSUBS 0.007679f
C340 B.n227 VSUBS 0.007679f
C341 B.n228 VSUBS 0.007679f
C342 B.n229 VSUBS 0.007679f
C343 B.n230 VSUBS 0.007679f
C344 B.n231 VSUBS 0.007679f
C345 B.n232 VSUBS 0.007679f
C346 B.n233 VSUBS 0.007679f
C347 B.n234 VSUBS 0.007679f
C348 B.n235 VSUBS 0.007679f
C349 B.n236 VSUBS 0.007679f
C350 B.n237 VSUBS 0.004291f
C351 B.n238 VSUBS 0.017791f
C352 B.n239 VSUBS 0.007227f
C353 B.n240 VSUBS 0.007679f
C354 B.n241 VSUBS 0.007679f
C355 B.n242 VSUBS 0.007679f
C356 B.n243 VSUBS 0.007679f
C357 B.n244 VSUBS 0.007679f
C358 B.n245 VSUBS 0.007679f
C359 B.n246 VSUBS 0.007679f
C360 B.n247 VSUBS 0.007679f
C361 B.n248 VSUBS 0.007679f
C362 B.n249 VSUBS 0.007679f
C363 B.n250 VSUBS 0.007679f
C364 B.n251 VSUBS 0.007679f
C365 B.n252 VSUBS 0.007679f
C366 B.n253 VSUBS 0.007679f
C367 B.n254 VSUBS 0.007679f
C368 B.n255 VSUBS 0.007679f
C369 B.n256 VSUBS 0.007679f
C370 B.n257 VSUBS 0.007679f
C371 B.n258 VSUBS 0.007679f
C372 B.n259 VSUBS 0.007679f
C373 B.n260 VSUBS 0.007679f
C374 B.n261 VSUBS 0.007679f
C375 B.n262 VSUBS 0.007679f
C376 B.n263 VSUBS 0.007679f
C377 B.n264 VSUBS 0.007679f
C378 B.n265 VSUBS 0.007679f
C379 B.n266 VSUBS 0.007679f
C380 B.n267 VSUBS 0.007679f
C381 B.n268 VSUBS 0.007679f
C382 B.n269 VSUBS 0.007679f
C383 B.n270 VSUBS 0.007679f
C384 B.n271 VSUBS 0.007679f
C385 B.n272 VSUBS 0.007679f
C386 B.n273 VSUBS 0.007679f
C387 B.n274 VSUBS 0.007679f
C388 B.n275 VSUBS 0.007679f
C389 B.n276 VSUBS 0.007679f
C390 B.n277 VSUBS 0.007679f
C391 B.n278 VSUBS 0.007679f
C392 B.n279 VSUBS 0.007679f
C393 B.n280 VSUBS 0.007679f
C394 B.n281 VSUBS 0.007679f
C395 B.n282 VSUBS 0.007679f
C396 B.n283 VSUBS 0.007679f
C397 B.n284 VSUBS 0.007679f
C398 B.n285 VSUBS 0.007679f
C399 B.n286 VSUBS 0.007679f
C400 B.n287 VSUBS 0.007679f
C401 B.n288 VSUBS 0.007679f
C402 B.n289 VSUBS 0.007679f
C403 B.n290 VSUBS 0.007679f
C404 B.n291 VSUBS 0.007679f
C405 B.n292 VSUBS 0.007679f
C406 B.n293 VSUBS 0.007679f
C407 B.n294 VSUBS 0.007679f
C408 B.n295 VSUBS 0.007679f
C409 B.n296 VSUBS 0.007679f
C410 B.n297 VSUBS 0.007679f
C411 B.n298 VSUBS 0.007679f
C412 B.n299 VSUBS 0.007679f
C413 B.n300 VSUBS 0.007679f
C414 B.n301 VSUBS 0.018366f
C415 B.n302 VSUBS 0.017996f
C416 B.n303 VSUBS 0.017996f
C417 B.n304 VSUBS 0.007679f
C418 B.n305 VSUBS 0.007679f
C419 B.n306 VSUBS 0.007679f
C420 B.n307 VSUBS 0.007679f
C421 B.n308 VSUBS 0.007679f
C422 B.n309 VSUBS 0.007679f
C423 B.n310 VSUBS 0.007679f
C424 B.n311 VSUBS 0.007679f
C425 B.n312 VSUBS 0.007679f
C426 B.n313 VSUBS 0.007679f
C427 B.n314 VSUBS 0.007679f
C428 B.n315 VSUBS 0.007679f
C429 B.n316 VSUBS 0.007679f
C430 B.n317 VSUBS 0.007679f
C431 B.n318 VSUBS 0.007679f
C432 B.n319 VSUBS 0.007679f
C433 B.n320 VSUBS 0.007679f
C434 B.n321 VSUBS 0.007679f
C435 B.n322 VSUBS 0.007679f
C436 B.n323 VSUBS 0.007679f
C437 B.n324 VSUBS 0.007679f
C438 B.n325 VSUBS 0.007679f
C439 B.n326 VSUBS 0.007679f
C440 B.n327 VSUBS 0.007679f
C441 B.n328 VSUBS 0.007679f
C442 B.n329 VSUBS 0.007679f
C443 B.n330 VSUBS 0.007679f
C444 B.n331 VSUBS 0.007679f
C445 B.n332 VSUBS 0.007679f
C446 B.n333 VSUBS 0.007679f
C447 B.n334 VSUBS 0.007679f
C448 B.n335 VSUBS 0.007679f
C449 B.n336 VSUBS 0.007679f
C450 B.n337 VSUBS 0.007679f
C451 B.n338 VSUBS 0.007679f
C452 B.n339 VSUBS 0.007679f
C453 B.n340 VSUBS 0.007679f
C454 B.n341 VSUBS 0.007679f
C455 B.n342 VSUBS 0.007679f
C456 B.n343 VSUBS 0.007679f
C457 B.n344 VSUBS 0.007679f
C458 B.n345 VSUBS 0.007679f
C459 B.n346 VSUBS 0.007679f
C460 B.n347 VSUBS 0.007679f
C461 B.n348 VSUBS 0.007679f
C462 B.n349 VSUBS 0.007679f
C463 B.n350 VSUBS 0.017996f
C464 B.n351 VSUBS 0.018887f
C465 B.n352 VSUBS 0.017475f
C466 B.n353 VSUBS 0.007679f
C467 B.n354 VSUBS 0.007679f
C468 B.n355 VSUBS 0.007679f
C469 B.n356 VSUBS 0.007679f
C470 B.n357 VSUBS 0.007679f
C471 B.n358 VSUBS 0.007679f
C472 B.n359 VSUBS 0.007679f
C473 B.n360 VSUBS 0.007679f
C474 B.n361 VSUBS 0.007679f
C475 B.n362 VSUBS 0.007679f
C476 B.n363 VSUBS 0.007679f
C477 B.n364 VSUBS 0.007679f
C478 B.n365 VSUBS 0.007679f
C479 B.n366 VSUBS 0.007679f
C480 B.n367 VSUBS 0.007679f
C481 B.n368 VSUBS 0.007679f
C482 B.n369 VSUBS 0.007679f
C483 B.n370 VSUBS 0.007679f
C484 B.n371 VSUBS 0.007679f
C485 B.n372 VSUBS 0.007679f
C486 B.n373 VSUBS 0.007679f
C487 B.n374 VSUBS 0.007679f
C488 B.n375 VSUBS 0.007679f
C489 B.n376 VSUBS 0.007679f
C490 B.n377 VSUBS 0.007679f
C491 B.n378 VSUBS 0.007679f
C492 B.n379 VSUBS 0.007679f
C493 B.n380 VSUBS 0.007679f
C494 B.n381 VSUBS 0.007679f
C495 B.n382 VSUBS 0.007679f
C496 B.n383 VSUBS 0.007679f
C497 B.n384 VSUBS 0.007679f
C498 B.n385 VSUBS 0.007679f
C499 B.n386 VSUBS 0.007679f
C500 B.n387 VSUBS 0.007679f
C501 B.n388 VSUBS 0.007679f
C502 B.n389 VSUBS 0.007679f
C503 B.n390 VSUBS 0.007679f
C504 B.n391 VSUBS 0.007679f
C505 B.n392 VSUBS 0.007679f
C506 B.n393 VSUBS 0.007679f
C507 B.n394 VSUBS 0.007679f
C508 B.n395 VSUBS 0.007679f
C509 B.n396 VSUBS 0.007679f
C510 B.n397 VSUBS 0.007679f
C511 B.n398 VSUBS 0.007679f
C512 B.n399 VSUBS 0.007679f
C513 B.n400 VSUBS 0.007679f
C514 B.n401 VSUBS 0.007679f
C515 B.n402 VSUBS 0.007679f
C516 B.n403 VSUBS 0.007679f
C517 B.n404 VSUBS 0.007679f
C518 B.n405 VSUBS 0.007679f
C519 B.n406 VSUBS 0.007679f
C520 B.n407 VSUBS 0.007679f
C521 B.n408 VSUBS 0.007679f
C522 B.n409 VSUBS 0.007679f
C523 B.n410 VSUBS 0.007679f
C524 B.n411 VSUBS 0.007679f
C525 B.n412 VSUBS 0.007679f
C526 B.n413 VSUBS 0.007227f
C527 B.n414 VSUBS 0.007679f
C528 B.n415 VSUBS 0.007679f
C529 B.n416 VSUBS 0.004291f
C530 B.n417 VSUBS 0.007679f
C531 B.n418 VSUBS 0.007679f
C532 B.n419 VSUBS 0.007679f
C533 B.n420 VSUBS 0.007679f
C534 B.n421 VSUBS 0.007679f
C535 B.n422 VSUBS 0.007679f
C536 B.n423 VSUBS 0.007679f
C537 B.n424 VSUBS 0.007679f
C538 B.n425 VSUBS 0.007679f
C539 B.n426 VSUBS 0.007679f
C540 B.n427 VSUBS 0.007679f
C541 B.n428 VSUBS 0.007679f
C542 B.n429 VSUBS 0.004291f
C543 B.n430 VSUBS 0.017791f
C544 B.n431 VSUBS 0.007227f
C545 B.n432 VSUBS 0.007679f
C546 B.n433 VSUBS 0.007679f
C547 B.n434 VSUBS 0.007679f
C548 B.n435 VSUBS 0.007679f
C549 B.n436 VSUBS 0.007679f
C550 B.n437 VSUBS 0.007679f
C551 B.n438 VSUBS 0.007679f
C552 B.n439 VSUBS 0.007679f
C553 B.n440 VSUBS 0.007679f
C554 B.n441 VSUBS 0.007679f
C555 B.n442 VSUBS 0.007679f
C556 B.n443 VSUBS 0.007679f
C557 B.n444 VSUBS 0.007679f
C558 B.n445 VSUBS 0.007679f
C559 B.n446 VSUBS 0.007679f
C560 B.n447 VSUBS 0.007679f
C561 B.n448 VSUBS 0.007679f
C562 B.n449 VSUBS 0.007679f
C563 B.n450 VSUBS 0.007679f
C564 B.n451 VSUBS 0.007679f
C565 B.n452 VSUBS 0.007679f
C566 B.n453 VSUBS 0.007679f
C567 B.n454 VSUBS 0.007679f
C568 B.n455 VSUBS 0.007679f
C569 B.n456 VSUBS 0.007679f
C570 B.n457 VSUBS 0.007679f
C571 B.n458 VSUBS 0.007679f
C572 B.n459 VSUBS 0.007679f
C573 B.n460 VSUBS 0.007679f
C574 B.n461 VSUBS 0.007679f
C575 B.n462 VSUBS 0.007679f
C576 B.n463 VSUBS 0.007679f
C577 B.n464 VSUBS 0.007679f
C578 B.n465 VSUBS 0.007679f
C579 B.n466 VSUBS 0.007679f
C580 B.n467 VSUBS 0.007679f
C581 B.n468 VSUBS 0.007679f
C582 B.n469 VSUBS 0.007679f
C583 B.n470 VSUBS 0.007679f
C584 B.n471 VSUBS 0.007679f
C585 B.n472 VSUBS 0.007679f
C586 B.n473 VSUBS 0.007679f
C587 B.n474 VSUBS 0.007679f
C588 B.n475 VSUBS 0.007679f
C589 B.n476 VSUBS 0.007679f
C590 B.n477 VSUBS 0.007679f
C591 B.n478 VSUBS 0.007679f
C592 B.n479 VSUBS 0.007679f
C593 B.n480 VSUBS 0.007679f
C594 B.n481 VSUBS 0.007679f
C595 B.n482 VSUBS 0.007679f
C596 B.n483 VSUBS 0.007679f
C597 B.n484 VSUBS 0.007679f
C598 B.n485 VSUBS 0.007679f
C599 B.n486 VSUBS 0.007679f
C600 B.n487 VSUBS 0.007679f
C601 B.n488 VSUBS 0.007679f
C602 B.n489 VSUBS 0.007679f
C603 B.n490 VSUBS 0.007679f
C604 B.n491 VSUBS 0.007679f
C605 B.n492 VSUBS 0.007679f
C606 B.n493 VSUBS 0.018366f
C607 B.n494 VSUBS 0.017996f
C608 B.n495 VSUBS 0.017996f
C609 B.n496 VSUBS 0.007679f
C610 B.n497 VSUBS 0.007679f
C611 B.n498 VSUBS 0.007679f
C612 B.n499 VSUBS 0.007679f
C613 B.n500 VSUBS 0.007679f
C614 B.n501 VSUBS 0.007679f
C615 B.n502 VSUBS 0.007679f
C616 B.n503 VSUBS 0.007679f
C617 B.n504 VSUBS 0.007679f
C618 B.n505 VSUBS 0.007679f
C619 B.n506 VSUBS 0.007679f
C620 B.n507 VSUBS 0.007679f
C621 B.n508 VSUBS 0.007679f
C622 B.n509 VSUBS 0.007679f
C623 B.n510 VSUBS 0.007679f
C624 B.n511 VSUBS 0.007679f
C625 B.n512 VSUBS 0.007679f
C626 B.n513 VSUBS 0.007679f
C627 B.n514 VSUBS 0.007679f
C628 B.n515 VSUBS 0.007679f
C629 B.n516 VSUBS 0.007679f
C630 B.n517 VSUBS 0.007679f
C631 B.n518 VSUBS 0.007679f
C632 B.n519 VSUBS 0.017388f
.ends

