* NGSPICE file created from diff_pair_sample_0117.ext - technology: sky130A

.subckt diff_pair_sample_0117 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=4.8789 pd=25.8 as=0 ps=0 w=12.51 l=1.09
X1 VDD2.t9 VN.t0 VTAIL.t13 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=2.06415 pd=12.84 as=2.06415 ps=12.84 w=12.51 l=1.09
X2 VTAIL.t9 VN.t1 VDD2.t8 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=2.06415 pd=12.84 as=2.06415 ps=12.84 w=12.51 l=1.09
X3 VDD1.t9 VP.t0 VTAIL.t0 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=2.06415 pd=12.84 as=4.8789 ps=25.8 w=12.51 l=1.09
X4 VTAIL.t7 VP.t1 VDD1.t8 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=2.06415 pd=12.84 as=2.06415 ps=12.84 w=12.51 l=1.09
X5 VTAIL.t11 VN.t2 VDD2.t7 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=2.06415 pd=12.84 as=2.06415 ps=12.84 w=12.51 l=1.09
X6 VTAIL.t6 VP.t2 VDD1.t7 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=2.06415 pd=12.84 as=2.06415 ps=12.84 w=12.51 l=1.09
X7 VTAIL.t14 VN.t3 VDD2.t6 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=2.06415 pd=12.84 as=2.06415 ps=12.84 w=12.51 l=1.09
X8 VDD2.t5 VN.t4 VTAIL.t10 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=2.06415 pd=12.84 as=2.06415 ps=12.84 w=12.51 l=1.09
X9 VDD1.t6 VP.t3 VTAIL.t3 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=4.8789 pd=25.8 as=2.06415 ps=12.84 w=12.51 l=1.09
X10 B.t8 B.t6 B.t7 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=4.8789 pd=25.8 as=0 ps=0 w=12.51 l=1.09
X11 VDD2.t4 VN.t5 VTAIL.t17 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=2.06415 pd=12.84 as=4.8789 ps=25.8 w=12.51 l=1.09
X12 VDD1.t5 VP.t4 VTAIL.t8 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=2.06415 pd=12.84 as=2.06415 ps=12.84 w=12.51 l=1.09
X13 VDD2.t3 VN.t6 VTAIL.t12 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=4.8789 pd=25.8 as=2.06415 ps=12.84 w=12.51 l=1.09
X14 VTAIL.t5 VP.t5 VDD1.t4 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=2.06415 pd=12.84 as=2.06415 ps=12.84 w=12.51 l=1.09
X15 VDD2.t2 VN.t7 VTAIL.t18 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=4.8789 pd=25.8 as=2.06415 ps=12.84 w=12.51 l=1.09
X16 B.t5 B.t3 B.t4 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=4.8789 pd=25.8 as=0 ps=0 w=12.51 l=1.09
X17 B.t2 B.t0 B.t1 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=4.8789 pd=25.8 as=0 ps=0 w=12.51 l=1.09
X18 VDD2.t1 VN.t8 VTAIL.t15 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=2.06415 pd=12.84 as=4.8789 ps=25.8 w=12.51 l=1.09
X19 VTAIL.t4 VP.t6 VDD1.t3 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=2.06415 pd=12.84 as=2.06415 ps=12.84 w=12.51 l=1.09
X20 VTAIL.t16 VN.t9 VDD2.t0 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=2.06415 pd=12.84 as=2.06415 ps=12.84 w=12.51 l=1.09
X21 VDD1.t2 VP.t7 VTAIL.t2 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=2.06415 pd=12.84 as=4.8789 ps=25.8 w=12.51 l=1.09
X22 VDD1.t1 VP.t8 VTAIL.t19 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=2.06415 pd=12.84 as=2.06415 ps=12.84 w=12.51 l=1.09
X23 VDD1.t0 VP.t9 VTAIL.t1 w_n2674_n3470# sky130_fd_pr__pfet_01v8 ad=4.8789 pd=25.8 as=2.06415 ps=12.84 w=12.51 l=1.09
R0 B.n468 B.n467 585
R1 B.n469 B.n70 585
R2 B.n471 B.n470 585
R3 B.n472 B.n69 585
R4 B.n474 B.n473 585
R5 B.n475 B.n68 585
R6 B.n477 B.n476 585
R7 B.n478 B.n67 585
R8 B.n480 B.n479 585
R9 B.n481 B.n66 585
R10 B.n483 B.n482 585
R11 B.n484 B.n65 585
R12 B.n486 B.n485 585
R13 B.n487 B.n64 585
R14 B.n489 B.n488 585
R15 B.n490 B.n63 585
R16 B.n492 B.n491 585
R17 B.n493 B.n62 585
R18 B.n495 B.n494 585
R19 B.n496 B.n61 585
R20 B.n498 B.n497 585
R21 B.n499 B.n60 585
R22 B.n501 B.n500 585
R23 B.n502 B.n59 585
R24 B.n504 B.n503 585
R25 B.n505 B.n58 585
R26 B.n507 B.n506 585
R27 B.n508 B.n57 585
R28 B.n510 B.n509 585
R29 B.n511 B.n56 585
R30 B.n513 B.n512 585
R31 B.n514 B.n55 585
R32 B.n516 B.n515 585
R33 B.n517 B.n54 585
R34 B.n519 B.n518 585
R35 B.n520 B.n53 585
R36 B.n522 B.n521 585
R37 B.n523 B.n52 585
R38 B.n525 B.n524 585
R39 B.n526 B.n51 585
R40 B.n528 B.n527 585
R41 B.n529 B.n50 585
R42 B.n531 B.n530 585
R43 B.n533 B.n47 585
R44 B.n535 B.n534 585
R45 B.n536 B.n46 585
R46 B.n538 B.n537 585
R47 B.n539 B.n45 585
R48 B.n541 B.n540 585
R49 B.n542 B.n44 585
R50 B.n544 B.n543 585
R51 B.n545 B.n43 585
R52 B.n547 B.n546 585
R53 B.n549 B.n548 585
R54 B.n550 B.n39 585
R55 B.n552 B.n551 585
R56 B.n553 B.n38 585
R57 B.n555 B.n554 585
R58 B.n556 B.n37 585
R59 B.n558 B.n557 585
R60 B.n559 B.n36 585
R61 B.n561 B.n560 585
R62 B.n562 B.n35 585
R63 B.n564 B.n563 585
R64 B.n565 B.n34 585
R65 B.n567 B.n566 585
R66 B.n568 B.n33 585
R67 B.n570 B.n569 585
R68 B.n571 B.n32 585
R69 B.n573 B.n572 585
R70 B.n574 B.n31 585
R71 B.n576 B.n575 585
R72 B.n577 B.n30 585
R73 B.n579 B.n578 585
R74 B.n580 B.n29 585
R75 B.n582 B.n581 585
R76 B.n583 B.n28 585
R77 B.n585 B.n584 585
R78 B.n586 B.n27 585
R79 B.n588 B.n587 585
R80 B.n589 B.n26 585
R81 B.n591 B.n590 585
R82 B.n592 B.n25 585
R83 B.n594 B.n593 585
R84 B.n595 B.n24 585
R85 B.n597 B.n596 585
R86 B.n598 B.n23 585
R87 B.n600 B.n599 585
R88 B.n601 B.n22 585
R89 B.n603 B.n602 585
R90 B.n604 B.n21 585
R91 B.n606 B.n605 585
R92 B.n607 B.n20 585
R93 B.n609 B.n608 585
R94 B.n610 B.n19 585
R95 B.n612 B.n611 585
R96 B.n466 B.n71 585
R97 B.n465 B.n464 585
R98 B.n463 B.n72 585
R99 B.n462 B.n461 585
R100 B.n460 B.n73 585
R101 B.n459 B.n458 585
R102 B.n457 B.n74 585
R103 B.n456 B.n455 585
R104 B.n454 B.n75 585
R105 B.n453 B.n452 585
R106 B.n451 B.n76 585
R107 B.n450 B.n449 585
R108 B.n448 B.n77 585
R109 B.n447 B.n446 585
R110 B.n445 B.n78 585
R111 B.n444 B.n443 585
R112 B.n442 B.n79 585
R113 B.n441 B.n440 585
R114 B.n439 B.n80 585
R115 B.n438 B.n437 585
R116 B.n436 B.n81 585
R117 B.n435 B.n434 585
R118 B.n433 B.n82 585
R119 B.n432 B.n431 585
R120 B.n430 B.n83 585
R121 B.n429 B.n428 585
R122 B.n427 B.n84 585
R123 B.n426 B.n425 585
R124 B.n424 B.n85 585
R125 B.n423 B.n422 585
R126 B.n421 B.n86 585
R127 B.n420 B.n419 585
R128 B.n418 B.n87 585
R129 B.n417 B.n416 585
R130 B.n415 B.n88 585
R131 B.n414 B.n413 585
R132 B.n412 B.n89 585
R133 B.n411 B.n410 585
R134 B.n409 B.n90 585
R135 B.n408 B.n407 585
R136 B.n406 B.n91 585
R137 B.n405 B.n404 585
R138 B.n403 B.n92 585
R139 B.n402 B.n401 585
R140 B.n400 B.n93 585
R141 B.n399 B.n398 585
R142 B.n397 B.n94 585
R143 B.n396 B.n395 585
R144 B.n394 B.n95 585
R145 B.n393 B.n392 585
R146 B.n391 B.n96 585
R147 B.n390 B.n389 585
R148 B.n388 B.n97 585
R149 B.n387 B.n386 585
R150 B.n385 B.n98 585
R151 B.n384 B.n383 585
R152 B.n382 B.n99 585
R153 B.n381 B.n380 585
R154 B.n379 B.n100 585
R155 B.n378 B.n377 585
R156 B.n376 B.n101 585
R157 B.n375 B.n374 585
R158 B.n373 B.n102 585
R159 B.n372 B.n371 585
R160 B.n370 B.n103 585
R161 B.n369 B.n368 585
R162 B.n367 B.n104 585
R163 B.n222 B.n221 585
R164 B.n223 B.n156 585
R165 B.n225 B.n224 585
R166 B.n226 B.n155 585
R167 B.n228 B.n227 585
R168 B.n229 B.n154 585
R169 B.n231 B.n230 585
R170 B.n232 B.n153 585
R171 B.n234 B.n233 585
R172 B.n235 B.n152 585
R173 B.n237 B.n236 585
R174 B.n238 B.n151 585
R175 B.n240 B.n239 585
R176 B.n241 B.n150 585
R177 B.n243 B.n242 585
R178 B.n244 B.n149 585
R179 B.n246 B.n245 585
R180 B.n247 B.n148 585
R181 B.n249 B.n248 585
R182 B.n250 B.n147 585
R183 B.n252 B.n251 585
R184 B.n253 B.n146 585
R185 B.n255 B.n254 585
R186 B.n256 B.n145 585
R187 B.n258 B.n257 585
R188 B.n259 B.n144 585
R189 B.n261 B.n260 585
R190 B.n262 B.n143 585
R191 B.n264 B.n263 585
R192 B.n265 B.n142 585
R193 B.n267 B.n266 585
R194 B.n268 B.n141 585
R195 B.n270 B.n269 585
R196 B.n271 B.n140 585
R197 B.n273 B.n272 585
R198 B.n274 B.n139 585
R199 B.n276 B.n275 585
R200 B.n277 B.n138 585
R201 B.n279 B.n278 585
R202 B.n280 B.n137 585
R203 B.n282 B.n281 585
R204 B.n283 B.n136 585
R205 B.n285 B.n284 585
R206 B.n287 B.n133 585
R207 B.n289 B.n288 585
R208 B.n290 B.n132 585
R209 B.n292 B.n291 585
R210 B.n293 B.n131 585
R211 B.n295 B.n294 585
R212 B.n296 B.n130 585
R213 B.n298 B.n297 585
R214 B.n299 B.n129 585
R215 B.n301 B.n300 585
R216 B.n303 B.n302 585
R217 B.n304 B.n125 585
R218 B.n306 B.n305 585
R219 B.n307 B.n124 585
R220 B.n309 B.n308 585
R221 B.n310 B.n123 585
R222 B.n312 B.n311 585
R223 B.n313 B.n122 585
R224 B.n315 B.n314 585
R225 B.n316 B.n121 585
R226 B.n318 B.n317 585
R227 B.n319 B.n120 585
R228 B.n321 B.n320 585
R229 B.n322 B.n119 585
R230 B.n324 B.n323 585
R231 B.n325 B.n118 585
R232 B.n327 B.n326 585
R233 B.n328 B.n117 585
R234 B.n330 B.n329 585
R235 B.n331 B.n116 585
R236 B.n333 B.n332 585
R237 B.n334 B.n115 585
R238 B.n336 B.n335 585
R239 B.n337 B.n114 585
R240 B.n339 B.n338 585
R241 B.n340 B.n113 585
R242 B.n342 B.n341 585
R243 B.n343 B.n112 585
R244 B.n345 B.n344 585
R245 B.n346 B.n111 585
R246 B.n348 B.n347 585
R247 B.n349 B.n110 585
R248 B.n351 B.n350 585
R249 B.n352 B.n109 585
R250 B.n354 B.n353 585
R251 B.n355 B.n108 585
R252 B.n357 B.n356 585
R253 B.n358 B.n107 585
R254 B.n360 B.n359 585
R255 B.n361 B.n106 585
R256 B.n363 B.n362 585
R257 B.n364 B.n105 585
R258 B.n366 B.n365 585
R259 B.n220 B.n157 585
R260 B.n219 B.n218 585
R261 B.n217 B.n158 585
R262 B.n216 B.n215 585
R263 B.n214 B.n159 585
R264 B.n213 B.n212 585
R265 B.n211 B.n160 585
R266 B.n210 B.n209 585
R267 B.n208 B.n161 585
R268 B.n207 B.n206 585
R269 B.n205 B.n162 585
R270 B.n204 B.n203 585
R271 B.n202 B.n163 585
R272 B.n201 B.n200 585
R273 B.n199 B.n164 585
R274 B.n198 B.n197 585
R275 B.n196 B.n165 585
R276 B.n195 B.n194 585
R277 B.n193 B.n166 585
R278 B.n192 B.n191 585
R279 B.n190 B.n167 585
R280 B.n189 B.n188 585
R281 B.n187 B.n168 585
R282 B.n186 B.n185 585
R283 B.n184 B.n169 585
R284 B.n183 B.n182 585
R285 B.n181 B.n170 585
R286 B.n180 B.n179 585
R287 B.n178 B.n171 585
R288 B.n177 B.n176 585
R289 B.n175 B.n172 585
R290 B.n174 B.n173 585
R291 B.n2 B.n0 585
R292 B.n661 B.n1 585
R293 B.n660 B.n659 585
R294 B.n658 B.n3 585
R295 B.n657 B.n656 585
R296 B.n655 B.n4 585
R297 B.n654 B.n653 585
R298 B.n652 B.n5 585
R299 B.n651 B.n650 585
R300 B.n649 B.n6 585
R301 B.n648 B.n647 585
R302 B.n646 B.n7 585
R303 B.n645 B.n644 585
R304 B.n643 B.n8 585
R305 B.n642 B.n641 585
R306 B.n640 B.n9 585
R307 B.n639 B.n638 585
R308 B.n637 B.n10 585
R309 B.n636 B.n635 585
R310 B.n634 B.n11 585
R311 B.n633 B.n632 585
R312 B.n631 B.n12 585
R313 B.n630 B.n629 585
R314 B.n628 B.n13 585
R315 B.n627 B.n626 585
R316 B.n625 B.n14 585
R317 B.n624 B.n623 585
R318 B.n622 B.n15 585
R319 B.n621 B.n620 585
R320 B.n619 B.n16 585
R321 B.n618 B.n617 585
R322 B.n616 B.n17 585
R323 B.n615 B.n614 585
R324 B.n613 B.n18 585
R325 B.n663 B.n662 585
R326 B.n222 B.n157 511.721
R327 B.n613 B.n612 511.721
R328 B.n367 B.n366 511.721
R329 B.n468 B.n71 511.721
R330 B.n126 B.t9 480.099
R331 B.n134 B.t6 480.099
R332 B.n40 B.t3 480.099
R333 B.n48 B.t0 480.099
R334 B.n218 B.n157 163.367
R335 B.n218 B.n217 163.367
R336 B.n217 B.n216 163.367
R337 B.n216 B.n159 163.367
R338 B.n212 B.n159 163.367
R339 B.n212 B.n211 163.367
R340 B.n211 B.n210 163.367
R341 B.n210 B.n161 163.367
R342 B.n206 B.n161 163.367
R343 B.n206 B.n205 163.367
R344 B.n205 B.n204 163.367
R345 B.n204 B.n163 163.367
R346 B.n200 B.n163 163.367
R347 B.n200 B.n199 163.367
R348 B.n199 B.n198 163.367
R349 B.n198 B.n165 163.367
R350 B.n194 B.n165 163.367
R351 B.n194 B.n193 163.367
R352 B.n193 B.n192 163.367
R353 B.n192 B.n167 163.367
R354 B.n188 B.n167 163.367
R355 B.n188 B.n187 163.367
R356 B.n187 B.n186 163.367
R357 B.n186 B.n169 163.367
R358 B.n182 B.n169 163.367
R359 B.n182 B.n181 163.367
R360 B.n181 B.n180 163.367
R361 B.n180 B.n171 163.367
R362 B.n176 B.n171 163.367
R363 B.n176 B.n175 163.367
R364 B.n175 B.n174 163.367
R365 B.n174 B.n2 163.367
R366 B.n662 B.n2 163.367
R367 B.n662 B.n661 163.367
R368 B.n661 B.n660 163.367
R369 B.n660 B.n3 163.367
R370 B.n656 B.n3 163.367
R371 B.n656 B.n655 163.367
R372 B.n655 B.n654 163.367
R373 B.n654 B.n5 163.367
R374 B.n650 B.n5 163.367
R375 B.n650 B.n649 163.367
R376 B.n649 B.n648 163.367
R377 B.n648 B.n7 163.367
R378 B.n644 B.n7 163.367
R379 B.n644 B.n643 163.367
R380 B.n643 B.n642 163.367
R381 B.n642 B.n9 163.367
R382 B.n638 B.n9 163.367
R383 B.n638 B.n637 163.367
R384 B.n637 B.n636 163.367
R385 B.n636 B.n11 163.367
R386 B.n632 B.n11 163.367
R387 B.n632 B.n631 163.367
R388 B.n631 B.n630 163.367
R389 B.n630 B.n13 163.367
R390 B.n626 B.n13 163.367
R391 B.n626 B.n625 163.367
R392 B.n625 B.n624 163.367
R393 B.n624 B.n15 163.367
R394 B.n620 B.n15 163.367
R395 B.n620 B.n619 163.367
R396 B.n619 B.n618 163.367
R397 B.n618 B.n17 163.367
R398 B.n614 B.n17 163.367
R399 B.n614 B.n613 163.367
R400 B.n223 B.n222 163.367
R401 B.n224 B.n223 163.367
R402 B.n224 B.n155 163.367
R403 B.n228 B.n155 163.367
R404 B.n229 B.n228 163.367
R405 B.n230 B.n229 163.367
R406 B.n230 B.n153 163.367
R407 B.n234 B.n153 163.367
R408 B.n235 B.n234 163.367
R409 B.n236 B.n235 163.367
R410 B.n236 B.n151 163.367
R411 B.n240 B.n151 163.367
R412 B.n241 B.n240 163.367
R413 B.n242 B.n241 163.367
R414 B.n242 B.n149 163.367
R415 B.n246 B.n149 163.367
R416 B.n247 B.n246 163.367
R417 B.n248 B.n247 163.367
R418 B.n248 B.n147 163.367
R419 B.n252 B.n147 163.367
R420 B.n253 B.n252 163.367
R421 B.n254 B.n253 163.367
R422 B.n254 B.n145 163.367
R423 B.n258 B.n145 163.367
R424 B.n259 B.n258 163.367
R425 B.n260 B.n259 163.367
R426 B.n260 B.n143 163.367
R427 B.n264 B.n143 163.367
R428 B.n265 B.n264 163.367
R429 B.n266 B.n265 163.367
R430 B.n266 B.n141 163.367
R431 B.n270 B.n141 163.367
R432 B.n271 B.n270 163.367
R433 B.n272 B.n271 163.367
R434 B.n272 B.n139 163.367
R435 B.n276 B.n139 163.367
R436 B.n277 B.n276 163.367
R437 B.n278 B.n277 163.367
R438 B.n278 B.n137 163.367
R439 B.n282 B.n137 163.367
R440 B.n283 B.n282 163.367
R441 B.n284 B.n283 163.367
R442 B.n284 B.n133 163.367
R443 B.n289 B.n133 163.367
R444 B.n290 B.n289 163.367
R445 B.n291 B.n290 163.367
R446 B.n291 B.n131 163.367
R447 B.n295 B.n131 163.367
R448 B.n296 B.n295 163.367
R449 B.n297 B.n296 163.367
R450 B.n297 B.n129 163.367
R451 B.n301 B.n129 163.367
R452 B.n302 B.n301 163.367
R453 B.n302 B.n125 163.367
R454 B.n306 B.n125 163.367
R455 B.n307 B.n306 163.367
R456 B.n308 B.n307 163.367
R457 B.n308 B.n123 163.367
R458 B.n312 B.n123 163.367
R459 B.n313 B.n312 163.367
R460 B.n314 B.n313 163.367
R461 B.n314 B.n121 163.367
R462 B.n318 B.n121 163.367
R463 B.n319 B.n318 163.367
R464 B.n320 B.n319 163.367
R465 B.n320 B.n119 163.367
R466 B.n324 B.n119 163.367
R467 B.n325 B.n324 163.367
R468 B.n326 B.n325 163.367
R469 B.n326 B.n117 163.367
R470 B.n330 B.n117 163.367
R471 B.n331 B.n330 163.367
R472 B.n332 B.n331 163.367
R473 B.n332 B.n115 163.367
R474 B.n336 B.n115 163.367
R475 B.n337 B.n336 163.367
R476 B.n338 B.n337 163.367
R477 B.n338 B.n113 163.367
R478 B.n342 B.n113 163.367
R479 B.n343 B.n342 163.367
R480 B.n344 B.n343 163.367
R481 B.n344 B.n111 163.367
R482 B.n348 B.n111 163.367
R483 B.n349 B.n348 163.367
R484 B.n350 B.n349 163.367
R485 B.n350 B.n109 163.367
R486 B.n354 B.n109 163.367
R487 B.n355 B.n354 163.367
R488 B.n356 B.n355 163.367
R489 B.n356 B.n107 163.367
R490 B.n360 B.n107 163.367
R491 B.n361 B.n360 163.367
R492 B.n362 B.n361 163.367
R493 B.n362 B.n105 163.367
R494 B.n366 B.n105 163.367
R495 B.n368 B.n367 163.367
R496 B.n368 B.n103 163.367
R497 B.n372 B.n103 163.367
R498 B.n373 B.n372 163.367
R499 B.n374 B.n373 163.367
R500 B.n374 B.n101 163.367
R501 B.n378 B.n101 163.367
R502 B.n379 B.n378 163.367
R503 B.n380 B.n379 163.367
R504 B.n380 B.n99 163.367
R505 B.n384 B.n99 163.367
R506 B.n385 B.n384 163.367
R507 B.n386 B.n385 163.367
R508 B.n386 B.n97 163.367
R509 B.n390 B.n97 163.367
R510 B.n391 B.n390 163.367
R511 B.n392 B.n391 163.367
R512 B.n392 B.n95 163.367
R513 B.n396 B.n95 163.367
R514 B.n397 B.n396 163.367
R515 B.n398 B.n397 163.367
R516 B.n398 B.n93 163.367
R517 B.n402 B.n93 163.367
R518 B.n403 B.n402 163.367
R519 B.n404 B.n403 163.367
R520 B.n404 B.n91 163.367
R521 B.n408 B.n91 163.367
R522 B.n409 B.n408 163.367
R523 B.n410 B.n409 163.367
R524 B.n410 B.n89 163.367
R525 B.n414 B.n89 163.367
R526 B.n415 B.n414 163.367
R527 B.n416 B.n415 163.367
R528 B.n416 B.n87 163.367
R529 B.n420 B.n87 163.367
R530 B.n421 B.n420 163.367
R531 B.n422 B.n421 163.367
R532 B.n422 B.n85 163.367
R533 B.n426 B.n85 163.367
R534 B.n427 B.n426 163.367
R535 B.n428 B.n427 163.367
R536 B.n428 B.n83 163.367
R537 B.n432 B.n83 163.367
R538 B.n433 B.n432 163.367
R539 B.n434 B.n433 163.367
R540 B.n434 B.n81 163.367
R541 B.n438 B.n81 163.367
R542 B.n439 B.n438 163.367
R543 B.n440 B.n439 163.367
R544 B.n440 B.n79 163.367
R545 B.n444 B.n79 163.367
R546 B.n445 B.n444 163.367
R547 B.n446 B.n445 163.367
R548 B.n446 B.n77 163.367
R549 B.n450 B.n77 163.367
R550 B.n451 B.n450 163.367
R551 B.n452 B.n451 163.367
R552 B.n452 B.n75 163.367
R553 B.n456 B.n75 163.367
R554 B.n457 B.n456 163.367
R555 B.n458 B.n457 163.367
R556 B.n458 B.n73 163.367
R557 B.n462 B.n73 163.367
R558 B.n463 B.n462 163.367
R559 B.n464 B.n463 163.367
R560 B.n464 B.n71 163.367
R561 B.n612 B.n19 163.367
R562 B.n608 B.n19 163.367
R563 B.n608 B.n607 163.367
R564 B.n607 B.n606 163.367
R565 B.n606 B.n21 163.367
R566 B.n602 B.n21 163.367
R567 B.n602 B.n601 163.367
R568 B.n601 B.n600 163.367
R569 B.n600 B.n23 163.367
R570 B.n596 B.n23 163.367
R571 B.n596 B.n595 163.367
R572 B.n595 B.n594 163.367
R573 B.n594 B.n25 163.367
R574 B.n590 B.n25 163.367
R575 B.n590 B.n589 163.367
R576 B.n589 B.n588 163.367
R577 B.n588 B.n27 163.367
R578 B.n584 B.n27 163.367
R579 B.n584 B.n583 163.367
R580 B.n583 B.n582 163.367
R581 B.n582 B.n29 163.367
R582 B.n578 B.n29 163.367
R583 B.n578 B.n577 163.367
R584 B.n577 B.n576 163.367
R585 B.n576 B.n31 163.367
R586 B.n572 B.n31 163.367
R587 B.n572 B.n571 163.367
R588 B.n571 B.n570 163.367
R589 B.n570 B.n33 163.367
R590 B.n566 B.n33 163.367
R591 B.n566 B.n565 163.367
R592 B.n565 B.n564 163.367
R593 B.n564 B.n35 163.367
R594 B.n560 B.n35 163.367
R595 B.n560 B.n559 163.367
R596 B.n559 B.n558 163.367
R597 B.n558 B.n37 163.367
R598 B.n554 B.n37 163.367
R599 B.n554 B.n553 163.367
R600 B.n553 B.n552 163.367
R601 B.n552 B.n39 163.367
R602 B.n548 B.n39 163.367
R603 B.n548 B.n547 163.367
R604 B.n547 B.n43 163.367
R605 B.n543 B.n43 163.367
R606 B.n543 B.n542 163.367
R607 B.n542 B.n541 163.367
R608 B.n541 B.n45 163.367
R609 B.n537 B.n45 163.367
R610 B.n537 B.n536 163.367
R611 B.n536 B.n535 163.367
R612 B.n535 B.n47 163.367
R613 B.n530 B.n47 163.367
R614 B.n530 B.n529 163.367
R615 B.n529 B.n528 163.367
R616 B.n528 B.n51 163.367
R617 B.n524 B.n51 163.367
R618 B.n524 B.n523 163.367
R619 B.n523 B.n522 163.367
R620 B.n522 B.n53 163.367
R621 B.n518 B.n53 163.367
R622 B.n518 B.n517 163.367
R623 B.n517 B.n516 163.367
R624 B.n516 B.n55 163.367
R625 B.n512 B.n55 163.367
R626 B.n512 B.n511 163.367
R627 B.n511 B.n510 163.367
R628 B.n510 B.n57 163.367
R629 B.n506 B.n57 163.367
R630 B.n506 B.n505 163.367
R631 B.n505 B.n504 163.367
R632 B.n504 B.n59 163.367
R633 B.n500 B.n59 163.367
R634 B.n500 B.n499 163.367
R635 B.n499 B.n498 163.367
R636 B.n498 B.n61 163.367
R637 B.n494 B.n61 163.367
R638 B.n494 B.n493 163.367
R639 B.n493 B.n492 163.367
R640 B.n492 B.n63 163.367
R641 B.n488 B.n63 163.367
R642 B.n488 B.n487 163.367
R643 B.n487 B.n486 163.367
R644 B.n486 B.n65 163.367
R645 B.n482 B.n65 163.367
R646 B.n482 B.n481 163.367
R647 B.n481 B.n480 163.367
R648 B.n480 B.n67 163.367
R649 B.n476 B.n67 163.367
R650 B.n476 B.n475 163.367
R651 B.n475 B.n474 163.367
R652 B.n474 B.n69 163.367
R653 B.n470 B.n69 163.367
R654 B.n470 B.n469 163.367
R655 B.n469 B.n468 163.367
R656 B.n126 B.t11 139.768
R657 B.n48 B.t1 139.768
R658 B.n134 B.t8 139.754
R659 B.n40 B.t4 139.754
R660 B.n127 B.t10 112.23
R661 B.n49 B.t2 112.23
R662 B.n135 B.t7 112.215
R663 B.n41 B.t5 112.215
R664 B.n128 B.n127 59.5399
R665 B.n286 B.n135 59.5399
R666 B.n42 B.n41 59.5399
R667 B.n532 B.n49 59.5399
R668 B.n611 B.n18 33.2493
R669 B.n467 B.n466 33.2493
R670 B.n365 B.n104 33.2493
R671 B.n221 B.n220 33.2493
R672 B.n127 B.n126 27.5399
R673 B.n135 B.n134 27.5399
R674 B.n41 B.n40 27.5399
R675 B.n49 B.n48 27.5399
R676 B B.n663 18.0485
R677 B.n611 B.n610 10.6151
R678 B.n610 B.n609 10.6151
R679 B.n609 B.n20 10.6151
R680 B.n605 B.n20 10.6151
R681 B.n605 B.n604 10.6151
R682 B.n604 B.n603 10.6151
R683 B.n603 B.n22 10.6151
R684 B.n599 B.n22 10.6151
R685 B.n599 B.n598 10.6151
R686 B.n598 B.n597 10.6151
R687 B.n597 B.n24 10.6151
R688 B.n593 B.n24 10.6151
R689 B.n593 B.n592 10.6151
R690 B.n592 B.n591 10.6151
R691 B.n591 B.n26 10.6151
R692 B.n587 B.n26 10.6151
R693 B.n587 B.n586 10.6151
R694 B.n586 B.n585 10.6151
R695 B.n585 B.n28 10.6151
R696 B.n581 B.n28 10.6151
R697 B.n581 B.n580 10.6151
R698 B.n580 B.n579 10.6151
R699 B.n579 B.n30 10.6151
R700 B.n575 B.n30 10.6151
R701 B.n575 B.n574 10.6151
R702 B.n574 B.n573 10.6151
R703 B.n573 B.n32 10.6151
R704 B.n569 B.n32 10.6151
R705 B.n569 B.n568 10.6151
R706 B.n568 B.n567 10.6151
R707 B.n567 B.n34 10.6151
R708 B.n563 B.n34 10.6151
R709 B.n563 B.n562 10.6151
R710 B.n562 B.n561 10.6151
R711 B.n561 B.n36 10.6151
R712 B.n557 B.n36 10.6151
R713 B.n557 B.n556 10.6151
R714 B.n556 B.n555 10.6151
R715 B.n555 B.n38 10.6151
R716 B.n551 B.n38 10.6151
R717 B.n551 B.n550 10.6151
R718 B.n550 B.n549 10.6151
R719 B.n546 B.n545 10.6151
R720 B.n545 B.n544 10.6151
R721 B.n544 B.n44 10.6151
R722 B.n540 B.n44 10.6151
R723 B.n540 B.n539 10.6151
R724 B.n539 B.n538 10.6151
R725 B.n538 B.n46 10.6151
R726 B.n534 B.n46 10.6151
R727 B.n534 B.n533 10.6151
R728 B.n531 B.n50 10.6151
R729 B.n527 B.n50 10.6151
R730 B.n527 B.n526 10.6151
R731 B.n526 B.n525 10.6151
R732 B.n525 B.n52 10.6151
R733 B.n521 B.n52 10.6151
R734 B.n521 B.n520 10.6151
R735 B.n520 B.n519 10.6151
R736 B.n519 B.n54 10.6151
R737 B.n515 B.n54 10.6151
R738 B.n515 B.n514 10.6151
R739 B.n514 B.n513 10.6151
R740 B.n513 B.n56 10.6151
R741 B.n509 B.n56 10.6151
R742 B.n509 B.n508 10.6151
R743 B.n508 B.n507 10.6151
R744 B.n507 B.n58 10.6151
R745 B.n503 B.n58 10.6151
R746 B.n503 B.n502 10.6151
R747 B.n502 B.n501 10.6151
R748 B.n501 B.n60 10.6151
R749 B.n497 B.n60 10.6151
R750 B.n497 B.n496 10.6151
R751 B.n496 B.n495 10.6151
R752 B.n495 B.n62 10.6151
R753 B.n491 B.n62 10.6151
R754 B.n491 B.n490 10.6151
R755 B.n490 B.n489 10.6151
R756 B.n489 B.n64 10.6151
R757 B.n485 B.n64 10.6151
R758 B.n485 B.n484 10.6151
R759 B.n484 B.n483 10.6151
R760 B.n483 B.n66 10.6151
R761 B.n479 B.n66 10.6151
R762 B.n479 B.n478 10.6151
R763 B.n478 B.n477 10.6151
R764 B.n477 B.n68 10.6151
R765 B.n473 B.n68 10.6151
R766 B.n473 B.n472 10.6151
R767 B.n472 B.n471 10.6151
R768 B.n471 B.n70 10.6151
R769 B.n467 B.n70 10.6151
R770 B.n369 B.n104 10.6151
R771 B.n370 B.n369 10.6151
R772 B.n371 B.n370 10.6151
R773 B.n371 B.n102 10.6151
R774 B.n375 B.n102 10.6151
R775 B.n376 B.n375 10.6151
R776 B.n377 B.n376 10.6151
R777 B.n377 B.n100 10.6151
R778 B.n381 B.n100 10.6151
R779 B.n382 B.n381 10.6151
R780 B.n383 B.n382 10.6151
R781 B.n383 B.n98 10.6151
R782 B.n387 B.n98 10.6151
R783 B.n388 B.n387 10.6151
R784 B.n389 B.n388 10.6151
R785 B.n389 B.n96 10.6151
R786 B.n393 B.n96 10.6151
R787 B.n394 B.n393 10.6151
R788 B.n395 B.n394 10.6151
R789 B.n395 B.n94 10.6151
R790 B.n399 B.n94 10.6151
R791 B.n400 B.n399 10.6151
R792 B.n401 B.n400 10.6151
R793 B.n401 B.n92 10.6151
R794 B.n405 B.n92 10.6151
R795 B.n406 B.n405 10.6151
R796 B.n407 B.n406 10.6151
R797 B.n407 B.n90 10.6151
R798 B.n411 B.n90 10.6151
R799 B.n412 B.n411 10.6151
R800 B.n413 B.n412 10.6151
R801 B.n413 B.n88 10.6151
R802 B.n417 B.n88 10.6151
R803 B.n418 B.n417 10.6151
R804 B.n419 B.n418 10.6151
R805 B.n419 B.n86 10.6151
R806 B.n423 B.n86 10.6151
R807 B.n424 B.n423 10.6151
R808 B.n425 B.n424 10.6151
R809 B.n425 B.n84 10.6151
R810 B.n429 B.n84 10.6151
R811 B.n430 B.n429 10.6151
R812 B.n431 B.n430 10.6151
R813 B.n431 B.n82 10.6151
R814 B.n435 B.n82 10.6151
R815 B.n436 B.n435 10.6151
R816 B.n437 B.n436 10.6151
R817 B.n437 B.n80 10.6151
R818 B.n441 B.n80 10.6151
R819 B.n442 B.n441 10.6151
R820 B.n443 B.n442 10.6151
R821 B.n443 B.n78 10.6151
R822 B.n447 B.n78 10.6151
R823 B.n448 B.n447 10.6151
R824 B.n449 B.n448 10.6151
R825 B.n449 B.n76 10.6151
R826 B.n453 B.n76 10.6151
R827 B.n454 B.n453 10.6151
R828 B.n455 B.n454 10.6151
R829 B.n455 B.n74 10.6151
R830 B.n459 B.n74 10.6151
R831 B.n460 B.n459 10.6151
R832 B.n461 B.n460 10.6151
R833 B.n461 B.n72 10.6151
R834 B.n465 B.n72 10.6151
R835 B.n466 B.n465 10.6151
R836 B.n221 B.n156 10.6151
R837 B.n225 B.n156 10.6151
R838 B.n226 B.n225 10.6151
R839 B.n227 B.n226 10.6151
R840 B.n227 B.n154 10.6151
R841 B.n231 B.n154 10.6151
R842 B.n232 B.n231 10.6151
R843 B.n233 B.n232 10.6151
R844 B.n233 B.n152 10.6151
R845 B.n237 B.n152 10.6151
R846 B.n238 B.n237 10.6151
R847 B.n239 B.n238 10.6151
R848 B.n239 B.n150 10.6151
R849 B.n243 B.n150 10.6151
R850 B.n244 B.n243 10.6151
R851 B.n245 B.n244 10.6151
R852 B.n245 B.n148 10.6151
R853 B.n249 B.n148 10.6151
R854 B.n250 B.n249 10.6151
R855 B.n251 B.n250 10.6151
R856 B.n251 B.n146 10.6151
R857 B.n255 B.n146 10.6151
R858 B.n256 B.n255 10.6151
R859 B.n257 B.n256 10.6151
R860 B.n257 B.n144 10.6151
R861 B.n261 B.n144 10.6151
R862 B.n262 B.n261 10.6151
R863 B.n263 B.n262 10.6151
R864 B.n263 B.n142 10.6151
R865 B.n267 B.n142 10.6151
R866 B.n268 B.n267 10.6151
R867 B.n269 B.n268 10.6151
R868 B.n269 B.n140 10.6151
R869 B.n273 B.n140 10.6151
R870 B.n274 B.n273 10.6151
R871 B.n275 B.n274 10.6151
R872 B.n275 B.n138 10.6151
R873 B.n279 B.n138 10.6151
R874 B.n280 B.n279 10.6151
R875 B.n281 B.n280 10.6151
R876 B.n281 B.n136 10.6151
R877 B.n285 B.n136 10.6151
R878 B.n288 B.n287 10.6151
R879 B.n288 B.n132 10.6151
R880 B.n292 B.n132 10.6151
R881 B.n293 B.n292 10.6151
R882 B.n294 B.n293 10.6151
R883 B.n294 B.n130 10.6151
R884 B.n298 B.n130 10.6151
R885 B.n299 B.n298 10.6151
R886 B.n300 B.n299 10.6151
R887 B.n304 B.n303 10.6151
R888 B.n305 B.n304 10.6151
R889 B.n305 B.n124 10.6151
R890 B.n309 B.n124 10.6151
R891 B.n310 B.n309 10.6151
R892 B.n311 B.n310 10.6151
R893 B.n311 B.n122 10.6151
R894 B.n315 B.n122 10.6151
R895 B.n316 B.n315 10.6151
R896 B.n317 B.n316 10.6151
R897 B.n317 B.n120 10.6151
R898 B.n321 B.n120 10.6151
R899 B.n322 B.n321 10.6151
R900 B.n323 B.n322 10.6151
R901 B.n323 B.n118 10.6151
R902 B.n327 B.n118 10.6151
R903 B.n328 B.n327 10.6151
R904 B.n329 B.n328 10.6151
R905 B.n329 B.n116 10.6151
R906 B.n333 B.n116 10.6151
R907 B.n334 B.n333 10.6151
R908 B.n335 B.n334 10.6151
R909 B.n335 B.n114 10.6151
R910 B.n339 B.n114 10.6151
R911 B.n340 B.n339 10.6151
R912 B.n341 B.n340 10.6151
R913 B.n341 B.n112 10.6151
R914 B.n345 B.n112 10.6151
R915 B.n346 B.n345 10.6151
R916 B.n347 B.n346 10.6151
R917 B.n347 B.n110 10.6151
R918 B.n351 B.n110 10.6151
R919 B.n352 B.n351 10.6151
R920 B.n353 B.n352 10.6151
R921 B.n353 B.n108 10.6151
R922 B.n357 B.n108 10.6151
R923 B.n358 B.n357 10.6151
R924 B.n359 B.n358 10.6151
R925 B.n359 B.n106 10.6151
R926 B.n363 B.n106 10.6151
R927 B.n364 B.n363 10.6151
R928 B.n365 B.n364 10.6151
R929 B.n220 B.n219 10.6151
R930 B.n219 B.n158 10.6151
R931 B.n215 B.n158 10.6151
R932 B.n215 B.n214 10.6151
R933 B.n214 B.n213 10.6151
R934 B.n213 B.n160 10.6151
R935 B.n209 B.n160 10.6151
R936 B.n209 B.n208 10.6151
R937 B.n208 B.n207 10.6151
R938 B.n207 B.n162 10.6151
R939 B.n203 B.n162 10.6151
R940 B.n203 B.n202 10.6151
R941 B.n202 B.n201 10.6151
R942 B.n201 B.n164 10.6151
R943 B.n197 B.n164 10.6151
R944 B.n197 B.n196 10.6151
R945 B.n196 B.n195 10.6151
R946 B.n195 B.n166 10.6151
R947 B.n191 B.n166 10.6151
R948 B.n191 B.n190 10.6151
R949 B.n190 B.n189 10.6151
R950 B.n189 B.n168 10.6151
R951 B.n185 B.n168 10.6151
R952 B.n185 B.n184 10.6151
R953 B.n184 B.n183 10.6151
R954 B.n183 B.n170 10.6151
R955 B.n179 B.n170 10.6151
R956 B.n179 B.n178 10.6151
R957 B.n178 B.n177 10.6151
R958 B.n177 B.n172 10.6151
R959 B.n173 B.n172 10.6151
R960 B.n173 B.n0 10.6151
R961 B.n659 B.n1 10.6151
R962 B.n659 B.n658 10.6151
R963 B.n658 B.n657 10.6151
R964 B.n657 B.n4 10.6151
R965 B.n653 B.n4 10.6151
R966 B.n653 B.n652 10.6151
R967 B.n652 B.n651 10.6151
R968 B.n651 B.n6 10.6151
R969 B.n647 B.n6 10.6151
R970 B.n647 B.n646 10.6151
R971 B.n646 B.n645 10.6151
R972 B.n645 B.n8 10.6151
R973 B.n641 B.n8 10.6151
R974 B.n641 B.n640 10.6151
R975 B.n640 B.n639 10.6151
R976 B.n639 B.n10 10.6151
R977 B.n635 B.n10 10.6151
R978 B.n635 B.n634 10.6151
R979 B.n634 B.n633 10.6151
R980 B.n633 B.n12 10.6151
R981 B.n629 B.n12 10.6151
R982 B.n629 B.n628 10.6151
R983 B.n628 B.n627 10.6151
R984 B.n627 B.n14 10.6151
R985 B.n623 B.n14 10.6151
R986 B.n623 B.n622 10.6151
R987 B.n622 B.n621 10.6151
R988 B.n621 B.n16 10.6151
R989 B.n617 B.n16 10.6151
R990 B.n617 B.n616 10.6151
R991 B.n616 B.n615 10.6151
R992 B.n615 B.n18 10.6151
R993 B.n549 B.n42 9.36635
R994 B.n532 B.n531 9.36635
R995 B.n286 B.n285 9.36635
R996 B.n303 B.n128 9.36635
R997 B.n663 B.n0 2.81026
R998 B.n663 B.n1 2.81026
R999 B.n546 B.n42 1.24928
R1000 B.n533 B.n532 1.24928
R1001 B.n287 B.n286 1.24928
R1002 B.n300 B.n128 1.24928
R1003 VN.n4 VN.t6 334.322
R1004 VN.n23 VN.t5 334.322
R1005 VN.n17 VN.t8 312.858
R1006 VN.n36 VN.t7 312.858
R1007 VN.n10 VN.t4 276.598
R1008 VN.n5 VN.t3 276.598
R1009 VN.n1 VN.t1 276.598
R1010 VN.n29 VN.t0 276.598
R1011 VN.n24 VN.t9 276.598
R1012 VN.n20 VN.t2 276.598
R1013 VN.n35 VN.n19 161.3
R1014 VN.n34 VN.n33 161.3
R1015 VN.n32 VN.n31 161.3
R1016 VN.n30 VN.n21 161.3
R1017 VN.n29 VN.n28 161.3
R1018 VN.n27 VN.n22 161.3
R1019 VN.n26 VN.n25 161.3
R1020 VN.n16 VN.n0 161.3
R1021 VN.n15 VN.n14 161.3
R1022 VN.n13 VN.n12 161.3
R1023 VN.n11 VN.n2 161.3
R1024 VN.n10 VN.n9 161.3
R1025 VN.n8 VN.n3 161.3
R1026 VN.n7 VN.n6 161.3
R1027 VN.n37 VN.n36 80.6037
R1028 VN.n18 VN.n17 80.6037
R1029 VN.n6 VN.n3 56.5193
R1030 VN.n12 VN.n11 56.5193
R1031 VN.n25 VN.n22 56.5193
R1032 VN.n31 VN.n30 56.5193
R1033 VN VN.n37 45.696
R1034 VN.n17 VN.n16 43.0884
R1035 VN.n36 VN.n35 43.0884
R1036 VN.n5 VN.n4 36.3862
R1037 VN.n24 VN.n23 36.3862
R1038 VN.n26 VN.n23 28.7416
R1039 VN.n7 VN.n4 28.7416
R1040 VN.n16 VN.n15 27.8669
R1041 VN.n35 VN.n34 27.8669
R1042 VN.n10 VN.n3 24.4675
R1043 VN.n11 VN.n10 24.4675
R1044 VN.n30 VN.n29 24.4675
R1045 VN.n29 VN.n22 24.4675
R1046 VN.n6 VN.n5 20.5528
R1047 VN.n12 VN.n1 20.5528
R1048 VN.n25 VN.n24 20.5528
R1049 VN.n31 VN.n20 20.5528
R1050 VN.n15 VN.n1 3.91522
R1051 VN.n34 VN.n20 3.91522
R1052 VN.n37 VN.n19 0.285035
R1053 VN.n18 VN.n0 0.285035
R1054 VN.n33 VN.n19 0.189894
R1055 VN.n33 VN.n32 0.189894
R1056 VN.n32 VN.n21 0.189894
R1057 VN.n28 VN.n21 0.189894
R1058 VN.n28 VN.n27 0.189894
R1059 VN.n27 VN.n26 0.189894
R1060 VN.n8 VN.n7 0.189894
R1061 VN.n9 VN.n8 0.189894
R1062 VN.n9 VN.n2 0.189894
R1063 VN.n13 VN.n2 0.189894
R1064 VN.n14 VN.n13 0.189894
R1065 VN.n14 VN.n0 0.189894
R1066 VN VN.n18 0.146778
R1067 VTAIL.n11 VTAIL.t17 59.913
R1068 VTAIL.n17 VTAIL.t15 59.9129
R1069 VTAIL.n2 VTAIL.t0 59.9129
R1070 VTAIL.n16 VTAIL.t2 59.9129
R1071 VTAIL.n15 VTAIL.n14 57.3148
R1072 VTAIL.n13 VTAIL.n12 57.3148
R1073 VTAIL.n10 VTAIL.n9 57.3148
R1074 VTAIL.n8 VTAIL.n7 57.3148
R1075 VTAIL.n19 VTAIL.n18 57.3145
R1076 VTAIL.n1 VTAIL.n0 57.3145
R1077 VTAIL.n4 VTAIL.n3 57.3145
R1078 VTAIL.n6 VTAIL.n5 57.3145
R1079 VTAIL.n8 VTAIL.n6 25.5996
R1080 VTAIL.n17 VTAIL.n16 24.3755
R1081 VTAIL.n18 VTAIL.t10 2.59882
R1082 VTAIL.n18 VTAIL.t9 2.59882
R1083 VTAIL.n0 VTAIL.t12 2.59882
R1084 VTAIL.n0 VTAIL.t14 2.59882
R1085 VTAIL.n3 VTAIL.t19 2.59882
R1086 VTAIL.n3 VTAIL.t7 2.59882
R1087 VTAIL.n5 VTAIL.t3 2.59882
R1088 VTAIL.n5 VTAIL.t5 2.59882
R1089 VTAIL.n14 VTAIL.t8 2.59882
R1090 VTAIL.n14 VTAIL.t4 2.59882
R1091 VTAIL.n12 VTAIL.t1 2.59882
R1092 VTAIL.n12 VTAIL.t6 2.59882
R1093 VTAIL.n9 VTAIL.t13 2.59882
R1094 VTAIL.n9 VTAIL.t16 2.59882
R1095 VTAIL.n7 VTAIL.t18 2.59882
R1096 VTAIL.n7 VTAIL.t11 2.59882
R1097 VTAIL.n10 VTAIL.n8 1.22464
R1098 VTAIL.n11 VTAIL.n10 1.22464
R1099 VTAIL.n15 VTAIL.n13 1.22464
R1100 VTAIL.n16 VTAIL.n15 1.22464
R1101 VTAIL.n6 VTAIL.n4 1.22464
R1102 VTAIL.n4 VTAIL.n2 1.22464
R1103 VTAIL.n19 VTAIL.n17 1.22464
R1104 VTAIL.n13 VTAIL.n11 1.0824
R1105 VTAIL.n2 VTAIL.n1 1.0824
R1106 VTAIL VTAIL.n1 0.976793
R1107 VTAIL VTAIL.n19 0.248345
R1108 VDD2.n1 VDD2.t3 77.8158
R1109 VDD2.n4 VDD2.t2 76.5918
R1110 VDD2.n3 VDD2.n2 74.8561
R1111 VDD2 VDD2.n7 74.8533
R1112 VDD2.n6 VDD2.n5 73.9936
R1113 VDD2.n1 VDD2.n0 73.9933
R1114 VDD2.n4 VDD2.n3 40.3144
R1115 VDD2.n7 VDD2.t0 2.59882
R1116 VDD2.n7 VDD2.t4 2.59882
R1117 VDD2.n5 VDD2.t7 2.59882
R1118 VDD2.n5 VDD2.t9 2.59882
R1119 VDD2.n2 VDD2.t8 2.59882
R1120 VDD2.n2 VDD2.t1 2.59882
R1121 VDD2.n0 VDD2.t6 2.59882
R1122 VDD2.n0 VDD2.t5 2.59882
R1123 VDD2.n6 VDD2.n4 1.22464
R1124 VDD2 VDD2.n6 0.364724
R1125 VDD2.n3 VDD2.n1 0.251188
R1126 VP.n10 VP.t9 334.322
R1127 VP.n5 VP.t3 312.858
R1128 VP.n41 VP.t0 312.858
R1129 VP.n23 VP.t7 312.858
R1130 VP.n34 VP.t8 276.598
R1131 VP.n29 VP.t5 276.598
R1132 VP.n1 VP.t1 276.598
R1133 VP.n16 VP.t4 276.598
R1134 VP.n7 VP.t6 276.598
R1135 VP.n11 VP.t2 276.598
R1136 VP.n13 VP.n12 161.3
R1137 VP.n14 VP.n9 161.3
R1138 VP.n16 VP.n15 161.3
R1139 VP.n17 VP.n8 161.3
R1140 VP.n19 VP.n18 161.3
R1141 VP.n21 VP.n20 161.3
R1142 VP.n22 VP.n6 161.3
R1143 VP.n40 VP.n0 161.3
R1144 VP.n39 VP.n38 161.3
R1145 VP.n37 VP.n36 161.3
R1146 VP.n35 VP.n2 161.3
R1147 VP.n34 VP.n33 161.3
R1148 VP.n32 VP.n3 161.3
R1149 VP.n31 VP.n30 161.3
R1150 VP.n28 VP.n4 161.3
R1151 VP.n27 VP.n26 161.3
R1152 VP.n24 VP.n23 80.6037
R1153 VP.n42 VP.n41 80.6037
R1154 VP.n25 VP.n5 80.6037
R1155 VP.n30 VP.n3 56.5193
R1156 VP.n36 VP.n35 56.5193
R1157 VP.n18 VP.n17 56.5193
R1158 VP.n12 VP.n9 56.5193
R1159 VP.n25 VP.n24 45.4105
R1160 VP.n27 VP.n5 43.0884
R1161 VP.n41 VP.n40 43.0884
R1162 VP.n23 VP.n22 43.0884
R1163 VP.n11 VP.n10 36.3862
R1164 VP.n13 VP.n10 28.7416
R1165 VP.n28 VP.n27 27.8669
R1166 VP.n40 VP.n39 27.8669
R1167 VP.n22 VP.n21 27.8669
R1168 VP.n34 VP.n3 24.4675
R1169 VP.n35 VP.n34 24.4675
R1170 VP.n16 VP.n9 24.4675
R1171 VP.n17 VP.n16 24.4675
R1172 VP.n30 VP.n29 20.5528
R1173 VP.n36 VP.n1 20.5528
R1174 VP.n18 VP.n7 20.5528
R1175 VP.n12 VP.n11 20.5528
R1176 VP.n29 VP.n28 3.91522
R1177 VP.n39 VP.n1 3.91522
R1178 VP.n21 VP.n7 3.91522
R1179 VP.n24 VP.n6 0.285035
R1180 VP.n26 VP.n25 0.285035
R1181 VP.n42 VP.n0 0.285035
R1182 VP.n14 VP.n13 0.189894
R1183 VP.n15 VP.n14 0.189894
R1184 VP.n15 VP.n8 0.189894
R1185 VP.n19 VP.n8 0.189894
R1186 VP.n20 VP.n19 0.189894
R1187 VP.n20 VP.n6 0.189894
R1188 VP.n26 VP.n4 0.189894
R1189 VP.n31 VP.n4 0.189894
R1190 VP.n32 VP.n31 0.189894
R1191 VP.n33 VP.n32 0.189894
R1192 VP.n33 VP.n2 0.189894
R1193 VP.n37 VP.n2 0.189894
R1194 VP.n38 VP.n37 0.189894
R1195 VP.n38 VP.n0 0.189894
R1196 VP VP.n42 0.146778
R1197 VDD1.n1 VDD1.t0 77.816
R1198 VDD1.n3 VDD1.t6 77.8158
R1199 VDD1.n5 VDD1.n4 74.8561
R1200 VDD1.n1 VDD1.n0 73.9936
R1201 VDD1.n7 VDD1.n6 73.9934
R1202 VDD1.n3 VDD1.n2 73.9933
R1203 VDD1.n7 VDD1.n5 41.5095
R1204 VDD1.n6 VDD1.t3 2.59882
R1205 VDD1.n6 VDD1.t2 2.59882
R1206 VDD1.n0 VDD1.t7 2.59882
R1207 VDD1.n0 VDD1.t5 2.59882
R1208 VDD1.n4 VDD1.t8 2.59882
R1209 VDD1.n4 VDD1.t9 2.59882
R1210 VDD1.n2 VDD1.t4 2.59882
R1211 VDD1.n2 VDD1.t1 2.59882
R1212 VDD1 VDD1.n7 0.860414
R1213 VDD1 VDD1.n1 0.364724
R1214 VDD1.n5 VDD1.n3 0.251188
C0 B w_n2674_n3470# 8.15036f
C1 VP B 1.47405f
C2 B VDD1 1.90891f
C3 VN B 0.904798f
C4 VTAIL B 3.07856f
C5 VDD2 B 1.96816f
C6 VP w_n2674_n3470# 5.61415f
C7 w_n2674_n3470# VDD1 2.2441f
C8 VP VDD1 8.80179f
C9 VN w_n2674_n3470# 5.27066f
C10 VN VP 6.26855f
C11 VTAIL w_n2674_n3470# 3.1193f
C12 VTAIL VP 8.57104f
C13 VDD2 w_n2674_n3470# 2.30914f
C14 VDD2 VP 0.391305f
C15 VN VDD1 0.149972f
C16 VTAIL VDD1 12.3309f
C17 VDD2 VDD1 1.21893f
C18 VTAIL VN 8.55653f
C19 VDD2 VN 8.56494f
C20 VDD2 VTAIL 12.368799f
C21 VDD2 VSUBS 1.558439f
C22 VDD1 VSUBS 1.323602f
C23 VTAIL VSUBS 0.925557f
C24 VN VSUBS 5.44368f
C25 VP VSUBS 2.350564f
C26 B VSUBS 3.535752f
C27 w_n2674_n3470# VSUBS 0.114137p
C28 VDD1.t0 VSUBS 2.6045f
C29 VDD1.t7 VSUBS 0.25266f
C30 VDD1.t5 VSUBS 0.25266f
C31 VDD1.n0 VSUBS 1.98701f
C32 VDD1.n1 VSUBS 1.27774f
C33 VDD1.t6 VSUBS 2.60449f
C34 VDD1.t4 VSUBS 0.25266f
C35 VDD1.t1 VSUBS 0.25266f
C36 VDD1.n2 VSUBS 1.98701f
C37 VDD1.n3 VSUBS 1.27077f
C38 VDD1.t8 VSUBS 0.25266f
C39 VDD1.t9 VSUBS 0.25266f
C40 VDD1.n4 VSUBS 1.99467f
C41 VDD1.n5 VSUBS 2.5479f
C42 VDD1.t3 VSUBS 0.25266f
C43 VDD1.t2 VSUBS 0.25266f
C44 VDD1.n6 VSUBS 1.98701f
C45 VDD1.n7 VSUBS 2.91681f
C46 VP.n0 VSUBS 0.059099f
C47 VP.t1 VSUBS 1.64741f
C48 VP.n1 VSUBS 0.604923f
C49 VP.n2 VSUBS 0.04429f
C50 VP.t8 VSUBS 1.64741f
C51 VP.n3 VSUBS 0.059719f
C52 VP.n4 VSUBS 0.04429f
C53 VP.t5 VSUBS 1.64741f
C54 VP.t3 VSUBS 1.72137f
C55 VP.n5 VSUBS 0.678027f
C56 VP.n6 VSUBS 0.059099f
C57 VP.t7 VSUBS 1.72137f
C58 VP.t6 VSUBS 1.64741f
C59 VP.n7 VSUBS 0.604923f
C60 VP.n8 VSUBS 0.04429f
C61 VP.t4 VSUBS 1.64741f
C62 VP.n9 VSUBS 0.059719f
C63 VP.t9 VSUBS 1.76555f
C64 VP.n10 VSUBS 0.665964f
C65 VP.t2 VSUBS 1.64741f
C66 VP.n11 VSUBS 0.669241f
C67 VP.n12 VSUBS 0.063072f
C68 VP.n13 VSUBS 0.22675f
C69 VP.n14 VSUBS 0.04429f
C70 VP.n15 VSUBS 0.04429f
C71 VP.n16 VSUBS 0.646715f
C72 VP.n17 VSUBS 0.059719f
C73 VP.n18 VSUBS 0.063072f
C74 VP.n19 VSUBS 0.04429f
C75 VP.n20 VSUBS 0.04429f
C76 VP.n21 VSUBS 0.052586f
C77 VP.n22 VSUBS 0.041777f
C78 VP.n23 VSUBS 0.678027f
C79 VP.n24 VSUBS 2.0912f
C80 VP.n25 VSUBS 2.12626f
C81 VP.n26 VSUBS 0.059099f
C82 VP.n27 VSUBS 0.041777f
C83 VP.n28 VSUBS 0.052586f
C84 VP.n29 VSUBS 0.604923f
C85 VP.n30 VSUBS 0.063072f
C86 VP.n31 VSUBS 0.04429f
C87 VP.n32 VSUBS 0.04429f
C88 VP.n33 VSUBS 0.04429f
C89 VP.n34 VSUBS 0.646715f
C90 VP.n35 VSUBS 0.059719f
C91 VP.n36 VSUBS 0.063072f
C92 VP.n37 VSUBS 0.04429f
C93 VP.n38 VSUBS 0.04429f
C94 VP.n39 VSUBS 0.052586f
C95 VP.n40 VSUBS 0.041777f
C96 VP.t0 VSUBS 1.72137f
C97 VP.n41 VSUBS 0.678027f
C98 VP.n42 VSUBS 0.041479f
C99 VDD2.t3 VSUBS 2.61509f
C100 VDD2.t6 VSUBS 0.253688f
C101 VDD2.t5 VSUBS 0.253688f
C102 VDD2.n0 VSUBS 1.99509f
C103 VDD2.n1 VSUBS 1.27594f
C104 VDD2.t8 VSUBS 0.253688f
C105 VDD2.t1 VSUBS 0.253688f
C106 VDD2.n2 VSUBS 2.00279f
C107 VDD2.n3 VSUBS 2.46945f
C108 VDD2.t2 VSUBS 2.60443f
C109 VDD2.n4 VSUBS 2.93413f
C110 VDD2.t7 VSUBS 0.253688f
C111 VDD2.t9 VSUBS 0.253688f
C112 VDD2.n5 VSUBS 1.9951f
C113 VDD2.n6 VSUBS 0.61542f
C114 VDD2.t0 VSUBS 0.253688f
C115 VDD2.t4 VSUBS 0.253688f
C116 VDD2.n7 VSUBS 2.00275f
C117 VTAIL.t12 VSUBS 0.279204f
C118 VTAIL.t14 VSUBS 0.279204f
C119 VTAIL.n0 VSUBS 2.04228f
C120 VTAIL.n1 VSUBS 0.835172f
C121 VTAIL.t0 VSUBS 2.69426f
C122 VTAIL.n2 VSUBS 0.967218f
C123 VTAIL.t19 VSUBS 0.279204f
C124 VTAIL.t7 VSUBS 0.279204f
C125 VTAIL.n3 VSUBS 2.04228f
C126 VTAIL.n4 VSUBS 0.870672f
C127 VTAIL.t3 VSUBS 0.279204f
C128 VTAIL.t5 VSUBS 0.279204f
C129 VTAIL.n5 VSUBS 2.04228f
C130 VTAIL.n6 VSUBS 2.34717f
C131 VTAIL.t18 VSUBS 0.279204f
C132 VTAIL.t11 VSUBS 0.279204f
C133 VTAIL.n7 VSUBS 2.04229f
C134 VTAIL.n8 VSUBS 2.34716f
C135 VTAIL.t13 VSUBS 0.279204f
C136 VTAIL.t16 VSUBS 0.279204f
C137 VTAIL.n9 VSUBS 2.04229f
C138 VTAIL.n10 VSUBS 0.870664f
C139 VTAIL.t17 VSUBS 2.69428f
C140 VTAIL.n11 VSUBS 0.9672f
C141 VTAIL.t1 VSUBS 0.279204f
C142 VTAIL.t6 VSUBS 0.279204f
C143 VTAIL.n12 VSUBS 2.04229f
C144 VTAIL.n13 VSUBS 0.857719f
C145 VTAIL.t8 VSUBS 0.279204f
C146 VTAIL.t4 VSUBS 0.279204f
C147 VTAIL.n14 VSUBS 2.04229f
C148 VTAIL.n15 VSUBS 0.870664f
C149 VTAIL.t2 VSUBS 2.69426f
C150 VTAIL.n16 VSUBS 2.34526f
C151 VTAIL.t15 VSUBS 2.69426f
C152 VTAIL.n17 VSUBS 2.34526f
C153 VTAIL.t10 VSUBS 0.279204f
C154 VTAIL.t9 VSUBS 0.279204f
C155 VTAIL.n18 VSUBS 2.04228f
C156 VTAIL.n19 VSUBS 0.781824f
C157 VN.n0 VSUBS 0.057968f
C158 VN.t1 VSUBS 1.61586f
C159 VN.n1 VSUBS 0.593339f
C160 VN.n2 VSUBS 0.043442f
C161 VN.t4 VSUBS 1.61586f
C162 VN.n3 VSUBS 0.058575f
C163 VN.t6 VSUBS 1.73174f
C164 VN.n4 VSUBS 0.653212f
C165 VN.t3 VSUBS 1.61586f
C166 VN.n5 VSUBS 0.656426f
C167 VN.n6 VSUBS 0.061864f
C168 VN.n7 VSUBS 0.222408f
C169 VN.n8 VSUBS 0.043442f
C170 VN.n9 VSUBS 0.043442f
C171 VN.n10 VSUBS 0.634331f
C172 VN.n11 VSUBS 0.058575f
C173 VN.n12 VSUBS 0.061864f
C174 VN.n13 VSUBS 0.043442f
C175 VN.n14 VSUBS 0.043442f
C176 VN.n15 VSUBS 0.051579f
C177 VN.n16 VSUBS 0.040977f
C178 VN.t8 VSUBS 1.68841f
C179 VN.n17 VSUBS 0.665044f
C180 VN.n18 VSUBS 0.040685f
C181 VN.n19 VSUBS 0.057968f
C182 VN.t2 VSUBS 1.61586f
C183 VN.n20 VSUBS 0.593339f
C184 VN.n21 VSUBS 0.043442f
C185 VN.t0 VSUBS 1.61586f
C186 VN.n22 VSUBS 0.058575f
C187 VN.t5 VSUBS 1.73174f
C188 VN.n23 VSUBS 0.653212f
C189 VN.t9 VSUBS 1.61586f
C190 VN.n24 VSUBS 0.656426f
C191 VN.n25 VSUBS 0.061864f
C192 VN.n26 VSUBS 0.222408f
C193 VN.n27 VSUBS 0.043442f
C194 VN.n28 VSUBS 0.043442f
C195 VN.n29 VSUBS 0.634331f
C196 VN.n30 VSUBS 0.058575f
C197 VN.n31 VSUBS 0.061864f
C198 VN.n32 VSUBS 0.043442f
C199 VN.n33 VSUBS 0.043442f
C200 VN.n34 VSUBS 0.051579f
C201 VN.n35 VSUBS 0.040977f
C202 VN.t7 VSUBS 1.68841f
C203 VN.n36 VSUBS 0.665044f
C204 VN.n37 VSUBS 2.07521f
C205 B.n0 VSUBS 0.004407f
C206 B.n1 VSUBS 0.004407f
C207 B.n2 VSUBS 0.00697f
C208 B.n3 VSUBS 0.00697f
C209 B.n4 VSUBS 0.00697f
C210 B.n5 VSUBS 0.00697f
C211 B.n6 VSUBS 0.00697f
C212 B.n7 VSUBS 0.00697f
C213 B.n8 VSUBS 0.00697f
C214 B.n9 VSUBS 0.00697f
C215 B.n10 VSUBS 0.00697f
C216 B.n11 VSUBS 0.00697f
C217 B.n12 VSUBS 0.00697f
C218 B.n13 VSUBS 0.00697f
C219 B.n14 VSUBS 0.00697f
C220 B.n15 VSUBS 0.00697f
C221 B.n16 VSUBS 0.00697f
C222 B.n17 VSUBS 0.00697f
C223 B.n18 VSUBS 0.01594f
C224 B.n19 VSUBS 0.00697f
C225 B.n20 VSUBS 0.00697f
C226 B.n21 VSUBS 0.00697f
C227 B.n22 VSUBS 0.00697f
C228 B.n23 VSUBS 0.00697f
C229 B.n24 VSUBS 0.00697f
C230 B.n25 VSUBS 0.00697f
C231 B.n26 VSUBS 0.00697f
C232 B.n27 VSUBS 0.00697f
C233 B.n28 VSUBS 0.00697f
C234 B.n29 VSUBS 0.00697f
C235 B.n30 VSUBS 0.00697f
C236 B.n31 VSUBS 0.00697f
C237 B.n32 VSUBS 0.00697f
C238 B.n33 VSUBS 0.00697f
C239 B.n34 VSUBS 0.00697f
C240 B.n35 VSUBS 0.00697f
C241 B.n36 VSUBS 0.00697f
C242 B.n37 VSUBS 0.00697f
C243 B.n38 VSUBS 0.00697f
C244 B.n39 VSUBS 0.00697f
C245 B.t5 VSUBS 0.407711f
C246 B.t4 VSUBS 0.418617f
C247 B.t3 VSUBS 0.577383f
C248 B.n40 VSUBS 0.165997f
C249 B.n41 VSUBS 0.065286f
C250 B.n42 VSUBS 0.016148f
C251 B.n43 VSUBS 0.00697f
C252 B.n44 VSUBS 0.00697f
C253 B.n45 VSUBS 0.00697f
C254 B.n46 VSUBS 0.00697f
C255 B.n47 VSUBS 0.00697f
C256 B.t2 VSUBS 0.407703f
C257 B.t1 VSUBS 0.418609f
C258 B.t0 VSUBS 0.577383f
C259 B.n48 VSUBS 0.166005f
C260 B.n49 VSUBS 0.065294f
C261 B.n50 VSUBS 0.00697f
C262 B.n51 VSUBS 0.00697f
C263 B.n52 VSUBS 0.00697f
C264 B.n53 VSUBS 0.00697f
C265 B.n54 VSUBS 0.00697f
C266 B.n55 VSUBS 0.00697f
C267 B.n56 VSUBS 0.00697f
C268 B.n57 VSUBS 0.00697f
C269 B.n58 VSUBS 0.00697f
C270 B.n59 VSUBS 0.00697f
C271 B.n60 VSUBS 0.00697f
C272 B.n61 VSUBS 0.00697f
C273 B.n62 VSUBS 0.00697f
C274 B.n63 VSUBS 0.00697f
C275 B.n64 VSUBS 0.00697f
C276 B.n65 VSUBS 0.00697f
C277 B.n66 VSUBS 0.00697f
C278 B.n67 VSUBS 0.00697f
C279 B.n68 VSUBS 0.00697f
C280 B.n69 VSUBS 0.00697f
C281 B.n70 VSUBS 0.00697f
C282 B.n71 VSUBS 0.01594f
C283 B.n72 VSUBS 0.00697f
C284 B.n73 VSUBS 0.00697f
C285 B.n74 VSUBS 0.00697f
C286 B.n75 VSUBS 0.00697f
C287 B.n76 VSUBS 0.00697f
C288 B.n77 VSUBS 0.00697f
C289 B.n78 VSUBS 0.00697f
C290 B.n79 VSUBS 0.00697f
C291 B.n80 VSUBS 0.00697f
C292 B.n81 VSUBS 0.00697f
C293 B.n82 VSUBS 0.00697f
C294 B.n83 VSUBS 0.00697f
C295 B.n84 VSUBS 0.00697f
C296 B.n85 VSUBS 0.00697f
C297 B.n86 VSUBS 0.00697f
C298 B.n87 VSUBS 0.00697f
C299 B.n88 VSUBS 0.00697f
C300 B.n89 VSUBS 0.00697f
C301 B.n90 VSUBS 0.00697f
C302 B.n91 VSUBS 0.00697f
C303 B.n92 VSUBS 0.00697f
C304 B.n93 VSUBS 0.00697f
C305 B.n94 VSUBS 0.00697f
C306 B.n95 VSUBS 0.00697f
C307 B.n96 VSUBS 0.00697f
C308 B.n97 VSUBS 0.00697f
C309 B.n98 VSUBS 0.00697f
C310 B.n99 VSUBS 0.00697f
C311 B.n100 VSUBS 0.00697f
C312 B.n101 VSUBS 0.00697f
C313 B.n102 VSUBS 0.00697f
C314 B.n103 VSUBS 0.00697f
C315 B.n104 VSUBS 0.01594f
C316 B.n105 VSUBS 0.00697f
C317 B.n106 VSUBS 0.00697f
C318 B.n107 VSUBS 0.00697f
C319 B.n108 VSUBS 0.00697f
C320 B.n109 VSUBS 0.00697f
C321 B.n110 VSUBS 0.00697f
C322 B.n111 VSUBS 0.00697f
C323 B.n112 VSUBS 0.00697f
C324 B.n113 VSUBS 0.00697f
C325 B.n114 VSUBS 0.00697f
C326 B.n115 VSUBS 0.00697f
C327 B.n116 VSUBS 0.00697f
C328 B.n117 VSUBS 0.00697f
C329 B.n118 VSUBS 0.00697f
C330 B.n119 VSUBS 0.00697f
C331 B.n120 VSUBS 0.00697f
C332 B.n121 VSUBS 0.00697f
C333 B.n122 VSUBS 0.00697f
C334 B.n123 VSUBS 0.00697f
C335 B.n124 VSUBS 0.00697f
C336 B.n125 VSUBS 0.00697f
C337 B.t10 VSUBS 0.407703f
C338 B.t11 VSUBS 0.418609f
C339 B.t9 VSUBS 0.577383f
C340 B.n126 VSUBS 0.166005f
C341 B.n127 VSUBS 0.065294f
C342 B.n128 VSUBS 0.016148f
C343 B.n129 VSUBS 0.00697f
C344 B.n130 VSUBS 0.00697f
C345 B.n131 VSUBS 0.00697f
C346 B.n132 VSUBS 0.00697f
C347 B.n133 VSUBS 0.00697f
C348 B.t7 VSUBS 0.407711f
C349 B.t8 VSUBS 0.418617f
C350 B.t6 VSUBS 0.577383f
C351 B.n134 VSUBS 0.165997f
C352 B.n135 VSUBS 0.065286f
C353 B.n136 VSUBS 0.00697f
C354 B.n137 VSUBS 0.00697f
C355 B.n138 VSUBS 0.00697f
C356 B.n139 VSUBS 0.00697f
C357 B.n140 VSUBS 0.00697f
C358 B.n141 VSUBS 0.00697f
C359 B.n142 VSUBS 0.00697f
C360 B.n143 VSUBS 0.00697f
C361 B.n144 VSUBS 0.00697f
C362 B.n145 VSUBS 0.00697f
C363 B.n146 VSUBS 0.00697f
C364 B.n147 VSUBS 0.00697f
C365 B.n148 VSUBS 0.00697f
C366 B.n149 VSUBS 0.00697f
C367 B.n150 VSUBS 0.00697f
C368 B.n151 VSUBS 0.00697f
C369 B.n152 VSUBS 0.00697f
C370 B.n153 VSUBS 0.00697f
C371 B.n154 VSUBS 0.00697f
C372 B.n155 VSUBS 0.00697f
C373 B.n156 VSUBS 0.00697f
C374 B.n157 VSUBS 0.01594f
C375 B.n158 VSUBS 0.00697f
C376 B.n159 VSUBS 0.00697f
C377 B.n160 VSUBS 0.00697f
C378 B.n161 VSUBS 0.00697f
C379 B.n162 VSUBS 0.00697f
C380 B.n163 VSUBS 0.00697f
C381 B.n164 VSUBS 0.00697f
C382 B.n165 VSUBS 0.00697f
C383 B.n166 VSUBS 0.00697f
C384 B.n167 VSUBS 0.00697f
C385 B.n168 VSUBS 0.00697f
C386 B.n169 VSUBS 0.00697f
C387 B.n170 VSUBS 0.00697f
C388 B.n171 VSUBS 0.00697f
C389 B.n172 VSUBS 0.00697f
C390 B.n173 VSUBS 0.00697f
C391 B.n174 VSUBS 0.00697f
C392 B.n175 VSUBS 0.00697f
C393 B.n176 VSUBS 0.00697f
C394 B.n177 VSUBS 0.00697f
C395 B.n178 VSUBS 0.00697f
C396 B.n179 VSUBS 0.00697f
C397 B.n180 VSUBS 0.00697f
C398 B.n181 VSUBS 0.00697f
C399 B.n182 VSUBS 0.00697f
C400 B.n183 VSUBS 0.00697f
C401 B.n184 VSUBS 0.00697f
C402 B.n185 VSUBS 0.00697f
C403 B.n186 VSUBS 0.00697f
C404 B.n187 VSUBS 0.00697f
C405 B.n188 VSUBS 0.00697f
C406 B.n189 VSUBS 0.00697f
C407 B.n190 VSUBS 0.00697f
C408 B.n191 VSUBS 0.00697f
C409 B.n192 VSUBS 0.00697f
C410 B.n193 VSUBS 0.00697f
C411 B.n194 VSUBS 0.00697f
C412 B.n195 VSUBS 0.00697f
C413 B.n196 VSUBS 0.00697f
C414 B.n197 VSUBS 0.00697f
C415 B.n198 VSUBS 0.00697f
C416 B.n199 VSUBS 0.00697f
C417 B.n200 VSUBS 0.00697f
C418 B.n201 VSUBS 0.00697f
C419 B.n202 VSUBS 0.00697f
C420 B.n203 VSUBS 0.00697f
C421 B.n204 VSUBS 0.00697f
C422 B.n205 VSUBS 0.00697f
C423 B.n206 VSUBS 0.00697f
C424 B.n207 VSUBS 0.00697f
C425 B.n208 VSUBS 0.00697f
C426 B.n209 VSUBS 0.00697f
C427 B.n210 VSUBS 0.00697f
C428 B.n211 VSUBS 0.00697f
C429 B.n212 VSUBS 0.00697f
C430 B.n213 VSUBS 0.00697f
C431 B.n214 VSUBS 0.00697f
C432 B.n215 VSUBS 0.00697f
C433 B.n216 VSUBS 0.00697f
C434 B.n217 VSUBS 0.00697f
C435 B.n218 VSUBS 0.00697f
C436 B.n219 VSUBS 0.00697f
C437 B.n220 VSUBS 0.01594f
C438 B.n221 VSUBS 0.017065f
C439 B.n222 VSUBS 0.017065f
C440 B.n223 VSUBS 0.00697f
C441 B.n224 VSUBS 0.00697f
C442 B.n225 VSUBS 0.00697f
C443 B.n226 VSUBS 0.00697f
C444 B.n227 VSUBS 0.00697f
C445 B.n228 VSUBS 0.00697f
C446 B.n229 VSUBS 0.00697f
C447 B.n230 VSUBS 0.00697f
C448 B.n231 VSUBS 0.00697f
C449 B.n232 VSUBS 0.00697f
C450 B.n233 VSUBS 0.00697f
C451 B.n234 VSUBS 0.00697f
C452 B.n235 VSUBS 0.00697f
C453 B.n236 VSUBS 0.00697f
C454 B.n237 VSUBS 0.00697f
C455 B.n238 VSUBS 0.00697f
C456 B.n239 VSUBS 0.00697f
C457 B.n240 VSUBS 0.00697f
C458 B.n241 VSUBS 0.00697f
C459 B.n242 VSUBS 0.00697f
C460 B.n243 VSUBS 0.00697f
C461 B.n244 VSUBS 0.00697f
C462 B.n245 VSUBS 0.00697f
C463 B.n246 VSUBS 0.00697f
C464 B.n247 VSUBS 0.00697f
C465 B.n248 VSUBS 0.00697f
C466 B.n249 VSUBS 0.00697f
C467 B.n250 VSUBS 0.00697f
C468 B.n251 VSUBS 0.00697f
C469 B.n252 VSUBS 0.00697f
C470 B.n253 VSUBS 0.00697f
C471 B.n254 VSUBS 0.00697f
C472 B.n255 VSUBS 0.00697f
C473 B.n256 VSUBS 0.00697f
C474 B.n257 VSUBS 0.00697f
C475 B.n258 VSUBS 0.00697f
C476 B.n259 VSUBS 0.00697f
C477 B.n260 VSUBS 0.00697f
C478 B.n261 VSUBS 0.00697f
C479 B.n262 VSUBS 0.00697f
C480 B.n263 VSUBS 0.00697f
C481 B.n264 VSUBS 0.00697f
C482 B.n265 VSUBS 0.00697f
C483 B.n266 VSUBS 0.00697f
C484 B.n267 VSUBS 0.00697f
C485 B.n268 VSUBS 0.00697f
C486 B.n269 VSUBS 0.00697f
C487 B.n270 VSUBS 0.00697f
C488 B.n271 VSUBS 0.00697f
C489 B.n272 VSUBS 0.00697f
C490 B.n273 VSUBS 0.00697f
C491 B.n274 VSUBS 0.00697f
C492 B.n275 VSUBS 0.00697f
C493 B.n276 VSUBS 0.00697f
C494 B.n277 VSUBS 0.00697f
C495 B.n278 VSUBS 0.00697f
C496 B.n279 VSUBS 0.00697f
C497 B.n280 VSUBS 0.00697f
C498 B.n281 VSUBS 0.00697f
C499 B.n282 VSUBS 0.00697f
C500 B.n283 VSUBS 0.00697f
C501 B.n284 VSUBS 0.00697f
C502 B.n285 VSUBS 0.00656f
C503 B.n286 VSUBS 0.016148f
C504 B.n287 VSUBS 0.003895f
C505 B.n288 VSUBS 0.00697f
C506 B.n289 VSUBS 0.00697f
C507 B.n290 VSUBS 0.00697f
C508 B.n291 VSUBS 0.00697f
C509 B.n292 VSUBS 0.00697f
C510 B.n293 VSUBS 0.00697f
C511 B.n294 VSUBS 0.00697f
C512 B.n295 VSUBS 0.00697f
C513 B.n296 VSUBS 0.00697f
C514 B.n297 VSUBS 0.00697f
C515 B.n298 VSUBS 0.00697f
C516 B.n299 VSUBS 0.00697f
C517 B.n300 VSUBS 0.003895f
C518 B.n301 VSUBS 0.00697f
C519 B.n302 VSUBS 0.00697f
C520 B.n303 VSUBS 0.00656f
C521 B.n304 VSUBS 0.00697f
C522 B.n305 VSUBS 0.00697f
C523 B.n306 VSUBS 0.00697f
C524 B.n307 VSUBS 0.00697f
C525 B.n308 VSUBS 0.00697f
C526 B.n309 VSUBS 0.00697f
C527 B.n310 VSUBS 0.00697f
C528 B.n311 VSUBS 0.00697f
C529 B.n312 VSUBS 0.00697f
C530 B.n313 VSUBS 0.00697f
C531 B.n314 VSUBS 0.00697f
C532 B.n315 VSUBS 0.00697f
C533 B.n316 VSUBS 0.00697f
C534 B.n317 VSUBS 0.00697f
C535 B.n318 VSUBS 0.00697f
C536 B.n319 VSUBS 0.00697f
C537 B.n320 VSUBS 0.00697f
C538 B.n321 VSUBS 0.00697f
C539 B.n322 VSUBS 0.00697f
C540 B.n323 VSUBS 0.00697f
C541 B.n324 VSUBS 0.00697f
C542 B.n325 VSUBS 0.00697f
C543 B.n326 VSUBS 0.00697f
C544 B.n327 VSUBS 0.00697f
C545 B.n328 VSUBS 0.00697f
C546 B.n329 VSUBS 0.00697f
C547 B.n330 VSUBS 0.00697f
C548 B.n331 VSUBS 0.00697f
C549 B.n332 VSUBS 0.00697f
C550 B.n333 VSUBS 0.00697f
C551 B.n334 VSUBS 0.00697f
C552 B.n335 VSUBS 0.00697f
C553 B.n336 VSUBS 0.00697f
C554 B.n337 VSUBS 0.00697f
C555 B.n338 VSUBS 0.00697f
C556 B.n339 VSUBS 0.00697f
C557 B.n340 VSUBS 0.00697f
C558 B.n341 VSUBS 0.00697f
C559 B.n342 VSUBS 0.00697f
C560 B.n343 VSUBS 0.00697f
C561 B.n344 VSUBS 0.00697f
C562 B.n345 VSUBS 0.00697f
C563 B.n346 VSUBS 0.00697f
C564 B.n347 VSUBS 0.00697f
C565 B.n348 VSUBS 0.00697f
C566 B.n349 VSUBS 0.00697f
C567 B.n350 VSUBS 0.00697f
C568 B.n351 VSUBS 0.00697f
C569 B.n352 VSUBS 0.00697f
C570 B.n353 VSUBS 0.00697f
C571 B.n354 VSUBS 0.00697f
C572 B.n355 VSUBS 0.00697f
C573 B.n356 VSUBS 0.00697f
C574 B.n357 VSUBS 0.00697f
C575 B.n358 VSUBS 0.00697f
C576 B.n359 VSUBS 0.00697f
C577 B.n360 VSUBS 0.00697f
C578 B.n361 VSUBS 0.00697f
C579 B.n362 VSUBS 0.00697f
C580 B.n363 VSUBS 0.00697f
C581 B.n364 VSUBS 0.00697f
C582 B.n365 VSUBS 0.017065f
C583 B.n366 VSUBS 0.017065f
C584 B.n367 VSUBS 0.01594f
C585 B.n368 VSUBS 0.00697f
C586 B.n369 VSUBS 0.00697f
C587 B.n370 VSUBS 0.00697f
C588 B.n371 VSUBS 0.00697f
C589 B.n372 VSUBS 0.00697f
C590 B.n373 VSUBS 0.00697f
C591 B.n374 VSUBS 0.00697f
C592 B.n375 VSUBS 0.00697f
C593 B.n376 VSUBS 0.00697f
C594 B.n377 VSUBS 0.00697f
C595 B.n378 VSUBS 0.00697f
C596 B.n379 VSUBS 0.00697f
C597 B.n380 VSUBS 0.00697f
C598 B.n381 VSUBS 0.00697f
C599 B.n382 VSUBS 0.00697f
C600 B.n383 VSUBS 0.00697f
C601 B.n384 VSUBS 0.00697f
C602 B.n385 VSUBS 0.00697f
C603 B.n386 VSUBS 0.00697f
C604 B.n387 VSUBS 0.00697f
C605 B.n388 VSUBS 0.00697f
C606 B.n389 VSUBS 0.00697f
C607 B.n390 VSUBS 0.00697f
C608 B.n391 VSUBS 0.00697f
C609 B.n392 VSUBS 0.00697f
C610 B.n393 VSUBS 0.00697f
C611 B.n394 VSUBS 0.00697f
C612 B.n395 VSUBS 0.00697f
C613 B.n396 VSUBS 0.00697f
C614 B.n397 VSUBS 0.00697f
C615 B.n398 VSUBS 0.00697f
C616 B.n399 VSUBS 0.00697f
C617 B.n400 VSUBS 0.00697f
C618 B.n401 VSUBS 0.00697f
C619 B.n402 VSUBS 0.00697f
C620 B.n403 VSUBS 0.00697f
C621 B.n404 VSUBS 0.00697f
C622 B.n405 VSUBS 0.00697f
C623 B.n406 VSUBS 0.00697f
C624 B.n407 VSUBS 0.00697f
C625 B.n408 VSUBS 0.00697f
C626 B.n409 VSUBS 0.00697f
C627 B.n410 VSUBS 0.00697f
C628 B.n411 VSUBS 0.00697f
C629 B.n412 VSUBS 0.00697f
C630 B.n413 VSUBS 0.00697f
C631 B.n414 VSUBS 0.00697f
C632 B.n415 VSUBS 0.00697f
C633 B.n416 VSUBS 0.00697f
C634 B.n417 VSUBS 0.00697f
C635 B.n418 VSUBS 0.00697f
C636 B.n419 VSUBS 0.00697f
C637 B.n420 VSUBS 0.00697f
C638 B.n421 VSUBS 0.00697f
C639 B.n422 VSUBS 0.00697f
C640 B.n423 VSUBS 0.00697f
C641 B.n424 VSUBS 0.00697f
C642 B.n425 VSUBS 0.00697f
C643 B.n426 VSUBS 0.00697f
C644 B.n427 VSUBS 0.00697f
C645 B.n428 VSUBS 0.00697f
C646 B.n429 VSUBS 0.00697f
C647 B.n430 VSUBS 0.00697f
C648 B.n431 VSUBS 0.00697f
C649 B.n432 VSUBS 0.00697f
C650 B.n433 VSUBS 0.00697f
C651 B.n434 VSUBS 0.00697f
C652 B.n435 VSUBS 0.00697f
C653 B.n436 VSUBS 0.00697f
C654 B.n437 VSUBS 0.00697f
C655 B.n438 VSUBS 0.00697f
C656 B.n439 VSUBS 0.00697f
C657 B.n440 VSUBS 0.00697f
C658 B.n441 VSUBS 0.00697f
C659 B.n442 VSUBS 0.00697f
C660 B.n443 VSUBS 0.00697f
C661 B.n444 VSUBS 0.00697f
C662 B.n445 VSUBS 0.00697f
C663 B.n446 VSUBS 0.00697f
C664 B.n447 VSUBS 0.00697f
C665 B.n448 VSUBS 0.00697f
C666 B.n449 VSUBS 0.00697f
C667 B.n450 VSUBS 0.00697f
C668 B.n451 VSUBS 0.00697f
C669 B.n452 VSUBS 0.00697f
C670 B.n453 VSUBS 0.00697f
C671 B.n454 VSUBS 0.00697f
C672 B.n455 VSUBS 0.00697f
C673 B.n456 VSUBS 0.00697f
C674 B.n457 VSUBS 0.00697f
C675 B.n458 VSUBS 0.00697f
C676 B.n459 VSUBS 0.00697f
C677 B.n460 VSUBS 0.00697f
C678 B.n461 VSUBS 0.00697f
C679 B.n462 VSUBS 0.00697f
C680 B.n463 VSUBS 0.00697f
C681 B.n464 VSUBS 0.00697f
C682 B.n465 VSUBS 0.00697f
C683 B.n466 VSUBS 0.016749f
C684 B.n467 VSUBS 0.016256f
C685 B.n468 VSUBS 0.017065f
C686 B.n469 VSUBS 0.00697f
C687 B.n470 VSUBS 0.00697f
C688 B.n471 VSUBS 0.00697f
C689 B.n472 VSUBS 0.00697f
C690 B.n473 VSUBS 0.00697f
C691 B.n474 VSUBS 0.00697f
C692 B.n475 VSUBS 0.00697f
C693 B.n476 VSUBS 0.00697f
C694 B.n477 VSUBS 0.00697f
C695 B.n478 VSUBS 0.00697f
C696 B.n479 VSUBS 0.00697f
C697 B.n480 VSUBS 0.00697f
C698 B.n481 VSUBS 0.00697f
C699 B.n482 VSUBS 0.00697f
C700 B.n483 VSUBS 0.00697f
C701 B.n484 VSUBS 0.00697f
C702 B.n485 VSUBS 0.00697f
C703 B.n486 VSUBS 0.00697f
C704 B.n487 VSUBS 0.00697f
C705 B.n488 VSUBS 0.00697f
C706 B.n489 VSUBS 0.00697f
C707 B.n490 VSUBS 0.00697f
C708 B.n491 VSUBS 0.00697f
C709 B.n492 VSUBS 0.00697f
C710 B.n493 VSUBS 0.00697f
C711 B.n494 VSUBS 0.00697f
C712 B.n495 VSUBS 0.00697f
C713 B.n496 VSUBS 0.00697f
C714 B.n497 VSUBS 0.00697f
C715 B.n498 VSUBS 0.00697f
C716 B.n499 VSUBS 0.00697f
C717 B.n500 VSUBS 0.00697f
C718 B.n501 VSUBS 0.00697f
C719 B.n502 VSUBS 0.00697f
C720 B.n503 VSUBS 0.00697f
C721 B.n504 VSUBS 0.00697f
C722 B.n505 VSUBS 0.00697f
C723 B.n506 VSUBS 0.00697f
C724 B.n507 VSUBS 0.00697f
C725 B.n508 VSUBS 0.00697f
C726 B.n509 VSUBS 0.00697f
C727 B.n510 VSUBS 0.00697f
C728 B.n511 VSUBS 0.00697f
C729 B.n512 VSUBS 0.00697f
C730 B.n513 VSUBS 0.00697f
C731 B.n514 VSUBS 0.00697f
C732 B.n515 VSUBS 0.00697f
C733 B.n516 VSUBS 0.00697f
C734 B.n517 VSUBS 0.00697f
C735 B.n518 VSUBS 0.00697f
C736 B.n519 VSUBS 0.00697f
C737 B.n520 VSUBS 0.00697f
C738 B.n521 VSUBS 0.00697f
C739 B.n522 VSUBS 0.00697f
C740 B.n523 VSUBS 0.00697f
C741 B.n524 VSUBS 0.00697f
C742 B.n525 VSUBS 0.00697f
C743 B.n526 VSUBS 0.00697f
C744 B.n527 VSUBS 0.00697f
C745 B.n528 VSUBS 0.00697f
C746 B.n529 VSUBS 0.00697f
C747 B.n530 VSUBS 0.00697f
C748 B.n531 VSUBS 0.00656f
C749 B.n532 VSUBS 0.016148f
C750 B.n533 VSUBS 0.003895f
C751 B.n534 VSUBS 0.00697f
C752 B.n535 VSUBS 0.00697f
C753 B.n536 VSUBS 0.00697f
C754 B.n537 VSUBS 0.00697f
C755 B.n538 VSUBS 0.00697f
C756 B.n539 VSUBS 0.00697f
C757 B.n540 VSUBS 0.00697f
C758 B.n541 VSUBS 0.00697f
C759 B.n542 VSUBS 0.00697f
C760 B.n543 VSUBS 0.00697f
C761 B.n544 VSUBS 0.00697f
C762 B.n545 VSUBS 0.00697f
C763 B.n546 VSUBS 0.003895f
C764 B.n547 VSUBS 0.00697f
C765 B.n548 VSUBS 0.00697f
C766 B.n549 VSUBS 0.00656f
C767 B.n550 VSUBS 0.00697f
C768 B.n551 VSUBS 0.00697f
C769 B.n552 VSUBS 0.00697f
C770 B.n553 VSUBS 0.00697f
C771 B.n554 VSUBS 0.00697f
C772 B.n555 VSUBS 0.00697f
C773 B.n556 VSUBS 0.00697f
C774 B.n557 VSUBS 0.00697f
C775 B.n558 VSUBS 0.00697f
C776 B.n559 VSUBS 0.00697f
C777 B.n560 VSUBS 0.00697f
C778 B.n561 VSUBS 0.00697f
C779 B.n562 VSUBS 0.00697f
C780 B.n563 VSUBS 0.00697f
C781 B.n564 VSUBS 0.00697f
C782 B.n565 VSUBS 0.00697f
C783 B.n566 VSUBS 0.00697f
C784 B.n567 VSUBS 0.00697f
C785 B.n568 VSUBS 0.00697f
C786 B.n569 VSUBS 0.00697f
C787 B.n570 VSUBS 0.00697f
C788 B.n571 VSUBS 0.00697f
C789 B.n572 VSUBS 0.00697f
C790 B.n573 VSUBS 0.00697f
C791 B.n574 VSUBS 0.00697f
C792 B.n575 VSUBS 0.00697f
C793 B.n576 VSUBS 0.00697f
C794 B.n577 VSUBS 0.00697f
C795 B.n578 VSUBS 0.00697f
C796 B.n579 VSUBS 0.00697f
C797 B.n580 VSUBS 0.00697f
C798 B.n581 VSUBS 0.00697f
C799 B.n582 VSUBS 0.00697f
C800 B.n583 VSUBS 0.00697f
C801 B.n584 VSUBS 0.00697f
C802 B.n585 VSUBS 0.00697f
C803 B.n586 VSUBS 0.00697f
C804 B.n587 VSUBS 0.00697f
C805 B.n588 VSUBS 0.00697f
C806 B.n589 VSUBS 0.00697f
C807 B.n590 VSUBS 0.00697f
C808 B.n591 VSUBS 0.00697f
C809 B.n592 VSUBS 0.00697f
C810 B.n593 VSUBS 0.00697f
C811 B.n594 VSUBS 0.00697f
C812 B.n595 VSUBS 0.00697f
C813 B.n596 VSUBS 0.00697f
C814 B.n597 VSUBS 0.00697f
C815 B.n598 VSUBS 0.00697f
C816 B.n599 VSUBS 0.00697f
C817 B.n600 VSUBS 0.00697f
C818 B.n601 VSUBS 0.00697f
C819 B.n602 VSUBS 0.00697f
C820 B.n603 VSUBS 0.00697f
C821 B.n604 VSUBS 0.00697f
C822 B.n605 VSUBS 0.00697f
C823 B.n606 VSUBS 0.00697f
C824 B.n607 VSUBS 0.00697f
C825 B.n608 VSUBS 0.00697f
C826 B.n609 VSUBS 0.00697f
C827 B.n610 VSUBS 0.00697f
C828 B.n611 VSUBS 0.017065f
C829 B.n612 VSUBS 0.017065f
C830 B.n613 VSUBS 0.01594f
C831 B.n614 VSUBS 0.00697f
C832 B.n615 VSUBS 0.00697f
C833 B.n616 VSUBS 0.00697f
C834 B.n617 VSUBS 0.00697f
C835 B.n618 VSUBS 0.00697f
C836 B.n619 VSUBS 0.00697f
C837 B.n620 VSUBS 0.00697f
C838 B.n621 VSUBS 0.00697f
C839 B.n622 VSUBS 0.00697f
C840 B.n623 VSUBS 0.00697f
C841 B.n624 VSUBS 0.00697f
C842 B.n625 VSUBS 0.00697f
C843 B.n626 VSUBS 0.00697f
C844 B.n627 VSUBS 0.00697f
C845 B.n628 VSUBS 0.00697f
C846 B.n629 VSUBS 0.00697f
C847 B.n630 VSUBS 0.00697f
C848 B.n631 VSUBS 0.00697f
C849 B.n632 VSUBS 0.00697f
C850 B.n633 VSUBS 0.00697f
C851 B.n634 VSUBS 0.00697f
C852 B.n635 VSUBS 0.00697f
C853 B.n636 VSUBS 0.00697f
C854 B.n637 VSUBS 0.00697f
C855 B.n638 VSUBS 0.00697f
C856 B.n639 VSUBS 0.00697f
C857 B.n640 VSUBS 0.00697f
C858 B.n641 VSUBS 0.00697f
C859 B.n642 VSUBS 0.00697f
C860 B.n643 VSUBS 0.00697f
C861 B.n644 VSUBS 0.00697f
C862 B.n645 VSUBS 0.00697f
C863 B.n646 VSUBS 0.00697f
C864 B.n647 VSUBS 0.00697f
C865 B.n648 VSUBS 0.00697f
C866 B.n649 VSUBS 0.00697f
C867 B.n650 VSUBS 0.00697f
C868 B.n651 VSUBS 0.00697f
C869 B.n652 VSUBS 0.00697f
C870 B.n653 VSUBS 0.00697f
C871 B.n654 VSUBS 0.00697f
C872 B.n655 VSUBS 0.00697f
C873 B.n656 VSUBS 0.00697f
C874 B.n657 VSUBS 0.00697f
C875 B.n658 VSUBS 0.00697f
C876 B.n659 VSUBS 0.00697f
C877 B.n660 VSUBS 0.00697f
C878 B.n661 VSUBS 0.00697f
C879 B.n662 VSUBS 0.00697f
C880 B.n663 VSUBS 0.015782f
.ends

