* NGSPICE file created from diff_pair_sample_1382.ext - technology: sky130A

.subckt diff_pair_sample_1382 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=4.2042 pd=22.34 as=1.7787 ps=11.11 w=10.78 l=2.22
X1 VTAIL.t2 VN.t0 VDD2.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=1.7787 pd=11.11 as=1.7787 ps=11.11 w=10.78 l=2.22
X2 VTAIL.t14 VP.t1 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=4.2042 pd=22.34 as=1.7787 ps=11.11 w=10.78 l=2.22
X3 VTAIL.t1 VN.t1 VDD2.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=4.2042 pd=22.34 as=1.7787 ps=11.11 w=10.78 l=2.22
X4 VDD1.t2 VP.t2 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=1.7787 pd=11.11 as=1.7787 ps=11.11 w=10.78 l=2.22
X5 VDD2.t5 VN.t2 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.7787 pd=11.11 as=1.7787 ps=11.11 w=10.78 l=2.22
X6 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=4.2042 pd=22.34 as=0 ps=0 w=10.78 l=2.22
X7 VDD2.t4 VN.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.7787 pd=11.11 as=4.2042 ps=22.34 w=10.78 l=2.22
X8 VDD1.t3 VP.t3 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=1.7787 pd=11.11 as=4.2042 ps=22.34 w=10.78 l=2.22
X9 VDD2.t3 VN.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.7787 pd=11.11 as=1.7787 ps=11.11 w=10.78 l=2.22
X10 VTAIL.t0 VN.t5 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=4.2042 pd=22.34 as=1.7787 ps=11.11 w=10.78 l=2.22
X11 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=4.2042 pd=22.34 as=0 ps=0 w=10.78 l=2.22
X12 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.2042 pd=22.34 as=0 ps=0 w=10.78 l=2.22
X13 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.2042 pd=22.34 as=0 ps=0 w=10.78 l=2.22
X14 VDD2.t1 VN.t6 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.7787 pd=11.11 as=4.2042 ps=22.34 w=10.78 l=2.22
X15 VTAIL.t11 VP.t4 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.7787 pd=11.11 as=1.7787 ps=11.11 w=10.78 l=2.22
X16 VDD1.t5 VP.t5 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=1.7787 pd=11.11 as=4.2042 ps=22.34 w=10.78 l=2.22
X17 VTAIL.t9 VP.t6 VDD1.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.7787 pd=11.11 as=1.7787 ps=11.11 w=10.78 l=2.22
X18 VDD1.t7 VP.t7 VTAIL.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.7787 pd=11.11 as=1.7787 ps=11.11 w=10.78 l=2.22
X19 VTAIL.t3 VN.t7 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.7787 pd=11.11 as=1.7787 ps=11.11 w=10.78 l=2.22
R0 VP.n16 VP.n15 161.3
R1 VP.n17 VP.n12 161.3
R2 VP.n19 VP.n18 161.3
R3 VP.n20 VP.n11 161.3
R4 VP.n22 VP.n21 161.3
R5 VP.n24 VP.n10 161.3
R6 VP.n26 VP.n25 161.3
R7 VP.n27 VP.n9 161.3
R8 VP.n29 VP.n28 161.3
R9 VP.n30 VP.n8 161.3
R10 VP.n58 VP.n0 161.3
R11 VP.n57 VP.n56 161.3
R12 VP.n55 VP.n1 161.3
R13 VP.n54 VP.n53 161.3
R14 VP.n52 VP.n2 161.3
R15 VP.n50 VP.n49 161.3
R16 VP.n48 VP.n3 161.3
R17 VP.n47 VP.n46 161.3
R18 VP.n45 VP.n4 161.3
R19 VP.n44 VP.n43 161.3
R20 VP.n42 VP.n41 161.3
R21 VP.n40 VP.n6 161.3
R22 VP.n39 VP.n38 161.3
R23 VP.n37 VP.n7 161.3
R24 VP.n36 VP.n35 161.3
R25 VP.n14 VP.t0 150.167
R26 VP.n34 VP.t1 117.026
R27 VP.n5 VP.t7 117.026
R28 VP.n51 VP.t4 117.026
R29 VP.n59 VP.t3 117.026
R30 VP.n31 VP.t5 117.026
R31 VP.n23 VP.t6 117.026
R32 VP.n13 VP.t2 117.026
R33 VP.n34 VP.n33 94.9235
R34 VP.n60 VP.n59 94.9235
R35 VP.n32 VP.n31 94.9235
R36 VP.n14 VP.n13 58.066
R37 VP.n33 VP.n32 48.2118
R38 VP.n39 VP.n7 45.4209
R39 VP.n57 VP.n1 45.4209
R40 VP.n29 VP.n9 45.4209
R41 VP.n46 VP.n45 40.577
R42 VP.n46 VP.n3 40.577
R43 VP.n18 VP.n11 40.577
R44 VP.n18 VP.n17 40.577
R45 VP.n40 VP.n39 35.7332
R46 VP.n53 VP.n1 35.7332
R47 VP.n25 VP.n9 35.7332
R48 VP.n35 VP.n7 24.5923
R49 VP.n41 VP.n40 24.5923
R50 VP.n45 VP.n44 24.5923
R51 VP.n50 VP.n3 24.5923
R52 VP.n53 VP.n52 24.5923
R53 VP.n58 VP.n57 24.5923
R54 VP.n30 VP.n29 24.5923
R55 VP.n22 VP.n11 24.5923
R56 VP.n25 VP.n24 24.5923
R57 VP.n17 VP.n16 24.5923
R58 VP.n35 VP.n34 15.9852
R59 VP.n59 VP.n58 15.9852
R60 VP.n31 VP.n30 15.9852
R61 VP.n44 VP.n5 13.526
R62 VP.n51 VP.n50 13.526
R63 VP.n23 VP.n22 13.526
R64 VP.n16 VP.n13 13.526
R65 VP.n41 VP.n5 11.0668
R66 VP.n52 VP.n51 11.0668
R67 VP.n24 VP.n23 11.0668
R68 VP.n15 VP.n14 9.34229
R69 VP.n32 VP.n8 0.278335
R70 VP.n36 VP.n33 0.278335
R71 VP.n60 VP.n0 0.278335
R72 VP.n15 VP.n12 0.189894
R73 VP.n19 VP.n12 0.189894
R74 VP.n20 VP.n19 0.189894
R75 VP.n21 VP.n20 0.189894
R76 VP.n21 VP.n10 0.189894
R77 VP.n26 VP.n10 0.189894
R78 VP.n27 VP.n26 0.189894
R79 VP.n28 VP.n27 0.189894
R80 VP.n28 VP.n8 0.189894
R81 VP.n37 VP.n36 0.189894
R82 VP.n38 VP.n37 0.189894
R83 VP.n38 VP.n6 0.189894
R84 VP.n42 VP.n6 0.189894
R85 VP.n43 VP.n42 0.189894
R86 VP.n43 VP.n4 0.189894
R87 VP.n47 VP.n4 0.189894
R88 VP.n48 VP.n47 0.189894
R89 VP.n49 VP.n48 0.189894
R90 VP.n49 VP.n2 0.189894
R91 VP.n54 VP.n2 0.189894
R92 VP.n55 VP.n54 0.189894
R93 VP.n56 VP.n55 0.189894
R94 VP.n56 VP.n0 0.189894
R95 VP VP.n60 0.153485
R96 VDD1 VDD1.n0 65.437
R97 VDD1.n3 VDD1.n2 65.3233
R98 VDD1.n3 VDD1.n1 65.3233
R99 VDD1.n5 VDD1.n4 64.2795
R100 VDD1.n5 VDD1.n3 43.4837
R101 VDD1.n4 VDD1.t6 1.83723
R102 VDD1.n4 VDD1.t5 1.83723
R103 VDD1.n0 VDD1.t0 1.83723
R104 VDD1.n0 VDD1.t2 1.83723
R105 VDD1.n2 VDD1.t4 1.83723
R106 VDD1.n2 VDD1.t3 1.83723
R107 VDD1.n1 VDD1.t1 1.83723
R108 VDD1.n1 VDD1.t7 1.83723
R109 VDD1 VDD1.n5 1.04145
R110 VTAIL.n466 VTAIL.n414 289.615
R111 VTAIL.n54 VTAIL.n2 289.615
R112 VTAIL.n112 VTAIL.n60 289.615
R113 VTAIL.n172 VTAIL.n120 289.615
R114 VTAIL.n408 VTAIL.n356 289.615
R115 VTAIL.n348 VTAIL.n296 289.615
R116 VTAIL.n290 VTAIL.n238 289.615
R117 VTAIL.n230 VTAIL.n178 289.615
R118 VTAIL.n433 VTAIL.n432 185
R119 VTAIL.n430 VTAIL.n429 185
R120 VTAIL.n439 VTAIL.n438 185
R121 VTAIL.n441 VTAIL.n440 185
R122 VTAIL.n426 VTAIL.n425 185
R123 VTAIL.n447 VTAIL.n446 185
R124 VTAIL.n450 VTAIL.n449 185
R125 VTAIL.n448 VTAIL.n422 185
R126 VTAIL.n455 VTAIL.n421 185
R127 VTAIL.n457 VTAIL.n456 185
R128 VTAIL.n459 VTAIL.n458 185
R129 VTAIL.n418 VTAIL.n417 185
R130 VTAIL.n465 VTAIL.n464 185
R131 VTAIL.n467 VTAIL.n466 185
R132 VTAIL.n21 VTAIL.n20 185
R133 VTAIL.n18 VTAIL.n17 185
R134 VTAIL.n27 VTAIL.n26 185
R135 VTAIL.n29 VTAIL.n28 185
R136 VTAIL.n14 VTAIL.n13 185
R137 VTAIL.n35 VTAIL.n34 185
R138 VTAIL.n38 VTAIL.n37 185
R139 VTAIL.n36 VTAIL.n10 185
R140 VTAIL.n43 VTAIL.n9 185
R141 VTAIL.n45 VTAIL.n44 185
R142 VTAIL.n47 VTAIL.n46 185
R143 VTAIL.n6 VTAIL.n5 185
R144 VTAIL.n53 VTAIL.n52 185
R145 VTAIL.n55 VTAIL.n54 185
R146 VTAIL.n79 VTAIL.n78 185
R147 VTAIL.n76 VTAIL.n75 185
R148 VTAIL.n85 VTAIL.n84 185
R149 VTAIL.n87 VTAIL.n86 185
R150 VTAIL.n72 VTAIL.n71 185
R151 VTAIL.n93 VTAIL.n92 185
R152 VTAIL.n96 VTAIL.n95 185
R153 VTAIL.n94 VTAIL.n68 185
R154 VTAIL.n101 VTAIL.n67 185
R155 VTAIL.n103 VTAIL.n102 185
R156 VTAIL.n105 VTAIL.n104 185
R157 VTAIL.n64 VTAIL.n63 185
R158 VTAIL.n111 VTAIL.n110 185
R159 VTAIL.n113 VTAIL.n112 185
R160 VTAIL.n139 VTAIL.n138 185
R161 VTAIL.n136 VTAIL.n135 185
R162 VTAIL.n145 VTAIL.n144 185
R163 VTAIL.n147 VTAIL.n146 185
R164 VTAIL.n132 VTAIL.n131 185
R165 VTAIL.n153 VTAIL.n152 185
R166 VTAIL.n156 VTAIL.n155 185
R167 VTAIL.n154 VTAIL.n128 185
R168 VTAIL.n161 VTAIL.n127 185
R169 VTAIL.n163 VTAIL.n162 185
R170 VTAIL.n165 VTAIL.n164 185
R171 VTAIL.n124 VTAIL.n123 185
R172 VTAIL.n171 VTAIL.n170 185
R173 VTAIL.n173 VTAIL.n172 185
R174 VTAIL.n409 VTAIL.n408 185
R175 VTAIL.n407 VTAIL.n406 185
R176 VTAIL.n360 VTAIL.n359 185
R177 VTAIL.n401 VTAIL.n400 185
R178 VTAIL.n399 VTAIL.n398 185
R179 VTAIL.n397 VTAIL.n363 185
R180 VTAIL.n367 VTAIL.n364 185
R181 VTAIL.n392 VTAIL.n391 185
R182 VTAIL.n390 VTAIL.n389 185
R183 VTAIL.n369 VTAIL.n368 185
R184 VTAIL.n384 VTAIL.n383 185
R185 VTAIL.n382 VTAIL.n381 185
R186 VTAIL.n373 VTAIL.n372 185
R187 VTAIL.n376 VTAIL.n375 185
R188 VTAIL.n349 VTAIL.n348 185
R189 VTAIL.n347 VTAIL.n346 185
R190 VTAIL.n300 VTAIL.n299 185
R191 VTAIL.n341 VTAIL.n340 185
R192 VTAIL.n339 VTAIL.n338 185
R193 VTAIL.n337 VTAIL.n303 185
R194 VTAIL.n307 VTAIL.n304 185
R195 VTAIL.n332 VTAIL.n331 185
R196 VTAIL.n330 VTAIL.n329 185
R197 VTAIL.n309 VTAIL.n308 185
R198 VTAIL.n324 VTAIL.n323 185
R199 VTAIL.n322 VTAIL.n321 185
R200 VTAIL.n313 VTAIL.n312 185
R201 VTAIL.n316 VTAIL.n315 185
R202 VTAIL.n291 VTAIL.n290 185
R203 VTAIL.n289 VTAIL.n288 185
R204 VTAIL.n242 VTAIL.n241 185
R205 VTAIL.n283 VTAIL.n282 185
R206 VTAIL.n281 VTAIL.n280 185
R207 VTAIL.n279 VTAIL.n245 185
R208 VTAIL.n249 VTAIL.n246 185
R209 VTAIL.n274 VTAIL.n273 185
R210 VTAIL.n272 VTAIL.n271 185
R211 VTAIL.n251 VTAIL.n250 185
R212 VTAIL.n266 VTAIL.n265 185
R213 VTAIL.n264 VTAIL.n263 185
R214 VTAIL.n255 VTAIL.n254 185
R215 VTAIL.n258 VTAIL.n257 185
R216 VTAIL.n231 VTAIL.n230 185
R217 VTAIL.n229 VTAIL.n228 185
R218 VTAIL.n182 VTAIL.n181 185
R219 VTAIL.n223 VTAIL.n222 185
R220 VTAIL.n221 VTAIL.n220 185
R221 VTAIL.n219 VTAIL.n185 185
R222 VTAIL.n189 VTAIL.n186 185
R223 VTAIL.n214 VTAIL.n213 185
R224 VTAIL.n212 VTAIL.n211 185
R225 VTAIL.n191 VTAIL.n190 185
R226 VTAIL.n206 VTAIL.n205 185
R227 VTAIL.n204 VTAIL.n203 185
R228 VTAIL.n195 VTAIL.n194 185
R229 VTAIL.n198 VTAIL.n197 185
R230 VTAIL.t6 VTAIL.n431 149.524
R231 VTAIL.t1 VTAIL.n19 149.524
R232 VTAIL.t12 VTAIL.n77 149.524
R233 VTAIL.t14 VTAIL.n137 149.524
R234 VTAIL.t10 VTAIL.n374 149.524
R235 VTAIL.t15 VTAIL.n314 149.524
R236 VTAIL.t4 VTAIL.n256 149.524
R237 VTAIL.t0 VTAIL.n196 149.524
R238 VTAIL.n432 VTAIL.n429 104.615
R239 VTAIL.n439 VTAIL.n429 104.615
R240 VTAIL.n440 VTAIL.n439 104.615
R241 VTAIL.n440 VTAIL.n425 104.615
R242 VTAIL.n447 VTAIL.n425 104.615
R243 VTAIL.n449 VTAIL.n447 104.615
R244 VTAIL.n449 VTAIL.n448 104.615
R245 VTAIL.n448 VTAIL.n421 104.615
R246 VTAIL.n457 VTAIL.n421 104.615
R247 VTAIL.n458 VTAIL.n457 104.615
R248 VTAIL.n458 VTAIL.n417 104.615
R249 VTAIL.n465 VTAIL.n417 104.615
R250 VTAIL.n466 VTAIL.n465 104.615
R251 VTAIL.n20 VTAIL.n17 104.615
R252 VTAIL.n27 VTAIL.n17 104.615
R253 VTAIL.n28 VTAIL.n27 104.615
R254 VTAIL.n28 VTAIL.n13 104.615
R255 VTAIL.n35 VTAIL.n13 104.615
R256 VTAIL.n37 VTAIL.n35 104.615
R257 VTAIL.n37 VTAIL.n36 104.615
R258 VTAIL.n36 VTAIL.n9 104.615
R259 VTAIL.n45 VTAIL.n9 104.615
R260 VTAIL.n46 VTAIL.n45 104.615
R261 VTAIL.n46 VTAIL.n5 104.615
R262 VTAIL.n53 VTAIL.n5 104.615
R263 VTAIL.n54 VTAIL.n53 104.615
R264 VTAIL.n78 VTAIL.n75 104.615
R265 VTAIL.n85 VTAIL.n75 104.615
R266 VTAIL.n86 VTAIL.n85 104.615
R267 VTAIL.n86 VTAIL.n71 104.615
R268 VTAIL.n93 VTAIL.n71 104.615
R269 VTAIL.n95 VTAIL.n93 104.615
R270 VTAIL.n95 VTAIL.n94 104.615
R271 VTAIL.n94 VTAIL.n67 104.615
R272 VTAIL.n103 VTAIL.n67 104.615
R273 VTAIL.n104 VTAIL.n103 104.615
R274 VTAIL.n104 VTAIL.n63 104.615
R275 VTAIL.n111 VTAIL.n63 104.615
R276 VTAIL.n112 VTAIL.n111 104.615
R277 VTAIL.n138 VTAIL.n135 104.615
R278 VTAIL.n145 VTAIL.n135 104.615
R279 VTAIL.n146 VTAIL.n145 104.615
R280 VTAIL.n146 VTAIL.n131 104.615
R281 VTAIL.n153 VTAIL.n131 104.615
R282 VTAIL.n155 VTAIL.n153 104.615
R283 VTAIL.n155 VTAIL.n154 104.615
R284 VTAIL.n154 VTAIL.n127 104.615
R285 VTAIL.n163 VTAIL.n127 104.615
R286 VTAIL.n164 VTAIL.n163 104.615
R287 VTAIL.n164 VTAIL.n123 104.615
R288 VTAIL.n171 VTAIL.n123 104.615
R289 VTAIL.n172 VTAIL.n171 104.615
R290 VTAIL.n408 VTAIL.n407 104.615
R291 VTAIL.n407 VTAIL.n359 104.615
R292 VTAIL.n400 VTAIL.n359 104.615
R293 VTAIL.n400 VTAIL.n399 104.615
R294 VTAIL.n399 VTAIL.n363 104.615
R295 VTAIL.n367 VTAIL.n363 104.615
R296 VTAIL.n391 VTAIL.n367 104.615
R297 VTAIL.n391 VTAIL.n390 104.615
R298 VTAIL.n390 VTAIL.n368 104.615
R299 VTAIL.n383 VTAIL.n368 104.615
R300 VTAIL.n383 VTAIL.n382 104.615
R301 VTAIL.n382 VTAIL.n372 104.615
R302 VTAIL.n375 VTAIL.n372 104.615
R303 VTAIL.n348 VTAIL.n347 104.615
R304 VTAIL.n347 VTAIL.n299 104.615
R305 VTAIL.n340 VTAIL.n299 104.615
R306 VTAIL.n340 VTAIL.n339 104.615
R307 VTAIL.n339 VTAIL.n303 104.615
R308 VTAIL.n307 VTAIL.n303 104.615
R309 VTAIL.n331 VTAIL.n307 104.615
R310 VTAIL.n331 VTAIL.n330 104.615
R311 VTAIL.n330 VTAIL.n308 104.615
R312 VTAIL.n323 VTAIL.n308 104.615
R313 VTAIL.n323 VTAIL.n322 104.615
R314 VTAIL.n322 VTAIL.n312 104.615
R315 VTAIL.n315 VTAIL.n312 104.615
R316 VTAIL.n290 VTAIL.n289 104.615
R317 VTAIL.n289 VTAIL.n241 104.615
R318 VTAIL.n282 VTAIL.n241 104.615
R319 VTAIL.n282 VTAIL.n281 104.615
R320 VTAIL.n281 VTAIL.n245 104.615
R321 VTAIL.n249 VTAIL.n245 104.615
R322 VTAIL.n273 VTAIL.n249 104.615
R323 VTAIL.n273 VTAIL.n272 104.615
R324 VTAIL.n272 VTAIL.n250 104.615
R325 VTAIL.n265 VTAIL.n250 104.615
R326 VTAIL.n265 VTAIL.n264 104.615
R327 VTAIL.n264 VTAIL.n254 104.615
R328 VTAIL.n257 VTAIL.n254 104.615
R329 VTAIL.n230 VTAIL.n229 104.615
R330 VTAIL.n229 VTAIL.n181 104.615
R331 VTAIL.n222 VTAIL.n181 104.615
R332 VTAIL.n222 VTAIL.n221 104.615
R333 VTAIL.n221 VTAIL.n185 104.615
R334 VTAIL.n189 VTAIL.n185 104.615
R335 VTAIL.n213 VTAIL.n189 104.615
R336 VTAIL.n213 VTAIL.n212 104.615
R337 VTAIL.n212 VTAIL.n190 104.615
R338 VTAIL.n205 VTAIL.n190 104.615
R339 VTAIL.n205 VTAIL.n204 104.615
R340 VTAIL.n204 VTAIL.n194 104.615
R341 VTAIL.n197 VTAIL.n194 104.615
R342 VTAIL.n432 VTAIL.t6 52.3082
R343 VTAIL.n20 VTAIL.t1 52.3082
R344 VTAIL.n78 VTAIL.t12 52.3082
R345 VTAIL.n138 VTAIL.t14 52.3082
R346 VTAIL.n375 VTAIL.t10 52.3082
R347 VTAIL.n315 VTAIL.t15 52.3082
R348 VTAIL.n257 VTAIL.t4 52.3082
R349 VTAIL.n197 VTAIL.t0 52.3082
R350 VTAIL.n355 VTAIL.n354 47.6009
R351 VTAIL.n237 VTAIL.n236 47.6009
R352 VTAIL.n1 VTAIL.n0 47.6007
R353 VTAIL.n119 VTAIL.n118 47.6007
R354 VTAIL.n471 VTAIL.n470 34.1247
R355 VTAIL.n59 VTAIL.n58 34.1247
R356 VTAIL.n117 VTAIL.n116 34.1247
R357 VTAIL.n177 VTAIL.n176 34.1247
R358 VTAIL.n413 VTAIL.n412 34.1247
R359 VTAIL.n353 VTAIL.n352 34.1247
R360 VTAIL.n295 VTAIL.n294 34.1247
R361 VTAIL.n235 VTAIL.n234 34.1247
R362 VTAIL.n471 VTAIL.n413 23.8583
R363 VTAIL.n235 VTAIL.n177 23.8583
R364 VTAIL.n456 VTAIL.n455 13.1884
R365 VTAIL.n44 VTAIL.n43 13.1884
R366 VTAIL.n102 VTAIL.n101 13.1884
R367 VTAIL.n162 VTAIL.n161 13.1884
R368 VTAIL.n398 VTAIL.n397 13.1884
R369 VTAIL.n338 VTAIL.n337 13.1884
R370 VTAIL.n280 VTAIL.n279 13.1884
R371 VTAIL.n220 VTAIL.n219 13.1884
R372 VTAIL.n454 VTAIL.n422 12.8005
R373 VTAIL.n459 VTAIL.n420 12.8005
R374 VTAIL.n42 VTAIL.n10 12.8005
R375 VTAIL.n47 VTAIL.n8 12.8005
R376 VTAIL.n100 VTAIL.n68 12.8005
R377 VTAIL.n105 VTAIL.n66 12.8005
R378 VTAIL.n160 VTAIL.n128 12.8005
R379 VTAIL.n165 VTAIL.n126 12.8005
R380 VTAIL.n401 VTAIL.n362 12.8005
R381 VTAIL.n396 VTAIL.n364 12.8005
R382 VTAIL.n341 VTAIL.n302 12.8005
R383 VTAIL.n336 VTAIL.n304 12.8005
R384 VTAIL.n283 VTAIL.n244 12.8005
R385 VTAIL.n278 VTAIL.n246 12.8005
R386 VTAIL.n223 VTAIL.n184 12.8005
R387 VTAIL.n218 VTAIL.n186 12.8005
R388 VTAIL.n451 VTAIL.n450 12.0247
R389 VTAIL.n460 VTAIL.n418 12.0247
R390 VTAIL.n39 VTAIL.n38 12.0247
R391 VTAIL.n48 VTAIL.n6 12.0247
R392 VTAIL.n97 VTAIL.n96 12.0247
R393 VTAIL.n106 VTAIL.n64 12.0247
R394 VTAIL.n157 VTAIL.n156 12.0247
R395 VTAIL.n166 VTAIL.n124 12.0247
R396 VTAIL.n402 VTAIL.n360 12.0247
R397 VTAIL.n393 VTAIL.n392 12.0247
R398 VTAIL.n342 VTAIL.n300 12.0247
R399 VTAIL.n333 VTAIL.n332 12.0247
R400 VTAIL.n284 VTAIL.n242 12.0247
R401 VTAIL.n275 VTAIL.n274 12.0247
R402 VTAIL.n224 VTAIL.n182 12.0247
R403 VTAIL.n215 VTAIL.n214 12.0247
R404 VTAIL.n446 VTAIL.n424 11.249
R405 VTAIL.n464 VTAIL.n463 11.249
R406 VTAIL.n34 VTAIL.n12 11.249
R407 VTAIL.n52 VTAIL.n51 11.249
R408 VTAIL.n92 VTAIL.n70 11.249
R409 VTAIL.n110 VTAIL.n109 11.249
R410 VTAIL.n152 VTAIL.n130 11.249
R411 VTAIL.n170 VTAIL.n169 11.249
R412 VTAIL.n406 VTAIL.n405 11.249
R413 VTAIL.n389 VTAIL.n366 11.249
R414 VTAIL.n346 VTAIL.n345 11.249
R415 VTAIL.n329 VTAIL.n306 11.249
R416 VTAIL.n288 VTAIL.n287 11.249
R417 VTAIL.n271 VTAIL.n248 11.249
R418 VTAIL.n228 VTAIL.n227 11.249
R419 VTAIL.n211 VTAIL.n188 11.249
R420 VTAIL.n445 VTAIL.n426 10.4732
R421 VTAIL.n467 VTAIL.n416 10.4732
R422 VTAIL.n33 VTAIL.n14 10.4732
R423 VTAIL.n55 VTAIL.n4 10.4732
R424 VTAIL.n91 VTAIL.n72 10.4732
R425 VTAIL.n113 VTAIL.n62 10.4732
R426 VTAIL.n151 VTAIL.n132 10.4732
R427 VTAIL.n173 VTAIL.n122 10.4732
R428 VTAIL.n409 VTAIL.n358 10.4732
R429 VTAIL.n388 VTAIL.n369 10.4732
R430 VTAIL.n349 VTAIL.n298 10.4732
R431 VTAIL.n328 VTAIL.n309 10.4732
R432 VTAIL.n291 VTAIL.n240 10.4732
R433 VTAIL.n270 VTAIL.n251 10.4732
R434 VTAIL.n231 VTAIL.n180 10.4732
R435 VTAIL.n210 VTAIL.n191 10.4732
R436 VTAIL.n433 VTAIL.n431 10.2747
R437 VTAIL.n21 VTAIL.n19 10.2747
R438 VTAIL.n79 VTAIL.n77 10.2747
R439 VTAIL.n139 VTAIL.n137 10.2747
R440 VTAIL.n376 VTAIL.n374 10.2747
R441 VTAIL.n316 VTAIL.n314 10.2747
R442 VTAIL.n258 VTAIL.n256 10.2747
R443 VTAIL.n198 VTAIL.n196 10.2747
R444 VTAIL.n442 VTAIL.n441 9.69747
R445 VTAIL.n468 VTAIL.n414 9.69747
R446 VTAIL.n30 VTAIL.n29 9.69747
R447 VTAIL.n56 VTAIL.n2 9.69747
R448 VTAIL.n88 VTAIL.n87 9.69747
R449 VTAIL.n114 VTAIL.n60 9.69747
R450 VTAIL.n148 VTAIL.n147 9.69747
R451 VTAIL.n174 VTAIL.n120 9.69747
R452 VTAIL.n410 VTAIL.n356 9.69747
R453 VTAIL.n385 VTAIL.n384 9.69747
R454 VTAIL.n350 VTAIL.n296 9.69747
R455 VTAIL.n325 VTAIL.n324 9.69747
R456 VTAIL.n292 VTAIL.n238 9.69747
R457 VTAIL.n267 VTAIL.n266 9.69747
R458 VTAIL.n232 VTAIL.n178 9.69747
R459 VTAIL.n207 VTAIL.n206 9.69747
R460 VTAIL.n470 VTAIL.n469 9.45567
R461 VTAIL.n58 VTAIL.n57 9.45567
R462 VTAIL.n116 VTAIL.n115 9.45567
R463 VTAIL.n176 VTAIL.n175 9.45567
R464 VTAIL.n412 VTAIL.n411 9.45567
R465 VTAIL.n352 VTAIL.n351 9.45567
R466 VTAIL.n294 VTAIL.n293 9.45567
R467 VTAIL.n234 VTAIL.n233 9.45567
R468 VTAIL.n469 VTAIL.n468 9.3005
R469 VTAIL.n416 VTAIL.n415 9.3005
R470 VTAIL.n463 VTAIL.n462 9.3005
R471 VTAIL.n461 VTAIL.n460 9.3005
R472 VTAIL.n420 VTAIL.n419 9.3005
R473 VTAIL.n435 VTAIL.n434 9.3005
R474 VTAIL.n437 VTAIL.n436 9.3005
R475 VTAIL.n428 VTAIL.n427 9.3005
R476 VTAIL.n443 VTAIL.n442 9.3005
R477 VTAIL.n445 VTAIL.n444 9.3005
R478 VTAIL.n424 VTAIL.n423 9.3005
R479 VTAIL.n452 VTAIL.n451 9.3005
R480 VTAIL.n454 VTAIL.n453 9.3005
R481 VTAIL.n57 VTAIL.n56 9.3005
R482 VTAIL.n4 VTAIL.n3 9.3005
R483 VTAIL.n51 VTAIL.n50 9.3005
R484 VTAIL.n49 VTAIL.n48 9.3005
R485 VTAIL.n8 VTAIL.n7 9.3005
R486 VTAIL.n23 VTAIL.n22 9.3005
R487 VTAIL.n25 VTAIL.n24 9.3005
R488 VTAIL.n16 VTAIL.n15 9.3005
R489 VTAIL.n31 VTAIL.n30 9.3005
R490 VTAIL.n33 VTAIL.n32 9.3005
R491 VTAIL.n12 VTAIL.n11 9.3005
R492 VTAIL.n40 VTAIL.n39 9.3005
R493 VTAIL.n42 VTAIL.n41 9.3005
R494 VTAIL.n115 VTAIL.n114 9.3005
R495 VTAIL.n62 VTAIL.n61 9.3005
R496 VTAIL.n109 VTAIL.n108 9.3005
R497 VTAIL.n107 VTAIL.n106 9.3005
R498 VTAIL.n66 VTAIL.n65 9.3005
R499 VTAIL.n81 VTAIL.n80 9.3005
R500 VTAIL.n83 VTAIL.n82 9.3005
R501 VTAIL.n74 VTAIL.n73 9.3005
R502 VTAIL.n89 VTAIL.n88 9.3005
R503 VTAIL.n91 VTAIL.n90 9.3005
R504 VTAIL.n70 VTAIL.n69 9.3005
R505 VTAIL.n98 VTAIL.n97 9.3005
R506 VTAIL.n100 VTAIL.n99 9.3005
R507 VTAIL.n175 VTAIL.n174 9.3005
R508 VTAIL.n122 VTAIL.n121 9.3005
R509 VTAIL.n169 VTAIL.n168 9.3005
R510 VTAIL.n167 VTAIL.n166 9.3005
R511 VTAIL.n126 VTAIL.n125 9.3005
R512 VTAIL.n141 VTAIL.n140 9.3005
R513 VTAIL.n143 VTAIL.n142 9.3005
R514 VTAIL.n134 VTAIL.n133 9.3005
R515 VTAIL.n149 VTAIL.n148 9.3005
R516 VTAIL.n151 VTAIL.n150 9.3005
R517 VTAIL.n130 VTAIL.n129 9.3005
R518 VTAIL.n158 VTAIL.n157 9.3005
R519 VTAIL.n160 VTAIL.n159 9.3005
R520 VTAIL.n378 VTAIL.n377 9.3005
R521 VTAIL.n380 VTAIL.n379 9.3005
R522 VTAIL.n371 VTAIL.n370 9.3005
R523 VTAIL.n386 VTAIL.n385 9.3005
R524 VTAIL.n388 VTAIL.n387 9.3005
R525 VTAIL.n366 VTAIL.n365 9.3005
R526 VTAIL.n394 VTAIL.n393 9.3005
R527 VTAIL.n396 VTAIL.n395 9.3005
R528 VTAIL.n411 VTAIL.n410 9.3005
R529 VTAIL.n358 VTAIL.n357 9.3005
R530 VTAIL.n405 VTAIL.n404 9.3005
R531 VTAIL.n403 VTAIL.n402 9.3005
R532 VTAIL.n362 VTAIL.n361 9.3005
R533 VTAIL.n318 VTAIL.n317 9.3005
R534 VTAIL.n320 VTAIL.n319 9.3005
R535 VTAIL.n311 VTAIL.n310 9.3005
R536 VTAIL.n326 VTAIL.n325 9.3005
R537 VTAIL.n328 VTAIL.n327 9.3005
R538 VTAIL.n306 VTAIL.n305 9.3005
R539 VTAIL.n334 VTAIL.n333 9.3005
R540 VTAIL.n336 VTAIL.n335 9.3005
R541 VTAIL.n351 VTAIL.n350 9.3005
R542 VTAIL.n298 VTAIL.n297 9.3005
R543 VTAIL.n345 VTAIL.n344 9.3005
R544 VTAIL.n343 VTAIL.n342 9.3005
R545 VTAIL.n302 VTAIL.n301 9.3005
R546 VTAIL.n260 VTAIL.n259 9.3005
R547 VTAIL.n262 VTAIL.n261 9.3005
R548 VTAIL.n253 VTAIL.n252 9.3005
R549 VTAIL.n268 VTAIL.n267 9.3005
R550 VTAIL.n270 VTAIL.n269 9.3005
R551 VTAIL.n248 VTAIL.n247 9.3005
R552 VTAIL.n276 VTAIL.n275 9.3005
R553 VTAIL.n278 VTAIL.n277 9.3005
R554 VTAIL.n293 VTAIL.n292 9.3005
R555 VTAIL.n240 VTAIL.n239 9.3005
R556 VTAIL.n287 VTAIL.n286 9.3005
R557 VTAIL.n285 VTAIL.n284 9.3005
R558 VTAIL.n244 VTAIL.n243 9.3005
R559 VTAIL.n200 VTAIL.n199 9.3005
R560 VTAIL.n202 VTAIL.n201 9.3005
R561 VTAIL.n193 VTAIL.n192 9.3005
R562 VTAIL.n208 VTAIL.n207 9.3005
R563 VTAIL.n210 VTAIL.n209 9.3005
R564 VTAIL.n188 VTAIL.n187 9.3005
R565 VTAIL.n216 VTAIL.n215 9.3005
R566 VTAIL.n218 VTAIL.n217 9.3005
R567 VTAIL.n233 VTAIL.n232 9.3005
R568 VTAIL.n180 VTAIL.n179 9.3005
R569 VTAIL.n227 VTAIL.n226 9.3005
R570 VTAIL.n225 VTAIL.n224 9.3005
R571 VTAIL.n184 VTAIL.n183 9.3005
R572 VTAIL.n438 VTAIL.n428 8.92171
R573 VTAIL.n26 VTAIL.n16 8.92171
R574 VTAIL.n84 VTAIL.n74 8.92171
R575 VTAIL.n144 VTAIL.n134 8.92171
R576 VTAIL.n381 VTAIL.n371 8.92171
R577 VTAIL.n321 VTAIL.n311 8.92171
R578 VTAIL.n263 VTAIL.n253 8.92171
R579 VTAIL.n203 VTAIL.n193 8.92171
R580 VTAIL.n437 VTAIL.n430 8.14595
R581 VTAIL.n25 VTAIL.n18 8.14595
R582 VTAIL.n83 VTAIL.n76 8.14595
R583 VTAIL.n143 VTAIL.n136 8.14595
R584 VTAIL.n380 VTAIL.n373 8.14595
R585 VTAIL.n320 VTAIL.n313 8.14595
R586 VTAIL.n262 VTAIL.n255 8.14595
R587 VTAIL.n202 VTAIL.n195 8.14595
R588 VTAIL.n434 VTAIL.n433 7.3702
R589 VTAIL.n22 VTAIL.n21 7.3702
R590 VTAIL.n80 VTAIL.n79 7.3702
R591 VTAIL.n140 VTAIL.n139 7.3702
R592 VTAIL.n377 VTAIL.n376 7.3702
R593 VTAIL.n317 VTAIL.n316 7.3702
R594 VTAIL.n259 VTAIL.n258 7.3702
R595 VTAIL.n199 VTAIL.n198 7.3702
R596 VTAIL.n434 VTAIL.n430 5.81868
R597 VTAIL.n22 VTAIL.n18 5.81868
R598 VTAIL.n80 VTAIL.n76 5.81868
R599 VTAIL.n140 VTAIL.n136 5.81868
R600 VTAIL.n377 VTAIL.n373 5.81868
R601 VTAIL.n317 VTAIL.n313 5.81868
R602 VTAIL.n259 VTAIL.n255 5.81868
R603 VTAIL.n199 VTAIL.n195 5.81868
R604 VTAIL.n438 VTAIL.n437 5.04292
R605 VTAIL.n26 VTAIL.n25 5.04292
R606 VTAIL.n84 VTAIL.n83 5.04292
R607 VTAIL.n144 VTAIL.n143 5.04292
R608 VTAIL.n381 VTAIL.n380 5.04292
R609 VTAIL.n321 VTAIL.n320 5.04292
R610 VTAIL.n263 VTAIL.n262 5.04292
R611 VTAIL.n203 VTAIL.n202 5.04292
R612 VTAIL.n441 VTAIL.n428 4.26717
R613 VTAIL.n470 VTAIL.n414 4.26717
R614 VTAIL.n29 VTAIL.n16 4.26717
R615 VTAIL.n58 VTAIL.n2 4.26717
R616 VTAIL.n87 VTAIL.n74 4.26717
R617 VTAIL.n116 VTAIL.n60 4.26717
R618 VTAIL.n147 VTAIL.n134 4.26717
R619 VTAIL.n176 VTAIL.n120 4.26717
R620 VTAIL.n412 VTAIL.n356 4.26717
R621 VTAIL.n384 VTAIL.n371 4.26717
R622 VTAIL.n352 VTAIL.n296 4.26717
R623 VTAIL.n324 VTAIL.n311 4.26717
R624 VTAIL.n294 VTAIL.n238 4.26717
R625 VTAIL.n266 VTAIL.n253 4.26717
R626 VTAIL.n234 VTAIL.n178 4.26717
R627 VTAIL.n206 VTAIL.n193 4.26717
R628 VTAIL.n442 VTAIL.n426 3.49141
R629 VTAIL.n468 VTAIL.n467 3.49141
R630 VTAIL.n30 VTAIL.n14 3.49141
R631 VTAIL.n56 VTAIL.n55 3.49141
R632 VTAIL.n88 VTAIL.n72 3.49141
R633 VTAIL.n114 VTAIL.n113 3.49141
R634 VTAIL.n148 VTAIL.n132 3.49141
R635 VTAIL.n174 VTAIL.n173 3.49141
R636 VTAIL.n410 VTAIL.n409 3.49141
R637 VTAIL.n385 VTAIL.n369 3.49141
R638 VTAIL.n350 VTAIL.n349 3.49141
R639 VTAIL.n325 VTAIL.n309 3.49141
R640 VTAIL.n292 VTAIL.n291 3.49141
R641 VTAIL.n267 VTAIL.n251 3.49141
R642 VTAIL.n232 VTAIL.n231 3.49141
R643 VTAIL.n207 VTAIL.n191 3.49141
R644 VTAIL.n435 VTAIL.n431 2.84303
R645 VTAIL.n23 VTAIL.n19 2.84303
R646 VTAIL.n81 VTAIL.n77 2.84303
R647 VTAIL.n141 VTAIL.n137 2.84303
R648 VTAIL.n378 VTAIL.n374 2.84303
R649 VTAIL.n318 VTAIL.n314 2.84303
R650 VTAIL.n260 VTAIL.n256 2.84303
R651 VTAIL.n200 VTAIL.n196 2.84303
R652 VTAIL.n446 VTAIL.n445 2.71565
R653 VTAIL.n464 VTAIL.n416 2.71565
R654 VTAIL.n34 VTAIL.n33 2.71565
R655 VTAIL.n52 VTAIL.n4 2.71565
R656 VTAIL.n92 VTAIL.n91 2.71565
R657 VTAIL.n110 VTAIL.n62 2.71565
R658 VTAIL.n152 VTAIL.n151 2.71565
R659 VTAIL.n170 VTAIL.n122 2.71565
R660 VTAIL.n406 VTAIL.n358 2.71565
R661 VTAIL.n389 VTAIL.n388 2.71565
R662 VTAIL.n346 VTAIL.n298 2.71565
R663 VTAIL.n329 VTAIL.n328 2.71565
R664 VTAIL.n288 VTAIL.n240 2.71565
R665 VTAIL.n271 VTAIL.n270 2.71565
R666 VTAIL.n228 VTAIL.n180 2.71565
R667 VTAIL.n211 VTAIL.n210 2.71565
R668 VTAIL.n237 VTAIL.n235 2.19878
R669 VTAIL.n295 VTAIL.n237 2.19878
R670 VTAIL.n355 VTAIL.n353 2.19878
R671 VTAIL.n413 VTAIL.n355 2.19878
R672 VTAIL.n177 VTAIL.n119 2.19878
R673 VTAIL.n119 VTAIL.n117 2.19878
R674 VTAIL.n59 VTAIL.n1 2.19878
R675 VTAIL VTAIL.n471 2.14059
R676 VTAIL.n450 VTAIL.n424 1.93989
R677 VTAIL.n463 VTAIL.n418 1.93989
R678 VTAIL.n38 VTAIL.n12 1.93989
R679 VTAIL.n51 VTAIL.n6 1.93989
R680 VTAIL.n96 VTAIL.n70 1.93989
R681 VTAIL.n109 VTAIL.n64 1.93989
R682 VTAIL.n156 VTAIL.n130 1.93989
R683 VTAIL.n169 VTAIL.n124 1.93989
R684 VTAIL.n405 VTAIL.n360 1.93989
R685 VTAIL.n392 VTAIL.n366 1.93989
R686 VTAIL.n345 VTAIL.n300 1.93989
R687 VTAIL.n332 VTAIL.n306 1.93989
R688 VTAIL.n287 VTAIL.n242 1.93989
R689 VTAIL.n274 VTAIL.n248 1.93989
R690 VTAIL.n227 VTAIL.n182 1.93989
R691 VTAIL.n214 VTAIL.n188 1.93989
R692 VTAIL.n0 VTAIL.t5 1.83723
R693 VTAIL.n0 VTAIL.t2 1.83723
R694 VTAIL.n118 VTAIL.t8 1.83723
R695 VTAIL.n118 VTAIL.t11 1.83723
R696 VTAIL.n354 VTAIL.t13 1.83723
R697 VTAIL.n354 VTAIL.t9 1.83723
R698 VTAIL.n236 VTAIL.t7 1.83723
R699 VTAIL.n236 VTAIL.t3 1.83723
R700 VTAIL.n451 VTAIL.n422 1.16414
R701 VTAIL.n460 VTAIL.n459 1.16414
R702 VTAIL.n39 VTAIL.n10 1.16414
R703 VTAIL.n48 VTAIL.n47 1.16414
R704 VTAIL.n97 VTAIL.n68 1.16414
R705 VTAIL.n106 VTAIL.n105 1.16414
R706 VTAIL.n157 VTAIL.n128 1.16414
R707 VTAIL.n166 VTAIL.n165 1.16414
R708 VTAIL.n402 VTAIL.n401 1.16414
R709 VTAIL.n393 VTAIL.n364 1.16414
R710 VTAIL.n342 VTAIL.n341 1.16414
R711 VTAIL.n333 VTAIL.n304 1.16414
R712 VTAIL.n284 VTAIL.n283 1.16414
R713 VTAIL.n275 VTAIL.n246 1.16414
R714 VTAIL.n224 VTAIL.n223 1.16414
R715 VTAIL.n215 VTAIL.n186 1.16414
R716 VTAIL.n353 VTAIL.n295 0.470328
R717 VTAIL.n117 VTAIL.n59 0.470328
R718 VTAIL.n455 VTAIL.n454 0.388379
R719 VTAIL.n456 VTAIL.n420 0.388379
R720 VTAIL.n43 VTAIL.n42 0.388379
R721 VTAIL.n44 VTAIL.n8 0.388379
R722 VTAIL.n101 VTAIL.n100 0.388379
R723 VTAIL.n102 VTAIL.n66 0.388379
R724 VTAIL.n161 VTAIL.n160 0.388379
R725 VTAIL.n162 VTAIL.n126 0.388379
R726 VTAIL.n398 VTAIL.n362 0.388379
R727 VTAIL.n397 VTAIL.n396 0.388379
R728 VTAIL.n338 VTAIL.n302 0.388379
R729 VTAIL.n337 VTAIL.n336 0.388379
R730 VTAIL.n280 VTAIL.n244 0.388379
R731 VTAIL.n279 VTAIL.n278 0.388379
R732 VTAIL.n220 VTAIL.n184 0.388379
R733 VTAIL.n219 VTAIL.n218 0.388379
R734 VTAIL.n436 VTAIL.n435 0.155672
R735 VTAIL.n436 VTAIL.n427 0.155672
R736 VTAIL.n443 VTAIL.n427 0.155672
R737 VTAIL.n444 VTAIL.n443 0.155672
R738 VTAIL.n444 VTAIL.n423 0.155672
R739 VTAIL.n452 VTAIL.n423 0.155672
R740 VTAIL.n453 VTAIL.n452 0.155672
R741 VTAIL.n453 VTAIL.n419 0.155672
R742 VTAIL.n461 VTAIL.n419 0.155672
R743 VTAIL.n462 VTAIL.n461 0.155672
R744 VTAIL.n462 VTAIL.n415 0.155672
R745 VTAIL.n469 VTAIL.n415 0.155672
R746 VTAIL.n24 VTAIL.n23 0.155672
R747 VTAIL.n24 VTAIL.n15 0.155672
R748 VTAIL.n31 VTAIL.n15 0.155672
R749 VTAIL.n32 VTAIL.n31 0.155672
R750 VTAIL.n32 VTAIL.n11 0.155672
R751 VTAIL.n40 VTAIL.n11 0.155672
R752 VTAIL.n41 VTAIL.n40 0.155672
R753 VTAIL.n41 VTAIL.n7 0.155672
R754 VTAIL.n49 VTAIL.n7 0.155672
R755 VTAIL.n50 VTAIL.n49 0.155672
R756 VTAIL.n50 VTAIL.n3 0.155672
R757 VTAIL.n57 VTAIL.n3 0.155672
R758 VTAIL.n82 VTAIL.n81 0.155672
R759 VTAIL.n82 VTAIL.n73 0.155672
R760 VTAIL.n89 VTAIL.n73 0.155672
R761 VTAIL.n90 VTAIL.n89 0.155672
R762 VTAIL.n90 VTAIL.n69 0.155672
R763 VTAIL.n98 VTAIL.n69 0.155672
R764 VTAIL.n99 VTAIL.n98 0.155672
R765 VTAIL.n99 VTAIL.n65 0.155672
R766 VTAIL.n107 VTAIL.n65 0.155672
R767 VTAIL.n108 VTAIL.n107 0.155672
R768 VTAIL.n108 VTAIL.n61 0.155672
R769 VTAIL.n115 VTAIL.n61 0.155672
R770 VTAIL.n142 VTAIL.n141 0.155672
R771 VTAIL.n142 VTAIL.n133 0.155672
R772 VTAIL.n149 VTAIL.n133 0.155672
R773 VTAIL.n150 VTAIL.n149 0.155672
R774 VTAIL.n150 VTAIL.n129 0.155672
R775 VTAIL.n158 VTAIL.n129 0.155672
R776 VTAIL.n159 VTAIL.n158 0.155672
R777 VTAIL.n159 VTAIL.n125 0.155672
R778 VTAIL.n167 VTAIL.n125 0.155672
R779 VTAIL.n168 VTAIL.n167 0.155672
R780 VTAIL.n168 VTAIL.n121 0.155672
R781 VTAIL.n175 VTAIL.n121 0.155672
R782 VTAIL.n411 VTAIL.n357 0.155672
R783 VTAIL.n404 VTAIL.n357 0.155672
R784 VTAIL.n404 VTAIL.n403 0.155672
R785 VTAIL.n403 VTAIL.n361 0.155672
R786 VTAIL.n395 VTAIL.n361 0.155672
R787 VTAIL.n395 VTAIL.n394 0.155672
R788 VTAIL.n394 VTAIL.n365 0.155672
R789 VTAIL.n387 VTAIL.n365 0.155672
R790 VTAIL.n387 VTAIL.n386 0.155672
R791 VTAIL.n386 VTAIL.n370 0.155672
R792 VTAIL.n379 VTAIL.n370 0.155672
R793 VTAIL.n379 VTAIL.n378 0.155672
R794 VTAIL.n351 VTAIL.n297 0.155672
R795 VTAIL.n344 VTAIL.n297 0.155672
R796 VTAIL.n344 VTAIL.n343 0.155672
R797 VTAIL.n343 VTAIL.n301 0.155672
R798 VTAIL.n335 VTAIL.n301 0.155672
R799 VTAIL.n335 VTAIL.n334 0.155672
R800 VTAIL.n334 VTAIL.n305 0.155672
R801 VTAIL.n327 VTAIL.n305 0.155672
R802 VTAIL.n327 VTAIL.n326 0.155672
R803 VTAIL.n326 VTAIL.n310 0.155672
R804 VTAIL.n319 VTAIL.n310 0.155672
R805 VTAIL.n319 VTAIL.n318 0.155672
R806 VTAIL.n293 VTAIL.n239 0.155672
R807 VTAIL.n286 VTAIL.n239 0.155672
R808 VTAIL.n286 VTAIL.n285 0.155672
R809 VTAIL.n285 VTAIL.n243 0.155672
R810 VTAIL.n277 VTAIL.n243 0.155672
R811 VTAIL.n277 VTAIL.n276 0.155672
R812 VTAIL.n276 VTAIL.n247 0.155672
R813 VTAIL.n269 VTAIL.n247 0.155672
R814 VTAIL.n269 VTAIL.n268 0.155672
R815 VTAIL.n268 VTAIL.n252 0.155672
R816 VTAIL.n261 VTAIL.n252 0.155672
R817 VTAIL.n261 VTAIL.n260 0.155672
R818 VTAIL.n233 VTAIL.n179 0.155672
R819 VTAIL.n226 VTAIL.n179 0.155672
R820 VTAIL.n226 VTAIL.n225 0.155672
R821 VTAIL.n225 VTAIL.n183 0.155672
R822 VTAIL.n217 VTAIL.n183 0.155672
R823 VTAIL.n217 VTAIL.n216 0.155672
R824 VTAIL.n216 VTAIL.n187 0.155672
R825 VTAIL.n209 VTAIL.n187 0.155672
R826 VTAIL.n209 VTAIL.n208 0.155672
R827 VTAIL.n208 VTAIL.n192 0.155672
R828 VTAIL.n201 VTAIL.n192 0.155672
R829 VTAIL.n201 VTAIL.n200 0.155672
R830 VTAIL VTAIL.n1 0.0586897
R831 B.n806 B.n805 585
R832 B.n302 B.n127 585
R833 B.n301 B.n300 585
R834 B.n299 B.n298 585
R835 B.n297 B.n296 585
R836 B.n295 B.n294 585
R837 B.n293 B.n292 585
R838 B.n291 B.n290 585
R839 B.n289 B.n288 585
R840 B.n287 B.n286 585
R841 B.n285 B.n284 585
R842 B.n283 B.n282 585
R843 B.n281 B.n280 585
R844 B.n279 B.n278 585
R845 B.n277 B.n276 585
R846 B.n275 B.n274 585
R847 B.n273 B.n272 585
R848 B.n271 B.n270 585
R849 B.n269 B.n268 585
R850 B.n267 B.n266 585
R851 B.n265 B.n264 585
R852 B.n263 B.n262 585
R853 B.n261 B.n260 585
R854 B.n259 B.n258 585
R855 B.n257 B.n256 585
R856 B.n255 B.n254 585
R857 B.n253 B.n252 585
R858 B.n251 B.n250 585
R859 B.n249 B.n248 585
R860 B.n247 B.n246 585
R861 B.n245 B.n244 585
R862 B.n243 B.n242 585
R863 B.n241 B.n240 585
R864 B.n239 B.n238 585
R865 B.n237 B.n236 585
R866 B.n235 B.n234 585
R867 B.n233 B.n232 585
R868 B.n231 B.n230 585
R869 B.n229 B.n228 585
R870 B.n227 B.n226 585
R871 B.n225 B.n224 585
R872 B.n223 B.n222 585
R873 B.n221 B.n220 585
R874 B.n219 B.n218 585
R875 B.n217 B.n216 585
R876 B.n215 B.n214 585
R877 B.n213 B.n212 585
R878 B.n211 B.n210 585
R879 B.n209 B.n208 585
R880 B.n207 B.n206 585
R881 B.n205 B.n204 585
R882 B.n203 B.n202 585
R883 B.n201 B.n200 585
R884 B.n199 B.n198 585
R885 B.n197 B.n196 585
R886 B.n195 B.n194 585
R887 B.n193 B.n192 585
R888 B.n191 B.n190 585
R889 B.n189 B.n188 585
R890 B.n187 B.n186 585
R891 B.n185 B.n184 585
R892 B.n183 B.n182 585
R893 B.n181 B.n180 585
R894 B.n179 B.n178 585
R895 B.n177 B.n176 585
R896 B.n175 B.n174 585
R897 B.n173 B.n172 585
R898 B.n171 B.n170 585
R899 B.n169 B.n168 585
R900 B.n167 B.n166 585
R901 B.n165 B.n164 585
R902 B.n163 B.n162 585
R903 B.n161 B.n160 585
R904 B.n159 B.n158 585
R905 B.n157 B.n156 585
R906 B.n155 B.n154 585
R907 B.n153 B.n152 585
R908 B.n151 B.n150 585
R909 B.n149 B.n148 585
R910 B.n147 B.n146 585
R911 B.n145 B.n144 585
R912 B.n143 B.n142 585
R913 B.n141 B.n140 585
R914 B.n139 B.n138 585
R915 B.n137 B.n136 585
R916 B.n135 B.n134 585
R917 B.n804 B.n84 585
R918 B.n809 B.n84 585
R919 B.n803 B.n83 585
R920 B.n810 B.n83 585
R921 B.n802 B.n801 585
R922 B.n801 B.n79 585
R923 B.n800 B.n78 585
R924 B.n816 B.n78 585
R925 B.n799 B.n77 585
R926 B.n817 B.n77 585
R927 B.n798 B.n76 585
R928 B.n818 B.n76 585
R929 B.n797 B.n796 585
R930 B.n796 B.n75 585
R931 B.n795 B.n71 585
R932 B.n824 B.n71 585
R933 B.n794 B.n70 585
R934 B.n825 B.n70 585
R935 B.n793 B.n69 585
R936 B.n826 B.n69 585
R937 B.n792 B.n791 585
R938 B.n791 B.n65 585
R939 B.n790 B.n64 585
R940 B.n832 B.n64 585
R941 B.n789 B.n63 585
R942 B.n833 B.n63 585
R943 B.n788 B.n62 585
R944 B.n834 B.n62 585
R945 B.n787 B.n786 585
R946 B.n786 B.n58 585
R947 B.n785 B.n57 585
R948 B.n840 B.n57 585
R949 B.n784 B.n56 585
R950 B.n841 B.n56 585
R951 B.n783 B.n55 585
R952 B.n842 B.n55 585
R953 B.n782 B.n781 585
R954 B.n781 B.n51 585
R955 B.n780 B.n50 585
R956 B.n848 B.n50 585
R957 B.n779 B.n49 585
R958 B.n849 B.n49 585
R959 B.n778 B.n48 585
R960 B.n850 B.n48 585
R961 B.n777 B.n776 585
R962 B.n776 B.n44 585
R963 B.n775 B.n43 585
R964 B.n856 B.n43 585
R965 B.n774 B.n42 585
R966 B.n857 B.n42 585
R967 B.n773 B.n41 585
R968 B.n858 B.n41 585
R969 B.n772 B.n771 585
R970 B.n771 B.n37 585
R971 B.n770 B.n36 585
R972 B.n864 B.n36 585
R973 B.n769 B.n35 585
R974 B.n865 B.n35 585
R975 B.n768 B.n34 585
R976 B.n866 B.n34 585
R977 B.n767 B.n766 585
R978 B.n766 B.n30 585
R979 B.n765 B.n29 585
R980 B.n872 B.n29 585
R981 B.n764 B.n28 585
R982 B.n873 B.n28 585
R983 B.n763 B.n27 585
R984 B.n874 B.n27 585
R985 B.n762 B.n761 585
R986 B.n761 B.n23 585
R987 B.n760 B.n22 585
R988 B.n880 B.n22 585
R989 B.n759 B.n21 585
R990 B.n881 B.n21 585
R991 B.n758 B.n20 585
R992 B.n882 B.n20 585
R993 B.n757 B.n756 585
R994 B.n756 B.n16 585
R995 B.n755 B.n15 585
R996 B.n888 B.n15 585
R997 B.n754 B.n14 585
R998 B.n889 B.n14 585
R999 B.n753 B.n13 585
R1000 B.n890 B.n13 585
R1001 B.n752 B.n751 585
R1002 B.n751 B.n12 585
R1003 B.n750 B.n749 585
R1004 B.n750 B.n8 585
R1005 B.n748 B.n7 585
R1006 B.n897 B.n7 585
R1007 B.n747 B.n6 585
R1008 B.n898 B.n6 585
R1009 B.n746 B.n5 585
R1010 B.n899 B.n5 585
R1011 B.n745 B.n744 585
R1012 B.n744 B.n4 585
R1013 B.n743 B.n303 585
R1014 B.n743 B.n742 585
R1015 B.n733 B.n304 585
R1016 B.n305 B.n304 585
R1017 B.n735 B.n734 585
R1018 B.n736 B.n735 585
R1019 B.n732 B.n309 585
R1020 B.n313 B.n309 585
R1021 B.n731 B.n730 585
R1022 B.n730 B.n729 585
R1023 B.n311 B.n310 585
R1024 B.n312 B.n311 585
R1025 B.n722 B.n721 585
R1026 B.n723 B.n722 585
R1027 B.n720 B.n318 585
R1028 B.n318 B.n317 585
R1029 B.n719 B.n718 585
R1030 B.n718 B.n717 585
R1031 B.n320 B.n319 585
R1032 B.n321 B.n320 585
R1033 B.n710 B.n709 585
R1034 B.n711 B.n710 585
R1035 B.n708 B.n325 585
R1036 B.n329 B.n325 585
R1037 B.n707 B.n706 585
R1038 B.n706 B.n705 585
R1039 B.n327 B.n326 585
R1040 B.n328 B.n327 585
R1041 B.n698 B.n697 585
R1042 B.n699 B.n698 585
R1043 B.n696 B.n334 585
R1044 B.n334 B.n333 585
R1045 B.n695 B.n694 585
R1046 B.n694 B.n693 585
R1047 B.n336 B.n335 585
R1048 B.n337 B.n336 585
R1049 B.n686 B.n685 585
R1050 B.n687 B.n686 585
R1051 B.n684 B.n342 585
R1052 B.n342 B.n341 585
R1053 B.n683 B.n682 585
R1054 B.n682 B.n681 585
R1055 B.n344 B.n343 585
R1056 B.n345 B.n344 585
R1057 B.n674 B.n673 585
R1058 B.n675 B.n674 585
R1059 B.n672 B.n350 585
R1060 B.n350 B.n349 585
R1061 B.n671 B.n670 585
R1062 B.n670 B.n669 585
R1063 B.n352 B.n351 585
R1064 B.n353 B.n352 585
R1065 B.n662 B.n661 585
R1066 B.n663 B.n662 585
R1067 B.n660 B.n358 585
R1068 B.n358 B.n357 585
R1069 B.n659 B.n658 585
R1070 B.n658 B.n657 585
R1071 B.n360 B.n359 585
R1072 B.n361 B.n360 585
R1073 B.n650 B.n649 585
R1074 B.n651 B.n650 585
R1075 B.n648 B.n366 585
R1076 B.n366 B.n365 585
R1077 B.n647 B.n646 585
R1078 B.n646 B.n645 585
R1079 B.n368 B.n367 585
R1080 B.n369 B.n368 585
R1081 B.n638 B.n637 585
R1082 B.n639 B.n638 585
R1083 B.n636 B.n374 585
R1084 B.n374 B.n373 585
R1085 B.n635 B.n634 585
R1086 B.n634 B.n633 585
R1087 B.n376 B.n375 585
R1088 B.n626 B.n376 585
R1089 B.n625 B.n624 585
R1090 B.n627 B.n625 585
R1091 B.n623 B.n381 585
R1092 B.n381 B.n380 585
R1093 B.n622 B.n621 585
R1094 B.n621 B.n620 585
R1095 B.n383 B.n382 585
R1096 B.n384 B.n383 585
R1097 B.n613 B.n612 585
R1098 B.n614 B.n613 585
R1099 B.n611 B.n389 585
R1100 B.n389 B.n388 585
R1101 B.n606 B.n605 585
R1102 B.n604 B.n434 585
R1103 B.n603 B.n433 585
R1104 B.n608 B.n433 585
R1105 B.n602 B.n601 585
R1106 B.n600 B.n599 585
R1107 B.n598 B.n597 585
R1108 B.n596 B.n595 585
R1109 B.n594 B.n593 585
R1110 B.n592 B.n591 585
R1111 B.n590 B.n589 585
R1112 B.n588 B.n587 585
R1113 B.n586 B.n585 585
R1114 B.n584 B.n583 585
R1115 B.n582 B.n581 585
R1116 B.n580 B.n579 585
R1117 B.n578 B.n577 585
R1118 B.n576 B.n575 585
R1119 B.n574 B.n573 585
R1120 B.n572 B.n571 585
R1121 B.n570 B.n569 585
R1122 B.n568 B.n567 585
R1123 B.n566 B.n565 585
R1124 B.n564 B.n563 585
R1125 B.n562 B.n561 585
R1126 B.n560 B.n559 585
R1127 B.n558 B.n557 585
R1128 B.n556 B.n555 585
R1129 B.n554 B.n553 585
R1130 B.n552 B.n551 585
R1131 B.n550 B.n549 585
R1132 B.n548 B.n547 585
R1133 B.n546 B.n545 585
R1134 B.n544 B.n543 585
R1135 B.n542 B.n541 585
R1136 B.n540 B.n539 585
R1137 B.n538 B.n537 585
R1138 B.n536 B.n535 585
R1139 B.n534 B.n533 585
R1140 B.n531 B.n530 585
R1141 B.n529 B.n528 585
R1142 B.n527 B.n526 585
R1143 B.n525 B.n524 585
R1144 B.n523 B.n522 585
R1145 B.n521 B.n520 585
R1146 B.n519 B.n518 585
R1147 B.n517 B.n516 585
R1148 B.n515 B.n514 585
R1149 B.n513 B.n512 585
R1150 B.n510 B.n509 585
R1151 B.n508 B.n507 585
R1152 B.n506 B.n505 585
R1153 B.n504 B.n503 585
R1154 B.n502 B.n501 585
R1155 B.n500 B.n499 585
R1156 B.n498 B.n497 585
R1157 B.n496 B.n495 585
R1158 B.n494 B.n493 585
R1159 B.n492 B.n491 585
R1160 B.n490 B.n489 585
R1161 B.n488 B.n487 585
R1162 B.n486 B.n485 585
R1163 B.n484 B.n483 585
R1164 B.n482 B.n481 585
R1165 B.n480 B.n479 585
R1166 B.n478 B.n477 585
R1167 B.n476 B.n475 585
R1168 B.n474 B.n473 585
R1169 B.n472 B.n471 585
R1170 B.n470 B.n469 585
R1171 B.n468 B.n467 585
R1172 B.n466 B.n465 585
R1173 B.n464 B.n463 585
R1174 B.n462 B.n461 585
R1175 B.n460 B.n459 585
R1176 B.n458 B.n457 585
R1177 B.n456 B.n455 585
R1178 B.n454 B.n453 585
R1179 B.n452 B.n451 585
R1180 B.n450 B.n449 585
R1181 B.n448 B.n447 585
R1182 B.n446 B.n445 585
R1183 B.n444 B.n443 585
R1184 B.n442 B.n441 585
R1185 B.n440 B.n439 585
R1186 B.n391 B.n390 585
R1187 B.n610 B.n609 585
R1188 B.n609 B.n608 585
R1189 B.n387 B.n386 585
R1190 B.n388 B.n387 585
R1191 B.n616 B.n615 585
R1192 B.n615 B.n614 585
R1193 B.n617 B.n385 585
R1194 B.n385 B.n384 585
R1195 B.n619 B.n618 585
R1196 B.n620 B.n619 585
R1197 B.n379 B.n378 585
R1198 B.n380 B.n379 585
R1199 B.n629 B.n628 585
R1200 B.n628 B.n627 585
R1201 B.n630 B.n377 585
R1202 B.n626 B.n377 585
R1203 B.n632 B.n631 585
R1204 B.n633 B.n632 585
R1205 B.n372 B.n371 585
R1206 B.n373 B.n372 585
R1207 B.n641 B.n640 585
R1208 B.n640 B.n639 585
R1209 B.n642 B.n370 585
R1210 B.n370 B.n369 585
R1211 B.n644 B.n643 585
R1212 B.n645 B.n644 585
R1213 B.n364 B.n363 585
R1214 B.n365 B.n364 585
R1215 B.n653 B.n652 585
R1216 B.n652 B.n651 585
R1217 B.n654 B.n362 585
R1218 B.n362 B.n361 585
R1219 B.n656 B.n655 585
R1220 B.n657 B.n656 585
R1221 B.n356 B.n355 585
R1222 B.n357 B.n356 585
R1223 B.n665 B.n664 585
R1224 B.n664 B.n663 585
R1225 B.n666 B.n354 585
R1226 B.n354 B.n353 585
R1227 B.n668 B.n667 585
R1228 B.n669 B.n668 585
R1229 B.n348 B.n347 585
R1230 B.n349 B.n348 585
R1231 B.n677 B.n676 585
R1232 B.n676 B.n675 585
R1233 B.n678 B.n346 585
R1234 B.n346 B.n345 585
R1235 B.n680 B.n679 585
R1236 B.n681 B.n680 585
R1237 B.n340 B.n339 585
R1238 B.n341 B.n340 585
R1239 B.n689 B.n688 585
R1240 B.n688 B.n687 585
R1241 B.n690 B.n338 585
R1242 B.n338 B.n337 585
R1243 B.n692 B.n691 585
R1244 B.n693 B.n692 585
R1245 B.n332 B.n331 585
R1246 B.n333 B.n332 585
R1247 B.n701 B.n700 585
R1248 B.n700 B.n699 585
R1249 B.n702 B.n330 585
R1250 B.n330 B.n328 585
R1251 B.n704 B.n703 585
R1252 B.n705 B.n704 585
R1253 B.n324 B.n323 585
R1254 B.n329 B.n324 585
R1255 B.n713 B.n712 585
R1256 B.n712 B.n711 585
R1257 B.n714 B.n322 585
R1258 B.n322 B.n321 585
R1259 B.n716 B.n715 585
R1260 B.n717 B.n716 585
R1261 B.n316 B.n315 585
R1262 B.n317 B.n316 585
R1263 B.n725 B.n724 585
R1264 B.n724 B.n723 585
R1265 B.n726 B.n314 585
R1266 B.n314 B.n312 585
R1267 B.n728 B.n727 585
R1268 B.n729 B.n728 585
R1269 B.n308 B.n307 585
R1270 B.n313 B.n308 585
R1271 B.n738 B.n737 585
R1272 B.n737 B.n736 585
R1273 B.n739 B.n306 585
R1274 B.n306 B.n305 585
R1275 B.n741 B.n740 585
R1276 B.n742 B.n741 585
R1277 B.n3 B.n0 585
R1278 B.n4 B.n3 585
R1279 B.n896 B.n1 585
R1280 B.n897 B.n896 585
R1281 B.n895 B.n894 585
R1282 B.n895 B.n8 585
R1283 B.n893 B.n9 585
R1284 B.n12 B.n9 585
R1285 B.n892 B.n891 585
R1286 B.n891 B.n890 585
R1287 B.n11 B.n10 585
R1288 B.n889 B.n11 585
R1289 B.n887 B.n886 585
R1290 B.n888 B.n887 585
R1291 B.n885 B.n17 585
R1292 B.n17 B.n16 585
R1293 B.n884 B.n883 585
R1294 B.n883 B.n882 585
R1295 B.n19 B.n18 585
R1296 B.n881 B.n19 585
R1297 B.n879 B.n878 585
R1298 B.n880 B.n879 585
R1299 B.n877 B.n24 585
R1300 B.n24 B.n23 585
R1301 B.n876 B.n875 585
R1302 B.n875 B.n874 585
R1303 B.n26 B.n25 585
R1304 B.n873 B.n26 585
R1305 B.n871 B.n870 585
R1306 B.n872 B.n871 585
R1307 B.n869 B.n31 585
R1308 B.n31 B.n30 585
R1309 B.n868 B.n867 585
R1310 B.n867 B.n866 585
R1311 B.n33 B.n32 585
R1312 B.n865 B.n33 585
R1313 B.n863 B.n862 585
R1314 B.n864 B.n863 585
R1315 B.n861 B.n38 585
R1316 B.n38 B.n37 585
R1317 B.n860 B.n859 585
R1318 B.n859 B.n858 585
R1319 B.n40 B.n39 585
R1320 B.n857 B.n40 585
R1321 B.n855 B.n854 585
R1322 B.n856 B.n855 585
R1323 B.n853 B.n45 585
R1324 B.n45 B.n44 585
R1325 B.n852 B.n851 585
R1326 B.n851 B.n850 585
R1327 B.n47 B.n46 585
R1328 B.n849 B.n47 585
R1329 B.n847 B.n846 585
R1330 B.n848 B.n847 585
R1331 B.n845 B.n52 585
R1332 B.n52 B.n51 585
R1333 B.n844 B.n843 585
R1334 B.n843 B.n842 585
R1335 B.n54 B.n53 585
R1336 B.n841 B.n54 585
R1337 B.n839 B.n838 585
R1338 B.n840 B.n839 585
R1339 B.n837 B.n59 585
R1340 B.n59 B.n58 585
R1341 B.n836 B.n835 585
R1342 B.n835 B.n834 585
R1343 B.n61 B.n60 585
R1344 B.n833 B.n61 585
R1345 B.n831 B.n830 585
R1346 B.n832 B.n831 585
R1347 B.n829 B.n66 585
R1348 B.n66 B.n65 585
R1349 B.n828 B.n827 585
R1350 B.n827 B.n826 585
R1351 B.n68 B.n67 585
R1352 B.n825 B.n68 585
R1353 B.n823 B.n822 585
R1354 B.n824 B.n823 585
R1355 B.n821 B.n72 585
R1356 B.n75 B.n72 585
R1357 B.n820 B.n819 585
R1358 B.n819 B.n818 585
R1359 B.n74 B.n73 585
R1360 B.n817 B.n74 585
R1361 B.n815 B.n814 585
R1362 B.n816 B.n815 585
R1363 B.n813 B.n80 585
R1364 B.n80 B.n79 585
R1365 B.n812 B.n811 585
R1366 B.n811 B.n810 585
R1367 B.n82 B.n81 585
R1368 B.n809 B.n82 585
R1369 B.n900 B.n899 585
R1370 B.n898 B.n2 585
R1371 B.n134 B.n82 487.695
R1372 B.n806 B.n84 487.695
R1373 B.n609 B.n389 487.695
R1374 B.n606 B.n387 487.695
R1375 B.n131 B.t12 324.418
R1376 B.n128 B.t16 324.418
R1377 B.n437 B.t8 324.418
R1378 B.n435 B.t19 324.418
R1379 B.n128 B.t17 310.753
R1380 B.n437 B.t11 310.753
R1381 B.n131 B.t14 310.753
R1382 B.n435 B.t21 310.753
R1383 B.n129 B.t18 261.298
R1384 B.n438 B.t10 261.298
R1385 B.n132 B.t15 261.298
R1386 B.n436 B.t20 261.298
R1387 B.n808 B.n807 256.663
R1388 B.n808 B.n126 256.663
R1389 B.n808 B.n125 256.663
R1390 B.n808 B.n124 256.663
R1391 B.n808 B.n123 256.663
R1392 B.n808 B.n122 256.663
R1393 B.n808 B.n121 256.663
R1394 B.n808 B.n120 256.663
R1395 B.n808 B.n119 256.663
R1396 B.n808 B.n118 256.663
R1397 B.n808 B.n117 256.663
R1398 B.n808 B.n116 256.663
R1399 B.n808 B.n115 256.663
R1400 B.n808 B.n114 256.663
R1401 B.n808 B.n113 256.663
R1402 B.n808 B.n112 256.663
R1403 B.n808 B.n111 256.663
R1404 B.n808 B.n110 256.663
R1405 B.n808 B.n109 256.663
R1406 B.n808 B.n108 256.663
R1407 B.n808 B.n107 256.663
R1408 B.n808 B.n106 256.663
R1409 B.n808 B.n105 256.663
R1410 B.n808 B.n104 256.663
R1411 B.n808 B.n103 256.663
R1412 B.n808 B.n102 256.663
R1413 B.n808 B.n101 256.663
R1414 B.n808 B.n100 256.663
R1415 B.n808 B.n99 256.663
R1416 B.n808 B.n98 256.663
R1417 B.n808 B.n97 256.663
R1418 B.n808 B.n96 256.663
R1419 B.n808 B.n95 256.663
R1420 B.n808 B.n94 256.663
R1421 B.n808 B.n93 256.663
R1422 B.n808 B.n92 256.663
R1423 B.n808 B.n91 256.663
R1424 B.n808 B.n90 256.663
R1425 B.n808 B.n89 256.663
R1426 B.n808 B.n88 256.663
R1427 B.n808 B.n87 256.663
R1428 B.n808 B.n86 256.663
R1429 B.n808 B.n85 256.663
R1430 B.n608 B.n607 256.663
R1431 B.n608 B.n392 256.663
R1432 B.n608 B.n393 256.663
R1433 B.n608 B.n394 256.663
R1434 B.n608 B.n395 256.663
R1435 B.n608 B.n396 256.663
R1436 B.n608 B.n397 256.663
R1437 B.n608 B.n398 256.663
R1438 B.n608 B.n399 256.663
R1439 B.n608 B.n400 256.663
R1440 B.n608 B.n401 256.663
R1441 B.n608 B.n402 256.663
R1442 B.n608 B.n403 256.663
R1443 B.n608 B.n404 256.663
R1444 B.n608 B.n405 256.663
R1445 B.n608 B.n406 256.663
R1446 B.n608 B.n407 256.663
R1447 B.n608 B.n408 256.663
R1448 B.n608 B.n409 256.663
R1449 B.n608 B.n410 256.663
R1450 B.n608 B.n411 256.663
R1451 B.n608 B.n412 256.663
R1452 B.n608 B.n413 256.663
R1453 B.n608 B.n414 256.663
R1454 B.n608 B.n415 256.663
R1455 B.n608 B.n416 256.663
R1456 B.n608 B.n417 256.663
R1457 B.n608 B.n418 256.663
R1458 B.n608 B.n419 256.663
R1459 B.n608 B.n420 256.663
R1460 B.n608 B.n421 256.663
R1461 B.n608 B.n422 256.663
R1462 B.n608 B.n423 256.663
R1463 B.n608 B.n424 256.663
R1464 B.n608 B.n425 256.663
R1465 B.n608 B.n426 256.663
R1466 B.n608 B.n427 256.663
R1467 B.n608 B.n428 256.663
R1468 B.n608 B.n429 256.663
R1469 B.n608 B.n430 256.663
R1470 B.n608 B.n431 256.663
R1471 B.n608 B.n432 256.663
R1472 B.n902 B.n901 256.663
R1473 B.n138 B.n137 163.367
R1474 B.n142 B.n141 163.367
R1475 B.n146 B.n145 163.367
R1476 B.n150 B.n149 163.367
R1477 B.n154 B.n153 163.367
R1478 B.n158 B.n157 163.367
R1479 B.n162 B.n161 163.367
R1480 B.n166 B.n165 163.367
R1481 B.n170 B.n169 163.367
R1482 B.n174 B.n173 163.367
R1483 B.n178 B.n177 163.367
R1484 B.n182 B.n181 163.367
R1485 B.n186 B.n185 163.367
R1486 B.n190 B.n189 163.367
R1487 B.n194 B.n193 163.367
R1488 B.n198 B.n197 163.367
R1489 B.n202 B.n201 163.367
R1490 B.n206 B.n205 163.367
R1491 B.n210 B.n209 163.367
R1492 B.n214 B.n213 163.367
R1493 B.n218 B.n217 163.367
R1494 B.n222 B.n221 163.367
R1495 B.n226 B.n225 163.367
R1496 B.n230 B.n229 163.367
R1497 B.n234 B.n233 163.367
R1498 B.n238 B.n237 163.367
R1499 B.n242 B.n241 163.367
R1500 B.n246 B.n245 163.367
R1501 B.n250 B.n249 163.367
R1502 B.n254 B.n253 163.367
R1503 B.n258 B.n257 163.367
R1504 B.n262 B.n261 163.367
R1505 B.n266 B.n265 163.367
R1506 B.n270 B.n269 163.367
R1507 B.n274 B.n273 163.367
R1508 B.n278 B.n277 163.367
R1509 B.n282 B.n281 163.367
R1510 B.n286 B.n285 163.367
R1511 B.n290 B.n289 163.367
R1512 B.n294 B.n293 163.367
R1513 B.n298 B.n297 163.367
R1514 B.n300 B.n127 163.367
R1515 B.n613 B.n389 163.367
R1516 B.n613 B.n383 163.367
R1517 B.n621 B.n383 163.367
R1518 B.n621 B.n381 163.367
R1519 B.n625 B.n381 163.367
R1520 B.n625 B.n376 163.367
R1521 B.n634 B.n376 163.367
R1522 B.n634 B.n374 163.367
R1523 B.n638 B.n374 163.367
R1524 B.n638 B.n368 163.367
R1525 B.n646 B.n368 163.367
R1526 B.n646 B.n366 163.367
R1527 B.n650 B.n366 163.367
R1528 B.n650 B.n360 163.367
R1529 B.n658 B.n360 163.367
R1530 B.n658 B.n358 163.367
R1531 B.n662 B.n358 163.367
R1532 B.n662 B.n352 163.367
R1533 B.n670 B.n352 163.367
R1534 B.n670 B.n350 163.367
R1535 B.n674 B.n350 163.367
R1536 B.n674 B.n344 163.367
R1537 B.n682 B.n344 163.367
R1538 B.n682 B.n342 163.367
R1539 B.n686 B.n342 163.367
R1540 B.n686 B.n336 163.367
R1541 B.n694 B.n336 163.367
R1542 B.n694 B.n334 163.367
R1543 B.n698 B.n334 163.367
R1544 B.n698 B.n327 163.367
R1545 B.n706 B.n327 163.367
R1546 B.n706 B.n325 163.367
R1547 B.n710 B.n325 163.367
R1548 B.n710 B.n320 163.367
R1549 B.n718 B.n320 163.367
R1550 B.n718 B.n318 163.367
R1551 B.n722 B.n318 163.367
R1552 B.n722 B.n311 163.367
R1553 B.n730 B.n311 163.367
R1554 B.n730 B.n309 163.367
R1555 B.n735 B.n309 163.367
R1556 B.n735 B.n304 163.367
R1557 B.n743 B.n304 163.367
R1558 B.n744 B.n743 163.367
R1559 B.n744 B.n5 163.367
R1560 B.n6 B.n5 163.367
R1561 B.n7 B.n6 163.367
R1562 B.n750 B.n7 163.367
R1563 B.n751 B.n750 163.367
R1564 B.n751 B.n13 163.367
R1565 B.n14 B.n13 163.367
R1566 B.n15 B.n14 163.367
R1567 B.n756 B.n15 163.367
R1568 B.n756 B.n20 163.367
R1569 B.n21 B.n20 163.367
R1570 B.n22 B.n21 163.367
R1571 B.n761 B.n22 163.367
R1572 B.n761 B.n27 163.367
R1573 B.n28 B.n27 163.367
R1574 B.n29 B.n28 163.367
R1575 B.n766 B.n29 163.367
R1576 B.n766 B.n34 163.367
R1577 B.n35 B.n34 163.367
R1578 B.n36 B.n35 163.367
R1579 B.n771 B.n36 163.367
R1580 B.n771 B.n41 163.367
R1581 B.n42 B.n41 163.367
R1582 B.n43 B.n42 163.367
R1583 B.n776 B.n43 163.367
R1584 B.n776 B.n48 163.367
R1585 B.n49 B.n48 163.367
R1586 B.n50 B.n49 163.367
R1587 B.n781 B.n50 163.367
R1588 B.n781 B.n55 163.367
R1589 B.n56 B.n55 163.367
R1590 B.n57 B.n56 163.367
R1591 B.n786 B.n57 163.367
R1592 B.n786 B.n62 163.367
R1593 B.n63 B.n62 163.367
R1594 B.n64 B.n63 163.367
R1595 B.n791 B.n64 163.367
R1596 B.n791 B.n69 163.367
R1597 B.n70 B.n69 163.367
R1598 B.n71 B.n70 163.367
R1599 B.n796 B.n71 163.367
R1600 B.n796 B.n76 163.367
R1601 B.n77 B.n76 163.367
R1602 B.n78 B.n77 163.367
R1603 B.n801 B.n78 163.367
R1604 B.n801 B.n83 163.367
R1605 B.n84 B.n83 163.367
R1606 B.n434 B.n433 163.367
R1607 B.n601 B.n433 163.367
R1608 B.n599 B.n598 163.367
R1609 B.n595 B.n594 163.367
R1610 B.n591 B.n590 163.367
R1611 B.n587 B.n586 163.367
R1612 B.n583 B.n582 163.367
R1613 B.n579 B.n578 163.367
R1614 B.n575 B.n574 163.367
R1615 B.n571 B.n570 163.367
R1616 B.n567 B.n566 163.367
R1617 B.n563 B.n562 163.367
R1618 B.n559 B.n558 163.367
R1619 B.n555 B.n554 163.367
R1620 B.n551 B.n550 163.367
R1621 B.n547 B.n546 163.367
R1622 B.n543 B.n542 163.367
R1623 B.n539 B.n538 163.367
R1624 B.n535 B.n534 163.367
R1625 B.n530 B.n529 163.367
R1626 B.n526 B.n525 163.367
R1627 B.n522 B.n521 163.367
R1628 B.n518 B.n517 163.367
R1629 B.n514 B.n513 163.367
R1630 B.n509 B.n508 163.367
R1631 B.n505 B.n504 163.367
R1632 B.n501 B.n500 163.367
R1633 B.n497 B.n496 163.367
R1634 B.n493 B.n492 163.367
R1635 B.n489 B.n488 163.367
R1636 B.n485 B.n484 163.367
R1637 B.n481 B.n480 163.367
R1638 B.n477 B.n476 163.367
R1639 B.n473 B.n472 163.367
R1640 B.n469 B.n468 163.367
R1641 B.n465 B.n464 163.367
R1642 B.n461 B.n460 163.367
R1643 B.n457 B.n456 163.367
R1644 B.n453 B.n452 163.367
R1645 B.n449 B.n448 163.367
R1646 B.n445 B.n444 163.367
R1647 B.n441 B.n440 163.367
R1648 B.n609 B.n391 163.367
R1649 B.n615 B.n387 163.367
R1650 B.n615 B.n385 163.367
R1651 B.n619 B.n385 163.367
R1652 B.n619 B.n379 163.367
R1653 B.n628 B.n379 163.367
R1654 B.n628 B.n377 163.367
R1655 B.n632 B.n377 163.367
R1656 B.n632 B.n372 163.367
R1657 B.n640 B.n372 163.367
R1658 B.n640 B.n370 163.367
R1659 B.n644 B.n370 163.367
R1660 B.n644 B.n364 163.367
R1661 B.n652 B.n364 163.367
R1662 B.n652 B.n362 163.367
R1663 B.n656 B.n362 163.367
R1664 B.n656 B.n356 163.367
R1665 B.n664 B.n356 163.367
R1666 B.n664 B.n354 163.367
R1667 B.n668 B.n354 163.367
R1668 B.n668 B.n348 163.367
R1669 B.n676 B.n348 163.367
R1670 B.n676 B.n346 163.367
R1671 B.n680 B.n346 163.367
R1672 B.n680 B.n340 163.367
R1673 B.n688 B.n340 163.367
R1674 B.n688 B.n338 163.367
R1675 B.n692 B.n338 163.367
R1676 B.n692 B.n332 163.367
R1677 B.n700 B.n332 163.367
R1678 B.n700 B.n330 163.367
R1679 B.n704 B.n330 163.367
R1680 B.n704 B.n324 163.367
R1681 B.n712 B.n324 163.367
R1682 B.n712 B.n322 163.367
R1683 B.n716 B.n322 163.367
R1684 B.n716 B.n316 163.367
R1685 B.n724 B.n316 163.367
R1686 B.n724 B.n314 163.367
R1687 B.n728 B.n314 163.367
R1688 B.n728 B.n308 163.367
R1689 B.n737 B.n308 163.367
R1690 B.n737 B.n306 163.367
R1691 B.n741 B.n306 163.367
R1692 B.n741 B.n3 163.367
R1693 B.n900 B.n3 163.367
R1694 B.n896 B.n2 163.367
R1695 B.n896 B.n895 163.367
R1696 B.n895 B.n9 163.367
R1697 B.n891 B.n9 163.367
R1698 B.n891 B.n11 163.367
R1699 B.n887 B.n11 163.367
R1700 B.n887 B.n17 163.367
R1701 B.n883 B.n17 163.367
R1702 B.n883 B.n19 163.367
R1703 B.n879 B.n19 163.367
R1704 B.n879 B.n24 163.367
R1705 B.n875 B.n24 163.367
R1706 B.n875 B.n26 163.367
R1707 B.n871 B.n26 163.367
R1708 B.n871 B.n31 163.367
R1709 B.n867 B.n31 163.367
R1710 B.n867 B.n33 163.367
R1711 B.n863 B.n33 163.367
R1712 B.n863 B.n38 163.367
R1713 B.n859 B.n38 163.367
R1714 B.n859 B.n40 163.367
R1715 B.n855 B.n40 163.367
R1716 B.n855 B.n45 163.367
R1717 B.n851 B.n45 163.367
R1718 B.n851 B.n47 163.367
R1719 B.n847 B.n47 163.367
R1720 B.n847 B.n52 163.367
R1721 B.n843 B.n52 163.367
R1722 B.n843 B.n54 163.367
R1723 B.n839 B.n54 163.367
R1724 B.n839 B.n59 163.367
R1725 B.n835 B.n59 163.367
R1726 B.n835 B.n61 163.367
R1727 B.n831 B.n61 163.367
R1728 B.n831 B.n66 163.367
R1729 B.n827 B.n66 163.367
R1730 B.n827 B.n68 163.367
R1731 B.n823 B.n68 163.367
R1732 B.n823 B.n72 163.367
R1733 B.n819 B.n72 163.367
R1734 B.n819 B.n74 163.367
R1735 B.n815 B.n74 163.367
R1736 B.n815 B.n80 163.367
R1737 B.n811 B.n80 163.367
R1738 B.n811 B.n82 163.367
R1739 B.n608 B.n388 89.7545
R1740 B.n809 B.n808 89.7545
R1741 B.n134 B.n85 71.676
R1742 B.n138 B.n86 71.676
R1743 B.n142 B.n87 71.676
R1744 B.n146 B.n88 71.676
R1745 B.n150 B.n89 71.676
R1746 B.n154 B.n90 71.676
R1747 B.n158 B.n91 71.676
R1748 B.n162 B.n92 71.676
R1749 B.n166 B.n93 71.676
R1750 B.n170 B.n94 71.676
R1751 B.n174 B.n95 71.676
R1752 B.n178 B.n96 71.676
R1753 B.n182 B.n97 71.676
R1754 B.n186 B.n98 71.676
R1755 B.n190 B.n99 71.676
R1756 B.n194 B.n100 71.676
R1757 B.n198 B.n101 71.676
R1758 B.n202 B.n102 71.676
R1759 B.n206 B.n103 71.676
R1760 B.n210 B.n104 71.676
R1761 B.n214 B.n105 71.676
R1762 B.n218 B.n106 71.676
R1763 B.n222 B.n107 71.676
R1764 B.n226 B.n108 71.676
R1765 B.n230 B.n109 71.676
R1766 B.n234 B.n110 71.676
R1767 B.n238 B.n111 71.676
R1768 B.n242 B.n112 71.676
R1769 B.n246 B.n113 71.676
R1770 B.n250 B.n114 71.676
R1771 B.n254 B.n115 71.676
R1772 B.n258 B.n116 71.676
R1773 B.n262 B.n117 71.676
R1774 B.n266 B.n118 71.676
R1775 B.n270 B.n119 71.676
R1776 B.n274 B.n120 71.676
R1777 B.n278 B.n121 71.676
R1778 B.n282 B.n122 71.676
R1779 B.n286 B.n123 71.676
R1780 B.n290 B.n124 71.676
R1781 B.n294 B.n125 71.676
R1782 B.n298 B.n126 71.676
R1783 B.n807 B.n127 71.676
R1784 B.n807 B.n806 71.676
R1785 B.n300 B.n126 71.676
R1786 B.n297 B.n125 71.676
R1787 B.n293 B.n124 71.676
R1788 B.n289 B.n123 71.676
R1789 B.n285 B.n122 71.676
R1790 B.n281 B.n121 71.676
R1791 B.n277 B.n120 71.676
R1792 B.n273 B.n119 71.676
R1793 B.n269 B.n118 71.676
R1794 B.n265 B.n117 71.676
R1795 B.n261 B.n116 71.676
R1796 B.n257 B.n115 71.676
R1797 B.n253 B.n114 71.676
R1798 B.n249 B.n113 71.676
R1799 B.n245 B.n112 71.676
R1800 B.n241 B.n111 71.676
R1801 B.n237 B.n110 71.676
R1802 B.n233 B.n109 71.676
R1803 B.n229 B.n108 71.676
R1804 B.n225 B.n107 71.676
R1805 B.n221 B.n106 71.676
R1806 B.n217 B.n105 71.676
R1807 B.n213 B.n104 71.676
R1808 B.n209 B.n103 71.676
R1809 B.n205 B.n102 71.676
R1810 B.n201 B.n101 71.676
R1811 B.n197 B.n100 71.676
R1812 B.n193 B.n99 71.676
R1813 B.n189 B.n98 71.676
R1814 B.n185 B.n97 71.676
R1815 B.n181 B.n96 71.676
R1816 B.n177 B.n95 71.676
R1817 B.n173 B.n94 71.676
R1818 B.n169 B.n93 71.676
R1819 B.n165 B.n92 71.676
R1820 B.n161 B.n91 71.676
R1821 B.n157 B.n90 71.676
R1822 B.n153 B.n89 71.676
R1823 B.n149 B.n88 71.676
R1824 B.n145 B.n87 71.676
R1825 B.n141 B.n86 71.676
R1826 B.n137 B.n85 71.676
R1827 B.n607 B.n606 71.676
R1828 B.n601 B.n392 71.676
R1829 B.n598 B.n393 71.676
R1830 B.n594 B.n394 71.676
R1831 B.n590 B.n395 71.676
R1832 B.n586 B.n396 71.676
R1833 B.n582 B.n397 71.676
R1834 B.n578 B.n398 71.676
R1835 B.n574 B.n399 71.676
R1836 B.n570 B.n400 71.676
R1837 B.n566 B.n401 71.676
R1838 B.n562 B.n402 71.676
R1839 B.n558 B.n403 71.676
R1840 B.n554 B.n404 71.676
R1841 B.n550 B.n405 71.676
R1842 B.n546 B.n406 71.676
R1843 B.n542 B.n407 71.676
R1844 B.n538 B.n408 71.676
R1845 B.n534 B.n409 71.676
R1846 B.n529 B.n410 71.676
R1847 B.n525 B.n411 71.676
R1848 B.n521 B.n412 71.676
R1849 B.n517 B.n413 71.676
R1850 B.n513 B.n414 71.676
R1851 B.n508 B.n415 71.676
R1852 B.n504 B.n416 71.676
R1853 B.n500 B.n417 71.676
R1854 B.n496 B.n418 71.676
R1855 B.n492 B.n419 71.676
R1856 B.n488 B.n420 71.676
R1857 B.n484 B.n421 71.676
R1858 B.n480 B.n422 71.676
R1859 B.n476 B.n423 71.676
R1860 B.n472 B.n424 71.676
R1861 B.n468 B.n425 71.676
R1862 B.n464 B.n426 71.676
R1863 B.n460 B.n427 71.676
R1864 B.n456 B.n428 71.676
R1865 B.n452 B.n429 71.676
R1866 B.n448 B.n430 71.676
R1867 B.n444 B.n431 71.676
R1868 B.n440 B.n432 71.676
R1869 B.n607 B.n434 71.676
R1870 B.n599 B.n392 71.676
R1871 B.n595 B.n393 71.676
R1872 B.n591 B.n394 71.676
R1873 B.n587 B.n395 71.676
R1874 B.n583 B.n396 71.676
R1875 B.n579 B.n397 71.676
R1876 B.n575 B.n398 71.676
R1877 B.n571 B.n399 71.676
R1878 B.n567 B.n400 71.676
R1879 B.n563 B.n401 71.676
R1880 B.n559 B.n402 71.676
R1881 B.n555 B.n403 71.676
R1882 B.n551 B.n404 71.676
R1883 B.n547 B.n405 71.676
R1884 B.n543 B.n406 71.676
R1885 B.n539 B.n407 71.676
R1886 B.n535 B.n408 71.676
R1887 B.n530 B.n409 71.676
R1888 B.n526 B.n410 71.676
R1889 B.n522 B.n411 71.676
R1890 B.n518 B.n412 71.676
R1891 B.n514 B.n413 71.676
R1892 B.n509 B.n414 71.676
R1893 B.n505 B.n415 71.676
R1894 B.n501 B.n416 71.676
R1895 B.n497 B.n417 71.676
R1896 B.n493 B.n418 71.676
R1897 B.n489 B.n419 71.676
R1898 B.n485 B.n420 71.676
R1899 B.n481 B.n421 71.676
R1900 B.n477 B.n422 71.676
R1901 B.n473 B.n423 71.676
R1902 B.n469 B.n424 71.676
R1903 B.n465 B.n425 71.676
R1904 B.n461 B.n426 71.676
R1905 B.n457 B.n427 71.676
R1906 B.n453 B.n428 71.676
R1907 B.n449 B.n429 71.676
R1908 B.n445 B.n430 71.676
R1909 B.n441 B.n431 71.676
R1910 B.n432 B.n391 71.676
R1911 B.n901 B.n900 71.676
R1912 B.n901 B.n2 71.676
R1913 B.n133 B.n132 59.5399
R1914 B.n130 B.n129 59.5399
R1915 B.n511 B.n438 59.5399
R1916 B.n532 B.n436 59.5399
R1917 B.n132 B.n131 49.455
R1918 B.n129 B.n128 49.455
R1919 B.n438 B.n437 49.455
R1920 B.n436 B.n435 49.455
R1921 B.n614 B.n388 46.5903
R1922 B.n614 B.n384 46.5903
R1923 B.n620 B.n384 46.5903
R1924 B.n620 B.n380 46.5903
R1925 B.n627 B.n380 46.5903
R1926 B.n627 B.n626 46.5903
R1927 B.n633 B.n373 46.5903
R1928 B.n639 B.n373 46.5903
R1929 B.n639 B.n369 46.5903
R1930 B.n645 B.n369 46.5903
R1931 B.n645 B.n365 46.5903
R1932 B.n651 B.n365 46.5903
R1933 B.n651 B.n361 46.5903
R1934 B.n657 B.n361 46.5903
R1935 B.n657 B.n357 46.5903
R1936 B.n663 B.n357 46.5903
R1937 B.n669 B.n353 46.5903
R1938 B.n669 B.n349 46.5903
R1939 B.n675 B.n349 46.5903
R1940 B.n675 B.n345 46.5903
R1941 B.n681 B.n345 46.5903
R1942 B.n681 B.n341 46.5903
R1943 B.n687 B.n341 46.5903
R1944 B.n693 B.n337 46.5903
R1945 B.n693 B.n333 46.5903
R1946 B.n699 B.n333 46.5903
R1947 B.n699 B.n328 46.5903
R1948 B.n705 B.n328 46.5903
R1949 B.n705 B.n329 46.5903
R1950 B.n711 B.n321 46.5903
R1951 B.n717 B.n321 46.5903
R1952 B.n717 B.n317 46.5903
R1953 B.n723 B.n317 46.5903
R1954 B.n723 B.n312 46.5903
R1955 B.n729 B.n312 46.5903
R1956 B.n729 B.n313 46.5903
R1957 B.n736 B.n305 46.5903
R1958 B.n742 B.n305 46.5903
R1959 B.n742 B.n4 46.5903
R1960 B.n899 B.n4 46.5903
R1961 B.n899 B.n898 46.5903
R1962 B.n898 B.n897 46.5903
R1963 B.n897 B.n8 46.5903
R1964 B.n12 B.n8 46.5903
R1965 B.n890 B.n12 46.5903
R1966 B.n889 B.n888 46.5903
R1967 B.n888 B.n16 46.5903
R1968 B.n882 B.n16 46.5903
R1969 B.n882 B.n881 46.5903
R1970 B.n881 B.n880 46.5903
R1971 B.n880 B.n23 46.5903
R1972 B.n874 B.n23 46.5903
R1973 B.n873 B.n872 46.5903
R1974 B.n872 B.n30 46.5903
R1975 B.n866 B.n30 46.5903
R1976 B.n866 B.n865 46.5903
R1977 B.n865 B.n864 46.5903
R1978 B.n864 B.n37 46.5903
R1979 B.n858 B.n857 46.5903
R1980 B.n857 B.n856 46.5903
R1981 B.n856 B.n44 46.5903
R1982 B.n850 B.n44 46.5903
R1983 B.n850 B.n849 46.5903
R1984 B.n849 B.n848 46.5903
R1985 B.n848 B.n51 46.5903
R1986 B.n842 B.n841 46.5903
R1987 B.n841 B.n840 46.5903
R1988 B.n840 B.n58 46.5903
R1989 B.n834 B.n58 46.5903
R1990 B.n834 B.n833 46.5903
R1991 B.n833 B.n832 46.5903
R1992 B.n832 B.n65 46.5903
R1993 B.n826 B.n65 46.5903
R1994 B.n826 B.n825 46.5903
R1995 B.n825 B.n824 46.5903
R1996 B.n818 B.n75 46.5903
R1997 B.n818 B.n817 46.5903
R1998 B.n817 B.n816 46.5903
R1999 B.n816 B.n79 46.5903
R2000 B.n810 B.n79 46.5903
R2001 B.n810 B.n809 46.5903
R2002 B.n626 B.t9 43.8498
R2003 B.n75 B.t13 43.8498
R2004 B.t7 B.n337 39.7389
R2005 B.n736 B.t4 39.7389
R2006 B.n890 B.t1 39.7389
R2007 B.t2 B.n37 39.7389
R2008 B.n605 B.n386 31.6883
R2009 B.n611 B.n610 31.6883
R2010 B.n805 B.n804 31.6883
R2011 B.n135 B.n81 31.6883
R2012 B.n663 B.t0 30.1469
R2013 B.n329 B.t3 30.1469
R2014 B.t5 B.n873 30.1469
R2015 B.n842 B.t6 30.1469
R2016 B B.n902 18.0485
R2017 B.t0 B.n353 16.444
R2018 B.n711 B.t3 16.444
R2019 B.n874 B.t5 16.444
R2020 B.t6 B.n51 16.444
R2021 B.n616 B.n386 10.6151
R2022 B.n617 B.n616 10.6151
R2023 B.n618 B.n617 10.6151
R2024 B.n618 B.n378 10.6151
R2025 B.n629 B.n378 10.6151
R2026 B.n630 B.n629 10.6151
R2027 B.n631 B.n630 10.6151
R2028 B.n631 B.n371 10.6151
R2029 B.n641 B.n371 10.6151
R2030 B.n642 B.n641 10.6151
R2031 B.n643 B.n642 10.6151
R2032 B.n643 B.n363 10.6151
R2033 B.n653 B.n363 10.6151
R2034 B.n654 B.n653 10.6151
R2035 B.n655 B.n654 10.6151
R2036 B.n655 B.n355 10.6151
R2037 B.n665 B.n355 10.6151
R2038 B.n666 B.n665 10.6151
R2039 B.n667 B.n666 10.6151
R2040 B.n667 B.n347 10.6151
R2041 B.n677 B.n347 10.6151
R2042 B.n678 B.n677 10.6151
R2043 B.n679 B.n678 10.6151
R2044 B.n679 B.n339 10.6151
R2045 B.n689 B.n339 10.6151
R2046 B.n690 B.n689 10.6151
R2047 B.n691 B.n690 10.6151
R2048 B.n691 B.n331 10.6151
R2049 B.n701 B.n331 10.6151
R2050 B.n702 B.n701 10.6151
R2051 B.n703 B.n702 10.6151
R2052 B.n703 B.n323 10.6151
R2053 B.n713 B.n323 10.6151
R2054 B.n714 B.n713 10.6151
R2055 B.n715 B.n714 10.6151
R2056 B.n715 B.n315 10.6151
R2057 B.n725 B.n315 10.6151
R2058 B.n726 B.n725 10.6151
R2059 B.n727 B.n726 10.6151
R2060 B.n727 B.n307 10.6151
R2061 B.n738 B.n307 10.6151
R2062 B.n739 B.n738 10.6151
R2063 B.n740 B.n739 10.6151
R2064 B.n740 B.n0 10.6151
R2065 B.n605 B.n604 10.6151
R2066 B.n604 B.n603 10.6151
R2067 B.n603 B.n602 10.6151
R2068 B.n602 B.n600 10.6151
R2069 B.n600 B.n597 10.6151
R2070 B.n597 B.n596 10.6151
R2071 B.n596 B.n593 10.6151
R2072 B.n593 B.n592 10.6151
R2073 B.n592 B.n589 10.6151
R2074 B.n589 B.n588 10.6151
R2075 B.n588 B.n585 10.6151
R2076 B.n585 B.n584 10.6151
R2077 B.n584 B.n581 10.6151
R2078 B.n581 B.n580 10.6151
R2079 B.n580 B.n577 10.6151
R2080 B.n577 B.n576 10.6151
R2081 B.n576 B.n573 10.6151
R2082 B.n573 B.n572 10.6151
R2083 B.n572 B.n569 10.6151
R2084 B.n569 B.n568 10.6151
R2085 B.n568 B.n565 10.6151
R2086 B.n565 B.n564 10.6151
R2087 B.n564 B.n561 10.6151
R2088 B.n561 B.n560 10.6151
R2089 B.n560 B.n557 10.6151
R2090 B.n557 B.n556 10.6151
R2091 B.n556 B.n553 10.6151
R2092 B.n553 B.n552 10.6151
R2093 B.n552 B.n549 10.6151
R2094 B.n549 B.n548 10.6151
R2095 B.n548 B.n545 10.6151
R2096 B.n545 B.n544 10.6151
R2097 B.n544 B.n541 10.6151
R2098 B.n541 B.n540 10.6151
R2099 B.n540 B.n537 10.6151
R2100 B.n537 B.n536 10.6151
R2101 B.n536 B.n533 10.6151
R2102 B.n531 B.n528 10.6151
R2103 B.n528 B.n527 10.6151
R2104 B.n527 B.n524 10.6151
R2105 B.n524 B.n523 10.6151
R2106 B.n523 B.n520 10.6151
R2107 B.n520 B.n519 10.6151
R2108 B.n519 B.n516 10.6151
R2109 B.n516 B.n515 10.6151
R2110 B.n515 B.n512 10.6151
R2111 B.n510 B.n507 10.6151
R2112 B.n507 B.n506 10.6151
R2113 B.n506 B.n503 10.6151
R2114 B.n503 B.n502 10.6151
R2115 B.n502 B.n499 10.6151
R2116 B.n499 B.n498 10.6151
R2117 B.n498 B.n495 10.6151
R2118 B.n495 B.n494 10.6151
R2119 B.n494 B.n491 10.6151
R2120 B.n491 B.n490 10.6151
R2121 B.n490 B.n487 10.6151
R2122 B.n487 B.n486 10.6151
R2123 B.n486 B.n483 10.6151
R2124 B.n483 B.n482 10.6151
R2125 B.n482 B.n479 10.6151
R2126 B.n479 B.n478 10.6151
R2127 B.n478 B.n475 10.6151
R2128 B.n475 B.n474 10.6151
R2129 B.n474 B.n471 10.6151
R2130 B.n471 B.n470 10.6151
R2131 B.n470 B.n467 10.6151
R2132 B.n467 B.n466 10.6151
R2133 B.n466 B.n463 10.6151
R2134 B.n463 B.n462 10.6151
R2135 B.n462 B.n459 10.6151
R2136 B.n459 B.n458 10.6151
R2137 B.n458 B.n455 10.6151
R2138 B.n455 B.n454 10.6151
R2139 B.n454 B.n451 10.6151
R2140 B.n451 B.n450 10.6151
R2141 B.n450 B.n447 10.6151
R2142 B.n447 B.n446 10.6151
R2143 B.n446 B.n443 10.6151
R2144 B.n443 B.n442 10.6151
R2145 B.n442 B.n439 10.6151
R2146 B.n439 B.n390 10.6151
R2147 B.n610 B.n390 10.6151
R2148 B.n612 B.n611 10.6151
R2149 B.n612 B.n382 10.6151
R2150 B.n622 B.n382 10.6151
R2151 B.n623 B.n622 10.6151
R2152 B.n624 B.n623 10.6151
R2153 B.n624 B.n375 10.6151
R2154 B.n635 B.n375 10.6151
R2155 B.n636 B.n635 10.6151
R2156 B.n637 B.n636 10.6151
R2157 B.n637 B.n367 10.6151
R2158 B.n647 B.n367 10.6151
R2159 B.n648 B.n647 10.6151
R2160 B.n649 B.n648 10.6151
R2161 B.n649 B.n359 10.6151
R2162 B.n659 B.n359 10.6151
R2163 B.n660 B.n659 10.6151
R2164 B.n661 B.n660 10.6151
R2165 B.n661 B.n351 10.6151
R2166 B.n671 B.n351 10.6151
R2167 B.n672 B.n671 10.6151
R2168 B.n673 B.n672 10.6151
R2169 B.n673 B.n343 10.6151
R2170 B.n683 B.n343 10.6151
R2171 B.n684 B.n683 10.6151
R2172 B.n685 B.n684 10.6151
R2173 B.n685 B.n335 10.6151
R2174 B.n695 B.n335 10.6151
R2175 B.n696 B.n695 10.6151
R2176 B.n697 B.n696 10.6151
R2177 B.n697 B.n326 10.6151
R2178 B.n707 B.n326 10.6151
R2179 B.n708 B.n707 10.6151
R2180 B.n709 B.n708 10.6151
R2181 B.n709 B.n319 10.6151
R2182 B.n719 B.n319 10.6151
R2183 B.n720 B.n719 10.6151
R2184 B.n721 B.n720 10.6151
R2185 B.n721 B.n310 10.6151
R2186 B.n731 B.n310 10.6151
R2187 B.n732 B.n731 10.6151
R2188 B.n734 B.n732 10.6151
R2189 B.n734 B.n733 10.6151
R2190 B.n733 B.n303 10.6151
R2191 B.n745 B.n303 10.6151
R2192 B.n746 B.n745 10.6151
R2193 B.n747 B.n746 10.6151
R2194 B.n748 B.n747 10.6151
R2195 B.n749 B.n748 10.6151
R2196 B.n752 B.n749 10.6151
R2197 B.n753 B.n752 10.6151
R2198 B.n754 B.n753 10.6151
R2199 B.n755 B.n754 10.6151
R2200 B.n757 B.n755 10.6151
R2201 B.n758 B.n757 10.6151
R2202 B.n759 B.n758 10.6151
R2203 B.n760 B.n759 10.6151
R2204 B.n762 B.n760 10.6151
R2205 B.n763 B.n762 10.6151
R2206 B.n764 B.n763 10.6151
R2207 B.n765 B.n764 10.6151
R2208 B.n767 B.n765 10.6151
R2209 B.n768 B.n767 10.6151
R2210 B.n769 B.n768 10.6151
R2211 B.n770 B.n769 10.6151
R2212 B.n772 B.n770 10.6151
R2213 B.n773 B.n772 10.6151
R2214 B.n774 B.n773 10.6151
R2215 B.n775 B.n774 10.6151
R2216 B.n777 B.n775 10.6151
R2217 B.n778 B.n777 10.6151
R2218 B.n779 B.n778 10.6151
R2219 B.n780 B.n779 10.6151
R2220 B.n782 B.n780 10.6151
R2221 B.n783 B.n782 10.6151
R2222 B.n784 B.n783 10.6151
R2223 B.n785 B.n784 10.6151
R2224 B.n787 B.n785 10.6151
R2225 B.n788 B.n787 10.6151
R2226 B.n789 B.n788 10.6151
R2227 B.n790 B.n789 10.6151
R2228 B.n792 B.n790 10.6151
R2229 B.n793 B.n792 10.6151
R2230 B.n794 B.n793 10.6151
R2231 B.n795 B.n794 10.6151
R2232 B.n797 B.n795 10.6151
R2233 B.n798 B.n797 10.6151
R2234 B.n799 B.n798 10.6151
R2235 B.n800 B.n799 10.6151
R2236 B.n802 B.n800 10.6151
R2237 B.n803 B.n802 10.6151
R2238 B.n804 B.n803 10.6151
R2239 B.n894 B.n1 10.6151
R2240 B.n894 B.n893 10.6151
R2241 B.n893 B.n892 10.6151
R2242 B.n892 B.n10 10.6151
R2243 B.n886 B.n10 10.6151
R2244 B.n886 B.n885 10.6151
R2245 B.n885 B.n884 10.6151
R2246 B.n884 B.n18 10.6151
R2247 B.n878 B.n18 10.6151
R2248 B.n878 B.n877 10.6151
R2249 B.n877 B.n876 10.6151
R2250 B.n876 B.n25 10.6151
R2251 B.n870 B.n25 10.6151
R2252 B.n870 B.n869 10.6151
R2253 B.n869 B.n868 10.6151
R2254 B.n868 B.n32 10.6151
R2255 B.n862 B.n32 10.6151
R2256 B.n862 B.n861 10.6151
R2257 B.n861 B.n860 10.6151
R2258 B.n860 B.n39 10.6151
R2259 B.n854 B.n39 10.6151
R2260 B.n854 B.n853 10.6151
R2261 B.n853 B.n852 10.6151
R2262 B.n852 B.n46 10.6151
R2263 B.n846 B.n46 10.6151
R2264 B.n846 B.n845 10.6151
R2265 B.n845 B.n844 10.6151
R2266 B.n844 B.n53 10.6151
R2267 B.n838 B.n53 10.6151
R2268 B.n838 B.n837 10.6151
R2269 B.n837 B.n836 10.6151
R2270 B.n836 B.n60 10.6151
R2271 B.n830 B.n60 10.6151
R2272 B.n830 B.n829 10.6151
R2273 B.n829 B.n828 10.6151
R2274 B.n828 B.n67 10.6151
R2275 B.n822 B.n67 10.6151
R2276 B.n822 B.n821 10.6151
R2277 B.n821 B.n820 10.6151
R2278 B.n820 B.n73 10.6151
R2279 B.n814 B.n73 10.6151
R2280 B.n814 B.n813 10.6151
R2281 B.n813 B.n812 10.6151
R2282 B.n812 B.n81 10.6151
R2283 B.n136 B.n135 10.6151
R2284 B.n139 B.n136 10.6151
R2285 B.n140 B.n139 10.6151
R2286 B.n143 B.n140 10.6151
R2287 B.n144 B.n143 10.6151
R2288 B.n147 B.n144 10.6151
R2289 B.n148 B.n147 10.6151
R2290 B.n151 B.n148 10.6151
R2291 B.n152 B.n151 10.6151
R2292 B.n155 B.n152 10.6151
R2293 B.n156 B.n155 10.6151
R2294 B.n159 B.n156 10.6151
R2295 B.n160 B.n159 10.6151
R2296 B.n163 B.n160 10.6151
R2297 B.n164 B.n163 10.6151
R2298 B.n167 B.n164 10.6151
R2299 B.n168 B.n167 10.6151
R2300 B.n171 B.n168 10.6151
R2301 B.n172 B.n171 10.6151
R2302 B.n175 B.n172 10.6151
R2303 B.n176 B.n175 10.6151
R2304 B.n179 B.n176 10.6151
R2305 B.n180 B.n179 10.6151
R2306 B.n183 B.n180 10.6151
R2307 B.n184 B.n183 10.6151
R2308 B.n187 B.n184 10.6151
R2309 B.n188 B.n187 10.6151
R2310 B.n191 B.n188 10.6151
R2311 B.n192 B.n191 10.6151
R2312 B.n195 B.n192 10.6151
R2313 B.n196 B.n195 10.6151
R2314 B.n199 B.n196 10.6151
R2315 B.n200 B.n199 10.6151
R2316 B.n203 B.n200 10.6151
R2317 B.n204 B.n203 10.6151
R2318 B.n207 B.n204 10.6151
R2319 B.n208 B.n207 10.6151
R2320 B.n212 B.n211 10.6151
R2321 B.n215 B.n212 10.6151
R2322 B.n216 B.n215 10.6151
R2323 B.n219 B.n216 10.6151
R2324 B.n220 B.n219 10.6151
R2325 B.n223 B.n220 10.6151
R2326 B.n224 B.n223 10.6151
R2327 B.n227 B.n224 10.6151
R2328 B.n228 B.n227 10.6151
R2329 B.n232 B.n231 10.6151
R2330 B.n235 B.n232 10.6151
R2331 B.n236 B.n235 10.6151
R2332 B.n239 B.n236 10.6151
R2333 B.n240 B.n239 10.6151
R2334 B.n243 B.n240 10.6151
R2335 B.n244 B.n243 10.6151
R2336 B.n247 B.n244 10.6151
R2337 B.n248 B.n247 10.6151
R2338 B.n251 B.n248 10.6151
R2339 B.n252 B.n251 10.6151
R2340 B.n255 B.n252 10.6151
R2341 B.n256 B.n255 10.6151
R2342 B.n259 B.n256 10.6151
R2343 B.n260 B.n259 10.6151
R2344 B.n263 B.n260 10.6151
R2345 B.n264 B.n263 10.6151
R2346 B.n267 B.n264 10.6151
R2347 B.n268 B.n267 10.6151
R2348 B.n271 B.n268 10.6151
R2349 B.n272 B.n271 10.6151
R2350 B.n275 B.n272 10.6151
R2351 B.n276 B.n275 10.6151
R2352 B.n279 B.n276 10.6151
R2353 B.n280 B.n279 10.6151
R2354 B.n283 B.n280 10.6151
R2355 B.n284 B.n283 10.6151
R2356 B.n287 B.n284 10.6151
R2357 B.n288 B.n287 10.6151
R2358 B.n291 B.n288 10.6151
R2359 B.n292 B.n291 10.6151
R2360 B.n295 B.n292 10.6151
R2361 B.n296 B.n295 10.6151
R2362 B.n299 B.n296 10.6151
R2363 B.n301 B.n299 10.6151
R2364 B.n302 B.n301 10.6151
R2365 B.n805 B.n302 10.6151
R2366 B.n533 B.n532 9.36635
R2367 B.n511 B.n510 9.36635
R2368 B.n208 B.n133 9.36635
R2369 B.n231 B.n130 9.36635
R2370 B.n902 B.n0 8.11757
R2371 B.n902 B.n1 8.11757
R2372 B.n687 B.t7 6.85195
R2373 B.n313 B.t4 6.85195
R2374 B.t1 B.n889 6.85195
R2375 B.n858 B.t2 6.85195
R2376 B.n633 B.t9 2.74108
R2377 B.n824 B.t13 2.74108
R2378 B.n532 B.n531 1.24928
R2379 B.n512 B.n511 1.24928
R2380 B.n211 B.n133 1.24928
R2381 B.n228 B.n130 1.24928
R2382 VN.n47 VN.n25 161.3
R2383 VN.n46 VN.n45 161.3
R2384 VN.n44 VN.n26 161.3
R2385 VN.n43 VN.n42 161.3
R2386 VN.n41 VN.n27 161.3
R2387 VN.n39 VN.n38 161.3
R2388 VN.n37 VN.n28 161.3
R2389 VN.n36 VN.n35 161.3
R2390 VN.n34 VN.n29 161.3
R2391 VN.n33 VN.n32 161.3
R2392 VN.n22 VN.n0 161.3
R2393 VN.n21 VN.n20 161.3
R2394 VN.n19 VN.n1 161.3
R2395 VN.n18 VN.n17 161.3
R2396 VN.n16 VN.n2 161.3
R2397 VN.n14 VN.n13 161.3
R2398 VN.n12 VN.n3 161.3
R2399 VN.n11 VN.n10 161.3
R2400 VN.n9 VN.n4 161.3
R2401 VN.n8 VN.n7 161.3
R2402 VN.n6 VN.t1 150.167
R2403 VN.n31 VN.t6 150.167
R2404 VN.n5 VN.t4 117.026
R2405 VN.n15 VN.t0 117.026
R2406 VN.n23 VN.t3 117.026
R2407 VN.n30 VN.t7 117.026
R2408 VN.n40 VN.t2 117.026
R2409 VN.n48 VN.t5 117.026
R2410 VN.n24 VN.n23 94.9235
R2411 VN.n49 VN.n48 94.9235
R2412 VN.n6 VN.n5 58.066
R2413 VN.n31 VN.n30 58.066
R2414 VN VN.n49 48.4906
R2415 VN.n21 VN.n1 45.4209
R2416 VN.n46 VN.n26 45.4209
R2417 VN.n10 VN.n9 40.577
R2418 VN.n10 VN.n3 40.577
R2419 VN.n35 VN.n34 40.577
R2420 VN.n35 VN.n28 40.577
R2421 VN.n17 VN.n1 35.7332
R2422 VN.n42 VN.n26 35.7332
R2423 VN.n9 VN.n8 24.5923
R2424 VN.n14 VN.n3 24.5923
R2425 VN.n17 VN.n16 24.5923
R2426 VN.n22 VN.n21 24.5923
R2427 VN.n34 VN.n33 24.5923
R2428 VN.n42 VN.n41 24.5923
R2429 VN.n39 VN.n28 24.5923
R2430 VN.n47 VN.n46 24.5923
R2431 VN.n23 VN.n22 15.9852
R2432 VN.n48 VN.n47 15.9852
R2433 VN.n8 VN.n5 13.526
R2434 VN.n15 VN.n14 13.526
R2435 VN.n33 VN.n30 13.526
R2436 VN.n40 VN.n39 13.526
R2437 VN.n16 VN.n15 11.0668
R2438 VN.n41 VN.n40 11.0668
R2439 VN.n32 VN.n31 9.34229
R2440 VN.n7 VN.n6 9.34229
R2441 VN.n49 VN.n25 0.278335
R2442 VN.n24 VN.n0 0.278335
R2443 VN.n45 VN.n25 0.189894
R2444 VN.n45 VN.n44 0.189894
R2445 VN.n44 VN.n43 0.189894
R2446 VN.n43 VN.n27 0.189894
R2447 VN.n38 VN.n27 0.189894
R2448 VN.n38 VN.n37 0.189894
R2449 VN.n37 VN.n36 0.189894
R2450 VN.n36 VN.n29 0.189894
R2451 VN.n32 VN.n29 0.189894
R2452 VN.n7 VN.n4 0.189894
R2453 VN.n11 VN.n4 0.189894
R2454 VN.n12 VN.n11 0.189894
R2455 VN.n13 VN.n12 0.189894
R2456 VN.n13 VN.n2 0.189894
R2457 VN.n18 VN.n2 0.189894
R2458 VN.n19 VN.n18 0.189894
R2459 VN.n20 VN.n19 0.189894
R2460 VN.n20 VN.n0 0.189894
R2461 VN VN.n24 0.153485
R2462 VDD2.n2 VDD2.n1 65.3233
R2463 VDD2.n2 VDD2.n0 65.3233
R2464 VDD2 VDD2.n5 65.3205
R2465 VDD2.n4 VDD2.n3 64.2797
R2466 VDD2.n4 VDD2.n2 42.9006
R2467 VDD2.n5 VDD2.t0 1.83723
R2468 VDD2.n5 VDD2.t1 1.83723
R2469 VDD2.n3 VDD2.t2 1.83723
R2470 VDD2.n3 VDD2.t5 1.83723
R2471 VDD2.n1 VDD2.t7 1.83723
R2472 VDD2.n1 VDD2.t4 1.83723
R2473 VDD2.n0 VDD2.t6 1.83723
R2474 VDD2.n0 VDD2.t3 1.83723
R2475 VDD2 VDD2.n4 1.15783
C0 VDD1 VDD2 1.57731f
C1 VN VTAIL 7.9272f
C2 VP VTAIL 7.94131f
C3 VP VN 6.96742f
C4 VDD1 VTAIL 7.60962f
C5 VDD2 VTAIL 7.66148f
C6 VDD1 VN 0.151043f
C7 VDD1 VP 7.93052f
C8 VDD2 VN 7.60353f
C9 VDD2 VP 0.479237f
C10 VDD2 B 4.88231f
C11 VDD1 B 5.276041f
C12 VTAIL B 9.487853f
C13 VN B 13.95968f
C14 VP B 12.51918f
C15 VDD2.t6 B 0.208652f
C16 VDD2.t3 B 0.208652f
C17 VDD2.n0 B 1.85577f
C18 VDD2.t7 B 0.208652f
C19 VDD2.t4 B 0.208652f
C20 VDD2.n1 B 1.85577f
C21 VDD2.n2 B 2.91726f
C22 VDD2.t2 B 0.208652f
C23 VDD2.t5 B 0.208652f
C24 VDD2.n3 B 1.84833f
C25 VDD2.n4 B 2.66695f
C26 VDD2.t0 B 0.208652f
C27 VDD2.t1 B 0.208652f
C28 VDD2.n5 B 1.85574f
C29 VN.n0 B 0.032668f
C30 VN.t3 B 1.61054f
C31 VN.n1 B 0.020815f
C32 VN.n2 B 0.02478f
C33 VN.t0 B 1.61054f
C34 VN.n3 B 0.04899f
C35 VN.n4 B 0.02478f
C36 VN.t4 B 1.61054f
C37 VN.n5 B 0.641582f
C38 VN.t1 B 1.76752f
C39 VN.n6 B 0.630602f
C40 VN.n7 B 0.211471f
C41 VN.n8 B 0.035744f
C42 VN.n9 B 0.04899f
C43 VN.n10 B 0.020014f
C44 VN.n11 B 0.02478f
C45 VN.n12 B 0.02478f
C46 VN.n13 B 0.02478f
C47 VN.n14 B 0.035744f
C48 VN.n15 B 0.57666f
C49 VN.n16 B 0.033475f
C50 VN.n17 B 0.049771f
C51 VN.n18 B 0.02478f
C52 VN.n19 B 0.02478f
C53 VN.n20 B 0.02478f
C54 VN.n21 B 0.047408f
C55 VN.n22 B 0.038012f
C56 VN.n23 B 0.65454f
C57 VN.n24 B 0.033851f
C58 VN.n25 B 0.032668f
C59 VN.t5 B 1.61054f
C60 VN.n26 B 0.020815f
C61 VN.n27 B 0.02478f
C62 VN.t2 B 1.61054f
C63 VN.n28 B 0.04899f
C64 VN.n29 B 0.02478f
C65 VN.t7 B 1.61054f
C66 VN.n30 B 0.641582f
C67 VN.t6 B 1.76752f
C68 VN.n31 B 0.630602f
C69 VN.n32 B 0.211471f
C70 VN.n33 B 0.035744f
C71 VN.n34 B 0.04899f
C72 VN.n35 B 0.020014f
C73 VN.n36 B 0.02478f
C74 VN.n37 B 0.02478f
C75 VN.n38 B 0.02478f
C76 VN.n39 B 0.035744f
C77 VN.n40 B 0.57666f
C78 VN.n41 B 0.033475f
C79 VN.n42 B 0.049771f
C80 VN.n43 B 0.02478f
C81 VN.n44 B 0.02478f
C82 VN.n45 B 0.02478f
C83 VN.n46 B 0.047408f
C84 VN.n47 B 0.038012f
C85 VN.n48 B 0.65454f
C86 VN.n49 B 1.31285f
C87 VTAIL.t5 B 0.169529f
C88 VTAIL.t2 B 0.169529f
C89 VTAIL.n0 B 1.44633f
C90 VTAIL.n1 B 0.335049f
C91 VTAIL.n2 B 0.028241f
C92 VTAIL.n3 B 0.019901f
C93 VTAIL.n4 B 0.010694f
C94 VTAIL.n5 B 0.025276f
C95 VTAIL.n6 B 0.011323f
C96 VTAIL.n7 B 0.019901f
C97 VTAIL.n8 B 0.010694f
C98 VTAIL.n9 B 0.025276f
C99 VTAIL.n10 B 0.011323f
C100 VTAIL.n11 B 0.019901f
C101 VTAIL.n12 B 0.010694f
C102 VTAIL.n13 B 0.025276f
C103 VTAIL.n14 B 0.011323f
C104 VTAIL.n15 B 0.019901f
C105 VTAIL.n16 B 0.010694f
C106 VTAIL.n17 B 0.025276f
C107 VTAIL.n18 B 0.011323f
C108 VTAIL.n19 B 0.134163f
C109 VTAIL.t1 B 0.04256f
C110 VTAIL.n20 B 0.018957f
C111 VTAIL.n21 B 0.017868f
C112 VTAIL.n22 B 0.010694f
C113 VTAIL.n23 B 0.89597f
C114 VTAIL.n24 B 0.019901f
C115 VTAIL.n25 B 0.010694f
C116 VTAIL.n26 B 0.011323f
C117 VTAIL.n27 B 0.025276f
C118 VTAIL.n28 B 0.025276f
C119 VTAIL.n29 B 0.011323f
C120 VTAIL.n30 B 0.010694f
C121 VTAIL.n31 B 0.019901f
C122 VTAIL.n32 B 0.019901f
C123 VTAIL.n33 B 0.010694f
C124 VTAIL.n34 B 0.011323f
C125 VTAIL.n35 B 0.025276f
C126 VTAIL.n36 B 0.025276f
C127 VTAIL.n37 B 0.025276f
C128 VTAIL.n38 B 0.011323f
C129 VTAIL.n39 B 0.010694f
C130 VTAIL.n40 B 0.019901f
C131 VTAIL.n41 B 0.019901f
C132 VTAIL.n42 B 0.010694f
C133 VTAIL.n43 B 0.011008f
C134 VTAIL.n44 B 0.011008f
C135 VTAIL.n45 B 0.025276f
C136 VTAIL.n46 B 0.025276f
C137 VTAIL.n47 B 0.011323f
C138 VTAIL.n48 B 0.010694f
C139 VTAIL.n49 B 0.019901f
C140 VTAIL.n50 B 0.019901f
C141 VTAIL.n51 B 0.010694f
C142 VTAIL.n52 B 0.011323f
C143 VTAIL.n53 B 0.025276f
C144 VTAIL.n54 B 0.055194f
C145 VTAIL.n55 B 0.011323f
C146 VTAIL.n56 B 0.010694f
C147 VTAIL.n57 B 0.048718f
C148 VTAIL.n58 B 0.031013f
C149 VTAIL.n59 B 0.189625f
C150 VTAIL.n60 B 0.028241f
C151 VTAIL.n61 B 0.019901f
C152 VTAIL.n62 B 0.010694f
C153 VTAIL.n63 B 0.025276f
C154 VTAIL.n64 B 0.011323f
C155 VTAIL.n65 B 0.019901f
C156 VTAIL.n66 B 0.010694f
C157 VTAIL.n67 B 0.025276f
C158 VTAIL.n68 B 0.011323f
C159 VTAIL.n69 B 0.019901f
C160 VTAIL.n70 B 0.010694f
C161 VTAIL.n71 B 0.025276f
C162 VTAIL.n72 B 0.011323f
C163 VTAIL.n73 B 0.019901f
C164 VTAIL.n74 B 0.010694f
C165 VTAIL.n75 B 0.025276f
C166 VTAIL.n76 B 0.011323f
C167 VTAIL.n77 B 0.134163f
C168 VTAIL.t12 B 0.04256f
C169 VTAIL.n78 B 0.018957f
C170 VTAIL.n79 B 0.017868f
C171 VTAIL.n80 B 0.010694f
C172 VTAIL.n81 B 0.89597f
C173 VTAIL.n82 B 0.019901f
C174 VTAIL.n83 B 0.010694f
C175 VTAIL.n84 B 0.011323f
C176 VTAIL.n85 B 0.025276f
C177 VTAIL.n86 B 0.025276f
C178 VTAIL.n87 B 0.011323f
C179 VTAIL.n88 B 0.010694f
C180 VTAIL.n89 B 0.019901f
C181 VTAIL.n90 B 0.019901f
C182 VTAIL.n91 B 0.010694f
C183 VTAIL.n92 B 0.011323f
C184 VTAIL.n93 B 0.025276f
C185 VTAIL.n94 B 0.025276f
C186 VTAIL.n95 B 0.025276f
C187 VTAIL.n96 B 0.011323f
C188 VTAIL.n97 B 0.010694f
C189 VTAIL.n98 B 0.019901f
C190 VTAIL.n99 B 0.019901f
C191 VTAIL.n100 B 0.010694f
C192 VTAIL.n101 B 0.011008f
C193 VTAIL.n102 B 0.011008f
C194 VTAIL.n103 B 0.025276f
C195 VTAIL.n104 B 0.025276f
C196 VTAIL.n105 B 0.011323f
C197 VTAIL.n106 B 0.010694f
C198 VTAIL.n107 B 0.019901f
C199 VTAIL.n108 B 0.019901f
C200 VTAIL.n109 B 0.010694f
C201 VTAIL.n110 B 0.011323f
C202 VTAIL.n111 B 0.025276f
C203 VTAIL.n112 B 0.055194f
C204 VTAIL.n113 B 0.011323f
C205 VTAIL.n114 B 0.010694f
C206 VTAIL.n115 B 0.048718f
C207 VTAIL.n116 B 0.031013f
C208 VTAIL.n117 B 0.189625f
C209 VTAIL.t8 B 0.169529f
C210 VTAIL.t11 B 0.169529f
C211 VTAIL.n118 B 1.44633f
C212 VTAIL.n119 B 0.472282f
C213 VTAIL.n120 B 0.028241f
C214 VTAIL.n121 B 0.019901f
C215 VTAIL.n122 B 0.010694f
C216 VTAIL.n123 B 0.025276f
C217 VTAIL.n124 B 0.011323f
C218 VTAIL.n125 B 0.019901f
C219 VTAIL.n126 B 0.010694f
C220 VTAIL.n127 B 0.025276f
C221 VTAIL.n128 B 0.011323f
C222 VTAIL.n129 B 0.019901f
C223 VTAIL.n130 B 0.010694f
C224 VTAIL.n131 B 0.025276f
C225 VTAIL.n132 B 0.011323f
C226 VTAIL.n133 B 0.019901f
C227 VTAIL.n134 B 0.010694f
C228 VTAIL.n135 B 0.025276f
C229 VTAIL.n136 B 0.011323f
C230 VTAIL.n137 B 0.134163f
C231 VTAIL.t14 B 0.04256f
C232 VTAIL.n138 B 0.018957f
C233 VTAIL.n139 B 0.017868f
C234 VTAIL.n140 B 0.010694f
C235 VTAIL.n141 B 0.89597f
C236 VTAIL.n142 B 0.019901f
C237 VTAIL.n143 B 0.010694f
C238 VTAIL.n144 B 0.011323f
C239 VTAIL.n145 B 0.025276f
C240 VTAIL.n146 B 0.025276f
C241 VTAIL.n147 B 0.011323f
C242 VTAIL.n148 B 0.010694f
C243 VTAIL.n149 B 0.019901f
C244 VTAIL.n150 B 0.019901f
C245 VTAIL.n151 B 0.010694f
C246 VTAIL.n152 B 0.011323f
C247 VTAIL.n153 B 0.025276f
C248 VTAIL.n154 B 0.025276f
C249 VTAIL.n155 B 0.025276f
C250 VTAIL.n156 B 0.011323f
C251 VTAIL.n157 B 0.010694f
C252 VTAIL.n158 B 0.019901f
C253 VTAIL.n159 B 0.019901f
C254 VTAIL.n160 B 0.010694f
C255 VTAIL.n161 B 0.011008f
C256 VTAIL.n162 B 0.011008f
C257 VTAIL.n163 B 0.025276f
C258 VTAIL.n164 B 0.025276f
C259 VTAIL.n165 B 0.011323f
C260 VTAIL.n166 B 0.010694f
C261 VTAIL.n167 B 0.019901f
C262 VTAIL.n168 B 0.019901f
C263 VTAIL.n169 B 0.010694f
C264 VTAIL.n170 B 0.011323f
C265 VTAIL.n171 B 0.025276f
C266 VTAIL.n172 B 0.055194f
C267 VTAIL.n173 B 0.011323f
C268 VTAIL.n174 B 0.010694f
C269 VTAIL.n175 B 0.048718f
C270 VTAIL.n176 B 0.031013f
C271 VTAIL.n177 B 1.16671f
C272 VTAIL.n178 B 0.028241f
C273 VTAIL.n179 B 0.019901f
C274 VTAIL.n180 B 0.010694f
C275 VTAIL.n181 B 0.025276f
C276 VTAIL.n182 B 0.011323f
C277 VTAIL.n183 B 0.019901f
C278 VTAIL.n184 B 0.010694f
C279 VTAIL.n185 B 0.025276f
C280 VTAIL.n186 B 0.011323f
C281 VTAIL.n187 B 0.019901f
C282 VTAIL.n188 B 0.010694f
C283 VTAIL.n189 B 0.025276f
C284 VTAIL.n190 B 0.025276f
C285 VTAIL.n191 B 0.011323f
C286 VTAIL.n192 B 0.019901f
C287 VTAIL.n193 B 0.010694f
C288 VTAIL.n194 B 0.025276f
C289 VTAIL.n195 B 0.011323f
C290 VTAIL.n196 B 0.134163f
C291 VTAIL.t0 B 0.04256f
C292 VTAIL.n197 B 0.018957f
C293 VTAIL.n198 B 0.017868f
C294 VTAIL.n199 B 0.010694f
C295 VTAIL.n200 B 0.89597f
C296 VTAIL.n201 B 0.019901f
C297 VTAIL.n202 B 0.010694f
C298 VTAIL.n203 B 0.011323f
C299 VTAIL.n204 B 0.025276f
C300 VTAIL.n205 B 0.025276f
C301 VTAIL.n206 B 0.011323f
C302 VTAIL.n207 B 0.010694f
C303 VTAIL.n208 B 0.019901f
C304 VTAIL.n209 B 0.019901f
C305 VTAIL.n210 B 0.010694f
C306 VTAIL.n211 B 0.011323f
C307 VTAIL.n212 B 0.025276f
C308 VTAIL.n213 B 0.025276f
C309 VTAIL.n214 B 0.011323f
C310 VTAIL.n215 B 0.010694f
C311 VTAIL.n216 B 0.019901f
C312 VTAIL.n217 B 0.019901f
C313 VTAIL.n218 B 0.010694f
C314 VTAIL.n219 B 0.011008f
C315 VTAIL.n220 B 0.011008f
C316 VTAIL.n221 B 0.025276f
C317 VTAIL.n222 B 0.025276f
C318 VTAIL.n223 B 0.011323f
C319 VTAIL.n224 B 0.010694f
C320 VTAIL.n225 B 0.019901f
C321 VTAIL.n226 B 0.019901f
C322 VTAIL.n227 B 0.010694f
C323 VTAIL.n228 B 0.011323f
C324 VTAIL.n229 B 0.025276f
C325 VTAIL.n230 B 0.055194f
C326 VTAIL.n231 B 0.011323f
C327 VTAIL.n232 B 0.010694f
C328 VTAIL.n233 B 0.048718f
C329 VTAIL.n234 B 0.031013f
C330 VTAIL.n235 B 1.16671f
C331 VTAIL.t7 B 0.169529f
C332 VTAIL.t3 B 0.169529f
C333 VTAIL.n236 B 1.44634f
C334 VTAIL.n237 B 0.472274f
C335 VTAIL.n238 B 0.028241f
C336 VTAIL.n239 B 0.019901f
C337 VTAIL.n240 B 0.010694f
C338 VTAIL.n241 B 0.025276f
C339 VTAIL.n242 B 0.011323f
C340 VTAIL.n243 B 0.019901f
C341 VTAIL.n244 B 0.010694f
C342 VTAIL.n245 B 0.025276f
C343 VTAIL.n246 B 0.011323f
C344 VTAIL.n247 B 0.019901f
C345 VTAIL.n248 B 0.010694f
C346 VTAIL.n249 B 0.025276f
C347 VTAIL.n250 B 0.025276f
C348 VTAIL.n251 B 0.011323f
C349 VTAIL.n252 B 0.019901f
C350 VTAIL.n253 B 0.010694f
C351 VTAIL.n254 B 0.025276f
C352 VTAIL.n255 B 0.011323f
C353 VTAIL.n256 B 0.134163f
C354 VTAIL.t4 B 0.04256f
C355 VTAIL.n257 B 0.018957f
C356 VTAIL.n258 B 0.017868f
C357 VTAIL.n259 B 0.010694f
C358 VTAIL.n260 B 0.89597f
C359 VTAIL.n261 B 0.019901f
C360 VTAIL.n262 B 0.010694f
C361 VTAIL.n263 B 0.011323f
C362 VTAIL.n264 B 0.025276f
C363 VTAIL.n265 B 0.025276f
C364 VTAIL.n266 B 0.011323f
C365 VTAIL.n267 B 0.010694f
C366 VTAIL.n268 B 0.019901f
C367 VTAIL.n269 B 0.019901f
C368 VTAIL.n270 B 0.010694f
C369 VTAIL.n271 B 0.011323f
C370 VTAIL.n272 B 0.025276f
C371 VTAIL.n273 B 0.025276f
C372 VTAIL.n274 B 0.011323f
C373 VTAIL.n275 B 0.010694f
C374 VTAIL.n276 B 0.019901f
C375 VTAIL.n277 B 0.019901f
C376 VTAIL.n278 B 0.010694f
C377 VTAIL.n279 B 0.011008f
C378 VTAIL.n280 B 0.011008f
C379 VTAIL.n281 B 0.025276f
C380 VTAIL.n282 B 0.025276f
C381 VTAIL.n283 B 0.011323f
C382 VTAIL.n284 B 0.010694f
C383 VTAIL.n285 B 0.019901f
C384 VTAIL.n286 B 0.019901f
C385 VTAIL.n287 B 0.010694f
C386 VTAIL.n288 B 0.011323f
C387 VTAIL.n289 B 0.025276f
C388 VTAIL.n290 B 0.055194f
C389 VTAIL.n291 B 0.011323f
C390 VTAIL.n292 B 0.010694f
C391 VTAIL.n293 B 0.048718f
C392 VTAIL.n294 B 0.031013f
C393 VTAIL.n295 B 0.189625f
C394 VTAIL.n296 B 0.028241f
C395 VTAIL.n297 B 0.019901f
C396 VTAIL.n298 B 0.010694f
C397 VTAIL.n299 B 0.025276f
C398 VTAIL.n300 B 0.011323f
C399 VTAIL.n301 B 0.019901f
C400 VTAIL.n302 B 0.010694f
C401 VTAIL.n303 B 0.025276f
C402 VTAIL.n304 B 0.011323f
C403 VTAIL.n305 B 0.019901f
C404 VTAIL.n306 B 0.010694f
C405 VTAIL.n307 B 0.025276f
C406 VTAIL.n308 B 0.025276f
C407 VTAIL.n309 B 0.011323f
C408 VTAIL.n310 B 0.019901f
C409 VTAIL.n311 B 0.010694f
C410 VTAIL.n312 B 0.025276f
C411 VTAIL.n313 B 0.011323f
C412 VTAIL.n314 B 0.134163f
C413 VTAIL.t15 B 0.04256f
C414 VTAIL.n315 B 0.018957f
C415 VTAIL.n316 B 0.017868f
C416 VTAIL.n317 B 0.010694f
C417 VTAIL.n318 B 0.89597f
C418 VTAIL.n319 B 0.019901f
C419 VTAIL.n320 B 0.010694f
C420 VTAIL.n321 B 0.011323f
C421 VTAIL.n322 B 0.025276f
C422 VTAIL.n323 B 0.025276f
C423 VTAIL.n324 B 0.011323f
C424 VTAIL.n325 B 0.010694f
C425 VTAIL.n326 B 0.019901f
C426 VTAIL.n327 B 0.019901f
C427 VTAIL.n328 B 0.010694f
C428 VTAIL.n329 B 0.011323f
C429 VTAIL.n330 B 0.025276f
C430 VTAIL.n331 B 0.025276f
C431 VTAIL.n332 B 0.011323f
C432 VTAIL.n333 B 0.010694f
C433 VTAIL.n334 B 0.019901f
C434 VTAIL.n335 B 0.019901f
C435 VTAIL.n336 B 0.010694f
C436 VTAIL.n337 B 0.011008f
C437 VTAIL.n338 B 0.011008f
C438 VTAIL.n339 B 0.025276f
C439 VTAIL.n340 B 0.025276f
C440 VTAIL.n341 B 0.011323f
C441 VTAIL.n342 B 0.010694f
C442 VTAIL.n343 B 0.019901f
C443 VTAIL.n344 B 0.019901f
C444 VTAIL.n345 B 0.010694f
C445 VTAIL.n346 B 0.011323f
C446 VTAIL.n347 B 0.025276f
C447 VTAIL.n348 B 0.055194f
C448 VTAIL.n349 B 0.011323f
C449 VTAIL.n350 B 0.010694f
C450 VTAIL.n351 B 0.048718f
C451 VTAIL.n352 B 0.031013f
C452 VTAIL.n353 B 0.189625f
C453 VTAIL.t13 B 0.169529f
C454 VTAIL.t9 B 0.169529f
C455 VTAIL.n354 B 1.44634f
C456 VTAIL.n355 B 0.472274f
C457 VTAIL.n356 B 0.028241f
C458 VTAIL.n357 B 0.019901f
C459 VTAIL.n358 B 0.010694f
C460 VTAIL.n359 B 0.025276f
C461 VTAIL.n360 B 0.011323f
C462 VTAIL.n361 B 0.019901f
C463 VTAIL.n362 B 0.010694f
C464 VTAIL.n363 B 0.025276f
C465 VTAIL.n364 B 0.011323f
C466 VTAIL.n365 B 0.019901f
C467 VTAIL.n366 B 0.010694f
C468 VTAIL.n367 B 0.025276f
C469 VTAIL.n368 B 0.025276f
C470 VTAIL.n369 B 0.011323f
C471 VTAIL.n370 B 0.019901f
C472 VTAIL.n371 B 0.010694f
C473 VTAIL.n372 B 0.025276f
C474 VTAIL.n373 B 0.011323f
C475 VTAIL.n374 B 0.134163f
C476 VTAIL.t10 B 0.04256f
C477 VTAIL.n375 B 0.018957f
C478 VTAIL.n376 B 0.017868f
C479 VTAIL.n377 B 0.010694f
C480 VTAIL.n378 B 0.89597f
C481 VTAIL.n379 B 0.019901f
C482 VTAIL.n380 B 0.010694f
C483 VTAIL.n381 B 0.011323f
C484 VTAIL.n382 B 0.025276f
C485 VTAIL.n383 B 0.025276f
C486 VTAIL.n384 B 0.011323f
C487 VTAIL.n385 B 0.010694f
C488 VTAIL.n386 B 0.019901f
C489 VTAIL.n387 B 0.019901f
C490 VTAIL.n388 B 0.010694f
C491 VTAIL.n389 B 0.011323f
C492 VTAIL.n390 B 0.025276f
C493 VTAIL.n391 B 0.025276f
C494 VTAIL.n392 B 0.011323f
C495 VTAIL.n393 B 0.010694f
C496 VTAIL.n394 B 0.019901f
C497 VTAIL.n395 B 0.019901f
C498 VTAIL.n396 B 0.010694f
C499 VTAIL.n397 B 0.011008f
C500 VTAIL.n398 B 0.011008f
C501 VTAIL.n399 B 0.025276f
C502 VTAIL.n400 B 0.025276f
C503 VTAIL.n401 B 0.011323f
C504 VTAIL.n402 B 0.010694f
C505 VTAIL.n403 B 0.019901f
C506 VTAIL.n404 B 0.019901f
C507 VTAIL.n405 B 0.010694f
C508 VTAIL.n406 B 0.011323f
C509 VTAIL.n407 B 0.025276f
C510 VTAIL.n408 B 0.055194f
C511 VTAIL.n409 B 0.011323f
C512 VTAIL.n410 B 0.010694f
C513 VTAIL.n411 B 0.048718f
C514 VTAIL.n412 B 0.031013f
C515 VTAIL.n413 B 1.16671f
C516 VTAIL.n414 B 0.028241f
C517 VTAIL.n415 B 0.019901f
C518 VTAIL.n416 B 0.010694f
C519 VTAIL.n417 B 0.025276f
C520 VTAIL.n418 B 0.011323f
C521 VTAIL.n419 B 0.019901f
C522 VTAIL.n420 B 0.010694f
C523 VTAIL.n421 B 0.025276f
C524 VTAIL.n422 B 0.011323f
C525 VTAIL.n423 B 0.019901f
C526 VTAIL.n424 B 0.010694f
C527 VTAIL.n425 B 0.025276f
C528 VTAIL.n426 B 0.011323f
C529 VTAIL.n427 B 0.019901f
C530 VTAIL.n428 B 0.010694f
C531 VTAIL.n429 B 0.025276f
C532 VTAIL.n430 B 0.011323f
C533 VTAIL.n431 B 0.134163f
C534 VTAIL.t6 B 0.04256f
C535 VTAIL.n432 B 0.018957f
C536 VTAIL.n433 B 0.017868f
C537 VTAIL.n434 B 0.010694f
C538 VTAIL.n435 B 0.89597f
C539 VTAIL.n436 B 0.019901f
C540 VTAIL.n437 B 0.010694f
C541 VTAIL.n438 B 0.011323f
C542 VTAIL.n439 B 0.025276f
C543 VTAIL.n440 B 0.025276f
C544 VTAIL.n441 B 0.011323f
C545 VTAIL.n442 B 0.010694f
C546 VTAIL.n443 B 0.019901f
C547 VTAIL.n444 B 0.019901f
C548 VTAIL.n445 B 0.010694f
C549 VTAIL.n446 B 0.011323f
C550 VTAIL.n447 B 0.025276f
C551 VTAIL.n448 B 0.025276f
C552 VTAIL.n449 B 0.025276f
C553 VTAIL.n450 B 0.011323f
C554 VTAIL.n451 B 0.010694f
C555 VTAIL.n452 B 0.019901f
C556 VTAIL.n453 B 0.019901f
C557 VTAIL.n454 B 0.010694f
C558 VTAIL.n455 B 0.011008f
C559 VTAIL.n456 B 0.011008f
C560 VTAIL.n457 B 0.025276f
C561 VTAIL.n458 B 0.025276f
C562 VTAIL.n459 B 0.011323f
C563 VTAIL.n460 B 0.010694f
C564 VTAIL.n461 B 0.019901f
C565 VTAIL.n462 B 0.019901f
C566 VTAIL.n463 B 0.010694f
C567 VTAIL.n464 B 0.011323f
C568 VTAIL.n465 B 0.025276f
C569 VTAIL.n466 B 0.055194f
C570 VTAIL.n467 B 0.011323f
C571 VTAIL.n468 B 0.010694f
C572 VTAIL.n469 B 0.048718f
C573 VTAIL.n470 B 0.031013f
C574 VTAIL.n471 B 1.16298f
C575 VDD1.t0 B 0.210137f
C576 VDD1.t2 B 0.210137f
C577 VDD1.n0 B 1.86993f
C578 VDD1.t1 B 0.210137f
C579 VDD1.t7 B 0.210137f
C580 VDD1.n1 B 1.86898f
C581 VDD1.t4 B 0.210137f
C582 VDD1.t3 B 0.210137f
C583 VDD1.n2 B 1.86898f
C584 VDD1.n3 B 2.98967f
C585 VDD1.t6 B 0.210137f
C586 VDD1.t5 B 0.210137f
C587 VDD1.n4 B 1.86148f
C588 VDD1.n5 B 2.71615f
C589 VP.n0 B 0.033155f
C590 VP.t3 B 1.63454f
C591 VP.n1 B 0.021125f
C592 VP.n2 B 0.025149f
C593 VP.t4 B 1.63454f
C594 VP.n3 B 0.049721f
C595 VP.n4 B 0.025149f
C596 VP.t7 B 1.63454f
C597 VP.n5 B 0.585255f
C598 VP.n6 B 0.025149f
C599 VP.n7 B 0.048115f
C600 VP.n8 B 0.033155f
C601 VP.t5 B 1.63454f
C602 VP.n9 B 0.021125f
C603 VP.n10 B 0.025149f
C604 VP.t6 B 1.63454f
C605 VP.n11 B 0.049721f
C606 VP.n12 B 0.025149f
C607 VP.t2 B 1.63454f
C608 VP.n13 B 0.651144f
C609 VP.t0 B 1.79387f
C610 VP.n14 B 0.64f
C611 VP.n15 B 0.214623f
C612 VP.n16 B 0.036276f
C613 VP.n17 B 0.049721f
C614 VP.n18 B 0.020312f
C615 VP.n19 B 0.025149f
C616 VP.n20 B 0.025149f
C617 VP.n21 B 0.025149f
C618 VP.n22 B 0.036276f
C619 VP.n23 B 0.585255f
C620 VP.n24 B 0.033974f
C621 VP.n25 B 0.050513f
C622 VP.n26 B 0.025149f
C623 VP.n27 B 0.025149f
C624 VP.n28 B 0.025149f
C625 VP.n29 B 0.048115f
C626 VP.n30 B 0.038579f
C627 VP.n31 B 0.664296f
C628 VP.n32 B 1.31883f
C629 VP.n33 B 1.33763f
C630 VP.t1 B 1.63454f
C631 VP.n34 B 0.664296f
C632 VP.n35 B 0.038579f
C633 VP.n36 B 0.033155f
C634 VP.n37 B 0.025149f
C635 VP.n38 B 0.025149f
C636 VP.n39 B 0.021125f
C637 VP.n40 B 0.050513f
C638 VP.n41 B 0.033974f
C639 VP.n42 B 0.025149f
C640 VP.n43 B 0.025149f
C641 VP.n44 B 0.036276f
C642 VP.n45 B 0.049721f
C643 VP.n46 B 0.020312f
C644 VP.n47 B 0.025149f
C645 VP.n48 B 0.025149f
C646 VP.n49 B 0.025149f
C647 VP.n50 B 0.036276f
C648 VP.n51 B 0.585255f
C649 VP.n52 B 0.033974f
C650 VP.n53 B 0.050513f
C651 VP.n54 B 0.025149f
C652 VP.n55 B 0.025149f
C653 VP.n56 B 0.025149f
C654 VP.n57 B 0.048115f
C655 VP.n58 B 0.038579f
C656 VP.n59 B 0.664296f
C657 VP.n60 B 0.034356f
.ends

