* NGSPICE file created from diff_pair_sample_1566.ext - technology: sky130A

.subckt diff_pair_sample_1566 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=2.8017 pd=17.31 as=2.8017 ps=17.31 w=16.98 l=2.78
X1 VTAIL.t8 VP.t1 VDD1.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=2.8017 pd=17.31 as=2.8017 ps=17.31 w=16.98 l=2.78
X2 VDD1.t5 VP.t2 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=2.8017 pd=17.31 as=2.8017 ps=17.31 w=16.98 l=2.78
X3 VTAIL.t0 VN.t0 VDD2.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=2.8017 pd=17.31 as=2.8017 ps=17.31 w=16.98 l=2.78
X4 VTAIL.t5 VN.t1 VDD2.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.6222 pd=34.74 as=2.8017 ps=17.31 w=16.98 l=2.78
X5 VDD2.t5 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.8017 pd=17.31 as=6.6222 ps=34.74 w=16.98 l=2.78
X6 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=6.6222 pd=34.74 as=0 ps=0 w=16.98 l=2.78
X7 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=6.6222 pd=34.74 as=0 ps=0 w=16.98 l=2.78
X8 VDD1.t4 VP.t3 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=2.8017 pd=17.31 as=6.6222 ps=34.74 w=16.98 l=2.78
X9 VTAIL.t12 VP.t4 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=6.6222 pd=34.74 as=2.8017 ps=17.31 w=16.98 l=2.78
X10 VDD2.t4 VN.t3 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.8017 pd=17.31 as=6.6222 ps=34.74 w=16.98 l=2.78
X11 VTAIL.t3 VN.t4 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.8017 pd=17.31 as=2.8017 ps=17.31 w=16.98 l=2.78
X12 VTAIL.t14 VP.t5 VDD1.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=6.6222 pd=34.74 as=2.8017 ps=17.31 w=16.98 l=2.78
X13 VDD2.t2 VN.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.8017 pd=17.31 as=2.8017 ps=17.31 w=16.98 l=2.78
X14 VTAIL.t13 VP.t6 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=2.8017 pd=17.31 as=2.8017 ps=17.31 w=16.98 l=2.78
X15 VDD1.t0 VP.t7 VTAIL.t15 B.t2 sky130_fd_pr__nfet_01v8 ad=2.8017 pd=17.31 as=6.6222 ps=34.74 w=16.98 l=2.78
X16 VTAIL.t4 VN.t6 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=6.6222 pd=34.74 as=2.8017 ps=17.31 w=16.98 l=2.78
X17 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=6.6222 pd=34.74 as=0 ps=0 w=16.98 l=2.78
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.6222 pd=34.74 as=0 ps=0 w=16.98 l=2.78
X19 VDD2.t0 VN.t7 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.8017 pd=17.31 as=2.8017 ps=17.31 w=16.98 l=2.78
R0 VP.n19 VP.t5 180.248
R1 VP.n21 VP.n20 161.3
R2 VP.n22 VP.n17 161.3
R3 VP.n24 VP.n23 161.3
R4 VP.n25 VP.n16 161.3
R5 VP.n27 VP.n26 161.3
R6 VP.n28 VP.n15 161.3
R7 VP.n30 VP.n29 161.3
R8 VP.n32 VP.n31 161.3
R9 VP.n33 VP.n13 161.3
R10 VP.n35 VP.n34 161.3
R11 VP.n36 VP.n12 161.3
R12 VP.n38 VP.n37 161.3
R13 VP.n39 VP.n11 161.3
R14 VP.n72 VP.n0 161.3
R15 VP.n71 VP.n70 161.3
R16 VP.n69 VP.n1 161.3
R17 VP.n68 VP.n67 161.3
R18 VP.n66 VP.n2 161.3
R19 VP.n65 VP.n64 161.3
R20 VP.n63 VP.n62 161.3
R21 VP.n61 VP.n4 161.3
R22 VP.n60 VP.n59 161.3
R23 VP.n58 VP.n5 161.3
R24 VP.n57 VP.n56 161.3
R25 VP.n55 VP.n6 161.3
R26 VP.n54 VP.n53 161.3
R27 VP.n52 VP.n51 161.3
R28 VP.n50 VP.n8 161.3
R29 VP.n49 VP.n48 161.3
R30 VP.n47 VP.n9 161.3
R31 VP.n46 VP.n45 161.3
R32 VP.n44 VP.n10 161.3
R33 VP.n43 VP.t4 147.202
R34 VP.n7 VP.t0 147.202
R35 VP.n3 VP.t6 147.202
R36 VP.n73 VP.t3 147.202
R37 VP.n40 VP.t7 147.202
R38 VP.n14 VP.t1 147.202
R39 VP.n18 VP.t2 147.202
R40 VP.n43 VP.n42 102.793
R41 VP.n74 VP.n73 102.793
R42 VP.n41 VP.n40 102.793
R43 VP.n19 VP.n18 70.4561
R44 VP.n42 VP.n41 55.5451
R45 VP.n49 VP.n9 51.2335
R46 VP.n67 VP.n1 51.2335
R47 VP.n34 VP.n12 51.2335
R48 VP.n56 VP.n5 40.577
R49 VP.n60 VP.n5 40.577
R50 VP.n27 VP.n16 40.577
R51 VP.n23 VP.n16 40.577
R52 VP.n50 VP.n49 29.9206
R53 VP.n67 VP.n66 29.9206
R54 VP.n34 VP.n33 29.9206
R55 VP.n45 VP.n44 24.5923
R56 VP.n45 VP.n9 24.5923
R57 VP.n51 VP.n50 24.5923
R58 VP.n55 VP.n54 24.5923
R59 VP.n56 VP.n55 24.5923
R60 VP.n61 VP.n60 24.5923
R61 VP.n62 VP.n61 24.5923
R62 VP.n66 VP.n65 24.5923
R63 VP.n71 VP.n1 24.5923
R64 VP.n72 VP.n71 24.5923
R65 VP.n38 VP.n12 24.5923
R66 VP.n39 VP.n38 24.5923
R67 VP.n28 VP.n27 24.5923
R68 VP.n29 VP.n28 24.5923
R69 VP.n33 VP.n32 24.5923
R70 VP.n22 VP.n21 24.5923
R71 VP.n23 VP.n22 24.5923
R72 VP.n51 VP.n7 21.8872
R73 VP.n65 VP.n3 21.8872
R74 VP.n32 VP.n14 21.8872
R75 VP.n44 VP.n43 8.11581
R76 VP.n73 VP.n72 8.11581
R77 VP.n40 VP.n39 8.11581
R78 VP.n20 VP.n19 6.95301
R79 VP.n54 VP.n7 2.7056
R80 VP.n62 VP.n3 2.7056
R81 VP.n29 VP.n14 2.7056
R82 VP.n21 VP.n18 2.7056
R83 VP.n41 VP.n11 0.278335
R84 VP.n42 VP.n10 0.278335
R85 VP.n74 VP.n0 0.278335
R86 VP.n20 VP.n17 0.189894
R87 VP.n24 VP.n17 0.189894
R88 VP.n25 VP.n24 0.189894
R89 VP.n26 VP.n25 0.189894
R90 VP.n26 VP.n15 0.189894
R91 VP.n30 VP.n15 0.189894
R92 VP.n31 VP.n30 0.189894
R93 VP.n31 VP.n13 0.189894
R94 VP.n35 VP.n13 0.189894
R95 VP.n36 VP.n35 0.189894
R96 VP.n37 VP.n36 0.189894
R97 VP.n37 VP.n11 0.189894
R98 VP.n46 VP.n10 0.189894
R99 VP.n47 VP.n46 0.189894
R100 VP.n48 VP.n47 0.189894
R101 VP.n48 VP.n8 0.189894
R102 VP.n52 VP.n8 0.189894
R103 VP.n53 VP.n52 0.189894
R104 VP.n53 VP.n6 0.189894
R105 VP.n57 VP.n6 0.189894
R106 VP.n58 VP.n57 0.189894
R107 VP.n59 VP.n58 0.189894
R108 VP.n59 VP.n4 0.189894
R109 VP.n63 VP.n4 0.189894
R110 VP.n64 VP.n63 0.189894
R111 VP.n64 VP.n2 0.189894
R112 VP.n68 VP.n2 0.189894
R113 VP.n69 VP.n68 0.189894
R114 VP.n70 VP.n69 0.189894
R115 VP.n70 VP.n0 0.189894
R116 VP VP.n74 0.153485
R117 VTAIL.n754 VTAIL.n666 289.615
R118 VTAIL.n90 VTAIL.n2 289.615
R119 VTAIL.n184 VTAIL.n96 289.615
R120 VTAIL.n280 VTAIL.n192 289.615
R121 VTAIL.n660 VTAIL.n572 289.615
R122 VTAIL.n564 VTAIL.n476 289.615
R123 VTAIL.n470 VTAIL.n382 289.615
R124 VTAIL.n374 VTAIL.n286 289.615
R125 VTAIL.n697 VTAIL.n696 185
R126 VTAIL.n694 VTAIL.n693 185
R127 VTAIL.n703 VTAIL.n702 185
R128 VTAIL.n705 VTAIL.n704 185
R129 VTAIL.n690 VTAIL.n689 185
R130 VTAIL.n711 VTAIL.n710 185
R131 VTAIL.n713 VTAIL.n712 185
R132 VTAIL.n686 VTAIL.n685 185
R133 VTAIL.n719 VTAIL.n718 185
R134 VTAIL.n721 VTAIL.n720 185
R135 VTAIL.n682 VTAIL.n681 185
R136 VTAIL.n727 VTAIL.n726 185
R137 VTAIL.n729 VTAIL.n728 185
R138 VTAIL.n678 VTAIL.n677 185
R139 VTAIL.n735 VTAIL.n734 185
R140 VTAIL.n738 VTAIL.n737 185
R141 VTAIL.n736 VTAIL.n674 185
R142 VTAIL.n743 VTAIL.n673 185
R143 VTAIL.n745 VTAIL.n744 185
R144 VTAIL.n747 VTAIL.n746 185
R145 VTAIL.n670 VTAIL.n669 185
R146 VTAIL.n753 VTAIL.n752 185
R147 VTAIL.n755 VTAIL.n754 185
R148 VTAIL.n33 VTAIL.n32 185
R149 VTAIL.n30 VTAIL.n29 185
R150 VTAIL.n39 VTAIL.n38 185
R151 VTAIL.n41 VTAIL.n40 185
R152 VTAIL.n26 VTAIL.n25 185
R153 VTAIL.n47 VTAIL.n46 185
R154 VTAIL.n49 VTAIL.n48 185
R155 VTAIL.n22 VTAIL.n21 185
R156 VTAIL.n55 VTAIL.n54 185
R157 VTAIL.n57 VTAIL.n56 185
R158 VTAIL.n18 VTAIL.n17 185
R159 VTAIL.n63 VTAIL.n62 185
R160 VTAIL.n65 VTAIL.n64 185
R161 VTAIL.n14 VTAIL.n13 185
R162 VTAIL.n71 VTAIL.n70 185
R163 VTAIL.n74 VTAIL.n73 185
R164 VTAIL.n72 VTAIL.n10 185
R165 VTAIL.n79 VTAIL.n9 185
R166 VTAIL.n81 VTAIL.n80 185
R167 VTAIL.n83 VTAIL.n82 185
R168 VTAIL.n6 VTAIL.n5 185
R169 VTAIL.n89 VTAIL.n88 185
R170 VTAIL.n91 VTAIL.n90 185
R171 VTAIL.n127 VTAIL.n126 185
R172 VTAIL.n124 VTAIL.n123 185
R173 VTAIL.n133 VTAIL.n132 185
R174 VTAIL.n135 VTAIL.n134 185
R175 VTAIL.n120 VTAIL.n119 185
R176 VTAIL.n141 VTAIL.n140 185
R177 VTAIL.n143 VTAIL.n142 185
R178 VTAIL.n116 VTAIL.n115 185
R179 VTAIL.n149 VTAIL.n148 185
R180 VTAIL.n151 VTAIL.n150 185
R181 VTAIL.n112 VTAIL.n111 185
R182 VTAIL.n157 VTAIL.n156 185
R183 VTAIL.n159 VTAIL.n158 185
R184 VTAIL.n108 VTAIL.n107 185
R185 VTAIL.n165 VTAIL.n164 185
R186 VTAIL.n168 VTAIL.n167 185
R187 VTAIL.n166 VTAIL.n104 185
R188 VTAIL.n173 VTAIL.n103 185
R189 VTAIL.n175 VTAIL.n174 185
R190 VTAIL.n177 VTAIL.n176 185
R191 VTAIL.n100 VTAIL.n99 185
R192 VTAIL.n183 VTAIL.n182 185
R193 VTAIL.n185 VTAIL.n184 185
R194 VTAIL.n223 VTAIL.n222 185
R195 VTAIL.n220 VTAIL.n219 185
R196 VTAIL.n229 VTAIL.n228 185
R197 VTAIL.n231 VTAIL.n230 185
R198 VTAIL.n216 VTAIL.n215 185
R199 VTAIL.n237 VTAIL.n236 185
R200 VTAIL.n239 VTAIL.n238 185
R201 VTAIL.n212 VTAIL.n211 185
R202 VTAIL.n245 VTAIL.n244 185
R203 VTAIL.n247 VTAIL.n246 185
R204 VTAIL.n208 VTAIL.n207 185
R205 VTAIL.n253 VTAIL.n252 185
R206 VTAIL.n255 VTAIL.n254 185
R207 VTAIL.n204 VTAIL.n203 185
R208 VTAIL.n261 VTAIL.n260 185
R209 VTAIL.n264 VTAIL.n263 185
R210 VTAIL.n262 VTAIL.n200 185
R211 VTAIL.n269 VTAIL.n199 185
R212 VTAIL.n271 VTAIL.n270 185
R213 VTAIL.n273 VTAIL.n272 185
R214 VTAIL.n196 VTAIL.n195 185
R215 VTAIL.n279 VTAIL.n278 185
R216 VTAIL.n281 VTAIL.n280 185
R217 VTAIL.n661 VTAIL.n660 185
R218 VTAIL.n659 VTAIL.n658 185
R219 VTAIL.n576 VTAIL.n575 185
R220 VTAIL.n653 VTAIL.n652 185
R221 VTAIL.n651 VTAIL.n650 185
R222 VTAIL.n649 VTAIL.n579 185
R223 VTAIL.n583 VTAIL.n580 185
R224 VTAIL.n644 VTAIL.n643 185
R225 VTAIL.n642 VTAIL.n641 185
R226 VTAIL.n585 VTAIL.n584 185
R227 VTAIL.n636 VTAIL.n635 185
R228 VTAIL.n634 VTAIL.n633 185
R229 VTAIL.n589 VTAIL.n588 185
R230 VTAIL.n628 VTAIL.n627 185
R231 VTAIL.n626 VTAIL.n625 185
R232 VTAIL.n593 VTAIL.n592 185
R233 VTAIL.n620 VTAIL.n619 185
R234 VTAIL.n618 VTAIL.n617 185
R235 VTAIL.n597 VTAIL.n596 185
R236 VTAIL.n612 VTAIL.n611 185
R237 VTAIL.n610 VTAIL.n609 185
R238 VTAIL.n601 VTAIL.n600 185
R239 VTAIL.n604 VTAIL.n603 185
R240 VTAIL.n565 VTAIL.n564 185
R241 VTAIL.n563 VTAIL.n562 185
R242 VTAIL.n480 VTAIL.n479 185
R243 VTAIL.n557 VTAIL.n556 185
R244 VTAIL.n555 VTAIL.n554 185
R245 VTAIL.n553 VTAIL.n483 185
R246 VTAIL.n487 VTAIL.n484 185
R247 VTAIL.n548 VTAIL.n547 185
R248 VTAIL.n546 VTAIL.n545 185
R249 VTAIL.n489 VTAIL.n488 185
R250 VTAIL.n540 VTAIL.n539 185
R251 VTAIL.n538 VTAIL.n537 185
R252 VTAIL.n493 VTAIL.n492 185
R253 VTAIL.n532 VTAIL.n531 185
R254 VTAIL.n530 VTAIL.n529 185
R255 VTAIL.n497 VTAIL.n496 185
R256 VTAIL.n524 VTAIL.n523 185
R257 VTAIL.n522 VTAIL.n521 185
R258 VTAIL.n501 VTAIL.n500 185
R259 VTAIL.n516 VTAIL.n515 185
R260 VTAIL.n514 VTAIL.n513 185
R261 VTAIL.n505 VTAIL.n504 185
R262 VTAIL.n508 VTAIL.n507 185
R263 VTAIL.n471 VTAIL.n470 185
R264 VTAIL.n469 VTAIL.n468 185
R265 VTAIL.n386 VTAIL.n385 185
R266 VTAIL.n463 VTAIL.n462 185
R267 VTAIL.n461 VTAIL.n460 185
R268 VTAIL.n459 VTAIL.n389 185
R269 VTAIL.n393 VTAIL.n390 185
R270 VTAIL.n454 VTAIL.n453 185
R271 VTAIL.n452 VTAIL.n451 185
R272 VTAIL.n395 VTAIL.n394 185
R273 VTAIL.n446 VTAIL.n445 185
R274 VTAIL.n444 VTAIL.n443 185
R275 VTAIL.n399 VTAIL.n398 185
R276 VTAIL.n438 VTAIL.n437 185
R277 VTAIL.n436 VTAIL.n435 185
R278 VTAIL.n403 VTAIL.n402 185
R279 VTAIL.n430 VTAIL.n429 185
R280 VTAIL.n428 VTAIL.n427 185
R281 VTAIL.n407 VTAIL.n406 185
R282 VTAIL.n422 VTAIL.n421 185
R283 VTAIL.n420 VTAIL.n419 185
R284 VTAIL.n411 VTAIL.n410 185
R285 VTAIL.n414 VTAIL.n413 185
R286 VTAIL.n375 VTAIL.n374 185
R287 VTAIL.n373 VTAIL.n372 185
R288 VTAIL.n290 VTAIL.n289 185
R289 VTAIL.n367 VTAIL.n366 185
R290 VTAIL.n365 VTAIL.n364 185
R291 VTAIL.n363 VTAIL.n293 185
R292 VTAIL.n297 VTAIL.n294 185
R293 VTAIL.n358 VTAIL.n357 185
R294 VTAIL.n356 VTAIL.n355 185
R295 VTAIL.n299 VTAIL.n298 185
R296 VTAIL.n350 VTAIL.n349 185
R297 VTAIL.n348 VTAIL.n347 185
R298 VTAIL.n303 VTAIL.n302 185
R299 VTAIL.n342 VTAIL.n341 185
R300 VTAIL.n340 VTAIL.n339 185
R301 VTAIL.n307 VTAIL.n306 185
R302 VTAIL.n334 VTAIL.n333 185
R303 VTAIL.n332 VTAIL.n331 185
R304 VTAIL.n311 VTAIL.n310 185
R305 VTAIL.n326 VTAIL.n325 185
R306 VTAIL.n324 VTAIL.n323 185
R307 VTAIL.n315 VTAIL.n314 185
R308 VTAIL.n318 VTAIL.n317 185
R309 VTAIL.t15 VTAIL.n602 147.659
R310 VTAIL.t14 VTAIL.n506 147.659
R311 VTAIL.t7 VTAIL.n412 147.659
R312 VTAIL.t4 VTAIL.n316 147.659
R313 VTAIL.t2 VTAIL.n695 147.659
R314 VTAIL.t5 VTAIL.n31 147.659
R315 VTAIL.t10 VTAIL.n125 147.659
R316 VTAIL.t12 VTAIL.n221 147.659
R317 VTAIL.n696 VTAIL.n693 104.615
R318 VTAIL.n703 VTAIL.n693 104.615
R319 VTAIL.n704 VTAIL.n703 104.615
R320 VTAIL.n704 VTAIL.n689 104.615
R321 VTAIL.n711 VTAIL.n689 104.615
R322 VTAIL.n712 VTAIL.n711 104.615
R323 VTAIL.n712 VTAIL.n685 104.615
R324 VTAIL.n719 VTAIL.n685 104.615
R325 VTAIL.n720 VTAIL.n719 104.615
R326 VTAIL.n720 VTAIL.n681 104.615
R327 VTAIL.n727 VTAIL.n681 104.615
R328 VTAIL.n728 VTAIL.n727 104.615
R329 VTAIL.n728 VTAIL.n677 104.615
R330 VTAIL.n735 VTAIL.n677 104.615
R331 VTAIL.n737 VTAIL.n735 104.615
R332 VTAIL.n737 VTAIL.n736 104.615
R333 VTAIL.n736 VTAIL.n673 104.615
R334 VTAIL.n745 VTAIL.n673 104.615
R335 VTAIL.n746 VTAIL.n745 104.615
R336 VTAIL.n746 VTAIL.n669 104.615
R337 VTAIL.n753 VTAIL.n669 104.615
R338 VTAIL.n754 VTAIL.n753 104.615
R339 VTAIL.n32 VTAIL.n29 104.615
R340 VTAIL.n39 VTAIL.n29 104.615
R341 VTAIL.n40 VTAIL.n39 104.615
R342 VTAIL.n40 VTAIL.n25 104.615
R343 VTAIL.n47 VTAIL.n25 104.615
R344 VTAIL.n48 VTAIL.n47 104.615
R345 VTAIL.n48 VTAIL.n21 104.615
R346 VTAIL.n55 VTAIL.n21 104.615
R347 VTAIL.n56 VTAIL.n55 104.615
R348 VTAIL.n56 VTAIL.n17 104.615
R349 VTAIL.n63 VTAIL.n17 104.615
R350 VTAIL.n64 VTAIL.n63 104.615
R351 VTAIL.n64 VTAIL.n13 104.615
R352 VTAIL.n71 VTAIL.n13 104.615
R353 VTAIL.n73 VTAIL.n71 104.615
R354 VTAIL.n73 VTAIL.n72 104.615
R355 VTAIL.n72 VTAIL.n9 104.615
R356 VTAIL.n81 VTAIL.n9 104.615
R357 VTAIL.n82 VTAIL.n81 104.615
R358 VTAIL.n82 VTAIL.n5 104.615
R359 VTAIL.n89 VTAIL.n5 104.615
R360 VTAIL.n90 VTAIL.n89 104.615
R361 VTAIL.n126 VTAIL.n123 104.615
R362 VTAIL.n133 VTAIL.n123 104.615
R363 VTAIL.n134 VTAIL.n133 104.615
R364 VTAIL.n134 VTAIL.n119 104.615
R365 VTAIL.n141 VTAIL.n119 104.615
R366 VTAIL.n142 VTAIL.n141 104.615
R367 VTAIL.n142 VTAIL.n115 104.615
R368 VTAIL.n149 VTAIL.n115 104.615
R369 VTAIL.n150 VTAIL.n149 104.615
R370 VTAIL.n150 VTAIL.n111 104.615
R371 VTAIL.n157 VTAIL.n111 104.615
R372 VTAIL.n158 VTAIL.n157 104.615
R373 VTAIL.n158 VTAIL.n107 104.615
R374 VTAIL.n165 VTAIL.n107 104.615
R375 VTAIL.n167 VTAIL.n165 104.615
R376 VTAIL.n167 VTAIL.n166 104.615
R377 VTAIL.n166 VTAIL.n103 104.615
R378 VTAIL.n175 VTAIL.n103 104.615
R379 VTAIL.n176 VTAIL.n175 104.615
R380 VTAIL.n176 VTAIL.n99 104.615
R381 VTAIL.n183 VTAIL.n99 104.615
R382 VTAIL.n184 VTAIL.n183 104.615
R383 VTAIL.n222 VTAIL.n219 104.615
R384 VTAIL.n229 VTAIL.n219 104.615
R385 VTAIL.n230 VTAIL.n229 104.615
R386 VTAIL.n230 VTAIL.n215 104.615
R387 VTAIL.n237 VTAIL.n215 104.615
R388 VTAIL.n238 VTAIL.n237 104.615
R389 VTAIL.n238 VTAIL.n211 104.615
R390 VTAIL.n245 VTAIL.n211 104.615
R391 VTAIL.n246 VTAIL.n245 104.615
R392 VTAIL.n246 VTAIL.n207 104.615
R393 VTAIL.n253 VTAIL.n207 104.615
R394 VTAIL.n254 VTAIL.n253 104.615
R395 VTAIL.n254 VTAIL.n203 104.615
R396 VTAIL.n261 VTAIL.n203 104.615
R397 VTAIL.n263 VTAIL.n261 104.615
R398 VTAIL.n263 VTAIL.n262 104.615
R399 VTAIL.n262 VTAIL.n199 104.615
R400 VTAIL.n271 VTAIL.n199 104.615
R401 VTAIL.n272 VTAIL.n271 104.615
R402 VTAIL.n272 VTAIL.n195 104.615
R403 VTAIL.n279 VTAIL.n195 104.615
R404 VTAIL.n280 VTAIL.n279 104.615
R405 VTAIL.n660 VTAIL.n659 104.615
R406 VTAIL.n659 VTAIL.n575 104.615
R407 VTAIL.n652 VTAIL.n575 104.615
R408 VTAIL.n652 VTAIL.n651 104.615
R409 VTAIL.n651 VTAIL.n579 104.615
R410 VTAIL.n583 VTAIL.n579 104.615
R411 VTAIL.n643 VTAIL.n583 104.615
R412 VTAIL.n643 VTAIL.n642 104.615
R413 VTAIL.n642 VTAIL.n584 104.615
R414 VTAIL.n635 VTAIL.n584 104.615
R415 VTAIL.n635 VTAIL.n634 104.615
R416 VTAIL.n634 VTAIL.n588 104.615
R417 VTAIL.n627 VTAIL.n588 104.615
R418 VTAIL.n627 VTAIL.n626 104.615
R419 VTAIL.n626 VTAIL.n592 104.615
R420 VTAIL.n619 VTAIL.n592 104.615
R421 VTAIL.n619 VTAIL.n618 104.615
R422 VTAIL.n618 VTAIL.n596 104.615
R423 VTAIL.n611 VTAIL.n596 104.615
R424 VTAIL.n611 VTAIL.n610 104.615
R425 VTAIL.n610 VTAIL.n600 104.615
R426 VTAIL.n603 VTAIL.n600 104.615
R427 VTAIL.n564 VTAIL.n563 104.615
R428 VTAIL.n563 VTAIL.n479 104.615
R429 VTAIL.n556 VTAIL.n479 104.615
R430 VTAIL.n556 VTAIL.n555 104.615
R431 VTAIL.n555 VTAIL.n483 104.615
R432 VTAIL.n487 VTAIL.n483 104.615
R433 VTAIL.n547 VTAIL.n487 104.615
R434 VTAIL.n547 VTAIL.n546 104.615
R435 VTAIL.n546 VTAIL.n488 104.615
R436 VTAIL.n539 VTAIL.n488 104.615
R437 VTAIL.n539 VTAIL.n538 104.615
R438 VTAIL.n538 VTAIL.n492 104.615
R439 VTAIL.n531 VTAIL.n492 104.615
R440 VTAIL.n531 VTAIL.n530 104.615
R441 VTAIL.n530 VTAIL.n496 104.615
R442 VTAIL.n523 VTAIL.n496 104.615
R443 VTAIL.n523 VTAIL.n522 104.615
R444 VTAIL.n522 VTAIL.n500 104.615
R445 VTAIL.n515 VTAIL.n500 104.615
R446 VTAIL.n515 VTAIL.n514 104.615
R447 VTAIL.n514 VTAIL.n504 104.615
R448 VTAIL.n507 VTAIL.n504 104.615
R449 VTAIL.n470 VTAIL.n469 104.615
R450 VTAIL.n469 VTAIL.n385 104.615
R451 VTAIL.n462 VTAIL.n385 104.615
R452 VTAIL.n462 VTAIL.n461 104.615
R453 VTAIL.n461 VTAIL.n389 104.615
R454 VTAIL.n393 VTAIL.n389 104.615
R455 VTAIL.n453 VTAIL.n393 104.615
R456 VTAIL.n453 VTAIL.n452 104.615
R457 VTAIL.n452 VTAIL.n394 104.615
R458 VTAIL.n445 VTAIL.n394 104.615
R459 VTAIL.n445 VTAIL.n444 104.615
R460 VTAIL.n444 VTAIL.n398 104.615
R461 VTAIL.n437 VTAIL.n398 104.615
R462 VTAIL.n437 VTAIL.n436 104.615
R463 VTAIL.n436 VTAIL.n402 104.615
R464 VTAIL.n429 VTAIL.n402 104.615
R465 VTAIL.n429 VTAIL.n428 104.615
R466 VTAIL.n428 VTAIL.n406 104.615
R467 VTAIL.n421 VTAIL.n406 104.615
R468 VTAIL.n421 VTAIL.n420 104.615
R469 VTAIL.n420 VTAIL.n410 104.615
R470 VTAIL.n413 VTAIL.n410 104.615
R471 VTAIL.n374 VTAIL.n373 104.615
R472 VTAIL.n373 VTAIL.n289 104.615
R473 VTAIL.n366 VTAIL.n289 104.615
R474 VTAIL.n366 VTAIL.n365 104.615
R475 VTAIL.n365 VTAIL.n293 104.615
R476 VTAIL.n297 VTAIL.n293 104.615
R477 VTAIL.n357 VTAIL.n297 104.615
R478 VTAIL.n357 VTAIL.n356 104.615
R479 VTAIL.n356 VTAIL.n298 104.615
R480 VTAIL.n349 VTAIL.n298 104.615
R481 VTAIL.n349 VTAIL.n348 104.615
R482 VTAIL.n348 VTAIL.n302 104.615
R483 VTAIL.n341 VTAIL.n302 104.615
R484 VTAIL.n341 VTAIL.n340 104.615
R485 VTAIL.n340 VTAIL.n306 104.615
R486 VTAIL.n333 VTAIL.n306 104.615
R487 VTAIL.n333 VTAIL.n332 104.615
R488 VTAIL.n332 VTAIL.n310 104.615
R489 VTAIL.n325 VTAIL.n310 104.615
R490 VTAIL.n325 VTAIL.n324 104.615
R491 VTAIL.n324 VTAIL.n314 104.615
R492 VTAIL.n317 VTAIL.n314 104.615
R493 VTAIL.n696 VTAIL.t2 52.3082
R494 VTAIL.n32 VTAIL.t5 52.3082
R495 VTAIL.n126 VTAIL.t10 52.3082
R496 VTAIL.n222 VTAIL.t12 52.3082
R497 VTAIL.n603 VTAIL.t15 52.3082
R498 VTAIL.n507 VTAIL.t14 52.3082
R499 VTAIL.n413 VTAIL.t7 52.3082
R500 VTAIL.n317 VTAIL.t4 52.3082
R501 VTAIL.n571 VTAIL.n570 47.5369
R502 VTAIL.n381 VTAIL.n380 47.5369
R503 VTAIL.n1 VTAIL.n0 47.5368
R504 VTAIL.n191 VTAIL.n190 47.5368
R505 VTAIL.n759 VTAIL.n758 35.6763
R506 VTAIL.n95 VTAIL.n94 35.6763
R507 VTAIL.n189 VTAIL.n188 35.6763
R508 VTAIL.n285 VTAIL.n284 35.6763
R509 VTAIL.n665 VTAIL.n664 35.6763
R510 VTAIL.n569 VTAIL.n568 35.6763
R511 VTAIL.n475 VTAIL.n474 35.6763
R512 VTAIL.n379 VTAIL.n378 35.6763
R513 VTAIL.n759 VTAIL.n665 29.6858
R514 VTAIL.n379 VTAIL.n285 29.6858
R515 VTAIL.n697 VTAIL.n695 15.6677
R516 VTAIL.n33 VTAIL.n31 15.6677
R517 VTAIL.n127 VTAIL.n125 15.6677
R518 VTAIL.n223 VTAIL.n221 15.6677
R519 VTAIL.n604 VTAIL.n602 15.6677
R520 VTAIL.n508 VTAIL.n506 15.6677
R521 VTAIL.n414 VTAIL.n412 15.6677
R522 VTAIL.n318 VTAIL.n316 15.6677
R523 VTAIL.n744 VTAIL.n743 13.1884
R524 VTAIL.n80 VTAIL.n79 13.1884
R525 VTAIL.n174 VTAIL.n173 13.1884
R526 VTAIL.n270 VTAIL.n269 13.1884
R527 VTAIL.n650 VTAIL.n649 13.1884
R528 VTAIL.n554 VTAIL.n553 13.1884
R529 VTAIL.n460 VTAIL.n459 13.1884
R530 VTAIL.n364 VTAIL.n363 13.1884
R531 VTAIL.n698 VTAIL.n694 12.8005
R532 VTAIL.n742 VTAIL.n674 12.8005
R533 VTAIL.n747 VTAIL.n672 12.8005
R534 VTAIL.n34 VTAIL.n30 12.8005
R535 VTAIL.n78 VTAIL.n10 12.8005
R536 VTAIL.n83 VTAIL.n8 12.8005
R537 VTAIL.n128 VTAIL.n124 12.8005
R538 VTAIL.n172 VTAIL.n104 12.8005
R539 VTAIL.n177 VTAIL.n102 12.8005
R540 VTAIL.n224 VTAIL.n220 12.8005
R541 VTAIL.n268 VTAIL.n200 12.8005
R542 VTAIL.n273 VTAIL.n198 12.8005
R543 VTAIL.n653 VTAIL.n578 12.8005
R544 VTAIL.n648 VTAIL.n580 12.8005
R545 VTAIL.n605 VTAIL.n601 12.8005
R546 VTAIL.n557 VTAIL.n482 12.8005
R547 VTAIL.n552 VTAIL.n484 12.8005
R548 VTAIL.n509 VTAIL.n505 12.8005
R549 VTAIL.n463 VTAIL.n388 12.8005
R550 VTAIL.n458 VTAIL.n390 12.8005
R551 VTAIL.n415 VTAIL.n411 12.8005
R552 VTAIL.n367 VTAIL.n292 12.8005
R553 VTAIL.n362 VTAIL.n294 12.8005
R554 VTAIL.n319 VTAIL.n315 12.8005
R555 VTAIL.n702 VTAIL.n701 12.0247
R556 VTAIL.n739 VTAIL.n738 12.0247
R557 VTAIL.n748 VTAIL.n670 12.0247
R558 VTAIL.n38 VTAIL.n37 12.0247
R559 VTAIL.n75 VTAIL.n74 12.0247
R560 VTAIL.n84 VTAIL.n6 12.0247
R561 VTAIL.n132 VTAIL.n131 12.0247
R562 VTAIL.n169 VTAIL.n168 12.0247
R563 VTAIL.n178 VTAIL.n100 12.0247
R564 VTAIL.n228 VTAIL.n227 12.0247
R565 VTAIL.n265 VTAIL.n264 12.0247
R566 VTAIL.n274 VTAIL.n196 12.0247
R567 VTAIL.n654 VTAIL.n576 12.0247
R568 VTAIL.n645 VTAIL.n644 12.0247
R569 VTAIL.n609 VTAIL.n608 12.0247
R570 VTAIL.n558 VTAIL.n480 12.0247
R571 VTAIL.n549 VTAIL.n548 12.0247
R572 VTAIL.n513 VTAIL.n512 12.0247
R573 VTAIL.n464 VTAIL.n386 12.0247
R574 VTAIL.n455 VTAIL.n454 12.0247
R575 VTAIL.n419 VTAIL.n418 12.0247
R576 VTAIL.n368 VTAIL.n290 12.0247
R577 VTAIL.n359 VTAIL.n358 12.0247
R578 VTAIL.n323 VTAIL.n322 12.0247
R579 VTAIL.n705 VTAIL.n692 11.249
R580 VTAIL.n734 VTAIL.n676 11.249
R581 VTAIL.n752 VTAIL.n751 11.249
R582 VTAIL.n41 VTAIL.n28 11.249
R583 VTAIL.n70 VTAIL.n12 11.249
R584 VTAIL.n88 VTAIL.n87 11.249
R585 VTAIL.n135 VTAIL.n122 11.249
R586 VTAIL.n164 VTAIL.n106 11.249
R587 VTAIL.n182 VTAIL.n181 11.249
R588 VTAIL.n231 VTAIL.n218 11.249
R589 VTAIL.n260 VTAIL.n202 11.249
R590 VTAIL.n278 VTAIL.n277 11.249
R591 VTAIL.n658 VTAIL.n657 11.249
R592 VTAIL.n641 VTAIL.n582 11.249
R593 VTAIL.n612 VTAIL.n599 11.249
R594 VTAIL.n562 VTAIL.n561 11.249
R595 VTAIL.n545 VTAIL.n486 11.249
R596 VTAIL.n516 VTAIL.n503 11.249
R597 VTAIL.n468 VTAIL.n467 11.249
R598 VTAIL.n451 VTAIL.n392 11.249
R599 VTAIL.n422 VTAIL.n409 11.249
R600 VTAIL.n372 VTAIL.n371 11.249
R601 VTAIL.n355 VTAIL.n296 11.249
R602 VTAIL.n326 VTAIL.n313 11.249
R603 VTAIL.n706 VTAIL.n690 10.4732
R604 VTAIL.n733 VTAIL.n678 10.4732
R605 VTAIL.n755 VTAIL.n668 10.4732
R606 VTAIL.n42 VTAIL.n26 10.4732
R607 VTAIL.n69 VTAIL.n14 10.4732
R608 VTAIL.n91 VTAIL.n4 10.4732
R609 VTAIL.n136 VTAIL.n120 10.4732
R610 VTAIL.n163 VTAIL.n108 10.4732
R611 VTAIL.n185 VTAIL.n98 10.4732
R612 VTAIL.n232 VTAIL.n216 10.4732
R613 VTAIL.n259 VTAIL.n204 10.4732
R614 VTAIL.n281 VTAIL.n194 10.4732
R615 VTAIL.n661 VTAIL.n574 10.4732
R616 VTAIL.n640 VTAIL.n585 10.4732
R617 VTAIL.n613 VTAIL.n597 10.4732
R618 VTAIL.n565 VTAIL.n478 10.4732
R619 VTAIL.n544 VTAIL.n489 10.4732
R620 VTAIL.n517 VTAIL.n501 10.4732
R621 VTAIL.n471 VTAIL.n384 10.4732
R622 VTAIL.n450 VTAIL.n395 10.4732
R623 VTAIL.n423 VTAIL.n407 10.4732
R624 VTAIL.n375 VTAIL.n288 10.4732
R625 VTAIL.n354 VTAIL.n299 10.4732
R626 VTAIL.n327 VTAIL.n311 10.4732
R627 VTAIL.n710 VTAIL.n709 9.69747
R628 VTAIL.n730 VTAIL.n729 9.69747
R629 VTAIL.n756 VTAIL.n666 9.69747
R630 VTAIL.n46 VTAIL.n45 9.69747
R631 VTAIL.n66 VTAIL.n65 9.69747
R632 VTAIL.n92 VTAIL.n2 9.69747
R633 VTAIL.n140 VTAIL.n139 9.69747
R634 VTAIL.n160 VTAIL.n159 9.69747
R635 VTAIL.n186 VTAIL.n96 9.69747
R636 VTAIL.n236 VTAIL.n235 9.69747
R637 VTAIL.n256 VTAIL.n255 9.69747
R638 VTAIL.n282 VTAIL.n192 9.69747
R639 VTAIL.n662 VTAIL.n572 9.69747
R640 VTAIL.n637 VTAIL.n636 9.69747
R641 VTAIL.n617 VTAIL.n616 9.69747
R642 VTAIL.n566 VTAIL.n476 9.69747
R643 VTAIL.n541 VTAIL.n540 9.69747
R644 VTAIL.n521 VTAIL.n520 9.69747
R645 VTAIL.n472 VTAIL.n382 9.69747
R646 VTAIL.n447 VTAIL.n446 9.69747
R647 VTAIL.n427 VTAIL.n426 9.69747
R648 VTAIL.n376 VTAIL.n286 9.69747
R649 VTAIL.n351 VTAIL.n350 9.69747
R650 VTAIL.n331 VTAIL.n330 9.69747
R651 VTAIL.n758 VTAIL.n757 9.45567
R652 VTAIL.n94 VTAIL.n93 9.45567
R653 VTAIL.n188 VTAIL.n187 9.45567
R654 VTAIL.n284 VTAIL.n283 9.45567
R655 VTAIL.n664 VTAIL.n663 9.45567
R656 VTAIL.n568 VTAIL.n567 9.45567
R657 VTAIL.n474 VTAIL.n473 9.45567
R658 VTAIL.n378 VTAIL.n377 9.45567
R659 VTAIL.n757 VTAIL.n756 9.3005
R660 VTAIL.n668 VTAIL.n667 9.3005
R661 VTAIL.n751 VTAIL.n750 9.3005
R662 VTAIL.n749 VTAIL.n748 9.3005
R663 VTAIL.n672 VTAIL.n671 9.3005
R664 VTAIL.n717 VTAIL.n716 9.3005
R665 VTAIL.n715 VTAIL.n714 9.3005
R666 VTAIL.n688 VTAIL.n687 9.3005
R667 VTAIL.n709 VTAIL.n708 9.3005
R668 VTAIL.n707 VTAIL.n706 9.3005
R669 VTAIL.n692 VTAIL.n691 9.3005
R670 VTAIL.n701 VTAIL.n700 9.3005
R671 VTAIL.n699 VTAIL.n698 9.3005
R672 VTAIL.n684 VTAIL.n683 9.3005
R673 VTAIL.n723 VTAIL.n722 9.3005
R674 VTAIL.n725 VTAIL.n724 9.3005
R675 VTAIL.n680 VTAIL.n679 9.3005
R676 VTAIL.n731 VTAIL.n730 9.3005
R677 VTAIL.n733 VTAIL.n732 9.3005
R678 VTAIL.n676 VTAIL.n675 9.3005
R679 VTAIL.n740 VTAIL.n739 9.3005
R680 VTAIL.n742 VTAIL.n741 9.3005
R681 VTAIL.n93 VTAIL.n92 9.3005
R682 VTAIL.n4 VTAIL.n3 9.3005
R683 VTAIL.n87 VTAIL.n86 9.3005
R684 VTAIL.n85 VTAIL.n84 9.3005
R685 VTAIL.n8 VTAIL.n7 9.3005
R686 VTAIL.n53 VTAIL.n52 9.3005
R687 VTAIL.n51 VTAIL.n50 9.3005
R688 VTAIL.n24 VTAIL.n23 9.3005
R689 VTAIL.n45 VTAIL.n44 9.3005
R690 VTAIL.n43 VTAIL.n42 9.3005
R691 VTAIL.n28 VTAIL.n27 9.3005
R692 VTAIL.n37 VTAIL.n36 9.3005
R693 VTAIL.n35 VTAIL.n34 9.3005
R694 VTAIL.n20 VTAIL.n19 9.3005
R695 VTAIL.n59 VTAIL.n58 9.3005
R696 VTAIL.n61 VTAIL.n60 9.3005
R697 VTAIL.n16 VTAIL.n15 9.3005
R698 VTAIL.n67 VTAIL.n66 9.3005
R699 VTAIL.n69 VTAIL.n68 9.3005
R700 VTAIL.n12 VTAIL.n11 9.3005
R701 VTAIL.n76 VTAIL.n75 9.3005
R702 VTAIL.n78 VTAIL.n77 9.3005
R703 VTAIL.n187 VTAIL.n186 9.3005
R704 VTAIL.n98 VTAIL.n97 9.3005
R705 VTAIL.n181 VTAIL.n180 9.3005
R706 VTAIL.n179 VTAIL.n178 9.3005
R707 VTAIL.n102 VTAIL.n101 9.3005
R708 VTAIL.n147 VTAIL.n146 9.3005
R709 VTAIL.n145 VTAIL.n144 9.3005
R710 VTAIL.n118 VTAIL.n117 9.3005
R711 VTAIL.n139 VTAIL.n138 9.3005
R712 VTAIL.n137 VTAIL.n136 9.3005
R713 VTAIL.n122 VTAIL.n121 9.3005
R714 VTAIL.n131 VTAIL.n130 9.3005
R715 VTAIL.n129 VTAIL.n128 9.3005
R716 VTAIL.n114 VTAIL.n113 9.3005
R717 VTAIL.n153 VTAIL.n152 9.3005
R718 VTAIL.n155 VTAIL.n154 9.3005
R719 VTAIL.n110 VTAIL.n109 9.3005
R720 VTAIL.n161 VTAIL.n160 9.3005
R721 VTAIL.n163 VTAIL.n162 9.3005
R722 VTAIL.n106 VTAIL.n105 9.3005
R723 VTAIL.n170 VTAIL.n169 9.3005
R724 VTAIL.n172 VTAIL.n171 9.3005
R725 VTAIL.n283 VTAIL.n282 9.3005
R726 VTAIL.n194 VTAIL.n193 9.3005
R727 VTAIL.n277 VTAIL.n276 9.3005
R728 VTAIL.n275 VTAIL.n274 9.3005
R729 VTAIL.n198 VTAIL.n197 9.3005
R730 VTAIL.n243 VTAIL.n242 9.3005
R731 VTAIL.n241 VTAIL.n240 9.3005
R732 VTAIL.n214 VTAIL.n213 9.3005
R733 VTAIL.n235 VTAIL.n234 9.3005
R734 VTAIL.n233 VTAIL.n232 9.3005
R735 VTAIL.n218 VTAIL.n217 9.3005
R736 VTAIL.n227 VTAIL.n226 9.3005
R737 VTAIL.n225 VTAIL.n224 9.3005
R738 VTAIL.n210 VTAIL.n209 9.3005
R739 VTAIL.n249 VTAIL.n248 9.3005
R740 VTAIL.n251 VTAIL.n250 9.3005
R741 VTAIL.n206 VTAIL.n205 9.3005
R742 VTAIL.n257 VTAIL.n256 9.3005
R743 VTAIL.n259 VTAIL.n258 9.3005
R744 VTAIL.n202 VTAIL.n201 9.3005
R745 VTAIL.n266 VTAIL.n265 9.3005
R746 VTAIL.n268 VTAIL.n267 9.3005
R747 VTAIL.n630 VTAIL.n629 9.3005
R748 VTAIL.n632 VTAIL.n631 9.3005
R749 VTAIL.n587 VTAIL.n586 9.3005
R750 VTAIL.n638 VTAIL.n637 9.3005
R751 VTAIL.n640 VTAIL.n639 9.3005
R752 VTAIL.n582 VTAIL.n581 9.3005
R753 VTAIL.n646 VTAIL.n645 9.3005
R754 VTAIL.n648 VTAIL.n647 9.3005
R755 VTAIL.n663 VTAIL.n662 9.3005
R756 VTAIL.n574 VTAIL.n573 9.3005
R757 VTAIL.n657 VTAIL.n656 9.3005
R758 VTAIL.n655 VTAIL.n654 9.3005
R759 VTAIL.n578 VTAIL.n577 9.3005
R760 VTAIL.n591 VTAIL.n590 9.3005
R761 VTAIL.n624 VTAIL.n623 9.3005
R762 VTAIL.n622 VTAIL.n621 9.3005
R763 VTAIL.n595 VTAIL.n594 9.3005
R764 VTAIL.n616 VTAIL.n615 9.3005
R765 VTAIL.n614 VTAIL.n613 9.3005
R766 VTAIL.n599 VTAIL.n598 9.3005
R767 VTAIL.n608 VTAIL.n607 9.3005
R768 VTAIL.n606 VTAIL.n605 9.3005
R769 VTAIL.n534 VTAIL.n533 9.3005
R770 VTAIL.n536 VTAIL.n535 9.3005
R771 VTAIL.n491 VTAIL.n490 9.3005
R772 VTAIL.n542 VTAIL.n541 9.3005
R773 VTAIL.n544 VTAIL.n543 9.3005
R774 VTAIL.n486 VTAIL.n485 9.3005
R775 VTAIL.n550 VTAIL.n549 9.3005
R776 VTAIL.n552 VTAIL.n551 9.3005
R777 VTAIL.n567 VTAIL.n566 9.3005
R778 VTAIL.n478 VTAIL.n477 9.3005
R779 VTAIL.n561 VTAIL.n560 9.3005
R780 VTAIL.n559 VTAIL.n558 9.3005
R781 VTAIL.n482 VTAIL.n481 9.3005
R782 VTAIL.n495 VTAIL.n494 9.3005
R783 VTAIL.n528 VTAIL.n527 9.3005
R784 VTAIL.n526 VTAIL.n525 9.3005
R785 VTAIL.n499 VTAIL.n498 9.3005
R786 VTAIL.n520 VTAIL.n519 9.3005
R787 VTAIL.n518 VTAIL.n517 9.3005
R788 VTAIL.n503 VTAIL.n502 9.3005
R789 VTAIL.n512 VTAIL.n511 9.3005
R790 VTAIL.n510 VTAIL.n509 9.3005
R791 VTAIL.n440 VTAIL.n439 9.3005
R792 VTAIL.n442 VTAIL.n441 9.3005
R793 VTAIL.n397 VTAIL.n396 9.3005
R794 VTAIL.n448 VTAIL.n447 9.3005
R795 VTAIL.n450 VTAIL.n449 9.3005
R796 VTAIL.n392 VTAIL.n391 9.3005
R797 VTAIL.n456 VTAIL.n455 9.3005
R798 VTAIL.n458 VTAIL.n457 9.3005
R799 VTAIL.n473 VTAIL.n472 9.3005
R800 VTAIL.n384 VTAIL.n383 9.3005
R801 VTAIL.n467 VTAIL.n466 9.3005
R802 VTAIL.n465 VTAIL.n464 9.3005
R803 VTAIL.n388 VTAIL.n387 9.3005
R804 VTAIL.n401 VTAIL.n400 9.3005
R805 VTAIL.n434 VTAIL.n433 9.3005
R806 VTAIL.n432 VTAIL.n431 9.3005
R807 VTAIL.n405 VTAIL.n404 9.3005
R808 VTAIL.n426 VTAIL.n425 9.3005
R809 VTAIL.n424 VTAIL.n423 9.3005
R810 VTAIL.n409 VTAIL.n408 9.3005
R811 VTAIL.n418 VTAIL.n417 9.3005
R812 VTAIL.n416 VTAIL.n415 9.3005
R813 VTAIL.n344 VTAIL.n343 9.3005
R814 VTAIL.n346 VTAIL.n345 9.3005
R815 VTAIL.n301 VTAIL.n300 9.3005
R816 VTAIL.n352 VTAIL.n351 9.3005
R817 VTAIL.n354 VTAIL.n353 9.3005
R818 VTAIL.n296 VTAIL.n295 9.3005
R819 VTAIL.n360 VTAIL.n359 9.3005
R820 VTAIL.n362 VTAIL.n361 9.3005
R821 VTAIL.n377 VTAIL.n376 9.3005
R822 VTAIL.n288 VTAIL.n287 9.3005
R823 VTAIL.n371 VTAIL.n370 9.3005
R824 VTAIL.n369 VTAIL.n368 9.3005
R825 VTAIL.n292 VTAIL.n291 9.3005
R826 VTAIL.n305 VTAIL.n304 9.3005
R827 VTAIL.n338 VTAIL.n337 9.3005
R828 VTAIL.n336 VTAIL.n335 9.3005
R829 VTAIL.n309 VTAIL.n308 9.3005
R830 VTAIL.n330 VTAIL.n329 9.3005
R831 VTAIL.n328 VTAIL.n327 9.3005
R832 VTAIL.n313 VTAIL.n312 9.3005
R833 VTAIL.n322 VTAIL.n321 9.3005
R834 VTAIL.n320 VTAIL.n319 9.3005
R835 VTAIL.n713 VTAIL.n688 8.92171
R836 VTAIL.n726 VTAIL.n680 8.92171
R837 VTAIL.n49 VTAIL.n24 8.92171
R838 VTAIL.n62 VTAIL.n16 8.92171
R839 VTAIL.n143 VTAIL.n118 8.92171
R840 VTAIL.n156 VTAIL.n110 8.92171
R841 VTAIL.n239 VTAIL.n214 8.92171
R842 VTAIL.n252 VTAIL.n206 8.92171
R843 VTAIL.n633 VTAIL.n587 8.92171
R844 VTAIL.n620 VTAIL.n595 8.92171
R845 VTAIL.n537 VTAIL.n491 8.92171
R846 VTAIL.n524 VTAIL.n499 8.92171
R847 VTAIL.n443 VTAIL.n397 8.92171
R848 VTAIL.n430 VTAIL.n405 8.92171
R849 VTAIL.n347 VTAIL.n301 8.92171
R850 VTAIL.n334 VTAIL.n309 8.92171
R851 VTAIL.n714 VTAIL.n686 8.14595
R852 VTAIL.n725 VTAIL.n682 8.14595
R853 VTAIL.n50 VTAIL.n22 8.14595
R854 VTAIL.n61 VTAIL.n18 8.14595
R855 VTAIL.n144 VTAIL.n116 8.14595
R856 VTAIL.n155 VTAIL.n112 8.14595
R857 VTAIL.n240 VTAIL.n212 8.14595
R858 VTAIL.n251 VTAIL.n208 8.14595
R859 VTAIL.n632 VTAIL.n589 8.14595
R860 VTAIL.n621 VTAIL.n593 8.14595
R861 VTAIL.n536 VTAIL.n493 8.14595
R862 VTAIL.n525 VTAIL.n497 8.14595
R863 VTAIL.n442 VTAIL.n399 8.14595
R864 VTAIL.n431 VTAIL.n403 8.14595
R865 VTAIL.n346 VTAIL.n303 8.14595
R866 VTAIL.n335 VTAIL.n307 8.14595
R867 VTAIL.n718 VTAIL.n717 7.3702
R868 VTAIL.n722 VTAIL.n721 7.3702
R869 VTAIL.n54 VTAIL.n53 7.3702
R870 VTAIL.n58 VTAIL.n57 7.3702
R871 VTAIL.n148 VTAIL.n147 7.3702
R872 VTAIL.n152 VTAIL.n151 7.3702
R873 VTAIL.n244 VTAIL.n243 7.3702
R874 VTAIL.n248 VTAIL.n247 7.3702
R875 VTAIL.n629 VTAIL.n628 7.3702
R876 VTAIL.n625 VTAIL.n624 7.3702
R877 VTAIL.n533 VTAIL.n532 7.3702
R878 VTAIL.n529 VTAIL.n528 7.3702
R879 VTAIL.n439 VTAIL.n438 7.3702
R880 VTAIL.n435 VTAIL.n434 7.3702
R881 VTAIL.n343 VTAIL.n342 7.3702
R882 VTAIL.n339 VTAIL.n338 7.3702
R883 VTAIL.n718 VTAIL.n684 6.59444
R884 VTAIL.n721 VTAIL.n684 6.59444
R885 VTAIL.n54 VTAIL.n20 6.59444
R886 VTAIL.n57 VTAIL.n20 6.59444
R887 VTAIL.n148 VTAIL.n114 6.59444
R888 VTAIL.n151 VTAIL.n114 6.59444
R889 VTAIL.n244 VTAIL.n210 6.59444
R890 VTAIL.n247 VTAIL.n210 6.59444
R891 VTAIL.n628 VTAIL.n591 6.59444
R892 VTAIL.n625 VTAIL.n591 6.59444
R893 VTAIL.n532 VTAIL.n495 6.59444
R894 VTAIL.n529 VTAIL.n495 6.59444
R895 VTAIL.n438 VTAIL.n401 6.59444
R896 VTAIL.n435 VTAIL.n401 6.59444
R897 VTAIL.n342 VTAIL.n305 6.59444
R898 VTAIL.n339 VTAIL.n305 6.59444
R899 VTAIL.n717 VTAIL.n686 5.81868
R900 VTAIL.n722 VTAIL.n682 5.81868
R901 VTAIL.n53 VTAIL.n22 5.81868
R902 VTAIL.n58 VTAIL.n18 5.81868
R903 VTAIL.n147 VTAIL.n116 5.81868
R904 VTAIL.n152 VTAIL.n112 5.81868
R905 VTAIL.n243 VTAIL.n212 5.81868
R906 VTAIL.n248 VTAIL.n208 5.81868
R907 VTAIL.n629 VTAIL.n589 5.81868
R908 VTAIL.n624 VTAIL.n593 5.81868
R909 VTAIL.n533 VTAIL.n493 5.81868
R910 VTAIL.n528 VTAIL.n497 5.81868
R911 VTAIL.n439 VTAIL.n399 5.81868
R912 VTAIL.n434 VTAIL.n403 5.81868
R913 VTAIL.n343 VTAIL.n303 5.81868
R914 VTAIL.n338 VTAIL.n307 5.81868
R915 VTAIL.n714 VTAIL.n713 5.04292
R916 VTAIL.n726 VTAIL.n725 5.04292
R917 VTAIL.n50 VTAIL.n49 5.04292
R918 VTAIL.n62 VTAIL.n61 5.04292
R919 VTAIL.n144 VTAIL.n143 5.04292
R920 VTAIL.n156 VTAIL.n155 5.04292
R921 VTAIL.n240 VTAIL.n239 5.04292
R922 VTAIL.n252 VTAIL.n251 5.04292
R923 VTAIL.n633 VTAIL.n632 5.04292
R924 VTAIL.n621 VTAIL.n620 5.04292
R925 VTAIL.n537 VTAIL.n536 5.04292
R926 VTAIL.n525 VTAIL.n524 5.04292
R927 VTAIL.n443 VTAIL.n442 5.04292
R928 VTAIL.n431 VTAIL.n430 5.04292
R929 VTAIL.n347 VTAIL.n346 5.04292
R930 VTAIL.n335 VTAIL.n334 5.04292
R931 VTAIL.n606 VTAIL.n602 4.38563
R932 VTAIL.n510 VTAIL.n506 4.38563
R933 VTAIL.n416 VTAIL.n412 4.38563
R934 VTAIL.n320 VTAIL.n316 4.38563
R935 VTAIL.n699 VTAIL.n695 4.38563
R936 VTAIL.n35 VTAIL.n31 4.38563
R937 VTAIL.n129 VTAIL.n125 4.38563
R938 VTAIL.n225 VTAIL.n221 4.38563
R939 VTAIL.n710 VTAIL.n688 4.26717
R940 VTAIL.n729 VTAIL.n680 4.26717
R941 VTAIL.n758 VTAIL.n666 4.26717
R942 VTAIL.n46 VTAIL.n24 4.26717
R943 VTAIL.n65 VTAIL.n16 4.26717
R944 VTAIL.n94 VTAIL.n2 4.26717
R945 VTAIL.n140 VTAIL.n118 4.26717
R946 VTAIL.n159 VTAIL.n110 4.26717
R947 VTAIL.n188 VTAIL.n96 4.26717
R948 VTAIL.n236 VTAIL.n214 4.26717
R949 VTAIL.n255 VTAIL.n206 4.26717
R950 VTAIL.n284 VTAIL.n192 4.26717
R951 VTAIL.n664 VTAIL.n572 4.26717
R952 VTAIL.n636 VTAIL.n587 4.26717
R953 VTAIL.n617 VTAIL.n595 4.26717
R954 VTAIL.n568 VTAIL.n476 4.26717
R955 VTAIL.n540 VTAIL.n491 4.26717
R956 VTAIL.n521 VTAIL.n499 4.26717
R957 VTAIL.n474 VTAIL.n382 4.26717
R958 VTAIL.n446 VTAIL.n397 4.26717
R959 VTAIL.n427 VTAIL.n405 4.26717
R960 VTAIL.n378 VTAIL.n286 4.26717
R961 VTAIL.n350 VTAIL.n301 4.26717
R962 VTAIL.n331 VTAIL.n309 4.26717
R963 VTAIL.n709 VTAIL.n690 3.49141
R964 VTAIL.n730 VTAIL.n678 3.49141
R965 VTAIL.n756 VTAIL.n755 3.49141
R966 VTAIL.n45 VTAIL.n26 3.49141
R967 VTAIL.n66 VTAIL.n14 3.49141
R968 VTAIL.n92 VTAIL.n91 3.49141
R969 VTAIL.n139 VTAIL.n120 3.49141
R970 VTAIL.n160 VTAIL.n108 3.49141
R971 VTAIL.n186 VTAIL.n185 3.49141
R972 VTAIL.n235 VTAIL.n216 3.49141
R973 VTAIL.n256 VTAIL.n204 3.49141
R974 VTAIL.n282 VTAIL.n281 3.49141
R975 VTAIL.n662 VTAIL.n661 3.49141
R976 VTAIL.n637 VTAIL.n585 3.49141
R977 VTAIL.n616 VTAIL.n597 3.49141
R978 VTAIL.n566 VTAIL.n565 3.49141
R979 VTAIL.n541 VTAIL.n489 3.49141
R980 VTAIL.n520 VTAIL.n501 3.49141
R981 VTAIL.n472 VTAIL.n471 3.49141
R982 VTAIL.n447 VTAIL.n395 3.49141
R983 VTAIL.n426 VTAIL.n407 3.49141
R984 VTAIL.n376 VTAIL.n375 3.49141
R985 VTAIL.n351 VTAIL.n299 3.49141
R986 VTAIL.n330 VTAIL.n311 3.49141
R987 VTAIL.n706 VTAIL.n705 2.71565
R988 VTAIL.n734 VTAIL.n733 2.71565
R989 VTAIL.n752 VTAIL.n668 2.71565
R990 VTAIL.n42 VTAIL.n41 2.71565
R991 VTAIL.n70 VTAIL.n69 2.71565
R992 VTAIL.n88 VTAIL.n4 2.71565
R993 VTAIL.n136 VTAIL.n135 2.71565
R994 VTAIL.n164 VTAIL.n163 2.71565
R995 VTAIL.n182 VTAIL.n98 2.71565
R996 VTAIL.n232 VTAIL.n231 2.71565
R997 VTAIL.n260 VTAIL.n259 2.71565
R998 VTAIL.n278 VTAIL.n194 2.71565
R999 VTAIL.n658 VTAIL.n574 2.71565
R1000 VTAIL.n641 VTAIL.n640 2.71565
R1001 VTAIL.n613 VTAIL.n612 2.71565
R1002 VTAIL.n562 VTAIL.n478 2.71565
R1003 VTAIL.n545 VTAIL.n544 2.71565
R1004 VTAIL.n517 VTAIL.n516 2.71565
R1005 VTAIL.n468 VTAIL.n384 2.71565
R1006 VTAIL.n451 VTAIL.n450 2.71565
R1007 VTAIL.n423 VTAIL.n422 2.71565
R1008 VTAIL.n372 VTAIL.n288 2.71565
R1009 VTAIL.n355 VTAIL.n354 2.71565
R1010 VTAIL.n327 VTAIL.n326 2.71565
R1011 VTAIL.n381 VTAIL.n379 2.68153
R1012 VTAIL.n475 VTAIL.n381 2.68153
R1013 VTAIL.n571 VTAIL.n569 2.68153
R1014 VTAIL.n665 VTAIL.n571 2.68153
R1015 VTAIL.n285 VTAIL.n191 2.68153
R1016 VTAIL.n191 VTAIL.n189 2.68153
R1017 VTAIL.n95 VTAIL.n1 2.68153
R1018 VTAIL VTAIL.n759 2.62334
R1019 VTAIL.n702 VTAIL.n692 1.93989
R1020 VTAIL.n738 VTAIL.n676 1.93989
R1021 VTAIL.n751 VTAIL.n670 1.93989
R1022 VTAIL.n38 VTAIL.n28 1.93989
R1023 VTAIL.n74 VTAIL.n12 1.93989
R1024 VTAIL.n87 VTAIL.n6 1.93989
R1025 VTAIL.n132 VTAIL.n122 1.93989
R1026 VTAIL.n168 VTAIL.n106 1.93989
R1027 VTAIL.n181 VTAIL.n100 1.93989
R1028 VTAIL.n228 VTAIL.n218 1.93989
R1029 VTAIL.n264 VTAIL.n202 1.93989
R1030 VTAIL.n277 VTAIL.n196 1.93989
R1031 VTAIL.n657 VTAIL.n576 1.93989
R1032 VTAIL.n644 VTAIL.n582 1.93989
R1033 VTAIL.n609 VTAIL.n599 1.93989
R1034 VTAIL.n561 VTAIL.n480 1.93989
R1035 VTAIL.n548 VTAIL.n486 1.93989
R1036 VTAIL.n513 VTAIL.n503 1.93989
R1037 VTAIL.n467 VTAIL.n386 1.93989
R1038 VTAIL.n454 VTAIL.n392 1.93989
R1039 VTAIL.n419 VTAIL.n409 1.93989
R1040 VTAIL.n371 VTAIL.n290 1.93989
R1041 VTAIL.n358 VTAIL.n296 1.93989
R1042 VTAIL.n323 VTAIL.n313 1.93989
R1043 VTAIL.n0 VTAIL.t6 1.16658
R1044 VTAIL.n0 VTAIL.t0 1.16658
R1045 VTAIL.n190 VTAIL.t9 1.16658
R1046 VTAIL.n190 VTAIL.t13 1.16658
R1047 VTAIL.n570 VTAIL.t11 1.16658
R1048 VTAIL.n570 VTAIL.t8 1.16658
R1049 VTAIL.n380 VTAIL.t1 1.16658
R1050 VTAIL.n380 VTAIL.t3 1.16658
R1051 VTAIL.n701 VTAIL.n694 1.16414
R1052 VTAIL.n739 VTAIL.n674 1.16414
R1053 VTAIL.n748 VTAIL.n747 1.16414
R1054 VTAIL.n37 VTAIL.n30 1.16414
R1055 VTAIL.n75 VTAIL.n10 1.16414
R1056 VTAIL.n84 VTAIL.n83 1.16414
R1057 VTAIL.n131 VTAIL.n124 1.16414
R1058 VTAIL.n169 VTAIL.n104 1.16414
R1059 VTAIL.n178 VTAIL.n177 1.16414
R1060 VTAIL.n227 VTAIL.n220 1.16414
R1061 VTAIL.n265 VTAIL.n200 1.16414
R1062 VTAIL.n274 VTAIL.n273 1.16414
R1063 VTAIL.n654 VTAIL.n653 1.16414
R1064 VTAIL.n645 VTAIL.n580 1.16414
R1065 VTAIL.n608 VTAIL.n601 1.16414
R1066 VTAIL.n558 VTAIL.n557 1.16414
R1067 VTAIL.n549 VTAIL.n484 1.16414
R1068 VTAIL.n512 VTAIL.n505 1.16414
R1069 VTAIL.n464 VTAIL.n463 1.16414
R1070 VTAIL.n455 VTAIL.n390 1.16414
R1071 VTAIL.n418 VTAIL.n411 1.16414
R1072 VTAIL.n368 VTAIL.n367 1.16414
R1073 VTAIL.n359 VTAIL.n294 1.16414
R1074 VTAIL.n322 VTAIL.n315 1.16414
R1075 VTAIL.n569 VTAIL.n475 0.470328
R1076 VTAIL.n189 VTAIL.n95 0.470328
R1077 VTAIL.n698 VTAIL.n697 0.388379
R1078 VTAIL.n743 VTAIL.n742 0.388379
R1079 VTAIL.n744 VTAIL.n672 0.388379
R1080 VTAIL.n34 VTAIL.n33 0.388379
R1081 VTAIL.n79 VTAIL.n78 0.388379
R1082 VTAIL.n80 VTAIL.n8 0.388379
R1083 VTAIL.n128 VTAIL.n127 0.388379
R1084 VTAIL.n173 VTAIL.n172 0.388379
R1085 VTAIL.n174 VTAIL.n102 0.388379
R1086 VTAIL.n224 VTAIL.n223 0.388379
R1087 VTAIL.n269 VTAIL.n268 0.388379
R1088 VTAIL.n270 VTAIL.n198 0.388379
R1089 VTAIL.n650 VTAIL.n578 0.388379
R1090 VTAIL.n649 VTAIL.n648 0.388379
R1091 VTAIL.n605 VTAIL.n604 0.388379
R1092 VTAIL.n554 VTAIL.n482 0.388379
R1093 VTAIL.n553 VTAIL.n552 0.388379
R1094 VTAIL.n509 VTAIL.n508 0.388379
R1095 VTAIL.n460 VTAIL.n388 0.388379
R1096 VTAIL.n459 VTAIL.n458 0.388379
R1097 VTAIL.n415 VTAIL.n414 0.388379
R1098 VTAIL.n364 VTAIL.n292 0.388379
R1099 VTAIL.n363 VTAIL.n362 0.388379
R1100 VTAIL.n319 VTAIL.n318 0.388379
R1101 VTAIL.n700 VTAIL.n699 0.155672
R1102 VTAIL.n700 VTAIL.n691 0.155672
R1103 VTAIL.n707 VTAIL.n691 0.155672
R1104 VTAIL.n708 VTAIL.n707 0.155672
R1105 VTAIL.n708 VTAIL.n687 0.155672
R1106 VTAIL.n715 VTAIL.n687 0.155672
R1107 VTAIL.n716 VTAIL.n715 0.155672
R1108 VTAIL.n716 VTAIL.n683 0.155672
R1109 VTAIL.n723 VTAIL.n683 0.155672
R1110 VTAIL.n724 VTAIL.n723 0.155672
R1111 VTAIL.n724 VTAIL.n679 0.155672
R1112 VTAIL.n731 VTAIL.n679 0.155672
R1113 VTAIL.n732 VTAIL.n731 0.155672
R1114 VTAIL.n732 VTAIL.n675 0.155672
R1115 VTAIL.n740 VTAIL.n675 0.155672
R1116 VTAIL.n741 VTAIL.n740 0.155672
R1117 VTAIL.n741 VTAIL.n671 0.155672
R1118 VTAIL.n749 VTAIL.n671 0.155672
R1119 VTAIL.n750 VTAIL.n749 0.155672
R1120 VTAIL.n750 VTAIL.n667 0.155672
R1121 VTAIL.n757 VTAIL.n667 0.155672
R1122 VTAIL.n36 VTAIL.n35 0.155672
R1123 VTAIL.n36 VTAIL.n27 0.155672
R1124 VTAIL.n43 VTAIL.n27 0.155672
R1125 VTAIL.n44 VTAIL.n43 0.155672
R1126 VTAIL.n44 VTAIL.n23 0.155672
R1127 VTAIL.n51 VTAIL.n23 0.155672
R1128 VTAIL.n52 VTAIL.n51 0.155672
R1129 VTAIL.n52 VTAIL.n19 0.155672
R1130 VTAIL.n59 VTAIL.n19 0.155672
R1131 VTAIL.n60 VTAIL.n59 0.155672
R1132 VTAIL.n60 VTAIL.n15 0.155672
R1133 VTAIL.n67 VTAIL.n15 0.155672
R1134 VTAIL.n68 VTAIL.n67 0.155672
R1135 VTAIL.n68 VTAIL.n11 0.155672
R1136 VTAIL.n76 VTAIL.n11 0.155672
R1137 VTAIL.n77 VTAIL.n76 0.155672
R1138 VTAIL.n77 VTAIL.n7 0.155672
R1139 VTAIL.n85 VTAIL.n7 0.155672
R1140 VTAIL.n86 VTAIL.n85 0.155672
R1141 VTAIL.n86 VTAIL.n3 0.155672
R1142 VTAIL.n93 VTAIL.n3 0.155672
R1143 VTAIL.n130 VTAIL.n129 0.155672
R1144 VTAIL.n130 VTAIL.n121 0.155672
R1145 VTAIL.n137 VTAIL.n121 0.155672
R1146 VTAIL.n138 VTAIL.n137 0.155672
R1147 VTAIL.n138 VTAIL.n117 0.155672
R1148 VTAIL.n145 VTAIL.n117 0.155672
R1149 VTAIL.n146 VTAIL.n145 0.155672
R1150 VTAIL.n146 VTAIL.n113 0.155672
R1151 VTAIL.n153 VTAIL.n113 0.155672
R1152 VTAIL.n154 VTAIL.n153 0.155672
R1153 VTAIL.n154 VTAIL.n109 0.155672
R1154 VTAIL.n161 VTAIL.n109 0.155672
R1155 VTAIL.n162 VTAIL.n161 0.155672
R1156 VTAIL.n162 VTAIL.n105 0.155672
R1157 VTAIL.n170 VTAIL.n105 0.155672
R1158 VTAIL.n171 VTAIL.n170 0.155672
R1159 VTAIL.n171 VTAIL.n101 0.155672
R1160 VTAIL.n179 VTAIL.n101 0.155672
R1161 VTAIL.n180 VTAIL.n179 0.155672
R1162 VTAIL.n180 VTAIL.n97 0.155672
R1163 VTAIL.n187 VTAIL.n97 0.155672
R1164 VTAIL.n226 VTAIL.n225 0.155672
R1165 VTAIL.n226 VTAIL.n217 0.155672
R1166 VTAIL.n233 VTAIL.n217 0.155672
R1167 VTAIL.n234 VTAIL.n233 0.155672
R1168 VTAIL.n234 VTAIL.n213 0.155672
R1169 VTAIL.n241 VTAIL.n213 0.155672
R1170 VTAIL.n242 VTAIL.n241 0.155672
R1171 VTAIL.n242 VTAIL.n209 0.155672
R1172 VTAIL.n249 VTAIL.n209 0.155672
R1173 VTAIL.n250 VTAIL.n249 0.155672
R1174 VTAIL.n250 VTAIL.n205 0.155672
R1175 VTAIL.n257 VTAIL.n205 0.155672
R1176 VTAIL.n258 VTAIL.n257 0.155672
R1177 VTAIL.n258 VTAIL.n201 0.155672
R1178 VTAIL.n266 VTAIL.n201 0.155672
R1179 VTAIL.n267 VTAIL.n266 0.155672
R1180 VTAIL.n267 VTAIL.n197 0.155672
R1181 VTAIL.n275 VTAIL.n197 0.155672
R1182 VTAIL.n276 VTAIL.n275 0.155672
R1183 VTAIL.n276 VTAIL.n193 0.155672
R1184 VTAIL.n283 VTAIL.n193 0.155672
R1185 VTAIL.n663 VTAIL.n573 0.155672
R1186 VTAIL.n656 VTAIL.n573 0.155672
R1187 VTAIL.n656 VTAIL.n655 0.155672
R1188 VTAIL.n655 VTAIL.n577 0.155672
R1189 VTAIL.n647 VTAIL.n577 0.155672
R1190 VTAIL.n647 VTAIL.n646 0.155672
R1191 VTAIL.n646 VTAIL.n581 0.155672
R1192 VTAIL.n639 VTAIL.n581 0.155672
R1193 VTAIL.n639 VTAIL.n638 0.155672
R1194 VTAIL.n638 VTAIL.n586 0.155672
R1195 VTAIL.n631 VTAIL.n586 0.155672
R1196 VTAIL.n631 VTAIL.n630 0.155672
R1197 VTAIL.n630 VTAIL.n590 0.155672
R1198 VTAIL.n623 VTAIL.n590 0.155672
R1199 VTAIL.n623 VTAIL.n622 0.155672
R1200 VTAIL.n622 VTAIL.n594 0.155672
R1201 VTAIL.n615 VTAIL.n594 0.155672
R1202 VTAIL.n615 VTAIL.n614 0.155672
R1203 VTAIL.n614 VTAIL.n598 0.155672
R1204 VTAIL.n607 VTAIL.n598 0.155672
R1205 VTAIL.n607 VTAIL.n606 0.155672
R1206 VTAIL.n567 VTAIL.n477 0.155672
R1207 VTAIL.n560 VTAIL.n477 0.155672
R1208 VTAIL.n560 VTAIL.n559 0.155672
R1209 VTAIL.n559 VTAIL.n481 0.155672
R1210 VTAIL.n551 VTAIL.n481 0.155672
R1211 VTAIL.n551 VTAIL.n550 0.155672
R1212 VTAIL.n550 VTAIL.n485 0.155672
R1213 VTAIL.n543 VTAIL.n485 0.155672
R1214 VTAIL.n543 VTAIL.n542 0.155672
R1215 VTAIL.n542 VTAIL.n490 0.155672
R1216 VTAIL.n535 VTAIL.n490 0.155672
R1217 VTAIL.n535 VTAIL.n534 0.155672
R1218 VTAIL.n534 VTAIL.n494 0.155672
R1219 VTAIL.n527 VTAIL.n494 0.155672
R1220 VTAIL.n527 VTAIL.n526 0.155672
R1221 VTAIL.n526 VTAIL.n498 0.155672
R1222 VTAIL.n519 VTAIL.n498 0.155672
R1223 VTAIL.n519 VTAIL.n518 0.155672
R1224 VTAIL.n518 VTAIL.n502 0.155672
R1225 VTAIL.n511 VTAIL.n502 0.155672
R1226 VTAIL.n511 VTAIL.n510 0.155672
R1227 VTAIL.n473 VTAIL.n383 0.155672
R1228 VTAIL.n466 VTAIL.n383 0.155672
R1229 VTAIL.n466 VTAIL.n465 0.155672
R1230 VTAIL.n465 VTAIL.n387 0.155672
R1231 VTAIL.n457 VTAIL.n387 0.155672
R1232 VTAIL.n457 VTAIL.n456 0.155672
R1233 VTAIL.n456 VTAIL.n391 0.155672
R1234 VTAIL.n449 VTAIL.n391 0.155672
R1235 VTAIL.n449 VTAIL.n448 0.155672
R1236 VTAIL.n448 VTAIL.n396 0.155672
R1237 VTAIL.n441 VTAIL.n396 0.155672
R1238 VTAIL.n441 VTAIL.n440 0.155672
R1239 VTAIL.n440 VTAIL.n400 0.155672
R1240 VTAIL.n433 VTAIL.n400 0.155672
R1241 VTAIL.n433 VTAIL.n432 0.155672
R1242 VTAIL.n432 VTAIL.n404 0.155672
R1243 VTAIL.n425 VTAIL.n404 0.155672
R1244 VTAIL.n425 VTAIL.n424 0.155672
R1245 VTAIL.n424 VTAIL.n408 0.155672
R1246 VTAIL.n417 VTAIL.n408 0.155672
R1247 VTAIL.n417 VTAIL.n416 0.155672
R1248 VTAIL.n377 VTAIL.n287 0.155672
R1249 VTAIL.n370 VTAIL.n287 0.155672
R1250 VTAIL.n370 VTAIL.n369 0.155672
R1251 VTAIL.n369 VTAIL.n291 0.155672
R1252 VTAIL.n361 VTAIL.n291 0.155672
R1253 VTAIL.n361 VTAIL.n360 0.155672
R1254 VTAIL.n360 VTAIL.n295 0.155672
R1255 VTAIL.n353 VTAIL.n295 0.155672
R1256 VTAIL.n353 VTAIL.n352 0.155672
R1257 VTAIL.n352 VTAIL.n300 0.155672
R1258 VTAIL.n345 VTAIL.n300 0.155672
R1259 VTAIL.n345 VTAIL.n344 0.155672
R1260 VTAIL.n344 VTAIL.n304 0.155672
R1261 VTAIL.n337 VTAIL.n304 0.155672
R1262 VTAIL.n337 VTAIL.n336 0.155672
R1263 VTAIL.n336 VTAIL.n308 0.155672
R1264 VTAIL.n329 VTAIL.n308 0.155672
R1265 VTAIL.n329 VTAIL.n328 0.155672
R1266 VTAIL.n328 VTAIL.n312 0.155672
R1267 VTAIL.n321 VTAIL.n312 0.155672
R1268 VTAIL.n321 VTAIL.n320 0.155672
R1269 VTAIL VTAIL.n1 0.0586897
R1270 VDD1 VDD1.n0 65.6144
R1271 VDD1.n3 VDD1.n2 65.5007
R1272 VDD1.n3 VDD1.n1 65.5007
R1273 VDD1.n5 VDD1.n4 64.2155
R1274 VDD1.n5 VDD1.n3 51.0009
R1275 VDD1 VDD1.n5 1.28283
R1276 VDD1.n4 VDD1.t6 1.16658
R1277 VDD1.n4 VDD1.t0 1.16658
R1278 VDD1.n0 VDD1.t2 1.16658
R1279 VDD1.n0 VDD1.t5 1.16658
R1280 VDD1.n2 VDD1.t1 1.16658
R1281 VDD1.n2 VDD1.t4 1.16658
R1282 VDD1.n1 VDD1.t3 1.16658
R1283 VDD1.n1 VDD1.t7 1.16658
R1284 B.n813 B.n812 585
R1285 B.n815 B.n165 585
R1286 B.n818 B.n817 585
R1287 B.n819 B.n164 585
R1288 B.n821 B.n820 585
R1289 B.n823 B.n163 585
R1290 B.n826 B.n825 585
R1291 B.n827 B.n162 585
R1292 B.n829 B.n828 585
R1293 B.n831 B.n161 585
R1294 B.n834 B.n833 585
R1295 B.n835 B.n160 585
R1296 B.n837 B.n836 585
R1297 B.n839 B.n159 585
R1298 B.n842 B.n841 585
R1299 B.n843 B.n158 585
R1300 B.n845 B.n844 585
R1301 B.n847 B.n157 585
R1302 B.n850 B.n849 585
R1303 B.n851 B.n156 585
R1304 B.n853 B.n852 585
R1305 B.n855 B.n155 585
R1306 B.n858 B.n857 585
R1307 B.n859 B.n154 585
R1308 B.n861 B.n860 585
R1309 B.n863 B.n153 585
R1310 B.n866 B.n865 585
R1311 B.n867 B.n152 585
R1312 B.n869 B.n868 585
R1313 B.n871 B.n151 585
R1314 B.n874 B.n873 585
R1315 B.n875 B.n150 585
R1316 B.n877 B.n876 585
R1317 B.n879 B.n149 585
R1318 B.n882 B.n881 585
R1319 B.n883 B.n148 585
R1320 B.n885 B.n884 585
R1321 B.n887 B.n147 585
R1322 B.n890 B.n889 585
R1323 B.n891 B.n146 585
R1324 B.n893 B.n892 585
R1325 B.n895 B.n145 585
R1326 B.n898 B.n897 585
R1327 B.n899 B.n144 585
R1328 B.n901 B.n900 585
R1329 B.n903 B.n143 585
R1330 B.n906 B.n905 585
R1331 B.n907 B.n142 585
R1332 B.n909 B.n908 585
R1333 B.n911 B.n141 585
R1334 B.n914 B.n913 585
R1335 B.n915 B.n140 585
R1336 B.n917 B.n916 585
R1337 B.n919 B.n139 585
R1338 B.n921 B.n920 585
R1339 B.n923 B.n922 585
R1340 B.n926 B.n925 585
R1341 B.n927 B.n134 585
R1342 B.n929 B.n928 585
R1343 B.n931 B.n133 585
R1344 B.n934 B.n933 585
R1345 B.n935 B.n132 585
R1346 B.n937 B.n936 585
R1347 B.n939 B.n131 585
R1348 B.n942 B.n941 585
R1349 B.n943 B.n128 585
R1350 B.n946 B.n945 585
R1351 B.n948 B.n127 585
R1352 B.n951 B.n950 585
R1353 B.n952 B.n126 585
R1354 B.n954 B.n953 585
R1355 B.n956 B.n125 585
R1356 B.n959 B.n958 585
R1357 B.n960 B.n124 585
R1358 B.n962 B.n961 585
R1359 B.n964 B.n123 585
R1360 B.n967 B.n966 585
R1361 B.n968 B.n122 585
R1362 B.n970 B.n969 585
R1363 B.n972 B.n121 585
R1364 B.n975 B.n974 585
R1365 B.n976 B.n120 585
R1366 B.n978 B.n977 585
R1367 B.n980 B.n119 585
R1368 B.n983 B.n982 585
R1369 B.n984 B.n118 585
R1370 B.n986 B.n985 585
R1371 B.n988 B.n117 585
R1372 B.n991 B.n990 585
R1373 B.n992 B.n116 585
R1374 B.n994 B.n993 585
R1375 B.n996 B.n115 585
R1376 B.n999 B.n998 585
R1377 B.n1000 B.n114 585
R1378 B.n1002 B.n1001 585
R1379 B.n1004 B.n113 585
R1380 B.n1007 B.n1006 585
R1381 B.n1008 B.n112 585
R1382 B.n1010 B.n1009 585
R1383 B.n1012 B.n111 585
R1384 B.n1015 B.n1014 585
R1385 B.n1016 B.n110 585
R1386 B.n1018 B.n1017 585
R1387 B.n1020 B.n109 585
R1388 B.n1023 B.n1022 585
R1389 B.n1024 B.n108 585
R1390 B.n1026 B.n1025 585
R1391 B.n1028 B.n107 585
R1392 B.n1031 B.n1030 585
R1393 B.n1032 B.n106 585
R1394 B.n1034 B.n1033 585
R1395 B.n1036 B.n105 585
R1396 B.n1039 B.n1038 585
R1397 B.n1040 B.n104 585
R1398 B.n1042 B.n1041 585
R1399 B.n1044 B.n103 585
R1400 B.n1047 B.n1046 585
R1401 B.n1048 B.n102 585
R1402 B.n1050 B.n1049 585
R1403 B.n1052 B.n101 585
R1404 B.n1055 B.n1054 585
R1405 B.n1056 B.n100 585
R1406 B.n811 B.n98 585
R1407 B.n1059 B.n98 585
R1408 B.n810 B.n97 585
R1409 B.n1060 B.n97 585
R1410 B.n809 B.n96 585
R1411 B.n1061 B.n96 585
R1412 B.n808 B.n807 585
R1413 B.n807 B.n92 585
R1414 B.n806 B.n91 585
R1415 B.n1067 B.n91 585
R1416 B.n805 B.n90 585
R1417 B.n1068 B.n90 585
R1418 B.n804 B.n89 585
R1419 B.n1069 B.n89 585
R1420 B.n803 B.n802 585
R1421 B.n802 B.n85 585
R1422 B.n801 B.n84 585
R1423 B.n1075 B.n84 585
R1424 B.n800 B.n83 585
R1425 B.n1076 B.n83 585
R1426 B.n799 B.n82 585
R1427 B.n1077 B.n82 585
R1428 B.n798 B.n797 585
R1429 B.n797 B.n78 585
R1430 B.n796 B.n77 585
R1431 B.n1083 B.n77 585
R1432 B.n795 B.n76 585
R1433 B.n1084 B.n76 585
R1434 B.n794 B.n75 585
R1435 B.n1085 B.n75 585
R1436 B.n793 B.n792 585
R1437 B.n792 B.n71 585
R1438 B.n791 B.n70 585
R1439 B.n1091 B.n70 585
R1440 B.n790 B.n69 585
R1441 B.n1092 B.n69 585
R1442 B.n789 B.n68 585
R1443 B.n1093 B.n68 585
R1444 B.n788 B.n787 585
R1445 B.n787 B.n64 585
R1446 B.n786 B.n63 585
R1447 B.n1099 B.n63 585
R1448 B.n785 B.n62 585
R1449 B.n1100 B.n62 585
R1450 B.n784 B.n61 585
R1451 B.n1101 B.n61 585
R1452 B.n783 B.n782 585
R1453 B.n782 B.n57 585
R1454 B.n781 B.n56 585
R1455 B.n1107 B.n56 585
R1456 B.n780 B.n55 585
R1457 B.n1108 B.n55 585
R1458 B.n779 B.n54 585
R1459 B.n1109 B.n54 585
R1460 B.n778 B.n777 585
R1461 B.n777 B.n50 585
R1462 B.n776 B.n49 585
R1463 B.n1115 B.n49 585
R1464 B.n775 B.n48 585
R1465 B.n1116 B.n48 585
R1466 B.n774 B.n47 585
R1467 B.n1117 B.n47 585
R1468 B.n773 B.n772 585
R1469 B.n772 B.n43 585
R1470 B.n771 B.n42 585
R1471 B.n1123 B.n42 585
R1472 B.n770 B.n41 585
R1473 B.n1124 B.n41 585
R1474 B.n769 B.n40 585
R1475 B.n1125 B.n40 585
R1476 B.n768 B.n767 585
R1477 B.n767 B.n36 585
R1478 B.n766 B.n35 585
R1479 B.n1131 B.n35 585
R1480 B.n765 B.n34 585
R1481 B.n1132 B.n34 585
R1482 B.n764 B.n33 585
R1483 B.n1133 B.n33 585
R1484 B.n763 B.n762 585
R1485 B.n762 B.n29 585
R1486 B.n761 B.n28 585
R1487 B.n1139 B.n28 585
R1488 B.n760 B.n27 585
R1489 B.n1140 B.n27 585
R1490 B.n759 B.n26 585
R1491 B.n1141 B.n26 585
R1492 B.n758 B.n757 585
R1493 B.n757 B.n22 585
R1494 B.n756 B.n21 585
R1495 B.n1147 B.n21 585
R1496 B.n755 B.n20 585
R1497 B.n1148 B.n20 585
R1498 B.n754 B.n19 585
R1499 B.n1149 B.n19 585
R1500 B.n753 B.n752 585
R1501 B.n752 B.n18 585
R1502 B.n751 B.n14 585
R1503 B.n1155 B.n14 585
R1504 B.n750 B.n13 585
R1505 B.n1156 B.n13 585
R1506 B.n749 B.n12 585
R1507 B.n1157 B.n12 585
R1508 B.n748 B.n747 585
R1509 B.n747 B.n8 585
R1510 B.n746 B.n7 585
R1511 B.n1163 B.n7 585
R1512 B.n745 B.n6 585
R1513 B.n1164 B.n6 585
R1514 B.n744 B.n5 585
R1515 B.n1165 B.n5 585
R1516 B.n743 B.n742 585
R1517 B.n742 B.n4 585
R1518 B.n741 B.n166 585
R1519 B.n741 B.n740 585
R1520 B.n731 B.n167 585
R1521 B.n168 B.n167 585
R1522 B.n733 B.n732 585
R1523 B.n734 B.n733 585
R1524 B.n730 B.n173 585
R1525 B.n173 B.n172 585
R1526 B.n729 B.n728 585
R1527 B.n728 B.n727 585
R1528 B.n175 B.n174 585
R1529 B.n720 B.n175 585
R1530 B.n719 B.n718 585
R1531 B.n721 B.n719 585
R1532 B.n717 B.n180 585
R1533 B.n180 B.n179 585
R1534 B.n716 B.n715 585
R1535 B.n715 B.n714 585
R1536 B.n182 B.n181 585
R1537 B.n183 B.n182 585
R1538 B.n707 B.n706 585
R1539 B.n708 B.n707 585
R1540 B.n705 B.n188 585
R1541 B.n188 B.n187 585
R1542 B.n704 B.n703 585
R1543 B.n703 B.n702 585
R1544 B.n190 B.n189 585
R1545 B.n191 B.n190 585
R1546 B.n695 B.n694 585
R1547 B.n696 B.n695 585
R1548 B.n693 B.n196 585
R1549 B.n196 B.n195 585
R1550 B.n692 B.n691 585
R1551 B.n691 B.n690 585
R1552 B.n198 B.n197 585
R1553 B.n199 B.n198 585
R1554 B.n683 B.n682 585
R1555 B.n684 B.n683 585
R1556 B.n681 B.n204 585
R1557 B.n204 B.n203 585
R1558 B.n680 B.n679 585
R1559 B.n679 B.n678 585
R1560 B.n206 B.n205 585
R1561 B.n207 B.n206 585
R1562 B.n671 B.n670 585
R1563 B.n672 B.n671 585
R1564 B.n669 B.n211 585
R1565 B.n215 B.n211 585
R1566 B.n668 B.n667 585
R1567 B.n667 B.n666 585
R1568 B.n213 B.n212 585
R1569 B.n214 B.n213 585
R1570 B.n659 B.n658 585
R1571 B.n660 B.n659 585
R1572 B.n657 B.n220 585
R1573 B.n220 B.n219 585
R1574 B.n656 B.n655 585
R1575 B.n655 B.n654 585
R1576 B.n222 B.n221 585
R1577 B.n223 B.n222 585
R1578 B.n647 B.n646 585
R1579 B.n648 B.n647 585
R1580 B.n645 B.n228 585
R1581 B.n228 B.n227 585
R1582 B.n644 B.n643 585
R1583 B.n643 B.n642 585
R1584 B.n230 B.n229 585
R1585 B.n231 B.n230 585
R1586 B.n635 B.n634 585
R1587 B.n636 B.n635 585
R1588 B.n633 B.n236 585
R1589 B.n236 B.n235 585
R1590 B.n632 B.n631 585
R1591 B.n631 B.n630 585
R1592 B.n238 B.n237 585
R1593 B.n239 B.n238 585
R1594 B.n623 B.n622 585
R1595 B.n624 B.n623 585
R1596 B.n621 B.n244 585
R1597 B.n244 B.n243 585
R1598 B.n620 B.n619 585
R1599 B.n619 B.n618 585
R1600 B.n246 B.n245 585
R1601 B.n247 B.n246 585
R1602 B.n611 B.n610 585
R1603 B.n612 B.n611 585
R1604 B.n609 B.n252 585
R1605 B.n252 B.n251 585
R1606 B.n608 B.n607 585
R1607 B.n607 B.n606 585
R1608 B.n254 B.n253 585
R1609 B.n255 B.n254 585
R1610 B.n599 B.n598 585
R1611 B.n600 B.n599 585
R1612 B.n597 B.n260 585
R1613 B.n260 B.n259 585
R1614 B.n596 B.n595 585
R1615 B.n595 B.n594 585
R1616 B.n262 B.n261 585
R1617 B.n263 B.n262 585
R1618 B.n587 B.n586 585
R1619 B.n588 B.n587 585
R1620 B.n585 B.n268 585
R1621 B.n268 B.n267 585
R1622 B.n584 B.n583 585
R1623 B.n583 B.n582 585
R1624 B.n579 B.n272 585
R1625 B.n578 B.n577 585
R1626 B.n575 B.n273 585
R1627 B.n575 B.n271 585
R1628 B.n574 B.n573 585
R1629 B.n572 B.n571 585
R1630 B.n570 B.n275 585
R1631 B.n568 B.n567 585
R1632 B.n566 B.n276 585
R1633 B.n565 B.n564 585
R1634 B.n562 B.n277 585
R1635 B.n560 B.n559 585
R1636 B.n558 B.n278 585
R1637 B.n557 B.n556 585
R1638 B.n554 B.n279 585
R1639 B.n552 B.n551 585
R1640 B.n550 B.n280 585
R1641 B.n549 B.n548 585
R1642 B.n546 B.n281 585
R1643 B.n544 B.n543 585
R1644 B.n542 B.n282 585
R1645 B.n541 B.n540 585
R1646 B.n538 B.n283 585
R1647 B.n536 B.n535 585
R1648 B.n534 B.n284 585
R1649 B.n533 B.n532 585
R1650 B.n530 B.n285 585
R1651 B.n528 B.n527 585
R1652 B.n526 B.n286 585
R1653 B.n525 B.n524 585
R1654 B.n522 B.n287 585
R1655 B.n520 B.n519 585
R1656 B.n518 B.n288 585
R1657 B.n517 B.n516 585
R1658 B.n514 B.n289 585
R1659 B.n512 B.n511 585
R1660 B.n510 B.n290 585
R1661 B.n509 B.n508 585
R1662 B.n506 B.n291 585
R1663 B.n504 B.n503 585
R1664 B.n502 B.n292 585
R1665 B.n501 B.n500 585
R1666 B.n498 B.n293 585
R1667 B.n496 B.n495 585
R1668 B.n494 B.n294 585
R1669 B.n493 B.n492 585
R1670 B.n490 B.n295 585
R1671 B.n488 B.n487 585
R1672 B.n486 B.n296 585
R1673 B.n485 B.n484 585
R1674 B.n482 B.n297 585
R1675 B.n480 B.n479 585
R1676 B.n478 B.n298 585
R1677 B.n477 B.n476 585
R1678 B.n474 B.n299 585
R1679 B.n472 B.n471 585
R1680 B.n470 B.n300 585
R1681 B.n468 B.n467 585
R1682 B.n465 B.n303 585
R1683 B.n463 B.n462 585
R1684 B.n461 B.n304 585
R1685 B.n460 B.n459 585
R1686 B.n457 B.n305 585
R1687 B.n455 B.n454 585
R1688 B.n453 B.n306 585
R1689 B.n452 B.n451 585
R1690 B.n449 B.n307 585
R1691 B.n447 B.n446 585
R1692 B.n445 B.n308 585
R1693 B.n444 B.n443 585
R1694 B.n441 B.n312 585
R1695 B.n439 B.n438 585
R1696 B.n437 B.n313 585
R1697 B.n436 B.n435 585
R1698 B.n433 B.n314 585
R1699 B.n431 B.n430 585
R1700 B.n429 B.n315 585
R1701 B.n428 B.n427 585
R1702 B.n425 B.n316 585
R1703 B.n423 B.n422 585
R1704 B.n421 B.n317 585
R1705 B.n420 B.n419 585
R1706 B.n417 B.n318 585
R1707 B.n415 B.n414 585
R1708 B.n413 B.n319 585
R1709 B.n412 B.n411 585
R1710 B.n409 B.n320 585
R1711 B.n407 B.n406 585
R1712 B.n405 B.n321 585
R1713 B.n404 B.n403 585
R1714 B.n401 B.n322 585
R1715 B.n399 B.n398 585
R1716 B.n397 B.n323 585
R1717 B.n396 B.n395 585
R1718 B.n393 B.n324 585
R1719 B.n391 B.n390 585
R1720 B.n389 B.n325 585
R1721 B.n388 B.n387 585
R1722 B.n385 B.n326 585
R1723 B.n383 B.n382 585
R1724 B.n381 B.n327 585
R1725 B.n380 B.n379 585
R1726 B.n377 B.n328 585
R1727 B.n375 B.n374 585
R1728 B.n373 B.n329 585
R1729 B.n372 B.n371 585
R1730 B.n369 B.n330 585
R1731 B.n367 B.n366 585
R1732 B.n365 B.n331 585
R1733 B.n364 B.n363 585
R1734 B.n361 B.n332 585
R1735 B.n359 B.n358 585
R1736 B.n357 B.n333 585
R1737 B.n356 B.n355 585
R1738 B.n353 B.n334 585
R1739 B.n351 B.n350 585
R1740 B.n349 B.n335 585
R1741 B.n348 B.n347 585
R1742 B.n345 B.n336 585
R1743 B.n343 B.n342 585
R1744 B.n341 B.n337 585
R1745 B.n340 B.n339 585
R1746 B.n270 B.n269 585
R1747 B.n271 B.n270 585
R1748 B.n581 B.n580 585
R1749 B.n582 B.n581 585
R1750 B.n266 B.n265 585
R1751 B.n267 B.n266 585
R1752 B.n590 B.n589 585
R1753 B.n589 B.n588 585
R1754 B.n591 B.n264 585
R1755 B.n264 B.n263 585
R1756 B.n593 B.n592 585
R1757 B.n594 B.n593 585
R1758 B.n258 B.n257 585
R1759 B.n259 B.n258 585
R1760 B.n602 B.n601 585
R1761 B.n601 B.n600 585
R1762 B.n603 B.n256 585
R1763 B.n256 B.n255 585
R1764 B.n605 B.n604 585
R1765 B.n606 B.n605 585
R1766 B.n250 B.n249 585
R1767 B.n251 B.n250 585
R1768 B.n614 B.n613 585
R1769 B.n613 B.n612 585
R1770 B.n615 B.n248 585
R1771 B.n248 B.n247 585
R1772 B.n617 B.n616 585
R1773 B.n618 B.n617 585
R1774 B.n242 B.n241 585
R1775 B.n243 B.n242 585
R1776 B.n626 B.n625 585
R1777 B.n625 B.n624 585
R1778 B.n627 B.n240 585
R1779 B.n240 B.n239 585
R1780 B.n629 B.n628 585
R1781 B.n630 B.n629 585
R1782 B.n234 B.n233 585
R1783 B.n235 B.n234 585
R1784 B.n638 B.n637 585
R1785 B.n637 B.n636 585
R1786 B.n639 B.n232 585
R1787 B.n232 B.n231 585
R1788 B.n641 B.n640 585
R1789 B.n642 B.n641 585
R1790 B.n226 B.n225 585
R1791 B.n227 B.n226 585
R1792 B.n650 B.n649 585
R1793 B.n649 B.n648 585
R1794 B.n651 B.n224 585
R1795 B.n224 B.n223 585
R1796 B.n653 B.n652 585
R1797 B.n654 B.n653 585
R1798 B.n218 B.n217 585
R1799 B.n219 B.n218 585
R1800 B.n662 B.n661 585
R1801 B.n661 B.n660 585
R1802 B.n663 B.n216 585
R1803 B.n216 B.n214 585
R1804 B.n665 B.n664 585
R1805 B.n666 B.n665 585
R1806 B.n210 B.n209 585
R1807 B.n215 B.n210 585
R1808 B.n674 B.n673 585
R1809 B.n673 B.n672 585
R1810 B.n675 B.n208 585
R1811 B.n208 B.n207 585
R1812 B.n677 B.n676 585
R1813 B.n678 B.n677 585
R1814 B.n202 B.n201 585
R1815 B.n203 B.n202 585
R1816 B.n686 B.n685 585
R1817 B.n685 B.n684 585
R1818 B.n687 B.n200 585
R1819 B.n200 B.n199 585
R1820 B.n689 B.n688 585
R1821 B.n690 B.n689 585
R1822 B.n194 B.n193 585
R1823 B.n195 B.n194 585
R1824 B.n698 B.n697 585
R1825 B.n697 B.n696 585
R1826 B.n699 B.n192 585
R1827 B.n192 B.n191 585
R1828 B.n701 B.n700 585
R1829 B.n702 B.n701 585
R1830 B.n186 B.n185 585
R1831 B.n187 B.n186 585
R1832 B.n710 B.n709 585
R1833 B.n709 B.n708 585
R1834 B.n711 B.n184 585
R1835 B.n184 B.n183 585
R1836 B.n713 B.n712 585
R1837 B.n714 B.n713 585
R1838 B.n178 B.n177 585
R1839 B.n179 B.n178 585
R1840 B.n723 B.n722 585
R1841 B.n722 B.n721 585
R1842 B.n724 B.n176 585
R1843 B.n720 B.n176 585
R1844 B.n726 B.n725 585
R1845 B.n727 B.n726 585
R1846 B.n171 B.n170 585
R1847 B.n172 B.n171 585
R1848 B.n736 B.n735 585
R1849 B.n735 B.n734 585
R1850 B.n737 B.n169 585
R1851 B.n169 B.n168 585
R1852 B.n739 B.n738 585
R1853 B.n740 B.n739 585
R1854 B.n2 B.n0 585
R1855 B.n4 B.n2 585
R1856 B.n3 B.n1 585
R1857 B.n1164 B.n3 585
R1858 B.n1162 B.n1161 585
R1859 B.n1163 B.n1162 585
R1860 B.n1160 B.n9 585
R1861 B.n9 B.n8 585
R1862 B.n1159 B.n1158 585
R1863 B.n1158 B.n1157 585
R1864 B.n11 B.n10 585
R1865 B.n1156 B.n11 585
R1866 B.n1154 B.n1153 585
R1867 B.n1155 B.n1154 585
R1868 B.n1152 B.n15 585
R1869 B.n18 B.n15 585
R1870 B.n1151 B.n1150 585
R1871 B.n1150 B.n1149 585
R1872 B.n17 B.n16 585
R1873 B.n1148 B.n17 585
R1874 B.n1146 B.n1145 585
R1875 B.n1147 B.n1146 585
R1876 B.n1144 B.n23 585
R1877 B.n23 B.n22 585
R1878 B.n1143 B.n1142 585
R1879 B.n1142 B.n1141 585
R1880 B.n25 B.n24 585
R1881 B.n1140 B.n25 585
R1882 B.n1138 B.n1137 585
R1883 B.n1139 B.n1138 585
R1884 B.n1136 B.n30 585
R1885 B.n30 B.n29 585
R1886 B.n1135 B.n1134 585
R1887 B.n1134 B.n1133 585
R1888 B.n32 B.n31 585
R1889 B.n1132 B.n32 585
R1890 B.n1130 B.n1129 585
R1891 B.n1131 B.n1130 585
R1892 B.n1128 B.n37 585
R1893 B.n37 B.n36 585
R1894 B.n1127 B.n1126 585
R1895 B.n1126 B.n1125 585
R1896 B.n39 B.n38 585
R1897 B.n1124 B.n39 585
R1898 B.n1122 B.n1121 585
R1899 B.n1123 B.n1122 585
R1900 B.n1120 B.n44 585
R1901 B.n44 B.n43 585
R1902 B.n1119 B.n1118 585
R1903 B.n1118 B.n1117 585
R1904 B.n46 B.n45 585
R1905 B.n1116 B.n46 585
R1906 B.n1114 B.n1113 585
R1907 B.n1115 B.n1114 585
R1908 B.n1112 B.n51 585
R1909 B.n51 B.n50 585
R1910 B.n1111 B.n1110 585
R1911 B.n1110 B.n1109 585
R1912 B.n53 B.n52 585
R1913 B.n1108 B.n53 585
R1914 B.n1106 B.n1105 585
R1915 B.n1107 B.n1106 585
R1916 B.n1104 B.n58 585
R1917 B.n58 B.n57 585
R1918 B.n1103 B.n1102 585
R1919 B.n1102 B.n1101 585
R1920 B.n60 B.n59 585
R1921 B.n1100 B.n60 585
R1922 B.n1098 B.n1097 585
R1923 B.n1099 B.n1098 585
R1924 B.n1096 B.n65 585
R1925 B.n65 B.n64 585
R1926 B.n1095 B.n1094 585
R1927 B.n1094 B.n1093 585
R1928 B.n67 B.n66 585
R1929 B.n1092 B.n67 585
R1930 B.n1090 B.n1089 585
R1931 B.n1091 B.n1090 585
R1932 B.n1088 B.n72 585
R1933 B.n72 B.n71 585
R1934 B.n1087 B.n1086 585
R1935 B.n1086 B.n1085 585
R1936 B.n74 B.n73 585
R1937 B.n1084 B.n74 585
R1938 B.n1082 B.n1081 585
R1939 B.n1083 B.n1082 585
R1940 B.n1080 B.n79 585
R1941 B.n79 B.n78 585
R1942 B.n1079 B.n1078 585
R1943 B.n1078 B.n1077 585
R1944 B.n81 B.n80 585
R1945 B.n1076 B.n81 585
R1946 B.n1074 B.n1073 585
R1947 B.n1075 B.n1074 585
R1948 B.n1072 B.n86 585
R1949 B.n86 B.n85 585
R1950 B.n1071 B.n1070 585
R1951 B.n1070 B.n1069 585
R1952 B.n88 B.n87 585
R1953 B.n1068 B.n88 585
R1954 B.n1066 B.n1065 585
R1955 B.n1067 B.n1066 585
R1956 B.n1064 B.n93 585
R1957 B.n93 B.n92 585
R1958 B.n1063 B.n1062 585
R1959 B.n1062 B.n1061 585
R1960 B.n95 B.n94 585
R1961 B.n1060 B.n95 585
R1962 B.n1058 B.n1057 585
R1963 B.n1059 B.n1058 585
R1964 B.n1167 B.n1166 585
R1965 B.n1166 B.n1165 585
R1966 B.n581 B.n272 482.89
R1967 B.n1058 B.n100 482.89
R1968 B.n583 B.n270 482.89
R1969 B.n813 B.n98 482.89
R1970 B.n309 B.t11 428.577
R1971 B.n135 B.t14 428.577
R1972 B.n301 B.t18 428.577
R1973 B.n129 B.t20 428.577
R1974 B.n310 B.t10 368.262
R1975 B.n136 B.t15 368.262
R1976 B.n302 B.t17 368.262
R1977 B.n130 B.t21 368.262
R1978 B.n309 B.t8 355.505
R1979 B.n301 B.t16 355.505
R1980 B.n129 B.t19 355.505
R1981 B.n135 B.t12 355.505
R1982 B.n814 B.n99 256.663
R1983 B.n816 B.n99 256.663
R1984 B.n822 B.n99 256.663
R1985 B.n824 B.n99 256.663
R1986 B.n830 B.n99 256.663
R1987 B.n832 B.n99 256.663
R1988 B.n838 B.n99 256.663
R1989 B.n840 B.n99 256.663
R1990 B.n846 B.n99 256.663
R1991 B.n848 B.n99 256.663
R1992 B.n854 B.n99 256.663
R1993 B.n856 B.n99 256.663
R1994 B.n862 B.n99 256.663
R1995 B.n864 B.n99 256.663
R1996 B.n870 B.n99 256.663
R1997 B.n872 B.n99 256.663
R1998 B.n878 B.n99 256.663
R1999 B.n880 B.n99 256.663
R2000 B.n886 B.n99 256.663
R2001 B.n888 B.n99 256.663
R2002 B.n894 B.n99 256.663
R2003 B.n896 B.n99 256.663
R2004 B.n902 B.n99 256.663
R2005 B.n904 B.n99 256.663
R2006 B.n910 B.n99 256.663
R2007 B.n912 B.n99 256.663
R2008 B.n918 B.n99 256.663
R2009 B.n138 B.n99 256.663
R2010 B.n924 B.n99 256.663
R2011 B.n930 B.n99 256.663
R2012 B.n932 B.n99 256.663
R2013 B.n938 B.n99 256.663
R2014 B.n940 B.n99 256.663
R2015 B.n947 B.n99 256.663
R2016 B.n949 B.n99 256.663
R2017 B.n955 B.n99 256.663
R2018 B.n957 B.n99 256.663
R2019 B.n963 B.n99 256.663
R2020 B.n965 B.n99 256.663
R2021 B.n971 B.n99 256.663
R2022 B.n973 B.n99 256.663
R2023 B.n979 B.n99 256.663
R2024 B.n981 B.n99 256.663
R2025 B.n987 B.n99 256.663
R2026 B.n989 B.n99 256.663
R2027 B.n995 B.n99 256.663
R2028 B.n997 B.n99 256.663
R2029 B.n1003 B.n99 256.663
R2030 B.n1005 B.n99 256.663
R2031 B.n1011 B.n99 256.663
R2032 B.n1013 B.n99 256.663
R2033 B.n1019 B.n99 256.663
R2034 B.n1021 B.n99 256.663
R2035 B.n1027 B.n99 256.663
R2036 B.n1029 B.n99 256.663
R2037 B.n1035 B.n99 256.663
R2038 B.n1037 B.n99 256.663
R2039 B.n1043 B.n99 256.663
R2040 B.n1045 B.n99 256.663
R2041 B.n1051 B.n99 256.663
R2042 B.n1053 B.n99 256.663
R2043 B.n576 B.n271 256.663
R2044 B.n274 B.n271 256.663
R2045 B.n569 B.n271 256.663
R2046 B.n563 B.n271 256.663
R2047 B.n561 B.n271 256.663
R2048 B.n555 B.n271 256.663
R2049 B.n553 B.n271 256.663
R2050 B.n547 B.n271 256.663
R2051 B.n545 B.n271 256.663
R2052 B.n539 B.n271 256.663
R2053 B.n537 B.n271 256.663
R2054 B.n531 B.n271 256.663
R2055 B.n529 B.n271 256.663
R2056 B.n523 B.n271 256.663
R2057 B.n521 B.n271 256.663
R2058 B.n515 B.n271 256.663
R2059 B.n513 B.n271 256.663
R2060 B.n507 B.n271 256.663
R2061 B.n505 B.n271 256.663
R2062 B.n499 B.n271 256.663
R2063 B.n497 B.n271 256.663
R2064 B.n491 B.n271 256.663
R2065 B.n489 B.n271 256.663
R2066 B.n483 B.n271 256.663
R2067 B.n481 B.n271 256.663
R2068 B.n475 B.n271 256.663
R2069 B.n473 B.n271 256.663
R2070 B.n466 B.n271 256.663
R2071 B.n464 B.n271 256.663
R2072 B.n458 B.n271 256.663
R2073 B.n456 B.n271 256.663
R2074 B.n450 B.n271 256.663
R2075 B.n448 B.n271 256.663
R2076 B.n442 B.n271 256.663
R2077 B.n440 B.n271 256.663
R2078 B.n434 B.n271 256.663
R2079 B.n432 B.n271 256.663
R2080 B.n426 B.n271 256.663
R2081 B.n424 B.n271 256.663
R2082 B.n418 B.n271 256.663
R2083 B.n416 B.n271 256.663
R2084 B.n410 B.n271 256.663
R2085 B.n408 B.n271 256.663
R2086 B.n402 B.n271 256.663
R2087 B.n400 B.n271 256.663
R2088 B.n394 B.n271 256.663
R2089 B.n392 B.n271 256.663
R2090 B.n386 B.n271 256.663
R2091 B.n384 B.n271 256.663
R2092 B.n378 B.n271 256.663
R2093 B.n376 B.n271 256.663
R2094 B.n370 B.n271 256.663
R2095 B.n368 B.n271 256.663
R2096 B.n362 B.n271 256.663
R2097 B.n360 B.n271 256.663
R2098 B.n354 B.n271 256.663
R2099 B.n352 B.n271 256.663
R2100 B.n346 B.n271 256.663
R2101 B.n344 B.n271 256.663
R2102 B.n338 B.n271 256.663
R2103 B.n581 B.n266 163.367
R2104 B.n589 B.n266 163.367
R2105 B.n589 B.n264 163.367
R2106 B.n593 B.n264 163.367
R2107 B.n593 B.n258 163.367
R2108 B.n601 B.n258 163.367
R2109 B.n601 B.n256 163.367
R2110 B.n605 B.n256 163.367
R2111 B.n605 B.n250 163.367
R2112 B.n613 B.n250 163.367
R2113 B.n613 B.n248 163.367
R2114 B.n617 B.n248 163.367
R2115 B.n617 B.n242 163.367
R2116 B.n625 B.n242 163.367
R2117 B.n625 B.n240 163.367
R2118 B.n629 B.n240 163.367
R2119 B.n629 B.n234 163.367
R2120 B.n637 B.n234 163.367
R2121 B.n637 B.n232 163.367
R2122 B.n641 B.n232 163.367
R2123 B.n641 B.n226 163.367
R2124 B.n649 B.n226 163.367
R2125 B.n649 B.n224 163.367
R2126 B.n653 B.n224 163.367
R2127 B.n653 B.n218 163.367
R2128 B.n661 B.n218 163.367
R2129 B.n661 B.n216 163.367
R2130 B.n665 B.n216 163.367
R2131 B.n665 B.n210 163.367
R2132 B.n673 B.n210 163.367
R2133 B.n673 B.n208 163.367
R2134 B.n677 B.n208 163.367
R2135 B.n677 B.n202 163.367
R2136 B.n685 B.n202 163.367
R2137 B.n685 B.n200 163.367
R2138 B.n689 B.n200 163.367
R2139 B.n689 B.n194 163.367
R2140 B.n697 B.n194 163.367
R2141 B.n697 B.n192 163.367
R2142 B.n701 B.n192 163.367
R2143 B.n701 B.n186 163.367
R2144 B.n709 B.n186 163.367
R2145 B.n709 B.n184 163.367
R2146 B.n713 B.n184 163.367
R2147 B.n713 B.n178 163.367
R2148 B.n722 B.n178 163.367
R2149 B.n722 B.n176 163.367
R2150 B.n726 B.n176 163.367
R2151 B.n726 B.n171 163.367
R2152 B.n735 B.n171 163.367
R2153 B.n735 B.n169 163.367
R2154 B.n739 B.n169 163.367
R2155 B.n739 B.n2 163.367
R2156 B.n1166 B.n2 163.367
R2157 B.n1166 B.n3 163.367
R2158 B.n1162 B.n3 163.367
R2159 B.n1162 B.n9 163.367
R2160 B.n1158 B.n9 163.367
R2161 B.n1158 B.n11 163.367
R2162 B.n1154 B.n11 163.367
R2163 B.n1154 B.n15 163.367
R2164 B.n1150 B.n15 163.367
R2165 B.n1150 B.n17 163.367
R2166 B.n1146 B.n17 163.367
R2167 B.n1146 B.n23 163.367
R2168 B.n1142 B.n23 163.367
R2169 B.n1142 B.n25 163.367
R2170 B.n1138 B.n25 163.367
R2171 B.n1138 B.n30 163.367
R2172 B.n1134 B.n30 163.367
R2173 B.n1134 B.n32 163.367
R2174 B.n1130 B.n32 163.367
R2175 B.n1130 B.n37 163.367
R2176 B.n1126 B.n37 163.367
R2177 B.n1126 B.n39 163.367
R2178 B.n1122 B.n39 163.367
R2179 B.n1122 B.n44 163.367
R2180 B.n1118 B.n44 163.367
R2181 B.n1118 B.n46 163.367
R2182 B.n1114 B.n46 163.367
R2183 B.n1114 B.n51 163.367
R2184 B.n1110 B.n51 163.367
R2185 B.n1110 B.n53 163.367
R2186 B.n1106 B.n53 163.367
R2187 B.n1106 B.n58 163.367
R2188 B.n1102 B.n58 163.367
R2189 B.n1102 B.n60 163.367
R2190 B.n1098 B.n60 163.367
R2191 B.n1098 B.n65 163.367
R2192 B.n1094 B.n65 163.367
R2193 B.n1094 B.n67 163.367
R2194 B.n1090 B.n67 163.367
R2195 B.n1090 B.n72 163.367
R2196 B.n1086 B.n72 163.367
R2197 B.n1086 B.n74 163.367
R2198 B.n1082 B.n74 163.367
R2199 B.n1082 B.n79 163.367
R2200 B.n1078 B.n79 163.367
R2201 B.n1078 B.n81 163.367
R2202 B.n1074 B.n81 163.367
R2203 B.n1074 B.n86 163.367
R2204 B.n1070 B.n86 163.367
R2205 B.n1070 B.n88 163.367
R2206 B.n1066 B.n88 163.367
R2207 B.n1066 B.n93 163.367
R2208 B.n1062 B.n93 163.367
R2209 B.n1062 B.n95 163.367
R2210 B.n1058 B.n95 163.367
R2211 B.n577 B.n575 163.367
R2212 B.n575 B.n574 163.367
R2213 B.n571 B.n570 163.367
R2214 B.n568 B.n276 163.367
R2215 B.n564 B.n562 163.367
R2216 B.n560 B.n278 163.367
R2217 B.n556 B.n554 163.367
R2218 B.n552 B.n280 163.367
R2219 B.n548 B.n546 163.367
R2220 B.n544 B.n282 163.367
R2221 B.n540 B.n538 163.367
R2222 B.n536 B.n284 163.367
R2223 B.n532 B.n530 163.367
R2224 B.n528 B.n286 163.367
R2225 B.n524 B.n522 163.367
R2226 B.n520 B.n288 163.367
R2227 B.n516 B.n514 163.367
R2228 B.n512 B.n290 163.367
R2229 B.n508 B.n506 163.367
R2230 B.n504 B.n292 163.367
R2231 B.n500 B.n498 163.367
R2232 B.n496 B.n294 163.367
R2233 B.n492 B.n490 163.367
R2234 B.n488 B.n296 163.367
R2235 B.n484 B.n482 163.367
R2236 B.n480 B.n298 163.367
R2237 B.n476 B.n474 163.367
R2238 B.n472 B.n300 163.367
R2239 B.n467 B.n465 163.367
R2240 B.n463 B.n304 163.367
R2241 B.n459 B.n457 163.367
R2242 B.n455 B.n306 163.367
R2243 B.n451 B.n449 163.367
R2244 B.n447 B.n308 163.367
R2245 B.n443 B.n441 163.367
R2246 B.n439 B.n313 163.367
R2247 B.n435 B.n433 163.367
R2248 B.n431 B.n315 163.367
R2249 B.n427 B.n425 163.367
R2250 B.n423 B.n317 163.367
R2251 B.n419 B.n417 163.367
R2252 B.n415 B.n319 163.367
R2253 B.n411 B.n409 163.367
R2254 B.n407 B.n321 163.367
R2255 B.n403 B.n401 163.367
R2256 B.n399 B.n323 163.367
R2257 B.n395 B.n393 163.367
R2258 B.n391 B.n325 163.367
R2259 B.n387 B.n385 163.367
R2260 B.n383 B.n327 163.367
R2261 B.n379 B.n377 163.367
R2262 B.n375 B.n329 163.367
R2263 B.n371 B.n369 163.367
R2264 B.n367 B.n331 163.367
R2265 B.n363 B.n361 163.367
R2266 B.n359 B.n333 163.367
R2267 B.n355 B.n353 163.367
R2268 B.n351 B.n335 163.367
R2269 B.n347 B.n345 163.367
R2270 B.n343 B.n337 163.367
R2271 B.n339 B.n270 163.367
R2272 B.n583 B.n268 163.367
R2273 B.n587 B.n268 163.367
R2274 B.n587 B.n262 163.367
R2275 B.n595 B.n262 163.367
R2276 B.n595 B.n260 163.367
R2277 B.n599 B.n260 163.367
R2278 B.n599 B.n254 163.367
R2279 B.n607 B.n254 163.367
R2280 B.n607 B.n252 163.367
R2281 B.n611 B.n252 163.367
R2282 B.n611 B.n246 163.367
R2283 B.n619 B.n246 163.367
R2284 B.n619 B.n244 163.367
R2285 B.n623 B.n244 163.367
R2286 B.n623 B.n238 163.367
R2287 B.n631 B.n238 163.367
R2288 B.n631 B.n236 163.367
R2289 B.n635 B.n236 163.367
R2290 B.n635 B.n230 163.367
R2291 B.n643 B.n230 163.367
R2292 B.n643 B.n228 163.367
R2293 B.n647 B.n228 163.367
R2294 B.n647 B.n222 163.367
R2295 B.n655 B.n222 163.367
R2296 B.n655 B.n220 163.367
R2297 B.n659 B.n220 163.367
R2298 B.n659 B.n213 163.367
R2299 B.n667 B.n213 163.367
R2300 B.n667 B.n211 163.367
R2301 B.n671 B.n211 163.367
R2302 B.n671 B.n206 163.367
R2303 B.n679 B.n206 163.367
R2304 B.n679 B.n204 163.367
R2305 B.n683 B.n204 163.367
R2306 B.n683 B.n198 163.367
R2307 B.n691 B.n198 163.367
R2308 B.n691 B.n196 163.367
R2309 B.n695 B.n196 163.367
R2310 B.n695 B.n190 163.367
R2311 B.n703 B.n190 163.367
R2312 B.n703 B.n188 163.367
R2313 B.n707 B.n188 163.367
R2314 B.n707 B.n182 163.367
R2315 B.n715 B.n182 163.367
R2316 B.n715 B.n180 163.367
R2317 B.n719 B.n180 163.367
R2318 B.n719 B.n175 163.367
R2319 B.n728 B.n175 163.367
R2320 B.n728 B.n173 163.367
R2321 B.n733 B.n173 163.367
R2322 B.n733 B.n167 163.367
R2323 B.n741 B.n167 163.367
R2324 B.n742 B.n741 163.367
R2325 B.n742 B.n5 163.367
R2326 B.n6 B.n5 163.367
R2327 B.n7 B.n6 163.367
R2328 B.n747 B.n7 163.367
R2329 B.n747 B.n12 163.367
R2330 B.n13 B.n12 163.367
R2331 B.n14 B.n13 163.367
R2332 B.n752 B.n14 163.367
R2333 B.n752 B.n19 163.367
R2334 B.n20 B.n19 163.367
R2335 B.n21 B.n20 163.367
R2336 B.n757 B.n21 163.367
R2337 B.n757 B.n26 163.367
R2338 B.n27 B.n26 163.367
R2339 B.n28 B.n27 163.367
R2340 B.n762 B.n28 163.367
R2341 B.n762 B.n33 163.367
R2342 B.n34 B.n33 163.367
R2343 B.n35 B.n34 163.367
R2344 B.n767 B.n35 163.367
R2345 B.n767 B.n40 163.367
R2346 B.n41 B.n40 163.367
R2347 B.n42 B.n41 163.367
R2348 B.n772 B.n42 163.367
R2349 B.n772 B.n47 163.367
R2350 B.n48 B.n47 163.367
R2351 B.n49 B.n48 163.367
R2352 B.n777 B.n49 163.367
R2353 B.n777 B.n54 163.367
R2354 B.n55 B.n54 163.367
R2355 B.n56 B.n55 163.367
R2356 B.n782 B.n56 163.367
R2357 B.n782 B.n61 163.367
R2358 B.n62 B.n61 163.367
R2359 B.n63 B.n62 163.367
R2360 B.n787 B.n63 163.367
R2361 B.n787 B.n68 163.367
R2362 B.n69 B.n68 163.367
R2363 B.n70 B.n69 163.367
R2364 B.n792 B.n70 163.367
R2365 B.n792 B.n75 163.367
R2366 B.n76 B.n75 163.367
R2367 B.n77 B.n76 163.367
R2368 B.n797 B.n77 163.367
R2369 B.n797 B.n82 163.367
R2370 B.n83 B.n82 163.367
R2371 B.n84 B.n83 163.367
R2372 B.n802 B.n84 163.367
R2373 B.n802 B.n89 163.367
R2374 B.n90 B.n89 163.367
R2375 B.n91 B.n90 163.367
R2376 B.n807 B.n91 163.367
R2377 B.n807 B.n96 163.367
R2378 B.n97 B.n96 163.367
R2379 B.n98 B.n97 163.367
R2380 B.n1054 B.n1052 163.367
R2381 B.n1050 B.n102 163.367
R2382 B.n1046 B.n1044 163.367
R2383 B.n1042 B.n104 163.367
R2384 B.n1038 B.n1036 163.367
R2385 B.n1034 B.n106 163.367
R2386 B.n1030 B.n1028 163.367
R2387 B.n1026 B.n108 163.367
R2388 B.n1022 B.n1020 163.367
R2389 B.n1018 B.n110 163.367
R2390 B.n1014 B.n1012 163.367
R2391 B.n1010 B.n112 163.367
R2392 B.n1006 B.n1004 163.367
R2393 B.n1002 B.n114 163.367
R2394 B.n998 B.n996 163.367
R2395 B.n994 B.n116 163.367
R2396 B.n990 B.n988 163.367
R2397 B.n986 B.n118 163.367
R2398 B.n982 B.n980 163.367
R2399 B.n978 B.n120 163.367
R2400 B.n974 B.n972 163.367
R2401 B.n970 B.n122 163.367
R2402 B.n966 B.n964 163.367
R2403 B.n962 B.n124 163.367
R2404 B.n958 B.n956 163.367
R2405 B.n954 B.n126 163.367
R2406 B.n950 B.n948 163.367
R2407 B.n946 B.n128 163.367
R2408 B.n941 B.n939 163.367
R2409 B.n937 B.n132 163.367
R2410 B.n933 B.n931 163.367
R2411 B.n929 B.n134 163.367
R2412 B.n925 B.n923 163.367
R2413 B.n920 B.n919 163.367
R2414 B.n917 B.n140 163.367
R2415 B.n913 B.n911 163.367
R2416 B.n909 B.n142 163.367
R2417 B.n905 B.n903 163.367
R2418 B.n901 B.n144 163.367
R2419 B.n897 B.n895 163.367
R2420 B.n893 B.n146 163.367
R2421 B.n889 B.n887 163.367
R2422 B.n885 B.n148 163.367
R2423 B.n881 B.n879 163.367
R2424 B.n877 B.n150 163.367
R2425 B.n873 B.n871 163.367
R2426 B.n869 B.n152 163.367
R2427 B.n865 B.n863 163.367
R2428 B.n861 B.n154 163.367
R2429 B.n857 B.n855 163.367
R2430 B.n853 B.n156 163.367
R2431 B.n849 B.n847 163.367
R2432 B.n845 B.n158 163.367
R2433 B.n841 B.n839 163.367
R2434 B.n837 B.n160 163.367
R2435 B.n833 B.n831 163.367
R2436 B.n829 B.n162 163.367
R2437 B.n825 B.n823 163.367
R2438 B.n821 B.n164 163.367
R2439 B.n817 B.n815 163.367
R2440 B.n576 B.n272 71.676
R2441 B.n574 B.n274 71.676
R2442 B.n570 B.n569 71.676
R2443 B.n563 B.n276 71.676
R2444 B.n562 B.n561 71.676
R2445 B.n555 B.n278 71.676
R2446 B.n554 B.n553 71.676
R2447 B.n547 B.n280 71.676
R2448 B.n546 B.n545 71.676
R2449 B.n539 B.n282 71.676
R2450 B.n538 B.n537 71.676
R2451 B.n531 B.n284 71.676
R2452 B.n530 B.n529 71.676
R2453 B.n523 B.n286 71.676
R2454 B.n522 B.n521 71.676
R2455 B.n515 B.n288 71.676
R2456 B.n514 B.n513 71.676
R2457 B.n507 B.n290 71.676
R2458 B.n506 B.n505 71.676
R2459 B.n499 B.n292 71.676
R2460 B.n498 B.n497 71.676
R2461 B.n491 B.n294 71.676
R2462 B.n490 B.n489 71.676
R2463 B.n483 B.n296 71.676
R2464 B.n482 B.n481 71.676
R2465 B.n475 B.n298 71.676
R2466 B.n474 B.n473 71.676
R2467 B.n466 B.n300 71.676
R2468 B.n465 B.n464 71.676
R2469 B.n458 B.n304 71.676
R2470 B.n457 B.n456 71.676
R2471 B.n450 B.n306 71.676
R2472 B.n449 B.n448 71.676
R2473 B.n442 B.n308 71.676
R2474 B.n441 B.n440 71.676
R2475 B.n434 B.n313 71.676
R2476 B.n433 B.n432 71.676
R2477 B.n426 B.n315 71.676
R2478 B.n425 B.n424 71.676
R2479 B.n418 B.n317 71.676
R2480 B.n417 B.n416 71.676
R2481 B.n410 B.n319 71.676
R2482 B.n409 B.n408 71.676
R2483 B.n402 B.n321 71.676
R2484 B.n401 B.n400 71.676
R2485 B.n394 B.n323 71.676
R2486 B.n393 B.n392 71.676
R2487 B.n386 B.n325 71.676
R2488 B.n385 B.n384 71.676
R2489 B.n378 B.n327 71.676
R2490 B.n377 B.n376 71.676
R2491 B.n370 B.n329 71.676
R2492 B.n369 B.n368 71.676
R2493 B.n362 B.n331 71.676
R2494 B.n361 B.n360 71.676
R2495 B.n354 B.n333 71.676
R2496 B.n353 B.n352 71.676
R2497 B.n346 B.n335 71.676
R2498 B.n345 B.n344 71.676
R2499 B.n338 B.n337 71.676
R2500 B.n1053 B.n100 71.676
R2501 B.n1052 B.n1051 71.676
R2502 B.n1045 B.n102 71.676
R2503 B.n1044 B.n1043 71.676
R2504 B.n1037 B.n104 71.676
R2505 B.n1036 B.n1035 71.676
R2506 B.n1029 B.n106 71.676
R2507 B.n1028 B.n1027 71.676
R2508 B.n1021 B.n108 71.676
R2509 B.n1020 B.n1019 71.676
R2510 B.n1013 B.n110 71.676
R2511 B.n1012 B.n1011 71.676
R2512 B.n1005 B.n112 71.676
R2513 B.n1004 B.n1003 71.676
R2514 B.n997 B.n114 71.676
R2515 B.n996 B.n995 71.676
R2516 B.n989 B.n116 71.676
R2517 B.n988 B.n987 71.676
R2518 B.n981 B.n118 71.676
R2519 B.n980 B.n979 71.676
R2520 B.n973 B.n120 71.676
R2521 B.n972 B.n971 71.676
R2522 B.n965 B.n122 71.676
R2523 B.n964 B.n963 71.676
R2524 B.n957 B.n124 71.676
R2525 B.n956 B.n955 71.676
R2526 B.n949 B.n126 71.676
R2527 B.n948 B.n947 71.676
R2528 B.n940 B.n128 71.676
R2529 B.n939 B.n938 71.676
R2530 B.n932 B.n132 71.676
R2531 B.n931 B.n930 71.676
R2532 B.n924 B.n134 71.676
R2533 B.n923 B.n138 71.676
R2534 B.n919 B.n918 71.676
R2535 B.n912 B.n140 71.676
R2536 B.n911 B.n910 71.676
R2537 B.n904 B.n142 71.676
R2538 B.n903 B.n902 71.676
R2539 B.n896 B.n144 71.676
R2540 B.n895 B.n894 71.676
R2541 B.n888 B.n146 71.676
R2542 B.n887 B.n886 71.676
R2543 B.n880 B.n148 71.676
R2544 B.n879 B.n878 71.676
R2545 B.n872 B.n150 71.676
R2546 B.n871 B.n870 71.676
R2547 B.n864 B.n152 71.676
R2548 B.n863 B.n862 71.676
R2549 B.n856 B.n154 71.676
R2550 B.n855 B.n854 71.676
R2551 B.n848 B.n156 71.676
R2552 B.n847 B.n846 71.676
R2553 B.n840 B.n158 71.676
R2554 B.n839 B.n838 71.676
R2555 B.n832 B.n160 71.676
R2556 B.n831 B.n830 71.676
R2557 B.n824 B.n162 71.676
R2558 B.n823 B.n822 71.676
R2559 B.n816 B.n164 71.676
R2560 B.n815 B.n814 71.676
R2561 B.n814 B.n813 71.676
R2562 B.n817 B.n816 71.676
R2563 B.n822 B.n821 71.676
R2564 B.n825 B.n824 71.676
R2565 B.n830 B.n829 71.676
R2566 B.n833 B.n832 71.676
R2567 B.n838 B.n837 71.676
R2568 B.n841 B.n840 71.676
R2569 B.n846 B.n845 71.676
R2570 B.n849 B.n848 71.676
R2571 B.n854 B.n853 71.676
R2572 B.n857 B.n856 71.676
R2573 B.n862 B.n861 71.676
R2574 B.n865 B.n864 71.676
R2575 B.n870 B.n869 71.676
R2576 B.n873 B.n872 71.676
R2577 B.n878 B.n877 71.676
R2578 B.n881 B.n880 71.676
R2579 B.n886 B.n885 71.676
R2580 B.n889 B.n888 71.676
R2581 B.n894 B.n893 71.676
R2582 B.n897 B.n896 71.676
R2583 B.n902 B.n901 71.676
R2584 B.n905 B.n904 71.676
R2585 B.n910 B.n909 71.676
R2586 B.n913 B.n912 71.676
R2587 B.n918 B.n917 71.676
R2588 B.n920 B.n138 71.676
R2589 B.n925 B.n924 71.676
R2590 B.n930 B.n929 71.676
R2591 B.n933 B.n932 71.676
R2592 B.n938 B.n937 71.676
R2593 B.n941 B.n940 71.676
R2594 B.n947 B.n946 71.676
R2595 B.n950 B.n949 71.676
R2596 B.n955 B.n954 71.676
R2597 B.n958 B.n957 71.676
R2598 B.n963 B.n962 71.676
R2599 B.n966 B.n965 71.676
R2600 B.n971 B.n970 71.676
R2601 B.n974 B.n973 71.676
R2602 B.n979 B.n978 71.676
R2603 B.n982 B.n981 71.676
R2604 B.n987 B.n986 71.676
R2605 B.n990 B.n989 71.676
R2606 B.n995 B.n994 71.676
R2607 B.n998 B.n997 71.676
R2608 B.n1003 B.n1002 71.676
R2609 B.n1006 B.n1005 71.676
R2610 B.n1011 B.n1010 71.676
R2611 B.n1014 B.n1013 71.676
R2612 B.n1019 B.n1018 71.676
R2613 B.n1022 B.n1021 71.676
R2614 B.n1027 B.n1026 71.676
R2615 B.n1030 B.n1029 71.676
R2616 B.n1035 B.n1034 71.676
R2617 B.n1038 B.n1037 71.676
R2618 B.n1043 B.n1042 71.676
R2619 B.n1046 B.n1045 71.676
R2620 B.n1051 B.n1050 71.676
R2621 B.n1054 B.n1053 71.676
R2622 B.n577 B.n576 71.676
R2623 B.n571 B.n274 71.676
R2624 B.n569 B.n568 71.676
R2625 B.n564 B.n563 71.676
R2626 B.n561 B.n560 71.676
R2627 B.n556 B.n555 71.676
R2628 B.n553 B.n552 71.676
R2629 B.n548 B.n547 71.676
R2630 B.n545 B.n544 71.676
R2631 B.n540 B.n539 71.676
R2632 B.n537 B.n536 71.676
R2633 B.n532 B.n531 71.676
R2634 B.n529 B.n528 71.676
R2635 B.n524 B.n523 71.676
R2636 B.n521 B.n520 71.676
R2637 B.n516 B.n515 71.676
R2638 B.n513 B.n512 71.676
R2639 B.n508 B.n507 71.676
R2640 B.n505 B.n504 71.676
R2641 B.n500 B.n499 71.676
R2642 B.n497 B.n496 71.676
R2643 B.n492 B.n491 71.676
R2644 B.n489 B.n488 71.676
R2645 B.n484 B.n483 71.676
R2646 B.n481 B.n480 71.676
R2647 B.n476 B.n475 71.676
R2648 B.n473 B.n472 71.676
R2649 B.n467 B.n466 71.676
R2650 B.n464 B.n463 71.676
R2651 B.n459 B.n458 71.676
R2652 B.n456 B.n455 71.676
R2653 B.n451 B.n450 71.676
R2654 B.n448 B.n447 71.676
R2655 B.n443 B.n442 71.676
R2656 B.n440 B.n439 71.676
R2657 B.n435 B.n434 71.676
R2658 B.n432 B.n431 71.676
R2659 B.n427 B.n426 71.676
R2660 B.n424 B.n423 71.676
R2661 B.n419 B.n418 71.676
R2662 B.n416 B.n415 71.676
R2663 B.n411 B.n410 71.676
R2664 B.n408 B.n407 71.676
R2665 B.n403 B.n402 71.676
R2666 B.n400 B.n399 71.676
R2667 B.n395 B.n394 71.676
R2668 B.n392 B.n391 71.676
R2669 B.n387 B.n386 71.676
R2670 B.n384 B.n383 71.676
R2671 B.n379 B.n378 71.676
R2672 B.n376 B.n375 71.676
R2673 B.n371 B.n370 71.676
R2674 B.n368 B.n367 71.676
R2675 B.n363 B.n362 71.676
R2676 B.n360 B.n359 71.676
R2677 B.n355 B.n354 71.676
R2678 B.n352 B.n351 71.676
R2679 B.n347 B.n346 71.676
R2680 B.n344 B.n343 71.676
R2681 B.n339 B.n338 71.676
R2682 B.n310 B.n309 60.3157
R2683 B.n302 B.n301 60.3157
R2684 B.n130 B.n129 60.3157
R2685 B.n136 B.n135 60.3157
R2686 B.n311 B.n310 59.5399
R2687 B.n469 B.n302 59.5399
R2688 B.n944 B.n130 59.5399
R2689 B.n137 B.n136 59.5399
R2690 B.n582 B.n271 55.8531
R2691 B.n1059 B.n99 55.8531
R2692 B.n582 B.n267 33.6109
R2693 B.n588 B.n267 33.6109
R2694 B.n588 B.n263 33.6109
R2695 B.n594 B.n263 33.6109
R2696 B.n594 B.n259 33.6109
R2697 B.n600 B.n259 33.6109
R2698 B.n600 B.n255 33.6109
R2699 B.n606 B.n255 33.6109
R2700 B.n612 B.n251 33.6109
R2701 B.n612 B.n247 33.6109
R2702 B.n618 B.n247 33.6109
R2703 B.n618 B.n243 33.6109
R2704 B.n624 B.n243 33.6109
R2705 B.n624 B.n239 33.6109
R2706 B.n630 B.n239 33.6109
R2707 B.n630 B.n235 33.6109
R2708 B.n636 B.n235 33.6109
R2709 B.n636 B.n231 33.6109
R2710 B.n642 B.n231 33.6109
R2711 B.n648 B.n227 33.6109
R2712 B.n648 B.n223 33.6109
R2713 B.n654 B.n223 33.6109
R2714 B.n654 B.n219 33.6109
R2715 B.n660 B.n219 33.6109
R2716 B.n660 B.n214 33.6109
R2717 B.n666 B.n214 33.6109
R2718 B.n666 B.n215 33.6109
R2719 B.n672 B.n207 33.6109
R2720 B.n678 B.n207 33.6109
R2721 B.n678 B.n203 33.6109
R2722 B.n684 B.n203 33.6109
R2723 B.n684 B.n199 33.6109
R2724 B.n690 B.n199 33.6109
R2725 B.n690 B.n195 33.6109
R2726 B.n696 B.n195 33.6109
R2727 B.n702 B.n191 33.6109
R2728 B.n702 B.n187 33.6109
R2729 B.n708 B.n187 33.6109
R2730 B.n708 B.n183 33.6109
R2731 B.n714 B.n183 33.6109
R2732 B.n714 B.n179 33.6109
R2733 B.n721 B.n179 33.6109
R2734 B.n721 B.n720 33.6109
R2735 B.n727 B.n172 33.6109
R2736 B.n734 B.n172 33.6109
R2737 B.n734 B.n168 33.6109
R2738 B.n740 B.n168 33.6109
R2739 B.n740 B.n4 33.6109
R2740 B.n1165 B.n4 33.6109
R2741 B.n1165 B.n1164 33.6109
R2742 B.n1164 B.n1163 33.6109
R2743 B.n1163 B.n8 33.6109
R2744 B.n1157 B.n8 33.6109
R2745 B.n1157 B.n1156 33.6109
R2746 B.n1156 B.n1155 33.6109
R2747 B.n1149 B.n18 33.6109
R2748 B.n1149 B.n1148 33.6109
R2749 B.n1148 B.n1147 33.6109
R2750 B.n1147 B.n22 33.6109
R2751 B.n1141 B.n22 33.6109
R2752 B.n1141 B.n1140 33.6109
R2753 B.n1140 B.n1139 33.6109
R2754 B.n1139 B.n29 33.6109
R2755 B.n1133 B.n1132 33.6109
R2756 B.n1132 B.n1131 33.6109
R2757 B.n1131 B.n36 33.6109
R2758 B.n1125 B.n36 33.6109
R2759 B.n1125 B.n1124 33.6109
R2760 B.n1124 B.n1123 33.6109
R2761 B.n1123 B.n43 33.6109
R2762 B.n1117 B.n43 33.6109
R2763 B.n1116 B.n1115 33.6109
R2764 B.n1115 B.n50 33.6109
R2765 B.n1109 B.n50 33.6109
R2766 B.n1109 B.n1108 33.6109
R2767 B.n1108 B.n1107 33.6109
R2768 B.n1107 B.n57 33.6109
R2769 B.n1101 B.n57 33.6109
R2770 B.n1101 B.n1100 33.6109
R2771 B.n1099 B.n64 33.6109
R2772 B.n1093 B.n64 33.6109
R2773 B.n1093 B.n1092 33.6109
R2774 B.n1092 B.n1091 33.6109
R2775 B.n1091 B.n71 33.6109
R2776 B.n1085 B.n71 33.6109
R2777 B.n1085 B.n1084 33.6109
R2778 B.n1084 B.n1083 33.6109
R2779 B.n1083 B.n78 33.6109
R2780 B.n1077 B.n78 33.6109
R2781 B.n1077 B.n1076 33.6109
R2782 B.n1075 B.n85 33.6109
R2783 B.n1069 B.n85 33.6109
R2784 B.n1069 B.n1068 33.6109
R2785 B.n1068 B.n1067 33.6109
R2786 B.n1067 B.n92 33.6109
R2787 B.n1061 B.n92 33.6109
R2788 B.n1061 B.n1060 33.6109
R2789 B.n1060 B.n1059 33.6109
R2790 B.t9 B.n251 32.6224
R2791 B.n1076 B.t13 32.6224
R2792 B.n1057 B.n1056 31.3761
R2793 B.n812 B.n811 31.3761
R2794 B.n584 B.n269 31.3761
R2795 B.n580 B.n579 31.3761
R2796 B.n720 B.t7 27.6797
R2797 B.n18 B.t5 27.6797
R2798 B.n696 B.t3 22.737
R2799 B.n1133 B.t6 22.737
R2800 B.t4 B.n227 20.7599
R2801 B.n1100 B.t2 20.7599
R2802 B B.n1167 18.0485
R2803 B.n215 B.t1 17.7943
R2804 B.t0 B.n1116 17.7943
R2805 B.n672 B.t1 15.8172
R2806 B.n1117 B.t0 15.8172
R2807 B.n642 B.t4 12.8515
R2808 B.t2 B.n1099 12.8515
R2809 B.t3 B.n191 10.8745
R2810 B.t6 B.n29 10.8745
R2811 B.n1056 B.n1055 10.6151
R2812 B.n1055 B.n101 10.6151
R2813 B.n1049 B.n101 10.6151
R2814 B.n1049 B.n1048 10.6151
R2815 B.n1048 B.n1047 10.6151
R2816 B.n1047 B.n103 10.6151
R2817 B.n1041 B.n103 10.6151
R2818 B.n1041 B.n1040 10.6151
R2819 B.n1040 B.n1039 10.6151
R2820 B.n1039 B.n105 10.6151
R2821 B.n1033 B.n105 10.6151
R2822 B.n1033 B.n1032 10.6151
R2823 B.n1032 B.n1031 10.6151
R2824 B.n1031 B.n107 10.6151
R2825 B.n1025 B.n107 10.6151
R2826 B.n1025 B.n1024 10.6151
R2827 B.n1024 B.n1023 10.6151
R2828 B.n1023 B.n109 10.6151
R2829 B.n1017 B.n109 10.6151
R2830 B.n1017 B.n1016 10.6151
R2831 B.n1016 B.n1015 10.6151
R2832 B.n1015 B.n111 10.6151
R2833 B.n1009 B.n111 10.6151
R2834 B.n1009 B.n1008 10.6151
R2835 B.n1008 B.n1007 10.6151
R2836 B.n1007 B.n113 10.6151
R2837 B.n1001 B.n113 10.6151
R2838 B.n1001 B.n1000 10.6151
R2839 B.n1000 B.n999 10.6151
R2840 B.n999 B.n115 10.6151
R2841 B.n993 B.n115 10.6151
R2842 B.n993 B.n992 10.6151
R2843 B.n992 B.n991 10.6151
R2844 B.n991 B.n117 10.6151
R2845 B.n985 B.n117 10.6151
R2846 B.n985 B.n984 10.6151
R2847 B.n984 B.n983 10.6151
R2848 B.n983 B.n119 10.6151
R2849 B.n977 B.n119 10.6151
R2850 B.n977 B.n976 10.6151
R2851 B.n976 B.n975 10.6151
R2852 B.n975 B.n121 10.6151
R2853 B.n969 B.n121 10.6151
R2854 B.n969 B.n968 10.6151
R2855 B.n968 B.n967 10.6151
R2856 B.n967 B.n123 10.6151
R2857 B.n961 B.n123 10.6151
R2858 B.n961 B.n960 10.6151
R2859 B.n960 B.n959 10.6151
R2860 B.n959 B.n125 10.6151
R2861 B.n953 B.n125 10.6151
R2862 B.n953 B.n952 10.6151
R2863 B.n952 B.n951 10.6151
R2864 B.n951 B.n127 10.6151
R2865 B.n945 B.n127 10.6151
R2866 B.n943 B.n942 10.6151
R2867 B.n942 B.n131 10.6151
R2868 B.n936 B.n131 10.6151
R2869 B.n936 B.n935 10.6151
R2870 B.n935 B.n934 10.6151
R2871 B.n934 B.n133 10.6151
R2872 B.n928 B.n133 10.6151
R2873 B.n928 B.n927 10.6151
R2874 B.n927 B.n926 10.6151
R2875 B.n922 B.n921 10.6151
R2876 B.n921 B.n139 10.6151
R2877 B.n916 B.n139 10.6151
R2878 B.n916 B.n915 10.6151
R2879 B.n915 B.n914 10.6151
R2880 B.n914 B.n141 10.6151
R2881 B.n908 B.n141 10.6151
R2882 B.n908 B.n907 10.6151
R2883 B.n907 B.n906 10.6151
R2884 B.n906 B.n143 10.6151
R2885 B.n900 B.n143 10.6151
R2886 B.n900 B.n899 10.6151
R2887 B.n899 B.n898 10.6151
R2888 B.n898 B.n145 10.6151
R2889 B.n892 B.n145 10.6151
R2890 B.n892 B.n891 10.6151
R2891 B.n891 B.n890 10.6151
R2892 B.n890 B.n147 10.6151
R2893 B.n884 B.n147 10.6151
R2894 B.n884 B.n883 10.6151
R2895 B.n883 B.n882 10.6151
R2896 B.n882 B.n149 10.6151
R2897 B.n876 B.n149 10.6151
R2898 B.n876 B.n875 10.6151
R2899 B.n875 B.n874 10.6151
R2900 B.n874 B.n151 10.6151
R2901 B.n868 B.n151 10.6151
R2902 B.n868 B.n867 10.6151
R2903 B.n867 B.n866 10.6151
R2904 B.n866 B.n153 10.6151
R2905 B.n860 B.n153 10.6151
R2906 B.n860 B.n859 10.6151
R2907 B.n859 B.n858 10.6151
R2908 B.n858 B.n155 10.6151
R2909 B.n852 B.n155 10.6151
R2910 B.n852 B.n851 10.6151
R2911 B.n851 B.n850 10.6151
R2912 B.n850 B.n157 10.6151
R2913 B.n844 B.n157 10.6151
R2914 B.n844 B.n843 10.6151
R2915 B.n843 B.n842 10.6151
R2916 B.n842 B.n159 10.6151
R2917 B.n836 B.n159 10.6151
R2918 B.n836 B.n835 10.6151
R2919 B.n835 B.n834 10.6151
R2920 B.n834 B.n161 10.6151
R2921 B.n828 B.n161 10.6151
R2922 B.n828 B.n827 10.6151
R2923 B.n827 B.n826 10.6151
R2924 B.n826 B.n163 10.6151
R2925 B.n820 B.n163 10.6151
R2926 B.n820 B.n819 10.6151
R2927 B.n819 B.n818 10.6151
R2928 B.n818 B.n165 10.6151
R2929 B.n812 B.n165 10.6151
R2930 B.n585 B.n584 10.6151
R2931 B.n586 B.n585 10.6151
R2932 B.n586 B.n261 10.6151
R2933 B.n596 B.n261 10.6151
R2934 B.n597 B.n596 10.6151
R2935 B.n598 B.n597 10.6151
R2936 B.n598 B.n253 10.6151
R2937 B.n608 B.n253 10.6151
R2938 B.n609 B.n608 10.6151
R2939 B.n610 B.n609 10.6151
R2940 B.n610 B.n245 10.6151
R2941 B.n620 B.n245 10.6151
R2942 B.n621 B.n620 10.6151
R2943 B.n622 B.n621 10.6151
R2944 B.n622 B.n237 10.6151
R2945 B.n632 B.n237 10.6151
R2946 B.n633 B.n632 10.6151
R2947 B.n634 B.n633 10.6151
R2948 B.n634 B.n229 10.6151
R2949 B.n644 B.n229 10.6151
R2950 B.n645 B.n644 10.6151
R2951 B.n646 B.n645 10.6151
R2952 B.n646 B.n221 10.6151
R2953 B.n656 B.n221 10.6151
R2954 B.n657 B.n656 10.6151
R2955 B.n658 B.n657 10.6151
R2956 B.n658 B.n212 10.6151
R2957 B.n668 B.n212 10.6151
R2958 B.n669 B.n668 10.6151
R2959 B.n670 B.n669 10.6151
R2960 B.n670 B.n205 10.6151
R2961 B.n680 B.n205 10.6151
R2962 B.n681 B.n680 10.6151
R2963 B.n682 B.n681 10.6151
R2964 B.n682 B.n197 10.6151
R2965 B.n692 B.n197 10.6151
R2966 B.n693 B.n692 10.6151
R2967 B.n694 B.n693 10.6151
R2968 B.n694 B.n189 10.6151
R2969 B.n704 B.n189 10.6151
R2970 B.n705 B.n704 10.6151
R2971 B.n706 B.n705 10.6151
R2972 B.n706 B.n181 10.6151
R2973 B.n716 B.n181 10.6151
R2974 B.n717 B.n716 10.6151
R2975 B.n718 B.n717 10.6151
R2976 B.n718 B.n174 10.6151
R2977 B.n729 B.n174 10.6151
R2978 B.n730 B.n729 10.6151
R2979 B.n732 B.n730 10.6151
R2980 B.n732 B.n731 10.6151
R2981 B.n731 B.n166 10.6151
R2982 B.n743 B.n166 10.6151
R2983 B.n744 B.n743 10.6151
R2984 B.n745 B.n744 10.6151
R2985 B.n746 B.n745 10.6151
R2986 B.n748 B.n746 10.6151
R2987 B.n749 B.n748 10.6151
R2988 B.n750 B.n749 10.6151
R2989 B.n751 B.n750 10.6151
R2990 B.n753 B.n751 10.6151
R2991 B.n754 B.n753 10.6151
R2992 B.n755 B.n754 10.6151
R2993 B.n756 B.n755 10.6151
R2994 B.n758 B.n756 10.6151
R2995 B.n759 B.n758 10.6151
R2996 B.n760 B.n759 10.6151
R2997 B.n761 B.n760 10.6151
R2998 B.n763 B.n761 10.6151
R2999 B.n764 B.n763 10.6151
R3000 B.n765 B.n764 10.6151
R3001 B.n766 B.n765 10.6151
R3002 B.n768 B.n766 10.6151
R3003 B.n769 B.n768 10.6151
R3004 B.n770 B.n769 10.6151
R3005 B.n771 B.n770 10.6151
R3006 B.n773 B.n771 10.6151
R3007 B.n774 B.n773 10.6151
R3008 B.n775 B.n774 10.6151
R3009 B.n776 B.n775 10.6151
R3010 B.n778 B.n776 10.6151
R3011 B.n779 B.n778 10.6151
R3012 B.n780 B.n779 10.6151
R3013 B.n781 B.n780 10.6151
R3014 B.n783 B.n781 10.6151
R3015 B.n784 B.n783 10.6151
R3016 B.n785 B.n784 10.6151
R3017 B.n786 B.n785 10.6151
R3018 B.n788 B.n786 10.6151
R3019 B.n789 B.n788 10.6151
R3020 B.n790 B.n789 10.6151
R3021 B.n791 B.n790 10.6151
R3022 B.n793 B.n791 10.6151
R3023 B.n794 B.n793 10.6151
R3024 B.n795 B.n794 10.6151
R3025 B.n796 B.n795 10.6151
R3026 B.n798 B.n796 10.6151
R3027 B.n799 B.n798 10.6151
R3028 B.n800 B.n799 10.6151
R3029 B.n801 B.n800 10.6151
R3030 B.n803 B.n801 10.6151
R3031 B.n804 B.n803 10.6151
R3032 B.n805 B.n804 10.6151
R3033 B.n806 B.n805 10.6151
R3034 B.n808 B.n806 10.6151
R3035 B.n809 B.n808 10.6151
R3036 B.n810 B.n809 10.6151
R3037 B.n811 B.n810 10.6151
R3038 B.n579 B.n578 10.6151
R3039 B.n578 B.n273 10.6151
R3040 B.n573 B.n273 10.6151
R3041 B.n573 B.n572 10.6151
R3042 B.n572 B.n275 10.6151
R3043 B.n567 B.n275 10.6151
R3044 B.n567 B.n566 10.6151
R3045 B.n566 B.n565 10.6151
R3046 B.n565 B.n277 10.6151
R3047 B.n559 B.n277 10.6151
R3048 B.n559 B.n558 10.6151
R3049 B.n558 B.n557 10.6151
R3050 B.n557 B.n279 10.6151
R3051 B.n551 B.n279 10.6151
R3052 B.n551 B.n550 10.6151
R3053 B.n550 B.n549 10.6151
R3054 B.n549 B.n281 10.6151
R3055 B.n543 B.n281 10.6151
R3056 B.n543 B.n542 10.6151
R3057 B.n542 B.n541 10.6151
R3058 B.n541 B.n283 10.6151
R3059 B.n535 B.n283 10.6151
R3060 B.n535 B.n534 10.6151
R3061 B.n534 B.n533 10.6151
R3062 B.n533 B.n285 10.6151
R3063 B.n527 B.n285 10.6151
R3064 B.n527 B.n526 10.6151
R3065 B.n526 B.n525 10.6151
R3066 B.n525 B.n287 10.6151
R3067 B.n519 B.n287 10.6151
R3068 B.n519 B.n518 10.6151
R3069 B.n518 B.n517 10.6151
R3070 B.n517 B.n289 10.6151
R3071 B.n511 B.n289 10.6151
R3072 B.n511 B.n510 10.6151
R3073 B.n510 B.n509 10.6151
R3074 B.n509 B.n291 10.6151
R3075 B.n503 B.n291 10.6151
R3076 B.n503 B.n502 10.6151
R3077 B.n502 B.n501 10.6151
R3078 B.n501 B.n293 10.6151
R3079 B.n495 B.n293 10.6151
R3080 B.n495 B.n494 10.6151
R3081 B.n494 B.n493 10.6151
R3082 B.n493 B.n295 10.6151
R3083 B.n487 B.n295 10.6151
R3084 B.n487 B.n486 10.6151
R3085 B.n486 B.n485 10.6151
R3086 B.n485 B.n297 10.6151
R3087 B.n479 B.n297 10.6151
R3088 B.n479 B.n478 10.6151
R3089 B.n478 B.n477 10.6151
R3090 B.n477 B.n299 10.6151
R3091 B.n471 B.n299 10.6151
R3092 B.n471 B.n470 10.6151
R3093 B.n468 B.n303 10.6151
R3094 B.n462 B.n303 10.6151
R3095 B.n462 B.n461 10.6151
R3096 B.n461 B.n460 10.6151
R3097 B.n460 B.n305 10.6151
R3098 B.n454 B.n305 10.6151
R3099 B.n454 B.n453 10.6151
R3100 B.n453 B.n452 10.6151
R3101 B.n452 B.n307 10.6151
R3102 B.n446 B.n445 10.6151
R3103 B.n445 B.n444 10.6151
R3104 B.n444 B.n312 10.6151
R3105 B.n438 B.n312 10.6151
R3106 B.n438 B.n437 10.6151
R3107 B.n437 B.n436 10.6151
R3108 B.n436 B.n314 10.6151
R3109 B.n430 B.n314 10.6151
R3110 B.n430 B.n429 10.6151
R3111 B.n429 B.n428 10.6151
R3112 B.n428 B.n316 10.6151
R3113 B.n422 B.n316 10.6151
R3114 B.n422 B.n421 10.6151
R3115 B.n421 B.n420 10.6151
R3116 B.n420 B.n318 10.6151
R3117 B.n414 B.n318 10.6151
R3118 B.n414 B.n413 10.6151
R3119 B.n413 B.n412 10.6151
R3120 B.n412 B.n320 10.6151
R3121 B.n406 B.n320 10.6151
R3122 B.n406 B.n405 10.6151
R3123 B.n405 B.n404 10.6151
R3124 B.n404 B.n322 10.6151
R3125 B.n398 B.n322 10.6151
R3126 B.n398 B.n397 10.6151
R3127 B.n397 B.n396 10.6151
R3128 B.n396 B.n324 10.6151
R3129 B.n390 B.n324 10.6151
R3130 B.n390 B.n389 10.6151
R3131 B.n389 B.n388 10.6151
R3132 B.n388 B.n326 10.6151
R3133 B.n382 B.n326 10.6151
R3134 B.n382 B.n381 10.6151
R3135 B.n381 B.n380 10.6151
R3136 B.n380 B.n328 10.6151
R3137 B.n374 B.n328 10.6151
R3138 B.n374 B.n373 10.6151
R3139 B.n373 B.n372 10.6151
R3140 B.n372 B.n330 10.6151
R3141 B.n366 B.n330 10.6151
R3142 B.n366 B.n365 10.6151
R3143 B.n365 B.n364 10.6151
R3144 B.n364 B.n332 10.6151
R3145 B.n358 B.n332 10.6151
R3146 B.n358 B.n357 10.6151
R3147 B.n357 B.n356 10.6151
R3148 B.n356 B.n334 10.6151
R3149 B.n350 B.n334 10.6151
R3150 B.n350 B.n349 10.6151
R3151 B.n349 B.n348 10.6151
R3152 B.n348 B.n336 10.6151
R3153 B.n342 B.n336 10.6151
R3154 B.n342 B.n341 10.6151
R3155 B.n341 B.n340 10.6151
R3156 B.n340 B.n269 10.6151
R3157 B.n580 B.n265 10.6151
R3158 B.n590 B.n265 10.6151
R3159 B.n591 B.n590 10.6151
R3160 B.n592 B.n591 10.6151
R3161 B.n592 B.n257 10.6151
R3162 B.n602 B.n257 10.6151
R3163 B.n603 B.n602 10.6151
R3164 B.n604 B.n603 10.6151
R3165 B.n604 B.n249 10.6151
R3166 B.n614 B.n249 10.6151
R3167 B.n615 B.n614 10.6151
R3168 B.n616 B.n615 10.6151
R3169 B.n616 B.n241 10.6151
R3170 B.n626 B.n241 10.6151
R3171 B.n627 B.n626 10.6151
R3172 B.n628 B.n627 10.6151
R3173 B.n628 B.n233 10.6151
R3174 B.n638 B.n233 10.6151
R3175 B.n639 B.n638 10.6151
R3176 B.n640 B.n639 10.6151
R3177 B.n640 B.n225 10.6151
R3178 B.n650 B.n225 10.6151
R3179 B.n651 B.n650 10.6151
R3180 B.n652 B.n651 10.6151
R3181 B.n652 B.n217 10.6151
R3182 B.n662 B.n217 10.6151
R3183 B.n663 B.n662 10.6151
R3184 B.n664 B.n663 10.6151
R3185 B.n664 B.n209 10.6151
R3186 B.n674 B.n209 10.6151
R3187 B.n675 B.n674 10.6151
R3188 B.n676 B.n675 10.6151
R3189 B.n676 B.n201 10.6151
R3190 B.n686 B.n201 10.6151
R3191 B.n687 B.n686 10.6151
R3192 B.n688 B.n687 10.6151
R3193 B.n688 B.n193 10.6151
R3194 B.n698 B.n193 10.6151
R3195 B.n699 B.n698 10.6151
R3196 B.n700 B.n699 10.6151
R3197 B.n700 B.n185 10.6151
R3198 B.n710 B.n185 10.6151
R3199 B.n711 B.n710 10.6151
R3200 B.n712 B.n711 10.6151
R3201 B.n712 B.n177 10.6151
R3202 B.n723 B.n177 10.6151
R3203 B.n724 B.n723 10.6151
R3204 B.n725 B.n724 10.6151
R3205 B.n725 B.n170 10.6151
R3206 B.n736 B.n170 10.6151
R3207 B.n737 B.n736 10.6151
R3208 B.n738 B.n737 10.6151
R3209 B.n738 B.n0 10.6151
R3210 B.n1161 B.n1 10.6151
R3211 B.n1161 B.n1160 10.6151
R3212 B.n1160 B.n1159 10.6151
R3213 B.n1159 B.n10 10.6151
R3214 B.n1153 B.n10 10.6151
R3215 B.n1153 B.n1152 10.6151
R3216 B.n1152 B.n1151 10.6151
R3217 B.n1151 B.n16 10.6151
R3218 B.n1145 B.n16 10.6151
R3219 B.n1145 B.n1144 10.6151
R3220 B.n1144 B.n1143 10.6151
R3221 B.n1143 B.n24 10.6151
R3222 B.n1137 B.n24 10.6151
R3223 B.n1137 B.n1136 10.6151
R3224 B.n1136 B.n1135 10.6151
R3225 B.n1135 B.n31 10.6151
R3226 B.n1129 B.n31 10.6151
R3227 B.n1129 B.n1128 10.6151
R3228 B.n1128 B.n1127 10.6151
R3229 B.n1127 B.n38 10.6151
R3230 B.n1121 B.n38 10.6151
R3231 B.n1121 B.n1120 10.6151
R3232 B.n1120 B.n1119 10.6151
R3233 B.n1119 B.n45 10.6151
R3234 B.n1113 B.n45 10.6151
R3235 B.n1113 B.n1112 10.6151
R3236 B.n1112 B.n1111 10.6151
R3237 B.n1111 B.n52 10.6151
R3238 B.n1105 B.n52 10.6151
R3239 B.n1105 B.n1104 10.6151
R3240 B.n1104 B.n1103 10.6151
R3241 B.n1103 B.n59 10.6151
R3242 B.n1097 B.n59 10.6151
R3243 B.n1097 B.n1096 10.6151
R3244 B.n1096 B.n1095 10.6151
R3245 B.n1095 B.n66 10.6151
R3246 B.n1089 B.n66 10.6151
R3247 B.n1089 B.n1088 10.6151
R3248 B.n1088 B.n1087 10.6151
R3249 B.n1087 B.n73 10.6151
R3250 B.n1081 B.n73 10.6151
R3251 B.n1081 B.n1080 10.6151
R3252 B.n1080 B.n1079 10.6151
R3253 B.n1079 B.n80 10.6151
R3254 B.n1073 B.n80 10.6151
R3255 B.n1073 B.n1072 10.6151
R3256 B.n1072 B.n1071 10.6151
R3257 B.n1071 B.n87 10.6151
R3258 B.n1065 B.n87 10.6151
R3259 B.n1065 B.n1064 10.6151
R3260 B.n1064 B.n1063 10.6151
R3261 B.n1063 B.n94 10.6151
R3262 B.n1057 B.n94 10.6151
R3263 B.n945 B.n944 9.36635
R3264 B.n922 B.n137 9.36635
R3265 B.n470 B.n469 9.36635
R3266 B.n446 B.n311 9.36635
R3267 B.n727 B.t7 5.93175
R3268 B.n1155 B.t5 5.93175
R3269 B.n1167 B.n0 2.81026
R3270 B.n1167 B.n1 2.81026
R3271 B.n944 B.n943 1.24928
R3272 B.n926 B.n137 1.24928
R3273 B.n469 B.n468 1.24928
R3274 B.n311 B.n307 1.24928
R3275 B.n606 B.t9 0.989042
R3276 B.t13 B.n1075 0.989042
R3277 VN.n8 VN.t1 180.248
R3278 VN.n39 VN.t3 180.248
R3279 VN.n59 VN.n31 161.3
R3280 VN.n58 VN.n57 161.3
R3281 VN.n56 VN.n32 161.3
R3282 VN.n55 VN.n54 161.3
R3283 VN.n53 VN.n33 161.3
R3284 VN.n52 VN.n51 161.3
R3285 VN.n50 VN.n49 161.3
R3286 VN.n48 VN.n35 161.3
R3287 VN.n47 VN.n46 161.3
R3288 VN.n45 VN.n36 161.3
R3289 VN.n44 VN.n43 161.3
R3290 VN.n42 VN.n37 161.3
R3291 VN.n41 VN.n40 161.3
R3292 VN.n28 VN.n0 161.3
R3293 VN.n27 VN.n26 161.3
R3294 VN.n25 VN.n1 161.3
R3295 VN.n24 VN.n23 161.3
R3296 VN.n22 VN.n2 161.3
R3297 VN.n21 VN.n20 161.3
R3298 VN.n19 VN.n18 161.3
R3299 VN.n17 VN.n4 161.3
R3300 VN.n16 VN.n15 161.3
R3301 VN.n14 VN.n5 161.3
R3302 VN.n13 VN.n12 161.3
R3303 VN.n11 VN.n6 161.3
R3304 VN.n10 VN.n9 161.3
R3305 VN.n7 VN.t7 147.202
R3306 VN.n3 VN.t0 147.202
R3307 VN.n29 VN.t2 147.202
R3308 VN.n38 VN.t4 147.202
R3309 VN.n34 VN.t5 147.202
R3310 VN.n60 VN.t6 147.202
R3311 VN.n30 VN.n29 102.793
R3312 VN.n61 VN.n60 102.793
R3313 VN.n8 VN.n7 70.4561
R3314 VN.n39 VN.n38 70.4561
R3315 VN VN.n61 55.8239
R3316 VN.n23 VN.n1 51.2335
R3317 VN.n54 VN.n32 51.2335
R3318 VN.n12 VN.n5 40.577
R3319 VN.n16 VN.n5 40.577
R3320 VN.n43 VN.n36 40.577
R3321 VN.n47 VN.n36 40.577
R3322 VN.n23 VN.n22 29.9206
R3323 VN.n54 VN.n53 29.9206
R3324 VN.n11 VN.n10 24.5923
R3325 VN.n12 VN.n11 24.5923
R3326 VN.n17 VN.n16 24.5923
R3327 VN.n18 VN.n17 24.5923
R3328 VN.n22 VN.n21 24.5923
R3329 VN.n27 VN.n1 24.5923
R3330 VN.n28 VN.n27 24.5923
R3331 VN.n43 VN.n42 24.5923
R3332 VN.n42 VN.n41 24.5923
R3333 VN.n53 VN.n52 24.5923
R3334 VN.n49 VN.n48 24.5923
R3335 VN.n48 VN.n47 24.5923
R3336 VN.n59 VN.n58 24.5923
R3337 VN.n58 VN.n32 24.5923
R3338 VN.n21 VN.n3 21.8872
R3339 VN.n52 VN.n34 21.8872
R3340 VN.n29 VN.n28 8.11581
R3341 VN.n60 VN.n59 8.11581
R3342 VN.n40 VN.n39 6.95301
R3343 VN.n9 VN.n8 6.95301
R3344 VN.n10 VN.n7 2.7056
R3345 VN.n18 VN.n3 2.7056
R3346 VN.n41 VN.n38 2.7056
R3347 VN.n49 VN.n34 2.7056
R3348 VN.n61 VN.n31 0.278335
R3349 VN.n30 VN.n0 0.278335
R3350 VN.n57 VN.n31 0.189894
R3351 VN.n57 VN.n56 0.189894
R3352 VN.n56 VN.n55 0.189894
R3353 VN.n55 VN.n33 0.189894
R3354 VN.n51 VN.n33 0.189894
R3355 VN.n51 VN.n50 0.189894
R3356 VN.n50 VN.n35 0.189894
R3357 VN.n46 VN.n35 0.189894
R3358 VN.n46 VN.n45 0.189894
R3359 VN.n45 VN.n44 0.189894
R3360 VN.n44 VN.n37 0.189894
R3361 VN.n40 VN.n37 0.189894
R3362 VN.n9 VN.n6 0.189894
R3363 VN.n13 VN.n6 0.189894
R3364 VN.n14 VN.n13 0.189894
R3365 VN.n15 VN.n14 0.189894
R3366 VN.n15 VN.n4 0.189894
R3367 VN.n19 VN.n4 0.189894
R3368 VN.n20 VN.n19 0.189894
R3369 VN.n20 VN.n2 0.189894
R3370 VN.n24 VN.n2 0.189894
R3371 VN.n25 VN.n24 0.189894
R3372 VN.n26 VN.n25 0.189894
R3373 VN.n26 VN.n0 0.189894
R3374 VN VN.n30 0.153485
R3375 VDD2.n2 VDD2.n1 65.5007
R3376 VDD2.n2 VDD2.n0 65.5007
R3377 VDD2 VDD2.n5 65.4979
R3378 VDD2.n4 VDD2.n3 64.2157
R3379 VDD2.n4 VDD2.n2 50.4179
R3380 VDD2 VDD2.n4 1.39921
R3381 VDD2.n5 VDD2.t3 1.16658
R3382 VDD2.n5 VDD2.t4 1.16658
R3383 VDD2.n3 VDD2.t1 1.16658
R3384 VDD2.n3 VDD2.t2 1.16658
R3385 VDD2.n1 VDD2.t7 1.16658
R3386 VDD2.n1 VDD2.t5 1.16658
R3387 VDD2.n0 VDD2.t6 1.16658
R3388 VDD2.n0 VDD2.t0 1.16658
C0 VDD1 VDD2 1.87042f
C1 VN VTAIL 12.5081f
C2 VN VP 8.796009f
C3 VTAIL VP 12.522201f
C4 VN VDD1 0.152286f
C5 VN VDD2 12.2731f
C6 VTAIL VDD1 9.73595f
C7 VDD1 VP 12.6584f
C8 VTAIL VDD2 9.79158f
C9 VDD2 VP 0.539058f
C10 VDD2 B 5.898353f
C11 VDD1 B 6.351901f
C12 VTAIL B 13.593126f
C13 VN B 16.590368f
C14 VP B 15.118764f
C15 VDD2.t6 B 0.32599f
C16 VDD2.t0 B 0.32599f
C17 VDD2.n0 B 2.97657f
C18 VDD2.t7 B 0.32599f
C19 VDD2.t5 B 0.32599f
C20 VDD2.n1 B 2.97657f
C21 VDD2.n2 B 3.58782f
C22 VDD2.t1 B 0.32599f
C23 VDD2.t2 B 0.32599f
C24 VDD2.n3 B 2.96642f
C25 VDD2.n4 B 3.2911f
C26 VDD2.t3 B 0.32599f
C27 VDD2.t4 B 0.32599f
C28 VDD2.n5 B 2.97653f
C29 VN.n0 B 0.026874f
C30 VN.t2 B 2.64378f
C31 VN.n1 B 0.036832f
C32 VN.n2 B 0.020385f
C33 VN.t0 B 2.64378f
C34 VN.n3 B 0.917568f
C35 VN.n4 B 0.020385f
C36 VN.n5 B 0.016464f
C37 VN.n6 B 0.020385f
C38 VN.t7 B 2.64378f
C39 VN.n7 B 0.972033f
C40 VN.t1 B 2.83599f
C41 VN.n8 B 0.949346f
C42 VN.n9 B 0.200804f
C43 VN.n10 B 0.021193f
C44 VN.n11 B 0.037802f
C45 VN.n12 B 0.040302f
C46 VN.n13 B 0.020385f
C47 VN.n14 B 0.020385f
C48 VN.n15 B 0.020385f
C49 VN.n16 B 0.040302f
C50 VN.n17 B 0.037802f
C51 VN.n18 B 0.021193f
C52 VN.n19 B 0.020385f
C53 VN.n20 B 0.020385f
C54 VN.n21 B 0.035749f
C55 VN.n22 B 0.040394f
C56 VN.n23 B 0.019842f
C57 VN.n24 B 0.020385f
C58 VN.n25 B 0.020385f
C59 VN.n26 B 0.020385f
C60 VN.n27 B 0.037802f
C61 VN.n28 B 0.025299f
C62 VN.n29 B 0.988272f
C63 VN.n30 B 0.035351f
C64 VN.n31 B 0.026874f
C65 VN.t6 B 2.64378f
C66 VN.n32 B 0.036832f
C67 VN.n33 B 0.020385f
C68 VN.t5 B 2.64378f
C69 VN.n34 B 0.917568f
C70 VN.n35 B 0.020385f
C71 VN.n36 B 0.016464f
C72 VN.n37 B 0.020385f
C73 VN.t4 B 2.64378f
C74 VN.n38 B 0.972033f
C75 VN.t3 B 2.83599f
C76 VN.n39 B 0.949346f
C77 VN.n40 B 0.200804f
C78 VN.n41 B 0.021193f
C79 VN.n42 B 0.037802f
C80 VN.n43 B 0.040302f
C81 VN.n44 B 0.020385f
C82 VN.n45 B 0.020385f
C83 VN.n46 B 0.020385f
C84 VN.n47 B 0.040302f
C85 VN.n48 B 0.037802f
C86 VN.n49 B 0.021193f
C87 VN.n50 B 0.020385f
C88 VN.n51 B 0.020385f
C89 VN.n52 B 0.035749f
C90 VN.n53 B 0.040394f
C91 VN.n54 B 0.019842f
C92 VN.n55 B 0.020385f
C93 VN.n56 B 0.020385f
C94 VN.n57 B 0.020385f
C95 VN.n58 B 0.037802f
C96 VN.n59 B 0.025299f
C97 VN.n60 B 0.988272f
C98 VN.n61 B 1.3324f
C99 VDD1.t2 B 0.329079f
C100 VDD1.t5 B 0.329079f
C101 VDD1.n0 B 3.00585f
C102 VDD1.t3 B 0.329079f
C103 VDD1.t7 B 0.329079f
C104 VDD1.n1 B 3.00478f
C105 VDD1.t1 B 0.329079f
C106 VDD1.t4 B 0.329079f
C107 VDD1.n2 B 3.00478f
C108 VDD1.n3 B 3.6726f
C109 VDD1.t6 B 0.329079f
C110 VDD1.t0 B 0.329079f
C111 VDD1.n4 B 2.99452f
C112 VDD1.n5 B 3.3529f
C113 VTAIL.t6 B 0.252128f
C114 VTAIL.t0 B 0.252128f
C115 VTAIL.n0 B 2.24201f
C116 VTAIL.n1 B 0.345149f
C117 VTAIL.n2 B 0.027679f
C118 VTAIL.n3 B 0.01879f
C119 VTAIL.n4 B 0.010097f
C120 VTAIL.n5 B 0.023866f
C121 VTAIL.n6 B 0.010691f
C122 VTAIL.n7 B 0.01879f
C123 VTAIL.n8 B 0.010097f
C124 VTAIL.n9 B 0.023866f
C125 VTAIL.n10 B 0.010691f
C126 VTAIL.n11 B 0.01879f
C127 VTAIL.n12 B 0.010097f
C128 VTAIL.n13 B 0.023866f
C129 VTAIL.n14 B 0.010691f
C130 VTAIL.n15 B 0.01879f
C131 VTAIL.n16 B 0.010097f
C132 VTAIL.n17 B 0.023866f
C133 VTAIL.n18 B 0.010691f
C134 VTAIL.n19 B 0.01879f
C135 VTAIL.n20 B 0.010097f
C136 VTAIL.n21 B 0.023866f
C137 VTAIL.n22 B 0.010691f
C138 VTAIL.n23 B 0.01879f
C139 VTAIL.n24 B 0.010097f
C140 VTAIL.n25 B 0.023866f
C141 VTAIL.n26 B 0.010691f
C142 VTAIL.n27 B 0.01879f
C143 VTAIL.n28 B 0.010097f
C144 VTAIL.n29 B 0.023866f
C145 VTAIL.n30 B 0.010691f
C146 VTAIL.n31 B 0.131881f
C147 VTAIL.t5 B 0.039479f
C148 VTAIL.n32 B 0.017899f
C149 VTAIL.n33 B 0.014098f
C150 VTAIL.n34 B 0.010097f
C151 VTAIL.n35 B 1.39302f
C152 VTAIL.n36 B 0.01879f
C153 VTAIL.n37 B 0.010097f
C154 VTAIL.n38 B 0.010691f
C155 VTAIL.n39 B 0.023866f
C156 VTAIL.n40 B 0.023866f
C157 VTAIL.n41 B 0.010691f
C158 VTAIL.n42 B 0.010097f
C159 VTAIL.n43 B 0.01879f
C160 VTAIL.n44 B 0.01879f
C161 VTAIL.n45 B 0.010097f
C162 VTAIL.n46 B 0.010691f
C163 VTAIL.n47 B 0.023866f
C164 VTAIL.n48 B 0.023866f
C165 VTAIL.n49 B 0.010691f
C166 VTAIL.n50 B 0.010097f
C167 VTAIL.n51 B 0.01879f
C168 VTAIL.n52 B 0.01879f
C169 VTAIL.n53 B 0.010097f
C170 VTAIL.n54 B 0.010691f
C171 VTAIL.n55 B 0.023866f
C172 VTAIL.n56 B 0.023866f
C173 VTAIL.n57 B 0.010691f
C174 VTAIL.n58 B 0.010097f
C175 VTAIL.n59 B 0.01879f
C176 VTAIL.n60 B 0.01879f
C177 VTAIL.n61 B 0.010097f
C178 VTAIL.n62 B 0.010691f
C179 VTAIL.n63 B 0.023866f
C180 VTAIL.n64 B 0.023866f
C181 VTAIL.n65 B 0.010691f
C182 VTAIL.n66 B 0.010097f
C183 VTAIL.n67 B 0.01879f
C184 VTAIL.n68 B 0.01879f
C185 VTAIL.n69 B 0.010097f
C186 VTAIL.n70 B 0.010691f
C187 VTAIL.n71 B 0.023866f
C188 VTAIL.n72 B 0.023866f
C189 VTAIL.n73 B 0.023866f
C190 VTAIL.n74 B 0.010691f
C191 VTAIL.n75 B 0.010097f
C192 VTAIL.n76 B 0.01879f
C193 VTAIL.n77 B 0.01879f
C194 VTAIL.n78 B 0.010097f
C195 VTAIL.n79 B 0.010394f
C196 VTAIL.n80 B 0.010394f
C197 VTAIL.n81 B 0.023866f
C198 VTAIL.n82 B 0.023866f
C199 VTAIL.n83 B 0.010691f
C200 VTAIL.n84 B 0.010097f
C201 VTAIL.n85 B 0.01879f
C202 VTAIL.n86 B 0.01879f
C203 VTAIL.n87 B 0.010097f
C204 VTAIL.n88 B 0.010691f
C205 VTAIL.n89 B 0.023866f
C206 VTAIL.n90 B 0.053907f
C207 VTAIL.n91 B 0.010691f
C208 VTAIL.n92 B 0.010097f
C209 VTAIL.n93 B 0.048053f
C210 VTAIL.n94 B 0.030529f
C211 VTAIL.n95 B 0.209434f
C212 VTAIL.n96 B 0.027679f
C213 VTAIL.n97 B 0.01879f
C214 VTAIL.n98 B 0.010097f
C215 VTAIL.n99 B 0.023866f
C216 VTAIL.n100 B 0.010691f
C217 VTAIL.n101 B 0.01879f
C218 VTAIL.n102 B 0.010097f
C219 VTAIL.n103 B 0.023866f
C220 VTAIL.n104 B 0.010691f
C221 VTAIL.n105 B 0.01879f
C222 VTAIL.n106 B 0.010097f
C223 VTAIL.n107 B 0.023866f
C224 VTAIL.n108 B 0.010691f
C225 VTAIL.n109 B 0.01879f
C226 VTAIL.n110 B 0.010097f
C227 VTAIL.n111 B 0.023866f
C228 VTAIL.n112 B 0.010691f
C229 VTAIL.n113 B 0.01879f
C230 VTAIL.n114 B 0.010097f
C231 VTAIL.n115 B 0.023866f
C232 VTAIL.n116 B 0.010691f
C233 VTAIL.n117 B 0.01879f
C234 VTAIL.n118 B 0.010097f
C235 VTAIL.n119 B 0.023866f
C236 VTAIL.n120 B 0.010691f
C237 VTAIL.n121 B 0.01879f
C238 VTAIL.n122 B 0.010097f
C239 VTAIL.n123 B 0.023866f
C240 VTAIL.n124 B 0.010691f
C241 VTAIL.n125 B 0.131881f
C242 VTAIL.t10 B 0.039479f
C243 VTAIL.n126 B 0.017899f
C244 VTAIL.n127 B 0.014098f
C245 VTAIL.n128 B 0.010097f
C246 VTAIL.n129 B 1.39302f
C247 VTAIL.n130 B 0.01879f
C248 VTAIL.n131 B 0.010097f
C249 VTAIL.n132 B 0.010691f
C250 VTAIL.n133 B 0.023866f
C251 VTAIL.n134 B 0.023866f
C252 VTAIL.n135 B 0.010691f
C253 VTAIL.n136 B 0.010097f
C254 VTAIL.n137 B 0.01879f
C255 VTAIL.n138 B 0.01879f
C256 VTAIL.n139 B 0.010097f
C257 VTAIL.n140 B 0.010691f
C258 VTAIL.n141 B 0.023866f
C259 VTAIL.n142 B 0.023866f
C260 VTAIL.n143 B 0.010691f
C261 VTAIL.n144 B 0.010097f
C262 VTAIL.n145 B 0.01879f
C263 VTAIL.n146 B 0.01879f
C264 VTAIL.n147 B 0.010097f
C265 VTAIL.n148 B 0.010691f
C266 VTAIL.n149 B 0.023866f
C267 VTAIL.n150 B 0.023866f
C268 VTAIL.n151 B 0.010691f
C269 VTAIL.n152 B 0.010097f
C270 VTAIL.n153 B 0.01879f
C271 VTAIL.n154 B 0.01879f
C272 VTAIL.n155 B 0.010097f
C273 VTAIL.n156 B 0.010691f
C274 VTAIL.n157 B 0.023866f
C275 VTAIL.n158 B 0.023866f
C276 VTAIL.n159 B 0.010691f
C277 VTAIL.n160 B 0.010097f
C278 VTAIL.n161 B 0.01879f
C279 VTAIL.n162 B 0.01879f
C280 VTAIL.n163 B 0.010097f
C281 VTAIL.n164 B 0.010691f
C282 VTAIL.n165 B 0.023866f
C283 VTAIL.n166 B 0.023866f
C284 VTAIL.n167 B 0.023866f
C285 VTAIL.n168 B 0.010691f
C286 VTAIL.n169 B 0.010097f
C287 VTAIL.n170 B 0.01879f
C288 VTAIL.n171 B 0.01879f
C289 VTAIL.n172 B 0.010097f
C290 VTAIL.n173 B 0.010394f
C291 VTAIL.n174 B 0.010394f
C292 VTAIL.n175 B 0.023866f
C293 VTAIL.n176 B 0.023866f
C294 VTAIL.n177 B 0.010691f
C295 VTAIL.n178 B 0.010097f
C296 VTAIL.n179 B 0.01879f
C297 VTAIL.n180 B 0.01879f
C298 VTAIL.n181 B 0.010097f
C299 VTAIL.n182 B 0.010691f
C300 VTAIL.n183 B 0.023866f
C301 VTAIL.n184 B 0.053907f
C302 VTAIL.n185 B 0.010691f
C303 VTAIL.n186 B 0.010097f
C304 VTAIL.n187 B 0.048053f
C305 VTAIL.n188 B 0.030529f
C306 VTAIL.n189 B 0.209434f
C307 VTAIL.t9 B 0.252128f
C308 VTAIL.t13 B 0.252128f
C309 VTAIL.n190 B 2.24201f
C310 VTAIL.n191 B 0.503951f
C311 VTAIL.n192 B 0.027679f
C312 VTAIL.n193 B 0.01879f
C313 VTAIL.n194 B 0.010097f
C314 VTAIL.n195 B 0.023866f
C315 VTAIL.n196 B 0.010691f
C316 VTAIL.n197 B 0.01879f
C317 VTAIL.n198 B 0.010097f
C318 VTAIL.n199 B 0.023866f
C319 VTAIL.n200 B 0.010691f
C320 VTAIL.n201 B 0.01879f
C321 VTAIL.n202 B 0.010097f
C322 VTAIL.n203 B 0.023866f
C323 VTAIL.n204 B 0.010691f
C324 VTAIL.n205 B 0.01879f
C325 VTAIL.n206 B 0.010097f
C326 VTAIL.n207 B 0.023866f
C327 VTAIL.n208 B 0.010691f
C328 VTAIL.n209 B 0.01879f
C329 VTAIL.n210 B 0.010097f
C330 VTAIL.n211 B 0.023866f
C331 VTAIL.n212 B 0.010691f
C332 VTAIL.n213 B 0.01879f
C333 VTAIL.n214 B 0.010097f
C334 VTAIL.n215 B 0.023866f
C335 VTAIL.n216 B 0.010691f
C336 VTAIL.n217 B 0.01879f
C337 VTAIL.n218 B 0.010097f
C338 VTAIL.n219 B 0.023866f
C339 VTAIL.n220 B 0.010691f
C340 VTAIL.n221 B 0.131881f
C341 VTAIL.t12 B 0.039479f
C342 VTAIL.n222 B 0.017899f
C343 VTAIL.n223 B 0.014098f
C344 VTAIL.n224 B 0.010097f
C345 VTAIL.n225 B 1.39302f
C346 VTAIL.n226 B 0.01879f
C347 VTAIL.n227 B 0.010097f
C348 VTAIL.n228 B 0.010691f
C349 VTAIL.n229 B 0.023866f
C350 VTAIL.n230 B 0.023866f
C351 VTAIL.n231 B 0.010691f
C352 VTAIL.n232 B 0.010097f
C353 VTAIL.n233 B 0.01879f
C354 VTAIL.n234 B 0.01879f
C355 VTAIL.n235 B 0.010097f
C356 VTAIL.n236 B 0.010691f
C357 VTAIL.n237 B 0.023866f
C358 VTAIL.n238 B 0.023866f
C359 VTAIL.n239 B 0.010691f
C360 VTAIL.n240 B 0.010097f
C361 VTAIL.n241 B 0.01879f
C362 VTAIL.n242 B 0.01879f
C363 VTAIL.n243 B 0.010097f
C364 VTAIL.n244 B 0.010691f
C365 VTAIL.n245 B 0.023866f
C366 VTAIL.n246 B 0.023866f
C367 VTAIL.n247 B 0.010691f
C368 VTAIL.n248 B 0.010097f
C369 VTAIL.n249 B 0.01879f
C370 VTAIL.n250 B 0.01879f
C371 VTAIL.n251 B 0.010097f
C372 VTAIL.n252 B 0.010691f
C373 VTAIL.n253 B 0.023866f
C374 VTAIL.n254 B 0.023866f
C375 VTAIL.n255 B 0.010691f
C376 VTAIL.n256 B 0.010097f
C377 VTAIL.n257 B 0.01879f
C378 VTAIL.n258 B 0.01879f
C379 VTAIL.n259 B 0.010097f
C380 VTAIL.n260 B 0.010691f
C381 VTAIL.n261 B 0.023866f
C382 VTAIL.n262 B 0.023866f
C383 VTAIL.n263 B 0.023866f
C384 VTAIL.n264 B 0.010691f
C385 VTAIL.n265 B 0.010097f
C386 VTAIL.n266 B 0.01879f
C387 VTAIL.n267 B 0.01879f
C388 VTAIL.n268 B 0.010097f
C389 VTAIL.n269 B 0.010394f
C390 VTAIL.n270 B 0.010394f
C391 VTAIL.n271 B 0.023866f
C392 VTAIL.n272 B 0.023866f
C393 VTAIL.n273 B 0.010691f
C394 VTAIL.n274 B 0.010097f
C395 VTAIL.n275 B 0.01879f
C396 VTAIL.n276 B 0.01879f
C397 VTAIL.n277 B 0.010097f
C398 VTAIL.n278 B 0.010691f
C399 VTAIL.n279 B 0.023866f
C400 VTAIL.n280 B 0.053907f
C401 VTAIL.n281 B 0.010691f
C402 VTAIL.n282 B 0.010097f
C403 VTAIL.n283 B 0.048053f
C404 VTAIL.n284 B 0.030529f
C405 VTAIL.n285 B 1.48482f
C406 VTAIL.n286 B 0.027679f
C407 VTAIL.n287 B 0.01879f
C408 VTAIL.n288 B 0.010097f
C409 VTAIL.n289 B 0.023866f
C410 VTAIL.n290 B 0.010691f
C411 VTAIL.n291 B 0.01879f
C412 VTAIL.n292 B 0.010097f
C413 VTAIL.n293 B 0.023866f
C414 VTAIL.n294 B 0.010691f
C415 VTAIL.n295 B 0.01879f
C416 VTAIL.n296 B 0.010097f
C417 VTAIL.n297 B 0.023866f
C418 VTAIL.n298 B 0.023866f
C419 VTAIL.n299 B 0.010691f
C420 VTAIL.n300 B 0.01879f
C421 VTAIL.n301 B 0.010097f
C422 VTAIL.n302 B 0.023866f
C423 VTAIL.n303 B 0.010691f
C424 VTAIL.n304 B 0.01879f
C425 VTAIL.n305 B 0.010097f
C426 VTAIL.n306 B 0.023866f
C427 VTAIL.n307 B 0.010691f
C428 VTAIL.n308 B 0.01879f
C429 VTAIL.n309 B 0.010097f
C430 VTAIL.n310 B 0.023866f
C431 VTAIL.n311 B 0.010691f
C432 VTAIL.n312 B 0.01879f
C433 VTAIL.n313 B 0.010097f
C434 VTAIL.n314 B 0.023866f
C435 VTAIL.n315 B 0.010691f
C436 VTAIL.n316 B 0.131881f
C437 VTAIL.t4 B 0.039479f
C438 VTAIL.n317 B 0.017899f
C439 VTAIL.n318 B 0.014098f
C440 VTAIL.n319 B 0.010097f
C441 VTAIL.n320 B 1.39302f
C442 VTAIL.n321 B 0.01879f
C443 VTAIL.n322 B 0.010097f
C444 VTAIL.n323 B 0.010691f
C445 VTAIL.n324 B 0.023866f
C446 VTAIL.n325 B 0.023866f
C447 VTAIL.n326 B 0.010691f
C448 VTAIL.n327 B 0.010097f
C449 VTAIL.n328 B 0.01879f
C450 VTAIL.n329 B 0.01879f
C451 VTAIL.n330 B 0.010097f
C452 VTAIL.n331 B 0.010691f
C453 VTAIL.n332 B 0.023866f
C454 VTAIL.n333 B 0.023866f
C455 VTAIL.n334 B 0.010691f
C456 VTAIL.n335 B 0.010097f
C457 VTAIL.n336 B 0.01879f
C458 VTAIL.n337 B 0.01879f
C459 VTAIL.n338 B 0.010097f
C460 VTAIL.n339 B 0.010691f
C461 VTAIL.n340 B 0.023866f
C462 VTAIL.n341 B 0.023866f
C463 VTAIL.n342 B 0.010691f
C464 VTAIL.n343 B 0.010097f
C465 VTAIL.n344 B 0.01879f
C466 VTAIL.n345 B 0.01879f
C467 VTAIL.n346 B 0.010097f
C468 VTAIL.n347 B 0.010691f
C469 VTAIL.n348 B 0.023866f
C470 VTAIL.n349 B 0.023866f
C471 VTAIL.n350 B 0.010691f
C472 VTAIL.n351 B 0.010097f
C473 VTAIL.n352 B 0.01879f
C474 VTAIL.n353 B 0.01879f
C475 VTAIL.n354 B 0.010097f
C476 VTAIL.n355 B 0.010691f
C477 VTAIL.n356 B 0.023866f
C478 VTAIL.n357 B 0.023866f
C479 VTAIL.n358 B 0.010691f
C480 VTAIL.n359 B 0.010097f
C481 VTAIL.n360 B 0.01879f
C482 VTAIL.n361 B 0.01879f
C483 VTAIL.n362 B 0.010097f
C484 VTAIL.n363 B 0.010394f
C485 VTAIL.n364 B 0.010394f
C486 VTAIL.n365 B 0.023866f
C487 VTAIL.n366 B 0.023866f
C488 VTAIL.n367 B 0.010691f
C489 VTAIL.n368 B 0.010097f
C490 VTAIL.n369 B 0.01879f
C491 VTAIL.n370 B 0.01879f
C492 VTAIL.n371 B 0.010097f
C493 VTAIL.n372 B 0.010691f
C494 VTAIL.n373 B 0.023866f
C495 VTAIL.n374 B 0.053907f
C496 VTAIL.n375 B 0.010691f
C497 VTAIL.n376 B 0.010097f
C498 VTAIL.n377 B 0.048053f
C499 VTAIL.n378 B 0.030529f
C500 VTAIL.n379 B 1.48482f
C501 VTAIL.t1 B 0.252128f
C502 VTAIL.t3 B 0.252128f
C503 VTAIL.n380 B 2.24202f
C504 VTAIL.n381 B 0.503942f
C505 VTAIL.n382 B 0.027679f
C506 VTAIL.n383 B 0.01879f
C507 VTAIL.n384 B 0.010097f
C508 VTAIL.n385 B 0.023866f
C509 VTAIL.n386 B 0.010691f
C510 VTAIL.n387 B 0.01879f
C511 VTAIL.n388 B 0.010097f
C512 VTAIL.n389 B 0.023866f
C513 VTAIL.n390 B 0.010691f
C514 VTAIL.n391 B 0.01879f
C515 VTAIL.n392 B 0.010097f
C516 VTAIL.n393 B 0.023866f
C517 VTAIL.n394 B 0.023866f
C518 VTAIL.n395 B 0.010691f
C519 VTAIL.n396 B 0.01879f
C520 VTAIL.n397 B 0.010097f
C521 VTAIL.n398 B 0.023866f
C522 VTAIL.n399 B 0.010691f
C523 VTAIL.n400 B 0.01879f
C524 VTAIL.n401 B 0.010097f
C525 VTAIL.n402 B 0.023866f
C526 VTAIL.n403 B 0.010691f
C527 VTAIL.n404 B 0.01879f
C528 VTAIL.n405 B 0.010097f
C529 VTAIL.n406 B 0.023866f
C530 VTAIL.n407 B 0.010691f
C531 VTAIL.n408 B 0.01879f
C532 VTAIL.n409 B 0.010097f
C533 VTAIL.n410 B 0.023866f
C534 VTAIL.n411 B 0.010691f
C535 VTAIL.n412 B 0.131881f
C536 VTAIL.t7 B 0.039479f
C537 VTAIL.n413 B 0.017899f
C538 VTAIL.n414 B 0.014098f
C539 VTAIL.n415 B 0.010097f
C540 VTAIL.n416 B 1.39302f
C541 VTAIL.n417 B 0.01879f
C542 VTAIL.n418 B 0.010097f
C543 VTAIL.n419 B 0.010691f
C544 VTAIL.n420 B 0.023866f
C545 VTAIL.n421 B 0.023866f
C546 VTAIL.n422 B 0.010691f
C547 VTAIL.n423 B 0.010097f
C548 VTAIL.n424 B 0.01879f
C549 VTAIL.n425 B 0.01879f
C550 VTAIL.n426 B 0.010097f
C551 VTAIL.n427 B 0.010691f
C552 VTAIL.n428 B 0.023866f
C553 VTAIL.n429 B 0.023866f
C554 VTAIL.n430 B 0.010691f
C555 VTAIL.n431 B 0.010097f
C556 VTAIL.n432 B 0.01879f
C557 VTAIL.n433 B 0.01879f
C558 VTAIL.n434 B 0.010097f
C559 VTAIL.n435 B 0.010691f
C560 VTAIL.n436 B 0.023866f
C561 VTAIL.n437 B 0.023866f
C562 VTAIL.n438 B 0.010691f
C563 VTAIL.n439 B 0.010097f
C564 VTAIL.n440 B 0.01879f
C565 VTAIL.n441 B 0.01879f
C566 VTAIL.n442 B 0.010097f
C567 VTAIL.n443 B 0.010691f
C568 VTAIL.n444 B 0.023866f
C569 VTAIL.n445 B 0.023866f
C570 VTAIL.n446 B 0.010691f
C571 VTAIL.n447 B 0.010097f
C572 VTAIL.n448 B 0.01879f
C573 VTAIL.n449 B 0.01879f
C574 VTAIL.n450 B 0.010097f
C575 VTAIL.n451 B 0.010691f
C576 VTAIL.n452 B 0.023866f
C577 VTAIL.n453 B 0.023866f
C578 VTAIL.n454 B 0.010691f
C579 VTAIL.n455 B 0.010097f
C580 VTAIL.n456 B 0.01879f
C581 VTAIL.n457 B 0.01879f
C582 VTAIL.n458 B 0.010097f
C583 VTAIL.n459 B 0.010394f
C584 VTAIL.n460 B 0.010394f
C585 VTAIL.n461 B 0.023866f
C586 VTAIL.n462 B 0.023866f
C587 VTAIL.n463 B 0.010691f
C588 VTAIL.n464 B 0.010097f
C589 VTAIL.n465 B 0.01879f
C590 VTAIL.n466 B 0.01879f
C591 VTAIL.n467 B 0.010097f
C592 VTAIL.n468 B 0.010691f
C593 VTAIL.n469 B 0.023866f
C594 VTAIL.n470 B 0.053907f
C595 VTAIL.n471 B 0.010691f
C596 VTAIL.n472 B 0.010097f
C597 VTAIL.n473 B 0.048053f
C598 VTAIL.n474 B 0.030529f
C599 VTAIL.n475 B 0.209434f
C600 VTAIL.n476 B 0.027679f
C601 VTAIL.n477 B 0.01879f
C602 VTAIL.n478 B 0.010097f
C603 VTAIL.n479 B 0.023866f
C604 VTAIL.n480 B 0.010691f
C605 VTAIL.n481 B 0.01879f
C606 VTAIL.n482 B 0.010097f
C607 VTAIL.n483 B 0.023866f
C608 VTAIL.n484 B 0.010691f
C609 VTAIL.n485 B 0.01879f
C610 VTAIL.n486 B 0.010097f
C611 VTAIL.n487 B 0.023866f
C612 VTAIL.n488 B 0.023866f
C613 VTAIL.n489 B 0.010691f
C614 VTAIL.n490 B 0.01879f
C615 VTAIL.n491 B 0.010097f
C616 VTAIL.n492 B 0.023866f
C617 VTAIL.n493 B 0.010691f
C618 VTAIL.n494 B 0.01879f
C619 VTAIL.n495 B 0.010097f
C620 VTAIL.n496 B 0.023866f
C621 VTAIL.n497 B 0.010691f
C622 VTAIL.n498 B 0.01879f
C623 VTAIL.n499 B 0.010097f
C624 VTAIL.n500 B 0.023866f
C625 VTAIL.n501 B 0.010691f
C626 VTAIL.n502 B 0.01879f
C627 VTAIL.n503 B 0.010097f
C628 VTAIL.n504 B 0.023866f
C629 VTAIL.n505 B 0.010691f
C630 VTAIL.n506 B 0.131881f
C631 VTAIL.t14 B 0.039479f
C632 VTAIL.n507 B 0.017899f
C633 VTAIL.n508 B 0.014098f
C634 VTAIL.n509 B 0.010097f
C635 VTAIL.n510 B 1.39302f
C636 VTAIL.n511 B 0.01879f
C637 VTAIL.n512 B 0.010097f
C638 VTAIL.n513 B 0.010691f
C639 VTAIL.n514 B 0.023866f
C640 VTAIL.n515 B 0.023866f
C641 VTAIL.n516 B 0.010691f
C642 VTAIL.n517 B 0.010097f
C643 VTAIL.n518 B 0.01879f
C644 VTAIL.n519 B 0.01879f
C645 VTAIL.n520 B 0.010097f
C646 VTAIL.n521 B 0.010691f
C647 VTAIL.n522 B 0.023866f
C648 VTAIL.n523 B 0.023866f
C649 VTAIL.n524 B 0.010691f
C650 VTAIL.n525 B 0.010097f
C651 VTAIL.n526 B 0.01879f
C652 VTAIL.n527 B 0.01879f
C653 VTAIL.n528 B 0.010097f
C654 VTAIL.n529 B 0.010691f
C655 VTAIL.n530 B 0.023866f
C656 VTAIL.n531 B 0.023866f
C657 VTAIL.n532 B 0.010691f
C658 VTAIL.n533 B 0.010097f
C659 VTAIL.n534 B 0.01879f
C660 VTAIL.n535 B 0.01879f
C661 VTAIL.n536 B 0.010097f
C662 VTAIL.n537 B 0.010691f
C663 VTAIL.n538 B 0.023866f
C664 VTAIL.n539 B 0.023866f
C665 VTAIL.n540 B 0.010691f
C666 VTAIL.n541 B 0.010097f
C667 VTAIL.n542 B 0.01879f
C668 VTAIL.n543 B 0.01879f
C669 VTAIL.n544 B 0.010097f
C670 VTAIL.n545 B 0.010691f
C671 VTAIL.n546 B 0.023866f
C672 VTAIL.n547 B 0.023866f
C673 VTAIL.n548 B 0.010691f
C674 VTAIL.n549 B 0.010097f
C675 VTAIL.n550 B 0.01879f
C676 VTAIL.n551 B 0.01879f
C677 VTAIL.n552 B 0.010097f
C678 VTAIL.n553 B 0.010394f
C679 VTAIL.n554 B 0.010394f
C680 VTAIL.n555 B 0.023866f
C681 VTAIL.n556 B 0.023866f
C682 VTAIL.n557 B 0.010691f
C683 VTAIL.n558 B 0.010097f
C684 VTAIL.n559 B 0.01879f
C685 VTAIL.n560 B 0.01879f
C686 VTAIL.n561 B 0.010097f
C687 VTAIL.n562 B 0.010691f
C688 VTAIL.n563 B 0.023866f
C689 VTAIL.n564 B 0.053907f
C690 VTAIL.n565 B 0.010691f
C691 VTAIL.n566 B 0.010097f
C692 VTAIL.n567 B 0.048053f
C693 VTAIL.n568 B 0.030529f
C694 VTAIL.n569 B 0.209434f
C695 VTAIL.t11 B 0.252128f
C696 VTAIL.t8 B 0.252128f
C697 VTAIL.n570 B 2.24202f
C698 VTAIL.n571 B 0.503942f
C699 VTAIL.n572 B 0.027679f
C700 VTAIL.n573 B 0.01879f
C701 VTAIL.n574 B 0.010097f
C702 VTAIL.n575 B 0.023866f
C703 VTAIL.n576 B 0.010691f
C704 VTAIL.n577 B 0.01879f
C705 VTAIL.n578 B 0.010097f
C706 VTAIL.n579 B 0.023866f
C707 VTAIL.n580 B 0.010691f
C708 VTAIL.n581 B 0.01879f
C709 VTAIL.n582 B 0.010097f
C710 VTAIL.n583 B 0.023866f
C711 VTAIL.n584 B 0.023866f
C712 VTAIL.n585 B 0.010691f
C713 VTAIL.n586 B 0.01879f
C714 VTAIL.n587 B 0.010097f
C715 VTAIL.n588 B 0.023866f
C716 VTAIL.n589 B 0.010691f
C717 VTAIL.n590 B 0.01879f
C718 VTAIL.n591 B 0.010097f
C719 VTAIL.n592 B 0.023866f
C720 VTAIL.n593 B 0.010691f
C721 VTAIL.n594 B 0.01879f
C722 VTAIL.n595 B 0.010097f
C723 VTAIL.n596 B 0.023866f
C724 VTAIL.n597 B 0.010691f
C725 VTAIL.n598 B 0.01879f
C726 VTAIL.n599 B 0.010097f
C727 VTAIL.n600 B 0.023866f
C728 VTAIL.n601 B 0.010691f
C729 VTAIL.n602 B 0.131881f
C730 VTAIL.t15 B 0.039479f
C731 VTAIL.n603 B 0.017899f
C732 VTAIL.n604 B 0.014098f
C733 VTAIL.n605 B 0.010097f
C734 VTAIL.n606 B 1.39302f
C735 VTAIL.n607 B 0.01879f
C736 VTAIL.n608 B 0.010097f
C737 VTAIL.n609 B 0.010691f
C738 VTAIL.n610 B 0.023866f
C739 VTAIL.n611 B 0.023866f
C740 VTAIL.n612 B 0.010691f
C741 VTAIL.n613 B 0.010097f
C742 VTAIL.n614 B 0.01879f
C743 VTAIL.n615 B 0.01879f
C744 VTAIL.n616 B 0.010097f
C745 VTAIL.n617 B 0.010691f
C746 VTAIL.n618 B 0.023866f
C747 VTAIL.n619 B 0.023866f
C748 VTAIL.n620 B 0.010691f
C749 VTAIL.n621 B 0.010097f
C750 VTAIL.n622 B 0.01879f
C751 VTAIL.n623 B 0.01879f
C752 VTAIL.n624 B 0.010097f
C753 VTAIL.n625 B 0.010691f
C754 VTAIL.n626 B 0.023866f
C755 VTAIL.n627 B 0.023866f
C756 VTAIL.n628 B 0.010691f
C757 VTAIL.n629 B 0.010097f
C758 VTAIL.n630 B 0.01879f
C759 VTAIL.n631 B 0.01879f
C760 VTAIL.n632 B 0.010097f
C761 VTAIL.n633 B 0.010691f
C762 VTAIL.n634 B 0.023866f
C763 VTAIL.n635 B 0.023866f
C764 VTAIL.n636 B 0.010691f
C765 VTAIL.n637 B 0.010097f
C766 VTAIL.n638 B 0.01879f
C767 VTAIL.n639 B 0.01879f
C768 VTAIL.n640 B 0.010097f
C769 VTAIL.n641 B 0.010691f
C770 VTAIL.n642 B 0.023866f
C771 VTAIL.n643 B 0.023866f
C772 VTAIL.n644 B 0.010691f
C773 VTAIL.n645 B 0.010097f
C774 VTAIL.n646 B 0.01879f
C775 VTAIL.n647 B 0.01879f
C776 VTAIL.n648 B 0.010097f
C777 VTAIL.n649 B 0.010394f
C778 VTAIL.n650 B 0.010394f
C779 VTAIL.n651 B 0.023866f
C780 VTAIL.n652 B 0.023866f
C781 VTAIL.n653 B 0.010691f
C782 VTAIL.n654 B 0.010097f
C783 VTAIL.n655 B 0.01879f
C784 VTAIL.n656 B 0.01879f
C785 VTAIL.n657 B 0.010097f
C786 VTAIL.n658 B 0.010691f
C787 VTAIL.n659 B 0.023866f
C788 VTAIL.n660 B 0.053907f
C789 VTAIL.n661 B 0.010691f
C790 VTAIL.n662 B 0.010097f
C791 VTAIL.n663 B 0.048053f
C792 VTAIL.n664 B 0.030529f
C793 VTAIL.n665 B 1.48482f
C794 VTAIL.n666 B 0.027679f
C795 VTAIL.n667 B 0.01879f
C796 VTAIL.n668 B 0.010097f
C797 VTAIL.n669 B 0.023866f
C798 VTAIL.n670 B 0.010691f
C799 VTAIL.n671 B 0.01879f
C800 VTAIL.n672 B 0.010097f
C801 VTAIL.n673 B 0.023866f
C802 VTAIL.n674 B 0.010691f
C803 VTAIL.n675 B 0.01879f
C804 VTAIL.n676 B 0.010097f
C805 VTAIL.n677 B 0.023866f
C806 VTAIL.n678 B 0.010691f
C807 VTAIL.n679 B 0.01879f
C808 VTAIL.n680 B 0.010097f
C809 VTAIL.n681 B 0.023866f
C810 VTAIL.n682 B 0.010691f
C811 VTAIL.n683 B 0.01879f
C812 VTAIL.n684 B 0.010097f
C813 VTAIL.n685 B 0.023866f
C814 VTAIL.n686 B 0.010691f
C815 VTAIL.n687 B 0.01879f
C816 VTAIL.n688 B 0.010097f
C817 VTAIL.n689 B 0.023866f
C818 VTAIL.n690 B 0.010691f
C819 VTAIL.n691 B 0.01879f
C820 VTAIL.n692 B 0.010097f
C821 VTAIL.n693 B 0.023866f
C822 VTAIL.n694 B 0.010691f
C823 VTAIL.n695 B 0.131881f
C824 VTAIL.t2 B 0.039479f
C825 VTAIL.n696 B 0.017899f
C826 VTAIL.n697 B 0.014098f
C827 VTAIL.n698 B 0.010097f
C828 VTAIL.n699 B 1.39302f
C829 VTAIL.n700 B 0.01879f
C830 VTAIL.n701 B 0.010097f
C831 VTAIL.n702 B 0.010691f
C832 VTAIL.n703 B 0.023866f
C833 VTAIL.n704 B 0.023866f
C834 VTAIL.n705 B 0.010691f
C835 VTAIL.n706 B 0.010097f
C836 VTAIL.n707 B 0.01879f
C837 VTAIL.n708 B 0.01879f
C838 VTAIL.n709 B 0.010097f
C839 VTAIL.n710 B 0.010691f
C840 VTAIL.n711 B 0.023866f
C841 VTAIL.n712 B 0.023866f
C842 VTAIL.n713 B 0.010691f
C843 VTAIL.n714 B 0.010097f
C844 VTAIL.n715 B 0.01879f
C845 VTAIL.n716 B 0.01879f
C846 VTAIL.n717 B 0.010097f
C847 VTAIL.n718 B 0.010691f
C848 VTAIL.n719 B 0.023866f
C849 VTAIL.n720 B 0.023866f
C850 VTAIL.n721 B 0.010691f
C851 VTAIL.n722 B 0.010097f
C852 VTAIL.n723 B 0.01879f
C853 VTAIL.n724 B 0.01879f
C854 VTAIL.n725 B 0.010097f
C855 VTAIL.n726 B 0.010691f
C856 VTAIL.n727 B 0.023866f
C857 VTAIL.n728 B 0.023866f
C858 VTAIL.n729 B 0.010691f
C859 VTAIL.n730 B 0.010097f
C860 VTAIL.n731 B 0.01879f
C861 VTAIL.n732 B 0.01879f
C862 VTAIL.n733 B 0.010097f
C863 VTAIL.n734 B 0.010691f
C864 VTAIL.n735 B 0.023866f
C865 VTAIL.n736 B 0.023866f
C866 VTAIL.n737 B 0.023866f
C867 VTAIL.n738 B 0.010691f
C868 VTAIL.n739 B 0.010097f
C869 VTAIL.n740 B 0.01879f
C870 VTAIL.n741 B 0.01879f
C871 VTAIL.n742 B 0.010097f
C872 VTAIL.n743 B 0.010394f
C873 VTAIL.n744 B 0.010394f
C874 VTAIL.n745 B 0.023866f
C875 VTAIL.n746 B 0.023866f
C876 VTAIL.n747 B 0.010691f
C877 VTAIL.n748 B 0.010097f
C878 VTAIL.n749 B 0.01879f
C879 VTAIL.n750 B 0.01879f
C880 VTAIL.n751 B 0.010097f
C881 VTAIL.n752 B 0.010691f
C882 VTAIL.n753 B 0.023866f
C883 VTAIL.n754 B 0.053907f
C884 VTAIL.n755 B 0.010691f
C885 VTAIL.n756 B 0.010097f
C886 VTAIL.n757 B 0.048053f
C887 VTAIL.n758 B 0.030529f
C888 VTAIL.n759 B 1.4813f
C889 VP.n0 B 0.027217f
C890 VP.t3 B 2.67754f
C891 VP.n1 B 0.037302f
C892 VP.n2 B 0.020645f
C893 VP.t6 B 2.67754f
C894 VP.n3 B 0.929284f
C895 VP.n4 B 0.020645f
C896 VP.n5 B 0.016674f
C897 VP.n6 B 0.020645f
C898 VP.t0 B 2.67754f
C899 VP.n7 B 0.929284f
C900 VP.n8 B 0.020645f
C901 VP.n9 B 0.037302f
C902 VP.n10 B 0.027217f
C903 VP.t4 B 2.67754f
C904 VP.n11 B 0.027217f
C905 VP.t7 B 2.67754f
C906 VP.n12 B 0.037302f
C907 VP.n13 B 0.020645f
C908 VP.t1 B 2.67754f
C909 VP.n14 B 0.929284f
C910 VP.n15 B 0.020645f
C911 VP.n16 B 0.016674f
C912 VP.n17 B 0.020645f
C913 VP.t2 B 2.67754f
C914 VP.n18 B 0.984444f
C915 VP.t5 B 2.87221f
C916 VP.n19 B 0.961468f
C917 VP.n20 B 0.203368f
C918 VP.n21 B 0.021464f
C919 VP.n22 B 0.038285f
C920 VP.n23 B 0.040816f
C921 VP.n24 B 0.020645f
C922 VP.n25 B 0.020645f
C923 VP.n26 B 0.020645f
C924 VP.n27 B 0.040816f
C925 VP.n28 B 0.038285f
C926 VP.n29 B 0.021464f
C927 VP.n30 B 0.020645f
C928 VP.n31 B 0.020645f
C929 VP.n32 B 0.036206f
C930 VP.n33 B 0.04091f
C931 VP.n34 B 0.020095f
C932 VP.n35 B 0.020645f
C933 VP.n36 B 0.020645f
C934 VP.n37 B 0.020645f
C935 VP.n38 B 0.038285f
C936 VP.n39 B 0.025622f
C937 VP.n40 B 1.00089f
C938 VP.n41 B 1.33849f
C939 VP.n42 B 1.35189f
C940 VP.n43 B 1.00089f
C941 VP.n44 B 0.025622f
C942 VP.n45 B 0.038285f
C943 VP.n46 B 0.020645f
C944 VP.n47 B 0.020645f
C945 VP.n48 B 0.020645f
C946 VP.n49 B 0.020095f
C947 VP.n50 B 0.04091f
C948 VP.n51 B 0.036206f
C949 VP.n52 B 0.020645f
C950 VP.n53 B 0.020645f
C951 VP.n54 B 0.021464f
C952 VP.n55 B 0.038285f
C953 VP.n56 B 0.040816f
C954 VP.n57 B 0.020645f
C955 VP.n58 B 0.020645f
C956 VP.n59 B 0.020645f
C957 VP.n60 B 0.040816f
C958 VP.n61 B 0.038285f
C959 VP.n62 B 0.021464f
C960 VP.n63 B 0.020645f
C961 VP.n64 B 0.020645f
C962 VP.n65 B 0.036206f
C963 VP.n66 B 0.04091f
C964 VP.n67 B 0.020095f
C965 VP.n68 B 0.020645f
C966 VP.n69 B 0.020645f
C967 VP.n70 B 0.020645f
C968 VP.n71 B 0.038285f
C969 VP.n72 B 0.025622f
C970 VP.n73 B 1.00089f
C971 VP.n74 B 0.035803f
.ends

