* NGSPICE file created from diff_pair_sample_1255.ext - technology: sky130A

.subckt diff_pair_sample_1255 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=1.0725 pd=6.28 as=0.45375 ps=3.08 w=2.75 l=2.05
X1 VDD2.t5 VN.t0 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=1.0725 pd=6.28 as=0.45375 ps=3.08 w=2.75 l=2.05
X2 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=1.0725 pd=6.28 as=0 ps=0 w=2.75 l=2.05
X3 VTAIL.t6 VP.t1 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=2.05
X4 VDD2.t4 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.45375 pd=3.08 as=1.0725 ps=6.28 w=2.75 l=2.05
X5 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=1.0725 pd=6.28 as=0 ps=0 w=2.75 l=2.05
X6 VDD1.t3 VP.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.0725 pd=6.28 as=0.45375 ps=3.08 w=2.75 l=2.05
X7 VDD1.t2 VP.t3 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=0.45375 pd=3.08 as=1.0725 ps=6.28 w=2.75 l=2.05
X8 VDD2.t3 VN.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.45375 pd=3.08 as=1.0725 ps=6.28 w=2.75 l=2.05
X9 VDD2.t2 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.0725 pd=6.28 as=0.45375 ps=3.08 w=2.75 l=2.05
X10 VDD1.t1 VP.t4 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=0.45375 pd=3.08 as=1.0725 ps=6.28 w=2.75 l=2.05
X11 VTAIL.t4 VN.t4 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=2.05
X12 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.0725 pd=6.28 as=0 ps=0 w=2.75 l=2.05
X13 VTAIL.t3 VN.t5 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=2.05
X14 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.0725 pd=6.28 as=0 ps=0 w=2.75 l=2.05
X15 VTAIL.t10 VP.t5 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=2.05
R0 VP.n10 VP.n9 161.3
R1 VP.n11 VP.n6 161.3
R2 VP.n13 VP.n12 161.3
R3 VP.n14 VP.n5 161.3
R4 VP.n31 VP.n0 161.3
R5 VP.n30 VP.n29 161.3
R6 VP.n28 VP.n1 161.3
R7 VP.n27 VP.n26 161.3
R8 VP.n25 VP.n2 161.3
R9 VP.n24 VP.n23 161.3
R10 VP.n22 VP.n3 161.3
R11 VP.n21 VP.n20 161.3
R12 VP.n19 VP.n4 161.3
R13 VP.n18 VP.n17 92.1615
R14 VP.n33 VP.n32 92.1615
R15 VP.n16 VP.n15 92.1615
R16 VP.n7 VP.t0 66.2423
R17 VP.n20 VP.n3 56.5193
R18 VP.n30 VP.n1 56.5193
R19 VP.n13 VP.n6 56.5193
R20 VP.n8 VP.n7 45.9387
R21 VP.n17 VP.n16 39.5299
R22 VP.n25 VP.t5 32.3298
R23 VP.n18 VP.t2 32.3298
R24 VP.n32 VP.t4 32.3298
R25 VP.n8 VP.t1 32.3298
R26 VP.n15 VP.t3 32.3298
R27 VP.n20 VP.n19 24.4675
R28 VP.n24 VP.n3 24.4675
R29 VP.n25 VP.n24 24.4675
R30 VP.n26 VP.n25 24.4675
R31 VP.n26 VP.n1 24.4675
R32 VP.n31 VP.n30 24.4675
R33 VP.n14 VP.n13 24.4675
R34 VP.n9 VP.n8 24.4675
R35 VP.n9 VP.n6 24.4675
R36 VP.n19 VP.n18 18.5954
R37 VP.n32 VP.n31 18.5954
R38 VP.n15 VP.n14 18.5954
R39 VP.n10 VP.n7 9.10166
R40 VP.n16 VP.n5 0.278367
R41 VP.n17 VP.n4 0.278367
R42 VP.n33 VP.n0 0.278367
R43 VP.n11 VP.n10 0.189894
R44 VP.n12 VP.n11 0.189894
R45 VP.n12 VP.n5 0.189894
R46 VP.n21 VP.n4 0.189894
R47 VP.n22 VP.n21 0.189894
R48 VP.n23 VP.n22 0.189894
R49 VP.n23 VP.n2 0.189894
R50 VP.n27 VP.n2 0.189894
R51 VP.n28 VP.n27 0.189894
R52 VP.n29 VP.n28 0.189894
R53 VP.n29 VP.n0 0.189894
R54 VP VP.n33 0.153454
R55 VTAIL.n7 VTAIL.t0 71.1559
R56 VTAIL.n11 VTAIL.t2 71.1556
R57 VTAIL.n2 VTAIL.t9 71.1556
R58 VTAIL.n10 VTAIL.t8 71.1556
R59 VTAIL.n9 VTAIL.n8 63.9559
R60 VTAIL.n6 VTAIL.n5 63.9559
R61 VTAIL.n1 VTAIL.n0 63.9556
R62 VTAIL.n4 VTAIL.n3 63.9556
R63 VTAIL.n6 VTAIL.n4 18.841
R64 VTAIL.n11 VTAIL.n10 16.7893
R65 VTAIL.n0 VTAIL.t1 7.2005
R66 VTAIL.n0 VTAIL.t4 7.2005
R67 VTAIL.n3 VTAIL.t5 7.2005
R68 VTAIL.n3 VTAIL.t10 7.2005
R69 VTAIL.n8 VTAIL.t7 7.2005
R70 VTAIL.n8 VTAIL.t6 7.2005
R71 VTAIL.n5 VTAIL.t11 7.2005
R72 VTAIL.n5 VTAIL.t3 7.2005
R73 VTAIL.n7 VTAIL.n6 2.05222
R74 VTAIL.n10 VTAIL.n9 2.05222
R75 VTAIL.n4 VTAIL.n2 2.05222
R76 VTAIL.n9 VTAIL.n7 1.49619
R77 VTAIL.n2 VTAIL.n1 1.49619
R78 VTAIL VTAIL.n11 1.4811
R79 VTAIL VTAIL.n1 0.571621
R80 VDD1 VDD1.t5 89.4316
R81 VDD1.n1 VDD1.t3 89.3179
R82 VDD1.n1 VDD1.n0 81.092
R83 VDD1.n3 VDD1.n2 80.6345
R84 VDD1.n3 VDD1.n1 34.363
R85 VDD1.n2 VDD1.t4 7.2005
R86 VDD1.n2 VDD1.t2 7.2005
R87 VDD1.n0 VDD1.t0 7.2005
R88 VDD1.n0 VDD1.t1 7.2005
R89 VDD1 VDD1.n3 0.455241
R90 B.n490 B.n489 585
R91 B.n164 B.n87 585
R92 B.n163 B.n162 585
R93 B.n161 B.n160 585
R94 B.n159 B.n158 585
R95 B.n157 B.n156 585
R96 B.n155 B.n154 585
R97 B.n153 B.n152 585
R98 B.n151 B.n150 585
R99 B.n149 B.n148 585
R100 B.n147 B.n146 585
R101 B.n145 B.n144 585
R102 B.n143 B.n142 585
R103 B.n141 B.n140 585
R104 B.n139 B.n138 585
R105 B.n137 B.n136 585
R106 B.n135 B.n134 585
R107 B.n133 B.n132 585
R108 B.n131 B.n130 585
R109 B.n129 B.n128 585
R110 B.n127 B.n126 585
R111 B.n125 B.n124 585
R112 B.n123 B.n122 585
R113 B.n121 B.n120 585
R114 B.n119 B.n118 585
R115 B.n117 B.n116 585
R116 B.n115 B.n114 585
R117 B.n113 B.n112 585
R118 B.n111 B.n110 585
R119 B.n109 B.n108 585
R120 B.n107 B.n106 585
R121 B.n105 B.n104 585
R122 B.n103 B.n102 585
R123 B.n101 B.n100 585
R124 B.n99 B.n98 585
R125 B.n97 B.n96 585
R126 B.n95 B.n94 585
R127 B.n67 B.n66 585
R128 B.n488 B.n68 585
R129 B.n493 B.n68 585
R130 B.n487 B.n486 585
R131 B.n486 B.n64 585
R132 B.n485 B.n63 585
R133 B.n499 B.n63 585
R134 B.n484 B.n62 585
R135 B.n500 B.n62 585
R136 B.n483 B.n61 585
R137 B.n501 B.n61 585
R138 B.n482 B.n481 585
R139 B.n481 B.n57 585
R140 B.n480 B.n56 585
R141 B.n507 B.n56 585
R142 B.n479 B.n55 585
R143 B.n508 B.n55 585
R144 B.n478 B.n54 585
R145 B.n509 B.n54 585
R146 B.n477 B.n476 585
R147 B.n476 B.n50 585
R148 B.n475 B.n49 585
R149 B.n515 B.n49 585
R150 B.n474 B.n48 585
R151 B.n516 B.n48 585
R152 B.n473 B.n47 585
R153 B.n517 B.n47 585
R154 B.n472 B.n471 585
R155 B.n471 B.n43 585
R156 B.n470 B.n42 585
R157 B.n523 B.n42 585
R158 B.n469 B.n41 585
R159 B.n524 B.n41 585
R160 B.n468 B.n40 585
R161 B.n525 B.n40 585
R162 B.n467 B.n466 585
R163 B.n466 B.n36 585
R164 B.n465 B.n35 585
R165 B.n531 B.n35 585
R166 B.n464 B.n34 585
R167 B.n532 B.n34 585
R168 B.n463 B.n33 585
R169 B.n533 B.n33 585
R170 B.n462 B.n461 585
R171 B.n461 B.n29 585
R172 B.n460 B.n28 585
R173 B.n539 B.n28 585
R174 B.n459 B.n27 585
R175 B.n540 B.n27 585
R176 B.n458 B.n26 585
R177 B.n541 B.n26 585
R178 B.n457 B.n456 585
R179 B.n456 B.n22 585
R180 B.n455 B.n21 585
R181 B.n547 B.n21 585
R182 B.n454 B.n20 585
R183 B.n548 B.n20 585
R184 B.n453 B.n19 585
R185 B.n549 B.n19 585
R186 B.n452 B.n451 585
R187 B.n451 B.n15 585
R188 B.n450 B.n14 585
R189 B.n555 B.n14 585
R190 B.n449 B.n13 585
R191 B.n556 B.n13 585
R192 B.n448 B.n12 585
R193 B.n557 B.n12 585
R194 B.n447 B.n446 585
R195 B.n446 B.n8 585
R196 B.n445 B.n7 585
R197 B.n563 B.n7 585
R198 B.n444 B.n6 585
R199 B.n564 B.n6 585
R200 B.n443 B.n5 585
R201 B.n565 B.n5 585
R202 B.n442 B.n441 585
R203 B.n441 B.n4 585
R204 B.n440 B.n165 585
R205 B.n440 B.n439 585
R206 B.n430 B.n166 585
R207 B.n167 B.n166 585
R208 B.n432 B.n431 585
R209 B.n433 B.n432 585
R210 B.n429 B.n172 585
R211 B.n172 B.n171 585
R212 B.n428 B.n427 585
R213 B.n427 B.n426 585
R214 B.n174 B.n173 585
R215 B.n175 B.n174 585
R216 B.n419 B.n418 585
R217 B.n420 B.n419 585
R218 B.n417 B.n180 585
R219 B.n180 B.n179 585
R220 B.n416 B.n415 585
R221 B.n415 B.n414 585
R222 B.n182 B.n181 585
R223 B.n183 B.n182 585
R224 B.n407 B.n406 585
R225 B.n408 B.n407 585
R226 B.n405 B.n187 585
R227 B.n191 B.n187 585
R228 B.n404 B.n403 585
R229 B.n403 B.n402 585
R230 B.n189 B.n188 585
R231 B.n190 B.n189 585
R232 B.n395 B.n394 585
R233 B.n396 B.n395 585
R234 B.n393 B.n196 585
R235 B.n196 B.n195 585
R236 B.n392 B.n391 585
R237 B.n391 B.n390 585
R238 B.n198 B.n197 585
R239 B.n199 B.n198 585
R240 B.n383 B.n382 585
R241 B.n384 B.n383 585
R242 B.n381 B.n204 585
R243 B.n204 B.n203 585
R244 B.n380 B.n379 585
R245 B.n379 B.n378 585
R246 B.n206 B.n205 585
R247 B.n207 B.n206 585
R248 B.n371 B.n370 585
R249 B.n372 B.n371 585
R250 B.n369 B.n212 585
R251 B.n212 B.n211 585
R252 B.n368 B.n367 585
R253 B.n367 B.n366 585
R254 B.n214 B.n213 585
R255 B.n215 B.n214 585
R256 B.n359 B.n358 585
R257 B.n360 B.n359 585
R258 B.n357 B.n220 585
R259 B.n220 B.n219 585
R260 B.n356 B.n355 585
R261 B.n355 B.n354 585
R262 B.n222 B.n221 585
R263 B.n223 B.n222 585
R264 B.n347 B.n346 585
R265 B.n348 B.n347 585
R266 B.n345 B.n228 585
R267 B.n228 B.n227 585
R268 B.n344 B.n343 585
R269 B.n343 B.n342 585
R270 B.n230 B.n229 585
R271 B.n231 B.n230 585
R272 B.n335 B.n334 585
R273 B.n336 B.n335 585
R274 B.n234 B.n233 585
R275 B.n259 B.n257 585
R276 B.n260 B.n256 585
R277 B.n260 B.n235 585
R278 B.n263 B.n262 585
R279 B.n264 B.n255 585
R280 B.n266 B.n265 585
R281 B.n268 B.n254 585
R282 B.n271 B.n270 585
R283 B.n272 B.n253 585
R284 B.n274 B.n273 585
R285 B.n276 B.n252 585
R286 B.n279 B.n278 585
R287 B.n280 B.n251 585
R288 B.n285 B.n284 585
R289 B.n287 B.n250 585
R290 B.n290 B.n289 585
R291 B.n291 B.n249 585
R292 B.n293 B.n292 585
R293 B.n295 B.n248 585
R294 B.n298 B.n297 585
R295 B.n299 B.n247 585
R296 B.n301 B.n300 585
R297 B.n303 B.n246 585
R298 B.n306 B.n305 585
R299 B.n308 B.n243 585
R300 B.n310 B.n309 585
R301 B.n312 B.n242 585
R302 B.n315 B.n314 585
R303 B.n316 B.n241 585
R304 B.n318 B.n317 585
R305 B.n320 B.n240 585
R306 B.n323 B.n322 585
R307 B.n324 B.n239 585
R308 B.n326 B.n325 585
R309 B.n328 B.n238 585
R310 B.n329 B.n237 585
R311 B.n332 B.n331 585
R312 B.n333 B.n236 585
R313 B.n236 B.n235 585
R314 B.n338 B.n337 585
R315 B.n337 B.n336 585
R316 B.n339 B.n232 585
R317 B.n232 B.n231 585
R318 B.n341 B.n340 585
R319 B.n342 B.n341 585
R320 B.n226 B.n225 585
R321 B.n227 B.n226 585
R322 B.n350 B.n349 585
R323 B.n349 B.n348 585
R324 B.n351 B.n224 585
R325 B.n224 B.n223 585
R326 B.n353 B.n352 585
R327 B.n354 B.n353 585
R328 B.n218 B.n217 585
R329 B.n219 B.n218 585
R330 B.n362 B.n361 585
R331 B.n361 B.n360 585
R332 B.n363 B.n216 585
R333 B.n216 B.n215 585
R334 B.n365 B.n364 585
R335 B.n366 B.n365 585
R336 B.n210 B.n209 585
R337 B.n211 B.n210 585
R338 B.n374 B.n373 585
R339 B.n373 B.n372 585
R340 B.n375 B.n208 585
R341 B.n208 B.n207 585
R342 B.n377 B.n376 585
R343 B.n378 B.n377 585
R344 B.n202 B.n201 585
R345 B.n203 B.n202 585
R346 B.n386 B.n385 585
R347 B.n385 B.n384 585
R348 B.n387 B.n200 585
R349 B.n200 B.n199 585
R350 B.n389 B.n388 585
R351 B.n390 B.n389 585
R352 B.n194 B.n193 585
R353 B.n195 B.n194 585
R354 B.n398 B.n397 585
R355 B.n397 B.n396 585
R356 B.n399 B.n192 585
R357 B.n192 B.n190 585
R358 B.n401 B.n400 585
R359 B.n402 B.n401 585
R360 B.n186 B.n185 585
R361 B.n191 B.n186 585
R362 B.n410 B.n409 585
R363 B.n409 B.n408 585
R364 B.n411 B.n184 585
R365 B.n184 B.n183 585
R366 B.n413 B.n412 585
R367 B.n414 B.n413 585
R368 B.n178 B.n177 585
R369 B.n179 B.n178 585
R370 B.n422 B.n421 585
R371 B.n421 B.n420 585
R372 B.n423 B.n176 585
R373 B.n176 B.n175 585
R374 B.n425 B.n424 585
R375 B.n426 B.n425 585
R376 B.n170 B.n169 585
R377 B.n171 B.n170 585
R378 B.n435 B.n434 585
R379 B.n434 B.n433 585
R380 B.n436 B.n168 585
R381 B.n168 B.n167 585
R382 B.n438 B.n437 585
R383 B.n439 B.n438 585
R384 B.n2 B.n0 585
R385 B.n4 B.n2 585
R386 B.n3 B.n1 585
R387 B.n564 B.n3 585
R388 B.n562 B.n561 585
R389 B.n563 B.n562 585
R390 B.n560 B.n9 585
R391 B.n9 B.n8 585
R392 B.n559 B.n558 585
R393 B.n558 B.n557 585
R394 B.n11 B.n10 585
R395 B.n556 B.n11 585
R396 B.n554 B.n553 585
R397 B.n555 B.n554 585
R398 B.n552 B.n16 585
R399 B.n16 B.n15 585
R400 B.n551 B.n550 585
R401 B.n550 B.n549 585
R402 B.n18 B.n17 585
R403 B.n548 B.n18 585
R404 B.n546 B.n545 585
R405 B.n547 B.n546 585
R406 B.n544 B.n23 585
R407 B.n23 B.n22 585
R408 B.n543 B.n542 585
R409 B.n542 B.n541 585
R410 B.n25 B.n24 585
R411 B.n540 B.n25 585
R412 B.n538 B.n537 585
R413 B.n539 B.n538 585
R414 B.n536 B.n30 585
R415 B.n30 B.n29 585
R416 B.n535 B.n534 585
R417 B.n534 B.n533 585
R418 B.n32 B.n31 585
R419 B.n532 B.n32 585
R420 B.n530 B.n529 585
R421 B.n531 B.n530 585
R422 B.n528 B.n37 585
R423 B.n37 B.n36 585
R424 B.n527 B.n526 585
R425 B.n526 B.n525 585
R426 B.n39 B.n38 585
R427 B.n524 B.n39 585
R428 B.n522 B.n521 585
R429 B.n523 B.n522 585
R430 B.n520 B.n44 585
R431 B.n44 B.n43 585
R432 B.n519 B.n518 585
R433 B.n518 B.n517 585
R434 B.n46 B.n45 585
R435 B.n516 B.n46 585
R436 B.n514 B.n513 585
R437 B.n515 B.n514 585
R438 B.n512 B.n51 585
R439 B.n51 B.n50 585
R440 B.n511 B.n510 585
R441 B.n510 B.n509 585
R442 B.n53 B.n52 585
R443 B.n508 B.n53 585
R444 B.n506 B.n505 585
R445 B.n507 B.n506 585
R446 B.n504 B.n58 585
R447 B.n58 B.n57 585
R448 B.n503 B.n502 585
R449 B.n502 B.n501 585
R450 B.n60 B.n59 585
R451 B.n500 B.n60 585
R452 B.n498 B.n497 585
R453 B.n499 B.n498 585
R454 B.n496 B.n65 585
R455 B.n65 B.n64 585
R456 B.n495 B.n494 585
R457 B.n494 B.n493 585
R458 B.n567 B.n566 585
R459 B.n566 B.n565 585
R460 B.n337 B.n234 550.159
R461 B.n494 B.n67 550.159
R462 B.n335 B.n236 550.159
R463 B.n490 B.n68 550.159
R464 B.n492 B.n491 256.663
R465 B.n492 B.n86 256.663
R466 B.n492 B.n85 256.663
R467 B.n492 B.n84 256.663
R468 B.n492 B.n83 256.663
R469 B.n492 B.n82 256.663
R470 B.n492 B.n81 256.663
R471 B.n492 B.n80 256.663
R472 B.n492 B.n79 256.663
R473 B.n492 B.n78 256.663
R474 B.n492 B.n77 256.663
R475 B.n492 B.n76 256.663
R476 B.n492 B.n75 256.663
R477 B.n492 B.n74 256.663
R478 B.n492 B.n73 256.663
R479 B.n492 B.n72 256.663
R480 B.n492 B.n71 256.663
R481 B.n492 B.n70 256.663
R482 B.n492 B.n69 256.663
R483 B.n258 B.n235 256.663
R484 B.n261 B.n235 256.663
R485 B.n267 B.n235 256.663
R486 B.n269 B.n235 256.663
R487 B.n275 B.n235 256.663
R488 B.n277 B.n235 256.663
R489 B.n286 B.n235 256.663
R490 B.n288 B.n235 256.663
R491 B.n294 B.n235 256.663
R492 B.n296 B.n235 256.663
R493 B.n302 B.n235 256.663
R494 B.n304 B.n235 256.663
R495 B.n311 B.n235 256.663
R496 B.n313 B.n235 256.663
R497 B.n319 B.n235 256.663
R498 B.n321 B.n235 256.663
R499 B.n327 B.n235 256.663
R500 B.n330 B.n235 256.663
R501 B.n244 B.t17 239.363
R502 B.n281 B.t6 239.363
R503 B.n91 B.t10 239.363
R504 B.n88 B.t14 239.363
R505 B.n336 B.n235 179.565
R506 B.n493 B.n492 179.565
R507 B.n337 B.n232 163.367
R508 B.n341 B.n232 163.367
R509 B.n341 B.n226 163.367
R510 B.n349 B.n226 163.367
R511 B.n349 B.n224 163.367
R512 B.n353 B.n224 163.367
R513 B.n353 B.n218 163.367
R514 B.n361 B.n218 163.367
R515 B.n361 B.n216 163.367
R516 B.n365 B.n216 163.367
R517 B.n365 B.n210 163.367
R518 B.n373 B.n210 163.367
R519 B.n373 B.n208 163.367
R520 B.n377 B.n208 163.367
R521 B.n377 B.n202 163.367
R522 B.n385 B.n202 163.367
R523 B.n385 B.n200 163.367
R524 B.n389 B.n200 163.367
R525 B.n389 B.n194 163.367
R526 B.n397 B.n194 163.367
R527 B.n397 B.n192 163.367
R528 B.n401 B.n192 163.367
R529 B.n401 B.n186 163.367
R530 B.n409 B.n186 163.367
R531 B.n409 B.n184 163.367
R532 B.n413 B.n184 163.367
R533 B.n413 B.n178 163.367
R534 B.n421 B.n178 163.367
R535 B.n421 B.n176 163.367
R536 B.n425 B.n176 163.367
R537 B.n425 B.n170 163.367
R538 B.n434 B.n170 163.367
R539 B.n434 B.n168 163.367
R540 B.n438 B.n168 163.367
R541 B.n438 B.n2 163.367
R542 B.n566 B.n2 163.367
R543 B.n566 B.n3 163.367
R544 B.n562 B.n3 163.367
R545 B.n562 B.n9 163.367
R546 B.n558 B.n9 163.367
R547 B.n558 B.n11 163.367
R548 B.n554 B.n11 163.367
R549 B.n554 B.n16 163.367
R550 B.n550 B.n16 163.367
R551 B.n550 B.n18 163.367
R552 B.n546 B.n18 163.367
R553 B.n546 B.n23 163.367
R554 B.n542 B.n23 163.367
R555 B.n542 B.n25 163.367
R556 B.n538 B.n25 163.367
R557 B.n538 B.n30 163.367
R558 B.n534 B.n30 163.367
R559 B.n534 B.n32 163.367
R560 B.n530 B.n32 163.367
R561 B.n530 B.n37 163.367
R562 B.n526 B.n37 163.367
R563 B.n526 B.n39 163.367
R564 B.n522 B.n39 163.367
R565 B.n522 B.n44 163.367
R566 B.n518 B.n44 163.367
R567 B.n518 B.n46 163.367
R568 B.n514 B.n46 163.367
R569 B.n514 B.n51 163.367
R570 B.n510 B.n51 163.367
R571 B.n510 B.n53 163.367
R572 B.n506 B.n53 163.367
R573 B.n506 B.n58 163.367
R574 B.n502 B.n58 163.367
R575 B.n502 B.n60 163.367
R576 B.n498 B.n60 163.367
R577 B.n498 B.n65 163.367
R578 B.n494 B.n65 163.367
R579 B.n260 B.n259 163.367
R580 B.n262 B.n260 163.367
R581 B.n266 B.n255 163.367
R582 B.n270 B.n268 163.367
R583 B.n274 B.n253 163.367
R584 B.n278 B.n276 163.367
R585 B.n285 B.n251 163.367
R586 B.n289 B.n287 163.367
R587 B.n293 B.n249 163.367
R588 B.n297 B.n295 163.367
R589 B.n301 B.n247 163.367
R590 B.n305 B.n303 163.367
R591 B.n310 B.n243 163.367
R592 B.n314 B.n312 163.367
R593 B.n318 B.n241 163.367
R594 B.n322 B.n320 163.367
R595 B.n326 B.n239 163.367
R596 B.n329 B.n328 163.367
R597 B.n331 B.n236 163.367
R598 B.n335 B.n230 163.367
R599 B.n343 B.n230 163.367
R600 B.n343 B.n228 163.367
R601 B.n347 B.n228 163.367
R602 B.n347 B.n222 163.367
R603 B.n355 B.n222 163.367
R604 B.n355 B.n220 163.367
R605 B.n359 B.n220 163.367
R606 B.n359 B.n214 163.367
R607 B.n367 B.n214 163.367
R608 B.n367 B.n212 163.367
R609 B.n371 B.n212 163.367
R610 B.n371 B.n206 163.367
R611 B.n379 B.n206 163.367
R612 B.n379 B.n204 163.367
R613 B.n383 B.n204 163.367
R614 B.n383 B.n198 163.367
R615 B.n391 B.n198 163.367
R616 B.n391 B.n196 163.367
R617 B.n395 B.n196 163.367
R618 B.n395 B.n189 163.367
R619 B.n403 B.n189 163.367
R620 B.n403 B.n187 163.367
R621 B.n407 B.n187 163.367
R622 B.n407 B.n182 163.367
R623 B.n415 B.n182 163.367
R624 B.n415 B.n180 163.367
R625 B.n419 B.n180 163.367
R626 B.n419 B.n174 163.367
R627 B.n427 B.n174 163.367
R628 B.n427 B.n172 163.367
R629 B.n432 B.n172 163.367
R630 B.n432 B.n166 163.367
R631 B.n440 B.n166 163.367
R632 B.n441 B.n440 163.367
R633 B.n441 B.n5 163.367
R634 B.n6 B.n5 163.367
R635 B.n7 B.n6 163.367
R636 B.n446 B.n7 163.367
R637 B.n446 B.n12 163.367
R638 B.n13 B.n12 163.367
R639 B.n14 B.n13 163.367
R640 B.n451 B.n14 163.367
R641 B.n451 B.n19 163.367
R642 B.n20 B.n19 163.367
R643 B.n21 B.n20 163.367
R644 B.n456 B.n21 163.367
R645 B.n456 B.n26 163.367
R646 B.n27 B.n26 163.367
R647 B.n28 B.n27 163.367
R648 B.n461 B.n28 163.367
R649 B.n461 B.n33 163.367
R650 B.n34 B.n33 163.367
R651 B.n35 B.n34 163.367
R652 B.n466 B.n35 163.367
R653 B.n466 B.n40 163.367
R654 B.n41 B.n40 163.367
R655 B.n42 B.n41 163.367
R656 B.n471 B.n42 163.367
R657 B.n471 B.n47 163.367
R658 B.n48 B.n47 163.367
R659 B.n49 B.n48 163.367
R660 B.n476 B.n49 163.367
R661 B.n476 B.n54 163.367
R662 B.n55 B.n54 163.367
R663 B.n56 B.n55 163.367
R664 B.n481 B.n56 163.367
R665 B.n481 B.n61 163.367
R666 B.n62 B.n61 163.367
R667 B.n63 B.n62 163.367
R668 B.n486 B.n63 163.367
R669 B.n486 B.n68 163.367
R670 B.n96 B.n95 163.367
R671 B.n100 B.n99 163.367
R672 B.n104 B.n103 163.367
R673 B.n108 B.n107 163.367
R674 B.n112 B.n111 163.367
R675 B.n116 B.n115 163.367
R676 B.n120 B.n119 163.367
R677 B.n124 B.n123 163.367
R678 B.n128 B.n127 163.367
R679 B.n132 B.n131 163.367
R680 B.n136 B.n135 163.367
R681 B.n140 B.n139 163.367
R682 B.n144 B.n143 163.367
R683 B.n148 B.n147 163.367
R684 B.n152 B.n151 163.367
R685 B.n156 B.n155 163.367
R686 B.n160 B.n159 163.367
R687 B.n162 B.n87 163.367
R688 B.n244 B.t19 122.523
R689 B.n88 B.t15 122.523
R690 B.n281 B.t9 122.522
R691 B.n91 B.t12 122.522
R692 B.n336 B.n231 93.2092
R693 B.n342 B.n231 93.2092
R694 B.n342 B.n227 93.2092
R695 B.n348 B.n227 93.2092
R696 B.n348 B.n223 93.2092
R697 B.n354 B.n223 93.2092
R698 B.n360 B.n219 93.2092
R699 B.n360 B.n215 93.2092
R700 B.n366 B.n215 93.2092
R701 B.n366 B.n211 93.2092
R702 B.n372 B.n211 93.2092
R703 B.n372 B.n207 93.2092
R704 B.n378 B.n207 93.2092
R705 B.n378 B.n203 93.2092
R706 B.n384 B.n203 93.2092
R707 B.n390 B.n199 93.2092
R708 B.n390 B.n195 93.2092
R709 B.n396 B.n195 93.2092
R710 B.n396 B.n190 93.2092
R711 B.n402 B.n190 93.2092
R712 B.n402 B.n191 93.2092
R713 B.n408 B.n183 93.2092
R714 B.n414 B.n183 93.2092
R715 B.n414 B.n179 93.2092
R716 B.n420 B.n179 93.2092
R717 B.n420 B.n175 93.2092
R718 B.n426 B.n175 93.2092
R719 B.n433 B.n171 93.2092
R720 B.n433 B.n167 93.2092
R721 B.n439 B.n167 93.2092
R722 B.n439 B.n4 93.2092
R723 B.n565 B.n4 93.2092
R724 B.n565 B.n564 93.2092
R725 B.n564 B.n563 93.2092
R726 B.n563 B.n8 93.2092
R727 B.n557 B.n8 93.2092
R728 B.n557 B.n556 93.2092
R729 B.n555 B.n15 93.2092
R730 B.n549 B.n15 93.2092
R731 B.n549 B.n548 93.2092
R732 B.n548 B.n547 93.2092
R733 B.n547 B.n22 93.2092
R734 B.n541 B.n22 93.2092
R735 B.n540 B.n539 93.2092
R736 B.n539 B.n29 93.2092
R737 B.n533 B.n29 93.2092
R738 B.n533 B.n532 93.2092
R739 B.n532 B.n531 93.2092
R740 B.n531 B.n36 93.2092
R741 B.n525 B.n524 93.2092
R742 B.n524 B.n523 93.2092
R743 B.n523 B.n43 93.2092
R744 B.n517 B.n43 93.2092
R745 B.n517 B.n516 93.2092
R746 B.n516 B.n515 93.2092
R747 B.n515 B.n50 93.2092
R748 B.n509 B.n50 93.2092
R749 B.n509 B.n508 93.2092
R750 B.n507 B.n57 93.2092
R751 B.n501 B.n57 93.2092
R752 B.n501 B.n500 93.2092
R753 B.n500 B.n499 93.2092
R754 B.n499 B.n64 93.2092
R755 B.n493 B.n64 93.2092
R756 B.n384 B.t5 83.6142
R757 B.n191 B.t3 83.6142
R758 B.n426 B.t0 83.6142
R759 B.t1 B.n555 83.6142
R760 B.t4 B.n540 83.6142
R761 B.n525 B.t2 83.6142
R762 B.n245 B.t18 76.3663
R763 B.n89 B.t16 76.3663
R764 B.n282 B.t8 76.3645
R765 B.n92 B.t13 76.3645
R766 B.n258 B.n234 71.676
R767 B.n262 B.n261 71.676
R768 B.n267 B.n266 71.676
R769 B.n270 B.n269 71.676
R770 B.n275 B.n274 71.676
R771 B.n278 B.n277 71.676
R772 B.n286 B.n285 71.676
R773 B.n289 B.n288 71.676
R774 B.n294 B.n293 71.676
R775 B.n297 B.n296 71.676
R776 B.n302 B.n301 71.676
R777 B.n305 B.n304 71.676
R778 B.n311 B.n310 71.676
R779 B.n314 B.n313 71.676
R780 B.n319 B.n318 71.676
R781 B.n322 B.n321 71.676
R782 B.n327 B.n326 71.676
R783 B.n330 B.n329 71.676
R784 B.n69 B.n67 71.676
R785 B.n96 B.n70 71.676
R786 B.n100 B.n71 71.676
R787 B.n104 B.n72 71.676
R788 B.n108 B.n73 71.676
R789 B.n112 B.n74 71.676
R790 B.n116 B.n75 71.676
R791 B.n120 B.n76 71.676
R792 B.n124 B.n77 71.676
R793 B.n128 B.n78 71.676
R794 B.n132 B.n79 71.676
R795 B.n136 B.n80 71.676
R796 B.n140 B.n81 71.676
R797 B.n144 B.n82 71.676
R798 B.n148 B.n83 71.676
R799 B.n152 B.n84 71.676
R800 B.n156 B.n85 71.676
R801 B.n160 B.n86 71.676
R802 B.n491 B.n87 71.676
R803 B.n491 B.n490 71.676
R804 B.n162 B.n86 71.676
R805 B.n159 B.n85 71.676
R806 B.n155 B.n84 71.676
R807 B.n151 B.n83 71.676
R808 B.n147 B.n82 71.676
R809 B.n143 B.n81 71.676
R810 B.n139 B.n80 71.676
R811 B.n135 B.n79 71.676
R812 B.n131 B.n78 71.676
R813 B.n127 B.n77 71.676
R814 B.n123 B.n76 71.676
R815 B.n119 B.n75 71.676
R816 B.n115 B.n74 71.676
R817 B.n111 B.n73 71.676
R818 B.n107 B.n72 71.676
R819 B.n103 B.n71 71.676
R820 B.n99 B.n70 71.676
R821 B.n95 B.n69 71.676
R822 B.n259 B.n258 71.676
R823 B.n261 B.n255 71.676
R824 B.n268 B.n267 71.676
R825 B.n269 B.n253 71.676
R826 B.n276 B.n275 71.676
R827 B.n277 B.n251 71.676
R828 B.n287 B.n286 71.676
R829 B.n288 B.n249 71.676
R830 B.n295 B.n294 71.676
R831 B.n296 B.n247 71.676
R832 B.n303 B.n302 71.676
R833 B.n304 B.n243 71.676
R834 B.n312 B.n311 71.676
R835 B.n313 B.n241 71.676
R836 B.n320 B.n319 71.676
R837 B.n321 B.n239 71.676
R838 B.n328 B.n327 71.676
R839 B.n331 B.n330 71.676
R840 B.n354 B.t7 64.4242
R841 B.t11 B.n507 64.4242
R842 B.n307 B.n245 59.5399
R843 B.n283 B.n282 59.5399
R844 B.n93 B.n92 59.5399
R845 B.n90 B.n89 59.5399
R846 B.n245 B.n244 46.1581
R847 B.n282 B.n281 46.1581
R848 B.n92 B.n91 46.1581
R849 B.n89 B.n88 46.1581
R850 B.n495 B.n66 35.7468
R851 B.n334 B.n333 35.7468
R852 B.n338 B.n233 35.7468
R853 B.n489 B.n488 35.7468
R854 B.t7 B.n219 28.7855
R855 B.n508 B.t11 28.7855
R856 B B.n567 18.0485
R857 B.n94 B.n66 10.6151
R858 B.n97 B.n94 10.6151
R859 B.n98 B.n97 10.6151
R860 B.n101 B.n98 10.6151
R861 B.n102 B.n101 10.6151
R862 B.n105 B.n102 10.6151
R863 B.n106 B.n105 10.6151
R864 B.n109 B.n106 10.6151
R865 B.n110 B.n109 10.6151
R866 B.n113 B.n110 10.6151
R867 B.n114 B.n113 10.6151
R868 B.n117 B.n114 10.6151
R869 B.n118 B.n117 10.6151
R870 B.n122 B.n121 10.6151
R871 B.n125 B.n122 10.6151
R872 B.n126 B.n125 10.6151
R873 B.n129 B.n126 10.6151
R874 B.n130 B.n129 10.6151
R875 B.n133 B.n130 10.6151
R876 B.n134 B.n133 10.6151
R877 B.n137 B.n134 10.6151
R878 B.n138 B.n137 10.6151
R879 B.n142 B.n141 10.6151
R880 B.n145 B.n142 10.6151
R881 B.n146 B.n145 10.6151
R882 B.n149 B.n146 10.6151
R883 B.n150 B.n149 10.6151
R884 B.n153 B.n150 10.6151
R885 B.n154 B.n153 10.6151
R886 B.n157 B.n154 10.6151
R887 B.n158 B.n157 10.6151
R888 B.n161 B.n158 10.6151
R889 B.n163 B.n161 10.6151
R890 B.n164 B.n163 10.6151
R891 B.n489 B.n164 10.6151
R892 B.n334 B.n229 10.6151
R893 B.n344 B.n229 10.6151
R894 B.n345 B.n344 10.6151
R895 B.n346 B.n345 10.6151
R896 B.n346 B.n221 10.6151
R897 B.n356 B.n221 10.6151
R898 B.n357 B.n356 10.6151
R899 B.n358 B.n357 10.6151
R900 B.n358 B.n213 10.6151
R901 B.n368 B.n213 10.6151
R902 B.n369 B.n368 10.6151
R903 B.n370 B.n369 10.6151
R904 B.n370 B.n205 10.6151
R905 B.n380 B.n205 10.6151
R906 B.n381 B.n380 10.6151
R907 B.n382 B.n381 10.6151
R908 B.n382 B.n197 10.6151
R909 B.n392 B.n197 10.6151
R910 B.n393 B.n392 10.6151
R911 B.n394 B.n393 10.6151
R912 B.n394 B.n188 10.6151
R913 B.n404 B.n188 10.6151
R914 B.n405 B.n404 10.6151
R915 B.n406 B.n405 10.6151
R916 B.n406 B.n181 10.6151
R917 B.n416 B.n181 10.6151
R918 B.n417 B.n416 10.6151
R919 B.n418 B.n417 10.6151
R920 B.n418 B.n173 10.6151
R921 B.n428 B.n173 10.6151
R922 B.n429 B.n428 10.6151
R923 B.n431 B.n429 10.6151
R924 B.n431 B.n430 10.6151
R925 B.n430 B.n165 10.6151
R926 B.n442 B.n165 10.6151
R927 B.n443 B.n442 10.6151
R928 B.n444 B.n443 10.6151
R929 B.n445 B.n444 10.6151
R930 B.n447 B.n445 10.6151
R931 B.n448 B.n447 10.6151
R932 B.n449 B.n448 10.6151
R933 B.n450 B.n449 10.6151
R934 B.n452 B.n450 10.6151
R935 B.n453 B.n452 10.6151
R936 B.n454 B.n453 10.6151
R937 B.n455 B.n454 10.6151
R938 B.n457 B.n455 10.6151
R939 B.n458 B.n457 10.6151
R940 B.n459 B.n458 10.6151
R941 B.n460 B.n459 10.6151
R942 B.n462 B.n460 10.6151
R943 B.n463 B.n462 10.6151
R944 B.n464 B.n463 10.6151
R945 B.n465 B.n464 10.6151
R946 B.n467 B.n465 10.6151
R947 B.n468 B.n467 10.6151
R948 B.n469 B.n468 10.6151
R949 B.n470 B.n469 10.6151
R950 B.n472 B.n470 10.6151
R951 B.n473 B.n472 10.6151
R952 B.n474 B.n473 10.6151
R953 B.n475 B.n474 10.6151
R954 B.n477 B.n475 10.6151
R955 B.n478 B.n477 10.6151
R956 B.n479 B.n478 10.6151
R957 B.n480 B.n479 10.6151
R958 B.n482 B.n480 10.6151
R959 B.n483 B.n482 10.6151
R960 B.n484 B.n483 10.6151
R961 B.n485 B.n484 10.6151
R962 B.n487 B.n485 10.6151
R963 B.n488 B.n487 10.6151
R964 B.n257 B.n233 10.6151
R965 B.n257 B.n256 10.6151
R966 B.n263 B.n256 10.6151
R967 B.n264 B.n263 10.6151
R968 B.n265 B.n264 10.6151
R969 B.n265 B.n254 10.6151
R970 B.n271 B.n254 10.6151
R971 B.n272 B.n271 10.6151
R972 B.n273 B.n272 10.6151
R973 B.n273 B.n252 10.6151
R974 B.n279 B.n252 10.6151
R975 B.n280 B.n279 10.6151
R976 B.n284 B.n280 10.6151
R977 B.n290 B.n250 10.6151
R978 B.n291 B.n290 10.6151
R979 B.n292 B.n291 10.6151
R980 B.n292 B.n248 10.6151
R981 B.n298 B.n248 10.6151
R982 B.n299 B.n298 10.6151
R983 B.n300 B.n299 10.6151
R984 B.n300 B.n246 10.6151
R985 B.n306 B.n246 10.6151
R986 B.n309 B.n308 10.6151
R987 B.n309 B.n242 10.6151
R988 B.n315 B.n242 10.6151
R989 B.n316 B.n315 10.6151
R990 B.n317 B.n316 10.6151
R991 B.n317 B.n240 10.6151
R992 B.n323 B.n240 10.6151
R993 B.n324 B.n323 10.6151
R994 B.n325 B.n324 10.6151
R995 B.n325 B.n238 10.6151
R996 B.n238 B.n237 10.6151
R997 B.n332 B.n237 10.6151
R998 B.n333 B.n332 10.6151
R999 B.n339 B.n338 10.6151
R1000 B.n340 B.n339 10.6151
R1001 B.n340 B.n225 10.6151
R1002 B.n350 B.n225 10.6151
R1003 B.n351 B.n350 10.6151
R1004 B.n352 B.n351 10.6151
R1005 B.n352 B.n217 10.6151
R1006 B.n362 B.n217 10.6151
R1007 B.n363 B.n362 10.6151
R1008 B.n364 B.n363 10.6151
R1009 B.n364 B.n209 10.6151
R1010 B.n374 B.n209 10.6151
R1011 B.n375 B.n374 10.6151
R1012 B.n376 B.n375 10.6151
R1013 B.n376 B.n201 10.6151
R1014 B.n386 B.n201 10.6151
R1015 B.n387 B.n386 10.6151
R1016 B.n388 B.n387 10.6151
R1017 B.n388 B.n193 10.6151
R1018 B.n398 B.n193 10.6151
R1019 B.n399 B.n398 10.6151
R1020 B.n400 B.n399 10.6151
R1021 B.n400 B.n185 10.6151
R1022 B.n410 B.n185 10.6151
R1023 B.n411 B.n410 10.6151
R1024 B.n412 B.n411 10.6151
R1025 B.n412 B.n177 10.6151
R1026 B.n422 B.n177 10.6151
R1027 B.n423 B.n422 10.6151
R1028 B.n424 B.n423 10.6151
R1029 B.n424 B.n169 10.6151
R1030 B.n435 B.n169 10.6151
R1031 B.n436 B.n435 10.6151
R1032 B.n437 B.n436 10.6151
R1033 B.n437 B.n0 10.6151
R1034 B.n561 B.n1 10.6151
R1035 B.n561 B.n560 10.6151
R1036 B.n560 B.n559 10.6151
R1037 B.n559 B.n10 10.6151
R1038 B.n553 B.n10 10.6151
R1039 B.n553 B.n552 10.6151
R1040 B.n552 B.n551 10.6151
R1041 B.n551 B.n17 10.6151
R1042 B.n545 B.n17 10.6151
R1043 B.n545 B.n544 10.6151
R1044 B.n544 B.n543 10.6151
R1045 B.n543 B.n24 10.6151
R1046 B.n537 B.n24 10.6151
R1047 B.n537 B.n536 10.6151
R1048 B.n536 B.n535 10.6151
R1049 B.n535 B.n31 10.6151
R1050 B.n529 B.n31 10.6151
R1051 B.n529 B.n528 10.6151
R1052 B.n528 B.n527 10.6151
R1053 B.n527 B.n38 10.6151
R1054 B.n521 B.n38 10.6151
R1055 B.n521 B.n520 10.6151
R1056 B.n520 B.n519 10.6151
R1057 B.n519 B.n45 10.6151
R1058 B.n513 B.n45 10.6151
R1059 B.n513 B.n512 10.6151
R1060 B.n512 B.n511 10.6151
R1061 B.n511 B.n52 10.6151
R1062 B.n505 B.n52 10.6151
R1063 B.n505 B.n504 10.6151
R1064 B.n504 B.n503 10.6151
R1065 B.n503 B.n59 10.6151
R1066 B.n497 B.n59 10.6151
R1067 B.n497 B.n496 10.6151
R1068 B.n496 B.n495 10.6151
R1069 B.t5 B.n199 9.59552
R1070 B.n408 B.t3 9.59552
R1071 B.t0 B.n171 9.59552
R1072 B.n556 B.t1 9.59552
R1073 B.n541 B.t4 9.59552
R1074 B.t2 B.n36 9.59552
R1075 B.n118 B.n93 9.36635
R1076 B.n141 B.n90 9.36635
R1077 B.n284 B.n283 9.36635
R1078 B.n308 B.n307 9.36635
R1079 B.n567 B.n0 2.81026
R1080 B.n567 B.n1 2.81026
R1081 B.n121 B.n93 1.24928
R1082 B.n138 B.n90 1.24928
R1083 B.n283 B.n250 1.24928
R1084 B.n307 B.n306 1.24928
R1085 VN.n21 VN.n12 161.3
R1086 VN.n20 VN.n19 161.3
R1087 VN.n18 VN.n13 161.3
R1088 VN.n17 VN.n16 161.3
R1089 VN.n9 VN.n0 161.3
R1090 VN.n8 VN.n7 161.3
R1091 VN.n6 VN.n1 161.3
R1092 VN.n5 VN.n4 161.3
R1093 VN.n11 VN.n10 92.1615
R1094 VN.n23 VN.n22 92.1615
R1095 VN.n2 VN.t3 66.2423
R1096 VN.n14 VN.t2 66.2423
R1097 VN.n8 VN.n1 56.5193
R1098 VN.n20 VN.n13 56.5193
R1099 VN.n15 VN.n14 45.9387
R1100 VN.n3 VN.n2 45.9387
R1101 VN VN.n23 39.8088
R1102 VN.n3 VN.t4 32.3298
R1103 VN.n10 VN.t1 32.3298
R1104 VN.n15 VN.t5 32.3298
R1105 VN.n22 VN.t0 32.3298
R1106 VN.n4 VN.n3 24.4675
R1107 VN.n4 VN.n1 24.4675
R1108 VN.n9 VN.n8 24.4675
R1109 VN.n16 VN.n13 24.4675
R1110 VN.n16 VN.n15 24.4675
R1111 VN.n21 VN.n20 24.4675
R1112 VN.n10 VN.n9 18.5954
R1113 VN.n22 VN.n21 18.5954
R1114 VN.n17 VN.n14 9.10166
R1115 VN.n5 VN.n2 9.10166
R1116 VN.n23 VN.n12 0.278367
R1117 VN.n11 VN.n0 0.278367
R1118 VN.n19 VN.n12 0.189894
R1119 VN.n19 VN.n18 0.189894
R1120 VN.n18 VN.n17 0.189894
R1121 VN.n6 VN.n5 0.189894
R1122 VN.n7 VN.n6 0.189894
R1123 VN.n7 VN.n0 0.189894
R1124 VN VN.n11 0.153454
R1125 VDD2.n1 VDD2.t2 89.3179
R1126 VDD2.n2 VDD2.t5 87.8346
R1127 VDD2.n1 VDD2.n0 81.092
R1128 VDD2 VDD2.n3 81.0893
R1129 VDD2.n2 VDD2.n1 32.7541
R1130 VDD2.n3 VDD2.t0 7.2005
R1131 VDD2.n3 VDD2.t3 7.2005
R1132 VDD2.n0 VDD2.t1 7.2005
R1133 VDD2.n0 VDD2.t4 7.2005
R1134 VDD2 VDD2.n2 1.59748
C0 VDD2 VN 1.75338f
C1 VTAIL VP 2.36838f
C2 VTAIL VDD1 4.03157f
C3 VP VDD1 2.01267f
C4 VTAIL VDD2 4.08069f
C5 VDD2 VP 0.417065f
C6 VDD2 VDD1 1.20077f
C7 VTAIL VN 2.35422f
C8 VP VN 4.68768f
C9 VDD1 VN 0.155475f
C10 VDD2 B 3.74458f
C11 VDD1 B 4.171769f
C12 VTAIL B 3.492687f
C13 VN B 10.2019f
C14 VP B 9.039652f
C15 VDD2.t2 B 0.321836f
C16 VDD2.t1 B 0.034238f
C17 VDD2.t4 B 0.034238f
C18 VDD2.n0 B 0.251517f
C19 VDD2.n1 B 1.29423f
C20 VDD2.t5 B 0.318133f
C21 VDD2.n2 B 1.17371f
C22 VDD2.t0 B 0.034238f
C23 VDD2.t3 B 0.034238f
C24 VDD2.n3 B 0.251502f
C25 VN.n0 B 0.035605f
C26 VN.t1 B 0.374951f
C27 VN.n1 B 0.034909f
C28 VN.t3 B 0.533115f
C29 VN.n2 B 0.220216f
C30 VN.t4 B 0.374951f
C31 VN.n3 B 0.247036f
C32 VN.n4 B 0.050333f
C33 VN.n5 B 0.226158f
C34 VN.n6 B 0.027006f
C35 VN.n7 B 0.027006f
C36 VN.n8 B 0.04394f
C37 VN.n9 B 0.044369f
C38 VN.n10 B 0.24996f
C39 VN.n11 B 0.03394f
C40 VN.n12 B 0.035605f
C41 VN.t0 B 0.374951f
C42 VN.n13 B 0.034909f
C43 VN.t2 B 0.533115f
C44 VN.n14 B 0.220216f
C45 VN.t5 B 0.374951f
C46 VN.n15 B 0.247036f
C47 VN.n16 B 0.050333f
C48 VN.n17 B 0.226158f
C49 VN.n18 B 0.027006f
C50 VN.n19 B 0.027006f
C51 VN.n20 B 0.04394f
C52 VN.n21 B 0.044369f
C53 VN.n22 B 0.24996f
C54 VN.n23 B 1.04431f
C55 VDD1.t5 B 0.464933f
C56 VDD1.t3 B 0.464388f
C57 VDD1.t0 B 0.049403f
C58 VDD1.t1 B 0.049403f
C59 VDD1.n0 B 0.362922f
C60 VDD1.n1 B 1.95976f
C61 VDD1.t4 B 0.049403f
C62 VDD1.t2 B 0.049403f
C63 VDD1.n2 B 0.360884f
C64 VDD1.n3 B 1.71533f
C65 VTAIL.t1 B 0.067924f
C66 VTAIL.t4 B 0.067924f
C67 VTAIL.n0 B 0.437827f
C68 VTAIL.n1 B 0.453681f
C69 VTAIL.t9 B 0.566899f
C70 VTAIL.n2 B 0.658972f
C71 VTAIL.t5 B 0.067924f
C72 VTAIL.t10 B 0.067924f
C73 VTAIL.n3 B 0.437827f
C74 VTAIL.n4 B 1.52877f
C75 VTAIL.t11 B 0.067924f
C76 VTAIL.t3 B 0.067924f
C77 VTAIL.n5 B 0.437829f
C78 VTAIL.n6 B 1.52877f
C79 VTAIL.t0 B 0.566901f
C80 VTAIL.n7 B 0.65897f
C81 VTAIL.t7 B 0.067924f
C82 VTAIL.t6 B 0.067924f
C83 VTAIL.n8 B 0.437829f
C84 VTAIL.n9 B 0.602796f
C85 VTAIL.t8 B 0.566899f
C86 VTAIL.n10 B 1.37831f
C87 VTAIL.t2 B 0.566899f
C88 VTAIL.n11 B 1.32079f
C89 VP.n0 B 0.04588f
C90 VP.t4 B 0.483154f
C91 VP.n1 B 0.044983f
C92 VP.n2 B 0.0348f
C93 VP.t5 B 0.483154f
C94 VP.n3 B 0.044983f
C95 VP.n4 B 0.04588f
C96 VP.t2 B 0.483154f
C97 VP.n5 B 0.04588f
C98 VP.t3 B 0.483154f
C99 VP.n6 B 0.044983f
C100 VP.t0 B 0.686961f
C101 VP.n7 B 0.283766f
C102 VP.t1 B 0.483154f
C103 VP.n8 B 0.318326f
C104 VP.n9 B 0.064858f
C105 VP.n10 B 0.291423f
C106 VP.n11 B 0.0348f
C107 VP.n12 B 0.0348f
C108 VP.n13 B 0.056619f
C109 VP.n14 B 0.057173f
C110 VP.n15 B 0.322093f
C111 VP.n16 B 1.32619f
C112 VP.n17 B 1.35783f
C113 VP.n18 B 0.322093f
C114 VP.n19 B 0.057173f
C115 VP.n20 B 0.056619f
C116 VP.n21 B 0.0348f
C117 VP.n22 B 0.0348f
C118 VP.n23 B 0.0348f
C119 VP.n24 B 0.064858f
C120 VP.n25 B 0.248123f
C121 VP.n26 B 0.064858f
C122 VP.n27 B 0.0348f
C123 VP.n28 B 0.0348f
C124 VP.n29 B 0.0348f
C125 VP.n30 B 0.056619f
C126 VP.n31 B 0.057173f
C127 VP.n32 B 0.322093f
C128 VP.n33 B 0.043734f
.ends

