* NGSPICE file created from diff_pair_sample_0637.ext - technology: sky130A

.subckt diff_pair_sample_0637 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=7.5426 pd=39.46 as=7.5426 ps=39.46 w=19.34 l=3.7
X1 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=7.5426 pd=39.46 as=7.5426 ps=39.46 w=19.34 l=3.7
X2 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.5426 pd=39.46 as=7.5426 ps=39.46 w=19.34 l=3.7
X3 VDD2.t0 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=7.5426 pd=39.46 as=7.5426 ps=39.46 w=19.34 l=3.7
X4 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=7.5426 pd=39.46 as=0 ps=0 w=19.34 l=3.7
X5 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=7.5426 pd=39.46 as=0 ps=0 w=19.34 l=3.7
X6 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.5426 pd=39.46 as=0 ps=0 w=19.34 l=3.7
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=7.5426 pd=39.46 as=0 ps=0 w=19.34 l=3.7
R0 VN VN.t1 214.01
R1 VN VN.t0 161.685
R2 VTAIL.n1 VTAIL.t3 45.344
R3 VTAIL.n3 VTAIL.t2 45.3438
R4 VTAIL.n0 VTAIL.t1 45.3438
R5 VTAIL.n2 VTAIL.t0 45.3438
R6 VTAIL.n1 VTAIL.n0 35.9876
R7 VTAIL.n3 VTAIL.n2 32.5134
R8 VTAIL.n2 VTAIL.n1 2.2074
R9 VTAIL VTAIL.n0 1.39705
R10 VTAIL VTAIL.n3 0.810845
R11 VDD2.n0 VDD2.t1 109.302
R12 VDD2.n0 VDD2.t0 62.0226
R13 VDD2 VDD2.n0 0.927224
R14 B.n948 B.n947 585
R15 B.n402 B.n129 585
R16 B.n401 B.n400 585
R17 B.n399 B.n398 585
R18 B.n397 B.n396 585
R19 B.n395 B.n394 585
R20 B.n393 B.n392 585
R21 B.n391 B.n390 585
R22 B.n389 B.n388 585
R23 B.n387 B.n386 585
R24 B.n385 B.n384 585
R25 B.n383 B.n382 585
R26 B.n381 B.n380 585
R27 B.n379 B.n378 585
R28 B.n377 B.n376 585
R29 B.n375 B.n374 585
R30 B.n373 B.n372 585
R31 B.n371 B.n370 585
R32 B.n369 B.n368 585
R33 B.n367 B.n366 585
R34 B.n365 B.n364 585
R35 B.n363 B.n362 585
R36 B.n361 B.n360 585
R37 B.n359 B.n358 585
R38 B.n357 B.n356 585
R39 B.n355 B.n354 585
R40 B.n353 B.n352 585
R41 B.n351 B.n350 585
R42 B.n349 B.n348 585
R43 B.n347 B.n346 585
R44 B.n345 B.n344 585
R45 B.n343 B.n342 585
R46 B.n341 B.n340 585
R47 B.n339 B.n338 585
R48 B.n337 B.n336 585
R49 B.n335 B.n334 585
R50 B.n333 B.n332 585
R51 B.n331 B.n330 585
R52 B.n329 B.n328 585
R53 B.n327 B.n326 585
R54 B.n325 B.n324 585
R55 B.n323 B.n322 585
R56 B.n321 B.n320 585
R57 B.n319 B.n318 585
R58 B.n317 B.n316 585
R59 B.n315 B.n314 585
R60 B.n313 B.n312 585
R61 B.n311 B.n310 585
R62 B.n309 B.n308 585
R63 B.n307 B.n306 585
R64 B.n305 B.n304 585
R65 B.n303 B.n302 585
R66 B.n301 B.n300 585
R67 B.n299 B.n298 585
R68 B.n297 B.n296 585
R69 B.n295 B.n294 585
R70 B.n293 B.n292 585
R71 B.n291 B.n290 585
R72 B.n289 B.n288 585
R73 B.n287 B.n286 585
R74 B.n285 B.n284 585
R75 B.n283 B.n282 585
R76 B.n281 B.n280 585
R77 B.n278 B.n277 585
R78 B.n276 B.n275 585
R79 B.n274 B.n273 585
R80 B.n272 B.n271 585
R81 B.n270 B.n269 585
R82 B.n268 B.n267 585
R83 B.n266 B.n265 585
R84 B.n264 B.n263 585
R85 B.n262 B.n261 585
R86 B.n260 B.n259 585
R87 B.n257 B.n256 585
R88 B.n255 B.n254 585
R89 B.n253 B.n252 585
R90 B.n251 B.n250 585
R91 B.n249 B.n248 585
R92 B.n247 B.n246 585
R93 B.n245 B.n244 585
R94 B.n243 B.n242 585
R95 B.n241 B.n240 585
R96 B.n239 B.n238 585
R97 B.n237 B.n236 585
R98 B.n235 B.n234 585
R99 B.n233 B.n232 585
R100 B.n231 B.n230 585
R101 B.n229 B.n228 585
R102 B.n227 B.n226 585
R103 B.n225 B.n224 585
R104 B.n223 B.n222 585
R105 B.n221 B.n220 585
R106 B.n219 B.n218 585
R107 B.n217 B.n216 585
R108 B.n215 B.n214 585
R109 B.n213 B.n212 585
R110 B.n211 B.n210 585
R111 B.n209 B.n208 585
R112 B.n207 B.n206 585
R113 B.n205 B.n204 585
R114 B.n203 B.n202 585
R115 B.n201 B.n200 585
R116 B.n199 B.n198 585
R117 B.n197 B.n196 585
R118 B.n195 B.n194 585
R119 B.n193 B.n192 585
R120 B.n191 B.n190 585
R121 B.n189 B.n188 585
R122 B.n187 B.n186 585
R123 B.n185 B.n184 585
R124 B.n183 B.n182 585
R125 B.n181 B.n180 585
R126 B.n179 B.n178 585
R127 B.n177 B.n176 585
R128 B.n175 B.n174 585
R129 B.n173 B.n172 585
R130 B.n171 B.n170 585
R131 B.n169 B.n168 585
R132 B.n167 B.n166 585
R133 B.n165 B.n164 585
R134 B.n163 B.n162 585
R135 B.n161 B.n160 585
R136 B.n159 B.n158 585
R137 B.n157 B.n156 585
R138 B.n155 B.n154 585
R139 B.n153 B.n152 585
R140 B.n151 B.n150 585
R141 B.n149 B.n148 585
R142 B.n147 B.n146 585
R143 B.n145 B.n144 585
R144 B.n143 B.n142 585
R145 B.n141 B.n140 585
R146 B.n139 B.n138 585
R147 B.n137 B.n136 585
R148 B.n135 B.n134 585
R149 B.n60 B.n59 585
R150 B.n946 B.n61 585
R151 B.n951 B.n61 585
R152 B.n945 B.n944 585
R153 B.n944 B.n57 585
R154 B.n943 B.n56 585
R155 B.n957 B.n56 585
R156 B.n942 B.n55 585
R157 B.n958 B.n55 585
R158 B.n941 B.n54 585
R159 B.n959 B.n54 585
R160 B.n940 B.n939 585
R161 B.n939 B.n50 585
R162 B.n938 B.n49 585
R163 B.n965 B.n49 585
R164 B.n937 B.n48 585
R165 B.n966 B.n48 585
R166 B.n936 B.n47 585
R167 B.n967 B.n47 585
R168 B.n935 B.n934 585
R169 B.n934 B.n46 585
R170 B.n933 B.n42 585
R171 B.n973 B.n42 585
R172 B.n932 B.n41 585
R173 B.n974 B.n41 585
R174 B.n931 B.n40 585
R175 B.n975 B.n40 585
R176 B.n930 B.n929 585
R177 B.n929 B.n36 585
R178 B.n928 B.n35 585
R179 B.n981 B.n35 585
R180 B.n927 B.n34 585
R181 B.n982 B.n34 585
R182 B.n926 B.n33 585
R183 B.n983 B.n33 585
R184 B.n925 B.n924 585
R185 B.n924 B.n29 585
R186 B.n923 B.n28 585
R187 B.n989 B.n28 585
R188 B.n922 B.n27 585
R189 B.n990 B.n27 585
R190 B.n921 B.n26 585
R191 B.n991 B.n26 585
R192 B.n920 B.n919 585
R193 B.n919 B.n22 585
R194 B.n918 B.n21 585
R195 B.n997 B.n21 585
R196 B.n917 B.n20 585
R197 B.n998 B.n20 585
R198 B.n916 B.n19 585
R199 B.n999 B.n19 585
R200 B.n915 B.n914 585
R201 B.n914 B.n15 585
R202 B.n913 B.n14 585
R203 B.n1005 B.n14 585
R204 B.n912 B.n13 585
R205 B.n1006 B.n13 585
R206 B.n911 B.n12 585
R207 B.n1007 B.n12 585
R208 B.n910 B.n909 585
R209 B.n909 B.n8 585
R210 B.n908 B.n7 585
R211 B.n1013 B.n7 585
R212 B.n907 B.n6 585
R213 B.n1014 B.n6 585
R214 B.n906 B.n5 585
R215 B.n1015 B.n5 585
R216 B.n905 B.n904 585
R217 B.n904 B.n4 585
R218 B.n903 B.n403 585
R219 B.n903 B.n902 585
R220 B.n893 B.n404 585
R221 B.n405 B.n404 585
R222 B.n895 B.n894 585
R223 B.n896 B.n895 585
R224 B.n892 B.n410 585
R225 B.n410 B.n409 585
R226 B.n891 B.n890 585
R227 B.n890 B.n889 585
R228 B.n412 B.n411 585
R229 B.n413 B.n412 585
R230 B.n882 B.n881 585
R231 B.n883 B.n882 585
R232 B.n880 B.n418 585
R233 B.n418 B.n417 585
R234 B.n879 B.n878 585
R235 B.n878 B.n877 585
R236 B.n420 B.n419 585
R237 B.n421 B.n420 585
R238 B.n870 B.n869 585
R239 B.n871 B.n870 585
R240 B.n868 B.n426 585
R241 B.n426 B.n425 585
R242 B.n867 B.n866 585
R243 B.n866 B.n865 585
R244 B.n428 B.n427 585
R245 B.n429 B.n428 585
R246 B.n858 B.n857 585
R247 B.n859 B.n858 585
R248 B.n856 B.n434 585
R249 B.n434 B.n433 585
R250 B.n855 B.n854 585
R251 B.n854 B.n853 585
R252 B.n436 B.n435 585
R253 B.n437 B.n436 585
R254 B.n846 B.n845 585
R255 B.n847 B.n846 585
R256 B.n844 B.n442 585
R257 B.n442 B.n441 585
R258 B.n843 B.n842 585
R259 B.n842 B.n841 585
R260 B.n444 B.n443 585
R261 B.n834 B.n444 585
R262 B.n833 B.n832 585
R263 B.n835 B.n833 585
R264 B.n831 B.n449 585
R265 B.n449 B.n448 585
R266 B.n830 B.n829 585
R267 B.n829 B.n828 585
R268 B.n451 B.n450 585
R269 B.n452 B.n451 585
R270 B.n821 B.n820 585
R271 B.n822 B.n821 585
R272 B.n819 B.n457 585
R273 B.n457 B.n456 585
R274 B.n818 B.n817 585
R275 B.n817 B.n816 585
R276 B.n459 B.n458 585
R277 B.n460 B.n459 585
R278 B.n809 B.n808 585
R279 B.n810 B.n809 585
R280 B.n463 B.n462 585
R281 B.n540 B.n539 585
R282 B.n541 B.n537 585
R283 B.n537 B.n464 585
R284 B.n543 B.n542 585
R285 B.n545 B.n536 585
R286 B.n548 B.n547 585
R287 B.n549 B.n535 585
R288 B.n551 B.n550 585
R289 B.n553 B.n534 585
R290 B.n556 B.n555 585
R291 B.n557 B.n533 585
R292 B.n559 B.n558 585
R293 B.n561 B.n532 585
R294 B.n564 B.n563 585
R295 B.n565 B.n531 585
R296 B.n567 B.n566 585
R297 B.n569 B.n530 585
R298 B.n572 B.n571 585
R299 B.n573 B.n529 585
R300 B.n575 B.n574 585
R301 B.n577 B.n528 585
R302 B.n580 B.n579 585
R303 B.n581 B.n527 585
R304 B.n583 B.n582 585
R305 B.n585 B.n526 585
R306 B.n588 B.n587 585
R307 B.n589 B.n525 585
R308 B.n591 B.n590 585
R309 B.n593 B.n524 585
R310 B.n596 B.n595 585
R311 B.n597 B.n523 585
R312 B.n599 B.n598 585
R313 B.n601 B.n522 585
R314 B.n604 B.n603 585
R315 B.n605 B.n521 585
R316 B.n607 B.n606 585
R317 B.n609 B.n520 585
R318 B.n612 B.n611 585
R319 B.n613 B.n519 585
R320 B.n615 B.n614 585
R321 B.n617 B.n518 585
R322 B.n620 B.n619 585
R323 B.n621 B.n517 585
R324 B.n623 B.n622 585
R325 B.n625 B.n516 585
R326 B.n628 B.n627 585
R327 B.n629 B.n515 585
R328 B.n631 B.n630 585
R329 B.n633 B.n514 585
R330 B.n636 B.n635 585
R331 B.n637 B.n513 585
R332 B.n639 B.n638 585
R333 B.n641 B.n512 585
R334 B.n644 B.n643 585
R335 B.n645 B.n511 585
R336 B.n647 B.n646 585
R337 B.n649 B.n510 585
R338 B.n652 B.n651 585
R339 B.n653 B.n509 585
R340 B.n655 B.n654 585
R341 B.n657 B.n508 585
R342 B.n660 B.n659 585
R343 B.n661 B.n505 585
R344 B.n664 B.n663 585
R345 B.n666 B.n504 585
R346 B.n669 B.n668 585
R347 B.n670 B.n503 585
R348 B.n672 B.n671 585
R349 B.n674 B.n502 585
R350 B.n677 B.n676 585
R351 B.n678 B.n501 585
R352 B.n680 B.n679 585
R353 B.n682 B.n500 585
R354 B.n685 B.n684 585
R355 B.n686 B.n496 585
R356 B.n688 B.n687 585
R357 B.n690 B.n495 585
R358 B.n693 B.n692 585
R359 B.n694 B.n494 585
R360 B.n696 B.n695 585
R361 B.n698 B.n493 585
R362 B.n701 B.n700 585
R363 B.n702 B.n492 585
R364 B.n704 B.n703 585
R365 B.n706 B.n491 585
R366 B.n709 B.n708 585
R367 B.n710 B.n490 585
R368 B.n712 B.n711 585
R369 B.n714 B.n489 585
R370 B.n717 B.n716 585
R371 B.n718 B.n488 585
R372 B.n720 B.n719 585
R373 B.n722 B.n487 585
R374 B.n725 B.n724 585
R375 B.n726 B.n486 585
R376 B.n728 B.n727 585
R377 B.n730 B.n485 585
R378 B.n733 B.n732 585
R379 B.n734 B.n484 585
R380 B.n736 B.n735 585
R381 B.n738 B.n483 585
R382 B.n741 B.n740 585
R383 B.n742 B.n482 585
R384 B.n744 B.n743 585
R385 B.n746 B.n481 585
R386 B.n749 B.n748 585
R387 B.n750 B.n480 585
R388 B.n752 B.n751 585
R389 B.n754 B.n479 585
R390 B.n757 B.n756 585
R391 B.n758 B.n478 585
R392 B.n760 B.n759 585
R393 B.n762 B.n477 585
R394 B.n765 B.n764 585
R395 B.n766 B.n476 585
R396 B.n768 B.n767 585
R397 B.n770 B.n475 585
R398 B.n773 B.n772 585
R399 B.n774 B.n474 585
R400 B.n776 B.n775 585
R401 B.n778 B.n473 585
R402 B.n781 B.n780 585
R403 B.n782 B.n472 585
R404 B.n784 B.n783 585
R405 B.n786 B.n471 585
R406 B.n789 B.n788 585
R407 B.n790 B.n470 585
R408 B.n792 B.n791 585
R409 B.n794 B.n469 585
R410 B.n797 B.n796 585
R411 B.n798 B.n468 585
R412 B.n800 B.n799 585
R413 B.n802 B.n467 585
R414 B.n803 B.n466 585
R415 B.n806 B.n805 585
R416 B.n807 B.n465 585
R417 B.n465 B.n464 585
R418 B.n812 B.n811 585
R419 B.n811 B.n810 585
R420 B.n813 B.n461 585
R421 B.n461 B.n460 585
R422 B.n815 B.n814 585
R423 B.n816 B.n815 585
R424 B.n455 B.n454 585
R425 B.n456 B.n455 585
R426 B.n824 B.n823 585
R427 B.n823 B.n822 585
R428 B.n825 B.n453 585
R429 B.n453 B.n452 585
R430 B.n827 B.n826 585
R431 B.n828 B.n827 585
R432 B.n447 B.n446 585
R433 B.n448 B.n447 585
R434 B.n837 B.n836 585
R435 B.n836 B.n835 585
R436 B.n838 B.n445 585
R437 B.n834 B.n445 585
R438 B.n840 B.n839 585
R439 B.n841 B.n840 585
R440 B.n440 B.n439 585
R441 B.n441 B.n440 585
R442 B.n849 B.n848 585
R443 B.n848 B.n847 585
R444 B.n850 B.n438 585
R445 B.n438 B.n437 585
R446 B.n852 B.n851 585
R447 B.n853 B.n852 585
R448 B.n432 B.n431 585
R449 B.n433 B.n432 585
R450 B.n861 B.n860 585
R451 B.n860 B.n859 585
R452 B.n862 B.n430 585
R453 B.n430 B.n429 585
R454 B.n864 B.n863 585
R455 B.n865 B.n864 585
R456 B.n424 B.n423 585
R457 B.n425 B.n424 585
R458 B.n873 B.n872 585
R459 B.n872 B.n871 585
R460 B.n874 B.n422 585
R461 B.n422 B.n421 585
R462 B.n876 B.n875 585
R463 B.n877 B.n876 585
R464 B.n416 B.n415 585
R465 B.n417 B.n416 585
R466 B.n885 B.n884 585
R467 B.n884 B.n883 585
R468 B.n886 B.n414 585
R469 B.n414 B.n413 585
R470 B.n888 B.n887 585
R471 B.n889 B.n888 585
R472 B.n408 B.n407 585
R473 B.n409 B.n408 585
R474 B.n898 B.n897 585
R475 B.n897 B.n896 585
R476 B.n899 B.n406 585
R477 B.n406 B.n405 585
R478 B.n901 B.n900 585
R479 B.n902 B.n901 585
R480 B.n2 B.n0 585
R481 B.n4 B.n2 585
R482 B.n3 B.n1 585
R483 B.n1014 B.n3 585
R484 B.n1012 B.n1011 585
R485 B.n1013 B.n1012 585
R486 B.n1010 B.n9 585
R487 B.n9 B.n8 585
R488 B.n1009 B.n1008 585
R489 B.n1008 B.n1007 585
R490 B.n11 B.n10 585
R491 B.n1006 B.n11 585
R492 B.n1004 B.n1003 585
R493 B.n1005 B.n1004 585
R494 B.n1002 B.n16 585
R495 B.n16 B.n15 585
R496 B.n1001 B.n1000 585
R497 B.n1000 B.n999 585
R498 B.n18 B.n17 585
R499 B.n998 B.n18 585
R500 B.n996 B.n995 585
R501 B.n997 B.n996 585
R502 B.n994 B.n23 585
R503 B.n23 B.n22 585
R504 B.n993 B.n992 585
R505 B.n992 B.n991 585
R506 B.n25 B.n24 585
R507 B.n990 B.n25 585
R508 B.n988 B.n987 585
R509 B.n989 B.n988 585
R510 B.n986 B.n30 585
R511 B.n30 B.n29 585
R512 B.n985 B.n984 585
R513 B.n984 B.n983 585
R514 B.n32 B.n31 585
R515 B.n982 B.n32 585
R516 B.n980 B.n979 585
R517 B.n981 B.n980 585
R518 B.n978 B.n37 585
R519 B.n37 B.n36 585
R520 B.n977 B.n976 585
R521 B.n976 B.n975 585
R522 B.n39 B.n38 585
R523 B.n974 B.n39 585
R524 B.n972 B.n971 585
R525 B.n973 B.n972 585
R526 B.n970 B.n43 585
R527 B.n46 B.n43 585
R528 B.n969 B.n968 585
R529 B.n968 B.n967 585
R530 B.n45 B.n44 585
R531 B.n966 B.n45 585
R532 B.n964 B.n963 585
R533 B.n965 B.n964 585
R534 B.n962 B.n51 585
R535 B.n51 B.n50 585
R536 B.n961 B.n960 585
R537 B.n960 B.n959 585
R538 B.n53 B.n52 585
R539 B.n958 B.n53 585
R540 B.n956 B.n955 585
R541 B.n957 B.n956 585
R542 B.n954 B.n58 585
R543 B.n58 B.n57 585
R544 B.n953 B.n952 585
R545 B.n952 B.n951 585
R546 B.n1017 B.n1016 585
R547 B.n1016 B.n1015 585
R548 B.n811 B.n463 468.476
R549 B.n952 B.n60 468.476
R550 B.n809 B.n465 468.476
R551 B.n948 B.n61 468.476
R552 B.n497 B.t10 335.236
R553 B.n506 B.t6 335.236
R554 B.n132 B.t13 335.236
R555 B.n130 B.t2 335.236
R556 B.n950 B.n949 256.663
R557 B.n950 B.n128 256.663
R558 B.n950 B.n127 256.663
R559 B.n950 B.n126 256.663
R560 B.n950 B.n125 256.663
R561 B.n950 B.n124 256.663
R562 B.n950 B.n123 256.663
R563 B.n950 B.n122 256.663
R564 B.n950 B.n121 256.663
R565 B.n950 B.n120 256.663
R566 B.n950 B.n119 256.663
R567 B.n950 B.n118 256.663
R568 B.n950 B.n117 256.663
R569 B.n950 B.n116 256.663
R570 B.n950 B.n115 256.663
R571 B.n950 B.n114 256.663
R572 B.n950 B.n113 256.663
R573 B.n950 B.n112 256.663
R574 B.n950 B.n111 256.663
R575 B.n950 B.n110 256.663
R576 B.n950 B.n109 256.663
R577 B.n950 B.n108 256.663
R578 B.n950 B.n107 256.663
R579 B.n950 B.n106 256.663
R580 B.n950 B.n105 256.663
R581 B.n950 B.n104 256.663
R582 B.n950 B.n103 256.663
R583 B.n950 B.n102 256.663
R584 B.n950 B.n101 256.663
R585 B.n950 B.n100 256.663
R586 B.n950 B.n99 256.663
R587 B.n950 B.n98 256.663
R588 B.n950 B.n97 256.663
R589 B.n950 B.n96 256.663
R590 B.n950 B.n95 256.663
R591 B.n950 B.n94 256.663
R592 B.n950 B.n93 256.663
R593 B.n950 B.n92 256.663
R594 B.n950 B.n91 256.663
R595 B.n950 B.n90 256.663
R596 B.n950 B.n89 256.663
R597 B.n950 B.n88 256.663
R598 B.n950 B.n87 256.663
R599 B.n950 B.n86 256.663
R600 B.n950 B.n85 256.663
R601 B.n950 B.n84 256.663
R602 B.n950 B.n83 256.663
R603 B.n950 B.n82 256.663
R604 B.n950 B.n81 256.663
R605 B.n950 B.n80 256.663
R606 B.n950 B.n79 256.663
R607 B.n950 B.n78 256.663
R608 B.n950 B.n77 256.663
R609 B.n950 B.n76 256.663
R610 B.n950 B.n75 256.663
R611 B.n950 B.n74 256.663
R612 B.n950 B.n73 256.663
R613 B.n950 B.n72 256.663
R614 B.n950 B.n71 256.663
R615 B.n950 B.n70 256.663
R616 B.n950 B.n69 256.663
R617 B.n950 B.n68 256.663
R618 B.n950 B.n67 256.663
R619 B.n950 B.n66 256.663
R620 B.n950 B.n65 256.663
R621 B.n950 B.n64 256.663
R622 B.n950 B.n63 256.663
R623 B.n950 B.n62 256.663
R624 B.n538 B.n464 256.663
R625 B.n544 B.n464 256.663
R626 B.n546 B.n464 256.663
R627 B.n552 B.n464 256.663
R628 B.n554 B.n464 256.663
R629 B.n560 B.n464 256.663
R630 B.n562 B.n464 256.663
R631 B.n568 B.n464 256.663
R632 B.n570 B.n464 256.663
R633 B.n576 B.n464 256.663
R634 B.n578 B.n464 256.663
R635 B.n584 B.n464 256.663
R636 B.n586 B.n464 256.663
R637 B.n592 B.n464 256.663
R638 B.n594 B.n464 256.663
R639 B.n600 B.n464 256.663
R640 B.n602 B.n464 256.663
R641 B.n608 B.n464 256.663
R642 B.n610 B.n464 256.663
R643 B.n616 B.n464 256.663
R644 B.n618 B.n464 256.663
R645 B.n624 B.n464 256.663
R646 B.n626 B.n464 256.663
R647 B.n632 B.n464 256.663
R648 B.n634 B.n464 256.663
R649 B.n640 B.n464 256.663
R650 B.n642 B.n464 256.663
R651 B.n648 B.n464 256.663
R652 B.n650 B.n464 256.663
R653 B.n656 B.n464 256.663
R654 B.n658 B.n464 256.663
R655 B.n665 B.n464 256.663
R656 B.n667 B.n464 256.663
R657 B.n673 B.n464 256.663
R658 B.n675 B.n464 256.663
R659 B.n681 B.n464 256.663
R660 B.n683 B.n464 256.663
R661 B.n689 B.n464 256.663
R662 B.n691 B.n464 256.663
R663 B.n697 B.n464 256.663
R664 B.n699 B.n464 256.663
R665 B.n705 B.n464 256.663
R666 B.n707 B.n464 256.663
R667 B.n713 B.n464 256.663
R668 B.n715 B.n464 256.663
R669 B.n721 B.n464 256.663
R670 B.n723 B.n464 256.663
R671 B.n729 B.n464 256.663
R672 B.n731 B.n464 256.663
R673 B.n737 B.n464 256.663
R674 B.n739 B.n464 256.663
R675 B.n745 B.n464 256.663
R676 B.n747 B.n464 256.663
R677 B.n753 B.n464 256.663
R678 B.n755 B.n464 256.663
R679 B.n761 B.n464 256.663
R680 B.n763 B.n464 256.663
R681 B.n769 B.n464 256.663
R682 B.n771 B.n464 256.663
R683 B.n777 B.n464 256.663
R684 B.n779 B.n464 256.663
R685 B.n785 B.n464 256.663
R686 B.n787 B.n464 256.663
R687 B.n793 B.n464 256.663
R688 B.n795 B.n464 256.663
R689 B.n801 B.n464 256.663
R690 B.n804 B.n464 256.663
R691 B.n811 B.n461 163.367
R692 B.n815 B.n461 163.367
R693 B.n815 B.n455 163.367
R694 B.n823 B.n455 163.367
R695 B.n823 B.n453 163.367
R696 B.n827 B.n453 163.367
R697 B.n827 B.n447 163.367
R698 B.n836 B.n447 163.367
R699 B.n836 B.n445 163.367
R700 B.n840 B.n445 163.367
R701 B.n840 B.n440 163.367
R702 B.n848 B.n440 163.367
R703 B.n848 B.n438 163.367
R704 B.n852 B.n438 163.367
R705 B.n852 B.n432 163.367
R706 B.n860 B.n432 163.367
R707 B.n860 B.n430 163.367
R708 B.n864 B.n430 163.367
R709 B.n864 B.n424 163.367
R710 B.n872 B.n424 163.367
R711 B.n872 B.n422 163.367
R712 B.n876 B.n422 163.367
R713 B.n876 B.n416 163.367
R714 B.n884 B.n416 163.367
R715 B.n884 B.n414 163.367
R716 B.n888 B.n414 163.367
R717 B.n888 B.n408 163.367
R718 B.n897 B.n408 163.367
R719 B.n897 B.n406 163.367
R720 B.n901 B.n406 163.367
R721 B.n901 B.n2 163.367
R722 B.n1016 B.n2 163.367
R723 B.n1016 B.n3 163.367
R724 B.n1012 B.n3 163.367
R725 B.n1012 B.n9 163.367
R726 B.n1008 B.n9 163.367
R727 B.n1008 B.n11 163.367
R728 B.n1004 B.n11 163.367
R729 B.n1004 B.n16 163.367
R730 B.n1000 B.n16 163.367
R731 B.n1000 B.n18 163.367
R732 B.n996 B.n18 163.367
R733 B.n996 B.n23 163.367
R734 B.n992 B.n23 163.367
R735 B.n992 B.n25 163.367
R736 B.n988 B.n25 163.367
R737 B.n988 B.n30 163.367
R738 B.n984 B.n30 163.367
R739 B.n984 B.n32 163.367
R740 B.n980 B.n32 163.367
R741 B.n980 B.n37 163.367
R742 B.n976 B.n37 163.367
R743 B.n976 B.n39 163.367
R744 B.n972 B.n39 163.367
R745 B.n972 B.n43 163.367
R746 B.n968 B.n43 163.367
R747 B.n968 B.n45 163.367
R748 B.n964 B.n45 163.367
R749 B.n964 B.n51 163.367
R750 B.n960 B.n51 163.367
R751 B.n960 B.n53 163.367
R752 B.n956 B.n53 163.367
R753 B.n956 B.n58 163.367
R754 B.n952 B.n58 163.367
R755 B.n539 B.n537 163.367
R756 B.n543 B.n537 163.367
R757 B.n547 B.n545 163.367
R758 B.n551 B.n535 163.367
R759 B.n555 B.n553 163.367
R760 B.n559 B.n533 163.367
R761 B.n563 B.n561 163.367
R762 B.n567 B.n531 163.367
R763 B.n571 B.n569 163.367
R764 B.n575 B.n529 163.367
R765 B.n579 B.n577 163.367
R766 B.n583 B.n527 163.367
R767 B.n587 B.n585 163.367
R768 B.n591 B.n525 163.367
R769 B.n595 B.n593 163.367
R770 B.n599 B.n523 163.367
R771 B.n603 B.n601 163.367
R772 B.n607 B.n521 163.367
R773 B.n611 B.n609 163.367
R774 B.n615 B.n519 163.367
R775 B.n619 B.n617 163.367
R776 B.n623 B.n517 163.367
R777 B.n627 B.n625 163.367
R778 B.n631 B.n515 163.367
R779 B.n635 B.n633 163.367
R780 B.n639 B.n513 163.367
R781 B.n643 B.n641 163.367
R782 B.n647 B.n511 163.367
R783 B.n651 B.n649 163.367
R784 B.n655 B.n509 163.367
R785 B.n659 B.n657 163.367
R786 B.n664 B.n505 163.367
R787 B.n668 B.n666 163.367
R788 B.n672 B.n503 163.367
R789 B.n676 B.n674 163.367
R790 B.n680 B.n501 163.367
R791 B.n684 B.n682 163.367
R792 B.n688 B.n496 163.367
R793 B.n692 B.n690 163.367
R794 B.n696 B.n494 163.367
R795 B.n700 B.n698 163.367
R796 B.n704 B.n492 163.367
R797 B.n708 B.n706 163.367
R798 B.n712 B.n490 163.367
R799 B.n716 B.n714 163.367
R800 B.n720 B.n488 163.367
R801 B.n724 B.n722 163.367
R802 B.n728 B.n486 163.367
R803 B.n732 B.n730 163.367
R804 B.n736 B.n484 163.367
R805 B.n740 B.n738 163.367
R806 B.n744 B.n482 163.367
R807 B.n748 B.n746 163.367
R808 B.n752 B.n480 163.367
R809 B.n756 B.n754 163.367
R810 B.n760 B.n478 163.367
R811 B.n764 B.n762 163.367
R812 B.n768 B.n476 163.367
R813 B.n772 B.n770 163.367
R814 B.n776 B.n474 163.367
R815 B.n780 B.n778 163.367
R816 B.n784 B.n472 163.367
R817 B.n788 B.n786 163.367
R818 B.n792 B.n470 163.367
R819 B.n796 B.n794 163.367
R820 B.n800 B.n468 163.367
R821 B.n803 B.n802 163.367
R822 B.n805 B.n465 163.367
R823 B.n809 B.n459 163.367
R824 B.n817 B.n459 163.367
R825 B.n817 B.n457 163.367
R826 B.n821 B.n457 163.367
R827 B.n821 B.n451 163.367
R828 B.n829 B.n451 163.367
R829 B.n829 B.n449 163.367
R830 B.n833 B.n449 163.367
R831 B.n833 B.n444 163.367
R832 B.n842 B.n444 163.367
R833 B.n842 B.n442 163.367
R834 B.n846 B.n442 163.367
R835 B.n846 B.n436 163.367
R836 B.n854 B.n436 163.367
R837 B.n854 B.n434 163.367
R838 B.n858 B.n434 163.367
R839 B.n858 B.n428 163.367
R840 B.n866 B.n428 163.367
R841 B.n866 B.n426 163.367
R842 B.n870 B.n426 163.367
R843 B.n870 B.n420 163.367
R844 B.n878 B.n420 163.367
R845 B.n878 B.n418 163.367
R846 B.n882 B.n418 163.367
R847 B.n882 B.n412 163.367
R848 B.n890 B.n412 163.367
R849 B.n890 B.n410 163.367
R850 B.n895 B.n410 163.367
R851 B.n895 B.n404 163.367
R852 B.n903 B.n404 163.367
R853 B.n904 B.n903 163.367
R854 B.n904 B.n5 163.367
R855 B.n6 B.n5 163.367
R856 B.n7 B.n6 163.367
R857 B.n909 B.n7 163.367
R858 B.n909 B.n12 163.367
R859 B.n13 B.n12 163.367
R860 B.n14 B.n13 163.367
R861 B.n914 B.n14 163.367
R862 B.n914 B.n19 163.367
R863 B.n20 B.n19 163.367
R864 B.n21 B.n20 163.367
R865 B.n919 B.n21 163.367
R866 B.n919 B.n26 163.367
R867 B.n27 B.n26 163.367
R868 B.n28 B.n27 163.367
R869 B.n924 B.n28 163.367
R870 B.n924 B.n33 163.367
R871 B.n34 B.n33 163.367
R872 B.n35 B.n34 163.367
R873 B.n929 B.n35 163.367
R874 B.n929 B.n40 163.367
R875 B.n41 B.n40 163.367
R876 B.n42 B.n41 163.367
R877 B.n934 B.n42 163.367
R878 B.n934 B.n47 163.367
R879 B.n48 B.n47 163.367
R880 B.n49 B.n48 163.367
R881 B.n939 B.n49 163.367
R882 B.n939 B.n54 163.367
R883 B.n55 B.n54 163.367
R884 B.n56 B.n55 163.367
R885 B.n944 B.n56 163.367
R886 B.n944 B.n61 163.367
R887 B.n136 B.n135 163.367
R888 B.n140 B.n139 163.367
R889 B.n144 B.n143 163.367
R890 B.n148 B.n147 163.367
R891 B.n152 B.n151 163.367
R892 B.n156 B.n155 163.367
R893 B.n160 B.n159 163.367
R894 B.n164 B.n163 163.367
R895 B.n168 B.n167 163.367
R896 B.n172 B.n171 163.367
R897 B.n176 B.n175 163.367
R898 B.n180 B.n179 163.367
R899 B.n184 B.n183 163.367
R900 B.n188 B.n187 163.367
R901 B.n192 B.n191 163.367
R902 B.n196 B.n195 163.367
R903 B.n200 B.n199 163.367
R904 B.n204 B.n203 163.367
R905 B.n208 B.n207 163.367
R906 B.n212 B.n211 163.367
R907 B.n216 B.n215 163.367
R908 B.n220 B.n219 163.367
R909 B.n224 B.n223 163.367
R910 B.n228 B.n227 163.367
R911 B.n232 B.n231 163.367
R912 B.n236 B.n235 163.367
R913 B.n240 B.n239 163.367
R914 B.n244 B.n243 163.367
R915 B.n248 B.n247 163.367
R916 B.n252 B.n251 163.367
R917 B.n256 B.n255 163.367
R918 B.n261 B.n260 163.367
R919 B.n265 B.n264 163.367
R920 B.n269 B.n268 163.367
R921 B.n273 B.n272 163.367
R922 B.n277 B.n276 163.367
R923 B.n282 B.n281 163.367
R924 B.n286 B.n285 163.367
R925 B.n290 B.n289 163.367
R926 B.n294 B.n293 163.367
R927 B.n298 B.n297 163.367
R928 B.n302 B.n301 163.367
R929 B.n306 B.n305 163.367
R930 B.n310 B.n309 163.367
R931 B.n314 B.n313 163.367
R932 B.n318 B.n317 163.367
R933 B.n322 B.n321 163.367
R934 B.n326 B.n325 163.367
R935 B.n330 B.n329 163.367
R936 B.n334 B.n333 163.367
R937 B.n338 B.n337 163.367
R938 B.n342 B.n341 163.367
R939 B.n346 B.n345 163.367
R940 B.n350 B.n349 163.367
R941 B.n354 B.n353 163.367
R942 B.n358 B.n357 163.367
R943 B.n362 B.n361 163.367
R944 B.n366 B.n365 163.367
R945 B.n370 B.n369 163.367
R946 B.n374 B.n373 163.367
R947 B.n378 B.n377 163.367
R948 B.n382 B.n381 163.367
R949 B.n386 B.n385 163.367
R950 B.n390 B.n389 163.367
R951 B.n394 B.n393 163.367
R952 B.n398 B.n397 163.367
R953 B.n400 B.n129 163.367
R954 B.n497 B.t12 151.15
R955 B.n130 B.t4 151.15
R956 B.n506 B.t9 151.125
R957 B.n132 B.t14 151.125
R958 B.n498 B.n497 78.1581
R959 B.n507 B.n506 78.1581
R960 B.n133 B.n132 78.1581
R961 B.n131 B.n130 78.1581
R962 B.n498 B.t11 72.9924
R963 B.n131 B.t5 72.9924
R964 B.n507 B.t8 72.9666
R965 B.n133 B.t15 72.9666
R966 B.n538 B.n463 71.676
R967 B.n544 B.n543 71.676
R968 B.n547 B.n546 71.676
R969 B.n552 B.n551 71.676
R970 B.n555 B.n554 71.676
R971 B.n560 B.n559 71.676
R972 B.n563 B.n562 71.676
R973 B.n568 B.n567 71.676
R974 B.n571 B.n570 71.676
R975 B.n576 B.n575 71.676
R976 B.n579 B.n578 71.676
R977 B.n584 B.n583 71.676
R978 B.n587 B.n586 71.676
R979 B.n592 B.n591 71.676
R980 B.n595 B.n594 71.676
R981 B.n600 B.n599 71.676
R982 B.n603 B.n602 71.676
R983 B.n608 B.n607 71.676
R984 B.n611 B.n610 71.676
R985 B.n616 B.n615 71.676
R986 B.n619 B.n618 71.676
R987 B.n624 B.n623 71.676
R988 B.n627 B.n626 71.676
R989 B.n632 B.n631 71.676
R990 B.n635 B.n634 71.676
R991 B.n640 B.n639 71.676
R992 B.n643 B.n642 71.676
R993 B.n648 B.n647 71.676
R994 B.n651 B.n650 71.676
R995 B.n656 B.n655 71.676
R996 B.n659 B.n658 71.676
R997 B.n665 B.n664 71.676
R998 B.n668 B.n667 71.676
R999 B.n673 B.n672 71.676
R1000 B.n676 B.n675 71.676
R1001 B.n681 B.n680 71.676
R1002 B.n684 B.n683 71.676
R1003 B.n689 B.n688 71.676
R1004 B.n692 B.n691 71.676
R1005 B.n697 B.n696 71.676
R1006 B.n700 B.n699 71.676
R1007 B.n705 B.n704 71.676
R1008 B.n708 B.n707 71.676
R1009 B.n713 B.n712 71.676
R1010 B.n716 B.n715 71.676
R1011 B.n721 B.n720 71.676
R1012 B.n724 B.n723 71.676
R1013 B.n729 B.n728 71.676
R1014 B.n732 B.n731 71.676
R1015 B.n737 B.n736 71.676
R1016 B.n740 B.n739 71.676
R1017 B.n745 B.n744 71.676
R1018 B.n748 B.n747 71.676
R1019 B.n753 B.n752 71.676
R1020 B.n756 B.n755 71.676
R1021 B.n761 B.n760 71.676
R1022 B.n764 B.n763 71.676
R1023 B.n769 B.n768 71.676
R1024 B.n772 B.n771 71.676
R1025 B.n777 B.n776 71.676
R1026 B.n780 B.n779 71.676
R1027 B.n785 B.n784 71.676
R1028 B.n788 B.n787 71.676
R1029 B.n793 B.n792 71.676
R1030 B.n796 B.n795 71.676
R1031 B.n801 B.n800 71.676
R1032 B.n804 B.n803 71.676
R1033 B.n62 B.n60 71.676
R1034 B.n136 B.n63 71.676
R1035 B.n140 B.n64 71.676
R1036 B.n144 B.n65 71.676
R1037 B.n148 B.n66 71.676
R1038 B.n152 B.n67 71.676
R1039 B.n156 B.n68 71.676
R1040 B.n160 B.n69 71.676
R1041 B.n164 B.n70 71.676
R1042 B.n168 B.n71 71.676
R1043 B.n172 B.n72 71.676
R1044 B.n176 B.n73 71.676
R1045 B.n180 B.n74 71.676
R1046 B.n184 B.n75 71.676
R1047 B.n188 B.n76 71.676
R1048 B.n192 B.n77 71.676
R1049 B.n196 B.n78 71.676
R1050 B.n200 B.n79 71.676
R1051 B.n204 B.n80 71.676
R1052 B.n208 B.n81 71.676
R1053 B.n212 B.n82 71.676
R1054 B.n216 B.n83 71.676
R1055 B.n220 B.n84 71.676
R1056 B.n224 B.n85 71.676
R1057 B.n228 B.n86 71.676
R1058 B.n232 B.n87 71.676
R1059 B.n236 B.n88 71.676
R1060 B.n240 B.n89 71.676
R1061 B.n244 B.n90 71.676
R1062 B.n248 B.n91 71.676
R1063 B.n252 B.n92 71.676
R1064 B.n256 B.n93 71.676
R1065 B.n261 B.n94 71.676
R1066 B.n265 B.n95 71.676
R1067 B.n269 B.n96 71.676
R1068 B.n273 B.n97 71.676
R1069 B.n277 B.n98 71.676
R1070 B.n282 B.n99 71.676
R1071 B.n286 B.n100 71.676
R1072 B.n290 B.n101 71.676
R1073 B.n294 B.n102 71.676
R1074 B.n298 B.n103 71.676
R1075 B.n302 B.n104 71.676
R1076 B.n306 B.n105 71.676
R1077 B.n310 B.n106 71.676
R1078 B.n314 B.n107 71.676
R1079 B.n318 B.n108 71.676
R1080 B.n322 B.n109 71.676
R1081 B.n326 B.n110 71.676
R1082 B.n330 B.n111 71.676
R1083 B.n334 B.n112 71.676
R1084 B.n338 B.n113 71.676
R1085 B.n342 B.n114 71.676
R1086 B.n346 B.n115 71.676
R1087 B.n350 B.n116 71.676
R1088 B.n354 B.n117 71.676
R1089 B.n358 B.n118 71.676
R1090 B.n362 B.n119 71.676
R1091 B.n366 B.n120 71.676
R1092 B.n370 B.n121 71.676
R1093 B.n374 B.n122 71.676
R1094 B.n378 B.n123 71.676
R1095 B.n382 B.n124 71.676
R1096 B.n386 B.n125 71.676
R1097 B.n390 B.n126 71.676
R1098 B.n394 B.n127 71.676
R1099 B.n398 B.n128 71.676
R1100 B.n949 B.n129 71.676
R1101 B.n949 B.n948 71.676
R1102 B.n400 B.n128 71.676
R1103 B.n397 B.n127 71.676
R1104 B.n393 B.n126 71.676
R1105 B.n389 B.n125 71.676
R1106 B.n385 B.n124 71.676
R1107 B.n381 B.n123 71.676
R1108 B.n377 B.n122 71.676
R1109 B.n373 B.n121 71.676
R1110 B.n369 B.n120 71.676
R1111 B.n365 B.n119 71.676
R1112 B.n361 B.n118 71.676
R1113 B.n357 B.n117 71.676
R1114 B.n353 B.n116 71.676
R1115 B.n349 B.n115 71.676
R1116 B.n345 B.n114 71.676
R1117 B.n341 B.n113 71.676
R1118 B.n337 B.n112 71.676
R1119 B.n333 B.n111 71.676
R1120 B.n329 B.n110 71.676
R1121 B.n325 B.n109 71.676
R1122 B.n321 B.n108 71.676
R1123 B.n317 B.n107 71.676
R1124 B.n313 B.n106 71.676
R1125 B.n309 B.n105 71.676
R1126 B.n305 B.n104 71.676
R1127 B.n301 B.n103 71.676
R1128 B.n297 B.n102 71.676
R1129 B.n293 B.n101 71.676
R1130 B.n289 B.n100 71.676
R1131 B.n285 B.n99 71.676
R1132 B.n281 B.n98 71.676
R1133 B.n276 B.n97 71.676
R1134 B.n272 B.n96 71.676
R1135 B.n268 B.n95 71.676
R1136 B.n264 B.n94 71.676
R1137 B.n260 B.n93 71.676
R1138 B.n255 B.n92 71.676
R1139 B.n251 B.n91 71.676
R1140 B.n247 B.n90 71.676
R1141 B.n243 B.n89 71.676
R1142 B.n239 B.n88 71.676
R1143 B.n235 B.n87 71.676
R1144 B.n231 B.n86 71.676
R1145 B.n227 B.n85 71.676
R1146 B.n223 B.n84 71.676
R1147 B.n219 B.n83 71.676
R1148 B.n215 B.n82 71.676
R1149 B.n211 B.n81 71.676
R1150 B.n207 B.n80 71.676
R1151 B.n203 B.n79 71.676
R1152 B.n199 B.n78 71.676
R1153 B.n195 B.n77 71.676
R1154 B.n191 B.n76 71.676
R1155 B.n187 B.n75 71.676
R1156 B.n183 B.n74 71.676
R1157 B.n179 B.n73 71.676
R1158 B.n175 B.n72 71.676
R1159 B.n171 B.n71 71.676
R1160 B.n167 B.n70 71.676
R1161 B.n163 B.n69 71.676
R1162 B.n159 B.n68 71.676
R1163 B.n155 B.n67 71.676
R1164 B.n151 B.n66 71.676
R1165 B.n147 B.n65 71.676
R1166 B.n143 B.n64 71.676
R1167 B.n139 B.n63 71.676
R1168 B.n135 B.n62 71.676
R1169 B.n539 B.n538 71.676
R1170 B.n545 B.n544 71.676
R1171 B.n546 B.n535 71.676
R1172 B.n553 B.n552 71.676
R1173 B.n554 B.n533 71.676
R1174 B.n561 B.n560 71.676
R1175 B.n562 B.n531 71.676
R1176 B.n569 B.n568 71.676
R1177 B.n570 B.n529 71.676
R1178 B.n577 B.n576 71.676
R1179 B.n578 B.n527 71.676
R1180 B.n585 B.n584 71.676
R1181 B.n586 B.n525 71.676
R1182 B.n593 B.n592 71.676
R1183 B.n594 B.n523 71.676
R1184 B.n601 B.n600 71.676
R1185 B.n602 B.n521 71.676
R1186 B.n609 B.n608 71.676
R1187 B.n610 B.n519 71.676
R1188 B.n617 B.n616 71.676
R1189 B.n618 B.n517 71.676
R1190 B.n625 B.n624 71.676
R1191 B.n626 B.n515 71.676
R1192 B.n633 B.n632 71.676
R1193 B.n634 B.n513 71.676
R1194 B.n641 B.n640 71.676
R1195 B.n642 B.n511 71.676
R1196 B.n649 B.n648 71.676
R1197 B.n650 B.n509 71.676
R1198 B.n657 B.n656 71.676
R1199 B.n658 B.n505 71.676
R1200 B.n666 B.n665 71.676
R1201 B.n667 B.n503 71.676
R1202 B.n674 B.n673 71.676
R1203 B.n675 B.n501 71.676
R1204 B.n682 B.n681 71.676
R1205 B.n683 B.n496 71.676
R1206 B.n690 B.n689 71.676
R1207 B.n691 B.n494 71.676
R1208 B.n698 B.n697 71.676
R1209 B.n699 B.n492 71.676
R1210 B.n706 B.n705 71.676
R1211 B.n707 B.n490 71.676
R1212 B.n714 B.n713 71.676
R1213 B.n715 B.n488 71.676
R1214 B.n722 B.n721 71.676
R1215 B.n723 B.n486 71.676
R1216 B.n730 B.n729 71.676
R1217 B.n731 B.n484 71.676
R1218 B.n738 B.n737 71.676
R1219 B.n739 B.n482 71.676
R1220 B.n746 B.n745 71.676
R1221 B.n747 B.n480 71.676
R1222 B.n754 B.n753 71.676
R1223 B.n755 B.n478 71.676
R1224 B.n762 B.n761 71.676
R1225 B.n763 B.n476 71.676
R1226 B.n770 B.n769 71.676
R1227 B.n771 B.n474 71.676
R1228 B.n778 B.n777 71.676
R1229 B.n779 B.n472 71.676
R1230 B.n786 B.n785 71.676
R1231 B.n787 B.n470 71.676
R1232 B.n794 B.n793 71.676
R1233 B.n795 B.n468 71.676
R1234 B.n802 B.n801 71.676
R1235 B.n805 B.n804 71.676
R1236 B.n499 B.n498 59.5399
R1237 B.n662 B.n507 59.5399
R1238 B.n258 B.n133 59.5399
R1239 B.n279 B.n131 59.5399
R1240 B.n810 B.n464 49.6044
R1241 B.n951 B.n950 49.6044
R1242 B.n953 B.n59 30.4395
R1243 B.n808 B.n807 30.4395
R1244 B.n812 B.n462 30.4395
R1245 B.n947 B.n946 30.4395
R1246 B.n810 B.n460 30.3885
R1247 B.n816 B.n460 30.3885
R1248 B.n816 B.n456 30.3885
R1249 B.n822 B.n456 30.3885
R1250 B.n822 B.n452 30.3885
R1251 B.n828 B.n452 30.3885
R1252 B.n828 B.n448 30.3885
R1253 B.n835 B.n448 30.3885
R1254 B.n835 B.n834 30.3885
R1255 B.n841 B.n441 30.3885
R1256 B.n847 B.n441 30.3885
R1257 B.n847 B.n437 30.3885
R1258 B.n853 B.n437 30.3885
R1259 B.n853 B.n433 30.3885
R1260 B.n859 B.n433 30.3885
R1261 B.n859 B.n429 30.3885
R1262 B.n865 B.n429 30.3885
R1263 B.n865 B.n425 30.3885
R1264 B.n871 B.n425 30.3885
R1265 B.n871 B.n421 30.3885
R1266 B.n877 B.n421 30.3885
R1267 B.n877 B.n417 30.3885
R1268 B.n883 B.n417 30.3885
R1269 B.n889 B.n413 30.3885
R1270 B.n889 B.n409 30.3885
R1271 B.n896 B.n409 30.3885
R1272 B.n896 B.n405 30.3885
R1273 B.n902 B.n405 30.3885
R1274 B.n902 B.n4 30.3885
R1275 B.n1015 B.n4 30.3885
R1276 B.n1015 B.n1014 30.3885
R1277 B.n1014 B.n1013 30.3885
R1278 B.n1013 B.n8 30.3885
R1279 B.n1007 B.n8 30.3885
R1280 B.n1007 B.n1006 30.3885
R1281 B.n1006 B.n1005 30.3885
R1282 B.n1005 B.n15 30.3885
R1283 B.n999 B.n998 30.3885
R1284 B.n998 B.n997 30.3885
R1285 B.n997 B.n22 30.3885
R1286 B.n991 B.n22 30.3885
R1287 B.n991 B.n990 30.3885
R1288 B.n990 B.n989 30.3885
R1289 B.n989 B.n29 30.3885
R1290 B.n983 B.n29 30.3885
R1291 B.n983 B.n982 30.3885
R1292 B.n982 B.n981 30.3885
R1293 B.n981 B.n36 30.3885
R1294 B.n975 B.n36 30.3885
R1295 B.n975 B.n974 30.3885
R1296 B.n974 B.n973 30.3885
R1297 B.n967 B.n46 30.3885
R1298 B.n967 B.n966 30.3885
R1299 B.n966 B.n965 30.3885
R1300 B.n965 B.n50 30.3885
R1301 B.n959 B.n50 30.3885
R1302 B.n959 B.n958 30.3885
R1303 B.n958 B.n957 30.3885
R1304 B.n957 B.n57 30.3885
R1305 B.n951 B.n57 30.3885
R1306 B B.n1017 18.0485
R1307 B.n841 B.t7 17.8758
R1308 B.n973 B.t3 17.8758
R1309 B.t1 B.n413 16.0883
R1310 B.t0 B.n15 16.0883
R1311 B.n883 B.t1 14.3007
R1312 B.n999 B.t0 14.3007
R1313 B.n834 B.t7 12.5132
R1314 B.n46 B.t3 12.5132
R1315 B.n134 B.n59 10.6151
R1316 B.n137 B.n134 10.6151
R1317 B.n138 B.n137 10.6151
R1318 B.n141 B.n138 10.6151
R1319 B.n142 B.n141 10.6151
R1320 B.n145 B.n142 10.6151
R1321 B.n146 B.n145 10.6151
R1322 B.n149 B.n146 10.6151
R1323 B.n150 B.n149 10.6151
R1324 B.n153 B.n150 10.6151
R1325 B.n154 B.n153 10.6151
R1326 B.n157 B.n154 10.6151
R1327 B.n158 B.n157 10.6151
R1328 B.n161 B.n158 10.6151
R1329 B.n162 B.n161 10.6151
R1330 B.n165 B.n162 10.6151
R1331 B.n166 B.n165 10.6151
R1332 B.n169 B.n166 10.6151
R1333 B.n170 B.n169 10.6151
R1334 B.n173 B.n170 10.6151
R1335 B.n174 B.n173 10.6151
R1336 B.n177 B.n174 10.6151
R1337 B.n178 B.n177 10.6151
R1338 B.n181 B.n178 10.6151
R1339 B.n182 B.n181 10.6151
R1340 B.n185 B.n182 10.6151
R1341 B.n186 B.n185 10.6151
R1342 B.n189 B.n186 10.6151
R1343 B.n190 B.n189 10.6151
R1344 B.n193 B.n190 10.6151
R1345 B.n194 B.n193 10.6151
R1346 B.n197 B.n194 10.6151
R1347 B.n198 B.n197 10.6151
R1348 B.n201 B.n198 10.6151
R1349 B.n202 B.n201 10.6151
R1350 B.n205 B.n202 10.6151
R1351 B.n206 B.n205 10.6151
R1352 B.n209 B.n206 10.6151
R1353 B.n210 B.n209 10.6151
R1354 B.n213 B.n210 10.6151
R1355 B.n214 B.n213 10.6151
R1356 B.n217 B.n214 10.6151
R1357 B.n218 B.n217 10.6151
R1358 B.n221 B.n218 10.6151
R1359 B.n222 B.n221 10.6151
R1360 B.n225 B.n222 10.6151
R1361 B.n226 B.n225 10.6151
R1362 B.n229 B.n226 10.6151
R1363 B.n230 B.n229 10.6151
R1364 B.n233 B.n230 10.6151
R1365 B.n234 B.n233 10.6151
R1366 B.n237 B.n234 10.6151
R1367 B.n238 B.n237 10.6151
R1368 B.n241 B.n238 10.6151
R1369 B.n242 B.n241 10.6151
R1370 B.n245 B.n242 10.6151
R1371 B.n246 B.n245 10.6151
R1372 B.n249 B.n246 10.6151
R1373 B.n250 B.n249 10.6151
R1374 B.n253 B.n250 10.6151
R1375 B.n254 B.n253 10.6151
R1376 B.n257 B.n254 10.6151
R1377 B.n262 B.n259 10.6151
R1378 B.n263 B.n262 10.6151
R1379 B.n266 B.n263 10.6151
R1380 B.n267 B.n266 10.6151
R1381 B.n270 B.n267 10.6151
R1382 B.n271 B.n270 10.6151
R1383 B.n274 B.n271 10.6151
R1384 B.n275 B.n274 10.6151
R1385 B.n278 B.n275 10.6151
R1386 B.n283 B.n280 10.6151
R1387 B.n284 B.n283 10.6151
R1388 B.n287 B.n284 10.6151
R1389 B.n288 B.n287 10.6151
R1390 B.n291 B.n288 10.6151
R1391 B.n292 B.n291 10.6151
R1392 B.n295 B.n292 10.6151
R1393 B.n296 B.n295 10.6151
R1394 B.n299 B.n296 10.6151
R1395 B.n300 B.n299 10.6151
R1396 B.n303 B.n300 10.6151
R1397 B.n304 B.n303 10.6151
R1398 B.n307 B.n304 10.6151
R1399 B.n308 B.n307 10.6151
R1400 B.n311 B.n308 10.6151
R1401 B.n312 B.n311 10.6151
R1402 B.n315 B.n312 10.6151
R1403 B.n316 B.n315 10.6151
R1404 B.n319 B.n316 10.6151
R1405 B.n320 B.n319 10.6151
R1406 B.n323 B.n320 10.6151
R1407 B.n324 B.n323 10.6151
R1408 B.n327 B.n324 10.6151
R1409 B.n328 B.n327 10.6151
R1410 B.n331 B.n328 10.6151
R1411 B.n332 B.n331 10.6151
R1412 B.n335 B.n332 10.6151
R1413 B.n336 B.n335 10.6151
R1414 B.n339 B.n336 10.6151
R1415 B.n340 B.n339 10.6151
R1416 B.n343 B.n340 10.6151
R1417 B.n344 B.n343 10.6151
R1418 B.n347 B.n344 10.6151
R1419 B.n348 B.n347 10.6151
R1420 B.n351 B.n348 10.6151
R1421 B.n352 B.n351 10.6151
R1422 B.n355 B.n352 10.6151
R1423 B.n356 B.n355 10.6151
R1424 B.n359 B.n356 10.6151
R1425 B.n360 B.n359 10.6151
R1426 B.n363 B.n360 10.6151
R1427 B.n364 B.n363 10.6151
R1428 B.n367 B.n364 10.6151
R1429 B.n368 B.n367 10.6151
R1430 B.n371 B.n368 10.6151
R1431 B.n372 B.n371 10.6151
R1432 B.n375 B.n372 10.6151
R1433 B.n376 B.n375 10.6151
R1434 B.n379 B.n376 10.6151
R1435 B.n380 B.n379 10.6151
R1436 B.n383 B.n380 10.6151
R1437 B.n384 B.n383 10.6151
R1438 B.n387 B.n384 10.6151
R1439 B.n388 B.n387 10.6151
R1440 B.n391 B.n388 10.6151
R1441 B.n392 B.n391 10.6151
R1442 B.n395 B.n392 10.6151
R1443 B.n396 B.n395 10.6151
R1444 B.n399 B.n396 10.6151
R1445 B.n401 B.n399 10.6151
R1446 B.n402 B.n401 10.6151
R1447 B.n947 B.n402 10.6151
R1448 B.n808 B.n458 10.6151
R1449 B.n818 B.n458 10.6151
R1450 B.n819 B.n818 10.6151
R1451 B.n820 B.n819 10.6151
R1452 B.n820 B.n450 10.6151
R1453 B.n830 B.n450 10.6151
R1454 B.n831 B.n830 10.6151
R1455 B.n832 B.n831 10.6151
R1456 B.n832 B.n443 10.6151
R1457 B.n843 B.n443 10.6151
R1458 B.n844 B.n843 10.6151
R1459 B.n845 B.n844 10.6151
R1460 B.n845 B.n435 10.6151
R1461 B.n855 B.n435 10.6151
R1462 B.n856 B.n855 10.6151
R1463 B.n857 B.n856 10.6151
R1464 B.n857 B.n427 10.6151
R1465 B.n867 B.n427 10.6151
R1466 B.n868 B.n867 10.6151
R1467 B.n869 B.n868 10.6151
R1468 B.n869 B.n419 10.6151
R1469 B.n879 B.n419 10.6151
R1470 B.n880 B.n879 10.6151
R1471 B.n881 B.n880 10.6151
R1472 B.n881 B.n411 10.6151
R1473 B.n891 B.n411 10.6151
R1474 B.n892 B.n891 10.6151
R1475 B.n894 B.n892 10.6151
R1476 B.n894 B.n893 10.6151
R1477 B.n893 B.n403 10.6151
R1478 B.n905 B.n403 10.6151
R1479 B.n906 B.n905 10.6151
R1480 B.n907 B.n906 10.6151
R1481 B.n908 B.n907 10.6151
R1482 B.n910 B.n908 10.6151
R1483 B.n911 B.n910 10.6151
R1484 B.n912 B.n911 10.6151
R1485 B.n913 B.n912 10.6151
R1486 B.n915 B.n913 10.6151
R1487 B.n916 B.n915 10.6151
R1488 B.n917 B.n916 10.6151
R1489 B.n918 B.n917 10.6151
R1490 B.n920 B.n918 10.6151
R1491 B.n921 B.n920 10.6151
R1492 B.n922 B.n921 10.6151
R1493 B.n923 B.n922 10.6151
R1494 B.n925 B.n923 10.6151
R1495 B.n926 B.n925 10.6151
R1496 B.n927 B.n926 10.6151
R1497 B.n928 B.n927 10.6151
R1498 B.n930 B.n928 10.6151
R1499 B.n931 B.n930 10.6151
R1500 B.n932 B.n931 10.6151
R1501 B.n933 B.n932 10.6151
R1502 B.n935 B.n933 10.6151
R1503 B.n936 B.n935 10.6151
R1504 B.n937 B.n936 10.6151
R1505 B.n938 B.n937 10.6151
R1506 B.n940 B.n938 10.6151
R1507 B.n941 B.n940 10.6151
R1508 B.n942 B.n941 10.6151
R1509 B.n943 B.n942 10.6151
R1510 B.n945 B.n943 10.6151
R1511 B.n946 B.n945 10.6151
R1512 B.n540 B.n462 10.6151
R1513 B.n541 B.n540 10.6151
R1514 B.n542 B.n541 10.6151
R1515 B.n542 B.n536 10.6151
R1516 B.n548 B.n536 10.6151
R1517 B.n549 B.n548 10.6151
R1518 B.n550 B.n549 10.6151
R1519 B.n550 B.n534 10.6151
R1520 B.n556 B.n534 10.6151
R1521 B.n557 B.n556 10.6151
R1522 B.n558 B.n557 10.6151
R1523 B.n558 B.n532 10.6151
R1524 B.n564 B.n532 10.6151
R1525 B.n565 B.n564 10.6151
R1526 B.n566 B.n565 10.6151
R1527 B.n566 B.n530 10.6151
R1528 B.n572 B.n530 10.6151
R1529 B.n573 B.n572 10.6151
R1530 B.n574 B.n573 10.6151
R1531 B.n574 B.n528 10.6151
R1532 B.n580 B.n528 10.6151
R1533 B.n581 B.n580 10.6151
R1534 B.n582 B.n581 10.6151
R1535 B.n582 B.n526 10.6151
R1536 B.n588 B.n526 10.6151
R1537 B.n589 B.n588 10.6151
R1538 B.n590 B.n589 10.6151
R1539 B.n590 B.n524 10.6151
R1540 B.n596 B.n524 10.6151
R1541 B.n597 B.n596 10.6151
R1542 B.n598 B.n597 10.6151
R1543 B.n598 B.n522 10.6151
R1544 B.n604 B.n522 10.6151
R1545 B.n605 B.n604 10.6151
R1546 B.n606 B.n605 10.6151
R1547 B.n606 B.n520 10.6151
R1548 B.n612 B.n520 10.6151
R1549 B.n613 B.n612 10.6151
R1550 B.n614 B.n613 10.6151
R1551 B.n614 B.n518 10.6151
R1552 B.n620 B.n518 10.6151
R1553 B.n621 B.n620 10.6151
R1554 B.n622 B.n621 10.6151
R1555 B.n622 B.n516 10.6151
R1556 B.n628 B.n516 10.6151
R1557 B.n629 B.n628 10.6151
R1558 B.n630 B.n629 10.6151
R1559 B.n630 B.n514 10.6151
R1560 B.n636 B.n514 10.6151
R1561 B.n637 B.n636 10.6151
R1562 B.n638 B.n637 10.6151
R1563 B.n638 B.n512 10.6151
R1564 B.n644 B.n512 10.6151
R1565 B.n645 B.n644 10.6151
R1566 B.n646 B.n645 10.6151
R1567 B.n646 B.n510 10.6151
R1568 B.n652 B.n510 10.6151
R1569 B.n653 B.n652 10.6151
R1570 B.n654 B.n653 10.6151
R1571 B.n654 B.n508 10.6151
R1572 B.n660 B.n508 10.6151
R1573 B.n661 B.n660 10.6151
R1574 B.n663 B.n504 10.6151
R1575 B.n669 B.n504 10.6151
R1576 B.n670 B.n669 10.6151
R1577 B.n671 B.n670 10.6151
R1578 B.n671 B.n502 10.6151
R1579 B.n677 B.n502 10.6151
R1580 B.n678 B.n677 10.6151
R1581 B.n679 B.n678 10.6151
R1582 B.n679 B.n500 10.6151
R1583 B.n686 B.n685 10.6151
R1584 B.n687 B.n686 10.6151
R1585 B.n687 B.n495 10.6151
R1586 B.n693 B.n495 10.6151
R1587 B.n694 B.n693 10.6151
R1588 B.n695 B.n694 10.6151
R1589 B.n695 B.n493 10.6151
R1590 B.n701 B.n493 10.6151
R1591 B.n702 B.n701 10.6151
R1592 B.n703 B.n702 10.6151
R1593 B.n703 B.n491 10.6151
R1594 B.n709 B.n491 10.6151
R1595 B.n710 B.n709 10.6151
R1596 B.n711 B.n710 10.6151
R1597 B.n711 B.n489 10.6151
R1598 B.n717 B.n489 10.6151
R1599 B.n718 B.n717 10.6151
R1600 B.n719 B.n718 10.6151
R1601 B.n719 B.n487 10.6151
R1602 B.n725 B.n487 10.6151
R1603 B.n726 B.n725 10.6151
R1604 B.n727 B.n726 10.6151
R1605 B.n727 B.n485 10.6151
R1606 B.n733 B.n485 10.6151
R1607 B.n734 B.n733 10.6151
R1608 B.n735 B.n734 10.6151
R1609 B.n735 B.n483 10.6151
R1610 B.n741 B.n483 10.6151
R1611 B.n742 B.n741 10.6151
R1612 B.n743 B.n742 10.6151
R1613 B.n743 B.n481 10.6151
R1614 B.n749 B.n481 10.6151
R1615 B.n750 B.n749 10.6151
R1616 B.n751 B.n750 10.6151
R1617 B.n751 B.n479 10.6151
R1618 B.n757 B.n479 10.6151
R1619 B.n758 B.n757 10.6151
R1620 B.n759 B.n758 10.6151
R1621 B.n759 B.n477 10.6151
R1622 B.n765 B.n477 10.6151
R1623 B.n766 B.n765 10.6151
R1624 B.n767 B.n766 10.6151
R1625 B.n767 B.n475 10.6151
R1626 B.n773 B.n475 10.6151
R1627 B.n774 B.n773 10.6151
R1628 B.n775 B.n774 10.6151
R1629 B.n775 B.n473 10.6151
R1630 B.n781 B.n473 10.6151
R1631 B.n782 B.n781 10.6151
R1632 B.n783 B.n782 10.6151
R1633 B.n783 B.n471 10.6151
R1634 B.n789 B.n471 10.6151
R1635 B.n790 B.n789 10.6151
R1636 B.n791 B.n790 10.6151
R1637 B.n791 B.n469 10.6151
R1638 B.n797 B.n469 10.6151
R1639 B.n798 B.n797 10.6151
R1640 B.n799 B.n798 10.6151
R1641 B.n799 B.n467 10.6151
R1642 B.n467 B.n466 10.6151
R1643 B.n806 B.n466 10.6151
R1644 B.n807 B.n806 10.6151
R1645 B.n813 B.n812 10.6151
R1646 B.n814 B.n813 10.6151
R1647 B.n814 B.n454 10.6151
R1648 B.n824 B.n454 10.6151
R1649 B.n825 B.n824 10.6151
R1650 B.n826 B.n825 10.6151
R1651 B.n826 B.n446 10.6151
R1652 B.n837 B.n446 10.6151
R1653 B.n838 B.n837 10.6151
R1654 B.n839 B.n838 10.6151
R1655 B.n839 B.n439 10.6151
R1656 B.n849 B.n439 10.6151
R1657 B.n850 B.n849 10.6151
R1658 B.n851 B.n850 10.6151
R1659 B.n851 B.n431 10.6151
R1660 B.n861 B.n431 10.6151
R1661 B.n862 B.n861 10.6151
R1662 B.n863 B.n862 10.6151
R1663 B.n863 B.n423 10.6151
R1664 B.n873 B.n423 10.6151
R1665 B.n874 B.n873 10.6151
R1666 B.n875 B.n874 10.6151
R1667 B.n875 B.n415 10.6151
R1668 B.n885 B.n415 10.6151
R1669 B.n886 B.n885 10.6151
R1670 B.n887 B.n886 10.6151
R1671 B.n887 B.n407 10.6151
R1672 B.n898 B.n407 10.6151
R1673 B.n899 B.n898 10.6151
R1674 B.n900 B.n899 10.6151
R1675 B.n900 B.n0 10.6151
R1676 B.n1011 B.n1 10.6151
R1677 B.n1011 B.n1010 10.6151
R1678 B.n1010 B.n1009 10.6151
R1679 B.n1009 B.n10 10.6151
R1680 B.n1003 B.n10 10.6151
R1681 B.n1003 B.n1002 10.6151
R1682 B.n1002 B.n1001 10.6151
R1683 B.n1001 B.n17 10.6151
R1684 B.n995 B.n17 10.6151
R1685 B.n995 B.n994 10.6151
R1686 B.n994 B.n993 10.6151
R1687 B.n993 B.n24 10.6151
R1688 B.n987 B.n24 10.6151
R1689 B.n987 B.n986 10.6151
R1690 B.n986 B.n985 10.6151
R1691 B.n985 B.n31 10.6151
R1692 B.n979 B.n31 10.6151
R1693 B.n979 B.n978 10.6151
R1694 B.n978 B.n977 10.6151
R1695 B.n977 B.n38 10.6151
R1696 B.n971 B.n38 10.6151
R1697 B.n971 B.n970 10.6151
R1698 B.n970 B.n969 10.6151
R1699 B.n969 B.n44 10.6151
R1700 B.n963 B.n44 10.6151
R1701 B.n963 B.n962 10.6151
R1702 B.n962 B.n961 10.6151
R1703 B.n961 B.n52 10.6151
R1704 B.n955 B.n52 10.6151
R1705 B.n955 B.n954 10.6151
R1706 B.n954 B.n953 10.6151
R1707 B.n258 B.n257 9.36635
R1708 B.n280 B.n279 9.36635
R1709 B.n662 B.n661 9.36635
R1710 B.n685 B.n499 9.36635
R1711 B.n1017 B.n0 2.81026
R1712 B.n1017 B.n1 2.81026
R1713 B.n259 B.n258 1.24928
R1714 B.n279 B.n278 1.24928
R1715 B.n663 B.n662 1.24928
R1716 B.n500 B.n499 1.24928
R1717 VP.n0 VP.t0 214.197
R1718 VP.n0 VP.t1 161.064
R1719 VP VP.n0 0.62124
R1720 VDD1 VDD1.t0 110.697
R1721 VDD1 VDD1.t1 62.9493
C0 VP VDD2 0.37959f
C1 VTAIL VDD1 7.12304f
C2 VN VDD1 0.148961f
C3 VDD2 VDD1 0.79587f
C4 VN VTAIL 3.92209f
C5 VP VDD1 4.76561f
C6 VTAIL VDD2 7.18075f
C7 VN VDD2 4.53756f
C8 VTAIL VP 3.93686f
C9 VN VP 7.331339f
C10 VDD2 B 6.144637f
C11 VDD1 B 10.03246f
C12 VTAIL B 10.909171f
C13 VN B 13.48288f
C14 VP B 8.267118f
C15 VDD1.t1 B 3.60521f
C16 VDD1.t0 B 4.46931f
C17 VP.t0 B 5.74192f
C18 VP.t1 B 4.9996f
C19 VP.n0 B 5.16208f
C20 VDD2.t1 B 4.3731f
C21 VDD2.t0 B 3.56269f
C22 VDD2.n0 B 3.59239f
C23 VTAIL.t1 B 3.45037f
C24 VTAIL.n0 B 2.13366f
C25 VTAIL.t3 B 3.45037f
C26 VTAIL.n1 B 2.18527f
C27 VTAIL.t0 B 3.45037f
C28 VTAIL.n2 B 1.96399f
C29 VTAIL.t2 B 3.45037f
C30 VTAIL.n3 B 1.87504f
C31 VN.t0 B 4.9017f
C32 VN.t1 B 5.62064f
.ends

