* NGSPICE file created from diff_pair_sample_1778.ext - technology: sky130A

.subckt diff_pair_sample_1778 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t10 w_n3482_n3776# sky130_fd_pr__pfet_01v8 ad=2.3166 pd=14.37 as=5.4756 ps=28.86 w=14.04 l=2.81
X1 VDD2.t5 VN.t0 VTAIL.t1 w_n3482_n3776# sky130_fd_pr__pfet_01v8 ad=2.3166 pd=14.37 as=5.4756 ps=28.86 w=14.04 l=2.81
X2 VDD1.t4 VP.t1 VTAIL.t8 w_n3482_n3776# sky130_fd_pr__pfet_01v8 ad=2.3166 pd=14.37 as=5.4756 ps=28.86 w=14.04 l=2.81
X3 B.t11 B.t9 B.t10 w_n3482_n3776# sky130_fd_pr__pfet_01v8 ad=5.4756 pd=28.86 as=0 ps=0 w=14.04 l=2.81
X4 VDD2.t4 VN.t1 VTAIL.t5 w_n3482_n3776# sky130_fd_pr__pfet_01v8 ad=5.4756 pd=28.86 as=2.3166 ps=14.37 w=14.04 l=2.81
X5 VDD2.t3 VN.t2 VTAIL.t2 w_n3482_n3776# sky130_fd_pr__pfet_01v8 ad=2.3166 pd=14.37 as=5.4756 ps=28.86 w=14.04 l=2.81
X6 B.t8 B.t6 B.t7 w_n3482_n3776# sky130_fd_pr__pfet_01v8 ad=5.4756 pd=28.86 as=0 ps=0 w=14.04 l=2.81
X7 VTAIL.t3 VN.t3 VDD2.t2 w_n3482_n3776# sky130_fd_pr__pfet_01v8 ad=2.3166 pd=14.37 as=2.3166 ps=14.37 w=14.04 l=2.81
X8 VTAIL.t11 VP.t2 VDD1.t3 w_n3482_n3776# sky130_fd_pr__pfet_01v8 ad=2.3166 pd=14.37 as=2.3166 ps=14.37 w=14.04 l=2.81
X9 B.t5 B.t3 B.t4 w_n3482_n3776# sky130_fd_pr__pfet_01v8 ad=5.4756 pd=28.86 as=0 ps=0 w=14.04 l=2.81
X10 VTAIL.t4 VN.t4 VDD2.t1 w_n3482_n3776# sky130_fd_pr__pfet_01v8 ad=2.3166 pd=14.37 as=2.3166 ps=14.37 w=14.04 l=2.81
X11 VDD2.t0 VN.t5 VTAIL.t0 w_n3482_n3776# sky130_fd_pr__pfet_01v8 ad=5.4756 pd=28.86 as=2.3166 ps=14.37 w=14.04 l=2.81
X12 B.t2 B.t0 B.t1 w_n3482_n3776# sky130_fd_pr__pfet_01v8 ad=5.4756 pd=28.86 as=0 ps=0 w=14.04 l=2.81
X13 VTAIL.t6 VP.t3 VDD1.t2 w_n3482_n3776# sky130_fd_pr__pfet_01v8 ad=2.3166 pd=14.37 as=2.3166 ps=14.37 w=14.04 l=2.81
X14 VDD1.t1 VP.t4 VTAIL.t7 w_n3482_n3776# sky130_fd_pr__pfet_01v8 ad=5.4756 pd=28.86 as=2.3166 ps=14.37 w=14.04 l=2.81
X15 VDD1.t0 VP.t5 VTAIL.t9 w_n3482_n3776# sky130_fd_pr__pfet_01v8 ad=5.4756 pd=28.86 as=2.3166 ps=14.37 w=14.04 l=2.81
R0 VP.n13 VP.n12 161.3
R1 VP.n14 VP.n9 161.3
R2 VP.n16 VP.n15 161.3
R3 VP.n17 VP.n8 161.3
R4 VP.n19 VP.n18 161.3
R5 VP.n20 VP.n7 161.3
R6 VP.n43 VP.n0 161.3
R7 VP.n42 VP.n41 161.3
R8 VP.n40 VP.n1 161.3
R9 VP.n39 VP.n38 161.3
R10 VP.n37 VP.n2 161.3
R11 VP.n36 VP.n35 161.3
R12 VP.n34 VP.n3 161.3
R13 VP.n33 VP.n32 161.3
R14 VP.n31 VP.n4 161.3
R15 VP.n30 VP.n29 161.3
R16 VP.n28 VP.n5 161.3
R17 VP.n27 VP.n26 161.3
R18 VP.n25 VP.n6 161.3
R19 VP.n11 VP.t4 155.148
R20 VP.n3 VP.t2 120.415
R21 VP.n24 VP.t5 120.415
R22 VP.n44 VP.t1 120.415
R23 VP.n10 VP.t3 120.415
R24 VP.n21 VP.t0 120.415
R25 VP.n24 VP.n23 104.022
R26 VP.n45 VP.n44 104.022
R27 VP.n22 VP.n21 104.022
R28 VP.n23 VP.n22 51.0678
R29 VP.n11 VP.n10 49.0208
R30 VP.n30 VP.n5 47.3584
R31 VP.n38 VP.n1 47.3584
R32 VP.n15 VP.n8 47.3584
R33 VP.n31 VP.n30 33.7956
R34 VP.n38 VP.n37 33.7956
R35 VP.n15 VP.n14 33.7956
R36 VP.n26 VP.n25 24.5923
R37 VP.n26 VP.n5 24.5923
R38 VP.n32 VP.n31 24.5923
R39 VP.n32 VP.n3 24.5923
R40 VP.n36 VP.n3 24.5923
R41 VP.n37 VP.n36 24.5923
R42 VP.n42 VP.n1 24.5923
R43 VP.n43 VP.n42 24.5923
R44 VP.n19 VP.n8 24.5923
R45 VP.n20 VP.n19 24.5923
R46 VP.n13 VP.n10 24.5923
R47 VP.n14 VP.n13 24.5923
R48 VP.n25 VP.n24 6.88621
R49 VP.n44 VP.n43 6.88621
R50 VP.n21 VP.n20 6.88621
R51 VP.n12 VP.n11 4.88317
R52 VP.n22 VP.n7 0.278335
R53 VP.n23 VP.n6 0.278335
R54 VP.n45 VP.n0 0.278335
R55 VP.n12 VP.n9 0.189894
R56 VP.n16 VP.n9 0.189894
R57 VP.n17 VP.n16 0.189894
R58 VP.n18 VP.n17 0.189894
R59 VP.n18 VP.n7 0.189894
R60 VP.n27 VP.n6 0.189894
R61 VP.n28 VP.n27 0.189894
R62 VP.n29 VP.n28 0.189894
R63 VP.n29 VP.n4 0.189894
R64 VP.n33 VP.n4 0.189894
R65 VP.n34 VP.n33 0.189894
R66 VP.n35 VP.n34 0.189894
R67 VP.n35 VP.n2 0.189894
R68 VP.n39 VP.n2 0.189894
R69 VP.n40 VP.n39 0.189894
R70 VP.n41 VP.n40 0.189894
R71 VP.n41 VP.n0 0.189894
R72 VP VP.n45 0.153485
R73 VTAIL.n314 VTAIL.n242 756.745
R74 VTAIL.n74 VTAIL.n2 756.745
R75 VTAIL.n236 VTAIL.n164 756.745
R76 VTAIL.n156 VTAIL.n84 756.745
R77 VTAIL.n266 VTAIL.n265 585
R78 VTAIL.n271 VTAIL.n270 585
R79 VTAIL.n273 VTAIL.n272 585
R80 VTAIL.n262 VTAIL.n261 585
R81 VTAIL.n279 VTAIL.n278 585
R82 VTAIL.n281 VTAIL.n280 585
R83 VTAIL.n258 VTAIL.n257 585
R84 VTAIL.n287 VTAIL.n286 585
R85 VTAIL.n289 VTAIL.n288 585
R86 VTAIL.n254 VTAIL.n253 585
R87 VTAIL.n295 VTAIL.n294 585
R88 VTAIL.n297 VTAIL.n296 585
R89 VTAIL.n250 VTAIL.n249 585
R90 VTAIL.n303 VTAIL.n302 585
R91 VTAIL.n305 VTAIL.n304 585
R92 VTAIL.n246 VTAIL.n245 585
R93 VTAIL.n312 VTAIL.n311 585
R94 VTAIL.n313 VTAIL.n244 585
R95 VTAIL.n315 VTAIL.n314 585
R96 VTAIL.n26 VTAIL.n25 585
R97 VTAIL.n31 VTAIL.n30 585
R98 VTAIL.n33 VTAIL.n32 585
R99 VTAIL.n22 VTAIL.n21 585
R100 VTAIL.n39 VTAIL.n38 585
R101 VTAIL.n41 VTAIL.n40 585
R102 VTAIL.n18 VTAIL.n17 585
R103 VTAIL.n47 VTAIL.n46 585
R104 VTAIL.n49 VTAIL.n48 585
R105 VTAIL.n14 VTAIL.n13 585
R106 VTAIL.n55 VTAIL.n54 585
R107 VTAIL.n57 VTAIL.n56 585
R108 VTAIL.n10 VTAIL.n9 585
R109 VTAIL.n63 VTAIL.n62 585
R110 VTAIL.n65 VTAIL.n64 585
R111 VTAIL.n6 VTAIL.n5 585
R112 VTAIL.n72 VTAIL.n71 585
R113 VTAIL.n73 VTAIL.n4 585
R114 VTAIL.n75 VTAIL.n74 585
R115 VTAIL.n237 VTAIL.n236 585
R116 VTAIL.n235 VTAIL.n166 585
R117 VTAIL.n234 VTAIL.n233 585
R118 VTAIL.n169 VTAIL.n167 585
R119 VTAIL.n228 VTAIL.n227 585
R120 VTAIL.n226 VTAIL.n225 585
R121 VTAIL.n173 VTAIL.n172 585
R122 VTAIL.n220 VTAIL.n219 585
R123 VTAIL.n218 VTAIL.n217 585
R124 VTAIL.n177 VTAIL.n176 585
R125 VTAIL.n212 VTAIL.n211 585
R126 VTAIL.n210 VTAIL.n209 585
R127 VTAIL.n181 VTAIL.n180 585
R128 VTAIL.n204 VTAIL.n203 585
R129 VTAIL.n202 VTAIL.n201 585
R130 VTAIL.n185 VTAIL.n184 585
R131 VTAIL.n196 VTAIL.n195 585
R132 VTAIL.n194 VTAIL.n193 585
R133 VTAIL.n189 VTAIL.n188 585
R134 VTAIL.n157 VTAIL.n156 585
R135 VTAIL.n155 VTAIL.n86 585
R136 VTAIL.n154 VTAIL.n153 585
R137 VTAIL.n89 VTAIL.n87 585
R138 VTAIL.n148 VTAIL.n147 585
R139 VTAIL.n146 VTAIL.n145 585
R140 VTAIL.n93 VTAIL.n92 585
R141 VTAIL.n140 VTAIL.n139 585
R142 VTAIL.n138 VTAIL.n137 585
R143 VTAIL.n97 VTAIL.n96 585
R144 VTAIL.n132 VTAIL.n131 585
R145 VTAIL.n130 VTAIL.n129 585
R146 VTAIL.n101 VTAIL.n100 585
R147 VTAIL.n124 VTAIL.n123 585
R148 VTAIL.n122 VTAIL.n121 585
R149 VTAIL.n105 VTAIL.n104 585
R150 VTAIL.n116 VTAIL.n115 585
R151 VTAIL.n114 VTAIL.n113 585
R152 VTAIL.n109 VTAIL.n108 585
R153 VTAIL.n267 VTAIL.t1 327.466
R154 VTAIL.n27 VTAIL.t8 327.466
R155 VTAIL.n190 VTAIL.t10 327.466
R156 VTAIL.n110 VTAIL.t2 327.466
R157 VTAIL.n271 VTAIL.n265 171.744
R158 VTAIL.n272 VTAIL.n271 171.744
R159 VTAIL.n272 VTAIL.n261 171.744
R160 VTAIL.n279 VTAIL.n261 171.744
R161 VTAIL.n280 VTAIL.n279 171.744
R162 VTAIL.n280 VTAIL.n257 171.744
R163 VTAIL.n287 VTAIL.n257 171.744
R164 VTAIL.n288 VTAIL.n287 171.744
R165 VTAIL.n288 VTAIL.n253 171.744
R166 VTAIL.n295 VTAIL.n253 171.744
R167 VTAIL.n296 VTAIL.n295 171.744
R168 VTAIL.n296 VTAIL.n249 171.744
R169 VTAIL.n303 VTAIL.n249 171.744
R170 VTAIL.n304 VTAIL.n303 171.744
R171 VTAIL.n304 VTAIL.n245 171.744
R172 VTAIL.n312 VTAIL.n245 171.744
R173 VTAIL.n313 VTAIL.n312 171.744
R174 VTAIL.n314 VTAIL.n313 171.744
R175 VTAIL.n31 VTAIL.n25 171.744
R176 VTAIL.n32 VTAIL.n31 171.744
R177 VTAIL.n32 VTAIL.n21 171.744
R178 VTAIL.n39 VTAIL.n21 171.744
R179 VTAIL.n40 VTAIL.n39 171.744
R180 VTAIL.n40 VTAIL.n17 171.744
R181 VTAIL.n47 VTAIL.n17 171.744
R182 VTAIL.n48 VTAIL.n47 171.744
R183 VTAIL.n48 VTAIL.n13 171.744
R184 VTAIL.n55 VTAIL.n13 171.744
R185 VTAIL.n56 VTAIL.n55 171.744
R186 VTAIL.n56 VTAIL.n9 171.744
R187 VTAIL.n63 VTAIL.n9 171.744
R188 VTAIL.n64 VTAIL.n63 171.744
R189 VTAIL.n64 VTAIL.n5 171.744
R190 VTAIL.n72 VTAIL.n5 171.744
R191 VTAIL.n73 VTAIL.n72 171.744
R192 VTAIL.n74 VTAIL.n73 171.744
R193 VTAIL.n236 VTAIL.n235 171.744
R194 VTAIL.n235 VTAIL.n234 171.744
R195 VTAIL.n234 VTAIL.n167 171.744
R196 VTAIL.n227 VTAIL.n167 171.744
R197 VTAIL.n227 VTAIL.n226 171.744
R198 VTAIL.n226 VTAIL.n172 171.744
R199 VTAIL.n219 VTAIL.n172 171.744
R200 VTAIL.n219 VTAIL.n218 171.744
R201 VTAIL.n218 VTAIL.n176 171.744
R202 VTAIL.n211 VTAIL.n176 171.744
R203 VTAIL.n211 VTAIL.n210 171.744
R204 VTAIL.n210 VTAIL.n180 171.744
R205 VTAIL.n203 VTAIL.n180 171.744
R206 VTAIL.n203 VTAIL.n202 171.744
R207 VTAIL.n202 VTAIL.n184 171.744
R208 VTAIL.n195 VTAIL.n184 171.744
R209 VTAIL.n195 VTAIL.n194 171.744
R210 VTAIL.n194 VTAIL.n188 171.744
R211 VTAIL.n156 VTAIL.n155 171.744
R212 VTAIL.n155 VTAIL.n154 171.744
R213 VTAIL.n154 VTAIL.n87 171.744
R214 VTAIL.n147 VTAIL.n87 171.744
R215 VTAIL.n147 VTAIL.n146 171.744
R216 VTAIL.n146 VTAIL.n92 171.744
R217 VTAIL.n139 VTAIL.n92 171.744
R218 VTAIL.n139 VTAIL.n138 171.744
R219 VTAIL.n138 VTAIL.n96 171.744
R220 VTAIL.n131 VTAIL.n96 171.744
R221 VTAIL.n131 VTAIL.n130 171.744
R222 VTAIL.n130 VTAIL.n100 171.744
R223 VTAIL.n123 VTAIL.n100 171.744
R224 VTAIL.n123 VTAIL.n122 171.744
R225 VTAIL.n122 VTAIL.n104 171.744
R226 VTAIL.n115 VTAIL.n104 171.744
R227 VTAIL.n115 VTAIL.n114 171.744
R228 VTAIL.n114 VTAIL.n108 171.744
R229 VTAIL.t1 VTAIL.n265 85.8723
R230 VTAIL.t8 VTAIL.n25 85.8723
R231 VTAIL.t10 VTAIL.n188 85.8723
R232 VTAIL.t2 VTAIL.n108 85.8723
R233 VTAIL.n163 VTAIL.n162 56.9828
R234 VTAIL.n83 VTAIL.n82 56.9828
R235 VTAIL.n1 VTAIL.n0 56.9826
R236 VTAIL.n81 VTAIL.n80 56.9826
R237 VTAIL.n319 VTAIL.n318 34.5126
R238 VTAIL.n79 VTAIL.n78 34.5126
R239 VTAIL.n241 VTAIL.n240 34.5126
R240 VTAIL.n161 VTAIL.n160 34.5126
R241 VTAIL.n83 VTAIL.n81 29.8841
R242 VTAIL.n319 VTAIL.n241 27.1772
R243 VTAIL.n267 VTAIL.n266 16.3895
R244 VTAIL.n27 VTAIL.n26 16.3895
R245 VTAIL.n190 VTAIL.n189 16.3895
R246 VTAIL.n110 VTAIL.n109 16.3895
R247 VTAIL.n315 VTAIL.n244 13.1884
R248 VTAIL.n75 VTAIL.n4 13.1884
R249 VTAIL.n237 VTAIL.n166 13.1884
R250 VTAIL.n157 VTAIL.n86 13.1884
R251 VTAIL.n270 VTAIL.n269 12.8005
R252 VTAIL.n311 VTAIL.n310 12.8005
R253 VTAIL.n316 VTAIL.n242 12.8005
R254 VTAIL.n30 VTAIL.n29 12.8005
R255 VTAIL.n71 VTAIL.n70 12.8005
R256 VTAIL.n76 VTAIL.n2 12.8005
R257 VTAIL.n238 VTAIL.n164 12.8005
R258 VTAIL.n233 VTAIL.n168 12.8005
R259 VTAIL.n193 VTAIL.n192 12.8005
R260 VTAIL.n158 VTAIL.n84 12.8005
R261 VTAIL.n153 VTAIL.n88 12.8005
R262 VTAIL.n113 VTAIL.n112 12.8005
R263 VTAIL.n273 VTAIL.n264 12.0247
R264 VTAIL.n309 VTAIL.n246 12.0247
R265 VTAIL.n33 VTAIL.n24 12.0247
R266 VTAIL.n69 VTAIL.n6 12.0247
R267 VTAIL.n232 VTAIL.n169 12.0247
R268 VTAIL.n196 VTAIL.n187 12.0247
R269 VTAIL.n152 VTAIL.n89 12.0247
R270 VTAIL.n116 VTAIL.n107 12.0247
R271 VTAIL.n274 VTAIL.n262 11.249
R272 VTAIL.n306 VTAIL.n305 11.249
R273 VTAIL.n34 VTAIL.n22 11.249
R274 VTAIL.n66 VTAIL.n65 11.249
R275 VTAIL.n229 VTAIL.n228 11.249
R276 VTAIL.n197 VTAIL.n185 11.249
R277 VTAIL.n149 VTAIL.n148 11.249
R278 VTAIL.n117 VTAIL.n105 11.249
R279 VTAIL.n278 VTAIL.n277 10.4732
R280 VTAIL.n302 VTAIL.n248 10.4732
R281 VTAIL.n38 VTAIL.n37 10.4732
R282 VTAIL.n62 VTAIL.n8 10.4732
R283 VTAIL.n225 VTAIL.n171 10.4732
R284 VTAIL.n201 VTAIL.n200 10.4732
R285 VTAIL.n145 VTAIL.n91 10.4732
R286 VTAIL.n121 VTAIL.n120 10.4732
R287 VTAIL.n281 VTAIL.n260 9.69747
R288 VTAIL.n301 VTAIL.n250 9.69747
R289 VTAIL.n41 VTAIL.n20 9.69747
R290 VTAIL.n61 VTAIL.n10 9.69747
R291 VTAIL.n224 VTAIL.n173 9.69747
R292 VTAIL.n204 VTAIL.n183 9.69747
R293 VTAIL.n144 VTAIL.n93 9.69747
R294 VTAIL.n124 VTAIL.n103 9.69747
R295 VTAIL.n318 VTAIL.n317 9.45567
R296 VTAIL.n78 VTAIL.n77 9.45567
R297 VTAIL.n240 VTAIL.n239 9.45567
R298 VTAIL.n160 VTAIL.n159 9.45567
R299 VTAIL.n317 VTAIL.n316 9.3005
R300 VTAIL.n256 VTAIL.n255 9.3005
R301 VTAIL.n285 VTAIL.n284 9.3005
R302 VTAIL.n283 VTAIL.n282 9.3005
R303 VTAIL.n260 VTAIL.n259 9.3005
R304 VTAIL.n277 VTAIL.n276 9.3005
R305 VTAIL.n275 VTAIL.n274 9.3005
R306 VTAIL.n264 VTAIL.n263 9.3005
R307 VTAIL.n269 VTAIL.n268 9.3005
R308 VTAIL.n291 VTAIL.n290 9.3005
R309 VTAIL.n293 VTAIL.n292 9.3005
R310 VTAIL.n252 VTAIL.n251 9.3005
R311 VTAIL.n299 VTAIL.n298 9.3005
R312 VTAIL.n301 VTAIL.n300 9.3005
R313 VTAIL.n248 VTAIL.n247 9.3005
R314 VTAIL.n307 VTAIL.n306 9.3005
R315 VTAIL.n309 VTAIL.n308 9.3005
R316 VTAIL.n310 VTAIL.n243 9.3005
R317 VTAIL.n77 VTAIL.n76 9.3005
R318 VTAIL.n16 VTAIL.n15 9.3005
R319 VTAIL.n45 VTAIL.n44 9.3005
R320 VTAIL.n43 VTAIL.n42 9.3005
R321 VTAIL.n20 VTAIL.n19 9.3005
R322 VTAIL.n37 VTAIL.n36 9.3005
R323 VTAIL.n35 VTAIL.n34 9.3005
R324 VTAIL.n24 VTAIL.n23 9.3005
R325 VTAIL.n29 VTAIL.n28 9.3005
R326 VTAIL.n51 VTAIL.n50 9.3005
R327 VTAIL.n53 VTAIL.n52 9.3005
R328 VTAIL.n12 VTAIL.n11 9.3005
R329 VTAIL.n59 VTAIL.n58 9.3005
R330 VTAIL.n61 VTAIL.n60 9.3005
R331 VTAIL.n8 VTAIL.n7 9.3005
R332 VTAIL.n67 VTAIL.n66 9.3005
R333 VTAIL.n69 VTAIL.n68 9.3005
R334 VTAIL.n70 VTAIL.n3 9.3005
R335 VTAIL.n216 VTAIL.n215 9.3005
R336 VTAIL.n175 VTAIL.n174 9.3005
R337 VTAIL.n222 VTAIL.n221 9.3005
R338 VTAIL.n224 VTAIL.n223 9.3005
R339 VTAIL.n171 VTAIL.n170 9.3005
R340 VTAIL.n230 VTAIL.n229 9.3005
R341 VTAIL.n232 VTAIL.n231 9.3005
R342 VTAIL.n168 VTAIL.n165 9.3005
R343 VTAIL.n239 VTAIL.n238 9.3005
R344 VTAIL.n214 VTAIL.n213 9.3005
R345 VTAIL.n179 VTAIL.n178 9.3005
R346 VTAIL.n208 VTAIL.n207 9.3005
R347 VTAIL.n206 VTAIL.n205 9.3005
R348 VTAIL.n183 VTAIL.n182 9.3005
R349 VTAIL.n200 VTAIL.n199 9.3005
R350 VTAIL.n198 VTAIL.n197 9.3005
R351 VTAIL.n187 VTAIL.n186 9.3005
R352 VTAIL.n192 VTAIL.n191 9.3005
R353 VTAIL.n136 VTAIL.n135 9.3005
R354 VTAIL.n95 VTAIL.n94 9.3005
R355 VTAIL.n142 VTAIL.n141 9.3005
R356 VTAIL.n144 VTAIL.n143 9.3005
R357 VTAIL.n91 VTAIL.n90 9.3005
R358 VTAIL.n150 VTAIL.n149 9.3005
R359 VTAIL.n152 VTAIL.n151 9.3005
R360 VTAIL.n88 VTAIL.n85 9.3005
R361 VTAIL.n159 VTAIL.n158 9.3005
R362 VTAIL.n134 VTAIL.n133 9.3005
R363 VTAIL.n99 VTAIL.n98 9.3005
R364 VTAIL.n128 VTAIL.n127 9.3005
R365 VTAIL.n126 VTAIL.n125 9.3005
R366 VTAIL.n103 VTAIL.n102 9.3005
R367 VTAIL.n120 VTAIL.n119 9.3005
R368 VTAIL.n118 VTAIL.n117 9.3005
R369 VTAIL.n107 VTAIL.n106 9.3005
R370 VTAIL.n112 VTAIL.n111 9.3005
R371 VTAIL.n282 VTAIL.n258 8.92171
R372 VTAIL.n298 VTAIL.n297 8.92171
R373 VTAIL.n42 VTAIL.n18 8.92171
R374 VTAIL.n58 VTAIL.n57 8.92171
R375 VTAIL.n221 VTAIL.n220 8.92171
R376 VTAIL.n205 VTAIL.n181 8.92171
R377 VTAIL.n141 VTAIL.n140 8.92171
R378 VTAIL.n125 VTAIL.n101 8.92171
R379 VTAIL.n286 VTAIL.n285 8.14595
R380 VTAIL.n294 VTAIL.n252 8.14595
R381 VTAIL.n46 VTAIL.n45 8.14595
R382 VTAIL.n54 VTAIL.n12 8.14595
R383 VTAIL.n217 VTAIL.n175 8.14595
R384 VTAIL.n209 VTAIL.n208 8.14595
R385 VTAIL.n137 VTAIL.n95 8.14595
R386 VTAIL.n129 VTAIL.n128 8.14595
R387 VTAIL.n289 VTAIL.n256 7.3702
R388 VTAIL.n293 VTAIL.n254 7.3702
R389 VTAIL.n49 VTAIL.n16 7.3702
R390 VTAIL.n53 VTAIL.n14 7.3702
R391 VTAIL.n216 VTAIL.n177 7.3702
R392 VTAIL.n212 VTAIL.n179 7.3702
R393 VTAIL.n136 VTAIL.n97 7.3702
R394 VTAIL.n132 VTAIL.n99 7.3702
R395 VTAIL.n290 VTAIL.n289 6.59444
R396 VTAIL.n290 VTAIL.n254 6.59444
R397 VTAIL.n50 VTAIL.n49 6.59444
R398 VTAIL.n50 VTAIL.n14 6.59444
R399 VTAIL.n213 VTAIL.n177 6.59444
R400 VTAIL.n213 VTAIL.n212 6.59444
R401 VTAIL.n133 VTAIL.n97 6.59444
R402 VTAIL.n133 VTAIL.n132 6.59444
R403 VTAIL.n286 VTAIL.n256 5.81868
R404 VTAIL.n294 VTAIL.n293 5.81868
R405 VTAIL.n46 VTAIL.n16 5.81868
R406 VTAIL.n54 VTAIL.n53 5.81868
R407 VTAIL.n217 VTAIL.n216 5.81868
R408 VTAIL.n209 VTAIL.n179 5.81868
R409 VTAIL.n137 VTAIL.n136 5.81868
R410 VTAIL.n129 VTAIL.n99 5.81868
R411 VTAIL.n285 VTAIL.n258 5.04292
R412 VTAIL.n297 VTAIL.n252 5.04292
R413 VTAIL.n45 VTAIL.n18 5.04292
R414 VTAIL.n57 VTAIL.n12 5.04292
R415 VTAIL.n220 VTAIL.n175 5.04292
R416 VTAIL.n208 VTAIL.n181 5.04292
R417 VTAIL.n140 VTAIL.n95 5.04292
R418 VTAIL.n128 VTAIL.n101 5.04292
R419 VTAIL.n282 VTAIL.n281 4.26717
R420 VTAIL.n298 VTAIL.n250 4.26717
R421 VTAIL.n42 VTAIL.n41 4.26717
R422 VTAIL.n58 VTAIL.n10 4.26717
R423 VTAIL.n221 VTAIL.n173 4.26717
R424 VTAIL.n205 VTAIL.n204 4.26717
R425 VTAIL.n141 VTAIL.n93 4.26717
R426 VTAIL.n125 VTAIL.n124 4.26717
R427 VTAIL.n268 VTAIL.n267 3.70982
R428 VTAIL.n28 VTAIL.n27 3.70982
R429 VTAIL.n191 VTAIL.n190 3.70982
R430 VTAIL.n111 VTAIL.n110 3.70982
R431 VTAIL.n278 VTAIL.n260 3.49141
R432 VTAIL.n302 VTAIL.n301 3.49141
R433 VTAIL.n38 VTAIL.n20 3.49141
R434 VTAIL.n62 VTAIL.n61 3.49141
R435 VTAIL.n225 VTAIL.n224 3.49141
R436 VTAIL.n201 VTAIL.n183 3.49141
R437 VTAIL.n145 VTAIL.n144 3.49141
R438 VTAIL.n121 VTAIL.n103 3.49141
R439 VTAIL.n277 VTAIL.n262 2.71565
R440 VTAIL.n305 VTAIL.n248 2.71565
R441 VTAIL.n37 VTAIL.n22 2.71565
R442 VTAIL.n65 VTAIL.n8 2.71565
R443 VTAIL.n228 VTAIL.n171 2.71565
R444 VTAIL.n200 VTAIL.n185 2.71565
R445 VTAIL.n148 VTAIL.n91 2.71565
R446 VTAIL.n120 VTAIL.n105 2.71565
R447 VTAIL.n161 VTAIL.n83 2.7074
R448 VTAIL.n241 VTAIL.n163 2.7074
R449 VTAIL.n81 VTAIL.n79 2.7074
R450 VTAIL.n0 VTAIL.t5 2.31567
R451 VTAIL.n0 VTAIL.t4 2.31567
R452 VTAIL.n80 VTAIL.t9 2.31567
R453 VTAIL.n80 VTAIL.t11 2.31567
R454 VTAIL.n162 VTAIL.t7 2.31567
R455 VTAIL.n162 VTAIL.t6 2.31567
R456 VTAIL.n82 VTAIL.t0 2.31567
R457 VTAIL.n82 VTAIL.t3 2.31567
R458 VTAIL VTAIL.n319 1.97248
R459 VTAIL.n274 VTAIL.n273 1.93989
R460 VTAIL.n306 VTAIL.n246 1.93989
R461 VTAIL.n34 VTAIL.n33 1.93989
R462 VTAIL.n66 VTAIL.n6 1.93989
R463 VTAIL.n229 VTAIL.n169 1.93989
R464 VTAIL.n197 VTAIL.n196 1.93989
R465 VTAIL.n149 VTAIL.n89 1.93989
R466 VTAIL.n117 VTAIL.n116 1.93989
R467 VTAIL.n163 VTAIL.n161 1.82378
R468 VTAIL.n79 VTAIL.n1 1.82378
R469 VTAIL.n270 VTAIL.n264 1.16414
R470 VTAIL.n311 VTAIL.n309 1.16414
R471 VTAIL.n318 VTAIL.n242 1.16414
R472 VTAIL.n30 VTAIL.n24 1.16414
R473 VTAIL.n71 VTAIL.n69 1.16414
R474 VTAIL.n78 VTAIL.n2 1.16414
R475 VTAIL.n240 VTAIL.n164 1.16414
R476 VTAIL.n233 VTAIL.n232 1.16414
R477 VTAIL.n193 VTAIL.n187 1.16414
R478 VTAIL.n160 VTAIL.n84 1.16414
R479 VTAIL.n153 VTAIL.n152 1.16414
R480 VTAIL.n113 VTAIL.n107 1.16414
R481 VTAIL VTAIL.n1 0.735414
R482 VTAIL.n269 VTAIL.n266 0.388379
R483 VTAIL.n310 VTAIL.n244 0.388379
R484 VTAIL.n316 VTAIL.n315 0.388379
R485 VTAIL.n29 VTAIL.n26 0.388379
R486 VTAIL.n70 VTAIL.n4 0.388379
R487 VTAIL.n76 VTAIL.n75 0.388379
R488 VTAIL.n238 VTAIL.n237 0.388379
R489 VTAIL.n168 VTAIL.n166 0.388379
R490 VTAIL.n192 VTAIL.n189 0.388379
R491 VTAIL.n158 VTAIL.n157 0.388379
R492 VTAIL.n88 VTAIL.n86 0.388379
R493 VTAIL.n112 VTAIL.n109 0.388379
R494 VTAIL.n268 VTAIL.n263 0.155672
R495 VTAIL.n275 VTAIL.n263 0.155672
R496 VTAIL.n276 VTAIL.n275 0.155672
R497 VTAIL.n276 VTAIL.n259 0.155672
R498 VTAIL.n283 VTAIL.n259 0.155672
R499 VTAIL.n284 VTAIL.n283 0.155672
R500 VTAIL.n284 VTAIL.n255 0.155672
R501 VTAIL.n291 VTAIL.n255 0.155672
R502 VTAIL.n292 VTAIL.n291 0.155672
R503 VTAIL.n292 VTAIL.n251 0.155672
R504 VTAIL.n299 VTAIL.n251 0.155672
R505 VTAIL.n300 VTAIL.n299 0.155672
R506 VTAIL.n300 VTAIL.n247 0.155672
R507 VTAIL.n307 VTAIL.n247 0.155672
R508 VTAIL.n308 VTAIL.n307 0.155672
R509 VTAIL.n308 VTAIL.n243 0.155672
R510 VTAIL.n317 VTAIL.n243 0.155672
R511 VTAIL.n28 VTAIL.n23 0.155672
R512 VTAIL.n35 VTAIL.n23 0.155672
R513 VTAIL.n36 VTAIL.n35 0.155672
R514 VTAIL.n36 VTAIL.n19 0.155672
R515 VTAIL.n43 VTAIL.n19 0.155672
R516 VTAIL.n44 VTAIL.n43 0.155672
R517 VTAIL.n44 VTAIL.n15 0.155672
R518 VTAIL.n51 VTAIL.n15 0.155672
R519 VTAIL.n52 VTAIL.n51 0.155672
R520 VTAIL.n52 VTAIL.n11 0.155672
R521 VTAIL.n59 VTAIL.n11 0.155672
R522 VTAIL.n60 VTAIL.n59 0.155672
R523 VTAIL.n60 VTAIL.n7 0.155672
R524 VTAIL.n67 VTAIL.n7 0.155672
R525 VTAIL.n68 VTAIL.n67 0.155672
R526 VTAIL.n68 VTAIL.n3 0.155672
R527 VTAIL.n77 VTAIL.n3 0.155672
R528 VTAIL.n239 VTAIL.n165 0.155672
R529 VTAIL.n231 VTAIL.n165 0.155672
R530 VTAIL.n231 VTAIL.n230 0.155672
R531 VTAIL.n230 VTAIL.n170 0.155672
R532 VTAIL.n223 VTAIL.n170 0.155672
R533 VTAIL.n223 VTAIL.n222 0.155672
R534 VTAIL.n222 VTAIL.n174 0.155672
R535 VTAIL.n215 VTAIL.n174 0.155672
R536 VTAIL.n215 VTAIL.n214 0.155672
R537 VTAIL.n214 VTAIL.n178 0.155672
R538 VTAIL.n207 VTAIL.n178 0.155672
R539 VTAIL.n207 VTAIL.n206 0.155672
R540 VTAIL.n206 VTAIL.n182 0.155672
R541 VTAIL.n199 VTAIL.n182 0.155672
R542 VTAIL.n199 VTAIL.n198 0.155672
R543 VTAIL.n198 VTAIL.n186 0.155672
R544 VTAIL.n191 VTAIL.n186 0.155672
R545 VTAIL.n159 VTAIL.n85 0.155672
R546 VTAIL.n151 VTAIL.n85 0.155672
R547 VTAIL.n151 VTAIL.n150 0.155672
R548 VTAIL.n150 VTAIL.n90 0.155672
R549 VTAIL.n143 VTAIL.n90 0.155672
R550 VTAIL.n143 VTAIL.n142 0.155672
R551 VTAIL.n142 VTAIL.n94 0.155672
R552 VTAIL.n135 VTAIL.n94 0.155672
R553 VTAIL.n135 VTAIL.n134 0.155672
R554 VTAIL.n134 VTAIL.n98 0.155672
R555 VTAIL.n127 VTAIL.n98 0.155672
R556 VTAIL.n127 VTAIL.n126 0.155672
R557 VTAIL.n126 VTAIL.n102 0.155672
R558 VTAIL.n119 VTAIL.n102 0.155672
R559 VTAIL.n119 VTAIL.n118 0.155672
R560 VTAIL.n118 VTAIL.n106 0.155672
R561 VTAIL.n111 VTAIL.n106 0.155672
R562 VDD1.n72 VDD1.n0 756.745
R563 VDD1.n149 VDD1.n77 756.745
R564 VDD1.n73 VDD1.n72 585
R565 VDD1.n71 VDD1.n2 585
R566 VDD1.n70 VDD1.n69 585
R567 VDD1.n5 VDD1.n3 585
R568 VDD1.n64 VDD1.n63 585
R569 VDD1.n62 VDD1.n61 585
R570 VDD1.n9 VDD1.n8 585
R571 VDD1.n56 VDD1.n55 585
R572 VDD1.n54 VDD1.n53 585
R573 VDD1.n13 VDD1.n12 585
R574 VDD1.n48 VDD1.n47 585
R575 VDD1.n46 VDD1.n45 585
R576 VDD1.n17 VDD1.n16 585
R577 VDD1.n40 VDD1.n39 585
R578 VDD1.n38 VDD1.n37 585
R579 VDD1.n21 VDD1.n20 585
R580 VDD1.n32 VDD1.n31 585
R581 VDD1.n30 VDD1.n29 585
R582 VDD1.n25 VDD1.n24 585
R583 VDD1.n101 VDD1.n100 585
R584 VDD1.n106 VDD1.n105 585
R585 VDD1.n108 VDD1.n107 585
R586 VDD1.n97 VDD1.n96 585
R587 VDD1.n114 VDD1.n113 585
R588 VDD1.n116 VDD1.n115 585
R589 VDD1.n93 VDD1.n92 585
R590 VDD1.n122 VDD1.n121 585
R591 VDD1.n124 VDD1.n123 585
R592 VDD1.n89 VDD1.n88 585
R593 VDD1.n130 VDD1.n129 585
R594 VDD1.n132 VDD1.n131 585
R595 VDD1.n85 VDD1.n84 585
R596 VDD1.n138 VDD1.n137 585
R597 VDD1.n140 VDD1.n139 585
R598 VDD1.n81 VDD1.n80 585
R599 VDD1.n147 VDD1.n146 585
R600 VDD1.n148 VDD1.n79 585
R601 VDD1.n150 VDD1.n149 585
R602 VDD1.n26 VDD1.t1 327.466
R603 VDD1.n102 VDD1.t0 327.466
R604 VDD1.n72 VDD1.n71 171.744
R605 VDD1.n71 VDD1.n70 171.744
R606 VDD1.n70 VDD1.n3 171.744
R607 VDD1.n63 VDD1.n3 171.744
R608 VDD1.n63 VDD1.n62 171.744
R609 VDD1.n62 VDD1.n8 171.744
R610 VDD1.n55 VDD1.n8 171.744
R611 VDD1.n55 VDD1.n54 171.744
R612 VDD1.n54 VDD1.n12 171.744
R613 VDD1.n47 VDD1.n12 171.744
R614 VDD1.n47 VDD1.n46 171.744
R615 VDD1.n46 VDD1.n16 171.744
R616 VDD1.n39 VDD1.n16 171.744
R617 VDD1.n39 VDD1.n38 171.744
R618 VDD1.n38 VDD1.n20 171.744
R619 VDD1.n31 VDD1.n20 171.744
R620 VDD1.n31 VDD1.n30 171.744
R621 VDD1.n30 VDD1.n24 171.744
R622 VDD1.n106 VDD1.n100 171.744
R623 VDD1.n107 VDD1.n106 171.744
R624 VDD1.n107 VDD1.n96 171.744
R625 VDD1.n114 VDD1.n96 171.744
R626 VDD1.n115 VDD1.n114 171.744
R627 VDD1.n115 VDD1.n92 171.744
R628 VDD1.n122 VDD1.n92 171.744
R629 VDD1.n123 VDD1.n122 171.744
R630 VDD1.n123 VDD1.n88 171.744
R631 VDD1.n130 VDD1.n88 171.744
R632 VDD1.n131 VDD1.n130 171.744
R633 VDD1.n131 VDD1.n84 171.744
R634 VDD1.n138 VDD1.n84 171.744
R635 VDD1.n139 VDD1.n138 171.744
R636 VDD1.n139 VDD1.n80 171.744
R637 VDD1.n147 VDD1.n80 171.744
R638 VDD1.n148 VDD1.n147 171.744
R639 VDD1.n149 VDD1.n148 171.744
R640 VDD1.t1 VDD1.n24 85.8723
R641 VDD1.t0 VDD1.n100 85.8723
R642 VDD1.n155 VDD1.n154 74.2828
R643 VDD1.n157 VDD1.n156 73.6614
R644 VDD1 VDD1.n76 53.2798
R645 VDD1.n155 VDD1.n153 53.1662
R646 VDD1.n157 VDD1.n155 46.5526
R647 VDD1.n26 VDD1.n25 16.3895
R648 VDD1.n102 VDD1.n101 16.3895
R649 VDD1.n73 VDD1.n2 13.1884
R650 VDD1.n150 VDD1.n79 13.1884
R651 VDD1.n74 VDD1.n0 12.8005
R652 VDD1.n69 VDD1.n4 12.8005
R653 VDD1.n29 VDD1.n28 12.8005
R654 VDD1.n105 VDD1.n104 12.8005
R655 VDD1.n146 VDD1.n145 12.8005
R656 VDD1.n151 VDD1.n77 12.8005
R657 VDD1.n68 VDD1.n5 12.0247
R658 VDD1.n32 VDD1.n23 12.0247
R659 VDD1.n108 VDD1.n99 12.0247
R660 VDD1.n144 VDD1.n81 12.0247
R661 VDD1.n65 VDD1.n64 11.249
R662 VDD1.n33 VDD1.n21 11.249
R663 VDD1.n109 VDD1.n97 11.249
R664 VDD1.n141 VDD1.n140 11.249
R665 VDD1.n61 VDD1.n7 10.4732
R666 VDD1.n37 VDD1.n36 10.4732
R667 VDD1.n113 VDD1.n112 10.4732
R668 VDD1.n137 VDD1.n83 10.4732
R669 VDD1.n60 VDD1.n9 9.69747
R670 VDD1.n40 VDD1.n19 9.69747
R671 VDD1.n116 VDD1.n95 9.69747
R672 VDD1.n136 VDD1.n85 9.69747
R673 VDD1.n76 VDD1.n75 9.45567
R674 VDD1.n153 VDD1.n152 9.45567
R675 VDD1.n52 VDD1.n51 9.3005
R676 VDD1.n11 VDD1.n10 9.3005
R677 VDD1.n58 VDD1.n57 9.3005
R678 VDD1.n60 VDD1.n59 9.3005
R679 VDD1.n7 VDD1.n6 9.3005
R680 VDD1.n66 VDD1.n65 9.3005
R681 VDD1.n68 VDD1.n67 9.3005
R682 VDD1.n4 VDD1.n1 9.3005
R683 VDD1.n75 VDD1.n74 9.3005
R684 VDD1.n50 VDD1.n49 9.3005
R685 VDD1.n15 VDD1.n14 9.3005
R686 VDD1.n44 VDD1.n43 9.3005
R687 VDD1.n42 VDD1.n41 9.3005
R688 VDD1.n19 VDD1.n18 9.3005
R689 VDD1.n36 VDD1.n35 9.3005
R690 VDD1.n34 VDD1.n33 9.3005
R691 VDD1.n23 VDD1.n22 9.3005
R692 VDD1.n28 VDD1.n27 9.3005
R693 VDD1.n152 VDD1.n151 9.3005
R694 VDD1.n91 VDD1.n90 9.3005
R695 VDD1.n120 VDD1.n119 9.3005
R696 VDD1.n118 VDD1.n117 9.3005
R697 VDD1.n95 VDD1.n94 9.3005
R698 VDD1.n112 VDD1.n111 9.3005
R699 VDD1.n110 VDD1.n109 9.3005
R700 VDD1.n99 VDD1.n98 9.3005
R701 VDD1.n104 VDD1.n103 9.3005
R702 VDD1.n126 VDD1.n125 9.3005
R703 VDD1.n128 VDD1.n127 9.3005
R704 VDD1.n87 VDD1.n86 9.3005
R705 VDD1.n134 VDD1.n133 9.3005
R706 VDD1.n136 VDD1.n135 9.3005
R707 VDD1.n83 VDD1.n82 9.3005
R708 VDD1.n142 VDD1.n141 9.3005
R709 VDD1.n144 VDD1.n143 9.3005
R710 VDD1.n145 VDD1.n78 9.3005
R711 VDD1.n57 VDD1.n56 8.92171
R712 VDD1.n41 VDD1.n17 8.92171
R713 VDD1.n117 VDD1.n93 8.92171
R714 VDD1.n133 VDD1.n132 8.92171
R715 VDD1.n53 VDD1.n11 8.14595
R716 VDD1.n45 VDD1.n44 8.14595
R717 VDD1.n121 VDD1.n120 8.14595
R718 VDD1.n129 VDD1.n87 8.14595
R719 VDD1.n52 VDD1.n13 7.3702
R720 VDD1.n48 VDD1.n15 7.3702
R721 VDD1.n124 VDD1.n91 7.3702
R722 VDD1.n128 VDD1.n89 7.3702
R723 VDD1.n49 VDD1.n13 6.59444
R724 VDD1.n49 VDD1.n48 6.59444
R725 VDD1.n125 VDD1.n124 6.59444
R726 VDD1.n125 VDD1.n89 6.59444
R727 VDD1.n53 VDD1.n52 5.81868
R728 VDD1.n45 VDD1.n15 5.81868
R729 VDD1.n121 VDD1.n91 5.81868
R730 VDD1.n129 VDD1.n128 5.81868
R731 VDD1.n56 VDD1.n11 5.04292
R732 VDD1.n44 VDD1.n17 5.04292
R733 VDD1.n120 VDD1.n93 5.04292
R734 VDD1.n132 VDD1.n87 5.04292
R735 VDD1.n57 VDD1.n9 4.26717
R736 VDD1.n41 VDD1.n40 4.26717
R737 VDD1.n117 VDD1.n116 4.26717
R738 VDD1.n133 VDD1.n85 4.26717
R739 VDD1.n27 VDD1.n26 3.70982
R740 VDD1.n103 VDD1.n102 3.70982
R741 VDD1.n61 VDD1.n60 3.49141
R742 VDD1.n37 VDD1.n19 3.49141
R743 VDD1.n113 VDD1.n95 3.49141
R744 VDD1.n137 VDD1.n136 3.49141
R745 VDD1.n64 VDD1.n7 2.71565
R746 VDD1.n36 VDD1.n21 2.71565
R747 VDD1.n112 VDD1.n97 2.71565
R748 VDD1.n140 VDD1.n83 2.71565
R749 VDD1.n156 VDD1.t2 2.31567
R750 VDD1.n156 VDD1.t5 2.31567
R751 VDD1.n154 VDD1.t3 2.31567
R752 VDD1.n154 VDD1.t4 2.31567
R753 VDD1.n65 VDD1.n5 1.93989
R754 VDD1.n33 VDD1.n32 1.93989
R755 VDD1.n109 VDD1.n108 1.93989
R756 VDD1.n141 VDD1.n81 1.93989
R757 VDD1.n76 VDD1.n0 1.16414
R758 VDD1.n69 VDD1.n68 1.16414
R759 VDD1.n29 VDD1.n23 1.16414
R760 VDD1.n105 VDD1.n99 1.16414
R761 VDD1.n146 VDD1.n144 1.16414
R762 VDD1.n153 VDD1.n77 1.16414
R763 VDD1 VDD1.n157 0.619035
R764 VDD1.n74 VDD1.n73 0.388379
R765 VDD1.n4 VDD1.n2 0.388379
R766 VDD1.n28 VDD1.n25 0.388379
R767 VDD1.n104 VDD1.n101 0.388379
R768 VDD1.n145 VDD1.n79 0.388379
R769 VDD1.n151 VDD1.n150 0.388379
R770 VDD1.n75 VDD1.n1 0.155672
R771 VDD1.n67 VDD1.n1 0.155672
R772 VDD1.n67 VDD1.n66 0.155672
R773 VDD1.n66 VDD1.n6 0.155672
R774 VDD1.n59 VDD1.n6 0.155672
R775 VDD1.n59 VDD1.n58 0.155672
R776 VDD1.n58 VDD1.n10 0.155672
R777 VDD1.n51 VDD1.n10 0.155672
R778 VDD1.n51 VDD1.n50 0.155672
R779 VDD1.n50 VDD1.n14 0.155672
R780 VDD1.n43 VDD1.n14 0.155672
R781 VDD1.n43 VDD1.n42 0.155672
R782 VDD1.n42 VDD1.n18 0.155672
R783 VDD1.n35 VDD1.n18 0.155672
R784 VDD1.n35 VDD1.n34 0.155672
R785 VDD1.n34 VDD1.n22 0.155672
R786 VDD1.n27 VDD1.n22 0.155672
R787 VDD1.n103 VDD1.n98 0.155672
R788 VDD1.n110 VDD1.n98 0.155672
R789 VDD1.n111 VDD1.n110 0.155672
R790 VDD1.n111 VDD1.n94 0.155672
R791 VDD1.n118 VDD1.n94 0.155672
R792 VDD1.n119 VDD1.n118 0.155672
R793 VDD1.n119 VDD1.n90 0.155672
R794 VDD1.n126 VDD1.n90 0.155672
R795 VDD1.n127 VDD1.n126 0.155672
R796 VDD1.n127 VDD1.n86 0.155672
R797 VDD1.n134 VDD1.n86 0.155672
R798 VDD1.n135 VDD1.n134 0.155672
R799 VDD1.n135 VDD1.n82 0.155672
R800 VDD1.n142 VDD1.n82 0.155672
R801 VDD1.n143 VDD1.n142 0.155672
R802 VDD1.n143 VDD1.n78 0.155672
R803 VDD1.n152 VDD1.n78 0.155672
R804 VN.n29 VN.n16 161.3
R805 VN.n28 VN.n27 161.3
R806 VN.n26 VN.n17 161.3
R807 VN.n25 VN.n24 161.3
R808 VN.n23 VN.n18 161.3
R809 VN.n22 VN.n21 161.3
R810 VN.n13 VN.n0 161.3
R811 VN.n12 VN.n11 161.3
R812 VN.n10 VN.n1 161.3
R813 VN.n9 VN.n8 161.3
R814 VN.n7 VN.n2 161.3
R815 VN.n6 VN.n5 161.3
R816 VN.n4 VN.t1 155.148
R817 VN.n20 VN.t2 155.148
R818 VN.n3 VN.t4 120.415
R819 VN.n14 VN.t0 120.415
R820 VN.n19 VN.t3 120.415
R821 VN.n30 VN.t5 120.415
R822 VN.n15 VN.n14 104.022
R823 VN.n31 VN.n30 104.022
R824 VN VN.n31 51.3467
R825 VN.n20 VN.n19 49.0208
R826 VN.n4 VN.n3 49.0208
R827 VN.n8 VN.n1 47.3584
R828 VN.n24 VN.n17 47.3584
R829 VN.n8 VN.n7 33.7956
R830 VN.n24 VN.n23 33.7956
R831 VN.n6 VN.n3 24.5923
R832 VN.n7 VN.n6 24.5923
R833 VN.n12 VN.n1 24.5923
R834 VN.n13 VN.n12 24.5923
R835 VN.n23 VN.n22 24.5923
R836 VN.n22 VN.n19 24.5923
R837 VN.n29 VN.n28 24.5923
R838 VN.n28 VN.n17 24.5923
R839 VN.n14 VN.n13 6.88621
R840 VN.n30 VN.n29 6.88621
R841 VN.n21 VN.n20 4.88317
R842 VN.n5 VN.n4 4.88317
R843 VN.n31 VN.n16 0.278335
R844 VN.n15 VN.n0 0.278335
R845 VN.n27 VN.n16 0.189894
R846 VN.n27 VN.n26 0.189894
R847 VN.n26 VN.n25 0.189894
R848 VN.n25 VN.n18 0.189894
R849 VN.n21 VN.n18 0.189894
R850 VN.n5 VN.n2 0.189894
R851 VN.n9 VN.n2 0.189894
R852 VN.n10 VN.n9 0.189894
R853 VN.n11 VN.n10 0.189894
R854 VN.n11 VN.n0 0.189894
R855 VN VN.n15 0.153485
R856 VDD2.n151 VDD2.n79 756.745
R857 VDD2.n72 VDD2.n0 756.745
R858 VDD2.n152 VDD2.n151 585
R859 VDD2.n150 VDD2.n81 585
R860 VDD2.n149 VDD2.n148 585
R861 VDD2.n84 VDD2.n82 585
R862 VDD2.n143 VDD2.n142 585
R863 VDD2.n141 VDD2.n140 585
R864 VDD2.n88 VDD2.n87 585
R865 VDD2.n135 VDD2.n134 585
R866 VDD2.n133 VDD2.n132 585
R867 VDD2.n92 VDD2.n91 585
R868 VDD2.n127 VDD2.n126 585
R869 VDD2.n125 VDD2.n124 585
R870 VDD2.n96 VDD2.n95 585
R871 VDD2.n119 VDD2.n118 585
R872 VDD2.n117 VDD2.n116 585
R873 VDD2.n100 VDD2.n99 585
R874 VDD2.n111 VDD2.n110 585
R875 VDD2.n109 VDD2.n108 585
R876 VDD2.n104 VDD2.n103 585
R877 VDD2.n24 VDD2.n23 585
R878 VDD2.n29 VDD2.n28 585
R879 VDD2.n31 VDD2.n30 585
R880 VDD2.n20 VDD2.n19 585
R881 VDD2.n37 VDD2.n36 585
R882 VDD2.n39 VDD2.n38 585
R883 VDD2.n16 VDD2.n15 585
R884 VDD2.n45 VDD2.n44 585
R885 VDD2.n47 VDD2.n46 585
R886 VDD2.n12 VDD2.n11 585
R887 VDD2.n53 VDD2.n52 585
R888 VDD2.n55 VDD2.n54 585
R889 VDD2.n8 VDD2.n7 585
R890 VDD2.n61 VDD2.n60 585
R891 VDD2.n63 VDD2.n62 585
R892 VDD2.n4 VDD2.n3 585
R893 VDD2.n70 VDD2.n69 585
R894 VDD2.n71 VDD2.n2 585
R895 VDD2.n73 VDD2.n72 585
R896 VDD2.n105 VDD2.t0 327.466
R897 VDD2.n25 VDD2.t4 327.466
R898 VDD2.n151 VDD2.n150 171.744
R899 VDD2.n150 VDD2.n149 171.744
R900 VDD2.n149 VDD2.n82 171.744
R901 VDD2.n142 VDD2.n82 171.744
R902 VDD2.n142 VDD2.n141 171.744
R903 VDD2.n141 VDD2.n87 171.744
R904 VDD2.n134 VDD2.n87 171.744
R905 VDD2.n134 VDD2.n133 171.744
R906 VDD2.n133 VDD2.n91 171.744
R907 VDD2.n126 VDD2.n91 171.744
R908 VDD2.n126 VDD2.n125 171.744
R909 VDD2.n125 VDD2.n95 171.744
R910 VDD2.n118 VDD2.n95 171.744
R911 VDD2.n118 VDD2.n117 171.744
R912 VDD2.n117 VDD2.n99 171.744
R913 VDD2.n110 VDD2.n99 171.744
R914 VDD2.n110 VDD2.n109 171.744
R915 VDD2.n109 VDD2.n103 171.744
R916 VDD2.n29 VDD2.n23 171.744
R917 VDD2.n30 VDD2.n29 171.744
R918 VDD2.n30 VDD2.n19 171.744
R919 VDD2.n37 VDD2.n19 171.744
R920 VDD2.n38 VDD2.n37 171.744
R921 VDD2.n38 VDD2.n15 171.744
R922 VDD2.n45 VDD2.n15 171.744
R923 VDD2.n46 VDD2.n45 171.744
R924 VDD2.n46 VDD2.n11 171.744
R925 VDD2.n53 VDD2.n11 171.744
R926 VDD2.n54 VDD2.n53 171.744
R927 VDD2.n54 VDD2.n7 171.744
R928 VDD2.n61 VDD2.n7 171.744
R929 VDD2.n62 VDD2.n61 171.744
R930 VDD2.n62 VDD2.n3 171.744
R931 VDD2.n70 VDD2.n3 171.744
R932 VDD2.n71 VDD2.n70 171.744
R933 VDD2.n72 VDD2.n71 171.744
R934 VDD2.t0 VDD2.n103 85.8723
R935 VDD2.t4 VDD2.n23 85.8723
R936 VDD2.n78 VDD2.n77 74.2828
R937 VDD2 VDD2.n157 74.2799
R938 VDD2.n78 VDD2.n76 53.1662
R939 VDD2.n156 VDD2.n155 51.1914
R940 VDD2.n156 VDD2.n78 44.6162
R941 VDD2.n105 VDD2.n104 16.3895
R942 VDD2.n25 VDD2.n24 16.3895
R943 VDD2.n152 VDD2.n81 13.1884
R944 VDD2.n73 VDD2.n2 13.1884
R945 VDD2.n153 VDD2.n79 12.8005
R946 VDD2.n148 VDD2.n83 12.8005
R947 VDD2.n108 VDD2.n107 12.8005
R948 VDD2.n28 VDD2.n27 12.8005
R949 VDD2.n69 VDD2.n68 12.8005
R950 VDD2.n74 VDD2.n0 12.8005
R951 VDD2.n147 VDD2.n84 12.0247
R952 VDD2.n111 VDD2.n102 12.0247
R953 VDD2.n31 VDD2.n22 12.0247
R954 VDD2.n67 VDD2.n4 12.0247
R955 VDD2.n144 VDD2.n143 11.249
R956 VDD2.n112 VDD2.n100 11.249
R957 VDD2.n32 VDD2.n20 11.249
R958 VDD2.n64 VDD2.n63 11.249
R959 VDD2.n140 VDD2.n86 10.4732
R960 VDD2.n116 VDD2.n115 10.4732
R961 VDD2.n36 VDD2.n35 10.4732
R962 VDD2.n60 VDD2.n6 10.4732
R963 VDD2.n139 VDD2.n88 9.69747
R964 VDD2.n119 VDD2.n98 9.69747
R965 VDD2.n39 VDD2.n18 9.69747
R966 VDD2.n59 VDD2.n8 9.69747
R967 VDD2.n155 VDD2.n154 9.45567
R968 VDD2.n76 VDD2.n75 9.45567
R969 VDD2.n131 VDD2.n130 9.3005
R970 VDD2.n90 VDD2.n89 9.3005
R971 VDD2.n137 VDD2.n136 9.3005
R972 VDD2.n139 VDD2.n138 9.3005
R973 VDD2.n86 VDD2.n85 9.3005
R974 VDD2.n145 VDD2.n144 9.3005
R975 VDD2.n147 VDD2.n146 9.3005
R976 VDD2.n83 VDD2.n80 9.3005
R977 VDD2.n154 VDD2.n153 9.3005
R978 VDD2.n129 VDD2.n128 9.3005
R979 VDD2.n94 VDD2.n93 9.3005
R980 VDD2.n123 VDD2.n122 9.3005
R981 VDD2.n121 VDD2.n120 9.3005
R982 VDD2.n98 VDD2.n97 9.3005
R983 VDD2.n115 VDD2.n114 9.3005
R984 VDD2.n113 VDD2.n112 9.3005
R985 VDD2.n102 VDD2.n101 9.3005
R986 VDD2.n107 VDD2.n106 9.3005
R987 VDD2.n75 VDD2.n74 9.3005
R988 VDD2.n14 VDD2.n13 9.3005
R989 VDD2.n43 VDD2.n42 9.3005
R990 VDD2.n41 VDD2.n40 9.3005
R991 VDD2.n18 VDD2.n17 9.3005
R992 VDD2.n35 VDD2.n34 9.3005
R993 VDD2.n33 VDD2.n32 9.3005
R994 VDD2.n22 VDD2.n21 9.3005
R995 VDD2.n27 VDD2.n26 9.3005
R996 VDD2.n49 VDD2.n48 9.3005
R997 VDD2.n51 VDD2.n50 9.3005
R998 VDD2.n10 VDD2.n9 9.3005
R999 VDD2.n57 VDD2.n56 9.3005
R1000 VDD2.n59 VDD2.n58 9.3005
R1001 VDD2.n6 VDD2.n5 9.3005
R1002 VDD2.n65 VDD2.n64 9.3005
R1003 VDD2.n67 VDD2.n66 9.3005
R1004 VDD2.n68 VDD2.n1 9.3005
R1005 VDD2.n136 VDD2.n135 8.92171
R1006 VDD2.n120 VDD2.n96 8.92171
R1007 VDD2.n40 VDD2.n16 8.92171
R1008 VDD2.n56 VDD2.n55 8.92171
R1009 VDD2.n132 VDD2.n90 8.14595
R1010 VDD2.n124 VDD2.n123 8.14595
R1011 VDD2.n44 VDD2.n43 8.14595
R1012 VDD2.n52 VDD2.n10 8.14595
R1013 VDD2.n131 VDD2.n92 7.3702
R1014 VDD2.n127 VDD2.n94 7.3702
R1015 VDD2.n47 VDD2.n14 7.3702
R1016 VDD2.n51 VDD2.n12 7.3702
R1017 VDD2.n128 VDD2.n92 6.59444
R1018 VDD2.n128 VDD2.n127 6.59444
R1019 VDD2.n48 VDD2.n47 6.59444
R1020 VDD2.n48 VDD2.n12 6.59444
R1021 VDD2.n132 VDD2.n131 5.81868
R1022 VDD2.n124 VDD2.n94 5.81868
R1023 VDD2.n44 VDD2.n14 5.81868
R1024 VDD2.n52 VDD2.n51 5.81868
R1025 VDD2.n135 VDD2.n90 5.04292
R1026 VDD2.n123 VDD2.n96 5.04292
R1027 VDD2.n43 VDD2.n16 5.04292
R1028 VDD2.n55 VDD2.n10 5.04292
R1029 VDD2.n136 VDD2.n88 4.26717
R1030 VDD2.n120 VDD2.n119 4.26717
R1031 VDD2.n40 VDD2.n39 4.26717
R1032 VDD2.n56 VDD2.n8 4.26717
R1033 VDD2.n106 VDD2.n105 3.70982
R1034 VDD2.n26 VDD2.n25 3.70982
R1035 VDD2.n140 VDD2.n139 3.49141
R1036 VDD2.n116 VDD2.n98 3.49141
R1037 VDD2.n36 VDD2.n18 3.49141
R1038 VDD2.n60 VDD2.n59 3.49141
R1039 VDD2.n143 VDD2.n86 2.71565
R1040 VDD2.n115 VDD2.n100 2.71565
R1041 VDD2.n35 VDD2.n20 2.71565
R1042 VDD2.n63 VDD2.n6 2.71565
R1043 VDD2.n157 VDD2.t2 2.31567
R1044 VDD2.n157 VDD2.t3 2.31567
R1045 VDD2.n77 VDD2.t1 2.31567
R1046 VDD2.n77 VDD2.t5 2.31567
R1047 VDD2 VDD2.n156 2.08886
R1048 VDD2.n144 VDD2.n84 1.93989
R1049 VDD2.n112 VDD2.n111 1.93989
R1050 VDD2.n32 VDD2.n31 1.93989
R1051 VDD2.n64 VDD2.n4 1.93989
R1052 VDD2.n155 VDD2.n79 1.16414
R1053 VDD2.n148 VDD2.n147 1.16414
R1054 VDD2.n108 VDD2.n102 1.16414
R1055 VDD2.n28 VDD2.n22 1.16414
R1056 VDD2.n69 VDD2.n67 1.16414
R1057 VDD2.n76 VDD2.n0 1.16414
R1058 VDD2.n153 VDD2.n152 0.388379
R1059 VDD2.n83 VDD2.n81 0.388379
R1060 VDD2.n107 VDD2.n104 0.388379
R1061 VDD2.n27 VDD2.n24 0.388379
R1062 VDD2.n68 VDD2.n2 0.388379
R1063 VDD2.n74 VDD2.n73 0.388379
R1064 VDD2.n154 VDD2.n80 0.155672
R1065 VDD2.n146 VDD2.n80 0.155672
R1066 VDD2.n146 VDD2.n145 0.155672
R1067 VDD2.n145 VDD2.n85 0.155672
R1068 VDD2.n138 VDD2.n85 0.155672
R1069 VDD2.n138 VDD2.n137 0.155672
R1070 VDD2.n137 VDD2.n89 0.155672
R1071 VDD2.n130 VDD2.n89 0.155672
R1072 VDD2.n130 VDD2.n129 0.155672
R1073 VDD2.n129 VDD2.n93 0.155672
R1074 VDD2.n122 VDD2.n93 0.155672
R1075 VDD2.n122 VDD2.n121 0.155672
R1076 VDD2.n121 VDD2.n97 0.155672
R1077 VDD2.n114 VDD2.n97 0.155672
R1078 VDD2.n114 VDD2.n113 0.155672
R1079 VDD2.n113 VDD2.n101 0.155672
R1080 VDD2.n106 VDD2.n101 0.155672
R1081 VDD2.n26 VDD2.n21 0.155672
R1082 VDD2.n33 VDD2.n21 0.155672
R1083 VDD2.n34 VDD2.n33 0.155672
R1084 VDD2.n34 VDD2.n17 0.155672
R1085 VDD2.n41 VDD2.n17 0.155672
R1086 VDD2.n42 VDD2.n41 0.155672
R1087 VDD2.n42 VDD2.n13 0.155672
R1088 VDD2.n49 VDD2.n13 0.155672
R1089 VDD2.n50 VDD2.n49 0.155672
R1090 VDD2.n50 VDD2.n9 0.155672
R1091 VDD2.n57 VDD2.n9 0.155672
R1092 VDD2.n58 VDD2.n57 0.155672
R1093 VDD2.n58 VDD2.n5 0.155672
R1094 VDD2.n65 VDD2.n5 0.155672
R1095 VDD2.n66 VDD2.n65 0.155672
R1096 VDD2.n66 VDD2.n1 0.155672
R1097 VDD2.n75 VDD2.n1 0.155672
R1098 B.n569 B.n568 585
R1099 B.n570 B.n81 585
R1100 B.n572 B.n571 585
R1101 B.n573 B.n80 585
R1102 B.n575 B.n574 585
R1103 B.n576 B.n79 585
R1104 B.n578 B.n577 585
R1105 B.n579 B.n78 585
R1106 B.n581 B.n580 585
R1107 B.n582 B.n77 585
R1108 B.n584 B.n583 585
R1109 B.n585 B.n76 585
R1110 B.n587 B.n586 585
R1111 B.n588 B.n75 585
R1112 B.n590 B.n589 585
R1113 B.n591 B.n74 585
R1114 B.n593 B.n592 585
R1115 B.n594 B.n73 585
R1116 B.n596 B.n595 585
R1117 B.n597 B.n72 585
R1118 B.n599 B.n598 585
R1119 B.n600 B.n71 585
R1120 B.n602 B.n601 585
R1121 B.n603 B.n70 585
R1122 B.n605 B.n604 585
R1123 B.n606 B.n69 585
R1124 B.n608 B.n607 585
R1125 B.n609 B.n68 585
R1126 B.n611 B.n610 585
R1127 B.n612 B.n67 585
R1128 B.n614 B.n613 585
R1129 B.n615 B.n66 585
R1130 B.n617 B.n616 585
R1131 B.n618 B.n65 585
R1132 B.n620 B.n619 585
R1133 B.n621 B.n64 585
R1134 B.n623 B.n622 585
R1135 B.n624 B.n63 585
R1136 B.n626 B.n625 585
R1137 B.n627 B.n62 585
R1138 B.n629 B.n628 585
R1139 B.n630 B.n61 585
R1140 B.n632 B.n631 585
R1141 B.n633 B.n60 585
R1142 B.n635 B.n634 585
R1143 B.n636 B.n59 585
R1144 B.n638 B.n637 585
R1145 B.n639 B.n56 585
R1146 B.n642 B.n641 585
R1147 B.n643 B.n55 585
R1148 B.n645 B.n644 585
R1149 B.n646 B.n54 585
R1150 B.n648 B.n647 585
R1151 B.n649 B.n53 585
R1152 B.n651 B.n650 585
R1153 B.n652 B.n49 585
R1154 B.n654 B.n653 585
R1155 B.n655 B.n48 585
R1156 B.n657 B.n656 585
R1157 B.n658 B.n47 585
R1158 B.n660 B.n659 585
R1159 B.n661 B.n46 585
R1160 B.n663 B.n662 585
R1161 B.n664 B.n45 585
R1162 B.n666 B.n665 585
R1163 B.n667 B.n44 585
R1164 B.n669 B.n668 585
R1165 B.n670 B.n43 585
R1166 B.n672 B.n671 585
R1167 B.n673 B.n42 585
R1168 B.n675 B.n674 585
R1169 B.n676 B.n41 585
R1170 B.n678 B.n677 585
R1171 B.n679 B.n40 585
R1172 B.n681 B.n680 585
R1173 B.n682 B.n39 585
R1174 B.n684 B.n683 585
R1175 B.n685 B.n38 585
R1176 B.n687 B.n686 585
R1177 B.n688 B.n37 585
R1178 B.n690 B.n689 585
R1179 B.n691 B.n36 585
R1180 B.n693 B.n692 585
R1181 B.n694 B.n35 585
R1182 B.n696 B.n695 585
R1183 B.n697 B.n34 585
R1184 B.n699 B.n698 585
R1185 B.n700 B.n33 585
R1186 B.n702 B.n701 585
R1187 B.n703 B.n32 585
R1188 B.n705 B.n704 585
R1189 B.n706 B.n31 585
R1190 B.n708 B.n707 585
R1191 B.n709 B.n30 585
R1192 B.n711 B.n710 585
R1193 B.n712 B.n29 585
R1194 B.n714 B.n713 585
R1195 B.n715 B.n28 585
R1196 B.n717 B.n716 585
R1197 B.n718 B.n27 585
R1198 B.n720 B.n719 585
R1199 B.n721 B.n26 585
R1200 B.n723 B.n722 585
R1201 B.n724 B.n25 585
R1202 B.n726 B.n725 585
R1203 B.n567 B.n82 585
R1204 B.n566 B.n565 585
R1205 B.n564 B.n83 585
R1206 B.n563 B.n562 585
R1207 B.n561 B.n84 585
R1208 B.n560 B.n559 585
R1209 B.n558 B.n85 585
R1210 B.n557 B.n556 585
R1211 B.n555 B.n86 585
R1212 B.n554 B.n553 585
R1213 B.n552 B.n87 585
R1214 B.n551 B.n550 585
R1215 B.n549 B.n88 585
R1216 B.n548 B.n547 585
R1217 B.n546 B.n89 585
R1218 B.n545 B.n544 585
R1219 B.n543 B.n90 585
R1220 B.n542 B.n541 585
R1221 B.n540 B.n91 585
R1222 B.n539 B.n538 585
R1223 B.n537 B.n92 585
R1224 B.n536 B.n535 585
R1225 B.n534 B.n93 585
R1226 B.n533 B.n532 585
R1227 B.n531 B.n94 585
R1228 B.n530 B.n529 585
R1229 B.n528 B.n95 585
R1230 B.n527 B.n526 585
R1231 B.n525 B.n96 585
R1232 B.n524 B.n523 585
R1233 B.n522 B.n97 585
R1234 B.n521 B.n520 585
R1235 B.n519 B.n98 585
R1236 B.n518 B.n517 585
R1237 B.n516 B.n99 585
R1238 B.n515 B.n514 585
R1239 B.n513 B.n100 585
R1240 B.n512 B.n511 585
R1241 B.n510 B.n101 585
R1242 B.n509 B.n508 585
R1243 B.n507 B.n102 585
R1244 B.n506 B.n505 585
R1245 B.n504 B.n103 585
R1246 B.n503 B.n502 585
R1247 B.n501 B.n104 585
R1248 B.n500 B.n499 585
R1249 B.n498 B.n105 585
R1250 B.n497 B.n496 585
R1251 B.n495 B.n106 585
R1252 B.n494 B.n493 585
R1253 B.n492 B.n107 585
R1254 B.n491 B.n490 585
R1255 B.n489 B.n108 585
R1256 B.n488 B.n487 585
R1257 B.n486 B.n109 585
R1258 B.n485 B.n484 585
R1259 B.n483 B.n110 585
R1260 B.n482 B.n481 585
R1261 B.n480 B.n111 585
R1262 B.n479 B.n478 585
R1263 B.n477 B.n112 585
R1264 B.n476 B.n475 585
R1265 B.n474 B.n113 585
R1266 B.n473 B.n472 585
R1267 B.n471 B.n114 585
R1268 B.n470 B.n469 585
R1269 B.n468 B.n115 585
R1270 B.n467 B.n466 585
R1271 B.n465 B.n116 585
R1272 B.n464 B.n463 585
R1273 B.n462 B.n117 585
R1274 B.n461 B.n460 585
R1275 B.n459 B.n118 585
R1276 B.n458 B.n457 585
R1277 B.n456 B.n119 585
R1278 B.n455 B.n454 585
R1279 B.n453 B.n120 585
R1280 B.n452 B.n451 585
R1281 B.n450 B.n121 585
R1282 B.n449 B.n448 585
R1283 B.n447 B.n122 585
R1284 B.n446 B.n445 585
R1285 B.n444 B.n123 585
R1286 B.n443 B.n442 585
R1287 B.n441 B.n124 585
R1288 B.n440 B.n439 585
R1289 B.n438 B.n125 585
R1290 B.n437 B.n436 585
R1291 B.n435 B.n126 585
R1292 B.n434 B.n433 585
R1293 B.n432 B.n127 585
R1294 B.n271 B.n270 585
R1295 B.n272 B.n181 585
R1296 B.n274 B.n273 585
R1297 B.n275 B.n180 585
R1298 B.n277 B.n276 585
R1299 B.n278 B.n179 585
R1300 B.n280 B.n279 585
R1301 B.n281 B.n178 585
R1302 B.n283 B.n282 585
R1303 B.n284 B.n177 585
R1304 B.n286 B.n285 585
R1305 B.n287 B.n176 585
R1306 B.n289 B.n288 585
R1307 B.n290 B.n175 585
R1308 B.n292 B.n291 585
R1309 B.n293 B.n174 585
R1310 B.n295 B.n294 585
R1311 B.n296 B.n173 585
R1312 B.n298 B.n297 585
R1313 B.n299 B.n172 585
R1314 B.n301 B.n300 585
R1315 B.n302 B.n171 585
R1316 B.n304 B.n303 585
R1317 B.n305 B.n170 585
R1318 B.n307 B.n306 585
R1319 B.n308 B.n169 585
R1320 B.n310 B.n309 585
R1321 B.n311 B.n168 585
R1322 B.n313 B.n312 585
R1323 B.n314 B.n167 585
R1324 B.n316 B.n315 585
R1325 B.n317 B.n166 585
R1326 B.n319 B.n318 585
R1327 B.n320 B.n165 585
R1328 B.n322 B.n321 585
R1329 B.n323 B.n164 585
R1330 B.n325 B.n324 585
R1331 B.n326 B.n163 585
R1332 B.n328 B.n327 585
R1333 B.n329 B.n162 585
R1334 B.n331 B.n330 585
R1335 B.n332 B.n161 585
R1336 B.n334 B.n333 585
R1337 B.n335 B.n160 585
R1338 B.n337 B.n336 585
R1339 B.n338 B.n159 585
R1340 B.n340 B.n339 585
R1341 B.n341 B.n156 585
R1342 B.n344 B.n343 585
R1343 B.n345 B.n155 585
R1344 B.n347 B.n346 585
R1345 B.n348 B.n154 585
R1346 B.n350 B.n349 585
R1347 B.n351 B.n153 585
R1348 B.n353 B.n352 585
R1349 B.n354 B.n152 585
R1350 B.n359 B.n358 585
R1351 B.n360 B.n151 585
R1352 B.n362 B.n361 585
R1353 B.n363 B.n150 585
R1354 B.n365 B.n364 585
R1355 B.n366 B.n149 585
R1356 B.n368 B.n367 585
R1357 B.n369 B.n148 585
R1358 B.n371 B.n370 585
R1359 B.n372 B.n147 585
R1360 B.n374 B.n373 585
R1361 B.n375 B.n146 585
R1362 B.n377 B.n376 585
R1363 B.n378 B.n145 585
R1364 B.n380 B.n379 585
R1365 B.n381 B.n144 585
R1366 B.n383 B.n382 585
R1367 B.n384 B.n143 585
R1368 B.n386 B.n385 585
R1369 B.n387 B.n142 585
R1370 B.n389 B.n388 585
R1371 B.n390 B.n141 585
R1372 B.n392 B.n391 585
R1373 B.n393 B.n140 585
R1374 B.n395 B.n394 585
R1375 B.n396 B.n139 585
R1376 B.n398 B.n397 585
R1377 B.n399 B.n138 585
R1378 B.n401 B.n400 585
R1379 B.n402 B.n137 585
R1380 B.n404 B.n403 585
R1381 B.n405 B.n136 585
R1382 B.n407 B.n406 585
R1383 B.n408 B.n135 585
R1384 B.n410 B.n409 585
R1385 B.n411 B.n134 585
R1386 B.n413 B.n412 585
R1387 B.n414 B.n133 585
R1388 B.n416 B.n415 585
R1389 B.n417 B.n132 585
R1390 B.n419 B.n418 585
R1391 B.n420 B.n131 585
R1392 B.n422 B.n421 585
R1393 B.n423 B.n130 585
R1394 B.n425 B.n424 585
R1395 B.n426 B.n129 585
R1396 B.n428 B.n427 585
R1397 B.n429 B.n128 585
R1398 B.n431 B.n430 585
R1399 B.n269 B.n182 585
R1400 B.n268 B.n267 585
R1401 B.n266 B.n183 585
R1402 B.n265 B.n264 585
R1403 B.n263 B.n184 585
R1404 B.n262 B.n261 585
R1405 B.n260 B.n185 585
R1406 B.n259 B.n258 585
R1407 B.n257 B.n186 585
R1408 B.n256 B.n255 585
R1409 B.n254 B.n187 585
R1410 B.n253 B.n252 585
R1411 B.n251 B.n188 585
R1412 B.n250 B.n249 585
R1413 B.n248 B.n189 585
R1414 B.n247 B.n246 585
R1415 B.n245 B.n190 585
R1416 B.n244 B.n243 585
R1417 B.n242 B.n191 585
R1418 B.n241 B.n240 585
R1419 B.n239 B.n192 585
R1420 B.n238 B.n237 585
R1421 B.n236 B.n193 585
R1422 B.n235 B.n234 585
R1423 B.n233 B.n194 585
R1424 B.n232 B.n231 585
R1425 B.n230 B.n195 585
R1426 B.n229 B.n228 585
R1427 B.n227 B.n196 585
R1428 B.n226 B.n225 585
R1429 B.n224 B.n197 585
R1430 B.n223 B.n222 585
R1431 B.n221 B.n198 585
R1432 B.n220 B.n219 585
R1433 B.n218 B.n199 585
R1434 B.n217 B.n216 585
R1435 B.n215 B.n200 585
R1436 B.n214 B.n213 585
R1437 B.n212 B.n201 585
R1438 B.n211 B.n210 585
R1439 B.n209 B.n202 585
R1440 B.n208 B.n207 585
R1441 B.n206 B.n203 585
R1442 B.n205 B.n204 585
R1443 B.n2 B.n0 585
R1444 B.n793 B.n1 585
R1445 B.n792 B.n791 585
R1446 B.n790 B.n3 585
R1447 B.n789 B.n788 585
R1448 B.n787 B.n4 585
R1449 B.n786 B.n785 585
R1450 B.n784 B.n5 585
R1451 B.n783 B.n782 585
R1452 B.n781 B.n6 585
R1453 B.n780 B.n779 585
R1454 B.n778 B.n7 585
R1455 B.n777 B.n776 585
R1456 B.n775 B.n8 585
R1457 B.n774 B.n773 585
R1458 B.n772 B.n9 585
R1459 B.n771 B.n770 585
R1460 B.n769 B.n10 585
R1461 B.n768 B.n767 585
R1462 B.n766 B.n11 585
R1463 B.n765 B.n764 585
R1464 B.n763 B.n12 585
R1465 B.n762 B.n761 585
R1466 B.n760 B.n13 585
R1467 B.n759 B.n758 585
R1468 B.n757 B.n14 585
R1469 B.n756 B.n755 585
R1470 B.n754 B.n15 585
R1471 B.n753 B.n752 585
R1472 B.n751 B.n16 585
R1473 B.n750 B.n749 585
R1474 B.n748 B.n17 585
R1475 B.n747 B.n746 585
R1476 B.n745 B.n18 585
R1477 B.n744 B.n743 585
R1478 B.n742 B.n19 585
R1479 B.n741 B.n740 585
R1480 B.n739 B.n20 585
R1481 B.n738 B.n737 585
R1482 B.n736 B.n21 585
R1483 B.n735 B.n734 585
R1484 B.n733 B.n22 585
R1485 B.n732 B.n731 585
R1486 B.n730 B.n23 585
R1487 B.n729 B.n728 585
R1488 B.n727 B.n24 585
R1489 B.n795 B.n794 585
R1490 B.n271 B.n182 492.5
R1491 B.n727 B.n726 492.5
R1492 B.n432 B.n431 492.5
R1493 B.n569 B.n82 492.5
R1494 B.n355 B.t8 473.17
R1495 B.n57 B.t1 473.17
R1496 B.n157 B.t11 473.17
R1497 B.n50 B.t4 473.17
R1498 B.n356 B.t7 412.272
R1499 B.n58 B.t2 412.272
R1500 B.n158 B.t10 412.272
R1501 B.n51 B.t5 412.272
R1502 B.n355 B.t6 328.757
R1503 B.n157 B.t9 328.757
R1504 B.n50 B.t3 328.757
R1505 B.n57 B.t0 328.757
R1506 B.n267 B.n182 163.367
R1507 B.n267 B.n266 163.367
R1508 B.n266 B.n265 163.367
R1509 B.n265 B.n184 163.367
R1510 B.n261 B.n184 163.367
R1511 B.n261 B.n260 163.367
R1512 B.n260 B.n259 163.367
R1513 B.n259 B.n186 163.367
R1514 B.n255 B.n186 163.367
R1515 B.n255 B.n254 163.367
R1516 B.n254 B.n253 163.367
R1517 B.n253 B.n188 163.367
R1518 B.n249 B.n188 163.367
R1519 B.n249 B.n248 163.367
R1520 B.n248 B.n247 163.367
R1521 B.n247 B.n190 163.367
R1522 B.n243 B.n190 163.367
R1523 B.n243 B.n242 163.367
R1524 B.n242 B.n241 163.367
R1525 B.n241 B.n192 163.367
R1526 B.n237 B.n192 163.367
R1527 B.n237 B.n236 163.367
R1528 B.n236 B.n235 163.367
R1529 B.n235 B.n194 163.367
R1530 B.n231 B.n194 163.367
R1531 B.n231 B.n230 163.367
R1532 B.n230 B.n229 163.367
R1533 B.n229 B.n196 163.367
R1534 B.n225 B.n196 163.367
R1535 B.n225 B.n224 163.367
R1536 B.n224 B.n223 163.367
R1537 B.n223 B.n198 163.367
R1538 B.n219 B.n198 163.367
R1539 B.n219 B.n218 163.367
R1540 B.n218 B.n217 163.367
R1541 B.n217 B.n200 163.367
R1542 B.n213 B.n200 163.367
R1543 B.n213 B.n212 163.367
R1544 B.n212 B.n211 163.367
R1545 B.n211 B.n202 163.367
R1546 B.n207 B.n202 163.367
R1547 B.n207 B.n206 163.367
R1548 B.n206 B.n205 163.367
R1549 B.n205 B.n2 163.367
R1550 B.n794 B.n2 163.367
R1551 B.n794 B.n793 163.367
R1552 B.n793 B.n792 163.367
R1553 B.n792 B.n3 163.367
R1554 B.n788 B.n3 163.367
R1555 B.n788 B.n787 163.367
R1556 B.n787 B.n786 163.367
R1557 B.n786 B.n5 163.367
R1558 B.n782 B.n5 163.367
R1559 B.n782 B.n781 163.367
R1560 B.n781 B.n780 163.367
R1561 B.n780 B.n7 163.367
R1562 B.n776 B.n7 163.367
R1563 B.n776 B.n775 163.367
R1564 B.n775 B.n774 163.367
R1565 B.n774 B.n9 163.367
R1566 B.n770 B.n9 163.367
R1567 B.n770 B.n769 163.367
R1568 B.n769 B.n768 163.367
R1569 B.n768 B.n11 163.367
R1570 B.n764 B.n11 163.367
R1571 B.n764 B.n763 163.367
R1572 B.n763 B.n762 163.367
R1573 B.n762 B.n13 163.367
R1574 B.n758 B.n13 163.367
R1575 B.n758 B.n757 163.367
R1576 B.n757 B.n756 163.367
R1577 B.n756 B.n15 163.367
R1578 B.n752 B.n15 163.367
R1579 B.n752 B.n751 163.367
R1580 B.n751 B.n750 163.367
R1581 B.n750 B.n17 163.367
R1582 B.n746 B.n17 163.367
R1583 B.n746 B.n745 163.367
R1584 B.n745 B.n744 163.367
R1585 B.n744 B.n19 163.367
R1586 B.n740 B.n19 163.367
R1587 B.n740 B.n739 163.367
R1588 B.n739 B.n738 163.367
R1589 B.n738 B.n21 163.367
R1590 B.n734 B.n21 163.367
R1591 B.n734 B.n733 163.367
R1592 B.n733 B.n732 163.367
R1593 B.n732 B.n23 163.367
R1594 B.n728 B.n23 163.367
R1595 B.n728 B.n727 163.367
R1596 B.n272 B.n271 163.367
R1597 B.n273 B.n272 163.367
R1598 B.n273 B.n180 163.367
R1599 B.n277 B.n180 163.367
R1600 B.n278 B.n277 163.367
R1601 B.n279 B.n278 163.367
R1602 B.n279 B.n178 163.367
R1603 B.n283 B.n178 163.367
R1604 B.n284 B.n283 163.367
R1605 B.n285 B.n284 163.367
R1606 B.n285 B.n176 163.367
R1607 B.n289 B.n176 163.367
R1608 B.n290 B.n289 163.367
R1609 B.n291 B.n290 163.367
R1610 B.n291 B.n174 163.367
R1611 B.n295 B.n174 163.367
R1612 B.n296 B.n295 163.367
R1613 B.n297 B.n296 163.367
R1614 B.n297 B.n172 163.367
R1615 B.n301 B.n172 163.367
R1616 B.n302 B.n301 163.367
R1617 B.n303 B.n302 163.367
R1618 B.n303 B.n170 163.367
R1619 B.n307 B.n170 163.367
R1620 B.n308 B.n307 163.367
R1621 B.n309 B.n308 163.367
R1622 B.n309 B.n168 163.367
R1623 B.n313 B.n168 163.367
R1624 B.n314 B.n313 163.367
R1625 B.n315 B.n314 163.367
R1626 B.n315 B.n166 163.367
R1627 B.n319 B.n166 163.367
R1628 B.n320 B.n319 163.367
R1629 B.n321 B.n320 163.367
R1630 B.n321 B.n164 163.367
R1631 B.n325 B.n164 163.367
R1632 B.n326 B.n325 163.367
R1633 B.n327 B.n326 163.367
R1634 B.n327 B.n162 163.367
R1635 B.n331 B.n162 163.367
R1636 B.n332 B.n331 163.367
R1637 B.n333 B.n332 163.367
R1638 B.n333 B.n160 163.367
R1639 B.n337 B.n160 163.367
R1640 B.n338 B.n337 163.367
R1641 B.n339 B.n338 163.367
R1642 B.n339 B.n156 163.367
R1643 B.n344 B.n156 163.367
R1644 B.n345 B.n344 163.367
R1645 B.n346 B.n345 163.367
R1646 B.n346 B.n154 163.367
R1647 B.n350 B.n154 163.367
R1648 B.n351 B.n350 163.367
R1649 B.n352 B.n351 163.367
R1650 B.n352 B.n152 163.367
R1651 B.n359 B.n152 163.367
R1652 B.n360 B.n359 163.367
R1653 B.n361 B.n360 163.367
R1654 B.n361 B.n150 163.367
R1655 B.n365 B.n150 163.367
R1656 B.n366 B.n365 163.367
R1657 B.n367 B.n366 163.367
R1658 B.n367 B.n148 163.367
R1659 B.n371 B.n148 163.367
R1660 B.n372 B.n371 163.367
R1661 B.n373 B.n372 163.367
R1662 B.n373 B.n146 163.367
R1663 B.n377 B.n146 163.367
R1664 B.n378 B.n377 163.367
R1665 B.n379 B.n378 163.367
R1666 B.n379 B.n144 163.367
R1667 B.n383 B.n144 163.367
R1668 B.n384 B.n383 163.367
R1669 B.n385 B.n384 163.367
R1670 B.n385 B.n142 163.367
R1671 B.n389 B.n142 163.367
R1672 B.n390 B.n389 163.367
R1673 B.n391 B.n390 163.367
R1674 B.n391 B.n140 163.367
R1675 B.n395 B.n140 163.367
R1676 B.n396 B.n395 163.367
R1677 B.n397 B.n396 163.367
R1678 B.n397 B.n138 163.367
R1679 B.n401 B.n138 163.367
R1680 B.n402 B.n401 163.367
R1681 B.n403 B.n402 163.367
R1682 B.n403 B.n136 163.367
R1683 B.n407 B.n136 163.367
R1684 B.n408 B.n407 163.367
R1685 B.n409 B.n408 163.367
R1686 B.n409 B.n134 163.367
R1687 B.n413 B.n134 163.367
R1688 B.n414 B.n413 163.367
R1689 B.n415 B.n414 163.367
R1690 B.n415 B.n132 163.367
R1691 B.n419 B.n132 163.367
R1692 B.n420 B.n419 163.367
R1693 B.n421 B.n420 163.367
R1694 B.n421 B.n130 163.367
R1695 B.n425 B.n130 163.367
R1696 B.n426 B.n425 163.367
R1697 B.n427 B.n426 163.367
R1698 B.n427 B.n128 163.367
R1699 B.n431 B.n128 163.367
R1700 B.n433 B.n432 163.367
R1701 B.n433 B.n126 163.367
R1702 B.n437 B.n126 163.367
R1703 B.n438 B.n437 163.367
R1704 B.n439 B.n438 163.367
R1705 B.n439 B.n124 163.367
R1706 B.n443 B.n124 163.367
R1707 B.n444 B.n443 163.367
R1708 B.n445 B.n444 163.367
R1709 B.n445 B.n122 163.367
R1710 B.n449 B.n122 163.367
R1711 B.n450 B.n449 163.367
R1712 B.n451 B.n450 163.367
R1713 B.n451 B.n120 163.367
R1714 B.n455 B.n120 163.367
R1715 B.n456 B.n455 163.367
R1716 B.n457 B.n456 163.367
R1717 B.n457 B.n118 163.367
R1718 B.n461 B.n118 163.367
R1719 B.n462 B.n461 163.367
R1720 B.n463 B.n462 163.367
R1721 B.n463 B.n116 163.367
R1722 B.n467 B.n116 163.367
R1723 B.n468 B.n467 163.367
R1724 B.n469 B.n468 163.367
R1725 B.n469 B.n114 163.367
R1726 B.n473 B.n114 163.367
R1727 B.n474 B.n473 163.367
R1728 B.n475 B.n474 163.367
R1729 B.n475 B.n112 163.367
R1730 B.n479 B.n112 163.367
R1731 B.n480 B.n479 163.367
R1732 B.n481 B.n480 163.367
R1733 B.n481 B.n110 163.367
R1734 B.n485 B.n110 163.367
R1735 B.n486 B.n485 163.367
R1736 B.n487 B.n486 163.367
R1737 B.n487 B.n108 163.367
R1738 B.n491 B.n108 163.367
R1739 B.n492 B.n491 163.367
R1740 B.n493 B.n492 163.367
R1741 B.n493 B.n106 163.367
R1742 B.n497 B.n106 163.367
R1743 B.n498 B.n497 163.367
R1744 B.n499 B.n498 163.367
R1745 B.n499 B.n104 163.367
R1746 B.n503 B.n104 163.367
R1747 B.n504 B.n503 163.367
R1748 B.n505 B.n504 163.367
R1749 B.n505 B.n102 163.367
R1750 B.n509 B.n102 163.367
R1751 B.n510 B.n509 163.367
R1752 B.n511 B.n510 163.367
R1753 B.n511 B.n100 163.367
R1754 B.n515 B.n100 163.367
R1755 B.n516 B.n515 163.367
R1756 B.n517 B.n516 163.367
R1757 B.n517 B.n98 163.367
R1758 B.n521 B.n98 163.367
R1759 B.n522 B.n521 163.367
R1760 B.n523 B.n522 163.367
R1761 B.n523 B.n96 163.367
R1762 B.n527 B.n96 163.367
R1763 B.n528 B.n527 163.367
R1764 B.n529 B.n528 163.367
R1765 B.n529 B.n94 163.367
R1766 B.n533 B.n94 163.367
R1767 B.n534 B.n533 163.367
R1768 B.n535 B.n534 163.367
R1769 B.n535 B.n92 163.367
R1770 B.n539 B.n92 163.367
R1771 B.n540 B.n539 163.367
R1772 B.n541 B.n540 163.367
R1773 B.n541 B.n90 163.367
R1774 B.n545 B.n90 163.367
R1775 B.n546 B.n545 163.367
R1776 B.n547 B.n546 163.367
R1777 B.n547 B.n88 163.367
R1778 B.n551 B.n88 163.367
R1779 B.n552 B.n551 163.367
R1780 B.n553 B.n552 163.367
R1781 B.n553 B.n86 163.367
R1782 B.n557 B.n86 163.367
R1783 B.n558 B.n557 163.367
R1784 B.n559 B.n558 163.367
R1785 B.n559 B.n84 163.367
R1786 B.n563 B.n84 163.367
R1787 B.n564 B.n563 163.367
R1788 B.n565 B.n564 163.367
R1789 B.n565 B.n82 163.367
R1790 B.n726 B.n25 163.367
R1791 B.n722 B.n25 163.367
R1792 B.n722 B.n721 163.367
R1793 B.n721 B.n720 163.367
R1794 B.n720 B.n27 163.367
R1795 B.n716 B.n27 163.367
R1796 B.n716 B.n715 163.367
R1797 B.n715 B.n714 163.367
R1798 B.n714 B.n29 163.367
R1799 B.n710 B.n29 163.367
R1800 B.n710 B.n709 163.367
R1801 B.n709 B.n708 163.367
R1802 B.n708 B.n31 163.367
R1803 B.n704 B.n31 163.367
R1804 B.n704 B.n703 163.367
R1805 B.n703 B.n702 163.367
R1806 B.n702 B.n33 163.367
R1807 B.n698 B.n33 163.367
R1808 B.n698 B.n697 163.367
R1809 B.n697 B.n696 163.367
R1810 B.n696 B.n35 163.367
R1811 B.n692 B.n35 163.367
R1812 B.n692 B.n691 163.367
R1813 B.n691 B.n690 163.367
R1814 B.n690 B.n37 163.367
R1815 B.n686 B.n37 163.367
R1816 B.n686 B.n685 163.367
R1817 B.n685 B.n684 163.367
R1818 B.n684 B.n39 163.367
R1819 B.n680 B.n39 163.367
R1820 B.n680 B.n679 163.367
R1821 B.n679 B.n678 163.367
R1822 B.n678 B.n41 163.367
R1823 B.n674 B.n41 163.367
R1824 B.n674 B.n673 163.367
R1825 B.n673 B.n672 163.367
R1826 B.n672 B.n43 163.367
R1827 B.n668 B.n43 163.367
R1828 B.n668 B.n667 163.367
R1829 B.n667 B.n666 163.367
R1830 B.n666 B.n45 163.367
R1831 B.n662 B.n45 163.367
R1832 B.n662 B.n661 163.367
R1833 B.n661 B.n660 163.367
R1834 B.n660 B.n47 163.367
R1835 B.n656 B.n47 163.367
R1836 B.n656 B.n655 163.367
R1837 B.n655 B.n654 163.367
R1838 B.n654 B.n49 163.367
R1839 B.n650 B.n49 163.367
R1840 B.n650 B.n649 163.367
R1841 B.n649 B.n648 163.367
R1842 B.n648 B.n54 163.367
R1843 B.n644 B.n54 163.367
R1844 B.n644 B.n643 163.367
R1845 B.n643 B.n642 163.367
R1846 B.n642 B.n56 163.367
R1847 B.n637 B.n56 163.367
R1848 B.n637 B.n636 163.367
R1849 B.n636 B.n635 163.367
R1850 B.n635 B.n60 163.367
R1851 B.n631 B.n60 163.367
R1852 B.n631 B.n630 163.367
R1853 B.n630 B.n629 163.367
R1854 B.n629 B.n62 163.367
R1855 B.n625 B.n62 163.367
R1856 B.n625 B.n624 163.367
R1857 B.n624 B.n623 163.367
R1858 B.n623 B.n64 163.367
R1859 B.n619 B.n64 163.367
R1860 B.n619 B.n618 163.367
R1861 B.n618 B.n617 163.367
R1862 B.n617 B.n66 163.367
R1863 B.n613 B.n66 163.367
R1864 B.n613 B.n612 163.367
R1865 B.n612 B.n611 163.367
R1866 B.n611 B.n68 163.367
R1867 B.n607 B.n68 163.367
R1868 B.n607 B.n606 163.367
R1869 B.n606 B.n605 163.367
R1870 B.n605 B.n70 163.367
R1871 B.n601 B.n70 163.367
R1872 B.n601 B.n600 163.367
R1873 B.n600 B.n599 163.367
R1874 B.n599 B.n72 163.367
R1875 B.n595 B.n72 163.367
R1876 B.n595 B.n594 163.367
R1877 B.n594 B.n593 163.367
R1878 B.n593 B.n74 163.367
R1879 B.n589 B.n74 163.367
R1880 B.n589 B.n588 163.367
R1881 B.n588 B.n587 163.367
R1882 B.n587 B.n76 163.367
R1883 B.n583 B.n76 163.367
R1884 B.n583 B.n582 163.367
R1885 B.n582 B.n581 163.367
R1886 B.n581 B.n78 163.367
R1887 B.n577 B.n78 163.367
R1888 B.n577 B.n576 163.367
R1889 B.n576 B.n575 163.367
R1890 B.n575 B.n80 163.367
R1891 B.n571 B.n80 163.367
R1892 B.n571 B.n570 163.367
R1893 B.n570 B.n569 163.367
R1894 B.n356 B.n355 60.8975
R1895 B.n158 B.n157 60.8975
R1896 B.n51 B.n50 60.8975
R1897 B.n58 B.n57 60.8975
R1898 B.n357 B.n356 59.5399
R1899 B.n342 B.n158 59.5399
R1900 B.n52 B.n51 59.5399
R1901 B.n640 B.n58 59.5399
R1902 B.n725 B.n24 32.0005
R1903 B.n568 B.n567 32.0005
R1904 B.n430 B.n127 32.0005
R1905 B.n270 B.n269 32.0005
R1906 B B.n795 18.0485
R1907 B.n725 B.n724 10.6151
R1908 B.n724 B.n723 10.6151
R1909 B.n723 B.n26 10.6151
R1910 B.n719 B.n26 10.6151
R1911 B.n719 B.n718 10.6151
R1912 B.n718 B.n717 10.6151
R1913 B.n717 B.n28 10.6151
R1914 B.n713 B.n28 10.6151
R1915 B.n713 B.n712 10.6151
R1916 B.n712 B.n711 10.6151
R1917 B.n711 B.n30 10.6151
R1918 B.n707 B.n30 10.6151
R1919 B.n707 B.n706 10.6151
R1920 B.n706 B.n705 10.6151
R1921 B.n705 B.n32 10.6151
R1922 B.n701 B.n32 10.6151
R1923 B.n701 B.n700 10.6151
R1924 B.n700 B.n699 10.6151
R1925 B.n699 B.n34 10.6151
R1926 B.n695 B.n34 10.6151
R1927 B.n695 B.n694 10.6151
R1928 B.n694 B.n693 10.6151
R1929 B.n693 B.n36 10.6151
R1930 B.n689 B.n36 10.6151
R1931 B.n689 B.n688 10.6151
R1932 B.n688 B.n687 10.6151
R1933 B.n687 B.n38 10.6151
R1934 B.n683 B.n38 10.6151
R1935 B.n683 B.n682 10.6151
R1936 B.n682 B.n681 10.6151
R1937 B.n681 B.n40 10.6151
R1938 B.n677 B.n40 10.6151
R1939 B.n677 B.n676 10.6151
R1940 B.n676 B.n675 10.6151
R1941 B.n675 B.n42 10.6151
R1942 B.n671 B.n42 10.6151
R1943 B.n671 B.n670 10.6151
R1944 B.n670 B.n669 10.6151
R1945 B.n669 B.n44 10.6151
R1946 B.n665 B.n44 10.6151
R1947 B.n665 B.n664 10.6151
R1948 B.n664 B.n663 10.6151
R1949 B.n663 B.n46 10.6151
R1950 B.n659 B.n46 10.6151
R1951 B.n659 B.n658 10.6151
R1952 B.n658 B.n657 10.6151
R1953 B.n657 B.n48 10.6151
R1954 B.n653 B.n652 10.6151
R1955 B.n652 B.n651 10.6151
R1956 B.n651 B.n53 10.6151
R1957 B.n647 B.n53 10.6151
R1958 B.n647 B.n646 10.6151
R1959 B.n646 B.n645 10.6151
R1960 B.n645 B.n55 10.6151
R1961 B.n641 B.n55 10.6151
R1962 B.n639 B.n638 10.6151
R1963 B.n638 B.n59 10.6151
R1964 B.n634 B.n59 10.6151
R1965 B.n634 B.n633 10.6151
R1966 B.n633 B.n632 10.6151
R1967 B.n632 B.n61 10.6151
R1968 B.n628 B.n61 10.6151
R1969 B.n628 B.n627 10.6151
R1970 B.n627 B.n626 10.6151
R1971 B.n626 B.n63 10.6151
R1972 B.n622 B.n63 10.6151
R1973 B.n622 B.n621 10.6151
R1974 B.n621 B.n620 10.6151
R1975 B.n620 B.n65 10.6151
R1976 B.n616 B.n65 10.6151
R1977 B.n616 B.n615 10.6151
R1978 B.n615 B.n614 10.6151
R1979 B.n614 B.n67 10.6151
R1980 B.n610 B.n67 10.6151
R1981 B.n610 B.n609 10.6151
R1982 B.n609 B.n608 10.6151
R1983 B.n608 B.n69 10.6151
R1984 B.n604 B.n69 10.6151
R1985 B.n604 B.n603 10.6151
R1986 B.n603 B.n602 10.6151
R1987 B.n602 B.n71 10.6151
R1988 B.n598 B.n71 10.6151
R1989 B.n598 B.n597 10.6151
R1990 B.n597 B.n596 10.6151
R1991 B.n596 B.n73 10.6151
R1992 B.n592 B.n73 10.6151
R1993 B.n592 B.n591 10.6151
R1994 B.n591 B.n590 10.6151
R1995 B.n590 B.n75 10.6151
R1996 B.n586 B.n75 10.6151
R1997 B.n586 B.n585 10.6151
R1998 B.n585 B.n584 10.6151
R1999 B.n584 B.n77 10.6151
R2000 B.n580 B.n77 10.6151
R2001 B.n580 B.n579 10.6151
R2002 B.n579 B.n578 10.6151
R2003 B.n578 B.n79 10.6151
R2004 B.n574 B.n79 10.6151
R2005 B.n574 B.n573 10.6151
R2006 B.n573 B.n572 10.6151
R2007 B.n572 B.n81 10.6151
R2008 B.n568 B.n81 10.6151
R2009 B.n434 B.n127 10.6151
R2010 B.n435 B.n434 10.6151
R2011 B.n436 B.n435 10.6151
R2012 B.n436 B.n125 10.6151
R2013 B.n440 B.n125 10.6151
R2014 B.n441 B.n440 10.6151
R2015 B.n442 B.n441 10.6151
R2016 B.n442 B.n123 10.6151
R2017 B.n446 B.n123 10.6151
R2018 B.n447 B.n446 10.6151
R2019 B.n448 B.n447 10.6151
R2020 B.n448 B.n121 10.6151
R2021 B.n452 B.n121 10.6151
R2022 B.n453 B.n452 10.6151
R2023 B.n454 B.n453 10.6151
R2024 B.n454 B.n119 10.6151
R2025 B.n458 B.n119 10.6151
R2026 B.n459 B.n458 10.6151
R2027 B.n460 B.n459 10.6151
R2028 B.n460 B.n117 10.6151
R2029 B.n464 B.n117 10.6151
R2030 B.n465 B.n464 10.6151
R2031 B.n466 B.n465 10.6151
R2032 B.n466 B.n115 10.6151
R2033 B.n470 B.n115 10.6151
R2034 B.n471 B.n470 10.6151
R2035 B.n472 B.n471 10.6151
R2036 B.n472 B.n113 10.6151
R2037 B.n476 B.n113 10.6151
R2038 B.n477 B.n476 10.6151
R2039 B.n478 B.n477 10.6151
R2040 B.n478 B.n111 10.6151
R2041 B.n482 B.n111 10.6151
R2042 B.n483 B.n482 10.6151
R2043 B.n484 B.n483 10.6151
R2044 B.n484 B.n109 10.6151
R2045 B.n488 B.n109 10.6151
R2046 B.n489 B.n488 10.6151
R2047 B.n490 B.n489 10.6151
R2048 B.n490 B.n107 10.6151
R2049 B.n494 B.n107 10.6151
R2050 B.n495 B.n494 10.6151
R2051 B.n496 B.n495 10.6151
R2052 B.n496 B.n105 10.6151
R2053 B.n500 B.n105 10.6151
R2054 B.n501 B.n500 10.6151
R2055 B.n502 B.n501 10.6151
R2056 B.n502 B.n103 10.6151
R2057 B.n506 B.n103 10.6151
R2058 B.n507 B.n506 10.6151
R2059 B.n508 B.n507 10.6151
R2060 B.n508 B.n101 10.6151
R2061 B.n512 B.n101 10.6151
R2062 B.n513 B.n512 10.6151
R2063 B.n514 B.n513 10.6151
R2064 B.n514 B.n99 10.6151
R2065 B.n518 B.n99 10.6151
R2066 B.n519 B.n518 10.6151
R2067 B.n520 B.n519 10.6151
R2068 B.n520 B.n97 10.6151
R2069 B.n524 B.n97 10.6151
R2070 B.n525 B.n524 10.6151
R2071 B.n526 B.n525 10.6151
R2072 B.n526 B.n95 10.6151
R2073 B.n530 B.n95 10.6151
R2074 B.n531 B.n530 10.6151
R2075 B.n532 B.n531 10.6151
R2076 B.n532 B.n93 10.6151
R2077 B.n536 B.n93 10.6151
R2078 B.n537 B.n536 10.6151
R2079 B.n538 B.n537 10.6151
R2080 B.n538 B.n91 10.6151
R2081 B.n542 B.n91 10.6151
R2082 B.n543 B.n542 10.6151
R2083 B.n544 B.n543 10.6151
R2084 B.n544 B.n89 10.6151
R2085 B.n548 B.n89 10.6151
R2086 B.n549 B.n548 10.6151
R2087 B.n550 B.n549 10.6151
R2088 B.n550 B.n87 10.6151
R2089 B.n554 B.n87 10.6151
R2090 B.n555 B.n554 10.6151
R2091 B.n556 B.n555 10.6151
R2092 B.n556 B.n85 10.6151
R2093 B.n560 B.n85 10.6151
R2094 B.n561 B.n560 10.6151
R2095 B.n562 B.n561 10.6151
R2096 B.n562 B.n83 10.6151
R2097 B.n566 B.n83 10.6151
R2098 B.n567 B.n566 10.6151
R2099 B.n270 B.n181 10.6151
R2100 B.n274 B.n181 10.6151
R2101 B.n275 B.n274 10.6151
R2102 B.n276 B.n275 10.6151
R2103 B.n276 B.n179 10.6151
R2104 B.n280 B.n179 10.6151
R2105 B.n281 B.n280 10.6151
R2106 B.n282 B.n281 10.6151
R2107 B.n282 B.n177 10.6151
R2108 B.n286 B.n177 10.6151
R2109 B.n287 B.n286 10.6151
R2110 B.n288 B.n287 10.6151
R2111 B.n288 B.n175 10.6151
R2112 B.n292 B.n175 10.6151
R2113 B.n293 B.n292 10.6151
R2114 B.n294 B.n293 10.6151
R2115 B.n294 B.n173 10.6151
R2116 B.n298 B.n173 10.6151
R2117 B.n299 B.n298 10.6151
R2118 B.n300 B.n299 10.6151
R2119 B.n300 B.n171 10.6151
R2120 B.n304 B.n171 10.6151
R2121 B.n305 B.n304 10.6151
R2122 B.n306 B.n305 10.6151
R2123 B.n306 B.n169 10.6151
R2124 B.n310 B.n169 10.6151
R2125 B.n311 B.n310 10.6151
R2126 B.n312 B.n311 10.6151
R2127 B.n312 B.n167 10.6151
R2128 B.n316 B.n167 10.6151
R2129 B.n317 B.n316 10.6151
R2130 B.n318 B.n317 10.6151
R2131 B.n318 B.n165 10.6151
R2132 B.n322 B.n165 10.6151
R2133 B.n323 B.n322 10.6151
R2134 B.n324 B.n323 10.6151
R2135 B.n324 B.n163 10.6151
R2136 B.n328 B.n163 10.6151
R2137 B.n329 B.n328 10.6151
R2138 B.n330 B.n329 10.6151
R2139 B.n330 B.n161 10.6151
R2140 B.n334 B.n161 10.6151
R2141 B.n335 B.n334 10.6151
R2142 B.n336 B.n335 10.6151
R2143 B.n336 B.n159 10.6151
R2144 B.n340 B.n159 10.6151
R2145 B.n341 B.n340 10.6151
R2146 B.n343 B.n155 10.6151
R2147 B.n347 B.n155 10.6151
R2148 B.n348 B.n347 10.6151
R2149 B.n349 B.n348 10.6151
R2150 B.n349 B.n153 10.6151
R2151 B.n353 B.n153 10.6151
R2152 B.n354 B.n353 10.6151
R2153 B.n358 B.n354 10.6151
R2154 B.n362 B.n151 10.6151
R2155 B.n363 B.n362 10.6151
R2156 B.n364 B.n363 10.6151
R2157 B.n364 B.n149 10.6151
R2158 B.n368 B.n149 10.6151
R2159 B.n369 B.n368 10.6151
R2160 B.n370 B.n369 10.6151
R2161 B.n370 B.n147 10.6151
R2162 B.n374 B.n147 10.6151
R2163 B.n375 B.n374 10.6151
R2164 B.n376 B.n375 10.6151
R2165 B.n376 B.n145 10.6151
R2166 B.n380 B.n145 10.6151
R2167 B.n381 B.n380 10.6151
R2168 B.n382 B.n381 10.6151
R2169 B.n382 B.n143 10.6151
R2170 B.n386 B.n143 10.6151
R2171 B.n387 B.n386 10.6151
R2172 B.n388 B.n387 10.6151
R2173 B.n388 B.n141 10.6151
R2174 B.n392 B.n141 10.6151
R2175 B.n393 B.n392 10.6151
R2176 B.n394 B.n393 10.6151
R2177 B.n394 B.n139 10.6151
R2178 B.n398 B.n139 10.6151
R2179 B.n399 B.n398 10.6151
R2180 B.n400 B.n399 10.6151
R2181 B.n400 B.n137 10.6151
R2182 B.n404 B.n137 10.6151
R2183 B.n405 B.n404 10.6151
R2184 B.n406 B.n405 10.6151
R2185 B.n406 B.n135 10.6151
R2186 B.n410 B.n135 10.6151
R2187 B.n411 B.n410 10.6151
R2188 B.n412 B.n411 10.6151
R2189 B.n412 B.n133 10.6151
R2190 B.n416 B.n133 10.6151
R2191 B.n417 B.n416 10.6151
R2192 B.n418 B.n417 10.6151
R2193 B.n418 B.n131 10.6151
R2194 B.n422 B.n131 10.6151
R2195 B.n423 B.n422 10.6151
R2196 B.n424 B.n423 10.6151
R2197 B.n424 B.n129 10.6151
R2198 B.n428 B.n129 10.6151
R2199 B.n429 B.n428 10.6151
R2200 B.n430 B.n429 10.6151
R2201 B.n269 B.n268 10.6151
R2202 B.n268 B.n183 10.6151
R2203 B.n264 B.n183 10.6151
R2204 B.n264 B.n263 10.6151
R2205 B.n263 B.n262 10.6151
R2206 B.n262 B.n185 10.6151
R2207 B.n258 B.n185 10.6151
R2208 B.n258 B.n257 10.6151
R2209 B.n257 B.n256 10.6151
R2210 B.n256 B.n187 10.6151
R2211 B.n252 B.n187 10.6151
R2212 B.n252 B.n251 10.6151
R2213 B.n251 B.n250 10.6151
R2214 B.n250 B.n189 10.6151
R2215 B.n246 B.n189 10.6151
R2216 B.n246 B.n245 10.6151
R2217 B.n245 B.n244 10.6151
R2218 B.n244 B.n191 10.6151
R2219 B.n240 B.n191 10.6151
R2220 B.n240 B.n239 10.6151
R2221 B.n239 B.n238 10.6151
R2222 B.n238 B.n193 10.6151
R2223 B.n234 B.n193 10.6151
R2224 B.n234 B.n233 10.6151
R2225 B.n233 B.n232 10.6151
R2226 B.n232 B.n195 10.6151
R2227 B.n228 B.n195 10.6151
R2228 B.n228 B.n227 10.6151
R2229 B.n227 B.n226 10.6151
R2230 B.n226 B.n197 10.6151
R2231 B.n222 B.n197 10.6151
R2232 B.n222 B.n221 10.6151
R2233 B.n221 B.n220 10.6151
R2234 B.n220 B.n199 10.6151
R2235 B.n216 B.n199 10.6151
R2236 B.n216 B.n215 10.6151
R2237 B.n215 B.n214 10.6151
R2238 B.n214 B.n201 10.6151
R2239 B.n210 B.n201 10.6151
R2240 B.n210 B.n209 10.6151
R2241 B.n209 B.n208 10.6151
R2242 B.n208 B.n203 10.6151
R2243 B.n204 B.n203 10.6151
R2244 B.n204 B.n0 10.6151
R2245 B.n791 B.n1 10.6151
R2246 B.n791 B.n790 10.6151
R2247 B.n790 B.n789 10.6151
R2248 B.n789 B.n4 10.6151
R2249 B.n785 B.n4 10.6151
R2250 B.n785 B.n784 10.6151
R2251 B.n784 B.n783 10.6151
R2252 B.n783 B.n6 10.6151
R2253 B.n779 B.n6 10.6151
R2254 B.n779 B.n778 10.6151
R2255 B.n778 B.n777 10.6151
R2256 B.n777 B.n8 10.6151
R2257 B.n773 B.n8 10.6151
R2258 B.n773 B.n772 10.6151
R2259 B.n772 B.n771 10.6151
R2260 B.n771 B.n10 10.6151
R2261 B.n767 B.n10 10.6151
R2262 B.n767 B.n766 10.6151
R2263 B.n766 B.n765 10.6151
R2264 B.n765 B.n12 10.6151
R2265 B.n761 B.n12 10.6151
R2266 B.n761 B.n760 10.6151
R2267 B.n760 B.n759 10.6151
R2268 B.n759 B.n14 10.6151
R2269 B.n755 B.n14 10.6151
R2270 B.n755 B.n754 10.6151
R2271 B.n754 B.n753 10.6151
R2272 B.n753 B.n16 10.6151
R2273 B.n749 B.n16 10.6151
R2274 B.n749 B.n748 10.6151
R2275 B.n748 B.n747 10.6151
R2276 B.n747 B.n18 10.6151
R2277 B.n743 B.n18 10.6151
R2278 B.n743 B.n742 10.6151
R2279 B.n742 B.n741 10.6151
R2280 B.n741 B.n20 10.6151
R2281 B.n737 B.n20 10.6151
R2282 B.n737 B.n736 10.6151
R2283 B.n736 B.n735 10.6151
R2284 B.n735 B.n22 10.6151
R2285 B.n731 B.n22 10.6151
R2286 B.n731 B.n730 10.6151
R2287 B.n730 B.n729 10.6151
R2288 B.n729 B.n24 10.6151
R2289 B.n653 B.n52 6.5566
R2290 B.n641 B.n640 6.5566
R2291 B.n343 B.n342 6.5566
R2292 B.n358 B.n357 6.5566
R2293 B.n52 B.n48 4.05904
R2294 B.n640 B.n639 4.05904
R2295 B.n342 B.n341 4.05904
R2296 B.n357 B.n151 4.05904
R2297 B.n795 B.n0 2.81026
R2298 B.n795 B.n1 2.81026
C0 B VP 1.993f
C1 VP VDD2 0.476517f
C2 VN VTAIL 8.03295f
C3 VTAIL w_n3482_n3776# 3.27099f
C4 VN w_n3482_n3776# 6.67225f
C5 VTAIL VDD1 8.49293f
C6 B VTAIL 4.24174f
C7 VTAIL VDD2 8.54495f
C8 VN VDD1 0.151267f
C9 VP VTAIL 8.04725f
C10 B VN 1.23935f
C11 w_n3482_n3776# VDD1 2.48184f
C12 VN VDD2 7.91679f
C13 B w_n3482_n3776# 10.5383f
C14 VP VN 7.50093f
C15 w_n3482_n3776# VDD2 2.5736f
C16 VP w_n3482_n3776# 7.12301f
C17 B VDD1 2.31008f
C18 VDD1 VDD2 1.48842f
C19 VP VDD1 8.238559f
C20 B VDD2 2.3892f
C21 VDD2 VSUBS 2.008355f
C22 VDD1 VSUBS 1.960518f
C23 VTAIL VSUBS 1.303317f
C24 VN VSUBS 6.09409f
C25 VP VSUBS 3.165581f
C26 B VSUBS 5.018094f
C27 w_n3482_n3776# VSUBS 0.161412p
C28 B.n0 VSUBS 0.004769f
C29 B.n1 VSUBS 0.004769f
C30 B.n2 VSUBS 0.007541f
C31 B.n3 VSUBS 0.007541f
C32 B.n4 VSUBS 0.007541f
C33 B.n5 VSUBS 0.007541f
C34 B.n6 VSUBS 0.007541f
C35 B.n7 VSUBS 0.007541f
C36 B.n8 VSUBS 0.007541f
C37 B.n9 VSUBS 0.007541f
C38 B.n10 VSUBS 0.007541f
C39 B.n11 VSUBS 0.007541f
C40 B.n12 VSUBS 0.007541f
C41 B.n13 VSUBS 0.007541f
C42 B.n14 VSUBS 0.007541f
C43 B.n15 VSUBS 0.007541f
C44 B.n16 VSUBS 0.007541f
C45 B.n17 VSUBS 0.007541f
C46 B.n18 VSUBS 0.007541f
C47 B.n19 VSUBS 0.007541f
C48 B.n20 VSUBS 0.007541f
C49 B.n21 VSUBS 0.007541f
C50 B.n22 VSUBS 0.007541f
C51 B.n23 VSUBS 0.007541f
C52 B.n24 VSUBS 0.016867f
C53 B.n25 VSUBS 0.007541f
C54 B.n26 VSUBS 0.007541f
C55 B.n27 VSUBS 0.007541f
C56 B.n28 VSUBS 0.007541f
C57 B.n29 VSUBS 0.007541f
C58 B.n30 VSUBS 0.007541f
C59 B.n31 VSUBS 0.007541f
C60 B.n32 VSUBS 0.007541f
C61 B.n33 VSUBS 0.007541f
C62 B.n34 VSUBS 0.007541f
C63 B.n35 VSUBS 0.007541f
C64 B.n36 VSUBS 0.007541f
C65 B.n37 VSUBS 0.007541f
C66 B.n38 VSUBS 0.007541f
C67 B.n39 VSUBS 0.007541f
C68 B.n40 VSUBS 0.007541f
C69 B.n41 VSUBS 0.007541f
C70 B.n42 VSUBS 0.007541f
C71 B.n43 VSUBS 0.007541f
C72 B.n44 VSUBS 0.007541f
C73 B.n45 VSUBS 0.007541f
C74 B.n46 VSUBS 0.007541f
C75 B.n47 VSUBS 0.007541f
C76 B.n48 VSUBS 0.005212f
C77 B.n49 VSUBS 0.007541f
C78 B.t5 VSUBS 0.277071f
C79 B.t4 VSUBS 0.314547f
C80 B.t3 VSUBS 1.92714f
C81 B.n50 VSUBS 0.494709f
C82 B.n51 VSUBS 0.30195f
C83 B.n52 VSUBS 0.017472f
C84 B.n53 VSUBS 0.007541f
C85 B.n54 VSUBS 0.007541f
C86 B.n55 VSUBS 0.007541f
C87 B.n56 VSUBS 0.007541f
C88 B.t2 VSUBS 0.277074f
C89 B.t1 VSUBS 0.314551f
C90 B.t0 VSUBS 1.92714f
C91 B.n57 VSUBS 0.494706f
C92 B.n58 VSUBS 0.301947f
C93 B.n59 VSUBS 0.007541f
C94 B.n60 VSUBS 0.007541f
C95 B.n61 VSUBS 0.007541f
C96 B.n62 VSUBS 0.007541f
C97 B.n63 VSUBS 0.007541f
C98 B.n64 VSUBS 0.007541f
C99 B.n65 VSUBS 0.007541f
C100 B.n66 VSUBS 0.007541f
C101 B.n67 VSUBS 0.007541f
C102 B.n68 VSUBS 0.007541f
C103 B.n69 VSUBS 0.007541f
C104 B.n70 VSUBS 0.007541f
C105 B.n71 VSUBS 0.007541f
C106 B.n72 VSUBS 0.007541f
C107 B.n73 VSUBS 0.007541f
C108 B.n74 VSUBS 0.007541f
C109 B.n75 VSUBS 0.007541f
C110 B.n76 VSUBS 0.007541f
C111 B.n77 VSUBS 0.007541f
C112 B.n78 VSUBS 0.007541f
C113 B.n79 VSUBS 0.007541f
C114 B.n80 VSUBS 0.007541f
C115 B.n81 VSUBS 0.007541f
C116 B.n82 VSUBS 0.016867f
C117 B.n83 VSUBS 0.007541f
C118 B.n84 VSUBS 0.007541f
C119 B.n85 VSUBS 0.007541f
C120 B.n86 VSUBS 0.007541f
C121 B.n87 VSUBS 0.007541f
C122 B.n88 VSUBS 0.007541f
C123 B.n89 VSUBS 0.007541f
C124 B.n90 VSUBS 0.007541f
C125 B.n91 VSUBS 0.007541f
C126 B.n92 VSUBS 0.007541f
C127 B.n93 VSUBS 0.007541f
C128 B.n94 VSUBS 0.007541f
C129 B.n95 VSUBS 0.007541f
C130 B.n96 VSUBS 0.007541f
C131 B.n97 VSUBS 0.007541f
C132 B.n98 VSUBS 0.007541f
C133 B.n99 VSUBS 0.007541f
C134 B.n100 VSUBS 0.007541f
C135 B.n101 VSUBS 0.007541f
C136 B.n102 VSUBS 0.007541f
C137 B.n103 VSUBS 0.007541f
C138 B.n104 VSUBS 0.007541f
C139 B.n105 VSUBS 0.007541f
C140 B.n106 VSUBS 0.007541f
C141 B.n107 VSUBS 0.007541f
C142 B.n108 VSUBS 0.007541f
C143 B.n109 VSUBS 0.007541f
C144 B.n110 VSUBS 0.007541f
C145 B.n111 VSUBS 0.007541f
C146 B.n112 VSUBS 0.007541f
C147 B.n113 VSUBS 0.007541f
C148 B.n114 VSUBS 0.007541f
C149 B.n115 VSUBS 0.007541f
C150 B.n116 VSUBS 0.007541f
C151 B.n117 VSUBS 0.007541f
C152 B.n118 VSUBS 0.007541f
C153 B.n119 VSUBS 0.007541f
C154 B.n120 VSUBS 0.007541f
C155 B.n121 VSUBS 0.007541f
C156 B.n122 VSUBS 0.007541f
C157 B.n123 VSUBS 0.007541f
C158 B.n124 VSUBS 0.007541f
C159 B.n125 VSUBS 0.007541f
C160 B.n126 VSUBS 0.007541f
C161 B.n127 VSUBS 0.016867f
C162 B.n128 VSUBS 0.007541f
C163 B.n129 VSUBS 0.007541f
C164 B.n130 VSUBS 0.007541f
C165 B.n131 VSUBS 0.007541f
C166 B.n132 VSUBS 0.007541f
C167 B.n133 VSUBS 0.007541f
C168 B.n134 VSUBS 0.007541f
C169 B.n135 VSUBS 0.007541f
C170 B.n136 VSUBS 0.007541f
C171 B.n137 VSUBS 0.007541f
C172 B.n138 VSUBS 0.007541f
C173 B.n139 VSUBS 0.007541f
C174 B.n140 VSUBS 0.007541f
C175 B.n141 VSUBS 0.007541f
C176 B.n142 VSUBS 0.007541f
C177 B.n143 VSUBS 0.007541f
C178 B.n144 VSUBS 0.007541f
C179 B.n145 VSUBS 0.007541f
C180 B.n146 VSUBS 0.007541f
C181 B.n147 VSUBS 0.007541f
C182 B.n148 VSUBS 0.007541f
C183 B.n149 VSUBS 0.007541f
C184 B.n150 VSUBS 0.007541f
C185 B.n151 VSUBS 0.005212f
C186 B.n152 VSUBS 0.007541f
C187 B.n153 VSUBS 0.007541f
C188 B.n154 VSUBS 0.007541f
C189 B.n155 VSUBS 0.007541f
C190 B.n156 VSUBS 0.007541f
C191 B.t10 VSUBS 0.277071f
C192 B.t11 VSUBS 0.314547f
C193 B.t9 VSUBS 1.92714f
C194 B.n157 VSUBS 0.494709f
C195 B.n158 VSUBS 0.30195f
C196 B.n159 VSUBS 0.007541f
C197 B.n160 VSUBS 0.007541f
C198 B.n161 VSUBS 0.007541f
C199 B.n162 VSUBS 0.007541f
C200 B.n163 VSUBS 0.007541f
C201 B.n164 VSUBS 0.007541f
C202 B.n165 VSUBS 0.007541f
C203 B.n166 VSUBS 0.007541f
C204 B.n167 VSUBS 0.007541f
C205 B.n168 VSUBS 0.007541f
C206 B.n169 VSUBS 0.007541f
C207 B.n170 VSUBS 0.007541f
C208 B.n171 VSUBS 0.007541f
C209 B.n172 VSUBS 0.007541f
C210 B.n173 VSUBS 0.007541f
C211 B.n174 VSUBS 0.007541f
C212 B.n175 VSUBS 0.007541f
C213 B.n176 VSUBS 0.007541f
C214 B.n177 VSUBS 0.007541f
C215 B.n178 VSUBS 0.007541f
C216 B.n179 VSUBS 0.007541f
C217 B.n180 VSUBS 0.007541f
C218 B.n181 VSUBS 0.007541f
C219 B.n182 VSUBS 0.016867f
C220 B.n183 VSUBS 0.007541f
C221 B.n184 VSUBS 0.007541f
C222 B.n185 VSUBS 0.007541f
C223 B.n186 VSUBS 0.007541f
C224 B.n187 VSUBS 0.007541f
C225 B.n188 VSUBS 0.007541f
C226 B.n189 VSUBS 0.007541f
C227 B.n190 VSUBS 0.007541f
C228 B.n191 VSUBS 0.007541f
C229 B.n192 VSUBS 0.007541f
C230 B.n193 VSUBS 0.007541f
C231 B.n194 VSUBS 0.007541f
C232 B.n195 VSUBS 0.007541f
C233 B.n196 VSUBS 0.007541f
C234 B.n197 VSUBS 0.007541f
C235 B.n198 VSUBS 0.007541f
C236 B.n199 VSUBS 0.007541f
C237 B.n200 VSUBS 0.007541f
C238 B.n201 VSUBS 0.007541f
C239 B.n202 VSUBS 0.007541f
C240 B.n203 VSUBS 0.007541f
C241 B.n204 VSUBS 0.007541f
C242 B.n205 VSUBS 0.007541f
C243 B.n206 VSUBS 0.007541f
C244 B.n207 VSUBS 0.007541f
C245 B.n208 VSUBS 0.007541f
C246 B.n209 VSUBS 0.007541f
C247 B.n210 VSUBS 0.007541f
C248 B.n211 VSUBS 0.007541f
C249 B.n212 VSUBS 0.007541f
C250 B.n213 VSUBS 0.007541f
C251 B.n214 VSUBS 0.007541f
C252 B.n215 VSUBS 0.007541f
C253 B.n216 VSUBS 0.007541f
C254 B.n217 VSUBS 0.007541f
C255 B.n218 VSUBS 0.007541f
C256 B.n219 VSUBS 0.007541f
C257 B.n220 VSUBS 0.007541f
C258 B.n221 VSUBS 0.007541f
C259 B.n222 VSUBS 0.007541f
C260 B.n223 VSUBS 0.007541f
C261 B.n224 VSUBS 0.007541f
C262 B.n225 VSUBS 0.007541f
C263 B.n226 VSUBS 0.007541f
C264 B.n227 VSUBS 0.007541f
C265 B.n228 VSUBS 0.007541f
C266 B.n229 VSUBS 0.007541f
C267 B.n230 VSUBS 0.007541f
C268 B.n231 VSUBS 0.007541f
C269 B.n232 VSUBS 0.007541f
C270 B.n233 VSUBS 0.007541f
C271 B.n234 VSUBS 0.007541f
C272 B.n235 VSUBS 0.007541f
C273 B.n236 VSUBS 0.007541f
C274 B.n237 VSUBS 0.007541f
C275 B.n238 VSUBS 0.007541f
C276 B.n239 VSUBS 0.007541f
C277 B.n240 VSUBS 0.007541f
C278 B.n241 VSUBS 0.007541f
C279 B.n242 VSUBS 0.007541f
C280 B.n243 VSUBS 0.007541f
C281 B.n244 VSUBS 0.007541f
C282 B.n245 VSUBS 0.007541f
C283 B.n246 VSUBS 0.007541f
C284 B.n247 VSUBS 0.007541f
C285 B.n248 VSUBS 0.007541f
C286 B.n249 VSUBS 0.007541f
C287 B.n250 VSUBS 0.007541f
C288 B.n251 VSUBS 0.007541f
C289 B.n252 VSUBS 0.007541f
C290 B.n253 VSUBS 0.007541f
C291 B.n254 VSUBS 0.007541f
C292 B.n255 VSUBS 0.007541f
C293 B.n256 VSUBS 0.007541f
C294 B.n257 VSUBS 0.007541f
C295 B.n258 VSUBS 0.007541f
C296 B.n259 VSUBS 0.007541f
C297 B.n260 VSUBS 0.007541f
C298 B.n261 VSUBS 0.007541f
C299 B.n262 VSUBS 0.007541f
C300 B.n263 VSUBS 0.007541f
C301 B.n264 VSUBS 0.007541f
C302 B.n265 VSUBS 0.007541f
C303 B.n266 VSUBS 0.007541f
C304 B.n267 VSUBS 0.007541f
C305 B.n268 VSUBS 0.007541f
C306 B.n269 VSUBS 0.016867f
C307 B.n270 VSUBS 0.017954f
C308 B.n271 VSUBS 0.017954f
C309 B.n272 VSUBS 0.007541f
C310 B.n273 VSUBS 0.007541f
C311 B.n274 VSUBS 0.007541f
C312 B.n275 VSUBS 0.007541f
C313 B.n276 VSUBS 0.007541f
C314 B.n277 VSUBS 0.007541f
C315 B.n278 VSUBS 0.007541f
C316 B.n279 VSUBS 0.007541f
C317 B.n280 VSUBS 0.007541f
C318 B.n281 VSUBS 0.007541f
C319 B.n282 VSUBS 0.007541f
C320 B.n283 VSUBS 0.007541f
C321 B.n284 VSUBS 0.007541f
C322 B.n285 VSUBS 0.007541f
C323 B.n286 VSUBS 0.007541f
C324 B.n287 VSUBS 0.007541f
C325 B.n288 VSUBS 0.007541f
C326 B.n289 VSUBS 0.007541f
C327 B.n290 VSUBS 0.007541f
C328 B.n291 VSUBS 0.007541f
C329 B.n292 VSUBS 0.007541f
C330 B.n293 VSUBS 0.007541f
C331 B.n294 VSUBS 0.007541f
C332 B.n295 VSUBS 0.007541f
C333 B.n296 VSUBS 0.007541f
C334 B.n297 VSUBS 0.007541f
C335 B.n298 VSUBS 0.007541f
C336 B.n299 VSUBS 0.007541f
C337 B.n300 VSUBS 0.007541f
C338 B.n301 VSUBS 0.007541f
C339 B.n302 VSUBS 0.007541f
C340 B.n303 VSUBS 0.007541f
C341 B.n304 VSUBS 0.007541f
C342 B.n305 VSUBS 0.007541f
C343 B.n306 VSUBS 0.007541f
C344 B.n307 VSUBS 0.007541f
C345 B.n308 VSUBS 0.007541f
C346 B.n309 VSUBS 0.007541f
C347 B.n310 VSUBS 0.007541f
C348 B.n311 VSUBS 0.007541f
C349 B.n312 VSUBS 0.007541f
C350 B.n313 VSUBS 0.007541f
C351 B.n314 VSUBS 0.007541f
C352 B.n315 VSUBS 0.007541f
C353 B.n316 VSUBS 0.007541f
C354 B.n317 VSUBS 0.007541f
C355 B.n318 VSUBS 0.007541f
C356 B.n319 VSUBS 0.007541f
C357 B.n320 VSUBS 0.007541f
C358 B.n321 VSUBS 0.007541f
C359 B.n322 VSUBS 0.007541f
C360 B.n323 VSUBS 0.007541f
C361 B.n324 VSUBS 0.007541f
C362 B.n325 VSUBS 0.007541f
C363 B.n326 VSUBS 0.007541f
C364 B.n327 VSUBS 0.007541f
C365 B.n328 VSUBS 0.007541f
C366 B.n329 VSUBS 0.007541f
C367 B.n330 VSUBS 0.007541f
C368 B.n331 VSUBS 0.007541f
C369 B.n332 VSUBS 0.007541f
C370 B.n333 VSUBS 0.007541f
C371 B.n334 VSUBS 0.007541f
C372 B.n335 VSUBS 0.007541f
C373 B.n336 VSUBS 0.007541f
C374 B.n337 VSUBS 0.007541f
C375 B.n338 VSUBS 0.007541f
C376 B.n339 VSUBS 0.007541f
C377 B.n340 VSUBS 0.007541f
C378 B.n341 VSUBS 0.005212f
C379 B.n342 VSUBS 0.017472f
C380 B.n343 VSUBS 0.006099f
C381 B.n344 VSUBS 0.007541f
C382 B.n345 VSUBS 0.007541f
C383 B.n346 VSUBS 0.007541f
C384 B.n347 VSUBS 0.007541f
C385 B.n348 VSUBS 0.007541f
C386 B.n349 VSUBS 0.007541f
C387 B.n350 VSUBS 0.007541f
C388 B.n351 VSUBS 0.007541f
C389 B.n352 VSUBS 0.007541f
C390 B.n353 VSUBS 0.007541f
C391 B.n354 VSUBS 0.007541f
C392 B.t7 VSUBS 0.277074f
C393 B.t8 VSUBS 0.314551f
C394 B.t6 VSUBS 1.92714f
C395 B.n355 VSUBS 0.494706f
C396 B.n356 VSUBS 0.301947f
C397 B.n357 VSUBS 0.017472f
C398 B.n358 VSUBS 0.006099f
C399 B.n359 VSUBS 0.007541f
C400 B.n360 VSUBS 0.007541f
C401 B.n361 VSUBS 0.007541f
C402 B.n362 VSUBS 0.007541f
C403 B.n363 VSUBS 0.007541f
C404 B.n364 VSUBS 0.007541f
C405 B.n365 VSUBS 0.007541f
C406 B.n366 VSUBS 0.007541f
C407 B.n367 VSUBS 0.007541f
C408 B.n368 VSUBS 0.007541f
C409 B.n369 VSUBS 0.007541f
C410 B.n370 VSUBS 0.007541f
C411 B.n371 VSUBS 0.007541f
C412 B.n372 VSUBS 0.007541f
C413 B.n373 VSUBS 0.007541f
C414 B.n374 VSUBS 0.007541f
C415 B.n375 VSUBS 0.007541f
C416 B.n376 VSUBS 0.007541f
C417 B.n377 VSUBS 0.007541f
C418 B.n378 VSUBS 0.007541f
C419 B.n379 VSUBS 0.007541f
C420 B.n380 VSUBS 0.007541f
C421 B.n381 VSUBS 0.007541f
C422 B.n382 VSUBS 0.007541f
C423 B.n383 VSUBS 0.007541f
C424 B.n384 VSUBS 0.007541f
C425 B.n385 VSUBS 0.007541f
C426 B.n386 VSUBS 0.007541f
C427 B.n387 VSUBS 0.007541f
C428 B.n388 VSUBS 0.007541f
C429 B.n389 VSUBS 0.007541f
C430 B.n390 VSUBS 0.007541f
C431 B.n391 VSUBS 0.007541f
C432 B.n392 VSUBS 0.007541f
C433 B.n393 VSUBS 0.007541f
C434 B.n394 VSUBS 0.007541f
C435 B.n395 VSUBS 0.007541f
C436 B.n396 VSUBS 0.007541f
C437 B.n397 VSUBS 0.007541f
C438 B.n398 VSUBS 0.007541f
C439 B.n399 VSUBS 0.007541f
C440 B.n400 VSUBS 0.007541f
C441 B.n401 VSUBS 0.007541f
C442 B.n402 VSUBS 0.007541f
C443 B.n403 VSUBS 0.007541f
C444 B.n404 VSUBS 0.007541f
C445 B.n405 VSUBS 0.007541f
C446 B.n406 VSUBS 0.007541f
C447 B.n407 VSUBS 0.007541f
C448 B.n408 VSUBS 0.007541f
C449 B.n409 VSUBS 0.007541f
C450 B.n410 VSUBS 0.007541f
C451 B.n411 VSUBS 0.007541f
C452 B.n412 VSUBS 0.007541f
C453 B.n413 VSUBS 0.007541f
C454 B.n414 VSUBS 0.007541f
C455 B.n415 VSUBS 0.007541f
C456 B.n416 VSUBS 0.007541f
C457 B.n417 VSUBS 0.007541f
C458 B.n418 VSUBS 0.007541f
C459 B.n419 VSUBS 0.007541f
C460 B.n420 VSUBS 0.007541f
C461 B.n421 VSUBS 0.007541f
C462 B.n422 VSUBS 0.007541f
C463 B.n423 VSUBS 0.007541f
C464 B.n424 VSUBS 0.007541f
C465 B.n425 VSUBS 0.007541f
C466 B.n426 VSUBS 0.007541f
C467 B.n427 VSUBS 0.007541f
C468 B.n428 VSUBS 0.007541f
C469 B.n429 VSUBS 0.007541f
C470 B.n430 VSUBS 0.017954f
C471 B.n431 VSUBS 0.017954f
C472 B.n432 VSUBS 0.016867f
C473 B.n433 VSUBS 0.007541f
C474 B.n434 VSUBS 0.007541f
C475 B.n435 VSUBS 0.007541f
C476 B.n436 VSUBS 0.007541f
C477 B.n437 VSUBS 0.007541f
C478 B.n438 VSUBS 0.007541f
C479 B.n439 VSUBS 0.007541f
C480 B.n440 VSUBS 0.007541f
C481 B.n441 VSUBS 0.007541f
C482 B.n442 VSUBS 0.007541f
C483 B.n443 VSUBS 0.007541f
C484 B.n444 VSUBS 0.007541f
C485 B.n445 VSUBS 0.007541f
C486 B.n446 VSUBS 0.007541f
C487 B.n447 VSUBS 0.007541f
C488 B.n448 VSUBS 0.007541f
C489 B.n449 VSUBS 0.007541f
C490 B.n450 VSUBS 0.007541f
C491 B.n451 VSUBS 0.007541f
C492 B.n452 VSUBS 0.007541f
C493 B.n453 VSUBS 0.007541f
C494 B.n454 VSUBS 0.007541f
C495 B.n455 VSUBS 0.007541f
C496 B.n456 VSUBS 0.007541f
C497 B.n457 VSUBS 0.007541f
C498 B.n458 VSUBS 0.007541f
C499 B.n459 VSUBS 0.007541f
C500 B.n460 VSUBS 0.007541f
C501 B.n461 VSUBS 0.007541f
C502 B.n462 VSUBS 0.007541f
C503 B.n463 VSUBS 0.007541f
C504 B.n464 VSUBS 0.007541f
C505 B.n465 VSUBS 0.007541f
C506 B.n466 VSUBS 0.007541f
C507 B.n467 VSUBS 0.007541f
C508 B.n468 VSUBS 0.007541f
C509 B.n469 VSUBS 0.007541f
C510 B.n470 VSUBS 0.007541f
C511 B.n471 VSUBS 0.007541f
C512 B.n472 VSUBS 0.007541f
C513 B.n473 VSUBS 0.007541f
C514 B.n474 VSUBS 0.007541f
C515 B.n475 VSUBS 0.007541f
C516 B.n476 VSUBS 0.007541f
C517 B.n477 VSUBS 0.007541f
C518 B.n478 VSUBS 0.007541f
C519 B.n479 VSUBS 0.007541f
C520 B.n480 VSUBS 0.007541f
C521 B.n481 VSUBS 0.007541f
C522 B.n482 VSUBS 0.007541f
C523 B.n483 VSUBS 0.007541f
C524 B.n484 VSUBS 0.007541f
C525 B.n485 VSUBS 0.007541f
C526 B.n486 VSUBS 0.007541f
C527 B.n487 VSUBS 0.007541f
C528 B.n488 VSUBS 0.007541f
C529 B.n489 VSUBS 0.007541f
C530 B.n490 VSUBS 0.007541f
C531 B.n491 VSUBS 0.007541f
C532 B.n492 VSUBS 0.007541f
C533 B.n493 VSUBS 0.007541f
C534 B.n494 VSUBS 0.007541f
C535 B.n495 VSUBS 0.007541f
C536 B.n496 VSUBS 0.007541f
C537 B.n497 VSUBS 0.007541f
C538 B.n498 VSUBS 0.007541f
C539 B.n499 VSUBS 0.007541f
C540 B.n500 VSUBS 0.007541f
C541 B.n501 VSUBS 0.007541f
C542 B.n502 VSUBS 0.007541f
C543 B.n503 VSUBS 0.007541f
C544 B.n504 VSUBS 0.007541f
C545 B.n505 VSUBS 0.007541f
C546 B.n506 VSUBS 0.007541f
C547 B.n507 VSUBS 0.007541f
C548 B.n508 VSUBS 0.007541f
C549 B.n509 VSUBS 0.007541f
C550 B.n510 VSUBS 0.007541f
C551 B.n511 VSUBS 0.007541f
C552 B.n512 VSUBS 0.007541f
C553 B.n513 VSUBS 0.007541f
C554 B.n514 VSUBS 0.007541f
C555 B.n515 VSUBS 0.007541f
C556 B.n516 VSUBS 0.007541f
C557 B.n517 VSUBS 0.007541f
C558 B.n518 VSUBS 0.007541f
C559 B.n519 VSUBS 0.007541f
C560 B.n520 VSUBS 0.007541f
C561 B.n521 VSUBS 0.007541f
C562 B.n522 VSUBS 0.007541f
C563 B.n523 VSUBS 0.007541f
C564 B.n524 VSUBS 0.007541f
C565 B.n525 VSUBS 0.007541f
C566 B.n526 VSUBS 0.007541f
C567 B.n527 VSUBS 0.007541f
C568 B.n528 VSUBS 0.007541f
C569 B.n529 VSUBS 0.007541f
C570 B.n530 VSUBS 0.007541f
C571 B.n531 VSUBS 0.007541f
C572 B.n532 VSUBS 0.007541f
C573 B.n533 VSUBS 0.007541f
C574 B.n534 VSUBS 0.007541f
C575 B.n535 VSUBS 0.007541f
C576 B.n536 VSUBS 0.007541f
C577 B.n537 VSUBS 0.007541f
C578 B.n538 VSUBS 0.007541f
C579 B.n539 VSUBS 0.007541f
C580 B.n540 VSUBS 0.007541f
C581 B.n541 VSUBS 0.007541f
C582 B.n542 VSUBS 0.007541f
C583 B.n543 VSUBS 0.007541f
C584 B.n544 VSUBS 0.007541f
C585 B.n545 VSUBS 0.007541f
C586 B.n546 VSUBS 0.007541f
C587 B.n547 VSUBS 0.007541f
C588 B.n548 VSUBS 0.007541f
C589 B.n549 VSUBS 0.007541f
C590 B.n550 VSUBS 0.007541f
C591 B.n551 VSUBS 0.007541f
C592 B.n552 VSUBS 0.007541f
C593 B.n553 VSUBS 0.007541f
C594 B.n554 VSUBS 0.007541f
C595 B.n555 VSUBS 0.007541f
C596 B.n556 VSUBS 0.007541f
C597 B.n557 VSUBS 0.007541f
C598 B.n558 VSUBS 0.007541f
C599 B.n559 VSUBS 0.007541f
C600 B.n560 VSUBS 0.007541f
C601 B.n561 VSUBS 0.007541f
C602 B.n562 VSUBS 0.007541f
C603 B.n563 VSUBS 0.007541f
C604 B.n564 VSUBS 0.007541f
C605 B.n565 VSUBS 0.007541f
C606 B.n566 VSUBS 0.007541f
C607 B.n567 VSUBS 0.017777f
C608 B.n568 VSUBS 0.017045f
C609 B.n569 VSUBS 0.017954f
C610 B.n570 VSUBS 0.007541f
C611 B.n571 VSUBS 0.007541f
C612 B.n572 VSUBS 0.007541f
C613 B.n573 VSUBS 0.007541f
C614 B.n574 VSUBS 0.007541f
C615 B.n575 VSUBS 0.007541f
C616 B.n576 VSUBS 0.007541f
C617 B.n577 VSUBS 0.007541f
C618 B.n578 VSUBS 0.007541f
C619 B.n579 VSUBS 0.007541f
C620 B.n580 VSUBS 0.007541f
C621 B.n581 VSUBS 0.007541f
C622 B.n582 VSUBS 0.007541f
C623 B.n583 VSUBS 0.007541f
C624 B.n584 VSUBS 0.007541f
C625 B.n585 VSUBS 0.007541f
C626 B.n586 VSUBS 0.007541f
C627 B.n587 VSUBS 0.007541f
C628 B.n588 VSUBS 0.007541f
C629 B.n589 VSUBS 0.007541f
C630 B.n590 VSUBS 0.007541f
C631 B.n591 VSUBS 0.007541f
C632 B.n592 VSUBS 0.007541f
C633 B.n593 VSUBS 0.007541f
C634 B.n594 VSUBS 0.007541f
C635 B.n595 VSUBS 0.007541f
C636 B.n596 VSUBS 0.007541f
C637 B.n597 VSUBS 0.007541f
C638 B.n598 VSUBS 0.007541f
C639 B.n599 VSUBS 0.007541f
C640 B.n600 VSUBS 0.007541f
C641 B.n601 VSUBS 0.007541f
C642 B.n602 VSUBS 0.007541f
C643 B.n603 VSUBS 0.007541f
C644 B.n604 VSUBS 0.007541f
C645 B.n605 VSUBS 0.007541f
C646 B.n606 VSUBS 0.007541f
C647 B.n607 VSUBS 0.007541f
C648 B.n608 VSUBS 0.007541f
C649 B.n609 VSUBS 0.007541f
C650 B.n610 VSUBS 0.007541f
C651 B.n611 VSUBS 0.007541f
C652 B.n612 VSUBS 0.007541f
C653 B.n613 VSUBS 0.007541f
C654 B.n614 VSUBS 0.007541f
C655 B.n615 VSUBS 0.007541f
C656 B.n616 VSUBS 0.007541f
C657 B.n617 VSUBS 0.007541f
C658 B.n618 VSUBS 0.007541f
C659 B.n619 VSUBS 0.007541f
C660 B.n620 VSUBS 0.007541f
C661 B.n621 VSUBS 0.007541f
C662 B.n622 VSUBS 0.007541f
C663 B.n623 VSUBS 0.007541f
C664 B.n624 VSUBS 0.007541f
C665 B.n625 VSUBS 0.007541f
C666 B.n626 VSUBS 0.007541f
C667 B.n627 VSUBS 0.007541f
C668 B.n628 VSUBS 0.007541f
C669 B.n629 VSUBS 0.007541f
C670 B.n630 VSUBS 0.007541f
C671 B.n631 VSUBS 0.007541f
C672 B.n632 VSUBS 0.007541f
C673 B.n633 VSUBS 0.007541f
C674 B.n634 VSUBS 0.007541f
C675 B.n635 VSUBS 0.007541f
C676 B.n636 VSUBS 0.007541f
C677 B.n637 VSUBS 0.007541f
C678 B.n638 VSUBS 0.007541f
C679 B.n639 VSUBS 0.005212f
C680 B.n640 VSUBS 0.017472f
C681 B.n641 VSUBS 0.006099f
C682 B.n642 VSUBS 0.007541f
C683 B.n643 VSUBS 0.007541f
C684 B.n644 VSUBS 0.007541f
C685 B.n645 VSUBS 0.007541f
C686 B.n646 VSUBS 0.007541f
C687 B.n647 VSUBS 0.007541f
C688 B.n648 VSUBS 0.007541f
C689 B.n649 VSUBS 0.007541f
C690 B.n650 VSUBS 0.007541f
C691 B.n651 VSUBS 0.007541f
C692 B.n652 VSUBS 0.007541f
C693 B.n653 VSUBS 0.006099f
C694 B.n654 VSUBS 0.007541f
C695 B.n655 VSUBS 0.007541f
C696 B.n656 VSUBS 0.007541f
C697 B.n657 VSUBS 0.007541f
C698 B.n658 VSUBS 0.007541f
C699 B.n659 VSUBS 0.007541f
C700 B.n660 VSUBS 0.007541f
C701 B.n661 VSUBS 0.007541f
C702 B.n662 VSUBS 0.007541f
C703 B.n663 VSUBS 0.007541f
C704 B.n664 VSUBS 0.007541f
C705 B.n665 VSUBS 0.007541f
C706 B.n666 VSUBS 0.007541f
C707 B.n667 VSUBS 0.007541f
C708 B.n668 VSUBS 0.007541f
C709 B.n669 VSUBS 0.007541f
C710 B.n670 VSUBS 0.007541f
C711 B.n671 VSUBS 0.007541f
C712 B.n672 VSUBS 0.007541f
C713 B.n673 VSUBS 0.007541f
C714 B.n674 VSUBS 0.007541f
C715 B.n675 VSUBS 0.007541f
C716 B.n676 VSUBS 0.007541f
C717 B.n677 VSUBS 0.007541f
C718 B.n678 VSUBS 0.007541f
C719 B.n679 VSUBS 0.007541f
C720 B.n680 VSUBS 0.007541f
C721 B.n681 VSUBS 0.007541f
C722 B.n682 VSUBS 0.007541f
C723 B.n683 VSUBS 0.007541f
C724 B.n684 VSUBS 0.007541f
C725 B.n685 VSUBS 0.007541f
C726 B.n686 VSUBS 0.007541f
C727 B.n687 VSUBS 0.007541f
C728 B.n688 VSUBS 0.007541f
C729 B.n689 VSUBS 0.007541f
C730 B.n690 VSUBS 0.007541f
C731 B.n691 VSUBS 0.007541f
C732 B.n692 VSUBS 0.007541f
C733 B.n693 VSUBS 0.007541f
C734 B.n694 VSUBS 0.007541f
C735 B.n695 VSUBS 0.007541f
C736 B.n696 VSUBS 0.007541f
C737 B.n697 VSUBS 0.007541f
C738 B.n698 VSUBS 0.007541f
C739 B.n699 VSUBS 0.007541f
C740 B.n700 VSUBS 0.007541f
C741 B.n701 VSUBS 0.007541f
C742 B.n702 VSUBS 0.007541f
C743 B.n703 VSUBS 0.007541f
C744 B.n704 VSUBS 0.007541f
C745 B.n705 VSUBS 0.007541f
C746 B.n706 VSUBS 0.007541f
C747 B.n707 VSUBS 0.007541f
C748 B.n708 VSUBS 0.007541f
C749 B.n709 VSUBS 0.007541f
C750 B.n710 VSUBS 0.007541f
C751 B.n711 VSUBS 0.007541f
C752 B.n712 VSUBS 0.007541f
C753 B.n713 VSUBS 0.007541f
C754 B.n714 VSUBS 0.007541f
C755 B.n715 VSUBS 0.007541f
C756 B.n716 VSUBS 0.007541f
C757 B.n717 VSUBS 0.007541f
C758 B.n718 VSUBS 0.007541f
C759 B.n719 VSUBS 0.007541f
C760 B.n720 VSUBS 0.007541f
C761 B.n721 VSUBS 0.007541f
C762 B.n722 VSUBS 0.007541f
C763 B.n723 VSUBS 0.007541f
C764 B.n724 VSUBS 0.007541f
C765 B.n725 VSUBS 0.017954f
C766 B.n726 VSUBS 0.017954f
C767 B.n727 VSUBS 0.016867f
C768 B.n728 VSUBS 0.007541f
C769 B.n729 VSUBS 0.007541f
C770 B.n730 VSUBS 0.007541f
C771 B.n731 VSUBS 0.007541f
C772 B.n732 VSUBS 0.007541f
C773 B.n733 VSUBS 0.007541f
C774 B.n734 VSUBS 0.007541f
C775 B.n735 VSUBS 0.007541f
C776 B.n736 VSUBS 0.007541f
C777 B.n737 VSUBS 0.007541f
C778 B.n738 VSUBS 0.007541f
C779 B.n739 VSUBS 0.007541f
C780 B.n740 VSUBS 0.007541f
C781 B.n741 VSUBS 0.007541f
C782 B.n742 VSUBS 0.007541f
C783 B.n743 VSUBS 0.007541f
C784 B.n744 VSUBS 0.007541f
C785 B.n745 VSUBS 0.007541f
C786 B.n746 VSUBS 0.007541f
C787 B.n747 VSUBS 0.007541f
C788 B.n748 VSUBS 0.007541f
C789 B.n749 VSUBS 0.007541f
C790 B.n750 VSUBS 0.007541f
C791 B.n751 VSUBS 0.007541f
C792 B.n752 VSUBS 0.007541f
C793 B.n753 VSUBS 0.007541f
C794 B.n754 VSUBS 0.007541f
C795 B.n755 VSUBS 0.007541f
C796 B.n756 VSUBS 0.007541f
C797 B.n757 VSUBS 0.007541f
C798 B.n758 VSUBS 0.007541f
C799 B.n759 VSUBS 0.007541f
C800 B.n760 VSUBS 0.007541f
C801 B.n761 VSUBS 0.007541f
C802 B.n762 VSUBS 0.007541f
C803 B.n763 VSUBS 0.007541f
C804 B.n764 VSUBS 0.007541f
C805 B.n765 VSUBS 0.007541f
C806 B.n766 VSUBS 0.007541f
C807 B.n767 VSUBS 0.007541f
C808 B.n768 VSUBS 0.007541f
C809 B.n769 VSUBS 0.007541f
C810 B.n770 VSUBS 0.007541f
C811 B.n771 VSUBS 0.007541f
C812 B.n772 VSUBS 0.007541f
C813 B.n773 VSUBS 0.007541f
C814 B.n774 VSUBS 0.007541f
C815 B.n775 VSUBS 0.007541f
C816 B.n776 VSUBS 0.007541f
C817 B.n777 VSUBS 0.007541f
C818 B.n778 VSUBS 0.007541f
C819 B.n779 VSUBS 0.007541f
C820 B.n780 VSUBS 0.007541f
C821 B.n781 VSUBS 0.007541f
C822 B.n782 VSUBS 0.007541f
C823 B.n783 VSUBS 0.007541f
C824 B.n784 VSUBS 0.007541f
C825 B.n785 VSUBS 0.007541f
C826 B.n786 VSUBS 0.007541f
C827 B.n787 VSUBS 0.007541f
C828 B.n788 VSUBS 0.007541f
C829 B.n789 VSUBS 0.007541f
C830 B.n790 VSUBS 0.007541f
C831 B.n791 VSUBS 0.007541f
C832 B.n792 VSUBS 0.007541f
C833 B.n793 VSUBS 0.007541f
C834 B.n794 VSUBS 0.007541f
C835 B.n795 VSUBS 0.017075f
C836 VDD2.n0 VSUBS 0.028886f
C837 VDD2.n1 VSUBS 0.027675f
C838 VDD2.n2 VSUBS 0.015309f
C839 VDD2.n3 VSUBS 0.035151f
C840 VDD2.n4 VSUBS 0.015746f
C841 VDD2.n5 VSUBS 0.027675f
C842 VDD2.n6 VSUBS 0.014871f
C843 VDD2.n7 VSUBS 0.035151f
C844 VDD2.n8 VSUBS 0.015746f
C845 VDD2.n9 VSUBS 0.027675f
C846 VDD2.n10 VSUBS 0.014871f
C847 VDD2.n11 VSUBS 0.035151f
C848 VDD2.n12 VSUBS 0.015746f
C849 VDD2.n13 VSUBS 0.027675f
C850 VDD2.n14 VSUBS 0.014871f
C851 VDD2.n15 VSUBS 0.035151f
C852 VDD2.n16 VSUBS 0.015746f
C853 VDD2.n17 VSUBS 0.027675f
C854 VDD2.n18 VSUBS 0.014871f
C855 VDD2.n19 VSUBS 0.035151f
C856 VDD2.n20 VSUBS 0.015746f
C857 VDD2.n21 VSUBS 0.027675f
C858 VDD2.n22 VSUBS 0.014871f
C859 VDD2.n23 VSUBS 0.026363f
C860 VDD2.n24 VSUBS 0.022361f
C861 VDD2.t4 VSUBS 0.075185f
C862 VDD2.n25 VSUBS 0.18725f
C863 VDD2.n26 VSUBS 1.6465f
C864 VDD2.n27 VSUBS 0.014871f
C865 VDD2.n28 VSUBS 0.015746f
C866 VDD2.n29 VSUBS 0.035151f
C867 VDD2.n30 VSUBS 0.035151f
C868 VDD2.n31 VSUBS 0.015746f
C869 VDD2.n32 VSUBS 0.014871f
C870 VDD2.n33 VSUBS 0.027675f
C871 VDD2.n34 VSUBS 0.027675f
C872 VDD2.n35 VSUBS 0.014871f
C873 VDD2.n36 VSUBS 0.015746f
C874 VDD2.n37 VSUBS 0.035151f
C875 VDD2.n38 VSUBS 0.035151f
C876 VDD2.n39 VSUBS 0.015746f
C877 VDD2.n40 VSUBS 0.014871f
C878 VDD2.n41 VSUBS 0.027675f
C879 VDD2.n42 VSUBS 0.027675f
C880 VDD2.n43 VSUBS 0.014871f
C881 VDD2.n44 VSUBS 0.015746f
C882 VDD2.n45 VSUBS 0.035151f
C883 VDD2.n46 VSUBS 0.035151f
C884 VDD2.n47 VSUBS 0.015746f
C885 VDD2.n48 VSUBS 0.014871f
C886 VDD2.n49 VSUBS 0.027675f
C887 VDD2.n50 VSUBS 0.027675f
C888 VDD2.n51 VSUBS 0.014871f
C889 VDD2.n52 VSUBS 0.015746f
C890 VDD2.n53 VSUBS 0.035151f
C891 VDD2.n54 VSUBS 0.035151f
C892 VDD2.n55 VSUBS 0.015746f
C893 VDD2.n56 VSUBS 0.014871f
C894 VDD2.n57 VSUBS 0.027675f
C895 VDD2.n58 VSUBS 0.027675f
C896 VDD2.n59 VSUBS 0.014871f
C897 VDD2.n60 VSUBS 0.015746f
C898 VDD2.n61 VSUBS 0.035151f
C899 VDD2.n62 VSUBS 0.035151f
C900 VDD2.n63 VSUBS 0.015746f
C901 VDD2.n64 VSUBS 0.014871f
C902 VDD2.n65 VSUBS 0.027675f
C903 VDD2.n66 VSUBS 0.027675f
C904 VDD2.n67 VSUBS 0.014871f
C905 VDD2.n68 VSUBS 0.014871f
C906 VDD2.n69 VSUBS 0.015746f
C907 VDD2.n70 VSUBS 0.035151f
C908 VDD2.n71 VSUBS 0.035151f
C909 VDD2.n72 VSUBS 0.079906f
C910 VDD2.n73 VSUBS 0.015309f
C911 VDD2.n74 VSUBS 0.014871f
C912 VDD2.n75 VSUBS 0.068507f
C913 VDD2.n76 VSUBS 0.067794f
C914 VDD2.t1 VSUBS 0.307051f
C915 VDD2.t5 VSUBS 0.307051f
C916 VDD2.n77 VSUBS 2.48417f
C917 VDD2.n78 VSUBS 3.49331f
C918 VDD2.n79 VSUBS 0.028886f
C919 VDD2.n80 VSUBS 0.027675f
C920 VDD2.n81 VSUBS 0.015309f
C921 VDD2.n82 VSUBS 0.035151f
C922 VDD2.n83 VSUBS 0.014871f
C923 VDD2.n84 VSUBS 0.015746f
C924 VDD2.n85 VSUBS 0.027675f
C925 VDD2.n86 VSUBS 0.014871f
C926 VDD2.n87 VSUBS 0.035151f
C927 VDD2.n88 VSUBS 0.015746f
C928 VDD2.n89 VSUBS 0.027675f
C929 VDD2.n90 VSUBS 0.014871f
C930 VDD2.n91 VSUBS 0.035151f
C931 VDD2.n92 VSUBS 0.015746f
C932 VDD2.n93 VSUBS 0.027675f
C933 VDD2.n94 VSUBS 0.014871f
C934 VDD2.n95 VSUBS 0.035151f
C935 VDD2.n96 VSUBS 0.015746f
C936 VDD2.n97 VSUBS 0.027675f
C937 VDD2.n98 VSUBS 0.014871f
C938 VDD2.n99 VSUBS 0.035151f
C939 VDD2.n100 VSUBS 0.015746f
C940 VDD2.n101 VSUBS 0.027675f
C941 VDD2.n102 VSUBS 0.014871f
C942 VDD2.n103 VSUBS 0.026363f
C943 VDD2.n104 VSUBS 0.022361f
C944 VDD2.t0 VSUBS 0.075185f
C945 VDD2.n105 VSUBS 0.18725f
C946 VDD2.n106 VSUBS 1.6465f
C947 VDD2.n107 VSUBS 0.014871f
C948 VDD2.n108 VSUBS 0.015746f
C949 VDD2.n109 VSUBS 0.035151f
C950 VDD2.n110 VSUBS 0.035151f
C951 VDD2.n111 VSUBS 0.015746f
C952 VDD2.n112 VSUBS 0.014871f
C953 VDD2.n113 VSUBS 0.027675f
C954 VDD2.n114 VSUBS 0.027675f
C955 VDD2.n115 VSUBS 0.014871f
C956 VDD2.n116 VSUBS 0.015746f
C957 VDD2.n117 VSUBS 0.035151f
C958 VDD2.n118 VSUBS 0.035151f
C959 VDD2.n119 VSUBS 0.015746f
C960 VDD2.n120 VSUBS 0.014871f
C961 VDD2.n121 VSUBS 0.027675f
C962 VDD2.n122 VSUBS 0.027675f
C963 VDD2.n123 VSUBS 0.014871f
C964 VDD2.n124 VSUBS 0.015746f
C965 VDD2.n125 VSUBS 0.035151f
C966 VDD2.n126 VSUBS 0.035151f
C967 VDD2.n127 VSUBS 0.015746f
C968 VDD2.n128 VSUBS 0.014871f
C969 VDD2.n129 VSUBS 0.027675f
C970 VDD2.n130 VSUBS 0.027675f
C971 VDD2.n131 VSUBS 0.014871f
C972 VDD2.n132 VSUBS 0.015746f
C973 VDD2.n133 VSUBS 0.035151f
C974 VDD2.n134 VSUBS 0.035151f
C975 VDD2.n135 VSUBS 0.015746f
C976 VDD2.n136 VSUBS 0.014871f
C977 VDD2.n137 VSUBS 0.027675f
C978 VDD2.n138 VSUBS 0.027675f
C979 VDD2.n139 VSUBS 0.014871f
C980 VDD2.n140 VSUBS 0.015746f
C981 VDD2.n141 VSUBS 0.035151f
C982 VDD2.n142 VSUBS 0.035151f
C983 VDD2.n143 VSUBS 0.015746f
C984 VDD2.n144 VSUBS 0.014871f
C985 VDD2.n145 VSUBS 0.027675f
C986 VDD2.n146 VSUBS 0.027675f
C987 VDD2.n147 VSUBS 0.014871f
C988 VDD2.n148 VSUBS 0.015746f
C989 VDD2.n149 VSUBS 0.035151f
C990 VDD2.n150 VSUBS 0.035151f
C991 VDD2.n151 VSUBS 0.079906f
C992 VDD2.n152 VSUBS 0.015309f
C993 VDD2.n153 VSUBS 0.014871f
C994 VDD2.n154 VSUBS 0.068507f
C995 VDD2.n155 VSUBS 0.059165f
C996 VDD2.n156 VSUBS 3.07511f
C997 VDD2.t2 VSUBS 0.307051f
C998 VDD2.t3 VSUBS 0.307051f
C999 VDD2.n157 VSUBS 2.48413f
C1000 VN.n0 VSUBS 0.036765f
C1001 VN.t0 VSUBS 3.01018f
C1002 VN.n1 VSUBS 0.052452f
C1003 VN.n2 VSUBS 0.027888f
C1004 VN.t4 VSUBS 3.01018f
C1005 VN.n3 VSUBS 1.15262f
C1006 VN.t1 VSUBS 3.28794f
C1007 VN.n4 VSUBS 1.09463f
C1008 VN.n5 VSUBS 0.29282f
C1009 VN.n6 VSUBS 0.051715f
C1010 VN.n7 VSUBS 0.056026f
C1011 VN.n8 VSUBS 0.024316f
C1012 VN.n9 VSUBS 0.027888f
C1013 VN.n10 VSUBS 0.027888f
C1014 VN.n11 VSUBS 0.027888f
C1015 VN.n12 VSUBS 0.051715f
C1016 VN.n13 VSUBS 0.033333f
C1017 VN.n14 VSUBS 1.14923f
C1018 VN.n15 VSUBS 0.049527f
C1019 VN.n16 VSUBS 0.036765f
C1020 VN.t5 VSUBS 3.01018f
C1021 VN.n17 VSUBS 0.052452f
C1022 VN.n18 VSUBS 0.027888f
C1023 VN.t3 VSUBS 3.01018f
C1024 VN.n19 VSUBS 1.15262f
C1025 VN.t2 VSUBS 3.28794f
C1026 VN.n20 VSUBS 1.09463f
C1027 VN.n21 VSUBS 0.29282f
C1028 VN.n22 VSUBS 0.051715f
C1029 VN.n23 VSUBS 0.056026f
C1030 VN.n24 VSUBS 0.024316f
C1031 VN.n25 VSUBS 0.027888f
C1032 VN.n26 VSUBS 0.027888f
C1033 VN.n27 VSUBS 0.027888f
C1034 VN.n28 VSUBS 0.051715f
C1035 VN.n29 VSUBS 0.033333f
C1036 VN.n30 VSUBS 1.14923f
C1037 VN.n31 VSUBS 1.62002f
C1038 VDD1.n0 VSUBS 0.028882f
C1039 VDD1.n1 VSUBS 0.027672f
C1040 VDD1.n2 VSUBS 0.015307f
C1041 VDD1.n3 VSUBS 0.035147f
C1042 VDD1.n4 VSUBS 0.01487f
C1043 VDD1.n5 VSUBS 0.015745f
C1044 VDD1.n6 VSUBS 0.027672f
C1045 VDD1.n7 VSUBS 0.01487f
C1046 VDD1.n8 VSUBS 0.035147f
C1047 VDD1.n9 VSUBS 0.015745f
C1048 VDD1.n10 VSUBS 0.027672f
C1049 VDD1.n11 VSUBS 0.01487f
C1050 VDD1.n12 VSUBS 0.035147f
C1051 VDD1.n13 VSUBS 0.015745f
C1052 VDD1.n14 VSUBS 0.027672f
C1053 VDD1.n15 VSUBS 0.01487f
C1054 VDD1.n16 VSUBS 0.035147f
C1055 VDD1.n17 VSUBS 0.015745f
C1056 VDD1.n18 VSUBS 0.027672f
C1057 VDD1.n19 VSUBS 0.01487f
C1058 VDD1.n20 VSUBS 0.035147f
C1059 VDD1.n21 VSUBS 0.015745f
C1060 VDD1.n22 VSUBS 0.027672f
C1061 VDD1.n23 VSUBS 0.01487f
C1062 VDD1.n24 VSUBS 0.02636f
C1063 VDD1.n25 VSUBS 0.022359f
C1064 VDD1.t1 VSUBS 0.075177f
C1065 VDD1.n26 VSUBS 0.18723f
C1066 VDD1.n27 VSUBS 1.64633f
C1067 VDD1.n28 VSUBS 0.01487f
C1068 VDD1.n29 VSUBS 0.015745f
C1069 VDD1.n30 VSUBS 0.035147f
C1070 VDD1.n31 VSUBS 0.035147f
C1071 VDD1.n32 VSUBS 0.015745f
C1072 VDD1.n33 VSUBS 0.01487f
C1073 VDD1.n34 VSUBS 0.027672f
C1074 VDD1.n35 VSUBS 0.027672f
C1075 VDD1.n36 VSUBS 0.01487f
C1076 VDD1.n37 VSUBS 0.015745f
C1077 VDD1.n38 VSUBS 0.035147f
C1078 VDD1.n39 VSUBS 0.035147f
C1079 VDD1.n40 VSUBS 0.015745f
C1080 VDD1.n41 VSUBS 0.01487f
C1081 VDD1.n42 VSUBS 0.027672f
C1082 VDD1.n43 VSUBS 0.027672f
C1083 VDD1.n44 VSUBS 0.01487f
C1084 VDD1.n45 VSUBS 0.015745f
C1085 VDD1.n46 VSUBS 0.035147f
C1086 VDD1.n47 VSUBS 0.035147f
C1087 VDD1.n48 VSUBS 0.015745f
C1088 VDD1.n49 VSUBS 0.01487f
C1089 VDD1.n50 VSUBS 0.027672f
C1090 VDD1.n51 VSUBS 0.027672f
C1091 VDD1.n52 VSUBS 0.01487f
C1092 VDD1.n53 VSUBS 0.015745f
C1093 VDD1.n54 VSUBS 0.035147f
C1094 VDD1.n55 VSUBS 0.035147f
C1095 VDD1.n56 VSUBS 0.015745f
C1096 VDD1.n57 VSUBS 0.01487f
C1097 VDD1.n58 VSUBS 0.027672f
C1098 VDD1.n59 VSUBS 0.027672f
C1099 VDD1.n60 VSUBS 0.01487f
C1100 VDD1.n61 VSUBS 0.015745f
C1101 VDD1.n62 VSUBS 0.035147f
C1102 VDD1.n63 VSUBS 0.035147f
C1103 VDD1.n64 VSUBS 0.015745f
C1104 VDD1.n65 VSUBS 0.01487f
C1105 VDD1.n66 VSUBS 0.027672f
C1106 VDD1.n67 VSUBS 0.027672f
C1107 VDD1.n68 VSUBS 0.01487f
C1108 VDD1.n69 VSUBS 0.015745f
C1109 VDD1.n70 VSUBS 0.035147f
C1110 VDD1.n71 VSUBS 0.035147f
C1111 VDD1.n72 VSUBS 0.079898f
C1112 VDD1.n73 VSUBS 0.015307f
C1113 VDD1.n74 VSUBS 0.01487f
C1114 VDD1.n75 VSUBS 0.068499f
C1115 VDD1.n76 VSUBS 0.068648f
C1116 VDD1.n77 VSUBS 0.028882f
C1117 VDD1.n78 VSUBS 0.027672f
C1118 VDD1.n79 VSUBS 0.015307f
C1119 VDD1.n80 VSUBS 0.035147f
C1120 VDD1.n81 VSUBS 0.015745f
C1121 VDD1.n82 VSUBS 0.027672f
C1122 VDD1.n83 VSUBS 0.01487f
C1123 VDD1.n84 VSUBS 0.035147f
C1124 VDD1.n85 VSUBS 0.015745f
C1125 VDD1.n86 VSUBS 0.027672f
C1126 VDD1.n87 VSUBS 0.01487f
C1127 VDD1.n88 VSUBS 0.035147f
C1128 VDD1.n89 VSUBS 0.015745f
C1129 VDD1.n90 VSUBS 0.027672f
C1130 VDD1.n91 VSUBS 0.01487f
C1131 VDD1.n92 VSUBS 0.035147f
C1132 VDD1.n93 VSUBS 0.015745f
C1133 VDD1.n94 VSUBS 0.027672f
C1134 VDD1.n95 VSUBS 0.01487f
C1135 VDD1.n96 VSUBS 0.035147f
C1136 VDD1.n97 VSUBS 0.015745f
C1137 VDD1.n98 VSUBS 0.027672f
C1138 VDD1.n99 VSUBS 0.01487f
C1139 VDD1.n100 VSUBS 0.02636f
C1140 VDD1.n101 VSUBS 0.022359f
C1141 VDD1.t0 VSUBS 0.075177f
C1142 VDD1.n102 VSUBS 0.18723f
C1143 VDD1.n103 VSUBS 1.64633f
C1144 VDD1.n104 VSUBS 0.01487f
C1145 VDD1.n105 VSUBS 0.015745f
C1146 VDD1.n106 VSUBS 0.035147f
C1147 VDD1.n107 VSUBS 0.035147f
C1148 VDD1.n108 VSUBS 0.015745f
C1149 VDD1.n109 VSUBS 0.01487f
C1150 VDD1.n110 VSUBS 0.027672f
C1151 VDD1.n111 VSUBS 0.027672f
C1152 VDD1.n112 VSUBS 0.01487f
C1153 VDD1.n113 VSUBS 0.015745f
C1154 VDD1.n114 VSUBS 0.035147f
C1155 VDD1.n115 VSUBS 0.035147f
C1156 VDD1.n116 VSUBS 0.015745f
C1157 VDD1.n117 VSUBS 0.01487f
C1158 VDD1.n118 VSUBS 0.027672f
C1159 VDD1.n119 VSUBS 0.027672f
C1160 VDD1.n120 VSUBS 0.01487f
C1161 VDD1.n121 VSUBS 0.015745f
C1162 VDD1.n122 VSUBS 0.035147f
C1163 VDD1.n123 VSUBS 0.035147f
C1164 VDD1.n124 VSUBS 0.015745f
C1165 VDD1.n125 VSUBS 0.01487f
C1166 VDD1.n126 VSUBS 0.027672f
C1167 VDD1.n127 VSUBS 0.027672f
C1168 VDD1.n128 VSUBS 0.01487f
C1169 VDD1.n129 VSUBS 0.015745f
C1170 VDD1.n130 VSUBS 0.035147f
C1171 VDD1.n131 VSUBS 0.035147f
C1172 VDD1.n132 VSUBS 0.015745f
C1173 VDD1.n133 VSUBS 0.01487f
C1174 VDD1.n134 VSUBS 0.027672f
C1175 VDD1.n135 VSUBS 0.027672f
C1176 VDD1.n136 VSUBS 0.01487f
C1177 VDD1.n137 VSUBS 0.015745f
C1178 VDD1.n138 VSUBS 0.035147f
C1179 VDD1.n139 VSUBS 0.035147f
C1180 VDD1.n140 VSUBS 0.015745f
C1181 VDD1.n141 VSUBS 0.01487f
C1182 VDD1.n142 VSUBS 0.027672f
C1183 VDD1.n143 VSUBS 0.027672f
C1184 VDD1.n144 VSUBS 0.01487f
C1185 VDD1.n145 VSUBS 0.01487f
C1186 VDD1.n146 VSUBS 0.015745f
C1187 VDD1.n147 VSUBS 0.035147f
C1188 VDD1.n148 VSUBS 0.035147f
C1189 VDD1.n149 VSUBS 0.079898f
C1190 VDD1.n150 VSUBS 0.015307f
C1191 VDD1.n151 VSUBS 0.01487f
C1192 VDD1.n152 VSUBS 0.068499f
C1193 VDD1.n153 VSUBS 0.067787f
C1194 VDD1.t3 VSUBS 0.307019f
C1195 VDD1.t4 VSUBS 0.307019f
C1196 VDD1.n154 VSUBS 2.48392f
C1197 VDD1.n155 VSUBS 3.63815f
C1198 VDD1.t2 VSUBS 0.307019f
C1199 VDD1.t5 VSUBS 0.307019f
C1200 VDD1.n156 VSUBS 2.47703f
C1201 VDD1.n157 VSUBS 3.61208f
C1202 VTAIL.t5 VSUBS 0.316487f
C1203 VTAIL.t4 VSUBS 0.316487f
C1204 VTAIL.n0 VSUBS 2.3997f
C1205 VTAIL.n1 VSUBS 0.880678f
C1206 VTAIL.n2 VSUBS 0.029773f
C1207 VTAIL.n3 VSUBS 0.028526f
C1208 VTAIL.n4 VSUBS 0.015779f
C1209 VTAIL.n5 VSUBS 0.036231f
C1210 VTAIL.n6 VSUBS 0.01623f
C1211 VTAIL.n7 VSUBS 0.028526f
C1212 VTAIL.n8 VSUBS 0.015328f
C1213 VTAIL.n9 VSUBS 0.036231f
C1214 VTAIL.n10 VSUBS 0.01623f
C1215 VTAIL.n11 VSUBS 0.028526f
C1216 VTAIL.n12 VSUBS 0.015328f
C1217 VTAIL.n13 VSUBS 0.036231f
C1218 VTAIL.n14 VSUBS 0.01623f
C1219 VTAIL.n15 VSUBS 0.028526f
C1220 VTAIL.n16 VSUBS 0.015328f
C1221 VTAIL.n17 VSUBS 0.036231f
C1222 VTAIL.n18 VSUBS 0.01623f
C1223 VTAIL.n19 VSUBS 0.028526f
C1224 VTAIL.n20 VSUBS 0.015328f
C1225 VTAIL.n21 VSUBS 0.036231f
C1226 VTAIL.n22 VSUBS 0.01623f
C1227 VTAIL.n23 VSUBS 0.028526f
C1228 VTAIL.n24 VSUBS 0.015328f
C1229 VTAIL.n25 VSUBS 0.027173f
C1230 VTAIL.n26 VSUBS 0.023048f
C1231 VTAIL.t8 VSUBS 0.077496f
C1232 VTAIL.n27 VSUBS 0.193004f
C1233 VTAIL.n28 VSUBS 1.6971f
C1234 VTAIL.n29 VSUBS 0.015328f
C1235 VTAIL.n30 VSUBS 0.01623f
C1236 VTAIL.n31 VSUBS 0.036231f
C1237 VTAIL.n32 VSUBS 0.036231f
C1238 VTAIL.n33 VSUBS 0.01623f
C1239 VTAIL.n34 VSUBS 0.015328f
C1240 VTAIL.n35 VSUBS 0.028526f
C1241 VTAIL.n36 VSUBS 0.028526f
C1242 VTAIL.n37 VSUBS 0.015328f
C1243 VTAIL.n38 VSUBS 0.01623f
C1244 VTAIL.n39 VSUBS 0.036231f
C1245 VTAIL.n40 VSUBS 0.036231f
C1246 VTAIL.n41 VSUBS 0.01623f
C1247 VTAIL.n42 VSUBS 0.015328f
C1248 VTAIL.n43 VSUBS 0.028526f
C1249 VTAIL.n44 VSUBS 0.028526f
C1250 VTAIL.n45 VSUBS 0.015328f
C1251 VTAIL.n46 VSUBS 0.01623f
C1252 VTAIL.n47 VSUBS 0.036231f
C1253 VTAIL.n48 VSUBS 0.036231f
C1254 VTAIL.n49 VSUBS 0.01623f
C1255 VTAIL.n50 VSUBS 0.015328f
C1256 VTAIL.n51 VSUBS 0.028526f
C1257 VTAIL.n52 VSUBS 0.028526f
C1258 VTAIL.n53 VSUBS 0.015328f
C1259 VTAIL.n54 VSUBS 0.01623f
C1260 VTAIL.n55 VSUBS 0.036231f
C1261 VTAIL.n56 VSUBS 0.036231f
C1262 VTAIL.n57 VSUBS 0.01623f
C1263 VTAIL.n58 VSUBS 0.015328f
C1264 VTAIL.n59 VSUBS 0.028526f
C1265 VTAIL.n60 VSUBS 0.028526f
C1266 VTAIL.n61 VSUBS 0.015328f
C1267 VTAIL.n62 VSUBS 0.01623f
C1268 VTAIL.n63 VSUBS 0.036231f
C1269 VTAIL.n64 VSUBS 0.036231f
C1270 VTAIL.n65 VSUBS 0.01623f
C1271 VTAIL.n66 VSUBS 0.015328f
C1272 VTAIL.n67 VSUBS 0.028526f
C1273 VTAIL.n68 VSUBS 0.028526f
C1274 VTAIL.n69 VSUBS 0.015328f
C1275 VTAIL.n70 VSUBS 0.015328f
C1276 VTAIL.n71 VSUBS 0.01623f
C1277 VTAIL.n72 VSUBS 0.036231f
C1278 VTAIL.n73 VSUBS 0.036231f
C1279 VTAIL.n74 VSUBS 0.082362f
C1280 VTAIL.n75 VSUBS 0.015779f
C1281 VTAIL.n76 VSUBS 0.015328f
C1282 VTAIL.n77 VSUBS 0.070612f
C1283 VTAIL.n78 VSUBS 0.041321f
C1284 VTAIL.n79 VSUBS 0.443402f
C1285 VTAIL.t9 VSUBS 0.316487f
C1286 VTAIL.t11 VSUBS 0.316487f
C1287 VTAIL.n80 VSUBS 2.3997f
C1288 VTAIL.n81 VSUBS 2.89195f
C1289 VTAIL.t0 VSUBS 0.316487f
C1290 VTAIL.t3 VSUBS 0.316487f
C1291 VTAIL.n82 VSUBS 2.39971f
C1292 VTAIL.n83 VSUBS 2.89193f
C1293 VTAIL.n84 VSUBS 0.029773f
C1294 VTAIL.n85 VSUBS 0.028526f
C1295 VTAIL.n86 VSUBS 0.015779f
C1296 VTAIL.n87 VSUBS 0.036231f
C1297 VTAIL.n88 VSUBS 0.015328f
C1298 VTAIL.n89 VSUBS 0.01623f
C1299 VTAIL.n90 VSUBS 0.028526f
C1300 VTAIL.n91 VSUBS 0.015328f
C1301 VTAIL.n92 VSUBS 0.036231f
C1302 VTAIL.n93 VSUBS 0.01623f
C1303 VTAIL.n94 VSUBS 0.028526f
C1304 VTAIL.n95 VSUBS 0.015328f
C1305 VTAIL.n96 VSUBS 0.036231f
C1306 VTAIL.n97 VSUBS 0.01623f
C1307 VTAIL.n98 VSUBS 0.028526f
C1308 VTAIL.n99 VSUBS 0.015328f
C1309 VTAIL.n100 VSUBS 0.036231f
C1310 VTAIL.n101 VSUBS 0.01623f
C1311 VTAIL.n102 VSUBS 0.028526f
C1312 VTAIL.n103 VSUBS 0.015328f
C1313 VTAIL.n104 VSUBS 0.036231f
C1314 VTAIL.n105 VSUBS 0.01623f
C1315 VTAIL.n106 VSUBS 0.028526f
C1316 VTAIL.n107 VSUBS 0.015328f
C1317 VTAIL.n108 VSUBS 0.027173f
C1318 VTAIL.n109 VSUBS 0.023048f
C1319 VTAIL.t2 VSUBS 0.077496f
C1320 VTAIL.n110 VSUBS 0.193004f
C1321 VTAIL.n111 VSUBS 1.6971f
C1322 VTAIL.n112 VSUBS 0.015328f
C1323 VTAIL.n113 VSUBS 0.01623f
C1324 VTAIL.n114 VSUBS 0.036231f
C1325 VTAIL.n115 VSUBS 0.036231f
C1326 VTAIL.n116 VSUBS 0.01623f
C1327 VTAIL.n117 VSUBS 0.015328f
C1328 VTAIL.n118 VSUBS 0.028526f
C1329 VTAIL.n119 VSUBS 0.028526f
C1330 VTAIL.n120 VSUBS 0.015328f
C1331 VTAIL.n121 VSUBS 0.01623f
C1332 VTAIL.n122 VSUBS 0.036231f
C1333 VTAIL.n123 VSUBS 0.036231f
C1334 VTAIL.n124 VSUBS 0.01623f
C1335 VTAIL.n125 VSUBS 0.015328f
C1336 VTAIL.n126 VSUBS 0.028526f
C1337 VTAIL.n127 VSUBS 0.028526f
C1338 VTAIL.n128 VSUBS 0.015328f
C1339 VTAIL.n129 VSUBS 0.01623f
C1340 VTAIL.n130 VSUBS 0.036231f
C1341 VTAIL.n131 VSUBS 0.036231f
C1342 VTAIL.n132 VSUBS 0.01623f
C1343 VTAIL.n133 VSUBS 0.015328f
C1344 VTAIL.n134 VSUBS 0.028526f
C1345 VTAIL.n135 VSUBS 0.028526f
C1346 VTAIL.n136 VSUBS 0.015328f
C1347 VTAIL.n137 VSUBS 0.01623f
C1348 VTAIL.n138 VSUBS 0.036231f
C1349 VTAIL.n139 VSUBS 0.036231f
C1350 VTAIL.n140 VSUBS 0.01623f
C1351 VTAIL.n141 VSUBS 0.015328f
C1352 VTAIL.n142 VSUBS 0.028526f
C1353 VTAIL.n143 VSUBS 0.028526f
C1354 VTAIL.n144 VSUBS 0.015328f
C1355 VTAIL.n145 VSUBS 0.01623f
C1356 VTAIL.n146 VSUBS 0.036231f
C1357 VTAIL.n147 VSUBS 0.036231f
C1358 VTAIL.n148 VSUBS 0.01623f
C1359 VTAIL.n149 VSUBS 0.015328f
C1360 VTAIL.n150 VSUBS 0.028526f
C1361 VTAIL.n151 VSUBS 0.028526f
C1362 VTAIL.n152 VSUBS 0.015328f
C1363 VTAIL.n153 VSUBS 0.01623f
C1364 VTAIL.n154 VSUBS 0.036231f
C1365 VTAIL.n155 VSUBS 0.036231f
C1366 VTAIL.n156 VSUBS 0.082362f
C1367 VTAIL.n157 VSUBS 0.015779f
C1368 VTAIL.n158 VSUBS 0.015328f
C1369 VTAIL.n159 VSUBS 0.070612f
C1370 VTAIL.n160 VSUBS 0.041321f
C1371 VTAIL.n161 VSUBS 0.443402f
C1372 VTAIL.t7 VSUBS 0.316487f
C1373 VTAIL.t6 VSUBS 0.316487f
C1374 VTAIL.n162 VSUBS 2.39971f
C1375 VTAIL.n163 VSUBS 1.06192f
C1376 VTAIL.n164 VSUBS 0.029773f
C1377 VTAIL.n165 VSUBS 0.028526f
C1378 VTAIL.n166 VSUBS 0.015779f
C1379 VTAIL.n167 VSUBS 0.036231f
C1380 VTAIL.n168 VSUBS 0.015328f
C1381 VTAIL.n169 VSUBS 0.01623f
C1382 VTAIL.n170 VSUBS 0.028526f
C1383 VTAIL.n171 VSUBS 0.015328f
C1384 VTAIL.n172 VSUBS 0.036231f
C1385 VTAIL.n173 VSUBS 0.01623f
C1386 VTAIL.n174 VSUBS 0.028526f
C1387 VTAIL.n175 VSUBS 0.015328f
C1388 VTAIL.n176 VSUBS 0.036231f
C1389 VTAIL.n177 VSUBS 0.01623f
C1390 VTAIL.n178 VSUBS 0.028526f
C1391 VTAIL.n179 VSUBS 0.015328f
C1392 VTAIL.n180 VSUBS 0.036231f
C1393 VTAIL.n181 VSUBS 0.01623f
C1394 VTAIL.n182 VSUBS 0.028526f
C1395 VTAIL.n183 VSUBS 0.015328f
C1396 VTAIL.n184 VSUBS 0.036231f
C1397 VTAIL.n185 VSUBS 0.01623f
C1398 VTAIL.n186 VSUBS 0.028526f
C1399 VTAIL.n187 VSUBS 0.015328f
C1400 VTAIL.n188 VSUBS 0.027173f
C1401 VTAIL.n189 VSUBS 0.023048f
C1402 VTAIL.t10 VSUBS 0.077496f
C1403 VTAIL.n190 VSUBS 0.193004f
C1404 VTAIL.n191 VSUBS 1.6971f
C1405 VTAIL.n192 VSUBS 0.015328f
C1406 VTAIL.n193 VSUBS 0.01623f
C1407 VTAIL.n194 VSUBS 0.036231f
C1408 VTAIL.n195 VSUBS 0.036231f
C1409 VTAIL.n196 VSUBS 0.01623f
C1410 VTAIL.n197 VSUBS 0.015328f
C1411 VTAIL.n198 VSUBS 0.028526f
C1412 VTAIL.n199 VSUBS 0.028526f
C1413 VTAIL.n200 VSUBS 0.015328f
C1414 VTAIL.n201 VSUBS 0.01623f
C1415 VTAIL.n202 VSUBS 0.036231f
C1416 VTAIL.n203 VSUBS 0.036231f
C1417 VTAIL.n204 VSUBS 0.01623f
C1418 VTAIL.n205 VSUBS 0.015328f
C1419 VTAIL.n206 VSUBS 0.028526f
C1420 VTAIL.n207 VSUBS 0.028526f
C1421 VTAIL.n208 VSUBS 0.015328f
C1422 VTAIL.n209 VSUBS 0.01623f
C1423 VTAIL.n210 VSUBS 0.036231f
C1424 VTAIL.n211 VSUBS 0.036231f
C1425 VTAIL.n212 VSUBS 0.01623f
C1426 VTAIL.n213 VSUBS 0.015328f
C1427 VTAIL.n214 VSUBS 0.028526f
C1428 VTAIL.n215 VSUBS 0.028526f
C1429 VTAIL.n216 VSUBS 0.015328f
C1430 VTAIL.n217 VSUBS 0.01623f
C1431 VTAIL.n218 VSUBS 0.036231f
C1432 VTAIL.n219 VSUBS 0.036231f
C1433 VTAIL.n220 VSUBS 0.01623f
C1434 VTAIL.n221 VSUBS 0.015328f
C1435 VTAIL.n222 VSUBS 0.028526f
C1436 VTAIL.n223 VSUBS 0.028526f
C1437 VTAIL.n224 VSUBS 0.015328f
C1438 VTAIL.n225 VSUBS 0.01623f
C1439 VTAIL.n226 VSUBS 0.036231f
C1440 VTAIL.n227 VSUBS 0.036231f
C1441 VTAIL.n228 VSUBS 0.01623f
C1442 VTAIL.n229 VSUBS 0.015328f
C1443 VTAIL.n230 VSUBS 0.028526f
C1444 VTAIL.n231 VSUBS 0.028526f
C1445 VTAIL.n232 VSUBS 0.015328f
C1446 VTAIL.n233 VSUBS 0.01623f
C1447 VTAIL.n234 VSUBS 0.036231f
C1448 VTAIL.n235 VSUBS 0.036231f
C1449 VTAIL.n236 VSUBS 0.082362f
C1450 VTAIL.n237 VSUBS 0.015779f
C1451 VTAIL.n238 VSUBS 0.015328f
C1452 VTAIL.n239 VSUBS 0.070612f
C1453 VTAIL.n240 VSUBS 0.041321f
C1454 VTAIL.n241 VSUBS 2.02461f
C1455 VTAIL.n242 VSUBS 0.029773f
C1456 VTAIL.n243 VSUBS 0.028526f
C1457 VTAIL.n244 VSUBS 0.015779f
C1458 VTAIL.n245 VSUBS 0.036231f
C1459 VTAIL.n246 VSUBS 0.01623f
C1460 VTAIL.n247 VSUBS 0.028526f
C1461 VTAIL.n248 VSUBS 0.015328f
C1462 VTAIL.n249 VSUBS 0.036231f
C1463 VTAIL.n250 VSUBS 0.01623f
C1464 VTAIL.n251 VSUBS 0.028526f
C1465 VTAIL.n252 VSUBS 0.015328f
C1466 VTAIL.n253 VSUBS 0.036231f
C1467 VTAIL.n254 VSUBS 0.01623f
C1468 VTAIL.n255 VSUBS 0.028526f
C1469 VTAIL.n256 VSUBS 0.015328f
C1470 VTAIL.n257 VSUBS 0.036231f
C1471 VTAIL.n258 VSUBS 0.01623f
C1472 VTAIL.n259 VSUBS 0.028526f
C1473 VTAIL.n260 VSUBS 0.015328f
C1474 VTAIL.n261 VSUBS 0.036231f
C1475 VTAIL.n262 VSUBS 0.01623f
C1476 VTAIL.n263 VSUBS 0.028526f
C1477 VTAIL.n264 VSUBS 0.015328f
C1478 VTAIL.n265 VSUBS 0.027173f
C1479 VTAIL.n266 VSUBS 0.023048f
C1480 VTAIL.t1 VSUBS 0.077496f
C1481 VTAIL.n267 VSUBS 0.193004f
C1482 VTAIL.n268 VSUBS 1.6971f
C1483 VTAIL.n269 VSUBS 0.015328f
C1484 VTAIL.n270 VSUBS 0.01623f
C1485 VTAIL.n271 VSUBS 0.036231f
C1486 VTAIL.n272 VSUBS 0.036231f
C1487 VTAIL.n273 VSUBS 0.01623f
C1488 VTAIL.n274 VSUBS 0.015328f
C1489 VTAIL.n275 VSUBS 0.028526f
C1490 VTAIL.n276 VSUBS 0.028526f
C1491 VTAIL.n277 VSUBS 0.015328f
C1492 VTAIL.n278 VSUBS 0.01623f
C1493 VTAIL.n279 VSUBS 0.036231f
C1494 VTAIL.n280 VSUBS 0.036231f
C1495 VTAIL.n281 VSUBS 0.01623f
C1496 VTAIL.n282 VSUBS 0.015328f
C1497 VTAIL.n283 VSUBS 0.028526f
C1498 VTAIL.n284 VSUBS 0.028526f
C1499 VTAIL.n285 VSUBS 0.015328f
C1500 VTAIL.n286 VSUBS 0.01623f
C1501 VTAIL.n287 VSUBS 0.036231f
C1502 VTAIL.n288 VSUBS 0.036231f
C1503 VTAIL.n289 VSUBS 0.01623f
C1504 VTAIL.n290 VSUBS 0.015328f
C1505 VTAIL.n291 VSUBS 0.028526f
C1506 VTAIL.n292 VSUBS 0.028526f
C1507 VTAIL.n293 VSUBS 0.015328f
C1508 VTAIL.n294 VSUBS 0.01623f
C1509 VTAIL.n295 VSUBS 0.036231f
C1510 VTAIL.n296 VSUBS 0.036231f
C1511 VTAIL.n297 VSUBS 0.01623f
C1512 VTAIL.n298 VSUBS 0.015328f
C1513 VTAIL.n299 VSUBS 0.028526f
C1514 VTAIL.n300 VSUBS 0.028526f
C1515 VTAIL.n301 VSUBS 0.015328f
C1516 VTAIL.n302 VSUBS 0.01623f
C1517 VTAIL.n303 VSUBS 0.036231f
C1518 VTAIL.n304 VSUBS 0.036231f
C1519 VTAIL.n305 VSUBS 0.01623f
C1520 VTAIL.n306 VSUBS 0.015328f
C1521 VTAIL.n307 VSUBS 0.028526f
C1522 VTAIL.n308 VSUBS 0.028526f
C1523 VTAIL.n309 VSUBS 0.015328f
C1524 VTAIL.n310 VSUBS 0.015328f
C1525 VTAIL.n311 VSUBS 0.01623f
C1526 VTAIL.n312 VSUBS 0.036231f
C1527 VTAIL.n313 VSUBS 0.036231f
C1528 VTAIL.n314 VSUBS 0.082362f
C1529 VTAIL.n315 VSUBS 0.015779f
C1530 VTAIL.n316 VSUBS 0.015328f
C1531 VTAIL.n317 VSUBS 0.070612f
C1532 VTAIL.n318 VSUBS 0.041321f
C1533 VTAIL.n319 VSUBS 1.95706f
C1534 VP.n0 VSUBS 0.037669f
C1535 VP.t1 VSUBS 3.0842f
C1536 VP.n1 VSUBS 0.053741f
C1537 VP.n2 VSUBS 0.028573f
C1538 VP.t2 VSUBS 3.0842f
C1539 VP.n3 VSUBS 1.10606f
C1540 VP.n4 VSUBS 0.028573f
C1541 VP.n5 VSUBS 0.053741f
C1542 VP.n6 VSUBS 0.037669f
C1543 VP.t5 VSUBS 3.0842f
C1544 VP.n7 VSUBS 0.037669f
C1545 VP.t0 VSUBS 3.0842f
C1546 VP.n8 VSUBS 0.053741f
C1547 VP.n9 VSUBS 0.028573f
C1548 VP.t3 VSUBS 3.0842f
C1549 VP.n10 VSUBS 1.18096f
C1550 VP.t4 VSUBS 3.36879f
C1551 VP.n11 VSUBS 1.12154f
C1552 VP.n12 VSUBS 0.30002f
C1553 VP.n13 VSUBS 0.052987f
C1554 VP.n14 VSUBS 0.057404f
C1555 VP.n15 VSUBS 0.024914f
C1556 VP.n16 VSUBS 0.028573f
C1557 VP.n17 VSUBS 0.028573f
C1558 VP.n18 VSUBS 0.028573f
C1559 VP.n19 VSUBS 0.052987f
C1560 VP.n20 VSUBS 0.034153f
C1561 VP.n21 VSUBS 1.17749f
C1562 VP.n22 VSUBS 1.64455f
C1563 VP.n23 VSUBS 1.66472f
C1564 VP.n24 VSUBS 1.17749f
C1565 VP.n25 VSUBS 0.034153f
C1566 VP.n26 VSUBS 0.052987f
C1567 VP.n27 VSUBS 0.028573f
C1568 VP.n28 VSUBS 0.028573f
C1569 VP.n29 VSUBS 0.028573f
C1570 VP.n30 VSUBS 0.024914f
C1571 VP.n31 VSUBS 0.057404f
C1572 VP.n32 VSUBS 0.052987f
C1573 VP.n33 VSUBS 0.028573f
C1574 VP.n34 VSUBS 0.028573f
C1575 VP.n35 VSUBS 0.028573f
C1576 VP.n36 VSUBS 0.052987f
C1577 VP.n37 VSUBS 0.057404f
C1578 VP.n38 VSUBS 0.024914f
C1579 VP.n39 VSUBS 0.028573f
C1580 VP.n40 VSUBS 0.028573f
C1581 VP.n41 VSUBS 0.028573f
C1582 VP.n42 VSUBS 0.052987f
C1583 VP.n43 VSUBS 0.034153f
C1584 VP.n44 VSUBS 1.17749f
C1585 VP.n45 VSUBS 0.050745f
.ends

