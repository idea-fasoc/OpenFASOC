* NGSPICE file created from diff_pair_sample_1346.ext - technology: sky130A

.subckt diff_pair_sample_1346 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=7.1253 pd=37.32 as=0 ps=0 w=18.27 l=1.89
X1 VDD1.t7 VP.t0 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=3.01455 pd=18.6 as=7.1253 ps=37.32 w=18.27 l=1.89
X2 VTAIL.t7 VN.t0 VDD2.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=3.01455 pd=18.6 as=3.01455 ps=18.6 w=18.27 l=1.89
X3 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=7.1253 pd=37.32 as=0 ps=0 w=18.27 l=1.89
X4 VDD1.t6 VP.t1 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=3.01455 pd=18.6 as=7.1253 ps=37.32 w=18.27 l=1.89
X5 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=7.1253 pd=37.32 as=0 ps=0 w=18.27 l=1.89
X6 VTAIL.t3 VN.t1 VDD2.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=7.1253 pd=37.32 as=3.01455 ps=18.6 w=18.27 l=1.89
X7 VTAIL.t2 VN.t2 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=3.01455 pd=18.6 as=3.01455 ps=18.6 w=18.27 l=1.89
X8 VTAIL.t5 VN.t3 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=7.1253 pd=37.32 as=3.01455 ps=18.6 w=18.27 l=1.89
X9 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.1253 pd=37.32 as=0 ps=0 w=18.27 l=1.89
X10 VTAIL.t10 VP.t2 VDD1.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=7.1253 pd=37.32 as=3.01455 ps=18.6 w=18.27 l=1.89
X11 VTAIL.t11 VP.t3 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=7.1253 pd=37.32 as=3.01455 ps=18.6 w=18.27 l=1.89
X12 VDD2.t3 VN.t4 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=3.01455 pd=18.6 as=7.1253 ps=37.32 w=18.27 l=1.89
X13 VDD2.t2 VN.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.01455 pd=18.6 as=3.01455 ps=18.6 w=18.27 l=1.89
X14 VTAIL.t14 VP.t4 VDD1.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=3.01455 pd=18.6 as=3.01455 ps=18.6 w=18.27 l=1.89
X15 VTAIL.t8 VP.t5 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.01455 pd=18.6 as=3.01455 ps=18.6 w=18.27 l=1.89
X16 VDD2.t1 VN.t6 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.01455 pd=18.6 as=7.1253 ps=37.32 w=18.27 l=1.89
X17 VDD2.t0 VN.t7 VTAIL.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=3.01455 pd=18.6 as=3.01455 ps=18.6 w=18.27 l=1.89
X18 VDD1.t1 VP.t6 VTAIL.t15 B.t1 sky130_fd_pr__nfet_01v8 ad=3.01455 pd=18.6 as=3.01455 ps=18.6 w=18.27 l=1.89
X19 VDD1.t0 VP.t7 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=3.01455 pd=18.6 as=3.01455 ps=18.6 w=18.27 l=1.89
R0 B.n985 B.n984 585
R1 B.n402 B.n141 585
R2 B.n401 B.n400 585
R3 B.n399 B.n398 585
R4 B.n397 B.n396 585
R5 B.n395 B.n394 585
R6 B.n393 B.n392 585
R7 B.n391 B.n390 585
R8 B.n389 B.n388 585
R9 B.n387 B.n386 585
R10 B.n385 B.n384 585
R11 B.n383 B.n382 585
R12 B.n381 B.n380 585
R13 B.n379 B.n378 585
R14 B.n377 B.n376 585
R15 B.n375 B.n374 585
R16 B.n373 B.n372 585
R17 B.n371 B.n370 585
R18 B.n369 B.n368 585
R19 B.n367 B.n366 585
R20 B.n365 B.n364 585
R21 B.n363 B.n362 585
R22 B.n361 B.n360 585
R23 B.n359 B.n358 585
R24 B.n357 B.n356 585
R25 B.n355 B.n354 585
R26 B.n353 B.n352 585
R27 B.n351 B.n350 585
R28 B.n349 B.n348 585
R29 B.n347 B.n346 585
R30 B.n345 B.n344 585
R31 B.n343 B.n342 585
R32 B.n341 B.n340 585
R33 B.n339 B.n338 585
R34 B.n337 B.n336 585
R35 B.n335 B.n334 585
R36 B.n333 B.n332 585
R37 B.n331 B.n330 585
R38 B.n329 B.n328 585
R39 B.n327 B.n326 585
R40 B.n325 B.n324 585
R41 B.n323 B.n322 585
R42 B.n321 B.n320 585
R43 B.n319 B.n318 585
R44 B.n317 B.n316 585
R45 B.n315 B.n314 585
R46 B.n313 B.n312 585
R47 B.n311 B.n310 585
R48 B.n309 B.n308 585
R49 B.n307 B.n306 585
R50 B.n305 B.n304 585
R51 B.n303 B.n302 585
R52 B.n301 B.n300 585
R53 B.n299 B.n298 585
R54 B.n297 B.n296 585
R55 B.n295 B.n294 585
R56 B.n293 B.n292 585
R57 B.n291 B.n290 585
R58 B.n289 B.n288 585
R59 B.n287 B.n286 585
R60 B.n285 B.n284 585
R61 B.n283 B.n282 585
R62 B.n281 B.n280 585
R63 B.n279 B.n278 585
R64 B.n277 B.n276 585
R65 B.n275 B.n274 585
R66 B.n273 B.n272 585
R67 B.n271 B.n270 585
R68 B.n269 B.n268 585
R69 B.n267 B.n266 585
R70 B.n265 B.n264 585
R71 B.n263 B.n262 585
R72 B.n261 B.n260 585
R73 B.n259 B.n258 585
R74 B.n257 B.n256 585
R75 B.n255 B.n254 585
R76 B.n253 B.n252 585
R77 B.n251 B.n250 585
R78 B.n249 B.n248 585
R79 B.n247 B.n246 585
R80 B.n245 B.n244 585
R81 B.n243 B.n242 585
R82 B.n241 B.n240 585
R83 B.n239 B.n238 585
R84 B.n237 B.n236 585
R85 B.n235 B.n234 585
R86 B.n233 B.n232 585
R87 B.n231 B.n230 585
R88 B.n229 B.n228 585
R89 B.n227 B.n226 585
R90 B.n225 B.n224 585
R91 B.n223 B.n222 585
R92 B.n221 B.n220 585
R93 B.n219 B.n218 585
R94 B.n217 B.n216 585
R95 B.n215 B.n214 585
R96 B.n213 B.n212 585
R97 B.n211 B.n210 585
R98 B.n209 B.n208 585
R99 B.n207 B.n206 585
R100 B.n205 B.n204 585
R101 B.n203 B.n202 585
R102 B.n201 B.n200 585
R103 B.n199 B.n198 585
R104 B.n197 B.n196 585
R105 B.n195 B.n194 585
R106 B.n193 B.n192 585
R107 B.n191 B.n190 585
R108 B.n189 B.n188 585
R109 B.n187 B.n186 585
R110 B.n185 B.n184 585
R111 B.n183 B.n182 585
R112 B.n181 B.n180 585
R113 B.n179 B.n178 585
R114 B.n177 B.n176 585
R115 B.n175 B.n174 585
R116 B.n173 B.n172 585
R117 B.n171 B.n170 585
R118 B.n169 B.n168 585
R119 B.n167 B.n166 585
R120 B.n165 B.n164 585
R121 B.n163 B.n162 585
R122 B.n161 B.n160 585
R123 B.n159 B.n158 585
R124 B.n157 B.n156 585
R125 B.n155 B.n154 585
R126 B.n153 B.n152 585
R127 B.n151 B.n150 585
R128 B.n149 B.n148 585
R129 B.n75 B.n74 585
R130 B.n983 B.n76 585
R131 B.n988 B.n76 585
R132 B.n982 B.n981 585
R133 B.n981 B.n72 585
R134 B.n980 B.n71 585
R135 B.n994 B.n71 585
R136 B.n979 B.n70 585
R137 B.n995 B.n70 585
R138 B.n978 B.n69 585
R139 B.n996 B.n69 585
R140 B.n977 B.n976 585
R141 B.n976 B.n65 585
R142 B.n975 B.n64 585
R143 B.n1002 B.n64 585
R144 B.n974 B.n63 585
R145 B.n1003 B.n63 585
R146 B.n973 B.n62 585
R147 B.n1004 B.n62 585
R148 B.n972 B.n971 585
R149 B.n971 B.n58 585
R150 B.n970 B.n57 585
R151 B.n1010 B.n57 585
R152 B.n969 B.n56 585
R153 B.n1011 B.n56 585
R154 B.n968 B.n55 585
R155 B.n1012 B.n55 585
R156 B.n967 B.n966 585
R157 B.n966 B.n51 585
R158 B.n965 B.n50 585
R159 B.n1018 B.n50 585
R160 B.n964 B.n49 585
R161 B.n1019 B.n49 585
R162 B.n963 B.n48 585
R163 B.n1020 B.n48 585
R164 B.n962 B.n961 585
R165 B.n961 B.n44 585
R166 B.n960 B.n43 585
R167 B.n1026 B.n43 585
R168 B.n959 B.n42 585
R169 B.n1027 B.n42 585
R170 B.n958 B.n41 585
R171 B.n1028 B.n41 585
R172 B.n957 B.n956 585
R173 B.n956 B.n37 585
R174 B.n955 B.n36 585
R175 B.n1034 B.n36 585
R176 B.n954 B.n35 585
R177 B.n1035 B.n35 585
R178 B.n953 B.n34 585
R179 B.n1036 B.n34 585
R180 B.n952 B.n951 585
R181 B.n951 B.n30 585
R182 B.n950 B.n29 585
R183 B.n1042 B.n29 585
R184 B.n949 B.n28 585
R185 B.n1043 B.n28 585
R186 B.n948 B.n27 585
R187 B.n1044 B.n27 585
R188 B.n947 B.n946 585
R189 B.n946 B.n26 585
R190 B.n945 B.n22 585
R191 B.n1050 B.n22 585
R192 B.n944 B.n21 585
R193 B.n1051 B.n21 585
R194 B.n943 B.n20 585
R195 B.n1052 B.n20 585
R196 B.n942 B.n941 585
R197 B.n941 B.n16 585
R198 B.n940 B.n15 585
R199 B.n1058 B.n15 585
R200 B.n939 B.n14 585
R201 B.n1059 B.n14 585
R202 B.n938 B.n13 585
R203 B.n1060 B.n13 585
R204 B.n937 B.n936 585
R205 B.n936 B.n12 585
R206 B.n935 B.n934 585
R207 B.n935 B.n8 585
R208 B.n933 B.n7 585
R209 B.n1067 B.n7 585
R210 B.n932 B.n6 585
R211 B.n1068 B.n6 585
R212 B.n931 B.n5 585
R213 B.n1069 B.n5 585
R214 B.n930 B.n929 585
R215 B.n929 B.n4 585
R216 B.n928 B.n403 585
R217 B.n928 B.n927 585
R218 B.n918 B.n404 585
R219 B.n405 B.n404 585
R220 B.n920 B.n919 585
R221 B.n921 B.n920 585
R222 B.n917 B.n409 585
R223 B.n413 B.n409 585
R224 B.n916 B.n915 585
R225 B.n915 B.n914 585
R226 B.n411 B.n410 585
R227 B.n412 B.n411 585
R228 B.n907 B.n906 585
R229 B.n908 B.n907 585
R230 B.n905 B.n418 585
R231 B.n418 B.n417 585
R232 B.n904 B.n903 585
R233 B.n903 B.n902 585
R234 B.n420 B.n419 585
R235 B.n895 B.n420 585
R236 B.n894 B.n893 585
R237 B.n896 B.n894 585
R238 B.n892 B.n425 585
R239 B.n425 B.n424 585
R240 B.n891 B.n890 585
R241 B.n890 B.n889 585
R242 B.n427 B.n426 585
R243 B.n428 B.n427 585
R244 B.n882 B.n881 585
R245 B.n883 B.n882 585
R246 B.n880 B.n433 585
R247 B.n433 B.n432 585
R248 B.n879 B.n878 585
R249 B.n878 B.n877 585
R250 B.n435 B.n434 585
R251 B.n436 B.n435 585
R252 B.n870 B.n869 585
R253 B.n871 B.n870 585
R254 B.n868 B.n441 585
R255 B.n441 B.n440 585
R256 B.n867 B.n866 585
R257 B.n866 B.n865 585
R258 B.n443 B.n442 585
R259 B.n444 B.n443 585
R260 B.n858 B.n857 585
R261 B.n859 B.n858 585
R262 B.n856 B.n449 585
R263 B.n449 B.n448 585
R264 B.n855 B.n854 585
R265 B.n854 B.n853 585
R266 B.n451 B.n450 585
R267 B.n452 B.n451 585
R268 B.n846 B.n845 585
R269 B.n847 B.n846 585
R270 B.n844 B.n457 585
R271 B.n457 B.n456 585
R272 B.n843 B.n842 585
R273 B.n842 B.n841 585
R274 B.n459 B.n458 585
R275 B.n460 B.n459 585
R276 B.n834 B.n833 585
R277 B.n835 B.n834 585
R278 B.n832 B.n465 585
R279 B.n465 B.n464 585
R280 B.n831 B.n830 585
R281 B.n830 B.n829 585
R282 B.n467 B.n466 585
R283 B.n468 B.n467 585
R284 B.n822 B.n821 585
R285 B.n823 B.n822 585
R286 B.n820 B.n473 585
R287 B.n473 B.n472 585
R288 B.n819 B.n818 585
R289 B.n818 B.n817 585
R290 B.n475 B.n474 585
R291 B.n476 B.n475 585
R292 B.n810 B.n809 585
R293 B.n811 B.n810 585
R294 B.n479 B.n478 585
R295 B.n550 B.n548 585
R296 B.n551 B.n547 585
R297 B.n551 B.n480 585
R298 B.n554 B.n553 585
R299 B.n555 B.n546 585
R300 B.n557 B.n556 585
R301 B.n559 B.n545 585
R302 B.n562 B.n561 585
R303 B.n563 B.n544 585
R304 B.n565 B.n564 585
R305 B.n567 B.n543 585
R306 B.n570 B.n569 585
R307 B.n571 B.n542 585
R308 B.n573 B.n572 585
R309 B.n575 B.n541 585
R310 B.n578 B.n577 585
R311 B.n579 B.n540 585
R312 B.n581 B.n580 585
R313 B.n583 B.n539 585
R314 B.n586 B.n585 585
R315 B.n587 B.n538 585
R316 B.n589 B.n588 585
R317 B.n591 B.n537 585
R318 B.n594 B.n593 585
R319 B.n595 B.n536 585
R320 B.n597 B.n596 585
R321 B.n599 B.n535 585
R322 B.n602 B.n601 585
R323 B.n603 B.n534 585
R324 B.n605 B.n604 585
R325 B.n607 B.n533 585
R326 B.n610 B.n609 585
R327 B.n611 B.n532 585
R328 B.n613 B.n612 585
R329 B.n615 B.n531 585
R330 B.n618 B.n617 585
R331 B.n619 B.n530 585
R332 B.n621 B.n620 585
R333 B.n623 B.n529 585
R334 B.n626 B.n625 585
R335 B.n627 B.n528 585
R336 B.n629 B.n628 585
R337 B.n631 B.n527 585
R338 B.n634 B.n633 585
R339 B.n635 B.n526 585
R340 B.n637 B.n636 585
R341 B.n639 B.n525 585
R342 B.n642 B.n641 585
R343 B.n643 B.n524 585
R344 B.n645 B.n644 585
R345 B.n647 B.n523 585
R346 B.n650 B.n649 585
R347 B.n651 B.n522 585
R348 B.n653 B.n652 585
R349 B.n655 B.n521 585
R350 B.n658 B.n657 585
R351 B.n659 B.n520 585
R352 B.n661 B.n660 585
R353 B.n663 B.n519 585
R354 B.n666 B.n665 585
R355 B.n668 B.n516 585
R356 B.n670 B.n669 585
R357 B.n672 B.n515 585
R358 B.n675 B.n674 585
R359 B.n676 B.n514 585
R360 B.n678 B.n677 585
R361 B.n680 B.n513 585
R362 B.n683 B.n682 585
R363 B.n684 B.n512 585
R364 B.n689 B.n688 585
R365 B.n691 B.n511 585
R366 B.n694 B.n693 585
R367 B.n695 B.n510 585
R368 B.n697 B.n696 585
R369 B.n699 B.n509 585
R370 B.n702 B.n701 585
R371 B.n703 B.n508 585
R372 B.n705 B.n704 585
R373 B.n707 B.n507 585
R374 B.n710 B.n709 585
R375 B.n711 B.n506 585
R376 B.n713 B.n712 585
R377 B.n715 B.n505 585
R378 B.n718 B.n717 585
R379 B.n719 B.n504 585
R380 B.n721 B.n720 585
R381 B.n723 B.n503 585
R382 B.n726 B.n725 585
R383 B.n727 B.n502 585
R384 B.n729 B.n728 585
R385 B.n731 B.n501 585
R386 B.n734 B.n733 585
R387 B.n735 B.n500 585
R388 B.n737 B.n736 585
R389 B.n739 B.n499 585
R390 B.n742 B.n741 585
R391 B.n743 B.n498 585
R392 B.n745 B.n744 585
R393 B.n747 B.n497 585
R394 B.n750 B.n749 585
R395 B.n751 B.n496 585
R396 B.n753 B.n752 585
R397 B.n755 B.n495 585
R398 B.n758 B.n757 585
R399 B.n759 B.n494 585
R400 B.n761 B.n760 585
R401 B.n763 B.n493 585
R402 B.n766 B.n765 585
R403 B.n767 B.n492 585
R404 B.n769 B.n768 585
R405 B.n771 B.n491 585
R406 B.n774 B.n773 585
R407 B.n775 B.n490 585
R408 B.n777 B.n776 585
R409 B.n779 B.n489 585
R410 B.n782 B.n781 585
R411 B.n783 B.n488 585
R412 B.n785 B.n784 585
R413 B.n787 B.n487 585
R414 B.n790 B.n789 585
R415 B.n791 B.n486 585
R416 B.n793 B.n792 585
R417 B.n795 B.n485 585
R418 B.n798 B.n797 585
R419 B.n799 B.n484 585
R420 B.n801 B.n800 585
R421 B.n803 B.n483 585
R422 B.n804 B.n482 585
R423 B.n807 B.n806 585
R424 B.n808 B.n481 585
R425 B.n481 B.n480 585
R426 B.n813 B.n812 585
R427 B.n812 B.n811 585
R428 B.n814 B.n477 585
R429 B.n477 B.n476 585
R430 B.n816 B.n815 585
R431 B.n817 B.n816 585
R432 B.n471 B.n470 585
R433 B.n472 B.n471 585
R434 B.n825 B.n824 585
R435 B.n824 B.n823 585
R436 B.n826 B.n469 585
R437 B.n469 B.n468 585
R438 B.n828 B.n827 585
R439 B.n829 B.n828 585
R440 B.n463 B.n462 585
R441 B.n464 B.n463 585
R442 B.n837 B.n836 585
R443 B.n836 B.n835 585
R444 B.n838 B.n461 585
R445 B.n461 B.n460 585
R446 B.n840 B.n839 585
R447 B.n841 B.n840 585
R448 B.n455 B.n454 585
R449 B.n456 B.n455 585
R450 B.n849 B.n848 585
R451 B.n848 B.n847 585
R452 B.n850 B.n453 585
R453 B.n453 B.n452 585
R454 B.n852 B.n851 585
R455 B.n853 B.n852 585
R456 B.n447 B.n446 585
R457 B.n448 B.n447 585
R458 B.n861 B.n860 585
R459 B.n860 B.n859 585
R460 B.n862 B.n445 585
R461 B.n445 B.n444 585
R462 B.n864 B.n863 585
R463 B.n865 B.n864 585
R464 B.n439 B.n438 585
R465 B.n440 B.n439 585
R466 B.n873 B.n872 585
R467 B.n872 B.n871 585
R468 B.n874 B.n437 585
R469 B.n437 B.n436 585
R470 B.n876 B.n875 585
R471 B.n877 B.n876 585
R472 B.n431 B.n430 585
R473 B.n432 B.n431 585
R474 B.n885 B.n884 585
R475 B.n884 B.n883 585
R476 B.n886 B.n429 585
R477 B.n429 B.n428 585
R478 B.n888 B.n887 585
R479 B.n889 B.n888 585
R480 B.n423 B.n422 585
R481 B.n424 B.n423 585
R482 B.n898 B.n897 585
R483 B.n897 B.n896 585
R484 B.n899 B.n421 585
R485 B.n895 B.n421 585
R486 B.n901 B.n900 585
R487 B.n902 B.n901 585
R488 B.n416 B.n415 585
R489 B.n417 B.n416 585
R490 B.n910 B.n909 585
R491 B.n909 B.n908 585
R492 B.n911 B.n414 585
R493 B.n414 B.n412 585
R494 B.n913 B.n912 585
R495 B.n914 B.n913 585
R496 B.n408 B.n407 585
R497 B.n413 B.n408 585
R498 B.n923 B.n922 585
R499 B.n922 B.n921 585
R500 B.n924 B.n406 585
R501 B.n406 B.n405 585
R502 B.n926 B.n925 585
R503 B.n927 B.n926 585
R504 B.n3 B.n0 585
R505 B.n4 B.n3 585
R506 B.n1066 B.n1 585
R507 B.n1067 B.n1066 585
R508 B.n1065 B.n1064 585
R509 B.n1065 B.n8 585
R510 B.n1063 B.n9 585
R511 B.n12 B.n9 585
R512 B.n1062 B.n1061 585
R513 B.n1061 B.n1060 585
R514 B.n11 B.n10 585
R515 B.n1059 B.n11 585
R516 B.n1057 B.n1056 585
R517 B.n1058 B.n1057 585
R518 B.n1055 B.n17 585
R519 B.n17 B.n16 585
R520 B.n1054 B.n1053 585
R521 B.n1053 B.n1052 585
R522 B.n19 B.n18 585
R523 B.n1051 B.n19 585
R524 B.n1049 B.n1048 585
R525 B.n1050 B.n1049 585
R526 B.n1047 B.n23 585
R527 B.n26 B.n23 585
R528 B.n1046 B.n1045 585
R529 B.n1045 B.n1044 585
R530 B.n25 B.n24 585
R531 B.n1043 B.n25 585
R532 B.n1041 B.n1040 585
R533 B.n1042 B.n1041 585
R534 B.n1039 B.n31 585
R535 B.n31 B.n30 585
R536 B.n1038 B.n1037 585
R537 B.n1037 B.n1036 585
R538 B.n33 B.n32 585
R539 B.n1035 B.n33 585
R540 B.n1033 B.n1032 585
R541 B.n1034 B.n1033 585
R542 B.n1031 B.n38 585
R543 B.n38 B.n37 585
R544 B.n1030 B.n1029 585
R545 B.n1029 B.n1028 585
R546 B.n40 B.n39 585
R547 B.n1027 B.n40 585
R548 B.n1025 B.n1024 585
R549 B.n1026 B.n1025 585
R550 B.n1023 B.n45 585
R551 B.n45 B.n44 585
R552 B.n1022 B.n1021 585
R553 B.n1021 B.n1020 585
R554 B.n47 B.n46 585
R555 B.n1019 B.n47 585
R556 B.n1017 B.n1016 585
R557 B.n1018 B.n1017 585
R558 B.n1015 B.n52 585
R559 B.n52 B.n51 585
R560 B.n1014 B.n1013 585
R561 B.n1013 B.n1012 585
R562 B.n54 B.n53 585
R563 B.n1011 B.n54 585
R564 B.n1009 B.n1008 585
R565 B.n1010 B.n1009 585
R566 B.n1007 B.n59 585
R567 B.n59 B.n58 585
R568 B.n1006 B.n1005 585
R569 B.n1005 B.n1004 585
R570 B.n61 B.n60 585
R571 B.n1003 B.n61 585
R572 B.n1001 B.n1000 585
R573 B.n1002 B.n1001 585
R574 B.n999 B.n66 585
R575 B.n66 B.n65 585
R576 B.n998 B.n997 585
R577 B.n997 B.n996 585
R578 B.n68 B.n67 585
R579 B.n995 B.n68 585
R580 B.n993 B.n992 585
R581 B.n994 B.n993 585
R582 B.n991 B.n73 585
R583 B.n73 B.n72 585
R584 B.n990 B.n989 585
R585 B.n989 B.n988 585
R586 B.n1070 B.n1069 585
R587 B.n1068 B.n2 585
R588 B.n989 B.n75 516.524
R589 B.n985 B.n76 516.524
R590 B.n810 B.n481 516.524
R591 B.n812 B.n479 516.524
R592 B.n145 B.t16 439.615
R593 B.n142 B.t12 439.615
R594 B.n685 B.t19 439.615
R595 B.n517 B.t8 439.615
R596 B.n142 B.t14 433.384
R597 B.n685 B.t21 433.384
R598 B.n145 B.t17 433.384
R599 B.n517 B.t11 433.384
R600 B.n143 B.t15 390.329
R601 B.n686 B.t20 390.329
R602 B.n146 B.t18 390.329
R603 B.n518 B.t10 390.329
R604 B.n987 B.n986 256.663
R605 B.n987 B.n140 256.663
R606 B.n987 B.n139 256.663
R607 B.n987 B.n138 256.663
R608 B.n987 B.n137 256.663
R609 B.n987 B.n136 256.663
R610 B.n987 B.n135 256.663
R611 B.n987 B.n134 256.663
R612 B.n987 B.n133 256.663
R613 B.n987 B.n132 256.663
R614 B.n987 B.n131 256.663
R615 B.n987 B.n130 256.663
R616 B.n987 B.n129 256.663
R617 B.n987 B.n128 256.663
R618 B.n987 B.n127 256.663
R619 B.n987 B.n126 256.663
R620 B.n987 B.n125 256.663
R621 B.n987 B.n124 256.663
R622 B.n987 B.n123 256.663
R623 B.n987 B.n122 256.663
R624 B.n987 B.n121 256.663
R625 B.n987 B.n120 256.663
R626 B.n987 B.n119 256.663
R627 B.n987 B.n118 256.663
R628 B.n987 B.n117 256.663
R629 B.n987 B.n116 256.663
R630 B.n987 B.n115 256.663
R631 B.n987 B.n114 256.663
R632 B.n987 B.n113 256.663
R633 B.n987 B.n112 256.663
R634 B.n987 B.n111 256.663
R635 B.n987 B.n110 256.663
R636 B.n987 B.n109 256.663
R637 B.n987 B.n108 256.663
R638 B.n987 B.n107 256.663
R639 B.n987 B.n106 256.663
R640 B.n987 B.n105 256.663
R641 B.n987 B.n104 256.663
R642 B.n987 B.n103 256.663
R643 B.n987 B.n102 256.663
R644 B.n987 B.n101 256.663
R645 B.n987 B.n100 256.663
R646 B.n987 B.n99 256.663
R647 B.n987 B.n98 256.663
R648 B.n987 B.n97 256.663
R649 B.n987 B.n96 256.663
R650 B.n987 B.n95 256.663
R651 B.n987 B.n94 256.663
R652 B.n987 B.n93 256.663
R653 B.n987 B.n92 256.663
R654 B.n987 B.n91 256.663
R655 B.n987 B.n90 256.663
R656 B.n987 B.n89 256.663
R657 B.n987 B.n88 256.663
R658 B.n987 B.n87 256.663
R659 B.n987 B.n86 256.663
R660 B.n987 B.n85 256.663
R661 B.n987 B.n84 256.663
R662 B.n987 B.n83 256.663
R663 B.n987 B.n82 256.663
R664 B.n987 B.n81 256.663
R665 B.n987 B.n80 256.663
R666 B.n987 B.n79 256.663
R667 B.n987 B.n78 256.663
R668 B.n987 B.n77 256.663
R669 B.n549 B.n480 256.663
R670 B.n552 B.n480 256.663
R671 B.n558 B.n480 256.663
R672 B.n560 B.n480 256.663
R673 B.n566 B.n480 256.663
R674 B.n568 B.n480 256.663
R675 B.n574 B.n480 256.663
R676 B.n576 B.n480 256.663
R677 B.n582 B.n480 256.663
R678 B.n584 B.n480 256.663
R679 B.n590 B.n480 256.663
R680 B.n592 B.n480 256.663
R681 B.n598 B.n480 256.663
R682 B.n600 B.n480 256.663
R683 B.n606 B.n480 256.663
R684 B.n608 B.n480 256.663
R685 B.n614 B.n480 256.663
R686 B.n616 B.n480 256.663
R687 B.n622 B.n480 256.663
R688 B.n624 B.n480 256.663
R689 B.n630 B.n480 256.663
R690 B.n632 B.n480 256.663
R691 B.n638 B.n480 256.663
R692 B.n640 B.n480 256.663
R693 B.n646 B.n480 256.663
R694 B.n648 B.n480 256.663
R695 B.n654 B.n480 256.663
R696 B.n656 B.n480 256.663
R697 B.n662 B.n480 256.663
R698 B.n664 B.n480 256.663
R699 B.n671 B.n480 256.663
R700 B.n673 B.n480 256.663
R701 B.n679 B.n480 256.663
R702 B.n681 B.n480 256.663
R703 B.n690 B.n480 256.663
R704 B.n692 B.n480 256.663
R705 B.n698 B.n480 256.663
R706 B.n700 B.n480 256.663
R707 B.n706 B.n480 256.663
R708 B.n708 B.n480 256.663
R709 B.n714 B.n480 256.663
R710 B.n716 B.n480 256.663
R711 B.n722 B.n480 256.663
R712 B.n724 B.n480 256.663
R713 B.n730 B.n480 256.663
R714 B.n732 B.n480 256.663
R715 B.n738 B.n480 256.663
R716 B.n740 B.n480 256.663
R717 B.n746 B.n480 256.663
R718 B.n748 B.n480 256.663
R719 B.n754 B.n480 256.663
R720 B.n756 B.n480 256.663
R721 B.n762 B.n480 256.663
R722 B.n764 B.n480 256.663
R723 B.n770 B.n480 256.663
R724 B.n772 B.n480 256.663
R725 B.n778 B.n480 256.663
R726 B.n780 B.n480 256.663
R727 B.n786 B.n480 256.663
R728 B.n788 B.n480 256.663
R729 B.n794 B.n480 256.663
R730 B.n796 B.n480 256.663
R731 B.n802 B.n480 256.663
R732 B.n805 B.n480 256.663
R733 B.n1072 B.n1071 256.663
R734 B.n150 B.n149 163.367
R735 B.n154 B.n153 163.367
R736 B.n158 B.n157 163.367
R737 B.n162 B.n161 163.367
R738 B.n166 B.n165 163.367
R739 B.n170 B.n169 163.367
R740 B.n174 B.n173 163.367
R741 B.n178 B.n177 163.367
R742 B.n182 B.n181 163.367
R743 B.n186 B.n185 163.367
R744 B.n190 B.n189 163.367
R745 B.n194 B.n193 163.367
R746 B.n198 B.n197 163.367
R747 B.n202 B.n201 163.367
R748 B.n206 B.n205 163.367
R749 B.n210 B.n209 163.367
R750 B.n214 B.n213 163.367
R751 B.n218 B.n217 163.367
R752 B.n222 B.n221 163.367
R753 B.n226 B.n225 163.367
R754 B.n230 B.n229 163.367
R755 B.n234 B.n233 163.367
R756 B.n238 B.n237 163.367
R757 B.n242 B.n241 163.367
R758 B.n246 B.n245 163.367
R759 B.n250 B.n249 163.367
R760 B.n254 B.n253 163.367
R761 B.n258 B.n257 163.367
R762 B.n262 B.n261 163.367
R763 B.n266 B.n265 163.367
R764 B.n270 B.n269 163.367
R765 B.n274 B.n273 163.367
R766 B.n278 B.n277 163.367
R767 B.n282 B.n281 163.367
R768 B.n286 B.n285 163.367
R769 B.n290 B.n289 163.367
R770 B.n294 B.n293 163.367
R771 B.n298 B.n297 163.367
R772 B.n302 B.n301 163.367
R773 B.n306 B.n305 163.367
R774 B.n310 B.n309 163.367
R775 B.n314 B.n313 163.367
R776 B.n318 B.n317 163.367
R777 B.n322 B.n321 163.367
R778 B.n326 B.n325 163.367
R779 B.n330 B.n329 163.367
R780 B.n334 B.n333 163.367
R781 B.n338 B.n337 163.367
R782 B.n342 B.n341 163.367
R783 B.n346 B.n345 163.367
R784 B.n350 B.n349 163.367
R785 B.n354 B.n353 163.367
R786 B.n358 B.n357 163.367
R787 B.n362 B.n361 163.367
R788 B.n366 B.n365 163.367
R789 B.n370 B.n369 163.367
R790 B.n374 B.n373 163.367
R791 B.n378 B.n377 163.367
R792 B.n382 B.n381 163.367
R793 B.n386 B.n385 163.367
R794 B.n390 B.n389 163.367
R795 B.n394 B.n393 163.367
R796 B.n398 B.n397 163.367
R797 B.n400 B.n141 163.367
R798 B.n810 B.n475 163.367
R799 B.n818 B.n475 163.367
R800 B.n818 B.n473 163.367
R801 B.n822 B.n473 163.367
R802 B.n822 B.n467 163.367
R803 B.n830 B.n467 163.367
R804 B.n830 B.n465 163.367
R805 B.n834 B.n465 163.367
R806 B.n834 B.n459 163.367
R807 B.n842 B.n459 163.367
R808 B.n842 B.n457 163.367
R809 B.n846 B.n457 163.367
R810 B.n846 B.n451 163.367
R811 B.n854 B.n451 163.367
R812 B.n854 B.n449 163.367
R813 B.n858 B.n449 163.367
R814 B.n858 B.n443 163.367
R815 B.n866 B.n443 163.367
R816 B.n866 B.n441 163.367
R817 B.n870 B.n441 163.367
R818 B.n870 B.n435 163.367
R819 B.n878 B.n435 163.367
R820 B.n878 B.n433 163.367
R821 B.n882 B.n433 163.367
R822 B.n882 B.n427 163.367
R823 B.n890 B.n427 163.367
R824 B.n890 B.n425 163.367
R825 B.n894 B.n425 163.367
R826 B.n894 B.n420 163.367
R827 B.n903 B.n420 163.367
R828 B.n903 B.n418 163.367
R829 B.n907 B.n418 163.367
R830 B.n907 B.n411 163.367
R831 B.n915 B.n411 163.367
R832 B.n915 B.n409 163.367
R833 B.n920 B.n409 163.367
R834 B.n920 B.n404 163.367
R835 B.n928 B.n404 163.367
R836 B.n929 B.n928 163.367
R837 B.n929 B.n5 163.367
R838 B.n6 B.n5 163.367
R839 B.n7 B.n6 163.367
R840 B.n935 B.n7 163.367
R841 B.n936 B.n935 163.367
R842 B.n936 B.n13 163.367
R843 B.n14 B.n13 163.367
R844 B.n15 B.n14 163.367
R845 B.n941 B.n15 163.367
R846 B.n941 B.n20 163.367
R847 B.n21 B.n20 163.367
R848 B.n22 B.n21 163.367
R849 B.n946 B.n22 163.367
R850 B.n946 B.n27 163.367
R851 B.n28 B.n27 163.367
R852 B.n29 B.n28 163.367
R853 B.n951 B.n29 163.367
R854 B.n951 B.n34 163.367
R855 B.n35 B.n34 163.367
R856 B.n36 B.n35 163.367
R857 B.n956 B.n36 163.367
R858 B.n956 B.n41 163.367
R859 B.n42 B.n41 163.367
R860 B.n43 B.n42 163.367
R861 B.n961 B.n43 163.367
R862 B.n961 B.n48 163.367
R863 B.n49 B.n48 163.367
R864 B.n50 B.n49 163.367
R865 B.n966 B.n50 163.367
R866 B.n966 B.n55 163.367
R867 B.n56 B.n55 163.367
R868 B.n57 B.n56 163.367
R869 B.n971 B.n57 163.367
R870 B.n971 B.n62 163.367
R871 B.n63 B.n62 163.367
R872 B.n64 B.n63 163.367
R873 B.n976 B.n64 163.367
R874 B.n976 B.n69 163.367
R875 B.n70 B.n69 163.367
R876 B.n71 B.n70 163.367
R877 B.n981 B.n71 163.367
R878 B.n981 B.n76 163.367
R879 B.n551 B.n550 163.367
R880 B.n553 B.n551 163.367
R881 B.n557 B.n546 163.367
R882 B.n561 B.n559 163.367
R883 B.n565 B.n544 163.367
R884 B.n569 B.n567 163.367
R885 B.n573 B.n542 163.367
R886 B.n577 B.n575 163.367
R887 B.n581 B.n540 163.367
R888 B.n585 B.n583 163.367
R889 B.n589 B.n538 163.367
R890 B.n593 B.n591 163.367
R891 B.n597 B.n536 163.367
R892 B.n601 B.n599 163.367
R893 B.n605 B.n534 163.367
R894 B.n609 B.n607 163.367
R895 B.n613 B.n532 163.367
R896 B.n617 B.n615 163.367
R897 B.n621 B.n530 163.367
R898 B.n625 B.n623 163.367
R899 B.n629 B.n528 163.367
R900 B.n633 B.n631 163.367
R901 B.n637 B.n526 163.367
R902 B.n641 B.n639 163.367
R903 B.n645 B.n524 163.367
R904 B.n649 B.n647 163.367
R905 B.n653 B.n522 163.367
R906 B.n657 B.n655 163.367
R907 B.n661 B.n520 163.367
R908 B.n665 B.n663 163.367
R909 B.n670 B.n516 163.367
R910 B.n674 B.n672 163.367
R911 B.n678 B.n514 163.367
R912 B.n682 B.n680 163.367
R913 B.n689 B.n512 163.367
R914 B.n693 B.n691 163.367
R915 B.n697 B.n510 163.367
R916 B.n701 B.n699 163.367
R917 B.n705 B.n508 163.367
R918 B.n709 B.n707 163.367
R919 B.n713 B.n506 163.367
R920 B.n717 B.n715 163.367
R921 B.n721 B.n504 163.367
R922 B.n725 B.n723 163.367
R923 B.n729 B.n502 163.367
R924 B.n733 B.n731 163.367
R925 B.n737 B.n500 163.367
R926 B.n741 B.n739 163.367
R927 B.n745 B.n498 163.367
R928 B.n749 B.n747 163.367
R929 B.n753 B.n496 163.367
R930 B.n757 B.n755 163.367
R931 B.n761 B.n494 163.367
R932 B.n765 B.n763 163.367
R933 B.n769 B.n492 163.367
R934 B.n773 B.n771 163.367
R935 B.n777 B.n490 163.367
R936 B.n781 B.n779 163.367
R937 B.n785 B.n488 163.367
R938 B.n789 B.n787 163.367
R939 B.n793 B.n486 163.367
R940 B.n797 B.n795 163.367
R941 B.n801 B.n484 163.367
R942 B.n804 B.n803 163.367
R943 B.n806 B.n481 163.367
R944 B.n812 B.n477 163.367
R945 B.n816 B.n477 163.367
R946 B.n816 B.n471 163.367
R947 B.n824 B.n471 163.367
R948 B.n824 B.n469 163.367
R949 B.n828 B.n469 163.367
R950 B.n828 B.n463 163.367
R951 B.n836 B.n463 163.367
R952 B.n836 B.n461 163.367
R953 B.n840 B.n461 163.367
R954 B.n840 B.n455 163.367
R955 B.n848 B.n455 163.367
R956 B.n848 B.n453 163.367
R957 B.n852 B.n453 163.367
R958 B.n852 B.n447 163.367
R959 B.n860 B.n447 163.367
R960 B.n860 B.n445 163.367
R961 B.n864 B.n445 163.367
R962 B.n864 B.n439 163.367
R963 B.n872 B.n439 163.367
R964 B.n872 B.n437 163.367
R965 B.n876 B.n437 163.367
R966 B.n876 B.n431 163.367
R967 B.n884 B.n431 163.367
R968 B.n884 B.n429 163.367
R969 B.n888 B.n429 163.367
R970 B.n888 B.n423 163.367
R971 B.n897 B.n423 163.367
R972 B.n897 B.n421 163.367
R973 B.n901 B.n421 163.367
R974 B.n901 B.n416 163.367
R975 B.n909 B.n416 163.367
R976 B.n909 B.n414 163.367
R977 B.n913 B.n414 163.367
R978 B.n913 B.n408 163.367
R979 B.n922 B.n408 163.367
R980 B.n922 B.n406 163.367
R981 B.n926 B.n406 163.367
R982 B.n926 B.n3 163.367
R983 B.n1070 B.n3 163.367
R984 B.n1066 B.n2 163.367
R985 B.n1066 B.n1065 163.367
R986 B.n1065 B.n9 163.367
R987 B.n1061 B.n9 163.367
R988 B.n1061 B.n11 163.367
R989 B.n1057 B.n11 163.367
R990 B.n1057 B.n17 163.367
R991 B.n1053 B.n17 163.367
R992 B.n1053 B.n19 163.367
R993 B.n1049 B.n19 163.367
R994 B.n1049 B.n23 163.367
R995 B.n1045 B.n23 163.367
R996 B.n1045 B.n25 163.367
R997 B.n1041 B.n25 163.367
R998 B.n1041 B.n31 163.367
R999 B.n1037 B.n31 163.367
R1000 B.n1037 B.n33 163.367
R1001 B.n1033 B.n33 163.367
R1002 B.n1033 B.n38 163.367
R1003 B.n1029 B.n38 163.367
R1004 B.n1029 B.n40 163.367
R1005 B.n1025 B.n40 163.367
R1006 B.n1025 B.n45 163.367
R1007 B.n1021 B.n45 163.367
R1008 B.n1021 B.n47 163.367
R1009 B.n1017 B.n47 163.367
R1010 B.n1017 B.n52 163.367
R1011 B.n1013 B.n52 163.367
R1012 B.n1013 B.n54 163.367
R1013 B.n1009 B.n54 163.367
R1014 B.n1009 B.n59 163.367
R1015 B.n1005 B.n59 163.367
R1016 B.n1005 B.n61 163.367
R1017 B.n1001 B.n61 163.367
R1018 B.n1001 B.n66 163.367
R1019 B.n997 B.n66 163.367
R1020 B.n997 B.n68 163.367
R1021 B.n993 B.n68 163.367
R1022 B.n993 B.n73 163.367
R1023 B.n989 B.n73 163.367
R1024 B.n77 B.n75 71.676
R1025 B.n150 B.n78 71.676
R1026 B.n154 B.n79 71.676
R1027 B.n158 B.n80 71.676
R1028 B.n162 B.n81 71.676
R1029 B.n166 B.n82 71.676
R1030 B.n170 B.n83 71.676
R1031 B.n174 B.n84 71.676
R1032 B.n178 B.n85 71.676
R1033 B.n182 B.n86 71.676
R1034 B.n186 B.n87 71.676
R1035 B.n190 B.n88 71.676
R1036 B.n194 B.n89 71.676
R1037 B.n198 B.n90 71.676
R1038 B.n202 B.n91 71.676
R1039 B.n206 B.n92 71.676
R1040 B.n210 B.n93 71.676
R1041 B.n214 B.n94 71.676
R1042 B.n218 B.n95 71.676
R1043 B.n222 B.n96 71.676
R1044 B.n226 B.n97 71.676
R1045 B.n230 B.n98 71.676
R1046 B.n234 B.n99 71.676
R1047 B.n238 B.n100 71.676
R1048 B.n242 B.n101 71.676
R1049 B.n246 B.n102 71.676
R1050 B.n250 B.n103 71.676
R1051 B.n254 B.n104 71.676
R1052 B.n258 B.n105 71.676
R1053 B.n262 B.n106 71.676
R1054 B.n266 B.n107 71.676
R1055 B.n270 B.n108 71.676
R1056 B.n274 B.n109 71.676
R1057 B.n278 B.n110 71.676
R1058 B.n282 B.n111 71.676
R1059 B.n286 B.n112 71.676
R1060 B.n290 B.n113 71.676
R1061 B.n294 B.n114 71.676
R1062 B.n298 B.n115 71.676
R1063 B.n302 B.n116 71.676
R1064 B.n306 B.n117 71.676
R1065 B.n310 B.n118 71.676
R1066 B.n314 B.n119 71.676
R1067 B.n318 B.n120 71.676
R1068 B.n322 B.n121 71.676
R1069 B.n326 B.n122 71.676
R1070 B.n330 B.n123 71.676
R1071 B.n334 B.n124 71.676
R1072 B.n338 B.n125 71.676
R1073 B.n342 B.n126 71.676
R1074 B.n346 B.n127 71.676
R1075 B.n350 B.n128 71.676
R1076 B.n354 B.n129 71.676
R1077 B.n358 B.n130 71.676
R1078 B.n362 B.n131 71.676
R1079 B.n366 B.n132 71.676
R1080 B.n370 B.n133 71.676
R1081 B.n374 B.n134 71.676
R1082 B.n378 B.n135 71.676
R1083 B.n382 B.n136 71.676
R1084 B.n386 B.n137 71.676
R1085 B.n390 B.n138 71.676
R1086 B.n394 B.n139 71.676
R1087 B.n398 B.n140 71.676
R1088 B.n986 B.n141 71.676
R1089 B.n986 B.n985 71.676
R1090 B.n400 B.n140 71.676
R1091 B.n397 B.n139 71.676
R1092 B.n393 B.n138 71.676
R1093 B.n389 B.n137 71.676
R1094 B.n385 B.n136 71.676
R1095 B.n381 B.n135 71.676
R1096 B.n377 B.n134 71.676
R1097 B.n373 B.n133 71.676
R1098 B.n369 B.n132 71.676
R1099 B.n365 B.n131 71.676
R1100 B.n361 B.n130 71.676
R1101 B.n357 B.n129 71.676
R1102 B.n353 B.n128 71.676
R1103 B.n349 B.n127 71.676
R1104 B.n345 B.n126 71.676
R1105 B.n341 B.n125 71.676
R1106 B.n337 B.n124 71.676
R1107 B.n333 B.n123 71.676
R1108 B.n329 B.n122 71.676
R1109 B.n325 B.n121 71.676
R1110 B.n321 B.n120 71.676
R1111 B.n317 B.n119 71.676
R1112 B.n313 B.n118 71.676
R1113 B.n309 B.n117 71.676
R1114 B.n305 B.n116 71.676
R1115 B.n301 B.n115 71.676
R1116 B.n297 B.n114 71.676
R1117 B.n293 B.n113 71.676
R1118 B.n289 B.n112 71.676
R1119 B.n285 B.n111 71.676
R1120 B.n281 B.n110 71.676
R1121 B.n277 B.n109 71.676
R1122 B.n273 B.n108 71.676
R1123 B.n269 B.n107 71.676
R1124 B.n265 B.n106 71.676
R1125 B.n261 B.n105 71.676
R1126 B.n257 B.n104 71.676
R1127 B.n253 B.n103 71.676
R1128 B.n249 B.n102 71.676
R1129 B.n245 B.n101 71.676
R1130 B.n241 B.n100 71.676
R1131 B.n237 B.n99 71.676
R1132 B.n233 B.n98 71.676
R1133 B.n229 B.n97 71.676
R1134 B.n225 B.n96 71.676
R1135 B.n221 B.n95 71.676
R1136 B.n217 B.n94 71.676
R1137 B.n213 B.n93 71.676
R1138 B.n209 B.n92 71.676
R1139 B.n205 B.n91 71.676
R1140 B.n201 B.n90 71.676
R1141 B.n197 B.n89 71.676
R1142 B.n193 B.n88 71.676
R1143 B.n189 B.n87 71.676
R1144 B.n185 B.n86 71.676
R1145 B.n181 B.n85 71.676
R1146 B.n177 B.n84 71.676
R1147 B.n173 B.n83 71.676
R1148 B.n169 B.n82 71.676
R1149 B.n165 B.n81 71.676
R1150 B.n161 B.n80 71.676
R1151 B.n157 B.n79 71.676
R1152 B.n153 B.n78 71.676
R1153 B.n149 B.n77 71.676
R1154 B.n549 B.n479 71.676
R1155 B.n553 B.n552 71.676
R1156 B.n558 B.n557 71.676
R1157 B.n561 B.n560 71.676
R1158 B.n566 B.n565 71.676
R1159 B.n569 B.n568 71.676
R1160 B.n574 B.n573 71.676
R1161 B.n577 B.n576 71.676
R1162 B.n582 B.n581 71.676
R1163 B.n585 B.n584 71.676
R1164 B.n590 B.n589 71.676
R1165 B.n593 B.n592 71.676
R1166 B.n598 B.n597 71.676
R1167 B.n601 B.n600 71.676
R1168 B.n606 B.n605 71.676
R1169 B.n609 B.n608 71.676
R1170 B.n614 B.n613 71.676
R1171 B.n617 B.n616 71.676
R1172 B.n622 B.n621 71.676
R1173 B.n625 B.n624 71.676
R1174 B.n630 B.n629 71.676
R1175 B.n633 B.n632 71.676
R1176 B.n638 B.n637 71.676
R1177 B.n641 B.n640 71.676
R1178 B.n646 B.n645 71.676
R1179 B.n649 B.n648 71.676
R1180 B.n654 B.n653 71.676
R1181 B.n657 B.n656 71.676
R1182 B.n662 B.n661 71.676
R1183 B.n665 B.n664 71.676
R1184 B.n671 B.n670 71.676
R1185 B.n674 B.n673 71.676
R1186 B.n679 B.n678 71.676
R1187 B.n682 B.n681 71.676
R1188 B.n690 B.n689 71.676
R1189 B.n693 B.n692 71.676
R1190 B.n698 B.n697 71.676
R1191 B.n701 B.n700 71.676
R1192 B.n706 B.n705 71.676
R1193 B.n709 B.n708 71.676
R1194 B.n714 B.n713 71.676
R1195 B.n717 B.n716 71.676
R1196 B.n722 B.n721 71.676
R1197 B.n725 B.n724 71.676
R1198 B.n730 B.n729 71.676
R1199 B.n733 B.n732 71.676
R1200 B.n738 B.n737 71.676
R1201 B.n741 B.n740 71.676
R1202 B.n746 B.n745 71.676
R1203 B.n749 B.n748 71.676
R1204 B.n754 B.n753 71.676
R1205 B.n757 B.n756 71.676
R1206 B.n762 B.n761 71.676
R1207 B.n765 B.n764 71.676
R1208 B.n770 B.n769 71.676
R1209 B.n773 B.n772 71.676
R1210 B.n778 B.n777 71.676
R1211 B.n781 B.n780 71.676
R1212 B.n786 B.n785 71.676
R1213 B.n789 B.n788 71.676
R1214 B.n794 B.n793 71.676
R1215 B.n797 B.n796 71.676
R1216 B.n802 B.n801 71.676
R1217 B.n805 B.n804 71.676
R1218 B.n550 B.n549 71.676
R1219 B.n552 B.n546 71.676
R1220 B.n559 B.n558 71.676
R1221 B.n560 B.n544 71.676
R1222 B.n567 B.n566 71.676
R1223 B.n568 B.n542 71.676
R1224 B.n575 B.n574 71.676
R1225 B.n576 B.n540 71.676
R1226 B.n583 B.n582 71.676
R1227 B.n584 B.n538 71.676
R1228 B.n591 B.n590 71.676
R1229 B.n592 B.n536 71.676
R1230 B.n599 B.n598 71.676
R1231 B.n600 B.n534 71.676
R1232 B.n607 B.n606 71.676
R1233 B.n608 B.n532 71.676
R1234 B.n615 B.n614 71.676
R1235 B.n616 B.n530 71.676
R1236 B.n623 B.n622 71.676
R1237 B.n624 B.n528 71.676
R1238 B.n631 B.n630 71.676
R1239 B.n632 B.n526 71.676
R1240 B.n639 B.n638 71.676
R1241 B.n640 B.n524 71.676
R1242 B.n647 B.n646 71.676
R1243 B.n648 B.n522 71.676
R1244 B.n655 B.n654 71.676
R1245 B.n656 B.n520 71.676
R1246 B.n663 B.n662 71.676
R1247 B.n664 B.n516 71.676
R1248 B.n672 B.n671 71.676
R1249 B.n673 B.n514 71.676
R1250 B.n680 B.n679 71.676
R1251 B.n681 B.n512 71.676
R1252 B.n691 B.n690 71.676
R1253 B.n692 B.n510 71.676
R1254 B.n699 B.n698 71.676
R1255 B.n700 B.n508 71.676
R1256 B.n707 B.n706 71.676
R1257 B.n708 B.n506 71.676
R1258 B.n715 B.n714 71.676
R1259 B.n716 B.n504 71.676
R1260 B.n723 B.n722 71.676
R1261 B.n724 B.n502 71.676
R1262 B.n731 B.n730 71.676
R1263 B.n732 B.n500 71.676
R1264 B.n739 B.n738 71.676
R1265 B.n740 B.n498 71.676
R1266 B.n747 B.n746 71.676
R1267 B.n748 B.n496 71.676
R1268 B.n755 B.n754 71.676
R1269 B.n756 B.n494 71.676
R1270 B.n763 B.n762 71.676
R1271 B.n764 B.n492 71.676
R1272 B.n771 B.n770 71.676
R1273 B.n772 B.n490 71.676
R1274 B.n779 B.n778 71.676
R1275 B.n780 B.n488 71.676
R1276 B.n787 B.n786 71.676
R1277 B.n788 B.n486 71.676
R1278 B.n795 B.n794 71.676
R1279 B.n796 B.n484 71.676
R1280 B.n803 B.n802 71.676
R1281 B.n806 B.n805 71.676
R1282 B.n1071 B.n1070 71.676
R1283 B.n1071 B.n2 71.676
R1284 B.n811 B.n480 65.8744
R1285 B.n988 B.n987 65.8744
R1286 B.n147 B.n146 59.5399
R1287 B.n144 B.n143 59.5399
R1288 B.n687 B.n686 59.5399
R1289 B.n667 B.n518 59.5399
R1290 B.n146 B.n145 43.055
R1291 B.n143 B.n142 43.055
R1292 B.n686 B.n685 43.055
R1293 B.n518 B.n517 43.055
R1294 B.n813 B.n478 33.5615
R1295 B.n809 B.n808 33.5615
R1296 B.n984 B.n983 33.5615
R1297 B.n990 B.n74 33.5615
R1298 B.n811 B.n476 31.7695
R1299 B.n817 B.n476 31.7695
R1300 B.n817 B.n472 31.7695
R1301 B.n823 B.n472 31.7695
R1302 B.n823 B.n468 31.7695
R1303 B.n829 B.n468 31.7695
R1304 B.n835 B.n464 31.7695
R1305 B.n835 B.n460 31.7695
R1306 B.n841 B.n460 31.7695
R1307 B.n841 B.n456 31.7695
R1308 B.n847 B.n456 31.7695
R1309 B.n847 B.n452 31.7695
R1310 B.n853 B.n452 31.7695
R1311 B.n853 B.n448 31.7695
R1312 B.n859 B.n448 31.7695
R1313 B.n865 B.n444 31.7695
R1314 B.n865 B.n440 31.7695
R1315 B.n871 B.n440 31.7695
R1316 B.n871 B.n436 31.7695
R1317 B.n877 B.n436 31.7695
R1318 B.n883 B.n432 31.7695
R1319 B.n883 B.n428 31.7695
R1320 B.n889 B.n428 31.7695
R1321 B.n889 B.n424 31.7695
R1322 B.n896 B.n424 31.7695
R1323 B.n896 B.n895 31.7695
R1324 B.n902 B.n417 31.7695
R1325 B.n908 B.n417 31.7695
R1326 B.n908 B.n412 31.7695
R1327 B.n914 B.n412 31.7695
R1328 B.n914 B.n413 31.7695
R1329 B.n921 B.n405 31.7695
R1330 B.n927 B.n405 31.7695
R1331 B.n927 B.n4 31.7695
R1332 B.n1069 B.n4 31.7695
R1333 B.n1069 B.n1068 31.7695
R1334 B.n1068 B.n1067 31.7695
R1335 B.n1067 B.n8 31.7695
R1336 B.n12 B.n8 31.7695
R1337 B.n1060 B.n12 31.7695
R1338 B.n1059 B.n1058 31.7695
R1339 B.n1058 B.n16 31.7695
R1340 B.n1052 B.n16 31.7695
R1341 B.n1052 B.n1051 31.7695
R1342 B.n1051 B.n1050 31.7695
R1343 B.n1044 B.n26 31.7695
R1344 B.n1044 B.n1043 31.7695
R1345 B.n1043 B.n1042 31.7695
R1346 B.n1042 B.n30 31.7695
R1347 B.n1036 B.n30 31.7695
R1348 B.n1036 B.n1035 31.7695
R1349 B.n1034 B.n37 31.7695
R1350 B.n1028 B.n37 31.7695
R1351 B.n1028 B.n1027 31.7695
R1352 B.n1027 B.n1026 31.7695
R1353 B.n1026 B.n44 31.7695
R1354 B.n1020 B.n1019 31.7695
R1355 B.n1019 B.n1018 31.7695
R1356 B.n1018 B.n51 31.7695
R1357 B.n1012 B.n51 31.7695
R1358 B.n1012 B.n1011 31.7695
R1359 B.n1011 B.n1010 31.7695
R1360 B.n1010 B.n58 31.7695
R1361 B.n1004 B.n58 31.7695
R1362 B.n1004 B.n1003 31.7695
R1363 B.n1002 B.n65 31.7695
R1364 B.n996 B.n65 31.7695
R1365 B.n996 B.n995 31.7695
R1366 B.n995 B.n994 31.7695
R1367 B.n994 B.n72 31.7695
R1368 B.n988 B.n72 31.7695
R1369 B.t3 B.n444 30.3679
R1370 B.t6 B.n44 30.3679
R1371 B.n902 B.t7 28.4991
R1372 B.n1050 B.t1 28.4991
R1373 B.t9 B.n464 21.9585
R1374 B.n1003 B.t13 21.9585
R1375 B.n413 B.t0 20.0897
R1376 B.t4 B.n1059 20.0897
R1377 B.n877 B.t5 18.2209
R1378 B.t2 B.n1034 18.2209
R1379 B B.n1072 18.0485
R1380 B.t5 B.n432 13.549
R1381 B.n1035 B.t2 13.549
R1382 B.n921 B.t0 11.6803
R1383 B.n1060 B.t4 11.6803
R1384 B.n814 B.n813 10.6151
R1385 B.n815 B.n814 10.6151
R1386 B.n815 B.n470 10.6151
R1387 B.n825 B.n470 10.6151
R1388 B.n826 B.n825 10.6151
R1389 B.n827 B.n826 10.6151
R1390 B.n827 B.n462 10.6151
R1391 B.n837 B.n462 10.6151
R1392 B.n838 B.n837 10.6151
R1393 B.n839 B.n838 10.6151
R1394 B.n839 B.n454 10.6151
R1395 B.n849 B.n454 10.6151
R1396 B.n850 B.n849 10.6151
R1397 B.n851 B.n850 10.6151
R1398 B.n851 B.n446 10.6151
R1399 B.n861 B.n446 10.6151
R1400 B.n862 B.n861 10.6151
R1401 B.n863 B.n862 10.6151
R1402 B.n863 B.n438 10.6151
R1403 B.n873 B.n438 10.6151
R1404 B.n874 B.n873 10.6151
R1405 B.n875 B.n874 10.6151
R1406 B.n875 B.n430 10.6151
R1407 B.n885 B.n430 10.6151
R1408 B.n886 B.n885 10.6151
R1409 B.n887 B.n886 10.6151
R1410 B.n887 B.n422 10.6151
R1411 B.n898 B.n422 10.6151
R1412 B.n899 B.n898 10.6151
R1413 B.n900 B.n899 10.6151
R1414 B.n900 B.n415 10.6151
R1415 B.n910 B.n415 10.6151
R1416 B.n911 B.n910 10.6151
R1417 B.n912 B.n911 10.6151
R1418 B.n912 B.n407 10.6151
R1419 B.n923 B.n407 10.6151
R1420 B.n924 B.n923 10.6151
R1421 B.n925 B.n924 10.6151
R1422 B.n925 B.n0 10.6151
R1423 B.n548 B.n478 10.6151
R1424 B.n548 B.n547 10.6151
R1425 B.n554 B.n547 10.6151
R1426 B.n555 B.n554 10.6151
R1427 B.n556 B.n555 10.6151
R1428 B.n556 B.n545 10.6151
R1429 B.n562 B.n545 10.6151
R1430 B.n563 B.n562 10.6151
R1431 B.n564 B.n563 10.6151
R1432 B.n564 B.n543 10.6151
R1433 B.n570 B.n543 10.6151
R1434 B.n571 B.n570 10.6151
R1435 B.n572 B.n571 10.6151
R1436 B.n572 B.n541 10.6151
R1437 B.n578 B.n541 10.6151
R1438 B.n579 B.n578 10.6151
R1439 B.n580 B.n579 10.6151
R1440 B.n580 B.n539 10.6151
R1441 B.n586 B.n539 10.6151
R1442 B.n587 B.n586 10.6151
R1443 B.n588 B.n587 10.6151
R1444 B.n588 B.n537 10.6151
R1445 B.n594 B.n537 10.6151
R1446 B.n595 B.n594 10.6151
R1447 B.n596 B.n595 10.6151
R1448 B.n596 B.n535 10.6151
R1449 B.n602 B.n535 10.6151
R1450 B.n603 B.n602 10.6151
R1451 B.n604 B.n603 10.6151
R1452 B.n604 B.n533 10.6151
R1453 B.n610 B.n533 10.6151
R1454 B.n611 B.n610 10.6151
R1455 B.n612 B.n611 10.6151
R1456 B.n612 B.n531 10.6151
R1457 B.n618 B.n531 10.6151
R1458 B.n619 B.n618 10.6151
R1459 B.n620 B.n619 10.6151
R1460 B.n620 B.n529 10.6151
R1461 B.n626 B.n529 10.6151
R1462 B.n627 B.n626 10.6151
R1463 B.n628 B.n627 10.6151
R1464 B.n628 B.n527 10.6151
R1465 B.n634 B.n527 10.6151
R1466 B.n635 B.n634 10.6151
R1467 B.n636 B.n635 10.6151
R1468 B.n636 B.n525 10.6151
R1469 B.n642 B.n525 10.6151
R1470 B.n643 B.n642 10.6151
R1471 B.n644 B.n643 10.6151
R1472 B.n644 B.n523 10.6151
R1473 B.n650 B.n523 10.6151
R1474 B.n651 B.n650 10.6151
R1475 B.n652 B.n651 10.6151
R1476 B.n652 B.n521 10.6151
R1477 B.n658 B.n521 10.6151
R1478 B.n659 B.n658 10.6151
R1479 B.n660 B.n659 10.6151
R1480 B.n660 B.n519 10.6151
R1481 B.n666 B.n519 10.6151
R1482 B.n669 B.n668 10.6151
R1483 B.n669 B.n515 10.6151
R1484 B.n675 B.n515 10.6151
R1485 B.n676 B.n675 10.6151
R1486 B.n677 B.n676 10.6151
R1487 B.n677 B.n513 10.6151
R1488 B.n683 B.n513 10.6151
R1489 B.n684 B.n683 10.6151
R1490 B.n688 B.n684 10.6151
R1491 B.n694 B.n511 10.6151
R1492 B.n695 B.n694 10.6151
R1493 B.n696 B.n695 10.6151
R1494 B.n696 B.n509 10.6151
R1495 B.n702 B.n509 10.6151
R1496 B.n703 B.n702 10.6151
R1497 B.n704 B.n703 10.6151
R1498 B.n704 B.n507 10.6151
R1499 B.n710 B.n507 10.6151
R1500 B.n711 B.n710 10.6151
R1501 B.n712 B.n711 10.6151
R1502 B.n712 B.n505 10.6151
R1503 B.n718 B.n505 10.6151
R1504 B.n719 B.n718 10.6151
R1505 B.n720 B.n719 10.6151
R1506 B.n720 B.n503 10.6151
R1507 B.n726 B.n503 10.6151
R1508 B.n727 B.n726 10.6151
R1509 B.n728 B.n727 10.6151
R1510 B.n728 B.n501 10.6151
R1511 B.n734 B.n501 10.6151
R1512 B.n735 B.n734 10.6151
R1513 B.n736 B.n735 10.6151
R1514 B.n736 B.n499 10.6151
R1515 B.n742 B.n499 10.6151
R1516 B.n743 B.n742 10.6151
R1517 B.n744 B.n743 10.6151
R1518 B.n744 B.n497 10.6151
R1519 B.n750 B.n497 10.6151
R1520 B.n751 B.n750 10.6151
R1521 B.n752 B.n751 10.6151
R1522 B.n752 B.n495 10.6151
R1523 B.n758 B.n495 10.6151
R1524 B.n759 B.n758 10.6151
R1525 B.n760 B.n759 10.6151
R1526 B.n760 B.n493 10.6151
R1527 B.n766 B.n493 10.6151
R1528 B.n767 B.n766 10.6151
R1529 B.n768 B.n767 10.6151
R1530 B.n768 B.n491 10.6151
R1531 B.n774 B.n491 10.6151
R1532 B.n775 B.n774 10.6151
R1533 B.n776 B.n775 10.6151
R1534 B.n776 B.n489 10.6151
R1535 B.n782 B.n489 10.6151
R1536 B.n783 B.n782 10.6151
R1537 B.n784 B.n783 10.6151
R1538 B.n784 B.n487 10.6151
R1539 B.n790 B.n487 10.6151
R1540 B.n791 B.n790 10.6151
R1541 B.n792 B.n791 10.6151
R1542 B.n792 B.n485 10.6151
R1543 B.n798 B.n485 10.6151
R1544 B.n799 B.n798 10.6151
R1545 B.n800 B.n799 10.6151
R1546 B.n800 B.n483 10.6151
R1547 B.n483 B.n482 10.6151
R1548 B.n807 B.n482 10.6151
R1549 B.n808 B.n807 10.6151
R1550 B.n809 B.n474 10.6151
R1551 B.n819 B.n474 10.6151
R1552 B.n820 B.n819 10.6151
R1553 B.n821 B.n820 10.6151
R1554 B.n821 B.n466 10.6151
R1555 B.n831 B.n466 10.6151
R1556 B.n832 B.n831 10.6151
R1557 B.n833 B.n832 10.6151
R1558 B.n833 B.n458 10.6151
R1559 B.n843 B.n458 10.6151
R1560 B.n844 B.n843 10.6151
R1561 B.n845 B.n844 10.6151
R1562 B.n845 B.n450 10.6151
R1563 B.n855 B.n450 10.6151
R1564 B.n856 B.n855 10.6151
R1565 B.n857 B.n856 10.6151
R1566 B.n857 B.n442 10.6151
R1567 B.n867 B.n442 10.6151
R1568 B.n868 B.n867 10.6151
R1569 B.n869 B.n868 10.6151
R1570 B.n869 B.n434 10.6151
R1571 B.n879 B.n434 10.6151
R1572 B.n880 B.n879 10.6151
R1573 B.n881 B.n880 10.6151
R1574 B.n881 B.n426 10.6151
R1575 B.n891 B.n426 10.6151
R1576 B.n892 B.n891 10.6151
R1577 B.n893 B.n892 10.6151
R1578 B.n893 B.n419 10.6151
R1579 B.n904 B.n419 10.6151
R1580 B.n905 B.n904 10.6151
R1581 B.n906 B.n905 10.6151
R1582 B.n906 B.n410 10.6151
R1583 B.n916 B.n410 10.6151
R1584 B.n917 B.n916 10.6151
R1585 B.n919 B.n917 10.6151
R1586 B.n919 B.n918 10.6151
R1587 B.n918 B.n403 10.6151
R1588 B.n930 B.n403 10.6151
R1589 B.n931 B.n930 10.6151
R1590 B.n932 B.n931 10.6151
R1591 B.n933 B.n932 10.6151
R1592 B.n934 B.n933 10.6151
R1593 B.n937 B.n934 10.6151
R1594 B.n938 B.n937 10.6151
R1595 B.n939 B.n938 10.6151
R1596 B.n940 B.n939 10.6151
R1597 B.n942 B.n940 10.6151
R1598 B.n943 B.n942 10.6151
R1599 B.n944 B.n943 10.6151
R1600 B.n945 B.n944 10.6151
R1601 B.n947 B.n945 10.6151
R1602 B.n948 B.n947 10.6151
R1603 B.n949 B.n948 10.6151
R1604 B.n950 B.n949 10.6151
R1605 B.n952 B.n950 10.6151
R1606 B.n953 B.n952 10.6151
R1607 B.n954 B.n953 10.6151
R1608 B.n955 B.n954 10.6151
R1609 B.n957 B.n955 10.6151
R1610 B.n958 B.n957 10.6151
R1611 B.n959 B.n958 10.6151
R1612 B.n960 B.n959 10.6151
R1613 B.n962 B.n960 10.6151
R1614 B.n963 B.n962 10.6151
R1615 B.n964 B.n963 10.6151
R1616 B.n965 B.n964 10.6151
R1617 B.n967 B.n965 10.6151
R1618 B.n968 B.n967 10.6151
R1619 B.n969 B.n968 10.6151
R1620 B.n970 B.n969 10.6151
R1621 B.n972 B.n970 10.6151
R1622 B.n973 B.n972 10.6151
R1623 B.n974 B.n973 10.6151
R1624 B.n975 B.n974 10.6151
R1625 B.n977 B.n975 10.6151
R1626 B.n978 B.n977 10.6151
R1627 B.n979 B.n978 10.6151
R1628 B.n980 B.n979 10.6151
R1629 B.n982 B.n980 10.6151
R1630 B.n983 B.n982 10.6151
R1631 B.n1064 B.n1 10.6151
R1632 B.n1064 B.n1063 10.6151
R1633 B.n1063 B.n1062 10.6151
R1634 B.n1062 B.n10 10.6151
R1635 B.n1056 B.n10 10.6151
R1636 B.n1056 B.n1055 10.6151
R1637 B.n1055 B.n1054 10.6151
R1638 B.n1054 B.n18 10.6151
R1639 B.n1048 B.n18 10.6151
R1640 B.n1048 B.n1047 10.6151
R1641 B.n1047 B.n1046 10.6151
R1642 B.n1046 B.n24 10.6151
R1643 B.n1040 B.n24 10.6151
R1644 B.n1040 B.n1039 10.6151
R1645 B.n1039 B.n1038 10.6151
R1646 B.n1038 B.n32 10.6151
R1647 B.n1032 B.n32 10.6151
R1648 B.n1032 B.n1031 10.6151
R1649 B.n1031 B.n1030 10.6151
R1650 B.n1030 B.n39 10.6151
R1651 B.n1024 B.n39 10.6151
R1652 B.n1024 B.n1023 10.6151
R1653 B.n1023 B.n1022 10.6151
R1654 B.n1022 B.n46 10.6151
R1655 B.n1016 B.n46 10.6151
R1656 B.n1016 B.n1015 10.6151
R1657 B.n1015 B.n1014 10.6151
R1658 B.n1014 B.n53 10.6151
R1659 B.n1008 B.n53 10.6151
R1660 B.n1008 B.n1007 10.6151
R1661 B.n1007 B.n1006 10.6151
R1662 B.n1006 B.n60 10.6151
R1663 B.n1000 B.n60 10.6151
R1664 B.n1000 B.n999 10.6151
R1665 B.n999 B.n998 10.6151
R1666 B.n998 B.n67 10.6151
R1667 B.n992 B.n67 10.6151
R1668 B.n992 B.n991 10.6151
R1669 B.n991 B.n990 10.6151
R1670 B.n148 B.n74 10.6151
R1671 B.n151 B.n148 10.6151
R1672 B.n152 B.n151 10.6151
R1673 B.n155 B.n152 10.6151
R1674 B.n156 B.n155 10.6151
R1675 B.n159 B.n156 10.6151
R1676 B.n160 B.n159 10.6151
R1677 B.n163 B.n160 10.6151
R1678 B.n164 B.n163 10.6151
R1679 B.n167 B.n164 10.6151
R1680 B.n168 B.n167 10.6151
R1681 B.n171 B.n168 10.6151
R1682 B.n172 B.n171 10.6151
R1683 B.n175 B.n172 10.6151
R1684 B.n176 B.n175 10.6151
R1685 B.n179 B.n176 10.6151
R1686 B.n180 B.n179 10.6151
R1687 B.n183 B.n180 10.6151
R1688 B.n184 B.n183 10.6151
R1689 B.n187 B.n184 10.6151
R1690 B.n188 B.n187 10.6151
R1691 B.n191 B.n188 10.6151
R1692 B.n192 B.n191 10.6151
R1693 B.n195 B.n192 10.6151
R1694 B.n196 B.n195 10.6151
R1695 B.n199 B.n196 10.6151
R1696 B.n200 B.n199 10.6151
R1697 B.n203 B.n200 10.6151
R1698 B.n204 B.n203 10.6151
R1699 B.n207 B.n204 10.6151
R1700 B.n208 B.n207 10.6151
R1701 B.n211 B.n208 10.6151
R1702 B.n212 B.n211 10.6151
R1703 B.n215 B.n212 10.6151
R1704 B.n216 B.n215 10.6151
R1705 B.n219 B.n216 10.6151
R1706 B.n220 B.n219 10.6151
R1707 B.n223 B.n220 10.6151
R1708 B.n224 B.n223 10.6151
R1709 B.n227 B.n224 10.6151
R1710 B.n228 B.n227 10.6151
R1711 B.n231 B.n228 10.6151
R1712 B.n232 B.n231 10.6151
R1713 B.n235 B.n232 10.6151
R1714 B.n236 B.n235 10.6151
R1715 B.n239 B.n236 10.6151
R1716 B.n240 B.n239 10.6151
R1717 B.n243 B.n240 10.6151
R1718 B.n244 B.n243 10.6151
R1719 B.n247 B.n244 10.6151
R1720 B.n248 B.n247 10.6151
R1721 B.n251 B.n248 10.6151
R1722 B.n252 B.n251 10.6151
R1723 B.n255 B.n252 10.6151
R1724 B.n256 B.n255 10.6151
R1725 B.n259 B.n256 10.6151
R1726 B.n260 B.n259 10.6151
R1727 B.n263 B.n260 10.6151
R1728 B.n264 B.n263 10.6151
R1729 B.n268 B.n267 10.6151
R1730 B.n271 B.n268 10.6151
R1731 B.n272 B.n271 10.6151
R1732 B.n275 B.n272 10.6151
R1733 B.n276 B.n275 10.6151
R1734 B.n279 B.n276 10.6151
R1735 B.n280 B.n279 10.6151
R1736 B.n283 B.n280 10.6151
R1737 B.n284 B.n283 10.6151
R1738 B.n288 B.n287 10.6151
R1739 B.n291 B.n288 10.6151
R1740 B.n292 B.n291 10.6151
R1741 B.n295 B.n292 10.6151
R1742 B.n296 B.n295 10.6151
R1743 B.n299 B.n296 10.6151
R1744 B.n300 B.n299 10.6151
R1745 B.n303 B.n300 10.6151
R1746 B.n304 B.n303 10.6151
R1747 B.n307 B.n304 10.6151
R1748 B.n308 B.n307 10.6151
R1749 B.n311 B.n308 10.6151
R1750 B.n312 B.n311 10.6151
R1751 B.n315 B.n312 10.6151
R1752 B.n316 B.n315 10.6151
R1753 B.n319 B.n316 10.6151
R1754 B.n320 B.n319 10.6151
R1755 B.n323 B.n320 10.6151
R1756 B.n324 B.n323 10.6151
R1757 B.n327 B.n324 10.6151
R1758 B.n328 B.n327 10.6151
R1759 B.n331 B.n328 10.6151
R1760 B.n332 B.n331 10.6151
R1761 B.n335 B.n332 10.6151
R1762 B.n336 B.n335 10.6151
R1763 B.n339 B.n336 10.6151
R1764 B.n340 B.n339 10.6151
R1765 B.n343 B.n340 10.6151
R1766 B.n344 B.n343 10.6151
R1767 B.n347 B.n344 10.6151
R1768 B.n348 B.n347 10.6151
R1769 B.n351 B.n348 10.6151
R1770 B.n352 B.n351 10.6151
R1771 B.n355 B.n352 10.6151
R1772 B.n356 B.n355 10.6151
R1773 B.n359 B.n356 10.6151
R1774 B.n360 B.n359 10.6151
R1775 B.n363 B.n360 10.6151
R1776 B.n364 B.n363 10.6151
R1777 B.n367 B.n364 10.6151
R1778 B.n368 B.n367 10.6151
R1779 B.n371 B.n368 10.6151
R1780 B.n372 B.n371 10.6151
R1781 B.n375 B.n372 10.6151
R1782 B.n376 B.n375 10.6151
R1783 B.n379 B.n376 10.6151
R1784 B.n380 B.n379 10.6151
R1785 B.n383 B.n380 10.6151
R1786 B.n384 B.n383 10.6151
R1787 B.n387 B.n384 10.6151
R1788 B.n388 B.n387 10.6151
R1789 B.n391 B.n388 10.6151
R1790 B.n392 B.n391 10.6151
R1791 B.n395 B.n392 10.6151
R1792 B.n396 B.n395 10.6151
R1793 B.n399 B.n396 10.6151
R1794 B.n401 B.n399 10.6151
R1795 B.n402 B.n401 10.6151
R1796 B.n984 B.n402 10.6151
R1797 B.n829 B.t9 9.8115
R1798 B.t13 B.n1002 9.8115
R1799 B.n667 B.n666 9.36635
R1800 B.n687 B.n511 9.36635
R1801 B.n264 B.n147 9.36635
R1802 B.n287 B.n144 9.36635
R1803 B.n1072 B.n0 8.11757
R1804 B.n1072 B.n1 8.11757
R1805 B.n895 B.t7 3.27083
R1806 B.n26 B.t1 3.27083
R1807 B.n859 B.t3 1.40207
R1808 B.n1020 B.t6 1.40207
R1809 B.n668 B.n667 1.24928
R1810 B.n688 B.n687 1.24928
R1811 B.n267 B.n147 1.24928
R1812 B.n284 B.n144 1.24928
R1813 VP.n13 VP.t3 267.307
R1814 VP.n7 VP.t2 232.968
R1815 VP.n40 VP.t7 232.968
R1816 VP.n47 VP.t4 232.968
R1817 VP.n55 VP.t1 232.968
R1818 VP.n29 VP.t0 232.968
R1819 VP.n21 VP.t5 232.968
R1820 VP.n14 VP.t6 232.968
R1821 VP.n31 VP.n7 181.852
R1822 VP.n56 VP.n55 181.852
R1823 VP.n30 VP.n29 181.852
R1824 VP.n15 VP.n12 161.3
R1825 VP.n17 VP.n16 161.3
R1826 VP.n18 VP.n11 161.3
R1827 VP.n20 VP.n19 161.3
R1828 VP.n22 VP.n10 161.3
R1829 VP.n24 VP.n23 161.3
R1830 VP.n25 VP.n9 161.3
R1831 VP.n27 VP.n26 161.3
R1832 VP.n28 VP.n8 161.3
R1833 VP.n54 VP.n0 161.3
R1834 VP.n53 VP.n52 161.3
R1835 VP.n51 VP.n1 161.3
R1836 VP.n50 VP.n49 161.3
R1837 VP.n48 VP.n2 161.3
R1838 VP.n46 VP.n45 161.3
R1839 VP.n44 VP.n3 161.3
R1840 VP.n43 VP.n42 161.3
R1841 VP.n41 VP.n4 161.3
R1842 VP.n39 VP.n38 161.3
R1843 VP.n37 VP.n5 161.3
R1844 VP.n36 VP.n35 161.3
R1845 VP.n34 VP.n6 161.3
R1846 VP.n33 VP.n32 161.3
R1847 VP.n42 VP.n3 56.5193
R1848 VP.n16 VP.n11 56.5193
R1849 VP.n31 VP.n30 52.2505
R1850 VP.n14 VP.n13 52.0405
R1851 VP.n35 VP.n5 43.4072
R1852 VP.n49 VP.n1 43.4072
R1853 VP.n23 VP.n9 43.4072
R1854 VP.n35 VP.n34 37.5796
R1855 VP.n53 VP.n1 37.5796
R1856 VP.n27 VP.n9 37.5796
R1857 VP.n34 VP.n33 24.4675
R1858 VP.n39 VP.n5 24.4675
R1859 VP.n42 VP.n41 24.4675
R1860 VP.n46 VP.n3 24.4675
R1861 VP.n49 VP.n48 24.4675
R1862 VP.n54 VP.n53 24.4675
R1863 VP.n28 VP.n27 24.4675
R1864 VP.n20 VP.n11 24.4675
R1865 VP.n23 VP.n22 24.4675
R1866 VP.n16 VP.n15 24.4675
R1867 VP.n41 VP.n40 17.6167
R1868 VP.n47 VP.n46 17.6167
R1869 VP.n21 VP.n20 17.6167
R1870 VP.n15 VP.n14 17.6167
R1871 VP.n13 VP.n12 12.2976
R1872 VP.n40 VP.n39 6.85126
R1873 VP.n48 VP.n47 6.85126
R1874 VP.n22 VP.n21 6.85126
R1875 VP.n33 VP.n7 3.91522
R1876 VP.n55 VP.n54 3.91522
R1877 VP.n29 VP.n28 3.91522
R1878 VP.n17 VP.n12 0.189894
R1879 VP.n18 VP.n17 0.189894
R1880 VP.n19 VP.n18 0.189894
R1881 VP.n19 VP.n10 0.189894
R1882 VP.n24 VP.n10 0.189894
R1883 VP.n25 VP.n24 0.189894
R1884 VP.n26 VP.n25 0.189894
R1885 VP.n26 VP.n8 0.189894
R1886 VP.n30 VP.n8 0.189894
R1887 VP.n32 VP.n31 0.189894
R1888 VP.n32 VP.n6 0.189894
R1889 VP.n36 VP.n6 0.189894
R1890 VP.n37 VP.n36 0.189894
R1891 VP.n38 VP.n37 0.189894
R1892 VP.n38 VP.n4 0.189894
R1893 VP.n43 VP.n4 0.189894
R1894 VP.n44 VP.n43 0.189894
R1895 VP.n45 VP.n44 0.189894
R1896 VP.n45 VP.n2 0.189894
R1897 VP.n50 VP.n2 0.189894
R1898 VP.n51 VP.n50 0.189894
R1899 VP.n52 VP.n51 0.189894
R1900 VP.n52 VP.n0 0.189894
R1901 VP.n56 VP.n0 0.189894
R1902 VP VP.n56 0.0516364
R1903 VTAIL.n818 VTAIL.n722 289.615
R1904 VTAIL.n98 VTAIL.n2 289.615
R1905 VTAIL.n200 VTAIL.n104 289.615
R1906 VTAIL.n304 VTAIL.n208 289.615
R1907 VTAIL.n716 VTAIL.n620 289.615
R1908 VTAIL.n612 VTAIL.n516 289.615
R1909 VTAIL.n510 VTAIL.n414 289.615
R1910 VTAIL.n406 VTAIL.n310 289.615
R1911 VTAIL.n754 VTAIL.n753 185
R1912 VTAIL.n759 VTAIL.n758 185
R1913 VTAIL.n761 VTAIL.n760 185
R1914 VTAIL.n750 VTAIL.n749 185
R1915 VTAIL.n767 VTAIL.n766 185
R1916 VTAIL.n769 VTAIL.n768 185
R1917 VTAIL.n746 VTAIL.n745 185
R1918 VTAIL.n775 VTAIL.n774 185
R1919 VTAIL.n777 VTAIL.n776 185
R1920 VTAIL.n742 VTAIL.n741 185
R1921 VTAIL.n783 VTAIL.n782 185
R1922 VTAIL.n785 VTAIL.n784 185
R1923 VTAIL.n738 VTAIL.n737 185
R1924 VTAIL.n791 VTAIL.n790 185
R1925 VTAIL.n793 VTAIL.n792 185
R1926 VTAIL.n734 VTAIL.n733 185
R1927 VTAIL.n800 VTAIL.n799 185
R1928 VTAIL.n801 VTAIL.n732 185
R1929 VTAIL.n803 VTAIL.n802 185
R1930 VTAIL.n730 VTAIL.n729 185
R1931 VTAIL.n809 VTAIL.n808 185
R1932 VTAIL.n811 VTAIL.n810 185
R1933 VTAIL.n726 VTAIL.n725 185
R1934 VTAIL.n817 VTAIL.n816 185
R1935 VTAIL.n819 VTAIL.n818 185
R1936 VTAIL.n34 VTAIL.n33 185
R1937 VTAIL.n39 VTAIL.n38 185
R1938 VTAIL.n41 VTAIL.n40 185
R1939 VTAIL.n30 VTAIL.n29 185
R1940 VTAIL.n47 VTAIL.n46 185
R1941 VTAIL.n49 VTAIL.n48 185
R1942 VTAIL.n26 VTAIL.n25 185
R1943 VTAIL.n55 VTAIL.n54 185
R1944 VTAIL.n57 VTAIL.n56 185
R1945 VTAIL.n22 VTAIL.n21 185
R1946 VTAIL.n63 VTAIL.n62 185
R1947 VTAIL.n65 VTAIL.n64 185
R1948 VTAIL.n18 VTAIL.n17 185
R1949 VTAIL.n71 VTAIL.n70 185
R1950 VTAIL.n73 VTAIL.n72 185
R1951 VTAIL.n14 VTAIL.n13 185
R1952 VTAIL.n80 VTAIL.n79 185
R1953 VTAIL.n81 VTAIL.n12 185
R1954 VTAIL.n83 VTAIL.n82 185
R1955 VTAIL.n10 VTAIL.n9 185
R1956 VTAIL.n89 VTAIL.n88 185
R1957 VTAIL.n91 VTAIL.n90 185
R1958 VTAIL.n6 VTAIL.n5 185
R1959 VTAIL.n97 VTAIL.n96 185
R1960 VTAIL.n99 VTAIL.n98 185
R1961 VTAIL.n136 VTAIL.n135 185
R1962 VTAIL.n141 VTAIL.n140 185
R1963 VTAIL.n143 VTAIL.n142 185
R1964 VTAIL.n132 VTAIL.n131 185
R1965 VTAIL.n149 VTAIL.n148 185
R1966 VTAIL.n151 VTAIL.n150 185
R1967 VTAIL.n128 VTAIL.n127 185
R1968 VTAIL.n157 VTAIL.n156 185
R1969 VTAIL.n159 VTAIL.n158 185
R1970 VTAIL.n124 VTAIL.n123 185
R1971 VTAIL.n165 VTAIL.n164 185
R1972 VTAIL.n167 VTAIL.n166 185
R1973 VTAIL.n120 VTAIL.n119 185
R1974 VTAIL.n173 VTAIL.n172 185
R1975 VTAIL.n175 VTAIL.n174 185
R1976 VTAIL.n116 VTAIL.n115 185
R1977 VTAIL.n182 VTAIL.n181 185
R1978 VTAIL.n183 VTAIL.n114 185
R1979 VTAIL.n185 VTAIL.n184 185
R1980 VTAIL.n112 VTAIL.n111 185
R1981 VTAIL.n191 VTAIL.n190 185
R1982 VTAIL.n193 VTAIL.n192 185
R1983 VTAIL.n108 VTAIL.n107 185
R1984 VTAIL.n199 VTAIL.n198 185
R1985 VTAIL.n201 VTAIL.n200 185
R1986 VTAIL.n240 VTAIL.n239 185
R1987 VTAIL.n245 VTAIL.n244 185
R1988 VTAIL.n247 VTAIL.n246 185
R1989 VTAIL.n236 VTAIL.n235 185
R1990 VTAIL.n253 VTAIL.n252 185
R1991 VTAIL.n255 VTAIL.n254 185
R1992 VTAIL.n232 VTAIL.n231 185
R1993 VTAIL.n261 VTAIL.n260 185
R1994 VTAIL.n263 VTAIL.n262 185
R1995 VTAIL.n228 VTAIL.n227 185
R1996 VTAIL.n269 VTAIL.n268 185
R1997 VTAIL.n271 VTAIL.n270 185
R1998 VTAIL.n224 VTAIL.n223 185
R1999 VTAIL.n277 VTAIL.n276 185
R2000 VTAIL.n279 VTAIL.n278 185
R2001 VTAIL.n220 VTAIL.n219 185
R2002 VTAIL.n286 VTAIL.n285 185
R2003 VTAIL.n287 VTAIL.n218 185
R2004 VTAIL.n289 VTAIL.n288 185
R2005 VTAIL.n216 VTAIL.n215 185
R2006 VTAIL.n295 VTAIL.n294 185
R2007 VTAIL.n297 VTAIL.n296 185
R2008 VTAIL.n212 VTAIL.n211 185
R2009 VTAIL.n303 VTAIL.n302 185
R2010 VTAIL.n305 VTAIL.n304 185
R2011 VTAIL.n717 VTAIL.n716 185
R2012 VTAIL.n715 VTAIL.n714 185
R2013 VTAIL.n624 VTAIL.n623 185
R2014 VTAIL.n709 VTAIL.n708 185
R2015 VTAIL.n707 VTAIL.n706 185
R2016 VTAIL.n628 VTAIL.n627 185
R2017 VTAIL.n701 VTAIL.n700 185
R2018 VTAIL.n699 VTAIL.n630 185
R2019 VTAIL.n698 VTAIL.n697 185
R2020 VTAIL.n633 VTAIL.n631 185
R2021 VTAIL.n692 VTAIL.n691 185
R2022 VTAIL.n690 VTAIL.n689 185
R2023 VTAIL.n637 VTAIL.n636 185
R2024 VTAIL.n684 VTAIL.n683 185
R2025 VTAIL.n682 VTAIL.n681 185
R2026 VTAIL.n641 VTAIL.n640 185
R2027 VTAIL.n676 VTAIL.n675 185
R2028 VTAIL.n674 VTAIL.n673 185
R2029 VTAIL.n645 VTAIL.n644 185
R2030 VTAIL.n668 VTAIL.n667 185
R2031 VTAIL.n666 VTAIL.n665 185
R2032 VTAIL.n649 VTAIL.n648 185
R2033 VTAIL.n660 VTAIL.n659 185
R2034 VTAIL.n658 VTAIL.n657 185
R2035 VTAIL.n653 VTAIL.n652 185
R2036 VTAIL.n613 VTAIL.n612 185
R2037 VTAIL.n611 VTAIL.n610 185
R2038 VTAIL.n520 VTAIL.n519 185
R2039 VTAIL.n605 VTAIL.n604 185
R2040 VTAIL.n603 VTAIL.n602 185
R2041 VTAIL.n524 VTAIL.n523 185
R2042 VTAIL.n597 VTAIL.n596 185
R2043 VTAIL.n595 VTAIL.n526 185
R2044 VTAIL.n594 VTAIL.n593 185
R2045 VTAIL.n529 VTAIL.n527 185
R2046 VTAIL.n588 VTAIL.n587 185
R2047 VTAIL.n586 VTAIL.n585 185
R2048 VTAIL.n533 VTAIL.n532 185
R2049 VTAIL.n580 VTAIL.n579 185
R2050 VTAIL.n578 VTAIL.n577 185
R2051 VTAIL.n537 VTAIL.n536 185
R2052 VTAIL.n572 VTAIL.n571 185
R2053 VTAIL.n570 VTAIL.n569 185
R2054 VTAIL.n541 VTAIL.n540 185
R2055 VTAIL.n564 VTAIL.n563 185
R2056 VTAIL.n562 VTAIL.n561 185
R2057 VTAIL.n545 VTAIL.n544 185
R2058 VTAIL.n556 VTAIL.n555 185
R2059 VTAIL.n554 VTAIL.n553 185
R2060 VTAIL.n549 VTAIL.n548 185
R2061 VTAIL.n511 VTAIL.n510 185
R2062 VTAIL.n509 VTAIL.n508 185
R2063 VTAIL.n418 VTAIL.n417 185
R2064 VTAIL.n503 VTAIL.n502 185
R2065 VTAIL.n501 VTAIL.n500 185
R2066 VTAIL.n422 VTAIL.n421 185
R2067 VTAIL.n495 VTAIL.n494 185
R2068 VTAIL.n493 VTAIL.n424 185
R2069 VTAIL.n492 VTAIL.n491 185
R2070 VTAIL.n427 VTAIL.n425 185
R2071 VTAIL.n486 VTAIL.n485 185
R2072 VTAIL.n484 VTAIL.n483 185
R2073 VTAIL.n431 VTAIL.n430 185
R2074 VTAIL.n478 VTAIL.n477 185
R2075 VTAIL.n476 VTAIL.n475 185
R2076 VTAIL.n435 VTAIL.n434 185
R2077 VTAIL.n470 VTAIL.n469 185
R2078 VTAIL.n468 VTAIL.n467 185
R2079 VTAIL.n439 VTAIL.n438 185
R2080 VTAIL.n462 VTAIL.n461 185
R2081 VTAIL.n460 VTAIL.n459 185
R2082 VTAIL.n443 VTAIL.n442 185
R2083 VTAIL.n454 VTAIL.n453 185
R2084 VTAIL.n452 VTAIL.n451 185
R2085 VTAIL.n447 VTAIL.n446 185
R2086 VTAIL.n407 VTAIL.n406 185
R2087 VTAIL.n405 VTAIL.n404 185
R2088 VTAIL.n314 VTAIL.n313 185
R2089 VTAIL.n399 VTAIL.n398 185
R2090 VTAIL.n397 VTAIL.n396 185
R2091 VTAIL.n318 VTAIL.n317 185
R2092 VTAIL.n391 VTAIL.n390 185
R2093 VTAIL.n389 VTAIL.n320 185
R2094 VTAIL.n388 VTAIL.n387 185
R2095 VTAIL.n323 VTAIL.n321 185
R2096 VTAIL.n382 VTAIL.n381 185
R2097 VTAIL.n380 VTAIL.n379 185
R2098 VTAIL.n327 VTAIL.n326 185
R2099 VTAIL.n374 VTAIL.n373 185
R2100 VTAIL.n372 VTAIL.n371 185
R2101 VTAIL.n331 VTAIL.n330 185
R2102 VTAIL.n366 VTAIL.n365 185
R2103 VTAIL.n364 VTAIL.n363 185
R2104 VTAIL.n335 VTAIL.n334 185
R2105 VTAIL.n358 VTAIL.n357 185
R2106 VTAIL.n356 VTAIL.n355 185
R2107 VTAIL.n339 VTAIL.n338 185
R2108 VTAIL.n350 VTAIL.n349 185
R2109 VTAIL.n348 VTAIL.n347 185
R2110 VTAIL.n343 VTAIL.n342 185
R2111 VTAIL.n755 VTAIL.t6 147.659
R2112 VTAIL.n35 VTAIL.t5 147.659
R2113 VTAIL.n137 VTAIL.t13 147.659
R2114 VTAIL.n241 VTAIL.t10 147.659
R2115 VTAIL.n654 VTAIL.t12 147.659
R2116 VTAIL.n550 VTAIL.t11 147.659
R2117 VTAIL.n448 VTAIL.t0 147.659
R2118 VTAIL.n344 VTAIL.t3 147.659
R2119 VTAIL.n759 VTAIL.n753 104.615
R2120 VTAIL.n760 VTAIL.n759 104.615
R2121 VTAIL.n760 VTAIL.n749 104.615
R2122 VTAIL.n767 VTAIL.n749 104.615
R2123 VTAIL.n768 VTAIL.n767 104.615
R2124 VTAIL.n768 VTAIL.n745 104.615
R2125 VTAIL.n775 VTAIL.n745 104.615
R2126 VTAIL.n776 VTAIL.n775 104.615
R2127 VTAIL.n776 VTAIL.n741 104.615
R2128 VTAIL.n783 VTAIL.n741 104.615
R2129 VTAIL.n784 VTAIL.n783 104.615
R2130 VTAIL.n784 VTAIL.n737 104.615
R2131 VTAIL.n791 VTAIL.n737 104.615
R2132 VTAIL.n792 VTAIL.n791 104.615
R2133 VTAIL.n792 VTAIL.n733 104.615
R2134 VTAIL.n800 VTAIL.n733 104.615
R2135 VTAIL.n801 VTAIL.n800 104.615
R2136 VTAIL.n802 VTAIL.n801 104.615
R2137 VTAIL.n802 VTAIL.n729 104.615
R2138 VTAIL.n809 VTAIL.n729 104.615
R2139 VTAIL.n810 VTAIL.n809 104.615
R2140 VTAIL.n810 VTAIL.n725 104.615
R2141 VTAIL.n817 VTAIL.n725 104.615
R2142 VTAIL.n818 VTAIL.n817 104.615
R2143 VTAIL.n39 VTAIL.n33 104.615
R2144 VTAIL.n40 VTAIL.n39 104.615
R2145 VTAIL.n40 VTAIL.n29 104.615
R2146 VTAIL.n47 VTAIL.n29 104.615
R2147 VTAIL.n48 VTAIL.n47 104.615
R2148 VTAIL.n48 VTAIL.n25 104.615
R2149 VTAIL.n55 VTAIL.n25 104.615
R2150 VTAIL.n56 VTAIL.n55 104.615
R2151 VTAIL.n56 VTAIL.n21 104.615
R2152 VTAIL.n63 VTAIL.n21 104.615
R2153 VTAIL.n64 VTAIL.n63 104.615
R2154 VTAIL.n64 VTAIL.n17 104.615
R2155 VTAIL.n71 VTAIL.n17 104.615
R2156 VTAIL.n72 VTAIL.n71 104.615
R2157 VTAIL.n72 VTAIL.n13 104.615
R2158 VTAIL.n80 VTAIL.n13 104.615
R2159 VTAIL.n81 VTAIL.n80 104.615
R2160 VTAIL.n82 VTAIL.n81 104.615
R2161 VTAIL.n82 VTAIL.n9 104.615
R2162 VTAIL.n89 VTAIL.n9 104.615
R2163 VTAIL.n90 VTAIL.n89 104.615
R2164 VTAIL.n90 VTAIL.n5 104.615
R2165 VTAIL.n97 VTAIL.n5 104.615
R2166 VTAIL.n98 VTAIL.n97 104.615
R2167 VTAIL.n141 VTAIL.n135 104.615
R2168 VTAIL.n142 VTAIL.n141 104.615
R2169 VTAIL.n142 VTAIL.n131 104.615
R2170 VTAIL.n149 VTAIL.n131 104.615
R2171 VTAIL.n150 VTAIL.n149 104.615
R2172 VTAIL.n150 VTAIL.n127 104.615
R2173 VTAIL.n157 VTAIL.n127 104.615
R2174 VTAIL.n158 VTAIL.n157 104.615
R2175 VTAIL.n158 VTAIL.n123 104.615
R2176 VTAIL.n165 VTAIL.n123 104.615
R2177 VTAIL.n166 VTAIL.n165 104.615
R2178 VTAIL.n166 VTAIL.n119 104.615
R2179 VTAIL.n173 VTAIL.n119 104.615
R2180 VTAIL.n174 VTAIL.n173 104.615
R2181 VTAIL.n174 VTAIL.n115 104.615
R2182 VTAIL.n182 VTAIL.n115 104.615
R2183 VTAIL.n183 VTAIL.n182 104.615
R2184 VTAIL.n184 VTAIL.n183 104.615
R2185 VTAIL.n184 VTAIL.n111 104.615
R2186 VTAIL.n191 VTAIL.n111 104.615
R2187 VTAIL.n192 VTAIL.n191 104.615
R2188 VTAIL.n192 VTAIL.n107 104.615
R2189 VTAIL.n199 VTAIL.n107 104.615
R2190 VTAIL.n200 VTAIL.n199 104.615
R2191 VTAIL.n245 VTAIL.n239 104.615
R2192 VTAIL.n246 VTAIL.n245 104.615
R2193 VTAIL.n246 VTAIL.n235 104.615
R2194 VTAIL.n253 VTAIL.n235 104.615
R2195 VTAIL.n254 VTAIL.n253 104.615
R2196 VTAIL.n254 VTAIL.n231 104.615
R2197 VTAIL.n261 VTAIL.n231 104.615
R2198 VTAIL.n262 VTAIL.n261 104.615
R2199 VTAIL.n262 VTAIL.n227 104.615
R2200 VTAIL.n269 VTAIL.n227 104.615
R2201 VTAIL.n270 VTAIL.n269 104.615
R2202 VTAIL.n270 VTAIL.n223 104.615
R2203 VTAIL.n277 VTAIL.n223 104.615
R2204 VTAIL.n278 VTAIL.n277 104.615
R2205 VTAIL.n278 VTAIL.n219 104.615
R2206 VTAIL.n286 VTAIL.n219 104.615
R2207 VTAIL.n287 VTAIL.n286 104.615
R2208 VTAIL.n288 VTAIL.n287 104.615
R2209 VTAIL.n288 VTAIL.n215 104.615
R2210 VTAIL.n295 VTAIL.n215 104.615
R2211 VTAIL.n296 VTAIL.n295 104.615
R2212 VTAIL.n296 VTAIL.n211 104.615
R2213 VTAIL.n303 VTAIL.n211 104.615
R2214 VTAIL.n304 VTAIL.n303 104.615
R2215 VTAIL.n716 VTAIL.n715 104.615
R2216 VTAIL.n715 VTAIL.n623 104.615
R2217 VTAIL.n708 VTAIL.n623 104.615
R2218 VTAIL.n708 VTAIL.n707 104.615
R2219 VTAIL.n707 VTAIL.n627 104.615
R2220 VTAIL.n700 VTAIL.n627 104.615
R2221 VTAIL.n700 VTAIL.n699 104.615
R2222 VTAIL.n699 VTAIL.n698 104.615
R2223 VTAIL.n698 VTAIL.n631 104.615
R2224 VTAIL.n691 VTAIL.n631 104.615
R2225 VTAIL.n691 VTAIL.n690 104.615
R2226 VTAIL.n690 VTAIL.n636 104.615
R2227 VTAIL.n683 VTAIL.n636 104.615
R2228 VTAIL.n683 VTAIL.n682 104.615
R2229 VTAIL.n682 VTAIL.n640 104.615
R2230 VTAIL.n675 VTAIL.n640 104.615
R2231 VTAIL.n675 VTAIL.n674 104.615
R2232 VTAIL.n674 VTAIL.n644 104.615
R2233 VTAIL.n667 VTAIL.n644 104.615
R2234 VTAIL.n667 VTAIL.n666 104.615
R2235 VTAIL.n666 VTAIL.n648 104.615
R2236 VTAIL.n659 VTAIL.n648 104.615
R2237 VTAIL.n659 VTAIL.n658 104.615
R2238 VTAIL.n658 VTAIL.n652 104.615
R2239 VTAIL.n612 VTAIL.n611 104.615
R2240 VTAIL.n611 VTAIL.n519 104.615
R2241 VTAIL.n604 VTAIL.n519 104.615
R2242 VTAIL.n604 VTAIL.n603 104.615
R2243 VTAIL.n603 VTAIL.n523 104.615
R2244 VTAIL.n596 VTAIL.n523 104.615
R2245 VTAIL.n596 VTAIL.n595 104.615
R2246 VTAIL.n595 VTAIL.n594 104.615
R2247 VTAIL.n594 VTAIL.n527 104.615
R2248 VTAIL.n587 VTAIL.n527 104.615
R2249 VTAIL.n587 VTAIL.n586 104.615
R2250 VTAIL.n586 VTAIL.n532 104.615
R2251 VTAIL.n579 VTAIL.n532 104.615
R2252 VTAIL.n579 VTAIL.n578 104.615
R2253 VTAIL.n578 VTAIL.n536 104.615
R2254 VTAIL.n571 VTAIL.n536 104.615
R2255 VTAIL.n571 VTAIL.n570 104.615
R2256 VTAIL.n570 VTAIL.n540 104.615
R2257 VTAIL.n563 VTAIL.n540 104.615
R2258 VTAIL.n563 VTAIL.n562 104.615
R2259 VTAIL.n562 VTAIL.n544 104.615
R2260 VTAIL.n555 VTAIL.n544 104.615
R2261 VTAIL.n555 VTAIL.n554 104.615
R2262 VTAIL.n554 VTAIL.n548 104.615
R2263 VTAIL.n510 VTAIL.n509 104.615
R2264 VTAIL.n509 VTAIL.n417 104.615
R2265 VTAIL.n502 VTAIL.n417 104.615
R2266 VTAIL.n502 VTAIL.n501 104.615
R2267 VTAIL.n501 VTAIL.n421 104.615
R2268 VTAIL.n494 VTAIL.n421 104.615
R2269 VTAIL.n494 VTAIL.n493 104.615
R2270 VTAIL.n493 VTAIL.n492 104.615
R2271 VTAIL.n492 VTAIL.n425 104.615
R2272 VTAIL.n485 VTAIL.n425 104.615
R2273 VTAIL.n485 VTAIL.n484 104.615
R2274 VTAIL.n484 VTAIL.n430 104.615
R2275 VTAIL.n477 VTAIL.n430 104.615
R2276 VTAIL.n477 VTAIL.n476 104.615
R2277 VTAIL.n476 VTAIL.n434 104.615
R2278 VTAIL.n469 VTAIL.n434 104.615
R2279 VTAIL.n469 VTAIL.n468 104.615
R2280 VTAIL.n468 VTAIL.n438 104.615
R2281 VTAIL.n461 VTAIL.n438 104.615
R2282 VTAIL.n461 VTAIL.n460 104.615
R2283 VTAIL.n460 VTAIL.n442 104.615
R2284 VTAIL.n453 VTAIL.n442 104.615
R2285 VTAIL.n453 VTAIL.n452 104.615
R2286 VTAIL.n452 VTAIL.n446 104.615
R2287 VTAIL.n406 VTAIL.n405 104.615
R2288 VTAIL.n405 VTAIL.n313 104.615
R2289 VTAIL.n398 VTAIL.n313 104.615
R2290 VTAIL.n398 VTAIL.n397 104.615
R2291 VTAIL.n397 VTAIL.n317 104.615
R2292 VTAIL.n390 VTAIL.n317 104.615
R2293 VTAIL.n390 VTAIL.n389 104.615
R2294 VTAIL.n389 VTAIL.n388 104.615
R2295 VTAIL.n388 VTAIL.n321 104.615
R2296 VTAIL.n381 VTAIL.n321 104.615
R2297 VTAIL.n381 VTAIL.n380 104.615
R2298 VTAIL.n380 VTAIL.n326 104.615
R2299 VTAIL.n373 VTAIL.n326 104.615
R2300 VTAIL.n373 VTAIL.n372 104.615
R2301 VTAIL.n372 VTAIL.n330 104.615
R2302 VTAIL.n365 VTAIL.n330 104.615
R2303 VTAIL.n365 VTAIL.n364 104.615
R2304 VTAIL.n364 VTAIL.n334 104.615
R2305 VTAIL.n357 VTAIL.n334 104.615
R2306 VTAIL.n357 VTAIL.n356 104.615
R2307 VTAIL.n356 VTAIL.n338 104.615
R2308 VTAIL.n349 VTAIL.n338 104.615
R2309 VTAIL.n349 VTAIL.n348 104.615
R2310 VTAIL.n348 VTAIL.n342 104.615
R2311 VTAIL.t6 VTAIL.n753 52.3082
R2312 VTAIL.t5 VTAIL.n33 52.3082
R2313 VTAIL.t13 VTAIL.n135 52.3082
R2314 VTAIL.t10 VTAIL.n239 52.3082
R2315 VTAIL.t12 VTAIL.n652 52.3082
R2316 VTAIL.t11 VTAIL.n548 52.3082
R2317 VTAIL.t0 VTAIL.n446 52.3082
R2318 VTAIL.t3 VTAIL.n342 52.3082
R2319 VTAIL.n619 VTAIL.n618 44.5513
R2320 VTAIL.n413 VTAIL.n412 44.5513
R2321 VTAIL.n1 VTAIL.n0 44.5511
R2322 VTAIL.n207 VTAIL.n206 44.5511
R2323 VTAIL.n823 VTAIL.n822 32.7672
R2324 VTAIL.n103 VTAIL.n102 32.7672
R2325 VTAIL.n205 VTAIL.n204 32.7672
R2326 VTAIL.n309 VTAIL.n308 32.7672
R2327 VTAIL.n721 VTAIL.n720 32.7672
R2328 VTAIL.n617 VTAIL.n616 32.7672
R2329 VTAIL.n515 VTAIL.n514 32.7672
R2330 VTAIL.n411 VTAIL.n410 32.7672
R2331 VTAIL.n823 VTAIL.n721 30.0307
R2332 VTAIL.n411 VTAIL.n309 30.0307
R2333 VTAIL.n755 VTAIL.n754 15.6677
R2334 VTAIL.n35 VTAIL.n34 15.6677
R2335 VTAIL.n137 VTAIL.n136 15.6677
R2336 VTAIL.n241 VTAIL.n240 15.6677
R2337 VTAIL.n654 VTAIL.n653 15.6677
R2338 VTAIL.n550 VTAIL.n549 15.6677
R2339 VTAIL.n448 VTAIL.n447 15.6677
R2340 VTAIL.n344 VTAIL.n343 15.6677
R2341 VTAIL.n803 VTAIL.n732 13.1884
R2342 VTAIL.n83 VTAIL.n12 13.1884
R2343 VTAIL.n185 VTAIL.n114 13.1884
R2344 VTAIL.n289 VTAIL.n218 13.1884
R2345 VTAIL.n701 VTAIL.n630 13.1884
R2346 VTAIL.n597 VTAIL.n526 13.1884
R2347 VTAIL.n495 VTAIL.n424 13.1884
R2348 VTAIL.n391 VTAIL.n320 13.1884
R2349 VTAIL.n758 VTAIL.n757 12.8005
R2350 VTAIL.n799 VTAIL.n798 12.8005
R2351 VTAIL.n804 VTAIL.n730 12.8005
R2352 VTAIL.n38 VTAIL.n37 12.8005
R2353 VTAIL.n79 VTAIL.n78 12.8005
R2354 VTAIL.n84 VTAIL.n10 12.8005
R2355 VTAIL.n140 VTAIL.n139 12.8005
R2356 VTAIL.n181 VTAIL.n180 12.8005
R2357 VTAIL.n186 VTAIL.n112 12.8005
R2358 VTAIL.n244 VTAIL.n243 12.8005
R2359 VTAIL.n285 VTAIL.n284 12.8005
R2360 VTAIL.n290 VTAIL.n216 12.8005
R2361 VTAIL.n702 VTAIL.n628 12.8005
R2362 VTAIL.n697 VTAIL.n632 12.8005
R2363 VTAIL.n657 VTAIL.n656 12.8005
R2364 VTAIL.n598 VTAIL.n524 12.8005
R2365 VTAIL.n593 VTAIL.n528 12.8005
R2366 VTAIL.n553 VTAIL.n552 12.8005
R2367 VTAIL.n496 VTAIL.n422 12.8005
R2368 VTAIL.n491 VTAIL.n426 12.8005
R2369 VTAIL.n451 VTAIL.n450 12.8005
R2370 VTAIL.n392 VTAIL.n318 12.8005
R2371 VTAIL.n387 VTAIL.n322 12.8005
R2372 VTAIL.n347 VTAIL.n346 12.8005
R2373 VTAIL.n761 VTAIL.n752 12.0247
R2374 VTAIL.n797 VTAIL.n734 12.0247
R2375 VTAIL.n808 VTAIL.n807 12.0247
R2376 VTAIL.n41 VTAIL.n32 12.0247
R2377 VTAIL.n77 VTAIL.n14 12.0247
R2378 VTAIL.n88 VTAIL.n87 12.0247
R2379 VTAIL.n143 VTAIL.n134 12.0247
R2380 VTAIL.n179 VTAIL.n116 12.0247
R2381 VTAIL.n190 VTAIL.n189 12.0247
R2382 VTAIL.n247 VTAIL.n238 12.0247
R2383 VTAIL.n283 VTAIL.n220 12.0247
R2384 VTAIL.n294 VTAIL.n293 12.0247
R2385 VTAIL.n706 VTAIL.n705 12.0247
R2386 VTAIL.n696 VTAIL.n633 12.0247
R2387 VTAIL.n660 VTAIL.n651 12.0247
R2388 VTAIL.n602 VTAIL.n601 12.0247
R2389 VTAIL.n592 VTAIL.n529 12.0247
R2390 VTAIL.n556 VTAIL.n547 12.0247
R2391 VTAIL.n500 VTAIL.n499 12.0247
R2392 VTAIL.n490 VTAIL.n427 12.0247
R2393 VTAIL.n454 VTAIL.n445 12.0247
R2394 VTAIL.n396 VTAIL.n395 12.0247
R2395 VTAIL.n386 VTAIL.n323 12.0247
R2396 VTAIL.n350 VTAIL.n341 12.0247
R2397 VTAIL.n762 VTAIL.n750 11.249
R2398 VTAIL.n794 VTAIL.n793 11.249
R2399 VTAIL.n811 VTAIL.n728 11.249
R2400 VTAIL.n42 VTAIL.n30 11.249
R2401 VTAIL.n74 VTAIL.n73 11.249
R2402 VTAIL.n91 VTAIL.n8 11.249
R2403 VTAIL.n144 VTAIL.n132 11.249
R2404 VTAIL.n176 VTAIL.n175 11.249
R2405 VTAIL.n193 VTAIL.n110 11.249
R2406 VTAIL.n248 VTAIL.n236 11.249
R2407 VTAIL.n280 VTAIL.n279 11.249
R2408 VTAIL.n297 VTAIL.n214 11.249
R2409 VTAIL.n709 VTAIL.n626 11.249
R2410 VTAIL.n693 VTAIL.n692 11.249
R2411 VTAIL.n661 VTAIL.n649 11.249
R2412 VTAIL.n605 VTAIL.n522 11.249
R2413 VTAIL.n589 VTAIL.n588 11.249
R2414 VTAIL.n557 VTAIL.n545 11.249
R2415 VTAIL.n503 VTAIL.n420 11.249
R2416 VTAIL.n487 VTAIL.n486 11.249
R2417 VTAIL.n455 VTAIL.n443 11.249
R2418 VTAIL.n399 VTAIL.n316 11.249
R2419 VTAIL.n383 VTAIL.n382 11.249
R2420 VTAIL.n351 VTAIL.n339 11.249
R2421 VTAIL.n766 VTAIL.n765 10.4732
R2422 VTAIL.n790 VTAIL.n736 10.4732
R2423 VTAIL.n812 VTAIL.n726 10.4732
R2424 VTAIL.n46 VTAIL.n45 10.4732
R2425 VTAIL.n70 VTAIL.n16 10.4732
R2426 VTAIL.n92 VTAIL.n6 10.4732
R2427 VTAIL.n148 VTAIL.n147 10.4732
R2428 VTAIL.n172 VTAIL.n118 10.4732
R2429 VTAIL.n194 VTAIL.n108 10.4732
R2430 VTAIL.n252 VTAIL.n251 10.4732
R2431 VTAIL.n276 VTAIL.n222 10.4732
R2432 VTAIL.n298 VTAIL.n212 10.4732
R2433 VTAIL.n710 VTAIL.n624 10.4732
R2434 VTAIL.n689 VTAIL.n635 10.4732
R2435 VTAIL.n665 VTAIL.n664 10.4732
R2436 VTAIL.n606 VTAIL.n520 10.4732
R2437 VTAIL.n585 VTAIL.n531 10.4732
R2438 VTAIL.n561 VTAIL.n560 10.4732
R2439 VTAIL.n504 VTAIL.n418 10.4732
R2440 VTAIL.n483 VTAIL.n429 10.4732
R2441 VTAIL.n459 VTAIL.n458 10.4732
R2442 VTAIL.n400 VTAIL.n314 10.4732
R2443 VTAIL.n379 VTAIL.n325 10.4732
R2444 VTAIL.n355 VTAIL.n354 10.4732
R2445 VTAIL.n769 VTAIL.n748 9.69747
R2446 VTAIL.n789 VTAIL.n738 9.69747
R2447 VTAIL.n816 VTAIL.n815 9.69747
R2448 VTAIL.n49 VTAIL.n28 9.69747
R2449 VTAIL.n69 VTAIL.n18 9.69747
R2450 VTAIL.n96 VTAIL.n95 9.69747
R2451 VTAIL.n151 VTAIL.n130 9.69747
R2452 VTAIL.n171 VTAIL.n120 9.69747
R2453 VTAIL.n198 VTAIL.n197 9.69747
R2454 VTAIL.n255 VTAIL.n234 9.69747
R2455 VTAIL.n275 VTAIL.n224 9.69747
R2456 VTAIL.n302 VTAIL.n301 9.69747
R2457 VTAIL.n714 VTAIL.n713 9.69747
R2458 VTAIL.n688 VTAIL.n637 9.69747
R2459 VTAIL.n668 VTAIL.n647 9.69747
R2460 VTAIL.n610 VTAIL.n609 9.69747
R2461 VTAIL.n584 VTAIL.n533 9.69747
R2462 VTAIL.n564 VTAIL.n543 9.69747
R2463 VTAIL.n508 VTAIL.n507 9.69747
R2464 VTAIL.n482 VTAIL.n431 9.69747
R2465 VTAIL.n462 VTAIL.n441 9.69747
R2466 VTAIL.n404 VTAIL.n403 9.69747
R2467 VTAIL.n378 VTAIL.n327 9.69747
R2468 VTAIL.n358 VTAIL.n337 9.69747
R2469 VTAIL.n822 VTAIL.n821 9.45567
R2470 VTAIL.n102 VTAIL.n101 9.45567
R2471 VTAIL.n204 VTAIL.n203 9.45567
R2472 VTAIL.n308 VTAIL.n307 9.45567
R2473 VTAIL.n720 VTAIL.n719 9.45567
R2474 VTAIL.n616 VTAIL.n615 9.45567
R2475 VTAIL.n514 VTAIL.n513 9.45567
R2476 VTAIL.n410 VTAIL.n409 9.45567
R2477 VTAIL.n821 VTAIL.n820 9.3005
R2478 VTAIL.n724 VTAIL.n723 9.3005
R2479 VTAIL.n815 VTAIL.n814 9.3005
R2480 VTAIL.n813 VTAIL.n812 9.3005
R2481 VTAIL.n728 VTAIL.n727 9.3005
R2482 VTAIL.n807 VTAIL.n806 9.3005
R2483 VTAIL.n805 VTAIL.n804 9.3005
R2484 VTAIL.n744 VTAIL.n743 9.3005
R2485 VTAIL.n773 VTAIL.n772 9.3005
R2486 VTAIL.n771 VTAIL.n770 9.3005
R2487 VTAIL.n748 VTAIL.n747 9.3005
R2488 VTAIL.n765 VTAIL.n764 9.3005
R2489 VTAIL.n763 VTAIL.n762 9.3005
R2490 VTAIL.n752 VTAIL.n751 9.3005
R2491 VTAIL.n757 VTAIL.n756 9.3005
R2492 VTAIL.n779 VTAIL.n778 9.3005
R2493 VTAIL.n781 VTAIL.n780 9.3005
R2494 VTAIL.n740 VTAIL.n739 9.3005
R2495 VTAIL.n787 VTAIL.n786 9.3005
R2496 VTAIL.n789 VTAIL.n788 9.3005
R2497 VTAIL.n736 VTAIL.n735 9.3005
R2498 VTAIL.n795 VTAIL.n794 9.3005
R2499 VTAIL.n797 VTAIL.n796 9.3005
R2500 VTAIL.n798 VTAIL.n731 9.3005
R2501 VTAIL.n101 VTAIL.n100 9.3005
R2502 VTAIL.n4 VTAIL.n3 9.3005
R2503 VTAIL.n95 VTAIL.n94 9.3005
R2504 VTAIL.n93 VTAIL.n92 9.3005
R2505 VTAIL.n8 VTAIL.n7 9.3005
R2506 VTAIL.n87 VTAIL.n86 9.3005
R2507 VTAIL.n85 VTAIL.n84 9.3005
R2508 VTAIL.n24 VTAIL.n23 9.3005
R2509 VTAIL.n53 VTAIL.n52 9.3005
R2510 VTAIL.n51 VTAIL.n50 9.3005
R2511 VTAIL.n28 VTAIL.n27 9.3005
R2512 VTAIL.n45 VTAIL.n44 9.3005
R2513 VTAIL.n43 VTAIL.n42 9.3005
R2514 VTAIL.n32 VTAIL.n31 9.3005
R2515 VTAIL.n37 VTAIL.n36 9.3005
R2516 VTAIL.n59 VTAIL.n58 9.3005
R2517 VTAIL.n61 VTAIL.n60 9.3005
R2518 VTAIL.n20 VTAIL.n19 9.3005
R2519 VTAIL.n67 VTAIL.n66 9.3005
R2520 VTAIL.n69 VTAIL.n68 9.3005
R2521 VTAIL.n16 VTAIL.n15 9.3005
R2522 VTAIL.n75 VTAIL.n74 9.3005
R2523 VTAIL.n77 VTAIL.n76 9.3005
R2524 VTAIL.n78 VTAIL.n11 9.3005
R2525 VTAIL.n203 VTAIL.n202 9.3005
R2526 VTAIL.n106 VTAIL.n105 9.3005
R2527 VTAIL.n197 VTAIL.n196 9.3005
R2528 VTAIL.n195 VTAIL.n194 9.3005
R2529 VTAIL.n110 VTAIL.n109 9.3005
R2530 VTAIL.n189 VTAIL.n188 9.3005
R2531 VTAIL.n187 VTAIL.n186 9.3005
R2532 VTAIL.n126 VTAIL.n125 9.3005
R2533 VTAIL.n155 VTAIL.n154 9.3005
R2534 VTAIL.n153 VTAIL.n152 9.3005
R2535 VTAIL.n130 VTAIL.n129 9.3005
R2536 VTAIL.n147 VTAIL.n146 9.3005
R2537 VTAIL.n145 VTAIL.n144 9.3005
R2538 VTAIL.n134 VTAIL.n133 9.3005
R2539 VTAIL.n139 VTAIL.n138 9.3005
R2540 VTAIL.n161 VTAIL.n160 9.3005
R2541 VTAIL.n163 VTAIL.n162 9.3005
R2542 VTAIL.n122 VTAIL.n121 9.3005
R2543 VTAIL.n169 VTAIL.n168 9.3005
R2544 VTAIL.n171 VTAIL.n170 9.3005
R2545 VTAIL.n118 VTAIL.n117 9.3005
R2546 VTAIL.n177 VTAIL.n176 9.3005
R2547 VTAIL.n179 VTAIL.n178 9.3005
R2548 VTAIL.n180 VTAIL.n113 9.3005
R2549 VTAIL.n307 VTAIL.n306 9.3005
R2550 VTAIL.n210 VTAIL.n209 9.3005
R2551 VTAIL.n301 VTAIL.n300 9.3005
R2552 VTAIL.n299 VTAIL.n298 9.3005
R2553 VTAIL.n214 VTAIL.n213 9.3005
R2554 VTAIL.n293 VTAIL.n292 9.3005
R2555 VTAIL.n291 VTAIL.n290 9.3005
R2556 VTAIL.n230 VTAIL.n229 9.3005
R2557 VTAIL.n259 VTAIL.n258 9.3005
R2558 VTAIL.n257 VTAIL.n256 9.3005
R2559 VTAIL.n234 VTAIL.n233 9.3005
R2560 VTAIL.n251 VTAIL.n250 9.3005
R2561 VTAIL.n249 VTAIL.n248 9.3005
R2562 VTAIL.n238 VTAIL.n237 9.3005
R2563 VTAIL.n243 VTAIL.n242 9.3005
R2564 VTAIL.n265 VTAIL.n264 9.3005
R2565 VTAIL.n267 VTAIL.n266 9.3005
R2566 VTAIL.n226 VTAIL.n225 9.3005
R2567 VTAIL.n273 VTAIL.n272 9.3005
R2568 VTAIL.n275 VTAIL.n274 9.3005
R2569 VTAIL.n222 VTAIL.n221 9.3005
R2570 VTAIL.n281 VTAIL.n280 9.3005
R2571 VTAIL.n283 VTAIL.n282 9.3005
R2572 VTAIL.n284 VTAIL.n217 9.3005
R2573 VTAIL.n680 VTAIL.n679 9.3005
R2574 VTAIL.n639 VTAIL.n638 9.3005
R2575 VTAIL.n686 VTAIL.n685 9.3005
R2576 VTAIL.n688 VTAIL.n687 9.3005
R2577 VTAIL.n635 VTAIL.n634 9.3005
R2578 VTAIL.n694 VTAIL.n693 9.3005
R2579 VTAIL.n696 VTAIL.n695 9.3005
R2580 VTAIL.n632 VTAIL.n629 9.3005
R2581 VTAIL.n719 VTAIL.n718 9.3005
R2582 VTAIL.n622 VTAIL.n621 9.3005
R2583 VTAIL.n713 VTAIL.n712 9.3005
R2584 VTAIL.n711 VTAIL.n710 9.3005
R2585 VTAIL.n626 VTAIL.n625 9.3005
R2586 VTAIL.n705 VTAIL.n704 9.3005
R2587 VTAIL.n703 VTAIL.n702 9.3005
R2588 VTAIL.n678 VTAIL.n677 9.3005
R2589 VTAIL.n643 VTAIL.n642 9.3005
R2590 VTAIL.n672 VTAIL.n671 9.3005
R2591 VTAIL.n670 VTAIL.n669 9.3005
R2592 VTAIL.n647 VTAIL.n646 9.3005
R2593 VTAIL.n664 VTAIL.n663 9.3005
R2594 VTAIL.n662 VTAIL.n661 9.3005
R2595 VTAIL.n651 VTAIL.n650 9.3005
R2596 VTAIL.n656 VTAIL.n655 9.3005
R2597 VTAIL.n576 VTAIL.n575 9.3005
R2598 VTAIL.n535 VTAIL.n534 9.3005
R2599 VTAIL.n582 VTAIL.n581 9.3005
R2600 VTAIL.n584 VTAIL.n583 9.3005
R2601 VTAIL.n531 VTAIL.n530 9.3005
R2602 VTAIL.n590 VTAIL.n589 9.3005
R2603 VTAIL.n592 VTAIL.n591 9.3005
R2604 VTAIL.n528 VTAIL.n525 9.3005
R2605 VTAIL.n615 VTAIL.n614 9.3005
R2606 VTAIL.n518 VTAIL.n517 9.3005
R2607 VTAIL.n609 VTAIL.n608 9.3005
R2608 VTAIL.n607 VTAIL.n606 9.3005
R2609 VTAIL.n522 VTAIL.n521 9.3005
R2610 VTAIL.n601 VTAIL.n600 9.3005
R2611 VTAIL.n599 VTAIL.n598 9.3005
R2612 VTAIL.n574 VTAIL.n573 9.3005
R2613 VTAIL.n539 VTAIL.n538 9.3005
R2614 VTAIL.n568 VTAIL.n567 9.3005
R2615 VTAIL.n566 VTAIL.n565 9.3005
R2616 VTAIL.n543 VTAIL.n542 9.3005
R2617 VTAIL.n560 VTAIL.n559 9.3005
R2618 VTAIL.n558 VTAIL.n557 9.3005
R2619 VTAIL.n547 VTAIL.n546 9.3005
R2620 VTAIL.n552 VTAIL.n551 9.3005
R2621 VTAIL.n474 VTAIL.n473 9.3005
R2622 VTAIL.n433 VTAIL.n432 9.3005
R2623 VTAIL.n480 VTAIL.n479 9.3005
R2624 VTAIL.n482 VTAIL.n481 9.3005
R2625 VTAIL.n429 VTAIL.n428 9.3005
R2626 VTAIL.n488 VTAIL.n487 9.3005
R2627 VTAIL.n490 VTAIL.n489 9.3005
R2628 VTAIL.n426 VTAIL.n423 9.3005
R2629 VTAIL.n513 VTAIL.n512 9.3005
R2630 VTAIL.n416 VTAIL.n415 9.3005
R2631 VTAIL.n507 VTAIL.n506 9.3005
R2632 VTAIL.n505 VTAIL.n504 9.3005
R2633 VTAIL.n420 VTAIL.n419 9.3005
R2634 VTAIL.n499 VTAIL.n498 9.3005
R2635 VTAIL.n497 VTAIL.n496 9.3005
R2636 VTAIL.n472 VTAIL.n471 9.3005
R2637 VTAIL.n437 VTAIL.n436 9.3005
R2638 VTAIL.n466 VTAIL.n465 9.3005
R2639 VTAIL.n464 VTAIL.n463 9.3005
R2640 VTAIL.n441 VTAIL.n440 9.3005
R2641 VTAIL.n458 VTAIL.n457 9.3005
R2642 VTAIL.n456 VTAIL.n455 9.3005
R2643 VTAIL.n445 VTAIL.n444 9.3005
R2644 VTAIL.n450 VTAIL.n449 9.3005
R2645 VTAIL.n370 VTAIL.n369 9.3005
R2646 VTAIL.n329 VTAIL.n328 9.3005
R2647 VTAIL.n376 VTAIL.n375 9.3005
R2648 VTAIL.n378 VTAIL.n377 9.3005
R2649 VTAIL.n325 VTAIL.n324 9.3005
R2650 VTAIL.n384 VTAIL.n383 9.3005
R2651 VTAIL.n386 VTAIL.n385 9.3005
R2652 VTAIL.n322 VTAIL.n319 9.3005
R2653 VTAIL.n409 VTAIL.n408 9.3005
R2654 VTAIL.n312 VTAIL.n311 9.3005
R2655 VTAIL.n403 VTAIL.n402 9.3005
R2656 VTAIL.n401 VTAIL.n400 9.3005
R2657 VTAIL.n316 VTAIL.n315 9.3005
R2658 VTAIL.n395 VTAIL.n394 9.3005
R2659 VTAIL.n393 VTAIL.n392 9.3005
R2660 VTAIL.n368 VTAIL.n367 9.3005
R2661 VTAIL.n333 VTAIL.n332 9.3005
R2662 VTAIL.n362 VTAIL.n361 9.3005
R2663 VTAIL.n360 VTAIL.n359 9.3005
R2664 VTAIL.n337 VTAIL.n336 9.3005
R2665 VTAIL.n354 VTAIL.n353 9.3005
R2666 VTAIL.n352 VTAIL.n351 9.3005
R2667 VTAIL.n341 VTAIL.n340 9.3005
R2668 VTAIL.n346 VTAIL.n345 9.3005
R2669 VTAIL.n770 VTAIL.n746 8.92171
R2670 VTAIL.n786 VTAIL.n785 8.92171
R2671 VTAIL.n819 VTAIL.n724 8.92171
R2672 VTAIL.n50 VTAIL.n26 8.92171
R2673 VTAIL.n66 VTAIL.n65 8.92171
R2674 VTAIL.n99 VTAIL.n4 8.92171
R2675 VTAIL.n152 VTAIL.n128 8.92171
R2676 VTAIL.n168 VTAIL.n167 8.92171
R2677 VTAIL.n201 VTAIL.n106 8.92171
R2678 VTAIL.n256 VTAIL.n232 8.92171
R2679 VTAIL.n272 VTAIL.n271 8.92171
R2680 VTAIL.n305 VTAIL.n210 8.92171
R2681 VTAIL.n717 VTAIL.n622 8.92171
R2682 VTAIL.n685 VTAIL.n684 8.92171
R2683 VTAIL.n669 VTAIL.n645 8.92171
R2684 VTAIL.n613 VTAIL.n518 8.92171
R2685 VTAIL.n581 VTAIL.n580 8.92171
R2686 VTAIL.n565 VTAIL.n541 8.92171
R2687 VTAIL.n511 VTAIL.n416 8.92171
R2688 VTAIL.n479 VTAIL.n478 8.92171
R2689 VTAIL.n463 VTAIL.n439 8.92171
R2690 VTAIL.n407 VTAIL.n312 8.92171
R2691 VTAIL.n375 VTAIL.n374 8.92171
R2692 VTAIL.n359 VTAIL.n335 8.92171
R2693 VTAIL.n774 VTAIL.n773 8.14595
R2694 VTAIL.n782 VTAIL.n740 8.14595
R2695 VTAIL.n820 VTAIL.n722 8.14595
R2696 VTAIL.n54 VTAIL.n53 8.14595
R2697 VTAIL.n62 VTAIL.n20 8.14595
R2698 VTAIL.n100 VTAIL.n2 8.14595
R2699 VTAIL.n156 VTAIL.n155 8.14595
R2700 VTAIL.n164 VTAIL.n122 8.14595
R2701 VTAIL.n202 VTAIL.n104 8.14595
R2702 VTAIL.n260 VTAIL.n259 8.14595
R2703 VTAIL.n268 VTAIL.n226 8.14595
R2704 VTAIL.n306 VTAIL.n208 8.14595
R2705 VTAIL.n718 VTAIL.n620 8.14595
R2706 VTAIL.n681 VTAIL.n639 8.14595
R2707 VTAIL.n673 VTAIL.n672 8.14595
R2708 VTAIL.n614 VTAIL.n516 8.14595
R2709 VTAIL.n577 VTAIL.n535 8.14595
R2710 VTAIL.n569 VTAIL.n568 8.14595
R2711 VTAIL.n512 VTAIL.n414 8.14595
R2712 VTAIL.n475 VTAIL.n433 8.14595
R2713 VTAIL.n467 VTAIL.n466 8.14595
R2714 VTAIL.n408 VTAIL.n310 8.14595
R2715 VTAIL.n371 VTAIL.n329 8.14595
R2716 VTAIL.n363 VTAIL.n362 8.14595
R2717 VTAIL.n777 VTAIL.n744 7.3702
R2718 VTAIL.n781 VTAIL.n742 7.3702
R2719 VTAIL.n57 VTAIL.n24 7.3702
R2720 VTAIL.n61 VTAIL.n22 7.3702
R2721 VTAIL.n159 VTAIL.n126 7.3702
R2722 VTAIL.n163 VTAIL.n124 7.3702
R2723 VTAIL.n263 VTAIL.n230 7.3702
R2724 VTAIL.n267 VTAIL.n228 7.3702
R2725 VTAIL.n680 VTAIL.n641 7.3702
R2726 VTAIL.n676 VTAIL.n643 7.3702
R2727 VTAIL.n576 VTAIL.n537 7.3702
R2728 VTAIL.n572 VTAIL.n539 7.3702
R2729 VTAIL.n474 VTAIL.n435 7.3702
R2730 VTAIL.n470 VTAIL.n437 7.3702
R2731 VTAIL.n370 VTAIL.n331 7.3702
R2732 VTAIL.n366 VTAIL.n333 7.3702
R2733 VTAIL.n778 VTAIL.n777 6.59444
R2734 VTAIL.n778 VTAIL.n742 6.59444
R2735 VTAIL.n58 VTAIL.n57 6.59444
R2736 VTAIL.n58 VTAIL.n22 6.59444
R2737 VTAIL.n160 VTAIL.n159 6.59444
R2738 VTAIL.n160 VTAIL.n124 6.59444
R2739 VTAIL.n264 VTAIL.n263 6.59444
R2740 VTAIL.n264 VTAIL.n228 6.59444
R2741 VTAIL.n677 VTAIL.n641 6.59444
R2742 VTAIL.n677 VTAIL.n676 6.59444
R2743 VTAIL.n573 VTAIL.n537 6.59444
R2744 VTAIL.n573 VTAIL.n572 6.59444
R2745 VTAIL.n471 VTAIL.n435 6.59444
R2746 VTAIL.n471 VTAIL.n470 6.59444
R2747 VTAIL.n367 VTAIL.n331 6.59444
R2748 VTAIL.n367 VTAIL.n366 6.59444
R2749 VTAIL.n774 VTAIL.n744 5.81868
R2750 VTAIL.n782 VTAIL.n781 5.81868
R2751 VTAIL.n822 VTAIL.n722 5.81868
R2752 VTAIL.n54 VTAIL.n24 5.81868
R2753 VTAIL.n62 VTAIL.n61 5.81868
R2754 VTAIL.n102 VTAIL.n2 5.81868
R2755 VTAIL.n156 VTAIL.n126 5.81868
R2756 VTAIL.n164 VTAIL.n163 5.81868
R2757 VTAIL.n204 VTAIL.n104 5.81868
R2758 VTAIL.n260 VTAIL.n230 5.81868
R2759 VTAIL.n268 VTAIL.n267 5.81868
R2760 VTAIL.n308 VTAIL.n208 5.81868
R2761 VTAIL.n720 VTAIL.n620 5.81868
R2762 VTAIL.n681 VTAIL.n680 5.81868
R2763 VTAIL.n673 VTAIL.n643 5.81868
R2764 VTAIL.n616 VTAIL.n516 5.81868
R2765 VTAIL.n577 VTAIL.n576 5.81868
R2766 VTAIL.n569 VTAIL.n539 5.81868
R2767 VTAIL.n514 VTAIL.n414 5.81868
R2768 VTAIL.n475 VTAIL.n474 5.81868
R2769 VTAIL.n467 VTAIL.n437 5.81868
R2770 VTAIL.n410 VTAIL.n310 5.81868
R2771 VTAIL.n371 VTAIL.n370 5.81868
R2772 VTAIL.n363 VTAIL.n333 5.81868
R2773 VTAIL.n773 VTAIL.n746 5.04292
R2774 VTAIL.n785 VTAIL.n740 5.04292
R2775 VTAIL.n820 VTAIL.n819 5.04292
R2776 VTAIL.n53 VTAIL.n26 5.04292
R2777 VTAIL.n65 VTAIL.n20 5.04292
R2778 VTAIL.n100 VTAIL.n99 5.04292
R2779 VTAIL.n155 VTAIL.n128 5.04292
R2780 VTAIL.n167 VTAIL.n122 5.04292
R2781 VTAIL.n202 VTAIL.n201 5.04292
R2782 VTAIL.n259 VTAIL.n232 5.04292
R2783 VTAIL.n271 VTAIL.n226 5.04292
R2784 VTAIL.n306 VTAIL.n305 5.04292
R2785 VTAIL.n718 VTAIL.n717 5.04292
R2786 VTAIL.n684 VTAIL.n639 5.04292
R2787 VTAIL.n672 VTAIL.n645 5.04292
R2788 VTAIL.n614 VTAIL.n613 5.04292
R2789 VTAIL.n580 VTAIL.n535 5.04292
R2790 VTAIL.n568 VTAIL.n541 5.04292
R2791 VTAIL.n512 VTAIL.n511 5.04292
R2792 VTAIL.n478 VTAIL.n433 5.04292
R2793 VTAIL.n466 VTAIL.n439 5.04292
R2794 VTAIL.n408 VTAIL.n407 5.04292
R2795 VTAIL.n374 VTAIL.n329 5.04292
R2796 VTAIL.n362 VTAIL.n335 5.04292
R2797 VTAIL.n756 VTAIL.n755 4.38563
R2798 VTAIL.n36 VTAIL.n35 4.38563
R2799 VTAIL.n138 VTAIL.n137 4.38563
R2800 VTAIL.n242 VTAIL.n241 4.38563
R2801 VTAIL.n655 VTAIL.n654 4.38563
R2802 VTAIL.n551 VTAIL.n550 4.38563
R2803 VTAIL.n449 VTAIL.n448 4.38563
R2804 VTAIL.n345 VTAIL.n344 4.38563
R2805 VTAIL.n770 VTAIL.n769 4.26717
R2806 VTAIL.n786 VTAIL.n738 4.26717
R2807 VTAIL.n816 VTAIL.n724 4.26717
R2808 VTAIL.n50 VTAIL.n49 4.26717
R2809 VTAIL.n66 VTAIL.n18 4.26717
R2810 VTAIL.n96 VTAIL.n4 4.26717
R2811 VTAIL.n152 VTAIL.n151 4.26717
R2812 VTAIL.n168 VTAIL.n120 4.26717
R2813 VTAIL.n198 VTAIL.n106 4.26717
R2814 VTAIL.n256 VTAIL.n255 4.26717
R2815 VTAIL.n272 VTAIL.n224 4.26717
R2816 VTAIL.n302 VTAIL.n210 4.26717
R2817 VTAIL.n714 VTAIL.n622 4.26717
R2818 VTAIL.n685 VTAIL.n637 4.26717
R2819 VTAIL.n669 VTAIL.n668 4.26717
R2820 VTAIL.n610 VTAIL.n518 4.26717
R2821 VTAIL.n581 VTAIL.n533 4.26717
R2822 VTAIL.n565 VTAIL.n564 4.26717
R2823 VTAIL.n508 VTAIL.n416 4.26717
R2824 VTAIL.n479 VTAIL.n431 4.26717
R2825 VTAIL.n463 VTAIL.n462 4.26717
R2826 VTAIL.n404 VTAIL.n312 4.26717
R2827 VTAIL.n375 VTAIL.n327 4.26717
R2828 VTAIL.n359 VTAIL.n358 4.26717
R2829 VTAIL.n766 VTAIL.n748 3.49141
R2830 VTAIL.n790 VTAIL.n789 3.49141
R2831 VTAIL.n815 VTAIL.n726 3.49141
R2832 VTAIL.n46 VTAIL.n28 3.49141
R2833 VTAIL.n70 VTAIL.n69 3.49141
R2834 VTAIL.n95 VTAIL.n6 3.49141
R2835 VTAIL.n148 VTAIL.n130 3.49141
R2836 VTAIL.n172 VTAIL.n171 3.49141
R2837 VTAIL.n197 VTAIL.n108 3.49141
R2838 VTAIL.n252 VTAIL.n234 3.49141
R2839 VTAIL.n276 VTAIL.n275 3.49141
R2840 VTAIL.n301 VTAIL.n212 3.49141
R2841 VTAIL.n713 VTAIL.n624 3.49141
R2842 VTAIL.n689 VTAIL.n688 3.49141
R2843 VTAIL.n665 VTAIL.n647 3.49141
R2844 VTAIL.n609 VTAIL.n520 3.49141
R2845 VTAIL.n585 VTAIL.n584 3.49141
R2846 VTAIL.n561 VTAIL.n543 3.49141
R2847 VTAIL.n507 VTAIL.n418 3.49141
R2848 VTAIL.n483 VTAIL.n482 3.49141
R2849 VTAIL.n459 VTAIL.n441 3.49141
R2850 VTAIL.n403 VTAIL.n314 3.49141
R2851 VTAIL.n379 VTAIL.n378 3.49141
R2852 VTAIL.n355 VTAIL.n337 3.49141
R2853 VTAIL.n765 VTAIL.n750 2.71565
R2854 VTAIL.n793 VTAIL.n736 2.71565
R2855 VTAIL.n812 VTAIL.n811 2.71565
R2856 VTAIL.n45 VTAIL.n30 2.71565
R2857 VTAIL.n73 VTAIL.n16 2.71565
R2858 VTAIL.n92 VTAIL.n91 2.71565
R2859 VTAIL.n147 VTAIL.n132 2.71565
R2860 VTAIL.n175 VTAIL.n118 2.71565
R2861 VTAIL.n194 VTAIL.n193 2.71565
R2862 VTAIL.n251 VTAIL.n236 2.71565
R2863 VTAIL.n279 VTAIL.n222 2.71565
R2864 VTAIL.n298 VTAIL.n297 2.71565
R2865 VTAIL.n710 VTAIL.n709 2.71565
R2866 VTAIL.n692 VTAIL.n635 2.71565
R2867 VTAIL.n664 VTAIL.n649 2.71565
R2868 VTAIL.n606 VTAIL.n605 2.71565
R2869 VTAIL.n588 VTAIL.n531 2.71565
R2870 VTAIL.n560 VTAIL.n545 2.71565
R2871 VTAIL.n504 VTAIL.n503 2.71565
R2872 VTAIL.n486 VTAIL.n429 2.71565
R2873 VTAIL.n458 VTAIL.n443 2.71565
R2874 VTAIL.n400 VTAIL.n399 2.71565
R2875 VTAIL.n382 VTAIL.n325 2.71565
R2876 VTAIL.n354 VTAIL.n339 2.71565
R2877 VTAIL.n762 VTAIL.n761 1.93989
R2878 VTAIL.n794 VTAIL.n734 1.93989
R2879 VTAIL.n808 VTAIL.n728 1.93989
R2880 VTAIL.n42 VTAIL.n41 1.93989
R2881 VTAIL.n74 VTAIL.n14 1.93989
R2882 VTAIL.n88 VTAIL.n8 1.93989
R2883 VTAIL.n144 VTAIL.n143 1.93989
R2884 VTAIL.n176 VTAIL.n116 1.93989
R2885 VTAIL.n190 VTAIL.n110 1.93989
R2886 VTAIL.n248 VTAIL.n247 1.93989
R2887 VTAIL.n280 VTAIL.n220 1.93989
R2888 VTAIL.n294 VTAIL.n214 1.93989
R2889 VTAIL.n706 VTAIL.n626 1.93989
R2890 VTAIL.n693 VTAIL.n633 1.93989
R2891 VTAIL.n661 VTAIL.n660 1.93989
R2892 VTAIL.n602 VTAIL.n522 1.93989
R2893 VTAIL.n589 VTAIL.n529 1.93989
R2894 VTAIL.n557 VTAIL.n556 1.93989
R2895 VTAIL.n500 VTAIL.n420 1.93989
R2896 VTAIL.n487 VTAIL.n427 1.93989
R2897 VTAIL.n455 VTAIL.n454 1.93989
R2898 VTAIL.n396 VTAIL.n316 1.93989
R2899 VTAIL.n383 VTAIL.n323 1.93989
R2900 VTAIL.n351 VTAIL.n350 1.93989
R2901 VTAIL.n413 VTAIL.n411 1.91429
R2902 VTAIL.n515 VTAIL.n413 1.91429
R2903 VTAIL.n619 VTAIL.n617 1.91429
R2904 VTAIL.n721 VTAIL.n619 1.91429
R2905 VTAIL.n309 VTAIL.n207 1.91429
R2906 VTAIL.n207 VTAIL.n205 1.91429
R2907 VTAIL.n103 VTAIL.n1 1.91429
R2908 VTAIL VTAIL.n823 1.8561
R2909 VTAIL.n758 VTAIL.n752 1.16414
R2910 VTAIL.n799 VTAIL.n797 1.16414
R2911 VTAIL.n807 VTAIL.n730 1.16414
R2912 VTAIL.n38 VTAIL.n32 1.16414
R2913 VTAIL.n79 VTAIL.n77 1.16414
R2914 VTAIL.n87 VTAIL.n10 1.16414
R2915 VTAIL.n140 VTAIL.n134 1.16414
R2916 VTAIL.n181 VTAIL.n179 1.16414
R2917 VTAIL.n189 VTAIL.n112 1.16414
R2918 VTAIL.n244 VTAIL.n238 1.16414
R2919 VTAIL.n285 VTAIL.n283 1.16414
R2920 VTAIL.n293 VTAIL.n216 1.16414
R2921 VTAIL.n705 VTAIL.n628 1.16414
R2922 VTAIL.n697 VTAIL.n696 1.16414
R2923 VTAIL.n657 VTAIL.n651 1.16414
R2924 VTAIL.n601 VTAIL.n524 1.16414
R2925 VTAIL.n593 VTAIL.n592 1.16414
R2926 VTAIL.n553 VTAIL.n547 1.16414
R2927 VTAIL.n499 VTAIL.n422 1.16414
R2928 VTAIL.n491 VTAIL.n490 1.16414
R2929 VTAIL.n451 VTAIL.n445 1.16414
R2930 VTAIL.n395 VTAIL.n318 1.16414
R2931 VTAIL.n387 VTAIL.n386 1.16414
R2932 VTAIL.n347 VTAIL.n341 1.16414
R2933 VTAIL.n0 VTAIL.t1 1.08424
R2934 VTAIL.n0 VTAIL.t2 1.08424
R2935 VTAIL.n206 VTAIL.t9 1.08424
R2936 VTAIL.n206 VTAIL.t14 1.08424
R2937 VTAIL.n618 VTAIL.t15 1.08424
R2938 VTAIL.n618 VTAIL.t8 1.08424
R2939 VTAIL.n412 VTAIL.t4 1.08424
R2940 VTAIL.n412 VTAIL.t7 1.08424
R2941 VTAIL.n617 VTAIL.n515 0.470328
R2942 VTAIL.n205 VTAIL.n103 0.470328
R2943 VTAIL.n757 VTAIL.n754 0.388379
R2944 VTAIL.n798 VTAIL.n732 0.388379
R2945 VTAIL.n804 VTAIL.n803 0.388379
R2946 VTAIL.n37 VTAIL.n34 0.388379
R2947 VTAIL.n78 VTAIL.n12 0.388379
R2948 VTAIL.n84 VTAIL.n83 0.388379
R2949 VTAIL.n139 VTAIL.n136 0.388379
R2950 VTAIL.n180 VTAIL.n114 0.388379
R2951 VTAIL.n186 VTAIL.n185 0.388379
R2952 VTAIL.n243 VTAIL.n240 0.388379
R2953 VTAIL.n284 VTAIL.n218 0.388379
R2954 VTAIL.n290 VTAIL.n289 0.388379
R2955 VTAIL.n702 VTAIL.n701 0.388379
R2956 VTAIL.n632 VTAIL.n630 0.388379
R2957 VTAIL.n656 VTAIL.n653 0.388379
R2958 VTAIL.n598 VTAIL.n597 0.388379
R2959 VTAIL.n528 VTAIL.n526 0.388379
R2960 VTAIL.n552 VTAIL.n549 0.388379
R2961 VTAIL.n496 VTAIL.n495 0.388379
R2962 VTAIL.n426 VTAIL.n424 0.388379
R2963 VTAIL.n450 VTAIL.n447 0.388379
R2964 VTAIL.n392 VTAIL.n391 0.388379
R2965 VTAIL.n322 VTAIL.n320 0.388379
R2966 VTAIL.n346 VTAIL.n343 0.388379
R2967 VTAIL.n756 VTAIL.n751 0.155672
R2968 VTAIL.n763 VTAIL.n751 0.155672
R2969 VTAIL.n764 VTAIL.n763 0.155672
R2970 VTAIL.n764 VTAIL.n747 0.155672
R2971 VTAIL.n771 VTAIL.n747 0.155672
R2972 VTAIL.n772 VTAIL.n771 0.155672
R2973 VTAIL.n772 VTAIL.n743 0.155672
R2974 VTAIL.n779 VTAIL.n743 0.155672
R2975 VTAIL.n780 VTAIL.n779 0.155672
R2976 VTAIL.n780 VTAIL.n739 0.155672
R2977 VTAIL.n787 VTAIL.n739 0.155672
R2978 VTAIL.n788 VTAIL.n787 0.155672
R2979 VTAIL.n788 VTAIL.n735 0.155672
R2980 VTAIL.n795 VTAIL.n735 0.155672
R2981 VTAIL.n796 VTAIL.n795 0.155672
R2982 VTAIL.n796 VTAIL.n731 0.155672
R2983 VTAIL.n805 VTAIL.n731 0.155672
R2984 VTAIL.n806 VTAIL.n805 0.155672
R2985 VTAIL.n806 VTAIL.n727 0.155672
R2986 VTAIL.n813 VTAIL.n727 0.155672
R2987 VTAIL.n814 VTAIL.n813 0.155672
R2988 VTAIL.n814 VTAIL.n723 0.155672
R2989 VTAIL.n821 VTAIL.n723 0.155672
R2990 VTAIL.n36 VTAIL.n31 0.155672
R2991 VTAIL.n43 VTAIL.n31 0.155672
R2992 VTAIL.n44 VTAIL.n43 0.155672
R2993 VTAIL.n44 VTAIL.n27 0.155672
R2994 VTAIL.n51 VTAIL.n27 0.155672
R2995 VTAIL.n52 VTAIL.n51 0.155672
R2996 VTAIL.n52 VTAIL.n23 0.155672
R2997 VTAIL.n59 VTAIL.n23 0.155672
R2998 VTAIL.n60 VTAIL.n59 0.155672
R2999 VTAIL.n60 VTAIL.n19 0.155672
R3000 VTAIL.n67 VTAIL.n19 0.155672
R3001 VTAIL.n68 VTAIL.n67 0.155672
R3002 VTAIL.n68 VTAIL.n15 0.155672
R3003 VTAIL.n75 VTAIL.n15 0.155672
R3004 VTAIL.n76 VTAIL.n75 0.155672
R3005 VTAIL.n76 VTAIL.n11 0.155672
R3006 VTAIL.n85 VTAIL.n11 0.155672
R3007 VTAIL.n86 VTAIL.n85 0.155672
R3008 VTAIL.n86 VTAIL.n7 0.155672
R3009 VTAIL.n93 VTAIL.n7 0.155672
R3010 VTAIL.n94 VTAIL.n93 0.155672
R3011 VTAIL.n94 VTAIL.n3 0.155672
R3012 VTAIL.n101 VTAIL.n3 0.155672
R3013 VTAIL.n138 VTAIL.n133 0.155672
R3014 VTAIL.n145 VTAIL.n133 0.155672
R3015 VTAIL.n146 VTAIL.n145 0.155672
R3016 VTAIL.n146 VTAIL.n129 0.155672
R3017 VTAIL.n153 VTAIL.n129 0.155672
R3018 VTAIL.n154 VTAIL.n153 0.155672
R3019 VTAIL.n154 VTAIL.n125 0.155672
R3020 VTAIL.n161 VTAIL.n125 0.155672
R3021 VTAIL.n162 VTAIL.n161 0.155672
R3022 VTAIL.n162 VTAIL.n121 0.155672
R3023 VTAIL.n169 VTAIL.n121 0.155672
R3024 VTAIL.n170 VTAIL.n169 0.155672
R3025 VTAIL.n170 VTAIL.n117 0.155672
R3026 VTAIL.n177 VTAIL.n117 0.155672
R3027 VTAIL.n178 VTAIL.n177 0.155672
R3028 VTAIL.n178 VTAIL.n113 0.155672
R3029 VTAIL.n187 VTAIL.n113 0.155672
R3030 VTAIL.n188 VTAIL.n187 0.155672
R3031 VTAIL.n188 VTAIL.n109 0.155672
R3032 VTAIL.n195 VTAIL.n109 0.155672
R3033 VTAIL.n196 VTAIL.n195 0.155672
R3034 VTAIL.n196 VTAIL.n105 0.155672
R3035 VTAIL.n203 VTAIL.n105 0.155672
R3036 VTAIL.n242 VTAIL.n237 0.155672
R3037 VTAIL.n249 VTAIL.n237 0.155672
R3038 VTAIL.n250 VTAIL.n249 0.155672
R3039 VTAIL.n250 VTAIL.n233 0.155672
R3040 VTAIL.n257 VTAIL.n233 0.155672
R3041 VTAIL.n258 VTAIL.n257 0.155672
R3042 VTAIL.n258 VTAIL.n229 0.155672
R3043 VTAIL.n265 VTAIL.n229 0.155672
R3044 VTAIL.n266 VTAIL.n265 0.155672
R3045 VTAIL.n266 VTAIL.n225 0.155672
R3046 VTAIL.n273 VTAIL.n225 0.155672
R3047 VTAIL.n274 VTAIL.n273 0.155672
R3048 VTAIL.n274 VTAIL.n221 0.155672
R3049 VTAIL.n281 VTAIL.n221 0.155672
R3050 VTAIL.n282 VTAIL.n281 0.155672
R3051 VTAIL.n282 VTAIL.n217 0.155672
R3052 VTAIL.n291 VTAIL.n217 0.155672
R3053 VTAIL.n292 VTAIL.n291 0.155672
R3054 VTAIL.n292 VTAIL.n213 0.155672
R3055 VTAIL.n299 VTAIL.n213 0.155672
R3056 VTAIL.n300 VTAIL.n299 0.155672
R3057 VTAIL.n300 VTAIL.n209 0.155672
R3058 VTAIL.n307 VTAIL.n209 0.155672
R3059 VTAIL.n719 VTAIL.n621 0.155672
R3060 VTAIL.n712 VTAIL.n621 0.155672
R3061 VTAIL.n712 VTAIL.n711 0.155672
R3062 VTAIL.n711 VTAIL.n625 0.155672
R3063 VTAIL.n704 VTAIL.n625 0.155672
R3064 VTAIL.n704 VTAIL.n703 0.155672
R3065 VTAIL.n703 VTAIL.n629 0.155672
R3066 VTAIL.n695 VTAIL.n629 0.155672
R3067 VTAIL.n695 VTAIL.n694 0.155672
R3068 VTAIL.n694 VTAIL.n634 0.155672
R3069 VTAIL.n687 VTAIL.n634 0.155672
R3070 VTAIL.n687 VTAIL.n686 0.155672
R3071 VTAIL.n686 VTAIL.n638 0.155672
R3072 VTAIL.n679 VTAIL.n638 0.155672
R3073 VTAIL.n679 VTAIL.n678 0.155672
R3074 VTAIL.n678 VTAIL.n642 0.155672
R3075 VTAIL.n671 VTAIL.n642 0.155672
R3076 VTAIL.n671 VTAIL.n670 0.155672
R3077 VTAIL.n670 VTAIL.n646 0.155672
R3078 VTAIL.n663 VTAIL.n646 0.155672
R3079 VTAIL.n663 VTAIL.n662 0.155672
R3080 VTAIL.n662 VTAIL.n650 0.155672
R3081 VTAIL.n655 VTAIL.n650 0.155672
R3082 VTAIL.n615 VTAIL.n517 0.155672
R3083 VTAIL.n608 VTAIL.n517 0.155672
R3084 VTAIL.n608 VTAIL.n607 0.155672
R3085 VTAIL.n607 VTAIL.n521 0.155672
R3086 VTAIL.n600 VTAIL.n521 0.155672
R3087 VTAIL.n600 VTAIL.n599 0.155672
R3088 VTAIL.n599 VTAIL.n525 0.155672
R3089 VTAIL.n591 VTAIL.n525 0.155672
R3090 VTAIL.n591 VTAIL.n590 0.155672
R3091 VTAIL.n590 VTAIL.n530 0.155672
R3092 VTAIL.n583 VTAIL.n530 0.155672
R3093 VTAIL.n583 VTAIL.n582 0.155672
R3094 VTAIL.n582 VTAIL.n534 0.155672
R3095 VTAIL.n575 VTAIL.n534 0.155672
R3096 VTAIL.n575 VTAIL.n574 0.155672
R3097 VTAIL.n574 VTAIL.n538 0.155672
R3098 VTAIL.n567 VTAIL.n538 0.155672
R3099 VTAIL.n567 VTAIL.n566 0.155672
R3100 VTAIL.n566 VTAIL.n542 0.155672
R3101 VTAIL.n559 VTAIL.n542 0.155672
R3102 VTAIL.n559 VTAIL.n558 0.155672
R3103 VTAIL.n558 VTAIL.n546 0.155672
R3104 VTAIL.n551 VTAIL.n546 0.155672
R3105 VTAIL.n513 VTAIL.n415 0.155672
R3106 VTAIL.n506 VTAIL.n415 0.155672
R3107 VTAIL.n506 VTAIL.n505 0.155672
R3108 VTAIL.n505 VTAIL.n419 0.155672
R3109 VTAIL.n498 VTAIL.n419 0.155672
R3110 VTAIL.n498 VTAIL.n497 0.155672
R3111 VTAIL.n497 VTAIL.n423 0.155672
R3112 VTAIL.n489 VTAIL.n423 0.155672
R3113 VTAIL.n489 VTAIL.n488 0.155672
R3114 VTAIL.n488 VTAIL.n428 0.155672
R3115 VTAIL.n481 VTAIL.n428 0.155672
R3116 VTAIL.n481 VTAIL.n480 0.155672
R3117 VTAIL.n480 VTAIL.n432 0.155672
R3118 VTAIL.n473 VTAIL.n432 0.155672
R3119 VTAIL.n473 VTAIL.n472 0.155672
R3120 VTAIL.n472 VTAIL.n436 0.155672
R3121 VTAIL.n465 VTAIL.n436 0.155672
R3122 VTAIL.n465 VTAIL.n464 0.155672
R3123 VTAIL.n464 VTAIL.n440 0.155672
R3124 VTAIL.n457 VTAIL.n440 0.155672
R3125 VTAIL.n457 VTAIL.n456 0.155672
R3126 VTAIL.n456 VTAIL.n444 0.155672
R3127 VTAIL.n449 VTAIL.n444 0.155672
R3128 VTAIL.n409 VTAIL.n311 0.155672
R3129 VTAIL.n402 VTAIL.n311 0.155672
R3130 VTAIL.n402 VTAIL.n401 0.155672
R3131 VTAIL.n401 VTAIL.n315 0.155672
R3132 VTAIL.n394 VTAIL.n315 0.155672
R3133 VTAIL.n394 VTAIL.n393 0.155672
R3134 VTAIL.n393 VTAIL.n319 0.155672
R3135 VTAIL.n385 VTAIL.n319 0.155672
R3136 VTAIL.n385 VTAIL.n384 0.155672
R3137 VTAIL.n384 VTAIL.n324 0.155672
R3138 VTAIL.n377 VTAIL.n324 0.155672
R3139 VTAIL.n377 VTAIL.n376 0.155672
R3140 VTAIL.n376 VTAIL.n328 0.155672
R3141 VTAIL.n369 VTAIL.n328 0.155672
R3142 VTAIL.n369 VTAIL.n368 0.155672
R3143 VTAIL.n368 VTAIL.n332 0.155672
R3144 VTAIL.n361 VTAIL.n332 0.155672
R3145 VTAIL.n361 VTAIL.n360 0.155672
R3146 VTAIL.n360 VTAIL.n336 0.155672
R3147 VTAIL.n353 VTAIL.n336 0.155672
R3148 VTAIL.n353 VTAIL.n352 0.155672
R3149 VTAIL.n352 VTAIL.n340 0.155672
R3150 VTAIL.n345 VTAIL.n340 0.155672
R3151 VTAIL VTAIL.n1 0.0586897
R3152 VDD1 VDD1.n0 62.2452
R3153 VDD1.n3 VDD1.n2 62.1315
R3154 VDD1.n3 VDD1.n1 62.1315
R3155 VDD1.n5 VDD1.n4 61.2299
R3156 VDD1.n5 VDD1.n3 48.6604
R3157 VDD1.n4 VDD1.t2 1.08424
R3158 VDD1.n4 VDD1.t7 1.08424
R3159 VDD1.n0 VDD1.t4 1.08424
R3160 VDD1.n0 VDD1.t1 1.08424
R3161 VDD1.n2 VDD1.t3 1.08424
R3162 VDD1.n2 VDD1.t6 1.08424
R3163 VDD1.n1 VDD1.t5 1.08424
R3164 VDD1.n1 VDD1.t0 1.08424
R3165 VDD1 VDD1.n5 0.899207
R3166 VN.n5 VN.t3 267.307
R3167 VN.n28 VN.t6 267.307
R3168 VN.n6 VN.t5 232.968
R3169 VN.n13 VN.t2 232.968
R3170 VN.n21 VN.t4 232.968
R3171 VN.n29 VN.t0 232.968
R3172 VN.n36 VN.t7 232.968
R3173 VN.n44 VN.t1 232.968
R3174 VN.n22 VN.n21 181.852
R3175 VN.n45 VN.n44 181.852
R3176 VN.n43 VN.n23 161.3
R3177 VN.n42 VN.n41 161.3
R3178 VN.n40 VN.n24 161.3
R3179 VN.n39 VN.n38 161.3
R3180 VN.n37 VN.n25 161.3
R3181 VN.n35 VN.n34 161.3
R3182 VN.n33 VN.n26 161.3
R3183 VN.n32 VN.n31 161.3
R3184 VN.n30 VN.n27 161.3
R3185 VN.n20 VN.n0 161.3
R3186 VN.n19 VN.n18 161.3
R3187 VN.n17 VN.n1 161.3
R3188 VN.n16 VN.n15 161.3
R3189 VN.n14 VN.n2 161.3
R3190 VN.n12 VN.n11 161.3
R3191 VN.n10 VN.n3 161.3
R3192 VN.n9 VN.n8 161.3
R3193 VN.n7 VN.n4 161.3
R3194 VN.n8 VN.n3 56.5193
R3195 VN.n31 VN.n26 56.5193
R3196 VN VN.n45 52.6312
R3197 VN.n6 VN.n5 52.0405
R3198 VN.n29 VN.n28 52.0405
R3199 VN.n15 VN.n1 43.4072
R3200 VN.n38 VN.n24 43.4072
R3201 VN.n19 VN.n1 37.5796
R3202 VN.n42 VN.n24 37.5796
R3203 VN.n8 VN.n7 24.4675
R3204 VN.n12 VN.n3 24.4675
R3205 VN.n15 VN.n14 24.4675
R3206 VN.n20 VN.n19 24.4675
R3207 VN.n31 VN.n30 24.4675
R3208 VN.n38 VN.n37 24.4675
R3209 VN.n35 VN.n26 24.4675
R3210 VN.n43 VN.n42 24.4675
R3211 VN.n7 VN.n6 17.6167
R3212 VN.n13 VN.n12 17.6167
R3213 VN.n30 VN.n29 17.6167
R3214 VN.n36 VN.n35 17.6167
R3215 VN.n28 VN.n27 12.2976
R3216 VN.n5 VN.n4 12.2976
R3217 VN.n14 VN.n13 6.85126
R3218 VN.n37 VN.n36 6.85126
R3219 VN.n21 VN.n20 3.91522
R3220 VN.n44 VN.n43 3.91522
R3221 VN.n45 VN.n23 0.189894
R3222 VN.n41 VN.n23 0.189894
R3223 VN.n41 VN.n40 0.189894
R3224 VN.n40 VN.n39 0.189894
R3225 VN.n39 VN.n25 0.189894
R3226 VN.n34 VN.n25 0.189894
R3227 VN.n34 VN.n33 0.189894
R3228 VN.n33 VN.n32 0.189894
R3229 VN.n32 VN.n27 0.189894
R3230 VN.n9 VN.n4 0.189894
R3231 VN.n10 VN.n9 0.189894
R3232 VN.n11 VN.n10 0.189894
R3233 VN.n11 VN.n2 0.189894
R3234 VN.n16 VN.n2 0.189894
R3235 VN.n17 VN.n16 0.189894
R3236 VN.n18 VN.n17 0.189894
R3237 VN.n18 VN.n0 0.189894
R3238 VN.n22 VN.n0 0.189894
R3239 VN VN.n22 0.0516364
R3240 VDD2.n2 VDD2.n1 62.1315
R3241 VDD2.n2 VDD2.n0 62.1315
R3242 VDD2 VDD2.n5 62.1286
R3243 VDD2.n4 VDD2.n3 61.2301
R3244 VDD2.n4 VDD2.n2 48.0774
R3245 VDD2.n5 VDD2.t7 1.08424
R3246 VDD2.n5 VDD2.t1 1.08424
R3247 VDD2.n3 VDD2.t6 1.08424
R3248 VDD2.n3 VDD2.t0 1.08424
R3249 VDD2.n1 VDD2.t5 1.08424
R3250 VDD2.n1 VDD2.t3 1.08424
R3251 VDD2.n0 VDD2.t4 1.08424
R3252 VDD2.n0 VDD2.t2 1.08424
R3253 VDD2 VDD2.n4 1.01559
C0 VN VDD2 12.094f
C1 VTAIL VDD1 10.6745f
C2 VTAIL VDD2 10.7242f
C3 VDD1 VP 12.3867f
C4 VDD2 VP 0.443706f
C5 VN VTAIL 11.9922f
C6 VDD1 VDD2 1.40507f
C7 VN VP 7.953f
C8 VTAIL VP 12.0063f
C9 VN VDD1 0.150031f
C10 VDD2 B 5.146651f
C11 VDD1 B 5.507319f
C12 VTAIL B 13.688592f
C13 VN B 13.389291f
C14 VP B 11.712229f
C15 VDD2.t4 B 0.356164f
C16 VDD2.t2 B 0.356164f
C17 VDD2.n0 B 3.25331f
C18 VDD2.t5 B 0.356164f
C19 VDD2.t3 B 0.356164f
C20 VDD2.n1 B 3.25331f
C21 VDD2.n2 B 3.22017f
C22 VDD2.t6 B 0.356164f
C23 VDD2.t0 B 0.356164f
C24 VDD2.n3 B 3.24695f
C25 VDD2.n4 B 3.13959f
C26 VDD2.t7 B 0.356164f
C27 VDD2.t1 B 0.356164f
C28 VDD2.n5 B 3.25328f
C29 VN.n0 B 0.026187f
C30 VN.t4 B 2.48789f
C31 VN.n1 B 0.021474f
C32 VN.n2 B 0.026187f
C33 VN.t2 B 2.48789f
C34 VN.n3 B 0.038229f
C35 VN.n4 B 0.194848f
C36 VN.t5 B 2.48789f
C37 VN.t3 B 2.61605f
C38 VN.n5 B 0.929475f
C39 VN.n6 B 0.934063f
C40 VN.n7 B 0.042059f
C41 VN.n8 B 0.038229f
C42 VN.n9 B 0.026187f
C43 VN.n10 B 0.026187f
C44 VN.n11 B 0.026187f
C45 VN.n12 B 0.042059f
C46 VN.n13 B 0.868806f
C47 VN.n14 B 0.031457f
C48 VN.n15 B 0.051117f
C49 VN.n16 B 0.026187f
C50 VN.n17 B 0.026187f
C51 VN.n18 B 0.026187f
C52 VN.n19 B 0.052672f
C53 VN.n20 B 0.028566f
C54 VN.n21 B 0.932186f
C55 VN.n22 B 0.02837f
C56 VN.n23 B 0.026187f
C57 VN.t1 B 2.48789f
C58 VN.n24 B 0.021474f
C59 VN.n25 B 0.026187f
C60 VN.t7 B 2.48789f
C61 VN.n26 B 0.038229f
C62 VN.n27 B 0.194848f
C63 VN.t0 B 2.48789f
C64 VN.t6 B 2.61605f
C65 VN.n28 B 0.929475f
C66 VN.n29 B 0.934063f
C67 VN.n30 B 0.042059f
C68 VN.n31 B 0.038229f
C69 VN.n32 B 0.026187f
C70 VN.n33 B 0.026187f
C71 VN.n34 B 0.026187f
C72 VN.n35 B 0.042059f
C73 VN.n36 B 0.868806f
C74 VN.n37 B 0.031457f
C75 VN.n38 B 0.051117f
C76 VN.n39 B 0.026187f
C77 VN.n40 B 0.026187f
C78 VN.n41 B 0.026187f
C79 VN.n42 B 0.052672f
C80 VN.n43 B 0.028566f
C81 VN.n44 B 0.932186f
C82 VN.n45 B 1.5451f
C83 VDD1.t4 B 0.359414f
C84 VDD1.t1 B 0.359414f
C85 VDD1.n0 B 3.28395f
C86 VDD1.t5 B 0.359414f
C87 VDD1.t0 B 0.359414f
C88 VDD1.n1 B 3.283f
C89 VDD1.t3 B 0.359414f
C90 VDD1.t6 B 0.359414f
C91 VDD1.n2 B 3.283f
C92 VDD1.n3 B 3.30153f
C93 VDD1.t2 B 0.359414f
C94 VDD1.t7 B 0.359414f
C95 VDD1.n4 B 3.27657f
C96 VDD1.n5 B 3.19888f
C97 VTAIL.t1 B 0.264305f
C98 VTAIL.t2 B 0.264305f
C99 VTAIL.n0 B 2.35393f
C100 VTAIL.n1 B 0.298996f
C101 VTAIL.n2 B 0.026102f
C102 VTAIL.n3 B 0.018307f
C103 VTAIL.n4 B 0.009837f
C104 VTAIL.n5 B 0.023252f
C105 VTAIL.n6 B 0.010416f
C106 VTAIL.n7 B 0.018307f
C107 VTAIL.n8 B 0.009837f
C108 VTAIL.n9 B 0.023252f
C109 VTAIL.n10 B 0.010416f
C110 VTAIL.n11 B 0.018307f
C111 VTAIL.n12 B 0.010127f
C112 VTAIL.n13 B 0.023252f
C113 VTAIL.n14 B 0.010416f
C114 VTAIL.n15 B 0.018307f
C115 VTAIL.n16 B 0.009837f
C116 VTAIL.n17 B 0.023252f
C117 VTAIL.n18 B 0.010416f
C118 VTAIL.n19 B 0.018307f
C119 VTAIL.n20 B 0.009837f
C120 VTAIL.n21 B 0.023252f
C121 VTAIL.n22 B 0.010416f
C122 VTAIL.n23 B 0.018307f
C123 VTAIL.n24 B 0.009837f
C124 VTAIL.n25 B 0.023252f
C125 VTAIL.n26 B 0.010416f
C126 VTAIL.n27 B 0.018307f
C127 VTAIL.n28 B 0.009837f
C128 VTAIL.n29 B 0.023252f
C129 VTAIL.n30 B 0.010416f
C130 VTAIL.n31 B 0.018307f
C131 VTAIL.n32 B 0.009837f
C132 VTAIL.n33 B 0.017439f
C133 VTAIL.n34 B 0.013736f
C134 VTAIL.t5 B 0.038545f
C135 VTAIL.n35 B 0.13441f
C136 VTAIL.n36 B 1.46542f
C137 VTAIL.n37 B 0.009837f
C138 VTAIL.n38 B 0.010416f
C139 VTAIL.n39 B 0.023252f
C140 VTAIL.n40 B 0.023252f
C141 VTAIL.n41 B 0.010416f
C142 VTAIL.n42 B 0.009837f
C143 VTAIL.n43 B 0.018307f
C144 VTAIL.n44 B 0.018307f
C145 VTAIL.n45 B 0.009837f
C146 VTAIL.n46 B 0.010416f
C147 VTAIL.n47 B 0.023252f
C148 VTAIL.n48 B 0.023252f
C149 VTAIL.n49 B 0.010416f
C150 VTAIL.n50 B 0.009837f
C151 VTAIL.n51 B 0.018307f
C152 VTAIL.n52 B 0.018307f
C153 VTAIL.n53 B 0.009837f
C154 VTAIL.n54 B 0.010416f
C155 VTAIL.n55 B 0.023252f
C156 VTAIL.n56 B 0.023252f
C157 VTAIL.n57 B 0.010416f
C158 VTAIL.n58 B 0.009837f
C159 VTAIL.n59 B 0.018307f
C160 VTAIL.n60 B 0.018307f
C161 VTAIL.n61 B 0.009837f
C162 VTAIL.n62 B 0.010416f
C163 VTAIL.n63 B 0.023252f
C164 VTAIL.n64 B 0.023252f
C165 VTAIL.n65 B 0.010416f
C166 VTAIL.n66 B 0.009837f
C167 VTAIL.n67 B 0.018307f
C168 VTAIL.n68 B 0.018307f
C169 VTAIL.n69 B 0.009837f
C170 VTAIL.n70 B 0.010416f
C171 VTAIL.n71 B 0.023252f
C172 VTAIL.n72 B 0.023252f
C173 VTAIL.n73 B 0.010416f
C174 VTAIL.n74 B 0.009837f
C175 VTAIL.n75 B 0.018307f
C176 VTAIL.n76 B 0.018307f
C177 VTAIL.n77 B 0.009837f
C178 VTAIL.n78 B 0.009837f
C179 VTAIL.n79 B 0.010416f
C180 VTAIL.n80 B 0.023252f
C181 VTAIL.n81 B 0.023252f
C182 VTAIL.n82 B 0.023252f
C183 VTAIL.n83 B 0.010127f
C184 VTAIL.n84 B 0.009837f
C185 VTAIL.n85 B 0.018307f
C186 VTAIL.n86 B 0.018307f
C187 VTAIL.n87 B 0.009837f
C188 VTAIL.n88 B 0.010416f
C189 VTAIL.n89 B 0.023252f
C190 VTAIL.n90 B 0.023252f
C191 VTAIL.n91 B 0.010416f
C192 VTAIL.n92 B 0.009837f
C193 VTAIL.n93 B 0.018307f
C194 VTAIL.n94 B 0.018307f
C195 VTAIL.n95 B 0.009837f
C196 VTAIL.n96 B 0.010416f
C197 VTAIL.n97 B 0.023252f
C198 VTAIL.n98 B 0.050991f
C199 VTAIL.n99 B 0.010416f
C200 VTAIL.n100 B 0.009837f
C201 VTAIL.n101 B 0.043066f
C202 VTAIL.n102 B 0.028622f
C203 VTAIL.n103 B 0.156666f
C204 VTAIL.n104 B 0.026102f
C205 VTAIL.n105 B 0.018307f
C206 VTAIL.n106 B 0.009837f
C207 VTAIL.n107 B 0.023252f
C208 VTAIL.n108 B 0.010416f
C209 VTAIL.n109 B 0.018307f
C210 VTAIL.n110 B 0.009837f
C211 VTAIL.n111 B 0.023252f
C212 VTAIL.n112 B 0.010416f
C213 VTAIL.n113 B 0.018307f
C214 VTAIL.n114 B 0.010127f
C215 VTAIL.n115 B 0.023252f
C216 VTAIL.n116 B 0.010416f
C217 VTAIL.n117 B 0.018307f
C218 VTAIL.n118 B 0.009837f
C219 VTAIL.n119 B 0.023252f
C220 VTAIL.n120 B 0.010416f
C221 VTAIL.n121 B 0.018307f
C222 VTAIL.n122 B 0.009837f
C223 VTAIL.n123 B 0.023252f
C224 VTAIL.n124 B 0.010416f
C225 VTAIL.n125 B 0.018307f
C226 VTAIL.n126 B 0.009837f
C227 VTAIL.n127 B 0.023252f
C228 VTAIL.n128 B 0.010416f
C229 VTAIL.n129 B 0.018307f
C230 VTAIL.n130 B 0.009837f
C231 VTAIL.n131 B 0.023252f
C232 VTAIL.n132 B 0.010416f
C233 VTAIL.n133 B 0.018307f
C234 VTAIL.n134 B 0.009837f
C235 VTAIL.n135 B 0.017439f
C236 VTAIL.n136 B 0.013736f
C237 VTAIL.t13 B 0.038545f
C238 VTAIL.n137 B 0.13441f
C239 VTAIL.n138 B 1.46542f
C240 VTAIL.n139 B 0.009837f
C241 VTAIL.n140 B 0.010416f
C242 VTAIL.n141 B 0.023252f
C243 VTAIL.n142 B 0.023252f
C244 VTAIL.n143 B 0.010416f
C245 VTAIL.n144 B 0.009837f
C246 VTAIL.n145 B 0.018307f
C247 VTAIL.n146 B 0.018307f
C248 VTAIL.n147 B 0.009837f
C249 VTAIL.n148 B 0.010416f
C250 VTAIL.n149 B 0.023252f
C251 VTAIL.n150 B 0.023252f
C252 VTAIL.n151 B 0.010416f
C253 VTAIL.n152 B 0.009837f
C254 VTAIL.n153 B 0.018307f
C255 VTAIL.n154 B 0.018307f
C256 VTAIL.n155 B 0.009837f
C257 VTAIL.n156 B 0.010416f
C258 VTAIL.n157 B 0.023252f
C259 VTAIL.n158 B 0.023252f
C260 VTAIL.n159 B 0.010416f
C261 VTAIL.n160 B 0.009837f
C262 VTAIL.n161 B 0.018307f
C263 VTAIL.n162 B 0.018307f
C264 VTAIL.n163 B 0.009837f
C265 VTAIL.n164 B 0.010416f
C266 VTAIL.n165 B 0.023252f
C267 VTAIL.n166 B 0.023252f
C268 VTAIL.n167 B 0.010416f
C269 VTAIL.n168 B 0.009837f
C270 VTAIL.n169 B 0.018307f
C271 VTAIL.n170 B 0.018307f
C272 VTAIL.n171 B 0.009837f
C273 VTAIL.n172 B 0.010416f
C274 VTAIL.n173 B 0.023252f
C275 VTAIL.n174 B 0.023252f
C276 VTAIL.n175 B 0.010416f
C277 VTAIL.n176 B 0.009837f
C278 VTAIL.n177 B 0.018307f
C279 VTAIL.n178 B 0.018307f
C280 VTAIL.n179 B 0.009837f
C281 VTAIL.n180 B 0.009837f
C282 VTAIL.n181 B 0.010416f
C283 VTAIL.n182 B 0.023252f
C284 VTAIL.n183 B 0.023252f
C285 VTAIL.n184 B 0.023252f
C286 VTAIL.n185 B 0.010127f
C287 VTAIL.n186 B 0.009837f
C288 VTAIL.n187 B 0.018307f
C289 VTAIL.n188 B 0.018307f
C290 VTAIL.n189 B 0.009837f
C291 VTAIL.n190 B 0.010416f
C292 VTAIL.n191 B 0.023252f
C293 VTAIL.n192 B 0.023252f
C294 VTAIL.n193 B 0.010416f
C295 VTAIL.n194 B 0.009837f
C296 VTAIL.n195 B 0.018307f
C297 VTAIL.n196 B 0.018307f
C298 VTAIL.n197 B 0.009837f
C299 VTAIL.n198 B 0.010416f
C300 VTAIL.n199 B 0.023252f
C301 VTAIL.n200 B 0.050991f
C302 VTAIL.n201 B 0.010416f
C303 VTAIL.n202 B 0.009837f
C304 VTAIL.n203 B 0.043066f
C305 VTAIL.n204 B 0.028622f
C306 VTAIL.n205 B 0.156666f
C307 VTAIL.t9 B 0.264305f
C308 VTAIL.t14 B 0.264305f
C309 VTAIL.n206 B 2.35393f
C310 VTAIL.n207 B 0.408455f
C311 VTAIL.n208 B 0.026102f
C312 VTAIL.n209 B 0.018307f
C313 VTAIL.n210 B 0.009837f
C314 VTAIL.n211 B 0.023252f
C315 VTAIL.n212 B 0.010416f
C316 VTAIL.n213 B 0.018307f
C317 VTAIL.n214 B 0.009837f
C318 VTAIL.n215 B 0.023252f
C319 VTAIL.n216 B 0.010416f
C320 VTAIL.n217 B 0.018307f
C321 VTAIL.n218 B 0.010127f
C322 VTAIL.n219 B 0.023252f
C323 VTAIL.n220 B 0.010416f
C324 VTAIL.n221 B 0.018307f
C325 VTAIL.n222 B 0.009837f
C326 VTAIL.n223 B 0.023252f
C327 VTAIL.n224 B 0.010416f
C328 VTAIL.n225 B 0.018307f
C329 VTAIL.n226 B 0.009837f
C330 VTAIL.n227 B 0.023252f
C331 VTAIL.n228 B 0.010416f
C332 VTAIL.n229 B 0.018307f
C333 VTAIL.n230 B 0.009837f
C334 VTAIL.n231 B 0.023252f
C335 VTAIL.n232 B 0.010416f
C336 VTAIL.n233 B 0.018307f
C337 VTAIL.n234 B 0.009837f
C338 VTAIL.n235 B 0.023252f
C339 VTAIL.n236 B 0.010416f
C340 VTAIL.n237 B 0.018307f
C341 VTAIL.n238 B 0.009837f
C342 VTAIL.n239 B 0.017439f
C343 VTAIL.n240 B 0.013736f
C344 VTAIL.t10 B 0.038545f
C345 VTAIL.n241 B 0.13441f
C346 VTAIL.n242 B 1.46542f
C347 VTAIL.n243 B 0.009837f
C348 VTAIL.n244 B 0.010416f
C349 VTAIL.n245 B 0.023252f
C350 VTAIL.n246 B 0.023252f
C351 VTAIL.n247 B 0.010416f
C352 VTAIL.n248 B 0.009837f
C353 VTAIL.n249 B 0.018307f
C354 VTAIL.n250 B 0.018307f
C355 VTAIL.n251 B 0.009837f
C356 VTAIL.n252 B 0.010416f
C357 VTAIL.n253 B 0.023252f
C358 VTAIL.n254 B 0.023252f
C359 VTAIL.n255 B 0.010416f
C360 VTAIL.n256 B 0.009837f
C361 VTAIL.n257 B 0.018307f
C362 VTAIL.n258 B 0.018307f
C363 VTAIL.n259 B 0.009837f
C364 VTAIL.n260 B 0.010416f
C365 VTAIL.n261 B 0.023252f
C366 VTAIL.n262 B 0.023252f
C367 VTAIL.n263 B 0.010416f
C368 VTAIL.n264 B 0.009837f
C369 VTAIL.n265 B 0.018307f
C370 VTAIL.n266 B 0.018307f
C371 VTAIL.n267 B 0.009837f
C372 VTAIL.n268 B 0.010416f
C373 VTAIL.n269 B 0.023252f
C374 VTAIL.n270 B 0.023252f
C375 VTAIL.n271 B 0.010416f
C376 VTAIL.n272 B 0.009837f
C377 VTAIL.n273 B 0.018307f
C378 VTAIL.n274 B 0.018307f
C379 VTAIL.n275 B 0.009837f
C380 VTAIL.n276 B 0.010416f
C381 VTAIL.n277 B 0.023252f
C382 VTAIL.n278 B 0.023252f
C383 VTAIL.n279 B 0.010416f
C384 VTAIL.n280 B 0.009837f
C385 VTAIL.n281 B 0.018307f
C386 VTAIL.n282 B 0.018307f
C387 VTAIL.n283 B 0.009837f
C388 VTAIL.n284 B 0.009837f
C389 VTAIL.n285 B 0.010416f
C390 VTAIL.n286 B 0.023252f
C391 VTAIL.n287 B 0.023252f
C392 VTAIL.n288 B 0.023252f
C393 VTAIL.n289 B 0.010127f
C394 VTAIL.n290 B 0.009837f
C395 VTAIL.n291 B 0.018307f
C396 VTAIL.n292 B 0.018307f
C397 VTAIL.n293 B 0.009837f
C398 VTAIL.n294 B 0.010416f
C399 VTAIL.n295 B 0.023252f
C400 VTAIL.n296 B 0.023252f
C401 VTAIL.n297 B 0.010416f
C402 VTAIL.n298 B 0.009837f
C403 VTAIL.n299 B 0.018307f
C404 VTAIL.n300 B 0.018307f
C405 VTAIL.n301 B 0.009837f
C406 VTAIL.n302 B 0.010416f
C407 VTAIL.n303 B 0.023252f
C408 VTAIL.n304 B 0.050991f
C409 VTAIL.n305 B 0.010416f
C410 VTAIL.n306 B 0.009837f
C411 VTAIL.n307 B 0.043066f
C412 VTAIL.n308 B 0.028622f
C413 VTAIL.n309 B 1.41959f
C414 VTAIL.n310 B 0.026102f
C415 VTAIL.n311 B 0.018307f
C416 VTAIL.n312 B 0.009837f
C417 VTAIL.n313 B 0.023252f
C418 VTAIL.n314 B 0.010416f
C419 VTAIL.n315 B 0.018307f
C420 VTAIL.n316 B 0.009837f
C421 VTAIL.n317 B 0.023252f
C422 VTAIL.n318 B 0.010416f
C423 VTAIL.n319 B 0.018307f
C424 VTAIL.n320 B 0.010127f
C425 VTAIL.n321 B 0.023252f
C426 VTAIL.n322 B 0.009837f
C427 VTAIL.n323 B 0.010416f
C428 VTAIL.n324 B 0.018307f
C429 VTAIL.n325 B 0.009837f
C430 VTAIL.n326 B 0.023252f
C431 VTAIL.n327 B 0.010416f
C432 VTAIL.n328 B 0.018307f
C433 VTAIL.n329 B 0.009837f
C434 VTAIL.n330 B 0.023252f
C435 VTAIL.n331 B 0.010416f
C436 VTAIL.n332 B 0.018307f
C437 VTAIL.n333 B 0.009837f
C438 VTAIL.n334 B 0.023252f
C439 VTAIL.n335 B 0.010416f
C440 VTAIL.n336 B 0.018307f
C441 VTAIL.n337 B 0.009837f
C442 VTAIL.n338 B 0.023252f
C443 VTAIL.n339 B 0.010416f
C444 VTAIL.n340 B 0.018307f
C445 VTAIL.n341 B 0.009837f
C446 VTAIL.n342 B 0.017439f
C447 VTAIL.n343 B 0.013736f
C448 VTAIL.t3 B 0.038545f
C449 VTAIL.n344 B 0.13441f
C450 VTAIL.n345 B 1.46542f
C451 VTAIL.n346 B 0.009837f
C452 VTAIL.n347 B 0.010416f
C453 VTAIL.n348 B 0.023252f
C454 VTAIL.n349 B 0.023252f
C455 VTAIL.n350 B 0.010416f
C456 VTAIL.n351 B 0.009837f
C457 VTAIL.n352 B 0.018307f
C458 VTAIL.n353 B 0.018307f
C459 VTAIL.n354 B 0.009837f
C460 VTAIL.n355 B 0.010416f
C461 VTAIL.n356 B 0.023252f
C462 VTAIL.n357 B 0.023252f
C463 VTAIL.n358 B 0.010416f
C464 VTAIL.n359 B 0.009837f
C465 VTAIL.n360 B 0.018307f
C466 VTAIL.n361 B 0.018307f
C467 VTAIL.n362 B 0.009837f
C468 VTAIL.n363 B 0.010416f
C469 VTAIL.n364 B 0.023252f
C470 VTAIL.n365 B 0.023252f
C471 VTAIL.n366 B 0.010416f
C472 VTAIL.n367 B 0.009837f
C473 VTAIL.n368 B 0.018307f
C474 VTAIL.n369 B 0.018307f
C475 VTAIL.n370 B 0.009837f
C476 VTAIL.n371 B 0.010416f
C477 VTAIL.n372 B 0.023252f
C478 VTAIL.n373 B 0.023252f
C479 VTAIL.n374 B 0.010416f
C480 VTAIL.n375 B 0.009837f
C481 VTAIL.n376 B 0.018307f
C482 VTAIL.n377 B 0.018307f
C483 VTAIL.n378 B 0.009837f
C484 VTAIL.n379 B 0.010416f
C485 VTAIL.n380 B 0.023252f
C486 VTAIL.n381 B 0.023252f
C487 VTAIL.n382 B 0.010416f
C488 VTAIL.n383 B 0.009837f
C489 VTAIL.n384 B 0.018307f
C490 VTAIL.n385 B 0.018307f
C491 VTAIL.n386 B 0.009837f
C492 VTAIL.n387 B 0.010416f
C493 VTAIL.n388 B 0.023252f
C494 VTAIL.n389 B 0.023252f
C495 VTAIL.n390 B 0.023252f
C496 VTAIL.n391 B 0.010127f
C497 VTAIL.n392 B 0.009837f
C498 VTAIL.n393 B 0.018307f
C499 VTAIL.n394 B 0.018307f
C500 VTAIL.n395 B 0.009837f
C501 VTAIL.n396 B 0.010416f
C502 VTAIL.n397 B 0.023252f
C503 VTAIL.n398 B 0.023252f
C504 VTAIL.n399 B 0.010416f
C505 VTAIL.n400 B 0.009837f
C506 VTAIL.n401 B 0.018307f
C507 VTAIL.n402 B 0.018307f
C508 VTAIL.n403 B 0.009837f
C509 VTAIL.n404 B 0.010416f
C510 VTAIL.n405 B 0.023252f
C511 VTAIL.n406 B 0.050991f
C512 VTAIL.n407 B 0.010416f
C513 VTAIL.n408 B 0.009837f
C514 VTAIL.n409 B 0.043066f
C515 VTAIL.n410 B 0.028622f
C516 VTAIL.n411 B 1.41959f
C517 VTAIL.t4 B 0.264305f
C518 VTAIL.t7 B 0.264305f
C519 VTAIL.n412 B 2.35394f
C520 VTAIL.n413 B 0.408445f
C521 VTAIL.n414 B 0.026102f
C522 VTAIL.n415 B 0.018307f
C523 VTAIL.n416 B 0.009837f
C524 VTAIL.n417 B 0.023252f
C525 VTAIL.n418 B 0.010416f
C526 VTAIL.n419 B 0.018307f
C527 VTAIL.n420 B 0.009837f
C528 VTAIL.n421 B 0.023252f
C529 VTAIL.n422 B 0.010416f
C530 VTAIL.n423 B 0.018307f
C531 VTAIL.n424 B 0.010127f
C532 VTAIL.n425 B 0.023252f
C533 VTAIL.n426 B 0.009837f
C534 VTAIL.n427 B 0.010416f
C535 VTAIL.n428 B 0.018307f
C536 VTAIL.n429 B 0.009837f
C537 VTAIL.n430 B 0.023252f
C538 VTAIL.n431 B 0.010416f
C539 VTAIL.n432 B 0.018307f
C540 VTAIL.n433 B 0.009837f
C541 VTAIL.n434 B 0.023252f
C542 VTAIL.n435 B 0.010416f
C543 VTAIL.n436 B 0.018307f
C544 VTAIL.n437 B 0.009837f
C545 VTAIL.n438 B 0.023252f
C546 VTAIL.n439 B 0.010416f
C547 VTAIL.n440 B 0.018307f
C548 VTAIL.n441 B 0.009837f
C549 VTAIL.n442 B 0.023252f
C550 VTAIL.n443 B 0.010416f
C551 VTAIL.n444 B 0.018307f
C552 VTAIL.n445 B 0.009837f
C553 VTAIL.n446 B 0.017439f
C554 VTAIL.n447 B 0.013736f
C555 VTAIL.t0 B 0.038545f
C556 VTAIL.n448 B 0.13441f
C557 VTAIL.n449 B 1.46542f
C558 VTAIL.n450 B 0.009837f
C559 VTAIL.n451 B 0.010416f
C560 VTAIL.n452 B 0.023252f
C561 VTAIL.n453 B 0.023252f
C562 VTAIL.n454 B 0.010416f
C563 VTAIL.n455 B 0.009837f
C564 VTAIL.n456 B 0.018307f
C565 VTAIL.n457 B 0.018307f
C566 VTAIL.n458 B 0.009837f
C567 VTAIL.n459 B 0.010416f
C568 VTAIL.n460 B 0.023252f
C569 VTAIL.n461 B 0.023252f
C570 VTAIL.n462 B 0.010416f
C571 VTAIL.n463 B 0.009837f
C572 VTAIL.n464 B 0.018307f
C573 VTAIL.n465 B 0.018307f
C574 VTAIL.n466 B 0.009837f
C575 VTAIL.n467 B 0.010416f
C576 VTAIL.n468 B 0.023252f
C577 VTAIL.n469 B 0.023252f
C578 VTAIL.n470 B 0.010416f
C579 VTAIL.n471 B 0.009837f
C580 VTAIL.n472 B 0.018307f
C581 VTAIL.n473 B 0.018307f
C582 VTAIL.n474 B 0.009837f
C583 VTAIL.n475 B 0.010416f
C584 VTAIL.n476 B 0.023252f
C585 VTAIL.n477 B 0.023252f
C586 VTAIL.n478 B 0.010416f
C587 VTAIL.n479 B 0.009837f
C588 VTAIL.n480 B 0.018307f
C589 VTAIL.n481 B 0.018307f
C590 VTAIL.n482 B 0.009837f
C591 VTAIL.n483 B 0.010416f
C592 VTAIL.n484 B 0.023252f
C593 VTAIL.n485 B 0.023252f
C594 VTAIL.n486 B 0.010416f
C595 VTAIL.n487 B 0.009837f
C596 VTAIL.n488 B 0.018307f
C597 VTAIL.n489 B 0.018307f
C598 VTAIL.n490 B 0.009837f
C599 VTAIL.n491 B 0.010416f
C600 VTAIL.n492 B 0.023252f
C601 VTAIL.n493 B 0.023252f
C602 VTAIL.n494 B 0.023252f
C603 VTAIL.n495 B 0.010127f
C604 VTAIL.n496 B 0.009837f
C605 VTAIL.n497 B 0.018307f
C606 VTAIL.n498 B 0.018307f
C607 VTAIL.n499 B 0.009837f
C608 VTAIL.n500 B 0.010416f
C609 VTAIL.n501 B 0.023252f
C610 VTAIL.n502 B 0.023252f
C611 VTAIL.n503 B 0.010416f
C612 VTAIL.n504 B 0.009837f
C613 VTAIL.n505 B 0.018307f
C614 VTAIL.n506 B 0.018307f
C615 VTAIL.n507 B 0.009837f
C616 VTAIL.n508 B 0.010416f
C617 VTAIL.n509 B 0.023252f
C618 VTAIL.n510 B 0.050991f
C619 VTAIL.n511 B 0.010416f
C620 VTAIL.n512 B 0.009837f
C621 VTAIL.n513 B 0.043066f
C622 VTAIL.n514 B 0.028622f
C623 VTAIL.n515 B 0.156666f
C624 VTAIL.n516 B 0.026102f
C625 VTAIL.n517 B 0.018307f
C626 VTAIL.n518 B 0.009837f
C627 VTAIL.n519 B 0.023252f
C628 VTAIL.n520 B 0.010416f
C629 VTAIL.n521 B 0.018307f
C630 VTAIL.n522 B 0.009837f
C631 VTAIL.n523 B 0.023252f
C632 VTAIL.n524 B 0.010416f
C633 VTAIL.n525 B 0.018307f
C634 VTAIL.n526 B 0.010127f
C635 VTAIL.n527 B 0.023252f
C636 VTAIL.n528 B 0.009837f
C637 VTAIL.n529 B 0.010416f
C638 VTAIL.n530 B 0.018307f
C639 VTAIL.n531 B 0.009837f
C640 VTAIL.n532 B 0.023252f
C641 VTAIL.n533 B 0.010416f
C642 VTAIL.n534 B 0.018307f
C643 VTAIL.n535 B 0.009837f
C644 VTAIL.n536 B 0.023252f
C645 VTAIL.n537 B 0.010416f
C646 VTAIL.n538 B 0.018307f
C647 VTAIL.n539 B 0.009837f
C648 VTAIL.n540 B 0.023252f
C649 VTAIL.n541 B 0.010416f
C650 VTAIL.n542 B 0.018307f
C651 VTAIL.n543 B 0.009837f
C652 VTAIL.n544 B 0.023252f
C653 VTAIL.n545 B 0.010416f
C654 VTAIL.n546 B 0.018307f
C655 VTAIL.n547 B 0.009837f
C656 VTAIL.n548 B 0.017439f
C657 VTAIL.n549 B 0.013736f
C658 VTAIL.t11 B 0.038545f
C659 VTAIL.n550 B 0.13441f
C660 VTAIL.n551 B 1.46542f
C661 VTAIL.n552 B 0.009837f
C662 VTAIL.n553 B 0.010416f
C663 VTAIL.n554 B 0.023252f
C664 VTAIL.n555 B 0.023252f
C665 VTAIL.n556 B 0.010416f
C666 VTAIL.n557 B 0.009837f
C667 VTAIL.n558 B 0.018307f
C668 VTAIL.n559 B 0.018307f
C669 VTAIL.n560 B 0.009837f
C670 VTAIL.n561 B 0.010416f
C671 VTAIL.n562 B 0.023252f
C672 VTAIL.n563 B 0.023252f
C673 VTAIL.n564 B 0.010416f
C674 VTAIL.n565 B 0.009837f
C675 VTAIL.n566 B 0.018307f
C676 VTAIL.n567 B 0.018307f
C677 VTAIL.n568 B 0.009837f
C678 VTAIL.n569 B 0.010416f
C679 VTAIL.n570 B 0.023252f
C680 VTAIL.n571 B 0.023252f
C681 VTAIL.n572 B 0.010416f
C682 VTAIL.n573 B 0.009837f
C683 VTAIL.n574 B 0.018307f
C684 VTAIL.n575 B 0.018307f
C685 VTAIL.n576 B 0.009837f
C686 VTAIL.n577 B 0.010416f
C687 VTAIL.n578 B 0.023252f
C688 VTAIL.n579 B 0.023252f
C689 VTAIL.n580 B 0.010416f
C690 VTAIL.n581 B 0.009837f
C691 VTAIL.n582 B 0.018307f
C692 VTAIL.n583 B 0.018307f
C693 VTAIL.n584 B 0.009837f
C694 VTAIL.n585 B 0.010416f
C695 VTAIL.n586 B 0.023252f
C696 VTAIL.n587 B 0.023252f
C697 VTAIL.n588 B 0.010416f
C698 VTAIL.n589 B 0.009837f
C699 VTAIL.n590 B 0.018307f
C700 VTAIL.n591 B 0.018307f
C701 VTAIL.n592 B 0.009837f
C702 VTAIL.n593 B 0.010416f
C703 VTAIL.n594 B 0.023252f
C704 VTAIL.n595 B 0.023252f
C705 VTAIL.n596 B 0.023252f
C706 VTAIL.n597 B 0.010127f
C707 VTAIL.n598 B 0.009837f
C708 VTAIL.n599 B 0.018307f
C709 VTAIL.n600 B 0.018307f
C710 VTAIL.n601 B 0.009837f
C711 VTAIL.n602 B 0.010416f
C712 VTAIL.n603 B 0.023252f
C713 VTAIL.n604 B 0.023252f
C714 VTAIL.n605 B 0.010416f
C715 VTAIL.n606 B 0.009837f
C716 VTAIL.n607 B 0.018307f
C717 VTAIL.n608 B 0.018307f
C718 VTAIL.n609 B 0.009837f
C719 VTAIL.n610 B 0.010416f
C720 VTAIL.n611 B 0.023252f
C721 VTAIL.n612 B 0.050991f
C722 VTAIL.n613 B 0.010416f
C723 VTAIL.n614 B 0.009837f
C724 VTAIL.n615 B 0.043066f
C725 VTAIL.n616 B 0.028622f
C726 VTAIL.n617 B 0.156666f
C727 VTAIL.t15 B 0.264305f
C728 VTAIL.t8 B 0.264305f
C729 VTAIL.n618 B 2.35394f
C730 VTAIL.n619 B 0.408445f
C731 VTAIL.n620 B 0.026102f
C732 VTAIL.n621 B 0.018307f
C733 VTAIL.n622 B 0.009837f
C734 VTAIL.n623 B 0.023252f
C735 VTAIL.n624 B 0.010416f
C736 VTAIL.n625 B 0.018307f
C737 VTAIL.n626 B 0.009837f
C738 VTAIL.n627 B 0.023252f
C739 VTAIL.n628 B 0.010416f
C740 VTAIL.n629 B 0.018307f
C741 VTAIL.n630 B 0.010127f
C742 VTAIL.n631 B 0.023252f
C743 VTAIL.n632 B 0.009837f
C744 VTAIL.n633 B 0.010416f
C745 VTAIL.n634 B 0.018307f
C746 VTAIL.n635 B 0.009837f
C747 VTAIL.n636 B 0.023252f
C748 VTAIL.n637 B 0.010416f
C749 VTAIL.n638 B 0.018307f
C750 VTAIL.n639 B 0.009837f
C751 VTAIL.n640 B 0.023252f
C752 VTAIL.n641 B 0.010416f
C753 VTAIL.n642 B 0.018307f
C754 VTAIL.n643 B 0.009837f
C755 VTAIL.n644 B 0.023252f
C756 VTAIL.n645 B 0.010416f
C757 VTAIL.n646 B 0.018307f
C758 VTAIL.n647 B 0.009837f
C759 VTAIL.n648 B 0.023252f
C760 VTAIL.n649 B 0.010416f
C761 VTAIL.n650 B 0.018307f
C762 VTAIL.n651 B 0.009837f
C763 VTAIL.n652 B 0.017439f
C764 VTAIL.n653 B 0.013736f
C765 VTAIL.t12 B 0.038545f
C766 VTAIL.n654 B 0.13441f
C767 VTAIL.n655 B 1.46542f
C768 VTAIL.n656 B 0.009837f
C769 VTAIL.n657 B 0.010416f
C770 VTAIL.n658 B 0.023252f
C771 VTAIL.n659 B 0.023252f
C772 VTAIL.n660 B 0.010416f
C773 VTAIL.n661 B 0.009837f
C774 VTAIL.n662 B 0.018307f
C775 VTAIL.n663 B 0.018307f
C776 VTAIL.n664 B 0.009837f
C777 VTAIL.n665 B 0.010416f
C778 VTAIL.n666 B 0.023252f
C779 VTAIL.n667 B 0.023252f
C780 VTAIL.n668 B 0.010416f
C781 VTAIL.n669 B 0.009837f
C782 VTAIL.n670 B 0.018307f
C783 VTAIL.n671 B 0.018307f
C784 VTAIL.n672 B 0.009837f
C785 VTAIL.n673 B 0.010416f
C786 VTAIL.n674 B 0.023252f
C787 VTAIL.n675 B 0.023252f
C788 VTAIL.n676 B 0.010416f
C789 VTAIL.n677 B 0.009837f
C790 VTAIL.n678 B 0.018307f
C791 VTAIL.n679 B 0.018307f
C792 VTAIL.n680 B 0.009837f
C793 VTAIL.n681 B 0.010416f
C794 VTAIL.n682 B 0.023252f
C795 VTAIL.n683 B 0.023252f
C796 VTAIL.n684 B 0.010416f
C797 VTAIL.n685 B 0.009837f
C798 VTAIL.n686 B 0.018307f
C799 VTAIL.n687 B 0.018307f
C800 VTAIL.n688 B 0.009837f
C801 VTAIL.n689 B 0.010416f
C802 VTAIL.n690 B 0.023252f
C803 VTAIL.n691 B 0.023252f
C804 VTAIL.n692 B 0.010416f
C805 VTAIL.n693 B 0.009837f
C806 VTAIL.n694 B 0.018307f
C807 VTAIL.n695 B 0.018307f
C808 VTAIL.n696 B 0.009837f
C809 VTAIL.n697 B 0.010416f
C810 VTAIL.n698 B 0.023252f
C811 VTAIL.n699 B 0.023252f
C812 VTAIL.n700 B 0.023252f
C813 VTAIL.n701 B 0.010127f
C814 VTAIL.n702 B 0.009837f
C815 VTAIL.n703 B 0.018307f
C816 VTAIL.n704 B 0.018307f
C817 VTAIL.n705 B 0.009837f
C818 VTAIL.n706 B 0.010416f
C819 VTAIL.n707 B 0.023252f
C820 VTAIL.n708 B 0.023252f
C821 VTAIL.n709 B 0.010416f
C822 VTAIL.n710 B 0.009837f
C823 VTAIL.n711 B 0.018307f
C824 VTAIL.n712 B 0.018307f
C825 VTAIL.n713 B 0.009837f
C826 VTAIL.n714 B 0.010416f
C827 VTAIL.n715 B 0.023252f
C828 VTAIL.n716 B 0.050991f
C829 VTAIL.n717 B 0.010416f
C830 VTAIL.n718 B 0.009837f
C831 VTAIL.n719 B 0.043066f
C832 VTAIL.n720 B 0.028622f
C833 VTAIL.n721 B 1.41959f
C834 VTAIL.n722 B 0.026102f
C835 VTAIL.n723 B 0.018307f
C836 VTAIL.n724 B 0.009837f
C837 VTAIL.n725 B 0.023252f
C838 VTAIL.n726 B 0.010416f
C839 VTAIL.n727 B 0.018307f
C840 VTAIL.n728 B 0.009837f
C841 VTAIL.n729 B 0.023252f
C842 VTAIL.n730 B 0.010416f
C843 VTAIL.n731 B 0.018307f
C844 VTAIL.n732 B 0.010127f
C845 VTAIL.n733 B 0.023252f
C846 VTAIL.n734 B 0.010416f
C847 VTAIL.n735 B 0.018307f
C848 VTAIL.n736 B 0.009837f
C849 VTAIL.n737 B 0.023252f
C850 VTAIL.n738 B 0.010416f
C851 VTAIL.n739 B 0.018307f
C852 VTAIL.n740 B 0.009837f
C853 VTAIL.n741 B 0.023252f
C854 VTAIL.n742 B 0.010416f
C855 VTAIL.n743 B 0.018307f
C856 VTAIL.n744 B 0.009837f
C857 VTAIL.n745 B 0.023252f
C858 VTAIL.n746 B 0.010416f
C859 VTAIL.n747 B 0.018307f
C860 VTAIL.n748 B 0.009837f
C861 VTAIL.n749 B 0.023252f
C862 VTAIL.n750 B 0.010416f
C863 VTAIL.n751 B 0.018307f
C864 VTAIL.n752 B 0.009837f
C865 VTAIL.n753 B 0.017439f
C866 VTAIL.n754 B 0.013736f
C867 VTAIL.t6 B 0.038545f
C868 VTAIL.n755 B 0.13441f
C869 VTAIL.n756 B 1.46542f
C870 VTAIL.n757 B 0.009837f
C871 VTAIL.n758 B 0.010416f
C872 VTAIL.n759 B 0.023252f
C873 VTAIL.n760 B 0.023252f
C874 VTAIL.n761 B 0.010416f
C875 VTAIL.n762 B 0.009837f
C876 VTAIL.n763 B 0.018307f
C877 VTAIL.n764 B 0.018307f
C878 VTAIL.n765 B 0.009837f
C879 VTAIL.n766 B 0.010416f
C880 VTAIL.n767 B 0.023252f
C881 VTAIL.n768 B 0.023252f
C882 VTAIL.n769 B 0.010416f
C883 VTAIL.n770 B 0.009837f
C884 VTAIL.n771 B 0.018307f
C885 VTAIL.n772 B 0.018307f
C886 VTAIL.n773 B 0.009837f
C887 VTAIL.n774 B 0.010416f
C888 VTAIL.n775 B 0.023252f
C889 VTAIL.n776 B 0.023252f
C890 VTAIL.n777 B 0.010416f
C891 VTAIL.n778 B 0.009837f
C892 VTAIL.n779 B 0.018307f
C893 VTAIL.n780 B 0.018307f
C894 VTAIL.n781 B 0.009837f
C895 VTAIL.n782 B 0.010416f
C896 VTAIL.n783 B 0.023252f
C897 VTAIL.n784 B 0.023252f
C898 VTAIL.n785 B 0.010416f
C899 VTAIL.n786 B 0.009837f
C900 VTAIL.n787 B 0.018307f
C901 VTAIL.n788 B 0.018307f
C902 VTAIL.n789 B 0.009837f
C903 VTAIL.n790 B 0.010416f
C904 VTAIL.n791 B 0.023252f
C905 VTAIL.n792 B 0.023252f
C906 VTAIL.n793 B 0.010416f
C907 VTAIL.n794 B 0.009837f
C908 VTAIL.n795 B 0.018307f
C909 VTAIL.n796 B 0.018307f
C910 VTAIL.n797 B 0.009837f
C911 VTAIL.n798 B 0.009837f
C912 VTAIL.n799 B 0.010416f
C913 VTAIL.n800 B 0.023252f
C914 VTAIL.n801 B 0.023252f
C915 VTAIL.n802 B 0.023252f
C916 VTAIL.n803 B 0.010127f
C917 VTAIL.n804 B 0.009837f
C918 VTAIL.n805 B 0.018307f
C919 VTAIL.n806 B 0.018307f
C920 VTAIL.n807 B 0.009837f
C921 VTAIL.n808 B 0.010416f
C922 VTAIL.n809 B 0.023252f
C923 VTAIL.n810 B 0.023252f
C924 VTAIL.n811 B 0.010416f
C925 VTAIL.n812 B 0.009837f
C926 VTAIL.n813 B 0.018307f
C927 VTAIL.n814 B 0.018307f
C928 VTAIL.n815 B 0.009837f
C929 VTAIL.n816 B 0.010416f
C930 VTAIL.n817 B 0.023252f
C931 VTAIL.n818 B 0.050991f
C932 VTAIL.n819 B 0.010416f
C933 VTAIL.n820 B 0.009837f
C934 VTAIL.n821 B 0.043066f
C935 VTAIL.n822 B 0.028622f
C936 VTAIL.n823 B 1.41616f
C937 VP.n0 B 0.026462f
C938 VP.t1 B 2.51403f
C939 VP.n1 B 0.0217f
C940 VP.n2 B 0.026462f
C941 VP.t4 B 2.51403f
C942 VP.n3 B 0.03863f
C943 VP.n4 B 0.026462f
C944 VP.t7 B 2.51403f
C945 VP.n5 B 0.051654f
C946 VP.n6 B 0.026462f
C947 VP.t2 B 2.51403f
C948 VP.n7 B 0.941978f
C949 VP.n8 B 0.026462f
C950 VP.t0 B 2.51403f
C951 VP.n9 B 0.0217f
C952 VP.n10 B 0.026462f
C953 VP.t5 B 2.51403f
C954 VP.n11 B 0.03863f
C955 VP.n12 B 0.196894f
C956 VP.t6 B 2.51403f
C957 VP.t3 B 2.64353f
C958 VP.n13 B 0.939239f
C959 VP.n14 B 0.943875f
C960 VP.n15 B 0.042501f
C961 VP.n16 B 0.03863f
C962 VP.n17 B 0.026462f
C963 VP.n18 B 0.026462f
C964 VP.n19 B 0.026462f
C965 VP.n20 B 0.042501f
C966 VP.n21 B 0.877932f
C967 VP.n22 B 0.031788f
C968 VP.n23 B 0.051654f
C969 VP.n24 B 0.026462f
C970 VP.n25 B 0.026462f
C971 VP.n26 B 0.026462f
C972 VP.n27 B 0.053225f
C973 VP.n28 B 0.028866f
C974 VP.n29 B 0.941978f
C975 VP.n30 B 1.54417f
C976 VP.n31 B 1.56237f
C977 VP.n32 B 0.026462f
C978 VP.n33 B 0.028866f
C979 VP.n34 B 0.053225f
C980 VP.n35 B 0.0217f
C981 VP.n36 B 0.026462f
C982 VP.n37 B 0.026462f
C983 VP.n38 B 0.026462f
C984 VP.n39 B 0.031788f
C985 VP.n40 B 0.877932f
C986 VP.n41 B 0.042501f
C987 VP.n42 B 0.03863f
C988 VP.n43 B 0.026462f
C989 VP.n44 B 0.026462f
C990 VP.n45 B 0.026462f
C991 VP.n46 B 0.042501f
C992 VP.n47 B 0.877932f
C993 VP.n48 B 0.031788f
C994 VP.n49 B 0.051654f
C995 VP.n50 B 0.026462f
C996 VP.n51 B 0.026462f
C997 VP.n52 B 0.026462f
C998 VP.n53 B 0.053225f
C999 VP.n54 B 0.028866f
C1000 VP.n55 B 0.941978f
C1001 VP.n56 B 0.028668f
.ends

