* NGSPICE file created from diff_pair_sample_1404.ext - technology: sky130A

.subckt diff_pair_sample_1404 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=4.5942 pd=24.34 as=1.9437 ps=12.11 w=11.78 l=2.1
X1 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=4.5942 pd=24.34 as=0 ps=0 w=11.78 l=2.1
X2 VDD2.t4 VN.t1 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9437 pd=12.11 as=4.5942 ps=24.34 w=11.78 l=2.1
X3 VTAIL.t7 VN.t2 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9437 pd=12.11 as=1.9437 ps=12.11 w=11.78 l=2.1
X4 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=4.5942 pd=24.34 as=0 ps=0 w=11.78 l=2.1
X5 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=4.5942 pd=24.34 as=0 ps=0 w=11.78 l=2.1
X6 VDD2.t2 VN.t3 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.9437 pd=12.11 as=4.5942 ps=24.34 w=11.78 l=2.1
X7 VTAIL.t10 VN.t4 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=1.9437 pd=12.11 as=1.9437 ps=12.11 w=11.78 l=2.1
X8 VDD1.t5 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.9437 pd=12.11 as=4.5942 ps=24.34 w=11.78 l=2.1
X9 VDD1.t4 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.5942 pd=24.34 as=1.9437 ps=12.11 w=11.78 l=2.1
X10 VDD1.t3 VP.t2 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=4.5942 pd=24.34 as=1.9437 ps=12.11 w=11.78 l=2.1
X11 VTAIL.t3 VP.t3 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9437 pd=12.11 as=1.9437 ps=12.11 w=11.78 l=2.1
X12 VDD1.t1 VP.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9437 pd=12.11 as=4.5942 ps=24.34 w=11.78 l=2.1
X13 VDD2.t0 VN.t5 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=4.5942 pd=24.34 as=1.9437 ps=12.11 w=11.78 l=2.1
X14 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.5942 pd=24.34 as=0 ps=0 w=11.78 l=2.1
X15 VTAIL.t5 VP.t5 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=1.9437 pd=12.11 as=1.9437 ps=12.11 w=11.78 l=2.1
R0 VN.n2 VN.t0 169.589
R1 VN.n14 VN.t3 169.589
R2 VN.n21 VN.n12 161.3
R3 VN.n20 VN.n19 161.3
R4 VN.n18 VN.n13 161.3
R5 VN.n17 VN.n16 161.3
R6 VN.n9 VN.n0 161.3
R7 VN.n8 VN.n7 161.3
R8 VN.n6 VN.n1 161.3
R9 VN.n5 VN.n4 161.3
R10 VN.n3 VN.t2 135.19
R11 VN.n10 VN.t1 135.19
R12 VN.n15 VN.t4 135.19
R13 VN.n22 VN.t5 135.19
R14 VN.n11 VN.n10 89.7593
R15 VN.n23 VN.n22 89.7593
R16 VN.n8 VN.n1 56.5617
R17 VN.n20 VN.n13 56.5617
R18 VN VN.n23 46.8959
R19 VN.n15 VN.n14 46.2728
R20 VN.n3 VN.n2 46.2728
R21 VN.n4 VN.n3 24.5923
R22 VN.n4 VN.n1 24.5923
R23 VN.n9 VN.n8 24.5923
R24 VN.n16 VN.n13 24.5923
R25 VN.n16 VN.n15 24.5923
R26 VN.n21 VN.n20 24.5923
R27 VN.n10 VN.n9 21.1495
R28 VN.n22 VN.n21 21.1495
R29 VN.n17 VN.n14 8.85089
R30 VN.n5 VN.n2 8.85089
R31 VN.n23 VN.n12 0.278335
R32 VN.n11 VN.n0 0.278335
R33 VN.n19 VN.n12 0.189894
R34 VN.n19 VN.n18 0.189894
R35 VN.n18 VN.n17 0.189894
R36 VN.n6 VN.n5 0.189894
R37 VN.n7 VN.n6 0.189894
R38 VN.n7 VN.n0 0.189894
R39 VN VN.n11 0.153485
R40 VTAIL.n7 VTAIL.t6 47.3699
R41 VTAIL.n11 VTAIL.t8 47.3697
R42 VTAIL.n2 VTAIL.t2 47.3697
R43 VTAIL.n10 VTAIL.t0 47.3697
R44 VTAIL.n9 VTAIL.n8 45.6891
R45 VTAIL.n6 VTAIL.n5 45.6891
R46 VTAIL.n1 VTAIL.n0 45.6889
R47 VTAIL.n4 VTAIL.n3 45.6889
R48 VTAIL.n6 VTAIL.n4 26.7117
R49 VTAIL.n11 VTAIL.n10 24.6169
R50 VTAIL.n7 VTAIL.n6 2.09533
R51 VTAIL.n10 VTAIL.n9 2.09533
R52 VTAIL.n4 VTAIL.n2 2.09533
R53 VTAIL.n0 VTAIL.t11 1.68131
R54 VTAIL.n0 VTAIL.t7 1.68131
R55 VTAIL.n3 VTAIL.t1 1.68131
R56 VTAIL.n3 VTAIL.t5 1.68131
R57 VTAIL.n8 VTAIL.t4 1.68131
R58 VTAIL.n8 VTAIL.t3 1.68131
R59 VTAIL.n5 VTAIL.t9 1.68131
R60 VTAIL.n5 VTAIL.t10 1.68131
R61 VTAIL.n9 VTAIL.n7 1.51774
R62 VTAIL.n2 VTAIL.n1 1.51774
R63 VTAIL VTAIL.n11 1.51343
R64 VTAIL VTAIL.n1 0.582397
R65 VDD2.n1 VDD2.t5 65.5643
R66 VDD2.n2 VDD2.t0 64.0487
R67 VDD2.n1 VDD2.n0 62.836
R68 VDD2 VDD2.n3 62.8332
R69 VDD2.n2 VDD2.n1 40.6787
R70 VDD2.n3 VDD2.t1 1.68131
R71 VDD2.n3 VDD2.t2 1.68131
R72 VDD2.n0 VDD2.t3 1.68131
R73 VDD2.n0 VDD2.t4 1.68131
R74 VDD2 VDD2.n2 1.62981
R75 B.n763 B.n762 585
R76 B.n300 B.n115 585
R77 B.n299 B.n298 585
R78 B.n297 B.n296 585
R79 B.n295 B.n294 585
R80 B.n293 B.n292 585
R81 B.n291 B.n290 585
R82 B.n289 B.n288 585
R83 B.n287 B.n286 585
R84 B.n285 B.n284 585
R85 B.n283 B.n282 585
R86 B.n281 B.n280 585
R87 B.n279 B.n278 585
R88 B.n277 B.n276 585
R89 B.n275 B.n274 585
R90 B.n273 B.n272 585
R91 B.n271 B.n270 585
R92 B.n269 B.n268 585
R93 B.n267 B.n266 585
R94 B.n265 B.n264 585
R95 B.n263 B.n262 585
R96 B.n261 B.n260 585
R97 B.n259 B.n258 585
R98 B.n257 B.n256 585
R99 B.n255 B.n254 585
R100 B.n253 B.n252 585
R101 B.n251 B.n250 585
R102 B.n249 B.n248 585
R103 B.n247 B.n246 585
R104 B.n245 B.n244 585
R105 B.n243 B.n242 585
R106 B.n241 B.n240 585
R107 B.n239 B.n238 585
R108 B.n237 B.n236 585
R109 B.n235 B.n234 585
R110 B.n233 B.n232 585
R111 B.n231 B.n230 585
R112 B.n229 B.n228 585
R113 B.n227 B.n226 585
R114 B.n225 B.n224 585
R115 B.n223 B.n222 585
R116 B.n220 B.n219 585
R117 B.n218 B.n217 585
R118 B.n216 B.n215 585
R119 B.n214 B.n213 585
R120 B.n212 B.n211 585
R121 B.n210 B.n209 585
R122 B.n208 B.n207 585
R123 B.n206 B.n205 585
R124 B.n204 B.n203 585
R125 B.n202 B.n201 585
R126 B.n199 B.n198 585
R127 B.n197 B.n196 585
R128 B.n195 B.n194 585
R129 B.n193 B.n192 585
R130 B.n191 B.n190 585
R131 B.n189 B.n188 585
R132 B.n187 B.n186 585
R133 B.n185 B.n184 585
R134 B.n183 B.n182 585
R135 B.n181 B.n180 585
R136 B.n179 B.n178 585
R137 B.n177 B.n176 585
R138 B.n175 B.n174 585
R139 B.n173 B.n172 585
R140 B.n171 B.n170 585
R141 B.n169 B.n168 585
R142 B.n167 B.n166 585
R143 B.n165 B.n164 585
R144 B.n163 B.n162 585
R145 B.n161 B.n160 585
R146 B.n159 B.n158 585
R147 B.n157 B.n156 585
R148 B.n155 B.n154 585
R149 B.n153 B.n152 585
R150 B.n151 B.n150 585
R151 B.n149 B.n148 585
R152 B.n147 B.n146 585
R153 B.n145 B.n144 585
R154 B.n143 B.n142 585
R155 B.n141 B.n140 585
R156 B.n139 B.n138 585
R157 B.n137 B.n136 585
R158 B.n135 B.n134 585
R159 B.n133 B.n132 585
R160 B.n131 B.n130 585
R161 B.n129 B.n128 585
R162 B.n127 B.n126 585
R163 B.n125 B.n124 585
R164 B.n123 B.n122 585
R165 B.n121 B.n120 585
R166 B.n68 B.n67 585
R167 B.n761 B.n69 585
R168 B.n766 B.n69 585
R169 B.n760 B.n759 585
R170 B.n759 B.n65 585
R171 B.n758 B.n64 585
R172 B.n772 B.n64 585
R173 B.n757 B.n63 585
R174 B.n773 B.n63 585
R175 B.n756 B.n62 585
R176 B.n774 B.n62 585
R177 B.n755 B.n754 585
R178 B.n754 B.n58 585
R179 B.n753 B.n57 585
R180 B.n780 B.n57 585
R181 B.n752 B.n56 585
R182 B.n781 B.n56 585
R183 B.n751 B.n55 585
R184 B.n782 B.n55 585
R185 B.n750 B.n749 585
R186 B.n749 B.n51 585
R187 B.n748 B.n50 585
R188 B.n788 B.n50 585
R189 B.n747 B.n49 585
R190 B.n789 B.n49 585
R191 B.n746 B.n48 585
R192 B.n790 B.n48 585
R193 B.n745 B.n744 585
R194 B.n744 B.n44 585
R195 B.n743 B.n43 585
R196 B.n796 B.n43 585
R197 B.n742 B.n42 585
R198 B.n797 B.n42 585
R199 B.n741 B.n41 585
R200 B.n798 B.n41 585
R201 B.n740 B.n739 585
R202 B.n739 B.n40 585
R203 B.n738 B.n36 585
R204 B.n804 B.n36 585
R205 B.n737 B.n35 585
R206 B.n805 B.n35 585
R207 B.n736 B.n34 585
R208 B.n806 B.n34 585
R209 B.n735 B.n734 585
R210 B.n734 B.n30 585
R211 B.n733 B.n29 585
R212 B.n812 B.n29 585
R213 B.n732 B.n28 585
R214 B.n813 B.n28 585
R215 B.n731 B.n27 585
R216 B.n814 B.n27 585
R217 B.n730 B.n729 585
R218 B.n729 B.n23 585
R219 B.n728 B.n22 585
R220 B.n820 B.n22 585
R221 B.n727 B.n21 585
R222 B.n821 B.n21 585
R223 B.n726 B.n20 585
R224 B.n822 B.n20 585
R225 B.n725 B.n724 585
R226 B.n724 B.n16 585
R227 B.n723 B.n15 585
R228 B.n828 B.n15 585
R229 B.n722 B.n14 585
R230 B.n829 B.n14 585
R231 B.n721 B.n13 585
R232 B.n830 B.n13 585
R233 B.n720 B.n719 585
R234 B.n719 B.n12 585
R235 B.n718 B.n717 585
R236 B.n718 B.n8 585
R237 B.n716 B.n7 585
R238 B.n837 B.n7 585
R239 B.n715 B.n6 585
R240 B.n838 B.n6 585
R241 B.n714 B.n5 585
R242 B.n839 B.n5 585
R243 B.n713 B.n712 585
R244 B.n712 B.n4 585
R245 B.n711 B.n301 585
R246 B.n711 B.n710 585
R247 B.n701 B.n302 585
R248 B.n303 B.n302 585
R249 B.n703 B.n702 585
R250 B.n704 B.n703 585
R251 B.n700 B.n307 585
R252 B.n311 B.n307 585
R253 B.n699 B.n698 585
R254 B.n698 B.n697 585
R255 B.n309 B.n308 585
R256 B.n310 B.n309 585
R257 B.n690 B.n689 585
R258 B.n691 B.n690 585
R259 B.n688 B.n316 585
R260 B.n316 B.n315 585
R261 B.n687 B.n686 585
R262 B.n686 B.n685 585
R263 B.n318 B.n317 585
R264 B.n319 B.n318 585
R265 B.n678 B.n677 585
R266 B.n679 B.n678 585
R267 B.n676 B.n324 585
R268 B.n324 B.n323 585
R269 B.n675 B.n674 585
R270 B.n674 B.n673 585
R271 B.n326 B.n325 585
R272 B.n327 B.n326 585
R273 B.n666 B.n665 585
R274 B.n667 B.n666 585
R275 B.n664 B.n332 585
R276 B.n332 B.n331 585
R277 B.n663 B.n662 585
R278 B.n662 B.n661 585
R279 B.n334 B.n333 585
R280 B.n654 B.n334 585
R281 B.n653 B.n652 585
R282 B.n655 B.n653 585
R283 B.n651 B.n339 585
R284 B.n339 B.n338 585
R285 B.n650 B.n649 585
R286 B.n649 B.n648 585
R287 B.n341 B.n340 585
R288 B.n342 B.n341 585
R289 B.n641 B.n640 585
R290 B.n642 B.n641 585
R291 B.n639 B.n347 585
R292 B.n347 B.n346 585
R293 B.n638 B.n637 585
R294 B.n637 B.n636 585
R295 B.n349 B.n348 585
R296 B.n350 B.n349 585
R297 B.n629 B.n628 585
R298 B.n630 B.n629 585
R299 B.n627 B.n355 585
R300 B.n355 B.n354 585
R301 B.n626 B.n625 585
R302 B.n625 B.n624 585
R303 B.n357 B.n356 585
R304 B.n358 B.n357 585
R305 B.n617 B.n616 585
R306 B.n618 B.n617 585
R307 B.n615 B.n363 585
R308 B.n363 B.n362 585
R309 B.n614 B.n613 585
R310 B.n613 B.n612 585
R311 B.n365 B.n364 585
R312 B.n366 B.n365 585
R313 B.n605 B.n604 585
R314 B.n606 B.n605 585
R315 B.n369 B.n368 585
R316 B.n424 B.n423 585
R317 B.n425 B.n421 585
R318 B.n421 B.n370 585
R319 B.n427 B.n426 585
R320 B.n429 B.n420 585
R321 B.n432 B.n431 585
R322 B.n433 B.n419 585
R323 B.n435 B.n434 585
R324 B.n437 B.n418 585
R325 B.n440 B.n439 585
R326 B.n441 B.n417 585
R327 B.n443 B.n442 585
R328 B.n445 B.n416 585
R329 B.n448 B.n447 585
R330 B.n449 B.n415 585
R331 B.n451 B.n450 585
R332 B.n453 B.n414 585
R333 B.n456 B.n455 585
R334 B.n457 B.n413 585
R335 B.n459 B.n458 585
R336 B.n461 B.n412 585
R337 B.n464 B.n463 585
R338 B.n465 B.n411 585
R339 B.n467 B.n466 585
R340 B.n469 B.n410 585
R341 B.n472 B.n471 585
R342 B.n473 B.n409 585
R343 B.n475 B.n474 585
R344 B.n477 B.n408 585
R345 B.n480 B.n479 585
R346 B.n481 B.n407 585
R347 B.n483 B.n482 585
R348 B.n485 B.n406 585
R349 B.n488 B.n487 585
R350 B.n489 B.n405 585
R351 B.n491 B.n490 585
R352 B.n493 B.n404 585
R353 B.n496 B.n495 585
R354 B.n497 B.n403 585
R355 B.n499 B.n498 585
R356 B.n501 B.n402 585
R357 B.n504 B.n503 585
R358 B.n505 B.n398 585
R359 B.n507 B.n506 585
R360 B.n509 B.n397 585
R361 B.n512 B.n511 585
R362 B.n513 B.n396 585
R363 B.n515 B.n514 585
R364 B.n517 B.n395 585
R365 B.n520 B.n519 585
R366 B.n521 B.n392 585
R367 B.n524 B.n523 585
R368 B.n526 B.n391 585
R369 B.n529 B.n528 585
R370 B.n530 B.n390 585
R371 B.n532 B.n531 585
R372 B.n534 B.n389 585
R373 B.n537 B.n536 585
R374 B.n538 B.n388 585
R375 B.n540 B.n539 585
R376 B.n542 B.n387 585
R377 B.n545 B.n544 585
R378 B.n546 B.n386 585
R379 B.n548 B.n547 585
R380 B.n550 B.n385 585
R381 B.n553 B.n552 585
R382 B.n554 B.n384 585
R383 B.n556 B.n555 585
R384 B.n558 B.n383 585
R385 B.n561 B.n560 585
R386 B.n562 B.n382 585
R387 B.n564 B.n563 585
R388 B.n566 B.n381 585
R389 B.n569 B.n568 585
R390 B.n570 B.n380 585
R391 B.n572 B.n571 585
R392 B.n574 B.n379 585
R393 B.n577 B.n576 585
R394 B.n578 B.n378 585
R395 B.n580 B.n579 585
R396 B.n582 B.n377 585
R397 B.n585 B.n584 585
R398 B.n586 B.n376 585
R399 B.n588 B.n587 585
R400 B.n590 B.n375 585
R401 B.n593 B.n592 585
R402 B.n594 B.n374 585
R403 B.n596 B.n595 585
R404 B.n598 B.n373 585
R405 B.n599 B.n372 585
R406 B.n602 B.n601 585
R407 B.n603 B.n371 585
R408 B.n371 B.n370 585
R409 B.n608 B.n607 585
R410 B.n607 B.n606 585
R411 B.n609 B.n367 585
R412 B.n367 B.n366 585
R413 B.n611 B.n610 585
R414 B.n612 B.n611 585
R415 B.n361 B.n360 585
R416 B.n362 B.n361 585
R417 B.n620 B.n619 585
R418 B.n619 B.n618 585
R419 B.n621 B.n359 585
R420 B.n359 B.n358 585
R421 B.n623 B.n622 585
R422 B.n624 B.n623 585
R423 B.n353 B.n352 585
R424 B.n354 B.n353 585
R425 B.n632 B.n631 585
R426 B.n631 B.n630 585
R427 B.n633 B.n351 585
R428 B.n351 B.n350 585
R429 B.n635 B.n634 585
R430 B.n636 B.n635 585
R431 B.n345 B.n344 585
R432 B.n346 B.n345 585
R433 B.n644 B.n643 585
R434 B.n643 B.n642 585
R435 B.n645 B.n343 585
R436 B.n343 B.n342 585
R437 B.n647 B.n646 585
R438 B.n648 B.n647 585
R439 B.n337 B.n336 585
R440 B.n338 B.n337 585
R441 B.n657 B.n656 585
R442 B.n656 B.n655 585
R443 B.n658 B.n335 585
R444 B.n654 B.n335 585
R445 B.n660 B.n659 585
R446 B.n661 B.n660 585
R447 B.n330 B.n329 585
R448 B.n331 B.n330 585
R449 B.n669 B.n668 585
R450 B.n668 B.n667 585
R451 B.n670 B.n328 585
R452 B.n328 B.n327 585
R453 B.n672 B.n671 585
R454 B.n673 B.n672 585
R455 B.n322 B.n321 585
R456 B.n323 B.n322 585
R457 B.n681 B.n680 585
R458 B.n680 B.n679 585
R459 B.n682 B.n320 585
R460 B.n320 B.n319 585
R461 B.n684 B.n683 585
R462 B.n685 B.n684 585
R463 B.n314 B.n313 585
R464 B.n315 B.n314 585
R465 B.n693 B.n692 585
R466 B.n692 B.n691 585
R467 B.n694 B.n312 585
R468 B.n312 B.n310 585
R469 B.n696 B.n695 585
R470 B.n697 B.n696 585
R471 B.n306 B.n305 585
R472 B.n311 B.n306 585
R473 B.n706 B.n705 585
R474 B.n705 B.n704 585
R475 B.n707 B.n304 585
R476 B.n304 B.n303 585
R477 B.n709 B.n708 585
R478 B.n710 B.n709 585
R479 B.n3 B.n0 585
R480 B.n4 B.n3 585
R481 B.n836 B.n1 585
R482 B.n837 B.n836 585
R483 B.n835 B.n834 585
R484 B.n835 B.n8 585
R485 B.n833 B.n9 585
R486 B.n12 B.n9 585
R487 B.n832 B.n831 585
R488 B.n831 B.n830 585
R489 B.n11 B.n10 585
R490 B.n829 B.n11 585
R491 B.n827 B.n826 585
R492 B.n828 B.n827 585
R493 B.n825 B.n17 585
R494 B.n17 B.n16 585
R495 B.n824 B.n823 585
R496 B.n823 B.n822 585
R497 B.n19 B.n18 585
R498 B.n821 B.n19 585
R499 B.n819 B.n818 585
R500 B.n820 B.n819 585
R501 B.n817 B.n24 585
R502 B.n24 B.n23 585
R503 B.n816 B.n815 585
R504 B.n815 B.n814 585
R505 B.n26 B.n25 585
R506 B.n813 B.n26 585
R507 B.n811 B.n810 585
R508 B.n812 B.n811 585
R509 B.n809 B.n31 585
R510 B.n31 B.n30 585
R511 B.n808 B.n807 585
R512 B.n807 B.n806 585
R513 B.n33 B.n32 585
R514 B.n805 B.n33 585
R515 B.n803 B.n802 585
R516 B.n804 B.n803 585
R517 B.n801 B.n37 585
R518 B.n40 B.n37 585
R519 B.n800 B.n799 585
R520 B.n799 B.n798 585
R521 B.n39 B.n38 585
R522 B.n797 B.n39 585
R523 B.n795 B.n794 585
R524 B.n796 B.n795 585
R525 B.n793 B.n45 585
R526 B.n45 B.n44 585
R527 B.n792 B.n791 585
R528 B.n791 B.n790 585
R529 B.n47 B.n46 585
R530 B.n789 B.n47 585
R531 B.n787 B.n786 585
R532 B.n788 B.n787 585
R533 B.n785 B.n52 585
R534 B.n52 B.n51 585
R535 B.n784 B.n783 585
R536 B.n783 B.n782 585
R537 B.n54 B.n53 585
R538 B.n781 B.n54 585
R539 B.n779 B.n778 585
R540 B.n780 B.n779 585
R541 B.n777 B.n59 585
R542 B.n59 B.n58 585
R543 B.n776 B.n775 585
R544 B.n775 B.n774 585
R545 B.n61 B.n60 585
R546 B.n773 B.n61 585
R547 B.n771 B.n770 585
R548 B.n772 B.n771 585
R549 B.n769 B.n66 585
R550 B.n66 B.n65 585
R551 B.n768 B.n767 585
R552 B.n767 B.n766 585
R553 B.n840 B.n839 585
R554 B.n838 B.n2 585
R555 B.n767 B.n68 492.5
R556 B.n763 B.n69 492.5
R557 B.n605 B.n371 492.5
R558 B.n607 B.n369 492.5
R559 B.n118 B.t17 342.332
R560 B.n116 B.t13 342.332
R561 B.n393 B.t6 342.332
R562 B.n399 B.t10 342.332
R563 B.n765 B.n764 256.663
R564 B.n765 B.n114 256.663
R565 B.n765 B.n113 256.663
R566 B.n765 B.n112 256.663
R567 B.n765 B.n111 256.663
R568 B.n765 B.n110 256.663
R569 B.n765 B.n109 256.663
R570 B.n765 B.n108 256.663
R571 B.n765 B.n107 256.663
R572 B.n765 B.n106 256.663
R573 B.n765 B.n105 256.663
R574 B.n765 B.n104 256.663
R575 B.n765 B.n103 256.663
R576 B.n765 B.n102 256.663
R577 B.n765 B.n101 256.663
R578 B.n765 B.n100 256.663
R579 B.n765 B.n99 256.663
R580 B.n765 B.n98 256.663
R581 B.n765 B.n97 256.663
R582 B.n765 B.n96 256.663
R583 B.n765 B.n95 256.663
R584 B.n765 B.n94 256.663
R585 B.n765 B.n93 256.663
R586 B.n765 B.n92 256.663
R587 B.n765 B.n91 256.663
R588 B.n765 B.n90 256.663
R589 B.n765 B.n89 256.663
R590 B.n765 B.n88 256.663
R591 B.n765 B.n87 256.663
R592 B.n765 B.n86 256.663
R593 B.n765 B.n85 256.663
R594 B.n765 B.n84 256.663
R595 B.n765 B.n83 256.663
R596 B.n765 B.n82 256.663
R597 B.n765 B.n81 256.663
R598 B.n765 B.n80 256.663
R599 B.n765 B.n79 256.663
R600 B.n765 B.n78 256.663
R601 B.n765 B.n77 256.663
R602 B.n765 B.n76 256.663
R603 B.n765 B.n75 256.663
R604 B.n765 B.n74 256.663
R605 B.n765 B.n73 256.663
R606 B.n765 B.n72 256.663
R607 B.n765 B.n71 256.663
R608 B.n765 B.n70 256.663
R609 B.n422 B.n370 256.663
R610 B.n428 B.n370 256.663
R611 B.n430 B.n370 256.663
R612 B.n436 B.n370 256.663
R613 B.n438 B.n370 256.663
R614 B.n444 B.n370 256.663
R615 B.n446 B.n370 256.663
R616 B.n452 B.n370 256.663
R617 B.n454 B.n370 256.663
R618 B.n460 B.n370 256.663
R619 B.n462 B.n370 256.663
R620 B.n468 B.n370 256.663
R621 B.n470 B.n370 256.663
R622 B.n476 B.n370 256.663
R623 B.n478 B.n370 256.663
R624 B.n484 B.n370 256.663
R625 B.n486 B.n370 256.663
R626 B.n492 B.n370 256.663
R627 B.n494 B.n370 256.663
R628 B.n500 B.n370 256.663
R629 B.n502 B.n370 256.663
R630 B.n508 B.n370 256.663
R631 B.n510 B.n370 256.663
R632 B.n516 B.n370 256.663
R633 B.n518 B.n370 256.663
R634 B.n525 B.n370 256.663
R635 B.n527 B.n370 256.663
R636 B.n533 B.n370 256.663
R637 B.n535 B.n370 256.663
R638 B.n541 B.n370 256.663
R639 B.n543 B.n370 256.663
R640 B.n549 B.n370 256.663
R641 B.n551 B.n370 256.663
R642 B.n557 B.n370 256.663
R643 B.n559 B.n370 256.663
R644 B.n565 B.n370 256.663
R645 B.n567 B.n370 256.663
R646 B.n573 B.n370 256.663
R647 B.n575 B.n370 256.663
R648 B.n581 B.n370 256.663
R649 B.n583 B.n370 256.663
R650 B.n589 B.n370 256.663
R651 B.n591 B.n370 256.663
R652 B.n597 B.n370 256.663
R653 B.n600 B.n370 256.663
R654 B.n842 B.n841 256.663
R655 B.n122 B.n121 163.367
R656 B.n126 B.n125 163.367
R657 B.n130 B.n129 163.367
R658 B.n134 B.n133 163.367
R659 B.n138 B.n137 163.367
R660 B.n142 B.n141 163.367
R661 B.n146 B.n145 163.367
R662 B.n150 B.n149 163.367
R663 B.n154 B.n153 163.367
R664 B.n158 B.n157 163.367
R665 B.n162 B.n161 163.367
R666 B.n166 B.n165 163.367
R667 B.n170 B.n169 163.367
R668 B.n174 B.n173 163.367
R669 B.n178 B.n177 163.367
R670 B.n182 B.n181 163.367
R671 B.n186 B.n185 163.367
R672 B.n190 B.n189 163.367
R673 B.n194 B.n193 163.367
R674 B.n198 B.n197 163.367
R675 B.n203 B.n202 163.367
R676 B.n207 B.n206 163.367
R677 B.n211 B.n210 163.367
R678 B.n215 B.n214 163.367
R679 B.n219 B.n218 163.367
R680 B.n224 B.n223 163.367
R681 B.n228 B.n227 163.367
R682 B.n232 B.n231 163.367
R683 B.n236 B.n235 163.367
R684 B.n240 B.n239 163.367
R685 B.n244 B.n243 163.367
R686 B.n248 B.n247 163.367
R687 B.n252 B.n251 163.367
R688 B.n256 B.n255 163.367
R689 B.n260 B.n259 163.367
R690 B.n264 B.n263 163.367
R691 B.n268 B.n267 163.367
R692 B.n272 B.n271 163.367
R693 B.n276 B.n275 163.367
R694 B.n280 B.n279 163.367
R695 B.n284 B.n283 163.367
R696 B.n288 B.n287 163.367
R697 B.n292 B.n291 163.367
R698 B.n296 B.n295 163.367
R699 B.n298 B.n115 163.367
R700 B.n605 B.n365 163.367
R701 B.n613 B.n365 163.367
R702 B.n613 B.n363 163.367
R703 B.n617 B.n363 163.367
R704 B.n617 B.n357 163.367
R705 B.n625 B.n357 163.367
R706 B.n625 B.n355 163.367
R707 B.n629 B.n355 163.367
R708 B.n629 B.n349 163.367
R709 B.n637 B.n349 163.367
R710 B.n637 B.n347 163.367
R711 B.n641 B.n347 163.367
R712 B.n641 B.n341 163.367
R713 B.n649 B.n341 163.367
R714 B.n649 B.n339 163.367
R715 B.n653 B.n339 163.367
R716 B.n653 B.n334 163.367
R717 B.n662 B.n334 163.367
R718 B.n662 B.n332 163.367
R719 B.n666 B.n332 163.367
R720 B.n666 B.n326 163.367
R721 B.n674 B.n326 163.367
R722 B.n674 B.n324 163.367
R723 B.n678 B.n324 163.367
R724 B.n678 B.n318 163.367
R725 B.n686 B.n318 163.367
R726 B.n686 B.n316 163.367
R727 B.n690 B.n316 163.367
R728 B.n690 B.n309 163.367
R729 B.n698 B.n309 163.367
R730 B.n698 B.n307 163.367
R731 B.n703 B.n307 163.367
R732 B.n703 B.n302 163.367
R733 B.n711 B.n302 163.367
R734 B.n712 B.n711 163.367
R735 B.n712 B.n5 163.367
R736 B.n6 B.n5 163.367
R737 B.n7 B.n6 163.367
R738 B.n718 B.n7 163.367
R739 B.n719 B.n718 163.367
R740 B.n719 B.n13 163.367
R741 B.n14 B.n13 163.367
R742 B.n15 B.n14 163.367
R743 B.n724 B.n15 163.367
R744 B.n724 B.n20 163.367
R745 B.n21 B.n20 163.367
R746 B.n22 B.n21 163.367
R747 B.n729 B.n22 163.367
R748 B.n729 B.n27 163.367
R749 B.n28 B.n27 163.367
R750 B.n29 B.n28 163.367
R751 B.n734 B.n29 163.367
R752 B.n734 B.n34 163.367
R753 B.n35 B.n34 163.367
R754 B.n36 B.n35 163.367
R755 B.n739 B.n36 163.367
R756 B.n739 B.n41 163.367
R757 B.n42 B.n41 163.367
R758 B.n43 B.n42 163.367
R759 B.n744 B.n43 163.367
R760 B.n744 B.n48 163.367
R761 B.n49 B.n48 163.367
R762 B.n50 B.n49 163.367
R763 B.n749 B.n50 163.367
R764 B.n749 B.n55 163.367
R765 B.n56 B.n55 163.367
R766 B.n57 B.n56 163.367
R767 B.n754 B.n57 163.367
R768 B.n754 B.n62 163.367
R769 B.n63 B.n62 163.367
R770 B.n64 B.n63 163.367
R771 B.n759 B.n64 163.367
R772 B.n759 B.n69 163.367
R773 B.n423 B.n421 163.367
R774 B.n427 B.n421 163.367
R775 B.n431 B.n429 163.367
R776 B.n435 B.n419 163.367
R777 B.n439 B.n437 163.367
R778 B.n443 B.n417 163.367
R779 B.n447 B.n445 163.367
R780 B.n451 B.n415 163.367
R781 B.n455 B.n453 163.367
R782 B.n459 B.n413 163.367
R783 B.n463 B.n461 163.367
R784 B.n467 B.n411 163.367
R785 B.n471 B.n469 163.367
R786 B.n475 B.n409 163.367
R787 B.n479 B.n477 163.367
R788 B.n483 B.n407 163.367
R789 B.n487 B.n485 163.367
R790 B.n491 B.n405 163.367
R791 B.n495 B.n493 163.367
R792 B.n499 B.n403 163.367
R793 B.n503 B.n501 163.367
R794 B.n507 B.n398 163.367
R795 B.n511 B.n509 163.367
R796 B.n515 B.n396 163.367
R797 B.n519 B.n517 163.367
R798 B.n524 B.n392 163.367
R799 B.n528 B.n526 163.367
R800 B.n532 B.n390 163.367
R801 B.n536 B.n534 163.367
R802 B.n540 B.n388 163.367
R803 B.n544 B.n542 163.367
R804 B.n548 B.n386 163.367
R805 B.n552 B.n550 163.367
R806 B.n556 B.n384 163.367
R807 B.n560 B.n558 163.367
R808 B.n564 B.n382 163.367
R809 B.n568 B.n566 163.367
R810 B.n572 B.n380 163.367
R811 B.n576 B.n574 163.367
R812 B.n580 B.n378 163.367
R813 B.n584 B.n582 163.367
R814 B.n588 B.n376 163.367
R815 B.n592 B.n590 163.367
R816 B.n596 B.n374 163.367
R817 B.n599 B.n598 163.367
R818 B.n601 B.n371 163.367
R819 B.n607 B.n367 163.367
R820 B.n611 B.n367 163.367
R821 B.n611 B.n361 163.367
R822 B.n619 B.n361 163.367
R823 B.n619 B.n359 163.367
R824 B.n623 B.n359 163.367
R825 B.n623 B.n353 163.367
R826 B.n631 B.n353 163.367
R827 B.n631 B.n351 163.367
R828 B.n635 B.n351 163.367
R829 B.n635 B.n345 163.367
R830 B.n643 B.n345 163.367
R831 B.n643 B.n343 163.367
R832 B.n647 B.n343 163.367
R833 B.n647 B.n337 163.367
R834 B.n656 B.n337 163.367
R835 B.n656 B.n335 163.367
R836 B.n660 B.n335 163.367
R837 B.n660 B.n330 163.367
R838 B.n668 B.n330 163.367
R839 B.n668 B.n328 163.367
R840 B.n672 B.n328 163.367
R841 B.n672 B.n322 163.367
R842 B.n680 B.n322 163.367
R843 B.n680 B.n320 163.367
R844 B.n684 B.n320 163.367
R845 B.n684 B.n314 163.367
R846 B.n692 B.n314 163.367
R847 B.n692 B.n312 163.367
R848 B.n696 B.n312 163.367
R849 B.n696 B.n306 163.367
R850 B.n705 B.n306 163.367
R851 B.n705 B.n304 163.367
R852 B.n709 B.n304 163.367
R853 B.n709 B.n3 163.367
R854 B.n840 B.n3 163.367
R855 B.n836 B.n2 163.367
R856 B.n836 B.n835 163.367
R857 B.n835 B.n9 163.367
R858 B.n831 B.n9 163.367
R859 B.n831 B.n11 163.367
R860 B.n827 B.n11 163.367
R861 B.n827 B.n17 163.367
R862 B.n823 B.n17 163.367
R863 B.n823 B.n19 163.367
R864 B.n819 B.n19 163.367
R865 B.n819 B.n24 163.367
R866 B.n815 B.n24 163.367
R867 B.n815 B.n26 163.367
R868 B.n811 B.n26 163.367
R869 B.n811 B.n31 163.367
R870 B.n807 B.n31 163.367
R871 B.n807 B.n33 163.367
R872 B.n803 B.n33 163.367
R873 B.n803 B.n37 163.367
R874 B.n799 B.n37 163.367
R875 B.n799 B.n39 163.367
R876 B.n795 B.n39 163.367
R877 B.n795 B.n45 163.367
R878 B.n791 B.n45 163.367
R879 B.n791 B.n47 163.367
R880 B.n787 B.n47 163.367
R881 B.n787 B.n52 163.367
R882 B.n783 B.n52 163.367
R883 B.n783 B.n54 163.367
R884 B.n779 B.n54 163.367
R885 B.n779 B.n59 163.367
R886 B.n775 B.n59 163.367
R887 B.n775 B.n61 163.367
R888 B.n771 B.n61 163.367
R889 B.n771 B.n66 163.367
R890 B.n767 B.n66 163.367
R891 B.n116 B.t15 119.215
R892 B.n393 B.t9 119.215
R893 B.n118 B.t18 119.2
R894 B.n399 B.t12 119.2
R895 B.n606 B.n370 88.3617
R896 B.n766 B.n765 88.3617
R897 B.n117 B.t16 72.0869
R898 B.n394 B.t8 72.0869
R899 B.n119 B.t19 72.0721
R900 B.n400 B.t11 72.0721
R901 B.n70 B.n68 71.676
R902 B.n122 B.n71 71.676
R903 B.n126 B.n72 71.676
R904 B.n130 B.n73 71.676
R905 B.n134 B.n74 71.676
R906 B.n138 B.n75 71.676
R907 B.n142 B.n76 71.676
R908 B.n146 B.n77 71.676
R909 B.n150 B.n78 71.676
R910 B.n154 B.n79 71.676
R911 B.n158 B.n80 71.676
R912 B.n162 B.n81 71.676
R913 B.n166 B.n82 71.676
R914 B.n170 B.n83 71.676
R915 B.n174 B.n84 71.676
R916 B.n178 B.n85 71.676
R917 B.n182 B.n86 71.676
R918 B.n186 B.n87 71.676
R919 B.n190 B.n88 71.676
R920 B.n194 B.n89 71.676
R921 B.n198 B.n90 71.676
R922 B.n203 B.n91 71.676
R923 B.n207 B.n92 71.676
R924 B.n211 B.n93 71.676
R925 B.n215 B.n94 71.676
R926 B.n219 B.n95 71.676
R927 B.n224 B.n96 71.676
R928 B.n228 B.n97 71.676
R929 B.n232 B.n98 71.676
R930 B.n236 B.n99 71.676
R931 B.n240 B.n100 71.676
R932 B.n244 B.n101 71.676
R933 B.n248 B.n102 71.676
R934 B.n252 B.n103 71.676
R935 B.n256 B.n104 71.676
R936 B.n260 B.n105 71.676
R937 B.n264 B.n106 71.676
R938 B.n268 B.n107 71.676
R939 B.n272 B.n108 71.676
R940 B.n276 B.n109 71.676
R941 B.n280 B.n110 71.676
R942 B.n284 B.n111 71.676
R943 B.n288 B.n112 71.676
R944 B.n292 B.n113 71.676
R945 B.n296 B.n114 71.676
R946 B.n764 B.n115 71.676
R947 B.n764 B.n763 71.676
R948 B.n298 B.n114 71.676
R949 B.n295 B.n113 71.676
R950 B.n291 B.n112 71.676
R951 B.n287 B.n111 71.676
R952 B.n283 B.n110 71.676
R953 B.n279 B.n109 71.676
R954 B.n275 B.n108 71.676
R955 B.n271 B.n107 71.676
R956 B.n267 B.n106 71.676
R957 B.n263 B.n105 71.676
R958 B.n259 B.n104 71.676
R959 B.n255 B.n103 71.676
R960 B.n251 B.n102 71.676
R961 B.n247 B.n101 71.676
R962 B.n243 B.n100 71.676
R963 B.n239 B.n99 71.676
R964 B.n235 B.n98 71.676
R965 B.n231 B.n97 71.676
R966 B.n227 B.n96 71.676
R967 B.n223 B.n95 71.676
R968 B.n218 B.n94 71.676
R969 B.n214 B.n93 71.676
R970 B.n210 B.n92 71.676
R971 B.n206 B.n91 71.676
R972 B.n202 B.n90 71.676
R973 B.n197 B.n89 71.676
R974 B.n193 B.n88 71.676
R975 B.n189 B.n87 71.676
R976 B.n185 B.n86 71.676
R977 B.n181 B.n85 71.676
R978 B.n177 B.n84 71.676
R979 B.n173 B.n83 71.676
R980 B.n169 B.n82 71.676
R981 B.n165 B.n81 71.676
R982 B.n161 B.n80 71.676
R983 B.n157 B.n79 71.676
R984 B.n153 B.n78 71.676
R985 B.n149 B.n77 71.676
R986 B.n145 B.n76 71.676
R987 B.n141 B.n75 71.676
R988 B.n137 B.n74 71.676
R989 B.n133 B.n73 71.676
R990 B.n129 B.n72 71.676
R991 B.n125 B.n71 71.676
R992 B.n121 B.n70 71.676
R993 B.n422 B.n369 71.676
R994 B.n428 B.n427 71.676
R995 B.n431 B.n430 71.676
R996 B.n436 B.n435 71.676
R997 B.n439 B.n438 71.676
R998 B.n444 B.n443 71.676
R999 B.n447 B.n446 71.676
R1000 B.n452 B.n451 71.676
R1001 B.n455 B.n454 71.676
R1002 B.n460 B.n459 71.676
R1003 B.n463 B.n462 71.676
R1004 B.n468 B.n467 71.676
R1005 B.n471 B.n470 71.676
R1006 B.n476 B.n475 71.676
R1007 B.n479 B.n478 71.676
R1008 B.n484 B.n483 71.676
R1009 B.n487 B.n486 71.676
R1010 B.n492 B.n491 71.676
R1011 B.n495 B.n494 71.676
R1012 B.n500 B.n499 71.676
R1013 B.n503 B.n502 71.676
R1014 B.n508 B.n507 71.676
R1015 B.n511 B.n510 71.676
R1016 B.n516 B.n515 71.676
R1017 B.n519 B.n518 71.676
R1018 B.n525 B.n524 71.676
R1019 B.n528 B.n527 71.676
R1020 B.n533 B.n532 71.676
R1021 B.n536 B.n535 71.676
R1022 B.n541 B.n540 71.676
R1023 B.n544 B.n543 71.676
R1024 B.n549 B.n548 71.676
R1025 B.n552 B.n551 71.676
R1026 B.n557 B.n556 71.676
R1027 B.n560 B.n559 71.676
R1028 B.n565 B.n564 71.676
R1029 B.n568 B.n567 71.676
R1030 B.n573 B.n572 71.676
R1031 B.n576 B.n575 71.676
R1032 B.n581 B.n580 71.676
R1033 B.n584 B.n583 71.676
R1034 B.n589 B.n588 71.676
R1035 B.n592 B.n591 71.676
R1036 B.n597 B.n596 71.676
R1037 B.n600 B.n599 71.676
R1038 B.n423 B.n422 71.676
R1039 B.n429 B.n428 71.676
R1040 B.n430 B.n419 71.676
R1041 B.n437 B.n436 71.676
R1042 B.n438 B.n417 71.676
R1043 B.n445 B.n444 71.676
R1044 B.n446 B.n415 71.676
R1045 B.n453 B.n452 71.676
R1046 B.n454 B.n413 71.676
R1047 B.n461 B.n460 71.676
R1048 B.n462 B.n411 71.676
R1049 B.n469 B.n468 71.676
R1050 B.n470 B.n409 71.676
R1051 B.n477 B.n476 71.676
R1052 B.n478 B.n407 71.676
R1053 B.n485 B.n484 71.676
R1054 B.n486 B.n405 71.676
R1055 B.n493 B.n492 71.676
R1056 B.n494 B.n403 71.676
R1057 B.n501 B.n500 71.676
R1058 B.n502 B.n398 71.676
R1059 B.n509 B.n508 71.676
R1060 B.n510 B.n396 71.676
R1061 B.n517 B.n516 71.676
R1062 B.n518 B.n392 71.676
R1063 B.n526 B.n525 71.676
R1064 B.n527 B.n390 71.676
R1065 B.n534 B.n533 71.676
R1066 B.n535 B.n388 71.676
R1067 B.n542 B.n541 71.676
R1068 B.n543 B.n386 71.676
R1069 B.n550 B.n549 71.676
R1070 B.n551 B.n384 71.676
R1071 B.n558 B.n557 71.676
R1072 B.n559 B.n382 71.676
R1073 B.n566 B.n565 71.676
R1074 B.n567 B.n380 71.676
R1075 B.n574 B.n573 71.676
R1076 B.n575 B.n378 71.676
R1077 B.n582 B.n581 71.676
R1078 B.n583 B.n376 71.676
R1079 B.n590 B.n589 71.676
R1080 B.n591 B.n374 71.676
R1081 B.n598 B.n597 71.676
R1082 B.n601 B.n600 71.676
R1083 B.n841 B.n840 71.676
R1084 B.n841 B.n2 71.676
R1085 B.n200 B.n119 59.5399
R1086 B.n221 B.n117 59.5399
R1087 B.n522 B.n394 59.5399
R1088 B.n401 B.n400 59.5399
R1089 B.n119 B.n118 47.1278
R1090 B.n117 B.n116 47.1278
R1091 B.n394 B.n393 47.1278
R1092 B.n400 B.n399 47.1278
R1093 B.n606 B.n366 43.8586
R1094 B.n612 B.n366 43.8586
R1095 B.n612 B.n362 43.8586
R1096 B.n618 B.n362 43.8586
R1097 B.n618 B.n358 43.8586
R1098 B.n624 B.n358 43.8586
R1099 B.n630 B.n354 43.8586
R1100 B.n630 B.n350 43.8586
R1101 B.n636 B.n350 43.8586
R1102 B.n636 B.n346 43.8586
R1103 B.n642 B.n346 43.8586
R1104 B.n642 B.n342 43.8586
R1105 B.n648 B.n342 43.8586
R1106 B.n648 B.n338 43.8586
R1107 B.n655 B.n338 43.8586
R1108 B.n655 B.n654 43.8586
R1109 B.n661 B.n331 43.8586
R1110 B.n667 B.n331 43.8586
R1111 B.n667 B.n327 43.8586
R1112 B.n673 B.n327 43.8586
R1113 B.n673 B.n323 43.8586
R1114 B.n679 B.n323 43.8586
R1115 B.n685 B.n319 43.8586
R1116 B.n685 B.n315 43.8586
R1117 B.n691 B.n315 43.8586
R1118 B.n691 B.n310 43.8586
R1119 B.n697 B.n310 43.8586
R1120 B.n697 B.n311 43.8586
R1121 B.n704 B.n303 43.8586
R1122 B.n710 B.n303 43.8586
R1123 B.n710 B.n4 43.8586
R1124 B.n839 B.n4 43.8586
R1125 B.n839 B.n838 43.8586
R1126 B.n838 B.n837 43.8586
R1127 B.n837 B.n8 43.8586
R1128 B.n12 B.n8 43.8586
R1129 B.n830 B.n12 43.8586
R1130 B.n829 B.n828 43.8586
R1131 B.n828 B.n16 43.8586
R1132 B.n822 B.n16 43.8586
R1133 B.n822 B.n821 43.8586
R1134 B.n821 B.n820 43.8586
R1135 B.n820 B.n23 43.8586
R1136 B.n814 B.n813 43.8586
R1137 B.n813 B.n812 43.8586
R1138 B.n812 B.n30 43.8586
R1139 B.n806 B.n30 43.8586
R1140 B.n806 B.n805 43.8586
R1141 B.n805 B.n804 43.8586
R1142 B.n798 B.n40 43.8586
R1143 B.n798 B.n797 43.8586
R1144 B.n797 B.n796 43.8586
R1145 B.n796 B.n44 43.8586
R1146 B.n790 B.n44 43.8586
R1147 B.n790 B.n789 43.8586
R1148 B.n789 B.n788 43.8586
R1149 B.n788 B.n51 43.8586
R1150 B.n782 B.n51 43.8586
R1151 B.n782 B.n781 43.8586
R1152 B.n780 B.n58 43.8586
R1153 B.n774 B.n58 43.8586
R1154 B.n774 B.n773 43.8586
R1155 B.n773 B.n772 43.8586
R1156 B.n772 B.n65 43.8586
R1157 B.n766 B.n65 43.8586
R1158 B.n661 B.t1 42.5687
R1159 B.n804 B.t0 42.5687
R1160 B.t5 B.n319 36.1189
R1161 B.t3 B.n23 36.1189
R1162 B.n608 B.n368 32.0005
R1163 B.n604 B.n603 32.0005
R1164 B.n762 B.n761 32.0005
R1165 B.n768 B.n67 32.0005
R1166 B.n624 B.t7 29.6692
R1167 B.n704 B.t2 29.6692
R1168 B.n830 B.t4 29.6692
R1169 B.t14 B.n780 29.6692
R1170 B B.n842 18.0485
R1171 B.t7 B.n354 14.1899
R1172 B.n311 B.t2 14.1899
R1173 B.t4 B.n829 14.1899
R1174 B.n781 B.t14 14.1899
R1175 B.n609 B.n608 10.6151
R1176 B.n610 B.n609 10.6151
R1177 B.n610 B.n360 10.6151
R1178 B.n620 B.n360 10.6151
R1179 B.n621 B.n620 10.6151
R1180 B.n622 B.n621 10.6151
R1181 B.n622 B.n352 10.6151
R1182 B.n632 B.n352 10.6151
R1183 B.n633 B.n632 10.6151
R1184 B.n634 B.n633 10.6151
R1185 B.n634 B.n344 10.6151
R1186 B.n644 B.n344 10.6151
R1187 B.n645 B.n644 10.6151
R1188 B.n646 B.n645 10.6151
R1189 B.n646 B.n336 10.6151
R1190 B.n657 B.n336 10.6151
R1191 B.n658 B.n657 10.6151
R1192 B.n659 B.n658 10.6151
R1193 B.n659 B.n329 10.6151
R1194 B.n669 B.n329 10.6151
R1195 B.n670 B.n669 10.6151
R1196 B.n671 B.n670 10.6151
R1197 B.n671 B.n321 10.6151
R1198 B.n681 B.n321 10.6151
R1199 B.n682 B.n681 10.6151
R1200 B.n683 B.n682 10.6151
R1201 B.n683 B.n313 10.6151
R1202 B.n693 B.n313 10.6151
R1203 B.n694 B.n693 10.6151
R1204 B.n695 B.n694 10.6151
R1205 B.n695 B.n305 10.6151
R1206 B.n706 B.n305 10.6151
R1207 B.n707 B.n706 10.6151
R1208 B.n708 B.n707 10.6151
R1209 B.n708 B.n0 10.6151
R1210 B.n424 B.n368 10.6151
R1211 B.n425 B.n424 10.6151
R1212 B.n426 B.n425 10.6151
R1213 B.n426 B.n420 10.6151
R1214 B.n432 B.n420 10.6151
R1215 B.n433 B.n432 10.6151
R1216 B.n434 B.n433 10.6151
R1217 B.n434 B.n418 10.6151
R1218 B.n440 B.n418 10.6151
R1219 B.n441 B.n440 10.6151
R1220 B.n442 B.n441 10.6151
R1221 B.n442 B.n416 10.6151
R1222 B.n448 B.n416 10.6151
R1223 B.n449 B.n448 10.6151
R1224 B.n450 B.n449 10.6151
R1225 B.n450 B.n414 10.6151
R1226 B.n456 B.n414 10.6151
R1227 B.n457 B.n456 10.6151
R1228 B.n458 B.n457 10.6151
R1229 B.n458 B.n412 10.6151
R1230 B.n464 B.n412 10.6151
R1231 B.n465 B.n464 10.6151
R1232 B.n466 B.n465 10.6151
R1233 B.n466 B.n410 10.6151
R1234 B.n472 B.n410 10.6151
R1235 B.n473 B.n472 10.6151
R1236 B.n474 B.n473 10.6151
R1237 B.n474 B.n408 10.6151
R1238 B.n480 B.n408 10.6151
R1239 B.n481 B.n480 10.6151
R1240 B.n482 B.n481 10.6151
R1241 B.n482 B.n406 10.6151
R1242 B.n488 B.n406 10.6151
R1243 B.n489 B.n488 10.6151
R1244 B.n490 B.n489 10.6151
R1245 B.n490 B.n404 10.6151
R1246 B.n496 B.n404 10.6151
R1247 B.n497 B.n496 10.6151
R1248 B.n498 B.n497 10.6151
R1249 B.n498 B.n402 10.6151
R1250 B.n505 B.n504 10.6151
R1251 B.n506 B.n505 10.6151
R1252 B.n506 B.n397 10.6151
R1253 B.n512 B.n397 10.6151
R1254 B.n513 B.n512 10.6151
R1255 B.n514 B.n513 10.6151
R1256 B.n514 B.n395 10.6151
R1257 B.n520 B.n395 10.6151
R1258 B.n521 B.n520 10.6151
R1259 B.n523 B.n391 10.6151
R1260 B.n529 B.n391 10.6151
R1261 B.n530 B.n529 10.6151
R1262 B.n531 B.n530 10.6151
R1263 B.n531 B.n389 10.6151
R1264 B.n537 B.n389 10.6151
R1265 B.n538 B.n537 10.6151
R1266 B.n539 B.n538 10.6151
R1267 B.n539 B.n387 10.6151
R1268 B.n545 B.n387 10.6151
R1269 B.n546 B.n545 10.6151
R1270 B.n547 B.n546 10.6151
R1271 B.n547 B.n385 10.6151
R1272 B.n553 B.n385 10.6151
R1273 B.n554 B.n553 10.6151
R1274 B.n555 B.n554 10.6151
R1275 B.n555 B.n383 10.6151
R1276 B.n561 B.n383 10.6151
R1277 B.n562 B.n561 10.6151
R1278 B.n563 B.n562 10.6151
R1279 B.n563 B.n381 10.6151
R1280 B.n569 B.n381 10.6151
R1281 B.n570 B.n569 10.6151
R1282 B.n571 B.n570 10.6151
R1283 B.n571 B.n379 10.6151
R1284 B.n577 B.n379 10.6151
R1285 B.n578 B.n577 10.6151
R1286 B.n579 B.n578 10.6151
R1287 B.n579 B.n377 10.6151
R1288 B.n585 B.n377 10.6151
R1289 B.n586 B.n585 10.6151
R1290 B.n587 B.n586 10.6151
R1291 B.n587 B.n375 10.6151
R1292 B.n593 B.n375 10.6151
R1293 B.n594 B.n593 10.6151
R1294 B.n595 B.n594 10.6151
R1295 B.n595 B.n373 10.6151
R1296 B.n373 B.n372 10.6151
R1297 B.n602 B.n372 10.6151
R1298 B.n603 B.n602 10.6151
R1299 B.n604 B.n364 10.6151
R1300 B.n614 B.n364 10.6151
R1301 B.n615 B.n614 10.6151
R1302 B.n616 B.n615 10.6151
R1303 B.n616 B.n356 10.6151
R1304 B.n626 B.n356 10.6151
R1305 B.n627 B.n626 10.6151
R1306 B.n628 B.n627 10.6151
R1307 B.n628 B.n348 10.6151
R1308 B.n638 B.n348 10.6151
R1309 B.n639 B.n638 10.6151
R1310 B.n640 B.n639 10.6151
R1311 B.n640 B.n340 10.6151
R1312 B.n650 B.n340 10.6151
R1313 B.n651 B.n650 10.6151
R1314 B.n652 B.n651 10.6151
R1315 B.n652 B.n333 10.6151
R1316 B.n663 B.n333 10.6151
R1317 B.n664 B.n663 10.6151
R1318 B.n665 B.n664 10.6151
R1319 B.n665 B.n325 10.6151
R1320 B.n675 B.n325 10.6151
R1321 B.n676 B.n675 10.6151
R1322 B.n677 B.n676 10.6151
R1323 B.n677 B.n317 10.6151
R1324 B.n687 B.n317 10.6151
R1325 B.n688 B.n687 10.6151
R1326 B.n689 B.n688 10.6151
R1327 B.n689 B.n308 10.6151
R1328 B.n699 B.n308 10.6151
R1329 B.n700 B.n699 10.6151
R1330 B.n702 B.n700 10.6151
R1331 B.n702 B.n701 10.6151
R1332 B.n701 B.n301 10.6151
R1333 B.n713 B.n301 10.6151
R1334 B.n714 B.n713 10.6151
R1335 B.n715 B.n714 10.6151
R1336 B.n716 B.n715 10.6151
R1337 B.n717 B.n716 10.6151
R1338 B.n720 B.n717 10.6151
R1339 B.n721 B.n720 10.6151
R1340 B.n722 B.n721 10.6151
R1341 B.n723 B.n722 10.6151
R1342 B.n725 B.n723 10.6151
R1343 B.n726 B.n725 10.6151
R1344 B.n727 B.n726 10.6151
R1345 B.n728 B.n727 10.6151
R1346 B.n730 B.n728 10.6151
R1347 B.n731 B.n730 10.6151
R1348 B.n732 B.n731 10.6151
R1349 B.n733 B.n732 10.6151
R1350 B.n735 B.n733 10.6151
R1351 B.n736 B.n735 10.6151
R1352 B.n737 B.n736 10.6151
R1353 B.n738 B.n737 10.6151
R1354 B.n740 B.n738 10.6151
R1355 B.n741 B.n740 10.6151
R1356 B.n742 B.n741 10.6151
R1357 B.n743 B.n742 10.6151
R1358 B.n745 B.n743 10.6151
R1359 B.n746 B.n745 10.6151
R1360 B.n747 B.n746 10.6151
R1361 B.n748 B.n747 10.6151
R1362 B.n750 B.n748 10.6151
R1363 B.n751 B.n750 10.6151
R1364 B.n752 B.n751 10.6151
R1365 B.n753 B.n752 10.6151
R1366 B.n755 B.n753 10.6151
R1367 B.n756 B.n755 10.6151
R1368 B.n757 B.n756 10.6151
R1369 B.n758 B.n757 10.6151
R1370 B.n760 B.n758 10.6151
R1371 B.n761 B.n760 10.6151
R1372 B.n834 B.n1 10.6151
R1373 B.n834 B.n833 10.6151
R1374 B.n833 B.n832 10.6151
R1375 B.n832 B.n10 10.6151
R1376 B.n826 B.n10 10.6151
R1377 B.n826 B.n825 10.6151
R1378 B.n825 B.n824 10.6151
R1379 B.n824 B.n18 10.6151
R1380 B.n818 B.n18 10.6151
R1381 B.n818 B.n817 10.6151
R1382 B.n817 B.n816 10.6151
R1383 B.n816 B.n25 10.6151
R1384 B.n810 B.n25 10.6151
R1385 B.n810 B.n809 10.6151
R1386 B.n809 B.n808 10.6151
R1387 B.n808 B.n32 10.6151
R1388 B.n802 B.n32 10.6151
R1389 B.n802 B.n801 10.6151
R1390 B.n801 B.n800 10.6151
R1391 B.n800 B.n38 10.6151
R1392 B.n794 B.n38 10.6151
R1393 B.n794 B.n793 10.6151
R1394 B.n793 B.n792 10.6151
R1395 B.n792 B.n46 10.6151
R1396 B.n786 B.n46 10.6151
R1397 B.n786 B.n785 10.6151
R1398 B.n785 B.n784 10.6151
R1399 B.n784 B.n53 10.6151
R1400 B.n778 B.n53 10.6151
R1401 B.n778 B.n777 10.6151
R1402 B.n777 B.n776 10.6151
R1403 B.n776 B.n60 10.6151
R1404 B.n770 B.n60 10.6151
R1405 B.n770 B.n769 10.6151
R1406 B.n769 B.n768 10.6151
R1407 B.n120 B.n67 10.6151
R1408 B.n123 B.n120 10.6151
R1409 B.n124 B.n123 10.6151
R1410 B.n127 B.n124 10.6151
R1411 B.n128 B.n127 10.6151
R1412 B.n131 B.n128 10.6151
R1413 B.n132 B.n131 10.6151
R1414 B.n135 B.n132 10.6151
R1415 B.n136 B.n135 10.6151
R1416 B.n139 B.n136 10.6151
R1417 B.n140 B.n139 10.6151
R1418 B.n143 B.n140 10.6151
R1419 B.n144 B.n143 10.6151
R1420 B.n147 B.n144 10.6151
R1421 B.n148 B.n147 10.6151
R1422 B.n151 B.n148 10.6151
R1423 B.n152 B.n151 10.6151
R1424 B.n155 B.n152 10.6151
R1425 B.n156 B.n155 10.6151
R1426 B.n159 B.n156 10.6151
R1427 B.n160 B.n159 10.6151
R1428 B.n163 B.n160 10.6151
R1429 B.n164 B.n163 10.6151
R1430 B.n167 B.n164 10.6151
R1431 B.n168 B.n167 10.6151
R1432 B.n171 B.n168 10.6151
R1433 B.n172 B.n171 10.6151
R1434 B.n175 B.n172 10.6151
R1435 B.n176 B.n175 10.6151
R1436 B.n179 B.n176 10.6151
R1437 B.n180 B.n179 10.6151
R1438 B.n183 B.n180 10.6151
R1439 B.n184 B.n183 10.6151
R1440 B.n187 B.n184 10.6151
R1441 B.n188 B.n187 10.6151
R1442 B.n191 B.n188 10.6151
R1443 B.n192 B.n191 10.6151
R1444 B.n195 B.n192 10.6151
R1445 B.n196 B.n195 10.6151
R1446 B.n199 B.n196 10.6151
R1447 B.n204 B.n201 10.6151
R1448 B.n205 B.n204 10.6151
R1449 B.n208 B.n205 10.6151
R1450 B.n209 B.n208 10.6151
R1451 B.n212 B.n209 10.6151
R1452 B.n213 B.n212 10.6151
R1453 B.n216 B.n213 10.6151
R1454 B.n217 B.n216 10.6151
R1455 B.n220 B.n217 10.6151
R1456 B.n225 B.n222 10.6151
R1457 B.n226 B.n225 10.6151
R1458 B.n229 B.n226 10.6151
R1459 B.n230 B.n229 10.6151
R1460 B.n233 B.n230 10.6151
R1461 B.n234 B.n233 10.6151
R1462 B.n237 B.n234 10.6151
R1463 B.n238 B.n237 10.6151
R1464 B.n241 B.n238 10.6151
R1465 B.n242 B.n241 10.6151
R1466 B.n245 B.n242 10.6151
R1467 B.n246 B.n245 10.6151
R1468 B.n249 B.n246 10.6151
R1469 B.n250 B.n249 10.6151
R1470 B.n253 B.n250 10.6151
R1471 B.n254 B.n253 10.6151
R1472 B.n257 B.n254 10.6151
R1473 B.n258 B.n257 10.6151
R1474 B.n261 B.n258 10.6151
R1475 B.n262 B.n261 10.6151
R1476 B.n265 B.n262 10.6151
R1477 B.n266 B.n265 10.6151
R1478 B.n269 B.n266 10.6151
R1479 B.n270 B.n269 10.6151
R1480 B.n273 B.n270 10.6151
R1481 B.n274 B.n273 10.6151
R1482 B.n277 B.n274 10.6151
R1483 B.n278 B.n277 10.6151
R1484 B.n281 B.n278 10.6151
R1485 B.n282 B.n281 10.6151
R1486 B.n285 B.n282 10.6151
R1487 B.n286 B.n285 10.6151
R1488 B.n289 B.n286 10.6151
R1489 B.n290 B.n289 10.6151
R1490 B.n293 B.n290 10.6151
R1491 B.n294 B.n293 10.6151
R1492 B.n297 B.n294 10.6151
R1493 B.n299 B.n297 10.6151
R1494 B.n300 B.n299 10.6151
R1495 B.n762 B.n300 10.6151
R1496 B.n402 B.n401 9.36635
R1497 B.n523 B.n522 9.36635
R1498 B.n200 B.n199 9.36635
R1499 B.n222 B.n221 9.36635
R1500 B.n842 B.n0 8.11757
R1501 B.n842 B.n1 8.11757
R1502 B.n679 B.t5 7.74017
R1503 B.n814 B.t3 7.74017
R1504 B.n654 B.t1 1.29044
R1505 B.n40 B.t0 1.29044
R1506 B.n504 B.n401 1.24928
R1507 B.n522 B.n521 1.24928
R1508 B.n201 B.n200 1.24928
R1509 B.n221 B.n220 1.24928
R1510 VP.n7 VP.t2 169.589
R1511 VP.n10 VP.n9 161.3
R1512 VP.n11 VP.n6 161.3
R1513 VP.n13 VP.n12 161.3
R1514 VP.n14 VP.n5 161.3
R1515 VP.n31 VP.n0 161.3
R1516 VP.n30 VP.n29 161.3
R1517 VP.n28 VP.n1 161.3
R1518 VP.n27 VP.n26 161.3
R1519 VP.n25 VP.n2 161.3
R1520 VP.n24 VP.n23 161.3
R1521 VP.n22 VP.n3 161.3
R1522 VP.n21 VP.n20 161.3
R1523 VP.n19 VP.n4 161.3
R1524 VP.n25 VP.t5 135.19
R1525 VP.n18 VP.t1 135.19
R1526 VP.n32 VP.t0 135.19
R1527 VP.n8 VP.t3 135.19
R1528 VP.n15 VP.t4 135.19
R1529 VP.n18 VP.n17 89.7593
R1530 VP.n33 VP.n32 89.7593
R1531 VP.n16 VP.n15 89.7593
R1532 VP.n20 VP.n3 56.5617
R1533 VP.n13 VP.n6 56.5617
R1534 VP.n30 VP.n1 56.5617
R1535 VP.n17 VP.n16 46.6171
R1536 VP.n8 VP.n7 46.2728
R1537 VP.n20 VP.n19 24.5923
R1538 VP.n24 VP.n3 24.5923
R1539 VP.n25 VP.n24 24.5923
R1540 VP.n26 VP.n25 24.5923
R1541 VP.n26 VP.n1 24.5923
R1542 VP.n31 VP.n30 24.5923
R1543 VP.n14 VP.n13 24.5923
R1544 VP.n9 VP.n8 24.5923
R1545 VP.n9 VP.n6 24.5923
R1546 VP.n19 VP.n18 21.1495
R1547 VP.n32 VP.n31 21.1495
R1548 VP.n15 VP.n14 21.1495
R1549 VP.n10 VP.n7 8.85089
R1550 VP.n16 VP.n5 0.278335
R1551 VP.n17 VP.n4 0.278335
R1552 VP.n33 VP.n0 0.278335
R1553 VP.n11 VP.n10 0.189894
R1554 VP.n12 VP.n11 0.189894
R1555 VP.n12 VP.n5 0.189894
R1556 VP.n21 VP.n4 0.189894
R1557 VP.n22 VP.n21 0.189894
R1558 VP.n23 VP.n22 0.189894
R1559 VP.n23 VP.n2 0.189894
R1560 VP.n27 VP.n2 0.189894
R1561 VP.n28 VP.n27 0.189894
R1562 VP.n29 VP.n28 0.189894
R1563 VP.n29 VP.n0 0.189894
R1564 VP VP.n33 0.153485
R1565 VDD1 VDD1.t3 65.678
R1566 VDD1.n1 VDD1.t4 65.5643
R1567 VDD1.n1 VDD1.n0 62.836
R1568 VDD1.n3 VDD1.n2 62.3677
R1569 VDD1.n3 VDD1.n1 42.3091
R1570 VDD1.n2 VDD1.t2 1.68131
R1571 VDD1.n2 VDD1.t1 1.68131
R1572 VDD1.n0 VDD1.t0 1.68131
R1573 VDD1.n0 VDD1.t5 1.68131
R1574 VDD1 VDD1.n3 0.466017
C0 VP VN 6.39497f
C1 VTAIL VN 6.36777f
C2 VDD1 VN 0.150463f
C3 VDD2 VP 0.416348f
C4 VDD2 VTAIL 7.673359f
C5 VDD2 VDD1 1.21513f
C6 VDD2 VN 6.31581f
C7 VP VTAIL 6.3821f
C8 VP VDD1 6.57838f
C9 VTAIL VDD1 7.62644f
C10 VDD2 B 5.568075f
C11 VDD1 B 5.866182f
C12 VTAIL B 7.394598f
C13 VN B 11.4339f
C14 VP B 9.983843f
C15 VDD1.t3 B 2.29985f
C16 VDD1.t4 B 2.29907f
C17 VDD1.t0 B 0.201847f
C18 VDD1.t5 B 0.201847f
C19 VDD1.n0 B 1.79952f
C20 VDD1.n1 B 2.41882f
C21 VDD1.t2 B 0.201847f
C22 VDD1.t1 B 0.201847f
C23 VDD1.n2 B 1.79678f
C24 VDD1.n3 B 2.28323f
C25 VP.n0 B 0.035841f
C26 VP.t0 B 1.83149f
C27 VP.n1 B 0.036888f
C28 VP.n2 B 0.027187f
C29 VP.t5 B 1.83149f
C30 VP.n3 B 0.036888f
C31 VP.n4 B 0.035841f
C32 VP.t1 B 1.83149f
C33 VP.n5 B 0.035841f
C34 VP.t4 B 1.83149f
C35 VP.n6 B 0.036888f
C36 VP.t2 B 1.9938f
C37 VP.n7 B 0.710284f
C38 VP.t3 B 1.83149f
C39 VP.n8 B 0.73447f
C40 VP.n9 B 0.050416f
C41 VP.n10 B 0.228709f
C42 VP.n11 B 0.027187f
C43 VP.n12 B 0.027187f
C44 VP.n13 B 0.042154f
C45 VP.n14 B 0.046932f
C46 VP.n15 B 0.742237f
C47 VP.n16 B 1.35041f
C48 VP.n17 B 1.37144f
C49 VP.n18 B 0.742237f
C50 VP.n19 B 0.046932f
C51 VP.n20 B 0.042154f
C52 VP.n21 B 0.027187f
C53 VP.n22 B 0.027187f
C54 VP.n23 B 0.027187f
C55 VP.n24 B 0.050416f
C56 VP.n25 B 0.67869f
C57 VP.n26 B 0.050416f
C58 VP.n27 B 0.027187f
C59 VP.n28 B 0.027187f
C60 VP.n29 B 0.027187f
C61 VP.n30 B 0.042154f
C62 VP.n31 B 0.046932f
C63 VP.n32 B 0.742237f
C64 VP.n33 B 0.03237f
C65 VDD2.t5 B 2.27954f
C66 VDD2.t3 B 0.200133f
C67 VDD2.t4 B 0.200133f
C68 VDD2.n0 B 1.78424f
C69 VDD2.n1 B 2.30273f
C70 VDD2.t0 B 2.27152f
C71 VDD2.n2 B 2.27129f
C72 VDD2.t1 B 0.200133f
C73 VDD2.t2 B 0.200133f
C74 VDD2.n3 B 1.78421f
C75 VTAIL.t11 B 0.219191f
C76 VTAIL.t7 B 0.219191f
C77 VTAIL.n0 B 1.88184f
C78 VTAIL.n1 B 0.390964f
C79 VTAIL.t2 B 2.39943f
C80 VTAIL.n2 B 0.58596f
C81 VTAIL.t1 B 0.219191f
C82 VTAIL.t5 B 0.219191f
C83 VTAIL.n3 B 1.88184f
C84 VTAIL.n4 B 1.79885f
C85 VTAIL.t9 B 0.219191f
C86 VTAIL.t10 B 0.219191f
C87 VTAIL.n5 B 1.88185f
C88 VTAIL.n6 B 1.79884f
C89 VTAIL.t6 B 2.39944f
C90 VTAIL.n7 B 0.585954f
C91 VTAIL.t4 B 0.219191f
C92 VTAIL.t3 B 0.219191f
C93 VTAIL.n8 B 1.88185f
C94 VTAIL.n9 B 0.505746f
C95 VTAIL.t0 B 2.39943f
C96 VTAIL.n10 B 1.72012f
C97 VTAIL.t8 B 2.39943f
C98 VTAIL.n11 B 1.67597f
C99 VN.n0 B 0.035218f
C100 VN.t1 B 1.79962f
C101 VN.n1 B 0.036246f
C102 VN.t0 B 1.95911f
C103 VN.n2 B 0.697925f
C104 VN.t2 B 1.79962f
C105 VN.n3 B 0.721691f
C106 VN.n4 B 0.049539f
C107 VN.n5 B 0.224729f
C108 VN.n6 B 0.026714f
C109 VN.n7 B 0.026714f
C110 VN.n8 B 0.04142f
C111 VN.n9 B 0.046115f
C112 VN.n10 B 0.729322f
C113 VN.n11 B 0.031807f
C114 VN.n12 B 0.035218f
C115 VN.t5 B 1.79962f
C116 VN.n13 B 0.036246f
C117 VN.t3 B 1.95911f
C118 VN.n14 B 0.697925f
C119 VN.t4 B 1.79962f
C120 VN.n15 B 0.721691f
C121 VN.n16 B 0.049539f
C122 VN.n17 B 0.224729f
C123 VN.n18 B 0.026714f
C124 VN.n19 B 0.026714f
C125 VN.n20 B 0.04142f
C126 VN.n21 B 0.046115f
C127 VN.n22 B 0.729322f
C128 VN.n23 B 1.34143f
.ends

