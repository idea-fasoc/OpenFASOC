* NGSPICE file created from diff_pair_sample_1052.ext - technology: sky130A

.subckt diff_pair_sample_1052 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t15 w_n2520_n4806# sky130_fd_pr__pfet_01v8 ad=3.16635 pd=19.52 as=7.4841 ps=39.16 w=19.19 l=1.22
X1 VTAIL.t9 VN.t1 VDD2.t6 w_n2520_n4806# sky130_fd_pr__pfet_01v8 ad=7.4841 pd=39.16 as=3.16635 ps=19.52 w=19.19 l=1.22
X2 VDD1.t7 VP.t0 VTAIL.t7 w_n2520_n4806# sky130_fd_pr__pfet_01v8 ad=3.16635 pd=19.52 as=7.4841 ps=39.16 w=19.19 l=1.22
X3 VDD2.t5 VN.t2 VTAIL.t8 w_n2520_n4806# sky130_fd_pr__pfet_01v8 ad=3.16635 pd=19.52 as=3.16635 ps=19.52 w=19.19 l=1.22
X4 VTAIL.t13 VN.t3 VDD2.t4 w_n2520_n4806# sky130_fd_pr__pfet_01v8 ad=7.4841 pd=39.16 as=3.16635 ps=19.52 w=19.19 l=1.22
X5 VDD1.t6 VP.t1 VTAIL.t6 w_n2520_n4806# sky130_fd_pr__pfet_01v8 ad=3.16635 pd=19.52 as=3.16635 ps=19.52 w=19.19 l=1.22
X6 VDD1.t5 VP.t2 VTAIL.t3 w_n2520_n4806# sky130_fd_pr__pfet_01v8 ad=3.16635 pd=19.52 as=3.16635 ps=19.52 w=19.19 l=1.22
X7 VTAIL.t1 VP.t3 VDD1.t4 w_n2520_n4806# sky130_fd_pr__pfet_01v8 ad=3.16635 pd=19.52 as=3.16635 ps=19.52 w=19.19 l=1.22
X8 VTAIL.t12 VN.t4 VDD2.t3 w_n2520_n4806# sky130_fd_pr__pfet_01v8 ad=3.16635 pd=19.52 as=3.16635 ps=19.52 w=19.19 l=1.22
X9 VDD1.t3 VP.t4 VTAIL.t5 w_n2520_n4806# sky130_fd_pr__pfet_01v8 ad=3.16635 pd=19.52 as=7.4841 ps=39.16 w=19.19 l=1.22
X10 B.t11 B.t9 B.t10 w_n2520_n4806# sky130_fd_pr__pfet_01v8 ad=7.4841 pd=39.16 as=0 ps=0 w=19.19 l=1.22
X11 VTAIL.t0 VP.t5 VDD1.t2 w_n2520_n4806# sky130_fd_pr__pfet_01v8 ad=7.4841 pd=39.16 as=3.16635 ps=19.52 w=19.19 l=1.22
X12 VDD2.t2 VN.t5 VTAIL.t14 w_n2520_n4806# sky130_fd_pr__pfet_01v8 ad=3.16635 pd=19.52 as=7.4841 ps=39.16 w=19.19 l=1.22
X13 B.t8 B.t6 B.t7 w_n2520_n4806# sky130_fd_pr__pfet_01v8 ad=7.4841 pd=39.16 as=0 ps=0 w=19.19 l=1.22
X14 B.t5 B.t3 B.t4 w_n2520_n4806# sky130_fd_pr__pfet_01v8 ad=7.4841 pd=39.16 as=0 ps=0 w=19.19 l=1.22
X15 VTAIL.t10 VN.t6 VDD2.t1 w_n2520_n4806# sky130_fd_pr__pfet_01v8 ad=3.16635 pd=19.52 as=3.16635 ps=19.52 w=19.19 l=1.22
X16 VTAIL.t4 VP.t6 VDD1.t1 w_n2520_n4806# sky130_fd_pr__pfet_01v8 ad=7.4841 pd=39.16 as=3.16635 ps=19.52 w=19.19 l=1.22
X17 B.t2 B.t0 B.t1 w_n2520_n4806# sky130_fd_pr__pfet_01v8 ad=7.4841 pd=39.16 as=0 ps=0 w=19.19 l=1.22
X18 VDD2.t0 VN.t7 VTAIL.t11 w_n2520_n4806# sky130_fd_pr__pfet_01v8 ad=3.16635 pd=19.52 as=3.16635 ps=19.52 w=19.19 l=1.22
X19 VTAIL.t2 VP.t7 VDD1.t0 w_n2520_n4806# sky130_fd_pr__pfet_01v8 ad=3.16635 pd=19.52 as=3.16635 ps=19.52 w=19.19 l=1.22
R0 VN.n4 VN.t3 430.61
R1 VN.n19 VN.t5 430.61
R2 VN.n13 VN.t0 411.478
R3 VN.n28 VN.t1 411.478
R4 VN.n3 VN.t7 379.082
R5 VN.n1 VN.t6 379.082
R6 VN.n18 VN.t4 379.082
R7 VN.n16 VN.t2 379.082
R8 VN.n27 VN.n15 161.3
R9 VN.n26 VN.n25 161.3
R10 VN.n24 VN.n23 161.3
R11 VN.n22 VN.n17 161.3
R12 VN.n21 VN.n20 161.3
R13 VN.n12 VN.n0 161.3
R14 VN.n11 VN.n10 161.3
R15 VN.n9 VN.n8 161.3
R16 VN.n7 VN.n2 161.3
R17 VN.n6 VN.n5 161.3
R18 VN.n29 VN.n28 80.6037
R19 VN.n14 VN.n13 80.6037
R20 VN VN.n29 50.3097
R21 VN.n4 VN.n3 44.1809
R22 VN.n19 VN.n18 44.1809
R23 VN.n7 VN.n6 40.4934
R24 VN.n8 VN.n7 40.4934
R25 VN.n22 VN.n21 40.4934
R26 VN.n23 VN.n22 40.4934
R27 VN.n12 VN.n11 35.6371
R28 VN.n27 VN.n26 35.6371
R29 VN.n13 VN.n12 31.4035
R30 VN.n28 VN.n27 31.4035
R31 VN.n20 VN.n19 29.5179
R32 VN.n5 VN.n4 29.5179
R33 VN.n6 VN.n3 13.4574
R34 VN.n8 VN.n1 13.4574
R35 VN.n21 VN.n18 13.4574
R36 VN.n23 VN.n16 13.4574
R37 VN.n11 VN.n1 11.0107
R38 VN.n26 VN.n16 11.0107
R39 VN.n29 VN.n15 0.285035
R40 VN.n14 VN.n0 0.285035
R41 VN.n25 VN.n15 0.189894
R42 VN.n25 VN.n24 0.189894
R43 VN.n24 VN.n17 0.189894
R44 VN.n20 VN.n17 0.189894
R45 VN.n5 VN.n2 0.189894
R46 VN.n9 VN.n2 0.189894
R47 VN.n10 VN.n9 0.189894
R48 VN.n10 VN.n0 0.189894
R49 VN VN.n14 0.146778
R50 VTAIL.n11 VTAIL.t0 57.4456
R51 VTAIL.n10 VTAIL.t14 57.4456
R52 VTAIL.n7 VTAIL.t9 57.4456
R53 VTAIL.n14 VTAIL.t7 57.4455
R54 VTAIL.n15 VTAIL.t15 57.4455
R55 VTAIL.n2 VTAIL.t13 57.4455
R56 VTAIL.n3 VTAIL.t5 57.4455
R57 VTAIL.n6 VTAIL.t4 57.4455
R58 VTAIL.n13 VTAIL.n12 55.7518
R59 VTAIL.n9 VTAIL.n8 55.7518
R60 VTAIL.n1 VTAIL.n0 55.7506
R61 VTAIL.n5 VTAIL.n4 55.7506
R62 VTAIL.n15 VTAIL.n14 30.2462
R63 VTAIL.n7 VTAIL.n6 30.2462
R64 VTAIL.n0 VTAIL.t11 1.69435
R65 VTAIL.n0 VTAIL.t10 1.69435
R66 VTAIL.n4 VTAIL.t3 1.69435
R67 VTAIL.n4 VTAIL.t2 1.69435
R68 VTAIL.n12 VTAIL.t6 1.69435
R69 VTAIL.n12 VTAIL.t1 1.69435
R70 VTAIL.n8 VTAIL.t8 1.69435
R71 VTAIL.n8 VTAIL.t12 1.69435
R72 VTAIL.n9 VTAIL.n7 1.33671
R73 VTAIL.n10 VTAIL.n9 1.33671
R74 VTAIL.n13 VTAIL.n11 1.33671
R75 VTAIL.n14 VTAIL.n13 1.33671
R76 VTAIL.n6 VTAIL.n5 1.33671
R77 VTAIL.n5 VTAIL.n3 1.33671
R78 VTAIL.n2 VTAIL.n1 1.33671
R79 VTAIL VTAIL.n15 1.27852
R80 VTAIL.n11 VTAIL.n10 0.470328
R81 VTAIL.n3 VTAIL.n2 0.470328
R82 VTAIL VTAIL.n1 0.0586897
R83 VDD2.n2 VDD2.n1 73.0421
R84 VDD2.n2 VDD2.n0 73.0421
R85 VDD2 VDD2.n5 73.0403
R86 VDD2.n4 VDD2.n3 72.4306
R87 VDD2.n4 VDD2.n2 46.2713
R88 VDD2.n5 VDD2.t3 1.69435
R89 VDD2.n5 VDD2.t2 1.69435
R90 VDD2.n3 VDD2.t6 1.69435
R91 VDD2.n3 VDD2.t5 1.69435
R92 VDD2.n1 VDD2.t1 1.69435
R93 VDD2.n1 VDD2.t7 1.69435
R94 VDD2.n0 VDD2.t4 1.69435
R95 VDD2.n0 VDD2.t0 1.69435
R96 VDD2 VDD2.n4 0.726793
R97 VP.n9 VP.t5 430.61
R98 VP.n21 VP.t6 411.478
R99 VP.n33 VP.t4 411.478
R100 VP.n18 VP.t0 411.478
R101 VP.n3 VP.t2 379.082
R102 VP.n1 VP.t7 379.082
R103 VP.n6 VP.t3 379.082
R104 VP.n8 VP.t1 379.082
R105 VP.n11 VP.n10 161.3
R106 VP.n12 VP.n7 161.3
R107 VP.n14 VP.n13 161.3
R108 VP.n16 VP.n15 161.3
R109 VP.n17 VP.n5 161.3
R110 VP.n32 VP.n0 161.3
R111 VP.n31 VP.n30 161.3
R112 VP.n29 VP.n28 161.3
R113 VP.n27 VP.n2 161.3
R114 VP.n26 VP.n25 161.3
R115 VP.n24 VP.n23 161.3
R116 VP.n22 VP.n4 161.3
R117 VP.n19 VP.n18 80.6037
R118 VP.n34 VP.n33 80.6037
R119 VP.n21 VP.n20 80.6037
R120 VP.n20 VP.n19 50.0241
R121 VP.n9 VP.n8 44.1809
R122 VP.n27 VP.n26 40.4934
R123 VP.n28 VP.n27 40.4934
R124 VP.n13 VP.n12 40.4934
R125 VP.n12 VP.n11 40.4934
R126 VP.n23 VP.n22 35.6371
R127 VP.n32 VP.n31 35.6371
R128 VP.n17 VP.n16 35.6371
R129 VP.n22 VP.n21 31.4035
R130 VP.n33 VP.n32 31.4035
R131 VP.n18 VP.n17 31.4035
R132 VP.n10 VP.n9 29.5179
R133 VP.n26 VP.n3 13.4574
R134 VP.n28 VP.n1 13.4574
R135 VP.n13 VP.n6 13.4574
R136 VP.n11 VP.n8 13.4574
R137 VP.n23 VP.n3 11.0107
R138 VP.n31 VP.n1 11.0107
R139 VP.n16 VP.n6 11.0107
R140 VP.n19 VP.n5 0.285035
R141 VP.n20 VP.n4 0.285035
R142 VP.n34 VP.n0 0.285035
R143 VP.n10 VP.n7 0.189894
R144 VP.n14 VP.n7 0.189894
R145 VP.n15 VP.n14 0.189894
R146 VP.n15 VP.n5 0.189894
R147 VP.n24 VP.n4 0.189894
R148 VP.n25 VP.n24 0.189894
R149 VP.n25 VP.n2 0.189894
R150 VP.n29 VP.n2 0.189894
R151 VP.n30 VP.n29 0.189894
R152 VP.n30 VP.n0 0.189894
R153 VP VP.n34 0.146778
R154 VDD1 VDD1.n0 73.1569
R155 VDD1.n3 VDD1.n2 73.0421
R156 VDD1.n3 VDD1.n1 73.0421
R157 VDD1.n5 VDD1.n4 72.4304
R158 VDD1.n5 VDD1.n3 46.8543
R159 VDD1.n4 VDD1.t4 1.69435
R160 VDD1.n4 VDD1.t7 1.69435
R161 VDD1.n0 VDD1.t2 1.69435
R162 VDD1.n0 VDD1.t6 1.69435
R163 VDD1.n2 VDD1.t0 1.69435
R164 VDD1.n2 VDD1.t3 1.69435
R165 VDD1.n1 VDD1.t1 1.69435
R166 VDD1.n1 VDD1.t5 1.69435
R167 VDD1 VDD1.n5 0.610414
R168 B.n552 B.n551 585
R169 B.n553 B.n88 585
R170 B.n555 B.n554 585
R171 B.n556 B.n87 585
R172 B.n558 B.n557 585
R173 B.n559 B.n86 585
R174 B.n561 B.n560 585
R175 B.n562 B.n85 585
R176 B.n564 B.n563 585
R177 B.n565 B.n84 585
R178 B.n567 B.n566 585
R179 B.n568 B.n83 585
R180 B.n570 B.n569 585
R181 B.n571 B.n82 585
R182 B.n573 B.n572 585
R183 B.n574 B.n81 585
R184 B.n576 B.n575 585
R185 B.n577 B.n80 585
R186 B.n579 B.n578 585
R187 B.n580 B.n79 585
R188 B.n582 B.n581 585
R189 B.n583 B.n78 585
R190 B.n585 B.n584 585
R191 B.n586 B.n77 585
R192 B.n588 B.n587 585
R193 B.n589 B.n76 585
R194 B.n591 B.n590 585
R195 B.n592 B.n75 585
R196 B.n594 B.n593 585
R197 B.n595 B.n74 585
R198 B.n597 B.n596 585
R199 B.n598 B.n73 585
R200 B.n600 B.n599 585
R201 B.n601 B.n72 585
R202 B.n603 B.n602 585
R203 B.n604 B.n71 585
R204 B.n606 B.n605 585
R205 B.n607 B.n70 585
R206 B.n609 B.n608 585
R207 B.n610 B.n69 585
R208 B.n612 B.n611 585
R209 B.n613 B.n68 585
R210 B.n615 B.n614 585
R211 B.n616 B.n67 585
R212 B.n618 B.n617 585
R213 B.n619 B.n66 585
R214 B.n621 B.n620 585
R215 B.n622 B.n65 585
R216 B.n624 B.n623 585
R217 B.n625 B.n64 585
R218 B.n627 B.n626 585
R219 B.n628 B.n63 585
R220 B.n630 B.n629 585
R221 B.n631 B.n62 585
R222 B.n633 B.n632 585
R223 B.n634 B.n61 585
R224 B.n636 B.n635 585
R225 B.n637 B.n60 585
R226 B.n639 B.n638 585
R227 B.n640 B.n59 585
R228 B.n642 B.n641 585
R229 B.n643 B.n58 585
R230 B.n645 B.n644 585
R231 B.n647 B.n55 585
R232 B.n649 B.n648 585
R233 B.n650 B.n54 585
R234 B.n652 B.n651 585
R235 B.n653 B.n53 585
R236 B.n655 B.n654 585
R237 B.n656 B.n52 585
R238 B.n658 B.n657 585
R239 B.n659 B.n49 585
R240 B.n662 B.n661 585
R241 B.n663 B.n48 585
R242 B.n665 B.n664 585
R243 B.n666 B.n47 585
R244 B.n668 B.n667 585
R245 B.n669 B.n46 585
R246 B.n671 B.n670 585
R247 B.n672 B.n45 585
R248 B.n674 B.n673 585
R249 B.n675 B.n44 585
R250 B.n677 B.n676 585
R251 B.n678 B.n43 585
R252 B.n680 B.n679 585
R253 B.n681 B.n42 585
R254 B.n683 B.n682 585
R255 B.n684 B.n41 585
R256 B.n686 B.n685 585
R257 B.n687 B.n40 585
R258 B.n689 B.n688 585
R259 B.n690 B.n39 585
R260 B.n692 B.n691 585
R261 B.n693 B.n38 585
R262 B.n695 B.n694 585
R263 B.n696 B.n37 585
R264 B.n698 B.n697 585
R265 B.n699 B.n36 585
R266 B.n701 B.n700 585
R267 B.n702 B.n35 585
R268 B.n704 B.n703 585
R269 B.n705 B.n34 585
R270 B.n707 B.n706 585
R271 B.n708 B.n33 585
R272 B.n710 B.n709 585
R273 B.n711 B.n32 585
R274 B.n713 B.n712 585
R275 B.n714 B.n31 585
R276 B.n716 B.n715 585
R277 B.n717 B.n30 585
R278 B.n719 B.n718 585
R279 B.n720 B.n29 585
R280 B.n722 B.n721 585
R281 B.n723 B.n28 585
R282 B.n725 B.n724 585
R283 B.n726 B.n27 585
R284 B.n728 B.n727 585
R285 B.n729 B.n26 585
R286 B.n731 B.n730 585
R287 B.n732 B.n25 585
R288 B.n734 B.n733 585
R289 B.n735 B.n24 585
R290 B.n737 B.n736 585
R291 B.n738 B.n23 585
R292 B.n740 B.n739 585
R293 B.n741 B.n22 585
R294 B.n743 B.n742 585
R295 B.n744 B.n21 585
R296 B.n746 B.n745 585
R297 B.n747 B.n20 585
R298 B.n749 B.n748 585
R299 B.n750 B.n19 585
R300 B.n752 B.n751 585
R301 B.n753 B.n18 585
R302 B.n755 B.n754 585
R303 B.n550 B.n89 585
R304 B.n549 B.n548 585
R305 B.n547 B.n90 585
R306 B.n546 B.n545 585
R307 B.n544 B.n91 585
R308 B.n543 B.n542 585
R309 B.n541 B.n92 585
R310 B.n540 B.n539 585
R311 B.n538 B.n93 585
R312 B.n537 B.n536 585
R313 B.n535 B.n94 585
R314 B.n534 B.n533 585
R315 B.n532 B.n95 585
R316 B.n531 B.n530 585
R317 B.n529 B.n96 585
R318 B.n528 B.n527 585
R319 B.n526 B.n97 585
R320 B.n525 B.n524 585
R321 B.n523 B.n98 585
R322 B.n522 B.n521 585
R323 B.n520 B.n99 585
R324 B.n519 B.n518 585
R325 B.n517 B.n100 585
R326 B.n516 B.n515 585
R327 B.n514 B.n101 585
R328 B.n513 B.n512 585
R329 B.n511 B.n102 585
R330 B.n510 B.n509 585
R331 B.n508 B.n103 585
R332 B.n507 B.n506 585
R333 B.n505 B.n104 585
R334 B.n504 B.n503 585
R335 B.n502 B.n105 585
R336 B.n501 B.n500 585
R337 B.n499 B.n106 585
R338 B.n498 B.n497 585
R339 B.n496 B.n107 585
R340 B.n495 B.n494 585
R341 B.n493 B.n108 585
R342 B.n492 B.n491 585
R343 B.n490 B.n109 585
R344 B.n489 B.n488 585
R345 B.n487 B.n110 585
R346 B.n486 B.n485 585
R347 B.n484 B.n111 585
R348 B.n483 B.n482 585
R349 B.n481 B.n112 585
R350 B.n480 B.n479 585
R351 B.n478 B.n113 585
R352 B.n477 B.n476 585
R353 B.n475 B.n114 585
R354 B.n474 B.n473 585
R355 B.n472 B.n115 585
R356 B.n471 B.n470 585
R357 B.n469 B.n116 585
R358 B.n468 B.n467 585
R359 B.n466 B.n117 585
R360 B.n465 B.n464 585
R361 B.n463 B.n118 585
R362 B.n462 B.n461 585
R363 B.n460 B.n119 585
R364 B.n459 B.n458 585
R365 B.n457 B.n120 585
R366 B.n253 B.n192 585
R367 B.n255 B.n254 585
R368 B.n256 B.n191 585
R369 B.n258 B.n257 585
R370 B.n259 B.n190 585
R371 B.n261 B.n260 585
R372 B.n262 B.n189 585
R373 B.n264 B.n263 585
R374 B.n265 B.n188 585
R375 B.n267 B.n266 585
R376 B.n268 B.n187 585
R377 B.n270 B.n269 585
R378 B.n271 B.n186 585
R379 B.n273 B.n272 585
R380 B.n274 B.n185 585
R381 B.n276 B.n275 585
R382 B.n277 B.n184 585
R383 B.n279 B.n278 585
R384 B.n280 B.n183 585
R385 B.n282 B.n281 585
R386 B.n283 B.n182 585
R387 B.n285 B.n284 585
R388 B.n286 B.n181 585
R389 B.n288 B.n287 585
R390 B.n289 B.n180 585
R391 B.n291 B.n290 585
R392 B.n292 B.n179 585
R393 B.n294 B.n293 585
R394 B.n295 B.n178 585
R395 B.n297 B.n296 585
R396 B.n298 B.n177 585
R397 B.n300 B.n299 585
R398 B.n301 B.n176 585
R399 B.n303 B.n302 585
R400 B.n304 B.n175 585
R401 B.n306 B.n305 585
R402 B.n307 B.n174 585
R403 B.n309 B.n308 585
R404 B.n310 B.n173 585
R405 B.n312 B.n311 585
R406 B.n313 B.n172 585
R407 B.n315 B.n314 585
R408 B.n316 B.n171 585
R409 B.n318 B.n317 585
R410 B.n319 B.n170 585
R411 B.n321 B.n320 585
R412 B.n322 B.n169 585
R413 B.n324 B.n323 585
R414 B.n325 B.n168 585
R415 B.n327 B.n326 585
R416 B.n328 B.n167 585
R417 B.n330 B.n329 585
R418 B.n331 B.n166 585
R419 B.n333 B.n332 585
R420 B.n334 B.n165 585
R421 B.n336 B.n335 585
R422 B.n337 B.n164 585
R423 B.n339 B.n338 585
R424 B.n340 B.n163 585
R425 B.n342 B.n341 585
R426 B.n343 B.n162 585
R427 B.n345 B.n344 585
R428 B.n346 B.n159 585
R429 B.n349 B.n348 585
R430 B.n350 B.n158 585
R431 B.n352 B.n351 585
R432 B.n353 B.n157 585
R433 B.n355 B.n354 585
R434 B.n356 B.n156 585
R435 B.n358 B.n357 585
R436 B.n359 B.n155 585
R437 B.n361 B.n360 585
R438 B.n363 B.n362 585
R439 B.n364 B.n151 585
R440 B.n366 B.n365 585
R441 B.n367 B.n150 585
R442 B.n369 B.n368 585
R443 B.n370 B.n149 585
R444 B.n372 B.n371 585
R445 B.n373 B.n148 585
R446 B.n375 B.n374 585
R447 B.n376 B.n147 585
R448 B.n378 B.n377 585
R449 B.n379 B.n146 585
R450 B.n381 B.n380 585
R451 B.n382 B.n145 585
R452 B.n384 B.n383 585
R453 B.n385 B.n144 585
R454 B.n387 B.n386 585
R455 B.n388 B.n143 585
R456 B.n390 B.n389 585
R457 B.n391 B.n142 585
R458 B.n393 B.n392 585
R459 B.n394 B.n141 585
R460 B.n396 B.n395 585
R461 B.n397 B.n140 585
R462 B.n399 B.n398 585
R463 B.n400 B.n139 585
R464 B.n402 B.n401 585
R465 B.n403 B.n138 585
R466 B.n405 B.n404 585
R467 B.n406 B.n137 585
R468 B.n408 B.n407 585
R469 B.n409 B.n136 585
R470 B.n411 B.n410 585
R471 B.n412 B.n135 585
R472 B.n414 B.n413 585
R473 B.n415 B.n134 585
R474 B.n417 B.n416 585
R475 B.n418 B.n133 585
R476 B.n420 B.n419 585
R477 B.n421 B.n132 585
R478 B.n423 B.n422 585
R479 B.n424 B.n131 585
R480 B.n426 B.n425 585
R481 B.n427 B.n130 585
R482 B.n429 B.n428 585
R483 B.n430 B.n129 585
R484 B.n432 B.n431 585
R485 B.n433 B.n128 585
R486 B.n435 B.n434 585
R487 B.n436 B.n127 585
R488 B.n438 B.n437 585
R489 B.n439 B.n126 585
R490 B.n441 B.n440 585
R491 B.n442 B.n125 585
R492 B.n444 B.n443 585
R493 B.n445 B.n124 585
R494 B.n447 B.n446 585
R495 B.n448 B.n123 585
R496 B.n450 B.n449 585
R497 B.n451 B.n122 585
R498 B.n453 B.n452 585
R499 B.n454 B.n121 585
R500 B.n456 B.n455 585
R501 B.n252 B.n251 585
R502 B.n250 B.n193 585
R503 B.n249 B.n248 585
R504 B.n247 B.n194 585
R505 B.n246 B.n245 585
R506 B.n244 B.n195 585
R507 B.n243 B.n242 585
R508 B.n241 B.n196 585
R509 B.n240 B.n239 585
R510 B.n238 B.n197 585
R511 B.n237 B.n236 585
R512 B.n235 B.n198 585
R513 B.n234 B.n233 585
R514 B.n232 B.n199 585
R515 B.n231 B.n230 585
R516 B.n229 B.n200 585
R517 B.n228 B.n227 585
R518 B.n226 B.n201 585
R519 B.n225 B.n224 585
R520 B.n223 B.n202 585
R521 B.n222 B.n221 585
R522 B.n220 B.n203 585
R523 B.n219 B.n218 585
R524 B.n217 B.n204 585
R525 B.n216 B.n215 585
R526 B.n214 B.n205 585
R527 B.n213 B.n212 585
R528 B.n211 B.n206 585
R529 B.n210 B.n209 585
R530 B.n208 B.n207 585
R531 B.n2 B.n0 585
R532 B.n801 B.n1 585
R533 B.n800 B.n799 585
R534 B.n798 B.n3 585
R535 B.n797 B.n796 585
R536 B.n795 B.n4 585
R537 B.n794 B.n793 585
R538 B.n792 B.n5 585
R539 B.n791 B.n790 585
R540 B.n789 B.n6 585
R541 B.n788 B.n787 585
R542 B.n786 B.n7 585
R543 B.n785 B.n784 585
R544 B.n783 B.n8 585
R545 B.n782 B.n781 585
R546 B.n780 B.n9 585
R547 B.n779 B.n778 585
R548 B.n777 B.n10 585
R549 B.n776 B.n775 585
R550 B.n774 B.n11 585
R551 B.n773 B.n772 585
R552 B.n771 B.n12 585
R553 B.n770 B.n769 585
R554 B.n768 B.n13 585
R555 B.n767 B.n766 585
R556 B.n765 B.n14 585
R557 B.n764 B.n763 585
R558 B.n762 B.n15 585
R559 B.n761 B.n760 585
R560 B.n759 B.n16 585
R561 B.n758 B.n757 585
R562 B.n756 B.n17 585
R563 B.n803 B.n802 585
R564 B.n152 B.t9 583.302
R565 B.n160 B.t0 583.302
R566 B.n50 B.t3 583.302
R567 B.n56 B.t6 583.302
R568 B.n253 B.n252 492.5
R569 B.n754 B.n17 492.5
R570 B.n457 B.n456 492.5
R571 B.n552 B.n89 492.5
R572 B.n252 B.n193 163.367
R573 B.n248 B.n193 163.367
R574 B.n248 B.n247 163.367
R575 B.n247 B.n246 163.367
R576 B.n246 B.n195 163.367
R577 B.n242 B.n195 163.367
R578 B.n242 B.n241 163.367
R579 B.n241 B.n240 163.367
R580 B.n240 B.n197 163.367
R581 B.n236 B.n197 163.367
R582 B.n236 B.n235 163.367
R583 B.n235 B.n234 163.367
R584 B.n234 B.n199 163.367
R585 B.n230 B.n199 163.367
R586 B.n230 B.n229 163.367
R587 B.n229 B.n228 163.367
R588 B.n228 B.n201 163.367
R589 B.n224 B.n201 163.367
R590 B.n224 B.n223 163.367
R591 B.n223 B.n222 163.367
R592 B.n222 B.n203 163.367
R593 B.n218 B.n203 163.367
R594 B.n218 B.n217 163.367
R595 B.n217 B.n216 163.367
R596 B.n216 B.n205 163.367
R597 B.n212 B.n205 163.367
R598 B.n212 B.n211 163.367
R599 B.n211 B.n210 163.367
R600 B.n210 B.n207 163.367
R601 B.n207 B.n2 163.367
R602 B.n802 B.n2 163.367
R603 B.n802 B.n801 163.367
R604 B.n801 B.n800 163.367
R605 B.n800 B.n3 163.367
R606 B.n796 B.n3 163.367
R607 B.n796 B.n795 163.367
R608 B.n795 B.n794 163.367
R609 B.n794 B.n5 163.367
R610 B.n790 B.n5 163.367
R611 B.n790 B.n789 163.367
R612 B.n789 B.n788 163.367
R613 B.n788 B.n7 163.367
R614 B.n784 B.n7 163.367
R615 B.n784 B.n783 163.367
R616 B.n783 B.n782 163.367
R617 B.n782 B.n9 163.367
R618 B.n778 B.n9 163.367
R619 B.n778 B.n777 163.367
R620 B.n777 B.n776 163.367
R621 B.n776 B.n11 163.367
R622 B.n772 B.n11 163.367
R623 B.n772 B.n771 163.367
R624 B.n771 B.n770 163.367
R625 B.n770 B.n13 163.367
R626 B.n766 B.n13 163.367
R627 B.n766 B.n765 163.367
R628 B.n765 B.n764 163.367
R629 B.n764 B.n15 163.367
R630 B.n760 B.n15 163.367
R631 B.n760 B.n759 163.367
R632 B.n759 B.n758 163.367
R633 B.n758 B.n17 163.367
R634 B.n254 B.n253 163.367
R635 B.n254 B.n191 163.367
R636 B.n258 B.n191 163.367
R637 B.n259 B.n258 163.367
R638 B.n260 B.n259 163.367
R639 B.n260 B.n189 163.367
R640 B.n264 B.n189 163.367
R641 B.n265 B.n264 163.367
R642 B.n266 B.n265 163.367
R643 B.n266 B.n187 163.367
R644 B.n270 B.n187 163.367
R645 B.n271 B.n270 163.367
R646 B.n272 B.n271 163.367
R647 B.n272 B.n185 163.367
R648 B.n276 B.n185 163.367
R649 B.n277 B.n276 163.367
R650 B.n278 B.n277 163.367
R651 B.n278 B.n183 163.367
R652 B.n282 B.n183 163.367
R653 B.n283 B.n282 163.367
R654 B.n284 B.n283 163.367
R655 B.n284 B.n181 163.367
R656 B.n288 B.n181 163.367
R657 B.n289 B.n288 163.367
R658 B.n290 B.n289 163.367
R659 B.n290 B.n179 163.367
R660 B.n294 B.n179 163.367
R661 B.n295 B.n294 163.367
R662 B.n296 B.n295 163.367
R663 B.n296 B.n177 163.367
R664 B.n300 B.n177 163.367
R665 B.n301 B.n300 163.367
R666 B.n302 B.n301 163.367
R667 B.n302 B.n175 163.367
R668 B.n306 B.n175 163.367
R669 B.n307 B.n306 163.367
R670 B.n308 B.n307 163.367
R671 B.n308 B.n173 163.367
R672 B.n312 B.n173 163.367
R673 B.n313 B.n312 163.367
R674 B.n314 B.n313 163.367
R675 B.n314 B.n171 163.367
R676 B.n318 B.n171 163.367
R677 B.n319 B.n318 163.367
R678 B.n320 B.n319 163.367
R679 B.n320 B.n169 163.367
R680 B.n324 B.n169 163.367
R681 B.n325 B.n324 163.367
R682 B.n326 B.n325 163.367
R683 B.n326 B.n167 163.367
R684 B.n330 B.n167 163.367
R685 B.n331 B.n330 163.367
R686 B.n332 B.n331 163.367
R687 B.n332 B.n165 163.367
R688 B.n336 B.n165 163.367
R689 B.n337 B.n336 163.367
R690 B.n338 B.n337 163.367
R691 B.n338 B.n163 163.367
R692 B.n342 B.n163 163.367
R693 B.n343 B.n342 163.367
R694 B.n344 B.n343 163.367
R695 B.n344 B.n159 163.367
R696 B.n349 B.n159 163.367
R697 B.n350 B.n349 163.367
R698 B.n351 B.n350 163.367
R699 B.n351 B.n157 163.367
R700 B.n355 B.n157 163.367
R701 B.n356 B.n355 163.367
R702 B.n357 B.n356 163.367
R703 B.n357 B.n155 163.367
R704 B.n361 B.n155 163.367
R705 B.n362 B.n361 163.367
R706 B.n362 B.n151 163.367
R707 B.n366 B.n151 163.367
R708 B.n367 B.n366 163.367
R709 B.n368 B.n367 163.367
R710 B.n368 B.n149 163.367
R711 B.n372 B.n149 163.367
R712 B.n373 B.n372 163.367
R713 B.n374 B.n373 163.367
R714 B.n374 B.n147 163.367
R715 B.n378 B.n147 163.367
R716 B.n379 B.n378 163.367
R717 B.n380 B.n379 163.367
R718 B.n380 B.n145 163.367
R719 B.n384 B.n145 163.367
R720 B.n385 B.n384 163.367
R721 B.n386 B.n385 163.367
R722 B.n386 B.n143 163.367
R723 B.n390 B.n143 163.367
R724 B.n391 B.n390 163.367
R725 B.n392 B.n391 163.367
R726 B.n392 B.n141 163.367
R727 B.n396 B.n141 163.367
R728 B.n397 B.n396 163.367
R729 B.n398 B.n397 163.367
R730 B.n398 B.n139 163.367
R731 B.n402 B.n139 163.367
R732 B.n403 B.n402 163.367
R733 B.n404 B.n403 163.367
R734 B.n404 B.n137 163.367
R735 B.n408 B.n137 163.367
R736 B.n409 B.n408 163.367
R737 B.n410 B.n409 163.367
R738 B.n410 B.n135 163.367
R739 B.n414 B.n135 163.367
R740 B.n415 B.n414 163.367
R741 B.n416 B.n415 163.367
R742 B.n416 B.n133 163.367
R743 B.n420 B.n133 163.367
R744 B.n421 B.n420 163.367
R745 B.n422 B.n421 163.367
R746 B.n422 B.n131 163.367
R747 B.n426 B.n131 163.367
R748 B.n427 B.n426 163.367
R749 B.n428 B.n427 163.367
R750 B.n428 B.n129 163.367
R751 B.n432 B.n129 163.367
R752 B.n433 B.n432 163.367
R753 B.n434 B.n433 163.367
R754 B.n434 B.n127 163.367
R755 B.n438 B.n127 163.367
R756 B.n439 B.n438 163.367
R757 B.n440 B.n439 163.367
R758 B.n440 B.n125 163.367
R759 B.n444 B.n125 163.367
R760 B.n445 B.n444 163.367
R761 B.n446 B.n445 163.367
R762 B.n446 B.n123 163.367
R763 B.n450 B.n123 163.367
R764 B.n451 B.n450 163.367
R765 B.n452 B.n451 163.367
R766 B.n452 B.n121 163.367
R767 B.n456 B.n121 163.367
R768 B.n458 B.n457 163.367
R769 B.n458 B.n119 163.367
R770 B.n462 B.n119 163.367
R771 B.n463 B.n462 163.367
R772 B.n464 B.n463 163.367
R773 B.n464 B.n117 163.367
R774 B.n468 B.n117 163.367
R775 B.n469 B.n468 163.367
R776 B.n470 B.n469 163.367
R777 B.n470 B.n115 163.367
R778 B.n474 B.n115 163.367
R779 B.n475 B.n474 163.367
R780 B.n476 B.n475 163.367
R781 B.n476 B.n113 163.367
R782 B.n480 B.n113 163.367
R783 B.n481 B.n480 163.367
R784 B.n482 B.n481 163.367
R785 B.n482 B.n111 163.367
R786 B.n486 B.n111 163.367
R787 B.n487 B.n486 163.367
R788 B.n488 B.n487 163.367
R789 B.n488 B.n109 163.367
R790 B.n492 B.n109 163.367
R791 B.n493 B.n492 163.367
R792 B.n494 B.n493 163.367
R793 B.n494 B.n107 163.367
R794 B.n498 B.n107 163.367
R795 B.n499 B.n498 163.367
R796 B.n500 B.n499 163.367
R797 B.n500 B.n105 163.367
R798 B.n504 B.n105 163.367
R799 B.n505 B.n504 163.367
R800 B.n506 B.n505 163.367
R801 B.n506 B.n103 163.367
R802 B.n510 B.n103 163.367
R803 B.n511 B.n510 163.367
R804 B.n512 B.n511 163.367
R805 B.n512 B.n101 163.367
R806 B.n516 B.n101 163.367
R807 B.n517 B.n516 163.367
R808 B.n518 B.n517 163.367
R809 B.n518 B.n99 163.367
R810 B.n522 B.n99 163.367
R811 B.n523 B.n522 163.367
R812 B.n524 B.n523 163.367
R813 B.n524 B.n97 163.367
R814 B.n528 B.n97 163.367
R815 B.n529 B.n528 163.367
R816 B.n530 B.n529 163.367
R817 B.n530 B.n95 163.367
R818 B.n534 B.n95 163.367
R819 B.n535 B.n534 163.367
R820 B.n536 B.n535 163.367
R821 B.n536 B.n93 163.367
R822 B.n540 B.n93 163.367
R823 B.n541 B.n540 163.367
R824 B.n542 B.n541 163.367
R825 B.n542 B.n91 163.367
R826 B.n546 B.n91 163.367
R827 B.n547 B.n546 163.367
R828 B.n548 B.n547 163.367
R829 B.n548 B.n89 163.367
R830 B.n754 B.n753 163.367
R831 B.n753 B.n752 163.367
R832 B.n752 B.n19 163.367
R833 B.n748 B.n19 163.367
R834 B.n748 B.n747 163.367
R835 B.n747 B.n746 163.367
R836 B.n746 B.n21 163.367
R837 B.n742 B.n21 163.367
R838 B.n742 B.n741 163.367
R839 B.n741 B.n740 163.367
R840 B.n740 B.n23 163.367
R841 B.n736 B.n23 163.367
R842 B.n736 B.n735 163.367
R843 B.n735 B.n734 163.367
R844 B.n734 B.n25 163.367
R845 B.n730 B.n25 163.367
R846 B.n730 B.n729 163.367
R847 B.n729 B.n728 163.367
R848 B.n728 B.n27 163.367
R849 B.n724 B.n27 163.367
R850 B.n724 B.n723 163.367
R851 B.n723 B.n722 163.367
R852 B.n722 B.n29 163.367
R853 B.n718 B.n29 163.367
R854 B.n718 B.n717 163.367
R855 B.n717 B.n716 163.367
R856 B.n716 B.n31 163.367
R857 B.n712 B.n31 163.367
R858 B.n712 B.n711 163.367
R859 B.n711 B.n710 163.367
R860 B.n710 B.n33 163.367
R861 B.n706 B.n33 163.367
R862 B.n706 B.n705 163.367
R863 B.n705 B.n704 163.367
R864 B.n704 B.n35 163.367
R865 B.n700 B.n35 163.367
R866 B.n700 B.n699 163.367
R867 B.n699 B.n698 163.367
R868 B.n698 B.n37 163.367
R869 B.n694 B.n37 163.367
R870 B.n694 B.n693 163.367
R871 B.n693 B.n692 163.367
R872 B.n692 B.n39 163.367
R873 B.n688 B.n39 163.367
R874 B.n688 B.n687 163.367
R875 B.n687 B.n686 163.367
R876 B.n686 B.n41 163.367
R877 B.n682 B.n41 163.367
R878 B.n682 B.n681 163.367
R879 B.n681 B.n680 163.367
R880 B.n680 B.n43 163.367
R881 B.n676 B.n43 163.367
R882 B.n676 B.n675 163.367
R883 B.n675 B.n674 163.367
R884 B.n674 B.n45 163.367
R885 B.n670 B.n45 163.367
R886 B.n670 B.n669 163.367
R887 B.n669 B.n668 163.367
R888 B.n668 B.n47 163.367
R889 B.n664 B.n47 163.367
R890 B.n664 B.n663 163.367
R891 B.n663 B.n662 163.367
R892 B.n662 B.n49 163.367
R893 B.n657 B.n49 163.367
R894 B.n657 B.n656 163.367
R895 B.n656 B.n655 163.367
R896 B.n655 B.n53 163.367
R897 B.n651 B.n53 163.367
R898 B.n651 B.n650 163.367
R899 B.n650 B.n649 163.367
R900 B.n649 B.n55 163.367
R901 B.n644 B.n55 163.367
R902 B.n644 B.n643 163.367
R903 B.n643 B.n642 163.367
R904 B.n642 B.n59 163.367
R905 B.n638 B.n59 163.367
R906 B.n638 B.n637 163.367
R907 B.n637 B.n636 163.367
R908 B.n636 B.n61 163.367
R909 B.n632 B.n61 163.367
R910 B.n632 B.n631 163.367
R911 B.n631 B.n630 163.367
R912 B.n630 B.n63 163.367
R913 B.n626 B.n63 163.367
R914 B.n626 B.n625 163.367
R915 B.n625 B.n624 163.367
R916 B.n624 B.n65 163.367
R917 B.n620 B.n65 163.367
R918 B.n620 B.n619 163.367
R919 B.n619 B.n618 163.367
R920 B.n618 B.n67 163.367
R921 B.n614 B.n67 163.367
R922 B.n614 B.n613 163.367
R923 B.n613 B.n612 163.367
R924 B.n612 B.n69 163.367
R925 B.n608 B.n69 163.367
R926 B.n608 B.n607 163.367
R927 B.n607 B.n606 163.367
R928 B.n606 B.n71 163.367
R929 B.n602 B.n71 163.367
R930 B.n602 B.n601 163.367
R931 B.n601 B.n600 163.367
R932 B.n600 B.n73 163.367
R933 B.n596 B.n73 163.367
R934 B.n596 B.n595 163.367
R935 B.n595 B.n594 163.367
R936 B.n594 B.n75 163.367
R937 B.n590 B.n75 163.367
R938 B.n590 B.n589 163.367
R939 B.n589 B.n588 163.367
R940 B.n588 B.n77 163.367
R941 B.n584 B.n77 163.367
R942 B.n584 B.n583 163.367
R943 B.n583 B.n582 163.367
R944 B.n582 B.n79 163.367
R945 B.n578 B.n79 163.367
R946 B.n578 B.n577 163.367
R947 B.n577 B.n576 163.367
R948 B.n576 B.n81 163.367
R949 B.n572 B.n81 163.367
R950 B.n572 B.n571 163.367
R951 B.n571 B.n570 163.367
R952 B.n570 B.n83 163.367
R953 B.n566 B.n83 163.367
R954 B.n566 B.n565 163.367
R955 B.n565 B.n564 163.367
R956 B.n564 B.n85 163.367
R957 B.n560 B.n85 163.367
R958 B.n560 B.n559 163.367
R959 B.n559 B.n558 163.367
R960 B.n558 B.n87 163.367
R961 B.n554 B.n87 163.367
R962 B.n554 B.n553 163.367
R963 B.n553 B.n552 163.367
R964 B.n152 B.t11 139.064
R965 B.n56 B.t7 139.064
R966 B.n160 B.t2 139.038
R967 B.n50 B.t4 139.038
R968 B.n153 B.t10 109.002
R969 B.n57 B.t8 109.002
R970 B.n161 B.t1 108.978
R971 B.n51 B.t5 108.978
R972 B.n154 B.n153 59.5399
R973 B.n347 B.n161 59.5399
R974 B.n660 B.n51 59.5399
R975 B.n646 B.n57 59.5399
R976 B.n756 B.n755 32.0005
R977 B.n551 B.n550 32.0005
R978 B.n455 B.n120 32.0005
R979 B.n251 B.n192 32.0005
R980 B.n153 B.n152 30.0611
R981 B.n161 B.n160 30.0611
R982 B.n51 B.n50 30.0611
R983 B.n57 B.n56 30.0611
R984 B B.n803 18.0485
R985 B.n755 B.n18 10.6151
R986 B.n751 B.n18 10.6151
R987 B.n751 B.n750 10.6151
R988 B.n750 B.n749 10.6151
R989 B.n749 B.n20 10.6151
R990 B.n745 B.n20 10.6151
R991 B.n745 B.n744 10.6151
R992 B.n744 B.n743 10.6151
R993 B.n743 B.n22 10.6151
R994 B.n739 B.n22 10.6151
R995 B.n739 B.n738 10.6151
R996 B.n738 B.n737 10.6151
R997 B.n737 B.n24 10.6151
R998 B.n733 B.n24 10.6151
R999 B.n733 B.n732 10.6151
R1000 B.n732 B.n731 10.6151
R1001 B.n731 B.n26 10.6151
R1002 B.n727 B.n26 10.6151
R1003 B.n727 B.n726 10.6151
R1004 B.n726 B.n725 10.6151
R1005 B.n725 B.n28 10.6151
R1006 B.n721 B.n28 10.6151
R1007 B.n721 B.n720 10.6151
R1008 B.n720 B.n719 10.6151
R1009 B.n719 B.n30 10.6151
R1010 B.n715 B.n30 10.6151
R1011 B.n715 B.n714 10.6151
R1012 B.n714 B.n713 10.6151
R1013 B.n713 B.n32 10.6151
R1014 B.n709 B.n32 10.6151
R1015 B.n709 B.n708 10.6151
R1016 B.n708 B.n707 10.6151
R1017 B.n707 B.n34 10.6151
R1018 B.n703 B.n34 10.6151
R1019 B.n703 B.n702 10.6151
R1020 B.n702 B.n701 10.6151
R1021 B.n701 B.n36 10.6151
R1022 B.n697 B.n36 10.6151
R1023 B.n697 B.n696 10.6151
R1024 B.n696 B.n695 10.6151
R1025 B.n695 B.n38 10.6151
R1026 B.n691 B.n38 10.6151
R1027 B.n691 B.n690 10.6151
R1028 B.n690 B.n689 10.6151
R1029 B.n689 B.n40 10.6151
R1030 B.n685 B.n40 10.6151
R1031 B.n685 B.n684 10.6151
R1032 B.n684 B.n683 10.6151
R1033 B.n683 B.n42 10.6151
R1034 B.n679 B.n42 10.6151
R1035 B.n679 B.n678 10.6151
R1036 B.n678 B.n677 10.6151
R1037 B.n677 B.n44 10.6151
R1038 B.n673 B.n44 10.6151
R1039 B.n673 B.n672 10.6151
R1040 B.n672 B.n671 10.6151
R1041 B.n671 B.n46 10.6151
R1042 B.n667 B.n46 10.6151
R1043 B.n667 B.n666 10.6151
R1044 B.n666 B.n665 10.6151
R1045 B.n665 B.n48 10.6151
R1046 B.n661 B.n48 10.6151
R1047 B.n659 B.n658 10.6151
R1048 B.n658 B.n52 10.6151
R1049 B.n654 B.n52 10.6151
R1050 B.n654 B.n653 10.6151
R1051 B.n653 B.n652 10.6151
R1052 B.n652 B.n54 10.6151
R1053 B.n648 B.n54 10.6151
R1054 B.n648 B.n647 10.6151
R1055 B.n645 B.n58 10.6151
R1056 B.n641 B.n58 10.6151
R1057 B.n641 B.n640 10.6151
R1058 B.n640 B.n639 10.6151
R1059 B.n639 B.n60 10.6151
R1060 B.n635 B.n60 10.6151
R1061 B.n635 B.n634 10.6151
R1062 B.n634 B.n633 10.6151
R1063 B.n633 B.n62 10.6151
R1064 B.n629 B.n62 10.6151
R1065 B.n629 B.n628 10.6151
R1066 B.n628 B.n627 10.6151
R1067 B.n627 B.n64 10.6151
R1068 B.n623 B.n64 10.6151
R1069 B.n623 B.n622 10.6151
R1070 B.n622 B.n621 10.6151
R1071 B.n621 B.n66 10.6151
R1072 B.n617 B.n66 10.6151
R1073 B.n617 B.n616 10.6151
R1074 B.n616 B.n615 10.6151
R1075 B.n615 B.n68 10.6151
R1076 B.n611 B.n68 10.6151
R1077 B.n611 B.n610 10.6151
R1078 B.n610 B.n609 10.6151
R1079 B.n609 B.n70 10.6151
R1080 B.n605 B.n70 10.6151
R1081 B.n605 B.n604 10.6151
R1082 B.n604 B.n603 10.6151
R1083 B.n603 B.n72 10.6151
R1084 B.n599 B.n72 10.6151
R1085 B.n599 B.n598 10.6151
R1086 B.n598 B.n597 10.6151
R1087 B.n597 B.n74 10.6151
R1088 B.n593 B.n74 10.6151
R1089 B.n593 B.n592 10.6151
R1090 B.n592 B.n591 10.6151
R1091 B.n591 B.n76 10.6151
R1092 B.n587 B.n76 10.6151
R1093 B.n587 B.n586 10.6151
R1094 B.n586 B.n585 10.6151
R1095 B.n585 B.n78 10.6151
R1096 B.n581 B.n78 10.6151
R1097 B.n581 B.n580 10.6151
R1098 B.n580 B.n579 10.6151
R1099 B.n579 B.n80 10.6151
R1100 B.n575 B.n80 10.6151
R1101 B.n575 B.n574 10.6151
R1102 B.n574 B.n573 10.6151
R1103 B.n573 B.n82 10.6151
R1104 B.n569 B.n82 10.6151
R1105 B.n569 B.n568 10.6151
R1106 B.n568 B.n567 10.6151
R1107 B.n567 B.n84 10.6151
R1108 B.n563 B.n84 10.6151
R1109 B.n563 B.n562 10.6151
R1110 B.n562 B.n561 10.6151
R1111 B.n561 B.n86 10.6151
R1112 B.n557 B.n86 10.6151
R1113 B.n557 B.n556 10.6151
R1114 B.n556 B.n555 10.6151
R1115 B.n555 B.n88 10.6151
R1116 B.n551 B.n88 10.6151
R1117 B.n459 B.n120 10.6151
R1118 B.n460 B.n459 10.6151
R1119 B.n461 B.n460 10.6151
R1120 B.n461 B.n118 10.6151
R1121 B.n465 B.n118 10.6151
R1122 B.n466 B.n465 10.6151
R1123 B.n467 B.n466 10.6151
R1124 B.n467 B.n116 10.6151
R1125 B.n471 B.n116 10.6151
R1126 B.n472 B.n471 10.6151
R1127 B.n473 B.n472 10.6151
R1128 B.n473 B.n114 10.6151
R1129 B.n477 B.n114 10.6151
R1130 B.n478 B.n477 10.6151
R1131 B.n479 B.n478 10.6151
R1132 B.n479 B.n112 10.6151
R1133 B.n483 B.n112 10.6151
R1134 B.n484 B.n483 10.6151
R1135 B.n485 B.n484 10.6151
R1136 B.n485 B.n110 10.6151
R1137 B.n489 B.n110 10.6151
R1138 B.n490 B.n489 10.6151
R1139 B.n491 B.n490 10.6151
R1140 B.n491 B.n108 10.6151
R1141 B.n495 B.n108 10.6151
R1142 B.n496 B.n495 10.6151
R1143 B.n497 B.n496 10.6151
R1144 B.n497 B.n106 10.6151
R1145 B.n501 B.n106 10.6151
R1146 B.n502 B.n501 10.6151
R1147 B.n503 B.n502 10.6151
R1148 B.n503 B.n104 10.6151
R1149 B.n507 B.n104 10.6151
R1150 B.n508 B.n507 10.6151
R1151 B.n509 B.n508 10.6151
R1152 B.n509 B.n102 10.6151
R1153 B.n513 B.n102 10.6151
R1154 B.n514 B.n513 10.6151
R1155 B.n515 B.n514 10.6151
R1156 B.n515 B.n100 10.6151
R1157 B.n519 B.n100 10.6151
R1158 B.n520 B.n519 10.6151
R1159 B.n521 B.n520 10.6151
R1160 B.n521 B.n98 10.6151
R1161 B.n525 B.n98 10.6151
R1162 B.n526 B.n525 10.6151
R1163 B.n527 B.n526 10.6151
R1164 B.n527 B.n96 10.6151
R1165 B.n531 B.n96 10.6151
R1166 B.n532 B.n531 10.6151
R1167 B.n533 B.n532 10.6151
R1168 B.n533 B.n94 10.6151
R1169 B.n537 B.n94 10.6151
R1170 B.n538 B.n537 10.6151
R1171 B.n539 B.n538 10.6151
R1172 B.n539 B.n92 10.6151
R1173 B.n543 B.n92 10.6151
R1174 B.n544 B.n543 10.6151
R1175 B.n545 B.n544 10.6151
R1176 B.n545 B.n90 10.6151
R1177 B.n549 B.n90 10.6151
R1178 B.n550 B.n549 10.6151
R1179 B.n255 B.n192 10.6151
R1180 B.n256 B.n255 10.6151
R1181 B.n257 B.n256 10.6151
R1182 B.n257 B.n190 10.6151
R1183 B.n261 B.n190 10.6151
R1184 B.n262 B.n261 10.6151
R1185 B.n263 B.n262 10.6151
R1186 B.n263 B.n188 10.6151
R1187 B.n267 B.n188 10.6151
R1188 B.n268 B.n267 10.6151
R1189 B.n269 B.n268 10.6151
R1190 B.n269 B.n186 10.6151
R1191 B.n273 B.n186 10.6151
R1192 B.n274 B.n273 10.6151
R1193 B.n275 B.n274 10.6151
R1194 B.n275 B.n184 10.6151
R1195 B.n279 B.n184 10.6151
R1196 B.n280 B.n279 10.6151
R1197 B.n281 B.n280 10.6151
R1198 B.n281 B.n182 10.6151
R1199 B.n285 B.n182 10.6151
R1200 B.n286 B.n285 10.6151
R1201 B.n287 B.n286 10.6151
R1202 B.n287 B.n180 10.6151
R1203 B.n291 B.n180 10.6151
R1204 B.n292 B.n291 10.6151
R1205 B.n293 B.n292 10.6151
R1206 B.n293 B.n178 10.6151
R1207 B.n297 B.n178 10.6151
R1208 B.n298 B.n297 10.6151
R1209 B.n299 B.n298 10.6151
R1210 B.n299 B.n176 10.6151
R1211 B.n303 B.n176 10.6151
R1212 B.n304 B.n303 10.6151
R1213 B.n305 B.n304 10.6151
R1214 B.n305 B.n174 10.6151
R1215 B.n309 B.n174 10.6151
R1216 B.n310 B.n309 10.6151
R1217 B.n311 B.n310 10.6151
R1218 B.n311 B.n172 10.6151
R1219 B.n315 B.n172 10.6151
R1220 B.n316 B.n315 10.6151
R1221 B.n317 B.n316 10.6151
R1222 B.n317 B.n170 10.6151
R1223 B.n321 B.n170 10.6151
R1224 B.n322 B.n321 10.6151
R1225 B.n323 B.n322 10.6151
R1226 B.n323 B.n168 10.6151
R1227 B.n327 B.n168 10.6151
R1228 B.n328 B.n327 10.6151
R1229 B.n329 B.n328 10.6151
R1230 B.n329 B.n166 10.6151
R1231 B.n333 B.n166 10.6151
R1232 B.n334 B.n333 10.6151
R1233 B.n335 B.n334 10.6151
R1234 B.n335 B.n164 10.6151
R1235 B.n339 B.n164 10.6151
R1236 B.n340 B.n339 10.6151
R1237 B.n341 B.n340 10.6151
R1238 B.n341 B.n162 10.6151
R1239 B.n345 B.n162 10.6151
R1240 B.n346 B.n345 10.6151
R1241 B.n348 B.n158 10.6151
R1242 B.n352 B.n158 10.6151
R1243 B.n353 B.n352 10.6151
R1244 B.n354 B.n353 10.6151
R1245 B.n354 B.n156 10.6151
R1246 B.n358 B.n156 10.6151
R1247 B.n359 B.n358 10.6151
R1248 B.n360 B.n359 10.6151
R1249 B.n364 B.n363 10.6151
R1250 B.n365 B.n364 10.6151
R1251 B.n365 B.n150 10.6151
R1252 B.n369 B.n150 10.6151
R1253 B.n370 B.n369 10.6151
R1254 B.n371 B.n370 10.6151
R1255 B.n371 B.n148 10.6151
R1256 B.n375 B.n148 10.6151
R1257 B.n376 B.n375 10.6151
R1258 B.n377 B.n376 10.6151
R1259 B.n377 B.n146 10.6151
R1260 B.n381 B.n146 10.6151
R1261 B.n382 B.n381 10.6151
R1262 B.n383 B.n382 10.6151
R1263 B.n383 B.n144 10.6151
R1264 B.n387 B.n144 10.6151
R1265 B.n388 B.n387 10.6151
R1266 B.n389 B.n388 10.6151
R1267 B.n389 B.n142 10.6151
R1268 B.n393 B.n142 10.6151
R1269 B.n394 B.n393 10.6151
R1270 B.n395 B.n394 10.6151
R1271 B.n395 B.n140 10.6151
R1272 B.n399 B.n140 10.6151
R1273 B.n400 B.n399 10.6151
R1274 B.n401 B.n400 10.6151
R1275 B.n401 B.n138 10.6151
R1276 B.n405 B.n138 10.6151
R1277 B.n406 B.n405 10.6151
R1278 B.n407 B.n406 10.6151
R1279 B.n407 B.n136 10.6151
R1280 B.n411 B.n136 10.6151
R1281 B.n412 B.n411 10.6151
R1282 B.n413 B.n412 10.6151
R1283 B.n413 B.n134 10.6151
R1284 B.n417 B.n134 10.6151
R1285 B.n418 B.n417 10.6151
R1286 B.n419 B.n418 10.6151
R1287 B.n419 B.n132 10.6151
R1288 B.n423 B.n132 10.6151
R1289 B.n424 B.n423 10.6151
R1290 B.n425 B.n424 10.6151
R1291 B.n425 B.n130 10.6151
R1292 B.n429 B.n130 10.6151
R1293 B.n430 B.n429 10.6151
R1294 B.n431 B.n430 10.6151
R1295 B.n431 B.n128 10.6151
R1296 B.n435 B.n128 10.6151
R1297 B.n436 B.n435 10.6151
R1298 B.n437 B.n436 10.6151
R1299 B.n437 B.n126 10.6151
R1300 B.n441 B.n126 10.6151
R1301 B.n442 B.n441 10.6151
R1302 B.n443 B.n442 10.6151
R1303 B.n443 B.n124 10.6151
R1304 B.n447 B.n124 10.6151
R1305 B.n448 B.n447 10.6151
R1306 B.n449 B.n448 10.6151
R1307 B.n449 B.n122 10.6151
R1308 B.n453 B.n122 10.6151
R1309 B.n454 B.n453 10.6151
R1310 B.n455 B.n454 10.6151
R1311 B.n251 B.n250 10.6151
R1312 B.n250 B.n249 10.6151
R1313 B.n249 B.n194 10.6151
R1314 B.n245 B.n194 10.6151
R1315 B.n245 B.n244 10.6151
R1316 B.n244 B.n243 10.6151
R1317 B.n243 B.n196 10.6151
R1318 B.n239 B.n196 10.6151
R1319 B.n239 B.n238 10.6151
R1320 B.n238 B.n237 10.6151
R1321 B.n237 B.n198 10.6151
R1322 B.n233 B.n198 10.6151
R1323 B.n233 B.n232 10.6151
R1324 B.n232 B.n231 10.6151
R1325 B.n231 B.n200 10.6151
R1326 B.n227 B.n200 10.6151
R1327 B.n227 B.n226 10.6151
R1328 B.n226 B.n225 10.6151
R1329 B.n225 B.n202 10.6151
R1330 B.n221 B.n202 10.6151
R1331 B.n221 B.n220 10.6151
R1332 B.n220 B.n219 10.6151
R1333 B.n219 B.n204 10.6151
R1334 B.n215 B.n204 10.6151
R1335 B.n215 B.n214 10.6151
R1336 B.n214 B.n213 10.6151
R1337 B.n213 B.n206 10.6151
R1338 B.n209 B.n206 10.6151
R1339 B.n209 B.n208 10.6151
R1340 B.n208 B.n0 10.6151
R1341 B.n799 B.n1 10.6151
R1342 B.n799 B.n798 10.6151
R1343 B.n798 B.n797 10.6151
R1344 B.n797 B.n4 10.6151
R1345 B.n793 B.n4 10.6151
R1346 B.n793 B.n792 10.6151
R1347 B.n792 B.n791 10.6151
R1348 B.n791 B.n6 10.6151
R1349 B.n787 B.n6 10.6151
R1350 B.n787 B.n786 10.6151
R1351 B.n786 B.n785 10.6151
R1352 B.n785 B.n8 10.6151
R1353 B.n781 B.n8 10.6151
R1354 B.n781 B.n780 10.6151
R1355 B.n780 B.n779 10.6151
R1356 B.n779 B.n10 10.6151
R1357 B.n775 B.n10 10.6151
R1358 B.n775 B.n774 10.6151
R1359 B.n774 B.n773 10.6151
R1360 B.n773 B.n12 10.6151
R1361 B.n769 B.n12 10.6151
R1362 B.n769 B.n768 10.6151
R1363 B.n768 B.n767 10.6151
R1364 B.n767 B.n14 10.6151
R1365 B.n763 B.n14 10.6151
R1366 B.n763 B.n762 10.6151
R1367 B.n762 B.n761 10.6151
R1368 B.n761 B.n16 10.6151
R1369 B.n757 B.n16 10.6151
R1370 B.n757 B.n756 10.6151
R1371 B.n660 B.n659 6.5566
R1372 B.n647 B.n646 6.5566
R1373 B.n348 B.n347 6.5566
R1374 B.n360 B.n154 6.5566
R1375 B.n661 B.n660 4.05904
R1376 B.n646 B.n645 4.05904
R1377 B.n347 B.n346 4.05904
R1378 B.n363 B.n154 4.05904
R1379 B.n803 B.n0 2.81026
R1380 B.n803 B.n1 2.81026
C0 w_n2520_n4806# VTAIL 5.87271f
C1 VN VDD1 0.148868f
C2 VN VDD2 11.033299f
C3 VDD1 VDD2 1.08418f
C4 VP B 1.52222f
C5 VP w_n2520_n4806# 5.20658f
C6 VN VTAIL 10.6995f
C7 VDD1 VTAIL 12.731f
C8 VDD2 VTAIL 12.7762f
C9 VN VP 7.306509f
C10 VDD1 VP 11.2561f
C11 VP VDD2 0.372459f
C12 w_n2520_n4806# B 10.0185f
C13 VP VTAIL 10.713599f
C14 VN B 0.98798f
C15 VDD1 B 1.42266f
C16 VN w_n2520_n4806# 4.8835f
C17 VDD2 B 1.47543f
C18 VDD1 w_n2520_n4806# 1.6806f
C19 VDD2 w_n2520_n4806# 1.73729f
C20 VTAIL B 6.3184f
C21 VDD2 VSUBS 1.59886f
C22 VDD1 VSUBS 1.998038f
C23 VTAIL VSUBS 1.39057f
C24 VN VSUBS 5.58698f
C25 VP VSUBS 2.451955f
C26 B VSUBS 4.07226f
C27 w_n2520_n4806# VSUBS 0.147964p
C28 B.n0 VSUBS 0.004446f
C29 B.n1 VSUBS 0.004446f
C30 B.n2 VSUBS 0.007032f
C31 B.n3 VSUBS 0.007032f
C32 B.n4 VSUBS 0.007032f
C33 B.n5 VSUBS 0.007032f
C34 B.n6 VSUBS 0.007032f
C35 B.n7 VSUBS 0.007032f
C36 B.n8 VSUBS 0.007032f
C37 B.n9 VSUBS 0.007032f
C38 B.n10 VSUBS 0.007032f
C39 B.n11 VSUBS 0.007032f
C40 B.n12 VSUBS 0.007032f
C41 B.n13 VSUBS 0.007032f
C42 B.n14 VSUBS 0.007032f
C43 B.n15 VSUBS 0.007032f
C44 B.n16 VSUBS 0.007032f
C45 B.n17 VSUBS 0.015935f
C46 B.n18 VSUBS 0.007032f
C47 B.n19 VSUBS 0.007032f
C48 B.n20 VSUBS 0.007032f
C49 B.n21 VSUBS 0.007032f
C50 B.n22 VSUBS 0.007032f
C51 B.n23 VSUBS 0.007032f
C52 B.n24 VSUBS 0.007032f
C53 B.n25 VSUBS 0.007032f
C54 B.n26 VSUBS 0.007032f
C55 B.n27 VSUBS 0.007032f
C56 B.n28 VSUBS 0.007032f
C57 B.n29 VSUBS 0.007032f
C58 B.n30 VSUBS 0.007032f
C59 B.n31 VSUBS 0.007032f
C60 B.n32 VSUBS 0.007032f
C61 B.n33 VSUBS 0.007032f
C62 B.n34 VSUBS 0.007032f
C63 B.n35 VSUBS 0.007032f
C64 B.n36 VSUBS 0.007032f
C65 B.n37 VSUBS 0.007032f
C66 B.n38 VSUBS 0.007032f
C67 B.n39 VSUBS 0.007032f
C68 B.n40 VSUBS 0.007032f
C69 B.n41 VSUBS 0.007032f
C70 B.n42 VSUBS 0.007032f
C71 B.n43 VSUBS 0.007032f
C72 B.n44 VSUBS 0.007032f
C73 B.n45 VSUBS 0.007032f
C74 B.n46 VSUBS 0.007032f
C75 B.n47 VSUBS 0.007032f
C76 B.n48 VSUBS 0.007032f
C77 B.n49 VSUBS 0.007032f
C78 B.t5 VSUBS 0.653602f
C79 B.t4 VSUBS 0.665863f
C80 B.t3 VSUBS 0.980432f
C81 B.n50 VSUBS 0.263355f
C82 B.n51 VSUBS 0.066737f
C83 B.n52 VSUBS 0.007032f
C84 B.n53 VSUBS 0.007032f
C85 B.n54 VSUBS 0.007032f
C86 B.n55 VSUBS 0.007032f
C87 B.t8 VSUBS 0.653576f
C88 B.t7 VSUBS 0.66584f
C89 B.t6 VSUBS 0.980432f
C90 B.n56 VSUBS 0.263379f
C91 B.n57 VSUBS 0.066764f
C92 B.n58 VSUBS 0.007032f
C93 B.n59 VSUBS 0.007032f
C94 B.n60 VSUBS 0.007032f
C95 B.n61 VSUBS 0.007032f
C96 B.n62 VSUBS 0.007032f
C97 B.n63 VSUBS 0.007032f
C98 B.n64 VSUBS 0.007032f
C99 B.n65 VSUBS 0.007032f
C100 B.n66 VSUBS 0.007032f
C101 B.n67 VSUBS 0.007032f
C102 B.n68 VSUBS 0.007032f
C103 B.n69 VSUBS 0.007032f
C104 B.n70 VSUBS 0.007032f
C105 B.n71 VSUBS 0.007032f
C106 B.n72 VSUBS 0.007032f
C107 B.n73 VSUBS 0.007032f
C108 B.n74 VSUBS 0.007032f
C109 B.n75 VSUBS 0.007032f
C110 B.n76 VSUBS 0.007032f
C111 B.n77 VSUBS 0.007032f
C112 B.n78 VSUBS 0.007032f
C113 B.n79 VSUBS 0.007032f
C114 B.n80 VSUBS 0.007032f
C115 B.n81 VSUBS 0.007032f
C116 B.n82 VSUBS 0.007032f
C117 B.n83 VSUBS 0.007032f
C118 B.n84 VSUBS 0.007032f
C119 B.n85 VSUBS 0.007032f
C120 B.n86 VSUBS 0.007032f
C121 B.n87 VSUBS 0.007032f
C122 B.n88 VSUBS 0.007032f
C123 B.n89 VSUBS 0.015935f
C124 B.n90 VSUBS 0.007032f
C125 B.n91 VSUBS 0.007032f
C126 B.n92 VSUBS 0.007032f
C127 B.n93 VSUBS 0.007032f
C128 B.n94 VSUBS 0.007032f
C129 B.n95 VSUBS 0.007032f
C130 B.n96 VSUBS 0.007032f
C131 B.n97 VSUBS 0.007032f
C132 B.n98 VSUBS 0.007032f
C133 B.n99 VSUBS 0.007032f
C134 B.n100 VSUBS 0.007032f
C135 B.n101 VSUBS 0.007032f
C136 B.n102 VSUBS 0.007032f
C137 B.n103 VSUBS 0.007032f
C138 B.n104 VSUBS 0.007032f
C139 B.n105 VSUBS 0.007032f
C140 B.n106 VSUBS 0.007032f
C141 B.n107 VSUBS 0.007032f
C142 B.n108 VSUBS 0.007032f
C143 B.n109 VSUBS 0.007032f
C144 B.n110 VSUBS 0.007032f
C145 B.n111 VSUBS 0.007032f
C146 B.n112 VSUBS 0.007032f
C147 B.n113 VSUBS 0.007032f
C148 B.n114 VSUBS 0.007032f
C149 B.n115 VSUBS 0.007032f
C150 B.n116 VSUBS 0.007032f
C151 B.n117 VSUBS 0.007032f
C152 B.n118 VSUBS 0.007032f
C153 B.n119 VSUBS 0.007032f
C154 B.n120 VSUBS 0.015935f
C155 B.n121 VSUBS 0.007032f
C156 B.n122 VSUBS 0.007032f
C157 B.n123 VSUBS 0.007032f
C158 B.n124 VSUBS 0.007032f
C159 B.n125 VSUBS 0.007032f
C160 B.n126 VSUBS 0.007032f
C161 B.n127 VSUBS 0.007032f
C162 B.n128 VSUBS 0.007032f
C163 B.n129 VSUBS 0.007032f
C164 B.n130 VSUBS 0.007032f
C165 B.n131 VSUBS 0.007032f
C166 B.n132 VSUBS 0.007032f
C167 B.n133 VSUBS 0.007032f
C168 B.n134 VSUBS 0.007032f
C169 B.n135 VSUBS 0.007032f
C170 B.n136 VSUBS 0.007032f
C171 B.n137 VSUBS 0.007032f
C172 B.n138 VSUBS 0.007032f
C173 B.n139 VSUBS 0.007032f
C174 B.n140 VSUBS 0.007032f
C175 B.n141 VSUBS 0.007032f
C176 B.n142 VSUBS 0.007032f
C177 B.n143 VSUBS 0.007032f
C178 B.n144 VSUBS 0.007032f
C179 B.n145 VSUBS 0.007032f
C180 B.n146 VSUBS 0.007032f
C181 B.n147 VSUBS 0.007032f
C182 B.n148 VSUBS 0.007032f
C183 B.n149 VSUBS 0.007032f
C184 B.n150 VSUBS 0.007032f
C185 B.n151 VSUBS 0.007032f
C186 B.t10 VSUBS 0.653576f
C187 B.t11 VSUBS 0.66584f
C188 B.t9 VSUBS 0.980432f
C189 B.n152 VSUBS 0.263379f
C190 B.n153 VSUBS 0.066764f
C191 B.n154 VSUBS 0.016292f
C192 B.n155 VSUBS 0.007032f
C193 B.n156 VSUBS 0.007032f
C194 B.n157 VSUBS 0.007032f
C195 B.n158 VSUBS 0.007032f
C196 B.n159 VSUBS 0.007032f
C197 B.t1 VSUBS 0.653602f
C198 B.t2 VSUBS 0.665863f
C199 B.t0 VSUBS 0.980432f
C200 B.n160 VSUBS 0.263355f
C201 B.n161 VSUBS 0.066737f
C202 B.n162 VSUBS 0.007032f
C203 B.n163 VSUBS 0.007032f
C204 B.n164 VSUBS 0.007032f
C205 B.n165 VSUBS 0.007032f
C206 B.n166 VSUBS 0.007032f
C207 B.n167 VSUBS 0.007032f
C208 B.n168 VSUBS 0.007032f
C209 B.n169 VSUBS 0.007032f
C210 B.n170 VSUBS 0.007032f
C211 B.n171 VSUBS 0.007032f
C212 B.n172 VSUBS 0.007032f
C213 B.n173 VSUBS 0.007032f
C214 B.n174 VSUBS 0.007032f
C215 B.n175 VSUBS 0.007032f
C216 B.n176 VSUBS 0.007032f
C217 B.n177 VSUBS 0.007032f
C218 B.n178 VSUBS 0.007032f
C219 B.n179 VSUBS 0.007032f
C220 B.n180 VSUBS 0.007032f
C221 B.n181 VSUBS 0.007032f
C222 B.n182 VSUBS 0.007032f
C223 B.n183 VSUBS 0.007032f
C224 B.n184 VSUBS 0.007032f
C225 B.n185 VSUBS 0.007032f
C226 B.n186 VSUBS 0.007032f
C227 B.n187 VSUBS 0.007032f
C228 B.n188 VSUBS 0.007032f
C229 B.n189 VSUBS 0.007032f
C230 B.n190 VSUBS 0.007032f
C231 B.n191 VSUBS 0.007032f
C232 B.n192 VSUBS 0.016535f
C233 B.n193 VSUBS 0.007032f
C234 B.n194 VSUBS 0.007032f
C235 B.n195 VSUBS 0.007032f
C236 B.n196 VSUBS 0.007032f
C237 B.n197 VSUBS 0.007032f
C238 B.n198 VSUBS 0.007032f
C239 B.n199 VSUBS 0.007032f
C240 B.n200 VSUBS 0.007032f
C241 B.n201 VSUBS 0.007032f
C242 B.n202 VSUBS 0.007032f
C243 B.n203 VSUBS 0.007032f
C244 B.n204 VSUBS 0.007032f
C245 B.n205 VSUBS 0.007032f
C246 B.n206 VSUBS 0.007032f
C247 B.n207 VSUBS 0.007032f
C248 B.n208 VSUBS 0.007032f
C249 B.n209 VSUBS 0.007032f
C250 B.n210 VSUBS 0.007032f
C251 B.n211 VSUBS 0.007032f
C252 B.n212 VSUBS 0.007032f
C253 B.n213 VSUBS 0.007032f
C254 B.n214 VSUBS 0.007032f
C255 B.n215 VSUBS 0.007032f
C256 B.n216 VSUBS 0.007032f
C257 B.n217 VSUBS 0.007032f
C258 B.n218 VSUBS 0.007032f
C259 B.n219 VSUBS 0.007032f
C260 B.n220 VSUBS 0.007032f
C261 B.n221 VSUBS 0.007032f
C262 B.n222 VSUBS 0.007032f
C263 B.n223 VSUBS 0.007032f
C264 B.n224 VSUBS 0.007032f
C265 B.n225 VSUBS 0.007032f
C266 B.n226 VSUBS 0.007032f
C267 B.n227 VSUBS 0.007032f
C268 B.n228 VSUBS 0.007032f
C269 B.n229 VSUBS 0.007032f
C270 B.n230 VSUBS 0.007032f
C271 B.n231 VSUBS 0.007032f
C272 B.n232 VSUBS 0.007032f
C273 B.n233 VSUBS 0.007032f
C274 B.n234 VSUBS 0.007032f
C275 B.n235 VSUBS 0.007032f
C276 B.n236 VSUBS 0.007032f
C277 B.n237 VSUBS 0.007032f
C278 B.n238 VSUBS 0.007032f
C279 B.n239 VSUBS 0.007032f
C280 B.n240 VSUBS 0.007032f
C281 B.n241 VSUBS 0.007032f
C282 B.n242 VSUBS 0.007032f
C283 B.n243 VSUBS 0.007032f
C284 B.n244 VSUBS 0.007032f
C285 B.n245 VSUBS 0.007032f
C286 B.n246 VSUBS 0.007032f
C287 B.n247 VSUBS 0.007032f
C288 B.n248 VSUBS 0.007032f
C289 B.n249 VSUBS 0.007032f
C290 B.n250 VSUBS 0.007032f
C291 B.n251 VSUBS 0.015935f
C292 B.n252 VSUBS 0.015935f
C293 B.n253 VSUBS 0.016535f
C294 B.n254 VSUBS 0.007032f
C295 B.n255 VSUBS 0.007032f
C296 B.n256 VSUBS 0.007032f
C297 B.n257 VSUBS 0.007032f
C298 B.n258 VSUBS 0.007032f
C299 B.n259 VSUBS 0.007032f
C300 B.n260 VSUBS 0.007032f
C301 B.n261 VSUBS 0.007032f
C302 B.n262 VSUBS 0.007032f
C303 B.n263 VSUBS 0.007032f
C304 B.n264 VSUBS 0.007032f
C305 B.n265 VSUBS 0.007032f
C306 B.n266 VSUBS 0.007032f
C307 B.n267 VSUBS 0.007032f
C308 B.n268 VSUBS 0.007032f
C309 B.n269 VSUBS 0.007032f
C310 B.n270 VSUBS 0.007032f
C311 B.n271 VSUBS 0.007032f
C312 B.n272 VSUBS 0.007032f
C313 B.n273 VSUBS 0.007032f
C314 B.n274 VSUBS 0.007032f
C315 B.n275 VSUBS 0.007032f
C316 B.n276 VSUBS 0.007032f
C317 B.n277 VSUBS 0.007032f
C318 B.n278 VSUBS 0.007032f
C319 B.n279 VSUBS 0.007032f
C320 B.n280 VSUBS 0.007032f
C321 B.n281 VSUBS 0.007032f
C322 B.n282 VSUBS 0.007032f
C323 B.n283 VSUBS 0.007032f
C324 B.n284 VSUBS 0.007032f
C325 B.n285 VSUBS 0.007032f
C326 B.n286 VSUBS 0.007032f
C327 B.n287 VSUBS 0.007032f
C328 B.n288 VSUBS 0.007032f
C329 B.n289 VSUBS 0.007032f
C330 B.n290 VSUBS 0.007032f
C331 B.n291 VSUBS 0.007032f
C332 B.n292 VSUBS 0.007032f
C333 B.n293 VSUBS 0.007032f
C334 B.n294 VSUBS 0.007032f
C335 B.n295 VSUBS 0.007032f
C336 B.n296 VSUBS 0.007032f
C337 B.n297 VSUBS 0.007032f
C338 B.n298 VSUBS 0.007032f
C339 B.n299 VSUBS 0.007032f
C340 B.n300 VSUBS 0.007032f
C341 B.n301 VSUBS 0.007032f
C342 B.n302 VSUBS 0.007032f
C343 B.n303 VSUBS 0.007032f
C344 B.n304 VSUBS 0.007032f
C345 B.n305 VSUBS 0.007032f
C346 B.n306 VSUBS 0.007032f
C347 B.n307 VSUBS 0.007032f
C348 B.n308 VSUBS 0.007032f
C349 B.n309 VSUBS 0.007032f
C350 B.n310 VSUBS 0.007032f
C351 B.n311 VSUBS 0.007032f
C352 B.n312 VSUBS 0.007032f
C353 B.n313 VSUBS 0.007032f
C354 B.n314 VSUBS 0.007032f
C355 B.n315 VSUBS 0.007032f
C356 B.n316 VSUBS 0.007032f
C357 B.n317 VSUBS 0.007032f
C358 B.n318 VSUBS 0.007032f
C359 B.n319 VSUBS 0.007032f
C360 B.n320 VSUBS 0.007032f
C361 B.n321 VSUBS 0.007032f
C362 B.n322 VSUBS 0.007032f
C363 B.n323 VSUBS 0.007032f
C364 B.n324 VSUBS 0.007032f
C365 B.n325 VSUBS 0.007032f
C366 B.n326 VSUBS 0.007032f
C367 B.n327 VSUBS 0.007032f
C368 B.n328 VSUBS 0.007032f
C369 B.n329 VSUBS 0.007032f
C370 B.n330 VSUBS 0.007032f
C371 B.n331 VSUBS 0.007032f
C372 B.n332 VSUBS 0.007032f
C373 B.n333 VSUBS 0.007032f
C374 B.n334 VSUBS 0.007032f
C375 B.n335 VSUBS 0.007032f
C376 B.n336 VSUBS 0.007032f
C377 B.n337 VSUBS 0.007032f
C378 B.n338 VSUBS 0.007032f
C379 B.n339 VSUBS 0.007032f
C380 B.n340 VSUBS 0.007032f
C381 B.n341 VSUBS 0.007032f
C382 B.n342 VSUBS 0.007032f
C383 B.n343 VSUBS 0.007032f
C384 B.n344 VSUBS 0.007032f
C385 B.n345 VSUBS 0.007032f
C386 B.n346 VSUBS 0.00486f
C387 B.n347 VSUBS 0.016292f
C388 B.n348 VSUBS 0.005687f
C389 B.n349 VSUBS 0.007032f
C390 B.n350 VSUBS 0.007032f
C391 B.n351 VSUBS 0.007032f
C392 B.n352 VSUBS 0.007032f
C393 B.n353 VSUBS 0.007032f
C394 B.n354 VSUBS 0.007032f
C395 B.n355 VSUBS 0.007032f
C396 B.n356 VSUBS 0.007032f
C397 B.n357 VSUBS 0.007032f
C398 B.n358 VSUBS 0.007032f
C399 B.n359 VSUBS 0.007032f
C400 B.n360 VSUBS 0.005687f
C401 B.n361 VSUBS 0.007032f
C402 B.n362 VSUBS 0.007032f
C403 B.n363 VSUBS 0.00486f
C404 B.n364 VSUBS 0.007032f
C405 B.n365 VSUBS 0.007032f
C406 B.n366 VSUBS 0.007032f
C407 B.n367 VSUBS 0.007032f
C408 B.n368 VSUBS 0.007032f
C409 B.n369 VSUBS 0.007032f
C410 B.n370 VSUBS 0.007032f
C411 B.n371 VSUBS 0.007032f
C412 B.n372 VSUBS 0.007032f
C413 B.n373 VSUBS 0.007032f
C414 B.n374 VSUBS 0.007032f
C415 B.n375 VSUBS 0.007032f
C416 B.n376 VSUBS 0.007032f
C417 B.n377 VSUBS 0.007032f
C418 B.n378 VSUBS 0.007032f
C419 B.n379 VSUBS 0.007032f
C420 B.n380 VSUBS 0.007032f
C421 B.n381 VSUBS 0.007032f
C422 B.n382 VSUBS 0.007032f
C423 B.n383 VSUBS 0.007032f
C424 B.n384 VSUBS 0.007032f
C425 B.n385 VSUBS 0.007032f
C426 B.n386 VSUBS 0.007032f
C427 B.n387 VSUBS 0.007032f
C428 B.n388 VSUBS 0.007032f
C429 B.n389 VSUBS 0.007032f
C430 B.n390 VSUBS 0.007032f
C431 B.n391 VSUBS 0.007032f
C432 B.n392 VSUBS 0.007032f
C433 B.n393 VSUBS 0.007032f
C434 B.n394 VSUBS 0.007032f
C435 B.n395 VSUBS 0.007032f
C436 B.n396 VSUBS 0.007032f
C437 B.n397 VSUBS 0.007032f
C438 B.n398 VSUBS 0.007032f
C439 B.n399 VSUBS 0.007032f
C440 B.n400 VSUBS 0.007032f
C441 B.n401 VSUBS 0.007032f
C442 B.n402 VSUBS 0.007032f
C443 B.n403 VSUBS 0.007032f
C444 B.n404 VSUBS 0.007032f
C445 B.n405 VSUBS 0.007032f
C446 B.n406 VSUBS 0.007032f
C447 B.n407 VSUBS 0.007032f
C448 B.n408 VSUBS 0.007032f
C449 B.n409 VSUBS 0.007032f
C450 B.n410 VSUBS 0.007032f
C451 B.n411 VSUBS 0.007032f
C452 B.n412 VSUBS 0.007032f
C453 B.n413 VSUBS 0.007032f
C454 B.n414 VSUBS 0.007032f
C455 B.n415 VSUBS 0.007032f
C456 B.n416 VSUBS 0.007032f
C457 B.n417 VSUBS 0.007032f
C458 B.n418 VSUBS 0.007032f
C459 B.n419 VSUBS 0.007032f
C460 B.n420 VSUBS 0.007032f
C461 B.n421 VSUBS 0.007032f
C462 B.n422 VSUBS 0.007032f
C463 B.n423 VSUBS 0.007032f
C464 B.n424 VSUBS 0.007032f
C465 B.n425 VSUBS 0.007032f
C466 B.n426 VSUBS 0.007032f
C467 B.n427 VSUBS 0.007032f
C468 B.n428 VSUBS 0.007032f
C469 B.n429 VSUBS 0.007032f
C470 B.n430 VSUBS 0.007032f
C471 B.n431 VSUBS 0.007032f
C472 B.n432 VSUBS 0.007032f
C473 B.n433 VSUBS 0.007032f
C474 B.n434 VSUBS 0.007032f
C475 B.n435 VSUBS 0.007032f
C476 B.n436 VSUBS 0.007032f
C477 B.n437 VSUBS 0.007032f
C478 B.n438 VSUBS 0.007032f
C479 B.n439 VSUBS 0.007032f
C480 B.n440 VSUBS 0.007032f
C481 B.n441 VSUBS 0.007032f
C482 B.n442 VSUBS 0.007032f
C483 B.n443 VSUBS 0.007032f
C484 B.n444 VSUBS 0.007032f
C485 B.n445 VSUBS 0.007032f
C486 B.n446 VSUBS 0.007032f
C487 B.n447 VSUBS 0.007032f
C488 B.n448 VSUBS 0.007032f
C489 B.n449 VSUBS 0.007032f
C490 B.n450 VSUBS 0.007032f
C491 B.n451 VSUBS 0.007032f
C492 B.n452 VSUBS 0.007032f
C493 B.n453 VSUBS 0.007032f
C494 B.n454 VSUBS 0.007032f
C495 B.n455 VSUBS 0.016535f
C496 B.n456 VSUBS 0.016535f
C497 B.n457 VSUBS 0.015935f
C498 B.n458 VSUBS 0.007032f
C499 B.n459 VSUBS 0.007032f
C500 B.n460 VSUBS 0.007032f
C501 B.n461 VSUBS 0.007032f
C502 B.n462 VSUBS 0.007032f
C503 B.n463 VSUBS 0.007032f
C504 B.n464 VSUBS 0.007032f
C505 B.n465 VSUBS 0.007032f
C506 B.n466 VSUBS 0.007032f
C507 B.n467 VSUBS 0.007032f
C508 B.n468 VSUBS 0.007032f
C509 B.n469 VSUBS 0.007032f
C510 B.n470 VSUBS 0.007032f
C511 B.n471 VSUBS 0.007032f
C512 B.n472 VSUBS 0.007032f
C513 B.n473 VSUBS 0.007032f
C514 B.n474 VSUBS 0.007032f
C515 B.n475 VSUBS 0.007032f
C516 B.n476 VSUBS 0.007032f
C517 B.n477 VSUBS 0.007032f
C518 B.n478 VSUBS 0.007032f
C519 B.n479 VSUBS 0.007032f
C520 B.n480 VSUBS 0.007032f
C521 B.n481 VSUBS 0.007032f
C522 B.n482 VSUBS 0.007032f
C523 B.n483 VSUBS 0.007032f
C524 B.n484 VSUBS 0.007032f
C525 B.n485 VSUBS 0.007032f
C526 B.n486 VSUBS 0.007032f
C527 B.n487 VSUBS 0.007032f
C528 B.n488 VSUBS 0.007032f
C529 B.n489 VSUBS 0.007032f
C530 B.n490 VSUBS 0.007032f
C531 B.n491 VSUBS 0.007032f
C532 B.n492 VSUBS 0.007032f
C533 B.n493 VSUBS 0.007032f
C534 B.n494 VSUBS 0.007032f
C535 B.n495 VSUBS 0.007032f
C536 B.n496 VSUBS 0.007032f
C537 B.n497 VSUBS 0.007032f
C538 B.n498 VSUBS 0.007032f
C539 B.n499 VSUBS 0.007032f
C540 B.n500 VSUBS 0.007032f
C541 B.n501 VSUBS 0.007032f
C542 B.n502 VSUBS 0.007032f
C543 B.n503 VSUBS 0.007032f
C544 B.n504 VSUBS 0.007032f
C545 B.n505 VSUBS 0.007032f
C546 B.n506 VSUBS 0.007032f
C547 B.n507 VSUBS 0.007032f
C548 B.n508 VSUBS 0.007032f
C549 B.n509 VSUBS 0.007032f
C550 B.n510 VSUBS 0.007032f
C551 B.n511 VSUBS 0.007032f
C552 B.n512 VSUBS 0.007032f
C553 B.n513 VSUBS 0.007032f
C554 B.n514 VSUBS 0.007032f
C555 B.n515 VSUBS 0.007032f
C556 B.n516 VSUBS 0.007032f
C557 B.n517 VSUBS 0.007032f
C558 B.n518 VSUBS 0.007032f
C559 B.n519 VSUBS 0.007032f
C560 B.n520 VSUBS 0.007032f
C561 B.n521 VSUBS 0.007032f
C562 B.n522 VSUBS 0.007032f
C563 B.n523 VSUBS 0.007032f
C564 B.n524 VSUBS 0.007032f
C565 B.n525 VSUBS 0.007032f
C566 B.n526 VSUBS 0.007032f
C567 B.n527 VSUBS 0.007032f
C568 B.n528 VSUBS 0.007032f
C569 B.n529 VSUBS 0.007032f
C570 B.n530 VSUBS 0.007032f
C571 B.n531 VSUBS 0.007032f
C572 B.n532 VSUBS 0.007032f
C573 B.n533 VSUBS 0.007032f
C574 B.n534 VSUBS 0.007032f
C575 B.n535 VSUBS 0.007032f
C576 B.n536 VSUBS 0.007032f
C577 B.n537 VSUBS 0.007032f
C578 B.n538 VSUBS 0.007032f
C579 B.n539 VSUBS 0.007032f
C580 B.n540 VSUBS 0.007032f
C581 B.n541 VSUBS 0.007032f
C582 B.n542 VSUBS 0.007032f
C583 B.n543 VSUBS 0.007032f
C584 B.n544 VSUBS 0.007032f
C585 B.n545 VSUBS 0.007032f
C586 B.n546 VSUBS 0.007032f
C587 B.n547 VSUBS 0.007032f
C588 B.n548 VSUBS 0.007032f
C589 B.n549 VSUBS 0.007032f
C590 B.n550 VSUBS 0.016783f
C591 B.n551 VSUBS 0.015687f
C592 B.n552 VSUBS 0.016535f
C593 B.n553 VSUBS 0.007032f
C594 B.n554 VSUBS 0.007032f
C595 B.n555 VSUBS 0.007032f
C596 B.n556 VSUBS 0.007032f
C597 B.n557 VSUBS 0.007032f
C598 B.n558 VSUBS 0.007032f
C599 B.n559 VSUBS 0.007032f
C600 B.n560 VSUBS 0.007032f
C601 B.n561 VSUBS 0.007032f
C602 B.n562 VSUBS 0.007032f
C603 B.n563 VSUBS 0.007032f
C604 B.n564 VSUBS 0.007032f
C605 B.n565 VSUBS 0.007032f
C606 B.n566 VSUBS 0.007032f
C607 B.n567 VSUBS 0.007032f
C608 B.n568 VSUBS 0.007032f
C609 B.n569 VSUBS 0.007032f
C610 B.n570 VSUBS 0.007032f
C611 B.n571 VSUBS 0.007032f
C612 B.n572 VSUBS 0.007032f
C613 B.n573 VSUBS 0.007032f
C614 B.n574 VSUBS 0.007032f
C615 B.n575 VSUBS 0.007032f
C616 B.n576 VSUBS 0.007032f
C617 B.n577 VSUBS 0.007032f
C618 B.n578 VSUBS 0.007032f
C619 B.n579 VSUBS 0.007032f
C620 B.n580 VSUBS 0.007032f
C621 B.n581 VSUBS 0.007032f
C622 B.n582 VSUBS 0.007032f
C623 B.n583 VSUBS 0.007032f
C624 B.n584 VSUBS 0.007032f
C625 B.n585 VSUBS 0.007032f
C626 B.n586 VSUBS 0.007032f
C627 B.n587 VSUBS 0.007032f
C628 B.n588 VSUBS 0.007032f
C629 B.n589 VSUBS 0.007032f
C630 B.n590 VSUBS 0.007032f
C631 B.n591 VSUBS 0.007032f
C632 B.n592 VSUBS 0.007032f
C633 B.n593 VSUBS 0.007032f
C634 B.n594 VSUBS 0.007032f
C635 B.n595 VSUBS 0.007032f
C636 B.n596 VSUBS 0.007032f
C637 B.n597 VSUBS 0.007032f
C638 B.n598 VSUBS 0.007032f
C639 B.n599 VSUBS 0.007032f
C640 B.n600 VSUBS 0.007032f
C641 B.n601 VSUBS 0.007032f
C642 B.n602 VSUBS 0.007032f
C643 B.n603 VSUBS 0.007032f
C644 B.n604 VSUBS 0.007032f
C645 B.n605 VSUBS 0.007032f
C646 B.n606 VSUBS 0.007032f
C647 B.n607 VSUBS 0.007032f
C648 B.n608 VSUBS 0.007032f
C649 B.n609 VSUBS 0.007032f
C650 B.n610 VSUBS 0.007032f
C651 B.n611 VSUBS 0.007032f
C652 B.n612 VSUBS 0.007032f
C653 B.n613 VSUBS 0.007032f
C654 B.n614 VSUBS 0.007032f
C655 B.n615 VSUBS 0.007032f
C656 B.n616 VSUBS 0.007032f
C657 B.n617 VSUBS 0.007032f
C658 B.n618 VSUBS 0.007032f
C659 B.n619 VSUBS 0.007032f
C660 B.n620 VSUBS 0.007032f
C661 B.n621 VSUBS 0.007032f
C662 B.n622 VSUBS 0.007032f
C663 B.n623 VSUBS 0.007032f
C664 B.n624 VSUBS 0.007032f
C665 B.n625 VSUBS 0.007032f
C666 B.n626 VSUBS 0.007032f
C667 B.n627 VSUBS 0.007032f
C668 B.n628 VSUBS 0.007032f
C669 B.n629 VSUBS 0.007032f
C670 B.n630 VSUBS 0.007032f
C671 B.n631 VSUBS 0.007032f
C672 B.n632 VSUBS 0.007032f
C673 B.n633 VSUBS 0.007032f
C674 B.n634 VSUBS 0.007032f
C675 B.n635 VSUBS 0.007032f
C676 B.n636 VSUBS 0.007032f
C677 B.n637 VSUBS 0.007032f
C678 B.n638 VSUBS 0.007032f
C679 B.n639 VSUBS 0.007032f
C680 B.n640 VSUBS 0.007032f
C681 B.n641 VSUBS 0.007032f
C682 B.n642 VSUBS 0.007032f
C683 B.n643 VSUBS 0.007032f
C684 B.n644 VSUBS 0.007032f
C685 B.n645 VSUBS 0.00486f
C686 B.n646 VSUBS 0.016292f
C687 B.n647 VSUBS 0.005687f
C688 B.n648 VSUBS 0.007032f
C689 B.n649 VSUBS 0.007032f
C690 B.n650 VSUBS 0.007032f
C691 B.n651 VSUBS 0.007032f
C692 B.n652 VSUBS 0.007032f
C693 B.n653 VSUBS 0.007032f
C694 B.n654 VSUBS 0.007032f
C695 B.n655 VSUBS 0.007032f
C696 B.n656 VSUBS 0.007032f
C697 B.n657 VSUBS 0.007032f
C698 B.n658 VSUBS 0.007032f
C699 B.n659 VSUBS 0.005687f
C700 B.n660 VSUBS 0.016292f
C701 B.n661 VSUBS 0.00486f
C702 B.n662 VSUBS 0.007032f
C703 B.n663 VSUBS 0.007032f
C704 B.n664 VSUBS 0.007032f
C705 B.n665 VSUBS 0.007032f
C706 B.n666 VSUBS 0.007032f
C707 B.n667 VSUBS 0.007032f
C708 B.n668 VSUBS 0.007032f
C709 B.n669 VSUBS 0.007032f
C710 B.n670 VSUBS 0.007032f
C711 B.n671 VSUBS 0.007032f
C712 B.n672 VSUBS 0.007032f
C713 B.n673 VSUBS 0.007032f
C714 B.n674 VSUBS 0.007032f
C715 B.n675 VSUBS 0.007032f
C716 B.n676 VSUBS 0.007032f
C717 B.n677 VSUBS 0.007032f
C718 B.n678 VSUBS 0.007032f
C719 B.n679 VSUBS 0.007032f
C720 B.n680 VSUBS 0.007032f
C721 B.n681 VSUBS 0.007032f
C722 B.n682 VSUBS 0.007032f
C723 B.n683 VSUBS 0.007032f
C724 B.n684 VSUBS 0.007032f
C725 B.n685 VSUBS 0.007032f
C726 B.n686 VSUBS 0.007032f
C727 B.n687 VSUBS 0.007032f
C728 B.n688 VSUBS 0.007032f
C729 B.n689 VSUBS 0.007032f
C730 B.n690 VSUBS 0.007032f
C731 B.n691 VSUBS 0.007032f
C732 B.n692 VSUBS 0.007032f
C733 B.n693 VSUBS 0.007032f
C734 B.n694 VSUBS 0.007032f
C735 B.n695 VSUBS 0.007032f
C736 B.n696 VSUBS 0.007032f
C737 B.n697 VSUBS 0.007032f
C738 B.n698 VSUBS 0.007032f
C739 B.n699 VSUBS 0.007032f
C740 B.n700 VSUBS 0.007032f
C741 B.n701 VSUBS 0.007032f
C742 B.n702 VSUBS 0.007032f
C743 B.n703 VSUBS 0.007032f
C744 B.n704 VSUBS 0.007032f
C745 B.n705 VSUBS 0.007032f
C746 B.n706 VSUBS 0.007032f
C747 B.n707 VSUBS 0.007032f
C748 B.n708 VSUBS 0.007032f
C749 B.n709 VSUBS 0.007032f
C750 B.n710 VSUBS 0.007032f
C751 B.n711 VSUBS 0.007032f
C752 B.n712 VSUBS 0.007032f
C753 B.n713 VSUBS 0.007032f
C754 B.n714 VSUBS 0.007032f
C755 B.n715 VSUBS 0.007032f
C756 B.n716 VSUBS 0.007032f
C757 B.n717 VSUBS 0.007032f
C758 B.n718 VSUBS 0.007032f
C759 B.n719 VSUBS 0.007032f
C760 B.n720 VSUBS 0.007032f
C761 B.n721 VSUBS 0.007032f
C762 B.n722 VSUBS 0.007032f
C763 B.n723 VSUBS 0.007032f
C764 B.n724 VSUBS 0.007032f
C765 B.n725 VSUBS 0.007032f
C766 B.n726 VSUBS 0.007032f
C767 B.n727 VSUBS 0.007032f
C768 B.n728 VSUBS 0.007032f
C769 B.n729 VSUBS 0.007032f
C770 B.n730 VSUBS 0.007032f
C771 B.n731 VSUBS 0.007032f
C772 B.n732 VSUBS 0.007032f
C773 B.n733 VSUBS 0.007032f
C774 B.n734 VSUBS 0.007032f
C775 B.n735 VSUBS 0.007032f
C776 B.n736 VSUBS 0.007032f
C777 B.n737 VSUBS 0.007032f
C778 B.n738 VSUBS 0.007032f
C779 B.n739 VSUBS 0.007032f
C780 B.n740 VSUBS 0.007032f
C781 B.n741 VSUBS 0.007032f
C782 B.n742 VSUBS 0.007032f
C783 B.n743 VSUBS 0.007032f
C784 B.n744 VSUBS 0.007032f
C785 B.n745 VSUBS 0.007032f
C786 B.n746 VSUBS 0.007032f
C787 B.n747 VSUBS 0.007032f
C788 B.n748 VSUBS 0.007032f
C789 B.n749 VSUBS 0.007032f
C790 B.n750 VSUBS 0.007032f
C791 B.n751 VSUBS 0.007032f
C792 B.n752 VSUBS 0.007032f
C793 B.n753 VSUBS 0.007032f
C794 B.n754 VSUBS 0.016535f
C795 B.n755 VSUBS 0.016535f
C796 B.n756 VSUBS 0.015935f
C797 B.n757 VSUBS 0.007032f
C798 B.n758 VSUBS 0.007032f
C799 B.n759 VSUBS 0.007032f
C800 B.n760 VSUBS 0.007032f
C801 B.n761 VSUBS 0.007032f
C802 B.n762 VSUBS 0.007032f
C803 B.n763 VSUBS 0.007032f
C804 B.n764 VSUBS 0.007032f
C805 B.n765 VSUBS 0.007032f
C806 B.n766 VSUBS 0.007032f
C807 B.n767 VSUBS 0.007032f
C808 B.n768 VSUBS 0.007032f
C809 B.n769 VSUBS 0.007032f
C810 B.n770 VSUBS 0.007032f
C811 B.n771 VSUBS 0.007032f
C812 B.n772 VSUBS 0.007032f
C813 B.n773 VSUBS 0.007032f
C814 B.n774 VSUBS 0.007032f
C815 B.n775 VSUBS 0.007032f
C816 B.n776 VSUBS 0.007032f
C817 B.n777 VSUBS 0.007032f
C818 B.n778 VSUBS 0.007032f
C819 B.n779 VSUBS 0.007032f
C820 B.n780 VSUBS 0.007032f
C821 B.n781 VSUBS 0.007032f
C822 B.n782 VSUBS 0.007032f
C823 B.n783 VSUBS 0.007032f
C824 B.n784 VSUBS 0.007032f
C825 B.n785 VSUBS 0.007032f
C826 B.n786 VSUBS 0.007032f
C827 B.n787 VSUBS 0.007032f
C828 B.n788 VSUBS 0.007032f
C829 B.n789 VSUBS 0.007032f
C830 B.n790 VSUBS 0.007032f
C831 B.n791 VSUBS 0.007032f
C832 B.n792 VSUBS 0.007032f
C833 B.n793 VSUBS 0.007032f
C834 B.n794 VSUBS 0.007032f
C835 B.n795 VSUBS 0.007032f
C836 B.n796 VSUBS 0.007032f
C837 B.n797 VSUBS 0.007032f
C838 B.n798 VSUBS 0.007032f
C839 B.n799 VSUBS 0.007032f
C840 B.n800 VSUBS 0.007032f
C841 B.n801 VSUBS 0.007032f
C842 B.n802 VSUBS 0.007032f
C843 B.n803 VSUBS 0.015922f
C844 VDD1.t2 VSUBS 0.388527f
C845 VDD1.t6 VSUBS 0.388527f
C846 VDD1.n0 VSUBS 3.28632f
C847 VDD1.t1 VSUBS 0.388527f
C848 VDD1.t5 VSUBS 0.388527f
C849 VDD1.n1 VSUBS 3.28521f
C850 VDD1.t0 VSUBS 0.388527f
C851 VDD1.t3 VSUBS 0.388527f
C852 VDD1.n2 VSUBS 3.28521f
C853 VDD1.n3 VSUBS 3.59199f
C854 VDD1.t4 VSUBS 0.388527f
C855 VDD1.t7 VSUBS 0.388527f
C856 VDD1.n4 VSUBS 3.27971f
C857 VDD1.n5 VSUBS 3.39665f
C858 VP.n0 VSUBS 0.053594f
C859 VP.t7 VSUBS 2.58942f
C860 VP.n1 VSUBS 0.915351f
C861 VP.n2 VSUBS 0.040164f
C862 VP.t2 VSUBS 2.58942f
C863 VP.n3 VSUBS 0.915351f
C864 VP.n4 VSUBS 0.053594f
C865 VP.n5 VSUBS 0.053594f
C866 VP.t0 VSUBS 2.66449f
C867 VP.t3 VSUBS 2.58942f
C868 VP.n6 VSUBS 0.915351f
C869 VP.n7 VSUBS 0.040164f
C870 VP.t1 VSUBS 2.58942f
C871 VP.n8 VSUBS 0.967571f
C872 VP.t5 VSUBS 2.70892f
C873 VP.n9 VSUBS 0.982539f
C874 VP.n10 VSUBS 0.208118f
C875 VP.n11 VSUBS 0.063193f
C876 VP.n12 VSUBS 0.032469f
C877 VP.n13 VSUBS 0.063193f
C878 VP.n14 VSUBS 0.040164f
C879 VP.n15 VSUBS 0.040164f
C880 VP.n16 VSUBS 0.06078f
C881 VP.n17 VSUBS 0.025662f
C882 VP.n18 VSUBS 0.990886f
C883 VP.n19 VSUBS 2.19947f
C884 VP.n20 VSUBS 2.22833f
C885 VP.t6 VSUBS 2.66449f
C886 VP.n21 VSUBS 0.990886f
C887 VP.n22 VSUBS 0.025662f
C888 VP.n23 VSUBS 0.06078f
C889 VP.n24 VSUBS 0.040164f
C890 VP.n25 VSUBS 0.040164f
C891 VP.n26 VSUBS 0.063193f
C892 VP.n27 VSUBS 0.032469f
C893 VP.n28 VSUBS 0.063193f
C894 VP.n29 VSUBS 0.040164f
C895 VP.n30 VSUBS 0.040164f
C896 VP.n31 VSUBS 0.06078f
C897 VP.n32 VSUBS 0.025662f
C898 VP.t4 VSUBS 2.66449f
C899 VP.n33 VSUBS 0.990886f
C900 VP.n34 VSUBS 0.037615f
C901 VDD2.t4 VSUBS 0.386815f
C902 VDD2.t0 VSUBS 0.386815f
C903 VDD2.n0 VSUBS 3.27073f
C904 VDD2.t1 VSUBS 0.386815f
C905 VDD2.t7 VSUBS 0.386815f
C906 VDD2.n1 VSUBS 3.27073f
C907 VDD2.n2 VSUBS 3.52253f
C908 VDD2.t6 VSUBS 0.386815f
C909 VDD2.t5 VSUBS 0.386815f
C910 VDD2.n3 VSUBS 3.26528f
C911 VDD2.n4 VSUBS 3.35064f
C912 VDD2.t3 VSUBS 0.386815f
C913 VDD2.t2 VSUBS 0.386815f
C914 VDD2.n5 VSUBS 3.27069f
C915 VTAIL.t11 VSUBS 0.35041f
C916 VTAIL.t10 VSUBS 0.35041f
C917 VTAIL.n0 VSUBS 2.82912f
C918 VTAIL.n1 VSUBS 0.636295f
C919 VTAIL.t13 VSUBS 3.68351f
C920 VTAIL.n2 VSUBS 0.768224f
C921 VTAIL.t5 VSUBS 3.68351f
C922 VTAIL.n3 VSUBS 0.768224f
C923 VTAIL.t3 VSUBS 0.35041f
C924 VTAIL.t2 VSUBS 0.35041f
C925 VTAIL.n4 VSUBS 2.82912f
C926 VTAIL.n5 VSUBS 0.731452f
C927 VTAIL.t4 VSUBS 3.68351f
C928 VTAIL.n6 VSUBS 2.37836f
C929 VTAIL.t9 VSUBS 3.68354f
C930 VTAIL.n7 VSUBS 2.37833f
C931 VTAIL.t8 VSUBS 0.35041f
C932 VTAIL.t12 VSUBS 0.35041f
C933 VTAIL.n8 VSUBS 2.82914f
C934 VTAIL.n9 VSUBS 0.731436f
C935 VTAIL.t14 VSUBS 3.68354f
C936 VTAIL.n10 VSUBS 0.768191f
C937 VTAIL.t0 VSUBS 3.68354f
C938 VTAIL.n11 VSUBS 0.768191f
C939 VTAIL.t6 VSUBS 0.35041f
C940 VTAIL.t1 VSUBS 0.35041f
C941 VTAIL.n12 VSUBS 2.82914f
C942 VTAIL.n13 VSUBS 0.731436f
C943 VTAIL.t7 VSUBS 3.68351f
C944 VTAIL.n14 VSUBS 2.37836f
C945 VTAIL.t15 VSUBS 3.68351f
C946 VTAIL.n15 VSUBS 2.37403f
C947 VN.n0 VSUBS 0.052576f
C948 VN.t6 VSUBS 2.54023f
C949 VN.n1 VSUBS 0.897962f
C950 VN.n2 VSUBS 0.039401f
C951 VN.t7 VSUBS 2.54023f
C952 VN.n3 VSUBS 0.949191f
C953 VN.t3 VSUBS 2.65746f
C954 VN.n4 VSUBS 0.963874f
C955 VN.n5 VSUBS 0.204165f
C956 VN.n6 VSUBS 0.061993f
C957 VN.n7 VSUBS 0.031852f
C958 VN.n8 VSUBS 0.061993f
C959 VN.n9 VSUBS 0.039401f
C960 VN.n10 VSUBS 0.039401f
C961 VN.n11 VSUBS 0.059625f
C962 VN.n12 VSUBS 0.025175f
C963 VN.t0 VSUBS 2.61387f
C964 VN.n13 VSUBS 0.972063f
C965 VN.n14 VSUBS 0.036901f
C966 VN.n15 VSUBS 0.052576f
C967 VN.t2 VSUBS 2.54023f
C968 VN.n16 VSUBS 0.897962f
C969 VN.n17 VSUBS 0.039401f
C970 VN.t4 VSUBS 2.54023f
C971 VN.n18 VSUBS 0.949191f
C972 VN.t5 VSUBS 2.65746f
C973 VN.n19 VSUBS 0.963874f
C974 VN.n20 VSUBS 0.204165f
C975 VN.n21 VSUBS 0.061993f
C976 VN.n22 VSUBS 0.031852f
C977 VN.n23 VSUBS 0.061993f
C978 VN.n24 VSUBS 0.039401f
C979 VN.n25 VSUBS 0.039401f
C980 VN.n26 VSUBS 0.059625f
C981 VN.n27 VSUBS 0.025175f
C982 VN.t1 VSUBS 2.61387f
C983 VN.n28 VSUBS 0.972063f
C984 VN.n29 VSUBS 2.17917f
.ends

