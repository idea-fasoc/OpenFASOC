* NGSPICE file created from diff_pair_sample_0415.ext - technology: sky130A

.subckt diff_pair_sample_0415 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t10 w_n3600_n4048# sky130_fd_pr__pfet_01v8 ad=2.541 pd=15.73 as=6.006 ps=31.58 w=15.4 l=2.3
X1 B.t11 B.t9 B.t10 w_n3600_n4048# sky130_fd_pr__pfet_01v8 ad=6.006 pd=31.58 as=0 ps=0 w=15.4 l=2.3
X2 VTAIL.t1 VN.t0 VDD2.t7 w_n3600_n4048# sky130_fd_pr__pfet_01v8 ad=2.541 pd=15.73 as=2.541 ps=15.73 w=15.4 l=2.3
X3 VDD2.t6 VN.t1 VTAIL.t2 w_n3600_n4048# sky130_fd_pr__pfet_01v8 ad=2.541 pd=15.73 as=2.541 ps=15.73 w=15.4 l=2.3
X4 VDD1.t6 VP.t1 VTAIL.t12 w_n3600_n4048# sky130_fd_pr__pfet_01v8 ad=2.541 pd=15.73 as=2.541 ps=15.73 w=15.4 l=2.3
X5 VDD2.t5 VN.t2 VTAIL.t0 w_n3600_n4048# sky130_fd_pr__pfet_01v8 ad=2.541 pd=15.73 as=6.006 ps=31.58 w=15.4 l=2.3
X6 VDD2.t4 VN.t3 VTAIL.t4 w_n3600_n4048# sky130_fd_pr__pfet_01v8 ad=2.541 pd=15.73 as=6.006 ps=31.58 w=15.4 l=2.3
X7 VTAIL.t15 VP.t2 VDD1.t5 w_n3600_n4048# sky130_fd_pr__pfet_01v8 ad=2.541 pd=15.73 as=2.541 ps=15.73 w=15.4 l=2.3
X8 B.t8 B.t6 B.t7 w_n3600_n4048# sky130_fd_pr__pfet_01v8 ad=6.006 pd=31.58 as=0 ps=0 w=15.4 l=2.3
X9 VTAIL.t7 VN.t4 VDD2.t3 w_n3600_n4048# sky130_fd_pr__pfet_01v8 ad=2.541 pd=15.73 as=2.541 ps=15.73 w=15.4 l=2.3
X10 VDD2.t2 VN.t5 VTAIL.t5 w_n3600_n4048# sky130_fd_pr__pfet_01v8 ad=2.541 pd=15.73 as=2.541 ps=15.73 w=15.4 l=2.3
X11 VTAIL.t9 VP.t3 VDD1.t4 w_n3600_n4048# sky130_fd_pr__pfet_01v8 ad=6.006 pd=31.58 as=2.541 ps=15.73 w=15.4 l=2.3
X12 VDD1.t3 VP.t4 VTAIL.t14 w_n3600_n4048# sky130_fd_pr__pfet_01v8 ad=2.541 pd=15.73 as=6.006 ps=31.58 w=15.4 l=2.3
X13 B.t5 B.t3 B.t4 w_n3600_n4048# sky130_fd_pr__pfet_01v8 ad=6.006 pd=31.58 as=0 ps=0 w=15.4 l=2.3
X14 B.t2 B.t0 B.t1 w_n3600_n4048# sky130_fd_pr__pfet_01v8 ad=6.006 pd=31.58 as=0 ps=0 w=15.4 l=2.3
X15 VDD1.t2 VP.t5 VTAIL.t8 w_n3600_n4048# sky130_fd_pr__pfet_01v8 ad=2.541 pd=15.73 as=2.541 ps=15.73 w=15.4 l=2.3
X16 VTAIL.t13 VP.t6 VDD1.t1 w_n3600_n4048# sky130_fd_pr__pfet_01v8 ad=2.541 pd=15.73 as=2.541 ps=15.73 w=15.4 l=2.3
X17 VTAIL.t11 VP.t7 VDD1.t0 w_n3600_n4048# sky130_fd_pr__pfet_01v8 ad=6.006 pd=31.58 as=2.541 ps=15.73 w=15.4 l=2.3
X18 VTAIL.t6 VN.t6 VDD2.t1 w_n3600_n4048# sky130_fd_pr__pfet_01v8 ad=6.006 pd=31.58 as=2.541 ps=15.73 w=15.4 l=2.3
X19 VTAIL.t3 VN.t7 VDD2.t0 w_n3600_n4048# sky130_fd_pr__pfet_01v8 ad=6.006 pd=31.58 as=2.541 ps=15.73 w=15.4 l=2.3
R0 VP.n15 VP.t7 192.149
R1 VP.n36 VP.t3 161.365
R2 VP.n43 VP.t1 161.365
R3 VP.n55 VP.t2 161.365
R4 VP.n63 VP.t0 161.365
R5 VP.n33 VP.t4 161.365
R6 VP.n25 VP.t6 161.365
R7 VP.n14 VP.t5 161.365
R8 VP.n16 VP.n13 161.3
R9 VP.n18 VP.n17 161.3
R10 VP.n19 VP.n12 161.3
R11 VP.n21 VP.n20 161.3
R12 VP.n22 VP.n11 161.3
R13 VP.n24 VP.n23 161.3
R14 VP.n26 VP.n10 161.3
R15 VP.n28 VP.n27 161.3
R16 VP.n29 VP.n9 161.3
R17 VP.n31 VP.n30 161.3
R18 VP.n32 VP.n8 161.3
R19 VP.n62 VP.n0 161.3
R20 VP.n61 VP.n60 161.3
R21 VP.n59 VP.n1 161.3
R22 VP.n58 VP.n57 161.3
R23 VP.n56 VP.n2 161.3
R24 VP.n54 VP.n53 161.3
R25 VP.n52 VP.n3 161.3
R26 VP.n51 VP.n50 161.3
R27 VP.n49 VP.n4 161.3
R28 VP.n48 VP.n47 161.3
R29 VP.n46 VP.n5 161.3
R30 VP.n45 VP.n44 161.3
R31 VP.n42 VP.n6 161.3
R32 VP.n41 VP.n40 161.3
R33 VP.n39 VP.n7 161.3
R34 VP.n38 VP.n37 161.3
R35 VP.n36 VP.n35 101.317
R36 VP.n64 VP.n63 101.317
R37 VP.n34 VP.n33 101.317
R38 VP.n15 VP.n14 69.2325
R39 VP.n50 VP.n49 56.5617
R40 VP.n20 VP.n19 56.5617
R41 VP.n42 VP.n41 52.2023
R42 VP.n57 VP.n1 52.2023
R43 VP.n27 VP.n9 52.2023
R44 VP.n35 VP.n34 52.0072
R45 VP.n41 VP.n7 28.9518
R46 VP.n61 VP.n1 28.9518
R47 VP.n31 VP.n9 28.9518
R48 VP.n37 VP.n7 24.5923
R49 VP.n44 VP.n42 24.5923
R50 VP.n48 VP.n5 24.5923
R51 VP.n49 VP.n48 24.5923
R52 VP.n50 VP.n3 24.5923
R53 VP.n54 VP.n3 24.5923
R54 VP.n57 VP.n56 24.5923
R55 VP.n62 VP.n61 24.5923
R56 VP.n32 VP.n31 24.5923
R57 VP.n20 VP.n11 24.5923
R58 VP.n24 VP.n11 24.5923
R59 VP.n27 VP.n26 24.5923
R60 VP.n18 VP.n13 24.5923
R61 VP.n19 VP.n18 24.5923
R62 VP.n44 VP.n43 21.3954
R63 VP.n56 VP.n55 21.3954
R64 VP.n26 VP.n25 21.3954
R65 VP.n16 VP.n15 10.0465
R66 VP.n37 VP.n36 9.59132
R67 VP.n63 VP.n62 9.59132
R68 VP.n33 VP.n32 9.59132
R69 VP.n43 VP.n5 3.19744
R70 VP.n55 VP.n54 3.19744
R71 VP.n25 VP.n24 3.19744
R72 VP.n14 VP.n13 3.19744
R73 VP.n34 VP.n8 0.278335
R74 VP.n38 VP.n35 0.278335
R75 VP.n64 VP.n0 0.278335
R76 VP.n17 VP.n16 0.189894
R77 VP.n17 VP.n12 0.189894
R78 VP.n21 VP.n12 0.189894
R79 VP.n22 VP.n21 0.189894
R80 VP.n23 VP.n22 0.189894
R81 VP.n23 VP.n10 0.189894
R82 VP.n28 VP.n10 0.189894
R83 VP.n29 VP.n28 0.189894
R84 VP.n30 VP.n29 0.189894
R85 VP.n30 VP.n8 0.189894
R86 VP.n39 VP.n38 0.189894
R87 VP.n40 VP.n39 0.189894
R88 VP.n40 VP.n6 0.189894
R89 VP.n45 VP.n6 0.189894
R90 VP.n46 VP.n45 0.189894
R91 VP.n47 VP.n46 0.189894
R92 VP.n47 VP.n4 0.189894
R93 VP.n51 VP.n4 0.189894
R94 VP.n52 VP.n51 0.189894
R95 VP.n53 VP.n52 0.189894
R96 VP.n53 VP.n2 0.189894
R97 VP.n58 VP.n2 0.189894
R98 VP.n59 VP.n58 0.189894
R99 VP.n60 VP.n59 0.189894
R100 VP.n60 VP.n0 0.189894
R101 VP VP.n64 0.153485
R102 VTAIL.n690 VTAIL.n610 756.745
R103 VTAIL.n82 VTAIL.n2 756.745
R104 VTAIL.n168 VTAIL.n88 756.745
R105 VTAIL.n256 VTAIL.n176 756.745
R106 VTAIL.n604 VTAIL.n524 756.745
R107 VTAIL.n516 VTAIL.n436 756.745
R108 VTAIL.n430 VTAIL.n350 756.745
R109 VTAIL.n342 VTAIL.n262 756.745
R110 VTAIL.n639 VTAIL.n638 585
R111 VTAIL.n641 VTAIL.n640 585
R112 VTAIL.n634 VTAIL.n633 585
R113 VTAIL.n647 VTAIL.n646 585
R114 VTAIL.n649 VTAIL.n648 585
R115 VTAIL.n630 VTAIL.n629 585
R116 VTAIL.n655 VTAIL.n654 585
R117 VTAIL.n657 VTAIL.n656 585
R118 VTAIL.n626 VTAIL.n625 585
R119 VTAIL.n663 VTAIL.n662 585
R120 VTAIL.n665 VTAIL.n664 585
R121 VTAIL.n622 VTAIL.n621 585
R122 VTAIL.n671 VTAIL.n670 585
R123 VTAIL.n673 VTAIL.n672 585
R124 VTAIL.n618 VTAIL.n617 585
R125 VTAIL.n680 VTAIL.n679 585
R126 VTAIL.n681 VTAIL.n616 585
R127 VTAIL.n683 VTAIL.n682 585
R128 VTAIL.n614 VTAIL.n613 585
R129 VTAIL.n689 VTAIL.n688 585
R130 VTAIL.n691 VTAIL.n690 585
R131 VTAIL.n31 VTAIL.n30 585
R132 VTAIL.n33 VTAIL.n32 585
R133 VTAIL.n26 VTAIL.n25 585
R134 VTAIL.n39 VTAIL.n38 585
R135 VTAIL.n41 VTAIL.n40 585
R136 VTAIL.n22 VTAIL.n21 585
R137 VTAIL.n47 VTAIL.n46 585
R138 VTAIL.n49 VTAIL.n48 585
R139 VTAIL.n18 VTAIL.n17 585
R140 VTAIL.n55 VTAIL.n54 585
R141 VTAIL.n57 VTAIL.n56 585
R142 VTAIL.n14 VTAIL.n13 585
R143 VTAIL.n63 VTAIL.n62 585
R144 VTAIL.n65 VTAIL.n64 585
R145 VTAIL.n10 VTAIL.n9 585
R146 VTAIL.n72 VTAIL.n71 585
R147 VTAIL.n73 VTAIL.n8 585
R148 VTAIL.n75 VTAIL.n74 585
R149 VTAIL.n6 VTAIL.n5 585
R150 VTAIL.n81 VTAIL.n80 585
R151 VTAIL.n83 VTAIL.n82 585
R152 VTAIL.n117 VTAIL.n116 585
R153 VTAIL.n119 VTAIL.n118 585
R154 VTAIL.n112 VTAIL.n111 585
R155 VTAIL.n125 VTAIL.n124 585
R156 VTAIL.n127 VTAIL.n126 585
R157 VTAIL.n108 VTAIL.n107 585
R158 VTAIL.n133 VTAIL.n132 585
R159 VTAIL.n135 VTAIL.n134 585
R160 VTAIL.n104 VTAIL.n103 585
R161 VTAIL.n141 VTAIL.n140 585
R162 VTAIL.n143 VTAIL.n142 585
R163 VTAIL.n100 VTAIL.n99 585
R164 VTAIL.n149 VTAIL.n148 585
R165 VTAIL.n151 VTAIL.n150 585
R166 VTAIL.n96 VTAIL.n95 585
R167 VTAIL.n158 VTAIL.n157 585
R168 VTAIL.n159 VTAIL.n94 585
R169 VTAIL.n161 VTAIL.n160 585
R170 VTAIL.n92 VTAIL.n91 585
R171 VTAIL.n167 VTAIL.n166 585
R172 VTAIL.n169 VTAIL.n168 585
R173 VTAIL.n205 VTAIL.n204 585
R174 VTAIL.n207 VTAIL.n206 585
R175 VTAIL.n200 VTAIL.n199 585
R176 VTAIL.n213 VTAIL.n212 585
R177 VTAIL.n215 VTAIL.n214 585
R178 VTAIL.n196 VTAIL.n195 585
R179 VTAIL.n221 VTAIL.n220 585
R180 VTAIL.n223 VTAIL.n222 585
R181 VTAIL.n192 VTAIL.n191 585
R182 VTAIL.n229 VTAIL.n228 585
R183 VTAIL.n231 VTAIL.n230 585
R184 VTAIL.n188 VTAIL.n187 585
R185 VTAIL.n237 VTAIL.n236 585
R186 VTAIL.n239 VTAIL.n238 585
R187 VTAIL.n184 VTAIL.n183 585
R188 VTAIL.n246 VTAIL.n245 585
R189 VTAIL.n247 VTAIL.n182 585
R190 VTAIL.n249 VTAIL.n248 585
R191 VTAIL.n180 VTAIL.n179 585
R192 VTAIL.n255 VTAIL.n254 585
R193 VTAIL.n257 VTAIL.n256 585
R194 VTAIL.n605 VTAIL.n604 585
R195 VTAIL.n603 VTAIL.n602 585
R196 VTAIL.n528 VTAIL.n527 585
R197 VTAIL.n532 VTAIL.n530 585
R198 VTAIL.n597 VTAIL.n596 585
R199 VTAIL.n595 VTAIL.n594 585
R200 VTAIL.n534 VTAIL.n533 585
R201 VTAIL.n589 VTAIL.n588 585
R202 VTAIL.n587 VTAIL.n586 585
R203 VTAIL.n538 VTAIL.n537 585
R204 VTAIL.n581 VTAIL.n580 585
R205 VTAIL.n579 VTAIL.n578 585
R206 VTAIL.n542 VTAIL.n541 585
R207 VTAIL.n573 VTAIL.n572 585
R208 VTAIL.n571 VTAIL.n570 585
R209 VTAIL.n546 VTAIL.n545 585
R210 VTAIL.n565 VTAIL.n564 585
R211 VTAIL.n563 VTAIL.n562 585
R212 VTAIL.n550 VTAIL.n549 585
R213 VTAIL.n557 VTAIL.n556 585
R214 VTAIL.n555 VTAIL.n554 585
R215 VTAIL.n517 VTAIL.n516 585
R216 VTAIL.n515 VTAIL.n514 585
R217 VTAIL.n440 VTAIL.n439 585
R218 VTAIL.n444 VTAIL.n442 585
R219 VTAIL.n509 VTAIL.n508 585
R220 VTAIL.n507 VTAIL.n506 585
R221 VTAIL.n446 VTAIL.n445 585
R222 VTAIL.n501 VTAIL.n500 585
R223 VTAIL.n499 VTAIL.n498 585
R224 VTAIL.n450 VTAIL.n449 585
R225 VTAIL.n493 VTAIL.n492 585
R226 VTAIL.n491 VTAIL.n490 585
R227 VTAIL.n454 VTAIL.n453 585
R228 VTAIL.n485 VTAIL.n484 585
R229 VTAIL.n483 VTAIL.n482 585
R230 VTAIL.n458 VTAIL.n457 585
R231 VTAIL.n477 VTAIL.n476 585
R232 VTAIL.n475 VTAIL.n474 585
R233 VTAIL.n462 VTAIL.n461 585
R234 VTAIL.n469 VTAIL.n468 585
R235 VTAIL.n467 VTAIL.n466 585
R236 VTAIL.n431 VTAIL.n430 585
R237 VTAIL.n429 VTAIL.n428 585
R238 VTAIL.n354 VTAIL.n353 585
R239 VTAIL.n358 VTAIL.n356 585
R240 VTAIL.n423 VTAIL.n422 585
R241 VTAIL.n421 VTAIL.n420 585
R242 VTAIL.n360 VTAIL.n359 585
R243 VTAIL.n415 VTAIL.n414 585
R244 VTAIL.n413 VTAIL.n412 585
R245 VTAIL.n364 VTAIL.n363 585
R246 VTAIL.n407 VTAIL.n406 585
R247 VTAIL.n405 VTAIL.n404 585
R248 VTAIL.n368 VTAIL.n367 585
R249 VTAIL.n399 VTAIL.n398 585
R250 VTAIL.n397 VTAIL.n396 585
R251 VTAIL.n372 VTAIL.n371 585
R252 VTAIL.n391 VTAIL.n390 585
R253 VTAIL.n389 VTAIL.n388 585
R254 VTAIL.n376 VTAIL.n375 585
R255 VTAIL.n383 VTAIL.n382 585
R256 VTAIL.n381 VTAIL.n380 585
R257 VTAIL.n343 VTAIL.n342 585
R258 VTAIL.n341 VTAIL.n340 585
R259 VTAIL.n266 VTAIL.n265 585
R260 VTAIL.n270 VTAIL.n268 585
R261 VTAIL.n335 VTAIL.n334 585
R262 VTAIL.n333 VTAIL.n332 585
R263 VTAIL.n272 VTAIL.n271 585
R264 VTAIL.n327 VTAIL.n326 585
R265 VTAIL.n325 VTAIL.n324 585
R266 VTAIL.n276 VTAIL.n275 585
R267 VTAIL.n319 VTAIL.n318 585
R268 VTAIL.n317 VTAIL.n316 585
R269 VTAIL.n280 VTAIL.n279 585
R270 VTAIL.n311 VTAIL.n310 585
R271 VTAIL.n309 VTAIL.n308 585
R272 VTAIL.n284 VTAIL.n283 585
R273 VTAIL.n303 VTAIL.n302 585
R274 VTAIL.n301 VTAIL.n300 585
R275 VTAIL.n288 VTAIL.n287 585
R276 VTAIL.n295 VTAIL.n294 585
R277 VTAIL.n293 VTAIL.n292 585
R278 VTAIL.n637 VTAIL.t0 327.466
R279 VTAIL.n29 VTAIL.t3 327.466
R280 VTAIL.n115 VTAIL.t10 327.466
R281 VTAIL.n203 VTAIL.t9 327.466
R282 VTAIL.n553 VTAIL.t14 327.466
R283 VTAIL.n465 VTAIL.t11 327.466
R284 VTAIL.n379 VTAIL.t4 327.466
R285 VTAIL.n291 VTAIL.t6 327.466
R286 VTAIL.n640 VTAIL.n639 171.744
R287 VTAIL.n640 VTAIL.n633 171.744
R288 VTAIL.n647 VTAIL.n633 171.744
R289 VTAIL.n648 VTAIL.n647 171.744
R290 VTAIL.n648 VTAIL.n629 171.744
R291 VTAIL.n655 VTAIL.n629 171.744
R292 VTAIL.n656 VTAIL.n655 171.744
R293 VTAIL.n656 VTAIL.n625 171.744
R294 VTAIL.n663 VTAIL.n625 171.744
R295 VTAIL.n664 VTAIL.n663 171.744
R296 VTAIL.n664 VTAIL.n621 171.744
R297 VTAIL.n671 VTAIL.n621 171.744
R298 VTAIL.n672 VTAIL.n671 171.744
R299 VTAIL.n672 VTAIL.n617 171.744
R300 VTAIL.n680 VTAIL.n617 171.744
R301 VTAIL.n681 VTAIL.n680 171.744
R302 VTAIL.n682 VTAIL.n681 171.744
R303 VTAIL.n682 VTAIL.n613 171.744
R304 VTAIL.n689 VTAIL.n613 171.744
R305 VTAIL.n690 VTAIL.n689 171.744
R306 VTAIL.n32 VTAIL.n31 171.744
R307 VTAIL.n32 VTAIL.n25 171.744
R308 VTAIL.n39 VTAIL.n25 171.744
R309 VTAIL.n40 VTAIL.n39 171.744
R310 VTAIL.n40 VTAIL.n21 171.744
R311 VTAIL.n47 VTAIL.n21 171.744
R312 VTAIL.n48 VTAIL.n47 171.744
R313 VTAIL.n48 VTAIL.n17 171.744
R314 VTAIL.n55 VTAIL.n17 171.744
R315 VTAIL.n56 VTAIL.n55 171.744
R316 VTAIL.n56 VTAIL.n13 171.744
R317 VTAIL.n63 VTAIL.n13 171.744
R318 VTAIL.n64 VTAIL.n63 171.744
R319 VTAIL.n64 VTAIL.n9 171.744
R320 VTAIL.n72 VTAIL.n9 171.744
R321 VTAIL.n73 VTAIL.n72 171.744
R322 VTAIL.n74 VTAIL.n73 171.744
R323 VTAIL.n74 VTAIL.n5 171.744
R324 VTAIL.n81 VTAIL.n5 171.744
R325 VTAIL.n82 VTAIL.n81 171.744
R326 VTAIL.n118 VTAIL.n117 171.744
R327 VTAIL.n118 VTAIL.n111 171.744
R328 VTAIL.n125 VTAIL.n111 171.744
R329 VTAIL.n126 VTAIL.n125 171.744
R330 VTAIL.n126 VTAIL.n107 171.744
R331 VTAIL.n133 VTAIL.n107 171.744
R332 VTAIL.n134 VTAIL.n133 171.744
R333 VTAIL.n134 VTAIL.n103 171.744
R334 VTAIL.n141 VTAIL.n103 171.744
R335 VTAIL.n142 VTAIL.n141 171.744
R336 VTAIL.n142 VTAIL.n99 171.744
R337 VTAIL.n149 VTAIL.n99 171.744
R338 VTAIL.n150 VTAIL.n149 171.744
R339 VTAIL.n150 VTAIL.n95 171.744
R340 VTAIL.n158 VTAIL.n95 171.744
R341 VTAIL.n159 VTAIL.n158 171.744
R342 VTAIL.n160 VTAIL.n159 171.744
R343 VTAIL.n160 VTAIL.n91 171.744
R344 VTAIL.n167 VTAIL.n91 171.744
R345 VTAIL.n168 VTAIL.n167 171.744
R346 VTAIL.n206 VTAIL.n205 171.744
R347 VTAIL.n206 VTAIL.n199 171.744
R348 VTAIL.n213 VTAIL.n199 171.744
R349 VTAIL.n214 VTAIL.n213 171.744
R350 VTAIL.n214 VTAIL.n195 171.744
R351 VTAIL.n221 VTAIL.n195 171.744
R352 VTAIL.n222 VTAIL.n221 171.744
R353 VTAIL.n222 VTAIL.n191 171.744
R354 VTAIL.n229 VTAIL.n191 171.744
R355 VTAIL.n230 VTAIL.n229 171.744
R356 VTAIL.n230 VTAIL.n187 171.744
R357 VTAIL.n237 VTAIL.n187 171.744
R358 VTAIL.n238 VTAIL.n237 171.744
R359 VTAIL.n238 VTAIL.n183 171.744
R360 VTAIL.n246 VTAIL.n183 171.744
R361 VTAIL.n247 VTAIL.n246 171.744
R362 VTAIL.n248 VTAIL.n247 171.744
R363 VTAIL.n248 VTAIL.n179 171.744
R364 VTAIL.n255 VTAIL.n179 171.744
R365 VTAIL.n256 VTAIL.n255 171.744
R366 VTAIL.n604 VTAIL.n603 171.744
R367 VTAIL.n603 VTAIL.n527 171.744
R368 VTAIL.n532 VTAIL.n527 171.744
R369 VTAIL.n596 VTAIL.n532 171.744
R370 VTAIL.n596 VTAIL.n595 171.744
R371 VTAIL.n595 VTAIL.n533 171.744
R372 VTAIL.n588 VTAIL.n533 171.744
R373 VTAIL.n588 VTAIL.n587 171.744
R374 VTAIL.n587 VTAIL.n537 171.744
R375 VTAIL.n580 VTAIL.n537 171.744
R376 VTAIL.n580 VTAIL.n579 171.744
R377 VTAIL.n579 VTAIL.n541 171.744
R378 VTAIL.n572 VTAIL.n541 171.744
R379 VTAIL.n572 VTAIL.n571 171.744
R380 VTAIL.n571 VTAIL.n545 171.744
R381 VTAIL.n564 VTAIL.n545 171.744
R382 VTAIL.n564 VTAIL.n563 171.744
R383 VTAIL.n563 VTAIL.n549 171.744
R384 VTAIL.n556 VTAIL.n549 171.744
R385 VTAIL.n556 VTAIL.n555 171.744
R386 VTAIL.n516 VTAIL.n515 171.744
R387 VTAIL.n515 VTAIL.n439 171.744
R388 VTAIL.n444 VTAIL.n439 171.744
R389 VTAIL.n508 VTAIL.n444 171.744
R390 VTAIL.n508 VTAIL.n507 171.744
R391 VTAIL.n507 VTAIL.n445 171.744
R392 VTAIL.n500 VTAIL.n445 171.744
R393 VTAIL.n500 VTAIL.n499 171.744
R394 VTAIL.n499 VTAIL.n449 171.744
R395 VTAIL.n492 VTAIL.n449 171.744
R396 VTAIL.n492 VTAIL.n491 171.744
R397 VTAIL.n491 VTAIL.n453 171.744
R398 VTAIL.n484 VTAIL.n453 171.744
R399 VTAIL.n484 VTAIL.n483 171.744
R400 VTAIL.n483 VTAIL.n457 171.744
R401 VTAIL.n476 VTAIL.n457 171.744
R402 VTAIL.n476 VTAIL.n475 171.744
R403 VTAIL.n475 VTAIL.n461 171.744
R404 VTAIL.n468 VTAIL.n461 171.744
R405 VTAIL.n468 VTAIL.n467 171.744
R406 VTAIL.n430 VTAIL.n429 171.744
R407 VTAIL.n429 VTAIL.n353 171.744
R408 VTAIL.n358 VTAIL.n353 171.744
R409 VTAIL.n422 VTAIL.n358 171.744
R410 VTAIL.n422 VTAIL.n421 171.744
R411 VTAIL.n421 VTAIL.n359 171.744
R412 VTAIL.n414 VTAIL.n359 171.744
R413 VTAIL.n414 VTAIL.n413 171.744
R414 VTAIL.n413 VTAIL.n363 171.744
R415 VTAIL.n406 VTAIL.n363 171.744
R416 VTAIL.n406 VTAIL.n405 171.744
R417 VTAIL.n405 VTAIL.n367 171.744
R418 VTAIL.n398 VTAIL.n367 171.744
R419 VTAIL.n398 VTAIL.n397 171.744
R420 VTAIL.n397 VTAIL.n371 171.744
R421 VTAIL.n390 VTAIL.n371 171.744
R422 VTAIL.n390 VTAIL.n389 171.744
R423 VTAIL.n389 VTAIL.n375 171.744
R424 VTAIL.n382 VTAIL.n375 171.744
R425 VTAIL.n382 VTAIL.n381 171.744
R426 VTAIL.n342 VTAIL.n341 171.744
R427 VTAIL.n341 VTAIL.n265 171.744
R428 VTAIL.n270 VTAIL.n265 171.744
R429 VTAIL.n334 VTAIL.n270 171.744
R430 VTAIL.n334 VTAIL.n333 171.744
R431 VTAIL.n333 VTAIL.n271 171.744
R432 VTAIL.n326 VTAIL.n271 171.744
R433 VTAIL.n326 VTAIL.n325 171.744
R434 VTAIL.n325 VTAIL.n275 171.744
R435 VTAIL.n318 VTAIL.n275 171.744
R436 VTAIL.n318 VTAIL.n317 171.744
R437 VTAIL.n317 VTAIL.n279 171.744
R438 VTAIL.n310 VTAIL.n279 171.744
R439 VTAIL.n310 VTAIL.n309 171.744
R440 VTAIL.n309 VTAIL.n283 171.744
R441 VTAIL.n302 VTAIL.n283 171.744
R442 VTAIL.n302 VTAIL.n301 171.744
R443 VTAIL.n301 VTAIL.n287 171.744
R444 VTAIL.n294 VTAIL.n287 171.744
R445 VTAIL.n294 VTAIL.n293 171.744
R446 VTAIL.n639 VTAIL.t0 85.8723
R447 VTAIL.n31 VTAIL.t3 85.8723
R448 VTAIL.n117 VTAIL.t10 85.8723
R449 VTAIL.n205 VTAIL.t9 85.8723
R450 VTAIL.n555 VTAIL.t14 85.8723
R451 VTAIL.n467 VTAIL.t11 85.8723
R452 VTAIL.n381 VTAIL.t4 85.8723
R453 VTAIL.n293 VTAIL.t6 85.8723
R454 VTAIL.n523 VTAIL.n522 54.3551
R455 VTAIL.n349 VTAIL.n348 54.3551
R456 VTAIL.n1 VTAIL.n0 54.3549
R457 VTAIL.n175 VTAIL.n174 54.3549
R458 VTAIL.n695 VTAIL.n694 32.9611
R459 VTAIL.n87 VTAIL.n86 32.9611
R460 VTAIL.n173 VTAIL.n172 32.9611
R461 VTAIL.n261 VTAIL.n260 32.9611
R462 VTAIL.n609 VTAIL.n608 32.9611
R463 VTAIL.n521 VTAIL.n520 32.9611
R464 VTAIL.n435 VTAIL.n434 32.9611
R465 VTAIL.n347 VTAIL.n346 32.9611
R466 VTAIL.n695 VTAIL.n609 27.91
R467 VTAIL.n347 VTAIL.n261 27.91
R468 VTAIL.n638 VTAIL.n637 16.3895
R469 VTAIL.n30 VTAIL.n29 16.3895
R470 VTAIL.n116 VTAIL.n115 16.3895
R471 VTAIL.n204 VTAIL.n203 16.3895
R472 VTAIL.n554 VTAIL.n553 16.3895
R473 VTAIL.n466 VTAIL.n465 16.3895
R474 VTAIL.n380 VTAIL.n379 16.3895
R475 VTAIL.n292 VTAIL.n291 16.3895
R476 VTAIL.n683 VTAIL.n614 13.1884
R477 VTAIL.n75 VTAIL.n6 13.1884
R478 VTAIL.n161 VTAIL.n92 13.1884
R479 VTAIL.n249 VTAIL.n180 13.1884
R480 VTAIL.n530 VTAIL.n528 13.1884
R481 VTAIL.n442 VTAIL.n440 13.1884
R482 VTAIL.n356 VTAIL.n354 13.1884
R483 VTAIL.n268 VTAIL.n266 13.1884
R484 VTAIL.n641 VTAIL.n636 12.8005
R485 VTAIL.n684 VTAIL.n616 12.8005
R486 VTAIL.n688 VTAIL.n687 12.8005
R487 VTAIL.n33 VTAIL.n28 12.8005
R488 VTAIL.n76 VTAIL.n8 12.8005
R489 VTAIL.n80 VTAIL.n79 12.8005
R490 VTAIL.n119 VTAIL.n114 12.8005
R491 VTAIL.n162 VTAIL.n94 12.8005
R492 VTAIL.n166 VTAIL.n165 12.8005
R493 VTAIL.n207 VTAIL.n202 12.8005
R494 VTAIL.n250 VTAIL.n182 12.8005
R495 VTAIL.n254 VTAIL.n253 12.8005
R496 VTAIL.n602 VTAIL.n601 12.8005
R497 VTAIL.n598 VTAIL.n597 12.8005
R498 VTAIL.n557 VTAIL.n552 12.8005
R499 VTAIL.n514 VTAIL.n513 12.8005
R500 VTAIL.n510 VTAIL.n509 12.8005
R501 VTAIL.n469 VTAIL.n464 12.8005
R502 VTAIL.n428 VTAIL.n427 12.8005
R503 VTAIL.n424 VTAIL.n423 12.8005
R504 VTAIL.n383 VTAIL.n378 12.8005
R505 VTAIL.n340 VTAIL.n339 12.8005
R506 VTAIL.n336 VTAIL.n335 12.8005
R507 VTAIL.n295 VTAIL.n290 12.8005
R508 VTAIL.n642 VTAIL.n634 12.0247
R509 VTAIL.n679 VTAIL.n678 12.0247
R510 VTAIL.n691 VTAIL.n612 12.0247
R511 VTAIL.n34 VTAIL.n26 12.0247
R512 VTAIL.n71 VTAIL.n70 12.0247
R513 VTAIL.n83 VTAIL.n4 12.0247
R514 VTAIL.n120 VTAIL.n112 12.0247
R515 VTAIL.n157 VTAIL.n156 12.0247
R516 VTAIL.n169 VTAIL.n90 12.0247
R517 VTAIL.n208 VTAIL.n200 12.0247
R518 VTAIL.n245 VTAIL.n244 12.0247
R519 VTAIL.n257 VTAIL.n178 12.0247
R520 VTAIL.n605 VTAIL.n526 12.0247
R521 VTAIL.n594 VTAIL.n531 12.0247
R522 VTAIL.n558 VTAIL.n550 12.0247
R523 VTAIL.n517 VTAIL.n438 12.0247
R524 VTAIL.n506 VTAIL.n443 12.0247
R525 VTAIL.n470 VTAIL.n462 12.0247
R526 VTAIL.n431 VTAIL.n352 12.0247
R527 VTAIL.n420 VTAIL.n357 12.0247
R528 VTAIL.n384 VTAIL.n376 12.0247
R529 VTAIL.n343 VTAIL.n264 12.0247
R530 VTAIL.n332 VTAIL.n269 12.0247
R531 VTAIL.n296 VTAIL.n288 12.0247
R532 VTAIL.n646 VTAIL.n645 11.249
R533 VTAIL.n677 VTAIL.n618 11.249
R534 VTAIL.n692 VTAIL.n610 11.249
R535 VTAIL.n38 VTAIL.n37 11.249
R536 VTAIL.n69 VTAIL.n10 11.249
R537 VTAIL.n84 VTAIL.n2 11.249
R538 VTAIL.n124 VTAIL.n123 11.249
R539 VTAIL.n155 VTAIL.n96 11.249
R540 VTAIL.n170 VTAIL.n88 11.249
R541 VTAIL.n212 VTAIL.n211 11.249
R542 VTAIL.n243 VTAIL.n184 11.249
R543 VTAIL.n258 VTAIL.n176 11.249
R544 VTAIL.n606 VTAIL.n524 11.249
R545 VTAIL.n593 VTAIL.n534 11.249
R546 VTAIL.n562 VTAIL.n561 11.249
R547 VTAIL.n518 VTAIL.n436 11.249
R548 VTAIL.n505 VTAIL.n446 11.249
R549 VTAIL.n474 VTAIL.n473 11.249
R550 VTAIL.n432 VTAIL.n350 11.249
R551 VTAIL.n419 VTAIL.n360 11.249
R552 VTAIL.n388 VTAIL.n387 11.249
R553 VTAIL.n344 VTAIL.n262 11.249
R554 VTAIL.n331 VTAIL.n272 11.249
R555 VTAIL.n300 VTAIL.n299 11.249
R556 VTAIL.n649 VTAIL.n632 10.4732
R557 VTAIL.n674 VTAIL.n673 10.4732
R558 VTAIL.n41 VTAIL.n24 10.4732
R559 VTAIL.n66 VTAIL.n65 10.4732
R560 VTAIL.n127 VTAIL.n110 10.4732
R561 VTAIL.n152 VTAIL.n151 10.4732
R562 VTAIL.n215 VTAIL.n198 10.4732
R563 VTAIL.n240 VTAIL.n239 10.4732
R564 VTAIL.n590 VTAIL.n589 10.4732
R565 VTAIL.n565 VTAIL.n548 10.4732
R566 VTAIL.n502 VTAIL.n501 10.4732
R567 VTAIL.n477 VTAIL.n460 10.4732
R568 VTAIL.n416 VTAIL.n415 10.4732
R569 VTAIL.n391 VTAIL.n374 10.4732
R570 VTAIL.n328 VTAIL.n327 10.4732
R571 VTAIL.n303 VTAIL.n286 10.4732
R572 VTAIL.n650 VTAIL.n630 9.69747
R573 VTAIL.n670 VTAIL.n620 9.69747
R574 VTAIL.n42 VTAIL.n22 9.69747
R575 VTAIL.n62 VTAIL.n12 9.69747
R576 VTAIL.n128 VTAIL.n108 9.69747
R577 VTAIL.n148 VTAIL.n98 9.69747
R578 VTAIL.n216 VTAIL.n196 9.69747
R579 VTAIL.n236 VTAIL.n186 9.69747
R580 VTAIL.n586 VTAIL.n536 9.69747
R581 VTAIL.n566 VTAIL.n546 9.69747
R582 VTAIL.n498 VTAIL.n448 9.69747
R583 VTAIL.n478 VTAIL.n458 9.69747
R584 VTAIL.n412 VTAIL.n362 9.69747
R585 VTAIL.n392 VTAIL.n372 9.69747
R586 VTAIL.n324 VTAIL.n274 9.69747
R587 VTAIL.n304 VTAIL.n284 9.69747
R588 VTAIL.n694 VTAIL.n693 9.45567
R589 VTAIL.n86 VTAIL.n85 9.45567
R590 VTAIL.n172 VTAIL.n171 9.45567
R591 VTAIL.n260 VTAIL.n259 9.45567
R592 VTAIL.n608 VTAIL.n607 9.45567
R593 VTAIL.n520 VTAIL.n519 9.45567
R594 VTAIL.n434 VTAIL.n433 9.45567
R595 VTAIL.n346 VTAIL.n345 9.45567
R596 VTAIL.n693 VTAIL.n692 9.3005
R597 VTAIL.n612 VTAIL.n611 9.3005
R598 VTAIL.n687 VTAIL.n686 9.3005
R599 VTAIL.n659 VTAIL.n658 9.3005
R600 VTAIL.n628 VTAIL.n627 9.3005
R601 VTAIL.n653 VTAIL.n652 9.3005
R602 VTAIL.n651 VTAIL.n650 9.3005
R603 VTAIL.n632 VTAIL.n631 9.3005
R604 VTAIL.n645 VTAIL.n644 9.3005
R605 VTAIL.n643 VTAIL.n642 9.3005
R606 VTAIL.n636 VTAIL.n635 9.3005
R607 VTAIL.n661 VTAIL.n660 9.3005
R608 VTAIL.n624 VTAIL.n623 9.3005
R609 VTAIL.n667 VTAIL.n666 9.3005
R610 VTAIL.n669 VTAIL.n668 9.3005
R611 VTAIL.n620 VTAIL.n619 9.3005
R612 VTAIL.n675 VTAIL.n674 9.3005
R613 VTAIL.n677 VTAIL.n676 9.3005
R614 VTAIL.n678 VTAIL.n615 9.3005
R615 VTAIL.n685 VTAIL.n684 9.3005
R616 VTAIL.n85 VTAIL.n84 9.3005
R617 VTAIL.n4 VTAIL.n3 9.3005
R618 VTAIL.n79 VTAIL.n78 9.3005
R619 VTAIL.n51 VTAIL.n50 9.3005
R620 VTAIL.n20 VTAIL.n19 9.3005
R621 VTAIL.n45 VTAIL.n44 9.3005
R622 VTAIL.n43 VTAIL.n42 9.3005
R623 VTAIL.n24 VTAIL.n23 9.3005
R624 VTAIL.n37 VTAIL.n36 9.3005
R625 VTAIL.n35 VTAIL.n34 9.3005
R626 VTAIL.n28 VTAIL.n27 9.3005
R627 VTAIL.n53 VTAIL.n52 9.3005
R628 VTAIL.n16 VTAIL.n15 9.3005
R629 VTAIL.n59 VTAIL.n58 9.3005
R630 VTAIL.n61 VTAIL.n60 9.3005
R631 VTAIL.n12 VTAIL.n11 9.3005
R632 VTAIL.n67 VTAIL.n66 9.3005
R633 VTAIL.n69 VTAIL.n68 9.3005
R634 VTAIL.n70 VTAIL.n7 9.3005
R635 VTAIL.n77 VTAIL.n76 9.3005
R636 VTAIL.n171 VTAIL.n170 9.3005
R637 VTAIL.n90 VTAIL.n89 9.3005
R638 VTAIL.n165 VTAIL.n164 9.3005
R639 VTAIL.n137 VTAIL.n136 9.3005
R640 VTAIL.n106 VTAIL.n105 9.3005
R641 VTAIL.n131 VTAIL.n130 9.3005
R642 VTAIL.n129 VTAIL.n128 9.3005
R643 VTAIL.n110 VTAIL.n109 9.3005
R644 VTAIL.n123 VTAIL.n122 9.3005
R645 VTAIL.n121 VTAIL.n120 9.3005
R646 VTAIL.n114 VTAIL.n113 9.3005
R647 VTAIL.n139 VTAIL.n138 9.3005
R648 VTAIL.n102 VTAIL.n101 9.3005
R649 VTAIL.n145 VTAIL.n144 9.3005
R650 VTAIL.n147 VTAIL.n146 9.3005
R651 VTAIL.n98 VTAIL.n97 9.3005
R652 VTAIL.n153 VTAIL.n152 9.3005
R653 VTAIL.n155 VTAIL.n154 9.3005
R654 VTAIL.n156 VTAIL.n93 9.3005
R655 VTAIL.n163 VTAIL.n162 9.3005
R656 VTAIL.n259 VTAIL.n258 9.3005
R657 VTAIL.n178 VTAIL.n177 9.3005
R658 VTAIL.n253 VTAIL.n252 9.3005
R659 VTAIL.n225 VTAIL.n224 9.3005
R660 VTAIL.n194 VTAIL.n193 9.3005
R661 VTAIL.n219 VTAIL.n218 9.3005
R662 VTAIL.n217 VTAIL.n216 9.3005
R663 VTAIL.n198 VTAIL.n197 9.3005
R664 VTAIL.n211 VTAIL.n210 9.3005
R665 VTAIL.n209 VTAIL.n208 9.3005
R666 VTAIL.n202 VTAIL.n201 9.3005
R667 VTAIL.n227 VTAIL.n226 9.3005
R668 VTAIL.n190 VTAIL.n189 9.3005
R669 VTAIL.n233 VTAIL.n232 9.3005
R670 VTAIL.n235 VTAIL.n234 9.3005
R671 VTAIL.n186 VTAIL.n185 9.3005
R672 VTAIL.n241 VTAIL.n240 9.3005
R673 VTAIL.n243 VTAIL.n242 9.3005
R674 VTAIL.n244 VTAIL.n181 9.3005
R675 VTAIL.n251 VTAIL.n250 9.3005
R676 VTAIL.n540 VTAIL.n539 9.3005
R677 VTAIL.n583 VTAIL.n582 9.3005
R678 VTAIL.n585 VTAIL.n584 9.3005
R679 VTAIL.n536 VTAIL.n535 9.3005
R680 VTAIL.n591 VTAIL.n590 9.3005
R681 VTAIL.n593 VTAIL.n592 9.3005
R682 VTAIL.n531 VTAIL.n529 9.3005
R683 VTAIL.n599 VTAIL.n598 9.3005
R684 VTAIL.n607 VTAIL.n606 9.3005
R685 VTAIL.n526 VTAIL.n525 9.3005
R686 VTAIL.n601 VTAIL.n600 9.3005
R687 VTAIL.n577 VTAIL.n576 9.3005
R688 VTAIL.n575 VTAIL.n574 9.3005
R689 VTAIL.n544 VTAIL.n543 9.3005
R690 VTAIL.n569 VTAIL.n568 9.3005
R691 VTAIL.n567 VTAIL.n566 9.3005
R692 VTAIL.n548 VTAIL.n547 9.3005
R693 VTAIL.n561 VTAIL.n560 9.3005
R694 VTAIL.n559 VTAIL.n558 9.3005
R695 VTAIL.n552 VTAIL.n551 9.3005
R696 VTAIL.n452 VTAIL.n451 9.3005
R697 VTAIL.n495 VTAIL.n494 9.3005
R698 VTAIL.n497 VTAIL.n496 9.3005
R699 VTAIL.n448 VTAIL.n447 9.3005
R700 VTAIL.n503 VTAIL.n502 9.3005
R701 VTAIL.n505 VTAIL.n504 9.3005
R702 VTAIL.n443 VTAIL.n441 9.3005
R703 VTAIL.n511 VTAIL.n510 9.3005
R704 VTAIL.n519 VTAIL.n518 9.3005
R705 VTAIL.n438 VTAIL.n437 9.3005
R706 VTAIL.n513 VTAIL.n512 9.3005
R707 VTAIL.n489 VTAIL.n488 9.3005
R708 VTAIL.n487 VTAIL.n486 9.3005
R709 VTAIL.n456 VTAIL.n455 9.3005
R710 VTAIL.n481 VTAIL.n480 9.3005
R711 VTAIL.n479 VTAIL.n478 9.3005
R712 VTAIL.n460 VTAIL.n459 9.3005
R713 VTAIL.n473 VTAIL.n472 9.3005
R714 VTAIL.n471 VTAIL.n470 9.3005
R715 VTAIL.n464 VTAIL.n463 9.3005
R716 VTAIL.n366 VTAIL.n365 9.3005
R717 VTAIL.n409 VTAIL.n408 9.3005
R718 VTAIL.n411 VTAIL.n410 9.3005
R719 VTAIL.n362 VTAIL.n361 9.3005
R720 VTAIL.n417 VTAIL.n416 9.3005
R721 VTAIL.n419 VTAIL.n418 9.3005
R722 VTAIL.n357 VTAIL.n355 9.3005
R723 VTAIL.n425 VTAIL.n424 9.3005
R724 VTAIL.n433 VTAIL.n432 9.3005
R725 VTAIL.n352 VTAIL.n351 9.3005
R726 VTAIL.n427 VTAIL.n426 9.3005
R727 VTAIL.n403 VTAIL.n402 9.3005
R728 VTAIL.n401 VTAIL.n400 9.3005
R729 VTAIL.n370 VTAIL.n369 9.3005
R730 VTAIL.n395 VTAIL.n394 9.3005
R731 VTAIL.n393 VTAIL.n392 9.3005
R732 VTAIL.n374 VTAIL.n373 9.3005
R733 VTAIL.n387 VTAIL.n386 9.3005
R734 VTAIL.n385 VTAIL.n384 9.3005
R735 VTAIL.n378 VTAIL.n377 9.3005
R736 VTAIL.n278 VTAIL.n277 9.3005
R737 VTAIL.n321 VTAIL.n320 9.3005
R738 VTAIL.n323 VTAIL.n322 9.3005
R739 VTAIL.n274 VTAIL.n273 9.3005
R740 VTAIL.n329 VTAIL.n328 9.3005
R741 VTAIL.n331 VTAIL.n330 9.3005
R742 VTAIL.n269 VTAIL.n267 9.3005
R743 VTAIL.n337 VTAIL.n336 9.3005
R744 VTAIL.n345 VTAIL.n344 9.3005
R745 VTAIL.n264 VTAIL.n263 9.3005
R746 VTAIL.n339 VTAIL.n338 9.3005
R747 VTAIL.n315 VTAIL.n314 9.3005
R748 VTAIL.n313 VTAIL.n312 9.3005
R749 VTAIL.n282 VTAIL.n281 9.3005
R750 VTAIL.n307 VTAIL.n306 9.3005
R751 VTAIL.n305 VTAIL.n304 9.3005
R752 VTAIL.n286 VTAIL.n285 9.3005
R753 VTAIL.n299 VTAIL.n298 9.3005
R754 VTAIL.n297 VTAIL.n296 9.3005
R755 VTAIL.n290 VTAIL.n289 9.3005
R756 VTAIL.n654 VTAIL.n653 8.92171
R757 VTAIL.n669 VTAIL.n622 8.92171
R758 VTAIL.n46 VTAIL.n45 8.92171
R759 VTAIL.n61 VTAIL.n14 8.92171
R760 VTAIL.n132 VTAIL.n131 8.92171
R761 VTAIL.n147 VTAIL.n100 8.92171
R762 VTAIL.n220 VTAIL.n219 8.92171
R763 VTAIL.n235 VTAIL.n188 8.92171
R764 VTAIL.n585 VTAIL.n538 8.92171
R765 VTAIL.n570 VTAIL.n569 8.92171
R766 VTAIL.n497 VTAIL.n450 8.92171
R767 VTAIL.n482 VTAIL.n481 8.92171
R768 VTAIL.n411 VTAIL.n364 8.92171
R769 VTAIL.n396 VTAIL.n395 8.92171
R770 VTAIL.n323 VTAIL.n276 8.92171
R771 VTAIL.n308 VTAIL.n307 8.92171
R772 VTAIL.n657 VTAIL.n628 8.14595
R773 VTAIL.n666 VTAIL.n665 8.14595
R774 VTAIL.n49 VTAIL.n20 8.14595
R775 VTAIL.n58 VTAIL.n57 8.14595
R776 VTAIL.n135 VTAIL.n106 8.14595
R777 VTAIL.n144 VTAIL.n143 8.14595
R778 VTAIL.n223 VTAIL.n194 8.14595
R779 VTAIL.n232 VTAIL.n231 8.14595
R780 VTAIL.n582 VTAIL.n581 8.14595
R781 VTAIL.n573 VTAIL.n544 8.14595
R782 VTAIL.n494 VTAIL.n493 8.14595
R783 VTAIL.n485 VTAIL.n456 8.14595
R784 VTAIL.n408 VTAIL.n407 8.14595
R785 VTAIL.n399 VTAIL.n370 8.14595
R786 VTAIL.n320 VTAIL.n319 8.14595
R787 VTAIL.n311 VTAIL.n282 8.14595
R788 VTAIL.n658 VTAIL.n626 7.3702
R789 VTAIL.n662 VTAIL.n624 7.3702
R790 VTAIL.n50 VTAIL.n18 7.3702
R791 VTAIL.n54 VTAIL.n16 7.3702
R792 VTAIL.n136 VTAIL.n104 7.3702
R793 VTAIL.n140 VTAIL.n102 7.3702
R794 VTAIL.n224 VTAIL.n192 7.3702
R795 VTAIL.n228 VTAIL.n190 7.3702
R796 VTAIL.n578 VTAIL.n540 7.3702
R797 VTAIL.n574 VTAIL.n542 7.3702
R798 VTAIL.n490 VTAIL.n452 7.3702
R799 VTAIL.n486 VTAIL.n454 7.3702
R800 VTAIL.n404 VTAIL.n366 7.3702
R801 VTAIL.n400 VTAIL.n368 7.3702
R802 VTAIL.n316 VTAIL.n278 7.3702
R803 VTAIL.n312 VTAIL.n280 7.3702
R804 VTAIL.n661 VTAIL.n626 6.59444
R805 VTAIL.n662 VTAIL.n661 6.59444
R806 VTAIL.n53 VTAIL.n18 6.59444
R807 VTAIL.n54 VTAIL.n53 6.59444
R808 VTAIL.n139 VTAIL.n104 6.59444
R809 VTAIL.n140 VTAIL.n139 6.59444
R810 VTAIL.n227 VTAIL.n192 6.59444
R811 VTAIL.n228 VTAIL.n227 6.59444
R812 VTAIL.n578 VTAIL.n577 6.59444
R813 VTAIL.n577 VTAIL.n542 6.59444
R814 VTAIL.n490 VTAIL.n489 6.59444
R815 VTAIL.n489 VTAIL.n454 6.59444
R816 VTAIL.n404 VTAIL.n403 6.59444
R817 VTAIL.n403 VTAIL.n368 6.59444
R818 VTAIL.n316 VTAIL.n315 6.59444
R819 VTAIL.n315 VTAIL.n280 6.59444
R820 VTAIL.n658 VTAIL.n657 5.81868
R821 VTAIL.n665 VTAIL.n624 5.81868
R822 VTAIL.n50 VTAIL.n49 5.81868
R823 VTAIL.n57 VTAIL.n16 5.81868
R824 VTAIL.n136 VTAIL.n135 5.81868
R825 VTAIL.n143 VTAIL.n102 5.81868
R826 VTAIL.n224 VTAIL.n223 5.81868
R827 VTAIL.n231 VTAIL.n190 5.81868
R828 VTAIL.n581 VTAIL.n540 5.81868
R829 VTAIL.n574 VTAIL.n573 5.81868
R830 VTAIL.n493 VTAIL.n452 5.81868
R831 VTAIL.n486 VTAIL.n485 5.81868
R832 VTAIL.n407 VTAIL.n366 5.81868
R833 VTAIL.n400 VTAIL.n399 5.81868
R834 VTAIL.n319 VTAIL.n278 5.81868
R835 VTAIL.n312 VTAIL.n311 5.81868
R836 VTAIL.n654 VTAIL.n628 5.04292
R837 VTAIL.n666 VTAIL.n622 5.04292
R838 VTAIL.n46 VTAIL.n20 5.04292
R839 VTAIL.n58 VTAIL.n14 5.04292
R840 VTAIL.n132 VTAIL.n106 5.04292
R841 VTAIL.n144 VTAIL.n100 5.04292
R842 VTAIL.n220 VTAIL.n194 5.04292
R843 VTAIL.n232 VTAIL.n188 5.04292
R844 VTAIL.n582 VTAIL.n538 5.04292
R845 VTAIL.n570 VTAIL.n544 5.04292
R846 VTAIL.n494 VTAIL.n450 5.04292
R847 VTAIL.n482 VTAIL.n456 5.04292
R848 VTAIL.n408 VTAIL.n364 5.04292
R849 VTAIL.n396 VTAIL.n370 5.04292
R850 VTAIL.n320 VTAIL.n276 5.04292
R851 VTAIL.n308 VTAIL.n282 5.04292
R852 VTAIL.n653 VTAIL.n630 4.26717
R853 VTAIL.n670 VTAIL.n669 4.26717
R854 VTAIL.n45 VTAIL.n22 4.26717
R855 VTAIL.n62 VTAIL.n61 4.26717
R856 VTAIL.n131 VTAIL.n108 4.26717
R857 VTAIL.n148 VTAIL.n147 4.26717
R858 VTAIL.n219 VTAIL.n196 4.26717
R859 VTAIL.n236 VTAIL.n235 4.26717
R860 VTAIL.n586 VTAIL.n585 4.26717
R861 VTAIL.n569 VTAIL.n546 4.26717
R862 VTAIL.n498 VTAIL.n497 4.26717
R863 VTAIL.n481 VTAIL.n458 4.26717
R864 VTAIL.n412 VTAIL.n411 4.26717
R865 VTAIL.n395 VTAIL.n372 4.26717
R866 VTAIL.n324 VTAIL.n323 4.26717
R867 VTAIL.n307 VTAIL.n284 4.26717
R868 VTAIL.n637 VTAIL.n635 3.70982
R869 VTAIL.n29 VTAIL.n27 3.70982
R870 VTAIL.n115 VTAIL.n113 3.70982
R871 VTAIL.n203 VTAIL.n201 3.70982
R872 VTAIL.n553 VTAIL.n551 3.70982
R873 VTAIL.n465 VTAIL.n463 3.70982
R874 VTAIL.n379 VTAIL.n377 3.70982
R875 VTAIL.n291 VTAIL.n289 3.70982
R876 VTAIL.n650 VTAIL.n649 3.49141
R877 VTAIL.n673 VTAIL.n620 3.49141
R878 VTAIL.n42 VTAIL.n41 3.49141
R879 VTAIL.n65 VTAIL.n12 3.49141
R880 VTAIL.n128 VTAIL.n127 3.49141
R881 VTAIL.n151 VTAIL.n98 3.49141
R882 VTAIL.n216 VTAIL.n215 3.49141
R883 VTAIL.n239 VTAIL.n186 3.49141
R884 VTAIL.n589 VTAIL.n536 3.49141
R885 VTAIL.n566 VTAIL.n565 3.49141
R886 VTAIL.n501 VTAIL.n448 3.49141
R887 VTAIL.n478 VTAIL.n477 3.49141
R888 VTAIL.n415 VTAIL.n362 3.49141
R889 VTAIL.n392 VTAIL.n391 3.49141
R890 VTAIL.n327 VTAIL.n274 3.49141
R891 VTAIL.n304 VTAIL.n303 3.49141
R892 VTAIL.n646 VTAIL.n632 2.71565
R893 VTAIL.n674 VTAIL.n618 2.71565
R894 VTAIL.n694 VTAIL.n610 2.71565
R895 VTAIL.n38 VTAIL.n24 2.71565
R896 VTAIL.n66 VTAIL.n10 2.71565
R897 VTAIL.n86 VTAIL.n2 2.71565
R898 VTAIL.n124 VTAIL.n110 2.71565
R899 VTAIL.n152 VTAIL.n96 2.71565
R900 VTAIL.n172 VTAIL.n88 2.71565
R901 VTAIL.n212 VTAIL.n198 2.71565
R902 VTAIL.n240 VTAIL.n184 2.71565
R903 VTAIL.n260 VTAIL.n176 2.71565
R904 VTAIL.n608 VTAIL.n524 2.71565
R905 VTAIL.n590 VTAIL.n534 2.71565
R906 VTAIL.n562 VTAIL.n548 2.71565
R907 VTAIL.n520 VTAIL.n436 2.71565
R908 VTAIL.n502 VTAIL.n446 2.71565
R909 VTAIL.n474 VTAIL.n460 2.71565
R910 VTAIL.n434 VTAIL.n350 2.71565
R911 VTAIL.n416 VTAIL.n360 2.71565
R912 VTAIL.n388 VTAIL.n374 2.71565
R913 VTAIL.n346 VTAIL.n262 2.71565
R914 VTAIL.n328 VTAIL.n272 2.71565
R915 VTAIL.n300 VTAIL.n286 2.71565
R916 VTAIL.n349 VTAIL.n347 2.26774
R917 VTAIL.n435 VTAIL.n349 2.26774
R918 VTAIL.n523 VTAIL.n521 2.26774
R919 VTAIL.n609 VTAIL.n523 2.26774
R920 VTAIL.n261 VTAIL.n175 2.26774
R921 VTAIL.n175 VTAIL.n173 2.26774
R922 VTAIL.n87 VTAIL.n1 2.26774
R923 VTAIL VTAIL.n695 2.20955
R924 VTAIL.n0 VTAIL.t2 2.11121
R925 VTAIL.n0 VTAIL.t1 2.11121
R926 VTAIL.n174 VTAIL.t12 2.11121
R927 VTAIL.n174 VTAIL.t15 2.11121
R928 VTAIL.n522 VTAIL.t8 2.11121
R929 VTAIL.n522 VTAIL.t13 2.11121
R930 VTAIL.n348 VTAIL.t5 2.11121
R931 VTAIL.n348 VTAIL.t7 2.11121
R932 VTAIL.n645 VTAIL.n634 1.93989
R933 VTAIL.n679 VTAIL.n677 1.93989
R934 VTAIL.n692 VTAIL.n691 1.93989
R935 VTAIL.n37 VTAIL.n26 1.93989
R936 VTAIL.n71 VTAIL.n69 1.93989
R937 VTAIL.n84 VTAIL.n83 1.93989
R938 VTAIL.n123 VTAIL.n112 1.93989
R939 VTAIL.n157 VTAIL.n155 1.93989
R940 VTAIL.n170 VTAIL.n169 1.93989
R941 VTAIL.n211 VTAIL.n200 1.93989
R942 VTAIL.n245 VTAIL.n243 1.93989
R943 VTAIL.n258 VTAIL.n257 1.93989
R944 VTAIL.n606 VTAIL.n605 1.93989
R945 VTAIL.n594 VTAIL.n593 1.93989
R946 VTAIL.n561 VTAIL.n550 1.93989
R947 VTAIL.n518 VTAIL.n517 1.93989
R948 VTAIL.n506 VTAIL.n505 1.93989
R949 VTAIL.n473 VTAIL.n462 1.93989
R950 VTAIL.n432 VTAIL.n431 1.93989
R951 VTAIL.n420 VTAIL.n419 1.93989
R952 VTAIL.n387 VTAIL.n376 1.93989
R953 VTAIL.n344 VTAIL.n343 1.93989
R954 VTAIL.n332 VTAIL.n331 1.93989
R955 VTAIL.n299 VTAIL.n288 1.93989
R956 VTAIL.n642 VTAIL.n641 1.16414
R957 VTAIL.n678 VTAIL.n616 1.16414
R958 VTAIL.n688 VTAIL.n612 1.16414
R959 VTAIL.n34 VTAIL.n33 1.16414
R960 VTAIL.n70 VTAIL.n8 1.16414
R961 VTAIL.n80 VTAIL.n4 1.16414
R962 VTAIL.n120 VTAIL.n119 1.16414
R963 VTAIL.n156 VTAIL.n94 1.16414
R964 VTAIL.n166 VTAIL.n90 1.16414
R965 VTAIL.n208 VTAIL.n207 1.16414
R966 VTAIL.n244 VTAIL.n182 1.16414
R967 VTAIL.n254 VTAIL.n178 1.16414
R968 VTAIL.n602 VTAIL.n526 1.16414
R969 VTAIL.n597 VTAIL.n531 1.16414
R970 VTAIL.n558 VTAIL.n557 1.16414
R971 VTAIL.n514 VTAIL.n438 1.16414
R972 VTAIL.n509 VTAIL.n443 1.16414
R973 VTAIL.n470 VTAIL.n469 1.16414
R974 VTAIL.n428 VTAIL.n352 1.16414
R975 VTAIL.n423 VTAIL.n357 1.16414
R976 VTAIL.n384 VTAIL.n383 1.16414
R977 VTAIL.n340 VTAIL.n264 1.16414
R978 VTAIL.n335 VTAIL.n269 1.16414
R979 VTAIL.n296 VTAIL.n295 1.16414
R980 VTAIL.n521 VTAIL.n435 0.470328
R981 VTAIL.n173 VTAIL.n87 0.470328
R982 VTAIL.n638 VTAIL.n636 0.388379
R983 VTAIL.n684 VTAIL.n683 0.388379
R984 VTAIL.n687 VTAIL.n614 0.388379
R985 VTAIL.n30 VTAIL.n28 0.388379
R986 VTAIL.n76 VTAIL.n75 0.388379
R987 VTAIL.n79 VTAIL.n6 0.388379
R988 VTAIL.n116 VTAIL.n114 0.388379
R989 VTAIL.n162 VTAIL.n161 0.388379
R990 VTAIL.n165 VTAIL.n92 0.388379
R991 VTAIL.n204 VTAIL.n202 0.388379
R992 VTAIL.n250 VTAIL.n249 0.388379
R993 VTAIL.n253 VTAIL.n180 0.388379
R994 VTAIL.n601 VTAIL.n528 0.388379
R995 VTAIL.n598 VTAIL.n530 0.388379
R996 VTAIL.n554 VTAIL.n552 0.388379
R997 VTAIL.n513 VTAIL.n440 0.388379
R998 VTAIL.n510 VTAIL.n442 0.388379
R999 VTAIL.n466 VTAIL.n464 0.388379
R1000 VTAIL.n427 VTAIL.n354 0.388379
R1001 VTAIL.n424 VTAIL.n356 0.388379
R1002 VTAIL.n380 VTAIL.n378 0.388379
R1003 VTAIL.n339 VTAIL.n266 0.388379
R1004 VTAIL.n336 VTAIL.n268 0.388379
R1005 VTAIL.n292 VTAIL.n290 0.388379
R1006 VTAIL.n643 VTAIL.n635 0.155672
R1007 VTAIL.n644 VTAIL.n643 0.155672
R1008 VTAIL.n644 VTAIL.n631 0.155672
R1009 VTAIL.n651 VTAIL.n631 0.155672
R1010 VTAIL.n652 VTAIL.n651 0.155672
R1011 VTAIL.n652 VTAIL.n627 0.155672
R1012 VTAIL.n659 VTAIL.n627 0.155672
R1013 VTAIL.n660 VTAIL.n659 0.155672
R1014 VTAIL.n660 VTAIL.n623 0.155672
R1015 VTAIL.n667 VTAIL.n623 0.155672
R1016 VTAIL.n668 VTAIL.n667 0.155672
R1017 VTAIL.n668 VTAIL.n619 0.155672
R1018 VTAIL.n675 VTAIL.n619 0.155672
R1019 VTAIL.n676 VTAIL.n675 0.155672
R1020 VTAIL.n676 VTAIL.n615 0.155672
R1021 VTAIL.n685 VTAIL.n615 0.155672
R1022 VTAIL.n686 VTAIL.n685 0.155672
R1023 VTAIL.n686 VTAIL.n611 0.155672
R1024 VTAIL.n693 VTAIL.n611 0.155672
R1025 VTAIL.n35 VTAIL.n27 0.155672
R1026 VTAIL.n36 VTAIL.n35 0.155672
R1027 VTAIL.n36 VTAIL.n23 0.155672
R1028 VTAIL.n43 VTAIL.n23 0.155672
R1029 VTAIL.n44 VTAIL.n43 0.155672
R1030 VTAIL.n44 VTAIL.n19 0.155672
R1031 VTAIL.n51 VTAIL.n19 0.155672
R1032 VTAIL.n52 VTAIL.n51 0.155672
R1033 VTAIL.n52 VTAIL.n15 0.155672
R1034 VTAIL.n59 VTAIL.n15 0.155672
R1035 VTAIL.n60 VTAIL.n59 0.155672
R1036 VTAIL.n60 VTAIL.n11 0.155672
R1037 VTAIL.n67 VTAIL.n11 0.155672
R1038 VTAIL.n68 VTAIL.n67 0.155672
R1039 VTAIL.n68 VTAIL.n7 0.155672
R1040 VTAIL.n77 VTAIL.n7 0.155672
R1041 VTAIL.n78 VTAIL.n77 0.155672
R1042 VTAIL.n78 VTAIL.n3 0.155672
R1043 VTAIL.n85 VTAIL.n3 0.155672
R1044 VTAIL.n121 VTAIL.n113 0.155672
R1045 VTAIL.n122 VTAIL.n121 0.155672
R1046 VTAIL.n122 VTAIL.n109 0.155672
R1047 VTAIL.n129 VTAIL.n109 0.155672
R1048 VTAIL.n130 VTAIL.n129 0.155672
R1049 VTAIL.n130 VTAIL.n105 0.155672
R1050 VTAIL.n137 VTAIL.n105 0.155672
R1051 VTAIL.n138 VTAIL.n137 0.155672
R1052 VTAIL.n138 VTAIL.n101 0.155672
R1053 VTAIL.n145 VTAIL.n101 0.155672
R1054 VTAIL.n146 VTAIL.n145 0.155672
R1055 VTAIL.n146 VTAIL.n97 0.155672
R1056 VTAIL.n153 VTAIL.n97 0.155672
R1057 VTAIL.n154 VTAIL.n153 0.155672
R1058 VTAIL.n154 VTAIL.n93 0.155672
R1059 VTAIL.n163 VTAIL.n93 0.155672
R1060 VTAIL.n164 VTAIL.n163 0.155672
R1061 VTAIL.n164 VTAIL.n89 0.155672
R1062 VTAIL.n171 VTAIL.n89 0.155672
R1063 VTAIL.n209 VTAIL.n201 0.155672
R1064 VTAIL.n210 VTAIL.n209 0.155672
R1065 VTAIL.n210 VTAIL.n197 0.155672
R1066 VTAIL.n217 VTAIL.n197 0.155672
R1067 VTAIL.n218 VTAIL.n217 0.155672
R1068 VTAIL.n218 VTAIL.n193 0.155672
R1069 VTAIL.n225 VTAIL.n193 0.155672
R1070 VTAIL.n226 VTAIL.n225 0.155672
R1071 VTAIL.n226 VTAIL.n189 0.155672
R1072 VTAIL.n233 VTAIL.n189 0.155672
R1073 VTAIL.n234 VTAIL.n233 0.155672
R1074 VTAIL.n234 VTAIL.n185 0.155672
R1075 VTAIL.n241 VTAIL.n185 0.155672
R1076 VTAIL.n242 VTAIL.n241 0.155672
R1077 VTAIL.n242 VTAIL.n181 0.155672
R1078 VTAIL.n251 VTAIL.n181 0.155672
R1079 VTAIL.n252 VTAIL.n251 0.155672
R1080 VTAIL.n252 VTAIL.n177 0.155672
R1081 VTAIL.n259 VTAIL.n177 0.155672
R1082 VTAIL.n607 VTAIL.n525 0.155672
R1083 VTAIL.n600 VTAIL.n525 0.155672
R1084 VTAIL.n600 VTAIL.n599 0.155672
R1085 VTAIL.n599 VTAIL.n529 0.155672
R1086 VTAIL.n592 VTAIL.n529 0.155672
R1087 VTAIL.n592 VTAIL.n591 0.155672
R1088 VTAIL.n591 VTAIL.n535 0.155672
R1089 VTAIL.n584 VTAIL.n535 0.155672
R1090 VTAIL.n584 VTAIL.n583 0.155672
R1091 VTAIL.n583 VTAIL.n539 0.155672
R1092 VTAIL.n576 VTAIL.n539 0.155672
R1093 VTAIL.n576 VTAIL.n575 0.155672
R1094 VTAIL.n575 VTAIL.n543 0.155672
R1095 VTAIL.n568 VTAIL.n543 0.155672
R1096 VTAIL.n568 VTAIL.n567 0.155672
R1097 VTAIL.n567 VTAIL.n547 0.155672
R1098 VTAIL.n560 VTAIL.n547 0.155672
R1099 VTAIL.n560 VTAIL.n559 0.155672
R1100 VTAIL.n559 VTAIL.n551 0.155672
R1101 VTAIL.n519 VTAIL.n437 0.155672
R1102 VTAIL.n512 VTAIL.n437 0.155672
R1103 VTAIL.n512 VTAIL.n511 0.155672
R1104 VTAIL.n511 VTAIL.n441 0.155672
R1105 VTAIL.n504 VTAIL.n441 0.155672
R1106 VTAIL.n504 VTAIL.n503 0.155672
R1107 VTAIL.n503 VTAIL.n447 0.155672
R1108 VTAIL.n496 VTAIL.n447 0.155672
R1109 VTAIL.n496 VTAIL.n495 0.155672
R1110 VTAIL.n495 VTAIL.n451 0.155672
R1111 VTAIL.n488 VTAIL.n451 0.155672
R1112 VTAIL.n488 VTAIL.n487 0.155672
R1113 VTAIL.n487 VTAIL.n455 0.155672
R1114 VTAIL.n480 VTAIL.n455 0.155672
R1115 VTAIL.n480 VTAIL.n479 0.155672
R1116 VTAIL.n479 VTAIL.n459 0.155672
R1117 VTAIL.n472 VTAIL.n459 0.155672
R1118 VTAIL.n472 VTAIL.n471 0.155672
R1119 VTAIL.n471 VTAIL.n463 0.155672
R1120 VTAIL.n433 VTAIL.n351 0.155672
R1121 VTAIL.n426 VTAIL.n351 0.155672
R1122 VTAIL.n426 VTAIL.n425 0.155672
R1123 VTAIL.n425 VTAIL.n355 0.155672
R1124 VTAIL.n418 VTAIL.n355 0.155672
R1125 VTAIL.n418 VTAIL.n417 0.155672
R1126 VTAIL.n417 VTAIL.n361 0.155672
R1127 VTAIL.n410 VTAIL.n361 0.155672
R1128 VTAIL.n410 VTAIL.n409 0.155672
R1129 VTAIL.n409 VTAIL.n365 0.155672
R1130 VTAIL.n402 VTAIL.n365 0.155672
R1131 VTAIL.n402 VTAIL.n401 0.155672
R1132 VTAIL.n401 VTAIL.n369 0.155672
R1133 VTAIL.n394 VTAIL.n369 0.155672
R1134 VTAIL.n394 VTAIL.n393 0.155672
R1135 VTAIL.n393 VTAIL.n373 0.155672
R1136 VTAIL.n386 VTAIL.n373 0.155672
R1137 VTAIL.n386 VTAIL.n385 0.155672
R1138 VTAIL.n385 VTAIL.n377 0.155672
R1139 VTAIL.n345 VTAIL.n263 0.155672
R1140 VTAIL.n338 VTAIL.n263 0.155672
R1141 VTAIL.n338 VTAIL.n337 0.155672
R1142 VTAIL.n337 VTAIL.n267 0.155672
R1143 VTAIL.n330 VTAIL.n267 0.155672
R1144 VTAIL.n330 VTAIL.n329 0.155672
R1145 VTAIL.n329 VTAIL.n273 0.155672
R1146 VTAIL.n322 VTAIL.n273 0.155672
R1147 VTAIL.n322 VTAIL.n321 0.155672
R1148 VTAIL.n321 VTAIL.n277 0.155672
R1149 VTAIL.n314 VTAIL.n277 0.155672
R1150 VTAIL.n314 VTAIL.n313 0.155672
R1151 VTAIL.n313 VTAIL.n281 0.155672
R1152 VTAIL.n306 VTAIL.n281 0.155672
R1153 VTAIL.n306 VTAIL.n305 0.155672
R1154 VTAIL.n305 VTAIL.n285 0.155672
R1155 VTAIL.n298 VTAIL.n285 0.155672
R1156 VTAIL.n298 VTAIL.n297 0.155672
R1157 VTAIL.n297 VTAIL.n289 0.155672
R1158 VTAIL VTAIL.n1 0.0586897
R1159 VDD1 VDD1.n0 72.2257
R1160 VDD1.n3 VDD1.n2 72.112
R1161 VDD1.n3 VDD1.n1 72.112
R1162 VDD1.n5 VDD1.n4 71.0337
R1163 VDD1.n5 VDD1.n3 47.7768
R1164 VDD1.n4 VDD1.t1 2.11121
R1165 VDD1.n4 VDD1.t3 2.11121
R1166 VDD1.n0 VDD1.t0 2.11121
R1167 VDD1.n0 VDD1.t2 2.11121
R1168 VDD1.n2 VDD1.t5 2.11121
R1169 VDD1.n2 VDD1.t7 2.11121
R1170 VDD1.n1 VDD1.t4 2.11121
R1171 VDD1.n1 VDD1.t6 2.11121
R1172 VDD1 VDD1.n5 1.07593
R1173 B.n601 B.n86 585
R1174 B.n603 B.n602 585
R1175 B.n604 B.n85 585
R1176 B.n606 B.n605 585
R1177 B.n607 B.n84 585
R1178 B.n609 B.n608 585
R1179 B.n610 B.n83 585
R1180 B.n612 B.n611 585
R1181 B.n613 B.n82 585
R1182 B.n615 B.n614 585
R1183 B.n616 B.n81 585
R1184 B.n618 B.n617 585
R1185 B.n619 B.n80 585
R1186 B.n621 B.n620 585
R1187 B.n622 B.n79 585
R1188 B.n624 B.n623 585
R1189 B.n625 B.n78 585
R1190 B.n627 B.n626 585
R1191 B.n628 B.n77 585
R1192 B.n630 B.n629 585
R1193 B.n631 B.n76 585
R1194 B.n633 B.n632 585
R1195 B.n634 B.n75 585
R1196 B.n636 B.n635 585
R1197 B.n637 B.n74 585
R1198 B.n639 B.n638 585
R1199 B.n640 B.n73 585
R1200 B.n642 B.n641 585
R1201 B.n643 B.n72 585
R1202 B.n645 B.n644 585
R1203 B.n646 B.n71 585
R1204 B.n648 B.n647 585
R1205 B.n649 B.n70 585
R1206 B.n651 B.n650 585
R1207 B.n652 B.n69 585
R1208 B.n654 B.n653 585
R1209 B.n655 B.n68 585
R1210 B.n657 B.n656 585
R1211 B.n658 B.n67 585
R1212 B.n660 B.n659 585
R1213 B.n661 B.n66 585
R1214 B.n663 B.n662 585
R1215 B.n664 B.n65 585
R1216 B.n666 B.n665 585
R1217 B.n667 B.n64 585
R1218 B.n669 B.n668 585
R1219 B.n670 B.n63 585
R1220 B.n672 B.n671 585
R1221 B.n673 B.n62 585
R1222 B.n675 B.n674 585
R1223 B.n676 B.n61 585
R1224 B.n678 B.n677 585
R1225 B.n680 B.n679 585
R1226 B.n681 B.n57 585
R1227 B.n683 B.n682 585
R1228 B.n684 B.n56 585
R1229 B.n686 B.n685 585
R1230 B.n687 B.n55 585
R1231 B.n689 B.n688 585
R1232 B.n690 B.n54 585
R1233 B.n692 B.n691 585
R1234 B.n694 B.n51 585
R1235 B.n696 B.n695 585
R1236 B.n697 B.n50 585
R1237 B.n699 B.n698 585
R1238 B.n700 B.n49 585
R1239 B.n702 B.n701 585
R1240 B.n703 B.n48 585
R1241 B.n705 B.n704 585
R1242 B.n706 B.n47 585
R1243 B.n708 B.n707 585
R1244 B.n709 B.n46 585
R1245 B.n711 B.n710 585
R1246 B.n712 B.n45 585
R1247 B.n714 B.n713 585
R1248 B.n715 B.n44 585
R1249 B.n717 B.n716 585
R1250 B.n718 B.n43 585
R1251 B.n720 B.n719 585
R1252 B.n721 B.n42 585
R1253 B.n723 B.n722 585
R1254 B.n724 B.n41 585
R1255 B.n726 B.n725 585
R1256 B.n727 B.n40 585
R1257 B.n729 B.n728 585
R1258 B.n730 B.n39 585
R1259 B.n732 B.n731 585
R1260 B.n733 B.n38 585
R1261 B.n735 B.n734 585
R1262 B.n736 B.n37 585
R1263 B.n738 B.n737 585
R1264 B.n739 B.n36 585
R1265 B.n741 B.n740 585
R1266 B.n742 B.n35 585
R1267 B.n744 B.n743 585
R1268 B.n745 B.n34 585
R1269 B.n747 B.n746 585
R1270 B.n748 B.n33 585
R1271 B.n750 B.n749 585
R1272 B.n751 B.n32 585
R1273 B.n753 B.n752 585
R1274 B.n754 B.n31 585
R1275 B.n756 B.n755 585
R1276 B.n757 B.n30 585
R1277 B.n759 B.n758 585
R1278 B.n760 B.n29 585
R1279 B.n762 B.n761 585
R1280 B.n763 B.n28 585
R1281 B.n765 B.n764 585
R1282 B.n766 B.n27 585
R1283 B.n768 B.n767 585
R1284 B.n769 B.n26 585
R1285 B.n771 B.n770 585
R1286 B.n600 B.n599 585
R1287 B.n598 B.n87 585
R1288 B.n597 B.n596 585
R1289 B.n595 B.n88 585
R1290 B.n594 B.n593 585
R1291 B.n592 B.n89 585
R1292 B.n591 B.n590 585
R1293 B.n589 B.n90 585
R1294 B.n588 B.n587 585
R1295 B.n586 B.n91 585
R1296 B.n585 B.n584 585
R1297 B.n583 B.n92 585
R1298 B.n582 B.n581 585
R1299 B.n580 B.n93 585
R1300 B.n579 B.n578 585
R1301 B.n577 B.n94 585
R1302 B.n576 B.n575 585
R1303 B.n574 B.n95 585
R1304 B.n573 B.n572 585
R1305 B.n571 B.n96 585
R1306 B.n570 B.n569 585
R1307 B.n568 B.n97 585
R1308 B.n567 B.n566 585
R1309 B.n565 B.n98 585
R1310 B.n564 B.n563 585
R1311 B.n562 B.n99 585
R1312 B.n561 B.n560 585
R1313 B.n559 B.n100 585
R1314 B.n558 B.n557 585
R1315 B.n556 B.n101 585
R1316 B.n555 B.n554 585
R1317 B.n553 B.n102 585
R1318 B.n552 B.n551 585
R1319 B.n550 B.n103 585
R1320 B.n549 B.n548 585
R1321 B.n547 B.n104 585
R1322 B.n546 B.n545 585
R1323 B.n544 B.n105 585
R1324 B.n543 B.n542 585
R1325 B.n541 B.n106 585
R1326 B.n540 B.n539 585
R1327 B.n538 B.n107 585
R1328 B.n537 B.n536 585
R1329 B.n535 B.n108 585
R1330 B.n534 B.n533 585
R1331 B.n532 B.n109 585
R1332 B.n531 B.n530 585
R1333 B.n529 B.n110 585
R1334 B.n528 B.n527 585
R1335 B.n526 B.n111 585
R1336 B.n525 B.n524 585
R1337 B.n523 B.n112 585
R1338 B.n522 B.n521 585
R1339 B.n520 B.n113 585
R1340 B.n519 B.n518 585
R1341 B.n517 B.n114 585
R1342 B.n516 B.n515 585
R1343 B.n514 B.n115 585
R1344 B.n513 B.n512 585
R1345 B.n511 B.n116 585
R1346 B.n510 B.n509 585
R1347 B.n508 B.n117 585
R1348 B.n507 B.n506 585
R1349 B.n505 B.n118 585
R1350 B.n504 B.n503 585
R1351 B.n502 B.n119 585
R1352 B.n501 B.n500 585
R1353 B.n499 B.n120 585
R1354 B.n498 B.n497 585
R1355 B.n496 B.n121 585
R1356 B.n495 B.n494 585
R1357 B.n493 B.n122 585
R1358 B.n492 B.n491 585
R1359 B.n490 B.n123 585
R1360 B.n489 B.n488 585
R1361 B.n487 B.n124 585
R1362 B.n486 B.n485 585
R1363 B.n484 B.n125 585
R1364 B.n483 B.n482 585
R1365 B.n481 B.n126 585
R1366 B.n480 B.n479 585
R1367 B.n478 B.n127 585
R1368 B.n477 B.n476 585
R1369 B.n475 B.n128 585
R1370 B.n474 B.n473 585
R1371 B.n472 B.n129 585
R1372 B.n471 B.n470 585
R1373 B.n469 B.n130 585
R1374 B.n468 B.n467 585
R1375 B.n466 B.n131 585
R1376 B.n465 B.n464 585
R1377 B.n463 B.n132 585
R1378 B.n462 B.n461 585
R1379 B.n460 B.n133 585
R1380 B.n459 B.n458 585
R1381 B.n288 B.n287 585
R1382 B.n289 B.n194 585
R1383 B.n291 B.n290 585
R1384 B.n292 B.n193 585
R1385 B.n294 B.n293 585
R1386 B.n295 B.n192 585
R1387 B.n297 B.n296 585
R1388 B.n298 B.n191 585
R1389 B.n300 B.n299 585
R1390 B.n301 B.n190 585
R1391 B.n303 B.n302 585
R1392 B.n304 B.n189 585
R1393 B.n306 B.n305 585
R1394 B.n307 B.n188 585
R1395 B.n309 B.n308 585
R1396 B.n310 B.n187 585
R1397 B.n312 B.n311 585
R1398 B.n313 B.n186 585
R1399 B.n315 B.n314 585
R1400 B.n316 B.n185 585
R1401 B.n318 B.n317 585
R1402 B.n319 B.n184 585
R1403 B.n321 B.n320 585
R1404 B.n322 B.n183 585
R1405 B.n324 B.n323 585
R1406 B.n325 B.n182 585
R1407 B.n327 B.n326 585
R1408 B.n328 B.n181 585
R1409 B.n330 B.n329 585
R1410 B.n331 B.n180 585
R1411 B.n333 B.n332 585
R1412 B.n334 B.n179 585
R1413 B.n336 B.n335 585
R1414 B.n337 B.n178 585
R1415 B.n339 B.n338 585
R1416 B.n340 B.n177 585
R1417 B.n342 B.n341 585
R1418 B.n343 B.n176 585
R1419 B.n345 B.n344 585
R1420 B.n346 B.n175 585
R1421 B.n348 B.n347 585
R1422 B.n349 B.n174 585
R1423 B.n351 B.n350 585
R1424 B.n352 B.n173 585
R1425 B.n354 B.n353 585
R1426 B.n355 B.n172 585
R1427 B.n357 B.n356 585
R1428 B.n358 B.n171 585
R1429 B.n360 B.n359 585
R1430 B.n361 B.n170 585
R1431 B.n363 B.n362 585
R1432 B.n364 B.n167 585
R1433 B.n367 B.n366 585
R1434 B.n368 B.n166 585
R1435 B.n370 B.n369 585
R1436 B.n371 B.n165 585
R1437 B.n373 B.n372 585
R1438 B.n374 B.n164 585
R1439 B.n376 B.n375 585
R1440 B.n377 B.n163 585
R1441 B.n379 B.n378 585
R1442 B.n381 B.n380 585
R1443 B.n382 B.n159 585
R1444 B.n384 B.n383 585
R1445 B.n385 B.n158 585
R1446 B.n387 B.n386 585
R1447 B.n388 B.n157 585
R1448 B.n390 B.n389 585
R1449 B.n391 B.n156 585
R1450 B.n393 B.n392 585
R1451 B.n394 B.n155 585
R1452 B.n396 B.n395 585
R1453 B.n397 B.n154 585
R1454 B.n399 B.n398 585
R1455 B.n400 B.n153 585
R1456 B.n402 B.n401 585
R1457 B.n403 B.n152 585
R1458 B.n405 B.n404 585
R1459 B.n406 B.n151 585
R1460 B.n408 B.n407 585
R1461 B.n409 B.n150 585
R1462 B.n411 B.n410 585
R1463 B.n412 B.n149 585
R1464 B.n414 B.n413 585
R1465 B.n415 B.n148 585
R1466 B.n417 B.n416 585
R1467 B.n418 B.n147 585
R1468 B.n420 B.n419 585
R1469 B.n421 B.n146 585
R1470 B.n423 B.n422 585
R1471 B.n424 B.n145 585
R1472 B.n426 B.n425 585
R1473 B.n427 B.n144 585
R1474 B.n429 B.n428 585
R1475 B.n430 B.n143 585
R1476 B.n432 B.n431 585
R1477 B.n433 B.n142 585
R1478 B.n435 B.n434 585
R1479 B.n436 B.n141 585
R1480 B.n438 B.n437 585
R1481 B.n439 B.n140 585
R1482 B.n441 B.n440 585
R1483 B.n442 B.n139 585
R1484 B.n444 B.n443 585
R1485 B.n445 B.n138 585
R1486 B.n447 B.n446 585
R1487 B.n448 B.n137 585
R1488 B.n450 B.n449 585
R1489 B.n451 B.n136 585
R1490 B.n453 B.n452 585
R1491 B.n454 B.n135 585
R1492 B.n456 B.n455 585
R1493 B.n457 B.n134 585
R1494 B.n286 B.n195 585
R1495 B.n285 B.n284 585
R1496 B.n283 B.n196 585
R1497 B.n282 B.n281 585
R1498 B.n280 B.n197 585
R1499 B.n279 B.n278 585
R1500 B.n277 B.n198 585
R1501 B.n276 B.n275 585
R1502 B.n274 B.n199 585
R1503 B.n273 B.n272 585
R1504 B.n271 B.n200 585
R1505 B.n270 B.n269 585
R1506 B.n268 B.n201 585
R1507 B.n267 B.n266 585
R1508 B.n265 B.n202 585
R1509 B.n264 B.n263 585
R1510 B.n262 B.n203 585
R1511 B.n261 B.n260 585
R1512 B.n259 B.n204 585
R1513 B.n258 B.n257 585
R1514 B.n256 B.n205 585
R1515 B.n255 B.n254 585
R1516 B.n253 B.n206 585
R1517 B.n252 B.n251 585
R1518 B.n250 B.n207 585
R1519 B.n249 B.n248 585
R1520 B.n247 B.n208 585
R1521 B.n246 B.n245 585
R1522 B.n244 B.n209 585
R1523 B.n243 B.n242 585
R1524 B.n241 B.n210 585
R1525 B.n240 B.n239 585
R1526 B.n238 B.n211 585
R1527 B.n237 B.n236 585
R1528 B.n235 B.n212 585
R1529 B.n234 B.n233 585
R1530 B.n232 B.n213 585
R1531 B.n231 B.n230 585
R1532 B.n229 B.n214 585
R1533 B.n228 B.n227 585
R1534 B.n226 B.n215 585
R1535 B.n225 B.n224 585
R1536 B.n223 B.n216 585
R1537 B.n222 B.n221 585
R1538 B.n220 B.n217 585
R1539 B.n219 B.n218 585
R1540 B.n2 B.n0 585
R1541 B.n841 B.n1 585
R1542 B.n840 B.n839 585
R1543 B.n838 B.n3 585
R1544 B.n837 B.n836 585
R1545 B.n835 B.n4 585
R1546 B.n834 B.n833 585
R1547 B.n832 B.n5 585
R1548 B.n831 B.n830 585
R1549 B.n829 B.n6 585
R1550 B.n828 B.n827 585
R1551 B.n826 B.n7 585
R1552 B.n825 B.n824 585
R1553 B.n823 B.n8 585
R1554 B.n822 B.n821 585
R1555 B.n820 B.n9 585
R1556 B.n819 B.n818 585
R1557 B.n817 B.n10 585
R1558 B.n816 B.n815 585
R1559 B.n814 B.n11 585
R1560 B.n813 B.n812 585
R1561 B.n811 B.n12 585
R1562 B.n810 B.n809 585
R1563 B.n808 B.n13 585
R1564 B.n807 B.n806 585
R1565 B.n805 B.n14 585
R1566 B.n804 B.n803 585
R1567 B.n802 B.n15 585
R1568 B.n801 B.n800 585
R1569 B.n799 B.n16 585
R1570 B.n798 B.n797 585
R1571 B.n796 B.n17 585
R1572 B.n795 B.n794 585
R1573 B.n793 B.n18 585
R1574 B.n792 B.n791 585
R1575 B.n790 B.n19 585
R1576 B.n789 B.n788 585
R1577 B.n787 B.n20 585
R1578 B.n786 B.n785 585
R1579 B.n784 B.n21 585
R1580 B.n783 B.n782 585
R1581 B.n781 B.n22 585
R1582 B.n780 B.n779 585
R1583 B.n778 B.n23 585
R1584 B.n777 B.n776 585
R1585 B.n775 B.n24 585
R1586 B.n774 B.n773 585
R1587 B.n772 B.n25 585
R1588 B.n843 B.n842 585
R1589 B.n160 B.t2 487.774
R1590 B.n58 B.t4 487.774
R1591 B.n168 B.t11 487.774
R1592 B.n52 B.t7 487.774
R1593 B.n288 B.n195 449.257
R1594 B.n770 B.n25 449.257
R1595 B.n458 B.n457 449.257
R1596 B.n601 B.n600 449.257
R1597 B.n161 B.t1 436.769
R1598 B.n59 B.t5 436.769
R1599 B.n169 B.t10 436.769
R1600 B.n53 B.t8 436.769
R1601 B.n160 B.t0 368.909
R1602 B.n168 B.t9 368.909
R1603 B.n52 B.t6 368.909
R1604 B.n58 B.t3 368.909
R1605 B.n284 B.n195 163.367
R1606 B.n284 B.n283 163.367
R1607 B.n283 B.n282 163.367
R1608 B.n282 B.n197 163.367
R1609 B.n278 B.n197 163.367
R1610 B.n278 B.n277 163.367
R1611 B.n277 B.n276 163.367
R1612 B.n276 B.n199 163.367
R1613 B.n272 B.n199 163.367
R1614 B.n272 B.n271 163.367
R1615 B.n271 B.n270 163.367
R1616 B.n270 B.n201 163.367
R1617 B.n266 B.n201 163.367
R1618 B.n266 B.n265 163.367
R1619 B.n265 B.n264 163.367
R1620 B.n264 B.n203 163.367
R1621 B.n260 B.n203 163.367
R1622 B.n260 B.n259 163.367
R1623 B.n259 B.n258 163.367
R1624 B.n258 B.n205 163.367
R1625 B.n254 B.n205 163.367
R1626 B.n254 B.n253 163.367
R1627 B.n253 B.n252 163.367
R1628 B.n252 B.n207 163.367
R1629 B.n248 B.n207 163.367
R1630 B.n248 B.n247 163.367
R1631 B.n247 B.n246 163.367
R1632 B.n246 B.n209 163.367
R1633 B.n242 B.n209 163.367
R1634 B.n242 B.n241 163.367
R1635 B.n241 B.n240 163.367
R1636 B.n240 B.n211 163.367
R1637 B.n236 B.n211 163.367
R1638 B.n236 B.n235 163.367
R1639 B.n235 B.n234 163.367
R1640 B.n234 B.n213 163.367
R1641 B.n230 B.n213 163.367
R1642 B.n230 B.n229 163.367
R1643 B.n229 B.n228 163.367
R1644 B.n228 B.n215 163.367
R1645 B.n224 B.n215 163.367
R1646 B.n224 B.n223 163.367
R1647 B.n223 B.n222 163.367
R1648 B.n222 B.n217 163.367
R1649 B.n218 B.n217 163.367
R1650 B.n218 B.n2 163.367
R1651 B.n842 B.n2 163.367
R1652 B.n842 B.n841 163.367
R1653 B.n841 B.n840 163.367
R1654 B.n840 B.n3 163.367
R1655 B.n836 B.n3 163.367
R1656 B.n836 B.n835 163.367
R1657 B.n835 B.n834 163.367
R1658 B.n834 B.n5 163.367
R1659 B.n830 B.n5 163.367
R1660 B.n830 B.n829 163.367
R1661 B.n829 B.n828 163.367
R1662 B.n828 B.n7 163.367
R1663 B.n824 B.n7 163.367
R1664 B.n824 B.n823 163.367
R1665 B.n823 B.n822 163.367
R1666 B.n822 B.n9 163.367
R1667 B.n818 B.n9 163.367
R1668 B.n818 B.n817 163.367
R1669 B.n817 B.n816 163.367
R1670 B.n816 B.n11 163.367
R1671 B.n812 B.n11 163.367
R1672 B.n812 B.n811 163.367
R1673 B.n811 B.n810 163.367
R1674 B.n810 B.n13 163.367
R1675 B.n806 B.n13 163.367
R1676 B.n806 B.n805 163.367
R1677 B.n805 B.n804 163.367
R1678 B.n804 B.n15 163.367
R1679 B.n800 B.n15 163.367
R1680 B.n800 B.n799 163.367
R1681 B.n799 B.n798 163.367
R1682 B.n798 B.n17 163.367
R1683 B.n794 B.n17 163.367
R1684 B.n794 B.n793 163.367
R1685 B.n793 B.n792 163.367
R1686 B.n792 B.n19 163.367
R1687 B.n788 B.n19 163.367
R1688 B.n788 B.n787 163.367
R1689 B.n787 B.n786 163.367
R1690 B.n786 B.n21 163.367
R1691 B.n782 B.n21 163.367
R1692 B.n782 B.n781 163.367
R1693 B.n781 B.n780 163.367
R1694 B.n780 B.n23 163.367
R1695 B.n776 B.n23 163.367
R1696 B.n776 B.n775 163.367
R1697 B.n775 B.n774 163.367
R1698 B.n774 B.n25 163.367
R1699 B.n289 B.n288 163.367
R1700 B.n290 B.n289 163.367
R1701 B.n290 B.n193 163.367
R1702 B.n294 B.n193 163.367
R1703 B.n295 B.n294 163.367
R1704 B.n296 B.n295 163.367
R1705 B.n296 B.n191 163.367
R1706 B.n300 B.n191 163.367
R1707 B.n301 B.n300 163.367
R1708 B.n302 B.n301 163.367
R1709 B.n302 B.n189 163.367
R1710 B.n306 B.n189 163.367
R1711 B.n307 B.n306 163.367
R1712 B.n308 B.n307 163.367
R1713 B.n308 B.n187 163.367
R1714 B.n312 B.n187 163.367
R1715 B.n313 B.n312 163.367
R1716 B.n314 B.n313 163.367
R1717 B.n314 B.n185 163.367
R1718 B.n318 B.n185 163.367
R1719 B.n319 B.n318 163.367
R1720 B.n320 B.n319 163.367
R1721 B.n320 B.n183 163.367
R1722 B.n324 B.n183 163.367
R1723 B.n325 B.n324 163.367
R1724 B.n326 B.n325 163.367
R1725 B.n326 B.n181 163.367
R1726 B.n330 B.n181 163.367
R1727 B.n331 B.n330 163.367
R1728 B.n332 B.n331 163.367
R1729 B.n332 B.n179 163.367
R1730 B.n336 B.n179 163.367
R1731 B.n337 B.n336 163.367
R1732 B.n338 B.n337 163.367
R1733 B.n338 B.n177 163.367
R1734 B.n342 B.n177 163.367
R1735 B.n343 B.n342 163.367
R1736 B.n344 B.n343 163.367
R1737 B.n344 B.n175 163.367
R1738 B.n348 B.n175 163.367
R1739 B.n349 B.n348 163.367
R1740 B.n350 B.n349 163.367
R1741 B.n350 B.n173 163.367
R1742 B.n354 B.n173 163.367
R1743 B.n355 B.n354 163.367
R1744 B.n356 B.n355 163.367
R1745 B.n356 B.n171 163.367
R1746 B.n360 B.n171 163.367
R1747 B.n361 B.n360 163.367
R1748 B.n362 B.n361 163.367
R1749 B.n362 B.n167 163.367
R1750 B.n367 B.n167 163.367
R1751 B.n368 B.n367 163.367
R1752 B.n369 B.n368 163.367
R1753 B.n369 B.n165 163.367
R1754 B.n373 B.n165 163.367
R1755 B.n374 B.n373 163.367
R1756 B.n375 B.n374 163.367
R1757 B.n375 B.n163 163.367
R1758 B.n379 B.n163 163.367
R1759 B.n380 B.n379 163.367
R1760 B.n380 B.n159 163.367
R1761 B.n384 B.n159 163.367
R1762 B.n385 B.n384 163.367
R1763 B.n386 B.n385 163.367
R1764 B.n386 B.n157 163.367
R1765 B.n390 B.n157 163.367
R1766 B.n391 B.n390 163.367
R1767 B.n392 B.n391 163.367
R1768 B.n392 B.n155 163.367
R1769 B.n396 B.n155 163.367
R1770 B.n397 B.n396 163.367
R1771 B.n398 B.n397 163.367
R1772 B.n398 B.n153 163.367
R1773 B.n402 B.n153 163.367
R1774 B.n403 B.n402 163.367
R1775 B.n404 B.n403 163.367
R1776 B.n404 B.n151 163.367
R1777 B.n408 B.n151 163.367
R1778 B.n409 B.n408 163.367
R1779 B.n410 B.n409 163.367
R1780 B.n410 B.n149 163.367
R1781 B.n414 B.n149 163.367
R1782 B.n415 B.n414 163.367
R1783 B.n416 B.n415 163.367
R1784 B.n416 B.n147 163.367
R1785 B.n420 B.n147 163.367
R1786 B.n421 B.n420 163.367
R1787 B.n422 B.n421 163.367
R1788 B.n422 B.n145 163.367
R1789 B.n426 B.n145 163.367
R1790 B.n427 B.n426 163.367
R1791 B.n428 B.n427 163.367
R1792 B.n428 B.n143 163.367
R1793 B.n432 B.n143 163.367
R1794 B.n433 B.n432 163.367
R1795 B.n434 B.n433 163.367
R1796 B.n434 B.n141 163.367
R1797 B.n438 B.n141 163.367
R1798 B.n439 B.n438 163.367
R1799 B.n440 B.n439 163.367
R1800 B.n440 B.n139 163.367
R1801 B.n444 B.n139 163.367
R1802 B.n445 B.n444 163.367
R1803 B.n446 B.n445 163.367
R1804 B.n446 B.n137 163.367
R1805 B.n450 B.n137 163.367
R1806 B.n451 B.n450 163.367
R1807 B.n452 B.n451 163.367
R1808 B.n452 B.n135 163.367
R1809 B.n456 B.n135 163.367
R1810 B.n457 B.n456 163.367
R1811 B.n458 B.n133 163.367
R1812 B.n462 B.n133 163.367
R1813 B.n463 B.n462 163.367
R1814 B.n464 B.n463 163.367
R1815 B.n464 B.n131 163.367
R1816 B.n468 B.n131 163.367
R1817 B.n469 B.n468 163.367
R1818 B.n470 B.n469 163.367
R1819 B.n470 B.n129 163.367
R1820 B.n474 B.n129 163.367
R1821 B.n475 B.n474 163.367
R1822 B.n476 B.n475 163.367
R1823 B.n476 B.n127 163.367
R1824 B.n480 B.n127 163.367
R1825 B.n481 B.n480 163.367
R1826 B.n482 B.n481 163.367
R1827 B.n482 B.n125 163.367
R1828 B.n486 B.n125 163.367
R1829 B.n487 B.n486 163.367
R1830 B.n488 B.n487 163.367
R1831 B.n488 B.n123 163.367
R1832 B.n492 B.n123 163.367
R1833 B.n493 B.n492 163.367
R1834 B.n494 B.n493 163.367
R1835 B.n494 B.n121 163.367
R1836 B.n498 B.n121 163.367
R1837 B.n499 B.n498 163.367
R1838 B.n500 B.n499 163.367
R1839 B.n500 B.n119 163.367
R1840 B.n504 B.n119 163.367
R1841 B.n505 B.n504 163.367
R1842 B.n506 B.n505 163.367
R1843 B.n506 B.n117 163.367
R1844 B.n510 B.n117 163.367
R1845 B.n511 B.n510 163.367
R1846 B.n512 B.n511 163.367
R1847 B.n512 B.n115 163.367
R1848 B.n516 B.n115 163.367
R1849 B.n517 B.n516 163.367
R1850 B.n518 B.n517 163.367
R1851 B.n518 B.n113 163.367
R1852 B.n522 B.n113 163.367
R1853 B.n523 B.n522 163.367
R1854 B.n524 B.n523 163.367
R1855 B.n524 B.n111 163.367
R1856 B.n528 B.n111 163.367
R1857 B.n529 B.n528 163.367
R1858 B.n530 B.n529 163.367
R1859 B.n530 B.n109 163.367
R1860 B.n534 B.n109 163.367
R1861 B.n535 B.n534 163.367
R1862 B.n536 B.n535 163.367
R1863 B.n536 B.n107 163.367
R1864 B.n540 B.n107 163.367
R1865 B.n541 B.n540 163.367
R1866 B.n542 B.n541 163.367
R1867 B.n542 B.n105 163.367
R1868 B.n546 B.n105 163.367
R1869 B.n547 B.n546 163.367
R1870 B.n548 B.n547 163.367
R1871 B.n548 B.n103 163.367
R1872 B.n552 B.n103 163.367
R1873 B.n553 B.n552 163.367
R1874 B.n554 B.n553 163.367
R1875 B.n554 B.n101 163.367
R1876 B.n558 B.n101 163.367
R1877 B.n559 B.n558 163.367
R1878 B.n560 B.n559 163.367
R1879 B.n560 B.n99 163.367
R1880 B.n564 B.n99 163.367
R1881 B.n565 B.n564 163.367
R1882 B.n566 B.n565 163.367
R1883 B.n566 B.n97 163.367
R1884 B.n570 B.n97 163.367
R1885 B.n571 B.n570 163.367
R1886 B.n572 B.n571 163.367
R1887 B.n572 B.n95 163.367
R1888 B.n576 B.n95 163.367
R1889 B.n577 B.n576 163.367
R1890 B.n578 B.n577 163.367
R1891 B.n578 B.n93 163.367
R1892 B.n582 B.n93 163.367
R1893 B.n583 B.n582 163.367
R1894 B.n584 B.n583 163.367
R1895 B.n584 B.n91 163.367
R1896 B.n588 B.n91 163.367
R1897 B.n589 B.n588 163.367
R1898 B.n590 B.n589 163.367
R1899 B.n590 B.n89 163.367
R1900 B.n594 B.n89 163.367
R1901 B.n595 B.n594 163.367
R1902 B.n596 B.n595 163.367
R1903 B.n596 B.n87 163.367
R1904 B.n600 B.n87 163.367
R1905 B.n770 B.n769 163.367
R1906 B.n769 B.n768 163.367
R1907 B.n768 B.n27 163.367
R1908 B.n764 B.n27 163.367
R1909 B.n764 B.n763 163.367
R1910 B.n763 B.n762 163.367
R1911 B.n762 B.n29 163.367
R1912 B.n758 B.n29 163.367
R1913 B.n758 B.n757 163.367
R1914 B.n757 B.n756 163.367
R1915 B.n756 B.n31 163.367
R1916 B.n752 B.n31 163.367
R1917 B.n752 B.n751 163.367
R1918 B.n751 B.n750 163.367
R1919 B.n750 B.n33 163.367
R1920 B.n746 B.n33 163.367
R1921 B.n746 B.n745 163.367
R1922 B.n745 B.n744 163.367
R1923 B.n744 B.n35 163.367
R1924 B.n740 B.n35 163.367
R1925 B.n740 B.n739 163.367
R1926 B.n739 B.n738 163.367
R1927 B.n738 B.n37 163.367
R1928 B.n734 B.n37 163.367
R1929 B.n734 B.n733 163.367
R1930 B.n733 B.n732 163.367
R1931 B.n732 B.n39 163.367
R1932 B.n728 B.n39 163.367
R1933 B.n728 B.n727 163.367
R1934 B.n727 B.n726 163.367
R1935 B.n726 B.n41 163.367
R1936 B.n722 B.n41 163.367
R1937 B.n722 B.n721 163.367
R1938 B.n721 B.n720 163.367
R1939 B.n720 B.n43 163.367
R1940 B.n716 B.n43 163.367
R1941 B.n716 B.n715 163.367
R1942 B.n715 B.n714 163.367
R1943 B.n714 B.n45 163.367
R1944 B.n710 B.n45 163.367
R1945 B.n710 B.n709 163.367
R1946 B.n709 B.n708 163.367
R1947 B.n708 B.n47 163.367
R1948 B.n704 B.n47 163.367
R1949 B.n704 B.n703 163.367
R1950 B.n703 B.n702 163.367
R1951 B.n702 B.n49 163.367
R1952 B.n698 B.n49 163.367
R1953 B.n698 B.n697 163.367
R1954 B.n697 B.n696 163.367
R1955 B.n696 B.n51 163.367
R1956 B.n691 B.n51 163.367
R1957 B.n691 B.n690 163.367
R1958 B.n690 B.n689 163.367
R1959 B.n689 B.n55 163.367
R1960 B.n685 B.n55 163.367
R1961 B.n685 B.n684 163.367
R1962 B.n684 B.n683 163.367
R1963 B.n683 B.n57 163.367
R1964 B.n679 B.n57 163.367
R1965 B.n679 B.n678 163.367
R1966 B.n678 B.n61 163.367
R1967 B.n674 B.n61 163.367
R1968 B.n674 B.n673 163.367
R1969 B.n673 B.n672 163.367
R1970 B.n672 B.n63 163.367
R1971 B.n668 B.n63 163.367
R1972 B.n668 B.n667 163.367
R1973 B.n667 B.n666 163.367
R1974 B.n666 B.n65 163.367
R1975 B.n662 B.n65 163.367
R1976 B.n662 B.n661 163.367
R1977 B.n661 B.n660 163.367
R1978 B.n660 B.n67 163.367
R1979 B.n656 B.n67 163.367
R1980 B.n656 B.n655 163.367
R1981 B.n655 B.n654 163.367
R1982 B.n654 B.n69 163.367
R1983 B.n650 B.n69 163.367
R1984 B.n650 B.n649 163.367
R1985 B.n649 B.n648 163.367
R1986 B.n648 B.n71 163.367
R1987 B.n644 B.n71 163.367
R1988 B.n644 B.n643 163.367
R1989 B.n643 B.n642 163.367
R1990 B.n642 B.n73 163.367
R1991 B.n638 B.n73 163.367
R1992 B.n638 B.n637 163.367
R1993 B.n637 B.n636 163.367
R1994 B.n636 B.n75 163.367
R1995 B.n632 B.n75 163.367
R1996 B.n632 B.n631 163.367
R1997 B.n631 B.n630 163.367
R1998 B.n630 B.n77 163.367
R1999 B.n626 B.n77 163.367
R2000 B.n626 B.n625 163.367
R2001 B.n625 B.n624 163.367
R2002 B.n624 B.n79 163.367
R2003 B.n620 B.n79 163.367
R2004 B.n620 B.n619 163.367
R2005 B.n619 B.n618 163.367
R2006 B.n618 B.n81 163.367
R2007 B.n614 B.n81 163.367
R2008 B.n614 B.n613 163.367
R2009 B.n613 B.n612 163.367
R2010 B.n612 B.n83 163.367
R2011 B.n608 B.n83 163.367
R2012 B.n608 B.n607 163.367
R2013 B.n607 B.n606 163.367
R2014 B.n606 B.n85 163.367
R2015 B.n602 B.n85 163.367
R2016 B.n602 B.n601 163.367
R2017 B.n162 B.n161 59.5399
R2018 B.n365 B.n169 59.5399
R2019 B.n693 B.n53 59.5399
R2020 B.n60 B.n59 59.5399
R2021 B.n161 B.n160 51.0066
R2022 B.n169 B.n168 51.0066
R2023 B.n53 B.n52 51.0066
R2024 B.n59 B.n58 51.0066
R2025 B.n772 B.n771 29.1907
R2026 B.n459 B.n134 29.1907
R2027 B.n287 B.n286 29.1907
R2028 B.n599 B.n86 29.1907
R2029 B B.n843 18.0485
R2030 B.n771 B.n26 10.6151
R2031 B.n767 B.n26 10.6151
R2032 B.n767 B.n766 10.6151
R2033 B.n766 B.n765 10.6151
R2034 B.n765 B.n28 10.6151
R2035 B.n761 B.n28 10.6151
R2036 B.n761 B.n760 10.6151
R2037 B.n760 B.n759 10.6151
R2038 B.n759 B.n30 10.6151
R2039 B.n755 B.n30 10.6151
R2040 B.n755 B.n754 10.6151
R2041 B.n754 B.n753 10.6151
R2042 B.n753 B.n32 10.6151
R2043 B.n749 B.n32 10.6151
R2044 B.n749 B.n748 10.6151
R2045 B.n748 B.n747 10.6151
R2046 B.n747 B.n34 10.6151
R2047 B.n743 B.n34 10.6151
R2048 B.n743 B.n742 10.6151
R2049 B.n742 B.n741 10.6151
R2050 B.n741 B.n36 10.6151
R2051 B.n737 B.n36 10.6151
R2052 B.n737 B.n736 10.6151
R2053 B.n736 B.n735 10.6151
R2054 B.n735 B.n38 10.6151
R2055 B.n731 B.n38 10.6151
R2056 B.n731 B.n730 10.6151
R2057 B.n730 B.n729 10.6151
R2058 B.n729 B.n40 10.6151
R2059 B.n725 B.n40 10.6151
R2060 B.n725 B.n724 10.6151
R2061 B.n724 B.n723 10.6151
R2062 B.n723 B.n42 10.6151
R2063 B.n719 B.n42 10.6151
R2064 B.n719 B.n718 10.6151
R2065 B.n718 B.n717 10.6151
R2066 B.n717 B.n44 10.6151
R2067 B.n713 B.n44 10.6151
R2068 B.n713 B.n712 10.6151
R2069 B.n712 B.n711 10.6151
R2070 B.n711 B.n46 10.6151
R2071 B.n707 B.n46 10.6151
R2072 B.n707 B.n706 10.6151
R2073 B.n706 B.n705 10.6151
R2074 B.n705 B.n48 10.6151
R2075 B.n701 B.n48 10.6151
R2076 B.n701 B.n700 10.6151
R2077 B.n700 B.n699 10.6151
R2078 B.n699 B.n50 10.6151
R2079 B.n695 B.n50 10.6151
R2080 B.n695 B.n694 10.6151
R2081 B.n692 B.n54 10.6151
R2082 B.n688 B.n54 10.6151
R2083 B.n688 B.n687 10.6151
R2084 B.n687 B.n686 10.6151
R2085 B.n686 B.n56 10.6151
R2086 B.n682 B.n56 10.6151
R2087 B.n682 B.n681 10.6151
R2088 B.n681 B.n680 10.6151
R2089 B.n677 B.n676 10.6151
R2090 B.n676 B.n675 10.6151
R2091 B.n675 B.n62 10.6151
R2092 B.n671 B.n62 10.6151
R2093 B.n671 B.n670 10.6151
R2094 B.n670 B.n669 10.6151
R2095 B.n669 B.n64 10.6151
R2096 B.n665 B.n64 10.6151
R2097 B.n665 B.n664 10.6151
R2098 B.n664 B.n663 10.6151
R2099 B.n663 B.n66 10.6151
R2100 B.n659 B.n66 10.6151
R2101 B.n659 B.n658 10.6151
R2102 B.n658 B.n657 10.6151
R2103 B.n657 B.n68 10.6151
R2104 B.n653 B.n68 10.6151
R2105 B.n653 B.n652 10.6151
R2106 B.n652 B.n651 10.6151
R2107 B.n651 B.n70 10.6151
R2108 B.n647 B.n70 10.6151
R2109 B.n647 B.n646 10.6151
R2110 B.n646 B.n645 10.6151
R2111 B.n645 B.n72 10.6151
R2112 B.n641 B.n72 10.6151
R2113 B.n641 B.n640 10.6151
R2114 B.n640 B.n639 10.6151
R2115 B.n639 B.n74 10.6151
R2116 B.n635 B.n74 10.6151
R2117 B.n635 B.n634 10.6151
R2118 B.n634 B.n633 10.6151
R2119 B.n633 B.n76 10.6151
R2120 B.n629 B.n76 10.6151
R2121 B.n629 B.n628 10.6151
R2122 B.n628 B.n627 10.6151
R2123 B.n627 B.n78 10.6151
R2124 B.n623 B.n78 10.6151
R2125 B.n623 B.n622 10.6151
R2126 B.n622 B.n621 10.6151
R2127 B.n621 B.n80 10.6151
R2128 B.n617 B.n80 10.6151
R2129 B.n617 B.n616 10.6151
R2130 B.n616 B.n615 10.6151
R2131 B.n615 B.n82 10.6151
R2132 B.n611 B.n82 10.6151
R2133 B.n611 B.n610 10.6151
R2134 B.n610 B.n609 10.6151
R2135 B.n609 B.n84 10.6151
R2136 B.n605 B.n84 10.6151
R2137 B.n605 B.n604 10.6151
R2138 B.n604 B.n603 10.6151
R2139 B.n603 B.n86 10.6151
R2140 B.n460 B.n459 10.6151
R2141 B.n461 B.n460 10.6151
R2142 B.n461 B.n132 10.6151
R2143 B.n465 B.n132 10.6151
R2144 B.n466 B.n465 10.6151
R2145 B.n467 B.n466 10.6151
R2146 B.n467 B.n130 10.6151
R2147 B.n471 B.n130 10.6151
R2148 B.n472 B.n471 10.6151
R2149 B.n473 B.n472 10.6151
R2150 B.n473 B.n128 10.6151
R2151 B.n477 B.n128 10.6151
R2152 B.n478 B.n477 10.6151
R2153 B.n479 B.n478 10.6151
R2154 B.n479 B.n126 10.6151
R2155 B.n483 B.n126 10.6151
R2156 B.n484 B.n483 10.6151
R2157 B.n485 B.n484 10.6151
R2158 B.n485 B.n124 10.6151
R2159 B.n489 B.n124 10.6151
R2160 B.n490 B.n489 10.6151
R2161 B.n491 B.n490 10.6151
R2162 B.n491 B.n122 10.6151
R2163 B.n495 B.n122 10.6151
R2164 B.n496 B.n495 10.6151
R2165 B.n497 B.n496 10.6151
R2166 B.n497 B.n120 10.6151
R2167 B.n501 B.n120 10.6151
R2168 B.n502 B.n501 10.6151
R2169 B.n503 B.n502 10.6151
R2170 B.n503 B.n118 10.6151
R2171 B.n507 B.n118 10.6151
R2172 B.n508 B.n507 10.6151
R2173 B.n509 B.n508 10.6151
R2174 B.n509 B.n116 10.6151
R2175 B.n513 B.n116 10.6151
R2176 B.n514 B.n513 10.6151
R2177 B.n515 B.n514 10.6151
R2178 B.n515 B.n114 10.6151
R2179 B.n519 B.n114 10.6151
R2180 B.n520 B.n519 10.6151
R2181 B.n521 B.n520 10.6151
R2182 B.n521 B.n112 10.6151
R2183 B.n525 B.n112 10.6151
R2184 B.n526 B.n525 10.6151
R2185 B.n527 B.n526 10.6151
R2186 B.n527 B.n110 10.6151
R2187 B.n531 B.n110 10.6151
R2188 B.n532 B.n531 10.6151
R2189 B.n533 B.n532 10.6151
R2190 B.n533 B.n108 10.6151
R2191 B.n537 B.n108 10.6151
R2192 B.n538 B.n537 10.6151
R2193 B.n539 B.n538 10.6151
R2194 B.n539 B.n106 10.6151
R2195 B.n543 B.n106 10.6151
R2196 B.n544 B.n543 10.6151
R2197 B.n545 B.n544 10.6151
R2198 B.n545 B.n104 10.6151
R2199 B.n549 B.n104 10.6151
R2200 B.n550 B.n549 10.6151
R2201 B.n551 B.n550 10.6151
R2202 B.n551 B.n102 10.6151
R2203 B.n555 B.n102 10.6151
R2204 B.n556 B.n555 10.6151
R2205 B.n557 B.n556 10.6151
R2206 B.n557 B.n100 10.6151
R2207 B.n561 B.n100 10.6151
R2208 B.n562 B.n561 10.6151
R2209 B.n563 B.n562 10.6151
R2210 B.n563 B.n98 10.6151
R2211 B.n567 B.n98 10.6151
R2212 B.n568 B.n567 10.6151
R2213 B.n569 B.n568 10.6151
R2214 B.n569 B.n96 10.6151
R2215 B.n573 B.n96 10.6151
R2216 B.n574 B.n573 10.6151
R2217 B.n575 B.n574 10.6151
R2218 B.n575 B.n94 10.6151
R2219 B.n579 B.n94 10.6151
R2220 B.n580 B.n579 10.6151
R2221 B.n581 B.n580 10.6151
R2222 B.n581 B.n92 10.6151
R2223 B.n585 B.n92 10.6151
R2224 B.n586 B.n585 10.6151
R2225 B.n587 B.n586 10.6151
R2226 B.n587 B.n90 10.6151
R2227 B.n591 B.n90 10.6151
R2228 B.n592 B.n591 10.6151
R2229 B.n593 B.n592 10.6151
R2230 B.n593 B.n88 10.6151
R2231 B.n597 B.n88 10.6151
R2232 B.n598 B.n597 10.6151
R2233 B.n599 B.n598 10.6151
R2234 B.n287 B.n194 10.6151
R2235 B.n291 B.n194 10.6151
R2236 B.n292 B.n291 10.6151
R2237 B.n293 B.n292 10.6151
R2238 B.n293 B.n192 10.6151
R2239 B.n297 B.n192 10.6151
R2240 B.n298 B.n297 10.6151
R2241 B.n299 B.n298 10.6151
R2242 B.n299 B.n190 10.6151
R2243 B.n303 B.n190 10.6151
R2244 B.n304 B.n303 10.6151
R2245 B.n305 B.n304 10.6151
R2246 B.n305 B.n188 10.6151
R2247 B.n309 B.n188 10.6151
R2248 B.n310 B.n309 10.6151
R2249 B.n311 B.n310 10.6151
R2250 B.n311 B.n186 10.6151
R2251 B.n315 B.n186 10.6151
R2252 B.n316 B.n315 10.6151
R2253 B.n317 B.n316 10.6151
R2254 B.n317 B.n184 10.6151
R2255 B.n321 B.n184 10.6151
R2256 B.n322 B.n321 10.6151
R2257 B.n323 B.n322 10.6151
R2258 B.n323 B.n182 10.6151
R2259 B.n327 B.n182 10.6151
R2260 B.n328 B.n327 10.6151
R2261 B.n329 B.n328 10.6151
R2262 B.n329 B.n180 10.6151
R2263 B.n333 B.n180 10.6151
R2264 B.n334 B.n333 10.6151
R2265 B.n335 B.n334 10.6151
R2266 B.n335 B.n178 10.6151
R2267 B.n339 B.n178 10.6151
R2268 B.n340 B.n339 10.6151
R2269 B.n341 B.n340 10.6151
R2270 B.n341 B.n176 10.6151
R2271 B.n345 B.n176 10.6151
R2272 B.n346 B.n345 10.6151
R2273 B.n347 B.n346 10.6151
R2274 B.n347 B.n174 10.6151
R2275 B.n351 B.n174 10.6151
R2276 B.n352 B.n351 10.6151
R2277 B.n353 B.n352 10.6151
R2278 B.n353 B.n172 10.6151
R2279 B.n357 B.n172 10.6151
R2280 B.n358 B.n357 10.6151
R2281 B.n359 B.n358 10.6151
R2282 B.n359 B.n170 10.6151
R2283 B.n363 B.n170 10.6151
R2284 B.n364 B.n363 10.6151
R2285 B.n366 B.n166 10.6151
R2286 B.n370 B.n166 10.6151
R2287 B.n371 B.n370 10.6151
R2288 B.n372 B.n371 10.6151
R2289 B.n372 B.n164 10.6151
R2290 B.n376 B.n164 10.6151
R2291 B.n377 B.n376 10.6151
R2292 B.n378 B.n377 10.6151
R2293 B.n382 B.n381 10.6151
R2294 B.n383 B.n382 10.6151
R2295 B.n383 B.n158 10.6151
R2296 B.n387 B.n158 10.6151
R2297 B.n388 B.n387 10.6151
R2298 B.n389 B.n388 10.6151
R2299 B.n389 B.n156 10.6151
R2300 B.n393 B.n156 10.6151
R2301 B.n394 B.n393 10.6151
R2302 B.n395 B.n394 10.6151
R2303 B.n395 B.n154 10.6151
R2304 B.n399 B.n154 10.6151
R2305 B.n400 B.n399 10.6151
R2306 B.n401 B.n400 10.6151
R2307 B.n401 B.n152 10.6151
R2308 B.n405 B.n152 10.6151
R2309 B.n406 B.n405 10.6151
R2310 B.n407 B.n406 10.6151
R2311 B.n407 B.n150 10.6151
R2312 B.n411 B.n150 10.6151
R2313 B.n412 B.n411 10.6151
R2314 B.n413 B.n412 10.6151
R2315 B.n413 B.n148 10.6151
R2316 B.n417 B.n148 10.6151
R2317 B.n418 B.n417 10.6151
R2318 B.n419 B.n418 10.6151
R2319 B.n419 B.n146 10.6151
R2320 B.n423 B.n146 10.6151
R2321 B.n424 B.n423 10.6151
R2322 B.n425 B.n424 10.6151
R2323 B.n425 B.n144 10.6151
R2324 B.n429 B.n144 10.6151
R2325 B.n430 B.n429 10.6151
R2326 B.n431 B.n430 10.6151
R2327 B.n431 B.n142 10.6151
R2328 B.n435 B.n142 10.6151
R2329 B.n436 B.n435 10.6151
R2330 B.n437 B.n436 10.6151
R2331 B.n437 B.n140 10.6151
R2332 B.n441 B.n140 10.6151
R2333 B.n442 B.n441 10.6151
R2334 B.n443 B.n442 10.6151
R2335 B.n443 B.n138 10.6151
R2336 B.n447 B.n138 10.6151
R2337 B.n448 B.n447 10.6151
R2338 B.n449 B.n448 10.6151
R2339 B.n449 B.n136 10.6151
R2340 B.n453 B.n136 10.6151
R2341 B.n454 B.n453 10.6151
R2342 B.n455 B.n454 10.6151
R2343 B.n455 B.n134 10.6151
R2344 B.n286 B.n285 10.6151
R2345 B.n285 B.n196 10.6151
R2346 B.n281 B.n196 10.6151
R2347 B.n281 B.n280 10.6151
R2348 B.n280 B.n279 10.6151
R2349 B.n279 B.n198 10.6151
R2350 B.n275 B.n198 10.6151
R2351 B.n275 B.n274 10.6151
R2352 B.n274 B.n273 10.6151
R2353 B.n273 B.n200 10.6151
R2354 B.n269 B.n200 10.6151
R2355 B.n269 B.n268 10.6151
R2356 B.n268 B.n267 10.6151
R2357 B.n267 B.n202 10.6151
R2358 B.n263 B.n202 10.6151
R2359 B.n263 B.n262 10.6151
R2360 B.n262 B.n261 10.6151
R2361 B.n261 B.n204 10.6151
R2362 B.n257 B.n204 10.6151
R2363 B.n257 B.n256 10.6151
R2364 B.n256 B.n255 10.6151
R2365 B.n255 B.n206 10.6151
R2366 B.n251 B.n206 10.6151
R2367 B.n251 B.n250 10.6151
R2368 B.n250 B.n249 10.6151
R2369 B.n249 B.n208 10.6151
R2370 B.n245 B.n208 10.6151
R2371 B.n245 B.n244 10.6151
R2372 B.n244 B.n243 10.6151
R2373 B.n243 B.n210 10.6151
R2374 B.n239 B.n210 10.6151
R2375 B.n239 B.n238 10.6151
R2376 B.n238 B.n237 10.6151
R2377 B.n237 B.n212 10.6151
R2378 B.n233 B.n212 10.6151
R2379 B.n233 B.n232 10.6151
R2380 B.n232 B.n231 10.6151
R2381 B.n231 B.n214 10.6151
R2382 B.n227 B.n214 10.6151
R2383 B.n227 B.n226 10.6151
R2384 B.n226 B.n225 10.6151
R2385 B.n225 B.n216 10.6151
R2386 B.n221 B.n216 10.6151
R2387 B.n221 B.n220 10.6151
R2388 B.n220 B.n219 10.6151
R2389 B.n219 B.n0 10.6151
R2390 B.n839 B.n1 10.6151
R2391 B.n839 B.n838 10.6151
R2392 B.n838 B.n837 10.6151
R2393 B.n837 B.n4 10.6151
R2394 B.n833 B.n4 10.6151
R2395 B.n833 B.n832 10.6151
R2396 B.n832 B.n831 10.6151
R2397 B.n831 B.n6 10.6151
R2398 B.n827 B.n6 10.6151
R2399 B.n827 B.n826 10.6151
R2400 B.n826 B.n825 10.6151
R2401 B.n825 B.n8 10.6151
R2402 B.n821 B.n8 10.6151
R2403 B.n821 B.n820 10.6151
R2404 B.n820 B.n819 10.6151
R2405 B.n819 B.n10 10.6151
R2406 B.n815 B.n10 10.6151
R2407 B.n815 B.n814 10.6151
R2408 B.n814 B.n813 10.6151
R2409 B.n813 B.n12 10.6151
R2410 B.n809 B.n12 10.6151
R2411 B.n809 B.n808 10.6151
R2412 B.n808 B.n807 10.6151
R2413 B.n807 B.n14 10.6151
R2414 B.n803 B.n14 10.6151
R2415 B.n803 B.n802 10.6151
R2416 B.n802 B.n801 10.6151
R2417 B.n801 B.n16 10.6151
R2418 B.n797 B.n16 10.6151
R2419 B.n797 B.n796 10.6151
R2420 B.n796 B.n795 10.6151
R2421 B.n795 B.n18 10.6151
R2422 B.n791 B.n18 10.6151
R2423 B.n791 B.n790 10.6151
R2424 B.n790 B.n789 10.6151
R2425 B.n789 B.n20 10.6151
R2426 B.n785 B.n20 10.6151
R2427 B.n785 B.n784 10.6151
R2428 B.n784 B.n783 10.6151
R2429 B.n783 B.n22 10.6151
R2430 B.n779 B.n22 10.6151
R2431 B.n779 B.n778 10.6151
R2432 B.n778 B.n777 10.6151
R2433 B.n777 B.n24 10.6151
R2434 B.n773 B.n24 10.6151
R2435 B.n773 B.n772 10.6151
R2436 B.n693 B.n692 6.5566
R2437 B.n680 B.n60 6.5566
R2438 B.n366 B.n365 6.5566
R2439 B.n378 B.n162 6.5566
R2440 B.n694 B.n693 4.05904
R2441 B.n677 B.n60 4.05904
R2442 B.n365 B.n364 4.05904
R2443 B.n381 B.n162 4.05904
R2444 B.n843 B.n0 2.81026
R2445 B.n843 B.n1 2.81026
R2446 VN.n7 VN.t7 192.149
R2447 VN.n34 VN.t3 192.149
R2448 VN.n6 VN.t1 161.365
R2449 VN.n17 VN.t0 161.365
R2450 VN.n25 VN.t2 161.365
R2451 VN.n33 VN.t4 161.365
R2452 VN.n44 VN.t5 161.365
R2453 VN.n52 VN.t6 161.365
R2454 VN.n51 VN.n27 161.3
R2455 VN.n50 VN.n49 161.3
R2456 VN.n48 VN.n28 161.3
R2457 VN.n47 VN.n46 161.3
R2458 VN.n45 VN.n29 161.3
R2459 VN.n43 VN.n42 161.3
R2460 VN.n41 VN.n30 161.3
R2461 VN.n40 VN.n39 161.3
R2462 VN.n38 VN.n31 161.3
R2463 VN.n37 VN.n36 161.3
R2464 VN.n35 VN.n32 161.3
R2465 VN.n24 VN.n0 161.3
R2466 VN.n23 VN.n22 161.3
R2467 VN.n21 VN.n1 161.3
R2468 VN.n20 VN.n19 161.3
R2469 VN.n18 VN.n2 161.3
R2470 VN.n16 VN.n15 161.3
R2471 VN.n14 VN.n3 161.3
R2472 VN.n13 VN.n12 161.3
R2473 VN.n11 VN.n4 161.3
R2474 VN.n10 VN.n9 161.3
R2475 VN.n8 VN.n5 161.3
R2476 VN.n26 VN.n25 101.317
R2477 VN.n53 VN.n52 101.317
R2478 VN.n7 VN.n6 69.2325
R2479 VN.n34 VN.n33 69.2325
R2480 VN.n12 VN.n11 56.5617
R2481 VN.n39 VN.n38 56.5617
R2482 VN VN.n53 52.2861
R2483 VN.n19 VN.n1 52.2023
R2484 VN.n46 VN.n28 52.2023
R2485 VN.n23 VN.n1 28.9518
R2486 VN.n50 VN.n28 28.9518
R2487 VN.n10 VN.n5 24.5923
R2488 VN.n11 VN.n10 24.5923
R2489 VN.n12 VN.n3 24.5923
R2490 VN.n16 VN.n3 24.5923
R2491 VN.n19 VN.n18 24.5923
R2492 VN.n24 VN.n23 24.5923
R2493 VN.n38 VN.n37 24.5923
R2494 VN.n37 VN.n32 24.5923
R2495 VN.n46 VN.n45 24.5923
R2496 VN.n43 VN.n30 24.5923
R2497 VN.n39 VN.n30 24.5923
R2498 VN.n51 VN.n50 24.5923
R2499 VN.n18 VN.n17 21.3954
R2500 VN.n45 VN.n44 21.3954
R2501 VN.n35 VN.n34 10.0465
R2502 VN.n8 VN.n7 10.0465
R2503 VN.n25 VN.n24 9.59132
R2504 VN.n52 VN.n51 9.59132
R2505 VN.n6 VN.n5 3.19744
R2506 VN.n17 VN.n16 3.19744
R2507 VN.n33 VN.n32 3.19744
R2508 VN.n44 VN.n43 3.19744
R2509 VN.n53 VN.n27 0.278335
R2510 VN.n26 VN.n0 0.278335
R2511 VN.n49 VN.n27 0.189894
R2512 VN.n49 VN.n48 0.189894
R2513 VN.n48 VN.n47 0.189894
R2514 VN.n47 VN.n29 0.189894
R2515 VN.n42 VN.n29 0.189894
R2516 VN.n42 VN.n41 0.189894
R2517 VN.n41 VN.n40 0.189894
R2518 VN.n40 VN.n31 0.189894
R2519 VN.n36 VN.n31 0.189894
R2520 VN.n36 VN.n35 0.189894
R2521 VN.n9 VN.n8 0.189894
R2522 VN.n9 VN.n4 0.189894
R2523 VN.n13 VN.n4 0.189894
R2524 VN.n14 VN.n13 0.189894
R2525 VN.n15 VN.n14 0.189894
R2526 VN.n15 VN.n2 0.189894
R2527 VN.n20 VN.n2 0.189894
R2528 VN.n21 VN.n20 0.189894
R2529 VN.n22 VN.n21 0.189894
R2530 VN.n22 VN.n0 0.189894
R2531 VN VN.n26 0.153485
R2532 VDD2.n2 VDD2.n1 72.112
R2533 VDD2.n2 VDD2.n0 72.112
R2534 VDD2 VDD2.n5 72.1092
R2535 VDD2.n4 VDD2.n3 71.0339
R2536 VDD2.n4 VDD2.n2 47.1937
R2537 VDD2.n5 VDD2.t3 2.11121
R2538 VDD2.n5 VDD2.t4 2.11121
R2539 VDD2.n3 VDD2.t1 2.11121
R2540 VDD2.n3 VDD2.t2 2.11121
R2541 VDD2.n1 VDD2.t7 2.11121
R2542 VDD2.n1 VDD2.t5 2.11121
R2543 VDD2.n0 VDD2.t0 2.11121
R2544 VDD2.n0 VDD2.t6 2.11121
R2545 VDD2 VDD2.n4 1.19231
C0 B VP 1.97925f
C1 VP VN 7.92368f
C2 VP VDD1 11.0871f
C3 w_n3600_n4048# B 10.6097f
C4 VP VDD2 0.487999f
C5 VP VTAIL 10.914401f
C6 w_n3600_n4048# VN 7.30487f
C7 B VN 1.19889f
C8 w_n3600_n4048# VDD1 1.94776f
C9 B VDD1 1.65068f
C10 VDD1 VN 0.151437f
C11 w_n3600_n4048# VDD2 2.04989f
C12 w_n3600_n4048# VTAIL 4.96573f
C13 B VDD2 1.73727f
C14 B VTAIL 5.93633f
C15 VDD2 VN 10.7517f
C16 VN VTAIL 10.9003f
C17 VDD1 VDD2 1.6207f
C18 VDD1 VTAIL 9.27602f
C19 VDD2 VTAIL 9.32843f
C20 w_n3600_n4048# VP 7.77135f
C21 VDD2 VSUBS 1.887643f
C22 VDD1 VSUBS 2.392503f
C23 VTAIL VSUBS 1.440321f
C24 VN VSUBS 6.49611f
C25 VP VSUBS 3.400721f
C26 B VSUBS 4.951468f
C27 w_n3600_n4048# VSUBS 0.178632p
C28 VDD2.t0 VSUBS 0.327171f
C29 VDD2.t6 VSUBS 0.327171f
C30 VDD2.n0 VSUBS 2.67912f
C31 VDD2.t7 VSUBS 0.327171f
C32 VDD2.t5 VSUBS 0.327171f
C33 VDD2.n1 VSUBS 2.67912f
C34 VDD2.n2 VSUBS 4.14726f
C35 VDD2.t1 VSUBS 0.327171f
C36 VDD2.t2 VSUBS 0.327171f
C37 VDD2.n3 VSUBS 2.66694f
C38 VDD2.n4 VSUBS 3.6319f
C39 VDD2.t3 VSUBS 0.327171f
C40 VDD2.t4 VSUBS 0.327171f
C41 VDD2.n5 VSUBS 2.67908f
C42 VN.n0 VSUBS 0.038384f
C43 VN.t2 VSUBS 2.8276f
C44 VN.n1 VSUBS 0.029339f
C45 VN.n2 VSUBS 0.029116f
C46 VN.t0 VSUBS 2.8276f
C47 VN.n3 VSUBS 0.053993f
C48 VN.n4 VSUBS 0.029116f
C49 VN.n5 VSUBS 0.030803f
C50 VN.t7 VSUBS 3.01119f
C51 VN.t1 VSUBS 2.8276f
C52 VN.n6 VSUBS 1.05861f
C53 VN.n7 VSUBS 1.05856f
C54 VN.n8 VSUBS 0.250278f
C55 VN.n9 VSUBS 0.029116f
C56 VN.n10 VSUBS 0.053993f
C57 VN.n11 VSUBS 0.042325f
C58 VN.n12 VSUBS 0.042325f
C59 VN.n13 VSUBS 0.029116f
C60 VN.n14 VSUBS 0.029116f
C61 VN.n15 VSUBS 0.029116f
C62 VN.n16 VSUBS 0.030803f
C63 VN.n17 VSUBS 0.99004f
C64 VN.n18 VSUBS 0.050528f
C65 VN.n19 VSUBS 0.052019f
C66 VN.n20 VSUBS 0.029116f
C67 VN.n21 VSUBS 0.029116f
C68 VN.n22 VSUBS 0.029116f
C69 VN.n23 VSUBS 0.057284f
C70 VN.n24 VSUBS 0.037734f
C71 VN.n25 VSUBS 1.07458f
C72 VN.n26 VSUBS 0.044918f
C73 VN.n27 VSUBS 0.038384f
C74 VN.t6 VSUBS 2.8276f
C75 VN.n28 VSUBS 0.029339f
C76 VN.n29 VSUBS 0.029116f
C77 VN.t5 VSUBS 2.8276f
C78 VN.n30 VSUBS 0.053993f
C79 VN.n31 VSUBS 0.029116f
C80 VN.n32 VSUBS 0.030803f
C81 VN.t3 VSUBS 3.01119f
C82 VN.t4 VSUBS 2.8276f
C83 VN.n33 VSUBS 1.05861f
C84 VN.n34 VSUBS 1.05856f
C85 VN.n35 VSUBS 0.250278f
C86 VN.n36 VSUBS 0.029116f
C87 VN.n37 VSUBS 0.053993f
C88 VN.n38 VSUBS 0.042325f
C89 VN.n39 VSUBS 0.042325f
C90 VN.n40 VSUBS 0.029116f
C91 VN.n41 VSUBS 0.029116f
C92 VN.n42 VSUBS 0.029116f
C93 VN.n43 VSUBS 0.030803f
C94 VN.n44 VSUBS 0.99004f
C95 VN.n45 VSUBS 0.050528f
C96 VN.n46 VSUBS 0.052019f
C97 VN.n47 VSUBS 0.029116f
C98 VN.n48 VSUBS 0.029116f
C99 VN.n49 VSUBS 0.029116f
C100 VN.n50 VSUBS 0.057284f
C101 VN.n51 VSUBS 0.037734f
C102 VN.n52 VSUBS 1.07458f
C103 VN.n53 VSUBS 1.72737f
C104 B.n0 VSUBS 0.004085f
C105 B.n1 VSUBS 0.004085f
C106 B.n2 VSUBS 0.00646f
C107 B.n3 VSUBS 0.00646f
C108 B.n4 VSUBS 0.00646f
C109 B.n5 VSUBS 0.00646f
C110 B.n6 VSUBS 0.00646f
C111 B.n7 VSUBS 0.00646f
C112 B.n8 VSUBS 0.00646f
C113 B.n9 VSUBS 0.00646f
C114 B.n10 VSUBS 0.00646f
C115 B.n11 VSUBS 0.00646f
C116 B.n12 VSUBS 0.00646f
C117 B.n13 VSUBS 0.00646f
C118 B.n14 VSUBS 0.00646f
C119 B.n15 VSUBS 0.00646f
C120 B.n16 VSUBS 0.00646f
C121 B.n17 VSUBS 0.00646f
C122 B.n18 VSUBS 0.00646f
C123 B.n19 VSUBS 0.00646f
C124 B.n20 VSUBS 0.00646f
C125 B.n21 VSUBS 0.00646f
C126 B.n22 VSUBS 0.00646f
C127 B.n23 VSUBS 0.00646f
C128 B.n24 VSUBS 0.00646f
C129 B.n25 VSUBS 0.013737f
C130 B.n26 VSUBS 0.00646f
C131 B.n27 VSUBS 0.00646f
C132 B.n28 VSUBS 0.00646f
C133 B.n29 VSUBS 0.00646f
C134 B.n30 VSUBS 0.00646f
C135 B.n31 VSUBS 0.00646f
C136 B.n32 VSUBS 0.00646f
C137 B.n33 VSUBS 0.00646f
C138 B.n34 VSUBS 0.00646f
C139 B.n35 VSUBS 0.00646f
C140 B.n36 VSUBS 0.00646f
C141 B.n37 VSUBS 0.00646f
C142 B.n38 VSUBS 0.00646f
C143 B.n39 VSUBS 0.00646f
C144 B.n40 VSUBS 0.00646f
C145 B.n41 VSUBS 0.00646f
C146 B.n42 VSUBS 0.00646f
C147 B.n43 VSUBS 0.00646f
C148 B.n44 VSUBS 0.00646f
C149 B.n45 VSUBS 0.00646f
C150 B.n46 VSUBS 0.00646f
C151 B.n47 VSUBS 0.00646f
C152 B.n48 VSUBS 0.00646f
C153 B.n49 VSUBS 0.00646f
C154 B.n50 VSUBS 0.00646f
C155 B.n51 VSUBS 0.00646f
C156 B.t8 VSUBS 0.266614f
C157 B.t7 VSUBS 0.294181f
C158 B.t6 VSUBS 1.45208f
C159 B.n52 VSUBS 0.450557f
C160 B.n53 VSUBS 0.272839f
C161 B.n54 VSUBS 0.00646f
C162 B.n55 VSUBS 0.00646f
C163 B.n56 VSUBS 0.00646f
C164 B.n57 VSUBS 0.00646f
C165 B.t5 VSUBS 0.266617f
C166 B.t4 VSUBS 0.294184f
C167 B.t3 VSUBS 1.45208f
C168 B.n58 VSUBS 0.450554f
C169 B.n59 VSUBS 0.272836f
C170 B.n60 VSUBS 0.014967f
C171 B.n61 VSUBS 0.00646f
C172 B.n62 VSUBS 0.00646f
C173 B.n63 VSUBS 0.00646f
C174 B.n64 VSUBS 0.00646f
C175 B.n65 VSUBS 0.00646f
C176 B.n66 VSUBS 0.00646f
C177 B.n67 VSUBS 0.00646f
C178 B.n68 VSUBS 0.00646f
C179 B.n69 VSUBS 0.00646f
C180 B.n70 VSUBS 0.00646f
C181 B.n71 VSUBS 0.00646f
C182 B.n72 VSUBS 0.00646f
C183 B.n73 VSUBS 0.00646f
C184 B.n74 VSUBS 0.00646f
C185 B.n75 VSUBS 0.00646f
C186 B.n76 VSUBS 0.00646f
C187 B.n77 VSUBS 0.00646f
C188 B.n78 VSUBS 0.00646f
C189 B.n79 VSUBS 0.00646f
C190 B.n80 VSUBS 0.00646f
C191 B.n81 VSUBS 0.00646f
C192 B.n82 VSUBS 0.00646f
C193 B.n83 VSUBS 0.00646f
C194 B.n84 VSUBS 0.00646f
C195 B.n85 VSUBS 0.00646f
C196 B.n86 VSUBS 0.013529f
C197 B.n87 VSUBS 0.00646f
C198 B.n88 VSUBS 0.00646f
C199 B.n89 VSUBS 0.00646f
C200 B.n90 VSUBS 0.00646f
C201 B.n91 VSUBS 0.00646f
C202 B.n92 VSUBS 0.00646f
C203 B.n93 VSUBS 0.00646f
C204 B.n94 VSUBS 0.00646f
C205 B.n95 VSUBS 0.00646f
C206 B.n96 VSUBS 0.00646f
C207 B.n97 VSUBS 0.00646f
C208 B.n98 VSUBS 0.00646f
C209 B.n99 VSUBS 0.00646f
C210 B.n100 VSUBS 0.00646f
C211 B.n101 VSUBS 0.00646f
C212 B.n102 VSUBS 0.00646f
C213 B.n103 VSUBS 0.00646f
C214 B.n104 VSUBS 0.00646f
C215 B.n105 VSUBS 0.00646f
C216 B.n106 VSUBS 0.00646f
C217 B.n107 VSUBS 0.00646f
C218 B.n108 VSUBS 0.00646f
C219 B.n109 VSUBS 0.00646f
C220 B.n110 VSUBS 0.00646f
C221 B.n111 VSUBS 0.00646f
C222 B.n112 VSUBS 0.00646f
C223 B.n113 VSUBS 0.00646f
C224 B.n114 VSUBS 0.00646f
C225 B.n115 VSUBS 0.00646f
C226 B.n116 VSUBS 0.00646f
C227 B.n117 VSUBS 0.00646f
C228 B.n118 VSUBS 0.00646f
C229 B.n119 VSUBS 0.00646f
C230 B.n120 VSUBS 0.00646f
C231 B.n121 VSUBS 0.00646f
C232 B.n122 VSUBS 0.00646f
C233 B.n123 VSUBS 0.00646f
C234 B.n124 VSUBS 0.00646f
C235 B.n125 VSUBS 0.00646f
C236 B.n126 VSUBS 0.00646f
C237 B.n127 VSUBS 0.00646f
C238 B.n128 VSUBS 0.00646f
C239 B.n129 VSUBS 0.00646f
C240 B.n130 VSUBS 0.00646f
C241 B.n131 VSUBS 0.00646f
C242 B.n132 VSUBS 0.00646f
C243 B.n133 VSUBS 0.00646f
C244 B.n134 VSUBS 0.014383f
C245 B.n135 VSUBS 0.00646f
C246 B.n136 VSUBS 0.00646f
C247 B.n137 VSUBS 0.00646f
C248 B.n138 VSUBS 0.00646f
C249 B.n139 VSUBS 0.00646f
C250 B.n140 VSUBS 0.00646f
C251 B.n141 VSUBS 0.00646f
C252 B.n142 VSUBS 0.00646f
C253 B.n143 VSUBS 0.00646f
C254 B.n144 VSUBS 0.00646f
C255 B.n145 VSUBS 0.00646f
C256 B.n146 VSUBS 0.00646f
C257 B.n147 VSUBS 0.00646f
C258 B.n148 VSUBS 0.00646f
C259 B.n149 VSUBS 0.00646f
C260 B.n150 VSUBS 0.00646f
C261 B.n151 VSUBS 0.00646f
C262 B.n152 VSUBS 0.00646f
C263 B.n153 VSUBS 0.00646f
C264 B.n154 VSUBS 0.00646f
C265 B.n155 VSUBS 0.00646f
C266 B.n156 VSUBS 0.00646f
C267 B.n157 VSUBS 0.00646f
C268 B.n158 VSUBS 0.00646f
C269 B.n159 VSUBS 0.00646f
C270 B.t1 VSUBS 0.266617f
C271 B.t2 VSUBS 0.294184f
C272 B.t0 VSUBS 1.45208f
C273 B.n160 VSUBS 0.450554f
C274 B.n161 VSUBS 0.272836f
C275 B.n162 VSUBS 0.014967f
C276 B.n163 VSUBS 0.00646f
C277 B.n164 VSUBS 0.00646f
C278 B.n165 VSUBS 0.00646f
C279 B.n166 VSUBS 0.00646f
C280 B.n167 VSUBS 0.00646f
C281 B.t10 VSUBS 0.266614f
C282 B.t11 VSUBS 0.294181f
C283 B.t9 VSUBS 1.45208f
C284 B.n168 VSUBS 0.450557f
C285 B.n169 VSUBS 0.272839f
C286 B.n170 VSUBS 0.00646f
C287 B.n171 VSUBS 0.00646f
C288 B.n172 VSUBS 0.00646f
C289 B.n173 VSUBS 0.00646f
C290 B.n174 VSUBS 0.00646f
C291 B.n175 VSUBS 0.00646f
C292 B.n176 VSUBS 0.00646f
C293 B.n177 VSUBS 0.00646f
C294 B.n178 VSUBS 0.00646f
C295 B.n179 VSUBS 0.00646f
C296 B.n180 VSUBS 0.00646f
C297 B.n181 VSUBS 0.00646f
C298 B.n182 VSUBS 0.00646f
C299 B.n183 VSUBS 0.00646f
C300 B.n184 VSUBS 0.00646f
C301 B.n185 VSUBS 0.00646f
C302 B.n186 VSUBS 0.00646f
C303 B.n187 VSUBS 0.00646f
C304 B.n188 VSUBS 0.00646f
C305 B.n189 VSUBS 0.00646f
C306 B.n190 VSUBS 0.00646f
C307 B.n191 VSUBS 0.00646f
C308 B.n192 VSUBS 0.00646f
C309 B.n193 VSUBS 0.00646f
C310 B.n194 VSUBS 0.00646f
C311 B.n195 VSUBS 0.013737f
C312 B.n196 VSUBS 0.00646f
C313 B.n197 VSUBS 0.00646f
C314 B.n198 VSUBS 0.00646f
C315 B.n199 VSUBS 0.00646f
C316 B.n200 VSUBS 0.00646f
C317 B.n201 VSUBS 0.00646f
C318 B.n202 VSUBS 0.00646f
C319 B.n203 VSUBS 0.00646f
C320 B.n204 VSUBS 0.00646f
C321 B.n205 VSUBS 0.00646f
C322 B.n206 VSUBS 0.00646f
C323 B.n207 VSUBS 0.00646f
C324 B.n208 VSUBS 0.00646f
C325 B.n209 VSUBS 0.00646f
C326 B.n210 VSUBS 0.00646f
C327 B.n211 VSUBS 0.00646f
C328 B.n212 VSUBS 0.00646f
C329 B.n213 VSUBS 0.00646f
C330 B.n214 VSUBS 0.00646f
C331 B.n215 VSUBS 0.00646f
C332 B.n216 VSUBS 0.00646f
C333 B.n217 VSUBS 0.00646f
C334 B.n218 VSUBS 0.00646f
C335 B.n219 VSUBS 0.00646f
C336 B.n220 VSUBS 0.00646f
C337 B.n221 VSUBS 0.00646f
C338 B.n222 VSUBS 0.00646f
C339 B.n223 VSUBS 0.00646f
C340 B.n224 VSUBS 0.00646f
C341 B.n225 VSUBS 0.00646f
C342 B.n226 VSUBS 0.00646f
C343 B.n227 VSUBS 0.00646f
C344 B.n228 VSUBS 0.00646f
C345 B.n229 VSUBS 0.00646f
C346 B.n230 VSUBS 0.00646f
C347 B.n231 VSUBS 0.00646f
C348 B.n232 VSUBS 0.00646f
C349 B.n233 VSUBS 0.00646f
C350 B.n234 VSUBS 0.00646f
C351 B.n235 VSUBS 0.00646f
C352 B.n236 VSUBS 0.00646f
C353 B.n237 VSUBS 0.00646f
C354 B.n238 VSUBS 0.00646f
C355 B.n239 VSUBS 0.00646f
C356 B.n240 VSUBS 0.00646f
C357 B.n241 VSUBS 0.00646f
C358 B.n242 VSUBS 0.00646f
C359 B.n243 VSUBS 0.00646f
C360 B.n244 VSUBS 0.00646f
C361 B.n245 VSUBS 0.00646f
C362 B.n246 VSUBS 0.00646f
C363 B.n247 VSUBS 0.00646f
C364 B.n248 VSUBS 0.00646f
C365 B.n249 VSUBS 0.00646f
C366 B.n250 VSUBS 0.00646f
C367 B.n251 VSUBS 0.00646f
C368 B.n252 VSUBS 0.00646f
C369 B.n253 VSUBS 0.00646f
C370 B.n254 VSUBS 0.00646f
C371 B.n255 VSUBS 0.00646f
C372 B.n256 VSUBS 0.00646f
C373 B.n257 VSUBS 0.00646f
C374 B.n258 VSUBS 0.00646f
C375 B.n259 VSUBS 0.00646f
C376 B.n260 VSUBS 0.00646f
C377 B.n261 VSUBS 0.00646f
C378 B.n262 VSUBS 0.00646f
C379 B.n263 VSUBS 0.00646f
C380 B.n264 VSUBS 0.00646f
C381 B.n265 VSUBS 0.00646f
C382 B.n266 VSUBS 0.00646f
C383 B.n267 VSUBS 0.00646f
C384 B.n268 VSUBS 0.00646f
C385 B.n269 VSUBS 0.00646f
C386 B.n270 VSUBS 0.00646f
C387 B.n271 VSUBS 0.00646f
C388 B.n272 VSUBS 0.00646f
C389 B.n273 VSUBS 0.00646f
C390 B.n274 VSUBS 0.00646f
C391 B.n275 VSUBS 0.00646f
C392 B.n276 VSUBS 0.00646f
C393 B.n277 VSUBS 0.00646f
C394 B.n278 VSUBS 0.00646f
C395 B.n279 VSUBS 0.00646f
C396 B.n280 VSUBS 0.00646f
C397 B.n281 VSUBS 0.00646f
C398 B.n282 VSUBS 0.00646f
C399 B.n283 VSUBS 0.00646f
C400 B.n284 VSUBS 0.00646f
C401 B.n285 VSUBS 0.00646f
C402 B.n286 VSUBS 0.013737f
C403 B.n287 VSUBS 0.014383f
C404 B.n288 VSUBS 0.014383f
C405 B.n289 VSUBS 0.00646f
C406 B.n290 VSUBS 0.00646f
C407 B.n291 VSUBS 0.00646f
C408 B.n292 VSUBS 0.00646f
C409 B.n293 VSUBS 0.00646f
C410 B.n294 VSUBS 0.00646f
C411 B.n295 VSUBS 0.00646f
C412 B.n296 VSUBS 0.00646f
C413 B.n297 VSUBS 0.00646f
C414 B.n298 VSUBS 0.00646f
C415 B.n299 VSUBS 0.00646f
C416 B.n300 VSUBS 0.00646f
C417 B.n301 VSUBS 0.00646f
C418 B.n302 VSUBS 0.00646f
C419 B.n303 VSUBS 0.00646f
C420 B.n304 VSUBS 0.00646f
C421 B.n305 VSUBS 0.00646f
C422 B.n306 VSUBS 0.00646f
C423 B.n307 VSUBS 0.00646f
C424 B.n308 VSUBS 0.00646f
C425 B.n309 VSUBS 0.00646f
C426 B.n310 VSUBS 0.00646f
C427 B.n311 VSUBS 0.00646f
C428 B.n312 VSUBS 0.00646f
C429 B.n313 VSUBS 0.00646f
C430 B.n314 VSUBS 0.00646f
C431 B.n315 VSUBS 0.00646f
C432 B.n316 VSUBS 0.00646f
C433 B.n317 VSUBS 0.00646f
C434 B.n318 VSUBS 0.00646f
C435 B.n319 VSUBS 0.00646f
C436 B.n320 VSUBS 0.00646f
C437 B.n321 VSUBS 0.00646f
C438 B.n322 VSUBS 0.00646f
C439 B.n323 VSUBS 0.00646f
C440 B.n324 VSUBS 0.00646f
C441 B.n325 VSUBS 0.00646f
C442 B.n326 VSUBS 0.00646f
C443 B.n327 VSUBS 0.00646f
C444 B.n328 VSUBS 0.00646f
C445 B.n329 VSUBS 0.00646f
C446 B.n330 VSUBS 0.00646f
C447 B.n331 VSUBS 0.00646f
C448 B.n332 VSUBS 0.00646f
C449 B.n333 VSUBS 0.00646f
C450 B.n334 VSUBS 0.00646f
C451 B.n335 VSUBS 0.00646f
C452 B.n336 VSUBS 0.00646f
C453 B.n337 VSUBS 0.00646f
C454 B.n338 VSUBS 0.00646f
C455 B.n339 VSUBS 0.00646f
C456 B.n340 VSUBS 0.00646f
C457 B.n341 VSUBS 0.00646f
C458 B.n342 VSUBS 0.00646f
C459 B.n343 VSUBS 0.00646f
C460 B.n344 VSUBS 0.00646f
C461 B.n345 VSUBS 0.00646f
C462 B.n346 VSUBS 0.00646f
C463 B.n347 VSUBS 0.00646f
C464 B.n348 VSUBS 0.00646f
C465 B.n349 VSUBS 0.00646f
C466 B.n350 VSUBS 0.00646f
C467 B.n351 VSUBS 0.00646f
C468 B.n352 VSUBS 0.00646f
C469 B.n353 VSUBS 0.00646f
C470 B.n354 VSUBS 0.00646f
C471 B.n355 VSUBS 0.00646f
C472 B.n356 VSUBS 0.00646f
C473 B.n357 VSUBS 0.00646f
C474 B.n358 VSUBS 0.00646f
C475 B.n359 VSUBS 0.00646f
C476 B.n360 VSUBS 0.00646f
C477 B.n361 VSUBS 0.00646f
C478 B.n362 VSUBS 0.00646f
C479 B.n363 VSUBS 0.00646f
C480 B.n364 VSUBS 0.004465f
C481 B.n365 VSUBS 0.014967f
C482 B.n366 VSUBS 0.005225f
C483 B.n367 VSUBS 0.00646f
C484 B.n368 VSUBS 0.00646f
C485 B.n369 VSUBS 0.00646f
C486 B.n370 VSUBS 0.00646f
C487 B.n371 VSUBS 0.00646f
C488 B.n372 VSUBS 0.00646f
C489 B.n373 VSUBS 0.00646f
C490 B.n374 VSUBS 0.00646f
C491 B.n375 VSUBS 0.00646f
C492 B.n376 VSUBS 0.00646f
C493 B.n377 VSUBS 0.00646f
C494 B.n378 VSUBS 0.005225f
C495 B.n379 VSUBS 0.00646f
C496 B.n380 VSUBS 0.00646f
C497 B.n381 VSUBS 0.004465f
C498 B.n382 VSUBS 0.00646f
C499 B.n383 VSUBS 0.00646f
C500 B.n384 VSUBS 0.00646f
C501 B.n385 VSUBS 0.00646f
C502 B.n386 VSUBS 0.00646f
C503 B.n387 VSUBS 0.00646f
C504 B.n388 VSUBS 0.00646f
C505 B.n389 VSUBS 0.00646f
C506 B.n390 VSUBS 0.00646f
C507 B.n391 VSUBS 0.00646f
C508 B.n392 VSUBS 0.00646f
C509 B.n393 VSUBS 0.00646f
C510 B.n394 VSUBS 0.00646f
C511 B.n395 VSUBS 0.00646f
C512 B.n396 VSUBS 0.00646f
C513 B.n397 VSUBS 0.00646f
C514 B.n398 VSUBS 0.00646f
C515 B.n399 VSUBS 0.00646f
C516 B.n400 VSUBS 0.00646f
C517 B.n401 VSUBS 0.00646f
C518 B.n402 VSUBS 0.00646f
C519 B.n403 VSUBS 0.00646f
C520 B.n404 VSUBS 0.00646f
C521 B.n405 VSUBS 0.00646f
C522 B.n406 VSUBS 0.00646f
C523 B.n407 VSUBS 0.00646f
C524 B.n408 VSUBS 0.00646f
C525 B.n409 VSUBS 0.00646f
C526 B.n410 VSUBS 0.00646f
C527 B.n411 VSUBS 0.00646f
C528 B.n412 VSUBS 0.00646f
C529 B.n413 VSUBS 0.00646f
C530 B.n414 VSUBS 0.00646f
C531 B.n415 VSUBS 0.00646f
C532 B.n416 VSUBS 0.00646f
C533 B.n417 VSUBS 0.00646f
C534 B.n418 VSUBS 0.00646f
C535 B.n419 VSUBS 0.00646f
C536 B.n420 VSUBS 0.00646f
C537 B.n421 VSUBS 0.00646f
C538 B.n422 VSUBS 0.00646f
C539 B.n423 VSUBS 0.00646f
C540 B.n424 VSUBS 0.00646f
C541 B.n425 VSUBS 0.00646f
C542 B.n426 VSUBS 0.00646f
C543 B.n427 VSUBS 0.00646f
C544 B.n428 VSUBS 0.00646f
C545 B.n429 VSUBS 0.00646f
C546 B.n430 VSUBS 0.00646f
C547 B.n431 VSUBS 0.00646f
C548 B.n432 VSUBS 0.00646f
C549 B.n433 VSUBS 0.00646f
C550 B.n434 VSUBS 0.00646f
C551 B.n435 VSUBS 0.00646f
C552 B.n436 VSUBS 0.00646f
C553 B.n437 VSUBS 0.00646f
C554 B.n438 VSUBS 0.00646f
C555 B.n439 VSUBS 0.00646f
C556 B.n440 VSUBS 0.00646f
C557 B.n441 VSUBS 0.00646f
C558 B.n442 VSUBS 0.00646f
C559 B.n443 VSUBS 0.00646f
C560 B.n444 VSUBS 0.00646f
C561 B.n445 VSUBS 0.00646f
C562 B.n446 VSUBS 0.00646f
C563 B.n447 VSUBS 0.00646f
C564 B.n448 VSUBS 0.00646f
C565 B.n449 VSUBS 0.00646f
C566 B.n450 VSUBS 0.00646f
C567 B.n451 VSUBS 0.00646f
C568 B.n452 VSUBS 0.00646f
C569 B.n453 VSUBS 0.00646f
C570 B.n454 VSUBS 0.00646f
C571 B.n455 VSUBS 0.00646f
C572 B.n456 VSUBS 0.00646f
C573 B.n457 VSUBS 0.014383f
C574 B.n458 VSUBS 0.013737f
C575 B.n459 VSUBS 0.013737f
C576 B.n460 VSUBS 0.00646f
C577 B.n461 VSUBS 0.00646f
C578 B.n462 VSUBS 0.00646f
C579 B.n463 VSUBS 0.00646f
C580 B.n464 VSUBS 0.00646f
C581 B.n465 VSUBS 0.00646f
C582 B.n466 VSUBS 0.00646f
C583 B.n467 VSUBS 0.00646f
C584 B.n468 VSUBS 0.00646f
C585 B.n469 VSUBS 0.00646f
C586 B.n470 VSUBS 0.00646f
C587 B.n471 VSUBS 0.00646f
C588 B.n472 VSUBS 0.00646f
C589 B.n473 VSUBS 0.00646f
C590 B.n474 VSUBS 0.00646f
C591 B.n475 VSUBS 0.00646f
C592 B.n476 VSUBS 0.00646f
C593 B.n477 VSUBS 0.00646f
C594 B.n478 VSUBS 0.00646f
C595 B.n479 VSUBS 0.00646f
C596 B.n480 VSUBS 0.00646f
C597 B.n481 VSUBS 0.00646f
C598 B.n482 VSUBS 0.00646f
C599 B.n483 VSUBS 0.00646f
C600 B.n484 VSUBS 0.00646f
C601 B.n485 VSUBS 0.00646f
C602 B.n486 VSUBS 0.00646f
C603 B.n487 VSUBS 0.00646f
C604 B.n488 VSUBS 0.00646f
C605 B.n489 VSUBS 0.00646f
C606 B.n490 VSUBS 0.00646f
C607 B.n491 VSUBS 0.00646f
C608 B.n492 VSUBS 0.00646f
C609 B.n493 VSUBS 0.00646f
C610 B.n494 VSUBS 0.00646f
C611 B.n495 VSUBS 0.00646f
C612 B.n496 VSUBS 0.00646f
C613 B.n497 VSUBS 0.00646f
C614 B.n498 VSUBS 0.00646f
C615 B.n499 VSUBS 0.00646f
C616 B.n500 VSUBS 0.00646f
C617 B.n501 VSUBS 0.00646f
C618 B.n502 VSUBS 0.00646f
C619 B.n503 VSUBS 0.00646f
C620 B.n504 VSUBS 0.00646f
C621 B.n505 VSUBS 0.00646f
C622 B.n506 VSUBS 0.00646f
C623 B.n507 VSUBS 0.00646f
C624 B.n508 VSUBS 0.00646f
C625 B.n509 VSUBS 0.00646f
C626 B.n510 VSUBS 0.00646f
C627 B.n511 VSUBS 0.00646f
C628 B.n512 VSUBS 0.00646f
C629 B.n513 VSUBS 0.00646f
C630 B.n514 VSUBS 0.00646f
C631 B.n515 VSUBS 0.00646f
C632 B.n516 VSUBS 0.00646f
C633 B.n517 VSUBS 0.00646f
C634 B.n518 VSUBS 0.00646f
C635 B.n519 VSUBS 0.00646f
C636 B.n520 VSUBS 0.00646f
C637 B.n521 VSUBS 0.00646f
C638 B.n522 VSUBS 0.00646f
C639 B.n523 VSUBS 0.00646f
C640 B.n524 VSUBS 0.00646f
C641 B.n525 VSUBS 0.00646f
C642 B.n526 VSUBS 0.00646f
C643 B.n527 VSUBS 0.00646f
C644 B.n528 VSUBS 0.00646f
C645 B.n529 VSUBS 0.00646f
C646 B.n530 VSUBS 0.00646f
C647 B.n531 VSUBS 0.00646f
C648 B.n532 VSUBS 0.00646f
C649 B.n533 VSUBS 0.00646f
C650 B.n534 VSUBS 0.00646f
C651 B.n535 VSUBS 0.00646f
C652 B.n536 VSUBS 0.00646f
C653 B.n537 VSUBS 0.00646f
C654 B.n538 VSUBS 0.00646f
C655 B.n539 VSUBS 0.00646f
C656 B.n540 VSUBS 0.00646f
C657 B.n541 VSUBS 0.00646f
C658 B.n542 VSUBS 0.00646f
C659 B.n543 VSUBS 0.00646f
C660 B.n544 VSUBS 0.00646f
C661 B.n545 VSUBS 0.00646f
C662 B.n546 VSUBS 0.00646f
C663 B.n547 VSUBS 0.00646f
C664 B.n548 VSUBS 0.00646f
C665 B.n549 VSUBS 0.00646f
C666 B.n550 VSUBS 0.00646f
C667 B.n551 VSUBS 0.00646f
C668 B.n552 VSUBS 0.00646f
C669 B.n553 VSUBS 0.00646f
C670 B.n554 VSUBS 0.00646f
C671 B.n555 VSUBS 0.00646f
C672 B.n556 VSUBS 0.00646f
C673 B.n557 VSUBS 0.00646f
C674 B.n558 VSUBS 0.00646f
C675 B.n559 VSUBS 0.00646f
C676 B.n560 VSUBS 0.00646f
C677 B.n561 VSUBS 0.00646f
C678 B.n562 VSUBS 0.00646f
C679 B.n563 VSUBS 0.00646f
C680 B.n564 VSUBS 0.00646f
C681 B.n565 VSUBS 0.00646f
C682 B.n566 VSUBS 0.00646f
C683 B.n567 VSUBS 0.00646f
C684 B.n568 VSUBS 0.00646f
C685 B.n569 VSUBS 0.00646f
C686 B.n570 VSUBS 0.00646f
C687 B.n571 VSUBS 0.00646f
C688 B.n572 VSUBS 0.00646f
C689 B.n573 VSUBS 0.00646f
C690 B.n574 VSUBS 0.00646f
C691 B.n575 VSUBS 0.00646f
C692 B.n576 VSUBS 0.00646f
C693 B.n577 VSUBS 0.00646f
C694 B.n578 VSUBS 0.00646f
C695 B.n579 VSUBS 0.00646f
C696 B.n580 VSUBS 0.00646f
C697 B.n581 VSUBS 0.00646f
C698 B.n582 VSUBS 0.00646f
C699 B.n583 VSUBS 0.00646f
C700 B.n584 VSUBS 0.00646f
C701 B.n585 VSUBS 0.00646f
C702 B.n586 VSUBS 0.00646f
C703 B.n587 VSUBS 0.00646f
C704 B.n588 VSUBS 0.00646f
C705 B.n589 VSUBS 0.00646f
C706 B.n590 VSUBS 0.00646f
C707 B.n591 VSUBS 0.00646f
C708 B.n592 VSUBS 0.00646f
C709 B.n593 VSUBS 0.00646f
C710 B.n594 VSUBS 0.00646f
C711 B.n595 VSUBS 0.00646f
C712 B.n596 VSUBS 0.00646f
C713 B.n597 VSUBS 0.00646f
C714 B.n598 VSUBS 0.00646f
C715 B.n599 VSUBS 0.014591f
C716 B.n600 VSUBS 0.013737f
C717 B.n601 VSUBS 0.014383f
C718 B.n602 VSUBS 0.00646f
C719 B.n603 VSUBS 0.00646f
C720 B.n604 VSUBS 0.00646f
C721 B.n605 VSUBS 0.00646f
C722 B.n606 VSUBS 0.00646f
C723 B.n607 VSUBS 0.00646f
C724 B.n608 VSUBS 0.00646f
C725 B.n609 VSUBS 0.00646f
C726 B.n610 VSUBS 0.00646f
C727 B.n611 VSUBS 0.00646f
C728 B.n612 VSUBS 0.00646f
C729 B.n613 VSUBS 0.00646f
C730 B.n614 VSUBS 0.00646f
C731 B.n615 VSUBS 0.00646f
C732 B.n616 VSUBS 0.00646f
C733 B.n617 VSUBS 0.00646f
C734 B.n618 VSUBS 0.00646f
C735 B.n619 VSUBS 0.00646f
C736 B.n620 VSUBS 0.00646f
C737 B.n621 VSUBS 0.00646f
C738 B.n622 VSUBS 0.00646f
C739 B.n623 VSUBS 0.00646f
C740 B.n624 VSUBS 0.00646f
C741 B.n625 VSUBS 0.00646f
C742 B.n626 VSUBS 0.00646f
C743 B.n627 VSUBS 0.00646f
C744 B.n628 VSUBS 0.00646f
C745 B.n629 VSUBS 0.00646f
C746 B.n630 VSUBS 0.00646f
C747 B.n631 VSUBS 0.00646f
C748 B.n632 VSUBS 0.00646f
C749 B.n633 VSUBS 0.00646f
C750 B.n634 VSUBS 0.00646f
C751 B.n635 VSUBS 0.00646f
C752 B.n636 VSUBS 0.00646f
C753 B.n637 VSUBS 0.00646f
C754 B.n638 VSUBS 0.00646f
C755 B.n639 VSUBS 0.00646f
C756 B.n640 VSUBS 0.00646f
C757 B.n641 VSUBS 0.00646f
C758 B.n642 VSUBS 0.00646f
C759 B.n643 VSUBS 0.00646f
C760 B.n644 VSUBS 0.00646f
C761 B.n645 VSUBS 0.00646f
C762 B.n646 VSUBS 0.00646f
C763 B.n647 VSUBS 0.00646f
C764 B.n648 VSUBS 0.00646f
C765 B.n649 VSUBS 0.00646f
C766 B.n650 VSUBS 0.00646f
C767 B.n651 VSUBS 0.00646f
C768 B.n652 VSUBS 0.00646f
C769 B.n653 VSUBS 0.00646f
C770 B.n654 VSUBS 0.00646f
C771 B.n655 VSUBS 0.00646f
C772 B.n656 VSUBS 0.00646f
C773 B.n657 VSUBS 0.00646f
C774 B.n658 VSUBS 0.00646f
C775 B.n659 VSUBS 0.00646f
C776 B.n660 VSUBS 0.00646f
C777 B.n661 VSUBS 0.00646f
C778 B.n662 VSUBS 0.00646f
C779 B.n663 VSUBS 0.00646f
C780 B.n664 VSUBS 0.00646f
C781 B.n665 VSUBS 0.00646f
C782 B.n666 VSUBS 0.00646f
C783 B.n667 VSUBS 0.00646f
C784 B.n668 VSUBS 0.00646f
C785 B.n669 VSUBS 0.00646f
C786 B.n670 VSUBS 0.00646f
C787 B.n671 VSUBS 0.00646f
C788 B.n672 VSUBS 0.00646f
C789 B.n673 VSUBS 0.00646f
C790 B.n674 VSUBS 0.00646f
C791 B.n675 VSUBS 0.00646f
C792 B.n676 VSUBS 0.00646f
C793 B.n677 VSUBS 0.004465f
C794 B.n678 VSUBS 0.00646f
C795 B.n679 VSUBS 0.00646f
C796 B.n680 VSUBS 0.005225f
C797 B.n681 VSUBS 0.00646f
C798 B.n682 VSUBS 0.00646f
C799 B.n683 VSUBS 0.00646f
C800 B.n684 VSUBS 0.00646f
C801 B.n685 VSUBS 0.00646f
C802 B.n686 VSUBS 0.00646f
C803 B.n687 VSUBS 0.00646f
C804 B.n688 VSUBS 0.00646f
C805 B.n689 VSUBS 0.00646f
C806 B.n690 VSUBS 0.00646f
C807 B.n691 VSUBS 0.00646f
C808 B.n692 VSUBS 0.005225f
C809 B.n693 VSUBS 0.014967f
C810 B.n694 VSUBS 0.004465f
C811 B.n695 VSUBS 0.00646f
C812 B.n696 VSUBS 0.00646f
C813 B.n697 VSUBS 0.00646f
C814 B.n698 VSUBS 0.00646f
C815 B.n699 VSUBS 0.00646f
C816 B.n700 VSUBS 0.00646f
C817 B.n701 VSUBS 0.00646f
C818 B.n702 VSUBS 0.00646f
C819 B.n703 VSUBS 0.00646f
C820 B.n704 VSUBS 0.00646f
C821 B.n705 VSUBS 0.00646f
C822 B.n706 VSUBS 0.00646f
C823 B.n707 VSUBS 0.00646f
C824 B.n708 VSUBS 0.00646f
C825 B.n709 VSUBS 0.00646f
C826 B.n710 VSUBS 0.00646f
C827 B.n711 VSUBS 0.00646f
C828 B.n712 VSUBS 0.00646f
C829 B.n713 VSUBS 0.00646f
C830 B.n714 VSUBS 0.00646f
C831 B.n715 VSUBS 0.00646f
C832 B.n716 VSUBS 0.00646f
C833 B.n717 VSUBS 0.00646f
C834 B.n718 VSUBS 0.00646f
C835 B.n719 VSUBS 0.00646f
C836 B.n720 VSUBS 0.00646f
C837 B.n721 VSUBS 0.00646f
C838 B.n722 VSUBS 0.00646f
C839 B.n723 VSUBS 0.00646f
C840 B.n724 VSUBS 0.00646f
C841 B.n725 VSUBS 0.00646f
C842 B.n726 VSUBS 0.00646f
C843 B.n727 VSUBS 0.00646f
C844 B.n728 VSUBS 0.00646f
C845 B.n729 VSUBS 0.00646f
C846 B.n730 VSUBS 0.00646f
C847 B.n731 VSUBS 0.00646f
C848 B.n732 VSUBS 0.00646f
C849 B.n733 VSUBS 0.00646f
C850 B.n734 VSUBS 0.00646f
C851 B.n735 VSUBS 0.00646f
C852 B.n736 VSUBS 0.00646f
C853 B.n737 VSUBS 0.00646f
C854 B.n738 VSUBS 0.00646f
C855 B.n739 VSUBS 0.00646f
C856 B.n740 VSUBS 0.00646f
C857 B.n741 VSUBS 0.00646f
C858 B.n742 VSUBS 0.00646f
C859 B.n743 VSUBS 0.00646f
C860 B.n744 VSUBS 0.00646f
C861 B.n745 VSUBS 0.00646f
C862 B.n746 VSUBS 0.00646f
C863 B.n747 VSUBS 0.00646f
C864 B.n748 VSUBS 0.00646f
C865 B.n749 VSUBS 0.00646f
C866 B.n750 VSUBS 0.00646f
C867 B.n751 VSUBS 0.00646f
C868 B.n752 VSUBS 0.00646f
C869 B.n753 VSUBS 0.00646f
C870 B.n754 VSUBS 0.00646f
C871 B.n755 VSUBS 0.00646f
C872 B.n756 VSUBS 0.00646f
C873 B.n757 VSUBS 0.00646f
C874 B.n758 VSUBS 0.00646f
C875 B.n759 VSUBS 0.00646f
C876 B.n760 VSUBS 0.00646f
C877 B.n761 VSUBS 0.00646f
C878 B.n762 VSUBS 0.00646f
C879 B.n763 VSUBS 0.00646f
C880 B.n764 VSUBS 0.00646f
C881 B.n765 VSUBS 0.00646f
C882 B.n766 VSUBS 0.00646f
C883 B.n767 VSUBS 0.00646f
C884 B.n768 VSUBS 0.00646f
C885 B.n769 VSUBS 0.00646f
C886 B.n770 VSUBS 0.014383f
C887 B.n771 VSUBS 0.014383f
C888 B.n772 VSUBS 0.013737f
C889 B.n773 VSUBS 0.00646f
C890 B.n774 VSUBS 0.00646f
C891 B.n775 VSUBS 0.00646f
C892 B.n776 VSUBS 0.00646f
C893 B.n777 VSUBS 0.00646f
C894 B.n778 VSUBS 0.00646f
C895 B.n779 VSUBS 0.00646f
C896 B.n780 VSUBS 0.00646f
C897 B.n781 VSUBS 0.00646f
C898 B.n782 VSUBS 0.00646f
C899 B.n783 VSUBS 0.00646f
C900 B.n784 VSUBS 0.00646f
C901 B.n785 VSUBS 0.00646f
C902 B.n786 VSUBS 0.00646f
C903 B.n787 VSUBS 0.00646f
C904 B.n788 VSUBS 0.00646f
C905 B.n789 VSUBS 0.00646f
C906 B.n790 VSUBS 0.00646f
C907 B.n791 VSUBS 0.00646f
C908 B.n792 VSUBS 0.00646f
C909 B.n793 VSUBS 0.00646f
C910 B.n794 VSUBS 0.00646f
C911 B.n795 VSUBS 0.00646f
C912 B.n796 VSUBS 0.00646f
C913 B.n797 VSUBS 0.00646f
C914 B.n798 VSUBS 0.00646f
C915 B.n799 VSUBS 0.00646f
C916 B.n800 VSUBS 0.00646f
C917 B.n801 VSUBS 0.00646f
C918 B.n802 VSUBS 0.00646f
C919 B.n803 VSUBS 0.00646f
C920 B.n804 VSUBS 0.00646f
C921 B.n805 VSUBS 0.00646f
C922 B.n806 VSUBS 0.00646f
C923 B.n807 VSUBS 0.00646f
C924 B.n808 VSUBS 0.00646f
C925 B.n809 VSUBS 0.00646f
C926 B.n810 VSUBS 0.00646f
C927 B.n811 VSUBS 0.00646f
C928 B.n812 VSUBS 0.00646f
C929 B.n813 VSUBS 0.00646f
C930 B.n814 VSUBS 0.00646f
C931 B.n815 VSUBS 0.00646f
C932 B.n816 VSUBS 0.00646f
C933 B.n817 VSUBS 0.00646f
C934 B.n818 VSUBS 0.00646f
C935 B.n819 VSUBS 0.00646f
C936 B.n820 VSUBS 0.00646f
C937 B.n821 VSUBS 0.00646f
C938 B.n822 VSUBS 0.00646f
C939 B.n823 VSUBS 0.00646f
C940 B.n824 VSUBS 0.00646f
C941 B.n825 VSUBS 0.00646f
C942 B.n826 VSUBS 0.00646f
C943 B.n827 VSUBS 0.00646f
C944 B.n828 VSUBS 0.00646f
C945 B.n829 VSUBS 0.00646f
C946 B.n830 VSUBS 0.00646f
C947 B.n831 VSUBS 0.00646f
C948 B.n832 VSUBS 0.00646f
C949 B.n833 VSUBS 0.00646f
C950 B.n834 VSUBS 0.00646f
C951 B.n835 VSUBS 0.00646f
C952 B.n836 VSUBS 0.00646f
C953 B.n837 VSUBS 0.00646f
C954 B.n838 VSUBS 0.00646f
C955 B.n839 VSUBS 0.00646f
C956 B.n840 VSUBS 0.00646f
C957 B.n841 VSUBS 0.00646f
C958 B.n842 VSUBS 0.00646f
C959 B.n843 VSUBS 0.014628f
C960 VDD1.t0 VSUBS 0.300653f
C961 VDD1.t2 VSUBS 0.300653f
C962 VDD1.n0 VSUBS 2.46329f
C963 VDD1.t4 VSUBS 0.300653f
C964 VDD1.t6 VSUBS 0.300653f
C965 VDD1.n1 VSUBS 2.46198f
C966 VDD1.t5 VSUBS 0.300653f
C967 VDD1.t7 VSUBS 0.300653f
C968 VDD1.n2 VSUBS 2.46198f
C969 VDD1.n3 VSUBS 3.8626f
C970 VDD1.t1 VSUBS 0.300653f
C971 VDD1.t3 VSUBS 0.300653f
C972 VDD1.n4 VSUBS 2.45077f
C973 VDD1.n5 VSUBS 3.36804f
C974 VTAIL.t2 VSUBS 0.291149f
C975 VTAIL.t1 VSUBS 0.291149f
C976 VTAIL.n0 VSUBS 2.23419f
C977 VTAIL.n1 VSUBS 0.743771f
C978 VTAIL.n2 VSUBS 0.024971f
C979 VTAIL.n3 VSUBS 0.023924f
C980 VTAIL.n4 VSUBS 0.012856f
C981 VTAIL.n5 VSUBS 0.030387f
C982 VTAIL.n6 VSUBS 0.013234f
C983 VTAIL.n7 VSUBS 0.023924f
C984 VTAIL.n8 VSUBS 0.013612f
C985 VTAIL.n9 VSUBS 0.030387f
C986 VTAIL.n10 VSUBS 0.013612f
C987 VTAIL.n11 VSUBS 0.023924f
C988 VTAIL.n12 VSUBS 0.012856f
C989 VTAIL.n13 VSUBS 0.030387f
C990 VTAIL.n14 VSUBS 0.013612f
C991 VTAIL.n15 VSUBS 0.023924f
C992 VTAIL.n16 VSUBS 0.012856f
C993 VTAIL.n17 VSUBS 0.030387f
C994 VTAIL.n18 VSUBS 0.013612f
C995 VTAIL.n19 VSUBS 0.023924f
C996 VTAIL.n20 VSUBS 0.012856f
C997 VTAIL.n21 VSUBS 0.030387f
C998 VTAIL.n22 VSUBS 0.013612f
C999 VTAIL.n23 VSUBS 0.023924f
C1000 VTAIL.n24 VSUBS 0.012856f
C1001 VTAIL.n25 VSUBS 0.030387f
C1002 VTAIL.n26 VSUBS 0.013612f
C1003 VTAIL.n27 VSUBS 1.57107f
C1004 VTAIL.n28 VSUBS 0.012856f
C1005 VTAIL.t3 VSUBS 0.065076f
C1006 VTAIL.n29 VSUBS 0.171469f
C1007 VTAIL.n30 VSUBS 0.019331f
C1008 VTAIL.n31 VSUBS 0.02279f
C1009 VTAIL.n32 VSUBS 0.030387f
C1010 VTAIL.n33 VSUBS 0.013612f
C1011 VTAIL.n34 VSUBS 0.012856f
C1012 VTAIL.n35 VSUBS 0.023924f
C1013 VTAIL.n36 VSUBS 0.023924f
C1014 VTAIL.n37 VSUBS 0.012856f
C1015 VTAIL.n38 VSUBS 0.013612f
C1016 VTAIL.n39 VSUBS 0.030387f
C1017 VTAIL.n40 VSUBS 0.030387f
C1018 VTAIL.n41 VSUBS 0.013612f
C1019 VTAIL.n42 VSUBS 0.012856f
C1020 VTAIL.n43 VSUBS 0.023924f
C1021 VTAIL.n44 VSUBS 0.023924f
C1022 VTAIL.n45 VSUBS 0.012856f
C1023 VTAIL.n46 VSUBS 0.013612f
C1024 VTAIL.n47 VSUBS 0.030387f
C1025 VTAIL.n48 VSUBS 0.030387f
C1026 VTAIL.n49 VSUBS 0.013612f
C1027 VTAIL.n50 VSUBS 0.012856f
C1028 VTAIL.n51 VSUBS 0.023924f
C1029 VTAIL.n52 VSUBS 0.023924f
C1030 VTAIL.n53 VSUBS 0.012856f
C1031 VTAIL.n54 VSUBS 0.013612f
C1032 VTAIL.n55 VSUBS 0.030387f
C1033 VTAIL.n56 VSUBS 0.030387f
C1034 VTAIL.n57 VSUBS 0.013612f
C1035 VTAIL.n58 VSUBS 0.012856f
C1036 VTAIL.n59 VSUBS 0.023924f
C1037 VTAIL.n60 VSUBS 0.023924f
C1038 VTAIL.n61 VSUBS 0.012856f
C1039 VTAIL.n62 VSUBS 0.013612f
C1040 VTAIL.n63 VSUBS 0.030387f
C1041 VTAIL.n64 VSUBS 0.030387f
C1042 VTAIL.n65 VSUBS 0.013612f
C1043 VTAIL.n66 VSUBS 0.012856f
C1044 VTAIL.n67 VSUBS 0.023924f
C1045 VTAIL.n68 VSUBS 0.023924f
C1046 VTAIL.n69 VSUBS 0.012856f
C1047 VTAIL.n70 VSUBS 0.012856f
C1048 VTAIL.n71 VSUBS 0.013612f
C1049 VTAIL.n72 VSUBS 0.030387f
C1050 VTAIL.n73 VSUBS 0.030387f
C1051 VTAIL.n74 VSUBS 0.030387f
C1052 VTAIL.n75 VSUBS 0.013234f
C1053 VTAIL.n76 VSUBS 0.012856f
C1054 VTAIL.n77 VSUBS 0.023924f
C1055 VTAIL.n78 VSUBS 0.023924f
C1056 VTAIL.n79 VSUBS 0.012856f
C1057 VTAIL.n80 VSUBS 0.013612f
C1058 VTAIL.n81 VSUBS 0.030387f
C1059 VTAIL.n82 VSUBS 0.069077f
C1060 VTAIL.n83 VSUBS 0.013612f
C1061 VTAIL.n84 VSUBS 0.012856f
C1062 VTAIL.n85 VSUBS 0.056607f
C1063 VTAIL.n86 VSUBS 0.034579f
C1064 VTAIL.n87 VSUBS 0.232172f
C1065 VTAIL.n88 VSUBS 0.024971f
C1066 VTAIL.n89 VSUBS 0.023924f
C1067 VTAIL.n90 VSUBS 0.012856f
C1068 VTAIL.n91 VSUBS 0.030387f
C1069 VTAIL.n92 VSUBS 0.013234f
C1070 VTAIL.n93 VSUBS 0.023924f
C1071 VTAIL.n94 VSUBS 0.013612f
C1072 VTAIL.n95 VSUBS 0.030387f
C1073 VTAIL.n96 VSUBS 0.013612f
C1074 VTAIL.n97 VSUBS 0.023924f
C1075 VTAIL.n98 VSUBS 0.012856f
C1076 VTAIL.n99 VSUBS 0.030387f
C1077 VTAIL.n100 VSUBS 0.013612f
C1078 VTAIL.n101 VSUBS 0.023924f
C1079 VTAIL.n102 VSUBS 0.012856f
C1080 VTAIL.n103 VSUBS 0.030387f
C1081 VTAIL.n104 VSUBS 0.013612f
C1082 VTAIL.n105 VSUBS 0.023924f
C1083 VTAIL.n106 VSUBS 0.012856f
C1084 VTAIL.n107 VSUBS 0.030387f
C1085 VTAIL.n108 VSUBS 0.013612f
C1086 VTAIL.n109 VSUBS 0.023924f
C1087 VTAIL.n110 VSUBS 0.012856f
C1088 VTAIL.n111 VSUBS 0.030387f
C1089 VTAIL.n112 VSUBS 0.013612f
C1090 VTAIL.n113 VSUBS 1.57107f
C1091 VTAIL.n114 VSUBS 0.012856f
C1092 VTAIL.t10 VSUBS 0.065076f
C1093 VTAIL.n115 VSUBS 0.171469f
C1094 VTAIL.n116 VSUBS 0.019331f
C1095 VTAIL.n117 VSUBS 0.02279f
C1096 VTAIL.n118 VSUBS 0.030387f
C1097 VTAIL.n119 VSUBS 0.013612f
C1098 VTAIL.n120 VSUBS 0.012856f
C1099 VTAIL.n121 VSUBS 0.023924f
C1100 VTAIL.n122 VSUBS 0.023924f
C1101 VTAIL.n123 VSUBS 0.012856f
C1102 VTAIL.n124 VSUBS 0.013612f
C1103 VTAIL.n125 VSUBS 0.030387f
C1104 VTAIL.n126 VSUBS 0.030387f
C1105 VTAIL.n127 VSUBS 0.013612f
C1106 VTAIL.n128 VSUBS 0.012856f
C1107 VTAIL.n129 VSUBS 0.023924f
C1108 VTAIL.n130 VSUBS 0.023924f
C1109 VTAIL.n131 VSUBS 0.012856f
C1110 VTAIL.n132 VSUBS 0.013612f
C1111 VTAIL.n133 VSUBS 0.030387f
C1112 VTAIL.n134 VSUBS 0.030387f
C1113 VTAIL.n135 VSUBS 0.013612f
C1114 VTAIL.n136 VSUBS 0.012856f
C1115 VTAIL.n137 VSUBS 0.023924f
C1116 VTAIL.n138 VSUBS 0.023924f
C1117 VTAIL.n139 VSUBS 0.012856f
C1118 VTAIL.n140 VSUBS 0.013612f
C1119 VTAIL.n141 VSUBS 0.030387f
C1120 VTAIL.n142 VSUBS 0.030387f
C1121 VTAIL.n143 VSUBS 0.013612f
C1122 VTAIL.n144 VSUBS 0.012856f
C1123 VTAIL.n145 VSUBS 0.023924f
C1124 VTAIL.n146 VSUBS 0.023924f
C1125 VTAIL.n147 VSUBS 0.012856f
C1126 VTAIL.n148 VSUBS 0.013612f
C1127 VTAIL.n149 VSUBS 0.030387f
C1128 VTAIL.n150 VSUBS 0.030387f
C1129 VTAIL.n151 VSUBS 0.013612f
C1130 VTAIL.n152 VSUBS 0.012856f
C1131 VTAIL.n153 VSUBS 0.023924f
C1132 VTAIL.n154 VSUBS 0.023924f
C1133 VTAIL.n155 VSUBS 0.012856f
C1134 VTAIL.n156 VSUBS 0.012856f
C1135 VTAIL.n157 VSUBS 0.013612f
C1136 VTAIL.n158 VSUBS 0.030387f
C1137 VTAIL.n159 VSUBS 0.030387f
C1138 VTAIL.n160 VSUBS 0.030387f
C1139 VTAIL.n161 VSUBS 0.013234f
C1140 VTAIL.n162 VSUBS 0.012856f
C1141 VTAIL.n163 VSUBS 0.023924f
C1142 VTAIL.n164 VSUBS 0.023924f
C1143 VTAIL.n165 VSUBS 0.012856f
C1144 VTAIL.n166 VSUBS 0.013612f
C1145 VTAIL.n167 VSUBS 0.030387f
C1146 VTAIL.n168 VSUBS 0.069077f
C1147 VTAIL.n169 VSUBS 0.013612f
C1148 VTAIL.n170 VSUBS 0.012856f
C1149 VTAIL.n171 VSUBS 0.056607f
C1150 VTAIL.n172 VSUBS 0.034579f
C1151 VTAIL.n173 VSUBS 0.232172f
C1152 VTAIL.t12 VSUBS 0.291149f
C1153 VTAIL.t15 VSUBS 0.291149f
C1154 VTAIL.n174 VSUBS 2.23419f
C1155 VTAIL.n175 VSUBS 0.914066f
C1156 VTAIL.n176 VSUBS 0.024971f
C1157 VTAIL.n177 VSUBS 0.023924f
C1158 VTAIL.n178 VSUBS 0.012856f
C1159 VTAIL.n179 VSUBS 0.030387f
C1160 VTAIL.n180 VSUBS 0.013234f
C1161 VTAIL.n181 VSUBS 0.023924f
C1162 VTAIL.n182 VSUBS 0.013612f
C1163 VTAIL.n183 VSUBS 0.030387f
C1164 VTAIL.n184 VSUBS 0.013612f
C1165 VTAIL.n185 VSUBS 0.023924f
C1166 VTAIL.n186 VSUBS 0.012856f
C1167 VTAIL.n187 VSUBS 0.030387f
C1168 VTAIL.n188 VSUBS 0.013612f
C1169 VTAIL.n189 VSUBS 0.023924f
C1170 VTAIL.n190 VSUBS 0.012856f
C1171 VTAIL.n191 VSUBS 0.030387f
C1172 VTAIL.n192 VSUBS 0.013612f
C1173 VTAIL.n193 VSUBS 0.023924f
C1174 VTAIL.n194 VSUBS 0.012856f
C1175 VTAIL.n195 VSUBS 0.030387f
C1176 VTAIL.n196 VSUBS 0.013612f
C1177 VTAIL.n197 VSUBS 0.023924f
C1178 VTAIL.n198 VSUBS 0.012856f
C1179 VTAIL.n199 VSUBS 0.030387f
C1180 VTAIL.n200 VSUBS 0.013612f
C1181 VTAIL.n201 VSUBS 1.57107f
C1182 VTAIL.n202 VSUBS 0.012856f
C1183 VTAIL.t9 VSUBS 0.065076f
C1184 VTAIL.n203 VSUBS 0.171469f
C1185 VTAIL.n204 VSUBS 0.019331f
C1186 VTAIL.n205 VSUBS 0.02279f
C1187 VTAIL.n206 VSUBS 0.030387f
C1188 VTAIL.n207 VSUBS 0.013612f
C1189 VTAIL.n208 VSUBS 0.012856f
C1190 VTAIL.n209 VSUBS 0.023924f
C1191 VTAIL.n210 VSUBS 0.023924f
C1192 VTAIL.n211 VSUBS 0.012856f
C1193 VTAIL.n212 VSUBS 0.013612f
C1194 VTAIL.n213 VSUBS 0.030387f
C1195 VTAIL.n214 VSUBS 0.030387f
C1196 VTAIL.n215 VSUBS 0.013612f
C1197 VTAIL.n216 VSUBS 0.012856f
C1198 VTAIL.n217 VSUBS 0.023924f
C1199 VTAIL.n218 VSUBS 0.023924f
C1200 VTAIL.n219 VSUBS 0.012856f
C1201 VTAIL.n220 VSUBS 0.013612f
C1202 VTAIL.n221 VSUBS 0.030387f
C1203 VTAIL.n222 VSUBS 0.030387f
C1204 VTAIL.n223 VSUBS 0.013612f
C1205 VTAIL.n224 VSUBS 0.012856f
C1206 VTAIL.n225 VSUBS 0.023924f
C1207 VTAIL.n226 VSUBS 0.023924f
C1208 VTAIL.n227 VSUBS 0.012856f
C1209 VTAIL.n228 VSUBS 0.013612f
C1210 VTAIL.n229 VSUBS 0.030387f
C1211 VTAIL.n230 VSUBS 0.030387f
C1212 VTAIL.n231 VSUBS 0.013612f
C1213 VTAIL.n232 VSUBS 0.012856f
C1214 VTAIL.n233 VSUBS 0.023924f
C1215 VTAIL.n234 VSUBS 0.023924f
C1216 VTAIL.n235 VSUBS 0.012856f
C1217 VTAIL.n236 VSUBS 0.013612f
C1218 VTAIL.n237 VSUBS 0.030387f
C1219 VTAIL.n238 VSUBS 0.030387f
C1220 VTAIL.n239 VSUBS 0.013612f
C1221 VTAIL.n240 VSUBS 0.012856f
C1222 VTAIL.n241 VSUBS 0.023924f
C1223 VTAIL.n242 VSUBS 0.023924f
C1224 VTAIL.n243 VSUBS 0.012856f
C1225 VTAIL.n244 VSUBS 0.012856f
C1226 VTAIL.n245 VSUBS 0.013612f
C1227 VTAIL.n246 VSUBS 0.030387f
C1228 VTAIL.n247 VSUBS 0.030387f
C1229 VTAIL.n248 VSUBS 0.030387f
C1230 VTAIL.n249 VSUBS 0.013234f
C1231 VTAIL.n250 VSUBS 0.012856f
C1232 VTAIL.n251 VSUBS 0.023924f
C1233 VTAIL.n252 VSUBS 0.023924f
C1234 VTAIL.n253 VSUBS 0.012856f
C1235 VTAIL.n254 VSUBS 0.013612f
C1236 VTAIL.n255 VSUBS 0.030387f
C1237 VTAIL.n256 VSUBS 0.069077f
C1238 VTAIL.n257 VSUBS 0.013612f
C1239 VTAIL.n258 VSUBS 0.012856f
C1240 VTAIL.n259 VSUBS 0.056607f
C1241 VTAIL.n260 VSUBS 0.034579f
C1242 VTAIL.n261 VSUBS 1.71915f
C1243 VTAIL.n262 VSUBS 0.024971f
C1244 VTAIL.n263 VSUBS 0.023924f
C1245 VTAIL.n264 VSUBS 0.012856f
C1246 VTAIL.n265 VSUBS 0.030387f
C1247 VTAIL.n266 VSUBS 0.013234f
C1248 VTAIL.n267 VSUBS 0.023924f
C1249 VTAIL.n268 VSUBS 0.013234f
C1250 VTAIL.n269 VSUBS 0.012856f
C1251 VTAIL.n270 VSUBS 0.030387f
C1252 VTAIL.n271 VSUBS 0.030387f
C1253 VTAIL.n272 VSUBS 0.013612f
C1254 VTAIL.n273 VSUBS 0.023924f
C1255 VTAIL.n274 VSUBS 0.012856f
C1256 VTAIL.n275 VSUBS 0.030387f
C1257 VTAIL.n276 VSUBS 0.013612f
C1258 VTAIL.n277 VSUBS 0.023924f
C1259 VTAIL.n278 VSUBS 0.012856f
C1260 VTAIL.n279 VSUBS 0.030387f
C1261 VTAIL.n280 VSUBS 0.013612f
C1262 VTAIL.n281 VSUBS 0.023924f
C1263 VTAIL.n282 VSUBS 0.012856f
C1264 VTAIL.n283 VSUBS 0.030387f
C1265 VTAIL.n284 VSUBS 0.013612f
C1266 VTAIL.n285 VSUBS 0.023924f
C1267 VTAIL.n286 VSUBS 0.012856f
C1268 VTAIL.n287 VSUBS 0.030387f
C1269 VTAIL.n288 VSUBS 0.013612f
C1270 VTAIL.n289 VSUBS 1.57107f
C1271 VTAIL.n290 VSUBS 0.012856f
C1272 VTAIL.t6 VSUBS 0.065076f
C1273 VTAIL.n291 VSUBS 0.171469f
C1274 VTAIL.n292 VSUBS 0.019331f
C1275 VTAIL.n293 VSUBS 0.02279f
C1276 VTAIL.n294 VSUBS 0.030387f
C1277 VTAIL.n295 VSUBS 0.013612f
C1278 VTAIL.n296 VSUBS 0.012856f
C1279 VTAIL.n297 VSUBS 0.023924f
C1280 VTAIL.n298 VSUBS 0.023924f
C1281 VTAIL.n299 VSUBS 0.012856f
C1282 VTAIL.n300 VSUBS 0.013612f
C1283 VTAIL.n301 VSUBS 0.030387f
C1284 VTAIL.n302 VSUBS 0.030387f
C1285 VTAIL.n303 VSUBS 0.013612f
C1286 VTAIL.n304 VSUBS 0.012856f
C1287 VTAIL.n305 VSUBS 0.023924f
C1288 VTAIL.n306 VSUBS 0.023924f
C1289 VTAIL.n307 VSUBS 0.012856f
C1290 VTAIL.n308 VSUBS 0.013612f
C1291 VTAIL.n309 VSUBS 0.030387f
C1292 VTAIL.n310 VSUBS 0.030387f
C1293 VTAIL.n311 VSUBS 0.013612f
C1294 VTAIL.n312 VSUBS 0.012856f
C1295 VTAIL.n313 VSUBS 0.023924f
C1296 VTAIL.n314 VSUBS 0.023924f
C1297 VTAIL.n315 VSUBS 0.012856f
C1298 VTAIL.n316 VSUBS 0.013612f
C1299 VTAIL.n317 VSUBS 0.030387f
C1300 VTAIL.n318 VSUBS 0.030387f
C1301 VTAIL.n319 VSUBS 0.013612f
C1302 VTAIL.n320 VSUBS 0.012856f
C1303 VTAIL.n321 VSUBS 0.023924f
C1304 VTAIL.n322 VSUBS 0.023924f
C1305 VTAIL.n323 VSUBS 0.012856f
C1306 VTAIL.n324 VSUBS 0.013612f
C1307 VTAIL.n325 VSUBS 0.030387f
C1308 VTAIL.n326 VSUBS 0.030387f
C1309 VTAIL.n327 VSUBS 0.013612f
C1310 VTAIL.n328 VSUBS 0.012856f
C1311 VTAIL.n329 VSUBS 0.023924f
C1312 VTAIL.n330 VSUBS 0.023924f
C1313 VTAIL.n331 VSUBS 0.012856f
C1314 VTAIL.n332 VSUBS 0.013612f
C1315 VTAIL.n333 VSUBS 0.030387f
C1316 VTAIL.n334 VSUBS 0.030387f
C1317 VTAIL.n335 VSUBS 0.013612f
C1318 VTAIL.n336 VSUBS 0.012856f
C1319 VTAIL.n337 VSUBS 0.023924f
C1320 VTAIL.n338 VSUBS 0.023924f
C1321 VTAIL.n339 VSUBS 0.012856f
C1322 VTAIL.n340 VSUBS 0.013612f
C1323 VTAIL.n341 VSUBS 0.030387f
C1324 VTAIL.n342 VSUBS 0.069077f
C1325 VTAIL.n343 VSUBS 0.013612f
C1326 VTAIL.n344 VSUBS 0.012856f
C1327 VTAIL.n345 VSUBS 0.056607f
C1328 VTAIL.n346 VSUBS 0.034579f
C1329 VTAIL.n347 VSUBS 1.71915f
C1330 VTAIL.t5 VSUBS 0.291149f
C1331 VTAIL.t7 VSUBS 0.291149f
C1332 VTAIL.n348 VSUBS 2.2342f
C1333 VTAIL.n349 VSUBS 0.914052f
C1334 VTAIL.n350 VSUBS 0.024971f
C1335 VTAIL.n351 VSUBS 0.023924f
C1336 VTAIL.n352 VSUBS 0.012856f
C1337 VTAIL.n353 VSUBS 0.030387f
C1338 VTAIL.n354 VSUBS 0.013234f
C1339 VTAIL.n355 VSUBS 0.023924f
C1340 VTAIL.n356 VSUBS 0.013234f
C1341 VTAIL.n357 VSUBS 0.012856f
C1342 VTAIL.n358 VSUBS 0.030387f
C1343 VTAIL.n359 VSUBS 0.030387f
C1344 VTAIL.n360 VSUBS 0.013612f
C1345 VTAIL.n361 VSUBS 0.023924f
C1346 VTAIL.n362 VSUBS 0.012856f
C1347 VTAIL.n363 VSUBS 0.030387f
C1348 VTAIL.n364 VSUBS 0.013612f
C1349 VTAIL.n365 VSUBS 0.023924f
C1350 VTAIL.n366 VSUBS 0.012856f
C1351 VTAIL.n367 VSUBS 0.030387f
C1352 VTAIL.n368 VSUBS 0.013612f
C1353 VTAIL.n369 VSUBS 0.023924f
C1354 VTAIL.n370 VSUBS 0.012856f
C1355 VTAIL.n371 VSUBS 0.030387f
C1356 VTAIL.n372 VSUBS 0.013612f
C1357 VTAIL.n373 VSUBS 0.023924f
C1358 VTAIL.n374 VSUBS 0.012856f
C1359 VTAIL.n375 VSUBS 0.030387f
C1360 VTAIL.n376 VSUBS 0.013612f
C1361 VTAIL.n377 VSUBS 1.57107f
C1362 VTAIL.n378 VSUBS 0.012856f
C1363 VTAIL.t4 VSUBS 0.065076f
C1364 VTAIL.n379 VSUBS 0.171469f
C1365 VTAIL.n380 VSUBS 0.019331f
C1366 VTAIL.n381 VSUBS 0.02279f
C1367 VTAIL.n382 VSUBS 0.030387f
C1368 VTAIL.n383 VSUBS 0.013612f
C1369 VTAIL.n384 VSUBS 0.012856f
C1370 VTAIL.n385 VSUBS 0.023924f
C1371 VTAIL.n386 VSUBS 0.023924f
C1372 VTAIL.n387 VSUBS 0.012856f
C1373 VTAIL.n388 VSUBS 0.013612f
C1374 VTAIL.n389 VSUBS 0.030387f
C1375 VTAIL.n390 VSUBS 0.030387f
C1376 VTAIL.n391 VSUBS 0.013612f
C1377 VTAIL.n392 VSUBS 0.012856f
C1378 VTAIL.n393 VSUBS 0.023924f
C1379 VTAIL.n394 VSUBS 0.023924f
C1380 VTAIL.n395 VSUBS 0.012856f
C1381 VTAIL.n396 VSUBS 0.013612f
C1382 VTAIL.n397 VSUBS 0.030387f
C1383 VTAIL.n398 VSUBS 0.030387f
C1384 VTAIL.n399 VSUBS 0.013612f
C1385 VTAIL.n400 VSUBS 0.012856f
C1386 VTAIL.n401 VSUBS 0.023924f
C1387 VTAIL.n402 VSUBS 0.023924f
C1388 VTAIL.n403 VSUBS 0.012856f
C1389 VTAIL.n404 VSUBS 0.013612f
C1390 VTAIL.n405 VSUBS 0.030387f
C1391 VTAIL.n406 VSUBS 0.030387f
C1392 VTAIL.n407 VSUBS 0.013612f
C1393 VTAIL.n408 VSUBS 0.012856f
C1394 VTAIL.n409 VSUBS 0.023924f
C1395 VTAIL.n410 VSUBS 0.023924f
C1396 VTAIL.n411 VSUBS 0.012856f
C1397 VTAIL.n412 VSUBS 0.013612f
C1398 VTAIL.n413 VSUBS 0.030387f
C1399 VTAIL.n414 VSUBS 0.030387f
C1400 VTAIL.n415 VSUBS 0.013612f
C1401 VTAIL.n416 VSUBS 0.012856f
C1402 VTAIL.n417 VSUBS 0.023924f
C1403 VTAIL.n418 VSUBS 0.023924f
C1404 VTAIL.n419 VSUBS 0.012856f
C1405 VTAIL.n420 VSUBS 0.013612f
C1406 VTAIL.n421 VSUBS 0.030387f
C1407 VTAIL.n422 VSUBS 0.030387f
C1408 VTAIL.n423 VSUBS 0.013612f
C1409 VTAIL.n424 VSUBS 0.012856f
C1410 VTAIL.n425 VSUBS 0.023924f
C1411 VTAIL.n426 VSUBS 0.023924f
C1412 VTAIL.n427 VSUBS 0.012856f
C1413 VTAIL.n428 VSUBS 0.013612f
C1414 VTAIL.n429 VSUBS 0.030387f
C1415 VTAIL.n430 VSUBS 0.069077f
C1416 VTAIL.n431 VSUBS 0.013612f
C1417 VTAIL.n432 VSUBS 0.012856f
C1418 VTAIL.n433 VSUBS 0.056607f
C1419 VTAIL.n434 VSUBS 0.034579f
C1420 VTAIL.n435 VSUBS 0.232172f
C1421 VTAIL.n436 VSUBS 0.024971f
C1422 VTAIL.n437 VSUBS 0.023924f
C1423 VTAIL.n438 VSUBS 0.012856f
C1424 VTAIL.n439 VSUBS 0.030387f
C1425 VTAIL.n440 VSUBS 0.013234f
C1426 VTAIL.n441 VSUBS 0.023924f
C1427 VTAIL.n442 VSUBS 0.013234f
C1428 VTAIL.n443 VSUBS 0.012856f
C1429 VTAIL.n444 VSUBS 0.030387f
C1430 VTAIL.n445 VSUBS 0.030387f
C1431 VTAIL.n446 VSUBS 0.013612f
C1432 VTAIL.n447 VSUBS 0.023924f
C1433 VTAIL.n448 VSUBS 0.012856f
C1434 VTAIL.n449 VSUBS 0.030387f
C1435 VTAIL.n450 VSUBS 0.013612f
C1436 VTAIL.n451 VSUBS 0.023924f
C1437 VTAIL.n452 VSUBS 0.012856f
C1438 VTAIL.n453 VSUBS 0.030387f
C1439 VTAIL.n454 VSUBS 0.013612f
C1440 VTAIL.n455 VSUBS 0.023924f
C1441 VTAIL.n456 VSUBS 0.012856f
C1442 VTAIL.n457 VSUBS 0.030387f
C1443 VTAIL.n458 VSUBS 0.013612f
C1444 VTAIL.n459 VSUBS 0.023924f
C1445 VTAIL.n460 VSUBS 0.012856f
C1446 VTAIL.n461 VSUBS 0.030387f
C1447 VTAIL.n462 VSUBS 0.013612f
C1448 VTAIL.n463 VSUBS 1.57107f
C1449 VTAIL.n464 VSUBS 0.012856f
C1450 VTAIL.t11 VSUBS 0.065076f
C1451 VTAIL.n465 VSUBS 0.171469f
C1452 VTAIL.n466 VSUBS 0.019331f
C1453 VTAIL.n467 VSUBS 0.02279f
C1454 VTAIL.n468 VSUBS 0.030387f
C1455 VTAIL.n469 VSUBS 0.013612f
C1456 VTAIL.n470 VSUBS 0.012856f
C1457 VTAIL.n471 VSUBS 0.023924f
C1458 VTAIL.n472 VSUBS 0.023924f
C1459 VTAIL.n473 VSUBS 0.012856f
C1460 VTAIL.n474 VSUBS 0.013612f
C1461 VTAIL.n475 VSUBS 0.030387f
C1462 VTAIL.n476 VSUBS 0.030387f
C1463 VTAIL.n477 VSUBS 0.013612f
C1464 VTAIL.n478 VSUBS 0.012856f
C1465 VTAIL.n479 VSUBS 0.023924f
C1466 VTAIL.n480 VSUBS 0.023924f
C1467 VTAIL.n481 VSUBS 0.012856f
C1468 VTAIL.n482 VSUBS 0.013612f
C1469 VTAIL.n483 VSUBS 0.030387f
C1470 VTAIL.n484 VSUBS 0.030387f
C1471 VTAIL.n485 VSUBS 0.013612f
C1472 VTAIL.n486 VSUBS 0.012856f
C1473 VTAIL.n487 VSUBS 0.023924f
C1474 VTAIL.n488 VSUBS 0.023924f
C1475 VTAIL.n489 VSUBS 0.012856f
C1476 VTAIL.n490 VSUBS 0.013612f
C1477 VTAIL.n491 VSUBS 0.030387f
C1478 VTAIL.n492 VSUBS 0.030387f
C1479 VTAIL.n493 VSUBS 0.013612f
C1480 VTAIL.n494 VSUBS 0.012856f
C1481 VTAIL.n495 VSUBS 0.023924f
C1482 VTAIL.n496 VSUBS 0.023924f
C1483 VTAIL.n497 VSUBS 0.012856f
C1484 VTAIL.n498 VSUBS 0.013612f
C1485 VTAIL.n499 VSUBS 0.030387f
C1486 VTAIL.n500 VSUBS 0.030387f
C1487 VTAIL.n501 VSUBS 0.013612f
C1488 VTAIL.n502 VSUBS 0.012856f
C1489 VTAIL.n503 VSUBS 0.023924f
C1490 VTAIL.n504 VSUBS 0.023924f
C1491 VTAIL.n505 VSUBS 0.012856f
C1492 VTAIL.n506 VSUBS 0.013612f
C1493 VTAIL.n507 VSUBS 0.030387f
C1494 VTAIL.n508 VSUBS 0.030387f
C1495 VTAIL.n509 VSUBS 0.013612f
C1496 VTAIL.n510 VSUBS 0.012856f
C1497 VTAIL.n511 VSUBS 0.023924f
C1498 VTAIL.n512 VSUBS 0.023924f
C1499 VTAIL.n513 VSUBS 0.012856f
C1500 VTAIL.n514 VSUBS 0.013612f
C1501 VTAIL.n515 VSUBS 0.030387f
C1502 VTAIL.n516 VSUBS 0.069077f
C1503 VTAIL.n517 VSUBS 0.013612f
C1504 VTAIL.n518 VSUBS 0.012856f
C1505 VTAIL.n519 VSUBS 0.056607f
C1506 VTAIL.n520 VSUBS 0.034579f
C1507 VTAIL.n521 VSUBS 0.232172f
C1508 VTAIL.t8 VSUBS 0.291149f
C1509 VTAIL.t13 VSUBS 0.291149f
C1510 VTAIL.n522 VSUBS 2.2342f
C1511 VTAIL.n523 VSUBS 0.914052f
C1512 VTAIL.n524 VSUBS 0.024971f
C1513 VTAIL.n525 VSUBS 0.023924f
C1514 VTAIL.n526 VSUBS 0.012856f
C1515 VTAIL.n527 VSUBS 0.030387f
C1516 VTAIL.n528 VSUBS 0.013234f
C1517 VTAIL.n529 VSUBS 0.023924f
C1518 VTAIL.n530 VSUBS 0.013234f
C1519 VTAIL.n531 VSUBS 0.012856f
C1520 VTAIL.n532 VSUBS 0.030387f
C1521 VTAIL.n533 VSUBS 0.030387f
C1522 VTAIL.n534 VSUBS 0.013612f
C1523 VTAIL.n535 VSUBS 0.023924f
C1524 VTAIL.n536 VSUBS 0.012856f
C1525 VTAIL.n537 VSUBS 0.030387f
C1526 VTAIL.n538 VSUBS 0.013612f
C1527 VTAIL.n539 VSUBS 0.023924f
C1528 VTAIL.n540 VSUBS 0.012856f
C1529 VTAIL.n541 VSUBS 0.030387f
C1530 VTAIL.n542 VSUBS 0.013612f
C1531 VTAIL.n543 VSUBS 0.023924f
C1532 VTAIL.n544 VSUBS 0.012856f
C1533 VTAIL.n545 VSUBS 0.030387f
C1534 VTAIL.n546 VSUBS 0.013612f
C1535 VTAIL.n547 VSUBS 0.023924f
C1536 VTAIL.n548 VSUBS 0.012856f
C1537 VTAIL.n549 VSUBS 0.030387f
C1538 VTAIL.n550 VSUBS 0.013612f
C1539 VTAIL.n551 VSUBS 1.57107f
C1540 VTAIL.n552 VSUBS 0.012856f
C1541 VTAIL.t14 VSUBS 0.065076f
C1542 VTAIL.n553 VSUBS 0.171469f
C1543 VTAIL.n554 VSUBS 0.019331f
C1544 VTAIL.n555 VSUBS 0.02279f
C1545 VTAIL.n556 VSUBS 0.030387f
C1546 VTAIL.n557 VSUBS 0.013612f
C1547 VTAIL.n558 VSUBS 0.012856f
C1548 VTAIL.n559 VSUBS 0.023924f
C1549 VTAIL.n560 VSUBS 0.023924f
C1550 VTAIL.n561 VSUBS 0.012856f
C1551 VTAIL.n562 VSUBS 0.013612f
C1552 VTAIL.n563 VSUBS 0.030387f
C1553 VTAIL.n564 VSUBS 0.030387f
C1554 VTAIL.n565 VSUBS 0.013612f
C1555 VTAIL.n566 VSUBS 0.012856f
C1556 VTAIL.n567 VSUBS 0.023924f
C1557 VTAIL.n568 VSUBS 0.023924f
C1558 VTAIL.n569 VSUBS 0.012856f
C1559 VTAIL.n570 VSUBS 0.013612f
C1560 VTAIL.n571 VSUBS 0.030387f
C1561 VTAIL.n572 VSUBS 0.030387f
C1562 VTAIL.n573 VSUBS 0.013612f
C1563 VTAIL.n574 VSUBS 0.012856f
C1564 VTAIL.n575 VSUBS 0.023924f
C1565 VTAIL.n576 VSUBS 0.023924f
C1566 VTAIL.n577 VSUBS 0.012856f
C1567 VTAIL.n578 VSUBS 0.013612f
C1568 VTAIL.n579 VSUBS 0.030387f
C1569 VTAIL.n580 VSUBS 0.030387f
C1570 VTAIL.n581 VSUBS 0.013612f
C1571 VTAIL.n582 VSUBS 0.012856f
C1572 VTAIL.n583 VSUBS 0.023924f
C1573 VTAIL.n584 VSUBS 0.023924f
C1574 VTAIL.n585 VSUBS 0.012856f
C1575 VTAIL.n586 VSUBS 0.013612f
C1576 VTAIL.n587 VSUBS 0.030387f
C1577 VTAIL.n588 VSUBS 0.030387f
C1578 VTAIL.n589 VSUBS 0.013612f
C1579 VTAIL.n590 VSUBS 0.012856f
C1580 VTAIL.n591 VSUBS 0.023924f
C1581 VTAIL.n592 VSUBS 0.023924f
C1582 VTAIL.n593 VSUBS 0.012856f
C1583 VTAIL.n594 VSUBS 0.013612f
C1584 VTAIL.n595 VSUBS 0.030387f
C1585 VTAIL.n596 VSUBS 0.030387f
C1586 VTAIL.n597 VSUBS 0.013612f
C1587 VTAIL.n598 VSUBS 0.012856f
C1588 VTAIL.n599 VSUBS 0.023924f
C1589 VTAIL.n600 VSUBS 0.023924f
C1590 VTAIL.n601 VSUBS 0.012856f
C1591 VTAIL.n602 VSUBS 0.013612f
C1592 VTAIL.n603 VSUBS 0.030387f
C1593 VTAIL.n604 VSUBS 0.069077f
C1594 VTAIL.n605 VSUBS 0.013612f
C1595 VTAIL.n606 VSUBS 0.012856f
C1596 VTAIL.n607 VSUBS 0.056607f
C1597 VTAIL.n608 VSUBS 0.034579f
C1598 VTAIL.n609 VSUBS 1.71915f
C1599 VTAIL.n610 VSUBS 0.024971f
C1600 VTAIL.n611 VSUBS 0.023924f
C1601 VTAIL.n612 VSUBS 0.012856f
C1602 VTAIL.n613 VSUBS 0.030387f
C1603 VTAIL.n614 VSUBS 0.013234f
C1604 VTAIL.n615 VSUBS 0.023924f
C1605 VTAIL.n616 VSUBS 0.013612f
C1606 VTAIL.n617 VSUBS 0.030387f
C1607 VTAIL.n618 VSUBS 0.013612f
C1608 VTAIL.n619 VSUBS 0.023924f
C1609 VTAIL.n620 VSUBS 0.012856f
C1610 VTAIL.n621 VSUBS 0.030387f
C1611 VTAIL.n622 VSUBS 0.013612f
C1612 VTAIL.n623 VSUBS 0.023924f
C1613 VTAIL.n624 VSUBS 0.012856f
C1614 VTAIL.n625 VSUBS 0.030387f
C1615 VTAIL.n626 VSUBS 0.013612f
C1616 VTAIL.n627 VSUBS 0.023924f
C1617 VTAIL.n628 VSUBS 0.012856f
C1618 VTAIL.n629 VSUBS 0.030387f
C1619 VTAIL.n630 VSUBS 0.013612f
C1620 VTAIL.n631 VSUBS 0.023924f
C1621 VTAIL.n632 VSUBS 0.012856f
C1622 VTAIL.n633 VSUBS 0.030387f
C1623 VTAIL.n634 VSUBS 0.013612f
C1624 VTAIL.n635 VSUBS 1.57107f
C1625 VTAIL.n636 VSUBS 0.012856f
C1626 VTAIL.t0 VSUBS 0.065076f
C1627 VTAIL.n637 VSUBS 0.171469f
C1628 VTAIL.n638 VSUBS 0.019331f
C1629 VTAIL.n639 VSUBS 0.02279f
C1630 VTAIL.n640 VSUBS 0.030387f
C1631 VTAIL.n641 VSUBS 0.013612f
C1632 VTAIL.n642 VSUBS 0.012856f
C1633 VTAIL.n643 VSUBS 0.023924f
C1634 VTAIL.n644 VSUBS 0.023924f
C1635 VTAIL.n645 VSUBS 0.012856f
C1636 VTAIL.n646 VSUBS 0.013612f
C1637 VTAIL.n647 VSUBS 0.030387f
C1638 VTAIL.n648 VSUBS 0.030387f
C1639 VTAIL.n649 VSUBS 0.013612f
C1640 VTAIL.n650 VSUBS 0.012856f
C1641 VTAIL.n651 VSUBS 0.023924f
C1642 VTAIL.n652 VSUBS 0.023924f
C1643 VTAIL.n653 VSUBS 0.012856f
C1644 VTAIL.n654 VSUBS 0.013612f
C1645 VTAIL.n655 VSUBS 0.030387f
C1646 VTAIL.n656 VSUBS 0.030387f
C1647 VTAIL.n657 VSUBS 0.013612f
C1648 VTAIL.n658 VSUBS 0.012856f
C1649 VTAIL.n659 VSUBS 0.023924f
C1650 VTAIL.n660 VSUBS 0.023924f
C1651 VTAIL.n661 VSUBS 0.012856f
C1652 VTAIL.n662 VSUBS 0.013612f
C1653 VTAIL.n663 VSUBS 0.030387f
C1654 VTAIL.n664 VSUBS 0.030387f
C1655 VTAIL.n665 VSUBS 0.013612f
C1656 VTAIL.n666 VSUBS 0.012856f
C1657 VTAIL.n667 VSUBS 0.023924f
C1658 VTAIL.n668 VSUBS 0.023924f
C1659 VTAIL.n669 VSUBS 0.012856f
C1660 VTAIL.n670 VSUBS 0.013612f
C1661 VTAIL.n671 VSUBS 0.030387f
C1662 VTAIL.n672 VSUBS 0.030387f
C1663 VTAIL.n673 VSUBS 0.013612f
C1664 VTAIL.n674 VSUBS 0.012856f
C1665 VTAIL.n675 VSUBS 0.023924f
C1666 VTAIL.n676 VSUBS 0.023924f
C1667 VTAIL.n677 VSUBS 0.012856f
C1668 VTAIL.n678 VSUBS 0.012856f
C1669 VTAIL.n679 VSUBS 0.013612f
C1670 VTAIL.n680 VSUBS 0.030387f
C1671 VTAIL.n681 VSUBS 0.030387f
C1672 VTAIL.n682 VSUBS 0.030387f
C1673 VTAIL.n683 VSUBS 0.013234f
C1674 VTAIL.n684 VSUBS 0.012856f
C1675 VTAIL.n685 VSUBS 0.023924f
C1676 VTAIL.n686 VSUBS 0.023924f
C1677 VTAIL.n687 VSUBS 0.012856f
C1678 VTAIL.n688 VSUBS 0.013612f
C1679 VTAIL.n689 VSUBS 0.030387f
C1680 VTAIL.n690 VSUBS 0.069077f
C1681 VTAIL.n691 VSUBS 0.013612f
C1682 VTAIL.n692 VSUBS 0.012856f
C1683 VTAIL.n693 VSUBS 0.056607f
C1684 VTAIL.n694 VSUBS 0.034579f
C1685 VTAIL.n695 VSUBS 1.71467f
C1686 VP.n0 VSUBS 0.03926f
C1687 VP.t0 VSUBS 2.89211f
C1688 VP.n1 VSUBS 0.030008f
C1689 VP.n2 VSUBS 0.02978f
C1690 VP.t2 VSUBS 2.89211f
C1691 VP.n3 VSUBS 0.055225f
C1692 VP.n4 VSUBS 0.02978f
C1693 VP.n5 VSUBS 0.031506f
C1694 VP.n6 VSUBS 0.02978f
C1695 VP.n7 VSUBS 0.058591f
C1696 VP.n8 VSUBS 0.03926f
C1697 VP.t4 VSUBS 2.89211f
C1698 VP.n9 VSUBS 0.030008f
C1699 VP.n10 VSUBS 0.02978f
C1700 VP.t6 VSUBS 2.89211f
C1701 VP.n11 VSUBS 0.055225f
C1702 VP.n12 VSUBS 0.02978f
C1703 VP.n13 VSUBS 0.031506f
C1704 VP.t7 VSUBS 3.07989f
C1705 VP.t5 VSUBS 2.89211f
C1706 VP.n14 VSUBS 1.08276f
C1707 VP.n15 VSUBS 1.08271f
C1708 VP.n16 VSUBS 0.255988f
C1709 VP.n17 VSUBS 0.02978f
C1710 VP.n18 VSUBS 0.055225f
C1711 VP.n19 VSUBS 0.04329f
C1712 VP.n20 VSUBS 0.04329f
C1713 VP.n21 VSUBS 0.02978f
C1714 VP.n22 VSUBS 0.02978f
C1715 VP.n23 VSUBS 0.02978f
C1716 VP.n24 VSUBS 0.031506f
C1717 VP.n25 VSUBS 1.01263f
C1718 VP.n26 VSUBS 0.051681f
C1719 VP.n27 VSUBS 0.053206f
C1720 VP.n28 VSUBS 0.02978f
C1721 VP.n29 VSUBS 0.02978f
C1722 VP.n30 VSUBS 0.02978f
C1723 VP.n31 VSUBS 0.058591f
C1724 VP.n32 VSUBS 0.038594f
C1725 VP.n33 VSUBS 1.0991f
C1726 VP.n34 VSUBS 1.75087f
C1727 VP.n35 VSUBS 1.77151f
C1728 VP.t3 VSUBS 2.89211f
C1729 VP.n36 VSUBS 1.0991f
C1730 VP.n37 VSUBS 0.038594f
C1731 VP.n38 VSUBS 0.03926f
C1732 VP.n39 VSUBS 0.02978f
C1733 VP.n40 VSUBS 0.02978f
C1734 VP.n41 VSUBS 0.030008f
C1735 VP.n42 VSUBS 0.053206f
C1736 VP.t1 VSUBS 2.89211f
C1737 VP.n43 VSUBS 1.01263f
C1738 VP.n44 VSUBS 0.051681f
C1739 VP.n45 VSUBS 0.02978f
C1740 VP.n46 VSUBS 0.02978f
C1741 VP.n47 VSUBS 0.02978f
C1742 VP.n48 VSUBS 0.055225f
C1743 VP.n49 VSUBS 0.04329f
C1744 VP.n50 VSUBS 0.04329f
C1745 VP.n51 VSUBS 0.02978f
C1746 VP.n52 VSUBS 0.02978f
C1747 VP.n53 VSUBS 0.02978f
C1748 VP.n54 VSUBS 0.031506f
C1749 VP.n55 VSUBS 1.01263f
C1750 VP.n56 VSUBS 0.051681f
C1751 VP.n57 VSUBS 0.053206f
C1752 VP.n58 VSUBS 0.02978f
C1753 VP.n59 VSUBS 0.02978f
C1754 VP.n60 VSUBS 0.02978f
C1755 VP.n61 VSUBS 0.058591f
C1756 VP.n62 VSUBS 0.038594f
C1757 VP.n63 VSUBS 1.0991f
C1758 VP.n64 VSUBS 0.045943f
.ends

