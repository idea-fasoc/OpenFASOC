* NGSPICE file created from diff_pair_sample_0338.ext - technology: sky130A

.subckt diff_pair_sample_0338 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t4 w_n3946_n2290# sky130_fd_pr__pfet_01v8 ad=1.09065 pd=6.94 as=1.09065 ps=6.94 w=6.61 l=3.39
X1 VTAIL.t4 VP.t0 VDD1.t5 w_n3946_n2290# sky130_fd_pr__pfet_01v8 ad=1.09065 pd=6.94 as=1.09065 ps=6.94 w=6.61 l=3.39
X2 VDD1.t4 VP.t1 VTAIL.t3 w_n3946_n2290# sky130_fd_pr__pfet_01v8 ad=2.5779 pd=14 as=1.09065 ps=6.94 w=6.61 l=3.39
X3 B.t11 B.t9 B.t10 w_n3946_n2290# sky130_fd_pr__pfet_01v8 ad=2.5779 pd=14 as=0 ps=0 w=6.61 l=3.39
X4 B.t8 B.t6 B.t7 w_n3946_n2290# sky130_fd_pr__pfet_01v8 ad=2.5779 pd=14 as=0 ps=0 w=6.61 l=3.39
X5 VDD2.t0 VN.t1 VTAIL.t10 w_n3946_n2290# sky130_fd_pr__pfet_01v8 ad=1.09065 pd=6.94 as=2.5779 ps=14 w=6.61 l=3.39
X6 B.t5 B.t3 B.t4 w_n3946_n2290# sky130_fd_pr__pfet_01v8 ad=2.5779 pd=14 as=0 ps=0 w=6.61 l=3.39
X7 VDD1.t3 VP.t2 VTAIL.t0 w_n3946_n2290# sky130_fd_pr__pfet_01v8 ad=2.5779 pd=14 as=1.09065 ps=6.94 w=6.61 l=3.39
X8 VDD2.t2 VN.t2 VTAIL.t9 w_n3946_n2290# sky130_fd_pr__pfet_01v8 ad=1.09065 pd=6.94 as=2.5779 ps=14 w=6.61 l=3.39
X9 VDD1.t2 VP.t3 VTAIL.t5 w_n3946_n2290# sky130_fd_pr__pfet_01v8 ad=1.09065 pd=6.94 as=2.5779 ps=14 w=6.61 l=3.39
X10 VTAIL.t8 VN.t3 VDD2.t5 w_n3946_n2290# sky130_fd_pr__pfet_01v8 ad=1.09065 pd=6.94 as=1.09065 ps=6.94 w=6.61 l=3.39
X11 B.t2 B.t0 B.t1 w_n3946_n2290# sky130_fd_pr__pfet_01v8 ad=2.5779 pd=14 as=0 ps=0 w=6.61 l=3.39
X12 VDD2.t3 VN.t4 VTAIL.t7 w_n3946_n2290# sky130_fd_pr__pfet_01v8 ad=2.5779 pd=14 as=1.09065 ps=6.94 w=6.61 l=3.39
X13 VDD1.t1 VP.t4 VTAIL.t2 w_n3946_n2290# sky130_fd_pr__pfet_01v8 ad=1.09065 pd=6.94 as=2.5779 ps=14 w=6.61 l=3.39
X14 VTAIL.t1 VP.t5 VDD1.t0 w_n3946_n2290# sky130_fd_pr__pfet_01v8 ad=1.09065 pd=6.94 as=1.09065 ps=6.94 w=6.61 l=3.39
X15 VDD2.t1 VN.t5 VTAIL.t6 w_n3946_n2290# sky130_fd_pr__pfet_01v8 ad=2.5779 pd=14 as=1.09065 ps=6.94 w=6.61 l=3.39
R0 VN.n34 VN.n33 161.3
R1 VN.n32 VN.n19 161.3
R2 VN.n31 VN.n30 161.3
R3 VN.n29 VN.n20 161.3
R4 VN.n28 VN.n27 161.3
R5 VN.n26 VN.n21 161.3
R6 VN.n25 VN.n24 161.3
R7 VN.n16 VN.n15 161.3
R8 VN.n14 VN.n1 161.3
R9 VN.n13 VN.n12 161.3
R10 VN.n11 VN.n2 161.3
R11 VN.n10 VN.n9 161.3
R12 VN.n8 VN.n3 161.3
R13 VN.n7 VN.n6 161.3
R14 VN.n23 VN.t2 80.5478
R15 VN.n5 VN.t4 80.5478
R16 VN.n17 VN.n0 79.3019
R17 VN.n35 VN.n18 79.3019
R18 VN.n9 VN.n2 54.0911
R19 VN.n27 VN.n20 54.0911
R20 VN.n23 VN.n22 50.1285
R21 VN.n5 VN.n4 50.1285
R22 VN VN.n35 47.9298
R23 VN.n4 VN.t3 46.9919
R24 VN.n0 VN.t1 46.9919
R25 VN.n22 VN.t0 46.9919
R26 VN.n18 VN.t5 46.9919
R27 VN.n13 VN.n2 26.8957
R28 VN.n31 VN.n20 26.8957
R29 VN.n7 VN.n4 24.4675
R30 VN.n8 VN.n7 24.4675
R31 VN.n9 VN.n8 24.4675
R32 VN.n14 VN.n13 24.4675
R33 VN.n15 VN.n14 24.4675
R34 VN.n27 VN.n26 24.4675
R35 VN.n26 VN.n25 24.4675
R36 VN.n25 VN.n22 24.4675
R37 VN.n33 VN.n32 24.4675
R38 VN.n32 VN.n31 24.4675
R39 VN.n15 VN.n0 10.766
R40 VN.n33 VN.n18 10.766
R41 VN.n24 VN.n23 3.12711
R42 VN.n6 VN.n5 3.12711
R43 VN.n35 VN.n34 0.354971
R44 VN.n17 VN.n16 0.354971
R45 VN VN.n17 0.26696
R46 VN.n34 VN.n19 0.189894
R47 VN.n30 VN.n19 0.189894
R48 VN.n30 VN.n29 0.189894
R49 VN.n29 VN.n28 0.189894
R50 VN.n28 VN.n21 0.189894
R51 VN.n24 VN.n21 0.189894
R52 VN.n6 VN.n3 0.189894
R53 VN.n10 VN.n3 0.189894
R54 VN.n11 VN.n10 0.189894
R55 VN.n12 VN.n11 0.189894
R56 VN.n12 VN.n1 0.189894
R57 VN.n16 VN.n1 0.189894
R58 VDD2.n67 VDD2.n37 756.745
R59 VDD2.n30 VDD2.n0 756.745
R60 VDD2.n68 VDD2.n67 585
R61 VDD2.n66 VDD2.n65 585
R62 VDD2.n41 VDD2.n40 585
R63 VDD2.n60 VDD2.n59 585
R64 VDD2.n58 VDD2.n57 585
R65 VDD2.n45 VDD2.n44 585
R66 VDD2.n52 VDD2.n51 585
R67 VDD2.n50 VDD2.n49 585
R68 VDD2.n13 VDD2.n12 585
R69 VDD2.n15 VDD2.n14 585
R70 VDD2.n8 VDD2.n7 585
R71 VDD2.n21 VDD2.n20 585
R72 VDD2.n23 VDD2.n22 585
R73 VDD2.n4 VDD2.n3 585
R74 VDD2.n29 VDD2.n28 585
R75 VDD2.n31 VDD2.n30 585
R76 VDD2.n48 VDD2.t1 327.514
R77 VDD2.n11 VDD2.t3 327.514
R78 VDD2.n67 VDD2.n66 171.744
R79 VDD2.n66 VDD2.n40 171.744
R80 VDD2.n59 VDD2.n40 171.744
R81 VDD2.n59 VDD2.n58 171.744
R82 VDD2.n58 VDD2.n44 171.744
R83 VDD2.n51 VDD2.n44 171.744
R84 VDD2.n51 VDD2.n50 171.744
R85 VDD2.n14 VDD2.n13 171.744
R86 VDD2.n14 VDD2.n7 171.744
R87 VDD2.n21 VDD2.n7 171.744
R88 VDD2.n22 VDD2.n21 171.744
R89 VDD2.n22 VDD2.n3 171.744
R90 VDD2.n29 VDD2.n3 171.744
R91 VDD2.n30 VDD2.n29 171.744
R92 VDD2.n36 VDD2.n35 87.0118
R93 VDD2 VDD2.n73 87.009
R94 VDD2.n50 VDD2.t1 85.8723
R95 VDD2.n13 VDD2.t3 85.8723
R96 VDD2.n36 VDD2.n34 49.0806
R97 VDD2.n72 VDD2.n71 46.7308
R98 VDD2.n72 VDD2.n36 39.836
R99 VDD2.n12 VDD2.n11 16.3884
R100 VDD2.n49 VDD2.n48 16.3884
R101 VDD2.n52 VDD2.n47 12.8005
R102 VDD2.n15 VDD2.n10 12.8005
R103 VDD2.n53 VDD2.n45 12.0247
R104 VDD2.n16 VDD2.n8 12.0247
R105 VDD2.n57 VDD2.n56 11.249
R106 VDD2.n20 VDD2.n19 11.249
R107 VDD2.n60 VDD2.n43 10.4732
R108 VDD2.n23 VDD2.n6 10.4732
R109 VDD2.n61 VDD2.n41 9.69747
R110 VDD2.n24 VDD2.n4 9.69747
R111 VDD2.n71 VDD2.n70 9.45567
R112 VDD2.n34 VDD2.n33 9.45567
R113 VDD2.n70 VDD2.n69 9.3005
R114 VDD2.n39 VDD2.n38 9.3005
R115 VDD2.n64 VDD2.n63 9.3005
R116 VDD2.n62 VDD2.n61 9.3005
R117 VDD2.n43 VDD2.n42 9.3005
R118 VDD2.n56 VDD2.n55 9.3005
R119 VDD2.n54 VDD2.n53 9.3005
R120 VDD2.n47 VDD2.n46 9.3005
R121 VDD2.n2 VDD2.n1 9.3005
R122 VDD2.n27 VDD2.n26 9.3005
R123 VDD2.n25 VDD2.n24 9.3005
R124 VDD2.n6 VDD2.n5 9.3005
R125 VDD2.n19 VDD2.n18 9.3005
R126 VDD2.n17 VDD2.n16 9.3005
R127 VDD2.n10 VDD2.n9 9.3005
R128 VDD2.n33 VDD2.n32 9.3005
R129 VDD2.n65 VDD2.n64 8.92171
R130 VDD2.n28 VDD2.n27 8.92171
R131 VDD2.n68 VDD2.n39 8.14595
R132 VDD2.n31 VDD2.n2 8.14595
R133 VDD2.n69 VDD2.n37 7.3702
R134 VDD2.n32 VDD2.n0 7.3702
R135 VDD2.n71 VDD2.n37 6.59444
R136 VDD2.n34 VDD2.n0 6.59444
R137 VDD2.n69 VDD2.n68 5.81868
R138 VDD2.n32 VDD2.n31 5.81868
R139 VDD2.n65 VDD2.n39 5.04292
R140 VDD2.n28 VDD2.n2 5.04292
R141 VDD2.n73 VDD2.t4 4.91805
R142 VDD2.n73 VDD2.t2 4.91805
R143 VDD2.n35 VDD2.t5 4.91805
R144 VDD2.n35 VDD2.t0 4.91805
R145 VDD2.n64 VDD2.n41 4.26717
R146 VDD2.n27 VDD2.n4 4.26717
R147 VDD2.n48 VDD2.n46 3.71088
R148 VDD2.n11 VDD2.n9 3.71088
R149 VDD2.n61 VDD2.n60 3.49141
R150 VDD2.n24 VDD2.n23 3.49141
R151 VDD2.n57 VDD2.n43 2.71565
R152 VDD2.n20 VDD2.n6 2.71565
R153 VDD2 VDD2.n72 2.46386
R154 VDD2.n56 VDD2.n45 1.93989
R155 VDD2.n19 VDD2.n8 1.93989
R156 VDD2.n53 VDD2.n52 1.16414
R157 VDD2.n16 VDD2.n15 1.16414
R158 VDD2.n49 VDD2.n47 0.388379
R159 VDD2.n12 VDD2.n10 0.388379
R160 VDD2.n70 VDD2.n38 0.155672
R161 VDD2.n63 VDD2.n38 0.155672
R162 VDD2.n63 VDD2.n62 0.155672
R163 VDD2.n62 VDD2.n42 0.155672
R164 VDD2.n55 VDD2.n42 0.155672
R165 VDD2.n55 VDD2.n54 0.155672
R166 VDD2.n54 VDD2.n46 0.155672
R167 VDD2.n17 VDD2.n9 0.155672
R168 VDD2.n18 VDD2.n17 0.155672
R169 VDD2.n18 VDD2.n5 0.155672
R170 VDD2.n25 VDD2.n5 0.155672
R171 VDD2.n26 VDD2.n25 0.155672
R172 VDD2.n26 VDD2.n1 0.155672
R173 VDD2.n33 VDD2.n1 0.155672
R174 VTAIL.n146 VTAIL.n116 756.745
R175 VTAIL.n32 VTAIL.n2 756.745
R176 VTAIL.n110 VTAIL.n80 756.745
R177 VTAIL.n72 VTAIL.n42 756.745
R178 VTAIL.n129 VTAIL.n128 585
R179 VTAIL.n131 VTAIL.n130 585
R180 VTAIL.n124 VTAIL.n123 585
R181 VTAIL.n137 VTAIL.n136 585
R182 VTAIL.n139 VTAIL.n138 585
R183 VTAIL.n120 VTAIL.n119 585
R184 VTAIL.n145 VTAIL.n144 585
R185 VTAIL.n147 VTAIL.n146 585
R186 VTAIL.n15 VTAIL.n14 585
R187 VTAIL.n17 VTAIL.n16 585
R188 VTAIL.n10 VTAIL.n9 585
R189 VTAIL.n23 VTAIL.n22 585
R190 VTAIL.n25 VTAIL.n24 585
R191 VTAIL.n6 VTAIL.n5 585
R192 VTAIL.n31 VTAIL.n30 585
R193 VTAIL.n33 VTAIL.n32 585
R194 VTAIL.n111 VTAIL.n110 585
R195 VTAIL.n109 VTAIL.n108 585
R196 VTAIL.n84 VTAIL.n83 585
R197 VTAIL.n103 VTAIL.n102 585
R198 VTAIL.n101 VTAIL.n100 585
R199 VTAIL.n88 VTAIL.n87 585
R200 VTAIL.n95 VTAIL.n94 585
R201 VTAIL.n93 VTAIL.n92 585
R202 VTAIL.n73 VTAIL.n72 585
R203 VTAIL.n71 VTAIL.n70 585
R204 VTAIL.n46 VTAIL.n45 585
R205 VTAIL.n65 VTAIL.n64 585
R206 VTAIL.n63 VTAIL.n62 585
R207 VTAIL.n50 VTAIL.n49 585
R208 VTAIL.n57 VTAIL.n56 585
R209 VTAIL.n55 VTAIL.n54 585
R210 VTAIL.n127 VTAIL.t10 327.514
R211 VTAIL.n13 VTAIL.t2 327.514
R212 VTAIL.n91 VTAIL.t5 327.514
R213 VTAIL.n53 VTAIL.t9 327.514
R214 VTAIL.n130 VTAIL.n129 171.744
R215 VTAIL.n130 VTAIL.n123 171.744
R216 VTAIL.n137 VTAIL.n123 171.744
R217 VTAIL.n138 VTAIL.n137 171.744
R218 VTAIL.n138 VTAIL.n119 171.744
R219 VTAIL.n145 VTAIL.n119 171.744
R220 VTAIL.n146 VTAIL.n145 171.744
R221 VTAIL.n16 VTAIL.n15 171.744
R222 VTAIL.n16 VTAIL.n9 171.744
R223 VTAIL.n23 VTAIL.n9 171.744
R224 VTAIL.n24 VTAIL.n23 171.744
R225 VTAIL.n24 VTAIL.n5 171.744
R226 VTAIL.n31 VTAIL.n5 171.744
R227 VTAIL.n32 VTAIL.n31 171.744
R228 VTAIL.n110 VTAIL.n109 171.744
R229 VTAIL.n109 VTAIL.n83 171.744
R230 VTAIL.n102 VTAIL.n83 171.744
R231 VTAIL.n102 VTAIL.n101 171.744
R232 VTAIL.n101 VTAIL.n87 171.744
R233 VTAIL.n94 VTAIL.n87 171.744
R234 VTAIL.n94 VTAIL.n93 171.744
R235 VTAIL.n72 VTAIL.n71 171.744
R236 VTAIL.n71 VTAIL.n45 171.744
R237 VTAIL.n64 VTAIL.n45 171.744
R238 VTAIL.n64 VTAIL.n63 171.744
R239 VTAIL.n63 VTAIL.n49 171.744
R240 VTAIL.n56 VTAIL.n49 171.744
R241 VTAIL.n56 VTAIL.n55 171.744
R242 VTAIL.n129 VTAIL.t10 85.8723
R243 VTAIL.n15 VTAIL.t2 85.8723
R244 VTAIL.n93 VTAIL.t5 85.8723
R245 VTAIL.n55 VTAIL.t9 85.8723
R246 VTAIL.n79 VTAIL.n78 69.5868
R247 VTAIL.n41 VTAIL.n40 69.5868
R248 VTAIL.n1 VTAIL.n0 69.5867
R249 VTAIL.n39 VTAIL.n38 69.5867
R250 VTAIL.n151 VTAIL.n150 30.052
R251 VTAIL.n37 VTAIL.n36 30.052
R252 VTAIL.n115 VTAIL.n114 30.052
R253 VTAIL.n77 VTAIL.n76 30.052
R254 VTAIL.n41 VTAIL.n39 24.4789
R255 VTAIL.n151 VTAIL.n115 21.2721
R256 VTAIL.n128 VTAIL.n127 16.3884
R257 VTAIL.n14 VTAIL.n13 16.3884
R258 VTAIL.n92 VTAIL.n91 16.3884
R259 VTAIL.n54 VTAIL.n53 16.3884
R260 VTAIL.n131 VTAIL.n126 12.8005
R261 VTAIL.n17 VTAIL.n12 12.8005
R262 VTAIL.n95 VTAIL.n90 12.8005
R263 VTAIL.n57 VTAIL.n52 12.8005
R264 VTAIL.n132 VTAIL.n124 12.0247
R265 VTAIL.n18 VTAIL.n10 12.0247
R266 VTAIL.n96 VTAIL.n88 12.0247
R267 VTAIL.n58 VTAIL.n50 12.0247
R268 VTAIL.n136 VTAIL.n135 11.249
R269 VTAIL.n22 VTAIL.n21 11.249
R270 VTAIL.n100 VTAIL.n99 11.249
R271 VTAIL.n62 VTAIL.n61 11.249
R272 VTAIL.n139 VTAIL.n122 10.4732
R273 VTAIL.n25 VTAIL.n8 10.4732
R274 VTAIL.n103 VTAIL.n86 10.4732
R275 VTAIL.n65 VTAIL.n48 10.4732
R276 VTAIL.n140 VTAIL.n120 9.69747
R277 VTAIL.n26 VTAIL.n6 9.69747
R278 VTAIL.n104 VTAIL.n84 9.69747
R279 VTAIL.n66 VTAIL.n46 9.69747
R280 VTAIL.n150 VTAIL.n149 9.45567
R281 VTAIL.n36 VTAIL.n35 9.45567
R282 VTAIL.n114 VTAIL.n113 9.45567
R283 VTAIL.n76 VTAIL.n75 9.45567
R284 VTAIL.n118 VTAIL.n117 9.3005
R285 VTAIL.n143 VTAIL.n142 9.3005
R286 VTAIL.n141 VTAIL.n140 9.3005
R287 VTAIL.n122 VTAIL.n121 9.3005
R288 VTAIL.n135 VTAIL.n134 9.3005
R289 VTAIL.n133 VTAIL.n132 9.3005
R290 VTAIL.n126 VTAIL.n125 9.3005
R291 VTAIL.n149 VTAIL.n148 9.3005
R292 VTAIL.n4 VTAIL.n3 9.3005
R293 VTAIL.n29 VTAIL.n28 9.3005
R294 VTAIL.n27 VTAIL.n26 9.3005
R295 VTAIL.n8 VTAIL.n7 9.3005
R296 VTAIL.n21 VTAIL.n20 9.3005
R297 VTAIL.n19 VTAIL.n18 9.3005
R298 VTAIL.n12 VTAIL.n11 9.3005
R299 VTAIL.n35 VTAIL.n34 9.3005
R300 VTAIL.n113 VTAIL.n112 9.3005
R301 VTAIL.n82 VTAIL.n81 9.3005
R302 VTAIL.n107 VTAIL.n106 9.3005
R303 VTAIL.n105 VTAIL.n104 9.3005
R304 VTAIL.n86 VTAIL.n85 9.3005
R305 VTAIL.n99 VTAIL.n98 9.3005
R306 VTAIL.n97 VTAIL.n96 9.3005
R307 VTAIL.n90 VTAIL.n89 9.3005
R308 VTAIL.n75 VTAIL.n74 9.3005
R309 VTAIL.n44 VTAIL.n43 9.3005
R310 VTAIL.n69 VTAIL.n68 9.3005
R311 VTAIL.n67 VTAIL.n66 9.3005
R312 VTAIL.n48 VTAIL.n47 9.3005
R313 VTAIL.n61 VTAIL.n60 9.3005
R314 VTAIL.n59 VTAIL.n58 9.3005
R315 VTAIL.n52 VTAIL.n51 9.3005
R316 VTAIL.n144 VTAIL.n143 8.92171
R317 VTAIL.n30 VTAIL.n29 8.92171
R318 VTAIL.n108 VTAIL.n107 8.92171
R319 VTAIL.n70 VTAIL.n69 8.92171
R320 VTAIL.n147 VTAIL.n118 8.14595
R321 VTAIL.n33 VTAIL.n4 8.14595
R322 VTAIL.n111 VTAIL.n82 8.14595
R323 VTAIL.n73 VTAIL.n44 8.14595
R324 VTAIL.n148 VTAIL.n116 7.3702
R325 VTAIL.n34 VTAIL.n2 7.3702
R326 VTAIL.n112 VTAIL.n80 7.3702
R327 VTAIL.n74 VTAIL.n42 7.3702
R328 VTAIL.n150 VTAIL.n116 6.59444
R329 VTAIL.n36 VTAIL.n2 6.59444
R330 VTAIL.n114 VTAIL.n80 6.59444
R331 VTAIL.n76 VTAIL.n42 6.59444
R332 VTAIL.n148 VTAIL.n147 5.81868
R333 VTAIL.n34 VTAIL.n33 5.81868
R334 VTAIL.n112 VTAIL.n111 5.81868
R335 VTAIL.n74 VTAIL.n73 5.81868
R336 VTAIL.n144 VTAIL.n118 5.04292
R337 VTAIL.n30 VTAIL.n4 5.04292
R338 VTAIL.n108 VTAIL.n82 5.04292
R339 VTAIL.n70 VTAIL.n44 5.04292
R340 VTAIL.n0 VTAIL.t7 4.91805
R341 VTAIL.n0 VTAIL.t8 4.91805
R342 VTAIL.n38 VTAIL.t3 4.91805
R343 VTAIL.n38 VTAIL.t4 4.91805
R344 VTAIL.n78 VTAIL.t0 4.91805
R345 VTAIL.n78 VTAIL.t1 4.91805
R346 VTAIL.n40 VTAIL.t6 4.91805
R347 VTAIL.n40 VTAIL.t11 4.91805
R348 VTAIL.n143 VTAIL.n120 4.26717
R349 VTAIL.n29 VTAIL.n6 4.26717
R350 VTAIL.n107 VTAIL.n84 4.26717
R351 VTAIL.n69 VTAIL.n46 4.26717
R352 VTAIL.n127 VTAIL.n125 3.71088
R353 VTAIL.n13 VTAIL.n11 3.71088
R354 VTAIL.n91 VTAIL.n89 3.71088
R355 VTAIL.n53 VTAIL.n51 3.71088
R356 VTAIL.n140 VTAIL.n139 3.49141
R357 VTAIL.n26 VTAIL.n25 3.49141
R358 VTAIL.n104 VTAIL.n103 3.49141
R359 VTAIL.n66 VTAIL.n65 3.49141
R360 VTAIL.n77 VTAIL.n41 3.2074
R361 VTAIL.n115 VTAIL.n79 3.2074
R362 VTAIL.n39 VTAIL.n37 3.2074
R363 VTAIL.n136 VTAIL.n122 2.71565
R364 VTAIL.n22 VTAIL.n8 2.71565
R365 VTAIL.n100 VTAIL.n86 2.71565
R366 VTAIL.n62 VTAIL.n48 2.71565
R367 VTAIL VTAIL.n151 2.34748
R368 VTAIL.n79 VTAIL.n77 2.07378
R369 VTAIL.n37 VTAIL.n1 2.07378
R370 VTAIL.n135 VTAIL.n124 1.93989
R371 VTAIL.n21 VTAIL.n10 1.93989
R372 VTAIL.n99 VTAIL.n88 1.93989
R373 VTAIL.n61 VTAIL.n50 1.93989
R374 VTAIL.n132 VTAIL.n131 1.16414
R375 VTAIL.n18 VTAIL.n17 1.16414
R376 VTAIL.n96 VTAIL.n95 1.16414
R377 VTAIL.n58 VTAIL.n57 1.16414
R378 VTAIL VTAIL.n1 0.860414
R379 VTAIL.n128 VTAIL.n126 0.388379
R380 VTAIL.n14 VTAIL.n12 0.388379
R381 VTAIL.n92 VTAIL.n90 0.388379
R382 VTAIL.n54 VTAIL.n52 0.388379
R383 VTAIL.n133 VTAIL.n125 0.155672
R384 VTAIL.n134 VTAIL.n133 0.155672
R385 VTAIL.n134 VTAIL.n121 0.155672
R386 VTAIL.n141 VTAIL.n121 0.155672
R387 VTAIL.n142 VTAIL.n141 0.155672
R388 VTAIL.n142 VTAIL.n117 0.155672
R389 VTAIL.n149 VTAIL.n117 0.155672
R390 VTAIL.n19 VTAIL.n11 0.155672
R391 VTAIL.n20 VTAIL.n19 0.155672
R392 VTAIL.n20 VTAIL.n7 0.155672
R393 VTAIL.n27 VTAIL.n7 0.155672
R394 VTAIL.n28 VTAIL.n27 0.155672
R395 VTAIL.n28 VTAIL.n3 0.155672
R396 VTAIL.n35 VTAIL.n3 0.155672
R397 VTAIL.n113 VTAIL.n81 0.155672
R398 VTAIL.n106 VTAIL.n81 0.155672
R399 VTAIL.n106 VTAIL.n105 0.155672
R400 VTAIL.n105 VTAIL.n85 0.155672
R401 VTAIL.n98 VTAIL.n85 0.155672
R402 VTAIL.n98 VTAIL.n97 0.155672
R403 VTAIL.n97 VTAIL.n89 0.155672
R404 VTAIL.n75 VTAIL.n43 0.155672
R405 VTAIL.n68 VTAIL.n43 0.155672
R406 VTAIL.n68 VTAIL.n67 0.155672
R407 VTAIL.n67 VTAIL.n47 0.155672
R408 VTAIL.n60 VTAIL.n47 0.155672
R409 VTAIL.n60 VTAIL.n59 0.155672
R410 VTAIL.n59 VTAIL.n51 0.155672
R411 VP.n16 VP.n15 161.3
R412 VP.n17 VP.n12 161.3
R413 VP.n19 VP.n18 161.3
R414 VP.n20 VP.n11 161.3
R415 VP.n22 VP.n21 161.3
R416 VP.n23 VP.n10 161.3
R417 VP.n25 VP.n24 161.3
R418 VP.n50 VP.n49 161.3
R419 VP.n48 VP.n1 161.3
R420 VP.n47 VP.n46 161.3
R421 VP.n45 VP.n2 161.3
R422 VP.n44 VP.n43 161.3
R423 VP.n42 VP.n3 161.3
R424 VP.n41 VP.n40 161.3
R425 VP.n39 VP.n4 161.3
R426 VP.n38 VP.n37 161.3
R427 VP.n36 VP.n5 161.3
R428 VP.n35 VP.n34 161.3
R429 VP.n33 VP.n6 161.3
R430 VP.n32 VP.n31 161.3
R431 VP.n30 VP.n7 161.3
R432 VP.n29 VP.n28 161.3
R433 VP.n14 VP.t2 80.5477
R434 VP.n27 VP.n8 79.3019
R435 VP.n51 VP.n0 79.3019
R436 VP.n26 VP.n9 79.3019
R437 VP.n35 VP.n6 54.0911
R438 VP.n43 VP.n2 54.0911
R439 VP.n18 VP.n11 54.0911
R440 VP.n14 VP.n13 50.1285
R441 VP.n27 VP.n26 47.7645
R442 VP.n4 VP.t0 46.9919
R443 VP.n8 VP.t1 46.9919
R444 VP.n0 VP.t4 46.9919
R445 VP.n13 VP.t5 46.9919
R446 VP.n9 VP.t3 46.9919
R447 VP.n31 VP.n6 26.8957
R448 VP.n47 VP.n2 26.8957
R449 VP.n22 VP.n11 26.8957
R450 VP.n30 VP.n29 24.4675
R451 VP.n31 VP.n30 24.4675
R452 VP.n36 VP.n35 24.4675
R453 VP.n37 VP.n36 24.4675
R454 VP.n37 VP.n4 24.4675
R455 VP.n41 VP.n4 24.4675
R456 VP.n42 VP.n41 24.4675
R457 VP.n43 VP.n42 24.4675
R458 VP.n48 VP.n47 24.4675
R459 VP.n49 VP.n48 24.4675
R460 VP.n23 VP.n22 24.4675
R461 VP.n24 VP.n23 24.4675
R462 VP.n16 VP.n13 24.4675
R463 VP.n17 VP.n16 24.4675
R464 VP.n18 VP.n17 24.4675
R465 VP.n29 VP.n8 10.766
R466 VP.n49 VP.n0 10.766
R467 VP.n24 VP.n9 10.766
R468 VP.n15 VP.n14 3.1271
R469 VP.n26 VP.n25 0.354971
R470 VP.n28 VP.n27 0.354971
R471 VP.n51 VP.n50 0.354971
R472 VP VP.n51 0.26696
R473 VP.n15 VP.n12 0.189894
R474 VP.n19 VP.n12 0.189894
R475 VP.n20 VP.n19 0.189894
R476 VP.n21 VP.n20 0.189894
R477 VP.n21 VP.n10 0.189894
R478 VP.n25 VP.n10 0.189894
R479 VP.n28 VP.n7 0.189894
R480 VP.n32 VP.n7 0.189894
R481 VP.n33 VP.n32 0.189894
R482 VP.n34 VP.n33 0.189894
R483 VP.n34 VP.n5 0.189894
R484 VP.n38 VP.n5 0.189894
R485 VP.n39 VP.n38 0.189894
R486 VP.n40 VP.n39 0.189894
R487 VP.n40 VP.n3 0.189894
R488 VP.n44 VP.n3 0.189894
R489 VP.n45 VP.n44 0.189894
R490 VP.n46 VP.n45 0.189894
R491 VP.n46 VP.n1 0.189894
R492 VP.n50 VP.n1 0.189894
R493 VDD1.n30 VDD1.n0 756.745
R494 VDD1.n65 VDD1.n35 756.745
R495 VDD1.n31 VDD1.n30 585
R496 VDD1.n29 VDD1.n28 585
R497 VDD1.n4 VDD1.n3 585
R498 VDD1.n23 VDD1.n22 585
R499 VDD1.n21 VDD1.n20 585
R500 VDD1.n8 VDD1.n7 585
R501 VDD1.n15 VDD1.n14 585
R502 VDD1.n13 VDD1.n12 585
R503 VDD1.n48 VDD1.n47 585
R504 VDD1.n50 VDD1.n49 585
R505 VDD1.n43 VDD1.n42 585
R506 VDD1.n56 VDD1.n55 585
R507 VDD1.n58 VDD1.n57 585
R508 VDD1.n39 VDD1.n38 585
R509 VDD1.n64 VDD1.n63 585
R510 VDD1.n66 VDD1.n65 585
R511 VDD1.n11 VDD1.t3 327.514
R512 VDD1.n46 VDD1.t4 327.514
R513 VDD1.n30 VDD1.n29 171.744
R514 VDD1.n29 VDD1.n3 171.744
R515 VDD1.n22 VDD1.n3 171.744
R516 VDD1.n22 VDD1.n21 171.744
R517 VDD1.n21 VDD1.n7 171.744
R518 VDD1.n14 VDD1.n7 171.744
R519 VDD1.n14 VDD1.n13 171.744
R520 VDD1.n49 VDD1.n48 171.744
R521 VDD1.n49 VDD1.n42 171.744
R522 VDD1.n56 VDD1.n42 171.744
R523 VDD1.n57 VDD1.n56 171.744
R524 VDD1.n57 VDD1.n38 171.744
R525 VDD1.n64 VDD1.n38 171.744
R526 VDD1.n65 VDD1.n64 171.744
R527 VDD1.n71 VDD1.n70 87.0118
R528 VDD1.n73 VDD1.n72 86.2655
R529 VDD1.n13 VDD1.t3 85.8723
R530 VDD1.n48 VDD1.t4 85.8723
R531 VDD1 VDD1.n34 49.1942
R532 VDD1.n71 VDD1.n69 49.0806
R533 VDD1.n73 VDD1.n71 42.0224
R534 VDD1.n47 VDD1.n46 16.3884
R535 VDD1.n12 VDD1.n11 16.3884
R536 VDD1.n15 VDD1.n10 12.8005
R537 VDD1.n50 VDD1.n45 12.8005
R538 VDD1.n16 VDD1.n8 12.0247
R539 VDD1.n51 VDD1.n43 12.0247
R540 VDD1.n20 VDD1.n19 11.249
R541 VDD1.n55 VDD1.n54 11.249
R542 VDD1.n23 VDD1.n6 10.4732
R543 VDD1.n58 VDD1.n41 10.4732
R544 VDD1.n24 VDD1.n4 9.69747
R545 VDD1.n59 VDD1.n39 9.69747
R546 VDD1.n34 VDD1.n33 9.45567
R547 VDD1.n69 VDD1.n68 9.45567
R548 VDD1.n33 VDD1.n32 9.3005
R549 VDD1.n2 VDD1.n1 9.3005
R550 VDD1.n27 VDD1.n26 9.3005
R551 VDD1.n25 VDD1.n24 9.3005
R552 VDD1.n6 VDD1.n5 9.3005
R553 VDD1.n19 VDD1.n18 9.3005
R554 VDD1.n17 VDD1.n16 9.3005
R555 VDD1.n10 VDD1.n9 9.3005
R556 VDD1.n37 VDD1.n36 9.3005
R557 VDD1.n62 VDD1.n61 9.3005
R558 VDD1.n60 VDD1.n59 9.3005
R559 VDD1.n41 VDD1.n40 9.3005
R560 VDD1.n54 VDD1.n53 9.3005
R561 VDD1.n52 VDD1.n51 9.3005
R562 VDD1.n45 VDD1.n44 9.3005
R563 VDD1.n68 VDD1.n67 9.3005
R564 VDD1.n28 VDD1.n27 8.92171
R565 VDD1.n63 VDD1.n62 8.92171
R566 VDD1.n31 VDD1.n2 8.14595
R567 VDD1.n66 VDD1.n37 8.14595
R568 VDD1.n32 VDD1.n0 7.3702
R569 VDD1.n67 VDD1.n35 7.3702
R570 VDD1.n34 VDD1.n0 6.59444
R571 VDD1.n69 VDD1.n35 6.59444
R572 VDD1.n32 VDD1.n31 5.81868
R573 VDD1.n67 VDD1.n66 5.81868
R574 VDD1.n28 VDD1.n2 5.04292
R575 VDD1.n63 VDD1.n37 5.04292
R576 VDD1.n72 VDD1.t0 4.91805
R577 VDD1.n72 VDD1.t2 4.91805
R578 VDD1.n70 VDD1.t5 4.91805
R579 VDD1.n70 VDD1.t1 4.91805
R580 VDD1.n27 VDD1.n4 4.26717
R581 VDD1.n62 VDD1.n39 4.26717
R582 VDD1.n11 VDD1.n9 3.71088
R583 VDD1.n46 VDD1.n44 3.71088
R584 VDD1.n24 VDD1.n23 3.49141
R585 VDD1.n59 VDD1.n58 3.49141
R586 VDD1.n20 VDD1.n6 2.71565
R587 VDD1.n55 VDD1.n41 2.71565
R588 VDD1.n19 VDD1.n8 1.93989
R589 VDD1.n54 VDD1.n43 1.93989
R590 VDD1.n16 VDD1.n15 1.16414
R591 VDD1.n51 VDD1.n50 1.16414
R592 VDD1 VDD1.n73 0.744035
R593 VDD1.n12 VDD1.n10 0.388379
R594 VDD1.n47 VDD1.n45 0.388379
R595 VDD1.n33 VDD1.n1 0.155672
R596 VDD1.n26 VDD1.n1 0.155672
R597 VDD1.n26 VDD1.n25 0.155672
R598 VDD1.n25 VDD1.n5 0.155672
R599 VDD1.n18 VDD1.n5 0.155672
R600 VDD1.n18 VDD1.n17 0.155672
R601 VDD1.n17 VDD1.n9 0.155672
R602 VDD1.n52 VDD1.n44 0.155672
R603 VDD1.n53 VDD1.n52 0.155672
R604 VDD1.n53 VDD1.n40 0.155672
R605 VDD1.n60 VDD1.n40 0.155672
R606 VDD1.n61 VDD1.n60 0.155672
R607 VDD1.n61 VDD1.n36 0.155672
R608 VDD1.n68 VDD1.n36 0.155672
R609 B.n503 B.n62 585
R610 B.n505 B.n504 585
R611 B.n506 B.n61 585
R612 B.n508 B.n507 585
R613 B.n509 B.n60 585
R614 B.n511 B.n510 585
R615 B.n512 B.n59 585
R616 B.n514 B.n513 585
R617 B.n515 B.n58 585
R618 B.n517 B.n516 585
R619 B.n518 B.n57 585
R620 B.n520 B.n519 585
R621 B.n521 B.n56 585
R622 B.n523 B.n522 585
R623 B.n524 B.n55 585
R624 B.n526 B.n525 585
R625 B.n527 B.n54 585
R626 B.n529 B.n528 585
R627 B.n530 B.n53 585
R628 B.n532 B.n531 585
R629 B.n533 B.n52 585
R630 B.n535 B.n534 585
R631 B.n536 B.n51 585
R632 B.n538 B.n537 585
R633 B.n539 B.n50 585
R634 B.n541 B.n540 585
R635 B.n543 B.n47 585
R636 B.n545 B.n544 585
R637 B.n546 B.n46 585
R638 B.n548 B.n547 585
R639 B.n549 B.n45 585
R640 B.n551 B.n550 585
R641 B.n552 B.n44 585
R642 B.n554 B.n553 585
R643 B.n555 B.n41 585
R644 B.n558 B.n557 585
R645 B.n559 B.n40 585
R646 B.n561 B.n560 585
R647 B.n562 B.n39 585
R648 B.n564 B.n563 585
R649 B.n565 B.n38 585
R650 B.n567 B.n566 585
R651 B.n568 B.n37 585
R652 B.n570 B.n569 585
R653 B.n571 B.n36 585
R654 B.n573 B.n572 585
R655 B.n574 B.n35 585
R656 B.n576 B.n575 585
R657 B.n577 B.n34 585
R658 B.n579 B.n578 585
R659 B.n580 B.n33 585
R660 B.n582 B.n581 585
R661 B.n583 B.n32 585
R662 B.n585 B.n584 585
R663 B.n586 B.n31 585
R664 B.n588 B.n587 585
R665 B.n589 B.n30 585
R666 B.n591 B.n590 585
R667 B.n592 B.n29 585
R668 B.n594 B.n593 585
R669 B.n595 B.n28 585
R670 B.n502 B.n501 585
R671 B.n500 B.n63 585
R672 B.n499 B.n498 585
R673 B.n497 B.n64 585
R674 B.n496 B.n495 585
R675 B.n494 B.n65 585
R676 B.n493 B.n492 585
R677 B.n491 B.n66 585
R678 B.n490 B.n489 585
R679 B.n488 B.n67 585
R680 B.n487 B.n486 585
R681 B.n485 B.n68 585
R682 B.n484 B.n483 585
R683 B.n482 B.n69 585
R684 B.n481 B.n480 585
R685 B.n479 B.n70 585
R686 B.n478 B.n477 585
R687 B.n476 B.n71 585
R688 B.n475 B.n474 585
R689 B.n473 B.n72 585
R690 B.n472 B.n471 585
R691 B.n470 B.n73 585
R692 B.n469 B.n468 585
R693 B.n467 B.n74 585
R694 B.n466 B.n465 585
R695 B.n464 B.n75 585
R696 B.n463 B.n462 585
R697 B.n461 B.n76 585
R698 B.n460 B.n459 585
R699 B.n458 B.n77 585
R700 B.n457 B.n456 585
R701 B.n455 B.n78 585
R702 B.n454 B.n453 585
R703 B.n452 B.n79 585
R704 B.n451 B.n450 585
R705 B.n449 B.n80 585
R706 B.n448 B.n447 585
R707 B.n446 B.n81 585
R708 B.n445 B.n444 585
R709 B.n443 B.n82 585
R710 B.n442 B.n441 585
R711 B.n440 B.n83 585
R712 B.n439 B.n438 585
R713 B.n437 B.n84 585
R714 B.n436 B.n435 585
R715 B.n434 B.n85 585
R716 B.n433 B.n432 585
R717 B.n431 B.n86 585
R718 B.n430 B.n429 585
R719 B.n428 B.n87 585
R720 B.n427 B.n426 585
R721 B.n425 B.n88 585
R722 B.n424 B.n423 585
R723 B.n422 B.n89 585
R724 B.n421 B.n420 585
R725 B.n419 B.n90 585
R726 B.n418 B.n417 585
R727 B.n416 B.n91 585
R728 B.n415 B.n414 585
R729 B.n413 B.n92 585
R730 B.n412 B.n411 585
R731 B.n410 B.n93 585
R732 B.n409 B.n408 585
R733 B.n407 B.n94 585
R734 B.n406 B.n405 585
R735 B.n404 B.n95 585
R736 B.n403 B.n402 585
R737 B.n401 B.n96 585
R738 B.n400 B.n399 585
R739 B.n398 B.n97 585
R740 B.n397 B.n396 585
R741 B.n395 B.n98 585
R742 B.n394 B.n393 585
R743 B.n392 B.n99 585
R744 B.n391 B.n390 585
R745 B.n389 B.n100 585
R746 B.n388 B.n387 585
R747 B.n386 B.n101 585
R748 B.n385 B.n384 585
R749 B.n383 B.n102 585
R750 B.n382 B.n381 585
R751 B.n380 B.n103 585
R752 B.n379 B.n378 585
R753 B.n377 B.n104 585
R754 B.n376 B.n375 585
R755 B.n374 B.n105 585
R756 B.n373 B.n372 585
R757 B.n371 B.n106 585
R758 B.n370 B.n369 585
R759 B.n368 B.n107 585
R760 B.n367 B.n366 585
R761 B.n365 B.n108 585
R762 B.n364 B.n363 585
R763 B.n362 B.n109 585
R764 B.n361 B.n360 585
R765 B.n359 B.n110 585
R766 B.n358 B.n357 585
R767 B.n356 B.n111 585
R768 B.n355 B.n354 585
R769 B.n353 B.n112 585
R770 B.n352 B.n351 585
R771 B.n350 B.n113 585
R772 B.n349 B.n348 585
R773 B.n347 B.n114 585
R774 B.n346 B.n345 585
R775 B.n253 B.n252 585
R776 B.n254 B.n149 585
R777 B.n256 B.n255 585
R778 B.n257 B.n148 585
R779 B.n259 B.n258 585
R780 B.n260 B.n147 585
R781 B.n262 B.n261 585
R782 B.n263 B.n146 585
R783 B.n265 B.n264 585
R784 B.n266 B.n145 585
R785 B.n268 B.n267 585
R786 B.n269 B.n144 585
R787 B.n271 B.n270 585
R788 B.n272 B.n143 585
R789 B.n274 B.n273 585
R790 B.n275 B.n142 585
R791 B.n277 B.n276 585
R792 B.n278 B.n141 585
R793 B.n280 B.n279 585
R794 B.n281 B.n140 585
R795 B.n283 B.n282 585
R796 B.n284 B.n139 585
R797 B.n286 B.n285 585
R798 B.n287 B.n138 585
R799 B.n289 B.n288 585
R800 B.n290 B.n135 585
R801 B.n293 B.n292 585
R802 B.n294 B.n134 585
R803 B.n296 B.n295 585
R804 B.n297 B.n133 585
R805 B.n299 B.n298 585
R806 B.n300 B.n132 585
R807 B.n302 B.n301 585
R808 B.n303 B.n131 585
R809 B.n305 B.n304 585
R810 B.n307 B.n306 585
R811 B.n308 B.n127 585
R812 B.n310 B.n309 585
R813 B.n311 B.n126 585
R814 B.n313 B.n312 585
R815 B.n314 B.n125 585
R816 B.n316 B.n315 585
R817 B.n317 B.n124 585
R818 B.n319 B.n318 585
R819 B.n320 B.n123 585
R820 B.n322 B.n321 585
R821 B.n323 B.n122 585
R822 B.n325 B.n324 585
R823 B.n326 B.n121 585
R824 B.n328 B.n327 585
R825 B.n329 B.n120 585
R826 B.n331 B.n330 585
R827 B.n332 B.n119 585
R828 B.n334 B.n333 585
R829 B.n335 B.n118 585
R830 B.n337 B.n336 585
R831 B.n338 B.n117 585
R832 B.n340 B.n339 585
R833 B.n341 B.n116 585
R834 B.n343 B.n342 585
R835 B.n344 B.n115 585
R836 B.n251 B.n150 585
R837 B.n250 B.n249 585
R838 B.n248 B.n151 585
R839 B.n247 B.n246 585
R840 B.n245 B.n152 585
R841 B.n244 B.n243 585
R842 B.n242 B.n153 585
R843 B.n241 B.n240 585
R844 B.n239 B.n154 585
R845 B.n238 B.n237 585
R846 B.n236 B.n155 585
R847 B.n235 B.n234 585
R848 B.n233 B.n156 585
R849 B.n232 B.n231 585
R850 B.n230 B.n157 585
R851 B.n229 B.n228 585
R852 B.n227 B.n158 585
R853 B.n226 B.n225 585
R854 B.n224 B.n159 585
R855 B.n223 B.n222 585
R856 B.n221 B.n160 585
R857 B.n220 B.n219 585
R858 B.n218 B.n161 585
R859 B.n217 B.n216 585
R860 B.n215 B.n162 585
R861 B.n214 B.n213 585
R862 B.n212 B.n163 585
R863 B.n211 B.n210 585
R864 B.n209 B.n164 585
R865 B.n208 B.n207 585
R866 B.n206 B.n165 585
R867 B.n205 B.n204 585
R868 B.n203 B.n166 585
R869 B.n202 B.n201 585
R870 B.n200 B.n167 585
R871 B.n199 B.n198 585
R872 B.n197 B.n168 585
R873 B.n196 B.n195 585
R874 B.n194 B.n169 585
R875 B.n193 B.n192 585
R876 B.n191 B.n170 585
R877 B.n190 B.n189 585
R878 B.n188 B.n171 585
R879 B.n187 B.n186 585
R880 B.n185 B.n172 585
R881 B.n184 B.n183 585
R882 B.n182 B.n173 585
R883 B.n181 B.n180 585
R884 B.n179 B.n174 585
R885 B.n178 B.n177 585
R886 B.n176 B.n175 585
R887 B.n2 B.n0 585
R888 B.n673 B.n1 585
R889 B.n672 B.n671 585
R890 B.n670 B.n3 585
R891 B.n669 B.n668 585
R892 B.n667 B.n4 585
R893 B.n666 B.n665 585
R894 B.n664 B.n5 585
R895 B.n663 B.n662 585
R896 B.n661 B.n6 585
R897 B.n660 B.n659 585
R898 B.n658 B.n7 585
R899 B.n657 B.n656 585
R900 B.n655 B.n8 585
R901 B.n654 B.n653 585
R902 B.n652 B.n9 585
R903 B.n651 B.n650 585
R904 B.n649 B.n10 585
R905 B.n648 B.n647 585
R906 B.n646 B.n11 585
R907 B.n645 B.n644 585
R908 B.n643 B.n12 585
R909 B.n642 B.n641 585
R910 B.n640 B.n13 585
R911 B.n639 B.n638 585
R912 B.n637 B.n14 585
R913 B.n636 B.n635 585
R914 B.n634 B.n15 585
R915 B.n633 B.n632 585
R916 B.n631 B.n16 585
R917 B.n630 B.n629 585
R918 B.n628 B.n17 585
R919 B.n627 B.n626 585
R920 B.n625 B.n18 585
R921 B.n624 B.n623 585
R922 B.n622 B.n19 585
R923 B.n621 B.n620 585
R924 B.n619 B.n20 585
R925 B.n618 B.n617 585
R926 B.n616 B.n21 585
R927 B.n615 B.n614 585
R928 B.n613 B.n22 585
R929 B.n612 B.n611 585
R930 B.n610 B.n23 585
R931 B.n609 B.n608 585
R932 B.n607 B.n24 585
R933 B.n606 B.n605 585
R934 B.n604 B.n25 585
R935 B.n603 B.n602 585
R936 B.n601 B.n26 585
R937 B.n600 B.n599 585
R938 B.n598 B.n27 585
R939 B.n597 B.n596 585
R940 B.n675 B.n674 585
R941 B.n252 B.n251 487.695
R942 B.n596 B.n595 487.695
R943 B.n346 B.n115 487.695
R944 B.n503 B.n502 487.695
R945 B.n128 B.t11 350.974
R946 B.n48 B.t7 350.974
R947 B.n136 B.t2 350.974
R948 B.n42 B.t4 350.974
R949 B.n129 B.t10 278.829
R950 B.n49 B.t8 278.829
R951 B.n137 B.t1 278.829
R952 B.n43 B.t5 278.829
R953 B.n128 B.t9 255.983
R954 B.n136 B.t0 255.983
R955 B.n42 B.t3 255.983
R956 B.n48 B.t6 255.983
R957 B.n251 B.n250 163.367
R958 B.n250 B.n151 163.367
R959 B.n246 B.n151 163.367
R960 B.n246 B.n245 163.367
R961 B.n245 B.n244 163.367
R962 B.n244 B.n153 163.367
R963 B.n240 B.n153 163.367
R964 B.n240 B.n239 163.367
R965 B.n239 B.n238 163.367
R966 B.n238 B.n155 163.367
R967 B.n234 B.n155 163.367
R968 B.n234 B.n233 163.367
R969 B.n233 B.n232 163.367
R970 B.n232 B.n157 163.367
R971 B.n228 B.n157 163.367
R972 B.n228 B.n227 163.367
R973 B.n227 B.n226 163.367
R974 B.n226 B.n159 163.367
R975 B.n222 B.n159 163.367
R976 B.n222 B.n221 163.367
R977 B.n221 B.n220 163.367
R978 B.n220 B.n161 163.367
R979 B.n216 B.n161 163.367
R980 B.n216 B.n215 163.367
R981 B.n215 B.n214 163.367
R982 B.n214 B.n163 163.367
R983 B.n210 B.n163 163.367
R984 B.n210 B.n209 163.367
R985 B.n209 B.n208 163.367
R986 B.n208 B.n165 163.367
R987 B.n204 B.n165 163.367
R988 B.n204 B.n203 163.367
R989 B.n203 B.n202 163.367
R990 B.n202 B.n167 163.367
R991 B.n198 B.n167 163.367
R992 B.n198 B.n197 163.367
R993 B.n197 B.n196 163.367
R994 B.n196 B.n169 163.367
R995 B.n192 B.n169 163.367
R996 B.n192 B.n191 163.367
R997 B.n191 B.n190 163.367
R998 B.n190 B.n171 163.367
R999 B.n186 B.n171 163.367
R1000 B.n186 B.n185 163.367
R1001 B.n185 B.n184 163.367
R1002 B.n184 B.n173 163.367
R1003 B.n180 B.n173 163.367
R1004 B.n180 B.n179 163.367
R1005 B.n179 B.n178 163.367
R1006 B.n178 B.n175 163.367
R1007 B.n175 B.n2 163.367
R1008 B.n674 B.n2 163.367
R1009 B.n674 B.n673 163.367
R1010 B.n673 B.n672 163.367
R1011 B.n672 B.n3 163.367
R1012 B.n668 B.n3 163.367
R1013 B.n668 B.n667 163.367
R1014 B.n667 B.n666 163.367
R1015 B.n666 B.n5 163.367
R1016 B.n662 B.n5 163.367
R1017 B.n662 B.n661 163.367
R1018 B.n661 B.n660 163.367
R1019 B.n660 B.n7 163.367
R1020 B.n656 B.n7 163.367
R1021 B.n656 B.n655 163.367
R1022 B.n655 B.n654 163.367
R1023 B.n654 B.n9 163.367
R1024 B.n650 B.n9 163.367
R1025 B.n650 B.n649 163.367
R1026 B.n649 B.n648 163.367
R1027 B.n648 B.n11 163.367
R1028 B.n644 B.n11 163.367
R1029 B.n644 B.n643 163.367
R1030 B.n643 B.n642 163.367
R1031 B.n642 B.n13 163.367
R1032 B.n638 B.n13 163.367
R1033 B.n638 B.n637 163.367
R1034 B.n637 B.n636 163.367
R1035 B.n636 B.n15 163.367
R1036 B.n632 B.n15 163.367
R1037 B.n632 B.n631 163.367
R1038 B.n631 B.n630 163.367
R1039 B.n630 B.n17 163.367
R1040 B.n626 B.n17 163.367
R1041 B.n626 B.n625 163.367
R1042 B.n625 B.n624 163.367
R1043 B.n624 B.n19 163.367
R1044 B.n620 B.n19 163.367
R1045 B.n620 B.n619 163.367
R1046 B.n619 B.n618 163.367
R1047 B.n618 B.n21 163.367
R1048 B.n614 B.n21 163.367
R1049 B.n614 B.n613 163.367
R1050 B.n613 B.n612 163.367
R1051 B.n612 B.n23 163.367
R1052 B.n608 B.n23 163.367
R1053 B.n608 B.n607 163.367
R1054 B.n607 B.n606 163.367
R1055 B.n606 B.n25 163.367
R1056 B.n602 B.n25 163.367
R1057 B.n602 B.n601 163.367
R1058 B.n601 B.n600 163.367
R1059 B.n600 B.n27 163.367
R1060 B.n596 B.n27 163.367
R1061 B.n252 B.n149 163.367
R1062 B.n256 B.n149 163.367
R1063 B.n257 B.n256 163.367
R1064 B.n258 B.n257 163.367
R1065 B.n258 B.n147 163.367
R1066 B.n262 B.n147 163.367
R1067 B.n263 B.n262 163.367
R1068 B.n264 B.n263 163.367
R1069 B.n264 B.n145 163.367
R1070 B.n268 B.n145 163.367
R1071 B.n269 B.n268 163.367
R1072 B.n270 B.n269 163.367
R1073 B.n270 B.n143 163.367
R1074 B.n274 B.n143 163.367
R1075 B.n275 B.n274 163.367
R1076 B.n276 B.n275 163.367
R1077 B.n276 B.n141 163.367
R1078 B.n280 B.n141 163.367
R1079 B.n281 B.n280 163.367
R1080 B.n282 B.n281 163.367
R1081 B.n282 B.n139 163.367
R1082 B.n286 B.n139 163.367
R1083 B.n287 B.n286 163.367
R1084 B.n288 B.n287 163.367
R1085 B.n288 B.n135 163.367
R1086 B.n293 B.n135 163.367
R1087 B.n294 B.n293 163.367
R1088 B.n295 B.n294 163.367
R1089 B.n295 B.n133 163.367
R1090 B.n299 B.n133 163.367
R1091 B.n300 B.n299 163.367
R1092 B.n301 B.n300 163.367
R1093 B.n301 B.n131 163.367
R1094 B.n305 B.n131 163.367
R1095 B.n306 B.n305 163.367
R1096 B.n306 B.n127 163.367
R1097 B.n310 B.n127 163.367
R1098 B.n311 B.n310 163.367
R1099 B.n312 B.n311 163.367
R1100 B.n312 B.n125 163.367
R1101 B.n316 B.n125 163.367
R1102 B.n317 B.n316 163.367
R1103 B.n318 B.n317 163.367
R1104 B.n318 B.n123 163.367
R1105 B.n322 B.n123 163.367
R1106 B.n323 B.n322 163.367
R1107 B.n324 B.n323 163.367
R1108 B.n324 B.n121 163.367
R1109 B.n328 B.n121 163.367
R1110 B.n329 B.n328 163.367
R1111 B.n330 B.n329 163.367
R1112 B.n330 B.n119 163.367
R1113 B.n334 B.n119 163.367
R1114 B.n335 B.n334 163.367
R1115 B.n336 B.n335 163.367
R1116 B.n336 B.n117 163.367
R1117 B.n340 B.n117 163.367
R1118 B.n341 B.n340 163.367
R1119 B.n342 B.n341 163.367
R1120 B.n342 B.n115 163.367
R1121 B.n347 B.n346 163.367
R1122 B.n348 B.n347 163.367
R1123 B.n348 B.n113 163.367
R1124 B.n352 B.n113 163.367
R1125 B.n353 B.n352 163.367
R1126 B.n354 B.n353 163.367
R1127 B.n354 B.n111 163.367
R1128 B.n358 B.n111 163.367
R1129 B.n359 B.n358 163.367
R1130 B.n360 B.n359 163.367
R1131 B.n360 B.n109 163.367
R1132 B.n364 B.n109 163.367
R1133 B.n365 B.n364 163.367
R1134 B.n366 B.n365 163.367
R1135 B.n366 B.n107 163.367
R1136 B.n370 B.n107 163.367
R1137 B.n371 B.n370 163.367
R1138 B.n372 B.n371 163.367
R1139 B.n372 B.n105 163.367
R1140 B.n376 B.n105 163.367
R1141 B.n377 B.n376 163.367
R1142 B.n378 B.n377 163.367
R1143 B.n378 B.n103 163.367
R1144 B.n382 B.n103 163.367
R1145 B.n383 B.n382 163.367
R1146 B.n384 B.n383 163.367
R1147 B.n384 B.n101 163.367
R1148 B.n388 B.n101 163.367
R1149 B.n389 B.n388 163.367
R1150 B.n390 B.n389 163.367
R1151 B.n390 B.n99 163.367
R1152 B.n394 B.n99 163.367
R1153 B.n395 B.n394 163.367
R1154 B.n396 B.n395 163.367
R1155 B.n396 B.n97 163.367
R1156 B.n400 B.n97 163.367
R1157 B.n401 B.n400 163.367
R1158 B.n402 B.n401 163.367
R1159 B.n402 B.n95 163.367
R1160 B.n406 B.n95 163.367
R1161 B.n407 B.n406 163.367
R1162 B.n408 B.n407 163.367
R1163 B.n408 B.n93 163.367
R1164 B.n412 B.n93 163.367
R1165 B.n413 B.n412 163.367
R1166 B.n414 B.n413 163.367
R1167 B.n414 B.n91 163.367
R1168 B.n418 B.n91 163.367
R1169 B.n419 B.n418 163.367
R1170 B.n420 B.n419 163.367
R1171 B.n420 B.n89 163.367
R1172 B.n424 B.n89 163.367
R1173 B.n425 B.n424 163.367
R1174 B.n426 B.n425 163.367
R1175 B.n426 B.n87 163.367
R1176 B.n430 B.n87 163.367
R1177 B.n431 B.n430 163.367
R1178 B.n432 B.n431 163.367
R1179 B.n432 B.n85 163.367
R1180 B.n436 B.n85 163.367
R1181 B.n437 B.n436 163.367
R1182 B.n438 B.n437 163.367
R1183 B.n438 B.n83 163.367
R1184 B.n442 B.n83 163.367
R1185 B.n443 B.n442 163.367
R1186 B.n444 B.n443 163.367
R1187 B.n444 B.n81 163.367
R1188 B.n448 B.n81 163.367
R1189 B.n449 B.n448 163.367
R1190 B.n450 B.n449 163.367
R1191 B.n450 B.n79 163.367
R1192 B.n454 B.n79 163.367
R1193 B.n455 B.n454 163.367
R1194 B.n456 B.n455 163.367
R1195 B.n456 B.n77 163.367
R1196 B.n460 B.n77 163.367
R1197 B.n461 B.n460 163.367
R1198 B.n462 B.n461 163.367
R1199 B.n462 B.n75 163.367
R1200 B.n466 B.n75 163.367
R1201 B.n467 B.n466 163.367
R1202 B.n468 B.n467 163.367
R1203 B.n468 B.n73 163.367
R1204 B.n472 B.n73 163.367
R1205 B.n473 B.n472 163.367
R1206 B.n474 B.n473 163.367
R1207 B.n474 B.n71 163.367
R1208 B.n478 B.n71 163.367
R1209 B.n479 B.n478 163.367
R1210 B.n480 B.n479 163.367
R1211 B.n480 B.n69 163.367
R1212 B.n484 B.n69 163.367
R1213 B.n485 B.n484 163.367
R1214 B.n486 B.n485 163.367
R1215 B.n486 B.n67 163.367
R1216 B.n490 B.n67 163.367
R1217 B.n491 B.n490 163.367
R1218 B.n492 B.n491 163.367
R1219 B.n492 B.n65 163.367
R1220 B.n496 B.n65 163.367
R1221 B.n497 B.n496 163.367
R1222 B.n498 B.n497 163.367
R1223 B.n498 B.n63 163.367
R1224 B.n502 B.n63 163.367
R1225 B.n595 B.n594 163.367
R1226 B.n594 B.n29 163.367
R1227 B.n590 B.n29 163.367
R1228 B.n590 B.n589 163.367
R1229 B.n589 B.n588 163.367
R1230 B.n588 B.n31 163.367
R1231 B.n584 B.n31 163.367
R1232 B.n584 B.n583 163.367
R1233 B.n583 B.n582 163.367
R1234 B.n582 B.n33 163.367
R1235 B.n578 B.n33 163.367
R1236 B.n578 B.n577 163.367
R1237 B.n577 B.n576 163.367
R1238 B.n576 B.n35 163.367
R1239 B.n572 B.n35 163.367
R1240 B.n572 B.n571 163.367
R1241 B.n571 B.n570 163.367
R1242 B.n570 B.n37 163.367
R1243 B.n566 B.n37 163.367
R1244 B.n566 B.n565 163.367
R1245 B.n565 B.n564 163.367
R1246 B.n564 B.n39 163.367
R1247 B.n560 B.n39 163.367
R1248 B.n560 B.n559 163.367
R1249 B.n559 B.n558 163.367
R1250 B.n558 B.n41 163.367
R1251 B.n553 B.n41 163.367
R1252 B.n553 B.n552 163.367
R1253 B.n552 B.n551 163.367
R1254 B.n551 B.n45 163.367
R1255 B.n547 B.n45 163.367
R1256 B.n547 B.n546 163.367
R1257 B.n546 B.n545 163.367
R1258 B.n545 B.n47 163.367
R1259 B.n540 B.n47 163.367
R1260 B.n540 B.n539 163.367
R1261 B.n539 B.n538 163.367
R1262 B.n538 B.n51 163.367
R1263 B.n534 B.n51 163.367
R1264 B.n534 B.n533 163.367
R1265 B.n533 B.n532 163.367
R1266 B.n532 B.n53 163.367
R1267 B.n528 B.n53 163.367
R1268 B.n528 B.n527 163.367
R1269 B.n527 B.n526 163.367
R1270 B.n526 B.n55 163.367
R1271 B.n522 B.n55 163.367
R1272 B.n522 B.n521 163.367
R1273 B.n521 B.n520 163.367
R1274 B.n520 B.n57 163.367
R1275 B.n516 B.n57 163.367
R1276 B.n516 B.n515 163.367
R1277 B.n515 B.n514 163.367
R1278 B.n514 B.n59 163.367
R1279 B.n510 B.n59 163.367
R1280 B.n510 B.n509 163.367
R1281 B.n509 B.n508 163.367
R1282 B.n508 B.n61 163.367
R1283 B.n504 B.n61 163.367
R1284 B.n504 B.n503 163.367
R1285 B.n129 B.n128 72.146
R1286 B.n137 B.n136 72.146
R1287 B.n43 B.n42 72.146
R1288 B.n49 B.n48 72.146
R1289 B.n130 B.n129 59.5399
R1290 B.n291 B.n137 59.5399
R1291 B.n556 B.n43 59.5399
R1292 B.n542 B.n49 59.5399
R1293 B.n597 B.n28 31.6883
R1294 B.n501 B.n62 31.6883
R1295 B.n345 B.n344 31.6883
R1296 B.n253 B.n150 31.6883
R1297 B B.n675 18.0485
R1298 B.n593 B.n28 10.6151
R1299 B.n593 B.n592 10.6151
R1300 B.n592 B.n591 10.6151
R1301 B.n591 B.n30 10.6151
R1302 B.n587 B.n30 10.6151
R1303 B.n587 B.n586 10.6151
R1304 B.n586 B.n585 10.6151
R1305 B.n585 B.n32 10.6151
R1306 B.n581 B.n32 10.6151
R1307 B.n581 B.n580 10.6151
R1308 B.n580 B.n579 10.6151
R1309 B.n579 B.n34 10.6151
R1310 B.n575 B.n34 10.6151
R1311 B.n575 B.n574 10.6151
R1312 B.n574 B.n573 10.6151
R1313 B.n573 B.n36 10.6151
R1314 B.n569 B.n36 10.6151
R1315 B.n569 B.n568 10.6151
R1316 B.n568 B.n567 10.6151
R1317 B.n567 B.n38 10.6151
R1318 B.n563 B.n38 10.6151
R1319 B.n563 B.n562 10.6151
R1320 B.n562 B.n561 10.6151
R1321 B.n561 B.n40 10.6151
R1322 B.n557 B.n40 10.6151
R1323 B.n555 B.n554 10.6151
R1324 B.n554 B.n44 10.6151
R1325 B.n550 B.n44 10.6151
R1326 B.n550 B.n549 10.6151
R1327 B.n549 B.n548 10.6151
R1328 B.n548 B.n46 10.6151
R1329 B.n544 B.n46 10.6151
R1330 B.n544 B.n543 10.6151
R1331 B.n541 B.n50 10.6151
R1332 B.n537 B.n50 10.6151
R1333 B.n537 B.n536 10.6151
R1334 B.n536 B.n535 10.6151
R1335 B.n535 B.n52 10.6151
R1336 B.n531 B.n52 10.6151
R1337 B.n531 B.n530 10.6151
R1338 B.n530 B.n529 10.6151
R1339 B.n529 B.n54 10.6151
R1340 B.n525 B.n54 10.6151
R1341 B.n525 B.n524 10.6151
R1342 B.n524 B.n523 10.6151
R1343 B.n523 B.n56 10.6151
R1344 B.n519 B.n56 10.6151
R1345 B.n519 B.n518 10.6151
R1346 B.n518 B.n517 10.6151
R1347 B.n517 B.n58 10.6151
R1348 B.n513 B.n58 10.6151
R1349 B.n513 B.n512 10.6151
R1350 B.n512 B.n511 10.6151
R1351 B.n511 B.n60 10.6151
R1352 B.n507 B.n60 10.6151
R1353 B.n507 B.n506 10.6151
R1354 B.n506 B.n505 10.6151
R1355 B.n505 B.n62 10.6151
R1356 B.n345 B.n114 10.6151
R1357 B.n349 B.n114 10.6151
R1358 B.n350 B.n349 10.6151
R1359 B.n351 B.n350 10.6151
R1360 B.n351 B.n112 10.6151
R1361 B.n355 B.n112 10.6151
R1362 B.n356 B.n355 10.6151
R1363 B.n357 B.n356 10.6151
R1364 B.n357 B.n110 10.6151
R1365 B.n361 B.n110 10.6151
R1366 B.n362 B.n361 10.6151
R1367 B.n363 B.n362 10.6151
R1368 B.n363 B.n108 10.6151
R1369 B.n367 B.n108 10.6151
R1370 B.n368 B.n367 10.6151
R1371 B.n369 B.n368 10.6151
R1372 B.n369 B.n106 10.6151
R1373 B.n373 B.n106 10.6151
R1374 B.n374 B.n373 10.6151
R1375 B.n375 B.n374 10.6151
R1376 B.n375 B.n104 10.6151
R1377 B.n379 B.n104 10.6151
R1378 B.n380 B.n379 10.6151
R1379 B.n381 B.n380 10.6151
R1380 B.n381 B.n102 10.6151
R1381 B.n385 B.n102 10.6151
R1382 B.n386 B.n385 10.6151
R1383 B.n387 B.n386 10.6151
R1384 B.n387 B.n100 10.6151
R1385 B.n391 B.n100 10.6151
R1386 B.n392 B.n391 10.6151
R1387 B.n393 B.n392 10.6151
R1388 B.n393 B.n98 10.6151
R1389 B.n397 B.n98 10.6151
R1390 B.n398 B.n397 10.6151
R1391 B.n399 B.n398 10.6151
R1392 B.n399 B.n96 10.6151
R1393 B.n403 B.n96 10.6151
R1394 B.n404 B.n403 10.6151
R1395 B.n405 B.n404 10.6151
R1396 B.n405 B.n94 10.6151
R1397 B.n409 B.n94 10.6151
R1398 B.n410 B.n409 10.6151
R1399 B.n411 B.n410 10.6151
R1400 B.n411 B.n92 10.6151
R1401 B.n415 B.n92 10.6151
R1402 B.n416 B.n415 10.6151
R1403 B.n417 B.n416 10.6151
R1404 B.n417 B.n90 10.6151
R1405 B.n421 B.n90 10.6151
R1406 B.n422 B.n421 10.6151
R1407 B.n423 B.n422 10.6151
R1408 B.n423 B.n88 10.6151
R1409 B.n427 B.n88 10.6151
R1410 B.n428 B.n427 10.6151
R1411 B.n429 B.n428 10.6151
R1412 B.n429 B.n86 10.6151
R1413 B.n433 B.n86 10.6151
R1414 B.n434 B.n433 10.6151
R1415 B.n435 B.n434 10.6151
R1416 B.n435 B.n84 10.6151
R1417 B.n439 B.n84 10.6151
R1418 B.n440 B.n439 10.6151
R1419 B.n441 B.n440 10.6151
R1420 B.n441 B.n82 10.6151
R1421 B.n445 B.n82 10.6151
R1422 B.n446 B.n445 10.6151
R1423 B.n447 B.n446 10.6151
R1424 B.n447 B.n80 10.6151
R1425 B.n451 B.n80 10.6151
R1426 B.n452 B.n451 10.6151
R1427 B.n453 B.n452 10.6151
R1428 B.n453 B.n78 10.6151
R1429 B.n457 B.n78 10.6151
R1430 B.n458 B.n457 10.6151
R1431 B.n459 B.n458 10.6151
R1432 B.n459 B.n76 10.6151
R1433 B.n463 B.n76 10.6151
R1434 B.n464 B.n463 10.6151
R1435 B.n465 B.n464 10.6151
R1436 B.n465 B.n74 10.6151
R1437 B.n469 B.n74 10.6151
R1438 B.n470 B.n469 10.6151
R1439 B.n471 B.n470 10.6151
R1440 B.n471 B.n72 10.6151
R1441 B.n475 B.n72 10.6151
R1442 B.n476 B.n475 10.6151
R1443 B.n477 B.n476 10.6151
R1444 B.n477 B.n70 10.6151
R1445 B.n481 B.n70 10.6151
R1446 B.n482 B.n481 10.6151
R1447 B.n483 B.n482 10.6151
R1448 B.n483 B.n68 10.6151
R1449 B.n487 B.n68 10.6151
R1450 B.n488 B.n487 10.6151
R1451 B.n489 B.n488 10.6151
R1452 B.n489 B.n66 10.6151
R1453 B.n493 B.n66 10.6151
R1454 B.n494 B.n493 10.6151
R1455 B.n495 B.n494 10.6151
R1456 B.n495 B.n64 10.6151
R1457 B.n499 B.n64 10.6151
R1458 B.n500 B.n499 10.6151
R1459 B.n501 B.n500 10.6151
R1460 B.n254 B.n253 10.6151
R1461 B.n255 B.n254 10.6151
R1462 B.n255 B.n148 10.6151
R1463 B.n259 B.n148 10.6151
R1464 B.n260 B.n259 10.6151
R1465 B.n261 B.n260 10.6151
R1466 B.n261 B.n146 10.6151
R1467 B.n265 B.n146 10.6151
R1468 B.n266 B.n265 10.6151
R1469 B.n267 B.n266 10.6151
R1470 B.n267 B.n144 10.6151
R1471 B.n271 B.n144 10.6151
R1472 B.n272 B.n271 10.6151
R1473 B.n273 B.n272 10.6151
R1474 B.n273 B.n142 10.6151
R1475 B.n277 B.n142 10.6151
R1476 B.n278 B.n277 10.6151
R1477 B.n279 B.n278 10.6151
R1478 B.n279 B.n140 10.6151
R1479 B.n283 B.n140 10.6151
R1480 B.n284 B.n283 10.6151
R1481 B.n285 B.n284 10.6151
R1482 B.n285 B.n138 10.6151
R1483 B.n289 B.n138 10.6151
R1484 B.n290 B.n289 10.6151
R1485 B.n292 B.n134 10.6151
R1486 B.n296 B.n134 10.6151
R1487 B.n297 B.n296 10.6151
R1488 B.n298 B.n297 10.6151
R1489 B.n298 B.n132 10.6151
R1490 B.n302 B.n132 10.6151
R1491 B.n303 B.n302 10.6151
R1492 B.n304 B.n303 10.6151
R1493 B.n308 B.n307 10.6151
R1494 B.n309 B.n308 10.6151
R1495 B.n309 B.n126 10.6151
R1496 B.n313 B.n126 10.6151
R1497 B.n314 B.n313 10.6151
R1498 B.n315 B.n314 10.6151
R1499 B.n315 B.n124 10.6151
R1500 B.n319 B.n124 10.6151
R1501 B.n320 B.n319 10.6151
R1502 B.n321 B.n320 10.6151
R1503 B.n321 B.n122 10.6151
R1504 B.n325 B.n122 10.6151
R1505 B.n326 B.n325 10.6151
R1506 B.n327 B.n326 10.6151
R1507 B.n327 B.n120 10.6151
R1508 B.n331 B.n120 10.6151
R1509 B.n332 B.n331 10.6151
R1510 B.n333 B.n332 10.6151
R1511 B.n333 B.n118 10.6151
R1512 B.n337 B.n118 10.6151
R1513 B.n338 B.n337 10.6151
R1514 B.n339 B.n338 10.6151
R1515 B.n339 B.n116 10.6151
R1516 B.n343 B.n116 10.6151
R1517 B.n344 B.n343 10.6151
R1518 B.n249 B.n150 10.6151
R1519 B.n249 B.n248 10.6151
R1520 B.n248 B.n247 10.6151
R1521 B.n247 B.n152 10.6151
R1522 B.n243 B.n152 10.6151
R1523 B.n243 B.n242 10.6151
R1524 B.n242 B.n241 10.6151
R1525 B.n241 B.n154 10.6151
R1526 B.n237 B.n154 10.6151
R1527 B.n237 B.n236 10.6151
R1528 B.n236 B.n235 10.6151
R1529 B.n235 B.n156 10.6151
R1530 B.n231 B.n156 10.6151
R1531 B.n231 B.n230 10.6151
R1532 B.n230 B.n229 10.6151
R1533 B.n229 B.n158 10.6151
R1534 B.n225 B.n158 10.6151
R1535 B.n225 B.n224 10.6151
R1536 B.n224 B.n223 10.6151
R1537 B.n223 B.n160 10.6151
R1538 B.n219 B.n160 10.6151
R1539 B.n219 B.n218 10.6151
R1540 B.n218 B.n217 10.6151
R1541 B.n217 B.n162 10.6151
R1542 B.n213 B.n162 10.6151
R1543 B.n213 B.n212 10.6151
R1544 B.n212 B.n211 10.6151
R1545 B.n211 B.n164 10.6151
R1546 B.n207 B.n164 10.6151
R1547 B.n207 B.n206 10.6151
R1548 B.n206 B.n205 10.6151
R1549 B.n205 B.n166 10.6151
R1550 B.n201 B.n166 10.6151
R1551 B.n201 B.n200 10.6151
R1552 B.n200 B.n199 10.6151
R1553 B.n199 B.n168 10.6151
R1554 B.n195 B.n168 10.6151
R1555 B.n195 B.n194 10.6151
R1556 B.n194 B.n193 10.6151
R1557 B.n193 B.n170 10.6151
R1558 B.n189 B.n170 10.6151
R1559 B.n189 B.n188 10.6151
R1560 B.n188 B.n187 10.6151
R1561 B.n187 B.n172 10.6151
R1562 B.n183 B.n172 10.6151
R1563 B.n183 B.n182 10.6151
R1564 B.n182 B.n181 10.6151
R1565 B.n181 B.n174 10.6151
R1566 B.n177 B.n174 10.6151
R1567 B.n177 B.n176 10.6151
R1568 B.n176 B.n0 10.6151
R1569 B.n671 B.n1 10.6151
R1570 B.n671 B.n670 10.6151
R1571 B.n670 B.n669 10.6151
R1572 B.n669 B.n4 10.6151
R1573 B.n665 B.n4 10.6151
R1574 B.n665 B.n664 10.6151
R1575 B.n664 B.n663 10.6151
R1576 B.n663 B.n6 10.6151
R1577 B.n659 B.n6 10.6151
R1578 B.n659 B.n658 10.6151
R1579 B.n658 B.n657 10.6151
R1580 B.n657 B.n8 10.6151
R1581 B.n653 B.n8 10.6151
R1582 B.n653 B.n652 10.6151
R1583 B.n652 B.n651 10.6151
R1584 B.n651 B.n10 10.6151
R1585 B.n647 B.n10 10.6151
R1586 B.n647 B.n646 10.6151
R1587 B.n646 B.n645 10.6151
R1588 B.n645 B.n12 10.6151
R1589 B.n641 B.n12 10.6151
R1590 B.n641 B.n640 10.6151
R1591 B.n640 B.n639 10.6151
R1592 B.n639 B.n14 10.6151
R1593 B.n635 B.n14 10.6151
R1594 B.n635 B.n634 10.6151
R1595 B.n634 B.n633 10.6151
R1596 B.n633 B.n16 10.6151
R1597 B.n629 B.n16 10.6151
R1598 B.n629 B.n628 10.6151
R1599 B.n628 B.n627 10.6151
R1600 B.n627 B.n18 10.6151
R1601 B.n623 B.n18 10.6151
R1602 B.n623 B.n622 10.6151
R1603 B.n622 B.n621 10.6151
R1604 B.n621 B.n20 10.6151
R1605 B.n617 B.n20 10.6151
R1606 B.n617 B.n616 10.6151
R1607 B.n616 B.n615 10.6151
R1608 B.n615 B.n22 10.6151
R1609 B.n611 B.n22 10.6151
R1610 B.n611 B.n610 10.6151
R1611 B.n610 B.n609 10.6151
R1612 B.n609 B.n24 10.6151
R1613 B.n605 B.n24 10.6151
R1614 B.n605 B.n604 10.6151
R1615 B.n604 B.n603 10.6151
R1616 B.n603 B.n26 10.6151
R1617 B.n599 B.n26 10.6151
R1618 B.n599 B.n598 10.6151
R1619 B.n598 B.n597 10.6151
R1620 B.n556 B.n555 6.5566
R1621 B.n543 B.n542 6.5566
R1622 B.n292 B.n291 6.5566
R1623 B.n304 B.n130 6.5566
R1624 B.n557 B.n556 4.05904
R1625 B.n542 B.n541 4.05904
R1626 B.n291 B.n290 4.05904
R1627 B.n307 B.n130 4.05904
R1628 B.n675 B.n0 2.81026
R1629 B.n675 B.n1 2.81026
C0 VDD2 VDD1 1.71497f
C1 VDD2 VP 0.525003f
C2 VDD2 B 1.95967f
C3 VDD2 w_n3946_n2290# 2.22431f
C4 VDD1 VP 4.42446f
C5 VDD1 B 1.86664f
C6 B VP 2.12744f
C7 VDD1 w_n3946_n2290# 2.11398f
C8 VDD2 VN 4.05363f
C9 VP w_n3946_n2290# 8.08367f
C10 B w_n3946_n2290# 9.26337f
C11 VDD1 VN 0.151859f
C12 VN VP 6.69852f
C13 VDD2 VTAIL 6.25289f
C14 VN B 1.26802f
C15 VN w_n3946_n2290# 7.57131f
C16 VDD1 VTAIL 6.19511f
C17 VTAIL VP 4.84188f
C18 VTAIL B 2.72421f
C19 VTAIL w_n3946_n2290# 2.30957f
C20 VN VTAIL 4.82771f
C21 VDD2 VSUBS 1.834136f
C22 VDD1 VSUBS 1.902195f
C23 VTAIL VSUBS 0.782475f
C24 VN VSUBS 6.37693f
C25 VP VSUBS 3.168071f
C26 B VSUBS 4.962208f
C27 w_n3946_n2290# VSUBS 0.112556p
C28 B.n0 VSUBS 0.005365f
C29 B.n1 VSUBS 0.005365f
C30 B.n2 VSUBS 0.008485f
C31 B.n3 VSUBS 0.008485f
C32 B.n4 VSUBS 0.008485f
C33 B.n5 VSUBS 0.008485f
C34 B.n6 VSUBS 0.008485f
C35 B.n7 VSUBS 0.008485f
C36 B.n8 VSUBS 0.008485f
C37 B.n9 VSUBS 0.008485f
C38 B.n10 VSUBS 0.008485f
C39 B.n11 VSUBS 0.008485f
C40 B.n12 VSUBS 0.008485f
C41 B.n13 VSUBS 0.008485f
C42 B.n14 VSUBS 0.008485f
C43 B.n15 VSUBS 0.008485f
C44 B.n16 VSUBS 0.008485f
C45 B.n17 VSUBS 0.008485f
C46 B.n18 VSUBS 0.008485f
C47 B.n19 VSUBS 0.008485f
C48 B.n20 VSUBS 0.008485f
C49 B.n21 VSUBS 0.008485f
C50 B.n22 VSUBS 0.008485f
C51 B.n23 VSUBS 0.008485f
C52 B.n24 VSUBS 0.008485f
C53 B.n25 VSUBS 0.008485f
C54 B.n26 VSUBS 0.008485f
C55 B.n27 VSUBS 0.008485f
C56 B.n28 VSUBS 0.019805f
C57 B.n29 VSUBS 0.008485f
C58 B.n30 VSUBS 0.008485f
C59 B.n31 VSUBS 0.008485f
C60 B.n32 VSUBS 0.008485f
C61 B.n33 VSUBS 0.008485f
C62 B.n34 VSUBS 0.008485f
C63 B.n35 VSUBS 0.008485f
C64 B.n36 VSUBS 0.008485f
C65 B.n37 VSUBS 0.008485f
C66 B.n38 VSUBS 0.008485f
C67 B.n39 VSUBS 0.008485f
C68 B.n40 VSUBS 0.008485f
C69 B.n41 VSUBS 0.008485f
C70 B.t5 VSUBS 0.121487f
C71 B.t4 VSUBS 0.161613f
C72 B.t3 VSUBS 1.29496f
C73 B.n42 VSUBS 0.26801f
C74 B.n43 VSUBS 0.207308f
C75 B.n44 VSUBS 0.008485f
C76 B.n45 VSUBS 0.008485f
C77 B.n46 VSUBS 0.008485f
C78 B.n47 VSUBS 0.008485f
C79 B.t8 VSUBS 0.12149f
C80 B.t7 VSUBS 0.161615f
C81 B.t6 VSUBS 1.29496f
C82 B.n48 VSUBS 0.268008f
C83 B.n49 VSUBS 0.207306f
C84 B.n50 VSUBS 0.008485f
C85 B.n51 VSUBS 0.008485f
C86 B.n52 VSUBS 0.008485f
C87 B.n53 VSUBS 0.008485f
C88 B.n54 VSUBS 0.008485f
C89 B.n55 VSUBS 0.008485f
C90 B.n56 VSUBS 0.008485f
C91 B.n57 VSUBS 0.008485f
C92 B.n58 VSUBS 0.008485f
C93 B.n59 VSUBS 0.008485f
C94 B.n60 VSUBS 0.008485f
C95 B.n61 VSUBS 0.008485f
C96 B.n62 VSUBS 0.018772f
C97 B.n63 VSUBS 0.008485f
C98 B.n64 VSUBS 0.008485f
C99 B.n65 VSUBS 0.008485f
C100 B.n66 VSUBS 0.008485f
C101 B.n67 VSUBS 0.008485f
C102 B.n68 VSUBS 0.008485f
C103 B.n69 VSUBS 0.008485f
C104 B.n70 VSUBS 0.008485f
C105 B.n71 VSUBS 0.008485f
C106 B.n72 VSUBS 0.008485f
C107 B.n73 VSUBS 0.008485f
C108 B.n74 VSUBS 0.008485f
C109 B.n75 VSUBS 0.008485f
C110 B.n76 VSUBS 0.008485f
C111 B.n77 VSUBS 0.008485f
C112 B.n78 VSUBS 0.008485f
C113 B.n79 VSUBS 0.008485f
C114 B.n80 VSUBS 0.008485f
C115 B.n81 VSUBS 0.008485f
C116 B.n82 VSUBS 0.008485f
C117 B.n83 VSUBS 0.008485f
C118 B.n84 VSUBS 0.008485f
C119 B.n85 VSUBS 0.008485f
C120 B.n86 VSUBS 0.008485f
C121 B.n87 VSUBS 0.008485f
C122 B.n88 VSUBS 0.008485f
C123 B.n89 VSUBS 0.008485f
C124 B.n90 VSUBS 0.008485f
C125 B.n91 VSUBS 0.008485f
C126 B.n92 VSUBS 0.008485f
C127 B.n93 VSUBS 0.008485f
C128 B.n94 VSUBS 0.008485f
C129 B.n95 VSUBS 0.008485f
C130 B.n96 VSUBS 0.008485f
C131 B.n97 VSUBS 0.008485f
C132 B.n98 VSUBS 0.008485f
C133 B.n99 VSUBS 0.008485f
C134 B.n100 VSUBS 0.008485f
C135 B.n101 VSUBS 0.008485f
C136 B.n102 VSUBS 0.008485f
C137 B.n103 VSUBS 0.008485f
C138 B.n104 VSUBS 0.008485f
C139 B.n105 VSUBS 0.008485f
C140 B.n106 VSUBS 0.008485f
C141 B.n107 VSUBS 0.008485f
C142 B.n108 VSUBS 0.008485f
C143 B.n109 VSUBS 0.008485f
C144 B.n110 VSUBS 0.008485f
C145 B.n111 VSUBS 0.008485f
C146 B.n112 VSUBS 0.008485f
C147 B.n113 VSUBS 0.008485f
C148 B.n114 VSUBS 0.008485f
C149 B.n115 VSUBS 0.019805f
C150 B.n116 VSUBS 0.008485f
C151 B.n117 VSUBS 0.008485f
C152 B.n118 VSUBS 0.008485f
C153 B.n119 VSUBS 0.008485f
C154 B.n120 VSUBS 0.008485f
C155 B.n121 VSUBS 0.008485f
C156 B.n122 VSUBS 0.008485f
C157 B.n123 VSUBS 0.008485f
C158 B.n124 VSUBS 0.008485f
C159 B.n125 VSUBS 0.008485f
C160 B.n126 VSUBS 0.008485f
C161 B.n127 VSUBS 0.008485f
C162 B.t10 VSUBS 0.12149f
C163 B.t11 VSUBS 0.161615f
C164 B.t9 VSUBS 1.29496f
C165 B.n128 VSUBS 0.268008f
C166 B.n129 VSUBS 0.207306f
C167 B.n130 VSUBS 0.019659f
C168 B.n131 VSUBS 0.008485f
C169 B.n132 VSUBS 0.008485f
C170 B.n133 VSUBS 0.008485f
C171 B.n134 VSUBS 0.008485f
C172 B.n135 VSUBS 0.008485f
C173 B.t1 VSUBS 0.121487f
C174 B.t2 VSUBS 0.161613f
C175 B.t0 VSUBS 1.29496f
C176 B.n136 VSUBS 0.26801f
C177 B.n137 VSUBS 0.207308f
C178 B.n138 VSUBS 0.008485f
C179 B.n139 VSUBS 0.008485f
C180 B.n140 VSUBS 0.008485f
C181 B.n141 VSUBS 0.008485f
C182 B.n142 VSUBS 0.008485f
C183 B.n143 VSUBS 0.008485f
C184 B.n144 VSUBS 0.008485f
C185 B.n145 VSUBS 0.008485f
C186 B.n146 VSUBS 0.008485f
C187 B.n147 VSUBS 0.008485f
C188 B.n148 VSUBS 0.008485f
C189 B.n149 VSUBS 0.008485f
C190 B.n150 VSUBS 0.019125f
C191 B.n151 VSUBS 0.008485f
C192 B.n152 VSUBS 0.008485f
C193 B.n153 VSUBS 0.008485f
C194 B.n154 VSUBS 0.008485f
C195 B.n155 VSUBS 0.008485f
C196 B.n156 VSUBS 0.008485f
C197 B.n157 VSUBS 0.008485f
C198 B.n158 VSUBS 0.008485f
C199 B.n159 VSUBS 0.008485f
C200 B.n160 VSUBS 0.008485f
C201 B.n161 VSUBS 0.008485f
C202 B.n162 VSUBS 0.008485f
C203 B.n163 VSUBS 0.008485f
C204 B.n164 VSUBS 0.008485f
C205 B.n165 VSUBS 0.008485f
C206 B.n166 VSUBS 0.008485f
C207 B.n167 VSUBS 0.008485f
C208 B.n168 VSUBS 0.008485f
C209 B.n169 VSUBS 0.008485f
C210 B.n170 VSUBS 0.008485f
C211 B.n171 VSUBS 0.008485f
C212 B.n172 VSUBS 0.008485f
C213 B.n173 VSUBS 0.008485f
C214 B.n174 VSUBS 0.008485f
C215 B.n175 VSUBS 0.008485f
C216 B.n176 VSUBS 0.008485f
C217 B.n177 VSUBS 0.008485f
C218 B.n178 VSUBS 0.008485f
C219 B.n179 VSUBS 0.008485f
C220 B.n180 VSUBS 0.008485f
C221 B.n181 VSUBS 0.008485f
C222 B.n182 VSUBS 0.008485f
C223 B.n183 VSUBS 0.008485f
C224 B.n184 VSUBS 0.008485f
C225 B.n185 VSUBS 0.008485f
C226 B.n186 VSUBS 0.008485f
C227 B.n187 VSUBS 0.008485f
C228 B.n188 VSUBS 0.008485f
C229 B.n189 VSUBS 0.008485f
C230 B.n190 VSUBS 0.008485f
C231 B.n191 VSUBS 0.008485f
C232 B.n192 VSUBS 0.008485f
C233 B.n193 VSUBS 0.008485f
C234 B.n194 VSUBS 0.008485f
C235 B.n195 VSUBS 0.008485f
C236 B.n196 VSUBS 0.008485f
C237 B.n197 VSUBS 0.008485f
C238 B.n198 VSUBS 0.008485f
C239 B.n199 VSUBS 0.008485f
C240 B.n200 VSUBS 0.008485f
C241 B.n201 VSUBS 0.008485f
C242 B.n202 VSUBS 0.008485f
C243 B.n203 VSUBS 0.008485f
C244 B.n204 VSUBS 0.008485f
C245 B.n205 VSUBS 0.008485f
C246 B.n206 VSUBS 0.008485f
C247 B.n207 VSUBS 0.008485f
C248 B.n208 VSUBS 0.008485f
C249 B.n209 VSUBS 0.008485f
C250 B.n210 VSUBS 0.008485f
C251 B.n211 VSUBS 0.008485f
C252 B.n212 VSUBS 0.008485f
C253 B.n213 VSUBS 0.008485f
C254 B.n214 VSUBS 0.008485f
C255 B.n215 VSUBS 0.008485f
C256 B.n216 VSUBS 0.008485f
C257 B.n217 VSUBS 0.008485f
C258 B.n218 VSUBS 0.008485f
C259 B.n219 VSUBS 0.008485f
C260 B.n220 VSUBS 0.008485f
C261 B.n221 VSUBS 0.008485f
C262 B.n222 VSUBS 0.008485f
C263 B.n223 VSUBS 0.008485f
C264 B.n224 VSUBS 0.008485f
C265 B.n225 VSUBS 0.008485f
C266 B.n226 VSUBS 0.008485f
C267 B.n227 VSUBS 0.008485f
C268 B.n228 VSUBS 0.008485f
C269 B.n229 VSUBS 0.008485f
C270 B.n230 VSUBS 0.008485f
C271 B.n231 VSUBS 0.008485f
C272 B.n232 VSUBS 0.008485f
C273 B.n233 VSUBS 0.008485f
C274 B.n234 VSUBS 0.008485f
C275 B.n235 VSUBS 0.008485f
C276 B.n236 VSUBS 0.008485f
C277 B.n237 VSUBS 0.008485f
C278 B.n238 VSUBS 0.008485f
C279 B.n239 VSUBS 0.008485f
C280 B.n240 VSUBS 0.008485f
C281 B.n241 VSUBS 0.008485f
C282 B.n242 VSUBS 0.008485f
C283 B.n243 VSUBS 0.008485f
C284 B.n244 VSUBS 0.008485f
C285 B.n245 VSUBS 0.008485f
C286 B.n246 VSUBS 0.008485f
C287 B.n247 VSUBS 0.008485f
C288 B.n248 VSUBS 0.008485f
C289 B.n249 VSUBS 0.008485f
C290 B.n250 VSUBS 0.008485f
C291 B.n251 VSUBS 0.019125f
C292 B.n252 VSUBS 0.019805f
C293 B.n253 VSUBS 0.019805f
C294 B.n254 VSUBS 0.008485f
C295 B.n255 VSUBS 0.008485f
C296 B.n256 VSUBS 0.008485f
C297 B.n257 VSUBS 0.008485f
C298 B.n258 VSUBS 0.008485f
C299 B.n259 VSUBS 0.008485f
C300 B.n260 VSUBS 0.008485f
C301 B.n261 VSUBS 0.008485f
C302 B.n262 VSUBS 0.008485f
C303 B.n263 VSUBS 0.008485f
C304 B.n264 VSUBS 0.008485f
C305 B.n265 VSUBS 0.008485f
C306 B.n266 VSUBS 0.008485f
C307 B.n267 VSUBS 0.008485f
C308 B.n268 VSUBS 0.008485f
C309 B.n269 VSUBS 0.008485f
C310 B.n270 VSUBS 0.008485f
C311 B.n271 VSUBS 0.008485f
C312 B.n272 VSUBS 0.008485f
C313 B.n273 VSUBS 0.008485f
C314 B.n274 VSUBS 0.008485f
C315 B.n275 VSUBS 0.008485f
C316 B.n276 VSUBS 0.008485f
C317 B.n277 VSUBS 0.008485f
C318 B.n278 VSUBS 0.008485f
C319 B.n279 VSUBS 0.008485f
C320 B.n280 VSUBS 0.008485f
C321 B.n281 VSUBS 0.008485f
C322 B.n282 VSUBS 0.008485f
C323 B.n283 VSUBS 0.008485f
C324 B.n284 VSUBS 0.008485f
C325 B.n285 VSUBS 0.008485f
C326 B.n286 VSUBS 0.008485f
C327 B.n287 VSUBS 0.008485f
C328 B.n288 VSUBS 0.008485f
C329 B.n289 VSUBS 0.008485f
C330 B.n290 VSUBS 0.005865f
C331 B.n291 VSUBS 0.019659f
C332 B.n292 VSUBS 0.006863f
C333 B.n293 VSUBS 0.008485f
C334 B.n294 VSUBS 0.008485f
C335 B.n295 VSUBS 0.008485f
C336 B.n296 VSUBS 0.008485f
C337 B.n297 VSUBS 0.008485f
C338 B.n298 VSUBS 0.008485f
C339 B.n299 VSUBS 0.008485f
C340 B.n300 VSUBS 0.008485f
C341 B.n301 VSUBS 0.008485f
C342 B.n302 VSUBS 0.008485f
C343 B.n303 VSUBS 0.008485f
C344 B.n304 VSUBS 0.006863f
C345 B.n305 VSUBS 0.008485f
C346 B.n306 VSUBS 0.008485f
C347 B.n307 VSUBS 0.005865f
C348 B.n308 VSUBS 0.008485f
C349 B.n309 VSUBS 0.008485f
C350 B.n310 VSUBS 0.008485f
C351 B.n311 VSUBS 0.008485f
C352 B.n312 VSUBS 0.008485f
C353 B.n313 VSUBS 0.008485f
C354 B.n314 VSUBS 0.008485f
C355 B.n315 VSUBS 0.008485f
C356 B.n316 VSUBS 0.008485f
C357 B.n317 VSUBS 0.008485f
C358 B.n318 VSUBS 0.008485f
C359 B.n319 VSUBS 0.008485f
C360 B.n320 VSUBS 0.008485f
C361 B.n321 VSUBS 0.008485f
C362 B.n322 VSUBS 0.008485f
C363 B.n323 VSUBS 0.008485f
C364 B.n324 VSUBS 0.008485f
C365 B.n325 VSUBS 0.008485f
C366 B.n326 VSUBS 0.008485f
C367 B.n327 VSUBS 0.008485f
C368 B.n328 VSUBS 0.008485f
C369 B.n329 VSUBS 0.008485f
C370 B.n330 VSUBS 0.008485f
C371 B.n331 VSUBS 0.008485f
C372 B.n332 VSUBS 0.008485f
C373 B.n333 VSUBS 0.008485f
C374 B.n334 VSUBS 0.008485f
C375 B.n335 VSUBS 0.008485f
C376 B.n336 VSUBS 0.008485f
C377 B.n337 VSUBS 0.008485f
C378 B.n338 VSUBS 0.008485f
C379 B.n339 VSUBS 0.008485f
C380 B.n340 VSUBS 0.008485f
C381 B.n341 VSUBS 0.008485f
C382 B.n342 VSUBS 0.008485f
C383 B.n343 VSUBS 0.008485f
C384 B.n344 VSUBS 0.019805f
C385 B.n345 VSUBS 0.019125f
C386 B.n346 VSUBS 0.019125f
C387 B.n347 VSUBS 0.008485f
C388 B.n348 VSUBS 0.008485f
C389 B.n349 VSUBS 0.008485f
C390 B.n350 VSUBS 0.008485f
C391 B.n351 VSUBS 0.008485f
C392 B.n352 VSUBS 0.008485f
C393 B.n353 VSUBS 0.008485f
C394 B.n354 VSUBS 0.008485f
C395 B.n355 VSUBS 0.008485f
C396 B.n356 VSUBS 0.008485f
C397 B.n357 VSUBS 0.008485f
C398 B.n358 VSUBS 0.008485f
C399 B.n359 VSUBS 0.008485f
C400 B.n360 VSUBS 0.008485f
C401 B.n361 VSUBS 0.008485f
C402 B.n362 VSUBS 0.008485f
C403 B.n363 VSUBS 0.008485f
C404 B.n364 VSUBS 0.008485f
C405 B.n365 VSUBS 0.008485f
C406 B.n366 VSUBS 0.008485f
C407 B.n367 VSUBS 0.008485f
C408 B.n368 VSUBS 0.008485f
C409 B.n369 VSUBS 0.008485f
C410 B.n370 VSUBS 0.008485f
C411 B.n371 VSUBS 0.008485f
C412 B.n372 VSUBS 0.008485f
C413 B.n373 VSUBS 0.008485f
C414 B.n374 VSUBS 0.008485f
C415 B.n375 VSUBS 0.008485f
C416 B.n376 VSUBS 0.008485f
C417 B.n377 VSUBS 0.008485f
C418 B.n378 VSUBS 0.008485f
C419 B.n379 VSUBS 0.008485f
C420 B.n380 VSUBS 0.008485f
C421 B.n381 VSUBS 0.008485f
C422 B.n382 VSUBS 0.008485f
C423 B.n383 VSUBS 0.008485f
C424 B.n384 VSUBS 0.008485f
C425 B.n385 VSUBS 0.008485f
C426 B.n386 VSUBS 0.008485f
C427 B.n387 VSUBS 0.008485f
C428 B.n388 VSUBS 0.008485f
C429 B.n389 VSUBS 0.008485f
C430 B.n390 VSUBS 0.008485f
C431 B.n391 VSUBS 0.008485f
C432 B.n392 VSUBS 0.008485f
C433 B.n393 VSUBS 0.008485f
C434 B.n394 VSUBS 0.008485f
C435 B.n395 VSUBS 0.008485f
C436 B.n396 VSUBS 0.008485f
C437 B.n397 VSUBS 0.008485f
C438 B.n398 VSUBS 0.008485f
C439 B.n399 VSUBS 0.008485f
C440 B.n400 VSUBS 0.008485f
C441 B.n401 VSUBS 0.008485f
C442 B.n402 VSUBS 0.008485f
C443 B.n403 VSUBS 0.008485f
C444 B.n404 VSUBS 0.008485f
C445 B.n405 VSUBS 0.008485f
C446 B.n406 VSUBS 0.008485f
C447 B.n407 VSUBS 0.008485f
C448 B.n408 VSUBS 0.008485f
C449 B.n409 VSUBS 0.008485f
C450 B.n410 VSUBS 0.008485f
C451 B.n411 VSUBS 0.008485f
C452 B.n412 VSUBS 0.008485f
C453 B.n413 VSUBS 0.008485f
C454 B.n414 VSUBS 0.008485f
C455 B.n415 VSUBS 0.008485f
C456 B.n416 VSUBS 0.008485f
C457 B.n417 VSUBS 0.008485f
C458 B.n418 VSUBS 0.008485f
C459 B.n419 VSUBS 0.008485f
C460 B.n420 VSUBS 0.008485f
C461 B.n421 VSUBS 0.008485f
C462 B.n422 VSUBS 0.008485f
C463 B.n423 VSUBS 0.008485f
C464 B.n424 VSUBS 0.008485f
C465 B.n425 VSUBS 0.008485f
C466 B.n426 VSUBS 0.008485f
C467 B.n427 VSUBS 0.008485f
C468 B.n428 VSUBS 0.008485f
C469 B.n429 VSUBS 0.008485f
C470 B.n430 VSUBS 0.008485f
C471 B.n431 VSUBS 0.008485f
C472 B.n432 VSUBS 0.008485f
C473 B.n433 VSUBS 0.008485f
C474 B.n434 VSUBS 0.008485f
C475 B.n435 VSUBS 0.008485f
C476 B.n436 VSUBS 0.008485f
C477 B.n437 VSUBS 0.008485f
C478 B.n438 VSUBS 0.008485f
C479 B.n439 VSUBS 0.008485f
C480 B.n440 VSUBS 0.008485f
C481 B.n441 VSUBS 0.008485f
C482 B.n442 VSUBS 0.008485f
C483 B.n443 VSUBS 0.008485f
C484 B.n444 VSUBS 0.008485f
C485 B.n445 VSUBS 0.008485f
C486 B.n446 VSUBS 0.008485f
C487 B.n447 VSUBS 0.008485f
C488 B.n448 VSUBS 0.008485f
C489 B.n449 VSUBS 0.008485f
C490 B.n450 VSUBS 0.008485f
C491 B.n451 VSUBS 0.008485f
C492 B.n452 VSUBS 0.008485f
C493 B.n453 VSUBS 0.008485f
C494 B.n454 VSUBS 0.008485f
C495 B.n455 VSUBS 0.008485f
C496 B.n456 VSUBS 0.008485f
C497 B.n457 VSUBS 0.008485f
C498 B.n458 VSUBS 0.008485f
C499 B.n459 VSUBS 0.008485f
C500 B.n460 VSUBS 0.008485f
C501 B.n461 VSUBS 0.008485f
C502 B.n462 VSUBS 0.008485f
C503 B.n463 VSUBS 0.008485f
C504 B.n464 VSUBS 0.008485f
C505 B.n465 VSUBS 0.008485f
C506 B.n466 VSUBS 0.008485f
C507 B.n467 VSUBS 0.008485f
C508 B.n468 VSUBS 0.008485f
C509 B.n469 VSUBS 0.008485f
C510 B.n470 VSUBS 0.008485f
C511 B.n471 VSUBS 0.008485f
C512 B.n472 VSUBS 0.008485f
C513 B.n473 VSUBS 0.008485f
C514 B.n474 VSUBS 0.008485f
C515 B.n475 VSUBS 0.008485f
C516 B.n476 VSUBS 0.008485f
C517 B.n477 VSUBS 0.008485f
C518 B.n478 VSUBS 0.008485f
C519 B.n479 VSUBS 0.008485f
C520 B.n480 VSUBS 0.008485f
C521 B.n481 VSUBS 0.008485f
C522 B.n482 VSUBS 0.008485f
C523 B.n483 VSUBS 0.008485f
C524 B.n484 VSUBS 0.008485f
C525 B.n485 VSUBS 0.008485f
C526 B.n486 VSUBS 0.008485f
C527 B.n487 VSUBS 0.008485f
C528 B.n488 VSUBS 0.008485f
C529 B.n489 VSUBS 0.008485f
C530 B.n490 VSUBS 0.008485f
C531 B.n491 VSUBS 0.008485f
C532 B.n492 VSUBS 0.008485f
C533 B.n493 VSUBS 0.008485f
C534 B.n494 VSUBS 0.008485f
C535 B.n495 VSUBS 0.008485f
C536 B.n496 VSUBS 0.008485f
C537 B.n497 VSUBS 0.008485f
C538 B.n498 VSUBS 0.008485f
C539 B.n499 VSUBS 0.008485f
C540 B.n500 VSUBS 0.008485f
C541 B.n501 VSUBS 0.020158f
C542 B.n502 VSUBS 0.019125f
C543 B.n503 VSUBS 0.019805f
C544 B.n504 VSUBS 0.008485f
C545 B.n505 VSUBS 0.008485f
C546 B.n506 VSUBS 0.008485f
C547 B.n507 VSUBS 0.008485f
C548 B.n508 VSUBS 0.008485f
C549 B.n509 VSUBS 0.008485f
C550 B.n510 VSUBS 0.008485f
C551 B.n511 VSUBS 0.008485f
C552 B.n512 VSUBS 0.008485f
C553 B.n513 VSUBS 0.008485f
C554 B.n514 VSUBS 0.008485f
C555 B.n515 VSUBS 0.008485f
C556 B.n516 VSUBS 0.008485f
C557 B.n517 VSUBS 0.008485f
C558 B.n518 VSUBS 0.008485f
C559 B.n519 VSUBS 0.008485f
C560 B.n520 VSUBS 0.008485f
C561 B.n521 VSUBS 0.008485f
C562 B.n522 VSUBS 0.008485f
C563 B.n523 VSUBS 0.008485f
C564 B.n524 VSUBS 0.008485f
C565 B.n525 VSUBS 0.008485f
C566 B.n526 VSUBS 0.008485f
C567 B.n527 VSUBS 0.008485f
C568 B.n528 VSUBS 0.008485f
C569 B.n529 VSUBS 0.008485f
C570 B.n530 VSUBS 0.008485f
C571 B.n531 VSUBS 0.008485f
C572 B.n532 VSUBS 0.008485f
C573 B.n533 VSUBS 0.008485f
C574 B.n534 VSUBS 0.008485f
C575 B.n535 VSUBS 0.008485f
C576 B.n536 VSUBS 0.008485f
C577 B.n537 VSUBS 0.008485f
C578 B.n538 VSUBS 0.008485f
C579 B.n539 VSUBS 0.008485f
C580 B.n540 VSUBS 0.008485f
C581 B.n541 VSUBS 0.005865f
C582 B.n542 VSUBS 0.019659f
C583 B.n543 VSUBS 0.006863f
C584 B.n544 VSUBS 0.008485f
C585 B.n545 VSUBS 0.008485f
C586 B.n546 VSUBS 0.008485f
C587 B.n547 VSUBS 0.008485f
C588 B.n548 VSUBS 0.008485f
C589 B.n549 VSUBS 0.008485f
C590 B.n550 VSUBS 0.008485f
C591 B.n551 VSUBS 0.008485f
C592 B.n552 VSUBS 0.008485f
C593 B.n553 VSUBS 0.008485f
C594 B.n554 VSUBS 0.008485f
C595 B.n555 VSUBS 0.006863f
C596 B.n556 VSUBS 0.019659f
C597 B.n557 VSUBS 0.005865f
C598 B.n558 VSUBS 0.008485f
C599 B.n559 VSUBS 0.008485f
C600 B.n560 VSUBS 0.008485f
C601 B.n561 VSUBS 0.008485f
C602 B.n562 VSUBS 0.008485f
C603 B.n563 VSUBS 0.008485f
C604 B.n564 VSUBS 0.008485f
C605 B.n565 VSUBS 0.008485f
C606 B.n566 VSUBS 0.008485f
C607 B.n567 VSUBS 0.008485f
C608 B.n568 VSUBS 0.008485f
C609 B.n569 VSUBS 0.008485f
C610 B.n570 VSUBS 0.008485f
C611 B.n571 VSUBS 0.008485f
C612 B.n572 VSUBS 0.008485f
C613 B.n573 VSUBS 0.008485f
C614 B.n574 VSUBS 0.008485f
C615 B.n575 VSUBS 0.008485f
C616 B.n576 VSUBS 0.008485f
C617 B.n577 VSUBS 0.008485f
C618 B.n578 VSUBS 0.008485f
C619 B.n579 VSUBS 0.008485f
C620 B.n580 VSUBS 0.008485f
C621 B.n581 VSUBS 0.008485f
C622 B.n582 VSUBS 0.008485f
C623 B.n583 VSUBS 0.008485f
C624 B.n584 VSUBS 0.008485f
C625 B.n585 VSUBS 0.008485f
C626 B.n586 VSUBS 0.008485f
C627 B.n587 VSUBS 0.008485f
C628 B.n588 VSUBS 0.008485f
C629 B.n589 VSUBS 0.008485f
C630 B.n590 VSUBS 0.008485f
C631 B.n591 VSUBS 0.008485f
C632 B.n592 VSUBS 0.008485f
C633 B.n593 VSUBS 0.008485f
C634 B.n594 VSUBS 0.008485f
C635 B.n595 VSUBS 0.019805f
C636 B.n596 VSUBS 0.019125f
C637 B.n597 VSUBS 0.019125f
C638 B.n598 VSUBS 0.008485f
C639 B.n599 VSUBS 0.008485f
C640 B.n600 VSUBS 0.008485f
C641 B.n601 VSUBS 0.008485f
C642 B.n602 VSUBS 0.008485f
C643 B.n603 VSUBS 0.008485f
C644 B.n604 VSUBS 0.008485f
C645 B.n605 VSUBS 0.008485f
C646 B.n606 VSUBS 0.008485f
C647 B.n607 VSUBS 0.008485f
C648 B.n608 VSUBS 0.008485f
C649 B.n609 VSUBS 0.008485f
C650 B.n610 VSUBS 0.008485f
C651 B.n611 VSUBS 0.008485f
C652 B.n612 VSUBS 0.008485f
C653 B.n613 VSUBS 0.008485f
C654 B.n614 VSUBS 0.008485f
C655 B.n615 VSUBS 0.008485f
C656 B.n616 VSUBS 0.008485f
C657 B.n617 VSUBS 0.008485f
C658 B.n618 VSUBS 0.008485f
C659 B.n619 VSUBS 0.008485f
C660 B.n620 VSUBS 0.008485f
C661 B.n621 VSUBS 0.008485f
C662 B.n622 VSUBS 0.008485f
C663 B.n623 VSUBS 0.008485f
C664 B.n624 VSUBS 0.008485f
C665 B.n625 VSUBS 0.008485f
C666 B.n626 VSUBS 0.008485f
C667 B.n627 VSUBS 0.008485f
C668 B.n628 VSUBS 0.008485f
C669 B.n629 VSUBS 0.008485f
C670 B.n630 VSUBS 0.008485f
C671 B.n631 VSUBS 0.008485f
C672 B.n632 VSUBS 0.008485f
C673 B.n633 VSUBS 0.008485f
C674 B.n634 VSUBS 0.008485f
C675 B.n635 VSUBS 0.008485f
C676 B.n636 VSUBS 0.008485f
C677 B.n637 VSUBS 0.008485f
C678 B.n638 VSUBS 0.008485f
C679 B.n639 VSUBS 0.008485f
C680 B.n640 VSUBS 0.008485f
C681 B.n641 VSUBS 0.008485f
C682 B.n642 VSUBS 0.008485f
C683 B.n643 VSUBS 0.008485f
C684 B.n644 VSUBS 0.008485f
C685 B.n645 VSUBS 0.008485f
C686 B.n646 VSUBS 0.008485f
C687 B.n647 VSUBS 0.008485f
C688 B.n648 VSUBS 0.008485f
C689 B.n649 VSUBS 0.008485f
C690 B.n650 VSUBS 0.008485f
C691 B.n651 VSUBS 0.008485f
C692 B.n652 VSUBS 0.008485f
C693 B.n653 VSUBS 0.008485f
C694 B.n654 VSUBS 0.008485f
C695 B.n655 VSUBS 0.008485f
C696 B.n656 VSUBS 0.008485f
C697 B.n657 VSUBS 0.008485f
C698 B.n658 VSUBS 0.008485f
C699 B.n659 VSUBS 0.008485f
C700 B.n660 VSUBS 0.008485f
C701 B.n661 VSUBS 0.008485f
C702 B.n662 VSUBS 0.008485f
C703 B.n663 VSUBS 0.008485f
C704 B.n664 VSUBS 0.008485f
C705 B.n665 VSUBS 0.008485f
C706 B.n666 VSUBS 0.008485f
C707 B.n667 VSUBS 0.008485f
C708 B.n668 VSUBS 0.008485f
C709 B.n669 VSUBS 0.008485f
C710 B.n670 VSUBS 0.008485f
C711 B.n671 VSUBS 0.008485f
C712 B.n672 VSUBS 0.008485f
C713 B.n673 VSUBS 0.008485f
C714 B.n674 VSUBS 0.008485f
C715 B.n675 VSUBS 0.019213f
C716 VDD1.n0 VSUBS 0.028363f
C717 VDD1.n1 VSUBS 0.026634f
C718 VDD1.n2 VSUBS 0.014312f
C719 VDD1.n3 VSUBS 0.033828f
C720 VDD1.n4 VSUBS 0.015154f
C721 VDD1.n5 VSUBS 0.026634f
C722 VDD1.n6 VSUBS 0.014312f
C723 VDD1.n7 VSUBS 0.033828f
C724 VDD1.n8 VSUBS 0.015154f
C725 VDD1.n9 VSUBS 0.685423f
C726 VDD1.n10 VSUBS 0.014312f
C727 VDD1.t3 VSUBS 0.072261f
C728 VDD1.n11 VSUBS 0.122216f
C729 VDD1.n12 VSUBS 0.021516f
C730 VDD1.n13 VSUBS 0.025371f
C731 VDD1.n14 VSUBS 0.033828f
C732 VDD1.n15 VSUBS 0.015154f
C733 VDD1.n16 VSUBS 0.014312f
C734 VDD1.n17 VSUBS 0.026634f
C735 VDD1.n18 VSUBS 0.026634f
C736 VDD1.n19 VSUBS 0.014312f
C737 VDD1.n20 VSUBS 0.015154f
C738 VDD1.n21 VSUBS 0.033828f
C739 VDD1.n22 VSUBS 0.033828f
C740 VDD1.n23 VSUBS 0.015154f
C741 VDD1.n24 VSUBS 0.014312f
C742 VDD1.n25 VSUBS 0.026634f
C743 VDD1.n26 VSUBS 0.026634f
C744 VDD1.n27 VSUBS 0.014312f
C745 VDD1.n28 VSUBS 0.015154f
C746 VDD1.n29 VSUBS 0.033828f
C747 VDD1.n30 VSUBS 0.078824f
C748 VDD1.n31 VSUBS 0.015154f
C749 VDD1.n32 VSUBS 0.014312f
C750 VDD1.n33 VSUBS 0.057561f
C751 VDD1.n34 VSUBS 0.070841f
C752 VDD1.n35 VSUBS 0.028363f
C753 VDD1.n36 VSUBS 0.026634f
C754 VDD1.n37 VSUBS 0.014312f
C755 VDD1.n38 VSUBS 0.033828f
C756 VDD1.n39 VSUBS 0.015154f
C757 VDD1.n40 VSUBS 0.026634f
C758 VDD1.n41 VSUBS 0.014312f
C759 VDD1.n42 VSUBS 0.033828f
C760 VDD1.n43 VSUBS 0.015154f
C761 VDD1.n44 VSUBS 0.685423f
C762 VDD1.n45 VSUBS 0.014312f
C763 VDD1.t4 VSUBS 0.072261f
C764 VDD1.n46 VSUBS 0.122216f
C765 VDD1.n47 VSUBS 0.021516f
C766 VDD1.n48 VSUBS 0.025371f
C767 VDD1.n49 VSUBS 0.033828f
C768 VDD1.n50 VSUBS 0.015154f
C769 VDD1.n51 VSUBS 0.014312f
C770 VDD1.n52 VSUBS 0.026634f
C771 VDD1.n53 VSUBS 0.026634f
C772 VDD1.n54 VSUBS 0.014312f
C773 VDD1.n55 VSUBS 0.015154f
C774 VDD1.n56 VSUBS 0.033828f
C775 VDD1.n57 VSUBS 0.033828f
C776 VDD1.n58 VSUBS 0.015154f
C777 VDD1.n59 VSUBS 0.014312f
C778 VDD1.n60 VSUBS 0.026634f
C779 VDD1.n61 VSUBS 0.026634f
C780 VDD1.n62 VSUBS 0.014312f
C781 VDD1.n63 VSUBS 0.015154f
C782 VDD1.n64 VSUBS 0.033828f
C783 VDD1.n65 VSUBS 0.078824f
C784 VDD1.n66 VSUBS 0.015154f
C785 VDD1.n67 VSUBS 0.014312f
C786 VDD1.n68 VSUBS 0.057561f
C787 VDD1.n69 VSUBS 0.069815f
C788 VDD1.t5 VSUBS 0.139121f
C789 VDD1.t1 VSUBS 0.139121f
C790 VDD1.n70 VSUBS 0.948896f
C791 VDD1.n71 VSUBS 3.24116f
C792 VDD1.t0 VSUBS 0.139121f
C793 VDD1.t2 VSUBS 0.139121f
C794 VDD1.n72 VSUBS 0.942031f
C795 VDD1.n73 VSUBS 2.99841f
C796 VP.t4 VSUBS 2.21693f
C797 VP.n0 VSUBS 0.953362f
C798 VP.n1 VSUBS 0.037178f
C799 VP.n2 VSUBS 0.040603f
C800 VP.n3 VSUBS 0.037178f
C801 VP.t0 VSUBS 2.21693f
C802 VP.n4 VSUBS 0.847511f
C803 VP.n5 VSUBS 0.037178f
C804 VP.n6 VSUBS 0.040603f
C805 VP.n7 VSUBS 0.037178f
C806 VP.t1 VSUBS 2.21693f
C807 VP.n8 VSUBS 0.953362f
C808 VP.t3 VSUBS 2.21693f
C809 VP.n9 VSUBS 0.953362f
C810 VP.n10 VSUBS 0.037178f
C811 VP.n11 VSUBS 0.040603f
C812 VP.n12 VSUBS 0.037178f
C813 VP.t5 VSUBS 2.21693f
C814 VP.n13 VSUBS 0.959093f
C815 VP.t2 VSUBS 2.66969f
C816 VP.n14 VSUBS 0.899116f
C817 VP.n15 VSUBS 0.453904f
C818 VP.n16 VSUBS 0.06929f
C819 VP.n17 VSUBS 0.06929f
C820 VP.n18 VSUBS 0.065165f
C821 VP.n19 VSUBS 0.037178f
C822 VP.n20 VSUBS 0.037178f
C823 VP.n21 VSUBS 0.037178f
C824 VP.n22 VSUBS 0.072067f
C825 VP.n23 VSUBS 0.06929f
C826 VP.n24 VSUBS 0.050133f
C827 VP.n25 VSUBS 0.060004f
C828 VP.n26 VSUBS 1.98526f
C829 VP.n27 VSUBS 2.01324f
C830 VP.n28 VSUBS 0.060004f
C831 VP.n29 VSUBS 0.050133f
C832 VP.n30 VSUBS 0.06929f
C833 VP.n31 VSUBS 0.072067f
C834 VP.n32 VSUBS 0.037178f
C835 VP.n33 VSUBS 0.037178f
C836 VP.n34 VSUBS 0.037178f
C837 VP.n35 VSUBS 0.065165f
C838 VP.n36 VSUBS 0.06929f
C839 VP.n37 VSUBS 0.06929f
C840 VP.n38 VSUBS 0.037178f
C841 VP.n39 VSUBS 0.037178f
C842 VP.n40 VSUBS 0.037178f
C843 VP.n41 VSUBS 0.06929f
C844 VP.n42 VSUBS 0.06929f
C845 VP.n43 VSUBS 0.065165f
C846 VP.n44 VSUBS 0.037178f
C847 VP.n45 VSUBS 0.037178f
C848 VP.n46 VSUBS 0.037178f
C849 VP.n47 VSUBS 0.072067f
C850 VP.n48 VSUBS 0.06929f
C851 VP.n49 VSUBS 0.050133f
C852 VP.n50 VSUBS 0.060004f
C853 VP.n51 VSUBS 0.096923f
C854 VTAIL.t7 VSUBS 0.175837f
C855 VTAIL.t8 VSUBS 0.175837f
C856 VTAIL.n0 VSUBS 1.05601f
C857 VTAIL.n1 VSUBS 0.975173f
C858 VTAIL.n2 VSUBS 0.035849f
C859 VTAIL.n3 VSUBS 0.033663f
C860 VTAIL.n4 VSUBS 0.018089f
C861 VTAIL.n5 VSUBS 0.042756f
C862 VTAIL.n6 VSUBS 0.019153f
C863 VTAIL.n7 VSUBS 0.033663f
C864 VTAIL.n8 VSUBS 0.018089f
C865 VTAIL.n9 VSUBS 0.042756f
C866 VTAIL.n10 VSUBS 0.019153f
C867 VTAIL.n11 VSUBS 0.866312f
C868 VTAIL.n12 VSUBS 0.018089f
C869 VTAIL.t2 VSUBS 0.091331f
C870 VTAIL.n13 VSUBS 0.15447f
C871 VTAIL.n14 VSUBS 0.027194f
C872 VTAIL.n15 VSUBS 0.032067f
C873 VTAIL.n16 VSUBS 0.042756f
C874 VTAIL.n17 VSUBS 0.019153f
C875 VTAIL.n18 VSUBS 0.018089f
C876 VTAIL.n19 VSUBS 0.033663f
C877 VTAIL.n20 VSUBS 0.033663f
C878 VTAIL.n21 VSUBS 0.018089f
C879 VTAIL.n22 VSUBS 0.019153f
C880 VTAIL.n23 VSUBS 0.042756f
C881 VTAIL.n24 VSUBS 0.042756f
C882 VTAIL.n25 VSUBS 0.019153f
C883 VTAIL.n26 VSUBS 0.018089f
C884 VTAIL.n27 VSUBS 0.033663f
C885 VTAIL.n28 VSUBS 0.033663f
C886 VTAIL.n29 VSUBS 0.018089f
C887 VTAIL.n30 VSUBS 0.019153f
C888 VTAIL.n31 VSUBS 0.042756f
C889 VTAIL.n32 VSUBS 0.099626f
C890 VTAIL.n33 VSUBS 0.019153f
C891 VTAIL.n34 VSUBS 0.018089f
C892 VTAIL.n35 VSUBS 0.072752f
C893 VTAIL.n36 VSUBS 0.049768f
C894 VTAIL.n37 VSUBS 0.598642f
C895 VTAIL.t3 VSUBS 0.175837f
C896 VTAIL.t4 VSUBS 0.175837f
C897 VTAIL.n38 VSUBS 1.05601f
C898 VTAIL.n39 VSUBS 2.77593f
C899 VTAIL.t6 VSUBS 0.175837f
C900 VTAIL.t11 VSUBS 0.175837f
C901 VTAIL.n40 VSUBS 1.05601f
C902 VTAIL.n41 VSUBS 2.77593f
C903 VTAIL.n42 VSUBS 0.035849f
C904 VTAIL.n43 VSUBS 0.033663f
C905 VTAIL.n44 VSUBS 0.018089f
C906 VTAIL.n45 VSUBS 0.042756f
C907 VTAIL.n46 VSUBS 0.019153f
C908 VTAIL.n47 VSUBS 0.033663f
C909 VTAIL.n48 VSUBS 0.018089f
C910 VTAIL.n49 VSUBS 0.042756f
C911 VTAIL.n50 VSUBS 0.019153f
C912 VTAIL.n51 VSUBS 0.866312f
C913 VTAIL.n52 VSUBS 0.018089f
C914 VTAIL.t9 VSUBS 0.091331f
C915 VTAIL.n53 VSUBS 0.15447f
C916 VTAIL.n54 VSUBS 0.027194f
C917 VTAIL.n55 VSUBS 0.032067f
C918 VTAIL.n56 VSUBS 0.042756f
C919 VTAIL.n57 VSUBS 0.019153f
C920 VTAIL.n58 VSUBS 0.018089f
C921 VTAIL.n59 VSUBS 0.033663f
C922 VTAIL.n60 VSUBS 0.033663f
C923 VTAIL.n61 VSUBS 0.018089f
C924 VTAIL.n62 VSUBS 0.019153f
C925 VTAIL.n63 VSUBS 0.042756f
C926 VTAIL.n64 VSUBS 0.042756f
C927 VTAIL.n65 VSUBS 0.019153f
C928 VTAIL.n66 VSUBS 0.018089f
C929 VTAIL.n67 VSUBS 0.033663f
C930 VTAIL.n68 VSUBS 0.033663f
C931 VTAIL.n69 VSUBS 0.018089f
C932 VTAIL.n70 VSUBS 0.019153f
C933 VTAIL.n71 VSUBS 0.042756f
C934 VTAIL.n72 VSUBS 0.099626f
C935 VTAIL.n73 VSUBS 0.019153f
C936 VTAIL.n74 VSUBS 0.018089f
C937 VTAIL.n75 VSUBS 0.072752f
C938 VTAIL.n76 VSUBS 0.049768f
C939 VTAIL.n77 VSUBS 0.598642f
C940 VTAIL.t0 VSUBS 0.175837f
C941 VTAIL.t1 VSUBS 0.175837f
C942 VTAIL.n78 VSUBS 1.05601f
C943 VTAIL.n79 VSUBS 1.22974f
C944 VTAIL.n80 VSUBS 0.035849f
C945 VTAIL.n81 VSUBS 0.033663f
C946 VTAIL.n82 VSUBS 0.018089f
C947 VTAIL.n83 VSUBS 0.042756f
C948 VTAIL.n84 VSUBS 0.019153f
C949 VTAIL.n85 VSUBS 0.033663f
C950 VTAIL.n86 VSUBS 0.018089f
C951 VTAIL.n87 VSUBS 0.042756f
C952 VTAIL.n88 VSUBS 0.019153f
C953 VTAIL.n89 VSUBS 0.866312f
C954 VTAIL.n90 VSUBS 0.018089f
C955 VTAIL.t5 VSUBS 0.091331f
C956 VTAIL.n91 VSUBS 0.15447f
C957 VTAIL.n92 VSUBS 0.027194f
C958 VTAIL.n93 VSUBS 0.032067f
C959 VTAIL.n94 VSUBS 0.042756f
C960 VTAIL.n95 VSUBS 0.019153f
C961 VTAIL.n96 VSUBS 0.018089f
C962 VTAIL.n97 VSUBS 0.033663f
C963 VTAIL.n98 VSUBS 0.033663f
C964 VTAIL.n99 VSUBS 0.018089f
C965 VTAIL.n100 VSUBS 0.019153f
C966 VTAIL.n101 VSUBS 0.042756f
C967 VTAIL.n102 VSUBS 0.042756f
C968 VTAIL.n103 VSUBS 0.019153f
C969 VTAIL.n104 VSUBS 0.018089f
C970 VTAIL.n105 VSUBS 0.033663f
C971 VTAIL.n106 VSUBS 0.033663f
C972 VTAIL.n107 VSUBS 0.018089f
C973 VTAIL.n108 VSUBS 0.019153f
C974 VTAIL.n109 VSUBS 0.042756f
C975 VTAIL.n110 VSUBS 0.099626f
C976 VTAIL.n111 VSUBS 0.019153f
C977 VTAIL.n112 VSUBS 0.018089f
C978 VTAIL.n113 VSUBS 0.072752f
C979 VTAIL.n114 VSUBS 0.049768f
C980 VTAIL.n115 VSUBS 1.79697f
C981 VTAIL.n116 VSUBS 0.035849f
C982 VTAIL.n117 VSUBS 0.033663f
C983 VTAIL.n118 VSUBS 0.018089f
C984 VTAIL.n119 VSUBS 0.042756f
C985 VTAIL.n120 VSUBS 0.019153f
C986 VTAIL.n121 VSUBS 0.033663f
C987 VTAIL.n122 VSUBS 0.018089f
C988 VTAIL.n123 VSUBS 0.042756f
C989 VTAIL.n124 VSUBS 0.019153f
C990 VTAIL.n125 VSUBS 0.866312f
C991 VTAIL.n126 VSUBS 0.018089f
C992 VTAIL.t10 VSUBS 0.091331f
C993 VTAIL.n127 VSUBS 0.15447f
C994 VTAIL.n128 VSUBS 0.027194f
C995 VTAIL.n129 VSUBS 0.032067f
C996 VTAIL.n130 VSUBS 0.042756f
C997 VTAIL.n131 VSUBS 0.019153f
C998 VTAIL.n132 VSUBS 0.018089f
C999 VTAIL.n133 VSUBS 0.033663f
C1000 VTAIL.n134 VSUBS 0.033663f
C1001 VTAIL.n135 VSUBS 0.018089f
C1002 VTAIL.n136 VSUBS 0.019153f
C1003 VTAIL.n137 VSUBS 0.042756f
C1004 VTAIL.n138 VSUBS 0.042756f
C1005 VTAIL.n139 VSUBS 0.019153f
C1006 VTAIL.n140 VSUBS 0.018089f
C1007 VTAIL.n141 VSUBS 0.033663f
C1008 VTAIL.n142 VSUBS 0.033663f
C1009 VTAIL.n143 VSUBS 0.018089f
C1010 VTAIL.n144 VSUBS 0.019153f
C1011 VTAIL.n145 VSUBS 0.042756f
C1012 VTAIL.n146 VSUBS 0.099626f
C1013 VTAIL.n147 VSUBS 0.019153f
C1014 VTAIL.n148 VSUBS 0.018089f
C1015 VTAIL.n149 VSUBS 0.072752f
C1016 VTAIL.n150 VSUBS 0.049768f
C1017 VTAIL.n151 VSUBS 1.7037f
C1018 VDD2.n0 VSUBS 0.02836f
C1019 VDD2.n1 VSUBS 0.026631f
C1020 VDD2.n2 VSUBS 0.01431f
C1021 VDD2.n3 VSUBS 0.033824f
C1022 VDD2.n4 VSUBS 0.015152f
C1023 VDD2.n5 VSUBS 0.026631f
C1024 VDD2.n6 VSUBS 0.01431f
C1025 VDD2.n7 VSUBS 0.033824f
C1026 VDD2.n8 VSUBS 0.015152f
C1027 VDD2.n9 VSUBS 0.685334f
C1028 VDD2.n10 VSUBS 0.01431f
C1029 VDD2.t3 VSUBS 0.072251f
C1030 VDD2.n11 VSUBS 0.1222f
C1031 VDD2.n12 VSUBS 0.021513f
C1032 VDD2.n13 VSUBS 0.025368f
C1033 VDD2.n14 VSUBS 0.033824f
C1034 VDD2.n15 VSUBS 0.015152f
C1035 VDD2.n16 VSUBS 0.01431f
C1036 VDD2.n17 VSUBS 0.026631f
C1037 VDD2.n18 VSUBS 0.026631f
C1038 VDD2.n19 VSUBS 0.01431f
C1039 VDD2.n20 VSUBS 0.015152f
C1040 VDD2.n21 VSUBS 0.033824f
C1041 VDD2.n22 VSUBS 0.033824f
C1042 VDD2.n23 VSUBS 0.015152f
C1043 VDD2.n24 VSUBS 0.01431f
C1044 VDD2.n25 VSUBS 0.026631f
C1045 VDD2.n26 VSUBS 0.026631f
C1046 VDD2.n27 VSUBS 0.01431f
C1047 VDD2.n28 VSUBS 0.015152f
C1048 VDD2.n29 VSUBS 0.033824f
C1049 VDD2.n30 VSUBS 0.078813f
C1050 VDD2.n31 VSUBS 0.015152f
C1051 VDD2.n32 VSUBS 0.01431f
C1052 VDD2.n33 VSUBS 0.057554f
C1053 VDD2.n34 VSUBS 0.069806f
C1054 VDD2.t5 VSUBS 0.139103f
C1055 VDD2.t0 VSUBS 0.139103f
C1056 VDD2.n35 VSUBS 0.948774f
C1057 VDD2.n36 VSUBS 3.09219f
C1058 VDD2.n37 VSUBS 0.02836f
C1059 VDD2.n38 VSUBS 0.026631f
C1060 VDD2.n39 VSUBS 0.01431f
C1061 VDD2.n40 VSUBS 0.033824f
C1062 VDD2.n41 VSUBS 0.015152f
C1063 VDD2.n42 VSUBS 0.026631f
C1064 VDD2.n43 VSUBS 0.01431f
C1065 VDD2.n44 VSUBS 0.033824f
C1066 VDD2.n45 VSUBS 0.015152f
C1067 VDD2.n46 VSUBS 0.685334f
C1068 VDD2.n47 VSUBS 0.01431f
C1069 VDD2.t1 VSUBS 0.072251f
C1070 VDD2.n48 VSUBS 0.1222f
C1071 VDD2.n49 VSUBS 0.021513f
C1072 VDD2.n50 VSUBS 0.025368f
C1073 VDD2.n51 VSUBS 0.033824f
C1074 VDD2.n52 VSUBS 0.015152f
C1075 VDD2.n53 VSUBS 0.01431f
C1076 VDD2.n54 VSUBS 0.026631f
C1077 VDD2.n55 VSUBS 0.026631f
C1078 VDD2.n56 VSUBS 0.01431f
C1079 VDD2.n57 VSUBS 0.015152f
C1080 VDD2.n58 VSUBS 0.033824f
C1081 VDD2.n59 VSUBS 0.033824f
C1082 VDD2.n60 VSUBS 0.015152f
C1083 VDD2.n61 VSUBS 0.01431f
C1084 VDD2.n62 VSUBS 0.026631f
C1085 VDD2.n63 VSUBS 0.026631f
C1086 VDD2.n64 VSUBS 0.01431f
C1087 VDD2.n65 VSUBS 0.015152f
C1088 VDD2.n66 VSUBS 0.033824f
C1089 VDD2.n67 VSUBS 0.078813f
C1090 VDD2.n68 VSUBS 0.015152f
C1091 VDD2.n69 VSUBS 0.01431f
C1092 VDD2.n70 VSUBS 0.057554f
C1093 VDD2.n71 VSUBS 0.057794f
C1094 VDD2.n72 VSUBS 2.50944f
C1095 VDD2.t4 VSUBS 0.139103f
C1096 VDD2.t2 VSUBS 0.139103f
C1097 VDD2.n73 VSUBS 0.948739f
C1098 VN.t1 VSUBS 1.96667f
C1099 VN.n0 VSUBS 0.845739f
C1100 VN.n1 VSUBS 0.032981f
C1101 VN.n2 VSUBS 0.036019f
C1102 VN.n3 VSUBS 0.032981f
C1103 VN.t3 VSUBS 1.96667f
C1104 VN.n4 VSUBS 0.850824f
C1105 VN.t4 VSUBS 2.36831f
C1106 VN.n5 VSUBS 0.797616f
C1107 VN.n6 VSUBS 0.402663f
C1108 VN.n7 VSUBS 0.061468f
C1109 VN.n8 VSUBS 0.061468f
C1110 VN.n9 VSUBS 0.057809f
C1111 VN.n10 VSUBS 0.032981f
C1112 VN.n11 VSUBS 0.032981f
C1113 VN.n12 VSUBS 0.032981f
C1114 VN.n13 VSUBS 0.063932f
C1115 VN.n14 VSUBS 0.061468f
C1116 VN.n15 VSUBS 0.044474f
C1117 VN.n16 VSUBS 0.05323f
C1118 VN.n17 VSUBS 0.085982f
C1119 VN.t5 VSUBS 1.96667f
C1120 VN.n18 VSUBS 0.845739f
C1121 VN.n19 VSUBS 0.032981f
C1122 VN.n20 VSUBS 0.036019f
C1123 VN.n21 VSUBS 0.032981f
C1124 VN.t0 VSUBS 1.96667f
C1125 VN.n22 VSUBS 0.850824f
C1126 VN.t2 VSUBS 2.36831f
C1127 VN.n23 VSUBS 0.797616f
C1128 VN.n24 VSUBS 0.402663f
C1129 VN.n25 VSUBS 0.061468f
C1130 VN.n26 VSUBS 0.061468f
C1131 VN.n27 VSUBS 0.057809f
C1132 VN.n28 VSUBS 0.032981f
C1133 VN.n29 VSUBS 0.032981f
C1134 VN.n30 VSUBS 0.032981f
C1135 VN.n31 VSUBS 0.063932f
C1136 VN.n32 VSUBS 0.061468f
C1137 VN.n33 VSUBS 0.044474f
C1138 VN.n34 VSUBS 0.05323f
C1139 VN.n35 VSUBS 1.77486f
.ends

