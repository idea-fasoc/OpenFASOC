* NGSPICE file created from diff_pair_sample_1378.ext - technology: sky130A

.subckt diff_pair_sample_1378 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.0085 pd=11.08 as=2.0085 ps=11.08 w=5.15 l=2.03
X1 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.0085 pd=11.08 as=2.0085 ps=11.08 w=5.15 l=2.03
X2 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=2.0085 pd=11.08 as=0 ps=0 w=5.15 l=2.03
X3 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=2.0085 pd=11.08 as=0 ps=0 w=5.15 l=2.03
X4 VDD2.t0 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.0085 pd=11.08 as=2.0085 ps=11.08 w=5.15 l=2.03
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.0085 pd=11.08 as=0 ps=0 w=5.15 l=2.03
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.0085 pd=11.08 as=0 ps=0 w=5.15 l=2.03
X7 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.0085 pd=11.08 as=2.0085 ps=11.08 w=5.15 l=2.03
R0 VN VN.t1 158.149
R1 VN VN.t0 120.243
R2 VTAIL.n102 VTAIL.n101 289.615
R3 VTAIL.n24 VTAIL.n23 289.615
R4 VTAIL.n76 VTAIL.n75 289.615
R5 VTAIL.n50 VTAIL.n49 289.615
R6 VTAIL.n87 VTAIL.n86 185
R7 VTAIL.n84 VTAIL.n83 185
R8 VTAIL.n93 VTAIL.n92 185
R9 VTAIL.n95 VTAIL.n94 185
R10 VTAIL.n80 VTAIL.n79 185
R11 VTAIL.n101 VTAIL.n100 185
R12 VTAIL.n9 VTAIL.n8 185
R13 VTAIL.n6 VTAIL.n5 185
R14 VTAIL.n15 VTAIL.n14 185
R15 VTAIL.n17 VTAIL.n16 185
R16 VTAIL.n2 VTAIL.n1 185
R17 VTAIL.n23 VTAIL.n22 185
R18 VTAIL.n75 VTAIL.n74 185
R19 VTAIL.n54 VTAIL.n53 185
R20 VTAIL.n69 VTAIL.n68 185
R21 VTAIL.n67 VTAIL.n66 185
R22 VTAIL.n58 VTAIL.n57 185
R23 VTAIL.n61 VTAIL.n60 185
R24 VTAIL.n49 VTAIL.n48 185
R25 VTAIL.n28 VTAIL.n27 185
R26 VTAIL.n43 VTAIL.n42 185
R27 VTAIL.n41 VTAIL.n40 185
R28 VTAIL.n32 VTAIL.n31 185
R29 VTAIL.n35 VTAIL.n34 185
R30 VTAIL.t2 VTAIL.n85 149.54
R31 VTAIL.t1 VTAIL.n7 149.54
R32 VTAIL.t3 VTAIL.n33 149.54
R33 VTAIL.t0 VTAIL.n59 149.54
R34 VTAIL.n86 VTAIL.n83 104.615
R35 VTAIL.n93 VTAIL.n83 104.615
R36 VTAIL.n94 VTAIL.n93 104.615
R37 VTAIL.n94 VTAIL.n79 104.615
R38 VTAIL.n101 VTAIL.n79 104.615
R39 VTAIL.n8 VTAIL.n5 104.615
R40 VTAIL.n15 VTAIL.n5 104.615
R41 VTAIL.n16 VTAIL.n15 104.615
R42 VTAIL.n16 VTAIL.n1 104.615
R43 VTAIL.n23 VTAIL.n1 104.615
R44 VTAIL.n75 VTAIL.n53 104.615
R45 VTAIL.n68 VTAIL.n53 104.615
R46 VTAIL.n68 VTAIL.n67 104.615
R47 VTAIL.n67 VTAIL.n57 104.615
R48 VTAIL.n60 VTAIL.n57 104.615
R49 VTAIL.n49 VTAIL.n27 104.615
R50 VTAIL.n42 VTAIL.n27 104.615
R51 VTAIL.n42 VTAIL.n41 104.615
R52 VTAIL.n41 VTAIL.n31 104.615
R53 VTAIL.n34 VTAIL.n31 104.615
R54 VTAIL.n86 VTAIL.t2 52.3082
R55 VTAIL.n8 VTAIL.t1 52.3082
R56 VTAIL.n60 VTAIL.t0 52.3082
R57 VTAIL.n34 VTAIL.t3 52.3082
R58 VTAIL.n103 VTAIL.n102 34.7066
R59 VTAIL.n25 VTAIL.n24 34.7066
R60 VTAIL.n77 VTAIL.n76 34.7066
R61 VTAIL.n51 VTAIL.n50 34.7066
R62 VTAIL.n51 VTAIL.n25 20.8755
R63 VTAIL.n103 VTAIL.n77 18.841
R64 VTAIL.n100 VTAIL.n78 11.249
R65 VTAIL.n22 VTAIL.n0 11.249
R66 VTAIL.n74 VTAIL.n52 11.249
R67 VTAIL.n48 VTAIL.n26 11.249
R68 VTAIL.n99 VTAIL.n80 10.4732
R69 VTAIL.n21 VTAIL.n2 10.4732
R70 VTAIL.n73 VTAIL.n54 10.4732
R71 VTAIL.n47 VTAIL.n28 10.4732
R72 VTAIL.n87 VTAIL.n85 10.2739
R73 VTAIL.n9 VTAIL.n7 10.2739
R74 VTAIL.n61 VTAIL.n59 10.2739
R75 VTAIL.n35 VTAIL.n33 10.2739
R76 VTAIL.n96 VTAIL.n95 9.69747
R77 VTAIL.n18 VTAIL.n17 9.69747
R78 VTAIL.n70 VTAIL.n69 9.69747
R79 VTAIL.n44 VTAIL.n43 9.69747
R80 VTAIL.n98 VTAIL.n78 9.45567
R81 VTAIL.n20 VTAIL.n0 9.45567
R82 VTAIL.n72 VTAIL.n52 9.45567
R83 VTAIL.n46 VTAIL.n26 9.45567
R84 VTAIL.n89 VTAIL.n88 9.3005
R85 VTAIL.n91 VTAIL.n90 9.3005
R86 VTAIL.n82 VTAIL.n81 9.3005
R87 VTAIL.n97 VTAIL.n96 9.3005
R88 VTAIL.n99 VTAIL.n98 9.3005
R89 VTAIL.n11 VTAIL.n10 9.3005
R90 VTAIL.n13 VTAIL.n12 9.3005
R91 VTAIL.n4 VTAIL.n3 9.3005
R92 VTAIL.n19 VTAIL.n18 9.3005
R93 VTAIL.n21 VTAIL.n20 9.3005
R94 VTAIL.n73 VTAIL.n72 9.3005
R95 VTAIL.n71 VTAIL.n70 9.3005
R96 VTAIL.n56 VTAIL.n55 9.3005
R97 VTAIL.n65 VTAIL.n64 9.3005
R98 VTAIL.n63 VTAIL.n62 9.3005
R99 VTAIL.n39 VTAIL.n38 9.3005
R100 VTAIL.n30 VTAIL.n29 9.3005
R101 VTAIL.n45 VTAIL.n44 9.3005
R102 VTAIL.n47 VTAIL.n46 9.3005
R103 VTAIL.n37 VTAIL.n36 9.3005
R104 VTAIL.n92 VTAIL.n82 8.92171
R105 VTAIL.n14 VTAIL.n4 8.92171
R106 VTAIL.n66 VTAIL.n56 8.92171
R107 VTAIL.n40 VTAIL.n30 8.92171
R108 VTAIL.n91 VTAIL.n84 8.14595
R109 VTAIL.n13 VTAIL.n6 8.14595
R110 VTAIL.n65 VTAIL.n58 8.14595
R111 VTAIL.n39 VTAIL.n32 8.14595
R112 VTAIL.n88 VTAIL.n87 7.3702
R113 VTAIL.n10 VTAIL.n9 7.3702
R114 VTAIL.n62 VTAIL.n61 7.3702
R115 VTAIL.n36 VTAIL.n35 7.3702
R116 VTAIL.n88 VTAIL.n84 5.81868
R117 VTAIL.n10 VTAIL.n6 5.81868
R118 VTAIL.n62 VTAIL.n58 5.81868
R119 VTAIL.n36 VTAIL.n32 5.81868
R120 VTAIL.n92 VTAIL.n91 5.04292
R121 VTAIL.n14 VTAIL.n13 5.04292
R122 VTAIL.n66 VTAIL.n65 5.04292
R123 VTAIL.n40 VTAIL.n39 5.04292
R124 VTAIL.n95 VTAIL.n82 4.26717
R125 VTAIL.n17 VTAIL.n4 4.26717
R126 VTAIL.n69 VTAIL.n56 4.26717
R127 VTAIL.n43 VTAIL.n30 4.26717
R128 VTAIL.n96 VTAIL.n80 3.49141
R129 VTAIL.n18 VTAIL.n2 3.49141
R130 VTAIL.n70 VTAIL.n54 3.49141
R131 VTAIL.n44 VTAIL.n28 3.49141
R132 VTAIL.n89 VTAIL.n85 2.84386
R133 VTAIL.n11 VTAIL.n7 2.84386
R134 VTAIL.n37 VTAIL.n33 2.84386
R135 VTAIL.n63 VTAIL.n59 2.84386
R136 VTAIL.n100 VTAIL.n99 2.71565
R137 VTAIL.n22 VTAIL.n21 2.71565
R138 VTAIL.n74 VTAIL.n73 2.71565
R139 VTAIL.n48 VTAIL.n47 2.71565
R140 VTAIL.n102 VTAIL.n78 1.93989
R141 VTAIL.n24 VTAIL.n0 1.93989
R142 VTAIL.n76 VTAIL.n52 1.93989
R143 VTAIL.n50 VTAIL.n26 1.93989
R144 VTAIL.n77 VTAIL.n51 1.48757
R145 VTAIL VTAIL.n25 1.03714
R146 VTAIL VTAIL.n103 0.450931
R147 VTAIL.n90 VTAIL.n89 0.155672
R148 VTAIL.n90 VTAIL.n81 0.155672
R149 VTAIL.n97 VTAIL.n81 0.155672
R150 VTAIL.n98 VTAIL.n97 0.155672
R151 VTAIL.n12 VTAIL.n11 0.155672
R152 VTAIL.n12 VTAIL.n3 0.155672
R153 VTAIL.n19 VTAIL.n3 0.155672
R154 VTAIL.n20 VTAIL.n19 0.155672
R155 VTAIL.n72 VTAIL.n71 0.155672
R156 VTAIL.n71 VTAIL.n55 0.155672
R157 VTAIL.n64 VTAIL.n55 0.155672
R158 VTAIL.n64 VTAIL.n63 0.155672
R159 VTAIL.n46 VTAIL.n45 0.155672
R160 VTAIL.n45 VTAIL.n29 0.155672
R161 VTAIL.n38 VTAIL.n29 0.155672
R162 VTAIL.n38 VTAIL.n37 0.155672
R163 VDD2.n49 VDD2.n48 289.615
R164 VDD2.n24 VDD2.n23 289.615
R165 VDD2.n48 VDD2.n47 185
R166 VDD2.n27 VDD2.n26 185
R167 VDD2.n42 VDD2.n41 185
R168 VDD2.n40 VDD2.n39 185
R169 VDD2.n31 VDD2.n30 185
R170 VDD2.n34 VDD2.n33 185
R171 VDD2.n9 VDD2.n8 185
R172 VDD2.n6 VDD2.n5 185
R173 VDD2.n15 VDD2.n14 185
R174 VDD2.n17 VDD2.n16 185
R175 VDD2.n2 VDD2.n1 185
R176 VDD2.n23 VDD2.n22 185
R177 VDD2.t1 VDD2.n7 149.54
R178 VDD2.t0 VDD2.n32 149.54
R179 VDD2.n48 VDD2.n26 104.615
R180 VDD2.n41 VDD2.n26 104.615
R181 VDD2.n41 VDD2.n40 104.615
R182 VDD2.n40 VDD2.n30 104.615
R183 VDD2.n33 VDD2.n30 104.615
R184 VDD2.n8 VDD2.n5 104.615
R185 VDD2.n15 VDD2.n5 104.615
R186 VDD2.n16 VDD2.n15 104.615
R187 VDD2.n16 VDD2.n1 104.615
R188 VDD2.n23 VDD2.n1 104.615
R189 VDD2.n50 VDD2.n24 83.5534
R190 VDD2.n33 VDD2.t0 52.3082
R191 VDD2.n8 VDD2.t1 52.3082
R192 VDD2.n50 VDD2.n49 51.3853
R193 VDD2.n47 VDD2.n25 11.249
R194 VDD2.n22 VDD2.n0 11.249
R195 VDD2.n46 VDD2.n27 10.4732
R196 VDD2.n21 VDD2.n2 10.4732
R197 VDD2.n34 VDD2.n32 10.2739
R198 VDD2.n9 VDD2.n7 10.2739
R199 VDD2.n43 VDD2.n42 9.69747
R200 VDD2.n18 VDD2.n17 9.69747
R201 VDD2.n45 VDD2.n25 9.45567
R202 VDD2.n20 VDD2.n0 9.45567
R203 VDD2.n46 VDD2.n45 9.3005
R204 VDD2.n44 VDD2.n43 9.3005
R205 VDD2.n29 VDD2.n28 9.3005
R206 VDD2.n38 VDD2.n37 9.3005
R207 VDD2.n36 VDD2.n35 9.3005
R208 VDD2.n11 VDD2.n10 9.3005
R209 VDD2.n13 VDD2.n12 9.3005
R210 VDD2.n4 VDD2.n3 9.3005
R211 VDD2.n19 VDD2.n18 9.3005
R212 VDD2.n21 VDD2.n20 9.3005
R213 VDD2.n39 VDD2.n29 8.92171
R214 VDD2.n14 VDD2.n4 8.92171
R215 VDD2.n38 VDD2.n31 8.14595
R216 VDD2.n13 VDD2.n6 8.14595
R217 VDD2.n35 VDD2.n34 7.3702
R218 VDD2.n10 VDD2.n9 7.3702
R219 VDD2.n35 VDD2.n31 5.81868
R220 VDD2.n10 VDD2.n6 5.81868
R221 VDD2.n39 VDD2.n38 5.04292
R222 VDD2.n14 VDD2.n13 5.04292
R223 VDD2.n42 VDD2.n29 4.26717
R224 VDD2.n17 VDD2.n4 4.26717
R225 VDD2.n43 VDD2.n27 3.49141
R226 VDD2.n18 VDD2.n2 3.49141
R227 VDD2.n11 VDD2.n7 2.84386
R228 VDD2.n36 VDD2.n32 2.84386
R229 VDD2.n47 VDD2.n46 2.71565
R230 VDD2.n22 VDD2.n21 2.71565
R231 VDD2.n49 VDD2.n25 1.93989
R232 VDD2.n24 VDD2.n0 1.93989
R233 VDD2 VDD2.n50 0.56731
R234 VDD2.n45 VDD2.n44 0.155672
R235 VDD2.n44 VDD2.n28 0.155672
R236 VDD2.n37 VDD2.n28 0.155672
R237 VDD2.n37 VDD2.n36 0.155672
R238 VDD2.n12 VDD2.n11 0.155672
R239 VDD2.n12 VDD2.n3 0.155672
R240 VDD2.n19 VDD2.n3 0.155672
R241 VDD2.n20 VDD2.n19 0.155672
R242 B.n347 B.n346 585
R243 B.n349 B.n74 585
R244 B.n352 B.n351 585
R245 B.n353 B.n73 585
R246 B.n355 B.n354 585
R247 B.n357 B.n72 585
R248 B.n360 B.n359 585
R249 B.n361 B.n71 585
R250 B.n363 B.n362 585
R251 B.n365 B.n70 585
R252 B.n368 B.n367 585
R253 B.n369 B.n69 585
R254 B.n371 B.n370 585
R255 B.n373 B.n68 585
R256 B.n376 B.n375 585
R257 B.n377 B.n67 585
R258 B.n379 B.n378 585
R259 B.n381 B.n66 585
R260 B.n384 B.n383 585
R261 B.n385 B.n62 585
R262 B.n387 B.n386 585
R263 B.n389 B.n61 585
R264 B.n392 B.n391 585
R265 B.n393 B.n60 585
R266 B.n395 B.n394 585
R267 B.n397 B.n59 585
R268 B.n400 B.n399 585
R269 B.n401 B.n58 585
R270 B.n403 B.n402 585
R271 B.n405 B.n57 585
R272 B.n408 B.n407 585
R273 B.n410 B.n54 585
R274 B.n412 B.n411 585
R275 B.n414 B.n53 585
R276 B.n417 B.n416 585
R277 B.n418 B.n52 585
R278 B.n420 B.n419 585
R279 B.n422 B.n51 585
R280 B.n425 B.n424 585
R281 B.n426 B.n50 585
R282 B.n428 B.n427 585
R283 B.n430 B.n49 585
R284 B.n433 B.n432 585
R285 B.n434 B.n48 585
R286 B.n436 B.n435 585
R287 B.n438 B.n47 585
R288 B.n441 B.n440 585
R289 B.n442 B.n46 585
R290 B.n444 B.n443 585
R291 B.n446 B.n45 585
R292 B.n449 B.n448 585
R293 B.n450 B.n44 585
R294 B.n345 B.n42 585
R295 B.n453 B.n42 585
R296 B.n344 B.n41 585
R297 B.n454 B.n41 585
R298 B.n343 B.n40 585
R299 B.n455 B.n40 585
R300 B.n342 B.n341 585
R301 B.n341 B.n36 585
R302 B.n340 B.n35 585
R303 B.n461 B.n35 585
R304 B.n339 B.n34 585
R305 B.n462 B.n34 585
R306 B.n338 B.n33 585
R307 B.n463 B.n33 585
R308 B.n337 B.n336 585
R309 B.n336 B.n29 585
R310 B.n335 B.n28 585
R311 B.n469 B.n28 585
R312 B.n334 B.n27 585
R313 B.n470 B.n27 585
R314 B.n333 B.n26 585
R315 B.n471 B.n26 585
R316 B.n332 B.n331 585
R317 B.n331 B.n22 585
R318 B.n330 B.n21 585
R319 B.n477 B.n21 585
R320 B.n329 B.n20 585
R321 B.n478 B.n20 585
R322 B.n328 B.n19 585
R323 B.n479 B.n19 585
R324 B.n327 B.n326 585
R325 B.n326 B.n15 585
R326 B.n325 B.n14 585
R327 B.n485 B.n14 585
R328 B.n324 B.n13 585
R329 B.n486 B.n13 585
R330 B.n323 B.n12 585
R331 B.n487 B.n12 585
R332 B.n322 B.n321 585
R333 B.n321 B.n8 585
R334 B.n320 B.n7 585
R335 B.n493 B.n7 585
R336 B.n319 B.n6 585
R337 B.n494 B.n6 585
R338 B.n318 B.n5 585
R339 B.n495 B.n5 585
R340 B.n317 B.n316 585
R341 B.n316 B.n4 585
R342 B.n315 B.n75 585
R343 B.n315 B.n314 585
R344 B.n305 B.n76 585
R345 B.n77 B.n76 585
R346 B.n307 B.n306 585
R347 B.n308 B.n307 585
R348 B.n304 B.n82 585
R349 B.n82 B.n81 585
R350 B.n303 B.n302 585
R351 B.n302 B.n301 585
R352 B.n84 B.n83 585
R353 B.n85 B.n84 585
R354 B.n294 B.n293 585
R355 B.n295 B.n294 585
R356 B.n292 B.n90 585
R357 B.n90 B.n89 585
R358 B.n291 B.n290 585
R359 B.n290 B.n289 585
R360 B.n92 B.n91 585
R361 B.n93 B.n92 585
R362 B.n282 B.n281 585
R363 B.n283 B.n282 585
R364 B.n280 B.n98 585
R365 B.n98 B.n97 585
R366 B.n279 B.n278 585
R367 B.n278 B.n277 585
R368 B.n100 B.n99 585
R369 B.n101 B.n100 585
R370 B.n270 B.n269 585
R371 B.n271 B.n270 585
R372 B.n268 B.n106 585
R373 B.n106 B.n105 585
R374 B.n267 B.n266 585
R375 B.n266 B.n265 585
R376 B.n108 B.n107 585
R377 B.n109 B.n108 585
R378 B.n258 B.n257 585
R379 B.n259 B.n258 585
R380 B.n256 B.n114 585
R381 B.n114 B.n113 585
R382 B.n255 B.n254 585
R383 B.n254 B.n253 585
R384 B.n250 B.n118 585
R385 B.n249 B.n248 585
R386 B.n246 B.n119 585
R387 B.n246 B.n117 585
R388 B.n245 B.n244 585
R389 B.n243 B.n242 585
R390 B.n241 B.n121 585
R391 B.n239 B.n238 585
R392 B.n237 B.n122 585
R393 B.n236 B.n235 585
R394 B.n233 B.n123 585
R395 B.n231 B.n230 585
R396 B.n229 B.n124 585
R397 B.n228 B.n227 585
R398 B.n225 B.n125 585
R399 B.n223 B.n222 585
R400 B.n221 B.n126 585
R401 B.n220 B.n219 585
R402 B.n217 B.n127 585
R403 B.n215 B.n214 585
R404 B.n213 B.n128 585
R405 B.n212 B.n211 585
R406 B.n209 B.n208 585
R407 B.n207 B.n206 585
R408 B.n205 B.n133 585
R409 B.n203 B.n202 585
R410 B.n201 B.n134 585
R411 B.n200 B.n199 585
R412 B.n197 B.n135 585
R413 B.n195 B.n194 585
R414 B.n193 B.n136 585
R415 B.n192 B.n191 585
R416 B.n189 B.n188 585
R417 B.n187 B.n186 585
R418 B.n185 B.n141 585
R419 B.n183 B.n182 585
R420 B.n181 B.n142 585
R421 B.n180 B.n179 585
R422 B.n177 B.n143 585
R423 B.n175 B.n174 585
R424 B.n173 B.n144 585
R425 B.n172 B.n171 585
R426 B.n169 B.n145 585
R427 B.n167 B.n166 585
R428 B.n165 B.n146 585
R429 B.n164 B.n163 585
R430 B.n161 B.n147 585
R431 B.n159 B.n158 585
R432 B.n157 B.n148 585
R433 B.n156 B.n155 585
R434 B.n153 B.n149 585
R435 B.n151 B.n150 585
R436 B.n116 B.n115 585
R437 B.n117 B.n116 585
R438 B.n252 B.n251 585
R439 B.n253 B.n252 585
R440 B.n112 B.n111 585
R441 B.n113 B.n112 585
R442 B.n261 B.n260 585
R443 B.n260 B.n259 585
R444 B.n262 B.n110 585
R445 B.n110 B.n109 585
R446 B.n264 B.n263 585
R447 B.n265 B.n264 585
R448 B.n104 B.n103 585
R449 B.n105 B.n104 585
R450 B.n273 B.n272 585
R451 B.n272 B.n271 585
R452 B.n274 B.n102 585
R453 B.n102 B.n101 585
R454 B.n276 B.n275 585
R455 B.n277 B.n276 585
R456 B.n96 B.n95 585
R457 B.n97 B.n96 585
R458 B.n285 B.n284 585
R459 B.n284 B.n283 585
R460 B.n286 B.n94 585
R461 B.n94 B.n93 585
R462 B.n288 B.n287 585
R463 B.n289 B.n288 585
R464 B.n88 B.n87 585
R465 B.n89 B.n88 585
R466 B.n297 B.n296 585
R467 B.n296 B.n295 585
R468 B.n298 B.n86 585
R469 B.n86 B.n85 585
R470 B.n300 B.n299 585
R471 B.n301 B.n300 585
R472 B.n80 B.n79 585
R473 B.n81 B.n80 585
R474 B.n310 B.n309 585
R475 B.n309 B.n308 585
R476 B.n311 B.n78 585
R477 B.n78 B.n77 585
R478 B.n313 B.n312 585
R479 B.n314 B.n313 585
R480 B.n2 B.n0 585
R481 B.n4 B.n2 585
R482 B.n3 B.n1 585
R483 B.n494 B.n3 585
R484 B.n492 B.n491 585
R485 B.n493 B.n492 585
R486 B.n490 B.n9 585
R487 B.n9 B.n8 585
R488 B.n489 B.n488 585
R489 B.n488 B.n487 585
R490 B.n11 B.n10 585
R491 B.n486 B.n11 585
R492 B.n484 B.n483 585
R493 B.n485 B.n484 585
R494 B.n482 B.n16 585
R495 B.n16 B.n15 585
R496 B.n481 B.n480 585
R497 B.n480 B.n479 585
R498 B.n18 B.n17 585
R499 B.n478 B.n18 585
R500 B.n476 B.n475 585
R501 B.n477 B.n476 585
R502 B.n474 B.n23 585
R503 B.n23 B.n22 585
R504 B.n473 B.n472 585
R505 B.n472 B.n471 585
R506 B.n25 B.n24 585
R507 B.n470 B.n25 585
R508 B.n468 B.n467 585
R509 B.n469 B.n468 585
R510 B.n466 B.n30 585
R511 B.n30 B.n29 585
R512 B.n465 B.n464 585
R513 B.n464 B.n463 585
R514 B.n32 B.n31 585
R515 B.n462 B.n32 585
R516 B.n460 B.n459 585
R517 B.n461 B.n460 585
R518 B.n458 B.n37 585
R519 B.n37 B.n36 585
R520 B.n457 B.n456 585
R521 B.n456 B.n455 585
R522 B.n39 B.n38 585
R523 B.n454 B.n39 585
R524 B.n452 B.n451 585
R525 B.n453 B.n452 585
R526 B.n497 B.n496 585
R527 B.n496 B.n495 585
R528 B.n252 B.n118 540.549
R529 B.n452 B.n44 540.549
R530 B.n254 B.n116 540.549
R531 B.n347 B.n42 540.549
R532 B.n137 B.t10 268.127
R533 B.n129 B.t2 268.127
R534 B.n55 B.t13 268.127
R535 B.n63 B.t6 268.127
R536 B.n348 B.n43 256.663
R537 B.n350 B.n43 256.663
R538 B.n356 B.n43 256.663
R539 B.n358 B.n43 256.663
R540 B.n364 B.n43 256.663
R541 B.n366 B.n43 256.663
R542 B.n372 B.n43 256.663
R543 B.n374 B.n43 256.663
R544 B.n380 B.n43 256.663
R545 B.n382 B.n43 256.663
R546 B.n388 B.n43 256.663
R547 B.n390 B.n43 256.663
R548 B.n396 B.n43 256.663
R549 B.n398 B.n43 256.663
R550 B.n404 B.n43 256.663
R551 B.n406 B.n43 256.663
R552 B.n413 B.n43 256.663
R553 B.n415 B.n43 256.663
R554 B.n421 B.n43 256.663
R555 B.n423 B.n43 256.663
R556 B.n429 B.n43 256.663
R557 B.n431 B.n43 256.663
R558 B.n437 B.n43 256.663
R559 B.n439 B.n43 256.663
R560 B.n445 B.n43 256.663
R561 B.n447 B.n43 256.663
R562 B.n247 B.n117 256.663
R563 B.n120 B.n117 256.663
R564 B.n240 B.n117 256.663
R565 B.n234 B.n117 256.663
R566 B.n232 B.n117 256.663
R567 B.n226 B.n117 256.663
R568 B.n224 B.n117 256.663
R569 B.n218 B.n117 256.663
R570 B.n216 B.n117 256.663
R571 B.n210 B.n117 256.663
R572 B.n132 B.n117 256.663
R573 B.n204 B.n117 256.663
R574 B.n198 B.n117 256.663
R575 B.n196 B.n117 256.663
R576 B.n190 B.n117 256.663
R577 B.n140 B.n117 256.663
R578 B.n184 B.n117 256.663
R579 B.n178 B.n117 256.663
R580 B.n176 B.n117 256.663
R581 B.n170 B.n117 256.663
R582 B.n168 B.n117 256.663
R583 B.n162 B.n117 256.663
R584 B.n160 B.n117 256.663
R585 B.n154 B.n117 256.663
R586 B.n152 B.n117 256.663
R587 B.n137 B.t12 209.822
R588 B.n63 B.t8 209.822
R589 B.n129 B.t5 209.822
R590 B.n55 B.t14 209.822
R591 B.n138 B.t11 164.053
R592 B.n64 B.t9 164.053
R593 B.n130 B.t4 164.053
R594 B.n56 B.t15 164.053
R595 B.n252 B.n112 163.367
R596 B.n260 B.n112 163.367
R597 B.n260 B.n110 163.367
R598 B.n264 B.n110 163.367
R599 B.n264 B.n104 163.367
R600 B.n272 B.n104 163.367
R601 B.n272 B.n102 163.367
R602 B.n276 B.n102 163.367
R603 B.n276 B.n96 163.367
R604 B.n284 B.n96 163.367
R605 B.n284 B.n94 163.367
R606 B.n288 B.n94 163.367
R607 B.n288 B.n88 163.367
R608 B.n296 B.n88 163.367
R609 B.n296 B.n86 163.367
R610 B.n300 B.n86 163.367
R611 B.n300 B.n80 163.367
R612 B.n309 B.n80 163.367
R613 B.n309 B.n78 163.367
R614 B.n313 B.n78 163.367
R615 B.n313 B.n2 163.367
R616 B.n496 B.n2 163.367
R617 B.n496 B.n3 163.367
R618 B.n492 B.n3 163.367
R619 B.n492 B.n9 163.367
R620 B.n488 B.n9 163.367
R621 B.n488 B.n11 163.367
R622 B.n484 B.n11 163.367
R623 B.n484 B.n16 163.367
R624 B.n480 B.n16 163.367
R625 B.n480 B.n18 163.367
R626 B.n476 B.n18 163.367
R627 B.n476 B.n23 163.367
R628 B.n472 B.n23 163.367
R629 B.n472 B.n25 163.367
R630 B.n468 B.n25 163.367
R631 B.n468 B.n30 163.367
R632 B.n464 B.n30 163.367
R633 B.n464 B.n32 163.367
R634 B.n460 B.n32 163.367
R635 B.n460 B.n37 163.367
R636 B.n456 B.n37 163.367
R637 B.n456 B.n39 163.367
R638 B.n452 B.n39 163.367
R639 B.n248 B.n246 163.367
R640 B.n246 B.n245 163.367
R641 B.n242 B.n241 163.367
R642 B.n239 B.n122 163.367
R643 B.n235 B.n233 163.367
R644 B.n231 B.n124 163.367
R645 B.n227 B.n225 163.367
R646 B.n223 B.n126 163.367
R647 B.n219 B.n217 163.367
R648 B.n215 B.n128 163.367
R649 B.n211 B.n209 163.367
R650 B.n206 B.n205 163.367
R651 B.n203 B.n134 163.367
R652 B.n199 B.n197 163.367
R653 B.n195 B.n136 163.367
R654 B.n191 B.n189 163.367
R655 B.n186 B.n185 163.367
R656 B.n183 B.n142 163.367
R657 B.n179 B.n177 163.367
R658 B.n175 B.n144 163.367
R659 B.n171 B.n169 163.367
R660 B.n167 B.n146 163.367
R661 B.n163 B.n161 163.367
R662 B.n159 B.n148 163.367
R663 B.n155 B.n153 163.367
R664 B.n151 B.n116 163.367
R665 B.n254 B.n114 163.367
R666 B.n258 B.n114 163.367
R667 B.n258 B.n108 163.367
R668 B.n266 B.n108 163.367
R669 B.n266 B.n106 163.367
R670 B.n270 B.n106 163.367
R671 B.n270 B.n100 163.367
R672 B.n278 B.n100 163.367
R673 B.n278 B.n98 163.367
R674 B.n282 B.n98 163.367
R675 B.n282 B.n92 163.367
R676 B.n290 B.n92 163.367
R677 B.n290 B.n90 163.367
R678 B.n294 B.n90 163.367
R679 B.n294 B.n84 163.367
R680 B.n302 B.n84 163.367
R681 B.n302 B.n82 163.367
R682 B.n307 B.n82 163.367
R683 B.n307 B.n76 163.367
R684 B.n315 B.n76 163.367
R685 B.n316 B.n315 163.367
R686 B.n316 B.n5 163.367
R687 B.n6 B.n5 163.367
R688 B.n7 B.n6 163.367
R689 B.n321 B.n7 163.367
R690 B.n321 B.n12 163.367
R691 B.n13 B.n12 163.367
R692 B.n14 B.n13 163.367
R693 B.n326 B.n14 163.367
R694 B.n326 B.n19 163.367
R695 B.n20 B.n19 163.367
R696 B.n21 B.n20 163.367
R697 B.n331 B.n21 163.367
R698 B.n331 B.n26 163.367
R699 B.n27 B.n26 163.367
R700 B.n28 B.n27 163.367
R701 B.n336 B.n28 163.367
R702 B.n336 B.n33 163.367
R703 B.n34 B.n33 163.367
R704 B.n35 B.n34 163.367
R705 B.n341 B.n35 163.367
R706 B.n341 B.n40 163.367
R707 B.n41 B.n40 163.367
R708 B.n42 B.n41 163.367
R709 B.n448 B.n446 163.367
R710 B.n444 B.n46 163.367
R711 B.n440 B.n438 163.367
R712 B.n436 B.n48 163.367
R713 B.n432 B.n430 163.367
R714 B.n428 B.n50 163.367
R715 B.n424 B.n422 163.367
R716 B.n420 B.n52 163.367
R717 B.n416 B.n414 163.367
R718 B.n412 B.n54 163.367
R719 B.n407 B.n405 163.367
R720 B.n403 B.n58 163.367
R721 B.n399 B.n397 163.367
R722 B.n395 B.n60 163.367
R723 B.n391 B.n389 163.367
R724 B.n387 B.n62 163.367
R725 B.n383 B.n381 163.367
R726 B.n379 B.n67 163.367
R727 B.n375 B.n373 163.367
R728 B.n371 B.n69 163.367
R729 B.n367 B.n365 163.367
R730 B.n363 B.n71 163.367
R731 B.n359 B.n357 163.367
R732 B.n355 B.n73 163.367
R733 B.n351 B.n349 163.367
R734 B.n253 B.n117 129.785
R735 B.n453 B.n43 129.785
R736 B.n253 B.n113 71.7511
R737 B.n259 B.n113 71.7511
R738 B.n259 B.n109 71.7511
R739 B.n265 B.n109 71.7511
R740 B.n265 B.n105 71.7511
R741 B.n271 B.n105 71.7511
R742 B.n277 B.n101 71.7511
R743 B.n277 B.n97 71.7511
R744 B.n283 B.n97 71.7511
R745 B.n283 B.n93 71.7511
R746 B.n289 B.n93 71.7511
R747 B.n289 B.n89 71.7511
R748 B.n295 B.n89 71.7511
R749 B.n295 B.n85 71.7511
R750 B.n301 B.n85 71.7511
R751 B.n308 B.n81 71.7511
R752 B.n308 B.n77 71.7511
R753 B.n314 B.n77 71.7511
R754 B.n314 B.n4 71.7511
R755 B.n495 B.n4 71.7511
R756 B.n495 B.n494 71.7511
R757 B.n494 B.n493 71.7511
R758 B.n493 B.n8 71.7511
R759 B.n487 B.n8 71.7511
R760 B.n487 B.n486 71.7511
R761 B.n485 B.n15 71.7511
R762 B.n479 B.n15 71.7511
R763 B.n479 B.n478 71.7511
R764 B.n478 B.n477 71.7511
R765 B.n477 B.n22 71.7511
R766 B.n471 B.n22 71.7511
R767 B.n471 B.n470 71.7511
R768 B.n470 B.n469 71.7511
R769 B.n469 B.n29 71.7511
R770 B.n463 B.n462 71.7511
R771 B.n462 B.n461 71.7511
R772 B.n461 B.n36 71.7511
R773 B.n455 B.n36 71.7511
R774 B.n455 B.n454 71.7511
R775 B.n454 B.n453 71.7511
R776 B.n247 B.n118 71.676
R777 B.n245 B.n120 71.676
R778 B.n241 B.n240 71.676
R779 B.n234 B.n122 71.676
R780 B.n233 B.n232 71.676
R781 B.n226 B.n124 71.676
R782 B.n225 B.n224 71.676
R783 B.n218 B.n126 71.676
R784 B.n217 B.n216 71.676
R785 B.n210 B.n128 71.676
R786 B.n209 B.n132 71.676
R787 B.n205 B.n204 71.676
R788 B.n198 B.n134 71.676
R789 B.n197 B.n196 71.676
R790 B.n190 B.n136 71.676
R791 B.n189 B.n140 71.676
R792 B.n185 B.n184 71.676
R793 B.n178 B.n142 71.676
R794 B.n177 B.n176 71.676
R795 B.n170 B.n144 71.676
R796 B.n169 B.n168 71.676
R797 B.n162 B.n146 71.676
R798 B.n161 B.n160 71.676
R799 B.n154 B.n148 71.676
R800 B.n153 B.n152 71.676
R801 B.n447 B.n44 71.676
R802 B.n446 B.n445 71.676
R803 B.n439 B.n46 71.676
R804 B.n438 B.n437 71.676
R805 B.n431 B.n48 71.676
R806 B.n430 B.n429 71.676
R807 B.n423 B.n50 71.676
R808 B.n422 B.n421 71.676
R809 B.n415 B.n52 71.676
R810 B.n414 B.n413 71.676
R811 B.n406 B.n54 71.676
R812 B.n405 B.n404 71.676
R813 B.n398 B.n58 71.676
R814 B.n397 B.n396 71.676
R815 B.n390 B.n60 71.676
R816 B.n389 B.n388 71.676
R817 B.n382 B.n62 71.676
R818 B.n381 B.n380 71.676
R819 B.n374 B.n67 71.676
R820 B.n373 B.n372 71.676
R821 B.n366 B.n69 71.676
R822 B.n365 B.n364 71.676
R823 B.n358 B.n71 71.676
R824 B.n357 B.n356 71.676
R825 B.n350 B.n73 71.676
R826 B.n349 B.n348 71.676
R827 B.n348 B.n347 71.676
R828 B.n351 B.n350 71.676
R829 B.n356 B.n355 71.676
R830 B.n359 B.n358 71.676
R831 B.n364 B.n363 71.676
R832 B.n367 B.n366 71.676
R833 B.n372 B.n371 71.676
R834 B.n375 B.n374 71.676
R835 B.n380 B.n379 71.676
R836 B.n383 B.n382 71.676
R837 B.n388 B.n387 71.676
R838 B.n391 B.n390 71.676
R839 B.n396 B.n395 71.676
R840 B.n399 B.n398 71.676
R841 B.n404 B.n403 71.676
R842 B.n407 B.n406 71.676
R843 B.n413 B.n412 71.676
R844 B.n416 B.n415 71.676
R845 B.n421 B.n420 71.676
R846 B.n424 B.n423 71.676
R847 B.n429 B.n428 71.676
R848 B.n432 B.n431 71.676
R849 B.n437 B.n436 71.676
R850 B.n440 B.n439 71.676
R851 B.n445 B.n444 71.676
R852 B.n448 B.n447 71.676
R853 B.n248 B.n247 71.676
R854 B.n242 B.n120 71.676
R855 B.n240 B.n239 71.676
R856 B.n235 B.n234 71.676
R857 B.n232 B.n231 71.676
R858 B.n227 B.n226 71.676
R859 B.n224 B.n223 71.676
R860 B.n219 B.n218 71.676
R861 B.n216 B.n215 71.676
R862 B.n211 B.n210 71.676
R863 B.n206 B.n132 71.676
R864 B.n204 B.n203 71.676
R865 B.n199 B.n198 71.676
R866 B.n196 B.n195 71.676
R867 B.n191 B.n190 71.676
R868 B.n186 B.n140 71.676
R869 B.n184 B.n183 71.676
R870 B.n179 B.n178 71.676
R871 B.n176 B.n175 71.676
R872 B.n171 B.n170 71.676
R873 B.n168 B.n167 71.676
R874 B.n163 B.n162 71.676
R875 B.n160 B.n159 71.676
R876 B.n155 B.n154 71.676
R877 B.n152 B.n151 71.676
R878 B.n301 B.t1 66.4753
R879 B.t0 B.n485 66.4753
R880 B.n139 B.n138 59.5399
R881 B.n131 B.n130 59.5399
R882 B.n409 B.n56 59.5399
R883 B.n65 B.n64 59.5399
R884 B.n271 B.t3 55.9238
R885 B.n463 B.t7 55.9238
R886 B.n138 B.n137 45.7702
R887 B.n130 B.n129 45.7702
R888 B.n56 B.n55 45.7702
R889 B.n64 B.n63 45.7702
R890 B.n451 B.n450 35.1225
R891 B.n346 B.n345 35.1225
R892 B.n255 B.n115 35.1225
R893 B.n251 B.n250 35.1225
R894 B B.n497 18.0485
R895 B.t3 B.n101 15.8278
R896 B.t7 B.n29 15.8278
R897 B.n450 B.n449 10.6151
R898 B.n449 B.n45 10.6151
R899 B.n443 B.n45 10.6151
R900 B.n443 B.n442 10.6151
R901 B.n442 B.n441 10.6151
R902 B.n441 B.n47 10.6151
R903 B.n435 B.n47 10.6151
R904 B.n435 B.n434 10.6151
R905 B.n434 B.n433 10.6151
R906 B.n433 B.n49 10.6151
R907 B.n427 B.n49 10.6151
R908 B.n427 B.n426 10.6151
R909 B.n426 B.n425 10.6151
R910 B.n425 B.n51 10.6151
R911 B.n419 B.n51 10.6151
R912 B.n419 B.n418 10.6151
R913 B.n418 B.n417 10.6151
R914 B.n417 B.n53 10.6151
R915 B.n411 B.n53 10.6151
R916 B.n411 B.n410 10.6151
R917 B.n408 B.n57 10.6151
R918 B.n402 B.n57 10.6151
R919 B.n402 B.n401 10.6151
R920 B.n401 B.n400 10.6151
R921 B.n400 B.n59 10.6151
R922 B.n394 B.n59 10.6151
R923 B.n394 B.n393 10.6151
R924 B.n393 B.n392 10.6151
R925 B.n392 B.n61 10.6151
R926 B.n386 B.n385 10.6151
R927 B.n385 B.n384 10.6151
R928 B.n384 B.n66 10.6151
R929 B.n378 B.n66 10.6151
R930 B.n378 B.n377 10.6151
R931 B.n377 B.n376 10.6151
R932 B.n376 B.n68 10.6151
R933 B.n370 B.n68 10.6151
R934 B.n370 B.n369 10.6151
R935 B.n369 B.n368 10.6151
R936 B.n368 B.n70 10.6151
R937 B.n362 B.n70 10.6151
R938 B.n362 B.n361 10.6151
R939 B.n361 B.n360 10.6151
R940 B.n360 B.n72 10.6151
R941 B.n354 B.n72 10.6151
R942 B.n354 B.n353 10.6151
R943 B.n353 B.n352 10.6151
R944 B.n352 B.n74 10.6151
R945 B.n346 B.n74 10.6151
R946 B.n256 B.n255 10.6151
R947 B.n257 B.n256 10.6151
R948 B.n257 B.n107 10.6151
R949 B.n267 B.n107 10.6151
R950 B.n268 B.n267 10.6151
R951 B.n269 B.n268 10.6151
R952 B.n269 B.n99 10.6151
R953 B.n279 B.n99 10.6151
R954 B.n280 B.n279 10.6151
R955 B.n281 B.n280 10.6151
R956 B.n281 B.n91 10.6151
R957 B.n291 B.n91 10.6151
R958 B.n292 B.n291 10.6151
R959 B.n293 B.n292 10.6151
R960 B.n293 B.n83 10.6151
R961 B.n303 B.n83 10.6151
R962 B.n304 B.n303 10.6151
R963 B.n306 B.n304 10.6151
R964 B.n306 B.n305 10.6151
R965 B.n305 B.n75 10.6151
R966 B.n317 B.n75 10.6151
R967 B.n318 B.n317 10.6151
R968 B.n319 B.n318 10.6151
R969 B.n320 B.n319 10.6151
R970 B.n322 B.n320 10.6151
R971 B.n323 B.n322 10.6151
R972 B.n324 B.n323 10.6151
R973 B.n325 B.n324 10.6151
R974 B.n327 B.n325 10.6151
R975 B.n328 B.n327 10.6151
R976 B.n329 B.n328 10.6151
R977 B.n330 B.n329 10.6151
R978 B.n332 B.n330 10.6151
R979 B.n333 B.n332 10.6151
R980 B.n334 B.n333 10.6151
R981 B.n335 B.n334 10.6151
R982 B.n337 B.n335 10.6151
R983 B.n338 B.n337 10.6151
R984 B.n339 B.n338 10.6151
R985 B.n340 B.n339 10.6151
R986 B.n342 B.n340 10.6151
R987 B.n343 B.n342 10.6151
R988 B.n344 B.n343 10.6151
R989 B.n345 B.n344 10.6151
R990 B.n250 B.n249 10.6151
R991 B.n249 B.n119 10.6151
R992 B.n244 B.n119 10.6151
R993 B.n244 B.n243 10.6151
R994 B.n243 B.n121 10.6151
R995 B.n238 B.n121 10.6151
R996 B.n238 B.n237 10.6151
R997 B.n237 B.n236 10.6151
R998 B.n236 B.n123 10.6151
R999 B.n230 B.n123 10.6151
R1000 B.n230 B.n229 10.6151
R1001 B.n229 B.n228 10.6151
R1002 B.n228 B.n125 10.6151
R1003 B.n222 B.n125 10.6151
R1004 B.n222 B.n221 10.6151
R1005 B.n221 B.n220 10.6151
R1006 B.n220 B.n127 10.6151
R1007 B.n214 B.n127 10.6151
R1008 B.n214 B.n213 10.6151
R1009 B.n213 B.n212 10.6151
R1010 B.n208 B.n207 10.6151
R1011 B.n207 B.n133 10.6151
R1012 B.n202 B.n133 10.6151
R1013 B.n202 B.n201 10.6151
R1014 B.n201 B.n200 10.6151
R1015 B.n200 B.n135 10.6151
R1016 B.n194 B.n135 10.6151
R1017 B.n194 B.n193 10.6151
R1018 B.n193 B.n192 10.6151
R1019 B.n188 B.n187 10.6151
R1020 B.n187 B.n141 10.6151
R1021 B.n182 B.n141 10.6151
R1022 B.n182 B.n181 10.6151
R1023 B.n181 B.n180 10.6151
R1024 B.n180 B.n143 10.6151
R1025 B.n174 B.n143 10.6151
R1026 B.n174 B.n173 10.6151
R1027 B.n173 B.n172 10.6151
R1028 B.n172 B.n145 10.6151
R1029 B.n166 B.n145 10.6151
R1030 B.n166 B.n165 10.6151
R1031 B.n165 B.n164 10.6151
R1032 B.n164 B.n147 10.6151
R1033 B.n158 B.n147 10.6151
R1034 B.n158 B.n157 10.6151
R1035 B.n157 B.n156 10.6151
R1036 B.n156 B.n149 10.6151
R1037 B.n150 B.n149 10.6151
R1038 B.n150 B.n115 10.6151
R1039 B.n251 B.n111 10.6151
R1040 B.n261 B.n111 10.6151
R1041 B.n262 B.n261 10.6151
R1042 B.n263 B.n262 10.6151
R1043 B.n263 B.n103 10.6151
R1044 B.n273 B.n103 10.6151
R1045 B.n274 B.n273 10.6151
R1046 B.n275 B.n274 10.6151
R1047 B.n275 B.n95 10.6151
R1048 B.n285 B.n95 10.6151
R1049 B.n286 B.n285 10.6151
R1050 B.n287 B.n286 10.6151
R1051 B.n287 B.n87 10.6151
R1052 B.n297 B.n87 10.6151
R1053 B.n298 B.n297 10.6151
R1054 B.n299 B.n298 10.6151
R1055 B.n299 B.n79 10.6151
R1056 B.n310 B.n79 10.6151
R1057 B.n311 B.n310 10.6151
R1058 B.n312 B.n311 10.6151
R1059 B.n312 B.n0 10.6151
R1060 B.n491 B.n1 10.6151
R1061 B.n491 B.n490 10.6151
R1062 B.n490 B.n489 10.6151
R1063 B.n489 B.n10 10.6151
R1064 B.n483 B.n10 10.6151
R1065 B.n483 B.n482 10.6151
R1066 B.n482 B.n481 10.6151
R1067 B.n481 B.n17 10.6151
R1068 B.n475 B.n17 10.6151
R1069 B.n475 B.n474 10.6151
R1070 B.n474 B.n473 10.6151
R1071 B.n473 B.n24 10.6151
R1072 B.n467 B.n24 10.6151
R1073 B.n467 B.n466 10.6151
R1074 B.n466 B.n465 10.6151
R1075 B.n465 B.n31 10.6151
R1076 B.n459 B.n31 10.6151
R1077 B.n459 B.n458 10.6151
R1078 B.n458 B.n457 10.6151
R1079 B.n457 B.n38 10.6151
R1080 B.n451 B.n38 10.6151
R1081 B.n410 B.n409 9.36635
R1082 B.n386 B.n65 9.36635
R1083 B.n212 B.n131 9.36635
R1084 B.n188 B.n139 9.36635
R1085 B.t1 B.n81 5.27628
R1086 B.n486 B.t0 5.27628
R1087 B.n497 B.n0 2.81026
R1088 B.n497 B.n1 2.81026
R1089 B.n409 B.n408 1.24928
R1090 B.n65 B.n61 1.24928
R1091 B.n208 B.n131 1.24928
R1092 B.n192 B.n139 1.24928
R1093 VP.n0 VP.t0 157.957
R1094 VP.n0 VP.t1 120.001
R1095 VP VP.n0 0.241678
R1096 VDD1.n24 VDD1.n23 289.615
R1097 VDD1.n49 VDD1.n48 289.615
R1098 VDD1.n23 VDD1.n22 185
R1099 VDD1.n2 VDD1.n1 185
R1100 VDD1.n17 VDD1.n16 185
R1101 VDD1.n15 VDD1.n14 185
R1102 VDD1.n6 VDD1.n5 185
R1103 VDD1.n9 VDD1.n8 185
R1104 VDD1.n34 VDD1.n33 185
R1105 VDD1.n31 VDD1.n30 185
R1106 VDD1.n40 VDD1.n39 185
R1107 VDD1.n42 VDD1.n41 185
R1108 VDD1.n27 VDD1.n26 185
R1109 VDD1.n48 VDD1.n47 185
R1110 VDD1.t0 VDD1.n32 149.54
R1111 VDD1.t1 VDD1.n7 149.54
R1112 VDD1.n23 VDD1.n1 104.615
R1113 VDD1.n16 VDD1.n1 104.615
R1114 VDD1.n16 VDD1.n15 104.615
R1115 VDD1.n15 VDD1.n5 104.615
R1116 VDD1.n8 VDD1.n5 104.615
R1117 VDD1.n33 VDD1.n30 104.615
R1118 VDD1.n40 VDD1.n30 104.615
R1119 VDD1.n41 VDD1.n40 104.615
R1120 VDD1.n41 VDD1.n26 104.615
R1121 VDD1.n48 VDD1.n26 104.615
R1122 VDD1 VDD1.n49 84.5869
R1123 VDD1.n8 VDD1.t1 52.3082
R1124 VDD1.n33 VDD1.t0 52.3082
R1125 VDD1 VDD1.n24 51.9522
R1126 VDD1.n22 VDD1.n0 11.249
R1127 VDD1.n47 VDD1.n25 11.249
R1128 VDD1.n21 VDD1.n2 10.4732
R1129 VDD1.n46 VDD1.n27 10.4732
R1130 VDD1.n9 VDD1.n7 10.2739
R1131 VDD1.n34 VDD1.n32 10.2739
R1132 VDD1.n18 VDD1.n17 9.69747
R1133 VDD1.n43 VDD1.n42 9.69747
R1134 VDD1.n20 VDD1.n0 9.45567
R1135 VDD1.n45 VDD1.n25 9.45567
R1136 VDD1.n21 VDD1.n20 9.3005
R1137 VDD1.n19 VDD1.n18 9.3005
R1138 VDD1.n4 VDD1.n3 9.3005
R1139 VDD1.n13 VDD1.n12 9.3005
R1140 VDD1.n11 VDD1.n10 9.3005
R1141 VDD1.n36 VDD1.n35 9.3005
R1142 VDD1.n38 VDD1.n37 9.3005
R1143 VDD1.n29 VDD1.n28 9.3005
R1144 VDD1.n44 VDD1.n43 9.3005
R1145 VDD1.n46 VDD1.n45 9.3005
R1146 VDD1.n14 VDD1.n4 8.92171
R1147 VDD1.n39 VDD1.n29 8.92171
R1148 VDD1.n13 VDD1.n6 8.14595
R1149 VDD1.n38 VDD1.n31 8.14595
R1150 VDD1.n10 VDD1.n9 7.3702
R1151 VDD1.n35 VDD1.n34 7.3702
R1152 VDD1.n10 VDD1.n6 5.81868
R1153 VDD1.n35 VDD1.n31 5.81868
R1154 VDD1.n14 VDD1.n13 5.04292
R1155 VDD1.n39 VDD1.n38 5.04292
R1156 VDD1.n17 VDD1.n4 4.26717
R1157 VDD1.n42 VDD1.n29 4.26717
R1158 VDD1.n18 VDD1.n2 3.49141
R1159 VDD1.n43 VDD1.n27 3.49141
R1160 VDD1.n36 VDD1.n32 2.84386
R1161 VDD1.n11 VDD1.n7 2.84386
R1162 VDD1.n22 VDD1.n21 2.71565
R1163 VDD1.n47 VDD1.n46 2.71565
R1164 VDD1.n24 VDD1.n0 1.93989
R1165 VDD1.n49 VDD1.n25 1.93989
R1166 VDD1.n20 VDD1.n19 0.155672
R1167 VDD1.n19 VDD1.n3 0.155672
R1168 VDD1.n12 VDD1.n3 0.155672
R1169 VDD1.n12 VDD1.n11 0.155672
R1170 VDD1.n37 VDD1.n36 0.155672
R1171 VDD1.n37 VDD1.n28 0.155672
R1172 VDD1.n44 VDD1.n28 0.155672
R1173 VDD1.n45 VDD1.n44 0.155672
C0 VN VP 3.91699f
C1 VN VTAIL 1.29223f
C2 VDD2 VDD1 0.605857f
C3 VTAIL VP 1.30644f
C4 VN VDD2 1.28747f
C5 VDD2 VP 0.312488f
C6 VDD2 VTAIL 3.16872f
C7 VN VDD1 0.147861f
C8 VDD1 VP 1.44668f
C9 VTAIL VDD1 3.12066f
C10 VDD2 B 2.962811f
C11 VDD1 B 4.4619f
C12 VTAIL B 4.150546f
C13 VN B 7.125051f
C14 VP B 5.096155f
C15 VDD1.n0 B 0.008109f
C16 VDD1.n1 B 0.018245f
C17 VDD1.n2 B 0.008173f
C18 VDD1.n3 B 0.014365f
C19 VDD1.n4 B 0.007719f
C20 VDD1.n5 B 0.018245f
C21 VDD1.n6 B 0.008173f
C22 VDD1.n7 B 0.066081f
C23 VDD1.t1 B 0.030443f
C24 VDD1.n8 B 0.013684f
C25 VDD1.n9 B 0.012895f
C26 VDD1.n10 B 0.007719f
C27 VDD1.n11 B 0.286566f
C28 VDD1.n12 B 0.014365f
C29 VDD1.n13 B 0.007719f
C30 VDD1.n14 B 0.008173f
C31 VDD1.n15 B 0.018245f
C32 VDD1.n16 B 0.018245f
C33 VDD1.n17 B 0.008173f
C34 VDD1.n18 B 0.007719f
C35 VDD1.n19 B 0.014365f
C36 VDD1.n20 B 0.037717f
C37 VDD1.n21 B 0.007719f
C38 VDD1.n22 B 0.008173f
C39 VDD1.n23 B 0.036583f
C40 VDD1.n24 B 0.041898f
C41 VDD1.n25 B 0.008109f
C42 VDD1.n26 B 0.018245f
C43 VDD1.n27 B 0.008173f
C44 VDD1.n28 B 0.014365f
C45 VDD1.n29 B 0.007719f
C46 VDD1.n30 B 0.018245f
C47 VDD1.n31 B 0.008173f
C48 VDD1.n32 B 0.066081f
C49 VDD1.t0 B 0.030443f
C50 VDD1.n33 B 0.013684f
C51 VDD1.n34 B 0.012895f
C52 VDD1.n35 B 0.007719f
C53 VDD1.n36 B 0.286566f
C54 VDD1.n37 B 0.014365f
C55 VDD1.n38 B 0.007719f
C56 VDD1.n39 B 0.008173f
C57 VDD1.n40 B 0.018245f
C58 VDD1.n41 B 0.018245f
C59 VDD1.n42 B 0.008173f
C60 VDD1.n43 B 0.007719f
C61 VDD1.n44 B 0.014365f
C62 VDD1.n45 B 0.037717f
C63 VDD1.n46 B 0.007719f
C64 VDD1.n47 B 0.008173f
C65 VDD1.n48 B 0.036583f
C66 VDD1.n49 B 0.29775f
C67 VP.t0 B 1.11126f
C68 VP.t1 B 0.849551f
C69 VP.n0 B 1.89834f
C70 VDD2.n0 B 0.008516f
C71 VDD2.n1 B 0.019161f
C72 VDD2.n2 B 0.008584f
C73 VDD2.n3 B 0.015086f
C74 VDD2.n4 B 0.008107f
C75 VDD2.n5 B 0.019161f
C76 VDD2.n6 B 0.008584f
C77 VDD2.n7 B 0.0694f
C78 VDD2.t1 B 0.031972f
C79 VDD2.n8 B 0.014371f
C80 VDD2.n9 B 0.013542f
C81 VDD2.n10 B 0.008107f
C82 VDD2.n11 B 0.30096f
C83 VDD2.n12 B 0.015086f
C84 VDD2.n13 B 0.008107f
C85 VDD2.n14 B 0.008584f
C86 VDD2.n15 B 0.019161f
C87 VDD2.n16 B 0.019161f
C88 VDD2.n17 B 0.008584f
C89 VDD2.n18 B 0.008107f
C90 VDD2.n19 B 0.015086f
C91 VDD2.n20 B 0.039611f
C92 VDD2.n21 B 0.008107f
C93 VDD2.n22 B 0.008584f
C94 VDD2.n23 B 0.038421f
C95 VDD2.n24 B 0.290225f
C96 VDD2.n25 B 0.008516f
C97 VDD2.n26 B 0.019161f
C98 VDD2.n27 B 0.008584f
C99 VDD2.n28 B 0.015086f
C100 VDD2.n29 B 0.008107f
C101 VDD2.n30 B 0.019161f
C102 VDD2.n31 B 0.008584f
C103 VDD2.n32 B 0.0694f
C104 VDD2.t0 B 0.031972f
C105 VDD2.n33 B 0.014371f
C106 VDD2.n34 B 0.013542f
C107 VDD2.n35 B 0.008107f
C108 VDD2.n36 B 0.30096f
C109 VDD2.n37 B 0.015086f
C110 VDD2.n38 B 0.008107f
C111 VDD2.n39 B 0.008584f
C112 VDD2.n40 B 0.019161f
C113 VDD2.n41 B 0.019161f
C114 VDD2.n42 B 0.008584f
C115 VDD2.n43 B 0.008107f
C116 VDD2.n44 B 0.015086f
C117 VDD2.n45 B 0.039611f
C118 VDD2.n46 B 0.008107f
C119 VDD2.n47 B 0.008584f
C120 VDD2.n48 B 0.038421f
C121 VDD2.n49 B 0.043369f
C122 VDD2.n50 B 1.34469f
C123 VTAIL.n0 B 0.009506f
C124 VTAIL.n1 B 0.02139f
C125 VTAIL.n2 B 0.009582f
C126 VTAIL.n3 B 0.016841f
C127 VTAIL.n4 B 0.00905f
C128 VTAIL.n5 B 0.02139f
C129 VTAIL.n6 B 0.009582f
C130 VTAIL.n7 B 0.077472f
C131 VTAIL.t1 B 0.035691f
C132 VTAIL.n8 B 0.016042f
C133 VTAIL.n9 B 0.015118f
C134 VTAIL.n10 B 0.00905f
C135 VTAIL.n11 B 0.335964f
C136 VTAIL.n12 B 0.016841f
C137 VTAIL.n13 B 0.00905f
C138 VTAIL.n14 B 0.009582f
C139 VTAIL.n15 B 0.02139f
C140 VTAIL.n16 B 0.02139f
C141 VTAIL.n17 B 0.009582f
C142 VTAIL.n18 B 0.00905f
C143 VTAIL.n19 B 0.016841f
C144 VTAIL.n20 B 0.044218f
C145 VTAIL.n21 B 0.00905f
C146 VTAIL.n22 B 0.009582f
C147 VTAIL.n23 B 0.04289f
C148 VTAIL.n24 B 0.036806f
C149 VTAIL.n25 B 0.762811f
C150 VTAIL.n26 B 0.009506f
C151 VTAIL.n27 B 0.02139f
C152 VTAIL.n28 B 0.009582f
C153 VTAIL.n29 B 0.016841f
C154 VTAIL.n30 B 0.00905f
C155 VTAIL.n31 B 0.02139f
C156 VTAIL.n32 B 0.009582f
C157 VTAIL.n33 B 0.077472f
C158 VTAIL.t3 B 0.035691f
C159 VTAIL.n34 B 0.016042f
C160 VTAIL.n35 B 0.015118f
C161 VTAIL.n36 B 0.00905f
C162 VTAIL.n37 B 0.335964f
C163 VTAIL.n38 B 0.016841f
C164 VTAIL.n39 B 0.00905f
C165 VTAIL.n40 B 0.009582f
C166 VTAIL.n41 B 0.02139f
C167 VTAIL.n42 B 0.02139f
C168 VTAIL.n43 B 0.009582f
C169 VTAIL.n44 B 0.00905f
C170 VTAIL.n45 B 0.016841f
C171 VTAIL.n46 B 0.044218f
C172 VTAIL.n47 B 0.00905f
C173 VTAIL.n48 B 0.009582f
C174 VTAIL.n49 B 0.04289f
C175 VTAIL.n50 B 0.036806f
C176 VTAIL.n51 B 0.787254f
C177 VTAIL.n52 B 0.009506f
C178 VTAIL.n53 B 0.02139f
C179 VTAIL.n54 B 0.009582f
C180 VTAIL.n55 B 0.016841f
C181 VTAIL.n56 B 0.00905f
C182 VTAIL.n57 B 0.02139f
C183 VTAIL.n58 B 0.009582f
C184 VTAIL.n59 B 0.077472f
C185 VTAIL.t0 B 0.035691f
C186 VTAIL.n60 B 0.016042f
C187 VTAIL.n61 B 0.015118f
C188 VTAIL.n62 B 0.00905f
C189 VTAIL.n63 B 0.335964f
C190 VTAIL.n64 B 0.016841f
C191 VTAIL.n65 B 0.00905f
C192 VTAIL.n66 B 0.009582f
C193 VTAIL.n67 B 0.02139f
C194 VTAIL.n68 B 0.02139f
C195 VTAIL.n69 B 0.009582f
C196 VTAIL.n70 B 0.00905f
C197 VTAIL.n71 B 0.016841f
C198 VTAIL.n72 B 0.044218f
C199 VTAIL.n73 B 0.00905f
C200 VTAIL.n74 B 0.009582f
C201 VTAIL.n75 B 0.04289f
C202 VTAIL.n76 B 0.036806f
C203 VTAIL.n77 B 0.676853f
C204 VTAIL.n78 B 0.009506f
C205 VTAIL.n79 B 0.02139f
C206 VTAIL.n80 B 0.009582f
C207 VTAIL.n81 B 0.016841f
C208 VTAIL.n82 B 0.00905f
C209 VTAIL.n83 B 0.02139f
C210 VTAIL.n84 B 0.009582f
C211 VTAIL.n85 B 0.077472f
C212 VTAIL.t2 B 0.035691f
C213 VTAIL.n86 B 0.016042f
C214 VTAIL.n87 B 0.015118f
C215 VTAIL.n88 B 0.00905f
C216 VTAIL.n89 B 0.335964f
C217 VTAIL.n90 B 0.016841f
C218 VTAIL.n91 B 0.00905f
C219 VTAIL.n92 B 0.009582f
C220 VTAIL.n93 B 0.02139f
C221 VTAIL.n94 B 0.02139f
C222 VTAIL.n95 B 0.009582f
C223 VTAIL.n96 B 0.00905f
C224 VTAIL.n97 B 0.016841f
C225 VTAIL.n98 B 0.044218f
C226 VTAIL.n99 B 0.00905f
C227 VTAIL.n100 B 0.009582f
C228 VTAIL.n101 B 0.04289f
C229 VTAIL.n102 B 0.036806f
C230 VTAIL.n103 B 0.620599f
C231 VN.t0 B 0.84282f
C232 VN.t1 B 1.1055f
.ends

