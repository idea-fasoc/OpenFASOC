* NGSPICE file created from diff_pair_sample_0470.ext - technology: sky130A

.subckt diff_pair_sample_0470 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t7 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=5.148 pd=27.18 as=2.178 ps=13.53 w=13.2 l=3.58
X1 B.t11 B.t9 B.t10 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=5.148 pd=27.18 as=0 ps=0 w=13.2 l=3.58
X2 VDD2.t9 VN.t0 VTAIL.t17 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=5.148 ps=27.18 w=13.2 l=3.58
X3 VDD1.t8 VP.t1 VTAIL.t8 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=5.148 ps=27.18 w=13.2 l=3.58
X4 VDD2.t8 VN.t1 VTAIL.t18 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=2.178 ps=13.53 w=13.2 l=3.58
X5 VTAIL.t19 VN.t2 VDD2.t7 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=2.178 ps=13.53 w=13.2 l=3.58
X6 VDD2.t6 VN.t3 VTAIL.t2 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=5.148 pd=27.18 as=2.178 ps=13.53 w=13.2 l=3.58
X7 VDD1.t7 VP.t2 VTAIL.t13 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=5.148 pd=27.18 as=2.178 ps=13.53 w=13.2 l=3.58
X8 B.t8 B.t6 B.t7 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=5.148 pd=27.18 as=0 ps=0 w=13.2 l=3.58
X9 B.t5 B.t3 B.t4 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=5.148 pd=27.18 as=0 ps=0 w=13.2 l=3.58
X10 VTAIL.t1 VN.t4 VDD2.t5 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=2.178 ps=13.53 w=13.2 l=3.58
X11 VDD2.t4 VN.t5 VTAIL.t6 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=5.148 ps=27.18 w=13.2 l=3.58
X12 VTAIL.t5 VN.t6 VDD2.t3 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=2.178 ps=13.53 w=13.2 l=3.58
X13 VTAIL.t16 VP.t3 VDD1.t6 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=2.178 ps=13.53 w=13.2 l=3.58
X14 VDD2.t2 VN.t7 VTAIL.t4 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=2.178 ps=13.53 w=13.2 l=3.58
X15 VTAIL.t14 VP.t4 VDD1.t5 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=2.178 ps=13.53 w=13.2 l=3.58
X16 VDD2.t1 VN.t8 VTAIL.t0 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=5.148 pd=27.18 as=2.178 ps=13.53 w=13.2 l=3.58
X17 VDD1.t4 VP.t5 VTAIL.t12 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=2.178 ps=13.53 w=13.2 l=3.58
X18 VDD1.t3 VP.t6 VTAIL.t10 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=5.148 ps=27.18 w=13.2 l=3.58
X19 VDD1.t2 VP.t7 VTAIL.t9 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=2.178 ps=13.53 w=13.2 l=3.58
X20 VTAIL.t11 VP.t8 VDD1.t1 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=2.178 ps=13.53 w=13.2 l=3.58
X21 B.t2 B.t0 B.t1 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=5.148 pd=27.18 as=0 ps=0 w=13.2 l=3.58
X22 VTAIL.t15 VP.t9 VDD1.t0 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=2.178 ps=13.53 w=13.2 l=3.58
X23 VTAIL.t3 VN.t9 VDD2.t0 w_n5662_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=2.178 ps=13.53 w=13.2 l=3.58
R0 VP.n32 VP.n29 161.3
R1 VP.n34 VP.n33 161.3
R2 VP.n35 VP.n28 161.3
R3 VP.n37 VP.n36 161.3
R4 VP.n38 VP.n27 161.3
R5 VP.n40 VP.n39 161.3
R6 VP.n41 VP.n26 161.3
R7 VP.n44 VP.n43 161.3
R8 VP.n45 VP.n25 161.3
R9 VP.n47 VP.n46 161.3
R10 VP.n48 VP.n24 161.3
R11 VP.n50 VP.n49 161.3
R12 VP.n51 VP.n23 161.3
R13 VP.n53 VP.n52 161.3
R14 VP.n54 VP.n22 161.3
R15 VP.n57 VP.n56 161.3
R16 VP.n58 VP.n21 161.3
R17 VP.n60 VP.n59 161.3
R18 VP.n61 VP.n20 161.3
R19 VP.n63 VP.n62 161.3
R20 VP.n64 VP.n19 161.3
R21 VP.n66 VP.n65 161.3
R22 VP.n67 VP.n18 161.3
R23 VP.n69 VP.n68 161.3
R24 VP.n123 VP.n122 161.3
R25 VP.n121 VP.n1 161.3
R26 VP.n120 VP.n119 161.3
R27 VP.n118 VP.n2 161.3
R28 VP.n117 VP.n116 161.3
R29 VP.n115 VP.n3 161.3
R30 VP.n114 VP.n113 161.3
R31 VP.n112 VP.n4 161.3
R32 VP.n111 VP.n110 161.3
R33 VP.n108 VP.n5 161.3
R34 VP.n107 VP.n106 161.3
R35 VP.n105 VP.n6 161.3
R36 VP.n104 VP.n103 161.3
R37 VP.n102 VP.n7 161.3
R38 VP.n101 VP.n100 161.3
R39 VP.n99 VP.n8 161.3
R40 VP.n98 VP.n97 161.3
R41 VP.n95 VP.n9 161.3
R42 VP.n94 VP.n93 161.3
R43 VP.n92 VP.n10 161.3
R44 VP.n91 VP.n90 161.3
R45 VP.n89 VP.n11 161.3
R46 VP.n88 VP.n87 161.3
R47 VP.n86 VP.n12 161.3
R48 VP.n85 VP.n84 161.3
R49 VP.n82 VP.n13 161.3
R50 VP.n81 VP.n80 161.3
R51 VP.n79 VP.n14 161.3
R52 VP.n78 VP.n77 161.3
R53 VP.n76 VP.n15 161.3
R54 VP.n75 VP.n74 161.3
R55 VP.n73 VP.n16 161.3
R56 VP.n31 VP.t0 120.98
R57 VP.n71 VP.t2 88.8608
R58 VP.n83 VP.t4 88.8608
R59 VP.n96 VP.t7 88.8608
R60 VP.n109 VP.t8 88.8608
R61 VP.n0 VP.t6 88.8608
R62 VP.n17 VP.t1 88.8608
R63 VP.n55 VP.t9 88.8608
R64 VP.n42 VP.t5 88.8608
R65 VP.n30 VP.t3 88.8608
R66 VP.n72 VP.n71 86.8027
R67 VP.n124 VP.n0 86.8027
R68 VP.n70 VP.n17 86.8027
R69 VP.n31 VP.n30 67.0059
R70 VP.n72 VP.n70 59.3594
R71 VP.n90 VP.n10 56.5617
R72 VP.n103 VP.n6 56.5617
R73 VP.n49 VP.n23 56.5617
R74 VP.n36 VP.n27 56.5617
R75 VP.n77 VP.n14 51.7179
R76 VP.n116 VP.n2 51.7179
R77 VP.n62 VP.n19 51.7179
R78 VP.n81 VP.n14 29.4362
R79 VP.n116 VP.n115 29.4362
R80 VP.n62 VP.n61 29.4362
R81 VP.n75 VP.n16 24.5923
R82 VP.n76 VP.n75 24.5923
R83 VP.n77 VP.n76 24.5923
R84 VP.n82 VP.n81 24.5923
R85 VP.n84 VP.n82 24.5923
R86 VP.n88 VP.n12 24.5923
R87 VP.n89 VP.n88 24.5923
R88 VP.n90 VP.n89 24.5923
R89 VP.n94 VP.n10 24.5923
R90 VP.n95 VP.n94 24.5923
R91 VP.n97 VP.n95 24.5923
R92 VP.n101 VP.n8 24.5923
R93 VP.n102 VP.n101 24.5923
R94 VP.n103 VP.n102 24.5923
R95 VP.n107 VP.n6 24.5923
R96 VP.n108 VP.n107 24.5923
R97 VP.n110 VP.n108 24.5923
R98 VP.n114 VP.n4 24.5923
R99 VP.n115 VP.n114 24.5923
R100 VP.n120 VP.n2 24.5923
R101 VP.n121 VP.n120 24.5923
R102 VP.n122 VP.n121 24.5923
R103 VP.n66 VP.n19 24.5923
R104 VP.n67 VP.n66 24.5923
R105 VP.n68 VP.n67 24.5923
R106 VP.n53 VP.n23 24.5923
R107 VP.n54 VP.n53 24.5923
R108 VP.n56 VP.n54 24.5923
R109 VP.n60 VP.n21 24.5923
R110 VP.n61 VP.n60 24.5923
R111 VP.n40 VP.n27 24.5923
R112 VP.n41 VP.n40 24.5923
R113 VP.n43 VP.n41 24.5923
R114 VP.n47 VP.n25 24.5923
R115 VP.n48 VP.n47 24.5923
R116 VP.n49 VP.n48 24.5923
R117 VP.n34 VP.n29 24.5923
R118 VP.n35 VP.n34 24.5923
R119 VP.n36 VP.n35 24.5923
R120 VP.n84 VP.n83 16.7229
R121 VP.n109 VP.n4 16.7229
R122 VP.n55 VP.n21 16.7229
R123 VP.n97 VP.n96 12.2964
R124 VP.n96 VP.n8 12.2964
R125 VP.n43 VP.n42 12.2964
R126 VP.n42 VP.n25 12.2964
R127 VP.n83 VP.n12 7.86989
R128 VP.n110 VP.n109 7.86989
R129 VP.n56 VP.n55 7.86989
R130 VP.n30 VP.n29 7.86989
R131 VP.n71 VP.n16 3.44336
R132 VP.n122 VP.n0 3.44336
R133 VP.n68 VP.n17 3.44336
R134 VP.n32 VP.n31 3.35171
R135 VP.n70 VP.n69 0.354861
R136 VP.n73 VP.n72 0.354861
R137 VP.n124 VP.n123 0.354861
R138 VP VP.n124 0.267071
R139 VP.n33 VP.n32 0.189894
R140 VP.n33 VP.n28 0.189894
R141 VP.n37 VP.n28 0.189894
R142 VP.n38 VP.n37 0.189894
R143 VP.n39 VP.n38 0.189894
R144 VP.n39 VP.n26 0.189894
R145 VP.n44 VP.n26 0.189894
R146 VP.n45 VP.n44 0.189894
R147 VP.n46 VP.n45 0.189894
R148 VP.n46 VP.n24 0.189894
R149 VP.n50 VP.n24 0.189894
R150 VP.n51 VP.n50 0.189894
R151 VP.n52 VP.n51 0.189894
R152 VP.n52 VP.n22 0.189894
R153 VP.n57 VP.n22 0.189894
R154 VP.n58 VP.n57 0.189894
R155 VP.n59 VP.n58 0.189894
R156 VP.n59 VP.n20 0.189894
R157 VP.n63 VP.n20 0.189894
R158 VP.n64 VP.n63 0.189894
R159 VP.n65 VP.n64 0.189894
R160 VP.n65 VP.n18 0.189894
R161 VP.n69 VP.n18 0.189894
R162 VP.n74 VP.n73 0.189894
R163 VP.n74 VP.n15 0.189894
R164 VP.n78 VP.n15 0.189894
R165 VP.n79 VP.n78 0.189894
R166 VP.n80 VP.n79 0.189894
R167 VP.n80 VP.n13 0.189894
R168 VP.n85 VP.n13 0.189894
R169 VP.n86 VP.n85 0.189894
R170 VP.n87 VP.n86 0.189894
R171 VP.n87 VP.n11 0.189894
R172 VP.n91 VP.n11 0.189894
R173 VP.n92 VP.n91 0.189894
R174 VP.n93 VP.n92 0.189894
R175 VP.n93 VP.n9 0.189894
R176 VP.n98 VP.n9 0.189894
R177 VP.n99 VP.n98 0.189894
R178 VP.n100 VP.n99 0.189894
R179 VP.n100 VP.n7 0.189894
R180 VP.n104 VP.n7 0.189894
R181 VP.n105 VP.n104 0.189894
R182 VP.n106 VP.n105 0.189894
R183 VP.n106 VP.n5 0.189894
R184 VP.n111 VP.n5 0.189894
R185 VP.n112 VP.n111 0.189894
R186 VP.n113 VP.n112 0.189894
R187 VP.n113 VP.n3 0.189894
R188 VP.n117 VP.n3 0.189894
R189 VP.n118 VP.n117 0.189894
R190 VP.n119 VP.n118 0.189894
R191 VP.n119 VP.n1 0.189894
R192 VP.n123 VP.n1 0.189894
R193 VTAIL.n11 VTAIL.t6 58.4184
R194 VTAIL.n17 VTAIL.t17 58.4181
R195 VTAIL.n2 VTAIL.t10 58.4181
R196 VTAIL.n16 VTAIL.t8 58.4181
R197 VTAIL.n15 VTAIL.n14 55.9559
R198 VTAIL.n13 VTAIL.n12 55.9559
R199 VTAIL.n10 VTAIL.n9 55.9559
R200 VTAIL.n8 VTAIL.n7 55.9559
R201 VTAIL.n19 VTAIL.n18 55.9558
R202 VTAIL.n1 VTAIL.n0 55.9558
R203 VTAIL.n4 VTAIL.n3 55.9558
R204 VTAIL.n6 VTAIL.n5 55.9558
R205 VTAIL.n8 VTAIL.n6 30.4876
R206 VTAIL.n17 VTAIL.n16 27.1169
R207 VTAIL.n10 VTAIL.n8 3.37119
R208 VTAIL.n11 VTAIL.n10 3.37119
R209 VTAIL.n15 VTAIL.n13 3.37119
R210 VTAIL.n16 VTAIL.n15 3.37119
R211 VTAIL.n6 VTAIL.n4 3.37119
R212 VTAIL.n4 VTAIL.n2 3.37119
R213 VTAIL.n19 VTAIL.n17 3.37119
R214 VTAIL VTAIL.n1 2.58671
R215 VTAIL.n18 VTAIL.t18 2.463
R216 VTAIL.n18 VTAIL.t19 2.463
R217 VTAIL.n0 VTAIL.t2 2.463
R218 VTAIL.n0 VTAIL.t1 2.463
R219 VTAIL.n3 VTAIL.t9 2.463
R220 VTAIL.n3 VTAIL.t11 2.463
R221 VTAIL.n5 VTAIL.t13 2.463
R222 VTAIL.n5 VTAIL.t14 2.463
R223 VTAIL.n14 VTAIL.t12 2.463
R224 VTAIL.n14 VTAIL.t15 2.463
R225 VTAIL.n12 VTAIL.t7 2.463
R226 VTAIL.n12 VTAIL.t16 2.463
R227 VTAIL.n9 VTAIL.t4 2.463
R228 VTAIL.n9 VTAIL.t3 2.463
R229 VTAIL.n7 VTAIL.t0 2.463
R230 VTAIL.n7 VTAIL.t5 2.463
R231 VTAIL.n13 VTAIL.n11 2.15567
R232 VTAIL.n2 VTAIL.n1 2.15567
R233 VTAIL VTAIL.n19 0.784983
R234 VDD1.n1 VDD1.t9 78.4679
R235 VDD1.n3 VDD1.t7 78.4676
R236 VDD1.n5 VDD1.n4 75.1073
R237 VDD1.n1 VDD1.n0 72.6347
R238 VDD1.n3 VDD1.n2 72.6346
R239 VDD1.n7 VDD1.n6 72.6345
R240 VDD1.n7 VDD1.n5 53.3737
R241 VDD1 VDD1.n7 2.47033
R242 VDD1.n6 VDD1.t0 2.463
R243 VDD1.n6 VDD1.t8 2.463
R244 VDD1.n0 VDD1.t6 2.463
R245 VDD1.n0 VDD1.t4 2.463
R246 VDD1.n4 VDD1.t1 2.463
R247 VDD1.n4 VDD1.t3 2.463
R248 VDD1.n2 VDD1.t5 2.463
R249 VDD1.n2 VDD1.t2 2.463
R250 VDD1 VDD1.n1 0.901362
R251 VDD1.n5 VDD1.n3 0.787826
R252 B.n764 B.n763 585
R253 B.n765 B.n94 585
R254 B.n767 B.n766 585
R255 B.n768 B.n93 585
R256 B.n770 B.n769 585
R257 B.n771 B.n92 585
R258 B.n773 B.n772 585
R259 B.n774 B.n91 585
R260 B.n776 B.n775 585
R261 B.n777 B.n90 585
R262 B.n779 B.n778 585
R263 B.n780 B.n89 585
R264 B.n782 B.n781 585
R265 B.n783 B.n88 585
R266 B.n785 B.n784 585
R267 B.n786 B.n87 585
R268 B.n788 B.n787 585
R269 B.n789 B.n86 585
R270 B.n791 B.n790 585
R271 B.n792 B.n85 585
R272 B.n794 B.n793 585
R273 B.n795 B.n84 585
R274 B.n797 B.n796 585
R275 B.n798 B.n83 585
R276 B.n800 B.n799 585
R277 B.n801 B.n82 585
R278 B.n803 B.n802 585
R279 B.n804 B.n81 585
R280 B.n806 B.n805 585
R281 B.n807 B.n80 585
R282 B.n809 B.n808 585
R283 B.n810 B.n79 585
R284 B.n812 B.n811 585
R285 B.n813 B.n78 585
R286 B.n815 B.n814 585
R287 B.n816 B.n77 585
R288 B.n818 B.n817 585
R289 B.n819 B.n76 585
R290 B.n821 B.n820 585
R291 B.n822 B.n75 585
R292 B.n824 B.n823 585
R293 B.n825 B.n74 585
R294 B.n827 B.n826 585
R295 B.n828 B.n73 585
R296 B.n830 B.n829 585
R297 B.n832 B.n831 585
R298 B.n833 B.n69 585
R299 B.n835 B.n834 585
R300 B.n836 B.n68 585
R301 B.n838 B.n837 585
R302 B.n839 B.n67 585
R303 B.n841 B.n840 585
R304 B.n842 B.n66 585
R305 B.n844 B.n843 585
R306 B.n845 B.n63 585
R307 B.n848 B.n847 585
R308 B.n849 B.n62 585
R309 B.n851 B.n850 585
R310 B.n852 B.n61 585
R311 B.n854 B.n853 585
R312 B.n855 B.n60 585
R313 B.n857 B.n856 585
R314 B.n858 B.n59 585
R315 B.n860 B.n859 585
R316 B.n861 B.n58 585
R317 B.n863 B.n862 585
R318 B.n864 B.n57 585
R319 B.n866 B.n865 585
R320 B.n867 B.n56 585
R321 B.n869 B.n868 585
R322 B.n870 B.n55 585
R323 B.n872 B.n871 585
R324 B.n873 B.n54 585
R325 B.n875 B.n874 585
R326 B.n876 B.n53 585
R327 B.n878 B.n877 585
R328 B.n879 B.n52 585
R329 B.n881 B.n880 585
R330 B.n882 B.n51 585
R331 B.n884 B.n883 585
R332 B.n885 B.n50 585
R333 B.n887 B.n886 585
R334 B.n888 B.n49 585
R335 B.n890 B.n889 585
R336 B.n891 B.n48 585
R337 B.n893 B.n892 585
R338 B.n894 B.n47 585
R339 B.n896 B.n895 585
R340 B.n897 B.n46 585
R341 B.n899 B.n898 585
R342 B.n900 B.n45 585
R343 B.n902 B.n901 585
R344 B.n903 B.n44 585
R345 B.n905 B.n904 585
R346 B.n906 B.n43 585
R347 B.n908 B.n907 585
R348 B.n909 B.n42 585
R349 B.n911 B.n910 585
R350 B.n912 B.n41 585
R351 B.n914 B.n913 585
R352 B.n762 B.n95 585
R353 B.n761 B.n760 585
R354 B.n759 B.n96 585
R355 B.n758 B.n757 585
R356 B.n756 B.n97 585
R357 B.n755 B.n754 585
R358 B.n753 B.n98 585
R359 B.n752 B.n751 585
R360 B.n750 B.n99 585
R361 B.n749 B.n748 585
R362 B.n747 B.n100 585
R363 B.n746 B.n745 585
R364 B.n744 B.n101 585
R365 B.n743 B.n742 585
R366 B.n741 B.n102 585
R367 B.n740 B.n739 585
R368 B.n738 B.n103 585
R369 B.n737 B.n736 585
R370 B.n735 B.n104 585
R371 B.n734 B.n733 585
R372 B.n732 B.n105 585
R373 B.n731 B.n730 585
R374 B.n729 B.n106 585
R375 B.n728 B.n727 585
R376 B.n726 B.n107 585
R377 B.n725 B.n724 585
R378 B.n723 B.n108 585
R379 B.n722 B.n721 585
R380 B.n720 B.n109 585
R381 B.n719 B.n718 585
R382 B.n717 B.n110 585
R383 B.n716 B.n715 585
R384 B.n714 B.n111 585
R385 B.n713 B.n712 585
R386 B.n711 B.n112 585
R387 B.n710 B.n709 585
R388 B.n708 B.n113 585
R389 B.n707 B.n706 585
R390 B.n705 B.n114 585
R391 B.n704 B.n703 585
R392 B.n702 B.n115 585
R393 B.n701 B.n700 585
R394 B.n699 B.n116 585
R395 B.n698 B.n697 585
R396 B.n696 B.n117 585
R397 B.n695 B.n694 585
R398 B.n693 B.n118 585
R399 B.n692 B.n691 585
R400 B.n690 B.n119 585
R401 B.n689 B.n688 585
R402 B.n687 B.n120 585
R403 B.n686 B.n685 585
R404 B.n684 B.n121 585
R405 B.n683 B.n682 585
R406 B.n681 B.n122 585
R407 B.n680 B.n679 585
R408 B.n678 B.n123 585
R409 B.n677 B.n676 585
R410 B.n675 B.n124 585
R411 B.n674 B.n673 585
R412 B.n672 B.n125 585
R413 B.n671 B.n670 585
R414 B.n669 B.n126 585
R415 B.n668 B.n667 585
R416 B.n666 B.n127 585
R417 B.n665 B.n664 585
R418 B.n663 B.n128 585
R419 B.n662 B.n661 585
R420 B.n660 B.n129 585
R421 B.n659 B.n658 585
R422 B.n657 B.n130 585
R423 B.n656 B.n655 585
R424 B.n654 B.n131 585
R425 B.n653 B.n652 585
R426 B.n651 B.n132 585
R427 B.n650 B.n649 585
R428 B.n648 B.n133 585
R429 B.n647 B.n646 585
R430 B.n645 B.n134 585
R431 B.n644 B.n643 585
R432 B.n642 B.n135 585
R433 B.n641 B.n640 585
R434 B.n639 B.n136 585
R435 B.n638 B.n637 585
R436 B.n636 B.n137 585
R437 B.n635 B.n634 585
R438 B.n633 B.n138 585
R439 B.n632 B.n631 585
R440 B.n630 B.n139 585
R441 B.n629 B.n628 585
R442 B.n627 B.n140 585
R443 B.n626 B.n625 585
R444 B.n624 B.n141 585
R445 B.n623 B.n622 585
R446 B.n621 B.n142 585
R447 B.n620 B.n619 585
R448 B.n618 B.n143 585
R449 B.n617 B.n616 585
R450 B.n615 B.n144 585
R451 B.n614 B.n613 585
R452 B.n612 B.n145 585
R453 B.n611 B.n610 585
R454 B.n609 B.n146 585
R455 B.n608 B.n607 585
R456 B.n606 B.n147 585
R457 B.n605 B.n604 585
R458 B.n603 B.n148 585
R459 B.n602 B.n601 585
R460 B.n600 B.n149 585
R461 B.n599 B.n598 585
R462 B.n597 B.n150 585
R463 B.n596 B.n595 585
R464 B.n594 B.n151 585
R465 B.n593 B.n592 585
R466 B.n591 B.n152 585
R467 B.n590 B.n589 585
R468 B.n588 B.n153 585
R469 B.n587 B.n586 585
R470 B.n585 B.n154 585
R471 B.n584 B.n583 585
R472 B.n582 B.n155 585
R473 B.n581 B.n580 585
R474 B.n579 B.n156 585
R475 B.n578 B.n577 585
R476 B.n576 B.n157 585
R477 B.n575 B.n574 585
R478 B.n573 B.n158 585
R479 B.n572 B.n571 585
R480 B.n570 B.n159 585
R481 B.n569 B.n568 585
R482 B.n567 B.n160 585
R483 B.n566 B.n565 585
R484 B.n564 B.n161 585
R485 B.n563 B.n562 585
R486 B.n561 B.n162 585
R487 B.n560 B.n559 585
R488 B.n558 B.n163 585
R489 B.n557 B.n556 585
R490 B.n555 B.n164 585
R491 B.n554 B.n553 585
R492 B.n552 B.n165 585
R493 B.n551 B.n550 585
R494 B.n549 B.n166 585
R495 B.n548 B.n547 585
R496 B.n546 B.n167 585
R497 B.n545 B.n544 585
R498 B.n543 B.n168 585
R499 B.n542 B.n541 585
R500 B.n540 B.n169 585
R501 B.n539 B.n538 585
R502 B.n537 B.n170 585
R503 B.n536 B.n535 585
R504 B.n534 B.n171 585
R505 B.n533 B.n532 585
R506 B.n531 B.n172 585
R507 B.n380 B.n379 585
R508 B.n381 B.n226 585
R509 B.n383 B.n382 585
R510 B.n384 B.n225 585
R511 B.n386 B.n385 585
R512 B.n387 B.n224 585
R513 B.n389 B.n388 585
R514 B.n390 B.n223 585
R515 B.n392 B.n391 585
R516 B.n393 B.n222 585
R517 B.n395 B.n394 585
R518 B.n396 B.n221 585
R519 B.n398 B.n397 585
R520 B.n399 B.n220 585
R521 B.n401 B.n400 585
R522 B.n402 B.n219 585
R523 B.n404 B.n403 585
R524 B.n405 B.n218 585
R525 B.n407 B.n406 585
R526 B.n408 B.n217 585
R527 B.n410 B.n409 585
R528 B.n411 B.n216 585
R529 B.n413 B.n412 585
R530 B.n414 B.n215 585
R531 B.n416 B.n415 585
R532 B.n417 B.n214 585
R533 B.n419 B.n418 585
R534 B.n420 B.n213 585
R535 B.n422 B.n421 585
R536 B.n423 B.n212 585
R537 B.n425 B.n424 585
R538 B.n426 B.n211 585
R539 B.n428 B.n427 585
R540 B.n429 B.n210 585
R541 B.n431 B.n430 585
R542 B.n432 B.n209 585
R543 B.n434 B.n433 585
R544 B.n435 B.n208 585
R545 B.n437 B.n436 585
R546 B.n438 B.n207 585
R547 B.n440 B.n439 585
R548 B.n441 B.n206 585
R549 B.n443 B.n442 585
R550 B.n444 B.n205 585
R551 B.n446 B.n445 585
R552 B.n448 B.n447 585
R553 B.n449 B.n201 585
R554 B.n451 B.n450 585
R555 B.n452 B.n200 585
R556 B.n454 B.n453 585
R557 B.n455 B.n199 585
R558 B.n457 B.n456 585
R559 B.n458 B.n198 585
R560 B.n460 B.n459 585
R561 B.n461 B.n195 585
R562 B.n464 B.n463 585
R563 B.n465 B.n194 585
R564 B.n467 B.n466 585
R565 B.n468 B.n193 585
R566 B.n470 B.n469 585
R567 B.n471 B.n192 585
R568 B.n473 B.n472 585
R569 B.n474 B.n191 585
R570 B.n476 B.n475 585
R571 B.n477 B.n190 585
R572 B.n479 B.n478 585
R573 B.n480 B.n189 585
R574 B.n482 B.n481 585
R575 B.n483 B.n188 585
R576 B.n485 B.n484 585
R577 B.n486 B.n187 585
R578 B.n488 B.n487 585
R579 B.n489 B.n186 585
R580 B.n491 B.n490 585
R581 B.n492 B.n185 585
R582 B.n494 B.n493 585
R583 B.n495 B.n184 585
R584 B.n497 B.n496 585
R585 B.n498 B.n183 585
R586 B.n500 B.n499 585
R587 B.n501 B.n182 585
R588 B.n503 B.n502 585
R589 B.n504 B.n181 585
R590 B.n506 B.n505 585
R591 B.n507 B.n180 585
R592 B.n509 B.n508 585
R593 B.n510 B.n179 585
R594 B.n512 B.n511 585
R595 B.n513 B.n178 585
R596 B.n515 B.n514 585
R597 B.n516 B.n177 585
R598 B.n518 B.n517 585
R599 B.n519 B.n176 585
R600 B.n521 B.n520 585
R601 B.n522 B.n175 585
R602 B.n524 B.n523 585
R603 B.n525 B.n174 585
R604 B.n527 B.n526 585
R605 B.n528 B.n173 585
R606 B.n530 B.n529 585
R607 B.n378 B.n227 585
R608 B.n377 B.n376 585
R609 B.n375 B.n228 585
R610 B.n374 B.n373 585
R611 B.n372 B.n229 585
R612 B.n371 B.n370 585
R613 B.n369 B.n230 585
R614 B.n368 B.n367 585
R615 B.n366 B.n231 585
R616 B.n365 B.n364 585
R617 B.n363 B.n232 585
R618 B.n362 B.n361 585
R619 B.n360 B.n233 585
R620 B.n359 B.n358 585
R621 B.n357 B.n234 585
R622 B.n356 B.n355 585
R623 B.n354 B.n235 585
R624 B.n353 B.n352 585
R625 B.n351 B.n236 585
R626 B.n350 B.n349 585
R627 B.n348 B.n237 585
R628 B.n347 B.n346 585
R629 B.n345 B.n238 585
R630 B.n344 B.n343 585
R631 B.n342 B.n239 585
R632 B.n341 B.n340 585
R633 B.n339 B.n240 585
R634 B.n338 B.n337 585
R635 B.n336 B.n241 585
R636 B.n335 B.n334 585
R637 B.n333 B.n242 585
R638 B.n332 B.n331 585
R639 B.n330 B.n243 585
R640 B.n329 B.n328 585
R641 B.n327 B.n244 585
R642 B.n326 B.n325 585
R643 B.n324 B.n245 585
R644 B.n323 B.n322 585
R645 B.n321 B.n246 585
R646 B.n320 B.n319 585
R647 B.n318 B.n247 585
R648 B.n317 B.n316 585
R649 B.n315 B.n248 585
R650 B.n314 B.n313 585
R651 B.n312 B.n249 585
R652 B.n311 B.n310 585
R653 B.n309 B.n250 585
R654 B.n308 B.n307 585
R655 B.n306 B.n251 585
R656 B.n305 B.n304 585
R657 B.n303 B.n252 585
R658 B.n302 B.n301 585
R659 B.n300 B.n253 585
R660 B.n299 B.n298 585
R661 B.n297 B.n254 585
R662 B.n296 B.n295 585
R663 B.n294 B.n255 585
R664 B.n293 B.n292 585
R665 B.n291 B.n256 585
R666 B.n290 B.n289 585
R667 B.n288 B.n257 585
R668 B.n287 B.n286 585
R669 B.n285 B.n258 585
R670 B.n284 B.n283 585
R671 B.n282 B.n259 585
R672 B.n281 B.n280 585
R673 B.n279 B.n260 585
R674 B.n278 B.n277 585
R675 B.n276 B.n261 585
R676 B.n275 B.n274 585
R677 B.n273 B.n262 585
R678 B.n272 B.n271 585
R679 B.n270 B.n263 585
R680 B.n269 B.n268 585
R681 B.n267 B.n264 585
R682 B.n266 B.n265 585
R683 B.n2 B.n0 585
R684 B.n1029 B.n1 585
R685 B.n1028 B.n1027 585
R686 B.n1026 B.n3 585
R687 B.n1025 B.n1024 585
R688 B.n1023 B.n4 585
R689 B.n1022 B.n1021 585
R690 B.n1020 B.n5 585
R691 B.n1019 B.n1018 585
R692 B.n1017 B.n6 585
R693 B.n1016 B.n1015 585
R694 B.n1014 B.n7 585
R695 B.n1013 B.n1012 585
R696 B.n1011 B.n8 585
R697 B.n1010 B.n1009 585
R698 B.n1008 B.n9 585
R699 B.n1007 B.n1006 585
R700 B.n1005 B.n10 585
R701 B.n1004 B.n1003 585
R702 B.n1002 B.n11 585
R703 B.n1001 B.n1000 585
R704 B.n999 B.n12 585
R705 B.n998 B.n997 585
R706 B.n996 B.n13 585
R707 B.n995 B.n994 585
R708 B.n993 B.n14 585
R709 B.n992 B.n991 585
R710 B.n990 B.n15 585
R711 B.n989 B.n988 585
R712 B.n987 B.n16 585
R713 B.n986 B.n985 585
R714 B.n984 B.n17 585
R715 B.n983 B.n982 585
R716 B.n981 B.n18 585
R717 B.n980 B.n979 585
R718 B.n978 B.n19 585
R719 B.n977 B.n976 585
R720 B.n975 B.n20 585
R721 B.n974 B.n973 585
R722 B.n972 B.n21 585
R723 B.n971 B.n970 585
R724 B.n969 B.n22 585
R725 B.n968 B.n967 585
R726 B.n966 B.n23 585
R727 B.n965 B.n964 585
R728 B.n963 B.n24 585
R729 B.n962 B.n961 585
R730 B.n960 B.n25 585
R731 B.n959 B.n958 585
R732 B.n957 B.n26 585
R733 B.n956 B.n955 585
R734 B.n954 B.n27 585
R735 B.n953 B.n952 585
R736 B.n951 B.n28 585
R737 B.n950 B.n949 585
R738 B.n948 B.n29 585
R739 B.n947 B.n946 585
R740 B.n945 B.n30 585
R741 B.n944 B.n943 585
R742 B.n942 B.n31 585
R743 B.n941 B.n940 585
R744 B.n939 B.n32 585
R745 B.n938 B.n937 585
R746 B.n936 B.n33 585
R747 B.n935 B.n934 585
R748 B.n933 B.n34 585
R749 B.n932 B.n931 585
R750 B.n930 B.n35 585
R751 B.n929 B.n928 585
R752 B.n927 B.n36 585
R753 B.n926 B.n925 585
R754 B.n924 B.n37 585
R755 B.n923 B.n922 585
R756 B.n921 B.n38 585
R757 B.n920 B.n919 585
R758 B.n918 B.n39 585
R759 B.n917 B.n916 585
R760 B.n915 B.n40 585
R761 B.n1031 B.n1030 585
R762 B.n380 B.n227 506.916
R763 B.n915 B.n914 506.916
R764 B.n531 B.n530 506.916
R765 B.n764 B.n95 506.916
R766 B.n196 B.t6 298.024
R767 B.n202 B.t3 298.024
R768 B.n64 B.t0 298.024
R769 B.n70 B.t9 298.024
R770 B.n196 B.t8 188.117
R771 B.n70 B.t10 188.117
R772 B.n202 B.t5 188.101
R773 B.n64 B.t1 188.101
R774 B.n376 B.n227 163.367
R775 B.n376 B.n375 163.367
R776 B.n375 B.n374 163.367
R777 B.n374 B.n229 163.367
R778 B.n370 B.n229 163.367
R779 B.n370 B.n369 163.367
R780 B.n369 B.n368 163.367
R781 B.n368 B.n231 163.367
R782 B.n364 B.n231 163.367
R783 B.n364 B.n363 163.367
R784 B.n363 B.n362 163.367
R785 B.n362 B.n233 163.367
R786 B.n358 B.n233 163.367
R787 B.n358 B.n357 163.367
R788 B.n357 B.n356 163.367
R789 B.n356 B.n235 163.367
R790 B.n352 B.n235 163.367
R791 B.n352 B.n351 163.367
R792 B.n351 B.n350 163.367
R793 B.n350 B.n237 163.367
R794 B.n346 B.n237 163.367
R795 B.n346 B.n345 163.367
R796 B.n345 B.n344 163.367
R797 B.n344 B.n239 163.367
R798 B.n340 B.n239 163.367
R799 B.n340 B.n339 163.367
R800 B.n339 B.n338 163.367
R801 B.n338 B.n241 163.367
R802 B.n334 B.n241 163.367
R803 B.n334 B.n333 163.367
R804 B.n333 B.n332 163.367
R805 B.n332 B.n243 163.367
R806 B.n328 B.n243 163.367
R807 B.n328 B.n327 163.367
R808 B.n327 B.n326 163.367
R809 B.n326 B.n245 163.367
R810 B.n322 B.n245 163.367
R811 B.n322 B.n321 163.367
R812 B.n321 B.n320 163.367
R813 B.n320 B.n247 163.367
R814 B.n316 B.n247 163.367
R815 B.n316 B.n315 163.367
R816 B.n315 B.n314 163.367
R817 B.n314 B.n249 163.367
R818 B.n310 B.n249 163.367
R819 B.n310 B.n309 163.367
R820 B.n309 B.n308 163.367
R821 B.n308 B.n251 163.367
R822 B.n304 B.n251 163.367
R823 B.n304 B.n303 163.367
R824 B.n303 B.n302 163.367
R825 B.n302 B.n253 163.367
R826 B.n298 B.n253 163.367
R827 B.n298 B.n297 163.367
R828 B.n297 B.n296 163.367
R829 B.n296 B.n255 163.367
R830 B.n292 B.n255 163.367
R831 B.n292 B.n291 163.367
R832 B.n291 B.n290 163.367
R833 B.n290 B.n257 163.367
R834 B.n286 B.n257 163.367
R835 B.n286 B.n285 163.367
R836 B.n285 B.n284 163.367
R837 B.n284 B.n259 163.367
R838 B.n280 B.n259 163.367
R839 B.n280 B.n279 163.367
R840 B.n279 B.n278 163.367
R841 B.n278 B.n261 163.367
R842 B.n274 B.n261 163.367
R843 B.n274 B.n273 163.367
R844 B.n273 B.n272 163.367
R845 B.n272 B.n263 163.367
R846 B.n268 B.n263 163.367
R847 B.n268 B.n267 163.367
R848 B.n267 B.n266 163.367
R849 B.n266 B.n2 163.367
R850 B.n1030 B.n2 163.367
R851 B.n1030 B.n1029 163.367
R852 B.n1029 B.n1028 163.367
R853 B.n1028 B.n3 163.367
R854 B.n1024 B.n3 163.367
R855 B.n1024 B.n1023 163.367
R856 B.n1023 B.n1022 163.367
R857 B.n1022 B.n5 163.367
R858 B.n1018 B.n5 163.367
R859 B.n1018 B.n1017 163.367
R860 B.n1017 B.n1016 163.367
R861 B.n1016 B.n7 163.367
R862 B.n1012 B.n7 163.367
R863 B.n1012 B.n1011 163.367
R864 B.n1011 B.n1010 163.367
R865 B.n1010 B.n9 163.367
R866 B.n1006 B.n9 163.367
R867 B.n1006 B.n1005 163.367
R868 B.n1005 B.n1004 163.367
R869 B.n1004 B.n11 163.367
R870 B.n1000 B.n11 163.367
R871 B.n1000 B.n999 163.367
R872 B.n999 B.n998 163.367
R873 B.n998 B.n13 163.367
R874 B.n994 B.n13 163.367
R875 B.n994 B.n993 163.367
R876 B.n993 B.n992 163.367
R877 B.n992 B.n15 163.367
R878 B.n988 B.n15 163.367
R879 B.n988 B.n987 163.367
R880 B.n987 B.n986 163.367
R881 B.n986 B.n17 163.367
R882 B.n982 B.n17 163.367
R883 B.n982 B.n981 163.367
R884 B.n981 B.n980 163.367
R885 B.n980 B.n19 163.367
R886 B.n976 B.n19 163.367
R887 B.n976 B.n975 163.367
R888 B.n975 B.n974 163.367
R889 B.n974 B.n21 163.367
R890 B.n970 B.n21 163.367
R891 B.n970 B.n969 163.367
R892 B.n969 B.n968 163.367
R893 B.n968 B.n23 163.367
R894 B.n964 B.n23 163.367
R895 B.n964 B.n963 163.367
R896 B.n963 B.n962 163.367
R897 B.n962 B.n25 163.367
R898 B.n958 B.n25 163.367
R899 B.n958 B.n957 163.367
R900 B.n957 B.n956 163.367
R901 B.n956 B.n27 163.367
R902 B.n952 B.n27 163.367
R903 B.n952 B.n951 163.367
R904 B.n951 B.n950 163.367
R905 B.n950 B.n29 163.367
R906 B.n946 B.n29 163.367
R907 B.n946 B.n945 163.367
R908 B.n945 B.n944 163.367
R909 B.n944 B.n31 163.367
R910 B.n940 B.n31 163.367
R911 B.n940 B.n939 163.367
R912 B.n939 B.n938 163.367
R913 B.n938 B.n33 163.367
R914 B.n934 B.n33 163.367
R915 B.n934 B.n933 163.367
R916 B.n933 B.n932 163.367
R917 B.n932 B.n35 163.367
R918 B.n928 B.n35 163.367
R919 B.n928 B.n927 163.367
R920 B.n927 B.n926 163.367
R921 B.n926 B.n37 163.367
R922 B.n922 B.n37 163.367
R923 B.n922 B.n921 163.367
R924 B.n921 B.n920 163.367
R925 B.n920 B.n39 163.367
R926 B.n916 B.n39 163.367
R927 B.n916 B.n915 163.367
R928 B.n381 B.n380 163.367
R929 B.n382 B.n381 163.367
R930 B.n382 B.n225 163.367
R931 B.n386 B.n225 163.367
R932 B.n387 B.n386 163.367
R933 B.n388 B.n387 163.367
R934 B.n388 B.n223 163.367
R935 B.n392 B.n223 163.367
R936 B.n393 B.n392 163.367
R937 B.n394 B.n393 163.367
R938 B.n394 B.n221 163.367
R939 B.n398 B.n221 163.367
R940 B.n399 B.n398 163.367
R941 B.n400 B.n399 163.367
R942 B.n400 B.n219 163.367
R943 B.n404 B.n219 163.367
R944 B.n405 B.n404 163.367
R945 B.n406 B.n405 163.367
R946 B.n406 B.n217 163.367
R947 B.n410 B.n217 163.367
R948 B.n411 B.n410 163.367
R949 B.n412 B.n411 163.367
R950 B.n412 B.n215 163.367
R951 B.n416 B.n215 163.367
R952 B.n417 B.n416 163.367
R953 B.n418 B.n417 163.367
R954 B.n418 B.n213 163.367
R955 B.n422 B.n213 163.367
R956 B.n423 B.n422 163.367
R957 B.n424 B.n423 163.367
R958 B.n424 B.n211 163.367
R959 B.n428 B.n211 163.367
R960 B.n429 B.n428 163.367
R961 B.n430 B.n429 163.367
R962 B.n430 B.n209 163.367
R963 B.n434 B.n209 163.367
R964 B.n435 B.n434 163.367
R965 B.n436 B.n435 163.367
R966 B.n436 B.n207 163.367
R967 B.n440 B.n207 163.367
R968 B.n441 B.n440 163.367
R969 B.n442 B.n441 163.367
R970 B.n442 B.n205 163.367
R971 B.n446 B.n205 163.367
R972 B.n447 B.n446 163.367
R973 B.n447 B.n201 163.367
R974 B.n451 B.n201 163.367
R975 B.n452 B.n451 163.367
R976 B.n453 B.n452 163.367
R977 B.n453 B.n199 163.367
R978 B.n457 B.n199 163.367
R979 B.n458 B.n457 163.367
R980 B.n459 B.n458 163.367
R981 B.n459 B.n195 163.367
R982 B.n464 B.n195 163.367
R983 B.n465 B.n464 163.367
R984 B.n466 B.n465 163.367
R985 B.n466 B.n193 163.367
R986 B.n470 B.n193 163.367
R987 B.n471 B.n470 163.367
R988 B.n472 B.n471 163.367
R989 B.n472 B.n191 163.367
R990 B.n476 B.n191 163.367
R991 B.n477 B.n476 163.367
R992 B.n478 B.n477 163.367
R993 B.n478 B.n189 163.367
R994 B.n482 B.n189 163.367
R995 B.n483 B.n482 163.367
R996 B.n484 B.n483 163.367
R997 B.n484 B.n187 163.367
R998 B.n488 B.n187 163.367
R999 B.n489 B.n488 163.367
R1000 B.n490 B.n489 163.367
R1001 B.n490 B.n185 163.367
R1002 B.n494 B.n185 163.367
R1003 B.n495 B.n494 163.367
R1004 B.n496 B.n495 163.367
R1005 B.n496 B.n183 163.367
R1006 B.n500 B.n183 163.367
R1007 B.n501 B.n500 163.367
R1008 B.n502 B.n501 163.367
R1009 B.n502 B.n181 163.367
R1010 B.n506 B.n181 163.367
R1011 B.n507 B.n506 163.367
R1012 B.n508 B.n507 163.367
R1013 B.n508 B.n179 163.367
R1014 B.n512 B.n179 163.367
R1015 B.n513 B.n512 163.367
R1016 B.n514 B.n513 163.367
R1017 B.n514 B.n177 163.367
R1018 B.n518 B.n177 163.367
R1019 B.n519 B.n518 163.367
R1020 B.n520 B.n519 163.367
R1021 B.n520 B.n175 163.367
R1022 B.n524 B.n175 163.367
R1023 B.n525 B.n524 163.367
R1024 B.n526 B.n525 163.367
R1025 B.n526 B.n173 163.367
R1026 B.n530 B.n173 163.367
R1027 B.n532 B.n531 163.367
R1028 B.n532 B.n171 163.367
R1029 B.n536 B.n171 163.367
R1030 B.n537 B.n536 163.367
R1031 B.n538 B.n537 163.367
R1032 B.n538 B.n169 163.367
R1033 B.n542 B.n169 163.367
R1034 B.n543 B.n542 163.367
R1035 B.n544 B.n543 163.367
R1036 B.n544 B.n167 163.367
R1037 B.n548 B.n167 163.367
R1038 B.n549 B.n548 163.367
R1039 B.n550 B.n549 163.367
R1040 B.n550 B.n165 163.367
R1041 B.n554 B.n165 163.367
R1042 B.n555 B.n554 163.367
R1043 B.n556 B.n555 163.367
R1044 B.n556 B.n163 163.367
R1045 B.n560 B.n163 163.367
R1046 B.n561 B.n560 163.367
R1047 B.n562 B.n561 163.367
R1048 B.n562 B.n161 163.367
R1049 B.n566 B.n161 163.367
R1050 B.n567 B.n566 163.367
R1051 B.n568 B.n567 163.367
R1052 B.n568 B.n159 163.367
R1053 B.n572 B.n159 163.367
R1054 B.n573 B.n572 163.367
R1055 B.n574 B.n573 163.367
R1056 B.n574 B.n157 163.367
R1057 B.n578 B.n157 163.367
R1058 B.n579 B.n578 163.367
R1059 B.n580 B.n579 163.367
R1060 B.n580 B.n155 163.367
R1061 B.n584 B.n155 163.367
R1062 B.n585 B.n584 163.367
R1063 B.n586 B.n585 163.367
R1064 B.n586 B.n153 163.367
R1065 B.n590 B.n153 163.367
R1066 B.n591 B.n590 163.367
R1067 B.n592 B.n591 163.367
R1068 B.n592 B.n151 163.367
R1069 B.n596 B.n151 163.367
R1070 B.n597 B.n596 163.367
R1071 B.n598 B.n597 163.367
R1072 B.n598 B.n149 163.367
R1073 B.n602 B.n149 163.367
R1074 B.n603 B.n602 163.367
R1075 B.n604 B.n603 163.367
R1076 B.n604 B.n147 163.367
R1077 B.n608 B.n147 163.367
R1078 B.n609 B.n608 163.367
R1079 B.n610 B.n609 163.367
R1080 B.n610 B.n145 163.367
R1081 B.n614 B.n145 163.367
R1082 B.n615 B.n614 163.367
R1083 B.n616 B.n615 163.367
R1084 B.n616 B.n143 163.367
R1085 B.n620 B.n143 163.367
R1086 B.n621 B.n620 163.367
R1087 B.n622 B.n621 163.367
R1088 B.n622 B.n141 163.367
R1089 B.n626 B.n141 163.367
R1090 B.n627 B.n626 163.367
R1091 B.n628 B.n627 163.367
R1092 B.n628 B.n139 163.367
R1093 B.n632 B.n139 163.367
R1094 B.n633 B.n632 163.367
R1095 B.n634 B.n633 163.367
R1096 B.n634 B.n137 163.367
R1097 B.n638 B.n137 163.367
R1098 B.n639 B.n638 163.367
R1099 B.n640 B.n639 163.367
R1100 B.n640 B.n135 163.367
R1101 B.n644 B.n135 163.367
R1102 B.n645 B.n644 163.367
R1103 B.n646 B.n645 163.367
R1104 B.n646 B.n133 163.367
R1105 B.n650 B.n133 163.367
R1106 B.n651 B.n650 163.367
R1107 B.n652 B.n651 163.367
R1108 B.n652 B.n131 163.367
R1109 B.n656 B.n131 163.367
R1110 B.n657 B.n656 163.367
R1111 B.n658 B.n657 163.367
R1112 B.n658 B.n129 163.367
R1113 B.n662 B.n129 163.367
R1114 B.n663 B.n662 163.367
R1115 B.n664 B.n663 163.367
R1116 B.n664 B.n127 163.367
R1117 B.n668 B.n127 163.367
R1118 B.n669 B.n668 163.367
R1119 B.n670 B.n669 163.367
R1120 B.n670 B.n125 163.367
R1121 B.n674 B.n125 163.367
R1122 B.n675 B.n674 163.367
R1123 B.n676 B.n675 163.367
R1124 B.n676 B.n123 163.367
R1125 B.n680 B.n123 163.367
R1126 B.n681 B.n680 163.367
R1127 B.n682 B.n681 163.367
R1128 B.n682 B.n121 163.367
R1129 B.n686 B.n121 163.367
R1130 B.n687 B.n686 163.367
R1131 B.n688 B.n687 163.367
R1132 B.n688 B.n119 163.367
R1133 B.n692 B.n119 163.367
R1134 B.n693 B.n692 163.367
R1135 B.n694 B.n693 163.367
R1136 B.n694 B.n117 163.367
R1137 B.n698 B.n117 163.367
R1138 B.n699 B.n698 163.367
R1139 B.n700 B.n699 163.367
R1140 B.n700 B.n115 163.367
R1141 B.n704 B.n115 163.367
R1142 B.n705 B.n704 163.367
R1143 B.n706 B.n705 163.367
R1144 B.n706 B.n113 163.367
R1145 B.n710 B.n113 163.367
R1146 B.n711 B.n710 163.367
R1147 B.n712 B.n711 163.367
R1148 B.n712 B.n111 163.367
R1149 B.n716 B.n111 163.367
R1150 B.n717 B.n716 163.367
R1151 B.n718 B.n717 163.367
R1152 B.n718 B.n109 163.367
R1153 B.n722 B.n109 163.367
R1154 B.n723 B.n722 163.367
R1155 B.n724 B.n723 163.367
R1156 B.n724 B.n107 163.367
R1157 B.n728 B.n107 163.367
R1158 B.n729 B.n728 163.367
R1159 B.n730 B.n729 163.367
R1160 B.n730 B.n105 163.367
R1161 B.n734 B.n105 163.367
R1162 B.n735 B.n734 163.367
R1163 B.n736 B.n735 163.367
R1164 B.n736 B.n103 163.367
R1165 B.n740 B.n103 163.367
R1166 B.n741 B.n740 163.367
R1167 B.n742 B.n741 163.367
R1168 B.n742 B.n101 163.367
R1169 B.n746 B.n101 163.367
R1170 B.n747 B.n746 163.367
R1171 B.n748 B.n747 163.367
R1172 B.n748 B.n99 163.367
R1173 B.n752 B.n99 163.367
R1174 B.n753 B.n752 163.367
R1175 B.n754 B.n753 163.367
R1176 B.n754 B.n97 163.367
R1177 B.n758 B.n97 163.367
R1178 B.n759 B.n758 163.367
R1179 B.n760 B.n759 163.367
R1180 B.n760 B.n95 163.367
R1181 B.n914 B.n41 163.367
R1182 B.n910 B.n41 163.367
R1183 B.n910 B.n909 163.367
R1184 B.n909 B.n908 163.367
R1185 B.n908 B.n43 163.367
R1186 B.n904 B.n43 163.367
R1187 B.n904 B.n903 163.367
R1188 B.n903 B.n902 163.367
R1189 B.n902 B.n45 163.367
R1190 B.n898 B.n45 163.367
R1191 B.n898 B.n897 163.367
R1192 B.n897 B.n896 163.367
R1193 B.n896 B.n47 163.367
R1194 B.n892 B.n47 163.367
R1195 B.n892 B.n891 163.367
R1196 B.n891 B.n890 163.367
R1197 B.n890 B.n49 163.367
R1198 B.n886 B.n49 163.367
R1199 B.n886 B.n885 163.367
R1200 B.n885 B.n884 163.367
R1201 B.n884 B.n51 163.367
R1202 B.n880 B.n51 163.367
R1203 B.n880 B.n879 163.367
R1204 B.n879 B.n878 163.367
R1205 B.n878 B.n53 163.367
R1206 B.n874 B.n53 163.367
R1207 B.n874 B.n873 163.367
R1208 B.n873 B.n872 163.367
R1209 B.n872 B.n55 163.367
R1210 B.n868 B.n55 163.367
R1211 B.n868 B.n867 163.367
R1212 B.n867 B.n866 163.367
R1213 B.n866 B.n57 163.367
R1214 B.n862 B.n57 163.367
R1215 B.n862 B.n861 163.367
R1216 B.n861 B.n860 163.367
R1217 B.n860 B.n59 163.367
R1218 B.n856 B.n59 163.367
R1219 B.n856 B.n855 163.367
R1220 B.n855 B.n854 163.367
R1221 B.n854 B.n61 163.367
R1222 B.n850 B.n61 163.367
R1223 B.n850 B.n849 163.367
R1224 B.n849 B.n848 163.367
R1225 B.n848 B.n63 163.367
R1226 B.n843 B.n63 163.367
R1227 B.n843 B.n842 163.367
R1228 B.n842 B.n841 163.367
R1229 B.n841 B.n67 163.367
R1230 B.n837 B.n67 163.367
R1231 B.n837 B.n836 163.367
R1232 B.n836 B.n835 163.367
R1233 B.n835 B.n69 163.367
R1234 B.n831 B.n69 163.367
R1235 B.n831 B.n830 163.367
R1236 B.n830 B.n73 163.367
R1237 B.n826 B.n73 163.367
R1238 B.n826 B.n825 163.367
R1239 B.n825 B.n824 163.367
R1240 B.n824 B.n75 163.367
R1241 B.n820 B.n75 163.367
R1242 B.n820 B.n819 163.367
R1243 B.n819 B.n818 163.367
R1244 B.n818 B.n77 163.367
R1245 B.n814 B.n77 163.367
R1246 B.n814 B.n813 163.367
R1247 B.n813 B.n812 163.367
R1248 B.n812 B.n79 163.367
R1249 B.n808 B.n79 163.367
R1250 B.n808 B.n807 163.367
R1251 B.n807 B.n806 163.367
R1252 B.n806 B.n81 163.367
R1253 B.n802 B.n81 163.367
R1254 B.n802 B.n801 163.367
R1255 B.n801 B.n800 163.367
R1256 B.n800 B.n83 163.367
R1257 B.n796 B.n83 163.367
R1258 B.n796 B.n795 163.367
R1259 B.n795 B.n794 163.367
R1260 B.n794 B.n85 163.367
R1261 B.n790 B.n85 163.367
R1262 B.n790 B.n789 163.367
R1263 B.n789 B.n788 163.367
R1264 B.n788 B.n87 163.367
R1265 B.n784 B.n87 163.367
R1266 B.n784 B.n783 163.367
R1267 B.n783 B.n782 163.367
R1268 B.n782 B.n89 163.367
R1269 B.n778 B.n89 163.367
R1270 B.n778 B.n777 163.367
R1271 B.n777 B.n776 163.367
R1272 B.n776 B.n91 163.367
R1273 B.n772 B.n91 163.367
R1274 B.n772 B.n771 163.367
R1275 B.n771 B.n770 163.367
R1276 B.n770 B.n93 163.367
R1277 B.n766 B.n93 163.367
R1278 B.n766 B.n765 163.367
R1279 B.n765 B.n764 163.367
R1280 B.n197 B.t7 112.287
R1281 B.n71 B.t11 112.287
R1282 B.n203 B.t4 112.27
R1283 B.n65 B.t2 112.27
R1284 B.n197 B.n196 75.8308
R1285 B.n203 B.n202 75.8308
R1286 B.n65 B.n64 75.8308
R1287 B.n71 B.n70 75.8308
R1288 B.n462 B.n197 59.5399
R1289 B.n204 B.n203 59.5399
R1290 B.n846 B.n65 59.5399
R1291 B.n72 B.n71 59.5399
R1292 B.n913 B.n40 32.9371
R1293 B.n763 B.n762 32.9371
R1294 B.n529 B.n172 32.9371
R1295 B.n379 B.n378 32.9371
R1296 B B.n1031 18.0485
R1297 B.n913 B.n912 10.6151
R1298 B.n912 B.n911 10.6151
R1299 B.n911 B.n42 10.6151
R1300 B.n907 B.n42 10.6151
R1301 B.n907 B.n906 10.6151
R1302 B.n906 B.n905 10.6151
R1303 B.n905 B.n44 10.6151
R1304 B.n901 B.n44 10.6151
R1305 B.n901 B.n900 10.6151
R1306 B.n900 B.n899 10.6151
R1307 B.n899 B.n46 10.6151
R1308 B.n895 B.n46 10.6151
R1309 B.n895 B.n894 10.6151
R1310 B.n894 B.n893 10.6151
R1311 B.n893 B.n48 10.6151
R1312 B.n889 B.n48 10.6151
R1313 B.n889 B.n888 10.6151
R1314 B.n888 B.n887 10.6151
R1315 B.n887 B.n50 10.6151
R1316 B.n883 B.n50 10.6151
R1317 B.n883 B.n882 10.6151
R1318 B.n882 B.n881 10.6151
R1319 B.n881 B.n52 10.6151
R1320 B.n877 B.n52 10.6151
R1321 B.n877 B.n876 10.6151
R1322 B.n876 B.n875 10.6151
R1323 B.n875 B.n54 10.6151
R1324 B.n871 B.n54 10.6151
R1325 B.n871 B.n870 10.6151
R1326 B.n870 B.n869 10.6151
R1327 B.n869 B.n56 10.6151
R1328 B.n865 B.n56 10.6151
R1329 B.n865 B.n864 10.6151
R1330 B.n864 B.n863 10.6151
R1331 B.n863 B.n58 10.6151
R1332 B.n859 B.n58 10.6151
R1333 B.n859 B.n858 10.6151
R1334 B.n858 B.n857 10.6151
R1335 B.n857 B.n60 10.6151
R1336 B.n853 B.n60 10.6151
R1337 B.n853 B.n852 10.6151
R1338 B.n852 B.n851 10.6151
R1339 B.n851 B.n62 10.6151
R1340 B.n847 B.n62 10.6151
R1341 B.n845 B.n844 10.6151
R1342 B.n844 B.n66 10.6151
R1343 B.n840 B.n66 10.6151
R1344 B.n840 B.n839 10.6151
R1345 B.n839 B.n838 10.6151
R1346 B.n838 B.n68 10.6151
R1347 B.n834 B.n68 10.6151
R1348 B.n834 B.n833 10.6151
R1349 B.n833 B.n832 10.6151
R1350 B.n829 B.n828 10.6151
R1351 B.n828 B.n827 10.6151
R1352 B.n827 B.n74 10.6151
R1353 B.n823 B.n74 10.6151
R1354 B.n823 B.n822 10.6151
R1355 B.n822 B.n821 10.6151
R1356 B.n821 B.n76 10.6151
R1357 B.n817 B.n76 10.6151
R1358 B.n817 B.n816 10.6151
R1359 B.n816 B.n815 10.6151
R1360 B.n815 B.n78 10.6151
R1361 B.n811 B.n78 10.6151
R1362 B.n811 B.n810 10.6151
R1363 B.n810 B.n809 10.6151
R1364 B.n809 B.n80 10.6151
R1365 B.n805 B.n80 10.6151
R1366 B.n805 B.n804 10.6151
R1367 B.n804 B.n803 10.6151
R1368 B.n803 B.n82 10.6151
R1369 B.n799 B.n82 10.6151
R1370 B.n799 B.n798 10.6151
R1371 B.n798 B.n797 10.6151
R1372 B.n797 B.n84 10.6151
R1373 B.n793 B.n84 10.6151
R1374 B.n793 B.n792 10.6151
R1375 B.n792 B.n791 10.6151
R1376 B.n791 B.n86 10.6151
R1377 B.n787 B.n86 10.6151
R1378 B.n787 B.n786 10.6151
R1379 B.n786 B.n785 10.6151
R1380 B.n785 B.n88 10.6151
R1381 B.n781 B.n88 10.6151
R1382 B.n781 B.n780 10.6151
R1383 B.n780 B.n779 10.6151
R1384 B.n779 B.n90 10.6151
R1385 B.n775 B.n90 10.6151
R1386 B.n775 B.n774 10.6151
R1387 B.n774 B.n773 10.6151
R1388 B.n773 B.n92 10.6151
R1389 B.n769 B.n92 10.6151
R1390 B.n769 B.n768 10.6151
R1391 B.n768 B.n767 10.6151
R1392 B.n767 B.n94 10.6151
R1393 B.n763 B.n94 10.6151
R1394 B.n533 B.n172 10.6151
R1395 B.n534 B.n533 10.6151
R1396 B.n535 B.n534 10.6151
R1397 B.n535 B.n170 10.6151
R1398 B.n539 B.n170 10.6151
R1399 B.n540 B.n539 10.6151
R1400 B.n541 B.n540 10.6151
R1401 B.n541 B.n168 10.6151
R1402 B.n545 B.n168 10.6151
R1403 B.n546 B.n545 10.6151
R1404 B.n547 B.n546 10.6151
R1405 B.n547 B.n166 10.6151
R1406 B.n551 B.n166 10.6151
R1407 B.n552 B.n551 10.6151
R1408 B.n553 B.n552 10.6151
R1409 B.n553 B.n164 10.6151
R1410 B.n557 B.n164 10.6151
R1411 B.n558 B.n557 10.6151
R1412 B.n559 B.n558 10.6151
R1413 B.n559 B.n162 10.6151
R1414 B.n563 B.n162 10.6151
R1415 B.n564 B.n563 10.6151
R1416 B.n565 B.n564 10.6151
R1417 B.n565 B.n160 10.6151
R1418 B.n569 B.n160 10.6151
R1419 B.n570 B.n569 10.6151
R1420 B.n571 B.n570 10.6151
R1421 B.n571 B.n158 10.6151
R1422 B.n575 B.n158 10.6151
R1423 B.n576 B.n575 10.6151
R1424 B.n577 B.n576 10.6151
R1425 B.n577 B.n156 10.6151
R1426 B.n581 B.n156 10.6151
R1427 B.n582 B.n581 10.6151
R1428 B.n583 B.n582 10.6151
R1429 B.n583 B.n154 10.6151
R1430 B.n587 B.n154 10.6151
R1431 B.n588 B.n587 10.6151
R1432 B.n589 B.n588 10.6151
R1433 B.n589 B.n152 10.6151
R1434 B.n593 B.n152 10.6151
R1435 B.n594 B.n593 10.6151
R1436 B.n595 B.n594 10.6151
R1437 B.n595 B.n150 10.6151
R1438 B.n599 B.n150 10.6151
R1439 B.n600 B.n599 10.6151
R1440 B.n601 B.n600 10.6151
R1441 B.n601 B.n148 10.6151
R1442 B.n605 B.n148 10.6151
R1443 B.n606 B.n605 10.6151
R1444 B.n607 B.n606 10.6151
R1445 B.n607 B.n146 10.6151
R1446 B.n611 B.n146 10.6151
R1447 B.n612 B.n611 10.6151
R1448 B.n613 B.n612 10.6151
R1449 B.n613 B.n144 10.6151
R1450 B.n617 B.n144 10.6151
R1451 B.n618 B.n617 10.6151
R1452 B.n619 B.n618 10.6151
R1453 B.n619 B.n142 10.6151
R1454 B.n623 B.n142 10.6151
R1455 B.n624 B.n623 10.6151
R1456 B.n625 B.n624 10.6151
R1457 B.n625 B.n140 10.6151
R1458 B.n629 B.n140 10.6151
R1459 B.n630 B.n629 10.6151
R1460 B.n631 B.n630 10.6151
R1461 B.n631 B.n138 10.6151
R1462 B.n635 B.n138 10.6151
R1463 B.n636 B.n635 10.6151
R1464 B.n637 B.n636 10.6151
R1465 B.n637 B.n136 10.6151
R1466 B.n641 B.n136 10.6151
R1467 B.n642 B.n641 10.6151
R1468 B.n643 B.n642 10.6151
R1469 B.n643 B.n134 10.6151
R1470 B.n647 B.n134 10.6151
R1471 B.n648 B.n647 10.6151
R1472 B.n649 B.n648 10.6151
R1473 B.n649 B.n132 10.6151
R1474 B.n653 B.n132 10.6151
R1475 B.n654 B.n653 10.6151
R1476 B.n655 B.n654 10.6151
R1477 B.n655 B.n130 10.6151
R1478 B.n659 B.n130 10.6151
R1479 B.n660 B.n659 10.6151
R1480 B.n661 B.n660 10.6151
R1481 B.n661 B.n128 10.6151
R1482 B.n665 B.n128 10.6151
R1483 B.n666 B.n665 10.6151
R1484 B.n667 B.n666 10.6151
R1485 B.n667 B.n126 10.6151
R1486 B.n671 B.n126 10.6151
R1487 B.n672 B.n671 10.6151
R1488 B.n673 B.n672 10.6151
R1489 B.n673 B.n124 10.6151
R1490 B.n677 B.n124 10.6151
R1491 B.n678 B.n677 10.6151
R1492 B.n679 B.n678 10.6151
R1493 B.n679 B.n122 10.6151
R1494 B.n683 B.n122 10.6151
R1495 B.n684 B.n683 10.6151
R1496 B.n685 B.n684 10.6151
R1497 B.n685 B.n120 10.6151
R1498 B.n689 B.n120 10.6151
R1499 B.n690 B.n689 10.6151
R1500 B.n691 B.n690 10.6151
R1501 B.n691 B.n118 10.6151
R1502 B.n695 B.n118 10.6151
R1503 B.n696 B.n695 10.6151
R1504 B.n697 B.n696 10.6151
R1505 B.n697 B.n116 10.6151
R1506 B.n701 B.n116 10.6151
R1507 B.n702 B.n701 10.6151
R1508 B.n703 B.n702 10.6151
R1509 B.n703 B.n114 10.6151
R1510 B.n707 B.n114 10.6151
R1511 B.n708 B.n707 10.6151
R1512 B.n709 B.n708 10.6151
R1513 B.n709 B.n112 10.6151
R1514 B.n713 B.n112 10.6151
R1515 B.n714 B.n713 10.6151
R1516 B.n715 B.n714 10.6151
R1517 B.n715 B.n110 10.6151
R1518 B.n719 B.n110 10.6151
R1519 B.n720 B.n719 10.6151
R1520 B.n721 B.n720 10.6151
R1521 B.n721 B.n108 10.6151
R1522 B.n725 B.n108 10.6151
R1523 B.n726 B.n725 10.6151
R1524 B.n727 B.n726 10.6151
R1525 B.n727 B.n106 10.6151
R1526 B.n731 B.n106 10.6151
R1527 B.n732 B.n731 10.6151
R1528 B.n733 B.n732 10.6151
R1529 B.n733 B.n104 10.6151
R1530 B.n737 B.n104 10.6151
R1531 B.n738 B.n737 10.6151
R1532 B.n739 B.n738 10.6151
R1533 B.n739 B.n102 10.6151
R1534 B.n743 B.n102 10.6151
R1535 B.n744 B.n743 10.6151
R1536 B.n745 B.n744 10.6151
R1537 B.n745 B.n100 10.6151
R1538 B.n749 B.n100 10.6151
R1539 B.n750 B.n749 10.6151
R1540 B.n751 B.n750 10.6151
R1541 B.n751 B.n98 10.6151
R1542 B.n755 B.n98 10.6151
R1543 B.n756 B.n755 10.6151
R1544 B.n757 B.n756 10.6151
R1545 B.n757 B.n96 10.6151
R1546 B.n761 B.n96 10.6151
R1547 B.n762 B.n761 10.6151
R1548 B.n379 B.n226 10.6151
R1549 B.n383 B.n226 10.6151
R1550 B.n384 B.n383 10.6151
R1551 B.n385 B.n384 10.6151
R1552 B.n385 B.n224 10.6151
R1553 B.n389 B.n224 10.6151
R1554 B.n390 B.n389 10.6151
R1555 B.n391 B.n390 10.6151
R1556 B.n391 B.n222 10.6151
R1557 B.n395 B.n222 10.6151
R1558 B.n396 B.n395 10.6151
R1559 B.n397 B.n396 10.6151
R1560 B.n397 B.n220 10.6151
R1561 B.n401 B.n220 10.6151
R1562 B.n402 B.n401 10.6151
R1563 B.n403 B.n402 10.6151
R1564 B.n403 B.n218 10.6151
R1565 B.n407 B.n218 10.6151
R1566 B.n408 B.n407 10.6151
R1567 B.n409 B.n408 10.6151
R1568 B.n409 B.n216 10.6151
R1569 B.n413 B.n216 10.6151
R1570 B.n414 B.n413 10.6151
R1571 B.n415 B.n414 10.6151
R1572 B.n415 B.n214 10.6151
R1573 B.n419 B.n214 10.6151
R1574 B.n420 B.n419 10.6151
R1575 B.n421 B.n420 10.6151
R1576 B.n421 B.n212 10.6151
R1577 B.n425 B.n212 10.6151
R1578 B.n426 B.n425 10.6151
R1579 B.n427 B.n426 10.6151
R1580 B.n427 B.n210 10.6151
R1581 B.n431 B.n210 10.6151
R1582 B.n432 B.n431 10.6151
R1583 B.n433 B.n432 10.6151
R1584 B.n433 B.n208 10.6151
R1585 B.n437 B.n208 10.6151
R1586 B.n438 B.n437 10.6151
R1587 B.n439 B.n438 10.6151
R1588 B.n439 B.n206 10.6151
R1589 B.n443 B.n206 10.6151
R1590 B.n444 B.n443 10.6151
R1591 B.n445 B.n444 10.6151
R1592 B.n449 B.n448 10.6151
R1593 B.n450 B.n449 10.6151
R1594 B.n450 B.n200 10.6151
R1595 B.n454 B.n200 10.6151
R1596 B.n455 B.n454 10.6151
R1597 B.n456 B.n455 10.6151
R1598 B.n456 B.n198 10.6151
R1599 B.n460 B.n198 10.6151
R1600 B.n461 B.n460 10.6151
R1601 B.n463 B.n194 10.6151
R1602 B.n467 B.n194 10.6151
R1603 B.n468 B.n467 10.6151
R1604 B.n469 B.n468 10.6151
R1605 B.n469 B.n192 10.6151
R1606 B.n473 B.n192 10.6151
R1607 B.n474 B.n473 10.6151
R1608 B.n475 B.n474 10.6151
R1609 B.n475 B.n190 10.6151
R1610 B.n479 B.n190 10.6151
R1611 B.n480 B.n479 10.6151
R1612 B.n481 B.n480 10.6151
R1613 B.n481 B.n188 10.6151
R1614 B.n485 B.n188 10.6151
R1615 B.n486 B.n485 10.6151
R1616 B.n487 B.n486 10.6151
R1617 B.n487 B.n186 10.6151
R1618 B.n491 B.n186 10.6151
R1619 B.n492 B.n491 10.6151
R1620 B.n493 B.n492 10.6151
R1621 B.n493 B.n184 10.6151
R1622 B.n497 B.n184 10.6151
R1623 B.n498 B.n497 10.6151
R1624 B.n499 B.n498 10.6151
R1625 B.n499 B.n182 10.6151
R1626 B.n503 B.n182 10.6151
R1627 B.n504 B.n503 10.6151
R1628 B.n505 B.n504 10.6151
R1629 B.n505 B.n180 10.6151
R1630 B.n509 B.n180 10.6151
R1631 B.n510 B.n509 10.6151
R1632 B.n511 B.n510 10.6151
R1633 B.n511 B.n178 10.6151
R1634 B.n515 B.n178 10.6151
R1635 B.n516 B.n515 10.6151
R1636 B.n517 B.n516 10.6151
R1637 B.n517 B.n176 10.6151
R1638 B.n521 B.n176 10.6151
R1639 B.n522 B.n521 10.6151
R1640 B.n523 B.n522 10.6151
R1641 B.n523 B.n174 10.6151
R1642 B.n527 B.n174 10.6151
R1643 B.n528 B.n527 10.6151
R1644 B.n529 B.n528 10.6151
R1645 B.n378 B.n377 10.6151
R1646 B.n377 B.n228 10.6151
R1647 B.n373 B.n228 10.6151
R1648 B.n373 B.n372 10.6151
R1649 B.n372 B.n371 10.6151
R1650 B.n371 B.n230 10.6151
R1651 B.n367 B.n230 10.6151
R1652 B.n367 B.n366 10.6151
R1653 B.n366 B.n365 10.6151
R1654 B.n365 B.n232 10.6151
R1655 B.n361 B.n232 10.6151
R1656 B.n361 B.n360 10.6151
R1657 B.n360 B.n359 10.6151
R1658 B.n359 B.n234 10.6151
R1659 B.n355 B.n234 10.6151
R1660 B.n355 B.n354 10.6151
R1661 B.n354 B.n353 10.6151
R1662 B.n353 B.n236 10.6151
R1663 B.n349 B.n236 10.6151
R1664 B.n349 B.n348 10.6151
R1665 B.n348 B.n347 10.6151
R1666 B.n347 B.n238 10.6151
R1667 B.n343 B.n238 10.6151
R1668 B.n343 B.n342 10.6151
R1669 B.n342 B.n341 10.6151
R1670 B.n341 B.n240 10.6151
R1671 B.n337 B.n240 10.6151
R1672 B.n337 B.n336 10.6151
R1673 B.n336 B.n335 10.6151
R1674 B.n335 B.n242 10.6151
R1675 B.n331 B.n242 10.6151
R1676 B.n331 B.n330 10.6151
R1677 B.n330 B.n329 10.6151
R1678 B.n329 B.n244 10.6151
R1679 B.n325 B.n244 10.6151
R1680 B.n325 B.n324 10.6151
R1681 B.n324 B.n323 10.6151
R1682 B.n323 B.n246 10.6151
R1683 B.n319 B.n246 10.6151
R1684 B.n319 B.n318 10.6151
R1685 B.n318 B.n317 10.6151
R1686 B.n317 B.n248 10.6151
R1687 B.n313 B.n248 10.6151
R1688 B.n313 B.n312 10.6151
R1689 B.n312 B.n311 10.6151
R1690 B.n311 B.n250 10.6151
R1691 B.n307 B.n250 10.6151
R1692 B.n307 B.n306 10.6151
R1693 B.n306 B.n305 10.6151
R1694 B.n305 B.n252 10.6151
R1695 B.n301 B.n252 10.6151
R1696 B.n301 B.n300 10.6151
R1697 B.n300 B.n299 10.6151
R1698 B.n299 B.n254 10.6151
R1699 B.n295 B.n254 10.6151
R1700 B.n295 B.n294 10.6151
R1701 B.n294 B.n293 10.6151
R1702 B.n293 B.n256 10.6151
R1703 B.n289 B.n256 10.6151
R1704 B.n289 B.n288 10.6151
R1705 B.n288 B.n287 10.6151
R1706 B.n287 B.n258 10.6151
R1707 B.n283 B.n258 10.6151
R1708 B.n283 B.n282 10.6151
R1709 B.n282 B.n281 10.6151
R1710 B.n281 B.n260 10.6151
R1711 B.n277 B.n260 10.6151
R1712 B.n277 B.n276 10.6151
R1713 B.n276 B.n275 10.6151
R1714 B.n275 B.n262 10.6151
R1715 B.n271 B.n262 10.6151
R1716 B.n271 B.n270 10.6151
R1717 B.n270 B.n269 10.6151
R1718 B.n269 B.n264 10.6151
R1719 B.n265 B.n264 10.6151
R1720 B.n265 B.n0 10.6151
R1721 B.n1027 B.n1 10.6151
R1722 B.n1027 B.n1026 10.6151
R1723 B.n1026 B.n1025 10.6151
R1724 B.n1025 B.n4 10.6151
R1725 B.n1021 B.n4 10.6151
R1726 B.n1021 B.n1020 10.6151
R1727 B.n1020 B.n1019 10.6151
R1728 B.n1019 B.n6 10.6151
R1729 B.n1015 B.n6 10.6151
R1730 B.n1015 B.n1014 10.6151
R1731 B.n1014 B.n1013 10.6151
R1732 B.n1013 B.n8 10.6151
R1733 B.n1009 B.n8 10.6151
R1734 B.n1009 B.n1008 10.6151
R1735 B.n1008 B.n1007 10.6151
R1736 B.n1007 B.n10 10.6151
R1737 B.n1003 B.n10 10.6151
R1738 B.n1003 B.n1002 10.6151
R1739 B.n1002 B.n1001 10.6151
R1740 B.n1001 B.n12 10.6151
R1741 B.n997 B.n12 10.6151
R1742 B.n997 B.n996 10.6151
R1743 B.n996 B.n995 10.6151
R1744 B.n995 B.n14 10.6151
R1745 B.n991 B.n14 10.6151
R1746 B.n991 B.n990 10.6151
R1747 B.n990 B.n989 10.6151
R1748 B.n989 B.n16 10.6151
R1749 B.n985 B.n16 10.6151
R1750 B.n985 B.n984 10.6151
R1751 B.n984 B.n983 10.6151
R1752 B.n983 B.n18 10.6151
R1753 B.n979 B.n18 10.6151
R1754 B.n979 B.n978 10.6151
R1755 B.n978 B.n977 10.6151
R1756 B.n977 B.n20 10.6151
R1757 B.n973 B.n20 10.6151
R1758 B.n973 B.n972 10.6151
R1759 B.n972 B.n971 10.6151
R1760 B.n971 B.n22 10.6151
R1761 B.n967 B.n22 10.6151
R1762 B.n967 B.n966 10.6151
R1763 B.n966 B.n965 10.6151
R1764 B.n965 B.n24 10.6151
R1765 B.n961 B.n24 10.6151
R1766 B.n961 B.n960 10.6151
R1767 B.n960 B.n959 10.6151
R1768 B.n959 B.n26 10.6151
R1769 B.n955 B.n26 10.6151
R1770 B.n955 B.n954 10.6151
R1771 B.n954 B.n953 10.6151
R1772 B.n953 B.n28 10.6151
R1773 B.n949 B.n28 10.6151
R1774 B.n949 B.n948 10.6151
R1775 B.n948 B.n947 10.6151
R1776 B.n947 B.n30 10.6151
R1777 B.n943 B.n30 10.6151
R1778 B.n943 B.n942 10.6151
R1779 B.n942 B.n941 10.6151
R1780 B.n941 B.n32 10.6151
R1781 B.n937 B.n32 10.6151
R1782 B.n937 B.n936 10.6151
R1783 B.n936 B.n935 10.6151
R1784 B.n935 B.n34 10.6151
R1785 B.n931 B.n34 10.6151
R1786 B.n931 B.n930 10.6151
R1787 B.n930 B.n929 10.6151
R1788 B.n929 B.n36 10.6151
R1789 B.n925 B.n36 10.6151
R1790 B.n925 B.n924 10.6151
R1791 B.n924 B.n923 10.6151
R1792 B.n923 B.n38 10.6151
R1793 B.n919 B.n38 10.6151
R1794 B.n919 B.n918 10.6151
R1795 B.n918 B.n917 10.6151
R1796 B.n917 B.n40 10.6151
R1797 B.n847 B.n846 9.36635
R1798 B.n829 B.n72 9.36635
R1799 B.n445 B.n204 9.36635
R1800 B.n463 B.n462 9.36635
R1801 B.n1031 B.n0 2.81026
R1802 B.n1031 B.n1 2.81026
R1803 B.n846 B.n845 1.24928
R1804 B.n832 B.n72 1.24928
R1805 B.n448 B.n204 1.24928
R1806 B.n462 B.n461 1.24928
R1807 VN.n106 VN.n105 161.3
R1808 VN.n104 VN.n55 161.3
R1809 VN.n103 VN.n102 161.3
R1810 VN.n101 VN.n56 161.3
R1811 VN.n100 VN.n99 161.3
R1812 VN.n98 VN.n57 161.3
R1813 VN.n97 VN.n96 161.3
R1814 VN.n95 VN.n58 161.3
R1815 VN.n94 VN.n93 161.3
R1816 VN.n92 VN.n59 161.3
R1817 VN.n91 VN.n90 161.3
R1818 VN.n89 VN.n61 161.3
R1819 VN.n88 VN.n87 161.3
R1820 VN.n86 VN.n62 161.3
R1821 VN.n85 VN.n84 161.3
R1822 VN.n83 VN.n63 161.3
R1823 VN.n82 VN.n81 161.3
R1824 VN.n80 VN.n64 161.3
R1825 VN.n79 VN.n78 161.3
R1826 VN.n77 VN.n66 161.3
R1827 VN.n76 VN.n75 161.3
R1828 VN.n74 VN.n67 161.3
R1829 VN.n73 VN.n72 161.3
R1830 VN.n71 VN.n68 161.3
R1831 VN.n52 VN.n51 161.3
R1832 VN.n50 VN.n1 161.3
R1833 VN.n49 VN.n48 161.3
R1834 VN.n47 VN.n2 161.3
R1835 VN.n46 VN.n45 161.3
R1836 VN.n44 VN.n3 161.3
R1837 VN.n43 VN.n42 161.3
R1838 VN.n41 VN.n4 161.3
R1839 VN.n40 VN.n39 161.3
R1840 VN.n37 VN.n5 161.3
R1841 VN.n36 VN.n35 161.3
R1842 VN.n34 VN.n6 161.3
R1843 VN.n33 VN.n32 161.3
R1844 VN.n31 VN.n7 161.3
R1845 VN.n30 VN.n29 161.3
R1846 VN.n28 VN.n8 161.3
R1847 VN.n27 VN.n26 161.3
R1848 VN.n24 VN.n9 161.3
R1849 VN.n23 VN.n22 161.3
R1850 VN.n21 VN.n10 161.3
R1851 VN.n20 VN.n19 161.3
R1852 VN.n18 VN.n11 161.3
R1853 VN.n17 VN.n16 161.3
R1854 VN.n15 VN.n12 161.3
R1855 VN.n70 VN.t5 120.981
R1856 VN.n14 VN.t3 120.981
R1857 VN.n13 VN.t4 88.8608
R1858 VN.n25 VN.t1 88.8608
R1859 VN.n38 VN.t2 88.8608
R1860 VN.n0 VN.t0 88.8608
R1861 VN.n69 VN.t9 88.8608
R1862 VN.n65 VN.t7 88.8608
R1863 VN.n60 VN.t6 88.8608
R1864 VN.n54 VN.t8 88.8608
R1865 VN.n53 VN.n0 86.8027
R1866 VN.n107 VN.n54 86.8027
R1867 VN.n14 VN.n13 67.0059
R1868 VN.n70 VN.n69 67.0059
R1869 VN VN.n107 59.5246
R1870 VN.n19 VN.n10 56.5617
R1871 VN.n32 VN.n6 56.5617
R1872 VN.n75 VN.n66 56.5617
R1873 VN.n87 VN.n61 56.5617
R1874 VN.n45 VN.n2 51.7179
R1875 VN.n99 VN.n56 51.7179
R1876 VN.n45 VN.n44 29.4362
R1877 VN.n99 VN.n98 29.4362
R1878 VN.n17 VN.n12 24.5923
R1879 VN.n18 VN.n17 24.5923
R1880 VN.n19 VN.n18 24.5923
R1881 VN.n23 VN.n10 24.5923
R1882 VN.n24 VN.n23 24.5923
R1883 VN.n26 VN.n24 24.5923
R1884 VN.n30 VN.n8 24.5923
R1885 VN.n31 VN.n30 24.5923
R1886 VN.n32 VN.n31 24.5923
R1887 VN.n36 VN.n6 24.5923
R1888 VN.n37 VN.n36 24.5923
R1889 VN.n39 VN.n37 24.5923
R1890 VN.n43 VN.n4 24.5923
R1891 VN.n44 VN.n43 24.5923
R1892 VN.n49 VN.n2 24.5923
R1893 VN.n50 VN.n49 24.5923
R1894 VN.n51 VN.n50 24.5923
R1895 VN.n75 VN.n74 24.5923
R1896 VN.n74 VN.n73 24.5923
R1897 VN.n73 VN.n68 24.5923
R1898 VN.n87 VN.n86 24.5923
R1899 VN.n86 VN.n85 24.5923
R1900 VN.n85 VN.n63 24.5923
R1901 VN.n81 VN.n80 24.5923
R1902 VN.n80 VN.n79 24.5923
R1903 VN.n79 VN.n66 24.5923
R1904 VN.n98 VN.n97 24.5923
R1905 VN.n97 VN.n58 24.5923
R1906 VN.n93 VN.n92 24.5923
R1907 VN.n92 VN.n91 24.5923
R1908 VN.n91 VN.n61 24.5923
R1909 VN.n105 VN.n104 24.5923
R1910 VN.n104 VN.n103 24.5923
R1911 VN.n103 VN.n56 24.5923
R1912 VN.n38 VN.n4 16.7229
R1913 VN.n60 VN.n58 16.7229
R1914 VN.n26 VN.n25 12.2964
R1915 VN.n25 VN.n8 12.2964
R1916 VN.n65 VN.n63 12.2964
R1917 VN.n81 VN.n65 12.2964
R1918 VN.n13 VN.n12 7.86989
R1919 VN.n39 VN.n38 7.86989
R1920 VN.n69 VN.n68 7.86989
R1921 VN.n93 VN.n60 7.86989
R1922 VN.n51 VN.n0 3.44336
R1923 VN.n105 VN.n54 3.44336
R1924 VN.n71 VN.n70 3.35172
R1925 VN.n15 VN.n14 3.35172
R1926 VN.n107 VN.n106 0.354861
R1927 VN.n53 VN.n52 0.354861
R1928 VN VN.n53 0.267071
R1929 VN.n106 VN.n55 0.189894
R1930 VN.n102 VN.n55 0.189894
R1931 VN.n102 VN.n101 0.189894
R1932 VN.n101 VN.n100 0.189894
R1933 VN.n100 VN.n57 0.189894
R1934 VN.n96 VN.n57 0.189894
R1935 VN.n96 VN.n95 0.189894
R1936 VN.n95 VN.n94 0.189894
R1937 VN.n94 VN.n59 0.189894
R1938 VN.n90 VN.n59 0.189894
R1939 VN.n90 VN.n89 0.189894
R1940 VN.n89 VN.n88 0.189894
R1941 VN.n88 VN.n62 0.189894
R1942 VN.n84 VN.n62 0.189894
R1943 VN.n84 VN.n83 0.189894
R1944 VN.n83 VN.n82 0.189894
R1945 VN.n82 VN.n64 0.189894
R1946 VN.n78 VN.n64 0.189894
R1947 VN.n78 VN.n77 0.189894
R1948 VN.n77 VN.n76 0.189894
R1949 VN.n76 VN.n67 0.189894
R1950 VN.n72 VN.n67 0.189894
R1951 VN.n72 VN.n71 0.189894
R1952 VN.n16 VN.n15 0.189894
R1953 VN.n16 VN.n11 0.189894
R1954 VN.n20 VN.n11 0.189894
R1955 VN.n21 VN.n20 0.189894
R1956 VN.n22 VN.n21 0.189894
R1957 VN.n22 VN.n9 0.189894
R1958 VN.n27 VN.n9 0.189894
R1959 VN.n28 VN.n27 0.189894
R1960 VN.n29 VN.n28 0.189894
R1961 VN.n29 VN.n7 0.189894
R1962 VN.n33 VN.n7 0.189894
R1963 VN.n34 VN.n33 0.189894
R1964 VN.n35 VN.n34 0.189894
R1965 VN.n35 VN.n5 0.189894
R1966 VN.n40 VN.n5 0.189894
R1967 VN.n41 VN.n40 0.189894
R1968 VN.n42 VN.n41 0.189894
R1969 VN.n42 VN.n3 0.189894
R1970 VN.n46 VN.n3 0.189894
R1971 VN.n47 VN.n46 0.189894
R1972 VN.n48 VN.n47 0.189894
R1973 VN.n48 VN.n1 0.189894
R1974 VN.n52 VN.n1 0.189894
R1975 VDD2.n1 VDD2.t6 78.4676
R1976 VDD2.n3 VDD2.n2 75.1073
R1977 VDD2 VDD2.n7 75.1043
R1978 VDD2.n4 VDD2.t1 75.0972
R1979 VDD2.n6 VDD2.n5 72.6347
R1980 VDD2.n1 VDD2.n0 72.6346
R1981 VDD2.n4 VDD2.n3 51.1054
R1982 VDD2.n6 VDD2.n4 3.37119
R1983 VDD2.n7 VDD2.t0 2.463
R1984 VDD2.n7 VDD2.t4 2.463
R1985 VDD2.n5 VDD2.t3 2.463
R1986 VDD2.n5 VDD2.t2 2.463
R1987 VDD2.n2 VDD2.t7 2.463
R1988 VDD2.n2 VDD2.t9 2.463
R1989 VDD2.n0 VDD2.t5 2.463
R1990 VDD2.n0 VDD2.t8 2.463
R1991 VDD2 VDD2.n6 0.901362
R1992 VDD2.n3 VDD2.n1 0.787826
C0 VN VP 10.061f
C1 VDD2 VDD1 2.81349f
C2 VTAIL VDD2 11.3905f
C3 VDD2 w_n5662_n3608# 3.43794f
C4 VTAIL VDD1 11.3324f
C5 w_n5662_n3608# VDD1 3.24345f
C6 VTAIL w_n5662_n3608# 3.51716f
C7 VDD2 VP 0.709064f
C8 VN B 1.55136f
C9 VP VDD1 12.895599f
C10 VTAIL VP 13.3665f
C11 w_n5662_n3608# VP 13.161201f
C12 B VDD2 3.11407f
C13 B VDD1 2.95799f
C14 VTAIL B 4.38911f
C15 B w_n5662_n3608# 12.5308f
C16 B VP 2.80143f
C17 VN VDD2 12.3466f
C18 VN VDD1 0.156012f
C19 VTAIL VN 13.352201f
C20 VN w_n5662_n3608# 12.421f
C21 VDD2 VSUBS 2.55197f
C22 VDD1 VSUBS 2.393872f
C23 VTAIL VSUBS 1.575726f
C24 VN VSUBS 9.35511f
C25 VP VSUBS 5.528338f
C26 B VSUBS 6.682472f
C27 w_n5662_n3608# VSUBS 0.251053p
C28 VDD2.t6 VSUBS 3.32245f
C29 VDD2.t5 VSUBS 0.317218f
C30 VDD2.t8 VSUBS 0.317218f
C31 VDD2.n0 VSUBS 2.51368f
C32 VDD2.n1 VSUBS 1.97143f
C33 VDD2.t7 VSUBS 0.317218f
C34 VDD2.t9 VSUBS 0.317218f
C35 VDD2.n2 VSUBS 2.5521f
C36 VDD2.n3 VSUBS 4.57074f
C37 VDD2.t1 VSUBS 3.27843f
C38 VDD2.n4 VSUBS 4.72847f
C39 VDD2.t3 VSUBS 0.317218f
C40 VDD2.t2 VSUBS 0.317218f
C41 VDD2.n5 VSUBS 2.51368f
C42 VDD2.n6 VSUBS 1.00066f
C43 VDD2.t0 VSUBS 0.317218f
C44 VDD2.t4 VSUBS 0.317218f
C45 VDD2.n7 VSUBS 2.55203f
C46 VN.t0 VSUBS 2.98756f
C47 VN.n0 VSUBS 1.125f
C48 VN.n1 VSUBS 0.023143f
C49 VN.n2 VSUBS 0.041584f
C50 VN.n3 VSUBS 0.023143f
C51 VN.n4 VSUBS 0.036137f
C52 VN.n5 VSUBS 0.023143f
C53 VN.n6 VSUBS 0.036524f
C54 VN.n7 VSUBS 0.023143f
C55 VN.n8 VSUBS 0.032324f
C56 VN.n9 VSUBS 0.023143f
C57 VN.n10 VSUBS 0.030761f
C58 VN.n11 VSUBS 0.023143f
C59 VN.n12 VSUBS 0.02851f
C60 VN.t4 VSUBS 2.98756f
C61 VN.n13 VSUBS 1.11913f
C62 VN.t3 VSUBS 3.31011f
C63 VN.n14 VSUBS 1.06967f
C64 VN.n15 VSUBS 0.290104f
C65 VN.n16 VSUBS 0.023143f
C66 VN.n17 VSUBS 0.042917f
C67 VN.n18 VSUBS 0.042917f
C68 VN.n19 VSUBS 0.036524f
C69 VN.n20 VSUBS 0.023143f
C70 VN.n21 VSUBS 0.023143f
C71 VN.n22 VSUBS 0.023143f
C72 VN.n23 VSUBS 0.042917f
C73 VN.n24 VSUBS 0.042917f
C74 VN.t1 VSUBS 2.98756f
C75 VN.n25 VSUBS 1.04284f
C76 VN.n26 VSUBS 0.032324f
C77 VN.n27 VSUBS 0.023143f
C78 VN.n28 VSUBS 0.023143f
C79 VN.n29 VSUBS 0.023143f
C80 VN.n30 VSUBS 0.042917f
C81 VN.n31 VSUBS 0.042917f
C82 VN.n32 VSUBS 0.030761f
C83 VN.n33 VSUBS 0.023143f
C84 VN.n34 VSUBS 0.023143f
C85 VN.n35 VSUBS 0.023143f
C86 VN.n36 VSUBS 0.042917f
C87 VN.n37 VSUBS 0.042917f
C88 VN.t2 VSUBS 2.98756f
C89 VN.n38 VSUBS 1.04284f
C90 VN.n39 VSUBS 0.02851f
C91 VN.n40 VSUBS 0.023143f
C92 VN.n41 VSUBS 0.023143f
C93 VN.n42 VSUBS 0.023143f
C94 VN.n43 VSUBS 0.042917f
C95 VN.n44 VSUBS 0.045706f
C96 VN.n45 VSUBS 0.022912f
C97 VN.n46 VSUBS 0.023143f
C98 VN.n47 VSUBS 0.023143f
C99 VN.n48 VSUBS 0.023143f
C100 VN.n49 VSUBS 0.042917f
C101 VN.n50 VSUBS 0.042917f
C102 VN.n51 VSUBS 0.024696f
C103 VN.n52 VSUBS 0.037347f
C104 VN.n53 VSUBS 0.067824f
C105 VN.t8 VSUBS 2.98756f
C106 VN.n54 VSUBS 1.125f
C107 VN.n55 VSUBS 0.023143f
C108 VN.n56 VSUBS 0.041584f
C109 VN.n57 VSUBS 0.023143f
C110 VN.n58 VSUBS 0.036137f
C111 VN.n59 VSUBS 0.023143f
C112 VN.t6 VSUBS 2.98756f
C113 VN.n60 VSUBS 1.04284f
C114 VN.n61 VSUBS 0.036524f
C115 VN.n62 VSUBS 0.023143f
C116 VN.n63 VSUBS 0.032324f
C117 VN.n64 VSUBS 0.023143f
C118 VN.t7 VSUBS 2.98756f
C119 VN.n65 VSUBS 1.04284f
C120 VN.n66 VSUBS 0.030761f
C121 VN.n67 VSUBS 0.023143f
C122 VN.n68 VSUBS 0.02851f
C123 VN.t5 VSUBS 3.31011f
C124 VN.t9 VSUBS 2.98756f
C125 VN.n69 VSUBS 1.11913f
C126 VN.n70 VSUBS 1.06967f
C127 VN.n71 VSUBS 0.290104f
C128 VN.n72 VSUBS 0.023143f
C129 VN.n73 VSUBS 0.042917f
C130 VN.n74 VSUBS 0.042917f
C131 VN.n75 VSUBS 0.036524f
C132 VN.n76 VSUBS 0.023143f
C133 VN.n77 VSUBS 0.023143f
C134 VN.n78 VSUBS 0.023143f
C135 VN.n79 VSUBS 0.042917f
C136 VN.n80 VSUBS 0.042917f
C137 VN.n81 VSUBS 0.032324f
C138 VN.n82 VSUBS 0.023143f
C139 VN.n83 VSUBS 0.023143f
C140 VN.n84 VSUBS 0.023143f
C141 VN.n85 VSUBS 0.042917f
C142 VN.n86 VSUBS 0.042917f
C143 VN.n87 VSUBS 0.030761f
C144 VN.n88 VSUBS 0.023143f
C145 VN.n89 VSUBS 0.023143f
C146 VN.n90 VSUBS 0.023143f
C147 VN.n91 VSUBS 0.042917f
C148 VN.n92 VSUBS 0.042917f
C149 VN.n93 VSUBS 0.02851f
C150 VN.n94 VSUBS 0.023143f
C151 VN.n95 VSUBS 0.023143f
C152 VN.n96 VSUBS 0.023143f
C153 VN.n97 VSUBS 0.042917f
C154 VN.n98 VSUBS 0.045706f
C155 VN.n99 VSUBS 0.022912f
C156 VN.n100 VSUBS 0.023143f
C157 VN.n101 VSUBS 0.023143f
C158 VN.n102 VSUBS 0.023143f
C159 VN.n103 VSUBS 0.042917f
C160 VN.n104 VSUBS 0.042917f
C161 VN.n105 VSUBS 0.024696f
C162 VN.n106 VSUBS 0.037347f
C163 VN.n107 VSUBS 1.68985f
C164 B.n0 VSUBS 0.005428f
C165 B.n1 VSUBS 0.005428f
C166 B.n2 VSUBS 0.008583f
C167 B.n3 VSUBS 0.008583f
C168 B.n4 VSUBS 0.008583f
C169 B.n5 VSUBS 0.008583f
C170 B.n6 VSUBS 0.008583f
C171 B.n7 VSUBS 0.008583f
C172 B.n8 VSUBS 0.008583f
C173 B.n9 VSUBS 0.008583f
C174 B.n10 VSUBS 0.008583f
C175 B.n11 VSUBS 0.008583f
C176 B.n12 VSUBS 0.008583f
C177 B.n13 VSUBS 0.008583f
C178 B.n14 VSUBS 0.008583f
C179 B.n15 VSUBS 0.008583f
C180 B.n16 VSUBS 0.008583f
C181 B.n17 VSUBS 0.008583f
C182 B.n18 VSUBS 0.008583f
C183 B.n19 VSUBS 0.008583f
C184 B.n20 VSUBS 0.008583f
C185 B.n21 VSUBS 0.008583f
C186 B.n22 VSUBS 0.008583f
C187 B.n23 VSUBS 0.008583f
C188 B.n24 VSUBS 0.008583f
C189 B.n25 VSUBS 0.008583f
C190 B.n26 VSUBS 0.008583f
C191 B.n27 VSUBS 0.008583f
C192 B.n28 VSUBS 0.008583f
C193 B.n29 VSUBS 0.008583f
C194 B.n30 VSUBS 0.008583f
C195 B.n31 VSUBS 0.008583f
C196 B.n32 VSUBS 0.008583f
C197 B.n33 VSUBS 0.008583f
C198 B.n34 VSUBS 0.008583f
C199 B.n35 VSUBS 0.008583f
C200 B.n36 VSUBS 0.008583f
C201 B.n37 VSUBS 0.008583f
C202 B.n38 VSUBS 0.008583f
C203 B.n39 VSUBS 0.008583f
C204 B.n40 VSUBS 0.019571f
C205 B.n41 VSUBS 0.008583f
C206 B.n42 VSUBS 0.008583f
C207 B.n43 VSUBS 0.008583f
C208 B.n44 VSUBS 0.008583f
C209 B.n45 VSUBS 0.008583f
C210 B.n46 VSUBS 0.008583f
C211 B.n47 VSUBS 0.008583f
C212 B.n48 VSUBS 0.008583f
C213 B.n49 VSUBS 0.008583f
C214 B.n50 VSUBS 0.008583f
C215 B.n51 VSUBS 0.008583f
C216 B.n52 VSUBS 0.008583f
C217 B.n53 VSUBS 0.008583f
C218 B.n54 VSUBS 0.008583f
C219 B.n55 VSUBS 0.008583f
C220 B.n56 VSUBS 0.008583f
C221 B.n57 VSUBS 0.008583f
C222 B.n58 VSUBS 0.008583f
C223 B.n59 VSUBS 0.008583f
C224 B.n60 VSUBS 0.008583f
C225 B.n61 VSUBS 0.008583f
C226 B.n62 VSUBS 0.008583f
C227 B.n63 VSUBS 0.008583f
C228 B.t2 VSUBS 0.53263f
C229 B.t1 VSUBS 0.565227f
C230 B.t0 VSUBS 2.67905f
C231 B.n64 VSUBS 0.325348f
C232 B.n65 VSUBS 0.0931f
C233 B.n66 VSUBS 0.008583f
C234 B.n67 VSUBS 0.008583f
C235 B.n68 VSUBS 0.008583f
C236 B.n69 VSUBS 0.008583f
C237 B.t11 VSUBS 0.532619f
C238 B.t10 VSUBS 0.565217f
C239 B.t9 VSUBS 2.67905f
C240 B.n70 VSUBS 0.325358f
C241 B.n71 VSUBS 0.093111f
C242 B.n72 VSUBS 0.019887f
C243 B.n73 VSUBS 0.008583f
C244 B.n74 VSUBS 0.008583f
C245 B.n75 VSUBS 0.008583f
C246 B.n76 VSUBS 0.008583f
C247 B.n77 VSUBS 0.008583f
C248 B.n78 VSUBS 0.008583f
C249 B.n79 VSUBS 0.008583f
C250 B.n80 VSUBS 0.008583f
C251 B.n81 VSUBS 0.008583f
C252 B.n82 VSUBS 0.008583f
C253 B.n83 VSUBS 0.008583f
C254 B.n84 VSUBS 0.008583f
C255 B.n85 VSUBS 0.008583f
C256 B.n86 VSUBS 0.008583f
C257 B.n87 VSUBS 0.008583f
C258 B.n88 VSUBS 0.008583f
C259 B.n89 VSUBS 0.008583f
C260 B.n90 VSUBS 0.008583f
C261 B.n91 VSUBS 0.008583f
C262 B.n92 VSUBS 0.008583f
C263 B.n93 VSUBS 0.008583f
C264 B.n94 VSUBS 0.008583f
C265 B.n95 VSUBS 0.019571f
C266 B.n96 VSUBS 0.008583f
C267 B.n97 VSUBS 0.008583f
C268 B.n98 VSUBS 0.008583f
C269 B.n99 VSUBS 0.008583f
C270 B.n100 VSUBS 0.008583f
C271 B.n101 VSUBS 0.008583f
C272 B.n102 VSUBS 0.008583f
C273 B.n103 VSUBS 0.008583f
C274 B.n104 VSUBS 0.008583f
C275 B.n105 VSUBS 0.008583f
C276 B.n106 VSUBS 0.008583f
C277 B.n107 VSUBS 0.008583f
C278 B.n108 VSUBS 0.008583f
C279 B.n109 VSUBS 0.008583f
C280 B.n110 VSUBS 0.008583f
C281 B.n111 VSUBS 0.008583f
C282 B.n112 VSUBS 0.008583f
C283 B.n113 VSUBS 0.008583f
C284 B.n114 VSUBS 0.008583f
C285 B.n115 VSUBS 0.008583f
C286 B.n116 VSUBS 0.008583f
C287 B.n117 VSUBS 0.008583f
C288 B.n118 VSUBS 0.008583f
C289 B.n119 VSUBS 0.008583f
C290 B.n120 VSUBS 0.008583f
C291 B.n121 VSUBS 0.008583f
C292 B.n122 VSUBS 0.008583f
C293 B.n123 VSUBS 0.008583f
C294 B.n124 VSUBS 0.008583f
C295 B.n125 VSUBS 0.008583f
C296 B.n126 VSUBS 0.008583f
C297 B.n127 VSUBS 0.008583f
C298 B.n128 VSUBS 0.008583f
C299 B.n129 VSUBS 0.008583f
C300 B.n130 VSUBS 0.008583f
C301 B.n131 VSUBS 0.008583f
C302 B.n132 VSUBS 0.008583f
C303 B.n133 VSUBS 0.008583f
C304 B.n134 VSUBS 0.008583f
C305 B.n135 VSUBS 0.008583f
C306 B.n136 VSUBS 0.008583f
C307 B.n137 VSUBS 0.008583f
C308 B.n138 VSUBS 0.008583f
C309 B.n139 VSUBS 0.008583f
C310 B.n140 VSUBS 0.008583f
C311 B.n141 VSUBS 0.008583f
C312 B.n142 VSUBS 0.008583f
C313 B.n143 VSUBS 0.008583f
C314 B.n144 VSUBS 0.008583f
C315 B.n145 VSUBS 0.008583f
C316 B.n146 VSUBS 0.008583f
C317 B.n147 VSUBS 0.008583f
C318 B.n148 VSUBS 0.008583f
C319 B.n149 VSUBS 0.008583f
C320 B.n150 VSUBS 0.008583f
C321 B.n151 VSUBS 0.008583f
C322 B.n152 VSUBS 0.008583f
C323 B.n153 VSUBS 0.008583f
C324 B.n154 VSUBS 0.008583f
C325 B.n155 VSUBS 0.008583f
C326 B.n156 VSUBS 0.008583f
C327 B.n157 VSUBS 0.008583f
C328 B.n158 VSUBS 0.008583f
C329 B.n159 VSUBS 0.008583f
C330 B.n160 VSUBS 0.008583f
C331 B.n161 VSUBS 0.008583f
C332 B.n162 VSUBS 0.008583f
C333 B.n163 VSUBS 0.008583f
C334 B.n164 VSUBS 0.008583f
C335 B.n165 VSUBS 0.008583f
C336 B.n166 VSUBS 0.008583f
C337 B.n167 VSUBS 0.008583f
C338 B.n168 VSUBS 0.008583f
C339 B.n169 VSUBS 0.008583f
C340 B.n170 VSUBS 0.008583f
C341 B.n171 VSUBS 0.008583f
C342 B.n172 VSUBS 0.019571f
C343 B.n173 VSUBS 0.008583f
C344 B.n174 VSUBS 0.008583f
C345 B.n175 VSUBS 0.008583f
C346 B.n176 VSUBS 0.008583f
C347 B.n177 VSUBS 0.008583f
C348 B.n178 VSUBS 0.008583f
C349 B.n179 VSUBS 0.008583f
C350 B.n180 VSUBS 0.008583f
C351 B.n181 VSUBS 0.008583f
C352 B.n182 VSUBS 0.008583f
C353 B.n183 VSUBS 0.008583f
C354 B.n184 VSUBS 0.008583f
C355 B.n185 VSUBS 0.008583f
C356 B.n186 VSUBS 0.008583f
C357 B.n187 VSUBS 0.008583f
C358 B.n188 VSUBS 0.008583f
C359 B.n189 VSUBS 0.008583f
C360 B.n190 VSUBS 0.008583f
C361 B.n191 VSUBS 0.008583f
C362 B.n192 VSUBS 0.008583f
C363 B.n193 VSUBS 0.008583f
C364 B.n194 VSUBS 0.008583f
C365 B.n195 VSUBS 0.008583f
C366 B.t7 VSUBS 0.532619f
C367 B.t8 VSUBS 0.565217f
C368 B.t6 VSUBS 2.67905f
C369 B.n196 VSUBS 0.325358f
C370 B.n197 VSUBS 0.093111f
C371 B.n198 VSUBS 0.008583f
C372 B.n199 VSUBS 0.008583f
C373 B.n200 VSUBS 0.008583f
C374 B.n201 VSUBS 0.008583f
C375 B.t4 VSUBS 0.53263f
C376 B.t5 VSUBS 0.565227f
C377 B.t3 VSUBS 2.67905f
C378 B.n202 VSUBS 0.325348f
C379 B.n203 VSUBS 0.0931f
C380 B.n204 VSUBS 0.019887f
C381 B.n205 VSUBS 0.008583f
C382 B.n206 VSUBS 0.008583f
C383 B.n207 VSUBS 0.008583f
C384 B.n208 VSUBS 0.008583f
C385 B.n209 VSUBS 0.008583f
C386 B.n210 VSUBS 0.008583f
C387 B.n211 VSUBS 0.008583f
C388 B.n212 VSUBS 0.008583f
C389 B.n213 VSUBS 0.008583f
C390 B.n214 VSUBS 0.008583f
C391 B.n215 VSUBS 0.008583f
C392 B.n216 VSUBS 0.008583f
C393 B.n217 VSUBS 0.008583f
C394 B.n218 VSUBS 0.008583f
C395 B.n219 VSUBS 0.008583f
C396 B.n220 VSUBS 0.008583f
C397 B.n221 VSUBS 0.008583f
C398 B.n222 VSUBS 0.008583f
C399 B.n223 VSUBS 0.008583f
C400 B.n224 VSUBS 0.008583f
C401 B.n225 VSUBS 0.008583f
C402 B.n226 VSUBS 0.008583f
C403 B.n227 VSUBS 0.019571f
C404 B.n228 VSUBS 0.008583f
C405 B.n229 VSUBS 0.008583f
C406 B.n230 VSUBS 0.008583f
C407 B.n231 VSUBS 0.008583f
C408 B.n232 VSUBS 0.008583f
C409 B.n233 VSUBS 0.008583f
C410 B.n234 VSUBS 0.008583f
C411 B.n235 VSUBS 0.008583f
C412 B.n236 VSUBS 0.008583f
C413 B.n237 VSUBS 0.008583f
C414 B.n238 VSUBS 0.008583f
C415 B.n239 VSUBS 0.008583f
C416 B.n240 VSUBS 0.008583f
C417 B.n241 VSUBS 0.008583f
C418 B.n242 VSUBS 0.008583f
C419 B.n243 VSUBS 0.008583f
C420 B.n244 VSUBS 0.008583f
C421 B.n245 VSUBS 0.008583f
C422 B.n246 VSUBS 0.008583f
C423 B.n247 VSUBS 0.008583f
C424 B.n248 VSUBS 0.008583f
C425 B.n249 VSUBS 0.008583f
C426 B.n250 VSUBS 0.008583f
C427 B.n251 VSUBS 0.008583f
C428 B.n252 VSUBS 0.008583f
C429 B.n253 VSUBS 0.008583f
C430 B.n254 VSUBS 0.008583f
C431 B.n255 VSUBS 0.008583f
C432 B.n256 VSUBS 0.008583f
C433 B.n257 VSUBS 0.008583f
C434 B.n258 VSUBS 0.008583f
C435 B.n259 VSUBS 0.008583f
C436 B.n260 VSUBS 0.008583f
C437 B.n261 VSUBS 0.008583f
C438 B.n262 VSUBS 0.008583f
C439 B.n263 VSUBS 0.008583f
C440 B.n264 VSUBS 0.008583f
C441 B.n265 VSUBS 0.008583f
C442 B.n266 VSUBS 0.008583f
C443 B.n267 VSUBS 0.008583f
C444 B.n268 VSUBS 0.008583f
C445 B.n269 VSUBS 0.008583f
C446 B.n270 VSUBS 0.008583f
C447 B.n271 VSUBS 0.008583f
C448 B.n272 VSUBS 0.008583f
C449 B.n273 VSUBS 0.008583f
C450 B.n274 VSUBS 0.008583f
C451 B.n275 VSUBS 0.008583f
C452 B.n276 VSUBS 0.008583f
C453 B.n277 VSUBS 0.008583f
C454 B.n278 VSUBS 0.008583f
C455 B.n279 VSUBS 0.008583f
C456 B.n280 VSUBS 0.008583f
C457 B.n281 VSUBS 0.008583f
C458 B.n282 VSUBS 0.008583f
C459 B.n283 VSUBS 0.008583f
C460 B.n284 VSUBS 0.008583f
C461 B.n285 VSUBS 0.008583f
C462 B.n286 VSUBS 0.008583f
C463 B.n287 VSUBS 0.008583f
C464 B.n288 VSUBS 0.008583f
C465 B.n289 VSUBS 0.008583f
C466 B.n290 VSUBS 0.008583f
C467 B.n291 VSUBS 0.008583f
C468 B.n292 VSUBS 0.008583f
C469 B.n293 VSUBS 0.008583f
C470 B.n294 VSUBS 0.008583f
C471 B.n295 VSUBS 0.008583f
C472 B.n296 VSUBS 0.008583f
C473 B.n297 VSUBS 0.008583f
C474 B.n298 VSUBS 0.008583f
C475 B.n299 VSUBS 0.008583f
C476 B.n300 VSUBS 0.008583f
C477 B.n301 VSUBS 0.008583f
C478 B.n302 VSUBS 0.008583f
C479 B.n303 VSUBS 0.008583f
C480 B.n304 VSUBS 0.008583f
C481 B.n305 VSUBS 0.008583f
C482 B.n306 VSUBS 0.008583f
C483 B.n307 VSUBS 0.008583f
C484 B.n308 VSUBS 0.008583f
C485 B.n309 VSUBS 0.008583f
C486 B.n310 VSUBS 0.008583f
C487 B.n311 VSUBS 0.008583f
C488 B.n312 VSUBS 0.008583f
C489 B.n313 VSUBS 0.008583f
C490 B.n314 VSUBS 0.008583f
C491 B.n315 VSUBS 0.008583f
C492 B.n316 VSUBS 0.008583f
C493 B.n317 VSUBS 0.008583f
C494 B.n318 VSUBS 0.008583f
C495 B.n319 VSUBS 0.008583f
C496 B.n320 VSUBS 0.008583f
C497 B.n321 VSUBS 0.008583f
C498 B.n322 VSUBS 0.008583f
C499 B.n323 VSUBS 0.008583f
C500 B.n324 VSUBS 0.008583f
C501 B.n325 VSUBS 0.008583f
C502 B.n326 VSUBS 0.008583f
C503 B.n327 VSUBS 0.008583f
C504 B.n328 VSUBS 0.008583f
C505 B.n329 VSUBS 0.008583f
C506 B.n330 VSUBS 0.008583f
C507 B.n331 VSUBS 0.008583f
C508 B.n332 VSUBS 0.008583f
C509 B.n333 VSUBS 0.008583f
C510 B.n334 VSUBS 0.008583f
C511 B.n335 VSUBS 0.008583f
C512 B.n336 VSUBS 0.008583f
C513 B.n337 VSUBS 0.008583f
C514 B.n338 VSUBS 0.008583f
C515 B.n339 VSUBS 0.008583f
C516 B.n340 VSUBS 0.008583f
C517 B.n341 VSUBS 0.008583f
C518 B.n342 VSUBS 0.008583f
C519 B.n343 VSUBS 0.008583f
C520 B.n344 VSUBS 0.008583f
C521 B.n345 VSUBS 0.008583f
C522 B.n346 VSUBS 0.008583f
C523 B.n347 VSUBS 0.008583f
C524 B.n348 VSUBS 0.008583f
C525 B.n349 VSUBS 0.008583f
C526 B.n350 VSUBS 0.008583f
C527 B.n351 VSUBS 0.008583f
C528 B.n352 VSUBS 0.008583f
C529 B.n353 VSUBS 0.008583f
C530 B.n354 VSUBS 0.008583f
C531 B.n355 VSUBS 0.008583f
C532 B.n356 VSUBS 0.008583f
C533 B.n357 VSUBS 0.008583f
C534 B.n358 VSUBS 0.008583f
C535 B.n359 VSUBS 0.008583f
C536 B.n360 VSUBS 0.008583f
C537 B.n361 VSUBS 0.008583f
C538 B.n362 VSUBS 0.008583f
C539 B.n363 VSUBS 0.008583f
C540 B.n364 VSUBS 0.008583f
C541 B.n365 VSUBS 0.008583f
C542 B.n366 VSUBS 0.008583f
C543 B.n367 VSUBS 0.008583f
C544 B.n368 VSUBS 0.008583f
C545 B.n369 VSUBS 0.008583f
C546 B.n370 VSUBS 0.008583f
C547 B.n371 VSUBS 0.008583f
C548 B.n372 VSUBS 0.008583f
C549 B.n373 VSUBS 0.008583f
C550 B.n374 VSUBS 0.008583f
C551 B.n375 VSUBS 0.008583f
C552 B.n376 VSUBS 0.008583f
C553 B.n377 VSUBS 0.008583f
C554 B.n378 VSUBS 0.019571f
C555 B.n379 VSUBS 0.020822f
C556 B.n380 VSUBS 0.020822f
C557 B.n381 VSUBS 0.008583f
C558 B.n382 VSUBS 0.008583f
C559 B.n383 VSUBS 0.008583f
C560 B.n384 VSUBS 0.008583f
C561 B.n385 VSUBS 0.008583f
C562 B.n386 VSUBS 0.008583f
C563 B.n387 VSUBS 0.008583f
C564 B.n388 VSUBS 0.008583f
C565 B.n389 VSUBS 0.008583f
C566 B.n390 VSUBS 0.008583f
C567 B.n391 VSUBS 0.008583f
C568 B.n392 VSUBS 0.008583f
C569 B.n393 VSUBS 0.008583f
C570 B.n394 VSUBS 0.008583f
C571 B.n395 VSUBS 0.008583f
C572 B.n396 VSUBS 0.008583f
C573 B.n397 VSUBS 0.008583f
C574 B.n398 VSUBS 0.008583f
C575 B.n399 VSUBS 0.008583f
C576 B.n400 VSUBS 0.008583f
C577 B.n401 VSUBS 0.008583f
C578 B.n402 VSUBS 0.008583f
C579 B.n403 VSUBS 0.008583f
C580 B.n404 VSUBS 0.008583f
C581 B.n405 VSUBS 0.008583f
C582 B.n406 VSUBS 0.008583f
C583 B.n407 VSUBS 0.008583f
C584 B.n408 VSUBS 0.008583f
C585 B.n409 VSUBS 0.008583f
C586 B.n410 VSUBS 0.008583f
C587 B.n411 VSUBS 0.008583f
C588 B.n412 VSUBS 0.008583f
C589 B.n413 VSUBS 0.008583f
C590 B.n414 VSUBS 0.008583f
C591 B.n415 VSUBS 0.008583f
C592 B.n416 VSUBS 0.008583f
C593 B.n417 VSUBS 0.008583f
C594 B.n418 VSUBS 0.008583f
C595 B.n419 VSUBS 0.008583f
C596 B.n420 VSUBS 0.008583f
C597 B.n421 VSUBS 0.008583f
C598 B.n422 VSUBS 0.008583f
C599 B.n423 VSUBS 0.008583f
C600 B.n424 VSUBS 0.008583f
C601 B.n425 VSUBS 0.008583f
C602 B.n426 VSUBS 0.008583f
C603 B.n427 VSUBS 0.008583f
C604 B.n428 VSUBS 0.008583f
C605 B.n429 VSUBS 0.008583f
C606 B.n430 VSUBS 0.008583f
C607 B.n431 VSUBS 0.008583f
C608 B.n432 VSUBS 0.008583f
C609 B.n433 VSUBS 0.008583f
C610 B.n434 VSUBS 0.008583f
C611 B.n435 VSUBS 0.008583f
C612 B.n436 VSUBS 0.008583f
C613 B.n437 VSUBS 0.008583f
C614 B.n438 VSUBS 0.008583f
C615 B.n439 VSUBS 0.008583f
C616 B.n440 VSUBS 0.008583f
C617 B.n441 VSUBS 0.008583f
C618 B.n442 VSUBS 0.008583f
C619 B.n443 VSUBS 0.008583f
C620 B.n444 VSUBS 0.008583f
C621 B.n445 VSUBS 0.008078f
C622 B.n446 VSUBS 0.008583f
C623 B.n447 VSUBS 0.008583f
C624 B.n448 VSUBS 0.004797f
C625 B.n449 VSUBS 0.008583f
C626 B.n450 VSUBS 0.008583f
C627 B.n451 VSUBS 0.008583f
C628 B.n452 VSUBS 0.008583f
C629 B.n453 VSUBS 0.008583f
C630 B.n454 VSUBS 0.008583f
C631 B.n455 VSUBS 0.008583f
C632 B.n456 VSUBS 0.008583f
C633 B.n457 VSUBS 0.008583f
C634 B.n458 VSUBS 0.008583f
C635 B.n459 VSUBS 0.008583f
C636 B.n460 VSUBS 0.008583f
C637 B.n461 VSUBS 0.004797f
C638 B.n462 VSUBS 0.019887f
C639 B.n463 VSUBS 0.008078f
C640 B.n464 VSUBS 0.008583f
C641 B.n465 VSUBS 0.008583f
C642 B.n466 VSUBS 0.008583f
C643 B.n467 VSUBS 0.008583f
C644 B.n468 VSUBS 0.008583f
C645 B.n469 VSUBS 0.008583f
C646 B.n470 VSUBS 0.008583f
C647 B.n471 VSUBS 0.008583f
C648 B.n472 VSUBS 0.008583f
C649 B.n473 VSUBS 0.008583f
C650 B.n474 VSUBS 0.008583f
C651 B.n475 VSUBS 0.008583f
C652 B.n476 VSUBS 0.008583f
C653 B.n477 VSUBS 0.008583f
C654 B.n478 VSUBS 0.008583f
C655 B.n479 VSUBS 0.008583f
C656 B.n480 VSUBS 0.008583f
C657 B.n481 VSUBS 0.008583f
C658 B.n482 VSUBS 0.008583f
C659 B.n483 VSUBS 0.008583f
C660 B.n484 VSUBS 0.008583f
C661 B.n485 VSUBS 0.008583f
C662 B.n486 VSUBS 0.008583f
C663 B.n487 VSUBS 0.008583f
C664 B.n488 VSUBS 0.008583f
C665 B.n489 VSUBS 0.008583f
C666 B.n490 VSUBS 0.008583f
C667 B.n491 VSUBS 0.008583f
C668 B.n492 VSUBS 0.008583f
C669 B.n493 VSUBS 0.008583f
C670 B.n494 VSUBS 0.008583f
C671 B.n495 VSUBS 0.008583f
C672 B.n496 VSUBS 0.008583f
C673 B.n497 VSUBS 0.008583f
C674 B.n498 VSUBS 0.008583f
C675 B.n499 VSUBS 0.008583f
C676 B.n500 VSUBS 0.008583f
C677 B.n501 VSUBS 0.008583f
C678 B.n502 VSUBS 0.008583f
C679 B.n503 VSUBS 0.008583f
C680 B.n504 VSUBS 0.008583f
C681 B.n505 VSUBS 0.008583f
C682 B.n506 VSUBS 0.008583f
C683 B.n507 VSUBS 0.008583f
C684 B.n508 VSUBS 0.008583f
C685 B.n509 VSUBS 0.008583f
C686 B.n510 VSUBS 0.008583f
C687 B.n511 VSUBS 0.008583f
C688 B.n512 VSUBS 0.008583f
C689 B.n513 VSUBS 0.008583f
C690 B.n514 VSUBS 0.008583f
C691 B.n515 VSUBS 0.008583f
C692 B.n516 VSUBS 0.008583f
C693 B.n517 VSUBS 0.008583f
C694 B.n518 VSUBS 0.008583f
C695 B.n519 VSUBS 0.008583f
C696 B.n520 VSUBS 0.008583f
C697 B.n521 VSUBS 0.008583f
C698 B.n522 VSUBS 0.008583f
C699 B.n523 VSUBS 0.008583f
C700 B.n524 VSUBS 0.008583f
C701 B.n525 VSUBS 0.008583f
C702 B.n526 VSUBS 0.008583f
C703 B.n527 VSUBS 0.008583f
C704 B.n528 VSUBS 0.008583f
C705 B.n529 VSUBS 0.020822f
C706 B.n530 VSUBS 0.020822f
C707 B.n531 VSUBS 0.019571f
C708 B.n532 VSUBS 0.008583f
C709 B.n533 VSUBS 0.008583f
C710 B.n534 VSUBS 0.008583f
C711 B.n535 VSUBS 0.008583f
C712 B.n536 VSUBS 0.008583f
C713 B.n537 VSUBS 0.008583f
C714 B.n538 VSUBS 0.008583f
C715 B.n539 VSUBS 0.008583f
C716 B.n540 VSUBS 0.008583f
C717 B.n541 VSUBS 0.008583f
C718 B.n542 VSUBS 0.008583f
C719 B.n543 VSUBS 0.008583f
C720 B.n544 VSUBS 0.008583f
C721 B.n545 VSUBS 0.008583f
C722 B.n546 VSUBS 0.008583f
C723 B.n547 VSUBS 0.008583f
C724 B.n548 VSUBS 0.008583f
C725 B.n549 VSUBS 0.008583f
C726 B.n550 VSUBS 0.008583f
C727 B.n551 VSUBS 0.008583f
C728 B.n552 VSUBS 0.008583f
C729 B.n553 VSUBS 0.008583f
C730 B.n554 VSUBS 0.008583f
C731 B.n555 VSUBS 0.008583f
C732 B.n556 VSUBS 0.008583f
C733 B.n557 VSUBS 0.008583f
C734 B.n558 VSUBS 0.008583f
C735 B.n559 VSUBS 0.008583f
C736 B.n560 VSUBS 0.008583f
C737 B.n561 VSUBS 0.008583f
C738 B.n562 VSUBS 0.008583f
C739 B.n563 VSUBS 0.008583f
C740 B.n564 VSUBS 0.008583f
C741 B.n565 VSUBS 0.008583f
C742 B.n566 VSUBS 0.008583f
C743 B.n567 VSUBS 0.008583f
C744 B.n568 VSUBS 0.008583f
C745 B.n569 VSUBS 0.008583f
C746 B.n570 VSUBS 0.008583f
C747 B.n571 VSUBS 0.008583f
C748 B.n572 VSUBS 0.008583f
C749 B.n573 VSUBS 0.008583f
C750 B.n574 VSUBS 0.008583f
C751 B.n575 VSUBS 0.008583f
C752 B.n576 VSUBS 0.008583f
C753 B.n577 VSUBS 0.008583f
C754 B.n578 VSUBS 0.008583f
C755 B.n579 VSUBS 0.008583f
C756 B.n580 VSUBS 0.008583f
C757 B.n581 VSUBS 0.008583f
C758 B.n582 VSUBS 0.008583f
C759 B.n583 VSUBS 0.008583f
C760 B.n584 VSUBS 0.008583f
C761 B.n585 VSUBS 0.008583f
C762 B.n586 VSUBS 0.008583f
C763 B.n587 VSUBS 0.008583f
C764 B.n588 VSUBS 0.008583f
C765 B.n589 VSUBS 0.008583f
C766 B.n590 VSUBS 0.008583f
C767 B.n591 VSUBS 0.008583f
C768 B.n592 VSUBS 0.008583f
C769 B.n593 VSUBS 0.008583f
C770 B.n594 VSUBS 0.008583f
C771 B.n595 VSUBS 0.008583f
C772 B.n596 VSUBS 0.008583f
C773 B.n597 VSUBS 0.008583f
C774 B.n598 VSUBS 0.008583f
C775 B.n599 VSUBS 0.008583f
C776 B.n600 VSUBS 0.008583f
C777 B.n601 VSUBS 0.008583f
C778 B.n602 VSUBS 0.008583f
C779 B.n603 VSUBS 0.008583f
C780 B.n604 VSUBS 0.008583f
C781 B.n605 VSUBS 0.008583f
C782 B.n606 VSUBS 0.008583f
C783 B.n607 VSUBS 0.008583f
C784 B.n608 VSUBS 0.008583f
C785 B.n609 VSUBS 0.008583f
C786 B.n610 VSUBS 0.008583f
C787 B.n611 VSUBS 0.008583f
C788 B.n612 VSUBS 0.008583f
C789 B.n613 VSUBS 0.008583f
C790 B.n614 VSUBS 0.008583f
C791 B.n615 VSUBS 0.008583f
C792 B.n616 VSUBS 0.008583f
C793 B.n617 VSUBS 0.008583f
C794 B.n618 VSUBS 0.008583f
C795 B.n619 VSUBS 0.008583f
C796 B.n620 VSUBS 0.008583f
C797 B.n621 VSUBS 0.008583f
C798 B.n622 VSUBS 0.008583f
C799 B.n623 VSUBS 0.008583f
C800 B.n624 VSUBS 0.008583f
C801 B.n625 VSUBS 0.008583f
C802 B.n626 VSUBS 0.008583f
C803 B.n627 VSUBS 0.008583f
C804 B.n628 VSUBS 0.008583f
C805 B.n629 VSUBS 0.008583f
C806 B.n630 VSUBS 0.008583f
C807 B.n631 VSUBS 0.008583f
C808 B.n632 VSUBS 0.008583f
C809 B.n633 VSUBS 0.008583f
C810 B.n634 VSUBS 0.008583f
C811 B.n635 VSUBS 0.008583f
C812 B.n636 VSUBS 0.008583f
C813 B.n637 VSUBS 0.008583f
C814 B.n638 VSUBS 0.008583f
C815 B.n639 VSUBS 0.008583f
C816 B.n640 VSUBS 0.008583f
C817 B.n641 VSUBS 0.008583f
C818 B.n642 VSUBS 0.008583f
C819 B.n643 VSUBS 0.008583f
C820 B.n644 VSUBS 0.008583f
C821 B.n645 VSUBS 0.008583f
C822 B.n646 VSUBS 0.008583f
C823 B.n647 VSUBS 0.008583f
C824 B.n648 VSUBS 0.008583f
C825 B.n649 VSUBS 0.008583f
C826 B.n650 VSUBS 0.008583f
C827 B.n651 VSUBS 0.008583f
C828 B.n652 VSUBS 0.008583f
C829 B.n653 VSUBS 0.008583f
C830 B.n654 VSUBS 0.008583f
C831 B.n655 VSUBS 0.008583f
C832 B.n656 VSUBS 0.008583f
C833 B.n657 VSUBS 0.008583f
C834 B.n658 VSUBS 0.008583f
C835 B.n659 VSUBS 0.008583f
C836 B.n660 VSUBS 0.008583f
C837 B.n661 VSUBS 0.008583f
C838 B.n662 VSUBS 0.008583f
C839 B.n663 VSUBS 0.008583f
C840 B.n664 VSUBS 0.008583f
C841 B.n665 VSUBS 0.008583f
C842 B.n666 VSUBS 0.008583f
C843 B.n667 VSUBS 0.008583f
C844 B.n668 VSUBS 0.008583f
C845 B.n669 VSUBS 0.008583f
C846 B.n670 VSUBS 0.008583f
C847 B.n671 VSUBS 0.008583f
C848 B.n672 VSUBS 0.008583f
C849 B.n673 VSUBS 0.008583f
C850 B.n674 VSUBS 0.008583f
C851 B.n675 VSUBS 0.008583f
C852 B.n676 VSUBS 0.008583f
C853 B.n677 VSUBS 0.008583f
C854 B.n678 VSUBS 0.008583f
C855 B.n679 VSUBS 0.008583f
C856 B.n680 VSUBS 0.008583f
C857 B.n681 VSUBS 0.008583f
C858 B.n682 VSUBS 0.008583f
C859 B.n683 VSUBS 0.008583f
C860 B.n684 VSUBS 0.008583f
C861 B.n685 VSUBS 0.008583f
C862 B.n686 VSUBS 0.008583f
C863 B.n687 VSUBS 0.008583f
C864 B.n688 VSUBS 0.008583f
C865 B.n689 VSUBS 0.008583f
C866 B.n690 VSUBS 0.008583f
C867 B.n691 VSUBS 0.008583f
C868 B.n692 VSUBS 0.008583f
C869 B.n693 VSUBS 0.008583f
C870 B.n694 VSUBS 0.008583f
C871 B.n695 VSUBS 0.008583f
C872 B.n696 VSUBS 0.008583f
C873 B.n697 VSUBS 0.008583f
C874 B.n698 VSUBS 0.008583f
C875 B.n699 VSUBS 0.008583f
C876 B.n700 VSUBS 0.008583f
C877 B.n701 VSUBS 0.008583f
C878 B.n702 VSUBS 0.008583f
C879 B.n703 VSUBS 0.008583f
C880 B.n704 VSUBS 0.008583f
C881 B.n705 VSUBS 0.008583f
C882 B.n706 VSUBS 0.008583f
C883 B.n707 VSUBS 0.008583f
C884 B.n708 VSUBS 0.008583f
C885 B.n709 VSUBS 0.008583f
C886 B.n710 VSUBS 0.008583f
C887 B.n711 VSUBS 0.008583f
C888 B.n712 VSUBS 0.008583f
C889 B.n713 VSUBS 0.008583f
C890 B.n714 VSUBS 0.008583f
C891 B.n715 VSUBS 0.008583f
C892 B.n716 VSUBS 0.008583f
C893 B.n717 VSUBS 0.008583f
C894 B.n718 VSUBS 0.008583f
C895 B.n719 VSUBS 0.008583f
C896 B.n720 VSUBS 0.008583f
C897 B.n721 VSUBS 0.008583f
C898 B.n722 VSUBS 0.008583f
C899 B.n723 VSUBS 0.008583f
C900 B.n724 VSUBS 0.008583f
C901 B.n725 VSUBS 0.008583f
C902 B.n726 VSUBS 0.008583f
C903 B.n727 VSUBS 0.008583f
C904 B.n728 VSUBS 0.008583f
C905 B.n729 VSUBS 0.008583f
C906 B.n730 VSUBS 0.008583f
C907 B.n731 VSUBS 0.008583f
C908 B.n732 VSUBS 0.008583f
C909 B.n733 VSUBS 0.008583f
C910 B.n734 VSUBS 0.008583f
C911 B.n735 VSUBS 0.008583f
C912 B.n736 VSUBS 0.008583f
C913 B.n737 VSUBS 0.008583f
C914 B.n738 VSUBS 0.008583f
C915 B.n739 VSUBS 0.008583f
C916 B.n740 VSUBS 0.008583f
C917 B.n741 VSUBS 0.008583f
C918 B.n742 VSUBS 0.008583f
C919 B.n743 VSUBS 0.008583f
C920 B.n744 VSUBS 0.008583f
C921 B.n745 VSUBS 0.008583f
C922 B.n746 VSUBS 0.008583f
C923 B.n747 VSUBS 0.008583f
C924 B.n748 VSUBS 0.008583f
C925 B.n749 VSUBS 0.008583f
C926 B.n750 VSUBS 0.008583f
C927 B.n751 VSUBS 0.008583f
C928 B.n752 VSUBS 0.008583f
C929 B.n753 VSUBS 0.008583f
C930 B.n754 VSUBS 0.008583f
C931 B.n755 VSUBS 0.008583f
C932 B.n756 VSUBS 0.008583f
C933 B.n757 VSUBS 0.008583f
C934 B.n758 VSUBS 0.008583f
C935 B.n759 VSUBS 0.008583f
C936 B.n760 VSUBS 0.008583f
C937 B.n761 VSUBS 0.008583f
C938 B.n762 VSUBS 0.020576f
C939 B.n763 VSUBS 0.019816f
C940 B.n764 VSUBS 0.020822f
C941 B.n765 VSUBS 0.008583f
C942 B.n766 VSUBS 0.008583f
C943 B.n767 VSUBS 0.008583f
C944 B.n768 VSUBS 0.008583f
C945 B.n769 VSUBS 0.008583f
C946 B.n770 VSUBS 0.008583f
C947 B.n771 VSUBS 0.008583f
C948 B.n772 VSUBS 0.008583f
C949 B.n773 VSUBS 0.008583f
C950 B.n774 VSUBS 0.008583f
C951 B.n775 VSUBS 0.008583f
C952 B.n776 VSUBS 0.008583f
C953 B.n777 VSUBS 0.008583f
C954 B.n778 VSUBS 0.008583f
C955 B.n779 VSUBS 0.008583f
C956 B.n780 VSUBS 0.008583f
C957 B.n781 VSUBS 0.008583f
C958 B.n782 VSUBS 0.008583f
C959 B.n783 VSUBS 0.008583f
C960 B.n784 VSUBS 0.008583f
C961 B.n785 VSUBS 0.008583f
C962 B.n786 VSUBS 0.008583f
C963 B.n787 VSUBS 0.008583f
C964 B.n788 VSUBS 0.008583f
C965 B.n789 VSUBS 0.008583f
C966 B.n790 VSUBS 0.008583f
C967 B.n791 VSUBS 0.008583f
C968 B.n792 VSUBS 0.008583f
C969 B.n793 VSUBS 0.008583f
C970 B.n794 VSUBS 0.008583f
C971 B.n795 VSUBS 0.008583f
C972 B.n796 VSUBS 0.008583f
C973 B.n797 VSUBS 0.008583f
C974 B.n798 VSUBS 0.008583f
C975 B.n799 VSUBS 0.008583f
C976 B.n800 VSUBS 0.008583f
C977 B.n801 VSUBS 0.008583f
C978 B.n802 VSUBS 0.008583f
C979 B.n803 VSUBS 0.008583f
C980 B.n804 VSUBS 0.008583f
C981 B.n805 VSUBS 0.008583f
C982 B.n806 VSUBS 0.008583f
C983 B.n807 VSUBS 0.008583f
C984 B.n808 VSUBS 0.008583f
C985 B.n809 VSUBS 0.008583f
C986 B.n810 VSUBS 0.008583f
C987 B.n811 VSUBS 0.008583f
C988 B.n812 VSUBS 0.008583f
C989 B.n813 VSUBS 0.008583f
C990 B.n814 VSUBS 0.008583f
C991 B.n815 VSUBS 0.008583f
C992 B.n816 VSUBS 0.008583f
C993 B.n817 VSUBS 0.008583f
C994 B.n818 VSUBS 0.008583f
C995 B.n819 VSUBS 0.008583f
C996 B.n820 VSUBS 0.008583f
C997 B.n821 VSUBS 0.008583f
C998 B.n822 VSUBS 0.008583f
C999 B.n823 VSUBS 0.008583f
C1000 B.n824 VSUBS 0.008583f
C1001 B.n825 VSUBS 0.008583f
C1002 B.n826 VSUBS 0.008583f
C1003 B.n827 VSUBS 0.008583f
C1004 B.n828 VSUBS 0.008583f
C1005 B.n829 VSUBS 0.008078f
C1006 B.n830 VSUBS 0.008583f
C1007 B.n831 VSUBS 0.008583f
C1008 B.n832 VSUBS 0.004797f
C1009 B.n833 VSUBS 0.008583f
C1010 B.n834 VSUBS 0.008583f
C1011 B.n835 VSUBS 0.008583f
C1012 B.n836 VSUBS 0.008583f
C1013 B.n837 VSUBS 0.008583f
C1014 B.n838 VSUBS 0.008583f
C1015 B.n839 VSUBS 0.008583f
C1016 B.n840 VSUBS 0.008583f
C1017 B.n841 VSUBS 0.008583f
C1018 B.n842 VSUBS 0.008583f
C1019 B.n843 VSUBS 0.008583f
C1020 B.n844 VSUBS 0.008583f
C1021 B.n845 VSUBS 0.004797f
C1022 B.n846 VSUBS 0.019887f
C1023 B.n847 VSUBS 0.008078f
C1024 B.n848 VSUBS 0.008583f
C1025 B.n849 VSUBS 0.008583f
C1026 B.n850 VSUBS 0.008583f
C1027 B.n851 VSUBS 0.008583f
C1028 B.n852 VSUBS 0.008583f
C1029 B.n853 VSUBS 0.008583f
C1030 B.n854 VSUBS 0.008583f
C1031 B.n855 VSUBS 0.008583f
C1032 B.n856 VSUBS 0.008583f
C1033 B.n857 VSUBS 0.008583f
C1034 B.n858 VSUBS 0.008583f
C1035 B.n859 VSUBS 0.008583f
C1036 B.n860 VSUBS 0.008583f
C1037 B.n861 VSUBS 0.008583f
C1038 B.n862 VSUBS 0.008583f
C1039 B.n863 VSUBS 0.008583f
C1040 B.n864 VSUBS 0.008583f
C1041 B.n865 VSUBS 0.008583f
C1042 B.n866 VSUBS 0.008583f
C1043 B.n867 VSUBS 0.008583f
C1044 B.n868 VSUBS 0.008583f
C1045 B.n869 VSUBS 0.008583f
C1046 B.n870 VSUBS 0.008583f
C1047 B.n871 VSUBS 0.008583f
C1048 B.n872 VSUBS 0.008583f
C1049 B.n873 VSUBS 0.008583f
C1050 B.n874 VSUBS 0.008583f
C1051 B.n875 VSUBS 0.008583f
C1052 B.n876 VSUBS 0.008583f
C1053 B.n877 VSUBS 0.008583f
C1054 B.n878 VSUBS 0.008583f
C1055 B.n879 VSUBS 0.008583f
C1056 B.n880 VSUBS 0.008583f
C1057 B.n881 VSUBS 0.008583f
C1058 B.n882 VSUBS 0.008583f
C1059 B.n883 VSUBS 0.008583f
C1060 B.n884 VSUBS 0.008583f
C1061 B.n885 VSUBS 0.008583f
C1062 B.n886 VSUBS 0.008583f
C1063 B.n887 VSUBS 0.008583f
C1064 B.n888 VSUBS 0.008583f
C1065 B.n889 VSUBS 0.008583f
C1066 B.n890 VSUBS 0.008583f
C1067 B.n891 VSUBS 0.008583f
C1068 B.n892 VSUBS 0.008583f
C1069 B.n893 VSUBS 0.008583f
C1070 B.n894 VSUBS 0.008583f
C1071 B.n895 VSUBS 0.008583f
C1072 B.n896 VSUBS 0.008583f
C1073 B.n897 VSUBS 0.008583f
C1074 B.n898 VSUBS 0.008583f
C1075 B.n899 VSUBS 0.008583f
C1076 B.n900 VSUBS 0.008583f
C1077 B.n901 VSUBS 0.008583f
C1078 B.n902 VSUBS 0.008583f
C1079 B.n903 VSUBS 0.008583f
C1080 B.n904 VSUBS 0.008583f
C1081 B.n905 VSUBS 0.008583f
C1082 B.n906 VSUBS 0.008583f
C1083 B.n907 VSUBS 0.008583f
C1084 B.n908 VSUBS 0.008583f
C1085 B.n909 VSUBS 0.008583f
C1086 B.n910 VSUBS 0.008583f
C1087 B.n911 VSUBS 0.008583f
C1088 B.n912 VSUBS 0.008583f
C1089 B.n913 VSUBS 0.020822f
C1090 B.n914 VSUBS 0.020822f
C1091 B.n915 VSUBS 0.019571f
C1092 B.n916 VSUBS 0.008583f
C1093 B.n917 VSUBS 0.008583f
C1094 B.n918 VSUBS 0.008583f
C1095 B.n919 VSUBS 0.008583f
C1096 B.n920 VSUBS 0.008583f
C1097 B.n921 VSUBS 0.008583f
C1098 B.n922 VSUBS 0.008583f
C1099 B.n923 VSUBS 0.008583f
C1100 B.n924 VSUBS 0.008583f
C1101 B.n925 VSUBS 0.008583f
C1102 B.n926 VSUBS 0.008583f
C1103 B.n927 VSUBS 0.008583f
C1104 B.n928 VSUBS 0.008583f
C1105 B.n929 VSUBS 0.008583f
C1106 B.n930 VSUBS 0.008583f
C1107 B.n931 VSUBS 0.008583f
C1108 B.n932 VSUBS 0.008583f
C1109 B.n933 VSUBS 0.008583f
C1110 B.n934 VSUBS 0.008583f
C1111 B.n935 VSUBS 0.008583f
C1112 B.n936 VSUBS 0.008583f
C1113 B.n937 VSUBS 0.008583f
C1114 B.n938 VSUBS 0.008583f
C1115 B.n939 VSUBS 0.008583f
C1116 B.n940 VSUBS 0.008583f
C1117 B.n941 VSUBS 0.008583f
C1118 B.n942 VSUBS 0.008583f
C1119 B.n943 VSUBS 0.008583f
C1120 B.n944 VSUBS 0.008583f
C1121 B.n945 VSUBS 0.008583f
C1122 B.n946 VSUBS 0.008583f
C1123 B.n947 VSUBS 0.008583f
C1124 B.n948 VSUBS 0.008583f
C1125 B.n949 VSUBS 0.008583f
C1126 B.n950 VSUBS 0.008583f
C1127 B.n951 VSUBS 0.008583f
C1128 B.n952 VSUBS 0.008583f
C1129 B.n953 VSUBS 0.008583f
C1130 B.n954 VSUBS 0.008583f
C1131 B.n955 VSUBS 0.008583f
C1132 B.n956 VSUBS 0.008583f
C1133 B.n957 VSUBS 0.008583f
C1134 B.n958 VSUBS 0.008583f
C1135 B.n959 VSUBS 0.008583f
C1136 B.n960 VSUBS 0.008583f
C1137 B.n961 VSUBS 0.008583f
C1138 B.n962 VSUBS 0.008583f
C1139 B.n963 VSUBS 0.008583f
C1140 B.n964 VSUBS 0.008583f
C1141 B.n965 VSUBS 0.008583f
C1142 B.n966 VSUBS 0.008583f
C1143 B.n967 VSUBS 0.008583f
C1144 B.n968 VSUBS 0.008583f
C1145 B.n969 VSUBS 0.008583f
C1146 B.n970 VSUBS 0.008583f
C1147 B.n971 VSUBS 0.008583f
C1148 B.n972 VSUBS 0.008583f
C1149 B.n973 VSUBS 0.008583f
C1150 B.n974 VSUBS 0.008583f
C1151 B.n975 VSUBS 0.008583f
C1152 B.n976 VSUBS 0.008583f
C1153 B.n977 VSUBS 0.008583f
C1154 B.n978 VSUBS 0.008583f
C1155 B.n979 VSUBS 0.008583f
C1156 B.n980 VSUBS 0.008583f
C1157 B.n981 VSUBS 0.008583f
C1158 B.n982 VSUBS 0.008583f
C1159 B.n983 VSUBS 0.008583f
C1160 B.n984 VSUBS 0.008583f
C1161 B.n985 VSUBS 0.008583f
C1162 B.n986 VSUBS 0.008583f
C1163 B.n987 VSUBS 0.008583f
C1164 B.n988 VSUBS 0.008583f
C1165 B.n989 VSUBS 0.008583f
C1166 B.n990 VSUBS 0.008583f
C1167 B.n991 VSUBS 0.008583f
C1168 B.n992 VSUBS 0.008583f
C1169 B.n993 VSUBS 0.008583f
C1170 B.n994 VSUBS 0.008583f
C1171 B.n995 VSUBS 0.008583f
C1172 B.n996 VSUBS 0.008583f
C1173 B.n997 VSUBS 0.008583f
C1174 B.n998 VSUBS 0.008583f
C1175 B.n999 VSUBS 0.008583f
C1176 B.n1000 VSUBS 0.008583f
C1177 B.n1001 VSUBS 0.008583f
C1178 B.n1002 VSUBS 0.008583f
C1179 B.n1003 VSUBS 0.008583f
C1180 B.n1004 VSUBS 0.008583f
C1181 B.n1005 VSUBS 0.008583f
C1182 B.n1006 VSUBS 0.008583f
C1183 B.n1007 VSUBS 0.008583f
C1184 B.n1008 VSUBS 0.008583f
C1185 B.n1009 VSUBS 0.008583f
C1186 B.n1010 VSUBS 0.008583f
C1187 B.n1011 VSUBS 0.008583f
C1188 B.n1012 VSUBS 0.008583f
C1189 B.n1013 VSUBS 0.008583f
C1190 B.n1014 VSUBS 0.008583f
C1191 B.n1015 VSUBS 0.008583f
C1192 B.n1016 VSUBS 0.008583f
C1193 B.n1017 VSUBS 0.008583f
C1194 B.n1018 VSUBS 0.008583f
C1195 B.n1019 VSUBS 0.008583f
C1196 B.n1020 VSUBS 0.008583f
C1197 B.n1021 VSUBS 0.008583f
C1198 B.n1022 VSUBS 0.008583f
C1199 B.n1023 VSUBS 0.008583f
C1200 B.n1024 VSUBS 0.008583f
C1201 B.n1025 VSUBS 0.008583f
C1202 B.n1026 VSUBS 0.008583f
C1203 B.n1027 VSUBS 0.008583f
C1204 B.n1028 VSUBS 0.008583f
C1205 B.n1029 VSUBS 0.008583f
C1206 B.n1030 VSUBS 0.008583f
C1207 B.n1031 VSUBS 0.019436f
C1208 VDD1.t9 VSUBS 3.33125f
C1209 VDD1.t6 VSUBS 0.318058f
C1210 VDD1.t4 VSUBS 0.318058f
C1211 VDD1.n0 VSUBS 2.52033f
C1212 VDD1.n1 VSUBS 1.98689f
C1213 VDD1.t7 VSUBS 3.33125f
C1214 VDD1.t5 VSUBS 0.318058f
C1215 VDD1.t2 VSUBS 0.318058f
C1216 VDD1.n2 VSUBS 2.52033f
C1217 VDD1.n3 VSUBS 1.97665f
C1218 VDD1.t1 VSUBS 0.318058f
C1219 VDD1.t3 VSUBS 0.318058f
C1220 VDD1.n4 VSUBS 2.55886f
C1221 VDD1.n5 VSUBS 4.76936f
C1222 VDD1.t0 VSUBS 0.318058f
C1223 VDD1.t8 VSUBS 0.318058f
C1224 VDD1.n6 VSUBS 2.52032f
C1225 VDD1.n7 VSUBS 4.80911f
C1226 VTAIL.t2 VSUBS 0.30647f
C1227 VTAIL.t1 VSUBS 0.30647f
C1228 VTAIL.n0 VSUBS 2.26254f
C1229 VTAIL.n1 VSUBS 1.13726f
C1230 VTAIL.t10 VSUBS 2.98068f
C1231 VTAIL.n2 VSUBS 1.32922f
C1232 VTAIL.t9 VSUBS 0.30647f
C1233 VTAIL.t11 VSUBS 0.30647f
C1234 VTAIL.n3 VSUBS 2.26254f
C1235 VTAIL.n4 VSUBS 1.3266f
C1236 VTAIL.t13 VSUBS 0.30647f
C1237 VTAIL.t14 VSUBS 0.30647f
C1238 VTAIL.n5 VSUBS 2.26254f
C1239 VTAIL.n6 VSUBS 3.12209f
C1240 VTAIL.t0 VSUBS 0.30647f
C1241 VTAIL.t5 VSUBS 0.30647f
C1242 VTAIL.n7 VSUBS 2.26255f
C1243 VTAIL.n8 VSUBS 3.12209f
C1244 VTAIL.t4 VSUBS 0.30647f
C1245 VTAIL.t3 VSUBS 0.30647f
C1246 VTAIL.n9 VSUBS 2.26255f
C1247 VTAIL.n10 VSUBS 1.32659f
C1248 VTAIL.t6 VSUBS 2.98069f
C1249 VTAIL.n11 VSUBS 1.32921f
C1250 VTAIL.t7 VSUBS 0.30647f
C1251 VTAIL.t16 VSUBS 0.30647f
C1252 VTAIL.n12 VSUBS 2.26255f
C1253 VTAIL.n13 VSUBS 1.21152f
C1254 VTAIL.t12 VSUBS 0.30647f
C1255 VTAIL.t15 VSUBS 0.30647f
C1256 VTAIL.n14 VSUBS 2.26255f
C1257 VTAIL.n15 VSUBS 1.32659f
C1258 VTAIL.t8 VSUBS 2.98068f
C1259 VTAIL.n16 VSUBS 2.92068f
C1260 VTAIL.t17 VSUBS 2.98068f
C1261 VTAIL.n17 VSUBS 2.92068f
C1262 VTAIL.t18 VSUBS 0.30647f
C1263 VTAIL.t19 VSUBS 0.30647f
C1264 VTAIL.n18 VSUBS 2.26254f
C1265 VTAIL.n19 VSUBS 1.08176f
C1266 VP.t6 VSUBS 3.25008f
C1267 VP.n0 VSUBS 1.22386f
C1268 VP.n1 VSUBS 0.025177f
C1269 VP.n2 VSUBS 0.045238f
C1270 VP.n3 VSUBS 0.025177f
C1271 VP.n4 VSUBS 0.039313f
C1272 VP.n5 VSUBS 0.025177f
C1273 VP.n6 VSUBS 0.039733f
C1274 VP.n7 VSUBS 0.025177f
C1275 VP.n8 VSUBS 0.035164f
C1276 VP.n9 VSUBS 0.025177f
C1277 VP.n10 VSUBS 0.033464f
C1278 VP.n11 VSUBS 0.025177f
C1279 VP.n12 VSUBS 0.031015f
C1280 VP.n13 VSUBS 0.025177f
C1281 VP.n14 VSUBS 0.024925f
C1282 VP.n15 VSUBS 0.025177f
C1283 VP.n16 VSUBS 0.026867f
C1284 VP.t1 VSUBS 3.25008f
C1285 VP.n17 VSUBS 1.22386f
C1286 VP.n18 VSUBS 0.025177f
C1287 VP.n19 VSUBS 0.045238f
C1288 VP.n20 VSUBS 0.025177f
C1289 VP.n21 VSUBS 0.039313f
C1290 VP.n22 VSUBS 0.025177f
C1291 VP.n23 VSUBS 0.039733f
C1292 VP.n24 VSUBS 0.025177f
C1293 VP.n25 VSUBS 0.035164f
C1294 VP.n26 VSUBS 0.025177f
C1295 VP.n27 VSUBS 0.033464f
C1296 VP.n28 VSUBS 0.025177f
C1297 VP.n29 VSUBS 0.031015f
C1298 VP.t0 VSUBS 3.60097f
C1299 VP.t3 VSUBS 3.25008f
C1300 VP.n30 VSUBS 1.21746f
C1301 VP.n31 VSUBS 1.16366f
C1302 VP.n32 VSUBS 0.315596f
C1303 VP.n33 VSUBS 0.025177f
C1304 VP.n34 VSUBS 0.046689f
C1305 VP.n35 VSUBS 0.046689f
C1306 VP.n36 VSUBS 0.039733f
C1307 VP.n37 VSUBS 0.025177f
C1308 VP.n38 VSUBS 0.025177f
C1309 VP.n39 VSUBS 0.025177f
C1310 VP.n40 VSUBS 0.046689f
C1311 VP.n41 VSUBS 0.046689f
C1312 VP.t5 VSUBS 3.25008f
C1313 VP.n42 VSUBS 1.13448f
C1314 VP.n43 VSUBS 0.035164f
C1315 VP.n44 VSUBS 0.025177f
C1316 VP.n45 VSUBS 0.025177f
C1317 VP.n46 VSUBS 0.025177f
C1318 VP.n47 VSUBS 0.046689f
C1319 VP.n48 VSUBS 0.046689f
C1320 VP.n49 VSUBS 0.033464f
C1321 VP.n50 VSUBS 0.025177f
C1322 VP.n51 VSUBS 0.025177f
C1323 VP.n52 VSUBS 0.025177f
C1324 VP.n53 VSUBS 0.046689f
C1325 VP.n54 VSUBS 0.046689f
C1326 VP.t9 VSUBS 3.25008f
C1327 VP.n55 VSUBS 1.13448f
C1328 VP.n56 VSUBS 0.031015f
C1329 VP.n57 VSUBS 0.025177f
C1330 VP.n58 VSUBS 0.025177f
C1331 VP.n59 VSUBS 0.025177f
C1332 VP.n60 VSUBS 0.046689f
C1333 VP.n61 VSUBS 0.049723f
C1334 VP.n62 VSUBS 0.024925f
C1335 VP.n63 VSUBS 0.025177f
C1336 VP.n64 VSUBS 0.025177f
C1337 VP.n65 VSUBS 0.025177f
C1338 VP.n66 VSUBS 0.046689f
C1339 VP.n67 VSUBS 0.046689f
C1340 VP.n68 VSUBS 0.026867f
C1341 VP.n69 VSUBS 0.040629f
C1342 VP.n70 VSUBS 1.82859f
C1343 VP.t2 VSUBS 3.25008f
C1344 VP.n71 VSUBS 1.22386f
C1345 VP.n72 VSUBS 1.84388f
C1346 VP.n73 VSUBS 0.040629f
C1347 VP.n74 VSUBS 0.025177f
C1348 VP.n75 VSUBS 0.046689f
C1349 VP.n76 VSUBS 0.046689f
C1350 VP.n77 VSUBS 0.045238f
C1351 VP.n78 VSUBS 0.025177f
C1352 VP.n79 VSUBS 0.025177f
C1353 VP.n80 VSUBS 0.025177f
C1354 VP.n81 VSUBS 0.049723f
C1355 VP.n82 VSUBS 0.046689f
C1356 VP.t4 VSUBS 3.25008f
C1357 VP.n83 VSUBS 1.13448f
C1358 VP.n84 VSUBS 0.039313f
C1359 VP.n85 VSUBS 0.025177f
C1360 VP.n86 VSUBS 0.025177f
C1361 VP.n87 VSUBS 0.025177f
C1362 VP.n88 VSUBS 0.046689f
C1363 VP.n89 VSUBS 0.046689f
C1364 VP.n90 VSUBS 0.039733f
C1365 VP.n91 VSUBS 0.025177f
C1366 VP.n92 VSUBS 0.025177f
C1367 VP.n93 VSUBS 0.025177f
C1368 VP.n94 VSUBS 0.046689f
C1369 VP.n95 VSUBS 0.046689f
C1370 VP.t7 VSUBS 3.25008f
C1371 VP.n96 VSUBS 1.13448f
C1372 VP.n97 VSUBS 0.035164f
C1373 VP.n98 VSUBS 0.025177f
C1374 VP.n99 VSUBS 0.025177f
C1375 VP.n100 VSUBS 0.025177f
C1376 VP.n101 VSUBS 0.046689f
C1377 VP.n102 VSUBS 0.046689f
C1378 VP.n103 VSUBS 0.033464f
C1379 VP.n104 VSUBS 0.025177f
C1380 VP.n105 VSUBS 0.025177f
C1381 VP.n106 VSUBS 0.025177f
C1382 VP.n107 VSUBS 0.046689f
C1383 VP.n108 VSUBS 0.046689f
C1384 VP.t8 VSUBS 3.25008f
C1385 VP.n109 VSUBS 1.13448f
C1386 VP.n110 VSUBS 0.031015f
C1387 VP.n111 VSUBS 0.025177f
C1388 VP.n112 VSUBS 0.025177f
C1389 VP.n113 VSUBS 0.025177f
C1390 VP.n114 VSUBS 0.046689f
C1391 VP.n115 VSUBS 0.049723f
C1392 VP.n116 VSUBS 0.024925f
C1393 VP.n117 VSUBS 0.025177f
C1394 VP.n118 VSUBS 0.025177f
C1395 VP.n119 VSUBS 0.025177f
C1396 VP.n120 VSUBS 0.046689f
C1397 VP.n121 VSUBS 0.046689f
C1398 VP.n122 VSUBS 0.026867f
C1399 VP.n123 VSUBS 0.040629f
C1400 VP.n124 VSUBS 0.073784f
.ends

