* NGSPICE file created from diff_pair_sample_1591.ext - technology: sky130A

.subckt diff_pair_sample_1591 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t9 VP.t0 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.60865 pd=16.14 as=2.60865 ps=16.14 w=15.81 l=2.54
X1 VDD2.t5 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.60865 pd=16.14 as=6.1659 ps=32.4 w=15.81 l=2.54
X2 VTAIL.t2 VN.t1 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=2.60865 pd=16.14 as=2.60865 ps=16.14 w=15.81 l=2.54
X3 VTAIL.t8 VP.t1 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.60865 pd=16.14 as=2.60865 ps=16.14 w=15.81 l=2.54
X4 VDD1.t1 VP.t2 VTAIL.t7 B.t19 sky130_fd_pr__nfet_01v8 ad=2.60865 pd=16.14 as=6.1659 ps=32.4 w=15.81 l=2.54
X5 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=6.1659 pd=32.4 as=0 ps=0 w=15.81 l=2.54
X6 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=6.1659 pd=32.4 as=0 ps=0 w=15.81 l=2.54
X7 VDD1.t5 VP.t3 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.60865 pd=16.14 as=6.1659 ps=32.4 w=15.81 l=2.54
X8 VDD1.t3 VP.t4 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=6.1659 pd=32.4 as=2.60865 ps=16.14 w=15.81 l=2.54
X9 VTAIL.t1 VN.t2 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.60865 pd=16.14 as=2.60865 ps=16.14 w=15.81 l=2.54
X10 VDD1.t4 VP.t5 VTAIL.t4 B.t18 sky130_fd_pr__nfet_01v8 ad=6.1659 pd=32.4 as=2.60865 ps=16.14 w=15.81 l=2.54
X11 VDD2.t2 VN.t3 VTAIL.t10 B.t19 sky130_fd_pr__nfet_01v8 ad=2.60865 pd=16.14 as=6.1659 ps=32.4 w=15.81 l=2.54
X12 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.1659 pd=32.4 as=0 ps=0 w=15.81 l=2.54
X13 VDD2.t1 VN.t4 VTAIL.t11 B.t18 sky130_fd_pr__nfet_01v8 ad=6.1659 pd=32.4 as=2.60865 ps=16.14 w=15.81 l=2.54
X14 VDD2.t0 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.1659 pd=32.4 as=2.60865 ps=16.14 w=15.81 l=2.54
X15 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.1659 pd=32.4 as=0 ps=0 w=15.81 l=2.54
R0 VP.n11 VP.t4 182.352
R1 VP.n13 VP.n12 161.3
R2 VP.n14 VP.n9 161.3
R3 VP.n16 VP.n15 161.3
R4 VP.n17 VP.n8 161.3
R5 VP.n19 VP.n18 161.3
R6 VP.n20 VP.n7 161.3
R7 VP.n42 VP.n0 161.3
R8 VP.n41 VP.n40 161.3
R9 VP.n39 VP.n1 161.3
R10 VP.n38 VP.n37 161.3
R11 VP.n36 VP.n2 161.3
R12 VP.n35 VP.n34 161.3
R13 VP.n33 VP.n32 161.3
R14 VP.n31 VP.n4 161.3
R15 VP.n30 VP.n29 161.3
R16 VP.n28 VP.n5 161.3
R17 VP.n27 VP.n26 161.3
R18 VP.n25 VP.n6 161.3
R19 VP.n24 VP.t5 150.008
R20 VP.n3 VP.t1 150.008
R21 VP.n43 VP.t2 150.008
R22 VP.n21 VP.t3 150.008
R23 VP.n10 VP.t0 150.008
R24 VP.n24 VP.n23 104.885
R25 VP.n44 VP.n43 104.885
R26 VP.n22 VP.n21 104.885
R27 VP.n11 VP.n10 59.9599
R28 VP.n30 VP.n5 56.5193
R29 VP.n37 VP.n1 56.5193
R30 VP.n15 VP.n8 56.5193
R31 VP.n23 VP.n22 51.2685
R32 VP.n26 VP.n25 24.4675
R33 VP.n26 VP.n5 24.4675
R34 VP.n31 VP.n30 24.4675
R35 VP.n32 VP.n31 24.4675
R36 VP.n36 VP.n35 24.4675
R37 VP.n37 VP.n36 24.4675
R38 VP.n41 VP.n1 24.4675
R39 VP.n42 VP.n41 24.4675
R40 VP.n19 VP.n8 24.4675
R41 VP.n20 VP.n19 24.4675
R42 VP.n14 VP.n13 24.4675
R43 VP.n15 VP.n14 24.4675
R44 VP.n32 VP.n3 12.234
R45 VP.n35 VP.n3 12.234
R46 VP.n13 VP.n10 12.234
R47 VP.n12 VP.n11 7.1096
R48 VP.n25 VP.n24 5.87258
R49 VP.n43 VP.n42 5.87258
R50 VP.n21 VP.n20 5.87258
R51 VP.n22 VP.n7 0.278367
R52 VP.n23 VP.n6 0.278367
R53 VP.n44 VP.n0 0.278367
R54 VP.n12 VP.n9 0.189894
R55 VP.n16 VP.n9 0.189894
R56 VP.n17 VP.n16 0.189894
R57 VP.n18 VP.n17 0.189894
R58 VP.n18 VP.n7 0.189894
R59 VP.n27 VP.n6 0.189894
R60 VP.n28 VP.n27 0.189894
R61 VP.n29 VP.n28 0.189894
R62 VP.n29 VP.n4 0.189894
R63 VP.n33 VP.n4 0.189894
R64 VP.n34 VP.n33 0.189894
R65 VP.n34 VP.n2 0.189894
R66 VP.n38 VP.n2 0.189894
R67 VP.n39 VP.n38 0.189894
R68 VP.n40 VP.n39 0.189894
R69 VP.n40 VP.n0 0.189894
R70 VP VP.n44 0.153454
R71 VDD1 VDD1.t3 65.7199
R72 VDD1.n1 VDD1.t4 65.6062
R73 VDD1.n1 VDD1.n0 63.1167
R74 VDD1.n3 VDD1.n2 62.5536
R75 VDD1.n3 VDD1.n1 47.2056
R76 VDD1.n2 VDD1.t2 1.25287
R77 VDD1.n2 VDD1.t5 1.25287
R78 VDD1.n0 VDD1.t0 1.25287
R79 VDD1.n0 VDD1.t1 1.25287
R80 VDD1 VDD1.n3 0.560845
R81 VTAIL.n7 VTAIL.t10 47.1273
R82 VTAIL.n11 VTAIL.t3 47.1272
R83 VTAIL.n2 VTAIL.t7 47.1272
R84 VTAIL.n10 VTAIL.t6 47.1272
R85 VTAIL.n9 VTAIL.n8 45.875
R86 VTAIL.n6 VTAIL.n5 45.875
R87 VTAIL.n1 VTAIL.n0 45.8747
R88 VTAIL.n4 VTAIL.n3 45.8747
R89 VTAIL.n6 VTAIL.n4 30.9445
R90 VTAIL.n11 VTAIL.n10 28.4703
R91 VTAIL.n7 VTAIL.n6 2.47464
R92 VTAIL.n10 VTAIL.n9 2.47464
R93 VTAIL.n4 VTAIL.n2 2.47464
R94 VTAIL VTAIL.n11 1.79791
R95 VTAIL.n9 VTAIL.n7 1.7074
R96 VTAIL.n2 VTAIL.n1 1.7074
R97 VTAIL.n0 VTAIL.t0 1.25287
R98 VTAIL.n0 VTAIL.t1 1.25287
R99 VTAIL.n3 VTAIL.t4 1.25287
R100 VTAIL.n3 VTAIL.t8 1.25287
R101 VTAIL.n8 VTAIL.t5 1.25287
R102 VTAIL.n8 VTAIL.t9 1.25287
R103 VTAIL.n5 VTAIL.t11 1.25287
R104 VTAIL.n5 VTAIL.t2 1.25287
R105 VTAIL VTAIL.n1 0.677224
R106 B.n696 B.n141 585
R107 B.n141 B.n78 585
R108 B.n698 B.n697 585
R109 B.n700 B.n140 585
R110 B.n703 B.n702 585
R111 B.n704 B.n139 585
R112 B.n706 B.n705 585
R113 B.n708 B.n138 585
R114 B.n711 B.n710 585
R115 B.n712 B.n137 585
R116 B.n714 B.n713 585
R117 B.n716 B.n136 585
R118 B.n719 B.n718 585
R119 B.n720 B.n135 585
R120 B.n722 B.n721 585
R121 B.n724 B.n134 585
R122 B.n727 B.n726 585
R123 B.n728 B.n133 585
R124 B.n730 B.n729 585
R125 B.n732 B.n132 585
R126 B.n735 B.n734 585
R127 B.n736 B.n131 585
R128 B.n738 B.n737 585
R129 B.n740 B.n130 585
R130 B.n743 B.n742 585
R131 B.n744 B.n129 585
R132 B.n746 B.n745 585
R133 B.n748 B.n128 585
R134 B.n751 B.n750 585
R135 B.n752 B.n127 585
R136 B.n754 B.n753 585
R137 B.n756 B.n126 585
R138 B.n759 B.n758 585
R139 B.n760 B.n125 585
R140 B.n762 B.n761 585
R141 B.n764 B.n124 585
R142 B.n767 B.n766 585
R143 B.n768 B.n123 585
R144 B.n770 B.n769 585
R145 B.n772 B.n122 585
R146 B.n775 B.n774 585
R147 B.n776 B.n121 585
R148 B.n778 B.n777 585
R149 B.n780 B.n120 585
R150 B.n783 B.n782 585
R151 B.n784 B.n119 585
R152 B.n786 B.n785 585
R153 B.n788 B.n118 585
R154 B.n791 B.n790 585
R155 B.n792 B.n117 585
R156 B.n794 B.n793 585
R157 B.n796 B.n116 585
R158 B.n798 B.n797 585
R159 B.n800 B.n799 585
R160 B.n803 B.n802 585
R161 B.n804 B.n111 585
R162 B.n806 B.n805 585
R163 B.n808 B.n110 585
R164 B.n811 B.n810 585
R165 B.n812 B.n109 585
R166 B.n814 B.n813 585
R167 B.n816 B.n108 585
R168 B.n819 B.n818 585
R169 B.n821 B.n105 585
R170 B.n823 B.n822 585
R171 B.n825 B.n104 585
R172 B.n828 B.n827 585
R173 B.n829 B.n103 585
R174 B.n831 B.n830 585
R175 B.n833 B.n102 585
R176 B.n836 B.n835 585
R177 B.n837 B.n101 585
R178 B.n839 B.n838 585
R179 B.n841 B.n100 585
R180 B.n844 B.n843 585
R181 B.n845 B.n99 585
R182 B.n847 B.n846 585
R183 B.n849 B.n98 585
R184 B.n852 B.n851 585
R185 B.n853 B.n97 585
R186 B.n855 B.n854 585
R187 B.n857 B.n96 585
R188 B.n860 B.n859 585
R189 B.n861 B.n95 585
R190 B.n863 B.n862 585
R191 B.n865 B.n94 585
R192 B.n868 B.n867 585
R193 B.n869 B.n93 585
R194 B.n871 B.n870 585
R195 B.n873 B.n92 585
R196 B.n876 B.n875 585
R197 B.n877 B.n91 585
R198 B.n879 B.n878 585
R199 B.n881 B.n90 585
R200 B.n884 B.n883 585
R201 B.n885 B.n89 585
R202 B.n887 B.n886 585
R203 B.n889 B.n88 585
R204 B.n892 B.n891 585
R205 B.n893 B.n87 585
R206 B.n895 B.n894 585
R207 B.n897 B.n86 585
R208 B.n900 B.n899 585
R209 B.n901 B.n85 585
R210 B.n903 B.n902 585
R211 B.n905 B.n84 585
R212 B.n908 B.n907 585
R213 B.n909 B.n83 585
R214 B.n911 B.n910 585
R215 B.n913 B.n82 585
R216 B.n916 B.n915 585
R217 B.n917 B.n81 585
R218 B.n919 B.n918 585
R219 B.n921 B.n80 585
R220 B.n924 B.n923 585
R221 B.n925 B.n79 585
R222 B.n695 B.n77 585
R223 B.n928 B.n77 585
R224 B.n694 B.n76 585
R225 B.n929 B.n76 585
R226 B.n693 B.n75 585
R227 B.n930 B.n75 585
R228 B.n692 B.n691 585
R229 B.n691 B.n71 585
R230 B.n690 B.n70 585
R231 B.n936 B.n70 585
R232 B.n689 B.n69 585
R233 B.n937 B.n69 585
R234 B.n688 B.n68 585
R235 B.n938 B.n68 585
R236 B.n687 B.n686 585
R237 B.n686 B.n67 585
R238 B.n685 B.n63 585
R239 B.n944 B.n63 585
R240 B.n684 B.n62 585
R241 B.n945 B.n62 585
R242 B.n683 B.n61 585
R243 B.n946 B.n61 585
R244 B.n682 B.n681 585
R245 B.n681 B.n57 585
R246 B.n680 B.n56 585
R247 B.n952 B.n56 585
R248 B.n679 B.n55 585
R249 B.n953 B.n55 585
R250 B.n678 B.n54 585
R251 B.n954 B.n54 585
R252 B.n677 B.n676 585
R253 B.n676 B.n50 585
R254 B.n675 B.n49 585
R255 B.n960 B.n49 585
R256 B.n674 B.n48 585
R257 B.n961 B.n48 585
R258 B.n673 B.n47 585
R259 B.n962 B.n47 585
R260 B.n672 B.n671 585
R261 B.n671 B.n46 585
R262 B.n670 B.n42 585
R263 B.n968 B.n42 585
R264 B.n669 B.n41 585
R265 B.n969 B.n41 585
R266 B.n668 B.n40 585
R267 B.n970 B.n40 585
R268 B.n667 B.n666 585
R269 B.n666 B.n36 585
R270 B.n665 B.n35 585
R271 B.n976 B.n35 585
R272 B.n664 B.n34 585
R273 B.n977 B.n34 585
R274 B.n663 B.n33 585
R275 B.n978 B.n33 585
R276 B.n662 B.n661 585
R277 B.n661 B.n32 585
R278 B.n660 B.n28 585
R279 B.n984 B.n28 585
R280 B.n659 B.n27 585
R281 B.n985 B.n27 585
R282 B.n658 B.n26 585
R283 B.n986 B.n26 585
R284 B.n657 B.n656 585
R285 B.n656 B.n22 585
R286 B.n655 B.n21 585
R287 B.n992 B.n21 585
R288 B.n654 B.n20 585
R289 B.n993 B.n20 585
R290 B.n653 B.n19 585
R291 B.n994 B.n19 585
R292 B.n652 B.n651 585
R293 B.n651 B.n15 585
R294 B.n650 B.n14 585
R295 B.n1000 B.n14 585
R296 B.n649 B.n13 585
R297 B.n1001 B.n13 585
R298 B.n648 B.n12 585
R299 B.n1002 B.n12 585
R300 B.n647 B.n646 585
R301 B.n646 B.n8 585
R302 B.n645 B.n7 585
R303 B.n1008 B.n7 585
R304 B.n644 B.n6 585
R305 B.n1009 B.n6 585
R306 B.n643 B.n5 585
R307 B.n1010 B.n5 585
R308 B.n642 B.n641 585
R309 B.n641 B.n4 585
R310 B.n640 B.n142 585
R311 B.n640 B.n639 585
R312 B.n630 B.n143 585
R313 B.n144 B.n143 585
R314 B.n632 B.n631 585
R315 B.n633 B.n632 585
R316 B.n629 B.n149 585
R317 B.n149 B.n148 585
R318 B.n628 B.n627 585
R319 B.n627 B.n626 585
R320 B.n151 B.n150 585
R321 B.n152 B.n151 585
R322 B.n619 B.n618 585
R323 B.n620 B.n619 585
R324 B.n617 B.n157 585
R325 B.n157 B.n156 585
R326 B.n616 B.n615 585
R327 B.n615 B.n614 585
R328 B.n159 B.n158 585
R329 B.n160 B.n159 585
R330 B.n607 B.n606 585
R331 B.n608 B.n607 585
R332 B.n605 B.n165 585
R333 B.n165 B.n164 585
R334 B.n604 B.n603 585
R335 B.n603 B.n602 585
R336 B.n167 B.n166 585
R337 B.n595 B.n167 585
R338 B.n594 B.n593 585
R339 B.n596 B.n594 585
R340 B.n592 B.n172 585
R341 B.n172 B.n171 585
R342 B.n591 B.n590 585
R343 B.n590 B.n589 585
R344 B.n174 B.n173 585
R345 B.n175 B.n174 585
R346 B.n582 B.n581 585
R347 B.n583 B.n582 585
R348 B.n580 B.n180 585
R349 B.n180 B.n179 585
R350 B.n579 B.n578 585
R351 B.n578 B.n577 585
R352 B.n182 B.n181 585
R353 B.n570 B.n182 585
R354 B.n569 B.n568 585
R355 B.n571 B.n569 585
R356 B.n567 B.n187 585
R357 B.n187 B.n186 585
R358 B.n566 B.n565 585
R359 B.n565 B.n564 585
R360 B.n189 B.n188 585
R361 B.n190 B.n189 585
R362 B.n557 B.n556 585
R363 B.n558 B.n557 585
R364 B.n555 B.n195 585
R365 B.n195 B.n194 585
R366 B.n554 B.n553 585
R367 B.n553 B.n552 585
R368 B.n197 B.n196 585
R369 B.n198 B.n197 585
R370 B.n545 B.n544 585
R371 B.n546 B.n545 585
R372 B.n543 B.n203 585
R373 B.n203 B.n202 585
R374 B.n542 B.n541 585
R375 B.n541 B.n540 585
R376 B.n205 B.n204 585
R377 B.n533 B.n205 585
R378 B.n532 B.n531 585
R379 B.n534 B.n532 585
R380 B.n530 B.n210 585
R381 B.n210 B.n209 585
R382 B.n529 B.n528 585
R383 B.n528 B.n527 585
R384 B.n212 B.n211 585
R385 B.n213 B.n212 585
R386 B.n520 B.n519 585
R387 B.n521 B.n520 585
R388 B.n518 B.n218 585
R389 B.n218 B.n217 585
R390 B.n517 B.n516 585
R391 B.n516 B.n515 585
R392 B.n512 B.n222 585
R393 B.n511 B.n510 585
R394 B.n508 B.n223 585
R395 B.n508 B.n221 585
R396 B.n507 B.n506 585
R397 B.n505 B.n504 585
R398 B.n503 B.n225 585
R399 B.n501 B.n500 585
R400 B.n499 B.n226 585
R401 B.n498 B.n497 585
R402 B.n495 B.n227 585
R403 B.n493 B.n492 585
R404 B.n491 B.n228 585
R405 B.n490 B.n489 585
R406 B.n487 B.n229 585
R407 B.n485 B.n484 585
R408 B.n483 B.n230 585
R409 B.n482 B.n481 585
R410 B.n479 B.n231 585
R411 B.n477 B.n476 585
R412 B.n475 B.n232 585
R413 B.n474 B.n473 585
R414 B.n471 B.n233 585
R415 B.n469 B.n468 585
R416 B.n467 B.n234 585
R417 B.n466 B.n465 585
R418 B.n463 B.n235 585
R419 B.n461 B.n460 585
R420 B.n459 B.n236 585
R421 B.n458 B.n457 585
R422 B.n455 B.n237 585
R423 B.n453 B.n452 585
R424 B.n451 B.n238 585
R425 B.n450 B.n449 585
R426 B.n447 B.n239 585
R427 B.n445 B.n444 585
R428 B.n443 B.n240 585
R429 B.n442 B.n441 585
R430 B.n439 B.n241 585
R431 B.n437 B.n436 585
R432 B.n435 B.n242 585
R433 B.n434 B.n433 585
R434 B.n431 B.n243 585
R435 B.n429 B.n428 585
R436 B.n427 B.n244 585
R437 B.n426 B.n425 585
R438 B.n423 B.n245 585
R439 B.n421 B.n420 585
R440 B.n419 B.n246 585
R441 B.n418 B.n417 585
R442 B.n415 B.n247 585
R443 B.n413 B.n412 585
R444 B.n411 B.n248 585
R445 B.n410 B.n409 585
R446 B.n407 B.n406 585
R447 B.n405 B.n404 585
R448 B.n403 B.n253 585
R449 B.n401 B.n400 585
R450 B.n399 B.n254 585
R451 B.n398 B.n397 585
R452 B.n395 B.n255 585
R453 B.n393 B.n392 585
R454 B.n391 B.n256 585
R455 B.n389 B.n388 585
R456 B.n386 B.n259 585
R457 B.n384 B.n383 585
R458 B.n382 B.n260 585
R459 B.n381 B.n380 585
R460 B.n378 B.n261 585
R461 B.n376 B.n375 585
R462 B.n374 B.n262 585
R463 B.n373 B.n372 585
R464 B.n370 B.n263 585
R465 B.n368 B.n367 585
R466 B.n366 B.n264 585
R467 B.n365 B.n364 585
R468 B.n362 B.n265 585
R469 B.n360 B.n359 585
R470 B.n358 B.n266 585
R471 B.n357 B.n356 585
R472 B.n354 B.n267 585
R473 B.n352 B.n351 585
R474 B.n350 B.n268 585
R475 B.n349 B.n348 585
R476 B.n346 B.n269 585
R477 B.n344 B.n343 585
R478 B.n342 B.n270 585
R479 B.n341 B.n340 585
R480 B.n338 B.n271 585
R481 B.n336 B.n335 585
R482 B.n334 B.n272 585
R483 B.n333 B.n332 585
R484 B.n330 B.n273 585
R485 B.n328 B.n327 585
R486 B.n326 B.n274 585
R487 B.n325 B.n324 585
R488 B.n322 B.n275 585
R489 B.n320 B.n319 585
R490 B.n318 B.n276 585
R491 B.n317 B.n316 585
R492 B.n314 B.n277 585
R493 B.n312 B.n311 585
R494 B.n310 B.n278 585
R495 B.n309 B.n308 585
R496 B.n306 B.n279 585
R497 B.n304 B.n303 585
R498 B.n302 B.n280 585
R499 B.n301 B.n300 585
R500 B.n298 B.n281 585
R501 B.n296 B.n295 585
R502 B.n294 B.n282 585
R503 B.n293 B.n292 585
R504 B.n290 B.n283 585
R505 B.n288 B.n287 585
R506 B.n286 B.n285 585
R507 B.n220 B.n219 585
R508 B.n514 B.n513 585
R509 B.n515 B.n514 585
R510 B.n216 B.n215 585
R511 B.n217 B.n216 585
R512 B.n523 B.n522 585
R513 B.n522 B.n521 585
R514 B.n524 B.n214 585
R515 B.n214 B.n213 585
R516 B.n526 B.n525 585
R517 B.n527 B.n526 585
R518 B.n208 B.n207 585
R519 B.n209 B.n208 585
R520 B.n536 B.n535 585
R521 B.n535 B.n534 585
R522 B.n537 B.n206 585
R523 B.n533 B.n206 585
R524 B.n539 B.n538 585
R525 B.n540 B.n539 585
R526 B.n201 B.n200 585
R527 B.n202 B.n201 585
R528 B.n548 B.n547 585
R529 B.n547 B.n546 585
R530 B.n549 B.n199 585
R531 B.n199 B.n198 585
R532 B.n551 B.n550 585
R533 B.n552 B.n551 585
R534 B.n193 B.n192 585
R535 B.n194 B.n193 585
R536 B.n560 B.n559 585
R537 B.n559 B.n558 585
R538 B.n561 B.n191 585
R539 B.n191 B.n190 585
R540 B.n563 B.n562 585
R541 B.n564 B.n563 585
R542 B.n185 B.n184 585
R543 B.n186 B.n185 585
R544 B.n573 B.n572 585
R545 B.n572 B.n571 585
R546 B.n574 B.n183 585
R547 B.n570 B.n183 585
R548 B.n576 B.n575 585
R549 B.n577 B.n576 585
R550 B.n178 B.n177 585
R551 B.n179 B.n178 585
R552 B.n585 B.n584 585
R553 B.n584 B.n583 585
R554 B.n586 B.n176 585
R555 B.n176 B.n175 585
R556 B.n588 B.n587 585
R557 B.n589 B.n588 585
R558 B.n170 B.n169 585
R559 B.n171 B.n170 585
R560 B.n598 B.n597 585
R561 B.n597 B.n596 585
R562 B.n599 B.n168 585
R563 B.n595 B.n168 585
R564 B.n601 B.n600 585
R565 B.n602 B.n601 585
R566 B.n163 B.n162 585
R567 B.n164 B.n163 585
R568 B.n610 B.n609 585
R569 B.n609 B.n608 585
R570 B.n611 B.n161 585
R571 B.n161 B.n160 585
R572 B.n613 B.n612 585
R573 B.n614 B.n613 585
R574 B.n155 B.n154 585
R575 B.n156 B.n155 585
R576 B.n622 B.n621 585
R577 B.n621 B.n620 585
R578 B.n623 B.n153 585
R579 B.n153 B.n152 585
R580 B.n625 B.n624 585
R581 B.n626 B.n625 585
R582 B.n147 B.n146 585
R583 B.n148 B.n147 585
R584 B.n635 B.n634 585
R585 B.n634 B.n633 585
R586 B.n636 B.n145 585
R587 B.n145 B.n144 585
R588 B.n638 B.n637 585
R589 B.n639 B.n638 585
R590 B.n2 B.n0 585
R591 B.n4 B.n2 585
R592 B.n3 B.n1 585
R593 B.n1009 B.n3 585
R594 B.n1007 B.n1006 585
R595 B.n1008 B.n1007 585
R596 B.n1005 B.n9 585
R597 B.n9 B.n8 585
R598 B.n1004 B.n1003 585
R599 B.n1003 B.n1002 585
R600 B.n11 B.n10 585
R601 B.n1001 B.n11 585
R602 B.n999 B.n998 585
R603 B.n1000 B.n999 585
R604 B.n997 B.n16 585
R605 B.n16 B.n15 585
R606 B.n996 B.n995 585
R607 B.n995 B.n994 585
R608 B.n18 B.n17 585
R609 B.n993 B.n18 585
R610 B.n991 B.n990 585
R611 B.n992 B.n991 585
R612 B.n989 B.n23 585
R613 B.n23 B.n22 585
R614 B.n988 B.n987 585
R615 B.n987 B.n986 585
R616 B.n25 B.n24 585
R617 B.n985 B.n25 585
R618 B.n983 B.n982 585
R619 B.n984 B.n983 585
R620 B.n981 B.n29 585
R621 B.n32 B.n29 585
R622 B.n980 B.n979 585
R623 B.n979 B.n978 585
R624 B.n31 B.n30 585
R625 B.n977 B.n31 585
R626 B.n975 B.n974 585
R627 B.n976 B.n975 585
R628 B.n973 B.n37 585
R629 B.n37 B.n36 585
R630 B.n972 B.n971 585
R631 B.n971 B.n970 585
R632 B.n39 B.n38 585
R633 B.n969 B.n39 585
R634 B.n967 B.n966 585
R635 B.n968 B.n967 585
R636 B.n965 B.n43 585
R637 B.n46 B.n43 585
R638 B.n964 B.n963 585
R639 B.n963 B.n962 585
R640 B.n45 B.n44 585
R641 B.n961 B.n45 585
R642 B.n959 B.n958 585
R643 B.n960 B.n959 585
R644 B.n957 B.n51 585
R645 B.n51 B.n50 585
R646 B.n956 B.n955 585
R647 B.n955 B.n954 585
R648 B.n53 B.n52 585
R649 B.n953 B.n53 585
R650 B.n951 B.n950 585
R651 B.n952 B.n951 585
R652 B.n949 B.n58 585
R653 B.n58 B.n57 585
R654 B.n948 B.n947 585
R655 B.n947 B.n946 585
R656 B.n60 B.n59 585
R657 B.n945 B.n60 585
R658 B.n943 B.n942 585
R659 B.n944 B.n943 585
R660 B.n941 B.n64 585
R661 B.n67 B.n64 585
R662 B.n940 B.n939 585
R663 B.n939 B.n938 585
R664 B.n66 B.n65 585
R665 B.n937 B.n66 585
R666 B.n935 B.n934 585
R667 B.n936 B.n935 585
R668 B.n933 B.n72 585
R669 B.n72 B.n71 585
R670 B.n932 B.n931 585
R671 B.n931 B.n930 585
R672 B.n74 B.n73 585
R673 B.n929 B.n74 585
R674 B.n927 B.n926 585
R675 B.n928 B.n927 585
R676 B.n1012 B.n1011 585
R677 B.n1011 B.n1010 585
R678 B.n514 B.n222 497.305
R679 B.n927 B.n79 497.305
R680 B.n516 B.n220 497.305
R681 B.n141 B.n77 497.305
R682 B.n257 B.t15 358.625
R683 B.n112 B.t4 358.625
R684 B.n249 B.t8 358.291
R685 B.n106 B.t12 358.291
R686 B.n699 B.n78 256.663
R687 B.n701 B.n78 256.663
R688 B.n707 B.n78 256.663
R689 B.n709 B.n78 256.663
R690 B.n715 B.n78 256.663
R691 B.n717 B.n78 256.663
R692 B.n723 B.n78 256.663
R693 B.n725 B.n78 256.663
R694 B.n731 B.n78 256.663
R695 B.n733 B.n78 256.663
R696 B.n739 B.n78 256.663
R697 B.n741 B.n78 256.663
R698 B.n747 B.n78 256.663
R699 B.n749 B.n78 256.663
R700 B.n755 B.n78 256.663
R701 B.n757 B.n78 256.663
R702 B.n763 B.n78 256.663
R703 B.n765 B.n78 256.663
R704 B.n771 B.n78 256.663
R705 B.n773 B.n78 256.663
R706 B.n779 B.n78 256.663
R707 B.n781 B.n78 256.663
R708 B.n787 B.n78 256.663
R709 B.n789 B.n78 256.663
R710 B.n795 B.n78 256.663
R711 B.n115 B.n78 256.663
R712 B.n801 B.n78 256.663
R713 B.n807 B.n78 256.663
R714 B.n809 B.n78 256.663
R715 B.n815 B.n78 256.663
R716 B.n817 B.n78 256.663
R717 B.n824 B.n78 256.663
R718 B.n826 B.n78 256.663
R719 B.n832 B.n78 256.663
R720 B.n834 B.n78 256.663
R721 B.n840 B.n78 256.663
R722 B.n842 B.n78 256.663
R723 B.n848 B.n78 256.663
R724 B.n850 B.n78 256.663
R725 B.n856 B.n78 256.663
R726 B.n858 B.n78 256.663
R727 B.n864 B.n78 256.663
R728 B.n866 B.n78 256.663
R729 B.n872 B.n78 256.663
R730 B.n874 B.n78 256.663
R731 B.n880 B.n78 256.663
R732 B.n882 B.n78 256.663
R733 B.n888 B.n78 256.663
R734 B.n890 B.n78 256.663
R735 B.n896 B.n78 256.663
R736 B.n898 B.n78 256.663
R737 B.n904 B.n78 256.663
R738 B.n906 B.n78 256.663
R739 B.n912 B.n78 256.663
R740 B.n914 B.n78 256.663
R741 B.n920 B.n78 256.663
R742 B.n922 B.n78 256.663
R743 B.n509 B.n221 256.663
R744 B.n224 B.n221 256.663
R745 B.n502 B.n221 256.663
R746 B.n496 B.n221 256.663
R747 B.n494 B.n221 256.663
R748 B.n488 B.n221 256.663
R749 B.n486 B.n221 256.663
R750 B.n480 B.n221 256.663
R751 B.n478 B.n221 256.663
R752 B.n472 B.n221 256.663
R753 B.n470 B.n221 256.663
R754 B.n464 B.n221 256.663
R755 B.n462 B.n221 256.663
R756 B.n456 B.n221 256.663
R757 B.n454 B.n221 256.663
R758 B.n448 B.n221 256.663
R759 B.n446 B.n221 256.663
R760 B.n440 B.n221 256.663
R761 B.n438 B.n221 256.663
R762 B.n432 B.n221 256.663
R763 B.n430 B.n221 256.663
R764 B.n424 B.n221 256.663
R765 B.n422 B.n221 256.663
R766 B.n416 B.n221 256.663
R767 B.n414 B.n221 256.663
R768 B.n408 B.n221 256.663
R769 B.n252 B.n221 256.663
R770 B.n402 B.n221 256.663
R771 B.n396 B.n221 256.663
R772 B.n394 B.n221 256.663
R773 B.n387 B.n221 256.663
R774 B.n385 B.n221 256.663
R775 B.n379 B.n221 256.663
R776 B.n377 B.n221 256.663
R777 B.n371 B.n221 256.663
R778 B.n369 B.n221 256.663
R779 B.n363 B.n221 256.663
R780 B.n361 B.n221 256.663
R781 B.n355 B.n221 256.663
R782 B.n353 B.n221 256.663
R783 B.n347 B.n221 256.663
R784 B.n345 B.n221 256.663
R785 B.n339 B.n221 256.663
R786 B.n337 B.n221 256.663
R787 B.n331 B.n221 256.663
R788 B.n329 B.n221 256.663
R789 B.n323 B.n221 256.663
R790 B.n321 B.n221 256.663
R791 B.n315 B.n221 256.663
R792 B.n313 B.n221 256.663
R793 B.n307 B.n221 256.663
R794 B.n305 B.n221 256.663
R795 B.n299 B.n221 256.663
R796 B.n297 B.n221 256.663
R797 B.n291 B.n221 256.663
R798 B.n289 B.n221 256.663
R799 B.n284 B.n221 256.663
R800 B.n514 B.n216 163.367
R801 B.n522 B.n216 163.367
R802 B.n522 B.n214 163.367
R803 B.n526 B.n214 163.367
R804 B.n526 B.n208 163.367
R805 B.n535 B.n208 163.367
R806 B.n535 B.n206 163.367
R807 B.n539 B.n206 163.367
R808 B.n539 B.n201 163.367
R809 B.n547 B.n201 163.367
R810 B.n547 B.n199 163.367
R811 B.n551 B.n199 163.367
R812 B.n551 B.n193 163.367
R813 B.n559 B.n193 163.367
R814 B.n559 B.n191 163.367
R815 B.n563 B.n191 163.367
R816 B.n563 B.n185 163.367
R817 B.n572 B.n185 163.367
R818 B.n572 B.n183 163.367
R819 B.n576 B.n183 163.367
R820 B.n576 B.n178 163.367
R821 B.n584 B.n178 163.367
R822 B.n584 B.n176 163.367
R823 B.n588 B.n176 163.367
R824 B.n588 B.n170 163.367
R825 B.n597 B.n170 163.367
R826 B.n597 B.n168 163.367
R827 B.n601 B.n168 163.367
R828 B.n601 B.n163 163.367
R829 B.n609 B.n163 163.367
R830 B.n609 B.n161 163.367
R831 B.n613 B.n161 163.367
R832 B.n613 B.n155 163.367
R833 B.n621 B.n155 163.367
R834 B.n621 B.n153 163.367
R835 B.n625 B.n153 163.367
R836 B.n625 B.n147 163.367
R837 B.n634 B.n147 163.367
R838 B.n634 B.n145 163.367
R839 B.n638 B.n145 163.367
R840 B.n638 B.n2 163.367
R841 B.n1011 B.n2 163.367
R842 B.n1011 B.n3 163.367
R843 B.n1007 B.n3 163.367
R844 B.n1007 B.n9 163.367
R845 B.n1003 B.n9 163.367
R846 B.n1003 B.n11 163.367
R847 B.n999 B.n11 163.367
R848 B.n999 B.n16 163.367
R849 B.n995 B.n16 163.367
R850 B.n995 B.n18 163.367
R851 B.n991 B.n18 163.367
R852 B.n991 B.n23 163.367
R853 B.n987 B.n23 163.367
R854 B.n987 B.n25 163.367
R855 B.n983 B.n25 163.367
R856 B.n983 B.n29 163.367
R857 B.n979 B.n29 163.367
R858 B.n979 B.n31 163.367
R859 B.n975 B.n31 163.367
R860 B.n975 B.n37 163.367
R861 B.n971 B.n37 163.367
R862 B.n971 B.n39 163.367
R863 B.n967 B.n39 163.367
R864 B.n967 B.n43 163.367
R865 B.n963 B.n43 163.367
R866 B.n963 B.n45 163.367
R867 B.n959 B.n45 163.367
R868 B.n959 B.n51 163.367
R869 B.n955 B.n51 163.367
R870 B.n955 B.n53 163.367
R871 B.n951 B.n53 163.367
R872 B.n951 B.n58 163.367
R873 B.n947 B.n58 163.367
R874 B.n947 B.n60 163.367
R875 B.n943 B.n60 163.367
R876 B.n943 B.n64 163.367
R877 B.n939 B.n64 163.367
R878 B.n939 B.n66 163.367
R879 B.n935 B.n66 163.367
R880 B.n935 B.n72 163.367
R881 B.n931 B.n72 163.367
R882 B.n931 B.n74 163.367
R883 B.n927 B.n74 163.367
R884 B.n510 B.n508 163.367
R885 B.n508 B.n507 163.367
R886 B.n504 B.n503 163.367
R887 B.n501 B.n226 163.367
R888 B.n497 B.n495 163.367
R889 B.n493 B.n228 163.367
R890 B.n489 B.n487 163.367
R891 B.n485 B.n230 163.367
R892 B.n481 B.n479 163.367
R893 B.n477 B.n232 163.367
R894 B.n473 B.n471 163.367
R895 B.n469 B.n234 163.367
R896 B.n465 B.n463 163.367
R897 B.n461 B.n236 163.367
R898 B.n457 B.n455 163.367
R899 B.n453 B.n238 163.367
R900 B.n449 B.n447 163.367
R901 B.n445 B.n240 163.367
R902 B.n441 B.n439 163.367
R903 B.n437 B.n242 163.367
R904 B.n433 B.n431 163.367
R905 B.n429 B.n244 163.367
R906 B.n425 B.n423 163.367
R907 B.n421 B.n246 163.367
R908 B.n417 B.n415 163.367
R909 B.n413 B.n248 163.367
R910 B.n409 B.n407 163.367
R911 B.n404 B.n403 163.367
R912 B.n401 B.n254 163.367
R913 B.n397 B.n395 163.367
R914 B.n393 B.n256 163.367
R915 B.n388 B.n386 163.367
R916 B.n384 B.n260 163.367
R917 B.n380 B.n378 163.367
R918 B.n376 B.n262 163.367
R919 B.n372 B.n370 163.367
R920 B.n368 B.n264 163.367
R921 B.n364 B.n362 163.367
R922 B.n360 B.n266 163.367
R923 B.n356 B.n354 163.367
R924 B.n352 B.n268 163.367
R925 B.n348 B.n346 163.367
R926 B.n344 B.n270 163.367
R927 B.n340 B.n338 163.367
R928 B.n336 B.n272 163.367
R929 B.n332 B.n330 163.367
R930 B.n328 B.n274 163.367
R931 B.n324 B.n322 163.367
R932 B.n320 B.n276 163.367
R933 B.n316 B.n314 163.367
R934 B.n312 B.n278 163.367
R935 B.n308 B.n306 163.367
R936 B.n304 B.n280 163.367
R937 B.n300 B.n298 163.367
R938 B.n296 B.n282 163.367
R939 B.n292 B.n290 163.367
R940 B.n288 B.n285 163.367
R941 B.n516 B.n218 163.367
R942 B.n520 B.n218 163.367
R943 B.n520 B.n212 163.367
R944 B.n528 B.n212 163.367
R945 B.n528 B.n210 163.367
R946 B.n532 B.n210 163.367
R947 B.n532 B.n205 163.367
R948 B.n541 B.n205 163.367
R949 B.n541 B.n203 163.367
R950 B.n545 B.n203 163.367
R951 B.n545 B.n197 163.367
R952 B.n553 B.n197 163.367
R953 B.n553 B.n195 163.367
R954 B.n557 B.n195 163.367
R955 B.n557 B.n189 163.367
R956 B.n565 B.n189 163.367
R957 B.n565 B.n187 163.367
R958 B.n569 B.n187 163.367
R959 B.n569 B.n182 163.367
R960 B.n578 B.n182 163.367
R961 B.n578 B.n180 163.367
R962 B.n582 B.n180 163.367
R963 B.n582 B.n174 163.367
R964 B.n590 B.n174 163.367
R965 B.n590 B.n172 163.367
R966 B.n594 B.n172 163.367
R967 B.n594 B.n167 163.367
R968 B.n603 B.n167 163.367
R969 B.n603 B.n165 163.367
R970 B.n607 B.n165 163.367
R971 B.n607 B.n159 163.367
R972 B.n615 B.n159 163.367
R973 B.n615 B.n157 163.367
R974 B.n619 B.n157 163.367
R975 B.n619 B.n151 163.367
R976 B.n627 B.n151 163.367
R977 B.n627 B.n149 163.367
R978 B.n632 B.n149 163.367
R979 B.n632 B.n143 163.367
R980 B.n640 B.n143 163.367
R981 B.n641 B.n640 163.367
R982 B.n641 B.n5 163.367
R983 B.n6 B.n5 163.367
R984 B.n7 B.n6 163.367
R985 B.n646 B.n7 163.367
R986 B.n646 B.n12 163.367
R987 B.n13 B.n12 163.367
R988 B.n14 B.n13 163.367
R989 B.n651 B.n14 163.367
R990 B.n651 B.n19 163.367
R991 B.n20 B.n19 163.367
R992 B.n21 B.n20 163.367
R993 B.n656 B.n21 163.367
R994 B.n656 B.n26 163.367
R995 B.n27 B.n26 163.367
R996 B.n28 B.n27 163.367
R997 B.n661 B.n28 163.367
R998 B.n661 B.n33 163.367
R999 B.n34 B.n33 163.367
R1000 B.n35 B.n34 163.367
R1001 B.n666 B.n35 163.367
R1002 B.n666 B.n40 163.367
R1003 B.n41 B.n40 163.367
R1004 B.n42 B.n41 163.367
R1005 B.n671 B.n42 163.367
R1006 B.n671 B.n47 163.367
R1007 B.n48 B.n47 163.367
R1008 B.n49 B.n48 163.367
R1009 B.n676 B.n49 163.367
R1010 B.n676 B.n54 163.367
R1011 B.n55 B.n54 163.367
R1012 B.n56 B.n55 163.367
R1013 B.n681 B.n56 163.367
R1014 B.n681 B.n61 163.367
R1015 B.n62 B.n61 163.367
R1016 B.n63 B.n62 163.367
R1017 B.n686 B.n63 163.367
R1018 B.n686 B.n68 163.367
R1019 B.n69 B.n68 163.367
R1020 B.n70 B.n69 163.367
R1021 B.n691 B.n70 163.367
R1022 B.n691 B.n75 163.367
R1023 B.n76 B.n75 163.367
R1024 B.n77 B.n76 163.367
R1025 B.n923 B.n921 163.367
R1026 B.n919 B.n81 163.367
R1027 B.n915 B.n913 163.367
R1028 B.n911 B.n83 163.367
R1029 B.n907 B.n905 163.367
R1030 B.n903 B.n85 163.367
R1031 B.n899 B.n897 163.367
R1032 B.n895 B.n87 163.367
R1033 B.n891 B.n889 163.367
R1034 B.n887 B.n89 163.367
R1035 B.n883 B.n881 163.367
R1036 B.n879 B.n91 163.367
R1037 B.n875 B.n873 163.367
R1038 B.n871 B.n93 163.367
R1039 B.n867 B.n865 163.367
R1040 B.n863 B.n95 163.367
R1041 B.n859 B.n857 163.367
R1042 B.n855 B.n97 163.367
R1043 B.n851 B.n849 163.367
R1044 B.n847 B.n99 163.367
R1045 B.n843 B.n841 163.367
R1046 B.n839 B.n101 163.367
R1047 B.n835 B.n833 163.367
R1048 B.n831 B.n103 163.367
R1049 B.n827 B.n825 163.367
R1050 B.n823 B.n105 163.367
R1051 B.n818 B.n816 163.367
R1052 B.n814 B.n109 163.367
R1053 B.n810 B.n808 163.367
R1054 B.n806 B.n111 163.367
R1055 B.n802 B.n800 163.367
R1056 B.n797 B.n796 163.367
R1057 B.n794 B.n117 163.367
R1058 B.n790 B.n788 163.367
R1059 B.n786 B.n119 163.367
R1060 B.n782 B.n780 163.367
R1061 B.n778 B.n121 163.367
R1062 B.n774 B.n772 163.367
R1063 B.n770 B.n123 163.367
R1064 B.n766 B.n764 163.367
R1065 B.n762 B.n125 163.367
R1066 B.n758 B.n756 163.367
R1067 B.n754 B.n127 163.367
R1068 B.n750 B.n748 163.367
R1069 B.n746 B.n129 163.367
R1070 B.n742 B.n740 163.367
R1071 B.n738 B.n131 163.367
R1072 B.n734 B.n732 163.367
R1073 B.n730 B.n133 163.367
R1074 B.n726 B.n724 163.367
R1075 B.n722 B.n135 163.367
R1076 B.n718 B.n716 163.367
R1077 B.n714 B.n137 163.367
R1078 B.n710 B.n708 163.367
R1079 B.n706 B.n139 163.367
R1080 B.n702 B.n700 163.367
R1081 B.n698 B.n141 163.367
R1082 B.n257 B.t17 126.549
R1083 B.n112 B.t6 126.549
R1084 B.n249 B.t11 126.528
R1085 B.n106 B.t13 126.528
R1086 B.n509 B.n222 71.676
R1087 B.n507 B.n224 71.676
R1088 B.n503 B.n502 71.676
R1089 B.n496 B.n226 71.676
R1090 B.n495 B.n494 71.676
R1091 B.n488 B.n228 71.676
R1092 B.n487 B.n486 71.676
R1093 B.n480 B.n230 71.676
R1094 B.n479 B.n478 71.676
R1095 B.n472 B.n232 71.676
R1096 B.n471 B.n470 71.676
R1097 B.n464 B.n234 71.676
R1098 B.n463 B.n462 71.676
R1099 B.n456 B.n236 71.676
R1100 B.n455 B.n454 71.676
R1101 B.n448 B.n238 71.676
R1102 B.n447 B.n446 71.676
R1103 B.n440 B.n240 71.676
R1104 B.n439 B.n438 71.676
R1105 B.n432 B.n242 71.676
R1106 B.n431 B.n430 71.676
R1107 B.n424 B.n244 71.676
R1108 B.n423 B.n422 71.676
R1109 B.n416 B.n246 71.676
R1110 B.n415 B.n414 71.676
R1111 B.n408 B.n248 71.676
R1112 B.n407 B.n252 71.676
R1113 B.n403 B.n402 71.676
R1114 B.n396 B.n254 71.676
R1115 B.n395 B.n394 71.676
R1116 B.n387 B.n256 71.676
R1117 B.n386 B.n385 71.676
R1118 B.n379 B.n260 71.676
R1119 B.n378 B.n377 71.676
R1120 B.n371 B.n262 71.676
R1121 B.n370 B.n369 71.676
R1122 B.n363 B.n264 71.676
R1123 B.n362 B.n361 71.676
R1124 B.n355 B.n266 71.676
R1125 B.n354 B.n353 71.676
R1126 B.n347 B.n268 71.676
R1127 B.n346 B.n345 71.676
R1128 B.n339 B.n270 71.676
R1129 B.n338 B.n337 71.676
R1130 B.n331 B.n272 71.676
R1131 B.n330 B.n329 71.676
R1132 B.n323 B.n274 71.676
R1133 B.n322 B.n321 71.676
R1134 B.n315 B.n276 71.676
R1135 B.n314 B.n313 71.676
R1136 B.n307 B.n278 71.676
R1137 B.n306 B.n305 71.676
R1138 B.n299 B.n280 71.676
R1139 B.n298 B.n297 71.676
R1140 B.n291 B.n282 71.676
R1141 B.n290 B.n289 71.676
R1142 B.n285 B.n284 71.676
R1143 B.n922 B.n79 71.676
R1144 B.n921 B.n920 71.676
R1145 B.n914 B.n81 71.676
R1146 B.n913 B.n912 71.676
R1147 B.n906 B.n83 71.676
R1148 B.n905 B.n904 71.676
R1149 B.n898 B.n85 71.676
R1150 B.n897 B.n896 71.676
R1151 B.n890 B.n87 71.676
R1152 B.n889 B.n888 71.676
R1153 B.n882 B.n89 71.676
R1154 B.n881 B.n880 71.676
R1155 B.n874 B.n91 71.676
R1156 B.n873 B.n872 71.676
R1157 B.n866 B.n93 71.676
R1158 B.n865 B.n864 71.676
R1159 B.n858 B.n95 71.676
R1160 B.n857 B.n856 71.676
R1161 B.n850 B.n97 71.676
R1162 B.n849 B.n848 71.676
R1163 B.n842 B.n99 71.676
R1164 B.n841 B.n840 71.676
R1165 B.n834 B.n101 71.676
R1166 B.n833 B.n832 71.676
R1167 B.n826 B.n103 71.676
R1168 B.n825 B.n824 71.676
R1169 B.n817 B.n105 71.676
R1170 B.n816 B.n815 71.676
R1171 B.n809 B.n109 71.676
R1172 B.n808 B.n807 71.676
R1173 B.n801 B.n111 71.676
R1174 B.n800 B.n115 71.676
R1175 B.n796 B.n795 71.676
R1176 B.n789 B.n117 71.676
R1177 B.n788 B.n787 71.676
R1178 B.n781 B.n119 71.676
R1179 B.n780 B.n779 71.676
R1180 B.n773 B.n121 71.676
R1181 B.n772 B.n771 71.676
R1182 B.n765 B.n123 71.676
R1183 B.n764 B.n763 71.676
R1184 B.n757 B.n125 71.676
R1185 B.n756 B.n755 71.676
R1186 B.n749 B.n127 71.676
R1187 B.n748 B.n747 71.676
R1188 B.n741 B.n129 71.676
R1189 B.n740 B.n739 71.676
R1190 B.n733 B.n131 71.676
R1191 B.n732 B.n731 71.676
R1192 B.n725 B.n133 71.676
R1193 B.n724 B.n723 71.676
R1194 B.n717 B.n135 71.676
R1195 B.n716 B.n715 71.676
R1196 B.n709 B.n137 71.676
R1197 B.n708 B.n707 71.676
R1198 B.n701 B.n139 71.676
R1199 B.n700 B.n699 71.676
R1200 B.n699 B.n698 71.676
R1201 B.n702 B.n701 71.676
R1202 B.n707 B.n706 71.676
R1203 B.n710 B.n709 71.676
R1204 B.n715 B.n714 71.676
R1205 B.n718 B.n717 71.676
R1206 B.n723 B.n722 71.676
R1207 B.n726 B.n725 71.676
R1208 B.n731 B.n730 71.676
R1209 B.n734 B.n733 71.676
R1210 B.n739 B.n738 71.676
R1211 B.n742 B.n741 71.676
R1212 B.n747 B.n746 71.676
R1213 B.n750 B.n749 71.676
R1214 B.n755 B.n754 71.676
R1215 B.n758 B.n757 71.676
R1216 B.n763 B.n762 71.676
R1217 B.n766 B.n765 71.676
R1218 B.n771 B.n770 71.676
R1219 B.n774 B.n773 71.676
R1220 B.n779 B.n778 71.676
R1221 B.n782 B.n781 71.676
R1222 B.n787 B.n786 71.676
R1223 B.n790 B.n789 71.676
R1224 B.n795 B.n794 71.676
R1225 B.n797 B.n115 71.676
R1226 B.n802 B.n801 71.676
R1227 B.n807 B.n806 71.676
R1228 B.n810 B.n809 71.676
R1229 B.n815 B.n814 71.676
R1230 B.n818 B.n817 71.676
R1231 B.n824 B.n823 71.676
R1232 B.n827 B.n826 71.676
R1233 B.n832 B.n831 71.676
R1234 B.n835 B.n834 71.676
R1235 B.n840 B.n839 71.676
R1236 B.n843 B.n842 71.676
R1237 B.n848 B.n847 71.676
R1238 B.n851 B.n850 71.676
R1239 B.n856 B.n855 71.676
R1240 B.n859 B.n858 71.676
R1241 B.n864 B.n863 71.676
R1242 B.n867 B.n866 71.676
R1243 B.n872 B.n871 71.676
R1244 B.n875 B.n874 71.676
R1245 B.n880 B.n879 71.676
R1246 B.n883 B.n882 71.676
R1247 B.n888 B.n887 71.676
R1248 B.n891 B.n890 71.676
R1249 B.n896 B.n895 71.676
R1250 B.n899 B.n898 71.676
R1251 B.n904 B.n903 71.676
R1252 B.n907 B.n906 71.676
R1253 B.n912 B.n911 71.676
R1254 B.n915 B.n914 71.676
R1255 B.n920 B.n919 71.676
R1256 B.n923 B.n922 71.676
R1257 B.n510 B.n509 71.676
R1258 B.n504 B.n224 71.676
R1259 B.n502 B.n501 71.676
R1260 B.n497 B.n496 71.676
R1261 B.n494 B.n493 71.676
R1262 B.n489 B.n488 71.676
R1263 B.n486 B.n485 71.676
R1264 B.n481 B.n480 71.676
R1265 B.n478 B.n477 71.676
R1266 B.n473 B.n472 71.676
R1267 B.n470 B.n469 71.676
R1268 B.n465 B.n464 71.676
R1269 B.n462 B.n461 71.676
R1270 B.n457 B.n456 71.676
R1271 B.n454 B.n453 71.676
R1272 B.n449 B.n448 71.676
R1273 B.n446 B.n445 71.676
R1274 B.n441 B.n440 71.676
R1275 B.n438 B.n437 71.676
R1276 B.n433 B.n432 71.676
R1277 B.n430 B.n429 71.676
R1278 B.n425 B.n424 71.676
R1279 B.n422 B.n421 71.676
R1280 B.n417 B.n416 71.676
R1281 B.n414 B.n413 71.676
R1282 B.n409 B.n408 71.676
R1283 B.n404 B.n252 71.676
R1284 B.n402 B.n401 71.676
R1285 B.n397 B.n396 71.676
R1286 B.n394 B.n393 71.676
R1287 B.n388 B.n387 71.676
R1288 B.n385 B.n384 71.676
R1289 B.n380 B.n379 71.676
R1290 B.n377 B.n376 71.676
R1291 B.n372 B.n371 71.676
R1292 B.n369 B.n368 71.676
R1293 B.n364 B.n363 71.676
R1294 B.n361 B.n360 71.676
R1295 B.n356 B.n355 71.676
R1296 B.n353 B.n352 71.676
R1297 B.n348 B.n347 71.676
R1298 B.n345 B.n344 71.676
R1299 B.n340 B.n339 71.676
R1300 B.n337 B.n336 71.676
R1301 B.n332 B.n331 71.676
R1302 B.n329 B.n328 71.676
R1303 B.n324 B.n323 71.676
R1304 B.n321 B.n320 71.676
R1305 B.n316 B.n315 71.676
R1306 B.n313 B.n312 71.676
R1307 B.n308 B.n307 71.676
R1308 B.n305 B.n304 71.676
R1309 B.n300 B.n299 71.676
R1310 B.n297 B.n296 71.676
R1311 B.n292 B.n291 71.676
R1312 B.n289 B.n288 71.676
R1313 B.n284 B.n220 71.676
R1314 B.n258 B.t16 70.8887
R1315 B.n113 B.t7 70.8887
R1316 B.n250 B.t10 70.8679
R1317 B.n107 B.t14 70.8679
R1318 B.n515 B.n221 59.9958
R1319 B.n928 B.n78 59.9958
R1320 B.n390 B.n258 59.5399
R1321 B.n251 B.n250 59.5399
R1322 B.n820 B.n107 59.5399
R1323 B.n114 B.n113 59.5399
R1324 B.n258 B.n257 55.6611
R1325 B.n250 B.n249 55.6611
R1326 B.n107 B.n106 55.6611
R1327 B.n113 B.n112 55.6611
R1328 B.n515 B.n217 35.476
R1329 B.n521 B.n217 35.476
R1330 B.n521 B.n213 35.476
R1331 B.n527 B.n213 35.476
R1332 B.n527 B.n209 35.476
R1333 B.n534 B.n209 35.476
R1334 B.n534 B.n533 35.476
R1335 B.n540 B.n202 35.476
R1336 B.n546 B.n202 35.476
R1337 B.n546 B.n198 35.476
R1338 B.n552 B.n198 35.476
R1339 B.n552 B.n194 35.476
R1340 B.n558 B.n194 35.476
R1341 B.n558 B.n190 35.476
R1342 B.n564 B.n190 35.476
R1343 B.n564 B.n186 35.476
R1344 B.n571 B.n186 35.476
R1345 B.n571 B.n570 35.476
R1346 B.n577 B.n179 35.476
R1347 B.n583 B.n179 35.476
R1348 B.n583 B.n175 35.476
R1349 B.n589 B.n175 35.476
R1350 B.n589 B.n171 35.476
R1351 B.n596 B.n171 35.476
R1352 B.n596 B.n595 35.476
R1353 B.n602 B.n164 35.476
R1354 B.n608 B.n164 35.476
R1355 B.n608 B.n160 35.476
R1356 B.n614 B.n160 35.476
R1357 B.n614 B.n156 35.476
R1358 B.n620 B.n156 35.476
R1359 B.n620 B.n152 35.476
R1360 B.n626 B.n152 35.476
R1361 B.n633 B.n148 35.476
R1362 B.n633 B.n144 35.476
R1363 B.n639 B.n144 35.476
R1364 B.n639 B.n4 35.476
R1365 B.n1010 B.n4 35.476
R1366 B.n1010 B.n1009 35.476
R1367 B.n1009 B.n1008 35.476
R1368 B.n1008 B.n8 35.476
R1369 B.n1002 B.n8 35.476
R1370 B.n1002 B.n1001 35.476
R1371 B.n1000 B.n15 35.476
R1372 B.n994 B.n15 35.476
R1373 B.n994 B.n993 35.476
R1374 B.n993 B.n992 35.476
R1375 B.n992 B.n22 35.476
R1376 B.n986 B.n22 35.476
R1377 B.n986 B.n985 35.476
R1378 B.n985 B.n984 35.476
R1379 B.n978 B.n32 35.476
R1380 B.n978 B.n977 35.476
R1381 B.n977 B.n976 35.476
R1382 B.n976 B.n36 35.476
R1383 B.n970 B.n36 35.476
R1384 B.n970 B.n969 35.476
R1385 B.n969 B.n968 35.476
R1386 B.n962 B.n46 35.476
R1387 B.n962 B.n961 35.476
R1388 B.n961 B.n960 35.476
R1389 B.n960 B.n50 35.476
R1390 B.n954 B.n50 35.476
R1391 B.n954 B.n953 35.476
R1392 B.n953 B.n952 35.476
R1393 B.n952 B.n57 35.476
R1394 B.n946 B.n57 35.476
R1395 B.n946 B.n945 35.476
R1396 B.n945 B.n944 35.476
R1397 B.n938 B.n67 35.476
R1398 B.n938 B.n937 35.476
R1399 B.n937 B.n936 35.476
R1400 B.n936 B.n71 35.476
R1401 B.n930 B.n71 35.476
R1402 B.n930 B.n929 35.476
R1403 B.n929 B.n928 35.476
R1404 B.n926 B.n925 32.3127
R1405 B.n696 B.n695 32.3127
R1406 B.n517 B.n219 32.3127
R1407 B.n513 B.n512 32.3127
R1408 B.t19 B.n148 29.2156
R1409 B.n1001 B.t0 29.2156
R1410 B.n595 B.t2 26.0854
R1411 B.n32 B.t1 26.0854
R1412 B.n577 B.t18 25.042
R1413 B.n968 B.t3 25.042
R1414 B.n533 B.t9 22.9552
R1415 B.n67 B.t5 22.9552
R1416 B B.n1012 18.0485
R1417 B.n540 B.t9 12.5212
R1418 B.n944 B.t5 12.5212
R1419 B.n925 B.n924 10.6151
R1420 B.n924 B.n80 10.6151
R1421 B.n918 B.n80 10.6151
R1422 B.n918 B.n917 10.6151
R1423 B.n917 B.n916 10.6151
R1424 B.n916 B.n82 10.6151
R1425 B.n910 B.n82 10.6151
R1426 B.n910 B.n909 10.6151
R1427 B.n909 B.n908 10.6151
R1428 B.n908 B.n84 10.6151
R1429 B.n902 B.n84 10.6151
R1430 B.n902 B.n901 10.6151
R1431 B.n901 B.n900 10.6151
R1432 B.n900 B.n86 10.6151
R1433 B.n894 B.n86 10.6151
R1434 B.n894 B.n893 10.6151
R1435 B.n893 B.n892 10.6151
R1436 B.n892 B.n88 10.6151
R1437 B.n886 B.n88 10.6151
R1438 B.n886 B.n885 10.6151
R1439 B.n885 B.n884 10.6151
R1440 B.n884 B.n90 10.6151
R1441 B.n878 B.n90 10.6151
R1442 B.n878 B.n877 10.6151
R1443 B.n877 B.n876 10.6151
R1444 B.n876 B.n92 10.6151
R1445 B.n870 B.n92 10.6151
R1446 B.n870 B.n869 10.6151
R1447 B.n869 B.n868 10.6151
R1448 B.n868 B.n94 10.6151
R1449 B.n862 B.n94 10.6151
R1450 B.n862 B.n861 10.6151
R1451 B.n861 B.n860 10.6151
R1452 B.n860 B.n96 10.6151
R1453 B.n854 B.n96 10.6151
R1454 B.n854 B.n853 10.6151
R1455 B.n853 B.n852 10.6151
R1456 B.n852 B.n98 10.6151
R1457 B.n846 B.n98 10.6151
R1458 B.n846 B.n845 10.6151
R1459 B.n845 B.n844 10.6151
R1460 B.n844 B.n100 10.6151
R1461 B.n838 B.n100 10.6151
R1462 B.n838 B.n837 10.6151
R1463 B.n837 B.n836 10.6151
R1464 B.n836 B.n102 10.6151
R1465 B.n830 B.n102 10.6151
R1466 B.n830 B.n829 10.6151
R1467 B.n829 B.n828 10.6151
R1468 B.n828 B.n104 10.6151
R1469 B.n822 B.n104 10.6151
R1470 B.n822 B.n821 10.6151
R1471 B.n819 B.n108 10.6151
R1472 B.n813 B.n108 10.6151
R1473 B.n813 B.n812 10.6151
R1474 B.n812 B.n811 10.6151
R1475 B.n811 B.n110 10.6151
R1476 B.n805 B.n110 10.6151
R1477 B.n805 B.n804 10.6151
R1478 B.n804 B.n803 10.6151
R1479 B.n799 B.n798 10.6151
R1480 B.n798 B.n116 10.6151
R1481 B.n793 B.n116 10.6151
R1482 B.n793 B.n792 10.6151
R1483 B.n792 B.n791 10.6151
R1484 B.n791 B.n118 10.6151
R1485 B.n785 B.n118 10.6151
R1486 B.n785 B.n784 10.6151
R1487 B.n784 B.n783 10.6151
R1488 B.n783 B.n120 10.6151
R1489 B.n777 B.n120 10.6151
R1490 B.n777 B.n776 10.6151
R1491 B.n776 B.n775 10.6151
R1492 B.n775 B.n122 10.6151
R1493 B.n769 B.n122 10.6151
R1494 B.n769 B.n768 10.6151
R1495 B.n768 B.n767 10.6151
R1496 B.n767 B.n124 10.6151
R1497 B.n761 B.n124 10.6151
R1498 B.n761 B.n760 10.6151
R1499 B.n760 B.n759 10.6151
R1500 B.n759 B.n126 10.6151
R1501 B.n753 B.n126 10.6151
R1502 B.n753 B.n752 10.6151
R1503 B.n752 B.n751 10.6151
R1504 B.n751 B.n128 10.6151
R1505 B.n745 B.n128 10.6151
R1506 B.n745 B.n744 10.6151
R1507 B.n744 B.n743 10.6151
R1508 B.n743 B.n130 10.6151
R1509 B.n737 B.n130 10.6151
R1510 B.n737 B.n736 10.6151
R1511 B.n736 B.n735 10.6151
R1512 B.n735 B.n132 10.6151
R1513 B.n729 B.n132 10.6151
R1514 B.n729 B.n728 10.6151
R1515 B.n728 B.n727 10.6151
R1516 B.n727 B.n134 10.6151
R1517 B.n721 B.n134 10.6151
R1518 B.n721 B.n720 10.6151
R1519 B.n720 B.n719 10.6151
R1520 B.n719 B.n136 10.6151
R1521 B.n713 B.n136 10.6151
R1522 B.n713 B.n712 10.6151
R1523 B.n712 B.n711 10.6151
R1524 B.n711 B.n138 10.6151
R1525 B.n705 B.n138 10.6151
R1526 B.n705 B.n704 10.6151
R1527 B.n704 B.n703 10.6151
R1528 B.n703 B.n140 10.6151
R1529 B.n697 B.n140 10.6151
R1530 B.n697 B.n696 10.6151
R1531 B.n518 B.n517 10.6151
R1532 B.n519 B.n518 10.6151
R1533 B.n519 B.n211 10.6151
R1534 B.n529 B.n211 10.6151
R1535 B.n530 B.n529 10.6151
R1536 B.n531 B.n530 10.6151
R1537 B.n531 B.n204 10.6151
R1538 B.n542 B.n204 10.6151
R1539 B.n543 B.n542 10.6151
R1540 B.n544 B.n543 10.6151
R1541 B.n544 B.n196 10.6151
R1542 B.n554 B.n196 10.6151
R1543 B.n555 B.n554 10.6151
R1544 B.n556 B.n555 10.6151
R1545 B.n556 B.n188 10.6151
R1546 B.n566 B.n188 10.6151
R1547 B.n567 B.n566 10.6151
R1548 B.n568 B.n567 10.6151
R1549 B.n568 B.n181 10.6151
R1550 B.n579 B.n181 10.6151
R1551 B.n580 B.n579 10.6151
R1552 B.n581 B.n580 10.6151
R1553 B.n581 B.n173 10.6151
R1554 B.n591 B.n173 10.6151
R1555 B.n592 B.n591 10.6151
R1556 B.n593 B.n592 10.6151
R1557 B.n593 B.n166 10.6151
R1558 B.n604 B.n166 10.6151
R1559 B.n605 B.n604 10.6151
R1560 B.n606 B.n605 10.6151
R1561 B.n606 B.n158 10.6151
R1562 B.n616 B.n158 10.6151
R1563 B.n617 B.n616 10.6151
R1564 B.n618 B.n617 10.6151
R1565 B.n618 B.n150 10.6151
R1566 B.n628 B.n150 10.6151
R1567 B.n629 B.n628 10.6151
R1568 B.n631 B.n629 10.6151
R1569 B.n631 B.n630 10.6151
R1570 B.n630 B.n142 10.6151
R1571 B.n642 B.n142 10.6151
R1572 B.n643 B.n642 10.6151
R1573 B.n644 B.n643 10.6151
R1574 B.n645 B.n644 10.6151
R1575 B.n647 B.n645 10.6151
R1576 B.n648 B.n647 10.6151
R1577 B.n649 B.n648 10.6151
R1578 B.n650 B.n649 10.6151
R1579 B.n652 B.n650 10.6151
R1580 B.n653 B.n652 10.6151
R1581 B.n654 B.n653 10.6151
R1582 B.n655 B.n654 10.6151
R1583 B.n657 B.n655 10.6151
R1584 B.n658 B.n657 10.6151
R1585 B.n659 B.n658 10.6151
R1586 B.n660 B.n659 10.6151
R1587 B.n662 B.n660 10.6151
R1588 B.n663 B.n662 10.6151
R1589 B.n664 B.n663 10.6151
R1590 B.n665 B.n664 10.6151
R1591 B.n667 B.n665 10.6151
R1592 B.n668 B.n667 10.6151
R1593 B.n669 B.n668 10.6151
R1594 B.n670 B.n669 10.6151
R1595 B.n672 B.n670 10.6151
R1596 B.n673 B.n672 10.6151
R1597 B.n674 B.n673 10.6151
R1598 B.n675 B.n674 10.6151
R1599 B.n677 B.n675 10.6151
R1600 B.n678 B.n677 10.6151
R1601 B.n679 B.n678 10.6151
R1602 B.n680 B.n679 10.6151
R1603 B.n682 B.n680 10.6151
R1604 B.n683 B.n682 10.6151
R1605 B.n684 B.n683 10.6151
R1606 B.n685 B.n684 10.6151
R1607 B.n687 B.n685 10.6151
R1608 B.n688 B.n687 10.6151
R1609 B.n689 B.n688 10.6151
R1610 B.n690 B.n689 10.6151
R1611 B.n692 B.n690 10.6151
R1612 B.n693 B.n692 10.6151
R1613 B.n694 B.n693 10.6151
R1614 B.n695 B.n694 10.6151
R1615 B.n512 B.n511 10.6151
R1616 B.n511 B.n223 10.6151
R1617 B.n506 B.n223 10.6151
R1618 B.n506 B.n505 10.6151
R1619 B.n505 B.n225 10.6151
R1620 B.n500 B.n225 10.6151
R1621 B.n500 B.n499 10.6151
R1622 B.n499 B.n498 10.6151
R1623 B.n498 B.n227 10.6151
R1624 B.n492 B.n227 10.6151
R1625 B.n492 B.n491 10.6151
R1626 B.n491 B.n490 10.6151
R1627 B.n490 B.n229 10.6151
R1628 B.n484 B.n229 10.6151
R1629 B.n484 B.n483 10.6151
R1630 B.n483 B.n482 10.6151
R1631 B.n482 B.n231 10.6151
R1632 B.n476 B.n231 10.6151
R1633 B.n476 B.n475 10.6151
R1634 B.n475 B.n474 10.6151
R1635 B.n474 B.n233 10.6151
R1636 B.n468 B.n233 10.6151
R1637 B.n468 B.n467 10.6151
R1638 B.n467 B.n466 10.6151
R1639 B.n466 B.n235 10.6151
R1640 B.n460 B.n235 10.6151
R1641 B.n460 B.n459 10.6151
R1642 B.n459 B.n458 10.6151
R1643 B.n458 B.n237 10.6151
R1644 B.n452 B.n237 10.6151
R1645 B.n452 B.n451 10.6151
R1646 B.n451 B.n450 10.6151
R1647 B.n450 B.n239 10.6151
R1648 B.n444 B.n239 10.6151
R1649 B.n444 B.n443 10.6151
R1650 B.n443 B.n442 10.6151
R1651 B.n442 B.n241 10.6151
R1652 B.n436 B.n241 10.6151
R1653 B.n436 B.n435 10.6151
R1654 B.n435 B.n434 10.6151
R1655 B.n434 B.n243 10.6151
R1656 B.n428 B.n243 10.6151
R1657 B.n428 B.n427 10.6151
R1658 B.n427 B.n426 10.6151
R1659 B.n426 B.n245 10.6151
R1660 B.n420 B.n245 10.6151
R1661 B.n420 B.n419 10.6151
R1662 B.n419 B.n418 10.6151
R1663 B.n418 B.n247 10.6151
R1664 B.n412 B.n247 10.6151
R1665 B.n412 B.n411 10.6151
R1666 B.n411 B.n410 10.6151
R1667 B.n406 B.n405 10.6151
R1668 B.n405 B.n253 10.6151
R1669 B.n400 B.n253 10.6151
R1670 B.n400 B.n399 10.6151
R1671 B.n399 B.n398 10.6151
R1672 B.n398 B.n255 10.6151
R1673 B.n392 B.n255 10.6151
R1674 B.n392 B.n391 10.6151
R1675 B.n389 B.n259 10.6151
R1676 B.n383 B.n259 10.6151
R1677 B.n383 B.n382 10.6151
R1678 B.n382 B.n381 10.6151
R1679 B.n381 B.n261 10.6151
R1680 B.n375 B.n261 10.6151
R1681 B.n375 B.n374 10.6151
R1682 B.n374 B.n373 10.6151
R1683 B.n373 B.n263 10.6151
R1684 B.n367 B.n263 10.6151
R1685 B.n367 B.n366 10.6151
R1686 B.n366 B.n365 10.6151
R1687 B.n365 B.n265 10.6151
R1688 B.n359 B.n265 10.6151
R1689 B.n359 B.n358 10.6151
R1690 B.n358 B.n357 10.6151
R1691 B.n357 B.n267 10.6151
R1692 B.n351 B.n267 10.6151
R1693 B.n351 B.n350 10.6151
R1694 B.n350 B.n349 10.6151
R1695 B.n349 B.n269 10.6151
R1696 B.n343 B.n269 10.6151
R1697 B.n343 B.n342 10.6151
R1698 B.n342 B.n341 10.6151
R1699 B.n341 B.n271 10.6151
R1700 B.n335 B.n271 10.6151
R1701 B.n335 B.n334 10.6151
R1702 B.n334 B.n333 10.6151
R1703 B.n333 B.n273 10.6151
R1704 B.n327 B.n273 10.6151
R1705 B.n327 B.n326 10.6151
R1706 B.n326 B.n325 10.6151
R1707 B.n325 B.n275 10.6151
R1708 B.n319 B.n275 10.6151
R1709 B.n319 B.n318 10.6151
R1710 B.n318 B.n317 10.6151
R1711 B.n317 B.n277 10.6151
R1712 B.n311 B.n277 10.6151
R1713 B.n311 B.n310 10.6151
R1714 B.n310 B.n309 10.6151
R1715 B.n309 B.n279 10.6151
R1716 B.n303 B.n279 10.6151
R1717 B.n303 B.n302 10.6151
R1718 B.n302 B.n301 10.6151
R1719 B.n301 B.n281 10.6151
R1720 B.n295 B.n281 10.6151
R1721 B.n295 B.n294 10.6151
R1722 B.n294 B.n293 10.6151
R1723 B.n293 B.n283 10.6151
R1724 B.n287 B.n283 10.6151
R1725 B.n287 B.n286 10.6151
R1726 B.n286 B.n219 10.6151
R1727 B.n513 B.n215 10.6151
R1728 B.n523 B.n215 10.6151
R1729 B.n524 B.n523 10.6151
R1730 B.n525 B.n524 10.6151
R1731 B.n525 B.n207 10.6151
R1732 B.n536 B.n207 10.6151
R1733 B.n537 B.n536 10.6151
R1734 B.n538 B.n537 10.6151
R1735 B.n538 B.n200 10.6151
R1736 B.n548 B.n200 10.6151
R1737 B.n549 B.n548 10.6151
R1738 B.n550 B.n549 10.6151
R1739 B.n550 B.n192 10.6151
R1740 B.n560 B.n192 10.6151
R1741 B.n561 B.n560 10.6151
R1742 B.n562 B.n561 10.6151
R1743 B.n562 B.n184 10.6151
R1744 B.n573 B.n184 10.6151
R1745 B.n574 B.n573 10.6151
R1746 B.n575 B.n574 10.6151
R1747 B.n575 B.n177 10.6151
R1748 B.n585 B.n177 10.6151
R1749 B.n586 B.n585 10.6151
R1750 B.n587 B.n586 10.6151
R1751 B.n587 B.n169 10.6151
R1752 B.n598 B.n169 10.6151
R1753 B.n599 B.n598 10.6151
R1754 B.n600 B.n599 10.6151
R1755 B.n600 B.n162 10.6151
R1756 B.n610 B.n162 10.6151
R1757 B.n611 B.n610 10.6151
R1758 B.n612 B.n611 10.6151
R1759 B.n612 B.n154 10.6151
R1760 B.n622 B.n154 10.6151
R1761 B.n623 B.n622 10.6151
R1762 B.n624 B.n623 10.6151
R1763 B.n624 B.n146 10.6151
R1764 B.n635 B.n146 10.6151
R1765 B.n636 B.n635 10.6151
R1766 B.n637 B.n636 10.6151
R1767 B.n637 B.n0 10.6151
R1768 B.n1006 B.n1 10.6151
R1769 B.n1006 B.n1005 10.6151
R1770 B.n1005 B.n1004 10.6151
R1771 B.n1004 B.n10 10.6151
R1772 B.n998 B.n10 10.6151
R1773 B.n998 B.n997 10.6151
R1774 B.n997 B.n996 10.6151
R1775 B.n996 B.n17 10.6151
R1776 B.n990 B.n17 10.6151
R1777 B.n990 B.n989 10.6151
R1778 B.n989 B.n988 10.6151
R1779 B.n988 B.n24 10.6151
R1780 B.n982 B.n24 10.6151
R1781 B.n982 B.n981 10.6151
R1782 B.n981 B.n980 10.6151
R1783 B.n980 B.n30 10.6151
R1784 B.n974 B.n30 10.6151
R1785 B.n974 B.n973 10.6151
R1786 B.n973 B.n972 10.6151
R1787 B.n972 B.n38 10.6151
R1788 B.n966 B.n38 10.6151
R1789 B.n966 B.n965 10.6151
R1790 B.n965 B.n964 10.6151
R1791 B.n964 B.n44 10.6151
R1792 B.n958 B.n44 10.6151
R1793 B.n958 B.n957 10.6151
R1794 B.n957 B.n956 10.6151
R1795 B.n956 B.n52 10.6151
R1796 B.n950 B.n52 10.6151
R1797 B.n950 B.n949 10.6151
R1798 B.n949 B.n948 10.6151
R1799 B.n948 B.n59 10.6151
R1800 B.n942 B.n59 10.6151
R1801 B.n942 B.n941 10.6151
R1802 B.n941 B.n940 10.6151
R1803 B.n940 B.n65 10.6151
R1804 B.n934 B.n65 10.6151
R1805 B.n934 B.n933 10.6151
R1806 B.n933 B.n932 10.6151
R1807 B.n932 B.n73 10.6151
R1808 B.n926 B.n73 10.6151
R1809 B.n570 B.t18 10.4345
R1810 B.n46 B.t3 10.4345
R1811 B.n602 B.t2 9.39106
R1812 B.n984 B.t1 9.39106
R1813 B.n820 B.n819 6.4005
R1814 B.n803 B.n114 6.4005
R1815 B.n406 B.n251 6.4005
R1816 B.n391 B.n390 6.4005
R1817 B.n626 B.t19 6.26087
R1818 B.t0 B.n1000 6.26087
R1819 B.n821 B.n820 4.21513
R1820 B.n799 B.n114 4.21513
R1821 B.n410 B.n251 4.21513
R1822 B.n390 B.n389 4.21513
R1823 B.n1012 B.n0 2.81026
R1824 B.n1012 B.n1 2.81026
R1825 VN.n4 VN.t5 182.352
R1826 VN.n20 VN.t3 182.352
R1827 VN.n29 VN.n16 161.3
R1828 VN.n28 VN.n27 161.3
R1829 VN.n26 VN.n17 161.3
R1830 VN.n25 VN.n24 161.3
R1831 VN.n23 VN.n18 161.3
R1832 VN.n22 VN.n21 161.3
R1833 VN.n13 VN.n0 161.3
R1834 VN.n12 VN.n11 161.3
R1835 VN.n10 VN.n1 161.3
R1836 VN.n9 VN.n8 161.3
R1837 VN.n7 VN.n2 161.3
R1838 VN.n6 VN.n5 161.3
R1839 VN.n3 VN.t2 150.008
R1840 VN.n14 VN.t0 150.008
R1841 VN.n19 VN.t1 150.008
R1842 VN.n30 VN.t4 150.008
R1843 VN.n15 VN.n14 104.885
R1844 VN.n31 VN.n30 104.885
R1845 VN.n4 VN.n3 59.9599
R1846 VN.n20 VN.n19 59.9599
R1847 VN.n8 VN.n1 56.5193
R1848 VN.n24 VN.n17 56.5193
R1849 VN VN.n31 51.5474
R1850 VN.n7 VN.n6 24.4675
R1851 VN.n8 VN.n7 24.4675
R1852 VN.n12 VN.n1 24.4675
R1853 VN.n13 VN.n12 24.4675
R1854 VN.n24 VN.n23 24.4675
R1855 VN.n23 VN.n22 24.4675
R1856 VN.n29 VN.n28 24.4675
R1857 VN.n28 VN.n17 24.4675
R1858 VN.n6 VN.n3 12.234
R1859 VN.n22 VN.n19 12.234
R1860 VN.n21 VN.n20 7.1096
R1861 VN.n5 VN.n4 7.1096
R1862 VN.n14 VN.n13 5.87258
R1863 VN.n30 VN.n29 5.87258
R1864 VN.n31 VN.n16 0.278367
R1865 VN.n15 VN.n0 0.278367
R1866 VN.n27 VN.n16 0.189894
R1867 VN.n27 VN.n26 0.189894
R1868 VN.n26 VN.n25 0.189894
R1869 VN.n25 VN.n18 0.189894
R1870 VN.n21 VN.n18 0.189894
R1871 VN.n5 VN.n2 0.189894
R1872 VN.n9 VN.n2 0.189894
R1873 VN.n10 VN.n9 0.189894
R1874 VN.n11 VN.n10 0.189894
R1875 VN.n11 VN.n0 0.189894
R1876 VN VN.n15 0.153454
R1877 VDD2.n1 VDD2.t0 65.6062
R1878 VDD2.n2 VDD2.t1 63.8061
R1879 VDD2.n1 VDD2.n0 63.1167
R1880 VDD2 VDD2.n3 63.1139
R1881 VDD2.n2 VDD2.n1 45.3856
R1882 VDD2 VDD2.n2 1.91429
R1883 VDD2.n3 VDD2.t4 1.25287
R1884 VDD2.n3 VDD2.t2 1.25287
R1885 VDD2.n0 VDD2.t3 1.25287
R1886 VDD2.n0 VDD2.t5 1.25287
C0 VDD2 VTAIL 9.16371f
C1 VN VDD1 0.150757f
C2 VP VDD2 0.45365f
C3 VN VDD2 8.69789f
C4 VP VTAIL 8.68818f
C5 VN VTAIL 8.67383f
C6 VN VP 7.57663f
C7 VDD2 VDD1 1.38462f
C8 VDD1 VTAIL 9.11425f
C9 VP VDD1 8.99689f
C10 VDD2 B 6.619783f
C11 VDD1 B 6.938702f
C12 VTAIL B 9.29318f
C13 VN B 13.05668f
C14 VP B 11.603004f
C15 VDD2.t0 B 3.09282f
C16 VDD2.t3 B 0.266176f
C17 VDD2.t5 B 0.266176f
C18 VDD2.n0 B 2.41684f
C19 VDD2.n1 B 2.65366f
C20 VDD2.t1 B 3.08289f
C21 VDD2.n2 B 2.61542f
C22 VDD2.t4 B 0.266176f
C23 VDD2.t2 B 0.266176f
C24 VDD2.n3 B 2.41681f
C25 VN.n0 B 0.030268f
C26 VN.t0 B 2.52814f
C27 VN.n1 B 0.037675f
C28 VN.n2 B 0.022958f
C29 VN.t2 B 2.52814f
C30 VN.n3 B 0.947592f
C31 VN.t5 B 2.70918f
C32 VN.n4 B 0.930333f
C33 VN.n5 B 0.220247f
C34 VN.n6 B 0.032226f
C35 VN.n7 B 0.042788f
C36 VN.n8 B 0.029359f
C37 VN.n9 B 0.022958f
C38 VN.n10 B 0.022958f
C39 VN.n11 B 0.022958f
C40 VN.n12 B 0.042788f
C41 VN.n13 B 0.026733f
C42 VN.n14 B 0.952408f
C43 VN.n15 B 0.039097f
C44 VN.n16 B 0.030268f
C45 VN.t4 B 2.52814f
C46 VN.n17 B 0.037675f
C47 VN.n18 B 0.022958f
C48 VN.t1 B 2.52814f
C49 VN.n19 B 0.947592f
C50 VN.t3 B 2.70918f
C51 VN.n20 B 0.930333f
C52 VN.n21 B 0.220247f
C53 VN.n22 B 0.032226f
C54 VN.n23 B 0.042788f
C55 VN.n24 B 0.029359f
C56 VN.n25 B 0.022958f
C57 VN.n26 B 0.022958f
C58 VN.n27 B 0.022958f
C59 VN.n28 B 0.042788f
C60 VN.n29 B 0.026733f
C61 VN.n30 B 0.952408f
C62 VN.n31 B 1.33838f
C63 VTAIL.t0 B 0.285844f
C64 VTAIL.t1 B 0.285844f
C65 VTAIL.n0 B 2.52549f
C66 VTAIL.n1 B 0.397206f
C67 VTAIL.t7 B 3.22482f
C68 VTAIL.n2 B 0.609959f
C69 VTAIL.t4 B 0.285844f
C70 VTAIL.t8 B 0.285844f
C71 VTAIL.n3 B 2.52549f
C72 VTAIL.n4 B 2.08425f
C73 VTAIL.t11 B 0.285844f
C74 VTAIL.t2 B 0.285844f
C75 VTAIL.n5 B 2.52549f
C76 VTAIL.n6 B 2.08425f
C77 VTAIL.t10 B 3.22484f
C78 VTAIL.n7 B 0.609938f
C79 VTAIL.t5 B 0.285844f
C80 VTAIL.t9 B 0.285844f
C81 VTAIL.n8 B 2.52549f
C82 VTAIL.n9 B 0.529712f
C83 VTAIL.t6 B 3.22482f
C84 VTAIL.n10 B 1.98209f
C85 VTAIL.t3 B 3.22482f
C86 VTAIL.n11 B 1.9322f
C87 VDD1.t3 B 3.11454f
C88 VDD1.t4 B 3.11369f
C89 VDD1.t0 B 0.267972f
C90 VDD1.t1 B 0.267972f
C91 VDD1.n0 B 2.43315f
C92 VDD1.n1 B 2.77897f
C93 VDD1.t2 B 0.267972f
C94 VDD1.t5 B 0.267972f
C95 VDD1.n2 B 2.42962f
C96 VDD1.n3 B 2.62558f
C97 VP.n0 B 0.030671f
C98 VP.t2 B 2.56179f
C99 VP.n1 B 0.038177f
C100 VP.n2 B 0.023264f
C101 VP.t1 B 2.56179f
C102 VP.n3 B 0.894103f
C103 VP.n4 B 0.023264f
C104 VP.n5 B 0.038177f
C105 VP.n6 B 0.030671f
C106 VP.t5 B 2.56179f
C107 VP.n7 B 0.030671f
C108 VP.t3 B 2.56179f
C109 VP.n8 B 0.038177f
C110 VP.n9 B 0.023264f
C111 VP.t0 B 2.56179f
C112 VP.n10 B 0.960203f
C113 VP.t4 B 2.74524f
C114 VP.n11 B 0.942714f
C115 VP.n12 B 0.223178f
C116 VP.n13 B 0.032655f
C117 VP.n14 B 0.043358f
C118 VP.n15 B 0.029749f
C119 VP.n16 B 0.023264f
C120 VP.n17 B 0.023264f
C121 VP.n18 B 0.023264f
C122 VP.n19 B 0.043358f
C123 VP.n20 B 0.027089f
C124 VP.n21 B 0.965083f
C125 VP.n22 B 1.34374f
C126 VP.n23 B 1.36005f
C127 VP.n24 B 0.965083f
C128 VP.n25 B 0.027089f
C129 VP.n26 B 0.043358f
C130 VP.n27 B 0.023264f
C131 VP.n28 B 0.023264f
C132 VP.n29 B 0.023264f
C133 VP.n30 B 0.029749f
C134 VP.n31 B 0.043358f
C135 VP.n32 B 0.032655f
C136 VP.n33 B 0.023264f
C137 VP.n34 B 0.023264f
C138 VP.n35 B 0.032655f
C139 VP.n36 B 0.043358f
C140 VP.n37 B 0.029749f
C141 VP.n38 B 0.023264f
C142 VP.n39 B 0.023264f
C143 VP.n40 B 0.023264f
C144 VP.n41 B 0.043358f
C145 VP.n42 B 0.027089f
C146 VP.n43 B 0.965083f
C147 VP.n44 B 0.039617f
.ends

