* NGSPICE file created from diff_pair_sample_1761.ext - technology: sky130A

.subckt diff_pair_sample_1761 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t3 w_n1790_n3530# sky130_fd_pr__pfet_01v8 ad=4.9959 pd=26.4 as=2.11365 ps=13.14 w=12.81 l=0.49
X1 VTAIL.t4 VP.t0 VDD1.t7 w_n1790_n3530# sky130_fd_pr__pfet_01v8 ad=4.9959 pd=26.4 as=2.11365 ps=13.14 w=12.81 l=0.49
X2 B.t11 B.t9 B.t10 w_n1790_n3530# sky130_fd_pr__pfet_01v8 ad=4.9959 pd=26.4 as=0 ps=0 w=12.81 l=0.49
X3 VDD2.t4 VN.t1 VTAIL.t14 w_n1790_n3530# sky130_fd_pr__pfet_01v8 ad=2.11365 pd=13.14 as=2.11365 ps=13.14 w=12.81 l=0.49
X4 B.t8 B.t6 B.t7 w_n1790_n3530# sky130_fd_pr__pfet_01v8 ad=4.9959 pd=26.4 as=0 ps=0 w=12.81 l=0.49
X5 VDD2.t1 VN.t2 VTAIL.t13 w_n1790_n3530# sky130_fd_pr__pfet_01v8 ad=2.11365 pd=13.14 as=4.9959 ps=26.4 w=12.81 l=0.49
X6 VDD2.t2 VN.t3 VTAIL.t12 w_n1790_n3530# sky130_fd_pr__pfet_01v8 ad=2.11365 pd=13.14 as=2.11365 ps=13.14 w=12.81 l=0.49
X7 B.t5 B.t3 B.t4 w_n1790_n3530# sky130_fd_pr__pfet_01v8 ad=4.9959 pd=26.4 as=0 ps=0 w=12.81 l=0.49
X8 B.t2 B.t0 B.t1 w_n1790_n3530# sky130_fd_pr__pfet_01v8 ad=4.9959 pd=26.4 as=0 ps=0 w=12.81 l=0.49
X9 VTAIL.t11 VN.t4 VDD2.t6 w_n1790_n3530# sky130_fd_pr__pfet_01v8 ad=4.9959 pd=26.4 as=2.11365 ps=13.14 w=12.81 l=0.49
X10 VTAIL.t3 VP.t1 VDD1.t6 w_n1790_n3530# sky130_fd_pr__pfet_01v8 ad=2.11365 pd=13.14 as=2.11365 ps=13.14 w=12.81 l=0.49
X11 VDD1.t5 VP.t2 VTAIL.t1 w_n1790_n3530# sky130_fd_pr__pfet_01v8 ad=2.11365 pd=13.14 as=2.11365 ps=13.14 w=12.81 l=0.49
X12 VTAIL.t10 VN.t5 VDD2.t5 w_n1790_n3530# sky130_fd_pr__pfet_01v8 ad=2.11365 pd=13.14 as=2.11365 ps=13.14 w=12.81 l=0.49
X13 VTAIL.t9 VN.t6 VDD2.t7 w_n1790_n3530# sky130_fd_pr__pfet_01v8 ad=2.11365 pd=13.14 as=2.11365 ps=13.14 w=12.81 l=0.49
X14 VTAIL.t6 VP.t3 VDD1.t4 w_n1790_n3530# sky130_fd_pr__pfet_01v8 ad=2.11365 pd=13.14 as=2.11365 ps=13.14 w=12.81 l=0.49
X15 VTAIL.t2 VP.t4 VDD1.t3 w_n1790_n3530# sky130_fd_pr__pfet_01v8 ad=4.9959 pd=26.4 as=2.11365 ps=13.14 w=12.81 l=0.49
X16 VDD1.t2 VP.t5 VTAIL.t7 w_n1790_n3530# sky130_fd_pr__pfet_01v8 ad=2.11365 pd=13.14 as=4.9959 ps=26.4 w=12.81 l=0.49
X17 VDD1.t1 VP.t6 VTAIL.t0 w_n1790_n3530# sky130_fd_pr__pfet_01v8 ad=2.11365 pd=13.14 as=2.11365 ps=13.14 w=12.81 l=0.49
X18 VDD2.t0 VN.t7 VTAIL.t8 w_n1790_n3530# sky130_fd_pr__pfet_01v8 ad=2.11365 pd=13.14 as=4.9959 ps=26.4 w=12.81 l=0.49
X19 VDD1.t0 VP.t7 VTAIL.t5 w_n1790_n3530# sky130_fd_pr__pfet_01v8 ad=2.11365 pd=13.14 as=4.9959 ps=26.4 w=12.81 l=0.49
R0 VN.n2 VN.t0 731.687
R1 VN.n10 VN.t2 731.687
R2 VN.n1 VN.t1 710.705
R3 VN.n5 VN.t6 710.705
R4 VN.n6 VN.t7 710.705
R5 VN.n9 VN.t5 710.705
R6 VN.n13 VN.t3 710.705
R7 VN.n14 VN.t4 710.705
R8 VN.n7 VN.n6 161.3
R9 VN.n15 VN.n14 161.3
R10 VN.n13 VN.n8 161.3
R11 VN.n12 VN.n11 161.3
R12 VN.n5 VN.n0 161.3
R13 VN.n4 VN.n3 161.3
R14 VN.n11 VN.n10 70.4033
R15 VN.n3 VN.n2 70.4033
R16 VN.n6 VN.n5 48.2005
R17 VN.n14 VN.n13 48.2005
R18 VN VN.n15 42.0933
R19 VN.n4 VN.n1 24.1005
R20 VN.n5 VN.n4 24.1005
R21 VN.n13 VN.n12 24.1005
R22 VN.n12 VN.n9 24.1005
R23 VN.n10 VN.n9 20.9576
R24 VN.n2 VN.n1 20.9576
R25 VN.n15 VN.n8 0.189894
R26 VN.n11 VN.n8 0.189894
R27 VN.n3 VN.n0 0.189894
R28 VN.n7 VN.n0 0.189894
R29 VN VN.n7 0.0516364
R30 VDD2.n2 VDD2.n1 72.7276
R31 VDD2.n2 VDD2.n0 72.7276
R32 VDD2 VDD2.n5 72.7246
R33 VDD2.n4 VDD2.n3 72.4295
R34 VDD2.n4 VDD2.n2 37.9394
R35 VDD2.n5 VDD2.t5 2.53797
R36 VDD2.n5 VDD2.t1 2.53797
R37 VDD2.n3 VDD2.t6 2.53797
R38 VDD2.n3 VDD2.t2 2.53797
R39 VDD2.n1 VDD2.t7 2.53797
R40 VDD2.n1 VDD2.t0 2.53797
R41 VDD2.n0 VDD2.t3 2.53797
R42 VDD2.n0 VDD2.t4 2.53797
R43 VDD2 VDD2.n4 0.412138
R44 VTAIL.n562 VTAIL.n498 756.745
R45 VTAIL.n66 VTAIL.n2 756.745
R46 VTAIL.n136 VTAIL.n72 756.745
R47 VTAIL.n208 VTAIL.n144 756.745
R48 VTAIL.n492 VTAIL.n428 756.745
R49 VTAIL.n420 VTAIL.n356 756.745
R50 VTAIL.n350 VTAIL.n286 756.745
R51 VTAIL.n278 VTAIL.n214 756.745
R52 VTAIL.n521 VTAIL.n520 585
R53 VTAIL.n518 VTAIL.n517 585
R54 VTAIL.n527 VTAIL.n526 585
R55 VTAIL.n529 VTAIL.n528 585
R56 VTAIL.n514 VTAIL.n513 585
R57 VTAIL.n535 VTAIL.n534 585
R58 VTAIL.n538 VTAIL.n537 585
R59 VTAIL.n536 VTAIL.n510 585
R60 VTAIL.n543 VTAIL.n509 585
R61 VTAIL.n545 VTAIL.n544 585
R62 VTAIL.n547 VTAIL.n546 585
R63 VTAIL.n506 VTAIL.n505 585
R64 VTAIL.n553 VTAIL.n552 585
R65 VTAIL.n555 VTAIL.n554 585
R66 VTAIL.n502 VTAIL.n501 585
R67 VTAIL.n561 VTAIL.n560 585
R68 VTAIL.n563 VTAIL.n562 585
R69 VTAIL.n25 VTAIL.n24 585
R70 VTAIL.n22 VTAIL.n21 585
R71 VTAIL.n31 VTAIL.n30 585
R72 VTAIL.n33 VTAIL.n32 585
R73 VTAIL.n18 VTAIL.n17 585
R74 VTAIL.n39 VTAIL.n38 585
R75 VTAIL.n42 VTAIL.n41 585
R76 VTAIL.n40 VTAIL.n14 585
R77 VTAIL.n47 VTAIL.n13 585
R78 VTAIL.n49 VTAIL.n48 585
R79 VTAIL.n51 VTAIL.n50 585
R80 VTAIL.n10 VTAIL.n9 585
R81 VTAIL.n57 VTAIL.n56 585
R82 VTAIL.n59 VTAIL.n58 585
R83 VTAIL.n6 VTAIL.n5 585
R84 VTAIL.n65 VTAIL.n64 585
R85 VTAIL.n67 VTAIL.n66 585
R86 VTAIL.n95 VTAIL.n94 585
R87 VTAIL.n92 VTAIL.n91 585
R88 VTAIL.n101 VTAIL.n100 585
R89 VTAIL.n103 VTAIL.n102 585
R90 VTAIL.n88 VTAIL.n87 585
R91 VTAIL.n109 VTAIL.n108 585
R92 VTAIL.n112 VTAIL.n111 585
R93 VTAIL.n110 VTAIL.n84 585
R94 VTAIL.n117 VTAIL.n83 585
R95 VTAIL.n119 VTAIL.n118 585
R96 VTAIL.n121 VTAIL.n120 585
R97 VTAIL.n80 VTAIL.n79 585
R98 VTAIL.n127 VTAIL.n126 585
R99 VTAIL.n129 VTAIL.n128 585
R100 VTAIL.n76 VTAIL.n75 585
R101 VTAIL.n135 VTAIL.n134 585
R102 VTAIL.n137 VTAIL.n136 585
R103 VTAIL.n167 VTAIL.n166 585
R104 VTAIL.n164 VTAIL.n163 585
R105 VTAIL.n173 VTAIL.n172 585
R106 VTAIL.n175 VTAIL.n174 585
R107 VTAIL.n160 VTAIL.n159 585
R108 VTAIL.n181 VTAIL.n180 585
R109 VTAIL.n184 VTAIL.n183 585
R110 VTAIL.n182 VTAIL.n156 585
R111 VTAIL.n189 VTAIL.n155 585
R112 VTAIL.n191 VTAIL.n190 585
R113 VTAIL.n193 VTAIL.n192 585
R114 VTAIL.n152 VTAIL.n151 585
R115 VTAIL.n199 VTAIL.n198 585
R116 VTAIL.n201 VTAIL.n200 585
R117 VTAIL.n148 VTAIL.n147 585
R118 VTAIL.n207 VTAIL.n206 585
R119 VTAIL.n209 VTAIL.n208 585
R120 VTAIL.n493 VTAIL.n492 585
R121 VTAIL.n491 VTAIL.n490 585
R122 VTAIL.n432 VTAIL.n431 585
R123 VTAIL.n485 VTAIL.n484 585
R124 VTAIL.n483 VTAIL.n482 585
R125 VTAIL.n436 VTAIL.n435 585
R126 VTAIL.n477 VTAIL.n476 585
R127 VTAIL.n475 VTAIL.n474 585
R128 VTAIL.n473 VTAIL.n439 585
R129 VTAIL.n443 VTAIL.n440 585
R130 VTAIL.n468 VTAIL.n467 585
R131 VTAIL.n466 VTAIL.n465 585
R132 VTAIL.n445 VTAIL.n444 585
R133 VTAIL.n460 VTAIL.n459 585
R134 VTAIL.n458 VTAIL.n457 585
R135 VTAIL.n449 VTAIL.n448 585
R136 VTAIL.n452 VTAIL.n451 585
R137 VTAIL.n421 VTAIL.n420 585
R138 VTAIL.n419 VTAIL.n418 585
R139 VTAIL.n360 VTAIL.n359 585
R140 VTAIL.n413 VTAIL.n412 585
R141 VTAIL.n411 VTAIL.n410 585
R142 VTAIL.n364 VTAIL.n363 585
R143 VTAIL.n405 VTAIL.n404 585
R144 VTAIL.n403 VTAIL.n402 585
R145 VTAIL.n401 VTAIL.n367 585
R146 VTAIL.n371 VTAIL.n368 585
R147 VTAIL.n396 VTAIL.n395 585
R148 VTAIL.n394 VTAIL.n393 585
R149 VTAIL.n373 VTAIL.n372 585
R150 VTAIL.n388 VTAIL.n387 585
R151 VTAIL.n386 VTAIL.n385 585
R152 VTAIL.n377 VTAIL.n376 585
R153 VTAIL.n380 VTAIL.n379 585
R154 VTAIL.n351 VTAIL.n350 585
R155 VTAIL.n349 VTAIL.n348 585
R156 VTAIL.n290 VTAIL.n289 585
R157 VTAIL.n343 VTAIL.n342 585
R158 VTAIL.n341 VTAIL.n340 585
R159 VTAIL.n294 VTAIL.n293 585
R160 VTAIL.n335 VTAIL.n334 585
R161 VTAIL.n333 VTAIL.n332 585
R162 VTAIL.n331 VTAIL.n297 585
R163 VTAIL.n301 VTAIL.n298 585
R164 VTAIL.n326 VTAIL.n325 585
R165 VTAIL.n324 VTAIL.n323 585
R166 VTAIL.n303 VTAIL.n302 585
R167 VTAIL.n318 VTAIL.n317 585
R168 VTAIL.n316 VTAIL.n315 585
R169 VTAIL.n307 VTAIL.n306 585
R170 VTAIL.n310 VTAIL.n309 585
R171 VTAIL.n279 VTAIL.n278 585
R172 VTAIL.n277 VTAIL.n276 585
R173 VTAIL.n218 VTAIL.n217 585
R174 VTAIL.n271 VTAIL.n270 585
R175 VTAIL.n269 VTAIL.n268 585
R176 VTAIL.n222 VTAIL.n221 585
R177 VTAIL.n263 VTAIL.n262 585
R178 VTAIL.n261 VTAIL.n260 585
R179 VTAIL.n259 VTAIL.n225 585
R180 VTAIL.n229 VTAIL.n226 585
R181 VTAIL.n254 VTAIL.n253 585
R182 VTAIL.n252 VTAIL.n251 585
R183 VTAIL.n231 VTAIL.n230 585
R184 VTAIL.n246 VTAIL.n245 585
R185 VTAIL.n244 VTAIL.n243 585
R186 VTAIL.n235 VTAIL.n234 585
R187 VTAIL.n238 VTAIL.n237 585
R188 VTAIL.t8 VTAIL.n519 329.036
R189 VTAIL.t15 VTAIL.n23 329.036
R190 VTAIL.t5 VTAIL.n93 329.036
R191 VTAIL.t4 VTAIL.n165 329.036
R192 VTAIL.t7 VTAIL.n450 329.036
R193 VTAIL.t2 VTAIL.n378 329.036
R194 VTAIL.t13 VTAIL.n308 329.036
R195 VTAIL.t11 VTAIL.n236 329.036
R196 VTAIL.n520 VTAIL.n517 171.744
R197 VTAIL.n527 VTAIL.n517 171.744
R198 VTAIL.n528 VTAIL.n527 171.744
R199 VTAIL.n528 VTAIL.n513 171.744
R200 VTAIL.n535 VTAIL.n513 171.744
R201 VTAIL.n537 VTAIL.n535 171.744
R202 VTAIL.n537 VTAIL.n536 171.744
R203 VTAIL.n536 VTAIL.n509 171.744
R204 VTAIL.n545 VTAIL.n509 171.744
R205 VTAIL.n546 VTAIL.n545 171.744
R206 VTAIL.n546 VTAIL.n505 171.744
R207 VTAIL.n553 VTAIL.n505 171.744
R208 VTAIL.n554 VTAIL.n553 171.744
R209 VTAIL.n554 VTAIL.n501 171.744
R210 VTAIL.n561 VTAIL.n501 171.744
R211 VTAIL.n562 VTAIL.n561 171.744
R212 VTAIL.n24 VTAIL.n21 171.744
R213 VTAIL.n31 VTAIL.n21 171.744
R214 VTAIL.n32 VTAIL.n31 171.744
R215 VTAIL.n32 VTAIL.n17 171.744
R216 VTAIL.n39 VTAIL.n17 171.744
R217 VTAIL.n41 VTAIL.n39 171.744
R218 VTAIL.n41 VTAIL.n40 171.744
R219 VTAIL.n40 VTAIL.n13 171.744
R220 VTAIL.n49 VTAIL.n13 171.744
R221 VTAIL.n50 VTAIL.n49 171.744
R222 VTAIL.n50 VTAIL.n9 171.744
R223 VTAIL.n57 VTAIL.n9 171.744
R224 VTAIL.n58 VTAIL.n57 171.744
R225 VTAIL.n58 VTAIL.n5 171.744
R226 VTAIL.n65 VTAIL.n5 171.744
R227 VTAIL.n66 VTAIL.n65 171.744
R228 VTAIL.n94 VTAIL.n91 171.744
R229 VTAIL.n101 VTAIL.n91 171.744
R230 VTAIL.n102 VTAIL.n101 171.744
R231 VTAIL.n102 VTAIL.n87 171.744
R232 VTAIL.n109 VTAIL.n87 171.744
R233 VTAIL.n111 VTAIL.n109 171.744
R234 VTAIL.n111 VTAIL.n110 171.744
R235 VTAIL.n110 VTAIL.n83 171.744
R236 VTAIL.n119 VTAIL.n83 171.744
R237 VTAIL.n120 VTAIL.n119 171.744
R238 VTAIL.n120 VTAIL.n79 171.744
R239 VTAIL.n127 VTAIL.n79 171.744
R240 VTAIL.n128 VTAIL.n127 171.744
R241 VTAIL.n128 VTAIL.n75 171.744
R242 VTAIL.n135 VTAIL.n75 171.744
R243 VTAIL.n136 VTAIL.n135 171.744
R244 VTAIL.n166 VTAIL.n163 171.744
R245 VTAIL.n173 VTAIL.n163 171.744
R246 VTAIL.n174 VTAIL.n173 171.744
R247 VTAIL.n174 VTAIL.n159 171.744
R248 VTAIL.n181 VTAIL.n159 171.744
R249 VTAIL.n183 VTAIL.n181 171.744
R250 VTAIL.n183 VTAIL.n182 171.744
R251 VTAIL.n182 VTAIL.n155 171.744
R252 VTAIL.n191 VTAIL.n155 171.744
R253 VTAIL.n192 VTAIL.n191 171.744
R254 VTAIL.n192 VTAIL.n151 171.744
R255 VTAIL.n199 VTAIL.n151 171.744
R256 VTAIL.n200 VTAIL.n199 171.744
R257 VTAIL.n200 VTAIL.n147 171.744
R258 VTAIL.n207 VTAIL.n147 171.744
R259 VTAIL.n208 VTAIL.n207 171.744
R260 VTAIL.n492 VTAIL.n491 171.744
R261 VTAIL.n491 VTAIL.n431 171.744
R262 VTAIL.n484 VTAIL.n431 171.744
R263 VTAIL.n484 VTAIL.n483 171.744
R264 VTAIL.n483 VTAIL.n435 171.744
R265 VTAIL.n476 VTAIL.n435 171.744
R266 VTAIL.n476 VTAIL.n475 171.744
R267 VTAIL.n475 VTAIL.n439 171.744
R268 VTAIL.n443 VTAIL.n439 171.744
R269 VTAIL.n467 VTAIL.n443 171.744
R270 VTAIL.n467 VTAIL.n466 171.744
R271 VTAIL.n466 VTAIL.n444 171.744
R272 VTAIL.n459 VTAIL.n444 171.744
R273 VTAIL.n459 VTAIL.n458 171.744
R274 VTAIL.n458 VTAIL.n448 171.744
R275 VTAIL.n451 VTAIL.n448 171.744
R276 VTAIL.n420 VTAIL.n419 171.744
R277 VTAIL.n419 VTAIL.n359 171.744
R278 VTAIL.n412 VTAIL.n359 171.744
R279 VTAIL.n412 VTAIL.n411 171.744
R280 VTAIL.n411 VTAIL.n363 171.744
R281 VTAIL.n404 VTAIL.n363 171.744
R282 VTAIL.n404 VTAIL.n403 171.744
R283 VTAIL.n403 VTAIL.n367 171.744
R284 VTAIL.n371 VTAIL.n367 171.744
R285 VTAIL.n395 VTAIL.n371 171.744
R286 VTAIL.n395 VTAIL.n394 171.744
R287 VTAIL.n394 VTAIL.n372 171.744
R288 VTAIL.n387 VTAIL.n372 171.744
R289 VTAIL.n387 VTAIL.n386 171.744
R290 VTAIL.n386 VTAIL.n376 171.744
R291 VTAIL.n379 VTAIL.n376 171.744
R292 VTAIL.n350 VTAIL.n349 171.744
R293 VTAIL.n349 VTAIL.n289 171.744
R294 VTAIL.n342 VTAIL.n289 171.744
R295 VTAIL.n342 VTAIL.n341 171.744
R296 VTAIL.n341 VTAIL.n293 171.744
R297 VTAIL.n334 VTAIL.n293 171.744
R298 VTAIL.n334 VTAIL.n333 171.744
R299 VTAIL.n333 VTAIL.n297 171.744
R300 VTAIL.n301 VTAIL.n297 171.744
R301 VTAIL.n325 VTAIL.n301 171.744
R302 VTAIL.n325 VTAIL.n324 171.744
R303 VTAIL.n324 VTAIL.n302 171.744
R304 VTAIL.n317 VTAIL.n302 171.744
R305 VTAIL.n317 VTAIL.n316 171.744
R306 VTAIL.n316 VTAIL.n306 171.744
R307 VTAIL.n309 VTAIL.n306 171.744
R308 VTAIL.n278 VTAIL.n277 171.744
R309 VTAIL.n277 VTAIL.n217 171.744
R310 VTAIL.n270 VTAIL.n217 171.744
R311 VTAIL.n270 VTAIL.n269 171.744
R312 VTAIL.n269 VTAIL.n221 171.744
R313 VTAIL.n262 VTAIL.n221 171.744
R314 VTAIL.n262 VTAIL.n261 171.744
R315 VTAIL.n261 VTAIL.n225 171.744
R316 VTAIL.n229 VTAIL.n225 171.744
R317 VTAIL.n253 VTAIL.n229 171.744
R318 VTAIL.n253 VTAIL.n252 171.744
R319 VTAIL.n252 VTAIL.n230 171.744
R320 VTAIL.n245 VTAIL.n230 171.744
R321 VTAIL.n245 VTAIL.n244 171.744
R322 VTAIL.n244 VTAIL.n234 171.744
R323 VTAIL.n237 VTAIL.n234 171.744
R324 VTAIL.n520 VTAIL.t8 85.8723
R325 VTAIL.n24 VTAIL.t15 85.8723
R326 VTAIL.n94 VTAIL.t5 85.8723
R327 VTAIL.n166 VTAIL.t4 85.8723
R328 VTAIL.n451 VTAIL.t7 85.8723
R329 VTAIL.n379 VTAIL.t2 85.8723
R330 VTAIL.n309 VTAIL.t13 85.8723
R331 VTAIL.n237 VTAIL.t11 85.8723
R332 VTAIL.n1 VTAIL.n0 55.7508
R333 VTAIL.n143 VTAIL.n142 55.7508
R334 VTAIL.n427 VTAIL.n426 55.7508
R335 VTAIL.n285 VTAIL.n284 55.7508
R336 VTAIL.n567 VTAIL.n566 31.6035
R337 VTAIL.n71 VTAIL.n70 31.6035
R338 VTAIL.n141 VTAIL.n140 31.6035
R339 VTAIL.n213 VTAIL.n212 31.6035
R340 VTAIL.n497 VTAIL.n496 31.6035
R341 VTAIL.n425 VTAIL.n424 31.6035
R342 VTAIL.n355 VTAIL.n354 31.6035
R343 VTAIL.n283 VTAIL.n282 31.6035
R344 VTAIL.n567 VTAIL.n497 24.1169
R345 VTAIL.n283 VTAIL.n213 24.1169
R346 VTAIL.n544 VTAIL.n543 13.1884
R347 VTAIL.n48 VTAIL.n47 13.1884
R348 VTAIL.n118 VTAIL.n117 13.1884
R349 VTAIL.n190 VTAIL.n189 13.1884
R350 VTAIL.n474 VTAIL.n473 13.1884
R351 VTAIL.n402 VTAIL.n401 13.1884
R352 VTAIL.n332 VTAIL.n331 13.1884
R353 VTAIL.n260 VTAIL.n259 13.1884
R354 VTAIL.n542 VTAIL.n510 12.8005
R355 VTAIL.n547 VTAIL.n508 12.8005
R356 VTAIL.n46 VTAIL.n14 12.8005
R357 VTAIL.n51 VTAIL.n12 12.8005
R358 VTAIL.n116 VTAIL.n84 12.8005
R359 VTAIL.n121 VTAIL.n82 12.8005
R360 VTAIL.n188 VTAIL.n156 12.8005
R361 VTAIL.n193 VTAIL.n154 12.8005
R362 VTAIL.n477 VTAIL.n438 12.8005
R363 VTAIL.n472 VTAIL.n440 12.8005
R364 VTAIL.n405 VTAIL.n366 12.8005
R365 VTAIL.n400 VTAIL.n368 12.8005
R366 VTAIL.n335 VTAIL.n296 12.8005
R367 VTAIL.n330 VTAIL.n298 12.8005
R368 VTAIL.n263 VTAIL.n224 12.8005
R369 VTAIL.n258 VTAIL.n226 12.8005
R370 VTAIL.n539 VTAIL.n538 12.0247
R371 VTAIL.n548 VTAIL.n506 12.0247
R372 VTAIL.n43 VTAIL.n42 12.0247
R373 VTAIL.n52 VTAIL.n10 12.0247
R374 VTAIL.n113 VTAIL.n112 12.0247
R375 VTAIL.n122 VTAIL.n80 12.0247
R376 VTAIL.n185 VTAIL.n184 12.0247
R377 VTAIL.n194 VTAIL.n152 12.0247
R378 VTAIL.n478 VTAIL.n436 12.0247
R379 VTAIL.n469 VTAIL.n468 12.0247
R380 VTAIL.n406 VTAIL.n364 12.0247
R381 VTAIL.n397 VTAIL.n396 12.0247
R382 VTAIL.n336 VTAIL.n294 12.0247
R383 VTAIL.n327 VTAIL.n326 12.0247
R384 VTAIL.n264 VTAIL.n222 12.0247
R385 VTAIL.n255 VTAIL.n254 12.0247
R386 VTAIL.n534 VTAIL.n512 11.249
R387 VTAIL.n552 VTAIL.n551 11.249
R388 VTAIL.n38 VTAIL.n16 11.249
R389 VTAIL.n56 VTAIL.n55 11.249
R390 VTAIL.n108 VTAIL.n86 11.249
R391 VTAIL.n126 VTAIL.n125 11.249
R392 VTAIL.n180 VTAIL.n158 11.249
R393 VTAIL.n198 VTAIL.n197 11.249
R394 VTAIL.n482 VTAIL.n481 11.249
R395 VTAIL.n465 VTAIL.n442 11.249
R396 VTAIL.n410 VTAIL.n409 11.249
R397 VTAIL.n393 VTAIL.n370 11.249
R398 VTAIL.n340 VTAIL.n339 11.249
R399 VTAIL.n323 VTAIL.n300 11.249
R400 VTAIL.n268 VTAIL.n267 11.249
R401 VTAIL.n251 VTAIL.n228 11.249
R402 VTAIL.n521 VTAIL.n519 10.7239
R403 VTAIL.n25 VTAIL.n23 10.7239
R404 VTAIL.n95 VTAIL.n93 10.7239
R405 VTAIL.n167 VTAIL.n165 10.7239
R406 VTAIL.n452 VTAIL.n450 10.7239
R407 VTAIL.n380 VTAIL.n378 10.7239
R408 VTAIL.n310 VTAIL.n308 10.7239
R409 VTAIL.n238 VTAIL.n236 10.7239
R410 VTAIL.n533 VTAIL.n514 10.4732
R411 VTAIL.n555 VTAIL.n504 10.4732
R412 VTAIL.n37 VTAIL.n18 10.4732
R413 VTAIL.n59 VTAIL.n8 10.4732
R414 VTAIL.n107 VTAIL.n88 10.4732
R415 VTAIL.n129 VTAIL.n78 10.4732
R416 VTAIL.n179 VTAIL.n160 10.4732
R417 VTAIL.n201 VTAIL.n150 10.4732
R418 VTAIL.n485 VTAIL.n434 10.4732
R419 VTAIL.n464 VTAIL.n445 10.4732
R420 VTAIL.n413 VTAIL.n362 10.4732
R421 VTAIL.n392 VTAIL.n373 10.4732
R422 VTAIL.n343 VTAIL.n292 10.4732
R423 VTAIL.n322 VTAIL.n303 10.4732
R424 VTAIL.n271 VTAIL.n220 10.4732
R425 VTAIL.n250 VTAIL.n231 10.4732
R426 VTAIL.n530 VTAIL.n529 9.69747
R427 VTAIL.n556 VTAIL.n502 9.69747
R428 VTAIL.n34 VTAIL.n33 9.69747
R429 VTAIL.n60 VTAIL.n6 9.69747
R430 VTAIL.n104 VTAIL.n103 9.69747
R431 VTAIL.n130 VTAIL.n76 9.69747
R432 VTAIL.n176 VTAIL.n175 9.69747
R433 VTAIL.n202 VTAIL.n148 9.69747
R434 VTAIL.n486 VTAIL.n432 9.69747
R435 VTAIL.n461 VTAIL.n460 9.69747
R436 VTAIL.n414 VTAIL.n360 9.69747
R437 VTAIL.n389 VTAIL.n388 9.69747
R438 VTAIL.n344 VTAIL.n290 9.69747
R439 VTAIL.n319 VTAIL.n318 9.69747
R440 VTAIL.n272 VTAIL.n218 9.69747
R441 VTAIL.n247 VTAIL.n246 9.69747
R442 VTAIL.n566 VTAIL.n565 9.45567
R443 VTAIL.n70 VTAIL.n69 9.45567
R444 VTAIL.n140 VTAIL.n139 9.45567
R445 VTAIL.n212 VTAIL.n211 9.45567
R446 VTAIL.n496 VTAIL.n495 9.45567
R447 VTAIL.n424 VTAIL.n423 9.45567
R448 VTAIL.n354 VTAIL.n353 9.45567
R449 VTAIL.n282 VTAIL.n281 9.45567
R450 VTAIL.n500 VTAIL.n499 9.3005
R451 VTAIL.n559 VTAIL.n558 9.3005
R452 VTAIL.n557 VTAIL.n556 9.3005
R453 VTAIL.n504 VTAIL.n503 9.3005
R454 VTAIL.n551 VTAIL.n550 9.3005
R455 VTAIL.n549 VTAIL.n548 9.3005
R456 VTAIL.n508 VTAIL.n507 9.3005
R457 VTAIL.n523 VTAIL.n522 9.3005
R458 VTAIL.n525 VTAIL.n524 9.3005
R459 VTAIL.n516 VTAIL.n515 9.3005
R460 VTAIL.n531 VTAIL.n530 9.3005
R461 VTAIL.n533 VTAIL.n532 9.3005
R462 VTAIL.n512 VTAIL.n511 9.3005
R463 VTAIL.n540 VTAIL.n539 9.3005
R464 VTAIL.n542 VTAIL.n541 9.3005
R465 VTAIL.n565 VTAIL.n564 9.3005
R466 VTAIL.n4 VTAIL.n3 9.3005
R467 VTAIL.n63 VTAIL.n62 9.3005
R468 VTAIL.n61 VTAIL.n60 9.3005
R469 VTAIL.n8 VTAIL.n7 9.3005
R470 VTAIL.n55 VTAIL.n54 9.3005
R471 VTAIL.n53 VTAIL.n52 9.3005
R472 VTAIL.n12 VTAIL.n11 9.3005
R473 VTAIL.n27 VTAIL.n26 9.3005
R474 VTAIL.n29 VTAIL.n28 9.3005
R475 VTAIL.n20 VTAIL.n19 9.3005
R476 VTAIL.n35 VTAIL.n34 9.3005
R477 VTAIL.n37 VTAIL.n36 9.3005
R478 VTAIL.n16 VTAIL.n15 9.3005
R479 VTAIL.n44 VTAIL.n43 9.3005
R480 VTAIL.n46 VTAIL.n45 9.3005
R481 VTAIL.n69 VTAIL.n68 9.3005
R482 VTAIL.n74 VTAIL.n73 9.3005
R483 VTAIL.n133 VTAIL.n132 9.3005
R484 VTAIL.n131 VTAIL.n130 9.3005
R485 VTAIL.n78 VTAIL.n77 9.3005
R486 VTAIL.n125 VTAIL.n124 9.3005
R487 VTAIL.n123 VTAIL.n122 9.3005
R488 VTAIL.n82 VTAIL.n81 9.3005
R489 VTAIL.n97 VTAIL.n96 9.3005
R490 VTAIL.n99 VTAIL.n98 9.3005
R491 VTAIL.n90 VTAIL.n89 9.3005
R492 VTAIL.n105 VTAIL.n104 9.3005
R493 VTAIL.n107 VTAIL.n106 9.3005
R494 VTAIL.n86 VTAIL.n85 9.3005
R495 VTAIL.n114 VTAIL.n113 9.3005
R496 VTAIL.n116 VTAIL.n115 9.3005
R497 VTAIL.n139 VTAIL.n138 9.3005
R498 VTAIL.n146 VTAIL.n145 9.3005
R499 VTAIL.n205 VTAIL.n204 9.3005
R500 VTAIL.n203 VTAIL.n202 9.3005
R501 VTAIL.n150 VTAIL.n149 9.3005
R502 VTAIL.n197 VTAIL.n196 9.3005
R503 VTAIL.n195 VTAIL.n194 9.3005
R504 VTAIL.n154 VTAIL.n153 9.3005
R505 VTAIL.n169 VTAIL.n168 9.3005
R506 VTAIL.n171 VTAIL.n170 9.3005
R507 VTAIL.n162 VTAIL.n161 9.3005
R508 VTAIL.n177 VTAIL.n176 9.3005
R509 VTAIL.n179 VTAIL.n178 9.3005
R510 VTAIL.n158 VTAIL.n157 9.3005
R511 VTAIL.n186 VTAIL.n185 9.3005
R512 VTAIL.n188 VTAIL.n187 9.3005
R513 VTAIL.n211 VTAIL.n210 9.3005
R514 VTAIL.n454 VTAIL.n453 9.3005
R515 VTAIL.n456 VTAIL.n455 9.3005
R516 VTAIL.n447 VTAIL.n446 9.3005
R517 VTAIL.n462 VTAIL.n461 9.3005
R518 VTAIL.n464 VTAIL.n463 9.3005
R519 VTAIL.n442 VTAIL.n441 9.3005
R520 VTAIL.n470 VTAIL.n469 9.3005
R521 VTAIL.n472 VTAIL.n471 9.3005
R522 VTAIL.n495 VTAIL.n494 9.3005
R523 VTAIL.n430 VTAIL.n429 9.3005
R524 VTAIL.n489 VTAIL.n488 9.3005
R525 VTAIL.n487 VTAIL.n486 9.3005
R526 VTAIL.n434 VTAIL.n433 9.3005
R527 VTAIL.n481 VTAIL.n480 9.3005
R528 VTAIL.n479 VTAIL.n478 9.3005
R529 VTAIL.n438 VTAIL.n437 9.3005
R530 VTAIL.n382 VTAIL.n381 9.3005
R531 VTAIL.n384 VTAIL.n383 9.3005
R532 VTAIL.n375 VTAIL.n374 9.3005
R533 VTAIL.n390 VTAIL.n389 9.3005
R534 VTAIL.n392 VTAIL.n391 9.3005
R535 VTAIL.n370 VTAIL.n369 9.3005
R536 VTAIL.n398 VTAIL.n397 9.3005
R537 VTAIL.n400 VTAIL.n399 9.3005
R538 VTAIL.n423 VTAIL.n422 9.3005
R539 VTAIL.n358 VTAIL.n357 9.3005
R540 VTAIL.n417 VTAIL.n416 9.3005
R541 VTAIL.n415 VTAIL.n414 9.3005
R542 VTAIL.n362 VTAIL.n361 9.3005
R543 VTAIL.n409 VTAIL.n408 9.3005
R544 VTAIL.n407 VTAIL.n406 9.3005
R545 VTAIL.n366 VTAIL.n365 9.3005
R546 VTAIL.n312 VTAIL.n311 9.3005
R547 VTAIL.n314 VTAIL.n313 9.3005
R548 VTAIL.n305 VTAIL.n304 9.3005
R549 VTAIL.n320 VTAIL.n319 9.3005
R550 VTAIL.n322 VTAIL.n321 9.3005
R551 VTAIL.n300 VTAIL.n299 9.3005
R552 VTAIL.n328 VTAIL.n327 9.3005
R553 VTAIL.n330 VTAIL.n329 9.3005
R554 VTAIL.n353 VTAIL.n352 9.3005
R555 VTAIL.n288 VTAIL.n287 9.3005
R556 VTAIL.n347 VTAIL.n346 9.3005
R557 VTAIL.n345 VTAIL.n344 9.3005
R558 VTAIL.n292 VTAIL.n291 9.3005
R559 VTAIL.n339 VTAIL.n338 9.3005
R560 VTAIL.n337 VTAIL.n336 9.3005
R561 VTAIL.n296 VTAIL.n295 9.3005
R562 VTAIL.n240 VTAIL.n239 9.3005
R563 VTAIL.n242 VTAIL.n241 9.3005
R564 VTAIL.n233 VTAIL.n232 9.3005
R565 VTAIL.n248 VTAIL.n247 9.3005
R566 VTAIL.n250 VTAIL.n249 9.3005
R567 VTAIL.n228 VTAIL.n227 9.3005
R568 VTAIL.n256 VTAIL.n255 9.3005
R569 VTAIL.n258 VTAIL.n257 9.3005
R570 VTAIL.n281 VTAIL.n280 9.3005
R571 VTAIL.n216 VTAIL.n215 9.3005
R572 VTAIL.n275 VTAIL.n274 9.3005
R573 VTAIL.n273 VTAIL.n272 9.3005
R574 VTAIL.n220 VTAIL.n219 9.3005
R575 VTAIL.n267 VTAIL.n266 9.3005
R576 VTAIL.n265 VTAIL.n264 9.3005
R577 VTAIL.n224 VTAIL.n223 9.3005
R578 VTAIL.n526 VTAIL.n516 8.92171
R579 VTAIL.n560 VTAIL.n559 8.92171
R580 VTAIL.n30 VTAIL.n20 8.92171
R581 VTAIL.n64 VTAIL.n63 8.92171
R582 VTAIL.n100 VTAIL.n90 8.92171
R583 VTAIL.n134 VTAIL.n133 8.92171
R584 VTAIL.n172 VTAIL.n162 8.92171
R585 VTAIL.n206 VTAIL.n205 8.92171
R586 VTAIL.n490 VTAIL.n489 8.92171
R587 VTAIL.n457 VTAIL.n447 8.92171
R588 VTAIL.n418 VTAIL.n417 8.92171
R589 VTAIL.n385 VTAIL.n375 8.92171
R590 VTAIL.n348 VTAIL.n347 8.92171
R591 VTAIL.n315 VTAIL.n305 8.92171
R592 VTAIL.n276 VTAIL.n275 8.92171
R593 VTAIL.n243 VTAIL.n233 8.92171
R594 VTAIL.n525 VTAIL.n518 8.14595
R595 VTAIL.n563 VTAIL.n500 8.14595
R596 VTAIL.n29 VTAIL.n22 8.14595
R597 VTAIL.n67 VTAIL.n4 8.14595
R598 VTAIL.n99 VTAIL.n92 8.14595
R599 VTAIL.n137 VTAIL.n74 8.14595
R600 VTAIL.n171 VTAIL.n164 8.14595
R601 VTAIL.n209 VTAIL.n146 8.14595
R602 VTAIL.n493 VTAIL.n430 8.14595
R603 VTAIL.n456 VTAIL.n449 8.14595
R604 VTAIL.n421 VTAIL.n358 8.14595
R605 VTAIL.n384 VTAIL.n377 8.14595
R606 VTAIL.n351 VTAIL.n288 8.14595
R607 VTAIL.n314 VTAIL.n307 8.14595
R608 VTAIL.n279 VTAIL.n216 8.14595
R609 VTAIL.n242 VTAIL.n235 8.14595
R610 VTAIL.n522 VTAIL.n521 7.3702
R611 VTAIL.n564 VTAIL.n498 7.3702
R612 VTAIL.n26 VTAIL.n25 7.3702
R613 VTAIL.n68 VTAIL.n2 7.3702
R614 VTAIL.n96 VTAIL.n95 7.3702
R615 VTAIL.n138 VTAIL.n72 7.3702
R616 VTAIL.n168 VTAIL.n167 7.3702
R617 VTAIL.n210 VTAIL.n144 7.3702
R618 VTAIL.n494 VTAIL.n428 7.3702
R619 VTAIL.n453 VTAIL.n452 7.3702
R620 VTAIL.n422 VTAIL.n356 7.3702
R621 VTAIL.n381 VTAIL.n380 7.3702
R622 VTAIL.n352 VTAIL.n286 7.3702
R623 VTAIL.n311 VTAIL.n310 7.3702
R624 VTAIL.n280 VTAIL.n214 7.3702
R625 VTAIL.n239 VTAIL.n238 7.3702
R626 VTAIL.n566 VTAIL.n498 6.59444
R627 VTAIL.n70 VTAIL.n2 6.59444
R628 VTAIL.n140 VTAIL.n72 6.59444
R629 VTAIL.n212 VTAIL.n144 6.59444
R630 VTAIL.n496 VTAIL.n428 6.59444
R631 VTAIL.n424 VTAIL.n356 6.59444
R632 VTAIL.n354 VTAIL.n286 6.59444
R633 VTAIL.n282 VTAIL.n214 6.59444
R634 VTAIL.n522 VTAIL.n518 5.81868
R635 VTAIL.n564 VTAIL.n563 5.81868
R636 VTAIL.n26 VTAIL.n22 5.81868
R637 VTAIL.n68 VTAIL.n67 5.81868
R638 VTAIL.n96 VTAIL.n92 5.81868
R639 VTAIL.n138 VTAIL.n137 5.81868
R640 VTAIL.n168 VTAIL.n164 5.81868
R641 VTAIL.n210 VTAIL.n209 5.81868
R642 VTAIL.n494 VTAIL.n493 5.81868
R643 VTAIL.n453 VTAIL.n449 5.81868
R644 VTAIL.n422 VTAIL.n421 5.81868
R645 VTAIL.n381 VTAIL.n377 5.81868
R646 VTAIL.n352 VTAIL.n351 5.81868
R647 VTAIL.n311 VTAIL.n307 5.81868
R648 VTAIL.n280 VTAIL.n279 5.81868
R649 VTAIL.n239 VTAIL.n235 5.81868
R650 VTAIL.n526 VTAIL.n525 5.04292
R651 VTAIL.n560 VTAIL.n500 5.04292
R652 VTAIL.n30 VTAIL.n29 5.04292
R653 VTAIL.n64 VTAIL.n4 5.04292
R654 VTAIL.n100 VTAIL.n99 5.04292
R655 VTAIL.n134 VTAIL.n74 5.04292
R656 VTAIL.n172 VTAIL.n171 5.04292
R657 VTAIL.n206 VTAIL.n146 5.04292
R658 VTAIL.n490 VTAIL.n430 5.04292
R659 VTAIL.n457 VTAIL.n456 5.04292
R660 VTAIL.n418 VTAIL.n358 5.04292
R661 VTAIL.n385 VTAIL.n384 5.04292
R662 VTAIL.n348 VTAIL.n288 5.04292
R663 VTAIL.n315 VTAIL.n314 5.04292
R664 VTAIL.n276 VTAIL.n216 5.04292
R665 VTAIL.n243 VTAIL.n242 5.04292
R666 VTAIL.n529 VTAIL.n516 4.26717
R667 VTAIL.n559 VTAIL.n502 4.26717
R668 VTAIL.n33 VTAIL.n20 4.26717
R669 VTAIL.n63 VTAIL.n6 4.26717
R670 VTAIL.n103 VTAIL.n90 4.26717
R671 VTAIL.n133 VTAIL.n76 4.26717
R672 VTAIL.n175 VTAIL.n162 4.26717
R673 VTAIL.n205 VTAIL.n148 4.26717
R674 VTAIL.n489 VTAIL.n432 4.26717
R675 VTAIL.n460 VTAIL.n447 4.26717
R676 VTAIL.n417 VTAIL.n360 4.26717
R677 VTAIL.n388 VTAIL.n375 4.26717
R678 VTAIL.n347 VTAIL.n290 4.26717
R679 VTAIL.n318 VTAIL.n305 4.26717
R680 VTAIL.n275 VTAIL.n218 4.26717
R681 VTAIL.n246 VTAIL.n233 4.26717
R682 VTAIL.n530 VTAIL.n514 3.49141
R683 VTAIL.n556 VTAIL.n555 3.49141
R684 VTAIL.n34 VTAIL.n18 3.49141
R685 VTAIL.n60 VTAIL.n59 3.49141
R686 VTAIL.n104 VTAIL.n88 3.49141
R687 VTAIL.n130 VTAIL.n129 3.49141
R688 VTAIL.n176 VTAIL.n160 3.49141
R689 VTAIL.n202 VTAIL.n201 3.49141
R690 VTAIL.n486 VTAIL.n485 3.49141
R691 VTAIL.n461 VTAIL.n445 3.49141
R692 VTAIL.n414 VTAIL.n413 3.49141
R693 VTAIL.n389 VTAIL.n373 3.49141
R694 VTAIL.n344 VTAIL.n343 3.49141
R695 VTAIL.n319 VTAIL.n303 3.49141
R696 VTAIL.n272 VTAIL.n271 3.49141
R697 VTAIL.n247 VTAIL.n231 3.49141
R698 VTAIL.n534 VTAIL.n533 2.71565
R699 VTAIL.n552 VTAIL.n504 2.71565
R700 VTAIL.n38 VTAIL.n37 2.71565
R701 VTAIL.n56 VTAIL.n8 2.71565
R702 VTAIL.n108 VTAIL.n107 2.71565
R703 VTAIL.n126 VTAIL.n78 2.71565
R704 VTAIL.n180 VTAIL.n179 2.71565
R705 VTAIL.n198 VTAIL.n150 2.71565
R706 VTAIL.n482 VTAIL.n434 2.71565
R707 VTAIL.n465 VTAIL.n464 2.71565
R708 VTAIL.n410 VTAIL.n362 2.71565
R709 VTAIL.n393 VTAIL.n392 2.71565
R710 VTAIL.n340 VTAIL.n292 2.71565
R711 VTAIL.n323 VTAIL.n322 2.71565
R712 VTAIL.n268 VTAIL.n220 2.71565
R713 VTAIL.n251 VTAIL.n250 2.71565
R714 VTAIL.n0 VTAIL.t14 2.53797
R715 VTAIL.n0 VTAIL.t9 2.53797
R716 VTAIL.n142 VTAIL.t1 2.53797
R717 VTAIL.n142 VTAIL.t3 2.53797
R718 VTAIL.n426 VTAIL.t0 2.53797
R719 VTAIL.n426 VTAIL.t6 2.53797
R720 VTAIL.n284 VTAIL.t12 2.53797
R721 VTAIL.n284 VTAIL.t10 2.53797
R722 VTAIL.n523 VTAIL.n519 2.41282
R723 VTAIL.n27 VTAIL.n23 2.41282
R724 VTAIL.n97 VTAIL.n93 2.41282
R725 VTAIL.n169 VTAIL.n165 2.41282
R726 VTAIL.n454 VTAIL.n450 2.41282
R727 VTAIL.n382 VTAIL.n378 2.41282
R728 VTAIL.n312 VTAIL.n308 2.41282
R729 VTAIL.n240 VTAIL.n236 2.41282
R730 VTAIL.n538 VTAIL.n512 1.93989
R731 VTAIL.n551 VTAIL.n506 1.93989
R732 VTAIL.n42 VTAIL.n16 1.93989
R733 VTAIL.n55 VTAIL.n10 1.93989
R734 VTAIL.n112 VTAIL.n86 1.93989
R735 VTAIL.n125 VTAIL.n80 1.93989
R736 VTAIL.n184 VTAIL.n158 1.93989
R737 VTAIL.n197 VTAIL.n152 1.93989
R738 VTAIL.n481 VTAIL.n436 1.93989
R739 VTAIL.n468 VTAIL.n442 1.93989
R740 VTAIL.n409 VTAIL.n364 1.93989
R741 VTAIL.n396 VTAIL.n370 1.93989
R742 VTAIL.n339 VTAIL.n294 1.93989
R743 VTAIL.n326 VTAIL.n300 1.93989
R744 VTAIL.n267 VTAIL.n222 1.93989
R745 VTAIL.n254 VTAIL.n228 1.93989
R746 VTAIL.n539 VTAIL.n510 1.16414
R747 VTAIL.n548 VTAIL.n547 1.16414
R748 VTAIL.n43 VTAIL.n14 1.16414
R749 VTAIL.n52 VTAIL.n51 1.16414
R750 VTAIL.n113 VTAIL.n84 1.16414
R751 VTAIL.n122 VTAIL.n121 1.16414
R752 VTAIL.n185 VTAIL.n156 1.16414
R753 VTAIL.n194 VTAIL.n193 1.16414
R754 VTAIL.n478 VTAIL.n477 1.16414
R755 VTAIL.n469 VTAIL.n440 1.16414
R756 VTAIL.n406 VTAIL.n405 1.16414
R757 VTAIL.n397 VTAIL.n368 1.16414
R758 VTAIL.n336 VTAIL.n335 1.16414
R759 VTAIL.n327 VTAIL.n298 1.16414
R760 VTAIL.n264 VTAIL.n263 1.16414
R761 VTAIL.n255 VTAIL.n226 1.16414
R762 VTAIL.n285 VTAIL.n283 0.707397
R763 VTAIL.n355 VTAIL.n285 0.707397
R764 VTAIL.n427 VTAIL.n425 0.707397
R765 VTAIL.n497 VTAIL.n427 0.707397
R766 VTAIL.n213 VTAIL.n143 0.707397
R767 VTAIL.n143 VTAIL.n141 0.707397
R768 VTAIL.n71 VTAIL.n1 0.707397
R769 VTAIL VTAIL.n567 0.649207
R770 VTAIL.n425 VTAIL.n355 0.470328
R771 VTAIL.n141 VTAIL.n71 0.470328
R772 VTAIL.n543 VTAIL.n542 0.388379
R773 VTAIL.n544 VTAIL.n508 0.388379
R774 VTAIL.n47 VTAIL.n46 0.388379
R775 VTAIL.n48 VTAIL.n12 0.388379
R776 VTAIL.n117 VTAIL.n116 0.388379
R777 VTAIL.n118 VTAIL.n82 0.388379
R778 VTAIL.n189 VTAIL.n188 0.388379
R779 VTAIL.n190 VTAIL.n154 0.388379
R780 VTAIL.n474 VTAIL.n438 0.388379
R781 VTAIL.n473 VTAIL.n472 0.388379
R782 VTAIL.n402 VTAIL.n366 0.388379
R783 VTAIL.n401 VTAIL.n400 0.388379
R784 VTAIL.n332 VTAIL.n296 0.388379
R785 VTAIL.n331 VTAIL.n330 0.388379
R786 VTAIL.n260 VTAIL.n224 0.388379
R787 VTAIL.n259 VTAIL.n258 0.388379
R788 VTAIL.n524 VTAIL.n523 0.155672
R789 VTAIL.n524 VTAIL.n515 0.155672
R790 VTAIL.n531 VTAIL.n515 0.155672
R791 VTAIL.n532 VTAIL.n531 0.155672
R792 VTAIL.n532 VTAIL.n511 0.155672
R793 VTAIL.n540 VTAIL.n511 0.155672
R794 VTAIL.n541 VTAIL.n540 0.155672
R795 VTAIL.n541 VTAIL.n507 0.155672
R796 VTAIL.n549 VTAIL.n507 0.155672
R797 VTAIL.n550 VTAIL.n549 0.155672
R798 VTAIL.n550 VTAIL.n503 0.155672
R799 VTAIL.n557 VTAIL.n503 0.155672
R800 VTAIL.n558 VTAIL.n557 0.155672
R801 VTAIL.n558 VTAIL.n499 0.155672
R802 VTAIL.n565 VTAIL.n499 0.155672
R803 VTAIL.n28 VTAIL.n27 0.155672
R804 VTAIL.n28 VTAIL.n19 0.155672
R805 VTAIL.n35 VTAIL.n19 0.155672
R806 VTAIL.n36 VTAIL.n35 0.155672
R807 VTAIL.n36 VTAIL.n15 0.155672
R808 VTAIL.n44 VTAIL.n15 0.155672
R809 VTAIL.n45 VTAIL.n44 0.155672
R810 VTAIL.n45 VTAIL.n11 0.155672
R811 VTAIL.n53 VTAIL.n11 0.155672
R812 VTAIL.n54 VTAIL.n53 0.155672
R813 VTAIL.n54 VTAIL.n7 0.155672
R814 VTAIL.n61 VTAIL.n7 0.155672
R815 VTAIL.n62 VTAIL.n61 0.155672
R816 VTAIL.n62 VTAIL.n3 0.155672
R817 VTAIL.n69 VTAIL.n3 0.155672
R818 VTAIL.n98 VTAIL.n97 0.155672
R819 VTAIL.n98 VTAIL.n89 0.155672
R820 VTAIL.n105 VTAIL.n89 0.155672
R821 VTAIL.n106 VTAIL.n105 0.155672
R822 VTAIL.n106 VTAIL.n85 0.155672
R823 VTAIL.n114 VTAIL.n85 0.155672
R824 VTAIL.n115 VTAIL.n114 0.155672
R825 VTAIL.n115 VTAIL.n81 0.155672
R826 VTAIL.n123 VTAIL.n81 0.155672
R827 VTAIL.n124 VTAIL.n123 0.155672
R828 VTAIL.n124 VTAIL.n77 0.155672
R829 VTAIL.n131 VTAIL.n77 0.155672
R830 VTAIL.n132 VTAIL.n131 0.155672
R831 VTAIL.n132 VTAIL.n73 0.155672
R832 VTAIL.n139 VTAIL.n73 0.155672
R833 VTAIL.n170 VTAIL.n169 0.155672
R834 VTAIL.n170 VTAIL.n161 0.155672
R835 VTAIL.n177 VTAIL.n161 0.155672
R836 VTAIL.n178 VTAIL.n177 0.155672
R837 VTAIL.n178 VTAIL.n157 0.155672
R838 VTAIL.n186 VTAIL.n157 0.155672
R839 VTAIL.n187 VTAIL.n186 0.155672
R840 VTAIL.n187 VTAIL.n153 0.155672
R841 VTAIL.n195 VTAIL.n153 0.155672
R842 VTAIL.n196 VTAIL.n195 0.155672
R843 VTAIL.n196 VTAIL.n149 0.155672
R844 VTAIL.n203 VTAIL.n149 0.155672
R845 VTAIL.n204 VTAIL.n203 0.155672
R846 VTAIL.n204 VTAIL.n145 0.155672
R847 VTAIL.n211 VTAIL.n145 0.155672
R848 VTAIL.n495 VTAIL.n429 0.155672
R849 VTAIL.n488 VTAIL.n429 0.155672
R850 VTAIL.n488 VTAIL.n487 0.155672
R851 VTAIL.n487 VTAIL.n433 0.155672
R852 VTAIL.n480 VTAIL.n433 0.155672
R853 VTAIL.n480 VTAIL.n479 0.155672
R854 VTAIL.n479 VTAIL.n437 0.155672
R855 VTAIL.n471 VTAIL.n437 0.155672
R856 VTAIL.n471 VTAIL.n470 0.155672
R857 VTAIL.n470 VTAIL.n441 0.155672
R858 VTAIL.n463 VTAIL.n441 0.155672
R859 VTAIL.n463 VTAIL.n462 0.155672
R860 VTAIL.n462 VTAIL.n446 0.155672
R861 VTAIL.n455 VTAIL.n446 0.155672
R862 VTAIL.n455 VTAIL.n454 0.155672
R863 VTAIL.n423 VTAIL.n357 0.155672
R864 VTAIL.n416 VTAIL.n357 0.155672
R865 VTAIL.n416 VTAIL.n415 0.155672
R866 VTAIL.n415 VTAIL.n361 0.155672
R867 VTAIL.n408 VTAIL.n361 0.155672
R868 VTAIL.n408 VTAIL.n407 0.155672
R869 VTAIL.n407 VTAIL.n365 0.155672
R870 VTAIL.n399 VTAIL.n365 0.155672
R871 VTAIL.n399 VTAIL.n398 0.155672
R872 VTAIL.n398 VTAIL.n369 0.155672
R873 VTAIL.n391 VTAIL.n369 0.155672
R874 VTAIL.n391 VTAIL.n390 0.155672
R875 VTAIL.n390 VTAIL.n374 0.155672
R876 VTAIL.n383 VTAIL.n374 0.155672
R877 VTAIL.n383 VTAIL.n382 0.155672
R878 VTAIL.n353 VTAIL.n287 0.155672
R879 VTAIL.n346 VTAIL.n287 0.155672
R880 VTAIL.n346 VTAIL.n345 0.155672
R881 VTAIL.n345 VTAIL.n291 0.155672
R882 VTAIL.n338 VTAIL.n291 0.155672
R883 VTAIL.n338 VTAIL.n337 0.155672
R884 VTAIL.n337 VTAIL.n295 0.155672
R885 VTAIL.n329 VTAIL.n295 0.155672
R886 VTAIL.n329 VTAIL.n328 0.155672
R887 VTAIL.n328 VTAIL.n299 0.155672
R888 VTAIL.n321 VTAIL.n299 0.155672
R889 VTAIL.n321 VTAIL.n320 0.155672
R890 VTAIL.n320 VTAIL.n304 0.155672
R891 VTAIL.n313 VTAIL.n304 0.155672
R892 VTAIL.n313 VTAIL.n312 0.155672
R893 VTAIL.n281 VTAIL.n215 0.155672
R894 VTAIL.n274 VTAIL.n215 0.155672
R895 VTAIL.n274 VTAIL.n273 0.155672
R896 VTAIL.n273 VTAIL.n219 0.155672
R897 VTAIL.n266 VTAIL.n219 0.155672
R898 VTAIL.n266 VTAIL.n265 0.155672
R899 VTAIL.n265 VTAIL.n223 0.155672
R900 VTAIL.n257 VTAIL.n223 0.155672
R901 VTAIL.n257 VTAIL.n256 0.155672
R902 VTAIL.n256 VTAIL.n227 0.155672
R903 VTAIL.n249 VTAIL.n227 0.155672
R904 VTAIL.n249 VTAIL.n248 0.155672
R905 VTAIL.n248 VTAIL.n232 0.155672
R906 VTAIL.n241 VTAIL.n232 0.155672
R907 VTAIL.n241 VTAIL.n240 0.155672
R908 VTAIL VTAIL.n1 0.0586897
R909 VP.n4 VP.t4 731.687
R910 VP.n10 VP.t0 710.705
R911 VP.n1 VP.t2 710.705
R912 VP.n15 VP.t1 710.705
R913 VP.n16 VP.t7 710.705
R914 VP.n8 VP.t5 710.705
R915 VP.n7 VP.t3 710.705
R916 VP.n3 VP.t6 710.705
R917 VP.n17 VP.n16 161.3
R918 VP.n6 VP.n5 161.3
R919 VP.n7 VP.n2 161.3
R920 VP.n9 VP.n8 161.3
R921 VP.n15 VP.n0 161.3
R922 VP.n14 VP.n13 161.3
R923 VP.n12 VP.n1 161.3
R924 VP.n11 VP.n10 161.3
R925 VP.n5 VP.n4 70.4033
R926 VP.n10 VP.n1 48.2005
R927 VP.n16 VP.n15 48.2005
R928 VP.n8 VP.n7 48.2005
R929 VP.n11 VP.n9 41.7126
R930 VP.n14 VP.n1 24.1005
R931 VP.n15 VP.n14 24.1005
R932 VP.n6 VP.n3 24.1005
R933 VP.n7 VP.n6 24.1005
R934 VP.n4 VP.n3 20.9576
R935 VP.n5 VP.n2 0.189894
R936 VP.n9 VP.n2 0.189894
R937 VP.n12 VP.n11 0.189894
R938 VP.n13 VP.n12 0.189894
R939 VP.n13 VP.n0 0.189894
R940 VP.n17 VP.n0 0.189894
R941 VP VP.n17 0.0516364
R942 VDD1 VDD1.n0 72.8412
R943 VDD1.n3 VDD1.n2 72.7276
R944 VDD1.n3 VDD1.n1 72.7276
R945 VDD1.n5 VDD1.n4 72.4293
R946 VDD1.n5 VDD1.n3 38.5224
R947 VDD1.n4 VDD1.t4 2.53797
R948 VDD1.n4 VDD1.t2 2.53797
R949 VDD1.n0 VDD1.t3 2.53797
R950 VDD1.n0 VDD1.t1 2.53797
R951 VDD1.n2 VDD1.t6 2.53797
R952 VDD1.n2 VDD1.t0 2.53797
R953 VDD1.n1 VDD1.t7 2.53797
R954 VDD1.n1 VDD1.t5 2.53797
R955 VDD1 VDD1.n5 0.295759
R956 B.n108 B.t0 836.697
R957 B.n116 B.t9 836.697
R958 B.n34 B.t6 836.697
R959 B.n42 B.t3 836.697
R960 B.n388 B.n65 585
R961 B.n390 B.n389 585
R962 B.n391 B.n64 585
R963 B.n393 B.n392 585
R964 B.n394 B.n63 585
R965 B.n396 B.n395 585
R966 B.n397 B.n62 585
R967 B.n399 B.n398 585
R968 B.n400 B.n61 585
R969 B.n402 B.n401 585
R970 B.n403 B.n60 585
R971 B.n405 B.n404 585
R972 B.n406 B.n59 585
R973 B.n408 B.n407 585
R974 B.n409 B.n58 585
R975 B.n411 B.n410 585
R976 B.n412 B.n57 585
R977 B.n414 B.n413 585
R978 B.n415 B.n56 585
R979 B.n417 B.n416 585
R980 B.n418 B.n55 585
R981 B.n420 B.n419 585
R982 B.n421 B.n54 585
R983 B.n423 B.n422 585
R984 B.n424 B.n53 585
R985 B.n426 B.n425 585
R986 B.n427 B.n52 585
R987 B.n429 B.n428 585
R988 B.n430 B.n51 585
R989 B.n432 B.n431 585
R990 B.n433 B.n50 585
R991 B.n435 B.n434 585
R992 B.n436 B.n49 585
R993 B.n438 B.n437 585
R994 B.n439 B.n48 585
R995 B.n441 B.n440 585
R996 B.n442 B.n47 585
R997 B.n444 B.n443 585
R998 B.n445 B.n46 585
R999 B.n447 B.n446 585
R1000 B.n448 B.n45 585
R1001 B.n450 B.n449 585
R1002 B.n451 B.n44 585
R1003 B.n453 B.n452 585
R1004 B.n455 B.n41 585
R1005 B.n457 B.n456 585
R1006 B.n458 B.n40 585
R1007 B.n460 B.n459 585
R1008 B.n461 B.n39 585
R1009 B.n463 B.n462 585
R1010 B.n464 B.n38 585
R1011 B.n466 B.n465 585
R1012 B.n467 B.n37 585
R1013 B.n469 B.n468 585
R1014 B.n471 B.n470 585
R1015 B.n472 B.n33 585
R1016 B.n474 B.n473 585
R1017 B.n475 B.n32 585
R1018 B.n477 B.n476 585
R1019 B.n478 B.n31 585
R1020 B.n480 B.n479 585
R1021 B.n481 B.n30 585
R1022 B.n483 B.n482 585
R1023 B.n484 B.n29 585
R1024 B.n486 B.n485 585
R1025 B.n487 B.n28 585
R1026 B.n489 B.n488 585
R1027 B.n490 B.n27 585
R1028 B.n492 B.n491 585
R1029 B.n493 B.n26 585
R1030 B.n495 B.n494 585
R1031 B.n496 B.n25 585
R1032 B.n498 B.n497 585
R1033 B.n499 B.n24 585
R1034 B.n501 B.n500 585
R1035 B.n502 B.n23 585
R1036 B.n504 B.n503 585
R1037 B.n505 B.n22 585
R1038 B.n507 B.n506 585
R1039 B.n508 B.n21 585
R1040 B.n510 B.n509 585
R1041 B.n511 B.n20 585
R1042 B.n513 B.n512 585
R1043 B.n514 B.n19 585
R1044 B.n516 B.n515 585
R1045 B.n517 B.n18 585
R1046 B.n519 B.n518 585
R1047 B.n520 B.n17 585
R1048 B.n522 B.n521 585
R1049 B.n523 B.n16 585
R1050 B.n525 B.n524 585
R1051 B.n526 B.n15 585
R1052 B.n528 B.n527 585
R1053 B.n529 B.n14 585
R1054 B.n531 B.n530 585
R1055 B.n532 B.n13 585
R1056 B.n534 B.n533 585
R1057 B.n535 B.n12 585
R1058 B.n387 B.n386 585
R1059 B.n385 B.n66 585
R1060 B.n384 B.n383 585
R1061 B.n382 B.n67 585
R1062 B.n381 B.n380 585
R1063 B.n379 B.n68 585
R1064 B.n378 B.n377 585
R1065 B.n376 B.n69 585
R1066 B.n375 B.n374 585
R1067 B.n373 B.n70 585
R1068 B.n372 B.n371 585
R1069 B.n370 B.n71 585
R1070 B.n369 B.n368 585
R1071 B.n367 B.n72 585
R1072 B.n366 B.n365 585
R1073 B.n364 B.n73 585
R1074 B.n363 B.n362 585
R1075 B.n361 B.n74 585
R1076 B.n360 B.n359 585
R1077 B.n358 B.n75 585
R1078 B.n357 B.n356 585
R1079 B.n355 B.n76 585
R1080 B.n354 B.n353 585
R1081 B.n352 B.n77 585
R1082 B.n351 B.n350 585
R1083 B.n349 B.n78 585
R1084 B.n348 B.n347 585
R1085 B.n346 B.n79 585
R1086 B.n345 B.n344 585
R1087 B.n343 B.n80 585
R1088 B.n342 B.n341 585
R1089 B.n340 B.n81 585
R1090 B.n339 B.n338 585
R1091 B.n337 B.n82 585
R1092 B.n336 B.n335 585
R1093 B.n334 B.n83 585
R1094 B.n333 B.n332 585
R1095 B.n331 B.n84 585
R1096 B.n330 B.n329 585
R1097 B.n328 B.n85 585
R1098 B.n327 B.n326 585
R1099 B.n178 B.n139 585
R1100 B.n180 B.n179 585
R1101 B.n181 B.n138 585
R1102 B.n183 B.n182 585
R1103 B.n184 B.n137 585
R1104 B.n186 B.n185 585
R1105 B.n187 B.n136 585
R1106 B.n189 B.n188 585
R1107 B.n190 B.n135 585
R1108 B.n192 B.n191 585
R1109 B.n193 B.n134 585
R1110 B.n195 B.n194 585
R1111 B.n196 B.n133 585
R1112 B.n198 B.n197 585
R1113 B.n199 B.n132 585
R1114 B.n201 B.n200 585
R1115 B.n202 B.n131 585
R1116 B.n204 B.n203 585
R1117 B.n205 B.n130 585
R1118 B.n207 B.n206 585
R1119 B.n208 B.n129 585
R1120 B.n210 B.n209 585
R1121 B.n211 B.n128 585
R1122 B.n213 B.n212 585
R1123 B.n214 B.n127 585
R1124 B.n216 B.n215 585
R1125 B.n217 B.n126 585
R1126 B.n219 B.n218 585
R1127 B.n220 B.n125 585
R1128 B.n222 B.n221 585
R1129 B.n223 B.n124 585
R1130 B.n225 B.n224 585
R1131 B.n226 B.n123 585
R1132 B.n228 B.n227 585
R1133 B.n229 B.n122 585
R1134 B.n231 B.n230 585
R1135 B.n232 B.n121 585
R1136 B.n234 B.n233 585
R1137 B.n235 B.n120 585
R1138 B.n237 B.n236 585
R1139 B.n238 B.n119 585
R1140 B.n240 B.n239 585
R1141 B.n241 B.n118 585
R1142 B.n243 B.n242 585
R1143 B.n245 B.n115 585
R1144 B.n247 B.n246 585
R1145 B.n248 B.n114 585
R1146 B.n250 B.n249 585
R1147 B.n251 B.n113 585
R1148 B.n253 B.n252 585
R1149 B.n254 B.n112 585
R1150 B.n256 B.n255 585
R1151 B.n257 B.n111 585
R1152 B.n259 B.n258 585
R1153 B.n261 B.n260 585
R1154 B.n262 B.n107 585
R1155 B.n264 B.n263 585
R1156 B.n265 B.n106 585
R1157 B.n267 B.n266 585
R1158 B.n268 B.n105 585
R1159 B.n270 B.n269 585
R1160 B.n271 B.n104 585
R1161 B.n273 B.n272 585
R1162 B.n274 B.n103 585
R1163 B.n276 B.n275 585
R1164 B.n277 B.n102 585
R1165 B.n279 B.n278 585
R1166 B.n280 B.n101 585
R1167 B.n282 B.n281 585
R1168 B.n283 B.n100 585
R1169 B.n285 B.n284 585
R1170 B.n286 B.n99 585
R1171 B.n288 B.n287 585
R1172 B.n289 B.n98 585
R1173 B.n291 B.n290 585
R1174 B.n292 B.n97 585
R1175 B.n294 B.n293 585
R1176 B.n295 B.n96 585
R1177 B.n297 B.n296 585
R1178 B.n298 B.n95 585
R1179 B.n300 B.n299 585
R1180 B.n301 B.n94 585
R1181 B.n303 B.n302 585
R1182 B.n304 B.n93 585
R1183 B.n306 B.n305 585
R1184 B.n307 B.n92 585
R1185 B.n309 B.n308 585
R1186 B.n310 B.n91 585
R1187 B.n312 B.n311 585
R1188 B.n313 B.n90 585
R1189 B.n315 B.n314 585
R1190 B.n316 B.n89 585
R1191 B.n318 B.n317 585
R1192 B.n319 B.n88 585
R1193 B.n321 B.n320 585
R1194 B.n322 B.n87 585
R1195 B.n324 B.n323 585
R1196 B.n325 B.n86 585
R1197 B.n177 B.n176 585
R1198 B.n175 B.n140 585
R1199 B.n174 B.n173 585
R1200 B.n172 B.n141 585
R1201 B.n171 B.n170 585
R1202 B.n169 B.n142 585
R1203 B.n168 B.n167 585
R1204 B.n166 B.n143 585
R1205 B.n165 B.n164 585
R1206 B.n163 B.n144 585
R1207 B.n162 B.n161 585
R1208 B.n160 B.n145 585
R1209 B.n159 B.n158 585
R1210 B.n157 B.n146 585
R1211 B.n156 B.n155 585
R1212 B.n154 B.n147 585
R1213 B.n153 B.n152 585
R1214 B.n151 B.n148 585
R1215 B.n150 B.n149 585
R1216 B.n2 B.n0 585
R1217 B.n565 B.n1 585
R1218 B.n564 B.n563 585
R1219 B.n562 B.n3 585
R1220 B.n561 B.n560 585
R1221 B.n559 B.n4 585
R1222 B.n558 B.n557 585
R1223 B.n556 B.n5 585
R1224 B.n555 B.n554 585
R1225 B.n553 B.n6 585
R1226 B.n552 B.n551 585
R1227 B.n550 B.n7 585
R1228 B.n549 B.n548 585
R1229 B.n547 B.n8 585
R1230 B.n546 B.n545 585
R1231 B.n544 B.n9 585
R1232 B.n543 B.n542 585
R1233 B.n541 B.n10 585
R1234 B.n540 B.n539 585
R1235 B.n538 B.n11 585
R1236 B.n537 B.n536 585
R1237 B.n567 B.n566 585
R1238 B.n176 B.n139 492.5
R1239 B.n536 B.n535 492.5
R1240 B.n326 B.n325 492.5
R1241 B.n386 B.n65 492.5
R1242 B.n108 B.t2 406.202
R1243 B.n42 B.t4 406.202
R1244 B.n116 B.t11 406.202
R1245 B.n34 B.t7 406.202
R1246 B.n109 B.t1 390.298
R1247 B.n43 B.t5 390.298
R1248 B.n117 B.t10 390.298
R1249 B.n35 B.t8 390.298
R1250 B.n176 B.n175 163.367
R1251 B.n175 B.n174 163.367
R1252 B.n174 B.n141 163.367
R1253 B.n170 B.n141 163.367
R1254 B.n170 B.n169 163.367
R1255 B.n169 B.n168 163.367
R1256 B.n168 B.n143 163.367
R1257 B.n164 B.n143 163.367
R1258 B.n164 B.n163 163.367
R1259 B.n163 B.n162 163.367
R1260 B.n162 B.n145 163.367
R1261 B.n158 B.n145 163.367
R1262 B.n158 B.n157 163.367
R1263 B.n157 B.n156 163.367
R1264 B.n156 B.n147 163.367
R1265 B.n152 B.n147 163.367
R1266 B.n152 B.n151 163.367
R1267 B.n151 B.n150 163.367
R1268 B.n150 B.n2 163.367
R1269 B.n566 B.n2 163.367
R1270 B.n566 B.n565 163.367
R1271 B.n565 B.n564 163.367
R1272 B.n564 B.n3 163.367
R1273 B.n560 B.n3 163.367
R1274 B.n560 B.n559 163.367
R1275 B.n559 B.n558 163.367
R1276 B.n558 B.n5 163.367
R1277 B.n554 B.n5 163.367
R1278 B.n554 B.n553 163.367
R1279 B.n553 B.n552 163.367
R1280 B.n552 B.n7 163.367
R1281 B.n548 B.n7 163.367
R1282 B.n548 B.n547 163.367
R1283 B.n547 B.n546 163.367
R1284 B.n546 B.n9 163.367
R1285 B.n542 B.n9 163.367
R1286 B.n542 B.n541 163.367
R1287 B.n541 B.n540 163.367
R1288 B.n540 B.n11 163.367
R1289 B.n536 B.n11 163.367
R1290 B.n180 B.n139 163.367
R1291 B.n181 B.n180 163.367
R1292 B.n182 B.n181 163.367
R1293 B.n182 B.n137 163.367
R1294 B.n186 B.n137 163.367
R1295 B.n187 B.n186 163.367
R1296 B.n188 B.n187 163.367
R1297 B.n188 B.n135 163.367
R1298 B.n192 B.n135 163.367
R1299 B.n193 B.n192 163.367
R1300 B.n194 B.n193 163.367
R1301 B.n194 B.n133 163.367
R1302 B.n198 B.n133 163.367
R1303 B.n199 B.n198 163.367
R1304 B.n200 B.n199 163.367
R1305 B.n200 B.n131 163.367
R1306 B.n204 B.n131 163.367
R1307 B.n205 B.n204 163.367
R1308 B.n206 B.n205 163.367
R1309 B.n206 B.n129 163.367
R1310 B.n210 B.n129 163.367
R1311 B.n211 B.n210 163.367
R1312 B.n212 B.n211 163.367
R1313 B.n212 B.n127 163.367
R1314 B.n216 B.n127 163.367
R1315 B.n217 B.n216 163.367
R1316 B.n218 B.n217 163.367
R1317 B.n218 B.n125 163.367
R1318 B.n222 B.n125 163.367
R1319 B.n223 B.n222 163.367
R1320 B.n224 B.n223 163.367
R1321 B.n224 B.n123 163.367
R1322 B.n228 B.n123 163.367
R1323 B.n229 B.n228 163.367
R1324 B.n230 B.n229 163.367
R1325 B.n230 B.n121 163.367
R1326 B.n234 B.n121 163.367
R1327 B.n235 B.n234 163.367
R1328 B.n236 B.n235 163.367
R1329 B.n236 B.n119 163.367
R1330 B.n240 B.n119 163.367
R1331 B.n241 B.n240 163.367
R1332 B.n242 B.n241 163.367
R1333 B.n242 B.n115 163.367
R1334 B.n247 B.n115 163.367
R1335 B.n248 B.n247 163.367
R1336 B.n249 B.n248 163.367
R1337 B.n249 B.n113 163.367
R1338 B.n253 B.n113 163.367
R1339 B.n254 B.n253 163.367
R1340 B.n255 B.n254 163.367
R1341 B.n255 B.n111 163.367
R1342 B.n259 B.n111 163.367
R1343 B.n260 B.n259 163.367
R1344 B.n260 B.n107 163.367
R1345 B.n264 B.n107 163.367
R1346 B.n265 B.n264 163.367
R1347 B.n266 B.n265 163.367
R1348 B.n266 B.n105 163.367
R1349 B.n270 B.n105 163.367
R1350 B.n271 B.n270 163.367
R1351 B.n272 B.n271 163.367
R1352 B.n272 B.n103 163.367
R1353 B.n276 B.n103 163.367
R1354 B.n277 B.n276 163.367
R1355 B.n278 B.n277 163.367
R1356 B.n278 B.n101 163.367
R1357 B.n282 B.n101 163.367
R1358 B.n283 B.n282 163.367
R1359 B.n284 B.n283 163.367
R1360 B.n284 B.n99 163.367
R1361 B.n288 B.n99 163.367
R1362 B.n289 B.n288 163.367
R1363 B.n290 B.n289 163.367
R1364 B.n290 B.n97 163.367
R1365 B.n294 B.n97 163.367
R1366 B.n295 B.n294 163.367
R1367 B.n296 B.n295 163.367
R1368 B.n296 B.n95 163.367
R1369 B.n300 B.n95 163.367
R1370 B.n301 B.n300 163.367
R1371 B.n302 B.n301 163.367
R1372 B.n302 B.n93 163.367
R1373 B.n306 B.n93 163.367
R1374 B.n307 B.n306 163.367
R1375 B.n308 B.n307 163.367
R1376 B.n308 B.n91 163.367
R1377 B.n312 B.n91 163.367
R1378 B.n313 B.n312 163.367
R1379 B.n314 B.n313 163.367
R1380 B.n314 B.n89 163.367
R1381 B.n318 B.n89 163.367
R1382 B.n319 B.n318 163.367
R1383 B.n320 B.n319 163.367
R1384 B.n320 B.n87 163.367
R1385 B.n324 B.n87 163.367
R1386 B.n325 B.n324 163.367
R1387 B.n326 B.n85 163.367
R1388 B.n330 B.n85 163.367
R1389 B.n331 B.n330 163.367
R1390 B.n332 B.n331 163.367
R1391 B.n332 B.n83 163.367
R1392 B.n336 B.n83 163.367
R1393 B.n337 B.n336 163.367
R1394 B.n338 B.n337 163.367
R1395 B.n338 B.n81 163.367
R1396 B.n342 B.n81 163.367
R1397 B.n343 B.n342 163.367
R1398 B.n344 B.n343 163.367
R1399 B.n344 B.n79 163.367
R1400 B.n348 B.n79 163.367
R1401 B.n349 B.n348 163.367
R1402 B.n350 B.n349 163.367
R1403 B.n350 B.n77 163.367
R1404 B.n354 B.n77 163.367
R1405 B.n355 B.n354 163.367
R1406 B.n356 B.n355 163.367
R1407 B.n356 B.n75 163.367
R1408 B.n360 B.n75 163.367
R1409 B.n361 B.n360 163.367
R1410 B.n362 B.n361 163.367
R1411 B.n362 B.n73 163.367
R1412 B.n366 B.n73 163.367
R1413 B.n367 B.n366 163.367
R1414 B.n368 B.n367 163.367
R1415 B.n368 B.n71 163.367
R1416 B.n372 B.n71 163.367
R1417 B.n373 B.n372 163.367
R1418 B.n374 B.n373 163.367
R1419 B.n374 B.n69 163.367
R1420 B.n378 B.n69 163.367
R1421 B.n379 B.n378 163.367
R1422 B.n380 B.n379 163.367
R1423 B.n380 B.n67 163.367
R1424 B.n384 B.n67 163.367
R1425 B.n385 B.n384 163.367
R1426 B.n386 B.n385 163.367
R1427 B.n535 B.n534 163.367
R1428 B.n534 B.n13 163.367
R1429 B.n530 B.n13 163.367
R1430 B.n530 B.n529 163.367
R1431 B.n529 B.n528 163.367
R1432 B.n528 B.n15 163.367
R1433 B.n524 B.n15 163.367
R1434 B.n524 B.n523 163.367
R1435 B.n523 B.n522 163.367
R1436 B.n522 B.n17 163.367
R1437 B.n518 B.n17 163.367
R1438 B.n518 B.n517 163.367
R1439 B.n517 B.n516 163.367
R1440 B.n516 B.n19 163.367
R1441 B.n512 B.n19 163.367
R1442 B.n512 B.n511 163.367
R1443 B.n511 B.n510 163.367
R1444 B.n510 B.n21 163.367
R1445 B.n506 B.n21 163.367
R1446 B.n506 B.n505 163.367
R1447 B.n505 B.n504 163.367
R1448 B.n504 B.n23 163.367
R1449 B.n500 B.n23 163.367
R1450 B.n500 B.n499 163.367
R1451 B.n499 B.n498 163.367
R1452 B.n498 B.n25 163.367
R1453 B.n494 B.n25 163.367
R1454 B.n494 B.n493 163.367
R1455 B.n493 B.n492 163.367
R1456 B.n492 B.n27 163.367
R1457 B.n488 B.n27 163.367
R1458 B.n488 B.n487 163.367
R1459 B.n487 B.n486 163.367
R1460 B.n486 B.n29 163.367
R1461 B.n482 B.n29 163.367
R1462 B.n482 B.n481 163.367
R1463 B.n481 B.n480 163.367
R1464 B.n480 B.n31 163.367
R1465 B.n476 B.n31 163.367
R1466 B.n476 B.n475 163.367
R1467 B.n475 B.n474 163.367
R1468 B.n474 B.n33 163.367
R1469 B.n470 B.n33 163.367
R1470 B.n470 B.n469 163.367
R1471 B.n469 B.n37 163.367
R1472 B.n465 B.n37 163.367
R1473 B.n465 B.n464 163.367
R1474 B.n464 B.n463 163.367
R1475 B.n463 B.n39 163.367
R1476 B.n459 B.n39 163.367
R1477 B.n459 B.n458 163.367
R1478 B.n458 B.n457 163.367
R1479 B.n457 B.n41 163.367
R1480 B.n452 B.n41 163.367
R1481 B.n452 B.n451 163.367
R1482 B.n451 B.n450 163.367
R1483 B.n450 B.n45 163.367
R1484 B.n446 B.n45 163.367
R1485 B.n446 B.n445 163.367
R1486 B.n445 B.n444 163.367
R1487 B.n444 B.n47 163.367
R1488 B.n440 B.n47 163.367
R1489 B.n440 B.n439 163.367
R1490 B.n439 B.n438 163.367
R1491 B.n438 B.n49 163.367
R1492 B.n434 B.n49 163.367
R1493 B.n434 B.n433 163.367
R1494 B.n433 B.n432 163.367
R1495 B.n432 B.n51 163.367
R1496 B.n428 B.n51 163.367
R1497 B.n428 B.n427 163.367
R1498 B.n427 B.n426 163.367
R1499 B.n426 B.n53 163.367
R1500 B.n422 B.n53 163.367
R1501 B.n422 B.n421 163.367
R1502 B.n421 B.n420 163.367
R1503 B.n420 B.n55 163.367
R1504 B.n416 B.n55 163.367
R1505 B.n416 B.n415 163.367
R1506 B.n415 B.n414 163.367
R1507 B.n414 B.n57 163.367
R1508 B.n410 B.n57 163.367
R1509 B.n410 B.n409 163.367
R1510 B.n409 B.n408 163.367
R1511 B.n408 B.n59 163.367
R1512 B.n404 B.n59 163.367
R1513 B.n404 B.n403 163.367
R1514 B.n403 B.n402 163.367
R1515 B.n402 B.n61 163.367
R1516 B.n398 B.n61 163.367
R1517 B.n398 B.n397 163.367
R1518 B.n397 B.n396 163.367
R1519 B.n396 B.n63 163.367
R1520 B.n392 B.n63 163.367
R1521 B.n392 B.n391 163.367
R1522 B.n391 B.n390 163.367
R1523 B.n390 B.n65 163.367
R1524 B.n110 B.n109 59.5399
R1525 B.n244 B.n117 59.5399
R1526 B.n36 B.n35 59.5399
R1527 B.n454 B.n43 59.5399
R1528 B.n537 B.n12 32.0005
R1529 B.n388 B.n387 32.0005
R1530 B.n327 B.n86 32.0005
R1531 B.n178 B.n177 32.0005
R1532 B B.n567 18.0485
R1533 B.n109 B.n108 15.9035
R1534 B.n117 B.n116 15.9035
R1535 B.n35 B.n34 15.9035
R1536 B.n43 B.n42 15.9035
R1537 B.n533 B.n12 10.6151
R1538 B.n533 B.n532 10.6151
R1539 B.n532 B.n531 10.6151
R1540 B.n531 B.n14 10.6151
R1541 B.n527 B.n14 10.6151
R1542 B.n527 B.n526 10.6151
R1543 B.n526 B.n525 10.6151
R1544 B.n525 B.n16 10.6151
R1545 B.n521 B.n16 10.6151
R1546 B.n521 B.n520 10.6151
R1547 B.n520 B.n519 10.6151
R1548 B.n519 B.n18 10.6151
R1549 B.n515 B.n18 10.6151
R1550 B.n515 B.n514 10.6151
R1551 B.n514 B.n513 10.6151
R1552 B.n513 B.n20 10.6151
R1553 B.n509 B.n20 10.6151
R1554 B.n509 B.n508 10.6151
R1555 B.n508 B.n507 10.6151
R1556 B.n507 B.n22 10.6151
R1557 B.n503 B.n22 10.6151
R1558 B.n503 B.n502 10.6151
R1559 B.n502 B.n501 10.6151
R1560 B.n501 B.n24 10.6151
R1561 B.n497 B.n24 10.6151
R1562 B.n497 B.n496 10.6151
R1563 B.n496 B.n495 10.6151
R1564 B.n495 B.n26 10.6151
R1565 B.n491 B.n26 10.6151
R1566 B.n491 B.n490 10.6151
R1567 B.n490 B.n489 10.6151
R1568 B.n489 B.n28 10.6151
R1569 B.n485 B.n28 10.6151
R1570 B.n485 B.n484 10.6151
R1571 B.n484 B.n483 10.6151
R1572 B.n483 B.n30 10.6151
R1573 B.n479 B.n30 10.6151
R1574 B.n479 B.n478 10.6151
R1575 B.n478 B.n477 10.6151
R1576 B.n477 B.n32 10.6151
R1577 B.n473 B.n32 10.6151
R1578 B.n473 B.n472 10.6151
R1579 B.n472 B.n471 10.6151
R1580 B.n468 B.n467 10.6151
R1581 B.n467 B.n466 10.6151
R1582 B.n466 B.n38 10.6151
R1583 B.n462 B.n38 10.6151
R1584 B.n462 B.n461 10.6151
R1585 B.n461 B.n460 10.6151
R1586 B.n460 B.n40 10.6151
R1587 B.n456 B.n40 10.6151
R1588 B.n456 B.n455 10.6151
R1589 B.n453 B.n44 10.6151
R1590 B.n449 B.n44 10.6151
R1591 B.n449 B.n448 10.6151
R1592 B.n448 B.n447 10.6151
R1593 B.n447 B.n46 10.6151
R1594 B.n443 B.n46 10.6151
R1595 B.n443 B.n442 10.6151
R1596 B.n442 B.n441 10.6151
R1597 B.n441 B.n48 10.6151
R1598 B.n437 B.n48 10.6151
R1599 B.n437 B.n436 10.6151
R1600 B.n436 B.n435 10.6151
R1601 B.n435 B.n50 10.6151
R1602 B.n431 B.n50 10.6151
R1603 B.n431 B.n430 10.6151
R1604 B.n430 B.n429 10.6151
R1605 B.n429 B.n52 10.6151
R1606 B.n425 B.n52 10.6151
R1607 B.n425 B.n424 10.6151
R1608 B.n424 B.n423 10.6151
R1609 B.n423 B.n54 10.6151
R1610 B.n419 B.n54 10.6151
R1611 B.n419 B.n418 10.6151
R1612 B.n418 B.n417 10.6151
R1613 B.n417 B.n56 10.6151
R1614 B.n413 B.n56 10.6151
R1615 B.n413 B.n412 10.6151
R1616 B.n412 B.n411 10.6151
R1617 B.n411 B.n58 10.6151
R1618 B.n407 B.n58 10.6151
R1619 B.n407 B.n406 10.6151
R1620 B.n406 B.n405 10.6151
R1621 B.n405 B.n60 10.6151
R1622 B.n401 B.n60 10.6151
R1623 B.n401 B.n400 10.6151
R1624 B.n400 B.n399 10.6151
R1625 B.n399 B.n62 10.6151
R1626 B.n395 B.n62 10.6151
R1627 B.n395 B.n394 10.6151
R1628 B.n394 B.n393 10.6151
R1629 B.n393 B.n64 10.6151
R1630 B.n389 B.n64 10.6151
R1631 B.n389 B.n388 10.6151
R1632 B.n328 B.n327 10.6151
R1633 B.n329 B.n328 10.6151
R1634 B.n329 B.n84 10.6151
R1635 B.n333 B.n84 10.6151
R1636 B.n334 B.n333 10.6151
R1637 B.n335 B.n334 10.6151
R1638 B.n335 B.n82 10.6151
R1639 B.n339 B.n82 10.6151
R1640 B.n340 B.n339 10.6151
R1641 B.n341 B.n340 10.6151
R1642 B.n341 B.n80 10.6151
R1643 B.n345 B.n80 10.6151
R1644 B.n346 B.n345 10.6151
R1645 B.n347 B.n346 10.6151
R1646 B.n347 B.n78 10.6151
R1647 B.n351 B.n78 10.6151
R1648 B.n352 B.n351 10.6151
R1649 B.n353 B.n352 10.6151
R1650 B.n353 B.n76 10.6151
R1651 B.n357 B.n76 10.6151
R1652 B.n358 B.n357 10.6151
R1653 B.n359 B.n358 10.6151
R1654 B.n359 B.n74 10.6151
R1655 B.n363 B.n74 10.6151
R1656 B.n364 B.n363 10.6151
R1657 B.n365 B.n364 10.6151
R1658 B.n365 B.n72 10.6151
R1659 B.n369 B.n72 10.6151
R1660 B.n370 B.n369 10.6151
R1661 B.n371 B.n370 10.6151
R1662 B.n371 B.n70 10.6151
R1663 B.n375 B.n70 10.6151
R1664 B.n376 B.n375 10.6151
R1665 B.n377 B.n376 10.6151
R1666 B.n377 B.n68 10.6151
R1667 B.n381 B.n68 10.6151
R1668 B.n382 B.n381 10.6151
R1669 B.n383 B.n382 10.6151
R1670 B.n383 B.n66 10.6151
R1671 B.n387 B.n66 10.6151
R1672 B.n179 B.n178 10.6151
R1673 B.n179 B.n138 10.6151
R1674 B.n183 B.n138 10.6151
R1675 B.n184 B.n183 10.6151
R1676 B.n185 B.n184 10.6151
R1677 B.n185 B.n136 10.6151
R1678 B.n189 B.n136 10.6151
R1679 B.n190 B.n189 10.6151
R1680 B.n191 B.n190 10.6151
R1681 B.n191 B.n134 10.6151
R1682 B.n195 B.n134 10.6151
R1683 B.n196 B.n195 10.6151
R1684 B.n197 B.n196 10.6151
R1685 B.n197 B.n132 10.6151
R1686 B.n201 B.n132 10.6151
R1687 B.n202 B.n201 10.6151
R1688 B.n203 B.n202 10.6151
R1689 B.n203 B.n130 10.6151
R1690 B.n207 B.n130 10.6151
R1691 B.n208 B.n207 10.6151
R1692 B.n209 B.n208 10.6151
R1693 B.n209 B.n128 10.6151
R1694 B.n213 B.n128 10.6151
R1695 B.n214 B.n213 10.6151
R1696 B.n215 B.n214 10.6151
R1697 B.n215 B.n126 10.6151
R1698 B.n219 B.n126 10.6151
R1699 B.n220 B.n219 10.6151
R1700 B.n221 B.n220 10.6151
R1701 B.n221 B.n124 10.6151
R1702 B.n225 B.n124 10.6151
R1703 B.n226 B.n225 10.6151
R1704 B.n227 B.n226 10.6151
R1705 B.n227 B.n122 10.6151
R1706 B.n231 B.n122 10.6151
R1707 B.n232 B.n231 10.6151
R1708 B.n233 B.n232 10.6151
R1709 B.n233 B.n120 10.6151
R1710 B.n237 B.n120 10.6151
R1711 B.n238 B.n237 10.6151
R1712 B.n239 B.n238 10.6151
R1713 B.n239 B.n118 10.6151
R1714 B.n243 B.n118 10.6151
R1715 B.n246 B.n245 10.6151
R1716 B.n246 B.n114 10.6151
R1717 B.n250 B.n114 10.6151
R1718 B.n251 B.n250 10.6151
R1719 B.n252 B.n251 10.6151
R1720 B.n252 B.n112 10.6151
R1721 B.n256 B.n112 10.6151
R1722 B.n257 B.n256 10.6151
R1723 B.n258 B.n257 10.6151
R1724 B.n262 B.n261 10.6151
R1725 B.n263 B.n262 10.6151
R1726 B.n263 B.n106 10.6151
R1727 B.n267 B.n106 10.6151
R1728 B.n268 B.n267 10.6151
R1729 B.n269 B.n268 10.6151
R1730 B.n269 B.n104 10.6151
R1731 B.n273 B.n104 10.6151
R1732 B.n274 B.n273 10.6151
R1733 B.n275 B.n274 10.6151
R1734 B.n275 B.n102 10.6151
R1735 B.n279 B.n102 10.6151
R1736 B.n280 B.n279 10.6151
R1737 B.n281 B.n280 10.6151
R1738 B.n281 B.n100 10.6151
R1739 B.n285 B.n100 10.6151
R1740 B.n286 B.n285 10.6151
R1741 B.n287 B.n286 10.6151
R1742 B.n287 B.n98 10.6151
R1743 B.n291 B.n98 10.6151
R1744 B.n292 B.n291 10.6151
R1745 B.n293 B.n292 10.6151
R1746 B.n293 B.n96 10.6151
R1747 B.n297 B.n96 10.6151
R1748 B.n298 B.n297 10.6151
R1749 B.n299 B.n298 10.6151
R1750 B.n299 B.n94 10.6151
R1751 B.n303 B.n94 10.6151
R1752 B.n304 B.n303 10.6151
R1753 B.n305 B.n304 10.6151
R1754 B.n305 B.n92 10.6151
R1755 B.n309 B.n92 10.6151
R1756 B.n310 B.n309 10.6151
R1757 B.n311 B.n310 10.6151
R1758 B.n311 B.n90 10.6151
R1759 B.n315 B.n90 10.6151
R1760 B.n316 B.n315 10.6151
R1761 B.n317 B.n316 10.6151
R1762 B.n317 B.n88 10.6151
R1763 B.n321 B.n88 10.6151
R1764 B.n322 B.n321 10.6151
R1765 B.n323 B.n322 10.6151
R1766 B.n323 B.n86 10.6151
R1767 B.n177 B.n140 10.6151
R1768 B.n173 B.n140 10.6151
R1769 B.n173 B.n172 10.6151
R1770 B.n172 B.n171 10.6151
R1771 B.n171 B.n142 10.6151
R1772 B.n167 B.n142 10.6151
R1773 B.n167 B.n166 10.6151
R1774 B.n166 B.n165 10.6151
R1775 B.n165 B.n144 10.6151
R1776 B.n161 B.n144 10.6151
R1777 B.n161 B.n160 10.6151
R1778 B.n160 B.n159 10.6151
R1779 B.n159 B.n146 10.6151
R1780 B.n155 B.n146 10.6151
R1781 B.n155 B.n154 10.6151
R1782 B.n154 B.n153 10.6151
R1783 B.n153 B.n148 10.6151
R1784 B.n149 B.n148 10.6151
R1785 B.n149 B.n0 10.6151
R1786 B.n563 B.n1 10.6151
R1787 B.n563 B.n562 10.6151
R1788 B.n562 B.n561 10.6151
R1789 B.n561 B.n4 10.6151
R1790 B.n557 B.n4 10.6151
R1791 B.n557 B.n556 10.6151
R1792 B.n556 B.n555 10.6151
R1793 B.n555 B.n6 10.6151
R1794 B.n551 B.n6 10.6151
R1795 B.n551 B.n550 10.6151
R1796 B.n550 B.n549 10.6151
R1797 B.n549 B.n8 10.6151
R1798 B.n545 B.n8 10.6151
R1799 B.n545 B.n544 10.6151
R1800 B.n544 B.n543 10.6151
R1801 B.n543 B.n10 10.6151
R1802 B.n539 B.n10 10.6151
R1803 B.n539 B.n538 10.6151
R1804 B.n538 B.n537 10.6151
R1805 B.n471 B.n36 9.36635
R1806 B.n454 B.n453 9.36635
R1807 B.n244 B.n243 9.36635
R1808 B.n261 B.n110 9.36635
R1809 B.n567 B.n0 2.81026
R1810 B.n567 B.n1 2.81026
R1811 B.n468 B.n36 1.24928
R1812 B.n455 B.n454 1.24928
R1813 B.n245 B.n244 1.24928
R1814 B.n258 B.n110 1.24928
C0 VP VTAIL 4.45572f
C1 VDD1 VN 0.14795f
C2 w_n1790_n3530# VN 3.06412f
C3 VDD2 VDD1 0.723577f
C4 VDD2 w_n1790_n3530# 1.26567f
C5 B VDD1 1.02771f
C6 B w_n1790_n3530# 7.115149f
C7 VDD1 VP 4.94413f
C8 w_n1790_n3530# VP 3.29028f
C9 VDD2 VN 4.79722f
C10 B VN 0.740932f
C11 VDD2 B 1.05789f
C12 VN VP 5.23043f
C13 VDD2 VP 0.295181f
C14 B VP 1.1088f
C15 VDD1 VTAIL 13.8138f
C16 w_n1790_n3530# VTAIL 4.439991f
C17 VN VTAIL 4.44161f
C18 VDD1 w_n1790_n3530# 1.23953f
C19 VDD2 VTAIL 13.854099f
C20 B VTAIL 3.87386f
C21 VDD2 VSUBS 1.36463f
C22 VDD1 VSUBS 1.629444f
C23 VTAIL VSUBS 0.85206f
C24 VN VSUBS 4.62468f
C25 VP VSUBS 1.468642f
C26 B VSUBS 2.713827f
C27 w_n1790_n3530# VSUBS 77.6932f
C28 B.n0 VSUBS 0.00527f
C29 B.n1 VSUBS 0.00527f
C30 B.n2 VSUBS 0.008334f
C31 B.n3 VSUBS 0.008334f
C32 B.n4 VSUBS 0.008334f
C33 B.n5 VSUBS 0.008334f
C34 B.n6 VSUBS 0.008334f
C35 B.n7 VSUBS 0.008334f
C36 B.n8 VSUBS 0.008334f
C37 B.n9 VSUBS 0.008334f
C38 B.n10 VSUBS 0.008334f
C39 B.n11 VSUBS 0.008334f
C40 B.n12 VSUBS 0.020039f
C41 B.n13 VSUBS 0.008334f
C42 B.n14 VSUBS 0.008334f
C43 B.n15 VSUBS 0.008334f
C44 B.n16 VSUBS 0.008334f
C45 B.n17 VSUBS 0.008334f
C46 B.n18 VSUBS 0.008334f
C47 B.n19 VSUBS 0.008334f
C48 B.n20 VSUBS 0.008334f
C49 B.n21 VSUBS 0.008334f
C50 B.n22 VSUBS 0.008334f
C51 B.n23 VSUBS 0.008334f
C52 B.n24 VSUBS 0.008334f
C53 B.n25 VSUBS 0.008334f
C54 B.n26 VSUBS 0.008334f
C55 B.n27 VSUBS 0.008334f
C56 B.n28 VSUBS 0.008334f
C57 B.n29 VSUBS 0.008334f
C58 B.n30 VSUBS 0.008334f
C59 B.n31 VSUBS 0.008334f
C60 B.n32 VSUBS 0.008334f
C61 B.n33 VSUBS 0.008334f
C62 B.t8 VSUBS 0.272985f
C63 B.t7 VSUBS 0.284364f
C64 B.t6 VSUBS 0.30023f
C65 B.n34 VSUBS 0.36892f
C66 B.n35 VSUBS 0.302549f
C67 B.n36 VSUBS 0.019309f
C68 B.n37 VSUBS 0.008334f
C69 B.n38 VSUBS 0.008334f
C70 B.n39 VSUBS 0.008334f
C71 B.n40 VSUBS 0.008334f
C72 B.n41 VSUBS 0.008334f
C73 B.t5 VSUBS 0.272988f
C74 B.t4 VSUBS 0.284368f
C75 B.t3 VSUBS 0.30023f
C76 B.n42 VSUBS 0.368917f
C77 B.n43 VSUBS 0.302545f
C78 B.n44 VSUBS 0.008334f
C79 B.n45 VSUBS 0.008334f
C80 B.n46 VSUBS 0.008334f
C81 B.n47 VSUBS 0.008334f
C82 B.n48 VSUBS 0.008334f
C83 B.n49 VSUBS 0.008334f
C84 B.n50 VSUBS 0.008334f
C85 B.n51 VSUBS 0.008334f
C86 B.n52 VSUBS 0.008334f
C87 B.n53 VSUBS 0.008334f
C88 B.n54 VSUBS 0.008334f
C89 B.n55 VSUBS 0.008334f
C90 B.n56 VSUBS 0.008334f
C91 B.n57 VSUBS 0.008334f
C92 B.n58 VSUBS 0.008334f
C93 B.n59 VSUBS 0.008334f
C94 B.n60 VSUBS 0.008334f
C95 B.n61 VSUBS 0.008334f
C96 B.n62 VSUBS 0.008334f
C97 B.n63 VSUBS 0.008334f
C98 B.n64 VSUBS 0.008334f
C99 B.n65 VSUBS 0.020039f
C100 B.n66 VSUBS 0.008334f
C101 B.n67 VSUBS 0.008334f
C102 B.n68 VSUBS 0.008334f
C103 B.n69 VSUBS 0.008334f
C104 B.n70 VSUBS 0.008334f
C105 B.n71 VSUBS 0.008334f
C106 B.n72 VSUBS 0.008334f
C107 B.n73 VSUBS 0.008334f
C108 B.n74 VSUBS 0.008334f
C109 B.n75 VSUBS 0.008334f
C110 B.n76 VSUBS 0.008334f
C111 B.n77 VSUBS 0.008334f
C112 B.n78 VSUBS 0.008334f
C113 B.n79 VSUBS 0.008334f
C114 B.n80 VSUBS 0.008334f
C115 B.n81 VSUBS 0.008334f
C116 B.n82 VSUBS 0.008334f
C117 B.n83 VSUBS 0.008334f
C118 B.n84 VSUBS 0.008334f
C119 B.n85 VSUBS 0.008334f
C120 B.n86 VSUBS 0.020039f
C121 B.n87 VSUBS 0.008334f
C122 B.n88 VSUBS 0.008334f
C123 B.n89 VSUBS 0.008334f
C124 B.n90 VSUBS 0.008334f
C125 B.n91 VSUBS 0.008334f
C126 B.n92 VSUBS 0.008334f
C127 B.n93 VSUBS 0.008334f
C128 B.n94 VSUBS 0.008334f
C129 B.n95 VSUBS 0.008334f
C130 B.n96 VSUBS 0.008334f
C131 B.n97 VSUBS 0.008334f
C132 B.n98 VSUBS 0.008334f
C133 B.n99 VSUBS 0.008334f
C134 B.n100 VSUBS 0.008334f
C135 B.n101 VSUBS 0.008334f
C136 B.n102 VSUBS 0.008334f
C137 B.n103 VSUBS 0.008334f
C138 B.n104 VSUBS 0.008334f
C139 B.n105 VSUBS 0.008334f
C140 B.n106 VSUBS 0.008334f
C141 B.n107 VSUBS 0.008334f
C142 B.t1 VSUBS 0.272988f
C143 B.t2 VSUBS 0.284368f
C144 B.t0 VSUBS 0.30023f
C145 B.n108 VSUBS 0.368917f
C146 B.n109 VSUBS 0.302545f
C147 B.n110 VSUBS 0.019309f
C148 B.n111 VSUBS 0.008334f
C149 B.n112 VSUBS 0.008334f
C150 B.n113 VSUBS 0.008334f
C151 B.n114 VSUBS 0.008334f
C152 B.n115 VSUBS 0.008334f
C153 B.t10 VSUBS 0.272985f
C154 B.t11 VSUBS 0.284364f
C155 B.t9 VSUBS 0.30023f
C156 B.n116 VSUBS 0.36892f
C157 B.n117 VSUBS 0.302549f
C158 B.n118 VSUBS 0.008334f
C159 B.n119 VSUBS 0.008334f
C160 B.n120 VSUBS 0.008334f
C161 B.n121 VSUBS 0.008334f
C162 B.n122 VSUBS 0.008334f
C163 B.n123 VSUBS 0.008334f
C164 B.n124 VSUBS 0.008334f
C165 B.n125 VSUBS 0.008334f
C166 B.n126 VSUBS 0.008334f
C167 B.n127 VSUBS 0.008334f
C168 B.n128 VSUBS 0.008334f
C169 B.n129 VSUBS 0.008334f
C170 B.n130 VSUBS 0.008334f
C171 B.n131 VSUBS 0.008334f
C172 B.n132 VSUBS 0.008334f
C173 B.n133 VSUBS 0.008334f
C174 B.n134 VSUBS 0.008334f
C175 B.n135 VSUBS 0.008334f
C176 B.n136 VSUBS 0.008334f
C177 B.n137 VSUBS 0.008334f
C178 B.n138 VSUBS 0.008334f
C179 B.n139 VSUBS 0.020039f
C180 B.n140 VSUBS 0.008334f
C181 B.n141 VSUBS 0.008334f
C182 B.n142 VSUBS 0.008334f
C183 B.n143 VSUBS 0.008334f
C184 B.n144 VSUBS 0.008334f
C185 B.n145 VSUBS 0.008334f
C186 B.n146 VSUBS 0.008334f
C187 B.n147 VSUBS 0.008334f
C188 B.n148 VSUBS 0.008334f
C189 B.n149 VSUBS 0.008334f
C190 B.n150 VSUBS 0.008334f
C191 B.n151 VSUBS 0.008334f
C192 B.n152 VSUBS 0.008334f
C193 B.n153 VSUBS 0.008334f
C194 B.n154 VSUBS 0.008334f
C195 B.n155 VSUBS 0.008334f
C196 B.n156 VSUBS 0.008334f
C197 B.n157 VSUBS 0.008334f
C198 B.n158 VSUBS 0.008334f
C199 B.n159 VSUBS 0.008334f
C200 B.n160 VSUBS 0.008334f
C201 B.n161 VSUBS 0.008334f
C202 B.n162 VSUBS 0.008334f
C203 B.n163 VSUBS 0.008334f
C204 B.n164 VSUBS 0.008334f
C205 B.n165 VSUBS 0.008334f
C206 B.n166 VSUBS 0.008334f
C207 B.n167 VSUBS 0.008334f
C208 B.n168 VSUBS 0.008334f
C209 B.n169 VSUBS 0.008334f
C210 B.n170 VSUBS 0.008334f
C211 B.n171 VSUBS 0.008334f
C212 B.n172 VSUBS 0.008334f
C213 B.n173 VSUBS 0.008334f
C214 B.n174 VSUBS 0.008334f
C215 B.n175 VSUBS 0.008334f
C216 B.n176 VSUBS 0.018445f
C217 B.n177 VSUBS 0.018445f
C218 B.n178 VSUBS 0.020039f
C219 B.n179 VSUBS 0.008334f
C220 B.n180 VSUBS 0.008334f
C221 B.n181 VSUBS 0.008334f
C222 B.n182 VSUBS 0.008334f
C223 B.n183 VSUBS 0.008334f
C224 B.n184 VSUBS 0.008334f
C225 B.n185 VSUBS 0.008334f
C226 B.n186 VSUBS 0.008334f
C227 B.n187 VSUBS 0.008334f
C228 B.n188 VSUBS 0.008334f
C229 B.n189 VSUBS 0.008334f
C230 B.n190 VSUBS 0.008334f
C231 B.n191 VSUBS 0.008334f
C232 B.n192 VSUBS 0.008334f
C233 B.n193 VSUBS 0.008334f
C234 B.n194 VSUBS 0.008334f
C235 B.n195 VSUBS 0.008334f
C236 B.n196 VSUBS 0.008334f
C237 B.n197 VSUBS 0.008334f
C238 B.n198 VSUBS 0.008334f
C239 B.n199 VSUBS 0.008334f
C240 B.n200 VSUBS 0.008334f
C241 B.n201 VSUBS 0.008334f
C242 B.n202 VSUBS 0.008334f
C243 B.n203 VSUBS 0.008334f
C244 B.n204 VSUBS 0.008334f
C245 B.n205 VSUBS 0.008334f
C246 B.n206 VSUBS 0.008334f
C247 B.n207 VSUBS 0.008334f
C248 B.n208 VSUBS 0.008334f
C249 B.n209 VSUBS 0.008334f
C250 B.n210 VSUBS 0.008334f
C251 B.n211 VSUBS 0.008334f
C252 B.n212 VSUBS 0.008334f
C253 B.n213 VSUBS 0.008334f
C254 B.n214 VSUBS 0.008334f
C255 B.n215 VSUBS 0.008334f
C256 B.n216 VSUBS 0.008334f
C257 B.n217 VSUBS 0.008334f
C258 B.n218 VSUBS 0.008334f
C259 B.n219 VSUBS 0.008334f
C260 B.n220 VSUBS 0.008334f
C261 B.n221 VSUBS 0.008334f
C262 B.n222 VSUBS 0.008334f
C263 B.n223 VSUBS 0.008334f
C264 B.n224 VSUBS 0.008334f
C265 B.n225 VSUBS 0.008334f
C266 B.n226 VSUBS 0.008334f
C267 B.n227 VSUBS 0.008334f
C268 B.n228 VSUBS 0.008334f
C269 B.n229 VSUBS 0.008334f
C270 B.n230 VSUBS 0.008334f
C271 B.n231 VSUBS 0.008334f
C272 B.n232 VSUBS 0.008334f
C273 B.n233 VSUBS 0.008334f
C274 B.n234 VSUBS 0.008334f
C275 B.n235 VSUBS 0.008334f
C276 B.n236 VSUBS 0.008334f
C277 B.n237 VSUBS 0.008334f
C278 B.n238 VSUBS 0.008334f
C279 B.n239 VSUBS 0.008334f
C280 B.n240 VSUBS 0.008334f
C281 B.n241 VSUBS 0.008334f
C282 B.n242 VSUBS 0.008334f
C283 B.n243 VSUBS 0.007844f
C284 B.n244 VSUBS 0.019309f
C285 B.n245 VSUBS 0.004657f
C286 B.n246 VSUBS 0.008334f
C287 B.n247 VSUBS 0.008334f
C288 B.n248 VSUBS 0.008334f
C289 B.n249 VSUBS 0.008334f
C290 B.n250 VSUBS 0.008334f
C291 B.n251 VSUBS 0.008334f
C292 B.n252 VSUBS 0.008334f
C293 B.n253 VSUBS 0.008334f
C294 B.n254 VSUBS 0.008334f
C295 B.n255 VSUBS 0.008334f
C296 B.n256 VSUBS 0.008334f
C297 B.n257 VSUBS 0.008334f
C298 B.n258 VSUBS 0.004657f
C299 B.n259 VSUBS 0.008334f
C300 B.n260 VSUBS 0.008334f
C301 B.n261 VSUBS 0.007844f
C302 B.n262 VSUBS 0.008334f
C303 B.n263 VSUBS 0.008334f
C304 B.n264 VSUBS 0.008334f
C305 B.n265 VSUBS 0.008334f
C306 B.n266 VSUBS 0.008334f
C307 B.n267 VSUBS 0.008334f
C308 B.n268 VSUBS 0.008334f
C309 B.n269 VSUBS 0.008334f
C310 B.n270 VSUBS 0.008334f
C311 B.n271 VSUBS 0.008334f
C312 B.n272 VSUBS 0.008334f
C313 B.n273 VSUBS 0.008334f
C314 B.n274 VSUBS 0.008334f
C315 B.n275 VSUBS 0.008334f
C316 B.n276 VSUBS 0.008334f
C317 B.n277 VSUBS 0.008334f
C318 B.n278 VSUBS 0.008334f
C319 B.n279 VSUBS 0.008334f
C320 B.n280 VSUBS 0.008334f
C321 B.n281 VSUBS 0.008334f
C322 B.n282 VSUBS 0.008334f
C323 B.n283 VSUBS 0.008334f
C324 B.n284 VSUBS 0.008334f
C325 B.n285 VSUBS 0.008334f
C326 B.n286 VSUBS 0.008334f
C327 B.n287 VSUBS 0.008334f
C328 B.n288 VSUBS 0.008334f
C329 B.n289 VSUBS 0.008334f
C330 B.n290 VSUBS 0.008334f
C331 B.n291 VSUBS 0.008334f
C332 B.n292 VSUBS 0.008334f
C333 B.n293 VSUBS 0.008334f
C334 B.n294 VSUBS 0.008334f
C335 B.n295 VSUBS 0.008334f
C336 B.n296 VSUBS 0.008334f
C337 B.n297 VSUBS 0.008334f
C338 B.n298 VSUBS 0.008334f
C339 B.n299 VSUBS 0.008334f
C340 B.n300 VSUBS 0.008334f
C341 B.n301 VSUBS 0.008334f
C342 B.n302 VSUBS 0.008334f
C343 B.n303 VSUBS 0.008334f
C344 B.n304 VSUBS 0.008334f
C345 B.n305 VSUBS 0.008334f
C346 B.n306 VSUBS 0.008334f
C347 B.n307 VSUBS 0.008334f
C348 B.n308 VSUBS 0.008334f
C349 B.n309 VSUBS 0.008334f
C350 B.n310 VSUBS 0.008334f
C351 B.n311 VSUBS 0.008334f
C352 B.n312 VSUBS 0.008334f
C353 B.n313 VSUBS 0.008334f
C354 B.n314 VSUBS 0.008334f
C355 B.n315 VSUBS 0.008334f
C356 B.n316 VSUBS 0.008334f
C357 B.n317 VSUBS 0.008334f
C358 B.n318 VSUBS 0.008334f
C359 B.n319 VSUBS 0.008334f
C360 B.n320 VSUBS 0.008334f
C361 B.n321 VSUBS 0.008334f
C362 B.n322 VSUBS 0.008334f
C363 B.n323 VSUBS 0.008334f
C364 B.n324 VSUBS 0.008334f
C365 B.n325 VSUBS 0.020039f
C366 B.n326 VSUBS 0.018445f
C367 B.n327 VSUBS 0.018445f
C368 B.n328 VSUBS 0.008334f
C369 B.n329 VSUBS 0.008334f
C370 B.n330 VSUBS 0.008334f
C371 B.n331 VSUBS 0.008334f
C372 B.n332 VSUBS 0.008334f
C373 B.n333 VSUBS 0.008334f
C374 B.n334 VSUBS 0.008334f
C375 B.n335 VSUBS 0.008334f
C376 B.n336 VSUBS 0.008334f
C377 B.n337 VSUBS 0.008334f
C378 B.n338 VSUBS 0.008334f
C379 B.n339 VSUBS 0.008334f
C380 B.n340 VSUBS 0.008334f
C381 B.n341 VSUBS 0.008334f
C382 B.n342 VSUBS 0.008334f
C383 B.n343 VSUBS 0.008334f
C384 B.n344 VSUBS 0.008334f
C385 B.n345 VSUBS 0.008334f
C386 B.n346 VSUBS 0.008334f
C387 B.n347 VSUBS 0.008334f
C388 B.n348 VSUBS 0.008334f
C389 B.n349 VSUBS 0.008334f
C390 B.n350 VSUBS 0.008334f
C391 B.n351 VSUBS 0.008334f
C392 B.n352 VSUBS 0.008334f
C393 B.n353 VSUBS 0.008334f
C394 B.n354 VSUBS 0.008334f
C395 B.n355 VSUBS 0.008334f
C396 B.n356 VSUBS 0.008334f
C397 B.n357 VSUBS 0.008334f
C398 B.n358 VSUBS 0.008334f
C399 B.n359 VSUBS 0.008334f
C400 B.n360 VSUBS 0.008334f
C401 B.n361 VSUBS 0.008334f
C402 B.n362 VSUBS 0.008334f
C403 B.n363 VSUBS 0.008334f
C404 B.n364 VSUBS 0.008334f
C405 B.n365 VSUBS 0.008334f
C406 B.n366 VSUBS 0.008334f
C407 B.n367 VSUBS 0.008334f
C408 B.n368 VSUBS 0.008334f
C409 B.n369 VSUBS 0.008334f
C410 B.n370 VSUBS 0.008334f
C411 B.n371 VSUBS 0.008334f
C412 B.n372 VSUBS 0.008334f
C413 B.n373 VSUBS 0.008334f
C414 B.n374 VSUBS 0.008334f
C415 B.n375 VSUBS 0.008334f
C416 B.n376 VSUBS 0.008334f
C417 B.n377 VSUBS 0.008334f
C418 B.n378 VSUBS 0.008334f
C419 B.n379 VSUBS 0.008334f
C420 B.n380 VSUBS 0.008334f
C421 B.n381 VSUBS 0.008334f
C422 B.n382 VSUBS 0.008334f
C423 B.n383 VSUBS 0.008334f
C424 B.n384 VSUBS 0.008334f
C425 B.n385 VSUBS 0.008334f
C426 B.n386 VSUBS 0.018445f
C427 B.n387 VSUBS 0.01945f
C428 B.n388 VSUBS 0.019034f
C429 B.n389 VSUBS 0.008334f
C430 B.n390 VSUBS 0.008334f
C431 B.n391 VSUBS 0.008334f
C432 B.n392 VSUBS 0.008334f
C433 B.n393 VSUBS 0.008334f
C434 B.n394 VSUBS 0.008334f
C435 B.n395 VSUBS 0.008334f
C436 B.n396 VSUBS 0.008334f
C437 B.n397 VSUBS 0.008334f
C438 B.n398 VSUBS 0.008334f
C439 B.n399 VSUBS 0.008334f
C440 B.n400 VSUBS 0.008334f
C441 B.n401 VSUBS 0.008334f
C442 B.n402 VSUBS 0.008334f
C443 B.n403 VSUBS 0.008334f
C444 B.n404 VSUBS 0.008334f
C445 B.n405 VSUBS 0.008334f
C446 B.n406 VSUBS 0.008334f
C447 B.n407 VSUBS 0.008334f
C448 B.n408 VSUBS 0.008334f
C449 B.n409 VSUBS 0.008334f
C450 B.n410 VSUBS 0.008334f
C451 B.n411 VSUBS 0.008334f
C452 B.n412 VSUBS 0.008334f
C453 B.n413 VSUBS 0.008334f
C454 B.n414 VSUBS 0.008334f
C455 B.n415 VSUBS 0.008334f
C456 B.n416 VSUBS 0.008334f
C457 B.n417 VSUBS 0.008334f
C458 B.n418 VSUBS 0.008334f
C459 B.n419 VSUBS 0.008334f
C460 B.n420 VSUBS 0.008334f
C461 B.n421 VSUBS 0.008334f
C462 B.n422 VSUBS 0.008334f
C463 B.n423 VSUBS 0.008334f
C464 B.n424 VSUBS 0.008334f
C465 B.n425 VSUBS 0.008334f
C466 B.n426 VSUBS 0.008334f
C467 B.n427 VSUBS 0.008334f
C468 B.n428 VSUBS 0.008334f
C469 B.n429 VSUBS 0.008334f
C470 B.n430 VSUBS 0.008334f
C471 B.n431 VSUBS 0.008334f
C472 B.n432 VSUBS 0.008334f
C473 B.n433 VSUBS 0.008334f
C474 B.n434 VSUBS 0.008334f
C475 B.n435 VSUBS 0.008334f
C476 B.n436 VSUBS 0.008334f
C477 B.n437 VSUBS 0.008334f
C478 B.n438 VSUBS 0.008334f
C479 B.n439 VSUBS 0.008334f
C480 B.n440 VSUBS 0.008334f
C481 B.n441 VSUBS 0.008334f
C482 B.n442 VSUBS 0.008334f
C483 B.n443 VSUBS 0.008334f
C484 B.n444 VSUBS 0.008334f
C485 B.n445 VSUBS 0.008334f
C486 B.n446 VSUBS 0.008334f
C487 B.n447 VSUBS 0.008334f
C488 B.n448 VSUBS 0.008334f
C489 B.n449 VSUBS 0.008334f
C490 B.n450 VSUBS 0.008334f
C491 B.n451 VSUBS 0.008334f
C492 B.n452 VSUBS 0.008334f
C493 B.n453 VSUBS 0.007844f
C494 B.n454 VSUBS 0.019309f
C495 B.n455 VSUBS 0.004657f
C496 B.n456 VSUBS 0.008334f
C497 B.n457 VSUBS 0.008334f
C498 B.n458 VSUBS 0.008334f
C499 B.n459 VSUBS 0.008334f
C500 B.n460 VSUBS 0.008334f
C501 B.n461 VSUBS 0.008334f
C502 B.n462 VSUBS 0.008334f
C503 B.n463 VSUBS 0.008334f
C504 B.n464 VSUBS 0.008334f
C505 B.n465 VSUBS 0.008334f
C506 B.n466 VSUBS 0.008334f
C507 B.n467 VSUBS 0.008334f
C508 B.n468 VSUBS 0.004657f
C509 B.n469 VSUBS 0.008334f
C510 B.n470 VSUBS 0.008334f
C511 B.n471 VSUBS 0.007844f
C512 B.n472 VSUBS 0.008334f
C513 B.n473 VSUBS 0.008334f
C514 B.n474 VSUBS 0.008334f
C515 B.n475 VSUBS 0.008334f
C516 B.n476 VSUBS 0.008334f
C517 B.n477 VSUBS 0.008334f
C518 B.n478 VSUBS 0.008334f
C519 B.n479 VSUBS 0.008334f
C520 B.n480 VSUBS 0.008334f
C521 B.n481 VSUBS 0.008334f
C522 B.n482 VSUBS 0.008334f
C523 B.n483 VSUBS 0.008334f
C524 B.n484 VSUBS 0.008334f
C525 B.n485 VSUBS 0.008334f
C526 B.n486 VSUBS 0.008334f
C527 B.n487 VSUBS 0.008334f
C528 B.n488 VSUBS 0.008334f
C529 B.n489 VSUBS 0.008334f
C530 B.n490 VSUBS 0.008334f
C531 B.n491 VSUBS 0.008334f
C532 B.n492 VSUBS 0.008334f
C533 B.n493 VSUBS 0.008334f
C534 B.n494 VSUBS 0.008334f
C535 B.n495 VSUBS 0.008334f
C536 B.n496 VSUBS 0.008334f
C537 B.n497 VSUBS 0.008334f
C538 B.n498 VSUBS 0.008334f
C539 B.n499 VSUBS 0.008334f
C540 B.n500 VSUBS 0.008334f
C541 B.n501 VSUBS 0.008334f
C542 B.n502 VSUBS 0.008334f
C543 B.n503 VSUBS 0.008334f
C544 B.n504 VSUBS 0.008334f
C545 B.n505 VSUBS 0.008334f
C546 B.n506 VSUBS 0.008334f
C547 B.n507 VSUBS 0.008334f
C548 B.n508 VSUBS 0.008334f
C549 B.n509 VSUBS 0.008334f
C550 B.n510 VSUBS 0.008334f
C551 B.n511 VSUBS 0.008334f
C552 B.n512 VSUBS 0.008334f
C553 B.n513 VSUBS 0.008334f
C554 B.n514 VSUBS 0.008334f
C555 B.n515 VSUBS 0.008334f
C556 B.n516 VSUBS 0.008334f
C557 B.n517 VSUBS 0.008334f
C558 B.n518 VSUBS 0.008334f
C559 B.n519 VSUBS 0.008334f
C560 B.n520 VSUBS 0.008334f
C561 B.n521 VSUBS 0.008334f
C562 B.n522 VSUBS 0.008334f
C563 B.n523 VSUBS 0.008334f
C564 B.n524 VSUBS 0.008334f
C565 B.n525 VSUBS 0.008334f
C566 B.n526 VSUBS 0.008334f
C567 B.n527 VSUBS 0.008334f
C568 B.n528 VSUBS 0.008334f
C569 B.n529 VSUBS 0.008334f
C570 B.n530 VSUBS 0.008334f
C571 B.n531 VSUBS 0.008334f
C572 B.n532 VSUBS 0.008334f
C573 B.n533 VSUBS 0.008334f
C574 B.n534 VSUBS 0.008334f
C575 B.n535 VSUBS 0.020039f
C576 B.n536 VSUBS 0.018445f
C577 B.n537 VSUBS 0.018445f
C578 B.n538 VSUBS 0.008334f
C579 B.n539 VSUBS 0.008334f
C580 B.n540 VSUBS 0.008334f
C581 B.n541 VSUBS 0.008334f
C582 B.n542 VSUBS 0.008334f
C583 B.n543 VSUBS 0.008334f
C584 B.n544 VSUBS 0.008334f
C585 B.n545 VSUBS 0.008334f
C586 B.n546 VSUBS 0.008334f
C587 B.n547 VSUBS 0.008334f
C588 B.n548 VSUBS 0.008334f
C589 B.n549 VSUBS 0.008334f
C590 B.n550 VSUBS 0.008334f
C591 B.n551 VSUBS 0.008334f
C592 B.n552 VSUBS 0.008334f
C593 B.n553 VSUBS 0.008334f
C594 B.n554 VSUBS 0.008334f
C595 B.n555 VSUBS 0.008334f
C596 B.n556 VSUBS 0.008334f
C597 B.n557 VSUBS 0.008334f
C598 B.n558 VSUBS 0.008334f
C599 B.n559 VSUBS 0.008334f
C600 B.n560 VSUBS 0.008334f
C601 B.n561 VSUBS 0.008334f
C602 B.n562 VSUBS 0.008334f
C603 B.n563 VSUBS 0.008334f
C604 B.n564 VSUBS 0.008334f
C605 B.n565 VSUBS 0.008334f
C606 B.n566 VSUBS 0.008334f
C607 B.n567 VSUBS 0.018871f
C608 VDD1.t3 VSUBS 0.297344f
C609 VDD1.t1 VSUBS 0.297344f
C610 VDD1.n0 VSUBS 2.34616f
C611 VDD1.t7 VSUBS 0.297344f
C612 VDD1.t5 VSUBS 0.297344f
C613 VDD1.n1 VSUBS 2.34507f
C614 VDD1.t6 VSUBS 0.297344f
C615 VDD1.t0 VSUBS 0.297344f
C616 VDD1.n2 VSUBS 2.34507f
C617 VDD1.n3 VSUBS 3.16635f
C618 VDD1.t4 VSUBS 0.297344f
C619 VDD1.t2 VSUBS 0.297344f
C620 VDD1.n4 VSUBS 2.34231f
C621 VDD1.n5 VSUBS 3.03382f
C622 VP.n0 VSUBS 0.061279f
C623 VP.t2 VSUBS 1.0959f
C624 VP.n1 VSUBS 0.443969f
C625 VP.n2 VSUBS 0.061279f
C626 VP.t5 VSUBS 1.0959f
C627 VP.t3 VSUBS 1.0959f
C628 VP.t6 VSUBS 1.0959f
C629 VP.n3 VSUBS 0.443969f
C630 VP.t4 VSUBS 1.10845f
C631 VP.n4 VSUBS 0.425647f
C632 VP.n5 VSUBS 0.200372f
C633 VP.n6 VSUBS 0.013906f
C634 VP.n7 VSUBS 0.443969f
C635 VP.n8 VSUBS 0.437736f
C636 VP.n9 VSUBS 2.50056f
C637 VP.t0 VSUBS 1.0959f
C638 VP.n10 VSUBS 0.437736f
C639 VP.n11 VSUBS 2.55337f
C640 VP.n12 VSUBS 0.061279f
C641 VP.n13 VSUBS 0.061279f
C642 VP.n14 VSUBS 0.013906f
C643 VP.t1 VSUBS 1.0959f
C644 VP.n15 VSUBS 0.443969f
C645 VP.t7 VSUBS 1.0959f
C646 VP.n16 VSUBS 0.437736f
C647 VP.n17 VSUBS 0.047489f
C648 VTAIL.t14 VSUBS 0.264224f
C649 VTAIL.t9 VSUBS 0.264224f
C650 VTAIL.n0 VSUBS 1.93357f
C651 VTAIL.n1 VSUBS 0.675844f
C652 VTAIL.n2 VSUBS 0.028682f
C653 VTAIL.n3 VSUBS 0.026102f
C654 VTAIL.n4 VSUBS 0.014026f
C655 VTAIL.n5 VSUBS 0.033152f
C656 VTAIL.n6 VSUBS 0.014851f
C657 VTAIL.n7 VSUBS 0.026102f
C658 VTAIL.n8 VSUBS 0.014026f
C659 VTAIL.n9 VSUBS 0.033152f
C660 VTAIL.n10 VSUBS 0.014851f
C661 VTAIL.n11 VSUBS 0.026102f
C662 VTAIL.n12 VSUBS 0.014026f
C663 VTAIL.n13 VSUBS 0.033152f
C664 VTAIL.n14 VSUBS 0.014851f
C665 VTAIL.n15 VSUBS 0.026102f
C666 VTAIL.n16 VSUBS 0.014026f
C667 VTAIL.n17 VSUBS 0.033152f
C668 VTAIL.n18 VSUBS 0.014851f
C669 VTAIL.n19 VSUBS 0.026102f
C670 VTAIL.n20 VSUBS 0.014026f
C671 VTAIL.n21 VSUBS 0.033152f
C672 VTAIL.n22 VSUBS 0.014851f
C673 VTAIL.n23 VSUBS 0.215124f
C674 VTAIL.t15 VSUBS 0.071509f
C675 VTAIL.n24 VSUBS 0.024864f
C676 VTAIL.n25 VSUBS 0.024939f
C677 VTAIL.n26 VSUBS 0.014026f
C678 VTAIL.n27 VSUBS 1.3751f
C679 VTAIL.n28 VSUBS 0.026102f
C680 VTAIL.n29 VSUBS 0.014026f
C681 VTAIL.n30 VSUBS 0.014851f
C682 VTAIL.n31 VSUBS 0.033152f
C683 VTAIL.n32 VSUBS 0.033152f
C684 VTAIL.n33 VSUBS 0.014851f
C685 VTAIL.n34 VSUBS 0.014026f
C686 VTAIL.n35 VSUBS 0.026102f
C687 VTAIL.n36 VSUBS 0.026102f
C688 VTAIL.n37 VSUBS 0.014026f
C689 VTAIL.n38 VSUBS 0.014851f
C690 VTAIL.n39 VSUBS 0.033152f
C691 VTAIL.n40 VSUBS 0.033152f
C692 VTAIL.n41 VSUBS 0.033152f
C693 VTAIL.n42 VSUBS 0.014851f
C694 VTAIL.n43 VSUBS 0.014026f
C695 VTAIL.n44 VSUBS 0.026102f
C696 VTAIL.n45 VSUBS 0.026102f
C697 VTAIL.n46 VSUBS 0.014026f
C698 VTAIL.n47 VSUBS 0.014438f
C699 VTAIL.n48 VSUBS 0.014438f
C700 VTAIL.n49 VSUBS 0.033152f
C701 VTAIL.n50 VSUBS 0.033152f
C702 VTAIL.n51 VSUBS 0.014851f
C703 VTAIL.n52 VSUBS 0.014026f
C704 VTAIL.n53 VSUBS 0.026102f
C705 VTAIL.n54 VSUBS 0.026102f
C706 VTAIL.n55 VSUBS 0.014026f
C707 VTAIL.n56 VSUBS 0.014851f
C708 VTAIL.n57 VSUBS 0.033152f
C709 VTAIL.n58 VSUBS 0.033152f
C710 VTAIL.n59 VSUBS 0.014851f
C711 VTAIL.n60 VSUBS 0.014026f
C712 VTAIL.n61 VSUBS 0.026102f
C713 VTAIL.n62 VSUBS 0.026102f
C714 VTAIL.n63 VSUBS 0.014026f
C715 VTAIL.n64 VSUBS 0.014851f
C716 VTAIL.n65 VSUBS 0.033152f
C717 VTAIL.n66 VSUBS 0.080263f
C718 VTAIL.n67 VSUBS 0.014851f
C719 VTAIL.n68 VSUBS 0.014026f
C720 VTAIL.n69 VSUBS 0.059263f
C721 VTAIL.n70 VSUBS 0.040331f
C722 VTAIL.n71 VSUBS 0.120658f
C723 VTAIL.n72 VSUBS 0.028682f
C724 VTAIL.n73 VSUBS 0.026102f
C725 VTAIL.n74 VSUBS 0.014026f
C726 VTAIL.n75 VSUBS 0.033152f
C727 VTAIL.n76 VSUBS 0.014851f
C728 VTAIL.n77 VSUBS 0.026102f
C729 VTAIL.n78 VSUBS 0.014026f
C730 VTAIL.n79 VSUBS 0.033152f
C731 VTAIL.n80 VSUBS 0.014851f
C732 VTAIL.n81 VSUBS 0.026102f
C733 VTAIL.n82 VSUBS 0.014026f
C734 VTAIL.n83 VSUBS 0.033152f
C735 VTAIL.n84 VSUBS 0.014851f
C736 VTAIL.n85 VSUBS 0.026102f
C737 VTAIL.n86 VSUBS 0.014026f
C738 VTAIL.n87 VSUBS 0.033152f
C739 VTAIL.n88 VSUBS 0.014851f
C740 VTAIL.n89 VSUBS 0.026102f
C741 VTAIL.n90 VSUBS 0.014026f
C742 VTAIL.n91 VSUBS 0.033152f
C743 VTAIL.n92 VSUBS 0.014851f
C744 VTAIL.n93 VSUBS 0.215124f
C745 VTAIL.t5 VSUBS 0.071509f
C746 VTAIL.n94 VSUBS 0.024864f
C747 VTAIL.n95 VSUBS 0.024939f
C748 VTAIL.n96 VSUBS 0.014026f
C749 VTAIL.n97 VSUBS 1.3751f
C750 VTAIL.n98 VSUBS 0.026102f
C751 VTAIL.n99 VSUBS 0.014026f
C752 VTAIL.n100 VSUBS 0.014851f
C753 VTAIL.n101 VSUBS 0.033152f
C754 VTAIL.n102 VSUBS 0.033152f
C755 VTAIL.n103 VSUBS 0.014851f
C756 VTAIL.n104 VSUBS 0.014026f
C757 VTAIL.n105 VSUBS 0.026102f
C758 VTAIL.n106 VSUBS 0.026102f
C759 VTAIL.n107 VSUBS 0.014026f
C760 VTAIL.n108 VSUBS 0.014851f
C761 VTAIL.n109 VSUBS 0.033152f
C762 VTAIL.n110 VSUBS 0.033152f
C763 VTAIL.n111 VSUBS 0.033152f
C764 VTAIL.n112 VSUBS 0.014851f
C765 VTAIL.n113 VSUBS 0.014026f
C766 VTAIL.n114 VSUBS 0.026102f
C767 VTAIL.n115 VSUBS 0.026102f
C768 VTAIL.n116 VSUBS 0.014026f
C769 VTAIL.n117 VSUBS 0.014438f
C770 VTAIL.n118 VSUBS 0.014438f
C771 VTAIL.n119 VSUBS 0.033152f
C772 VTAIL.n120 VSUBS 0.033152f
C773 VTAIL.n121 VSUBS 0.014851f
C774 VTAIL.n122 VSUBS 0.014026f
C775 VTAIL.n123 VSUBS 0.026102f
C776 VTAIL.n124 VSUBS 0.026102f
C777 VTAIL.n125 VSUBS 0.014026f
C778 VTAIL.n126 VSUBS 0.014851f
C779 VTAIL.n127 VSUBS 0.033152f
C780 VTAIL.n128 VSUBS 0.033152f
C781 VTAIL.n129 VSUBS 0.014851f
C782 VTAIL.n130 VSUBS 0.014026f
C783 VTAIL.n131 VSUBS 0.026102f
C784 VTAIL.n132 VSUBS 0.026102f
C785 VTAIL.n133 VSUBS 0.014026f
C786 VTAIL.n134 VSUBS 0.014851f
C787 VTAIL.n135 VSUBS 0.033152f
C788 VTAIL.n136 VSUBS 0.080263f
C789 VTAIL.n137 VSUBS 0.014851f
C790 VTAIL.n138 VSUBS 0.014026f
C791 VTAIL.n139 VSUBS 0.059263f
C792 VTAIL.n140 VSUBS 0.040331f
C793 VTAIL.n141 VSUBS 0.120658f
C794 VTAIL.t1 VSUBS 0.264224f
C795 VTAIL.t3 VSUBS 0.264224f
C796 VTAIL.n142 VSUBS 1.93357f
C797 VTAIL.n143 VSUBS 0.730404f
C798 VTAIL.n144 VSUBS 0.028682f
C799 VTAIL.n145 VSUBS 0.026102f
C800 VTAIL.n146 VSUBS 0.014026f
C801 VTAIL.n147 VSUBS 0.033152f
C802 VTAIL.n148 VSUBS 0.014851f
C803 VTAIL.n149 VSUBS 0.026102f
C804 VTAIL.n150 VSUBS 0.014026f
C805 VTAIL.n151 VSUBS 0.033152f
C806 VTAIL.n152 VSUBS 0.014851f
C807 VTAIL.n153 VSUBS 0.026102f
C808 VTAIL.n154 VSUBS 0.014026f
C809 VTAIL.n155 VSUBS 0.033152f
C810 VTAIL.n156 VSUBS 0.014851f
C811 VTAIL.n157 VSUBS 0.026102f
C812 VTAIL.n158 VSUBS 0.014026f
C813 VTAIL.n159 VSUBS 0.033152f
C814 VTAIL.n160 VSUBS 0.014851f
C815 VTAIL.n161 VSUBS 0.026102f
C816 VTAIL.n162 VSUBS 0.014026f
C817 VTAIL.n163 VSUBS 0.033152f
C818 VTAIL.n164 VSUBS 0.014851f
C819 VTAIL.n165 VSUBS 0.215124f
C820 VTAIL.t4 VSUBS 0.071509f
C821 VTAIL.n166 VSUBS 0.024864f
C822 VTAIL.n167 VSUBS 0.024939f
C823 VTAIL.n168 VSUBS 0.014026f
C824 VTAIL.n169 VSUBS 1.3751f
C825 VTAIL.n170 VSUBS 0.026102f
C826 VTAIL.n171 VSUBS 0.014026f
C827 VTAIL.n172 VSUBS 0.014851f
C828 VTAIL.n173 VSUBS 0.033152f
C829 VTAIL.n174 VSUBS 0.033152f
C830 VTAIL.n175 VSUBS 0.014851f
C831 VTAIL.n176 VSUBS 0.014026f
C832 VTAIL.n177 VSUBS 0.026102f
C833 VTAIL.n178 VSUBS 0.026102f
C834 VTAIL.n179 VSUBS 0.014026f
C835 VTAIL.n180 VSUBS 0.014851f
C836 VTAIL.n181 VSUBS 0.033152f
C837 VTAIL.n182 VSUBS 0.033152f
C838 VTAIL.n183 VSUBS 0.033152f
C839 VTAIL.n184 VSUBS 0.014851f
C840 VTAIL.n185 VSUBS 0.014026f
C841 VTAIL.n186 VSUBS 0.026102f
C842 VTAIL.n187 VSUBS 0.026102f
C843 VTAIL.n188 VSUBS 0.014026f
C844 VTAIL.n189 VSUBS 0.014438f
C845 VTAIL.n190 VSUBS 0.014438f
C846 VTAIL.n191 VSUBS 0.033152f
C847 VTAIL.n192 VSUBS 0.033152f
C848 VTAIL.n193 VSUBS 0.014851f
C849 VTAIL.n194 VSUBS 0.014026f
C850 VTAIL.n195 VSUBS 0.026102f
C851 VTAIL.n196 VSUBS 0.026102f
C852 VTAIL.n197 VSUBS 0.014026f
C853 VTAIL.n198 VSUBS 0.014851f
C854 VTAIL.n199 VSUBS 0.033152f
C855 VTAIL.n200 VSUBS 0.033152f
C856 VTAIL.n201 VSUBS 0.014851f
C857 VTAIL.n202 VSUBS 0.014026f
C858 VTAIL.n203 VSUBS 0.026102f
C859 VTAIL.n204 VSUBS 0.026102f
C860 VTAIL.n205 VSUBS 0.014026f
C861 VTAIL.n206 VSUBS 0.014851f
C862 VTAIL.n207 VSUBS 0.033152f
C863 VTAIL.n208 VSUBS 0.080263f
C864 VTAIL.n209 VSUBS 0.014851f
C865 VTAIL.n210 VSUBS 0.014026f
C866 VTAIL.n211 VSUBS 0.059263f
C867 VTAIL.n212 VSUBS 0.040331f
C868 VTAIL.n213 VSUBS 1.42394f
C869 VTAIL.n214 VSUBS 0.028682f
C870 VTAIL.n215 VSUBS 0.026102f
C871 VTAIL.n216 VSUBS 0.014026f
C872 VTAIL.n217 VSUBS 0.033152f
C873 VTAIL.n218 VSUBS 0.014851f
C874 VTAIL.n219 VSUBS 0.026102f
C875 VTAIL.n220 VSUBS 0.014026f
C876 VTAIL.n221 VSUBS 0.033152f
C877 VTAIL.n222 VSUBS 0.014851f
C878 VTAIL.n223 VSUBS 0.026102f
C879 VTAIL.n224 VSUBS 0.014026f
C880 VTAIL.n225 VSUBS 0.033152f
C881 VTAIL.n226 VSUBS 0.014851f
C882 VTAIL.n227 VSUBS 0.026102f
C883 VTAIL.n228 VSUBS 0.014026f
C884 VTAIL.n229 VSUBS 0.033152f
C885 VTAIL.n230 VSUBS 0.033152f
C886 VTAIL.n231 VSUBS 0.014851f
C887 VTAIL.n232 VSUBS 0.026102f
C888 VTAIL.n233 VSUBS 0.014026f
C889 VTAIL.n234 VSUBS 0.033152f
C890 VTAIL.n235 VSUBS 0.014851f
C891 VTAIL.n236 VSUBS 0.215124f
C892 VTAIL.t11 VSUBS 0.071509f
C893 VTAIL.n237 VSUBS 0.024864f
C894 VTAIL.n238 VSUBS 0.024939f
C895 VTAIL.n239 VSUBS 0.014026f
C896 VTAIL.n240 VSUBS 1.3751f
C897 VTAIL.n241 VSUBS 0.026102f
C898 VTAIL.n242 VSUBS 0.014026f
C899 VTAIL.n243 VSUBS 0.014851f
C900 VTAIL.n244 VSUBS 0.033152f
C901 VTAIL.n245 VSUBS 0.033152f
C902 VTAIL.n246 VSUBS 0.014851f
C903 VTAIL.n247 VSUBS 0.014026f
C904 VTAIL.n248 VSUBS 0.026102f
C905 VTAIL.n249 VSUBS 0.026102f
C906 VTAIL.n250 VSUBS 0.014026f
C907 VTAIL.n251 VSUBS 0.014851f
C908 VTAIL.n252 VSUBS 0.033152f
C909 VTAIL.n253 VSUBS 0.033152f
C910 VTAIL.n254 VSUBS 0.014851f
C911 VTAIL.n255 VSUBS 0.014026f
C912 VTAIL.n256 VSUBS 0.026102f
C913 VTAIL.n257 VSUBS 0.026102f
C914 VTAIL.n258 VSUBS 0.014026f
C915 VTAIL.n259 VSUBS 0.014438f
C916 VTAIL.n260 VSUBS 0.014438f
C917 VTAIL.n261 VSUBS 0.033152f
C918 VTAIL.n262 VSUBS 0.033152f
C919 VTAIL.n263 VSUBS 0.014851f
C920 VTAIL.n264 VSUBS 0.014026f
C921 VTAIL.n265 VSUBS 0.026102f
C922 VTAIL.n266 VSUBS 0.026102f
C923 VTAIL.n267 VSUBS 0.014026f
C924 VTAIL.n268 VSUBS 0.014851f
C925 VTAIL.n269 VSUBS 0.033152f
C926 VTAIL.n270 VSUBS 0.033152f
C927 VTAIL.n271 VSUBS 0.014851f
C928 VTAIL.n272 VSUBS 0.014026f
C929 VTAIL.n273 VSUBS 0.026102f
C930 VTAIL.n274 VSUBS 0.026102f
C931 VTAIL.n275 VSUBS 0.014026f
C932 VTAIL.n276 VSUBS 0.014851f
C933 VTAIL.n277 VSUBS 0.033152f
C934 VTAIL.n278 VSUBS 0.080263f
C935 VTAIL.n279 VSUBS 0.014851f
C936 VTAIL.n280 VSUBS 0.014026f
C937 VTAIL.n281 VSUBS 0.059263f
C938 VTAIL.n282 VSUBS 0.040331f
C939 VTAIL.n283 VSUBS 1.42394f
C940 VTAIL.t12 VSUBS 0.264224f
C941 VTAIL.t10 VSUBS 0.264224f
C942 VTAIL.n284 VSUBS 1.93358f
C943 VTAIL.n285 VSUBS 0.730394f
C944 VTAIL.n286 VSUBS 0.028682f
C945 VTAIL.n287 VSUBS 0.026102f
C946 VTAIL.n288 VSUBS 0.014026f
C947 VTAIL.n289 VSUBS 0.033152f
C948 VTAIL.n290 VSUBS 0.014851f
C949 VTAIL.n291 VSUBS 0.026102f
C950 VTAIL.n292 VSUBS 0.014026f
C951 VTAIL.n293 VSUBS 0.033152f
C952 VTAIL.n294 VSUBS 0.014851f
C953 VTAIL.n295 VSUBS 0.026102f
C954 VTAIL.n296 VSUBS 0.014026f
C955 VTAIL.n297 VSUBS 0.033152f
C956 VTAIL.n298 VSUBS 0.014851f
C957 VTAIL.n299 VSUBS 0.026102f
C958 VTAIL.n300 VSUBS 0.014026f
C959 VTAIL.n301 VSUBS 0.033152f
C960 VTAIL.n302 VSUBS 0.033152f
C961 VTAIL.n303 VSUBS 0.014851f
C962 VTAIL.n304 VSUBS 0.026102f
C963 VTAIL.n305 VSUBS 0.014026f
C964 VTAIL.n306 VSUBS 0.033152f
C965 VTAIL.n307 VSUBS 0.014851f
C966 VTAIL.n308 VSUBS 0.215124f
C967 VTAIL.t13 VSUBS 0.071509f
C968 VTAIL.n309 VSUBS 0.024864f
C969 VTAIL.n310 VSUBS 0.024939f
C970 VTAIL.n311 VSUBS 0.014026f
C971 VTAIL.n312 VSUBS 1.3751f
C972 VTAIL.n313 VSUBS 0.026102f
C973 VTAIL.n314 VSUBS 0.014026f
C974 VTAIL.n315 VSUBS 0.014851f
C975 VTAIL.n316 VSUBS 0.033152f
C976 VTAIL.n317 VSUBS 0.033152f
C977 VTAIL.n318 VSUBS 0.014851f
C978 VTAIL.n319 VSUBS 0.014026f
C979 VTAIL.n320 VSUBS 0.026102f
C980 VTAIL.n321 VSUBS 0.026102f
C981 VTAIL.n322 VSUBS 0.014026f
C982 VTAIL.n323 VSUBS 0.014851f
C983 VTAIL.n324 VSUBS 0.033152f
C984 VTAIL.n325 VSUBS 0.033152f
C985 VTAIL.n326 VSUBS 0.014851f
C986 VTAIL.n327 VSUBS 0.014026f
C987 VTAIL.n328 VSUBS 0.026102f
C988 VTAIL.n329 VSUBS 0.026102f
C989 VTAIL.n330 VSUBS 0.014026f
C990 VTAIL.n331 VSUBS 0.014438f
C991 VTAIL.n332 VSUBS 0.014438f
C992 VTAIL.n333 VSUBS 0.033152f
C993 VTAIL.n334 VSUBS 0.033152f
C994 VTAIL.n335 VSUBS 0.014851f
C995 VTAIL.n336 VSUBS 0.014026f
C996 VTAIL.n337 VSUBS 0.026102f
C997 VTAIL.n338 VSUBS 0.026102f
C998 VTAIL.n339 VSUBS 0.014026f
C999 VTAIL.n340 VSUBS 0.014851f
C1000 VTAIL.n341 VSUBS 0.033152f
C1001 VTAIL.n342 VSUBS 0.033152f
C1002 VTAIL.n343 VSUBS 0.014851f
C1003 VTAIL.n344 VSUBS 0.014026f
C1004 VTAIL.n345 VSUBS 0.026102f
C1005 VTAIL.n346 VSUBS 0.026102f
C1006 VTAIL.n347 VSUBS 0.014026f
C1007 VTAIL.n348 VSUBS 0.014851f
C1008 VTAIL.n349 VSUBS 0.033152f
C1009 VTAIL.n350 VSUBS 0.080263f
C1010 VTAIL.n351 VSUBS 0.014851f
C1011 VTAIL.n352 VSUBS 0.014026f
C1012 VTAIL.n353 VSUBS 0.059263f
C1013 VTAIL.n354 VSUBS 0.040331f
C1014 VTAIL.n355 VSUBS 0.120658f
C1015 VTAIL.n356 VSUBS 0.028682f
C1016 VTAIL.n357 VSUBS 0.026102f
C1017 VTAIL.n358 VSUBS 0.014026f
C1018 VTAIL.n359 VSUBS 0.033152f
C1019 VTAIL.n360 VSUBS 0.014851f
C1020 VTAIL.n361 VSUBS 0.026102f
C1021 VTAIL.n362 VSUBS 0.014026f
C1022 VTAIL.n363 VSUBS 0.033152f
C1023 VTAIL.n364 VSUBS 0.014851f
C1024 VTAIL.n365 VSUBS 0.026102f
C1025 VTAIL.n366 VSUBS 0.014026f
C1026 VTAIL.n367 VSUBS 0.033152f
C1027 VTAIL.n368 VSUBS 0.014851f
C1028 VTAIL.n369 VSUBS 0.026102f
C1029 VTAIL.n370 VSUBS 0.014026f
C1030 VTAIL.n371 VSUBS 0.033152f
C1031 VTAIL.n372 VSUBS 0.033152f
C1032 VTAIL.n373 VSUBS 0.014851f
C1033 VTAIL.n374 VSUBS 0.026102f
C1034 VTAIL.n375 VSUBS 0.014026f
C1035 VTAIL.n376 VSUBS 0.033152f
C1036 VTAIL.n377 VSUBS 0.014851f
C1037 VTAIL.n378 VSUBS 0.215124f
C1038 VTAIL.t2 VSUBS 0.071509f
C1039 VTAIL.n379 VSUBS 0.024864f
C1040 VTAIL.n380 VSUBS 0.024939f
C1041 VTAIL.n381 VSUBS 0.014026f
C1042 VTAIL.n382 VSUBS 1.3751f
C1043 VTAIL.n383 VSUBS 0.026102f
C1044 VTAIL.n384 VSUBS 0.014026f
C1045 VTAIL.n385 VSUBS 0.014851f
C1046 VTAIL.n386 VSUBS 0.033152f
C1047 VTAIL.n387 VSUBS 0.033152f
C1048 VTAIL.n388 VSUBS 0.014851f
C1049 VTAIL.n389 VSUBS 0.014026f
C1050 VTAIL.n390 VSUBS 0.026102f
C1051 VTAIL.n391 VSUBS 0.026102f
C1052 VTAIL.n392 VSUBS 0.014026f
C1053 VTAIL.n393 VSUBS 0.014851f
C1054 VTAIL.n394 VSUBS 0.033152f
C1055 VTAIL.n395 VSUBS 0.033152f
C1056 VTAIL.n396 VSUBS 0.014851f
C1057 VTAIL.n397 VSUBS 0.014026f
C1058 VTAIL.n398 VSUBS 0.026102f
C1059 VTAIL.n399 VSUBS 0.026102f
C1060 VTAIL.n400 VSUBS 0.014026f
C1061 VTAIL.n401 VSUBS 0.014438f
C1062 VTAIL.n402 VSUBS 0.014438f
C1063 VTAIL.n403 VSUBS 0.033152f
C1064 VTAIL.n404 VSUBS 0.033152f
C1065 VTAIL.n405 VSUBS 0.014851f
C1066 VTAIL.n406 VSUBS 0.014026f
C1067 VTAIL.n407 VSUBS 0.026102f
C1068 VTAIL.n408 VSUBS 0.026102f
C1069 VTAIL.n409 VSUBS 0.014026f
C1070 VTAIL.n410 VSUBS 0.014851f
C1071 VTAIL.n411 VSUBS 0.033152f
C1072 VTAIL.n412 VSUBS 0.033152f
C1073 VTAIL.n413 VSUBS 0.014851f
C1074 VTAIL.n414 VSUBS 0.014026f
C1075 VTAIL.n415 VSUBS 0.026102f
C1076 VTAIL.n416 VSUBS 0.026102f
C1077 VTAIL.n417 VSUBS 0.014026f
C1078 VTAIL.n418 VSUBS 0.014851f
C1079 VTAIL.n419 VSUBS 0.033152f
C1080 VTAIL.n420 VSUBS 0.080263f
C1081 VTAIL.n421 VSUBS 0.014851f
C1082 VTAIL.n422 VSUBS 0.014026f
C1083 VTAIL.n423 VSUBS 0.059263f
C1084 VTAIL.n424 VSUBS 0.040331f
C1085 VTAIL.n425 VSUBS 0.120658f
C1086 VTAIL.t0 VSUBS 0.264224f
C1087 VTAIL.t6 VSUBS 0.264224f
C1088 VTAIL.n426 VSUBS 1.93358f
C1089 VTAIL.n427 VSUBS 0.730394f
C1090 VTAIL.n428 VSUBS 0.028682f
C1091 VTAIL.n429 VSUBS 0.026102f
C1092 VTAIL.n430 VSUBS 0.014026f
C1093 VTAIL.n431 VSUBS 0.033152f
C1094 VTAIL.n432 VSUBS 0.014851f
C1095 VTAIL.n433 VSUBS 0.026102f
C1096 VTAIL.n434 VSUBS 0.014026f
C1097 VTAIL.n435 VSUBS 0.033152f
C1098 VTAIL.n436 VSUBS 0.014851f
C1099 VTAIL.n437 VSUBS 0.026102f
C1100 VTAIL.n438 VSUBS 0.014026f
C1101 VTAIL.n439 VSUBS 0.033152f
C1102 VTAIL.n440 VSUBS 0.014851f
C1103 VTAIL.n441 VSUBS 0.026102f
C1104 VTAIL.n442 VSUBS 0.014026f
C1105 VTAIL.n443 VSUBS 0.033152f
C1106 VTAIL.n444 VSUBS 0.033152f
C1107 VTAIL.n445 VSUBS 0.014851f
C1108 VTAIL.n446 VSUBS 0.026102f
C1109 VTAIL.n447 VSUBS 0.014026f
C1110 VTAIL.n448 VSUBS 0.033152f
C1111 VTAIL.n449 VSUBS 0.014851f
C1112 VTAIL.n450 VSUBS 0.215124f
C1113 VTAIL.t7 VSUBS 0.071509f
C1114 VTAIL.n451 VSUBS 0.024864f
C1115 VTAIL.n452 VSUBS 0.024939f
C1116 VTAIL.n453 VSUBS 0.014026f
C1117 VTAIL.n454 VSUBS 1.3751f
C1118 VTAIL.n455 VSUBS 0.026102f
C1119 VTAIL.n456 VSUBS 0.014026f
C1120 VTAIL.n457 VSUBS 0.014851f
C1121 VTAIL.n458 VSUBS 0.033152f
C1122 VTAIL.n459 VSUBS 0.033152f
C1123 VTAIL.n460 VSUBS 0.014851f
C1124 VTAIL.n461 VSUBS 0.014026f
C1125 VTAIL.n462 VSUBS 0.026102f
C1126 VTAIL.n463 VSUBS 0.026102f
C1127 VTAIL.n464 VSUBS 0.014026f
C1128 VTAIL.n465 VSUBS 0.014851f
C1129 VTAIL.n466 VSUBS 0.033152f
C1130 VTAIL.n467 VSUBS 0.033152f
C1131 VTAIL.n468 VSUBS 0.014851f
C1132 VTAIL.n469 VSUBS 0.014026f
C1133 VTAIL.n470 VSUBS 0.026102f
C1134 VTAIL.n471 VSUBS 0.026102f
C1135 VTAIL.n472 VSUBS 0.014026f
C1136 VTAIL.n473 VSUBS 0.014438f
C1137 VTAIL.n474 VSUBS 0.014438f
C1138 VTAIL.n475 VSUBS 0.033152f
C1139 VTAIL.n476 VSUBS 0.033152f
C1140 VTAIL.n477 VSUBS 0.014851f
C1141 VTAIL.n478 VSUBS 0.014026f
C1142 VTAIL.n479 VSUBS 0.026102f
C1143 VTAIL.n480 VSUBS 0.026102f
C1144 VTAIL.n481 VSUBS 0.014026f
C1145 VTAIL.n482 VSUBS 0.014851f
C1146 VTAIL.n483 VSUBS 0.033152f
C1147 VTAIL.n484 VSUBS 0.033152f
C1148 VTAIL.n485 VSUBS 0.014851f
C1149 VTAIL.n486 VSUBS 0.014026f
C1150 VTAIL.n487 VSUBS 0.026102f
C1151 VTAIL.n488 VSUBS 0.026102f
C1152 VTAIL.n489 VSUBS 0.014026f
C1153 VTAIL.n490 VSUBS 0.014851f
C1154 VTAIL.n491 VSUBS 0.033152f
C1155 VTAIL.n492 VSUBS 0.080263f
C1156 VTAIL.n493 VSUBS 0.014851f
C1157 VTAIL.n494 VSUBS 0.014026f
C1158 VTAIL.n495 VSUBS 0.059263f
C1159 VTAIL.n496 VSUBS 0.040331f
C1160 VTAIL.n497 VSUBS 1.42394f
C1161 VTAIL.n498 VSUBS 0.028682f
C1162 VTAIL.n499 VSUBS 0.026102f
C1163 VTAIL.n500 VSUBS 0.014026f
C1164 VTAIL.n501 VSUBS 0.033152f
C1165 VTAIL.n502 VSUBS 0.014851f
C1166 VTAIL.n503 VSUBS 0.026102f
C1167 VTAIL.n504 VSUBS 0.014026f
C1168 VTAIL.n505 VSUBS 0.033152f
C1169 VTAIL.n506 VSUBS 0.014851f
C1170 VTAIL.n507 VSUBS 0.026102f
C1171 VTAIL.n508 VSUBS 0.014026f
C1172 VTAIL.n509 VSUBS 0.033152f
C1173 VTAIL.n510 VSUBS 0.014851f
C1174 VTAIL.n511 VSUBS 0.026102f
C1175 VTAIL.n512 VSUBS 0.014026f
C1176 VTAIL.n513 VSUBS 0.033152f
C1177 VTAIL.n514 VSUBS 0.014851f
C1178 VTAIL.n515 VSUBS 0.026102f
C1179 VTAIL.n516 VSUBS 0.014026f
C1180 VTAIL.n517 VSUBS 0.033152f
C1181 VTAIL.n518 VSUBS 0.014851f
C1182 VTAIL.n519 VSUBS 0.215124f
C1183 VTAIL.t8 VSUBS 0.071509f
C1184 VTAIL.n520 VSUBS 0.024864f
C1185 VTAIL.n521 VSUBS 0.024939f
C1186 VTAIL.n522 VSUBS 0.014026f
C1187 VTAIL.n523 VSUBS 1.3751f
C1188 VTAIL.n524 VSUBS 0.026102f
C1189 VTAIL.n525 VSUBS 0.014026f
C1190 VTAIL.n526 VSUBS 0.014851f
C1191 VTAIL.n527 VSUBS 0.033152f
C1192 VTAIL.n528 VSUBS 0.033152f
C1193 VTAIL.n529 VSUBS 0.014851f
C1194 VTAIL.n530 VSUBS 0.014026f
C1195 VTAIL.n531 VSUBS 0.026102f
C1196 VTAIL.n532 VSUBS 0.026102f
C1197 VTAIL.n533 VSUBS 0.014026f
C1198 VTAIL.n534 VSUBS 0.014851f
C1199 VTAIL.n535 VSUBS 0.033152f
C1200 VTAIL.n536 VSUBS 0.033152f
C1201 VTAIL.n537 VSUBS 0.033152f
C1202 VTAIL.n538 VSUBS 0.014851f
C1203 VTAIL.n539 VSUBS 0.014026f
C1204 VTAIL.n540 VSUBS 0.026102f
C1205 VTAIL.n541 VSUBS 0.026102f
C1206 VTAIL.n542 VSUBS 0.014026f
C1207 VTAIL.n543 VSUBS 0.014438f
C1208 VTAIL.n544 VSUBS 0.014438f
C1209 VTAIL.n545 VSUBS 0.033152f
C1210 VTAIL.n546 VSUBS 0.033152f
C1211 VTAIL.n547 VSUBS 0.014851f
C1212 VTAIL.n548 VSUBS 0.014026f
C1213 VTAIL.n549 VSUBS 0.026102f
C1214 VTAIL.n550 VSUBS 0.026102f
C1215 VTAIL.n551 VSUBS 0.014026f
C1216 VTAIL.n552 VSUBS 0.014851f
C1217 VTAIL.n553 VSUBS 0.033152f
C1218 VTAIL.n554 VSUBS 0.033152f
C1219 VTAIL.n555 VSUBS 0.014851f
C1220 VTAIL.n556 VSUBS 0.014026f
C1221 VTAIL.n557 VSUBS 0.026102f
C1222 VTAIL.n558 VSUBS 0.026102f
C1223 VTAIL.n559 VSUBS 0.014026f
C1224 VTAIL.n560 VSUBS 0.014851f
C1225 VTAIL.n561 VSUBS 0.033152f
C1226 VTAIL.n562 VSUBS 0.080263f
C1227 VTAIL.n563 VSUBS 0.014851f
C1228 VTAIL.n564 VSUBS 0.014026f
C1229 VTAIL.n565 VSUBS 0.059263f
C1230 VTAIL.n566 VSUBS 0.040331f
C1231 VTAIL.n567 VSUBS 1.41905f
C1232 VDD2.t3 VSUBS 0.299079f
C1233 VDD2.t4 VSUBS 0.299079f
C1234 VDD2.n0 VSUBS 2.35875f
C1235 VDD2.t7 VSUBS 0.299079f
C1236 VDD2.t0 VSUBS 0.299079f
C1237 VDD2.n1 VSUBS 2.35875f
C1238 VDD2.n2 VSUBS 3.12164f
C1239 VDD2.t6 VSUBS 0.299079f
C1240 VDD2.t2 VSUBS 0.299079f
C1241 VDD2.n3 VSUBS 2.35599f
C1242 VDD2.n4 VSUBS 3.01667f
C1243 VDD2.t5 VSUBS 0.299079f
C1244 VDD2.t1 VSUBS 0.299079f
C1245 VDD2.n5 VSUBS 2.35871f
C1246 VN.n0 VSUBS 0.059623f
C1247 VN.t1 VSUBS 1.06628f
C1248 VN.n1 VSUBS 0.43197f
C1249 VN.t0 VSUBS 1.07849f
C1250 VN.n2 VSUBS 0.414143f
C1251 VN.n3 VSUBS 0.194956f
C1252 VN.n4 VSUBS 0.01353f
C1253 VN.t6 VSUBS 1.06628f
C1254 VN.n5 VSUBS 0.43197f
C1255 VN.t7 VSUBS 1.06628f
C1256 VN.n6 VSUBS 0.425904f
C1257 VN.n7 VSUBS 0.046205f
C1258 VN.n8 VSUBS 0.059623f
C1259 VN.t5 VSUBS 1.06628f
C1260 VN.n9 VSUBS 0.43197f
C1261 VN.t2 VSUBS 1.07849f
C1262 VN.n10 VSUBS 0.414143f
C1263 VN.n11 VSUBS 0.194956f
C1264 VN.n12 VSUBS 0.01353f
C1265 VN.t3 VSUBS 1.06628f
C1266 VN.n13 VSUBS 0.43197f
C1267 VN.t4 VSUBS 1.06628f
C1268 VN.n14 VSUBS 0.425904f
C1269 VN.n15 VSUBS 2.47213f
.ends

