* NGSPICE file created from diff_pair_sample_0961.ext - technology: sky130A

.subckt diff_pair_sample_0961 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VN.t0 VDD2.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9569 pd=12.19 as=1.9569 ps=12.19 w=11.86 l=2.28
X1 VTAIL.t19 VP.t0 VDD1.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=1.9569 pd=12.19 as=1.9569 ps=12.19 w=11.86 l=2.28
X2 VDD2.t1 VN.t1 VTAIL.t17 B.t8 sky130_fd_pr__nfet_01v8 ad=4.6254 pd=24.5 as=1.9569 ps=12.19 w=11.86 l=2.28
X3 VDD1.t8 VP.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=4.6254 pd=24.5 as=1.9569 ps=12.19 w=11.86 l=2.28
X4 VDD1.t7 VP.t2 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=4.6254 pd=24.5 as=1.9569 ps=12.19 w=11.86 l=2.28
X5 VDD2.t0 VN.t2 VTAIL.t16 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9569 pd=12.19 as=4.6254 ps=24.5 w=11.86 l=2.28
X6 VTAIL.t15 VN.t3 VDD2.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=1.9569 pd=12.19 as=1.9569 ps=12.19 w=11.86 l=2.28
X7 VDD1.t6 VP.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.9569 pd=12.19 as=1.9569 ps=12.19 w=11.86 l=2.28
X8 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=4.6254 pd=24.5 as=0 ps=0 w=11.86 l=2.28
X9 VDD2.t2 VN.t4 VTAIL.t14 B.t5 sky130_fd_pr__nfet_01v8 ad=1.9569 pd=12.19 as=1.9569 ps=12.19 w=11.86 l=2.28
X10 VDD1.t5 VP.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9569 pd=12.19 as=4.6254 ps=24.5 w=11.86 l=2.28
X11 VDD2.t5 VN.t5 VTAIL.t13 B.t4 sky130_fd_pr__nfet_01v8 ad=4.6254 pd=24.5 as=1.9569 ps=12.19 w=11.86 l=2.28
X12 VDD2.t4 VN.t6 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=1.9569 pd=12.19 as=1.9569 ps=12.19 w=11.86 l=2.28
X13 VDD1.t4 VP.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9569 pd=12.19 as=4.6254 ps=24.5 w=11.86 l=2.28
X14 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=4.6254 pd=24.5 as=0 ps=0 w=11.86 l=2.28
X15 VTAIL.t7 VP.t6 VDD1.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=1.9569 pd=12.19 as=1.9569 ps=12.19 w=11.86 l=2.28
X16 VDD2.t7 VN.t7 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9569 pd=12.19 as=4.6254 ps=24.5 w=11.86 l=2.28
X17 VTAIL.t10 VN.t8 VDD2.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=1.9569 pd=12.19 as=1.9569 ps=12.19 w=11.86 l=2.28
X18 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=4.6254 pd=24.5 as=0 ps=0 w=11.86 l=2.28
X19 VTAIL.t2 VP.t7 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.9569 pd=12.19 as=1.9569 ps=12.19 w=11.86 l=2.28
X20 VDD1.t1 VP.t8 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.9569 pd=12.19 as=1.9569 ps=12.19 w=11.86 l=2.28
X21 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.6254 pd=24.5 as=0 ps=0 w=11.86 l=2.28
X22 VTAIL.t9 VN.t9 VDD2.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=1.9569 pd=12.19 as=1.9569 ps=12.19 w=11.86 l=2.28
X23 VTAIL.t0 VP.t9 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9569 pd=12.19 as=1.9569 ps=12.19 w=11.86 l=2.28
R0 VN.n71 VN.n37 161.3
R1 VN.n70 VN.n69 161.3
R2 VN.n68 VN.n38 161.3
R3 VN.n67 VN.n66 161.3
R4 VN.n65 VN.n39 161.3
R5 VN.n63 VN.n62 161.3
R6 VN.n61 VN.n40 161.3
R7 VN.n60 VN.n59 161.3
R8 VN.n58 VN.n41 161.3
R9 VN.n57 VN.n56 161.3
R10 VN.n55 VN.n42 161.3
R11 VN.n54 VN.n53 161.3
R12 VN.n52 VN.n43 161.3
R13 VN.n51 VN.n50 161.3
R14 VN.n49 VN.n44 161.3
R15 VN.n48 VN.n47 161.3
R16 VN.n34 VN.n0 161.3
R17 VN.n33 VN.n32 161.3
R18 VN.n31 VN.n1 161.3
R19 VN.n30 VN.n29 161.3
R20 VN.n28 VN.n2 161.3
R21 VN.n26 VN.n25 161.3
R22 VN.n24 VN.n3 161.3
R23 VN.n23 VN.n22 161.3
R24 VN.n21 VN.n4 161.3
R25 VN.n20 VN.n19 161.3
R26 VN.n18 VN.n5 161.3
R27 VN.n17 VN.n16 161.3
R28 VN.n15 VN.n6 161.3
R29 VN.n14 VN.n13 161.3
R30 VN.n12 VN.n7 161.3
R31 VN.n11 VN.n10 161.3
R32 VN.n8 VN.t5 156.679
R33 VN.n45 VN.t7 156.679
R34 VN.n5 VN.t4 125.362
R35 VN.n9 VN.t3 125.362
R36 VN.n27 VN.t8 125.362
R37 VN.n35 VN.t2 125.362
R38 VN.n42 VN.t6 125.362
R39 VN.n46 VN.t9 125.362
R40 VN.n64 VN.t0 125.362
R41 VN.n72 VN.t1 125.362
R42 VN.n36 VN.n35 100.088
R43 VN.n73 VN.n72 100.088
R44 VN.n9 VN.n8 66.8721
R45 VN.n46 VN.n45 66.8721
R46 VN.n15 VN.n14 56.5617
R47 VN.n22 VN.n21 56.5617
R48 VN.n52 VN.n51 56.5617
R49 VN.n59 VN.n58 56.5617
R50 VN VN.n73 51.502
R51 VN.n29 VN.n1 48.8116
R52 VN.n66 VN.n38 48.8116
R53 VN.n33 VN.n1 32.3425
R54 VN.n70 VN.n38 32.3425
R55 VN.n10 VN.n7 24.5923
R56 VN.n14 VN.n7 24.5923
R57 VN.n16 VN.n15 24.5923
R58 VN.n16 VN.n5 24.5923
R59 VN.n20 VN.n5 24.5923
R60 VN.n21 VN.n20 24.5923
R61 VN.n22 VN.n3 24.5923
R62 VN.n26 VN.n3 24.5923
R63 VN.n29 VN.n28 24.5923
R64 VN.n34 VN.n33 24.5923
R65 VN.n51 VN.n44 24.5923
R66 VN.n47 VN.n44 24.5923
R67 VN.n58 VN.n57 24.5923
R68 VN.n57 VN.n42 24.5923
R69 VN.n53 VN.n42 24.5923
R70 VN.n53 VN.n52 24.5923
R71 VN.n66 VN.n65 24.5923
R72 VN.n63 VN.n40 24.5923
R73 VN.n59 VN.n40 24.5923
R74 VN.n71 VN.n70 24.5923
R75 VN.n28 VN.n27 19.1821
R76 VN.n65 VN.n64 19.1821
R77 VN.n35 VN.n34 10.8209
R78 VN.n72 VN.n71 10.8209
R79 VN.n48 VN.n45 9.89957
R80 VN.n11 VN.n8 9.89957
R81 VN.n10 VN.n9 5.4107
R82 VN.n27 VN.n26 5.4107
R83 VN.n47 VN.n46 5.4107
R84 VN.n64 VN.n63 5.4107
R85 VN.n73 VN.n37 0.278335
R86 VN.n36 VN.n0 0.278335
R87 VN.n69 VN.n37 0.189894
R88 VN.n69 VN.n68 0.189894
R89 VN.n68 VN.n67 0.189894
R90 VN.n67 VN.n39 0.189894
R91 VN.n62 VN.n39 0.189894
R92 VN.n62 VN.n61 0.189894
R93 VN.n61 VN.n60 0.189894
R94 VN.n60 VN.n41 0.189894
R95 VN.n56 VN.n41 0.189894
R96 VN.n56 VN.n55 0.189894
R97 VN.n55 VN.n54 0.189894
R98 VN.n54 VN.n43 0.189894
R99 VN.n50 VN.n43 0.189894
R100 VN.n50 VN.n49 0.189894
R101 VN.n49 VN.n48 0.189894
R102 VN.n12 VN.n11 0.189894
R103 VN.n13 VN.n12 0.189894
R104 VN.n13 VN.n6 0.189894
R105 VN.n17 VN.n6 0.189894
R106 VN.n18 VN.n17 0.189894
R107 VN.n19 VN.n18 0.189894
R108 VN.n19 VN.n4 0.189894
R109 VN.n23 VN.n4 0.189894
R110 VN.n24 VN.n23 0.189894
R111 VN.n25 VN.n24 0.189894
R112 VN.n25 VN.n2 0.189894
R113 VN.n30 VN.n2 0.189894
R114 VN.n31 VN.n30 0.189894
R115 VN.n32 VN.n31 0.189894
R116 VN.n32 VN.n0 0.189894
R117 VN VN.n36 0.153485
R118 VDD2.n1 VDD2.t5 67.8387
R119 VDD2.n4 VDD2.t1 65.5889
R120 VDD2.n3 VDD2.n2 65.5513
R121 VDD2 VDD2.n7 65.5486
R122 VDD2.n6 VDD2.n5 63.9194
R123 VDD2.n1 VDD2.n0 63.9192
R124 VDD2.n4 VDD2.n3 44.6269
R125 VDD2.n6 VDD2.n4 2.2505
R126 VDD2.n7 VDD2.t9 1.66998
R127 VDD2.n7 VDD2.t7 1.66998
R128 VDD2.n5 VDD2.t8 1.66998
R129 VDD2.n5 VDD2.t4 1.66998
R130 VDD2.n2 VDD2.t6 1.66998
R131 VDD2.n2 VDD2.t0 1.66998
R132 VDD2.n0 VDD2.t3 1.66998
R133 VDD2.n0 VDD2.t2 1.66998
R134 VDD2 VDD2.n6 0.62119
R135 VDD2.n3 VDD2.n1 0.507654
R136 VTAIL.n11 VTAIL.t11 48.9101
R137 VTAIL.n17 VTAIL.t16 48.9099
R138 VTAIL.n2 VTAIL.t1 48.9099
R139 VTAIL.n16 VTAIL.t3 48.9099
R140 VTAIL.n15 VTAIL.n14 47.2406
R141 VTAIL.n13 VTAIL.n12 47.2406
R142 VTAIL.n10 VTAIL.n9 47.2406
R143 VTAIL.n8 VTAIL.n7 47.2406
R144 VTAIL.n19 VTAIL.n18 47.2404
R145 VTAIL.n1 VTAIL.n0 47.2404
R146 VTAIL.n4 VTAIL.n3 47.2404
R147 VTAIL.n6 VTAIL.n5 47.2404
R148 VTAIL.n8 VTAIL.n6 27.091
R149 VTAIL.n17 VTAIL.n16 24.841
R150 VTAIL.n10 VTAIL.n8 2.2505
R151 VTAIL.n11 VTAIL.n10 2.2505
R152 VTAIL.n15 VTAIL.n13 2.2505
R153 VTAIL.n16 VTAIL.n15 2.2505
R154 VTAIL.n6 VTAIL.n4 2.2505
R155 VTAIL.n4 VTAIL.n2 2.2505
R156 VTAIL.n19 VTAIL.n17 2.2505
R157 VTAIL VTAIL.n1 1.74619
R158 VTAIL.n18 VTAIL.t14 1.66998
R159 VTAIL.n18 VTAIL.t10 1.66998
R160 VTAIL.n0 VTAIL.t13 1.66998
R161 VTAIL.n0 VTAIL.t15 1.66998
R162 VTAIL.n3 VTAIL.t6 1.66998
R163 VTAIL.n3 VTAIL.t2 1.66998
R164 VTAIL.n5 VTAIL.t8 1.66998
R165 VTAIL.n5 VTAIL.t0 1.66998
R166 VTAIL.n14 VTAIL.t5 1.66998
R167 VTAIL.n14 VTAIL.t19 1.66998
R168 VTAIL.n12 VTAIL.t4 1.66998
R169 VTAIL.n12 VTAIL.t7 1.66998
R170 VTAIL.n9 VTAIL.t12 1.66998
R171 VTAIL.n9 VTAIL.t9 1.66998
R172 VTAIL.n7 VTAIL.t17 1.66998
R173 VTAIL.n7 VTAIL.t18 1.66998
R174 VTAIL.n13 VTAIL.n11 1.59533
R175 VTAIL.n2 VTAIL.n1 1.59533
R176 VTAIL VTAIL.n19 0.50481
R177 B.n723 B.n722 585
R178 B.n725 B.n150 585
R179 B.n728 B.n727 585
R180 B.n729 B.n149 585
R181 B.n731 B.n730 585
R182 B.n733 B.n148 585
R183 B.n736 B.n735 585
R184 B.n737 B.n147 585
R185 B.n739 B.n738 585
R186 B.n741 B.n146 585
R187 B.n744 B.n743 585
R188 B.n745 B.n145 585
R189 B.n747 B.n746 585
R190 B.n749 B.n144 585
R191 B.n752 B.n751 585
R192 B.n753 B.n143 585
R193 B.n755 B.n754 585
R194 B.n757 B.n142 585
R195 B.n760 B.n759 585
R196 B.n761 B.n141 585
R197 B.n763 B.n762 585
R198 B.n765 B.n140 585
R199 B.n768 B.n767 585
R200 B.n769 B.n139 585
R201 B.n771 B.n770 585
R202 B.n773 B.n138 585
R203 B.n776 B.n775 585
R204 B.n777 B.n137 585
R205 B.n779 B.n778 585
R206 B.n781 B.n136 585
R207 B.n784 B.n783 585
R208 B.n785 B.n135 585
R209 B.n787 B.n786 585
R210 B.n789 B.n134 585
R211 B.n792 B.n791 585
R212 B.n793 B.n133 585
R213 B.n795 B.n794 585
R214 B.n797 B.n132 585
R215 B.n800 B.n799 585
R216 B.n801 B.n128 585
R217 B.n803 B.n802 585
R218 B.n805 B.n127 585
R219 B.n808 B.n807 585
R220 B.n809 B.n126 585
R221 B.n811 B.n810 585
R222 B.n813 B.n125 585
R223 B.n816 B.n815 585
R224 B.n817 B.n124 585
R225 B.n819 B.n818 585
R226 B.n821 B.n123 585
R227 B.n824 B.n823 585
R228 B.n826 B.n120 585
R229 B.n828 B.n827 585
R230 B.n830 B.n119 585
R231 B.n833 B.n832 585
R232 B.n834 B.n118 585
R233 B.n836 B.n835 585
R234 B.n838 B.n117 585
R235 B.n841 B.n840 585
R236 B.n842 B.n116 585
R237 B.n844 B.n843 585
R238 B.n846 B.n115 585
R239 B.n849 B.n848 585
R240 B.n850 B.n114 585
R241 B.n852 B.n851 585
R242 B.n854 B.n113 585
R243 B.n857 B.n856 585
R244 B.n858 B.n112 585
R245 B.n860 B.n859 585
R246 B.n862 B.n111 585
R247 B.n865 B.n864 585
R248 B.n866 B.n110 585
R249 B.n868 B.n867 585
R250 B.n870 B.n109 585
R251 B.n873 B.n872 585
R252 B.n874 B.n108 585
R253 B.n876 B.n875 585
R254 B.n878 B.n107 585
R255 B.n881 B.n880 585
R256 B.n882 B.n106 585
R257 B.n884 B.n883 585
R258 B.n886 B.n105 585
R259 B.n889 B.n888 585
R260 B.n890 B.n104 585
R261 B.n892 B.n891 585
R262 B.n894 B.n103 585
R263 B.n897 B.n896 585
R264 B.n898 B.n102 585
R265 B.n900 B.n899 585
R266 B.n902 B.n101 585
R267 B.n905 B.n904 585
R268 B.n906 B.n100 585
R269 B.n721 B.n98 585
R270 B.n909 B.n98 585
R271 B.n720 B.n97 585
R272 B.n910 B.n97 585
R273 B.n719 B.n96 585
R274 B.n911 B.n96 585
R275 B.n718 B.n717 585
R276 B.n717 B.n92 585
R277 B.n716 B.n91 585
R278 B.n917 B.n91 585
R279 B.n715 B.n90 585
R280 B.n918 B.n90 585
R281 B.n714 B.n89 585
R282 B.n919 B.n89 585
R283 B.n713 B.n712 585
R284 B.n712 B.n85 585
R285 B.n711 B.n84 585
R286 B.n925 B.n84 585
R287 B.n710 B.n83 585
R288 B.n926 B.n83 585
R289 B.n709 B.n82 585
R290 B.n927 B.n82 585
R291 B.n708 B.n707 585
R292 B.n707 B.n78 585
R293 B.n706 B.n77 585
R294 B.n933 B.n77 585
R295 B.n705 B.n76 585
R296 B.n934 B.n76 585
R297 B.n704 B.n75 585
R298 B.n935 B.n75 585
R299 B.n703 B.n702 585
R300 B.n702 B.n71 585
R301 B.n701 B.n70 585
R302 B.n941 B.n70 585
R303 B.n700 B.n69 585
R304 B.n942 B.n69 585
R305 B.n699 B.n68 585
R306 B.n943 B.n68 585
R307 B.n698 B.n697 585
R308 B.n697 B.n64 585
R309 B.n696 B.n63 585
R310 B.n949 B.n63 585
R311 B.n695 B.n62 585
R312 B.n950 B.n62 585
R313 B.n694 B.n61 585
R314 B.n951 B.n61 585
R315 B.n693 B.n692 585
R316 B.n692 B.n57 585
R317 B.n691 B.n56 585
R318 B.n957 B.n56 585
R319 B.n690 B.n55 585
R320 B.n958 B.n55 585
R321 B.n689 B.n54 585
R322 B.n959 B.n54 585
R323 B.n688 B.n687 585
R324 B.n687 B.n50 585
R325 B.n686 B.n49 585
R326 B.n965 B.n49 585
R327 B.n685 B.n48 585
R328 B.n966 B.n48 585
R329 B.n684 B.n47 585
R330 B.n967 B.n47 585
R331 B.n683 B.n682 585
R332 B.n682 B.n43 585
R333 B.n681 B.n42 585
R334 B.n973 B.n42 585
R335 B.n680 B.n41 585
R336 B.n974 B.n41 585
R337 B.n679 B.n40 585
R338 B.n975 B.n40 585
R339 B.n678 B.n677 585
R340 B.n677 B.n36 585
R341 B.n676 B.n35 585
R342 B.n981 B.n35 585
R343 B.n675 B.n34 585
R344 B.n982 B.n34 585
R345 B.n674 B.n33 585
R346 B.n983 B.n33 585
R347 B.n673 B.n672 585
R348 B.n672 B.n29 585
R349 B.n671 B.n28 585
R350 B.n989 B.n28 585
R351 B.n670 B.n27 585
R352 B.n990 B.n27 585
R353 B.n669 B.n26 585
R354 B.n991 B.n26 585
R355 B.n668 B.n667 585
R356 B.n667 B.n22 585
R357 B.n666 B.n21 585
R358 B.n997 B.n21 585
R359 B.n665 B.n20 585
R360 B.n998 B.n20 585
R361 B.n664 B.n19 585
R362 B.n999 B.n19 585
R363 B.n663 B.n662 585
R364 B.n662 B.n15 585
R365 B.n661 B.n14 585
R366 B.n1005 B.n14 585
R367 B.n660 B.n13 585
R368 B.n1006 B.n13 585
R369 B.n659 B.n12 585
R370 B.n1007 B.n12 585
R371 B.n658 B.n657 585
R372 B.n657 B.n8 585
R373 B.n656 B.n7 585
R374 B.n1013 B.n7 585
R375 B.n655 B.n6 585
R376 B.n1014 B.n6 585
R377 B.n654 B.n5 585
R378 B.n1015 B.n5 585
R379 B.n653 B.n652 585
R380 B.n652 B.n4 585
R381 B.n651 B.n151 585
R382 B.n651 B.n650 585
R383 B.n641 B.n152 585
R384 B.n153 B.n152 585
R385 B.n643 B.n642 585
R386 B.n644 B.n643 585
R387 B.n640 B.n158 585
R388 B.n158 B.n157 585
R389 B.n639 B.n638 585
R390 B.n638 B.n637 585
R391 B.n160 B.n159 585
R392 B.n161 B.n160 585
R393 B.n630 B.n629 585
R394 B.n631 B.n630 585
R395 B.n628 B.n166 585
R396 B.n166 B.n165 585
R397 B.n627 B.n626 585
R398 B.n626 B.n625 585
R399 B.n168 B.n167 585
R400 B.n169 B.n168 585
R401 B.n618 B.n617 585
R402 B.n619 B.n618 585
R403 B.n616 B.n174 585
R404 B.n174 B.n173 585
R405 B.n615 B.n614 585
R406 B.n614 B.n613 585
R407 B.n176 B.n175 585
R408 B.n177 B.n176 585
R409 B.n606 B.n605 585
R410 B.n607 B.n606 585
R411 B.n604 B.n182 585
R412 B.n182 B.n181 585
R413 B.n603 B.n602 585
R414 B.n602 B.n601 585
R415 B.n184 B.n183 585
R416 B.n185 B.n184 585
R417 B.n594 B.n593 585
R418 B.n595 B.n594 585
R419 B.n592 B.n189 585
R420 B.n193 B.n189 585
R421 B.n591 B.n590 585
R422 B.n590 B.n589 585
R423 B.n191 B.n190 585
R424 B.n192 B.n191 585
R425 B.n582 B.n581 585
R426 B.n583 B.n582 585
R427 B.n580 B.n198 585
R428 B.n198 B.n197 585
R429 B.n579 B.n578 585
R430 B.n578 B.n577 585
R431 B.n200 B.n199 585
R432 B.n201 B.n200 585
R433 B.n570 B.n569 585
R434 B.n571 B.n570 585
R435 B.n568 B.n205 585
R436 B.n209 B.n205 585
R437 B.n567 B.n566 585
R438 B.n566 B.n565 585
R439 B.n207 B.n206 585
R440 B.n208 B.n207 585
R441 B.n558 B.n557 585
R442 B.n559 B.n558 585
R443 B.n556 B.n214 585
R444 B.n214 B.n213 585
R445 B.n555 B.n554 585
R446 B.n554 B.n553 585
R447 B.n216 B.n215 585
R448 B.n217 B.n216 585
R449 B.n546 B.n545 585
R450 B.n547 B.n546 585
R451 B.n544 B.n221 585
R452 B.n225 B.n221 585
R453 B.n543 B.n542 585
R454 B.n542 B.n541 585
R455 B.n223 B.n222 585
R456 B.n224 B.n223 585
R457 B.n534 B.n533 585
R458 B.n535 B.n534 585
R459 B.n532 B.n230 585
R460 B.n230 B.n229 585
R461 B.n531 B.n530 585
R462 B.n530 B.n529 585
R463 B.n232 B.n231 585
R464 B.n233 B.n232 585
R465 B.n522 B.n521 585
R466 B.n523 B.n522 585
R467 B.n520 B.n238 585
R468 B.n238 B.n237 585
R469 B.n519 B.n518 585
R470 B.n518 B.n517 585
R471 B.n240 B.n239 585
R472 B.n241 B.n240 585
R473 B.n510 B.n509 585
R474 B.n511 B.n510 585
R475 B.n508 B.n246 585
R476 B.n246 B.n245 585
R477 B.n507 B.n506 585
R478 B.n506 B.n505 585
R479 B.n248 B.n247 585
R480 B.n249 B.n248 585
R481 B.n498 B.n497 585
R482 B.n499 B.n498 585
R483 B.n496 B.n254 585
R484 B.n254 B.n253 585
R485 B.n495 B.n494 585
R486 B.n494 B.n493 585
R487 B.n490 B.n258 585
R488 B.n489 B.n488 585
R489 B.n486 B.n259 585
R490 B.n486 B.n257 585
R491 B.n485 B.n484 585
R492 B.n483 B.n482 585
R493 B.n481 B.n261 585
R494 B.n479 B.n478 585
R495 B.n477 B.n262 585
R496 B.n476 B.n475 585
R497 B.n473 B.n263 585
R498 B.n471 B.n470 585
R499 B.n469 B.n264 585
R500 B.n468 B.n467 585
R501 B.n465 B.n265 585
R502 B.n463 B.n462 585
R503 B.n461 B.n266 585
R504 B.n460 B.n459 585
R505 B.n457 B.n267 585
R506 B.n455 B.n454 585
R507 B.n453 B.n268 585
R508 B.n452 B.n451 585
R509 B.n449 B.n269 585
R510 B.n447 B.n446 585
R511 B.n445 B.n270 585
R512 B.n444 B.n443 585
R513 B.n441 B.n271 585
R514 B.n439 B.n438 585
R515 B.n437 B.n272 585
R516 B.n436 B.n435 585
R517 B.n433 B.n273 585
R518 B.n431 B.n430 585
R519 B.n429 B.n274 585
R520 B.n428 B.n427 585
R521 B.n425 B.n275 585
R522 B.n423 B.n422 585
R523 B.n421 B.n276 585
R524 B.n420 B.n419 585
R525 B.n417 B.n277 585
R526 B.n415 B.n414 585
R527 B.n413 B.n278 585
R528 B.n412 B.n411 585
R529 B.n409 B.n408 585
R530 B.n407 B.n406 585
R531 B.n405 B.n283 585
R532 B.n403 B.n402 585
R533 B.n401 B.n284 585
R534 B.n400 B.n399 585
R535 B.n397 B.n285 585
R536 B.n395 B.n394 585
R537 B.n393 B.n286 585
R538 B.n392 B.n391 585
R539 B.n389 B.n388 585
R540 B.n387 B.n386 585
R541 B.n385 B.n291 585
R542 B.n383 B.n382 585
R543 B.n381 B.n292 585
R544 B.n380 B.n379 585
R545 B.n377 B.n293 585
R546 B.n375 B.n374 585
R547 B.n373 B.n294 585
R548 B.n372 B.n371 585
R549 B.n369 B.n295 585
R550 B.n367 B.n366 585
R551 B.n365 B.n296 585
R552 B.n364 B.n363 585
R553 B.n361 B.n297 585
R554 B.n359 B.n358 585
R555 B.n357 B.n298 585
R556 B.n356 B.n355 585
R557 B.n353 B.n299 585
R558 B.n351 B.n350 585
R559 B.n349 B.n300 585
R560 B.n348 B.n347 585
R561 B.n345 B.n301 585
R562 B.n343 B.n342 585
R563 B.n341 B.n302 585
R564 B.n340 B.n339 585
R565 B.n337 B.n303 585
R566 B.n335 B.n334 585
R567 B.n333 B.n304 585
R568 B.n332 B.n331 585
R569 B.n329 B.n305 585
R570 B.n327 B.n326 585
R571 B.n325 B.n306 585
R572 B.n324 B.n323 585
R573 B.n321 B.n307 585
R574 B.n319 B.n318 585
R575 B.n317 B.n308 585
R576 B.n316 B.n315 585
R577 B.n313 B.n309 585
R578 B.n311 B.n310 585
R579 B.n256 B.n255 585
R580 B.n257 B.n256 585
R581 B.n492 B.n491 585
R582 B.n493 B.n492 585
R583 B.n252 B.n251 585
R584 B.n253 B.n252 585
R585 B.n501 B.n500 585
R586 B.n500 B.n499 585
R587 B.n502 B.n250 585
R588 B.n250 B.n249 585
R589 B.n504 B.n503 585
R590 B.n505 B.n504 585
R591 B.n244 B.n243 585
R592 B.n245 B.n244 585
R593 B.n513 B.n512 585
R594 B.n512 B.n511 585
R595 B.n514 B.n242 585
R596 B.n242 B.n241 585
R597 B.n516 B.n515 585
R598 B.n517 B.n516 585
R599 B.n236 B.n235 585
R600 B.n237 B.n236 585
R601 B.n525 B.n524 585
R602 B.n524 B.n523 585
R603 B.n526 B.n234 585
R604 B.n234 B.n233 585
R605 B.n528 B.n527 585
R606 B.n529 B.n528 585
R607 B.n228 B.n227 585
R608 B.n229 B.n228 585
R609 B.n537 B.n536 585
R610 B.n536 B.n535 585
R611 B.n538 B.n226 585
R612 B.n226 B.n224 585
R613 B.n540 B.n539 585
R614 B.n541 B.n540 585
R615 B.n220 B.n219 585
R616 B.n225 B.n220 585
R617 B.n549 B.n548 585
R618 B.n548 B.n547 585
R619 B.n550 B.n218 585
R620 B.n218 B.n217 585
R621 B.n552 B.n551 585
R622 B.n553 B.n552 585
R623 B.n212 B.n211 585
R624 B.n213 B.n212 585
R625 B.n561 B.n560 585
R626 B.n560 B.n559 585
R627 B.n562 B.n210 585
R628 B.n210 B.n208 585
R629 B.n564 B.n563 585
R630 B.n565 B.n564 585
R631 B.n204 B.n203 585
R632 B.n209 B.n204 585
R633 B.n573 B.n572 585
R634 B.n572 B.n571 585
R635 B.n574 B.n202 585
R636 B.n202 B.n201 585
R637 B.n576 B.n575 585
R638 B.n577 B.n576 585
R639 B.n196 B.n195 585
R640 B.n197 B.n196 585
R641 B.n585 B.n584 585
R642 B.n584 B.n583 585
R643 B.n586 B.n194 585
R644 B.n194 B.n192 585
R645 B.n588 B.n587 585
R646 B.n589 B.n588 585
R647 B.n188 B.n187 585
R648 B.n193 B.n188 585
R649 B.n597 B.n596 585
R650 B.n596 B.n595 585
R651 B.n598 B.n186 585
R652 B.n186 B.n185 585
R653 B.n600 B.n599 585
R654 B.n601 B.n600 585
R655 B.n180 B.n179 585
R656 B.n181 B.n180 585
R657 B.n609 B.n608 585
R658 B.n608 B.n607 585
R659 B.n610 B.n178 585
R660 B.n178 B.n177 585
R661 B.n612 B.n611 585
R662 B.n613 B.n612 585
R663 B.n172 B.n171 585
R664 B.n173 B.n172 585
R665 B.n621 B.n620 585
R666 B.n620 B.n619 585
R667 B.n622 B.n170 585
R668 B.n170 B.n169 585
R669 B.n624 B.n623 585
R670 B.n625 B.n624 585
R671 B.n164 B.n163 585
R672 B.n165 B.n164 585
R673 B.n633 B.n632 585
R674 B.n632 B.n631 585
R675 B.n634 B.n162 585
R676 B.n162 B.n161 585
R677 B.n636 B.n635 585
R678 B.n637 B.n636 585
R679 B.n156 B.n155 585
R680 B.n157 B.n156 585
R681 B.n646 B.n645 585
R682 B.n645 B.n644 585
R683 B.n647 B.n154 585
R684 B.n154 B.n153 585
R685 B.n649 B.n648 585
R686 B.n650 B.n649 585
R687 B.n2 B.n0 585
R688 B.n4 B.n2 585
R689 B.n3 B.n1 585
R690 B.n1014 B.n3 585
R691 B.n1012 B.n1011 585
R692 B.n1013 B.n1012 585
R693 B.n1010 B.n9 585
R694 B.n9 B.n8 585
R695 B.n1009 B.n1008 585
R696 B.n1008 B.n1007 585
R697 B.n11 B.n10 585
R698 B.n1006 B.n11 585
R699 B.n1004 B.n1003 585
R700 B.n1005 B.n1004 585
R701 B.n1002 B.n16 585
R702 B.n16 B.n15 585
R703 B.n1001 B.n1000 585
R704 B.n1000 B.n999 585
R705 B.n18 B.n17 585
R706 B.n998 B.n18 585
R707 B.n996 B.n995 585
R708 B.n997 B.n996 585
R709 B.n994 B.n23 585
R710 B.n23 B.n22 585
R711 B.n993 B.n992 585
R712 B.n992 B.n991 585
R713 B.n25 B.n24 585
R714 B.n990 B.n25 585
R715 B.n988 B.n987 585
R716 B.n989 B.n988 585
R717 B.n986 B.n30 585
R718 B.n30 B.n29 585
R719 B.n985 B.n984 585
R720 B.n984 B.n983 585
R721 B.n32 B.n31 585
R722 B.n982 B.n32 585
R723 B.n980 B.n979 585
R724 B.n981 B.n980 585
R725 B.n978 B.n37 585
R726 B.n37 B.n36 585
R727 B.n977 B.n976 585
R728 B.n976 B.n975 585
R729 B.n39 B.n38 585
R730 B.n974 B.n39 585
R731 B.n972 B.n971 585
R732 B.n973 B.n972 585
R733 B.n970 B.n44 585
R734 B.n44 B.n43 585
R735 B.n969 B.n968 585
R736 B.n968 B.n967 585
R737 B.n46 B.n45 585
R738 B.n966 B.n46 585
R739 B.n964 B.n963 585
R740 B.n965 B.n964 585
R741 B.n962 B.n51 585
R742 B.n51 B.n50 585
R743 B.n961 B.n960 585
R744 B.n960 B.n959 585
R745 B.n53 B.n52 585
R746 B.n958 B.n53 585
R747 B.n956 B.n955 585
R748 B.n957 B.n956 585
R749 B.n954 B.n58 585
R750 B.n58 B.n57 585
R751 B.n953 B.n952 585
R752 B.n952 B.n951 585
R753 B.n60 B.n59 585
R754 B.n950 B.n60 585
R755 B.n948 B.n947 585
R756 B.n949 B.n948 585
R757 B.n946 B.n65 585
R758 B.n65 B.n64 585
R759 B.n945 B.n944 585
R760 B.n944 B.n943 585
R761 B.n67 B.n66 585
R762 B.n942 B.n67 585
R763 B.n940 B.n939 585
R764 B.n941 B.n940 585
R765 B.n938 B.n72 585
R766 B.n72 B.n71 585
R767 B.n937 B.n936 585
R768 B.n936 B.n935 585
R769 B.n74 B.n73 585
R770 B.n934 B.n74 585
R771 B.n932 B.n931 585
R772 B.n933 B.n932 585
R773 B.n930 B.n79 585
R774 B.n79 B.n78 585
R775 B.n929 B.n928 585
R776 B.n928 B.n927 585
R777 B.n81 B.n80 585
R778 B.n926 B.n81 585
R779 B.n924 B.n923 585
R780 B.n925 B.n924 585
R781 B.n922 B.n86 585
R782 B.n86 B.n85 585
R783 B.n921 B.n920 585
R784 B.n920 B.n919 585
R785 B.n88 B.n87 585
R786 B.n918 B.n88 585
R787 B.n916 B.n915 585
R788 B.n917 B.n916 585
R789 B.n914 B.n93 585
R790 B.n93 B.n92 585
R791 B.n913 B.n912 585
R792 B.n912 B.n911 585
R793 B.n95 B.n94 585
R794 B.n910 B.n95 585
R795 B.n908 B.n907 585
R796 B.n909 B.n908 585
R797 B.n1017 B.n1016 585
R798 B.n1016 B.n1015 585
R799 B.n492 B.n258 526.135
R800 B.n908 B.n100 526.135
R801 B.n494 B.n256 526.135
R802 B.n723 B.n98 526.135
R803 B.n287 B.t18 332.87
R804 B.n279 B.t10 332.87
R805 B.n121 B.t21 332.87
R806 B.n129 B.t14 332.87
R807 B.n724 B.n99 256.663
R808 B.n726 B.n99 256.663
R809 B.n732 B.n99 256.663
R810 B.n734 B.n99 256.663
R811 B.n740 B.n99 256.663
R812 B.n742 B.n99 256.663
R813 B.n748 B.n99 256.663
R814 B.n750 B.n99 256.663
R815 B.n756 B.n99 256.663
R816 B.n758 B.n99 256.663
R817 B.n764 B.n99 256.663
R818 B.n766 B.n99 256.663
R819 B.n772 B.n99 256.663
R820 B.n774 B.n99 256.663
R821 B.n780 B.n99 256.663
R822 B.n782 B.n99 256.663
R823 B.n788 B.n99 256.663
R824 B.n790 B.n99 256.663
R825 B.n796 B.n99 256.663
R826 B.n798 B.n99 256.663
R827 B.n804 B.n99 256.663
R828 B.n806 B.n99 256.663
R829 B.n812 B.n99 256.663
R830 B.n814 B.n99 256.663
R831 B.n820 B.n99 256.663
R832 B.n822 B.n99 256.663
R833 B.n829 B.n99 256.663
R834 B.n831 B.n99 256.663
R835 B.n837 B.n99 256.663
R836 B.n839 B.n99 256.663
R837 B.n845 B.n99 256.663
R838 B.n847 B.n99 256.663
R839 B.n853 B.n99 256.663
R840 B.n855 B.n99 256.663
R841 B.n861 B.n99 256.663
R842 B.n863 B.n99 256.663
R843 B.n869 B.n99 256.663
R844 B.n871 B.n99 256.663
R845 B.n877 B.n99 256.663
R846 B.n879 B.n99 256.663
R847 B.n885 B.n99 256.663
R848 B.n887 B.n99 256.663
R849 B.n893 B.n99 256.663
R850 B.n895 B.n99 256.663
R851 B.n901 B.n99 256.663
R852 B.n903 B.n99 256.663
R853 B.n487 B.n257 256.663
R854 B.n260 B.n257 256.663
R855 B.n480 B.n257 256.663
R856 B.n474 B.n257 256.663
R857 B.n472 B.n257 256.663
R858 B.n466 B.n257 256.663
R859 B.n464 B.n257 256.663
R860 B.n458 B.n257 256.663
R861 B.n456 B.n257 256.663
R862 B.n450 B.n257 256.663
R863 B.n448 B.n257 256.663
R864 B.n442 B.n257 256.663
R865 B.n440 B.n257 256.663
R866 B.n434 B.n257 256.663
R867 B.n432 B.n257 256.663
R868 B.n426 B.n257 256.663
R869 B.n424 B.n257 256.663
R870 B.n418 B.n257 256.663
R871 B.n416 B.n257 256.663
R872 B.n410 B.n257 256.663
R873 B.n282 B.n257 256.663
R874 B.n404 B.n257 256.663
R875 B.n398 B.n257 256.663
R876 B.n396 B.n257 256.663
R877 B.n390 B.n257 256.663
R878 B.n290 B.n257 256.663
R879 B.n384 B.n257 256.663
R880 B.n378 B.n257 256.663
R881 B.n376 B.n257 256.663
R882 B.n370 B.n257 256.663
R883 B.n368 B.n257 256.663
R884 B.n362 B.n257 256.663
R885 B.n360 B.n257 256.663
R886 B.n354 B.n257 256.663
R887 B.n352 B.n257 256.663
R888 B.n346 B.n257 256.663
R889 B.n344 B.n257 256.663
R890 B.n338 B.n257 256.663
R891 B.n336 B.n257 256.663
R892 B.n330 B.n257 256.663
R893 B.n328 B.n257 256.663
R894 B.n322 B.n257 256.663
R895 B.n320 B.n257 256.663
R896 B.n314 B.n257 256.663
R897 B.n312 B.n257 256.663
R898 B.n492 B.n252 163.367
R899 B.n500 B.n252 163.367
R900 B.n500 B.n250 163.367
R901 B.n504 B.n250 163.367
R902 B.n504 B.n244 163.367
R903 B.n512 B.n244 163.367
R904 B.n512 B.n242 163.367
R905 B.n516 B.n242 163.367
R906 B.n516 B.n236 163.367
R907 B.n524 B.n236 163.367
R908 B.n524 B.n234 163.367
R909 B.n528 B.n234 163.367
R910 B.n528 B.n228 163.367
R911 B.n536 B.n228 163.367
R912 B.n536 B.n226 163.367
R913 B.n540 B.n226 163.367
R914 B.n540 B.n220 163.367
R915 B.n548 B.n220 163.367
R916 B.n548 B.n218 163.367
R917 B.n552 B.n218 163.367
R918 B.n552 B.n212 163.367
R919 B.n560 B.n212 163.367
R920 B.n560 B.n210 163.367
R921 B.n564 B.n210 163.367
R922 B.n564 B.n204 163.367
R923 B.n572 B.n204 163.367
R924 B.n572 B.n202 163.367
R925 B.n576 B.n202 163.367
R926 B.n576 B.n196 163.367
R927 B.n584 B.n196 163.367
R928 B.n584 B.n194 163.367
R929 B.n588 B.n194 163.367
R930 B.n588 B.n188 163.367
R931 B.n596 B.n188 163.367
R932 B.n596 B.n186 163.367
R933 B.n600 B.n186 163.367
R934 B.n600 B.n180 163.367
R935 B.n608 B.n180 163.367
R936 B.n608 B.n178 163.367
R937 B.n612 B.n178 163.367
R938 B.n612 B.n172 163.367
R939 B.n620 B.n172 163.367
R940 B.n620 B.n170 163.367
R941 B.n624 B.n170 163.367
R942 B.n624 B.n164 163.367
R943 B.n632 B.n164 163.367
R944 B.n632 B.n162 163.367
R945 B.n636 B.n162 163.367
R946 B.n636 B.n156 163.367
R947 B.n645 B.n156 163.367
R948 B.n645 B.n154 163.367
R949 B.n649 B.n154 163.367
R950 B.n649 B.n2 163.367
R951 B.n1016 B.n2 163.367
R952 B.n1016 B.n3 163.367
R953 B.n1012 B.n3 163.367
R954 B.n1012 B.n9 163.367
R955 B.n1008 B.n9 163.367
R956 B.n1008 B.n11 163.367
R957 B.n1004 B.n11 163.367
R958 B.n1004 B.n16 163.367
R959 B.n1000 B.n16 163.367
R960 B.n1000 B.n18 163.367
R961 B.n996 B.n18 163.367
R962 B.n996 B.n23 163.367
R963 B.n992 B.n23 163.367
R964 B.n992 B.n25 163.367
R965 B.n988 B.n25 163.367
R966 B.n988 B.n30 163.367
R967 B.n984 B.n30 163.367
R968 B.n984 B.n32 163.367
R969 B.n980 B.n32 163.367
R970 B.n980 B.n37 163.367
R971 B.n976 B.n37 163.367
R972 B.n976 B.n39 163.367
R973 B.n972 B.n39 163.367
R974 B.n972 B.n44 163.367
R975 B.n968 B.n44 163.367
R976 B.n968 B.n46 163.367
R977 B.n964 B.n46 163.367
R978 B.n964 B.n51 163.367
R979 B.n960 B.n51 163.367
R980 B.n960 B.n53 163.367
R981 B.n956 B.n53 163.367
R982 B.n956 B.n58 163.367
R983 B.n952 B.n58 163.367
R984 B.n952 B.n60 163.367
R985 B.n948 B.n60 163.367
R986 B.n948 B.n65 163.367
R987 B.n944 B.n65 163.367
R988 B.n944 B.n67 163.367
R989 B.n940 B.n67 163.367
R990 B.n940 B.n72 163.367
R991 B.n936 B.n72 163.367
R992 B.n936 B.n74 163.367
R993 B.n932 B.n74 163.367
R994 B.n932 B.n79 163.367
R995 B.n928 B.n79 163.367
R996 B.n928 B.n81 163.367
R997 B.n924 B.n81 163.367
R998 B.n924 B.n86 163.367
R999 B.n920 B.n86 163.367
R1000 B.n920 B.n88 163.367
R1001 B.n916 B.n88 163.367
R1002 B.n916 B.n93 163.367
R1003 B.n912 B.n93 163.367
R1004 B.n912 B.n95 163.367
R1005 B.n908 B.n95 163.367
R1006 B.n488 B.n486 163.367
R1007 B.n486 B.n485 163.367
R1008 B.n482 B.n481 163.367
R1009 B.n479 B.n262 163.367
R1010 B.n475 B.n473 163.367
R1011 B.n471 B.n264 163.367
R1012 B.n467 B.n465 163.367
R1013 B.n463 B.n266 163.367
R1014 B.n459 B.n457 163.367
R1015 B.n455 B.n268 163.367
R1016 B.n451 B.n449 163.367
R1017 B.n447 B.n270 163.367
R1018 B.n443 B.n441 163.367
R1019 B.n439 B.n272 163.367
R1020 B.n435 B.n433 163.367
R1021 B.n431 B.n274 163.367
R1022 B.n427 B.n425 163.367
R1023 B.n423 B.n276 163.367
R1024 B.n419 B.n417 163.367
R1025 B.n415 B.n278 163.367
R1026 B.n411 B.n409 163.367
R1027 B.n406 B.n405 163.367
R1028 B.n403 B.n284 163.367
R1029 B.n399 B.n397 163.367
R1030 B.n395 B.n286 163.367
R1031 B.n391 B.n389 163.367
R1032 B.n386 B.n385 163.367
R1033 B.n383 B.n292 163.367
R1034 B.n379 B.n377 163.367
R1035 B.n375 B.n294 163.367
R1036 B.n371 B.n369 163.367
R1037 B.n367 B.n296 163.367
R1038 B.n363 B.n361 163.367
R1039 B.n359 B.n298 163.367
R1040 B.n355 B.n353 163.367
R1041 B.n351 B.n300 163.367
R1042 B.n347 B.n345 163.367
R1043 B.n343 B.n302 163.367
R1044 B.n339 B.n337 163.367
R1045 B.n335 B.n304 163.367
R1046 B.n331 B.n329 163.367
R1047 B.n327 B.n306 163.367
R1048 B.n323 B.n321 163.367
R1049 B.n319 B.n308 163.367
R1050 B.n315 B.n313 163.367
R1051 B.n311 B.n256 163.367
R1052 B.n494 B.n254 163.367
R1053 B.n498 B.n254 163.367
R1054 B.n498 B.n248 163.367
R1055 B.n506 B.n248 163.367
R1056 B.n506 B.n246 163.367
R1057 B.n510 B.n246 163.367
R1058 B.n510 B.n240 163.367
R1059 B.n518 B.n240 163.367
R1060 B.n518 B.n238 163.367
R1061 B.n522 B.n238 163.367
R1062 B.n522 B.n232 163.367
R1063 B.n530 B.n232 163.367
R1064 B.n530 B.n230 163.367
R1065 B.n534 B.n230 163.367
R1066 B.n534 B.n223 163.367
R1067 B.n542 B.n223 163.367
R1068 B.n542 B.n221 163.367
R1069 B.n546 B.n221 163.367
R1070 B.n546 B.n216 163.367
R1071 B.n554 B.n216 163.367
R1072 B.n554 B.n214 163.367
R1073 B.n558 B.n214 163.367
R1074 B.n558 B.n207 163.367
R1075 B.n566 B.n207 163.367
R1076 B.n566 B.n205 163.367
R1077 B.n570 B.n205 163.367
R1078 B.n570 B.n200 163.367
R1079 B.n578 B.n200 163.367
R1080 B.n578 B.n198 163.367
R1081 B.n582 B.n198 163.367
R1082 B.n582 B.n191 163.367
R1083 B.n590 B.n191 163.367
R1084 B.n590 B.n189 163.367
R1085 B.n594 B.n189 163.367
R1086 B.n594 B.n184 163.367
R1087 B.n602 B.n184 163.367
R1088 B.n602 B.n182 163.367
R1089 B.n606 B.n182 163.367
R1090 B.n606 B.n176 163.367
R1091 B.n614 B.n176 163.367
R1092 B.n614 B.n174 163.367
R1093 B.n618 B.n174 163.367
R1094 B.n618 B.n168 163.367
R1095 B.n626 B.n168 163.367
R1096 B.n626 B.n166 163.367
R1097 B.n630 B.n166 163.367
R1098 B.n630 B.n160 163.367
R1099 B.n638 B.n160 163.367
R1100 B.n638 B.n158 163.367
R1101 B.n643 B.n158 163.367
R1102 B.n643 B.n152 163.367
R1103 B.n651 B.n152 163.367
R1104 B.n652 B.n651 163.367
R1105 B.n652 B.n5 163.367
R1106 B.n6 B.n5 163.367
R1107 B.n7 B.n6 163.367
R1108 B.n657 B.n7 163.367
R1109 B.n657 B.n12 163.367
R1110 B.n13 B.n12 163.367
R1111 B.n14 B.n13 163.367
R1112 B.n662 B.n14 163.367
R1113 B.n662 B.n19 163.367
R1114 B.n20 B.n19 163.367
R1115 B.n21 B.n20 163.367
R1116 B.n667 B.n21 163.367
R1117 B.n667 B.n26 163.367
R1118 B.n27 B.n26 163.367
R1119 B.n28 B.n27 163.367
R1120 B.n672 B.n28 163.367
R1121 B.n672 B.n33 163.367
R1122 B.n34 B.n33 163.367
R1123 B.n35 B.n34 163.367
R1124 B.n677 B.n35 163.367
R1125 B.n677 B.n40 163.367
R1126 B.n41 B.n40 163.367
R1127 B.n42 B.n41 163.367
R1128 B.n682 B.n42 163.367
R1129 B.n682 B.n47 163.367
R1130 B.n48 B.n47 163.367
R1131 B.n49 B.n48 163.367
R1132 B.n687 B.n49 163.367
R1133 B.n687 B.n54 163.367
R1134 B.n55 B.n54 163.367
R1135 B.n56 B.n55 163.367
R1136 B.n692 B.n56 163.367
R1137 B.n692 B.n61 163.367
R1138 B.n62 B.n61 163.367
R1139 B.n63 B.n62 163.367
R1140 B.n697 B.n63 163.367
R1141 B.n697 B.n68 163.367
R1142 B.n69 B.n68 163.367
R1143 B.n70 B.n69 163.367
R1144 B.n702 B.n70 163.367
R1145 B.n702 B.n75 163.367
R1146 B.n76 B.n75 163.367
R1147 B.n77 B.n76 163.367
R1148 B.n707 B.n77 163.367
R1149 B.n707 B.n82 163.367
R1150 B.n83 B.n82 163.367
R1151 B.n84 B.n83 163.367
R1152 B.n712 B.n84 163.367
R1153 B.n712 B.n89 163.367
R1154 B.n90 B.n89 163.367
R1155 B.n91 B.n90 163.367
R1156 B.n717 B.n91 163.367
R1157 B.n717 B.n96 163.367
R1158 B.n97 B.n96 163.367
R1159 B.n98 B.n97 163.367
R1160 B.n904 B.n902 163.367
R1161 B.n900 B.n102 163.367
R1162 B.n896 B.n894 163.367
R1163 B.n892 B.n104 163.367
R1164 B.n888 B.n886 163.367
R1165 B.n884 B.n106 163.367
R1166 B.n880 B.n878 163.367
R1167 B.n876 B.n108 163.367
R1168 B.n872 B.n870 163.367
R1169 B.n868 B.n110 163.367
R1170 B.n864 B.n862 163.367
R1171 B.n860 B.n112 163.367
R1172 B.n856 B.n854 163.367
R1173 B.n852 B.n114 163.367
R1174 B.n848 B.n846 163.367
R1175 B.n844 B.n116 163.367
R1176 B.n840 B.n838 163.367
R1177 B.n836 B.n118 163.367
R1178 B.n832 B.n830 163.367
R1179 B.n828 B.n120 163.367
R1180 B.n823 B.n821 163.367
R1181 B.n819 B.n124 163.367
R1182 B.n815 B.n813 163.367
R1183 B.n811 B.n126 163.367
R1184 B.n807 B.n805 163.367
R1185 B.n803 B.n128 163.367
R1186 B.n799 B.n797 163.367
R1187 B.n795 B.n133 163.367
R1188 B.n791 B.n789 163.367
R1189 B.n787 B.n135 163.367
R1190 B.n783 B.n781 163.367
R1191 B.n779 B.n137 163.367
R1192 B.n775 B.n773 163.367
R1193 B.n771 B.n139 163.367
R1194 B.n767 B.n765 163.367
R1195 B.n763 B.n141 163.367
R1196 B.n759 B.n757 163.367
R1197 B.n755 B.n143 163.367
R1198 B.n751 B.n749 163.367
R1199 B.n747 B.n145 163.367
R1200 B.n743 B.n741 163.367
R1201 B.n739 B.n147 163.367
R1202 B.n735 B.n733 163.367
R1203 B.n731 B.n149 163.367
R1204 B.n727 B.n725 163.367
R1205 B.n287 B.t20 124.246
R1206 B.n129 B.t16 124.246
R1207 B.n279 B.t13 124.231
R1208 B.n121 B.t22 124.231
R1209 B.n493 B.n257 86.6652
R1210 B.n909 B.n99 86.6652
R1211 B.n288 B.t19 73.6271
R1212 B.n130 B.t17 73.6271
R1213 B.n280 B.t12 73.6123
R1214 B.n122 B.t23 73.6123
R1215 B.n487 B.n258 71.676
R1216 B.n485 B.n260 71.676
R1217 B.n481 B.n480 71.676
R1218 B.n474 B.n262 71.676
R1219 B.n473 B.n472 71.676
R1220 B.n466 B.n264 71.676
R1221 B.n465 B.n464 71.676
R1222 B.n458 B.n266 71.676
R1223 B.n457 B.n456 71.676
R1224 B.n450 B.n268 71.676
R1225 B.n449 B.n448 71.676
R1226 B.n442 B.n270 71.676
R1227 B.n441 B.n440 71.676
R1228 B.n434 B.n272 71.676
R1229 B.n433 B.n432 71.676
R1230 B.n426 B.n274 71.676
R1231 B.n425 B.n424 71.676
R1232 B.n418 B.n276 71.676
R1233 B.n417 B.n416 71.676
R1234 B.n410 B.n278 71.676
R1235 B.n409 B.n282 71.676
R1236 B.n405 B.n404 71.676
R1237 B.n398 B.n284 71.676
R1238 B.n397 B.n396 71.676
R1239 B.n390 B.n286 71.676
R1240 B.n389 B.n290 71.676
R1241 B.n385 B.n384 71.676
R1242 B.n378 B.n292 71.676
R1243 B.n377 B.n376 71.676
R1244 B.n370 B.n294 71.676
R1245 B.n369 B.n368 71.676
R1246 B.n362 B.n296 71.676
R1247 B.n361 B.n360 71.676
R1248 B.n354 B.n298 71.676
R1249 B.n353 B.n352 71.676
R1250 B.n346 B.n300 71.676
R1251 B.n345 B.n344 71.676
R1252 B.n338 B.n302 71.676
R1253 B.n337 B.n336 71.676
R1254 B.n330 B.n304 71.676
R1255 B.n329 B.n328 71.676
R1256 B.n322 B.n306 71.676
R1257 B.n321 B.n320 71.676
R1258 B.n314 B.n308 71.676
R1259 B.n313 B.n312 71.676
R1260 B.n903 B.n100 71.676
R1261 B.n902 B.n901 71.676
R1262 B.n895 B.n102 71.676
R1263 B.n894 B.n893 71.676
R1264 B.n887 B.n104 71.676
R1265 B.n886 B.n885 71.676
R1266 B.n879 B.n106 71.676
R1267 B.n878 B.n877 71.676
R1268 B.n871 B.n108 71.676
R1269 B.n870 B.n869 71.676
R1270 B.n863 B.n110 71.676
R1271 B.n862 B.n861 71.676
R1272 B.n855 B.n112 71.676
R1273 B.n854 B.n853 71.676
R1274 B.n847 B.n114 71.676
R1275 B.n846 B.n845 71.676
R1276 B.n839 B.n116 71.676
R1277 B.n838 B.n837 71.676
R1278 B.n831 B.n118 71.676
R1279 B.n830 B.n829 71.676
R1280 B.n822 B.n120 71.676
R1281 B.n821 B.n820 71.676
R1282 B.n814 B.n124 71.676
R1283 B.n813 B.n812 71.676
R1284 B.n806 B.n126 71.676
R1285 B.n805 B.n804 71.676
R1286 B.n798 B.n128 71.676
R1287 B.n797 B.n796 71.676
R1288 B.n790 B.n133 71.676
R1289 B.n789 B.n788 71.676
R1290 B.n782 B.n135 71.676
R1291 B.n781 B.n780 71.676
R1292 B.n774 B.n137 71.676
R1293 B.n773 B.n772 71.676
R1294 B.n766 B.n139 71.676
R1295 B.n765 B.n764 71.676
R1296 B.n758 B.n141 71.676
R1297 B.n757 B.n756 71.676
R1298 B.n750 B.n143 71.676
R1299 B.n749 B.n748 71.676
R1300 B.n742 B.n145 71.676
R1301 B.n741 B.n740 71.676
R1302 B.n734 B.n147 71.676
R1303 B.n733 B.n732 71.676
R1304 B.n726 B.n149 71.676
R1305 B.n725 B.n724 71.676
R1306 B.n724 B.n723 71.676
R1307 B.n727 B.n726 71.676
R1308 B.n732 B.n731 71.676
R1309 B.n735 B.n734 71.676
R1310 B.n740 B.n739 71.676
R1311 B.n743 B.n742 71.676
R1312 B.n748 B.n747 71.676
R1313 B.n751 B.n750 71.676
R1314 B.n756 B.n755 71.676
R1315 B.n759 B.n758 71.676
R1316 B.n764 B.n763 71.676
R1317 B.n767 B.n766 71.676
R1318 B.n772 B.n771 71.676
R1319 B.n775 B.n774 71.676
R1320 B.n780 B.n779 71.676
R1321 B.n783 B.n782 71.676
R1322 B.n788 B.n787 71.676
R1323 B.n791 B.n790 71.676
R1324 B.n796 B.n795 71.676
R1325 B.n799 B.n798 71.676
R1326 B.n804 B.n803 71.676
R1327 B.n807 B.n806 71.676
R1328 B.n812 B.n811 71.676
R1329 B.n815 B.n814 71.676
R1330 B.n820 B.n819 71.676
R1331 B.n823 B.n822 71.676
R1332 B.n829 B.n828 71.676
R1333 B.n832 B.n831 71.676
R1334 B.n837 B.n836 71.676
R1335 B.n840 B.n839 71.676
R1336 B.n845 B.n844 71.676
R1337 B.n848 B.n847 71.676
R1338 B.n853 B.n852 71.676
R1339 B.n856 B.n855 71.676
R1340 B.n861 B.n860 71.676
R1341 B.n864 B.n863 71.676
R1342 B.n869 B.n868 71.676
R1343 B.n872 B.n871 71.676
R1344 B.n877 B.n876 71.676
R1345 B.n880 B.n879 71.676
R1346 B.n885 B.n884 71.676
R1347 B.n888 B.n887 71.676
R1348 B.n893 B.n892 71.676
R1349 B.n896 B.n895 71.676
R1350 B.n901 B.n900 71.676
R1351 B.n904 B.n903 71.676
R1352 B.n488 B.n487 71.676
R1353 B.n482 B.n260 71.676
R1354 B.n480 B.n479 71.676
R1355 B.n475 B.n474 71.676
R1356 B.n472 B.n471 71.676
R1357 B.n467 B.n466 71.676
R1358 B.n464 B.n463 71.676
R1359 B.n459 B.n458 71.676
R1360 B.n456 B.n455 71.676
R1361 B.n451 B.n450 71.676
R1362 B.n448 B.n447 71.676
R1363 B.n443 B.n442 71.676
R1364 B.n440 B.n439 71.676
R1365 B.n435 B.n434 71.676
R1366 B.n432 B.n431 71.676
R1367 B.n427 B.n426 71.676
R1368 B.n424 B.n423 71.676
R1369 B.n419 B.n418 71.676
R1370 B.n416 B.n415 71.676
R1371 B.n411 B.n410 71.676
R1372 B.n406 B.n282 71.676
R1373 B.n404 B.n403 71.676
R1374 B.n399 B.n398 71.676
R1375 B.n396 B.n395 71.676
R1376 B.n391 B.n390 71.676
R1377 B.n386 B.n290 71.676
R1378 B.n384 B.n383 71.676
R1379 B.n379 B.n378 71.676
R1380 B.n376 B.n375 71.676
R1381 B.n371 B.n370 71.676
R1382 B.n368 B.n367 71.676
R1383 B.n363 B.n362 71.676
R1384 B.n360 B.n359 71.676
R1385 B.n355 B.n354 71.676
R1386 B.n352 B.n351 71.676
R1387 B.n347 B.n346 71.676
R1388 B.n344 B.n343 71.676
R1389 B.n339 B.n338 71.676
R1390 B.n336 B.n335 71.676
R1391 B.n331 B.n330 71.676
R1392 B.n328 B.n327 71.676
R1393 B.n323 B.n322 71.676
R1394 B.n320 B.n319 71.676
R1395 B.n315 B.n314 71.676
R1396 B.n312 B.n311 71.676
R1397 B.n289 B.n288 59.5399
R1398 B.n281 B.n280 59.5399
R1399 B.n825 B.n122 59.5399
R1400 B.n131 B.n130 59.5399
R1401 B.n288 B.n287 50.6187
R1402 B.n280 B.n279 50.6187
R1403 B.n122 B.n121 50.6187
R1404 B.n130 B.n129 50.6187
R1405 B.n493 B.n253 43.6538
R1406 B.n499 B.n253 43.6538
R1407 B.n499 B.n249 43.6538
R1408 B.n505 B.n249 43.6538
R1409 B.n505 B.n245 43.6538
R1410 B.n511 B.n245 43.6538
R1411 B.n517 B.n241 43.6538
R1412 B.n517 B.n237 43.6538
R1413 B.n523 B.n237 43.6538
R1414 B.n523 B.n233 43.6538
R1415 B.n529 B.n233 43.6538
R1416 B.n529 B.n229 43.6538
R1417 B.n535 B.n229 43.6538
R1418 B.n535 B.n224 43.6538
R1419 B.n541 B.n224 43.6538
R1420 B.n541 B.n225 43.6538
R1421 B.n547 B.n217 43.6538
R1422 B.n553 B.n217 43.6538
R1423 B.n553 B.n213 43.6538
R1424 B.n559 B.n213 43.6538
R1425 B.n559 B.n208 43.6538
R1426 B.n565 B.n208 43.6538
R1427 B.n565 B.n209 43.6538
R1428 B.n571 B.n201 43.6538
R1429 B.n577 B.n201 43.6538
R1430 B.n577 B.n197 43.6538
R1431 B.n583 B.n197 43.6538
R1432 B.n583 B.n192 43.6538
R1433 B.n589 B.n192 43.6538
R1434 B.n589 B.n193 43.6538
R1435 B.n595 B.n185 43.6538
R1436 B.n601 B.n185 43.6538
R1437 B.n601 B.n181 43.6538
R1438 B.n607 B.n181 43.6538
R1439 B.n607 B.n177 43.6538
R1440 B.n613 B.n177 43.6538
R1441 B.n619 B.n173 43.6538
R1442 B.n619 B.n169 43.6538
R1443 B.n625 B.n169 43.6538
R1444 B.n625 B.n165 43.6538
R1445 B.n631 B.n165 43.6538
R1446 B.n631 B.n161 43.6538
R1447 B.n637 B.n161 43.6538
R1448 B.n644 B.n157 43.6538
R1449 B.n644 B.n153 43.6538
R1450 B.n650 B.n153 43.6538
R1451 B.n650 B.n4 43.6538
R1452 B.n1015 B.n4 43.6538
R1453 B.n1015 B.n1014 43.6538
R1454 B.n1014 B.n1013 43.6538
R1455 B.n1013 B.n8 43.6538
R1456 B.n1007 B.n8 43.6538
R1457 B.n1007 B.n1006 43.6538
R1458 B.n1005 B.n15 43.6538
R1459 B.n999 B.n15 43.6538
R1460 B.n999 B.n998 43.6538
R1461 B.n998 B.n997 43.6538
R1462 B.n997 B.n22 43.6538
R1463 B.n991 B.n22 43.6538
R1464 B.n991 B.n990 43.6538
R1465 B.n989 B.n29 43.6538
R1466 B.n983 B.n29 43.6538
R1467 B.n983 B.n982 43.6538
R1468 B.n982 B.n981 43.6538
R1469 B.n981 B.n36 43.6538
R1470 B.n975 B.n36 43.6538
R1471 B.n974 B.n973 43.6538
R1472 B.n973 B.n43 43.6538
R1473 B.n967 B.n43 43.6538
R1474 B.n967 B.n966 43.6538
R1475 B.n966 B.n965 43.6538
R1476 B.n965 B.n50 43.6538
R1477 B.n959 B.n50 43.6538
R1478 B.n958 B.n957 43.6538
R1479 B.n957 B.n57 43.6538
R1480 B.n951 B.n57 43.6538
R1481 B.n951 B.n950 43.6538
R1482 B.n950 B.n949 43.6538
R1483 B.n949 B.n64 43.6538
R1484 B.n943 B.n64 43.6538
R1485 B.n942 B.n941 43.6538
R1486 B.n941 B.n71 43.6538
R1487 B.n935 B.n71 43.6538
R1488 B.n935 B.n934 43.6538
R1489 B.n934 B.n933 43.6538
R1490 B.n933 B.n78 43.6538
R1491 B.n927 B.n78 43.6538
R1492 B.n927 B.n926 43.6538
R1493 B.n926 B.n925 43.6538
R1494 B.n925 B.n85 43.6538
R1495 B.n919 B.n918 43.6538
R1496 B.n918 B.n917 43.6538
R1497 B.n917 B.n92 43.6538
R1498 B.n911 B.n92 43.6538
R1499 B.n911 B.n910 43.6538
R1500 B.n910 B.n909 43.6538
R1501 B.n511 B.t11 42.3699
R1502 B.n919 B.t15 42.3699
R1503 B.n613 B.t2 38.5182
R1504 B.t7 B.n989 38.5182
R1505 B.n225 B.t8 37.2342
R1506 B.t3 B.n942 37.2342
R1507 B.n595 B.t6 34.6664
R1508 B.n975 B.t5 34.6664
R1509 B.n907 B.n906 34.1859
R1510 B.n722 B.n721 34.1859
R1511 B.n495 B.n255 34.1859
R1512 B.n491 B.n490 34.1859
R1513 B.n637 B.t1 24.395
R1514 B.t4 B.n1005 24.395
R1515 B.n209 B.t0 23.1111
R1516 B.t9 B.n958 23.1111
R1517 B.n571 B.t0 20.5432
R1518 B.n959 B.t9 20.5432
R1519 B.t1 B.n157 19.2593
R1520 B.n1006 B.t4 19.2593
R1521 B B.n1017 18.0485
R1522 B.n906 B.n905 10.6151
R1523 B.n905 B.n101 10.6151
R1524 B.n899 B.n101 10.6151
R1525 B.n899 B.n898 10.6151
R1526 B.n898 B.n897 10.6151
R1527 B.n897 B.n103 10.6151
R1528 B.n891 B.n103 10.6151
R1529 B.n891 B.n890 10.6151
R1530 B.n890 B.n889 10.6151
R1531 B.n889 B.n105 10.6151
R1532 B.n883 B.n105 10.6151
R1533 B.n883 B.n882 10.6151
R1534 B.n882 B.n881 10.6151
R1535 B.n881 B.n107 10.6151
R1536 B.n875 B.n107 10.6151
R1537 B.n875 B.n874 10.6151
R1538 B.n874 B.n873 10.6151
R1539 B.n873 B.n109 10.6151
R1540 B.n867 B.n109 10.6151
R1541 B.n867 B.n866 10.6151
R1542 B.n866 B.n865 10.6151
R1543 B.n865 B.n111 10.6151
R1544 B.n859 B.n111 10.6151
R1545 B.n859 B.n858 10.6151
R1546 B.n858 B.n857 10.6151
R1547 B.n857 B.n113 10.6151
R1548 B.n851 B.n113 10.6151
R1549 B.n851 B.n850 10.6151
R1550 B.n850 B.n849 10.6151
R1551 B.n849 B.n115 10.6151
R1552 B.n843 B.n115 10.6151
R1553 B.n843 B.n842 10.6151
R1554 B.n842 B.n841 10.6151
R1555 B.n841 B.n117 10.6151
R1556 B.n835 B.n117 10.6151
R1557 B.n835 B.n834 10.6151
R1558 B.n834 B.n833 10.6151
R1559 B.n833 B.n119 10.6151
R1560 B.n827 B.n119 10.6151
R1561 B.n827 B.n826 10.6151
R1562 B.n824 B.n123 10.6151
R1563 B.n818 B.n123 10.6151
R1564 B.n818 B.n817 10.6151
R1565 B.n817 B.n816 10.6151
R1566 B.n816 B.n125 10.6151
R1567 B.n810 B.n125 10.6151
R1568 B.n810 B.n809 10.6151
R1569 B.n809 B.n808 10.6151
R1570 B.n808 B.n127 10.6151
R1571 B.n802 B.n801 10.6151
R1572 B.n801 B.n800 10.6151
R1573 B.n800 B.n132 10.6151
R1574 B.n794 B.n132 10.6151
R1575 B.n794 B.n793 10.6151
R1576 B.n793 B.n792 10.6151
R1577 B.n792 B.n134 10.6151
R1578 B.n786 B.n134 10.6151
R1579 B.n786 B.n785 10.6151
R1580 B.n785 B.n784 10.6151
R1581 B.n784 B.n136 10.6151
R1582 B.n778 B.n136 10.6151
R1583 B.n778 B.n777 10.6151
R1584 B.n777 B.n776 10.6151
R1585 B.n776 B.n138 10.6151
R1586 B.n770 B.n138 10.6151
R1587 B.n770 B.n769 10.6151
R1588 B.n769 B.n768 10.6151
R1589 B.n768 B.n140 10.6151
R1590 B.n762 B.n140 10.6151
R1591 B.n762 B.n761 10.6151
R1592 B.n761 B.n760 10.6151
R1593 B.n760 B.n142 10.6151
R1594 B.n754 B.n142 10.6151
R1595 B.n754 B.n753 10.6151
R1596 B.n753 B.n752 10.6151
R1597 B.n752 B.n144 10.6151
R1598 B.n746 B.n144 10.6151
R1599 B.n746 B.n745 10.6151
R1600 B.n745 B.n744 10.6151
R1601 B.n744 B.n146 10.6151
R1602 B.n738 B.n146 10.6151
R1603 B.n738 B.n737 10.6151
R1604 B.n737 B.n736 10.6151
R1605 B.n736 B.n148 10.6151
R1606 B.n730 B.n148 10.6151
R1607 B.n730 B.n729 10.6151
R1608 B.n729 B.n728 10.6151
R1609 B.n728 B.n150 10.6151
R1610 B.n722 B.n150 10.6151
R1611 B.n496 B.n495 10.6151
R1612 B.n497 B.n496 10.6151
R1613 B.n497 B.n247 10.6151
R1614 B.n507 B.n247 10.6151
R1615 B.n508 B.n507 10.6151
R1616 B.n509 B.n508 10.6151
R1617 B.n509 B.n239 10.6151
R1618 B.n519 B.n239 10.6151
R1619 B.n520 B.n519 10.6151
R1620 B.n521 B.n520 10.6151
R1621 B.n521 B.n231 10.6151
R1622 B.n531 B.n231 10.6151
R1623 B.n532 B.n531 10.6151
R1624 B.n533 B.n532 10.6151
R1625 B.n533 B.n222 10.6151
R1626 B.n543 B.n222 10.6151
R1627 B.n544 B.n543 10.6151
R1628 B.n545 B.n544 10.6151
R1629 B.n545 B.n215 10.6151
R1630 B.n555 B.n215 10.6151
R1631 B.n556 B.n555 10.6151
R1632 B.n557 B.n556 10.6151
R1633 B.n557 B.n206 10.6151
R1634 B.n567 B.n206 10.6151
R1635 B.n568 B.n567 10.6151
R1636 B.n569 B.n568 10.6151
R1637 B.n569 B.n199 10.6151
R1638 B.n579 B.n199 10.6151
R1639 B.n580 B.n579 10.6151
R1640 B.n581 B.n580 10.6151
R1641 B.n581 B.n190 10.6151
R1642 B.n591 B.n190 10.6151
R1643 B.n592 B.n591 10.6151
R1644 B.n593 B.n592 10.6151
R1645 B.n593 B.n183 10.6151
R1646 B.n603 B.n183 10.6151
R1647 B.n604 B.n603 10.6151
R1648 B.n605 B.n604 10.6151
R1649 B.n605 B.n175 10.6151
R1650 B.n615 B.n175 10.6151
R1651 B.n616 B.n615 10.6151
R1652 B.n617 B.n616 10.6151
R1653 B.n617 B.n167 10.6151
R1654 B.n627 B.n167 10.6151
R1655 B.n628 B.n627 10.6151
R1656 B.n629 B.n628 10.6151
R1657 B.n629 B.n159 10.6151
R1658 B.n639 B.n159 10.6151
R1659 B.n640 B.n639 10.6151
R1660 B.n642 B.n640 10.6151
R1661 B.n642 B.n641 10.6151
R1662 B.n641 B.n151 10.6151
R1663 B.n653 B.n151 10.6151
R1664 B.n654 B.n653 10.6151
R1665 B.n655 B.n654 10.6151
R1666 B.n656 B.n655 10.6151
R1667 B.n658 B.n656 10.6151
R1668 B.n659 B.n658 10.6151
R1669 B.n660 B.n659 10.6151
R1670 B.n661 B.n660 10.6151
R1671 B.n663 B.n661 10.6151
R1672 B.n664 B.n663 10.6151
R1673 B.n665 B.n664 10.6151
R1674 B.n666 B.n665 10.6151
R1675 B.n668 B.n666 10.6151
R1676 B.n669 B.n668 10.6151
R1677 B.n670 B.n669 10.6151
R1678 B.n671 B.n670 10.6151
R1679 B.n673 B.n671 10.6151
R1680 B.n674 B.n673 10.6151
R1681 B.n675 B.n674 10.6151
R1682 B.n676 B.n675 10.6151
R1683 B.n678 B.n676 10.6151
R1684 B.n679 B.n678 10.6151
R1685 B.n680 B.n679 10.6151
R1686 B.n681 B.n680 10.6151
R1687 B.n683 B.n681 10.6151
R1688 B.n684 B.n683 10.6151
R1689 B.n685 B.n684 10.6151
R1690 B.n686 B.n685 10.6151
R1691 B.n688 B.n686 10.6151
R1692 B.n689 B.n688 10.6151
R1693 B.n690 B.n689 10.6151
R1694 B.n691 B.n690 10.6151
R1695 B.n693 B.n691 10.6151
R1696 B.n694 B.n693 10.6151
R1697 B.n695 B.n694 10.6151
R1698 B.n696 B.n695 10.6151
R1699 B.n698 B.n696 10.6151
R1700 B.n699 B.n698 10.6151
R1701 B.n700 B.n699 10.6151
R1702 B.n701 B.n700 10.6151
R1703 B.n703 B.n701 10.6151
R1704 B.n704 B.n703 10.6151
R1705 B.n705 B.n704 10.6151
R1706 B.n706 B.n705 10.6151
R1707 B.n708 B.n706 10.6151
R1708 B.n709 B.n708 10.6151
R1709 B.n710 B.n709 10.6151
R1710 B.n711 B.n710 10.6151
R1711 B.n713 B.n711 10.6151
R1712 B.n714 B.n713 10.6151
R1713 B.n715 B.n714 10.6151
R1714 B.n716 B.n715 10.6151
R1715 B.n718 B.n716 10.6151
R1716 B.n719 B.n718 10.6151
R1717 B.n720 B.n719 10.6151
R1718 B.n721 B.n720 10.6151
R1719 B.n490 B.n489 10.6151
R1720 B.n489 B.n259 10.6151
R1721 B.n484 B.n259 10.6151
R1722 B.n484 B.n483 10.6151
R1723 B.n483 B.n261 10.6151
R1724 B.n478 B.n261 10.6151
R1725 B.n478 B.n477 10.6151
R1726 B.n477 B.n476 10.6151
R1727 B.n476 B.n263 10.6151
R1728 B.n470 B.n263 10.6151
R1729 B.n470 B.n469 10.6151
R1730 B.n469 B.n468 10.6151
R1731 B.n468 B.n265 10.6151
R1732 B.n462 B.n265 10.6151
R1733 B.n462 B.n461 10.6151
R1734 B.n461 B.n460 10.6151
R1735 B.n460 B.n267 10.6151
R1736 B.n454 B.n267 10.6151
R1737 B.n454 B.n453 10.6151
R1738 B.n453 B.n452 10.6151
R1739 B.n452 B.n269 10.6151
R1740 B.n446 B.n269 10.6151
R1741 B.n446 B.n445 10.6151
R1742 B.n445 B.n444 10.6151
R1743 B.n444 B.n271 10.6151
R1744 B.n438 B.n271 10.6151
R1745 B.n438 B.n437 10.6151
R1746 B.n437 B.n436 10.6151
R1747 B.n436 B.n273 10.6151
R1748 B.n430 B.n273 10.6151
R1749 B.n430 B.n429 10.6151
R1750 B.n429 B.n428 10.6151
R1751 B.n428 B.n275 10.6151
R1752 B.n422 B.n275 10.6151
R1753 B.n422 B.n421 10.6151
R1754 B.n421 B.n420 10.6151
R1755 B.n420 B.n277 10.6151
R1756 B.n414 B.n277 10.6151
R1757 B.n414 B.n413 10.6151
R1758 B.n413 B.n412 10.6151
R1759 B.n408 B.n407 10.6151
R1760 B.n407 B.n283 10.6151
R1761 B.n402 B.n283 10.6151
R1762 B.n402 B.n401 10.6151
R1763 B.n401 B.n400 10.6151
R1764 B.n400 B.n285 10.6151
R1765 B.n394 B.n285 10.6151
R1766 B.n394 B.n393 10.6151
R1767 B.n393 B.n392 10.6151
R1768 B.n388 B.n387 10.6151
R1769 B.n387 B.n291 10.6151
R1770 B.n382 B.n291 10.6151
R1771 B.n382 B.n381 10.6151
R1772 B.n381 B.n380 10.6151
R1773 B.n380 B.n293 10.6151
R1774 B.n374 B.n293 10.6151
R1775 B.n374 B.n373 10.6151
R1776 B.n373 B.n372 10.6151
R1777 B.n372 B.n295 10.6151
R1778 B.n366 B.n295 10.6151
R1779 B.n366 B.n365 10.6151
R1780 B.n365 B.n364 10.6151
R1781 B.n364 B.n297 10.6151
R1782 B.n358 B.n297 10.6151
R1783 B.n358 B.n357 10.6151
R1784 B.n357 B.n356 10.6151
R1785 B.n356 B.n299 10.6151
R1786 B.n350 B.n299 10.6151
R1787 B.n350 B.n349 10.6151
R1788 B.n349 B.n348 10.6151
R1789 B.n348 B.n301 10.6151
R1790 B.n342 B.n301 10.6151
R1791 B.n342 B.n341 10.6151
R1792 B.n341 B.n340 10.6151
R1793 B.n340 B.n303 10.6151
R1794 B.n334 B.n303 10.6151
R1795 B.n334 B.n333 10.6151
R1796 B.n333 B.n332 10.6151
R1797 B.n332 B.n305 10.6151
R1798 B.n326 B.n305 10.6151
R1799 B.n326 B.n325 10.6151
R1800 B.n325 B.n324 10.6151
R1801 B.n324 B.n307 10.6151
R1802 B.n318 B.n307 10.6151
R1803 B.n318 B.n317 10.6151
R1804 B.n317 B.n316 10.6151
R1805 B.n316 B.n309 10.6151
R1806 B.n310 B.n309 10.6151
R1807 B.n310 B.n255 10.6151
R1808 B.n491 B.n251 10.6151
R1809 B.n501 B.n251 10.6151
R1810 B.n502 B.n501 10.6151
R1811 B.n503 B.n502 10.6151
R1812 B.n503 B.n243 10.6151
R1813 B.n513 B.n243 10.6151
R1814 B.n514 B.n513 10.6151
R1815 B.n515 B.n514 10.6151
R1816 B.n515 B.n235 10.6151
R1817 B.n525 B.n235 10.6151
R1818 B.n526 B.n525 10.6151
R1819 B.n527 B.n526 10.6151
R1820 B.n527 B.n227 10.6151
R1821 B.n537 B.n227 10.6151
R1822 B.n538 B.n537 10.6151
R1823 B.n539 B.n538 10.6151
R1824 B.n539 B.n219 10.6151
R1825 B.n549 B.n219 10.6151
R1826 B.n550 B.n549 10.6151
R1827 B.n551 B.n550 10.6151
R1828 B.n551 B.n211 10.6151
R1829 B.n561 B.n211 10.6151
R1830 B.n562 B.n561 10.6151
R1831 B.n563 B.n562 10.6151
R1832 B.n563 B.n203 10.6151
R1833 B.n573 B.n203 10.6151
R1834 B.n574 B.n573 10.6151
R1835 B.n575 B.n574 10.6151
R1836 B.n575 B.n195 10.6151
R1837 B.n585 B.n195 10.6151
R1838 B.n586 B.n585 10.6151
R1839 B.n587 B.n586 10.6151
R1840 B.n587 B.n187 10.6151
R1841 B.n597 B.n187 10.6151
R1842 B.n598 B.n597 10.6151
R1843 B.n599 B.n598 10.6151
R1844 B.n599 B.n179 10.6151
R1845 B.n609 B.n179 10.6151
R1846 B.n610 B.n609 10.6151
R1847 B.n611 B.n610 10.6151
R1848 B.n611 B.n171 10.6151
R1849 B.n621 B.n171 10.6151
R1850 B.n622 B.n621 10.6151
R1851 B.n623 B.n622 10.6151
R1852 B.n623 B.n163 10.6151
R1853 B.n633 B.n163 10.6151
R1854 B.n634 B.n633 10.6151
R1855 B.n635 B.n634 10.6151
R1856 B.n635 B.n155 10.6151
R1857 B.n646 B.n155 10.6151
R1858 B.n647 B.n646 10.6151
R1859 B.n648 B.n647 10.6151
R1860 B.n648 B.n0 10.6151
R1861 B.n1011 B.n1 10.6151
R1862 B.n1011 B.n1010 10.6151
R1863 B.n1010 B.n1009 10.6151
R1864 B.n1009 B.n10 10.6151
R1865 B.n1003 B.n10 10.6151
R1866 B.n1003 B.n1002 10.6151
R1867 B.n1002 B.n1001 10.6151
R1868 B.n1001 B.n17 10.6151
R1869 B.n995 B.n17 10.6151
R1870 B.n995 B.n994 10.6151
R1871 B.n994 B.n993 10.6151
R1872 B.n993 B.n24 10.6151
R1873 B.n987 B.n24 10.6151
R1874 B.n987 B.n986 10.6151
R1875 B.n986 B.n985 10.6151
R1876 B.n985 B.n31 10.6151
R1877 B.n979 B.n31 10.6151
R1878 B.n979 B.n978 10.6151
R1879 B.n978 B.n977 10.6151
R1880 B.n977 B.n38 10.6151
R1881 B.n971 B.n38 10.6151
R1882 B.n971 B.n970 10.6151
R1883 B.n970 B.n969 10.6151
R1884 B.n969 B.n45 10.6151
R1885 B.n963 B.n45 10.6151
R1886 B.n963 B.n962 10.6151
R1887 B.n962 B.n961 10.6151
R1888 B.n961 B.n52 10.6151
R1889 B.n955 B.n52 10.6151
R1890 B.n955 B.n954 10.6151
R1891 B.n954 B.n953 10.6151
R1892 B.n953 B.n59 10.6151
R1893 B.n947 B.n59 10.6151
R1894 B.n947 B.n946 10.6151
R1895 B.n946 B.n945 10.6151
R1896 B.n945 B.n66 10.6151
R1897 B.n939 B.n66 10.6151
R1898 B.n939 B.n938 10.6151
R1899 B.n938 B.n937 10.6151
R1900 B.n937 B.n73 10.6151
R1901 B.n931 B.n73 10.6151
R1902 B.n931 B.n930 10.6151
R1903 B.n930 B.n929 10.6151
R1904 B.n929 B.n80 10.6151
R1905 B.n923 B.n80 10.6151
R1906 B.n923 B.n922 10.6151
R1907 B.n922 B.n921 10.6151
R1908 B.n921 B.n87 10.6151
R1909 B.n915 B.n87 10.6151
R1910 B.n915 B.n914 10.6151
R1911 B.n914 B.n913 10.6151
R1912 B.n913 B.n94 10.6151
R1913 B.n907 B.n94 10.6151
R1914 B.n826 B.n825 9.36635
R1915 B.n802 B.n131 9.36635
R1916 B.n412 B.n281 9.36635
R1917 B.n388 B.n289 9.36635
R1918 B.n193 B.t6 8.98795
R1919 B.t5 B.n974 8.98795
R1920 B.n547 B.t8 6.42011
R1921 B.n943 B.t3 6.42011
R1922 B.t2 B.n173 5.13619
R1923 B.n990 B.t7 5.13619
R1924 B.n1017 B.n0 2.81026
R1925 B.n1017 B.n1 2.81026
R1926 B.t11 B.n241 1.28442
R1927 B.t15 B.n85 1.28442
R1928 B.n825 B.n824 1.24928
R1929 B.n131 B.n127 1.24928
R1930 B.n408 B.n281 1.24928
R1931 B.n392 B.n289 1.24928
R1932 VP.n22 VP.n21 161.3
R1933 VP.n23 VP.n18 161.3
R1934 VP.n25 VP.n24 161.3
R1935 VP.n26 VP.n17 161.3
R1936 VP.n28 VP.n27 161.3
R1937 VP.n29 VP.n16 161.3
R1938 VP.n31 VP.n30 161.3
R1939 VP.n32 VP.n15 161.3
R1940 VP.n34 VP.n33 161.3
R1941 VP.n35 VP.n14 161.3
R1942 VP.n37 VP.n36 161.3
R1943 VP.n39 VP.n13 161.3
R1944 VP.n41 VP.n40 161.3
R1945 VP.n42 VP.n12 161.3
R1946 VP.n44 VP.n43 161.3
R1947 VP.n45 VP.n11 161.3
R1948 VP.n82 VP.n0 161.3
R1949 VP.n81 VP.n80 161.3
R1950 VP.n79 VP.n1 161.3
R1951 VP.n78 VP.n77 161.3
R1952 VP.n76 VP.n2 161.3
R1953 VP.n74 VP.n73 161.3
R1954 VP.n72 VP.n3 161.3
R1955 VP.n71 VP.n70 161.3
R1956 VP.n69 VP.n4 161.3
R1957 VP.n68 VP.n67 161.3
R1958 VP.n66 VP.n5 161.3
R1959 VP.n65 VP.n64 161.3
R1960 VP.n63 VP.n6 161.3
R1961 VP.n62 VP.n61 161.3
R1962 VP.n60 VP.n7 161.3
R1963 VP.n59 VP.n58 161.3
R1964 VP.n56 VP.n8 161.3
R1965 VP.n55 VP.n54 161.3
R1966 VP.n53 VP.n9 161.3
R1967 VP.n52 VP.n51 161.3
R1968 VP.n50 VP.n10 161.3
R1969 VP.n19 VP.t1 156.679
R1970 VP.n5 VP.t3 125.362
R1971 VP.n49 VP.t2 125.362
R1972 VP.n57 VP.t9 125.362
R1973 VP.n75 VP.t7 125.362
R1974 VP.n83 VP.t5 125.362
R1975 VP.n16 VP.t8 125.362
R1976 VP.n46 VP.t4 125.362
R1977 VP.n38 VP.t0 125.362
R1978 VP.n20 VP.t6 125.362
R1979 VP.n49 VP.n48 100.088
R1980 VP.n84 VP.n83 100.088
R1981 VP.n47 VP.n46 100.088
R1982 VP.n20 VP.n19 66.8721
R1983 VP.n63 VP.n62 56.5617
R1984 VP.n70 VP.n69 56.5617
R1985 VP.n33 VP.n32 56.5617
R1986 VP.n26 VP.n25 56.5617
R1987 VP.n48 VP.n47 51.2231
R1988 VP.n55 VP.n9 48.8116
R1989 VP.n77 VP.n1 48.8116
R1990 VP.n40 VP.n12 48.8116
R1991 VP.n51 VP.n9 32.3425
R1992 VP.n81 VP.n1 32.3425
R1993 VP.n44 VP.n12 32.3425
R1994 VP.n51 VP.n50 24.5923
R1995 VP.n56 VP.n55 24.5923
R1996 VP.n58 VP.n7 24.5923
R1997 VP.n62 VP.n7 24.5923
R1998 VP.n64 VP.n63 24.5923
R1999 VP.n64 VP.n5 24.5923
R2000 VP.n68 VP.n5 24.5923
R2001 VP.n69 VP.n68 24.5923
R2002 VP.n70 VP.n3 24.5923
R2003 VP.n74 VP.n3 24.5923
R2004 VP.n77 VP.n76 24.5923
R2005 VP.n82 VP.n81 24.5923
R2006 VP.n45 VP.n44 24.5923
R2007 VP.n33 VP.n14 24.5923
R2008 VP.n37 VP.n14 24.5923
R2009 VP.n40 VP.n39 24.5923
R2010 VP.n27 VP.n26 24.5923
R2011 VP.n27 VP.n16 24.5923
R2012 VP.n31 VP.n16 24.5923
R2013 VP.n32 VP.n31 24.5923
R2014 VP.n21 VP.n18 24.5923
R2015 VP.n25 VP.n18 24.5923
R2016 VP.n57 VP.n56 19.1821
R2017 VP.n76 VP.n75 19.1821
R2018 VP.n39 VP.n38 19.1821
R2019 VP.n50 VP.n49 10.8209
R2020 VP.n83 VP.n82 10.8209
R2021 VP.n46 VP.n45 10.8209
R2022 VP.n22 VP.n19 9.89957
R2023 VP.n58 VP.n57 5.4107
R2024 VP.n75 VP.n74 5.4107
R2025 VP.n38 VP.n37 5.4107
R2026 VP.n21 VP.n20 5.4107
R2027 VP.n47 VP.n11 0.278335
R2028 VP.n48 VP.n10 0.278335
R2029 VP.n84 VP.n0 0.278335
R2030 VP.n23 VP.n22 0.189894
R2031 VP.n24 VP.n23 0.189894
R2032 VP.n24 VP.n17 0.189894
R2033 VP.n28 VP.n17 0.189894
R2034 VP.n29 VP.n28 0.189894
R2035 VP.n30 VP.n29 0.189894
R2036 VP.n30 VP.n15 0.189894
R2037 VP.n34 VP.n15 0.189894
R2038 VP.n35 VP.n34 0.189894
R2039 VP.n36 VP.n35 0.189894
R2040 VP.n36 VP.n13 0.189894
R2041 VP.n41 VP.n13 0.189894
R2042 VP.n42 VP.n41 0.189894
R2043 VP.n43 VP.n42 0.189894
R2044 VP.n43 VP.n11 0.189894
R2045 VP.n52 VP.n10 0.189894
R2046 VP.n53 VP.n52 0.189894
R2047 VP.n54 VP.n53 0.189894
R2048 VP.n54 VP.n8 0.189894
R2049 VP.n59 VP.n8 0.189894
R2050 VP.n60 VP.n59 0.189894
R2051 VP.n61 VP.n60 0.189894
R2052 VP.n61 VP.n6 0.189894
R2053 VP.n65 VP.n6 0.189894
R2054 VP.n66 VP.n65 0.189894
R2055 VP.n67 VP.n66 0.189894
R2056 VP.n67 VP.n4 0.189894
R2057 VP.n71 VP.n4 0.189894
R2058 VP.n72 VP.n71 0.189894
R2059 VP.n73 VP.n72 0.189894
R2060 VP.n73 VP.n2 0.189894
R2061 VP.n78 VP.n2 0.189894
R2062 VP.n79 VP.n78 0.189894
R2063 VP.n80 VP.n79 0.189894
R2064 VP.n80 VP.n0 0.189894
R2065 VP VP.n84 0.153485
R2066 VDD1.n1 VDD1.t8 67.8389
R2067 VDD1.n3 VDD1.t7 67.8387
R2068 VDD1.n5 VDD1.n4 65.5513
R2069 VDD1.n1 VDD1.n0 63.9194
R2070 VDD1.n7 VDD1.n6 63.9192
R2071 VDD1.n3 VDD1.n2 63.9192
R2072 VDD1.n7 VDD1.n5 46.3349
R2073 VDD1.n6 VDD1.t9 1.66998
R2074 VDD1.n6 VDD1.t5 1.66998
R2075 VDD1.n0 VDD1.t3 1.66998
R2076 VDD1.n0 VDD1.t1 1.66998
R2077 VDD1.n4 VDD1.t2 1.66998
R2078 VDD1.n4 VDD1.t4 1.66998
R2079 VDD1.n2 VDD1.t0 1.66998
R2080 VDD1.n2 VDD1.t6 1.66998
R2081 VDD1 VDD1.n7 1.62981
R2082 VDD1 VDD1.n1 0.62119
R2083 VDD1.n5 VDD1.n3 0.507654
C0 VDD1 VP 10.6447f
C1 VDD2 VDD1 1.96619f
C2 VN VP 7.89784f
C3 VDD2 VN 10.258401f
C4 VDD2 VP 0.543094f
C5 VTAIL VDD1 10.3039f
C6 VTAIL VN 10.7725f
C7 VTAIL VP 10.786799f
C8 VDD2 VTAIL 10.3524f
C9 VN VDD1 0.152964f
C10 VDD2 B 6.775081f
C11 VDD1 B 6.7717f
C12 VTAIL B 7.903029f
C13 VN B 16.62003f
C14 VP B 15.11545f
C15 VDD1.t8 B 2.392f
C16 VDD1.t3 B 0.209212f
C17 VDD1.t1 B 0.209212f
C18 VDD1.n0 B 1.86447f
C19 VDD1.n1 B 0.786388f
C20 VDD1.t7 B 2.392f
C21 VDD1.t0 B 0.209212f
C22 VDD1.t6 B 0.209212f
C23 VDD1.n2 B 1.86446f
C24 VDD1.n3 B 0.779249f
C25 VDD1.t2 B 0.209212f
C26 VDD1.t4 B 0.209212f
C27 VDD1.n4 B 1.8762f
C28 VDD1.n5 B 2.54062f
C29 VDD1.t9 B 0.209212f
C30 VDD1.t5 B 0.209212f
C31 VDD1.n6 B 1.86446f
C32 VDD1.n7 B 2.70462f
C33 VP.n0 B 0.031199f
C34 VP.t5 B 1.74301f
C35 VP.n1 B 0.021387f
C36 VP.n2 B 0.023666f
C37 VP.t7 B 1.74301f
C38 VP.n3 B 0.043886f
C39 VP.n4 B 0.023666f
C40 VP.t3 B 1.74301f
C41 VP.n5 B 0.64169f
C42 VP.n6 B 0.023666f
C43 VP.n7 B 0.043886f
C44 VP.n8 B 0.023666f
C45 VP.t9 B 1.74301f
C46 VP.n9 B 0.021387f
C47 VP.n10 B 0.031199f
C48 VP.t2 B 1.74301f
C49 VP.n11 B 0.031199f
C50 VP.t4 B 1.74301f
C51 VP.n12 B 0.021387f
C52 VP.n13 B 0.023666f
C53 VP.t0 B 1.74301f
C54 VP.n14 B 0.043886f
C55 VP.n15 B 0.023666f
C56 VP.t8 B 1.74301f
C57 VP.n16 B 0.64169f
C58 VP.n17 B 0.023666f
C59 VP.n18 B 0.043886f
C60 VP.t1 B 1.89218f
C61 VP.n19 B 0.674166f
C62 VP.t6 B 1.74301f
C63 VP.n20 B 0.676384f
C64 VP.n21 B 0.026987f
C65 VP.n22 B 0.203087f
C66 VP.n23 B 0.023666f
C67 VP.n24 B 0.023666f
C68 VP.n25 B 0.030801f
C69 VP.n26 B 0.038003f
C70 VP.n27 B 0.043886f
C71 VP.n28 B 0.023666f
C72 VP.n29 B 0.023666f
C73 VP.n30 B 0.023666f
C74 VP.n31 B 0.043886f
C75 VP.n32 B 0.038003f
C76 VP.n33 B 0.030801f
C77 VP.n34 B 0.023666f
C78 VP.n35 B 0.023666f
C79 VP.n36 B 0.023666f
C80 VP.n37 B 0.026987f
C81 VP.n38 B 0.61947f
C82 VP.n39 B 0.03912f
C83 VP.n40 B 0.043886f
C84 VP.n41 B 0.023666f
C85 VP.n42 B 0.023666f
C86 VP.n43 B 0.023666f
C87 VP.n44 B 0.047416f
C88 VP.n45 B 0.031753f
C89 VP.n46 B 0.68907f
C90 VP.n47 B 1.36038f
C91 VP.n48 B 1.37704f
C92 VP.n49 B 0.68907f
C93 VP.n50 B 0.031753f
C94 VP.n51 B 0.047416f
C95 VP.n52 B 0.023666f
C96 VP.n53 B 0.023666f
C97 VP.n54 B 0.023666f
C98 VP.n55 B 0.043886f
C99 VP.n56 B 0.03912f
C100 VP.n57 B 0.61947f
C101 VP.n58 B 0.026987f
C102 VP.n59 B 0.023666f
C103 VP.n60 B 0.023666f
C104 VP.n61 B 0.023666f
C105 VP.n62 B 0.030801f
C106 VP.n63 B 0.038003f
C107 VP.n64 B 0.043886f
C108 VP.n65 B 0.023666f
C109 VP.n66 B 0.023666f
C110 VP.n67 B 0.023666f
C111 VP.n68 B 0.043886f
C112 VP.n69 B 0.038003f
C113 VP.n70 B 0.030801f
C114 VP.n71 B 0.023666f
C115 VP.n72 B 0.023666f
C116 VP.n73 B 0.023666f
C117 VP.n74 B 0.026987f
C118 VP.n75 B 0.61947f
C119 VP.n76 B 0.03912f
C120 VP.n77 B 0.043886f
C121 VP.n78 B 0.023666f
C122 VP.n79 B 0.023666f
C123 VP.n80 B 0.023666f
C124 VP.n81 B 0.047416f
C125 VP.n82 B 0.031753f
C126 VP.n83 B 0.68907f
C127 VP.n84 B 0.035729f
C128 VTAIL.t13 B 0.232829f
C129 VTAIL.t15 B 0.232829f
C130 VTAIL.n0 B 2.00469f
C131 VTAIL.n1 B 0.50756f
C132 VTAIL.t1 B 2.55752f
C133 VTAIL.n2 B 0.630085f
C134 VTAIL.t6 B 0.232829f
C135 VTAIL.t2 B 0.232829f
C136 VTAIL.n3 B 2.00469f
C137 VTAIL.n4 B 0.600375f
C138 VTAIL.t8 B 0.232829f
C139 VTAIL.t0 B 0.232829f
C140 VTAIL.n5 B 2.00469f
C141 VTAIL.n6 B 1.93637f
C142 VTAIL.t17 B 0.232829f
C143 VTAIL.t18 B 0.232829f
C144 VTAIL.n7 B 2.0047f
C145 VTAIL.n8 B 1.93637f
C146 VTAIL.t12 B 0.232829f
C147 VTAIL.t9 B 0.232829f
C148 VTAIL.n9 B 2.0047f
C149 VTAIL.n10 B 0.600369f
C150 VTAIL.t11 B 2.55753f
C151 VTAIL.n11 B 0.630079f
C152 VTAIL.t4 B 0.232829f
C153 VTAIL.t7 B 0.232829f
C154 VTAIL.n12 B 2.0047f
C155 VTAIL.n13 B 0.547923f
C156 VTAIL.t5 B 0.232829f
C157 VTAIL.t19 B 0.232829f
C158 VTAIL.n14 B 2.0047f
C159 VTAIL.n15 B 0.600369f
C160 VTAIL.t3 B 2.55752f
C161 VTAIL.n16 B 1.83842f
C162 VTAIL.t16 B 2.55752f
C163 VTAIL.n17 B 1.83842f
C164 VTAIL.t14 B 0.232829f
C165 VTAIL.t10 B 0.232829f
C166 VTAIL.n18 B 2.00469f
C167 VTAIL.n19 B 0.460635f
C168 VDD2.t5 B 2.37849f
C169 VDD2.t3 B 0.20803f
C170 VDD2.t2 B 0.20803f
C171 VDD2.n0 B 1.85393f
C172 VDD2.n1 B 0.774849f
C173 VDD2.t6 B 0.20803f
C174 VDD2.t0 B 0.20803f
C175 VDD2.n2 B 1.86561f
C176 VDD2.n3 B 2.42288f
C177 VDD2.t1 B 2.36496f
C178 VDD2.n4 B 2.65056f
C179 VDD2.t8 B 0.20803f
C180 VDD2.t4 B 0.20803f
C181 VDD2.n5 B 1.85394f
C182 VDD2.n6 B 0.387301f
C183 VDD2.t9 B 0.20803f
C184 VDD2.t7 B 0.20803f
C185 VDD2.n7 B 1.86557f
C186 VN.n0 B 0.030845f
C187 VN.t2 B 1.72321f
C188 VN.n1 B 0.021144f
C189 VN.n2 B 0.023397f
C190 VN.t8 B 1.72321f
C191 VN.n3 B 0.043387f
C192 VN.n4 B 0.023397f
C193 VN.t4 B 1.72321f
C194 VN.n5 B 0.6344f
C195 VN.n6 B 0.023397f
C196 VN.n7 B 0.043387f
C197 VN.t5 B 1.87068f
C198 VN.n8 B 0.666506f
C199 VN.t3 B 1.72321f
C200 VN.n9 B 0.6687f
C201 VN.n10 B 0.02668f
C202 VN.n11 B 0.20078f
C203 VN.n12 B 0.023397f
C204 VN.n13 B 0.023397f
C205 VN.n14 B 0.030451f
C206 VN.n15 B 0.037571f
C207 VN.n16 B 0.043387f
C208 VN.n17 B 0.023397f
C209 VN.n18 B 0.023397f
C210 VN.n19 B 0.023397f
C211 VN.n20 B 0.043387f
C212 VN.n21 B 0.037571f
C213 VN.n22 B 0.030451f
C214 VN.n23 B 0.023397f
C215 VN.n24 B 0.023397f
C216 VN.n25 B 0.023397f
C217 VN.n26 B 0.02668f
C218 VN.n27 B 0.612432f
C219 VN.n28 B 0.038675f
C220 VN.n29 B 0.043387f
C221 VN.n30 B 0.023397f
C222 VN.n31 B 0.023397f
C223 VN.n32 B 0.023397f
C224 VN.n33 B 0.046878f
C225 VN.n34 B 0.031393f
C226 VN.n35 B 0.681242f
C227 VN.n36 B 0.035323f
C228 VN.n37 B 0.030845f
C229 VN.t1 B 1.72321f
C230 VN.n38 B 0.021144f
C231 VN.n39 B 0.023397f
C232 VN.t0 B 1.72321f
C233 VN.n40 B 0.043387f
C234 VN.n41 B 0.023397f
C235 VN.t6 B 1.72321f
C236 VN.n42 B 0.6344f
C237 VN.n43 B 0.023397f
C238 VN.n44 B 0.043387f
C239 VN.t7 B 1.87068f
C240 VN.n45 B 0.666506f
C241 VN.t9 B 1.72321f
C242 VN.n46 B 0.6687f
C243 VN.n47 B 0.02668f
C244 VN.n48 B 0.20078f
C245 VN.n49 B 0.023397f
C246 VN.n50 B 0.023397f
C247 VN.n51 B 0.030451f
C248 VN.n52 B 0.037571f
C249 VN.n53 B 0.043387f
C250 VN.n54 B 0.023397f
C251 VN.n55 B 0.023397f
C252 VN.n56 B 0.023397f
C253 VN.n57 B 0.043387f
C254 VN.n58 B 0.037571f
C255 VN.n59 B 0.030451f
C256 VN.n60 B 0.023397f
C257 VN.n61 B 0.023397f
C258 VN.n62 B 0.023397f
C259 VN.n63 B 0.02668f
C260 VN.n64 B 0.612432f
C261 VN.n65 B 0.038675f
C262 VN.n66 B 0.043387f
C263 VN.n67 B 0.023397f
C264 VN.n68 B 0.023397f
C265 VN.n69 B 0.023397f
C266 VN.n70 B 0.046878f
C267 VN.n71 B 0.031393f
C268 VN.n72 B 0.681242f
C269 VN.n73 B 1.35745f
.ends

