* NGSPICE file created from diff_pair_sample_1162.ext - technology: sky130A

.subckt diff_pair_sample_1162 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t16 B.t4 sky130_fd_pr__nfet_01v8 ad=3.11025 pd=19.18 as=3.11025 ps=19.18 w=18.85 l=2.37
X1 VTAIL.t19 VN.t1 VDD2.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=3.11025 pd=19.18 as=3.11025 ps=19.18 w=18.85 l=2.37
X2 VTAIL.t8 VP.t0 VDD1.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=3.11025 pd=19.18 as=3.11025 ps=19.18 w=18.85 l=2.37
X3 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=7.3515 pd=38.48 as=0 ps=0 w=18.85 l=2.37
X4 VDD1.t8 VP.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=7.3515 pd=38.48 as=3.11025 ps=19.18 w=18.85 l=2.37
X5 VDD1.t7 VP.t2 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=3.11025 pd=19.18 as=7.3515 ps=38.48 w=18.85 l=2.37
X6 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=7.3515 pd=38.48 as=0 ps=0 w=18.85 l=2.37
X7 VDD1.t6 VP.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.11025 pd=19.18 as=3.11025 ps=19.18 w=18.85 l=2.37
X8 VTAIL.t15 VN.t2 VDD2.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=3.11025 pd=19.18 as=3.11025 ps=19.18 w=18.85 l=2.37
X9 VDD2.t6 VN.t3 VTAIL.t11 B.t9 sky130_fd_pr__nfet_01v8 ad=3.11025 pd=19.18 as=7.3515 ps=38.48 w=18.85 l=2.37
X10 VTAIL.t3 VP.t4 VDD1.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=3.11025 pd=19.18 as=3.11025 ps=19.18 w=18.85 l=2.37
X11 VTAIL.t14 VN.t4 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=3.11025 pd=19.18 as=3.11025 ps=19.18 w=18.85 l=2.37
X12 VDD1.t4 VP.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.3515 pd=38.48 as=3.11025 ps=19.18 w=18.85 l=2.37
X13 VDD1.t3 VP.t6 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=3.11025 pd=19.18 as=7.3515 ps=38.48 w=18.85 l=2.37
X14 VDD2.t4 VN.t5 VTAIL.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=3.11025 pd=19.18 as=7.3515 ps=38.48 w=18.85 l=2.37
X15 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=7.3515 pd=38.48 as=0 ps=0 w=18.85 l=2.37
X16 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.3515 pd=38.48 as=0 ps=0 w=18.85 l=2.37
X17 VTAIL.t12 VN.t6 VDD2.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=3.11025 pd=19.18 as=3.11025 ps=19.18 w=18.85 l=2.37
X18 VDD1.t2 VP.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.11025 pd=19.18 as=3.11025 ps=19.18 w=18.85 l=2.37
X19 VTAIL.t6 VP.t8 VDD1.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=3.11025 pd=19.18 as=3.11025 ps=19.18 w=18.85 l=2.37
X20 VDD2.t2 VN.t7 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=7.3515 pd=38.48 as=3.11025 ps=19.18 w=18.85 l=2.37
X21 VTAIL.t2 VP.t9 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=3.11025 pd=19.18 as=3.11025 ps=19.18 w=18.85 l=2.37
X22 VDD2.t1 VN.t8 VTAIL.t17 B.t0 sky130_fd_pr__nfet_01v8 ad=3.11025 pd=19.18 as=3.11025 ps=19.18 w=18.85 l=2.37
X23 VDD2.t0 VN.t9 VTAIL.t13 B.t1 sky130_fd_pr__nfet_01v8 ad=7.3515 pd=38.48 as=3.11025 ps=19.18 w=18.85 l=2.37
R0 VN.n9 VN.t9 224.499
R1 VN.n47 VN.t5 224.499
R2 VN.n10 VN.t4 191.681
R3 VN.n18 VN.t0 191.681
R4 VN.n3 VN.t6 191.681
R5 VN.n36 VN.t3 191.681
R6 VN.n48 VN.t1 191.681
R7 VN.n56 VN.t8 191.681
R8 VN.n41 VN.t2 191.681
R9 VN.n74 VN.t7 191.681
R10 VN.n73 VN.n38 161.3
R11 VN.n72 VN.n71 161.3
R12 VN.n70 VN.n39 161.3
R13 VN.n69 VN.n68 161.3
R14 VN.n67 VN.n40 161.3
R15 VN.n66 VN.n65 161.3
R16 VN.n64 VN.n63 161.3
R17 VN.n62 VN.n42 161.3
R18 VN.n61 VN.n60 161.3
R19 VN.n59 VN.n43 161.3
R20 VN.n58 VN.n57 161.3
R21 VN.n55 VN.n44 161.3
R22 VN.n54 VN.n53 161.3
R23 VN.n52 VN.n45 161.3
R24 VN.n51 VN.n50 161.3
R25 VN.n49 VN.n46 161.3
R26 VN.n35 VN.n0 161.3
R27 VN.n34 VN.n33 161.3
R28 VN.n32 VN.n1 161.3
R29 VN.n31 VN.n30 161.3
R30 VN.n29 VN.n2 161.3
R31 VN.n28 VN.n27 161.3
R32 VN.n26 VN.n25 161.3
R33 VN.n24 VN.n4 161.3
R34 VN.n23 VN.n22 161.3
R35 VN.n21 VN.n5 161.3
R36 VN.n20 VN.n19 161.3
R37 VN.n17 VN.n6 161.3
R38 VN.n16 VN.n15 161.3
R39 VN.n14 VN.n7 161.3
R40 VN.n13 VN.n12 161.3
R41 VN.n11 VN.n8 161.3
R42 VN.n37 VN.n36 103.416
R43 VN.n75 VN.n74 103.416
R44 VN VN.n75 57.2557
R45 VN.n30 VN.n1 56.5193
R46 VN.n68 VN.n39 56.5193
R47 VN.n10 VN.n9 50.2654
R48 VN.n48 VN.n47 50.2654
R49 VN.n12 VN.n7 50.2061
R50 VN.n24 VN.n23 50.2061
R51 VN.n50 VN.n45 50.2061
R52 VN.n62 VN.n61 50.2061
R53 VN.n16 VN.n7 30.7807
R54 VN.n23 VN.n5 30.7807
R55 VN.n54 VN.n45 30.7807
R56 VN.n61 VN.n43 30.7807
R57 VN.n12 VN.n11 24.4675
R58 VN.n17 VN.n16 24.4675
R59 VN.n19 VN.n5 24.4675
R60 VN.n25 VN.n24 24.4675
R61 VN.n29 VN.n28 24.4675
R62 VN.n30 VN.n29 24.4675
R63 VN.n34 VN.n1 24.4675
R64 VN.n35 VN.n34 24.4675
R65 VN.n50 VN.n49 24.4675
R66 VN.n57 VN.n43 24.4675
R67 VN.n55 VN.n54 24.4675
R68 VN.n68 VN.n67 24.4675
R69 VN.n67 VN.n66 24.4675
R70 VN.n63 VN.n62 24.4675
R71 VN.n73 VN.n72 24.4675
R72 VN.n72 VN.n39 24.4675
R73 VN.n11 VN.n10 22.0208
R74 VN.n25 VN.n3 22.0208
R75 VN.n49 VN.n48 22.0208
R76 VN.n63 VN.n41 22.0208
R77 VN.n18 VN.n17 12.234
R78 VN.n19 VN.n18 12.234
R79 VN.n57 VN.n56 12.234
R80 VN.n56 VN.n55 12.234
R81 VN.n36 VN.n35 7.3406
R82 VN.n74 VN.n73 7.3406
R83 VN.n47 VN.n46 7.01727
R84 VN.n9 VN.n8 7.01727
R85 VN.n28 VN.n3 2.4472
R86 VN.n66 VN.n41 2.4472
R87 VN.n75 VN.n38 0.278367
R88 VN.n37 VN.n0 0.278367
R89 VN.n71 VN.n38 0.189894
R90 VN.n71 VN.n70 0.189894
R91 VN.n70 VN.n69 0.189894
R92 VN.n69 VN.n40 0.189894
R93 VN.n65 VN.n40 0.189894
R94 VN.n65 VN.n64 0.189894
R95 VN.n64 VN.n42 0.189894
R96 VN.n60 VN.n42 0.189894
R97 VN.n60 VN.n59 0.189894
R98 VN.n59 VN.n58 0.189894
R99 VN.n58 VN.n44 0.189894
R100 VN.n53 VN.n44 0.189894
R101 VN.n53 VN.n52 0.189894
R102 VN.n52 VN.n51 0.189894
R103 VN.n51 VN.n46 0.189894
R104 VN.n13 VN.n8 0.189894
R105 VN.n14 VN.n13 0.189894
R106 VN.n15 VN.n14 0.189894
R107 VN.n15 VN.n6 0.189894
R108 VN.n20 VN.n6 0.189894
R109 VN.n21 VN.n20 0.189894
R110 VN.n22 VN.n21 0.189894
R111 VN.n22 VN.n4 0.189894
R112 VN.n26 VN.n4 0.189894
R113 VN.n27 VN.n26 0.189894
R114 VN.n27 VN.n2 0.189894
R115 VN.n31 VN.n2 0.189894
R116 VN.n32 VN.n31 0.189894
R117 VN.n33 VN.n32 0.189894
R118 VN.n33 VN.n0 0.189894
R119 VN VN.n37 0.153454
R120 VTAIL.n432 VTAIL.n332 289.615
R121 VTAIL.n102 VTAIL.n2 289.615
R122 VTAIL.n326 VTAIL.n226 289.615
R123 VTAIL.n216 VTAIL.n116 289.615
R124 VTAIL.n367 VTAIL.n366 185
R125 VTAIL.n364 VTAIL.n363 185
R126 VTAIL.n373 VTAIL.n372 185
R127 VTAIL.n375 VTAIL.n374 185
R128 VTAIL.n360 VTAIL.n359 185
R129 VTAIL.n381 VTAIL.n380 185
R130 VTAIL.n383 VTAIL.n382 185
R131 VTAIL.n356 VTAIL.n355 185
R132 VTAIL.n389 VTAIL.n388 185
R133 VTAIL.n391 VTAIL.n390 185
R134 VTAIL.n352 VTAIL.n351 185
R135 VTAIL.n397 VTAIL.n396 185
R136 VTAIL.n399 VTAIL.n398 185
R137 VTAIL.n348 VTAIL.n347 185
R138 VTAIL.n405 VTAIL.n404 185
R139 VTAIL.n408 VTAIL.n407 185
R140 VTAIL.n406 VTAIL.n344 185
R141 VTAIL.n413 VTAIL.n343 185
R142 VTAIL.n415 VTAIL.n414 185
R143 VTAIL.n417 VTAIL.n416 185
R144 VTAIL.n340 VTAIL.n339 185
R145 VTAIL.n423 VTAIL.n422 185
R146 VTAIL.n425 VTAIL.n424 185
R147 VTAIL.n336 VTAIL.n335 185
R148 VTAIL.n431 VTAIL.n430 185
R149 VTAIL.n433 VTAIL.n432 185
R150 VTAIL.n37 VTAIL.n36 185
R151 VTAIL.n34 VTAIL.n33 185
R152 VTAIL.n43 VTAIL.n42 185
R153 VTAIL.n45 VTAIL.n44 185
R154 VTAIL.n30 VTAIL.n29 185
R155 VTAIL.n51 VTAIL.n50 185
R156 VTAIL.n53 VTAIL.n52 185
R157 VTAIL.n26 VTAIL.n25 185
R158 VTAIL.n59 VTAIL.n58 185
R159 VTAIL.n61 VTAIL.n60 185
R160 VTAIL.n22 VTAIL.n21 185
R161 VTAIL.n67 VTAIL.n66 185
R162 VTAIL.n69 VTAIL.n68 185
R163 VTAIL.n18 VTAIL.n17 185
R164 VTAIL.n75 VTAIL.n74 185
R165 VTAIL.n78 VTAIL.n77 185
R166 VTAIL.n76 VTAIL.n14 185
R167 VTAIL.n83 VTAIL.n13 185
R168 VTAIL.n85 VTAIL.n84 185
R169 VTAIL.n87 VTAIL.n86 185
R170 VTAIL.n10 VTAIL.n9 185
R171 VTAIL.n93 VTAIL.n92 185
R172 VTAIL.n95 VTAIL.n94 185
R173 VTAIL.n6 VTAIL.n5 185
R174 VTAIL.n101 VTAIL.n100 185
R175 VTAIL.n103 VTAIL.n102 185
R176 VTAIL.n327 VTAIL.n326 185
R177 VTAIL.n325 VTAIL.n324 185
R178 VTAIL.n230 VTAIL.n229 185
R179 VTAIL.n319 VTAIL.n318 185
R180 VTAIL.n317 VTAIL.n316 185
R181 VTAIL.n234 VTAIL.n233 185
R182 VTAIL.n311 VTAIL.n310 185
R183 VTAIL.n309 VTAIL.n308 185
R184 VTAIL.n307 VTAIL.n237 185
R185 VTAIL.n241 VTAIL.n238 185
R186 VTAIL.n302 VTAIL.n301 185
R187 VTAIL.n300 VTAIL.n299 185
R188 VTAIL.n243 VTAIL.n242 185
R189 VTAIL.n294 VTAIL.n293 185
R190 VTAIL.n292 VTAIL.n291 185
R191 VTAIL.n247 VTAIL.n246 185
R192 VTAIL.n286 VTAIL.n285 185
R193 VTAIL.n284 VTAIL.n283 185
R194 VTAIL.n251 VTAIL.n250 185
R195 VTAIL.n278 VTAIL.n277 185
R196 VTAIL.n276 VTAIL.n275 185
R197 VTAIL.n255 VTAIL.n254 185
R198 VTAIL.n270 VTAIL.n269 185
R199 VTAIL.n268 VTAIL.n267 185
R200 VTAIL.n259 VTAIL.n258 185
R201 VTAIL.n262 VTAIL.n261 185
R202 VTAIL.n217 VTAIL.n216 185
R203 VTAIL.n215 VTAIL.n214 185
R204 VTAIL.n120 VTAIL.n119 185
R205 VTAIL.n209 VTAIL.n208 185
R206 VTAIL.n207 VTAIL.n206 185
R207 VTAIL.n124 VTAIL.n123 185
R208 VTAIL.n201 VTAIL.n200 185
R209 VTAIL.n199 VTAIL.n198 185
R210 VTAIL.n197 VTAIL.n127 185
R211 VTAIL.n131 VTAIL.n128 185
R212 VTAIL.n192 VTAIL.n191 185
R213 VTAIL.n190 VTAIL.n189 185
R214 VTAIL.n133 VTAIL.n132 185
R215 VTAIL.n184 VTAIL.n183 185
R216 VTAIL.n182 VTAIL.n181 185
R217 VTAIL.n137 VTAIL.n136 185
R218 VTAIL.n176 VTAIL.n175 185
R219 VTAIL.n174 VTAIL.n173 185
R220 VTAIL.n141 VTAIL.n140 185
R221 VTAIL.n168 VTAIL.n167 185
R222 VTAIL.n166 VTAIL.n165 185
R223 VTAIL.n145 VTAIL.n144 185
R224 VTAIL.n160 VTAIL.n159 185
R225 VTAIL.n158 VTAIL.n157 185
R226 VTAIL.n149 VTAIL.n148 185
R227 VTAIL.n152 VTAIL.n151 185
R228 VTAIL.t9 VTAIL.n260 147.659
R229 VTAIL.t18 VTAIL.n150 147.659
R230 VTAIL.t11 VTAIL.n365 147.659
R231 VTAIL.t7 VTAIL.n35 147.659
R232 VTAIL.n366 VTAIL.n363 104.615
R233 VTAIL.n373 VTAIL.n363 104.615
R234 VTAIL.n374 VTAIL.n373 104.615
R235 VTAIL.n374 VTAIL.n359 104.615
R236 VTAIL.n381 VTAIL.n359 104.615
R237 VTAIL.n382 VTAIL.n381 104.615
R238 VTAIL.n382 VTAIL.n355 104.615
R239 VTAIL.n389 VTAIL.n355 104.615
R240 VTAIL.n390 VTAIL.n389 104.615
R241 VTAIL.n390 VTAIL.n351 104.615
R242 VTAIL.n397 VTAIL.n351 104.615
R243 VTAIL.n398 VTAIL.n397 104.615
R244 VTAIL.n398 VTAIL.n347 104.615
R245 VTAIL.n405 VTAIL.n347 104.615
R246 VTAIL.n407 VTAIL.n405 104.615
R247 VTAIL.n407 VTAIL.n406 104.615
R248 VTAIL.n406 VTAIL.n343 104.615
R249 VTAIL.n415 VTAIL.n343 104.615
R250 VTAIL.n416 VTAIL.n415 104.615
R251 VTAIL.n416 VTAIL.n339 104.615
R252 VTAIL.n423 VTAIL.n339 104.615
R253 VTAIL.n424 VTAIL.n423 104.615
R254 VTAIL.n424 VTAIL.n335 104.615
R255 VTAIL.n431 VTAIL.n335 104.615
R256 VTAIL.n432 VTAIL.n431 104.615
R257 VTAIL.n36 VTAIL.n33 104.615
R258 VTAIL.n43 VTAIL.n33 104.615
R259 VTAIL.n44 VTAIL.n43 104.615
R260 VTAIL.n44 VTAIL.n29 104.615
R261 VTAIL.n51 VTAIL.n29 104.615
R262 VTAIL.n52 VTAIL.n51 104.615
R263 VTAIL.n52 VTAIL.n25 104.615
R264 VTAIL.n59 VTAIL.n25 104.615
R265 VTAIL.n60 VTAIL.n59 104.615
R266 VTAIL.n60 VTAIL.n21 104.615
R267 VTAIL.n67 VTAIL.n21 104.615
R268 VTAIL.n68 VTAIL.n67 104.615
R269 VTAIL.n68 VTAIL.n17 104.615
R270 VTAIL.n75 VTAIL.n17 104.615
R271 VTAIL.n77 VTAIL.n75 104.615
R272 VTAIL.n77 VTAIL.n76 104.615
R273 VTAIL.n76 VTAIL.n13 104.615
R274 VTAIL.n85 VTAIL.n13 104.615
R275 VTAIL.n86 VTAIL.n85 104.615
R276 VTAIL.n86 VTAIL.n9 104.615
R277 VTAIL.n93 VTAIL.n9 104.615
R278 VTAIL.n94 VTAIL.n93 104.615
R279 VTAIL.n94 VTAIL.n5 104.615
R280 VTAIL.n101 VTAIL.n5 104.615
R281 VTAIL.n102 VTAIL.n101 104.615
R282 VTAIL.n326 VTAIL.n325 104.615
R283 VTAIL.n325 VTAIL.n229 104.615
R284 VTAIL.n318 VTAIL.n229 104.615
R285 VTAIL.n318 VTAIL.n317 104.615
R286 VTAIL.n317 VTAIL.n233 104.615
R287 VTAIL.n310 VTAIL.n233 104.615
R288 VTAIL.n310 VTAIL.n309 104.615
R289 VTAIL.n309 VTAIL.n237 104.615
R290 VTAIL.n241 VTAIL.n237 104.615
R291 VTAIL.n301 VTAIL.n241 104.615
R292 VTAIL.n301 VTAIL.n300 104.615
R293 VTAIL.n300 VTAIL.n242 104.615
R294 VTAIL.n293 VTAIL.n242 104.615
R295 VTAIL.n293 VTAIL.n292 104.615
R296 VTAIL.n292 VTAIL.n246 104.615
R297 VTAIL.n285 VTAIL.n246 104.615
R298 VTAIL.n285 VTAIL.n284 104.615
R299 VTAIL.n284 VTAIL.n250 104.615
R300 VTAIL.n277 VTAIL.n250 104.615
R301 VTAIL.n277 VTAIL.n276 104.615
R302 VTAIL.n276 VTAIL.n254 104.615
R303 VTAIL.n269 VTAIL.n254 104.615
R304 VTAIL.n269 VTAIL.n268 104.615
R305 VTAIL.n268 VTAIL.n258 104.615
R306 VTAIL.n261 VTAIL.n258 104.615
R307 VTAIL.n216 VTAIL.n215 104.615
R308 VTAIL.n215 VTAIL.n119 104.615
R309 VTAIL.n208 VTAIL.n119 104.615
R310 VTAIL.n208 VTAIL.n207 104.615
R311 VTAIL.n207 VTAIL.n123 104.615
R312 VTAIL.n200 VTAIL.n123 104.615
R313 VTAIL.n200 VTAIL.n199 104.615
R314 VTAIL.n199 VTAIL.n127 104.615
R315 VTAIL.n131 VTAIL.n127 104.615
R316 VTAIL.n191 VTAIL.n131 104.615
R317 VTAIL.n191 VTAIL.n190 104.615
R318 VTAIL.n190 VTAIL.n132 104.615
R319 VTAIL.n183 VTAIL.n132 104.615
R320 VTAIL.n183 VTAIL.n182 104.615
R321 VTAIL.n182 VTAIL.n136 104.615
R322 VTAIL.n175 VTAIL.n136 104.615
R323 VTAIL.n175 VTAIL.n174 104.615
R324 VTAIL.n174 VTAIL.n140 104.615
R325 VTAIL.n167 VTAIL.n140 104.615
R326 VTAIL.n167 VTAIL.n166 104.615
R327 VTAIL.n166 VTAIL.n144 104.615
R328 VTAIL.n159 VTAIL.n144 104.615
R329 VTAIL.n159 VTAIL.n158 104.615
R330 VTAIL.n158 VTAIL.n148 104.615
R331 VTAIL.n151 VTAIL.n148 104.615
R332 VTAIL.n366 VTAIL.t11 52.3082
R333 VTAIL.n36 VTAIL.t7 52.3082
R334 VTAIL.n261 VTAIL.t9 52.3082
R335 VTAIL.n151 VTAIL.t18 52.3082
R336 VTAIL.n439 VTAIL.n438 41.8099
R337 VTAIL.n1 VTAIL.n0 41.8099
R338 VTAIL.n109 VTAIL.n108 41.8099
R339 VTAIL.n111 VTAIL.n110 41.8099
R340 VTAIL.n225 VTAIL.n224 41.8099
R341 VTAIL.n223 VTAIL.n222 41.8099
R342 VTAIL.n115 VTAIL.n114 41.8099
R343 VTAIL.n113 VTAIL.n112 41.8099
R344 VTAIL.n113 VTAIL.n111 33.272
R345 VTAIL.n437 VTAIL.n331 30.9445
R346 VTAIL.n437 VTAIL.n436 30.052
R347 VTAIL.n107 VTAIL.n106 30.052
R348 VTAIL.n331 VTAIL.n330 30.052
R349 VTAIL.n221 VTAIL.n220 30.052
R350 VTAIL.n367 VTAIL.n365 15.6677
R351 VTAIL.n37 VTAIL.n35 15.6677
R352 VTAIL.n262 VTAIL.n260 15.6677
R353 VTAIL.n152 VTAIL.n150 15.6677
R354 VTAIL.n414 VTAIL.n413 13.1884
R355 VTAIL.n84 VTAIL.n83 13.1884
R356 VTAIL.n308 VTAIL.n307 13.1884
R357 VTAIL.n198 VTAIL.n197 13.1884
R358 VTAIL.n368 VTAIL.n364 12.8005
R359 VTAIL.n412 VTAIL.n344 12.8005
R360 VTAIL.n417 VTAIL.n342 12.8005
R361 VTAIL.n38 VTAIL.n34 12.8005
R362 VTAIL.n82 VTAIL.n14 12.8005
R363 VTAIL.n87 VTAIL.n12 12.8005
R364 VTAIL.n311 VTAIL.n236 12.8005
R365 VTAIL.n306 VTAIL.n238 12.8005
R366 VTAIL.n263 VTAIL.n259 12.8005
R367 VTAIL.n201 VTAIL.n126 12.8005
R368 VTAIL.n196 VTAIL.n128 12.8005
R369 VTAIL.n153 VTAIL.n149 12.8005
R370 VTAIL.n372 VTAIL.n371 12.0247
R371 VTAIL.n409 VTAIL.n408 12.0247
R372 VTAIL.n418 VTAIL.n340 12.0247
R373 VTAIL.n42 VTAIL.n41 12.0247
R374 VTAIL.n79 VTAIL.n78 12.0247
R375 VTAIL.n88 VTAIL.n10 12.0247
R376 VTAIL.n312 VTAIL.n234 12.0247
R377 VTAIL.n303 VTAIL.n302 12.0247
R378 VTAIL.n267 VTAIL.n266 12.0247
R379 VTAIL.n202 VTAIL.n124 12.0247
R380 VTAIL.n193 VTAIL.n192 12.0247
R381 VTAIL.n157 VTAIL.n156 12.0247
R382 VTAIL.n375 VTAIL.n362 11.249
R383 VTAIL.n404 VTAIL.n346 11.249
R384 VTAIL.n422 VTAIL.n421 11.249
R385 VTAIL.n45 VTAIL.n32 11.249
R386 VTAIL.n74 VTAIL.n16 11.249
R387 VTAIL.n92 VTAIL.n91 11.249
R388 VTAIL.n316 VTAIL.n315 11.249
R389 VTAIL.n299 VTAIL.n240 11.249
R390 VTAIL.n270 VTAIL.n257 11.249
R391 VTAIL.n206 VTAIL.n205 11.249
R392 VTAIL.n189 VTAIL.n130 11.249
R393 VTAIL.n160 VTAIL.n147 11.249
R394 VTAIL.n376 VTAIL.n360 10.4732
R395 VTAIL.n403 VTAIL.n348 10.4732
R396 VTAIL.n425 VTAIL.n338 10.4732
R397 VTAIL.n46 VTAIL.n30 10.4732
R398 VTAIL.n73 VTAIL.n18 10.4732
R399 VTAIL.n95 VTAIL.n8 10.4732
R400 VTAIL.n319 VTAIL.n232 10.4732
R401 VTAIL.n298 VTAIL.n243 10.4732
R402 VTAIL.n271 VTAIL.n255 10.4732
R403 VTAIL.n209 VTAIL.n122 10.4732
R404 VTAIL.n188 VTAIL.n133 10.4732
R405 VTAIL.n161 VTAIL.n145 10.4732
R406 VTAIL.n380 VTAIL.n379 9.69747
R407 VTAIL.n400 VTAIL.n399 9.69747
R408 VTAIL.n426 VTAIL.n336 9.69747
R409 VTAIL.n50 VTAIL.n49 9.69747
R410 VTAIL.n70 VTAIL.n69 9.69747
R411 VTAIL.n96 VTAIL.n6 9.69747
R412 VTAIL.n320 VTAIL.n230 9.69747
R413 VTAIL.n295 VTAIL.n294 9.69747
R414 VTAIL.n275 VTAIL.n274 9.69747
R415 VTAIL.n210 VTAIL.n120 9.69747
R416 VTAIL.n185 VTAIL.n184 9.69747
R417 VTAIL.n165 VTAIL.n164 9.69747
R418 VTAIL.n436 VTAIL.n435 9.45567
R419 VTAIL.n106 VTAIL.n105 9.45567
R420 VTAIL.n330 VTAIL.n329 9.45567
R421 VTAIL.n220 VTAIL.n219 9.45567
R422 VTAIL.n334 VTAIL.n333 9.3005
R423 VTAIL.n429 VTAIL.n428 9.3005
R424 VTAIL.n427 VTAIL.n426 9.3005
R425 VTAIL.n338 VTAIL.n337 9.3005
R426 VTAIL.n421 VTAIL.n420 9.3005
R427 VTAIL.n419 VTAIL.n418 9.3005
R428 VTAIL.n342 VTAIL.n341 9.3005
R429 VTAIL.n387 VTAIL.n386 9.3005
R430 VTAIL.n385 VTAIL.n384 9.3005
R431 VTAIL.n358 VTAIL.n357 9.3005
R432 VTAIL.n379 VTAIL.n378 9.3005
R433 VTAIL.n377 VTAIL.n376 9.3005
R434 VTAIL.n362 VTAIL.n361 9.3005
R435 VTAIL.n371 VTAIL.n370 9.3005
R436 VTAIL.n369 VTAIL.n368 9.3005
R437 VTAIL.n354 VTAIL.n353 9.3005
R438 VTAIL.n393 VTAIL.n392 9.3005
R439 VTAIL.n395 VTAIL.n394 9.3005
R440 VTAIL.n350 VTAIL.n349 9.3005
R441 VTAIL.n401 VTAIL.n400 9.3005
R442 VTAIL.n403 VTAIL.n402 9.3005
R443 VTAIL.n346 VTAIL.n345 9.3005
R444 VTAIL.n410 VTAIL.n409 9.3005
R445 VTAIL.n412 VTAIL.n411 9.3005
R446 VTAIL.n435 VTAIL.n434 9.3005
R447 VTAIL.n4 VTAIL.n3 9.3005
R448 VTAIL.n99 VTAIL.n98 9.3005
R449 VTAIL.n97 VTAIL.n96 9.3005
R450 VTAIL.n8 VTAIL.n7 9.3005
R451 VTAIL.n91 VTAIL.n90 9.3005
R452 VTAIL.n89 VTAIL.n88 9.3005
R453 VTAIL.n12 VTAIL.n11 9.3005
R454 VTAIL.n57 VTAIL.n56 9.3005
R455 VTAIL.n55 VTAIL.n54 9.3005
R456 VTAIL.n28 VTAIL.n27 9.3005
R457 VTAIL.n49 VTAIL.n48 9.3005
R458 VTAIL.n47 VTAIL.n46 9.3005
R459 VTAIL.n32 VTAIL.n31 9.3005
R460 VTAIL.n41 VTAIL.n40 9.3005
R461 VTAIL.n39 VTAIL.n38 9.3005
R462 VTAIL.n24 VTAIL.n23 9.3005
R463 VTAIL.n63 VTAIL.n62 9.3005
R464 VTAIL.n65 VTAIL.n64 9.3005
R465 VTAIL.n20 VTAIL.n19 9.3005
R466 VTAIL.n71 VTAIL.n70 9.3005
R467 VTAIL.n73 VTAIL.n72 9.3005
R468 VTAIL.n16 VTAIL.n15 9.3005
R469 VTAIL.n80 VTAIL.n79 9.3005
R470 VTAIL.n82 VTAIL.n81 9.3005
R471 VTAIL.n105 VTAIL.n104 9.3005
R472 VTAIL.n288 VTAIL.n287 9.3005
R473 VTAIL.n290 VTAIL.n289 9.3005
R474 VTAIL.n245 VTAIL.n244 9.3005
R475 VTAIL.n296 VTAIL.n295 9.3005
R476 VTAIL.n298 VTAIL.n297 9.3005
R477 VTAIL.n240 VTAIL.n239 9.3005
R478 VTAIL.n304 VTAIL.n303 9.3005
R479 VTAIL.n306 VTAIL.n305 9.3005
R480 VTAIL.n329 VTAIL.n328 9.3005
R481 VTAIL.n228 VTAIL.n227 9.3005
R482 VTAIL.n323 VTAIL.n322 9.3005
R483 VTAIL.n321 VTAIL.n320 9.3005
R484 VTAIL.n232 VTAIL.n231 9.3005
R485 VTAIL.n315 VTAIL.n314 9.3005
R486 VTAIL.n313 VTAIL.n312 9.3005
R487 VTAIL.n236 VTAIL.n235 9.3005
R488 VTAIL.n249 VTAIL.n248 9.3005
R489 VTAIL.n282 VTAIL.n281 9.3005
R490 VTAIL.n280 VTAIL.n279 9.3005
R491 VTAIL.n253 VTAIL.n252 9.3005
R492 VTAIL.n274 VTAIL.n273 9.3005
R493 VTAIL.n272 VTAIL.n271 9.3005
R494 VTAIL.n257 VTAIL.n256 9.3005
R495 VTAIL.n266 VTAIL.n265 9.3005
R496 VTAIL.n264 VTAIL.n263 9.3005
R497 VTAIL.n178 VTAIL.n177 9.3005
R498 VTAIL.n180 VTAIL.n179 9.3005
R499 VTAIL.n135 VTAIL.n134 9.3005
R500 VTAIL.n186 VTAIL.n185 9.3005
R501 VTAIL.n188 VTAIL.n187 9.3005
R502 VTAIL.n130 VTAIL.n129 9.3005
R503 VTAIL.n194 VTAIL.n193 9.3005
R504 VTAIL.n196 VTAIL.n195 9.3005
R505 VTAIL.n219 VTAIL.n218 9.3005
R506 VTAIL.n118 VTAIL.n117 9.3005
R507 VTAIL.n213 VTAIL.n212 9.3005
R508 VTAIL.n211 VTAIL.n210 9.3005
R509 VTAIL.n122 VTAIL.n121 9.3005
R510 VTAIL.n205 VTAIL.n204 9.3005
R511 VTAIL.n203 VTAIL.n202 9.3005
R512 VTAIL.n126 VTAIL.n125 9.3005
R513 VTAIL.n139 VTAIL.n138 9.3005
R514 VTAIL.n172 VTAIL.n171 9.3005
R515 VTAIL.n170 VTAIL.n169 9.3005
R516 VTAIL.n143 VTAIL.n142 9.3005
R517 VTAIL.n164 VTAIL.n163 9.3005
R518 VTAIL.n162 VTAIL.n161 9.3005
R519 VTAIL.n147 VTAIL.n146 9.3005
R520 VTAIL.n156 VTAIL.n155 9.3005
R521 VTAIL.n154 VTAIL.n153 9.3005
R522 VTAIL.n383 VTAIL.n358 8.92171
R523 VTAIL.n396 VTAIL.n350 8.92171
R524 VTAIL.n430 VTAIL.n429 8.92171
R525 VTAIL.n53 VTAIL.n28 8.92171
R526 VTAIL.n66 VTAIL.n20 8.92171
R527 VTAIL.n100 VTAIL.n99 8.92171
R528 VTAIL.n324 VTAIL.n323 8.92171
R529 VTAIL.n291 VTAIL.n245 8.92171
R530 VTAIL.n278 VTAIL.n253 8.92171
R531 VTAIL.n214 VTAIL.n213 8.92171
R532 VTAIL.n181 VTAIL.n135 8.92171
R533 VTAIL.n168 VTAIL.n143 8.92171
R534 VTAIL.n384 VTAIL.n356 8.14595
R535 VTAIL.n395 VTAIL.n352 8.14595
R536 VTAIL.n433 VTAIL.n334 8.14595
R537 VTAIL.n54 VTAIL.n26 8.14595
R538 VTAIL.n65 VTAIL.n22 8.14595
R539 VTAIL.n103 VTAIL.n4 8.14595
R540 VTAIL.n327 VTAIL.n228 8.14595
R541 VTAIL.n290 VTAIL.n247 8.14595
R542 VTAIL.n279 VTAIL.n251 8.14595
R543 VTAIL.n217 VTAIL.n118 8.14595
R544 VTAIL.n180 VTAIL.n137 8.14595
R545 VTAIL.n169 VTAIL.n141 8.14595
R546 VTAIL.n388 VTAIL.n387 7.3702
R547 VTAIL.n392 VTAIL.n391 7.3702
R548 VTAIL.n434 VTAIL.n332 7.3702
R549 VTAIL.n58 VTAIL.n57 7.3702
R550 VTAIL.n62 VTAIL.n61 7.3702
R551 VTAIL.n104 VTAIL.n2 7.3702
R552 VTAIL.n328 VTAIL.n226 7.3702
R553 VTAIL.n287 VTAIL.n286 7.3702
R554 VTAIL.n283 VTAIL.n282 7.3702
R555 VTAIL.n218 VTAIL.n116 7.3702
R556 VTAIL.n177 VTAIL.n176 7.3702
R557 VTAIL.n173 VTAIL.n172 7.3702
R558 VTAIL.n388 VTAIL.n354 6.59444
R559 VTAIL.n391 VTAIL.n354 6.59444
R560 VTAIL.n436 VTAIL.n332 6.59444
R561 VTAIL.n58 VTAIL.n24 6.59444
R562 VTAIL.n61 VTAIL.n24 6.59444
R563 VTAIL.n106 VTAIL.n2 6.59444
R564 VTAIL.n330 VTAIL.n226 6.59444
R565 VTAIL.n286 VTAIL.n249 6.59444
R566 VTAIL.n283 VTAIL.n249 6.59444
R567 VTAIL.n220 VTAIL.n116 6.59444
R568 VTAIL.n176 VTAIL.n139 6.59444
R569 VTAIL.n173 VTAIL.n139 6.59444
R570 VTAIL.n387 VTAIL.n356 5.81868
R571 VTAIL.n392 VTAIL.n352 5.81868
R572 VTAIL.n434 VTAIL.n433 5.81868
R573 VTAIL.n57 VTAIL.n26 5.81868
R574 VTAIL.n62 VTAIL.n22 5.81868
R575 VTAIL.n104 VTAIL.n103 5.81868
R576 VTAIL.n328 VTAIL.n327 5.81868
R577 VTAIL.n287 VTAIL.n247 5.81868
R578 VTAIL.n282 VTAIL.n251 5.81868
R579 VTAIL.n218 VTAIL.n217 5.81868
R580 VTAIL.n177 VTAIL.n137 5.81868
R581 VTAIL.n172 VTAIL.n141 5.81868
R582 VTAIL.n384 VTAIL.n383 5.04292
R583 VTAIL.n396 VTAIL.n395 5.04292
R584 VTAIL.n430 VTAIL.n334 5.04292
R585 VTAIL.n54 VTAIL.n53 5.04292
R586 VTAIL.n66 VTAIL.n65 5.04292
R587 VTAIL.n100 VTAIL.n4 5.04292
R588 VTAIL.n324 VTAIL.n228 5.04292
R589 VTAIL.n291 VTAIL.n290 5.04292
R590 VTAIL.n279 VTAIL.n278 5.04292
R591 VTAIL.n214 VTAIL.n118 5.04292
R592 VTAIL.n181 VTAIL.n180 5.04292
R593 VTAIL.n169 VTAIL.n168 5.04292
R594 VTAIL.n264 VTAIL.n260 4.38563
R595 VTAIL.n154 VTAIL.n150 4.38563
R596 VTAIL.n369 VTAIL.n365 4.38563
R597 VTAIL.n39 VTAIL.n35 4.38563
R598 VTAIL.n380 VTAIL.n358 4.26717
R599 VTAIL.n399 VTAIL.n350 4.26717
R600 VTAIL.n429 VTAIL.n336 4.26717
R601 VTAIL.n50 VTAIL.n28 4.26717
R602 VTAIL.n69 VTAIL.n20 4.26717
R603 VTAIL.n99 VTAIL.n6 4.26717
R604 VTAIL.n323 VTAIL.n230 4.26717
R605 VTAIL.n294 VTAIL.n245 4.26717
R606 VTAIL.n275 VTAIL.n253 4.26717
R607 VTAIL.n213 VTAIL.n120 4.26717
R608 VTAIL.n184 VTAIL.n135 4.26717
R609 VTAIL.n165 VTAIL.n143 4.26717
R610 VTAIL.n379 VTAIL.n360 3.49141
R611 VTAIL.n400 VTAIL.n348 3.49141
R612 VTAIL.n426 VTAIL.n425 3.49141
R613 VTAIL.n49 VTAIL.n30 3.49141
R614 VTAIL.n70 VTAIL.n18 3.49141
R615 VTAIL.n96 VTAIL.n95 3.49141
R616 VTAIL.n320 VTAIL.n319 3.49141
R617 VTAIL.n295 VTAIL.n243 3.49141
R618 VTAIL.n274 VTAIL.n255 3.49141
R619 VTAIL.n210 VTAIL.n209 3.49141
R620 VTAIL.n185 VTAIL.n133 3.49141
R621 VTAIL.n164 VTAIL.n145 3.49141
R622 VTAIL.n376 VTAIL.n375 2.71565
R623 VTAIL.n404 VTAIL.n403 2.71565
R624 VTAIL.n422 VTAIL.n338 2.71565
R625 VTAIL.n46 VTAIL.n45 2.71565
R626 VTAIL.n74 VTAIL.n73 2.71565
R627 VTAIL.n92 VTAIL.n8 2.71565
R628 VTAIL.n316 VTAIL.n232 2.71565
R629 VTAIL.n299 VTAIL.n298 2.71565
R630 VTAIL.n271 VTAIL.n270 2.71565
R631 VTAIL.n206 VTAIL.n122 2.71565
R632 VTAIL.n189 VTAIL.n188 2.71565
R633 VTAIL.n161 VTAIL.n160 2.71565
R634 VTAIL.n115 VTAIL.n113 2.32809
R635 VTAIL.n221 VTAIL.n115 2.32809
R636 VTAIL.n225 VTAIL.n223 2.32809
R637 VTAIL.n331 VTAIL.n225 2.32809
R638 VTAIL.n111 VTAIL.n109 2.32809
R639 VTAIL.n109 VTAIL.n107 2.32809
R640 VTAIL.n439 VTAIL.n437 2.32809
R641 VTAIL.n372 VTAIL.n362 1.93989
R642 VTAIL.n408 VTAIL.n346 1.93989
R643 VTAIL.n421 VTAIL.n340 1.93989
R644 VTAIL.n42 VTAIL.n32 1.93989
R645 VTAIL.n78 VTAIL.n16 1.93989
R646 VTAIL.n91 VTAIL.n10 1.93989
R647 VTAIL.n315 VTAIL.n234 1.93989
R648 VTAIL.n302 VTAIL.n240 1.93989
R649 VTAIL.n267 VTAIL.n257 1.93989
R650 VTAIL.n205 VTAIL.n124 1.93989
R651 VTAIL.n192 VTAIL.n130 1.93989
R652 VTAIL.n157 VTAIL.n147 1.93989
R653 VTAIL VTAIL.n1 1.80438
R654 VTAIL.n223 VTAIL.n221 1.63412
R655 VTAIL.n107 VTAIL.n1 1.63412
R656 VTAIL.n371 VTAIL.n364 1.16414
R657 VTAIL.n409 VTAIL.n344 1.16414
R658 VTAIL.n418 VTAIL.n417 1.16414
R659 VTAIL.n41 VTAIL.n34 1.16414
R660 VTAIL.n79 VTAIL.n14 1.16414
R661 VTAIL.n88 VTAIL.n87 1.16414
R662 VTAIL.n312 VTAIL.n311 1.16414
R663 VTAIL.n303 VTAIL.n238 1.16414
R664 VTAIL.n266 VTAIL.n259 1.16414
R665 VTAIL.n202 VTAIL.n201 1.16414
R666 VTAIL.n193 VTAIL.n128 1.16414
R667 VTAIL.n156 VTAIL.n149 1.16414
R668 VTAIL.n438 VTAIL.t16 1.0509
R669 VTAIL.n438 VTAIL.t12 1.0509
R670 VTAIL.n0 VTAIL.t13 1.0509
R671 VTAIL.n0 VTAIL.t14 1.0509
R672 VTAIL.n108 VTAIL.t0 1.0509
R673 VTAIL.n108 VTAIL.t8 1.0509
R674 VTAIL.n110 VTAIL.t5 1.0509
R675 VTAIL.n110 VTAIL.t3 1.0509
R676 VTAIL.n224 VTAIL.t4 1.0509
R677 VTAIL.n224 VTAIL.t6 1.0509
R678 VTAIL.n222 VTAIL.t1 1.0509
R679 VTAIL.n222 VTAIL.t2 1.0509
R680 VTAIL.n114 VTAIL.t17 1.0509
R681 VTAIL.n114 VTAIL.t19 1.0509
R682 VTAIL.n112 VTAIL.t10 1.0509
R683 VTAIL.n112 VTAIL.t15 1.0509
R684 VTAIL VTAIL.n439 0.524207
R685 VTAIL.n368 VTAIL.n367 0.388379
R686 VTAIL.n413 VTAIL.n412 0.388379
R687 VTAIL.n414 VTAIL.n342 0.388379
R688 VTAIL.n38 VTAIL.n37 0.388379
R689 VTAIL.n83 VTAIL.n82 0.388379
R690 VTAIL.n84 VTAIL.n12 0.388379
R691 VTAIL.n308 VTAIL.n236 0.388379
R692 VTAIL.n307 VTAIL.n306 0.388379
R693 VTAIL.n263 VTAIL.n262 0.388379
R694 VTAIL.n198 VTAIL.n126 0.388379
R695 VTAIL.n197 VTAIL.n196 0.388379
R696 VTAIL.n153 VTAIL.n152 0.388379
R697 VTAIL.n370 VTAIL.n369 0.155672
R698 VTAIL.n370 VTAIL.n361 0.155672
R699 VTAIL.n377 VTAIL.n361 0.155672
R700 VTAIL.n378 VTAIL.n377 0.155672
R701 VTAIL.n378 VTAIL.n357 0.155672
R702 VTAIL.n385 VTAIL.n357 0.155672
R703 VTAIL.n386 VTAIL.n385 0.155672
R704 VTAIL.n386 VTAIL.n353 0.155672
R705 VTAIL.n393 VTAIL.n353 0.155672
R706 VTAIL.n394 VTAIL.n393 0.155672
R707 VTAIL.n394 VTAIL.n349 0.155672
R708 VTAIL.n401 VTAIL.n349 0.155672
R709 VTAIL.n402 VTAIL.n401 0.155672
R710 VTAIL.n402 VTAIL.n345 0.155672
R711 VTAIL.n410 VTAIL.n345 0.155672
R712 VTAIL.n411 VTAIL.n410 0.155672
R713 VTAIL.n411 VTAIL.n341 0.155672
R714 VTAIL.n419 VTAIL.n341 0.155672
R715 VTAIL.n420 VTAIL.n419 0.155672
R716 VTAIL.n420 VTAIL.n337 0.155672
R717 VTAIL.n427 VTAIL.n337 0.155672
R718 VTAIL.n428 VTAIL.n427 0.155672
R719 VTAIL.n428 VTAIL.n333 0.155672
R720 VTAIL.n435 VTAIL.n333 0.155672
R721 VTAIL.n40 VTAIL.n39 0.155672
R722 VTAIL.n40 VTAIL.n31 0.155672
R723 VTAIL.n47 VTAIL.n31 0.155672
R724 VTAIL.n48 VTAIL.n47 0.155672
R725 VTAIL.n48 VTAIL.n27 0.155672
R726 VTAIL.n55 VTAIL.n27 0.155672
R727 VTAIL.n56 VTAIL.n55 0.155672
R728 VTAIL.n56 VTAIL.n23 0.155672
R729 VTAIL.n63 VTAIL.n23 0.155672
R730 VTAIL.n64 VTAIL.n63 0.155672
R731 VTAIL.n64 VTAIL.n19 0.155672
R732 VTAIL.n71 VTAIL.n19 0.155672
R733 VTAIL.n72 VTAIL.n71 0.155672
R734 VTAIL.n72 VTAIL.n15 0.155672
R735 VTAIL.n80 VTAIL.n15 0.155672
R736 VTAIL.n81 VTAIL.n80 0.155672
R737 VTAIL.n81 VTAIL.n11 0.155672
R738 VTAIL.n89 VTAIL.n11 0.155672
R739 VTAIL.n90 VTAIL.n89 0.155672
R740 VTAIL.n90 VTAIL.n7 0.155672
R741 VTAIL.n97 VTAIL.n7 0.155672
R742 VTAIL.n98 VTAIL.n97 0.155672
R743 VTAIL.n98 VTAIL.n3 0.155672
R744 VTAIL.n105 VTAIL.n3 0.155672
R745 VTAIL.n329 VTAIL.n227 0.155672
R746 VTAIL.n322 VTAIL.n227 0.155672
R747 VTAIL.n322 VTAIL.n321 0.155672
R748 VTAIL.n321 VTAIL.n231 0.155672
R749 VTAIL.n314 VTAIL.n231 0.155672
R750 VTAIL.n314 VTAIL.n313 0.155672
R751 VTAIL.n313 VTAIL.n235 0.155672
R752 VTAIL.n305 VTAIL.n235 0.155672
R753 VTAIL.n305 VTAIL.n304 0.155672
R754 VTAIL.n304 VTAIL.n239 0.155672
R755 VTAIL.n297 VTAIL.n239 0.155672
R756 VTAIL.n297 VTAIL.n296 0.155672
R757 VTAIL.n296 VTAIL.n244 0.155672
R758 VTAIL.n289 VTAIL.n244 0.155672
R759 VTAIL.n289 VTAIL.n288 0.155672
R760 VTAIL.n288 VTAIL.n248 0.155672
R761 VTAIL.n281 VTAIL.n248 0.155672
R762 VTAIL.n281 VTAIL.n280 0.155672
R763 VTAIL.n280 VTAIL.n252 0.155672
R764 VTAIL.n273 VTAIL.n252 0.155672
R765 VTAIL.n273 VTAIL.n272 0.155672
R766 VTAIL.n272 VTAIL.n256 0.155672
R767 VTAIL.n265 VTAIL.n256 0.155672
R768 VTAIL.n265 VTAIL.n264 0.155672
R769 VTAIL.n219 VTAIL.n117 0.155672
R770 VTAIL.n212 VTAIL.n117 0.155672
R771 VTAIL.n212 VTAIL.n211 0.155672
R772 VTAIL.n211 VTAIL.n121 0.155672
R773 VTAIL.n204 VTAIL.n121 0.155672
R774 VTAIL.n204 VTAIL.n203 0.155672
R775 VTAIL.n203 VTAIL.n125 0.155672
R776 VTAIL.n195 VTAIL.n125 0.155672
R777 VTAIL.n195 VTAIL.n194 0.155672
R778 VTAIL.n194 VTAIL.n129 0.155672
R779 VTAIL.n187 VTAIL.n129 0.155672
R780 VTAIL.n187 VTAIL.n186 0.155672
R781 VTAIL.n186 VTAIL.n134 0.155672
R782 VTAIL.n179 VTAIL.n134 0.155672
R783 VTAIL.n179 VTAIL.n178 0.155672
R784 VTAIL.n178 VTAIL.n138 0.155672
R785 VTAIL.n171 VTAIL.n138 0.155672
R786 VTAIL.n171 VTAIL.n170 0.155672
R787 VTAIL.n170 VTAIL.n142 0.155672
R788 VTAIL.n163 VTAIL.n142 0.155672
R789 VTAIL.n163 VTAIL.n162 0.155672
R790 VTAIL.n162 VTAIL.n146 0.155672
R791 VTAIL.n155 VTAIL.n146 0.155672
R792 VTAIL.n155 VTAIL.n154 0.155672
R793 VDD2.n209 VDD2.n109 289.615
R794 VDD2.n100 VDD2.n0 289.615
R795 VDD2.n210 VDD2.n209 185
R796 VDD2.n208 VDD2.n207 185
R797 VDD2.n113 VDD2.n112 185
R798 VDD2.n202 VDD2.n201 185
R799 VDD2.n200 VDD2.n199 185
R800 VDD2.n117 VDD2.n116 185
R801 VDD2.n194 VDD2.n193 185
R802 VDD2.n192 VDD2.n191 185
R803 VDD2.n190 VDD2.n120 185
R804 VDD2.n124 VDD2.n121 185
R805 VDD2.n185 VDD2.n184 185
R806 VDD2.n183 VDD2.n182 185
R807 VDD2.n126 VDD2.n125 185
R808 VDD2.n177 VDD2.n176 185
R809 VDD2.n175 VDD2.n174 185
R810 VDD2.n130 VDD2.n129 185
R811 VDD2.n169 VDD2.n168 185
R812 VDD2.n167 VDD2.n166 185
R813 VDD2.n134 VDD2.n133 185
R814 VDD2.n161 VDD2.n160 185
R815 VDD2.n159 VDD2.n158 185
R816 VDD2.n138 VDD2.n137 185
R817 VDD2.n153 VDD2.n152 185
R818 VDD2.n151 VDD2.n150 185
R819 VDD2.n142 VDD2.n141 185
R820 VDD2.n145 VDD2.n144 185
R821 VDD2.n35 VDD2.n34 185
R822 VDD2.n32 VDD2.n31 185
R823 VDD2.n41 VDD2.n40 185
R824 VDD2.n43 VDD2.n42 185
R825 VDD2.n28 VDD2.n27 185
R826 VDD2.n49 VDD2.n48 185
R827 VDD2.n51 VDD2.n50 185
R828 VDD2.n24 VDD2.n23 185
R829 VDD2.n57 VDD2.n56 185
R830 VDD2.n59 VDD2.n58 185
R831 VDD2.n20 VDD2.n19 185
R832 VDD2.n65 VDD2.n64 185
R833 VDD2.n67 VDD2.n66 185
R834 VDD2.n16 VDD2.n15 185
R835 VDD2.n73 VDD2.n72 185
R836 VDD2.n76 VDD2.n75 185
R837 VDD2.n74 VDD2.n12 185
R838 VDD2.n81 VDD2.n11 185
R839 VDD2.n83 VDD2.n82 185
R840 VDD2.n85 VDD2.n84 185
R841 VDD2.n8 VDD2.n7 185
R842 VDD2.n91 VDD2.n90 185
R843 VDD2.n93 VDD2.n92 185
R844 VDD2.n4 VDD2.n3 185
R845 VDD2.n99 VDD2.n98 185
R846 VDD2.n101 VDD2.n100 185
R847 VDD2.t2 VDD2.n143 147.659
R848 VDD2.t0 VDD2.n33 147.659
R849 VDD2.n209 VDD2.n208 104.615
R850 VDD2.n208 VDD2.n112 104.615
R851 VDD2.n201 VDD2.n112 104.615
R852 VDD2.n201 VDD2.n200 104.615
R853 VDD2.n200 VDD2.n116 104.615
R854 VDD2.n193 VDD2.n116 104.615
R855 VDD2.n193 VDD2.n192 104.615
R856 VDD2.n192 VDD2.n120 104.615
R857 VDD2.n124 VDD2.n120 104.615
R858 VDD2.n184 VDD2.n124 104.615
R859 VDD2.n184 VDD2.n183 104.615
R860 VDD2.n183 VDD2.n125 104.615
R861 VDD2.n176 VDD2.n125 104.615
R862 VDD2.n176 VDD2.n175 104.615
R863 VDD2.n175 VDD2.n129 104.615
R864 VDD2.n168 VDD2.n129 104.615
R865 VDD2.n168 VDD2.n167 104.615
R866 VDD2.n167 VDD2.n133 104.615
R867 VDD2.n160 VDD2.n133 104.615
R868 VDD2.n160 VDD2.n159 104.615
R869 VDD2.n159 VDD2.n137 104.615
R870 VDD2.n152 VDD2.n137 104.615
R871 VDD2.n152 VDD2.n151 104.615
R872 VDD2.n151 VDD2.n141 104.615
R873 VDD2.n144 VDD2.n141 104.615
R874 VDD2.n34 VDD2.n31 104.615
R875 VDD2.n41 VDD2.n31 104.615
R876 VDD2.n42 VDD2.n41 104.615
R877 VDD2.n42 VDD2.n27 104.615
R878 VDD2.n49 VDD2.n27 104.615
R879 VDD2.n50 VDD2.n49 104.615
R880 VDD2.n50 VDD2.n23 104.615
R881 VDD2.n57 VDD2.n23 104.615
R882 VDD2.n58 VDD2.n57 104.615
R883 VDD2.n58 VDD2.n19 104.615
R884 VDD2.n65 VDD2.n19 104.615
R885 VDD2.n66 VDD2.n65 104.615
R886 VDD2.n66 VDD2.n15 104.615
R887 VDD2.n73 VDD2.n15 104.615
R888 VDD2.n75 VDD2.n73 104.615
R889 VDD2.n75 VDD2.n74 104.615
R890 VDD2.n74 VDD2.n11 104.615
R891 VDD2.n83 VDD2.n11 104.615
R892 VDD2.n84 VDD2.n83 104.615
R893 VDD2.n84 VDD2.n7 104.615
R894 VDD2.n91 VDD2.n7 104.615
R895 VDD2.n92 VDD2.n91 104.615
R896 VDD2.n92 VDD2.n3 104.615
R897 VDD2.n99 VDD2.n3 104.615
R898 VDD2.n100 VDD2.n99 104.615
R899 VDD2.n108 VDD2.n107 60.179
R900 VDD2 VDD2.n217 60.176
R901 VDD2.n216 VDD2.n215 58.4887
R902 VDD2.n106 VDD2.n105 58.4887
R903 VDD2.n144 VDD2.t2 52.3082
R904 VDD2.n34 VDD2.t0 52.3082
R905 VDD2.n214 VDD2.n108 51.0213
R906 VDD2.n106 VDD2.n104 49.0584
R907 VDD2.n214 VDD2.n213 46.7308
R908 VDD2.n145 VDD2.n143 15.6677
R909 VDD2.n35 VDD2.n33 15.6677
R910 VDD2.n191 VDD2.n190 13.1884
R911 VDD2.n82 VDD2.n81 13.1884
R912 VDD2.n194 VDD2.n119 12.8005
R913 VDD2.n189 VDD2.n121 12.8005
R914 VDD2.n146 VDD2.n142 12.8005
R915 VDD2.n36 VDD2.n32 12.8005
R916 VDD2.n80 VDD2.n12 12.8005
R917 VDD2.n85 VDD2.n10 12.8005
R918 VDD2.n195 VDD2.n117 12.0247
R919 VDD2.n186 VDD2.n185 12.0247
R920 VDD2.n150 VDD2.n149 12.0247
R921 VDD2.n40 VDD2.n39 12.0247
R922 VDD2.n77 VDD2.n76 12.0247
R923 VDD2.n86 VDD2.n8 12.0247
R924 VDD2.n199 VDD2.n198 11.249
R925 VDD2.n182 VDD2.n123 11.249
R926 VDD2.n153 VDD2.n140 11.249
R927 VDD2.n43 VDD2.n30 11.249
R928 VDD2.n72 VDD2.n14 11.249
R929 VDD2.n90 VDD2.n89 11.249
R930 VDD2.n202 VDD2.n115 10.4732
R931 VDD2.n181 VDD2.n126 10.4732
R932 VDD2.n154 VDD2.n138 10.4732
R933 VDD2.n44 VDD2.n28 10.4732
R934 VDD2.n71 VDD2.n16 10.4732
R935 VDD2.n93 VDD2.n6 10.4732
R936 VDD2.n203 VDD2.n113 9.69747
R937 VDD2.n178 VDD2.n177 9.69747
R938 VDD2.n158 VDD2.n157 9.69747
R939 VDD2.n48 VDD2.n47 9.69747
R940 VDD2.n68 VDD2.n67 9.69747
R941 VDD2.n94 VDD2.n4 9.69747
R942 VDD2.n213 VDD2.n212 9.45567
R943 VDD2.n104 VDD2.n103 9.45567
R944 VDD2.n171 VDD2.n170 9.3005
R945 VDD2.n173 VDD2.n172 9.3005
R946 VDD2.n128 VDD2.n127 9.3005
R947 VDD2.n179 VDD2.n178 9.3005
R948 VDD2.n181 VDD2.n180 9.3005
R949 VDD2.n123 VDD2.n122 9.3005
R950 VDD2.n187 VDD2.n186 9.3005
R951 VDD2.n189 VDD2.n188 9.3005
R952 VDD2.n212 VDD2.n211 9.3005
R953 VDD2.n111 VDD2.n110 9.3005
R954 VDD2.n206 VDD2.n205 9.3005
R955 VDD2.n204 VDD2.n203 9.3005
R956 VDD2.n115 VDD2.n114 9.3005
R957 VDD2.n198 VDD2.n197 9.3005
R958 VDD2.n196 VDD2.n195 9.3005
R959 VDD2.n119 VDD2.n118 9.3005
R960 VDD2.n132 VDD2.n131 9.3005
R961 VDD2.n165 VDD2.n164 9.3005
R962 VDD2.n163 VDD2.n162 9.3005
R963 VDD2.n136 VDD2.n135 9.3005
R964 VDD2.n157 VDD2.n156 9.3005
R965 VDD2.n155 VDD2.n154 9.3005
R966 VDD2.n140 VDD2.n139 9.3005
R967 VDD2.n149 VDD2.n148 9.3005
R968 VDD2.n147 VDD2.n146 9.3005
R969 VDD2.n2 VDD2.n1 9.3005
R970 VDD2.n97 VDD2.n96 9.3005
R971 VDD2.n95 VDD2.n94 9.3005
R972 VDD2.n6 VDD2.n5 9.3005
R973 VDD2.n89 VDD2.n88 9.3005
R974 VDD2.n87 VDD2.n86 9.3005
R975 VDD2.n10 VDD2.n9 9.3005
R976 VDD2.n55 VDD2.n54 9.3005
R977 VDD2.n53 VDD2.n52 9.3005
R978 VDD2.n26 VDD2.n25 9.3005
R979 VDD2.n47 VDD2.n46 9.3005
R980 VDD2.n45 VDD2.n44 9.3005
R981 VDD2.n30 VDD2.n29 9.3005
R982 VDD2.n39 VDD2.n38 9.3005
R983 VDD2.n37 VDD2.n36 9.3005
R984 VDD2.n22 VDD2.n21 9.3005
R985 VDD2.n61 VDD2.n60 9.3005
R986 VDD2.n63 VDD2.n62 9.3005
R987 VDD2.n18 VDD2.n17 9.3005
R988 VDD2.n69 VDD2.n68 9.3005
R989 VDD2.n71 VDD2.n70 9.3005
R990 VDD2.n14 VDD2.n13 9.3005
R991 VDD2.n78 VDD2.n77 9.3005
R992 VDD2.n80 VDD2.n79 9.3005
R993 VDD2.n103 VDD2.n102 9.3005
R994 VDD2.n207 VDD2.n206 8.92171
R995 VDD2.n174 VDD2.n128 8.92171
R996 VDD2.n161 VDD2.n136 8.92171
R997 VDD2.n51 VDD2.n26 8.92171
R998 VDD2.n64 VDD2.n18 8.92171
R999 VDD2.n98 VDD2.n97 8.92171
R1000 VDD2.n210 VDD2.n111 8.14595
R1001 VDD2.n173 VDD2.n130 8.14595
R1002 VDD2.n162 VDD2.n134 8.14595
R1003 VDD2.n52 VDD2.n24 8.14595
R1004 VDD2.n63 VDD2.n20 8.14595
R1005 VDD2.n101 VDD2.n2 8.14595
R1006 VDD2.n211 VDD2.n109 7.3702
R1007 VDD2.n170 VDD2.n169 7.3702
R1008 VDD2.n166 VDD2.n165 7.3702
R1009 VDD2.n56 VDD2.n55 7.3702
R1010 VDD2.n60 VDD2.n59 7.3702
R1011 VDD2.n102 VDD2.n0 7.3702
R1012 VDD2.n213 VDD2.n109 6.59444
R1013 VDD2.n169 VDD2.n132 6.59444
R1014 VDD2.n166 VDD2.n132 6.59444
R1015 VDD2.n56 VDD2.n22 6.59444
R1016 VDD2.n59 VDD2.n22 6.59444
R1017 VDD2.n104 VDD2.n0 6.59444
R1018 VDD2.n211 VDD2.n210 5.81868
R1019 VDD2.n170 VDD2.n130 5.81868
R1020 VDD2.n165 VDD2.n134 5.81868
R1021 VDD2.n55 VDD2.n24 5.81868
R1022 VDD2.n60 VDD2.n20 5.81868
R1023 VDD2.n102 VDD2.n101 5.81868
R1024 VDD2.n207 VDD2.n111 5.04292
R1025 VDD2.n174 VDD2.n173 5.04292
R1026 VDD2.n162 VDD2.n161 5.04292
R1027 VDD2.n52 VDD2.n51 5.04292
R1028 VDD2.n64 VDD2.n63 5.04292
R1029 VDD2.n98 VDD2.n2 5.04292
R1030 VDD2.n147 VDD2.n143 4.38563
R1031 VDD2.n37 VDD2.n33 4.38563
R1032 VDD2.n206 VDD2.n113 4.26717
R1033 VDD2.n177 VDD2.n128 4.26717
R1034 VDD2.n158 VDD2.n136 4.26717
R1035 VDD2.n48 VDD2.n26 4.26717
R1036 VDD2.n67 VDD2.n18 4.26717
R1037 VDD2.n97 VDD2.n4 4.26717
R1038 VDD2.n203 VDD2.n202 3.49141
R1039 VDD2.n178 VDD2.n126 3.49141
R1040 VDD2.n157 VDD2.n138 3.49141
R1041 VDD2.n47 VDD2.n28 3.49141
R1042 VDD2.n68 VDD2.n16 3.49141
R1043 VDD2.n94 VDD2.n93 3.49141
R1044 VDD2.n199 VDD2.n115 2.71565
R1045 VDD2.n182 VDD2.n181 2.71565
R1046 VDD2.n154 VDD2.n153 2.71565
R1047 VDD2.n44 VDD2.n43 2.71565
R1048 VDD2.n72 VDD2.n71 2.71565
R1049 VDD2.n90 VDD2.n6 2.71565
R1050 VDD2.n216 VDD2.n214 2.32809
R1051 VDD2.n198 VDD2.n117 1.93989
R1052 VDD2.n185 VDD2.n123 1.93989
R1053 VDD2.n150 VDD2.n140 1.93989
R1054 VDD2.n40 VDD2.n30 1.93989
R1055 VDD2.n76 VDD2.n14 1.93989
R1056 VDD2.n89 VDD2.n8 1.93989
R1057 VDD2.n195 VDD2.n194 1.16414
R1058 VDD2.n186 VDD2.n121 1.16414
R1059 VDD2.n149 VDD2.n142 1.16414
R1060 VDD2.n39 VDD2.n32 1.16414
R1061 VDD2.n77 VDD2.n12 1.16414
R1062 VDD2.n86 VDD2.n85 1.16414
R1063 VDD2.n217 VDD2.t8 1.0509
R1064 VDD2.n217 VDD2.t4 1.0509
R1065 VDD2.n215 VDD2.t7 1.0509
R1066 VDD2.n215 VDD2.t1 1.0509
R1067 VDD2.n107 VDD2.t3 1.0509
R1068 VDD2.n107 VDD2.t6 1.0509
R1069 VDD2.n105 VDD2.t5 1.0509
R1070 VDD2.n105 VDD2.t9 1.0509
R1071 VDD2 VDD2.n216 0.640586
R1072 VDD2.n108 VDD2.n106 0.527051
R1073 VDD2.n191 VDD2.n119 0.388379
R1074 VDD2.n190 VDD2.n189 0.388379
R1075 VDD2.n146 VDD2.n145 0.388379
R1076 VDD2.n36 VDD2.n35 0.388379
R1077 VDD2.n81 VDD2.n80 0.388379
R1078 VDD2.n82 VDD2.n10 0.388379
R1079 VDD2.n212 VDD2.n110 0.155672
R1080 VDD2.n205 VDD2.n110 0.155672
R1081 VDD2.n205 VDD2.n204 0.155672
R1082 VDD2.n204 VDD2.n114 0.155672
R1083 VDD2.n197 VDD2.n114 0.155672
R1084 VDD2.n197 VDD2.n196 0.155672
R1085 VDD2.n196 VDD2.n118 0.155672
R1086 VDD2.n188 VDD2.n118 0.155672
R1087 VDD2.n188 VDD2.n187 0.155672
R1088 VDD2.n187 VDD2.n122 0.155672
R1089 VDD2.n180 VDD2.n122 0.155672
R1090 VDD2.n180 VDD2.n179 0.155672
R1091 VDD2.n179 VDD2.n127 0.155672
R1092 VDD2.n172 VDD2.n127 0.155672
R1093 VDD2.n172 VDD2.n171 0.155672
R1094 VDD2.n171 VDD2.n131 0.155672
R1095 VDD2.n164 VDD2.n131 0.155672
R1096 VDD2.n164 VDD2.n163 0.155672
R1097 VDD2.n163 VDD2.n135 0.155672
R1098 VDD2.n156 VDD2.n135 0.155672
R1099 VDD2.n156 VDD2.n155 0.155672
R1100 VDD2.n155 VDD2.n139 0.155672
R1101 VDD2.n148 VDD2.n139 0.155672
R1102 VDD2.n148 VDD2.n147 0.155672
R1103 VDD2.n38 VDD2.n37 0.155672
R1104 VDD2.n38 VDD2.n29 0.155672
R1105 VDD2.n45 VDD2.n29 0.155672
R1106 VDD2.n46 VDD2.n45 0.155672
R1107 VDD2.n46 VDD2.n25 0.155672
R1108 VDD2.n53 VDD2.n25 0.155672
R1109 VDD2.n54 VDD2.n53 0.155672
R1110 VDD2.n54 VDD2.n21 0.155672
R1111 VDD2.n61 VDD2.n21 0.155672
R1112 VDD2.n62 VDD2.n61 0.155672
R1113 VDD2.n62 VDD2.n17 0.155672
R1114 VDD2.n69 VDD2.n17 0.155672
R1115 VDD2.n70 VDD2.n69 0.155672
R1116 VDD2.n70 VDD2.n13 0.155672
R1117 VDD2.n78 VDD2.n13 0.155672
R1118 VDD2.n79 VDD2.n78 0.155672
R1119 VDD2.n79 VDD2.n9 0.155672
R1120 VDD2.n87 VDD2.n9 0.155672
R1121 VDD2.n88 VDD2.n87 0.155672
R1122 VDD2.n88 VDD2.n5 0.155672
R1123 VDD2.n95 VDD2.n5 0.155672
R1124 VDD2.n96 VDD2.n95 0.155672
R1125 VDD2.n96 VDD2.n1 0.155672
R1126 VDD2.n103 VDD2.n1 0.155672
R1127 B.n1119 B.n1118 585
R1128 B.n1120 B.n1119 585
R1129 B.n435 B.n169 585
R1130 B.n434 B.n433 585
R1131 B.n432 B.n431 585
R1132 B.n430 B.n429 585
R1133 B.n428 B.n427 585
R1134 B.n426 B.n425 585
R1135 B.n424 B.n423 585
R1136 B.n422 B.n421 585
R1137 B.n420 B.n419 585
R1138 B.n418 B.n417 585
R1139 B.n416 B.n415 585
R1140 B.n414 B.n413 585
R1141 B.n412 B.n411 585
R1142 B.n410 B.n409 585
R1143 B.n408 B.n407 585
R1144 B.n406 B.n405 585
R1145 B.n404 B.n403 585
R1146 B.n402 B.n401 585
R1147 B.n400 B.n399 585
R1148 B.n398 B.n397 585
R1149 B.n396 B.n395 585
R1150 B.n394 B.n393 585
R1151 B.n392 B.n391 585
R1152 B.n390 B.n389 585
R1153 B.n388 B.n387 585
R1154 B.n386 B.n385 585
R1155 B.n384 B.n383 585
R1156 B.n382 B.n381 585
R1157 B.n380 B.n379 585
R1158 B.n378 B.n377 585
R1159 B.n376 B.n375 585
R1160 B.n374 B.n373 585
R1161 B.n372 B.n371 585
R1162 B.n370 B.n369 585
R1163 B.n368 B.n367 585
R1164 B.n366 B.n365 585
R1165 B.n364 B.n363 585
R1166 B.n362 B.n361 585
R1167 B.n360 B.n359 585
R1168 B.n358 B.n357 585
R1169 B.n356 B.n355 585
R1170 B.n354 B.n353 585
R1171 B.n352 B.n351 585
R1172 B.n350 B.n349 585
R1173 B.n348 B.n347 585
R1174 B.n346 B.n345 585
R1175 B.n344 B.n343 585
R1176 B.n342 B.n341 585
R1177 B.n340 B.n339 585
R1178 B.n338 B.n337 585
R1179 B.n336 B.n335 585
R1180 B.n334 B.n333 585
R1181 B.n332 B.n331 585
R1182 B.n330 B.n329 585
R1183 B.n328 B.n327 585
R1184 B.n326 B.n325 585
R1185 B.n324 B.n323 585
R1186 B.n322 B.n321 585
R1187 B.n320 B.n319 585
R1188 B.n318 B.n317 585
R1189 B.n316 B.n315 585
R1190 B.n313 B.n312 585
R1191 B.n311 B.n310 585
R1192 B.n309 B.n308 585
R1193 B.n307 B.n306 585
R1194 B.n305 B.n304 585
R1195 B.n303 B.n302 585
R1196 B.n301 B.n300 585
R1197 B.n299 B.n298 585
R1198 B.n297 B.n296 585
R1199 B.n295 B.n294 585
R1200 B.n293 B.n292 585
R1201 B.n291 B.n290 585
R1202 B.n289 B.n288 585
R1203 B.n287 B.n286 585
R1204 B.n285 B.n284 585
R1205 B.n283 B.n282 585
R1206 B.n281 B.n280 585
R1207 B.n279 B.n278 585
R1208 B.n277 B.n276 585
R1209 B.n275 B.n274 585
R1210 B.n273 B.n272 585
R1211 B.n271 B.n270 585
R1212 B.n269 B.n268 585
R1213 B.n267 B.n266 585
R1214 B.n265 B.n264 585
R1215 B.n263 B.n262 585
R1216 B.n261 B.n260 585
R1217 B.n259 B.n258 585
R1218 B.n257 B.n256 585
R1219 B.n255 B.n254 585
R1220 B.n253 B.n252 585
R1221 B.n251 B.n250 585
R1222 B.n249 B.n248 585
R1223 B.n247 B.n246 585
R1224 B.n245 B.n244 585
R1225 B.n243 B.n242 585
R1226 B.n241 B.n240 585
R1227 B.n239 B.n238 585
R1228 B.n237 B.n236 585
R1229 B.n235 B.n234 585
R1230 B.n233 B.n232 585
R1231 B.n231 B.n230 585
R1232 B.n229 B.n228 585
R1233 B.n227 B.n226 585
R1234 B.n225 B.n224 585
R1235 B.n223 B.n222 585
R1236 B.n221 B.n220 585
R1237 B.n219 B.n218 585
R1238 B.n217 B.n216 585
R1239 B.n215 B.n214 585
R1240 B.n213 B.n212 585
R1241 B.n211 B.n210 585
R1242 B.n209 B.n208 585
R1243 B.n207 B.n206 585
R1244 B.n205 B.n204 585
R1245 B.n203 B.n202 585
R1246 B.n201 B.n200 585
R1247 B.n199 B.n198 585
R1248 B.n197 B.n196 585
R1249 B.n195 B.n194 585
R1250 B.n193 B.n192 585
R1251 B.n191 B.n190 585
R1252 B.n189 B.n188 585
R1253 B.n187 B.n186 585
R1254 B.n185 B.n184 585
R1255 B.n183 B.n182 585
R1256 B.n181 B.n180 585
R1257 B.n179 B.n178 585
R1258 B.n177 B.n176 585
R1259 B.n103 B.n102 585
R1260 B.n1123 B.n1122 585
R1261 B.n1117 B.n170 585
R1262 B.n170 B.n100 585
R1263 B.n1116 B.n99 585
R1264 B.n1127 B.n99 585
R1265 B.n1115 B.n98 585
R1266 B.n1128 B.n98 585
R1267 B.n1114 B.n97 585
R1268 B.n1129 B.n97 585
R1269 B.n1113 B.n1112 585
R1270 B.n1112 B.n93 585
R1271 B.n1111 B.n92 585
R1272 B.n1135 B.n92 585
R1273 B.n1110 B.n91 585
R1274 B.n1136 B.n91 585
R1275 B.n1109 B.n90 585
R1276 B.n1137 B.n90 585
R1277 B.n1108 B.n1107 585
R1278 B.n1107 B.n86 585
R1279 B.n1106 B.n85 585
R1280 B.n1143 B.n85 585
R1281 B.n1105 B.n84 585
R1282 B.n1144 B.n84 585
R1283 B.n1104 B.n83 585
R1284 B.n1145 B.n83 585
R1285 B.n1103 B.n1102 585
R1286 B.n1102 B.n79 585
R1287 B.n1101 B.n78 585
R1288 B.n1151 B.n78 585
R1289 B.n1100 B.n77 585
R1290 B.n1152 B.n77 585
R1291 B.n1099 B.n76 585
R1292 B.n1153 B.n76 585
R1293 B.n1098 B.n1097 585
R1294 B.n1097 B.n72 585
R1295 B.n1096 B.n71 585
R1296 B.n1159 B.n71 585
R1297 B.n1095 B.n70 585
R1298 B.n1160 B.n70 585
R1299 B.n1094 B.n69 585
R1300 B.n1161 B.n69 585
R1301 B.n1093 B.n1092 585
R1302 B.n1092 B.n65 585
R1303 B.n1091 B.n64 585
R1304 B.n1167 B.n64 585
R1305 B.n1090 B.n63 585
R1306 B.n1168 B.n63 585
R1307 B.n1089 B.n62 585
R1308 B.n1169 B.n62 585
R1309 B.n1088 B.n1087 585
R1310 B.n1087 B.n58 585
R1311 B.n1086 B.n57 585
R1312 B.n1175 B.n57 585
R1313 B.n1085 B.n56 585
R1314 B.n1176 B.n56 585
R1315 B.n1084 B.n55 585
R1316 B.n1177 B.n55 585
R1317 B.n1083 B.n1082 585
R1318 B.n1082 B.n51 585
R1319 B.n1081 B.n50 585
R1320 B.n1183 B.n50 585
R1321 B.n1080 B.n49 585
R1322 B.n1184 B.n49 585
R1323 B.n1079 B.n48 585
R1324 B.n1185 B.n48 585
R1325 B.n1078 B.n1077 585
R1326 B.n1077 B.n44 585
R1327 B.n1076 B.n43 585
R1328 B.n1191 B.n43 585
R1329 B.n1075 B.n42 585
R1330 B.n1192 B.n42 585
R1331 B.n1074 B.n41 585
R1332 B.n1193 B.n41 585
R1333 B.n1073 B.n1072 585
R1334 B.n1072 B.n37 585
R1335 B.n1071 B.n36 585
R1336 B.n1199 B.n36 585
R1337 B.n1070 B.n35 585
R1338 B.n1200 B.n35 585
R1339 B.n1069 B.n34 585
R1340 B.n1201 B.n34 585
R1341 B.n1068 B.n1067 585
R1342 B.n1067 B.n30 585
R1343 B.n1066 B.n29 585
R1344 B.n1207 B.n29 585
R1345 B.n1065 B.n28 585
R1346 B.n1208 B.n28 585
R1347 B.n1064 B.n27 585
R1348 B.n1209 B.n27 585
R1349 B.n1063 B.n1062 585
R1350 B.n1062 B.n23 585
R1351 B.n1061 B.n22 585
R1352 B.n1215 B.n22 585
R1353 B.n1060 B.n21 585
R1354 B.n1216 B.n21 585
R1355 B.n1059 B.n20 585
R1356 B.n1217 B.n20 585
R1357 B.n1058 B.n1057 585
R1358 B.n1057 B.n16 585
R1359 B.n1056 B.n15 585
R1360 B.n1223 B.n15 585
R1361 B.n1055 B.n14 585
R1362 B.n1224 B.n14 585
R1363 B.n1054 B.n13 585
R1364 B.n1225 B.n13 585
R1365 B.n1053 B.n1052 585
R1366 B.n1052 B.n12 585
R1367 B.n1051 B.n1050 585
R1368 B.n1051 B.n8 585
R1369 B.n1049 B.n7 585
R1370 B.n1232 B.n7 585
R1371 B.n1048 B.n6 585
R1372 B.n1233 B.n6 585
R1373 B.n1047 B.n5 585
R1374 B.n1234 B.n5 585
R1375 B.n1046 B.n1045 585
R1376 B.n1045 B.n4 585
R1377 B.n1044 B.n436 585
R1378 B.n1044 B.n1043 585
R1379 B.n1034 B.n437 585
R1380 B.n438 B.n437 585
R1381 B.n1036 B.n1035 585
R1382 B.n1037 B.n1036 585
R1383 B.n1033 B.n443 585
R1384 B.n443 B.n442 585
R1385 B.n1032 B.n1031 585
R1386 B.n1031 B.n1030 585
R1387 B.n445 B.n444 585
R1388 B.n446 B.n445 585
R1389 B.n1023 B.n1022 585
R1390 B.n1024 B.n1023 585
R1391 B.n1021 B.n451 585
R1392 B.n451 B.n450 585
R1393 B.n1020 B.n1019 585
R1394 B.n1019 B.n1018 585
R1395 B.n453 B.n452 585
R1396 B.n454 B.n453 585
R1397 B.n1011 B.n1010 585
R1398 B.n1012 B.n1011 585
R1399 B.n1009 B.n459 585
R1400 B.n459 B.n458 585
R1401 B.n1008 B.n1007 585
R1402 B.n1007 B.n1006 585
R1403 B.n461 B.n460 585
R1404 B.n462 B.n461 585
R1405 B.n999 B.n998 585
R1406 B.n1000 B.n999 585
R1407 B.n997 B.n467 585
R1408 B.n467 B.n466 585
R1409 B.n996 B.n995 585
R1410 B.n995 B.n994 585
R1411 B.n469 B.n468 585
R1412 B.n470 B.n469 585
R1413 B.n987 B.n986 585
R1414 B.n988 B.n987 585
R1415 B.n985 B.n474 585
R1416 B.n478 B.n474 585
R1417 B.n984 B.n983 585
R1418 B.n983 B.n982 585
R1419 B.n476 B.n475 585
R1420 B.n477 B.n476 585
R1421 B.n975 B.n974 585
R1422 B.n976 B.n975 585
R1423 B.n973 B.n483 585
R1424 B.n483 B.n482 585
R1425 B.n972 B.n971 585
R1426 B.n971 B.n970 585
R1427 B.n485 B.n484 585
R1428 B.n486 B.n485 585
R1429 B.n963 B.n962 585
R1430 B.n964 B.n963 585
R1431 B.n961 B.n490 585
R1432 B.n494 B.n490 585
R1433 B.n960 B.n959 585
R1434 B.n959 B.n958 585
R1435 B.n492 B.n491 585
R1436 B.n493 B.n492 585
R1437 B.n951 B.n950 585
R1438 B.n952 B.n951 585
R1439 B.n949 B.n499 585
R1440 B.n499 B.n498 585
R1441 B.n948 B.n947 585
R1442 B.n947 B.n946 585
R1443 B.n501 B.n500 585
R1444 B.n502 B.n501 585
R1445 B.n939 B.n938 585
R1446 B.n940 B.n939 585
R1447 B.n937 B.n506 585
R1448 B.n510 B.n506 585
R1449 B.n936 B.n935 585
R1450 B.n935 B.n934 585
R1451 B.n508 B.n507 585
R1452 B.n509 B.n508 585
R1453 B.n927 B.n926 585
R1454 B.n928 B.n927 585
R1455 B.n925 B.n515 585
R1456 B.n515 B.n514 585
R1457 B.n924 B.n923 585
R1458 B.n923 B.n922 585
R1459 B.n517 B.n516 585
R1460 B.n518 B.n517 585
R1461 B.n915 B.n914 585
R1462 B.n916 B.n915 585
R1463 B.n913 B.n523 585
R1464 B.n523 B.n522 585
R1465 B.n912 B.n911 585
R1466 B.n911 B.n910 585
R1467 B.n525 B.n524 585
R1468 B.n526 B.n525 585
R1469 B.n903 B.n902 585
R1470 B.n904 B.n903 585
R1471 B.n901 B.n531 585
R1472 B.n531 B.n530 585
R1473 B.n900 B.n899 585
R1474 B.n899 B.n898 585
R1475 B.n533 B.n532 585
R1476 B.n534 B.n533 585
R1477 B.n891 B.n890 585
R1478 B.n892 B.n891 585
R1479 B.n889 B.n539 585
R1480 B.n539 B.n538 585
R1481 B.n888 B.n887 585
R1482 B.n887 B.n886 585
R1483 B.n541 B.n540 585
R1484 B.n542 B.n541 585
R1485 B.n882 B.n881 585
R1486 B.n545 B.n544 585
R1487 B.n878 B.n877 585
R1488 B.n879 B.n878 585
R1489 B.n876 B.n611 585
R1490 B.n875 B.n874 585
R1491 B.n873 B.n872 585
R1492 B.n871 B.n870 585
R1493 B.n869 B.n868 585
R1494 B.n867 B.n866 585
R1495 B.n865 B.n864 585
R1496 B.n863 B.n862 585
R1497 B.n861 B.n860 585
R1498 B.n859 B.n858 585
R1499 B.n857 B.n856 585
R1500 B.n855 B.n854 585
R1501 B.n853 B.n852 585
R1502 B.n851 B.n850 585
R1503 B.n849 B.n848 585
R1504 B.n847 B.n846 585
R1505 B.n845 B.n844 585
R1506 B.n843 B.n842 585
R1507 B.n841 B.n840 585
R1508 B.n839 B.n838 585
R1509 B.n837 B.n836 585
R1510 B.n835 B.n834 585
R1511 B.n833 B.n832 585
R1512 B.n831 B.n830 585
R1513 B.n829 B.n828 585
R1514 B.n827 B.n826 585
R1515 B.n825 B.n824 585
R1516 B.n823 B.n822 585
R1517 B.n821 B.n820 585
R1518 B.n819 B.n818 585
R1519 B.n817 B.n816 585
R1520 B.n815 B.n814 585
R1521 B.n813 B.n812 585
R1522 B.n811 B.n810 585
R1523 B.n809 B.n808 585
R1524 B.n807 B.n806 585
R1525 B.n805 B.n804 585
R1526 B.n803 B.n802 585
R1527 B.n801 B.n800 585
R1528 B.n799 B.n798 585
R1529 B.n797 B.n796 585
R1530 B.n795 B.n794 585
R1531 B.n793 B.n792 585
R1532 B.n791 B.n790 585
R1533 B.n789 B.n788 585
R1534 B.n787 B.n786 585
R1535 B.n785 B.n784 585
R1536 B.n783 B.n782 585
R1537 B.n781 B.n780 585
R1538 B.n779 B.n778 585
R1539 B.n777 B.n776 585
R1540 B.n775 B.n774 585
R1541 B.n773 B.n772 585
R1542 B.n771 B.n770 585
R1543 B.n769 B.n768 585
R1544 B.n767 B.n766 585
R1545 B.n765 B.n764 585
R1546 B.n763 B.n762 585
R1547 B.n761 B.n760 585
R1548 B.n758 B.n757 585
R1549 B.n756 B.n755 585
R1550 B.n754 B.n753 585
R1551 B.n752 B.n751 585
R1552 B.n750 B.n749 585
R1553 B.n748 B.n747 585
R1554 B.n746 B.n745 585
R1555 B.n744 B.n743 585
R1556 B.n742 B.n741 585
R1557 B.n740 B.n739 585
R1558 B.n738 B.n737 585
R1559 B.n736 B.n735 585
R1560 B.n734 B.n733 585
R1561 B.n732 B.n731 585
R1562 B.n730 B.n729 585
R1563 B.n728 B.n727 585
R1564 B.n726 B.n725 585
R1565 B.n724 B.n723 585
R1566 B.n722 B.n721 585
R1567 B.n720 B.n719 585
R1568 B.n718 B.n717 585
R1569 B.n716 B.n715 585
R1570 B.n714 B.n713 585
R1571 B.n712 B.n711 585
R1572 B.n710 B.n709 585
R1573 B.n708 B.n707 585
R1574 B.n706 B.n705 585
R1575 B.n704 B.n703 585
R1576 B.n702 B.n701 585
R1577 B.n700 B.n699 585
R1578 B.n698 B.n697 585
R1579 B.n696 B.n695 585
R1580 B.n694 B.n693 585
R1581 B.n692 B.n691 585
R1582 B.n690 B.n689 585
R1583 B.n688 B.n687 585
R1584 B.n686 B.n685 585
R1585 B.n684 B.n683 585
R1586 B.n682 B.n681 585
R1587 B.n680 B.n679 585
R1588 B.n678 B.n677 585
R1589 B.n676 B.n675 585
R1590 B.n674 B.n673 585
R1591 B.n672 B.n671 585
R1592 B.n670 B.n669 585
R1593 B.n668 B.n667 585
R1594 B.n666 B.n665 585
R1595 B.n664 B.n663 585
R1596 B.n662 B.n661 585
R1597 B.n660 B.n659 585
R1598 B.n658 B.n657 585
R1599 B.n656 B.n655 585
R1600 B.n654 B.n653 585
R1601 B.n652 B.n651 585
R1602 B.n650 B.n649 585
R1603 B.n648 B.n647 585
R1604 B.n646 B.n645 585
R1605 B.n644 B.n643 585
R1606 B.n642 B.n641 585
R1607 B.n640 B.n639 585
R1608 B.n638 B.n637 585
R1609 B.n636 B.n635 585
R1610 B.n634 B.n633 585
R1611 B.n632 B.n631 585
R1612 B.n630 B.n629 585
R1613 B.n628 B.n627 585
R1614 B.n626 B.n625 585
R1615 B.n624 B.n623 585
R1616 B.n622 B.n621 585
R1617 B.n620 B.n619 585
R1618 B.n618 B.n617 585
R1619 B.n883 B.n543 585
R1620 B.n543 B.n542 585
R1621 B.n885 B.n884 585
R1622 B.n886 B.n885 585
R1623 B.n537 B.n536 585
R1624 B.n538 B.n537 585
R1625 B.n894 B.n893 585
R1626 B.n893 B.n892 585
R1627 B.n895 B.n535 585
R1628 B.n535 B.n534 585
R1629 B.n897 B.n896 585
R1630 B.n898 B.n897 585
R1631 B.n529 B.n528 585
R1632 B.n530 B.n529 585
R1633 B.n906 B.n905 585
R1634 B.n905 B.n904 585
R1635 B.n907 B.n527 585
R1636 B.n527 B.n526 585
R1637 B.n909 B.n908 585
R1638 B.n910 B.n909 585
R1639 B.n521 B.n520 585
R1640 B.n522 B.n521 585
R1641 B.n918 B.n917 585
R1642 B.n917 B.n916 585
R1643 B.n919 B.n519 585
R1644 B.n519 B.n518 585
R1645 B.n921 B.n920 585
R1646 B.n922 B.n921 585
R1647 B.n513 B.n512 585
R1648 B.n514 B.n513 585
R1649 B.n930 B.n929 585
R1650 B.n929 B.n928 585
R1651 B.n931 B.n511 585
R1652 B.n511 B.n509 585
R1653 B.n933 B.n932 585
R1654 B.n934 B.n933 585
R1655 B.n505 B.n504 585
R1656 B.n510 B.n505 585
R1657 B.n942 B.n941 585
R1658 B.n941 B.n940 585
R1659 B.n943 B.n503 585
R1660 B.n503 B.n502 585
R1661 B.n945 B.n944 585
R1662 B.n946 B.n945 585
R1663 B.n497 B.n496 585
R1664 B.n498 B.n497 585
R1665 B.n954 B.n953 585
R1666 B.n953 B.n952 585
R1667 B.n955 B.n495 585
R1668 B.n495 B.n493 585
R1669 B.n957 B.n956 585
R1670 B.n958 B.n957 585
R1671 B.n489 B.n488 585
R1672 B.n494 B.n489 585
R1673 B.n966 B.n965 585
R1674 B.n965 B.n964 585
R1675 B.n967 B.n487 585
R1676 B.n487 B.n486 585
R1677 B.n969 B.n968 585
R1678 B.n970 B.n969 585
R1679 B.n481 B.n480 585
R1680 B.n482 B.n481 585
R1681 B.n978 B.n977 585
R1682 B.n977 B.n976 585
R1683 B.n979 B.n479 585
R1684 B.n479 B.n477 585
R1685 B.n981 B.n980 585
R1686 B.n982 B.n981 585
R1687 B.n473 B.n472 585
R1688 B.n478 B.n473 585
R1689 B.n990 B.n989 585
R1690 B.n989 B.n988 585
R1691 B.n991 B.n471 585
R1692 B.n471 B.n470 585
R1693 B.n993 B.n992 585
R1694 B.n994 B.n993 585
R1695 B.n465 B.n464 585
R1696 B.n466 B.n465 585
R1697 B.n1002 B.n1001 585
R1698 B.n1001 B.n1000 585
R1699 B.n1003 B.n463 585
R1700 B.n463 B.n462 585
R1701 B.n1005 B.n1004 585
R1702 B.n1006 B.n1005 585
R1703 B.n457 B.n456 585
R1704 B.n458 B.n457 585
R1705 B.n1014 B.n1013 585
R1706 B.n1013 B.n1012 585
R1707 B.n1015 B.n455 585
R1708 B.n455 B.n454 585
R1709 B.n1017 B.n1016 585
R1710 B.n1018 B.n1017 585
R1711 B.n449 B.n448 585
R1712 B.n450 B.n449 585
R1713 B.n1026 B.n1025 585
R1714 B.n1025 B.n1024 585
R1715 B.n1027 B.n447 585
R1716 B.n447 B.n446 585
R1717 B.n1029 B.n1028 585
R1718 B.n1030 B.n1029 585
R1719 B.n441 B.n440 585
R1720 B.n442 B.n441 585
R1721 B.n1039 B.n1038 585
R1722 B.n1038 B.n1037 585
R1723 B.n1040 B.n439 585
R1724 B.n439 B.n438 585
R1725 B.n1042 B.n1041 585
R1726 B.n1043 B.n1042 585
R1727 B.n3 B.n0 585
R1728 B.n4 B.n3 585
R1729 B.n1231 B.n1 585
R1730 B.n1232 B.n1231 585
R1731 B.n1230 B.n1229 585
R1732 B.n1230 B.n8 585
R1733 B.n1228 B.n9 585
R1734 B.n12 B.n9 585
R1735 B.n1227 B.n1226 585
R1736 B.n1226 B.n1225 585
R1737 B.n11 B.n10 585
R1738 B.n1224 B.n11 585
R1739 B.n1222 B.n1221 585
R1740 B.n1223 B.n1222 585
R1741 B.n1220 B.n17 585
R1742 B.n17 B.n16 585
R1743 B.n1219 B.n1218 585
R1744 B.n1218 B.n1217 585
R1745 B.n19 B.n18 585
R1746 B.n1216 B.n19 585
R1747 B.n1214 B.n1213 585
R1748 B.n1215 B.n1214 585
R1749 B.n1212 B.n24 585
R1750 B.n24 B.n23 585
R1751 B.n1211 B.n1210 585
R1752 B.n1210 B.n1209 585
R1753 B.n26 B.n25 585
R1754 B.n1208 B.n26 585
R1755 B.n1206 B.n1205 585
R1756 B.n1207 B.n1206 585
R1757 B.n1204 B.n31 585
R1758 B.n31 B.n30 585
R1759 B.n1203 B.n1202 585
R1760 B.n1202 B.n1201 585
R1761 B.n33 B.n32 585
R1762 B.n1200 B.n33 585
R1763 B.n1198 B.n1197 585
R1764 B.n1199 B.n1198 585
R1765 B.n1196 B.n38 585
R1766 B.n38 B.n37 585
R1767 B.n1195 B.n1194 585
R1768 B.n1194 B.n1193 585
R1769 B.n40 B.n39 585
R1770 B.n1192 B.n40 585
R1771 B.n1190 B.n1189 585
R1772 B.n1191 B.n1190 585
R1773 B.n1188 B.n45 585
R1774 B.n45 B.n44 585
R1775 B.n1187 B.n1186 585
R1776 B.n1186 B.n1185 585
R1777 B.n47 B.n46 585
R1778 B.n1184 B.n47 585
R1779 B.n1182 B.n1181 585
R1780 B.n1183 B.n1182 585
R1781 B.n1180 B.n52 585
R1782 B.n52 B.n51 585
R1783 B.n1179 B.n1178 585
R1784 B.n1178 B.n1177 585
R1785 B.n54 B.n53 585
R1786 B.n1176 B.n54 585
R1787 B.n1174 B.n1173 585
R1788 B.n1175 B.n1174 585
R1789 B.n1172 B.n59 585
R1790 B.n59 B.n58 585
R1791 B.n1171 B.n1170 585
R1792 B.n1170 B.n1169 585
R1793 B.n61 B.n60 585
R1794 B.n1168 B.n61 585
R1795 B.n1166 B.n1165 585
R1796 B.n1167 B.n1166 585
R1797 B.n1164 B.n66 585
R1798 B.n66 B.n65 585
R1799 B.n1163 B.n1162 585
R1800 B.n1162 B.n1161 585
R1801 B.n68 B.n67 585
R1802 B.n1160 B.n68 585
R1803 B.n1158 B.n1157 585
R1804 B.n1159 B.n1158 585
R1805 B.n1156 B.n73 585
R1806 B.n73 B.n72 585
R1807 B.n1155 B.n1154 585
R1808 B.n1154 B.n1153 585
R1809 B.n75 B.n74 585
R1810 B.n1152 B.n75 585
R1811 B.n1150 B.n1149 585
R1812 B.n1151 B.n1150 585
R1813 B.n1148 B.n80 585
R1814 B.n80 B.n79 585
R1815 B.n1147 B.n1146 585
R1816 B.n1146 B.n1145 585
R1817 B.n82 B.n81 585
R1818 B.n1144 B.n82 585
R1819 B.n1142 B.n1141 585
R1820 B.n1143 B.n1142 585
R1821 B.n1140 B.n87 585
R1822 B.n87 B.n86 585
R1823 B.n1139 B.n1138 585
R1824 B.n1138 B.n1137 585
R1825 B.n89 B.n88 585
R1826 B.n1136 B.n89 585
R1827 B.n1134 B.n1133 585
R1828 B.n1135 B.n1134 585
R1829 B.n1132 B.n94 585
R1830 B.n94 B.n93 585
R1831 B.n1131 B.n1130 585
R1832 B.n1130 B.n1129 585
R1833 B.n96 B.n95 585
R1834 B.n1128 B.n96 585
R1835 B.n1126 B.n1125 585
R1836 B.n1127 B.n1126 585
R1837 B.n1124 B.n101 585
R1838 B.n101 B.n100 585
R1839 B.n1235 B.n1234 585
R1840 B.n1233 B.n2 585
R1841 B.n1122 B.n101 550.159
R1842 B.n1119 B.n170 550.159
R1843 B.n617 B.n541 550.159
R1844 B.n881 B.n543 550.159
R1845 B.n171 B.t22 452.466
R1846 B.n614 B.t16 452.466
R1847 B.n173 B.t19 452.466
R1848 B.n612 B.t13 452.466
R1849 B.n172 B.t23 400.101
R1850 B.n615 B.t15 400.101
R1851 B.n174 B.t20 400.101
R1852 B.n613 B.t12 400.101
R1853 B.n173 B.t17 399.353
R1854 B.n171 B.t21 399.353
R1855 B.n614 B.t14 399.353
R1856 B.n612 B.t10 399.353
R1857 B.n1120 B.n168 256.663
R1858 B.n1120 B.n167 256.663
R1859 B.n1120 B.n166 256.663
R1860 B.n1120 B.n165 256.663
R1861 B.n1120 B.n164 256.663
R1862 B.n1120 B.n163 256.663
R1863 B.n1120 B.n162 256.663
R1864 B.n1120 B.n161 256.663
R1865 B.n1120 B.n160 256.663
R1866 B.n1120 B.n159 256.663
R1867 B.n1120 B.n158 256.663
R1868 B.n1120 B.n157 256.663
R1869 B.n1120 B.n156 256.663
R1870 B.n1120 B.n155 256.663
R1871 B.n1120 B.n154 256.663
R1872 B.n1120 B.n153 256.663
R1873 B.n1120 B.n152 256.663
R1874 B.n1120 B.n151 256.663
R1875 B.n1120 B.n150 256.663
R1876 B.n1120 B.n149 256.663
R1877 B.n1120 B.n148 256.663
R1878 B.n1120 B.n147 256.663
R1879 B.n1120 B.n146 256.663
R1880 B.n1120 B.n145 256.663
R1881 B.n1120 B.n144 256.663
R1882 B.n1120 B.n143 256.663
R1883 B.n1120 B.n142 256.663
R1884 B.n1120 B.n141 256.663
R1885 B.n1120 B.n140 256.663
R1886 B.n1120 B.n139 256.663
R1887 B.n1120 B.n138 256.663
R1888 B.n1120 B.n137 256.663
R1889 B.n1120 B.n136 256.663
R1890 B.n1120 B.n135 256.663
R1891 B.n1120 B.n134 256.663
R1892 B.n1120 B.n133 256.663
R1893 B.n1120 B.n132 256.663
R1894 B.n1120 B.n131 256.663
R1895 B.n1120 B.n130 256.663
R1896 B.n1120 B.n129 256.663
R1897 B.n1120 B.n128 256.663
R1898 B.n1120 B.n127 256.663
R1899 B.n1120 B.n126 256.663
R1900 B.n1120 B.n125 256.663
R1901 B.n1120 B.n124 256.663
R1902 B.n1120 B.n123 256.663
R1903 B.n1120 B.n122 256.663
R1904 B.n1120 B.n121 256.663
R1905 B.n1120 B.n120 256.663
R1906 B.n1120 B.n119 256.663
R1907 B.n1120 B.n118 256.663
R1908 B.n1120 B.n117 256.663
R1909 B.n1120 B.n116 256.663
R1910 B.n1120 B.n115 256.663
R1911 B.n1120 B.n114 256.663
R1912 B.n1120 B.n113 256.663
R1913 B.n1120 B.n112 256.663
R1914 B.n1120 B.n111 256.663
R1915 B.n1120 B.n110 256.663
R1916 B.n1120 B.n109 256.663
R1917 B.n1120 B.n108 256.663
R1918 B.n1120 B.n107 256.663
R1919 B.n1120 B.n106 256.663
R1920 B.n1120 B.n105 256.663
R1921 B.n1120 B.n104 256.663
R1922 B.n1121 B.n1120 256.663
R1923 B.n880 B.n879 256.663
R1924 B.n879 B.n546 256.663
R1925 B.n879 B.n547 256.663
R1926 B.n879 B.n548 256.663
R1927 B.n879 B.n549 256.663
R1928 B.n879 B.n550 256.663
R1929 B.n879 B.n551 256.663
R1930 B.n879 B.n552 256.663
R1931 B.n879 B.n553 256.663
R1932 B.n879 B.n554 256.663
R1933 B.n879 B.n555 256.663
R1934 B.n879 B.n556 256.663
R1935 B.n879 B.n557 256.663
R1936 B.n879 B.n558 256.663
R1937 B.n879 B.n559 256.663
R1938 B.n879 B.n560 256.663
R1939 B.n879 B.n561 256.663
R1940 B.n879 B.n562 256.663
R1941 B.n879 B.n563 256.663
R1942 B.n879 B.n564 256.663
R1943 B.n879 B.n565 256.663
R1944 B.n879 B.n566 256.663
R1945 B.n879 B.n567 256.663
R1946 B.n879 B.n568 256.663
R1947 B.n879 B.n569 256.663
R1948 B.n879 B.n570 256.663
R1949 B.n879 B.n571 256.663
R1950 B.n879 B.n572 256.663
R1951 B.n879 B.n573 256.663
R1952 B.n879 B.n574 256.663
R1953 B.n879 B.n575 256.663
R1954 B.n879 B.n576 256.663
R1955 B.n879 B.n577 256.663
R1956 B.n879 B.n578 256.663
R1957 B.n879 B.n579 256.663
R1958 B.n879 B.n580 256.663
R1959 B.n879 B.n581 256.663
R1960 B.n879 B.n582 256.663
R1961 B.n879 B.n583 256.663
R1962 B.n879 B.n584 256.663
R1963 B.n879 B.n585 256.663
R1964 B.n879 B.n586 256.663
R1965 B.n879 B.n587 256.663
R1966 B.n879 B.n588 256.663
R1967 B.n879 B.n589 256.663
R1968 B.n879 B.n590 256.663
R1969 B.n879 B.n591 256.663
R1970 B.n879 B.n592 256.663
R1971 B.n879 B.n593 256.663
R1972 B.n879 B.n594 256.663
R1973 B.n879 B.n595 256.663
R1974 B.n879 B.n596 256.663
R1975 B.n879 B.n597 256.663
R1976 B.n879 B.n598 256.663
R1977 B.n879 B.n599 256.663
R1978 B.n879 B.n600 256.663
R1979 B.n879 B.n601 256.663
R1980 B.n879 B.n602 256.663
R1981 B.n879 B.n603 256.663
R1982 B.n879 B.n604 256.663
R1983 B.n879 B.n605 256.663
R1984 B.n879 B.n606 256.663
R1985 B.n879 B.n607 256.663
R1986 B.n879 B.n608 256.663
R1987 B.n879 B.n609 256.663
R1988 B.n879 B.n610 256.663
R1989 B.n1237 B.n1236 256.663
R1990 B.n176 B.n103 163.367
R1991 B.n180 B.n179 163.367
R1992 B.n184 B.n183 163.367
R1993 B.n188 B.n187 163.367
R1994 B.n192 B.n191 163.367
R1995 B.n196 B.n195 163.367
R1996 B.n200 B.n199 163.367
R1997 B.n204 B.n203 163.367
R1998 B.n208 B.n207 163.367
R1999 B.n212 B.n211 163.367
R2000 B.n216 B.n215 163.367
R2001 B.n220 B.n219 163.367
R2002 B.n224 B.n223 163.367
R2003 B.n228 B.n227 163.367
R2004 B.n232 B.n231 163.367
R2005 B.n236 B.n235 163.367
R2006 B.n240 B.n239 163.367
R2007 B.n244 B.n243 163.367
R2008 B.n248 B.n247 163.367
R2009 B.n252 B.n251 163.367
R2010 B.n256 B.n255 163.367
R2011 B.n260 B.n259 163.367
R2012 B.n264 B.n263 163.367
R2013 B.n268 B.n267 163.367
R2014 B.n272 B.n271 163.367
R2015 B.n276 B.n275 163.367
R2016 B.n280 B.n279 163.367
R2017 B.n284 B.n283 163.367
R2018 B.n288 B.n287 163.367
R2019 B.n292 B.n291 163.367
R2020 B.n296 B.n295 163.367
R2021 B.n300 B.n299 163.367
R2022 B.n304 B.n303 163.367
R2023 B.n308 B.n307 163.367
R2024 B.n312 B.n311 163.367
R2025 B.n317 B.n316 163.367
R2026 B.n321 B.n320 163.367
R2027 B.n325 B.n324 163.367
R2028 B.n329 B.n328 163.367
R2029 B.n333 B.n332 163.367
R2030 B.n337 B.n336 163.367
R2031 B.n341 B.n340 163.367
R2032 B.n345 B.n344 163.367
R2033 B.n349 B.n348 163.367
R2034 B.n353 B.n352 163.367
R2035 B.n357 B.n356 163.367
R2036 B.n361 B.n360 163.367
R2037 B.n365 B.n364 163.367
R2038 B.n369 B.n368 163.367
R2039 B.n373 B.n372 163.367
R2040 B.n377 B.n376 163.367
R2041 B.n381 B.n380 163.367
R2042 B.n385 B.n384 163.367
R2043 B.n389 B.n388 163.367
R2044 B.n393 B.n392 163.367
R2045 B.n397 B.n396 163.367
R2046 B.n401 B.n400 163.367
R2047 B.n405 B.n404 163.367
R2048 B.n409 B.n408 163.367
R2049 B.n413 B.n412 163.367
R2050 B.n417 B.n416 163.367
R2051 B.n421 B.n420 163.367
R2052 B.n425 B.n424 163.367
R2053 B.n429 B.n428 163.367
R2054 B.n433 B.n432 163.367
R2055 B.n1119 B.n169 163.367
R2056 B.n887 B.n541 163.367
R2057 B.n887 B.n539 163.367
R2058 B.n891 B.n539 163.367
R2059 B.n891 B.n533 163.367
R2060 B.n899 B.n533 163.367
R2061 B.n899 B.n531 163.367
R2062 B.n903 B.n531 163.367
R2063 B.n903 B.n525 163.367
R2064 B.n911 B.n525 163.367
R2065 B.n911 B.n523 163.367
R2066 B.n915 B.n523 163.367
R2067 B.n915 B.n517 163.367
R2068 B.n923 B.n517 163.367
R2069 B.n923 B.n515 163.367
R2070 B.n927 B.n515 163.367
R2071 B.n927 B.n508 163.367
R2072 B.n935 B.n508 163.367
R2073 B.n935 B.n506 163.367
R2074 B.n939 B.n506 163.367
R2075 B.n939 B.n501 163.367
R2076 B.n947 B.n501 163.367
R2077 B.n947 B.n499 163.367
R2078 B.n951 B.n499 163.367
R2079 B.n951 B.n492 163.367
R2080 B.n959 B.n492 163.367
R2081 B.n959 B.n490 163.367
R2082 B.n963 B.n490 163.367
R2083 B.n963 B.n485 163.367
R2084 B.n971 B.n485 163.367
R2085 B.n971 B.n483 163.367
R2086 B.n975 B.n483 163.367
R2087 B.n975 B.n476 163.367
R2088 B.n983 B.n476 163.367
R2089 B.n983 B.n474 163.367
R2090 B.n987 B.n474 163.367
R2091 B.n987 B.n469 163.367
R2092 B.n995 B.n469 163.367
R2093 B.n995 B.n467 163.367
R2094 B.n999 B.n467 163.367
R2095 B.n999 B.n461 163.367
R2096 B.n1007 B.n461 163.367
R2097 B.n1007 B.n459 163.367
R2098 B.n1011 B.n459 163.367
R2099 B.n1011 B.n453 163.367
R2100 B.n1019 B.n453 163.367
R2101 B.n1019 B.n451 163.367
R2102 B.n1023 B.n451 163.367
R2103 B.n1023 B.n445 163.367
R2104 B.n1031 B.n445 163.367
R2105 B.n1031 B.n443 163.367
R2106 B.n1036 B.n443 163.367
R2107 B.n1036 B.n437 163.367
R2108 B.n1044 B.n437 163.367
R2109 B.n1045 B.n1044 163.367
R2110 B.n1045 B.n5 163.367
R2111 B.n6 B.n5 163.367
R2112 B.n7 B.n6 163.367
R2113 B.n1051 B.n7 163.367
R2114 B.n1052 B.n1051 163.367
R2115 B.n1052 B.n13 163.367
R2116 B.n14 B.n13 163.367
R2117 B.n15 B.n14 163.367
R2118 B.n1057 B.n15 163.367
R2119 B.n1057 B.n20 163.367
R2120 B.n21 B.n20 163.367
R2121 B.n22 B.n21 163.367
R2122 B.n1062 B.n22 163.367
R2123 B.n1062 B.n27 163.367
R2124 B.n28 B.n27 163.367
R2125 B.n29 B.n28 163.367
R2126 B.n1067 B.n29 163.367
R2127 B.n1067 B.n34 163.367
R2128 B.n35 B.n34 163.367
R2129 B.n36 B.n35 163.367
R2130 B.n1072 B.n36 163.367
R2131 B.n1072 B.n41 163.367
R2132 B.n42 B.n41 163.367
R2133 B.n43 B.n42 163.367
R2134 B.n1077 B.n43 163.367
R2135 B.n1077 B.n48 163.367
R2136 B.n49 B.n48 163.367
R2137 B.n50 B.n49 163.367
R2138 B.n1082 B.n50 163.367
R2139 B.n1082 B.n55 163.367
R2140 B.n56 B.n55 163.367
R2141 B.n57 B.n56 163.367
R2142 B.n1087 B.n57 163.367
R2143 B.n1087 B.n62 163.367
R2144 B.n63 B.n62 163.367
R2145 B.n64 B.n63 163.367
R2146 B.n1092 B.n64 163.367
R2147 B.n1092 B.n69 163.367
R2148 B.n70 B.n69 163.367
R2149 B.n71 B.n70 163.367
R2150 B.n1097 B.n71 163.367
R2151 B.n1097 B.n76 163.367
R2152 B.n77 B.n76 163.367
R2153 B.n78 B.n77 163.367
R2154 B.n1102 B.n78 163.367
R2155 B.n1102 B.n83 163.367
R2156 B.n84 B.n83 163.367
R2157 B.n85 B.n84 163.367
R2158 B.n1107 B.n85 163.367
R2159 B.n1107 B.n90 163.367
R2160 B.n91 B.n90 163.367
R2161 B.n92 B.n91 163.367
R2162 B.n1112 B.n92 163.367
R2163 B.n1112 B.n97 163.367
R2164 B.n98 B.n97 163.367
R2165 B.n99 B.n98 163.367
R2166 B.n170 B.n99 163.367
R2167 B.n878 B.n545 163.367
R2168 B.n878 B.n611 163.367
R2169 B.n874 B.n873 163.367
R2170 B.n870 B.n869 163.367
R2171 B.n866 B.n865 163.367
R2172 B.n862 B.n861 163.367
R2173 B.n858 B.n857 163.367
R2174 B.n854 B.n853 163.367
R2175 B.n850 B.n849 163.367
R2176 B.n846 B.n845 163.367
R2177 B.n842 B.n841 163.367
R2178 B.n838 B.n837 163.367
R2179 B.n834 B.n833 163.367
R2180 B.n830 B.n829 163.367
R2181 B.n826 B.n825 163.367
R2182 B.n822 B.n821 163.367
R2183 B.n818 B.n817 163.367
R2184 B.n814 B.n813 163.367
R2185 B.n810 B.n809 163.367
R2186 B.n806 B.n805 163.367
R2187 B.n802 B.n801 163.367
R2188 B.n798 B.n797 163.367
R2189 B.n794 B.n793 163.367
R2190 B.n790 B.n789 163.367
R2191 B.n786 B.n785 163.367
R2192 B.n782 B.n781 163.367
R2193 B.n778 B.n777 163.367
R2194 B.n774 B.n773 163.367
R2195 B.n770 B.n769 163.367
R2196 B.n766 B.n765 163.367
R2197 B.n762 B.n761 163.367
R2198 B.n757 B.n756 163.367
R2199 B.n753 B.n752 163.367
R2200 B.n749 B.n748 163.367
R2201 B.n745 B.n744 163.367
R2202 B.n741 B.n740 163.367
R2203 B.n737 B.n736 163.367
R2204 B.n733 B.n732 163.367
R2205 B.n729 B.n728 163.367
R2206 B.n725 B.n724 163.367
R2207 B.n721 B.n720 163.367
R2208 B.n717 B.n716 163.367
R2209 B.n713 B.n712 163.367
R2210 B.n709 B.n708 163.367
R2211 B.n705 B.n704 163.367
R2212 B.n701 B.n700 163.367
R2213 B.n697 B.n696 163.367
R2214 B.n693 B.n692 163.367
R2215 B.n689 B.n688 163.367
R2216 B.n685 B.n684 163.367
R2217 B.n681 B.n680 163.367
R2218 B.n677 B.n676 163.367
R2219 B.n673 B.n672 163.367
R2220 B.n669 B.n668 163.367
R2221 B.n665 B.n664 163.367
R2222 B.n661 B.n660 163.367
R2223 B.n657 B.n656 163.367
R2224 B.n653 B.n652 163.367
R2225 B.n649 B.n648 163.367
R2226 B.n645 B.n644 163.367
R2227 B.n641 B.n640 163.367
R2228 B.n637 B.n636 163.367
R2229 B.n633 B.n632 163.367
R2230 B.n629 B.n628 163.367
R2231 B.n625 B.n624 163.367
R2232 B.n621 B.n620 163.367
R2233 B.n885 B.n543 163.367
R2234 B.n885 B.n537 163.367
R2235 B.n893 B.n537 163.367
R2236 B.n893 B.n535 163.367
R2237 B.n897 B.n535 163.367
R2238 B.n897 B.n529 163.367
R2239 B.n905 B.n529 163.367
R2240 B.n905 B.n527 163.367
R2241 B.n909 B.n527 163.367
R2242 B.n909 B.n521 163.367
R2243 B.n917 B.n521 163.367
R2244 B.n917 B.n519 163.367
R2245 B.n921 B.n519 163.367
R2246 B.n921 B.n513 163.367
R2247 B.n929 B.n513 163.367
R2248 B.n929 B.n511 163.367
R2249 B.n933 B.n511 163.367
R2250 B.n933 B.n505 163.367
R2251 B.n941 B.n505 163.367
R2252 B.n941 B.n503 163.367
R2253 B.n945 B.n503 163.367
R2254 B.n945 B.n497 163.367
R2255 B.n953 B.n497 163.367
R2256 B.n953 B.n495 163.367
R2257 B.n957 B.n495 163.367
R2258 B.n957 B.n489 163.367
R2259 B.n965 B.n489 163.367
R2260 B.n965 B.n487 163.367
R2261 B.n969 B.n487 163.367
R2262 B.n969 B.n481 163.367
R2263 B.n977 B.n481 163.367
R2264 B.n977 B.n479 163.367
R2265 B.n981 B.n479 163.367
R2266 B.n981 B.n473 163.367
R2267 B.n989 B.n473 163.367
R2268 B.n989 B.n471 163.367
R2269 B.n993 B.n471 163.367
R2270 B.n993 B.n465 163.367
R2271 B.n1001 B.n465 163.367
R2272 B.n1001 B.n463 163.367
R2273 B.n1005 B.n463 163.367
R2274 B.n1005 B.n457 163.367
R2275 B.n1013 B.n457 163.367
R2276 B.n1013 B.n455 163.367
R2277 B.n1017 B.n455 163.367
R2278 B.n1017 B.n449 163.367
R2279 B.n1025 B.n449 163.367
R2280 B.n1025 B.n447 163.367
R2281 B.n1029 B.n447 163.367
R2282 B.n1029 B.n441 163.367
R2283 B.n1038 B.n441 163.367
R2284 B.n1038 B.n439 163.367
R2285 B.n1042 B.n439 163.367
R2286 B.n1042 B.n3 163.367
R2287 B.n1235 B.n3 163.367
R2288 B.n1231 B.n2 163.367
R2289 B.n1231 B.n1230 163.367
R2290 B.n1230 B.n9 163.367
R2291 B.n1226 B.n9 163.367
R2292 B.n1226 B.n11 163.367
R2293 B.n1222 B.n11 163.367
R2294 B.n1222 B.n17 163.367
R2295 B.n1218 B.n17 163.367
R2296 B.n1218 B.n19 163.367
R2297 B.n1214 B.n19 163.367
R2298 B.n1214 B.n24 163.367
R2299 B.n1210 B.n24 163.367
R2300 B.n1210 B.n26 163.367
R2301 B.n1206 B.n26 163.367
R2302 B.n1206 B.n31 163.367
R2303 B.n1202 B.n31 163.367
R2304 B.n1202 B.n33 163.367
R2305 B.n1198 B.n33 163.367
R2306 B.n1198 B.n38 163.367
R2307 B.n1194 B.n38 163.367
R2308 B.n1194 B.n40 163.367
R2309 B.n1190 B.n40 163.367
R2310 B.n1190 B.n45 163.367
R2311 B.n1186 B.n45 163.367
R2312 B.n1186 B.n47 163.367
R2313 B.n1182 B.n47 163.367
R2314 B.n1182 B.n52 163.367
R2315 B.n1178 B.n52 163.367
R2316 B.n1178 B.n54 163.367
R2317 B.n1174 B.n54 163.367
R2318 B.n1174 B.n59 163.367
R2319 B.n1170 B.n59 163.367
R2320 B.n1170 B.n61 163.367
R2321 B.n1166 B.n61 163.367
R2322 B.n1166 B.n66 163.367
R2323 B.n1162 B.n66 163.367
R2324 B.n1162 B.n68 163.367
R2325 B.n1158 B.n68 163.367
R2326 B.n1158 B.n73 163.367
R2327 B.n1154 B.n73 163.367
R2328 B.n1154 B.n75 163.367
R2329 B.n1150 B.n75 163.367
R2330 B.n1150 B.n80 163.367
R2331 B.n1146 B.n80 163.367
R2332 B.n1146 B.n82 163.367
R2333 B.n1142 B.n82 163.367
R2334 B.n1142 B.n87 163.367
R2335 B.n1138 B.n87 163.367
R2336 B.n1138 B.n89 163.367
R2337 B.n1134 B.n89 163.367
R2338 B.n1134 B.n94 163.367
R2339 B.n1130 B.n94 163.367
R2340 B.n1130 B.n96 163.367
R2341 B.n1126 B.n96 163.367
R2342 B.n1126 B.n101 163.367
R2343 B.n1122 B.n1121 71.676
R2344 B.n176 B.n104 71.676
R2345 B.n180 B.n105 71.676
R2346 B.n184 B.n106 71.676
R2347 B.n188 B.n107 71.676
R2348 B.n192 B.n108 71.676
R2349 B.n196 B.n109 71.676
R2350 B.n200 B.n110 71.676
R2351 B.n204 B.n111 71.676
R2352 B.n208 B.n112 71.676
R2353 B.n212 B.n113 71.676
R2354 B.n216 B.n114 71.676
R2355 B.n220 B.n115 71.676
R2356 B.n224 B.n116 71.676
R2357 B.n228 B.n117 71.676
R2358 B.n232 B.n118 71.676
R2359 B.n236 B.n119 71.676
R2360 B.n240 B.n120 71.676
R2361 B.n244 B.n121 71.676
R2362 B.n248 B.n122 71.676
R2363 B.n252 B.n123 71.676
R2364 B.n256 B.n124 71.676
R2365 B.n260 B.n125 71.676
R2366 B.n264 B.n126 71.676
R2367 B.n268 B.n127 71.676
R2368 B.n272 B.n128 71.676
R2369 B.n276 B.n129 71.676
R2370 B.n280 B.n130 71.676
R2371 B.n284 B.n131 71.676
R2372 B.n288 B.n132 71.676
R2373 B.n292 B.n133 71.676
R2374 B.n296 B.n134 71.676
R2375 B.n300 B.n135 71.676
R2376 B.n304 B.n136 71.676
R2377 B.n308 B.n137 71.676
R2378 B.n312 B.n138 71.676
R2379 B.n317 B.n139 71.676
R2380 B.n321 B.n140 71.676
R2381 B.n325 B.n141 71.676
R2382 B.n329 B.n142 71.676
R2383 B.n333 B.n143 71.676
R2384 B.n337 B.n144 71.676
R2385 B.n341 B.n145 71.676
R2386 B.n345 B.n146 71.676
R2387 B.n349 B.n147 71.676
R2388 B.n353 B.n148 71.676
R2389 B.n357 B.n149 71.676
R2390 B.n361 B.n150 71.676
R2391 B.n365 B.n151 71.676
R2392 B.n369 B.n152 71.676
R2393 B.n373 B.n153 71.676
R2394 B.n377 B.n154 71.676
R2395 B.n381 B.n155 71.676
R2396 B.n385 B.n156 71.676
R2397 B.n389 B.n157 71.676
R2398 B.n393 B.n158 71.676
R2399 B.n397 B.n159 71.676
R2400 B.n401 B.n160 71.676
R2401 B.n405 B.n161 71.676
R2402 B.n409 B.n162 71.676
R2403 B.n413 B.n163 71.676
R2404 B.n417 B.n164 71.676
R2405 B.n421 B.n165 71.676
R2406 B.n425 B.n166 71.676
R2407 B.n429 B.n167 71.676
R2408 B.n433 B.n168 71.676
R2409 B.n169 B.n168 71.676
R2410 B.n432 B.n167 71.676
R2411 B.n428 B.n166 71.676
R2412 B.n424 B.n165 71.676
R2413 B.n420 B.n164 71.676
R2414 B.n416 B.n163 71.676
R2415 B.n412 B.n162 71.676
R2416 B.n408 B.n161 71.676
R2417 B.n404 B.n160 71.676
R2418 B.n400 B.n159 71.676
R2419 B.n396 B.n158 71.676
R2420 B.n392 B.n157 71.676
R2421 B.n388 B.n156 71.676
R2422 B.n384 B.n155 71.676
R2423 B.n380 B.n154 71.676
R2424 B.n376 B.n153 71.676
R2425 B.n372 B.n152 71.676
R2426 B.n368 B.n151 71.676
R2427 B.n364 B.n150 71.676
R2428 B.n360 B.n149 71.676
R2429 B.n356 B.n148 71.676
R2430 B.n352 B.n147 71.676
R2431 B.n348 B.n146 71.676
R2432 B.n344 B.n145 71.676
R2433 B.n340 B.n144 71.676
R2434 B.n336 B.n143 71.676
R2435 B.n332 B.n142 71.676
R2436 B.n328 B.n141 71.676
R2437 B.n324 B.n140 71.676
R2438 B.n320 B.n139 71.676
R2439 B.n316 B.n138 71.676
R2440 B.n311 B.n137 71.676
R2441 B.n307 B.n136 71.676
R2442 B.n303 B.n135 71.676
R2443 B.n299 B.n134 71.676
R2444 B.n295 B.n133 71.676
R2445 B.n291 B.n132 71.676
R2446 B.n287 B.n131 71.676
R2447 B.n283 B.n130 71.676
R2448 B.n279 B.n129 71.676
R2449 B.n275 B.n128 71.676
R2450 B.n271 B.n127 71.676
R2451 B.n267 B.n126 71.676
R2452 B.n263 B.n125 71.676
R2453 B.n259 B.n124 71.676
R2454 B.n255 B.n123 71.676
R2455 B.n251 B.n122 71.676
R2456 B.n247 B.n121 71.676
R2457 B.n243 B.n120 71.676
R2458 B.n239 B.n119 71.676
R2459 B.n235 B.n118 71.676
R2460 B.n231 B.n117 71.676
R2461 B.n227 B.n116 71.676
R2462 B.n223 B.n115 71.676
R2463 B.n219 B.n114 71.676
R2464 B.n215 B.n113 71.676
R2465 B.n211 B.n112 71.676
R2466 B.n207 B.n111 71.676
R2467 B.n203 B.n110 71.676
R2468 B.n199 B.n109 71.676
R2469 B.n195 B.n108 71.676
R2470 B.n191 B.n107 71.676
R2471 B.n187 B.n106 71.676
R2472 B.n183 B.n105 71.676
R2473 B.n179 B.n104 71.676
R2474 B.n1121 B.n103 71.676
R2475 B.n881 B.n880 71.676
R2476 B.n611 B.n546 71.676
R2477 B.n873 B.n547 71.676
R2478 B.n869 B.n548 71.676
R2479 B.n865 B.n549 71.676
R2480 B.n861 B.n550 71.676
R2481 B.n857 B.n551 71.676
R2482 B.n853 B.n552 71.676
R2483 B.n849 B.n553 71.676
R2484 B.n845 B.n554 71.676
R2485 B.n841 B.n555 71.676
R2486 B.n837 B.n556 71.676
R2487 B.n833 B.n557 71.676
R2488 B.n829 B.n558 71.676
R2489 B.n825 B.n559 71.676
R2490 B.n821 B.n560 71.676
R2491 B.n817 B.n561 71.676
R2492 B.n813 B.n562 71.676
R2493 B.n809 B.n563 71.676
R2494 B.n805 B.n564 71.676
R2495 B.n801 B.n565 71.676
R2496 B.n797 B.n566 71.676
R2497 B.n793 B.n567 71.676
R2498 B.n789 B.n568 71.676
R2499 B.n785 B.n569 71.676
R2500 B.n781 B.n570 71.676
R2501 B.n777 B.n571 71.676
R2502 B.n773 B.n572 71.676
R2503 B.n769 B.n573 71.676
R2504 B.n765 B.n574 71.676
R2505 B.n761 B.n575 71.676
R2506 B.n756 B.n576 71.676
R2507 B.n752 B.n577 71.676
R2508 B.n748 B.n578 71.676
R2509 B.n744 B.n579 71.676
R2510 B.n740 B.n580 71.676
R2511 B.n736 B.n581 71.676
R2512 B.n732 B.n582 71.676
R2513 B.n728 B.n583 71.676
R2514 B.n724 B.n584 71.676
R2515 B.n720 B.n585 71.676
R2516 B.n716 B.n586 71.676
R2517 B.n712 B.n587 71.676
R2518 B.n708 B.n588 71.676
R2519 B.n704 B.n589 71.676
R2520 B.n700 B.n590 71.676
R2521 B.n696 B.n591 71.676
R2522 B.n692 B.n592 71.676
R2523 B.n688 B.n593 71.676
R2524 B.n684 B.n594 71.676
R2525 B.n680 B.n595 71.676
R2526 B.n676 B.n596 71.676
R2527 B.n672 B.n597 71.676
R2528 B.n668 B.n598 71.676
R2529 B.n664 B.n599 71.676
R2530 B.n660 B.n600 71.676
R2531 B.n656 B.n601 71.676
R2532 B.n652 B.n602 71.676
R2533 B.n648 B.n603 71.676
R2534 B.n644 B.n604 71.676
R2535 B.n640 B.n605 71.676
R2536 B.n636 B.n606 71.676
R2537 B.n632 B.n607 71.676
R2538 B.n628 B.n608 71.676
R2539 B.n624 B.n609 71.676
R2540 B.n620 B.n610 71.676
R2541 B.n880 B.n545 71.676
R2542 B.n874 B.n546 71.676
R2543 B.n870 B.n547 71.676
R2544 B.n866 B.n548 71.676
R2545 B.n862 B.n549 71.676
R2546 B.n858 B.n550 71.676
R2547 B.n854 B.n551 71.676
R2548 B.n850 B.n552 71.676
R2549 B.n846 B.n553 71.676
R2550 B.n842 B.n554 71.676
R2551 B.n838 B.n555 71.676
R2552 B.n834 B.n556 71.676
R2553 B.n830 B.n557 71.676
R2554 B.n826 B.n558 71.676
R2555 B.n822 B.n559 71.676
R2556 B.n818 B.n560 71.676
R2557 B.n814 B.n561 71.676
R2558 B.n810 B.n562 71.676
R2559 B.n806 B.n563 71.676
R2560 B.n802 B.n564 71.676
R2561 B.n798 B.n565 71.676
R2562 B.n794 B.n566 71.676
R2563 B.n790 B.n567 71.676
R2564 B.n786 B.n568 71.676
R2565 B.n782 B.n569 71.676
R2566 B.n778 B.n570 71.676
R2567 B.n774 B.n571 71.676
R2568 B.n770 B.n572 71.676
R2569 B.n766 B.n573 71.676
R2570 B.n762 B.n574 71.676
R2571 B.n757 B.n575 71.676
R2572 B.n753 B.n576 71.676
R2573 B.n749 B.n577 71.676
R2574 B.n745 B.n578 71.676
R2575 B.n741 B.n579 71.676
R2576 B.n737 B.n580 71.676
R2577 B.n733 B.n581 71.676
R2578 B.n729 B.n582 71.676
R2579 B.n725 B.n583 71.676
R2580 B.n721 B.n584 71.676
R2581 B.n717 B.n585 71.676
R2582 B.n713 B.n586 71.676
R2583 B.n709 B.n587 71.676
R2584 B.n705 B.n588 71.676
R2585 B.n701 B.n589 71.676
R2586 B.n697 B.n590 71.676
R2587 B.n693 B.n591 71.676
R2588 B.n689 B.n592 71.676
R2589 B.n685 B.n593 71.676
R2590 B.n681 B.n594 71.676
R2591 B.n677 B.n595 71.676
R2592 B.n673 B.n596 71.676
R2593 B.n669 B.n597 71.676
R2594 B.n665 B.n598 71.676
R2595 B.n661 B.n599 71.676
R2596 B.n657 B.n600 71.676
R2597 B.n653 B.n601 71.676
R2598 B.n649 B.n602 71.676
R2599 B.n645 B.n603 71.676
R2600 B.n641 B.n604 71.676
R2601 B.n637 B.n605 71.676
R2602 B.n633 B.n606 71.676
R2603 B.n629 B.n607 71.676
R2604 B.n625 B.n608 71.676
R2605 B.n621 B.n609 71.676
R2606 B.n617 B.n610 71.676
R2607 B.n1236 B.n1235 71.676
R2608 B.n1236 B.n2 71.676
R2609 B.n879 B.n542 64.2907
R2610 B.n1120 B.n100 64.2907
R2611 B.n175 B.n174 59.5399
R2612 B.n314 B.n172 59.5399
R2613 B.n616 B.n615 59.5399
R2614 B.n759 B.n613 59.5399
R2615 B.n174 B.n173 52.3641
R2616 B.n172 B.n171 52.3641
R2617 B.n615 B.n614 52.3641
R2618 B.n613 B.n612 52.3641
R2619 B.n1118 B.n1117 35.7468
R2620 B.n883 B.n882 35.7468
R2621 B.n618 B.n540 35.7468
R2622 B.n1124 B.n1123 35.7468
R2623 B.n886 B.n542 31.0057
R2624 B.n886 B.n538 31.0057
R2625 B.n892 B.n538 31.0057
R2626 B.n892 B.n534 31.0057
R2627 B.n898 B.n534 31.0057
R2628 B.n898 B.n530 31.0057
R2629 B.n904 B.n530 31.0057
R2630 B.n910 B.n526 31.0057
R2631 B.n910 B.n522 31.0057
R2632 B.n916 B.n522 31.0057
R2633 B.n916 B.n518 31.0057
R2634 B.n922 B.n518 31.0057
R2635 B.n922 B.n514 31.0057
R2636 B.n928 B.n514 31.0057
R2637 B.n928 B.n509 31.0057
R2638 B.n934 B.n509 31.0057
R2639 B.n934 B.n510 31.0057
R2640 B.n940 B.n502 31.0057
R2641 B.n946 B.n502 31.0057
R2642 B.n946 B.n498 31.0057
R2643 B.n952 B.n498 31.0057
R2644 B.n952 B.n493 31.0057
R2645 B.n958 B.n493 31.0057
R2646 B.n958 B.n494 31.0057
R2647 B.n964 B.n486 31.0057
R2648 B.n970 B.n486 31.0057
R2649 B.n970 B.n482 31.0057
R2650 B.n976 B.n482 31.0057
R2651 B.n976 B.n477 31.0057
R2652 B.n982 B.n477 31.0057
R2653 B.n982 B.n478 31.0057
R2654 B.n988 B.n470 31.0057
R2655 B.n994 B.n470 31.0057
R2656 B.n994 B.n466 31.0057
R2657 B.n1000 B.n466 31.0057
R2658 B.n1000 B.n462 31.0057
R2659 B.n1006 B.n462 31.0057
R2660 B.n1012 B.n458 31.0057
R2661 B.n1012 B.n454 31.0057
R2662 B.n1018 B.n454 31.0057
R2663 B.n1018 B.n450 31.0057
R2664 B.n1024 B.n450 31.0057
R2665 B.n1024 B.n446 31.0057
R2666 B.n1030 B.n446 31.0057
R2667 B.n1037 B.n442 31.0057
R2668 B.n1037 B.n438 31.0057
R2669 B.n1043 B.n438 31.0057
R2670 B.n1043 B.n4 31.0057
R2671 B.n1234 B.n4 31.0057
R2672 B.n1234 B.n1233 31.0057
R2673 B.n1233 B.n1232 31.0057
R2674 B.n1232 B.n8 31.0057
R2675 B.n12 B.n8 31.0057
R2676 B.n1225 B.n12 31.0057
R2677 B.n1225 B.n1224 31.0057
R2678 B.n1223 B.n16 31.0057
R2679 B.n1217 B.n16 31.0057
R2680 B.n1217 B.n1216 31.0057
R2681 B.n1216 B.n1215 31.0057
R2682 B.n1215 B.n23 31.0057
R2683 B.n1209 B.n23 31.0057
R2684 B.n1209 B.n1208 31.0057
R2685 B.n1207 B.n30 31.0057
R2686 B.n1201 B.n30 31.0057
R2687 B.n1201 B.n1200 31.0057
R2688 B.n1200 B.n1199 31.0057
R2689 B.n1199 B.n37 31.0057
R2690 B.n1193 B.n37 31.0057
R2691 B.n1192 B.n1191 31.0057
R2692 B.n1191 B.n44 31.0057
R2693 B.n1185 B.n44 31.0057
R2694 B.n1185 B.n1184 31.0057
R2695 B.n1184 B.n1183 31.0057
R2696 B.n1183 B.n51 31.0057
R2697 B.n1177 B.n51 31.0057
R2698 B.n1176 B.n1175 31.0057
R2699 B.n1175 B.n58 31.0057
R2700 B.n1169 B.n58 31.0057
R2701 B.n1169 B.n1168 31.0057
R2702 B.n1168 B.n1167 31.0057
R2703 B.n1167 B.n65 31.0057
R2704 B.n1161 B.n65 31.0057
R2705 B.n1160 B.n1159 31.0057
R2706 B.n1159 B.n72 31.0057
R2707 B.n1153 B.n72 31.0057
R2708 B.n1153 B.n1152 31.0057
R2709 B.n1152 B.n1151 31.0057
R2710 B.n1151 B.n79 31.0057
R2711 B.n1145 B.n79 31.0057
R2712 B.n1145 B.n1144 31.0057
R2713 B.n1144 B.n1143 31.0057
R2714 B.n1143 B.n86 31.0057
R2715 B.n1137 B.n1136 31.0057
R2716 B.n1136 B.n1135 31.0057
R2717 B.n1135 B.n93 31.0057
R2718 B.n1129 B.n93 31.0057
R2719 B.n1129 B.n1128 31.0057
R2720 B.n1128 B.n1127 31.0057
R2721 B.n1127 B.n100 31.0057
R2722 B.t11 B.n526 30.5497
R2723 B.n1006 B.t8 30.5497
R2724 B.t2 B.n1207 30.5497
R2725 B.t18 B.n86 30.5497
R2726 B.n988 B.t0 29.6378
R2727 B.n1193 B.t4 29.6378
R2728 B.n1030 B.t7 28.7259
R2729 B.t1 B.n1223 28.7259
R2730 B.n964 B.t3 27.814
R2731 B.n1177 B.t6 27.814
R2732 B.n940 B.t5 25.9901
R2733 B.n1161 B.t9 25.9901
R2734 B B.n1237 18.0485
R2735 B.n884 B.n883 10.6151
R2736 B.n884 B.n536 10.6151
R2737 B.n894 B.n536 10.6151
R2738 B.n895 B.n894 10.6151
R2739 B.n896 B.n895 10.6151
R2740 B.n896 B.n528 10.6151
R2741 B.n906 B.n528 10.6151
R2742 B.n907 B.n906 10.6151
R2743 B.n908 B.n907 10.6151
R2744 B.n908 B.n520 10.6151
R2745 B.n918 B.n520 10.6151
R2746 B.n919 B.n918 10.6151
R2747 B.n920 B.n919 10.6151
R2748 B.n920 B.n512 10.6151
R2749 B.n930 B.n512 10.6151
R2750 B.n931 B.n930 10.6151
R2751 B.n932 B.n931 10.6151
R2752 B.n932 B.n504 10.6151
R2753 B.n942 B.n504 10.6151
R2754 B.n943 B.n942 10.6151
R2755 B.n944 B.n943 10.6151
R2756 B.n944 B.n496 10.6151
R2757 B.n954 B.n496 10.6151
R2758 B.n955 B.n954 10.6151
R2759 B.n956 B.n955 10.6151
R2760 B.n956 B.n488 10.6151
R2761 B.n966 B.n488 10.6151
R2762 B.n967 B.n966 10.6151
R2763 B.n968 B.n967 10.6151
R2764 B.n968 B.n480 10.6151
R2765 B.n978 B.n480 10.6151
R2766 B.n979 B.n978 10.6151
R2767 B.n980 B.n979 10.6151
R2768 B.n980 B.n472 10.6151
R2769 B.n990 B.n472 10.6151
R2770 B.n991 B.n990 10.6151
R2771 B.n992 B.n991 10.6151
R2772 B.n992 B.n464 10.6151
R2773 B.n1002 B.n464 10.6151
R2774 B.n1003 B.n1002 10.6151
R2775 B.n1004 B.n1003 10.6151
R2776 B.n1004 B.n456 10.6151
R2777 B.n1014 B.n456 10.6151
R2778 B.n1015 B.n1014 10.6151
R2779 B.n1016 B.n1015 10.6151
R2780 B.n1016 B.n448 10.6151
R2781 B.n1026 B.n448 10.6151
R2782 B.n1027 B.n1026 10.6151
R2783 B.n1028 B.n1027 10.6151
R2784 B.n1028 B.n440 10.6151
R2785 B.n1039 B.n440 10.6151
R2786 B.n1040 B.n1039 10.6151
R2787 B.n1041 B.n1040 10.6151
R2788 B.n1041 B.n0 10.6151
R2789 B.n882 B.n544 10.6151
R2790 B.n877 B.n544 10.6151
R2791 B.n877 B.n876 10.6151
R2792 B.n876 B.n875 10.6151
R2793 B.n875 B.n872 10.6151
R2794 B.n872 B.n871 10.6151
R2795 B.n871 B.n868 10.6151
R2796 B.n868 B.n867 10.6151
R2797 B.n867 B.n864 10.6151
R2798 B.n864 B.n863 10.6151
R2799 B.n863 B.n860 10.6151
R2800 B.n860 B.n859 10.6151
R2801 B.n859 B.n856 10.6151
R2802 B.n856 B.n855 10.6151
R2803 B.n855 B.n852 10.6151
R2804 B.n852 B.n851 10.6151
R2805 B.n851 B.n848 10.6151
R2806 B.n848 B.n847 10.6151
R2807 B.n847 B.n844 10.6151
R2808 B.n844 B.n843 10.6151
R2809 B.n843 B.n840 10.6151
R2810 B.n840 B.n839 10.6151
R2811 B.n839 B.n836 10.6151
R2812 B.n836 B.n835 10.6151
R2813 B.n835 B.n832 10.6151
R2814 B.n832 B.n831 10.6151
R2815 B.n831 B.n828 10.6151
R2816 B.n828 B.n827 10.6151
R2817 B.n827 B.n824 10.6151
R2818 B.n824 B.n823 10.6151
R2819 B.n823 B.n820 10.6151
R2820 B.n820 B.n819 10.6151
R2821 B.n819 B.n816 10.6151
R2822 B.n816 B.n815 10.6151
R2823 B.n815 B.n812 10.6151
R2824 B.n812 B.n811 10.6151
R2825 B.n811 B.n808 10.6151
R2826 B.n808 B.n807 10.6151
R2827 B.n807 B.n804 10.6151
R2828 B.n804 B.n803 10.6151
R2829 B.n803 B.n800 10.6151
R2830 B.n800 B.n799 10.6151
R2831 B.n799 B.n796 10.6151
R2832 B.n796 B.n795 10.6151
R2833 B.n795 B.n792 10.6151
R2834 B.n792 B.n791 10.6151
R2835 B.n791 B.n788 10.6151
R2836 B.n788 B.n787 10.6151
R2837 B.n787 B.n784 10.6151
R2838 B.n784 B.n783 10.6151
R2839 B.n783 B.n780 10.6151
R2840 B.n780 B.n779 10.6151
R2841 B.n779 B.n776 10.6151
R2842 B.n776 B.n775 10.6151
R2843 B.n775 B.n772 10.6151
R2844 B.n772 B.n771 10.6151
R2845 B.n771 B.n768 10.6151
R2846 B.n768 B.n767 10.6151
R2847 B.n767 B.n764 10.6151
R2848 B.n764 B.n763 10.6151
R2849 B.n763 B.n760 10.6151
R2850 B.n758 B.n755 10.6151
R2851 B.n755 B.n754 10.6151
R2852 B.n754 B.n751 10.6151
R2853 B.n751 B.n750 10.6151
R2854 B.n750 B.n747 10.6151
R2855 B.n747 B.n746 10.6151
R2856 B.n746 B.n743 10.6151
R2857 B.n743 B.n742 10.6151
R2858 B.n739 B.n738 10.6151
R2859 B.n738 B.n735 10.6151
R2860 B.n735 B.n734 10.6151
R2861 B.n734 B.n731 10.6151
R2862 B.n731 B.n730 10.6151
R2863 B.n730 B.n727 10.6151
R2864 B.n727 B.n726 10.6151
R2865 B.n726 B.n723 10.6151
R2866 B.n723 B.n722 10.6151
R2867 B.n722 B.n719 10.6151
R2868 B.n719 B.n718 10.6151
R2869 B.n718 B.n715 10.6151
R2870 B.n715 B.n714 10.6151
R2871 B.n714 B.n711 10.6151
R2872 B.n711 B.n710 10.6151
R2873 B.n710 B.n707 10.6151
R2874 B.n707 B.n706 10.6151
R2875 B.n706 B.n703 10.6151
R2876 B.n703 B.n702 10.6151
R2877 B.n702 B.n699 10.6151
R2878 B.n699 B.n698 10.6151
R2879 B.n698 B.n695 10.6151
R2880 B.n695 B.n694 10.6151
R2881 B.n694 B.n691 10.6151
R2882 B.n691 B.n690 10.6151
R2883 B.n690 B.n687 10.6151
R2884 B.n687 B.n686 10.6151
R2885 B.n686 B.n683 10.6151
R2886 B.n683 B.n682 10.6151
R2887 B.n682 B.n679 10.6151
R2888 B.n679 B.n678 10.6151
R2889 B.n678 B.n675 10.6151
R2890 B.n675 B.n674 10.6151
R2891 B.n674 B.n671 10.6151
R2892 B.n671 B.n670 10.6151
R2893 B.n670 B.n667 10.6151
R2894 B.n667 B.n666 10.6151
R2895 B.n666 B.n663 10.6151
R2896 B.n663 B.n662 10.6151
R2897 B.n662 B.n659 10.6151
R2898 B.n659 B.n658 10.6151
R2899 B.n658 B.n655 10.6151
R2900 B.n655 B.n654 10.6151
R2901 B.n654 B.n651 10.6151
R2902 B.n651 B.n650 10.6151
R2903 B.n650 B.n647 10.6151
R2904 B.n647 B.n646 10.6151
R2905 B.n646 B.n643 10.6151
R2906 B.n643 B.n642 10.6151
R2907 B.n642 B.n639 10.6151
R2908 B.n639 B.n638 10.6151
R2909 B.n638 B.n635 10.6151
R2910 B.n635 B.n634 10.6151
R2911 B.n634 B.n631 10.6151
R2912 B.n631 B.n630 10.6151
R2913 B.n630 B.n627 10.6151
R2914 B.n627 B.n626 10.6151
R2915 B.n626 B.n623 10.6151
R2916 B.n623 B.n622 10.6151
R2917 B.n622 B.n619 10.6151
R2918 B.n619 B.n618 10.6151
R2919 B.n888 B.n540 10.6151
R2920 B.n889 B.n888 10.6151
R2921 B.n890 B.n889 10.6151
R2922 B.n890 B.n532 10.6151
R2923 B.n900 B.n532 10.6151
R2924 B.n901 B.n900 10.6151
R2925 B.n902 B.n901 10.6151
R2926 B.n902 B.n524 10.6151
R2927 B.n912 B.n524 10.6151
R2928 B.n913 B.n912 10.6151
R2929 B.n914 B.n913 10.6151
R2930 B.n914 B.n516 10.6151
R2931 B.n924 B.n516 10.6151
R2932 B.n925 B.n924 10.6151
R2933 B.n926 B.n925 10.6151
R2934 B.n926 B.n507 10.6151
R2935 B.n936 B.n507 10.6151
R2936 B.n937 B.n936 10.6151
R2937 B.n938 B.n937 10.6151
R2938 B.n938 B.n500 10.6151
R2939 B.n948 B.n500 10.6151
R2940 B.n949 B.n948 10.6151
R2941 B.n950 B.n949 10.6151
R2942 B.n950 B.n491 10.6151
R2943 B.n960 B.n491 10.6151
R2944 B.n961 B.n960 10.6151
R2945 B.n962 B.n961 10.6151
R2946 B.n962 B.n484 10.6151
R2947 B.n972 B.n484 10.6151
R2948 B.n973 B.n972 10.6151
R2949 B.n974 B.n973 10.6151
R2950 B.n974 B.n475 10.6151
R2951 B.n984 B.n475 10.6151
R2952 B.n985 B.n984 10.6151
R2953 B.n986 B.n985 10.6151
R2954 B.n986 B.n468 10.6151
R2955 B.n996 B.n468 10.6151
R2956 B.n997 B.n996 10.6151
R2957 B.n998 B.n997 10.6151
R2958 B.n998 B.n460 10.6151
R2959 B.n1008 B.n460 10.6151
R2960 B.n1009 B.n1008 10.6151
R2961 B.n1010 B.n1009 10.6151
R2962 B.n1010 B.n452 10.6151
R2963 B.n1020 B.n452 10.6151
R2964 B.n1021 B.n1020 10.6151
R2965 B.n1022 B.n1021 10.6151
R2966 B.n1022 B.n444 10.6151
R2967 B.n1032 B.n444 10.6151
R2968 B.n1033 B.n1032 10.6151
R2969 B.n1035 B.n1033 10.6151
R2970 B.n1035 B.n1034 10.6151
R2971 B.n1034 B.n436 10.6151
R2972 B.n1046 B.n436 10.6151
R2973 B.n1047 B.n1046 10.6151
R2974 B.n1048 B.n1047 10.6151
R2975 B.n1049 B.n1048 10.6151
R2976 B.n1050 B.n1049 10.6151
R2977 B.n1053 B.n1050 10.6151
R2978 B.n1054 B.n1053 10.6151
R2979 B.n1055 B.n1054 10.6151
R2980 B.n1056 B.n1055 10.6151
R2981 B.n1058 B.n1056 10.6151
R2982 B.n1059 B.n1058 10.6151
R2983 B.n1060 B.n1059 10.6151
R2984 B.n1061 B.n1060 10.6151
R2985 B.n1063 B.n1061 10.6151
R2986 B.n1064 B.n1063 10.6151
R2987 B.n1065 B.n1064 10.6151
R2988 B.n1066 B.n1065 10.6151
R2989 B.n1068 B.n1066 10.6151
R2990 B.n1069 B.n1068 10.6151
R2991 B.n1070 B.n1069 10.6151
R2992 B.n1071 B.n1070 10.6151
R2993 B.n1073 B.n1071 10.6151
R2994 B.n1074 B.n1073 10.6151
R2995 B.n1075 B.n1074 10.6151
R2996 B.n1076 B.n1075 10.6151
R2997 B.n1078 B.n1076 10.6151
R2998 B.n1079 B.n1078 10.6151
R2999 B.n1080 B.n1079 10.6151
R3000 B.n1081 B.n1080 10.6151
R3001 B.n1083 B.n1081 10.6151
R3002 B.n1084 B.n1083 10.6151
R3003 B.n1085 B.n1084 10.6151
R3004 B.n1086 B.n1085 10.6151
R3005 B.n1088 B.n1086 10.6151
R3006 B.n1089 B.n1088 10.6151
R3007 B.n1090 B.n1089 10.6151
R3008 B.n1091 B.n1090 10.6151
R3009 B.n1093 B.n1091 10.6151
R3010 B.n1094 B.n1093 10.6151
R3011 B.n1095 B.n1094 10.6151
R3012 B.n1096 B.n1095 10.6151
R3013 B.n1098 B.n1096 10.6151
R3014 B.n1099 B.n1098 10.6151
R3015 B.n1100 B.n1099 10.6151
R3016 B.n1101 B.n1100 10.6151
R3017 B.n1103 B.n1101 10.6151
R3018 B.n1104 B.n1103 10.6151
R3019 B.n1105 B.n1104 10.6151
R3020 B.n1106 B.n1105 10.6151
R3021 B.n1108 B.n1106 10.6151
R3022 B.n1109 B.n1108 10.6151
R3023 B.n1110 B.n1109 10.6151
R3024 B.n1111 B.n1110 10.6151
R3025 B.n1113 B.n1111 10.6151
R3026 B.n1114 B.n1113 10.6151
R3027 B.n1115 B.n1114 10.6151
R3028 B.n1116 B.n1115 10.6151
R3029 B.n1117 B.n1116 10.6151
R3030 B.n1229 B.n1 10.6151
R3031 B.n1229 B.n1228 10.6151
R3032 B.n1228 B.n1227 10.6151
R3033 B.n1227 B.n10 10.6151
R3034 B.n1221 B.n10 10.6151
R3035 B.n1221 B.n1220 10.6151
R3036 B.n1220 B.n1219 10.6151
R3037 B.n1219 B.n18 10.6151
R3038 B.n1213 B.n18 10.6151
R3039 B.n1213 B.n1212 10.6151
R3040 B.n1212 B.n1211 10.6151
R3041 B.n1211 B.n25 10.6151
R3042 B.n1205 B.n25 10.6151
R3043 B.n1205 B.n1204 10.6151
R3044 B.n1204 B.n1203 10.6151
R3045 B.n1203 B.n32 10.6151
R3046 B.n1197 B.n32 10.6151
R3047 B.n1197 B.n1196 10.6151
R3048 B.n1196 B.n1195 10.6151
R3049 B.n1195 B.n39 10.6151
R3050 B.n1189 B.n39 10.6151
R3051 B.n1189 B.n1188 10.6151
R3052 B.n1188 B.n1187 10.6151
R3053 B.n1187 B.n46 10.6151
R3054 B.n1181 B.n46 10.6151
R3055 B.n1181 B.n1180 10.6151
R3056 B.n1180 B.n1179 10.6151
R3057 B.n1179 B.n53 10.6151
R3058 B.n1173 B.n53 10.6151
R3059 B.n1173 B.n1172 10.6151
R3060 B.n1172 B.n1171 10.6151
R3061 B.n1171 B.n60 10.6151
R3062 B.n1165 B.n60 10.6151
R3063 B.n1165 B.n1164 10.6151
R3064 B.n1164 B.n1163 10.6151
R3065 B.n1163 B.n67 10.6151
R3066 B.n1157 B.n67 10.6151
R3067 B.n1157 B.n1156 10.6151
R3068 B.n1156 B.n1155 10.6151
R3069 B.n1155 B.n74 10.6151
R3070 B.n1149 B.n74 10.6151
R3071 B.n1149 B.n1148 10.6151
R3072 B.n1148 B.n1147 10.6151
R3073 B.n1147 B.n81 10.6151
R3074 B.n1141 B.n81 10.6151
R3075 B.n1141 B.n1140 10.6151
R3076 B.n1140 B.n1139 10.6151
R3077 B.n1139 B.n88 10.6151
R3078 B.n1133 B.n88 10.6151
R3079 B.n1133 B.n1132 10.6151
R3080 B.n1132 B.n1131 10.6151
R3081 B.n1131 B.n95 10.6151
R3082 B.n1125 B.n95 10.6151
R3083 B.n1125 B.n1124 10.6151
R3084 B.n1123 B.n102 10.6151
R3085 B.n177 B.n102 10.6151
R3086 B.n178 B.n177 10.6151
R3087 B.n181 B.n178 10.6151
R3088 B.n182 B.n181 10.6151
R3089 B.n185 B.n182 10.6151
R3090 B.n186 B.n185 10.6151
R3091 B.n189 B.n186 10.6151
R3092 B.n190 B.n189 10.6151
R3093 B.n193 B.n190 10.6151
R3094 B.n194 B.n193 10.6151
R3095 B.n197 B.n194 10.6151
R3096 B.n198 B.n197 10.6151
R3097 B.n201 B.n198 10.6151
R3098 B.n202 B.n201 10.6151
R3099 B.n205 B.n202 10.6151
R3100 B.n206 B.n205 10.6151
R3101 B.n209 B.n206 10.6151
R3102 B.n210 B.n209 10.6151
R3103 B.n213 B.n210 10.6151
R3104 B.n214 B.n213 10.6151
R3105 B.n217 B.n214 10.6151
R3106 B.n218 B.n217 10.6151
R3107 B.n221 B.n218 10.6151
R3108 B.n222 B.n221 10.6151
R3109 B.n225 B.n222 10.6151
R3110 B.n226 B.n225 10.6151
R3111 B.n229 B.n226 10.6151
R3112 B.n230 B.n229 10.6151
R3113 B.n233 B.n230 10.6151
R3114 B.n234 B.n233 10.6151
R3115 B.n237 B.n234 10.6151
R3116 B.n238 B.n237 10.6151
R3117 B.n241 B.n238 10.6151
R3118 B.n242 B.n241 10.6151
R3119 B.n245 B.n242 10.6151
R3120 B.n246 B.n245 10.6151
R3121 B.n249 B.n246 10.6151
R3122 B.n250 B.n249 10.6151
R3123 B.n253 B.n250 10.6151
R3124 B.n254 B.n253 10.6151
R3125 B.n257 B.n254 10.6151
R3126 B.n258 B.n257 10.6151
R3127 B.n261 B.n258 10.6151
R3128 B.n262 B.n261 10.6151
R3129 B.n265 B.n262 10.6151
R3130 B.n266 B.n265 10.6151
R3131 B.n269 B.n266 10.6151
R3132 B.n270 B.n269 10.6151
R3133 B.n273 B.n270 10.6151
R3134 B.n274 B.n273 10.6151
R3135 B.n277 B.n274 10.6151
R3136 B.n278 B.n277 10.6151
R3137 B.n281 B.n278 10.6151
R3138 B.n282 B.n281 10.6151
R3139 B.n285 B.n282 10.6151
R3140 B.n286 B.n285 10.6151
R3141 B.n289 B.n286 10.6151
R3142 B.n290 B.n289 10.6151
R3143 B.n293 B.n290 10.6151
R3144 B.n294 B.n293 10.6151
R3145 B.n298 B.n297 10.6151
R3146 B.n301 B.n298 10.6151
R3147 B.n302 B.n301 10.6151
R3148 B.n305 B.n302 10.6151
R3149 B.n306 B.n305 10.6151
R3150 B.n309 B.n306 10.6151
R3151 B.n310 B.n309 10.6151
R3152 B.n313 B.n310 10.6151
R3153 B.n318 B.n315 10.6151
R3154 B.n319 B.n318 10.6151
R3155 B.n322 B.n319 10.6151
R3156 B.n323 B.n322 10.6151
R3157 B.n326 B.n323 10.6151
R3158 B.n327 B.n326 10.6151
R3159 B.n330 B.n327 10.6151
R3160 B.n331 B.n330 10.6151
R3161 B.n334 B.n331 10.6151
R3162 B.n335 B.n334 10.6151
R3163 B.n338 B.n335 10.6151
R3164 B.n339 B.n338 10.6151
R3165 B.n342 B.n339 10.6151
R3166 B.n343 B.n342 10.6151
R3167 B.n346 B.n343 10.6151
R3168 B.n347 B.n346 10.6151
R3169 B.n350 B.n347 10.6151
R3170 B.n351 B.n350 10.6151
R3171 B.n354 B.n351 10.6151
R3172 B.n355 B.n354 10.6151
R3173 B.n358 B.n355 10.6151
R3174 B.n359 B.n358 10.6151
R3175 B.n362 B.n359 10.6151
R3176 B.n363 B.n362 10.6151
R3177 B.n366 B.n363 10.6151
R3178 B.n367 B.n366 10.6151
R3179 B.n370 B.n367 10.6151
R3180 B.n371 B.n370 10.6151
R3181 B.n374 B.n371 10.6151
R3182 B.n375 B.n374 10.6151
R3183 B.n378 B.n375 10.6151
R3184 B.n379 B.n378 10.6151
R3185 B.n382 B.n379 10.6151
R3186 B.n383 B.n382 10.6151
R3187 B.n386 B.n383 10.6151
R3188 B.n387 B.n386 10.6151
R3189 B.n390 B.n387 10.6151
R3190 B.n391 B.n390 10.6151
R3191 B.n394 B.n391 10.6151
R3192 B.n395 B.n394 10.6151
R3193 B.n398 B.n395 10.6151
R3194 B.n399 B.n398 10.6151
R3195 B.n402 B.n399 10.6151
R3196 B.n403 B.n402 10.6151
R3197 B.n406 B.n403 10.6151
R3198 B.n407 B.n406 10.6151
R3199 B.n410 B.n407 10.6151
R3200 B.n411 B.n410 10.6151
R3201 B.n414 B.n411 10.6151
R3202 B.n415 B.n414 10.6151
R3203 B.n418 B.n415 10.6151
R3204 B.n419 B.n418 10.6151
R3205 B.n422 B.n419 10.6151
R3206 B.n423 B.n422 10.6151
R3207 B.n426 B.n423 10.6151
R3208 B.n427 B.n426 10.6151
R3209 B.n430 B.n427 10.6151
R3210 B.n431 B.n430 10.6151
R3211 B.n434 B.n431 10.6151
R3212 B.n435 B.n434 10.6151
R3213 B.n1118 B.n435 10.6151
R3214 B.n1237 B.n0 8.11757
R3215 B.n1237 B.n1 8.11757
R3216 B.n759 B.n758 6.5566
R3217 B.n742 B.n616 6.5566
R3218 B.n297 B.n175 6.5566
R3219 B.n314 B.n313 6.5566
R3220 B.n510 B.t5 5.01604
R3221 B.t9 B.n1160 5.01604
R3222 B.n760 B.n759 4.05904
R3223 B.n739 B.n616 4.05904
R3224 B.n294 B.n175 4.05904
R3225 B.n315 B.n314 4.05904
R3226 B.n494 B.t3 3.19221
R3227 B.t6 B.n1176 3.19221
R3228 B.t7 B.n442 2.28029
R3229 B.n1224 B.t1 2.28029
R3230 B.n478 B.t0 1.36838
R3231 B.t4 B.n1192 1.36838
R3232 B.n904 B.t11 0.456459
R3233 B.t8 B.n458 0.456459
R3234 B.n1208 B.t2 0.456459
R3235 B.n1137 B.t18 0.456459
R3236 VP.n21 VP.t5 224.499
R3237 VP.n50 VP.t1 191.681
R3238 VP.n61 VP.t4 191.681
R3239 VP.n69 VP.t7 191.681
R3240 VP.n3 VP.t0 191.681
R3241 VP.n87 VP.t6 191.681
R3242 VP.n48 VP.t2 191.681
R3243 VP.n15 VP.t8 191.681
R3244 VP.n30 VP.t3 191.681
R3245 VP.n22 VP.t9 191.681
R3246 VP.n23 VP.n20 161.3
R3247 VP.n25 VP.n24 161.3
R3248 VP.n26 VP.n19 161.3
R3249 VP.n28 VP.n27 161.3
R3250 VP.n29 VP.n18 161.3
R3251 VP.n32 VP.n31 161.3
R3252 VP.n33 VP.n17 161.3
R3253 VP.n35 VP.n34 161.3
R3254 VP.n36 VP.n16 161.3
R3255 VP.n38 VP.n37 161.3
R3256 VP.n40 VP.n39 161.3
R3257 VP.n41 VP.n14 161.3
R3258 VP.n43 VP.n42 161.3
R3259 VP.n44 VP.n13 161.3
R3260 VP.n46 VP.n45 161.3
R3261 VP.n47 VP.n12 161.3
R3262 VP.n86 VP.n0 161.3
R3263 VP.n85 VP.n84 161.3
R3264 VP.n83 VP.n1 161.3
R3265 VP.n82 VP.n81 161.3
R3266 VP.n80 VP.n2 161.3
R3267 VP.n79 VP.n78 161.3
R3268 VP.n77 VP.n76 161.3
R3269 VP.n75 VP.n4 161.3
R3270 VP.n74 VP.n73 161.3
R3271 VP.n72 VP.n5 161.3
R3272 VP.n71 VP.n70 161.3
R3273 VP.n68 VP.n6 161.3
R3274 VP.n67 VP.n66 161.3
R3275 VP.n65 VP.n7 161.3
R3276 VP.n64 VP.n63 161.3
R3277 VP.n62 VP.n8 161.3
R3278 VP.n60 VP.n59 161.3
R3279 VP.n58 VP.n9 161.3
R3280 VP.n57 VP.n56 161.3
R3281 VP.n55 VP.n10 161.3
R3282 VP.n54 VP.n53 161.3
R3283 VP.n52 VP.n11 161.3
R3284 VP.n51 VP.n50 103.416
R3285 VP.n88 VP.n87 103.416
R3286 VP.n49 VP.n48 103.416
R3287 VP.n51 VP.n49 56.9769
R3288 VP.n56 VP.n55 56.5193
R3289 VP.n81 VP.n1 56.5193
R3290 VP.n42 VP.n13 56.5193
R3291 VP.n22 VP.n21 50.2654
R3292 VP.n63 VP.n7 50.2061
R3293 VP.n75 VP.n74 50.2061
R3294 VP.n36 VP.n35 50.2061
R3295 VP.n24 VP.n19 50.2061
R3296 VP.n67 VP.n7 30.7807
R3297 VP.n74 VP.n5 30.7807
R3298 VP.n35 VP.n17 30.7807
R3299 VP.n28 VP.n19 30.7807
R3300 VP.n54 VP.n11 24.4675
R3301 VP.n55 VP.n54 24.4675
R3302 VP.n56 VP.n9 24.4675
R3303 VP.n60 VP.n9 24.4675
R3304 VP.n63 VP.n62 24.4675
R3305 VP.n68 VP.n67 24.4675
R3306 VP.n70 VP.n5 24.4675
R3307 VP.n76 VP.n75 24.4675
R3308 VP.n80 VP.n79 24.4675
R3309 VP.n81 VP.n80 24.4675
R3310 VP.n85 VP.n1 24.4675
R3311 VP.n86 VP.n85 24.4675
R3312 VP.n46 VP.n13 24.4675
R3313 VP.n47 VP.n46 24.4675
R3314 VP.n37 VP.n36 24.4675
R3315 VP.n41 VP.n40 24.4675
R3316 VP.n42 VP.n41 24.4675
R3317 VP.n29 VP.n28 24.4675
R3318 VP.n31 VP.n17 24.4675
R3319 VP.n24 VP.n23 24.4675
R3320 VP.n62 VP.n61 22.0208
R3321 VP.n76 VP.n3 22.0208
R3322 VP.n37 VP.n15 22.0208
R3323 VP.n23 VP.n22 22.0208
R3324 VP.n69 VP.n68 12.234
R3325 VP.n70 VP.n69 12.234
R3326 VP.n30 VP.n29 12.234
R3327 VP.n31 VP.n30 12.234
R3328 VP.n50 VP.n11 7.3406
R3329 VP.n87 VP.n86 7.3406
R3330 VP.n48 VP.n47 7.3406
R3331 VP.n21 VP.n20 7.01727
R3332 VP.n61 VP.n60 2.4472
R3333 VP.n79 VP.n3 2.4472
R3334 VP.n40 VP.n15 2.4472
R3335 VP.n49 VP.n12 0.278367
R3336 VP.n52 VP.n51 0.278367
R3337 VP.n88 VP.n0 0.278367
R3338 VP.n25 VP.n20 0.189894
R3339 VP.n26 VP.n25 0.189894
R3340 VP.n27 VP.n26 0.189894
R3341 VP.n27 VP.n18 0.189894
R3342 VP.n32 VP.n18 0.189894
R3343 VP.n33 VP.n32 0.189894
R3344 VP.n34 VP.n33 0.189894
R3345 VP.n34 VP.n16 0.189894
R3346 VP.n38 VP.n16 0.189894
R3347 VP.n39 VP.n38 0.189894
R3348 VP.n39 VP.n14 0.189894
R3349 VP.n43 VP.n14 0.189894
R3350 VP.n44 VP.n43 0.189894
R3351 VP.n45 VP.n44 0.189894
R3352 VP.n45 VP.n12 0.189894
R3353 VP.n53 VP.n52 0.189894
R3354 VP.n53 VP.n10 0.189894
R3355 VP.n57 VP.n10 0.189894
R3356 VP.n58 VP.n57 0.189894
R3357 VP.n59 VP.n58 0.189894
R3358 VP.n59 VP.n8 0.189894
R3359 VP.n64 VP.n8 0.189894
R3360 VP.n65 VP.n64 0.189894
R3361 VP.n66 VP.n65 0.189894
R3362 VP.n66 VP.n6 0.189894
R3363 VP.n71 VP.n6 0.189894
R3364 VP.n72 VP.n71 0.189894
R3365 VP.n73 VP.n72 0.189894
R3366 VP.n73 VP.n4 0.189894
R3367 VP.n77 VP.n4 0.189894
R3368 VP.n78 VP.n77 0.189894
R3369 VP.n78 VP.n2 0.189894
R3370 VP.n82 VP.n2 0.189894
R3371 VP.n83 VP.n82 0.189894
R3372 VP.n84 VP.n83 0.189894
R3373 VP.n84 VP.n0 0.189894
R3374 VP VP.n88 0.153454
R3375 VDD1.n100 VDD1.n0 289.615
R3376 VDD1.n207 VDD1.n107 289.615
R3377 VDD1.n101 VDD1.n100 185
R3378 VDD1.n99 VDD1.n98 185
R3379 VDD1.n4 VDD1.n3 185
R3380 VDD1.n93 VDD1.n92 185
R3381 VDD1.n91 VDD1.n90 185
R3382 VDD1.n8 VDD1.n7 185
R3383 VDD1.n85 VDD1.n84 185
R3384 VDD1.n83 VDD1.n82 185
R3385 VDD1.n81 VDD1.n11 185
R3386 VDD1.n15 VDD1.n12 185
R3387 VDD1.n76 VDD1.n75 185
R3388 VDD1.n74 VDD1.n73 185
R3389 VDD1.n17 VDD1.n16 185
R3390 VDD1.n68 VDD1.n67 185
R3391 VDD1.n66 VDD1.n65 185
R3392 VDD1.n21 VDD1.n20 185
R3393 VDD1.n60 VDD1.n59 185
R3394 VDD1.n58 VDD1.n57 185
R3395 VDD1.n25 VDD1.n24 185
R3396 VDD1.n52 VDD1.n51 185
R3397 VDD1.n50 VDD1.n49 185
R3398 VDD1.n29 VDD1.n28 185
R3399 VDD1.n44 VDD1.n43 185
R3400 VDD1.n42 VDD1.n41 185
R3401 VDD1.n33 VDD1.n32 185
R3402 VDD1.n36 VDD1.n35 185
R3403 VDD1.n142 VDD1.n141 185
R3404 VDD1.n139 VDD1.n138 185
R3405 VDD1.n148 VDD1.n147 185
R3406 VDD1.n150 VDD1.n149 185
R3407 VDD1.n135 VDD1.n134 185
R3408 VDD1.n156 VDD1.n155 185
R3409 VDD1.n158 VDD1.n157 185
R3410 VDD1.n131 VDD1.n130 185
R3411 VDD1.n164 VDD1.n163 185
R3412 VDD1.n166 VDD1.n165 185
R3413 VDD1.n127 VDD1.n126 185
R3414 VDD1.n172 VDD1.n171 185
R3415 VDD1.n174 VDD1.n173 185
R3416 VDD1.n123 VDD1.n122 185
R3417 VDD1.n180 VDD1.n179 185
R3418 VDD1.n183 VDD1.n182 185
R3419 VDD1.n181 VDD1.n119 185
R3420 VDD1.n188 VDD1.n118 185
R3421 VDD1.n190 VDD1.n189 185
R3422 VDD1.n192 VDD1.n191 185
R3423 VDD1.n115 VDD1.n114 185
R3424 VDD1.n198 VDD1.n197 185
R3425 VDD1.n200 VDD1.n199 185
R3426 VDD1.n111 VDD1.n110 185
R3427 VDD1.n206 VDD1.n205 185
R3428 VDD1.n208 VDD1.n207 185
R3429 VDD1.t4 VDD1.n34 147.659
R3430 VDD1.t8 VDD1.n140 147.659
R3431 VDD1.n100 VDD1.n99 104.615
R3432 VDD1.n99 VDD1.n3 104.615
R3433 VDD1.n92 VDD1.n3 104.615
R3434 VDD1.n92 VDD1.n91 104.615
R3435 VDD1.n91 VDD1.n7 104.615
R3436 VDD1.n84 VDD1.n7 104.615
R3437 VDD1.n84 VDD1.n83 104.615
R3438 VDD1.n83 VDD1.n11 104.615
R3439 VDD1.n15 VDD1.n11 104.615
R3440 VDD1.n75 VDD1.n15 104.615
R3441 VDD1.n75 VDD1.n74 104.615
R3442 VDD1.n74 VDD1.n16 104.615
R3443 VDD1.n67 VDD1.n16 104.615
R3444 VDD1.n67 VDD1.n66 104.615
R3445 VDD1.n66 VDD1.n20 104.615
R3446 VDD1.n59 VDD1.n20 104.615
R3447 VDD1.n59 VDD1.n58 104.615
R3448 VDD1.n58 VDD1.n24 104.615
R3449 VDD1.n51 VDD1.n24 104.615
R3450 VDD1.n51 VDD1.n50 104.615
R3451 VDD1.n50 VDD1.n28 104.615
R3452 VDD1.n43 VDD1.n28 104.615
R3453 VDD1.n43 VDD1.n42 104.615
R3454 VDD1.n42 VDD1.n32 104.615
R3455 VDD1.n35 VDD1.n32 104.615
R3456 VDD1.n141 VDD1.n138 104.615
R3457 VDD1.n148 VDD1.n138 104.615
R3458 VDD1.n149 VDD1.n148 104.615
R3459 VDD1.n149 VDD1.n134 104.615
R3460 VDD1.n156 VDD1.n134 104.615
R3461 VDD1.n157 VDD1.n156 104.615
R3462 VDD1.n157 VDD1.n130 104.615
R3463 VDD1.n164 VDD1.n130 104.615
R3464 VDD1.n165 VDD1.n164 104.615
R3465 VDD1.n165 VDD1.n126 104.615
R3466 VDD1.n172 VDD1.n126 104.615
R3467 VDD1.n173 VDD1.n172 104.615
R3468 VDD1.n173 VDD1.n122 104.615
R3469 VDD1.n180 VDD1.n122 104.615
R3470 VDD1.n182 VDD1.n180 104.615
R3471 VDD1.n182 VDD1.n181 104.615
R3472 VDD1.n181 VDD1.n118 104.615
R3473 VDD1.n190 VDD1.n118 104.615
R3474 VDD1.n191 VDD1.n190 104.615
R3475 VDD1.n191 VDD1.n114 104.615
R3476 VDD1.n198 VDD1.n114 104.615
R3477 VDD1.n199 VDD1.n198 104.615
R3478 VDD1.n199 VDD1.n110 104.615
R3479 VDD1.n206 VDD1.n110 104.615
R3480 VDD1.n207 VDD1.n206 104.615
R3481 VDD1.n215 VDD1.n214 60.179
R3482 VDD1.n106 VDD1.n105 58.4887
R3483 VDD1.n213 VDD1.n212 58.4887
R3484 VDD1.n217 VDD1.n216 58.4885
R3485 VDD1.n217 VDD1.n215 52.7681
R3486 VDD1.n35 VDD1.t4 52.3082
R3487 VDD1.n141 VDD1.t8 52.3082
R3488 VDD1.n106 VDD1.n104 49.0584
R3489 VDD1.n213 VDD1.n211 49.0584
R3490 VDD1.n36 VDD1.n34 15.6677
R3491 VDD1.n142 VDD1.n140 15.6677
R3492 VDD1.n82 VDD1.n81 13.1884
R3493 VDD1.n189 VDD1.n188 13.1884
R3494 VDD1.n85 VDD1.n10 12.8005
R3495 VDD1.n80 VDD1.n12 12.8005
R3496 VDD1.n37 VDD1.n33 12.8005
R3497 VDD1.n143 VDD1.n139 12.8005
R3498 VDD1.n187 VDD1.n119 12.8005
R3499 VDD1.n192 VDD1.n117 12.8005
R3500 VDD1.n86 VDD1.n8 12.0247
R3501 VDD1.n77 VDD1.n76 12.0247
R3502 VDD1.n41 VDD1.n40 12.0247
R3503 VDD1.n147 VDD1.n146 12.0247
R3504 VDD1.n184 VDD1.n183 12.0247
R3505 VDD1.n193 VDD1.n115 12.0247
R3506 VDD1.n90 VDD1.n89 11.249
R3507 VDD1.n73 VDD1.n14 11.249
R3508 VDD1.n44 VDD1.n31 11.249
R3509 VDD1.n150 VDD1.n137 11.249
R3510 VDD1.n179 VDD1.n121 11.249
R3511 VDD1.n197 VDD1.n196 11.249
R3512 VDD1.n93 VDD1.n6 10.4732
R3513 VDD1.n72 VDD1.n17 10.4732
R3514 VDD1.n45 VDD1.n29 10.4732
R3515 VDD1.n151 VDD1.n135 10.4732
R3516 VDD1.n178 VDD1.n123 10.4732
R3517 VDD1.n200 VDD1.n113 10.4732
R3518 VDD1.n94 VDD1.n4 9.69747
R3519 VDD1.n69 VDD1.n68 9.69747
R3520 VDD1.n49 VDD1.n48 9.69747
R3521 VDD1.n155 VDD1.n154 9.69747
R3522 VDD1.n175 VDD1.n174 9.69747
R3523 VDD1.n201 VDD1.n111 9.69747
R3524 VDD1.n104 VDD1.n103 9.45567
R3525 VDD1.n211 VDD1.n210 9.45567
R3526 VDD1.n62 VDD1.n61 9.3005
R3527 VDD1.n64 VDD1.n63 9.3005
R3528 VDD1.n19 VDD1.n18 9.3005
R3529 VDD1.n70 VDD1.n69 9.3005
R3530 VDD1.n72 VDD1.n71 9.3005
R3531 VDD1.n14 VDD1.n13 9.3005
R3532 VDD1.n78 VDD1.n77 9.3005
R3533 VDD1.n80 VDD1.n79 9.3005
R3534 VDD1.n103 VDD1.n102 9.3005
R3535 VDD1.n2 VDD1.n1 9.3005
R3536 VDD1.n97 VDD1.n96 9.3005
R3537 VDD1.n95 VDD1.n94 9.3005
R3538 VDD1.n6 VDD1.n5 9.3005
R3539 VDD1.n89 VDD1.n88 9.3005
R3540 VDD1.n87 VDD1.n86 9.3005
R3541 VDD1.n10 VDD1.n9 9.3005
R3542 VDD1.n23 VDD1.n22 9.3005
R3543 VDD1.n56 VDD1.n55 9.3005
R3544 VDD1.n54 VDD1.n53 9.3005
R3545 VDD1.n27 VDD1.n26 9.3005
R3546 VDD1.n48 VDD1.n47 9.3005
R3547 VDD1.n46 VDD1.n45 9.3005
R3548 VDD1.n31 VDD1.n30 9.3005
R3549 VDD1.n40 VDD1.n39 9.3005
R3550 VDD1.n38 VDD1.n37 9.3005
R3551 VDD1.n109 VDD1.n108 9.3005
R3552 VDD1.n204 VDD1.n203 9.3005
R3553 VDD1.n202 VDD1.n201 9.3005
R3554 VDD1.n113 VDD1.n112 9.3005
R3555 VDD1.n196 VDD1.n195 9.3005
R3556 VDD1.n194 VDD1.n193 9.3005
R3557 VDD1.n117 VDD1.n116 9.3005
R3558 VDD1.n162 VDD1.n161 9.3005
R3559 VDD1.n160 VDD1.n159 9.3005
R3560 VDD1.n133 VDD1.n132 9.3005
R3561 VDD1.n154 VDD1.n153 9.3005
R3562 VDD1.n152 VDD1.n151 9.3005
R3563 VDD1.n137 VDD1.n136 9.3005
R3564 VDD1.n146 VDD1.n145 9.3005
R3565 VDD1.n144 VDD1.n143 9.3005
R3566 VDD1.n129 VDD1.n128 9.3005
R3567 VDD1.n168 VDD1.n167 9.3005
R3568 VDD1.n170 VDD1.n169 9.3005
R3569 VDD1.n125 VDD1.n124 9.3005
R3570 VDD1.n176 VDD1.n175 9.3005
R3571 VDD1.n178 VDD1.n177 9.3005
R3572 VDD1.n121 VDD1.n120 9.3005
R3573 VDD1.n185 VDD1.n184 9.3005
R3574 VDD1.n187 VDD1.n186 9.3005
R3575 VDD1.n210 VDD1.n209 9.3005
R3576 VDD1.n98 VDD1.n97 8.92171
R3577 VDD1.n65 VDD1.n19 8.92171
R3578 VDD1.n52 VDD1.n27 8.92171
R3579 VDD1.n158 VDD1.n133 8.92171
R3580 VDD1.n171 VDD1.n125 8.92171
R3581 VDD1.n205 VDD1.n204 8.92171
R3582 VDD1.n101 VDD1.n2 8.14595
R3583 VDD1.n64 VDD1.n21 8.14595
R3584 VDD1.n53 VDD1.n25 8.14595
R3585 VDD1.n159 VDD1.n131 8.14595
R3586 VDD1.n170 VDD1.n127 8.14595
R3587 VDD1.n208 VDD1.n109 8.14595
R3588 VDD1.n102 VDD1.n0 7.3702
R3589 VDD1.n61 VDD1.n60 7.3702
R3590 VDD1.n57 VDD1.n56 7.3702
R3591 VDD1.n163 VDD1.n162 7.3702
R3592 VDD1.n167 VDD1.n166 7.3702
R3593 VDD1.n209 VDD1.n107 7.3702
R3594 VDD1.n104 VDD1.n0 6.59444
R3595 VDD1.n60 VDD1.n23 6.59444
R3596 VDD1.n57 VDD1.n23 6.59444
R3597 VDD1.n163 VDD1.n129 6.59444
R3598 VDD1.n166 VDD1.n129 6.59444
R3599 VDD1.n211 VDD1.n107 6.59444
R3600 VDD1.n102 VDD1.n101 5.81868
R3601 VDD1.n61 VDD1.n21 5.81868
R3602 VDD1.n56 VDD1.n25 5.81868
R3603 VDD1.n162 VDD1.n131 5.81868
R3604 VDD1.n167 VDD1.n127 5.81868
R3605 VDD1.n209 VDD1.n208 5.81868
R3606 VDD1.n98 VDD1.n2 5.04292
R3607 VDD1.n65 VDD1.n64 5.04292
R3608 VDD1.n53 VDD1.n52 5.04292
R3609 VDD1.n159 VDD1.n158 5.04292
R3610 VDD1.n171 VDD1.n170 5.04292
R3611 VDD1.n205 VDD1.n109 5.04292
R3612 VDD1.n38 VDD1.n34 4.38563
R3613 VDD1.n144 VDD1.n140 4.38563
R3614 VDD1.n97 VDD1.n4 4.26717
R3615 VDD1.n68 VDD1.n19 4.26717
R3616 VDD1.n49 VDD1.n27 4.26717
R3617 VDD1.n155 VDD1.n133 4.26717
R3618 VDD1.n174 VDD1.n125 4.26717
R3619 VDD1.n204 VDD1.n111 4.26717
R3620 VDD1.n94 VDD1.n93 3.49141
R3621 VDD1.n69 VDD1.n17 3.49141
R3622 VDD1.n48 VDD1.n29 3.49141
R3623 VDD1.n154 VDD1.n135 3.49141
R3624 VDD1.n175 VDD1.n123 3.49141
R3625 VDD1.n201 VDD1.n200 3.49141
R3626 VDD1.n90 VDD1.n6 2.71565
R3627 VDD1.n73 VDD1.n72 2.71565
R3628 VDD1.n45 VDD1.n44 2.71565
R3629 VDD1.n151 VDD1.n150 2.71565
R3630 VDD1.n179 VDD1.n178 2.71565
R3631 VDD1.n197 VDD1.n113 2.71565
R3632 VDD1.n89 VDD1.n8 1.93989
R3633 VDD1.n76 VDD1.n14 1.93989
R3634 VDD1.n41 VDD1.n31 1.93989
R3635 VDD1.n147 VDD1.n137 1.93989
R3636 VDD1.n183 VDD1.n121 1.93989
R3637 VDD1.n196 VDD1.n115 1.93989
R3638 VDD1 VDD1.n217 1.688
R3639 VDD1.n86 VDD1.n85 1.16414
R3640 VDD1.n77 VDD1.n12 1.16414
R3641 VDD1.n40 VDD1.n33 1.16414
R3642 VDD1.n146 VDD1.n139 1.16414
R3643 VDD1.n184 VDD1.n119 1.16414
R3644 VDD1.n193 VDD1.n192 1.16414
R3645 VDD1.n216 VDD1.t1 1.0509
R3646 VDD1.n216 VDD1.t7 1.0509
R3647 VDD1.n105 VDD1.t0 1.0509
R3648 VDD1.n105 VDD1.t6 1.0509
R3649 VDD1.n214 VDD1.t9 1.0509
R3650 VDD1.n214 VDD1.t3 1.0509
R3651 VDD1.n212 VDD1.t5 1.0509
R3652 VDD1.n212 VDD1.t2 1.0509
R3653 VDD1 VDD1.n106 0.640586
R3654 VDD1.n215 VDD1.n213 0.527051
R3655 VDD1.n82 VDD1.n10 0.388379
R3656 VDD1.n81 VDD1.n80 0.388379
R3657 VDD1.n37 VDD1.n36 0.388379
R3658 VDD1.n143 VDD1.n142 0.388379
R3659 VDD1.n188 VDD1.n187 0.388379
R3660 VDD1.n189 VDD1.n117 0.388379
R3661 VDD1.n103 VDD1.n1 0.155672
R3662 VDD1.n96 VDD1.n1 0.155672
R3663 VDD1.n96 VDD1.n95 0.155672
R3664 VDD1.n95 VDD1.n5 0.155672
R3665 VDD1.n88 VDD1.n5 0.155672
R3666 VDD1.n88 VDD1.n87 0.155672
R3667 VDD1.n87 VDD1.n9 0.155672
R3668 VDD1.n79 VDD1.n9 0.155672
R3669 VDD1.n79 VDD1.n78 0.155672
R3670 VDD1.n78 VDD1.n13 0.155672
R3671 VDD1.n71 VDD1.n13 0.155672
R3672 VDD1.n71 VDD1.n70 0.155672
R3673 VDD1.n70 VDD1.n18 0.155672
R3674 VDD1.n63 VDD1.n18 0.155672
R3675 VDD1.n63 VDD1.n62 0.155672
R3676 VDD1.n62 VDD1.n22 0.155672
R3677 VDD1.n55 VDD1.n22 0.155672
R3678 VDD1.n55 VDD1.n54 0.155672
R3679 VDD1.n54 VDD1.n26 0.155672
R3680 VDD1.n47 VDD1.n26 0.155672
R3681 VDD1.n47 VDD1.n46 0.155672
R3682 VDD1.n46 VDD1.n30 0.155672
R3683 VDD1.n39 VDD1.n30 0.155672
R3684 VDD1.n39 VDD1.n38 0.155672
R3685 VDD1.n145 VDD1.n144 0.155672
R3686 VDD1.n145 VDD1.n136 0.155672
R3687 VDD1.n152 VDD1.n136 0.155672
R3688 VDD1.n153 VDD1.n152 0.155672
R3689 VDD1.n153 VDD1.n132 0.155672
R3690 VDD1.n160 VDD1.n132 0.155672
R3691 VDD1.n161 VDD1.n160 0.155672
R3692 VDD1.n161 VDD1.n128 0.155672
R3693 VDD1.n168 VDD1.n128 0.155672
R3694 VDD1.n169 VDD1.n168 0.155672
R3695 VDD1.n169 VDD1.n124 0.155672
R3696 VDD1.n176 VDD1.n124 0.155672
R3697 VDD1.n177 VDD1.n176 0.155672
R3698 VDD1.n177 VDD1.n120 0.155672
R3699 VDD1.n185 VDD1.n120 0.155672
R3700 VDD1.n186 VDD1.n185 0.155672
R3701 VDD1.n186 VDD1.n116 0.155672
R3702 VDD1.n194 VDD1.n116 0.155672
R3703 VDD1.n195 VDD1.n194 0.155672
R3704 VDD1.n195 VDD1.n112 0.155672
R3705 VDD1.n202 VDD1.n112 0.155672
R3706 VDD1.n203 VDD1.n202 0.155672
R3707 VDD1.n203 VDD1.n108 0.155672
R3708 VDD1.n210 VDD1.n108 0.155672
C0 VDD1 VN 0.152866f
C1 VTAIL VDD1 13.6783f
C2 VP VDD2 0.554863f
C3 VN VDD2 16.1463f
C4 VTAIL VDD2 13.7257f
C5 VP VN 9.33215f
C6 VTAIL VP 16.4059f
C7 VDD1 VDD2 2.02583f
C8 VTAIL VN 16.3915f
C9 VDD1 VP 16.543098f
C10 VDD2 B 8.15519f
C11 VDD1 B 8.127254f
C12 VTAIL B 10.740474f
C13 VN B 17.648548f
C14 VP B 16.029875f
C15 VDD1.n0 B 0.031935f
C16 VDD1.n1 B 0.02351f
C17 VDD1.n2 B 0.012633f
C18 VDD1.n3 B 0.02986f
C19 VDD1.n4 B 0.013376f
C20 VDD1.n5 B 0.02351f
C21 VDD1.n6 B 0.012633f
C22 VDD1.n7 B 0.02986f
C23 VDD1.n8 B 0.013376f
C24 VDD1.n9 B 0.02351f
C25 VDD1.n10 B 0.012633f
C26 VDD1.n11 B 0.02986f
C27 VDD1.n12 B 0.013376f
C28 VDD1.n13 B 0.02351f
C29 VDD1.n14 B 0.012633f
C30 VDD1.n15 B 0.02986f
C31 VDD1.n16 B 0.02986f
C32 VDD1.n17 B 0.013376f
C33 VDD1.n18 B 0.02351f
C34 VDD1.n19 B 0.012633f
C35 VDD1.n20 B 0.02986f
C36 VDD1.n21 B 0.013376f
C37 VDD1.n22 B 0.02351f
C38 VDD1.n23 B 0.012633f
C39 VDD1.n24 B 0.02986f
C40 VDD1.n25 B 0.013376f
C41 VDD1.n26 B 0.02351f
C42 VDD1.n27 B 0.012633f
C43 VDD1.n28 B 0.02986f
C44 VDD1.n29 B 0.013376f
C45 VDD1.n30 B 0.02351f
C46 VDD1.n31 B 0.012633f
C47 VDD1.n32 B 0.02986f
C48 VDD1.n33 B 0.013376f
C49 VDD1.n34 B 0.176029f
C50 VDD1.t4 B 0.049546f
C51 VDD1.n35 B 0.022395f
C52 VDD1.n36 B 0.017639f
C53 VDD1.n37 B 0.012633f
C54 VDD1.n38 B 1.9444f
C55 VDD1.n39 B 0.02351f
C56 VDD1.n40 B 0.012633f
C57 VDD1.n41 B 0.013376f
C58 VDD1.n42 B 0.02986f
C59 VDD1.n43 B 0.02986f
C60 VDD1.n44 B 0.013376f
C61 VDD1.n45 B 0.012633f
C62 VDD1.n46 B 0.02351f
C63 VDD1.n47 B 0.02351f
C64 VDD1.n48 B 0.012633f
C65 VDD1.n49 B 0.013376f
C66 VDD1.n50 B 0.02986f
C67 VDD1.n51 B 0.02986f
C68 VDD1.n52 B 0.013376f
C69 VDD1.n53 B 0.012633f
C70 VDD1.n54 B 0.02351f
C71 VDD1.n55 B 0.02351f
C72 VDD1.n56 B 0.012633f
C73 VDD1.n57 B 0.013376f
C74 VDD1.n58 B 0.02986f
C75 VDD1.n59 B 0.02986f
C76 VDD1.n60 B 0.013376f
C77 VDD1.n61 B 0.012633f
C78 VDD1.n62 B 0.02351f
C79 VDD1.n63 B 0.02351f
C80 VDD1.n64 B 0.012633f
C81 VDD1.n65 B 0.013376f
C82 VDD1.n66 B 0.02986f
C83 VDD1.n67 B 0.02986f
C84 VDD1.n68 B 0.013376f
C85 VDD1.n69 B 0.012633f
C86 VDD1.n70 B 0.02351f
C87 VDD1.n71 B 0.02351f
C88 VDD1.n72 B 0.012633f
C89 VDD1.n73 B 0.013376f
C90 VDD1.n74 B 0.02986f
C91 VDD1.n75 B 0.02986f
C92 VDD1.n76 B 0.013376f
C93 VDD1.n77 B 0.012633f
C94 VDD1.n78 B 0.02351f
C95 VDD1.n79 B 0.02351f
C96 VDD1.n80 B 0.012633f
C97 VDD1.n81 B 0.013005f
C98 VDD1.n82 B 0.013005f
C99 VDD1.n83 B 0.02986f
C100 VDD1.n84 B 0.02986f
C101 VDD1.n85 B 0.013376f
C102 VDD1.n86 B 0.012633f
C103 VDD1.n87 B 0.02351f
C104 VDD1.n88 B 0.02351f
C105 VDD1.n89 B 0.012633f
C106 VDD1.n90 B 0.013376f
C107 VDD1.n91 B 0.02986f
C108 VDD1.n92 B 0.02986f
C109 VDD1.n93 B 0.013376f
C110 VDD1.n94 B 0.012633f
C111 VDD1.n95 B 0.02351f
C112 VDD1.n96 B 0.02351f
C113 VDD1.n97 B 0.012633f
C114 VDD1.n98 B 0.013376f
C115 VDD1.n99 B 0.02986f
C116 VDD1.n100 B 0.062679f
C117 VDD1.n101 B 0.013376f
C118 VDD1.n102 B 0.012633f
C119 VDD1.n103 B 0.050809f
C120 VDD1.n104 B 0.061438f
C121 VDD1.t0 B 0.350197f
C122 VDD1.t6 B 0.350197f
C123 VDD1.n105 B 3.19278f
C124 VDD1.n106 B 0.633188f
C125 VDD1.n107 B 0.031935f
C126 VDD1.n108 B 0.02351f
C127 VDD1.n109 B 0.012633f
C128 VDD1.n110 B 0.02986f
C129 VDD1.n111 B 0.013376f
C130 VDD1.n112 B 0.02351f
C131 VDD1.n113 B 0.012633f
C132 VDD1.n114 B 0.02986f
C133 VDD1.n115 B 0.013376f
C134 VDD1.n116 B 0.02351f
C135 VDD1.n117 B 0.012633f
C136 VDD1.n118 B 0.02986f
C137 VDD1.n119 B 0.013376f
C138 VDD1.n120 B 0.02351f
C139 VDD1.n121 B 0.012633f
C140 VDD1.n122 B 0.02986f
C141 VDD1.n123 B 0.013376f
C142 VDD1.n124 B 0.02351f
C143 VDD1.n125 B 0.012633f
C144 VDD1.n126 B 0.02986f
C145 VDD1.n127 B 0.013376f
C146 VDD1.n128 B 0.02351f
C147 VDD1.n129 B 0.012633f
C148 VDD1.n130 B 0.02986f
C149 VDD1.n131 B 0.013376f
C150 VDD1.n132 B 0.02351f
C151 VDD1.n133 B 0.012633f
C152 VDD1.n134 B 0.02986f
C153 VDD1.n135 B 0.013376f
C154 VDD1.n136 B 0.02351f
C155 VDD1.n137 B 0.012633f
C156 VDD1.n138 B 0.02986f
C157 VDD1.n139 B 0.013376f
C158 VDD1.n140 B 0.176029f
C159 VDD1.t8 B 0.049546f
C160 VDD1.n141 B 0.022395f
C161 VDD1.n142 B 0.017639f
C162 VDD1.n143 B 0.012633f
C163 VDD1.n144 B 1.9444f
C164 VDD1.n145 B 0.02351f
C165 VDD1.n146 B 0.012633f
C166 VDD1.n147 B 0.013376f
C167 VDD1.n148 B 0.02986f
C168 VDD1.n149 B 0.02986f
C169 VDD1.n150 B 0.013376f
C170 VDD1.n151 B 0.012633f
C171 VDD1.n152 B 0.02351f
C172 VDD1.n153 B 0.02351f
C173 VDD1.n154 B 0.012633f
C174 VDD1.n155 B 0.013376f
C175 VDD1.n156 B 0.02986f
C176 VDD1.n157 B 0.02986f
C177 VDD1.n158 B 0.013376f
C178 VDD1.n159 B 0.012633f
C179 VDD1.n160 B 0.02351f
C180 VDD1.n161 B 0.02351f
C181 VDD1.n162 B 0.012633f
C182 VDD1.n163 B 0.013376f
C183 VDD1.n164 B 0.02986f
C184 VDD1.n165 B 0.02986f
C185 VDD1.n166 B 0.013376f
C186 VDD1.n167 B 0.012633f
C187 VDD1.n168 B 0.02351f
C188 VDD1.n169 B 0.02351f
C189 VDD1.n170 B 0.012633f
C190 VDD1.n171 B 0.013376f
C191 VDD1.n172 B 0.02986f
C192 VDD1.n173 B 0.02986f
C193 VDD1.n174 B 0.013376f
C194 VDD1.n175 B 0.012633f
C195 VDD1.n176 B 0.02351f
C196 VDD1.n177 B 0.02351f
C197 VDD1.n178 B 0.012633f
C198 VDD1.n179 B 0.013376f
C199 VDD1.n180 B 0.02986f
C200 VDD1.n181 B 0.02986f
C201 VDD1.n182 B 0.02986f
C202 VDD1.n183 B 0.013376f
C203 VDD1.n184 B 0.012633f
C204 VDD1.n185 B 0.02351f
C205 VDD1.n186 B 0.02351f
C206 VDD1.n187 B 0.012633f
C207 VDD1.n188 B 0.013005f
C208 VDD1.n189 B 0.013005f
C209 VDD1.n190 B 0.02986f
C210 VDD1.n191 B 0.02986f
C211 VDD1.n192 B 0.013376f
C212 VDD1.n193 B 0.012633f
C213 VDD1.n194 B 0.02351f
C214 VDD1.n195 B 0.02351f
C215 VDD1.n196 B 0.012633f
C216 VDD1.n197 B 0.013376f
C217 VDD1.n198 B 0.02986f
C218 VDD1.n199 B 0.02986f
C219 VDD1.n200 B 0.013376f
C220 VDD1.n201 B 0.012633f
C221 VDD1.n202 B 0.02351f
C222 VDD1.n203 B 0.02351f
C223 VDD1.n204 B 0.012633f
C224 VDD1.n205 B 0.013376f
C225 VDD1.n206 B 0.02986f
C226 VDD1.n207 B 0.062679f
C227 VDD1.n208 B 0.013376f
C228 VDD1.n209 B 0.012633f
C229 VDD1.n210 B 0.050809f
C230 VDD1.n211 B 0.061438f
C231 VDD1.t5 B 0.350197f
C232 VDD1.t2 B 0.350197f
C233 VDD1.n212 B 3.19278f
C234 VDD1.n213 B 0.625624f
C235 VDD1.t9 B 0.350197f
C236 VDD1.t3 B 0.350197f
C237 VDD1.n214 B 3.2072f
C238 VDD1.n215 B 3.1427f
C239 VDD1.t1 B 0.350197f
C240 VDD1.t7 B 0.350197f
C241 VDD1.n216 B 3.19277f
C242 VDD1.n217 B 3.38763f
C243 VP.n0 B 0.028968f
C244 VP.t6 B 2.70227f
C245 VP.n1 B 0.029014f
C246 VP.n2 B 0.021972f
C247 VP.t0 B 2.70227f
C248 VP.n3 B 0.93719f
C249 VP.n4 B 0.021972f
C250 VP.n5 B 0.044018f
C251 VP.n6 B 0.021972f
C252 VP.t7 B 2.70227f
C253 VP.n7 B 0.020757f
C254 VP.n8 B 0.021972f
C255 VP.t4 B 2.70227f
C256 VP.n9 B 0.040951f
C257 VP.n10 B 0.021972f
C258 VP.n11 B 0.026799f
C259 VP.n12 B 0.028968f
C260 VP.t2 B 2.70227f
C261 VP.n13 B 0.029014f
C262 VP.n14 B 0.021972f
C263 VP.t8 B 2.70227f
C264 VP.n15 B 0.93719f
C265 VP.n16 B 0.021972f
C266 VP.n17 B 0.044018f
C267 VP.n18 B 0.021972f
C268 VP.t3 B 2.70227f
C269 VP.n19 B 0.020757f
C270 VP.n20 B 0.207045f
C271 VP.t9 B 2.70227f
C272 VP.t5 B 2.85776f
C273 VP.n21 B 0.983888f
C274 VP.n22 B 1.00633f
C275 VP.n23 B 0.038929f
C276 VP.n24 B 0.040327f
C277 VP.n25 B 0.021972f
C278 VP.n26 B 0.021972f
C279 VP.n27 B 0.021972f
C280 VP.n28 B 0.044018f
C281 VP.n29 B 0.030842f
C282 VP.n30 B 0.93719f
C283 VP.n31 B 0.030842f
C284 VP.n32 B 0.021972f
C285 VP.n33 B 0.021972f
C286 VP.n34 B 0.021972f
C287 VP.n35 B 0.020757f
C288 VP.n36 B 0.040327f
C289 VP.n37 B 0.038929f
C290 VP.n38 B 0.021972f
C291 VP.n39 B 0.021972f
C292 VP.n40 B 0.022755f
C293 VP.n41 B 0.040951f
C294 VP.n42 B 0.035137f
C295 VP.n43 B 0.021972f
C296 VP.n44 B 0.021972f
C297 VP.n45 B 0.021972f
C298 VP.n46 B 0.040951f
C299 VP.n47 B 0.026799f
C300 VP.n48 B 1.00095f
C301 VP.n49 B 1.4717f
C302 VP.t1 B 2.70227f
C303 VP.n50 B 1.00095f
C304 VP.n51 B 1.48556f
C305 VP.n52 B 0.028968f
C306 VP.n53 B 0.021972f
C307 VP.n54 B 0.040951f
C308 VP.n55 B 0.029014f
C309 VP.n56 B 0.035137f
C310 VP.n57 B 0.021972f
C311 VP.n58 B 0.021972f
C312 VP.n59 B 0.021972f
C313 VP.n60 B 0.022755f
C314 VP.n61 B 0.93719f
C315 VP.n62 B 0.038929f
C316 VP.n63 B 0.040327f
C317 VP.n64 B 0.021972f
C318 VP.n65 B 0.021972f
C319 VP.n66 B 0.021972f
C320 VP.n67 B 0.044018f
C321 VP.n68 B 0.030842f
C322 VP.n69 B 0.93719f
C323 VP.n70 B 0.030842f
C324 VP.n71 B 0.021972f
C325 VP.n72 B 0.021972f
C326 VP.n73 B 0.021972f
C327 VP.n74 B 0.020757f
C328 VP.n75 B 0.040327f
C329 VP.n76 B 0.038929f
C330 VP.n77 B 0.021972f
C331 VP.n78 B 0.021972f
C332 VP.n79 B 0.022755f
C333 VP.n80 B 0.040951f
C334 VP.n81 B 0.035137f
C335 VP.n82 B 0.021972f
C336 VP.n83 B 0.021972f
C337 VP.n84 B 0.021972f
C338 VP.n85 B 0.040951f
C339 VP.n86 B 0.026799f
C340 VP.n87 B 1.00095f
C341 VP.n88 B 0.03543f
C342 VDD2.n0 B 0.031623f
C343 VDD2.n1 B 0.02328f
C344 VDD2.n2 B 0.01251f
C345 VDD2.n3 B 0.029569f
C346 VDD2.n4 B 0.013246f
C347 VDD2.n5 B 0.02328f
C348 VDD2.n6 B 0.01251f
C349 VDD2.n7 B 0.029569f
C350 VDD2.n8 B 0.013246f
C351 VDD2.n9 B 0.02328f
C352 VDD2.n10 B 0.01251f
C353 VDD2.n11 B 0.029569f
C354 VDD2.n12 B 0.013246f
C355 VDD2.n13 B 0.02328f
C356 VDD2.n14 B 0.01251f
C357 VDD2.n15 B 0.029569f
C358 VDD2.n16 B 0.013246f
C359 VDD2.n17 B 0.02328f
C360 VDD2.n18 B 0.01251f
C361 VDD2.n19 B 0.029569f
C362 VDD2.n20 B 0.013246f
C363 VDD2.n21 B 0.02328f
C364 VDD2.n22 B 0.01251f
C365 VDD2.n23 B 0.029569f
C366 VDD2.n24 B 0.013246f
C367 VDD2.n25 B 0.02328f
C368 VDD2.n26 B 0.01251f
C369 VDD2.n27 B 0.029569f
C370 VDD2.n28 B 0.013246f
C371 VDD2.n29 B 0.02328f
C372 VDD2.n30 B 0.01251f
C373 VDD2.n31 B 0.029569f
C374 VDD2.n32 B 0.013246f
C375 VDD2.n33 B 0.174312f
C376 VDD2.t0 B 0.049063f
C377 VDD2.n34 B 0.022177f
C378 VDD2.n35 B 0.017467f
C379 VDD2.n36 B 0.01251f
C380 VDD2.n37 B 1.92543f
C381 VDD2.n38 B 0.02328f
C382 VDD2.n39 B 0.01251f
C383 VDD2.n40 B 0.013246f
C384 VDD2.n41 B 0.029569f
C385 VDD2.n42 B 0.029569f
C386 VDD2.n43 B 0.013246f
C387 VDD2.n44 B 0.01251f
C388 VDD2.n45 B 0.02328f
C389 VDD2.n46 B 0.02328f
C390 VDD2.n47 B 0.01251f
C391 VDD2.n48 B 0.013246f
C392 VDD2.n49 B 0.029569f
C393 VDD2.n50 B 0.029569f
C394 VDD2.n51 B 0.013246f
C395 VDD2.n52 B 0.01251f
C396 VDD2.n53 B 0.02328f
C397 VDD2.n54 B 0.02328f
C398 VDD2.n55 B 0.01251f
C399 VDD2.n56 B 0.013246f
C400 VDD2.n57 B 0.029569f
C401 VDD2.n58 B 0.029569f
C402 VDD2.n59 B 0.013246f
C403 VDD2.n60 B 0.01251f
C404 VDD2.n61 B 0.02328f
C405 VDD2.n62 B 0.02328f
C406 VDD2.n63 B 0.01251f
C407 VDD2.n64 B 0.013246f
C408 VDD2.n65 B 0.029569f
C409 VDD2.n66 B 0.029569f
C410 VDD2.n67 B 0.013246f
C411 VDD2.n68 B 0.01251f
C412 VDD2.n69 B 0.02328f
C413 VDD2.n70 B 0.02328f
C414 VDD2.n71 B 0.01251f
C415 VDD2.n72 B 0.013246f
C416 VDD2.n73 B 0.029569f
C417 VDD2.n74 B 0.029569f
C418 VDD2.n75 B 0.029569f
C419 VDD2.n76 B 0.013246f
C420 VDD2.n77 B 0.01251f
C421 VDD2.n78 B 0.02328f
C422 VDD2.n79 B 0.02328f
C423 VDD2.n80 B 0.01251f
C424 VDD2.n81 B 0.012878f
C425 VDD2.n82 B 0.012878f
C426 VDD2.n83 B 0.029569f
C427 VDD2.n84 B 0.029569f
C428 VDD2.n85 B 0.013246f
C429 VDD2.n86 B 0.01251f
C430 VDD2.n87 B 0.02328f
C431 VDD2.n88 B 0.02328f
C432 VDD2.n89 B 0.01251f
C433 VDD2.n90 B 0.013246f
C434 VDD2.n91 B 0.029569f
C435 VDD2.n92 B 0.029569f
C436 VDD2.n93 B 0.013246f
C437 VDD2.n94 B 0.01251f
C438 VDD2.n95 B 0.02328f
C439 VDD2.n96 B 0.02328f
C440 VDD2.n97 B 0.01251f
C441 VDD2.n98 B 0.013246f
C442 VDD2.n99 B 0.029569f
C443 VDD2.n100 B 0.062067f
C444 VDD2.n101 B 0.013246f
C445 VDD2.n102 B 0.01251f
C446 VDD2.n103 B 0.050313f
C447 VDD2.n104 B 0.060839f
C448 VDD2.t5 B 0.346782f
C449 VDD2.t9 B 0.346782f
C450 VDD2.n105 B 3.16164f
C451 VDD2.n106 B 0.619523f
C452 VDD2.t3 B 0.346782f
C453 VDD2.t6 B 0.346782f
C454 VDD2.n107 B 3.17592f
C455 VDD2.n108 B 2.99776f
C456 VDD2.n109 B 0.031623f
C457 VDD2.n110 B 0.02328f
C458 VDD2.n111 B 0.01251f
C459 VDD2.n112 B 0.029569f
C460 VDD2.n113 B 0.013246f
C461 VDD2.n114 B 0.02328f
C462 VDD2.n115 B 0.01251f
C463 VDD2.n116 B 0.029569f
C464 VDD2.n117 B 0.013246f
C465 VDD2.n118 B 0.02328f
C466 VDD2.n119 B 0.01251f
C467 VDD2.n120 B 0.029569f
C468 VDD2.n121 B 0.013246f
C469 VDD2.n122 B 0.02328f
C470 VDD2.n123 B 0.01251f
C471 VDD2.n124 B 0.029569f
C472 VDD2.n125 B 0.029569f
C473 VDD2.n126 B 0.013246f
C474 VDD2.n127 B 0.02328f
C475 VDD2.n128 B 0.01251f
C476 VDD2.n129 B 0.029569f
C477 VDD2.n130 B 0.013246f
C478 VDD2.n131 B 0.02328f
C479 VDD2.n132 B 0.01251f
C480 VDD2.n133 B 0.029569f
C481 VDD2.n134 B 0.013246f
C482 VDD2.n135 B 0.02328f
C483 VDD2.n136 B 0.01251f
C484 VDD2.n137 B 0.029569f
C485 VDD2.n138 B 0.013246f
C486 VDD2.n139 B 0.02328f
C487 VDD2.n140 B 0.01251f
C488 VDD2.n141 B 0.029569f
C489 VDD2.n142 B 0.013246f
C490 VDD2.n143 B 0.174312f
C491 VDD2.t2 B 0.049063f
C492 VDD2.n144 B 0.022177f
C493 VDD2.n145 B 0.017467f
C494 VDD2.n146 B 0.01251f
C495 VDD2.n147 B 1.92543f
C496 VDD2.n148 B 0.02328f
C497 VDD2.n149 B 0.01251f
C498 VDD2.n150 B 0.013246f
C499 VDD2.n151 B 0.029569f
C500 VDD2.n152 B 0.029569f
C501 VDD2.n153 B 0.013246f
C502 VDD2.n154 B 0.01251f
C503 VDD2.n155 B 0.02328f
C504 VDD2.n156 B 0.02328f
C505 VDD2.n157 B 0.01251f
C506 VDD2.n158 B 0.013246f
C507 VDD2.n159 B 0.029569f
C508 VDD2.n160 B 0.029569f
C509 VDD2.n161 B 0.013246f
C510 VDD2.n162 B 0.01251f
C511 VDD2.n163 B 0.02328f
C512 VDD2.n164 B 0.02328f
C513 VDD2.n165 B 0.01251f
C514 VDD2.n166 B 0.013246f
C515 VDD2.n167 B 0.029569f
C516 VDD2.n168 B 0.029569f
C517 VDD2.n169 B 0.013246f
C518 VDD2.n170 B 0.01251f
C519 VDD2.n171 B 0.02328f
C520 VDD2.n172 B 0.02328f
C521 VDD2.n173 B 0.01251f
C522 VDD2.n174 B 0.013246f
C523 VDD2.n175 B 0.029569f
C524 VDD2.n176 B 0.029569f
C525 VDD2.n177 B 0.013246f
C526 VDD2.n178 B 0.01251f
C527 VDD2.n179 B 0.02328f
C528 VDD2.n180 B 0.02328f
C529 VDD2.n181 B 0.01251f
C530 VDD2.n182 B 0.013246f
C531 VDD2.n183 B 0.029569f
C532 VDD2.n184 B 0.029569f
C533 VDD2.n185 B 0.013246f
C534 VDD2.n186 B 0.01251f
C535 VDD2.n187 B 0.02328f
C536 VDD2.n188 B 0.02328f
C537 VDD2.n189 B 0.01251f
C538 VDD2.n190 B 0.012878f
C539 VDD2.n191 B 0.012878f
C540 VDD2.n192 B 0.029569f
C541 VDD2.n193 B 0.029569f
C542 VDD2.n194 B 0.013246f
C543 VDD2.n195 B 0.01251f
C544 VDD2.n196 B 0.02328f
C545 VDD2.n197 B 0.02328f
C546 VDD2.n198 B 0.01251f
C547 VDD2.n199 B 0.013246f
C548 VDD2.n200 B 0.029569f
C549 VDD2.n201 B 0.029569f
C550 VDD2.n202 B 0.013246f
C551 VDD2.n203 B 0.01251f
C552 VDD2.n204 B 0.02328f
C553 VDD2.n205 B 0.02328f
C554 VDD2.n206 B 0.01251f
C555 VDD2.n207 B 0.013246f
C556 VDD2.n208 B 0.029569f
C557 VDD2.n209 B 0.062067f
C558 VDD2.n210 B 0.013246f
C559 VDD2.n211 B 0.01251f
C560 VDD2.n212 B 0.050313f
C561 VDD2.n213 B 0.050523f
C562 VDD2.n214 B 3.09248f
C563 VDD2.t7 B 0.346782f
C564 VDD2.t1 B 0.346782f
C565 VDD2.n215 B 3.16164f
C566 VDD2.n216 B 0.419899f
C567 VDD2.t8 B 0.346782f
C568 VDD2.t4 B 0.346782f
C569 VDD2.n217 B 3.17587f
C570 VTAIL.t13 B 0.349503f
C571 VTAIL.t14 B 0.349503f
C572 VTAIL.n0 B 3.10891f
C573 VTAIL.n1 B 0.50436f
C574 VTAIL.n2 B 0.031871f
C575 VTAIL.n3 B 0.023463f
C576 VTAIL.n4 B 0.012608f
C577 VTAIL.n5 B 0.029801f
C578 VTAIL.n6 B 0.01335f
C579 VTAIL.n7 B 0.023463f
C580 VTAIL.n8 B 0.012608f
C581 VTAIL.n9 B 0.029801f
C582 VTAIL.n10 B 0.01335f
C583 VTAIL.n11 B 0.023463f
C584 VTAIL.n12 B 0.012608f
C585 VTAIL.n13 B 0.029801f
C586 VTAIL.n14 B 0.01335f
C587 VTAIL.n15 B 0.023463f
C588 VTAIL.n16 B 0.012608f
C589 VTAIL.n17 B 0.029801f
C590 VTAIL.n18 B 0.01335f
C591 VTAIL.n19 B 0.023463f
C592 VTAIL.n20 B 0.012608f
C593 VTAIL.n21 B 0.029801f
C594 VTAIL.n22 B 0.01335f
C595 VTAIL.n23 B 0.023463f
C596 VTAIL.n24 B 0.012608f
C597 VTAIL.n25 B 0.029801f
C598 VTAIL.n26 B 0.01335f
C599 VTAIL.n27 B 0.023463f
C600 VTAIL.n28 B 0.012608f
C601 VTAIL.n29 B 0.029801f
C602 VTAIL.n30 B 0.01335f
C603 VTAIL.n31 B 0.023463f
C604 VTAIL.n32 B 0.012608f
C605 VTAIL.n33 B 0.029801f
C606 VTAIL.n34 B 0.01335f
C607 VTAIL.n35 B 0.17568f
C608 VTAIL.t7 B 0.049448f
C609 VTAIL.n36 B 0.022351f
C610 VTAIL.n37 B 0.017604f
C611 VTAIL.n38 B 0.012608f
C612 VTAIL.n39 B 1.94054f
C613 VTAIL.n40 B 0.023463f
C614 VTAIL.n41 B 0.012608f
C615 VTAIL.n42 B 0.01335f
C616 VTAIL.n43 B 0.029801f
C617 VTAIL.n44 B 0.029801f
C618 VTAIL.n45 B 0.01335f
C619 VTAIL.n46 B 0.012608f
C620 VTAIL.n47 B 0.023463f
C621 VTAIL.n48 B 0.023463f
C622 VTAIL.n49 B 0.012608f
C623 VTAIL.n50 B 0.01335f
C624 VTAIL.n51 B 0.029801f
C625 VTAIL.n52 B 0.029801f
C626 VTAIL.n53 B 0.01335f
C627 VTAIL.n54 B 0.012608f
C628 VTAIL.n55 B 0.023463f
C629 VTAIL.n56 B 0.023463f
C630 VTAIL.n57 B 0.012608f
C631 VTAIL.n58 B 0.01335f
C632 VTAIL.n59 B 0.029801f
C633 VTAIL.n60 B 0.029801f
C634 VTAIL.n61 B 0.01335f
C635 VTAIL.n62 B 0.012608f
C636 VTAIL.n63 B 0.023463f
C637 VTAIL.n64 B 0.023463f
C638 VTAIL.n65 B 0.012608f
C639 VTAIL.n66 B 0.01335f
C640 VTAIL.n67 B 0.029801f
C641 VTAIL.n68 B 0.029801f
C642 VTAIL.n69 B 0.01335f
C643 VTAIL.n70 B 0.012608f
C644 VTAIL.n71 B 0.023463f
C645 VTAIL.n72 B 0.023463f
C646 VTAIL.n73 B 0.012608f
C647 VTAIL.n74 B 0.01335f
C648 VTAIL.n75 B 0.029801f
C649 VTAIL.n76 B 0.029801f
C650 VTAIL.n77 B 0.029801f
C651 VTAIL.n78 B 0.01335f
C652 VTAIL.n79 B 0.012608f
C653 VTAIL.n80 B 0.023463f
C654 VTAIL.n81 B 0.023463f
C655 VTAIL.n82 B 0.012608f
C656 VTAIL.n83 B 0.012979f
C657 VTAIL.n84 B 0.012979f
C658 VTAIL.n85 B 0.029801f
C659 VTAIL.n86 B 0.029801f
C660 VTAIL.n87 B 0.01335f
C661 VTAIL.n88 B 0.012608f
C662 VTAIL.n89 B 0.023463f
C663 VTAIL.n90 B 0.023463f
C664 VTAIL.n91 B 0.012608f
C665 VTAIL.n92 B 0.01335f
C666 VTAIL.n93 B 0.029801f
C667 VTAIL.n94 B 0.029801f
C668 VTAIL.n95 B 0.01335f
C669 VTAIL.n96 B 0.012608f
C670 VTAIL.n97 B 0.023463f
C671 VTAIL.n98 B 0.023463f
C672 VTAIL.n99 B 0.012608f
C673 VTAIL.n100 B 0.01335f
C674 VTAIL.n101 B 0.029801f
C675 VTAIL.n102 B 0.062554f
C676 VTAIL.n103 B 0.01335f
C677 VTAIL.n104 B 0.012608f
C678 VTAIL.n105 B 0.050708f
C679 VTAIL.n106 B 0.034688f
C680 VTAIL.n107 B 0.317534f
C681 VTAIL.t0 B 0.349503f
C682 VTAIL.t8 B 0.349503f
C683 VTAIL.n108 B 3.10891f
C684 VTAIL.n109 B 0.59642f
C685 VTAIL.t5 B 0.349503f
C686 VTAIL.t3 B 0.349503f
C687 VTAIL.n110 B 3.10891f
C688 VTAIL.n111 B 2.31967f
C689 VTAIL.t10 B 0.349503f
C690 VTAIL.t15 B 0.349503f
C691 VTAIL.n112 B 3.10892f
C692 VTAIL.n113 B 2.31967f
C693 VTAIL.t17 B 0.349503f
C694 VTAIL.t19 B 0.349503f
C695 VTAIL.n114 B 3.10892f
C696 VTAIL.n115 B 0.596418f
C697 VTAIL.n116 B 0.031871f
C698 VTAIL.n117 B 0.023463f
C699 VTAIL.n118 B 0.012608f
C700 VTAIL.n119 B 0.029801f
C701 VTAIL.n120 B 0.01335f
C702 VTAIL.n121 B 0.023463f
C703 VTAIL.n122 B 0.012608f
C704 VTAIL.n123 B 0.029801f
C705 VTAIL.n124 B 0.01335f
C706 VTAIL.n125 B 0.023463f
C707 VTAIL.n126 B 0.012608f
C708 VTAIL.n127 B 0.029801f
C709 VTAIL.n128 B 0.01335f
C710 VTAIL.n129 B 0.023463f
C711 VTAIL.n130 B 0.012608f
C712 VTAIL.n131 B 0.029801f
C713 VTAIL.n132 B 0.029801f
C714 VTAIL.n133 B 0.01335f
C715 VTAIL.n134 B 0.023463f
C716 VTAIL.n135 B 0.012608f
C717 VTAIL.n136 B 0.029801f
C718 VTAIL.n137 B 0.01335f
C719 VTAIL.n138 B 0.023463f
C720 VTAIL.n139 B 0.012608f
C721 VTAIL.n140 B 0.029801f
C722 VTAIL.n141 B 0.01335f
C723 VTAIL.n142 B 0.023463f
C724 VTAIL.n143 B 0.012608f
C725 VTAIL.n144 B 0.029801f
C726 VTAIL.n145 B 0.01335f
C727 VTAIL.n146 B 0.023463f
C728 VTAIL.n147 B 0.012608f
C729 VTAIL.n148 B 0.029801f
C730 VTAIL.n149 B 0.01335f
C731 VTAIL.n150 B 0.17568f
C732 VTAIL.t18 B 0.049448f
C733 VTAIL.n151 B 0.022351f
C734 VTAIL.n152 B 0.017604f
C735 VTAIL.n153 B 0.012608f
C736 VTAIL.n154 B 1.94054f
C737 VTAIL.n155 B 0.023463f
C738 VTAIL.n156 B 0.012608f
C739 VTAIL.n157 B 0.01335f
C740 VTAIL.n158 B 0.029801f
C741 VTAIL.n159 B 0.029801f
C742 VTAIL.n160 B 0.01335f
C743 VTAIL.n161 B 0.012608f
C744 VTAIL.n162 B 0.023463f
C745 VTAIL.n163 B 0.023463f
C746 VTAIL.n164 B 0.012608f
C747 VTAIL.n165 B 0.01335f
C748 VTAIL.n166 B 0.029801f
C749 VTAIL.n167 B 0.029801f
C750 VTAIL.n168 B 0.01335f
C751 VTAIL.n169 B 0.012608f
C752 VTAIL.n170 B 0.023463f
C753 VTAIL.n171 B 0.023463f
C754 VTAIL.n172 B 0.012608f
C755 VTAIL.n173 B 0.01335f
C756 VTAIL.n174 B 0.029801f
C757 VTAIL.n175 B 0.029801f
C758 VTAIL.n176 B 0.01335f
C759 VTAIL.n177 B 0.012608f
C760 VTAIL.n178 B 0.023463f
C761 VTAIL.n179 B 0.023463f
C762 VTAIL.n180 B 0.012608f
C763 VTAIL.n181 B 0.01335f
C764 VTAIL.n182 B 0.029801f
C765 VTAIL.n183 B 0.029801f
C766 VTAIL.n184 B 0.01335f
C767 VTAIL.n185 B 0.012608f
C768 VTAIL.n186 B 0.023463f
C769 VTAIL.n187 B 0.023463f
C770 VTAIL.n188 B 0.012608f
C771 VTAIL.n189 B 0.01335f
C772 VTAIL.n190 B 0.029801f
C773 VTAIL.n191 B 0.029801f
C774 VTAIL.n192 B 0.01335f
C775 VTAIL.n193 B 0.012608f
C776 VTAIL.n194 B 0.023463f
C777 VTAIL.n195 B 0.023463f
C778 VTAIL.n196 B 0.012608f
C779 VTAIL.n197 B 0.012979f
C780 VTAIL.n198 B 0.012979f
C781 VTAIL.n199 B 0.029801f
C782 VTAIL.n200 B 0.029801f
C783 VTAIL.n201 B 0.01335f
C784 VTAIL.n202 B 0.012608f
C785 VTAIL.n203 B 0.023463f
C786 VTAIL.n204 B 0.023463f
C787 VTAIL.n205 B 0.012608f
C788 VTAIL.n206 B 0.01335f
C789 VTAIL.n207 B 0.029801f
C790 VTAIL.n208 B 0.029801f
C791 VTAIL.n209 B 0.01335f
C792 VTAIL.n210 B 0.012608f
C793 VTAIL.n211 B 0.023463f
C794 VTAIL.n212 B 0.023463f
C795 VTAIL.n213 B 0.012608f
C796 VTAIL.n214 B 0.01335f
C797 VTAIL.n215 B 0.029801f
C798 VTAIL.n216 B 0.062554f
C799 VTAIL.n217 B 0.01335f
C800 VTAIL.n218 B 0.012608f
C801 VTAIL.n219 B 0.050708f
C802 VTAIL.n220 B 0.034688f
C803 VTAIL.n221 B 0.317534f
C804 VTAIL.t1 B 0.349503f
C805 VTAIL.t2 B 0.349503f
C806 VTAIL.n222 B 3.10892f
C807 VTAIL.n223 B 0.543952f
C808 VTAIL.t4 B 0.349503f
C809 VTAIL.t6 B 0.349503f
C810 VTAIL.n224 B 3.10892f
C811 VTAIL.n225 B 0.596418f
C812 VTAIL.n226 B 0.031871f
C813 VTAIL.n227 B 0.023463f
C814 VTAIL.n228 B 0.012608f
C815 VTAIL.n229 B 0.029801f
C816 VTAIL.n230 B 0.01335f
C817 VTAIL.n231 B 0.023463f
C818 VTAIL.n232 B 0.012608f
C819 VTAIL.n233 B 0.029801f
C820 VTAIL.n234 B 0.01335f
C821 VTAIL.n235 B 0.023463f
C822 VTAIL.n236 B 0.012608f
C823 VTAIL.n237 B 0.029801f
C824 VTAIL.n238 B 0.01335f
C825 VTAIL.n239 B 0.023463f
C826 VTAIL.n240 B 0.012608f
C827 VTAIL.n241 B 0.029801f
C828 VTAIL.n242 B 0.029801f
C829 VTAIL.n243 B 0.01335f
C830 VTAIL.n244 B 0.023463f
C831 VTAIL.n245 B 0.012608f
C832 VTAIL.n246 B 0.029801f
C833 VTAIL.n247 B 0.01335f
C834 VTAIL.n248 B 0.023463f
C835 VTAIL.n249 B 0.012608f
C836 VTAIL.n250 B 0.029801f
C837 VTAIL.n251 B 0.01335f
C838 VTAIL.n252 B 0.023463f
C839 VTAIL.n253 B 0.012608f
C840 VTAIL.n254 B 0.029801f
C841 VTAIL.n255 B 0.01335f
C842 VTAIL.n256 B 0.023463f
C843 VTAIL.n257 B 0.012608f
C844 VTAIL.n258 B 0.029801f
C845 VTAIL.n259 B 0.01335f
C846 VTAIL.n260 B 0.17568f
C847 VTAIL.t9 B 0.049448f
C848 VTAIL.n261 B 0.022351f
C849 VTAIL.n262 B 0.017604f
C850 VTAIL.n263 B 0.012608f
C851 VTAIL.n264 B 1.94054f
C852 VTAIL.n265 B 0.023463f
C853 VTAIL.n266 B 0.012608f
C854 VTAIL.n267 B 0.01335f
C855 VTAIL.n268 B 0.029801f
C856 VTAIL.n269 B 0.029801f
C857 VTAIL.n270 B 0.01335f
C858 VTAIL.n271 B 0.012608f
C859 VTAIL.n272 B 0.023463f
C860 VTAIL.n273 B 0.023463f
C861 VTAIL.n274 B 0.012608f
C862 VTAIL.n275 B 0.01335f
C863 VTAIL.n276 B 0.029801f
C864 VTAIL.n277 B 0.029801f
C865 VTAIL.n278 B 0.01335f
C866 VTAIL.n279 B 0.012608f
C867 VTAIL.n280 B 0.023463f
C868 VTAIL.n281 B 0.023463f
C869 VTAIL.n282 B 0.012608f
C870 VTAIL.n283 B 0.01335f
C871 VTAIL.n284 B 0.029801f
C872 VTAIL.n285 B 0.029801f
C873 VTAIL.n286 B 0.01335f
C874 VTAIL.n287 B 0.012608f
C875 VTAIL.n288 B 0.023463f
C876 VTAIL.n289 B 0.023463f
C877 VTAIL.n290 B 0.012608f
C878 VTAIL.n291 B 0.01335f
C879 VTAIL.n292 B 0.029801f
C880 VTAIL.n293 B 0.029801f
C881 VTAIL.n294 B 0.01335f
C882 VTAIL.n295 B 0.012608f
C883 VTAIL.n296 B 0.023463f
C884 VTAIL.n297 B 0.023463f
C885 VTAIL.n298 B 0.012608f
C886 VTAIL.n299 B 0.01335f
C887 VTAIL.n300 B 0.029801f
C888 VTAIL.n301 B 0.029801f
C889 VTAIL.n302 B 0.01335f
C890 VTAIL.n303 B 0.012608f
C891 VTAIL.n304 B 0.023463f
C892 VTAIL.n305 B 0.023463f
C893 VTAIL.n306 B 0.012608f
C894 VTAIL.n307 B 0.012979f
C895 VTAIL.n308 B 0.012979f
C896 VTAIL.n309 B 0.029801f
C897 VTAIL.n310 B 0.029801f
C898 VTAIL.n311 B 0.01335f
C899 VTAIL.n312 B 0.012608f
C900 VTAIL.n313 B 0.023463f
C901 VTAIL.n314 B 0.023463f
C902 VTAIL.n315 B 0.012608f
C903 VTAIL.n316 B 0.01335f
C904 VTAIL.n317 B 0.029801f
C905 VTAIL.n318 B 0.029801f
C906 VTAIL.n319 B 0.01335f
C907 VTAIL.n320 B 0.012608f
C908 VTAIL.n321 B 0.023463f
C909 VTAIL.n322 B 0.023463f
C910 VTAIL.n323 B 0.012608f
C911 VTAIL.n324 B 0.01335f
C912 VTAIL.n325 B 0.029801f
C913 VTAIL.n326 B 0.062554f
C914 VTAIL.n327 B 0.01335f
C915 VTAIL.n328 B 0.012608f
C916 VTAIL.n329 B 0.050708f
C917 VTAIL.n330 B 0.034688f
C918 VTAIL.n331 B 1.91727f
C919 VTAIL.n332 B 0.031871f
C920 VTAIL.n333 B 0.023463f
C921 VTAIL.n334 B 0.012608f
C922 VTAIL.n335 B 0.029801f
C923 VTAIL.n336 B 0.01335f
C924 VTAIL.n337 B 0.023463f
C925 VTAIL.n338 B 0.012608f
C926 VTAIL.n339 B 0.029801f
C927 VTAIL.n340 B 0.01335f
C928 VTAIL.n341 B 0.023463f
C929 VTAIL.n342 B 0.012608f
C930 VTAIL.n343 B 0.029801f
C931 VTAIL.n344 B 0.01335f
C932 VTAIL.n345 B 0.023463f
C933 VTAIL.n346 B 0.012608f
C934 VTAIL.n347 B 0.029801f
C935 VTAIL.n348 B 0.01335f
C936 VTAIL.n349 B 0.023463f
C937 VTAIL.n350 B 0.012608f
C938 VTAIL.n351 B 0.029801f
C939 VTAIL.n352 B 0.01335f
C940 VTAIL.n353 B 0.023463f
C941 VTAIL.n354 B 0.012608f
C942 VTAIL.n355 B 0.029801f
C943 VTAIL.n356 B 0.01335f
C944 VTAIL.n357 B 0.023463f
C945 VTAIL.n358 B 0.012608f
C946 VTAIL.n359 B 0.029801f
C947 VTAIL.n360 B 0.01335f
C948 VTAIL.n361 B 0.023463f
C949 VTAIL.n362 B 0.012608f
C950 VTAIL.n363 B 0.029801f
C951 VTAIL.n364 B 0.01335f
C952 VTAIL.n365 B 0.17568f
C953 VTAIL.t11 B 0.049448f
C954 VTAIL.n366 B 0.022351f
C955 VTAIL.n367 B 0.017604f
C956 VTAIL.n368 B 0.012608f
C957 VTAIL.n369 B 1.94054f
C958 VTAIL.n370 B 0.023463f
C959 VTAIL.n371 B 0.012608f
C960 VTAIL.n372 B 0.01335f
C961 VTAIL.n373 B 0.029801f
C962 VTAIL.n374 B 0.029801f
C963 VTAIL.n375 B 0.01335f
C964 VTAIL.n376 B 0.012608f
C965 VTAIL.n377 B 0.023463f
C966 VTAIL.n378 B 0.023463f
C967 VTAIL.n379 B 0.012608f
C968 VTAIL.n380 B 0.01335f
C969 VTAIL.n381 B 0.029801f
C970 VTAIL.n382 B 0.029801f
C971 VTAIL.n383 B 0.01335f
C972 VTAIL.n384 B 0.012608f
C973 VTAIL.n385 B 0.023463f
C974 VTAIL.n386 B 0.023463f
C975 VTAIL.n387 B 0.012608f
C976 VTAIL.n388 B 0.01335f
C977 VTAIL.n389 B 0.029801f
C978 VTAIL.n390 B 0.029801f
C979 VTAIL.n391 B 0.01335f
C980 VTAIL.n392 B 0.012608f
C981 VTAIL.n393 B 0.023463f
C982 VTAIL.n394 B 0.023463f
C983 VTAIL.n395 B 0.012608f
C984 VTAIL.n396 B 0.01335f
C985 VTAIL.n397 B 0.029801f
C986 VTAIL.n398 B 0.029801f
C987 VTAIL.n399 B 0.01335f
C988 VTAIL.n400 B 0.012608f
C989 VTAIL.n401 B 0.023463f
C990 VTAIL.n402 B 0.023463f
C991 VTAIL.n403 B 0.012608f
C992 VTAIL.n404 B 0.01335f
C993 VTAIL.n405 B 0.029801f
C994 VTAIL.n406 B 0.029801f
C995 VTAIL.n407 B 0.029801f
C996 VTAIL.n408 B 0.01335f
C997 VTAIL.n409 B 0.012608f
C998 VTAIL.n410 B 0.023463f
C999 VTAIL.n411 B 0.023463f
C1000 VTAIL.n412 B 0.012608f
C1001 VTAIL.n413 B 0.012979f
C1002 VTAIL.n414 B 0.012979f
C1003 VTAIL.n415 B 0.029801f
C1004 VTAIL.n416 B 0.029801f
C1005 VTAIL.n417 B 0.01335f
C1006 VTAIL.n418 B 0.012608f
C1007 VTAIL.n419 B 0.023463f
C1008 VTAIL.n420 B 0.023463f
C1009 VTAIL.n421 B 0.012608f
C1010 VTAIL.n422 B 0.01335f
C1011 VTAIL.n423 B 0.029801f
C1012 VTAIL.n424 B 0.029801f
C1013 VTAIL.n425 B 0.01335f
C1014 VTAIL.n426 B 0.012608f
C1015 VTAIL.n427 B 0.023463f
C1016 VTAIL.n428 B 0.023463f
C1017 VTAIL.n429 B 0.012608f
C1018 VTAIL.n430 B 0.01335f
C1019 VTAIL.n431 B 0.029801f
C1020 VTAIL.n432 B 0.062554f
C1021 VTAIL.n433 B 0.01335f
C1022 VTAIL.n434 B 0.012608f
C1023 VTAIL.n435 B 0.050708f
C1024 VTAIL.n436 B 0.034688f
C1025 VTAIL.n437 B 1.91727f
C1026 VTAIL.t16 B 0.349503f
C1027 VTAIL.t12 B 0.349503f
C1028 VTAIL.n438 B 3.10891f
C1029 VTAIL.n439 B 0.460041f
C1030 VN.n0 B 0.028673f
C1031 VN.t3 B 2.6747f
C1032 VN.n1 B 0.028718f
C1033 VN.n2 B 0.021748f
C1034 VN.t6 B 2.6747f
C1035 VN.n3 B 0.927627f
C1036 VN.n4 B 0.021748f
C1037 VN.n5 B 0.043569f
C1038 VN.n6 B 0.021748f
C1039 VN.t0 B 2.6747f
C1040 VN.n7 B 0.020545f
C1041 VN.n8 B 0.204932f
C1042 VN.t4 B 2.6747f
C1043 VN.t9 B 2.8286f
C1044 VN.n9 B 0.973849f
C1045 VN.n10 B 0.996066f
C1046 VN.n11 B 0.038532f
C1047 VN.n12 B 0.039916f
C1048 VN.n13 B 0.021748f
C1049 VN.n14 B 0.021748f
C1050 VN.n15 B 0.021748f
C1051 VN.n16 B 0.043569f
C1052 VN.n17 B 0.030527f
C1053 VN.n18 B 0.927627f
C1054 VN.n19 B 0.030527f
C1055 VN.n20 B 0.021748f
C1056 VN.n21 B 0.021748f
C1057 VN.n22 B 0.021748f
C1058 VN.n23 B 0.020545f
C1059 VN.n24 B 0.039916f
C1060 VN.n25 B 0.038532f
C1061 VN.n26 B 0.021748f
C1062 VN.n27 B 0.021748f
C1063 VN.n28 B 0.022523f
C1064 VN.n29 B 0.040533f
C1065 VN.n30 B 0.034779f
C1066 VN.n31 B 0.021748f
C1067 VN.n32 B 0.021748f
C1068 VN.n33 B 0.021748f
C1069 VN.n34 B 0.040533f
C1070 VN.n35 B 0.026525f
C1071 VN.n36 B 0.990734f
C1072 VN.n37 B 0.035068f
C1073 VN.n38 B 0.028673f
C1074 VN.t7 B 2.6747f
C1075 VN.n39 B 0.028718f
C1076 VN.n40 B 0.021748f
C1077 VN.t2 B 2.6747f
C1078 VN.n41 B 0.927627f
C1079 VN.n42 B 0.021748f
C1080 VN.n43 B 0.043569f
C1081 VN.n44 B 0.021748f
C1082 VN.t8 B 2.6747f
C1083 VN.n45 B 0.020545f
C1084 VN.n46 B 0.204932f
C1085 VN.t1 B 2.6747f
C1086 VN.t5 B 2.8286f
C1087 VN.n47 B 0.973849f
C1088 VN.n48 B 0.996066f
C1089 VN.n49 B 0.038532f
C1090 VN.n50 B 0.039916f
C1091 VN.n51 B 0.021748f
C1092 VN.n52 B 0.021748f
C1093 VN.n53 B 0.021748f
C1094 VN.n54 B 0.043569f
C1095 VN.n55 B 0.030527f
C1096 VN.n56 B 0.927627f
C1097 VN.n57 B 0.030527f
C1098 VN.n58 B 0.021748f
C1099 VN.n59 B 0.021748f
C1100 VN.n60 B 0.021748f
C1101 VN.n61 B 0.020545f
C1102 VN.n62 B 0.039916f
C1103 VN.n63 B 0.038532f
C1104 VN.n64 B 0.021748f
C1105 VN.n65 B 0.021748f
C1106 VN.n66 B 0.022523f
C1107 VN.n67 B 0.040533f
C1108 VN.n68 B 0.034779f
C1109 VN.n69 B 0.021748f
C1110 VN.n70 B 0.021748f
C1111 VN.n71 B 0.021748f
C1112 VN.n72 B 0.040533f
C1113 VN.n73 B 0.026525f
C1114 VN.n74 B 0.990734f
C1115 VN.n75 B 1.46815f
.ends

