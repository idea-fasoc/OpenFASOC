* NGSPICE file created from diff_pair_sample_1076.ext - technology: sky130A

.subckt diff_pair_sample_1076 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t0 w_n2110_n4366# sky130_fd_pr__pfet_01v8 ad=6.6261 pd=34.76 as=2.80335 ps=17.32 w=16.99 l=1.57
X1 VDD1.t3 VP.t1 VTAIL.t6 w_n2110_n4366# sky130_fd_pr__pfet_01v8 ad=2.80335 pd=17.32 as=6.6261 ps=34.76 w=16.99 l=1.57
X2 VDD2.t3 VN.t0 VTAIL.t2 w_n2110_n4366# sky130_fd_pr__pfet_01v8 ad=2.80335 pd=17.32 as=6.6261 ps=34.76 w=16.99 l=1.57
X3 VTAIL.t1 VN.t1 VDD2.t2 w_n2110_n4366# sky130_fd_pr__pfet_01v8 ad=6.6261 pd=34.76 as=2.80335 ps=17.32 w=16.99 l=1.57
X4 B.t11 B.t9 B.t10 w_n2110_n4366# sky130_fd_pr__pfet_01v8 ad=6.6261 pd=34.76 as=0 ps=0 w=16.99 l=1.57
X5 B.t8 B.t6 B.t7 w_n2110_n4366# sky130_fd_pr__pfet_01v8 ad=6.6261 pd=34.76 as=0 ps=0 w=16.99 l=1.57
X6 VDD2.t1 VN.t2 VTAIL.t3 w_n2110_n4366# sky130_fd_pr__pfet_01v8 ad=2.80335 pd=17.32 as=6.6261 ps=34.76 w=16.99 l=1.57
X7 VTAIL.t0 VN.t3 VDD2.t0 w_n2110_n4366# sky130_fd_pr__pfet_01v8 ad=6.6261 pd=34.76 as=2.80335 ps=17.32 w=16.99 l=1.57
X8 VTAIL.t5 VP.t2 VDD1.t1 w_n2110_n4366# sky130_fd_pr__pfet_01v8 ad=6.6261 pd=34.76 as=2.80335 ps=17.32 w=16.99 l=1.57
X9 VDD1.t2 VP.t3 VTAIL.t4 w_n2110_n4366# sky130_fd_pr__pfet_01v8 ad=2.80335 pd=17.32 as=6.6261 ps=34.76 w=16.99 l=1.57
X10 B.t5 B.t3 B.t4 w_n2110_n4366# sky130_fd_pr__pfet_01v8 ad=6.6261 pd=34.76 as=0 ps=0 w=16.99 l=1.57
X11 B.t2 B.t0 B.t1 w_n2110_n4366# sky130_fd_pr__pfet_01v8 ad=6.6261 pd=34.76 as=0 ps=0 w=16.99 l=1.57
R0 VP.n2 VP.t2 298.171
R1 VP.n2 VP.t1 297.848
R2 VP.n4 VP.t0 260.803
R3 VP.n11 VP.t3 260.803
R4 VP.n4 VP.n3 175.981
R5 VP.n12 VP.n11 175.981
R6 VP.n10 VP.n0 161.3
R7 VP.n9 VP.n8 161.3
R8 VP.n7 VP.n1 161.3
R9 VP.n6 VP.n5 161.3
R10 VP.n3 VP.n2 59.6833
R11 VP.n9 VP.n1 56.5193
R12 VP.n5 VP.n1 24.4675
R13 VP.n10 VP.n9 24.4675
R14 VP.n5 VP.n4 9.7873
R15 VP.n11 VP.n10 9.7873
R16 VP.n6 VP.n3 0.189894
R17 VP.n7 VP.n6 0.189894
R18 VP.n8 VP.n7 0.189894
R19 VP.n8 VP.n0 0.189894
R20 VP.n12 VP.n0 0.189894
R21 VP VP.n12 0.0516364
R22 VDD1 VDD1.n1 116.876
R23 VDD1 VDD1.n0 73.1349
R24 VDD1.n0 VDD1.t1 1.91368
R25 VDD1.n0 VDD1.t3 1.91368
R26 VDD1.n1 VDD1.t0 1.91368
R27 VDD1.n1 VDD1.t2 1.91368
R28 VTAIL.n746 VTAIL.n658 756.745
R29 VTAIL.n88 VTAIL.n0 756.745
R30 VTAIL.n182 VTAIL.n94 756.745
R31 VTAIL.n276 VTAIL.n188 756.745
R32 VTAIL.n652 VTAIL.n564 756.745
R33 VTAIL.n558 VTAIL.n470 756.745
R34 VTAIL.n464 VTAIL.n376 756.745
R35 VTAIL.n370 VTAIL.n282 756.745
R36 VTAIL.n689 VTAIL.n688 585
R37 VTAIL.n686 VTAIL.n685 585
R38 VTAIL.n695 VTAIL.n694 585
R39 VTAIL.n697 VTAIL.n696 585
R40 VTAIL.n682 VTAIL.n681 585
R41 VTAIL.n703 VTAIL.n702 585
R42 VTAIL.n705 VTAIL.n704 585
R43 VTAIL.n678 VTAIL.n677 585
R44 VTAIL.n711 VTAIL.n710 585
R45 VTAIL.n713 VTAIL.n712 585
R46 VTAIL.n674 VTAIL.n673 585
R47 VTAIL.n719 VTAIL.n718 585
R48 VTAIL.n721 VTAIL.n720 585
R49 VTAIL.n670 VTAIL.n669 585
R50 VTAIL.n727 VTAIL.n726 585
R51 VTAIL.n730 VTAIL.n729 585
R52 VTAIL.n728 VTAIL.n666 585
R53 VTAIL.n735 VTAIL.n665 585
R54 VTAIL.n737 VTAIL.n736 585
R55 VTAIL.n739 VTAIL.n738 585
R56 VTAIL.n662 VTAIL.n661 585
R57 VTAIL.n745 VTAIL.n744 585
R58 VTAIL.n747 VTAIL.n746 585
R59 VTAIL.n31 VTAIL.n30 585
R60 VTAIL.n28 VTAIL.n27 585
R61 VTAIL.n37 VTAIL.n36 585
R62 VTAIL.n39 VTAIL.n38 585
R63 VTAIL.n24 VTAIL.n23 585
R64 VTAIL.n45 VTAIL.n44 585
R65 VTAIL.n47 VTAIL.n46 585
R66 VTAIL.n20 VTAIL.n19 585
R67 VTAIL.n53 VTAIL.n52 585
R68 VTAIL.n55 VTAIL.n54 585
R69 VTAIL.n16 VTAIL.n15 585
R70 VTAIL.n61 VTAIL.n60 585
R71 VTAIL.n63 VTAIL.n62 585
R72 VTAIL.n12 VTAIL.n11 585
R73 VTAIL.n69 VTAIL.n68 585
R74 VTAIL.n72 VTAIL.n71 585
R75 VTAIL.n70 VTAIL.n8 585
R76 VTAIL.n77 VTAIL.n7 585
R77 VTAIL.n79 VTAIL.n78 585
R78 VTAIL.n81 VTAIL.n80 585
R79 VTAIL.n4 VTAIL.n3 585
R80 VTAIL.n87 VTAIL.n86 585
R81 VTAIL.n89 VTAIL.n88 585
R82 VTAIL.n125 VTAIL.n124 585
R83 VTAIL.n122 VTAIL.n121 585
R84 VTAIL.n131 VTAIL.n130 585
R85 VTAIL.n133 VTAIL.n132 585
R86 VTAIL.n118 VTAIL.n117 585
R87 VTAIL.n139 VTAIL.n138 585
R88 VTAIL.n141 VTAIL.n140 585
R89 VTAIL.n114 VTAIL.n113 585
R90 VTAIL.n147 VTAIL.n146 585
R91 VTAIL.n149 VTAIL.n148 585
R92 VTAIL.n110 VTAIL.n109 585
R93 VTAIL.n155 VTAIL.n154 585
R94 VTAIL.n157 VTAIL.n156 585
R95 VTAIL.n106 VTAIL.n105 585
R96 VTAIL.n163 VTAIL.n162 585
R97 VTAIL.n166 VTAIL.n165 585
R98 VTAIL.n164 VTAIL.n102 585
R99 VTAIL.n171 VTAIL.n101 585
R100 VTAIL.n173 VTAIL.n172 585
R101 VTAIL.n175 VTAIL.n174 585
R102 VTAIL.n98 VTAIL.n97 585
R103 VTAIL.n181 VTAIL.n180 585
R104 VTAIL.n183 VTAIL.n182 585
R105 VTAIL.n219 VTAIL.n218 585
R106 VTAIL.n216 VTAIL.n215 585
R107 VTAIL.n225 VTAIL.n224 585
R108 VTAIL.n227 VTAIL.n226 585
R109 VTAIL.n212 VTAIL.n211 585
R110 VTAIL.n233 VTAIL.n232 585
R111 VTAIL.n235 VTAIL.n234 585
R112 VTAIL.n208 VTAIL.n207 585
R113 VTAIL.n241 VTAIL.n240 585
R114 VTAIL.n243 VTAIL.n242 585
R115 VTAIL.n204 VTAIL.n203 585
R116 VTAIL.n249 VTAIL.n248 585
R117 VTAIL.n251 VTAIL.n250 585
R118 VTAIL.n200 VTAIL.n199 585
R119 VTAIL.n257 VTAIL.n256 585
R120 VTAIL.n260 VTAIL.n259 585
R121 VTAIL.n258 VTAIL.n196 585
R122 VTAIL.n265 VTAIL.n195 585
R123 VTAIL.n267 VTAIL.n266 585
R124 VTAIL.n269 VTAIL.n268 585
R125 VTAIL.n192 VTAIL.n191 585
R126 VTAIL.n275 VTAIL.n274 585
R127 VTAIL.n277 VTAIL.n276 585
R128 VTAIL.n653 VTAIL.n652 585
R129 VTAIL.n651 VTAIL.n650 585
R130 VTAIL.n568 VTAIL.n567 585
R131 VTAIL.n645 VTAIL.n644 585
R132 VTAIL.n643 VTAIL.n642 585
R133 VTAIL.n641 VTAIL.n571 585
R134 VTAIL.n575 VTAIL.n572 585
R135 VTAIL.n636 VTAIL.n635 585
R136 VTAIL.n634 VTAIL.n633 585
R137 VTAIL.n577 VTAIL.n576 585
R138 VTAIL.n628 VTAIL.n627 585
R139 VTAIL.n626 VTAIL.n625 585
R140 VTAIL.n581 VTAIL.n580 585
R141 VTAIL.n620 VTAIL.n619 585
R142 VTAIL.n618 VTAIL.n617 585
R143 VTAIL.n585 VTAIL.n584 585
R144 VTAIL.n612 VTAIL.n611 585
R145 VTAIL.n610 VTAIL.n609 585
R146 VTAIL.n589 VTAIL.n588 585
R147 VTAIL.n604 VTAIL.n603 585
R148 VTAIL.n602 VTAIL.n601 585
R149 VTAIL.n593 VTAIL.n592 585
R150 VTAIL.n596 VTAIL.n595 585
R151 VTAIL.n559 VTAIL.n558 585
R152 VTAIL.n557 VTAIL.n556 585
R153 VTAIL.n474 VTAIL.n473 585
R154 VTAIL.n551 VTAIL.n550 585
R155 VTAIL.n549 VTAIL.n548 585
R156 VTAIL.n547 VTAIL.n477 585
R157 VTAIL.n481 VTAIL.n478 585
R158 VTAIL.n542 VTAIL.n541 585
R159 VTAIL.n540 VTAIL.n539 585
R160 VTAIL.n483 VTAIL.n482 585
R161 VTAIL.n534 VTAIL.n533 585
R162 VTAIL.n532 VTAIL.n531 585
R163 VTAIL.n487 VTAIL.n486 585
R164 VTAIL.n526 VTAIL.n525 585
R165 VTAIL.n524 VTAIL.n523 585
R166 VTAIL.n491 VTAIL.n490 585
R167 VTAIL.n518 VTAIL.n517 585
R168 VTAIL.n516 VTAIL.n515 585
R169 VTAIL.n495 VTAIL.n494 585
R170 VTAIL.n510 VTAIL.n509 585
R171 VTAIL.n508 VTAIL.n507 585
R172 VTAIL.n499 VTAIL.n498 585
R173 VTAIL.n502 VTAIL.n501 585
R174 VTAIL.n465 VTAIL.n464 585
R175 VTAIL.n463 VTAIL.n462 585
R176 VTAIL.n380 VTAIL.n379 585
R177 VTAIL.n457 VTAIL.n456 585
R178 VTAIL.n455 VTAIL.n454 585
R179 VTAIL.n453 VTAIL.n383 585
R180 VTAIL.n387 VTAIL.n384 585
R181 VTAIL.n448 VTAIL.n447 585
R182 VTAIL.n446 VTAIL.n445 585
R183 VTAIL.n389 VTAIL.n388 585
R184 VTAIL.n440 VTAIL.n439 585
R185 VTAIL.n438 VTAIL.n437 585
R186 VTAIL.n393 VTAIL.n392 585
R187 VTAIL.n432 VTAIL.n431 585
R188 VTAIL.n430 VTAIL.n429 585
R189 VTAIL.n397 VTAIL.n396 585
R190 VTAIL.n424 VTAIL.n423 585
R191 VTAIL.n422 VTAIL.n421 585
R192 VTAIL.n401 VTAIL.n400 585
R193 VTAIL.n416 VTAIL.n415 585
R194 VTAIL.n414 VTAIL.n413 585
R195 VTAIL.n405 VTAIL.n404 585
R196 VTAIL.n408 VTAIL.n407 585
R197 VTAIL.n371 VTAIL.n370 585
R198 VTAIL.n369 VTAIL.n368 585
R199 VTAIL.n286 VTAIL.n285 585
R200 VTAIL.n363 VTAIL.n362 585
R201 VTAIL.n361 VTAIL.n360 585
R202 VTAIL.n359 VTAIL.n289 585
R203 VTAIL.n293 VTAIL.n290 585
R204 VTAIL.n354 VTAIL.n353 585
R205 VTAIL.n352 VTAIL.n351 585
R206 VTAIL.n295 VTAIL.n294 585
R207 VTAIL.n346 VTAIL.n345 585
R208 VTAIL.n344 VTAIL.n343 585
R209 VTAIL.n299 VTAIL.n298 585
R210 VTAIL.n338 VTAIL.n337 585
R211 VTAIL.n336 VTAIL.n335 585
R212 VTAIL.n303 VTAIL.n302 585
R213 VTAIL.n330 VTAIL.n329 585
R214 VTAIL.n328 VTAIL.n327 585
R215 VTAIL.n307 VTAIL.n306 585
R216 VTAIL.n322 VTAIL.n321 585
R217 VTAIL.n320 VTAIL.n319 585
R218 VTAIL.n311 VTAIL.n310 585
R219 VTAIL.n314 VTAIL.n313 585
R220 VTAIL.t6 VTAIL.n594 327.466
R221 VTAIL.t5 VTAIL.n500 327.466
R222 VTAIL.t2 VTAIL.n406 327.466
R223 VTAIL.t0 VTAIL.n312 327.466
R224 VTAIL.t3 VTAIL.n687 327.466
R225 VTAIL.t1 VTAIL.n29 327.466
R226 VTAIL.t4 VTAIL.n123 327.466
R227 VTAIL.t7 VTAIL.n217 327.466
R228 VTAIL.n688 VTAIL.n685 171.744
R229 VTAIL.n695 VTAIL.n685 171.744
R230 VTAIL.n696 VTAIL.n695 171.744
R231 VTAIL.n696 VTAIL.n681 171.744
R232 VTAIL.n703 VTAIL.n681 171.744
R233 VTAIL.n704 VTAIL.n703 171.744
R234 VTAIL.n704 VTAIL.n677 171.744
R235 VTAIL.n711 VTAIL.n677 171.744
R236 VTAIL.n712 VTAIL.n711 171.744
R237 VTAIL.n712 VTAIL.n673 171.744
R238 VTAIL.n719 VTAIL.n673 171.744
R239 VTAIL.n720 VTAIL.n719 171.744
R240 VTAIL.n720 VTAIL.n669 171.744
R241 VTAIL.n727 VTAIL.n669 171.744
R242 VTAIL.n729 VTAIL.n727 171.744
R243 VTAIL.n729 VTAIL.n728 171.744
R244 VTAIL.n728 VTAIL.n665 171.744
R245 VTAIL.n737 VTAIL.n665 171.744
R246 VTAIL.n738 VTAIL.n737 171.744
R247 VTAIL.n738 VTAIL.n661 171.744
R248 VTAIL.n745 VTAIL.n661 171.744
R249 VTAIL.n746 VTAIL.n745 171.744
R250 VTAIL.n30 VTAIL.n27 171.744
R251 VTAIL.n37 VTAIL.n27 171.744
R252 VTAIL.n38 VTAIL.n37 171.744
R253 VTAIL.n38 VTAIL.n23 171.744
R254 VTAIL.n45 VTAIL.n23 171.744
R255 VTAIL.n46 VTAIL.n45 171.744
R256 VTAIL.n46 VTAIL.n19 171.744
R257 VTAIL.n53 VTAIL.n19 171.744
R258 VTAIL.n54 VTAIL.n53 171.744
R259 VTAIL.n54 VTAIL.n15 171.744
R260 VTAIL.n61 VTAIL.n15 171.744
R261 VTAIL.n62 VTAIL.n61 171.744
R262 VTAIL.n62 VTAIL.n11 171.744
R263 VTAIL.n69 VTAIL.n11 171.744
R264 VTAIL.n71 VTAIL.n69 171.744
R265 VTAIL.n71 VTAIL.n70 171.744
R266 VTAIL.n70 VTAIL.n7 171.744
R267 VTAIL.n79 VTAIL.n7 171.744
R268 VTAIL.n80 VTAIL.n79 171.744
R269 VTAIL.n80 VTAIL.n3 171.744
R270 VTAIL.n87 VTAIL.n3 171.744
R271 VTAIL.n88 VTAIL.n87 171.744
R272 VTAIL.n124 VTAIL.n121 171.744
R273 VTAIL.n131 VTAIL.n121 171.744
R274 VTAIL.n132 VTAIL.n131 171.744
R275 VTAIL.n132 VTAIL.n117 171.744
R276 VTAIL.n139 VTAIL.n117 171.744
R277 VTAIL.n140 VTAIL.n139 171.744
R278 VTAIL.n140 VTAIL.n113 171.744
R279 VTAIL.n147 VTAIL.n113 171.744
R280 VTAIL.n148 VTAIL.n147 171.744
R281 VTAIL.n148 VTAIL.n109 171.744
R282 VTAIL.n155 VTAIL.n109 171.744
R283 VTAIL.n156 VTAIL.n155 171.744
R284 VTAIL.n156 VTAIL.n105 171.744
R285 VTAIL.n163 VTAIL.n105 171.744
R286 VTAIL.n165 VTAIL.n163 171.744
R287 VTAIL.n165 VTAIL.n164 171.744
R288 VTAIL.n164 VTAIL.n101 171.744
R289 VTAIL.n173 VTAIL.n101 171.744
R290 VTAIL.n174 VTAIL.n173 171.744
R291 VTAIL.n174 VTAIL.n97 171.744
R292 VTAIL.n181 VTAIL.n97 171.744
R293 VTAIL.n182 VTAIL.n181 171.744
R294 VTAIL.n218 VTAIL.n215 171.744
R295 VTAIL.n225 VTAIL.n215 171.744
R296 VTAIL.n226 VTAIL.n225 171.744
R297 VTAIL.n226 VTAIL.n211 171.744
R298 VTAIL.n233 VTAIL.n211 171.744
R299 VTAIL.n234 VTAIL.n233 171.744
R300 VTAIL.n234 VTAIL.n207 171.744
R301 VTAIL.n241 VTAIL.n207 171.744
R302 VTAIL.n242 VTAIL.n241 171.744
R303 VTAIL.n242 VTAIL.n203 171.744
R304 VTAIL.n249 VTAIL.n203 171.744
R305 VTAIL.n250 VTAIL.n249 171.744
R306 VTAIL.n250 VTAIL.n199 171.744
R307 VTAIL.n257 VTAIL.n199 171.744
R308 VTAIL.n259 VTAIL.n257 171.744
R309 VTAIL.n259 VTAIL.n258 171.744
R310 VTAIL.n258 VTAIL.n195 171.744
R311 VTAIL.n267 VTAIL.n195 171.744
R312 VTAIL.n268 VTAIL.n267 171.744
R313 VTAIL.n268 VTAIL.n191 171.744
R314 VTAIL.n275 VTAIL.n191 171.744
R315 VTAIL.n276 VTAIL.n275 171.744
R316 VTAIL.n652 VTAIL.n651 171.744
R317 VTAIL.n651 VTAIL.n567 171.744
R318 VTAIL.n644 VTAIL.n567 171.744
R319 VTAIL.n644 VTAIL.n643 171.744
R320 VTAIL.n643 VTAIL.n571 171.744
R321 VTAIL.n575 VTAIL.n571 171.744
R322 VTAIL.n635 VTAIL.n575 171.744
R323 VTAIL.n635 VTAIL.n634 171.744
R324 VTAIL.n634 VTAIL.n576 171.744
R325 VTAIL.n627 VTAIL.n576 171.744
R326 VTAIL.n627 VTAIL.n626 171.744
R327 VTAIL.n626 VTAIL.n580 171.744
R328 VTAIL.n619 VTAIL.n580 171.744
R329 VTAIL.n619 VTAIL.n618 171.744
R330 VTAIL.n618 VTAIL.n584 171.744
R331 VTAIL.n611 VTAIL.n584 171.744
R332 VTAIL.n611 VTAIL.n610 171.744
R333 VTAIL.n610 VTAIL.n588 171.744
R334 VTAIL.n603 VTAIL.n588 171.744
R335 VTAIL.n603 VTAIL.n602 171.744
R336 VTAIL.n602 VTAIL.n592 171.744
R337 VTAIL.n595 VTAIL.n592 171.744
R338 VTAIL.n558 VTAIL.n557 171.744
R339 VTAIL.n557 VTAIL.n473 171.744
R340 VTAIL.n550 VTAIL.n473 171.744
R341 VTAIL.n550 VTAIL.n549 171.744
R342 VTAIL.n549 VTAIL.n477 171.744
R343 VTAIL.n481 VTAIL.n477 171.744
R344 VTAIL.n541 VTAIL.n481 171.744
R345 VTAIL.n541 VTAIL.n540 171.744
R346 VTAIL.n540 VTAIL.n482 171.744
R347 VTAIL.n533 VTAIL.n482 171.744
R348 VTAIL.n533 VTAIL.n532 171.744
R349 VTAIL.n532 VTAIL.n486 171.744
R350 VTAIL.n525 VTAIL.n486 171.744
R351 VTAIL.n525 VTAIL.n524 171.744
R352 VTAIL.n524 VTAIL.n490 171.744
R353 VTAIL.n517 VTAIL.n490 171.744
R354 VTAIL.n517 VTAIL.n516 171.744
R355 VTAIL.n516 VTAIL.n494 171.744
R356 VTAIL.n509 VTAIL.n494 171.744
R357 VTAIL.n509 VTAIL.n508 171.744
R358 VTAIL.n508 VTAIL.n498 171.744
R359 VTAIL.n501 VTAIL.n498 171.744
R360 VTAIL.n464 VTAIL.n463 171.744
R361 VTAIL.n463 VTAIL.n379 171.744
R362 VTAIL.n456 VTAIL.n379 171.744
R363 VTAIL.n456 VTAIL.n455 171.744
R364 VTAIL.n455 VTAIL.n383 171.744
R365 VTAIL.n387 VTAIL.n383 171.744
R366 VTAIL.n447 VTAIL.n387 171.744
R367 VTAIL.n447 VTAIL.n446 171.744
R368 VTAIL.n446 VTAIL.n388 171.744
R369 VTAIL.n439 VTAIL.n388 171.744
R370 VTAIL.n439 VTAIL.n438 171.744
R371 VTAIL.n438 VTAIL.n392 171.744
R372 VTAIL.n431 VTAIL.n392 171.744
R373 VTAIL.n431 VTAIL.n430 171.744
R374 VTAIL.n430 VTAIL.n396 171.744
R375 VTAIL.n423 VTAIL.n396 171.744
R376 VTAIL.n423 VTAIL.n422 171.744
R377 VTAIL.n422 VTAIL.n400 171.744
R378 VTAIL.n415 VTAIL.n400 171.744
R379 VTAIL.n415 VTAIL.n414 171.744
R380 VTAIL.n414 VTAIL.n404 171.744
R381 VTAIL.n407 VTAIL.n404 171.744
R382 VTAIL.n370 VTAIL.n369 171.744
R383 VTAIL.n369 VTAIL.n285 171.744
R384 VTAIL.n362 VTAIL.n285 171.744
R385 VTAIL.n362 VTAIL.n361 171.744
R386 VTAIL.n361 VTAIL.n289 171.744
R387 VTAIL.n293 VTAIL.n289 171.744
R388 VTAIL.n353 VTAIL.n293 171.744
R389 VTAIL.n353 VTAIL.n352 171.744
R390 VTAIL.n352 VTAIL.n294 171.744
R391 VTAIL.n345 VTAIL.n294 171.744
R392 VTAIL.n345 VTAIL.n344 171.744
R393 VTAIL.n344 VTAIL.n298 171.744
R394 VTAIL.n337 VTAIL.n298 171.744
R395 VTAIL.n337 VTAIL.n336 171.744
R396 VTAIL.n336 VTAIL.n302 171.744
R397 VTAIL.n329 VTAIL.n302 171.744
R398 VTAIL.n329 VTAIL.n328 171.744
R399 VTAIL.n328 VTAIL.n306 171.744
R400 VTAIL.n321 VTAIL.n306 171.744
R401 VTAIL.n321 VTAIL.n320 171.744
R402 VTAIL.n320 VTAIL.n310 171.744
R403 VTAIL.n313 VTAIL.n310 171.744
R404 VTAIL.n688 VTAIL.t3 85.8723
R405 VTAIL.n30 VTAIL.t1 85.8723
R406 VTAIL.n124 VTAIL.t4 85.8723
R407 VTAIL.n218 VTAIL.t7 85.8723
R408 VTAIL.n595 VTAIL.t6 85.8723
R409 VTAIL.n501 VTAIL.t5 85.8723
R410 VTAIL.n407 VTAIL.t2 85.8723
R411 VTAIL.n313 VTAIL.t0 85.8723
R412 VTAIL.n751 VTAIL.n750 35.8702
R413 VTAIL.n93 VTAIL.n92 35.8702
R414 VTAIL.n187 VTAIL.n186 35.8702
R415 VTAIL.n281 VTAIL.n280 35.8702
R416 VTAIL.n657 VTAIL.n656 35.8702
R417 VTAIL.n563 VTAIL.n562 35.8702
R418 VTAIL.n469 VTAIL.n468 35.8702
R419 VTAIL.n375 VTAIL.n374 35.8702
R420 VTAIL.n751 VTAIL.n657 28.6514
R421 VTAIL.n375 VTAIL.n281 28.6514
R422 VTAIL.n689 VTAIL.n687 16.3895
R423 VTAIL.n31 VTAIL.n29 16.3895
R424 VTAIL.n125 VTAIL.n123 16.3895
R425 VTAIL.n219 VTAIL.n217 16.3895
R426 VTAIL.n596 VTAIL.n594 16.3895
R427 VTAIL.n502 VTAIL.n500 16.3895
R428 VTAIL.n408 VTAIL.n406 16.3895
R429 VTAIL.n314 VTAIL.n312 16.3895
R430 VTAIL.n736 VTAIL.n735 13.1884
R431 VTAIL.n78 VTAIL.n77 13.1884
R432 VTAIL.n172 VTAIL.n171 13.1884
R433 VTAIL.n266 VTAIL.n265 13.1884
R434 VTAIL.n642 VTAIL.n641 13.1884
R435 VTAIL.n548 VTAIL.n547 13.1884
R436 VTAIL.n454 VTAIL.n453 13.1884
R437 VTAIL.n360 VTAIL.n359 13.1884
R438 VTAIL.n690 VTAIL.n686 12.8005
R439 VTAIL.n734 VTAIL.n666 12.8005
R440 VTAIL.n739 VTAIL.n664 12.8005
R441 VTAIL.n32 VTAIL.n28 12.8005
R442 VTAIL.n76 VTAIL.n8 12.8005
R443 VTAIL.n81 VTAIL.n6 12.8005
R444 VTAIL.n126 VTAIL.n122 12.8005
R445 VTAIL.n170 VTAIL.n102 12.8005
R446 VTAIL.n175 VTAIL.n100 12.8005
R447 VTAIL.n220 VTAIL.n216 12.8005
R448 VTAIL.n264 VTAIL.n196 12.8005
R449 VTAIL.n269 VTAIL.n194 12.8005
R450 VTAIL.n645 VTAIL.n570 12.8005
R451 VTAIL.n640 VTAIL.n572 12.8005
R452 VTAIL.n597 VTAIL.n593 12.8005
R453 VTAIL.n551 VTAIL.n476 12.8005
R454 VTAIL.n546 VTAIL.n478 12.8005
R455 VTAIL.n503 VTAIL.n499 12.8005
R456 VTAIL.n457 VTAIL.n382 12.8005
R457 VTAIL.n452 VTAIL.n384 12.8005
R458 VTAIL.n409 VTAIL.n405 12.8005
R459 VTAIL.n363 VTAIL.n288 12.8005
R460 VTAIL.n358 VTAIL.n290 12.8005
R461 VTAIL.n315 VTAIL.n311 12.8005
R462 VTAIL.n694 VTAIL.n693 12.0247
R463 VTAIL.n731 VTAIL.n730 12.0247
R464 VTAIL.n740 VTAIL.n662 12.0247
R465 VTAIL.n36 VTAIL.n35 12.0247
R466 VTAIL.n73 VTAIL.n72 12.0247
R467 VTAIL.n82 VTAIL.n4 12.0247
R468 VTAIL.n130 VTAIL.n129 12.0247
R469 VTAIL.n167 VTAIL.n166 12.0247
R470 VTAIL.n176 VTAIL.n98 12.0247
R471 VTAIL.n224 VTAIL.n223 12.0247
R472 VTAIL.n261 VTAIL.n260 12.0247
R473 VTAIL.n270 VTAIL.n192 12.0247
R474 VTAIL.n646 VTAIL.n568 12.0247
R475 VTAIL.n637 VTAIL.n636 12.0247
R476 VTAIL.n601 VTAIL.n600 12.0247
R477 VTAIL.n552 VTAIL.n474 12.0247
R478 VTAIL.n543 VTAIL.n542 12.0247
R479 VTAIL.n507 VTAIL.n506 12.0247
R480 VTAIL.n458 VTAIL.n380 12.0247
R481 VTAIL.n449 VTAIL.n448 12.0247
R482 VTAIL.n413 VTAIL.n412 12.0247
R483 VTAIL.n364 VTAIL.n286 12.0247
R484 VTAIL.n355 VTAIL.n354 12.0247
R485 VTAIL.n319 VTAIL.n318 12.0247
R486 VTAIL.n697 VTAIL.n684 11.249
R487 VTAIL.n726 VTAIL.n668 11.249
R488 VTAIL.n744 VTAIL.n743 11.249
R489 VTAIL.n39 VTAIL.n26 11.249
R490 VTAIL.n68 VTAIL.n10 11.249
R491 VTAIL.n86 VTAIL.n85 11.249
R492 VTAIL.n133 VTAIL.n120 11.249
R493 VTAIL.n162 VTAIL.n104 11.249
R494 VTAIL.n180 VTAIL.n179 11.249
R495 VTAIL.n227 VTAIL.n214 11.249
R496 VTAIL.n256 VTAIL.n198 11.249
R497 VTAIL.n274 VTAIL.n273 11.249
R498 VTAIL.n650 VTAIL.n649 11.249
R499 VTAIL.n633 VTAIL.n574 11.249
R500 VTAIL.n604 VTAIL.n591 11.249
R501 VTAIL.n556 VTAIL.n555 11.249
R502 VTAIL.n539 VTAIL.n480 11.249
R503 VTAIL.n510 VTAIL.n497 11.249
R504 VTAIL.n462 VTAIL.n461 11.249
R505 VTAIL.n445 VTAIL.n386 11.249
R506 VTAIL.n416 VTAIL.n403 11.249
R507 VTAIL.n368 VTAIL.n367 11.249
R508 VTAIL.n351 VTAIL.n292 11.249
R509 VTAIL.n322 VTAIL.n309 11.249
R510 VTAIL.n698 VTAIL.n682 10.4732
R511 VTAIL.n725 VTAIL.n670 10.4732
R512 VTAIL.n747 VTAIL.n660 10.4732
R513 VTAIL.n40 VTAIL.n24 10.4732
R514 VTAIL.n67 VTAIL.n12 10.4732
R515 VTAIL.n89 VTAIL.n2 10.4732
R516 VTAIL.n134 VTAIL.n118 10.4732
R517 VTAIL.n161 VTAIL.n106 10.4732
R518 VTAIL.n183 VTAIL.n96 10.4732
R519 VTAIL.n228 VTAIL.n212 10.4732
R520 VTAIL.n255 VTAIL.n200 10.4732
R521 VTAIL.n277 VTAIL.n190 10.4732
R522 VTAIL.n653 VTAIL.n566 10.4732
R523 VTAIL.n632 VTAIL.n577 10.4732
R524 VTAIL.n605 VTAIL.n589 10.4732
R525 VTAIL.n559 VTAIL.n472 10.4732
R526 VTAIL.n538 VTAIL.n483 10.4732
R527 VTAIL.n511 VTAIL.n495 10.4732
R528 VTAIL.n465 VTAIL.n378 10.4732
R529 VTAIL.n444 VTAIL.n389 10.4732
R530 VTAIL.n417 VTAIL.n401 10.4732
R531 VTAIL.n371 VTAIL.n284 10.4732
R532 VTAIL.n350 VTAIL.n295 10.4732
R533 VTAIL.n323 VTAIL.n307 10.4732
R534 VTAIL.n702 VTAIL.n701 9.69747
R535 VTAIL.n722 VTAIL.n721 9.69747
R536 VTAIL.n748 VTAIL.n658 9.69747
R537 VTAIL.n44 VTAIL.n43 9.69747
R538 VTAIL.n64 VTAIL.n63 9.69747
R539 VTAIL.n90 VTAIL.n0 9.69747
R540 VTAIL.n138 VTAIL.n137 9.69747
R541 VTAIL.n158 VTAIL.n157 9.69747
R542 VTAIL.n184 VTAIL.n94 9.69747
R543 VTAIL.n232 VTAIL.n231 9.69747
R544 VTAIL.n252 VTAIL.n251 9.69747
R545 VTAIL.n278 VTAIL.n188 9.69747
R546 VTAIL.n654 VTAIL.n564 9.69747
R547 VTAIL.n629 VTAIL.n628 9.69747
R548 VTAIL.n609 VTAIL.n608 9.69747
R549 VTAIL.n560 VTAIL.n470 9.69747
R550 VTAIL.n535 VTAIL.n534 9.69747
R551 VTAIL.n515 VTAIL.n514 9.69747
R552 VTAIL.n466 VTAIL.n376 9.69747
R553 VTAIL.n441 VTAIL.n440 9.69747
R554 VTAIL.n421 VTAIL.n420 9.69747
R555 VTAIL.n372 VTAIL.n282 9.69747
R556 VTAIL.n347 VTAIL.n346 9.69747
R557 VTAIL.n327 VTAIL.n326 9.69747
R558 VTAIL.n750 VTAIL.n749 9.45567
R559 VTAIL.n92 VTAIL.n91 9.45567
R560 VTAIL.n186 VTAIL.n185 9.45567
R561 VTAIL.n280 VTAIL.n279 9.45567
R562 VTAIL.n656 VTAIL.n655 9.45567
R563 VTAIL.n562 VTAIL.n561 9.45567
R564 VTAIL.n468 VTAIL.n467 9.45567
R565 VTAIL.n374 VTAIL.n373 9.45567
R566 VTAIL.n749 VTAIL.n748 9.3005
R567 VTAIL.n660 VTAIL.n659 9.3005
R568 VTAIL.n743 VTAIL.n742 9.3005
R569 VTAIL.n741 VTAIL.n740 9.3005
R570 VTAIL.n664 VTAIL.n663 9.3005
R571 VTAIL.n709 VTAIL.n708 9.3005
R572 VTAIL.n707 VTAIL.n706 9.3005
R573 VTAIL.n680 VTAIL.n679 9.3005
R574 VTAIL.n701 VTAIL.n700 9.3005
R575 VTAIL.n699 VTAIL.n698 9.3005
R576 VTAIL.n684 VTAIL.n683 9.3005
R577 VTAIL.n693 VTAIL.n692 9.3005
R578 VTAIL.n691 VTAIL.n690 9.3005
R579 VTAIL.n676 VTAIL.n675 9.3005
R580 VTAIL.n715 VTAIL.n714 9.3005
R581 VTAIL.n717 VTAIL.n716 9.3005
R582 VTAIL.n672 VTAIL.n671 9.3005
R583 VTAIL.n723 VTAIL.n722 9.3005
R584 VTAIL.n725 VTAIL.n724 9.3005
R585 VTAIL.n668 VTAIL.n667 9.3005
R586 VTAIL.n732 VTAIL.n731 9.3005
R587 VTAIL.n734 VTAIL.n733 9.3005
R588 VTAIL.n91 VTAIL.n90 9.3005
R589 VTAIL.n2 VTAIL.n1 9.3005
R590 VTAIL.n85 VTAIL.n84 9.3005
R591 VTAIL.n83 VTAIL.n82 9.3005
R592 VTAIL.n6 VTAIL.n5 9.3005
R593 VTAIL.n51 VTAIL.n50 9.3005
R594 VTAIL.n49 VTAIL.n48 9.3005
R595 VTAIL.n22 VTAIL.n21 9.3005
R596 VTAIL.n43 VTAIL.n42 9.3005
R597 VTAIL.n41 VTAIL.n40 9.3005
R598 VTAIL.n26 VTAIL.n25 9.3005
R599 VTAIL.n35 VTAIL.n34 9.3005
R600 VTAIL.n33 VTAIL.n32 9.3005
R601 VTAIL.n18 VTAIL.n17 9.3005
R602 VTAIL.n57 VTAIL.n56 9.3005
R603 VTAIL.n59 VTAIL.n58 9.3005
R604 VTAIL.n14 VTAIL.n13 9.3005
R605 VTAIL.n65 VTAIL.n64 9.3005
R606 VTAIL.n67 VTAIL.n66 9.3005
R607 VTAIL.n10 VTAIL.n9 9.3005
R608 VTAIL.n74 VTAIL.n73 9.3005
R609 VTAIL.n76 VTAIL.n75 9.3005
R610 VTAIL.n185 VTAIL.n184 9.3005
R611 VTAIL.n96 VTAIL.n95 9.3005
R612 VTAIL.n179 VTAIL.n178 9.3005
R613 VTAIL.n177 VTAIL.n176 9.3005
R614 VTAIL.n100 VTAIL.n99 9.3005
R615 VTAIL.n145 VTAIL.n144 9.3005
R616 VTAIL.n143 VTAIL.n142 9.3005
R617 VTAIL.n116 VTAIL.n115 9.3005
R618 VTAIL.n137 VTAIL.n136 9.3005
R619 VTAIL.n135 VTAIL.n134 9.3005
R620 VTAIL.n120 VTAIL.n119 9.3005
R621 VTAIL.n129 VTAIL.n128 9.3005
R622 VTAIL.n127 VTAIL.n126 9.3005
R623 VTAIL.n112 VTAIL.n111 9.3005
R624 VTAIL.n151 VTAIL.n150 9.3005
R625 VTAIL.n153 VTAIL.n152 9.3005
R626 VTAIL.n108 VTAIL.n107 9.3005
R627 VTAIL.n159 VTAIL.n158 9.3005
R628 VTAIL.n161 VTAIL.n160 9.3005
R629 VTAIL.n104 VTAIL.n103 9.3005
R630 VTAIL.n168 VTAIL.n167 9.3005
R631 VTAIL.n170 VTAIL.n169 9.3005
R632 VTAIL.n279 VTAIL.n278 9.3005
R633 VTAIL.n190 VTAIL.n189 9.3005
R634 VTAIL.n273 VTAIL.n272 9.3005
R635 VTAIL.n271 VTAIL.n270 9.3005
R636 VTAIL.n194 VTAIL.n193 9.3005
R637 VTAIL.n239 VTAIL.n238 9.3005
R638 VTAIL.n237 VTAIL.n236 9.3005
R639 VTAIL.n210 VTAIL.n209 9.3005
R640 VTAIL.n231 VTAIL.n230 9.3005
R641 VTAIL.n229 VTAIL.n228 9.3005
R642 VTAIL.n214 VTAIL.n213 9.3005
R643 VTAIL.n223 VTAIL.n222 9.3005
R644 VTAIL.n221 VTAIL.n220 9.3005
R645 VTAIL.n206 VTAIL.n205 9.3005
R646 VTAIL.n245 VTAIL.n244 9.3005
R647 VTAIL.n247 VTAIL.n246 9.3005
R648 VTAIL.n202 VTAIL.n201 9.3005
R649 VTAIL.n253 VTAIL.n252 9.3005
R650 VTAIL.n255 VTAIL.n254 9.3005
R651 VTAIL.n198 VTAIL.n197 9.3005
R652 VTAIL.n262 VTAIL.n261 9.3005
R653 VTAIL.n264 VTAIL.n263 9.3005
R654 VTAIL.n622 VTAIL.n621 9.3005
R655 VTAIL.n624 VTAIL.n623 9.3005
R656 VTAIL.n579 VTAIL.n578 9.3005
R657 VTAIL.n630 VTAIL.n629 9.3005
R658 VTAIL.n632 VTAIL.n631 9.3005
R659 VTAIL.n574 VTAIL.n573 9.3005
R660 VTAIL.n638 VTAIL.n637 9.3005
R661 VTAIL.n640 VTAIL.n639 9.3005
R662 VTAIL.n655 VTAIL.n654 9.3005
R663 VTAIL.n566 VTAIL.n565 9.3005
R664 VTAIL.n649 VTAIL.n648 9.3005
R665 VTAIL.n647 VTAIL.n646 9.3005
R666 VTAIL.n570 VTAIL.n569 9.3005
R667 VTAIL.n583 VTAIL.n582 9.3005
R668 VTAIL.n616 VTAIL.n615 9.3005
R669 VTAIL.n614 VTAIL.n613 9.3005
R670 VTAIL.n587 VTAIL.n586 9.3005
R671 VTAIL.n608 VTAIL.n607 9.3005
R672 VTAIL.n606 VTAIL.n605 9.3005
R673 VTAIL.n591 VTAIL.n590 9.3005
R674 VTAIL.n600 VTAIL.n599 9.3005
R675 VTAIL.n598 VTAIL.n597 9.3005
R676 VTAIL.n528 VTAIL.n527 9.3005
R677 VTAIL.n530 VTAIL.n529 9.3005
R678 VTAIL.n485 VTAIL.n484 9.3005
R679 VTAIL.n536 VTAIL.n535 9.3005
R680 VTAIL.n538 VTAIL.n537 9.3005
R681 VTAIL.n480 VTAIL.n479 9.3005
R682 VTAIL.n544 VTAIL.n543 9.3005
R683 VTAIL.n546 VTAIL.n545 9.3005
R684 VTAIL.n561 VTAIL.n560 9.3005
R685 VTAIL.n472 VTAIL.n471 9.3005
R686 VTAIL.n555 VTAIL.n554 9.3005
R687 VTAIL.n553 VTAIL.n552 9.3005
R688 VTAIL.n476 VTAIL.n475 9.3005
R689 VTAIL.n489 VTAIL.n488 9.3005
R690 VTAIL.n522 VTAIL.n521 9.3005
R691 VTAIL.n520 VTAIL.n519 9.3005
R692 VTAIL.n493 VTAIL.n492 9.3005
R693 VTAIL.n514 VTAIL.n513 9.3005
R694 VTAIL.n512 VTAIL.n511 9.3005
R695 VTAIL.n497 VTAIL.n496 9.3005
R696 VTAIL.n506 VTAIL.n505 9.3005
R697 VTAIL.n504 VTAIL.n503 9.3005
R698 VTAIL.n434 VTAIL.n433 9.3005
R699 VTAIL.n436 VTAIL.n435 9.3005
R700 VTAIL.n391 VTAIL.n390 9.3005
R701 VTAIL.n442 VTAIL.n441 9.3005
R702 VTAIL.n444 VTAIL.n443 9.3005
R703 VTAIL.n386 VTAIL.n385 9.3005
R704 VTAIL.n450 VTAIL.n449 9.3005
R705 VTAIL.n452 VTAIL.n451 9.3005
R706 VTAIL.n467 VTAIL.n466 9.3005
R707 VTAIL.n378 VTAIL.n377 9.3005
R708 VTAIL.n461 VTAIL.n460 9.3005
R709 VTAIL.n459 VTAIL.n458 9.3005
R710 VTAIL.n382 VTAIL.n381 9.3005
R711 VTAIL.n395 VTAIL.n394 9.3005
R712 VTAIL.n428 VTAIL.n427 9.3005
R713 VTAIL.n426 VTAIL.n425 9.3005
R714 VTAIL.n399 VTAIL.n398 9.3005
R715 VTAIL.n420 VTAIL.n419 9.3005
R716 VTAIL.n418 VTAIL.n417 9.3005
R717 VTAIL.n403 VTAIL.n402 9.3005
R718 VTAIL.n412 VTAIL.n411 9.3005
R719 VTAIL.n410 VTAIL.n409 9.3005
R720 VTAIL.n340 VTAIL.n339 9.3005
R721 VTAIL.n342 VTAIL.n341 9.3005
R722 VTAIL.n297 VTAIL.n296 9.3005
R723 VTAIL.n348 VTAIL.n347 9.3005
R724 VTAIL.n350 VTAIL.n349 9.3005
R725 VTAIL.n292 VTAIL.n291 9.3005
R726 VTAIL.n356 VTAIL.n355 9.3005
R727 VTAIL.n358 VTAIL.n357 9.3005
R728 VTAIL.n373 VTAIL.n372 9.3005
R729 VTAIL.n284 VTAIL.n283 9.3005
R730 VTAIL.n367 VTAIL.n366 9.3005
R731 VTAIL.n365 VTAIL.n364 9.3005
R732 VTAIL.n288 VTAIL.n287 9.3005
R733 VTAIL.n301 VTAIL.n300 9.3005
R734 VTAIL.n334 VTAIL.n333 9.3005
R735 VTAIL.n332 VTAIL.n331 9.3005
R736 VTAIL.n305 VTAIL.n304 9.3005
R737 VTAIL.n326 VTAIL.n325 9.3005
R738 VTAIL.n324 VTAIL.n323 9.3005
R739 VTAIL.n309 VTAIL.n308 9.3005
R740 VTAIL.n318 VTAIL.n317 9.3005
R741 VTAIL.n316 VTAIL.n315 9.3005
R742 VTAIL.n705 VTAIL.n680 8.92171
R743 VTAIL.n718 VTAIL.n672 8.92171
R744 VTAIL.n47 VTAIL.n22 8.92171
R745 VTAIL.n60 VTAIL.n14 8.92171
R746 VTAIL.n141 VTAIL.n116 8.92171
R747 VTAIL.n154 VTAIL.n108 8.92171
R748 VTAIL.n235 VTAIL.n210 8.92171
R749 VTAIL.n248 VTAIL.n202 8.92171
R750 VTAIL.n625 VTAIL.n579 8.92171
R751 VTAIL.n612 VTAIL.n587 8.92171
R752 VTAIL.n531 VTAIL.n485 8.92171
R753 VTAIL.n518 VTAIL.n493 8.92171
R754 VTAIL.n437 VTAIL.n391 8.92171
R755 VTAIL.n424 VTAIL.n399 8.92171
R756 VTAIL.n343 VTAIL.n297 8.92171
R757 VTAIL.n330 VTAIL.n305 8.92171
R758 VTAIL.n706 VTAIL.n678 8.14595
R759 VTAIL.n717 VTAIL.n674 8.14595
R760 VTAIL.n48 VTAIL.n20 8.14595
R761 VTAIL.n59 VTAIL.n16 8.14595
R762 VTAIL.n142 VTAIL.n114 8.14595
R763 VTAIL.n153 VTAIL.n110 8.14595
R764 VTAIL.n236 VTAIL.n208 8.14595
R765 VTAIL.n247 VTAIL.n204 8.14595
R766 VTAIL.n624 VTAIL.n581 8.14595
R767 VTAIL.n613 VTAIL.n585 8.14595
R768 VTAIL.n530 VTAIL.n487 8.14595
R769 VTAIL.n519 VTAIL.n491 8.14595
R770 VTAIL.n436 VTAIL.n393 8.14595
R771 VTAIL.n425 VTAIL.n397 8.14595
R772 VTAIL.n342 VTAIL.n299 8.14595
R773 VTAIL.n331 VTAIL.n303 8.14595
R774 VTAIL.n710 VTAIL.n709 7.3702
R775 VTAIL.n714 VTAIL.n713 7.3702
R776 VTAIL.n52 VTAIL.n51 7.3702
R777 VTAIL.n56 VTAIL.n55 7.3702
R778 VTAIL.n146 VTAIL.n145 7.3702
R779 VTAIL.n150 VTAIL.n149 7.3702
R780 VTAIL.n240 VTAIL.n239 7.3702
R781 VTAIL.n244 VTAIL.n243 7.3702
R782 VTAIL.n621 VTAIL.n620 7.3702
R783 VTAIL.n617 VTAIL.n616 7.3702
R784 VTAIL.n527 VTAIL.n526 7.3702
R785 VTAIL.n523 VTAIL.n522 7.3702
R786 VTAIL.n433 VTAIL.n432 7.3702
R787 VTAIL.n429 VTAIL.n428 7.3702
R788 VTAIL.n339 VTAIL.n338 7.3702
R789 VTAIL.n335 VTAIL.n334 7.3702
R790 VTAIL.n710 VTAIL.n676 6.59444
R791 VTAIL.n713 VTAIL.n676 6.59444
R792 VTAIL.n52 VTAIL.n18 6.59444
R793 VTAIL.n55 VTAIL.n18 6.59444
R794 VTAIL.n146 VTAIL.n112 6.59444
R795 VTAIL.n149 VTAIL.n112 6.59444
R796 VTAIL.n240 VTAIL.n206 6.59444
R797 VTAIL.n243 VTAIL.n206 6.59444
R798 VTAIL.n620 VTAIL.n583 6.59444
R799 VTAIL.n617 VTAIL.n583 6.59444
R800 VTAIL.n526 VTAIL.n489 6.59444
R801 VTAIL.n523 VTAIL.n489 6.59444
R802 VTAIL.n432 VTAIL.n395 6.59444
R803 VTAIL.n429 VTAIL.n395 6.59444
R804 VTAIL.n338 VTAIL.n301 6.59444
R805 VTAIL.n335 VTAIL.n301 6.59444
R806 VTAIL.n709 VTAIL.n678 5.81868
R807 VTAIL.n714 VTAIL.n674 5.81868
R808 VTAIL.n51 VTAIL.n20 5.81868
R809 VTAIL.n56 VTAIL.n16 5.81868
R810 VTAIL.n145 VTAIL.n114 5.81868
R811 VTAIL.n150 VTAIL.n110 5.81868
R812 VTAIL.n239 VTAIL.n208 5.81868
R813 VTAIL.n244 VTAIL.n204 5.81868
R814 VTAIL.n621 VTAIL.n581 5.81868
R815 VTAIL.n616 VTAIL.n585 5.81868
R816 VTAIL.n527 VTAIL.n487 5.81868
R817 VTAIL.n522 VTAIL.n491 5.81868
R818 VTAIL.n433 VTAIL.n393 5.81868
R819 VTAIL.n428 VTAIL.n397 5.81868
R820 VTAIL.n339 VTAIL.n299 5.81868
R821 VTAIL.n334 VTAIL.n303 5.81868
R822 VTAIL.n706 VTAIL.n705 5.04292
R823 VTAIL.n718 VTAIL.n717 5.04292
R824 VTAIL.n48 VTAIL.n47 5.04292
R825 VTAIL.n60 VTAIL.n59 5.04292
R826 VTAIL.n142 VTAIL.n141 5.04292
R827 VTAIL.n154 VTAIL.n153 5.04292
R828 VTAIL.n236 VTAIL.n235 5.04292
R829 VTAIL.n248 VTAIL.n247 5.04292
R830 VTAIL.n625 VTAIL.n624 5.04292
R831 VTAIL.n613 VTAIL.n612 5.04292
R832 VTAIL.n531 VTAIL.n530 5.04292
R833 VTAIL.n519 VTAIL.n518 5.04292
R834 VTAIL.n437 VTAIL.n436 5.04292
R835 VTAIL.n425 VTAIL.n424 5.04292
R836 VTAIL.n343 VTAIL.n342 5.04292
R837 VTAIL.n331 VTAIL.n330 5.04292
R838 VTAIL.n702 VTAIL.n680 4.26717
R839 VTAIL.n721 VTAIL.n672 4.26717
R840 VTAIL.n750 VTAIL.n658 4.26717
R841 VTAIL.n44 VTAIL.n22 4.26717
R842 VTAIL.n63 VTAIL.n14 4.26717
R843 VTAIL.n92 VTAIL.n0 4.26717
R844 VTAIL.n138 VTAIL.n116 4.26717
R845 VTAIL.n157 VTAIL.n108 4.26717
R846 VTAIL.n186 VTAIL.n94 4.26717
R847 VTAIL.n232 VTAIL.n210 4.26717
R848 VTAIL.n251 VTAIL.n202 4.26717
R849 VTAIL.n280 VTAIL.n188 4.26717
R850 VTAIL.n656 VTAIL.n564 4.26717
R851 VTAIL.n628 VTAIL.n579 4.26717
R852 VTAIL.n609 VTAIL.n587 4.26717
R853 VTAIL.n562 VTAIL.n470 4.26717
R854 VTAIL.n534 VTAIL.n485 4.26717
R855 VTAIL.n515 VTAIL.n493 4.26717
R856 VTAIL.n468 VTAIL.n376 4.26717
R857 VTAIL.n440 VTAIL.n391 4.26717
R858 VTAIL.n421 VTAIL.n399 4.26717
R859 VTAIL.n374 VTAIL.n282 4.26717
R860 VTAIL.n346 VTAIL.n297 4.26717
R861 VTAIL.n327 VTAIL.n305 4.26717
R862 VTAIL.n691 VTAIL.n687 3.70982
R863 VTAIL.n33 VTAIL.n29 3.70982
R864 VTAIL.n127 VTAIL.n123 3.70982
R865 VTAIL.n221 VTAIL.n217 3.70982
R866 VTAIL.n598 VTAIL.n594 3.70982
R867 VTAIL.n504 VTAIL.n500 3.70982
R868 VTAIL.n410 VTAIL.n406 3.70982
R869 VTAIL.n316 VTAIL.n312 3.70982
R870 VTAIL.n701 VTAIL.n682 3.49141
R871 VTAIL.n722 VTAIL.n670 3.49141
R872 VTAIL.n748 VTAIL.n747 3.49141
R873 VTAIL.n43 VTAIL.n24 3.49141
R874 VTAIL.n64 VTAIL.n12 3.49141
R875 VTAIL.n90 VTAIL.n89 3.49141
R876 VTAIL.n137 VTAIL.n118 3.49141
R877 VTAIL.n158 VTAIL.n106 3.49141
R878 VTAIL.n184 VTAIL.n183 3.49141
R879 VTAIL.n231 VTAIL.n212 3.49141
R880 VTAIL.n252 VTAIL.n200 3.49141
R881 VTAIL.n278 VTAIL.n277 3.49141
R882 VTAIL.n654 VTAIL.n653 3.49141
R883 VTAIL.n629 VTAIL.n577 3.49141
R884 VTAIL.n608 VTAIL.n589 3.49141
R885 VTAIL.n560 VTAIL.n559 3.49141
R886 VTAIL.n535 VTAIL.n483 3.49141
R887 VTAIL.n514 VTAIL.n495 3.49141
R888 VTAIL.n466 VTAIL.n465 3.49141
R889 VTAIL.n441 VTAIL.n389 3.49141
R890 VTAIL.n420 VTAIL.n401 3.49141
R891 VTAIL.n372 VTAIL.n371 3.49141
R892 VTAIL.n347 VTAIL.n295 3.49141
R893 VTAIL.n326 VTAIL.n307 3.49141
R894 VTAIL.n698 VTAIL.n697 2.71565
R895 VTAIL.n726 VTAIL.n725 2.71565
R896 VTAIL.n744 VTAIL.n660 2.71565
R897 VTAIL.n40 VTAIL.n39 2.71565
R898 VTAIL.n68 VTAIL.n67 2.71565
R899 VTAIL.n86 VTAIL.n2 2.71565
R900 VTAIL.n134 VTAIL.n133 2.71565
R901 VTAIL.n162 VTAIL.n161 2.71565
R902 VTAIL.n180 VTAIL.n96 2.71565
R903 VTAIL.n228 VTAIL.n227 2.71565
R904 VTAIL.n256 VTAIL.n255 2.71565
R905 VTAIL.n274 VTAIL.n190 2.71565
R906 VTAIL.n650 VTAIL.n566 2.71565
R907 VTAIL.n633 VTAIL.n632 2.71565
R908 VTAIL.n605 VTAIL.n604 2.71565
R909 VTAIL.n556 VTAIL.n472 2.71565
R910 VTAIL.n539 VTAIL.n538 2.71565
R911 VTAIL.n511 VTAIL.n510 2.71565
R912 VTAIL.n462 VTAIL.n378 2.71565
R913 VTAIL.n445 VTAIL.n444 2.71565
R914 VTAIL.n417 VTAIL.n416 2.71565
R915 VTAIL.n368 VTAIL.n284 2.71565
R916 VTAIL.n351 VTAIL.n350 2.71565
R917 VTAIL.n323 VTAIL.n322 2.71565
R918 VTAIL.n694 VTAIL.n684 1.93989
R919 VTAIL.n730 VTAIL.n668 1.93989
R920 VTAIL.n743 VTAIL.n662 1.93989
R921 VTAIL.n36 VTAIL.n26 1.93989
R922 VTAIL.n72 VTAIL.n10 1.93989
R923 VTAIL.n85 VTAIL.n4 1.93989
R924 VTAIL.n130 VTAIL.n120 1.93989
R925 VTAIL.n166 VTAIL.n104 1.93989
R926 VTAIL.n179 VTAIL.n98 1.93989
R927 VTAIL.n224 VTAIL.n214 1.93989
R928 VTAIL.n260 VTAIL.n198 1.93989
R929 VTAIL.n273 VTAIL.n192 1.93989
R930 VTAIL.n649 VTAIL.n568 1.93989
R931 VTAIL.n636 VTAIL.n574 1.93989
R932 VTAIL.n601 VTAIL.n591 1.93989
R933 VTAIL.n555 VTAIL.n474 1.93989
R934 VTAIL.n542 VTAIL.n480 1.93989
R935 VTAIL.n507 VTAIL.n497 1.93989
R936 VTAIL.n461 VTAIL.n380 1.93989
R937 VTAIL.n448 VTAIL.n386 1.93989
R938 VTAIL.n413 VTAIL.n403 1.93989
R939 VTAIL.n367 VTAIL.n286 1.93989
R940 VTAIL.n354 VTAIL.n292 1.93989
R941 VTAIL.n319 VTAIL.n309 1.93989
R942 VTAIL.n469 VTAIL.n375 1.63843
R943 VTAIL.n657 VTAIL.n563 1.63843
R944 VTAIL.n281 VTAIL.n187 1.63843
R945 VTAIL.n693 VTAIL.n686 1.16414
R946 VTAIL.n731 VTAIL.n666 1.16414
R947 VTAIL.n740 VTAIL.n739 1.16414
R948 VTAIL.n35 VTAIL.n28 1.16414
R949 VTAIL.n73 VTAIL.n8 1.16414
R950 VTAIL.n82 VTAIL.n81 1.16414
R951 VTAIL.n129 VTAIL.n122 1.16414
R952 VTAIL.n167 VTAIL.n102 1.16414
R953 VTAIL.n176 VTAIL.n175 1.16414
R954 VTAIL.n223 VTAIL.n216 1.16414
R955 VTAIL.n261 VTAIL.n196 1.16414
R956 VTAIL.n270 VTAIL.n269 1.16414
R957 VTAIL.n646 VTAIL.n645 1.16414
R958 VTAIL.n637 VTAIL.n572 1.16414
R959 VTAIL.n600 VTAIL.n593 1.16414
R960 VTAIL.n552 VTAIL.n551 1.16414
R961 VTAIL.n543 VTAIL.n478 1.16414
R962 VTAIL.n506 VTAIL.n499 1.16414
R963 VTAIL.n458 VTAIL.n457 1.16414
R964 VTAIL.n449 VTAIL.n384 1.16414
R965 VTAIL.n412 VTAIL.n405 1.16414
R966 VTAIL.n364 VTAIL.n363 1.16414
R967 VTAIL.n355 VTAIL.n290 1.16414
R968 VTAIL.n318 VTAIL.n311 1.16414
R969 VTAIL VTAIL.n93 0.877655
R970 VTAIL VTAIL.n751 0.761276
R971 VTAIL.n563 VTAIL.n469 0.470328
R972 VTAIL.n187 VTAIL.n93 0.470328
R973 VTAIL.n690 VTAIL.n689 0.388379
R974 VTAIL.n735 VTAIL.n734 0.388379
R975 VTAIL.n736 VTAIL.n664 0.388379
R976 VTAIL.n32 VTAIL.n31 0.388379
R977 VTAIL.n77 VTAIL.n76 0.388379
R978 VTAIL.n78 VTAIL.n6 0.388379
R979 VTAIL.n126 VTAIL.n125 0.388379
R980 VTAIL.n171 VTAIL.n170 0.388379
R981 VTAIL.n172 VTAIL.n100 0.388379
R982 VTAIL.n220 VTAIL.n219 0.388379
R983 VTAIL.n265 VTAIL.n264 0.388379
R984 VTAIL.n266 VTAIL.n194 0.388379
R985 VTAIL.n642 VTAIL.n570 0.388379
R986 VTAIL.n641 VTAIL.n640 0.388379
R987 VTAIL.n597 VTAIL.n596 0.388379
R988 VTAIL.n548 VTAIL.n476 0.388379
R989 VTAIL.n547 VTAIL.n546 0.388379
R990 VTAIL.n503 VTAIL.n502 0.388379
R991 VTAIL.n454 VTAIL.n382 0.388379
R992 VTAIL.n453 VTAIL.n452 0.388379
R993 VTAIL.n409 VTAIL.n408 0.388379
R994 VTAIL.n360 VTAIL.n288 0.388379
R995 VTAIL.n359 VTAIL.n358 0.388379
R996 VTAIL.n315 VTAIL.n314 0.388379
R997 VTAIL.n692 VTAIL.n691 0.155672
R998 VTAIL.n692 VTAIL.n683 0.155672
R999 VTAIL.n699 VTAIL.n683 0.155672
R1000 VTAIL.n700 VTAIL.n699 0.155672
R1001 VTAIL.n700 VTAIL.n679 0.155672
R1002 VTAIL.n707 VTAIL.n679 0.155672
R1003 VTAIL.n708 VTAIL.n707 0.155672
R1004 VTAIL.n708 VTAIL.n675 0.155672
R1005 VTAIL.n715 VTAIL.n675 0.155672
R1006 VTAIL.n716 VTAIL.n715 0.155672
R1007 VTAIL.n716 VTAIL.n671 0.155672
R1008 VTAIL.n723 VTAIL.n671 0.155672
R1009 VTAIL.n724 VTAIL.n723 0.155672
R1010 VTAIL.n724 VTAIL.n667 0.155672
R1011 VTAIL.n732 VTAIL.n667 0.155672
R1012 VTAIL.n733 VTAIL.n732 0.155672
R1013 VTAIL.n733 VTAIL.n663 0.155672
R1014 VTAIL.n741 VTAIL.n663 0.155672
R1015 VTAIL.n742 VTAIL.n741 0.155672
R1016 VTAIL.n742 VTAIL.n659 0.155672
R1017 VTAIL.n749 VTAIL.n659 0.155672
R1018 VTAIL.n34 VTAIL.n33 0.155672
R1019 VTAIL.n34 VTAIL.n25 0.155672
R1020 VTAIL.n41 VTAIL.n25 0.155672
R1021 VTAIL.n42 VTAIL.n41 0.155672
R1022 VTAIL.n42 VTAIL.n21 0.155672
R1023 VTAIL.n49 VTAIL.n21 0.155672
R1024 VTAIL.n50 VTAIL.n49 0.155672
R1025 VTAIL.n50 VTAIL.n17 0.155672
R1026 VTAIL.n57 VTAIL.n17 0.155672
R1027 VTAIL.n58 VTAIL.n57 0.155672
R1028 VTAIL.n58 VTAIL.n13 0.155672
R1029 VTAIL.n65 VTAIL.n13 0.155672
R1030 VTAIL.n66 VTAIL.n65 0.155672
R1031 VTAIL.n66 VTAIL.n9 0.155672
R1032 VTAIL.n74 VTAIL.n9 0.155672
R1033 VTAIL.n75 VTAIL.n74 0.155672
R1034 VTAIL.n75 VTAIL.n5 0.155672
R1035 VTAIL.n83 VTAIL.n5 0.155672
R1036 VTAIL.n84 VTAIL.n83 0.155672
R1037 VTAIL.n84 VTAIL.n1 0.155672
R1038 VTAIL.n91 VTAIL.n1 0.155672
R1039 VTAIL.n128 VTAIL.n127 0.155672
R1040 VTAIL.n128 VTAIL.n119 0.155672
R1041 VTAIL.n135 VTAIL.n119 0.155672
R1042 VTAIL.n136 VTAIL.n135 0.155672
R1043 VTAIL.n136 VTAIL.n115 0.155672
R1044 VTAIL.n143 VTAIL.n115 0.155672
R1045 VTAIL.n144 VTAIL.n143 0.155672
R1046 VTAIL.n144 VTAIL.n111 0.155672
R1047 VTAIL.n151 VTAIL.n111 0.155672
R1048 VTAIL.n152 VTAIL.n151 0.155672
R1049 VTAIL.n152 VTAIL.n107 0.155672
R1050 VTAIL.n159 VTAIL.n107 0.155672
R1051 VTAIL.n160 VTAIL.n159 0.155672
R1052 VTAIL.n160 VTAIL.n103 0.155672
R1053 VTAIL.n168 VTAIL.n103 0.155672
R1054 VTAIL.n169 VTAIL.n168 0.155672
R1055 VTAIL.n169 VTAIL.n99 0.155672
R1056 VTAIL.n177 VTAIL.n99 0.155672
R1057 VTAIL.n178 VTAIL.n177 0.155672
R1058 VTAIL.n178 VTAIL.n95 0.155672
R1059 VTAIL.n185 VTAIL.n95 0.155672
R1060 VTAIL.n222 VTAIL.n221 0.155672
R1061 VTAIL.n222 VTAIL.n213 0.155672
R1062 VTAIL.n229 VTAIL.n213 0.155672
R1063 VTAIL.n230 VTAIL.n229 0.155672
R1064 VTAIL.n230 VTAIL.n209 0.155672
R1065 VTAIL.n237 VTAIL.n209 0.155672
R1066 VTAIL.n238 VTAIL.n237 0.155672
R1067 VTAIL.n238 VTAIL.n205 0.155672
R1068 VTAIL.n245 VTAIL.n205 0.155672
R1069 VTAIL.n246 VTAIL.n245 0.155672
R1070 VTAIL.n246 VTAIL.n201 0.155672
R1071 VTAIL.n253 VTAIL.n201 0.155672
R1072 VTAIL.n254 VTAIL.n253 0.155672
R1073 VTAIL.n254 VTAIL.n197 0.155672
R1074 VTAIL.n262 VTAIL.n197 0.155672
R1075 VTAIL.n263 VTAIL.n262 0.155672
R1076 VTAIL.n263 VTAIL.n193 0.155672
R1077 VTAIL.n271 VTAIL.n193 0.155672
R1078 VTAIL.n272 VTAIL.n271 0.155672
R1079 VTAIL.n272 VTAIL.n189 0.155672
R1080 VTAIL.n279 VTAIL.n189 0.155672
R1081 VTAIL.n655 VTAIL.n565 0.155672
R1082 VTAIL.n648 VTAIL.n565 0.155672
R1083 VTAIL.n648 VTAIL.n647 0.155672
R1084 VTAIL.n647 VTAIL.n569 0.155672
R1085 VTAIL.n639 VTAIL.n569 0.155672
R1086 VTAIL.n639 VTAIL.n638 0.155672
R1087 VTAIL.n638 VTAIL.n573 0.155672
R1088 VTAIL.n631 VTAIL.n573 0.155672
R1089 VTAIL.n631 VTAIL.n630 0.155672
R1090 VTAIL.n630 VTAIL.n578 0.155672
R1091 VTAIL.n623 VTAIL.n578 0.155672
R1092 VTAIL.n623 VTAIL.n622 0.155672
R1093 VTAIL.n622 VTAIL.n582 0.155672
R1094 VTAIL.n615 VTAIL.n582 0.155672
R1095 VTAIL.n615 VTAIL.n614 0.155672
R1096 VTAIL.n614 VTAIL.n586 0.155672
R1097 VTAIL.n607 VTAIL.n586 0.155672
R1098 VTAIL.n607 VTAIL.n606 0.155672
R1099 VTAIL.n606 VTAIL.n590 0.155672
R1100 VTAIL.n599 VTAIL.n590 0.155672
R1101 VTAIL.n599 VTAIL.n598 0.155672
R1102 VTAIL.n561 VTAIL.n471 0.155672
R1103 VTAIL.n554 VTAIL.n471 0.155672
R1104 VTAIL.n554 VTAIL.n553 0.155672
R1105 VTAIL.n553 VTAIL.n475 0.155672
R1106 VTAIL.n545 VTAIL.n475 0.155672
R1107 VTAIL.n545 VTAIL.n544 0.155672
R1108 VTAIL.n544 VTAIL.n479 0.155672
R1109 VTAIL.n537 VTAIL.n479 0.155672
R1110 VTAIL.n537 VTAIL.n536 0.155672
R1111 VTAIL.n536 VTAIL.n484 0.155672
R1112 VTAIL.n529 VTAIL.n484 0.155672
R1113 VTAIL.n529 VTAIL.n528 0.155672
R1114 VTAIL.n528 VTAIL.n488 0.155672
R1115 VTAIL.n521 VTAIL.n488 0.155672
R1116 VTAIL.n521 VTAIL.n520 0.155672
R1117 VTAIL.n520 VTAIL.n492 0.155672
R1118 VTAIL.n513 VTAIL.n492 0.155672
R1119 VTAIL.n513 VTAIL.n512 0.155672
R1120 VTAIL.n512 VTAIL.n496 0.155672
R1121 VTAIL.n505 VTAIL.n496 0.155672
R1122 VTAIL.n505 VTAIL.n504 0.155672
R1123 VTAIL.n467 VTAIL.n377 0.155672
R1124 VTAIL.n460 VTAIL.n377 0.155672
R1125 VTAIL.n460 VTAIL.n459 0.155672
R1126 VTAIL.n459 VTAIL.n381 0.155672
R1127 VTAIL.n451 VTAIL.n381 0.155672
R1128 VTAIL.n451 VTAIL.n450 0.155672
R1129 VTAIL.n450 VTAIL.n385 0.155672
R1130 VTAIL.n443 VTAIL.n385 0.155672
R1131 VTAIL.n443 VTAIL.n442 0.155672
R1132 VTAIL.n442 VTAIL.n390 0.155672
R1133 VTAIL.n435 VTAIL.n390 0.155672
R1134 VTAIL.n435 VTAIL.n434 0.155672
R1135 VTAIL.n434 VTAIL.n394 0.155672
R1136 VTAIL.n427 VTAIL.n394 0.155672
R1137 VTAIL.n427 VTAIL.n426 0.155672
R1138 VTAIL.n426 VTAIL.n398 0.155672
R1139 VTAIL.n419 VTAIL.n398 0.155672
R1140 VTAIL.n419 VTAIL.n418 0.155672
R1141 VTAIL.n418 VTAIL.n402 0.155672
R1142 VTAIL.n411 VTAIL.n402 0.155672
R1143 VTAIL.n411 VTAIL.n410 0.155672
R1144 VTAIL.n373 VTAIL.n283 0.155672
R1145 VTAIL.n366 VTAIL.n283 0.155672
R1146 VTAIL.n366 VTAIL.n365 0.155672
R1147 VTAIL.n365 VTAIL.n287 0.155672
R1148 VTAIL.n357 VTAIL.n287 0.155672
R1149 VTAIL.n357 VTAIL.n356 0.155672
R1150 VTAIL.n356 VTAIL.n291 0.155672
R1151 VTAIL.n349 VTAIL.n291 0.155672
R1152 VTAIL.n349 VTAIL.n348 0.155672
R1153 VTAIL.n348 VTAIL.n296 0.155672
R1154 VTAIL.n341 VTAIL.n296 0.155672
R1155 VTAIL.n341 VTAIL.n340 0.155672
R1156 VTAIL.n340 VTAIL.n300 0.155672
R1157 VTAIL.n333 VTAIL.n300 0.155672
R1158 VTAIL.n333 VTAIL.n332 0.155672
R1159 VTAIL.n332 VTAIL.n304 0.155672
R1160 VTAIL.n325 VTAIL.n304 0.155672
R1161 VTAIL.n325 VTAIL.n324 0.155672
R1162 VTAIL.n324 VTAIL.n308 0.155672
R1163 VTAIL.n317 VTAIL.n308 0.155672
R1164 VTAIL.n317 VTAIL.n316 0.155672
R1165 VN.n0 VN.t1 298.171
R1166 VN.n1 VN.t0 298.171
R1167 VN.n0 VN.t2 297.848
R1168 VN.n1 VN.t3 297.848
R1169 VN VN.n1 60.064
R1170 VN VN.n0 12.8178
R1171 VDD2.n2 VDD2.n0 116.352
R1172 VDD2.n2 VDD2.n1 73.0767
R1173 VDD2.n1 VDD2.t0 1.91368
R1174 VDD2.n1 VDD2.t3 1.91368
R1175 VDD2.n0 VDD2.t2 1.91368
R1176 VDD2.n0 VDD2.t1 1.91368
R1177 VDD2 VDD2.n2 0.0586897
R1178 B.n481 B.n80 585
R1179 B.n483 B.n482 585
R1180 B.n484 B.n79 585
R1181 B.n486 B.n485 585
R1182 B.n487 B.n78 585
R1183 B.n489 B.n488 585
R1184 B.n490 B.n77 585
R1185 B.n492 B.n491 585
R1186 B.n493 B.n76 585
R1187 B.n495 B.n494 585
R1188 B.n496 B.n75 585
R1189 B.n498 B.n497 585
R1190 B.n499 B.n74 585
R1191 B.n501 B.n500 585
R1192 B.n502 B.n73 585
R1193 B.n504 B.n503 585
R1194 B.n505 B.n72 585
R1195 B.n507 B.n506 585
R1196 B.n508 B.n71 585
R1197 B.n510 B.n509 585
R1198 B.n511 B.n70 585
R1199 B.n513 B.n512 585
R1200 B.n514 B.n69 585
R1201 B.n516 B.n515 585
R1202 B.n517 B.n68 585
R1203 B.n519 B.n518 585
R1204 B.n520 B.n67 585
R1205 B.n522 B.n521 585
R1206 B.n523 B.n66 585
R1207 B.n525 B.n524 585
R1208 B.n526 B.n65 585
R1209 B.n528 B.n527 585
R1210 B.n529 B.n64 585
R1211 B.n531 B.n530 585
R1212 B.n532 B.n63 585
R1213 B.n534 B.n533 585
R1214 B.n535 B.n62 585
R1215 B.n537 B.n536 585
R1216 B.n538 B.n61 585
R1217 B.n540 B.n539 585
R1218 B.n541 B.n60 585
R1219 B.n543 B.n542 585
R1220 B.n544 B.n59 585
R1221 B.n546 B.n545 585
R1222 B.n547 B.n58 585
R1223 B.n549 B.n548 585
R1224 B.n550 B.n57 585
R1225 B.n552 B.n551 585
R1226 B.n553 B.n56 585
R1227 B.n555 B.n554 585
R1228 B.n556 B.n55 585
R1229 B.n558 B.n557 585
R1230 B.n559 B.n54 585
R1231 B.n561 B.n560 585
R1232 B.n562 B.n53 585
R1233 B.n564 B.n563 585
R1234 B.n566 B.n50 585
R1235 B.n568 B.n567 585
R1236 B.n569 B.n49 585
R1237 B.n571 B.n570 585
R1238 B.n572 B.n48 585
R1239 B.n574 B.n573 585
R1240 B.n575 B.n47 585
R1241 B.n577 B.n576 585
R1242 B.n578 B.n43 585
R1243 B.n580 B.n579 585
R1244 B.n581 B.n42 585
R1245 B.n583 B.n582 585
R1246 B.n584 B.n41 585
R1247 B.n586 B.n585 585
R1248 B.n587 B.n40 585
R1249 B.n589 B.n588 585
R1250 B.n590 B.n39 585
R1251 B.n592 B.n591 585
R1252 B.n593 B.n38 585
R1253 B.n595 B.n594 585
R1254 B.n596 B.n37 585
R1255 B.n598 B.n597 585
R1256 B.n599 B.n36 585
R1257 B.n601 B.n600 585
R1258 B.n602 B.n35 585
R1259 B.n604 B.n603 585
R1260 B.n605 B.n34 585
R1261 B.n607 B.n606 585
R1262 B.n608 B.n33 585
R1263 B.n610 B.n609 585
R1264 B.n611 B.n32 585
R1265 B.n613 B.n612 585
R1266 B.n614 B.n31 585
R1267 B.n616 B.n615 585
R1268 B.n617 B.n30 585
R1269 B.n619 B.n618 585
R1270 B.n620 B.n29 585
R1271 B.n622 B.n621 585
R1272 B.n623 B.n28 585
R1273 B.n625 B.n624 585
R1274 B.n626 B.n27 585
R1275 B.n628 B.n627 585
R1276 B.n629 B.n26 585
R1277 B.n631 B.n630 585
R1278 B.n632 B.n25 585
R1279 B.n634 B.n633 585
R1280 B.n635 B.n24 585
R1281 B.n637 B.n636 585
R1282 B.n638 B.n23 585
R1283 B.n640 B.n639 585
R1284 B.n641 B.n22 585
R1285 B.n643 B.n642 585
R1286 B.n644 B.n21 585
R1287 B.n646 B.n645 585
R1288 B.n647 B.n20 585
R1289 B.n649 B.n648 585
R1290 B.n650 B.n19 585
R1291 B.n652 B.n651 585
R1292 B.n653 B.n18 585
R1293 B.n655 B.n654 585
R1294 B.n656 B.n17 585
R1295 B.n658 B.n657 585
R1296 B.n659 B.n16 585
R1297 B.n661 B.n660 585
R1298 B.n662 B.n15 585
R1299 B.n664 B.n663 585
R1300 B.n480 B.n479 585
R1301 B.n478 B.n81 585
R1302 B.n477 B.n476 585
R1303 B.n475 B.n82 585
R1304 B.n474 B.n473 585
R1305 B.n472 B.n83 585
R1306 B.n471 B.n470 585
R1307 B.n469 B.n84 585
R1308 B.n468 B.n467 585
R1309 B.n466 B.n85 585
R1310 B.n465 B.n464 585
R1311 B.n463 B.n86 585
R1312 B.n462 B.n461 585
R1313 B.n460 B.n87 585
R1314 B.n459 B.n458 585
R1315 B.n457 B.n88 585
R1316 B.n456 B.n455 585
R1317 B.n454 B.n89 585
R1318 B.n453 B.n452 585
R1319 B.n451 B.n90 585
R1320 B.n450 B.n449 585
R1321 B.n448 B.n91 585
R1322 B.n447 B.n446 585
R1323 B.n445 B.n92 585
R1324 B.n444 B.n443 585
R1325 B.n442 B.n93 585
R1326 B.n441 B.n440 585
R1327 B.n439 B.n94 585
R1328 B.n438 B.n437 585
R1329 B.n436 B.n95 585
R1330 B.n435 B.n434 585
R1331 B.n433 B.n96 585
R1332 B.n432 B.n431 585
R1333 B.n430 B.n97 585
R1334 B.n429 B.n428 585
R1335 B.n427 B.n98 585
R1336 B.n426 B.n425 585
R1337 B.n424 B.n99 585
R1338 B.n423 B.n422 585
R1339 B.n421 B.n100 585
R1340 B.n420 B.n419 585
R1341 B.n418 B.n101 585
R1342 B.n417 B.n416 585
R1343 B.n415 B.n102 585
R1344 B.n414 B.n413 585
R1345 B.n412 B.n103 585
R1346 B.n411 B.n410 585
R1347 B.n409 B.n104 585
R1348 B.n408 B.n407 585
R1349 B.n406 B.n105 585
R1350 B.n405 B.n404 585
R1351 B.n220 B.n171 585
R1352 B.n222 B.n221 585
R1353 B.n223 B.n170 585
R1354 B.n225 B.n224 585
R1355 B.n226 B.n169 585
R1356 B.n228 B.n227 585
R1357 B.n229 B.n168 585
R1358 B.n231 B.n230 585
R1359 B.n232 B.n167 585
R1360 B.n234 B.n233 585
R1361 B.n235 B.n166 585
R1362 B.n237 B.n236 585
R1363 B.n238 B.n165 585
R1364 B.n240 B.n239 585
R1365 B.n241 B.n164 585
R1366 B.n243 B.n242 585
R1367 B.n244 B.n163 585
R1368 B.n246 B.n245 585
R1369 B.n247 B.n162 585
R1370 B.n249 B.n248 585
R1371 B.n250 B.n161 585
R1372 B.n252 B.n251 585
R1373 B.n253 B.n160 585
R1374 B.n255 B.n254 585
R1375 B.n256 B.n159 585
R1376 B.n258 B.n257 585
R1377 B.n259 B.n158 585
R1378 B.n261 B.n260 585
R1379 B.n262 B.n157 585
R1380 B.n264 B.n263 585
R1381 B.n265 B.n156 585
R1382 B.n267 B.n266 585
R1383 B.n268 B.n155 585
R1384 B.n270 B.n269 585
R1385 B.n271 B.n154 585
R1386 B.n273 B.n272 585
R1387 B.n274 B.n153 585
R1388 B.n276 B.n275 585
R1389 B.n277 B.n152 585
R1390 B.n279 B.n278 585
R1391 B.n280 B.n151 585
R1392 B.n282 B.n281 585
R1393 B.n283 B.n150 585
R1394 B.n285 B.n284 585
R1395 B.n286 B.n149 585
R1396 B.n288 B.n287 585
R1397 B.n289 B.n148 585
R1398 B.n291 B.n290 585
R1399 B.n292 B.n147 585
R1400 B.n294 B.n293 585
R1401 B.n295 B.n146 585
R1402 B.n297 B.n296 585
R1403 B.n298 B.n145 585
R1404 B.n300 B.n299 585
R1405 B.n301 B.n144 585
R1406 B.n303 B.n302 585
R1407 B.n305 B.n304 585
R1408 B.n306 B.n140 585
R1409 B.n308 B.n307 585
R1410 B.n309 B.n139 585
R1411 B.n311 B.n310 585
R1412 B.n312 B.n138 585
R1413 B.n314 B.n313 585
R1414 B.n315 B.n137 585
R1415 B.n317 B.n316 585
R1416 B.n318 B.n134 585
R1417 B.n321 B.n320 585
R1418 B.n322 B.n133 585
R1419 B.n324 B.n323 585
R1420 B.n325 B.n132 585
R1421 B.n327 B.n326 585
R1422 B.n328 B.n131 585
R1423 B.n330 B.n329 585
R1424 B.n331 B.n130 585
R1425 B.n333 B.n332 585
R1426 B.n334 B.n129 585
R1427 B.n336 B.n335 585
R1428 B.n337 B.n128 585
R1429 B.n339 B.n338 585
R1430 B.n340 B.n127 585
R1431 B.n342 B.n341 585
R1432 B.n343 B.n126 585
R1433 B.n345 B.n344 585
R1434 B.n346 B.n125 585
R1435 B.n348 B.n347 585
R1436 B.n349 B.n124 585
R1437 B.n351 B.n350 585
R1438 B.n352 B.n123 585
R1439 B.n354 B.n353 585
R1440 B.n355 B.n122 585
R1441 B.n357 B.n356 585
R1442 B.n358 B.n121 585
R1443 B.n360 B.n359 585
R1444 B.n361 B.n120 585
R1445 B.n363 B.n362 585
R1446 B.n364 B.n119 585
R1447 B.n366 B.n365 585
R1448 B.n367 B.n118 585
R1449 B.n369 B.n368 585
R1450 B.n370 B.n117 585
R1451 B.n372 B.n371 585
R1452 B.n373 B.n116 585
R1453 B.n375 B.n374 585
R1454 B.n376 B.n115 585
R1455 B.n378 B.n377 585
R1456 B.n379 B.n114 585
R1457 B.n381 B.n380 585
R1458 B.n382 B.n113 585
R1459 B.n384 B.n383 585
R1460 B.n385 B.n112 585
R1461 B.n387 B.n386 585
R1462 B.n388 B.n111 585
R1463 B.n390 B.n389 585
R1464 B.n391 B.n110 585
R1465 B.n393 B.n392 585
R1466 B.n394 B.n109 585
R1467 B.n396 B.n395 585
R1468 B.n397 B.n108 585
R1469 B.n399 B.n398 585
R1470 B.n400 B.n107 585
R1471 B.n402 B.n401 585
R1472 B.n403 B.n106 585
R1473 B.n219 B.n218 585
R1474 B.n217 B.n172 585
R1475 B.n216 B.n215 585
R1476 B.n214 B.n173 585
R1477 B.n213 B.n212 585
R1478 B.n211 B.n174 585
R1479 B.n210 B.n209 585
R1480 B.n208 B.n175 585
R1481 B.n207 B.n206 585
R1482 B.n205 B.n176 585
R1483 B.n204 B.n203 585
R1484 B.n202 B.n177 585
R1485 B.n201 B.n200 585
R1486 B.n199 B.n178 585
R1487 B.n198 B.n197 585
R1488 B.n196 B.n179 585
R1489 B.n195 B.n194 585
R1490 B.n193 B.n180 585
R1491 B.n192 B.n191 585
R1492 B.n190 B.n181 585
R1493 B.n189 B.n188 585
R1494 B.n187 B.n182 585
R1495 B.n186 B.n185 585
R1496 B.n184 B.n183 585
R1497 B.n2 B.n0 585
R1498 B.n701 B.n1 585
R1499 B.n700 B.n699 585
R1500 B.n698 B.n3 585
R1501 B.n697 B.n696 585
R1502 B.n695 B.n4 585
R1503 B.n694 B.n693 585
R1504 B.n692 B.n5 585
R1505 B.n691 B.n690 585
R1506 B.n689 B.n6 585
R1507 B.n688 B.n687 585
R1508 B.n686 B.n7 585
R1509 B.n685 B.n684 585
R1510 B.n683 B.n8 585
R1511 B.n682 B.n681 585
R1512 B.n680 B.n9 585
R1513 B.n679 B.n678 585
R1514 B.n677 B.n10 585
R1515 B.n676 B.n675 585
R1516 B.n674 B.n11 585
R1517 B.n673 B.n672 585
R1518 B.n671 B.n12 585
R1519 B.n670 B.n669 585
R1520 B.n668 B.n13 585
R1521 B.n667 B.n666 585
R1522 B.n665 B.n14 585
R1523 B.n703 B.n702 585
R1524 B.n135 B.t5 502.575
R1525 B.n51 B.t7 502.575
R1526 B.n141 B.t11 502.574
R1527 B.n44 B.t1 502.574
R1528 B.n220 B.n219 492.5
R1529 B.n665 B.n664 492.5
R1530 B.n405 B.n106 492.5
R1531 B.n479 B.n80 492.5
R1532 B.n135 B.t3 466.493
R1533 B.n141 B.t9 466.493
R1534 B.n44 B.t0 466.493
R1535 B.n51 B.t6 466.493
R1536 B.n136 B.t4 465.726
R1537 B.n52 B.t8 465.726
R1538 B.n142 B.t10 465.726
R1539 B.n45 B.t2 465.726
R1540 B.n219 B.n172 163.367
R1541 B.n215 B.n172 163.367
R1542 B.n215 B.n214 163.367
R1543 B.n214 B.n213 163.367
R1544 B.n213 B.n174 163.367
R1545 B.n209 B.n174 163.367
R1546 B.n209 B.n208 163.367
R1547 B.n208 B.n207 163.367
R1548 B.n207 B.n176 163.367
R1549 B.n203 B.n176 163.367
R1550 B.n203 B.n202 163.367
R1551 B.n202 B.n201 163.367
R1552 B.n201 B.n178 163.367
R1553 B.n197 B.n178 163.367
R1554 B.n197 B.n196 163.367
R1555 B.n196 B.n195 163.367
R1556 B.n195 B.n180 163.367
R1557 B.n191 B.n180 163.367
R1558 B.n191 B.n190 163.367
R1559 B.n190 B.n189 163.367
R1560 B.n189 B.n182 163.367
R1561 B.n185 B.n182 163.367
R1562 B.n185 B.n184 163.367
R1563 B.n184 B.n2 163.367
R1564 B.n702 B.n2 163.367
R1565 B.n702 B.n701 163.367
R1566 B.n701 B.n700 163.367
R1567 B.n700 B.n3 163.367
R1568 B.n696 B.n3 163.367
R1569 B.n696 B.n695 163.367
R1570 B.n695 B.n694 163.367
R1571 B.n694 B.n5 163.367
R1572 B.n690 B.n5 163.367
R1573 B.n690 B.n689 163.367
R1574 B.n689 B.n688 163.367
R1575 B.n688 B.n7 163.367
R1576 B.n684 B.n7 163.367
R1577 B.n684 B.n683 163.367
R1578 B.n683 B.n682 163.367
R1579 B.n682 B.n9 163.367
R1580 B.n678 B.n9 163.367
R1581 B.n678 B.n677 163.367
R1582 B.n677 B.n676 163.367
R1583 B.n676 B.n11 163.367
R1584 B.n672 B.n11 163.367
R1585 B.n672 B.n671 163.367
R1586 B.n671 B.n670 163.367
R1587 B.n670 B.n13 163.367
R1588 B.n666 B.n13 163.367
R1589 B.n666 B.n665 163.367
R1590 B.n221 B.n220 163.367
R1591 B.n221 B.n170 163.367
R1592 B.n225 B.n170 163.367
R1593 B.n226 B.n225 163.367
R1594 B.n227 B.n226 163.367
R1595 B.n227 B.n168 163.367
R1596 B.n231 B.n168 163.367
R1597 B.n232 B.n231 163.367
R1598 B.n233 B.n232 163.367
R1599 B.n233 B.n166 163.367
R1600 B.n237 B.n166 163.367
R1601 B.n238 B.n237 163.367
R1602 B.n239 B.n238 163.367
R1603 B.n239 B.n164 163.367
R1604 B.n243 B.n164 163.367
R1605 B.n244 B.n243 163.367
R1606 B.n245 B.n244 163.367
R1607 B.n245 B.n162 163.367
R1608 B.n249 B.n162 163.367
R1609 B.n250 B.n249 163.367
R1610 B.n251 B.n250 163.367
R1611 B.n251 B.n160 163.367
R1612 B.n255 B.n160 163.367
R1613 B.n256 B.n255 163.367
R1614 B.n257 B.n256 163.367
R1615 B.n257 B.n158 163.367
R1616 B.n261 B.n158 163.367
R1617 B.n262 B.n261 163.367
R1618 B.n263 B.n262 163.367
R1619 B.n263 B.n156 163.367
R1620 B.n267 B.n156 163.367
R1621 B.n268 B.n267 163.367
R1622 B.n269 B.n268 163.367
R1623 B.n269 B.n154 163.367
R1624 B.n273 B.n154 163.367
R1625 B.n274 B.n273 163.367
R1626 B.n275 B.n274 163.367
R1627 B.n275 B.n152 163.367
R1628 B.n279 B.n152 163.367
R1629 B.n280 B.n279 163.367
R1630 B.n281 B.n280 163.367
R1631 B.n281 B.n150 163.367
R1632 B.n285 B.n150 163.367
R1633 B.n286 B.n285 163.367
R1634 B.n287 B.n286 163.367
R1635 B.n287 B.n148 163.367
R1636 B.n291 B.n148 163.367
R1637 B.n292 B.n291 163.367
R1638 B.n293 B.n292 163.367
R1639 B.n293 B.n146 163.367
R1640 B.n297 B.n146 163.367
R1641 B.n298 B.n297 163.367
R1642 B.n299 B.n298 163.367
R1643 B.n299 B.n144 163.367
R1644 B.n303 B.n144 163.367
R1645 B.n304 B.n303 163.367
R1646 B.n304 B.n140 163.367
R1647 B.n308 B.n140 163.367
R1648 B.n309 B.n308 163.367
R1649 B.n310 B.n309 163.367
R1650 B.n310 B.n138 163.367
R1651 B.n314 B.n138 163.367
R1652 B.n315 B.n314 163.367
R1653 B.n316 B.n315 163.367
R1654 B.n316 B.n134 163.367
R1655 B.n321 B.n134 163.367
R1656 B.n322 B.n321 163.367
R1657 B.n323 B.n322 163.367
R1658 B.n323 B.n132 163.367
R1659 B.n327 B.n132 163.367
R1660 B.n328 B.n327 163.367
R1661 B.n329 B.n328 163.367
R1662 B.n329 B.n130 163.367
R1663 B.n333 B.n130 163.367
R1664 B.n334 B.n333 163.367
R1665 B.n335 B.n334 163.367
R1666 B.n335 B.n128 163.367
R1667 B.n339 B.n128 163.367
R1668 B.n340 B.n339 163.367
R1669 B.n341 B.n340 163.367
R1670 B.n341 B.n126 163.367
R1671 B.n345 B.n126 163.367
R1672 B.n346 B.n345 163.367
R1673 B.n347 B.n346 163.367
R1674 B.n347 B.n124 163.367
R1675 B.n351 B.n124 163.367
R1676 B.n352 B.n351 163.367
R1677 B.n353 B.n352 163.367
R1678 B.n353 B.n122 163.367
R1679 B.n357 B.n122 163.367
R1680 B.n358 B.n357 163.367
R1681 B.n359 B.n358 163.367
R1682 B.n359 B.n120 163.367
R1683 B.n363 B.n120 163.367
R1684 B.n364 B.n363 163.367
R1685 B.n365 B.n364 163.367
R1686 B.n365 B.n118 163.367
R1687 B.n369 B.n118 163.367
R1688 B.n370 B.n369 163.367
R1689 B.n371 B.n370 163.367
R1690 B.n371 B.n116 163.367
R1691 B.n375 B.n116 163.367
R1692 B.n376 B.n375 163.367
R1693 B.n377 B.n376 163.367
R1694 B.n377 B.n114 163.367
R1695 B.n381 B.n114 163.367
R1696 B.n382 B.n381 163.367
R1697 B.n383 B.n382 163.367
R1698 B.n383 B.n112 163.367
R1699 B.n387 B.n112 163.367
R1700 B.n388 B.n387 163.367
R1701 B.n389 B.n388 163.367
R1702 B.n389 B.n110 163.367
R1703 B.n393 B.n110 163.367
R1704 B.n394 B.n393 163.367
R1705 B.n395 B.n394 163.367
R1706 B.n395 B.n108 163.367
R1707 B.n399 B.n108 163.367
R1708 B.n400 B.n399 163.367
R1709 B.n401 B.n400 163.367
R1710 B.n401 B.n106 163.367
R1711 B.n406 B.n405 163.367
R1712 B.n407 B.n406 163.367
R1713 B.n407 B.n104 163.367
R1714 B.n411 B.n104 163.367
R1715 B.n412 B.n411 163.367
R1716 B.n413 B.n412 163.367
R1717 B.n413 B.n102 163.367
R1718 B.n417 B.n102 163.367
R1719 B.n418 B.n417 163.367
R1720 B.n419 B.n418 163.367
R1721 B.n419 B.n100 163.367
R1722 B.n423 B.n100 163.367
R1723 B.n424 B.n423 163.367
R1724 B.n425 B.n424 163.367
R1725 B.n425 B.n98 163.367
R1726 B.n429 B.n98 163.367
R1727 B.n430 B.n429 163.367
R1728 B.n431 B.n430 163.367
R1729 B.n431 B.n96 163.367
R1730 B.n435 B.n96 163.367
R1731 B.n436 B.n435 163.367
R1732 B.n437 B.n436 163.367
R1733 B.n437 B.n94 163.367
R1734 B.n441 B.n94 163.367
R1735 B.n442 B.n441 163.367
R1736 B.n443 B.n442 163.367
R1737 B.n443 B.n92 163.367
R1738 B.n447 B.n92 163.367
R1739 B.n448 B.n447 163.367
R1740 B.n449 B.n448 163.367
R1741 B.n449 B.n90 163.367
R1742 B.n453 B.n90 163.367
R1743 B.n454 B.n453 163.367
R1744 B.n455 B.n454 163.367
R1745 B.n455 B.n88 163.367
R1746 B.n459 B.n88 163.367
R1747 B.n460 B.n459 163.367
R1748 B.n461 B.n460 163.367
R1749 B.n461 B.n86 163.367
R1750 B.n465 B.n86 163.367
R1751 B.n466 B.n465 163.367
R1752 B.n467 B.n466 163.367
R1753 B.n467 B.n84 163.367
R1754 B.n471 B.n84 163.367
R1755 B.n472 B.n471 163.367
R1756 B.n473 B.n472 163.367
R1757 B.n473 B.n82 163.367
R1758 B.n477 B.n82 163.367
R1759 B.n478 B.n477 163.367
R1760 B.n479 B.n478 163.367
R1761 B.n664 B.n15 163.367
R1762 B.n660 B.n15 163.367
R1763 B.n660 B.n659 163.367
R1764 B.n659 B.n658 163.367
R1765 B.n658 B.n17 163.367
R1766 B.n654 B.n17 163.367
R1767 B.n654 B.n653 163.367
R1768 B.n653 B.n652 163.367
R1769 B.n652 B.n19 163.367
R1770 B.n648 B.n19 163.367
R1771 B.n648 B.n647 163.367
R1772 B.n647 B.n646 163.367
R1773 B.n646 B.n21 163.367
R1774 B.n642 B.n21 163.367
R1775 B.n642 B.n641 163.367
R1776 B.n641 B.n640 163.367
R1777 B.n640 B.n23 163.367
R1778 B.n636 B.n23 163.367
R1779 B.n636 B.n635 163.367
R1780 B.n635 B.n634 163.367
R1781 B.n634 B.n25 163.367
R1782 B.n630 B.n25 163.367
R1783 B.n630 B.n629 163.367
R1784 B.n629 B.n628 163.367
R1785 B.n628 B.n27 163.367
R1786 B.n624 B.n27 163.367
R1787 B.n624 B.n623 163.367
R1788 B.n623 B.n622 163.367
R1789 B.n622 B.n29 163.367
R1790 B.n618 B.n29 163.367
R1791 B.n618 B.n617 163.367
R1792 B.n617 B.n616 163.367
R1793 B.n616 B.n31 163.367
R1794 B.n612 B.n31 163.367
R1795 B.n612 B.n611 163.367
R1796 B.n611 B.n610 163.367
R1797 B.n610 B.n33 163.367
R1798 B.n606 B.n33 163.367
R1799 B.n606 B.n605 163.367
R1800 B.n605 B.n604 163.367
R1801 B.n604 B.n35 163.367
R1802 B.n600 B.n35 163.367
R1803 B.n600 B.n599 163.367
R1804 B.n599 B.n598 163.367
R1805 B.n598 B.n37 163.367
R1806 B.n594 B.n37 163.367
R1807 B.n594 B.n593 163.367
R1808 B.n593 B.n592 163.367
R1809 B.n592 B.n39 163.367
R1810 B.n588 B.n39 163.367
R1811 B.n588 B.n587 163.367
R1812 B.n587 B.n586 163.367
R1813 B.n586 B.n41 163.367
R1814 B.n582 B.n41 163.367
R1815 B.n582 B.n581 163.367
R1816 B.n581 B.n580 163.367
R1817 B.n580 B.n43 163.367
R1818 B.n576 B.n43 163.367
R1819 B.n576 B.n575 163.367
R1820 B.n575 B.n574 163.367
R1821 B.n574 B.n48 163.367
R1822 B.n570 B.n48 163.367
R1823 B.n570 B.n569 163.367
R1824 B.n569 B.n568 163.367
R1825 B.n568 B.n50 163.367
R1826 B.n563 B.n50 163.367
R1827 B.n563 B.n562 163.367
R1828 B.n562 B.n561 163.367
R1829 B.n561 B.n54 163.367
R1830 B.n557 B.n54 163.367
R1831 B.n557 B.n556 163.367
R1832 B.n556 B.n555 163.367
R1833 B.n555 B.n56 163.367
R1834 B.n551 B.n56 163.367
R1835 B.n551 B.n550 163.367
R1836 B.n550 B.n549 163.367
R1837 B.n549 B.n58 163.367
R1838 B.n545 B.n58 163.367
R1839 B.n545 B.n544 163.367
R1840 B.n544 B.n543 163.367
R1841 B.n543 B.n60 163.367
R1842 B.n539 B.n60 163.367
R1843 B.n539 B.n538 163.367
R1844 B.n538 B.n537 163.367
R1845 B.n537 B.n62 163.367
R1846 B.n533 B.n62 163.367
R1847 B.n533 B.n532 163.367
R1848 B.n532 B.n531 163.367
R1849 B.n531 B.n64 163.367
R1850 B.n527 B.n64 163.367
R1851 B.n527 B.n526 163.367
R1852 B.n526 B.n525 163.367
R1853 B.n525 B.n66 163.367
R1854 B.n521 B.n66 163.367
R1855 B.n521 B.n520 163.367
R1856 B.n520 B.n519 163.367
R1857 B.n519 B.n68 163.367
R1858 B.n515 B.n68 163.367
R1859 B.n515 B.n514 163.367
R1860 B.n514 B.n513 163.367
R1861 B.n513 B.n70 163.367
R1862 B.n509 B.n70 163.367
R1863 B.n509 B.n508 163.367
R1864 B.n508 B.n507 163.367
R1865 B.n507 B.n72 163.367
R1866 B.n503 B.n72 163.367
R1867 B.n503 B.n502 163.367
R1868 B.n502 B.n501 163.367
R1869 B.n501 B.n74 163.367
R1870 B.n497 B.n74 163.367
R1871 B.n497 B.n496 163.367
R1872 B.n496 B.n495 163.367
R1873 B.n495 B.n76 163.367
R1874 B.n491 B.n76 163.367
R1875 B.n491 B.n490 163.367
R1876 B.n490 B.n489 163.367
R1877 B.n489 B.n78 163.367
R1878 B.n485 B.n78 163.367
R1879 B.n485 B.n484 163.367
R1880 B.n484 B.n483 163.367
R1881 B.n483 B.n80 163.367
R1882 B.n319 B.n136 59.5399
R1883 B.n143 B.n142 59.5399
R1884 B.n46 B.n45 59.5399
R1885 B.n565 B.n52 59.5399
R1886 B.n136 B.n135 36.849
R1887 B.n142 B.n141 36.849
R1888 B.n45 B.n44 36.849
R1889 B.n52 B.n51 36.849
R1890 B.n663 B.n14 32.0005
R1891 B.n481 B.n480 32.0005
R1892 B.n404 B.n403 32.0005
R1893 B.n218 B.n171 32.0005
R1894 B B.n703 18.0485
R1895 B.n663 B.n662 10.6151
R1896 B.n662 B.n661 10.6151
R1897 B.n661 B.n16 10.6151
R1898 B.n657 B.n16 10.6151
R1899 B.n657 B.n656 10.6151
R1900 B.n656 B.n655 10.6151
R1901 B.n655 B.n18 10.6151
R1902 B.n651 B.n18 10.6151
R1903 B.n651 B.n650 10.6151
R1904 B.n650 B.n649 10.6151
R1905 B.n649 B.n20 10.6151
R1906 B.n645 B.n20 10.6151
R1907 B.n645 B.n644 10.6151
R1908 B.n644 B.n643 10.6151
R1909 B.n643 B.n22 10.6151
R1910 B.n639 B.n22 10.6151
R1911 B.n639 B.n638 10.6151
R1912 B.n638 B.n637 10.6151
R1913 B.n637 B.n24 10.6151
R1914 B.n633 B.n24 10.6151
R1915 B.n633 B.n632 10.6151
R1916 B.n632 B.n631 10.6151
R1917 B.n631 B.n26 10.6151
R1918 B.n627 B.n26 10.6151
R1919 B.n627 B.n626 10.6151
R1920 B.n626 B.n625 10.6151
R1921 B.n625 B.n28 10.6151
R1922 B.n621 B.n28 10.6151
R1923 B.n621 B.n620 10.6151
R1924 B.n620 B.n619 10.6151
R1925 B.n619 B.n30 10.6151
R1926 B.n615 B.n30 10.6151
R1927 B.n615 B.n614 10.6151
R1928 B.n614 B.n613 10.6151
R1929 B.n613 B.n32 10.6151
R1930 B.n609 B.n32 10.6151
R1931 B.n609 B.n608 10.6151
R1932 B.n608 B.n607 10.6151
R1933 B.n607 B.n34 10.6151
R1934 B.n603 B.n34 10.6151
R1935 B.n603 B.n602 10.6151
R1936 B.n602 B.n601 10.6151
R1937 B.n601 B.n36 10.6151
R1938 B.n597 B.n36 10.6151
R1939 B.n597 B.n596 10.6151
R1940 B.n596 B.n595 10.6151
R1941 B.n595 B.n38 10.6151
R1942 B.n591 B.n38 10.6151
R1943 B.n591 B.n590 10.6151
R1944 B.n590 B.n589 10.6151
R1945 B.n589 B.n40 10.6151
R1946 B.n585 B.n40 10.6151
R1947 B.n585 B.n584 10.6151
R1948 B.n584 B.n583 10.6151
R1949 B.n583 B.n42 10.6151
R1950 B.n579 B.n578 10.6151
R1951 B.n578 B.n577 10.6151
R1952 B.n577 B.n47 10.6151
R1953 B.n573 B.n47 10.6151
R1954 B.n573 B.n572 10.6151
R1955 B.n572 B.n571 10.6151
R1956 B.n571 B.n49 10.6151
R1957 B.n567 B.n49 10.6151
R1958 B.n567 B.n566 10.6151
R1959 B.n564 B.n53 10.6151
R1960 B.n560 B.n53 10.6151
R1961 B.n560 B.n559 10.6151
R1962 B.n559 B.n558 10.6151
R1963 B.n558 B.n55 10.6151
R1964 B.n554 B.n55 10.6151
R1965 B.n554 B.n553 10.6151
R1966 B.n553 B.n552 10.6151
R1967 B.n552 B.n57 10.6151
R1968 B.n548 B.n57 10.6151
R1969 B.n548 B.n547 10.6151
R1970 B.n547 B.n546 10.6151
R1971 B.n546 B.n59 10.6151
R1972 B.n542 B.n59 10.6151
R1973 B.n542 B.n541 10.6151
R1974 B.n541 B.n540 10.6151
R1975 B.n540 B.n61 10.6151
R1976 B.n536 B.n61 10.6151
R1977 B.n536 B.n535 10.6151
R1978 B.n535 B.n534 10.6151
R1979 B.n534 B.n63 10.6151
R1980 B.n530 B.n63 10.6151
R1981 B.n530 B.n529 10.6151
R1982 B.n529 B.n528 10.6151
R1983 B.n528 B.n65 10.6151
R1984 B.n524 B.n65 10.6151
R1985 B.n524 B.n523 10.6151
R1986 B.n523 B.n522 10.6151
R1987 B.n522 B.n67 10.6151
R1988 B.n518 B.n67 10.6151
R1989 B.n518 B.n517 10.6151
R1990 B.n517 B.n516 10.6151
R1991 B.n516 B.n69 10.6151
R1992 B.n512 B.n69 10.6151
R1993 B.n512 B.n511 10.6151
R1994 B.n511 B.n510 10.6151
R1995 B.n510 B.n71 10.6151
R1996 B.n506 B.n71 10.6151
R1997 B.n506 B.n505 10.6151
R1998 B.n505 B.n504 10.6151
R1999 B.n504 B.n73 10.6151
R2000 B.n500 B.n73 10.6151
R2001 B.n500 B.n499 10.6151
R2002 B.n499 B.n498 10.6151
R2003 B.n498 B.n75 10.6151
R2004 B.n494 B.n75 10.6151
R2005 B.n494 B.n493 10.6151
R2006 B.n493 B.n492 10.6151
R2007 B.n492 B.n77 10.6151
R2008 B.n488 B.n77 10.6151
R2009 B.n488 B.n487 10.6151
R2010 B.n487 B.n486 10.6151
R2011 B.n486 B.n79 10.6151
R2012 B.n482 B.n79 10.6151
R2013 B.n482 B.n481 10.6151
R2014 B.n404 B.n105 10.6151
R2015 B.n408 B.n105 10.6151
R2016 B.n409 B.n408 10.6151
R2017 B.n410 B.n409 10.6151
R2018 B.n410 B.n103 10.6151
R2019 B.n414 B.n103 10.6151
R2020 B.n415 B.n414 10.6151
R2021 B.n416 B.n415 10.6151
R2022 B.n416 B.n101 10.6151
R2023 B.n420 B.n101 10.6151
R2024 B.n421 B.n420 10.6151
R2025 B.n422 B.n421 10.6151
R2026 B.n422 B.n99 10.6151
R2027 B.n426 B.n99 10.6151
R2028 B.n427 B.n426 10.6151
R2029 B.n428 B.n427 10.6151
R2030 B.n428 B.n97 10.6151
R2031 B.n432 B.n97 10.6151
R2032 B.n433 B.n432 10.6151
R2033 B.n434 B.n433 10.6151
R2034 B.n434 B.n95 10.6151
R2035 B.n438 B.n95 10.6151
R2036 B.n439 B.n438 10.6151
R2037 B.n440 B.n439 10.6151
R2038 B.n440 B.n93 10.6151
R2039 B.n444 B.n93 10.6151
R2040 B.n445 B.n444 10.6151
R2041 B.n446 B.n445 10.6151
R2042 B.n446 B.n91 10.6151
R2043 B.n450 B.n91 10.6151
R2044 B.n451 B.n450 10.6151
R2045 B.n452 B.n451 10.6151
R2046 B.n452 B.n89 10.6151
R2047 B.n456 B.n89 10.6151
R2048 B.n457 B.n456 10.6151
R2049 B.n458 B.n457 10.6151
R2050 B.n458 B.n87 10.6151
R2051 B.n462 B.n87 10.6151
R2052 B.n463 B.n462 10.6151
R2053 B.n464 B.n463 10.6151
R2054 B.n464 B.n85 10.6151
R2055 B.n468 B.n85 10.6151
R2056 B.n469 B.n468 10.6151
R2057 B.n470 B.n469 10.6151
R2058 B.n470 B.n83 10.6151
R2059 B.n474 B.n83 10.6151
R2060 B.n475 B.n474 10.6151
R2061 B.n476 B.n475 10.6151
R2062 B.n476 B.n81 10.6151
R2063 B.n480 B.n81 10.6151
R2064 B.n222 B.n171 10.6151
R2065 B.n223 B.n222 10.6151
R2066 B.n224 B.n223 10.6151
R2067 B.n224 B.n169 10.6151
R2068 B.n228 B.n169 10.6151
R2069 B.n229 B.n228 10.6151
R2070 B.n230 B.n229 10.6151
R2071 B.n230 B.n167 10.6151
R2072 B.n234 B.n167 10.6151
R2073 B.n235 B.n234 10.6151
R2074 B.n236 B.n235 10.6151
R2075 B.n236 B.n165 10.6151
R2076 B.n240 B.n165 10.6151
R2077 B.n241 B.n240 10.6151
R2078 B.n242 B.n241 10.6151
R2079 B.n242 B.n163 10.6151
R2080 B.n246 B.n163 10.6151
R2081 B.n247 B.n246 10.6151
R2082 B.n248 B.n247 10.6151
R2083 B.n248 B.n161 10.6151
R2084 B.n252 B.n161 10.6151
R2085 B.n253 B.n252 10.6151
R2086 B.n254 B.n253 10.6151
R2087 B.n254 B.n159 10.6151
R2088 B.n258 B.n159 10.6151
R2089 B.n259 B.n258 10.6151
R2090 B.n260 B.n259 10.6151
R2091 B.n260 B.n157 10.6151
R2092 B.n264 B.n157 10.6151
R2093 B.n265 B.n264 10.6151
R2094 B.n266 B.n265 10.6151
R2095 B.n266 B.n155 10.6151
R2096 B.n270 B.n155 10.6151
R2097 B.n271 B.n270 10.6151
R2098 B.n272 B.n271 10.6151
R2099 B.n272 B.n153 10.6151
R2100 B.n276 B.n153 10.6151
R2101 B.n277 B.n276 10.6151
R2102 B.n278 B.n277 10.6151
R2103 B.n278 B.n151 10.6151
R2104 B.n282 B.n151 10.6151
R2105 B.n283 B.n282 10.6151
R2106 B.n284 B.n283 10.6151
R2107 B.n284 B.n149 10.6151
R2108 B.n288 B.n149 10.6151
R2109 B.n289 B.n288 10.6151
R2110 B.n290 B.n289 10.6151
R2111 B.n290 B.n147 10.6151
R2112 B.n294 B.n147 10.6151
R2113 B.n295 B.n294 10.6151
R2114 B.n296 B.n295 10.6151
R2115 B.n296 B.n145 10.6151
R2116 B.n300 B.n145 10.6151
R2117 B.n301 B.n300 10.6151
R2118 B.n302 B.n301 10.6151
R2119 B.n306 B.n305 10.6151
R2120 B.n307 B.n306 10.6151
R2121 B.n307 B.n139 10.6151
R2122 B.n311 B.n139 10.6151
R2123 B.n312 B.n311 10.6151
R2124 B.n313 B.n312 10.6151
R2125 B.n313 B.n137 10.6151
R2126 B.n317 B.n137 10.6151
R2127 B.n318 B.n317 10.6151
R2128 B.n320 B.n133 10.6151
R2129 B.n324 B.n133 10.6151
R2130 B.n325 B.n324 10.6151
R2131 B.n326 B.n325 10.6151
R2132 B.n326 B.n131 10.6151
R2133 B.n330 B.n131 10.6151
R2134 B.n331 B.n330 10.6151
R2135 B.n332 B.n331 10.6151
R2136 B.n332 B.n129 10.6151
R2137 B.n336 B.n129 10.6151
R2138 B.n337 B.n336 10.6151
R2139 B.n338 B.n337 10.6151
R2140 B.n338 B.n127 10.6151
R2141 B.n342 B.n127 10.6151
R2142 B.n343 B.n342 10.6151
R2143 B.n344 B.n343 10.6151
R2144 B.n344 B.n125 10.6151
R2145 B.n348 B.n125 10.6151
R2146 B.n349 B.n348 10.6151
R2147 B.n350 B.n349 10.6151
R2148 B.n350 B.n123 10.6151
R2149 B.n354 B.n123 10.6151
R2150 B.n355 B.n354 10.6151
R2151 B.n356 B.n355 10.6151
R2152 B.n356 B.n121 10.6151
R2153 B.n360 B.n121 10.6151
R2154 B.n361 B.n360 10.6151
R2155 B.n362 B.n361 10.6151
R2156 B.n362 B.n119 10.6151
R2157 B.n366 B.n119 10.6151
R2158 B.n367 B.n366 10.6151
R2159 B.n368 B.n367 10.6151
R2160 B.n368 B.n117 10.6151
R2161 B.n372 B.n117 10.6151
R2162 B.n373 B.n372 10.6151
R2163 B.n374 B.n373 10.6151
R2164 B.n374 B.n115 10.6151
R2165 B.n378 B.n115 10.6151
R2166 B.n379 B.n378 10.6151
R2167 B.n380 B.n379 10.6151
R2168 B.n380 B.n113 10.6151
R2169 B.n384 B.n113 10.6151
R2170 B.n385 B.n384 10.6151
R2171 B.n386 B.n385 10.6151
R2172 B.n386 B.n111 10.6151
R2173 B.n390 B.n111 10.6151
R2174 B.n391 B.n390 10.6151
R2175 B.n392 B.n391 10.6151
R2176 B.n392 B.n109 10.6151
R2177 B.n396 B.n109 10.6151
R2178 B.n397 B.n396 10.6151
R2179 B.n398 B.n397 10.6151
R2180 B.n398 B.n107 10.6151
R2181 B.n402 B.n107 10.6151
R2182 B.n403 B.n402 10.6151
R2183 B.n218 B.n217 10.6151
R2184 B.n217 B.n216 10.6151
R2185 B.n216 B.n173 10.6151
R2186 B.n212 B.n173 10.6151
R2187 B.n212 B.n211 10.6151
R2188 B.n211 B.n210 10.6151
R2189 B.n210 B.n175 10.6151
R2190 B.n206 B.n175 10.6151
R2191 B.n206 B.n205 10.6151
R2192 B.n205 B.n204 10.6151
R2193 B.n204 B.n177 10.6151
R2194 B.n200 B.n177 10.6151
R2195 B.n200 B.n199 10.6151
R2196 B.n199 B.n198 10.6151
R2197 B.n198 B.n179 10.6151
R2198 B.n194 B.n179 10.6151
R2199 B.n194 B.n193 10.6151
R2200 B.n193 B.n192 10.6151
R2201 B.n192 B.n181 10.6151
R2202 B.n188 B.n181 10.6151
R2203 B.n188 B.n187 10.6151
R2204 B.n187 B.n186 10.6151
R2205 B.n186 B.n183 10.6151
R2206 B.n183 B.n0 10.6151
R2207 B.n699 B.n1 10.6151
R2208 B.n699 B.n698 10.6151
R2209 B.n698 B.n697 10.6151
R2210 B.n697 B.n4 10.6151
R2211 B.n693 B.n4 10.6151
R2212 B.n693 B.n692 10.6151
R2213 B.n692 B.n691 10.6151
R2214 B.n691 B.n6 10.6151
R2215 B.n687 B.n6 10.6151
R2216 B.n687 B.n686 10.6151
R2217 B.n686 B.n685 10.6151
R2218 B.n685 B.n8 10.6151
R2219 B.n681 B.n8 10.6151
R2220 B.n681 B.n680 10.6151
R2221 B.n680 B.n679 10.6151
R2222 B.n679 B.n10 10.6151
R2223 B.n675 B.n10 10.6151
R2224 B.n675 B.n674 10.6151
R2225 B.n674 B.n673 10.6151
R2226 B.n673 B.n12 10.6151
R2227 B.n669 B.n12 10.6151
R2228 B.n669 B.n668 10.6151
R2229 B.n668 B.n667 10.6151
R2230 B.n667 B.n14 10.6151
R2231 B.n46 B.n42 9.36635
R2232 B.n565 B.n564 9.36635
R2233 B.n302 B.n143 9.36635
R2234 B.n320 B.n319 9.36635
R2235 B.n703 B.n0 2.81026
R2236 B.n703 B.n1 2.81026
R2237 B.n579 B.n46 1.24928
R2238 B.n566 B.n565 1.24928
R2239 B.n305 B.n143 1.24928
R2240 B.n319 B.n318 1.24928
C0 VDD2 VP 0.328884f
C1 w_n2110_n4366# B 9.37739f
C2 VP VN 6.37152f
C3 VDD2 B 1.25028f
C4 B VN 0.971771f
C5 VDD1 VP 6.05497f
C6 VDD1 B 1.21495f
C7 B VP 1.41278f
C8 VTAIL w_n2110_n4366# 5.18417f
C9 VTAIL VDD2 7.01573f
C10 VTAIL VN 5.43108f
C11 VDD2 w_n2110_n4366# 1.41896f
C12 VTAIL VDD1 6.96842f
C13 w_n2110_n4366# VN 3.47168f
C14 VDD2 VN 5.87475f
C15 VDD1 w_n2110_n4366# 1.38588f
C16 VDD1 VDD2 0.776947f
C17 VDD1 VN 0.148188f
C18 VTAIL VP 5.44518f
C19 VTAIL B 5.9285f
C20 w_n2110_n4366# VP 3.74033f
C21 VDD2 VSUBS 0.910093f
C22 VDD1 VSUBS 5.885f
C23 VTAIL VSUBS 1.296889f
C24 VN VSUBS 5.46432f
C25 VP VSUBS 1.91967f
C26 B VSUBS 3.807018f
C27 w_n2110_n4366# VSUBS 0.11275p
C28 B.n0 VSUBS 0.00435f
C29 B.n1 VSUBS 0.00435f
C30 B.n2 VSUBS 0.006879f
C31 B.n3 VSUBS 0.006879f
C32 B.n4 VSUBS 0.006879f
C33 B.n5 VSUBS 0.006879f
C34 B.n6 VSUBS 0.006879f
C35 B.n7 VSUBS 0.006879f
C36 B.n8 VSUBS 0.006879f
C37 B.n9 VSUBS 0.006879f
C38 B.n10 VSUBS 0.006879f
C39 B.n11 VSUBS 0.006879f
C40 B.n12 VSUBS 0.006879f
C41 B.n13 VSUBS 0.006879f
C42 B.n14 VSUBS 0.01563f
C43 B.n15 VSUBS 0.006879f
C44 B.n16 VSUBS 0.006879f
C45 B.n17 VSUBS 0.006879f
C46 B.n18 VSUBS 0.006879f
C47 B.n19 VSUBS 0.006879f
C48 B.n20 VSUBS 0.006879f
C49 B.n21 VSUBS 0.006879f
C50 B.n22 VSUBS 0.006879f
C51 B.n23 VSUBS 0.006879f
C52 B.n24 VSUBS 0.006879f
C53 B.n25 VSUBS 0.006879f
C54 B.n26 VSUBS 0.006879f
C55 B.n27 VSUBS 0.006879f
C56 B.n28 VSUBS 0.006879f
C57 B.n29 VSUBS 0.006879f
C58 B.n30 VSUBS 0.006879f
C59 B.n31 VSUBS 0.006879f
C60 B.n32 VSUBS 0.006879f
C61 B.n33 VSUBS 0.006879f
C62 B.n34 VSUBS 0.006879f
C63 B.n35 VSUBS 0.006879f
C64 B.n36 VSUBS 0.006879f
C65 B.n37 VSUBS 0.006879f
C66 B.n38 VSUBS 0.006879f
C67 B.n39 VSUBS 0.006879f
C68 B.n40 VSUBS 0.006879f
C69 B.n41 VSUBS 0.006879f
C70 B.n42 VSUBS 0.006474f
C71 B.n43 VSUBS 0.006879f
C72 B.t2 VSUBS 0.321354f
C73 B.t1 VSUBS 0.343116f
C74 B.t0 VSUBS 1.12314f
C75 B.n44 VSUBS 0.489086f
C76 B.n45 VSUBS 0.306619f
C77 B.n46 VSUBS 0.015938f
C78 B.n47 VSUBS 0.006879f
C79 B.n48 VSUBS 0.006879f
C80 B.n49 VSUBS 0.006879f
C81 B.n50 VSUBS 0.006879f
C82 B.t8 VSUBS 0.321357f
C83 B.t7 VSUBS 0.343119f
C84 B.t6 VSUBS 1.12314f
C85 B.n51 VSUBS 0.489082f
C86 B.n52 VSUBS 0.306616f
C87 B.n53 VSUBS 0.006879f
C88 B.n54 VSUBS 0.006879f
C89 B.n55 VSUBS 0.006879f
C90 B.n56 VSUBS 0.006879f
C91 B.n57 VSUBS 0.006879f
C92 B.n58 VSUBS 0.006879f
C93 B.n59 VSUBS 0.006879f
C94 B.n60 VSUBS 0.006879f
C95 B.n61 VSUBS 0.006879f
C96 B.n62 VSUBS 0.006879f
C97 B.n63 VSUBS 0.006879f
C98 B.n64 VSUBS 0.006879f
C99 B.n65 VSUBS 0.006879f
C100 B.n66 VSUBS 0.006879f
C101 B.n67 VSUBS 0.006879f
C102 B.n68 VSUBS 0.006879f
C103 B.n69 VSUBS 0.006879f
C104 B.n70 VSUBS 0.006879f
C105 B.n71 VSUBS 0.006879f
C106 B.n72 VSUBS 0.006879f
C107 B.n73 VSUBS 0.006879f
C108 B.n74 VSUBS 0.006879f
C109 B.n75 VSUBS 0.006879f
C110 B.n76 VSUBS 0.006879f
C111 B.n77 VSUBS 0.006879f
C112 B.n78 VSUBS 0.006879f
C113 B.n79 VSUBS 0.006879f
C114 B.n80 VSUBS 0.016136f
C115 B.n81 VSUBS 0.006879f
C116 B.n82 VSUBS 0.006879f
C117 B.n83 VSUBS 0.006879f
C118 B.n84 VSUBS 0.006879f
C119 B.n85 VSUBS 0.006879f
C120 B.n86 VSUBS 0.006879f
C121 B.n87 VSUBS 0.006879f
C122 B.n88 VSUBS 0.006879f
C123 B.n89 VSUBS 0.006879f
C124 B.n90 VSUBS 0.006879f
C125 B.n91 VSUBS 0.006879f
C126 B.n92 VSUBS 0.006879f
C127 B.n93 VSUBS 0.006879f
C128 B.n94 VSUBS 0.006879f
C129 B.n95 VSUBS 0.006879f
C130 B.n96 VSUBS 0.006879f
C131 B.n97 VSUBS 0.006879f
C132 B.n98 VSUBS 0.006879f
C133 B.n99 VSUBS 0.006879f
C134 B.n100 VSUBS 0.006879f
C135 B.n101 VSUBS 0.006879f
C136 B.n102 VSUBS 0.006879f
C137 B.n103 VSUBS 0.006879f
C138 B.n104 VSUBS 0.006879f
C139 B.n105 VSUBS 0.006879f
C140 B.n106 VSUBS 0.016136f
C141 B.n107 VSUBS 0.006879f
C142 B.n108 VSUBS 0.006879f
C143 B.n109 VSUBS 0.006879f
C144 B.n110 VSUBS 0.006879f
C145 B.n111 VSUBS 0.006879f
C146 B.n112 VSUBS 0.006879f
C147 B.n113 VSUBS 0.006879f
C148 B.n114 VSUBS 0.006879f
C149 B.n115 VSUBS 0.006879f
C150 B.n116 VSUBS 0.006879f
C151 B.n117 VSUBS 0.006879f
C152 B.n118 VSUBS 0.006879f
C153 B.n119 VSUBS 0.006879f
C154 B.n120 VSUBS 0.006879f
C155 B.n121 VSUBS 0.006879f
C156 B.n122 VSUBS 0.006879f
C157 B.n123 VSUBS 0.006879f
C158 B.n124 VSUBS 0.006879f
C159 B.n125 VSUBS 0.006879f
C160 B.n126 VSUBS 0.006879f
C161 B.n127 VSUBS 0.006879f
C162 B.n128 VSUBS 0.006879f
C163 B.n129 VSUBS 0.006879f
C164 B.n130 VSUBS 0.006879f
C165 B.n131 VSUBS 0.006879f
C166 B.n132 VSUBS 0.006879f
C167 B.n133 VSUBS 0.006879f
C168 B.n134 VSUBS 0.006879f
C169 B.t4 VSUBS 0.321357f
C170 B.t5 VSUBS 0.343119f
C171 B.t3 VSUBS 1.12314f
C172 B.n135 VSUBS 0.489082f
C173 B.n136 VSUBS 0.306616f
C174 B.n137 VSUBS 0.006879f
C175 B.n138 VSUBS 0.006879f
C176 B.n139 VSUBS 0.006879f
C177 B.n140 VSUBS 0.006879f
C178 B.t10 VSUBS 0.321354f
C179 B.t11 VSUBS 0.343116f
C180 B.t9 VSUBS 1.12314f
C181 B.n141 VSUBS 0.489086f
C182 B.n142 VSUBS 0.306619f
C183 B.n143 VSUBS 0.015938f
C184 B.n144 VSUBS 0.006879f
C185 B.n145 VSUBS 0.006879f
C186 B.n146 VSUBS 0.006879f
C187 B.n147 VSUBS 0.006879f
C188 B.n148 VSUBS 0.006879f
C189 B.n149 VSUBS 0.006879f
C190 B.n150 VSUBS 0.006879f
C191 B.n151 VSUBS 0.006879f
C192 B.n152 VSUBS 0.006879f
C193 B.n153 VSUBS 0.006879f
C194 B.n154 VSUBS 0.006879f
C195 B.n155 VSUBS 0.006879f
C196 B.n156 VSUBS 0.006879f
C197 B.n157 VSUBS 0.006879f
C198 B.n158 VSUBS 0.006879f
C199 B.n159 VSUBS 0.006879f
C200 B.n160 VSUBS 0.006879f
C201 B.n161 VSUBS 0.006879f
C202 B.n162 VSUBS 0.006879f
C203 B.n163 VSUBS 0.006879f
C204 B.n164 VSUBS 0.006879f
C205 B.n165 VSUBS 0.006879f
C206 B.n166 VSUBS 0.006879f
C207 B.n167 VSUBS 0.006879f
C208 B.n168 VSUBS 0.006879f
C209 B.n169 VSUBS 0.006879f
C210 B.n170 VSUBS 0.006879f
C211 B.n171 VSUBS 0.016136f
C212 B.n172 VSUBS 0.006879f
C213 B.n173 VSUBS 0.006879f
C214 B.n174 VSUBS 0.006879f
C215 B.n175 VSUBS 0.006879f
C216 B.n176 VSUBS 0.006879f
C217 B.n177 VSUBS 0.006879f
C218 B.n178 VSUBS 0.006879f
C219 B.n179 VSUBS 0.006879f
C220 B.n180 VSUBS 0.006879f
C221 B.n181 VSUBS 0.006879f
C222 B.n182 VSUBS 0.006879f
C223 B.n183 VSUBS 0.006879f
C224 B.n184 VSUBS 0.006879f
C225 B.n185 VSUBS 0.006879f
C226 B.n186 VSUBS 0.006879f
C227 B.n187 VSUBS 0.006879f
C228 B.n188 VSUBS 0.006879f
C229 B.n189 VSUBS 0.006879f
C230 B.n190 VSUBS 0.006879f
C231 B.n191 VSUBS 0.006879f
C232 B.n192 VSUBS 0.006879f
C233 B.n193 VSUBS 0.006879f
C234 B.n194 VSUBS 0.006879f
C235 B.n195 VSUBS 0.006879f
C236 B.n196 VSUBS 0.006879f
C237 B.n197 VSUBS 0.006879f
C238 B.n198 VSUBS 0.006879f
C239 B.n199 VSUBS 0.006879f
C240 B.n200 VSUBS 0.006879f
C241 B.n201 VSUBS 0.006879f
C242 B.n202 VSUBS 0.006879f
C243 B.n203 VSUBS 0.006879f
C244 B.n204 VSUBS 0.006879f
C245 B.n205 VSUBS 0.006879f
C246 B.n206 VSUBS 0.006879f
C247 B.n207 VSUBS 0.006879f
C248 B.n208 VSUBS 0.006879f
C249 B.n209 VSUBS 0.006879f
C250 B.n210 VSUBS 0.006879f
C251 B.n211 VSUBS 0.006879f
C252 B.n212 VSUBS 0.006879f
C253 B.n213 VSUBS 0.006879f
C254 B.n214 VSUBS 0.006879f
C255 B.n215 VSUBS 0.006879f
C256 B.n216 VSUBS 0.006879f
C257 B.n217 VSUBS 0.006879f
C258 B.n218 VSUBS 0.01563f
C259 B.n219 VSUBS 0.01563f
C260 B.n220 VSUBS 0.016136f
C261 B.n221 VSUBS 0.006879f
C262 B.n222 VSUBS 0.006879f
C263 B.n223 VSUBS 0.006879f
C264 B.n224 VSUBS 0.006879f
C265 B.n225 VSUBS 0.006879f
C266 B.n226 VSUBS 0.006879f
C267 B.n227 VSUBS 0.006879f
C268 B.n228 VSUBS 0.006879f
C269 B.n229 VSUBS 0.006879f
C270 B.n230 VSUBS 0.006879f
C271 B.n231 VSUBS 0.006879f
C272 B.n232 VSUBS 0.006879f
C273 B.n233 VSUBS 0.006879f
C274 B.n234 VSUBS 0.006879f
C275 B.n235 VSUBS 0.006879f
C276 B.n236 VSUBS 0.006879f
C277 B.n237 VSUBS 0.006879f
C278 B.n238 VSUBS 0.006879f
C279 B.n239 VSUBS 0.006879f
C280 B.n240 VSUBS 0.006879f
C281 B.n241 VSUBS 0.006879f
C282 B.n242 VSUBS 0.006879f
C283 B.n243 VSUBS 0.006879f
C284 B.n244 VSUBS 0.006879f
C285 B.n245 VSUBS 0.006879f
C286 B.n246 VSUBS 0.006879f
C287 B.n247 VSUBS 0.006879f
C288 B.n248 VSUBS 0.006879f
C289 B.n249 VSUBS 0.006879f
C290 B.n250 VSUBS 0.006879f
C291 B.n251 VSUBS 0.006879f
C292 B.n252 VSUBS 0.006879f
C293 B.n253 VSUBS 0.006879f
C294 B.n254 VSUBS 0.006879f
C295 B.n255 VSUBS 0.006879f
C296 B.n256 VSUBS 0.006879f
C297 B.n257 VSUBS 0.006879f
C298 B.n258 VSUBS 0.006879f
C299 B.n259 VSUBS 0.006879f
C300 B.n260 VSUBS 0.006879f
C301 B.n261 VSUBS 0.006879f
C302 B.n262 VSUBS 0.006879f
C303 B.n263 VSUBS 0.006879f
C304 B.n264 VSUBS 0.006879f
C305 B.n265 VSUBS 0.006879f
C306 B.n266 VSUBS 0.006879f
C307 B.n267 VSUBS 0.006879f
C308 B.n268 VSUBS 0.006879f
C309 B.n269 VSUBS 0.006879f
C310 B.n270 VSUBS 0.006879f
C311 B.n271 VSUBS 0.006879f
C312 B.n272 VSUBS 0.006879f
C313 B.n273 VSUBS 0.006879f
C314 B.n274 VSUBS 0.006879f
C315 B.n275 VSUBS 0.006879f
C316 B.n276 VSUBS 0.006879f
C317 B.n277 VSUBS 0.006879f
C318 B.n278 VSUBS 0.006879f
C319 B.n279 VSUBS 0.006879f
C320 B.n280 VSUBS 0.006879f
C321 B.n281 VSUBS 0.006879f
C322 B.n282 VSUBS 0.006879f
C323 B.n283 VSUBS 0.006879f
C324 B.n284 VSUBS 0.006879f
C325 B.n285 VSUBS 0.006879f
C326 B.n286 VSUBS 0.006879f
C327 B.n287 VSUBS 0.006879f
C328 B.n288 VSUBS 0.006879f
C329 B.n289 VSUBS 0.006879f
C330 B.n290 VSUBS 0.006879f
C331 B.n291 VSUBS 0.006879f
C332 B.n292 VSUBS 0.006879f
C333 B.n293 VSUBS 0.006879f
C334 B.n294 VSUBS 0.006879f
C335 B.n295 VSUBS 0.006879f
C336 B.n296 VSUBS 0.006879f
C337 B.n297 VSUBS 0.006879f
C338 B.n298 VSUBS 0.006879f
C339 B.n299 VSUBS 0.006879f
C340 B.n300 VSUBS 0.006879f
C341 B.n301 VSUBS 0.006879f
C342 B.n302 VSUBS 0.006474f
C343 B.n303 VSUBS 0.006879f
C344 B.n304 VSUBS 0.006879f
C345 B.n305 VSUBS 0.003844f
C346 B.n306 VSUBS 0.006879f
C347 B.n307 VSUBS 0.006879f
C348 B.n308 VSUBS 0.006879f
C349 B.n309 VSUBS 0.006879f
C350 B.n310 VSUBS 0.006879f
C351 B.n311 VSUBS 0.006879f
C352 B.n312 VSUBS 0.006879f
C353 B.n313 VSUBS 0.006879f
C354 B.n314 VSUBS 0.006879f
C355 B.n315 VSUBS 0.006879f
C356 B.n316 VSUBS 0.006879f
C357 B.n317 VSUBS 0.006879f
C358 B.n318 VSUBS 0.003844f
C359 B.n319 VSUBS 0.015938f
C360 B.n320 VSUBS 0.006474f
C361 B.n321 VSUBS 0.006879f
C362 B.n322 VSUBS 0.006879f
C363 B.n323 VSUBS 0.006879f
C364 B.n324 VSUBS 0.006879f
C365 B.n325 VSUBS 0.006879f
C366 B.n326 VSUBS 0.006879f
C367 B.n327 VSUBS 0.006879f
C368 B.n328 VSUBS 0.006879f
C369 B.n329 VSUBS 0.006879f
C370 B.n330 VSUBS 0.006879f
C371 B.n331 VSUBS 0.006879f
C372 B.n332 VSUBS 0.006879f
C373 B.n333 VSUBS 0.006879f
C374 B.n334 VSUBS 0.006879f
C375 B.n335 VSUBS 0.006879f
C376 B.n336 VSUBS 0.006879f
C377 B.n337 VSUBS 0.006879f
C378 B.n338 VSUBS 0.006879f
C379 B.n339 VSUBS 0.006879f
C380 B.n340 VSUBS 0.006879f
C381 B.n341 VSUBS 0.006879f
C382 B.n342 VSUBS 0.006879f
C383 B.n343 VSUBS 0.006879f
C384 B.n344 VSUBS 0.006879f
C385 B.n345 VSUBS 0.006879f
C386 B.n346 VSUBS 0.006879f
C387 B.n347 VSUBS 0.006879f
C388 B.n348 VSUBS 0.006879f
C389 B.n349 VSUBS 0.006879f
C390 B.n350 VSUBS 0.006879f
C391 B.n351 VSUBS 0.006879f
C392 B.n352 VSUBS 0.006879f
C393 B.n353 VSUBS 0.006879f
C394 B.n354 VSUBS 0.006879f
C395 B.n355 VSUBS 0.006879f
C396 B.n356 VSUBS 0.006879f
C397 B.n357 VSUBS 0.006879f
C398 B.n358 VSUBS 0.006879f
C399 B.n359 VSUBS 0.006879f
C400 B.n360 VSUBS 0.006879f
C401 B.n361 VSUBS 0.006879f
C402 B.n362 VSUBS 0.006879f
C403 B.n363 VSUBS 0.006879f
C404 B.n364 VSUBS 0.006879f
C405 B.n365 VSUBS 0.006879f
C406 B.n366 VSUBS 0.006879f
C407 B.n367 VSUBS 0.006879f
C408 B.n368 VSUBS 0.006879f
C409 B.n369 VSUBS 0.006879f
C410 B.n370 VSUBS 0.006879f
C411 B.n371 VSUBS 0.006879f
C412 B.n372 VSUBS 0.006879f
C413 B.n373 VSUBS 0.006879f
C414 B.n374 VSUBS 0.006879f
C415 B.n375 VSUBS 0.006879f
C416 B.n376 VSUBS 0.006879f
C417 B.n377 VSUBS 0.006879f
C418 B.n378 VSUBS 0.006879f
C419 B.n379 VSUBS 0.006879f
C420 B.n380 VSUBS 0.006879f
C421 B.n381 VSUBS 0.006879f
C422 B.n382 VSUBS 0.006879f
C423 B.n383 VSUBS 0.006879f
C424 B.n384 VSUBS 0.006879f
C425 B.n385 VSUBS 0.006879f
C426 B.n386 VSUBS 0.006879f
C427 B.n387 VSUBS 0.006879f
C428 B.n388 VSUBS 0.006879f
C429 B.n389 VSUBS 0.006879f
C430 B.n390 VSUBS 0.006879f
C431 B.n391 VSUBS 0.006879f
C432 B.n392 VSUBS 0.006879f
C433 B.n393 VSUBS 0.006879f
C434 B.n394 VSUBS 0.006879f
C435 B.n395 VSUBS 0.006879f
C436 B.n396 VSUBS 0.006879f
C437 B.n397 VSUBS 0.006879f
C438 B.n398 VSUBS 0.006879f
C439 B.n399 VSUBS 0.006879f
C440 B.n400 VSUBS 0.006879f
C441 B.n401 VSUBS 0.006879f
C442 B.n402 VSUBS 0.006879f
C443 B.n403 VSUBS 0.016136f
C444 B.n404 VSUBS 0.01563f
C445 B.n405 VSUBS 0.01563f
C446 B.n406 VSUBS 0.006879f
C447 B.n407 VSUBS 0.006879f
C448 B.n408 VSUBS 0.006879f
C449 B.n409 VSUBS 0.006879f
C450 B.n410 VSUBS 0.006879f
C451 B.n411 VSUBS 0.006879f
C452 B.n412 VSUBS 0.006879f
C453 B.n413 VSUBS 0.006879f
C454 B.n414 VSUBS 0.006879f
C455 B.n415 VSUBS 0.006879f
C456 B.n416 VSUBS 0.006879f
C457 B.n417 VSUBS 0.006879f
C458 B.n418 VSUBS 0.006879f
C459 B.n419 VSUBS 0.006879f
C460 B.n420 VSUBS 0.006879f
C461 B.n421 VSUBS 0.006879f
C462 B.n422 VSUBS 0.006879f
C463 B.n423 VSUBS 0.006879f
C464 B.n424 VSUBS 0.006879f
C465 B.n425 VSUBS 0.006879f
C466 B.n426 VSUBS 0.006879f
C467 B.n427 VSUBS 0.006879f
C468 B.n428 VSUBS 0.006879f
C469 B.n429 VSUBS 0.006879f
C470 B.n430 VSUBS 0.006879f
C471 B.n431 VSUBS 0.006879f
C472 B.n432 VSUBS 0.006879f
C473 B.n433 VSUBS 0.006879f
C474 B.n434 VSUBS 0.006879f
C475 B.n435 VSUBS 0.006879f
C476 B.n436 VSUBS 0.006879f
C477 B.n437 VSUBS 0.006879f
C478 B.n438 VSUBS 0.006879f
C479 B.n439 VSUBS 0.006879f
C480 B.n440 VSUBS 0.006879f
C481 B.n441 VSUBS 0.006879f
C482 B.n442 VSUBS 0.006879f
C483 B.n443 VSUBS 0.006879f
C484 B.n444 VSUBS 0.006879f
C485 B.n445 VSUBS 0.006879f
C486 B.n446 VSUBS 0.006879f
C487 B.n447 VSUBS 0.006879f
C488 B.n448 VSUBS 0.006879f
C489 B.n449 VSUBS 0.006879f
C490 B.n450 VSUBS 0.006879f
C491 B.n451 VSUBS 0.006879f
C492 B.n452 VSUBS 0.006879f
C493 B.n453 VSUBS 0.006879f
C494 B.n454 VSUBS 0.006879f
C495 B.n455 VSUBS 0.006879f
C496 B.n456 VSUBS 0.006879f
C497 B.n457 VSUBS 0.006879f
C498 B.n458 VSUBS 0.006879f
C499 B.n459 VSUBS 0.006879f
C500 B.n460 VSUBS 0.006879f
C501 B.n461 VSUBS 0.006879f
C502 B.n462 VSUBS 0.006879f
C503 B.n463 VSUBS 0.006879f
C504 B.n464 VSUBS 0.006879f
C505 B.n465 VSUBS 0.006879f
C506 B.n466 VSUBS 0.006879f
C507 B.n467 VSUBS 0.006879f
C508 B.n468 VSUBS 0.006879f
C509 B.n469 VSUBS 0.006879f
C510 B.n470 VSUBS 0.006879f
C511 B.n471 VSUBS 0.006879f
C512 B.n472 VSUBS 0.006879f
C513 B.n473 VSUBS 0.006879f
C514 B.n474 VSUBS 0.006879f
C515 B.n475 VSUBS 0.006879f
C516 B.n476 VSUBS 0.006879f
C517 B.n477 VSUBS 0.006879f
C518 B.n478 VSUBS 0.006879f
C519 B.n479 VSUBS 0.01563f
C520 B.n480 VSUBS 0.016459f
C521 B.n481 VSUBS 0.015306f
C522 B.n482 VSUBS 0.006879f
C523 B.n483 VSUBS 0.006879f
C524 B.n484 VSUBS 0.006879f
C525 B.n485 VSUBS 0.006879f
C526 B.n486 VSUBS 0.006879f
C527 B.n487 VSUBS 0.006879f
C528 B.n488 VSUBS 0.006879f
C529 B.n489 VSUBS 0.006879f
C530 B.n490 VSUBS 0.006879f
C531 B.n491 VSUBS 0.006879f
C532 B.n492 VSUBS 0.006879f
C533 B.n493 VSUBS 0.006879f
C534 B.n494 VSUBS 0.006879f
C535 B.n495 VSUBS 0.006879f
C536 B.n496 VSUBS 0.006879f
C537 B.n497 VSUBS 0.006879f
C538 B.n498 VSUBS 0.006879f
C539 B.n499 VSUBS 0.006879f
C540 B.n500 VSUBS 0.006879f
C541 B.n501 VSUBS 0.006879f
C542 B.n502 VSUBS 0.006879f
C543 B.n503 VSUBS 0.006879f
C544 B.n504 VSUBS 0.006879f
C545 B.n505 VSUBS 0.006879f
C546 B.n506 VSUBS 0.006879f
C547 B.n507 VSUBS 0.006879f
C548 B.n508 VSUBS 0.006879f
C549 B.n509 VSUBS 0.006879f
C550 B.n510 VSUBS 0.006879f
C551 B.n511 VSUBS 0.006879f
C552 B.n512 VSUBS 0.006879f
C553 B.n513 VSUBS 0.006879f
C554 B.n514 VSUBS 0.006879f
C555 B.n515 VSUBS 0.006879f
C556 B.n516 VSUBS 0.006879f
C557 B.n517 VSUBS 0.006879f
C558 B.n518 VSUBS 0.006879f
C559 B.n519 VSUBS 0.006879f
C560 B.n520 VSUBS 0.006879f
C561 B.n521 VSUBS 0.006879f
C562 B.n522 VSUBS 0.006879f
C563 B.n523 VSUBS 0.006879f
C564 B.n524 VSUBS 0.006879f
C565 B.n525 VSUBS 0.006879f
C566 B.n526 VSUBS 0.006879f
C567 B.n527 VSUBS 0.006879f
C568 B.n528 VSUBS 0.006879f
C569 B.n529 VSUBS 0.006879f
C570 B.n530 VSUBS 0.006879f
C571 B.n531 VSUBS 0.006879f
C572 B.n532 VSUBS 0.006879f
C573 B.n533 VSUBS 0.006879f
C574 B.n534 VSUBS 0.006879f
C575 B.n535 VSUBS 0.006879f
C576 B.n536 VSUBS 0.006879f
C577 B.n537 VSUBS 0.006879f
C578 B.n538 VSUBS 0.006879f
C579 B.n539 VSUBS 0.006879f
C580 B.n540 VSUBS 0.006879f
C581 B.n541 VSUBS 0.006879f
C582 B.n542 VSUBS 0.006879f
C583 B.n543 VSUBS 0.006879f
C584 B.n544 VSUBS 0.006879f
C585 B.n545 VSUBS 0.006879f
C586 B.n546 VSUBS 0.006879f
C587 B.n547 VSUBS 0.006879f
C588 B.n548 VSUBS 0.006879f
C589 B.n549 VSUBS 0.006879f
C590 B.n550 VSUBS 0.006879f
C591 B.n551 VSUBS 0.006879f
C592 B.n552 VSUBS 0.006879f
C593 B.n553 VSUBS 0.006879f
C594 B.n554 VSUBS 0.006879f
C595 B.n555 VSUBS 0.006879f
C596 B.n556 VSUBS 0.006879f
C597 B.n557 VSUBS 0.006879f
C598 B.n558 VSUBS 0.006879f
C599 B.n559 VSUBS 0.006879f
C600 B.n560 VSUBS 0.006879f
C601 B.n561 VSUBS 0.006879f
C602 B.n562 VSUBS 0.006879f
C603 B.n563 VSUBS 0.006879f
C604 B.n564 VSUBS 0.006474f
C605 B.n565 VSUBS 0.015938f
C606 B.n566 VSUBS 0.003844f
C607 B.n567 VSUBS 0.006879f
C608 B.n568 VSUBS 0.006879f
C609 B.n569 VSUBS 0.006879f
C610 B.n570 VSUBS 0.006879f
C611 B.n571 VSUBS 0.006879f
C612 B.n572 VSUBS 0.006879f
C613 B.n573 VSUBS 0.006879f
C614 B.n574 VSUBS 0.006879f
C615 B.n575 VSUBS 0.006879f
C616 B.n576 VSUBS 0.006879f
C617 B.n577 VSUBS 0.006879f
C618 B.n578 VSUBS 0.006879f
C619 B.n579 VSUBS 0.003844f
C620 B.n580 VSUBS 0.006879f
C621 B.n581 VSUBS 0.006879f
C622 B.n582 VSUBS 0.006879f
C623 B.n583 VSUBS 0.006879f
C624 B.n584 VSUBS 0.006879f
C625 B.n585 VSUBS 0.006879f
C626 B.n586 VSUBS 0.006879f
C627 B.n587 VSUBS 0.006879f
C628 B.n588 VSUBS 0.006879f
C629 B.n589 VSUBS 0.006879f
C630 B.n590 VSUBS 0.006879f
C631 B.n591 VSUBS 0.006879f
C632 B.n592 VSUBS 0.006879f
C633 B.n593 VSUBS 0.006879f
C634 B.n594 VSUBS 0.006879f
C635 B.n595 VSUBS 0.006879f
C636 B.n596 VSUBS 0.006879f
C637 B.n597 VSUBS 0.006879f
C638 B.n598 VSUBS 0.006879f
C639 B.n599 VSUBS 0.006879f
C640 B.n600 VSUBS 0.006879f
C641 B.n601 VSUBS 0.006879f
C642 B.n602 VSUBS 0.006879f
C643 B.n603 VSUBS 0.006879f
C644 B.n604 VSUBS 0.006879f
C645 B.n605 VSUBS 0.006879f
C646 B.n606 VSUBS 0.006879f
C647 B.n607 VSUBS 0.006879f
C648 B.n608 VSUBS 0.006879f
C649 B.n609 VSUBS 0.006879f
C650 B.n610 VSUBS 0.006879f
C651 B.n611 VSUBS 0.006879f
C652 B.n612 VSUBS 0.006879f
C653 B.n613 VSUBS 0.006879f
C654 B.n614 VSUBS 0.006879f
C655 B.n615 VSUBS 0.006879f
C656 B.n616 VSUBS 0.006879f
C657 B.n617 VSUBS 0.006879f
C658 B.n618 VSUBS 0.006879f
C659 B.n619 VSUBS 0.006879f
C660 B.n620 VSUBS 0.006879f
C661 B.n621 VSUBS 0.006879f
C662 B.n622 VSUBS 0.006879f
C663 B.n623 VSUBS 0.006879f
C664 B.n624 VSUBS 0.006879f
C665 B.n625 VSUBS 0.006879f
C666 B.n626 VSUBS 0.006879f
C667 B.n627 VSUBS 0.006879f
C668 B.n628 VSUBS 0.006879f
C669 B.n629 VSUBS 0.006879f
C670 B.n630 VSUBS 0.006879f
C671 B.n631 VSUBS 0.006879f
C672 B.n632 VSUBS 0.006879f
C673 B.n633 VSUBS 0.006879f
C674 B.n634 VSUBS 0.006879f
C675 B.n635 VSUBS 0.006879f
C676 B.n636 VSUBS 0.006879f
C677 B.n637 VSUBS 0.006879f
C678 B.n638 VSUBS 0.006879f
C679 B.n639 VSUBS 0.006879f
C680 B.n640 VSUBS 0.006879f
C681 B.n641 VSUBS 0.006879f
C682 B.n642 VSUBS 0.006879f
C683 B.n643 VSUBS 0.006879f
C684 B.n644 VSUBS 0.006879f
C685 B.n645 VSUBS 0.006879f
C686 B.n646 VSUBS 0.006879f
C687 B.n647 VSUBS 0.006879f
C688 B.n648 VSUBS 0.006879f
C689 B.n649 VSUBS 0.006879f
C690 B.n650 VSUBS 0.006879f
C691 B.n651 VSUBS 0.006879f
C692 B.n652 VSUBS 0.006879f
C693 B.n653 VSUBS 0.006879f
C694 B.n654 VSUBS 0.006879f
C695 B.n655 VSUBS 0.006879f
C696 B.n656 VSUBS 0.006879f
C697 B.n657 VSUBS 0.006879f
C698 B.n658 VSUBS 0.006879f
C699 B.n659 VSUBS 0.006879f
C700 B.n660 VSUBS 0.006879f
C701 B.n661 VSUBS 0.006879f
C702 B.n662 VSUBS 0.006879f
C703 B.n663 VSUBS 0.016136f
C704 B.n664 VSUBS 0.016136f
C705 B.n665 VSUBS 0.01563f
C706 B.n666 VSUBS 0.006879f
C707 B.n667 VSUBS 0.006879f
C708 B.n668 VSUBS 0.006879f
C709 B.n669 VSUBS 0.006879f
C710 B.n670 VSUBS 0.006879f
C711 B.n671 VSUBS 0.006879f
C712 B.n672 VSUBS 0.006879f
C713 B.n673 VSUBS 0.006879f
C714 B.n674 VSUBS 0.006879f
C715 B.n675 VSUBS 0.006879f
C716 B.n676 VSUBS 0.006879f
C717 B.n677 VSUBS 0.006879f
C718 B.n678 VSUBS 0.006879f
C719 B.n679 VSUBS 0.006879f
C720 B.n680 VSUBS 0.006879f
C721 B.n681 VSUBS 0.006879f
C722 B.n682 VSUBS 0.006879f
C723 B.n683 VSUBS 0.006879f
C724 B.n684 VSUBS 0.006879f
C725 B.n685 VSUBS 0.006879f
C726 B.n686 VSUBS 0.006879f
C727 B.n687 VSUBS 0.006879f
C728 B.n688 VSUBS 0.006879f
C729 B.n689 VSUBS 0.006879f
C730 B.n690 VSUBS 0.006879f
C731 B.n691 VSUBS 0.006879f
C732 B.n692 VSUBS 0.006879f
C733 B.n693 VSUBS 0.006879f
C734 B.n694 VSUBS 0.006879f
C735 B.n695 VSUBS 0.006879f
C736 B.n696 VSUBS 0.006879f
C737 B.n697 VSUBS 0.006879f
C738 B.n698 VSUBS 0.006879f
C739 B.n699 VSUBS 0.006879f
C740 B.n700 VSUBS 0.006879f
C741 B.n701 VSUBS 0.006879f
C742 B.n702 VSUBS 0.006879f
C743 B.n703 VSUBS 0.015577f
C744 VDD2.t2 VSUBS 0.357304f
C745 VDD2.t1 VSUBS 0.357304f
C746 VDD2.n0 VSUBS 3.78455f
C747 VDD2.t0 VSUBS 0.357304f
C748 VDD2.t3 VSUBS 0.357304f
C749 VDD2.n1 VSUBS 2.96273f
C750 VDD2.n2 VSUBS 4.57731f
C751 VN.t1 VSUBS 3.09126f
C752 VN.t2 VSUBS 3.08994f
C753 VN.n0 VSUBS 2.17373f
C754 VN.t0 VSUBS 3.09126f
C755 VN.t3 VSUBS 3.08994f
C756 VN.n1 VSUBS 3.92771f
C757 VTAIL.n0 VSUBS 0.025029f
C758 VTAIL.n1 VSUBS 0.021931f
C759 VTAIL.n2 VSUBS 0.011785f
C760 VTAIL.n3 VSUBS 0.027855f
C761 VTAIL.n4 VSUBS 0.012478f
C762 VTAIL.n5 VSUBS 0.021931f
C763 VTAIL.n6 VSUBS 0.011785f
C764 VTAIL.n7 VSUBS 0.027855f
C765 VTAIL.n8 VSUBS 0.012478f
C766 VTAIL.n9 VSUBS 0.021931f
C767 VTAIL.n10 VSUBS 0.011785f
C768 VTAIL.n11 VSUBS 0.027855f
C769 VTAIL.n12 VSUBS 0.012478f
C770 VTAIL.n13 VSUBS 0.021931f
C771 VTAIL.n14 VSUBS 0.011785f
C772 VTAIL.n15 VSUBS 0.027855f
C773 VTAIL.n16 VSUBS 0.012478f
C774 VTAIL.n17 VSUBS 0.021931f
C775 VTAIL.n18 VSUBS 0.011785f
C776 VTAIL.n19 VSUBS 0.027855f
C777 VTAIL.n20 VSUBS 0.012478f
C778 VTAIL.n21 VSUBS 0.021931f
C779 VTAIL.n22 VSUBS 0.011785f
C780 VTAIL.n23 VSUBS 0.027855f
C781 VTAIL.n24 VSUBS 0.012478f
C782 VTAIL.n25 VSUBS 0.021931f
C783 VTAIL.n26 VSUBS 0.011785f
C784 VTAIL.n27 VSUBS 0.027855f
C785 VTAIL.n28 VSUBS 0.012478f
C786 VTAIL.n29 VSUBS 0.16747f
C787 VTAIL.t1 VSUBS 0.059741f
C788 VTAIL.n30 VSUBS 0.020892f
C789 VTAIL.n31 VSUBS 0.01772f
C790 VTAIL.n32 VSUBS 0.011785f
C791 VTAIL.n33 VSUBS 1.5985f
C792 VTAIL.n34 VSUBS 0.021931f
C793 VTAIL.n35 VSUBS 0.011785f
C794 VTAIL.n36 VSUBS 0.012478f
C795 VTAIL.n37 VSUBS 0.027855f
C796 VTAIL.n38 VSUBS 0.027855f
C797 VTAIL.n39 VSUBS 0.012478f
C798 VTAIL.n40 VSUBS 0.011785f
C799 VTAIL.n41 VSUBS 0.021931f
C800 VTAIL.n42 VSUBS 0.021931f
C801 VTAIL.n43 VSUBS 0.011785f
C802 VTAIL.n44 VSUBS 0.012478f
C803 VTAIL.n45 VSUBS 0.027855f
C804 VTAIL.n46 VSUBS 0.027855f
C805 VTAIL.n47 VSUBS 0.012478f
C806 VTAIL.n48 VSUBS 0.011785f
C807 VTAIL.n49 VSUBS 0.021931f
C808 VTAIL.n50 VSUBS 0.021931f
C809 VTAIL.n51 VSUBS 0.011785f
C810 VTAIL.n52 VSUBS 0.012478f
C811 VTAIL.n53 VSUBS 0.027855f
C812 VTAIL.n54 VSUBS 0.027855f
C813 VTAIL.n55 VSUBS 0.012478f
C814 VTAIL.n56 VSUBS 0.011785f
C815 VTAIL.n57 VSUBS 0.021931f
C816 VTAIL.n58 VSUBS 0.021931f
C817 VTAIL.n59 VSUBS 0.011785f
C818 VTAIL.n60 VSUBS 0.012478f
C819 VTAIL.n61 VSUBS 0.027855f
C820 VTAIL.n62 VSUBS 0.027855f
C821 VTAIL.n63 VSUBS 0.012478f
C822 VTAIL.n64 VSUBS 0.011785f
C823 VTAIL.n65 VSUBS 0.021931f
C824 VTAIL.n66 VSUBS 0.021931f
C825 VTAIL.n67 VSUBS 0.011785f
C826 VTAIL.n68 VSUBS 0.012478f
C827 VTAIL.n69 VSUBS 0.027855f
C828 VTAIL.n70 VSUBS 0.027855f
C829 VTAIL.n71 VSUBS 0.027855f
C830 VTAIL.n72 VSUBS 0.012478f
C831 VTAIL.n73 VSUBS 0.011785f
C832 VTAIL.n74 VSUBS 0.021931f
C833 VTAIL.n75 VSUBS 0.021931f
C834 VTAIL.n76 VSUBS 0.011785f
C835 VTAIL.n77 VSUBS 0.012132f
C836 VTAIL.n78 VSUBS 0.012132f
C837 VTAIL.n79 VSUBS 0.027855f
C838 VTAIL.n80 VSUBS 0.027855f
C839 VTAIL.n81 VSUBS 0.012478f
C840 VTAIL.n82 VSUBS 0.011785f
C841 VTAIL.n83 VSUBS 0.021931f
C842 VTAIL.n84 VSUBS 0.021931f
C843 VTAIL.n85 VSUBS 0.011785f
C844 VTAIL.n86 VSUBS 0.012478f
C845 VTAIL.n87 VSUBS 0.027855f
C846 VTAIL.n88 VSUBS 0.070606f
C847 VTAIL.n89 VSUBS 0.012478f
C848 VTAIL.n90 VSUBS 0.011785f
C849 VTAIL.n91 VSUBS 0.056386f
C850 VTAIL.n92 VSUBS 0.035815f
C851 VTAIL.n93 VSUBS 0.117141f
C852 VTAIL.n94 VSUBS 0.025029f
C853 VTAIL.n95 VSUBS 0.021931f
C854 VTAIL.n96 VSUBS 0.011785f
C855 VTAIL.n97 VSUBS 0.027855f
C856 VTAIL.n98 VSUBS 0.012478f
C857 VTAIL.n99 VSUBS 0.021931f
C858 VTAIL.n100 VSUBS 0.011785f
C859 VTAIL.n101 VSUBS 0.027855f
C860 VTAIL.n102 VSUBS 0.012478f
C861 VTAIL.n103 VSUBS 0.021931f
C862 VTAIL.n104 VSUBS 0.011785f
C863 VTAIL.n105 VSUBS 0.027855f
C864 VTAIL.n106 VSUBS 0.012478f
C865 VTAIL.n107 VSUBS 0.021931f
C866 VTAIL.n108 VSUBS 0.011785f
C867 VTAIL.n109 VSUBS 0.027855f
C868 VTAIL.n110 VSUBS 0.012478f
C869 VTAIL.n111 VSUBS 0.021931f
C870 VTAIL.n112 VSUBS 0.011785f
C871 VTAIL.n113 VSUBS 0.027855f
C872 VTAIL.n114 VSUBS 0.012478f
C873 VTAIL.n115 VSUBS 0.021931f
C874 VTAIL.n116 VSUBS 0.011785f
C875 VTAIL.n117 VSUBS 0.027855f
C876 VTAIL.n118 VSUBS 0.012478f
C877 VTAIL.n119 VSUBS 0.021931f
C878 VTAIL.n120 VSUBS 0.011785f
C879 VTAIL.n121 VSUBS 0.027855f
C880 VTAIL.n122 VSUBS 0.012478f
C881 VTAIL.n123 VSUBS 0.16747f
C882 VTAIL.t4 VSUBS 0.059741f
C883 VTAIL.n124 VSUBS 0.020892f
C884 VTAIL.n125 VSUBS 0.01772f
C885 VTAIL.n126 VSUBS 0.011785f
C886 VTAIL.n127 VSUBS 1.5985f
C887 VTAIL.n128 VSUBS 0.021931f
C888 VTAIL.n129 VSUBS 0.011785f
C889 VTAIL.n130 VSUBS 0.012478f
C890 VTAIL.n131 VSUBS 0.027855f
C891 VTAIL.n132 VSUBS 0.027855f
C892 VTAIL.n133 VSUBS 0.012478f
C893 VTAIL.n134 VSUBS 0.011785f
C894 VTAIL.n135 VSUBS 0.021931f
C895 VTAIL.n136 VSUBS 0.021931f
C896 VTAIL.n137 VSUBS 0.011785f
C897 VTAIL.n138 VSUBS 0.012478f
C898 VTAIL.n139 VSUBS 0.027855f
C899 VTAIL.n140 VSUBS 0.027855f
C900 VTAIL.n141 VSUBS 0.012478f
C901 VTAIL.n142 VSUBS 0.011785f
C902 VTAIL.n143 VSUBS 0.021931f
C903 VTAIL.n144 VSUBS 0.021931f
C904 VTAIL.n145 VSUBS 0.011785f
C905 VTAIL.n146 VSUBS 0.012478f
C906 VTAIL.n147 VSUBS 0.027855f
C907 VTAIL.n148 VSUBS 0.027855f
C908 VTAIL.n149 VSUBS 0.012478f
C909 VTAIL.n150 VSUBS 0.011785f
C910 VTAIL.n151 VSUBS 0.021931f
C911 VTAIL.n152 VSUBS 0.021931f
C912 VTAIL.n153 VSUBS 0.011785f
C913 VTAIL.n154 VSUBS 0.012478f
C914 VTAIL.n155 VSUBS 0.027855f
C915 VTAIL.n156 VSUBS 0.027855f
C916 VTAIL.n157 VSUBS 0.012478f
C917 VTAIL.n158 VSUBS 0.011785f
C918 VTAIL.n159 VSUBS 0.021931f
C919 VTAIL.n160 VSUBS 0.021931f
C920 VTAIL.n161 VSUBS 0.011785f
C921 VTAIL.n162 VSUBS 0.012478f
C922 VTAIL.n163 VSUBS 0.027855f
C923 VTAIL.n164 VSUBS 0.027855f
C924 VTAIL.n165 VSUBS 0.027855f
C925 VTAIL.n166 VSUBS 0.012478f
C926 VTAIL.n167 VSUBS 0.011785f
C927 VTAIL.n168 VSUBS 0.021931f
C928 VTAIL.n169 VSUBS 0.021931f
C929 VTAIL.n170 VSUBS 0.011785f
C930 VTAIL.n171 VSUBS 0.012132f
C931 VTAIL.n172 VSUBS 0.012132f
C932 VTAIL.n173 VSUBS 0.027855f
C933 VTAIL.n174 VSUBS 0.027855f
C934 VTAIL.n175 VSUBS 0.012478f
C935 VTAIL.n176 VSUBS 0.011785f
C936 VTAIL.n177 VSUBS 0.021931f
C937 VTAIL.n178 VSUBS 0.021931f
C938 VTAIL.n179 VSUBS 0.011785f
C939 VTAIL.n180 VSUBS 0.012478f
C940 VTAIL.n181 VSUBS 0.027855f
C941 VTAIL.n182 VSUBS 0.070606f
C942 VTAIL.n183 VSUBS 0.012478f
C943 VTAIL.n184 VSUBS 0.011785f
C944 VTAIL.n185 VSUBS 0.056386f
C945 VTAIL.n186 VSUBS 0.035815f
C946 VTAIL.n187 VSUBS 0.170903f
C947 VTAIL.n188 VSUBS 0.025029f
C948 VTAIL.n189 VSUBS 0.021931f
C949 VTAIL.n190 VSUBS 0.011785f
C950 VTAIL.n191 VSUBS 0.027855f
C951 VTAIL.n192 VSUBS 0.012478f
C952 VTAIL.n193 VSUBS 0.021931f
C953 VTAIL.n194 VSUBS 0.011785f
C954 VTAIL.n195 VSUBS 0.027855f
C955 VTAIL.n196 VSUBS 0.012478f
C956 VTAIL.n197 VSUBS 0.021931f
C957 VTAIL.n198 VSUBS 0.011785f
C958 VTAIL.n199 VSUBS 0.027855f
C959 VTAIL.n200 VSUBS 0.012478f
C960 VTAIL.n201 VSUBS 0.021931f
C961 VTAIL.n202 VSUBS 0.011785f
C962 VTAIL.n203 VSUBS 0.027855f
C963 VTAIL.n204 VSUBS 0.012478f
C964 VTAIL.n205 VSUBS 0.021931f
C965 VTAIL.n206 VSUBS 0.011785f
C966 VTAIL.n207 VSUBS 0.027855f
C967 VTAIL.n208 VSUBS 0.012478f
C968 VTAIL.n209 VSUBS 0.021931f
C969 VTAIL.n210 VSUBS 0.011785f
C970 VTAIL.n211 VSUBS 0.027855f
C971 VTAIL.n212 VSUBS 0.012478f
C972 VTAIL.n213 VSUBS 0.021931f
C973 VTAIL.n214 VSUBS 0.011785f
C974 VTAIL.n215 VSUBS 0.027855f
C975 VTAIL.n216 VSUBS 0.012478f
C976 VTAIL.n217 VSUBS 0.16747f
C977 VTAIL.t7 VSUBS 0.059741f
C978 VTAIL.n218 VSUBS 0.020892f
C979 VTAIL.n219 VSUBS 0.01772f
C980 VTAIL.n220 VSUBS 0.011785f
C981 VTAIL.n221 VSUBS 1.5985f
C982 VTAIL.n222 VSUBS 0.021931f
C983 VTAIL.n223 VSUBS 0.011785f
C984 VTAIL.n224 VSUBS 0.012478f
C985 VTAIL.n225 VSUBS 0.027855f
C986 VTAIL.n226 VSUBS 0.027855f
C987 VTAIL.n227 VSUBS 0.012478f
C988 VTAIL.n228 VSUBS 0.011785f
C989 VTAIL.n229 VSUBS 0.021931f
C990 VTAIL.n230 VSUBS 0.021931f
C991 VTAIL.n231 VSUBS 0.011785f
C992 VTAIL.n232 VSUBS 0.012478f
C993 VTAIL.n233 VSUBS 0.027855f
C994 VTAIL.n234 VSUBS 0.027855f
C995 VTAIL.n235 VSUBS 0.012478f
C996 VTAIL.n236 VSUBS 0.011785f
C997 VTAIL.n237 VSUBS 0.021931f
C998 VTAIL.n238 VSUBS 0.021931f
C999 VTAIL.n239 VSUBS 0.011785f
C1000 VTAIL.n240 VSUBS 0.012478f
C1001 VTAIL.n241 VSUBS 0.027855f
C1002 VTAIL.n242 VSUBS 0.027855f
C1003 VTAIL.n243 VSUBS 0.012478f
C1004 VTAIL.n244 VSUBS 0.011785f
C1005 VTAIL.n245 VSUBS 0.021931f
C1006 VTAIL.n246 VSUBS 0.021931f
C1007 VTAIL.n247 VSUBS 0.011785f
C1008 VTAIL.n248 VSUBS 0.012478f
C1009 VTAIL.n249 VSUBS 0.027855f
C1010 VTAIL.n250 VSUBS 0.027855f
C1011 VTAIL.n251 VSUBS 0.012478f
C1012 VTAIL.n252 VSUBS 0.011785f
C1013 VTAIL.n253 VSUBS 0.021931f
C1014 VTAIL.n254 VSUBS 0.021931f
C1015 VTAIL.n255 VSUBS 0.011785f
C1016 VTAIL.n256 VSUBS 0.012478f
C1017 VTAIL.n257 VSUBS 0.027855f
C1018 VTAIL.n258 VSUBS 0.027855f
C1019 VTAIL.n259 VSUBS 0.027855f
C1020 VTAIL.n260 VSUBS 0.012478f
C1021 VTAIL.n261 VSUBS 0.011785f
C1022 VTAIL.n262 VSUBS 0.021931f
C1023 VTAIL.n263 VSUBS 0.021931f
C1024 VTAIL.n264 VSUBS 0.011785f
C1025 VTAIL.n265 VSUBS 0.012132f
C1026 VTAIL.n266 VSUBS 0.012132f
C1027 VTAIL.n267 VSUBS 0.027855f
C1028 VTAIL.n268 VSUBS 0.027855f
C1029 VTAIL.n269 VSUBS 0.012478f
C1030 VTAIL.n270 VSUBS 0.011785f
C1031 VTAIL.n271 VSUBS 0.021931f
C1032 VTAIL.n272 VSUBS 0.021931f
C1033 VTAIL.n273 VSUBS 0.011785f
C1034 VTAIL.n274 VSUBS 0.012478f
C1035 VTAIL.n275 VSUBS 0.027855f
C1036 VTAIL.n276 VSUBS 0.070606f
C1037 VTAIL.n277 VSUBS 0.012478f
C1038 VTAIL.n278 VSUBS 0.011785f
C1039 VTAIL.n279 VSUBS 0.056386f
C1040 VTAIL.n280 VSUBS 0.035815f
C1041 VTAIL.n281 VSUBS 1.5864f
C1042 VTAIL.n282 VSUBS 0.025029f
C1043 VTAIL.n283 VSUBS 0.021931f
C1044 VTAIL.n284 VSUBS 0.011785f
C1045 VTAIL.n285 VSUBS 0.027855f
C1046 VTAIL.n286 VSUBS 0.012478f
C1047 VTAIL.n287 VSUBS 0.021931f
C1048 VTAIL.n288 VSUBS 0.011785f
C1049 VTAIL.n289 VSUBS 0.027855f
C1050 VTAIL.n290 VSUBS 0.012478f
C1051 VTAIL.n291 VSUBS 0.021931f
C1052 VTAIL.n292 VSUBS 0.011785f
C1053 VTAIL.n293 VSUBS 0.027855f
C1054 VTAIL.n294 VSUBS 0.027855f
C1055 VTAIL.n295 VSUBS 0.012478f
C1056 VTAIL.n296 VSUBS 0.021931f
C1057 VTAIL.n297 VSUBS 0.011785f
C1058 VTAIL.n298 VSUBS 0.027855f
C1059 VTAIL.n299 VSUBS 0.012478f
C1060 VTAIL.n300 VSUBS 0.021931f
C1061 VTAIL.n301 VSUBS 0.011785f
C1062 VTAIL.n302 VSUBS 0.027855f
C1063 VTAIL.n303 VSUBS 0.012478f
C1064 VTAIL.n304 VSUBS 0.021931f
C1065 VTAIL.n305 VSUBS 0.011785f
C1066 VTAIL.n306 VSUBS 0.027855f
C1067 VTAIL.n307 VSUBS 0.012478f
C1068 VTAIL.n308 VSUBS 0.021931f
C1069 VTAIL.n309 VSUBS 0.011785f
C1070 VTAIL.n310 VSUBS 0.027855f
C1071 VTAIL.n311 VSUBS 0.012478f
C1072 VTAIL.n312 VSUBS 0.16747f
C1073 VTAIL.t0 VSUBS 0.059741f
C1074 VTAIL.n313 VSUBS 0.020892f
C1075 VTAIL.n314 VSUBS 0.01772f
C1076 VTAIL.n315 VSUBS 0.011785f
C1077 VTAIL.n316 VSUBS 1.5985f
C1078 VTAIL.n317 VSUBS 0.021931f
C1079 VTAIL.n318 VSUBS 0.011785f
C1080 VTAIL.n319 VSUBS 0.012478f
C1081 VTAIL.n320 VSUBS 0.027855f
C1082 VTAIL.n321 VSUBS 0.027855f
C1083 VTAIL.n322 VSUBS 0.012478f
C1084 VTAIL.n323 VSUBS 0.011785f
C1085 VTAIL.n324 VSUBS 0.021931f
C1086 VTAIL.n325 VSUBS 0.021931f
C1087 VTAIL.n326 VSUBS 0.011785f
C1088 VTAIL.n327 VSUBS 0.012478f
C1089 VTAIL.n328 VSUBS 0.027855f
C1090 VTAIL.n329 VSUBS 0.027855f
C1091 VTAIL.n330 VSUBS 0.012478f
C1092 VTAIL.n331 VSUBS 0.011785f
C1093 VTAIL.n332 VSUBS 0.021931f
C1094 VTAIL.n333 VSUBS 0.021931f
C1095 VTAIL.n334 VSUBS 0.011785f
C1096 VTAIL.n335 VSUBS 0.012478f
C1097 VTAIL.n336 VSUBS 0.027855f
C1098 VTAIL.n337 VSUBS 0.027855f
C1099 VTAIL.n338 VSUBS 0.012478f
C1100 VTAIL.n339 VSUBS 0.011785f
C1101 VTAIL.n340 VSUBS 0.021931f
C1102 VTAIL.n341 VSUBS 0.021931f
C1103 VTAIL.n342 VSUBS 0.011785f
C1104 VTAIL.n343 VSUBS 0.012478f
C1105 VTAIL.n344 VSUBS 0.027855f
C1106 VTAIL.n345 VSUBS 0.027855f
C1107 VTAIL.n346 VSUBS 0.012478f
C1108 VTAIL.n347 VSUBS 0.011785f
C1109 VTAIL.n348 VSUBS 0.021931f
C1110 VTAIL.n349 VSUBS 0.021931f
C1111 VTAIL.n350 VSUBS 0.011785f
C1112 VTAIL.n351 VSUBS 0.012478f
C1113 VTAIL.n352 VSUBS 0.027855f
C1114 VTAIL.n353 VSUBS 0.027855f
C1115 VTAIL.n354 VSUBS 0.012478f
C1116 VTAIL.n355 VSUBS 0.011785f
C1117 VTAIL.n356 VSUBS 0.021931f
C1118 VTAIL.n357 VSUBS 0.021931f
C1119 VTAIL.n358 VSUBS 0.011785f
C1120 VTAIL.n359 VSUBS 0.012132f
C1121 VTAIL.n360 VSUBS 0.012132f
C1122 VTAIL.n361 VSUBS 0.027855f
C1123 VTAIL.n362 VSUBS 0.027855f
C1124 VTAIL.n363 VSUBS 0.012478f
C1125 VTAIL.n364 VSUBS 0.011785f
C1126 VTAIL.n365 VSUBS 0.021931f
C1127 VTAIL.n366 VSUBS 0.021931f
C1128 VTAIL.n367 VSUBS 0.011785f
C1129 VTAIL.n368 VSUBS 0.012478f
C1130 VTAIL.n369 VSUBS 0.027855f
C1131 VTAIL.n370 VSUBS 0.070606f
C1132 VTAIL.n371 VSUBS 0.012478f
C1133 VTAIL.n372 VSUBS 0.011785f
C1134 VTAIL.n373 VSUBS 0.056386f
C1135 VTAIL.n374 VSUBS 0.035815f
C1136 VTAIL.n375 VSUBS 1.5864f
C1137 VTAIL.n376 VSUBS 0.025029f
C1138 VTAIL.n377 VSUBS 0.021931f
C1139 VTAIL.n378 VSUBS 0.011785f
C1140 VTAIL.n379 VSUBS 0.027855f
C1141 VTAIL.n380 VSUBS 0.012478f
C1142 VTAIL.n381 VSUBS 0.021931f
C1143 VTAIL.n382 VSUBS 0.011785f
C1144 VTAIL.n383 VSUBS 0.027855f
C1145 VTAIL.n384 VSUBS 0.012478f
C1146 VTAIL.n385 VSUBS 0.021931f
C1147 VTAIL.n386 VSUBS 0.011785f
C1148 VTAIL.n387 VSUBS 0.027855f
C1149 VTAIL.n388 VSUBS 0.027855f
C1150 VTAIL.n389 VSUBS 0.012478f
C1151 VTAIL.n390 VSUBS 0.021931f
C1152 VTAIL.n391 VSUBS 0.011785f
C1153 VTAIL.n392 VSUBS 0.027855f
C1154 VTAIL.n393 VSUBS 0.012478f
C1155 VTAIL.n394 VSUBS 0.021931f
C1156 VTAIL.n395 VSUBS 0.011785f
C1157 VTAIL.n396 VSUBS 0.027855f
C1158 VTAIL.n397 VSUBS 0.012478f
C1159 VTAIL.n398 VSUBS 0.021931f
C1160 VTAIL.n399 VSUBS 0.011785f
C1161 VTAIL.n400 VSUBS 0.027855f
C1162 VTAIL.n401 VSUBS 0.012478f
C1163 VTAIL.n402 VSUBS 0.021931f
C1164 VTAIL.n403 VSUBS 0.011785f
C1165 VTAIL.n404 VSUBS 0.027855f
C1166 VTAIL.n405 VSUBS 0.012478f
C1167 VTAIL.n406 VSUBS 0.16747f
C1168 VTAIL.t2 VSUBS 0.059741f
C1169 VTAIL.n407 VSUBS 0.020892f
C1170 VTAIL.n408 VSUBS 0.01772f
C1171 VTAIL.n409 VSUBS 0.011785f
C1172 VTAIL.n410 VSUBS 1.5985f
C1173 VTAIL.n411 VSUBS 0.021931f
C1174 VTAIL.n412 VSUBS 0.011785f
C1175 VTAIL.n413 VSUBS 0.012478f
C1176 VTAIL.n414 VSUBS 0.027855f
C1177 VTAIL.n415 VSUBS 0.027855f
C1178 VTAIL.n416 VSUBS 0.012478f
C1179 VTAIL.n417 VSUBS 0.011785f
C1180 VTAIL.n418 VSUBS 0.021931f
C1181 VTAIL.n419 VSUBS 0.021931f
C1182 VTAIL.n420 VSUBS 0.011785f
C1183 VTAIL.n421 VSUBS 0.012478f
C1184 VTAIL.n422 VSUBS 0.027855f
C1185 VTAIL.n423 VSUBS 0.027855f
C1186 VTAIL.n424 VSUBS 0.012478f
C1187 VTAIL.n425 VSUBS 0.011785f
C1188 VTAIL.n426 VSUBS 0.021931f
C1189 VTAIL.n427 VSUBS 0.021931f
C1190 VTAIL.n428 VSUBS 0.011785f
C1191 VTAIL.n429 VSUBS 0.012478f
C1192 VTAIL.n430 VSUBS 0.027855f
C1193 VTAIL.n431 VSUBS 0.027855f
C1194 VTAIL.n432 VSUBS 0.012478f
C1195 VTAIL.n433 VSUBS 0.011785f
C1196 VTAIL.n434 VSUBS 0.021931f
C1197 VTAIL.n435 VSUBS 0.021931f
C1198 VTAIL.n436 VSUBS 0.011785f
C1199 VTAIL.n437 VSUBS 0.012478f
C1200 VTAIL.n438 VSUBS 0.027855f
C1201 VTAIL.n439 VSUBS 0.027855f
C1202 VTAIL.n440 VSUBS 0.012478f
C1203 VTAIL.n441 VSUBS 0.011785f
C1204 VTAIL.n442 VSUBS 0.021931f
C1205 VTAIL.n443 VSUBS 0.021931f
C1206 VTAIL.n444 VSUBS 0.011785f
C1207 VTAIL.n445 VSUBS 0.012478f
C1208 VTAIL.n446 VSUBS 0.027855f
C1209 VTAIL.n447 VSUBS 0.027855f
C1210 VTAIL.n448 VSUBS 0.012478f
C1211 VTAIL.n449 VSUBS 0.011785f
C1212 VTAIL.n450 VSUBS 0.021931f
C1213 VTAIL.n451 VSUBS 0.021931f
C1214 VTAIL.n452 VSUBS 0.011785f
C1215 VTAIL.n453 VSUBS 0.012132f
C1216 VTAIL.n454 VSUBS 0.012132f
C1217 VTAIL.n455 VSUBS 0.027855f
C1218 VTAIL.n456 VSUBS 0.027855f
C1219 VTAIL.n457 VSUBS 0.012478f
C1220 VTAIL.n458 VSUBS 0.011785f
C1221 VTAIL.n459 VSUBS 0.021931f
C1222 VTAIL.n460 VSUBS 0.021931f
C1223 VTAIL.n461 VSUBS 0.011785f
C1224 VTAIL.n462 VSUBS 0.012478f
C1225 VTAIL.n463 VSUBS 0.027855f
C1226 VTAIL.n464 VSUBS 0.070606f
C1227 VTAIL.n465 VSUBS 0.012478f
C1228 VTAIL.n466 VSUBS 0.011785f
C1229 VTAIL.n467 VSUBS 0.056386f
C1230 VTAIL.n468 VSUBS 0.035815f
C1231 VTAIL.n469 VSUBS 0.170903f
C1232 VTAIL.n470 VSUBS 0.025029f
C1233 VTAIL.n471 VSUBS 0.021931f
C1234 VTAIL.n472 VSUBS 0.011785f
C1235 VTAIL.n473 VSUBS 0.027855f
C1236 VTAIL.n474 VSUBS 0.012478f
C1237 VTAIL.n475 VSUBS 0.021931f
C1238 VTAIL.n476 VSUBS 0.011785f
C1239 VTAIL.n477 VSUBS 0.027855f
C1240 VTAIL.n478 VSUBS 0.012478f
C1241 VTAIL.n479 VSUBS 0.021931f
C1242 VTAIL.n480 VSUBS 0.011785f
C1243 VTAIL.n481 VSUBS 0.027855f
C1244 VTAIL.n482 VSUBS 0.027855f
C1245 VTAIL.n483 VSUBS 0.012478f
C1246 VTAIL.n484 VSUBS 0.021931f
C1247 VTAIL.n485 VSUBS 0.011785f
C1248 VTAIL.n486 VSUBS 0.027855f
C1249 VTAIL.n487 VSUBS 0.012478f
C1250 VTAIL.n488 VSUBS 0.021931f
C1251 VTAIL.n489 VSUBS 0.011785f
C1252 VTAIL.n490 VSUBS 0.027855f
C1253 VTAIL.n491 VSUBS 0.012478f
C1254 VTAIL.n492 VSUBS 0.021931f
C1255 VTAIL.n493 VSUBS 0.011785f
C1256 VTAIL.n494 VSUBS 0.027855f
C1257 VTAIL.n495 VSUBS 0.012478f
C1258 VTAIL.n496 VSUBS 0.021931f
C1259 VTAIL.n497 VSUBS 0.011785f
C1260 VTAIL.n498 VSUBS 0.027855f
C1261 VTAIL.n499 VSUBS 0.012478f
C1262 VTAIL.n500 VSUBS 0.16747f
C1263 VTAIL.t5 VSUBS 0.059741f
C1264 VTAIL.n501 VSUBS 0.020892f
C1265 VTAIL.n502 VSUBS 0.01772f
C1266 VTAIL.n503 VSUBS 0.011785f
C1267 VTAIL.n504 VSUBS 1.5985f
C1268 VTAIL.n505 VSUBS 0.021931f
C1269 VTAIL.n506 VSUBS 0.011785f
C1270 VTAIL.n507 VSUBS 0.012478f
C1271 VTAIL.n508 VSUBS 0.027855f
C1272 VTAIL.n509 VSUBS 0.027855f
C1273 VTAIL.n510 VSUBS 0.012478f
C1274 VTAIL.n511 VSUBS 0.011785f
C1275 VTAIL.n512 VSUBS 0.021931f
C1276 VTAIL.n513 VSUBS 0.021931f
C1277 VTAIL.n514 VSUBS 0.011785f
C1278 VTAIL.n515 VSUBS 0.012478f
C1279 VTAIL.n516 VSUBS 0.027855f
C1280 VTAIL.n517 VSUBS 0.027855f
C1281 VTAIL.n518 VSUBS 0.012478f
C1282 VTAIL.n519 VSUBS 0.011785f
C1283 VTAIL.n520 VSUBS 0.021931f
C1284 VTAIL.n521 VSUBS 0.021931f
C1285 VTAIL.n522 VSUBS 0.011785f
C1286 VTAIL.n523 VSUBS 0.012478f
C1287 VTAIL.n524 VSUBS 0.027855f
C1288 VTAIL.n525 VSUBS 0.027855f
C1289 VTAIL.n526 VSUBS 0.012478f
C1290 VTAIL.n527 VSUBS 0.011785f
C1291 VTAIL.n528 VSUBS 0.021931f
C1292 VTAIL.n529 VSUBS 0.021931f
C1293 VTAIL.n530 VSUBS 0.011785f
C1294 VTAIL.n531 VSUBS 0.012478f
C1295 VTAIL.n532 VSUBS 0.027855f
C1296 VTAIL.n533 VSUBS 0.027855f
C1297 VTAIL.n534 VSUBS 0.012478f
C1298 VTAIL.n535 VSUBS 0.011785f
C1299 VTAIL.n536 VSUBS 0.021931f
C1300 VTAIL.n537 VSUBS 0.021931f
C1301 VTAIL.n538 VSUBS 0.011785f
C1302 VTAIL.n539 VSUBS 0.012478f
C1303 VTAIL.n540 VSUBS 0.027855f
C1304 VTAIL.n541 VSUBS 0.027855f
C1305 VTAIL.n542 VSUBS 0.012478f
C1306 VTAIL.n543 VSUBS 0.011785f
C1307 VTAIL.n544 VSUBS 0.021931f
C1308 VTAIL.n545 VSUBS 0.021931f
C1309 VTAIL.n546 VSUBS 0.011785f
C1310 VTAIL.n547 VSUBS 0.012132f
C1311 VTAIL.n548 VSUBS 0.012132f
C1312 VTAIL.n549 VSUBS 0.027855f
C1313 VTAIL.n550 VSUBS 0.027855f
C1314 VTAIL.n551 VSUBS 0.012478f
C1315 VTAIL.n552 VSUBS 0.011785f
C1316 VTAIL.n553 VSUBS 0.021931f
C1317 VTAIL.n554 VSUBS 0.021931f
C1318 VTAIL.n555 VSUBS 0.011785f
C1319 VTAIL.n556 VSUBS 0.012478f
C1320 VTAIL.n557 VSUBS 0.027855f
C1321 VTAIL.n558 VSUBS 0.070606f
C1322 VTAIL.n559 VSUBS 0.012478f
C1323 VTAIL.n560 VSUBS 0.011785f
C1324 VTAIL.n561 VSUBS 0.056386f
C1325 VTAIL.n562 VSUBS 0.035815f
C1326 VTAIL.n563 VSUBS 0.170903f
C1327 VTAIL.n564 VSUBS 0.025029f
C1328 VTAIL.n565 VSUBS 0.021931f
C1329 VTAIL.n566 VSUBS 0.011785f
C1330 VTAIL.n567 VSUBS 0.027855f
C1331 VTAIL.n568 VSUBS 0.012478f
C1332 VTAIL.n569 VSUBS 0.021931f
C1333 VTAIL.n570 VSUBS 0.011785f
C1334 VTAIL.n571 VSUBS 0.027855f
C1335 VTAIL.n572 VSUBS 0.012478f
C1336 VTAIL.n573 VSUBS 0.021931f
C1337 VTAIL.n574 VSUBS 0.011785f
C1338 VTAIL.n575 VSUBS 0.027855f
C1339 VTAIL.n576 VSUBS 0.027855f
C1340 VTAIL.n577 VSUBS 0.012478f
C1341 VTAIL.n578 VSUBS 0.021931f
C1342 VTAIL.n579 VSUBS 0.011785f
C1343 VTAIL.n580 VSUBS 0.027855f
C1344 VTAIL.n581 VSUBS 0.012478f
C1345 VTAIL.n582 VSUBS 0.021931f
C1346 VTAIL.n583 VSUBS 0.011785f
C1347 VTAIL.n584 VSUBS 0.027855f
C1348 VTAIL.n585 VSUBS 0.012478f
C1349 VTAIL.n586 VSUBS 0.021931f
C1350 VTAIL.n587 VSUBS 0.011785f
C1351 VTAIL.n588 VSUBS 0.027855f
C1352 VTAIL.n589 VSUBS 0.012478f
C1353 VTAIL.n590 VSUBS 0.021931f
C1354 VTAIL.n591 VSUBS 0.011785f
C1355 VTAIL.n592 VSUBS 0.027855f
C1356 VTAIL.n593 VSUBS 0.012478f
C1357 VTAIL.n594 VSUBS 0.16747f
C1358 VTAIL.t6 VSUBS 0.059741f
C1359 VTAIL.n595 VSUBS 0.020892f
C1360 VTAIL.n596 VSUBS 0.01772f
C1361 VTAIL.n597 VSUBS 0.011785f
C1362 VTAIL.n598 VSUBS 1.5985f
C1363 VTAIL.n599 VSUBS 0.021931f
C1364 VTAIL.n600 VSUBS 0.011785f
C1365 VTAIL.n601 VSUBS 0.012478f
C1366 VTAIL.n602 VSUBS 0.027855f
C1367 VTAIL.n603 VSUBS 0.027855f
C1368 VTAIL.n604 VSUBS 0.012478f
C1369 VTAIL.n605 VSUBS 0.011785f
C1370 VTAIL.n606 VSUBS 0.021931f
C1371 VTAIL.n607 VSUBS 0.021931f
C1372 VTAIL.n608 VSUBS 0.011785f
C1373 VTAIL.n609 VSUBS 0.012478f
C1374 VTAIL.n610 VSUBS 0.027855f
C1375 VTAIL.n611 VSUBS 0.027855f
C1376 VTAIL.n612 VSUBS 0.012478f
C1377 VTAIL.n613 VSUBS 0.011785f
C1378 VTAIL.n614 VSUBS 0.021931f
C1379 VTAIL.n615 VSUBS 0.021931f
C1380 VTAIL.n616 VSUBS 0.011785f
C1381 VTAIL.n617 VSUBS 0.012478f
C1382 VTAIL.n618 VSUBS 0.027855f
C1383 VTAIL.n619 VSUBS 0.027855f
C1384 VTAIL.n620 VSUBS 0.012478f
C1385 VTAIL.n621 VSUBS 0.011785f
C1386 VTAIL.n622 VSUBS 0.021931f
C1387 VTAIL.n623 VSUBS 0.021931f
C1388 VTAIL.n624 VSUBS 0.011785f
C1389 VTAIL.n625 VSUBS 0.012478f
C1390 VTAIL.n626 VSUBS 0.027855f
C1391 VTAIL.n627 VSUBS 0.027855f
C1392 VTAIL.n628 VSUBS 0.012478f
C1393 VTAIL.n629 VSUBS 0.011785f
C1394 VTAIL.n630 VSUBS 0.021931f
C1395 VTAIL.n631 VSUBS 0.021931f
C1396 VTAIL.n632 VSUBS 0.011785f
C1397 VTAIL.n633 VSUBS 0.012478f
C1398 VTAIL.n634 VSUBS 0.027855f
C1399 VTAIL.n635 VSUBS 0.027855f
C1400 VTAIL.n636 VSUBS 0.012478f
C1401 VTAIL.n637 VSUBS 0.011785f
C1402 VTAIL.n638 VSUBS 0.021931f
C1403 VTAIL.n639 VSUBS 0.021931f
C1404 VTAIL.n640 VSUBS 0.011785f
C1405 VTAIL.n641 VSUBS 0.012132f
C1406 VTAIL.n642 VSUBS 0.012132f
C1407 VTAIL.n643 VSUBS 0.027855f
C1408 VTAIL.n644 VSUBS 0.027855f
C1409 VTAIL.n645 VSUBS 0.012478f
C1410 VTAIL.n646 VSUBS 0.011785f
C1411 VTAIL.n647 VSUBS 0.021931f
C1412 VTAIL.n648 VSUBS 0.021931f
C1413 VTAIL.n649 VSUBS 0.011785f
C1414 VTAIL.n650 VSUBS 0.012478f
C1415 VTAIL.n651 VSUBS 0.027855f
C1416 VTAIL.n652 VSUBS 0.070606f
C1417 VTAIL.n653 VSUBS 0.012478f
C1418 VTAIL.n654 VSUBS 0.011785f
C1419 VTAIL.n655 VSUBS 0.056386f
C1420 VTAIL.n656 VSUBS 0.035815f
C1421 VTAIL.n657 VSUBS 1.5864f
C1422 VTAIL.n658 VSUBS 0.025029f
C1423 VTAIL.n659 VSUBS 0.021931f
C1424 VTAIL.n660 VSUBS 0.011785f
C1425 VTAIL.n661 VSUBS 0.027855f
C1426 VTAIL.n662 VSUBS 0.012478f
C1427 VTAIL.n663 VSUBS 0.021931f
C1428 VTAIL.n664 VSUBS 0.011785f
C1429 VTAIL.n665 VSUBS 0.027855f
C1430 VTAIL.n666 VSUBS 0.012478f
C1431 VTAIL.n667 VSUBS 0.021931f
C1432 VTAIL.n668 VSUBS 0.011785f
C1433 VTAIL.n669 VSUBS 0.027855f
C1434 VTAIL.n670 VSUBS 0.012478f
C1435 VTAIL.n671 VSUBS 0.021931f
C1436 VTAIL.n672 VSUBS 0.011785f
C1437 VTAIL.n673 VSUBS 0.027855f
C1438 VTAIL.n674 VSUBS 0.012478f
C1439 VTAIL.n675 VSUBS 0.021931f
C1440 VTAIL.n676 VSUBS 0.011785f
C1441 VTAIL.n677 VSUBS 0.027855f
C1442 VTAIL.n678 VSUBS 0.012478f
C1443 VTAIL.n679 VSUBS 0.021931f
C1444 VTAIL.n680 VSUBS 0.011785f
C1445 VTAIL.n681 VSUBS 0.027855f
C1446 VTAIL.n682 VSUBS 0.012478f
C1447 VTAIL.n683 VSUBS 0.021931f
C1448 VTAIL.n684 VSUBS 0.011785f
C1449 VTAIL.n685 VSUBS 0.027855f
C1450 VTAIL.n686 VSUBS 0.012478f
C1451 VTAIL.n687 VSUBS 0.16747f
C1452 VTAIL.t3 VSUBS 0.059741f
C1453 VTAIL.n688 VSUBS 0.020892f
C1454 VTAIL.n689 VSUBS 0.01772f
C1455 VTAIL.n690 VSUBS 0.011785f
C1456 VTAIL.n691 VSUBS 1.5985f
C1457 VTAIL.n692 VSUBS 0.021931f
C1458 VTAIL.n693 VSUBS 0.011785f
C1459 VTAIL.n694 VSUBS 0.012478f
C1460 VTAIL.n695 VSUBS 0.027855f
C1461 VTAIL.n696 VSUBS 0.027855f
C1462 VTAIL.n697 VSUBS 0.012478f
C1463 VTAIL.n698 VSUBS 0.011785f
C1464 VTAIL.n699 VSUBS 0.021931f
C1465 VTAIL.n700 VSUBS 0.021931f
C1466 VTAIL.n701 VSUBS 0.011785f
C1467 VTAIL.n702 VSUBS 0.012478f
C1468 VTAIL.n703 VSUBS 0.027855f
C1469 VTAIL.n704 VSUBS 0.027855f
C1470 VTAIL.n705 VSUBS 0.012478f
C1471 VTAIL.n706 VSUBS 0.011785f
C1472 VTAIL.n707 VSUBS 0.021931f
C1473 VTAIL.n708 VSUBS 0.021931f
C1474 VTAIL.n709 VSUBS 0.011785f
C1475 VTAIL.n710 VSUBS 0.012478f
C1476 VTAIL.n711 VSUBS 0.027855f
C1477 VTAIL.n712 VSUBS 0.027855f
C1478 VTAIL.n713 VSUBS 0.012478f
C1479 VTAIL.n714 VSUBS 0.011785f
C1480 VTAIL.n715 VSUBS 0.021931f
C1481 VTAIL.n716 VSUBS 0.021931f
C1482 VTAIL.n717 VSUBS 0.011785f
C1483 VTAIL.n718 VSUBS 0.012478f
C1484 VTAIL.n719 VSUBS 0.027855f
C1485 VTAIL.n720 VSUBS 0.027855f
C1486 VTAIL.n721 VSUBS 0.012478f
C1487 VTAIL.n722 VSUBS 0.011785f
C1488 VTAIL.n723 VSUBS 0.021931f
C1489 VTAIL.n724 VSUBS 0.021931f
C1490 VTAIL.n725 VSUBS 0.011785f
C1491 VTAIL.n726 VSUBS 0.012478f
C1492 VTAIL.n727 VSUBS 0.027855f
C1493 VTAIL.n728 VSUBS 0.027855f
C1494 VTAIL.n729 VSUBS 0.027855f
C1495 VTAIL.n730 VSUBS 0.012478f
C1496 VTAIL.n731 VSUBS 0.011785f
C1497 VTAIL.n732 VSUBS 0.021931f
C1498 VTAIL.n733 VSUBS 0.021931f
C1499 VTAIL.n734 VSUBS 0.011785f
C1500 VTAIL.n735 VSUBS 0.012132f
C1501 VTAIL.n736 VSUBS 0.012132f
C1502 VTAIL.n737 VSUBS 0.027855f
C1503 VTAIL.n738 VSUBS 0.027855f
C1504 VTAIL.n739 VSUBS 0.012478f
C1505 VTAIL.n740 VSUBS 0.011785f
C1506 VTAIL.n741 VSUBS 0.021931f
C1507 VTAIL.n742 VSUBS 0.021931f
C1508 VTAIL.n743 VSUBS 0.011785f
C1509 VTAIL.n744 VSUBS 0.012478f
C1510 VTAIL.n745 VSUBS 0.027855f
C1511 VTAIL.n746 VSUBS 0.070606f
C1512 VTAIL.n747 VSUBS 0.012478f
C1513 VTAIL.n748 VSUBS 0.011785f
C1514 VTAIL.n749 VSUBS 0.056386f
C1515 VTAIL.n750 VSUBS 0.035815f
C1516 VTAIL.n751 VSUBS 1.52442f
C1517 VDD1.t1 VSUBS 0.3601f
C1518 VDD1.t3 VSUBS 0.3601f
C1519 VDD1.n0 VSUBS 2.98645f
C1520 VDD1.t0 VSUBS 0.3601f
C1521 VDD1.t2 VSUBS 0.3601f
C1522 VDD1.n1 VSUBS 3.84043f
C1523 VP.n0 VSUBS 0.040985f
C1524 VP.t3 VSUBS 3.00365f
C1525 VP.n1 VSUBS 0.05983f
C1526 VP.t2 VSUBS 3.15799f
C1527 VP.t1 VSUBS 3.15664f
C1528 VP.n2 VSUBS 3.98839f
C1529 VP.n3 VSUBS 2.54234f
C1530 VP.t0 VSUBS 3.00365f
C1531 VP.n4 VSUBS 1.14765f
C1532 VP.n5 VSUBS 0.053758f
C1533 VP.n6 VSUBS 0.040985f
C1534 VP.n7 VSUBS 0.040985f
C1535 VP.n8 VSUBS 0.040985f
C1536 VP.n9 VSUBS 0.05983f
C1537 VP.n10 VSUBS 0.053758f
C1538 VP.n11 VSUBS 1.14765f
C1539 VP.n12 VSUBS 0.039832f
.ends

