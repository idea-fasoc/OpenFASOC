* NGSPICE file created from diff_pair_sample_0094.ext - technology: sky130A

.subckt diff_pair_sample_0094 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=7.6947 pd=40.24 as=3.25545 ps=20.06 w=19.73 l=3.56
X1 VDD1.t3 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.25545 pd=20.06 as=7.6947 ps=40.24 w=19.73 l=3.56
X2 VDD1.t2 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.25545 pd=20.06 as=7.6947 ps=40.24 w=19.73 l=3.56
X3 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=7.6947 pd=40.24 as=0 ps=0 w=19.73 l=3.56
X4 VDD2.t1 VN.t1 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=3.25545 pd=20.06 as=7.6947 ps=40.24 w=19.73 l=3.56
X5 VTAIL.t5 VN.t2 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=7.6947 pd=40.24 as=3.25545 ps=20.06 w=19.73 l=3.56
X6 VTAIL.t3 VP.t2 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=7.6947 pd=40.24 as=3.25545 ps=20.06 w=19.73 l=3.56
X7 VTAIL.t0 VP.t3 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=7.6947 pd=40.24 as=3.25545 ps=20.06 w=19.73 l=3.56
X8 VDD2.t3 VN.t3 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=3.25545 pd=20.06 as=7.6947 ps=40.24 w=19.73 l=3.56
X9 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=7.6947 pd=40.24 as=0 ps=0 w=19.73 l=3.56
X10 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=7.6947 pd=40.24 as=0 ps=0 w=19.73 l=3.56
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.6947 pd=40.24 as=0 ps=0 w=19.73 l=3.56
R0 VN.n1 VN.t3 168.275
R1 VN.n0 VN.t0 168.275
R2 VN.n0 VN.t1 167.041
R3 VN.n1 VN.t2 167.041
R4 VN VN.n1 57.4841
R5 VN VN.n0 2.13941
R6 VDD2.n2 VDD2.n0 111.959
R7 VDD2.n2 VDD2.n1 61.1744
R8 VDD2.n1 VDD2.t0 1.00405
R9 VDD2.n1 VDD2.t3 1.00405
R10 VDD2.n0 VDD2.t2 1.00405
R11 VDD2.n0 VDD2.t1 1.00405
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t3 45.4993
R14 VTAIL.n4 VTAIL.t4 45.4993
R15 VTAIL.n3 VTAIL.t5 45.4993
R16 VTAIL.n6 VTAIL.t1 45.4991
R17 VTAIL.n7 VTAIL.t6 45.4991
R18 VTAIL.n0 VTAIL.t7 45.4991
R19 VTAIL.n1 VTAIL.t2 45.4991
R20 VTAIL.n2 VTAIL.t0 45.4991
R21 VTAIL.n7 VTAIL.n6 32.729
R22 VTAIL.n3 VTAIL.n2 32.729
R23 VTAIL.n4 VTAIL.n3 3.35395
R24 VTAIL.n6 VTAIL.n5 3.35395
R25 VTAIL.n2 VTAIL.n1 3.35395
R26 VTAIL VTAIL.n0 1.73541
R27 VTAIL VTAIL.n7 1.61903
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 B.n768 B.n767 585
R31 B.n770 B.n153 585
R32 B.n773 B.n772 585
R33 B.n774 B.n152 585
R34 B.n776 B.n775 585
R35 B.n778 B.n151 585
R36 B.n781 B.n780 585
R37 B.n782 B.n150 585
R38 B.n784 B.n783 585
R39 B.n786 B.n149 585
R40 B.n789 B.n788 585
R41 B.n790 B.n148 585
R42 B.n792 B.n791 585
R43 B.n794 B.n147 585
R44 B.n797 B.n796 585
R45 B.n798 B.n146 585
R46 B.n800 B.n799 585
R47 B.n802 B.n145 585
R48 B.n805 B.n804 585
R49 B.n806 B.n144 585
R50 B.n808 B.n807 585
R51 B.n810 B.n143 585
R52 B.n813 B.n812 585
R53 B.n814 B.n142 585
R54 B.n816 B.n815 585
R55 B.n818 B.n141 585
R56 B.n821 B.n820 585
R57 B.n822 B.n140 585
R58 B.n824 B.n823 585
R59 B.n826 B.n139 585
R60 B.n829 B.n828 585
R61 B.n830 B.n138 585
R62 B.n832 B.n831 585
R63 B.n834 B.n137 585
R64 B.n837 B.n836 585
R65 B.n838 B.n136 585
R66 B.n840 B.n839 585
R67 B.n842 B.n135 585
R68 B.n845 B.n844 585
R69 B.n846 B.n134 585
R70 B.n848 B.n847 585
R71 B.n850 B.n133 585
R72 B.n853 B.n852 585
R73 B.n854 B.n132 585
R74 B.n856 B.n855 585
R75 B.n858 B.n131 585
R76 B.n861 B.n860 585
R77 B.n862 B.n130 585
R78 B.n864 B.n863 585
R79 B.n866 B.n129 585
R80 B.n869 B.n868 585
R81 B.n870 B.n128 585
R82 B.n872 B.n871 585
R83 B.n874 B.n127 585
R84 B.n877 B.n876 585
R85 B.n878 B.n126 585
R86 B.n880 B.n879 585
R87 B.n882 B.n125 585
R88 B.n885 B.n884 585
R89 B.n886 B.n124 585
R90 B.n888 B.n887 585
R91 B.n890 B.n123 585
R92 B.n892 B.n891 585
R93 B.n894 B.n893 585
R94 B.n897 B.n896 585
R95 B.n898 B.n118 585
R96 B.n900 B.n899 585
R97 B.n902 B.n117 585
R98 B.n905 B.n904 585
R99 B.n906 B.n116 585
R100 B.n908 B.n907 585
R101 B.n910 B.n115 585
R102 B.n913 B.n912 585
R103 B.n914 B.n112 585
R104 B.n917 B.n916 585
R105 B.n919 B.n111 585
R106 B.n922 B.n921 585
R107 B.n923 B.n110 585
R108 B.n925 B.n924 585
R109 B.n927 B.n109 585
R110 B.n930 B.n929 585
R111 B.n931 B.n108 585
R112 B.n933 B.n932 585
R113 B.n935 B.n107 585
R114 B.n938 B.n937 585
R115 B.n939 B.n106 585
R116 B.n941 B.n940 585
R117 B.n943 B.n105 585
R118 B.n946 B.n945 585
R119 B.n947 B.n104 585
R120 B.n949 B.n948 585
R121 B.n951 B.n103 585
R122 B.n954 B.n953 585
R123 B.n955 B.n102 585
R124 B.n957 B.n956 585
R125 B.n959 B.n101 585
R126 B.n962 B.n961 585
R127 B.n963 B.n100 585
R128 B.n965 B.n964 585
R129 B.n967 B.n99 585
R130 B.n970 B.n969 585
R131 B.n971 B.n98 585
R132 B.n973 B.n972 585
R133 B.n975 B.n97 585
R134 B.n978 B.n977 585
R135 B.n979 B.n96 585
R136 B.n981 B.n980 585
R137 B.n983 B.n95 585
R138 B.n986 B.n985 585
R139 B.n987 B.n94 585
R140 B.n989 B.n988 585
R141 B.n991 B.n93 585
R142 B.n994 B.n993 585
R143 B.n995 B.n92 585
R144 B.n997 B.n996 585
R145 B.n999 B.n91 585
R146 B.n1002 B.n1001 585
R147 B.n1003 B.n90 585
R148 B.n1005 B.n1004 585
R149 B.n1007 B.n89 585
R150 B.n1010 B.n1009 585
R151 B.n1011 B.n88 585
R152 B.n1013 B.n1012 585
R153 B.n1015 B.n87 585
R154 B.n1018 B.n1017 585
R155 B.n1019 B.n86 585
R156 B.n1021 B.n1020 585
R157 B.n1023 B.n85 585
R158 B.n1026 B.n1025 585
R159 B.n1027 B.n84 585
R160 B.n1029 B.n1028 585
R161 B.n1031 B.n83 585
R162 B.n1034 B.n1033 585
R163 B.n1035 B.n82 585
R164 B.n1037 B.n1036 585
R165 B.n1039 B.n81 585
R166 B.n1042 B.n1041 585
R167 B.n1043 B.n80 585
R168 B.n766 B.n78 585
R169 B.n1046 B.n78 585
R170 B.n765 B.n77 585
R171 B.n1047 B.n77 585
R172 B.n764 B.n76 585
R173 B.n1048 B.n76 585
R174 B.n763 B.n762 585
R175 B.n762 B.n72 585
R176 B.n761 B.n71 585
R177 B.n1054 B.n71 585
R178 B.n760 B.n70 585
R179 B.n1055 B.n70 585
R180 B.n759 B.n69 585
R181 B.n1056 B.n69 585
R182 B.n758 B.n757 585
R183 B.n757 B.n65 585
R184 B.n756 B.n64 585
R185 B.n1062 B.n64 585
R186 B.n755 B.n63 585
R187 B.n1063 B.n63 585
R188 B.n754 B.n62 585
R189 B.n1064 B.n62 585
R190 B.n753 B.n752 585
R191 B.n752 B.n58 585
R192 B.n751 B.n57 585
R193 B.n1070 B.n57 585
R194 B.n750 B.n56 585
R195 B.n1071 B.n56 585
R196 B.n749 B.n55 585
R197 B.n1072 B.n55 585
R198 B.n748 B.n747 585
R199 B.n747 B.n51 585
R200 B.n746 B.n50 585
R201 B.n1078 B.n50 585
R202 B.n745 B.n49 585
R203 B.n1079 B.n49 585
R204 B.n744 B.n48 585
R205 B.n1080 B.n48 585
R206 B.n743 B.n742 585
R207 B.n742 B.n44 585
R208 B.n741 B.n43 585
R209 B.n1086 B.n43 585
R210 B.n740 B.n42 585
R211 B.n1087 B.n42 585
R212 B.n739 B.n41 585
R213 B.n1088 B.n41 585
R214 B.n738 B.n737 585
R215 B.n737 B.n40 585
R216 B.n736 B.n36 585
R217 B.n1094 B.n36 585
R218 B.n735 B.n35 585
R219 B.n1095 B.n35 585
R220 B.n734 B.n34 585
R221 B.n1096 B.n34 585
R222 B.n733 B.n732 585
R223 B.n732 B.n30 585
R224 B.n731 B.n29 585
R225 B.n1102 B.n29 585
R226 B.n730 B.n28 585
R227 B.n1103 B.n28 585
R228 B.n729 B.n27 585
R229 B.n1104 B.n27 585
R230 B.n728 B.n727 585
R231 B.n727 B.n23 585
R232 B.n726 B.n22 585
R233 B.n1110 B.n22 585
R234 B.n725 B.n21 585
R235 B.n1111 B.n21 585
R236 B.n724 B.n20 585
R237 B.n1112 B.n20 585
R238 B.n723 B.n722 585
R239 B.n722 B.n19 585
R240 B.n721 B.n15 585
R241 B.n1118 B.n15 585
R242 B.n720 B.n14 585
R243 B.n1119 B.n14 585
R244 B.n719 B.n13 585
R245 B.n1120 B.n13 585
R246 B.n718 B.n717 585
R247 B.n717 B.n12 585
R248 B.n716 B.n715 585
R249 B.n716 B.n8 585
R250 B.n714 B.n7 585
R251 B.n1127 B.n7 585
R252 B.n713 B.n6 585
R253 B.n1128 B.n6 585
R254 B.n712 B.n5 585
R255 B.n1129 B.n5 585
R256 B.n711 B.n710 585
R257 B.n710 B.n4 585
R258 B.n709 B.n154 585
R259 B.n709 B.n708 585
R260 B.n699 B.n155 585
R261 B.n156 B.n155 585
R262 B.n701 B.n700 585
R263 B.n702 B.n701 585
R264 B.n698 B.n161 585
R265 B.n161 B.n160 585
R266 B.n697 B.n696 585
R267 B.n696 B.n695 585
R268 B.n163 B.n162 585
R269 B.n688 B.n163 585
R270 B.n687 B.n686 585
R271 B.n689 B.n687 585
R272 B.n685 B.n168 585
R273 B.n168 B.n167 585
R274 B.n684 B.n683 585
R275 B.n683 B.n682 585
R276 B.n170 B.n169 585
R277 B.n171 B.n170 585
R278 B.n675 B.n674 585
R279 B.n676 B.n675 585
R280 B.n673 B.n176 585
R281 B.n176 B.n175 585
R282 B.n672 B.n671 585
R283 B.n671 B.n670 585
R284 B.n178 B.n177 585
R285 B.n179 B.n178 585
R286 B.n663 B.n662 585
R287 B.n664 B.n663 585
R288 B.n661 B.n184 585
R289 B.n184 B.n183 585
R290 B.n660 B.n659 585
R291 B.n659 B.n658 585
R292 B.n186 B.n185 585
R293 B.n651 B.n186 585
R294 B.n650 B.n649 585
R295 B.n652 B.n650 585
R296 B.n648 B.n191 585
R297 B.n191 B.n190 585
R298 B.n647 B.n646 585
R299 B.n646 B.n645 585
R300 B.n193 B.n192 585
R301 B.n194 B.n193 585
R302 B.n638 B.n637 585
R303 B.n639 B.n638 585
R304 B.n636 B.n199 585
R305 B.n199 B.n198 585
R306 B.n635 B.n634 585
R307 B.n634 B.n633 585
R308 B.n201 B.n200 585
R309 B.n202 B.n201 585
R310 B.n626 B.n625 585
R311 B.n627 B.n626 585
R312 B.n624 B.n207 585
R313 B.n207 B.n206 585
R314 B.n623 B.n622 585
R315 B.n622 B.n621 585
R316 B.n209 B.n208 585
R317 B.n210 B.n209 585
R318 B.n614 B.n613 585
R319 B.n615 B.n614 585
R320 B.n612 B.n214 585
R321 B.n218 B.n214 585
R322 B.n611 B.n610 585
R323 B.n610 B.n609 585
R324 B.n216 B.n215 585
R325 B.n217 B.n216 585
R326 B.n602 B.n601 585
R327 B.n603 B.n602 585
R328 B.n600 B.n223 585
R329 B.n223 B.n222 585
R330 B.n599 B.n598 585
R331 B.n598 B.n597 585
R332 B.n225 B.n224 585
R333 B.n226 B.n225 585
R334 B.n590 B.n589 585
R335 B.n591 B.n590 585
R336 B.n588 B.n231 585
R337 B.n231 B.n230 585
R338 B.n587 B.n586 585
R339 B.n586 B.n585 585
R340 B.n582 B.n235 585
R341 B.n581 B.n580 585
R342 B.n578 B.n236 585
R343 B.n578 B.n234 585
R344 B.n577 B.n576 585
R345 B.n575 B.n574 585
R346 B.n573 B.n238 585
R347 B.n571 B.n570 585
R348 B.n569 B.n239 585
R349 B.n568 B.n567 585
R350 B.n565 B.n240 585
R351 B.n563 B.n562 585
R352 B.n561 B.n241 585
R353 B.n560 B.n559 585
R354 B.n557 B.n242 585
R355 B.n555 B.n554 585
R356 B.n553 B.n243 585
R357 B.n552 B.n551 585
R358 B.n549 B.n244 585
R359 B.n547 B.n546 585
R360 B.n545 B.n245 585
R361 B.n544 B.n543 585
R362 B.n541 B.n246 585
R363 B.n539 B.n538 585
R364 B.n537 B.n247 585
R365 B.n536 B.n535 585
R366 B.n533 B.n248 585
R367 B.n531 B.n530 585
R368 B.n529 B.n249 585
R369 B.n528 B.n527 585
R370 B.n525 B.n250 585
R371 B.n523 B.n522 585
R372 B.n521 B.n251 585
R373 B.n520 B.n519 585
R374 B.n517 B.n252 585
R375 B.n515 B.n514 585
R376 B.n513 B.n253 585
R377 B.n512 B.n511 585
R378 B.n509 B.n254 585
R379 B.n507 B.n506 585
R380 B.n505 B.n255 585
R381 B.n504 B.n503 585
R382 B.n501 B.n256 585
R383 B.n499 B.n498 585
R384 B.n497 B.n257 585
R385 B.n496 B.n495 585
R386 B.n493 B.n258 585
R387 B.n491 B.n490 585
R388 B.n489 B.n259 585
R389 B.n488 B.n487 585
R390 B.n485 B.n260 585
R391 B.n483 B.n482 585
R392 B.n481 B.n261 585
R393 B.n480 B.n479 585
R394 B.n477 B.n262 585
R395 B.n475 B.n474 585
R396 B.n473 B.n263 585
R397 B.n472 B.n471 585
R398 B.n469 B.n264 585
R399 B.n467 B.n466 585
R400 B.n465 B.n265 585
R401 B.n464 B.n463 585
R402 B.n461 B.n266 585
R403 B.n459 B.n458 585
R404 B.n457 B.n267 585
R405 B.n455 B.n454 585
R406 B.n452 B.n270 585
R407 B.n450 B.n449 585
R408 B.n448 B.n271 585
R409 B.n447 B.n446 585
R410 B.n444 B.n272 585
R411 B.n442 B.n441 585
R412 B.n440 B.n273 585
R413 B.n439 B.n438 585
R414 B.n436 B.n274 585
R415 B.n434 B.n433 585
R416 B.n432 B.n275 585
R417 B.n431 B.n430 585
R418 B.n428 B.n279 585
R419 B.n426 B.n425 585
R420 B.n424 B.n280 585
R421 B.n423 B.n422 585
R422 B.n420 B.n281 585
R423 B.n418 B.n417 585
R424 B.n416 B.n282 585
R425 B.n415 B.n414 585
R426 B.n412 B.n283 585
R427 B.n410 B.n409 585
R428 B.n408 B.n284 585
R429 B.n407 B.n406 585
R430 B.n404 B.n285 585
R431 B.n402 B.n401 585
R432 B.n400 B.n286 585
R433 B.n399 B.n398 585
R434 B.n396 B.n287 585
R435 B.n394 B.n393 585
R436 B.n392 B.n288 585
R437 B.n391 B.n390 585
R438 B.n388 B.n289 585
R439 B.n386 B.n385 585
R440 B.n384 B.n290 585
R441 B.n383 B.n382 585
R442 B.n380 B.n291 585
R443 B.n378 B.n377 585
R444 B.n376 B.n292 585
R445 B.n375 B.n374 585
R446 B.n372 B.n293 585
R447 B.n370 B.n369 585
R448 B.n368 B.n294 585
R449 B.n367 B.n366 585
R450 B.n364 B.n295 585
R451 B.n362 B.n361 585
R452 B.n360 B.n296 585
R453 B.n359 B.n358 585
R454 B.n356 B.n297 585
R455 B.n354 B.n353 585
R456 B.n352 B.n298 585
R457 B.n351 B.n350 585
R458 B.n348 B.n299 585
R459 B.n346 B.n345 585
R460 B.n344 B.n300 585
R461 B.n343 B.n342 585
R462 B.n340 B.n301 585
R463 B.n338 B.n337 585
R464 B.n336 B.n302 585
R465 B.n335 B.n334 585
R466 B.n332 B.n303 585
R467 B.n330 B.n329 585
R468 B.n328 B.n304 585
R469 B.n327 B.n326 585
R470 B.n324 B.n305 585
R471 B.n322 B.n321 585
R472 B.n320 B.n306 585
R473 B.n319 B.n318 585
R474 B.n316 B.n307 585
R475 B.n314 B.n313 585
R476 B.n312 B.n308 585
R477 B.n311 B.n310 585
R478 B.n233 B.n232 585
R479 B.n234 B.n233 585
R480 B.n584 B.n583 585
R481 B.n585 B.n584 585
R482 B.n229 B.n228 585
R483 B.n230 B.n229 585
R484 B.n593 B.n592 585
R485 B.n592 B.n591 585
R486 B.n594 B.n227 585
R487 B.n227 B.n226 585
R488 B.n596 B.n595 585
R489 B.n597 B.n596 585
R490 B.n221 B.n220 585
R491 B.n222 B.n221 585
R492 B.n605 B.n604 585
R493 B.n604 B.n603 585
R494 B.n606 B.n219 585
R495 B.n219 B.n217 585
R496 B.n608 B.n607 585
R497 B.n609 B.n608 585
R498 B.n213 B.n212 585
R499 B.n218 B.n213 585
R500 B.n617 B.n616 585
R501 B.n616 B.n615 585
R502 B.n618 B.n211 585
R503 B.n211 B.n210 585
R504 B.n620 B.n619 585
R505 B.n621 B.n620 585
R506 B.n205 B.n204 585
R507 B.n206 B.n205 585
R508 B.n629 B.n628 585
R509 B.n628 B.n627 585
R510 B.n630 B.n203 585
R511 B.n203 B.n202 585
R512 B.n632 B.n631 585
R513 B.n633 B.n632 585
R514 B.n197 B.n196 585
R515 B.n198 B.n197 585
R516 B.n641 B.n640 585
R517 B.n640 B.n639 585
R518 B.n642 B.n195 585
R519 B.n195 B.n194 585
R520 B.n644 B.n643 585
R521 B.n645 B.n644 585
R522 B.n189 B.n188 585
R523 B.n190 B.n189 585
R524 B.n654 B.n653 585
R525 B.n653 B.n652 585
R526 B.n655 B.n187 585
R527 B.n651 B.n187 585
R528 B.n657 B.n656 585
R529 B.n658 B.n657 585
R530 B.n182 B.n181 585
R531 B.n183 B.n182 585
R532 B.n666 B.n665 585
R533 B.n665 B.n664 585
R534 B.n667 B.n180 585
R535 B.n180 B.n179 585
R536 B.n669 B.n668 585
R537 B.n670 B.n669 585
R538 B.n174 B.n173 585
R539 B.n175 B.n174 585
R540 B.n678 B.n677 585
R541 B.n677 B.n676 585
R542 B.n679 B.n172 585
R543 B.n172 B.n171 585
R544 B.n681 B.n680 585
R545 B.n682 B.n681 585
R546 B.n166 B.n165 585
R547 B.n167 B.n166 585
R548 B.n691 B.n690 585
R549 B.n690 B.n689 585
R550 B.n692 B.n164 585
R551 B.n688 B.n164 585
R552 B.n694 B.n693 585
R553 B.n695 B.n694 585
R554 B.n159 B.n158 585
R555 B.n160 B.n159 585
R556 B.n704 B.n703 585
R557 B.n703 B.n702 585
R558 B.n705 B.n157 585
R559 B.n157 B.n156 585
R560 B.n707 B.n706 585
R561 B.n708 B.n707 585
R562 B.n3 B.n0 585
R563 B.n4 B.n3 585
R564 B.n1126 B.n1 585
R565 B.n1127 B.n1126 585
R566 B.n1125 B.n1124 585
R567 B.n1125 B.n8 585
R568 B.n1123 B.n9 585
R569 B.n12 B.n9 585
R570 B.n1122 B.n1121 585
R571 B.n1121 B.n1120 585
R572 B.n11 B.n10 585
R573 B.n1119 B.n11 585
R574 B.n1117 B.n1116 585
R575 B.n1118 B.n1117 585
R576 B.n1115 B.n16 585
R577 B.n19 B.n16 585
R578 B.n1114 B.n1113 585
R579 B.n1113 B.n1112 585
R580 B.n18 B.n17 585
R581 B.n1111 B.n18 585
R582 B.n1109 B.n1108 585
R583 B.n1110 B.n1109 585
R584 B.n1107 B.n24 585
R585 B.n24 B.n23 585
R586 B.n1106 B.n1105 585
R587 B.n1105 B.n1104 585
R588 B.n26 B.n25 585
R589 B.n1103 B.n26 585
R590 B.n1101 B.n1100 585
R591 B.n1102 B.n1101 585
R592 B.n1099 B.n31 585
R593 B.n31 B.n30 585
R594 B.n1098 B.n1097 585
R595 B.n1097 B.n1096 585
R596 B.n33 B.n32 585
R597 B.n1095 B.n33 585
R598 B.n1093 B.n1092 585
R599 B.n1094 B.n1093 585
R600 B.n1091 B.n37 585
R601 B.n40 B.n37 585
R602 B.n1090 B.n1089 585
R603 B.n1089 B.n1088 585
R604 B.n39 B.n38 585
R605 B.n1087 B.n39 585
R606 B.n1085 B.n1084 585
R607 B.n1086 B.n1085 585
R608 B.n1083 B.n45 585
R609 B.n45 B.n44 585
R610 B.n1082 B.n1081 585
R611 B.n1081 B.n1080 585
R612 B.n47 B.n46 585
R613 B.n1079 B.n47 585
R614 B.n1077 B.n1076 585
R615 B.n1078 B.n1077 585
R616 B.n1075 B.n52 585
R617 B.n52 B.n51 585
R618 B.n1074 B.n1073 585
R619 B.n1073 B.n1072 585
R620 B.n54 B.n53 585
R621 B.n1071 B.n54 585
R622 B.n1069 B.n1068 585
R623 B.n1070 B.n1069 585
R624 B.n1067 B.n59 585
R625 B.n59 B.n58 585
R626 B.n1066 B.n1065 585
R627 B.n1065 B.n1064 585
R628 B.n61 B.n60 585
R629 B.n1063 B.n61 585
R630 B.n1061 B.n1060 585
R631 B.n1062 B.n1061 585
R632 B.n1059 B.n66 585
R633 B.n66 B.n65 585
R634 B.n1058 B.n1057 585
R635 B.n1057 B.n1056 585
R636 B.n68 B.n67 585
R637 B.n1055 B.n68 585
R638 B.n1053 B.n1052 585
R639 B.n1054 B.n1053 585
R640 B.n1051 B.n73 585
R641 B.n73 B.n72 585
R642 B.n1050 B.n1049 585
R643 B.n1049 B.n1048 585
R644 B.n75 B.n74 585
R645 B.n1047 B.n75 585
R646 B.n1045 B.n1044 585
R647 B.n1046 B.n1045 585
R648 B.n1130 B.n1129 585
R649 B.n1128 B.n2 585
R650 B.n1045 B.n80 511.721
R651 B.n768 B.n78 511.721
R652 B.n586 B.n233 511.721
R653 B.n584 B.n235 511.721
R654 B.n113 B.t15 342.712
R655 B.n119 B.t11 342.712
R656 B.n276 B.t4 342.712
R657 B.n268 B.t8 342.712
R658 B.n769 B.n79 256.663
R659 B.n771 B.n79 256.663
R660 B.n777 B.n79 256.663
R661 B.n779 B.n79 256.663
R662 B.n785 B.n79 256.663
R663 B.n787 B.n79 256.663
R664 B.n793 B.n79 256.663
R665 B.n795 B.n79 256.663
R666 B.n801 B.n79 256.663
R667 B.n803 B.n79 256.663
R668 B.n809 B.n79 256.663
R669 B.n811 B.n79 256.663
R670 B.n817 B.n79 256.663
R671 B.n819 B.n79 256.663
R672 B.n825 B.n79 256.663
R673 B.n827 B.n79 256.663
R674 B.n833 B.n79 256.663
R675 B.n835 B.n79 256.663
R676 B.n841 B.n79 256.663
R677 B.n843 B.n79 256.663
R678 B.n849 B.n79 256.663
R679 B.n851 B.n79 256.663
R680 B.n857 B.n79 256.663
R681 B.n859 B.n79 256.663
R682 B.n865 B.n79 256.663
R683 B.n867 B.n79 256.663
R684 B.n873 B.n79 256.663
R685 B.n875 B.n79 256.663
R686 B.n881 B.n79 256.663
R687 B.n883 B.n79 256.663
R688 B.n889 B.n79 256.663
R689 B.n122 B.n79 256.663
R690 B.n895 B.n79 256.663
R691 B.n901 B.n79 256.663
R692 B.n903 B.n79 256.663
R693 B.n909 B.n79 256.663
R694 B.n911 B.n79 256.663
R695 B.n918 B.n79 256.663
R696 B.n920 B.n79 256.663
R697 B.n926 B.n79 256.663
R698 B.n928 B.n79 256.663
R699 B.n934 B.n79 256.663
R700 B.n936 B.n79 256.663
R701 B.n942 B.n79 256.663
R702 B.n944 B.n79 256.663
R703 B.n950 B.n79 256.663
R704 B.n952 B.n79 256.663
R705 B.n958 B.n79 256.663
R706 B.n960 B.n79 256.663
R707 B.n966 B.n79 256.663
R708 B.n968 B.n79 256.663
R709 B.n974 B.n79 256.663
R710 B.n976 B.n79 256.663
R711 B.n982 B.n79 256.663
R712 B.n984 B.n79 256.663
R713 B.n990 B.n79 256.663
R714 B.n992 B.n79 256.663
R715 B.n998 B.n79 256.663
R716 B.n1000 B.n79 256.663
R717 B.n1006 B.n79 256.663
R718 B.n1008 B.n79 256.663
R719 B.n1014 B.n79 256.663
R720 B.n1016 B.n79 256.663
R721 B.n1022 B.n79 256.663
R722 B.n1024 B.n79 256.663
R723 B.n1030 B.n79 256.663
R724 B.n1032 B.n79 256.663
R725 B.n1038 B.n79 256.663
R726 B.n1040 B.n79 256.663
R727 B.n579 B.n234 256.663
R728 B.n237 B.n234 256.663
R729 B.n572 B.n234 256.663
R730 B.n566 B.n234 256.663
R731 B.n564 B.n234 256.663
R732 B.n558 B.n234 256.663
R733 B.n556 B.n234 256.663
R734 B.n550 B.n234 256.663
R735 B.n548 B.n234 256.663
R736 B.n542 B.n234 256.663
R737 B.n540 B.n234 256.663
R738 B.n534 B.n234 256.663
R739 B.n532 B.n234 256.663
R740 B.n526 B.n234 256.663
R741 B.n524 B.n234 256.663
R742 B.n518 B.n234 256.663
R743 B.n516 B.n234 256.663
R744 B.n510 B.n234 256.663
R745 B.n508 B.n234 256.663
R746 B.n502 B.n234 256.663
R747 B.n500 B.n234 256.663
R748 B.n494 B.n234 256.663
R749 B.n492 B.n234 256.663
R750 B.n486 B.n234 256.663
R751 B.n484 B.n234 256.663
R752 B.n478 B.n234 256.663
R753 B.n476 B.n234 256.663
R754 B.n470 B.n234 256.663
R755 B.n468 B.n234 256.663
R756 B.n462 B.n234 256.663
R757 B.n460 B.n234 256.663
R758 B.n453 B.n234 256.663
R759 B.n451 B.n234 256.663
R760 B.n445 B.n234 256.663
R761 B.n443 B.n234 256.663
R762 B.n437 B.n234 256.663
R763 B.n435 B.n234 256.663
R764 B.n429 B.n234 256.663
R765 B.n427 B.n234 256.663
R766 B.n421 B.n234 256.663
R767 B.n419 B.n234 256.663
R768 B.n413 B.n234 256.663
R769 B.n411 B.n234 256.663
R770 B.n405 B.n234 256.663
R771 B.n403 B.n234 256.663
R772 B.n397 B.n234 256.663
R773 B.n395 B.n234 256.663
R774 B.n389 B.n234 256.663
R775 B.n387 B.n234 256.663
R776 B.n381 B.n234 256.663
R777 B.n379 B.n234 256.663
R778 B.n373 B.n234 256.663
R779 B.n371 B.n234 256.663
R780 B.n365 B.n234 256.663
R781 B.n363 B.n234 256.663
R782 B.n357 B.n234 256.663
R783 B.n355 B.n234 256.663
R784 B.n349 B.n234 256.663
R785 B.n347 B.n234 256.663
R786 B.n341 B.n234 256.663
R787 B.n339 B.n234 256.663
R788 B.n333 B.n234 256.663
R789 B.n331 B.n234 256.663
R790 B.n325 B.n234 256.663
R791 B.n323 B.n234 256.663
R792 B.n317 B.n234 256.663
R793 B.n315 B.n234 256.663
R794 B.n309 B.n234 256.663
R795 B.n1132 B.n1131 256.663
R796 B.n1041 B.n1039 163.367
R797 B.n1037 B.n82 163.367
R798 B.n1033 B.n1031 163.367
R799 B.n1029 B.n84 163.367
R800 B.n1025 B.n1023 163.367
R801 B.n1021 B.n86 163.367
R802 B.n1017 B.n1015 163.367
R803 B.n1013 B.n88 163.367
R804 B.n1009 B.n1007 163.367
R805 B.n1005 B.n90 163.367
R806 B.n1001 B.n999 163.367
R807 B.n997 B.n92 163.367
R808 B.n993 B.n991 163.367
R809 B.n989 B.n94 163.367
R810 B.n985 B.n983 163.367
R811 B.n981 B.n96 163.367
R812 B.n977 B.n975 163.367
R813 B.n973 B.n98 163.367
R814 B.n969 B.n967 163.367
R815 B.n965 B.n100 163.367
R816 B.n961 B.n959 163.367
R817 B.n957 B.n102 163.367
R818 B.n953 B.n951 163.367
R819 B.n949 B.n104 163.367
R820 B.n945 B.n943 163.367
R821 B.n941 B.n106 163.367
R822 B.n937 B.n935 163.367
R823 B.n933 B.n108 163.367
R824 B.n929 B.n927 163.367
R825 B.n925 B.n110 163.367
R826 B.n921 B.n919 163.367
R827 B.n917 B.n112 163.367
R828 B.n912 B.n910 163.367
R829 B.n908 B.n116 163.367
R830 B.n904 B.n902 163.367
R831 B.n900 B.n118 163.367
R832 B.n896 B.n894 163.367
R833 B.n891 B.n890 163.367
R834 B.n888 B.n124 163.367
R835 B.n884 B.n882 163.367
R836 B.n880 B.n126 163.367
R837 B.n876 B.n874 163.367
R838 B.n872 B.n128 163.367
R839 B.n868 B.n866 163.367
R840 B.n864 B.n130 163.367
R841 B.n860 B.n858 163.367
R842 B.n856 B.n132 163.367
R843 B.n852 B.n850 163.367
R844 B.n848 B.n134 163.367
R845 B.n844 B.n842 163.367
R846 B.n840 B.n136 163.367
R847 B.n836 B.n834 163.367
R848 B.n832 B.n138 163.367
R849 B.n828 B.n826 163.367
R850 B.n824 B.n140 163.367
R851 B.n820 B.n818 163.367
R852 B.n816 B.n142 163.367
R853 B.n812 B.n810 163.367
R854 B.n808 B.n144 163.367
R855 B.n804 B.n802 163.367
R856 B.n800 B.n146 163.367
R857 B.n796 B.n794 163.367
R858 B.n792 B.n148 163.367
R859 B.n788 B.n786 163.367
R860 B.n784 B.n150 163.367
R861 B.n780 B.n778 163.367
R862 B.n776 B.n152 163.367
R863 B.n772 B.n770 163.367
R864 B.n586 B.n231 163.367
R865 B.n590 B.n231 163.367
R866 B.n590 B.n225 163.367
R867 B.n598 B.n225 163.367
R868 B.n598 B.n223 163.367
R869 B.n602 B.n223 163.367
R870 B.n602 B.n216 163.367
R871 B.n610 B.n216 163.367
R872 B.n610 B.n214 163.367
R873 B.n614 B.n214 163.367
R874 B.n614 B.n209 163.367
R875 B.n622 B.n209 163.367
R876 B.n622 B.n207 163.367
R877 B.n626 B.n207 163.367
R878 B.n626 B.n201 163.367
R879 B.n634 B.n201 163.367
R880 B.n634 B.n199 163.367
R881 B.n638 B.n199 163.367
R882 B.n638 B.n193 163.367
R883 B.n646 B.n193 163.367
R884 B.n646 B.n191 163.367
R885 B.n650 B.n191 163.367
R886 B.n650 B.n186 163.367
R887 B.n659 B.n186 163.367
R888 B.n659 B.n184 163.367
R889 B.n663 B.n184 163.367
R890 B.n663 B.n178 163.367
R891 B.n671 B.n178 163.367
R892 B.n671 B.n176 163.367
R893 B.n675 B.n176 163.367
R894 B.n675 B.n170 163.367
R895 B.n683 B.n170 163.367
R896 B.n683 B.n168 163.367
R897 B.n687 B.n168 163.367
R898 B.n687 B.n163 163.367
R899 B.n696 B.n163 163.367
R900 B.n696 B.n161 163.367
R901 B.n701 B.n161 163.367
R902 B.n701 B.n155 163.367
R903 B.n709 B.n155 163.367
R904 B.n710 B.n709 163.367
R905 B.n710 B.n5 163.367
R906 B.n6 B.n5 163.367
R907 B.n7 B.n6 163.367
R908 B.n716 B.n7 163.367
R909 B.n717 B.n716 163.367
R910 B.n717 B.n13 163.367
R911 B.n14 B.n13 163.367
R912 B.n15 B.n14 163.367
R913 B.n722 B.n15 163.367
R914 B.n722 B.n20 163.367
R915 B.n21 B.n20 163.367
R916 B.n22 B.n21 163.367
R917 B.n727 B.n22 163.367
R918 B.n727 B.n27 163.367
R919 B.n28 B.n27 163.367
R920 B.n29 B.n28 163.367
R921 B.n732 B.n29 163.367
R922 B.n732 B.n34 163.367
R923 B.n35 B.n34 163.367
R924 B.n36 B.n35 163.367
R925 B.n737 B.n36 163.367
R926 B.n737 B.n41 163.367
R927 B.n42 B.n41 163.367
R928 B.n43 B.n42 163.367
R929 B.n742 B.n43 163.367
R930 B.n742 B.n48 163.367
R931 B.n49 B.n48 163.367
R932 B.n50 B.n49 163.367
R933 B.n747 B.n50 163.367
R934 B.n747 B.n55 163.367
R935 B.n56 B.n55 163.367
R936 B.n57 B.n56 163.367
R937 B.n752 B.n57 163.367
R938 B.n752 B.n62 163.367
R939 B.n63 B.n62 163.367
R940 B.n64 B.n63 163.367
R941 B.n757 B.n64 163.367
R942 B.n757 B.n69 163.367
R943 B.n70 B.n69 163.367
R944 B.n71 B.n70 163.367
R945 B.n762 B.n71 163.367
R946 B.n762 B.n76 163.367
R947 B.n77 B.n76 163.367
R948 B.n78 B.n77 163.367
R949 B.n580 B.n578 163.367
R950 B.n578 B.n577 163.367
R951 B.n574 B.n573 163.367
R952 B.n571 B.n239 163.367
R953 B.n567 B.n565 163.367
R954 B.n563 B.n241 163.367
R955 B.n559 B.n557 163.367
R956 B.n555 B.n243 163.367
R957 B.n551 B.n549 163.367
R958 B.n547 B.n245 163.367
R959 B.n543 B.n541 163.367
R960 B.n539 B.n247 163.367
R961 B.n535 B.n533 163.367
R962 B.n531 B.n249 163.367
R963 B.n527 B.n525 163.367
R964 B.n523 B.n251 163.367
R965 B.n519 B.n517 163.367
R966 B.n515 B.n253 163.367
R967 B.n511 B.n509 163.367
R968 B.n507 B.n255 163.367
R969 B.n503 B.n501 163.367
R970 B.n499 B.n257 163.367
R971 B.n495 B.n493 163.367
R972 B.n491 B.n259 163.367
R973 B.n487 B.n485 163.367
R974 B.n483 B.n261 163.367
R975 B.n479 B.n477 163.367
R976 B.n475 B.n263 163.367
R977 B.n471 B.n469 163.367
R978 B.n467 B.n265 163.367
R979 B.n463 B.n461 163.367
R980 B.n459 B.n267 163.367
R981 B.n454 B.n452 163.367
R982 B.n450 B.n271 163.367
R983 B.n446 B.n444 163.367
R984 B.n442 B.n273 163.367
R985 B.n438 B.n436 163.367
R986 B.n434 B.n275 163.367
R987 B.n430 B.n428 163.367
R988 B.n426 B.n280 163.367
R989 B.n422 B.n420 163.367
R990 B.n418 B.n282 163.367
R991 B.n414 B.n412 163.367
R992 B.n410 B.n284 163.367
R993 B.n406 B.n404 163.367
R994 B.n402 B.n286 163.367
R995 B.n398 B.n396 163.367
R996 B.n394 B.n288 163.367
R997 B.n390 B.n388 163.367
R998 B.n386 B.n290 163.367
R999 B.n382 B.n380 163.367
R1000 B.n378 B.n292 163.367
R1001 B.n374 B.n372 163.367
R1002 B.n370 B.n294 163.367
R1003 B.n366 B.n364 163.367
R1004 B.n362 B.n296 163.367
R1005 B.n358 B.n356 163.367
R1006 B.n354 B.n298 163.367
R1007 B.n350 B.n348 163.367
R1008 B.n346 B.n300 163.367
R1009 B.n342 B.n340 163.367
R1010 B.n338 B.n302 163.367
R1011 B.n334 B.n332 163.367
R1012 B.n330 B.n304 163.367
R1013 B.n326 B.n324 163.367
R1014 B.n322 B.n306 163.367
R1015 B.n318 B.n316 163.367
R1016 B.n314 B.n308 163.367
R1017 B.n310 B.n233 163.367
R1018 B.n584 B.n229 163.367
R1019 B.n592 B.n229 163.367
R1020 B.n592 B.n227 163.367
R1021 B.n596 B.n227 163.367
R1022 B.n596 B.n221 163.367
R1023 B.n604 B.n221 163.367
R1024 B.n604 B.n219 163.367
R1025 B.n608 B.n219 163.367
R1026 B.n608 B.n213 163.367
R1027 B.n616 B.n213 163.367
R1028 B.n616 B.n211 163.367
R1029 B.n620 B.n211 163.367
R1030 B.n620 B.n205 163.367
R1031 B.n628 B.n205 163.367
R1032 B.n628 B.n203 163.367
R1033 B.n632 B.n203 163.367
R1034 B.n632 B.n197 163.367
R1035 B.n640 B.n197 163.367
R1036 B.n640 B.n195 163.367
R1037 B.n644 B.n195 163.367
R1038 B.n644 B.n189 163.367
R1039 B.n653 B.n189 163.367
R1040 B.n653 B.n187 163.367
R1041 B.n657 B.n187 163.367
R1042 B.n657 B.n182 163.367
R1043 B.n665 B.n182 163.367
R1044 B.n665 B.n180 163.367
R1045 B.n669 B.n180 163.367
R1046 B.n669 B.n174 163.367
R1047 B.n677 B.n174 163.367
R1048 B.n677 B.n172 163.367
R1049 B.n681 B.n172 163.367
R1050 B.n681 B.n166 163.367
R1051 B.n690 B.n166 163.367
R1052 B.n690 B.n164 163.367
R1053 B.n694 B.n164 163.367
R1054 B.n694 B.n159 163.367
R1055 B.n703 B.n159 163.367
R1056 B.n703 B.n157 163.367
R1057 B.n707 B.n157 163.367
R1058 B.n707 B.n3 163.367
R1059 B.n1130 B.n3 163.367
R1060 B.n1126 B.n2 163.367
R1061 B.n1126 B.n1125 163.367
R1062 B.n1125 B.n9 163.367
R1063 B.n1121 B.n9 163.367
R1064 B.n1121 B.n11 163.367
R1065 B.n1117 B.n11 163.367
R1066 B.n1117 B.n16 163.367
R1067 B.n1113 B.n16 163.367
R1068 B.n1113 B.n18 163.367
R1069 B.n1109 B.n18 163.367
R1070 B.n1109 B.n24 163.367
R1071 B.n1105 B.n24 163.367
R1072 B.n1105 B.n26 163.367
R1073 B.n1101 B.n26 163.367
R1074 B.n1101 B.n31 163.367
R1075 B.n1097 B.n31 163.367
R1076 B.n1097 B.n33 163.367
R1077 B.n1093 B.n33 163.367
R1078 B.n1093 B.n37 163.367
R1079 B.n1089 B.n37 163.367
R1080 B.n1089 B.n39 163.367
R1081 B.n1085 B.n39 163.367
R1082 B.n1085 B.n45 163.367
R1083 B.n1081 B.n45 163.367
R1084 B.n1081 B.n47 163.367
R1085 B.n1077 B.n47 163.367
R1086 B.n1077 B.n52 163.367
R1087 B.n1073 B.n52 163.367
R1088 B.n1073 B.n54 163.367
R1089 B.n1069 B.n54 163.367
R1090 B.n1069 B.n59 163.367
R1091 B.n1065 B.n59 163.367
R1092 B.n1065 B.n61 163.367
R1093 B.n1061 B.n61 163.367
R1094 B.n1061 B.n66 163.367
R1095 B.n1057 B.n66 163.367
R1096 B.n1057 B.n68 163.367
R1097 B.n1053 B.n68 163.367
R1098 B.n1053 B.n73 163.367
R1099 B.n1049 B.n73 163.367
R1100 B.n1049 B.n75 163.367
R1101 B.n1045 B.n75 163.367
R1102 B.n119 B.t13 142.792
R1103 B.n276 B.t7 142.792
R1104 B.n113 B.t16 142.764
R1105 B.n268 B.t10 142.764
R1106 B.n114 B.n113 75.4429
R1107 B.n120 B.n119 75.4429
R1108 B.n277 B.n276 75.4429
R1109 B.n269 B.n268 75.4429
R1110 B.n1040 B.n80 71.676
R1111 B.n1039 B.n1038 71.676
R1112 B.n1032 B.n82 71.676
R1113 B.n1031 B.n1030 71.676
R1114 B.n1024 B.n84 71.676
R1115 B.n1023 B.n1022 71.676
R1116 B.n1016 B.n86 71.676
R1117 B.n1015 B.n1014 71.676
R1118 B.n1008 B.n88 71.676
R1119 B.n1007 B.n1006 71.676
R1120 B.n1000 B.n90 71.676
R1121 B.n999 B.n998 71.676
R1122 B.n992 B.n92 71.676
R1123 B.n991 B.n990 71.676
R1124 B.n984 B.n94 71.676
R1125 B.n983 B.n982 71.676
R1126 B.n976 B.n96 71.676
R1127 B.n975 B.n974 71.676
R1128 B.n968 B.n98 71.676
R1129 B.n967 B.n966 71.676
R1130 B.n960 B.n100 71.676
R1131 B.n959 B.n958 71.676
R1132 B.n952 B.n102 71.676
R1133 B.n951 B.n950 71.676
R1134 B.n944 B.n104 71.676
R1135 B.n943 B.n942 71.676
R1136 B.n936 B.n106 71.676
R1137 B.n935 B.n934 71.676
R1138 B.n928 B.n108 71.676
R1139 B.n927 B.n926 71.676
R1140 B.n920 B.n110 71.676
R1141 B.n919 B.n918 71.676
R1142 B.n911 B.n112 71.676
R1143 B.n910 B.n909 71.676
R1144 B.n903 B.n116 71.676
R1145 B.n902 B.n901 71.676
R1146 B.n895 B.n118 71.676
R1147 B.n894 B.n122 71.676
R1148 B.n890 B.n889 71.676
R1149 B.n883 B.n124 71.676
R1150 B.n882 B.n881 71.676
R1151 B.n875 B.n126 71.676
R1152 B.n874 B.n873 71.676
R1153 B.n867 B.n128 71.676
R1154 B.n866 B.n865 71.676
R1155 B.n859 B.n130 71.676
R1156 B.n858 B.n857 71.676
R1157 B.n851 B.n132 71.676
R1158 B.n850 B.n849 71.676
R1159 B.n843 B.n134 71.676
R1160 B.n842 B.n841 71.676
R1161 B.n835 B.n136 71.676
R1162 B.n834 B.n833 71.676
R1163 B.n827 B.n138 71.676
R1164 B.n826 B.n825 71.676
R1165 B.n819 B.n140 71.676
R1166 B.n818 B.n817 71.676
R1167 B.n811 B.n142 71.676
R1168 B.n810 B.n809 71.676
R1169 B.n803 B.n144 71.676
R1170 B.n802 B.n801 71.676
R1171 B.n795 B.n146 71.676
R1172 B.n794 B.n793 71.676
R1173 B.n787 B.n148 71.676
R1174 B.n786 B.n785 71.676
R1175 B.n779 B.n150 71.676
R1176 B.n778 B.n777 71.676
R1177 B.n771 B.n152 71.676
R1178 B.n770 B.n769 71.676
R1179 B.n769 B.n768 71.676
R1180 B.n772 B.n771 71.676
R1181 B.n777 B.n776 71.676
R1182 B.n780 B.n779 71.676
R1183 B.n785 B.n784 71.676
R1184 B.n788 B.n787 71.676
R1185 B.n793 B.n792 71.676
R1186 B.n796 B.n795 71.676
R1187 B.n801 B.n800 71.676
R1188 B.n804 B.n803 71.676
R1189 B.n809 B.n808 71.676
R1190 B.n812 B.n811 71.676
R1191 B.n817 B.n816 71.676
R1192 B.n820 B.n819 71.676
R1193 B.n825 B.n824 71.676
R1194 B.n828 B.n827 71.676
R1195 B.n833 B.n832 71.676
R1196 B.n836 B.n835 71.676
R1197 B.n841 B.n840 71.676
R1198 B.n844 B.n843 71.676
R1199 B.n849 B.n848 71.676
R1200 B.n852 B.n851 71.676
R1201 B.n857 B.n856 71.676
R1202 B.n860 B.n859 71.676
R1203 B.n865 B.n864 71.676
R1204 B.n868 B.n867 71.676
R1205 B.n873 B.n872 71.676
R1206 B.n876 B.n875 71.676
R1207 B.n881 B.n880 71.676
R1208 B.n884 B.n883 71.676
R1209 B.n889 B.n888 71.676
R1210 B.n891 B.n122 71.676
R1211 B.n896 B.n895 71.676
R1212 B.n901 B.n900 71.676
R1213 B.n904 B.n903 71.676
R1214 B.n909 B.n908 71.676
R1215 B.n912 B.n911 71.676
R1216 B.n918 B.n917 71.676
R1217 B.n921 B.n920 71.676
R1218 B.n926 B.n925 71.676
R1219 B.n929 B.n928 71.676
R1220 B.n934 B.n933 71.676
R1221 B.n937 B.n936 71.676
R1222 B.n942 B.n941 71.676
R1223 B.n945 B.n944 71.676
R1224 B.n950 B.n949 71.676
R1225 B.n953 B.n952 71.676
R1226 B.n958 B.n957 71.676
R1227 B.n961 B.n960 71.676
R1228 B.n966 B.n965 71.676
R1229 B.n969 B.n968 71.676
R1230 B.n974 B.n973 71.676
R1231 B.n977 B.n976 71.676
R1232 B.n982 B.n981 71.676
R1233 B.n985 B.n984 71.676
R1234 B.n990 B.n989 71.676
R1235 B.n993 B.n992 71.676
R1236 B.n998 B.n997 71.676
R1237 B.n1001 B.n1000 71.676
R1238 B.n1006 B.n1005 71.676
R1239 B.n1009 B.n1008 71.676
R1240 B.n1014 B.n1013 71.676
R1241 B.n1017 B.n1016 71.676
R1242 B.n1022 B.n1021 71.676
R1243 B.n1025 B.n1024 71.676
R1244 B.n1030 B.n1029 71.676
R1245 B.n1033 B.n1032 71.676
R1246 B.n1038 B.n1037 71.676
R1247 B.n1041 B.n1040 71.676
R1248 B.n579 B.n235 71.676
R1249 B.n577 B.n237 71.676
R1250 B.n573 B.n572 71.676
R1251 B.n566 B.n239 71.676
R1252 B.n565 B.n564 71.676
R1253 B.n558 B.n241 71.676
R1254 B.n557 B.n556 71.676
R1255 B.n550 B.n243 71.676
R1256 B.n549 B.n548 71.676
R1257 B.n542 B.n245 71.676
R1258 B.n541 B.n540 71.676
R1259 B.n534 B.n247 71.676
R1260 B.n533 B.n532 71.676
R1261 B.n526 B.n249 71.676
R1262 B.n525 B.n524 71.676
R1263 B.n518 B.n251 71.676
R1264 B.n517 B.n516 71.676
R1265 B.n510 B.n253 71.676
R1266 B.n509 B.n508 71.676
R1267 B.n502 B.n255 71.676
R1268 B.n501 B.n500 71.676
R1269 B.n494 B.n257 71.676
R1270 B.n493 B.n492 71.676
R1271 B.n486 B.n259 71.676
R1272 B.n485 B.n484 71.676
R1273 B.n478 B.n261 71.676
R1274 B.n477 B.n476 71.676
R1275 B.n470 B.n263 71.676
R1276 B.n469 B.n468 71.676
R1277 B.n462 B.n265 71.676
R1278 B.n461 B.n460 71.676
R1279 B.n453 B.n267 71.676
R1280 B.n452 B.n451 71.676
R1281 B.n445 B.n271 71.676
R1282 B.n444 B.n443 71.676
R1283 B.n437 B.n273 71.676
R1284 B.n436 B.n435 71.676
R1285 B.n429 B.n275 71.676
R1286 B.n428 B.n427 71.676
R1287 B.n421 B.n280 71.676
R1288 B.n420 B.n419 71.676
R1289 B.n413 B.n282 71.676
R1290 B.n412 B.n411 71.676
R1291 B.n405 B.n284 71.676
R1292 B.n404 B.n403 71.676
R1293 B.n397 B.n286 71.676
R1294 B.n396 B.n395 71.676
R1295 B.n389 B.n288 71.676
R1296 B.n388 B.n387 71.676
R1297 B.n381 B.n290 71.676
R1298 B.n380 B.n379 71.676
R1299 B.n373 B.n292 71.676
R1300 B.n372 B.n371 71.676
R1301 B.n365 B.n294 71.676
R1302 B.n364 B.n363 71.676
R1303 B.n357 B.n296 71.676
R1304 B.n356 B.n355 71.676
R1305 B.n349 B.n298 71.676
R1306 B.n348 B.n347 71.676
R1307 B.n341 B.n300 71.676
R1308 B.n340 B.n339 71.676
R1309 B.n333 B.n302 71.676
R1310 B.n332 B.n331 71.676
R1311 B.n325 B.n304 71.676
R1312 B.n324 B.n323 71.676
R1313 B.n317 B.n306 71.676
R1314 B.n316 B.n315 71.676
R1315 B.n309 B.n308 71.676
R1316 B.n580 B.n579 71.676
R1317 B.n574 B.n237 71.676
R1318 B.n572 B.n571 71.676
R1319 B.n567 B.n566 71.676
R1320 B.n564 B.n563 71.676
R1321 B.n559 B.n558 71.676
R1322 B.n556 B.n555 71.676
R1323 B.n551 B.n550 71.676
R1324 B.n548 B.n547 71.676
R1325 B.n543 B.n542 71.676
R1326 B.n540 B.n539 71.676
R1327 B.n535 B.n534 71.676
R1328 B.n532 B.n531 71.676
R1329 B.n527 B.n526 71.676
R1330 B.n524 B.n523 71.676
R1331 B.n519 B.n518 71.676
R1332 B.n516 B.n515 71.676
R1333 B.n511 B.n510 71.676
R1334 B.n508 B.n507 71.676
R1335 B.n503 B.n502 71.676
R1336 B.n500 B.n499 71.676
R1337 B.n495 B.n494 71.676
R1338 B.n492 B.n491 71.676
R1339 B.n487 B.n486 71.676
R1340 B.n484 B.n483 71.676
R1341 B.n479 B.n478 71.676
R1342 B.n476 B.n475 71.676
R1343 B.n471 B.n470 71.676
R1344 B.n468 B.n467 71.676
R1345 B.n463 B.n462 71.676
R1346 B.n460 B.n459 71.676
R1347 B.n454 B.n453 71.676
R1348 B.n451 B.n450 71.676
R1349 B.n446 B.n445 71.676
R1350 B.n443 B.n442 71.676
R1351 B.n438 B.n437 71.676
R1352 B.n435 B.n434 71.676
R1353 B.n430 B.n429 71.676
R1354 B.n427 B.n426 71.676
R1355 B.n422 B.n421 71.676
R1356 B.n419 B.n418 71.676
R1357 B.n414 B.n413 71.676
R1358 B.n411 B.n410 71.676
R1359 B.n406 B.n405 71.676
R1360 B.n403 B.n402 71.676
R1361 B.n398 B.n397 71.676
R1362 B.n395 B.n394 71.676
R1363 B.n390 B.n389 71.676
R1364 B.n387 B.n386 71.676
R1365 B.n382 B.n381 71.676
R1366 B.n379 B.n378 71.676
R1367 B.n374 B.n373 71.676
R1368 B.n371 B.n370 71.676
R1369 B.n366 B.n365 71.676
R1370 B.n363 B.n362 71.676
R1371 B.n358 B.n357 71.676
R1372 B.n355 B.n354 71.676
R1373 B.n350 B.n349 71.676
R1374 B.n347 B.n346 71.676
R1375 B.n342 B.n341 71.676
R1376 B.n339 B.n338 71.676
R1377 B.n334 B.n333 71.676
R1378 B.n331 B.n330 71.676
R1379 B.n326 B.n325 71.676
R1380 B.n323 B.n322 71.676
R1381 B.n318 B.n317 71.676
R1382 B.n315 B.n314 71.676
R1383 B.n310 B.n309 71.676
R1384 B.n1131 B.n1130 71.676
R1385 B.n1131 B.n2 71.676
R1386 B.n120 B.t14 67.3489
R1387 B.n277 B.t6 67.3489
R1388 B.n114 B.t17 67.3221
R1389 B.n269 B.t9 67.3221
R1390 B.n915 B.n114 59.5399
R1391 B.n121 B.n120 59.5399
R1392 B.n278 B.n277 59.5399
R1393 B.n456 B.n269 59.5399
R1394 B.n585 B.n234 52.35
R1395 B.n1046 B.n79 52.35
R1396 B.n583 B.n582 33.2493
R1397 B.n587 B.n232 33.2493
R1398 B.n767 B.n766 33.2493
R1399 B.n1044 B.n1043 33.2493
R1400 B.n585 B.n230 29.9145
R1401 B.n591 B.n230 29.9145
R1402 B.n591 B.n226 29.9145
R1403 B.n597 B.n226 29.9145
R1404 B.n597 B.n222 29.9145
R1405 B.n603 B.n222 29.9145
R1406 B.n603 B.n217 29.9145
R1407 B.n609 B.n217 29.9145
R1408 B.n609 B.n218 29.9145
R1409 B.n615 B.n210 29.9145
R1410 B.n621 B.n210 29.9145
R1411 B.n621 B.n206 29.9145
R1412 B.n627 B.n206 29.9145
R1413 B.n627 B.n202 29.9145
R1414 B.n633 B.n202 29.9145
R1415 B.n633 B.n198 29.9145
R1416 B.n639 B.n198 29.9145
R1417 B.n639 B.n194 29.9145
R1418 B.n645 B.n194 29.9145
R1419 B.n645 B.n190 29.9145
R1420 B.n652 B.n190 29.9145
R1421 B.n652 B.n651 29.9145
R1422 B.n658 B.n183 29.9145
R1423 B.n664 B.n183 29.9145
R1424 B.n664 B.n179 29.9145
R1425 B.n670 B.n179 29.9145
R1426 B.n670 B.n175 29.9145
R1427 B.n676 B.n175 29.9145
R1428 B.n676 B.n171 29.9145
R1429 B.n682 B.n171 29.9145
R1430 B.n682 B.n167 29.9145
R1431 B.n689 B.n167 29.9145
R1432 B.n689 B.n688 29.9145
R1433 B.n695 B.n160 29.9145
R1434 B.n702 B.n160 29.9145
R1435 B.n702 B.n156 29.9145
R1436 B.n708 B.n156 29.9145
R1437 B.n708 B.n4 29.9145
R1438 B.n1129 B.n4 29.9145
R1439 B.n1129 B.n1128 29.9145
R1440 B.n1128 B.n1127 29.9145
R1441 B.n1127 B.n8 29.9145
R1442 B.n12 B.n8 29.9145
R1443 B.n1120 B.n12 29.9145
R1444 B.n1120 B.n1119 29.9145
R1445 B.n1119 B.n1118 29.9145
R1446 B.n1112 B.n19 29.9145
R1447 B.n1112 B.n1111 29.9145
R1448 B.n1111 B.n1110 29.9145
R1449 B.n1110 B.n23 29.9145
R1450 B.n1104 B.n23 29.9145
R1451 B.n1104 B.n1103 29.9145
R1452 B.n1103 B.n1102 29.9145
R1453 B.n1102 B.n30 29.9145
R1454 B.n1096 B.n30 29.9145
R1455 B.n1096 B.n1095 29.9145
R1456 B.n1095 B.n1094 29.9145
R1457 B.n1088 B.n40 29.9145
R1458 B.n1088 B.n1087 29.9145
R1459 B.n1087 B.n1086 29.9145
R1460 B.n1086 B.n44 29.9145
R1461 B.n1080 B.n44 29.9145
R1462 B.n1080 B.n1079 29.9145
R1463 B.n1079 B.n1078 29.9145
R1464 B.n1078 B.n51 29.9145
R1465 B.n1072 B.n51 29.9145
R1466 B.n1072 B.n1071 29.9145
R1467 B.n1071 B.n1070 29.9145
R1468 B.n1070 B.n58 29.9145
R1469 B.n1064 B.n58 29.9145
R1470 B.n1063 B.n1062 29.9145
R1471 B.n1062 B.n65 29.9145
R1472 B.n1056 B.n65 29.9145
R1473 B.n1056 B.n1055 29.9145
R1474 B.n1055 B.n1054 29.9145
R1475 B.n1054 B.n72 29.9145
R1476 B.n1048 B.n72 29.9145
R1477 B.n1048 B.n1047 29.9145
R1478 B.n1047 B.n1046 29.9145
R1479 B.n615 B.t5 27.275
R1480 B.n1064 B.t12 27.275
R1481 B.n695 B.t2 24.6356
R1482 B.n1118 B.t3 24.6356
R1483 B.n651 B.t0 21.9961
R1484 B.n40 B.t1 21.9961
R1485 B B.n1132 18.0485
R1486 B.n583 B.n228 10.6151
R1487 B.n593 B.n228 10.6151
R1488 B.n594 B.n593 10.6151
R1489 B.n595 B.n594 10.6151
R1490 B.n595 B.n220 10.6151
R1491 B.n605 B.n220 10.6151
R1492 B.n606 B.n605 10.6151
R1493 B.n607 B.n606 10.6151
R1494 B.n607 B.n212 10.6151
R1495 B.n617 B.n212 10.6151
R1496 B.n618 B.n617 10.6151
R1497 B.n619 B.n618 10.6151
R1498 B.n619 B.n204 10.6151
R1499 B.n629 B.n204 10.6151
R1500 B.n630 B.n629 10.6151
R1501 B.n631 B.n630 10.6151
R1502 B.n631 B.n196 10.6151
R1503 B.n641 B.n196 10.6151
R1504 B.n642 B.n641 10.6151
R1505 B.n643 B.n642 10.6151
R1506 B.n643 B.n188 10.6151
R1507 B.n654 B.n188 10.6151
R1508 B.n655 B.n654 10.6151
R1509 B.n656 B.n655 10.6151
R1510 B.n656 B.n181 10.6151
R1511 B.n666 B.n181 10.6151
R1512 B.n667 B.n666 10.6151
R1513 B.n668 B.n667 10.6151
R1514 B.n668 B.n173 10.6151
R1515 B.n678 B.n173 10.6151
R1516 B.n679 B.n678 10.6151
R1517 B.n680 B.n679 10.6151
R1518 B.n680 B.n165 10.6151
R1519 B.n691 B.n165 10.6151
R1520 B.n692 B.n691 10.6151
R1521 B.n693 B.n692 10.6151
R1522 B.n693 B.n158 10.6151
R1523 B.n704 B.n158 10.6151
R1524 B.n705 B.n704 10.6151
R1525 B.n706 B.n705 10.6151
R1526 B.n706 B.n0 10.6151
R1527 B.n582 B.n581 10.6151
R1528 B.n581 B.n236 10.6151
R1529 B.n576 B.n236 10.6151
R1530 B.n576 B.n575 10.6151
R1531 B.n575 B.n238 10.6151
R1532 B.n570 B.n238 10.6151
R1533 B.n570 B.n569 10.6151
R1534 B.n569 B.n568 10.6151
R1535 B.n568 B.n240 10.6151
R1536 B.n562 B.n240 10.6151
R1537 B.n562 B.n561 10.6151
R1538 B.n561 B.n560 10.6151
R1539 B.n560 B.n242 10.6151
R1540 B.n554 B.n242 10.6151
R1541 B.n554 B.n553 10.6151
R1542 B.n553 B.n552 10.6151
R1543 B.n552 B.n244 10.6151
R1544 B.n546 B.n244 10.6151
R1545 B.n546 B.n545 10.6151
R1546 B.n545 B.n544 10.6151
R1547 B.n544 B.n246 10.6151
R1548 B.n538 B.n246 10.6151
R1549 B.n538 B.n537 10.6151
R1550 B.n537 B.n536 10.6151
R1551 B.n536 B.n248 10.6151
R1552 B.n530 B.n248 10.6151
R1553 B.n530 B.n529 10.6151
R1554 B.n529 B.n528 10.6151
R1555 B.n528 B.n250 10.6151
R1556 B.n522 B.n250 10.6151
R1557 B.n522 B.n521 10.6151
R1558 B.n521 B.n520 10.6151
R1559 B.n520 B.n252 10.6151
R1560 B.n514 B.n252 10.6151
R1561 B.n514 B.n513 10.6151
R1562 B.n513 B.n512 10.6151
R1563 B.n512 B.n254 10.6151
R1564 B.n506 B.n254 10.6151
R1565 B.n506 B.n505 10.6151
R1566 B.n505 B.n504 10.6151
R1567 B.n504 B.n256 10.6151
R1568 B.n498 B.n256 10.6151
R1569 B.n498 B.n497 10.6151
R1570 B.n497 B.n496 10.6151
R1571 B.n496 B.n258 10.6151
R1572 B.n490 B.n258 10.6151
R1573 B.n490 B.n489 10.6151
R1574 B.n489 B.n488 10.6151
R1575 B.n488 B.n260 10.6151
R1576 B.n482 B.n260 10.6151
R1577 B.n482 B.n481 10.6151
R1578 B.n481 B.n480 10.6151
R1579 B.n480 B.n262 10.6151
R1580 B.n474 B.n262 10.6151
R1581 B.n474 B.n473 10.6151
R1582 B.n473 B.n472 10.6151
R1583 B.n472 B.n264 10.6151
R1584 B.n466 B.n264 10.6151
R1585 B.n466 B.n465 10.6151
R1586 B.n465 B.n464 10.6151
R1587 B.n464 B.n266 10.6151
R1588 B.n458 B.n266 10.6151
R1589 B.n458 B.n457 10.6151
R1590 B.n455 B.n270 10.6151
R1591 B.n449 B.n270 10.6151
R1592 B.n449 B.n448 10.6151
R1593 B.n448 B.n447 10.6151
R1594 B.n447 B.n272 10.6151
R1595 B.n441 B.n272 10.6151
R1596 B.n441 B.n440 10.6151
R1597 B.n440 B.n439 10.6151
R1598 B.n439 B.n274 10.6151
R1599 B.n433 B.n432 10.6151
R1600 B.n432 B.n431 10.6151
R1601 B.n431 B.n279 10.6151
R1602 B.n425 B.n279 10.6151
R1603 B.n425 B.n424 10.6151
R1604 B.n424 B.n423 10.6151
R1605 B.n423 B.n281 10.6151
R1606 B.n417 B.n281 10.6151
R1607 B.n417 B.n416 10.6151
R1608 B.n416 B.n415 10.6151
R1609 B.n415 B.n283 10.6151
R1610 B.n409 B.n283 10.6151
R1611 B.n409 B.n408 10.6151
R1612 B.n408 B.n407 10.6151
R1613 B.n407 B.n285 10.6151
R1614 B.n401 B.n285 10.6151
R1615 B.n401 B.n400 10.6151
R1616 B.n400 B.n399 10.6151
R1617 B.n399 B.n287 10.6151
R1618 B.n393 B.n287 10.6151
R1619 B.n393 B.n392 10.6151
R1620 B.n392 B.n391 10.6151
R1621 B.n391 B.n289 10.6151
R1622 B.n385 B.n289 10.6151
R1623 B.n385 B.n384 10.6151
R1624 B.n384 B.n383 10.6151
R1625 B.n383 B.n291 10.6151
R1626 B.n377 B.n291 10.6151
R1627 B.n377 B.n376 10.6151
R1628 B.n376 B.n375 10.6151
R1629 B.n375 B.n293 10.6151
R1630 B.n369 B.n293 10.6151
R1631 B.n369 B.n368 10.6151
R1632 B.n368 B.n367 10.6151
R1633 B.n367 B.n295 10.6151
R1634 B.n361 B.n295 10.6151
R1635 B.n361 B.n360 10.6151
R1636 B.n360 B.n359 10.6151
R1637 B.n359 B.n297 10.6151
R1638 B.n353 B.n297 10.6151
R1639 B.n353 B.n352 10.6151
R1640 B.n352 B.n351 10.6151
R1641 B.n351 B.n299 10.6151
R1642 B.n345 B.n299 10.6151
R1643 B.n345 B.n344 10.6151
R1644 B.n344 B.n343 10.6151
R1645 B.n343 B.n301 10.6151
R1646 B.n337 B.n301 10.6151
R1647 B.n337 B.n336 10.6151
R1648 B.n336 B.n335 10.6151
R1649 B.n335 B.n303 10.6151
R1650 B.n329 B.n303 10.6151
R1651 B.n329 B.n328 10.6151
R1652 B.n328 B.n327 10.6151
R1653 B.n327 B.n305 10.6151
R1654 B.n321 B.n305 10.6151
R1655 B.n321 B.n320 10.6151
R1656 B.n320 B.n319 10.6151
R1657 B.n319 B.n307 10.6151
R1658 B.n313 B.n307 10.6151
R1659 B.n313 B.n312 10.6151
R1660 B.n312 B.n311 10.6151
R1661 B.n311 B.n232 10.6151
R1662 B.n588 B.n587 10.6151
R1663 B.n589 B.n588 10.6151
R1664 B.n589 B.n224 10.6151
R1665 B.n599 B.n224 10.6151
R1666 B.n600 B.n599 10.6151
R1667 B.n601 B.n600 10.6151
R1668 B.n601 B.n215 10.6151
R1669 B.n611 B.n215 10.6151
R1670 B.n612 B.n611 10.6151
R1671 B.n613 B.n612 10.6151
R1672 B.n613 B.n208 10.6151
R1673 B.n623 B.n208 10.6151
R1674 B.n624 B.n623 10.6151
R1675 B.n625 B.n624 10.6151
R1676 B.n625 B.n200 10.6151
R1677 B.n635 B.n200 10.6151
R1678 B.n636 B.n635 10.6151
R1679 B.n637 B.n636 10.6151
R1680 B.n637 B.n192 10.6151
R1681 B.n647 B.n192 10.6151
R1682 B.n648 B.n647 10.6151
R1683 B.n649 B.n648 10.6151
R1684 B.n649 B.n185 10.6151
R1685 B.n660 B.n185 10.6151
R1686 B.n661 B.n660 10.6151
R1687 B.n662 B.n661 10.6151
R1688 B.n662 B.n177 10.6151
R1689 B.n672 B.n177 10.6151
R1690 B.n673 B.n672 10.6151
R1691 B.n674 B.n673 10.6151
R1692 B.n674 B.n169 10.6151
R1693 B.n684 B.n169 10.6151
R1694 B.n685 B.n684 10.6151
R1695 B.n686 B.n685 10.6151
R1696 B.n686 B.n162 10.6151
R1697 B.n697 B.n162 10.6151
R1698 B.n698 B.n697 10.6151
R1699 B.n700 B.n698 10.6151
R1700 B.n700 B.n699 10.6151
R1701 B.n699 B.n154 10.6151
R1702 B.n711 B.n154 10.6151
R1703 B.n712 B.n711 10.6151
R1704 B.n713 B.n712 10.6151
R1705 B.n714 B.n713 10.6151
R1706 B.n715 B.n714 10.6151
R1707 B.n718 B.n715 10.6151
R1708 B.n719 B.n718 10.6151
R1709 B.n720 B.n719 10.6151
R1710 B.n721 B.n720 10.6151
R1711 B.n723 B.n721 10.6151
R1712 B.n724 B.n723 10.6151
R1713 B.n725 B.n724 10.6151
R1714 B.n726 B.n725 10.6151
R1715 B.n728 B.n726 10.6151
R1716 B.n729 B.n728 10.6151
R1717 B.n730 B.n729 10.6151
R1718 B.n731 B.n730 10.6151
R1719 B.n733 B.n731 10.6151
R1720 B.n734 B.n733 10.6151
R1721 B.n735 B.n734 10.6151
R1722 B.n736 B.n735 10.6151
R1723 B.n738 B.n736 10.6151
R1724 B.n739 B.n738 10.6151
R1725 B.n740 B.n739 10.6151
R1726 B.n741 B.n740 10.6151
R1727 B.n743 B.n741 10.6151
R1728 B.n744 B.n743 10.6151
R1729 B.n745 B.n744 10.6151
R1730 B.n746 B.n745 10.6151
R1731 B.n748 B.n746 10.6151
R1732 B.n749 B.n748 10.6151
R1733 B.n750 B.n749 10.6151
R1734 B.n751 B.n750 10.6151
R1735 B.n753 B.n751 10.6151
R1736 B.n754 B.n753 10.6151
R1737 B.n755 B.n754 10.6151
R1738 B.n756 B.n755 10.6151
R1739 B.n758 B.n756 10.6151
R1740 B.n759 B.n758 10.6151
R1741 B.n760 B.n759 10.6151
R1742 B.n761 B.n760 10.6151
R1743 B.n763 B.n761 10.6151
R1744 B.n764 B.n763 10.6151
R1745 B.n765 B.n764 10.6151
R1746 B.n766 B.n765 10.6151
R1747 B.n1124 B.n1 10.6151
R1748 B.n1124 B.n1123 10.6151
R1749 B.n1123 B.n1122 10.6151
R1750 B.n1122 B.n10 10.6151
R1751 B.n1116 B.n10 10.6151
R1752 B.n1116 B.n1115 10.6151
R1753 B.n1115 B.n1114 10.6151
R1754 B.n1114 B.n17 10.6151
R1755 B.n1108 B.n17 10.6151
R1756 B.n1108 B.n1107 10.6151
R1757 B.n1107 B.n1106 10.6151
R1758 B.n1106 B.n25 10.6151
R1759 B.n1100 B.n25 10.6151
R1760 B.n1100 B.n1099 10.6151
R1761 B.n1099 B.n1098 10.6151
R1762 B.n1098 B.n32 10.6151
R1763 B.n1092 B.n32 10.6151
R1764 B.n1092 B.n1091 10.6151
R1765 B.n1091 B.n1090 10.6151
R1766 B.n1090 B.n38 10.6151
R1767 B.n1084 B.n38 10.6151
R1768 B.n1084 B.n1083 10.6151
R1769 B.n1083 B.n1082 10.6151
R1770 B.n1082 B.n46 10.6151
R1771 B.n1076 B.n46 10.6151
R1772 B.n1076 B.n1075 10.6151
R1773 B.n1075 B.n1074 10.6151
R1774 B.n1074 B.n53 10.6151
R1775 B.n1068 B.n53 10.6151
R1776 B.n1068 B.n1067 10.6151
R1777 B.n1067 B.n1066 10.6151
R1778 B.n1066 B.n60 10.6151
R1779 B.n1060 B.n60 10.6151
R1780 B.n1060 B.n1059 10.6151
R1781 B.n1059 B.n1058 10.6151
R1782 B.n1058 B.n67 10.6151
R1783 B.n1052 B.n67 10.6151
R1784 B.n1052 B.n1051 10.6151
R1785 B.n1051 B.n1050 10.6151
R1786 B.n1050 B.n74 10.6151
R1787 B.n1044 B.n74 10.6151
R1788 B.n1043 B.n1042 10.6151
R1789 B.n1042 B.n81 10.6151
R1790 B.n1036 B.n81 10.6151
R1791 B.n1036 B.n1035 10.6151
R1792 B.n1035 B.n1034 10.6151
R1793 B.n1034 B.n83 10.6151
R1794 B.n1028 B.n83 10.6151
R1795 B.n1028 B.n1027 10.6151
R1796 B.n1027 B.n1026 10.6151
R1797 B.n1026 B.n85 10.6151
R1798 B.n1020 B.n85 10.6151
R1799 B.n1020 B.n1019 10.6151
R1800 B.n1019 B.n1018 10.6151
R1801 B.n1018 B.n87 10.6151
R1802 B.n1012 B.n87 10.6151
R1803 B.n1012 B.n1011 10.6151
R1804 B.n1011 B.n1010 10.6151
R1805 B.n1010 B.n89 10.6151
R1806 B.n1004 B.n89 10.6151
R1807 B.n1004 B.n1003 10.6151
R1808 B.n1003 B.n1002 10.6151
R1809 B.n1002 B.n91 10.6151
R1810 B.n996 B.n91 10.6151
R1811 B.n996 B.n995 10.6151
R1812 B.n995 B.n994 10.6151
R1813 B.n994 B.n93 10.6151
R1814 B.n988 B.n93 10.6151
R1815 B.n988 B.n987 10.6151
R1816 B.n987 B.n986 10.6151
R1817 B.n986 B.n95 10.6151
R1818 B.n980 B.n95 10.6151
R1819 B.n980 B.n979 10.6151
R1820 B.n979 B.n978 10.6151
R1821 B.n978 B.n97 10.6151
R1822 B.n972 B.n97 10.6151
R1823 B.n972 B.n971 10.6151
R1824 B.n971 B.n970 10.6151
R1825 B.n970 B.n99 10.6151
R1826 B.n964 B.n99 10.6151
R1827 B.n964 B.n963 10.6151
R1828 B.n963 B.n962 10.6151
R1829 B.n962 B.n101 10.6151
R1830 B.n956 B.n101 10.6151
R1831 B.n956 B.n955 10.6151
R1832 B.n955 B.n954 10.6151
R1833 B.n954 B.n103 10.6151
R1834 B.n948 B.n103 10.6151
R1835 B.n948 B.n947 10.6151
R1836 B.n947 B.n946 10.6151
R1837 B.n946 B.n105 10.6151
R1838 B.n940 B.n105 10.6151
R1839 B.n940 B.n939 10.6151
R1840 B.n939 B.n938 10.6151
R1841 B.n938 B.n107 10.6151
R1842 B.n932 B.n107 10.6151
R1843 B.n932 B.n931 10.6151
R1844 B.n931 B.n930 10.6151
R1845 B.n930 B.n109 10.6151
R1846 B.n924 B.n109 10.6151
R1847 B.n924 B.n923 10.6151
R1848 B.n923 B.n922 10.6151
R1849 B.n922 B.n111 10.6151
R1850 B.n916 B.n111 10.6151
R1851 B.n914 B.n913 10.6151
R1852 B.n913 B.n115 10.6151
R1853 B.n907 B.n115 10.6151
R1854 B.n907 B.n906 10.6151
R1855 B.n906 B.n905 10.6151
R1856 B.n905 B.n117 10.6151
R1857 B.n899 B.n117 10.6151
R1858 B.n899 B.n898 10.6151
R1859 B.n898 B.n897 10.6151
R1860 B.n893 B.n892 10.6151
R1861 B.n892 B.n123 10.6151
R1862 B.n887 B.n123 10.6151
R1863 B.n887 B.n886 10.6151
R1864 B.n886 B.n885 10.6151
R1865 B.n885 B.n125 10.6151
R1866 B.n879 B.n125 10.6151
R1867 B.n879 B.n878 10.6151
R1868 B.n878 B.n877 10.6151
R1869 B.n877 B.n127 10.6151
R1870 B.n871 B.n127 10.6151
R1871 B.n871 B.n870 10.6151
R1872 B.n870 B.n869 10.6151
R1873 B.n869 B.n129 10.6151
R1874 B.n863 B.n129 10.6151
R1875 B.n863 B.n862 10.6151
R1876 B.n862 B.n861 10.6151
R1877 B.n861 B.n131 10.6151
R1878 B.n855 B.n131 10.6151
R1879 B.n855 B.n854 10.6151
R1880 B.n854 B.n853 10.6151
R1881 B.n853 B.n133 10.6151
R1882 B.n847 B.n133 10.6151
R1883 B.n847 B.n846 10.6151
R1884 B.n846 B.n845 10.6151
R1885 B.n845 B.n135 10.6151
R1886 B.n839 B.n135 10.6151
R1887 B.n839 B.n838 10.6151
R1888 B.n838 B.n837 10.6151
R1889 B.n837 B.n137 10.6151
R1890 B.n831 B.n137 10.6151
R1891 B.n831 B.n830 10.6151
R1892 B.n830 B.n829 10.6151
R1893 B.n829 B.n139 10.6151
R1894 B.n823 B.n139 10.6151
R1895 B.n823 B.n822 10.6151
R1896 B.n822 B.n821 10.6151
R1897 B.n821 B.n141 10.6151
R1898 B.n815 B.n141 10.6151
R1899 B.n815 B.n814 10.6151
R1900 B.n814 B.n813 10.6151
R1901 B.n813 B.n143 10.6151
R1902 B.n807 B.n143 10.6151
R1903 B.n807 B.n806 10.6151
R1904 B.n806 B.n805 10.6151
R1905 B.n805 B.n145 10.6151
R1906 B.n799 B.n145 10.6151
R1907 B.n799 B.n798 10.6151
R1908 B.n798 B.n797 10.6151
R1909 B.n797 B.n147 10.6151
R1910 B.n791 B.n147 10.6151
R1911 B.n791 B.n790 10.6151
R1912 B.n790 B.n789 10.6151
R1913 B.n789 B.n149 10.6151
R1914 B.n783 B.n149 10.6151
R1915 B.n783 B.n782 10.6151
R1916 B.n782 B.n781 10.6151
R1917 B.n781 B.n151 10.6151
R1918 B.n775 B.n151 10.6151
R1919 B.n775 B.n774 10.6151
R1920 B.n774 B.n773 10.6151
R1921 B.n773 B.n153 10.6151
R1922 B.n767 B.n153 10.6151
R1923 B.n457 B.n456 9.36635
R1924 B.n433 B.n278 9.36635
R1925 B.n916 B.n915 9.36635
R1926 B.n893 B.n121 9.36635
R1927 B.n1132 B.n0 8.11757
R1928 B.n1132 B.n1 8.11757
R1929 B.n658 B.t0 7.91892
R1930 B.n1094 B.t1 7.91892
R1931 B.n688 B.t2 5.27944
R1932 B.n19 B.t3 5.27944
R1933 B.n218 B.t5 2.63997
R1934 B.t12 B.n1063 2.63997
R1935 B.n456 B.n455 1.24928
R1936 B.n278 B.n274 1.24928
R1937 B.n915 B.n914 1.24928
R1938 B.n897 B.n121 1.24928
R1939 VP.n5 VP.t2 168.275
R1940 VP.n5 VP.t0 167.041
R1941 VP.n19 VP.n18 161.3
R1942 VP.n17 VP.n1 161.3
R1943 VP.n16 VP.n15 161.3
R1944 VP.n14 VP.n2 161.3
R1945 VP.n13 VP.n12 161.3
R1946 VP.n11 VP.n3 161.3
R1947 VP.n10 VP.n9 161.3
R1948 VP.n8 VP.n4 161.3
R1949 VP.n6 VP.t3 133.565
R1950 VP.n0 VP.t1 133.565
R1951 VP.n7 VP.n6 80.5253
R1952 VP.n20 VP.n0 80.5253
R1953 VP.n7 VP.n5 57.3187
R1954 VP.n12 VP.n2 56.5193
R1955 VP.n10 VP.n4 24.4675
R1956 VP.n11 VP.n10 24.4675
R1957 VP.n12 VP.n11 24.4675
R1958 VP.n16 VP.n2 24.4675
R1959 VP.n17 VP.n16 24.4675
R1960 VP.n18 VP.n17 24.4675
R1961 VP.n6 VP.n4 9.54263
R1962 VP.n18 VP.n0 9.54263
R1963 VP.n8 VP.n7 0.354971
R1964 VP.n20 VP.n19 0.354971
R1965 VP VP.n20 0.26696
R1966 VP.n9 VP.n8 0.189894
R1967 VP.n9 VP.n3 0.189894
R1968 VP.n13 VP.n3 0.189894
R1969 VP.n14 VP.n13 0.189894
R1970 VP.n15 VP.n14 0.189894
R1971 VP.n15 VP.n1 0.189894
R1972 VP.n19 VP.n1 0.189894
R1973 VDD1 VDD1.n1 112.483
R1974 VDD1 VDD1.n0 61.2326
R1975 VDD1.n0 VDD1.t1 1.00405
R1976 VDD1.n0 VDD1.t3 1.00405
R1977 VDD1.n1 VDD1.t0 1.00405
R1978 VDD1.n1 VDD1.t2 1.00405
C0 VDD2 VDD1 1.25721f
C1 VTAIL VDD1 7.30433f
C2 VDD2 VTAIL 7.36497f
C3 VP VDD1 8.29559f
C4 VN VDD1 0.150019f
C5 VDD2 VP 0.455543f
C6 VDD2 VN 7.991049f
C7 VTAIL VP 7.69669f
C8 VN VTAIL 7.68258f
C9 VN VP 8.314361f
C10 VDD2 B 4.916161f
C11 VDD1 B 10.15166f
C12 VTAIL B 15.303256f
C13 VN B 13.15784f
C14 VP B 11.49858f
C15 VDD1.t1 B 0.418521f
C16 VDD1.t3 B 0.418521f
C17 VDD1.n0 B 3.83294f
C18 VDD1.t0 B 0.418521f
C19 VDD1.t2 B 0.418521f
C20 VDD1.n1 B 4.8893f
C21 VP.t1 B 3.78394f
C22 VP.n0 B 1.37709f
C23 VP.n1 B 0.019554f
C24 VP.n2 B 0.028545f
C25 VP.n3 B 0.019554f
C26 VP.n4 B 0.025467f
C27 VP.t2 B 4.08413f
C28 VP.t0 B 4.07388f
C29 VP.n5 B 3.93612f
C30 VP.t3 B 3.78394f
C31 VP.n6 B 1.37709f
C32 VP.n7 B 1.35509f
C33 VP.n8 B 0.031559f
C34 VP.n9 B 0.019554f
C35 VP.n10 B 0.036443f
C36 VP.n11 B 0.036443f
C37 VP.n12 B 0.028545f
C38 VP.n13 B 0.019554f
C39 VP.n14 B 0.019554f
C40 VP.n15 B 0.019554f
C41 VP.n16 B 0.036443f
C42 VP.n17 B 0.036443f
C43 VP.n18 B 0.025467f
C44 VP.n19 B 0.031559f
C45 VP.n20 B 0.053395f
C46 VTAIL.t7 B 2.76348f
C47 VTAIL.n0 B 0.317493f
C48 VTAIL.t2 B 2.76348f
C49 VTAIL.n1 B 0.398171f
C50 VTAIL.t0 B 2.76348f
C51 VTAIL.n2 B 1.59986f
C52 VTAIL.t5 B 2.76348f
C53 VTAIL.n3 B 1.59986f
C54 VTAIL.t4 B 2.76348f
C55 VTAIL.n4 B 0.398171f
C56 VTAIL.t3 B 2.76348f
C57 VTAIL.n5 B 0.398171f
C58 VTAIL.t1 B 2.76348f
C59 VTAIL.n6 B 1.59986f
C60 VTAIL.t6 B 2.76348f
C61 VTAIL.n7 B 1.51338f
C62 VDD2.t2 B 0.415798f
C63 VDD2.t1 B 0.415798f
C64 VDD2.n0 B 4.82808f
C65 VDD2.t0 B 0.415798f
C66 VDD2.t3 B 0.415798f
C67 VDD2.n1 B 3.80751f
C68 VDD2.n2 B 4.8073f
C69 VN.t1 B 4.01904f
C70 VN.t0 B 4.02915f
C71 VN.n0 B 2.47022f
C72 VN.t3 B 4.02915f
C73 VN.t2 B 4.01904f
C74 VN.n1 B 3.89065f
.ends

