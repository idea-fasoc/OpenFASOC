* NGSPICE file created from diff_pair_sample_0171.ext - technology: sky130A

.subckt diff_pair_sample_0171 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2100_n3922# sky130_fd_pr__pfet_01v8 ad=5.7603 pd=30.32 as=0 ps=0 w=14.77 l=0.8
X1 VDD1.t7 VP.t0 VTAIL.t14 w_n2100_n3922# sky130_fd_pr__pfet_01v8 ad=2.43705 pd=15.1 as=5.7603 ps=30.32 w=14.77 l=0.8
X2 B.t8 B.t6 B.t7 w_n2100_n3922# sky130_fd_pr__pfet_01v8 ad=5.7603 pd=30.32 as=0 ps=0 w=14.77 l=0.8
X3 VTAIL.t5 VN.t0 VDD2.t7 w_n2100_n3922# sky130_fd_pr__pfet_01v8 ad=5.7603 pd=30.32 as=2.43705 ps=15.1 w=14.77 l=0.8
X4 B.t5 B.t3 B.t4 w_n2100_n3922# sky130_fd_pr__pfet_01v8 ad=5.7603 pd=30.32 as=0 ps=0 w=14.77 l=0.8
X5 VDD2.t6 VN.t1 VTAIL.t6 w_n2100_n3922# sky130_fd_pr__pfet_01v8 ad=2.43705 pd=15.1 as=2.43705 ps=15.1 w=14.77 l=0.8
X6 VTAIL.t7 VN.t2 VDD2.t5 w_n2100_n3922# sky130_fd_pr__pfet_01v8 ad=2.43705 pd=15.1 as=2.43705 ps=15.1 w=14.77 l=0.8
X7 VDD2.t4 VN.t3 VTAIL.t3 w_n2100_n3922# sky130_fd_pr__pfet_01v8 ad=2.43705 pd=15.1 as=5.7603 ps=30.32 w=14.77 l=0.8
X8 VTAIL.t2 VN.t4 VDD2.t3 w_n2100_n3922# sky130_fd_pr__pfet_01v8 ad=5.7603 pd=30.32 as=2.43705 ps=15.1 w=14.77 l=0.8
X9 VDD2.t2 VN.t5 VTAIL.t4 w_n2100_n3922# sky130_fd_pr__pfet_01v8 ad=2.43705 pd=15.1 as=5.7603 ps=30.32 w=14.77 l=0.8
X10 VTAIL.t13 VP.t1 VDD1.t6 w_n2100_n3922# sky130_fd_pr__pfet_01v8 ad=5.7603 pd=30.32 as=2.43705 ps=15.1 w=14.77 l=0.8
X11 VDD1.t5 VP.t2 VTAIL.t8 w_n2100_n3922# sky130_fd_pr__pfet_01v8 ad=2.43705 pd=15.1 as=5.7603 ps=30.32 w=14.77 l=0.8
X12 VTAIL.t11 VP.t3 VDD1.t4 w_n2100_n3922# sky130_fd_pr__pfet_01v8 ad=2.43705 pd=15.1 as=2.43705 ps=15.1 w=14.77 l=0.8
X13 VTAIL.t9 VP.t4 VDD1.t3 w_n2100_n3922# sky130_fd_pr__pfet_01v8 ad=2.43705 pd=15.1 as=2.43705 ps=15.1 w=14.77 l=0.8
X14 VDD2.t1 VN.t6 VTAIL.t0 w_n2100_n3922# sky130_fd_pr__pfet_01v8 ad=2.43705 pd=15.1 as=2.43705 ps=15.1 w=14.77 l=0.8
X15 VDD1.t2 VP.t5 VTAIL.t10 w_n2100_n3922# sky130_fd_pr__pfet_01v8 ad=2.43705 pd=15.1 as=2.43705 ps=15.1 w=14.77 l=0.8
X16 VTAIL.t12 VP.t6 VDD1.t1 w_n2100_n3922# sky130_fd_pr__pfet_01v8 ad=5.7603 pd=30.32 as=2.43705 ps=15.1 w=14.77 l=0.8
X17 B.t2 B.t0 B.t1 w_n2100_n3922# sky130_fd_pr__pfet_01v8 ad=5.7603 pd=30.32 as=0 ps=0 w=14.77 l=0.8
X18 VDD1.t0 VP.t7 VTAIL.t15 w_n2100_n3922# sky130_fd_pr__pfet_01v8 ad=2.43705 pd=15.1 as=2.43705 ps=15.1 w=14.77 l=0.8
X19 VTAIL.t1 VN.t7 VDD2.t0 w_n2100_n3922# sky130_fd_pr__pfet_01v8 ad=2.43705 pd=15.1 as=2.43705 ps=15.1 w=14.77 l=0.8
R0 B.n128 B.t3 646.836
R1 B.n288 B.t9 646.836
R2 B.n46 B.t0 646.836
R3 B.n40 B.t6 646.836
R4 B.n367 B.n366 585
R5 B.n365 B.n98 585
R6 B.n364 B.n363 585
R7 B.n362 B.n99 585
R8 B.n361 B.n360 585
R9 B.n359 B.n100 585
R10 B.n358 B.n357 585
R11 B.n356 B.n101 585
R12 B.n355 B.n354 585
R13 B.n353 B.n102 585
R14 B.n352 B.n351 585
R15 B.n350 B.n103 585
R16 B.n349 B.n348 585
R17 B.n347 B.n104 585
R18 B.n346 B.n345 585
R19 B.n344 B.n105 585
R20 B.n343 B.n342 585
R21 B.n341 B.n106 585
R22 B.n340 B.n339 585
R23 B.n338 B.n107 585
R24 B.n337 B.n336 585
R25 B.n335 B.n108 585
R26 B.n334 B.n333 585
R27 B.n332 B.n109 585
R28 B.n331 B.n330 585
R29 B.n329 B.n110 585
R30 B.n328 B.n327 585
R31 B.n326 B.n111 585
R32 B.n325 B.n324 585
R33 B.n323 B.n112 585
R34 B.n322 B.n321 585
R35 B.n320 B.n113 585
R36 B.n319 B.n318 585
R37 B.n317 B.n114 585
R38 B.n316 B.n315 585
R39 B.n314 B.n115 585
R40 B.n313 B.n312 585
R41 B.n311 B.n116 585
R42 B.n310 B.n309 585
R43 B.n308 B.n117 585
R44 B.n307 B.n306 585
R45 B.n305 B.n118 585
R46 B.n304 B.n303 585
R47 B.n302 B.n119 585
R48 B.n301 B.n300 585
R49 B.n299 B.n120 585
R50 B.n298 B.n297 585
R51 B.n296 B.n121 585
R52 B.n295 B.n294 585
R53 B.n293 B.n122 585
R54 B.n292 B.n291 585
R55 B.n287 B.n123 585
R56 B.n286 B.n285 585
R57 B.n284 B.n124 585
R58 B.n283 B.n282 585
R59 B.n281 B.n125 585
R60 B.n280 B.n279 585
R61 B.n278 B.n126 585
R62 B.n277 B.n276 585
R63 B.n274 B.n127 585
R64 B.n273 B.n272 585
R65 B.n271 B.n130 585
R66 B.n270 B.n269 585
R67 B.n268 B.n131 585
R68 B.n267 B.n266 585
R69 B.n265 B.n132 585
R70 B.n264 B.n263 585
R71 B.n262 B.n133 585
R72 B.n261 B.n260 585
R73 B.n259 B.n134 585
R74 B.n258 B.n257 585
R75 B.n256 B.n135 585
R76 B.n255 B.n254 585
R77 B.n253 B.n136 585
R78 B.n252 B.n251 585
R79 B.n250 B.n137 585
R80 B.n249 B.n248 585
R81 B.n247 B.n138 585
R82 B.n246 B.n245 585
R83 B.n244 B.n139 585
R84 B.n243 B.n242 585
R85 B.n241 B.n140 585
R86 B.n240 B.n239 585
R87 B.n238 B.n141 585
R88 B.n237 B.n236 585
R89 B.n235 B.n142 585
R90 B.n234 B.n233 585
R91 B.n232 B.n143 585
R92 B.n231 B.n230 585
R93 B.n229 B.n144 585
R94 B.n228 B.n227 585
R95 B.n226 B.n145 585
R96 B.n225 B.n224 585
R97 B.n223 B.n146 585
R98 B.n222 B.n221 585
R99 B.n220 B.n147 585
R100 B.n219 B.n218 585
R101 B.n217 B.n148 585
R102 B.n216 B.n215 585
R103 B.n214 B.n149 585
R104 B.n213 B.n212 585
R105 B.n211 B.n150 585
R106 B.n210 B.n209 585
R107 B.n208 B.n151 585
R108 B.n207 B.n206 585
R109 B.n205 B.n152 585
R110 B.n204 B.n203 585
R111 B.n202 B.n153 585
R112 B.n201 B.n200 585
R113 B.n368 B.n97 585
R114 B.n370 B.n369 585
R115 B.n371 B.n96 585
R116 B.n373 B.n372 585
R117 B.n374 B.n95 585
R118 B.n376 B.n375 585
R119 B.n377 B.n94 585
R120 B.n379 B.n378 585
R121 B.n380 B.n93 585
R122 B.n382 B.n381 585
R123 B.n383 B.n92 585
R124 B.n385 B.n384 585
R125 B.n386 B.n91 585
R126 B.n388 B.n387 585
R127 B.n389 B.n90 585
R128 B.n391 B.n390 585
R129 B.n392 B.n89 585
R130 B.n394 B.n393 585
R131 B.n395 B.n88 585
R132 B.n397 B.n396 585
R133 B.n398 B.n87 585
R134 B.n400 B.n399 585
R135 B.n401 B.n86 585
R136 B.n403 B.n402 585
R137 B.n404 B.n85 585
R138 B.n406 B.n405 585
R139 B.n407 B.n84 585
R140 B.n409 B.n408 585
R141 B.n410 B.n83 585
R142 B.n412 B.n411 585
R143 B.n413 B.n82 585
R144 B.n415 B.n414 585
R145 B.n416 B.n81 585
R146 B.n418 B.n417 585
R147 B.n419 B.n80 585
R148 B.n421 B.n420 585
R149 B.n422 B.n79 585
R150 B.n424 B.n423 585
R151 B.n425 B.n78 585
R152 B.n427 B.n426 585
R153 B.n428 B.n77 585
R154 B.n430 B.n429 585
R155 B.n431 B.n76 585
R156 B.n433 B.n432 585
R157 B.n434 B.n75 585
R158 B.n436 B.n435 585
R159 B.n437 B.n74 585
R160 B.n439 B.n438 585
R161 B.n440 B.n73 585
R162 B.n442 B.n441 585
R163 B.n607 B.n14 585
R164 B.n606 B.n605 585
R165 B.n604 B.n15 585
R166 B.n603 B.n602 585
R167 B.n601 B.n16 585
R168 B.n600 B.n599 585
R169 B.n598 B.n17 585
R170 B.n597 B.n596 585
R171 B.n595 B.n18 585
R172 B.n594 B.n593 585
R173 B.n592 B.n19 585
R174 B.n591 B.n590 585
R175 B.n589 B.n20 585
R176 B.n588 B.n587 585
R177 B.n586 B.n21 585
R178 B.n585 B.n584 585
R179 B.n583 B.n22 585
R180 B.n582 B.n581 585
R181 B.n580 B.n23 585
R182 B.n579 B.n578 585
R183 B.n577 B.n24 585
R184 B.n576 B.n575 585
R185 B.n574 B.n25 585
R186 B.n573 B.n572 585
R187 B.n571 B.n26 585
R188 B.n570 B.n569 585
R189 B.n568 B.n27 585
R190 B.n567 B.n566 585
R191 B.n565 B.n28 585
R192 B.n564 B.n563 585
R193 B.n562 B.n29 585
R194 B.n561 B.n560 585
R195 B.n559 B.n30 585
R196 B.n558 B.n557 585
R197 B.n556 B.n31 585
R198 B.n555 B.n554 585
R199 B.n553 B.n32 585
R200 B.n552 B.n551 585
R201 B.n550 B.n33 585
R202 B.n549 B.n548 585
R203 B.n547 B.n34 585
R204 B.n546 B.n545 585
R205 B.n544 B.n35 585
R206 B.n543 B.n542 585
R207 B.n541 B.n36 585
R208 B.n540 B.n539 585
R209 B.n538 B.n37 585
R210 B.n537 B.n536 585
R211 B.n535 B.n38 585
R212 B.n534 B.n533 585
R213 B.n531 B.n39 585
R214 B.n530 B.n529 585
R215 B.n528 B.n42 585
R216 B.n527 B.n526 585
R217 B.n525 B.n43 585
R218 B.n524 B.n523 585
R219 B.n522 B.n44 585
R220 B.n521 B.n520 585
R221 B.n519 B.n45 585
R222 B.n517 B.n516 585
R223 B.n515 B.n48 585
R224 B.n514 B.n513 585
R225 B.n512 B.n49 585
R226 B.n511 B.n510 585
R227 B.n509 B.n50 585
R228 B.n508 B.n507 585
R229 B.n506 B.n51 585
R230 B.n505 B.n504 585
R231 B.n503 B.n52 585
R232 B.n502 B.n501 585
R233 B.n500 B.n53 585
R234 B.n499 B.n498 585
R235 B.n497 B.n54 585
R236 B.n496 B.n495 585
R237 B.n494 B.n55 585
R238 B.n493 B.n492 585
R239 B.n491 B.n56 585
R240 B.n490 B.n489 585
R241 B.n488 B.n57 585
R242 B.n487 B.n486 585
R243 B.n485 B.n58 585
R244 B.n484 B.n483 585
R245 B.n482 B.n59 585
R246 B.n481 B.n480 585
R247 B.n479 B.n60 585
R248 B.n478 B.n477 585
R249 B.n476 B.n61 585
R250 B.n475 B.n474 585
R251 B.n473 B.n62 585
R252 B.n472 B.n471 585
R253 B.n470 B.n63 585
R254 B.n469 B.n468 585
R255 B.n467 B.n64 585
R256 B.n466 B.n465 585
R257 B.n464 B.n65 585
R258 B.n463 B.n462 585
R259 B.n461 B.n66 585
R260 B.n460 B.n459 585
R261 B.n458 B.n67 585
R262 B.n457 B.n456 585
R263 B.n455 B.n68 585
R264 B.n454 B.n453 585
R265 B.n452 B.n69 585
R266 B.n451 B.n450 585
R267 B.n449 B.n70 585
R268 B.n448 B.n447 585
R269 B.n446 B.n71 585
R270 B.n445 B.n444 585
R271 B.n443 B.n72 585
R272 B.n609 B.n608 585
R273 B.n610 B.n13 585
R274 B.n612 B.n611 585
R275 B.n613 B.n12 585
R276 B.n615 B.n614 585
R277 B.n616 B.n11 585
R278 B.n618 B.n617 585
R279 B.n619 B.n10 585
R280 B.n621 B.n620 585
R281 B.n622 B.n9 585
R282 B.n624 B.n623 585
R283 B.n625 B.n8 585
R284 B.n627 B.n626 585
R285 B.n628 B.n7 585
R286 B.n630 B.n629 585
R287 B.n631 B.n6 585
R288 B.n633 B.n632 585
R289 B.n634 B.n5 585
R290 B.n636 B.n635 585
R291 B.n637 B.n4 585
R292 B.n639 B.n638 585
R293 B.n640 B.n3 585
R294 B.n642 B.n641 585
R295 B.n643 B.n0 585
R296 B.n2 B.n1 585
R297 B.n166 B.n165 585
R298 B.n168 B.n167 585
R299 B.n169 B.n164 585
R300 B.n171 B.n170 585
R301 B.n172 B.n163 585
R302 B.n174 B.n173 585
R303 B.n175 B.n162 585
R304 B.n177 B.n176 585
R305 B.n178 B.n161 585
R306 B.n180 B.n179 585
R307 B.n181 B.n160 585
R308 B.n183 B.n182 585
R309 B.n184 B.n159 585
R310 B.n186 B.n185 585
R311 B.n187 B.n158 585
R312 B.n189 B.n188 585
R313 B.n190 B.n157 585
R314 B.n192 B.n191 585
R315 B.n193 B.n156 585
R316 B.n195 B.n194 585
R317 B.n196 B.n155 585
R318 B.n198 B.n197 585
R319 B.n199 B.n154 585
R320 B.n200 B.n199 545.355
R321 B.n366 B.n97 545.355
R322 B.n443 B.n442 545.355
R323 B.n608 B.n607 545.355
R324 B.n288 B.t10 447.406
R325 B.n46 B.t2 447.406
R326 B.n128 B.t4 447.406
R327 B.n40 B.t8 447.406
R328 B.n289 B.t11 425.49
R329 B.n47 B.t1 425.49
R330 B.n129 B.t5 425.49
R331 B.n41 B.t7 425.49
R332 B.n645 B.n644 256.663
R333 B.n644 B.n643 235.042
R334 B.n644 B.n2 235.042
R335 B.n200 B.n153 163.367
R336 B.n204 B.n153 163.367
R337 B.n205 B.n204 163.367
R338 B.n206 B.n205 163.367
R339 B.n206 B.n151 163.367
R340 B.n210 B.n151 163.367
R341 B.n211 B.n210 163.367
R342 B.n212 B.n211 163.367
R343 B.n212 B.n149 163.367
R344 B.n216 B.n149 163.367
R345 B.n217 B.n216 163.367
R346 B.n218 B.n217 163.367
R347 B.n218 B.n147 163.367
R348 B.n222 B.n147 163.367
R349 B.n223 B.n222 163.367
R350 B.n224 B.n223 163.367
R351 B.n224 B.n145 163.367
R352 B.n228 B.n145 163.367
R353 B.n229 B.n228 163.367
R354 B.n230 B.n229 163.367
R355 B.n230 B.n143 163.367
R356 B.n234 B.n143 163.367
R357 B.n235 B.n234 163.367
R358 B.n236 B.n235 163.367
R359 B.n236 B.n141 163.367
R360 B.n240 B.n141 163.367
R361 B.n241 B.n240 163.367
R362 B.n242 B.n241 163.367
R363 B.n242 B.n139 163.367
R364 B.n246 B.n139 163.367
R365 B.n247 B.n246 163.367
R366 B.n248 B.n247 163.367
R367 B.n248 B.n137 163.367
R368 B.n252 B.n137 163.367
R369 B.n253 B.n252 163.367
R370 B.n254 B.n253 163.367
R371 B.n254 B.n135 163.367
R372 B.n258 B.n135 163.367
R373 B.n259 B.n258 163.367
R374 B.n260 B.n259 163.367
R375 B.n260 B.n133 163.367
R376 B.n264 B.n133 163.367
R377 B.n265 B.n264 163.367
R378 B.n266 B.n265 163.367
R379 B.n266 B.n131 163.367
R380 B.n270 B.n131 163.367
R381 B.n271 B.n270 163.367
R382 B.n272 B.n271 163.367
R383 B.n272 B.n127 163.367
R384 B.n277 B.n127 163.367
R385 B.n278 B.n277 163.367
R386 B.n279 B.n278 163.367
R387 B.n279 B.n125 163.367
R388 B.n283 B.n125 163.367
R389 B.n284 B.n283 163.367
R390 B.n285 B.n284 163.367
R391 B.n285 B.n123 163.367
R392 B.n292 B.n123 163.367
R393 B.n293 B.n292 163.367
R394 B.n294 B.n293 163.367
R395 B.n294 B.n121 163.367
R396 B.n298 B.n121 163.367
R397 B.n299 B.n298 163.367
R398 B.n300 B.n299 163.367
R399 B.n300 B.n119 163.367
R400 B.n304 B.n119 163.367
R401 B.n305 B.n304 163.367
R402 B.n306 B.n305 163.367
R403 B.n306 B.n117 163.367
R404 B.n310 B.n117 163.367
R405 B.n311 B.n310 163.367
R406 B.n312 B.n311 163.367
R407 B.n312 B.n115 163.367
R408 B.n316 B.n115 163.367
R409 B.n317 B.n316 163.367
R410 B.n318 B.n317 163.367
R411 B.n318 B.n113 163.367
R412 B.n322 B.n113 163.367
R413 B.n323 B.n322 163.367
R414 B.n324 B.n323 163.367
R415 B.n324 B.n111 163.367
R416 B.n328 B.n111 163.367
R417 B.n329 B.n328 163.367
R418 B.n330 B.n329 163.367
R419 B.n330 B.n109 163.367
R420 B.n334 B.n109 163.367
R421 B.n335 B.n334 163.367
R422 B.n336 B.n335 163.367
R423 B.n336 B.n107 163.367
R424 B.n340 B.n107 163.367
R425 B.n341 B.n340 163.367
R426 B.n342 B.n341 163.367
R427 B.n342 B.n105 163.367
R428 B.n346 B.n105 163.367
R429 B.n347 B.n346 163.367
R430 B.n348 B.n347 163.367
R431 B.n348 B.n103 163.367
R432 B.n352 B.n103 163.367
R433 B.n353 B.n352 163.367
R434 B.n354 B.n353 163.367
R435 B.n354 B.n101 163.367
R436 B.n358 B.n101 163.367
R437 B.n359 B.n358 163.367
R438 B.n360 B.n359 163.367
R439 B.n360 B.n99 163.367
R440 B.n364 B.n99 163.367
R441 B.n365 B.n364 163.367
R442 B.n366 B.n365 163.367
R443 B.n442 B.n73 163.367
R444 B.n438 B.n73 163.367
R445 B.n438 B.n437 163.367
R446 B.n437 B.n436 163.367
R447 B.n436 B.n75 163.367
R448 B.n432 B.n75 163.367
R449 B.n432 B.n431 163.367
R450 B.n431 B.n430 163.367
R451 B.n430 B.n77 163.367
R452 B.n426 B.n77 163.367
R453 B.n426 B.n425 163.367
R454 B.n425 B.n424 163.367
R455 B.n424 B.n79 163.367
R456 B.n420 B.n79 163.367
R457 B.n420 B.n419 163.367
R458 B.n419 B.n418 163.367
R459 B.n418 B.n81 163.367
R460 B.n414 B.n81 163.367
R461 B.n414 B.n413 163.367
R462 B.n413 B.n412 163.367
R463 B.n412 B.n83 163.367
R464 B.n408 B.n83 163.367
R465 B.n408 B.n407 163.367
R466 B.n407 B.n406 163.367
R467 B.n406 B.n85 163.367
R468 B.n402 B.n85 163.367
R469 B.n402 B.n401 163.367
R470 B.n401 B.n400 163.367
R471 B.n400 B.n87 163.367
R472 B.n396 B.n87 163.367
R473 B.n396 B.n395 163.367
R474 B.n395 B.n394 163.367
R475 B.n394 B.n89 163.367
R476 B.n390 B.n89 163.367
R477 B.n390 B.n389 163.367
R478 B.n389 B.n388 163.367
R479 B.n388 B.n91 163.367
R480 B.n384 B.n91 163.367
R481 B.n384 B.n383 163.367
R482 B.n383 B.n382 163.367
R483 B.n382 B.n93 163.367
R484 B.n378 B.n93 163.367
R485 B.n378 B.n377 163.367
R486 B.n377 B.n376 163.367
R487 B.n376 B.n95 163.367
R488 B.n372 B.n95 163.367
R489 B.n372 B.n371 163.367
R490 B.n371 B.n370 163.367
R491 B.n370 B.n97 163.367
R492 B.n607 B.n606 163.367
R493 B.n606 B.n15 163.367
R494 B.n602 B.n15 163.367
R495 B.n602 B.n601 163.367
R496 B.n601 B.n600 163.367
R497 B.n600 B.n17 163.367
R498 B.n596 B.n17 163.367
R499 B.n596 B.n595 163.367
R500 B.n595 B.n594 163.367
R501 B.n594 B.n19 163.367
R502 B.n590 B.n19 163.367
R503 B.n590 B.n589 163.367
R504 B.n589 B.n588 163.367
R505 B.n588 B.n21 163.367
R506 B.n584 B.n21 163.367
R507 B.n584 B.n583 163.367
R508 B.n583 B.n582 163.367
R509 B.n582 B.n23 163.367
R510 B.n578 B.n23 163.367
R511 B.n578 B.n577 163.367
R512 B.n577 B.n576 163.367
R513 B.n576 B.n25 163.367
R514 B.n572 B.n25 163.367
R515 B.n572 B.n571 163.367
R516 B.n571 B.n570 163.367
R517 B.n570 B.n27 163.367
R518 B.n566 B.n27 163.367
R519 B.n566 B.n565 163.367
R520 B.n565 B.n564 163.367
R521 B.n564 B.n29 163.367
R522 B.n560 B.n29 163.367
R523 B.n560 B.n559 163.367
R524 B.n559 B.n558 163.367
R525 B.n558 B.n31 163.367
R526 B.n554 B.n31 163.367
R527 B.n554 B.n553 163.367
R528 B.n553 B.n552 163.367
R529 B.n552 B.n33 163.367
R530 B.n548 B.n33 163.367
R531 B.n548 B.n547 163.367
R532 B.n547 B.n546 163.367
R533 B.n546 B.n35 163.367
R534 B.n542 B.n35 163.367
R535 B.n542 B.n541 163.367
R536 B.n541 B.n540 163.367
R537 B.n540 B.n37 163.367
R538 B.n536 B.n37 163.367
R539 B.n536 B.n535 163.367
R540 B.n535 B.n534 163.367
R541 B.n534 B.n39 163.367
R542 B.n529 B.n39 163.367
R543 B.n529 B.n528 163.367
R544 B.n528 B.n527 163.367
R545 B.n527 B.n43 163.367
R546 B.n523 B.n43 163.367
R547 B.n523 B.n522 163.367
R548 B.n522 B.n521 163.367
R549 B.n521 B.n45 163.367
R550 B.n516 B.n45 163.367
R551 B.n516 B.n515 163.367
R552 B.n515 B.n514 163.367
R553 B.n514 B.n49 163.367
R554 B.n510 B.n49 163.367
R555 B.n510 B.n509 163.367
R556 B.n509 B.n508 163.367
R557 B.n508 B.n51 163.367
R558 B.n504 B.n51 163.367
R559 B.n504 B.n503 163.367
R560 B.n503 B.n502 163.367
R561 B.n502 B.n53 163.367
R562 B.n498 B.n53 163.367
R563 B.n498 B.n497 163.367
R564 B.n497 B.n496 163.367
R565 B.n496 B.n55 163.367
R566 B.n492 B.n55 163.367
R567 B.n492 B.n491 163.367
R568 B.n491 B.n490 163.367
R569 B.n490 B.n57 163.367
R570 B.n486 B.n57 163.367
R571 B.n486 B.n485 163.367
R572 B.n485 B.n484 163.367
R573 B.n484 B.n59 163.367
R574 B.n480 B.n59 163.367
R575 B.n480 B.n479 163.367
R576 B.n479 B.n478 163.367
R577 B.n478 B.n61 163.367
R578 B.n474 B.n61 163.367
R579 B.n474 B.n473 163.367
R580 B.n473 B.n472 163.367
R581 B.n472 B.n63 163.367
R582 B.n468 B.n63 163.367
R583 B.n468 B.n467 163.367
R584 B.n467 B.n466 163.367
R585 B.n466 B.n65 163.367
R586 B.n462 B.n65 163.367
R587 B.n462 B.n461 163.367
R588 B.n461 B.n460 163.367
R589 B.n460 B.n67 163.367
R590 B.n456 B.n67 163.367
R591 B.n456 B.n455 163.367
R592 B.n455 B.n454 163.367
R593 B.n454 B.n69 163.367
R594 B.n450 B.n69 163.367
R595 B.n450 B.n449 163.367
R596 B.n449 B.n448 163.367
R597 B.n448 B.n71 163.367
R598 B.n444 B.n71 163.367
R599 B.n444 B.n443 163.367
R600 B.n608 B.n13 163.367
R601 B.n612 B.n13 163.367
R602 B.n613 B.n612 163.367
R603 B.n614 B.n613 163.367
R604 B.n614 B.n11 163.367
R605 B.n618 B.n11 163.367
R606 B.n619 B.n618 163.367
R607 B.n620 B.n619 163.367
R608 B.n620 B.n9 163.367
R609 B.n624 B.n9 163.367
R610 B.n625 B.n624 163.367
R611 B.n626 B.n625 163.367
R612 B.n626 B.n7 163.367
R613 B.n630 B.n7 163.367
R614 B.n631 B.n630 163.367
R615 B.n632 B.n631 163.367
R616 B.n632 B.n5 163.367
R617 B.n636 B.n5 163.367
R618 B.n637 B.n636 163.367
R619 B.n638 B.n637 163.367
R620 B.n638 B.n3 163.367
R621 B.n642 B.n3 163.367
R622 B.n643 B.n642 163.367
R623 B.n165 B.n2 163.367
R624 B.n168 B.n165 163.367
R625 B.n169 B.n168 163.367
R626 B.n170 B.n169 163.367
R627 B.n170 B.n163 163.367
R628 B.n174 B.n163 163.367
R629 B.n175 B.n174 163.367
R630 B.n176 B.n175 163.367
R631 B.n176 B.n161 163.367
R632 B.n180 B.n161 163.367
R633 B.n181 B.n180 163.367
R634 B.n182 B.n181 163.367
R635 B.n182 B.n159 163.367
R636 B.n186 B.n159 163.367
R637 B.n187 B.n186 163.367
R638 B.n188 B.n187 163.367
R639 B.n188 B.n157 163.367
R640 B.n192 B.n157 163.367
R641 B.n193 B.n192 163.367
R642 B.n194 B.n193 163.367
R643 B.n194 B.n155 163.367
R644 B.n198 B.n155 163.367
R645 B.n199 B.n198 163.367
R646 B.n275 B.n129 59.5399
R647 B.n290 B.n289 59.5399
R648 B.n518 B.n47 59.5399
R649 B.n532 B.n41 59.5399
R650 B.n368 B.n367 35.4346
R651 B.n609 B.n14 35.4346
R652 B.n441 B.n72 35.4346
R653 B.n201 B.n154 35.4346
R654 B.n129 B.n128 21.9157
R655 B.n289 B.n288 21.9157
R656 B.n47 B.n46 21.9157
R657 B.n41 B.n40 21.9157
R658 B B.n645 18.0485
R659 B.n610 B.n609 10.6151
R660 B.n611 B.n610 10.6151
R661 B.n611 B.n12 10.6151
R662 B.n615 B.n12 10.6151
R663 B.n616 B.n615 10.6151
R664 B.n617 B.n616 10.6151
R665 B.n617 B.n10 10.6151
R666 B.n621 B.n10 10.6151
R667 B.n622 B.n621 10.6151
R668 B.n623 B.n622 10.6151
R669 B.n623 B.n8 10.6151
R670 B.n627 B.n8 10.6151
R671 B.n628 B.n627 10.6151
R672 B.n629 B.n628 10.6151
R673 B.n629 B.n6 10.6151
R674 B.n633 B.n6 10.6151
R675 B.n634 B.n633 10.6151
R676 B.n635 B.n634 10.6151
R677 B.n635 B.n4 10.6151
R678 B.n639 B.n4 10.6151
R679 B.n640 B.n639 10.6151
R680 B.n641 B.n640 10.6151
R681 B.n641 B.n0 10.6151
R682 B.n605 B.n14 10.6151
R683 B.n605 B.n604 10.6151
R684 B.n604 B.n603 10.6151
R685 B.n603 B.n16 10.6151
R686 B.n599 B.n16 10.6151
R687 B.n599 B.n598 10.6151
R688 B.n598 B.n597 10.6151
R689 B.n597 B.n18 10.6151
R690 B.n593 B.n18 10.6151
R691 B.n593 B.n592 10.6151
R692 B.n592 B.n591 10.6151
R693 B.n591 B.n20 10.6151
R694 B.n587 B.n20 10.6151
R695 B.n587 B.n586 10.6151
R696 B.n586 B.n585 10.6151
R697 B.n585 B.n22 10.6151
R698 B.n581 B.n22 10.6151
R699 B.n581 B.n580 10.6151
R700 B.n580 B.n579 10.6151
R701 B.n579 B.n24 10.6151
R702 B.n575 B.n24 10.6151
R703 B.n575 B.n574 10.6151
R704 B.n574 B.n573 10.6151
R705 B.n573 B.n26 10.6151
R706 B.n569 B.n26 10.6151
R707 B.n569 B.n568 10.6151
R708 B.n568 B.n567 10.6151
R709 B.n567 B.n28 10.6151
R710 B.n563 B.n28 10.6151
R711 B.n563 B.n562 10.6151
R712 B.n562 B.n561 10.6151
R713 B.n561 B.n30 10.6151
R714 B.n557 B.n30 10.6151
R715 B.n557 B.n556 10.6151
R716 B.n556 B.n555 10.6151
R717 B.n555 B.n32 10.6151
R718 B.n551 B.n32 10.6151
R719 B.n551 B.n550 10.6151
R720 B.n550 B.n549 10.6151
R721 B.n549 B.n34 10.6151
R722 B.n545 B.n34 10.6151
R723 B.n545 B.n544 10.6151
R724 B.n544 B.n543 10.6151
R725 B.n543 B.n36 10.6151
R726 B.n539 B.n36 10.6151
R727 B.n539 B.n538 10.6151
R728 B.n538 B.n537 10.6151
R729 B.n537 B.n38 10.6151
R730 B.n533 B.n38 10.6151
R731 B.n531 B.n530 10.6151
R732 B.n530 B.n42 10.6151
R733 B.n526 B.n42 10.6151
R734 B.n526 B.n525 10.6151
R735 B.n525 B.n524 10.6151
R736 B.n524 B.n44 10.6151
R737 B.n520 B.n44 10.6151
R738 B.n520 B.n519 10.6151
R739 B.n517 B.n48 10.6151
R740 B.n513 B.n48 10.6151
R741 B.n513 B.n512 10.6151
R742 B.n512 B.n511 10.6151
R743 B.n511 B.n50 10.6151
R744 B.n507 B.n50 10.6151
R745 B.n507 B.n506 10.6151
R746 B.n506 B.n505 10.6151
R747 B.n505 B.n52 10.6151
R748 B.n501 B.n52 10.6151
R749 B.n501 B.n500 10.6151
R750 B.n500 B.n499 10.6151
R751 B.n499 B.n54 10.6151
R752 B.n495 B.n54 10.6151
R753 B.n495 B.n494 10.6151
R754 B.n494 B.n493 10.6151
R755 B.n493 B.n56 10.6151
R756 B.n489 B.n56 10.6151
R757 B.n489 B.n488 10.6151
R758 B.n488 B.n487 10.6151
R759 B.n487 B.n58 10.6151
R760 B.n483 B.n58 10.6151
R761 B.n483 B.n482 10.6151
R762 B.n482 B.n481 10.6151
R763 B.n481 B.n60 10.6151
R764 B.n477 B.n60 10.6151
R765 B.n477 B.n476 10.6151
R766 B.n476 B.n475 10.6151
R767 B.n475 B.n62 10.6151
R768 B.n471 B.n62 10.6151
R769 B.n471 B.n470 10.6151
R770 B.n470 B.n469 10.6151
R771 B.n469 B.n64 10.6151
R772 B.n465 B.n64 10.6151
R773 B.n465 B.n464 10.6151
R774 B.n464 B.n463 10.6151
R775 B.n463 B.n66 10.6151
R776 B.n459 B.n66 10.6151
R777 B.n459 B.n458 10.6151
R778 B.n458 B.n457 10.6151
R779 B.n457 B.n68 10.6151
R780 B.n453 B.n68 10.6151
R781 B.n453 B.n452 10.6151
R782 B.n452 B.n451 10.6151
R783 B.n451 B.n70 10.6151
R784 B.n447 B.n70 10.6151
R785 B.n447 B.n446 10.6151
R786 B.n446 B.n445 10.6151
R787 B.n445 B.n72 10.6151
R788 B.n441 B.n440 10.6151
R789 B.n440 B.n439 10.6151
R790 B.n439 B.n74 10.6151
R791 B.n435 B.n74 10.6151
R792 B.n435 B.n434 10.6151
R793 B.n434 B.n433 10.6151
R794 B.n433 B.n76 10.6151
R795 B.n429 B.n76 10.6151
R796 B.n429 B.n428 10.6151
R797 B.n428 B.n427 10.6151
R798 B.n427 B.n78 10.6151
R799 B.n423 B.n78 10.6151
R800 B.n423 B.n422 10.6151
R801 B.n422 B.n421 10.6151
R802 B.n421 B.n80 10.6151
R803 B.n417 B.n80 10.6151
R804 B.n417 B.n416 10.6151
R805 B.n416 B.n415 10.6151
R806 B.n415 B.n82 10.6151
R807 B.n411 B.n82 10.6151
R808 B.n411 B.n410 10.6151
R809 B.n410 B.n409 10.6151
R810 B.n409 B.n84 10.6151
R811 B.n405 B.n84 10.6151
R812 B.n405 B.n404 10.6151
R813 B.n404 B.n403 10.6151
R814 B.n403 B.n86 10.6151
R815 B.n399 B.n86 10.6151
R816 B.n399 B.n398 10.6151
R817 B.n398 B.n397 10.6151
R818 B.n397 B.n88 10.6151
R819 B.n393 B.n88 10.6151
R820 B.n393 B.n392 10.6151
R821 B.n392 B.n391 10.6151
R822 B.n391 B.n90 10.6151
R823 B.n387 B.n90 10.6151
R824 B.n387 B.n386 10.6151
R825 B.n386 B.n385 10.6151
R826 B.n385 B.n92 10.6151
R827 B.n381 B.n92 10.6151
R828 B.n381 B.n380 10.6151
R829 B.n380 B.n379 10.6151
R830 B.n379 B.n94 10.6151
R831 B.n375 B.n94 10.6151
R832 B.n375 B.n374 10.6151
R833 B.n374 B.n373 10.6151
R834 B.n373 B.n96 10.6151
R835 B.n369 B.n96 10.6151
R836 B.n369 B.n368 10.6151
R837 B.n166 B.n1 10.6151
R838 B.n167 B.n166 10.6151
R839 B.n167 B.n164 10.6151
R840 B.n171 B.n164 10.6151
R841 B.n172 B.n171 10.6151
R842 B.n173 B.n172 10.6151
R843 B.n173 B.n162 10.6151
R844 B.n177 B.n162 10.6151
R845 B.n178 B.n177 10.6151
R846 B.n179 B.n178 10.6151
R847 B.n179 B.n160 10.6151
R848 B.n183 B.n160 10.6151
R849 B.n184 B.n183 10.6151
R850 B.n185 B.n184 10.6151
R851 B.n185 B.n158 10.6151
R852 B.n189 B.n158 10.6151
R853 B.n190 B.n189 10.6151
R854 B.n191 B.n190 10.6151
R855 B.n191 B.n156 10.6151
R856 B.n195 B.n156 10.6151
R857 B.n196 B.n195 10.6151
R858 B.n197 B.n196 10.6151
R859 B.n197 B.n154 10.6151
R860 B.n202 B.n201 10.6151
R861 B.n203 B.n202 10.6151
R862 B.n203 B.n152 10.6151
R863 B.n207 B.n152 10.6151
R864 B.n208 B.n207 10.6151
R865 B.n209 B.n208 10.6151
R866 B.n209 B.n150 10.6151
R867 B.n213 B.n150 10.6151
R868 B.n214 B.n213 10.6151
R869 B.n215 B.n214 10.6151
R870 B.n215 B.n148 10.6151
R871 B.n219 B.n148 10.6151
R872 B.n220 B.n219 10.6151
R873 B.n221 B.n220 10.6151
R874 B.n221 B.n146 10.6151
R875 B.n225 B.n146 10.6151
R876 B.n226 B.n225 10.6151
R877 B.n227 B.n226 10.6151
R878 B.n227 B.n144 10.6151
R879 B.n231 B.n144 10.6151
R880 B.n232 B.n231 10.6151
R881 B.n233 B.n232 10.6151
R882 B.n233 B.n142 10.6151
R883 B.n237 B.n142 10.6151
R884 B.n238 B.n237 10.6151
R885 B.n239 B.n238 10.6151
R886 B.n239 B.n140 10.6151
R887 B.n243 B.n140 10.6151
R888 B.n244 B.n243 10.6151
R889 B.n245 B.n244 10.6151
R890 B.n245 B.n138 10.6151
R891 B.n249 B.n138 10.6151
R892 B.n250 B.n249 10.6151
R893 B.n251 B.n250 10.6151
R894 B.n251 B.n136 10.6151
R895 B.n255 B.n136 10.6151
R896 B.n256 B.n255 10.6151
R897 B.n257 B.n256 10.6151
R898 B.n257 B.n134 10.6151
R899 B.n261 B.n134 10.6151
R900 B.n262 B.n261 10.6151
R901 B.n263 B.n262 10.6151
R902 B.n263 B.n132 10.6151
R903 B.n267 B.n132 10.6151
R904 B.n268 B.n267 10.6151
R905 B.n269 B.n268 10.6151
R906 B.n269 B.n130 10.6151
R907 B.n273 B.n130 10.6151
R908 B.n274 B.n273 10.6151
R909 B.n276 B.n126 10.6151
R910 B.n280 B.n126 10.6151
R911 B.n281 B.n280 10.6151
R912 B.n282 B.n281 10.6151
R913 B.n282 B.n124 10.6151
R914 B.n286 B.n124 10.6151
R915 B.n287 B.n286 10.6151
R916 B.n291 B.n287 10.6151
R917 B.n295 B.n122 10.6151
R918 B.n296 B.n295 10.6151
R919 B.n297 B.n296 10.6151
R920 B.n297 B.n120 10.6151
R921 B.n301 B.n120 10.6151
R922 B.n302 B.n301 10.6151
R923 B.n303 B.n302 10.6151
R924 B.n303 B.n118 10.6151
R925 B.n307 B.n118 10.6151
R926 B.n308 B.n307 10.6151
R927 B.n309 B.n308 10.6151
R928 B.n309 B.n116 10.6151
R929 B.n313 B.n116 10.6151
R930 B.n314 B.n313 10.6151
R931 B.n315 B.n314 10.6151
R932 B.n315 B.n114 10.6151
R933 B.n319 B.n114 10.6151
R934 B.n320 B.n319 10.6151
R935 B.n321 B.n320 10.6151
R936 B.n321 B.n112 10.6151
R937 B.n325 B.n112 10.6151
R938 B.n326 B.n325 10.6151
R939 B.n327 B.n326 10.6151
R940 B.n327 B.n110 10.6151
R941 B.n331 B.n110 10.6151
R942 B.n332 B.n331 10.6151
R943 B.n333 B.n332 10.6151
R944 B.n333 B.n108 10.6151
R945 B.n337 B.n108 10.6151
R946 B.n338 B.n337 10.6151
R947 B.n339 B.n338 10.6151
R948 B.n339 B.n106 10.6151
R949 B.n343 B.n106 10.6151
R950 B.n344 B.n343 10.6151
R951 B.n345 B.n344 10.6151
R952 B.n345 B.n104 10.6151
R953 B.n349 B.n104 10.6151
R954 B.n350 B.n349 10.6151
R955 B.n351 B.n350 10.6151
R956 B.n351 B.n102 10.6151
R957 B.n355 B.n102 10.6151
R958 B.n356 B.n355 10.6151
R959 B.n357 B.n356 10.6151
R960 B.n357 B.n100 10.6151
R961 B.n361 B.n100 10.6151
R962 B.n362 B.n361 10.6151
R963 B.n363 B.n362 10.6151
R964 B.n363 B.n98 10.6151
R965 B.n367 B.n98 10.6151
R966 B.n645 B.n0 8.11757
R967 B.n645 B.n1 8.11757
R968 B.n532 B.n531 6.5566
R969 B.n519 B.n518 6.5566
R970 B.n276 B.n275 6.5566
R971 B.n291 B.n290 6.5566
R972 B.n533 B.n532 4.05904
R973 B.n518 B.n517 4.05904
R974 B.n275 B.n274 4.05904
R975 B.n290 B.n122 4.05904
R976 VP.n4 VP.t6 514.955
R977 VP.n11 VP.t1 494.351
R978 VP.n1 VP.t7 494.351
R979 VP.n16 VP.t3 494.351
R980 VP.n18 VP.t0 494.351
R981 VP.n8 VP.t2 494.351
R982 VP.n6 VP.t4 494.351
R983 VP.n5 VP.t5 494.351
R984 VP.n19 VP.n18 161.3
R985 VP.n7 VP.n2 161.3
R986 VP.n9 VP.n8 161.3
R987 VP.n17 VP.n0 161.3
R988 VP.n13 VP.n12 161.3
R989 VP.n11 VP.n10 161.3
R990 VP.n6 VP.n3 80.6037
R991 VP.n16 VP.n15 80.6037
R992 VP.n14 VP.n1 80.6037
R993 VP.n16 VP.n1 48.2005
R994 VP.n6 VP.n5 48.2005
R995 VP.n10 VP.n9 44.5081
R996 VP.n12 VP.n1 41.6278
R997 VP.n17 VP.n16 41.6278
R998 VP.n7 VP.n6 41.6278
R999 VP.n4 VP.n3 31.6158
R1000 VP.n5 VP.n4 17.6494
R1001 VP.n12 VP.n11 6.57323
R1002 VP.n18 VP.n17 6.57323
R1003 VP.n8 VP.n7 6.57323
R1004 VP.n15 VP.n14 0.380177
R1005 VP.n3 VP.n2 0.285035
R1006 VP.n14 VP.n13 0.285035
R1007 VP.n15 VP.n0 0.285035
R1008 VP.n9 VP.n2 0.189894
R1009 VP.n13 VP.n10 0.189894
R1010 VP.n19 VP.n0 0.189894
R1011 VP VP.n19 0.0516364
R1012 VTAIL.n658 VTAIL.n582 756.745
R1013 VTAIL.n78 VTAIL.n2 756.745
R1014 VTAIL.n160 VTAIL.n84 756.745
R1015 VTAIL.n244 VTAIL.n168 756.745
R1016 VTAIL.n576 VTAIL.n500 756.745
R1017 VTAIL.n492 VTAIL.n416 756.745
R1018 VTAIL.n410 VTAIL.n334 756.745
R1019 VTAIL.n326 VTAIL.n250 756.745
R1020 VTAIL.n609 VTAIL.n608 585
R1021 VTAIL.n606 VTAIL.n605 585
R1022 VTAIL.n615 VTAIL.n614 585
R1023 VTAIL.n617 VTAIL.n616 585
R1024 VTAIL.n602 VTAIL.n601 585
R1025 VTAIL.n623 VTAIL.n622 585
R1026 VTAIL.n625 VTAIL.n624 585
R1027 VTAIL.n598 VTAIL.n597 585
R1028 VTAIL.n631 VTAIL.n630 585
R1029 VTAIL.n633 VTAIL.n632 585
R1030 VTAIL.n594 VTAIL.n593 585
R1031 VTAIL.n639 VTAIL.n638 585
R1032 VTAIL.n641 VTAIL.n640 585
R1033 VTAIL.n590 VTAIL.n589 585
R1034 VTAIL.n647 VTAIL.n646 585
R1035 VTAIL.n650 VTAIL.n649 585
R1036 VTAIL.n648 VTAIL.n586 585
R1037 VTAIL.n655 VTAIL.n585 585
R1038 VTAIL.n657 VTAIL.n656 585
R1039 VTAIL.n659 VTAIL.n658 585
R1040 VTAIL.n29 VTAIL.n28 585
R1041 VTAIL.n26 VTAIL.n25 585
R1042 VTAIL.n35 VTAIL.n34 585
R1043 VTAIL.n37 VTAIL.n36 585
R1044 VTAIL.n22 VTAIL.n21 585
R1045 VTAIL.n43 VTAIL.n42 585
R1046 VTAIL.n45 VTAIL.n44 585
R1047 VTAIL.n18 VTAIL.n17 585
R1048 VTAIL.n51 VTAIL.n50 585
R1049 VTAIL.n53 VTAIL.n52 585
R1050 VTAIL.n14 VTAIL.n13 585
R1051 VTAIL.n59 VTAIL.n58 585
R1052 VTAIL.n61 VTAIL.n60 585
R1053 VTAIL.n10 VTAIL.n9 585
R1054 VTAIL.n67 VTAIL.n66 585
R1055 VTAIL.n70 VTAIL.n69 585
R1056 VTAIL.n68 VTAIL.n6 585
R1057 VTAIL.n75 VTAIL.n5 585
R1058 VTAIL.n77 VTAIL.n76 585
R1059 VTAIL.n79 VTAIL.n78 585
R1060 VTAIL.n111 VTAIL.n110 585
R1061 VTAIL.n108 VTAIL.n107 585
R1062 VTAIL.n117 VTAIL.n116 585
R1063 VTAIL.n119 VTAIL.n118 585
R1064 VTAIL.n104 VTAIL.n103 585
R1065 VTAIL.n125 VTAIL.n124 585
R1066 VTAIL.n127 VTAIL.n126 585
R1067 VTAIL.n100 VTAIL.n99 585
R1068 VTAIL.n133 VTAIL.n132 585
R1069 VTAIL.n135 VTAIL.n134 585
R1070 VTAIL.n96 VTAIL.n95 585
R1071 VTAIL.n141 VTAIL.n140 585
R1072 VTAIL.n143 VTAIL.n142 585
R1073 VTAIL.n92 VTAIL.n91 585
R1074 VTAIL.n149 VTAIL.n148 585
R1075 VTAIL.n152 VTAIL.n151 585
R1076 VTAIL.n150 VTAIL.n88 585
R1077 VTAIL.n157 VTAIL.n87 585
R1078 VTAIL.n159 VTAIL.n158 585
R1079 VTAIL.n161 VTAIL.n160 585
R1080 VTAIL.n195 VTAIL.n194 585
R1081 VTAIL.n192 VTAIL.n191 585
R1082 VTAIL.n201 VTAIL.n200 585
R1083 VTAIL.n203 VTAIL.n202 585
R1084 VTAIL.n188 VTAIL.n187 585
R1085 VTAIL.n209 VTAIL.n208 585
R1086 VTAIL.n211 VTAIL.n210 585
R1087 VTAIL.n184 VTAIL.n183 585
R1088 VTAIL.n217 VTAIL.n216 585
R1089 VTAIL.n219 VTAIL.n218 585
R1090 VTAIL.n180 VTAIL.n179 585
R1091 VTAIL.n225 VTAIL.n224 585
R1092 VTAIL.n227 VTAIL.n226 585
R1093 VTAIL.n176 VTAIL.n175 585
R1094 VTAIL.n233 VTAIL.n232 585
R1095 VTAIL.n236 VTAIL.n235 585
R1096 VTAIL.n234 VTAIL.n172 585
R1097 VTAIL.n241 VTAIL.n171 585
R1098 VTAIL.n243 VTAIL.n242 585
R1099 VTAIL.n245 VTAIL.n244 585
R1100 VTAIL.n577 VTAIL.n576 585
R1101 VTAIL.n575 VTAIL.n574 585
R1102 VTAIL.n573 VTAIL.n503 585
R1103 VTAIL.n507 VTAIL.n504 585
R1104 VTAIL.n568 VTAIL.n567 585
R1105 VTAIL.n566 VTAIL.n565 585
R1106 VTAIL.n509 VTAIL.n508 585
R1107 VTAIL.n560 VTAIL.n559 585
R1108 VTAIL.n558 VTAIL.n557 585
R1109 VTAIL.n513 VTAIL.n512 585
R1110 VTAIL.n552 VTAIL.n551 585
R1111 VTAIL.n550 VTAIL.n549 585
R1112 VTAIL.n517 VTAIL.n516 585
R1113 VTAIL.n544 VTAIL.n543 585
R1114 VTAIL.n542 VTAIL.n541 585
R1115 VTAIL.n521 VTAIL.n520 585
R1116 VTAIL.n536 VTAIL.n535 585
R1117 VTAIL.n534 VTAIL.n533 585
R1118 VTAIL.n525 VTAIL.n524 585
R1119 VTAIL.n528 VTAIL.n527 585
R1120 VTAIL.n493 VTAIL.n492 585
R1121 VTAIL.n491 VTAIL.n490 585
R1122 VTAIL.n489 VTAIL.n419 585
R1123 VTAIL.n423 VTAIL.n420 585
R1124 VTAIL.n484 VTAIL.n483 585
R1125 VTAIL.n482 VTAIL.n481 585
R1126 VTAIL.n425 VTAIL.n424 585
R1127 VTAIL.n476 VTAIL.n475 585
R1128 VTAIL.n474 VTAIL.n473 585
R1129 VTAIL.n429 VTAIL.n428 585
R1130 VTAIL.n468 VTAIL.n467 585
R1131 VTAIL.n466 VTAIL.n465 585
R1132 VTAIL.n433 VTAIL.n432 585
R1133 VTAIL.n460 VTAIL.n459 585
R1134 VTAIL.n458 VTAIL.n457 585
R1135 VTAIL.n437 VTAIL.n436 585
R1136 VTAIL.n452 VTAIL.n451 585
R1137 VTAIL.n450 VTAIL.n449 585
R1138 VTAIL.n441 VTAIL.n440 585
R1139 VTAIL.n444 VTAIL.n443 585
R1140 VTAIL.n411 VTAIL.n410 585
R1141 VTAIL.n409 VTAIL.n408 585
R1142 VTAIL.n407 VTAIL.n337 585
R1143 VTAIL.n341 VTAIL.n338 585
R1144 VTAIL.n402 VTAIL.n401 585
R1145 VTAIL.n400 VTAIL.n399 585
R1146 VTAIL.n343 VTAIL.n342 585
R1147 VTAIL.n394 VTAIL.n393 585
R1148 VTAIL.n392 VTAIL.n391 585
R1149 VTAIL.n347 VTAIL.n346 585
R1150 VTAIL.n386 VTAIL.n385 585
R1151 VTAIL.n384 VTAIL.n383 585
R1152 VTAIL.n351 VTAIL.n350 585
R1153 VTAIL.n378 VTAIL.n377 585
R1154 VTAIL.n376 VTAIL.n375 585
R1155 VTAIL.n355 VTAIL.n354 585
R1156 VTAIL.n370 VTAIL.n369 585
R1157 VTAIL.n368 VTAIL.n367 585
R1158 VTAIL.n359 VTAIL.n358 585
R1159 VTAIL.n362 VTAIL.n361 585
R1160 VTAIL.n327 VTAIL.n326 585
R1161 VTAIL.n325 VTAIL.n324 585
R1162 VTAIL.n323 VTAIL.n253 585
R1163 VTAIL.n257 VTAIL.n254 585
R1164 VTAIL.n318 VTAIL.n317 585
R1165 VTAIL.n316 VTAIL.n315 585
R1166 VTAIL.n259 VTAIL.n258 585
R1167 VTAIL.n310 VTAIL.n309 585
R1168 VTAIL.n308 VTAIL.n307 585
R1169 VTAIL.n263 VTAIL.n262 585
R1170 VTAIL.n302 VTAIL.n301 585
R1171 VTAIL.n300 VTAIL.n299 585
R1172 VTAIL.n267 VTAIL.n266 585
R1173 VTAIL.n294 VTAIL.n293 585
R1174 VTAIL.n292 VTAIL.n291 585
R1175 VTAIL.n271 VTAIL.n270 585
R1176 VTAIL.n286 VTAIL.n285 585
R1177 VTAIL.n284 VTAIL.n283 585
R1178 VTAIL.n275 VTAIL.n274 585
R1179 VTAIL.n278 VTAIL.n277 585
R1180 VTAIL.t8 VTAIL.n526 327.466
R1181 VTAIL.t12 VTAIL.n442 327.466
R1182 VTAIL.t3 VTAIL.n360 327.466
R1183 VTAIL.t2 VTAIL.n276 327.466
R1184 VTAIL.t4 VTAIL.n607 327.466
R1185 VTAIL.t5 VTAIL.n27 327.466
R1186 VTAIL.t14 VTAIL.n109 327.466
R1187 VTAIL.t13 VTAIL.n193 327.466
R1188 VTAIL.n608 VTAIL.n605 171.744
R1189 VTAIL.n615 VTAIL.n605 171.744
R1190 VTAIL.n616 VTAIL.n615 171.744
R1191 VTAIL.n616 VTAIL.n601 171.744
R1192 VTAIL.n623 VTAIL.n601 171.744
R1193 VTAIL.n624 VTAIL.n623 171.744
R1194 VTAIL.n624 VTAIL.n597 171.744
R1195 VTAIL.n631 VTAIL.n597 171.744
R1196 VTAIL.n632 VTAIL.n631 171.744
R1197 VTAIL.n632 VTAIL.n593 171.744
R1198 VTAIL.n639 VTAIL.n593 171.744
R1199 VTAIL.n640 VTAIL.n639 171.744
R1200 VTAIL.n640 VTAIL.n589 171.744
R1201 VTAIL.n647 VTAIL.n589 171.744
R1202 VTAIL.n649 VTAIL.n647 171.744
R1203 VTAIL.n649 VTAIL.n648 171.744
R1204 VTAIL.n648 VTAIL.n585 171.744
R1205 VTAIL.n657 VTAIL.n585 171.744
R1206 VTAIL.n658 VTAIL.n657 171.744
R1207 VTAIL.n28 VTAIL.n25 171.744
R1208 VTAIL.n35 VTAIL.n25 171.744
R1209 VTAIL.n36 VTAIL.n35 171.744
R1210 VTAIL.n36 VTAIL.n21 171.744
R1211 VTAIL.n43 VTAIL.n21 171.744
R1212 VTAIL.n44 VTAIL.n43 171.744
R1213 VTAIL.n44 VTAIL.n17 171.744
R1214 VTAIL.n51 VTAIL.n17 171.744
R1215 VTAIL.n52 VTAIL.n51 171.744
R1216 VTAIL.n52 VTAIL.n13 171.744
R1217 VTAIL.n59 VTAIL.n13 171.744
R1218 VTAIL.n60 VTAIL.n59 171.744
R1219 VTAIL.n60 VTAIL.n9 171.744
R1220 VTAIL.n67 VTAIL.n9 171.744
R1221 VTAIL.n69 VTAIL.n67 171.744
R1222 VTAIL.n69 VTAIL.n68 171.744
R1223 VTAIL.n68 VTAIL.n5 171.744
R1224 VTAIL.n77 VTAIL.n5 171.744
R1225 VTAIL.n78 VTAIL.n77 171.744
R1226 VTAIL.n110 VTAIL.n107 171.744
R1227 VTAIL.n117 VTAIL.n107 171.744
R1228 VTAIL.n118 VTAIL.n117 171.744
R1229 VTAIL.n118 VTAIL.n103 171.744
R1230 VTAIL.n125 VTAIL.n103 171.744
R1231 VTAIL.n126 VTAIL.n125 171.744
R1232 VTAIL.n126 VTAIL.n99 171.744
R1233 VTAIL.n133 VTAIL.n99 171.744
R1234 VTAIL.n134 VTAIL.n133 171.744
R1235 VTAIL.n134 VTAIL.n95 171.744
R1236 VTAIL.n141 VTAIL.n95 171.744
R1237 VTAIL.n142 VTAIL.n141 171.744
R1238 VTAIL.n142 VTAIL.n91 171.744
R1239 VTAIL.n149 VTAIL.n91 171.744
R1240 VTAIL.n151 VTAIL.n149 171.744
R1241 VTAIL.n151 VTAIL.n150 171.744
R1242 VTAIL.n150 VTAIL.n87 171.744
R1243 VTAIL.n159 VTAIL.n87 171.744
R1244 VTAIL.n160 VTAIL.n159 171.744
R1245 VTAIL.n194 VTAIL.n191 171.744
R1246 VTAIL.n201 VTAIL.n191 171.744
R1247 VTAIL.n202 VTAIL.n201 171.744
R1248 VTAIL.n202 VTAIL.n187 171.744
R1249 VTAIL.n209 VTAIL.n187 171.744
R1250 VTAIL.n210 VTAIL.n209 171.744
R1251 VTAIL.n210 VTAIL.n183 171.744
R1252 VTAIL.n217 VTAIL.n183 171.744
R1253 VTAIL.n218 VTAIL.n217 171.744
R1254 VTAIL.n218 VTAIL.n179 171.744
R1255 VTAIL.n225 VTAIL.n179 171.744
R1256 VTAIL.n226 VTAIL.n225 171.744
R1257 VTAIL.n226 VTAIL.n175 171.744
R1258 VTAIL.n233 VTAIL.n175 171.744
R1259 VTAIL.n235 VTAIL.n233 171.744
R1260 VTAIL.n235 VTAIL.n234 171.744
R1261 VTAIL.n234 VTAIL.n171 171.744
R1262 VTAIL.n243 VTAIL.n171 171.744
R1263 VTAIL.n244 VTAIL.n243 171.744
R1264 VTAIL.n576 VTAIL.n575 171.744
R1265 VTAIL.n575 VTAIL.n503 171.744
R1266 VTAIL.n507 VTAIL.n503 171.744
R1267 VTAIL.n567 VTAIL.n507 171.744
R1268 VTAIL.n567 VTAIL.n566 171.744
R1269 VTAIL.n566 VTAIL.n508 171.744
R1270 VTAIL.n559 VTAIL.n508 171.744
R1271 VTAIL.n559 VTAIL.n558 171.744
R1272 VTAIL.n558 VTAIL.n512 171.744
R1273 VTAIL.n551 VTAIL.n512 171.744
R1274 VTAIL.n551 VTAIL.n550 171.744
R1275 VTAIL.n550 VTAIL.n516 171.744
R1276 VTAIL.n543 VTAIL.n516 171.744
R1277 VTAIL.n543 VTAIL.n542 171.744
R1278 VTAIL.n542 VTAIL.n520 171.744
R1279 VTAIL.n535 VTAIL.n520 171.744
R1280 VTAIL.n535 VTAIL.n534 171.744
R1281 VTAIL.n534 VTAIL.n524 171.744
R1282 VTAIL.n527 VTAIL.n524 171.744
R1283 VTAIL.n492 VTAIL.n491 171.744
R1284 VTAIL.n491 VTAIL.n419 171.744
R1285 VTAIL.n423 VTAIL.n419 171.744
R1286 VTAIL.n483 VTAIL.n423 171.744
R1287 VTAIL.n483 VTAIL.n482 171.744
R1288 VTAIL.n482 VTAIL.n424 171.744
R1289 VTAIL.n475 VTAIL.n424 171.744
R1290 VTAIL.n475 VTAIL.n474 171.744
R1291 VTAIL.n474 VTAIL.n428 171.744
R1292 VTAIL.n467 VTAIL.n428 171.744
R1293 VTAIL.n467 VTAIL.n466 171.744
R1294 VTAIL.n466 VTAIL.n432 171.744
R1295 VTAIL.n459 VTAIL.n432 171.744
R1296 VTAIL.n459 VTAIL.n458 171.744
R1297 VTAIL.n458 VTAIL.n436 171.744
R1298 VTAIL.n451 VTAIL.n436 171.744
R1299 VTAIL.n451 VTAIL.n450 171.744
R1300 VTAIL.n450 VTAIL.n440 171.744
R1301 VTAIL.n443 VTAIL.n440 171.744
R1302 VTAIL.n410 VTAIL.n409 171.744
R1303 VTAIL.n409 VTAIL.n337 171.744
R1304 VTAIL.n341 VTAIL.n337 171.744
R1305 VTAIL.n401 VTAIL.n341 171.744
R1306 VTAIL.n401 VTAIL.n400 171.744
R1307 VTAIL.n400 VTAIL.n342 171.744
R1308 VTAIL.n393 VTAIL.n342 171.744
R1309 VTAIL.n393 VTAIL.n392 171.744
R1310 VTAIL.n392 VTAIL.n346 171.744
R1311 VTAIL.n385 VTAIL.n346 171.744
R1312 VTAIL.n385 VTAIL.n384 171.744
R1313 VTAIL.n384 VTAIL.n350 171.744
R1314 VTAIL.n377 VTAIL.n350 171.744
R1315 VTAIL.n377 VTAIL.n376 171.744
R1316 VTAIL.n376 VTAIL.n354 171.744
R1317 VTAIL.n369 VTAIL.n354 171.744
R1318 VTAIL.n369 VTAIL.n368 171.744
R1319 VTAIL.n368 VTAIL.n358 171.744
R1320 VTAIL.n361 VTAIL.n358 171.744
R1321 VTAIL.n326 VTAIL.n325 171.744
R1322 VTAIL.n325 VTAIL.n253 171.744
R1323 VTAIL.n257 VTAIL.n253 171.744
R1324 VTAIL.n317 VTAIL.n257 171.744
R1325 VTAIL.n317 VTAIL.n316 171.744
R1326 VTAIL.n316 VTAIL.n258 171.744
R1327 VTAIL.n309 VTAIL.n258 171.744
R1328 VTAIL.n309 VTAIL.n308 171.744
R1329 VTAIL.n308 VTAIL.n262 171.744
R1330 VTAIL.n301 VTAIL.n262 171.744
R1331 VTAIL.n301 VTAIL.n300 171.744
R1332 VTAIL.n300 VTAIL.n266 171.744
R1333 VTAIL.n293 VTAIL.n266 171.744
R1334 VTAIL.n293 VTAIL.n292 171.744
R1335 VTAIL.n292 VTAIL.n270 171.744
R1336 VTAIL.n285 VTAIL.n270 171.744
R1337 VTAIL.n285 VTAIL.n284 171.744
R1338 VTAIL.n284 VTAIL.n274 171.744
R1339 VTAIL.n277 VTAIL.n274 171.744
R1340 VTAIL.n608 VTAIL.t4 85.8723
R1341 VTAIL.n28 VTAIL.t5 85.8723
R1342 VTAIL.n110 VTAIL.t14 85.8723
R1343 VTAIL.n194 VTAIL.t13 85.8723
R1344 VTAIL.n527 VTAIL.t8 85.8723
R1345 VTAIL.n443 VTAIL.t12 85.8723
R1346 VTAIL.n361 VTAIL.t3 85.8723
R1347 VTAIL.n277 VTAIL.t2 85.8723
R1348 VTAIL.n499 VTAIL.n498 56.609
R1349 VTAIL.n333 VTAIL.n332 56.609
R1350 VTAIL.n1 VTAIL.n0 56.6088
R1351 VTAIL.n167 VTAIL.n166 56.6088
R1352 VTAIL.n663 VTAIL.n662 34.7066
R1353 VTAIL.n83 VTAIL.n82 34.7066
R1354 VTAIL.n165 VTAIL.n164 34.7066
R1355 VTAIL.n249 VTAIL.n248 34.7066
R1356 VTAIL.n581 VTAIL.n580 34.7066
R1357 VTAIL.n497 VTAIL.n496 34.7066
R1358 VTAIL.n415 VTAIL.n414 34.7066
R1359 VTAIL.n331 VTAIL.n330 34.7066
R1360 VTAIL.n663 VTAIL.n581 26.0738
R1361 VTAIL.n331 VTAIL.n249 26.0738
R1362 VTAIL.n609 VTAIL.n607 16.3895
R1363 VTAIL.n29 VTAIL.n27 16.3895
R1364 VTAIL.n111 VTAIL.n109 16.3895
R1365 VTAIL.n195 VTAIL.n193 16.3895
R1366 VTAIL.n528 VTAIL.n526 16.3895
R1367 VTAIL.n444 VTAIL.n442 16.3895
R1368 VTAIL.n362 VTAIL.n360 16.3895
R1369 VTAIL.n278 VTAIL.n276 16.3895
R1370 VTAIL.n656 VTAIL.n655 13.1884
R1371 VTAIL.n76 VTAIL.n75 13.1884
R1372 VTAIL.n158 VTAIL.n157 13.1884
R1373 VTAIL.n242 VTAIL.n241 13.1884
R1374 VTAIL.n574 VTAIL.n573 13.1884
R1375 VTAIL.n490 VTAIL.n489 13.1884
R1376 VTAIL.n408 VTAIL.n407 13.1884
R1377 VTAIL.n324 VTAIL.n323 13.1884
R1378 VTAIL.n610 VTAIL.n606 12.8005
R1379 VTAIL.n654 VTAIL.n586 12.8005
R1380 VTAIL.n659 VTAIL.n584 12.8005
R1381 VTAIL.n30 VTAIL.n26 12.8005
R1382 VTAIL.n74 VTAIL.n6 12.8005
R1383 VTAIL.n79 VTAIL.n4 12.8005
R1384 VTAIL.n112 VTAIL.n108 12.8005
R1385 VTAIL.n156 VTAIL.n88 12.8005
R1386 VTAIL.n161 VTAIL.n86 12.8005
R1387 VTAIL.n196 VTAIL.n192 12.8005
R1388 VTAIL.n240 VTAIL.n172 12.8005
R1389 VTAIL.n245 VTAIL.n170 12.8005
R1390 VTAIL.n577 VTAIL.n502 12.8005
R1391 VTAIL.n572 VTAIL.n504 12.8005
R1392 VTAIL.n529 VTAIL.n525 12.8005
R1393 VTAIL.n493 VTAIL.n418 12.8005
R1394 VTAIL.n488 VTAIL.n420 12.8005
R1395 VTAIL.n445 VTAIL.n441 12.8005
R1396 VTAIL.n411 VTAIL.n336 12.8005
R1397 VTAIL.n406 VTAIL.n338 12.8005
R1398 VTAIL.n363 VTAIL.n359 12.8005
R1399 VTAIL.n327 VTAIL.n252 12.8005
R1400 VTAIL.n322 VTAIL.n254 12.8005
R1401 VTAIL.n279 VTAIL.n275 12.8005
R1402 VTAIL.n614 VTAIL.n613 12.0247
R1403 VTAIL.n651 VTAIL.n650 12.0247
R1404 VTAIL.n660 VTAIL.n582 12.0247
R1405 VTAIL.n34 VTAIL.n33 12.0247
R1406 VTAIL.n71 VTAIL.n70 12.0247
R1407 VTAIL.n80 VTAIL.n2 12.0247
R1408 VTAIL.n116 VTAIL.n115 12.0247
R1409 VTAIL.n153 VTAIL.n152 12.0247
R1410 VTAIL.n162 VTAIL.n84 12.0247
R1411 VTAIL.n200 VTAIL.n199 12.0247
R1412 VTAIL.n237 VTAIL.n236 12.0247
R1413 VTAIL.n246 VTAIL.n168 12.0247
R1414 VTAIL.n578 VTAIL.n500 12.0247
R1415 VTAIL.n569 VTAIL.n568 12.0247
R1416 VTAIL.n533 VTAIL.n532 12.0247
R1417 VTAIL.n494 VTAIL.n416 12.0247
R1418 VTAIL.n485 VTAIL.n484 12.0247
R1419 VTAIL.n449 VTAIL.n448 12.0247
R1420 VTAIL.n412 VTAIL.n334 12.0247
R1421 VTAIL.n403 VTAIL.n402 12.0247
R1422 VTAIL.n367 VTAIL.n366 12.0247
R1423 VTAIL.n328 VTAIL.n250 12.0247
R1424 VTAIL.n319 VTAIL.n318 12.0247
R1425 VTAIL.n283 VTAIL.n282 12.0247
R1426 VTAIL.n617 VTAIL.n604 11.249
R1427 VTAIL.n646 VTAIL.n588 11.249
R1428 VTAIL.n37 VTAIL.n24 11.249
R1429 VTAIL.n66 VTAIL.n8 11.249
R1430 VTAIL.n119 VTAIL.n106 11.249
R1431 VTAIL.n148 VTAIL.n90 11.249
R1432 VTAIL.n203 VTAIL.n190 11.249
R1433 VTAIL.n232 VTAIL.n174 11.249
R1434 VTAIL.n565 VTAIL.n506 11.249
R1435 VTAIL.n536 VTAIL.n523 11.249
R1436 VTAIL.n481 VTAIL.n422 11.249
R1437 VTAIL.n452 VTAIL.n439 11.249
R1438 VTAIL.n399 VTAIL.n340 11.249
R1439 VTAIL.n370 VTAIL.n357 11.249
R1440 VTAIL.n315 VTAIL.n256 11.249
R1441 VTAIL.n286 VTAIL.n273 11.249
R1442 VTAIL.n618 VTAIL.n602 10.4732
R1443 VTAIL.n645 VTAIL.n590 10.4732
R1444 VTAIL.n38 VTAIL.n22 10.4732
R1445 VTAIL.n65 VTAIL.n10 10.4732
R1446 VTAIL.n120 VTAIL.n104 10.4732
R1447 VTAIL.n147 VTAIL.n92 10.4732
R1448 VTAIL.n204 VTAIL.n188 10.4732
R1449 VTAIL.n231 VTAIL.n176 10.4732
R1450 VTAIL.n564 VTAIL.n509 10.4732
R1451 VTAIL.n537 VTAIL.n521 10.4732
R1452 VTAIL.n480 VTAIL.n425 10.4732
R1453 VTAIL.n453 VTAIL.n437 10.4732
R1454 VTAIL.n398 VTAIL.n343 10.4732
R1455 VTAIL.n371 VTAIL.n355 10.4732
R1456 VTAIL.n314 VTAIL.n259 10.4732
R1457 VTAIL.n287 VTAIL.n271 10.4732
R1458 VTAIL.n622 VTAIL.n621 9.69747
R1459 VTAIL.n642 VTAIL.n641 9.69747
R1460 VTAIL.n42 VTAIL.n41 9.69747
R1461 VTAIL.n62 VTAIL.n61 9.69747
R1462 VTAIL.n124 VTAIL.n123 9.69747
R1463 VTAIL.n144 VTAIL.n143 9.69747
R1464 VTAIL.n208 VTAIL.n207 9.69747
R1465 VTAIL.n228 VTAIL.n227 9.69747
R1466 VTAIL.n561 VTAIL.n560 9.69747
R1467 VTAIL.n541 VTAIL.n540 9.69747
R1468 VTAIL.n477 VTAIL.n476 9.69747
R1469 VTAIL.n457 VTAIL.n456 9.69747
R1470 VTAIL.n395 VTAIL.n394 9.69747
R1471 VTAIL.n375 VTAIL.n374 9.69747
R1472 VTAIL.n311 VTAIL.n310 9.69747
R1473 VTAIL.n291 VTAIL.n290 9.69747
R1474 VTAIL.n662 VTAIL.n661 9.45567
R1475 VTAIL.n82 VTAIL.n81 9.45567
R1476 VTAIL.n164 VTAIL.n163 9.45567
R1477 VTAIL.n248 VTAIL.n247 9.45567
R1478 VTAIL.n580 VTAIL.n579 9.45567
R1479 VTAIL.n496 VTAIL.n495 9.45567
R1480 VTAIL.n414 VTAIL.n413 9.45567
R1481 VTAIL.n330 VTAIL.n329 9.45567
R1482 VTAIL.n661 VTAIL.n660 9.3005
R1483 VTAIL.n584 VTAIL.n583 9.3005
R1484 VTAIL.n629 VTAIL.n628 9.3005
R1485 VTAIL.n627 VTAIL.n626 9.3005
R1486 VTAIL.n600 VTAIL.n599 9.3005
R1487 VTAIL.n621 VTAIL.n620 9.3005
R1488 VTAIL.n619 VTAIL.n618 9.3005
R1489 VTAIL.n604 VTAIL.n603 9.3005
R1490 VTAIL.n613 VTAIL.n612 9.3005
R1491 VTAIL.n611 VTAIL.n610 9.3005
R1492 VTAIL.n596 VTAIL.n595 9.3005
R1493 VTAIL.n635 VTAIL.n634 9.3005
R1494 VTAIL.n637 VTAIL.n636 9.3005
R1495 VTAIL.n592 VTAIL.n591 9.3005
R1496 VTAIL.n643 VTAIL.n642 9.3005
R1497 VTAIL.n645 VTAIL.n644 9.3005
R1498 VTAIL.n588 VTAIL.n587 9.3005
R1499 VTAIL.n652 VTAIL.n651 9.3005
R1500 VTAIL.n654 VTAIL.n653 9.3005
R1501 VTAIL.n81 VTAIL.n80 9.3005
R1502 VTAIL.n4 VTAIL.n3 9.3005
R1503 VTAIL.n49 VTAIL.n48 9.3005
R1504 VTAIL.n47 VTAIL.n46 9.3005
R1505 VTAIL.n20 VTAIL.n19 9.3005
R1506 VTAIL.n41 VTAIL.n40 9.3005
R1507 VTAIL.n39 VTAIL.n38 9.3005
R1508 VTAIL.n24 VTAIL.n23 9.3005
R1509 VTAIL.n33 VTAIL.n32 9.3005
R1510 VTAIL.n31 VTAIL.n30 9.3005
R1511 VTAIL.n16 VTAIL.n15 9.3005
R1512 VTAIL.n55 VTAIL.n54 9.3005
R1513 VTAIL.n57 VTAIL.n56 9.3005
R1514 VTAIL.n12 VTAIL.n11 9.3005
R1515 VTAIL.n63 VTAIL.n62 9.3005
R1516 VTAIL.n65 VTAIL.n64 9.3005
R1517 VTAIL.n8 VTAIL.n7 9.3005
R1518 VTAIL.n72 VTAIL.n71 9.3005
R1519 VTAIL.n74 VTAIL.n73 9.3005
R1520 VTAIL.n163 VTAIL.n162 9.3005
R1521 VTAIL.n86 VTAIL.n85 9.3005
R1522 VTAIL.n131 VTAIL.n130 9.3005
R1523 VTAIL.n129 VTAIL.n128 9.3005
R1524 VTAIL.n102 VTAIL.n101 9.3005
R1525 VTAIL.n123 VTAIL.n122 9.3005
R1526 VTAIL.n121 VTAIL.n120 9.3005
R1527 VTAIL.n106 VTAIL.n105 9.3005
R1528 VTAIL.n115 VTAIL.n114 9.3005
R1529 VTAIL.n113 VTAIL.n112 9.3005
R1530 VTAIL.n98 VTAIL.n97 9.3005
R1531 VTAIL.n137 VTAIL.n136 9.3005
R1532 VTAIL.n139 VTAIL.n138 9.3005
R1533 VTAIL.n94 VTAIL.n93 9.3005
R1534 VTAIL.n145 VTAIL.n144 9.3005
R1535 VTAIL.n147 VTAIL.n146 9.3005
R1536 VTAIL.n90 VTAIL.n89 9.3005
R1537 VTAIL.n154 VTAIL.n153 9.3005
R1538 VTAIL.n156 VTAIL.n155 9.3005
R1539 VTAIL.n247 VTAIL.n246 9.3005
R1540 VTAIL.n170 VTAIL.n169 9.3005
R1541 VTAIL.n215 VTAIL.n214 9.3005
R1542 VTAIL.n213 VTAIL.n212 9.3005
R1543 VTAIL.n186 VTAIL.n185 9.3005
R1544 VTAIL.n207 VTAIL.n206 9.3005
R1545 VTAIL.n205 VTAIL.n204 9.3005
R1546 VTAIL.n190 VTAIL.n189 9.3005
R1547 VTAIL.n199 VTAIL.n198 9.3005
R1548 VTAIL.n197 VTAIL.n196 9.3005
R1549 VTAIL.n182 VTAIL.n181 9.3005
R1550 VTAIL.n221 VTAIL.n220 9.3005
R1551 VTAIL.n223 VTAIL.n222 9.3005
R1552 VTAIL.n178 VTAIL.n177 9.3005
R1553 VTAIL.n229 VTAIL.n228 9.3005
R1554 VTAIL.n231 VTAIL.n230 9.3005
R1555 VTAIL.n174 VTAIL.n173 9.3005
R1556 VTAIL.n238 VTAIL.n237 9.3005
R1557 VTAIL.n240 VTAIL.n239 9.3005
R1558 VTAIL.n554 VTAIL.n553 9.3005
R1559 VTAIL.n556 VTAIL.n555 9.3005
R1560 VTAIL.n511 VTAIL.n510 9.3005
R1561 VTAIL.n562 VTAIL.n561 9.3005
R1562 VTAIL.n564 VTAIL.n563 9.3005
R1563 VTAIL.n506 VTAIL.n505 9.3005
R1564 VTAIL.n570 VTAIL.n569 9.3005
R1565 VTAIL.n572 VTAIL.n571 9.3005
R1566 VTAIL.n579 VTAIL.n578 9.3005
R1567 VTAIL.n502 VTAIL.n501 9.3005
R1568 VTAIL.n515 VTAIL.n514 9.3005
R1569 VTAIL.n548 VTAIL.n547 9.3005
R1570 VTAIL.n546 VTAIL.n545 9.3005
R1571 VTAIL.n519 VTAIL.n518 9.3005
R1572 VTAIL.n540 VTAIL.n539 9.3005
R1573 VTAIL.n538 VTAIL.n537 9.3005
R1574 VTAIL.n523 VTAIL.n522 9.3005
R1575 VTAIL.n532 VTAIL.n531 9.3005
R1576 VTAIL.n530 VTAIL.n529 9.3005
R1577 VTAIL.n470 VTAIL.n469 9.3005
R1578 VTAIL.n472 VTAIL.n471 9.3005
R1579 VTAIL.n427 VTAIL.n426 9.3005
R1580 VTAIL.n478 VTAIL.n477 9.3005
R1581 VTAIL.n480 VTAIL.n479 9.3005
R1582 VTAIL.n422 VTAIL.n421 9.3005
R1583 VTAIL.n486 VTAIL.n485 9.3005
R1584 VTAIL.n488 VTAIL.n487 9.3005
R1585 VTAIL.n495 VTAIL.n494 9.3005
R1586 VTAIL.n418 VTAIL.n417 9.3005
R1587 VTAIL.n431 VTAIL.n430 9.3005
R1588 VTAIL.n464 VTAIL.n463 9.3005
R1589 VTAIL.n462 VTAIL.n461 9.3005
R1590 VTAIL.n435 VTAIL.n434 9.3005
R1591 VTAIL.n456 VTAIL.n455 9.3005
R1592 VTAIL.n454 VTAIL.n453 9.3005
R1593 VTAIL.n439 VTAIL.n438 9.3005
R1594 VTAIL.n448 VTAIL.n447 9.3005
R1595 VTAIL.n446 VTAIL.n445 9.3005
R1596 VTAIL.n388 VTAIL.n387 9.3005
R1597 VTAIL.n390 VTAIL.n389 9.3005
R1598 VTAIL.n345 VTAIL.n344 9.3005
R1599 VTAIL.n396 VTAIL.n395 9.3005
R1600 VTAIL.n398 VTAIL.n397 9.3005
R1601 VTAIL.n340 VTAIL.n339 9.3005
R1602 VTAIL.n404 VTAIL.n403 9.3005
R1603 VTAIL.n406 VTAIL.n405 9.3005
R1604 VTAIL.n413 VTAIL.n412 9.3005
R1605 VTAIL.n336 VTAIL.n335 9.3005
R1606 VTAIL.n349 VTAIL.n348 9.3005
R1607 VTAIL.n382 VTAIL.n381 9.3005
R1608 VTAIL.n380 VTAIL.n379 9.3005
R1609 VTAIL.n353 VTAIL.n352 9.3005
R1610 VTAIL.n374 VTAIL.n373 9.3005
R1611 VTAIL.n372 VTAIL.n371 9.3005
R1612 VTAIL.n357 VTAIL.n356 9.3005
R1613 VTAIL.n366 VTAIL.n365 9.3005
R1614 VTAIL.n364 VTAIL.n363 9.3005
R1615 VTAIL.n304 VTAIL.n303 9.3005
R1616 VTAIL.n306 VTAIL.n305 9.3005
R1617 VTAIL.n261 VTAIL.n260 9.3005
R1618 VTAIL.n312 VTAIL.n311 9.3005
R1619 VTAIL.n314 VTAIL.n313 9.3005
R1620 VTAIL.n256 VTAIL.n255 9.3005
R1621 VTAIL.n320 VTAIL.n319 9.3005
R1622 VTAIL.n322 VTAIL.n321 9.3005
R1623 VTAIL.n329 VTAIL.n328 9.3005
R1624 VTAIL.n252 VTAIL.n251 9.3005
R1625 VTAIL.n265 VTAIL.n264 9.3005
R1626 VTAIL.n298 VTAIL.n297 9.3005
R1627 VTAIL.n296 VTAIL.n295 9.3005
R1628 VTAIL.n269 VTAIL.n268 9.3005
R1629 VTAIL.n290 VTAIL.n289 9.3005
R1630 VTAIL.n288 VTAIL.n287 9.3005
R1631 VTAIL.n273 VTAIL.n272 9.3005
R1632 VTAIL.n282 VTAIL.n281 9.3005
R1633 VTAIL.n280 VTAIL.n279 9.3005
R1634 VTAIL.n625 VTAIL.n600 8.92171
R1635 VTAIL.n638 VTAIL.n592 8.92171
R1636 VTAIL.n45 VTAIL.n20 8.92171
R1637 VTAIL.n58 VTAIL.n12 8.92171
R1638 VTAIL.n127 VTAIL.n102 8.92171
R1639 VTAIL.n140 VTAIL.n94 8.92171
R1640 VTAIL.n211 VTAIL.n186 8.92171
R1641 VTAIL.n224 VTAIL.n178 8.92171
R1642 VTAIL.n557 VTAIL.n511 8.92171
R1643 VTAIL.n544 VTAIL.n519 8.92171
R1644 VTAIL.n473 VTAIL.n427 8.92171
R1645 VTAIL.n460 VTAIL.n435 8.92171
R1646 VTAIL.n391 VTAIL.n345 8.92171
R1647 VTAIL.n378 VTAIL.n353 8.92171
R1648 VTAIL.n307 VTAIL.n261 8.92171
R1649 VTAIL.n294 VTAIL.n269 8.92171
R1650 VTAIL.n626 VTAIL.n598 8.14595
R1651 VTAIL.n637 VTAIL.n594 8.14595
R1652 VTAIL.n46 VTAIL.n18 8.14595
R1653 VTAIL.n57 VTAIL.n14 8.14595
R1654 VTAIL.n128 VTAIL.n100 8.14595
R1655 VTAIL.n139 VTAIL.n96 8.14595
R1656 VTAIL.n212 VTAIL.n184 8.14595
R1657 VTAIL.n223 VTAIL.n180 8.14595
R1658 VTAIL.n556 VTAIL.n513 8.14595
R1659 VTAIL.n545 VTAIL.n517 8.14595
R1660 VTAIL.n472 VTAIL.n429 8.14595
R1661 VTAIL.n461 VTAIL.n433 8.14595
R1662 VTAIL.n390 VTAIL.n347 8.14595
R1663 VTAIL.n379 VTAIL.n351 8.14595
R1664 VTAIL.n306 VTAIL.n263 8.14595
R1665 VTAIL.n295 VTAIL.n267 8.14595
R1666 VTAIL.n630 VTAIL.n629 7.3702
R1667 VTAIL.n634 VTAIL.n633 7.3702
R1668 VTAIL.n50 VTAIL.n49 7.3702
R1669 VTAIL.n54 VTAIL.n53 7.3702
R1670 VTAIL.n132 VTAIL.n131 7.3702
R1671 VTAIL.n136 VTAIL.n135 7.3702
R1672 VTAIL.n216 VTAIL.n215 7.3702
R1673 VTAIL.n220 VTAIL.n219 7.3702
R1674 VTAIL.n553 VTAIL.n552 7.3702
R1675 VTAIL.n549 VTAIL.n548 7.3702
R1676 VTAIL.n469 VTAIL.n468 7.3702
R1677 VTAIL.n465 VTAIL.n464 7.3702
R1678 VTAIL.n387 VTAIL.n386 7.3702
R1679 VTAIL.n383 VTAIL.n382 7.3702
R1680 VTAIL.n303 VTAIL.n302 7.3702
R1681 VTAIL.n299 VTAIL.n298 7.3702
R1682 VTAIL.n630 VTAIL.n596 6.59444
R1683 VTAIL.n633 VTAIL.n596 6.59444
R1684 VTAIL.n50 VTAIL.n16 6.59444
R1685 VTAIL.n53 VTAIL.n16 6.59444
R1686 VTAIL.n132 VTAIL.n98 6.59444
R1687 VTAIL.n135 VTAIL.n98 6.59444
R1688 VTAIL.n216 VTAIL.n182 6.59444
R1689 VTAIL.n219 VTAIL.n182 6.59444
R1690 VTAIL.n552 VTAIL.n515 6.59444
R1691 VTAIL.n549 VTAIL.n515 6.59444
R1692 VTAIL.n468 VTAIL.n431 6.59444
R1693 VTAIL.n465 VTAIL.n431 6.59444
R1694 VTAIL.n386 VTAIL.n349 6.59444
R1695 VTAIL.n383 VTAIL.n349 6.59444
R1696 VTAIL.n302 VTAIL.n265 6.59444
R1697 VTAIL.n299 VTAIL.n265 6.59444
R1698 VTAIL.n629 VTAIL.n598 5.81868
R1699 VTAIL.n634 VTAIL.n594 5.81868
R1700 VTAIL.n49 VTAIL.n18 5.81868
R1701 VTAIL.n54 VTAIL.n14 5.81868
R1702 VTAIL.n131 VTAIL.n100 5.81868
R1703 VTAIL.n136 VTAIL.n96 5.81868
R1704 VTAIL.n215 VTAIL.n184 5.81868
R1705 VTAIL.n220 VTAIL.n180 5.81868
R1706 VTAIL.n553 VTAIL.n513 5.81868
R1707 VTAIL.n548 VTAIL.n517 5.81868
R1708 VTAIL.n469 VTAIL.n429 5.81868
R1709 VTAIL.n464 VTAIL.n433 5.81868
R1710 VTAIL.n387 VTAIL.n347 5.81868
R1711 VTAIL.n382 VTAIL.n351 5.81868
R1712 VTAIL.n303 VTAIL.n263 5.81868
R1713 VTAIL.n298 VTAIL.n267 5.81868
R1714 VTAIL.n626 VTAIL.n625 5.04292
R1715 VTAIL.n638 VTAIL.n637 5.04292
R1716 VTAIL.n46 VTAIL.n45 5.04292
R1717 VTAIL.n58 VTAIL.n57 5.04292
R1718 VTAIL.n128 VTAIL.n127 5.04292
R1719 VTAIL.n140 VTAIL.n139 5.04292
R1720 VTAIL.n212 VTAIL.n211 5.04292
R1721 VTAIL.n224 VTAIL.n223 5.04292
R1722 VTAIL.n557 VTAIL.n556 5.04292
R1723 VTAIL.n545 VTAIL.n544 5.04292
R1724 VTAIL.n473 VTAIL.n472 5.04292
R1725 VTAIL.n461 VTAIL.n460 5.04292
R1726 VTAIL.n391 VTAIL.n390 5.04292
R1727 VTAIL.n379 VTAIL.n378 5.04292
R1728 VTAIL.n307 VTAIL.n306 5.04292
R1729 VTAIL.n295 VTAIL.n294 5.04292
R1730 VTAIL.n622 VTAIL.n600 4.26717
R1731 VTAIL.n641 VTAIL.n592 4.26717
R1732 VTAIL.n42 VTAIL.n20 4.26717
R1733 VTAIL.n61 VTAIL.n12 4.26717
R1734 VTAIL.n124 VTAIL.n102 4.26717
R1735 VTAIL.n143 VTAIL.n94 4.26717
R1736 VTAIL.n208 VTAIL.n186 4.26717
R1737 VTAIL.n227 VTAIL.n178 4.26717
R1738 VTAIL.n560 VTAIL.n511 4.26717
R1739 VTAIL.n541 VTAIL.n519 4.26717
R1740 VTAIL.n476 VTAIL.n427 4.26717
R1741 VTAIL.n457 VTAIL.n435 4.26717
R1742 VTAIL.n394 VTAIL.n345 4.26717
R1743 VTAIL.n375 VTAIL.n353 4.26717
R1744 VTAIL.n310 VTAIL.n261 4.26717
R1745 VTAIL.n291 VTAIL.n269 4.26717
R1746 VTAIL.n611 VTAIL.n607 3.70982
R1747 VTAIL.n31 VTAIL.n27 3.70982
R1748 VTAIL.n113 VTAIL.n109 3.70982
R1749 VTAIL.n197 VTAIL.n193 3.70982
R1750 VTAIL.n530 VTAIL.n526 3.70982
R1751 VTAIL.n446 VTAIL.n442 3.70982
R1752 VTAIL.n364 VTAIL.n360 3.70982
R1753 VTAIL.n280 VTAIL.n276 3.70982
R1754 VTAIL.n621 VTAIL.n602 3.49141
R1755 VTAIL.n642 VTAIL.n590 3.49141
R1756 VTAIL.n41 VTAIL.n22 3.49141
R1757 VTAIL.n62 VTAIL.n10 3.49141
R1758 VTAIL.n123 VTAIL.n104 3.49141
R1759 VTAIL.n144 VTAIL.n92 3.49141
R1760 VTAIL.n207 VTAIL.n188 3.49141
R1761 VTAIL.n228 VTAIL.n176 3.49141
R1762 VTAIL.n561 VTAIL.n509 3.49141
R1763 VTAIL.n540 VTAIL.n521 3.49141
R1764 VTAIL.n477 VTAIL.n425 3.49141
R1765 VTAIL.n456 VTAIL.n437 3.49141
R1766 VTAIL.n395 VTAIL.n343 3.49141
R1767 VTAIL.n374 VTAIL.n355 3.49141
R1768 VTAIL.n311 VTAIL.n259 3.49141
R1769 VTAIL.n290 VTAIL.n271 3.49141
R1770 VTAIL.n618 VTAIL.n617 2.71565
R1771 VTAIL.n646 VTAIL.n645 2.71565
R1772 VTAIL.n38 VTAIL.n37 2.71565
R1773 VTAIL.n66 VTAIL.n65 2.71565
R1774 VTAIL.n120 VTAIL.n119 2.71565
R1775 VTAIL.n148 VTAIL.n147 2.71565
R1776 VTAIL.n204 VTAIL.n203 2.71565
R1777 VTAIL.n232 VTAIL.n231 2.71565
R1778 VTAIL.n565 VTAIL.n564 2.71565
R1779 VTAIL.n537 VTAIL.n536 2.71565
R1780 VTAIL.n481 VTAIL.n480 2.71565
R1781 VTAIL.n453 VTAIL.n452 2.71565
R1782 VTAIL.n399 VTAIL.n398 2.71565
R1783 VTAIL.n371 VTAIL.n370 2.71565
R1784 VTAIL.n315 VTAIL.n314 2.71565
R1785 VTAIL.n287 VTAIL.n286 2.71565
R1786 VTAIL.n0 VTAIL.t0 2.20124
R1787 VTAIL.n0 VTAIL.t1 2.20124
R1788 VTAIL.n166 VTAIL.t15 2.20124
R1789 VTAIL.n166 VTAIL.t11 2.20124
R1790 VTAIL.n498 VTAIL.t10 2.20124
R1791 VTAIL.n498 VTAIL.t9 2.20124
R1792 VTAIL.n332 VTAIL.t6 2.20124
R1793 VTAIL.n332 VTAIL.t7 2.20124
R1794 VTAIL.n614 VTAIL.n604 1.93989
R1795 VTAIL.n650 VTAIL.n588 1.93989
R1796 VTAIL.n662 VTAIL.n582 1.93989
R1797 VTAIL.n34 VTAIL.n24 1.93989
R1798 VTAIL.n70 VTAIL.n8 1.93989
R1799 VTAIL.n82 VTAIL.n2 1.93989
R1800 VTAIL.n116 VTAIL.n106 1.93989
R1801 VTAIL.n152 VTAIL.n90 1.93989
R1802 VTAIL.n164 VTAIL.n84 1.93989
R1803 VTAIL.n200 VTAIL.n190 1.93989
R1804 VTAIL.n236 VTAIL.n174 1.93989
R1805 VTAIL.n248 VTAIL.n168 1.93989
R1806 VTAIL.n580 VTAIL.n500 1.93989
R1807 VTAIL.n568 VTAIL.n506 1.93989
R1808 VTAIL.n533 VTAIL.n523 1.93989
R1809 VTAIL.n496 VTAIL.n416 1.93989
R1810 VTAIL.n484 VTAIL.n422 1.93989
R1811 VTAIL.n449 VTAIL.n439 1.93989
R1812 VTAIL.n414 VTAIL.n334 1.93989
R1813 VTAIL.n402 VTAIL.n340 1.93989
R1814 VTAIL.n367 VTAIL.n357 1.93989
R1815 VTAIL.n330 VTAIL.n250 1.93989
R1816 VTAIL.n318 VTAIL.n256 1.93989
R1817 VTAIL.n283 VTAIL.n273 1.93989
R1818 VTAIL.n613 VTAIL.n606 1.16414
R1819 VTAIL.n651 VTAIL.n586 1.16414
R1820 VTAIL.n660 VTAIL.n659 1.16414
R1821 VTAIL.n33 VTAIL.n26 1.16414
R1822 VTAIL.n71 VTAIL.n6 1.16414
R1823 VTAIL.n80 VTAIL.n79 1.16414
R1824 VTAIL.n115 VTAIL.n108 1.16414
R1825 VTAIL.n153 VTAIL.n88 1.16414
R1826 VTAIL.n162 VTAIL.n161 1.16414
R1827 VTAIL.n199 VTAIL.n192 1.16414
R1828 VTAIL.n237 VTAIL.n172 1.16414
R1829 VTAIL.n246 VTAIL.n245 1.16414
R1830 VTAIL.n578 VTAIL.n577 1.16414
R1831 VTAIL.n569 VTAIL.n504 1.16414
R1832 VTAIL.n532 VTAIL.n525 1.16414
R1833 VTAIL.n494 VTAIL.n493 1.16414
R1834 VTAIL.n485 VTAIL.n420 1.16414
R1835 VTAIL.n448 VTAIL.n441 1.16414
R1836 VTAIL.n412 VTAIL.n411 1.16414
R1837 VTAIL.n403 VTAIL.n338 1.16414
R1838 VTAIL.n366 VTAIL.n359 1.16414
R1839 VTAIL.n328 VTAIL.n327 1.16414
R1840 VTAIL.n319 VTAIL.n254 1.16414
R1841 VTAIL.n282 VTAIL.n275 1.16414
R1842 VTAIL.n333 VTAIL.n331 0.974638
R1843 VTAIL.n415 VTAIL.n333 0.974638
R1844 VTAIL.n499 VTAIL.n497 0.974638
R1845 VTAIL.n581 VTAIL.n499 0.974638
R1846 VTAIL.n249 VTAIL.n167 0.974638
R1847 VTAIL.n167 VTAIL.n165 0.974638
R1848 VTAIL.n83 VTAIL.n1 0.974638
R1849 VTAIL VTAIL.n663 0.916448
R1850 VTAIL.n497 VTAIL.n415 0.470328
R1851 VTAIL.n165 VTAIL.n83 0.470328
R1852 VTAIL.n610 VTAIL.n609 0.388379
R1853 VTAIL.n655 VTAIL.n654 0.388379
R1854 VTAIL.n656 VTAIL.n584 0.388379
R1855 VTAIL.n30 VTAIL.n29 0.388379
R1856 VTAIL.n75 VTAIL.n74 0.388379
R1857 VTAIL.n76 VTAIL.n4 0.388379
R1858 VTAIL.n112 VTAIL.n111 0.388379
R1859 VTAIL.n157 VTAIL.n156 0.388379
R1860 VTAIL.n158 VTAIL.n86 0.388379
R1861 VTAIL.n196 VTAIL.n195 0.388379
R1862 VTAIL.n241 VTAIL.n240 0.388379
R1863 VTAIL.n242 VTAIL.n170 0.388379
R1864 VTAIL.n574 VTAIL.n502 0.388379
R1865 VTAIL.n573 VTAIL.n572 0.388379
R1866 VTAIL.n529 VTAIL.n528 0.388379
R1867 VTAIL.n490 VTAIL.n418 0.388379
R1868 VTAIL.n489 VTAIL.n488 0.388379
R1869 VTAIL.n445 VTAIL.n444 0.388379
R1870 VTAIL.n408 VTAIL.n336 0.388379
R1871 VTAIL.n407 VTAIL.n406 0.388379
R1872 VTAIL.n363 VTAIL.n362 0.388379
R1873 VTAIL.n324 VTAIL.n252 0.388379
R1874 VTAIL.n323 VTAIL.n322 0.388379
R1875 VTAIL.n279 VTAIL.n278 0.388379
R1876 VTAIL.n612 VTAIL.n611 0.155672
R1877 VTAIL.n612 VTAIL.n603 0.155672
R1878 VTAIL.n619 VTAIL.n603 0.155672
R1879 VTAIL.n620 VTAIL.n619 0.155672
R1880 VTAIL.n620 VTAIL.n599 0.155672
R1881 VTAIL.n627 VTAIL.n599 0.155672
R1882 VTAIL.n628 VTAIL.n627 0.155672
R1883 VTAIL.n628 VTAIL.n595 0.155672
R1884 VTAIL.n635 VTAIL.n595 0.155672
R1885 VTAIL.n636 VTAIL.n635 0.155672
R1886 VTAIL.n636 VTAIL.n591 0.155672
R1887 VTAIL.n643 VTAIL.n591 0.155672
R1888 VTAIL.n644 VTAIL.n643 0.155672
R1889 VTAIL.n644 VTAIL.n587 0.155672
R1890 VTAIL.n652 VTAIL.n587 0.155672
R1891 VTAIL.n653 VTAIL.n652 0.155672
R1892 VTAIL.n653 VTAIL.n583 0.155672
R1893 VTAIL.n661 VTAIL.n583 0.155672
R1894 VTAIL.n32 VTAIL.n31 0.155672
R1895 VTAIL.n32 VTAIL.n23 0.155672
R1896 VTAIL.n39 VTAIL.n23 0.155672
R1897 VTAIL.n40 VTAIL.n39 0.155672
R1898 VTAIL.n40 VTAIL.n19 0.155672
R1899 VTAIL.n47 VTAIL.n19 0.155672
R1900 VTAIL.n48 VTAIL.n47 0.155672
R1901 VTAIL.n48 VTAIL.n15 0.155672
R1902 VTAIL.n55 VTAIL.n15 0.155672
R1903 VTAIL.n56 VTAIL.n55 0.155672
R1904 VTAIL.n56 VTAIL.n11 0.155672
R1905 VTAIL.n63 VTAIL.n11 0.155672
R1906 VTAIL.n64 VTAIL.n63 0.155672
R1907 VTAIL.n64 VTAIL.n7 0.155672
R1908 VTAIL.n72 VTAIL.n7 0.155672
R1909 VTAIL.n73 VTAIL.n72 0.155672
R1910 VTAIL.n73 VTAIL.n3 0.155672
R1911 VTAIL.n81 VTAIL.n3 0.155672
R1912 VTAIL.n114 VTAIL.n113 0.155672
R1913 VTAIL.n114 VTAIL.n105 0.155672
R1914 VTAIL.n121 VTAIL.n105 0.155672
R1915 VTAIL.n122 VTAIL.n121 0.155672
R1916 VTAIL.n122 VTAIL.n101 0.155672
R1917 VTAIL.n129 VTAIL.n101 0.155672
R1918 VTAIL.n130 VTAIL.n129 0.155672
R1919 VTAIL.n130 VTAIL.n97 0.155672
R1920 VTAIL.n137 VTAIL.n97 0.155672
R1921 VTAIL.n138 VTAIL.n137 0.155672
R1922 VTAIL.n138 VTAIL.n93 0.155672
R1923 VTAIL.n145 VTAIL.n93 0.155672
R1924 VTAIL.n146 VTAIL.n145 0.155672
R1925 VTAIL.n146 VTAIL.n89 0.155672
R1926 VTAIL.n154 VTAIL.n89 0.155672
R1927 VTAIL.n155 VTAIL.n154 0.155672
R1928 VTAIL.n155 VTAIL.n85 0.155672
R1929 VTAIL.n163 VTAIL.n85 0.155672
R1930 VTAIL.n198 VTAIL.n197 0.155672
R1931 VTAIL.n198 VTAIL.n189 0.155672
R1932 VTAIL.n205 VTAIL.n189 0.155672
R1933 VTAIL.n206 VTAIL.n205 0.155672
R1934 VTAIL.n206 VTAIL.n185 0.155672
R1935 VTAIL.n213 VTAIL.n185 0.155672
R1936 VTAIL.n214 VTAIL.n213 0.155672
R1937 VTAIL.n214 VTAIL.n181 0.155672
R1938 VTAIL.n221 VTAIL.n181 0.155672
R1939 VTAIL.n222 VTAIL.n221 0.155672
R1940 VTAIL.n222 VTAIL.n177 0.155672
R1941 VTAIL.n229 VTAIL.n177 0.155672
R1942 VTAIL.n230 VTAIL.n229 0.155672
R1943 VTAIL.n230 VTAIL.n173 0.155672
R1944 VTAIL.n238 VTAIL.n173 0.155672
R1945 VTAIL.n239 VTAIL.n238 0.155672
R1946 VTAIL.n239 VTAIL.n169 0.155672
R1947 VTAIL.n247 VTAIL.n169 0.155672
R1948 VTAIL.n579 VTAIL.n501 0.155672
R1949 VTAIL.n571 VTAIL.n501 0.155672
R1950 VTAIL.n571 VTAIL.n570 0.155672
R1951 VTAIL.n570 VTAIL.n505 0.155672
R1952 VTAIL.n563 VTAIL.n505 0.155672
R1953 VTAIL.n563 VTAIL.n562 0.155672
R1954 VTAIL.n562 VTAIL.n510 0.155672
R1955 VTAIL.n555 VTAIL.n510 0.155672
R1956 VTAIL.n555 VTAIL.n554 0.155672
R1957 VTAIL.n554 VTAIL.n514 0.155672
R1958 VTAIL.n547 VTAIL.n514 0.155672
R1959 VTAIL.n547 VTAIL.n546 0.155672
R1960 VTAIL.n546 VTAIL.n518 0.155672
R1961 VTAIL.n539 VTAIL.n518 0.155672
R1962 VTAIL.n539 VTAIL.n538 0.155672
R1963 VTAIL.n538 VTAIL.n522 0.155672
R1964 VTAIL.n531 VTAIL.n522 0.155672
R1965 VTAIL.n531 VTAIL.n530 0.155672
R1966 VTAIL.n495 VTAIL.n417 0.155672
R1967 VTAIL.n487 VTAIL.n417 0.155672
R1968 VTAIL.n487 VTAIL.n486 0.155672
R1969 VTAIL.n486 VTAIL.n421 0.155672
R1970 VTAIL.n479 VTAIL.n421 0.155672
R1971 VTAIL.n479 VTAIL.n478 0.155672
R1972 VTAIL.n478 VTAIL.n426 0.155672
R1973 VTAIL.n471 VTAIL.n426 0.155672
R1974 VTAIL.n471 VTAIL.n470 0.155672
R1975 VTAIL.n470 VTAIL.n430 0.155672
R1976 VTAIL.n463 VTAIL.n430 0.155672
R1977 VTAIL.n463 VTAIL.n462 0.155672
R1978 VTAIL.n462 VTAIL.n434 0.155672
R1979 VTAIL.n455 VTAIL.n434 0.155672
R1980 VTAIL.n455 VTAIL.n454 0.155672
R1981 VTAIL.n454 VTAIL.n438 0.155672
R1982 VTAIL.n447 VTAIL.n438 0.155672
R1983 VTAIL.n447 VTAIL.n446 0.155672
R1984 VTAIL.n413 VTAIL.n335 0.155672
R1985 VTAIL.n405 VTAIL.n335 0.155672
R1986 VTAIL.n405 VTAIL.n404 0.155672
R1987 VTAIL.n404 VTAIL.n339 0.155672
R1988 VTAIL.n397 VTAIL.n339 0.155672
R1989 VTAIL.n397 VTAIL.n396 0.155672
R1990 VTAIL.n396 VTAIL.n344 0.155672
R1991 VTAIL.n389 VTAIL.n344 0.155672
R1992 VTAIL.n389 VTAIL.n388 0.155672
R1993 VTAIL.n388 VTAIL.n348 0.155672
R1994 VTAIL.n381 VTAIL.n348 0.155672
R1995 VTAIL.n381 VTAIL.n380 0.155672
R1996 VTAIL.n380 VTAIL.n352 0.155672
R1997 VTAIL.n373 VTAIL.n352 0.155672
R1998 VTAIL.n373 VTAIL.n372 0.155672
R1999 VTAIL.n372 VTAIL.n356 0.155672
R2000 VTAIL.n365 VTAIL.n356 0.155672
R2001 VTAIL.n365 VTAIL.n364 0.155672
R2002 VTAIL.n329 VTAIL.n251 0.155672
R2003 VTAIL.n321 VTAIL.n251 0.155672
R2004 VTAIL.n321 VTAIL.n320 0.155672
R2005 VTAIL.n320 VTAIL.n255 0.155672
R2006 VTAIL.n313 VTAIL.n255 0.155672
R2007 VTAIL.n313 VTAIL.n312 0.155672
R2008 VTAIL.n312 VTAIL.n260 0.155672
R2009 VTAIL.n305 VTAIL.n260 0.155672
R2010 VTAIL.n305 VTAIL.n304 0.155672
R2011 VTAIL.n304 VTAIL.n264 0.155672
R2012 VTAIL.n297 VTAIL.n264 0.155672
R2013 VTAIL.n297 VTAIL.n296 0.155672
R2014 VTAIL.n296 VTAIL.n268 0.155672
R2015 VTAIL.n289 VTAIL.n268 0.155672
R2016 VTAIL.n289 VTAIL.n288 0.155672
R2017 VTAIL.n288 VTAIL.n272 0.155672
R2018 VTAIL.n281 VTAIL.n272 0.155672
R2019 VTAIL.n281 VTAIL.n280 0.155672
R2020 VTAIL VTAIL.n1 0.0586897
R2021 VDD1 VDD1.n0 73.833
R2022 VDD1.n3 VDD1.n2 73.7193
R2023 VDD1.n3 VDD1.n1 73.7193
R2024 VDD1.n5 VDD1.n4 73.2876
R2025 VDD1.n5 VDD1.n3 41.4147
R2026 VDD1.n4 VDD1.t3 2.20124
R2027 VDD1.n4 VDD1.t5 2.20124
R2028 VDD1.n0 VDD1.t1 2.20124
R2029 VDD1.n0 VDD1.t2 2.20124
R2030 VDD1.n2 VDD1.t4 2.20124
R2031 VDD1.n2 VDD1.t7 2.20124
R2032 VDD1.n1 VDD1.t6 2.20124
R2033 VDD1.n1 VDD1.t0 2.20124
R2034 VDD1 VDD1.n5 0.429379
R2035 VN.n2 VN.t0 514.955
R2036 VN.n10 VN.t3 514.955
R2037 VN.n1 VN.t6 494.351
R2038 VN.n4 VN.t7 494.351
R2039 VN.n6 VN.t5 494.351
R2040 VN.n9 VN.t2 494.351
R2041 VN.n12 VN.t1 494.351
R2042 VN.n14 VN.t4 494.351
R2043 VN.n7 VN.n6 161.3
R2044 VN.n15 VN.n14 161.3
R2045 VN.n13 VN.n8 161.3
R2046 VN.n5 VN.n0 161.3
R2047 VN.n12 VN.n11 80.6037
R2048 VN.n4 VN.n3 80.6037
R2049 VN.n4 VN.n1 48.2005
R2050 VN.n12 VN.n9 48.2005
R2051 VN VN.n15 44.8888
R2052 VN.n5 VN.n4 41.6278
R2053 VN.n13 VN.n12 41.6278
R2054 VN.n11 VN.n10 31.6158
R2055 VN.n3 VN.n2 31.6158
R2056 VN.n2 VN.n1 17.6494
R2057 VN.n10 VN.n9 17.6494
R2058 VN.n6 VN.n5 6.57323
R2059 VN.n14 VN.n13 6.57323
R2060 VN.n11 VN.n8 0.285035
R2061 VN.n3 VN.n0 0.285035
R2062 VN.n15 VN.n8 0.189894
R2063 VN.n7 VN.n0 0.189894
R2064 VN VN.n7 0.0516364
R2065 VDD2.n2 VDD2.n1 73.7193
R2066 VDD2.n2 VDD2.n0 73.7193
R2067 VDD2 VDD2.n5 73.7165
R2068 VDD2.n4 VDD2.n3 73.2878
R2069 VDD2.n4 VDD2.n2 40.8317
R2070 VDD2.n5 VDD2.t5 2.20124
R2071 VDD2.n5 VDD2.t4 2.20124
R2072 VDD2.n3 VDD2.t3 2.20124
R2073 VDD2.n3 VDD2.t6 2.20124
R2074 VDD2.n1 VDD2.t0 2.20124
R2075 VDD2.n1 VDD2.t2 2.20124
R2076 VDD2.n0 VDD2.t7 2.20124
R2077 VDD2.n0 VDD2.t1 2.20124
R2078 VDD2 VDD2.n4 0.545759
C0 VP w_n2100_n3922# 4.09581f
C1 VDD1 w_n2100_n3922# 1.4113f
C2 VDD2 w_n2100_n3922# 1.45029f
C3 VTAIL w_n2100_n3922# 4.88253f
C4 VP B 1.27598f
C5 VDD1 B 1.17519f
C6 w_n2100_n3922# VN 3.82849f
C7 VDD2 B 1.21494f
C8 VTAIL B 4.67953f
C9 B VN 0.83746f
C10 VDD1 VP 7.33705f
C11 VDD2 VP 0.328001f
C12 VTAIL VP 6.8614f
C13 VDD1 VDD2 0.874934f
C14 VDD1 VTAIL 12.3577f
C15 B w_n2100_n3922# 8.13756f
C16 VDD2 VTAIL 12.4001f
C17 VP VN 5.977f
C18 VDD1 VN 0.148343f
C19 VDD2 VN 7.15787f
C20 VTAIL VN 6.8473f
C21 VDD2 VSUBS 1.4186f
C22 VDD1 VSUBS 1.741089f
C23 VTAIL VSUBS 1.060532f
C24 VN VSUBS 4.93785f
C25 VP VSUBS 1.844314f
C26 B VSUBS 3.232256f
C27 w_n2100_n3922# VSUBS 0.101027p
C28 VDD2.t7 VSUBS 0.313832f
C29 VDD2.t1 VSUBS 0.313832f
C30 VDD2.n0 VSUBS 2.55458f
C31 VDD2.t0 VSUBS 0.313832f
C32 VDD2.t2 VSUBS 0.313832f
C33 VDD2.n1 VSUBS 2.55458f
C34 VDD2.n2 VSUBS 3.14509f
C35 VDD2.t3 VSUBS 0.313832f
C36 VDD2.t6 VSUBS 0.313832f
C37 VDD2.n3 VSUBS 2.55086f
C38 VDD2.n4 VSUBS 3.01286f
C39 VDD2.t5 VSUBS 0.313832f
C40 VDD2.t4 VSUBS 0.313832f
C41 VDD2.n5 VSUBS 2.55455f
C42 VN.n0 VSUBS 0.066049f
C43 VN.t6 VSUBS 1.66276f
C44 VN.n1 VSUBS 0.65334f
C45 VN.t0 VSUBS 1.6885f
C46 VN.n2 VSUBS 0.62161f
C47 VN.n3 VSUBS 0.283297f
C48 VN.t7 VSUBS 1.66276f
C49 VN.n4 VSUBS 0.652534f
C50 VN.n5 VSUBS 0.011232f
C51 VN.t5 VSUBS 1.66276f
C52 VN.n6 VSUBS 0.633977f
C53 VN.n7 VSUBS 0.038359f
C54 VN.n8 VSUBS 0.066049f
C55 VN.t2 VSUBS 1.66276f
C56 VN.n9 VSUBS 0.65334f
C57 VN.t1 VSUBS 1.66276f
C58 VN.t3 VSUBS 1.6885f
C59 VN.n10 VSUBS 0.62161f
C60 VN.n11 VSUBS 0.283297f
C61 VN.n12 VSUBS 0.652534f
C62 VN.n13 VSUBS 0.011232f
C63 VN.t4 VSUBS 1.66276f
C64 VN.n14 VSUBS 0.633977f
C65 VN.n15 VSUBS 2.27878f
C66 VDD1.t1 VSUBS 0.313843f
C67 VDD1.t2 VSUBS 0.313843f
C68 VDD1.n0 VSUBS 2.55572f
C69 VDD1.t6 VSUBS 0.313843f
C70 VDD1.t0 VSUBS 0.313843f
C71 VDD1.n1 VSUBS 2.55467f
C72 VDD1.t4 VSUBS 0.313843f
C73 VDD1.t7 VSUBS 0.313843f
C74 VDD1.n2 VSUBS 2.55467f
C75 VDD1.n3 VSUBS 3.20233f
C76 VDD1.t3 VSUBS 0.313843f
C77 VDD1.t5 VSUBS 0.313843f
C78 VDD1.n4 VSUBS 2.55094f
C79 VDD1.n5 VSUBS 3.04508f
C80 VTAIL.t0 VSUBS 0.283221f
C81 VTAIL.t1 VSUBS 0.283221f
C82 VTAIL.n0 VSUBS 2.16945f
C83 VTAIL.n1 VSUBS 0.634916f
C84 VTAIL.n2 VSUBS 0.025841f
C85 VTAIL.n3 VSUBS 0.024266f
C86 VTAIL.n4 VSUBS 0.013039f
C87 VTAIL.n5 VSUBS 0.03082f
C88 VTAIL.n6 VSUBS 0.013806f
C89 VTAIL.n7 VSUBS 0.024266f
C90 VTAIL.n8 VSUBS 0.013039f
C91 VTAIL.n9 VSUBS 0.03082f
C92 VTAIL.n10 VSUBS 0.013806f
C93 VTAIL.n11 VSUBS 0.024266f
C94 VTAIL.n12 VSUBS 0.013039f
C95 VTAIL.n13 VSUBS 0.03082f
C96 VTAIL.n14 VSUBS 0.013806f
C97 VTAIL.n15 VSUBS 0.024266f
C98 VTAIL.n16 VSUBS 0.013039f
C99 VTAIL.n17 VSUBS 0.03082f
C100 VTAIL.n18 VSUBS 0.013806f
C101 VTAIL.n19 VSUBS 0.024266f
C102 VTAIL.n20 VSUBS 0.013039f
C103 VTAIL.n21 VSUBS 0.03082f
C104 VTAIL.n22 VSUBS 0.013806f
C105 VTAIL.n23 VSUBS 0.024266f
C106 VTAIL.n24 VSUBS 0.013039f
C107 VTAIL.n25 VSUBS 0.03082f
C108 VTAIL.n26 VSUBS 0.013806f
C109 VTAIL.n27 VSUBS 0.169406f
C110 VTAIL.t5 VSUBS 0.065966f
C111 VTAIL.n28 VSUBS 0.023115f
C112 VTAIL.n29 VSUBS 0.019606f
C113 VTAIL.n30 VSUBS 0.013039f
C114 VTAIL.n31 VSUBS 1.52407f
C115 VTAIL.n32 VSUBS 0.024266f
C116 VTAIL.n33 VSUBS 0.013039f
C117 VTAIL.n34 VSUBS 0.013806f
C118 VTAIL.n35 VSUBS 0.03082f
C119 VTAIL.n36 VSUBS 0.03082f
C120 VTAIL.n37 VSUBS 0.013806f
C121 VTAIL.n38 VSUBS 0.013039f
C122 VTAIL.n39 VSUBS 0.024266f
C123 VTAIL.n40 VSUBS 0.024266f
C124 VTAIL.n41 VSUBS 0.013039f
C125 VTAIL.n42 VSUBS 0.013806f
C126 VTAIL.n43 VSUBS 0.03082f
C127 VTAIL.n44 VSUBS 0.03082f
C128 VTAIL.n45 VSUBS 0.013806f
C129 VTAIL.n46 VSUBS 0.013039f
C130 VTAIL.n47 VSUBS 0.024266f
C131 VTAIL.n48 VSUBS 0.024266f
C132 VTAIL.n49 VSUBS 0.013039f
C133 VTAIL.n50 VSUBS 0.013806f
C134 VTAIL.n51 VSUBS 0.03082f
C135 VTAIL.n52 VSUBS 0.03082f
C136 VTAIL.n53 VSUBS 0.013806f
C137 VTAIL.n54 VSUBS 0.013039f
C138 VTAIL.n55 VSUBS 0.024266f
C139 VTAIL.n56 VSUBS 0.024266f
C140 VTAIL.n57 VSUBS 0.013039f
C141 VTAIL.n58 VSUBS 0.013806f
C142 VTAIL.n59 VSUBS 0.03082f
C143 VTAIL.n60 VSUBS 0.03082f
C144 VTAIL.n61 VSUBS 0.013806f
C145 VTAIL.n62 VSUBS 0.013039f
C146 VTAIL.n63 VSUBS 0.024266f
C147 VTAIL.n64 VSUBS 0.024266f
C148 VTAIL.n65 VSUBS 0.013039f
C149 VTAIL.n66 VSUBS 0.013806f
C150 VTAIL.n67 VSUBS 0.03082f
C151 VTAIL.n68 VSUBS 0.03082f
C152 VTAIL.n69 VSUBS 0.03082f
C153 VTAIL.n70 VSUBS 0.013806f
C154 VTAIL.n71 VSUBS 0.013039f
C155 VTAIL.n72 VSUBS 0.024266f
C156 VTAIL.n73 VSUBS 0.024266f
C157 VTAIL.n74 VSUBS 0.013039f
C158 VTAIL.n75 VSUBS 0.013423f
C159 VTAIL.n76 VSUBS 0.013423f
C160 VTAIL.n77 VSUBS 0.03082f
C161 VTAIL.n78 VSUBS 0.071814f
C162 VTAIL.n79 VSUBS 0.013806f
C163 VTAIL.n80 VSUBS 0.013039f
C164 VTAIL.n81 VSUBS 0.060398f
C165 VTAIL.n82 VSUBS 0.036118f
C166 VTAIL.n83 VSUBS 0.136064f
C167 VTAIL.n84 VSUBS 0.025841f
C168 VTAIL.n85 VSUBS 0.024266f
C169 VTAIL.n86 VSUBS 0.013039f
C170 VTAIL.n87 VSUBS 0.03082f
C171 VTAIL.n88 VSUBS 0.013806f
C172 VTAIL.n89 VSUBS 0.024266f
C173 VTAIL.n90 VSUBS 0.013039f
C174 VTAIL.n91 VSUBS 0.03082f
C175 VTAIL.n92 VSUBS 0.013806f
C176 VTAIL.n93 VSUBS 0.024266f
C177 VTAIL.n94 VSUBS 0.013039f
C178 VTAIL.n95 VSUBS 0.03082f
C179 VTAIL.n96 VSUBS 0.013806f
C180 VTAIL.n97 VSUBS 0.024266f
C181 VTAIL.n98 VSUBS 0.013039f
C182 VTAIL.n99 VSUBS 0.03082f
C183 VTAIL.n100 VSUBS 0.013806f
C184 VTAIL.n101 VSUBS 0.024266f
C185 VTAIL.n102 VSUBS 0.013039f
C186 VTAIL.n103 VSUBS 0.03082f
C187 VTAIL.n104 VSUBS 0.013806f
C188 VTAIL.n105 VSUBS 0.024266f
C189 VTAIL.n106 VSUBS 0.013039f
C190 VTAIL.n107 VSUBS 0.03082f
C191 VTAIL.n108 VSUBS 0.013806f
C192 VTAIL.n109 VSUBS 0.169406f
C193 VTAIL.t14 VSUBS 0.065966f
C194 VTAIL.n110 VSUBS 0.023115f
C195 VTAIL.n111 VSUBS 0.019606f
C196 VTAIL.n112 VSUBS 0.013039f
C197 VTAIL.n113 VSUBS 1.52407f
C198 VTAIL.n114 VSUBS 0.024266f
C199 VTAIL.n115 VSUBS 0.013039f
C200 VTAIL.n116 VSUBS 0.013806f
C201 VTAIL.n117 VSUBS 0.03082f
C202 VTAIL.n118 VSUBS 0.03082f
C203 VTAIL.n119 VSUBS 0.013806f
C204 VTAIL.n120 VSUBS 0.013039f
C205 VTAIL.n121 VSUBS 0.024266f
C206 VTAIL.n122 VSUBS 0.024266f
C207 VTAIL.n123 VSUBS 0.013039f
C208 VTAIL.n124 VSUBS 0.013806f
C209 VTAIL.n125 VSUBS 0.03082f
C210 VTAIL.n126 VSUBS 0.03082f
C211 VTAIL.n127 VSUBS 0.013806f
C212 VTAIL.n128 VSUBS 0.013039f
C213 VTAIL.n129 VSUBS 0.024266f
C214 VTAIL.n130 VSUBS 0.024266f
C215 VTAIL.n131 VSUBS 0.013039f
C216 VTAIL.n132 VSUBS 0.013806f
C217 VTAIL.n133 VSUBS 0.03082f
C218 VTAIL.n134 VSUBS 0.03082f
C219 VTAIL.n135 VSUBS 0.013806f
C220 VTAIL.n136 VSUBS 0.013039f
C221 VTAIL.n137 VSUBS 0.024266f
C222 VTAIL.n138 VSUBS 0.024266f
C223 VTAIL.n139 VSUBS 0.013039f
C224 VTAIL.n140 VSUBS 0.013806f
C225 VTAIL.n141 VSUBS 0.03082f
C226 VTAIL.n142 VSUBS 0.03082f
C227 VTAIL.n143 VSUBS 0.013806f
C228 VTAIL.n144 VSUBS 0.013039f
C229 VTAIL.n145 VSUBS 0.024266f
C230 VTAIL.n146 VSUBS 0.024266f
C231 VTAIL.n147 VSUBS 0.013039f
C232 VTAIL.n148 VSUBS 0.013806f
C233 VTAIL.n149 VSUBS 0.03082f
C234 VTAIL.n150 VSUBS 0.03082f
C235 VTAIL.n151 VSUBS 0.03082f
C236 VTAIL.n152 VSUBS 0.013806f
C237 VTAIL.n153 VSUBS 0.013039f
C238 VTAIL.n154 VSUBS 0.024266f
C239 VTAIL.n155 VSUBS 0.024266f
C240 VTAIL.n156 VSUBS 0.013039f
C241 VTAIL.n157 VSUBS 0.013423f
C242 VTAIL.n158 VSUBS 0.013423f
C243 VTAIL.n159 VSUBS 0.03082f
C244 VTAIL.n160 VSUBS 0.071814f
C245 VTAIL.n161 VSUBS 0.013806f
C246 VTAIL.n162 VSUBS 0.013039f
C247 VTAIL.n163 VSUBS 0.060398f
C248 VTAIL.n164 VSUBS 0.036118f
C249 VTAIL.n165 VSUBS 0.136064f
C250 VTAIL.t15 VSUBS 0.283221f
C251 VTAIL.t11 VSUBS 0.283221f
C252 VTAIL.n166 VSUBS 2.16945f
C253 VTAIL.n167 VSUBS 0.706534f
C254 VTAIL.n168 VSUBS 0.025841f
C255 VTAIL.n169 VSUBS 0.024266f
C256 VTAIL.n170 VSUBS 0.013039f
C257 VTAIL.n171 VSUBS 0.03082f
C258 VTAIL.n172 VSUBS 0.013806f
C259 VTAIL.n173 VSUBS 0.024266f
C260 VTAIL.n174 VSUBS 0.013039f
C261 VTAIL.n175 VSUBS 0.03082f
C262 VTAIL.n176 VSUBS 0.013806f
C263 VTAIL.n177 VSUBS 0.024266f
C264 VTAIL.n178 VSUBS 0.013039f
C265 VTAIL.n179 VSUBS 0.03082f
C266 VTAIL.n180 VSUBS 0.013806f
C267 VTAIL.n181 VSUBS 0.024266f
C268 VTAIL.n182 VSUBS 0.013039f
C269 VTAIL.n183 VSUBS 0.03082f
C270 VTAIL.n184 VSUBS 0.013806f
C271 VTAIL.n185 VSUBS 0.024266f
C272 VTAIL.n186 VSUBS 0.013039f
C273 VTAIL.n187 VSUBS 0.03082f
C274 VTAIL.n188 VSUBS 0.013806f
C275 VTAIL.n189 VSUBS 0.024266f
C276 VTAIL.n190 VSUBS 0.013039f
C277 VTAIL.n191 VSUBS 0.03082f
C278 VTAIL.n192 VSUBS 0.013806f
C279 VTAIL.n193 VSUBS 0.169406f
C280 VTAIL.t13 VSUBS 0.065966f
C281 VTAIL.n194 VSUBS 0.023115f
C282 VTAIL.n195 VSUBS 0.019606f
C283 VTAIL.n196 VSUBS 0.013039f
C284 VTAIL.n197 VSUBS 1.52407f
C285 VTAIL.n198 VSUBS 0.024266f
C286 VTAIL.n199 VSUBS 0.013039f
C287 VTAIL.n200 VSUBS 0.013806f
C288 VTAIL.n201 VSUBS 0.03082f
C289 VTAIL.n202 VSUBS 0.03082f
C290 VTAIL.n203 VSUBS 0.013806f
C291 VTAIL.n204 VSUBS 0.013039f
C292 VTAIL.n205 VSUBS 0.024266f
C293 VTAIL.n206 VSUBS 0.024266f
C294 VTAIL.n207 VSUBS 0.013039f
C295 VTAIL.n208 VSUBS 0.013806f
C296 VTAIL.n209 VSUBS 0.03082f
C297 VTAIL.n210 VSUBS 0.03082f
C298 VTAIL.n211 VSUBS 0.013806f
C299 VTAIL.n212 VSUBS 0.013039f
C300 VTAIL.n213 VSUBS 0.024266f
C301 VTAIL.n214 VSUBS 0.024266f
C302 VTAIL.n215 VSUBS 0.013039f
C303 VTAIL.n216 VSUBS 0.013806f
C304 VTAIL.n217 VSUBS 0.03082f
C305 VTAIL.n218 VSUBS 0.03082f
C306 VTAIL.n219 VSUBS 0.013806f
C307 VTAIL.n220 VSUBS 0.013039f
C308 VTAIL.n221 VSUBS 0.024266f
C309 VTAIL.n222 VSUBS 0.024266f
C310 VTAIL.n223 VSUBS 0.013039f
C311 VTAIL.n224 VSUBS 0.013806f
C312 VTAIL.n225 VSUBS 0.03082f
C313 VTAIL.n226 VSUBS 0.03082f
C314 VTAIL.n227 VSUBS 0.013806f
C315 VTAIL.n228 VSUBS 0.013039f
C316 VTAIL.n229 VSUBS 0.024266f
C317 VTAIL.n230 VSUBS 0.024266f
C318 VTAIL.n231 VSUBS 0.013039f
C319 VTAIL.n232 VSUBS 0.013806f
C320 VTAIL.n233 VSUBS 0.03082f
C321 VTAIL.n234 VSUBS 0.03082f
C322 VTAIL.n235 VSUBS 0.03082f
C323 VTAIL.n236 VSUBS 0.013806f
C324 VTAIL.n237 VSUBS 0.013039f
C325 VTAIL.n238 VSUBS 0.024266f
C326 VTAIL.n239 VSUBS 0.024266f
C327 VTAIL.n240 VSUBS 0.013039f
C328 VTAIL.n241 VSUBS 0.013423f
C329 VTAIL.n242 VSUBS 0.013423f
C330 VTAIL.n243 VSUBS 0.03082f
C331 VTAIL.n244 VSUBS 0.071814f
C332 VTAIL.n245 VSUBS 0.013806f
C333 VTAIL.n246 VSUBS 0.013039f
C334 VTAIL.n247 VSUBS 0.060398f
C335 VTAIL.n248 VSUBS 0.036118f
C336 VTAIL.n249 VSUBS 1.50068f
C337 VTAIL.n250 VSUBS 0.025841f
C338 VTAIL.n251 VSUBS 0.024266f
C339 VTAIL.n252 VSUBS 0.013039f
C340 VTAIL.n253 VSUBS 0.03082f
C341 VTAIL.n254 VSUBS 0.013806f
C342 VTAIL.n255 VSUBS 0.024266f
C343 VTAIL.n256 VSUBS 0.013039f
C344 VTAIL.n257 VSUBS 0.03082f
C345 VTAIL.n258 VSUBS 0.03082f
C346 VTAIL.n259 VSUBS 0.013806f
C347 VTAIL.n260 VSUBS 0.024266f
C348 VTAIL.n261 VSUBS 0.013039f
C349 VTAIL.n262 VSUBS 0.03082f
C350 VTAIL.n263 VSUBS 0.013806f
C351 VTAIL.n264 VSUBS 0.024266f
C352 VTAIL.n265 VSUBS 0.013039f
C353 VTAIL.n266 VSUBS 0.03082f
C354 VTAIL.n267 VSUBS 0.013806f
C355 VTAIL.n268 VSUBS 0.024266f
C356 VTAIL.n269 VSUBS 0.013039f
C357 VTAIL.n270 VSUBS 0.03082f
C358 VTAIL.n271 VSUBS 0.013806f
C359 VTAIL.n272 VSUBS 0.024266f
C360 VTAIL.n273 VSUBS 0.013039f
C361 VTAIL.n274 VSUBS 0.03082f
C362 VTAIL.n275 VSUBS 0.013806f
C363 VTAIL.n276 VSUBS 0.169406f
C364 VTAIL.t2 VSUBS 0.065966f
C365 VTAIL.n277 VSUBS 0.023115f
C366 VTAIL.n278 VSUBS 0.019606f
C367 VTAIL.n279 VSUBS 0.013039f
C368 VTAIL.n280 VSUBS 1.52407f
C369 VTAIL.n281 VSUBS 0.024266f
C370 VTAIL.n282 VSUBS 0.013039f
C371 VTAIL.n283 VSUBS 0.013806f
C372 VTAIL.n284 VSUBS 0.03082f
C373 VTAIL.n285 VSUBS 0.03082f
C374 VTAIL.n286 VSUBS 0.013806f
C375 VTAIL.n287 VSUBS 0.013039f
C376 VTAIL.n288 VSUBS 0.024266f
C377 VTAIL.n289 VSUBS 0.024266f
C378 VTAIL.n290 VSUBS 0.013039f
C379 VTAIL.n291 VSUBS 0.013806f
C380 VTAIL.n292 VSUBS 0.03082f
C381 VTAIL.n293 VSUBS 0.03082f
C382 VTAIL.n294 VSUBS 0.013806f
C383 VTAIL.n295 VSUBS 0.013039f
C384 VTAIL.n296 VSUBS 0.024266f
C385 VTAIL.n297 VSUBS 0.024266f
C386 VTAIL.n298 VSUBS 0.013039f
C387 VTAIL.n299 VSUBS 0.013806f
C388 VTAIL.n300 VSUBS 0.03082f
C389 VTAIL.n301 VSUBS 0.03082f
C390 VTAIL.n302 VSUBS 0.013806f
C391 VTAIL.n303 VSUBS 0.013039f
C392 VTAIL.n304 VSUBS 0.024266f
C393 VTAIL.n305 VSUBS 0.024266f
C394 VTAIL.n306 VSUBS 0.013039f
C395 VTAIL.n307 VSUBS 0.013806f
C396 VTAIL.n308 VSUBS 0.03082f
C397 VTAIL.n309 VSUBS 0.03082f
C398 VTAIL.n310 VSUBS 0.013806f
C399 VTAIL.n311 VSUBS 0.013039f
C400 VTAIL.n312 VSUBS 0.024266f
C401 VTAIL.n313 VSUBS 0.024266f
C402 VTAIL.n314 VSUBS 0.013039f
C403 VTAIL.n315 VSUBS 0.013806f
C404 VTAIL.n316 VSUBS 0.03082f
C405 VTAIL.n317 VSUBS 0.03082f
C406 VTAIL.n318 VSUBS 0.013806f
C407 VTAIL.n319 VSUBS 0.013039f
C408 VTAIL.n320 VSUBS 0.024266f
C409 VTAIL.n321 VSUBS 0.024266f
C410 VTAIL.n322 VSUBS 0.013039f
C411 VTAIL.n323 VSUBS 0.013423f
C412 VTAIL.n324 VSUBS 0.013423f
C413 VTAIL.n325 VSUBS 0.03082f
C414 VTAIL.n326 VSUBS 0.071814f
C415 VTAIL.n327 VSUBS 0.013806f
C416 VTAIL.n328 VSUBS 0.013039f
C417 VTAIL.n329 VSUBS 0.060398f
C418 VTAIL.n330 VSUBS 0.036118f
C419 VTAIL.n331 VSUBS 1.50068f
C420 VTAIL.t6 VSUBS 0.283221f
C421 VTAIL.t7 VSUBS 0.283221f
C422 VTAIL.n332 VSUBS 2.16947f
C423 VTAIL.n333 VSUBS 0.706521f
C424 VTAIL.n334 VSUBS 0.025841f
C425 VTAIL.n335 VSUBS 0.024266f
C426 VTAIL.n336 VSUBS 0.013039f
C427 VTAIL.n337 VSUBS 0.03082f
C428 VTAIL.n338 VSUBS 0.013806f
C429 VTAIL.n339 VSUBS 0.024266f
C430 VTAIL.n340 VSUBS 0.013039f
C431 VTAIL.n341 VSUBS 0.03082f
C432 VTAIL.n342 VSUBS 0.03082f
C433 VTAIL.n343 VSUBS 0.013806f
C434 VTAIL.n344 VSUBS 0.024266f
C435 VTAIL.n345 VSUBS 0.013039f
C436 VTAIL.n346 VSUBS 0.03082f
C437 VTAIL.n347 VSUBS 0.013806f
C438 VTAIL.n348 VSUBS 0.024266f
C439 VTAIL.n349 VSUBS 0.013039f
C440 VTAIL.n350 VSUBS 0.03082f
C441 VTAIL.n351 VSUBS 0.013806f
C442 VTAIL.n352 VSUBS 0.024266f
C443 VTAIL.n353 VSUBS 0.013039f
C444 VTAIL.n354 VSUBS 0.03082f
C445 VTAIL.n355 VSUBS 0.013806f
C446 VTAIL.n356 VSUBS 0.024266f
C447 VTAIL.n357 VSUBS 0.013039f
C448 VTAIL.n358 VSUBS 0.03082f
C449 VTAIL.n359 VSUBS 0.013806f
C450 VTAIL.n360 VSUBS 0.169406f
C451 VTAIL.t3 VSUBS 0.065966f
C452 VTAIL.n361 VSUBS 0.023115f
C453 VTAIL.n362 VSUBS 0.019606f
C454 VTAIL.n363 VSUBS 0.013039f
C455 VTAIL.n364 VSUBS 1.52407f
C456 VTAIL.n365 VSUBS 0.024266f
C457 VTAIL.n366 VSUBS 0.013039f
C458 VTAIL.n367 VSUBS 0.013806f
C459 VTAIL.n368 VSUBS 0.03082f
C460 VTAIL.n369 VSUBS 0.03082f
C461 VTAIL.n370 VSUBS 0.013806f
C462 VTAIL.n371 VSUBS 0.013039f
C463 VTAIL.n372 VSUBS 0.024266f
C464 VTAIL.n373 VSUBS 0.024266f
C465 VTAIL.n374 VSUBS 0.013039f
C466 VTAIL.n375 VSUBS 0.013806f
C467 VTAIL.n376 VSUBS 0.03082f
C468 VTAIL.n377 VSUBS 0.03082f
C469 VTAIL.n378 VSUBS 0.013806f
C470 VTAIL.n379 VSUBS 0.013039f
C471 VTAIL.n380 VSUBS 0.024266f
C472 VTAIL.n381 VSUBS 0.024266f
C473 VTAIL.n382 VSUBS 0.013039f
C474 VTAIL.n383 VSUBS 0.013806f
C475 VTAIL.n384 VSUBS 0.03082f
C476 VTAIL.n385 VSUBS 0.03082f
C477 VTAIL.n386 VSUBS 0.013806f
C478 VTAIL.n387 VSUBS 0.013039f
C479 VTAIL.n388 VSUBS 0.024266f
C480 VTAIL.n389 VSUBS 0.024266f
C481 VTAIL.n390 VSUBS 0.013039f
C482 VTAIL.n391 VSUBS 0.013806f
C483 VTAIL.n392 VSUBS 0.03082f
C484 VTAIL.n393 VSUBS 0.03082f
C485 VTAIL.n394 VSUBS 0.013806f
C486 VTAIL.n395 VSUBS 0.013039f
C487 VTAIL.n396 VSUBS 0.024266f
C488 VTAIL.n397 VSUBS 0.024266f
C489 VTAIL.n398 VSUBS 0.013039f
C490 VTAIL.n399 VSUBS 0.013806f
C491 VTAIL.n400 VSUBS 0.03082f
C492 VTAIL.n401 VSUBS 0.03082f
C493 VTAIL.n402 VSUBS 0.013806f
C494 VTAIL.n403 VSUBS 0.013039f
C495 VTAIL.n404 VSUBS 0.024266f
C496 VTAIL.n405 VSUBS 0.024266f
C497 VTAIL.n406 VSUBS 0.013039f
C498 VTAIL.n407 VSUBS 0.013423f
C499 VTAIL.n408 VSUBS 0.013423f
C500 VTAIL.n409 VSUBS 0.03082f
C501 VTAIL.n410 VSUBS 0.071814f
C502 VTAIL.n411 VSUBS 0.013806f
C503 VTAIL.n412 VSUBS 0.013039f
C504 VTAIL.n413 VSUBS 0.060398f
C505 VTAIL.n414 VSUBS 0.036118f
C506 VTAIL.n415 VSUBS 0.136064f
C507 VTAIL.n416 VSUBS 0.025841f
C508 VTAIL.n417 VSUBS 0.024266f
C509 VTAIL.n418 VSUBS 0.013039f
C510 VTAIL.n419 VSUBS 0.03082f
C511 VTAIL.n420 VSUBS 0.013806f
C512 VTAIL.n421 VSUBS 0.024266f
C513 VTAIL.n422 VSUBS 0.013039f
C514 VTAIL.n423 VSUBS 0.03082f
C515 VTAIL.n424 VSUBS 0.03082f
C516 VTAIL.n425 VSUBS 0.013806f
C517 VTAIL.n426 VSUBS 0.024266f
C518 VTAIL.n427 VSUBS 0.013039f
C519 VTAIL.n428 VSUBS 0.03082f
C520 VTAIL.n429 VSUBS 0.013806f
C521 VTAIL.n430 VSUBS 0.024266f
C522 VTAIL.n431 VSUBS 0.013039f
C523 VTAIL.n432 VSUBS 0.03082f
C524 VTAIL.n433 VSUBS 0.013806f
C525 VTAIL.n434 VSUBS 0.024266f
C526 VTAIL.n435 VSUBS 0.013039f
C527 VTAIL.n436 VSUBS 0.03082f
C528 VTAIL.n437 VSUBS 0.013806f
C529 VTAIL.n438 VSUBS 0.024266f
C530 VTAIL.n439 VSUBS 0.013039f
C531 VTAIL.n440 VSUBS 0.03082f
C532 VTAIL.n441 VSUBS 0.013806f
C533 VTAIL.n442 VSUBS 0.169406f
C534 VTAIL.t12 VSUBS 0.065966f
C535 VTAIL.n443 VSUBS 0.023115f
C536 VTAIL.n444 VSUBS 0.019606f
C537 VTAIL.n445 VSUBS 0.013039f
C538 VTAIL.n446 VSUBS 1.52407f
C539 VTAIL.n447 VSUBS 0.024266f
C540 VTAIL.n448 VSUBS 0.013039f
C541 VTAIL.n449 VSUBS 0.013806f
C542 VTAIL.n450 VSUBS 0.03082f
C543 VTAIL.n451 VSUBS 0.03082f
C544 VTAIL.n452 VSUBS 0.013806f
C545 VTAIL.n453 VSUBS 0.013039f
C546 VTAIL.n454 VSUBS 0.024266f
C547 VTAIL.n455 VSUBS 0.024266f
C548 VTAIL.n456 VSUBS 0.013039f
C549 VTAIL.n457 VSUBS 0.013806f
C550 VTAIL.n458 VSUBS 0.03082f
C551 VTAIL.n459 VSUBS 0.03082f
C552 VTAIL.n460 VSUBS 0.013806f
C553 VTAIL.n461 VSUBS 0.013039f
C554 VTAIL.n462 VSUBS 0.024266f
C555 VTAIL.n463 VSUBS 0.024266f
C556 VTAIL.n464 VSUBS 0.013039f
C557 VTAIL.n465 VSUBS 0.013806f
C558 VTAIL.n466 VSUBS 0.03082f
C559 VTAIL.n467 VSUBS 0.03082f
C560 VTAIL.n468 VSUBS 0.013806f
C561 VTAIL.n469 VSUBS 0.013039f
C562 VTAIL.n470 VSUBS 0.024266f
C563 VTAIL.n471 VSUBS 0.024266f
C564 VTAIL.n472 VSUBS 0.013039f
C565 VTAIL.n473 VSUBS 0.013806f
C566 VTAIL.n474 VSUBS 0.03082f
C567 VTAIL.n475 VSUBS 0.03082f
C568 VTAIL.n476 VSUBS 0.013806f
C569 VTAIL.n477 VSUBS 0.013039f
C570 VTAIL.n478 VSUBS 0.024266f
C571 VTAIL.n479 VSUBS 0.024266f
C572 VTAIL.n480 VSUBS 0.013039f
C573 VTAIL.n481 VSUBS 0.013806f
C574 VTAIL.n482 VSUBS 0.03082f
C575 VTAIL.n483 VSUBS 0.03082f
C576 VTAIL.n484 VSUBS 0.013806f
C577 VTAIL.n485 VSUBS 0.013039f
C578 VTAIL.n486 VSUBS 0.024266f
C579 VTAIL.n487 VSUBS 0.024266f
C580 VTAIL.n488 VSUBS 0.013039f
C581 VTAIL.n489 VSUBS 0.013423f
C582 VTAIL.n490 VSUBS 0.013423f
C583 VTAIL.n491 VSUBS 0.03082f
C584 VTAIL.n492 VSUBS 0.071814f
C585 VTAIL.n493 VSUBS 0.013806f
C586 VTAIL.n494 VSUBS 0.013039f
C587 VTAIL.n495 VSUBS 0.060398f
C588 VTAIL.n496 VSUBS 0.036118f
C589 VTAIL.n497 VSUBS 0.136064f
C590 VTAIL.t10 VSUBS 0.283221f
C591 VTAIL.t9 VSUBS 0.283221f
C592 VTAIL.n498 VSUBS 2.16947f
C593 VTAIL.n499 VSUBS 0.706521f
C594 VTAIL.n500 VSUBS 0.025841f
C595 VTAIL.n501 VSUBS 0.024266f
C596 VTAIL.n502 VSUBS 0.013039f
C597 VTAIL.n503 VSUBS 0.03082f
C598 VTAIL.n504 VSUBS 0.013806f
C599 VTAIL.n505 VSUBS 0.024266f
C600 VTAIL.n506 VSUBS 0.013039f
C601 VTAIL.n507 VSUBS 0.03082f
C602 VTAIL.n508 VSUBS 0.03082f
C603 VTAIL.n509 VSUBS 0.013806f
C604 VTAIL.n510 VSUBS 0.024266f
C605 VTAIL.n511 VSUBS 0.013039f
C606 VTAIL.n512 VSUBS 0.03082f
C607 VTAIL.n513 VSUBS 0.013806f
C608 VTAIL.n514 VSUBS 0.024266f
C609 VTAIL.n515 VSUBS 0.013039f
C610 VTAIL.n516 VSUBS 0.03082f
C611 VTAIL.n517 VSUBS 0.013806f
C612 VTAIL.n518 VSUBS 0.024266f
C613 VTAIL.n519 VSUBS 0.013039f
C614 VTAIL.n520 VSUBS 0.03082f
C615 VTAIL.n521 VSUBS 0.013806f
C616 VTAIL.n522 VSUBS 0.024266f
C617 VTAIL.n523 VSUBS 0.013039f
C618 VTAIL.n524 VSUBS 0.03082f
C619 VTAIL.n525 VSUBS 0.013806f
C620 VTAIL.n526 VSUBS 0.169406f
C621 VTAIL.t8 VSUBS 0.065966f
C622 VTAIL.n527 VSUBS 0.023115f
C623 VTAIL.n528 VSUBS 0.019606f
C624 VTAIL.n529 VSUBS 0.013039f
C625 VTAIL.n530 VSUBS 1.52407f
C626 VTAIL.n531 VSUBS 0.024266f
C627 VTAIL.n532 VSUBS 0.013039f
C628 VTAIL.n533 VSUBS 0.013806f
C629 VTAIL.n534 VSUBS 0.03082f
C630 VTAIL.n535 VSUBS 0.03082f
C631 VTAIL.n536 VSUBS 0.013806f
C632 VTAIL.n537 VSUBS 0.013039f
C633 VTAIL.n538 VSUBS 0.024266f
C634 VTAIL.n539 VSUBS 0.024266f
C635 VTAIL.n540 VSUBS 0.013039f
C636 VTAIL.n541 VSUBS 0.013806f
C637 VTAIL.n542 VSUBS 0.03082f
C638 VTAIL.n543 VSUBS 0.03082f
C639 VTAIL.n544 VSUBS 0.013806f
C640 VTAIL.n545 VSUBS 0.013039f
C641 VTAIL.n546 VSUBS 0.024266f
C642 VTAIL.n547 VSUBS 0.024266f
C643 VTAIL.n548 VSUBS 0.013039f
C644 VTAIL.n549 VSUBS 0.013806f
C645 VTAIL.n550 VSUBS 0.03082f
C646 VTAIL.n551 VSUBS 0.03082f
C647 VTAIL.n552 VSUBS 0.013806f
C648 VTAIL.n553 VSUBS 0.013039f
C649 VTAIL.n554 VSUBS 0.024266f
C650 VTAIL.n555 VSUBS 0.024266f
C651 VTAIL.n556 VSUBS 0.013039f
C652 VTAIL.n557 VSUBS 0.013806f
C653 VTAIL.n558 VSUBS 0.03082f
C654 VTAIL.n559 VSUBS 0.03082f
C655 VTAIL.n560 VSUBS 0.013806f
C656 VTAIL.n561 VSUBS 0.013039f
C657 VTAIL.n562 VSUBS 0.024266f
C658 VTAIL.n563 VSUBS 0.024266f
C659 VTAIL.n564 VSUBS 0.013039f
C660 VTAIL.n565 VSUBS 0.013806f
C661 VTAIL.n566 VSUBS 0.03082f
C662 VTAIL.n567 VSUBS 0.03082f
C663 VTAIL.n568 VSUBS 0.013806f
C664 VTAIL.n569 VSUBS 0.013039f
C665 VTAIL.n570 VSUBS 0.024266f
C666 VTAIL.n571 VSUBS 0.024266f
C667 VTAIL.n572 VSUBS 0.013039f
C668 VTAIL.n573 VSUBS 0.013423f
C669 VTAIL.n574 VSUBS 0.013423f
C670 VTAIL.n575 VSUBS 0.03082f
C671 VTAIL.n576 VSUBS 0.071814f
C672 VTAIL.n577 VSUBS 0.013806f
C673 VTAIL.n578 VSUBS 0.013039f
C674 VTAIL.n579 VSUBS 0.060398f
C675 VTAIL.n580 VSUBS 0.036118f
C676 VTAIL.n581 VSUBS 1.50068f
C677 VTAIL.n582 VSUBS 0.025841f
C678 VTAIL.n583 VSUBS 0.024266f
C679 VTAIL.n584 VSUBS 0.013039f
C680 VTAIL.n585 VSUBS 0.03082f
C681 VTAIL.n586 VSUBS 0.013806f
C682 VTAIL.n587 VSUBS 0.024266f
C683 VTAIL.n588 VSUBS 0.013039f
C684 VTAIL.n589 VSUBS 0.03082f
C685 VTAIL.n590 VSUBS 0.013806f
C686 VTAIL.n591 VSUBS 0.024266f
C687 VTAIL.n592 VSUBS 0.013039f
C688 VTAIL.n593 VSUBS 0.03082f
C689 VTAIL.n594 VSUBS 0.013806f
C690 VTAIL.n595 VSUBS 0.024266f
C691 VTAIL.n596 VSUBS 0.013039f
C692 VTAIL.n597 VSUBS 0.03082f
C693 VTAIL.n598 VSUBS 0.013806f
C694 VTAIL.n599 VSUBS 0.024266f
C695 VTAIL.n600 VSUBS 0.013039f
C696 VTAIL.n601 VSUBS 0.03082f
C697 VTAIL.n602 VSUBS 0.013806f
C698 VTAIL.n603 VSUBS 0.024266f
C699 VTAIL.n604 VSUBS 0.013039f
C700 VTAIL.n605 VSUBS 0.03082f
C701 VTAIL.n606 VSUBS 0.013806f
C702 VTAIL.n607 VSUBS 0.169406f
C703 VTAIL.t4 VSUBS 0.065966f
C704 VTAIL.n608 VSUBS 0.023115f
C705 VTAIL.n609 VSUBS 0.019606f
C706 VTAIL.n610 VSUBS 0.013039f
C707 VTAIL.n611 VSUBS 1.52407f
C708 VTAIL.n612 VSUBS 0.024266f
C709 VTAIL.n613 VSUBS 0.013039f
C710 VTAIL.n614 VSUBS 0.013806f
C711 VTAIL.n615 VSUBS 0.03082f
C712 VTAIL.n616 VSUBS 0.03082f
C713 VTAIL.n617 VSUBS 0.013806f
C714 VTAIL.n618 VSUBS 0.013039f
C715 VTAIL.n619 VSUBS 0.024266f
C716 VTAIL.n620 VSUBS 0.024266f
C717 VTAIL.n621 VSUBS 0.013039f
C718 VTAIL.n622 VSUBS 0.013806f
C719 VTAIL.n623 VSUBS 0.03082f
C720 VTAIL.n624 VSUBS 0.03082f
C721 VTAIL.n625 VSUBS 0.013806f
C722 VTAIL.n626 VSUBS 0.013039f
C723 VTAIL.n627 VSUBS 0.024266f
C724 VTAIL.n628 VSUBS 0.024266f
C725 VTAIL.n629 VSUBS 0.013039f
C726 VTAIL.n630 VSUBS 0.013806f
C727 VTAIL.n631 VSUBS 0.03082f
C728 VTAIL.n632 VSUBS 0.03082f
C729 VTAIL.n633 VSUBS 0.013806f
C730 VTAIL.n634 VSUBS 0.013039f
C731 VTAIL.n635 VSUBS 0.024266f
C732 VTAIL.n636 VSUBS 0.024266f
C733 VTAIL.n637 VSUBS 0.013039f
C734 VTAIL.n638 VSUBS 0.013806f
C735 VTAIL.n639 VSUBS 0.03082f
C736 VTAIL.n640 VSUBS 0.03082f
C737 VTAIL.n641 VSUBS 0.013806f
C738 VTAIL.n642 VSUBS 0.013039f
C739 VTAIL.n643 VSUBS 0.024266f
C740 VTAIL.n644 VSUBS 0.024266f
C741 VTAIL.n645 VSUBS 0.013039f
C742 VTAIL.n646 VSUBS 0.013806f
C743 VTAIL.n647 VSUBS 0.03082f
C744 VTAIL.n648 VSUBS 0.03082f
C745 VTAIL.n649 VSUBS 0.03082f
C746 VTAIL.n650 VSUBS 0.013806f
C747 VTAIL.n651 VSUBS 0.013039f
C748 VTAIL.n652 VSUBS 0.024266f
C749 VTAIL.n653 VSUBS 0.024266f
C750 VTAIL.n654 VSUBS 0.013039f
C751 VTAIL.n655 VSUBS 0.013423f
C752 VTAIL.n656 VSUBS 0.013423f
C753 VTAIL.n657 VSUBS 0.03082f
C754 VTAIL.n658 VSUBS 0.071814f
C755 VTAIL.n659 VSUBS 0.013806f
C756 VTAIL.n660 VSUBS 0.013039f
C757 VTAIL.n661 VSUBS 0.060398f
C758 VTAIL.n662 VSUBS 0.036118f
C759 VTAIL.n663 VSUBS 1.49613f
C760 VP.n0 VSUBS 0.067635f
C761 VP.t7 VSUBS 1.70267f
C762 VP.n1 VSUBS 0.668196f
C763 VP.n2 VSUBS 0.067635f
C764 VP.t2 VSUBS 1.70267f
C765 VP.t4 VSUBS 1.70267f
C766 VP.n3 VSUBS 0.290096f
C767 VP.t5 VSUBS 1.70267f
C768 VP.t6 VSUBS 1.72902f
C769 VP.n4 VSUBS 0.63653f
C770 VP.n5 VSUBS 0.669022f
C771 VP.n6 VSUBS 0.668196f
C772 VP.n7 VSUBS 0.011502f
C773 VP.n8 VSUBS 0.649194f
C774 VP.n9 VSUBS 2.30032f
C775 VP.n10 VSUBS 2.34126f
C776 VP.t1 VSUBS 1.70267f
C777 VP.n11 VSUBS 0.649194f
C778 VP.n12 VSUBS 0.011502f
C779 VP.n13 VSUBS 0.067635f
C780 VP.n14 VSUBS 0.084425f
C781 VP.n15 VSUBS 0.084425f
C782 VP.t3 VSUBS 1.70267f
C783 VP.n16 VSUBS 0.668196f
C784 VP.n17 VSUBS 0.011502f
C785 VP.t0 VSUBS 1.70267f
C786 VP.n18 VSUBS 0.649194f
C787 VP.n19 VSUBS 0.03928f
C788 B.n0 VSUBS 0.006864f
C789 B.n1 VSUBS 0.006864f
C790 B.n2 VSUBS 0.010152f
C791 B.n3 VSUBS 0.00778f
C792 B.n4 VSUBS 0.00778f
C793 B.n5 VSUBS 0.00778f
C794 B.n6 VSUBS 0.00778f
C795 B.n7 VSUBS 0.00778f
C796 B.n8 VSUBS 0.00778f
C797 B.n9 VSUBS 0.00778f
C798 B.n10 VSUBS 0.00778f
C799 B.n11 VSUBS 0.00778f
C800 B.n12 VSUBS 0.00778f
C801 B.n13 VSUBS 0.00778f
C802 B.n14 VSUBS 0.019747f
C803 B.n15 VSUBS 0.00778f
C804 B.n16 VSUBS 0.00778f
C805 B.n17 VSUBS 0.00778f
C806 B.n18 VSUBS 0.00778f
C807 B.n19 VSUBS 0.00778f
C808 B.n20 VSUBS 0.00778f
C809 B.n21 VSUBS 0.00778f
C810 B.n22 VSUBS 0.00778f
C811 B.n23 VSUBS 0.00778f
C812 B.n24 VSUBS 0.00778f
C813 B.n25 VSUBS 0.00778f
C814 B.n26 VSUBS 0.00778f
C815 B.n27 VSUBS 0.00778f
C816 B.n28 VSUBS 0.00778f
C817 B.n29 VSUBS 0.00778f
C818 B.n30 VSUBS 0.00778f
C819 B.n31 VSUBS 0.00778f
C820 B.n32 VSUBS 0.00778f
C821 B.n33 VSUBS 0.00778f
C822 B.n34 VSUBS 0.00778f
C823 B.n35 VSUBS 0.00778f
C824 B.n36 VSUBS 0.00778f
C825 B.n37 VSUBS 0.00778f
C826 B.n38 VSUBS 0.00778f
C827 B.n39 VSUBS 0.00778f
C828 B.t7 VSUBS 0.304754f
C829 B.t8 VSUBS 0.319526f
C830 B.t6 VSUBS 0.5397f
C831 B.n40 VSUBS 0.423008f
C832 B.n41 VSUBS 0.31267f
C833 B.n42 VSUBS 0.00778f
C834 B.n43 VSUBS 0.00778f
C835 B.n44 VSUBS 0.00778f
C836 B.n45 VSUBS 0.00778f
C837 B.t1 VSUBS 0.304758f
C838 B.t2 VSUBS 0.319529f
C839 B.t0 VSUBS 0.5397f
C840 B.n46 VSUBS 0.423004f
C841 B.n47 VSUBS 0.312667f
C842 B.n48 VSUBS 0.00778f
C843 B.n49 VSUBS 0.00778f
C844 B.n50 VSUBS 0.00778f
C845 B.n51 VSUBS 0.00778f
C846 B.n52 VSUBS 0.00778f
C847 B.n53 VSUBS 0.00778f
C848 B.n54 VSUBS 0.00778f
C849 B.n55 VSUBS 0.00778f
C850 B.n56 VSUBS 0.00778f
C851 B.n57 VSUBS 0.00778f
C852 B.n58 VSUBS 0.00778f
C853 B.n59 VSUBS 0.00778f
C854 B.n60 VSUBS 0.00778f
C855 B.n61 VSUBS 0.00778f
C856 B.n62 VSUBS 0.00778f
C857 B.n63 VSUBS 0.00778f
C858 B.n64 VSUBS 0.00778f
C859 B.n65 VSUBS 0.00778f
C860 B.n66 VSUBS 0.00778f
C861 B.n67 VSUBS 0.00778f
C862 B.n68 VSUBS 0.00778f
C863 B.n69 VSUBS 0.00778f
C864 B.n70 VSUBS 0.00778f
C865 B.n71 VSUBS 0.00778f
C866 B.n72 VSUBS 0.019747f
C867 B.n73 VSUBS 0.00778f
C868 B.n74 VSUBS 0.00778f
C869 B.n75 VSUBS 0.00778f
C870 B.n76 VSUBS 0.00778f
C871 B.n77 VSUBS 0.00778f
C872 B.n78 VSUBS 0.00778f
C873 B.n79 VSUBS 0.00778f
C874 B.n80 VSUBS 0.00778f
C875 B.n81 VSUBS 0.00778f
C876 B.n82 VSUBS 0.00778f
C877 B.n83 VSUBS 0.00778f
C878 B.n84 VSUBS 0.00778f
C879 B.n85 VSUBS 0.00778f
C880 B.n86 VSUBS 0.00778f
C881 B.n87 VSUBS 0.00778f
C882 B.n88 VSUBS 0.00778f
C883 B.n89 VSUBS 0.00778f
C884 B.n90 VSUBS 0.00778f
C885 B.n91 VSUBS 0.00778f
C886 B.n92 VSUBS 0.00778f
C887 B.n93 VSUBS 0.00778f
C888 B.n94 VSUBS 0.00778f
C889 B.n95 VSUBS 0.00778f
C890 B.n96 VSUBS 0.00778f
C891 B.n97 VSUBS 0.018693f
C892 B.n98 VSUBS 0.00778f
C893 B.n99 VSUBS 0.00778f
C894 B.n100 VSUBS 0.00778f
C895 B.n101 VSUBS 0.00778f
C896 B.n102 VSUBS 0.00778f
C897 B.n103 VSUBS 0.00778f
C898 B.n104 VSUBS 0.00778f
C899 B.n105 VSUBS 0.00778f
C900 B.n106 VSUBS 0.00778f
C901 B.n107 VSUBS 0.00778f
C902 B.n108 VSUBS 0.00778f
C903 B.n109 VSUBS 0.00778f
C904 B.n110 VSUBS 0.00778f
C905 B.n111 VSUBS 0.00778f
C906 B.n112 VSUBS 0.00778f
C907 B.n113 VSUBS 0.00778f
C908 B.n114 VSUBS 0.00778f
C909 B.n115 VSUBS 0.00778f
C910 B.n116 VSUBS 0.00778f
C911 B.n117 VSUBS 0.00778f
C912 B.n118 VSUBS 0.00778f
C913 B.n119 VSUBS 0.00778f
C914 B.n120 VSUBS 0.00778f
C915 B.n121 VSUBS 0.00778f
C916 B.n122 VSUBS 0.005377f
C917 B.n123 VSUBS 0.00778f
C918 B.n124 VSUBS 0.00778f
C919 B.n125 VSUBS 0.00778f
C920 B.n126 VSUBS 0.00778f
C921 B.n127 VSUBS 0.00778f
C922 B.t5 VSUBS 0.304754f
C923 B.t4 VSUBS 0.319526f
C924 B.t3 VSUBS 0.5397f
C925 B.n128 VSUBS 0.423008f
C926 B.n129 VSUBS 0.31267f
C927 B.n130 VSUBS 0.00778f
C928 B.n131 VSUBS 0.00778f
C929 B.n132 VSUBS 0.00778f
C930 B.n133 VSUBS 0.00778f
C931 B.n134 VSUBS 0.00778f
C932 B.n135 VSUBS 0.00778f
C933 B.n136 VSUBS 0.00778f
C934 B.n137 VSUBS 0.00778f
C935 B.n138 VSUBS 0.00778f
C936 B.n139 VSUBS 0.00778f
C937 B.n140 VSUBS 0.00778f
C938 B.n141 VSUBS 0.00778f
C939 B.n142 VSUBS 0.00778f
C940 B.n143 VSUBS 0.00778f
C941 B.n144 VSUBS 0.00778f
C942 B.n145 VSUBS 0.00778f
C943 B.n146 VSUBS 0.00778f
C944 B.n147 VSUBS 0.00778f
C945 B.n148 VSUBS 0.00778f
C946 B.n149 VSUBS 0.00778f
C947 B.n150 VSUBS 0.00778f
C948 B.n151 VSUBS 0.00778f
C949 B.n152 VSUBS 0.00778f
C950 B.n153 VSUBS 0.00778f
C951 B.n154 VSUBS 0.018693f
C952 B.n155 VSUBS 0.00778f
C953 B.n156 VSUBS 0.00778f
C954 B.n157 VSUBS 0.00778f
C955 B.n158 VSUBS 0.00778f
C956 B.n159 VSUBS 0.00778f
C957 B.n160 VSUBS 0.00778f
C958 B.n161 VSUBS 0.00778f
C959 B.n162 VSUBS 0.00778f
C960 B.n163 VSUBS 0.00778f
C961 B.n164 VSUBS 0.00778f
C962 B.n165 VSUBS 0.00778f
C963 B.n166 VSUBS 0.00778f
C964 B.n167 VSUBS 0.00778f
C965 B.n168 VSUBS 0.00778f
C966 B.n169 VSUBS 0.00778f
C967 B.n170 VSUBS 0.00778f
C968 B.n171 VSUBS 0.00778f
C969 B.n172 VSUBS 0.00778f
C970 B.n173 VSUBS 0.00778f
C971 B.n174 VSUBS 0.00778f
C972 B.n175 VSUBS 0.00778f
C973 B.n176 VSUBS 0.00778f
C974 B.n177 VSUBS 0.00778f
C975 B.n178 VSUBS 0.00778f
C976 B.n179 VSUBS 0.00778f
C977 B.n180 VSUBS 0.00778f
C978 B.n181 VSUBS 0.00778f
C979 B.n182 VSUBS 0.00778f
C980 B.n183 VSUBS 0.00778f
C981 B.n184 VSUBS 0.00778f
C982 B.n185 VSUBS 0.00778f
C983 B.n186 VSUBS 0.00778f
C984 B.n187 VSUBS 0.00778f
C985 B.n188 VSUBS 0.00778f
C986 B.n189 VSUBS 0.00778f
C987 B.n190 VSUBS 0.00778f
C988 B.n191 VSUBS 0.00778f
C989 B.n192 VSUBS 0.00778f
C990 B.n193 VSUBS 0.00778f
C991 B.n194 VSUBS 0.00778f
C992 B.n195 VSUBS 0.00778f
C993 B.n196 VSUBS 0.00778f
C994 B.n197 VSUBS 0.00778f
C995 B.n198 VSUBS 0.00778f
C996 B.n199 VSUBS 0.018693f
C997 B.n200 VSUBS 0.019747f
C998 B.n201 VSUBS 0.019747f
C999 B.n202 VSUBS 0.00778f
C1000 B.n203 VSUBS 0.00778f
C1001 B.n204 VSUBS 0.00778f
C1002 B.n205 VSUBS 0.00778f
C1003 B.n206 VSUBS 0.00778f
C1004 B.n207 VSUBS 0.00778f
C1005 B.n208 VSUBS 0.00778f
C1006 B.n209 VSUBS 0.00778f
C1007 B.n210 VSUBS 0.00778f
C1008 B.n211 VSUBS 0.00778f
C1009 B.n212 VSUBS 0.00778f
C1010 B.n213 VSUBS 0.00778f
C1011 B.n214 VSUBS 0.00778f
C1012 B.n215 VSUBS 0.00778f
C1013 B.n216 VSUBS 0.00778f
C1014 B.n217 VSUBS 0.00778f
C1015 B.n218 VSUBS 0.00778f
C1016 B.n219 VSUBS 0.00778f
C1017 B.n220 VSUBS 0.00778f
C1018 B.n221 VSUBS 0.00778f
C1019 B.n222 VSUBS 0.00778f
C1020 B.n223 VSUBS 0.00778f
C1021 B.n224 VSUBS 0.00778f
C1022 B.n225 VSUBS 0.00778f
C1023 B.n226 VSUBS 0.00778f
C1024 B.n227 VSUBS 0.00778f
C1025 B.n228 VSUBS 0.00778f
C1026 B.n229 VSUBS 0.00778f
C1027 B.n230 VSUBS 0.00778f
C1028 B.n231 VSUBS 0.00778f
C1029 B.n232 VSUBS 0.00778f
C1030 B.n233 VSUBS 0.00778f
C1031 B.n234 VSUBS 0.00778f
C1032 B.n235 VSUBS 0.00778f
C1033 B.n236 VSUBS 0.00778f
C1034 B.n237 VSUBS 0.00778f
C1035 B.n238 VSUBS 0.00778f
C1036 B.n239 VSUBS 0.00778f
C1037 B.n240 VSUBS 0.00778f
C1038 B.n241 VSUBS 0.00778f
C1039 B.n242 VSUBS 0.00778f
C1040 B.n243 VSUBS 0.00778f
C1041 B.n244 VSUBS 0.00778f
C1042 B.n245 VSUBS 0.00778f
C1043 B.n246 VSUBS 0.00778f
C1044 B.n247 VSUBS 0.00778f
C1045 B.n248 VSUBS 0.00778f
C1046 B.n249 VSUBS 0.00778f
C1047 B.n250 VSUBS 0.00778f
C1048 B.n251 VSUBS 0.00778f
C1049 B.n252 VSUBS 0.00778f
C1050 B.n253 VSUBS 0.00778f
C1051 B.n254 VSUBS 0.00778f
C1052 B.n255 VSUBS 0.00778f
C1053 B.n256 VSUBS 0.00778f
C1054 B.n257 VSUBS 0.00778f
C1055 B.n258 VSUBS 0.00778f
C1056 B.n259 VSUBS 0.00778f
C1057 B.n260 VSUBS 0.00778f
C1058 B.n261 VSUBS 0.00778f
C1059 B.n262 VSUBS 0.00778f
C1060 B.n263 VSUBS 0.00778f
C1061 B.n264 VSUBS 0.00778f
C1062 B.n265 VSUBS 0.00778f
C1063 B.n266 VSUBS 0.00778f
C1064 B.n267 VSUBS 0.00778f
C1065 B.n268 VSUBS 0.00778f
C1066 B.n269 VSUBS 0.00778f
C1067 B.n270 VSUBS 0.00778f
C1068 B.n271 VSUBS 0.00778f
C1069 B.n272 VSUBS 0.00778f
C1070 B.n273 VSUBS 0.00778f
C1071 B.n274 VSUBS 0.005377f
C1072 B.n275 VSUBS 0.018025f
C1073 B.n276 VSUBS 0.006292f
C1074 B.n277 VSUBS 0.00778f
C1075 B.n278 VSUBS 0.00778f
C1076 B.n279 VSUBS 0.00778f
C1077 B.n280 VSUBS 0.00778f
C1078 B.n281 VSUBS 0.00778f
C1079 B.n282 VSUBS 0.00778f
C1080 B.n283 VSUBS 0.00778f
C1081 B.n284 VSUBS 0.00778f
C1082 B.n285 VSUBS 0.00778f
C1083 B.n286 VSUBS 0.00778f
C1084 B.n287 VSUBS 0.00778f
C1085 B.t11 VSUBS 0.304758f
C1086 B.t10 VSUBS 0.319529f
C1087 B.t9 VSUBS 0.5397f
C1088 B.n288 VSUBS 0.423004f
C1089 B.n289 VSUBS 0.312667f
C1090 B.n290 VSUBS 0.018025f
C1091 B.n291 VSUBS 0.006292f
C1092 B.n292 VSUBS 0.00778f
C1093 B.n293 VSUBS 0.00778f
C1094 B.n294 VSUBS 0.00778f
C1095 B.n295 VSUBS 0.00778f
C1096 B.n296 VSUBS 0.00778f
C1097 B.n297 VSUBS 0.00778f
C1098 B.n298 VSUBS 0.00778f
C1099 B.n299 VSUBS 0.00778f
C1100 B.n300 VSUBS 0.00778f
C1101 B.n301 VSUBS 0.00778f
C1102 B.n302 VSUBS 0.00778f
C1103 B.n303 VSUBS 0.00778f
C1104 B.n304 VSUBS 0.00778f
C1105 B.n305 VSUBS 0.00778f
C1106 B.n306 VSUBS 0.00778f
C1107 B.n307 VSUBS 0.00778f
C1108 B.n308 VSUBS 0.00778f
C1109 B.n309 VSUBS 0.00778f
C1110 B.n310 VSUBS 0.00778f
C1111 B.n311 VSUBS 0.00778f
C1112 B.n312 VSUBS 0.00778f
C1113 B.n313 VSUBS 0.00778f
C1114 B.n314 VSUBS 0.00778f
C1115 B.n315 VSUBS 0.00778f
C1116 B.n316 VSUBS 0.00778f
C1117 B.n317 VSUBS 0.00778f
C1118 B.n318 VSUBS 0.00778f
C1119 B.n319 VSUBS 0.00778f
C1120 B.n320 VSUBS 0.00778f
C1121 B.n321 VSUBS 0.00778f
C1122 B.n322 VSUBS 0.00778f
C1123 B.n323 VSUBS 0.00778f
C1124 B.n324 VSUBS 0.00778f
C1125 B.n325 VSUBS 0.00778f
C1126 B.n326 VSUBS 0.00778f
C1127 B.n327 VSUBS 0.00778f
C1128 B.n328 VSUBS 0.00778f
C1129 B.n329 VSUBS 0.00778f
C1130 B.n330 VSUBS 0.00778f
C1131 B.n331 VSUBS 0.00778f
C1132 B.n332 VSUBS 0.00778f
C1133 B.n333 VSUBS 0.00778f
C1134 B.n334 VSUBS 0.00778f
C1135 B.n335 VSUBS 0.00778f
C1136 B.n336 VSUBS 0.00778f
C1137 B.n337 VSUBS 0.00778f
C1138 B.n338 VSUBS 0.00778f
C1139 B.n339 VSUBS 0.00778f
C1140 B.n340 VSUBS 0.00778f
C1141 B.n341 VSUBS 0.00778f
C1142 B.n342 VSUBS 0.00778f
C1143 B.n343 VSUBS 0.00778f
C1144 B.n344 VSUBS 0.00778f
C1145 B.n345 VSUBS 0.00778f
C1146 B.n346 VSUBS 0.00778f
C1147 B.n347 VSUBS 0.00778f
C1148 B.n348 VSUBS 0.00778f
C1149 B.n349 VSUBS 0.00778f
C1150 B.n350 VSUBS 0.00778f
C1151 B.n351 VSUBS 0.00778f
C1152 B.n352 VSUBS 0.00778f
C1153 B.n353 VSUBS 0.00778f
C1154 B.n354 VSUBS 0.00778f
C1155 B.n355 VSUBS 0.00778f
C1156 B.n356 VSUBS 0.00778f
C1157 B.n357 VSUBS 0.00778f
C1158 B.n358 VSUBS 0.00778f
C1159 B.n359 VSUBS 0.00778f
C1160 B.n360 VSUBS 0.00778f
C1161 B.n361 VSUBS 0.00778f
C1162 B.n362 VSUBS 0.00778f
C1163 B.n363 VSUBS 0.00778f
C1164 B.n364 VSUBS 0.00778f
C1165 B.n365 VSUBS 0.00778f
C1166 B.n366 VSUBS 0.019747f
C1167 B.n367 VSUBS 0.0189f
C1168 B.n368 VSUBS 0.019541f
C1169 B.n369 VSUBS 0.00778f
C1170 B.n370 VSUBS 0.00778f
C1171 B.n371 VSUBS 0.00778f
C1172 B.n372 VSUBS 0.00778f
C1173 B.n373 VSUBS 0.00778f
C1174 B.n374 VSUBS 0.00778f
C1175 B.n375 VSUBS 0.00778f
C1176 B.n376 VSUBS 0.00778f
C1177 B.n377 VSUBS 0.00778f
C1178 B.n378 VSUBS 0.00778f
C1179 B.n379 VSUBS 0.00778f
C1180 B.n380 VSUBS 0.00778f
C1181 B.n381 VSUBS 0.00778f
C1182 B.n382 VSUBS 0.00778f
C1183 B.n383 VSUBS 0.00778f
C1184 B.n384 VSUBS 0.00778f
C1185 B.n385 VSUBS 0.00778f
C1186 B.n386 VSUBS 0.00778f
C1187 B.n387 VSUBS 0.00778f
C1188 B.n388 VSUBS 0.00778f
C1189 B.n389 VSUBS 0.00778f
C1190 B.n390 VSUBS 0.00778f
C1191 B.n391 VSUBS 0.00778f
C1192 B.n392 VSUBS 0.00778f
C1193 B.n393 VSUBS 0.00778f
C1194 B.n394 VSUBS 0.00778f
C1195 B.n395 VSUBS 0.00778f
C1196 B.n396 VSUBS 0.00778f
C1197 B.n397 VSUBS 0.00778f
C1198 B.n398 VSUBS 0.00778f
C1199 B.n399 VSUBS 0.00778f
C1200 B.n400 VSUBS 0.00778f
C1201 B.n401 VSUBS 0.00778f
C1202 B.n402 VSUBS 0.00778f
C1203 B.n403 VSUBS 0.00778f
C1204 B.n404 VSUBS 0.00778f
C1205 B.n405 VSUBS 0.00778f
C1206 B.n406 VSUBS 0.00778f
C1207 B.n407 VSUBS 0.00778f
C1208 B.n408 VSUBS 0.00778f
C1209 B.n409 VSUBS 0.00778f
C1210 B.n410 VSUBS 0.00778f
C1211 B.n411 VSUBS 0.00778f
C1212 B.n412 VSUBS 0.00778f
C1213 B.n413 VSUBS 0.00778f
C1214 B.n414 VSUBS 0.00778f
C1215 B.n415 VSUBS 0.00778f
C1216 B.n416 VSUBS 0.00778f
C1217 B.n417 VSUBS 0.00778f
C1218 B.n418 VSUBS 0.00778f
C1219 B.n419 VSUBS 0.00778f
C1220 B.n420 VSUBS 0.00778f
C1221 B.n421 VSUBS 0.00778f
C1222 B.n422 VSUBS 0.00778f
C1223 B.n423 VSUBS 0.00778f
C1224 B.n424 VSUBS 0.00778f
C1225 B.n425 VSUBS 0.00778f
C1226 B.n426 VSUBS 0.00778f
C1227 B.n427 VSUBS 0.00778f
C1228 B.n428 VSUBS 0.00778f
C1229 B.n429 VSUBS 0.00778f
C1230 B.n430 VSUBS 0.00778f
C1231 B.n431 VSUBS 0.00778f
C1232 B.n432 VSUBS 0.00778f
C1233 B.n433 VSUBS 0.00778f
C1234 B.n434 VSUBS 0.00778f
C1235 B.n435 VSUBS 0.00778f
C1236 B.n436 VSUBS 0.00778f
C1237 B.n437 VSUBS 0.00778f
C1238 B.n438 VSUBS 0.00778f
C1239 B.n439 VSUBS 0.00778f
C1240 B.n440 VSUBS 0.00778f
C1241 B.n441 VSUBS 0.018693f
C1242 B.n442 VSUBS 0.018693f
C1243 B.n443 VSUBS 0.019747f
C1244 B.n444 VSUBS 0.00778f
C1245 B.n445 VSUBS 0.00778f
C1246 B.n446 VSUBS 0.00778f
C1247 B.n447 VSUBS 0.00778f
C1248 B.n448 VSUBS 0.00778f
C1249 B.n449 VSUBS 0.00778f
C1250 B.n450 VSUBS 0.00778f
C1251 B.n451 VSUBS 0.00778f
C1252 B.n452 VSUBS 0.00778f
C1253 B.n453 VSUBS 0.00778f
C1254 B.n454 VSUBS 0.00778f
C1255 B.n455 VSUBS 0.00778f
C1256 B.n456 VSUBS 0.00778f
C1257 B.n457 VSUBS 0.00778f
C1258 B.n458 VSUBS 0.00778f
C1259 B.n459 VSUBS 0.00778f
C1260 B.n460 VSUBS 0.00778f
C1261 B.n461 VSUBS 0.00778f
C1262 B.n462 VSUBS 0.00778f
C1263 B.n463 VSUBS 0.00778f
C1264 B.n464 VSUBS 0.00778f
C1265 B.n465 VSUBS 0.00778f
C1266 B.n466 VSUBS 0.00778f
C1267 B.n467 VSUBS 0.00778f
C1268 B.n468 VSUBS 0.00778f
C1269 B.n469 VSUBS 0.00778f
C1270 B.n470 VSUBS 0.00778f
C1271 B.n471 VSUBS 0.00778f
C1272 B.n472 VSUBS 0.00778f
C1273 B.n473 VSUBS 0.00778f
C1274 B.n474 VSUBS 0.00778f
C1275 B.n475 VSUBS 0.00778f
C1276 B.n476 VSUBS 0.00778f
C1277 B.n477 VSUBS 0.00778f
C1278 B.n478 VSUBS 0.00778f
C1279 B.n479 VSUBS 0.00778f
C1280 B.n480 VSUBS 0.00778f
C1281 B.n481 VSUBS 0.00778f
C1282 B.n482 VSUBS 0.00778f
C1283 B.n483 VSUBS 0.00778f
C1284 B.n484 VSUBS 0.00778f
C1285 B.n485 VSUBS 0.00778f
C1286 B.n486 VSUBS 0.00778f
C1287 B.n487 VSUBS 0.00778f
C1288 B.n488 VSUBS 0.00778f
C1289 B.n489 VSUBS 0.00778f
C1290 B.n490 VSUBS 0.00778f
C1291 B.n491 VSUBS 0.00778f
C1292 B.n492 VSUBS 0.00778f
C1293 B.n493 VSUBS 0.00778f
C1294 B.n494 VSUBS 0.00778f
C1295 B.n495 VSUBS 0.00778f
C1296 B.n496 VSUBS 0.00778f
C1297 B.n497 VSUBS 0.00778f
C1298 B.n498 VSUBS 0.00778f
C1299 B.n499 VSUBS 0.00778f
C1300 B.n500 VSUBS 0.00778f
C1301 B.n501 VSUBS 0.00778f
C1302 B.n502 VSUBS 0.00778f
C1303 B.n503 VSUBS 0.00778f
C1304 B.n504 VSUBS 0.00778f
C1305 B.n505 VSUBS 0.00778f
C1306 B.n506 VSUBS 0.00778f
C1307 B.n507 VSUBS 0.00778f
C1308 B.n508 VSUBS 0.00778f
C1309 B.n509 VSUBS 0.00778f
C1310 B.n510 VSUBS 0.00778f
C1311 B.n511 VSUBS 0.00778f
C1312 B.n512 VSUBS 0.00778f
C1313 B.n513 VSUBS 0.00778f
C1314 B.n514 VSUBS 0.00778f
C1315 B.n515 VSUBS 0.00778f
C1316 B.n516 VSUBS 0.00778f
C1317 B.n517 VSUBS 0.005377f
C1318 B.n518 VSUBS 0.018025f
C1319 B.n519 VSUBS 0.006292f
C1320 B.n520 VSUBS 0.00778f
C1321 B.n521 VSUBS 0.00778f
C1322 B.n522 VSUBS 0.00778f
C1323 B.n523 VSUBS 0.00778f
C1324 B.n524 VSUBS 0.00778f
C1325 B.n525 VSUBS 0.00778f
C1326 B.n526 VSUBS 0.00778f
C1327 B.n527 VSUBS 0.00778f
C1328 B.n528 VSUBS 0.00778f
C1329 B.n529 VSUBS 0.00778f
C1330 B.n530 VSUBS 0.00778f
C1331 B.n531 VSUBS 0.006292f
C1332 B.n532 VSUBS 0.018025f
C1333 B.n533 VSUBS 0.005377f
C1334 B.n534 VSUBS 0.00778f
C1335 B.n535 VSUBS 0.00778f
C1336 B.n536 VSUBS 0.00778f
C1337 B.n537 VSUBS 0.00778f
C1338 B.n538 VSUBS 0.00778f
C1339 B.n539 VSUBS 0.00778f
C1340 B.n540 VSUBS 0.00778f
C1341 B.n541 VSUBS 0.00778f
C1342 B.n542 VSUBS 0.00778f
C1343 B.n543 VSUBS 0.00778f
C1344 B.n544 VSUBS 0.00778f
C1345 B.n545 VSUBS 0.00778f
C1346 B.n546 VSUBS 0.00778f
C1347 B.n547 VSUBS 0.00778f
C1348 B.n548 VSUBS 0.00778f
C1349 B.n549 VSUBS 0.00778f
C1350 B.n550 VSUBS 0.00778f
C1351 B.n551 VSUBS 0.00778f
C1352 B.n552 VSUBS 0.00778f
C1353 B.n553 VSUBS 0.00778f
C1354 B.n554 VSUBS 0.00778f
C1355 B.n555 VSUBS 0.00778f
C1356 B.n556 VSUBS 0.00778f
C1357 B.n557 VSUBS 0.00778f
C1358 B.n558 VSUBS 0.00778f
C1359 B.n559 VSUBS 0.00778f
C1360 B.n560 VSUBS 0.00778f
C1361 B.n561 VSUBS 0.00778f
C1362 B.n562 VSUBS 0.00778f
C1363 B.n563 VSUBS 0.00778f
C1364 B.n564 VSUBS 0.00778f
C1365 B.n565 VSUBS 0.00778f
C1366 B.n566 VSUBS 0.00778f
C1367 B.n567 VSUBS 0.00778f
C1368 B.n568 VSUBS 0.00778f
C1369 B.n569 VSUBS 0.00778f
C1370 B.n570 VSUBS 0.00778f
C1371 B.n571 VSUBS 0.00778f
C1372 B.n572 VSUBS 0.00778f
C1373 B.n573 VSUBS 0.00778f
C1374 B.n574 VSUBS 0.00778f
C1375 B.n575 VSUBS 0.00778f
C1376 B.n576 VSUBS 0.00778f
C1377 B.n577 VSUBS 0.00778f
C1378 B.n578 VSUBS 0.00778f
C1379 B.n579 VSUBS 0.00778f
C1380 B.n580 VSUBS 0.00778f
C1381 B.n581 VSUBS 0.00778f
C1382 B.n582 VSUBS 0.00778f
C1383 B.n583 VSUBS 0.00778f
C1384 B.n584 VSUBS 0.00778f
C1385 B.n585 VSUBS 0.00778f
C1386 B.n586 VSUBS 0.00778f
C1387 B.n587 VSUBS 0.00778f
C1388 B.n588 VSUBS 0.00778f
C1389 B.n589 VSUBS 0.00778f
C1390 B.n590 VSUBS 0.00778f
C1391 B.n591 VSUBS 0.00778f
C1392 B.n592 VSUBS 0.00778f
C1393 B.n593 VSUBS 0.00778f
C1394 B.n594 VSUBS 0.00778f
C1395 B.n595 VSUBS 0.00778f
C1396 B.n596 VSUBS 0.00778f
C1397 B.n597 VSUBS 0.00778f
C1398 B.n598 VSUBS 0.00778f
C1399 B.n599 VSUBS 0.00778f
C1400 B.n600 VSUBS 0.00778f
C1401 B.n601 VSUBS 0.00778f
C1402 B.n602 VSUBS 0.00778f
C1403 B.n603 VSUBS 0.00778f
C1404 B.n604 VSUBS 0.00778f
C1405 B.n605 VSUBS 0.00778f
C1406 B.n606 VSUBS 0.00778f
C1407 B.n607 VSUBS 0.019747f
C1408 B.n608 VSUBS 0.018693f
C1409 B.n609 VSUBS 0.018693f
C1410 B.n610 VSUBS 0.00778f
C1411 B.n611 VSUBS 0.00778f
C1412 B.n612 VSUBS 0.00778f
C1413 B.n613 VSUBS 0.00778f
C1414 B.n614 VSUBS 0.00778f
C1415 B.n615 VSUBS 0.00778f
C1416 B.n616 VSUBS 0.00778f
C1417 B.n617 VSUBS 0.00778f
C1418 B.n618 VSUBS 0.00778f
C1419 B.n619 VSUBS 0.00778f
C1420 B.n620 VSUBS 0.00778f
C1421 B.n621 VSUBS 0.00778f
C1422 B.n622 VSUBS 0.00778f
C1423 B.n623 VSUBS 0.00778f
C1424 B.n624 VSUBS 0.00778f
C1425 B.n625 VSUBS 0.00778f
C1426 B.n626 VSUBS 0.00778f
C1427 B.n627 VSUBS 0.00778f
C1428 B.n628 VSUBS 0.00778f
C1429 B.n629 VSUBS 0.00778f
C1430 B.n630 VSUBS 0.00778f
C1431 B.n631 VSUBS 0.00778f
C1432 B.n632 VSUBS 0.00778f
C1433 B.n633 VSUBS 0.00778f
C1434 B.n634 VSUBS 0.00778f
C1435 B.n635 VSUBS 0.00778f
C1436 B.n636 VSUBS 0.00778f
C1437 B.n637 VSUBS 0.00778f
C1438 B.n638 VSUBS 0.00778f
C1439 B.n639 VSUBS 0.00778f
C1440 B.n640 VSUBS 0.00778f
C1441 B.n641 VSUBS 0.00778f
C1442 B.n642 VSUBS 0.00778f
C1443 B.n643 VSUBS 0.010152f
C1444 B.n644 VSUBS 0.010815f
C1445 B.n645 VSUBS 0.021506f
.ends

