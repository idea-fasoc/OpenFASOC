* NGSPICE file created from diff_pair_sample_0510.ext - technology: sky130A

.subckt diff_pair_sample_0510 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4530_n4070# sky130_fd_pr__pfet_01v8 ad=6.0489 pd=31.8 as=0 ps=0 w=15.51 l=3.23
X1 VDD1.t7 VP.t0 VTAIL.t8 w_n4530_n4070# sky130_fd_pr__pfet_01v8 ad=2.55915 pd=15.84 as=2.55915 ps=15.84 w=15.51 l=3.23
X2 B.t8 B.t6 B.t7 w_n4530_n4070# sky130_fd_pr__pfet_01v8 ad=6.0489 pd=31.8 as=0 ps=0 w=15.51 l=3.23
X3 VTAIL.t3 VN.t0 VDD2.t7 w_n4530_n4070# sky130_fd_pr__pfet_01v8 ad=2.55915 pd=15.84 as=2.55915 ps=15.84 w=15.51 l=3.23
X4 VTAIL.t2 VN.t1 VDD2.t6 w_n4530_n4070# sky130_fd_pr__pfet_01v8 ad=6.0489 pd=31.8 as=2.55915 ps=15.84 w=15.51 l=3.23
X5 VDD1.t6 VP.t1 VTAIL.t9 w_n4530_n4070# sky130_fd_pr__pfet_01v8 ad=2.55915 pd=15.84 as=6.0489 ps=31.8 w=15.51 l=3.23
X6 VTAIL.t6 VN.t2 VDD2.t5 w_n4530_n4070# sky130_fd_pr__pfet_01v8 ad=6.0489 pd=31.8 as=2.55915 ps=15.84 w=15.51 l=3.23
X7 VDD2.t4 VN.t3 VTAIL.t1 w_n4530_n4070# sky130_fd_pr__pfet_01v8 ad=2.55915 pd=15.84 as=6.0489 ps=31.8 w=15.51 l=3.23
X8 VTAIL.t7 VN.t4 VDD2.t3 w_n4530_n4070# sky130_fd_pr__pfet_01v8 ad=2.55915 pd=15.84 as=2.55915 ps=15.84 w=15.51 l=3.23
X9 VDD1.t5 VP.t2 VTAIL.t10 w_n4530_n4070# sky130_fd_pr__pfet_01v8 ad=2.55915 pd=15.84 as=6.0489 ps=31.8 w=15.51 l=3.23
X10 VTAIL.t11 VP.t3 VDD1.t4 w_n4530_n4070# sky130_fd_pr__pfet_01v8 ad=2.55915 pd=15.84 as=2.55915 ps=15.84 w=15.51 l=3.23
X11 VDD1.t3 VP.t4 VTAIL.t12 w_n4530_n4070# sky130_fd_pr__pfet_01v8 ad=2.55915 pd=15.84 as=2.55915 ps=15.84 w=15.51 l=3.23
X12 VTAIL.t13 VP.t5 VDD1.t2 w_n4530_n4070# sky130_fd_pr__pfet_01v8 ad=6.0489 pd=31.8 as=2.55915 ps=15.84 w=15.51 l=3.23
X13 VDD2.t2 VN.t5 VTAIL.t0 w_n4530_n4070# sky130_fd_pr__pfet_01v8 ad=2.55915 pd=15.84 as=2.55915 ps=15.84 w=15.51 l=3.23
X14 VTAIL.t14 VP.t6 VDD1.t1 w_n4530_n4070# sky130_fd_pr__pfet_01v8 ad=6.0489 pd=31.8 as=2.55915 ps=15.84 w=15.51 l=3.23
X15 VDD2.t1 VN.t6 VTAIL.t5 w_n4530_n4070# sky130_fd_pr__pfet_01v8 ad=2.55915 pd=15.84 as=2.55915 ps=15.84 w=15.51 l=3.23
X16 VDD2.t0 VN.t7 VTAIL.t4 w_n4530_n4070# sky130_fd_pr__pfet_01v8 ad=2.55915 pd=15.84 as=6.0489 ps=31.8 w=15.51 l=3.23
X17 B.t5 B.t3 B.t4 w_n4530_n4070# sky130_fd_pr__pfet_01v8 ad=6.0489 pd=31.8 as=0 ps=0 w=15.51 l=3.23
X18 VTAIL.t15 VP.t7 VDD1.t0 w_n4530_n4070# sky130_fd_pr__pfet_01v8 ad=2.55915 pd=15.84 as=2.55915 ps=15.84 w=15.51 l=3.23
X19 B.t2 B.t0 B.t1 w_n4530_n4070# sky130_fd_pr__pfet_01v8 ad=6.0489 pd=31.8 as=0 ps=0 w=15.51 l=3.23
R0 B.n503 B.n154 585
R1 B.n502 B.n501 585
R2 B.n500 B.n155 585
R3 B.n499 B.n498 585
R4 B.n497 B.n156 585
R5 B.n496 B.n495 585
R6 B.n494 B.n157 585
R7 B.n493 B.n492 585
R8 B.n491 B.n158 585
R9 B.n490 B.n489 585
R10 B.n488 B.n159 585
R11 B.n487 B.n486 585
R12 B.n485 B.n160 585
R13 B.n484 B.n483 585
R14 B.n482 B.n161 585
R15 B.n481 B.n480 585
R16 B.n479 B.n162 585
R17 B.n478 B.n477 585
R18 B.n476 B.n163 585
R19 B.n475 B.n474 585
R20 B.n473 B.n164 585
R21 B.n472 B.n471 585
R22 B.n470 B.n165 585
R23 B.n469 B.n468 585
R24 B.n467 B.n166 585
R25 B.n466 B.n465 585
R26 B.n464 B.n167 585
R27 B.n463 B.n462 585
R28 B.n461 B.n168 585
R29 B.n460 B.n459 585
R30 B.n458 B.n169 585
R31 B.n457 B.n456 585
R32 B.n455 B.n170 585
R33 B.n454 B.n453 585
R34 B.n452 B.n171 585
R35 B.n451 B.n450 585
R36 B.n449 B.n172 585
R37 B.n448 B.n447 585
R38 B.n446 B.n173 585
R39 B.n445 B.n444 585
R40 B.n443 B.n174 585
R41 B.n442 B.n441 585
R42 B.n440 B.n175 585
R43 B.n439 B.n438 585
R44 B.n437 B.n176 585
R45 B.n436 B.n435 585
R46 B.n434 B.n177 585
R47 B.n433 B.n432 585
R48 B.n431 B.n178 585
R49 B.n430 B.n429 585
R50 B.n428 B.n179 585
R51 B.n427 B.n426 585
R52 B.n425 B.n424 585
R53 B.n423 B.n183 585
R54 B.n422 B.n421 585
R55 B.n420 B.n184 585
R56 B.n419 B.n418 585
R57 B.n417 B.n185 585
R58 B.n416 B.n415 585
R59 B.n414 B.n186 585
R60 B.n413 B.n412 585
R61 B.n410 B.n187 585
R62 B.n409 B.n408 585
R63 B.n407 B.n190 585
R64 B.n406 B.n405 585
R65 B.n404 B.n191 585
R66 B.n403 B.n402 585
R67 B.n401 B.n192 585
R68 B.n400 B.n399 585
R69 B.n398 B.n193 585
R70 B.n397 B.n396 585
R71 B.n395 B.n194 585
R72 B.n394 B.n393 585
R73 B.n392 B.n195 585
R74 B.n391 B.n390 585
R75 B.n389 B.n196 585
R76 B.n388 B.n387 585
R77 B.n386 B.n197 585
R78 B.n385 B.n384 585
R79 B.n383 B.n198 585
R80 B.n382 B.n381 585
R81 B.n380 B.n199 585
R82 B.n379 B.n378 585
R83 B.n377 B.n200 585
R84 B.n376 B.n375 585
R85 B.n374 B.n201 585
R86 B.n373 B.n372 585
R87 B.n371 B.n202 585
R88 B.n370 B.n369 585
R89 B.n368 B.n203 585
R90 B.n367 B.n366 585
R91 B.n365 B.n204 585
R92 B.n364 B.n363 585
R93 B.n362 B.n205 585
R94 B.n361 B.n360 585
R95 B.n359 B.n206 585
R96 B.n358 B.n357 585
R97 B.n356 B.n207 585
R98 B.n355 B.n354 585
R99 B.n353 B.n208 585
R100 B.n352 B.n351 585
R101 B.n350 B.n209 585
R102 B.n349 B.n348 585
R103 B.n347 B.n210 585
R104 B.n346 B.n345 585
R105 B.n344 B.n211 585
R106 B.n343 B.n342 585
R107 B.n341 B.n212 585
R108 B.n340 B.n339 585
R109 B.n338 B.n213 585
R110 B.n337 B.n336 585
R111 B.n335 B.n214 585
R112 B.n334 B.n333 585
R113 B.n505 B.n504 585
R114 B.n506 B.n153 585
R115 B.n508 B.n507 585
R116 B.n509 B.n152 585
R117 B.n511 B.n510 585
R118 B.n512 B.n151 585
R119 B.n514 B.n513 585
R120 B.n515 B.n150 585
R121 B.n517 B.n516 585
R122 B.n518 B.n149 585
R123 B.n520 B.n519 585
R124 B.n521 B.n148 585
R125 B.n523 B.n522 585
R126 B.n524 B.n147 585
R127 B.n526 B.n525 585
R128 B.n527 B.n146 585
R129 B.n529 B.n528 585
R130 B.n530 B.n145 585
R131 B.n532 B.n531 585
R132 B.n533 B.n144 585
R133 B.n535 B.n534 585
R134 B.n536 B.n143 585
R135 B.n538 B.n537 585
R136 B.n539 B.n142 585
R137 B.n541 B.n540 585
R138 B.n542 B.n141 585
R139 B.n544 B.n543 585
R140 B.n545 B.n140 585
R141 B.n547 B.n546 585
R142 B.n548 B.n139 585
R143 B.n550 B.n549 585
R144 B.n551 B.n138 585
R145 B.n553 B.n552 585
R146 B.n554 B.n137 585
R147 B.n556 B.n555 585
R148 B.n557 B.n136 585
R149 B.n559 B.n558 585
R150 B.n560 B.n135 585
R151 B.n562 B.n561 585
R152 B.n563 B.n134 585
R153 B.n565 B.n564 585
R154 B.n566 B.n133 585
R155 B.n568 B.n567 585
R156 B.n569 B.n132 585
R157 B.n571 B.n570 585
R158 B.n572 B.n131 585
R159 B.n574 B.n573 585
R160 B.n575 B.n130 585
R161 B.n577 B.n576 585
R162 B.n578 B.n129 585
R163 B.n580 B.n579 585
R164 B.n581 B.n128 585
R165 B.n583 B.n582 585
R166 B.n584 B.n127 585
R167 B.n586 B.n585 585
R168 B.n587 B.n126 585
R169 B.n589 B.n588 585
R170 B.n590 B.n125 585
R171 B.n592 B.n591 585
R172 B.n593 B.n124 585
R173 B.n595 B.n594 585
R174 B.n596 B.n123 585
R175 B.n598 B.n597 585
R176 B.n599 B.n122 585
R177 B.n601 B.n600 585
R178 B.n602 B.n121 585
R179 B.n604 B.n603 585
R180 B.n605 B.n120 585
R181 B.n607 B.n606 585
R182 B.n608 B.n119 585
R183 B.n610 B.n609 585
R184 B.n611 B.n118 585
R185 B.n613 B.n612 585
R186 B.n614 B.n117 585
R187 B.n616 B.n615 585
R188 B.n617 B.n116 585
R189 B.n619 B.n618 585
R190 B.n620 B.n115 585
R191 B.n622 B.n621 585
R192 B.n623 B.n114 585
R193 B.n625 B.n624 585
R194 B.n626 B.n113 585
R195 B.n628 B.n627 585
R196 B.n629 B.n112 585
R197 B.n631 B.n630 585
R198 B.n632 B.n111 585
R199 B.n634 B.n633 585
R200 B.n635 B.n110 585
R201 B.n637 B.n636 585
R202 B.n638 B.n109 585
R203 B.n640 B.n639 585
R204 B.n641 B.n108 585
R205 B.n643 B.n642 585
R206 B.n644 B.n107 585
R207 B.n646 B.n645 585
R208 B.n647 B.n106 585
R209 B.n649 B.n648 585
R210 B.n650 B.n105 585
R211 B.n652 B.n651 585
R212 B.n653 B.n104 585
R213 B.n655 B.n654 585
R214 B.n656 B.n103 585
R215 B.n658 B.n657 585
R216 B.n659 B.n102 585
R217 B.n661 B.n660 585
R218 B.n662 B.n101 585
R219 B.n664 B.n663 585
R220 B.n665 B.n100 585
R221 B.n667 B.n666 585
R222 B.n668 B.n99 585
R223 B.n670 B.n669 585
R224 B.n671 B.n98 585
R225 B.n673 B.n672 585
R226 B.n674 B.n97 585
R227 B.n676 B.n675 585
R228 B.n677 B.n96 585
R229 B.n679 B.n678 585
R230 B.n680 B.n95 585
R231 B.n682 B.n681 585
R232 B.n683 B.n94 585
R233 B.n685 B.n684 585
R234 B.n686 B.n93 585
R235 B.n857 B.n32 585
R236 B.n856 B.n855 585
R237 B.n854 B.n33 585
R238 B.n853 B.n852 585
R239 B.n851 B.n34 585
R240 B.n850 B.n849 585
R241 B.n848 B.n35 585
R242 B.n847 B.n846 585
R243 B.n845 B.n36 585
R244 B.n844 B.n843 585
R245 B.n842 B.n37 585
R246 B.n841 B.n840 585
R247 B.n839 B.n38 585
R248 B.n838 B.n837 585
R249 B.n836 B.n39 585
R250 B.n835 B.n834 585
R251 B.n833 B.n40 585
R252 B.n832 B.n831 585
R253 B.n830 B.n41 585
R254 B.n829 B.n828 585
R255 B.n827 B.n42 585
R256 B.n826 B.n825 585
R257 B.n824 B.n43 585
R258 B.n823 B.n822 585
R259 B.n821 B.n44 585
R260 B.n820 B.n819 585
R261 B.n818 B.n45 585
R262 B.n817 B.n816 585
R263 B.n815 B.n46 585
R264 B.n814 B.n813 585
R265 B.n812 B.n47 585
R266 B.n811 B.n810 585
R267 B.n809 B.n48 585
R268 B.n808 B.n807 585
R269 B.n806 B.n49 585
R270 B.n805 B.n804 585
R271 B.n803 B.n50 585
R272 B.n802 B.n801 585
R273 B.n800 B.n51 585
R274 B.n799 B.n798 585
R275 B.n797 B.n52 585
R276 B.n796 B.n795 585
R277 B.n794 B.n53 585
R278 B.n793 B.n792 585
R279 B.n791 B.n54 585
R280 B.n790 B.n789 585
R281 B.n788 B.n55 585
R282 B.n787 B.n786 585
R283 B.n785 B.n56 585
R284 B.n784 B.n783 585
R285 B.n782 B.n57 585
R286 B.n781 B.n780 585
R287 B.n779 B.n778 585
R288 B.n777 B.n61 585
R289 B.n776 B.n775 585
R290 B.n774 B.n62 585
R291 B.n773 B.n772 585
R292 B.n771 B.n63 585
R293 B.n770 B.n769 585
R294 B.n768 B.n64 585
R295 B.n767 B.n766 585
R296 B.n764 B.n65 585
R297 B.n763 B.n762 585
R298 B.n761 B.n68 585
R299 B.n760 B.n759 585
R300 B.n758 B.n69 585
R301 B.n757 B.n756 585
R302 B.n755 B.n70 585
R303 B.n754 B.n753 585
R304 B.n752 B.n71 585
R305 B.n751 B.n750 585
R306 B.n749 B.n72 585
R307 B.n748 B.n747 585
R308 B.n746 B.n73 585
R309 B.n745 B.n744 585
R310 B.n743 B.n74 585
R311 B.n742 B.n741 585
R312 B.n740 B.n75 585
R313 B.n739 B.n738 585
R314 B.n737 B.n76 585
R315 B.n736 B.n735 585
R316 B.n734 B.n77 585
R317 B.n733 B.n732 585
R318 B.n731 B.n78 585
R319 B.n730 B.n729 585
R320 B.n728 B.n79 585
R321 B.n727 B.n726 585
R322 B.n725 B.n80 585
R323 B.n724 B.n723 585
R324 B.n722 B.n81 585
R325 B.n721 B.n720 585
R326 B.n719 B.n82 585
R327 B.n718 B.n717 585
R328 B.n716 B.n83 585
R329 B.n715 B.n714 585
R330 B.n713 B.n84 585
R331 B.n712 B.n711 585
R332 B.n710 B.n85 585
R333 B.n709 B.n708 585
R334 B.n707 B.n86 585
R335 B.n706 B.n705 585
R336 B.n704 B.n87 585
R337 B.n703 B.n702 585
R338 B.n701 B.n88 585
R339 B.n700 B.n699 585
R340 B.n698 B.n89 585
R341 B.n697 B.n696 585
R342 B.n695 B.n90 585
R343 B.n694 B.n693 585
R344 B.n692 B.n91 585
R345 B.n691 B.n690 585
R346 B.n689 B.n92 585
R347 B.n688 B.n687 585
R348 B.n859 B.n858 585
R349 B.n860 B.n31 585
R350 B.n862 B.n861 585
R351 B.n863 B.n30 585
R352 B.n865 B.n864 585
R353 B.n866 B.n29 585
R354 B.n868 B.n867 585
R355 B.n869 B.n28 585
R356 B.n871 B.n870 585
R357 B.n872 B.n27 585
R358 B.n874 B.n873 585
R359 B.n875 B.n26 585
R360 B.n877 B.n876 585
R361 B.n878 B.n25 585
R362 B.n880 B.n879 585
R363 B.n881 B.n24 585
R364 B.n883 B.n882 585
R365 B.n884 B.n23 585
R366 B.n886 B.n885 585
R367 B.n887 B.n22 585
R368 B.n889 B.n888 585
R369 B.n890 B.n21 585
R370 B.n892 B.n891 585
R371 B.n893 B.n20 585
R372 B.n895 B.n894 585
R373 B.n896 B.n19 585
R374 B.n898 B.n897 585
R375 B.n899 B.n18 585
R376 B.n901 B.n900 585
R377 B.n902 B.n17 585
R378 B.n904 B.n903 585
R379 B.n905 B.n16 585
R380 B.n907 B.n906 585
R381 B.n908 B.n15 585
R382 B.n910 B.n909 585
R383 B.n911 B.n14 585
R384 B.n913 B.n912 585
R385 B.n914 B.n13 585
R386 B.n916 B.n915 585
R387 B.n917 B.n12 585
R388 B.n919 B.n918 585
R389 B.n920 B.n11 585
R390 B.n922 B.n921 585
R391 B.n923 B.n10 585
R392 B.n925 B.n924 585
R393 B.n926 B.n9 585
R394 B.n928 B.n927 585
R395 B.n929 B.n8 585
R396 B.n931 B.n930 585
R397 B.n932 B.n7 585
R398 B.n934 B.n933 585
R399 B.n935 B.n6 585
R400 B.n937 B.n936 585
R401 B.n938 B.n5 585
R402 B.n940 B.n939 585
R403 B.n941 B.n4 585
R404 B.n943 B.n942 585
R405 B.n944 B.n3 585
R406 B.n946 B.n945 585
R407 B.n947 B.n0 585
R408 B.n2 B.n1 585
R409 B.n245 B.n244 585
R410 B.n247 B.n246 585
R411 B.n248 B.n243 585
R412 B.n250 B.n249 585
R413 B.n251 B.n242 585
R414 B.n253 B.n252 585
R415 B.n254 B.n241 585
R416 B.n256 B.n255 585
R417 B.n257 B.n240 585
R418 B.n259 B.n258 585
R419 B.n260 B.n239 585
R420 B.n262 B.n261 585
R421 B.n263 B.n238 585
R422 B.n265 B.n264 585
R423 B.n266 B.n237 585
R424 B.n268 B.n267 585
R425 B.n269 B.n236 585
R426 B.n271 B.n270 585
R427 B.n272 B.n235 585
R428 B.n274 B.n273 585
R429 B.n275 B.n234 585
R430 B.n277 B.n276 585
R431 B.n278 B.n233 585
R432 B.n280 B.n279 585
R433 B.n281 B.n232 585
R434 B.n283 B.n282 585
R435 B.n284 B.n231 585
R436 B.n286 B.n285 585
R437 B.n287 B.n230 585
R438 B.n289 B.n288 585
R439 B.n290 B.n229 585
R440 B.n292 B.n291 585
R441 B.n293 B.n228 585
R442 B.n295 B.n294 585
R443 B.n296 B.n227 585
R444 B.n298 B.n297 585
R445 B.n299 B.n226 585
R446 B.n301 B.n300 585
R447 B.n302 B.n225 585
R448 B.n304 B.n303 585
R449 B.n305 B.n224 585
R450 B.n307 B.n306 585
R451 B.n308 B.n223 585
R452 B.n310 B.n309 585
R453 B.n311 B.n222 585
R454 B.n313 B.n312 585
R455 B.n314 B.n221 585
R456 B.n316 B.n315 585
R457 B.n317 B.n220 585
R458 B.n319 B.n318 585
R459 B.n320 B.n219 585
R460 B.n322 B.n321 585
R461 B.n323 B.n218 585
R462 B.n325 B.n324 585
R463 B.n326 B.n217 585
R464 B.n328 B.n327 585
R465 B.n329 B.n216 585
R466 B.n331 B.n330 585
R467 B.n332 B.n215 585
R468 B.n334 B.n215 530.939
R469 B.n504 B.n503 530.939
R470 B.n688 B.n93 530.939
R471 B.n858 B.n857 530.939
R472 B.n180 B.t10 507.945
R473 B.n66 B.t8 507.945
R474 B.n188 B.t4 507.945
R475 B.n58 B.t2 507.945
R476 B.n181 B.t11 438.901
R477 B.n67 B.t7 438.901
R478 B.n189 B.t5 438.901
R479 B.n59 B.t1 438.901
R480 B.n188 B.t3 324.558
R481 B.n180 B.t9 324.558
R482 B.n66 B.t6 324.558
R483 B.n58 B.t0 324.558
R484 B.n949 B.n948 256.663
R485 B.n948 B.n947 235.042
R486 B.n948 B.n2 235.042
R487 B.n335 B.n334 163.367
R488 B.n336 B.n335 163.367
R489 B.n336 B.n213 163.367
R490 B.n340 B.n213 163.367
R491 B.n341 B.n340 163.367
R492 B.n342 B.n341 163.367
R493 B.n342 B.n211 163.367
R494 B.n346 B.n211 163.367
R495 B.n347 B.n346 163.367
R496 B.n348 B.n347 163.367
R497 B.n348 B.n209 163.367
R498 B.n352 B.n209 163.367
R499 B.n353 B.n352 163.367
R500 B.n354 B.n353 163.367
R501 B.n354 B.n207 163.367
R502 B.n358 B.n207 163.367
R503 B.n359 B.n358 163.367
R504 B.n360 B.n359 163.367
R505 B.n360 B.n205 163.367
R506 B.n364 B.n205 163.367
R507 B.n365 B.n364 163.367
R508 B.n366 B.n365 163.367
R509 B.n366 B.n203 163.367
R510 B.n370 B.n203 163.367
R511 B.n371 B.n370 163.367
R512 B.n372 B.n371 163.367
R513 B.n372 B.n201 163.367
R514 B.n376 B.n201 163.367
R515 B.n377 B.n376 163.367
R516 B.n378 B.n377 163.367
R517 B.n378 B.n199 163.367
R518 B.n382 B.n199 163.367
R519 B.n383 B.n382 163.367
R520 B.n384 B.n383 163.367
R521 B.n384 B.n197 163.367
R522 B.n388 B.n197 163.367
R523 B.n389 B.n388 163.367
R524 B.n390 B.n389 163.367
R525 B.n390 B.n195 163.367
R526 B.n394 B.n195 163.367
R527 B.n395 B.n394 163.367
R528 B.n396 B.n395 163.367
R529 B.n396 B.n193 163.367
R530 B.n400 B.n193 163.367
R531 B.n401 B.n400 163.367
R532 B.n402 B.n401 163.367
R533 B.n402 B.n191 163.367
R534 B.n406 B.n191 163.367
R535 B.n407 B.n406 163.367
R536 B.n408 B.n407 163.367
R537 B.n408 B.n187 163.367
R538 B.n413 B.n187 163.367
R539 B.n414 B.n413 163.367
R540 B.n415 B.n414 163.367
R541 B.n415 B.n185 163.367
R542 B.n419 B.n185 163.367
R543 B.n420 B.n419 163.367
R544 B.n421 B.n420 163.367
R545 B.n421 B.n183 163.367
R546 B.n425 B.n183 163.367
R547 B.n426 B.n425 163.367
R548 B.n426 B.n179 163.367
R549 B.n430 B.n179 163.367
R550 B.n431 B.n430 163.367
R551 B.n432 B.n431 163.367
R552 B.n432 B.n177 163.367
R553 B.n436 B.n177 163.367
R554 B.n437 B.n436 163.367
R555 B.n438 B.n437 163.367
R556 B.n438 B.n175 163.367
R557 B.n442 B.n175 163.367
R558 B.n443 B.n442 163.367
R559 B.n444 B.n443 163.367
R560 B.n444 B.n173 163.367
R561 B.n448 B.n173 163.367
R562 B.n449 B.n448 163.367
R563 B.n450 B.n449 163.367
R564 B.n450 B.n171 163.367
R565 B.n454 B.n171 163.367
R566 B.n455 B.n454 163.367
R567 B.n456 B.n455 163.367
R568 B.n456 B.n169 163.367
R569 B.n460 B.n169 163.367
R570 B.n461 B.n460 163.367
R571 B.n462 B.n461 163.367
R572 B.n462 B.n167 163.367
R573 B.n466 B.n167 163.367
R574 B.n467 B.n466 163.367
R575 B.n468 B.n467 163.367
R576 B.n468 B.n165 163.367
R577 B.n472 B.n165 163.367
R578 B.n473 B.n472 163.367
R579 B.n474 B.n473 163.367
R580 B.n474 B.n163 163.367
R581 B.n478 B.n163 163.367
R582 B.n479 B.n478 163.367
R583 B.n480 B.n479 163.367
R584 B.n480 B.n161 163.367
R585 B.n484 B.n161 163.367
R586 B.n485 B.n484 163.367
R587 B.n486 B.n485 163.367
R588 B.n486 B.n159 163.367
R589 B.n490 B.n159 163.367
R590 B.n491 B.n490 163.367
R591 B.n492 B.n491 163.367
R592 B.n492 B.n157 163.367
R593 B.n496 B.n157 163.367
R594 B.n497 B.n496 163.367
R595 B.n498 B.n497 163.367
R596 B.n498 B.n155 163.367
R597 B.n502 B.n155 163.367
R598 B.n503 B.n502 163.367
R599 B.n684 B.n93 163.367
R600 B.n684 B.n683 163.367
R601 B.n683 B.n682 163.367
R602 B.n682 B.n95 163.367
R603 B.n678 B.n95 163.367
R604 B.n678 B.n677 163.367
R605 B.n677 B.n676 163.367
R606 B.n676 B.n97 163.367
R607 B.n672 B.n97 163.367
R608 B.n672 B.n671 163.367
R609 B.n671 B.n670 163.367
R610 B.n670 B.n99 163.367
R611 B.n666 B.n99 163.367
R612 B.n666 B.n665 163.367
R613 B.n665 B.n664 163.367
R614 B.n664 B.n101 163.367
R615 B.n660 B.n101 163.367
R616 B.n660 B.n659 163.367
R617 B.n659 B.n658 163.367
R618 B.n658 B.n103 163.367
R619 B.n654 B.n103 163.367
R620 B.n654 B.n653 163.367
R621 B.n653 B.n652 163.367
R622 B.n652 B.n105 163.367
R623 B.n648 B.n105 163.367
R624 B.n648 B.n647 163.367
R625 B.n647 B.n646 163.367
R626 B.n646 B.n107 163.367
R627 B.n642 B.n107 163.367
R628 B.n642 B.n641 163.367
R629 B.n641 B.n640 163.367
R630 B.n640 B.n109 163.367
R631 B.n636 B.n109 163.367
R632 B.n636 B.n635 163.367
R633 B.n635 B.n634 163.367
R634 B.n634 B.n111 163.367
R635 B.n630 B.n111 163.367
R636 B.n630 B.n629 163.367
R637 B.n629 B.n628 163.367
R638 B.n628 B.n113 163.367
R639 B.n624 B.n113 163.367
R640 B.n624 B.n623 163.367
R641 B.n623 B.n622 163.367
R642 B.n622 B.n115 163.367
R643 B.n618 B.n115 163.367
R644 B.n618 B.n617 163.367
R645 B.n617 B.n616 163.367
R646 B.n616 B.n117 163.367
R647 B.n612 B.n117 163.367
R648 B.n612 B.n611 163.367
R649 B.n611 B.n610 163.367
R650 B.n610 B.n119 163.367
R651 B.n606 B.n119 163.367
R652 B.n606 B.n605 163.367
R653 B.n605 B.n604 163.367
R654 B.n604 B.n121 163.367
R655 B.n600 B.n121 163.367
R656 B.n600 B.n599 163.367
R657 B.n599 B.n598 163.367
R658 B.n598 B.n123 163.367
R659 B.n594 B.n123 163.367
R660 B.n594 B.n593 163.367
R661 B.n593 B.n592 163.367
R662 B.n592 B.n125 163.367
R663 B.n588 B.n125 163.367
R664 B.n588 B.n587 163.367
R665 B.n587 B.n586 163.367
R666 B.n586 B.n127 163.367
R667 B.n582 B.n127 163.367
R668 B.n582 B.n581 163.367
R669 B.n581 B.n580 163.367
R670 B.n580 B.n129 163.367
R671 B.n576 B.n129 163.367
R672 B.n576 B.n575 163.367
R673 B.n575 B.n574 163.367
R674 B.n574 B.n131 163.367
R675 B.n570 B.n131 163.367
R676 B.n570 B.n569 163.367
R677 B.n569 B.n568 163.367
R678 B.n568 B.n133 163.367
R679 B.n564 B.n133 163.367
R680 B.n564 B.n563 163.367
R681 B.n563 B.n562 163.367
R682 B.n562 B.n135 163.367
R683 B.n558 B.n135 163.367
R684 B.n558 B.n557 163.367
R685 B.n557 B.n556 163.367
R686 B.n556 B.n137 163.367
R687 B.n552 B.n137 163.367
R688 B.n552 B.n551 163.367
R689 B.n551 B.n550 163.367
R690 B.n550 B.n139 163.367
R691 B.n546 B.n139 163.367
R692 B.n546 B.n545 163.367
R693 B.n545 B.n544 163.367
R694 B.n544 B.n141 163.367
R695 B.n540 B.n141 163.367
R696 B.n540 B.n539 163.367
R697 B.n539 B.n538 163.367
R698 B.n538 B.n143 163.367
R699 B.n534 B.n143 163.367
R700 B.n534 B.n533 163.367
R701 B.n533 B.n532 163.367
R702 B.n532 B.n145 163.367
R703 B.n528 B.n145 163.367
R704 B.n528 B.n527 163.367
R705 B.n527 B.n526 163.367
R706 B.n526 B.n147 163.367
R707 B.n522 B.n147 163.367
R708 B.n522 B.n521 163.367
R709 B.n521 B.n520 163.367
R710 B.n520 B.n149 163.367
R711 B.n516 B.n149 163.367
R712 B.n516 B.n515 163.367
R713 B.n515 B.n514 163.367
R714 B.n514 B.n151 163.367
R715 B.n510 B.n151 163.367
R716 B.n510 B.n509 163.367
R717 B.n509 B.n508 163.367
R718 B.n508 B.n153 163.367
R719 B.n504 B.n153 163.367
R720 B.n857 B.n856 163.367
R721 B.n856 B.n33 163.367
R722 B.n852 B.n33 163.367
R723 B.n852 B.n851 163.367
R724 B.n851 B.n850 163.367
R725 B.n850 B.n35 163.367
R726 B.n846 B.n35 163.367
R727 B.n846 B.n845 163.367
R728 B.n845 B.n844 163.367
R729 B.n844 B.n37 163.367
R730 B.n840 B.n37 163.367
R731 B.n840 B.n839 163.367
R732 B.n839 B.n838 163.367
R733 B.n838 B.n39 163.367
R734 B.n834 B.n39 163.367
R735 B.n834 B.n833 163.367
R736 B.n833 B.n832 163.367
R737 B.n832 B.n41 163.367
R738 B.n828 B.n41 163.367
R739 B.n828 B.n827 163.367
R740 B.n827 B.n826 163.367
R741 B.n826 B.n43 163.367
R742 B.n822 B.n43 163.367
R743 B.n822 B.n821 163.367
R744 B.n821 B.n820 163.367
R745 B.n820 B.n45 163.367
R746 B.n816 B.n45 163.367
R747 B.n816 B.n815 163.367
R748 B.n815 B.n814 163.367
R749 B.n814 B.n47 163.367
R750 B.n810 B.n47 163.367
R751 B.n810 B.n809 163.367
R752 B.n809 B.n808 163.367
R753 B.n808 B.n49 163.367
R754 B.n804 B.n49 163.367
R755 B.n804 B.n803 163.367
R756 B.n803 B.n802 163.367
R757 B.n802 B.n51 163.367
R758 B.n798 B.n51 163.367
R759 B.n798 B.n797 163.367
R760 B.n797 B.n796 163.367
R761 B.n796 B.n53 163.367
R762 B.n792 B.n53 163.367
R763 B.n792 B.n791 163.367
R764 B.n791 B.n790 163.367
R765 B.n790 B.n55 163.367
R766 B.n786 B.n55 163.367
R767 B.n786 B.n785 163.367
R768 B.n785 B.n784 163.367
R769 B.n784 B.n57 163.367
R770 B.n780 B.n57 163.367
R771 B.n780 B.n779 163.367
R772 B.n779 B.n61 163.367
R773 B.n775 B.n61 163.367
R774 B.n775 B.n774 163.367
R775 B.n774 B.n773 163.367
R776 B.n773 B.n63 163.367
R777 B.n769 B.n63 163.367
R778 B.n769 B.n768 163.367
R779 B.n768 B.n767 163.367
R780 B.n767 B.n65 163.367
R781 B.n762 B.n65 163.367
R782 B.n762 B.n761 163.367
R783 B.n761 B.n760 163.367
R784 B.n760 B.n69 163.367
R785 B.n756 B.n69 163.367
R786 B.n756 B.n755 163.367
R787 B.n755 B.n754 163.367
R788 B.n754 B.n71 163.367
R789 B.n750 B.n71 163.367
R790 B.n750 B.n749 163.367
R791 B.n749 B.n748 163.367
R792 B.n748 B.n73 163.367
R793 B.n744 B.n73 163.367
R794 B.n744 B.n743 163.367
R795 B.n743 B.n742 163.367
R796 B.n742 B.n75 163.367
R797 B.n738 B.n75 163.367
R798 B.n738 B.n737 163.367
R799 B.n737 B.n736 163.367
R800 B.n736 B.n77 163.367
R801 B.n732 B.n77 163.367
R802 B.n732 B.n731 163.367
R803 B.n731 B.n730 163.367
R804 B.n730 B.n79 163.367
R805 B.n726 B.n79 163.367
R806 B.n726 B.n725 163.367
R807 B.n725 B.n724 163.367
R808 B.n724 B.n81 163.367
R809 B.n720 B.n81 163.367
R810 B.n720 B.n719 163.367
R811 B.n719 B.n718 163.367
R812 B.n718 B.n83 163.367
R813 B.n714 B.n83 163.367
R814 B.n714 B.n713 163.367
R815 B.n713 B.n712 163.367
R816 B.n712 B.n85 163.367
R817 B.n708 B.n85 163.367
R818 B.n708 B.n707 163.367
R819 B.n707 B.n706 163.367
R820 B.n706 B.n87 163.367
R821 B.n702 B.n87 163.367
R822 B.n702 B.n701 163.367
R823 B.n701 B.n700 163.367
R824 B.n700 B.n89 163.367
R825 B.n696 B.n89 163.367
R826 B.n696 B.n695 163.367
R827 B.n695 B.n694 163.367
R828 B.n694 B.n91 163.367
R829 B.n690 B.n91 163.367
R830 B.n690 B.n689 163.367
R831 B.n689 B.n688 163.367
R832 B.n858 B.n31 163.367
R833 B.n862 B.n31 163.367
R834 B.n863 B.n862 163.367
R835 B.n864 B.n863 163.367
R836 B.n864 B.n29 163.367
R837 B.n868 B.n29 163.367
R838 B.n869 B.n868 163.367
R839 B.n870 B.n869 163.367
R840 B.n870 B.n27 163.367
R841 B.n874 B.n27 163.367
R842 B.n875 B.n874 163.367
R843 B.n876 B.n875 163.367
R844 B.n876 B.n25 163.367
R845 B.n880 B.n25 163.367
R846 B.n881 B.n880 163.367
R847 B.n882 B.n881 163.367
R848 B.n882 B.n23 163.367
R849 B.n886 B.n23 163.367
R850 B.n887 B.n886 163.367
R851 B.n888 B.n887 163.367
R852 B.n888 B.n21 163.367
R853 B.n892 B.n21 163.367
R854 B.n893 B.n892 163.367
R855 B.n894 B.n893 163.367
R856 B.n894 B.n19 163.367
R857 B.n898 B.n19 163.367
R858 B.n899 B.n898 163.367
R859 B.n900 B.n899 163.367
R860 B.n900 B.n17 163.367
R861 B.n904 B.n17 163.367
R862 B.n905 B.n904 163.367
R863 B.n906 B.n905 163.367
R864 B.n906 B.n15 163.367
R865 B.n910 B.n15 163.367
R866 B.n911 B.n910 163.367
R867 B.n912 B.n911 163.367
R868 B.n912 B.n13 163.367
R869 B.n916 B.n13 163.367
R870 B.n917 B.n916 163.367
R871 B.n918 B.n917 163.367
R872 B.n918 B.n11 163.367
R873 B.n922 B.n11 163.367
R874 B.n923 B.n922 163.367
R875 B.n924 B.n923 163.367
R876 B.n924 B.n9 163.367
R877 B.n928 B.n9 163.367
R878 B.n929 B.n928 163.367
R879 B.n930 B.n929 163.367
R880 B.n930 B.n7 163.367
R881 B.n934 B.n7 163.367
R882 B.n935 B.n934 163.367
R883 B.n936 B.n935 163.367
R884 B.n936 B.n5 163.367
R885 B.n940 B.n5 163.367
R886 B.n941 B.n940 163.367
R887 B.n942 B.n941 163.367
R888 B.n942 B.n3 163.367
R889 B.n946 B.n3 163.367
R890 B.n947 B.n946 163.367
R891 B.n245 B.n2 163.367
R892 B.n246 B.n245 163.367
R893 B.n246 B.n243 163.367
R894 B.n250 B.n243 163.367
R895 B.n251 B.n250 163.367
R896 B.n252 B.n251 163.367
R897 B.n252 B.n241 163.367
R898 B.n256 B.n241 163.367
R899 B.n257 B.n256 163.367
R900 B.n258 B.n257 163.367
R901 B.n258 B.n239 163.367
R902 B.n262 B.n239 163.367
R903 B.n263 B.n262 163.367
R904 B.n264 B.n263 163.367
R905 B.n264 B.n237 163.367
R906 B.n268 B.n237 163.367
R907 B.n269 B.n268 163.367
R908 B.n270 B.n269 163.367
R909 B.n270 B.n235 163.367
R910 B.n274 B.n235 163.367
R911 B.n275 B.n274 163.367
R912 B.n276 B.n275 163.367
R913 B.n276 B.n233 163.367
R914 B.n280 B.n233 163.367
R915 B.n281 B.n280 163.367
R916 B.n282 B.n281 163.367
R917 B.n282 B.n231 163.367
R918 B.n286 B.n231 163.367
R919 B.n287 B.n286 163.367
R920 B.n288 B.n287 163.367
R921 B.n288 B.n229 163.367
R922 B.n292 B.n229 163.367
R923 B.n293 B.n292 163.367
R924 B.n294 B.n293 163.367
R925 B.n294 B.n227 163.367
R926 B.n298 B.n227 163.367
R927 B.n299 B.n298 163.367
R928 B.n300 B.n299 163.367
R929 B.n300 B.n225 163.367
R930 B.n304 B.n225 163.367
R931 B.n305 B.n304 163.367
R932 B.n306 B.n305 163.367
R933 B.n306 B.n223 163.367
R934 B.n310 B.n223 163.367
R935 B.n311 B.n310 163.367
R936 B.n312 B.n311 163.367
R937 B.n312 B.n221 163.367
R938 B.n316 B.n221 163.367
R939 B.n317 B.n316 163.367
R940 B.n318 B.n317 163.367
R941 B.n318 B.n219 163.367
R942 B.n322 B.n219 163.367
R943 B.n323 B.n322 163.367
R944 B.n324 B.n323 163.367
R945 B.n324 B.n217 163.367
R946 B.n328 B.n217 163.367
R947 B.n329 B.n328 163.367
R948 B.n330 B.n329 163.367
R949 B.n330 B.n215 163.367
R950 B.n189 B.n188 69.0429
R951 B.n181 B.n180 69.0429
R952 B.n67 B.n66 69.0429
R953 B.n59 B.n58 69.0429
R954 B.n411 B.n189 59.5399
R955 B.n182 B.n181 59.5399
R956 B.n765 B.n67 59.5399
R957 B.n60 B.n59 59.5399
R958 B.n859 B.n32 34.4981
R959 B.n687 B.n686 34.4981
R960 B.n505 B.n154 34.4981
R961 B.n333 B.n332 34.4981
R962 B B.n949 18.0485
R963 B.n860 B.n859 10.6151
R964 B.n861 B.n860 10.6151
R965 B.n861 B.n30 10.6151
R966 B.n865 B.n30 10.6151
R967 B.n866 B.n865 10.6151
R968 B.n867 B.n866 10.6151
R969 B.n867 B.n28 10.6151
R970 B.n871 B.n28 10.6151
R971 B.n872 B.n871 10.6151
R972 B.n873 B.n872 10.6151
R973 B.n873 B.n26 10.6151
R974 B.n877 B.n26 10.6151
R975 B.n878 B.n877 10.6151
R976 B.n879 B.n878 10.6151
R977 B.n879 B.n24 10.6151
R978 B.n883 B.n24 10.6151
R979 B.n884 B.n883 10.6151
R980 B.n885 B.n884 10.6151
R981 B.n885 B.n22 10.6151
R982 B.n889 B.n22 10.6151
R983 B.n890 B.n889 10.6151
R984 B.n891 B.n890 10.6151
R985 B.n891 B.n20 10.6151
R986 B.n895 B.n20 10.6151
R987 B.n896 B.n895 10.6151
R988 B.n897 B.n896 10.6151
R989 B.n897 B.n18 10.6151
R990 B.n901 B.n18 10.6151
R991 B.n902 B.n901 10.6151
R992 B.n903 B.n902 10.6151
R993 B.n903 B.n16 10.6151
R994 B.n907 B.n16 10.6151
R995 B.n908 B.n907 10.6151
R996 B.n909 B.n908 10.6151
R997 B.n909 B.n14 10.6151
R998 B.n913 B.n14 10.6151
R999 B.n914 B.n913 10.6151
R1000 B.n915 B.n914 10.6151
R1001 B.n915 B.n12 10.6151
R1002 B.n919 B.n12 10.6151
R1003 B.n920 B.n919 10.6151
R1004 B.n921 B.n920 10.6151
R1005 B.n921 B.n10 10.6151
R1006 B.n925 B.n10 10.6151
R1007 B.n926 B.n925 10.6151
R1008 B.n927 B.n926 10.6151
R1009 B.n927 B.n8 10.6151
R1010 B.n931 B.n8 10.6151
R1011 B.n932 B.n931 10.6151
R1012 B.n933 B.n932 10.6151
R1013 B.n933 B.n6 10.6151
R1014 B.n937 B.n6 10.6151
R1015 B.n938 B.n937 10.6151
R1016 B.n939 B.n938 10.6151
R1017 B.n939 B.n4 10.6151
R1018 B.n943 B.n4 10.6151
R1019 B.n944 B.n943 10.6151
R1020 B.n945 B.n944 10.6151
R1021 B.n945 B.n0 10.6151
R1022 B.n855 B.n32 10.6151
R1023 B.n855 B.n854 10.6151
R1024 B.n854 B.n853 10.6151
R1025 B.n853 B.n34 10.6151
R1026 B.n849 B.n34 10.6151
R1027 B.n849 B.n848 10.6151
R1028 B.n848 B.n847 10.6151
R1029 B.n847 B.n36 10.6151
R1030 B.n843 B.n36 10.6151
R1031 B.n843 B.n842 10.6151
R1032 B.n842 B.n841 10.6151
R1033 B.n841 B.n38 10.6151
R1034 B.n837 B.n38 10.6151
R1035 B.n837 B.n836 10.6151
R1036 B.n836 B.n835 10.6151
R1037 B.n835 B.n40 10.6151
R1038 B.n831 B.n40 10.6151
R1039 B.n831 B.n830 10.6151
R1040 B.n830 B.n829 10.6151
R1041 B.n829 B.n42 10.6151
R1042 B.n825 B.n42 10.6151
R1043 B.n825 B.n824 10.6151
R1044 B.n824 B.n823 10.6151
R1045 B.n823 B.n44 10.6151
R1046 B.n819 B.n44 10.6151
R1047 B.n819 B.n818 10.6151
R1048 B.n818 B.n817 10.6151
R1049 B.n817 B.n46 10.6151
R1050 B.n813 B.n46 10.6151
R1051 B.n813 B.n812 10.6151
R1052 B.n812 B.n811 10.6151
R1053 B.n811 B.n48 10.6151
R1054 B.n807 B.n48 10.6151
R1055 B.n807 B.n806 10.6151
R1056 B.n806 B.n805 10.6151
R1057 B.n805 B.n50 10.6151
R1058 B.n801 B.n50 10.6151
R1059 B.n801 B.n800 10.6151
R1060 B.n800 B.n799 10.6151
R1061 B.n799 B.n52 10.6151
R1062 B.n795 B.n52 10.6151
R1063 B.n795 B.n794 10.6151
R1064 B.n794 B.n793 10.6151
R1065 B.n793 B.n54 10.6151
R1066 B.n789 B.n54 10.6151
R1067 B.n789 B.n788 10.6151
R1068 B.n788 B.n787 10.6151
R1069 B.n787 B.n56 10.6151
R1070 B.n783 B.n56 10.6151
R1071 B.n783 B.n782 10.6151
R1072 B.n782 B.n781 10.6151
R1073 B.n778 B.n777 10.6151
R1074 B.n777 B.n776 10.6151
R1075 B.n776 B.n62 10.6151
R1076 B.n772 B.n62 10.6151
R1077 B.n772 B.n771 10.6151
R1078 B.n771 B.n770 10.6151
R1079 B.n770 B.n64 10.6151
R1080 B.n766 B.n64 10.6151
R1081 B.n764 B.n763 10.6151
R1082 B.n763 B.n68 10.6151
R1083 B.n759 B.n68 10.6151
R1084 B.n759 B.n758 10.6151
R1085 B.n758 B.n757 10.6151
R1086 B.n757 B.n70 10.6151
R1087 B.n753 B.n70 10.6151
R1088 B.n753 B.n752 10.6151
R1089 B.n752 B.n751 10.6151
R1090 B.n751 B.n72 10.6151
R1091 B.n747 B.n72 10.6151
R1092 B.n747 B.n746 10.6151
R1093 B.n746 B.n745 10.6151
R1094 B.n745 B.n74 10.6151
R1095 B.n741 B.n74 10.6151
R1096 B.n741 B.n740 10.6151
R1097 B.n740 B.n739 10.6151
R1098 B.n739 B.n76 10.6151
R1099 B.n735 B.n76 10.6151
R1100 B.n735 B.n734 10.6151
R1101 B.n734 B.n733 10.6151
R1102 B.n733 B.n78 10.6151
R1103 B.n729 B.n78 10.6151
R1104 B.n729 B.n728 10.6151
R1105 B.n728 B.n727 10.6151
R1106 B.n727 B.n80 10.6151
R1107 B.n723 B.n80 10.6151
R1108 B.n723 B.n722 10.6151
R1109 B.n722 B.n721 10.6151
R1110 B.n721 B.n82 10.6151
R1111 B.n717 B.n82 10.6151
R1112 B.n717 B.n716 10.6151
R1113 B.n716 B.n715 10.6151
R1114 B.n715 B.n84 10.6151
R1115 B.n711 B.n84 10.6151
R1116 B.n711 B.n710 10.6151
R1117 B.n710 B.n709 10.6151
R1118 B.n709 B.n86 10.6151
R1119 B.n705 B.n86 10.6151
R1120 B.n705 B.n704 10.6151
R1121 B.n704 B.n703 10.6151
R1122 B.n703 B.n88 10.6151
R1123 B.n699 B.n88 10.6151
R1124 B.n699 B.n698 10.6151
R1125 B.n698 B.n697 10.6151
R1126 B.n697 B.n90 10.6151
R1127 B.n693 B.n90 10.6151
R1128 B.n693 B.n692 10.6151
R1129 B.n692 B.n691 10.6151
R1130 B.n691 B.n92 10.6151
R1131 B.n687 B.n92 10.6151
R1132 B.n686 B.n685 10.6151
R1133 B.n685 B.n94 10.6151
R1134 B.n681 B.n94 10.6151
R1135 B.n681 B.n680 10.6151
R1136 B.n680 B.n679 10.6151
R1137 B.n679 B.n96 10.6151
R1138 B.n675 B.n96 10.6151
R1139 B.n675 B.n674 10.6151
R1140 B.n674 B.n673 10.6151
R1141 B.n673 B.n98 10.6151
R1142 B.n669 B.n98 10.6151
R1143 B.n669 B.n668 10.6151
R1144 B.n668 B.n667 10.6151
R1145 B.n667 B.n100 10.6151
R1146 B.n663 B.n100 10.6151
R1147 B.n663 B.n662 10.6151
R1148 B.n662 B.n661 10.6151
R1149 B.n661 B.n102 10.6151
R1150 B.n657 B.n102 10.6151
R1151 B.n657 B.n656 10.6151
R1152 B.n656 B.n655 10.6151
R1153 B.n655 B.n104 10.6151
R1154 B.n651 B.n104 10.6151
R1155 B.n651 B.n650 10.6151
R1156 B.n650 B.n649 10.6151
R1157 B.n649 B.n106 10.6151
R1158 B.n645 B.n106 10.6151
R1159 B.n645 B.n644 10.6151
R1160 B.n644 B.n643 10.6151
R1161 B.n643 B.n108 10.6151
R1162 B.n639 B.n108 10.6151
R1163 B.n639 B.n638 10.6151
R1164 B.n638 B.n637 10.6151
R1165 B.n637 B.n110 10.6151
R1166 B.n633 B.n110 10.6151
R1167 B.n633 B.n632 10.6151
R1168 B.n632 B.n631 10.6151
R1169 B.n631 B.n112 10.6151
R1170 B.n627 B.n112 10.6151
R1171 B.n627 B.n626 10.6151
R1172 B.n626 B.n625 10.6151
R1173 B.n625 B.n114 10.6151
R1174 B.n621 B.n114 10.6151
R1175 B.n621 B.n620 10.6151
R1176 B.n620 B.n619 10.6151
R1177 B.n619 B.n116 10.6151
R1178 B.n615 B.n116 10.6151
R1179 B.n615 B.n614 10.6151
R1180 B.n614 B.n613 10.6151
R1181 B.n613 B.n118 10.6151
R1182 B.n609 B.n118 10.6151
R1183 B.n609 B.n608 10.6151
R1184 B.n608 B.n607 10.6151
R1185 B.n607 B.n120 10.6151
R1186 B.n603 B.n120 10.6151
R1187 B.n603 B.n602 10.6151
R1188 B.n602 B.n601 10.6151
R1189 B.n601 B.n122 10.6151
R1190 B.n597 B.n122 10.6151
R1191 B.n597 B.n596 10.6151
R1192 B.n596 B.n595 10.6151
R1193 B.n595 B.n124 10.6151
R1194 B.n591 B.n124 10.6151
R1195 B.n591 B.n590 10.6151
R1196 B.n590 B.n589 10.6151
R1197 B.n589 B.n126 10.6151
R1198 B.n585 B.n126 10.6151
R1199 B.n585 B.n584 10.6151
R1200 B.n584 B.n583 10.6151
R1201 B.n583 B.n128 10.6151
R1202 B.n579 B.n128 10.6151
R1203 B.n579 B.n578 10.6151
R1204 B.n578 B.n577 10.6151
R1205 B.n577 B.n130 10.6151
R1206 B.n573 B.n130 10.6151
R1207 B.n573 B.n572 10.6151
R1208 B.n572 B.n571 10.6151
R1209 B.n571 B.n132 10.6151
R1210 B.n567 B.n132 10.6151
R1211 B.n567 B.n566 10.6151
R1212 B.n566 B.n565 10.6151
R1213 B.n565 B.n134 10.6151
R1214 B.n561 B.n134 10.6151
R1215 B.n561 B.n560 10.6151
R1216 B.n560 B.n559 10.6151
R1217 B.n559 B.n136 10.6151
R1218 B.n555 B.n136 10.6151
R1219 B.n555 B.n554 10.6151
R1220 B.n554 B.n553 10.6151
R1221 B.n553 B.n138 10.6151
R1222 B.n549 B.n138 10.6151
R1223 B.n549 B.n548 10.6151
R1224 B.n548 B.n547 10.6151
R1225 B.n547 B.n140 10.6151
R1226 B.n543 B.n140 10.6151
R1227 B.n543 B.n542 10.6151
R1228 B.n542 B.n541 10.6151
R1229 B.n541 B.n142 10.6151
R1230 B.n537 B.n142 10.6151
R1231 B.n537 B.n536 10.6151
R1232 B.n536 B.n535 10.6151
R1233 B.n535 B.n144 10.6151
R1234 B.n531 B.n144 10.6151
R1235 B.n531 B.n530 10.6151
R1236 B.n530 B.n529 10.6151
R1237 B.n529 B.n146 10.6151
R1238 B.n525 B.n146 10.6151
R1239 B.n525 B.n524 10.6151
R1240 B.n524 B.n523 10.6151
R1241 B.n523 B.n148 10.6151
R1242 B.n519 B.n148 10.6151
R1243 B.n519 B.n518 10.6151
R1244 B.n518 B.n517 10.6151
R1245 B.n517 B.n150 10.6151
R1246 B.n513 B.n150 10.6151
R1247 B.n513 B.n512 10.6151
R1248 B.n512 B.n511 10.6151
R1249 B.n511 B.n152 10.6151
R1250 B.n507 B.n152 10.6151
R1251 B.n507 B.n506 10.6151
R1252 B.n506 B.n505 10.6151
R1253 B.n244 B.n1 10.6151
R1254 B.n247 B.n244 10.6151
R1255 B.n248 B.n247 10.6151
R1256 B.n249 B.n248 10.6151
R1257 B.n249 B.n242 10.6151
R1258 B.n253 B.n242 10.6151
R1259 B.n254 B.n253 10.6151
R1260 B.n255 B.n254 10.6151
R1261 B.n255 B.n240 10.6151
R1262 B.n259 B.n240 10.6151
R1263 B.n260 B.n259 10.6151
R1264 B.n261 B.n260 10.6151
R1265 B.n261 B.n238 10.6151
R1266 B.n265 B.n238 10.6151
R1267 B.n266 B.n265 10.6151
R1268 B.n267 B.n266 10.6151
R1269 B.n267 B.n236 10.6151
R1270 B.n271 B.n236 10.6151
R1271 B.n272 B.n271 10.6151
R1272 B.n273 B.n272 10.6151
R1273 B.n273 B.n234 10.6151
R1274 B.n277 B.n234 10.6151
R1275 B.n278 B.n277 10.6151
R1276 B.n279 B.n278 10.6151
R1277 B.n279 B.n232 10.6151
R1278 B.n283 B.n232 10.6151
R1279 B.n284 B.n283 10.6151
R1280 B.n285 B.n284 10.6151
R1281 B.n285 B.n230 10.6151
R1282 B.n289 B.n230 10.6151
R1283 B.n290 B.n289 10.6151
R1284 B.n291 B.n290 10.6151
R1285 B.n291 B.n228 10.6151
R1286 B.n295 B.n228 10.6151
R1287 B.n296 B.n295 10.6151
R1288 B.n297 B.n296 10.6151
R1289 B.n297 B.n226 10.6151
R1290 B.n301 B.n226 10.6151
R1291 B.n302 B.n301 10.6151
R1292 B.n303 B.n302 10.6151
R1293 B.n303 B.n224 10.6151
R1294 B.n307 B.n224 10.6151
R1295 B.n308 B.n307 10.6151
R1296 B.n309 B.n308 10.6151
R1297 B.n309 B.n222 10.6151
R1298 B.n313 B.n222 10.6151
R1299 B.n314 B.n313 10.6151
R1300 B.n315 B.n314 10.6151
R1301 B.n315 B.n220 10.6151
R1302 B.n319 B.n220 10.6151
R1303 B.n320 B.n319 10.6151
R1304 B.n321 B.n320 10.6151
R1305 B.n321 B.n218 10.6151
R1306 B.n325 B.n218 10.6151
R1307 B.n326 B.n325 10.6151
R1308 B.n327 B.n326 10.6151
R1309 B.n327 B.n216 10.6151
R1310 B.n331 B.n216 10.6151
R1311 B.n332 B.n331 10.6151
R1312 B.n333 B.n214 10.6151
R1313 B.n337 B.n214 10.6151
R1314 B.n338 B.n337 10.6151
R1315 B.n339 B.n338 10.6151
R1316 B.n339 B.n212 10.6151
R1317 B.n343 B.n212 10.6151
R1318 B.n344 B.n343 10.6151
R1319 B.n345 B.n344 10.6151
R1320 B.n345 B.n210 10.6151
R1321 B.n349 B.n210 10.6151
R1322 B.n350 B.n349 10.6151
R1323 B.n351 B.n350 10.6151
R1324 B.n351 B.n208 10.6151
R1325 B.n355 B.n208 10.6151
R1326 B.n356 B.n355 10.6151
R1327 B.n357 B.n356 10.6151
R1328 B.n357 B.n206 10.6151
R1329 B.n361 B.n206 10.6151
R1330 B.n362 B.n361 10.6151
R1331 B.n363 B.n362 10.6151
R1332 B.n363 B.n204 10.6151
R1333 B.n367 B.n204 10.6151
R1334 B.n368 B.n367 10.6151
R1335 B.n369 B.n368 10.6151
R1336 B.n369 B.n202 10.6151
R1337 B.n373 B.n202 10.6151
R1338 B.n374 B.n373 10.6151
R1339 B.n375 B.n374 10.6151
R1340 B.n375 B.n200 10.6151
R1341 B.n379 B.n200 10.6151
R1342 B.n380 B.n379 10.6151
R1343 B.n381 B.n380 10.6151
R1344 B.n381 B.n198 10.6151
R1345 B.n385 B.n198 10.6151
R1346 B.n386 B.n385 10.6151
R1347 B.n387 B.n386 10.6151
R1348 B.n387 B.n196 10.6151
R1349 B.n391 B.n196 10.6151
R1350 B.n392 B.n391 10.6151
R1351 B.n393 B.n392 10.6151
R1352 B.n393 B.n194 10.6151
R1353 B.n397 B.n194 10.6151
R1354 B.n398 B.n397 10.6151
R1355 B.n399 B.n398 10.6151
R1356 B.n399 B.n192 10.6151
R1357 B.n403 B.n192 10.6151
R1358 B.n404 B.n403 10.6151
R1359 B.n405 B.n404 10.6151
R1360 B.n405 B.n190 10.6151
R1361 B.n409 B.n190 10.6151
R1362 B.n410 B.n409 10.6151
R1363 B.n412 B.n186 10.6151
R1364 B.n416 B.n186 10.6151
R1365 B.n417 B.n416 10.6151
R1366 B.n418 B.n417 10.6151
R1367 B.n418 B.n184 10.6151
R1368 B.n422 B.n184 10.6151
R1369 B.n423 B.n422 10.6151
R1370 B.n424 B.n423 10.6151
R1371 B.n428 B.n427 10.6151
R1372 B.n429 B.n428 10.6151
R1373 B.n429 B.n178 10.6151
R1374 B.n433 B.n178 10.6151
R1375 B.n434 B.n433 10.6151
R1376 B.n435 B.n434 10.6151
R1377 B.n435 B.n176 10.6151
R1378 B.n439 B.n176 10.6151
R1379 B.n440 B.n439 10.6151
R1380 B.n441 B.n440 10.6151
R1381 B.n441 B.n174 10.6151
R1382 B.n445 B.n174 10.6151
R1383 B.n446 B.n445 10.6151
R1384 B.n447 B.n446 10.6151
R1385 B.n447 B.n172 10.6151
R1386 B.n451 B.n172 10.6151
R1387 B.n452 B.n451 10.6151
R1388 B.n453 B.n452 10.6151
R1389 B.n453 B.n170 10.6151
R1390 B.n457 B.n170 10.6151
R1391 B.n458 B.n457 10.6151
R1392 B.n459 B.n458 10.6151
R1393 B.n459 B.n168 10.6151
R1394 B.n463 B.n168 10.6151
R1395 B.n464 B.n463 10.6151
R1396 B.n465 B.n464 10.6151
R1397 B.n465 B.n166 10.6151
R1398 B.n469 B.n166 10.6151
R1399 B.n470 B.n469 10.6151
R1400 B.n471 B.n470 10.6151
R1401 B.n471 B.n164 10.6151
R1402 B.n475 B.n164 10.6151
R1403 B.n476 B.n475 10.6151
R1404 B.n477 B.n476 10.6151
R1405 B.n477 B.n162 10.6151
R1406 B.n481 B.n162 10.6151
R1407 B.n482 B.n481 10.6151
R1408 B.n483 B.n482 10.6151
R1409 B.n483 B.n160 10.6151
R1410 B.n487 B.n160 10.6151
R1411 B.n488 B.n487 10.6151
R1412 B.n489 B.n488 10.6151
R1413 B.n489 B.n158 10.6151
R1414 B.n493 B.n158 10.6151
R1415 B.n494 B.n493 10.6151
R1416 B.n495 B.n494 10.6151
R1417 B.n495 B.n156 10.6151
R1418 B.n499 B.n156 10.6151
R1419 B.n500 B.n499 10.6151
R1420 B.n501 B.n500 10.6151
R1421 B.n501 B.n154 10.6151
R1422 B.n949 B.n0 8.11757
R1423 B.n949 B.n1 8.11757
R1424 B.n778 B.n60 6.5566
R1425 B.n766 B.n765 6.5566
R1426 B.n412 B.n411 6.5566
R1427 B.n424 B.n182 6.5566
R1428 B.n781 B.n60 4.05904
R1429 B.n765 B.n764 4.05904
R1430 B.n411 B.n410 4.05904
R1431 B.n427 B.n182 4.05904
R1432 VP.n24 VP.n23 161.3
R1433 VP.n25 VP.n20 161.3
R1434 VP.n27 VP.n26 161.3
R1435 VP.n28 VP.n19 161.3
R1436 VP.n30 VP.n29 161.3
R1437 VP.n31 VP.n18 161.3
R1438 VP.n33 VP.n32 161.3
R1439 VP.n35 VP.n34 161.3
R1440 VP.n36 VP.n16 161.3
R1441 VP.n38 VP.n37 161.3
R1442 VP.n39 VP.n15 161.3
R1443 VP.n41 VP.n40 161.3
R1444 VP.n42 VP.n14 161.3
R1445 VP.n44 VP.n43 161.3
R1446 VP.n79 VP.n78 161.3
R1447 VP.n77 VP.n1 161.3
R1448 VP.n76 VP.n75 161.3
R1449 VP.n74 VP.n2 161.3
R1450 VP.n73 VP.n72 161.3
R1451 VP.n71 VP.n3 161.3
R1452 VP.n70 VP.n69 161.3
R1453 VP.n68 VP.n67 161.3
R1454 VP.n66 VP.n5 161.3
R1455 VP.n65 VP.n64 161.3
R1456 VP.n63 VP.n6 161.3
R1457 VP.n62 VP.n61 161.3
R1458 VP.n60 VP.n7 161.3
R1459 VP.n59 VP.n58 161.3
R1460 VP.n57 VP.n56 161.3
R1461 VP.n55 VP.n9 161.3
R1462 VP.n54 VP.n53 161.3
R1463 VP.n52 VP.n10 161.3
R1464 VP.n51 VP.n50 161.3
R1465 VP.n49 VP.n11 161.3
R1466 VP.n48 VP.n47 161.3
R1467 VP.n22 VP.t6 148.882
R1468 VP.n12 VP.t5 115.725
R1469 VP.n8 VP.t0 115.725
R1470 VP.n4 VP.t7 115.725
R1471 VP.n0 VP.t1 115.725
R1472 VP.n13 VP.t2 115.725
R1473 VP.n17 VP.t3 115.725
R1474 VP.n21 VP.t4 115.725
R1475 VP.n46 VP.n12 73.4298
R1476 VP.n80 VP.n0 73.4298
R1477 VP.n45 VP.n13 73.4298
R1478 VP.n22 VP.n21 60.5173
R1479 VP.n46 VP.n45 56.6281
R1480 VP.n50 VP.n10 46.321
R1481 VP.n76 VP.n2 46.321
R1482 VP.n41 VP.n15 46.321
R1483 VP.n61 VP.n6 40.4934
R1484 VP.n65 VP.n6 40.4934
R1485 VP.n30 VP.n19 40.4934
R1486 VP.n26 VP.n19 40.4934
R1487 VP.n54 VP.n10 34.6658
R1488 VP.n72 VP.n2 34.6658
R1489 VP.n37 VP.n15 34.6658
R1490 VP.n49 VP.n48 24.4675
R1491 VP.n50 VP.n49 24.4675
R1492 VP.n55 VP.n54 24.4675
R1493 VP.n56 VP.n55 24.4675
R1494 VP.n60 VP.n59 24.4675
R1495 VP.n61 VP.n60 24.4675
R1496 VP.n66 VP.n65 24.4675
R1497 VP.n67 VP.n66 24.4675
R1498 VP.n71 VP.n70 24.4675
R1499 VP.n72 VP.n71 24.4675
R1500 VP.n77 VP.n76 24.4675
R1501 VP.n78 VP.n77 24.4675
R1502 VP.n42 VP.n41 24.4675
R1503 VP.n43 VP.n42 24.4675
R1504 VP.n31 VP.n30 24.4675
R1505 VP.n32 VP.n31 24.4675
R1506 VP.n36 VP.n35 24.4675
R1507 VP.n37 VP.n36 24.4675
R1508 VP.n25 VP.n24 24.4675
R1509 VP.n26 VP.n25 24.4675
R1510 VP.n48 VP.n12 16.6381
R1511 VP.n78 VP.n0 16.6381
R1512 VP.n43 VP.n13 16.6381
R1513 VP.n59 VP.n8 13.702
R1514 VP.n67 VP.n4 13.702
R1515 VP.n32 VP.n17 13.702
R1516 VP.n24 VP.n21 13.702
R1517 VP.n56 VP.n8 10.766
R1518 VP.n70 VP.n4 10.766
R1519 VP.n35 VP.n17 10.766
R1520 VP.n23 VP.n22 4.06449
R1521 VP.n45 VP.n44 0.354971
R1522 VP.n47 VP.n46 0.354971
R1523 VP.n80 VP.n79 0.354971
R1524 VP VP.n80 0.26696
R1525 VP.n23 VP.n20 0.189894
R1526 VP.n27 VP.n20 0.189894
R1527 VP.n28 VP.n27 0.189894
R1528 VP.n29 VP.n28 0.189894
R1529 VP.n29 VP.n18 0.189894
R1530 VP.n33 VP.n18 0.189894
R1531 VP.n34 VP.n33 0.189894
R1532 VP.n34 VP.n16 0.189894
R1533 VP.n38 VP.n16 0.189894
R1534 VP.n39 VP.n38 0.189894
R1535 VP.n40 VP.n39 0.189894
R1536 VP.n40 VP.n14 0.189894
R1537 VP.n44 VP.n14 0.189894
R1538 VP.n47 VP.n11 0.189894
R1539 VP.n51 VP.n11 0.189894
R1540 VP.n52 VP.n51 0.189894
R1541 VP.n53 VP.n52 0.189894
R1542 VP.n53 VP.n9 0.189894
R1543 VP.n57 VP.n9 0.189894
R1544 VP.n58 VP.n57 0.189894
R1545 VP.n58 VP.n7 0.189894
R1546 VP.n62 VP.n7 0.189894
R1547 VP.n63 VP.n62 0.189894
R1548 VP.n64 VP.n63 0.189894
R1549 VP.n64 VP.n5 0.189894
R1550 VP.n68 VP.n5 0.189894
R1551 VP.n69 VP.n68 0.189894
R1552 VP.n69 VP.n3 0.189894
R1553 VP.n73 VP.n3 0.189894
R1554 VP.n74 VP.n73 0.189894
R1555 VP.n75 VP.n74 0.189894
R1556 VP.n75 VP.n1 0.189894
R1557 VP.n79 VP.n1 0.189894
R1558 VTAIL.n690 VTAIL.n610 756.745
R1559 VTAIL.n82 VTAIL.n2 756.745
R1560 VTAIL.n168 VTAIL.n88 756.745
R1561 VTAIL.n256 VTAIL.n176 756.745
R1562 VTAIL.n604 VTAIL.n524 756.745
R1563 VTAIL.n516 VTAIL.n436 756.745
R1564 VTAIL.n430 VTAIL.n350 756.745
R1565 VTAIL.n342 VTAIL.n262 756.745
R1566 VTAIL.n639 VTAIL.n638 585
R1567 VTAIL.n641 VTAIL.n640 585
R1568 VTAIL.n634 VTAIL.n633 585
R1569 VTAIL.n647 VTAIL.n646 585
R1570 VTAIL.n649 VTAIL.n648 585
R1571 VTAIL.n630 VTAIL.n629 585
R1572 VTAIL.n655 VTAIL.n654 585
R1573 VTAIL.n657 VTAIL.n656 585
R1574 VTAIL.n626 VTAIL.n625 585
R1575 VTAIL.n663 VTAIL.n662 585
R1576 VTAIL.n665 VTAIL.n664 585
R1577 VTAIL.n622 VTAIL.n621 585
R1578 VTAIL.n671 VTAIL.n670 585
R1579 VTAIL.n673 VTAIL.n672 585
R1580 VTAIL.n618 VTAIL.n617 585
R1581 VTAIL.n680 VTAIL.n679 585
R1582 VTAIL.n681 VTAIL.n616 585
R1583 VTAIL.n683 VTAIL.n682 585
R1584 VTAIL.n614 VTAIL.n613 585
R1585 VTAIL.n689 VTAIL.n688 585
R1586 VTAIL.n691 VTAIL.n690 585
R1587 VTAIL.n31 VTAIL.n30 585
R1588 VTAIL.n33 VTAIL.n32 585
R1589 VTAIL.n26 VTAIL.n25 585
R1590 VTAIL.n39 VTAIL.n38 585
R1591 VTAIL.n41 VTAIL.n40 585
R1592 VTAIL.n22 VTAIL.n21 585
R1593 VTAIL.n47 VTAIL.n46 585
R1594 VTAIL.n49 VTAIL.n48 585
R1595 VTAIL.n18 VTAIL.n17 585
R1596 VTAIL.n55 VTAIL.n54 585
R1597 VTAIL.n57 VTAIL.n56 585
R1598 VTAIL.n14 VTAIL.n13 585
R1599 VTAIL.n63 VTAIL.n62 585
R1600 VTAIL.n65 VTAIL.n64 585
R1601 VTAIL.n10 VTAIL.n9 585
R1602 VTAIL.n72 VTAIL.n71 585
R1603 VTAIL.n73 VTAIL.n8 585
R1604 VTAIL.n75 VTAIL.n74 585
R1605 VTAIL.n6 VTAIL.n5 585
R1606 VTAIL.n81 VTAIL.n80 585
R1607 VTAIL.n83 VTAIL.n82 585
R1608 VTAIL.n117 VTAIL.n116 585
R1609 VTAIL.n119 VTAIL.n118 585
R1610 VTAIL.n112 VTAIL.n111 585
R1611 VTAIL.n125 VTAIL.n124 585
R1612 VTAIL.n127 VTAIL.n126 585
R1613 VTAIL.n108 VTAIL.n107 585
R1614 VTAIL.n133 VTAIL.n132 585
R1615 VTAIL.n135 VTAIL.n134 585
R1616 VTAIL.n104 VTAIL.n103 585
R1617 VTAIL.n141 VTAIL.n140 585
R1618 VTAIL.n143 VTAIL.n142 585
R1619 VTAIL.n100 VTAIL.n99 585
R1620 VTAIL.n149 VTAIL.n148 585
R1621 VTAIL.n151 VTAIL.n150 585
R1622 VTAIL.n96 VTAIL.n95 585
R1623 VTAIL.n158 VTAIL.n157 585
R1624 VTAIL.n159 VTAIL.n94 585
R1625 VTAIL.n161 VTAIL.n160 585
R1626 VTAIL.n92 VTAIL.n91 585
R1627 VTAIL.n167 VTAIL.n166 585
R1628 VTAIL.n169 VTAIL.n168 585
R1629 VTAIL.n205 VTAIL.n204 585
R1630 VTAIL.n207 VTAIL.n206 585
R1631 VTAIL.n200 VTAIL.n199 585
R1632 VTAIL.n213 VTAIL.n212 585
R1633 VTAIL.n215 VTAIL.n214 585
R1634 VTAIL.n196 VTAIL.n195 585
R1635 VTAIL.n221 VTAIL.n220 585
R1636 VTAIL.n223 VTAIL.n222 585
R1637 VTAIL.n192 VTAIL.n191 585
R1638 VTAIL.n229 VTAIL.n228 585
R1639 VTAIL.n231 VTAIL.n230 585
R1640 VTAIL.n188 VTAIL.n187 585
R1641 VTAIL.n237 VTAIL.n236 585
R1642 VTAIL.n239 VTAIL.n238 585
R1643 VTAIL.n184 VTAIL.n183 585
R1644 VTAIL.n246 VTAIL.n245 585
R1645 VTAIL.n247 VTAIL.n182 585
R1646 VTAIL.n249 VTAIL.n248 585
R1647 VTAIL.n180 VTAIL.n179 585
R1648 VTAIL.n255 VTAIL.n254 585
R1649 VTAIL.n257 VTAIL.n256 585
R1650 VTAIL.n605 VTAIL.n604 585
R1651 VTAIL.n603 VTAIL.n602 585
R1652 VTAIL.n528 VTAIL.n527 585
R1653 VTAIL.n532 VTAIL.n530 585
R1654 VTAIL.n597 VTAIL.n596 585
R1655 VTAIL.n595 VTAIL.n594 585
R1656 VTAIL.n534 VTAIL.n533 585
R1657 VTAIL.n589 VTAIL.n588 585
R1658 VTAIL.n587 VTAIL.n586 585
R1659 VTAIL.n538 VTAIL.n537 585
R1660 VTAIL.n581 VTAIL.n580 585
R1661 VTAIL.n579 VTAIL.n578 585
R1662 VTAIL.n542 VTAIL.n541 585
R1663 VTAIL.n573 VTAIL.n572 585
R1664 VTAIL.n571 VTAIL.n570 585
R1665 VTAIL.n546 VTAIL.n545 585
R1666 VTAIL.n565 VTAIL.n564 585
R1667 VTAIL.n563 VTAIL.n562 585
R1668 VTAIL.n550 VTAIL.n549 585
R1669 VTAIL.n557 VTAIL.n556 585
R1670 VTAIL.n555 VTAIL.n554 585
R1671 VTAIL.n517 VTAIL.n516 585
R1672 VTAIL.n515 VTAIL.n514 585
R1673 VTAIL.n440 VTAIL.n439 585
R1674 VTAIL.n444 VTAIL.n442 585
R1675 VTAIL.n509 VTAIL.n508 585
R1676 VTAIL.n507 VTAIL.n506 585
R1677 VTAIL.n446 VTAIL.n445 585
R1678 VTAIL.n501 VTAIL.n500 585
R1679 VTAIL.n499 VTAIL.n498 585
R1680 VTAIL.n450 VTAIL.n449 585
R1681 VTAIL.n493 VTAIL.n492 585
R1682 VTAIL.n491 VTAIL.n490 585
R1683 VTAIL.n454 VTAIL.n453 585
R1684 VTAIL.n485 VTAIL.n484 585
R1685 VTAIL.n483 VTAIL.n482 585
R1686 VTAIL.n458 VTAIL.n457 585
R1687 VTAIL.n477 VTAIL.n476 585
R1688 VTAIL.n475 VTAIL.n474 585
R1689 VTAIL.n462 VTAIL.n461 585
R1690 VTAIL.n469 VTAIL.n468 585
R1691 VTAIL.n467 VTAIL.n466 585
R1692 VTAIL.n431 VTAIL.n430 585
R1693 VTAIL.n429 VTAIL.n428 585
R1694 VTAIL.n354 VTAIL.n353 585
R1695 VTAIL.n358 VTAIL.n356 585
R1696 VTAIL.n423 VTAIL.n422 585
R1697 VTAIL.n421 VTAIL.n420 585
R1698 VTAIL.n360 VTAIL.n359 585
R1699 VTAIL.n415 VTAIL.n414 585
R1700 VTAIL.n413 VTAIL.n412 585
R1701 VTAIL.n364 VTAIL.n363 585
R1702 VTAIL.n407 VTAIL.n406 585
R1703 VTAIL.n405 VTAIL.n404 585
R1704 VTAIL.n368 VTAIL.n367 585
R1705 VTAIL.n399 VTAIL.n398 585
R1706 VTAIL.n397 VTAIL.n396 585
R1707 VTAIL.n372 VTAIL.n371 585
R1708 VTAIL.n391 VTAIL.n390 585
R1709 VTAIL.n389 VTAIL.n388 585
R1710 VTAIL.n376 VTAIL.n375 585
R1711 VTAIL.n383 VTAIL.n382 585
R1712 VTAIL.n381 VTAIL.n380 585
R1713 VTAIL.n343 VTAIL.n342 585
R1714 VTAIL.n341 VTAIL.n340 585
R1715 VTAIL.n266 VTAIL.n265 585
R1716 VTAIL.n270 VTAIL.n268 585
R1717 VTAIL.n335 VTAIL.n334 585
R1718 VTAIL.n333 VTAIL.n332 585
R1719 VTAIL.n272 VTAIL.n271 585
R1720 VTAIL.n327 VTAIL.n326 585
R1721 VTAIL.n325 VTAIL.n324 585
R1722 VTAIL.n276 VTAIL.n275 585
R1723 VTAIL.n319 VTAIL.n318 585
R1724 VTAIL.n317 VTAIL.n316 585
R1725 VTAIL.n280 VTAIL.n279 585
R1726 VTAIL.n311 VTAIL.n310 585
R1727 VTAIL.n309 VTAIL.n308 585
R1728 VTAIL.n284 VTAIL.n283 585
R1729 VTAIL.n303 VTAIL.n302 585
R1730 VTAIL.n301 VTAIL.n300 585
R1731 VTAIL.n288 VTAIL.n287 585
R1732 VTAIL.n295 VTAIL.n294 585
R1733 VTAIL.n293 VTAIL.n292 585
R1734 VTAIL.n637 VTAIL.t4 327.466
R1735 VTAIL.n29 VTAIL.t2 327.466
R1736 VTAIL.n115 VTAIL.t9 327.466
R1737 VTAIL.n203 VTAIL.t13 327.466
R1738 VTAIL.n553 VTAIL.t10 327.466
R1739 VTAIL.n465 VTAIL.t14 327.466
R1740 VTAIL.n379 VTAIL.t1 327.466
R1741 VTAIL.n291 VTAIL.t6 327.466
R1742 VTAIL.n640 VTAIL.n639 171.744
R1743 VTAIL.n640 VTAIL.n633 171.744
R1744 VTAIL.n647 VTAIL.n633 171.744
R1745 VTAIL.n648 VTAIL.n647 171.744
R1746 VTAIL.n648 VTAIL.n629 171.744
R1747 VTAIL.n655 VTAIL.n629 171.744
R1748 VTAIL.n656 VTAIL.n655 171.744
R1749 VTAIL.n656 VTAIL.n625 171.744
R1750 VTAIL.n663 VTAIL.n625 171.744
R1751 VTAIL.n664 VTAIL.n663 171.744
R1752 VTAIL.n664 VTAIL.n621 171.744
R1753 VTAIL.n671 VTAIL.n621 171.744
R1754 VTAIL.n672 VTAIL.n671 171.744
R1755 VTAIL.n672 VTAIL.n617 171.744
R1756 VTAIL.n680 VTAIL.n617 171.744
R1757 VTAIL.n681 VTAIL.n680 171.744
R1758 VTAIL.n682 VTAIL.n681 171.744
R1759 VTAIL.n682 VTAIL.n613 171.744
R1760 VTAIL.n689 VTAIL.n613 171.744
R1761 VTAIL.n690 VTAIL.n689 171.744
R1762 VTAIL.n32 VTAIL.n31 171.744
R1763 VTAIL.n32 VTAIL.n25 171.744
R1764 VTAIL.n39 VTAIL.n25 171.744
R1765 VTAIL.n40 VTAIL.n39 171.744
R1766 VTAIL.n40 VTAIL.n21 171.744
R1767 VTAIL.n47 VTAIL.n21 171.744
R1768 VTAIL.n48 VTAIL.n47 171.744
R1769 VTAIL.n48 VTAIL.n17 171.744
R1770 VTAIL.n55 VTAIL.n17 171.744
R1771 VTAIL.n56 VTAIL.n55 171.744
R1772 VTAIL.n56 VTAIL.n13 171.744
R1773 VTAIL.n63 VTAIL.n13 171.744
R1774 VTAIL.n64 VTAIL.n63 171.744
R1775 VTAIL.n64 VTAIL.n9 171.744
R1776 VTAIL.n72 VTAIL.n9 171.744
R1777 VTAIL.n73 VTAIL.n72 171.744
R1778 VTAIL.n74 VTAIL.n73 171.744
R1779 VTAIL.n74 VTAIL.n5 171.744
R1780 VTAIL.n81 VTAIL.n5 171.744
R1781 VTAIL.n82 VTAIL.n81 171.744
R1782 VTAIL.n118 VTAIL.n117 171.744
R1783 VTAIL.n118 VTAIL.n111 171.744
R1784 VTAIL.n125 VTAIL.n111 171.744
R1785 VTAIL.n126 VTAIL.n125 171.744
R1786 VTAIL.n126 VTAIL.n107 171.744
R1787 VTAIL.n133 VTAIL.n107 171.744
R1788 VTAIL.n134 VTAIL.n133 171.744
R1789 VTAIL.n134 VTAIL.n103 171.744
R1790 VTAIL.n141 VTAIL.n103 171.744
R1791 VTAIL.n142 VTAIL.n141 171.744
R1792 VTAIL.n142 VTAIL.n99 171.744
R1793 VTAIL.n149 VTAIL.n99 171.744
R1794 VTAIL.n150 VTAIL.n149 171.744
R1795 VTAIL.n150 VTAIL.n95 171.744
R1796 VTAIL.n158 VTAIL.n95 171.744
R1797 VTAIL.n159 VTAIL.n158 171.744
R1798 VTAIL.n160 VTAIL.n159 171.744
R1799 VTAIL.n160 VTAIL.n91 171.744
R1800 VTAIL.n167 VTAIL.n91 171.744
R1801 VTAIL.n168 VTAIL.n167 171.744
R1802 VTAIL.n206 VTAIL.n205 171.744
R1803 VTAIL.n206 VTAIL.n199 171.744
R1804 VTAIL.n213 VTAIL.n199 171.744
R1805 VTAIL.n214 VTAIL.n213 171.744
R1806 VTAIL.n214 VTAIL.n195 171.744
R1807 VTAIL.n221 VTAIL.n195 171.744
R1808 VTAIL.n222 VTAIL.n221 171.744
R1809 VTAIL.n222 VTAIL.n191 171.744
R1810 VTAIL.n229 VTAIL.n191 171.744
R1811 VTAIL.n230 VTAIL.n229 171.744
R1812 VTAIL.n230 VTAIL.n187 171.744
R1813 VTAIL.n237 VTAIL.n187 171.744
R1814 VTAIL.n238 VTAIL.n237 171.744
R1815 VTAIL.n238 VTAIL.n183 171.744
R1816 VTAIL.n246 VTAIL.n183 171.744
R1817 VTAIL.n247 VTAIL.n246 171.744
R1818 VTAIL.n248 VTAIL.n247 171.744
R1819 VTAIL.n248 VTAIL.n179 171.744
R1820 VTAIL.n255 VTAIL.n179 171.744
R1821 VTAIL.n256 VTAIL.n255 171.744
R1822 VTAIL.n604 VTAIL.n603 171.744
R1823 VTAIL.n603 VTAIL.n527 171.744
R1824 VTAIL.n532 VTAIL.n527 171.744
R1825 VTAIL.n596 VTAIL.n532 171.744
R1826 VTAIL.n596 VTAIL.n595 171.744
R1827 VTAIL.n595 VTAIL.n533 171.744
R1828 VTAIL.n588 VTAIL.n533 171.744
R1829 VTAIL.n588 VTAIL.n587 171.744
R1830 VTAIL.n587 VTAIL.n537 171.744
R1831 VTAIL.n580 VTAIL.n537 171.744
R1832 VTAIL.n580 VTAIL.n579 171.744
R1833 VTAIL.n579 VTAIL.n541 171.744
R1834 VTAIL.n572 VTAIL.n541 171.744
R1835 VTAIL.n572 VTAIL.n571 171.744
R1836 VTAIL.n571 VTAIL.n545 171.744
R1837 VTAIL.n564 VTAIL.n545 171.744
R1838 VTAIL.n564 VTAIL.n563 171.744
R1839 VTAIL.n563 VTAIL.n549 171.744
R1840 VTAIL.n556 VTAIL.n549 171.744
R1841 VTAIL.n556 VTAIL.n555 171.744
R1842 VTAIL.n516 VTAIL.n515 171.744
R1843 VTAIL.n515 VTAIL.n439 171.744
R1844 VTAIL.n444 VTAIL.n439 171.744
R1845 VTAIL.n508 VTAIL.n444 171.744
R1846 VTAIL.n508 VTAIL.n507 171.744
R1847 VTAIL.n507 VTAIL.n445 171.744
R1848 VTAIL.n500 VTAIL.n445 171.744
R1849 VTAIL.n500 VTAIL.n499 171.744
R1850 VTAIL.n499 VTAIL.n449 171.744
R1851 VTAIL.n492 VTAIL.n449 171.744
R1852 VTAIL.n492 VTAIL.n491 171.744
R1853 VTAIL.n491 VTAIL.n453 171.744
R1854 VTAIL.n484 VTAIL.n453 171.744
R1855 VTAIL.n484 VTAIL.n483 171.744
R1856 VTAIL.n483 VTAIL.n457 171.744
R1857 VTAIL.n476 VTAIL.n457 171.744
R1858 VTAIL.n476 VTAIL.n475 171.744
R1859 VTAIL.n475 VTAIL.n461 171.744
R1860 VTAIL.n468 VTAIL.n461 171.744
R1861 VTAIL.n468 VTAIL.n467 171.744
R1862 VTAIL.n430 VTAIL.n429 171.744
R1863 VTAIL.n429 VTAIL.n353 171.744
R1864 VTAIL.n358 VTAIL.n353 171.744
R1865 VTAIL.n422 VTAIL.n358 171.744
R1866 VTAIL.n422 VTAIL.n421 171.744
R1867 VTAIL.n421 VTAIL.n359 171.744
R1868 VTAIL.n414 VTAIL.n359 171.744
R1869 VTAIL.n414 VTAIL.n413 171.744
R1870 VTAIL.n413 VTAIL.n363 171.744
R1871 VTAIL.n406 VTAIL.n363 171.744
R1872 VTAIL.n406 VTAIL.n405 171.744
R1873 VTAIL.n405 VTAIL.n367 171.744
R1874 VTAIL.n398 VTAIL.n367 171.744
R1875 VTAIL.n398 VTAIL.n397 171.744
R1876 VTAIL.n397 VTAIL.n371 171.744
R1877 VTAIL.n390 VTAIL.n371 171.744
R1878 VTAIL.n390 VTAIL.n389 171.744
R1879 VTAIL.n389 VTAIL.n375 171.744
R1880 VTAIL.n382 VTAIL.n375 171.744
R1881 VTAIL.n382 VTAIL.n381 171.744
R1882 VTAIL.n342 VTAIL.n341 171.744
R1883 VTAIL.n341 VTAIL.n265 171.744
R1884 VTAIL.n270 VTAIL.n265 171.744
R1885 VTAIL.n334 VTAIL.n270 171.744
R1886 VTAIL.n334 VTAIL.n333 171.744
R1887 VTAIL.n333 VTAIL.n271 171.744
R1888 VTAIL.n326 VTAIL.n271 171.744
R1889 VTAIL.n326 VTAIL.n325 171.744
R1890 VTAIL.n325 VTAIL.n275 171.744
R1891 VTAIL.n318 VTAIL.n275 171.744
R1892 VTAIL.n318 VTAIL.n317 171.744
R1893 VTAIL.n317 VTAIL.n279 171.744
R1894 VTAIL.n310 VTAIL.n279 171.744
R1895 VTAIL.n310 VTAIL.n309 171.744
R1896 VTAIL.n309 VTAIL.n283 171.744
R1897 VTAIL.n302 VTAIL.n283 171.744
R1898 VTAIL.n302 VTAIL.n301 171.744
R1899 VTAIL.n301 VTAIL.n287 171.744
R1900 VTAIL.n294 VTAIL.n287 171.744
R1901 VTAIL.n294 VTAIL.n293 171.744
R1902 VTAIL.n639 VTAIL.t4 85.8723
R1903 VTAIL.n31 VTAIL.t2 85.8723
R1904 VTAIL.n117 VTAIL.t9 85.8723
R1905 VTAIL.n205 VTAIL.t13 85.8723
R1906 VTAIL.n555 VTAIL.t10 85.8723
R1907 VTAIL.n467 VTAIL.t14 85.8723
R1908 VTAIL.n381 VTAIL.t1 85.8723
R1909 VTAIL.n293 VTAIL.t6 85.8723
R1910 VTAIL.n523 VTAIL.n522 56.4885
R1911 VTAIL.n349 VTAIL.n348 56.4885
R1912 VTAIL.n1 VTAIL.n0 56.4883
R1913 VTAIL.n175 VTAIL.n174 56.4883
R1914 VTAIL.n695 VTAIL.n694 35.0944
R1915 VTAIL.n87 VTAIL.n86 35.0944
R1916 VTAIL.n173 VTAIL.n172 35.0944
R1917 VTAIL.n261 VTAIL.n260 35.0944
R1918 VTAIL.n609 VTAIL.n608 35.0944
R1919 VTAIL.n521 VTAIL.n520 35.0944
R1920 VTAIL.n435 VTAIL.n434 35.0944
R1921 VTAIL.n347 VTAIL.n346 35.0944
R1922 VTAIL.n695 VTAIL.n609 28.8065
R1923 VTAIL.n347 VTAIL.n261 28.8065
R1924 VTAIL.n638 VTAIL.n637 16.3895
R1925 VTAIL.n30 VTAIL.n29 16.3895
R1926 VTAIL.n116 VTAIL.n115 16.3895
R1927 VTAIL.n204 VTAIL.n203 16.3895
R1928 VTAIL.n554 VTAIL.n553 16.3895
R1929 VTAIL.n466 VTAIL.n465 16.3895
R1930 VTAIL.n380 VTAIL.n379 16.3895
R1931 VTAIL.n292 VTAIL.n291 16.3895
R1932 VTAIL.n683 VTAIL.n614 13.1884
R1933 VTAIL.n75 VTAIL.n6 13.1884
R1934 VTAIL.n161 VTAIL.n92 13.1884
R1935 VTAIL.n249 VTAIL.n180 13.1884
R1936 VTAIL.n530 VTAIL.n528 13.1884
R1937 VTAIL.n442 VTAIL.n440 13.1884
R1938 VTAIL.n356 VTAIL.n354 13.1884
R1939 VTAIL.n268 VTAIL.n266 13.1884
R1940 VTAIL.n641 VTAIL.n636 12.8005
R1941 VTAIL.n684 VTAIL.n616 12.8005
R1942 VTAIL.n688 VTAIL.n687 12.8005
R1943 VTAIL.n33 VTAIL.n28 12.8005
R1944 VTAIL.n76 VTAIL.n8 12.8005
R1945 VTAIL.n80 VTAIL.n79 12.8005
R1946 VTAIL.n119 VTAIL.n114 12.8005
R1947 VTAIL.n162 VTAIL.n94 12.8005
R1948 VTAIL.n166 VTAIL.n165 12.8005
R1949 VTAIL.n207 VTAIL.n202 12.8005
R1950 VTAIL.n250 VTAIL.n182 12.8005
R1951 VTAIL.n254 VTAIL.n253 12.8005
R1952 VTAIL.n602 VTAIL.n601 12.8005
R1953 VTAIL.n598 VTAIL.n597 12.8005
R1954 VTAIL.n557 VTAIL.n552 12.8005
R1955 VTAIL.n514 VTAIL.n513 12.8005
R1956 VTAIL.n510 VTAIL.n509 12.8005
R1957 VTAIL.n469 VTAIL.n464 12.8005
R1958 VTAIL.n428 VTAIL.n427 12.8005
R1959 VTAIL.n424 VTAIL.n423 12.8005
R1960 VTAIL.n383 VTAIL.n378 12.8005
R1961 VTAIL.n340 VTAIL.n339 12.8005
R1962 VTAIL.n336 VTAIL.n335 12.8005
R1963 VTAIL.n295 VTAIL.n290 12.8005
R1964 VTAIL.n642 VTAIL.n634 12.0247
R1965 VTAIL.n679 VTAIL.n678 12.0247
R1966 VTAIL.n691 VTAIL.n612 12.0247
R1967 VTAIL.n34 VTAIL.n26 12.0247
R1968 VTAIL.n71 VTAIL.n70 12.0247
R1969 VTAIL.n83 VTAIL.n4 12.0247
R1970 VTAIL.n120 VTAIL.n112 12.0247
R1971 VTAIL.n157 VTAIL.n156 12.0247
R1972 VTAIL.n169 VTAIL.n90 12.0247
R1973 VTAIL.n208 VTAIL.n200 12.0247
R1974 VTAIL.n245 VTAIL.n244 12.0247
R1975 VTAIL.n257 VTAIL.n178 12.0247
R1976 VTAIL.n605 VTAIL.n526 12.0247
R1977 VTAIL.n594 VTAIL.n531 12.0247
R1978 VTAIL.n558 VTAIL.n550 12.0247
R1979 VTAIL.n517 VTAIL.n438 12.0247
R1980 VTAIL.n506 VTAIL.n443 12.0247
R1981 VTAIL.n470 VTAIL.n462 12.0247
R1982 VTAIL.n431 VTAIL.n352 12.0247
R1983 VTAIL.n420 VTAIL.n357 12.0247
R1984 VTAIL.n384 VTAIL.n376 12.0247
R1985 VTAIL.n343 VTAIL.n264 12.0247
R1986 VTAIL.n332 VTAIL.n269 12.0247
R1987 VTAIL.n296 VTAIL.n288 12.0247
R1988 VTAIL.n646 VTAIL.n645 11.249
R1989 VTAIL.n677 VTAIL.n618 11.249
R1990 VTAIL.n692 VTAIL.n610 11.249
R1991 VTAIL.n38 VTAIL.n37 11.249
R1992 VTAIL.n69 VTAIL.n10 11.249
R1993 VTAIL.n84 VTAIL.n2 11.249
R1994 VTAIL.n124 VTAIL.n123 11.249
R1995 VTAIL.n155 VTAIL.n96 11.249
R1996 VTAIL.n170 VTAIL.n88 11.249
R1997 VTAIL.n212 VTAIL.n211 11.249
R1998 VTAIL.n243 VTAIL.n184 11.249
R1999 VTAIL.n258 VTAIL.n176 11.249
R2000 VTAIL.n606 VTAIL.n524 11.249
R2001 VTAIL.n593 VTAIL.n534 11.249
R2002 VTAIL.n562 VTAIL.n561 11.249
R2003 VTAIL.n518 VTAIL.n436 11.249
R2004 VTAIL.n505 VTAIL.n446 11.249
R2005 VTAIL.n474 VTAIL.n473 11.249
R2006 VTAIL.n432 VTAIL.n350 11.249
R2007 VTAIL.n419 VTAIL.n360 11.249
R2008 VTAIL.n388 VTAIL.n387 11.249
R2009 VTAIL.n344 VTAIL.n262 11.249
R2010 VTAIL.n331 VTAIL.n272 11.249
R2011 VTAIL.n300 VTAIL.n299 11.249
R2012 VTAIL.n649 VTAIL.n632 10.4732
R2013 VTAIL.n674 VTAIL.n673 10.4732
R2014 VTAIL.n41 VTAIL.n24 10.4732
R2015 VTAIL.n66 VTAIL.n65 10.4732
R2016 VTAIL.n127 VTAIL.n110 10.4732
R2017 VTAIL.n152 VTAIL.n151 10.4732
R2018 VTAIL.n215 VTAIL.n198 10.4732
R2019 VTAIL.n240 VTAIL.n239 10.4732
R2020 VTAIL.n590 VTAIL.n589 10.4732
R2021 VTAIL.n565 VTAIL.n548 10.4732
R2022 VTAIL.n502 VTAIL.n501 10.4732
R2023 VTAIL.n477 VTAIL.n460 10.4732
R2024 VTAIL.n416 VTAIL.n415 10.4732
R2025 VTAIL.n391 VTAIL.n374 10.4732
R2026 VTAIL.n328 VTAIL.n327 10.4732
R2027 VTAIL.n303 VTAIL.n286 10.4732
R2028 VTAIL.n650 VTAIL.n630 9.69747
R2029 VTAIL.n670 VTAIL.n620 9.69747
R2030 VTAIL.n42 VTAIL.n22 9.69747
R2031 VTAIL.n62 VTAIL.n12 9.69747
R2032 VTAIL.n128 VTAIL.n108 9.69747
R2033 VTAIL.n148 VTAIL.n98 9.69747
R2034 VTAIL.n216 VTAIL.n196 9.69747
R2035 VTAIL.n236 VTAIL.n186 9.69747
R2036 VTAIL.n586 VTAIL.n536 9.69747
R2037 VTAIL.n566 VTAIL.n546 9.69747
R2038 VTAIL.n498 VTAIL.n448 9.69747
R2039 VTAIL.n478 VTAIL.n458 9.69747
R2040 VTAIL.n412 VTAIL.n362 9.69747
R2041 VTAIL.n392 VTAIL.n372 9.69747
R2042 VTAIL.n324 VTAIL.n274 9.69747
R2043 VTAIL.n304 VTAIL.n284 9.69747
R2044 VTAIL.n694 VTAIL.n693 9.45567
R2045 VTAIL.n86 VTAIL.n85 9.45567
R2046 VTAIL.n172 VTAIL.n171 9.45567
R2047 VTAIL.n260 VTAIL.n259 9.45567
R2048 VTAIL.n608 VTAIL.n607 9.45567
R2049 VTAIL.n520 VTAIL.n519 9.45567
R2050 VTAIL.n434 VTAIL.n433 9.45567
R2051 VTAIL.n346 VTAIL.n345 9.45567
R2052 VTAIL.n693 VTAIL.n692 9.3005
R2053 VTAIL.n612 VTAIL.n611 9.3005
R2054 VTAIL.n687 VTAIL.n686 9.3005
R2055 VTAIL.n659 VTAIL.n658 9.3005
R2056 VTAIL.n628 VTAIL.n627 9.3005
R2057 VTAIL.n653 VTAIL.n652 9.3005
R2058 VTAIL.n651 VTAIL.n650 9.3005
R2059 VTAIL.n632 VTAIL.n631 9.3005
R2060 VTAIL.n645 VTAIL.n644 9.3005
R2061 VTAIL.n643 VTAIL.n642 9.3005
R2062 VTAIL.n636 VTAIL.n635 9.3005
R2063 VTAIL.n661 VTAIL.n660 9.3005
R2064 VTAIL.n624 VTAIL.n623 9.3005
R2065 VTAIL.n667 VTAIL.n666 9.3005
R2066 VTAIL.n669 VTAIL.n668 9.3005
R2067 VTAIL.n620 VTAIL.n619 9.3005
R2068 VTAIL.n675 VTAIL.n674 9.3005
R2069 VTAIL.n677 VTAIL.n676 9.3005
R2070 VTAIL.n678 VTAIL.n615 9.3005
R2071 VTAIL.n685 VTAIL.n684 9.3005
R2072 VTAIL.n85 VTAIL.n84 9.3005
R2073 VTAIL.n4 VTAIL.n3 9.3005
R2074 VTAIL.n79 VTAIL.n78 9.3005
R2075 VTAIL.n51 VTAIL.n50 9.3005
R2076 VTAIL.n20 VTAIL.n19 9.3005
R2077 VTAIL.n45 VTAIL.n44 9.3005
R2078 VTAIL.n43 VTAIL.n42 9.3005
R2079 VTAIL.n24 VTAIL.n23 9.3005
R2080 VTAIL.n37 VTAIL.n36 9.3005
R2081 VTAIL.n35 VTAIL.n34 9.3005
R2082 VTAIL.n28 VTAIL.n27 9.3005
R2083 VTAIL.n53 VTAIL.n52 9.3005
R2084 VTAIL.n16 VTAIL.n15 9.3005
R2085 VTAIL.n59 VTAIL.n58 9.3005
R2086 VTAIL.n61 VTAIL.n60 9.3005
R2087 VTAIL.n12 VTAIL.n11 9.3005
R2088 VTAIL.n67 VTAIL.n66 9.3005
R2089 VTAIL.n69 VTAIL.n68 9.3005
R2090 VTAIL.n70 VTAIL.n7 9.3005
R2091 VTAIL.n77 VTAIL.n76 9.3005
R2092 VTAIL.n171 VTAIL.n170 9.3005
R2093 VTAIL.n90 VTAIL.n89 9.3005
R2094 VTAIL.n165 VTAIL.n164 9.3005
R2095 VTAIL.n137 VTAIL.n136 9.3005
R2096 VTAIL.n106 VTAIL.n105 9.3005
R2097 VTAIL.n131 VTAIL.n130 9.3005
R2098 VTAIL.n129 VTAIL.n128 9.3005
R2099 VTAIL.n110 VTAIL.n109 9.3005
R2100 VTAIL.n123 VTAIL.n122 9.3005
R2101 VTAIL.n121 VTAIL.n120 9.3005
R2102 VTAIL.n114 VTAIL.n113 9.3005
R2103 VTAIL.n139 VTAIL.n138 9.3005
R2104 VTAIL.n102 VTAIL.n101 9.3005
R2105 VTAIL.n145 VTAIL.n144 9.3005
R2106 VTAIL.n147 VTAIL.n146 9.3005
R2107 VTAIL.n98 VTAIL.n97 9.3005
R2108 VTAIL.n153 VTAIL.n152 9.3005
R2109 VTAIL.n155 VTAIL.n154 9.3005
R2110 VTAIL.n156 VTAIL.n93 9.3005
R2111 VTAIL.n163 VTAIL.n162 9.3005
R2112 VTAIL.n259 VTAIL.n258 9.3005
R2113 VTAIL.n178 VTAIL.n177 9.3005
R2114 VTAIL.n253 VTAIL.n252 9.3005
R2115 VTAIL.n225 VTAIL.n224 9.3005
R2116 VTAIL.n194 VTAIL.n193 9.3005
R2117 VTAIL.n219 VTAIL.n218 9.3005
R2118 VTAIL.n217 VTAIL.n216 9.3005
R2119 VTAIL.n198 VTAIL.n197 9.3005
R2120 VTAIL.n211 VTAIL.n210 9.3005
R2121 VTAIL.n209 VTAIL.n208 9.3005
R2122 VTAIL.n202 VTAIL.n201 9.3005
R2123 VTAIL.n227 VTAIL.n226 9.3005
R2124 VTAIL.n190 VTAIL.n189 9.3005
R2125 VTAIL.n233 VTAIL.n232 9.3005
R2126 VTAIL.n235 VTAIL.n234 9.3005
R2127 VTAIL.n186 VTAIL.n185 9.3005
R2128 VTAIL.n241 VTAIL.n240 9.3005
R2129 VTAIL.n243 VTAIL.n242 9.3005
R2130 VTAIL.n244 VTAIL.n181 9.3005
R2131 VTAIL.n251 VTAIL.n250 9.3005
R2132 VTAIL.n540 VTAIL.n539 9.3005
R2133 VTAIL.n583 VTAIL.n582 9.3005
R2134 VTAIL.n585 VTAIL.n584 9.3005
R2135 VTAIL.n536 VTAIL.n535 9.3005
R2136 VTAIL.n591 VTAIL.n590 9.3005
R2137 VTAIL.n593 VTAIL.n592 9.3005
R2138 VTAIL.n531 VTAIL.n529 9.3005
R2139 VTAIL.n599 VTAIL.n598 9.3005
R2140 VTAIL.n607 VTAIL.n606 9.3005
R2141 VTAIL.n526 VTAIL.n525 9.3005
R2142 VTAIL.n601 VTAIL.n600 9.3005
R2143 VTAIL.n577 VTAIL.n576 9.3005
R2144 VTAIL.n575 VTAIL.n574 9.3005
R2145 VTAIL.n544 VTAIL.n543 9.3005
R2146 VTAIL.n569 VTAIL.n568 9.3005
R2147 VTAIL.n567 VTAIL.n566 9.3005
R2148 VTAIL.n548 VTAIL.n547 9.3005
R2149 VTAIL.n561 VTAIL.n560 9.3005
R2150 VTAIL.n559 VTAIL.n558 9.3005
R2151 VTAIL.n552 VTAIL.n551 9.3005
R2152 VTAIL.n452 VTAIL.n451 9.3005
R2153 VTAIL.n495 VTAIL.n494 9.3005
R2154 VTAIL.n497 VTAIL.n496 9.3005
R2155 VTAIL.n448 VTAIL.n447 9.3005
R2156 VTAIL.n503 VTAIL.n502 9.3005
R2157 VTAIL.n505 VTAIL.n504 9.3005
R2158 VTAIL.n443 VTAIL.n441 9.3005
R2159 VTAIL.n511 VTAIL.n510 9.3005
R2160 VTAIL.n519 VTAIL.n518 9.3005
R2161 VTAIL.n438 VTAIL.n437 9.3005
R2162 VTAIL.n513 VTAIL.n512 9.3005
R2163 VTAIL.n489 VTAIL.n488 9.3005
R2164 VTAIL.n487 VTAIL.n486 9.3005
R2165 VTAIL.n456 VTAIL.n455 9.3005
R2166 VTAIL.n481 VTAIL.n480 9.3005
R2167 VTAIL.n479 VTAIL.n478 9.3005
R2168 VTAIL.n460 VTAIL.n459 9.3005
R2169 VTAIL.n473 VTAIL.n472 9.3005
R2170 VTAIL.n471 VTAIL.n470 9.3005
R2171 VTAIL.n464 VTAIL.n463 9.3005
R2172 VTAIL.n366 VTAIL.n365 9.3005
R2173 VTAIL.n409 VTAIL.n408 9.3005
R2174 VTAIL.n411 VTAIL.n410 9.3005
R2175 VTAIL.n362 VTAIL.n361 9.3005
R2176 VTAIL.n417 VTAIL.n416 9.3005
R2177 VTAIL.n419 VTAIL.n418 9.3005
R2178 VTAIL.n357 VTAIL.n355 9.3005
R2179 VTAIL.n425 VTAIL.n424 9.3005
R2180 VTAIL.n433 VTAIL.n432 9.3005
R2181 VTAIL.n352 VTAIL.n351 9.3005
R2182 VTAIL.n427 VTAIL.n426 9.3005
R2183 VTAIL.n403 VTAIL.n402 9.3005
R2184 VTAIL.n401 VTAIL.n400 9.3005
R2185 VTAIL.n370 VTAIL.n369 9.3005
R2186 VTAIL.n395 VTAIL.n394 9.3005
R2187 VTAIL.n393 VTAIL.n392 9.3005
R2188 VTAIL.n374 VTAIL.n373 9.3005
R2189 VTAIL.n387 VTAIL.n386 9.3005
R2190 VTAIL.n385 VTAIL.n384 9.3005
R2191 VTAIL.n378 VTAIL.n377 9.3005
R2192 VTAIL.n278 VTAIL.n277 9.3005
R2193 VTAIL.n321 VTAIL.n320 9.3005
R2194 VTAIL.n323 VTAIL.n322 9.3005
R2195 VTAIL.n274 VTAIL.n273 9.3005
R2196 VTAIL.n329 VTAIL.n328 9.3005
R2197 VTAIL.n331 VTAIL.n330 9.3005
R2198 VTAIL.n269 VTAIL.n267 9.3005
R2199 VTAIL.n337 VTAIL.n336 9.3005
R2200 VTAIL.n345 VTAIL.n344 9.3005
R2201 VTAIL.n264 VTAIL.n263 9.3005
R2202 VTAIL.n339 VTAIL.n338 9.3005
R2203 VTAIL.n315 VTAIL.n314 9.3005
R2204 VTAIL.n313 VTAIL.n312 9.3005
R2205 VTAIL.n282 VTAIL.n281 9.3005
R2206 VTAIL.n307 VTAIL.n306 9.3005
R2207 VTAIL.n305 VTAIL.n304 9.3005
R2208 VTAIL.n286 VTAIL.n285 9.3005
R2209 VTAIL.n299 VTAIL.n298 9.3005
R2210 VTAIL.n297 VTAIL.n296 9.3005
R2211 VTAIL.n290 VTAIL.n289 9.3005
R2212 VTAIL.n654 VTAIL.n653 8.92171
R2213 VTAIL.n669 VTAIL.n622 8.92171
R2214 VTAIL.n46 VTAIL.n45 8.92171
R2215 VTAIL.n61 VTAIL.n14 8.92171
R2216 VTAIL.n132 VTAIL.n131 8.92171
R2217 VTAIL.n147 VTAIL.n100 8.92171
R2218 VTAIL.n220 VTAIL.n219 8.92171
R2219 VTAIL.n235 VTAIL.n188 8.92171
R2220 VTAIL.n585 VTAIL.n538 8.92171
R2221 VTAIL.n570 VTAIL.n569 8.92171
R2222 VTAIL.n497 VTAIL.n450 8.92171
R2223 VTAIL.n482 VTAIL.n481 8.92171
R2224 VTAIL.n411 VTAIL.n364 8.92171
R2225 VTAIL.n396 VTAIL.n395 8.92171
R2226 VTAIL.n323 VTAIL.n276 8.92171
R2227 VTAIL.n308 VTAIL.n307 8.92171
R2228 VTAIL.n657 VTAIL.n628 8.14595
R2229 VTAIL.n666 VTAIL.n665 8.14595
R2230 VTAIL.n49 VTAIL.n20 8.14595
R2231 VTAIL.n58 VTAIL.n57 8.14595
R2232 VTAIL.n135 VTAIL.n106 8.14595
R2233 VTAIL.n144 VTAIL.n143 8.14595
R2234 VTAIL.n223 VTAIL.n194 8.14595
R2235 VTAIL.n232 VTAIL.n231 8.14595
R2236 VTAIL.n582 VTAIL.n581 8.14595
R2237 VTAIL.n573 VTAIL.n544 8.14595
R2238 VTAIL.n494 VTAIL.n493 8.14595
R2239 VTAIL.n485 VTAIL.n456 8.14595
R2240 VTAIL.n408 VTAIL.n407 8.14595
R2241 VTAIL.n399 VTAIL.n370 8.14595
R2242 VTAIL.n320 VTAIL.n319 8.14595
R2243 VTAIL.n311 VTAIL.n282 8.14595
R2244 VTAIL.n658 VTAIL.n626 7.3702
R2245 VTAIL.n662 VTAIL.n624 7.3702
R2246 VTAIL.n50 VTAIL.n18 7.3702
R2247 VTAIL.n54 VTAIL.n16 7.3702
R2248 VTAIL.n136 VTAIL.n104 7.3702
R2249 VTAIL.n140 VTAIL.n102 7.3702
R2250 VTAIL.n224 VTAIL.n192 7.3702
R2251 VTAIL.n228 VTAIL.n190 7.3702
R2252 VTAIL.n578 VTAIL.n540 7.3702
R2253 VTAIL.n574 VTAIL.n542 7.3702
R2254 VTAIL.n490 VTAIL.n452 7.3702
R2255 VTAIL.n486 VTAIL.n454 7.3702
R2256 VTAIL.n404 VTAIL.n366 7.3702
R2257 VTAIL.n400 VTAIL.n368 7.3702
R2258 VTAIL.n316 VTAIL.n278 7.3702
R2259 VTAIL.n312 VTAIL.n280 7.3702
R2260 VTAIL.n661 VTAIL.n626 6.59444
R2261 VTAIL.n662 VTAIL.n661 6.59444
R2262 VTAIL.n53 VTAIL.n18 6.59444
R2263 VTAIL.n54 VTAIL.n53 6.59444
R2264 VTAIL.n139 VTAIL.n104 6.59444
R2265 VTAIL.n140 VTAIL.n139 6.59444
R2266 VTAIL.n227 VTAIL.n192 6.59444
R2267 VTAIL.n228 VTAIL.n227 6.59444
R2268 VTAIL.n578 VTAIL.n577 6.59444
R2269 VTAIL.n577 VTAIL.n542 6.59444
R2270 VTAIL.n490 VTAIL.n489 6.59444
R2271 VTAIL.n489 VTAIL.n454 6.59444
R2272 VTAIL.n404 VTAIL.n403 6.59444
R2273 VTAIL.n403 VTAIL.n368 6.59444
R2274 VTAIL.n316 VTAIL.n315 6.59444
R2275 VTAIL.n315 VTAIL.n280 6.59444
R2276 VTAIL.n658 VTAIL.n657 5.81868
R2277 VTAIL.n665 VTAIL.n624 5.81868
R2278 VTAIL.n50 VTAIL.n49 5.81868
R2279 VTAIL.n57 VTAIL.n16 5.81868
R2280 VTAIL.n136 VTAIL.n135 5.81868
R2281 VTAIL.n143 VTAIL.n102 5.81868
R2282 VTAIL.n224 VTAIL.n223 5.81868
R2283 VTAIL.n231 VTAIL.n190 5.81868
R2284 VTAIL.n581 VTAIL.n540 5.81868
R2285 VTAIL.n574 VTAIL.n573 5.81868
R2286 VTAIL.n493 VTAIL.n452 5.81868
R2287 VTAIL.n486 VTAIL.n485 5.81868
R2288 VTAIL.n407 VTAIL.n366 5.81868
R2289 VTAIL.n400 VTAIL.n399 5.81868
R2290 VTAIL.n319 VTAIL.n278 5.81868
R2291 VTAIL.n312 VTAIL.n311 5.81868
R2292 VTAIL.n654 VTAIL.n628 5.04292
R2293 VTAIL.n666 VTAIL.n622 5.04292
R2294 VTAIL.n46 VTAIL.n20 5.04292
R2295 VTAIL.n58 VTAIL.n14 5.04292
R2296 VTAIL.n132 VTAIL.n106 5.04292
R2297 VTAIL.n144 VTAIL.n100 5.04292
R2298 VTAIL.n220 VTAIL.n194 5.04292
R2299 VTAIL.n232 VTAIL.n188 5.04292
R2300 VTAIL.n582 VTAIL.n538 5.04292
R2301 VTAIL.n570 VTAIL.n544 5.04292
R2302 VTAIL.n494 VTAIL.n450 5.04292
R2303 VTAIL.n482 VTAIL.n456 5.04292
R2304 VTAIL.n408 VTAIL.n364 5.04292
R2305 VTAIL.n396 VTAIL.n370 5.04292
R2306 VTAIL.n320 VTAIL.n276 5.04292
R2307 VTAIL.n308 VTAIL.n282 5.04292
R2308 VTAIL.n653 VTAIL.n630 4.26717
R2309 VTAIL.n670 VTAIL.n669 4.26717
R2310 VTAIL.n45 VTAIL.n22 4.26717
R2311 VTAIL.n62 VTAIL.n61 4.26717
R2312 VTAIL.n131 VTAIL.n108 4.26717
R2313 VTAIL.n148 VTAIL.n147 4.26717
R2314 VTAIL.n219 VTAIL.n196 4.26717
R2315 VTAIL.n236 VTAIL.n235 4.26717
R2316 VTAIL.n586 VTAIL.n585 4.26717
R2317 VTAIL.n569 VTAIL.n546 4.26717
R2318 VTAIL.n498 VTAIL.n497 4.26717
R2319 VTAIL.n481 VTAIL.n458 4.26717
R2320 VTAIL.n412 VTAIL.n411 4.26717
R2321 VTAIL.n395 VTAIL.n372 4.26717
R2322 VTAIL.n324 VTAIL.n323 4.26717
R2323 VTAIL.n307 VTAIL.n284 4.26717
R2324 VTAIL.n637 VTAIL.n635 3.70982
R2325 VTAIL.n29 VTAIL.n27 3.70982
R2326 VTAIL.n115 VTAIL.n113 3.70982
R2327 VTAIL.n203 VTAIL.n201 3.70982
R2328 VTAIL.n553 VTAIL.n551 3.70982
R2329 VTAIL.n465 VTAIL.n463 3.70982
R2330 VTAIL.n379 VTAIL.n377 3.70982
R2331 VTAIL.n291 VTAIL.n289 3.70982
R2332 VTAIL.n650 VTAIL.n649 3.49141
R2333 VTAIL.n673 VTAIL.n620 3.49141
R2334 VTAIL.n42 VTAIL.n41 3.49141
R2335 VTAIL.n65 VTAIL.n12 3.49141
R2336 VTAIL.n128 VTAIL.n127 3.49141
R2337 VTAIL.n151 VTAIL.n98 3.49141
R2338 VTAIL.n216 VTAIL.n215 3.49141
R2339 VTAIL.n239 VTAIL.n186 3.49141
R2340 VTAIL.n589 VTAIL.n536 3.49141
R2341 VTAIL.n566 VTAIL.n565 3.49141
R2342 VTAIL.n501 VTAIL.n448 3.49141
R2343 VTAIL.n478 VTAIL.n477 3.49141
R2344 VTAIL.n415 VTAIL.n362 3.49141
R2345 VTAIL.n392 VTAIL.n391 3.49141
R2346 VTAIL.n327 VTAIL.n274 3.49141
R2347 VTAIL.n304 VTAIL.n303 3.49141
R2348 VTAIL.n349 VTAIL.n347 3.06947
R2349 VTAIL.n435 VTAIL.n349 3.06947
R2350 VTAIL.n523 VTAIL.n521 3.06947
R2351 VTAIL.n609 VTAIL.n523 3.06947
R2352 VTAIL.n261 VTAIL.n175 3.06947
R2353 VTAIL.n175 VTAIL.n173 3.06947
R2354 VTAIL.n87 VTAIL.n1 3.06947
R2355 VTAIL VTAIL.n695 3.01128
R2356 VTAIL.n646 VTAIL.n632 2.71565
R2357 VTAIL.n674 VTAIL.n618 2.71565
R2358 VTAIL.n694 VTAIL.n610 2.71565
R2359 VTAIL.n38 VTAIL.n24 2.71565
R2360 VTAIL.n66 VTAIL.n10 2.71565
R2361 VTAIL.n86 VTAIL.n2 2.71565
R2362 VTAIL.n124 VTAIL.n110 2.71565
R2363 VTAIL.n152 VTAIL.n96 2.71565
R2364 VTAIL.n172 VTAIL.n88 2.71565
R2365 VTAIL.n212 VTAIL.n198 2.71565
R2366 VTAIL.n240 VTAIL.n184 2.71565
R2367 VTAIL.n260 VTAIL.n176 2.71565
R2368 VTAIL.n608 VTAIL.n524 2.71565
R2369 VTAIL.n590 VTAIL.n534 2.71565
R2370 VTAIL.n562 VTAIL.n548 2.71565
R2371 VTAIL.n520 VTAIL.n436 2.71565
R2372 VTAIL.n502 VTAIL.n446 2.71565
R2373 VTAIL.n474 VTAIL.n460 2.71565
R2374 VTAIL.n434 VTAIL.n350 2.71565
R2375 VTAIL.n416 VTAIL.n360 2.71565
R2376 VTAIL.n388 VTAIL.n374 2.71565
R2377 VTAIL.n346 VTAIL.n262 2.71565
R2378 VTAIL.n328 VTAIL.n272 2.71565
R2379 VTAIL.n300 VTAIL.n286 2.71565
R2380 VTAIL.n0 VTAIL.t5 2.09624
R2381 VTAIL.n0 VTAIL.t3 2.09624
R2382 VTAIL.n174 VTAIL.t8 2.09624
R2383 VTAIL.n174 VTAIL.t15 2.09624
R2384 VTAIL.n522 VTAIL.t12 2.09624
R2385 VTAIL.n522 VTAIL.t11 2.09624
R2386 VTAIL.n348 VTAIL.t0 2.09624
R2387 VTAIL.n348 VTAIL.t7 2.09624
R2388 VTAIL.n645 VTAIL.n634 1.93989
R2389 VTAIL.n679 VTAIL.n677 1.93989
R2390 VTAIL.n692 VTAIL.n691 1.93989
R2391 VTAIL.n37 VTAIL.n26 1.93989
R2392 VTAIL.n71 VTAIL.n69 1.93989
R2393 VTAIL.n84 VTAIL.n83 1.93989
R2394 VTAIL.n123 VTAIL.n112 1.93989
R2395 VTAIL.n157 VTAIL.n155 1.93989
R2396 VTAIL.n170 VTAIL.n169 1.93989
R2397 VTAIL.n211 VTAIL.n200 1.93989
R2398 VTAIL.n245 VTAIL.n243 1.93989
R2399 VTAIL.n258 VTAIL.n257 1.93989
R2400 VTAIL.n606 VTAIL.n605 1.93989
R2401 VTAIL.n594 VTAIL.n593 1.93989
R2402 VTAIL.n561 VTAIL.n550 1.93989
R2403 VTAIL.n518 VTAIL.n517 1.93989
R2404 VTAIL.n506 VTAIL.n505 1.93989
R2405 VTAIL.n473 VTAIL.n462 1.93989
R2406 VTAIL.n432 VTAIL.n431 1.93989
R2407 VTAIL.n420 VTAIL.n419 1.93989
R2408 VTAIL.n387 VTAIL.n376 1.93989
R2409 VTAIL.n344 VTAIL.n343 1.93989
R2410 VTAIL.n332 VTAIL.n331 1.93989
R2411 VTAIL.n299 VTAIL.n288 1.93989
R2412 VTAIL.n642 VTAIL.n641 1.16414
R2413 VTAIL.n678 VTAIL.n616 1.16414
R2414 VTAIL.n688 VTAIL.n612 1.16414
R2415 VTAIL.n34 VTAIL.n33 1.16414
R2416 VTAIL.n70 VTAIL.n8 1.16414
R2417 VTAIL.n80 VTAIL.n4 1.16414
R2418 VTAIL.n120 VTAIL.n119 1.16414
R2419 VTAIL.n156 VTAIL.n94 1.16414
R2420 VTAIL.n166 VTAIL.n90 1.16414
R2421 VTAIL.n208 VTAIL.n207 1.16414
R2422 VTAIL.n244 VTAIL.n182 1.16414
R2423 VTAIL.n254 VTAIL.n178 1.16414
R2424 VTAIL.n602 VTAIL.n526 1.16414
R2425 VTAIL.n597 VTAIL.n531 1.16414
R2426 VTAIL.n558 VTAIL.n557 1.16414
R2427 VTAIL.n514 VTAIL.n438 1.16414
R2428 VTAIL.n509 VTAIL.n443 1.16414
R2429 VTAIL.n470 VTAIL.n469 1.16414
R2430 VTAIL.n428 VTAIL.n352 1.16414
R2431 VTAIL.n423 VTAIL.n357 1.16414
R2432 VTAIL.n384 VTAIL.n383 1.16414
R2433 VTAIL.n340 VTAIL.n264 1.16414
R2434 VTAIL.n335 VTAIL.n269 1.16414
R2435 VTAIL.n296 VTAIL.n295 1.16414
R2436 VTAIL.n521 VTAIL.n435 0.470328
R2437 VTAIL.n173 VTAIL.n87 0.470328
R2438 VTAIL.n638 VTAIL.n636 0.388379
R2439 VTAIL.n684 VTAIL.n683 0.388379
R2440 VTAIL.n687 VTAIL.n614 0.388379
R2441 VTAIL.n30 VTAIL.n28 0.388379
R2442 VTAIL.n76 VTAIL.n75 0.388379
R2443 VTAIL.n79 VTAIL.n6 0.388379
R2444 VTAIL.n116 VTAIL.n114 0.388379
R2445 VTAIL.n162 VTAIL.n161 0.388379
R2446 VTAIL.n165 VTAIL.n92 0.388379
R2447 VTAIL.n204 VTAIL.n202 0.388379
R2448 VTAIL.n250 VTAIL.n249 0.388379
R2449 VTAIL.n253 VTAIL.n180 0.388379
R2450 VTAIL.n601 VTAIL.n528 0.388379
R2451 VTAIL.n598 VTAIL.n530 0.388379
R2452 VTAIL.n554 VTAIL.n552 0.388379
R2453 VTAIL.n513 VTAIL.n440 0.388379
R2454 VTAIL.n510 VTAIL.n442 0.388379
R2455 VTAIL.n466 VTAIL.n464 0.388379
R2456 VTAIL.n427 VTAIL.n354 0.388379
R2457 VTAIL.n424 VTAIL.n356 0.388379
R2458 VTAIL.n380 VTAIL.n378 0.388379
R2459 VTAIL.n339 VTAIL.n266 0.388379
R2460 VTAIL.n336 VTAIL.n268 0.388379
R2461 VTAIL.n292 VTAIL.n290 0.388379
R2462 VTAIL.n643 VTAIL.n635 0.155672
R2463 VTAIL.n644 VTAIL.n643 0.155672
R2464 VTAIL.n644 VTAIL.n631 0.155672
R2465 VTAIL.n651 VTAIL.n631 0.155672
R2466 VTAIL.n652 VTAIL.n651 0.155672
R2467 VTAIL.n652 VTAIL.n627 0.155672
R2468 VTAIL.n659 VTAIL.n627 0.155672
R2469 VTAIL.n660 VTAIL.n659 0.155672
R2470 VTAIL.n660 VTAIL.n623 0.155672
R2471 VTAIL.n667 VTAIL.n623 0.155672
R2472 VTAIL.n668 VTAIL.n667 0.155672
R2473 VTAIL.n668 VTAIL.n619 0.155672
R2474 VTAIL.n675 VTAIL.n619 0.155672
R2475 VTAIL.n676 VTAIL.n675 0.155672
R2476 VTAIL.n676 VTAIL.n615 0.155672
R2477 VTAIL.n685 VTAIL.n615 0.155672
R2478 VTAIL.n686 VTAIL.n685 0.155672
R2479 VTAIL.n686 VTAIL.n611 0.155672
R2480 VTAIL.n693 VTAIL.n611 0.155672
R2481 VTAIL.n35 VTAIL.n27 0.155672
R2482 VTAIL.n36 VTAIL.n35 0.155672
R2483 VTAIL.n36 VTAIL.n23 0.155672
R2484 VTAIL.n43 VTAIL.n23 0.155672
R2485 VTAIL.n44 VTAIL.n43 0.155672
R2486 VTAIL.n44 VTAIL.n19 0.155672
R2487 VTAIL.n51 VTAIL.n19 0.155672
R2488 VTAIL.n52 VTAIL.n51 0.155672
R2489 VTAIL.n52 VTAIL.n15 0.155672
R2490 VTAIL.n59 VTAIL.n15 0.155672
R2491 VTAIL.n60 VTAIL.n59 0.155672
R2492 VTAIL.n60 VTAIL.n11 0.155672
R2493 VTAIL.n67 VTAIL.n11 0.155672
R2494 VTAIL.n68 VTAIL.n67 0.155672
R2495 VTAIL.n68 VTAIL.n7 0.155672
R2496 VTAIL.n77 VTAIL.n7 0.155672
R2497 VTAIL.n78 VTAIL.n77 0.155672
R2498 VTAIL.n78 VTAIL.n3 0.155672
R2499 VTAIL.n85 VTAIL.n3 0.155672
R2500 VTAIL.n121 VTAIL.n113 0.155672
R2501 VTAIL.n122 VTAIL.n121 0.155672
R2502 VTAIL.n122 VTAIL.n109 0.155672
R2503 VTAIL.n129 VTAIL.n109 0.155672
R2504 VTAIL.n130 VTAIL.n129 0.155672
R2505 VTAIL.n130 VTAIL.n105 0.155672
R2506 VTAIL.n137 VTAIL.n105 0.155672
R2507 VTAIL.n138 VTAIL.n137 0.155672
R2508 VTAIL.n138 VTAIL.n101 0.155672
R2509 VTAIL.n145 VTAIL.n101 0.155672
R2510 VTAIL.n146 VTAIL.n145 0.155672
R2511 VTAIL.n146 VTAIL.n97 0.155672
R2512 VTAIL.n153 VTAIL.n97 0.155672
R2513 VTAIL.n154 VTAIL.n153 0.155672
R2514 VTAIL.n154 VTAIL.n93 0.155672
R2515 VTAIL.n163 VTAIL.n93 0.155672
R2516 VTAIL.n164 VTAIL.n163 0.155672
R2517 VTAIL.n164 VTAIL.n89 0.155672
R2518 VTAIL.n171 VTAIL.n89 0.155672
R2519 VTAIL.n209 VTAIL.n201 0.155672
R2520 VTAIL.n210 VTAIL.n209 0.155672
R2521 VTAIL.n210 VTAIL.n197 0.155672
R2522 VTAIL.n217 VTAIL.n197 0.155672
R2523 VTAIL.n218 VTAIL.n217 0.155672
R2524 VTAIL.n218 VTAIL.n193 0.155672
R2525 VTAIL.n225 VTAIL.n193 0.155672
R2526 VTAIL.n226 VTAIL.n225 0.155672
R2527 VTAIL.n226 VTAIL.n189 0.155672
R2528 VTAIL.n233 VTAIL.n189 0.155672
R2529 VTAIL.n234 VTAIL.n233 0.155672
R2530 VTAIL.n234 VTAIL.n185 0.155672
R2531 VTAIL.n241 VTAIL.n185 0.155672
R2532 VTAIL.n242 VTAIL.n241 0.155672
R2533 VTAIL.n242 VTAIL.n181 0.155672
R2534 VTAIL.n251 VTAIL.n181 0.155672
R2535 VTAIL.n252 VTAIL.n251 0.155672
R2536 VTAIL.n252 VTAIL.n177 0.155672
R2537 VTAIL.n259 VTAIL.n177 0.155672
R2538 VTAIL.n607 VTAIL.n525 0.155672
R2539 VTAIL.n600 VTAIL.n525 0.155672
R2540 VTAIL.n600 VTAIL.n599 0.155672
R2541 VTAIL.n599 VTAIL.n529 0.155672
R2542 VTAIL.n592 VTAIL.n529 0.155672
R2543 VTAIL.n592 VTAIL.n591 0.155672
R2544 VTAIL.n591 VTAIL.n535 0.155672
R2545 VTAIL.n584 VTAIL.n535 0.155672
R2546 VTAIL.n584 VTAIL.n583 0.155672
R2547 VTAIL.n583 VTAIL.n539 0.155672
R2548 VTAIL.n576 VTAIL.n539 0.155672
R2549 VTAIL.n576 VTAIL.n575 0.155672
R2550 VTAIL.n575 VTAIL.n543 0.155672
R2551 VTAIL.n568 VTAIL.n543 0.155672
R2552 VTAIL.n568 VTAIL.n567 0.155672
R2553 VTAIL.n567 VTAIL.n547 0.155672
R2554 VTAIL.n560 VTAIL.n547 0.155672
R2555 VTAIL.n560 VTAIL.n559 0.155672
R2556 VTAIL.n559 VTAIL.n551 0.155672
R2557 VTAIL.n519 VTAIL.n437 0.155672
R2558 VTAIL.n512 VTAIL.n437 0.155672
R2559 VTAIL.n512 VTAIL.n511 0.155672
R2560 VTAIL.n511 VTAIL.n441 0.155672
R2561 VTAIL.n504 VTAIL.n441 0.155672
R2562 VTAIL.n504 VTAIL.n503 0.155672
R2563 VTAIL.n503 VTAIL.n447 0.155672
R2564 VTAIL.n496 VTAIL.n447 0.155672
R2565 VTAIL.n496 VTAIL.n495 0.155672
R2566 VTAIL.n495 VTAIL.n451 0.155672
R2567 VTAIL.n488 VTAIL.n451 0.155672
R2568 VTAIL.n488 VTAIL.n487 0.155672
R2569 VTAIL.n487 VTAIL.n455 0.155672
R2570 VTAIL.n480 VTAIL.n455 0.155672
R2571 VTAIL.n480 VTAIL.n479 0.155672
R2572 VTAIL.n479 VTAIL.n459 0.155672
R2573 VTAIL.n472 VTAIL.n459 0.155672
R2574 VTAIL.n472 VTAIL.n471 0.155672
R2575 VTAIL.n471 VTAIL.n463 0.155672
R2576 VTAIL.n433 VTAIL.n351 0.155672
R2577 VTAIL.n426 VTAIL.n351 0.155672
R2578 VTAIL.n426 VTAIL.n425 0.155672
R2579 VTAIL.n425 VTAIL.n355 0.155672
R2580 VTAIL.n418 VTAIL.n355 0.155672
R2581 VTAIL.n418 VTAIL.n417 0.155672
R2582 VTAIL.n417 VTAIL.n361 0.155672
R2583 VTAIL.n410 VTAIL.n361 0.155672
R2584 VTAIL.n410 VTAIL.n409 0.155672
R2585 VTAIL.n409 VTAIL.n365 0.155672
R2586 VTAIL.n402 VTAIL.n365 0.155672
R2587 VTAIL.n402 VTAIL.n401 0.155672
R2588 VTAIL.n401 VTAIL.n369 0.155672
R2589 VTAIL.n394 VTAIL.n369 0.155672
R2590 VTAIL.n394 VTAIL.n393 0.155672
R2591 VTAIL.n393 VTAIL.n373 0.155672
R2592 VTAIL.n386 VTAIL.n373 0.155672
R2593 VTAIL.n386 VTAIL.n385 0.155672
R2594 VTAIL.n385 VTAIL.n377 0.155672
R2595 VTAIL.n345 VTAIL.n263 0.155672
R2596 VTAIL.n338 VTAIL.n263 0.155672
R2597 VTAIL.n338 VTAIL.n337 0.155672
R2598 VTAIL.n337 VTAIL.n267 0.155672
R2599 VTAIL.n330 VTAIL.n267 0.155672
R2600 VTAIL.n330 VTAIL.n329 0.155672
R2601 VTAIL.n329 VTAIL.n273 0.155672
R2602 VTAIL.n322 VTAIL.n273 0.155672
R2603 VTAIL.n322 VTAIL.n321 0.155672
R2604 VTAIL.n321 VTAIL.n277 0.155672
R2605 VTAIL.n314 VTAIL.n277 0.155672
R2606 VTAIL.n314 VTAIL.n313 0.155672
R2607 VTAIL.n313 VTAIL.n281 0.155672
R2608 VTAIL.n306 VTAIL.n281 0.155672
R2609 VTAIL.n306 VTAIL.n305 0.155672
R2610 VTAIL.n305 VTAIL.n285 0.155672
R2611 VTAIL.n298 VTAIL.n285 0.155672
R2612 VTAIL.n298 VTAIL.n297 0.155672
R2613 VTAIL.n297 VTAIL.n289 0.155672
R2614 VTAIL VTAIL.n1 0.0586897
R2615 VDD1 VDD1.n0 74.7599
R2616 VDD1.n3 VDD1.n2 74.6462
R2617 VDD1.n3 VDD1.n1 74.6462
R2618 VDD1.n5 VDD1.n4 73.167
R2619 VDD1.n5 VDD1.n3 51.4793
R2620 VDD1.n4 VDD1.t4 2.09624
R2621 VDD1.n4 VDD1.t5 2.09624
R2622 VDD1.n0 VDD1.t1 2.09624
R2623 VDD1.n0 VDD1.t3 2.09624
R2624 VDD1.n2 VDD1.t0 2.09624
R2625 VDD1.n2 VDD1.t6 2.09624
R2626 VDD1.n1 VDD1.t2 2.09624
R2627 VDD1.n1 VDD1.t7 2.09624
R2628 VDD1 VDD1.n5 1.47679
R2629 VN.n64 VN.n63 161.3
R2630 VN.n62 VN.n34 161.3
R2631 VN.n61 VN.n60 161.3
R2632 VN.n59 VN.n35 161.3
R2633 VN.n58 VN.n57 161.3
R2634 VN.n56 VN.n36 161.3
R2635 VN.n55 VN.n54 161.3
R2636 VN.n53 VN.n52 161.3
R2637 VN.n51 VN.n38 161.3
R2638 VN.n50 VN.n49 161.3
R2639 VN.n48 VN.n39 161.3
R2640 VN.n47 VN.n46 161.3
R2641 VN.n45 VN.n40 161.3
R2642 VN.n44 VN.n43 161.3
R2643 VN.n31 VN.n30 161.3
R2644 VN.n29 VN.n1 161.3
R2645 VN.n28 VN.n27 161.3
R2646 VN.n26 VN.n2 161.3
R2647 VN.n25 VN.n24 161.3
R2648 VN.n23 VN.n3 161.3
R2649 VN.n22 VN.n21 161.3
R2650 VN.n20 VN.n19 161.3
R2651 VN.n18 VN.n5 161.3
R2652 VN.n17 VN.n16 161.3
R2653 VN.n15 VN.n6 161.3
R2654 VN.n14 VN.n13 161.3
R2655 VN.n12 VN.n7 161.3
R2656 VN.n11 VN.n10 161.3
R2657 VN.n42 VN.t3 148.882
R2658 VN.n9 VN.t1 148.882
R2659 VN.n8 VN.t6 115.725
R2660 VN.n4 VN.t0 115.725
R2661 VN.n0 VN.t7 115.725
R2662 VN.n41 VN.t4 115.725
R2663 VN.n37 VN.t5 115.725
R2664 VN.n33 VN.t2 115.725
R2665 VN.n32 VN.n0 73.4298
R2666 VN.n65 VN.n33 73.4298
R2667 VN.n9 VN.n8 60.5173
R2668 VN.n42 VN.n41 60.5173
R2669 VN VN.n65 56.7935
R2670 VN.n28 VN.n2 46.321
R2671 VN.n61 VN.n35 46.321
R2672 VN.n13 VN.n6 40.4934
R2673 VN.n17 VN.n6 40.4934
R2674 VN.n46 VN.n39 40.4934
R2675 VN.n50 VN.n39 40.4934
R2676 VN.n24 VN.n2 34.6658
R2677 VN.n57 VN.n35 34.6658
R2678 VN.n12 VN.n11 24.4675
R2679 VN.n13 VN.n12 24.4675
R2680 VN.n18 VN.n17 24.4675
R2681 VN.n19 VN.n18 24.4675
R2682 VN.n23 VN.n22 24.4675
R2683 VN.n24 VN.n23 24.4675
R2684 VN.n29 VN.n28 24.4675
R2685 VN.n30 VN.n29 24.4675
R2686 VN.n46 VN.n45 24.4675
R2687 VN.n45 VN.n44 24.4675
R2688 VN.n57 VN.n56 24.4675
R2689 VN.n56 VN.n55 24.4675
R2690 VN.n52 VN.n51 24.4675
R2691 VN.n51 VN.n50 24.4675
R2692 VN.n63 VN.n62 24.4675
R2693 VN.n62 VN.n61 24.4675
R2694 VN.n30 VN.n0 16.6381
R2695 VN.n63 VN.n33 16.6381
R2696 VN.n11 VN.n8 13.702
R2697 VN.n19 VN.n4 13.702
R2698 VN.n44 VN.n41 13.702
R2699 VN.n52 VN.n37 13.702
R2700 VN.n22 VN.n4 10.766
R2701 VN.n55 VN.n37 10.766
R2702 VN.n43 VN.n42 4.06451
R2703 VN.n10 VN.n9 4.06451
R2704 VN.n65 VN.n64 0.354971
R2705 VN.n32 VN.n31 0.354971
R2706 VN VN.n32 0.26696
R2707 VN.n64 VN.n34 0.189894
R2708 VN.n60 VN.n34 0.189894
R2709 VN.n60 VN.n59 0.189894
R2710 VN.n59 VN.n58 0.189894
R2711 VN.n58 VN.n36 0.189894
R2712 VN.n54 VN.n36 0.189894
R2713 VN.n54 VN.n53 0.189894
R2714 VN.n53 VN.n38 0.189894
R2715 VN.n49 VN.n38 0.189894
R2716 VN.n49 VN.n48 0.189894
R2717 VN.n48 VN.n47 0.189894
R2718 VN.n47 VN.n40 0.189894
R2719 VN.n43 VN.n40 0.189894
R2720 VN.n10 VN.n7 0.189894
R2721 VN.n14 VN.n7 0.189894
R2722 VN.n15 VN.n14 0.189894
R2723 VN.n16 VN.n15 0.189894
R2724 VN.n16 VN.n5 0.189894
R2725 VN.n20 VN.n5 0.189894
R2726 VN.n21 VN.n20 0.189894
R2727 VN.n21 VN.n3 0.189894
R2728 VN.n25 VN.n3 0.189894
R2729 VN.n26 VN.n25 0.189894
R2730 VN.n27 VN.n26 0.189894
R2731 VN.n27 VN.n1 0.189894
R2732 VN.n31 VN.n1 0.189894
R2733 VDD2.n2 VDD2.n1 74.6462
R2734 VDD2.n2 VDD2.n0 74.6462
R2735 VDD2 VDD2.n5 74.6433
R2736 VDD2.n4 VDD2.n3 73.1672
R2737 VDD2.n4 VDD2.n2 50.8963
R2738 VDD2.n5 VDD2.t3 2.09624
R2739 VDD2.n5 VDD2.t4 2.09624
R2740 VDD2.n3 VDD2.t5 2.09624
R2741 VDD2.n3 VDD2.t2 2.09624
R2742 VDD2.n1 VDD2.t7 2.09624
R2743 VDD2.n1 VDD2.t0 2.09624
R2744 VDD2.n0 VDD2.t6 2.09624
R2745 VDD2.n0 VDD2.t1 2.09624
R2746 VDD2 VDD2.n4 1.59317
C0 VDD1 VDD2 2.10379f
C1 B VP 2.40539f
C2 B w_n4530_n4070# 12.064f
C3 VTAIL B 6.44301f
C4 VP w_n4530_n4070# 10.0561f
C5 VTAIL VP 12.0081f
C6 VN B 1.41308f
C7 VTAIL w_n4530_n4070# 5.03247f
C8 VN VP 9.08396f
C9 VN w_n4530_n4070# 9.46612f
C10 VN VTAIL 11.994f
C11 B VDD1 1.93587f
C12 B VDD2 2.05172f
C13 VP VDD1 11.981f
C14 VDD1 w_n4530_n4070# 2.2481f
C15 VTAIL VDD1 9.34485f
C16 VP VDD2 0.586448f
C17 VDD2 w_n4530_n4070# 2.38923f
C18 VTAIL VDD2 9.40349f
C19 VN VDD1 0.152606f
C20 VN VDD2 11.548901f
C21 VDD2 VSUBS 2.347898f
C22 VDD1 VSUBS 2.99946f
C23 VTAIL VSUBS 1.600494f
C24 VN VSUBS 7.695879f
C25 VP VSUBS 4.364876f
C26 B VSUBS 6.003489f
C27 w_n4530_n4070# VSUBS 0.225975p
C28 VDD2.t6 VSUBS 0.388316f
C29 VDD2.t1 VSUBS 0.388316f
C30 VDD2.n0 VSUBS 3.20033f
C31 VDD2.t7 VSUBS 0.388316f
C32 VDD2.t0 VSUBS 0.388316f
C33 VDD2.n1 VSUBS 3.20033f
C34 VDD2.n2 VSUBS 5.56031f
C35 VDD2.t5 VSUBS 0.388316f
C36 VDD2.t2 VSUBS 0.388316f
C37 VDD2.n3 VSUBS 3.17907f
C38 VDD2.n4 VSUBS 4.68785f
C39 VDD2.t3 VSUBS 0.388316f
C40 VDD2.t4 VSUBS 0.388316f
C41 VDD2.n5 VSUBS 3.20028f
C42 VN.t7 VSUBS 3.29408f
C43 VN.n0 VSUBS 1.23977f
C44 VN.n1 VSUBS 0.023978f
C45 VN.n2 VSUBS 0.020516f
C46 VN.n3 VSUBS 0.023978f
C47 VN.t0 VSUBS 3.29408f
C48 VN.n4 VSUBS 1.14421f
C49 VN.n5 VSUBS 0.023978f
C50 VN.n6 VSUBS 0.019384f
C51 VN.n7 VSUBS 0.023978f
C52 VN.t6 VSUBS 3.29408f
C53 VN.n8 VSUBS 1.22467f
C54 VN.t1 VSUBS 3.58704f
C55 VN.n9 VSUBS 1.17293f
C56 VN.n10 VSUBS 0.278853f
C57 VN.n11 VSUBS 0.034981f
C58 VN.n12 VSUBS 0.044689f
C59 VN.n13 VSUBS 0.047656f
C60 VN.n14 VSUBS 0.023978f
C61 VN.n15 VSUBS 0.023978f
C62 VN.n16 VSUBS 0.023978f
C63 VN.n17 VSUBS 0.047656f
C64 VN.n18 VSUBS 0.044689f
C65 VN.n19 VSUBS 0.034981f
C66 VN.n20 VSUBS 0.023978f
C67 VN.n21 VSUBS 0.023978f
C68 VN.n22 VSUBS 0.032334f
C69 VN.n23 VSUBS 0.044689f
C70 VN.n24 VSUBS 0.048452f
C71 VN.n25 VSUBS 0.023978f
C72 VN.n26 VSUBS 0.023978f
C73 VN.n27 VSUBS 0.023978f
C74 VN.n28 VSUBS 0.045728f
C75 VN.n29 VSUBS 0.044689f
C76 VN.n30 VSUBS 0.037629f
C77 VN.n31 VSUBS 0.0387f
C78 VN.n32 VSUBS 0.055411f
C79 VN.t2 VSUBS 3.29408f
C80 VN.n33 VSUBS 1.23977f
C81 VN.n34 VSUBS 0.023978f
C82 VN.n35 VSUBS 0.020516f
C83 VN.n36 VSUBS 0.023978f
C84 VN.t5 VSUBS 3.29408f
C85 VN.n37 VSUBS 1.14421f
C86 VN.n38 VSUBS 0.023978f
C87 VN.n39 VSUBS 0.019384f
C88 VN.n40 VSUBS 0.023978f
C89 VN.t4 VSUBS 3.29408f
C90 VN.n41 VSUBS 1.22467f
C91 VN.t3 VSUBS 3.58704f
C92 VN.n42 VSUBS 1.17293f
C93 VN.n43 VSUBS 0.278853f
C94 VN.n44 VSUBS 0.034981f
C95 VN.n45 VSUBS 0.044689f
C96 VN.n46 VSUBS 0.047656f
C97 VN.n47 VSUBS 0.023978f
C98 VN.n48 VSUBS 0.023978f
C99 VN.n49 VSUBS 0.023978f
C100 VN.n50 VSUBS 0.047656f
C101 VN.n51 VSUBS 0.044689f
C102 VN.n52 VSUBS 0.034981f
C103 VN.n53 VSUBS 0.023978f
C104 VN.n54 VSUBS 0.023978f
C105 VN.n55 VSUBS 0.032334f
C106 VN.n56 VSUBS 0.044689f
C107 VN.n57 VSUBS 0.048452f
C108 VN.n58 VSUBS 0.023978f
C109 VN.n59 VSUBS 0.023978f
C110 VN.n60 VSUBS 0.023978f
C111 VN.n61 VSUBS 0.045728f
C112 VN.n62 VSUBS 0.044689f
C113 VN.n63 VSUBS 0.037629f
C114 VN.n64 VSUBS 0.0387f
C115 VN.n65 VSUBS 1.63073f
C116 VDD1.t1 VSUBS 0.359955f
C117 VDD1.t3 VSUBS 0.359955f
C118 VDD1.n0 VSUBS 2.96831f
C119 VDD1.t2 VSUBS 0.359955f
C120 VDD1.t7 VSUBS 0.359955f
C121 VDD1.n1 VSUBS 2.9666f
C122 VDD1.t0 VSUBS 0.359955f
C123 VDD1.t6 VSUBS 0.359955f
C124 VDD1.n2 VSUBS 2.9666f
C125 VDD1.n3 VSUBS 5.21483f
C126 VDD1.t4 VSUBS 0.359955f
C127 VDD1.t5 VSUBS 0.359955f
C128 VDD1.n4 VSUBS 2.94687f
C129 VDD1.n5 VSUBS 4.38232f
C130 VTAIL.t5 VSUBS 0.30008f
C131 VTAIL.t3 VSUBS 0.30008f
C132 VTAIL.n0 VSUBS 2.32197f
C133 VTAIL.n1 VSUBS 0.809063f
C134 VTAIL.n2 VSUBS 0.026696f
C135 VTAIL.n3 VSUBS 0.024483f
C136 VTAIL.n4 VSUBS 0.013156f
C137 VTAIL.n5 VSUBS 0.031097f
C138 VTAIL.n6 VSUBS 0.013543f
C139 VTAIL.n7 VSUBS 0.024483f
C140 VTAIL.n8 VSUBS 0.01393f
C141 VTAIL.n9 VSUBS 0.031097f
C142 VTAIL.n10 VSUBS 0.01393f
C143 VTAIL.n11 VSUBS 0.024483f
C144 VTAIL.n12 VSUBS 0.013156f
C145 VTAIL.n13 VSUBS 0.031097f
C146 VTAIL.n14 VSUBS 0.01393f
C147 VTAIL.n15 VSUBS 0.024483f
C148 VTAIL.n16 VSUBS 0.013156f
C149 VTAIL.n17 VSUBS 0.031097f
C150 VTAIL.n18 VSUBS 0.01393f
C151 VTAIL.n19 VSUBS 0.024483f
C152 VTAIL.n20 VSUBS 0.013156f
C153 VTAIL.n21 VSUBS 0.031097f
C154 VTAIL.n22 VSUBS 0.01393f
C155 VTAIL.n23 VSUBS 0.024483f
C156 VTAIL.n24 VSUBS 0.013156f
C157 VTAIL.n25 VSUBS 0.031097f
C158 VTAIL.n26 VSUBS 0.01393f
C159 VTAIL.n27 VSUBS 1.62f
C160 VTAIL.n28 VSUBS 0.013156f
C161 VTAIL.t2 VSUBS 0.066603f
C162 VTAIL.n29 VSUBS 0.17627f
C163 VTAIL.n30 VSUBS 0.019782f
C164 VTAIL.n31 VSUBS 0.023323f
C165 VTAIL.n32 VSUBS 0.031097f
C166 VTAIL.n33 VSUBS 0.01393f
C167 VTAIL.n34 VSUBS 0.013156f
C168 VTAIL.n35 VSUBS 0.024483f
C169 VTAIL.n36 VSUBS 0.024483f
C170 VTAIL.n37 VSUBS 0.013156f
C171 VTAIL.n38 VSUBS 0.01393f
C172 VTAIL.n39 VSUBS 0.031097f
C173 VTAIL.n40 VSUBS 0.031097f
C174 VTAIL.n41 VSUBS 0.01393f
C175 VTAIL.n42 VSUBS 0.013156f
C176 VTAIL.n43 VSUBS 0.024483f
C177 VTAIL.n44 VSUBS 0.024483f
C178 VTAIL.n45 VSUBS 0.013156f
C179 VTAIL.n46 VSUBS 0.01393f
C180 VTAIL.n47 VSUBS 0.031097f
C181 VTAIL.n48 VSUBS 0.031097f
C182 VTAIL.n49 VSUBS 0.01393f
C183 VTAIL.n50 VSUBS 0.013156f
C184 VTAIL.n51 VSUBS 0.024483f
C185 VTAIL.n52 VSUBS 0.024483f
C186 VTAIL.n53 VSUBS 0.013156f
C187 VTAIL.n54 VSUBS 0.01393f
C188 VTAIL.n55 VSUBS 0.031097f
C189 VTAIL.n56 VSUBS 0.031097f
C190 VTAIL.n57 VSUBS 0.01393f
C191 VTAIL.n58 VSUBS 0.013156f
C192 VTAIL.n59 VSUBS 0.024483f
C193 VTAIL.n60 VSUBS 0.024483f
C194 VTAIL.n61 VSUBS 0.013156f
C195 VTAIL.n62 VSUBS 0.01393f
C196 VTAIL.n63 VSUBS 0.031097f
C197 VTAIL.n64 VSUBS 0.031097f
C198 VTAIL.n65 VSUBS 0.01393f
C199 VTAIL.n66 VSUBS 0.013156f
C200 VTAIL.n67 VSUBS 0.024483f
C201 VTAIL.n68 VSUBS 0.024483f
C202 VTAIL.n69 VSUBS 0.013156f
C203 VTAIL.n70 VSUBS 0.013156f
C204 VTAIL.n71 VSUBS 0.01393f
C205 VTAIL.n72 VSUBS 0.031097f
C206 VTAIL.n73 VSUBS 0.031097f
C207 VTAIL.n74 VSUBS 0.031097f
C208 VTAIL.n75 VSUBS 0.013543f
C209 VTAIL.n76 VSUBS 0.013156f
C210 VTAIL.n77 VSUBS 0.024483f
C211 VTAIL.n78 VSUBS 0.024483f
C212 VTAIL.n79 VSUBS 0.013156f
C213 VTAIL.n80 VSUBS 0.01393f
C214 VTAIL.n81 VSUBS 0.031097f
C215 VTAIL.n82 VSUBS 0.07458f
C216 VTAIL.n83 VSUBS 0.01393f
C217 VTAIL.n84 VSUBS 0.013156f
C218 VTAIL.n85 VSUBS 0.061609f
C219 VTAIL.n86 VSUBS 0.037623f
C220 VTAIL.n87 VSUBS 0.302927f
C221 VTAIL.n88 VSUBS 0.026696f
C222 VTAIL.n89 VSUBS 0.024483f
C223 VTAIL.n90 VSUBS 0.013156f
C224 VTAIL.n91 VSUBS 0.031097f
C225 VTAIL.n92 VSUBS 0.013543f
C226 VTAIL.n93 VSUBS 0.024483f
C227 VTAIL.n94 VSUBS 0.01393f
C228 VTAIL.n95 VSUBS 0.031097f
C229 VTAIL.n96 VSUBS 0.01393f
C230 VTAIL.n97 VSUBS 0.024483f
C231 VTAIL.n98 VSUBS 0.013156f
C232 VTAIL.n99 VSUBS 0.031097f
C233 VTAIL.n100 VSUBS 0.01393f
C234 VTAIL.n101 VSUBS 0.024483f
C235 VTAIL.n102 VSUBS 0.013156f
C236 VTAIL.n103 VSUBS 0.031097f
C237 VTAIL.n104 VSUBS 0.01393f
C238 VTAIL.n105 VSUBS 0.024483f
C239 VTAIL.n106 VSUBS 0.013156f
C240 VTAIL.n107 VSUBS 0.031097f
C241 VTAIL.n108 VSUBS 0.01393f
C242 VTAIL.n109 VSUBS 0.024483f
C243 VTAIL.n110 VSUBS 0.013156f
C244 VTAIL.n111 VSUBS 0.031097f
C245 VTAIL.n112 VSUBS 0.01393f
C246 VTAIL.n113 VSUBS 1.62f
C247 VTAIL.n114 VSUBS 0.013156f
C248 VTAIL.t9 VSUBS 0.066603f
C249 VTAIL.n115 VSUBS 0.17627f
C250 VTAIL.n116 VSUBS 0.019782f
C251 VTAIL.n117 VSUBS 0.023323f
C252 VTAIL.n118 VSUBS 0.031097f
C253 VTAIL.n119 VSUBS 0.01393f
C254 VTAIL.n120 VSUBS 0.013156f
C255 VTAIL.n121 VSUBS 0.024483f
C256 VTAIL.n122 VSUBS 0.024483f
C257 VTAIL.n123 VSUBS 0.013156f
C258 VTAIL.n124 VSUBS 0.01393f
C259 VTAIL.n125 VSUBS 0.031097f
C260 VTAIL.n126 VSUBS 0.031097f
C261 VTAIL.n127 VSUBS 0.01393f
C262 VTAIL.n128 VSUBS 0.013156f
C263 VTAIL.n129 VSUBS 0.024483f
C264 VTAIL.n130 VSUBS 0.024483f
C265 VTAIL.n131 VSUBS 0.013156f
C266 VTAIL.n132 VSUBS 0.01393f
C267 VTAIL.n133 VSUBS 0.031097f
C268 VTAIL.n134 VSUBS 0.031097f
C269 VTAIL.n135 VSUBS 0.01393f
C270 VTAIL.n136 VSUBS 0.013156f
C271 VTAIL.n137 VSUBS 0.024483f
C272 VTAIL.n138 VSUBS 0.024483f
C273 VTAIL.n139 VSUBS 0.013156f
C274 VTAIL.n140 VSUBS 0.01393f
C275 VTAIL.n141 VSUBS 0.031097f
C276 VTAIL.n142 VSUBS 0.031097f
C277 VTAIL.n143 VSUBS 0.01393f
C278 VTAIL.n144 VSUBS 0.013156f
C279 VTAIL.n145 VSUBS 0.024483f
C280 VTAIL.n146 VSUBS 0.024483f
C281 VTAIL.n147 VSUBS 0.013156f
C282 VTAIL.n148 VSUBS 0.01393f
C283 VTAIL.n149 VSUBS 0.031097f
C284 VTAIL.n150 VSUBS 0.031097f
C285 VTAIL.n151 VSUBS 0.01393f
C286 VTAIL.n152 VSUBS 0.013156f
C287 VTAIL.n153 VSUBS 0.024483f
C288 VTAIL.n154 VSUBS 0.024483f
C289 VTAIL.n155 VSUBS 0.013156f
C290 VTAIL.n156 VSUBS 0.013156f
C291 VTAIL.n157 VSUBS 0.01393f
C292 VTAIL.n158 VSUBS 0.031097f
C293 VTAIL.n159 VSUBS 0.031097f
C294 VTAIL.n160 VSUBS 0.031097f
C295 VTAIL.n161 VSUBS 0.013543f
C296 VTAIL.n162 VSUBS 0.013156f
C297 VTAIL.n163 VSUBS 0.024483f
C298 VTAIL.n164 VSUBS 0.024483f
C299 VTAIL.n165 VSUBS 0.013156f
C300 VTAIL.n166 VSUBS 0.01393f
C301 VTAIL.n167 VSUBS 0.031097f
C302 VTAIL.n168 VSUBS 0.07458f
C303 VTAIL.n169 VSUBS 0.01393f
C304 VTAIL.n170 VSUBS 0.013156f
C305 VTAIL.n171 VSUBS 0.061609f
C306 VTAIL.n172 VSUBS 0.037623f
C307 VTAIL.n173 VSUBS 0.302927f
C308 VTAIL.t8 VSUBS 0.30008f
C309 VTAIL.t15 VSUBS 0.30008f
C310 VTAIL.n174 VSUBS 2.32197f
C311 VTAIL.n175 VSUBS 1.04659f
C312 VTAIL.n176 VSUBS 0.026696f
C313 VTAIL.n177 VSUBS 0.024483f
C314 VTAIL.n178 VSUBS 0.013156f
C315 VTAIL.n179 VSUBS 0.031097f
C316 VTAIL.n180 VSUBS 0.013543f
C317 VTAIL.n181 VSUBS 0.024483f
C318 VTAIL.n182 VSUBS 0.01393f
C319 VTAIL.n183 VSUBS 0.031097f
C320 VTAIL.n184 VSUBS 0.01393f
C321 VTAIL.n185 VSUBS 0.024483f
C322 VTAIL.n186 VSUBS 0.013156f
C323 VTAIL.n187 VSUBS 0.031097f
C324 VTAIL.n188 VSUBS 0.01393f
C325 VTAIL.n189 VSUBS 0.024483f
C326 VTAIL.n190 VSUBS 0.013156f
C327 VTAIL.n191 VSUBS 0.031097f
C328 VTAIL.n192 VSUBS 0.01393f
C329 VTAIL.n193 VSUBS 0.024483f
C330 VTAIL.n194 VSUBS 0.013156f
C331 VTAIL.n195 VSUBS 0.031097f
C332 VTAIL.n196 VSUBS 0.01393f
C333 VTAIL.n197 VSUBS 0.024483f
C334 VTAIL.n198 VSUBS 0.013156f
C335 VTAIL.n199 VSUBS 0.031097f
C336 VTAIL.n200 VSUBS 0.01393f
C337 VTAIL.n201 VSUBS 1.62f
C338 VTAIL.n202 VSUBS 0.013156f
C339 VTAIL.t13 VSUBS 0.066603f
C340 VTAIL.n203 VSUBS 0.17627f
C341 VTAIL.n204 VSUBS 0.019782f
C342 VTAIL.n205 VSUBS 0.023323f
C343 VTAIL.n206 VSUBS 0.031097f
C344 VTAIL.n207 VSUBS 0.01393f
C345 VTAIL.n208 VSUBS 0.013156f
C346 VTAIL.n209 VSUBS 0.024483f
C347 VTAIL.n210 VSUBS 0.024483f
C348 VTAIL.n211 VSUBS 0.013156f
C349 VTAIL.n212 VSUBS 0.01393f
C350 VTAIL.n213 VSUBS 0.031097f
C351 VTAIL.n214 VSUBS 0.031097f
C352 VTAIL.n215 VSUBS 0.01393f
C353 VTAIL.n216 VSUBS 0.013156f
C354 VTAIL.n217 VSUBS 0.024483f
C355 VTAIL.n218 VSUBS 0.024483f
C356 VTAIL.n219 VSUBS 0.013156f
C357 VTAIL.n220 VSUBS 0.01393f
C358 VTAIL.n221 VSUBS 0.031097f
C359 VTAIL.n222 VSUBS 0.031097f
C360 VTAIL.n223 VSUBS 0.01393f
C361 VTAIL.n224 VSUBS 0.013156f
C362 VTAIL.n225 VSUBS 0.024483f
C363 VTAIL.n226 VSUBS 0.024483f
C364 VTAIL.n227 VSUBS 0.013156f
C365 VTAIL.n228 VSUBS 0.01393f
C366 VTAIL.n229 VSUBS 0.031097f
C367 VTAIL.n230 VSUBS 0.031097f
C368 VTAIL.n231 VSUBS 0.01393f
C369 VTAIL.n232 VSUBS 0.013156f
C370 VTAIL.n233 VSUBS 0.024483f
C371 VTAIL.n234 VSUBS 0.024483f
C372 VTAIL.n235 VSUBS 0.013156f
C373 VTAIL.n236 VSUBS 0.01393f
C374 VTAIL.n237 VSUBS 0.031097f
C375 VTAIL.n238 VSUBS 0.031097f
C376 VTAIL.n239 VSUBS 0.01393f
C377 VTAIL.n240 VSUBS 0.013156f
C378 VTAIL.n241 VSUBS 0.024483f
C379 VTAIL.n242 VSUBS 0.024483f
C380 VTAIL.n243 VSUBS 0.013156f
C381 VTAIL.n244 VSUBS 0.013156f
C382 VTAIL.n245 VSUBS 0.01393f
C383 VTAIL.n246 VSUBS 0.031097f
C384 VTAIL.n247 VSUBS 0.031097f
C385 VTAIL.n248 VSUBS 0.031097f
C386 VTAIL.n249 VSUBS 0.013543f
C387 VTAIL.n250 VSUBS 0.013156f
C388 VTAIL.n251 VSUBS 0.024483f
C389 VTAIL.n252 VSUBS 0.024483f
C390 VTAIL.n253 VSUBS 0.013156f
C391 VTAIL.n254 VSUBS 0.01393f
C392 VTAIL.n255 VSUBS 0.031097f
C393 VTAIL.n256 VSUBS 0.07458f
C394 VTAIL.n257 VSUBS 0.01393f
C395 VTAIL.n258 VSUBS 0.013156f
C396 VTAIL.n259 VSUBS 0.061609f
C397 VTAIL.n260 VSUBS 0.037623f
C398 VTAIL.n261 VSUBS 1.89538f
C399 VTAIL.n262 VSUBS 0.026696f
C400 VTAIL.n263 VSUBS 0.024483f
C401 VTAIL.n264 VSUBS 0.013156f
C402 VTAIL.n265 VSUBS 0.031097f
C403 VTAIL.n266 VSUBS 0.013543f
C404 VTAIL.n267 VSUBS 0.024483f
C405 VTAIL.n268 VSUBS 0.013543f
C406 VTAIL.n269 VSUBS 0.013156f
C407 VTAIL.n270 VSUBS 0.031097f
C408 VTAIL.n271 VSUBS 0.031097f
C409 VTAIL.n272 VSUBS 0.01393f
C410 VTAIL.n273 VSUBS 0.024483f
C411 VTAIL.n274 VSUBS 0.013156f
C412 VTAIL.n275 VSUBS 0.031097f
C413 VTAIL.n276 VSUBS 0.01393f
C414 VTAIL.n277 VSUBS 0.024483f
C415 VTAIL.n278 VSUBS 0.013156f
C416 VTAIL.n279 VSUBS 0.031097f
C417 VTAIL.n280 VSUBS 0.01393f
C418 VTAIL.n281 VSUBS 0.024483f
C419 VTAIL.n282 VSUBS 0.013156f
C420 VTAIL.n283 VSUBS 0.031097f
C421 VTAIL.n284 VSUBS 0.01393f
C422 VTAIL.n285 VSUBS 0.024483f
C423 VTAIL.n286 VSUBS 0.013156f
C424 VTAIL.n287 VSUBS 0.031097f
C425 VTAIL.n288 VSUBS 0.01393f
C426 VTAIL.n289 VSUBS 1.62f
C427 VTAIL.n290 VSUBS 0.013156f
C428 VTAIL.t6 VSUBS 0.066603f
C429 VTAIL.n291 VSUBS 0.17627f
C430 VTAIL.n292 VSUBS 0.019782f
C431 VTAIL.n293 VSUBS 0.023323f
C432 VTAIL.n294 VSUBS 0.031097f
C433 VTAIL.n295 VSUBS 0.01393f
C434 VTAIL.n296 VSUBS 0.013156f
C435 VTAIL.n297 VSUBS 0.024483f
C436 VTAIL.n298 VSUBS 0.024483f
C437 VTAIL.n299 VSUBS 0.013156f
C438 VTAIL.n300 VSUBS 0.01393f
C439 VTAIL.n301 VSUBS 0.031097f
C440 VTAIL.n302 VSUBS 0.031097f
C441 VTAIL.n303 VSUBS 0.01393f
C442 VTAIL.n304 VSUBS 0.013156f
C443 VTAIL.n305 VSUBS 0.024483f
C444 VTAIL.n306 VSUBS 0.024483f
C445 VTAIL.n307 VSUBS 0.013156f
C446 VTAIL.n308 VSUBS 0.01393f
C447 VTAIL.n309 VSUBS 0.031097f
C448 VTAIL.n310 VSUBS 0.031097f
C449 VTAIL.n311 VSUBS 0.01393f
C450 VTAIL.n312 VSUBS 0.013156f
C451 VTAIL.n313 VSUBS 0.024483f
C452 VTAIL.n314 VSUBS 0.024483f
C453 VTAIL.n315 VSUBS 0.013156f
C454 VTAIL.n316 VSUBS 0.01393f
C455 VTAIL.n317 VSUBS 0.031097f
C456 VTAIL.n318 VSUBS 0.031097f
C457 VTAIL.n319 VSUBS 0.01393f
C458 VTAIL.n320 VSUBS 0.013156f
C459 VTAIL.n321 VSUBS 0.024483f
C460 VTAIL.n322 VSUBS 0.024483f
C461 VTAIL.n323 VSUBS 0.013156f
C462 VTAIL.n324 VSUBS 0.01393f
C463 VTAIL.n325 VSUBS 0.031097f
C464 VTAIL.n326 VSUBS 0.031097f
C465 VTAIL.n327 VSUBS 0.01393f
C466 VTAIL.n328 VSUBS 0.013156f
C467 VTAIL.n329 VSUBS 0.024483f
C468 VTAIL.n330 VSUBS 0.024483f
C469 VTAIL.n331 VSUBS 0.013156f
C470 VTAIL.n332 VSUBS 0.01393f
C471 VTAIL.n333 VSUBS 0.031097f
C472 VTAIL.n334 VSUBS 0.031097f
C473 VTAIL.n335 VSUBS 0.01393f
C474 VTAIL.n336 VSUBS 0.013156f
C475 VTAIL.n337 VSUBS 0.024483f
C476 VTAIL.n338 VSUBS 0.024483f
C477 VTAIL.n339 VSUBS 0.013156f
C478 VTAIL.n340 VSUBS 0.01393f
C479 VTAIL.n341 VSUBS 0.031097f
C480 VTAIL.n342 VSUBS 0.07458f
C481 VTAIL.n343 VSUBS 0.01393f
C482 VTAIL.n344 VSUBS 0.013156f
C483 VTAIL.n345 VSUBS 0.061609f
C484 VTAIL.n346 VSUBS 0.037623f
C485 VTAIL.n347 VSUBS 1.89538f
C486 VTAIL.t0 VSUBS 0.30008f
C487 VTAIL.t7 VSUBS 0.30008f
C488 VTAIL.n348 VSUBS 2.32199f
C489 VTAIL.n349 VSUBS 1.04657f
C490 VTAIL.n350 VSUBS 0.026696f
C491 VTAIL.n351 VSUBS 0.024483f
C492 VTAIL.n352 VSUBS 0.013156f
C493 VTAIL.n353 VSUBS 0.031097f
C494 VTAIL.n354 VSUBS 0.013543f
C495 VTAIL.n355 VSUBS 0.024483f
C496 VTAIL.n356 VSUBS 0.013543f
C497 VTAIL.n357 VSUBS 0.013156f
C498 VTAIL.n358 VSUBS 0.031097f
C499 VTAIL.n359 VSUBS 0.031097f
C500 VTAIL.n360 VSUBS 0.01393f
C501 VTAIL.n361 VSUBS 0.024483f
C502 VTAIL.n362 VSUBS 0.013156f
C503 VTAIL.n363 VSUBS 0.031097f
C504 VTAIL.n364 VSUBS 0.01393f
C505 VTAIL.n365 VSUBS 0.024483f
C506 VTAIL.n366 VSUBS 0.013156f
C507 VTAIL.n367 VSUBS 0.031097f
C508 VTAIL.n368 VSUBS 0.01393f
C509 VTAIL.n369 VSUBS 0.024483f
C510 VTAIL.n370 VSUBS 0.013156f
C511 VTAIL.n371 VSUBS 0.031097f
C512 VTAIL.n372 VSUBS 0.01393f
C513 VTAIL.n373 VSUBS 0.024483f
C514 VTAIL.n374 VSUBS 0.013156f
C515 VTAIL.n375 VSUBS 0.031097f
C516 VTAIL.n376 VSUBS 0.01393f
C517 VTAIL.n377 VSUBS 1.62f
C518 VTAIL.n378 VSUBS 0.013156f
C519 VTAIL.t1 VSUBS 0.066603f
C520 VTAIL.n379 VSUBS 0.17627f
C521 VTAIL.n380 VSUBS 0.019782f
C522 VTAIL.n381 VSUBS 0.023323f
C523 VTAIL.n382 VSUBS 0.031097f
C524 VTAIL.n383 VSUBS 0.01393f
C525 VTAIL.n384 VSUBS 0.013156f
C526 VTAIL.n385 VSUBS 0.024483f
C527 VTAIL.n386 VSUBS 0.024483f
C528 VTAIL.n387 VSUBS 0.013156f
C529 VTAIL.n388 VSUBS 0.01393f
C530 VTAIL.n389 VSUBS 0.031097f
C531 VTAIL.n390 VSUBS 0.031097f
C532 VTAIL.n391 VSUBS 0.01393f
C533 VTAIL.n392 VSUBS 0.013156f
C534 VTAIL.n393 VSUBS 0.024483f
C535 VTAIL.n394 VSUBS 0.024483f
C536 VTAIL.n395 VSUBS 0.013156f
C537 VTAIL.n396 VSUBS 0.01393f
C538 VTAIL.n397 VSUBS 0.031097f
C539 VTAIL.n398 VSUBS 0.031097f
C540 VTAIL.n399 VSUBS 0.01393f
C541 VTAIL.n400 VSUBS 0.013156f
C542 VTAIL.n401 VSUBS 0.024483f
C543 VTAIL.n402 VSUBS 0.024483f
C544 VTAIL.n403 VSUBS 0.013156f
C545 VTAIL.n404 VSUBS 0.01393f
C546 VTAIL.n405 VSUBS 0.031097f
C547 VTAIL.n406 VSUBS 0.031097f
C548 VTAIL.n407 VSUBS 0.01393f
C549 VTAIL.n408 VSUBS 0.013156f
C550 VTAIL.n409 VSUBS 0.024483f
C551 VTAIL.n410 VSUBS 0.024483f
C552 VTAIL.n411 VSUBS 0.013156f
C553 VTAIL.n412 VSUBS 0.01393f
C554 VTAIL.n413 VSUBS 0.031097f
C555 VTAIL.n414 VSUBS 0.031097f
C556 VTAIL.n415 VSUBS 0.01393f
C557 VTAIL.n416 VSUBS 0.013156f
C558 VTAIL.n417 VSUBS 0.024483f
C559 VTAIL.n418 VSUBS 0.024483f
C560 VTAIL.n419 VSUBS 0.013156f
C561 VTAIL.n420 VSUBS 0.01393f
C562 VTAIL.n421 VSUBS 0.031097f
C563 VTAIL.n422 VSUBS 0.031097f
C564 VTAIL.n423 VSUBS 0.01393f
C565 VTAIL.n424 VSUBS 0.013156f
C566 VTAIL.n425 VSUBS 0.024483f
C567 VTAIL.n426 VSUBS 0.024483f
C568 VTAIL.n427 VSUBS 0.013156f
C569 VTAIL.n428 VSUBS 0.01393f
C570 VTAIL.n429 VSUBS 0.031097f
C571 VTAIL.n430 VSUBS 0.07458f
C572 VTAIL.n431 VSUBS 0.01393f
C573 VTAIL.n432 VSUBS 0.013156f
C574 VTAIL.n433 VSUBS 0.061609f
C575 VTAIL.n434 VSUBS 0.037623f
C576 VTAIL.n435 VSUBS 0.302927f
C577 VTAIL.n436 VSUBS 0.026696f
C578 VTAIL.n437 VSUBS 0.024483f
C579 VTAIL.n438 VSUBS 0.013156f
C580 VTAIL.n439 VSUBS 0.031097f
C581 VTAIL.n440 VSUBS 0.013543f
C582 VTAIL.n441 VSUBS 0.024483f
C583 VTAIL.n442 VSUBS 0.013543f
C584 VTAIL.n443 VSUBS 0.013156f
C585 VTAIL.n444 VSUBS 0.031097f
C586 VTAIL.n445 VSUBS 0.031097f
C587 VTAIL.n446 VSUBS 0.01393f
C588 VTAIL.n447 VSUBS 0.024483f
C589 VTAIL.n448 VSUBS 0.013156f
C590 VTAIL.n449 VSUBS 0.031097f
C591 VTAIL.n450 VSUBS 0.01393f
C592 VTAIL.n451 VSUBS 0.024483f
C593 VTAIL.n452 VSUBS 0.013156f
C594 VTAIL.n453 VSUBS 0.031097f
C595 VTAIL.n454 VSUBS 0.01393f
C596 VTAIL.n455 VSUBS 0.024483f
C597 VTAIL.n456 VSUBS 0.013156f
C598 VTAIL.n457 VSUBS 0.031097f
C599 VTAIL.n458 VSUBS 0.01393f
C600 VTAIL.n459 VSUBS 0.024483f
C601 VTAIL.n460 VSUBS 0.013156f
C602 VTAIL.n461 VSUBS 0.031097f
C603 VTAIL.n462 VSUBS 0.01393f
C604 VTAIL.n463 VSUBS 1.62f
C605 VTAIL.n464 VSUBS 0.013156f
C606 VTAIL.t14 VSUBS 0.066603f
C607 VTAIL.n465 VSUBS 0.17627f
C608 VTAIL.n466 VSUBS 0.019782f
C609 VTAIL.n467 VSUBS 0.023323f
C610 VTAIL.n468 VSUBS 0.031097f
C611 VTAIL.n469 VSUBS 0.01393f
C612 VTAIL.n470 VSUBS 0.013156f
C613 VTAIL.n471 VSUBS 0.024483f
C614 VTAIL.n472 VSUBS 0.024483f
C615 VTAIL.n473 VSUBS 0.013156f
C616 VTAIL.n474 VSUBS 0.01393f
C617 VTAIL.n475 VSUBS 0.031097f
C618 VTAIL.n476 VSUBS 0.031097f
C619 VTAIL.n477 VSUBS 0.01393f
C620 VTAIL.n478 VSUBS 0.013156f
C621 VTAIL.n479 VSUBS 0.024483f
C622 VTAIL.n480 VSUBS 0.024483f
C623 VTAIL.n481 VSUBS 0.013156f
C624 VTAIL.n482 VSUBS 0.01393f
C625 VTAIL.n483 VSUBS 0.031097f
C626 VTAIL.n484 VSUBS 0.031097f
C627 VTAIL.n485 VSUBS 0.01393f
C628 VTAIL.n486 VSUBS 0.013156f
C629 VTAIL.n487 VSUBS 0.024483f
C630 VTAIL.n488 VSUBS 0.024483f
C631 VTAIL.n489 VSUBS 0.013156f
C632 VTAIL.n490 VSUBS 0.01393f
C633 VTAIL.n491 VSUBS 0.031097f
C634 VTAIL.n492 VSUBS 0.031097f
C635 VTAIL.n493 VSUBS 0.01393f
C636 VTAIL.n494 VSUBS 0.013156f
C637 VTAIL.n495 VSUBS 0.024483f
C638 VTAIL.n496 VSUBS 0.024483f
C639 VTAIL.n497 VSUBS 0.013156f
C640 VTAIL.n498 VSUBS 0.01393f
C641 VTAIL.n499 VSUBS 0.031097f
C642 VTAIL.n500 VSUBS 0.031097f
C643 VTAIL.n501 VSUBS 0.01393f
C644 VTAIL.n502 VSUBS 0.013156f
C645 VTAIL.n503 VSUBS 0.024483f
C646 VTAIL.n504 VSUBS 0.024483f
C647 VTAIL.n505 VSUBS 0.013156f
C648 VTAIL.n506 VSUBS 0.01393f
C649 VTAIL.n507 VSUBS 0.031097f
C650 VTAIL.n508 VSUBS 0.031097f
C651 VTAIL.n509 VSUBS 0.01393f
C652 VTAIL.n510 VSUBS 0.013156f
C653 VTAIL.n511 VSUBS 0.024483f
C654 VTAIL.n512 VSUBS 0.024483f
C655 VTAIL.n513 VSUBS 0.013156f
C656 VTAIL.n514 VSUBS 0.01393f
C657 VTAIL.n515 VSUBS 0.031097f
C658 VTAIL.n516 VSUBS 0.07458f
C659 VTAIL.n517 VSUBS 0.01393f
C660 VTAIL.n518 VSUBS 0.013156f
C661 VTAIL.n519 VSUBS 0.061609f
C662 VTAIL.n520 VSUBS 0.037623f
C663 VTAIL.n521 VSUBS 0.302927f
C664 VTAIL.t12 VSUBS 0.30008f
C665 VTAIL.t11 VSUBS 0.30008f
C666 VTAIL.n522 VSUBS 2.32199f
C667 VTAIL.n523 VSUBS 1.04657f
C668 VTAIL.n524 VSUBS 0.026696f
C669 VTAIL.n525 VSUBS 0.024483f
C670 VTAIL.n526 VSUBS 0.013156f
C671 VTAIL.n527 VSUBS 0.031097f
C672 VTAIL.n528 VSUBS 0.013543f
C673 VTAIL.n529 VSUBS 0.024483f
C674 VTAIL.n530 VSUBS 0.013543f
C675 VTAIL.n531 VSUBS 0.013156f
C676 VTAIL.n532 VSUBS 0.031097f
C677 VTAIL.n533 VSUBS 0.031097f
C678 VTAIL.n534 VSUBS 0.01393f
C679 VTAIL.n535 VSUBS 0.024483f
C680 VTAIL.n536 VSUBS 0.013156f
C681 VTAIL.n537 VSUBS 0.031097f
C682 VTAIL.n538 VSUBS 0.01393f
C683 VTAIL.n539 VSUBS 0.024483f
C684 VTAIL.n540 VSUBS 0.013156f
C685 VTAIL.n541 VSUBS 0.031097f
C686 VTAIL.n542 VSUBS 0.01393f
C687 VTAIL.n543 VSUBS 0.024483f
C688 VTAIL.n544 VSUBS 0.013156f
C689 VTAIL.n545 VSUBS 0.031097f
C690 VTAIL.n546 VSUBS 0.01393f
C691 VTAIL.n547 VSUBS 0.024483f
C692 VTAIL.n548 VSUBS 0.013156f
C693 VTAIL.n549 VSUBS 0.031097f
C694 VTAIL.n550 VSUBS 0.01393f
C695 VTAIL.n551 VSUBS 1.62f
C696 VTAIL.n552 VSUBS 0.013156f
C697 VTAIL.t10 VSUBS 0.066603f
C698 VTAIL.n553 VSUBS 0.17627f
C699 VTAIL.n554 VSUBS 0.019782f
C700 VTAIL.n555 VSUBS 0.023323f
C701 VTAIL.n556 VSUBS 0.031097f
C702 VTAIL.n557 VSUBS 0.01393f
C703 VTAIL.n558 VSUBS 0.013156f
C704 VTAIL.n559 VSUBS 0.024483f
C705 VTAIL.n560 VSUBS 0.024483f
C706 VTAIL.n561 VSUBS 0.013156f
C707 VTAIL.n562 VSUBS 0.01393f
C708 VTAIL.n563 VSUBS 0.031097f
C709 VTAIL.n564 VSUBS 0.031097f
C710 VTAIL.n565 VSUBS 0.01393f
C711 VTAIL.n566 VSUBS 0.013156f
C712 VTAIL.n567 VSUBS 0.024483f
C713 VTAIL.n568 VSUBS 0.024483f
C714 VTAIL.n569 VSUBS 0.013156f
C715 VTAIL.n570 VSUBS 0.01393f
C716 VTAIL.n571 VSUBS 0.031097f
C717 VTAIL.n572 VSUBS 0.031097f
C718 VTAIL.n573 VSUBS 0.01393f
C719 VTAIL.n574 VSUBS 0.013156f
C720 VTAIL.n575 VSUBS 0.024483f
C721 VTAIL.n576 VSUBS 0.024483f
C722 VTAIL.n577 VSUBS 0.013156f
C723 VTAIL.n578 VSUBS 0.01393f
C724 VTAIL.n579 VSUBS 0.031097f
C725 VTAIL.n580 VSUBS 0.031097f
C726 VTAIL.n581 VSUBS 0.01393f
C727 VTAIL.n582 VSUBS 0.013156f
C728 VTAIL.n583 VSUBS 0.024483f
C729 VTAIL.n584 VSUBS 0.024483f
C730 VTAIL.n585 VSUBS 0.013156f
C731 VTAIL.n586 VSUBS 0.01393f
C732 VTAIL.n587 VSUBS 0.031097f
C733 VTAIL.n588 VSUBS 0.031097f
C734 VTAIL.n589 VSUBS 0.01393f
C735 VTAIL.n590 VSUBS 0.013156f
C736 VTAIL.n591 VSUBS 0.024483f
C737 VTAIL.n592 VSUBS 0.024483f
C738 VTAIL.n593 VSUBS 0.013156f
C739 VTAIL.n594 VSUBS 0.01393f
C740 VTAIL.n595 VSUBS 0.031097f
C741 VTAIL.n596 VSUBS 0.031097f
C742 VTAIL.n597 VSUBS 0.01393f
C743 VTAIL.n598 VSUBS 0.013156f
C744 VTAIL.n599 VSUBS 0.024483f
C745 VTAIL.n600 VSUBS 0.024483f
C746 VTAIL.n601 VSUBS 0.013156f
C747 VTAIL.n602 VSUBS 0.01393f
C748 VTAIL.n603 VSUBS 0.031097f
C749 VTAIL.n604 VSUBS 0.07458f
C750 VTAIL.n605 VSUBS 0.01393f
C751 VTAIL.n606 VSUBS 0.013156f
C752 VTAIL.n607 VSUBS 0.061609f
C753 VTAIL.n608 VSUBS 0.037623f
C754 VTAIL.n609 VSUBS 1.89538f
C755 VTAIL.n610 VSUBS 0.026696f
C756 VTAIL.n611 VSUBS 0.024483f
C757 VTAIL.n612 VSUBS 0.013156f
C758 VTAIL.n613 VSUBS 0.031097f
C759 VTAIL.n614 VSUBS 0.013543f
C760 VTAIL.n615 VSUBS 0.024483f
C761 VTAIL.n616 VSUBS 0.01393f
C762 VTAIL.n617 VSUBS 0.031097f
C763 VTAIL.n618 VSUBS 0.01393f
C764 VTAIL.n619 VSUBS 0.024483f
C765 VTAIL.n620 VSUBS 0.013156f
C766 VTAIL.n621 VSUBS 0.031097f
C767 VTAIL.n622 VSUBS 0.01393f
C768 VTAIL.n623 VSUBS 0.024483f
C769 VTAIL.n624 VSUBS 0.013156f
C770 VTAIL.n625 VSUBS 0.031097f
C771 VTAIL.n626 VSUBS 0.01393f
C772 VTAIL.n627 VSUBS 0.024483f
C773 VTAIL.n628 VSUBS 0.013156f
C774 VTAIL.n629 VSUBS 0.031097f
C775 VTAIL.n630 VSUBS 0.01393f
C776 VTAIL.n631 VSUBS 0.024483f
C777 VTAIL.n632 VSUBS 0.013156f
C778 VTAIL.n633 VSUBS 0.031097f
C779 VTAIL.n634 VSUBS 0.01393f
C780 VTAIL.n635 VSUBS 1.62f
C781 VTAIL.n636 VSUBS 0.013156f
C782 VTAIL.t4 VSUBS 0.066603f
C783 VTAIL.n637 VSUBS 0.17627f
C784 VTAIL.n638 VSUBS 0.019782f
C785 VTAIL.n639 VSUBS 0.023323f
C786 VTAIL.n640 VSUBS 0.031097f
C787 VTAIL.n641 VSUBS 0.01393f
C788 VTAIL.n642 VSUBS 0.013156f
C789 VTAIL.n643 VSUBS 0.024483f
C790 VTAIL.n644 VSUBS 0.024483f
C791 VTAIL.n645 VSUBS 0.013156f
C792 VTAIL.n646 VSUBS 0.01393f
C793 VTAIL.n647 VSUBS 0.031097f
C794 VTAIL.n648 VSUBS 0.031097f
C795 VTAIL.n649 VSUBS 0.01393f
C796 VTAIL.n650 VSUBS 0.013156f
C797 VTAIL.n651 VSUBS 0.024483f
C798 VTAIL.n652 VSUBS 0.024483f
C799 VTAIL.n653 VSUBS 0.013156f
C800 VTAIL.n654 VSUBS 0.01393f
C801 VTAIL.n655 VSUBS 0.031097f
C802 VTAIL.n656 VSUBS 0.031097f
C803 VTAIL.n657 VSUBS 0.01393f
C804 VTAIL.n658 VSUBS 0.013156f
C805 VTAIL.n659 VSUBS 0.024483f
C806 VTAIL.n660 VSUBS 0.024483f
C807 VTAIL.n661 VSUBS 0.013156f
C808 VTAIL.n662 VSUBS 0.01393f
C809 VTAIL.n663 VSUBS 0.031097f
C810 VTAIL.n664 VSUBS 0.031097f
C811 VTAIL.n665 VSUBS 0.01393f
C812 VTAIL.n666 VSUBS 0.013156f
C813 VTAIL.n667 VSUBS 0.024483f
C814 VTAIL.n668 VSUBS 0.024483f
C815 VTAIL.n669 VSUBS 0.013156f
C816 VTAIL.n670 VSUBS 0.01393f
C817 VTAIL.n671 VSUBS 0.031097f
C818 VTAIL.n672 VSUBS 0.031097f
C819 VTAIL.n673 VSUBS 0.01393f
C820 VTAIL.n674 VSUBS 0.013156f
C821 VTAIL.n675 VSUBS 0.024483f
C822 VTAIL.n676 VSUBS 0.024483f
C823 VTAIL.n677 VSUBS 0.013156f
C824 VTAIL.n678 VSUBS 0.013156f
C825 VTAIL.n679 VSUBS 0.01393f
C826 VTAIL.n680 VSUBS 0.031097f
C827 VTAIL.n681 VSUBS 0.031097f
C828 VTAIL.n682 VSUBS 0.031097f
C829 VTAIL.n683 VSUBS 0.013543f
C830 VTAIL.n684 VSUBS 0.013156f
C831 VTAIL.n685 VSUBS 0.024483f
C832 VTAIL.n686 VSUBS 0.024483f
C833 VTAIL.n687 VSUBS 0.013156f
C834 VTAIL.n688 VSUBS 0.01393f
C835 VTAIL.n689 VSUBS 0.031097f
C836 VTAIL.n690 VSUBS 0.07458f
C837 VTAIL.n691 VSUBS 0.01393f
C838 VTAIL.n692 VSUBS 0.013156f
C839 VTAIL.n693 VSUBS 0.061609f
C840 VTAIL.n694 VSUBS 0.037623f
C841 VTAIL.n695 VSUBS 1.89079f
C842 VP.t1 VSUBS 3.57079f
C843 VP.n0 VSUBS 1.34392f
C844 VP.n1 VSUBS 0.025992f
C845 VP.n2 VSUBS 0.02224f
C846 VP.n3 VSUBS 0.025992f
C847 VP.t7 VSUBS 3.57079f
C848 VP.n4 VSUBS 1.24032f
C849 VP.n5 VSUBS 0.025992f
C850 VP.n6 VSUBS 0.021012f
C851 VP.n7 VSUBS 0.025992f
C852 VP.t0 VSUBS 3.57079f
C853 VP.n8 VSUBS 1.24032f
C854 VP.n9 VSUBS 0.025992f
C855 VP.n10 VSUBS 0.02224f
C856 VP.n11 VSUBS 0.025992f
C857 VP.t5 VSUBS 3.57079f
C858 VP.n12 VSUBS 1.34392f
C859 VP.t2 VSUBS 3.57079f
C860 VP.n13 VSUBS 1.34392f
C861 VP.n14 VSUBS 0.025992f
C862 VP.n15 VSUBS 0.02224f
C863 VP.n16 VSUBS 0.025992f
C864 VP.t3 VSUBS 3.57079f
C865 VP.n17 VSUBS 1.24032f
C866 VP.n18 VSUBS 0.025992f
C867 VP.n19 VSUBS 0.021012f
C868 VP.n20 VSUBS 0.025992f
C869 VP.t4 VSUBS 3.57079f
C870 VP.n21 VSUBS 1.32755f
C871 VP.t6 VSUBS 3.88837f
C872 VP.n22 VSUBS 1.27146f
C873 VP.n23 VSUBS 0.302278f
C874 VP.n24 VSUBS 0.03792f
C875 VP.n25 VSUBS 0.048443f
C876 VP.n26 VSUBS 0.051659f
C877 VP.n27 VSUBS 0.025992f
C878 VP.n28 VSUBS 0.025992f
C879 VP.n29 VSUBS 0.025992f
C880 VP.n30 VSUBS 0.051659f
C881 VP.n31 VSUBS 0.048443f
C882 VP.n32 VSUBS 0.03792f
C883 VP.n33 VSUBS 0.025992f
C884 VP.n34 VSUBS 0.025992f
C885 VP.n35 VSUBS 0.03505f
C886 VP.n36 VSUBS 0.048443f
C887 VP.n37 VSUBS 0.052522f
C888 VP.n38 VSUBS 0.025992f
C889 VP.n39 VSUBS 0.025992f
C890 VP.n40 VSUBS 0.025992f
C891 VP.n41 VSUBS 0.049569f
C892 VP.n42 VSUBS 0.048443f
C893 VP.n43 VSUBS 0.04079f
C894 VP.n44 VSUBS 0.041951f
C895 VP.n45 VSUBS 1.75752f
C896 VP.n46 VSUBS 1.77402f
C897 VP.n47 VSUBS 0.041951f
C898 VP.n48 VSUBS 0.04079f
C899 VP.n49 VSUBS 0.048443f
C900 VP.n50 VSUBS 0.049569f
C901 VP.n51 VSUBS 0.025992f
C902 VP.n52 VSUBS 0.025992f
C903 VP.n53 VSUBS 0.025992f
C904 VP.n54 VSUBS 0.052522f
C905 VP.n55 VSUBS 0.048443f
C906 VP.n56 VSUBS 0.03505f
C907 VP.n57 VSUBS 0.025992f
C908 VP.n58 VSUBS 0.025992f
C909 VP.n59 VSUBS 0.03792f
C910 VP.n60 VSUBS 0.048443f
C911 VP.n61 VSUBS 0.051659f
C912 VP.n62 VSUBS 0.025992f
C913 VP.n63 VSUBS 0.025992f
C914 VP.n64 VSUBS 0.025992f
C915 VP.n65 VSUBS 0.051659f
C916 VP.n66 VSUBS 0.048443f
C917 VP.n67 VSUBS 0.03792f
C918 VP.n68 VSUBS 0.025992f
C919 VP.n69 VSUBS 0.025992f
C920 VP.n70 VSUBS 0.03505f
C921 VP.n71 VSUBS 0.048443f
C922 VP.n72 VSUBS 0.052522f
C923 VP.n73 VSUBS 0.025992f
C924 VP.n74 VSUBS 0.025992f
C925 VP.n75 VSUBS 0.025992f
C926 VP.n76 VSUBS 0.049569f
C927 VP.n77 VSUBS 0.048443f
C928 VP.n78 VSUBS 0.04079f
C929 VP.n79 VSUBS 0.041951f
C930 VP.n80 VSUBS 0.060065f
C931 B.n0 VSUBS 0.006545f
C932 B.n1 VSUBS 0.006545f
C933 B.n2 VSUBS 0.00968f
C934 B.n3 VSUBS 0.007418f
C935 B.n4 VSUBS 0.007418f
C936 B.n5 VSUBS 0.007418f
C937 B.n6 VSUBS 0.007418f
C938 B.n7 VSUBS 0.007418f
C939 B.n8 VSUBS 0.007418f
C940 B.n9 VSUBS 0.007418f
C941 B.n10 VSUBS 0.007418f
C942 B.n11 VSUBS 0.007418f
C943 B.n12 VSUBS 0.007418f
C944 B.n13 VSUBS 0.007418f
C945 B.n14 VSUBS 0.007418f
C946 B.n15 VSUBS 0.007418f
C947 B.n16 VSUBS 0.007418f
C948 B.n17 VSUBS 0.007418f
C949 B.n18 VSUBS 0.007418f
C950 B.n19 VSUBS 0.007418f
C951 B.n20 VSUBS 0.007418f
C952 B.n21 VSUBS 0.007418f
C953 B.n22 VSUBS 0.007418f
C954 B.n23 VSUBS 0.007418f
C955 B.n24 VSUBS 0.007418f
C956 B.n25 VSUBS 0.007418f
C957 B.n26 VSUBS 0.007418f
C958 B.n27 VSUBS 0.007418f
C959 B.n28 VSUBS 0.007418f
C960 B.n29 VSUBS 0.007418f
C961 B.n30 VSUBS 0.007418f
C962 B.n31 VSUBS 0.007418f
C963 B.n32 VSUBS 0.018211f
C964 B.n33 VSUBS 0.007418f
C965 B.n34 VSUBS 0.007418f
C966 B.n35 VSUBS 0.007418f
C967 B.n36 VSUBS 0.007418f
C968 B.n37 VSUBS 0.007418f
C969 B.n38 VSUBS 0.007418f
C970 B.n39 VSUBS 0.007418f
C971 B.n40 VSUBS 0.007418f
C972 B.n41 VSUBS 0.007418f
C973 B.n42 VSUBS 0.007418f
C974 B.n43 VSUBS 0.007418f
C975 B.n44 VSUBS 0.007418f
C976 B.n45 VSUBS 0.007418f
C977 B.n46 VSUBS 0.007418f
C978 B.n47 VSUBS 0.007418f
C979 B.n48 VSUBS 0.007418f
C980 B.n49 VSUBS 0.007418f
C981 B.n50 VSUBS 0.007418f
C982 B.n51 VSUBS 0.007418f
C983 B.n52 VSUBS 0.007418f
C984 B.n53 VSUBS 0.007418f
C985 B.n54 VSUBS 0.007418f
C986 B.n55 VSUBS 0.007418f
C987 B.n56 VSUBS 0.007418f
C988 B.n57 VSUBS 0.007418f
C989 B.t1 VSUBS 0.30906f
C990 B.t2 VSUBS 0.350936f
C991 B.t0 VSUBS 2.41501f
C992 B.n58 VSUBS 0.554026f
C993 B.n59 VSUBS 0.318665f
C994 B.n60 VSUBS 0.017186f
C995 B.n61 VSUBS 0.007418f
C996 B.n62 VSUBS 0.007418f
C997 B.n63 VSUBS 0.007418f
C998 B.n64 VSUBS 0.007418f
C999 B.n65 VSUBS 0.007418f
C1000 B.t7 VSUBS 0.309063f
C1001 B.t8 VSUBS 0.350939f
C1002 B.t6 VSUBS 2.41501f
C1003 B.n66 VSUBS 0.554023f
C1004 B.n67 VSUBS 0.318661f
C1005 B.n68 VSUBS 0.007418f
C1006 B.n69 VSUBS 0.007418f
C1007 B.n70 VSUBS 0.007418f
C1008 B.n71 VSUBS 0.007418f
C1009 B.n72 VSUBS 0.007418f
C1010 B.n73 VSUBS 0.007418f
C1011 B.n74 VSUBS 0.007418f
C1012 B.n75 VSUBS 0.007418f
C1013 B.n76 VSUBS 0.007418f
C1014 B.n77 VSUBS 0.007418f
C1015 B.n78 VSUBS 0.007418f
C1016 B.n79 VSUBS 0.007418f
C1017 B.n80 VSUBS 0.007418f
C1018 B.n81 VSUBS 0.007418f
C1019 B.n82 VSUBS 0.007418f
C1020 B.n83 VSUBS 0.007418f
C1021 B.n84 VSUBS 0.007418f
C1022 B.n85 VSUBS 0.007418f
C1023 B.n86 VSUBS 0.007418f
C1024 B.n87 VSUBS 0.007418f
C1025 B.n88 VSUBS 0.007418f
C1026 B.n89 VSUBS 0.007418f
C1027 B.n90 VSUBS 0.007418f
C1028 B.n91 VSUBS 0.007418f
C1029 B.n92 VSUBS 0.007418f
C1030 B.n93 VSUBS 0.017787f
C1031 B.n94 VSUBS 0.007418f
C1032 B.n95 VSUBS 0.007418f
C1033 B.n96 VSUBS 0.007418f
C1034 B.n97 VSUBS 0.007418f
C1035 B.n98 VSUBS 0.007418f
C1036 B.n99 VSUBS 0.007418f
C1037 B.n100 VSUBS 0.007418f
C1038 B.n101 VSUBS 0.007418f
C1039 B.n102 VSUBS 0.007418f
C1040 B.n103 VSUBS 0.007418f
C1041 B.n104 VSUBS 0.007418f
C1042 B.n105 VSUBS 0.007418f
C1043 B.n106 VSUBS 0.007418f
C1044 B.n107 VSUBS 0.007418f
C1045 B.n108 VSUBS 0.007418f
C1046 B.n109 VSUBS 0.007418f
C1047 B.n110 VSUBS 0.007418f
C1048 B.n111 VSUBS 0.007418f
C1049 B.n112 VSUBS 0.007418f
C1050 B.n113 VSUBS 0.007418f
C1051 B.n114 VSUBS 0.007418f
C1052 B.n115 VSUBS 0.007418f
C1053 B.n116 VSUBS 0.007418f
C1054 B.n117 VSUBS 0.007418f
C1055 B.n118 VSUBS 0.007418f
C1056 B.n119 VSUBS 0.007418f
C1057 B.n120 VSUBS 0.007418f
C1058 B.n121 VSUBS 0.007418f
C1059 B.n122 VSUBS 0.007418f
C1060 B.n123 VSUBS 0.007418f
C1061 B.n124 VSUBS 0.007418f
C1062 B.n125 VSUBS 0.007418f
C1063 B.n126 VSUBS 0.007418f
C1064 B.n127 VSUBS 0.007418f
C1065 B.n128 VSUBS 0.007418f
C1066 B.n129 VSUBS 0.007418f
C1067 B.n130 VSUBS 0.007418f
C1068 B.n131 VSUBS 0.007418f
C1069 B.n132 VSUBS 0.007418f
C1070 B.n133 VSUBS 0.007418f
C1071 B.n134 VSUBS 0.007418f
C1072 B.n135 VSUBS 0.007418f
C1073 B.n136 VSUBS 0.007418f
C1074 B.n137 VSUBS 0.007418f
C1075 B.n138 VSUBS 0.007418f
C1076 B.n139 VSUBS 0.007418f
C1077 B.n140 VSUBS 0.007418f
C1078 B.n141 VSUBS 0.007418f
C1079 B.n142 VSUBS 0.007418f
C1080 B.n143 VSUBS 0.007418f
C1081 B.n144 VSUBS 0.007418f
C1082 B.n145 VSUBS 0.007418f
C1083 B.n146 VSUBS 0.007418f
C1084 B.n147 VSUBS 0.007418f
C1085 B.n148 VSUBS 0.007418f
C1086 B.n149 VSUBS 0.007418f
C1087 B.n150 VSUBS 0.007418f
C1088 B.n151 VSUBS 0.007418f
C1089 B.n152 VSUBS 0.007418f
C1090 B.n153 VSUBS 0.007418f
C1091 B.n154 VSUBS 0.017382f
C1092 B.n155 VSUBS 0.007418f
C1093 B.n156 VSUBS 0.007418f
C1094 B.n157 VSUBS 0.007418f
C1095 B.n158 VSUBS 0.007418f
C1096 B.n159 VSUBS 0.007418f
C1097 B.n160 VSUBS 0.007418f
C1098 B.n161 VSUBS 0.007418f
C1099 B.n162 VSUBS 0.007418f
C1100 B.n163 VSUBS 0.007418f
C1101 B.n164 VSUBS 0.007418f
C1102 B.n165 VSUBS 0.007418f
C1103 B.n166 VSUBS 0.007418f
C1104 B.n167 VSUBS 0.007418f
C1105 B.n168 VSUBS 0.007418f
C1106 B.n169 VSUBS 0.007418f
C1107 B.n170 VSUBS 0.007418f
C1108 B.n171 VSUBS 0.007418f
C1109 B.n172 VSUBS 0.007418f
C1110 B.n173 VSUBS 0.007418f
C1111 B.n174 VSUBS 0.007418f
C1112 B.n175 VSUBS 0.007418f
C1113 B.n176 VSUBS 0.007418f
C1114 B.n177 VSUBS 0.007418f
C1115 B.n178 VSUBS 0.007418f
C1116 B.n179 VSUBS 0.007418f
C1117 B.t11 VSUBS 0.309063f
C1118 B.t10 VSUBS 0.350939f
C1119 B.t9 VSUBS 2.41501f
C1120 B.n180 VSUBS 0.554023f
C1121 B.n181 VSUBS 0.318661f
C1122 B.n182 VSUBS 0.017186f
C1123 B.n183 VSUBS 0.007418f
C1124 B.n184 VSUBS 0.007418f
C1125 B.n185 VSUBS 0.007418f
C1126 B.n186 VSUBS 0.007418f
C1127 B.n187 VSUBS 0.007418f
C1128 B.t5 VSUBS 0.30906f
C1129 B.t4 VSUBS 0.350936f
C1130 B.t3 VSUBS 2.41501f
C1131 B.n188 VSUBS 0.554026f
C1132 B.n189 VSUBS 0.318665f
C1133 B.n190 VSUBS 0.007418f
C1134 B.n191 VSUBS 0.007418f
C1135 B.n192 VSUBS 0.007418f
C1136 B.n193 VSUBS 0.007418f
C1137 B.n194 VSUBS 0.007418f
C1138 B.n195 VSUBS 0.007418f
C1139 B.n196 VSUBS 0.007418f
C1140 B.n197 VSUBS 0.007418f
C1141 B.n198 VSUBS 0.007418f
C1142 B.n199 VSUBS 0.007418f
C1143 B.n200 VSUBS 0.007418f
C1144 B.n201 VSUBS 0.007418f
C1145 B.n202 VSUBS 0.007418f
C1146 B.n203 VSUBS 0.007418f
C1147 B.n204 VSUBS 0.007418f
C1148 B.n205 VSUBS 0.007418f
C1149 B.n206 VSUBS 0.007418f
C1150 B.n207 VSUBS 0.007418f
C1151 B.n208 VSUBS 0.007418f
C1152 B.n209 VSUBS 0.007418f
C1153 B.n210 VSUBS 0.007418f
C1154 B.n211 VSUBS 0.007418f
C1155 B.n212 VSUBS 0.007418f
C1156 B.n213 VSUBS 0.007418f
C1157 B.n214 VSUBS 0.007418f
C1158 B.n215 VSUBS 0.017787f
C1159 B.n216 VSUBS 0.007418f
C1160 B.n217 VSUBS 0.007418f
C1161 B.n218 VSUBS 0.007418f
C1162 B.n219 VSUBS 0.007418f
C1163 B.n220 VSUBS 0.007418f
C1164 B.n221 VSUBS 0.007418f
C1165 B.n222 VSUBS 0.007418f
C1166 B.n223 VSUBS 0.007418f
C1167 B.n224 VSUBS 0.007418f
C1168 B.n225 VSUBS 0.007418f
C1169 B.n226 VSUBS 0.007418f
C1170 B.n227 VSUBS 0.007418f
C1171 B.n228 VSUBS 0.007418f
C1172 B.n229 VSUBS 0.007418f
C1173 B.n230 VSUBS 0.007418f
C1174 B.n231 VSUBS 0.007418f
C1175 B.n232 VSUBS 0.007418f
C1176 B.n233 VSUBS 0.007418f
C1177 B.n234 VSUBS 0.007418f
C1178 B.n235 VSUBS 0.007418f
C1179 B.n236 VSUBS 0.007418f
C1180 B.n237 VSUBS 0.007418f
C1181 B.n238 VSUBS 0.007418f
C1182 B.n239 VSUBS 0.007418f
C1183 B.n240 VSUBS 0.007418f
C1184 B.n241 VSUBS 0.007418f
C1185 B.n242 VSUBS 0.007418f
C1186 B.n243 VSUBS 0.007418f
C1187 B.n244 VSUBS 0.007418f
C1188 B.n245 VSUBS 0.007418f
C1189 B.n246 VSUBS 0.007418f
C1190 B.n247 VSUBS 0.007418f
C1191 B.n248 VSUBS 0.007418f
C1192 B.n249 VSUBS 0.007418f
C1193 B.n250 VSUBS 0.007418f
C1194 B.n251 VSUBS 0.007418f
C1195 B.n252 VSUBS 0.007418f
C1196 B.n253 VSUBS 0.007418f
C1197 B.n254 VSUBS 0.007418f
C1198 B.n255 VSUBS 0.007418f
C1199 B.n256 VSUBS 0.007418f
C1200 B.n257 VSUBS 0.007418f
C1201 B.n258 VSUBS 0.007418f
C1202 B.n259 VSUBS 0.007418f
C1203 B.n260 VSUBS 0.007418f
C1204 B.n261 VSUBS 0.007418f
C1205 B.n262 VSUBS 0.007418f
C1206 B.n263 VSUBS 0.007418f
C1207 B.n264 VSUBS 0.007418f
C1208 B.n265 VSUBS 0.007418f
C1209 B.n266 VSUBS 0.007418f
C1210 B.n267 VSUBS 0.007418f
C1211 B.n268 VSUBS 0.007418f
C1212 B.n269 VSUBS 0.007418f
C1213 B.n270 VSUBS 0.007418f
C1214 B.n271 VSUBS 0.007418f
C1215 B.n272 VSUBS 0.007418f
C1216 B.n273 VSUBS 0.007418f
C1217 B.n274 VSUBS 0.007418f
C1218 B.n275 VSUBS 0.007418f
C1219 B.n276 VSUBS 0.007418f
C1220 B.n277 VSUBS 0.007418f
C1221 B.n278 VSUBS 0.007418f
C1222 B.n279 VSUBS 0.007418f
C1223 B.n280 VSUBS 0.007418f
C1224 B.n281 VSUBS 0.007418f
C1225 B.n282 VSUBS 0.007418f
C1226 B.n283 VSUBS 0.007418f
C1227 B.n284 VSUBS 0.007418f
C1228 B.n285 VSUBS 0.007418f
C1229 B.n286 VSUBS 0.007418f
C1230 B.n287 VSUBS 0.007418f
C1231 B.n288 VSUBS 0.007418f
C1232 B.n289 VSUBS 0.007418f
C1233 B.n290 VSUBS 0.007418f
C1234 B.n291 VSUBS 0.007418f
C1235 B.n292 VSUBS 0.007418f
C1236 B.n293 VSUBS 0.007418f
C1237 B.n294 VSUBS 0.007418f
C1238 B.n295 VSUBS 0.007418f
C1239 B.n296 VSUBS 0.007418f
C1240 B.n297 VSUBS 0.007418f
C1241 B.n298 VSUBS 0.007418f
C1242 B.n299 VSUBS 0.007418f
C1243 B.n300 VSUBS 0.007418f
C1244 B.n301 VSUBS 0.007418f
C1245 B.n302 VSUBS 0.007418f
C1246 B.n303 VSUBS 0.007418f
C1247 B.n304 VSUBS 0.007418f
C1248 B.n305 VSUBS 0.007418f
C1249 B.n306 VSUBS 0.007418f
C1250 B.n307 VSUBS 0.007418f
C1251 B.n308 VSUBS 0.007418f
C1252 B.n309 VSUBS 0.007418f
C1253 B.n310 VSUBS 0.007418f
C1254 B.n311 VSUBS 0.007418f
C1255 B.n312 VSUBS 0.007418f
C1256 B.n313 VSUBS 0.007418f
C1257 B.n314 VSUBS 0.007418f
C1258 B.n315 VSUBS 0.007418f
C1259 B.n316 VSUBS 0.007418f
C1260 B.n317 VSUBS 0.007418f
C1261 B.n318 VSUBS 0.007418f
C1262 B.n319 VSUBS 0.007418f
C1263 B.n320 VSUBS 0.007418f
C1264 B.n321 VSUBS 0.007418f
C1265 B.n322 VSUBS 0.007418f
C1266 B.n323 VSUBS 0.007418f
C1267 B.n324 VSUBS 0.007418f
C1268 B.n325 VSUBS 0.007418f
C1269 B.n326 VSUBS 0.007418f
C1270 B.n327 VSUBS 0.007418f
C1271 B.n328 VSUBS 0.007418f
C1272 B.n329 VSUBS 0.007418f
C1273 B.n330 VSUBS 0.007418f
C1274 B.n331 VSUBS 0.007418f
C1275 B.n332 VSUBS 0.017787f
C1276 B.n333 VSUBS 0.018211f
C1277 B.n334 VSUBS 0.018211f
C1278 B.n335 VSUBS 0.007418f
C1279 B.n336 VSUBS 0.007418f
C1280 B.n337 VSUBS 0.007418f
C1281 B.n338 VSUBS 0.007418f
C1282 B.n339 VSUBS 0.007418f
C1283 B.n340 VSUBS 0.007418f
C1284 B.n341 VSUBS 0.007418f
C1285 B.n342 VSUBS 0.007418f
C1286 B.n343 VSUBS 0.007418f
C1287 B.n344 VSUBS 0.007418f
C1288 B.n345 VSUBS 0.007418f
C1289 B.n346 VSUBS 0.007418f
C1290 B.n347 VSUBS 0.007418f
C1291 B.n348 VSUBS 0.007418f
C1292 B.n349 VSUBS 0.007418f
C1293 B.n350 VSUBS 0.007418f
C1294 B.n351 VSUBS 0.007418f
C1295 B.n352 VSUBS 0.007418f
C1296 B.n353 VSUBS 0.007418f
C1297 B.n354 VSUBS 0.007418f
C1298 B.n355 VSUBS 0.007418f
C1299 B.n356 VSUBS 0.007418f
C1300 B.n357 VSUBS 0.007418f
C1301 B.n358 VSUBS 0.007418f
C1302 B.n359 VSUBS 0.007418f
C1303 B.n360 VSUBS 0.007418f
C1304 B.n361 VSUBS 0.007418f
C1305 B.n362 VSUBS 0.007418f
C1306 B.n363 VSUBS 0.007418f
C1307 B.n364 VSUBS 0.007418f
C1308 B.n365 VSUBS 0.007418f
C1309 B.n366 VSUBS 0.007418f
C1310 B.n367 VSUBS 0.007418f
C1311 B.n368 VSUBS 0.007418f
C1312 B.n369 VSUBS 0.007418f
C1313 B.n370 VSUBS 0.007418f
C1314 B.n371 VSUBS 0.007418f
C1315 B.n372 VSUBS 0.007418f
C1316 B.n373 VSUBS 0.007418f
C1317 B.n374 VSUBS 0.007418f
C1318 B.n375 VSUBS 0.007418f
C1319 B.n376 VSUBS 0.007418f
C1320 B.n377 VSUBS 0.007418f
C1321 B.n378 VSUBS 0.007418f
C1322 B.n379 VSUBS 0.007418f
C1323 B.n380 VSUBS 0.007418f
C1324 B.n381 VSUBS 0.007418f
C1325 B.n382 VSUBS 0.007418f
C1326 B.n383 VSUBS 0.007418f
C1327 B.n384 VSUBS 0.007418f
C1328 B.n385 VSUBS 0.007418f
C1329 B.n386 VSUBS 0.007418f
C1330 B.n387 VSUBS 0.007418f
C1331 B.n388 VSUBS 0.007418f
C1332 B.n389 VSUBS 0.007418f
C1333 B.n390 VSUBS 0.007418f
C1334 B.n391 VSUBS 0.007418f
C1335 B.n392 VSUBS 0.007418f
C1336 B.n393 VSUBS 0.007418f
C1337 B.n394 VSUBS 0.007418f
C1338 B.n395 VSUBS 0.007418f
C1339 B.n396 VSUBS 0.007418f
C1340 B.n397 VSUBS 0.007418f
C1341 B.n398 VSUBS 0.007418f
C1342 B.n399 VSUBS 0.007418f
C1343 B.n400 VSUBS 0.007418f
C1344 B.n401 VSUBS 0.007418f
C1345 B.n402 VSUBS 0.007418f
C1346 B.n403 VSUBS 0.007418f
C1347 B.n404 VSUBS 0.007418f
C1348 B.n405 VSUBS 0.007418f
C1349 B.n406 VSUBS 0.007418f
C1350 B.n407 VSUBS 0.007418f
C1351 B.n408 VSUBS 0.007418f
C1352 B.n409 VSUBS 0.007418f
C1353 B.n410 VSUBS 0.005127f
C1354 B.n411 VSUBS 0.017186f
C1355 B.n412 VSUBS 0.006f
C1356 B.n413 VSUBS 0.007418f
C1357 B.n414 VSUBS 0.007418f
C1358 B.n415 VSUBS 0.007418f
C1359 B.n416 VSUBS 0.007418f
C1360 B.n417 VSUBS 0.007418f
C1361 B.n418 VSUBS 0.007418f
C1362 B.n419 VSUBS 0.007418f
C1363 B.n420 VSUBS 0.007418f
C1364 B.n421 VSUBS 0.007418f
C1365 B.n422 VSUBS 0.007418f
C1366 B.n423 VSUBS 0.007418f
C1367 B.n424 VSUBS 0.006f
C1368 B.n425 VSUBS 0.007418f
C1369 B.n426 VSUBS 0.007418f
C1370 B.n427 VSUBS 0.005127f
C1371 B.n428 VSUBS 0.007418f
C1372 B.n429 VSUBS 0.007418f
C1373 B.n430 VSUBS 0.007418f
C1374 B.n431 VSUBS 0.007418f
C1375 B.n432 VSUBS 0.007418f
C1376 B.n433 VSUBS 0.007418f
C1377 B.n434 VSUBS 0.007418f
C1378 B.n435 VSUBS 0.007418f
C1379 B.n436 VSUBS 0.007418f
C1380 B.n437 VSUBS 0.007418f
C1381 B.n438 VSUBS 0.007418f
C1382 B.n439 VSUBS 0.007418f
C1383 B.n440 VSUBS 0.007418f
C1384 B.n441 VSUBS 0.007418f
C1385 B.n442 VSUBS 0.007418f
C1386 B.n443 VSUBS 0.007418f
C1387 B.n444 VSUBS 0.007418f
C1388 B.n445 VSUBS 0.007418f
C1389 B.n446 VSUBS 0.007418f
C1390 B.n447 VSUBS 0.007418f
C1391 B.n448 VSUBS 0.007418f
C1392 B.n449 VSUBS 0.007418f
C1393 B.n450 VSUBS 0.007418f
C1394 B.n451 VSUBS 0.007418f
C1395 B.n452 VSUBS 0.007418f
C1396 B.n453 VSUBS 0.007418f
C1397 B.n454 VSUBS 0.007418f
C1398 B.n455 VSUBS 0.007418f
C1399 B.n456 VSUBS 0.007418f
C1400 B.n457 VSUBS 0.007418f
C1401 B.n458 VSUBS 0.007418f
C1402 B.n459 VSUBS 0.007418f
C1403 B.n460 VSUBS 0.007418f
C1404 B.n461 VSUBS 0.007418f
C1405 B.n462 VSUBS 0.007418f
C1406 B.n463 VSUBS 0.007418f
C1407 B.n464 VSUBS 0.007418f
C1408 B.n465 VSUBS 0.007418f
C1409 B.n466 VSUBS 0.007418f
C1410 B.n467 VSUBS 0.007418f
C1411 B.n468 VSUBS 0.007418f
C1412 B.n469 VSUBS 0.007418f
C1413 B.n470 VSUBS 0.007418f
C1414 B.n471 VSUBS 0.007418f
C1415 B.n472 VSUBS 0.007418f
C1416 B.n473 VSUBS 0.007418f
C1417 B.n474 VSUBS 0.007418f
C1418 B.n475 VSUBS 0.007418f
C1419 B.n476 VSUBS 0.007418f
C1420 B.n477 VSUBS 0.007418f
C1421 B.n478 VSUBS 0.007418f
C1422 B.n479 VSUBS 0.007418f
C1423 B.n480 VSUBS 0.007418f
C1424 B.n481 VSUBS 0.007418f
C1425 B.n482 VSUBS 0.007418f
C1426 B.n483 VSUBS 0.007418f
C1427 B.n484 VSUBS 0.007418f
C1428 B.n485 VSUBS 0.007418f
C1429 B.n486 VSUBS 0.007418f
C1430 B.n487 VSUBS 0.007418f
C1431 B.n488 VSUBS 0.007418f
C1432 B.n489 VSUBS 0.007418f
C1433 B.n490 VSUBS 0.007418f
C1434 B.n491 VSUBS 0.007418f
C1435 B.n492 VSUBS 0.007418f
C1436 B.n493 VSUBS 0.007418f
C1437 B.n494 VSUBS 0.007418f
C1438 B.n495 VSUBS 0.007418f
C1439 B.n496 VSUBS 0.007418f
C1440 B.n497 VSUBS 0.007418f
C1441 B.n498 VSUBS 0.007418f
C1442 B.n499 VSUBS 0.007418f
C1443 B.n500 VSUBS 0.007418f
C1444 B.n501 VSUBS 0.007418f
C1445 B.n502 VSUBS 0.007418f
C1446 B.n503 VSUBS 0.018211f
C1447 B.n504 VSUBS 0.017787f
C1448 B.n505 VSUBS 0.018616f
C1449 B.n506 VSUBS 0.007418f
C1450 B.n507 VSUBS 0.007418f
C1451 B.n508 VSUBS 0.007418f
C1452 B.n509 VSUBS 0.007418f
C1453 B.n510 VSUBS 0.007418f
C1454 B.n511 VSUBS 0.007418f
C1455 B.n512 VSUBS 0.007418f
C1456 B.n513 VSUBS 0.007418f
C1457 B.n514 VSUBS 0.007418f
C1458 B.n515 VSUBS 0.007418f
C1459 B.n516 VSUBS 0.007418f
C1460 B.n517 VSUBS 0.007418f
C1461 B.n518 VSUBS 0.007418f
C1462 B.n519 VSUBS 0.007418f
C1463 B.n520 VSUBS 0.007418f
C1464 B.n521 VSUBS 0.007418f
C1465 B.n522 VSUBS 0.007418f
C1466 B.n523 VSUBS 0.007418f
C1467 B.n524 VSUBS 0.007418f
C1468 B.n525 VSUBS 0.007418f
C1469 B.n526 VSUBS 0.007418f
C1470 B.n527 VSUBS 0.007418f
C1471 B.n528 VSUBS 0.007418f
C1472 B.n529 VSUBS 0.007418f
C1473 B.n530 VSUBS 0.007418f
C1474 B.n531 VSUBS 0.007418f
C1475 B.n532 VSUBS 0.007418f
C1476 B.n533 VSUBS 0.007418f
C1477 B.n534 VSUBS 0.007418f
C1478 B.n535 VSUBS 0.007418f
C1479 B.n536 VSUBS 0.007418f
C1480 B.n537 VSUBS 0.007418f
C1481 B.n538 VSUBS 0.007418f
C1482 B.n539 VSUBS 0.007418f
C1483 B.n540 VSUBS 0.007418f
C1484 B.n541 VSUBS 0.007418f
C1485 B.n542 VSUBS 0.007418f
C1486 B.n543 VSUBS 0.007418f
C1487 B.n544 VSUBS 0.007418f
C1488 B.n545 VSUBS 0.007418f
C1489 B.n546 VSUBS 0.007418f
C1490 B.n547 VSUBS 0.007418f
C1491 B.n548 VSUBS 0.007418f
C1492 B.n549 VSUBS 0.007418f
C1493 B.n550 VSUBS 0.007418f
C1494 B.n551 VSUBS 0.007418f
C1495 B.n552 VSUBS 0.007418f
C1496 B.n553 VSUBS 0.007418f
C1497 B.n554 VSUBS 0.007418f
C1498 B.n555 VSUBS 0.007418f
C1499 B.n556 VSUBS 0.007418f
C1500 B.n557 VSUBS 0.007418f
C1501 B.n558 VSUBS 0.007418f
C1502 B.n559 VSUBS 0.007418f
C1503 B.n560 VSUBS 0.007418f
C1504 B.n561 VSUBS 0.007418f
C1505 B.n562 VSUBS 0.007418f
C1506 B.n563 VSUBS 0.007418f
C1507 B.n564 VSUBS 0.007418f
C1508 B.n565 VSUBS 0.007418f
C1509 B.n566 VSUBS 0.007418f
C1510 B.n567 VSUBS 0.007418f
C1511 B.n568 VSUBS 0.007418f
C1512 B.n569 VSUBS 0.007418f
C1513 B.n570 VSUBS 0.007418f
C1514 B.n571 VSUBS 0.007418f
C1515 B.n572 VSUBS 0.007418f
C1516 B.n573 VSUBS 0.007418f
C1517 B.n574 VSUBS 0.007418f
C1518 B.n575 VSUBS 0.007418f
C1519 B.n576 VSUBS 0.007418f
C1520 B.n577 VSUBS 0.007418f
C1521 B.n578 VSUBS 0.007418f
C1522 B.n579 VSUBS 0.007418f
C1523 B.n580 VSUBS 0.007418f
C1524 B.n581 VSUBS 0.007418f
C1525 B.n582 VSUBS 0.007418f
C1526 B.n583 VSUBS 0.007418f
C1527 B.n584 VSUBS 0.007418f
C1528 B.n585 VSUBS 0.007418f
C1529 B.n586 VSUBS 0.007418f
C1530 B.n587 VSUBS 0.007418f
C1531 B.n588 VSUBS 0.007418f
C1532 B.n589 VSUBS 0.007418f
C1533 B.n590 VSUBS 0.007418f
C1534 B.n591 VSUBS 0.007418f
C1535 B.n592 VSUBS 0.007418f
C1536 B.n593 VSUBS 0.007418f
C1537 B.n594 VSUBS 0.007418f
C1538 B.n595 VSUBS 0.007418f
C1539 B.n596 VSUBS 0.007418f
C1540 B.n597 VSUBS 0.007418f
C1541 B.n598 VSUBS 0.007418f
C1542 B.n599 VSUBS 0.007418f
C1543 B.n600 VSUBS 0.007418f
C1544 B.n601 VSUBS 0.007418f
C1545 B.n602 VSUBS 0.007418f
C1546 B.n603 VSUBS 0.007418f
C1547 B.n604 VSUBS 0.007418f
C1548 B.n605 VSUBS 0.007418f
C1549 B.n606 VSUBS 0.007418f
C1550 B.n607 VSUBS 0.007418f
C1551 B.n608 VSUBS 0.007418f
C1552 B.n609 VSUBS 0.007418f
C1553 B.n610 VSUBS 0.007418f
C1554 B.n611 VSUBS 0.007418f
C1555 B.n612 VSUBS 0.007418f
C1556 B.n613 VSUBS 0.007418f
C1557 B.n614 VSUBS 0.007418f
C1558 B.n615 VSUBS 0.007418f
C1559 B.n616 VSUBS 0.007418f
C1560 B.n617 VSUBS 0.007418f
C1561 B.n618 VSUBS 0.007418f
C1562 B.n619 VSUBS 0.007418f
C1563 B.n620 VSUBS 0.007418f
C1564 B.n621 VSUBS 0.007418f
C1565 B.n622 VSUBS 0.007418f
C1566 B.n623 VSUBS 0.007418f
C1567 B.n624 VSUBS 0.007418f
C1568 B.n625 VSUBS 0.007418f
C1569 B.n626 VSUBS 0.007418f
C1570 B.n627 VSUBS 0.007418f
C1571 B.n628 VSUBS 0.007418f
C1572 B.n629 VSUBS 0.007418f
C1573 B.n630 VSUBS 0.007418f
C1574 B.n631 VSUBS 0.007418f
C1575 B.n632 VSUBS 0.007418f
C1576 B.n633 VSUBS 0.007418f
C1577 B.n634 VSUBS 0.007418f
C1578 B.n635 VSUBS 0.007418f
C1579 B.n636 VSUBS 0.007418f
C1580 B.n637 VSUBS 0.007418f
C1581 B.n638 VSUBS 0.007418f
C1582 B.n639 VSUBS 0.007418f
C1583 B.n640 VSUBS 0.007418f
C1584 B.n641 VSUBS 0.007418f
C1585 B.n642 VSUBS 0.007418f
C1586 B.n643 VSUBS 0.007418f
C1587 B.n644 VSUBS 0.007418f
C1588 B.n645 VSUBS 0.007418f
C1589 B.n646 VSUBS 0.007418f
C1590 B.n647 VSUBS 0.007418f
C1591 B.n648 VSUBS 0.007418f
C1592 B.n649 VSUBS 0.007418f
C1593 B.n650 VSUBS 0.007418f
C1594 B.n651 VSUBS 0.007418f
C1595 B.n652 VSUBS 0.007418f
C1596 B.n653 VSUBS 0.007418f
C1597 B.n654 VSUBS 0.007418f
C1598 B.n655 VSUBS 0.007418f
C1599 B.n656 VSUBS 0.007418f
C1600 B.n657 VSUBS 0.007418f
C1601 B.n658 VSUBS 0.007418f
C1602 B.n659 VSUBS 0.007418f
C1603 B.n660 VSUBS 0.007418f
C1604 B.n661 VSUBS 0.007418f
C1605 B.n662 VSUBS 0.007418f
C1606 B.n663 VSUBS 0.007418f
C1607 B.n664 VSUBS 0.007418f
C1608 B.n665 VSUBS 0.007418f
C1609 B.n666 VSUBS 0.007418f
C1610 B.n667 VSUBS 0.007418f
C1611 B.n668 VSUBS 0.007418f
C1612 B.n669 VSUBS 0.007418f
C1613 B.n670 VSUBS 0.007418f
C1614 B.n671 VSUBS 0.007418f
C1615 B.n672 VSUBS 0.007418f
C1616 B.n673 VSUBS 0.007418f
C1617 B.n674 VSUBS 0.007418f
C1618 B.n675 VSUBS 0.007418f
C1619 B.n676 VSUBS 0.007418f
C1620 B.n677 VSUBS 0.007418f
C1621 B.n678 VSUBS 0.007418f
C1622 B.n679 VSUBS 0.007418f
C1623 B.n680 VSUBS 0.007418f
C1624 B.n681 VSUBS 0.007418f
C1625 B.n682 VSUBS 0.007418f
C1626 B.n683 VSUBS 0.007418f
C1627 B.n684 VSUBS 0.007418f
C1628 B.n685 VSUBS 0.007418f
C1629 B.n686 VSUBS 0.017787f
C1630 B.n687 VSUBS 0.018211f
C1631 B.n688 VSUBS 0.018211f
C1632 B.n689 VSUBS 0.007418f
C1633 B.n690 VSUBS 0.007418f
C1634 B.n691 VSUBS 0.007418f
C1635 B.n692 VSUBS 0.007418f
C1636 B.n693 VSUBS 0.007418f
C1637 B.n694 VSUBS 0.007418f
C1638 B.n695 VSUBS 0.007418f
C1639 B.n696 VSUBS 0.007418f
C1640 B.n697 VSUBS 0.007418f
C1641 B.n698 VSUBS 0.007418f
C1642 B.n699 VSUBS 0.007418f
C1643 B.n700 VSUBS 0.007418f
C1644 B.n701 VSUBS 0.007418f
C1645 B.n702 VSUBS 0.007418f
C1646 B.n703 VSUBS 0.007418f
C1647 B.n704 VSUBS 0.007418f
C1648 B.n705 VSUBS 0.007418f
C1649 B.n706 VSUBS 0.007418f
C1650 B.n707 VSUBS 0.007418f
C1651 B.n708 VSUBS 0.007418f
C1652 B.n709 VSUBS 0.007418f
C1653 B.n710 VSUBS 0.007418f
C1654 B.n711 VSUBS 0.007418f
C1655 B.n712 VSUBS 0.007418f
C1656 B.n713 VSUBS 0.007418f
C1657 B.n714 VSUBS 0.007418f
C1658 B.n715 VSUBS 0.007418f
C1659 B.n716 VSUBS 0.007418f
C1660 B.n717 VSUBS 0.007418f
C1661 B.n718 VSUBS 0.007418f
C1662 B.n719 VSUBS 0.007418f
C1663 B.n720 VSUBS 0.007418f
C1664 B.n721 VSUBS 0.007418f
C1665 B.n722 VSUBS 0.007418f
C1666 B.n723 VSUBS 0.007418f
C1667 B.n724 VSUBS 0.007418f
C1668 B.n725 VSUBS 0.007418f
C1669 B.n726 VSUBS 0.007418f
C1670 B.n727 VSUBS 0.007418f
C1671 B.n728 VSUBS 0.007418f
C1672 B.n729 VSUBS 0.007418f
C1673 B.n730 VSUBS 0.007418f
C1674 B.n731 VSUBS 0.007418f
C1675 B.n732 VSUBS 0.007418f
C1676 B.n733 VSUBS 0.007418f
C1677 B.n734 VSUBS 0.007418f
C1678 B.n735 VSUBS 0.007418f
C1679 B.n736 VSUBS 0.007418f
C1680 B.n737 VSUBS 0.007418f
C1681 B.n738 VSUBS 0.007418f
C1682 B.n739 VSUBS 0.007418f
C1683 B.n740 VSUBS 0.007418f
C1684 B.n741 VSUBS 0.007418f
C1685 B.n742 VSUBS 0.007418f
C1686 B.n743 VSUBS 0.007418f
C1687 B.n744 VSUBS 0.007418f
C1688 B.n745 VSUBS 0.007418f
C1689 B.n746 VSUBS 0.007418f
C1690 B.n747 VSUBS 0.007418f
C1691 B.n748 VSUBS 0.007418f
C1692 B.n749 VSUBS 0.007418f
C1693 B.n750 VSUBS 0.007418f
C1694 B.n751 VSUBS 0.007418f
C1695 B.n752 VSUBS 0.007418f
C1696 B.n753 VSUBS 0.007418f
C1697 B.n754 VSUBS 0.007418f
C1698 B.n755 VSUBS 0.007418f
C1699 B.n756 VSUBS 0.007418f
C1700 B.n757 VSUBS 0.007418f
C1701 B.n758 VSUBS 0.007418f
C1702 B.n759 VSUBS 0.007418f
C1703 B.n760 VSUBS 0.007418f
C1704 B.n761 VSUBS 0.007418f
C1705 B.n762 VSUBS 0.007418f
C1706 B.n763 VSUBS 0.007418f
C1707 B.n764 VSUBS 0.005127f
C1708 B.n765 VSUBS 0.017186f
C1709 B.n766 VSUBS 0.006f
C1710 B.n767 VSUBS 0.007418f
C1711 B.n768 VSUBS 0.007418f
C1712 B.n769 VSUBS 0.007418f
C1713 B.n770 VSUBS 0.007418f
C1714 B.n771 VSUBS 0.007418f
C1715 B.n772 VSUBS 0.007418f
C1716 B.n773 VSUBS 0.007418f
C1717 B.n774 VSUBS 0.007418f
C1718 B.n775 VSUBS 0.007418f
C1719 B.n776 VSUBS 0.007418f
C1720 B.n777 VSUBS 0.007418f
C1721 B.n778 VSUBS 0.006f
C1722 B.n779 VSUBS 0.007418f
C1723 B.n780 VSUBS 0.007418f
C1724 B.n781 VSUBS 0.005127f
C1725 B.n782 VSUBS 0.007418f
C1726 B.n783 VSUBS 0.007418f
C1727 B.n784 VSUBS 0.007418f
C1728 B.n785 VSUBS 0.007418f
C1729 B.n786 VSUBS 0.007418f
C1730 B.n787 VSUBS 0.007418f
C1731 B.n788 VSUBS 0.007418f
C1732 B.n789 VSUBS 0.007418f
C1733 B.n790 VSUBS 0.007418f
C1734 B.n791 VSUBS 0.007418f
C1735 B.n792 VSUBS 0.007418f
C1736 B.n793 VSUBS 0.007418f
C1737 B.n794 VSUBS 0.007418f
C1738 B.n795 VSUBS 0.007418f
C1739 B.n796 VSUBS 0.007418f
C1740 B.n797 VSUBS 0.007418f
C1741 B.n798 VSUBS 0.007418f
C1742 B.n799 VSUBS 0.007418f
C1743 B.n800 VSUBS 0.007418f
C1744 B.n801 VSUBS 0.007418f
C1745 B.n802 VSUBS 0.007418f
C1746 B.n803 VSUBS 0.007418f
C1747 B.n804 VSUBS 0.007418f
C1748 B.n805 VSUBS 0.007418f
C1749 B.n806 VSUBS 0.007418f
C1750 B.n807 VSUBS 0.007418f
C1751 B.n808 VSUBS 0.007418f
C1752 B.n809 VSUBS 0.007418f
C1753 B.n810 VSUBS 0.007418f
C1754 B.n811 VSUBS 0.007418f
C1755 B.n812 VSUBS 0.007418f
C1756 B.n813 VSUBS 0.007418f
C1757 B.n814 VSUBS 0.007418f
C1758 B.n815 VSUBS 0.007418f
C1759 B.n816 VSUBS 0.007418f
C1760 B.n817 VSUBS 0.007418f
C1761 B.n818 VSUBS 0.007418f
C1762 B.n819 VSUBS 0.007418f
C1763 B.n820 VSUBS 0.007418f
C1764 B.n821 VSUBS 0.007418f
C1765 B.n822 VSUBS 0.007418f
C1766 B.n823 VSUBS 0.007418f
C1767 B.n824 VSUBS 0.007418f
C1768 B.n825 VSUBS 0.007418f
C1769 B.n826 VSUBS 0.007418f
C1770 B.n827 VSUBS 0.007418f
C1771 B.n828 VSUBS 0.007418f
C1772 B.n829 VSUBS 0.007418f
C1773 B.n830 VSUBS 0.007418f
C1774 B.n831 VSUBS 0.007418f
C1775 B.n832 VSUBS 0.007418f
C1776 B.n833 VSUBS 0.007418f
C1777 B.n834 VSUBS 0.007418f
C1778 B.n835 VSUBS 0.007418f
C1779 B.n836 VSUBS 0.007418f
C1780 B.n837 VSUBS 0.007418f
C1781 B.n838 VSUBS 0.007418f
C1782 B.n839 VSUBS 0.007418f
C1783 B.n840 VSUBS 0.007418f
C1784 B.n841 VSUBS 0.007418f
C1785 B.n842 VSUBS 0.007418f
C1786 B.n843 VSUBS 0.007418f
C1787 B.n844 VSUBS 0.007418f
C1788 B.n845 VSUBS 0.007418f
C1789 B.n846 VSUBS 0.007418f
C1790 B.n847 VSUBS 0.007418f
C1791 B.n848 VSUBS 0.007418f
C1792 B.n849 VSUBS 0.007418f
C1793 B.n850 VSUBS 0.007418f
C1794 B.n851 VSUBS 0.007418f
C1795 B.n852 VSUBS 0.007418f
C1796 B.n853 VSUBS 0.007418f
C1797 B.n854 VSUBS 0.007418f
C1798 B.n855 VSUBS 0.007418f
C1799 B.n856 VSUBS 0.007418f
C1800 B.n857 VSUBS 0.018211f
C1801 B.n858 VSUBS 0.017787f
C1802 B.n859 VSUBS 0.017787f
C1803 B.n860 VSUBS 0.007418f
C1804 B.n861 VSUBS 0.007418f
C1805 B.n862 VSUBS 0.007418f
C1806 B.n863 VSUBS 0.007418f
C1807 B.n864 VSUBS 0.007418f
C1808 B.n865 VSUBS 0.007418f
C1809 B.n866 VSUBS 0.007418f
C1810 B.n867 VSUBS 0.007418f
C1811 B.n868 VSUBS 0.007418f
C1812 B.n869 VSUBS 0.007418f
C1813 B.n870 VSUBS 0.007418f
C1814 B.n871 VSUBS 0.007418f
C1815 B.n872 VSUBS 0.007418f
C1816 B.n873 VSUBS 0.007418f
C1817 B.n874 VSUBS 0.007418f
C1818 B.n875 VSUBS 0.007418f
C1819 B.n876 VSUBS 0.007418f
C1820 B.n877 VSUBS 0.007418f
C1821 B.n878 VSUBS 0.007418f
C1822 B.n879 VSUBS 0.007418f
C1823 B.n880 VSUBS 0.007418f
C1824 B.n881 VSUBS 0.007418f
C1825 B.n882 VSUBS 0.007418f
C1826 B.n883 VSUBS 0.007418f
C1827 B.n884 VSUBS 0.007418f
C1828 B.n885 VSUBS 0.007418f
C1829 B.n886 VSUBS 0.007418f
C1830 B.n887 VSUBS 0.007418f
C1831 B.n888 VSUBS 0.007418f
C1832 B.n889 VSUBS 0.007418f
C1833 B.n890 VSUBS 0.007418f
C1834 B.n891 VSUBS 0.007418f
C1835 B.n892 VSUBS 0.007418f
C1836 B.n893 VSUBS 0.007418f
C1837 B.n894 VSUBS 0.007418f
C1838 B.n895 VSUBS 0.007418f
C1839 B.n896 VSUBS 0.007418f
C1840 B.n897 VSUBS 0.007418f
C1841 B.n898 VSUBS 0.007418f
C1842 B.n899 VSUBS 0.007418f
C1843 B.n900 VSUBS 0.007418f
C1844 B.n901 VSUBS 0.007418f
C1845 B.n902 VSUBS 0.007418f
C1846 B.n903 VSUBS 0.007418f
C1847 B.n904 VSUBS 0.007418f
C1848 B.n905 VSUBS 0.007418f
C1849 B.n906 VSUBS 0.007418f
C1850 B.n907 VSUBS 0.007418f
C1851 B.n908 VSUBS 0.007418f
C1852 B.n909 VSUBS 0.007418f
C1853 B.n910 VSUBS 0.007418f
C1854 B.n911 VSUBS 0.007418f
C1855 B.n912 VSUBS 0.007418f
C1856 B.n913 VSUBS 0.007418f
C1857 B.n914 VSUBS 0.007418f
C1858 B.n915 VSUBS 0.007418f
C1859 B.n916 VSUBS 0.007418f
C1860 B.n917 VSUBS 0.007418f
C1861 B.n918 VSUBS 0.007418f
C1862 B.n919 VSUBS 0.007418f
C1863 B.n920 VSUBS 0.007418f
C1864 B.n921 VSUBS 0.007418f
C1865 B.n922 VSUBS 0.007418f
C1866 B.n923 VSUBS 0.007418f
C1867 B.n924 VSUBS 0.007418f
C1868 B.n925 VSUBS 0.007418f
C1869 B.n926 VSUBS 0.007418f
C1870 B.n927 VSUBS 0.007418f
C1871 B.n928 VSUBS 0.007418f
C1872 B.n929 VSUBS 0.007418f
C1873 B.n930 VSUBS 0.007418f
C1874 B.n931 VSUBS 0.007418f
C1875 B.n932 VSUBS 0.007418f
C1876 B.n933 VSUBS 0.007418f
C1877 B.n934 VSUBS 0.007418f
C1878 B.n935 VSUBS 0.007418f
C1879 B.n936 VSUBS 0.007418f
C1880 B.n937 VSUBS 0.007418f
C1881 B.n938 VSUBS 0.007418f
C1882 B.n939 VSUBS 0.007418f
C1883 B.n940 VSUBS 0.007418f
C1884 B.n941 VSUBS 0.007418f
C1885 B.n942 VSUBS 0.007418f
C1886 B.n943 VSUBS 0.007418f
C1887 B.n944 VSUBS 0.007418f
C1888 B.n945 VSUBS 0.007418f
C1889 B.n946 VSUBS 0.007418f
C1890 B.n947 VSUBS 0.00968f
C1891 B.n948 VSUBS 0.010311f
C1892 B.n949 VSUBS 0.020505f
.ends

