* NGSPICE file created from diff_pair_sample_1093.ext - technology: sky130A

.subckt diff_pair_sample_1093 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=5.1129 pd=27 as=2.16315 ps=13.44 w=13.11 l=0.82
X1 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=5.1129 pd=27 as=0 ps=0 w=13.11 l=0.82
X2 VDD2.t1 VN.t1 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=2.16315 pd=13.44 as=2.16315 ps=13.44 w=13.11 l=0.82
X3 VDD1.t7 VP.t0 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.16315 pd=13.44 as=5.1129 ps=27 w=13.11 l=0.82
X4 VDD2.t6 VN.t2 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=2.16315 pd=13.44 as=2.16315 ps=13.44 w=13.11 l=0.82
X5 VTAIL.t12 VN.t3 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=2.16315 pd=13.44 as=2.16315 ps=13.44 w=13.11 l=0.82
X6 VTAIL.t6 VP.t1 VDD1.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.16315 pd=13.44 as=2.16315 ps=13.44 w=13.11 l=0.82
X7 VTAIL.t11 VN.t4 VDD2.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=2.16315 pd=13.44 as=2.16315 ps=13.44 w=13.11 l=0.82
X8 VDD2.t4 VN.t5 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=2.16315 pd=13.44 as=5.1129 ps=27 w=13.11 l=0.82
X9 VDD1.t5 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.16315 pd=13.44 as=2.16315 ps=13.44 w=13.11 l=0.82
X10 VDD1.t4 VP.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.16315 pd=13.44 as=5.1129 ps=27 w=13.11 l=0.82
X11 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=5.1129 pd=27 as=0 ps=0 w=13.11 l=0.82
X12 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=5.1129 pd=27 as=0 ps=0 w=13.11 l=0.82
X13 VTAIL.t5 VP.t4 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=5.1129 pd=27 as=2.16315 ps=13.44 w=13.11 l=0.82
X14 VDD2.t2 VN.t6 VTAIL.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=2.16315 pd=13.44 as=5.1129 ps=27 w=13.11 l=0.82
X15 VDD1.t2 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.16315 pd=13.44 as=2.16315 ps=13.44 w=13.11 l=0.82
X16 VTAIL.t2 VP.t6 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=5.1129 pd=27 as=2.16315 ps=13.44 w=13.11 l=0.82
X17 VTAIL.t8 VN.t7 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=5.1129 pd=27 as=2.16315 ps=13.44 w=13.11 l=0.82
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.1129 pd=27 as=0 ps=0 w=13.11 l=0.82
X19 VTAIL.t0 VP.t7 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.16315 pd=13.44 as=2.16315 ps=13.44 w=13.11 l=0.82
R0 VN.n3 VN.t0 452.738
R1 VN.n16 VN.t6 452.738
R2 VN.n11 VN.t5 433.507
R3 VN.n24 VN.t7 433.507
R4 VN.n4 VN.t1 385.307
R5 VN.n1 VN.t3 385.307
R6 VN.n17 VN.t4 385.307
R7 VN.n14 VN.t2 385.307
R8 VN.n12 VN.n11 161.3
R9 VN.n25 VN.n24 161.3
R10 VN.n23 VN.n13 161.3
R11 VN.n22 VN.n21 161.3
R12 VN.n20 VN.n19 161.3
R13 VN.n18 VN.n15 161.3
R14 VN.n10 VN.n0 161.3
R15 VN.n9 VN.n8 161.3
R16 VN.n7 VN.n6 161.3
R17 VN.n5 VN.n2 161.3
R18 VN.n6 VN.n5 56.5193
R19 VN.n19 VN.n18 56.5193
R20 VN.n10 VN.n9 50.2061
R21 VN.n23 VN.n22 50.2061
R22 VN VN.n25 43.7524
R23 VN.n16 VN.n15 43.2015
R24 VN.n3 VN.n2 43.2015
R25 VN.n4 VN.n3 38.5669
R26 VN.n17 VN.n16 38.5669
R27 VN.n5 VN.n4 15.9041
R28 VN.n6 VN.n1 15.9041
R29 VN.n18 VN.n17 15.9041
R30 VN.n19 VN.n14 15.9041
R31 VN.n11 VN.n10 9.49444
R32 VN.n24 VN.n23 9.49444
R33 VN.n9 VN.n1 8.56395
R34 VN.n22 VN.n14 8.56395
R35 VN.n25 VN.n13 0.189894
R36 VN.n21 VN.n13 0.189894
R37 VN.n21 VN.n20 0.189894
R38 VN.n20 VN.n15 0.189894
R39 VN.n7 VN.n2 0.189894
R40 VN.n8 VN.n7 0.189894
R41 VN.n8 VN.n0 0.189894
R42 VN.n12 VN.n0 0.189894
R43 VN VN.n12 0.0516364
R44 VDD2.n2 VDD2.n1 60.3201
R45 VDD2.n2 VDD2.n0 60.3201
R46 VDD2 VDD2.n5 60.3172
R47 VDD2.n4 VDD2.n3 59.8799
R48 VDD2.n4 VDD2.n2 39.4782
R49 VDD2.n5 VDD2.t0 1.5108
R50 VDD2.n5 VDD2.t2 1.5108
R51 VDD2.n3 VDD2.t3 1.5108
R52 VDD2.n3 VDD2.t6 1.5108
R53 VDD2.n1 VDD2.t5 1.5108
R54 VDD2.n1 VDD2.t4 1.5108
R55 VDD2.n0 VDD2.t7 1.5108
R56 VDD2.n0 VDD2.t1 1.5108
R57 VDD2 VDD2.n4 0.554379
R58 VTAIL.n11 VTAIL.t5 44.7114
R59 VTAIL.n10 VTAIL.t9 44.7114
R60 VTAIL.n7 VTAIL.t8 44.7114
R61 VTAIL.n15 VTAIL.t10 44.7111
R62 VTAIL.n2 VTAIL.t15 44.7111
R63 VTAIL.n3 VTAIL.t7 44.7111
R64 VTAIL.n6 VTAIL.t2 44.7111
R65 VTAIL.n14 VTAIL.t4 44.7111
R66 VTAIL.n13 VTAIL.n12 43.2011
R67 VTAIL.n9 VTAIL.n8 43.2011
R68 VTAIL.n1 VTAIL.n0 43.201
R69 VTAIL.n5 VTAIL.n4 43.201
R70 VTAIL.n15 VTAIL.n14 24.66
R71 VTAIL.n7 VTAIL.n6 24.66
R72 VTAIL.n0 VTAIL.t14 1.5108
R73 VTAIL.n0 VTAIL.t12 1.5108
R74 VTAIL.n4 VTAIL.t3 1.5108
R75 VTAIL.n4 VTAIL.t6 1.5108
R76 VTAIL.n12 VTAIL.t1 1.5108
R77 VTAIL.n12 VTAIL.t0 1.5108
R78 VTAIL.n8 VTAIL.t13 1.5108
R79 VTAIL.n8 VTAIL.t11 1.5108
R80 VTAIL.n9 VTAIL.n7 0.991879
R81 VTAIL.n10 VTAIL.n9 0.991879
R82 VTAIL.n13 VTAIL.n11 0.991879
R83 VTAIL.n14 VTAIL.n13 0.991879
R84 VTAIL.n6 VTAIL.n5 0.991879
R85 VTAIL.n5 VTAIL.n3 0.991879
R86 VTAIL.n2 VTAIL.n1 0.991879
R87 VTAIL VTAIL.n15 0.93369
R88 VTAIL.n11 VTAIL.n10 0.470328
R89 VTAIL.n3 VTAIL.n2 0.470328
R90 VTAIL VTAIL.n1 0.0586897
R91 B.n400 B.t15 586.967
R92 B.n397 B.t19 586.967
R93 B.n102 B.t8 586.967
R94 B.n99 B.t12 586.967
R95 B.n709 B.n708 585
R96 B.n710 B.n709 585
R97 B.n299 B.n98 585
R98 B.n298 B.n297 585
R99 B.n296 B.n295 585
R100 B.n294 B.n293 585
R101 B.n292 B.n291 585
R102 B.n290 B.n289 585
R103 B.n288 B.n287 585
R104 B.n286 B.n285 585
R105 B.n284 B.n283 585
R106 B.n282 B.n281 585
R107 B.n280 B.n279 585
R108 B.n278 B.n277 585
R109 B.n276 B.n275 585
R110 B.n274 B.n273 585
R111 B.n272 B.n271 585
R112 B.n270 B.n269 585
R113 B.n268 B.n267 585
R114 B.n266 B.n265 585
R115 B.n264 B.n263 585
R116 B.n262 B.n261 585
R117 B.n260 B.n259 585
R118 B.n258 B.n257 585
R119 B.n256 B.n255 585
R120 B.n254 B.n253 585
R121 B.n252 B.n251 585
R122 B.n250 B.n249 585
R123 B.n248 B.n247 585
R124 B.n246 B.n245 585
R125 B.n244 B.n243 585
R126 B.n242 B.n241 585
R127 B.n240 B.n239 585
R128 B.n238 B.n237 585
R129 B.n236 B.n235 585
R130 B.n234 B.n233 585
R131 B.n232 B.n231 585
R132 B.n230 B.n229 585
R133 B.n228 B.n227 585
R134 B.n226 B.n225 585
R135 B.n224 B.n223 585
R136 B.n222 B.n221 585
R137 B.n220 B.n219 585
R138 B.n218 B.n217 585
R139 B.n216 B.n215 585
R140 B.n214 B.n213 585
R141 B.n212 B.n211 585
R142 B.n210 B.n209 585
R143 B.n208 B.n207 585
R144 B.n206 B.n205 585
R145 B.n204 B.n203 585
R146 B.n202 B.n201 585
R147 B.n200 B.n199 585
R148 B.n198 B.n197 585
R149 B.n196 B.n195 585
R150 B.n193 B.n192 585
R151 B.n191 B.n190 585
R152 B.n189 B.n188 585
R153 B.n187 B.n186 585
R154 B.n185 B.n184 585
R155 B.n183 B.n182 585
R156 B.n181 B.n180 585
R157 B.n179 B.n178 585
R158 B.n177 B.n176 585
R159 B.n175 B.n174 585
R160 B.n173 B.n172 585
R161 B.n171 B.n170 585
R162 B.n169 B.n168 585
R163 B.n167 B.n166 585
R164 B.n165 B.n164 585
R165 B.n163 B.n162 585
R166 B.n161 B.n160 585
R167 B.n159 B.n158 585
R168 B.n157 B.n156 585
R169 B.n155 B.n154 585
R170 B.n153 B.n152 585
R171 B.n151 B.n150 585
R172 B.n149 B.n148 585
R173 B.n147 B.n146 585
R174 B.n145 B.n144 585
R175 B.n143 B.n142 585
R176 B.n141 B.n140 585
R177 B.n139 B.n138 585
R178 B.n137 B.n136 585
R179 B.n135 B.n134 585
R180 B.n133 B.n132 585
R181 B.n131 B.n130 585
R182 B.n129 B.n128 585
R183 B.n127 B.n126 585
R184 B.n125 B.n124 585
R185 B.n123 B.n122 585
R186 B.n121 B.n120 585
R187 B.n119 B.n118 585
R188 B.n117 B.n116 585
R189 B.n115 B.n114 585
R190 B.n113 B.n112 585
R191 B.n111 B.n110 585
R192 B.n109 B.n108 585
R193 B.n107 B.n106 585
R194 B.n105 B.n104 585
R195 B.n707 B.n48 585
R196 B.n711 B.n48 585
R197 B.n706 B.n47 585
R198 B.n712 B.n47 585
R199 B.n705 B.n704 585
R200 B.n704 B.n43 585
R201 B.n703 B.n42 585
R202 B.n718 B.n42 585
R203 B.n702 B.n41 585
R204 B.n719 B.n41 585
R205 B.n701 B.n40 585
R206 B.n720 B.n40 585
R207 B.n700 B.n699 585
R208 B.n699 B.n36 585
R209 B.n698 B.n35 585
R210 B.n726 B.n35 585
R211 B.n697 B.n34 585
R212 B.n727 B.n34 585
R213 B.n696 B.n33 585
R214 B.n728 B.n33 585
R215 B.n695 B.n694 585
R216 B.n694 B.n29 585
R217 B.n693 B.n28 585
R218 B.n734 B.n28 585
R219 B.n692 B.n27 585
R220 B.n735 B.n27 585
R221 B.n691 B.n26 585
R222 B.n736 B.n26 585
R223 B.n690 B.n689 585
R224 B.n689 B.n25 585
R225 B.n688 B.n21 585
R226 B.n742 B.n21 585
R227 B.n687 B.n20 585
R228 B.n743 B.n20 585
R229 B.n686 B.n19 585
R230 B.n744 B.n19 585
R231 B.n685 B.n684 585
R232 B.n684 B.n18 585
R233 B.n683 B.n14 585
R234 B.n750 B.n14 585
R235 B.n682 B.n13 585
R236 B.n751 B.n13 585
R237 B.n681 B.n12 585
R238 B.n752 B.n12 585
R239 B.n680 B.n679 585
R240 B.n679 B.n8 585
R241 B.n678 B.n7 585
R242 B.n758 B.n7 585
R243 B.n677 B.n6 585
R244 B.n759 B.n6 585
R245 B.n676 B.n5 585
R246 B.n760 B.n5 585
R247 B.n675 B.n674 585
R248 B.n674 B.n4 585
R249 B.n673 B.n300 585
R250 B.n673 B.n672 585
R251 B.n663 B.n301 585
R252 B.n302 B.n301 585
R253 B.n665 B.n664 585
R254 B.n666 B.n665 585
R255 B.n662 B.n307 585
R256 B.n307 B.n306 585
R257 B.n661 B.n660 585
R258 B.n660 B.n659 585
R259 B.n309 B.n308 585
R260 B.n652 B.n309 585
R261 B.n651 B.n650 585
R262 B.n653 B.n651 585
R263 B.n649 B.n314 585
R264 B.n314 B.n313 585
R265 B.n648 B.n647 585
R266 B.n647 B.n646 585
R267 B.n316 B.n315 585
R268 B.n639 B.n316 585
R269 B.n638 B.n637 585
R270 B.n640 B.n638 585
R271 B.n636 B.n321 585
R272 B.n321 B.n320 585
R273 B.n635 B.n634 585
R274 B.n634 B.n633 585
R275 B.n323 B.n322 585
R276 B.n324 B.n323 585
R277 B.n626 B.n625 585
R278 B.n627 B.n626 585
R279 B.n624 B.n329 585
R280 B.n329 B.n328 585
R281 B.n623 B.n622 585
R282 B.n622 B.n621 585
R283 B.n331 B.n330 585
R284 B.n332 B.n331 585
R285 B.n614 B.n613 585
R286 B.n615 B.n614 585
R287 B.n612 B.n336 585
R288 B.n340 B.n336 585
R289 B.n611 B.n610 585
R290 B.n610 B.n609 585
R291 B.n338 B.n337 585
R292 B.n339 B.n338 585
R293 B.n602 B.n601 585
R294 B.n603 B.n602 585
R295 B.n600 B.n345 585
R296 B.n345 B.n344 585
R297 B.n594 B.n593 585
R298 B.n592 B.n396 585
R299 B.n591 B.n395 585
R300 B.n596 B.n395 585
R301 B.n590 B.n589 585
R302 B.n588 B.n587 585
R303 B.n586 B.n585 585
R304 B.n584 B.n583 585
R305 B.n582 B.n581 585
R306 B.n580 B.n579 585
R307 B.n578 B.n577 585
R308 B.n576 B.n575 585
R309 B.n574 B.n573 585
R310 B.n572 B.n571 585
R311 B.n570 B.n569 585
R312 B.n568 B.n567 585
R313 B.n566 B.n565 585
R314 B.n564 B.n563 585
R315 B.n562 B.n561 585
R316 B.n560 B.n559 585
R317 B.n558 B.n557 585
R318 B.n556 B.n555 585
R319 B.n554 B.n553 585
R320 B.n552 B.n551 585
R321 B.n550 B.n549 585
R322 B.n548 B.n547 585
R323 B.n546 B.n545 585
R324 B.n544 B.n543 585
R325 B.n542 B.n541 585
R326 B.n540 B.n539 585
R327 B.n538 B.n537 585
R328 B.n536 B.n535 585
R329 B.n534 B.n533 585
R330 B.n532 B.n531 585
R331 B.n530 B.n529 585
R332 B.n528 B.n527 585
R333 B.n526 B.n525 585
R334 B.n524 B.n523 585
R335 B.n522 B.n521 585
R336 B.n520 B.n519 585
R337 B.n518 B.n517 585
R338 B.n516 B.n515 585
R339 B.n514 B.n513 585
R340 B.n512 B.n511 585
R341 B.n510 B.n509 585
R342 B.n508 B.n507 585
R343 B.n506 B.n505 585
R344 B.n504 B.n503 585
R345 B.n502 B.n501 585
R346 B.n500 B.n499 585
R347 B.n498 B.n497 585
R348 B.n496 B.n495 585
R349 B.n494 B.n493 585
R350 B.n492 B.n491 585
R351 B.n490 B.n489 585
R352 B.n487 B.n486 585
R353 B.n485 B.n484 585
R354 B.n483 B.n482 585
R355 B.n481 B.n480 585
R356 B.n479 B.n478 585
R357 B.n477 B.n476 585
R358 B.n475 B.n474 585
R359 B.n473 B.n472 585
R360 B.n471 B.n470 585
R361 B.n469 B.n468 585
R362 B.n467 B.n466 585
R363 B.n465 B.n464 585
R364 B.n463 B.n462 585
R365 B.n461 B.n460 585
R366 B.n459 B.n458 585
R367 B.n457 B.n456 585
R368 B.n455 B.n454 585
R369 B.n453 B.n452 585
R370 B.n451 B.n450 585
R371 B.n449 B.n448 585
R372 B.n447 B.n446 585
R373 B.n445 B.n444 585
R374 B.n443 B.n442 585
R375 B.n441 B.n440 585
R376 B.n439 B.n438 585
R377 B.n437 B.n436 585
R378 B.n435 B.n434 585
R379 B.n433 B.n432 585
R380 B.n431 B.n430 585
R381 B.n429 B.n428 585
R382 B.n427 B.n426 585
R383 B.n425 B.n424 585
R384 B.n423 B.n422 585
R385 B.n421 B.n420 585
R386 B.n419 B.n418 585
R387 B.n417 B.n416 585
R388 B.n415 B.n414 585
R389 B.n413 B.n412 585
R390 B.n411 B.n410 585
R391 B.n409 B.n408 585
R392 B.n407 B.n406 585
R393 B.n405 B.n404 585
R394 B.n403 B.n402 585
R395 B.n347 B.n346 585
R396 B.n599 B.n598 585
R397 B.n343 B.n342 585
R398 B.n344 B.n343 585
R399 B.n605 B.n604 585
R400 B.n604 B.n603 585
R401 B.n606 B.n341 585
R402 B.n341 B.n339 585
R403 B.n608 B.n607 585
R404 B.n609 B.n608 585
R405 B.n335 B.n334 585
R406 B.n340 B.n335 585
R407 B.n617 B.n616 585
R408 B.n616 B.n615 585
R409 B.n618 B.n333 585
R410 B.n333 B.n332 585
R411 B.n620 B.n619 585
R412 B.n621 B.n620 585
R413 B.n327 B.n326 585
R414 B.n328 B.n327 585
R415 B.n629 B.n628 585
R416 B.n628 B.n627 585
R417 B.n630 B.n325 585
R418 B.n325 B.n324 585
R419 B.n632 B.n631 585
R420 B.n633 B.n632 585
R421 B.n319 B.n318 585
R422 B.n320 B.n319 585
R423 B.n642 B.n641 585
R424 B.n641 B.n640 585
R425 B.n643 B.n317 585
R426 B.n639 B.n317 585
R427 B.n645 B.n644 585
R428 B.n646 B.n645 585
R429 B.n312 B.n311 585
R430 B.n313 B.n312 585
R431 B.n655 B.n654 585
R432 B.n654 B.n653 585
R433 B.n656 B.n310 585
R434 B.n652 B.n310 585
R435 B.n658 B.n657 585
R436 B.n659 B.n658 585
R437 B.n305 B.n304 585
R438 B.n306 B.n305 585
R439 B.n668 B.n667 585
R440 B.n667 B.n666 585
R441 B.n669 B.n303 585
R442 B.n303 B.n302 585
R443 B.n671 B.n670 585
R444 B.n672 B.n671 585
R445 B.n2 B.n0 585
R446 B.n4 B.n2 585
R447 B.n3 B.n1 585
R448 B.n759 B.n3 585
R449 B.n757 B.n756 585
R450 B.n758 B.n757 585
R451 B.n755 B.n9 585
R452 B.n9 B.n8 585
R453 B.n754 B.n753 585
R454 B.n753 B.n752 585
R455 B.n11 B.n10 585
R456 B.n751 B.n11 585
R457 B.n749 B.n748 585
R458 B.n750 B.n749 585
R459 B.n747 B.n15 585
R460 B.n18 B.n15 585
R461 B.n746 B.n745 585
R462 B.n745 B.n744 585
R463 B.n17 B.n16 585
R464 B.n743 B.n17 585
R465 B.n741 B.n740 585
R466 B.n742 B.n741 585
R467 B.n739 B.n22 585
R468 B.n25 B.n22 585
R469 B.n738 B.n737 585
R470 B.n737 B.n736 585
R471 B.n24 B.n23 585
R472 B.n735 B.n24 585
R473 B.n733 B.n732 585
R474 B.n734 B.n733 585
R475 B.n731 B.n30 585
R476 B.n30 B.n29 585
R477 B.n730 B.n729 585
R478 B.n729 B.n728 585
R479 B.n32 B.n31 585
R480 B.n727 B.n32 585
R481 B.n725 B.n724 585
R482 B.n726 B.n725 585
R483 B.n723 B.n37 585
R484 B.n37 B.n36 585
R485 B.n722 B.n721 585
R486 B.n721 B.n720 585
R487 B.n39 B.n38 585
R488 B.n719 B.n39 585
R489 B.n717 B.n716 585
R490 B.n718 B.n717 585
R491 B.n715 B.n44 585
R492 B.n44 B.n43 585
R493 B.n714 B.n713 585
R494 B.n713 B.n712 585
R495 B.n46 B.n45 585
R496 B.n711 B.n46 585
R497 B.n762 B.n761 585
R498 B.n761 B.n760 585
R499 B.n594 B.n343 530.939
R500 B.n104 B.n46 530.939
R501 B.n598 B.n345 530.939
R502 B.n709 B.n48 530.939
R503 B.n710 B.n97 256.663
R504 B.n710 B.n96 256.663
R505 B.n710 B.n95 256.663
R506 B.n710 B.n94 256.663
R507 B.n710 B.n93 256.663
R508 B.n710 B.n92 256.663
R509 B.n710 B.n91 256.663
R510 B.n710 B.n90 256.663
R511 B.n710 B.n89 256.663
R512 B.n710 B.n88 256.663
R513 B.n710 B.n87 256.663
R514 B.n710 B.n86 256.663
R515 B.n710 B.n85 256.663
R516 B.n710 B.n84 256.663
R517 B.n710 B.n83 256.663
R518 B.n710 B.n82 256.663
R519 B.n710 B.n81 256.663
R520 B.n710 B.n80 256.663
R521 B.n710 B.n79 256.663
R522 B.n710 B.n78 256.663
R523 B.n710 B.n77 256.663
R524 B.n710 B.n76 256.663
R525 B.n710 B.n75 256.663
R526 B.n710 B.n74 256.663
R527 B.n710 B.n73 256.663
R528 B.n710 B.n72 256.663
R529 B.n710 B.n71 256.663
R530 B.n710 B.n70 256.663
R531 B.n710 B.n69 256.663
R532 B.n710 B.n68 256.663
R533 B.n710 B.n67 256.663
R534 B.n710 B.n66 256.663
R535 B.n710 B.n65 256.663
R536 B.n710 B.n64 256.663
R537 B.n710 B.n63 256.663
R538 B.n710 B.n62 256.663
R539 B.n710 B.n61 256.663
R540 B.n710 B.n60 256.663
R541 B.n710 B.n59 256.663
R542 B.n710 B.n58 256.663
R543 B.n710 B.n57 256.663
R544 B.n710 B.n56 256.663
R545 B.n710 B.n55 256.663
R546 B.n710 B.n54 256.663
R547 B.n710 B.n53 256.663
R548 B.n710 B.n52 256.663
R549 B.n710 B.n51 256.663
R550 B.n710 B.n50 256.663
R551 B.n710 B.n49 256.663
R552 B.n596 B.n595 256.663
R553 B.n596 B.n348 256.663
R554 B.n596 B.n349 256.663
R555 B.n596 B.n350 256.663
R556 B.n596 B.n351 256.663
R557 B.n596 B.n352 256.663
R558 B.n596 B.n353 256.663
R559 B.n596 B.n354 256.663
R560 B.n596 B.n355 256.663
R561 B.n596 B.n356 256.663
R562 B.n596 B.n357 256.663
R563 B.n596 B.n358 256.663
R564 B.n596 B.n359 256.663
R565 B.n596 B.n360 256.663
R566 B.n596 B.n361 256.663
R567 B.n596 B.n362 256.663
R568 B.n596 B.n363 256.663
R569 B.n596 B.n364 256.663
R570 B.n596 B.n365 256.663
R571 B.n596 B.n366 256.663
R572 B.n596 B.n367 256.663
R573 B.n596 B.n368 256.663
R574 B.n596 B.n369 256.663
R575 B.n596 B.n370 256.663
R576 B.n596 B.n371 256.663
R577 B.n596 B.n372 256.663
R578 B.n596 B.n373 256.663
R579 B.n596 B.n374 256.663
R580 B.n596 B.n375 256.663
R581 B.n596 B.n376 256.663
R582 B.n596 B.n377 256.663
R583 B.n596 B.n378 256.663
R584 B.n596 B.n379 256.663
R585 B.n596 B.n380 256.663
R586 B.n596 B.n381 256.663
R587 B.n596 B.n382 256.663
R588 B.n596 B.n383 256.663
R589 B.n596 B.n384 256.663
R590 B.n596 B.n385 256.663
R591 B.n596 B.n386 256.663
R592 B.n596 B.n387 256.663
R593 B.n596 B.n388 256.663
R594 B.n596 B.n389 256.663
R595 B.n596 B.n390 256.663
R596 B.n596 B.n391 256.663
R597 B.n596 B.n392 256.663
R598 B.n596 B.n393 256.663
R599 B.n596 B.n394 256.663
R600 B.n597 B.n596 256.663
R601 B.n604 B.n343 163.367
R602 B.n604 B.n341 163.367
R603 B.n608 B.n341 163.367
R604 B.n608 B.n335 163.367
R605 B.n616 B.n335 163.367
R606 B.n616 B.n333 163.367
R607 B.n620 B.n333 163.367
R608 B.n620 B.n327 163.367
R609 B.n628 B.n327 163.367
R610 B.n628 B.n325 163.367
R611 B.n632 B.n325 163.367
R612 B.n632 B.n319 163.367
R613 B.n641 B.n319 163.367
R614 B.n641 B.n317 163.367
R615 B.n645 B.n317 163.367
R616 B.n645 B.n312 163.367
R617 B.n654 B.n312 163.367
R618 B.n654 B.n310 163.367
R619 B.n658 B.n310 163.367
R620 B.n658 B.n305 163.367
R621 B.n667 B.n305 163.367
R622 B.n667 B.n303 163.367
R623 B.n671 B.n303 163.367
R624 B.n671 B.n2 163.367
R625 B.n761 B.n2 163.367
R626 B.n761 B.n3 163.367
R627 B.n757 B.n3 163.367
R628 B.n757 B.n9 163.367
R629 B.n753 B.n9 163.367
R630 B.n753 B.n11 163.367
R631 B.n749 B.n11 163.367
R632 B.n749 B.n15 163.367
R633 B.n745 B.n15 163.367
R634 B.n745 B.n17 163.367
R635 B.n741 B.n17 163.367
R636 B.n741 B.n22 163.367
R637 B.n737 B.n22 163.367
R638 B.n737 B.n24 163.367
R639 B.n733 B.n24 163.367
R640 B.n733 B.n30 163.367
R641 B.n729 B.n30 163.367
R642 B.n729 B.n32 163.367
R643 B.n725 B.n32 163.367
R644 B.n725 B.n37 163.367
R645 B.n721 B.n37 163.367
R646 B.n721 B.n39 163.367
R647 B.n717 B.n39 163.367
R648 B.n717 B.n44 163.367
R649 B.n713 B.n44 163.367
R650 B.n713 B.n46 163.367
R651 B.n396 B.n395 163.367
R652 B.n589 B.n395 163.367
R653 B.n587 B.n586 163.367
R654 B.n583 B.n582 163.367
R655 B.n579 B.n578 163.367
R656 B.n575 B.n574 163.367
R657 B.n571 B.n570 163.367
R658 B.n567 B.n566 163.367
R659 B.n563 B.n562 163.367
R660 B.n559 B.n558 163.367
R661 B.n555 B.n554 163.367
R662 B.n551 B.n550 163.367
R663 B.n547 B.n546 163.367
R664 B.n543 B.n542 163.367
R665 B.n539 B.n538 163.367
R666 B.n535 B.n534 163.367
R667 B.n531 B.n530 163.367
R668 B.n527 B.n526 163.367
R669 B.n523 B.n522 163.367
R670 B.n519 B.n518 163.367
R671 B.n515 B.n514 163.367
R672 B.n511 B.n510 163.367
R673 B.n507 B.n506 163.367
R674 B.n503 B.n502 163.367
R675 B.n499 B.n498 163.367
R676 B.n495 B.n494 163.367
R677 B.n491 B.n490 163.367
R678 B.n486 B.n485 163.367
R679 B.n482 B.n481 163.367
R680 B.n478 B.n477 163.367
R681 B.n474 B.n473 163.367
R682 B.n470 B.n469 163.367
R683 B.n466 B.n465 163.367
R684 B.n462 B.n461 163.367
R685 B.n458 B.n457 163.367
R686 B.n454 B.n453 163.367
R687 B.n450 B.n449 163.367
R688 B.n446 B.n445 163.367
R689 B.n442 B.n441 163.367
R690 B.n438 B.n437 163.367
R691 B.n434 B.n433 163.367
R692 B.n430 B.n429 163.367
R693 B.n426 B.n425 163.367
R694 B.n422 B.n421 163.367
R695 B.n418 B.n417 163.367
R696 B.n414 B.n413 163.367
R697 B.n410 B.n409 163.367
R698 B.n406 B.n405 163.367
R699 B.n402 B.n347 163.367
R700 B.n602 B.n345 163.367
R701 B.n602 B.n338 163.367
R702 B.n610 B.n338 163.367
R703 B.n610 B.n336 163.367
R704 B.n614 B.n336 163.367
R705 B.n614 B.n331 163.367
R706 B.n622 B.n331 163.367
R707 B.n622 B.n329 163.367
R708 B.n626 B.n329 163.367
R709 B.n626 B.n323 163.367
R710 B.n634 B.n323 163.367
R711 B.n634 B.n321 163.367
R712 B.n638 B.n321 163.367
R713 B.n638 B.n316 163.367
R714 B.n647 B.n316 163.367
R715 B.n647 B.n314 163.367
R716 B.n651 B.n314 163.367
R717 B.n651 B.n309 163.367
R718 B.n660 B.n309 163.367
R719 B.n660 B.n307 163.367
R720 B.n665 B.n307 163.367
R721 B.n665 B.n301 163.367
R722 B.n673 B.n301 163.367
R723 B.n674 B.n673 163.367
R724 B.n674 B.n5 163.367
R725 B.n6 B.n5 163.367
R726 B.n7 B.n6 163.367
R727 B.n679 B.n7 163.367
R728 B.n679 B.n12 163.367
R729 B.n13 B.n12 163.367
R730 B.n14 B.n13 163.367
R731 B.n684 B.n14 163.367
R732 B.n684 B.n19 163.367
R733 B.n20 B.n19 163.367
R734 B.n21 B.n20 163.367
R735 B.n689 B.n21 163.367
R736 B.n689 B.n26 163.367
R737 B.n27 B.n26 163.367
R738 B.n28 B.n27 163.367
R739 B.n694 B.n28 163.367
R740 B.n694 B.n33 163.367
R741 B.n34 B.n33 163.367
R742 B.n35 B.n34 163.367
R743 B.n699 B.n35 163.367
R744 B.n699 B.n40 163.367
R745 B.n41 B.n40 163.367
R746 B.n42 B.n41 163.367
R747 B.n704 B.n42 163.367
R748 B.n704 B.n47 163.367
R749 B.n48 B.n47 163.367
R750 B.n108 B.n107 163.367
R751 B.n112 B.n111 163.367
R752 B.n116 B.n115 163.367
R753 B.n120 B.n119 163.367
R754 B.n124 B.n123 163.367
R755 B.n128 B.n127 163.367
R756 B.n132 B.n131 163.367
R757 B.n136 B.n135 163.367
R758 B.n140 B.n139 163.367
R759 B.n144 B.n143 163.367
R760 B.n148 B.n147 163.367
R761 B.n152 B.n151 163.367
R762 B.n156 B.n155 163.367
R763 B.n160 B.n159 163.367
R764 B.n164 B.n163 163.367
R765 B.n168 B.n167 163.367
R766 B.n172 B.n171 163.367
R767 B.n176 B.n175 163.367
R768 B.n180 B.n179 163.367
R769 B.n184 B.n183 163.367
R770 B.n188 B.n187 163.367
R771 B.n192 B.n191 163.367
R772 B.n197 B.n196 163.367
R773 B.n201 B.n200 163.367
R774 B.n205 B.n204 163.367
R775 B.n209 B.n208 163.367
R776 B.n213 B.n212 163.367
R777 B.n217 B.n216 163.367
R778 B.n221 B.n220 163.367
R779 B.n225 B.n224 163.367
R780 B.n229 B.n228 163.367
R781 B.n233 B.n232 163.367
R782 B.n237 B.n236 163.367
R783 B.n241 B.n240 163.367
R784 B.n245 B.n244 163.367
R785 B.n249 B.n248 163.367
R786 B.n253 B.n252 163.367
R787 B.n257 B.n256 163.367
R788 B.n261 B.n260 163.367
R789 B.n265 B.n264 163.367
R790 B.n269 B.n268 163.367
R791 B.n273 B.n272 163.367
R792 B.n277 B.n276 163.367
R793 B.n281 B.n280 163.367
R794 B.n285 B.n284 163.367
R795 B.n289 B.n288 163.367
R796 B.n293 B.n292 163.367
R797 B.n297 B.n296 163.367
R798 B.n709 B.n98 163.367
R799 B.n400 B.t18 93.6396
R800 B.n99 B.t13 93.6396
R801 B.n397 B.t21 93.6228
R802 B.n102 B.t10 93.6228
R803 B.n596 B.n344 74.7897
R804 B.n711 B.n710 74.7897
R805 B.n595 B.n594 71.676
R806 B.n589 B.n348 71.676
R807 B.n586 B.n349 71.676
R808 B.n582 B.n350 71.676
R809 B.n578 B.n351 71.676
R810 B.n574 B.n352 71.676
R811 B.n570 B.n353 71.676
R812 B.n566 B.n354 71.676
R813 B.n562 B.n355 71.676
R814 B.n558 B.n356 71.676
R815 B.n554 B.n357 71.676
R816 B.n550 B.n358 71.676
R817 B.n546 B.n359 71.676
R818 B.n542 B.n360 71.676
R819 B.n538 B.n361 71.676
R820 B.n534 B.n362 71.676
R821 B.n530 B.n363 71.676
R822 B.n526 B.n364 71.676
R823 B.n522 B.n365 71.676
R824 B.n518 B.n366 71.676
R825 B.n514 B.n367 71.676
R826 B.n510 B.n368 71.676
R827 B.n506 B.n369 71.676
R828 B.n502 B.n370 71.676
R829 B.n498 B.n371 71.676
R830 B.n494 B.n372 71.676
R831 B.n490 B.n373 71.676
R832 B.n485 B.n374 71.676
R833 B.n481 B.n375 71.676
R834 B.n477 B.n376 71.676
R835 B.n473 B.n377 71.676
R836 B.n469 B.n378 71.676
R837 B.n465 B.n379 71.676
R838 B.n461 B.n380 71.676
R839 B.n457 B.n381 71.676
R840 B.n453 B.n382 71.676
R841 B.n449 B.n383 71.676
R842 B.n445 B.n384 71.676
R843 B.n441 B.n385 71.676
R844 B.n437 B.n386 71.676
R845 B.n433 B.n387 71.676
R846 B.n429 B.n388 71.676
R847 B.n425 B.n389 71.676
R848 B.n421 B.n390 71.676
R849 B.n417 B.n391 71.676
R850 B.n413 B.n392 71.676
R851 B.n409 B.n393 71.676
R852 B.n405 B.n394 71.676
R853 B.n597 B.n347 71.676
R854 B.n104 B.n49 71.676
R855 B.n108 B.n50 71.676
R856 B.n112 B.n51 71.676
R857 B.n116 B.n52 71.676
R858 B.n120 B.n53 71.676
R859 B.n124 B.n54 71.676
R860 B.n128 B.n55 71.676
R861 B.n132 B.n56 71.676
R862 B.n136 B.n57 71.676
R863 B.n140 B.n58 71.676
R864 B.n144 B.n59 71.676
R865 B.n148 B.n60 71.676
R866 B.n152 B.n61 71.676
R867 B.n156 B.n62 71.676
R868 B.n160 B.n63 71.676
R869 B.n164 B.n64 71.676
R870 B.n168 B.n65 71.676
R871 B.n172 B.n66 71.676
R872 B.n176 B.n67 71.676
R873 B.n180 B.n68 71.676
R874 B.n184 B.n69 71.676
R875 B.n188 B.n70 71.676
R876 B.n192 B.n71 71.676
R877 B.n197 B.n72 71.676
R878 B.n201 B.n73 71.676
R879 B.n205 B.n74 71.676
R880 B.n209 B.n75 71.676
R881 B.n213 B.n76 71.676
R882 B.n217 B.n77 71.676
R883 B.n221 B.n78 71.676
R884 B.n225 B.n79 71.676
R885 B.n229 B.n80 71.676
R886 B.n233 B.n81 71.676
R887 B.n237 B.n82 71.676
R888 B.n241 B.n83 71.676
R889 B.n245 B.n84 71.676
R890 B.n249 B.n85 71.676
R891 B.n253 B.n86 71.676
R892 B.n257 B.n87 71.676
R893 B.n261 B.n88 71.676
R894 B.n265 B.n89 71.676
R895 B.n269 B.n90 71.676
R896 B.n273 B.n91 71.676
R897 B.n277 B.n92 71.676
R898 B.n281 B.n93 71.676
R899 B.n285 B.n94 71.676
R900 B.n289 B.n95 71.676
R901 B.n293 B.n96 71.676
R902 B.n297 B.n97 71.676
R903 B.n98 B.n97 71.676
R904 B.n296 B.n96 71.676
R905 B.n292 B.n95 71.676
R906 B.n288 B.n94 71.676
R907 B.n284 B.n93 71.676
R908 B.n280 B.n92 71.676
R909 B.n276 B.n91 71.676
R910 B.n272 B.n90 71.676
R911 B.n268 B.n89 71.676
R912 B.n264 B.n88 71.676
R913 B.n260 B.n87 71.676
R914 B.n256 B.n86 71.676
R915 B.n252 B.n85 71.676
R916 B.n248 B.n84 71.676
R917 B.n244 B.n83 71.676
R918 B.n240 B.n82 71.676
R919 B.n236 B.n81 71.676
R920 B.n232 B.n80 71.676
R921 B.n228 B.n79 71.676
R922 B.n224 B.n78 71.676
R923 B.n220 B.n77 71.676
R924 B.n216 B.n76 71.676
R925 B.n212 B.n75 71.676
R926 B.n208 B.n74 71.676
R927 B.n204 B.n73 71.676
R928 B.n200 B.n72 71.676
R929 B.n196 B.n71 71.676
R930 B.n191 B.n70 71.676
R931 B.n187 B.n69 71.676
R932 B.n183 B.n68 71.676
R933 B.n179 B.n67 71.676
R934 B.n175 B.n66 71.676
R935 B.n171 B.n65 71.676
R936 B.n167 B.n64 71.676
R937 B.n163 B.n63 71.676
R938 B.n159 B.n62 71.676
R939 B.n155 B.n61 71.676
R940 B.n151 B.n60 71.676
R941 B.n147 B.n59 71.676
R942 B.n143 B.n58 71.676
R943 B.n139 B.n57 71.676
R944 B.n135 B.n56 71.676
R945 B.n131 B.n55 71.676
R946 B.n127 B.n54 71.676
R947 B.n123 B.n53 71.676
R948 B.n119 B.n52 71.676
R949 B.n115 B.n51 71.676
R950 B.n111 B.n50 71.676
R951 B.n107 B.n49 71.676
R952 B.n595 B.n396 71.676
R953 B.n587 B.n348 71.676
R954 B.n583 B.n349 71.676
R955 B.n579 B.n350 71.676
R956 B.n575 B.n351 71.676
R957 B.n571 B.n352 71.676
R958 B.n567 B.n353 71.676
R959 B.n563 B.n354 71.676
R960 B.n559 B.n355 71.676
R961 B.n555 B.n356 71.676
R962 B.n551 B.n357 71.676
R963 B.n547 B.n358 71.676
R964 B.n543 B.n359 71.676
R965 B.n539 B.n360 71.676
R966 B.n535 B.n361 71.676
R967 B.n531 B.n362 71.676
R968 B.n527 B.n363 71.676
R969 B.n523 B.n364 71.676
R970 B.n519 B.n365 71.676
R971 B.n515 B.n366 71.676
R972 B.n511 B.n367 71.676
R973 B.n507 B.n368 71.676
R974 B.n503 B.n369 71.676
R975 B.n499 B.n370 71.676
R976 B.n495 B.n371 71.676
R977 B.n491 B.n372 71.676
R978 B.n486 B.n373 71.676
R979 B.n482 B.n374 71.676
R980 B.n478 B.n375 71.676
R981 B.n474 B.n376 71.676
R982 B.n470 B.n377 71.676
R983 B.n466 B.n378 71.676
R984 B.n462 B.n379 71.676
R985 B.n458 B.n380 71.676
R986 B.n454 B.n381 71.676
R987 B.n450 B.n382 71.676
R988 B.n446 B.n383 71.676
R989 B.n442 B.n384 71.676
R990 B.n438 B.n385 71.676
R991 B.n434 B.n386 71.676
R992 B.n430 B.n387 71.676
R993 B.n426 B.n388 71.676
R994 B.n422 B.n389 71.676
R995 B.n418 B.n390 71.676
R996 B.n414 B.n391 71.676
R997 B.n410 B.n392 71.676
R998 B.n406 B.n393 71.676
R999 B.n402 B.n394 71.676
R1000 B.n598 B.n597 71.676
R1001 B.n401 B.t17 71.3365
R1002 B.n100 B.t14 71.3365
R1003 B.n398 B.t20 71.3198
R1004 B.n103 B.t11 71.3198
R1005 B.n488 B.n401 59.5399
R1006 B.n399 B.n398 59.5399
R1007 B.n194 B.n103 59.5399
R1008 B.n101 B.n100 59.5399
R1009 B.n603 B.n344 40.6858
R1010 B.n603 B.n339 40.6858
R1011 B.n609 B.n339 40.6858
R1012 B.n609 B.n340 40.6858
R1013 B.n615 B.n332 40.6858
R1014 B.n621 B.n332 40.6858
R1015 B.n621 B.n328 40.6858
R1016 B.n627 B.n328 40.6858
R1017 B.n627 B.n324 40.6858
R1018 B.n633 B.n324 40.6858
R1019 B.n640 B.n320 40.6858
R1020 B.n640 B.n639 40.6858
R1021 B.n646 B.n313 40.6858
R1022 B.n653 B.n313 40.6858
R1023 B.n653 B.n652 40.6858
R1024 B.n659 B.n306 40.6858
R1025 B.n666 B.n306 40.6858
R1026 B.n672 B.n302 40.6858
R1027 B.n672 B.n4 40.6858
R1028 B.n760 B.n4 40.6858
R1029 B.n760 B.n759 40.6858
R1030 B.n759 B.n758 40.6858
R1031 B.n758 B.n8 40.6858
R1032 B.n752 B.n751 40.6858
R1033 B.n751 B.n750 40.6858
R1034 B.n744 B.n18 40.6858
R1035 B.n744 B.n743 40.6858
R1036 B.n743 B.n742 40.6858
R1037 B.n736 B.n25 40.6858
R1038 B.n736 B.n735 40.6858
R1039 B.n734 B.n29 40.6858
R1040 B.n728 B.n29 40.6858
R1041 B.n728 B.n727 40.6858
R1042 B.n727 B.n726 40.6858
R1043 B.n726 B.n36 40.6858
R1044 B.n720 B.n36 40.6858
R1045 B.n719 B.n718 40.6858
R1046 B.n718 B.n43 40.6858
R1047 B.n712 B.n43 40.6858
R1048 B.n712 B.n711 40.6858
R1049 B.n340 B.t16 39.4892
R1050 B.t9 B.n719 39.4892
R1051 B.n639 B.t3 38.2926
R1052 B.n25 B.t0 38.2926
R1053 B.n105 B.n45 34.4981
R1054 B.n708 B.n707 34.4981
R1055 B.n600 B.n599 34.4981
R1056 B.n593 B.n342 34.4981
R1057 B.n666 B.t7 28.7196
R1058 B.n752 B.t5 28.7196
R1059 B.n659 B.t6 27.5229
R1060 B.n750 B.t1 27.5229
R1061 B.n633 B.t2 22.7364
R1062 B.t4 B.n734 22.7364
R1063 B.n401 B.n400 22.3035
R1064 B.n398 B.n397 22.3035
R1065 B.n103 B.n102 22.3035
R1066 B.n100 B.n99 22.3035
R1067 B B.n762 18.0485
R1068 B.t2 B.n320 17.9499
R1069 B.n735 B.t4 17.9499
R1070 B.n652 B.t6 13.1634
R1071 B.n18 B.t1 13.1634
R1072 B.t7 B.n302 11.9668
R1073 B.t5 B.n8 11.9668
R1074 B.n106 B.n105 10.6151
R1075 B.n109 B.n106 10.6151
R1076 B.n110 B.n109 10.6151
R1077 B.n113 B.n110 10.6151
R1078 B.n114 B.n113 10.6151
R1079 B.n117 B.n114 10.6151
R1080 B.n118 B.n117 10.6151
R1081 B.n121 B.n118 10.6151
R1082 B.n122 B.n121 10.6151
R1083 B.n125 B.n122 10.6151
R1084 B.n126 B.n125 10.6151
R1085 B.n129 B.n126 10.6151
R1086 B.n130 B.n129 10.6151
R1087 B.n133 B.n130 10.6151
R1088 B.n134 B.n133 10.6151
R1089 B.n137 B.n134 10.6151
R1090 B.n138 B.n137 10.6151
R1091 B.n141 B.n138 10.6151
R1092 B.n142 B.n141 10.6151
R1093 B.n145 B.n142 10.6151
R1094 B.n146 B.n145 10.6151
R1095 B.n149 B.n146 10.6151
R1096 B.n150 B.n149 10.6151
R1097 B.n153 B.n150 10.6151
R1098 B.n154 B.n153 10.6151
R1099 B.n157 B.n154 10.6151
R1100 B.n158 B.n157 10.6151
R1101 B.n161 B.n158 10.6151
R1102 B.n162 B.n161 10.6151
R1103 B.n165 B.n162 10.6151
R1104 B.n166 B.n165 10.6151
R1105 B.n169 B.n166 10.6151
R1106 B.n170 B.n169 10.6151
R1107 B.n173 B.n170 10.6151
R1108 B.n174 B.n173 10.6151
R1109 B.n177 B.n174 10.6151
R1110 B.n178 B.n177 10.6151
R1111 B.n181 B.n178 10.6151
R1112 B.n182 B.n181 10.6151
R1113 B.n185 B.n182 10.6151
R1114 B.n186 B.n185 10.6151
R1115 B.n189 B.n186 10.6151
R1116 B.n190 B.n189 10.6151
R1117 B.n193 B.n190 10.6151
R1118 B.n198 B.n195 10.6151
R1119 B.n199 B.n198 10.6151
R1120 B.n202 B.n199 10.6151
R1121 B.n203 B.n202 10.6151
R1122 B.n206 B.n203 10.6151
R1123 B.n207 B.n206 10.6151
R1124 B.n210 B.n207 10.6151
R1125 B.n211 B.n210 10.6151
R1126 B.n215 B.n214 10.6151
R1127 B.n218 B.n215 10.6151
R1128 B.n219 B.n218 10.6151
R1129 B.n222 B.n219 10.6151
R1130 B.n223 B.n222 10.6151
R1131 B.n226 B.n223 10.6151
R1132 B.n227 B.n226 10.6151
R1133 B.n230 B.n227 10.6151
R1134 B.n231 B.n230 10.6151
R1135 B.n234 B.n231 10.6151
R1136 B.n235 B.n234 10.6151
R1137 B.n238 B.n235 10.6151
R1138 B.n239 B.n238 10.6151
R1139 B.n242 B.n239 10.6151
R1140 B.n243 B.n242 10.6151
R1141 B.n246 B.n243 10.6151
R1142 B.n247 B.n246 10.6151
R1143 B.n250 B.n247 10.6151
R1144 B.n251 B.n250 10.6151
R1145 B.n254 B.n251 10.6151
R1146 B.n255 B.n254 10.6151
R1147 B.n258 B.n255 10.6151
R1148 B.n259 B.n258 10.6151
R1149 B.n262 B.n259 10.6151
R1150 B.n263 B.n262 10.6151
R1151 B.n266 B.n263 10.6151
R1152 B.n267 B.n266 10.6151
R1153 B.n270 B.n267 10.6151
R1154 B.n271 B.n270 10.6151
R1155 B.n274 B.n271 10.6151
R1156 B.n275 B.n274 10.6151
R1157 B.n278 B.n275 10.6151
R1158 B.n279 B.n278 10.6151
R1159 B.n282 B.n279 10.6151
R1160 B.n283 B.n282 10.6151
R1161 B.n286 B.n283 10.6151
R1162 B.n287 B.n286 10.6151
R1163 B.n290 B.n287 10.6151
R1164 B.n291 B.n290 10.6151
R1165 B.n294 B.n291 10.6151
R1166 B.n295 B.n294 10.6151
R1167 B.n298 B.n295 10.6151
R1168 B.n299 B.n298 10.6151
R1169 B.n708 B.n299 10.6151
R1170 B.n601 B.n600 10.6151
R1171 B.n601 B.n337 10.6151
R1172 B.n611 B.n337 10.6151
R1173 B.n612 B.n611 10.6151
R1174 B.n613 B.n612 10.6151
R1175 B.n613 B.n330 10.6151
R1176 B.n623 B.n330 10.6151
R1177 B.n624 B.n623 10.6151
R1178 B.n625 B.n624 10.6151
R1179 B.n625 B.n322 10.6151
R1180 B.n635 B.n322 10.6151
R1181 B.n636 B.n635 10.6151
R1182 B.n637 B.n636 10.6151
R1183 B.n637 B.n315 10.6151
R1184 B.n648 B.n315 10.6151
R1185 B.n649 B.n648 10.6151
R1186 B.n650 B.n649 10.6151
R1187 B.n650 B.n308 10.6151
R1188 B.n661 B.n308 10.6151
R1189 B.n662 B.n661 10.6151
R1190 B.n664 B.n662 10.6151
R1191 B.n664 B.n663 10.6151
R1192 B.n663 B.n300 10.6151
R1193 B.n675 B.n300 10.6151
R1194 B.n676 B.n675 10.6151
R1195 B.n677 B.n676 10.6151
R1196 B.n678 B.n677 10.6151
R1197 B.n680 B.n678 10.6151
R1198 B.n681 B.n680 10.6151
R1199 B.n682 B.n681 10.6151
R1200 B.n683 B.n682 10.6151
R1201 B.n685 B.n683 10.6151
R1202 B.n686 B.n685 10.6151
R1203 B.n687 B.n686 10.6151
R1204 B.n688 B.n687 10.6151
R1205 B.n690 B.n688 10.6151
R1206 B.n691 B.n690 10.6151
R1207 B.n692 B.n691 10.6151
R1208 B.n693 B.n692 10.6151
R1209 B.n695 B.n693 10.6151
R1210 B.n696 B.n695 10.6151
R1211 B.n697 B.n696 10.6151
R1212 B.n698 B.n697 10.6151
R1213 B.n700 B.n698 10.6151
R1214 B.n701 B.n700 10.6151
R1215 B.n702 B.n701 10.6151
R1216 B.n703 B.n702 10.6151
R1217 B.n705 B.n703 10.6151
R1218 B.n706 B.n705 10.6151
R1219 B.n707 B.n706 10.6151
R1220 B.n593 B.n592 10.6151
R1221 B.n592 B.n591 10.6151
R1222 B.n591 B.n590 10.6151
R1223 B.n590 B.n588 10.6151
R1224 B.n588 B.n585 10.6151
R1225 B.n585 B.n584 10.6151
R1226 B.n584 B.n581 10.6151
R1227 B.n581 B.n580 10.6151
R1228 B.n580 B.n577 10.6151
R1229 B.n577 B.n576 10.6151
R1230 B.n576 B.n573 10.6151
R1231 B.n573 B.n572 10.6151
R1232 B.n572 B.n569 10.6151
R1233 B.n569 B.n568 10.6151
R1234 B.n568 B.n565 10.6151
R1235 B.n565 B.n564 10.6151
R1236 B.n564 B.n561 10.6151
R1237 B.n561 B.n560 10.6151
R1238 B.n560 B.n557 10.6151
R1239 B.n557 B.n556 10.6151
R1240 B.n556 B.n553 10.6151
R1241 B.n553 B.n552 10.6151
R1242 B.n552 B.n549 10.6151
R1243 B.n549 B.n548 10.6151
R1244 B.n548 B.n545 10.6151
R1245 B.n545 B.n544 10.6151
R1246 B.n544 B.n541 10.6151
R1247 B.n541 B.n540 10.6151
R1248 B.n540 B.n537 10.6151
R1249 B.n537 B.n536 10.6151
R1250 B.n536 B.n533 10.6151
R1251 B.n533 B.n532 10.6151
R1252 B.n532 B.n529 10.6151
R1253 B.n529 B.n528 10.6151
R1254 B.n528 B.n525 10.6151
R1255 B.n525 B.n524 10.6151
R1256 B.n524 B.n521 10.6151
R1257 B.n521 B.n520 10.6151
R1258 B.n520 B.n517 10.6151
R1259 B.n517 B.n516 10.6151
R1260 B.n516 B.n513 10.6151
R1261 B.n513 B.n512 10.6151
R1262 B.n512 B.n509 10.6151
R1263 B.n509 B.n508 10.6151
R1264 B.n505 B.n504 10.6151
R1265 B.n504 B.n501 10.6151
R1266 B.n501 B.n500 10.6151
R1267 B.n500 B.n497 10.6151
R1268 B.n497 B.n496 10.6151
R1269 B.n496 B.n493 10.6151
R1270 B.n493 B.n492 10.6151
R1271 B.n492 B.n489 10.6151
R1272 B.n487 B.n484 10.6151
R1273 B.n484 B.n483 10.6151
R1274 B.n483 B.n480 10.6151
R1275 B.n480 B.n479 10.6151
R1276 B.n479 B.n476 10.6151
R1277 B.n476 B.n475 10.6151
R1278 B.n475 B.n472 10.6151
R1279 B.n472 B.n471 10.6151
R1280 B.n471 B.n468 10.6151
R1281 B.n468 B.n467 10.6151
R1282 B.n467 B.n464 10.6151
R1283 B.n464 B.n463 10.6151
R1284 B.n463 B.n460 10.6151
R1285 B.n460 B.n459 10.6151
R1286 B.n459 B.n456 10.6151
R1287 B.n456 B.n455 10.6151
R1288 B.n455 B.n452 10.6151
R1289 B.n452 B.n451 10.6151
R1290 B.n451 B.n448 10.6151
R1291 B.n448 B.n447 10.6151
R1292 B.n447 B.n444 10.6151
R1293 B.n444 B.n443 10.6151
R1294 B.n443 B.n440 10.6151
R1295 B.n440 B.n439 10.6151
R1296 B.n439 B.n436 10.6151
R1297 B.n436 B.n435 10.6151
R1298 B.n435 B.n432 10.6151
R1299 B.n432 B.n431 10.6151
R1300 B.n431 B.n428 10.6151
R1301 B.n428 B.n427 10.6151
R1302 B.n427 B.n424 10.6151
R1303 B.n424 B.n423 10.6151
R1304 B.n423 B.n420 10.6151
R1305 B.n420 B.n419 10.6151
R1306 B.n419 B.n416 10.6151
R1307 B.n416 B.n415 10.6151
R1308 B.n415 B.n412 10.6151
R1309 B.n412 B.n411 10.6151
R1310 B.n411 B.n408 10.6151
R1311 B.n408 B.n407 10.6151
R1312 B.n407 B.n404 10.6151
R1313 B.n404 B.n403 10.6151
R1314 B.n403 B.n346 10.6151
R1315 B.n599 B.n346 10.6151
R1316 B.n605 B.n342 10.6151
R1317 B.n606 B.n605 10.6151
R1318 B.n607 B.n606 10.6151
R1319 B.n607 B.n334 10.6151
R1320 B.n617 B.n334 10.6151
R1321 B.n618 B.n617 10.6151
R1322 B.n619 B.n618 10.6151
R1323 B.n619 B.n326 10.6151
R1324 B.n629 B.n326 10.6151
R1325 B.n630 B.n629 10.6151
R1326 B.n631 B.n630 10.6151
R1327 B.n631 B.n318 10.6151
R1328 B.n642 B.n318 10.6151
R1329 B.n643 B.n642 10.6151
R1330 B.n644 B.n643 10.6151
R1331 B.n644 B.n311 10.6151
R1332 B.n655 B.n311 10.6151
R1333 B.n656 B.n655 10.6151
R1334 B.n657 B.n656 10.6151
R1335 B.n657 B.n304 10.6151
R1336 B.n668 B.n304 10.6151
R1337 B.n669 B.n668 10.6151
R1338 B.n670 B.n669 10.6151
R1339 B.n670 B.n0 10.6151
R1340 B.n756 B.n1 10.6151
R1341 B.n756 B.n755 10.6151
R1342 B.n755 B.n754 10.6151
R1343 B.n754 B.n10 10.6151
R1344 B.n748 B.n10 10.6151
R1345 B.n748 B.n747 10.6151
R1346 B.n747 B.n746 10.6151
R1347 B.n746 B.n16 10.6151
R1348 B.n740 B.n16 10.6151
R1349 B.n740 B.n739 10.6151
R1350 B.n739 B.n738 10.6151
R1351 B.n738 B.n23 10.6151
R1352 B.n732 B.n23 10.6151
R1353 B.n732 B.n731 10.6151
R1354 B.n731 B.n730 10.6151
R1355 B.n730 B.n31 10.6151
R1356 B.n724 B.n31 10.6151
R1357 B.n724 B.n723 10.6151
R1358 B.n723 B.n722 10.6151
R1359 B.n722 B.n38 10.6151
R1360 B.n716 B.n38 10.6151
R1361 B.n716 B.n715 10.6151
R1362 B.n715 B.n714 10.6151
R1363 B.n714 B.n45 10.6151
R1364 B.n195 B.n194 6.5566
R1365 B.n211 B.n101 6.5566
R1366 B.n505 B.n399 6.5566
R1367 B.n489 B.n488 6.5566
R1368 B.n194 B.n193 4.05904
R1369 B.n214 B.n101 4.05904
R1370 B.n508 B.n399 4.05904
R1371 B.n488 B.n487 4.05904
R1372 B.n762 B.n0 2.81026
R1373 B.n762 B.n1 2.81026
R1374 B.n646 B.t3 2.39376
R1375 B.n742 B.t0 2.39376
R1376 B.n615 B.t16 1.19713
R1377 B.n720 B.t9 1.19713
R1378 VP.n7 VP.t4 452.738
R1379 VP.n17 VP.t6 433.507
R1380 VP.n29 VP.t0 433.507
R1381 VP.n15 VP.t3 433.507
R1382 VP.n22 VP.t5 385.307
R1383 VP.n1 VP.t1 385.307
R1384 VP.n5 VP.t7 385.307
R1385 VP.n8 VP.t2 385.307
R1386 VP.n30 VP.n29 161.3
R1387 VP.n9 VP.n6 161.3
R1388 VP.n11 VP.n10 161.3
R1389 VP.n13 VP.n12 161.3
R1390 VP.n14 VP.n4 161.3
R1391 VP.n16 VP.n15 161.3
R1392 VP.n28 VP.n0 161.3
R1393 VP.n27 VP.n26 161.3
R1394 VP.n25 VP.n24 161.3
R1395 VP.n23 VP.n2 161.3
R1396 VP.n21 VP.n20 161.3
R1397 VP.n19 VP.n3 161.3
R1398 VP.n18 VP.n17 161.3
R1399 VP.n24 VP.n23 56.5193
R1400 VP.n10 VP.n9 56.5193
R1401 VP.n21 VP.n3 50.2061
R1402 VP.n28 VP.n27 50.2061
R1403 VP.n14 VP.n13 50.2061
R1404 VP.n18 VP.n16 43.3717
R1405 VP.n7 VP.n6 43.2015
R1406 VP.n8 VP.n7 38.5669
R1407 VP.n23 VP.n22 15.9041
R1408 VP.n24 VP.n1 15.9041
R1409 VP.n10 VP.n5 15.9041
R1410 VP.n9 VP.n8 15.9041
R1411 VP.n17 VP.n3 9.49444
R1412 VP.n29 VP.n28 9.49444
R1413 VP.n15 VP.n14 9.49444
R1414 VP.n22 VP.n21 8.56395
R1415 VP.n27 VP.n1 8.56395
R1416 VP.n13 VP.n5 8.56395
R1417 VP.n11 VP.n6 0.189894
R1418 VP.n12 VP.n11 0.189894
R1419 VP.n12 VP.n4 0.189894
R1420 VP.n16 VP.n4 0.189894
R1421 VP.n19 VP.n18 0.189894
R1422 VP.n20 VP.n19 0.189894
R1423 VP.n20 VP.n2 0.189894
R1424 VP.n25 VP.n2 0.189894
R1425 VP.n26 VP.n25 0.189894
R1426 VP.n26 VP.n0 0.189894
R1427 VP.n30 VP.n0 0.189894
R1428 VP VP.n30 0.0516364
R1429 VDD1 VDD1.n0 60.4337
R1430 VDD1.n3 VDD1.n2 60.3201
R1431 VDD1.n3 VDD1.n1 60.3201
R1432 VDD1.n5 VDD1.n4 59.8797
R1433 VDD1.n5 VDD1.n3 40.0612
R1434 VDD1.n4 VDD1.t0 1.5108
R1435 VDD1.n4 VDD1.t4 1.5108
R1436 VDD1.n0 VDD1.t3 1.5108
R1437 VDD1.n0 VDD1.t5 1.5108
R1438 VDD1.n2 VDD1.t6 1.5108
R1439 VDD1.n2 VDD1.t7 1.5108
R1440 VDD1.n1 VDD1.t1 1.5108
R1441 VDD1.n1 VDD1.t2 1.5108
R1442 VDD1 VDD1.n5 0.438
C0 VDD2 VTAIL 11.141299f
C1 VDD2 VDD1 0.884393f
C2 VDD2 VN 6.4746f
C3 VDD2 VP 0.330059f
C4 VTAIL VDD1 11.0988f
C5 VN VTAIL 6.2352f
C6 VTAIL VP 6.24931f
C7 VN VDD1 0.148309f
C8 VDD1 VP 6.65585f
C9 VN VP 5.69277f
C10 VDD2 B 3.69569f
C11 VDD1 B 3.944253f
C12 VTAIL B 9.681495f
C13 VN B 9.11153f
C14 VP B 7.177876f
C15 VDD1.t3 B 0.277771f
C16 VDD1.t5 B 0.277771f
C17 VDD1.n0 B 2.48869f
C18 VDD1.t1 B 0.277771f
C19 VDD1.t2 B 0.277771f
C20 VDD1.n1 B 2.48794f
C21 VDD1.t6 B 0.277771f
C22 VDD1.t7 B 0.277771f
C23 VDD1.n2 B 2.48794f
C24 VDD1.n3 B 2.54513f
C25 VDD1.t0 B 0.277771f
C26 VDD1.t4 B 0.277771f
C27 VDD1.n4 B 2.48528f
C28 VDD1.n5 B 2.63034f
C29 VP.n0 B 0.041855f
C30 VP.t1 B 1.2289f
C31 VP.n1 B 0.458827f
C32 VP.n2 B 0.041855f
C33 VP.t5 B 1.2289f
C34 VP.n3 B 0.01521f
C35 VP.n4 B 0.041855f
C36 VP.t3 B 1.28148f
C37 VP.t7 B 1.2289f
C38 VP.n5 B 0.458827f
C39 VP.n6 B 0.17353f
C40 VP.t2 B 1.2289f
C41 VP.t4 B 1.30304f
C42 VP.n7 B 0.501728f
C43 VP.n8 B 0.500108f
C44 VP.n9 B 0.047619f
C45 VP.n10 B 0.047619f
C46 VP.n11 B 0.041855f
C47 VP.n12 B 0.041855f
C48 VP.n13 B 0.051784f
C49 VP.n14 B 0.01521f
C50 VP.n15 B 0.496719f
C51 VP.n16 B 1.82164f
C52 VP.t6 B 1.28148f
C53 VP.n17 B 0.496719f
C54 VP.n18 B 1.85633f
C55 VP.n19 B 0.041855f
C56 VP.n20 B 0.041855f
C57 VP.n21 B 0.051784f
C58 VP.n22 B 0.458827f
C59 VP.n23 B 0.047619f
C60 VP.n24 B 0.047619f
C61 VP.n25 B 0.041855f
C62 VP.n26 B 0.041855f
C63 VP.n27 B 0.051784f
C64 VP.n28 B 0.01521f
C65 VP.t0 B 1.28148f
C66 VP.n29 B 0.496719f
C67 VP.n30 B 0.032436f
C68 VTAIL.t14 B 0.201832f
C69 VTAIL.t12 B 0.201832f
C70 VTAIL.n0 B 1.74389f
C71 VTAIL.n1 B 0.265552f
C72 VTAIL.t15 B 2.22365f
C73 VTAIL.n2 B 0.362084f
C74 VTAIL.t7 B 2.22365f
C75 VTAIL.n3 B 0.362084f
C76 VTAIL.t3 B 0.201832f
C77 VTAIL.t6 B 0.201832f
C78 VTAIL.n4 B 1.74389f
C79 VTAIL.n5 B 0.324134f
C80 VTAIL.t2 B 2.22365f
C81 VTAIL.n6 B 1.36893f
C82 VTAIL.t8 B 2.22365f
C83 VTAIL.n7 B 1.36893f
C84 VTAIL.t13 B 0.201832f
C85 VTAIL.t11 B 0.201832f
C86 VTAIL.n8 B 1.74389f
C87 VTAIL.n9 B 0.324135f
C88 VTAIL.t9 B 2.22365f
C89 VTAIL.n10 B 0.362078f
C90 VTAIL.t5 B 2.22365f
C91 VTAIL.n11 B 0.362078f
C92 VTAIL.t1 B 0.201832f
C93 VTAIL.t0 B 0.201832f
C94 VTAIL.n12 B 1.74389f
C95 VTAIL.n13 B 0.324135f
C96 VTAIL.t4 B 2.22365f
C97 VTAIL.n14 B 1.36893f
C98 VTAIL.t10 B 2.22365f
C99 VTAIL.n15 B 1.36528f
C100 VDD2.t7 B 0.276187f
C101 VDD2.t1 B 0.276187f
C102 VDD2.n0 B 2.47375f
C103 VDD2.t5 B 0.276187f
C104 VDD2.t4 B 0.276187f
C105 VDD2.n1 B 2.47375f
C106 VDD2.n2 B 2.47389f
C107 VDD2.t3 B 0.276187f
C108 VDD2.t6 B 0.276187f
C109 VDD2.n3 B 2.47112f
C110 VDD2.n4 B 2.58358f
C111 VDD2.t0 B 0.276187f
C112 VDD2.t2 B 0.276187f
C113 VDD2.n5 B 2.47371f
C114 VN.n0 B 0.041274f
C115 VN.t3 B 1.21185f
C116 VN.n1 B 0.452463f
C117 VN.n2 B 0.171123f
C118 VN.t1 B 1.21185f
C119 VN.t0 B 1.28496f
C120 VN.n3 B 0.494768f
C121 VN.n4 B 0.49317f
C122 VN.n5 B 0.046958f
C123 VN.n6 B 0.046958f
C124 VN.n7 B 0.041274f
C125 VN.n8 B 0.041274f
C126 VN.n9 B 0.051065f
C127 VN.n10 B 0.014999f
C128 VN.t5 B 1.2637f
C129 VN.n11 B 0.489828f
C130 VN.n12 B 0.031986f
C131 VN.n13 B 0.041274f
C132 VN.t2 B 1.21185f
C133 VN.n14 B 0.452463f
C134 VN.n15 B 0.171123f
C135 VN.t4 B 1.21185f
C136 VN.t6 B 1.28496f
C137 VN.n16 B 0.494768f
C138 VN.n17 B 0.49317f
C139 VN.n18 B 0.046958f
C140 VN.n19 B 0.046958f
C141 VN.n20 B 0.041274f
C142 VN.n21 B 0.041274f
C143 VN.n22 B 0.051065f
C144 VN.n23 B 0.014999f
C145 VN.t7 B 1.2637f
C146 VN.n24 B 0.489828f
C147 VN.n25 B 1.82342f
.ends

