* NGSPICE file created from diff_pair_sample_1284.ext - technology: sky130A

.subckt diff_pair_sample_1284 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1636_n1732# sky130_fd_pr__pfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=0.78
X1 VTAIL.t7 VP.t0 VDD1.t3 w_n1636_n1732# sky130_fd_pr__pfet_01v8 ad=1.4898 pd=8.42 as=0.6303 ps=4.15 w=3.82 l=0.78
X2 B.t8 B.t6 B.t7 w_n1636_n1732# sky130_fd_pr__pfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=0.78
X3 VDD1.t0 VP.t1 VTAIL.t6 w_n1636_n1732# sky130_fd_pr__pfet_01v8 ad=0.6303 pd=4.15 as=1.4898 ps=8.42 w=3.82 l=0.78
X4 B.t5 B.t3 B.t4 w_n1636_n1732# sky130_fd_pr__pfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=0.78
X5 VDD2.t3 VN.t0 VTAIL.t3 w_n1636_n1732# sky130_fd_pr__pfet_01v8 ad=0.6303 pd=4.15 as=1.4898 ps=8.42 w=3.82 l=0.78
X6 VDD1.t2 VP.t2 VTAIL.t5 w_n1636_n1732# sky130_fd_pr__pfet_01v8 ad=0.6303 pd=4.15 as=1.4898 ps=8.42 w=3.82 l=0.78
X7 VTAIL.t0 VN.t1 VDD2.t2 w_n1636_n1732# sky130_fd_pr__pfet_01v8 ad=1.4898 pd=8.42 as=0.6303 ps=4.15 w=3.82 l=0.78
X8 VTAIL.t1 VN.t2 VDD2.t1 w_n1636_n1732# sky130_fd_pr__pfet_01v8 ad=1.4898 pd=8.42 as=0.6303 ps=4.15 w=3.82 l=0.78
X9 VDD2.t0 VN.t3 VTAIL.t2 w_n1636_n1732# sky130_fd_pr__pfet_01v8 ad=0.6303 pd=4.15 as=1.4898 ps=8.42 w=3.82 l=0.78
X10 B.t2 B.t0 B.t1 w_n1636_n1732# sky130_fd_pr__pfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=0.78
X11 VTAIL.t4 VP.t3 VDD1.t1 w_n1636_n1732# sky130_fd_pr__pfet_01v8 ad=1.4898 pd=8.42 as=0.6303 ps=4.15 w=3.82 l=0.78
R0 B.n243 B.n242 585
R1 B.n244 B.n37 585
R2 B.n246 B.n245 585
R3 B.n247 B.n36 585
R4 B.n249 B.n248 585
R5 B.n250 B.n35 585
R6 B.n252 B.n251 585
R7 B.n253 B.n34 585
R8 B.n255 B.n254 585
R9 B.n256 B.n33 585
R10 B.n258 B.n257 585
R11 B.n259 B.n32 585
R12 B.n261 B.n260 585
R13 B.n262 B.n31 585
R14 B.n264 B.n263 585
R15 B.n265 B.n30 585
R16 B.n267 B.n266 585
R17 B.n268 B.n27 585
R18 B.n271 B.n270 585
R19 B.n272 B.n26 585
R20 B.n274 B.n273 585
R21 B.n275 B.n25 585
R22 B.n277 B.n276 585
R23 B.n278 B.n24 585
R24 B.n280 B.n279 585
R25 B.n281 B.n23 585
R26 B.n283 B.n282 585
R27 B.n285 B.n284 585
R28 B.n286 B.n19 585
R29 B.n288 B.n287 585
R30 B.n289 B.n18 585
R31 B.n291 B.n290 585
R32 B.n292 B.n17 585
R33 B.n294 B.n293 585
R34 B.n295 B.n16 585
R35 B.n297 B.n296 585
R36 B.n298 B.n15 585
R37 B.n300 B.n299 585
R38 B.n301 B.n14 585
R39 B.n303 B.n302 585
R40 B.n304 B.n13 585
R41 B.n306 B.n305 585
R42 B.n307 B.n12 585
R43 B.n309 B.n308 585
R44 B.n310 B.n11 585
R45 B.n241 B.n38 585
R46 B.n240 B.n239 585
R47 B.n238 B.n39 585
R48 B.n237 B.n236 585
R49 B.n235 B.n40 585
R50 B.n234 B.n233 585
R51 B.n232 B.n41 585
R52 B.n231 B.n230 585
R53 B.n229 B.n42 585
R54 B.n228 B.n227 585
R55 B.n226 B.n43 585
R56 B.n225 B.n224 585
R57 B.n223 B.n44 585
R58 B.n222 B.n221 585
R59 B.n220 B.n45 585
R60 B.n219 B.n218 585
R61 B.n217 B.n46 585
R62 B.n216 B.n215 585
R63 B.n214 B.n47 585
R64 B.n213 B.n212 585
R65 B.n211 B.n48 585
R66 B.n210 B.n209 585
R67 B.n208 B.n49 585
R68 B.n207 B.n206 585
R69 B.n205 B.n50 585
R70 B.n204 B.n203 585
R71 B.n202 B.n51 585
R72 B.n201 B.n200 585
R73 B.n199 B.n52 585
R74 B.n198 B.n197 585
R75 B.n196 B.n53 585
R76 B.n195 B.n194 585
R77 B.n193 B.n54 585
R78 B.n192 B.n191 585
R79 B.n190 B.n55 585
R80 B.n189 B.n188 585
R81 B.n187 B.n56 585
R82 B.n118 B.n83 585
R83 B.n120 B.n119 585
R84 B.n121 B.n82 585
R85 B.n123 B.n122 585
R86 B.n124 B.n81 585
R87 B.n126 B.n125 585
R88 B.n127 B.n80 585
R89 B.n129 B.n128 585
R90 B.n130 B.n79 585
R91 B.n132 B.n131 585
R92 B.n133 B.n78 585
R93 B.n135 B.n134 585
R94 B.n136 B.n77 585
R95 B.n138 B.n137 585
R96 B.n139 B.n76 585
R97 B.n141 B.n140 585
R98 B.n142 B.n75 585
R99 B.n144 B.n143 585
R100 B.n146 B.n145 585
R101 B.n147 B.n71 585
R102 B.n149 B.n148 585
R103 B.n150 B.n70 585
R104 B.n152 B.n151 585
R105 B.n153 B.n69 585
R106 B.n155 B.n154 585
R107 B.n156 B.n68 585
R108 B.n158 B.n157 585
R109 B.n160 B.n65 585
R110 B.n162 B.n161 585
R111 B.n163 B.n64 585
R112 B.n165 B.n164 585
R113 B.n166 B.n63 585
R114 B.n168 B.n167 585
R115 B.n169 B.n62 585
R116 B.n171 B.n170 585
R117 B.n172 B.n61 585
R118 B.n174 B.n173 585
R119 B.n175 B.n60 585
R120 B.n177 B.n176 585
R121 B.n178 B.n59 585
R122 B.n180 B.n179 585
R123 B.n181 B.n58 585
R124 B.n183 B.n182 585
R125 B.n184 B.n57 585
R126 B.n186 B.n185 585
R127 B.n117 B.n116 585
R128 B.n115 B.n84 585
R129 B.n114 B.n113 585
R130 B.n112 B.n85 585
R131 B.n111 B.n110 585
R132 B.n109 B.n86 585
R133 B.n108 B.n107 585
R134 B.n106 B.n87 585
R135 B.n105 B.n104 585
R136 B.n103 B.n88 585
R137 B.n102 B.n101 585
R138 B.n100 B.n89 585
R139 B.n99 B.n98 585
R140 B.n97 B.n90 585
R141 B.n96 B.n95 585
R142 B.n94 B.n91 585
R143 B.n93 B.n92 585
R144 B.n2 B.n0 585
R145 B.n337 B.n1 585
R146 B.n336 B.n335 585
R147 B.n334 B.n3 585
R148 B.n333 B.n332 585
R149 B.n331 B.n4 585
R150 B.n330 B.n329 585
R151 B.n328 B.n5 585
R152 B.n327 B.n326 585
R153 B.n325 B.n6 585
R154 B.n324 B.n323 585
R155 B.n322 B.n7 585
R156 B.n321 B.n320 585
R157 B.n319 B.n8 585
R158 B.n318 B.n317 585
R159 B.n316 B.n9 585
R160 B.n315 B.n314 585
R161 B.n313 B.n10 585
R162 B.n312 B.n311 585
R163 B.n339 B.n338 585
R164 B.n116 B.n83 458.866
R165 B.n312 B.n11 458.866
R166 B.n187 B.n186 458.866
R167 B.n242 B.n241 458.866
R168 B.n66 B.t6 320.111
R169 B.n72 B.t0 320.111
R170 B.n20 B.t9 320.111
R171 B.n28 B.t3 320.111
R172 B.n66 B.t8 253.666
R173 B.n28 B.t4 253.666
R174 B.n72 B.t2 253.666
R175 B.n20 B.t10 253.666
R176 B.n67 B.t7 232.138
R177 B.n29 B.t5 232.138
R178 B.n73 B.t1 232.138
R179 B.n21 B.t11 232.138
R180 B.n116 B.n115 163.367
R181 B.n115 B.n114 163.367
R182 B.n114 B.n85 163.367
R183 B.n110 B.n85 163.367
R184 B.n110 B.n109 163.367
R185 B.n109 B.n108 163.367
R186 B.n108 B.n87 163.367
R187 B.n104 B.n87 163.367
R188 B.n104 B.n103 163.367
R189 B.n103 B.n102 163.367
R190 B.n102 B.n89 163.367
R191 B.n98 B.n89 163.367
R192 B.n98 B.n97 163.367
R193 B.n97 B.n96 163.367
R194 B.n96 B.n91 163.367
R195 B.n92 B.n91 163.367
R196 B.n92 B.n2 163.367
R197 B.n338 B.n2 163.367
R198 B.n338 B.n337 163.367
R199 B.n337 B.n336 163.367
R200 B.n336 B.n3 163.367
R201 B.n332 B.n3 163.367
R202 B.n332 B.n331 163.367
R203 B.n331 B.n330 163.367
R204 B.n330 B.n5 163.367
R205 B.n326 B.n5 163.367
R206 B.n326 B.n325 163.367
R207 B.n325 B.n324 163.367
R208 B.n324 B.n7 163.367
R209 B.n320 B.n7 163.367
R210 B.n320 B.n319 163.367
R211 B.n319 B.n318 163.367
R212 B.n318 B.n9 163.367
R213 B.n314 B.n9 163.367
R214 B.n314 B.n313 163.367
R215 B.n313 B.n312 163.367
R216 B.n120 B.n83 163.367
R217 B.n121 B.n120 163.367
R218 B.n122 B.n121 163.367
R219 B.n122 B.n81 163.367
R220 B.n126 B.n81 163.367
R221 B.n127 B.n126 163.367
R222 B.n128 B.n127 163.367
R223 B.n128 B.n79 163.367
R224 B.n132 B.n79 163.367
R225 B.n133 B.n132 163.367
R226 B.n134 B.n133 163.367
R227 B.n134 B.n77 163.367
R228 B.n138 B.n77 163.367
R229 B.n139 B.n138 163.367
R230 B.n140 B.n139 163.367
R231 B.n140 B.n75 163.367
R232 B.n144 B.n75 163.367
R233 B.n145 B.n144 163.367
R234 B.n145 B.n71 163.367
R235 B.n149 B.n71 163.367
R236 B.n150 B.n149 163.367
R237 B.n151 B.n150 163.367
R238 B.n151 B.n69 163.367
R239 B.n155 B.n69 163.367
R240 B.n156 B.n155 163.367
R241 B.n157 B.n156 163.367
R242 B.n157 B.n65 163.367
R243 B.n162 B.n65 163.367
R244 B.n163 B.n162 163.367
R245 B.n164 B.n163 163.367
R246 B.n164 B.n63 163.367
R247 B.n168 B.n63 163.367
R248 B.n169 B.n168 163.367
R249 B.n170 B.n169 163.367
R250 B.n170 B.n61 163.367
R251 B.n174 B.n61 163.367
R252 B.n175 B.n174 163.367
R253 B.n176 B.n175 163.367
R254 B.n176 B.n59 163.367
R255 B.n180 B.n59 163.367
R256 B.n181 B.n180 163.367
R257 B.n182 B.n181 163.367
R258 B.n182 B.n57 163.367
R259 B.n186 B.n57 163.367
R260 B.n188 B.n187 163.367
R261 B.n188 B.n55 163.367
R262 B.n192 B.n55 163.367
R263 B.n193 B.n192 163.367
R264 B.n194 B.n193 163.367
R265 B.n194 B.n53 163.367
R266 B.n198 B.n53 163.367
R267 B.n199 B.n198 163.367
R268 B.n200 B.n199 163.367
R269 B.n200 B.n51 163.367
R270 B.n204 B.n51 163.367
R271 B.n205 B.n204 163.367
R272 B.n206 B.n205 163.367
R273 B.n206 B.n49 163.367
R274 B.n210 B.n49 163.367
R275 B.n211 B.n210 163.367
R276 B.n212 B.n211 163.367
R277 B.n212 B.n47 163.367
R278 B.n216 B.n47 163.367
R279 B.n217 B.n216 163.367
R280 B.n218 B.n217 163.367
R281 B.n218 B.n45 163.367
R282 B.n222 B.n45 163.367
R283 B.n223 B.n222 163.367
R284 B.n224 B.n223 163.367
R285 B.n224 B.n43 163.367
R286 B.n228 B.n43 163.367
R287 B.n229 B.n228 163.367
R288 B.n230 B.n229 163.367
R289 B.n230 B.n41 163.367
R290 B.n234 B.n41 163.367
R291 B.n235 B.n234 163.367
R292 B.n236 B.n235 163.367
R293 B.n236 B.n39 163.367
R294 B.n240 B.n39 163.367
R295 B.n241 B.n240 163.367
R296 B.n308 B.n11 163.367
R297 B.n308 B.n307 163.367
R298 B.n307 B.n306 163.367
R299 B.n306 B.n13 163.367
R300 B.n302 B.n13 163.367
R301 B.n302 B.n301 163.367
R302 B.n301 B.n300 163.367
R303 B.n300 B.n15 163.367
R304 B.n296 B.n15 163.367
R305 B.n296 B.n295 163.367
R306 B.n295 B.n294 163.367
R307 B.n294 B.n17 163.367
R308 B.n290 B.n17 163.367
R309 B.n290 B.n289 163.367
R310 B.n289 B.n288 163.367
R311 B.n288 B.n19 163.367
R312 B.n284 B.n19 163.367
R313 B.n284 B.n283 163.367
R314 B.n283 B.n23 163.367
R315 B.n279 B.n23 163.367
R316 B.n279 B.n278 163.367
R317 B.n278 B.n277 163.367
R318 B.n277 B.n25 163.367
R319 B.n273 B.n25 163.367
R320 B.n273 B.n272 163.367
R321 B.n272 B.n271 163.367
R322 B.n271 B.n27 163.367
R323 B.n266 B.n27 163.367
R324 B.n266 B.n265 163.367
R325 B.n265 B.n264 163.367
R326 B.n264 B.n31 163.367
R327 B.n260 B.n31 163.367
R328 B.n260 B.n259 163.367
R329 B.n259 B.n258 163.367
R330 B.n258 B.n33 163.367
R331 B.n254 B.n33 163.367
R332 B.n254 B.n253 163.367
R333 B.n253 B.n252 163.367
R334 B.n252 B.n35 163.367
R335 B.n248 B.n35 163.367
R336 B.n248 B.n247 163.367
R337 B.n247 B.n246 163.367
R338 B.n246 B.n37 163.367
R339 B.n242 B.n37 163.367
R340 B.n159 B.n67 59.5399
R341 B.n74 B.n73 59.5399
R342 B.n22 B.n21 59.5399
R343 B.n269 B.n29 59.5399
R344 B.n311 B.n310 29.8151
R345 B.n243 B.n38 29.8151
R346 B.n185 B.n56 29.8151
R347 B.n118 B.n117 29.8151
R348 B.n67 B.n66 21.5278
R349 B.n73 B.n72 21.5278
R350 B.n21 B.n20 21.5278
R351 B.n29 B.n28 21.5278
R352 B B.n339 18.0485
R353 B.n310 B.n309 10.6151
R354 B.n309 B.n12 10.6151
R355 B.n305 B.n12 10.6151
R356 B.n305 B.n304 10.6151
R357 B.n304 B.n303 10.6151
R358 B.n303 B.n14 10.6151
R359 B.n299 B.n14 10.6151
R360 B.n299 B.n298 10.6151
R361 B.n298 B.n297 10.6151
R362 B.n297 B.n16 10.6151
R363 B.n293 B.n16 10.6151
R364 B.n293 B.n292 10.6151
R365 B.n292 B.n291 10.6151
R366 B.n291 B.n18 10.6151
R367 B.n287 B.n18 10.6151
R368 B.n287 B.n286 10.6151
R369 B.n286 B.n285 10.6151
R370 B.n282 B.n281 10.6151
R371 B.n281 B.n280 10.6151
R372 B.n280 B.n24 10.6151
R373 B.n276 B.n24 10.6151
R374 B.n276 B.n275 10.6151
R375 B.n275 B.n274 10.6151
R376 B.n274 B.n26 10.6151
R377 B.n270 B.n26 10.6151
R378 B.n268 B.n267 10.6151
R379 B.n267 B.n30 10.6151
R380 B.n263 B.n30 10.6151
R381 B.n263 B.n262 10.6151
R382 B.n262 B.n261 10.6151
R383 B.n261 B.n32 10.6151
R384 B.n257 B.n32 10.6151
R385 B.n257 B.n256 10.6151
R386 B.n256 B.n255 10.6151
R387 B.n255 B.n34 10.6151
R388 B.n251 B.n34 10.6151
R389 B.n251 B.n250 10.6151
R390 B.n250 B.n249 10.6151
R391 B.n249 B.n36 10.6151
R392 B.n245 B.n36 10.6151
R393 B.n245 B.n244 10.6151
R394 B.n244 B.n243 10.6151
R395 B.n189 B.n56 10.6151
R396 B.n190 B.n189 10.6151
R397 B.n191 B.n190 10.6151
R398 B.n191 B.n54 10.6151
R399 B.n195 B.n54 10.6151
R400 B.n196 B.n195 10.6151
R401 B.n197 B.n196 10.6151
R402 B.n197 B.n52 10.6151
R403 B.n201 B.n52 10.6151
R404 B.n202 B.n201 10.6151
R405 B.n203 B.n202 10.6151
R406 B.n203 B.n50 10.6151
R407 B.n207 B.n50 10.6151
R408 B.n208 B.n207 10.6151
R409 B.n209 B.n208 10.6151
R410 B.n209 B.n48 10.6151
R411 B.n213 B.n48 10.6151
R412 B.n214 B.n213 10.6151
R413 B.n215 B.n214 10.6151
R414 B.n215 B.n46 10.6151
R415 B.n219 B.n46 10.6151
R416 B.n220 B.n219 10.6151
R417 B.n221 B.n220 10.6151
R418 B.n221 B.n44 10.6151
R419 B.n225 B.n44 10.6151
R420 B.n226 B.n225 10.6151
R421 B.n227 B.n226 10.6151
R422 B.n227 B.n42 10.6151
R423 B.n231 B.n42 10.6151
R424 B.n232 B.n231 10.6151
R425 B.n233 B.n232 10.6151
R426 B.n233 B.n40 10.6151
R427 B.n237 B.n40 10.6151
R428 B.n238 B.n237 10.6151
R429 B.n239 B.n238 10.6151
R430 B.n239 B.n38 10.6151
R431 B.n119 B.n118 10.6151
R432 B.n119 B.n82 10.6151
R433 B.n123 B.n82 10.6151
R434 B.n124 B.n123 10.6151
R435 B.n125 B.n124 10.6151
R436 B.n125 B.n80 10.6151
R437 B.n129 B.n80 10.6151
R438 B.n130 B.n129 10.6151
R439 B.n131 B.n130 10.6151
R440 B.n131 B.n78 10.6151
R441 B.n135 B.n78 10.6151
R442 B.n136 B.n135 10.6151
R443 B.n137 B.n136 10.6151
R444 B.n137 B.n76 10.6151
R445 B.n141 B.n76 10.6151
R446 B.n142 B.n141 10.6151
R447 B.n143 B.n142 10.6151
R448 B.n147 B.n146 10.6151
R449 B.n148 B.n147 10.6151
R450 B.n148 B.n70 10.6151
R451 B.n152 B.n70 10.6151
R452 B.n153 B.n152 10.6151
R453 B.n154 B.n153 10.6151
R454 B.n154 B.n68 10.6151
R455 B.n158 B.n68 10.6151
R456 B.n161 B.n160 10.6151
R457 B.n161 B.n64 10.6151
R458 B.n165 B.n64 10.6151
R459 B.n166 B.n165 10.6151
R460 B.n167 B.n166 10.6151
R461 B.n167 B.n62 10.6151
R462 B.n171 B.n62 10.6151
R463 B.n172 B.n171 10.6151
R464 B.n173 B.n172 10.6151
R465 B.n173 B.n60 10.6151
R466 B.n177 B.n60 10.6151
R467 B.n178 B.n177 10.6151
R468 B.n179 B.n178 10.6151
R469 B.n179 B.n58 10.6151
R470 B.n183 B.n58 10.6151
R471 B.n184 B.n183 10.6151
R472 B.n185 B.n184 10.6151
R473 B.n117 B.n84 10.6151
R474 B.n113 B.n84 10.6151
R475 B.n113 B.n112 10.6151
R476 B.n112 B.n111 10.6151
R477 B.n111 B.n86 10.6151
R478 B.n107 B.n86 10.6151
R479 B.n107 B.n106 10.6151
R480 B.n106 B.n105 10.6151
R481 B.n105 B.n88 10.6151
R482 B.n101 B.n88 10.6151
R483 B.n101 B.n100 10.6151
R484 B.n100 B.n99 10.6151
R485 B.n99 B.n90 10.6151
R486 B.n95 B.n90 10.6151
R487 B.n95 B.n94 10.6151
R488 B.n94 B.n93 10.6151
R489 B.n93 B.n0 10.6151
R490 B.n335 B.n1 10.6151
R491 B.n335 B.n334 10.6151
R492 B.n334 B.n333 10.6151
R493 B.n333 B.n4 10.6151
R494 B.n329 B.n4 10.6151
R495 B.n329 B.n328 10.6151
R496 B.n328 B.n327 10.6151
R497 B.n327 B.n6 10.6151
R498 B.n323 B.n6 10.6151
R499 B.n323 B.n322 10.6151
R500 B.n322 B.n321 10.6151
R501 B.n321 B.n8 10.6151
R502 B.n317 B.n8 10.6151
R503 B.n317 B.n316 10.6151
R504 B.n316 B.n315 10.6151
R505 B.n315 B.n10 10.6151
R506 B.n311 B.n10 10.6151
R507 B.n282 B.n22 6.5566
R508 B.n270 B.n269 6.5566
R509 B.n146 B.n74 6.5566
R510 B.n159 B.n158 6.5566
R511 B.n285 B.n22 4.05904
R512 B.n269 B.n268 4.05904
R513 B.n143 B.n74 4.05904
R514 B.n160 B.n159 4.05904
R515 B.n339 B.n0 2.81026
R516 B.n339 B.n1 2.81026
R517 VP.n1 VP.t3 189.387
R518 VP.n1 VP.t1 189.339
R519 VP.n3 VP.t0 168.392
R520 VP.n5 VP.t2 168.392
R521 VP.n6 VP.n5 161.3
R522 VP.n4 VP.n0 161.3
R523 VP.n3 VP.n2 161.3
R524 VP.n2 VP.n1 79.1772
R525 VP.n4 VP.n3 24.1005
R526 VP.n5 VP.n4 24.1005
R527 VP.n2 VP.n0 0.189894
R528 VP.n6 VP.n0 0.189894
R529 VP VP.n6 0.0516364
R530 VDD1 VDD1.n1 143.583
R531 VDD1 VDD1.n0 113.239
R532 VDD1.n0 VDD1.t1 8.50966
R533 VDD1.n0 VDD1.t0 8.50966
R534 VDD1.n1 VDD1.t3 8.50966
R535 VDD1.n1 VDD1.t2 8.50966
R536 VTAIL.n154 VTAIL.n140 756.745
R537 VTAIL.n14 VTAIL.n0 756.745
R538 VTAIL.n34 VTAIL.n20 756.745
R539 VTAIL.n54 VTAIL.n40 756.745
R540 VTAIL.n134 VTAIL.n120 756.745
R541 VTAIL.n114 VTAIL.n100 756.745
R542 VTAIL.n94 VTAIL.n80 756.745
R543 VTAIL.n74 VTAIL.n60 756.745
R544 VTAIL.n147 VTAIL.n146 585
R545 VTAIL.n144 VTAIL.n143 585
R546 VTAIL.n153 VTAIL.n152 585
R547 VTAIL.n155 VTAIL.n154 585
R548 VTAIL.n7 VTAIL.n6 585
R549 VTAIL.n4 VTAIL.n3 585
R550 VTAIL.n13 VTAIL.n12 585
R551 VTAIL.n15 VTAIL.n14 585
R552 VTAIL.n27 VTAIL.n26 585
R553 VTAIL.n24 VTAIL.n23 585
R554 VTAIL.n33 VTAIL.n32 585
R555 VTAIL.n35 VTAIL.n34 585
R556 VTAIL.n47 VTAIL.n46 585
R557 VTAIL.n44 VTAIL.n43 585
R558 VTAIL.n53 VTAIL.n52 585
R559 VTAIL.n55 VTAIL.n54 585
R560 VTAIL.n135 VTAIL.n134 585
R561 VTAIL.n133 VTAIL.n132 585
R562 VTAIL.n124 VTAIL.n123 585
R563 VTAIL.n127 VTAIL.n126 585
R564 VTAIL.n115 VTAIL.n114 585
R565 VTAIL.n113 VTAIL.n112 585
R566 VTAIL.n104 VTAIL.n103 585
R567 VTAIL.n107 VTAIL.n106 585
R568 VTAIL.n95 VTAIL.n94 585
R569 VTAIL.n93 VTAIL.n92 585
R570 VTAIL.n84 VTAIL.n83 585
R571 VTAIL.n87 VTAIL.n86 585
R572 VTAIL.n75 VTAIL.n74 585
R573 VTAIL.n73 VTAIL.n72 585
R574 VTAIL.n64 VTAIL.n63 585
R575 VTAIL.n67 VTAIL.n66 585
R576 VTAIL.t2 VTAIL.n145 330.707
R577 VTAIL.t0 VTAIL.n5 330.707
R578 VTAIL.t5 VTAIL.n25 330.707
R579 VTAIL.t7 VTAIL.n45 330.707
R580 VTAIL.t6 VTAIL.n125 330.707
R581 VTAIL.t4 VTAIL.n105 330.707
R582 VTAIL.t3 VTAIL.n85 330.707
R583 VTAIL.t1 VTAIL.n65 330.707
R584 VTAIL.n146 VTAIL.n143 171.744
R585 VTAIL.n153 VTAIL.n143 171.744
R586 VTAIL.n154 VTAIL.n153 171.744
R587 VTAIL.n6 VTAIL.n3 171.744
R588 VTAIL.n13 VTAIL.n3 171.744
R589 VTAIL.n14 VTAIL.n13 171.744
R590 VTAIL.n26 VTAIL.n23 171.744
R591 VTAIL.n33 VTAIL.n23 171.744
R592 VTAIL.n34 VTAIL.n33 171.744
R593 VTAIL.n46 VTAIL.n43 171.744
R594 VTAIL.n53 VTAIL.n43 171.744
R595 VTAIL.n54 VTAIL.n53 171.744
R596 VTAIL.n134 VTAIL.n133 171.744
R597 VTAIL.n133 VTAIL.n123 171.744
R598 VTAIL.n126 VTAIL.n123 171.744
R599 VTAIL.n114 VTAIL.n113 171.744
R600 VTAIL.n113 VTAIL.n103 171.744
R601 VTAIL.n106 VTAIL.n103 171.744
R602 VTAIL.n94 VTAIL.n93 171.744
R603 VTAIL.n93 VTAIL.n83 171.744
R604 VTAIL.n86 VTAIL.n83 171.744
R605 VTAIL.n74 VTAIL.n73 171.744
R606 VTAIL.n73 VTAIL.n63 171.744
R607 VTAIL.n66 VTAIL.n63 171.744
R608 VTAIL.n146 VTAIL.t2 85.8723
R609 VTAIL.n6 VTAIL.t0 85.8723
R610 VTAIL.n26 VTAIL.t5 85.8723
R611 VTAIL.n46 VTAIL.t7 85.8723
R612 VTAIL.n126 VTAIL.t6 85.8723
R613 VTAIL.n106 VTAIL.t4 85.8723
R614 VTAIL.n86 VTAIL.t3 85.8723
R615 VTAIL.n66 VTAIL.t1 85.8723
R616 VTAIL.n159 VTAIL.n158 31.7975
R617 VTAIL.n19 VTAIL.n18 31.7975
R618 VTAIL.n39 VTAIL.n38 31.7975
R619 VTAIL.n59 VTAIL.n58 31.7975
R620 VTAIL.n139 VTAIL.n138 31.7975
R621 VTAIL.n119 VTAIL.n118 31.7975
R622 VTAIL.n99 VTAIL.n98 31.7975
R623 VTAIL.n79 VTAIL.n78 31.7975
R624 VTAIL.n159 VTAIL.n139 16.6169
R625 VTAIL.n79 VTAIL.n59 16.6169
R626 VTAIL.n147 VTAIL.n145 16.3201
R627 VTAIL.n7 VTAIL.n5 16.3201
R628 VTAIL.n27 VTAIL.n25 16.3201
R629 VTAIL.n47 VTAIL.n45 16.3201
R630 VTAIL.n127 VTAIL.n125 16.3201
R631 VTAIL.n107 VTAIL.n105 16.3201
R632 VTAIL.n87 VTAIL.n85 16.3201
R633 VTAIL.n67 VTAIL.n65 16.3201
R634 VTAIL.n148 VTAIL.n144 12.8005
R635 VTAIL.n8 VTAIL.n4 12.8005
R636 VTAIL.n28 VTAIL.n24 12.8005
R637 VTAIL.n48 VTAIL.n44 12.8005
R638 VTAIL.n128 VTAIL.n124 12.8005
R639 VTAIL.n108 VTAIL.n104 12.8005
R640 VTAIL.n88 VTAIL.n84 12.8005
R641 VTAIL.n68 VTAIL.n64 12.8005
R642 VTAIL.n152 VTAIL.n151 12.0247
R643 VTAIL.n12 VTAIL.n11 12.0247
R644 VTAIL.n32 VTAIL.n31 12.0247
R645 VTAIL.n52 VTAIL.n51 12.0247
R646 VTAIL.n132 VTAIL.n131 12.0247
R647 VTAIL.n112 VTAIL.n111 12.0247
R648 VTAIL.n92 VTAIL.n91 12.0247
R649 VTAIL.n72 VTAIL.n71 12.0247
R650 VTAIL.n155 VTAIL.n142 11.249
R651 VTAIL.n15 VTAIL.n2 11.249
R652 VTAIL.n35 VTAIL.n22 11.249
R653 VTAIL.n55 VTAIL.n42 11.249
R654 VTAIL.n135 VTAIL.n122 11.249
R655 VTAIL.n115 VTAIL.n102 11.249
R656 VTAIL.n95 VTAIL.n82 11.249
R657 VTAIL.n75 VTAIL.n62 11.249
R658 VTAIL.n156 VTAIL.n140 10.4732
R659 VTAIL.n16 VTAIL.n0 10.4732
R660 VTAIL.n36 VTAIL.n20 10.4732
R661 VTAIL.n56 VTAIL.n40 10.4732
R662 VTAIL.n136 VTAIL.n120 10.4732
R663 VTAIL.n116 VTAIL.n100 10.4732
R664 VTAIL.n96 VTAIL.n80 10.4732
R665 VTAIL.n76 VTAIL.n60 10.4732
R666 VTAIL.n158 VTAIL.n157 9.45567
R667 VTAIL.n18 VTAIL.n17 9.45567
R668 VTAIL.n38 VTAIL.n37 9.45567
R669 VTAIL.n58 VTAIL.n57 9.45567
R670 VTAIL.n138 VTAIL.n137 9.45567
R671 VTAIL.n118 VTAIL.n117 9.45567
R672 VTAIL.n98 VTAIL.n97 9.45567
R673 VTAIL.n78 VTAIL.n77 9.45567
R674 VTAIL.n157 VTAIL.n156 9.3005
R675 VTAIL.n142 VTAIL.n141 9.3005
R676 VTAIL.n151 VTAIL.n150 9.3005
R677 VTAIL.n149 VTAIL.n148 9.3005
R678 VTAIL.n17 VTAIL.n16 9.3005
R679 VTAIL.n2 VTAIL.n1 9.3005
R680 VTAIL.n11 VTAIL.n10 9.3005
R681 VTAIL.n9 VTAIL.n8 9.3005
R682 VTAIL.n37 VTAIL.n36 9.3005
R683 VTAIL.n22 VTAIL.n21 9.3005
R684 VTAIL.n31 VTAIL.n30 9.3005
R685 VTAIL.n29 VTAIL.n28 9.3005
R686 VTAIL.n57 VTAIL.n56 9.3005
R687 VTAIL.n42 VTAIL.n41 9.3005
R688 VTAIL.n51 VTAIL.n50 9.3005
R689 VTAIL.n49 VTAIL.n48 9.3005
R690 VTAIL.n137 VTAIL.n136 9.3005
R691 VTAIL.n122 VTAIL.n121 9.3005
R692 VTAIL.n131 VTAIL.n130 9.3005
R693 VTAIL.n129 VTAIL.n128 9.3005
R694 VTAIL.n117 VTAIL.n116 9.3005
R695 VTAIL.n102 VTAIL.n101 9.3005
R696 VTAIL.n111 VTAIL.n110 9.3005
R697 VTAIL.n109 VTAIL.n108 9.3005
R698 VTAIL.n97 VTAIL.n96 9.3005
R699 VTAIL.n82 VTAIL.n81 9.3005
R700 VTAIL.n91 VTAIL.n90 9.3005
R701 VTAIL.n89 VTAIL.n88 9.3005
R702 VTAIL.n77 VTAIL.n76 9.3005
R703 VTAIL.n62 VTAIL.n61 9.3005
R704 VTAIL.n71 VTAIL.n70 9.3005
R705 VTAIL.n69 VTAIL.n68 9.3005
R706 VTAIL.n149 VTAIL.n145 3.78097
R707 VTAIL.n9 VTAIL.n5 3.78097
R708 VTAIL.n29 VTAIL.n25 3.78097
R709 VTAIL.n49 VTAIL.n45 3.78097
R710 VTAIL.n129 VTAIL.n125 3.78097
R711 VTAIL.n109 VTAIL.n105 3.78097
R712 VTAIL.n89 VTAIL.n85 3.78097
R713 VTAIL.n69 VTAIL.n65 3.78097
R714 VTAIL.n158 VTAIL.n140 3.49141
R715 VTAIL.n18 VTAIL.n0 3.49141
R716 VTAIL.n38 VTAIL.n20 3.49141
R717 VTAIL.n58 VTAIL.n40 3.49141
R718 VTAIL.n138 VTAIL.n120 3.49141
R719 VTAIL.n118 VTAIL.n100 3.49141
R720 VTAIL.n98 VTAIL.n80 3.49141
R721 VTAIL.n78 VTAIL.n60 3.49141
R722 VTAIL.n156 VTAIL.n155 2.71565
R723 VTAIL.n16 VTAIL.n15 2.71565
R724 VTAIL.n36 VTAIL.n35 2.71565
R725 VTAIL.n56 VTAIL.n55 2.71565
R726 VTAIL.n136 VTAIL.n135 2.71565
R727 VTAIL.n116 VTAIL.n115 2.71565
R728 VTAIL.n96 VTAIL.n95 2.71565
R729 VTAIL.n76 VTAIL.n75 2.71565
R730 VTAIL.n152 VTAIL.n142 1.93989
R731 VTAIL.n12 VTAIL.n2 1.93989
R732 VTAIL.n32 VTAIL.n22 1.93989
R733 VTAIL.n52 VTAIL.n42 1.93989
R734 VTAIL.n132 VTAIL.n122 1.93989
R735 VTAIL.n112 VTAIL.n102 1.93989
R736 VTAIL.n92 VTAIL.n82 1.93989
R737 VTAIL.n72 VTAIL.n62 1.93989
R738 VTAIL.n151 VTAIL.n144 1.16414
R739 VTAIL.n11 VTAIL.n4 1.16414
R740 VTAIL.n31 VTAIL.n24 1.16414
R741 VTAIL.n51 VTAIL.n44 1.16414
R742 VTAIL.n131 VTAIL.n124 1.16414
R743 VTAIL.n111 VTAIL.n104 1.16414
R744 VTAIL.n91 VTAIL.n84 1.16414
R745 VTAIL.n71 VTAIL.n64 1.16414
R746 VTAIL.n99 VTAIL.n79 0.957397
R747 VTAIL.n139 VTAIL.n119 0.957397
R748 VTAIL.n59 VTAIL.n39 0.957397
R749 VTAIL VTAIL.n19 0.537138
R750 VTAIL.n119 VTAIL.n99 0.470328
R751 VTAIL.n39 VTAIL.n19 0.470328
R752 VTAIL VTAIL.n159 0.420759
R753 VTAIL.n148 VTAIL.n147 0.388379
R754 VTAIL.n8 VTAIL.n7 0.388379
R755 VTAIL.n28 VTAIL.n27 0.388379
R756 VTAIL.n48 VTAIL.n47 0.388379
R757 VTAIL.n128 VTAIL.n127 0.388379
R758 VTAIL.n108 VTAIL.n107 0.388379
R759 VTAIL.n88 VTAIL.n87 0.388379
R760 VTAIL.n68 VTAIL.n67 0.388379
R761 VTAIL.n150 VTAIL.n149 0.155672
R762 VTAIL.n150 VTAIL.n141 0.155672
R763 VTAIL.n157 VTAIL.n141 0.155672
R764 VTAIL.n10 VTAIL.n9 0.155672
R765 VTAIL.n10 VTAIL.n1 0.155672
R766 VTAIL.n17 VTAIL.n1 0.155672
R767 VTAIL.n30 VTAIL.n29 0.155672
R768 VTAIL.n30 VTAIL.n21 0.155672
R769 VTAIL.n37 VTAIL.n21 0.155672
R770 VTAIL.n50 VTAIL.n49 0.155672
R771 VTAIL.n50 VTAIL.n41 0.155672
R772 VTAIL.n57 VTAIL.n41 0.155672
R773 VTAIL.n137 VTAIL.n121 0.155672
R774 VTAIL.n130 VTAIL.n121 0.155672
R775 VTAIL.n130 VTAIL.n129 0.155672
R776 VTAIL.n117 VTAIL.n101 0.155672
R777 VTAIL.n110 VTAIL.n101 0.155672
R778 VTAIL.n110 VTAIL.n109 0.155672
R779 VTAIL.n97 VTAIL.n81 0.155672
R780 VTAIL.n90 VTAIL.n81 0.155672
R781 VTAIL.n90 VTAIL.n89 0.155672
R782 VTAIL.n77 VTAIL.n61 0.155672
R783 VTAIL.n70 VTAIL.n61 0.155672
R784 VTAIL.n70 VTAIL.n69 0.155672
R785 VN.n0 VN.t1 189.387
R786 VN.n1 VN.t0 189.387
R787 VN.n0 VN.t3 189.339
R788 VN.n1 VN.t2 189.339
R789 VN VN.n1 79.5579
R790 VN VN.n0 44.7132
R791 VDD2.n2 VDD2.n0 143.059
R792 VDD2.n2 VDD2.n1 113.18
R793 VDD2.n1 VDD2.t1 8.50966
R794 VDD2.n1 VDD2.t3 8.50966
R795 VDD2.n0 VDD2.t2 8.50966
R796 VDD2.n0 VDD2.t0 8.50966
R797 VDD2 VDD2.n2 0.0586897
C0 B VN 0.664189f
C1 VTAIL VN 1.27448f
C2 w_n1636_n1732# VN 2.26753f
C3 B VP 0.996853f
C4 VTAIL VP 1.28859f
C5 w_n1636_n1732# VP 2.47212f
C6 B VDD2 0.742128f
C7 VDD2 VTAIL 3.15374f
C8 VDD2 w_n1636_n1732# 0.873516f
C9 B VDD1 0.719386f
C10 VTAIL VDD1 3.11174f
C11 VDD1 w_n1636_n1732# 0.857764f
C12 VP VN 3.36746f
C13 VDD2 VN 1.25658f
C14 VDD2 VP 0.283379f
C15 B VTAIL 1.62402f
C16 B w_n1636_n1732# 4.7104f
C17 VTAIL w_n1636_n1732# 2.0272f
C18 VDD1 VN 0.151873f
C19 VDD1 VP 1.38745f
C20 VDD2 VDD1 0.584849f
C21 VDD2 VSUBS 0.454718f
C22 VDD1 VSUBS 2.623691f
C23 VTAIL VSUBS 0.405204f
C24 VN VSUBS 4.00767f
C25 VP VSUBS 0.93498f
C26 B VSUBS 1.909519f
C27 w_n1636_n1732# VSUBS 35.7106f
C28 VDD2.t2 VSUBS 0.060034f
C29 VDD2.t0 VSUBS 0.060034f
C30 VDD2.n0 VSUBS 0.528944f
C31 VDD2.t1 VSUBS 0.060034f
C32 VDD2.t3 VSUBS 0.060034f
C33 VDD2.n1 VSUBS 0.345449f
C34 VDD2.n2 VSUBS 2.01987f
C35 VN.t1 VSUBS 0.446924f
C36 VN.t3 VSUBS 0.44685f
C37 VN.n0 VSUBS 0.400743f
C38 VN.t0 VSUBS 0.446924f
C39 VN.t2 VSUBS 0.44685f
C40 VN.n1 VSUBS 1.07116f
C41 VTAIL.n0 VSUBS 0.019311f
C42 VTAIL.n1 VSUBS 0.018653f
C43 VTAIL.n2 VSUBS 0.010023f
C44 VTAIL.n3 VSUBS 0.023692f
C45 VTAIL.n4 VSUBS 0.010613f
C46 VTAIL.n5 VSUBS 0.07099f
C47 VTAIL.t0 VSUBS 0.05178f
C48 VTAIL.n6 VSUBS 0.017769f
C49 VTAIL.n7 VSUBS 0.014902f
C50 VTAIL.n8 VSUBS 0.010023f
C51 VTAIL.n9 VSUBS 0.241895f
C52 VTAIL.n10 VSUBS 0.018653f
C53 VTAIL.n11 VSUBS 0.010023f
C54 VTAIL.n12 VSUBS 0.010613f
C55 VTAIL.n13 VSUBS 0.023692f
C56 VTAIL.n14 VSUBS 0.053319f
C57 VTAIL.n15 VSUBS 0.010613f
C58 VTAIL.n16 VSUBS 0.010023f
C59 VTAIL.n17 VSUBS 0.042606f
C60 VTAIL.n18 VSUBS 0.026618f
C61 VTAIL.n19 VSUBS 0.076137f
C62 VTAIL.n20 VSUBS 0.019311f
C63 VTAIL.n21 VSUBS 0.018653f
C64 VTAIL.n22 VSUBS 0.010023f
C65 VTAIL.n23 VSUBS 0.023692f
C66 VTAIL.n24 VSUBS 0.010613f
C67 VTAIL.n25 VSUBS 0.07099f
C68 VTAIL.t5 VSUBS 0.05178f
C69 VTAIL.n26 VSUBS 0.017769f
C70 VTAIL.n27 VSUBS 0.014902f
C71 VTAIL.n28 VSUBS 0.010023f
C72 VTAIL.n29 VSUBS 0.241895f
C73 VTAIL.n30 VSUBS 0.018653f
C74 VTAIL.n31 VSUBS 0.010023f
C75 VTAIL.n32 VSUBS 0.010613f
C76 VTAIL.n33 VSUBS 0.023692f
C77 VTAIL.n34 VSUBS 0.053319f
C78 VTAIL.n35 VSUBS 0.010613f
C79 VTAIL.n36 VSUBS 0.010023f
C80 VTAIL.n37 VSUBS 0.042606f
C81 VTAIL.n38 VSUBS 0.026618f
C82 VTAIL.n39 VSUBS 0.101396f
C83 VTAIL.n40 VSUBS 0.019311f
C84 VTAIL.n41 VSUBS 0.018653f
C85 VTAIL.n42 VSUBS 0.010023f
C86 VTAIL.n43 VSUBS 0.023692f
C87 VTAIL.n44 VSUBS 0.010613f
C88 VTAIL.n45 VSUBS 0.07099f
C89 VTAIL.t7 VSUBS 0.05178f
C90 VTAIL.n46 VSUBS 0.017769f
C91 VTAIL.n47 VSUBS 0.014902f
C92 VTAIL.n48 VSUBS 0.010023f
C93 VTAIL.n49 VSUBS 0.241895f
C94 VTAIL.n50 VSUBS 0.018653f
C95 VTAIL.n51 VSUBS 0.010023f
C96 VTAIL.n52 VSUBS 0.010613f
C97 VTAIL.n53 VSUBS 0.023692f
C98 VTAIL.n54 VSUBS 0.053319f
C99 VTAIL.n55 VSUBS 0.010613f
C100 VTAIL.n56 VSUBS 0.010023f
C101 VTAIL.n57 VSUBS 0.042606f
C102 VTAIL.n58 VSUBS 0.026618f
C103 VTAIL.n59 VSUBS 0.581982f
C104 VTAIL.n60 VSUBS 0.019311f
C105 VTAIL.n61 VSUBS 0.018653f
C106 VTAIL.n62 VSUBS 0.010023f
C107 VTAIL.n63 VSUBS 0.023692f
C108 VTAIL.n64 VSUBS 0.010613f
C109 VTAIL.n65 VSUBS 0.07099f
C110 VTAIL.t1 VSUBS 0.05178f
C111 VTAIL.n66 VSUBS 0.017769f
C112 VTAIL.n67 VSUBS 0.014902f
C113 VTAIL.n68 VSUBS 0.010023f
C114 VTAIL.n69 VSUBS 0.241895f
C115 VTAIL.n70 VSUBS 0.018653f
C116 VTAIL.n71 VSUBS 0.010023f
C117 VTAIL.n72 VSUBS 0.010613f
C118 VTAIL.n73 VSUBS 0.023692f
C119 VTAIL.n74 VSUBS 0.053319f
C120 VTAIL.n75 VSUBS 0.010613f
C121 VTAIL.n76 VSUBS 0.010023f
C122 VTAIL.n77 VSUBS 0.042606f
C123 VTAIL.n78 VSUBS 0.026618f
C124 VTAIL.n79 VSUBS 0.581982f
C125 VTAIL.n80 VSUBS 0.019311f
C126 VTAIL.n81 VSUBS 0.018653f
C127 VTAIL.n82 VSUBS 0.010023f
C128 VTAIL.n83 VSUBS 0.023692f
C129 VTAIL.n84 VSUBS 0.010613f
C130 VTAIL.n85 VSUBS 0.07099f
C131 VTAIL.t3 VSUBS 0.05178f
C132 VTAIL.n86 VSUBS 0.017769f
C133 VTAIL.n87 VSUBS 0.014902f
C134 VTAIL.n88 VSUBS 0.010023f
C135 VTAIL.n89 VSUBS 0.241895f
C136 VTAIL.n90 VSUBS 0.018653f
C137 VTAIL.n91 VSUBS 0.010023f
C138 VTAIL.n92 VSUBS 0.010613f
C139 VTAIL.n93 VSUBS 0.023692f
C140 VTAIL.n94 VSUBS 0.053319f
C141 VTAIL.n95 VSUBS 0.010613f
C142 VTAIL.n96 VSUBS 0.010023f
C143 VTAIL.n97 VSUBS 0.042606f
C144 VTAIL.n98 VSUBS 0.026618f
C145 VTAIL.n99 VSUBS 0.101396f
C146 VTAIL.n100 VSUBS 0.019311f
C147 VTAIL.n101 VSUBS 0.018653f
C148 VTAIL.n102 VSUBS 0.010023f
C149 VTAIL.n103 VSUBS 0.023692f
C150 VTAIL.n104 VSUBS 0.010613f
C151 VTAIL.n105 VSUBS 0.07099f
C152 VTAIL.t4 VSUBS 0.05178f
C153 VTAIL.n106 VSUBS 0.017769f
C154 VTAIL.n107 VSUBS 0.014902f
C155 VTAIL.n108 VSUBS 0.010023f
C156 VTAIL.n109 VSUBS 0.241895f
C157 VTAIL.n110 VSUBS 0.018653f
C158 VTAIL.n111 VSUBS 0.010023f
C159 VTAIL.n112 VSUBS 0.010613f
C160 VTAIL.n113 VSUBS 0.023692f
C161 VTAIL.n114 VSUBS 0.053319f
C162 VTAIL.n115 VSUBS 0.010613f
C163 VTAIL.n116 VSUBS 0.010023f
C164 VTAIL.n117 VSUBS 0.042606f
C165 VTAIL.n118 VSUBS 0.026618f
C166 VTAIL.n119 VSUBS 0.101396f
C167 VTAIL.n120 VSUBS 0.019311f
C168 VTAIL.n121 VSUBS 0.018653f
C169 VTAIL.n122 VSUBS 0.010023f
C170 VTAIL.n123 VSUBS 0.023692f
C171 VTAIL.n124 VSUBS 0.010613f
C172 VTAIL.n125 VSUBS 0.07099f
C173 VTAIL.t6 VSUBS 0.05178f
C174 VTAIL.n126 VSUBS 0.017769f
C175 VTAIL.n127 VSUBS 0.014902f
C176 VTAIL.n128 VSUBS 0.010023f
C177 VTAIL.n129 VSUBS 0.241895f
C178 VTAIL.n130 VSUBS 0.018653f
C179 VTAIL.n131 VSUBS 0.010023f
C180 VTAIL.n132 VSUBS 0.010613f
C181 VTAIL.n133 VSUBS 0.023692f
C182 VTAIL.n134 VSUBS 0.053319f
C183 VTAIL.n135 VSUBS 0.010613f
C184 VTAIL.n136 VSUBS 0.010023f
C185 VTAIL.n137 VSUBS 0.042606f
C186 VTAIL.n138 VSUBS 0.026618f
C187 VTAIL.n139 VSUBS 0.581982f
C188 VTAIL.n140 VSUBS 0.019311f
C189 VTAIL.n141 VSUBS 0.018653f
C190 VTAIL.n142 VSUBS 0.010023f
C191 VTAIL.n143 VSUBS 0.023692f
C192 VTAIL.n144 VSUBS 0.010613f
C193 VTAIL.n145 VSUBS 0.07099f
C194 VTAIL.t2 VSUBS 0.05178f
C195 VTAIL.n146 VSUBS 0.017769f
C196 VTAIL.n147 VSUBS 0.014902f
C197 VTAIL.n148 VSUBS 0.010023f
C198 VTAIL.n149 VSUBS 0.241895f
C199 VTAIL.n150 VSUBS 0.018653f
C200 VTAIL.n151 VSUBS 0.010023f
C201 VTAIL.n152 VSUBS 0.010613f
C202 VTAIL.n153 VSUBS 0.023692f
C203 VTAIL.n154 VSUBS 0.053319f
C204 VTAIL.n155 VSUBS 0.010613f
C205 VTAIL.n156 VSUBS 0.010023f
C206 VTAIL.n157 VSUBS 0.042606f
C207 VTAIL.n158 VSUBS 0.026618f
C208 VTAIL.n159 VSUBS 0.549728f
C209 VDD1.t1 VSUBS 0.056853f
C210 VDD1.t0 VSUBS 0.056853f
C211 VDD1.n0 VSUBS 0.327314f
C212 VDD1.t3 VSUBS 0.056853f
C213 VDD1.t2 VSUBS 0.056853f
C214 VDD1.n1 VSUBS 0.511543f
C215 VP.n0 VSUBS 0.050202f
C216 VP.t1 VSUBS 0.468061f
C217 VP.t3 VSUBS 0.468138f
C218 VP.n1 VSUBS 1.10312f
C219 VP.n2 VSUBS 2.39277f
C220 VP.t0 VSUBS 0.44224f
C221 VP.n3 VSUBS 0.229782f
C222 VP.n4 VSUBS 0.011392f
C223 VP.t2 VSUBS 0.44224f
C224 VP.n5 VSUBS 0.229782f
C225 VP.n6 VSUBS 0.038904f
C226 B.n0 VSUBS 0.004741f
C227 B.n1 VSUBS 0.004741f
C228 B.n2 VSUBS 0.007497f
C229 B.n3 VSUBS 0.007497f
C230 B.n4 VSUBS 0.007497f
C231 B.n5 VSUBS 0.007497f
C232 B.n6 VSUBS 0.007497f
C233 B.n7 VSUBS 0.007497f
C234 B.n8 VSUBS 0.007497f
C235 B.n9 VSUBS 0.007497f
C236 B.n10 VSUBS 0.007497f
C237 B.n11 VSUBS 0.017047f
C238 B.n12 VSUBS 0.007497f
C239 B.n13 VSUBS 0.007497f
C240 B.n14 VSUBS 0.007497f
C241 B.n15 VSUBS 0.007497f
C242 B.n16 VSUBS 0.007497f
C243 B.n17 VSUBS 0.007497f
C244 B.n18 VSUBS 0.007497f
C245 B.n19 VSUBS 0.007497f
C246 B.t11 VSUBS 0.058882f
C247 B.t10 VSUBS 0.067482f
C248 B.t9 VSUBS 0.144249f
C249 B.n20 VSUBS 0.124439f
C250 B.n21 VSUBS 0.112025f
C251 B.n22 VSUBS 0.01737f
C252 B.n23 VSUBS 0.007497f
C253 B.n24 VSUBS 0.007497f
C254 B.n25 VSUBS 0.007497f
C255 B.n26 VSUBS 0.007497f
C256 B.n27 VSUBS 0.007497f
C257 B.t5 VSUBS 0.058883f
C258 B.t4 VSUBS 0.067483f
C259 B.t3 VSUBS 0.144249f
C260 B.n28 VSUBS 0.124438f
C261 B.n29 VSUBS 0.112024f
C262 B.n30 VSUBS 0.007497f
C263 B.n31 VSUBS 0.007497f
C264 B.n32 VSUBS 0.007497f
C265 B.n33 VSUBS 0.007497f
C266 B.n34 VSUBS 0.007497f
C267 B.n35 VSUBS 0.007497f
C268 B.n36 VSUBS 0.007497f
C269 B.n37 VSUBS 0.007497f
C270 B.n38 VSUBS 0.017f
C271 B.n39 VSUBS 0.007497f
C272 B.n40 VSUBS 0.007497f
C273 B.n41 VSUBS 0.007497f
C274 B.n42 VSUBS 0.007497f
C275 B.n43 VSUBS 0.007497f
C276 B.n44 VSUBS 0.007497f
C277 B.n45 VSUBS 0.007497f
C278 B.n46 VSUBS 0.007497f
C279 B.n47 VSUBS 0.007497f
C280 B.n48 VSUBS 0.007497f
C281 B.n49 VSUBS 0.007497f
C282 B.n50 VSUBS 0.007497f
C283 B.n51 VSUBS 0.007497f
C284 B.n52 VSUBS 0.007497f
C285 B.n53 VSUBS 0.007497f
C286 B.n54 VSUBS 0.007497f
C287 B.n55 VSUBS 0.007497f
C288 B.n56 VSUBS 0.016029f
C289 B.n57 VSUBS 0.007497f
C290 B.n58 VSUBS 0.007497f
C291 B.n59 VSUBS 0.007497f
C292 B.n60 VSUBS 0.007497f
C293 B.n61 VSUBS 0.007497f
C294 B.n62 VSUBS 0.007497f
C295 B.n63 VSUBS 0.007497f
C296 B.n64 VSUBS 0.007497f
C297 B.n65 VSUBS 0.007497f
C298 B.t7 VSUBS 0.058883f
C299 B.t8 VSUBS 0.067483f
C300 B.t6 VSUBS 0.144249f
C301 B.n66 VSUBS 0.124438f
C302 B.n67 VSUBS 0.112024f
C303 B.n68 VSUBS 0.007497f
C304 B.n69 VSUBS 0.007497f
C305 B.n70 VSUBS 0.007497f
C306 B.n71 VSUBS 0.007497f
C307 B.t1 VSUBS 0.058882f
C308 B.t2 VSUBS 0.067482f
C309 B.t0 VSUBS 0.144249f
C310 B.n72 VSUBS 0.124439f
C311 B.n73 VSUBS 0.112025f
C312 B.n74 VSUBS 0.01737f
C313 B.n75 VSUBS 0.007497f
C314 B.n76 VSUBS 0.007497f
C315 B.n77 VSUBS 0.007497f
C316 B.n78 VSUBS 0.007497f
C317 B.n79 VSUBS 0.007497f
C318 B.n80 VSUBS 0.007497f
C319 B.n81 VSUBS 0.007497f
C320 B.n82 VSUBS 0.007497f
C321 B.n83 VSUBS 0.017047f
C322 B.n84 VSUBS 0.007497f
C323 B.n85 VSUBS 0.007497f
C324 B.n86 VSUBS 0.007497f
C325 B.n87 VSUBS 0.007497f
C326 B.n88 VSUBS 0.007497f
C327 B.n89 VSUBS 0.007497f
C328 B.n90 VSUBS 0.007497f
C329 B.n91 VSUBS 0.007497f
C330 B.n92 VSUBS 0.007497f
C331 B.n93 VSUBS 0.007497f
C332 B.n94 VSUBS 0.007497f
C333 B.n95 VSUBS 0.007497f
C334 B.n96 VSUBS 0.007497f
C335 B.n97 VSUBS 0.007497f
C336 B.n98 VSUBS 0.007497f
C337 B.n99 VSUBS 0.007497f
C338 B.n100 VSUBS 0.007497f
C339 B.n101 VSUBS 0.007497f
C340 B.n102 VSUBS 0.007497f
C341 B.n103 VSUBS 0.007497f
C342 B.n104 VSUBS 0.007497f
C343 B.n105 VSUBS 0.007497f
C344 B.n106 VSUBS 0.007497f
C345 B.n107 VSUBS 0.007497f
C346 B.n108 VSUBS 0.007497f
C347 B.n109 VSUBS 0.007497f
C348 B.n110 VSUBS 0.007497f
C349 B.n111 VSUBS 0.007497f
C350 B.n112 VSUBS 0.007497f
C351 B.n113 VSUBS 0.007497f
C352 B.n114 VSUBS 0.007497f
C353 B.n115 VSUBS 0.007497f
C354 B.n116 VSUBS 0.016029f
C355 B.n117 VSUBS 0.016029f
C356 B.n118 VSUBS 0.017047f
C357 B.n119 VSUBS 0.007497f
C358 B.n120 VSUBS 0.007497f
C359 B.n121 VSUBS 0.007497f
C360 B.n122 VSUBS 0.007497f
C361 B.n123 VSUBS 0.007497f
C362 B.n124 VSUBS 0.007497f
C363 B.n125 VSUBS 0.007497f
C364 B.n126 VSUBS 0.007497f
C365 B.n127 VSUBS 0.007497f
C366 B.n128 VSUBS 0.007497f
C367 B.n129 VSUBS 0.007497f
C368 B.n130 VSUBS 0.007497f
C369 B.n131 VSUBS 0.007497f
C370 B.n132 VSUBS 0.007497f
C371 B.n133 VSUBS 0.007497f
C372 B.n134 VSUBS 0.007497f
C373 B.n135 VSUBS 0.007497f
C374 B.n136 VSUBS 0.007497f
C375 B.n137 VSUBS 0.007497f
C376 B.n138 VSUBS 0.007497f
C377 B.n139 VSUBS 0.007497f
C378 B.n140 VSUBS 0.007497f
C379 B.n141 VSUBS 0.007497f
C380 B.n142 VSUBS 0.007497f
C381 B.n143 VSUBS 0.005182f
C382 B.n144 VSUBS 0.007497f
C383 B.n145 VSUBS 0.007497f
C384 B.n146 VSUBS 0.006064f
C385 B.n147 VSUBS 0.007497f
C386 B.n148 VSUBS 0.007497f
C387 B.n149 VSUBS 0.007497f
C388 B.n150 VSUBS 0.007497f
C389 B.n151 VSUBS 0.007497f
C390 B.n152 VSUBS 0.007497f
C391 B.n153 VSUBS 0.007497f
C392 B.n154 VSUBS 0.007497f
C393 B.n155 VSUBS 0.007497f
C394 B.n156 VSUBS 0.007497f
C395 B.n157 VSUBS 0.007497f
C396 B.n158 VSUBS 0.006064f
C397 B.n159 VSUBS 0.01737f
C398 B.n160 VSUBS 0.005182f
C399 B.n161 VSUBS 0.007497f
C400 B.n162 VSUBS 0.007497f
C401 B.n163 VSUBS 0.007497f
C402 B.n164 VSUBS 0.007497f
C403 B.n165 VSUBS 0.007497f
C404 B.n166 VSUBS 0.007497f
C405 B.n167 VSUBS 0.007497f
C406 B.n168 VSUBS 0.007497f
C407 B.n169 VSUBS 0.007497f
C408 B.n170 VSUBS 0.007497f
C409 B.n171 VSUBS 0.007497f
C410 B.n172 VSUBS 0.007497f
C411 B.n173 VSUBS 0.007497f
C412 B.n174 VSUBS 0.007497f
C413 B.n175 VSUBS 0.007497f
C414 B.n176 VSUBS 0.007497f
C415 B.n177 VSUBS 0.007497f
C416 B.n178 VSUBS 0.007497f
C417 B.n179 VSUBS 0.007497f
C418 B.n180 VSUBS 0.007497f
C419 B.n181 VSUBS 0.007497f
C420 B.n182 VSUBS 0.007497f
C421 B.n183 VSUBS 0.007497f
C422 B.n184 VSUBS 0.007497f
C423 B.n185 VSUBS 0.017047f
C424 B.n186 VSUBS 0.017047f
C425 B.n187 VSUBS 0.016029f
C426 B.n188 VSUBS 0.007497f
C427 B.n189 VSUBS 0.007497f
C428 B.n190 VSUBS 0.007497f
C429 B.n191 VSUBS 0.007497f
C430 B.n192 VSUBS 0.007497f
C431 B.n193 VSUBS 0.007497f
C432 B.n194 VSUBS 0.007497f
C433 B.n195 VSUBS 0.007497f
C434 B.n196 VSUBS 0.007497f
C435 B.n197 VSUBS 0.007497f
C436 B.n198 VSUBS 0.007497f
C437 B.n199 VSUBS 0.007497f
C438 B.n200 VSUBS 0.007497f
C439 B.n201 VSUBS 0.007497f
C440 B.n202 VSUBS 0.007497f
C441 B.n203 VSUBS 0.007497f
C442 B.n204 VSUBS 0.007497f
C443 B.n205 VSUBS 0.007497f
C444 B.n206 VSUBS 0.007497f
C445 B.n207 VSUBS 0.007497f
C446 B.n208 VSUBS 0.007497f
C447 B.n209 VSUBS 0.007497f
C448 B.n210 VSUBS 0.007497f
C449 B.n211 VSUBS 0.007497f
C450 B.n212 VSUBS 0.007497f
C451 B.n213 VSUBS 0.007497f
C452 B.n214 VSUBS 0.007497f
C453 B.n215 VSUBS 0.007497f
C454 B.n216 VSUBS 0.007497f
C455 B.n217 VSUBS 0.007497f
C456 B.n218 VSUBS 0.007497f
C457 B.n219 VSUBS 0.007497f
C458 B.n220 VSUBS 0.007497f
C459 B.n221 VSUBS 0.007497f
C460 B.n222 VSUBS 0.007497f
C461 B.n223 VSUBS 0.007497f
C462 B.n224 VSUBS 0.007497f
C463 B.n225 VSUBS 0.007497f
C464 B.n226 VSUBS 0.007497f
C465 B.n227 VSUBS 0.007497f
C466 B.n228 VSUBS 0.007497f
C467 B.n229 VSUBS 0.007497f
C468 B.n230 VSUBS 0.007497f
C469 B.n231 VSUBS 0.007497f
C470 B.n232 VSUBS 0.007497f
C471 B.n233 VSUBS 0.007497f
C472 B.n234 VSUBS 0.007497f
C473 B.n235 VSUBS 0.007497f
C474 B.n236 VSUBS 0.007497f
C475 B.n237 VSUBS 0.007497f
C476 B.n238 VSUBS 0.007497f
C477 B.n239 VSUBS 0.007497f
C478 B.n240 VSUBS 0.007497f
C479 B.n241 VSUBS 0.016029f
C480 B.n242 VSUBS 0.017047f
C481 B.n243 VSUBS 0.016077f
C482 B.n244 VSUBS 0.007497f
C483 B.n245 VSUBS 0.007497f
C484 B.n246 VSUBS 0.007497f
C485 B.n247 VSUBS 0.007497f
C486 B.n248 VSUBS 0.007497f
C487 B.n249 VSUBS 0.007497f
C488 B.n250 VSUBS 0.007497f
C489 B.n251 VSUBS 0.007497f
C490 B.n252 VSUBS 0.007497f
C491 B.n253 VSUBS 0.007497f
C492 B.n254 VSUBS 0.007497f
C493 B.n255 VSUBS 0.007497f
C494 B.n256 VSUBS 0.007497f
C495 B.n257 VSUBS 0.007497f
C496 B.n258 VSUBS 0.007497f
C497 B.n259 VSUBS 0.007497f
C498 B.n260 VSUBS 0.007497f
C499 B.n261 VSUBS 0.007497f
C500 B.n262 VSUBS 0.007497f
C501 B.n263 VSUBS 0.007497f
C502 B.n264 VSUBS 0.007497f
C503 B.n265 VSUBS 0.007497f
C504 B.n266 VSUBS 0.007497f
C505 B.n267 VSUBS 0.007497f
C506 B.n268 VSUBS 0.005182f
C507 B.n269 VSUBS 0.01737f
C508 B.n270 VSUBS 0.006064f
C509 B.n271 VSUBS 0.007497f
C510 B.n272 VSUBS 0.007497f
C511 B.n273 VSUBS 0.007497f
C512 B.n274 VSUBS 0.007497f
C513 B.n275 VSUBS 0.007497f
C514 B.n276 VSUBS 0.007497f
C515 B.n277 VSUBS 0.007497f
C516 B.n278 VSUBS 0.007497f
C517 B.n279 VSUBS 0.007497f
C518 B.n280 VSUBS 0.007497f
C519 B.n281 VSUBS 0.007497f
C520 B.n282 VSUBS 0.006064f
C521 B.n283 VSUBS 0.007497f
C522 B.n284 VSUBS 0.007497f
C523 B.n285 VSUBS 0.005182f
C524 B.n286 VSUBS 0.007497f
C525 B.n287 VSUBS 0.007497f
C526 B.n288 VSUBS 0.007497f
C527 B.n289 VSUBS 0.007497f
C528 B.n290 VSUBS 0.007497f
C529 B.n291 VSUBS 0.007497f
C530 B.n292 VSUBS 0.007497f
C531 B.n293 VSUBS 0.007497f
C532 B.n294 VSUBS 0.007497f
C533 B.n295 VSUBS 0.007497f
C534 B.n296 VSUBS 0.007497f
C535 B.n297 VSUBS 0.007497f
C536 B.n298 VSUBS 0.007497f
C537 B.n299 VSUBS 0.007497f
C538 B.n300 VSUBS 0.007497f
C539 B.n301 VSUBS 0.007497f
C540 B.n302 VSUBS 0.007497f
C541 B.n303 VSUBS 0.007497f
C542 B.n304 VSUBS 0.007497f
C543 B.n305 VSUBS 0.007497f
C544 B.n306 VSUBS 0.007497f
C545 B.n307 VSUBS 0.007497f
C546 B.n308 VSUBS 0.007497f
C547 B.n309 VSUBS 0.007497f
C548 B.n310 VSUBS 0.017047f
C549 B.n311 VSUBS 0.016029f
C550 B.n312 VSUBS 0.016029f
C551 B.n313 VSUBS 0.007497f
C552 B.n314 VSUBS 0.007497f
C553 B.n315 VSUBS 0.007497f
C554 B.n316 VSUBS 0.007497f
C555 B.n317 VSUBS 0.007497f
C556 B.n318 VSUBS 0.007497f
C557 B.n319 VSUBS 0.007497f
C558 B.n320 VSUBS 0.007497f
C559 B.n321 VSUBS 0.007497f
C560 B.n322 VSUBS 0.007497f
C561 B.n323 VSUBS 0.007497f
C562 B.n324 VSUBS 0.007497f
C563 B.n325 VSUBS 0.007497f
C564 B.n326 VSUBS 0.007497f
C565 B.n327 VSUBS 0.007497f
C566 B.n328 VSUBS 0.007497f
C567 B.n329 VSUBS 0.007497f
C568 B.n330 VSUBS 0.007497f
C569 B.n331 VSUBS 0.007497f
C570 B.n332 VSUBS 0.007497f
C571 B.n333 VSUBS 0.007497f
C572 B.n334 VSUBS 0.007497f
C573 B.n335 VSUBS 0.007497f
C574 B.n336 VSUBS 0.007497f
C575 B.n337 VSUBS 0.007497f
C576 B.n338 VSUBS 0.007497f
C577 B.n339 VSUBS 0.016976f
.ends

