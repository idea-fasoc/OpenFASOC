* NGSPICE file created from diff_pair_sample_0173.ext - technology: sky130A

.subckt diff_pair_sample_0173 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=2.7885 pd=15.08 as=0 ps=0 w=7.15 l=2.04
X1 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=2.7885 pd=15.08 as=0 ps=0 w=7.15 l=2.04
X2 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7885 pd=15.08 as=0 ps=0 w=7.15 l=2.04
X3 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7885 pd=15.08 as=2.7885 ps=15.08 w=7.15 l=2.04
X4 VDD2.t0 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7885 pd=15.08 as=2.7885 ps=15.08 w=7.15 l=2.04
X5 VDD1.t1 VP.t0 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7885 pd=15.08 as=2.7885 ps=15.08 w=7.15 l=2.04
X6 VDD1.t0 VP.t1 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7885 pd=15.08 as=2.7885 ps=15.08 w=7.15 l=2.04
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7885 pd=15.08 as=0 ps=0 w=7.15 l=2.04
R0 B.n383 B.n382 585
R1 B.n385 B.n80 585
R2 B.n388 B.n387 585
R3 B.n389 B.n79 585
R4 B.n391 B.n390 585
R5 B.n393 B.n78 585
R6 B.n396 B.n395 585
R7 B.n397 B.n77 585
R8 B.n399 B.n398 585
R9 B.n401 B.n76 585
R10 B.n404 B.n403 585
R11 B.n405 B.n75 585
R12 B.n407 B.n406 585
R13 B.n409 B.n74 585
R14 B.n412 B.n411 585
R15 B.n413 B.n73 585
R16 B.n415 B.n414 585
R17 B.n417 B.n72 585
R18 B.n420 B.n419 585
R19 B.n421 B.n71 585
R20 B.n423 B.n422 585
R21 B.n425 B.n70 585
R22 B.n428 B.n427 585
R23 B.n429 B.n69 585
R24 B.n431 B.n430 585
R25 B.n433 B.n68 585
R26 B.n436 B.n435 585
R27 B.n438 B.n65 585
R28 B.n440 B.n439 585
R29 B.n442 B.n64 585
R30 B.n445 B.n444 585
R31 B.n446 B.n63 585
R32 B.n448 B.n447 585
R33 B.n450 B.n62 585
R34 B.n453 B.n452 585
R35 B.n454 B.n58 585
R36 B.n456 B.n455 585
R37 B.n458 B.n57 585
R38 B.n461 B.n460 585
R39 B.n462 B.n56 585
R40 B.n464 B.n463 585
R41 B.n466 B.n55 585
R42 B.n469 B.n468 585
R43 B.n470 B.n54 585
R44 B.n472 B.n471 585
R45 B.n474 B.n53 585
R46 B.n477 B.n476 585
R47 B.n478 B.n52 585
R48 B.n480 B.n479 585
R49 B.n482 B.n51 585
R50 B.n485 B.n484 585
R51 B.n486 B.n50 585
R52 B.n488 B.n487 585
R53 B.n490 B.n49 585
R54 B.n493 B.n492 585
R55 B.n494 B.n48 585
R56 B.n496 B.n495 585
R57 B.n498 B.n47 585
R58 B.n501 B.n500 585
R59 B.n502 B.n46 585
R60 B.n504 B.n503 585
R61 B.n506 B.n45 585
R62 B.n509 B.n508 585
R63 B.n510 B.n44 585
R64 B.n381 B.n42 585
R65 B.n513 B.n42 585
R66 B.n380 B.n41 585
R67 B.n514 B.n41 585
R68 B.n379 B.n40 585
R69 B.n515 B.n40 585
R70 B.n378 B.n377 585
R71 B.n377 B.n36 585
R72 B.n376 B.n35 585
R73 B.n521 B.n35 585
R74 B.n375 B.n34 585
R75 B.n522 B.n34 585
R76 B.n374 B.n33 585
R77 B.n523 B.n33 585
R78 B.n373 B.n372 585
R79 B.n372 B.n29 585
R80 B.n371 B.n28 585
R81 B.n529 B.n28 585
R82 B.n370 B.n27 585
R83 B.n530 B.n27 585
R84 B.n369 B.n26 585
R85 B.n531 B.n26 585
R86 B.n368 B.n367 585
R87 B.n367 B.n22 585
R88 B.n366 B.n21 585
R89 B.n537 B.n21 585
R90 B.n365 B.n20 585
R91 B.n538 B.n20 585
R92 B.n364 B.n19 585
R93 B.n539 B.n19 585
R94 B.n363 B.n362 585
R95 B.n362 B.n15 585
R96 B.n361 B.n14 585
R97 B.n545 B.n14 585
R98 B.n360 B.n13 585
R99 B.n546 B.n13 585
R100 B.n359 B.n12 585
R101 B.n547 B.n12 585
R102 B.n358 B.n357 585
R103 B.n357 B.n8 585
R104 B.n356 B.n7 585
R105 B.n553 B.n7 585
R106 B.n355 B.n6 585
R107 B.n554 B.n6 585
R108 B.n354 B.n5 585
R109 B.n555 B.n5 585
R110 B.n353 B.n352 585
R111 B.n352 B.n4 585
R112 B.n351 B.n81 585
R113 B.n351 B.n350 585
R114 B.n341 B.n82 585
R115 B.n83 B.n82 585
R116 B.n343 B.n342 585
R117 B.n344 B.n343 585
R118 B.n340 B.n88 585
R119 B.n88 B.n87 585
R120 B.n339 B.n338 585
R121 B.n338 B.n337 585
R122 B.n90 B.n89 585
R123 B.n91 B.n90 585
R124 B.n330 B.n329 585
R125 B.n331 B.n330 585
R126 B.n328 B.n96 585
R127 B.n96 B.n95 585
R128 B.n327 B.n326 585
R129 B.n326 B.n325 585
R130 B.n98 B.n97 585
R131 B.n99 B.n98 585
R132 B.n318 B.n317 585
R133 B.n319 B.n318 585
R134 B.n316 B.n104 585
R135 B.n104 B.n103 585
R136 B.n315 B.n314 585
R137 B.n314 B.n313 585
R138 B.n106 B.n105 585
R139 B.n107 B.n106 585
R140 B.n306 B.n305 585
R141 B.n307 B.n306 585
R142 B.n304 B.n112 585
R143 B.n112 B.n111 585
R144 B.n303 B.n302 585
R145 B.n302 B.n301 585
R146 B.n114 B.n113 585
R147 B.n115 B.n114 585
R148 B.n294 B.n293 585
R149 B.n295 B.n294 585
R150 B.n292 B.n120 585
R151 B.n120 B.n119 585
R152 B.n291 B.n290 585
R153 B.n290 B.n289 585
R154 B.n286 B.n124 585
R155 B.n285 B.n284 585
R156 B.n282 B.n125 585
R157 B.n282 B.n123 585
R158 B.n281 B.n280 585
R159 B.n279 B.n278 585
R160 B.n277 B.n127 585
R161 B.n275 B.n274 585
R162 B.n273 B.n128 585
R163 B.n272 B.n271 585
R164 B.n269 B.n129 585
R165 B.n267 B.n266 585
R166 B.n265 B.n130 585
R167 B.n264 B.n263 585
R168 B.n261 B.n131 585
R169 B.n259 B.n258 585
R170 B.n257 B.n132 585
R171 B.n256 B.n255 585
R172 B.n253 B.n133 585
R173 B.n251 B.n250 585
R174 B.n249 B.n134 585
R175 B.n248 B.n247 585
R176 B.n245 B.n135 585
R177 B.n243 B.n242 585
R178 B.n241 B.n136 585
R179 B.n240 B.n239 585
R180 B.n237 B.n137 585
R181 B.n235 B.n234 585
R182 B.n232 B.n138 585
R183 B.n231 B.n230 585
R184 B.n228 B.n141 585
R185 B.n226 B.n225 585
R186 B.n224 B.n142 585
R187 B.n223 B.n222 585
R188 B.n220 B.n143 585
R189 B.n218 B.n217 585
R190 B.n216 B.n144 585
R191 B.n215 B.n214 585
R192 B.n212 B.n211 585
R193 B.n210 B.n209 585
R194 B.n208 B.n149 585
R195 B.n206 B.n205 585
R196 B.n204 B.n150 585
R197 B.n203 B.n202 585
R198 B.n200 B.n151 585
R199 B.n198 B.n197 585
R200 B.n196 B.n152 585
R201 B.n195 B.n194 585
R202 B.n192 B.n153 585
R203 B.n190 B.n189 585
R204 B.n188 B.n154 585
R205 B.n187 B.n186 585
R206 B.n184 B.n155 585
R207 B.n182 B.n181 585
R208 B.n180 B.n156 585
R209 B.n179 B.n178 585
R210 B.n176 B.n157 585
R211 B.n174 B.n173 585
R212 B.n172 B.n158 585
R213 B.n171 B.n170 585
R214 B.n168 B.n159 585
R215 B.n166 B.n165 585
R216 B.n164 B.n160 585
R217 B.n163 B.n162 585
R218 B.n122 B.n121 585
R219 B.n123 B.n122 585
R220 B.n288 B.n287 585
R221 B.n289 B.n288 585
R222 B.n118 B.n117 585
R223 B.n119 B.n118 585
R224 B.n297 B.n296 585
R225 B.n296 B.n295 585
R226 B.n298 B.n116 585
R227 B.n116 B.n115 585
R228 B.n300 B.n299 585
R229 B.n301 B.n300 585
R230 B.n110 B.n109 585
R231 B.n111 B.n110 585
R232 B.n309 B.n308 585
R233 B.n308 B.n307 585
R234 B.n310 B.n108 585
R235 B.n108 B.n107 585
R236 B.n312 B.n311 585
R237 B.n313 B.n312 585
R238 B.n102 B.n101 585
R239 B.n103 B.n102 585
R240 B.n321 B.n320 585
R241 B.n320 B.n319 585
R242 B.n322 B.n100 585
R243 B.n100 B.n99 585
R244 B.n324 B.n323 585
R245 B.n325 B.n324 585
R246 B.n94 B.n93 585
R247 B.n95 B.n94 585
R248 B.n333 B.n332 585
R249 B.n332 B.n331 585
R250 B.n334 B.n92 585
R251 B.n92 B.n91 585
R252 B.n336 B.n335 585
R253 B.n337 B.n336 585
R254 B.n86 B.n85 585
R255 B.n87 B.n86 585
R256 B.n346 B.n345 585
R257 B.n345 B.n344 585
R258 B.n347 B.n84 585
R259 B.n84 B.n83 585
R260 B.n349 B.n348 585
R261 B.n350 B.n349 585
R262 B.n2 B.n0 585
R263 B.n4 B.n2 585
R264 B.n3 B.n1 585
R265 B.n554 B.n3 585
R266 B.n552 B.n551 585
R267 B.n553 B.n552 585
R268 B.n550 B.n9 585
R269 B.n9 B.n8 585
R270 B.n549 B.n548 585
R271 B.n548 B.n547 585
R272 B.n11 B.n10 585
R273 B.n546 B.n11 585
R274 B.n544 B.n543 585
R275 B.n545 B.n544 585
R276 B.n542 B.n16 585
R277 B.n16 B.n15 585
R278 B.n541 B.n540 585
R279 B.n540 B.n539 585
R280 B.n18 B.n17 585
R281 B.n538 B.n18 585
R282 B.n536 B.n535 585
R283 B.n537 B.n536 585
R284 B.n534 B.n23 585
R285 B.n23 B.n22 585
R286 B.n533 B.n532 585
R287 B.n532 B.n531 585
R288 B.n25 B.n24 585
R289 B.n530 B.n25 585
R290 B.n528 B.n527 585
R291 B.n529 B.n528 585
R292 B.n526 B.n30 585
R293 B.n30 B.n29 585
R294 B.n525 B.n524 585
R295 B.n524 B.n523 585
R296 B.n32 B.n31 585
R297 B.n522 B.n32 585
R298 B.n520 B.n519 585
R299 B.n521 B.n520 585
R300 B.n518 B.n37 585
R301 B.n37 B.n36 585
R302 B.n517 B.n516 585
R303 B.n516 B.n515 585
R304 B.n39 B.n38 585
R305 B.n514 B.n39 585
R306 B.n512 B.n511 585
R307 B.n513 B.n512 585
R308 B.n557 B.n556 585
R309 B.n556 B.n555 585
R310 B.n288 B.n124 530.939
R311 B.n512 B.n44 530.939
R312 B.n290 B.n122 530.939
R313 B.n383 B.n42 530.939
R314 B.n145 B.t2 291.478
R315 B.n139 B.t6 291.478
R316 B.n59 B.t9 291.478
R317 B.n66 B.t13 291.478
R318 B.n384 B.n43 256.663
R319 B.n386 B.n43 256.663
R320 B.n392 B.n43 256.663
R321 B.n394 B.n43 256.663
R322 B.n400 B.n43 256.663
R323 B.n402 B.n43 256.663
R324 B.n408 B.n43 256.663
R325 B.n410 B.n43 256.663
R326 B.n416 B.n43 256.663
R327 B.n418 B.n43 256.663
R328 B.n424 B.n43 256.663
R329 B.n426 B.n43 256.663
R330 B.n432 B.n43 256.663
R331 B.n434 B.n43 256.663
R332 B.n441 B.n43 256.663
R333 B.n443 B.n43 256.663
R334 B.n449 B.n43 256.663
R335 B.n451 B.n43 256.663
R336 B.n457 B.n43 256.663
R337 B.n459 B.n43 256.663
R338 B.n465 B.n43 256.663
R339 B.n467 B.n43 256.663
R340 B.n473 B.n43 256.663
R341 B.n475 B.n43 256.663
R342 B.n481 B.n43 256.663
R343 B.n483 B.n43 256.663
R344 B.n489 B.n43 256.663
R345 B.n491 B.n43 256.663
R346 B.n497 B.n43 256.663
R347 B.n499 B.n43 256.663
R348 B.n505 B.n43 256.663
R349 B.n507 B.n43 256.663
R350 B.n283 B.n123 256.663
R351 B.n126 B.n123 256.663
R352 B.n276 B.n123 256.663
R353 B.n270 B.n123 256.663
R354 B.n268 B.n123 256.663
R355 B.n262 B.n123 256.663
R356 B.n260 B.n123 256.663
R357 B.n254 B.n123 256.663
R358 B.n252 B.n123 256.663
R359 B.n246 B.n123 256.663
R360 B.n244 B.n123 256.663
R361 B.n238 B.n123 256.663
R362 B.n236 B.n123 256.663
R363 B.n229 B.n123 256.663
R364 B.n227 B.n123 256.663
R365 B.n221 B.n123 256.663
R366 B.n219 B.n123 256.663
R367 B.n213 B.n123 256.663
R368 B.n148 B.n123 256.663
R369 B.n207 B.n123 256.663
R370 B.n201 B.n123 256.663
R371 B.n199 B.n123 256.663
R372 B.n193 B.n123 256.663
R373 B.n191 B.n123 256.663
R374 B.n185 B.n123 256.663
R375 B.n183 B.n123 256.663
R376 B.n177 B.n123 256.663
R377 B.n175 B.n123 256.663
R378 B.n169 B.n123 256.663
R379 B.n167 B.n123 256.663
R380 B.n161 B.n123 256.663
R381 B.n145 B.t5 244.252
R382 B.n66 B.t14 244.252
R383 B.n139 B.t8 244.252
R384 B.n59 B.t11 244.252
R385 B.n146 B.t4 198.288
R386 B.n67 B.t15 198.288
R387 B.n140 B.t7 198.288
R388 B.n60 B.t12 198.288
R389 B.n288 B.n118 163.367
R390 B.n296 B.n118 163.367
R391 B.n296 B.n116 163.367
R392 B.n300 B.n116 163.367
R393 B.n300 B.n110 163.367
R394 B.n308 B.n110 163.367
R395 B.n308 B.n108 163.367
R396 B.n312 B.n108 163.367
R397 B.n312 B.n102 163.367
R398 B.n320 B.n102 163.367
R399 B.n320 B.n100 163.367
R400 B.n324 B.n100 163.367
R401 B.n324 B.n94 163.367
R402 B.n332 B.n94 163.367
R403 B.n332 B.n92 163.367
R404 B.n336 B.n92 163.367
R405 B.n336 B.n86 163.367
R406 B.n345 B.n86 163.367
R407 B.n345 B.n84 163.367
R408 B.n349 B.n84 163.367
R409 B.n349 B.n2 163.367
R410 B.n556 B.n2 163.367
R411 B.n556 B.n3 163.367
R412 B.n552 B.n3 163.367
R413 B.n552 B.n9 163.367
R414 B.n548 B.n9 163.367
R415 B.n548 B.n11 163.367
R416 B.n544 B.n11 163.367
R417 B.n544 B.n16 163.367
R418 B.n540 B.n16 163.367
R419 B.n540 B.n18 163.367
R420 B.n536 B.n18 163.367
R421 B.n536 B.n23 163.367
R422 B.n532 B.n23 163.367
R423 B.n532 B.n25 163.367
R424 B.n528 B.n25 163.367
R425 B.n528 B.n30 163.367
R426 B.n524 B.n30 163.367
R427 B.n524 B.n32 163.367
R428 B.n520 B.n32 163.367
R429 B.n520 B.n37 163.367
R430 B.n516 B.n37 163.367
R431 B.n516 B.n39 163.367
R432 B.n512 B.n39 163.367
R433 B.n284 B.n282 163.367
R434 B.n282 B.n281 163.367
R435 B.n278 B.n277 163.367
R436 B.n275 B.n128 163.367
R437 B.n271 B.n269 163.367
R438 B.n267 B.n130 163.367
R439 B.n263 B.n261 163.367
R440 B.n259 B.n132 163.367
R441 B.n255 B.n253 163.367
R442 B.n251 B.n134 163.367
R443 B.n247 B.n245 163.367
R444 B.n243 B.n136 163.367
R445 B.n239 B.n237 163.367
R446 B.n235 B.n138 163.367
R447 B.n230 B.n228 163.367
R448 B.n226 B.n142 163.367
R449 B.n222 B.n220 163.367
R450 B.n218 B.n144 163.367
R451 B.n214 B.n212 163.367
R452 B.n209 B.n208 163.367
R453 B.n206 B.n150 163.367
R454 B.n202 B.n200 163.367
R455 B.n198 B.n152 163.367
R456 B.n194 B.n192 163.367
R457 B.n190 B.n154 163.367
R458 B.n186 B.n184 163.367
R459 B.n182 B.n156 163.367
R460 B.n178 B.n176 163.367
R461 B.n174 B.n158 163.367
R462 B.n170 B.n168 163.367
R463 B.n166 B.n160 163.367
R464 B.n162 B.n122 163.367
R465 B.n290 B.n120 163.367
R466 B.n294 B.n120 163.367
R467 B.n294 B.n114 163.367
R468 B.n302 B.n114 163.367
R469 B.n302 B.n112 163.367
R470 B.n306 B.n112 163.367
R471 B.n306 B.n106 163.367
R472 B.n314 B.n106 163.367
R473 B.n314 B.n104 163.367
R474 B.n318 B.n104 163.367
R475 B.n318 B.n98 163.367
R476 B.n326 B.n98 163.367
R477 B.n326 B.n96 163.367
R478 B.n330 B.n96 163.367
R479 B.n330 B.n90 163.367
R480 B.n338 B.n90 163.367
R481 B.n338 B.n88 163.367
R482 B.n343 B.n88 163.367
R483 B.n343 B.n82 163.367
R484 B.n351 B.n82 163.367
R485 B.n352 B.n351 163.367
R486 B.n352 B.n5 163.367
R487 B.n6 B.n5 163.367
R488 B.n7 B.n6 163.367
R489 B.n357 B.n7 163.367
R490 B.n357 B.n12 163.367
R491 B.n13 B.n12 163.367
R492 B.n14 B.n13 163.367
R493 B.n362 B.n14 163.367
R494 B.n362 B.n19 163.367
R495 B.n20 B.n19 163.367
R496 B.n21 B.n20 163.367
R497 B.n367 B.n21 163.367
R498 B.n367 B.n26 163.367
R499 B.n27 B.n26 163.367
R500 B.n28 B.n27 163.367
R501 B.n372 B.n28 163.367
R502 B.n372 B.n33 163.367
R503 B.n34 B.n33 163.367
R504 B.n35 B.n34 163.367
R505 B.n377 B.n35 163.367
R506 B.n377 B.n40 163.367
R507 B.n41 B.n40 163.367
R508 B.n42 B.n41 163.367
R509 B.n508 B.n506 163.367
R510 B.n504 B.n46 163.367
R511 B.n500 B.n498 163.367
R512 B.n496 B.n48 163.367
R513 B.n492 B.n490 163.367
R514 B.n488 B.n50 163.367
R515 B.n484 B.n482 163.367
R516 B.n480 B.n52 163.367
R517 B.n476 B.n474 163.367
R518 B.n472 B.n54 163.367
R519 B.n468 B.n466 163.367
R520 B.n464 B.n56 163.367
R521 B.n460 B.n458 163.367
R522 B.n456 B.n58 163.367
R523 B.n452 B.n450 163.367
R524 B.n448 B.n63 163.367
R525 B.n444 B.n442 163.367
R526 B.n440 B.n65 163.367
R527 B.n435 B.n433 163.367
R528 B.n431 B.n69 163.367
R529 B.n427 B.n425 163.367
R530 B.n423 B.n71 163.367
R531 B.n419 B.n417 163.367
R532 B.n415 B.n73 163.367
R533 B.n411 B.n409 163.367
R534 B.n407 B.n75 163.367
R535 B.n403 B.n401 163.367
R536 B.n399 B.n77 163.367
R537 B.n395 B.n393 163.367
R538 B.n391 B.n79 163.367
R539 B.n387 B.n385 163.367
R540 B.n289 B.n123 112.436
R541 B.n513 B.n43 112.436
R542 B.n283 B.n124 71.676
R543 B.n281 B.n126 71.676
R544 B.n277 B.n276 71.676
R545 B.n270 B.n128 71.676
R546 B.n269 B.n268 71.676
R547 B.n262 B.n130 71.676
R548 B.n261 B.n260 71.676
R549 B.n254 B.n132 71.676
R550 B.n253 B.n252 71.676
R551 B.n246 B.n134 71.676
R552 B.n245 B.n244 71.676
R553 B.n238 B.n136 71.676
R554 B.n237 B.n236 71.676
R555 B.n229 B.n138 71.676
R556 B.n228 B.n227 71.676
R557 B.n221 B.n142 71.676
R558 B.n220 B.n219 71.676
R559 B.n213 B.n144 71.676
R560 B.n212 B.n148 71.676
R561 B.n208 B.n207 71.676
R562 B.n201 B.n150 71.676
R563 B.n200 B.n199 71.676
R564 B.n193 B.n152 71.676
R565 B.n192 B.n191 71.676
R566 B.n185 B.n154 71.676
R567 B.n184 B.n183 71.676
R568 B.n177 B.n156 71.676
R569 B.n176 B.n175 71.676
R570 B.n169 B.n158 71.676
R571 B.n168 B.n167 71.676
R572 B.n161 B.n160 71.676
R573 B.n507 B.n44 71.676
R574 B.n506 B.n505 71.676
R575 B.n499 B.n46 71.676
R576 B.n498 B.n497 71.676
R577 B.n491 B.n48 71.676
R578 B.n490 B.n489 71.676
R579 B.n483 B.n50 71.676
R580 B.n482 B.n481 71.676
R581 B.n475 B.n52 71.676
R582 B.n474 B.n473 71.676
R583 B.n467 B.n54 71.676
R584 B.n466 B.n465 71.676
R585 B.n459 B.n56 71.676
R586 B.n458 B.n457 71.676
R587 B.n451 B.n58 71.676
R588 B.n450 B.n449 71.676
R589 B.n443 B.n63 71.676
R590 B.n442 B.n441 71.676
R591 B.n434 B.n65 71.676
R592 B.n433 B.n432 71.676
R593 B.n426 B.n69 71.676
R594 B.n425 B.n424 71.676
R595 B.n418 B.n71 71.676
R596 B.n417 B.n416 71.676
R597 B.n410 B.n73 71.676
R598 B.n409 B.n408 71.676
R599 B.n402 B.n75 71.676
R600 B.n401 B.n400 71.676
R601 B.n394 B.n77 71.676
R602 B.n393 B.n392 71.676
R603 B.n386 B.n79 71.676
R604 B.n385 B.n384 71.676
R605 B.n384 B.n383 71.676
R606 B.n387 B.n386 71.676
R607 B.n392 B.n391 71.676
R608 B.n395 B.n394 71.676
R609 B.n400 B.n399 71.676
R610 B.n403 B.n402 71.676
R611 B.n408 B.n407 71.676
R612 B.n411 B.n410 71.676
R613 B.n416 B.n415 71.676
R614 B.n419 B.n418 71.676
R615 B.n424 B.n423 71.676
R616 B.n427 B.n426 71.676
R617 B.n432 B.n431 71.676
R618 B.n435 B.n434 71.676
R619 B.n441 B.n440 71.676
R620 B.n444 B.n443 71.676
R621 B.n449 B.n448 71.676
R622 B.n452 B.n451 71.676
R623 B.n457 B.n456 71.676
R624 B.n460 B.n459 71.676
R625 B.n465 B.n464 71.676
R626 B.n468 B.n467 71.676
R627 B.n473 B.n472 71.676
R628 B.n476 B.n475 71.676
R629 B.n481 B.n480 71.676
R630 B.n484 B.n483 71.676
R631 B.n489 B.n488 71.676
R632 B.n492 B.n491 71.676
R633 B.n497 B.n496 71.676
R634 B.n500 B.n499 71.676
R635 B.n505 B.n504 71.676
R636 B.n508 B.n507 71.676
R637 B.n284 B.n283 71.676
R638 B.n278 B.n126 71.676
R639 B.n276 B.n275 71.676
R640 B.n271 B.n270 71.676
R641 B.n268 B.n267 71.676
R642 B.n263 B.n262 71.676
R643 B.n260 B.n259 71.676
R644 B.n255 B.n254 71.676
R645 B.n252 B.n251 71.676
R646 B.n247 B.n246 71.676
R647 B.n244 B.n243 71.676
R648 B.n239 B.n238 71.676
R649 B.n236 B.n235 71.676
R650 B.n230 B.n229 71.676
R651 B.n227 B.n226 71.676
R652 B.n222 B.n221 71.676
R653 B.n219 B.n218 71.676
R654 B.n214 B.n213 71.676
R655 B.n209 B.n148 71.676
R656 B.n207 B.n206 71.676
R657 B.n202 B.n201 71.676
R658 B.n199 B.n198 71.676
R659 B.n194 B.n193 71.676
R660 B.n191 B.n190 71.676
R661 B.n186 B.n185 71.676
R662 B.n183 B.n182 71.676
R663 B.n178 B.n177 71.676
R664 B.n175 B.n174 71.676
R665 B.n170 B.n169 71.676
R666 B.n167 B.n166 71.676
R667 B.n162 B.n161 71.676
R668 B.n289 B.n119 60.2017
R669 B.n295 B.n119 60.2017
R670 B.n295 B.n115 60.2017
R671 B.n301 B.n115 60.2017
R672 B.n301 B.n111 60.2017
R673 B.n307 B.n111 60.2017
R674 B.n313 B.n107 60.2017
R675 B.n313 B.n103 60.2017
R676 B.n319 B.n103 60.2017
R677 B.n319 B.n99 60.2017
R678 B.n325 B.n99 60.2017
R679 B.n325 B.n95 60.2017
R680 B.n331 B.n95 60.2017
R681 B.n331 B.n91 60.2017
R682 B.n337 B.n91 60.2017
R683 B.n344 B.n87 60.2017
R684 B.n344 B.n83 60.2017
R685 B.n350 B.n83 60.2017
R686 B.n350 B.n4 60.2017
R687 B.n555 B.n4 60.2017
R688 B.n555 B.n554 60.2017
R689 B.n554 B.n553 60.2017
R690 B.n553 B.n8 60.2017
R691 B.n547 B.n8 60.2017
R692 B.n547 B.n546 60.2017
R693 B.n545 B.n15 60.2017
R694 B.n539 B.n15 60.2017
R695 B.n539 B.n538 60.2017
R696 B.n538 B.n537 60.2017
R697 B.n537 B.n22 60.2017
R698 B.n531 B.n22 60.2017
R699 B.n531 B.n530 60.2017
R700 B.n530 B.n529 60.2017
R701 B.n529 B.n29 60.2017
R702 B.n523 B.n522 60.2017
R703 B.n522 B.n521 60.2017
R704 B.n521 B.n36 60.2017
R705 B.n515 B.n36 60.2017
R706 B.n515 B.n514 60.2017
R707 B.n514 B.n513 60.2017
R708 B.n147 B.n146 59.5399
R709 B.n233 B.n140 59.5399
R710 B.n61 B.n60 59.5399
R711 B.n437 B.n67 59.5399
R712 B.n337 B.t1 54.8898
R713 B.t0 B.n545 54.8898
R714 B.n146 B.n145 45.9641
R715 B.n140 B.n139 45.9641
R716 B.n60 B.n59 45.9641
R717 B.n67 B.n66 45.9641
R718 B.n307 B.t3 44.2661
R719 B.n523 B.t10 44.2661
R720 B.n511 B.n510 34.4981
R721 B.n382 B.n381 34.4981
R722 B.n291 B.n121 34.4981
R723 B.n287 B.n286 34.4981
R724 B B.n557 18.0485
R725 B.t3 B.n107 15.9361
R726 B.t10 B.n29 15.9361
R727 B.n510 B.n509 10.6151
R728 B.n509 B.n45 10.6151
R729 B.n503 B.n45 10.6151
R730 B.n503 B.n502 10.6151
R731 B.n502 B.n501 10.6151
R732 B.n501 B.n47 10.6151
R733 B.n495 B.n47 10.6151
R734 B.n495 B.n494 10.6151
R735 B.n494 B.n493 10.6151
R736 B.n493 B.n49 10.6151
R737 B.n487 B.n49 10.6151
R738 B.n487 B.n486 10.6151
R739 B.n486 B.n485 10.6151
R740 B.n485 B.n51 10.6151
R741 B.n479 B.n51 10.6151
R742 B.n479 B.n478 10.6151
R743 B.n478 B.n477 10.6151
R744 B.n477 B.n53 10.6151
R745 B.n471 B.n53 10.6151
R746 B.n471 B.n470 10.6151
R747 B.n470 B.n469 10.6151
R748 B.n469 B.n55 10.6151
R749 B.n463 B.n55 10.6151
R750 B.n463 B.n462 10.6151
R751 B.n462 B.n461 10.6151
R752 B.n461 B.n57 10.6151
R753 B.n455 B.n454 10.6151
R754 B.n454 B.n453 10.6151
R755 B.n453 B.n62 10.6151
R756 B.n447 B.n62 10.6151
R757 B.n447 B.n446 10.6151
R758 B.n446 B.n445 10.6151
R759 B.n445 B.n64 10.6151
R760 B.n439 B.n64 10.6151
R761 B.n439 B.n438 10.6151
R762 B.n436 B.n68 10.6151
R763 B.n430 B.n68 10.6151
R764 B.n430 B.n429 10.6151
R765 B.n429 B.n428 10.6151
R766 B.n428 B.n70 10.6151
R767 B.n422 B.n70 10.6151
R768 B.n422 B.n421 10.6151
R769 B.n421 B.n420 10.6151
R770 B.n420 B.n72 10.6151
R771 B.n414 B.n72 10.6151
R772 B.n414 B.n413 10.6151
R773 B.n413 B.n412 10.6151
R774 B.n412 B.n74 10.6151
R775 B.n406 B.n74 10.6151
R776 B.n406 B.n405 10.6151
R777 B.n405 B.n404 10.6151
R778 B.n404 B.n76 10.6151
R779 B.n398 B.n76 10.6151
R780 B.n398 B.n397 10.6151
R781 B.n397 B.n396 10.6151
R782 B.n396 B.n78 10.6151
R783 B.n390 B.n78 10.6151
R784 B.n390 B.n389 10.6151
R785 B.n389 B.n388 10.6151
R786 B.n388 B.n80 10.6151
R787 B.n382 B.n80 10.6151
R788 B.n292 B.n291 10.6151
R789 B.n293 B.n292 10.6151
R790 B.n293 B.n113 10.6151
R791 B.n303 B.n113 10.6151
R792 B.n304 B.n303 10.6151
R793 B.n305 B.n304 10.6151
R794 B.n305 B.n105 10.6151
R795 B.n315 B.n105 10.6151
R796 B.n316 B.n315 10.6151
R797 B.n317 B.n316 10.6151
R798 B.n317 B.n97 10.6151
R799 B.n327 B.n97 10.6151
R800 B.n328 B.n327 10.6151
R801 B.n329 B.n328 10.6151
R802 B.n329 B.n89 10.6151
R803 B.n339 B.n89 10.6151
R804 B.n340 B.n339 10.6151
R805 B.n342 B.n340 10.6151
R806 B.n342 B.n341 10.6151
R807 B.n341 B.n81 10.6151
R808 B.n353 B.n81 10.6151
R809 B.n354 B.n353 10.6151
R810 B.n355 B.n354 10.6151
R811 B.n356 B.n355 10.6151
R812 B.n358 B.n356 10.6151
R813 B.n359 B.n358 10.6151
R814 B.n360 B.n359 10.6151
R815 B.n361 B.n360 10.6151
R816 B.n363 B.n361 10.6151
R817 B.n364 B.n363 10.6151
R818 B.n365 B.n364 10.6151
R819 B.n366 B.n365 10.6151
R820 B.n368 B.n366 10.6151
R821 B.n369 B.n368 10.6151
R822 B.n370 B.n369 10.6151
R823 B.n371 B.n370 10.6151
R824 B.n373 B.n371 10.6151
R825 B.n374 B.n373 10.6151
R826 B.n375 B.n374 10.6151
R827 B.n376 B.n375 10.6151
R828 B.n378 B.n376 10.6151
R829 B.n379 B.n378 10.6151
R830 B.n380 B.n379 10.6151
R831 B.n381 B.n380 10.6151
R832 B.n286 B.n285 10.6151
R833 B.n285 B.n125 10.6151
R834 B.n280 B.n125 10.6151
R835 B.n280 B.n279 10.6151
R836 B.n279 B.n127 10.6151
R837 B.n274 B.n127 10.6151
R838 B.n274 B.n273 10.6151
R839 B.n273 B.n272 10.6151
R840 B.n272 B.n129 10.6151
R841 B.n266 B.n129 10.6151
R842 B.n266 B.n265 10.6151
R843 B.n265 B.n264 10.6151
R844 B.n264 B.n131 10.6151
R845 B.n258 B.n131 10.6151
R846 B.n258 B.n257 10.6151
R847 B.n257 B.n256 10.6151
R848 B.n256 B.n133 10.6151
R849 B.n250 B.n133 10.6151
R850 B.n250 B.n249 10.6151
R851 B.n249 B.n248 10.6151
R852 B.n248 B.n135 10.6151
R853 B.n242 B.n135 10.6151
R854 B.n242 B.n241 10.6151
R855 B.n241 B.n240 10.6151
R856 B.n240 B.n137 10.6151
R857 B.n234 B.n137 10.6151
R858 B.n232 B.n231 10.6151
R859 B.n231 B.n141 10.6151
R860 B.n225 B.n141 10.6151
R861 B.n225 B.n224 10.6151
R862 B.n224 B.n223 10.6151
R863 B.n223 B.n143 10.6151
R864 B.n217 B.n143 10.6151
R865 B.n217 B.n216 10.6151
R866 B.n216 B.n215 10.6151
R867 B.n211 B.n210 10.6151
R868 B.n210 B.n149 10.6151
R869 B.n205 B.n149 10.6151
R870 B.n205 B.n204 10.6151
R871 B.n204 B.n203 10.6151
R872 B.n203 B.n151 10.6151
R873 B.n197 B.n151 10.6151
R874 B.n197 B.n196 10.6151
R875 B.n196 B.n195 10.6151
R876 B.n195 B.n153 10.6151
R877 B.n189 B.n153 10.6151
R878 B.n189 B.n188 10.6151
R879 B.n188 B.n187 10.6151
R880 B.n187 B.n155 10.6151
R881 B.n181 B.n155 10.6151
R882 B.n181 B.n180 10.6151
R883 B.n180 B.n179 10.6151
R884 B.n179 B.n157 10.6151
R885 B.n173 B.n157 10.6151
R886 B.n173 B.n172 10.6151
R887 B.n172 B.n171 10.6151
R888 B.n171 B.n159 10.6151
R889 B.n165 B.n159 10.6151
R890 B.n165 B.n164 10.6151
R891 B.n164 B.n163 10.6151
R892 B.n163 B.n121 10.6151
R893 B.n287 B.n117 10.6151
R894 B.n297 B.n117 10.6151
R895 B.n298 B.n297 10.6151
R896 B.n299 B.n298 10.6151
R897 B.n299 B.n109 10.6151
R898 B.n309 B.n109 10.6151
R899 B.n310 B.n309 10.6151
R900 B.n311 B.n310 10.6151
R901 B.n311 B.n101 10.6151
R902 B.n321 B.n101 10.6151
R903 B.n322 B.n321 10.6151
R904 B.n323 B.n322 10.6151
R905 B.n323 B.n93 10.6151
R906 B.n333 B.n93 10.6151
R907 B.n334 B.n333 10.6151
R908 B.n335 B.n334 10.6151
R909 B.n335 B.n85 10.6151
R910 B.n346 B.n85 10.6151
R911 B.n347 B.n346 10.6151
R912 B.n348 B.n347 10.6151
R913 B.n348 B.n0 10.6151
R914 B.n551 B.n1 10.6151
R915 B.n551 B.n550 10.6151
R916 B.n550 B.n549 10.6151
R917 B.n549 B.n10 10.6151
R918 B.n543 B.n10 10.6151
R919 B.n543 B.n542 10.6151
R920 B.n542 B.n541 10.6151
R921 B.n541 B.n17 10.6151
R922 B.n535 B.n17 10.6151
R923 B.n535 B.n534 10.6151
R924 B.n534 B.n533 10.6151
R925 B.n533 B.n24 10.6151
R926 B.n527 B.n24 10.6151
R927 B.n527 B.n526 10.6151
R928 B.n526 B.n525 10.6151
R929 B.n525 B.n31 10.6151
R930 B.n519 B.n31 10.6151
R931 B.n519 B.n518 10.6151
R932 B.n518 B.n517 10.6151
R933 B.n517 B.n38 10.6151
R934 B.n511 B.n38 10.6151
R935 B.n61 B.n57 9.36635
R936 B.n437 B.n436 9.36635
R937 B.n234 B.n233 9.36635
R938 B.n211 B.n147 9.36635
R939 B.t1 B.n87 5.31237
R940 B.n546 B.t0 5.31237
R941 B.n557 B.n0 2.81026
R942 B.n557 B.n1 2.81026
R943 B.n455 B.n61 1.24928
R944 B.n438 B.n437 1.24928
R945 B.n233 B.n232 1.24928
R946 B.n215 B.n147 1.24928
R947 VN VN.t1 183.018
R948 VN VN.t0 143.571
R949 VTAIL.n138 VTAIL.n108 214.453
R950 VTAIL.n30 VTAIL.n0 214.453
R951 VTAIL.n102 VTAIL.n72 214.453
R952 VTAIL.n66 VTAIL.n36 214.453
R953 VTAIL.n121 VTAIL.n120 185
R954 VTAIL.n123 VTAIL.n122 185
R955 VTAIL.n116 VTAIL.n115 185
R956 VTAIL.n129 VTAIL.n128 185
R957 VTAIL.n131 VTAIL.n130 185
R958 VTAIL.n112 VTAIL.n111 185
R959 VTAIL.n137 VTAIL.n136 185
R960 VTAIL.n139 VTAIL.n138 185
R961 VTAIL.n13 VTAIL.n12 185
R962 VTAIL.n15 VTAIL.n14 185
R963 VTAIL.n8 VTAIL.n7 185
R964 VTAIL.n21 VTAIL.n20 185
R965 VTAIL.n23 VTAIL.n22 185
R966 VTAIL.n4 VTAIL.n3 185
R967 VTAIL.n29 VTAIL.n28 185
R968 VTAIL.n31 VTAIL.n30 185
R969 VTAIL.n103 VTAIL.n102 185
R970 VTAIL.n101 VTAIL.n100 185
R971 VTAIL.n76 VTAIL.n75 185
R972 VTAIL.n95 VTAIL.n94 185
R973 VTAIL.n93 VTAIL.n92 185
R974 VTAIL.n80 VTAIL.n79 185
R975 VTAIL.n87 VTAIL.n86 185
R976 VTAIL.n85 VTAIL.n84 185
R977 VTAIL.n67 VTAIL.n66 185
R978 VTAIL.n65 VTAIL.n64 185
R979 VTAIL.n40 VTAIL.n39 185
R980 VTAIL.n59 VTAIL.n58 185
R981 VTAIL.n57 VTAIL.n56 185
R982 VTAIL.n44 VTAIL.n43 185
R983 VTAIL.n51 VTAIL.n50 185
R984 VTAIL.n49 VTAIL.n48 185
R985 VTAIL.n119 VTAIL.t2 149.524
R986 VTAIL.n11 VTAIL.t0 149.524
R987 VTAIL.n83 VTAIL.t1 149.524
R988 VTAIL.n47 VTAIL.t3 149.524
R989 VTAIL.n122 VTAIL.n121 104.615
R990 VTAIL.n122 VTAIL.n115 104.615
R991 VTAIL.n129 VTAIL.n115 104.615
R992 VTAIL.n130 VTAIL.n129 104.615
R993 VTAIL.n130 VTAIL.n111 104.615
R994 VTAIL.n137 VTAIL.n111 104.615
R995 VTAIL.n138 VTAIL.n137 104.615
R996 VTAIL.n14 VTAIL.n13 104.615
R997 VTAIL.n14 VTAIL.n7 104.615
R998 VTAIL.n21 VTAIL.n7 104.615
R999 VTAIL.n22 VTAIL.n21 104.615
R1000 VTAIL.n22 VTAIL.n3 104.615
R1001 VTAIL.n29 VTAIL.n3 104.615
R1002 VTAIL.n30 VTAIL.n29 104.615
R1003 VTAIL.n102 VTAIL.n101 104.615
R1004 VTAIL.n101 VTAIL.n75 104.615
R1005 VTAIL.n94 VTAIL.n75 104.615
R1006 VTAIL.n94 VTAIL.n93 104.615
R1007 VTAIL.n93 VTAIL.n79 104.615
R1008 VTAIL.n86 VTAIL.n79 104.615
R1009 VTAIL.n86 VTAIL.n85 104.615
R1010 VTAIL.n66 VTAIL.n65 104.615
R1011 VTAIL.n65 VTAIL.n39 104.615
R1012 VTAIL.n58 VTAIL.n39 104.615
R1013 VTAIL.n58 VTAIL.n57 104.615
R1014 VTAIL.n57 VTAIL.n43 104.615
R1015 VTAIL.n50 VTAIL.n43 104.615
R1016 VTAIL.n50 VTAIL.n49 104.615
R1017 VTAIL.n121 VTAIL.t2 52.3082
R1018 VTAIL.n13 VTAIL.t0 52.3082
R1019 VTAIL.n85 VTAIL.t1 52.3082
R1020 VTAIL.n49 VTAIL.t3 52.3082
R1021 VTAIL.n143 VTAIL.n142 33.5429
R1022 VTAIL.n35 VTAIL.n34 33.5429
R1023 VTAIL.n107 VTAIL.n106 33.5429
R1024 VTAIL.n71 VTAIL.n70 33.5429
R1025 VTAIL.n71 VTAIL.n35 22.6169
R1026 VTAIL.n143 VTAIL.n107 20.5738
R1027 VTAIL.n140 VTAIL.n139 12.8005
R1028 VTAIL.n32 VTAIL.n31 12.8005
R1029 VTAIL.n104 VTAIL.n103 12.8005
R1030 VTAIL.n68 VTAIL.n67 12.8005
R1031 VTAIL.n136 VTAIL.n110 12.0247
R1032 VTAIL.n28 VTAIL.n2 12.0247
R1033 VTAIL.n100 VTAIL.n74 12.0247
R1034 VTAIL.n64 VTAIL.n38 12.0247
R1035 VTAIL.n135 VTAIL.n112 11.249
R1036 VTAIL.n27 VTAIL.n4 11.249
R1037 VTAIL.n99 VTAIL.n76 11.249
R1038 VTAIL.n63 VTAIL.n40 11.249
R1039 VTAIL.n132 VTAIL.n131 10.4732
R1040 VTAIL.n24 VTAIL.n23 10.4732
R1041 VTAIL.n96 VTAIL.n95 10.4732
R1042 VTAIL.n60 VTAIL.n59 10.4732
R1043 VTAIL.n120 VTAIL.n119 10.2747
R1044 VTAIL.n12 VTAIL.n11 10.2747
R1045 VTAIL.n84 VTAIL.n83 10.2747
R1046 VTAIL.n48 VTAIL.n47 10.2747
R1047 VTAIL.n128 VTAIL.n114 9.69747
R1048 VTAIL.n20 VTAIL.n6 9.69747
R1049 VTAIL.n92 VTAIL.n78 9.69747
R1050 VTAIL.n56 VTAIL.n42 9.69747
R1051 VTAIL.n142 VTAIL.n141 9.45567
R1052 VTAIL.n34 VTAIL.n33 9.45567
R1053 VTAIL.n106 VTAIL.n105 9.45567
R1054 VTAIL.n70 VTAIL.n69 9.45567
R1055 VTAIL.n118 VTAIL.n117 9.3005
R1056 VTAIL.n125 VTAIL.n124 9.3005
R1057 VTAIL.n127 VTAIL.n126 9.3005
R1058 VTAIL.n114 VTAIL.n113 9.3005
R1059 VTAIL.n133 VTAIL.n132 9.3005
R1060 VTAIL.n135 VTAIL.n134 9.3005
R1061 VTAIL.n110 VTAIL.n109 9.3005
R1062 VTAIL.n141 VTAIL.n140 9.3005
R1063 VTAIL.n10 VTAIL.n9 9.3005
R1064 VTAIL.n17 VTAIL.n16 9.3005
R1065 VTAIL.n19 VTAIL.n18 9.3005
R1066 VTAIL.n6 VTAIL.n5 9.3005
R1067 VTAIL.n25 VTAIL.n24 9.3005
R1068 VTAIL.n27 VTAIL.n26 9.3005
R1069 VTAIL.n2 VTAIL.n1 9.3005
R1070 VTAIL.n33 VTAIL.n32 9.3005
R1071 VTAIL.n82 VTAIL.n81 9.3005
R1072 VTAIL.n89 VTAIL.n88 9.3005
R1073 VTAIL.n91 VTAIL.n90 9.3005
R1074 VTAIL.n78 VTAIL.n77 9.3005
R1075 VTAIL.n97 VTAIL.n96 9.3005
R1076 VTAIL.n99 VTAIL.n98 9.3005
R1077 VTAIL.n74 VTAIL.n73 9.3005
R1078 VTAIL.n105 VTAIL.n104 9.3005
R1079 VTAIL.n46 VTAIL.n45 9.3005
R1080 VTAIL.n53 VTAIL.n52 9.3005
R1081 VTAIL.n55 VTAIL.n54 9.3005
R1082 VTAIL.n42 VTAIL.n41 9.3005
R1083 VTAIL.n61 VTAIL.n60 9.3005
R1084 VTAIL.n63 VTAIL.n62 9.3005
R1085 VTAIL.n38 VTAIL.n37 9.3005
R1086 VTAIL.n69 VTAIL.n68 9.3005
R1087 VTAIL.n127 VTAIL.n116 8.92171
R1088 VTAIL.n19 VTAIL.n8 8.92171
R1089 VTAIL.n91 VTAIL.n80 8.92171
R1090 VTAIL.n55 VTAIL.n44 8.92171
R1091 VTAIL.n142 VTAIL.n108 8.2187
R1092 VTAIL.n34 VTAIL.n0 8.2187
R1093 VTAIL.n106 VTAIL.n72 8.2187
R1094 VTAIL.n70 VTAIL.n36 8.2187
R1095 VTAIL.n124 VTAIL.n123 8.14595
R1096 VTAIL.n16 VTAIL.n15 8.14595
R1097 VTAIL.n88 VTAIL.n87 8.14595
R1098 VTAIL.n52 VTAIL.n51 8.14595
R1099 VTAIL.n120 VTAIL.n118 7.3702
R1100 VTAIL.n12 VTAIL.n10 7.3702
R1101 VTAIL.n84 VTAIL.n82 7.3702
R1102 VTAIL.n48 VTAIL.n46 7.3702
R1103 VTAIL.n123 VTAIL.n118 5.81868
R1104 VTAIL.n15 VTAIL.n10 5.81868
R1105 VTAIL.n87 VTAIL.n82 5.81868
R1106 VTAIL.n51 VTAIL.n46 5.81868
R1107 VTAIL.n140 VTAIL.n108 5.3904
R1108 VTAIL.n32 VTAIL.n0 5.3904
R1109 VTAIL.n104 VTAIL.n72 5.3904
R1110 VTAIL.n68 VTAIL.n36 5.3904
R1111 VTAIL.n124 VTAIL.n116 5.04292
R1112 VTAIL.n16 VTAIL.n8 5.04292
R1113 VTAIL.n88 VTAIL.n80 5.04292
R1114 VTAIL.n52 VTAIL.n44 5.04292
R1115 VTAIL.n128 VTAIL.n127 4.26717
R1116 VTAIL.n20 VTAIL.n19 4.26717
R1117 VTAIL.n92 VTAIL.n91 4.26717
R1118 VTAIL.n56 VTAIL.n55 4.26717
R1119 VTAIL.n131 VTAIL.n114 3.49141
R1120 VTAIL.n23 VTAIL.n6 3.49141
R1121 VTAIL.n95 VTAIL.n78 3.49141
R1122 VTAIL.n59 VTAIL.n42 3.49141
R1123 VTAIL.n119 VTAIL.n117 2.84305
R1124 VTAIL.n11 VTAIL.n9 2.84305
R1125 VTAIL.n83 VTAIL.n81 2.84305
R1126 VTAIL.n47 VTAIL.n45 2.84305
R1127 VTAIL.n132 VTAIL.n112 2.71565
R1128 VTAIL.n24 VTAIL.n4 2.71565
R1129 VTAIL.n96 VTAIL.n76 2.71565
R1130 VTAIL.n60 VTAIL.n40 2.71565
R1131 VTAIL.n136 VTAIL.n135 1.93989
R1132 VTAIL.n28 VTAIL.n27 1.93989
R1133 VTAIL.n100 VTAIL.n99 1.93989
R1134 VTAIL.n64 VTAIL.n63 1.93989
R1135 VTAIL.n107 VTAIL.n71 1.49188
R1136 VTAIL.n139 VTAIL.n110 1.16414
R1137 VTAIL.n31 VTAIL.n2 1.16414
R1138 VTAIL.n103 VTAIL.n74 1.16414
R1139 VTAIL.n67 VTAIL.n38 1.16414
R1140 VTAIL VTAIL.n35 1.03929
R1141 VTAIL VTAIL.n143 0.453086
R1142 VTAIL.n125 VTAIL.n117 0.155672
R1143 VTAIL.n126 VTAIL.n125 0.155672
R1144 VTAIL.n126 VTAIL.n113 0.155672
R1145 VTAIL.n133 VTAIL.n113 0.155672
R1146 VTAIL.n134 VTAIL.n133 0.155672
R1147 VTAIL.n134 VTAIL.n109 0.155672
R1148 VTAIL.n141 VTAIL.n109 0.155672
R1149 VTAIL.n17 VTAIL.n9 0.155672
R1150 VTAIL.n18 VTAIL.n17 0.155672
R1151 VTAIL.n18 VTAIL.n5 0.155672
R1152 VTAIL.n25 VTAIL.n5 0.155672
R1153 VTAIL.n26 VTAIL.n25 0.155672
R1154 VTAIL.n26 VTAIL.n1 0.155672
R1155 VTAIL.n33 VTAIL.n1 0.155672
R1156 VTAIL.n105 VTAIL.n73 0.155672
R1157 VTAIL.n98 VTAIL.n73 0.155672
R1158 VTAIL.n98 VTAIL.n97 0.155672
R1159 VTAIL.n97 VTAIL.n77 0.155672
R1160 VTAIL.n90 VTAIL.n77 0.155672
R1161 VTAIL.n90 VTAIL.n89 0.155672
R1162 VTAIL.n89 VTAIL.n81 0.155672
R1163 VTAIL.n69 VTAIL.n37 0.155672
R1164 VTAIL.n62 VTAIL.n37 0.155672
R1165 VTAIL.n62 VTAIL.n61 0.155672
R1166 VTAIL.n61 VTAIL.n41 0.155672
R1167 VTAIL.n54 VTAIL.n41 0.155672
R1168 VTAIL.n54 VTAIL.n53 0.155672
R1169 VTAIL.n53 VTAIL.n45 0.155672
R1170 VDD2.n65 VDD2.n35 214.453
R1171 VDD2.n30 VDD2.n0 214.453
R1172 VDD2.n66 VDD2.n65 185
R1173 VDD2.n64 VDD2.n63 185
R1174 VDD2.n39 VDD2.n38 185
R1175 VDD2.n58 VDD2.n57 185
R1176 VDD2.n56 VDD2.n55 185
R1177 VDD2.n43 VDD2.n42 185
R1178 VDD2.n50 VDD2.n49 185
R1179 VDD2.n48 VDD2.n47 185
R1180 VDD2.n13 VDD2.n12 185
R1181 VDD2.n15 VDD2.n14 185
R1182 VDD2.n8 VDD2.n7 185
R1183 VDD2.n21 VDD2.n20 185
R1184 VDD2.n23 VDD2.n22 185
R1185 VDD2.n4 VDD2.n3 185
R1186 VDD2.n29 VDD2.n28 185
R1187 VDD2.n31 VDD2.n30 185
R1188 VDD2.n11 VDD2.t1 149.524
R1189 VDD2.n46 VDD2.t0 149.524
R1190 VDD2.n65 VDD2.n64 104.615
R1191 VDD2.n64 VDD2.n38 104.615
R1192 VDD2.n57 VDD2.n38 104.615
R1193 VDD2.n57 VDD2.n56 104.615
R1194 VDD2.n56 VDD2.n42 104.615
R1195 VDD2.n49 VDD2.n42 104.615
R1196 VDD2.n49 VDD2.n48 104.615
R1197 VDD2.n14 VDD2.n13 104.615
R1198 VDD2.n14 VDD2.n7 104.615
R1199 VDD2.n21 VDD2.n7 104.615
R1200 VDD2.n22 VDD2.n21 104.615
R1201 VDD2.n22 VDD2.n3 104.615
R1202 VDD2.n29 VDD2.n3 104.615
R1203 VDD2.n30 VDD2.n29 104.615
R1204 VDD2.n70 VDD2.n34 84.1312
R1205 VDD2.n48 VDD2.t0 52.3082
R1206 VDD2.n13 VDD2.t1 52.3082
R1207 VDD2.n70 VDD2.n69 50.2217
R1208 VDD2.n67 VDD2.n66 12.8005
R1209 VDD2.n32 VDD2.n31 12.8005
R1210 VDD2.n63 VDD2.n37 12.0247
R1211 VDD2.n28 VDD2.n2 12.0247
R1212 VDD2.n62 VDD2.n39 11.249
R1213 VDD2.n27 VDD2.n4 11.249
R1214 VDD2.n59 VDD2.n58 10.4732
R1215 VDD2.n24 VDD2.n23 10.4732
R1216 VDD2.n47 VDD2.n46 10.2747
R1217 VDD2.n12 VDD2.n11 10.2747
R1218 VDD2.n55 VDD2.n41 9.69747
R1219 VDD2.n20 VDD2.n6 9.69747
R1220 VDD2.n69 VDD2.n68 9.45567
R1221 VDD2.n34 VDD2.n33 9.45567
R1222 VDD2.n45 VDD2.n44 9.3005
R1223 VDD2.n52 VDD2.n51 9.3005
R1224 VDD2.n54 VDD2.n53 9.3005
R1225 VDD2.n41 VDD2.n40 9.3005
R1226 VDD2.n60 VDD2.n59 9.3005
R1227 VDD2.n62 VDD2.n61 9.3005
R1228 VDD2.n37 VDD2.n36 9.3005
R1229 VDD2.n68 VDD2.n67 9.3005
R1230 VDD2.n10 VDD2.n9 9.3005
R1231 VDD2.n17 VDD2.n16 9.3005
R1232 VDD2.n19 VDD2.n18 9.3005
R1233 VDD2.n6 VDD2.n5 9.3005
R1234 VDD2.n25 VDD2.n24 9.3005
R1235 VDD2.n27 VDD2.n26 9.3005
R1236 VDD2.n2 VDD2.n1 9.3005
R1237 VDD2.n33 VDD2.n32 9.3005
R1238 VDD2.n54 VDD2.n43 8.92171
R1239 VDD2.n19 VDD2.n8 8.92171
R1240 VDD2.n69 VDD2.n35 8.2187
R1241 VDD2.n34 VDD2.n0 8.2187
R1242 VDD2.n51 VDD2.n50 8.14595
R1243 VDD2.n16 VDD2.n15 8.14595
R1244 VDD2.n47 VDD2.n45 7.3702
R1245 VDD2.n12 VDD2.n10 7.3702
R1246 VDD2.n50 VDD2.n45 5.81868
R1247 VDD2.n15 VDD2.n10 5.81868
R1248 VDD2.n67 VDD2.n35 5.3904
R1249 VDD2.n32 VDD2.n0 5.3904
R1250 VDD2.n51 VDD2.n43 5.04292
R1251 VDD2.n16 VDD2.n8 5.04292
R1252 VDD2.n55 VDD2.n54 4.26717
R1253 VDD2.n20 VDD2.n19 4.26717
R1254 VDD2.n58 VDD2.n41 3.49141
R1255 VDD2.n23 VDD2.n6 3.49141
R1256 VDD2.n46 VDD2.n44 2.84305
R1257 VDD2.n11 VDD2.n9 2.84305
R1258 VDD2.n59 VDD2.n39 2.71565
R1259 VDD2.n24 VDD2.n4 2.71565
R1260 VDD2.n63 VDD2.n62 1.93989
R1261 VDD2.n28 VDD2.n27 1.93989
R1262 VDD2.n66 VDD2.n37 1.16414
R1263 VDD2.n31 VDD2.n2 1.16414
R1264 VDD2 VDD2.n70 0.569465
R1265 VDD2.n68 VDD2.n36 0.155672
R1266 VDD2.n61 VDD2.n36 0.155672
R1267 VDD2.n61 VDD2.n60 0.155672
R1268 VDD2.n60 VDD2.n40 0.155672
R1269 VDD2.n53 VDD2.n40 0.155672
R1270 VDD2.n53 VDD2.n52 0.155672
R1271 VDD2.n52 VDD2.n44 0.155672
R1272 VDD2.n17 VDD2.n9 0.155672
R1273 VDD2.n18 VDD2.n17 0.155672
R1274 VDD2.n18 VDD2.n5 0.155672
R1275 VDD2.n25 VDD2.n5 0.155672
R1276 VDD2.n26 VDD2.n25 0.155672
R1277 VDD2.n26 VDD2.n1 0.155672
R1278 VDD2.n33 VDD2.n1 0.155672
R1279 VP.n0 VP.t0 182.827
R1280 VP.n0 VP.t1 143.329
R1281 VP VP.n0 0.241678
R1282 VDD1.n30 VDD1.n0 214.453
R1283 VDD1.n65 VDD1.n35 214.453
R1284 VDD1.n31 VDD1.n30 185
R1285 VDD1.n29 VDD1.n28 185
R1286 VDD1.n4 VDD1.n3 185
R1287 VDD1.n23 VDD1.n22 185
R1288 VDD1.n21 VDD1.n20 185
R1289 VDD1.n8 VDD1.n7 185
R1290 VDD1.n15 VDD1.n14 185
R1291 VDD1.n13 VDD1.n12 185
R1292 VDD1.n48 VDD1.n47 185
R1293 VDD1.n50 VDD1.n49 185
R1294 VDD1.n43 VDD1.n42 185
R1295 VDD1.n56 VDD1.n55 185
R1296 VDD1.n58 VDD1.n57 185
R1297 VDD1.n39 VDD1.n38 185
R1298 VDD1.n64 VDD1.n63 185
R1299 VDD1.n66 VDD1.n65 185
R1300 VDD1.n46 VDD1.t0 149.524
R1301 VDD1.n11 VDD1.t1 149.524
R1302 VDD1.n30 VDD1.n29 104.615
R1303 VDD1.n29 VDD1.n3 104.615
R1304 VDD1.n22 VDD1.n3 104.615
R1305 VDD1.n22 VDD1.n21 104.615
R1306 VDD1.n21 VDD1.n7 104.615
R1307 VDD1.n14 VDD1.n7 104.615
R1308 VDD1.n14 VDD1.n13 104.615
R1309 VDD1.n49 VDD1.n48 104.615
R1310 VDD1.n49 VDD1.n42 104.615
R1311 VDD1.n56 VDD1.n42 104.615
R1312 VDD1.n57 VDD1.n56 104.615
R1313 VDD1.n57 VDD1.n38 104.615
R1314 VDD1.n64 VDD1.n38 104.615
R1315 VDD1.n65 VDD1.n64 104.615
R1316 VDD1 VDD1.n69 85.1668
R1317 VDD1.n13 VDD1.t1 52.3082
R1318 VDD1.n48 VDD1.t0 52.3082
R1319 VDD1 VDD1.n34 50.7907
R1320 VDD1.n32 VDD1.n31 12.8005
R1321 VDD1.n67 VDD1.n66 12.8005
R1322 VDD1.n28 VDD1.n2 12.0247
R1323 VDD1.n63 VDD1.n37 12.0247
R1324 VDD1.n27 VDD1.n4 11.249
R1325 VDD1.n62 VDD1.n39 11.249
R1326 VDD1.n24 VDD1.n23 10.4732
R1327 VDD1.n59 VDD1.n58 10.4732
R1328 VDD1.n12 VDD1.n11 10.2747
R1329 VDD1.n47 VDD1.n46 10.2747
R1330 VDD1.n20 VDD1.n6 9.69747
R1331 VDD1.n55 VDD1.n41 9.69747
R1332 VDD1.n34 VDD1.n33 9.45567
R1333 VDD1.n69 VDD1.n68 9.45567
R1334 VDD1.n10 VDD1.n9 9.3005
R1335 VDD1.n17 VDD1.n16 9.3005
R1336 VDD1.n19 VDD1.n18 9.3005
R1337 VDD1.n6 VDD1.n5 9.3005
R1338 VDD1.n25 VDD1.n24 9.3005
R1339 VDD1.n27 VDD1.n26 9.3005
R1340 VDD1.n2 VDD1.n1 9.3005
R1341 VDD1.n33 VDD1.n32 9.3005
R1342 VDD1.n45 VDD1.n44 9.3005
R1343 VDD1.n52 VDD1.n51 9.3005
R1344 VDD1.n54 VDD1.n53 9.3005
R1345 VDD1.n41 VDD1.n40 9.3005
R1346 VDD1.n60 VDD1.n59 9.3005
R1347 VDD1.n62 VDD1.n61 9.3005
R1348 VDD1.n37 VDD1.n36 9.3005
R1349 VDD1.n68 VDD1.n67 9.3005
R1350 VDD1.n19 VDD1.n8 8.92171
R1351 VDD1.n54 VDD1.n43 8.92171
R1352 VDD1.n34 VDD1.n0 8.2187
R1353 VDD1.n69 VDD1.n35 8.2187
R1354 VDD1.n16 VDD1.n15 8.14595
R1355 VDD1.n51 VDD1.n50 8.14595
R1356 VDD1.n12 VDD1.n10 7.3702
R1357 VDD1.n47 VDD1.n45 7.3702
R1358 VDD1.n15 VDD1.n10 5.81868
R1359 VDD1.n50 VDD1.n45 5.81868
R1360 VDD1.n32 VDD1.n0 5.3904
R1361 VDD1.n67 VDD1.n35 5.3904
R1362 VDD1.n16 VDD1.n8 5.04292
R1363 VDD1.n51 VDD1.n43 5.04292
R1364 VDD1.n20 VDD1.n19 4.26717
R1365 VDD1.n55 VDD1.n54 4.26717
R1366 VDD1.n23 VDD1.n6 3.49141
R1367 VDD1.n58 VDD1.n41 3.49141
R1368 VDD1.n11 VDD1.n9 2.84305
R1369 VDD1.n46 VDD1.n44 2.84305
R1370 VDD1.n24 VDD1.n4 2.71565
R1371 VDD1.n59 VDD1.n39 2.71565
R1372 VDD1.n28 VDD1.n27 1.93989
R1373 VDD1.n63 VDD1.n62 1.93989
R1374 VDD1.n31 VDD1.n2 1.16414
R1375 VDD1.n66 VDD1.n37 1.16414
R1376 VDD1.n33 VDD1.n1 0.155672
R1377 VDD1.n26 VDD1.n1 0.155672
R1378 VDD1.n26 VDD1.n25 0.155672
R1379 VDD1.n25 VDD1.n5 0.155672
R1380 VDD1.n18 VDD1.n5 0.155672
R1381 VDD1.n18 VDD1.n17 0.155672
R1382 VDD1.n17 VDD1.n9 0.155672
R1383 VDD1.n52 VDD1.n44 0.155672
R1384 VDD1.n53 VDD1.n52 0.155672
R1385 VDD1.n53 VDD1.n40 0.155672
R1386 VDD1.n60 VDD1.n40 0.155672
R1387 VDD1.n61 VDD1.n60 0.155672
R1388 VDD1.n61 VDD1.n36 0.155672
R1389 VDD1.n68 VDD1.n36 0.155672
C0 VTAIL VP 1.60721f
C1 VDD2 VN 1.68806f
C2 VN VDD1 0.147865f
C3 VDD2 VDD1 0.607321f
C4 VN VTAIL 1.59296f
C5 VDD2 VTAIL 3.72433f
C6 VDD1 VTAIL 3.67677f
C7 VN VP 4.29189f
C8 VDD2 VP 0.309125f
C9 VDD1 VP 1.84746f
C10 VDD2 B 3.330865f
C11 VDD1 B 4.90489f
C12 VTAIL B 4.971925f
C13 VN B 7.36227f
C14 VP B 5.261202f
C15 VDD1.n0 B 0.018348f
C16 VDD1.n1 B 0.013923f
C17 VDD1.n2 B 0.007482f
C18 VDD1.n3 B 0.017684f
C19 VDD1.n4 B 0.007922f
C20 VDD1.n5 B 0.013923f
C21 VDD1.n6 B 0.007482f
C22 VDD1.n7 B 0.017684f
C23 VDD1.n8 B 0.007922f
C24 VDD1.n9 B 0.40201f
C25 VDD1.n10 B 0.007482f
C26 VDD1.t1 B 0.029519f
C27 VDD1.n11 B 0.074487f
C28 VDD1.n12 B 0.012501f
C29 VDD1.n13 B 0.013263f
C30 VDD1.n14 B 0.017684f
C31 VDD1.n15 B 0.007922f
C32 VDD1.n16 B 0.007482f
C33 VDD1.n17 B 0.013923f
C34 VDD1.n18 B 0.013923f
C35 VDD1.n19 B 0.007482f
C36 VDD1.n20 B 0.007922f
C37 VDD1.n21 B 0.017684f
C38 VDD1.n22 B 0.017684f
C39 VDD1.n23 B 0.007922f
C40 VDD1.n24 B 0.007482f
C41 VDD1.n25 B 0.013923f
C42 VDD1.n26 B 0.013923f
C43 VDD1.n27 B 0.007482f
C44 VDD1.n28 B 0.007922f
C45 VDD1.n29 B 0.017684f
C46 VDD1.n30 B 0.035505f
C47 VDD1.n31 B 0.007922f
C48 VDD1.n32 B 0.014629f
C49 VDD1.n33 B 0.033515f
C50 VDD1.n34 B 0.045907f
C51 VDD1.n35 B 0.018348f
C52 VDD1.n36 B 0.013923f
C53 VDD1.n37 B 0.007482f
C54 VDD1.n38 B 0.017684f
C55 VDD1.n39 B 0.007922f
C56 VDD1.n40 B 0.013923f
C57 VDD1.n41 B 0.007482f
C58 VDD1.n42 B 0.017684f
C59 VDD1.n43 B 0.007922f
C60 VDD1.n44 B 0.40201f
C61 VDD1.n45 B 0.007482f
C62 VDD1.t0 B 0.029519f
C63 VDD1.n46 B 0.074487f
C64 VDD1.n47 B 0.012501f
C65 VDD1.n48 B 0.013263f
C66 VDD1.n49 B 0.017684f
C67 VDD1.n50 B 0.007922f
C68 VDD1.n51 B 0.007482f
C69 VDD1.n52 B 0.013923f
C70 VDD1.n53 B 0.013923f
C71 VDD1.n54 B 0.007482f
C72 VDD1.n55 B 0.007922f
C73 VDD1.n56 B 0.017684f
C74 VDD1.n57 B 0.017684f
C75 VDD1.n58 B 0.007922f
C76 VDD1.n59 B 0.007482f
C77 VDD1.n60 B 0.013923f
C78 VDD1.n61 B 0.013923f
C79 VDD1.n62 B 0.007482f
C80 VDD1.n63 B 0.007922f
C81 VDD1.n64 B 0.017684f
C82 VDD1.n65 B 0.035505f
C83 VDD1.n66 B 0.007922f
C84 VDD1.n67 B 0.014629f
C85 VDD1.n68 B 0.033515f
C86 VDD1.n69 B 0.331951f
C87 VP.t0 B 1.26462f
C88 VP.t1 B 1.02334f
C89 VP.n0 B 1.97496f
C90 VDD2.n0 B 0.018607f
C91 VDD2.n1 B 0.01412f
C92 VDD2.n2 B 0.007587f
C93 VDD2.n3 B 0.017934f
C94 VDD2.n4 B 0.008034f
C95 VDD2.n5 B 0.01412f
C96 VDD2.n6 B 0.007587f
C97 VDD2.n7 B 0.017934f
C98 VDD2.n8 B 0.008034f
C99 VDD2.n9 B 0.407676f
C100 VDD2.n10 B 0.007587f
C101 VDD2.t1 B 0.029935f
C102 VDD2.n11 B 0.075537f
C103 VDD2.n12 B 0.012678f
C104 VDD2.n13 B 0.01345f
C105 VDD2.n14 B 0.017934f
C106 VDD2.n15 B 0.008034f
C107 VDD2.n16 B 0.007587f
C108 VDD2.n17 B 0.01412f
C109 VDD2.n18 B 0.01412f
C110 VDD2.n19 B 0.007587f
C111 VDD2.n20 B 0.008034f
C112 VDD2.n21 B 0.017934f
C113 VDD2.n22 B 0.017934f
C114 VDD2.n23 B 0.008034f
C115 VDD2.n24 B 0.007587f
C116 VDD2.n25 B 0.01412f
C117 VDD2.n26 B 0.01412f
C118 VDD2.n27 B 0.007587f
C119 VDD2.n28 B 0.008034f
C120 VDD2.n29 B 0.017934f
C121 VDD2.n30 B 0.036006f
C122 VDD2.n31 B 0.008034f
C123 VDD2.n32 B 0.014836f
C124 VDD2.n33 B 0.033987f
C125 VDD2.n34 B 0.314254f
C126 VDD2.n35 B 0.018607f
C127 VDD2.n36 B 0.01412f
C128 VDD2.n37 B 0.007587f
C129 VDD2.n38 B 0.017934f
C130 VDD2.n39 B 0.008034f
C131 VDD2.n40 B 0.01412f
C132 VDD2.n41 B 0.007587f
C133 VDD2.n42 B 0.017934f
C134 VDD2.n43 B 0.008034f
C135 VDD2.n44 B 0.407676f
C136 VDD2.n45 B 0.007587f
C137 VDD2.t0 B 0.029935f
C138 VDD2.n46 B 0.075537f
C139 VDD2.n47 B 0.012678f
C140 VDD2.n48 B 0.01345f
C141 VDD2.n49 B 0.017934f
C142 VDD2.n50 B 0.008034f
C143 VDD2.n51 B 0.007587f
C144 VDD2.n52 B 0.01412f
C145 VDD2.n53 B 0.01412f
C146 VDD2.n54 B 0.007587f
C147 VDD2.n55 B 0.008034f
C148 VDD2.n56 B 0.017934f
C149 VDD2.n57 B 0.017934f
C150 VDD2.n58 B 0.008034f
C151 VDD2.n59 B 0.007587f
C152 VDD2.n60 B 0.01412f
C153 VDD2.n61 B 0.01412f
C154 VDD2.n62 B 0.007587f
C155 VDD2.n63 B 0.008034f
C156 VDD2.n64 B 0.017934f
C157 VDD2.n65 B 0.036006f
C158 VDD2.n66 B 0.008034f
C159 VDD2.n67 B 0.014836f
C160 VDD2.n68 B 0.033987f
C161 VDD2.n69 B 0.045951f
C162 VDD2.n70 B 1.37829f
C163 VTAIL.n0 B 0.020576f
C164 VTAIL.n1 B 0.015614f
C165 VTAIL.n2 B 0.00839f
C166 VTAIL.n3 B 0.019832f
C167 VTAIL.n4 B 0.008884f
C168 VTAIL.n5 B 0.015614f
C169 VTAIL.n6 B 0.00839f
C170 VTAIL.n7 B 0.019832f
C171 VTAIL.n8 B 0.008884f
C172 VTAIL.n9 B 0.450829f
C173 VTAIL.n10 B 0.00839f
C174 VTAIL.t0 B 0.033104f
C175 VTAIL.n11 B 0.083533f
C176 VTAIL.n12 B 0.01402f
C177 VTAIL.n13 B 0.014874f
C178 VTAIL.n14 B 0.019832f
C179 VTAIL.n15 B 0.008884f
C180 VTAIL.n16 B 0.00839f
C181 VTAIL.n17 B 0.015614f
C182 VTAIL.n18 B 0.015614f
C183 VTAIL.n19 B 0.00839f
C184 VTAIL.n20 B 0.008884f
C185 VTAIL.n21 B 0.019832f
C186 VTAIL.n22 B 0.019832f
C187 VTAIL.n23 B 0.008884f
C188 VTAIL.n24 B 0.00839f
C189 VTAIL.n25 B 0.015614f
C190 VTAIL.n26 B 0.015614f
C191 VTAIL.n27 B 0.00839f
C192 VTAIL.n28 B 0.008884f
C193 VTAIL.n29 B 0.019832f
C194 VTAIL.n30 B 0.039817f
C195 VTAIL.n31 B 0.008884f
C196 VTAIL.n32 B 0.016406f
C197 VTAIL.n33 B 0.037584f
C198 VTAIL.n34 B 0.040044f
C199 VTAIL.n35 B 0.794244f
C200 VTAIL.n36 B 0.020576f
C201 VTAIL.n37 B 0.015614f
C202 VTAIL.n38 B 0.00839f
C203 VTAIL.n39 B 0.019832f
C204 VTAIL.n40 B 0.008884f
C205 VTAIL.n41 B 0.015614f
C206 VTAIL.n42 B 0.00839f
C207 VTAIL.n43 B 0.019832f
C208 VTAIL.n44 B 0.008884f
C209 VTAIL.n45 B 0.450829f
C210 VTAIL.n46 B 0.00839f
C211 VTAIL.t3 B 0.033104f
C212 VTAIL.n47 B 0.083533f
C213 VTAIL.n48 B 0.01402f
C214 VTAIL.n49 B 0.014874f
C215 VTAIL.n50 B 0.019832f
C216 VTAIL.n51 B 0.008884f
C217 VTAIL.n52 B 0.00839f
C218 VTAIL.n53 B 0.015614f
C219 VTAIL.n54 B 0.015614f
C220 VTAIL.n55 B 0.00839f
C221 VTAIL.n56 B 0.008884f
C222 VTAIL.n57 B 0.019832f
C223 VTAIL.n58 B 0.019832f
C224 VTAIL.n59 B 0.008884f
C225 VTAIL.n60 B 0.00839f
C226 VTAIL.n61 B 0.015614f
C227 VTAIL.n62 B 0.015614f
C228 VTAIL.n63 B 0.00839f
C229 VTAIL.n64 B 0.008884f
C230 VTAIL.n65 B 0.019832f
C231 VTAIL.n66 B 0.039817f
C232 VTAIL.n67 B 0.008884f
C233 VTAIL.n68 B 0.016406f
C234 VTAIL.n69 B 0.037584f
C235 VTAIL.n70 B 0.040044f
C236 VTAIL.n71 B 0.817014f
C237 VTAIL.n72 B 0.020576f
C238 VTAIL.n73 B 0.015614f
C239 VTAIL.n74 B 0.00839f
C240 VTAIL.n75 B 0.019832f
C241 VTAIL.n76 B 0.008884f
C242 VTAIL.n77 B 0.015614f
C243 VTAIL.n78 B 0.00839f
C244 VTAIL.n79 B 0.019832f
C245 VTAIL.n80 B 0.008884f
C246 VTAIL.n81 B 0.450829f
C247 VTAIL.n82 B 0.00839f
C248 VTAIL.t1 B 0.033104f
C249 VTAIL.n83 B 0.083533f
C250 VTAIL.n84 B 0.01402f
C251 VTAIL.n85 B 0.014874f
C252 VTAIL.n86 B 0.019832f
C253 VTAIL.n87 B 0.008884f
C254 VTAIL.n88 B 0.00839f
C255 VTAIL.n89 B 0.015614f
C256 VTAIL.n90 B 0.015614f
C257 VTAIL.n91 B 0.00839f
C258 VTAIL.n92 B 0.008884f
C259 VTAIL.n93 B 0.019832f
C260 VTAIL.n94 B 0.019832f
C261 VTAIL.n95 B 0.008884f
C262 VTAIL.n96 B 0.00839f
C263 VTAIL.n97 B 0.015614f
C264 VTAIL.n98 B 0.015614f
C265 VTAIL.n99 B 0.00839f
C266 VTAIL.n100 B 0.008884f
C267 VTAIL.n101 B 0.019832f
C268 VTAIL.n102 B 0.039817f
C269 VTAIL.n103 B 0.008884f
C270 VTAIL.n104 B 0.016406f
C271 VTAIL.n105 B 0.037584f
C272 VTAIL.n106 B 0.040044f
C273 VTAIL.n107 B 0.714221f
C274 VTAIL.n108 B 0.020576f
C275 VTAIL.n109 B 0.015614f
C276 VTAIL.n110 B 0.00839f
C277 VTAIL.n111 B 0.019832f
C278 VTAIL.n112 B 0.008884f
C279 VTAIL.n113 B 0.015614f
C280 VTAIL.n114 B 0.00839f
C281 VTAIL.n115 B 0.019832f
C282 VTAIL.n116 B 0.008884f
C283 VTAIL.n117 B 0.450829f
C284 VTAIL.n118 B 0.00839f
C285 VTAIL.t2 B 0.033104f
C286 VTAIL.n119 B 0.083533f
C287 VTAIL.n120 B 0.01402f
C288 VTAIL.n121 B 0.014874f
C289 VTAIL.n122 B 0.019832f
C290 VTAIL.n123 B 0.008884f
C291 VTAIL.n124 B 0.00839f
C292 VTAIL.n125 B 0.015614f
C293 VTAIL.n126 B 0.015614f
C294 VTAIL.n127 B 0.00839f
C295 VTAIL.n128 B 0.008884f
C296 VTAIL.n129 B 0.019832f
C297 VTAIL.n130 B 0.019832f
C298 VTAIL.n131 B 0.008884f
C299 VTAIL.n132 B 0.00839f
C300 VTAIL.n133 B 0.015614f
C301 VTAIL.n134 B 0.015614f
C302 VTAIL.n135 B 0.00839f
C303 VTAIL.n136 B 0.008884f
C304 VTAIL.n137 B 0.019832f
C305 VTAIL.n138 B 0.039817f
C306 VTAIL.n139 B 0.008884f
C307 VTAIL.n140 B 0.016406f
C308 VTAIL.n141 B 0.037584f
C309 VTAIL.n142 B 0.040044f
C310 VTAIL.n143 B 0.661957f
C311 VN.t0 B 1.0167f
C312 VN.t1 B 1.25886f
.ends

