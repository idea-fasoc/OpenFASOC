* NGSPICE file created from diff_pair_sample_0141.ext - technology: sky130A

.subckt diff_pair_sample_0141 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t11 w_n4122_n4204# sky130_fd_pr__pfet_01v8 ad=6.3102 pd=33.14 as=2.6697 ps=16.51 w=16.18 l=3.61
X1 VTAIL.t3 VN.t0 VDD2.t5 w_n4122_n4204# sky130_fd_pr__pfet_01v8 ad=2.6697 pd=16.51 as=2.6697 ps=16.51 w=16.18 l=3.61
X2 B.t11 B.t9 B.t10 w_n4122_n4204# sky130_fd_pr__pfet_01v8 ad=6.3102 pd=33.14 as=0 ps=0 w=16.18 l=3.61
X3 VDD2.t4 VN.t1 VTAIL.t4 w_n4122_n4204# sky130_fd_pr__pfet_01v8 ad=2.6697 pd=16.51 as=6.3102 ps=33.14 w=16.18 l=3.61
X4 B.t8 B.t6 B.t7 w_n4122_n4204# sky130_fd_pr__pfet_01v8 ad=6.3102 pd=33.14 as=0 ps=0 w=16.18 l=3.61
X5 VDD2.t3 VN.t2 VTAIL.t2 w_n4122_n4204# sky130_fd_pr__pfet_01v8 ad=2.6697 pd=16.51 as=6.3102 ps=33.14 w=16.18 l=3.61
X6 VDD1.t4 VP.t1 VTAIL.t10 w_n4122_n4204# sky130_fd_pr__pfet_01v8 ad=2.6697 pd=16.51 as=6.3102 ps=33.14 w=16.18 l=3.61
X7 VTAIL.t6 VP.t2 VDD1.t3 w_n4122_n4204# sky130_fd_pr__pfet_01v8 ad=2.6697 pd=16.51 as=2.6697 ps=16.51 w=16.18 l=3.61
X8 VTAIL.t8 VP.t3 VDD1.t2 w_n4122_n4204# sky130_fd_pr__pfet_01v8 ad=2.6697 pd=16.51 as=2.6697 ps=16.51 w=16.18 l=3.61
X9 B.t5 B.t3 B.t4 w_n4122_n4204# sky130_fd_pr__pfet_01v8 ad=6.3102 pd=33.14 as=0 ps=0 w=16.18 l=3.61
X10 VDD2.t2 VN.t3 VTAIL.t5 w_n4122_n4204# sky130_fd_pr__pfet_01v8 ad=6.3102 pd=33.14 as=2.6697 ps=16.51 w=16.18 l=3.61
X11 B.t2 B.t0 B.t1 w_n4122_n4204# sky130_fd_pr__pfet_01v8 ad=6.3102 pd=33.14 as=0 ps=0 w=16.18 l=3.61
X12 VDD1.t1 VP.t4 VTAIL.t7 w_n4122_n4204# sky130_fd_pr__pfet_01v8 ad=6.3102 pd=33.14 as=2.6697 ps=16.51 w=16.18 l=3.61
X13 VDD1.t0 VP.t5 VTAIL.t9 w_n4122_n4204# sky130_fd_pr__pfet_01v8 ad=2.6697 pd=16.51 as=6.3102 ps=33.14 w=16.18 l=3.61
X14 VTAIL.t0 VN.t4 VDD2.t1 w_n4122_n4204# sky130_fd_pr__pfet_01v8 ad=2.6697 pd=16.51 as=2.6697 ps=16.51 w=16.18 l=3.61
X15 VDD2.t0 VN.t5 VTAIL.t1 w_n4122_n4204# sky130_fd_pr__pfet_01v8 ad=6.3102 pd=33.14 as=2.6697 ps=16.51 w=16.18 l=3.61
R0 VP.n16 VP.n13 161.3
R1 VP.n18 VP.n17 161.3
R2 VP.n19 VP.n12 161.3
R3 VP.n21 VP.n20 161.3
R4 VP.n22 VP.n11 161.3
R5 VP.n24 VP.n23 161.3
R6 VP.n25 VP.n10 161.3
R7 VP.n27 VP.n26 161.3
R8 VP.n55 VP.n54 161.3
R9 VP.n53 VP.n1 161.3
R10 VP.n52 VP.n51 161.3
R11 VP.n50 VP.n2 161.3
R12 VP.n49 VP.n48 161.3
R13 VP.n47 VP.n3 161.3
R14 VP.n46 VP.n45 161.3
R15 VP.n44 VP.n4 161.3
R16 VP.n43 VP.n42 161.3
R17 VP.n40 VP.n5 161.3
R18 VP.n39 VP.n38 161.3
R19 VP.n37 VP.n6 161.3
R20 VP.n36 VP.n35 161.3
R21 VP.n34 VP.n7 161.3
R22 VP.n33 VP.n32 161.3
R23 VP.n31 VP.n8 161.3
R24 VP.n15 VP.t0 141.381
R25 VP.n29 VP.t4 108.016
R26 VP.n41 VP.t3 108.016
R27 VP.n0 VP.t1 108.016
R28 VP.n9 VP.t5 108.016
R29 VP.n14 VP.t2 108.016
R30 VP.n30 VP.n29 80.9007
R31 VP.n56 VP.n0 80.9007
R32 VP.n28 VP.n9 80.9007
R33 VP.n15 VP.n14 62.5184
R34 VP.n35 VP.n6 56.5617
R35 VP.n48 VP.n2 56.5617
R36 VP.n20 VP.n11 56.5617
R37 VP.n30 VP.n28 55.9086
R38 VP.n33 VP.n8 24.5923
R39 VP.n34 VP.n33 24.5923
R40 VP.n35 VP.n34 24.5923
R41 VP.n39 VP.n6 24.5923
R42 VP.n40 VP.n39 24.5923
R43 VP.n42 VP.n40 24.5923
R44 VP.n46 VP.n4 24.5923
R45 VP.n47 VP.n46 24.5923
R46 VP.n48 VP.n47 24.5923
R47 VP.n52 VP.n2 24.5923
R48 VP.n53 VP.n52 24.5923
R49 VP.n54 VP.n53 24.5923
R50 VP.n24 VP.n11 24.5923
R51 VP.n25 VP.n24 24.5923
R52 VP.n26 VP.n25 24.5923
R53 VP.n18 VP.n13 24.5923
R54 VP.n19 VP.n18 24.5923
R55 VP.n20 VP.n19 24.5923
R56 VP.n42 VP.n41 12.2964
R57 VP.n41 VP.n4 12.2964
R58 VP.n14 VP.n13 12.2964
R59 VP.n29 VP.n8 9.3454
R60 VP.n54 VP.n0 9.3454
R61 VP.n26 VP.n9 9.3454
R62 VP.n16 VP.n15 3.16704
R63 VP.n28 VP.n27 0.354861
R64 VP.n31 VP.n30 0.354861
R65 VP.n56 VP.n55 0.354861
R66 VP VP.n56 0.267071
R67 VP.n17 VP.n16 0.189894
R68 VP.n17 VP.n12 0.189894
R69 VP.n21 VP.n12 0.189894
R70 VP.n22 VP.n21 0.189894
R71 VP.n23 VP.n22 0.189894
R72 VP.n23 VP.n10 0.189894
R73 VP.n27 VP.n10 0.189894
R74 VP.n32 VP.n31 0.189894
R75 VP.n32 VP.n7 0.189894
R76 VP.n36 VP.n7 0.189894
R77 VP.n37 VP.n36 0.189894
R78 VP.n38 VP.n37 0.189894
R79 VP.n38 VP.n5 0.189894
R80 VP.n43 VP.n5 0.189894
R81 VP.n44 VP.n43 0.189894
R82 VP.n45 VP.n44 0.189894
R83 VP.n45 VP.n3 0.189894
R84 VP.n49 VP.n3 0.189894
R85 VP.n50 VP.n49 0.189894
R86 VP.n51 VP.n50 0.189894
R87 VP.n51 VP.n1 0.189894
R88 VP.n55 VP.n1 0.189894
R89 VTAIL.n362 VTAIL.n278 756.745
R90 VTAIL.n86 VTAIL.n2 756.745
R91 VTAIL.n272 VTAIL.n188 756.745
R92 VTAIL.n180 VTAIL.n96 756.745
R93 VTAIL.n306 VTAIL.n305 585
R94 VTAIL.n311 VTAIL.n310 585
R95 VTAIL.n313 VTAIL.n312 585
R96 VTAIL.n302 VTAIL.n301 585
R97 VTAIL.n319 VTAIL.n318 585
R98 VTAIL.n321 VTAIL.n320 585
R99 VTAIL.n298 VTAIL.n297 585
R100 VTAIL.n327 VTAIL.n326 585
R101 VTAIL.n329 VTAIL.n328 585
R102 VTAIL.n294 VTAIL.n293 585
R103 VTAIL.n335 VTAIL.n334 585
R104 VTAIL.n337 VTAIL.n336 585
R105 VTAIL.n290 VTAIL.n289 585
R106 VTAIL.n343 VTAIL.n342 585
R107 VTAIL.n345 VTAIL.n344 585
R108 VTAIL.n286 VTAIL.n285 585
R109 VTAIL.n352 VTAIL.n351 585
R110 VTAIL.n353 VTAIL.n284 585
R111 VTAIL.n355 VTAIL.n354 585
R112 VTAIL.n282 VTAIL.n281 585
R113 VTAIL.n361 VTAIL.n360 585
R114 VTAIL.n363 VTAIL.n362 585
R115 VTAIL.n30 VTAIL.n29 585
R116 VTAIL.n35 VTAIL.n34 585
R117 VTAIL.n37 VTAIL.n36 585
R118 VTAIL.n26 VTAIL.n25 585
R119 VTAIL.n43 VTAIL.n42 585
R120 VTAIL.n45 VTAIL.n44 585
R121 VTAIL.n22 VTAIL.n21 585
R122 VTAIL.n51 VTAIL.n50 585
R123 VTAIL.n53 VTAIL.n52 585
R124 VTAIL.n18 VTAIL.n17 585
R125 VTAIL.n59 VTAIL.n58 585
R126 VTAIL.n61 VTAIL.n60 585
R127 VTAIL.n14 VTAIL.n13 585
R128 VTAIL.n67 VTAIL.n66 585
R129 VTAIL.n69 VTAIL.n68 585
R130 VTAIL.n10 VTAIL.n9 585
R131 VTAIL.n76 VTAIL.n75 585
R132 VTAIL.n77 VTAIL.n8 585
R133 VTAIL.n79 VTAIL.n78 585
R134 VTAIL.n6 VTAIL.n5 585
R135 VTAIL.n85 VTAIL.n84 585
R136 VTAIL.n87 VTAIL.n86 585
R137 VTAIL.n273 VTAIL.n272 585
R138 VTAIL.n271 VTAIL.n270 585
R139 VTAIL.n192 VTAIL.n191 585
R140 VTAIL.n265 VTAIL.n264 585
R141 VTAIL.n263 VTAIL.n194 585
R142 VTAIL.n262 VTAIL.n261 585
R143 VTAIL.n197 VTAIL.n195 585
R144 VTAIL.n256 VTAIL.n255 585
R145 VTAIL.n254 VTAIL.n253 585
R146 VTAIL.n201 VTAIL.n200 585
R147 VTAIL.n248 VTAIL.n247 585
R148 VTAIL.n246 VTAIL.n245 585
R149 VTAIL.n205 VTAIL.n204 585
R150 VTAIL.n240 VTAIL.n239 585
R151 VTAIL.n238 VTAIL.n237 585
R152 VTAIL.n209 VTAIL.n208 585
R153 VTAIL.n232 VTAIL.n231 585
R154 VTAIL.n230 VTAIL.n229 585
R155 VTAIL.n213 VTAIL.n212 585
R156 VTAIL.n224 VTAIL.n223 585
R157 VTAIL.n222 VTAIL.n221 585
R158 VTAIL.n217 VTAIL.n216 585
R159 VTAIL.n181 VTAIL.n180 585
R160 VTAIL.n179 VTAIL.n178 585
R161 VTAIL.n100 VTAIL.n99 585
R162 VTAIL.n173 VTAIL.n172 585
R163 VTAIL.n171 VTAIL.n102 585
R164 VTAIL.n170 VTAIL.n169 585
R165 VTAIL.n105 VTAIL.n103 585
R166 VTAIL.n164 VTAIL.n163 585
R167 VTAIL.n162 VTAIL.n161 585
R168 VTAIL.n109 VTAIL.n108 585
R169 VTAIL.n156 VTAIL.n155 585
R170 VTAIL.n154 VTAIL.n153 585
R171 VTAIL.n113 VTAIL.n112 585
R172 VTAIL.n148 VTAIL.n147 585
R173 VTAIL.n146 VTAIL.n145 585
R174 VTAIL.n117 VTAIL.n116 585
R175 VTAIL.n140 VTAIL.n139 585
R176 VTAIL.n138 VTAIL.n137 585
R177 VTAIL.n121 VTAIL.n120 585
R178 VTAIL.n132 VTAIL.n131 585
R179 VTAIL.n130 VTAIL.n129 585
R180 VTAIL.n125 VTAIL.n124 585
R181 VTAIL.n307 VTAIL.t4 327.466
R182 VTAIL.n31 VTAIL.t10 327.466
R183 VTAIL.n218 VTAIL.t9 327.466
R184 VTAIL.n126 VTAIL.t2 327.466
R185 VTAIL.n311 VTAIL.n305 171.744
R186 VTAIL.n312 VTAIL.n311 171.744
R187 VTAIL.n312 VTAIL.n301 171.744
R188 VTAIL.n319 VTAIL.n301 171.744
R189 VTAIL.n320 VTAIL.n319 171.744
R190 VTAIL.n320 VTAIL.n297 171.744
R191 VTAIL.n327 VTAIL.n297 171.744
R192 VTAIL.n328 VTAIL.n327 171.744
R193 VTAIL.n328 VTAIL.n293 171.744
R194 VTAIL.n335 VTAIL.n293 171.744
R195 VTAIL.n336 VTAIL.n335 171.744
R196 VTAIL.n336 VTAIL.n289 171.744
R197 VTAIL.n343 VTAIL.n289 171.744
R198 VTAIL.n344 VTAIL.n343 171.744
R199 VTAIL.n344 VTAIL.n285 171.744
R200 VTAIL.n352 VTAIL.n285 171.744
R201 VTAIL.n353 VTAIL.n352 171.744
R202 VTAIL.n354 VTAIL.n353 171.744
R203 VTAIL.n354 VTAIL.n281 171.744
R204 VTAIL.n361 VTAIL.n281 171.744
R205 VTAIL.n362 VTAIL.n361 171.744
R206 VTAIL.n35 VTAIL.n29 171.744
R207 VTAIL.n36 VTAIL.n35 171.744
R208 VTAIL.n36 VTAIL.n25 171.744
R209 VTAIL.n43 VTAIL.n25 171.744
R210 VTAIL.n44 VTAIL.n43 171.744
R211 VTAIL.n44 VTAIL.n21 171.744
R212 VTAIL.n51 VTAIL.n21 171.744
R213 VTAIL.n52 VTAIL.n51 171.744
R214 VTAIL.n52 VTAIL.n17 171.744
R215 VTAIL.n59 VTAIL.n17 171.744
R216 VTAIL.n60 VTAIL.n59 171.744
R217 VTAIL.n60 VTAIL.n13 171.744
R218 VTAIL.n67 VTAIL.n13 171.744
R219 VTAIL.n68 VTAIL.n67 171.744
R220 VTAIL.n68 VTAIL.n9 171.744
R221 VTAIL.n76 VTAIL.n9 171.744
R222 VTAIL.n77 VTAIL.n76 171.744
R223 VTAIL.n78 VTAIL.n77 171.744
R224 VTAIL.n78 VTAIL.n5 171.744
R225 VTAIL.n85 VTAIL.n5 171.744
R226 VTAIL.n86 VTAIL.n85 171.744
R227 VTAIL.n272 VTAIL.n271 171.744
R228 VTAIL.n271 VTAIL.n191 171.744
R229 VTAIL.n264 VTAIL.n191 171.744
R230 VTAIL.n264 VTAIL.n263 171.744
R231 VTAIL.n263 VTAIL.n262 171.744
R232 VTAIL.n262 VTAIL.n195 171.744
R233 VTAIL.n255 VTAIL.n195 171.744
R234 VTAIL.n255 VTAIL.n254 171.744
R235 VTAIL.n254 VTAIL.n200 171.744
R236 VTAIL.n247 VTAIL.n200 171.744
R237 VTAIL.n247 VTAIL.n246 171.744
R238 VTAIL.n246 VTAIL.n204 171.744
R239 VTAIL.n239 VTAIL.n204 171.744
R240 VTAIL.n239 VTAIL.n238 171.744
R241 VTAIL.n238 VTAIL.n208 171.744
R242 VTAIL.n231 VTAIL.n208 171.744
R243 VTAIL.n231 VTAIL.n230 171.744
R244 VTAIL.n230 VTAIL.n212 171.744
R245 VTAIL.n223 VTAIL.n212 171.744
R246 VTAIL.n223 VTAIL.n222 171.744
R247 VTAIL.n222 VTAIL.n216 171.744
R248 VTAIL.n180 VTAIL.n179 171.744
R249 VTAIL.n179 VTAIL.n99 171.744
R250 VTAIL.n172 VTAIL.n99 171.744
R251 VTAIL.n172 VTAIL.n171 171.744
R252 VTAIL.n171 VTAIL.n170 171.744
R253 VTAIL.n170 VTAIL.n103 171.744
R254 VTAIL.n163 VTAIL.n103 171.744
R255 VTAIL.n163 VTAIL.n162 171.744
R256 VTAIL.n162 VTAIL.n108 171.744
R257 VTAIL.n155 VTAIL.n108 171.744
R258 VTAIL.n155 VTAIL.n154 171.744
R259 VTAIL.n154 VTAIL.n112 171.744
R260 VTAIL.n147 VTAIL.n112 171.744
R261 VTAIL.n147 VTAIL.n146 171.744
R262 VTAIL.n146 VTAIL.n116 171.744
R263 VTAIL.n139 VTAIL.n116 171.744
R264 VTAIL.n139 VTAIL.n138 171.744
R265 VTAIL.n138 VTAIL.n120 171.744
R266 VTAIL.n131 VTAIL.n120 171.744
R267 VTAIL.n131 VTAIL.n130 171.744
R268 VTAIL.n130 VTAIL.n124 171.744
R269 VTAIL.t4 VTAIL.n305 85.8723
R270 VTAIL.t10 VTAIL.n29 85.8723
R271 VTAIL.t9 VTAIL.n216 85.8723
R272 VTAIL.t2 VTAIL.n124 85.8723
R273 VTAIL.n187 VTAIL.n186 55.0627
R274 VTAIL.n95 VTAIL.n94 55.0627
R275 VTAIL.n1 VTAIL.n0 55.0625
R276 VTAIL.n93 VTAIL.n92 55.0625
R277 VTAIL.n367 VTAIL.n366 34.1247
R278 VTAIL.n91 VTAIL.n90 34.1247
R279 VTAIL.n277 VTAIL.n276 34.1247
R280 VTAIL.n185 VTAIL.n184 34.1247
R281 VTAIL.n95 VTAIL.n93 33.1083
R282 VTAIL.n367 VTAIL.n277 29.7117
R283 VTAIL.n307 VTAIL.n306 16.3895
R284 VTAIL.n31 VTAIL.n30 16.3895
R285 VTAIL.n218 VTAIL.n217 16.3895
R286 VTAIL.n126 VTAIL.n125 16.3895
R287 VTAIL.n355 VTAIL.n284 13.1884
R288 VTAIL.n79 VTAIL.n8 13.1884
R289 VTAIL.n265 VTAIL.n194 13.1884
R290 VTAIL.n173 VTAIL.n102 13.1884
R291 VTAIL.n310 VTAIL.n309 12.8005
R292 VTAIL.n351 VTAIL.n350 12.8005
R293 VTAIL.n356 VTAIL.n282 12.8005
R294 VTAIL.n34 VTAIL.n33 12.8005
R295 VTAIL.n75 VTAIL.n74 12.8005
R296 VTAIL.n80 VTAIL.n6 12.8005
R297 VTAIL.n266 VTAIL.n192 12.8005
R298 VTAIL.n261 VTAIL.n196 12.8005
R299 VTAIL.n221 VTAIL.n220 12.8005
R300 VTAIL.n174 VTAIL.n100 12.8005
R301 VTAIL.n169 VTAIL.n104 12.8005
R302 VTAIL.n129 VTAIL.n128 12.8005
R303 VTAIL.n313 VTAIL.n304 12.0247
R304 VTAIL.n349 VTAIL.n286 12.0247
R305 VTAIL.n360 VTAIL.n359 12.0247
R306 VTAIL.n37 VTAIL.n28 12.0247
R307 VTAIL.n73 VTAIL.n10 12.0247
R308 VTAIL.n84 VTAIL.n83 12.0247
R309 VTAIL.n270 VTAIL.n269 12.0247
R310 VTAIL.n260 VTAIL.n197 12.0247
R311 VTAIL.n224 VTAIL.n215 12.0247
R312 VTAIL.n178 VTAIL.n177 12.0247
R313 VTAIL.n168 VTAIL.n105 12.0247
R314 VTAIL.n132 VTAIL.n123 12.0247
R315 VTAIL.n314 VTAIL.n302 11.249
R316 VTAIL.n346 VTAIL.n345 11.249
R317 VTAIL.n363 VTAIL.n280 11.249
R318 VTAIL.n38 VTAIL.n26 11.249
R319 VTAIL.n70 VTAIL.n69 11.249
R320 VTAIL.n87 VTAIL.n4 11.249
R321 VTAIL.n273 VTAIL.n190 11.249
R322 VTAIL.n257 VTAIL.n256 11.249
R323 VTAIL.n225 VTAIL.n213 11.249
R324 VTAIL.n181 VTAIL.n98 11.249
R325 VTAIL.n165 VTAIL.n164 11.249
R326 VTAIL.n133 VTAIL.n121 11.249
R327 VTAIL.n318 VTAIL.n317 10.4732
R328 VTAIL.n342 VTAIL.n288 10.4732
R329 VTAIL.n364 VTAIL.n278 10.4732
R330 VTAIL.n42 VTAIL.n41 10.4732
R331 VTAIL.n66 VTAIL.n12 10.4732
R332 VTAIL.n88 VTAIL.n2 10.4732
R333 VTAIL.n274 VTAIL.n188 10.4732
R334 VTAIL.n253 VTAIL.n199 10.4732
R335 VTAIL.n229 VTAIL.n228 10.4732
R336 VTAIL.n182 VTAIL.n96 10.4732
R337 VTAIL.n161 VTAIL.n107 10.4732
R338 VTAIL.n137 VTAIL.n136 10.4732
R339 VTAIL.n321 VTAIL.n300 9.69747
R340 VTAIL.n341 VTAIL.n290 9.69747
R341 VTAIL.n45 VTAIL.n24 9.69747
R342 VTAIL.n65 VTAIL.n14 9.69747
R343 VTAIL.n252 VTAIL.n201 9.69747
R344 VTAIL.n232 VTAIL.n211 9.69747
R345 VTAIL.n160 VTAIL.n109 9.69747
R346 VTAIL.n140 VTAIL.n119 9.69747
R347 VTAIL.n366 VTAIL.n365 9.45567
R348 VTAIL.n90 VTAIL.n89 9.45567
R349 VTAIL.n276 VTAIL.n275 9.45567
R350 VTAIL.n184 VTAIL.n183 9.45567
R351 VTAIL.n365 VTAIL.n364 9.3005
R352 VTAIL.n280 VTAIL.n279 9.3005
R353 VTAIL.n359 VTAIL.n358 9.3005
R354 VTAIL.n357 VTAIL.n356 9.3005
R355 VTAIL.n296 VTAIL.n295 9.3005
R356 VTAIL.n325 VTAIL.n324 9.3005
R357 VTAIL.n323 VTAIL.n322 9.3005
R358 VTAIL.n300 VTAIL.n299 9.3005
R359 VTAIL.n317 VTAIL.n316 9.3005
R360 VTAIL.n315 VTAIL.n314 9.3005
R361 VTAIL.n304 VTAIL.n303 9.3005
R362 VTAIL.n309 VTAIL.n308 9.3005
R363 VTAIL.n331 VTAIL.n330 9.3005
R364 VTAIL.n333 VTAIL.n332 9.3005
R365 VTAIL.n292 VTAIL.n291 9.3005
R366 VTAIL.n339 VTAIL.n338 9.3005
R367 VTAIL.n341 VTAIL.n340 9.3005
R368 VTAIL.n288 VTAIL.n287 9.3005
R369 VTAIL.n347 VTAIL.n346 9.3005
R370 VTAIL.n349 VTAIL.n348 9.3005
R371 VTAIL.n350 VTAIL.n283 9.3005
R372 VTAIL.n89 VTAIL.n88 9.3005
R373 VTAIL.n4 VTAIL.n3 9.3005
R374 VTAIL.n83 VTAIL.n82 9.3005
R375 VTAIL.n81 VTAIL.n80 9.3005
R376 VTAIL.n20 VTAIL.n19 9.3005
R377 VTAIL.n49 VTAIL.n48 9.3005
R378 VTAIL.n47 VTAIL.n46 9.3005
R379 VTAIL.n24 VTAIL.n23 9.3005
R380 VTAIL.n41 VTAIL.n40 9.3005
R381 VTAIL.n39 VTAIL.n38 9.3005
R382 VTAIL.n28 VTAIL.n27 9.3005
R383 VTAIL.n33 VTAIL.n32 9.3005
R384 VTAIL.n55 VTAIL.n54 9.3005
R385 VTAIL.n57 VTAIL.n56 9.3005
R386 VTAIL.n16 VTAIL.n15 9.3005
R387 VTAIL.n63 VTAIL.n62 9.3005
R388 VTAIL.n65 VTAIL.n64 9.3005
R389 VTAIL.n12 VTAIL.n11 9.3005
R390 VTAIL.n71 VTAIL.n70 9.3005
R391 VTAIL.n73 VTAIL.n72 9.3005
R392 VTAIL.n74 VTAIL.n7 9.3005
R393 VTAIL.n244 VTAIL.n243 9.3005
R394 VTAIL.n203 VTAIL.n202 9.3005
R395 VTAIL.n250 VTAIL.n249 9.3005
R396 VTAIL.n252 VTAIL.n251 9.3005
R397 VTAIL.n199 VTAIL.n198 9.3005
R398 VTAIL.n258 VTAIL.n257 9.3005
R399 VTAIL.n260 VTAIL.n259 9.3005
R400 VTAIL.n196 VTAIL.n193 9.3005
R401 VTAIL.n275 VTAIL.n274 9.3005
R402 VTAIL.n190 VTAIL.n189 9.3005
R403 VTAIL.n269 VTAIL.n268 9.3005
R404 VTAIL.n267 VTAIL.n266 9.3005
R405 VTAIL.n242 VTAIL.n241 9.3005
R406 VTAIL.n207 VTAIL.n206 9.3005
R407 VTAIL.n236 VTAIL.n235 9.3005
R408 VTAIL.n234 VTAIL.n233 9.3005
R409 VTAIL.n211 VTAIL.n210 9.3005
R410 VTAIL.n228 VTAIL.n227 9.3005
R411 VTAIL.n226 VTAIL.n225 9.3005
R412 VTAIL.n215 VTAIL.n214 9.3005
R413 VTAIL.n220 VTAIL.n219 9.3005
R414 VTAIL.n152 VTAIL.n151 9.3005
R415 VTAIL.n111 VTAIL.n110 9.3005
R416 VTAIL.n158 VTAIL.n157 9.3005
R417 VTAIL.n160 VTAIL.n159 9.3005
R418 VTAIL.n107 VTAIL.n106 9.3005
R419 VTAIL.n166 VTAIL.n165 9.3005
R420 VTAIL.n168 VTAIL.n167 9.3005
R421 VTAIL.n104 VTAIL.n101 9.3005
R422 VTAIL.n183 VTAIL.n182 9.3005
R423 VTAIL.n98 VTAIL.n97 9.3005
R424 VTAIL.n177 VTAIL.n176 9.3005
R425 VTAIL.n175 VTAIL.n174 9.3005
R426 VTAIL.n150 VTAIL.n149 9.3005
R427 VTAIL.n115 VTAIL.n114 9.3005
R428 VTAIL.n144 VTAIL.n143 9.3005
R429 VTAIL.n142 VTAIL.n141 9.3005
R430 VTAIL.n119 VTAIL.n118 9.3005
R431 VTAIL.n136 VTAIL.n135 9.3005
R432 VTAIL.n134 VTAIL.n133 9.3005
R433 VTAIL.n123 VTAIL.n122 9.3005
R434 VTAIL.n128 VTAIL.n127 9.3005
R435 VTAIL.n322 VTAIL.n298 8.92171
R436 VTAIL.n338 VTAIL.n337 8.92171
R437 VTAIL.n46 VTAIL.n22 8.92171
R438 VTAIL.n62 VTAIL.n61 8.92171
R439 VTAIL.n249 VTAIL.n248 8.92171
R440 VTAIL.n233 VTAIL.n209 8.92171
R441 VTAIL.n157 VTAIL.n156 8.92171
R442 VTAIL.n141 VTAIL.n117 8.92171
R443 VTAIL.n326 VTAIL.n325 8.14595
R444 VTAIL.n334 VTAIL.n292 8.14595
R445 VTAIL.n50 VTAIL.n49 8.14595
R446 VTAIL.n58 VTAIL.n16 8.14595
R447 VTAIL.n245 VTAIL.n203 8.14595
R448 VTAIL.n237 VTAIL.n236 8.14595
R449 VTAIL.n153 VTAIL.n111 8.14595
R450 VTAIL.n145 VTAIL.n144 8.14595
R451 VTAIL.n329 VTAIL.n296 7.3702
R452 VTAIL.n333 VTAIL.n294 7.3702
R453 VTAIL.n53 VTAIL.n20 7.3702
R454 VTAIL.n57 VTAIL.n18 7.3702
R455 VTAIL.n244 VTAIL.n205 7.3702
R456 VTAIL.n240 VTAIL.n207 7.3702
R457 VTAIL.n152 VTAIL.n113 7.3702
R458 VTAIL.n148 VTAIL.n115 7.3702
R459 VTAIL.n330 VTAIL.n329 6.59444
R460 VTAIL.n330 VTAIL.n294 6.59444
R461 VTAIL.n54 VTAIL.n53 6.59444
R462 VTAIL.n54 VTAIL.n18 6.59444
R463 VTAIL.n241 VTAIL.n205 6.59444
R464 VTAIL.n241 VTAIL.n240 6.59444
R465 VTAIL.n149 VTAIL.n113 6.59444
R466 VTAIL.n149 VTAIL.n148 6.59444
R467 VTAIL.n326 VTAIL.n296 5.81868
R468 VTAIL.n334 VTAIL.n333 5.81868
R469 VTAIL.n50 VTAIL.n20 5.81868
R470 VTAIL.n58 VTAIL.n57 5.81868
R471 VTAIL.n245 VTAIL.n244 5.81868
R472 VTAIL.n237 VTAIL.n207 5.81868
R473 VTAIL.n153 VTAIL.n152 5.81868
R474 VTAIL.n145 VTAIL.n115 5.81868
R475 VTAIL.n325 VTAIL.n298 5.04292
R476 VTAIL.n337 VTAIL.n292 5.04292
R477 VTAIL.n49 VTAIL.n22 5.04292
R478 VTAIL.n61 VTAIL.n16 5.04292
R479 VTAIL.n248 VTAIL.n203 5.04292
R480 VTAIL.n236 VTAIL.n209 5.04292
R481 VTAIL.n156 VTAIL.n111 5.04292
R482 VTAIL.n144 VTAIL.n117 5.04292
R483 VTAIL.n322 VTAIL.n321 4.26717
R484 VTAIL.n338 VTAIL.n290 4.26717
R485 VTAIL.n46 VTAIL.n45 4.26717
R486 VTAIL.n62 VTAIL.n14 4.26717
R487 VTAIL.n249 VTAIL.n201 4.26717
R488 VTAIL.n233 VTAIL.n232 4.26717
R489 VTAIL.n157 VTAIL.n109 4.26717
R490 VTAIL.n141 VTAIL.n140 4.26717
R491 VTAIL.n308 VTAIL.n307 3.70982
R492 VTAIL.n32 VTAIL.n31 3.70982
R493 VTAIL.n219 VTAIL.n218 3.70982
R494 VTAIL.n127 VTAIL.n126 3.70982
R495 VTAIL.n318 VTAIL.n300 3.49141
R496 VTAIL.n342 VTAIL.n341 3.49141
R497 VTAIL.n366 VTAIL.n278 3.49141
R498 VTAIL.n42 VTAIL.n24 3.49141
R499 VTAIL.n66 VTAIL.n65 3.49141
R500 VTAIL.n90 VTAIL.n2 3.49141
R501 VTAIL.n276 VTAIL.n188 3.49141
R502 VTAIL.n253 VTAIL.n252 3.49141
R503 VTAIL.n229 VTAIL.n211 3.49141
R504 VTAIL.n184 VTAIL.n96 3.49141
R505 VTAIL.n161 VTAIL.n160 3.49141
R506 VTAIL.n137 VTAIL.n119 3.49141
R507 VTAIL.n185 VTAIL.n95 3.39705
R508 VTAIL.n277 VTAIL.n187 3.39705
R509 VTAIL.n93 VTAIL.n91 3.39705
R510 VTAIL.n317 VTAIL.n302 2.71565
R511 VTAIL.n345 VTAIL.n288 2.71565
R512 VTAIL.n364 VTAIL.n363 2.71565
R513 VTAIL.n41 VTAIL.n26 2.71565
R514 VTAIL.n69 VTAIL.n12 2.71565
R515 VTAIL.n88 VTAIL.n87 2.71565
R516 VTAIL.n274 VTAIL.n273 2.71565
R517 VTAIL.n256 VTAIL.n199 2.71565
R518 VTAIL.n228 VTAIL.n213 2.71565
R519 VTAIL.n182 VTAIL.n181 2.71565
R520 VTAIL.n164 VTAIL.n107 2.71565
R521 VTAIL.n136 VTAIL.n121 2.71565
R522 VTAIL VTAIL.n367 2.48972
R523 VTAIL.n187 VTAIL.n185 2.1686
R524 VTAIL.n91 VTAIL.n1 2.1686
R525 VTAIL.n0 VTAIL.t1 2.00946
R526 VTAIL.n0 VTAIL.t3 2.00946
R527 VTAIL.n92 VTAIL.t7 2.00946
R528 VTAIL.n92 VTAIL.t8 2.00946
R529 VTAIL.n186 VTAIL.t11 2.00946
R530 VTAIL.n186 VTAIL.t6 2.00946
R531 VTAIL.n94 VTAIL.t5 2.00946
R532 VTAIL.n94 VTAIL.t0 2.00946
R533 VTAIL.n314 VTAIL.n313 1.93989
R534 VTAIL.n346 VTAIL.n286 1.93989
R535 VTAIL.n360 VTAIL.n280 1.93989
R536 VTAIL.n38 VTAIL.n37 1.93989
R537 VTAIL.n70 VTAIL.n10 1.93989
R538 VTAIL.n84 VTAIL.n4 1.93989
R539 VTAIL.n270 VTAIL.n190 1.93989
R540 VTAIL.n257 VTAIL.n197 1.93989
R541 VTAIL.n225 VTAIL.n224 1.93989
R542 VTAIL.n178 VTAIL.n98 1.93989
R543 VTAIL.n165 VTAIL.n105 1.93989
R544 VTAIL.n133 VTAIL.n132 1.93989
R545 VTAIL.n310 VTAIL.n304 1.16414
R546 VTAIL.n351 VTAIL.n349 1.16414
R547 VTAIL.n359 VTAIL.n282 1.16414
R548 VTAIL.n34 VTAIL.n28 1.16414
R549 VTAIL.n75 VTAIL.n73 1.16414
R550 VTAIL.n83 VTAIL.n6 1.16414
R551 VTAIL.n269 VTAIL.n192 1.16414
R552 VTAIL.n261 VTAIL.n260 1.16414
R553 VTAIL.n221 VTAIL.n215 1.16414
R554 VTAIL.n177 VTAIL.n100 1.16414
R555 VTAIL.n169 VTAIL.n168 1.16414
R556 VTAIL.n129 VTAIL.n123 1.16414
R557 VTAIL VTAIL.n1 0.907828
R558 VTAIL.n309 VTAIL.n306 0.388379
R559 VTAIL.n350 VTAIL.n284 0.388379
R560 VTAIL.n356 VTAIL.n355 0.388379
R561 VTAIL.n33 VTAIL.n30 0.388379
R562 VTAIL.n74 VTAIL.n8 0.388379
R563 VTAIL.n80 VTAIL.n79 0.388379
R564 VTAIL.n266 VTAIL.n265 0.388379
R565 VTAIL.n196 VTAIL.n194 0.388379
R566 VTAIL.n220 VTAIL.n217 0.388379
R567 VTAIL.n174 VTAIL.n173 0.388379
R568 VTAIL.n104 VTAIL.n102 0.388379
R569 VTAIL.n128 VTAIL.n125 0.388379
R570 VTAIL.n308 VTAIL.n303 0.155672
R571 VTAIL.n315 VTAIL.n303 0.155672
R572 VTAIL.n316 VTAIL.n315 0.155672
R573 VTAIL.n316 VTAIL.n299 0.155672
R574 VTAIL.n323 VTAIL.n299 0.155672
R575 VTAIL.n324 VTAIL.n323 0.155672
R576 VTAIL.n324 VTAIL.n295 0.155672
R577 VTAIL.n331 VTAIL.n295 0.155672
R578 VTAIL.n332 VTAIL.n331 0.155672
R579 VTAIL.n332 VTAIL.n291 0.155672
R580 VTAIL.n339 VTAIL.n291 0.155672
R581 VTAIL.n340 VTAIL.n339 0.155672
R582 VTAIL.n340 VTAIL.n287 0.155672
R583 VTAIL.n347 VTAIL.n287 0.155672
R584 VTAIL.n348 VTAIL.n347 0.155672
R585 VTAIL.n348 VTAIL.n283 0.155672
R586 VTAIL.n357 VTAIL.n283 0.155672
R587 VTAIL.n358 VTAIL.n357 0.155672
R588 VTAIL.n358 VTAIL.n279 0.155672
R589 VTAIL.n365 VTAIL.n279 0.155672
R590 VTAIL.n32 VTAIL.n27 0.155672
R591 VTAIL.n39 VTAIL.n27 0.155672
R592 VTAIL.n40 VTAIL.n39 0.155672
R593 VTAIL.n40 VTAIL.n23 0.155672
R594 VTAIL.n47 VTAIL.n23 0.155672
R595 VTAIL.n48 VTAIL.n47 0.155672
R596 VTAIL.n48 VTAIL.n19 0.155672
R597 VTAIL.n55 VTAIL.n19 0.155672
R598 VTAIL.n56 VTAIL.n55 0.155672
R599 VTAIL.n56 VTAIL.n15 0.155672
R600 VTAIL.n63 VTAIL.n15 0.155672
R601 VTAIL.n64 VTAIL.n63 0.155672
R602 VTAIL.n64 VTAIL.n11 0.155672
R603 VTAIL.n71 VTAIL.n11 0.155672
R604 VTAIL.n72 VTAIL.n71 0.155672
R605 VTAIL.n72 VTAIL.n7 0.155672
R606 VTAIL.n81 VTAIL.n7 0.155672
R607 VTAIL.n82 VTAIL.n81 0.155672
R608 VTAIL.n82 VTAIL.n3 0.155672
R609 VTAIL.n89 VTAIL.n3 0.155672
R610 VTAIL.n275 VTAIL.n189 0.155672
R611 VTAIL.n268 VTAIL.n189 0.155672
R612 VTAIL.n268 VTAIL.n267 0.155672
R613 VTAIL.n267 VTAIL.n193 0.155672
R614 VTAIL.n259 VTAIL.n193 0.155672
R615 VTAIL.n259 VTAIL.n258 0.155672
R616 VTAIL.n258 VTAIL.n198 0.155672
R617 VTAIL.n251 VTAIL.n198 0.155672
R618 VTAIL.n251 VTAIL.n250 0.155672
R619 VTAIL.n250 VTAIL.n202 0.155672
R620 VTAIL.n243 VTAIL.n202 0.155672
R621 VTAIL.n243 VTAIL.n242 0.155672
R622 VTAIL.n242 VTAIL.n206 0.155672
R623 VTAIL.n235 VTAIL.n206 0.155672
R624 VTAIL.n235 VTAIL.n234 0.155672
R625 VTAIL.n234 VTAIL.n210 0.155672
R626 VTAIL.n227 VTAIL.n210 0.155672
R627 VTAIL.n227 VTAIL.n226 0.155672
R628 VTAIL.n226 VTAIL.n214 0.155672
R629 VTAIL.n219 VTAIL.n214 0.155672
R630 VTAIL.n183 VTAIL.n97 0.155672
R631 VTAIL.n176 VTAIL.n97 0.155672
R632 VTAIL.n176 VTAIL.n175 0.155672
R633 VTAIL.n175 VTAIL.n101 0.155672
R634 VTAIL.n167 VTAIL.n101 0.155672
R635 VTAIL.n167 VTAIL.n166 0.155672
R636 VTAIL.n166 VTAIL.n106 0.155672
R637 VTAIL.n159 VTAIL.n106 0.155672
R638 VTAIL.n159 VTAIL.n158 0.155672
R639 VTAIL.n158 VTAIL.n110 0.155672
R640 VTAIL.n151 VTAIL.n110 0.155672
R641 VTAIL.n151 VTAIL.n150 0.155672
R642 VTAIL.n150 VTAIL.n114 0.155672
R643 VTAIL.n143 VTAIL.n114 0.155672
R644 VTAIL.n143 VTAIL.n142 0.155672
R645 VTAIL.n142 VTAIL.n118 0.155672
R646 VTAIL.n135 VTAIL.n118 0.155672
R647 VTAIL.n135 VTAIL.n134 0.155672
R648 VTAIL.n134 VTAIL.n122 0.155672
R649 VTAIL.n127 VTAIL.n122 0.155672
R650 VDD1.n84 VDD1.n0 756.745
R651 VDD1.n173 VDD1.n89 756.745
R652 VDD1.n85 VDD1.n84 585
R653 VDD1.n83 VDD1.n82 585
R654 VDD1.n4 VDD1.n3 585
R655 VDD1.n77 VDD1.n76 585
R656 VDD1.n75 VDD1.n6 585
R657 VDD1.n74 VDD1.n73 585
R658 VDD1.n9 VDD1.n7 585
R659 VDD1.n68 VDD1.n67 585
R660 VDD1.n66 VDD1.n65 585
R661 VDD1.n13 VDD1.n12 585
R662 VDD1.n60 VDD1.n59 585
R663 VDD1.n58 VDD1.n57 585
R664 VDD1.n17 VDD1.n16 585
R665 VDD1.n52 VDD1.n51 585
R666 VDD1.n50 VDD1.n49 585
R667 VDD1.n21 VDD1.n20 585
R668 VDD1.n44 VDD1.n43 585
R669 VDD1.n42 VDD1.n41 585
R670 VDD1.n25 VDD1.n24 585
R671 VDD1.n36 VDD1.n35 585
R672 VDD1.n34 VDD1.n33 585
R673 VDD1.n29 VDD1.n28 585
R674 VDD1.n117 VDD1.n116 585
R675 VDD1.n122 VDD1.n121 585
R676 VDD1.n124 VDD1.n123 585
R677 VDD1.n113 VDD1.n112 585
R678 VDD1.n130 VDD1.n129 585
R679 VDD1.n132 VDD1.n131 585
R680 VDD1.n109 VDD1.n108 585
R681 VDD1.n138 VDD1.n137 585
R682 VDD1.n140 VDD1.n139 585
R683 VDD1.n105 VDD1.n104 585
R684 VDD1.n146 VDD1.n145 585
R685 VDD1.n148 VDD1.n147 585
R686 VDD1.n101 VDD1.n100 585
R687 VDD1.n154 VDD1.n153 585
R688 VDD1.n156 VDD1.n155 585
R689 VDD1.n97 VDD1.n96 585
R690 VDD1.n163 VDD1.n162 585
R691 VDD1.n164 VDD1.n95 585
R692 VDD1.n166 VDD1.n165 585
R693 VDD1.n93 VDD1.n92 585
R694 VDD1.n172 VDD1.n171 585
R695 VDD1.n174 VDD1.n173 585
R696 VDD1.n30 VDD1.t5 327.466
R697 VDD1.n118 VDD1.t1 327.466
R698 VDD1.n84 VDD1.n83 171.744
R699 VDD1.n83 VDD1.n3 171.744
R700 VDD1.n76 VDD1.n3 171.744
R701 VDD1.n76 VDD1.n75 171.744
R702 VDD1.n75 VDD1.n74 171.744
R703 VDD1.n74 VDD1.n7 171.744
R704 VDD1.n67 VDD1.n7 171.744
R705 VDD1.n67 VDD1.n66 171.744
R706 VDD1.n66 VDD1.n12 171.744
R707 VDD1.n59 VDD1.n12 171.744
R708 VDD1.n59 VDD1.n58 171.744
R709 VDD1.n58 VDD1.n16 171.744
R710 VDD1.n51 VDD1.n16 171.744
R711 VDD1.n51 VDD1.n50 171.744
R712 VDD1.n50 VDD1.n20 171.744
R713 VDD1.n43 VDD1.n20 171.744
R714 VDD1.n43 VDD1.n42 171.744
R715 VDD1.n42 VDD1.n24 171.744
R716 VDD1.n35 VDD1.n24 171.744
R717 VDD1.n35 VDD1.n34 171.744
R718 VDD1.n34 VDD1.n28 171.744
R719 VDD1.n122 VDD1.n116 171.744
R720 VDD1.n123 VDD1.n122 171.744
R721 VDD1.n123 VDD1.n112 171.744
R722 VDD1.n130 VDD1.n112 171.744
R723 VDD1.n131 VDD1.n130 171.744
R724 VDD1.n131 VDD1.n108 171.744
R725 VDD1.n138 VDD1.n108 171.744
R726 VDD1.n139 VDD1.n138 171.744
R727 VDD1.n139 VDD1.n104 171.744
R728 VDD1.n146 VDD1.n104 171.744
R729 VDD1.n147 VDD1.n146 171.744
R730 VDD1.n147 VDD1.n100 171.744
R731 VDD1.n154 VDD1.n100 171.744
R732 VDD1.n155 VDD1.n154 171.744
R733 VDD1.n155 VDD1.n96 171.744
R734 VDD1.n163 VDD1.n96 171.744
R735 VDD1.n164 VDD1.n163 171.744
R736 VDD1.n165 VDD1.n164 171.744
R737 VDD1.n165 VDD1.n92 171.744
R738 VDD1.n172 VDD1.n92 171.744
R739 VDD1.n173 VDD1.n172 171.744
R740 VDD1.t5 VDD1.n28 85.8723
R741 VDD1.t1 VDD1.n116 85.8723
R742 VDD1.n179 VDD1.n178 72.5351
R743 VDD1.n181 VDD1.n180 71.7413
R744 VDD1 VDD1.n88 53.4091
R745 VDD1.n179 VDD1.n177 53.2956
R746 VDD1.n181 VDD1.n179 50.9836
R747 VDD1.n30 VDD1.n29 16.3895
R748 VDD1.n118 VDD1.n117 16.3895
R749 VDD1.n77 VDD1.n6 13.1884
R750 VDD1.n166 VDD1.n95 13.1884
R751 VDD1.n78 VDD1.n4 12.8005
R752 VDD1.n73 VDD1.n8 12.8005
R753 VDD1.n33 VDD1.n32 12.8005
R754 VDD1.n121 VDD1.n120 12.8005
R755 VDD1.n162 VDD1.n161 12.8005
R756 VDD1.n167 VDD1.n93 12.8005
R757 VDD1.n82 VDD1.n81 12.0247
R758 VDD1.n72 VDD1.n9 12.0247
R759 VDD1.n36 VDD1.n27 12.0247
R760 VDD1.n124 VDD1.n115 12.0247
R761 VDD1.n160 VDD1.n97 12.0247
R762 VDD1.n171 VDD1.n170 12.0247
R763 VDD1.n85 VDD1.n2 11.249
R764 VDD1.n69 VDD1.n68 11.249
R765 VDD1.n37 VDD1.n25 11.249
R766 VDD1.n125 VDD1.n113 11.249
R767 VDD1.n157 VDD1.n156 11.249
R768 VDD1.n174 VDD1.n91 11.249
R769 VDD1.n86 VDD1.n0 10.4732
R770 VDD1.n65 VDD1.n11 10.4732
R771 VDD1.n41 VDD1.n40 10.4732
R772 VDD1.n129 VDD1.n128 10.4732
R773 VDD1.n153 VDD1.n99 10.4732
R774 VDD1.n175 VDD1.n89 10.4732
R775 VDD1.n64 VDD1.n13 9.69747
R776 VDD1.n44 VDD1.n23 9.69747
R777 VDD1.n132 VDD1.n111 9.69747
R778 VDD1.n152 VDD1.n101 9.69747
R779 VDD1.n88 VDD1.n87 9.45567
R780 VDD1.n177 VDD1.n176 9.45567
R781 VDD1.n56 VDD1.n55 9.3005
R782 VDD1.n15 VDD1.n14 9.3005
R783 VDD1.n62 VDD1.n61 9.3005
R784 VDD1.n64 VDD1.n63 9.3005
R785 VDD1.n11 VDD1.n10 9.3005
R786 VDD1.n70 VDD1.n69 9.3005
R787 VDD1.n72 VDD1.n71 9.3005
R788 VDD1.n8 VDD1.n5 9.3005
R789 VDD1.n87 VDD1.n86 9.3005
R790 VDD1.n2 VDD1.n1 9.3005
R791 VDD1.n81 VDD1.n80 9.3005
R792 VDD1.n79 VDD1.n78 9.3005
R793 VDD1.n54 VDD1.n53 9.3005
R794 VDD1.n19 VDD1.n18 9.3005
R795 VDD1.n48 VDD1.n47 9.3005
R796 VDD1.n46 VDD1.n45 9.3005
R797 VDD1.n23 VDD1.n22 9.3005
R798 VDD1.n40 VDD1.n39 9.3005
R799 VDD1.n38 VDD1.n37 9.3005
R800 VDD1.n27 VDD1.n26 9.3005
R801 VDD1.n32 VDD1.n31 9.3005
R802 VDD1.n176 VDD1.n175 9.3005
R803 VDD1.n91 VDD1.n90 9.3005
R804 VDD1.n170 VDD1.n169 9.3005
R805 VDD1.n168 VDD1.n167 9.3005
R806 VDD1.n107 VDD1.n106 9.3005
R807 VDD1.n136 VDD1.n135 9.3005
R808 VDD1.n134 VDD1.n133 9.3005
R809 VDD1.n111 VDD1.n110 9.3005
R810 VDD1.n128 VDD1.n127 9.3005
R811 VDD1.n126 VDD1.n125 9.3005
R812 VDD1.n115 VDD1.n114 9.3005
R813 VDD1.n120 VDD1.n119 9.3005
R814 VDD1.n142 VDD1.n141 9.3005
R815 VDD1.n144 VDD1.n143 9.3005
R816 VDD1.n103 VDD1.n102 9.3005
R817 VDD1.n150 VDD1.n149 9.3005
R818 VDD1.n152 VDD1.n151 9.3005
R819 VDD1.n99 VDD1.n98 9.3005
R820 VDD1.n158 VDD1.n157 9.3005
R821 VDD1.n160 VDD1.n159 9.3005
R822 VDD1.n161 VDD1.n94 9.3005
R823 VDD1.n61 VDD1.n60 8.92171
R824 VDD1.n45 VDD1.n21 8.92171
R825 VDD1.n133 VDD1.n109 8.92171
R826 VDD1.n149 VDD1.n148 8.92171
R827 VDD1.n57 VDD1.n15 8.14595
R828 VDD1.n49 VDD1.n48 8.14595
R829 VDD1.n137 VDD1.n136 8.14595
R830 VDD1.n145 VDD1.n103 8.14595
R831 VDD1.n56 VDD1.n17 7.3702
R832 VDD1.n52 VDD1.n19 7.3702
R833 VDD1.n140 VDD1.n107 7.3702
R834 VDD1.n144 VDD1.n105 7.3702
R835 VDD1.n53 VDD1.n17 6.59444
R836 VDD1.n53 VDD1.n52 6.59444
R837 VDD1.n141 VDD1.n140 6.59444
R838 VDD1.n141 VDD1.n105 6.59444
R839 VDD1.n57 VDD1.n56 5.81868
R840 VDD1.n49 VDD1.n19 5.81868
R841 VDD1.n137 VDD1.n107 5.81868
R842 VDD1.n145 VDD1.n144 5.81868
R843 VDD1.n60 VDD1.n15 5.04292
R844 VDD1.n48 VDD1.n21 5.04292
R845 VDD1.n136 VDD1.n109 5.04292
R846 VDD1.n148 VDD1.n103 5.04292
R847 VDD1.n61 VDD1.n13 4.26717
R848 VDD1.n45 VDD1.n44 4.26717
R849 VDD1.n133 VDD1.n132 4.26717
R850 VDD1.n149 VDD1.n101 4.26717
R851 VDD1.n31 VDD1.n30 3.70982
R852 VDD1.n119 VDD1.n118 3.70982
R853 VDD1.n88 VDD1.n0 3.49141
R854 VDD1.n65 VDD1.n64 3.49141
R855 VDD1.n41 VDD1.n23 3.49141
R856 VDD1.n129 VDD1.n111 3.49141
R857 VDD1.n153 VDD1.n152 3.49141
R858 VDD1.n177 VDD1.n89 3.49141
R859 VDD1.n86 VDD1.n85 2.71565
R860 VDD1.n68 VDD1.n11 2.71565
R861 VDD1.n40 VDD1.n25 2.71565
R862 VDD1.n128 VDD1.n113 2.71565
R863 VDD1.n156 VDD1.n99 2.71565
R864 VDD1.n175 VDD1.n174 2.71565
R865 VDD1.n180 VDD1.t3 2.00946
R866 VDD1.n180 VDD1.t0 2.00946
R867 VDD1.n178 VDD1.t2 2.00946
R868 VDD1.n178 VDD1.t4 2.00946
R869 VDD1.n82 VDD1.n2 1.93989
R870 VDD1.n69 VDD1.n9 1.93989
R871 VDD1.n37 VDD1.n36 1.93989
R872 VDD1.n125 VDD1.n124 1.93989
R873 VDD1.n157 VDD1.n97 1.93989
R874 VDD1.n171 VDD1.n91 1.93989
R875 VDD1.n81 VDD1.n4 1.16414
R876 VDD1.n73 VDD1.n72 1.16414
R877 VDD1.n33 VDD1.n27 1.16414
R878 VDD1.n121 VDD1.n115 1.16414
R879 VDD1.n162 VDD1.n160 1.16414
R880 VDD1.n170 VDD1.n93 1.16414
R881 VDD1 VDD1.n181 0.791448
R882 VDD1.n78 VDD1.n77 0.388379
R883 VDD1.n8 VDD1.n6 0.388379
R884 VDD1.n32 VDD1.n29 0.388379
R885 VDD1.n120 VDD1.n117 0.388379
R886 VDD1.n161 VDD1.n95 0.388379
R887 VDD1.n167 VDD1.n166 0.388379
R888 VDD1.n87 VDD1.n1 0.155672
R889 VDD1.n80 VDD1.n1 0.155672
R890 VDD1.n80 VDD1.n79 0.155672
R891 VDD1.n79 VDD1.n5 0.155672
R892 VDD1.n71 VDD1.n5 0.155672
R893 VDD1.n71 VDD1.n70 0.155672
R894 VDD1.n70 VDD1.n10 0.155672
R895 VDD1.n63 VDD1.n10 0.155672
R896 VDD1.n63 VDD1.n62 0.155672
R897 VDD1.n62 VDD1.n14 0.155672
R898 VDD1.n55 VDD1.n14 0.155672
R899 VDD1.n55 VDD1.n54 0.155672
R900 VDD1.n54 VDD1.n18 0.155672
R901 VDD1.n47 VDD1.n18 0.155672
R902 VDD1.n47 VDD1.n46 0.155672
R903 VDD1.n46 VDD1.n22 0.155672
R904 VDD1.n39 VDD1.n22 0.155672
R905 VDD1.n39 VDD1.n38 0.155672
R906 VDD1.n38 VDD1.n26 0.155672
R907 VDD1.n31 VDD1.n26 0.155672
R908 VDD1.n119 VDD1.n114 0.155672
R909 VDD1.n126 VDD1.n114 0.155672
R910 VDD1.n127 VDD1.n126 0.155672
R911 VDD1.n127 VDD1.n110 0.155672
R912 VDD1.n134 VDD1.n110 0.155672
R913 VDD1.n135 VDD1.n134 0.155672
R914 VDD1.n135 VDD1.n106 0.155672
R915 VDD1.n142 VDD1.n106 0.155672
R916 VDD1.n143 VDD1.n142 0.155672
R917 VDD1.n143 VDD1.n102 0.155672
R918 VDD1.n150 VDD1.n102 0.155672
R919 VDD1.n151 VDD1.n150 0.155672
R920 VDD1.n151 VDD1.n98 0.155672
R921 VDD1.n158 VDD1.n98 0.155672
R922 VDD1.n159 VDD1.n158 0.155672
R923 VDD1.n159 VDD1.n94 0.155672
R924 VDD1.n168 VDD1.n94 0.155672
R925 VDD1.n169 VDD1.n168 0.155672
R926 VDD1.n169 VDD1.n90 0.155672
R927 VDD1.n176 VDD1.n90 0.155672
R928 VN.n38 VN.n37 161.3
R929 VN.n36 VN.n21 161.3
R930 VN.n35 VN.n34 161.3
R931 VN.n33 VN.n22 161.3
R932 VN.n32 VN.n31 161.3
R933 VN.n30 VN.n23 161.3
R934 VN.n29 VN.n28 161.3
R935 VN.n27 VN.n24 161.3
R936 VN.n18 VN.n17 161.3
R937 VN.n16 VN.n1 161.3
R938 VN.n15 VN.n14 161.3
R939 VN.n13 VN.n2 161.3
R940 VN.n12 VN.n11 161.3
R941 VN.n10 VN.n3 161.3
R942 VN.n9 VN.n8 161.3
R943 VN.n7 VN.n4 161.3
R944 VN.n26 VN.t2 141.381
R945 VN.n6 VN.t5 141.381
R946 VN.n5 VN.t0 108.016
R947 VN.n0 VN.t1 108.016
R948 VN.n25 VN.t4 108.016
R949 VN.n20 VN.t3 108.016
R950 VN.n19 VN.n0 80.9007
R951 VN.n39 VN.n20 80.9007
R952 VN.n6 VN.n5 62.5184
R953 VN.n26 VN.n25 62.5184
R954 VN.n11 VN.n2 56.5617
R955 VN.n31 VN.n22 56.5617
R956 VN VN.n39 56.0739
R957 VN.n9 VN.n4 24.5923
R958 VN.n10 VN.n9 24.5923
R959 VN.n11 VN.n10 24.5923
R960 VN.n15 VN.n2 24.5923
R961 VN.n16 VN.n15 24.5923
R962 VN.n17 VN.n16 24.5923
R963 VN.n31 VN.n30 24.5923
R964 VN.n30 VN.n29 24.5923
R965 VN.n29 VN.n24 24.5923
R966 VN.n37 VN.n36 24.5923
R967 VN.n36 VN.n35 24.5923
R968 VN.n35 VN.n22 24.5923
R969 VN.n5 VN.n4 12.2964
R970 VN.n25 VN.n24 12.2964
R971 VN.n17 VN.n0 9.3454
R972 VN.n37 VN.n20 9.3454
R973 VN.n27 VN.n26 3.16706
R974 VN.n7 VN.n6 3.16706
R975 VN.n39 VN.n38 0.354861
R976 VN.n19 VN.n18 0.354861
R977 VN VN.n19 0.267071
R978 VN.n38 VN.n21 0.189894
R979 VN.n34 VN.n21 0.189894
R980 VN.n34 VN.n33 0.189894
R981 VN.n33 VN.n32 0.189894
R982 VN.n32 VN.n23 0.189894
R983 VN.n28 VN.n23 0.189894
R984 VN.n28 VN.n27 0.189894
R985 VN.n8 VN.n7 0.189894
R986 VN.n8 VN.n3 0.189894
R987 VN.n12 VN.n3 0.189894
R988 VN.n13 VN.n12 0.189894
R989 VN.n14 VN.n13 0.189894
R990 VN.n14 VN.n1 0.189894
R991 VN.n18 VN.n1 0.189894
R992 VDD2.n175 VDD2.n91 756.745
R993 VDD2.n84 VDD2.n0 756.745
R994 VDD2.n176 VDD2.n175 585
R995 VDD2.n174 VDD2.n173 585
R996 VDD2.n95 VDD2.n94 585
R997 VDD2.n168 VDD2.n167 585
R998 VDD2.n166 VDD2.n97 585
R999 VDD2.n165 VDD2.n164 585
R1000 VDD2.n100 VDD2.n98 585
R1001 VDD2.n159 VDD2.n158 585
R1002 VDD2.n157 VDD2.n156 585
R1003 VDD2.n104 VDD2.n103 585
R1004 VDD2.n151 VDD2.n150 585
R1005 VDD2.n149 VDD2.n148 585
R1006 VDD2.n108 VDD2.n107 585
R1007 VDD2.n143 VDD2.n142 585
R1008 VDD2.n141 VDD2.n140 585
R1009 VDD2.n112 VDD2.n111 585
R1010 VDD2.n135 VDD2.n134 585
R1011 VDD2.n133 VDD2.n132 585
R1012 VDD2.n116 VDD2.n115 585
R1013 VDD2.n127 VDD2.n126 585
R1014 VDD2.n125 VDD2.n124 585
R1015 VDD2.n120 VDD2.n119 585
R1016 VDD2.n28 VDD2.n27 585
R1017 VDD2.n33 VDD2.n32 585
R1018 VDD2.n35 VDD2.n34 585
R1019 VDD2.n24 VDD2.n23 585
R1020 VDD2.n41 VDD2.n40 585
R1021 VDD2.n43 VDD2.n42 585
R1022 VDD2.n20 VDD2.n19 585
R1023 VDD2.n49 VDD2.n48 585
R1024 VDD2.n51 VDD2.n50 585
R1025 VDD2.n16 VDD2.n15 585
R1026 VDD2.n57 VDD2.n56 585
R1027 VDD2.n59 VDD2.n58 585
R1028 VDD2.n12 VDD2.n11 585
R1029 VDD2.n65 VDD2.n64 585
R1030 VDD2.n67 VDD2.n66 585
R1031 VDD2.n8 VDD2.n7 585
R1032 VDD2.n74 VDD2.n73 585
R1033 VDD2.n75 VDD2.n6 585
R1034 VDD2.n77 VDD2.n76 585
R1035 VDD2.n4 VDD2.n3 585
R1036 VDD2.n83 VDD2.n82 585
R1037 VDD2.n85 VDD2.n84 585
R1038 VDD2.n121 VDD2.t2 327.466
R1039 VDD2.n29 VDD2.t0 327.466
R1040 VDD2.n175 VDD2.n174 171.744
R1041 VDD2.n174 VDD2.n94 171.744
R1042 VDD2.n167 VDD2.n94 171.744
R1043 VDD2.n167 VDD2.n166 171.744
R1044 VDD2.n166 VDD2.n165 171.744
R1045 VDD2.n165 VDD2.n98 171.744
R1046 VDD2.n158 VDD2.n98 171.744
R1047 VDD2.n158 VDD2.n157 171.744
R1048 VDD2.n157 VDD2.n103 171.744
R1049 VDD2.n150 VDD2.n103 171.744
R1050 VDD2.n150 VDD2.n149 171.744
R1051 VDD2.n149 VDD2.n107 171.744
R1052 VDD2.n142 VDD2.n107 171.744
R1053 VDD2.n142 VDD2.n141 171.744
R1054 VDD2.n141 VDD2.n111 171.744
R1055 VDD2.n134 VDD2.n111 171.744
R1056 VDD2.n134 VDD2.n133 171.744
R1057 VDD2.n133 VDD2.n115 171.744
R1058 VDD2.n126 VDD2.n115 171.744
R1059 VDD2.n126 VDD2.n125 171.744
R1060 VDD2.n125 VDD2.n119 171.744
R1061 VDD2.n33 VDD2.n27 171.744
R1062 VDD2.n34 VDD2.n33 171.744
R1063 VDD2.n34 VDD2.n23 171.744
R1064 VDD2.n41 VDD2.n23 171.744
R1065 VDD2.n42 VDD2.n41 171.744
R1066 VDD2.n42 VDD2.n19 171.744
R1067 VDD2.n49 VDD2.n19 171.744
R1068 VDD2.n50 VDD2.n49 171.744
R1069 VDD2.n50 VDD2.n15 171.744
R1070 VDD2.n57 VDD2.n15 171.744
R1071 VDD2.n58 VDD2.n57 171.744
R1072 VDD2.n58 VDD2.n11 171.744
R1073 VDD2.n65 VDD2.n11 171.744
R1074 VDD2.n66 VDD2.n65 171.744
R1075 VDD2.n66 VDD2.n7 171.744
R1076 VDD2.n74 VDD2.n7 171.744
R1077 VDD2.n75 VDD2.n74 171.744
R1078 VDD2.n76 VDD2.n75 171.744
R1079 VDD2.n76 VDD2.n3 171.744
R1080 VDD2.n83 VDD2.n3 171.744
R1081 VDD2.n84 VDD2.n83 171.744
R1082 VDD2.t2 VDD2.n119 85.8723
R1083 VDD2.t0 VDD2.n27 85.8723
R1084 VDD2.n90 VDD2.n89 72.5351
R1085 VDD2 VDD2.n181 72.5323
R1086 VDD2.n90 VDD2.n88 53.2956
R1087 VDD2.n180 VDD2.n179 50.8035
R1088 VDD2.n180 VDD2.n90 48.7024
R1089 VDD2.n121 VDD2.n120 16.3895
R1090 VDD2.n29 VDD2.n28 16.3895
R1091 VDD2.n168 VDD2.n97 13.1884
R1092 VDD2.n77 VDD2.n6 13.1884
R1093 VDD2.n169 VDD2.n95 12.8005
R1094 VDD2.n164 VDD2.n99 12.8005
R1095 VDD2.n124 VDD2.n123 12.8005
R1096 VDD2.n32 VDD2.n31 12.8005
R1097 VDD2.n73 VDD2.n72 12.8005
R1098 VDD2.n78 VDD2.n4 12.8005
R1099 VDD2.n173 VDD2.n172 12.0247
R1100 VDD2.n163 VDD2.n100 12.0247
R1101 VDD2.n127 VDD2.n118 12.0247
R1102 VDD2.n35 VDD2.n26 12.0247
R1103 VDD2.n71 VDD2.n8 12.0247
R1104 VDD2.n82 VDD2.n81 12.0247
R1105 VDD2.n176 VDD2.n93 11.249
R1106 VDD2.n160 VDD2.n159 11.249
R1107 VDD2.n128 VDD2.n116 11.249
R1108 VDD2.n36 VDD2.n24 11.249
R1109 VDD2.n68 VDD2.n67 11.249
R1110 VDD2.n85 VDD2.n2 11.249
R1111 VDD2.n177 VDD2.n91 10.4732
R1112 VDD2.n156 VDD2.n102 10.4732
R1113 VDD2.n132 VDD2.n131 10.4732
R1114 VDD2.n40 VDD2.n39 10.4732
R1115 VDD2.n64 VDD2.n10 10.4732
R1116 VDD2.n86 VDD2.n0 10.4732
R1117 VDD2.n155 VDD2.n104 9.69747
R1118 VDD2.n135 VDD2.n114 9.69747
R1119 VDD2.n43 VDD2.n22 9.69747
R1120 VDD2.n63 VDD2.n12 9.69747
R1121 VDD2.n179 VDD2.n178 9.45567
R1122 VDD2.n88 VDD2.n87 9.45567
R1123 VDD2.n147 VDD2.n146 9.3005
R1124 VDD2.n106 VDD2.n105 9.3005
R1125 VDD2.n153 VDD2.n152 9.3005
R1126 VDD2.n155 VDD2.n154 9.3005
R1127 VDD2.n102 VDD2.n101 9.3005
R1128 VDD2.n161 VDD2.n160 9.3005
R1129 VDD2.n163 VDD2.n162 9.3005
R1130 VDD2.n99 VDD2.n96 9.3005
R1131 VDD2.n178 VDD2.n177 9.3005
R1132 VDD2.n93 VDD2.n92 9.3005
R1133 VDD2.n172 VDD2.n171 9.3005
R1134 VDD2.n170 VDD2.n169 9.3005
R1135 VDD2.n145 VDD2.n144 9.3005
R1136 VDD2.n110 VDD2.n109 9.3005
R1137 VDD2.n139 VDD2.n138 9.3005
R1138 VDD2.n137 VDD2.n136 9.3005
R1139 VDD2.n114 VDD2.n113 9.3005
R1140 VDD2.n131 VDD2.n130 9.3005
R1141 VDD2.n129 VDD2.n128 9.3005
R1142 VDD2.n118 VDD2.n117 9.3005
R1143 VDD2.n123 VDD2.n122 9.3005
R1144 VDD2.n87 VDD2.n86 9.3005
R1145 VDD2.n2 VDD2.n1 9.3005
R1146 VDD2.n81 VDD2.n80 9.3005
R1147 VDD2.n79 VDD2.n78 9.3005
R1148 VDD2.n18 VDD2.n17 9.3005
R1149 VDD2.n47 VDD2.n46 9.3005
R1150 VDD2.n45 VDD2.n44 9.3005
R1151 VDD2.n22 VDD2.n21 9.3005
R1152 VDD2.n39 VDD2.n38 9.3005
R1153 VDD2.n37 VDD2.n36 9.3005
R1154 VDD2.n26 VDD2.n25 9.3005
R1155 VDD2.n31 VDD2.n30 9.3005
R1156 VDD2.n53 VDD2.n52 9.3005
R1157 VDD2.n55 VDD2.n54 9.3005
R1158 VDD2.n14 VDD2.n13 9.3005
R1159 VDD2.n61 VDD2.n60 9.3005
R1160 VDD2.n63 VDD2.n62 9.3005
R1161 VDD2.n10 VDD2.n9 9.3005
R1162 VDD2.n69 VDD2.n68 9.3005
R1163 VDD2.n71 VDD2.n70 9.3005
R1164 VDD2.n72 VDD2.n5 9.3005
R1165 VDD2.n152 VDD2.n151 8.92171
R1166 VDD2.n136 VDD2.n112 8.92171
R1167 VDD2.n44 VDD2.n20 8.92171
R1168 VDD2.n60 VDD2.n59 8.92171
R1169 VDD2.n148 VDD2.n106 8.14595
R1170 VDD2.n140 VDD2.n139 8.14595
R1171 VDD2.n48 VDD2.n47 8.14595
R1172 VDD2.n56 VDD2.n14 8.14595
R1173 VDD2.n147 VDD2.n108 7.3702
R1174 VDD2.n143 VDD2.n110 7.3702
R1175 VDD2.n51 VDD2.n18 7.3702
R1176 VDD2.n55 VDD2.n16 7.3702
R1177 VDD2.n144 VDD2.n108 6.59444
R1178 VDD2.n144 VDD2.n143 6.59444
R1179 VDD2.n52 VDD2.n51 6.59444
R1180 VDD2.n52 VDD2.n16 6.59444
R1181 VDD2.n148 VDD2.n147 5.81868
R1182 VDD2.n140 VDD2.n110 5.81868
R1183 VDD2.n48 VDD2.n18 5.81868
R1184 VDD2.n56 VDD2.n55 5.81868
R1185 VDD2.n151 VDD2.n106 5.04292
R1186 VDD2.n139 VDD2.n112 5.04292
R1187 VDD2.n47 VDD2.n20 5.04292
R1188 VDD2.n59 VDD2.n14 5.04292
R1189 VDD2.n152 VDD2.n104 4.26717
R1190 VDD2.n136 VDD2.n135 4.26717
R1191 VDD2.n44 VDD2.n43 4.26717
R1192 VDD2.n60 VDD2.n12 4.26717
R1193 VDD2.n122 VDD2.n121 3.70982
R1194 VDD2.n30 VDD2.n29 3.70982
R1195 VDD2.n179 VDD2.n91 3.49141
R1196 VDD2.n156 VDD2.n155 3.49141
R1197 VDD2.n132 VDD2.n114 3.49141
R1198 VDD2.n40 VDD2.n22 3.49141
R1199 VDD2.n64 VDD2.n63 3.49141
R1200 VDD2.n88 VDD2.n0 3.49141
R1201 VDD2.n177 VDD2.n176 2.71565
R1202 VDD2.n159 VDD2.n102 2.71565
R1203 VDD2.n131 VDD2.n116 2.71565
R1204 VDD2.n39 VDD2.n24 2.71565
R1205 VDD2.n67 VDD2.n10 2.71565
R1206 VDD2.n86 VDD2.n85 2.71565
R1207 VDD2 VDD2.n180 2.6061
R1208 VDD2.n181 VDD2.t1 2.00946
R1209 VDD2.n181 VDD2.t3 2.00946
R1210 VDD2.n89 VDD2.t5 2.00946
R1211 VDD2.n89 VDD2.t4 2.00946
R1212 VDD2.n173 VDD2.n93 1.93989
R1213 VDD2.n160 VDD2.n100 1.93989
R1214 VDD2.n128 VDD2.n127 1.93989
R1215 VDD2.n36 VDD2.n35 1.93989
R1216 VDD2.n68 VDD2.n8 1.93989
R1217 VDD2.n82 VDD2.n2 1.93989
R1218 VDD2.n172 VDD2.n95 1.16414
R1219 VDD2.n164 VDD2.n163 1.16414
R1220 VDD2.n124 VDD2.n118 1.16414
R1221 VDD2.n32 VDD2.n26 1.16414
R1222 VDD2.n73 VDD2.n71 1.16414
R1223 VDD2.n81 VDD2.n4 1.16414
R1224 VDD2.n169 VDD2.n168 0.388379
R1225 VDD2.n99 VDD2.n97 0.388379
R1226 VDD2.n123 VDD2.n120 0.388379
R1227 VDD2.n31 VDD2.n28 0.388379
R1228 VDD2.n72 VDD2.n6 0.388379
R1229 VDD2.n78 VDD2.n77 0.388379
R1230 VDD2.n178 VDD2.n92 0.155672
R1231 VDD2.n171 VDD2.n92 0.155672
R1232 VDD2.n171 VDD2.n170 0.155672
R1233 VDD2.n170 VDD2.n96 0.155672
R1234 VDD2.n162 VDD2.n96 0.155672
R1235 VDD2.n162 VDD2.n161 0.155672
R1236 VDD2.n161 VDD2.n101 0.155672
R1237 VDD2.n154 VDD2.n101 0.155672
R1238 VDD2.n154 VDD2.n153 0.155672
R1239 VDD2.n153 VDD2.n105 0.155672
R1240 VDD2.n146 VDD2.n105 0.155672
R1241 VDD2.n146 VDD2.n145 0.155672
R1242 VDD2.n145 VDD2.n109 0.155672
R1243 VDD2.n138 VDD2.n109 0.155672
R1244 VDD2.n138 VDD2.n137 0.155672
R1245 VDD2.n137 VDD2.n113 0.155672
R1246 VDD2.n130 VDD2.n113 0.155672
R1247 VDD2.n130 VDD2.n129 0.155672
R1248 VDD2.n129 VDD2.n117 0.155672
R1249 VDD2.n122 VDD2.n117 0.155672
R1250 VDD2.n30 VDD2.n25 0.155672
R1251 VDD2.n37 VDD2.n25 0.155672
R1252 VDD2.n38 VDD2.n37 0.155672
R1253 VDD2.n38 VDD2.n21 0.155672
R1254 VDD2.n45 VDD2.n21 0.155672
R1255 VDD2.n46 VDD2.n45 0.155672
R1256 VDD2.n46 VDD2.n17 0.155672
R1257 VDD2.n53 VDD2.n17 0.155672
R1258 VDD2.n54 VDD2.n53 0.155672
R1259 VDD2.n54 VDD2.n13 0.155672
R1260 VDD2.n61 VDD2.n13 0.155672
R1261 VDD2.n62 VDD2.n61 0.155672
R1262 VDD2.n62 VDD2.n9 0.155672
R1263 VDD2.n69 VDD2.n9 0.155672
R1264 VDD2.n70 VDD2.n69 0.155672
R1265 VDD2.n70 VDD2.n5 0.155672
R1266 VDD2.n79 VDD2.n5 0.155672
R1267 VDD2.n80 VDD2.n79 0.155672
R1268 VDD2.n80 VDD2.n1 0.155672
R1269 VDD2.n87 VDD2.n1 0.155672
R1270 B.n492 B.n147 585
R1271 B.n491 B.n490 585
R1272 B.n489 B.n148 585
R1273 B.n488 B.n487 585
R1274 B.n486 B.n149 585
R1275 B.n485 B.n484 585
R1276 B.n483 B.n150 585
R1277 B.n482 B.n481 585
R1278 B.n480 B.n151 585
R1279 B.n479 B.n478 585
R1280 B.n477 B.n152 585
R1281 B.n476 B.n475 585
R1282 B.n474 B.n153 585
R1283 B.n473 B.n472 585
R1284 B.n471 B.n154 585
R1285 B.n470 B.n469 585
R1286 B.n468 B.n155 585
R1287 B.n467 B.n466 585
R1288 B.n465 B.n156 585
R1289 B.n464 B.n463 585
R1290 B.n462 B.n157 585
R1291 B.n461 B.n460 585
R1292 B.n459 B.n158 585
R1293 B.n458 B.n457 585
R1294 B.n456 B.n159 585
R1295 B.n455 B.n454 585
R1296 B.n453 B.n160 585
R1297 B.n452 B.n451 585
R1298 B.n450 B.n161 585
R1299 B.n449 B.n448 585
R1300 B.n447 B.n162 585
R1301 B.n446 B.n445 585
R1302 B.n444 B.n163 585
R1303 B.n443 B.n442 585
R1304 B.n441 B.n164 585
R1305 B.n440 B.n439 585
R1306 B.n438 B.n165 585
R1307 B.n437 B.n436 585
R1308 B.n435 B.n166 585
R1309 B.n434 B.n433 585
R1310 B.n432 B.n167 585
R1311 B.n431 B.n430 585
R1312 B.n429 B.n168 585
R1313 B.n428 B.n427 585
R1314 B.n426 B.n169 585
R1315 B.n425 B.n424 585
R1316 B.n423 B.n170 585
R1317 B.n422 B.n421 585
R1318 B.n420 B.n171 585
R1319 B.n419 B.n418 585
R1320 B.n417 B.n172 585
R1321 B.n416 B.n415 585
R1322 B.n414 B.n173 585
R1323 B.n413 B.n412 585
R1324 B.n411 B.n410 585
R1325 B.n409 B.n177 585
R1326 B.n408 B.n407 585
R1327 B.n406 B.n178 585
R1328 B.n405 B.n404 585
R1329 B.n403 B.n179 585
R1330 B.n402 B.n401 585
R1331 B.n400 B.n180 585
R1332 B.n399 B.n398 585
R1333 B.n396 B.n181 585
R1334 B.n395 B.n394 585
R1335 B.n393 B.n184 585
R1336 B.n392 B.n391 585
R1337 B.n390 B.n185 585
R1338 B.n389 B.n388 585
R1339 B.n387 B.n186 585
R1340 B.n386 B.n385 585
R1341 B.n384 B.n187 585
R1342 B.n383 B.n382 585
R1343 B.n381 B.n188 585
R1344 B.n380 B.n379 585
R1345 B.n378 B.n189 585
R1346 B.n377 B.n376 585
R1347 B.n375 B.n190 585
R1348 B.n374 B.n373 585
R1349 B.n372 B.n191 585
R1350 B.n371 B.n370 585
R1351 B.n369 B.n192 585
R1352 B.n368 B.n367 585
R1353 B.n366 B.n193 585
R1354 B.n365 B.n364 585
R1355 B.n363 B.n194 585
R1356 B.n362 B.n361 585
R1357 B.n360 B.n195 585
R1358 B.n359 B.n358 585
R1359 B.n357 B.n196 585
R1360 B.n356 B.n355 585
R1361 B.n354 B.n197 585
R1362 B.n353 B.n352 585
R1363 B.n351 B.n198 585
R1364 B.n350 B.n349 585
R1365 B.n348 B.n199 585
R1366 B.n347 B.n346 585
R1367 B.n345 B.n200 585
R1368 B.n344 B.n343 585
R1369 B.n342 B.n201 585
R1370 B.n341 B.n340 585
R1371 B.n339 B.n202 585
R1372 B.n338 B.n337 585
R1373 B.n336 B.n203 585
R1374 B.n335 B.n334 585
R1375 B.n333 B.n204 585
R1376 B.n332 B.n331 585
R1377 B.n330 B.n205 585
R1378 B.n329 B.n328 585
R1379 B.n327 B.n206 585
R1380 B.n326 B.n325 585
R1381 B.n324 B.n207 585
R1382 B.n323 B.n322 585
R1383 B.n321 B.n208 585
R1384 B.n320 B.n319 585
R1385 B.n318 B.n209 585
R1386 B.n317 B.n316 585
R1387 B.n494 B.n493 585
R1388 B.n495 B.n146 585
R1389 B.n497 B.n496 585
R1390 B.n498 B.n145 585
R1391 B.n500 B.n499 585
R1392 B.n501 B.n144 585
R1393 B.n503 B.n502 585
R1394 B.n504 B.n143 585
R1395 B.n506 B.n505 585
R1396 B.n507 B.n142 585
R1397 B.n509 B.n508 585
R1398 B.n510 B.n141 585
R1399 B.n512 B.n511 585
R1400 B.n513 B.n140 585
R1401 B.n515 B.n514 585
R1402 B.n516 B.n139 585
R1403 B.n518 B.n517 585
R1404 B.n519 B.n138 585
R1405 B.n521 B.n520 585
R1406 B.n522 B.n137 585
R1407 B.n524 B.n523 585
R1408 B.n525 B.n136 585
R1409 B.n527 B.n526 585
R1410 B.n528 B.n135 585
R1411 B.n530 B.n529 585
R1412 B.n531 B.n134 585
R1413 B.n533 B.n532 585
R1414 B.n534 B.n133 585
R1415 B.n536 B.n535 585
R1416 B.n537 B.n132 585
R1417 B.n539 B.n538 585
R1418 B.n540 B.n131 585
R1419 B.n542 B.n541 585
R1420 B.n543 B.n130 585
R1421 B.n545 B.n544 585
R1422 B.n546 B.n129 585
R1423 B.n548 B.n547 585
R1424 B.n549 B.n128 585
R1425 B.n551 B.n550 585
R1426 B.n552 B.n127 585
R1427 B.n554 B.n553 585
R1428 B.n555 B.n126 585
R1429 B.n557 B.n556 585
R1430 B.n558 B.n125 585
R1431 B.n560 B.n559 585
R1432 B.n561 B.n124 585
R1433 B.n563 B.n562 585
R1434 B.n564 B.n123 585
R1435 B.n566 B.n565 585
R1436 B.n567 B.n122 585
R1437 B.n569 B.n568 585
R1438 B.n570 B.n121 585
R1439 B.n572 B.n571 585
R1440 B.n573 B.n120 585
R1441 B.n575 B.n574 585
R1442 B.n576 B.n119 585
R1443 B.n578 B.n577 585
R1444 B.n579 B.n118 585
R1445 B.n581 B.n580 585
R1446 B.n582 B.n117 585
R1447 B.n584 B.n583 585
R1448 B.n585 B.n116 585
R1449 B.n587 B.n586 585
R1450 B.n588 B.n115 585
R1451 B.n590 B.n589 585
R1452 B.n591 B.n114 585
R1453 B.n593 B.n592 585
R1454 B.n594 B.n113 585
R1455 B.n596 B.n595 585
R1456 B.n597 B.n112 585
R1457 B.n599 B.n598 585
R1458 B.n600 B.n111 585
R1459 B.n602 B.n601 585
R1460 B.n603 B.n110 585
R1461 B.n605 B.n604 585
R1462 B.n606 B.n109 585
R1463 B.n608 B.n607 585
R1464 B.n609 B.n108 585
R1465 B.n611 B.n610 585
R1466 B.n612 B.n107 585
R1467 B.n614 B.n613 585
R1468 B.n615 B.n106 585
R1469 B.n617 B.n616 585
R1470 B.n618 B.n105 585
R1471 B.n620 B.n619 585
R1472 B.n621 B.n104 585
R1473 B.n623 B.n622 585
R1474 B.n624 B.n103 585
R1475 B.n626 B.n625 585
R1476 B.n627 B.n102 585
R1477 B.n629 B.n628 585
R1478 B.n630 B.n101 585
R1479 B.n632 B.n631 585
R1480 B.n633 B.n100 585
R1481 B.n635 B.n634 585
R1482 B.n636 B.n99 585
R1483 B.n638 B.n637 585
R1484 B.n639 B.n98 585
R1485 B.n641 B.n640 585
R1486 B.n642 B.n97 585
R1487 B.n644 B.n643 585
R1488 B.n645 B.n96 585
R1489 B.n647 B.n646 585
R1490 B.n648 B.n95 585
R1491 B.n650 B.n649 585
R1492 B.n651 B.n94 585
R1493 B.n653 B.n652 585
R1494 B.n654 B.n93 585
R1495 B.n656 B.n655 585
R1496 B.n657 B.n92 585
R1497 B.n834 B.n29 585
R1498 B.n833 B.n832 585
R1499 B.n831 B.n30 585
R1500 B.n830 B.n829 585
R1501 B.n828 B.n31 585
R1502 B.n827 B.n826 585
R1503 B.n825 B.n32 585
R1504 B.n824 B.n823 585
R1505 B.n822 B.n33 585
R1506 B.n821 B.n820 585
R1507 B.n819 B.n34 585
R1508 B.n818 B.n817 585
R1509 B.n816 B.n35 585
R1510 B.n815 B.n814 585
R1511 B.n813 B.n36 585
R1512 B.n812 B.n811 585
R1513 B.n810 B.n37 585
R1514 B.n809 B.n808 585
R1515 B.n807 B.n38 585
R1516 B.n806 B.n805 585
R1517 B.n804 B.n39 585
R1518 B.n803 B.n802 585
R1519 B.n801 B.n40 585
R1520 B.n800 B.n799 585
R1521 B.n798 B.n41 585
R1522 B.n797 B.n796 585
R1523 B.n795 B.n42 585
R1524 B.n794 B.n793 585
R1525 B.n792 B.n43 585
R1526 B.n791 B.n790 585
R1527 B.n789 B.n44 585
R1528 B.n788 B.n787 585
R1529 B.n786 B.n45 585
R1530 B.n785 B.n784 585
R1531 B.n783 B.n46 585
R1532 B.n782 B.n781 585
R1533 B.n780 B.n47 585
R1534 B.n779 B.n778 585
R1535 B.n777 B.n48 585
R1536 B.n776 B.n775 585
R1537 B.n774 B.n49 585
R1538 B.n773 B.n772 585
R1539 B.n771 B.n50 585
R1540 B.n770 B.n769 585
R1541 B.n768 B.n51 585
R1542 B.n767 B.n766 585
R1543 B.n765 B.n52 585
R1544 B.n764 B.n763 585
R1545 B.n762 B.n53 585
R1546 B.n761 B.n760 585
R1547 B.n759 B.n54 585
R1548 B.n758 B.n757 585
R1549 B.n756 B.n55 585
R1550 B.n755 B.n754 585
R1551 B.n753 B.n752 585
R1552 B.n751 B.n59 585
R1553 B.n750 B.n749 585
R1554 B.n748 B.n60 585
R1555 B.n747 B.n746 585
R1556 B.n745 B.n61 585
R1557 B.n744 B.n743 585
R1558 B.n742 B.n62 585
R1559 B.n741 B.n740 585
R1560 B.n738 B.n63 585
R1561 B.n737 B.n736 585
R1562 B.n735 B.n66 585
R1563 B.n734 B.n733 585
R1564 B.n732 B.n67 585
R1565 B.n731 B.n730 585
R1566 B.n729 B.n68 585
R1567 B.n728 B.n727 585
R1568 B.n726 B.n69 585
R1569 B.n725 B.n724 585
R1570 B.n723 B.n70 585
R1571 B.n722 B.n721 585
R1572 B.n720 B.n71 585
R1573 B.n719 B.n718 585
R1574 B.n717 B.n72 585
R1575 B.n716 B.n715 585
R1576 B.n714 B.n73 585
R1577 B.n713 B.n712 585
R1578 B.n711 B.n74 585
R1579 B.n710 B.n709 585
R1580 B.n708 B.n75 585
R1581 B.n707 B.n706 585
R1582 B.n705 B.n76 585
R1583 B.n704 B.n703 585
R1584 B.n702 B.n77 585
R1585 B.n701 B.n700 585
R1586 B.n699 B.n78 585
R1587 B.n698 B.n697 585
R1588 B.n696 B.n79 585
R1589 B.n695 B.n694 585
R1590 B.n693 B.n80 585
R1591 B.n692 B.n691 585
R1592 B.n690 B.n81 585
R1593 B.n689 B.n688 585
R1594 B.n687 B.n82 585
R1595 B.n686 B.n685 585
R1596 B.n684 B.n83 585
R1597 B.n683 B.n682 585
R1598 B.n681 B.n84 585
R1599 B.n680 B.n679 585
R1600 B.n678 B.n85 585
R1601 B.n677 B.n676 585
R1602 B.n675 B.n86 585
R1603 B.n674 B.n673 585
R1604 B.n672 B.n87 585
R1605 B.n671 B.n670 585
R1606 B.n669 B.n88 585
R1607 B.n668 B.n667 585
R1608 B.n666 B.n89 585
R1609 B.n665 B.n664 585
R1610 B.n663 B.n90 585
R1611 B.n662 B.n661 585
R1612 B.n660 B.n91 585
R1613 B.n659 B.n658 585
R1614 B.n836 B.n835 585
R1615 B.n837 B.n28 585
R1616 B.n839 B.n838 585
R1617 B.n840 B.n27 585
R1618 B.n842 B.n841 585
R1619 B.n843 B.n26 585
R1620 B.n845 B.n844 585
R1621 B.n846 B.n25 585
R1622 B.n848 B.n847 585
R1623 B.n849 B.n24 585
R1624 B.n851 B.n850 585
R1625 B.n852 B.n23 585
R1626 B.n854 B.n853 585
R1627 B.n855 B.n22 585
R1628 B.n857 B.n856 585
R1629 B.n858 B.n21 585
R1630 B.n860 B.n859 585
R1631 B.n861 B.n20 585
R1632 B.n863 B.n862 585
R1633 B.n864 B.n19 585
R1634 B.n866 B.n865 585
R1635 B.n867 B.n18 585
R1636 B.n869 B.n868 585
R1637 B.n870 B.n17 585
R1638 B.n872 B.n871 585
R1639 B.n873 B.n16 585
R1640 B.n875 B.n874 585
R1641 B.n876 B.n15 585
R1642 B.n878 B.n877 585
R1643 B.n879 B.n14 585
R1644 B.n881 B.n880 585
R1645 B.n882 B.n13 585
R1646 B.n884 B.n883 585
R1647 B.n885 B.n12 585
R1648 B.n887 B.n886 585
R1649 B.n888 B.n11 585
R1650 B.n890 B.n889 585
R1651 B.n891 B.n10 585
R1652 B.n893 B.n892 585
R1653 B.n894 B.n9 585
R1654 B.n896 B.n895 585
R1655 B.n897 B.n8 585
R1656 B.n899 B.n898 585
R1657 B.n900 B.n7 585
R1658 B.n902 B.n901 585
R1659 B.n903 B.n6 585
R1660 B.n905 B.n904 585
R1661 B.n906 B.n5 585
R1662 B.n908 B.n907 585
R1663 B.n909 B.n4 585
R1664 B.n911 B.n910 585
R1665 B.n912 B.n3 585
R1666 B.n914 B.n913 585
R1667 B.n915 B.n0 585
R1668 B.n2 B.n1 585
R1669 B.n237 B.n236 585
R1670 B.n239 B.n238 585
R1671 B.n240 B.n235 585
R1672 B.n242 B.n241 585
R1673 B.n243 B.n234 585
R1674 B.n245 B.n244 585
R1675 B.n246 B.n233 585
R1676 B.n248 B.n247 585
R1677 B.n249 B.n232 585
R1678 B.n251 B.n250 585
R1679 B.n252 B.n231 585
R1680 B.n254 B.n253 585
R1681 B.n255 B.n230 585
R1682 B.n257 B.n256 585
R1683 B.n258 B.n229 585
R1684 B.n260 B.n259 585
R1685 B.n261 B.n228 585
R1686 B.n263 B.n262 585
R1687 B.n264 B.n227 585
R1688 B.n266 B.n265 585
R1689 B.n267 B.n226 585
R1690 B.n269 B.n268 585
R1691 B.n270 B.n225 585
R1692 B.n272 B.n271 585
R1693 B.n273 B.n224 585
R1694 B.n275 B.n274 585
R1695 B.n276 B.n223 585
R1696 B.n278 B.n277 585
R1697 B.n279 B.n222 585
R1698 B.n281 B.n280 585
R1699 B.n282 B.n221 585
R1700 B.n284 B.n283 585
R1701 B.n285 B.n220 585
R1702 B.n287 B.n286 585
R1703 B.n288 B.n219 585
R1704 B.n290 B.n289 585
R1705 B.n291 B.n218 585
R1706 B.n293 B.n292 585
R1707 B.n294 B.n217 585
R1708 B.n296 B.n295 585
R1709 B.n297 B.n216 585
R1710 B.n299 B.n298 585
R1711 B.n300 B.n215 585
R1712 B.n302 B.n301 585
R1713 B.n303 B.n214 585
R1714 B.n305 B.n304 585
R1715 B.n306 B.n213 585
R1716 B.n308 B.n307 585
R1717 B.n309 B.n212 585
R1718 B.n311 B.n310 585
R1719 B.n312 B.n211 585
R1720 B.n314 B.n313 585
R1721 B.n315 B.n210 585
R1722 B.n174 B.t10 527.369
R1723 B.n64 B.t2 527.369
R1724 B.n182 B.t4 527.369
R1725 B.n56 B.t8 527.369
R1726 B.n316 B.n315 526.135
R1727 B.n494 B.n147 526.135
R1728 B.n658 B.n657 526.135
R1729 B.n836 B.n29 526.135
R1730 B.n175 B.t11 450.957
R1731 B.n65 B.t1 450.957
R1732 B.n183 B.t5 450.955
R1733 B.n57 B.t7 450.955
R1734 B.n182 B.t3 317.207
R1735 B.n174 B.t9 317.207
R1736 B.n64 B.t0 317.207
R1737 B.n56 B.t6 317.207
R1738 B.n917 B.n916 256.663
R1739 B.n916 B.n915 235.042
R1740 B.n916 B.n2 235.042
R1741 B.n316 B.n209 163.367
R1742 B.n320 B.n209 163.367
R1743 B.n321 B.n320 163.367
R1744 B.n322 B.n321 163.367
R1745 B.n322 B.n207 163.367
R1746 B.n326 B.n207 163.367
R1747 B.n327 B.n326 163.367
R1748 B.n328 B.n327 163.367
R1749 B.n328 B.n205 163.367
R1750 B.n332 B.n205 163.367
R1751 B.n333 B.n332 163.367
R1752 B.n334 B.n333 163.367
R1753 B.n334 B.n203 163.367
R1754 B.n338 B.n203 163.367
R1755 B.n339 B.n338 163.367
R1756 B.n340 B.n339 163.367
R1757 B.n340 B.n201 163.367
R1758 B.n344 B.n201 163.367
R1759 B.n345 B.n344 163.367
R1760 B.n346 B.n345 163.367
R1761 B.n346 B.n199 163.367
R1762 B.n350 B.n199 163.367
R1763 B.n351 B.n350 163.367
R1764 B.n352 B.n351 163.367
R1765 B.n352 B.n197 163.367
R1766 B.n356 B.n197 163.367
R1767 B.n357 B.n356 163.367
R1768 B.n358 B.n357 163.367
R1769 B.n358 B.n195 163.367
R1770 B.n362 B.n195 163.367
R1771 B.n363 B.n362 163.367
R1772 B.n364 B.n363 163.367
R1773 B.n364 B.n193 163.367
R1774 B.n368 B.n193 163.367
R1775 B.n369 B.n368 163.367
R1776 B.n370 B.n369 163.367
R1777 B.n370 B.n191 163.367
R1778 B.n374 B.n191 163.367
R1779 B.n375 B.n374 163.367
R1780 B.n376 B.n375 163.367
R1781 B.n376 B.n189 163.367
R1782 B.n380 B.n189 163.367
R1783 B.n381 B.n380 163.367
R1784 B.n382 B.n381 163.367
R1785 B.n382 B.n187 163.367
R1786 B.n386 B.n187 163.367
R1787 B.n387 B.n386 163.367
R1788 B.n388 B.n387 163.367
R1789 B.n388 B.n185 163.367
R1790 B.n392 B.n185 163.367
R1791 B.n393 B.n392 163.367
R1792 B.n394 B.n393 163.367
R1793 B.n394 B.n181 163.367
R1794 B.n399 B.n181 163.367
R1795 B.n400 B.n399 163.367
R1796 B.n401 B.n400 163.367
R1797 B.n401 B.n179 163.367
R1798 B.n405 B.n179 163.367
R1799 B.n406 B.n405 163.367
R1800 B.n407 B.n406 163.367
R1801 B.n407 B.n177 163.367
R1802 B.n411 B.n177 163.367
R1803 B.n412 B.n411 163.367
R1804 B.n412 B.n173 163.367
R1805 B.n416 B.n173 163.367
R1806 B.n417 B.n416 163.367
R1807 B.n418 B.n417 163.367
R1808 B.n418 B.n171 163.367
R1809 B.n422 B.n171 163.367
R1810 B.n423 B.n422 163.367
R1811 B.n424 B.n423 163.367
R1812 B.n424 B.n169 163.367
R1813 B.n428 B.n169 163.367
R1814 B.n429 B.n428 163.367
R1815 B.n430 B.n429 163.367
R1816 B.n430 B.n167 163.367
R1817 B.n434 B.n167 163.367
R1818 B.n435 B.n434 163.367
R1819 B.n436 B.n435 163.367
R1820 B.n436 B.n165 163.367
R1821 B.n440 B.n165 163.367
R1822 B.n441 B.n440 163.367
R1823 B.n442 B.n441 163.367
R1824 B.n442 B.n163 163.367
R1825 B.n446 B.n163 163.367
R1826 B.n447 B.n446 163.367
R1827 B.n448 B.n447 163.367
R1828 B.n448 B.n161 163.367
R1829 B.n452 B.n161 163.367
R1830 B.n453 B.n452 163.367
R1831 B.n454 B.n453 163.367
R1832 B.n454 B.n159 163.367
R1833 B.n458 B.n159 163.367
R1834 B.n459 B.n458 163.367
R1835 B.n460 B.n459 163.367
R1836 B.n460 B.n157 163.367
R1837 B.n464 B.n157 163.367
R1838 B.n465 B.n464 163.367
R1839 B.n466 B.n465 163.367
R1840 B.n466 B.n155 163.367
R1841 B.n470 B.n155 163.367
R1842 B.n471 B.n470 163.367
R1843 B.n472 B.n471 163.367
R1844 B.n472 B.n153 163.367
R1845 B.n476 B.n153 163.367
R1846 B.n477 B.n476 163.367
R1847 B.n478 B.n477 163.367
R1848 B.n478 B.n151 163.367
R1849 B.n482 B.n151 163.367
R1850 B.n483 B.n482 163.367
R1851 B.n484 B.n483 163.367
R1852 B.n484 B.n149 163.367
R1853 B.n488 B.n149 163.367
R1854 B.n489 B.n488 163.367
R1855 B.n490 B.n489 163.367
R1856 B.n490 B.n147 163.367
R1857 B.n657 B.n656 163.367
R1858 B.n656 B.n93 163.367
R1859 B.n652 B.n93 163.367
R1860 B.n652 B.n651 163.367
R1861 B.n651 B.n650 163.367
R1862 B.n650 B.n95 163.367
R1863 B.n646 B.n95 163.367
R1864 B.n646 B.n645 163.367
R1865 B.n645 B.n644 163.367
R1866 B.n644 B.n97 163.367
R1867 B.n640 B.n97 163.367
R1868 B.n640 B.n639 163.367
R1869 B.n639 B.n638 163.367
R1870 B.n638 B.n99 163.367
R1871 B.n634 B.n99 163.367
R1872 B.n634 B.n633 163.367
R1873 B.n633 B.n632 163.367
R1874 B.n632 B.n101 163.367
R1875 B.n628 B.n101 163.367
R1876 B.n628 B.n627 163.367
R1877 B.n627 B.n626 163.367
R1878 B.n626 B.n103 163.367
R1879 B.n622 B.n103 163.367
R1880 B.n622 B.n621 163.367
R1881 B.n621 B.n620 163.367
R1882 B.n620 B.n105 163.367
R1883 B.n616 B.n105 163.367
R1884 B.n616 B.n615 163.367
R1885 B.n615 B.n614 163.367
R1886 B.n614 B.n107 163.367
R1887 B.n610 B.n107 163.367
R1888 B.n610 B.n609 163.367
R1889 B.n609 B.n608 163.367
R1890 B.n608 B.n109 163.367
R1891 B.n604 B.n109 163.367
R1892 B.n604 B.n603 163.367
R1893 B.n603 B.n602 163.367
R1894 B.n602 B.n111 163.367
R1895 B.n598 B.n111 163.367
R1896 B.n598 B.n597 163.367
R1897 B.n597 B.n596 163.367
R1898 B.n596 B.n113 163.367
R1899 B.n592 B.n113 163.367
R1900 B.n592 B.n591 163.367
R1901 B.n591 B.n590 163.367
R1902 B.n590 B.n115 163.367
R1903 B.n586 B.n115 163.367
R1904 B.n586 B.n585 163.367
R1905 B.n585 B.n584 163.367
R1906 B.n584 B.n117 163.367
R1907 B.n580 B.n117 163.367
R1908 B.n580 B.n579 163.367
R1909 B.n579 B.n578 163.367
R1910 B.n578 B.n119 163.367
R1911 B.n574 B.n119 163.367
R1912 B.n574 B.n573 163.367
R1913 B.n573 B.n572 163.367
R1914 B.n572 B.n121 163.367
R1915 B.n568 B.n121 163.367
R1916 B.n568 B.n567 163.367
R1917 B.n567 B.n566 163.367
R1918 B.n566 B.n123 163.367
R1919 B.n562 B.n123 163.367
R1920 B.n562 B.n561 163.367
R1921 B.n561 B.n560 163.367
R1922 B.n560 B.n125 163.367
R1923 B.n556 B.n125 163.367
R1924 B.n556 B.n555 163.367
R1925 B.n555 B.n554 163.367
R1926 B.n554 B.n127 163.367
R1927 B.n550 B.n127 163.367
R1928 B.n550 B.n549 163.367
R1929 B.n549 B.n548 163.367
R1930 B.n548 B.n129 163.367
R1931 B.n544 B.n129 163.367
R1932 B.n544 B.n543 163.367
R1933 B.n543 B.n542 163.367
R1934 B.n542 B.n131 163.367
R1935 B.n538 B.n131 163.367
R1936 B.n538 B.n537 163.367
R1937 B.n537 B.n536 163.367
R1938 B.n536 B.n133 163.367
R1939 B.n532 B.n133 163.367
R1940 B.n532 B.n531 163.367
R1941 B.n531 B.n530 163.367
R1942 B.n530 B.n135 163.367
R1943 B.n526 B.n135 163.367
R1944 B.n526 B.n525 163.367
R1945 B.n525 B.n524 163.367
R1946 B.n524 B.n137 163.367
R1947 B.n520 B.n137 163.367
R1948 B.n520 B.n519 163.367
R1949 B.n519 B.n518 163.367
R1950 B.n518 B.n139 163.367
R1951 B.n514 B.n139 163.367
R1952 B.n514 B.n513 163.367
R1953 B.n513 B.n512 163.367
R1954 B.n512 B.n141 163.367
R1955 B.n508 B.n141 163.367
R1956 B.n508 B.n507 163.367
R1957 B.n507 B.n506 163.367
R1958 B.n506 B.n143 163.367
R1959 B.n502 B.n143 163.367
R1960 B.n502 B.n501 163.367
R1961 B.n501 B.n500 163.367
R1962 B.n500 B.n145 163.367
R1963 B.n496 B.n145 163.367
R1964 B.n496 B.n495 163.367
R1965 B.n495 B.n494 163.367
R1966 B.n832 B.n29 163.367
R1967 B.n832 B.n831 163.367
R1968 B.n831 B.n830 163.367
R1969 B.n830 B.n31 163.367
R1970 B.n826 B.n31 163.367
R1971 B.n826 B.n825 163.367
R1972 B.n825 B.n824 163.367
R1973 B.n824 B.n33 163.367
R1974 B.n820 B.n33 163.367
R1975 B.n820 B.n819 163.367
R1976 B.n819 B.n818 163.367
R1977 B.n818 B.n35 163.367
R1978 B.n814 B.n35 163.367
R1979 B.n814 B.n813 163.367
R1980 B.n813 B.n812 163.367
R1981 B.n812 B.n37 163.367
R1982 B.n808 B.n37 163.367
R1983 B.n808 B.n807 163.367
R1984 B.n807 B.n806 163.367
R1985 B.n806 B.n39 163.367
R1986 B.n802 B.n39 163.367
R1987 B.n802 B.n801 163.367
R1988 B.n801 B.n800 163.367
R1989 B.n800 B.n41 163.367
R1990 B.n796 B.n41 163.367
R1991 B.n796 B.n795 163.367
R1992 B.n795 B.n794 163.367
R1993 B.n794 B.n43 163.367
R1994 B.n790 B.n43 163.367
R1995 B.n790 B.n789 163.367
R1996 B.n789 B.n788 163.367
R1997 B.n788 B.n45 163.367
R1998 B.n784 B.n45 163.367
R1999 B.n784 B.n783 163.367
R2000 B.n783 B.n782 163.367
R2001 B.n782 B.n47 163.367
R2002 B.n778 B.n47 163.367
R2003 B.n778 B.n777 163.367
R2004 B.n777 B.n776 163.367
R2005 B.n776 B.n49 163.367
R2006 B.n772 B.n49 163.367
R2007 B.n772 B.n771 163.367
R2008 B.n771 B.n770 163.367
R2009 B.n770 B.n51 163.367
R2010 B.n766 B.n51 163.367
R2011 B.n766 B.n765 163.367
R2012 B.n765 B.n764 163.367
R2013 B.n764 B.n53 163.367
R2014 B.n760 B.n53 163.367
R2015 B.n760 B.n759 163.367
R2016 B.n759 B.n758 163.367
R2017 B.n758 B.n55 163.367
R2018 B.n754 B.n55 163.367
R2019 B.n754 B.n753 163.367
R2020 B.n753 B.n59 163.367
R2021 B.n749 B.n59 163.367
R2022 B.n749 B.n748 163.367
R2023 B.n748 B.n747 163.367
R2024 B.n747 B.n61 163.367
R2025 B.n743 B.n61 163.367
R2026 B.n743 B.n742 163.367
R2027 B.n742 B.n741 163.367
R2028 B.n741 B.n63 163.367
R2029 B.n736 B.n63 163.367
R2030 B.n736 B.n735 163.367
R2031 B.n735 B.n734 163.367
R2032 B.n734 B.n67 163.367
R2033 B.n730 B.n67 163.367
R2034 B.n730 B.n729 163.367
R2035 B.n729 B.n728 163.367
R2036 B.n728 B.n69 163.367
R2037 B.n724 B.n69 163.367
R2038 B.n724 B.n723 163.367
R2039 B.n723 B.n722 163.367
R2040 B.n722 B.n71 163.367
R2041 B.n718 B.n71 163.367
R2042 B.n718 B.n717 163.367
R2043 B.n717 B.n716 163.367
R2044 B.n716 B.n73 163.367
R2045 B.n712 B.n73 163.367
R2046 B.n712 B.n711 163.367
R2047 B.n711 B.n710 163.367
R2048 B.n710 B.n75 163.367
R2049 B.n706 B.n75 163.367
R2050 B.n706 B.n705 163.367
R2051 B.n705 B.n704 163.367
R2052 B.n704 B.n77 163.367
R2053 B.n700 B.n77 163.367
R2054 B.n700 B.n699 163.367
R2055 B.n699 B.n698 163.367
R2056 B.n698 B.n79 163.367
R2057 B.n694 B.n79 163.367
R2058 B.n694 B.n693 163.367
R2059 B.n693 B.n692 163.367
R2060 B.n692 B.n81 163.367
R2061 B.n688 B.n81 163.367
R2062 B.n688 B.n687 163.367
R2063 B.n687 B.n686 163.367
R2064 B.n686 B.n83 163.367
R2065 B.n682 B.n83 163.367
R2066 B.n682 B.n681 163.367
R2067 B.n681 B.n680 163.367
R2068 B.n680 B.n85 163.367
R2069 B.n676 B.n85 163.367
R2070 B.n676 B.n675 163.367
R2071 B.n675 B.n674 163.367
R2072 B.n674 B.n87 163.367
R2073 B.n670 B.n87 163.367
R2074 B.n670 B.n669 163.367
R2075 B.n669 B.n668 163.367
R2076 B.n668 B.n89 163.367
R2077 B.n664 B.n89 163.367
R2078 B.n664 B.n663 163.367
R2079 B.n663 B.n662 163.367
R2080 B.n662 B.n91 163.367
R2081 B.n658 B.n91 163.367
R2082 B.n837 B.n836 163.367
R2083 B.n838 B.n837 163.367
R2084 B.n838 B.n27 163.367
R2085 B.n842 B.n27 163.367
R2086 B.n843 B.n842 163.367
R2087 B.n844 B.n843 163.367
R2088 B.n844 B.n25 163.367
R2089 B.n848 B.n25 163.367
R2090 B.n849 B.n848 163.367
R2091 B.n850 B.n849 163.367
R2092 B.n850 B.n23 163.367
R2093 B.n854 B.n23 163.367
R2094 B.n855 B.n854 163.367
R2095 B.n856 B.n855 163.367
R2096 B.n856 B.n21 163.367
R2097 B.n860 B.n21 163.367
R2098 B.n861 B.n860 163.367
R2099 B.n862 B.n861 163.367
R2100 B.n862 B.n19 163.367
R2101 B.n866 B.n19 163.367
R2102 B.n867 B.n866 163.367
R2103 B.n868 B.n867 163.367
R2104 B.n868 B.n17 163.367
R2105 B.n872 B.n17 163.367
R2106 B.n873 B.n872 163.367
R2107 B.n874 B.n873 163.367
R2108 B.n874 B.n15 163.367
R2109 B.n878 B.n15 163.367
R2110 B.n879 B.n878 163.367
R2111 B.n880 B.n879 163.367
R2112 B.n880 B.n13 163.367
R2113 B.n884 B.n13 163.367
R2114 B.n885 B.n884 163.367
R2115 B.n886 B.n885 163.367
R2116 B.n886 B.n11 163.367
R2117 B.n890 B.n11 163.367
R2118 B.n891 B.n890 163.367
R2119 B.n892 B.n891 163.367
R2120 B.n892 B.n9 163.367
R2121 B.n896 B.n9 163.367
R2122 B.n897 B.n896 163.367
R2123 B.n898 B.n897 163.367
R2124 B.n898 B.n7 163.367
R2125 B.n902 B.n7 163.367
R2126 B.n903 B.n902 163.367
R2127 B.n904 B.n903 163.367
R2128 B.n904 B.n5 163.367
R2129 B.n908 B.n5 163.367
R2130 B.n909 B.n908 163.367
R2131 B.n910 B.n909 163.367
R2132 B.n910 B.n3 163.367
R2133 B.n914 B.n3 163.367
R2134 B.n915 B.n914 163.367
R2135 B.n237 B.n2 163.367
R2136 B.n238 B.n237 163.367
R2137 B.n238 B.n235 163.367
R2138 B.n242 B.n235 163.367
R2139 B.n243 B.n242 163.367
R2140 B.n244 B.n243 163.367
R2141 B.n244 B.n233 163.367
R2142 B.n248 B.n233 163.367
R2143 B.n249 B.n248 163.367
R2144 B.n250 B.n249 163.367
R2145 B.n250 B.n231 163.367
R2146 B.n254 B.n231 163.367
R2147 B.n255 B.n254 163.367
R2148 B.n256 B.n255 163.367
R2149 B.n256 B.n229 163.367
R2150 B.n260 B.n229 163.367
R2151 B.n261 B.n260 163.367
R2152 B.n262 B.n261 163.367
R2153 B.n262 B.n227 163.367
R2154 B.n266 B.n227 163.367
R2155 B.n267 B.n266 163.367
R2156 B.n268 B.n267 163.367
R2157 B.n268 B.n225 163.367
R2158 B.n272 B.n225 163.367
R2159 B.n273 B.n272 163.367
R2160 B.n274 B.n273 163.367
R2161 B.n274 B.n223 163.367
R2162 B.n278 B.n223 163.367
R2163 B.n279 B.n278 163.367
R2164 B.n280 B.n279 163.367
R2165 B.n280 B.n221 163.367
R2166 B.n284 B.n221 163.367
R2167 B.n285 B.n284 163.367
R2168 B.n286 B.n285 163.367
R2169 B.n286 B.n219 163.367
R2170 B.n290 B.n219 163.367
R2171 B.n291 B.n290 163.367
R2172 B.n292 B.n291 163.367
R2173 B.n292 B.n217 163.367
R2174 B.n296 B.n217 163.367
R2175 B.n297 B.n296 163.367
R2176 B.n298 B.n297 163.367
R2177 B.n298 B.n215 163.367
R2178 B.n302 B.n215 163.367
R2179 B.n303 B.n302 163.367
R2180 B.n304 B.n303 163.367
R2181 B.n304 B.n213 163.367
R2182 B.n308 B.n213 163.367
R2183 B.n309 B.n308 163.367
R2184 B.n310 B.n309 163.367
R2185 B.n310 B.n211 163.367
R2186 B.n314 B.n211 163.367
R2187 B.n315 B.n314 163.367
R2188 B.n183 B.n182 76.4126
R2189 B.n175 B.n174 76.4126
R2190 B.n65 B.n64 76.4126
R2191 B.n57 B.n56 76.4126
R2192 B.n397 B.n183 59.5399
R2193 B.n176 B.n175 59.5399
R2194 B.n739 B.n65 59.5399
R2195 B.n58 B.n57 59.5399
R2196 B.n835 B.n834 34.1859
R2197 B.n659 B.n92 34.1859
R2198 B.n493 B.n492 34.1859
R2199 B.n317 B.n210 34.1859
R2200 B B.n917 18.0485
R2201 B.n835 B.n28 10.6151
R2202 B.n839 B.n28 10.6151
R2203 B.n840 B.n839 10.6151
R2204 B.n841 B.n840 10.6151
R2205 B.n841 B.n26 10.6151
R2206 B.n845 B.n26 10.6151
R2207 B.n846 B.n845 10.6151
R2208 B.n847 B.n846 10.6151
R2209 B.n847 B.n24 10.6151
R2210 B.n851 B.n24 10.6151
R2211 B.n852 B.n851 10.6151
R2212 B.n853 B.n852 10.6151
R2213 B.n853 B.n22 10.6151
R2214 B.n857 B.n22 10.6151
R2215 B.n858 B.n857 10.6151
R2216 B.n859 B.n858 10.6151
R2217 B.n859 B.n20 10.6151
R2218 B.n863 B.n20 10.6151
R2219 B.n864 B.n863 10.6151
R2220 B.n865 B.n864 10.6151
R2221 B.n865 B.n18 10.6151
R2222 B.n869 B.n18 10.6151
R2223 B.n870 B.n869 10.6151
R2224 B.n871 B.n870 10.6151
R2225 B.n871 B.n16 10.6151
R2226 B.n875 B.n16 10.6151
R2227 B.n876 B.n875 10.6151
R2228 B.n877 B.n876 10.6151
R2229 B.n877 B.n14 10.6151
R2230 B.n881 B.n14 10.6151
R2231 B.n882 B.n881 10.6151
R2232 B.n883 B.n882 10.6151
R2233 B.n883 B.n12 10.6151
R2234 B.n887 B.n12 10.6151
R2235 B.n888 B.n887 10.6151
R2236 B.n889 B.n888 10.6151
R2237 B.n889 B.n10 10.6151
R2238 B.n893 B.n10 10.6151
R2239 B.n894 B.n893 10.6151
R2240 B.n895 B.n894 10.6151
R2241 B.n895 B.n8 10.6151
R2242 B.n899 B.n8 10.6151
R2243 B.n900 B.n899 10.6151
R2244 B.n901 B.n900 10.6151
R2245 B.n901 B.n6 10.6151
R2246 B.n905 B.n6 10.6151
R2247 B.n906 B.n905 10.6151
R2248 B.n907 B.n906 10.6151
R2249 B.n907 B.n4 10.6151
R2250 B.n911 B.n4 10.6151
R2251 B.n912 B.n911 10.6151
R2252 B.n913 B.n912 10.6151
R2253 B.n913 B.n0 10.6151
R2254 B.n834 B.n833 10.6151
R2255 B.n833 B.n30 10.6151
R2256 B.n829 B.n30 10.6151
R2257 B.n829 B.n828 10.6151
R2258 B.n828 B.n827 10.6151
R2259 B.n827 B.n32 10.6151
R2260 B.n823 B.n32 10.6151
R2261 B.n823 B.n822 10.6151
R2262 B.n822 B.n821 10.6151
R2263 B.n821 B.n34 10.6151
R2264 B.n817 B.n34 10.6151
R2265 B.n817 B.n816 10.6151
R2266 B.n816 B.n815 10.6151
R2267 B.n815 B.n36 10.6151
R2268 B.n811 B.n36 10.6151
R2269 B.n811 B.n810 10.6151
R2270 B.n810 B.n809 10.6151
R2271 B.n809 B.n38 10.6151
R2272 B.n805 B.n38 10.6151
R2273 B.n805 B.n804 10.6151
R2274 B.n804 B.n803 10.6151
R2275 B.n803 B.n40 10.6151
R2276 B.n799 B.n40 10.6151
R2277 B.n799 B.n798 10.6151
R2278 B.n798 B.n797 10.6151
R2279 B.n797 B.n42 10.6151
R2280 B.n793 B.n42 10.6151
R2281 B.n793 B.n792 10.6151
R2282 B.n792 B.n791 10.6151
R2283 B.n791 B.n44 10.6151
R2284 B.n787 B.n44 10.6151
R2285 B.n787 B.n786 10.6151
R2286 B.n786 B.n785 10.6151
R2287 B.n785 B.n46 10.6151
R2288 B.n781 B.n46 10.6151
R2289 B.n781 B.n780 10.6151
R2290 B.n780 B.n779 10.6151
R2291 B.n779 B.n48 10.6151
R2292 B.n775 B.n48 10.6151
R2293 B.n775 B.n774 10.6151
R2294 B.n774 B.n773 10.6151
R2295 B.n773 B.n50 10.6151
R2296 B.n769 B.n50 10.6151
R2297 B.n769 B.n768 10.6151
R2298 B.n768 B.n767 10.6151
R2299 B.n767 B.n52 10.6151
R2300 B.n763 B.n52 10.6151
R2301 B.n763 B.n762 10.6151
R2302 B.n762 B.n761 10.6151
R2303 B.n761 B.n54 10.6151
R2304 B.n757 B.n54 10.6151
R2305 B.n757 B.n756 10.6151
R2306 B.n756 B.n755 10.6151
R2307 B.n752 B.n751 10.6151
R2308 B.n751 B.n750 10.6151
R2309 B.n750 B.n60 10.6151
R2310 B.n746 B.n60 10.6151
R2311 B.n746 B.n745 10.6151
R2312 B.n745 B.n744 10.6151
R2313 B.n744 B.n62 10.6151
R2314 B.n740 B.n62 10.6151
R2315 B.n738 B.n737 10.6151
R2316 B.n737 B.n66 10.6151
R2317 B.n733 B.n66 10.6151
R2318 B.n733 B.n732 10.6151
R2319 B.n732 B.n731 10.6151
R2320 B.n731 B.n68 10.6151
R2321 B.n727 B.n68 10.6151
R2322 B.n727 B.n726 10.6151
R2323 B.n726 B.n725 10.6151
R2324 B.n725 B.n70 10.6151
R2325 B.n721 B.n70 10.6151
R2326 B.n721 B.n720 10.6151
R2327 B.n720 B.n719 10.6151
R2328 B.n719 B.n72 10.6151
R2329 B.n715 B.n72 10.6151
R2330 B.n715 B.n714 10.6151
R2331 B.n714 B.n713 10.6151
R2332 B.n713 B.n74 10.6151
R2333 B.n709 B.n74 10.6151
R2334 B.n709 B.n708 10.6151
R2335 B.n708 B.n707 10.6151
R2336 B.n707 B.n76 10.6151
R2337 B.n703 B.n76 10.6151
R2338 B.n703 B.n702 10.6151
R2339 B.n702 B.n701 10.6151
R2340 B.n701 B.n78 10.6151
R2341 B.n697 B.n78 10.6151
R2342 B.n697 B.n696 10.6151
R2343 B.n696 B.n695 10.6151
R2344 B.n695 B.n80 10.6151
R2345 B.n691 B.n80 10.6151
R2346 B.n691 B.n690 10.6151
R2347 B.n690 B.n689 10.6151
R2348 B.n689 B.n82 10.6151
R2349 B.n685 B.n82 10.6151
R2350 B.n685 B.n684 10.6151
R2351 B.n684 B.n683 10.6151
R2352 B.n683 B.n84 10.6151
R2353 B.n679 B.n84 10.6151
R2354 B.n679 B.n678 10.6151
R2355 B.n678 B.n677 10.6151
R2356 B.n677 B.n86 10.6151
R2357 B.n673 B.n86 10.6151
R2358 B.n673 B.n672 10.6151
R2359 B.n672 B.n671 10.6151
R2360 B.n671 B.n88 10.6151
R2361 B.n667 B.n88 10.6151
R2362 B.n667 B.n666 10.6151
R2363 B.n666 B.n665 10.6151
R2364 B.n665 B.n90 10.6151
R2365 B.n661 B.n90 10.6151
R2366 B.n661 B.n660 10.6151
R2367 B.n660 B.n659 10.6151
R2368 B.n655 B.n92 10.6151
R2369 B.n655 B.n654 10.6151
R2370 B.n654 B.n653 10.6151
R2371 B.n653 B.n94 10.6151
R2372 B.n649 B.n94 10.6151
R2373 B.n649 B.n648 10.6151
R2374 B.n648 B.n647 10.6151
R2375 B.n647 B.n96 10.6151
R2376 B.n643 B.n96 10.6151
R2377 B.n643 B.n642 10.6151
R2378 B.n642 B.n641 10.6151
R2379 B.n641 B.n98 10.6151
R2380 B.n637 B.n98 10.6151
R2381 B.n637 B.n636 10.6151
R2382 B.n636 B.n635 10.6151
R2383 B.n635 B.n100 10.6151
R2384 B.n631 B.n100 10.6151
R2385 B.n631 B.n630 10.6151
R2386 B.n630 B.n629 10.6151
R2387 B.n629 B.n102 10.6151
R2388 B.n625 B.n102 10.6151
R2389 B.n625 B.n624 10.6151
R2390 B.n624 B.n623 10.6151
R2391 B.n623 B.n104 10.6151
R2392 B.n619 B.n104 10.6151
R2393 B.n619 B.n618 10.6151
R2394 B.n618 B.n617 10.6151
R2395 B.n617 B.n106 10.6151
R2396 B.n613 B.n106 10.6151
R2397 B.n613 B.n612 10.6151
R2398 B.n612 B.n611 10.6151
R2399 B.n611 B.n108 10.6151
R2400 B.n607 B.n108 10.6151
R2401 B.n607 B.n606 10.6151
R2402 B.n606 B.n605 10.6151
R2403 B.n605 B.n110 10.6151
R2404 B.n601 B.n110 10.6151
R2405 B.n601 B.n600 10.6151
R2406 B.n600 B.n599 10.6151
R2407 B.n599 B.n112 10.6151
R2408 B.n595 B.n112 10.6151
R2409 B.n595 B.n594 10.6151
R2410 B.n594 B.n593 10.6151
R2411 B.n593 B.n114 10.6151
R2412 B.n589 B.n114 10.6151
R2413 B.n589 B.n588 10.6151
R2414 B.n588 B.n587 10.6151
R2415 B.n587 B.n116 10.6151
R2416 B.n583 B.n116 10.6151
R2417 B.n583 B.n582 10.6151
R2418 B.n582 B.n581 10.6151
R2419 B.n581 B.n118 10.6151
R2420 B.n577 B.n118 10.6151
R2421 B.n577 B.n576 10.6151
R2422 B.n576 B.n575 10.6151
R2423 B.n575 B.n120 10.6151
R2424 B.n571 B.n120 10.6151
R2425 B.n571 B.n570 10.6151
R2426 B.n570 B.n569 10.6151
R2427 B.n569 B.n122 10.6151
R2428 B.n565 B.n122 10.6151
R2429 B.n565 B.n564 10.6151
R2430 B.n564 B.n563 10.6151
R2431 B.n563 B.n124 10.6151
R2432 B.n559 B.n124 10.6151
R2433 B.n559 B.n558 10.6151
R2434 B.n558 B.n557 10.6151
R2435 B.n557 B.n126 10.6151
R2436 B.n553 B.n126 10.6151
R2437 B.n553 B.n552 10.6151
R2438 B.n552 B.n551 10.6151
R2439 B.n551 B.n128 10.6151
R2440 B.n547 B.n128 10.6151
R2441 B.n547 B.n546 10.6151
R2442 B.n546 B.n545 10.6151
R2443 B.n545 B.n130 10.6151
R2444 B.n541 B.n130 10.6151
R2445 B.n541 B.n540 10.6151
R2446 B.n540 B.n539 10.6151
R2447 B.n539 B.n132 10.6151
R2448 B.n535 B.n132 10.6151
R2449 B.n535 B.n534 10.6151
R2450 B.n534 B.n533 10.6151
R2451 B.n533 B.n134 10.6151
R2452 B.n529 B.n134 10.6151
R2453 B.n529 B.n528 10.6151
R2454 B.n528 B.n527 10.6151
R2455 B.n527 B.n136 10.6151
R2456 B.n523 B.n136 10.6151
R2457 B.n523 B.n522 10.6151
R2458 B.n522 B.n521 10.6151
R2459 B.n521 B.n138 10.6151
R2460 B.n517 B.n138 10.6151
R2461 B.n517 B.n516 10.6151
R2462 B.n516 B.n515 10.6151
R2463 B.n515 B.n140 10.6151
R2464 B.n511 B.n140 10.6151
R2465 B.n511 B.n510 10.6151
R2466 B.n510 B.n509 10.6151
R2467 B.n509 B.n142 10.6151
R2468 B.n505 B.n142 10.6151
R2469 B.n505 B.n504 10.6151
R2470 B.n504 B.n503 10.6151
R2471 B.n503 B.n144 10.6151
R2472 B.n499 B.n144 10.6151
R2473 B.n499 B.n498 10.6151
R2474 B.n498 B.n497 10.6151
R2475 B.n497 B.n146 10.6151
R2476 B.n493 B.n146 10.6151
R2477 B.n236 B.n1 10.6151
R2478 B.n239 B.n236 10.6151
R2479 B.n240 B.n239 10.6151
R2480 B.n241 B.n240 10.6151
R2481 B.n241 B.n234 10.6151
R2482 B.n245 B.n234 10.6151
R2483 B.n246 B.n245 10.6151
R2484 B.n247 B.n246 10.6151
R2485 B.n247 B.n232 10.6151
R2486 B.n251 B.n232 10.6151
R2487 B.n252 B.n251 10.6151
R2488 B.n253 B.n252 10.6151
R2489 B.n253 B.n230 10.6151
R2490 B.n257 B.n230 10.6151
R2491 B.n258 B.n257 10.6151
R2492 B.n259 B.n258 10.6151
R2493 B.n259 B.n228 10.6151
R2494 B.n263 B.n228 10.6151
R2495 B.n264 B.n263 10.6151
R2496 B.n265 B.n264 10.6151
R2497 B.n265 B.n226 10.6151
R2498 B.n269 B.n226 10.6151
R2499 B.n270 B.n269 10.6151
R2500 B.n271 B.n270 10.6151
R2501 B.n271 B.n224 10.6151
R2502 B.n275 B.n224 10.6151
R2503 B.n276 B.n275 10.6151
R2504 B.n277 B.n276 10.6151
R2505 B.n277 B.n222 10.6151
R2506 B.n281 B.n222 10.6151
R2507 B.n282 B.n281 10.6151
R2508 B.n283 B.n282 10.6151
R2509 B.n283 B.n220 10.6151
R2510 B.n287 B.n220 10.6151
R2511 B.n288 B.n287 10.6151
R2512 B.n289 B.n288 10.6151
R2513 B.n289 B.n218 10.6151
R2514 B.n293 B.n218 10.6151
R2515 B.n294 B.n293 10.6151
R2516 B.n295 B.n294 10.6151
R2517 B.n295 B.n216 10.6151
R2518 B.n299 B.n216 10.6151
R2519 B.n300 B.n299 10.6151
R2520 B.n301 B.n300 10.6151
R2521 B.n301 B.n214 10.6151
R2522 B.n305 B.n214 10.6151
R2523 B.n306 B.n305 10.6151
R2524 B.n307 B.n306 10.6151
R2525 B.n307 B.n212 10.6151
R2526 B.n311 B.n212 10.6151
R2527 B.n312 B.n311 10.6151
R2528 B.n313 B.n312 10.6151
R2529 B.n313 B.n210 10.6151
R2530 B.n318 B.n317 10.6151
R2531 B.n319 B.n318 10.6151
R2532 B.n319 B.n208 10.6151
R2533 B.n323 B.n208 10.6151
R2534 B.n324 B.n323 10.6151
R2535 B.n325 B.n324 10.6151
R2536 B.n325 B.n206 10.6151
R2537 B.n329 B.n206 10.6151
R2538 B.n330 B.n329 10.6151
R2539 B.n331 B.n330 10.6151
R2540 B.n331 B.n204 10.6151
R2541 B.n335 B.n204 10.6151
R2542 B.n336 B.n335 10.6151
R2543 B.n337 B.n336 10.6151
R2544 B.n337 B.n202 10.6151
R2545 B.n341 B.n202 10.6151
R2546 B.n342 B.n341 10.6151
R2547 B.n343 B.n342 10.6151
R2548 B.n343 B.n200 10.6151
R2549 B.n347 B.n200 10.6151
R2550 B.n348 B.n347 10.6151
R2551 B.n349 B.n348 10.6151
R2552 B.n349 B.n198 10.6151
R2553 B.n353 B.n198 10.6151
R2554 B.n354 B.n353 10.6151
R2555 B.n355 B.n354 10.6151
R2556 B.n355 B.n196 10.6151
R2557 B.n359 B.n196 10.6151
R2558 B.n360 B.n359 10.6151
R2559 B.n361 B.n360 10.6151
R2560 B.n361 B.n194 10.6151
R2561 B.n365 B.n194 10.6151
R2562 B.n366 B.n365 10.6151
R2563 B.n367 B.n366 10.6151
R2564 B.n367 B.n192 10.6151
R2565 B.n371 B.n192 10.6151
R2566 B.n372 B.n371 10.6151
R2567 B.n373 B.n372 10.6151
R2568 B.n373 B.n190 10.6151
R2569 B.n377 B.n190 10.6151
R2570 B.n378 B.n377 10.6151
R2571 B.n379 B.n378 10.6151
R2572 B.n379 B.n188 10.6151
R2573 B.n383 B.n188 10.6151
R2574 B.n384 B.n383 10.6151
R2575 B.n385 B.n384 10.6151
R2576 B.n385 B.n186 10.6151
R2577 B.n389 B.n186 10.6151
R2578 B.n390 B.n389 10.6151
R2579 B.n391 B.n390 10.6151
R2580 B.n391 B.n184 10.6151
R2581 B.n395 B.n184 10.6151
R2582 B.n396 B.n395 10.6151
R2583 B.n398 B.n180 10.6151
R2584 B.n402 B.n180 10.6151
R2585 B.n403 B.n402 10.6151
R2586 B.n404 B.n403 10.6151
R2587 B.n404 B.n178 10.6151
R2588 B.n408 B.n178 10.6151
R2589 B.n409 B.n408 10.6151
R2590 B.n410 B.n409 10.6151
R2591 B.n414 B.n413 10.6151
R2592 B.n415 B.n414 10.6151
R2593 B.n415 B.n172 10.6151
R2594 B.n419 B.n172 10.6151
R2595 B.n420 B.n419 10.6151
R2596 B.n421 B.n420 10.6151
R2597 B.n421 B.n170 10.6151
R2598 B.n425 B.n170 10.6151
R2599 B.n426 B.n425 10.6151
R2600 B.n427 B.n426 10.6151
R2601 B.n427 B.n168 10.6151
R2602 B.n431 B.n168 10.6151
R2603 B.n432 B.n431 10.6151
R2604 B.n433 B.n432 10.6151
R2605 B.n433 B.n166 10.6151
R2606 B.n437 B.n166 10.6151
R2607 B.n438 B.n437 10.6151
R2608 B.n439 B.n438 10.6151
R2609 B.n439 B.n164 10.6151
R2610 B.n443 B.n164 10.6151
R2611 B.n444 B.n443 10.6151
R2612 B.n445 B.n444 10.6151
R2613 B.n445 B.n162 10.6151
R2614 B.n449 B.n162 10.6151
R2615 B.n450 B.n449 10.6151
R2616 B.n451 B.n450 10.6151
R2617 B.n451 B.n160 10.6151
R2618 B.n455 B.n160 10.6151
R2619 B.n456 B.n455 10.6151
R2620 B.n457 B.n456 10.6151
R2621 B.n457 B.n158 10.6151
R2622 B.n461 B.n158 10.6151
R2623 B.n462 B.n461 10.6151
R2624 B.n463 B.n462 10.6151
R2625 B.n463 B.n156 10.6151
R2626 B.n467 B.n156 10.6151
R2627 B.n468 B.n467 10.6151
R2628 B.n469 B.n468 10.6151
R2629 B.n469 B.n154 10.6151
R2630 B.n473 B.n154 10.6151
R2631 B.n474 B.n473 10.6151
R2632 B.n475 B.n474 10.6151
R2633 B.n475 B.n152 10.6151
R2634 B.n479 B.n152 10.6151
R2635 B.n480 B.n479 10.6151
R2636 B.n481 B.n480 10.6151
R2637 B.n481 B.n150 10.6151
R2638 B.n485 B.n150 10.6151
R2639 B.n486 B.n485 10.6151
R2640 B.n487 B.n486 10.6151
R2641 B.n487 B.n148 10.6151
R2642 B.n491 B.n148 10.6151
R2643 B.n492 B.n491 10.6151
R2644 B.n917 B.n0 8.11757
R2645 B.n917 B.n1 8.11757
R2646 B.n752 B.n58 6.5566
R2647 B.n740 B.n739 6.5566
R2648 B.n398 B.n397 6.5566
R2649 B.n410 B.n176 6.5566
R2650 B.n755 B.n58 4.05904
R2651 B.n739 B.n738 4.05904
R2652 B.n397 B.n396 4.05904
R2653 B.n413 B.n176 4.05904
C0 w_n4122_n4204# B 12.243f
C1 VP B 2.33359f
C2 VTAIL VDD1 9.42274f
C3 VTAIL VN 9.631861f
C4 VDD1 VDD2 1.80209f
C5 VN VDD2 9.42759f
C6 VTAIL w_n4122_n4204# 3.63162f
C7 VDD1 VN 0.152549f
C8 w_n4122_n4204# VDD2 2.94024f
C9 VTAIL VP 9.64627f
C10 VP VDD2 0.544514f
C11 VDD1 w_n4122_n4204# 2.82288f
C12 VN w_n4122_n4204# 8.11623f
C13 VDD1 VP 9.8161f
C14 VP VN 8.675871f
C15 VTAIL B 5.06251f
C16 B VDD2 2.79086f
C17 VP w_n4122_n4204# 8.651959f
C18 VDD1 B 2.69255f
C19 VN B 1.43404f
C20 VTAIL VDD2 9.48051f
C21 VDD2 VSUBS 2.26958f
C22 VDD1 VSUBS 2.285563f
C23 VTAIL VSUBS 1.530843f
C24 VN VSUBS 6.96539f
C25 VP VSUBS 3.873174f
C26 B VSUBS 5.987786f
C27 w_n4122_n4204# VSUBS 0.21225p
C28 B.n0 VSUBS 0.006634f
C29 B.n1 VSUBS 0.006634f
C30 B.n2 VSUBS 0.009812f
C31 B.n3 VSUBS 0.007519f
C32 B.n4 VSUBS 0.007519f
C33 B.n5 VSUBS 0.007519f
C34 B.n6 VSUBS 0.007519f
C35 B.n7 VSUBS 0.007519f
C36 B.n8 VSUBS 0.007519f
C37 B.n9 VSUBS 0.007519f
C38 B.n10 VSUBS 0.007519f
C39 B.n11 VSUBS 0.007519f
C40 B.n12 VSUBS 0.007519f
C41 B.n13 VSUBS 0.007519f
C42 B.n14 VSUBS 0.007519f
C43 B.n15 VSUBS 0.007519f
C44 B.n16 VSUBS 0.007519f
C45 B.n17 VSUBS 0.007519f
C46 B.n18 VSUBS 0.007519f
C47 B.n19 VSUBS 0.007519f
C48 B.n20 VSUBS 0.007519f
C49 B.n21 VSUBS 0.007519f
C50 B.n22 VSUBS 0.007519f
C51 B.n23 VSUBS 0.007519f
C52 B.n24 VSUBS 0.007519f
C53 B.n25 VSUBS 0.007519f
C54 B.n26 VSUBS 0.007519f
C55 B.n27 VSUBS 0.007519f
C56 B.n28 VSUBS 0.007519f
C57 B.n29 VSUBS 0.018372f
C58 B.n30 VSUBS 0.007519f
C59 B.n31 VSUBS 0.007519f
C60 B.n32 VSUBS 0.007519f
C61 B.n33 VSUBS 0.007519f
C62 B.n34 VSUBS 0.007519f
C63 B.n35 VSUBS 0.007519f
C64 B.n36 VSUBS 0.007519f
C65 B.n37 VSUBS 0.007519f
C66 B.n38 VSUBS 0.007519f
C67 B.n39 VSUBS 0.007519f
C68 B.n40 VSUBS 0.007519f
C69 B.n41 VSUBS 0.007519f
C70 B.n42 VSUBS 0.007519f
C71 B.n43 VSUBS 0.007519f
C72 B.n44 VSUBS 0.007519f
C73 B.n45 VSUBS 0.007519f
C74 B.n46 VSUBS 0.007519f
C75 B.n47 VSUBS 0.007519f
C76 B.n48 VSUBS 0.007519f
C77 B.n49 VSUBS 0.007519f
C78 B.n50 VSUBS 0.007519f
C79 B.n51 VSUBS 0.007519f
C80 B.n52 VSUBS 0.007519f
C81 B.n53 VSUBS 0.007519f
C82 B.n54 VSUBS 0.007519f
C83 B.n55 VSUBS 0.007519f
C84 B.t7 VSUBS 0.33028f
C85 B.t8 VSUBS 0.377079f
C86 B.t6 VSUBS 2.86791f
C87 B.n56 VSUBS 0.599725f
C88 B.n57 VSUBS 0.333718f
C89 B.n58 VSUBS 0.017421f
C90 B.n59 VSUBS 0.007519f
C91 B.n60 VSUBS 0.007519f
C92 B.n61 VSUBS 0.007519f
C93 B.n62 VSUBS 0.007519f
C94 B.n63 VSUBS 0.007519f
C95 B.t1 VSUBS 0.330283f
C96 B.t2 VSUBS 0.377083f
C97 B.t0 VSUBS 2.86791f
C98 B.n64 VSUBS 0.599722f
C99 B.n65 VSUBS 0.333714f
C100 B.n66 VSUBS 0.007519f
C101 B.n67 VSUBS 0.007519f
C102 B.n68 VSUBS 0.007519f
C103 B.n69 VSUBS 0.007519f
C104 B.n70 VSUBS 0.007519f
C105 B.n71 VSUBS 0.007519f
C106 B.n72 VSUBS 0.007519f
C107 B.n73 VSUBS 0.007519f
C108 B.n74 VSUBS 0.007519f
C109 B.n75 VSUBS 0.007519f
C110 B.n76 VSUBS 0.007519f
C111 B.n77 VSUBS 0.007519f
C112 B.n78 VSUBS 0.007519f
C113 B.n79 VSUBS 0.007519f
C114 B.n80 VSUBS 0.007519f
C115 B.n81 VSUBS 0.007519f
C116 B.n82 VSUBS 0.007519f
C117 B.n83 VSUBS 0.007519f
C118 B.n84 VSUBS 0.007519f
C119 B.n85 VSUBS 0.007519f
C120 B.n86 VSUBS 0.007519f
C121 B.n87 VSUBS 0.007519f
C122 B.n88 VSUBS 0.007519f
C123 B.n89 VSUBS 0.007519f
C124 B.n90 VSUBS 0.007519f
C125 B.n91 VSUBS 0.007519f
C126 B.n92 VSUBS 0.017896f
C127 B.n93 VSUBS 0.007519f
C128 B.n94 VSUBS 0.007519f
C129 B.n95 VSUBS 0.007519f
C130 B.n96 VSUBS 0.007519f
C131 B.n97 VSUBS 0.007519f
C132 B.n98 VSUBS 0.007519f
C133 B.n99 VSUBS 0.007519f
C134 B.n100 VSUBS 0.007519f
C135 B.n101 VSUBS 0.007519f
C136 B.n102 VSUBS 0.007519f
C137 B.n103 VSUBS 0.007519f
C138 B.n104 VSUBS 0.007519f
C139 B.n105 VSUBS 0.007519f
C140 B.n106 VSUBS 0.007519f
C141 B.n107 VSUBS 0.007519f
C142 B.n108 VSUBS 0.007519f
C143 B.n109 VSUBS 0.007519f
C144 B.n110 VSUBS 0.007519f
C145 B.n111 VSUBS 0.007519f
C146 B.n112 VSUBS 0.007519f
C147 B.n113 VSUBS 0.007519f
C148 B.n114 VSUBS 0.007519f
C149 B.n115 VSUBS 0.007519f
C150 B.n116 VSUBS 0.007519f
C151 B.n117 VSUBS 0.007519f
C152 B.n118 VSUBS 0.007519f
C153 B.n119 VSUBS 0.007519f
C154 B.n120 VSUBS 0.007519f
C155 B.n121 VSUBS 0.007519f
C156 B.n122 VSUBS 0.007519f
C157 B.n123 VSUBS 0.007519f
C158 B.n124 VSUBS 0.007519f
C159 B.n125 VSUBS 0.007519f
C160 B.n126 VSUBS 0.007519f
C161 B.n127 VSUBS 0.007519f
C162 B.n128 VSUBS 0.007519f
C163 B.n129 VSUBS 0.007519f
C164 B.n130 VSUBS 0.007519f
C165 B.n131 VSUBS 0.007519f
C166 B.n132 VSUBS 0.007519f
C167 B.n133 VSUBS 0.007519f
C168 B.n134 VSUBS 0.007519f
C169 B.n135 VSUBS 0.007519f
C170 B.n136 VSUBS 0.007519f
C171 B.n137 VSUBS 0.007519f
C172 B.n138 VSUBS 0.007519f
C173 B.n139 VSUBS 0.007519f
C174 B.n140 VSUBS 0.007519f
C175 B.n141 VSUBS 0.007519f
C176 B.n142 VSUBS 0.007519f
C177 B.n143 VSUBS 0.007519f
C178 B.n144 VSUBS 0.007519f
C179 B.n145 VSUBS 0.007519f
C180 B.n146 VSUBS 0.007519f
C181 B.n147 VSUBS 0.018372f
C182 B.n148 VSUBS 0.007519f
C183 B.n149 VSUBS 0.007519f
C184 B.n150 VSUBS 0.007519f
C185 B.n151 VSUBS 0.007519f
C186 B.n152 VSUBS 0.007519f
C187 B.n153 VSUBS 0.007519f
C188 B.n154 VSUBS 0.007519f
C189 B.n155 VSUBS 0.007519f
C190 B.n156 VSUBS 0.007519f
C191 B.n157 VSUBS 0.007519f
C192 B.n158 VSUBS 0.007519f
C193 B.n159 VSUBS 0.007519f
C194 B.n160 VSUBS 0.007519f
C195 B.n161 VSUBS 0.007519f
C196 B.n162 VSUBS 0.007519f
C197 B.n163 VSUBS 0.007519f
C198 B.n164 VSUBS 0.007519f
C199 B.n165 VSUBS 0.007519f
C200 B.n166 VSUBS 0.007519f
C201 B.n167 VSUBS 0.007519f
C202 B.n168 VSUBS 0.007519f
C203 B.n169 VSUBS 0.007519f
C204 B.n170 VSUBS 0.007519f
C205 B.n171 VSUBS 0.007519f
C206 B.n172 VSUBS 0.007519f
C207 B.n173 VSUBS 0.007519f
C208 B.t11 VSUBS 0.330283f
C209 B.t10 VSUBS 0.377083f
C210 B.t9 VSUBS 2.86791f
C211 B.n174 VSUBS 0.599722f
C212 B.n175 VSUBS 0.333714f
C213 B.n176 VSUBS 0.017421f
C214 B.n177 VSUBS 0.007519f
C215 B.n178 VSUBS 0.007519f
C216 B.n179 VSUBS 0.007519f
C217 B.n180 VSUBS 0.007519f
C218 B.n181 VSUBS 0.007519f
C219 B.t5 VSUBS 0.33028f
C220 B.t4 VSUBS 0.377079f
C221 B.t3 VSUBS 2.86791f
C222 B.n182 VSUBS 0.599725f
C223 B.n183 VSUBS 0.333718f
C224 B.n184 VSUBS 0.007519f
C225 B.n185 VSUBS 0.007519f
C226 B.n186 VSUBS 0.007519f
C227 B.n187 VSUBS 0.007519f
C228 B.n188 VSUBS 0.007519f
C229 B.n189 VSUBS 0.007519f
C230 B.n190 VSUBS 0.007519f
C231 B.n191 VSUBS 0.007519f
C232 B.n192 VSUBS 0.007519f
C233 B.n193 VSUBS 0.007519f
C234 B.n194 VSUBS 0.007519f
C235 B.n195 VSUBS 0.007519f
C236 B.n196 VSUBS 0.007519f
C237 B.n197 VSUBS 0.007519f
C238 B.n198 VSUBS 0.007519f
C239 B.n199 VSUBS 0.007519f
C240 B.n200 VSUBS 0.007519f
C241 B.n201 VSUBS 0.007519f
C242 B.n202 VSUBS 0.007519f
C243 B.n203 VSUBS 0.007519f
C244 B.n204 VSUBS 0.007519f
C245 B.n205 VSUBS 0.007519f
C246 B.n206 VSUBS 0.007519f
C247 B.n207 VSUBS 0.007519f
C248 B.n208 VSUBS 0.007519f
C249 B.n209 VSUBS 0.007519f
C250 B.n210 VSUBS 0.017896f
C251 B.n211 VSUBS 0.007519f
C252 B.n212 VSUBS 0.007519f
C253 B.n213 VSUBS 0.007519f
C254 B.n214 VSUBS 0.007519f
C255 B.n215 VSUBS 0.007519f
C256 B.n216 VSUBS 0.007519f
C257 B.n217 VSUBS 0.007519f
C258 B.n218 VSUBS 0.007519f
C259 B.n219 VSUBS 0.007519f
C260 B.n220 VSUBS 0.007519f
C261 B.n221 VSUBS 0.007519f
C262 B.n222 VSUBS 0.007519f
C263 B.n223 VSUBS 0.007519f
C264 B.n224 VSUBS 0.007519f
C265 B.n225 VSUBS 0.007519f
C266 B.n226 VSUBS 0.007519f
C267 B.n227 VSUBS 0.007519f
C268 B.n228 VSUBS 0.007519f
C269 B.n229 VSUBS 0.007519f
C270 B.n230 VSUBS 0.007519f
C271 B.n231 VSUBS 0.007519f
C272 B.n232 VSUBS 0.007519f
C273 B.n233 VSUBS 0.007519f
C274 B.n234 VSUBS 0.007519f
C275 B.n235 VSUBS 0.007519f
C276 B.n236 VSUBS 0.007519f
C277 B.n237 VSUBS 0.007519f
C278 B.n238 VSUBS 0.007519f
C279 B.n239 VSUBS 0.007519f
C280 B.n240 VSUBS 0.007519f
C281 B.n241 VSUBS 0.007519f
C282 B.n242 VSUBS 0.007519f
C283 B.n243 VSUBS 0.007519f
C284 B.n244 VSUBS 0.007519f
C285 B.n245 VSUBS 0.007519f
C286 B.n246 VSUBS 0.007519f
C287 B.n247 VSUBS 0.007519f
C288 B.n248 VSUBS 0.007519f
C289 B.n249 VSUBS 0.007519f
C290 B.n250 VSUBS 0.007519f
C291 B.n251 VSUBS 0.007519f
C292 B.n252 VSUBS 0.007519f
C293 B.n253 VSUBS 0.007519f
C294 B.n254 VSUBS 0.007519f
C295 B.n255 VSUBS 0.007519f
C296 B.n256 VSUBS 0.007519f
C297 B.n257 VSUBS 0.007519f
C298 B.n258 VSUBS 0.007519f
C299 B.n259 VSUBS 0.007519f
C300 B.n260 VSUBS 0.007519f
C301 B.n261 VSUBS 0.007519f
C302 B.n262 VSUBS 0.007519f
C303 B.n263 VSUBS 0.007519f
C304 B.n264 VSUBS 0.007519f
C305 B.n265 VSUBS 0.007519f
C306 B.n266 VSUBS 0.007519f
C307 B.n267 VSUBS 0.007519f
C308 B.n268 VSUBS 0.007519f
C309 B.n269 VSUBS 0.007519f
C310 B.n270 VSUBS 0.007519f
C311 B.n271 VSUBS 0.007519f
C312 B.n272 VSUBS 0.007519f
C313 B.n273 VSUBS 0.007519f
C314 B.n274 VSUBS 0.007519f
C315 B.n275 VSUBS 0.007519f
C316 B.n276 VSUBS 0.007519f
C317 B.n277 VSUBS 0.007519f
C318 B.n278 VSUBS 0.007519f
C319 B.n279 VSUBS 0.007519f
C320 B.n280 VSUBS 0.007519f
C321 B.n281 VSUBS 0.007519f
C322 B.n282 VSUBS 0.007519f
C323 B.n283 VSUBS 0.007519f
C324 B.n284 VSUBS 0.007519f
C325 B.n285 VSUBS 0.007519f
C326 B.n286 VSUBS 0.007519f
C327 B.n287 VSUBS 0.007519f
C328 B.n288 VSUBS 0.007519f
C329 B.n289 VSUBS 0.007519f
C330 B.n290 VSUBS 0.007519f
C331 B.n291 VSUBS 0.007519f
C332 B.n292 VSUBS 0.007519f
C333 B.n293 VSUBS 0.007519f
C334 B.n294 VSUBS 0.007519f
C335 B.n295 VSUBS 0.007519f
C336 B.n296 VSUBS 0.007519f
C337 B.n297 VSUBS 0.007519f
C338 B.n298 VSUBS 0.007519f
C339 B.n299 VSUBS 0.007519f
C340 B.n300 VSUBS 0.007519f
C341 B.n301 VSUBS 0.007519f
C342 B.n302 VSUBS 0.007519f
C343 B.n303 VSUBS 0.007519f
C344 B.n304 VSUBS 0.007519f
C345 B.n305 VSUBS 0.007519f
C346 B.n306 VSUBS 0.007519f
C347 B.n307 VSUBS 0.007519f
C348 B.n308 VSUBS 0.007519f
C349 B.n309 VSUBS 0.007519f
C350 B.n310 VSUBS 0.007519f
C351 B.n311 VSUBS 0.007519f
C352 B.n312 VSUBS 0.007519f
C353 B.n313 VSUBS 0.007519f
C354 B.n314 VSUBS 0.007519f
C355 B.n315 VSUBS 0.017896f
C356 B.n316 VSUBS 0.018372f
C357 B.n317 VSUBS 0.018372f
C358 B.n318 VSUBS 0.007519f
C359 B.n319 VSUBS 0.007519f
C360 B.n320 VSUBS 0.007519f
C361 B.n321 VSUBS 0.007519f
C362 B.n322 VSUBS 0.007519f
C363 B.n323 VSUBS 0.007519f
C364 B.n324 VSUBS 0.007519f
C365 B.n325 VSUBS 0.007519f
C366 B.n326 VSUBS 0.007519f
C367 B.n327 VSUBS 0.007519f
C368 B.n328 VSUBS 0.007519f
C369 B.n329 VSUBS 0.007519f
C370 B.n330 VSUBS 0.007519f
C371 B.n331 VSUBS 0.007519f
C372 B.n332 VSUBS 0.007519f
C373 B.n333 VSUBS 0.007519f
C374 B.n334 VSUBS 0.007519f
C375 B.n335 VSUBS 0.007519f
C376 B.n336 VSUBS 0.007519f
C377 B.n337 VSUBS 0.007519f
C378 B.n338 VSUBS 0.007519f
C379 B.n339 VSUBS 0.007519f
C380 B.n340 VSUBS 0.007519f
C381 B.n341 VSUBS 0.007519f
C382 B.n342 VSUBS 0.007519f
C383 B.n343 VSUBS 0.007519f
C384 B.n344 VSUBS 0.007519f
C385 B.n345 VSUBS 0.007519f
C386 B.n346 VSUBS 0.007519f
C387 B.n347 VSUBS 0.007519f
C388 B.n348 VSUBS 0.007519f
C389 B.n349 VSUBS 0.007519f
C390 B.n350 VSUBS 0.007519f
C391 B.n351 VSUBS 0.007519f
C392 B.n352 VSUBS 0.007519f
C393 B.n353 VSUBS 0.007519f
C394 B.n354 VSUBS 0.007519f
C395 B.n355 VSUBS 0.007519f
C396 B.n356 VSUBS 0.007519f
C397 B.n357 VSUBS 0.007519f
C398 B.n358 VSUBS 0.007519f
C399 B.n359 VSUBS 0.007519f
C400 B.n360 VSUBS 0.007519f
C401 B.n361 VSUBS 0.007519f
C402 B.n362 VSUBS 0.007519f
C403 B.n363 VSUBS 0.007519f
C404 B.n364 VSUBS 0.007519f
C405 B.n365 VSUBS 0.007519f
C406 B.n366 VSUBS 0.007519f
C407 B.n367 VSUBS 0.007519f
C408 B.n368 VSUBS 0.007519f
C409 B.n369 VSUBS 0.007519f
C410 B.n370 VSUBS 0.007519f
C411 B.n371 VSUBS 0.007519f
C412 B.n372 VSUBS 0.007519f
C413 B.n373 VSUBS 0.007519f
C414 B.n374 VSUBS 0.007519f
C415 B.n375 VSUBS 0.007519f
C416 B.n376 VSUBS 0.007519f
C417 B.n377 VSUBS 0.007519f
C418 B.n378 VSUBS 0.007519f
C419 B.n379 VSUBS 0.007519f
C420 B.n380 VSUBS 0.007519f
C421 B.n381 VSUBS 0.007519f
C422 B.n382 VSUBS 0.007519f
C423 B.n383 VSUBS 0.007519f
C424 B.n384 VSUBS 0.007519f
C425 B.n385 VSUBS 0.007519f
C426 B.n386 VSUBS 0.007519f
C427 B.n387 VSUBS 0.007519f
C428 B.n388 VSUBS 0.007519f
C429 B.n389 VSUBS 0.007519f
C430 B.n390 VSUBS 0.007519f
C431 B.n391 VSUBS 0.007519f
C432 B.n392 VSUBS 0.007519f
C433 B.n393 VSUBS 0.007519f
C434 B.n394 VSUBS 0.007519f
C435 B.n395 VSUBS 0.007519f
C436 B.n396 VSUBS 0.005197f
C437 B.n397 VSUBS 0.017421f
C438 B.n398 VSUBS 0.006081f
C439 B.n399 VSUBS 0.007519f
C440 B.n400 VSUBS 0.007519f
C441 B.n401 VSUBS 0.007519f
C442 B.n402 VSUBS 0.007519f
C443 B.n403 VSUBS 0.007519f
C444 B.n404 VSUBS 0.007519f
C445 B.n405 VSUBS 0.007519f
C446 B.n406 VSUBS 0.007519f
C447 B.n407 VSUBS 0.007519f
C448 B.n408 VSUBS 0.007519f
C449 B.n409 VSUBS 0.007519f
C450 B.n410 VSUBS 0.006081f
C451 B.n411 VSUBS 0.007519f
C452 B.n412 VSUBS 0.007519f
C453 B.n413 VSUBS 0.005197f
C454 B.n414 VSUBS 0.007519f
C455 B.n415 VSUBS 0.007519f
C456 B.n416 VSUBS 0.007519f
C457 B.n417 VSUBS 0.007519f
C458 B.n418 VSUBS 0.007519f
C459 B.n419 VSUBS 0.007519f
C460 B.n420 VSUBS 0.007519f
C461 B.n421 VSUBS 0.007519f
C462 B.n422 VSUBS 0.007519f
C463 B.n423 VSUBS 0.007519f
C464 B.n424 VSUBS 0.007519f
C465 B.n425 VSUBS 0.007519f
C466 B.n426 VSUBS 0.007519f
C467 B.n427 VSUBS 0.007519f
C468 B.n428 VSUBS 0.007519f
C469 B.n429 VSUBS 0.007519f
C470 B.n430 VSUBS 0.007519f
C471 B.n431 VSUBS 0.007519f
C472 B.n432 VSUBS 0.007519f
C473 B.n433 VSUBS 0.007519f
C474 B.n434 VSUBS 0.007519f
C475 B.n435 VSUBS 0.007519f
C476 B.n436 VSUBS 0.007519f
C477 B.n437 VSUBS 0.007519f
C478 B.n438 VSUBS 0.007519f
C479 B.n439 VSUBS 0.007519f
C480 B.n440 VSUBS 0.007519f
C481 B.n441 VSUBS 0.007519f
C482 B.n442 VSUBS 0.007519f
C483 B.n443 VSUBS 0.007519f
C484 B.n444 VSUBS 0.007519f
C485 B.n445 VSUBS 0.007519f
C486 B.n446 VSUBS 0.007519f
C487 B.n447 VSUBS 0.007519f
C488 B.n448 VSUBS 0.007519f
C489 B.n449 VSUBS 0.007519f
C490 B.n450 VSUBS 0.007519f
C491 B.n451 VSUBS 0.007519f
C492 B.n452 VSUBS 0.007519f
C493 B.n453 VSUBS 0.007519f
C494 B.n454 VSUBS 0.007519f
C495 B.n455 VSUBS 0.007519f
C496 B.n456 VSUBS 0.007519f
C497 B.n457 VSUBS 0.007519f
C498 B.n458 VSUBS 0.007519f
C499 B.n459 VSUBS 0.007519f
C500 B.n460 VSUBS 0.007519f
C501 B.n461 VSUBS 0.007519f
C502 B.n462 VSUBS 0.007519f
C503 B.n463 VSUBS 0.007519f
C504 B.n464 VSUBS 0.007519f
C505 B.n465 VSUBS 0.007519f
C506 B.n466 VSUBS 0.007519f
C507 B.n467 VSUBS 0.007519f
C508 B.n468 VSUBS 0.007519f
C509 B.n469 VSUBS 0.007519f
C510 B.n470 VSUBS 0.007519f
C511 B.n471 VSUBS 0.007519f
C512 B.n472 VSUBS 0.007519f
C513 B.n473 VSUBS 0.007519f
C514 B.n474 VSUBS 0.007519f
C515 B.n475 VSUBS 0.007519f
C516 B.n476 VSUBS 0.007519f
C517 B.n477 VSUBS 0.007519f
C518 B.n478 VSUBS 0.007519f
C519 B.n479 VSUBS 0.007519f
C520 B.n480 VSUBS 0.007519f
C521 B.n481 VSUBS 0.007519f
C522 B.n482 VSUBS 0.007519f
C523 B.n483 VSUBS 0.007519f
C524 B.n484 VSUBS 0.007519f
C525 B.n485 VSUBS 0.007519f
C526 B.n486 VSUBS 0.007519f
C527 B.n487 VSUBS 0.007519f
C528 B.n488 VSUBS 0.007519f
C529 B.n489 VSUBS 0.007519f
C530 B.n490 VSUBS 0.007519f
C531 B.n491 VSUBS 0.007519f
C532 B.n492 VSUBS 0.017523f
C533 B.n493 VSUBS 0.018745f
C534 B.n494 VSUBS 0.017896f
C535 B.n495 VSUBS 0.007519f
C536 B.n496 VSUBS 0.007519f
C537 B.n497 VSUBS 0.007519f
C538 B.n498 VSUBS 0.007519f
C539 B.n499 VSUBS 0.007519f
C540 B.n500 VSUBS 0.007519f
C541 B.n501 VSUBS 0.007519f
C542 B.n502 VSUBS 0.007519f
C543 B.n503 VSUBS 0.007519f
C544 B.n504 VSUBS 0.007519f
C545 B.n505 VSUBS 0.007519f
C546 B.n506 VSUBS 0.007519f
C547 B.n507 VSUBS 0.007519f
C548 B.n508 VSUBS 0.007519f
C549 B.n509 VSUBS 0.007519f
C550 B.n510 VSUBS 0.007519f
C551 B.n511 VSUBS 0.007519f
C552 B.n512 VSUBS 0.007519f
C553 B.n513 VSUBS 0.007519f
C554 B.n514 VSUBS 0.007519f
C555 B.n515 VSUBS 0.007519f
C556 B.n516 VSUBS 0.007519f
C557 B.n517 VSUBS 0.007519f
C558 B.n518 VSUBS 0.007519f
C559 B.n519 VSUBS 0.007519f
C560 B.n520 VSUBS 0.007519f
C561 B.n521 VSUBS 0.007519f
C562 B.n522 VSUBS 0.007519f
C563 B.n523 VSUBS 0.007519f
C564 B.n524 VSUBS 0.007519f
C565 B.n525 VSUBS 0.007519f
C566 B.n526 VSUBS 0.007519f
C567 B.n527 VSUBS 0.007519f
C568 B.n528 VSUBS 0.007519f
C569 B.n529 VSUBS 0.007519f
C570 B.n530 VSUBS 0.007519f
C571 B.n531 VSUBS 0.007519f
C572 B.n532 VSUBS 0.007519f
C573 B.n533 VSUBS 0.007519f
C574 B.n534 VSUBS 0.007519f
C575 B.n535 VSUBS 0.007519f
C576 B.n536 VSUBS 0.007519f
C577 B.n537 VSUBS 0.007519f
C578 B.n538 VSUBS 0.007519f
C579 B.n539 VSUBS 0.007519f
C580 B.n540 VSUBS 0.007519f
C581 B.n541 VSUBS 0.007519f
C582 B.n542 VSUBS 0.007519f
C583 B.n543 VSUBS 0.007519f
C584 B.n544 VSUBS 0.007519f
C585 B.n545 VSUBS 0.007519f
C586 B.n546 VSUBS 0.007519f
C587 B.n547 VSUBS 0.007519f
C588 B.n548 VSUBS 0.007519f
C589 B.n549 VSUBS 0.007519f
C590 B.n550 VSUBS 0.007519f
C591 B.n551 VSUBS 0.007519f
C592 B.n552 VSUBS 0.007519f
C593 B.n553 VSUBS 0.007519f
C594 B.n554 VSUBS 0.007519f
C595 B.n555 VSUBS 0.007519f
C596 B.n556 VSUBS 0.007519f
C597 B.n557 VSUBS 0.007519f
C598 B.n558 VSUBS 0.007519f
C599 B.n559 VSUBS 0.007519f
C600 B.n560 VSUBS 0.007519f
C601 B.n561 VSUBS 0.007519f
C602 B.n562 VSUBS 0.007519f
C603 B.n563 VSUBS 0.007519f
C604 B.n564 VSUBS 0.007519f
C605 B.n565 VSUBS 0.007519f
C606 B.n566 VSUBS 0.007519f
C607 B.n567 VSUBS 0.007519f
C608 B.n568 VSUBS 0.007519f
C609 B.n569 VSUBS 0.007519f
C610 B.n570 VSUBS 0.007519f
C611 B.n571 VSUBS 0.007519f
C612 B.n572 VSUBS 0.007519f
C613 B.n573 VSUBS 0.007519f
C614 B.n574 VSUBS 0.007519f
C615 B.n575 VSUBS 0.007519f
C616 B.n576 VSUBS 0.007519f
C617 B.n577 VSUBS 0.007519f
C618 B.n578 VSUBS 0.007519f
C619 B.n579 VSUBS 0.007519f
C620 B.n580 VSUBS 0.007519f
C621 B.n581 VSUBS 0.007519f
C622 B.n582 VSUBS 0.007519f
C623 B.n583 VSUBS 0.007519f
C624 B.n584 VSUBS 0.007519f
C625 B.n585 VSUBS 0.007519f
C626 B.n586 VSUBS 0.007519f
C627 B.n587 VSUBS 0.007519f
C628 B.n588 VSUBS 0.007519f
C629 B.n589 VSUBS 0.007519f
C630 B.n590 VSUBS 0.007519f
C631 B.n591 VSUBS 0.007519f
C632 B.n592 VSUBS 0.007519f
C633 B.n593 VSUBS 0.007519f
C634 B.n594 VSUBS 0.007519f
C635 B.n595 VSUBS 0.007519f
C636 B.n596 VSUBS 0.007519f
C637 B.n597 VSUBS 0.007519f
C638 B.n598 VSUBS 0.007519f
C639 B.n599 VSUBS 0.007519f
C640 B.n600 VSUBS 0.007519f
C641 B.n601 VSUBS 0.007519f
C642 B.n602 VSUBS 0.007519f
C643 B.n603 VSUBS 0.007519f
C644 B.n604 VSUBS 0.007519f
C645 B.n605 VSUBS 0.007519f
C646 B.n606 VSUBS 0.007519f
C647 B.n607 VSUBS 0.007519f
C648 B.n608 VSUBS 0.007519f
C649 B.n609 VSUBS 0.007519f
C650 B.n610 VSUBS 0.007519f
C651 B.n611 VSUBS 0.007519f
C652 B.n612 VSUBS 0.007519f
C653 B.n613 VSUBS 0.007519f
C654 B.n614 VSUBS 0.007519f
C655 B.n615 VSUBS 0.007519f
C656 B.n616 VSUBS 0.007519f
C657 B.n617 VSUBS 0.007519f
C658 B.n618 VSUBS 0.007519f
C659 B.n619 VSUBS 0.007519f
C660 B.n620 VSUBS 0.007519f
C661 B.n621 VSUBS 0.007519f
C662 B.n622 VSUBS 0.007519f
C663 B.n623 VSUBS 0.007519f
C664 B.n624 VSUBS 0.007519f
C665 B.n625 VSUBS 0.007519f
C666 B.n626 VSUBS 0.007519f
C667 B.n627 VSUBS 0.007519f
C668 B.n628 VSUBS 0.007519f
C669 B.n629 VSUBS 0.007519f
C670 B.n630 VSUBS 0.007519f
C671 B.n631 VSUBS 0.007519f
C672 B.n632 VSUBS 0.007519f
C673 B.n633 VSUBS 0.007519f
C674 B.n634 VSUBS 0.007519f
C675 B.n635 VSUBS 0.007519f
C676 B.n636 VSUBS 0.007519f
C677 B.n637 VSUBS 0.007519f
C678 B.n638 VSUBS 0.007519f
C679 B.n639 VSUBS 0.007519f
C680 B.n640 VSUBS 0.007519f
C681 B.n641 VSUBS 0.007519f
C682 B.n642 VSUBS 0.007519f
C683 B.n643 VSUBS 0.007519f
C684 B.n644 VSUBS 0.007519f
C685 B.n645 VSUBS 0.007519f
C686 B.n646 VSUBS 0.007519f
C687 B.n647 VSUBS 0.007519f
C688 B.n648 VSUBS 0.007519f
C689 B.n649 VSUBS 0.007519f
C690 B.n650 VSUBS 0.007519f
C691 B.n651 VSUBS 0.007519f
C692 B.n652 VSUBS 0.007519f
C693 B.n653 VSUBS 0.007519f
C694 B.n654 VSUBS 0.007519f
C695 B.n655 VSUBS 0.007519f
C696 B.n656 VSUBS 0.007519f
C697 B.n657 VSUBS 0.017896f
C698 B.n658 VSUBS 0.018372f
C699 B.n659 VSUBS 0.018372f
C700 B.n660 VSUBS 0.007519f
C701 B.n661 VSUBS 0.007519f
C702 B.n662 VSUBS 0.007519f
C703 B.n663 VSUBS 0.007519f
C704 B.n664 VSUBS 0.007519f
C705 B.n665 VSUBS 0.007519f
C706 B.n666 VSUBS 0.007519f
C707 B.n667 VSUBS 0.007519f
C708 B.n668 VSUBS 0.007519f
C709 B.n669 VSUBS 0.007519f
C710 B.n670 VSUBS 0.007519f
C711 B.n671 VSUBS 0.007519f
C712 B.n672 VSUBS 0.007519f
C713 B.n673 VSUBS 0.007519f
C714 B.n674 VSUBS 0.007519f
C715 B.n675 VSUBS 0.007519f
C716 B.n676 VSUBS 0.007519f
C717 B.n677 VSUBS 0.007519f
C718 B.n678 VSUBS 0.007519f
C719 B.n679 VSUBS 0.007519f
C720 B.n680 VSUBS 0.007519f
C721 B.n681 VSUBS 0.007519f
C722 B.n682 VSUBS 0.007519f
C723 B.n683 VSUBS 0.007519f
C724 B.n684 VSUBS 0.007519f
C725 B.n685 VSUBS 0.007519f
C726 B.n686 VSUBS 0.007519f
C727 B.n687 VSUBS 0.007519f
C728 B.n688 VSUBS 0.007519f
C729 B.n689 VSUBS 0.007519f
C730 B.n690 VSUBS 0.007519f
C731 B.n691 VSUBS 0.007519f
C732 B.n692 VSUBS 0.007519f
C733 B.n693 VSUBS 0.007519f
C734 B.n694 VSUBS 0.007519f
C735 B.n695 VSUBS 0.007519f
C736 B.n696 VSUBS 0.007519f
C737 B.n697 VSUBS 0.007519f
C738 B.n698 VSUBS 0.007519f
C739 B.n699 VSUBS 0.007519f
C740 B.n700 VSUBS 0.007519f
C741 B.n701 VSUBS 0.007519f
C742 B.n702 VSUBS 0.007519f
C743 B.n703 VSUBS 0.007519f
C744 B.n704 VSUBS 0.007519f
C745 B.n705 VSUBS 0.007519f
C746 B.n706 VSUBS 0.007519f
C747 B.n707 VSUBS 0.007519f
C748 B.n708 VSUBS 0.007519f
C749 B.n709 VSUBS 0.007519f
C750 B.n710 VSUBS 0.007519f
C751 B.n711 VSUBS 0.007519f
C752 B.n712 VSUBS 0.007519f
C753 B.n713 VSUBS 0.007519f
C754 B.n714 VSUBS 0.007519f
C755 B.n715 VSUBS 0.007519f
C756 B.n716 VSUBS 0.007519f
C757 B.n717 VSUBS 0.007519f
C758 B.n718 VSUBS 0.007519f
C759 B.n719 VSUBS 0.007519f
C760 B.n720 VSUBS 0.007519f
C761 B.n721 VSUBS 0.007519f
C762 B.n722 VSUBS 0.007519f
C763 B.n723 VSUBS 0.007519f
C764 B.n724 VSUBS 0.007519f
C765 B.n725 VSUBS 0.007519f
C766 B.n726 VSUBS 0.007519f
C767 B.n727 VSUBS 0.007519f
C768 B.n728 VSUBS 0.007519f
C769 B.n729 VSUBS 0.007519f
C770 B.n730 VSUBS 0.007519f
C771 B.n731 VSUBS 0.007519f
C772 B.n732 VSUBS 0.007519f
C773 B.n733 VSUBS 0.007519f
C774 B.n734 VSUBS 0.007519f
C775 B.n735 VSUBS 0.007519f
C776 B.n736 VSUBS 0.007519f
C777 B.n737 VSUBS 0.007519f
C778 B.n738 VSUBS 0.005197f
C779 B.n739 VSUBS 0.017421f
C780 B.n740 VSUBS 0.006081f
C781 B.n741 VSUBS 0.007519f
C782 B.n742 VSUBS 0.007519f
C783 B.n743 VSUBS 0.007519f
C784 B.n744 VSUBS 0.007519f
C785 B.n745 VSUBS 0.007519f
C786 B.n746 VSUBS 0.007519f
C787 B.n747 VSUBS 0.007519f
C788 B.n748 VSUBS 0.007519f
C789 B.n749 VSUBS 0.007519f
C790 B.n750 VSUBS 0.007519f
C791 B.n751 VSUBS 0.007519f
C792 B.n752 VSUBS 0.006081f
C793 B.n753 VSUBS 0.007519f
C794 B.n754 VSUBS 0.007519f
C795 B.n755 VSUBS 0.005197f
C796 B.n756 VSUBS 0.007519f
C797 B.n757 VSUBS 0.007519f
C798 B.n758 VSUBS 0.007519f
C799 B.n759 VSUBS 0.007519f
C800 B.n760 VSUBS 0.007519f
C801 B.n761 VSUBS 0.007519f
C802 B.n762 VSUBS 0.007519f
C803 B.n763 VSUBS 0.007519f
C804 B.n764 VSUBS 0.007519f
C805 B.n765 VSUBS 0.007519f
C806 B.n766 VSUBS 0.007519f
C807 B.n767 VSUBS 0.007519f
C808 B.n768 VSUBS 0.007519f
C809 B.n769 VSUBS 0.007519f
C810 B.n770 VSUBS 0.007519f
C811 B.n771 VSUBS 0.007519f
C812 B.n772 VSUBS 0.007519f
C813 B.n773 VSUBS 0.007519f
C814 B.n774 VSUBS 0.007519f
C815 B.n775 VSUBS 0.007519f
C816 B.n776 VSUBS 0.007519f
C817 B.n777 VSUBS 0.007519f
C818 B.n778 VSUBS 0.007519f
C819 B.n779 VSUBS 0.007519f
C820 B.n780 VSUBS 0.007519f
C821 B.n781 VSUBS 0.007519f
C822 B.n782 VSUBS 0.007519f
C823 B.n783 VSUBS 0.007519f
C824 B.n784 VSUBS 0.007519f
C825 B.n785 VSUBS 0.007519f
C826 B.n786 VSUBS 0.007519f
C827 B.n787 VSUBS 0.007519f
C828 B.n788 VSUBS 0.007519f
C829 B.n789 VSUBS 0.007519f
C830 B.n790 VSUBS 0.007519f
C831 B.n791 VSUBS 0.007519f
C832 B.n792 VSUBS 0.007519f
C833 B.n793 VSUBS 0.007519f
C834 B.n794 VSUBS 0.007519f
C835 B.n795 VSUBS 0.007519f
C836 B.n796 VSUBS 0.007519f
C837 B.n797 VSUBS 0.007519f
C838 B.n798 VSUBS 0.007519f
C839 B.n799 VSUBS 0.007519f
C840 B.n800 VSUBS 0.007519f
C841 B.n801 VSUBS 0.007519f
C842 B.n802 VSUBS 0.007519f
C843 B.n803 VSUBS 0.007519f
C844 B.n804 VSUBS 0.007519f
C845 B.n805 VSUBS 0.007519f
C846 B.n806 VSUBS 0.007519f
C847 B.n807 VSUBS 0.007519f
C848 B.n808 VSUBS 0.007519f
C849 B.n809 VSUBS 0.007519f
C850 B.n810 VSUBS 0.007519f
C851 B.n811 VSUBS 0.007519f
C852 B.n812 VSUBS 0.007519f
C853 B.n813 VSUBS 0.007519f
C854 B.n814 VSUBS 0.007519f
C855 B.n815 VSUBS 0.007519f
C856 B.n816 VSUBS 0.007519f
C857 B.n817 VSUBS 0.007519f
C858 B.n818 VSUBS 0.007519f
C859 B.n819 VSUBS 0.007519f
C860 B.n820 VSUBS 0.007519f
C861 B.n821 VSUBS 0.007519f
C862 B.n822 VSUBS 0.007519f
C863 B.n823 VSUBS 0.007519f
C864 B.n824 VSUBS 0.007519f
C865 B.n825 VSUBS 0.007519f
C866 B.n826 VSUBS 0.007519f
C867 B.n827 VSUBS 0.007519f
C868 B.n828 VSUBS 0.007519f
C869 B.n829 VSUBS 0.007519f
C870 B.n830 VSUBS 0.007519f
C871 B.n831 VSUBS 0.007519f
C872 B.n832 VSUBS 0.007519f
C873 B.n833 VSUBS 0.007519f
C874 B.n834 VSUBS 0.018372f
C875 B.n835 VSUBS 0.017896f
C876 B.n836 VSUBS 0.017896f
C877 B.n837 VSUBS 0.007519f
C878 B.n838 VSUBS 0.007519f
C879 B.n839 VSUBS 0.007519f
C880 B.n840 VSUBS 0.007519f
C881 B.n841 VSUBS 0.007519f
C882 B.n842 VSUBS 0.007519f
C883 B.n843 VSUBS 0.007519f
C884 B.n844 VSUBS 0.007519f
C885 B.n845 VSUBS 0.007519f
C886 B.n846 VSUBS 0.007519f
C887 B.n847 VSUBS 0.007519f
C888 B.n848 VSUBS 0.007519f
C889 B.n849 VSUBS 0.007519f
C890 B.n850 VSUBS 0.007519f
C891 B.n851 VSUBS 0.007519f
C892 B.n852 VSUBS 0.007519f
C893 B.n853 VSUBS 0.007519f
C894 B.n854 VSUBS 0.007519f
C895 B.n855 VSUBS 0.007519f
C896 B.n856 VSUBS 0.007519f
C897 B.n857 VSUBS 0.007519f
C898 B.n858 VSUBS 0.007519f
C899 B.n859 VSUBS 0.007519f
C900 B.n860 VSUBS 0.007519f
C901 B.n861 VSUBS 0.007519f
C902 B.n862 VSUBS 0.007519f
C903 B.n863 VSUBS 0.007519f
C904 B.n864 VSUBS 0.007519f
C905 B.n865 VSUBS 0.007519f
C906 B.n866 VSUBS 0.007519f
C907 B.n867 VSUBS 0.007519f
C908 B.n868 VSUBS 0.007519f
C909 B.n869 VSUBS 0.007519f
C910 B.n870 VSUBS 0.007519f
C911 B.n871 VSUBS 0.007519f
C912 B.n872 VSUBS 0.007519f
C913 B.n873 VSUBS 0.007519f
C914 B.n874 VSUBS 0.007519f
C915 B.n875 VSUBS 0.007519f
C916 B.n876 VSUBS 0.007519f
C917 B.n877 VSUBS 0.007519f
C918 B.n878 VSUBS 0.007519f
C919 B.n879 VSUBS 0.007519f
C920 B.n880 VSUBS 0.007519f
C921 B.n881 VSUBS 0.007519f
C922 B.n882 VSUBS 0.007519f
C923 B.n883 VSUBS 0.007519f
C924 B.n884 VSUBS 0.007519f
C925 B.n885 VSUBS 0.007519f
C926 B.n886 VSUBS 0.007519f
C927 B.n887 VSUBS 0.007519f
C928 B.n888 VSUBS 0.007519f
C929 B.n889 VSUBS 0.007519f
C930 B.n890 VSUBS 0.007519f
C931 B.n891 VSUBS 0.007519f
C932 B.n892 VSUBS 0.007519f
C933 B.n893 VSUBS 0.007519f
C934 B.n894 VSUBS 0.007519f
C935 B.n895 VSUBS 0.007519f
C936 B.n896 VSUBS 0.007519f
C937 B.n897 VSUBS 0.007519f
C938 B.n898 VSUBS 0.007519f
C939 B.n899 VSUBS 0.007519f
C940 B.n900 VSUBS 0.007519f
C941 B.n901 VSUBS 0.007519f
C942 B.n902 VSUBS 0.007519f
C943 B.n903 VSUBS 0.007519f
C944 B.n904 VSUBS 0.007519f
C945 B.n905 VSUBS 0.007519f
C946 B.n906 VSUBS 0.007519f
C947 B.n907 VSUBS 0.007519f
C948 B.n908 VSUBS 0.007519f
C949 B.n909 VSUBS 0.007519f
C950 B.n910 VSUBS 0.007519f
C951 B.n911 VSUBS 0.007519f
C952 B.n912 VSUBS 0.007519f
C953 B.n913 VSUBS 0.007519f
C954 B.n914 VSUBS 0.007519f
C955 B.n915 VSUBS 0.009812f
C956 B.n916 VSUBS 0.010452f
C957 B.n917 VSUBS 0.020785f
C958 VDD2.n0 VSUBS 0.029911f
C959 VDD2.n1 VSUBS 0.027539f
C960 VDD2.n2 VSUBS 0.014798f
C961 VDD2.n3 VSUBS 0.034978f
C962 VDD2.n4 VSUBS 0.015669f
C963 VDD2.n5 VSUBS 0.027539f
C964 VDD2.n6 VSUBS 0.015233f
C965 VDD2.n7 VSUBS 0.034978f
C966 VDD2.n8 VSUBS 0.015669f
C967 VDD2.n9 VSUBS 0.027539f
C968 VDD2.n10 VSUBS 0.014798f
C969 VDD2.n11 VSUBS 0.034978f
C970 VDD2.n12 VSUBS 0.015669f
C971 VDD2.n13 VSUBS 0.027539f
C972 VDD2.n14 VSUBS 0.014798f
C973 VDD2.n15 VSUBS 0.034978f
C974 VDD2.n16 VSUBS 0.015669f
C975 VDD2.n17 VSUBS 0.027539f
C976 VDD2.n18 VSUBS 0.014798f
C977 VDD2.n19 VSUBS 0.034978f
C978 VDD2.n20 VSUBS 0.015669f
C979 VDD2.n21 VSUBS 0.027539f
C980 VDD2.n22 VSUBS 0.014798f
C981 VDD2.n23 VSUBS 0.034978f
C982 VDD2.n24 VSUBS 0.015669f
C983 VDD2.n25 VSUBS 0.027539f
C984 VDD2.n26 VSUBS 0.014798f
C985 VDD2.n27 VSUBS 0.026233f
C986 VDD2.n28 VSUBS 0.022251f
C987 VDD2.t0 VSUBS 0.074961f
C988 VDD2.n29 VSUBS 0.203711f
C989 VDD2.n30 VSUBS 1.90595f
C990 VDD2.n31 VSUBS 0.014798f
C991 VDD2.n32 VSUBS 0.015669f
C992 VDD2.n33 VSUBS 0.034978f
C993 VDD2.n34 VSUBS 0.034978f
C994 VDD2.n35 VSUBS 0.015669f
C995 VDD2.n36 VSUBS 0.014798f
C996 VDD2.n37 VSUBS 0.027539f
C997 VDD2.n38 VSUBS 0.027539f
C998 VDD2.n39 VSUBS 0.014798f
C999 VDD2.n40 VSUBS 0.015669f
C1000 VDD2.n41 VSUBS 0.034978f
C1001 VDD2.n42 VSUBS 0.034978f
C1002 VDD2.n43 VSUBS 0.015669f
C1003 VDD2.n44 VSUBS 0.014798f
C1004 VDD2.n45 VSUBS 0.027539f
C1005 VDD2.n46 VSUBS 0.027539f
C1006 VDD2.n47 VSUBS 0.014798f
C1007 VDD2.n48 VSUBS 0.015669f
C1008 VDD2.n49 VSUBS 0.034978f
C1009 VDD2.n50 VSUBS 0.034978f
C1010 VDD2.n51 VSUBS 0.015669f
C1011 VDD2.n52 VSUBS 0.014798f
C1012 VDD2.n53 VSUBS 0.027539f
C1013 VDD2.n54 VSUBS 0.027539f
C1014 VDD2.n55 VSUBS 0.014798f
C1015 VDD2.n56 VSUBS 0.015669f
C1016 VDD2.n57 VSUBS 0.034978f
C1017 VDD2.n58 VSUBS 0.034978f
C1018 VDD2.n59 VSUBS 0.015669f
C1019 VDD2.n60 VSUBS 0.014798f
C1020 VDD2.n61 VSUBS 0.027539f
C1021 VDD2.n62 VSUBS 0.027539f
C1022 VDD2.n63 VSUBS 0.014798f
C1023 VDD2.n64 VSUBS 0.015669f
C1024 VDD2.n65 VSUBS 0.034978f
C1025 VDD2.n66 VSUBS 0.034978f
C1026 VDD2.n67 VSUBS 0.015669f
C1027 VDD2.n68 VSUBS 0.014798f
C1028 VDD2.n69 VSUBS 0.027539f
C1029 VDD2.n70 VSUBS 0.027539f
C1030 VDD2.n71 VSUBS 0.014798f
C1031 VDD2.n72 VSUBS 0.014798f
C1032 VDD2.n73 VSUBS 0.015669f
C1033 VDD2.n74 VSUBS 0.034978f
C1034 VDD2.n75 VSUBS 0.034978f
C1035 VDD2.n76 VSUBS 0.034978f
C1036 VDD2.n77 VSUBS 0.015233f
C1037 VDD2.n78 VSUBS 0.014798f
C1038 VDD2.n79 VSUBS 0.027539f
C1039 VDD2.n80 VSUBS 0.027539f
C1040 VDD2.n81 VSUBS 0.014798f
C1041 VDD2.n82 VSUBS 0.015669f
C1042 VDD2.n83 VSUBS 0.034978f
C1043 VDD2.n84 VSUBS 0.08349f
C1044 VDD2.n85 VSUBS 0.015669f
C1045 VDD2.n86 VSUBS 0.014798f
C1046 VDD2.n87 VSUBS 0.067417f
C1047 VDD2.n88 VSUBS 0.073966f
C1048 VDD2.t5 VSUBS 0.352112f
C1049 VDD2.t4 VSUBS 0.352112f
C1050 VDD2.n89 VSUBS 2.90432f
C1051 VDD2.n90 VSUBS 4.01732f
C1052 VDD2.n91 VSUBS 0.029911f
C1053 VDD2.n92 VSUBS 0.027539f
C1054 VDD2.n93 VSUBS 0.014798f
C1055 VDD2.n94 VSUBS 0.034978f
C1056 VDD2.n95 VSUBS 0.015669f
C1057 VDD2.n96 VSUBS 0.027539f
C1058 VDD2.n97 VSUBS 0.015233f
C1059 VDD2.n98 VSUBS 0.034978f
C1060 VDD2.n99 VSUBS 0.014798f
C1061 VDD2.n100 VSUBS 0.015669f
C1062 VDD2.n101 VSUBS 0.027539f
C1063 VDD2.n102 VSUBS 0.014798f
C1064 VDD2.n103 VSUBS 0.034978f
C1065 VDD2.n104 VSUBS 0.015669f
C1066 VDD2.n105 VSUBS 0.027539f
C1067 VDD2.n106 VSUBS 0.014798f
C1068 VDD2.n107 VSUBS 0.034978f
C1069 VDD2.n108 VSUBS 0.015669f
C1070 VDD2.n109 VSUBS 0.027539f
C1071 VDD2.n110 VSUBS 0.014798f
C1072 VDD2.n111 VSUBS 0.034978f
C1073 VDD2.n112 VSUBS 0.015669f
C1074 VDD2.n113 VSUBS 0.027539f
C1075 VDD2.n114 VSUBS 0.014798f
C1076 VDD2.n115 VSUBS 0.034978f
C1077 VDD2.n116 VSUBS 0.015669f
C1078 VDD2.n117 VSUBS 0.027539f
C1079 VDD2.n118 VSUBS 0.014798f
C1080 VDD2.n119 VSUBS 0.026233f
C1081 VDD2.n120 VSUBS 0.022251f
C1082 VDD2.t2 VSUBS 0.074961f
C1083 VDD2.n121 VSUBS 0.203711f
C1084 VDD2.n122 VSUBS 1.90595f
C1085 VDD2.n123 VSUBS 0.014798f
C1086 VDD2.n124 VSUBS 0.015669f
C1087 VDD2.n125 VSUBS 0.034978f
C1088 VDD2.n126 VSUBS 0.034978f
C1089 VDD2.n127 VSUBS 0.015669f
C1090 VDD2.n128 VSUBS 0.014798f
C1091 VDD2.n129 VSUBS 0.027539f
C1092 VDD2.n130 VSUBS 0.027539f
C1093 VDD2.n131 VSUBS 0.014798f
C1094 VDD2.n132 VSUBS 0.015669f
C1095 VDD2.n133 VSUBS 0.034978f
C1096 VDD2.n134 VSUBS 0.034978f
C1097 VDD2.n135 VSUBS 0.015669f
C1098 VDD2.n136 VSUBS 0.014798f
C1099 VDD2.n137 VSUBS 0.027539f
C1100 VDD2.n138 VSUBS 0.027539f
C1101 VDD2.n139 VSUBS 0.014798f
C1102 VDD2.n140 VSUBS 0.015669f
C1103 VDD2.n141 VSUBS 0.034978f
C1104 VDD2.n142 VSUBS 0.034978f
C1105 VDD2.n143 VSUBS 0.015669f
C1106 VDD2.n144 VSUBS 0.014798f
C1107 VDD2.n145 VSUBS 0.027539f
C1108 VDD2.n146 VSUBS 0.027539f
C1109 VDD2.n147 VSUBS 0.014798f
C1110 VDD2.n148 VSUBS 0.015669f
C1111 VDD2.n149 VSUBS 0.034978f
C1112 VDD2.n150 VSUBS 0.034978f
C1113 VDD2.n151 VSUBS 0.015669f
C1114 VDD2.n152 VSUBS 0.014798f
C1115 VDD2.n153 VSUBS 0.027539f
C1116 VDD2.n154 VSUBS 0.027539f
C1117 VDD2.n155 VSUBS 0.014798f
C1118 VDD2.n156 VSUBS 0.015669f
C1119 VDD2.n157 VSUBS 0.034978f
C1120 VDD2.n158 VSUBS 0.034978f
C1121 VDD2.n159 VSUBS 0.015669f
C1122 VDD2.n160 VSUBS 0.014798f
C1123 VDD2.n161 VSUBS 0.027539f
C1124 VDD2.n162 VSUBS 0.027539f
C1125 VDD2.n163 VSUBS 0.014798f
C1126 VDD2.n164 VSUBS 0.015669f
C1127 VDD2.n165 VSUBS 0.034978f
C1128 VDD2.n166 VSUBS 0.034978f
C1129 VDD2.n167 VSUBS 0.034978f
C1130 VDD2.n168 VSUBS 0.015233f
C1131 VDD2.n169 VSUBS 0.014798f
C1132 VDD2.n170 VSUBS 0.027539f
C1133 VDD2.n171 VSUBS 0.027539f
C1134 VDD2.n172 VSUBS 0.014798f
C1135 VDD2.n173 VSUBS 0.015669f
C1136 VDD2.n174 VSUBS 0.034978f
C1137 VDD2.n175 VSUBS 0.08349f
C1138 VDD2.n176 VSUBS 0.015669f
C1139 VDD2.n177 VSUBS 0.014798f
C1140 VDD2.n178 VSUBS 0.067417f
C1141 VDD2.n179 VSUBS 0.061033f
C1142 VDD2.n180 VSUBS 3.47904f
C1143 VDD2.t1 VSUBS 0.352112f
C1144 VDD2.t3 VSUBS 0.352112f
C1145 VDD2.n181 VSUBS 2.90427f
C1146 VN.t1 VSUBS 3.72069f
C1147 VN.n0 VSUBS 1.37812f
C1148 VN.n1 VSUBS 0.023208f
C1149 VN.n2 VSUBS 0.035663f
C1150 VN.n3 VSUBS 0.023208f
C1151 VN.n4 VSUBS 0.032414f
C1152 VN.t0 VSUBS 3.72069f
C1153 VN.n5 VSUBS 1.36774f
C1154 VN.t5 VSUBS 4.066f
C1155 VN.n6 VSUBS 1.30143f
C1156 VN.n7 VSUBS 0.289911f
C1157 VN.n8 VSUBS 0.023208f
C1158 VN.n9 VSUBS 0.043037f
C1159 VN.n10 VSUBS 0.043037f
C1160 VN.n11 VSUBS 0.03181f
C1161 VN.n12 VSUBS 0.023208f
C1162 VN.n13 VSUBS 0.023208f
C1163 VN.n14 VSUBS 0.023208f
C1164 VN.n15 VSUBS 0.043037f
C1165 VN.n16 VSUBS 0.043037f
C1166 VN.n17 VSUBS 0.029864f
C1167 VN.n18 VSUBS 0.037451f
C1168 VN.n19 VSUBS 0.06406f
C1169 VN.t3 VSUBS 3.72069f
C1170 VN.n20 VSUBS 1.37812f
C1171 VN.n21 VSUBS 0.023208f
C1172 VN.n22 VSUBS 0.035663f
C1173 VN.n23 VSUBS 0.023208f
C1174 VN.n24 VSUBS 0.032414f
C1175 VN.t2 VSUBS 4.066f
C1176 VN.t4 VSUBS 3.72069f
C1177 VN.n25 VSUBS 1.36774f
C1178 VN.n26 VSUBS 1.30143f
C1179 VN.n27 VSUBS 0.289911f
C1180 VN.n28 VSUBS 0.023208f
C1181 VN.n29 VSUBS 0.043037f
C1182 VN.n30 VSUBS 0.043037f
C1183 VN.n31 VSUBS 0.03181f
C1184 VN.n32 VSUBS 0.023208f
C1185 VN.n33 VSUBS 0.023208f
C1186 VN.n34 VSUBS 0.023208f
C1187 VN.n35 VSUBS 0.043037f
C1188 VN.n36 VSUBS 0.043037f
C1189 VN.n37 VSUBS 0.029864f
C1190 VN.n38 VSUBS 0.037451f
C1191 VN.n39 VSUBS 1.56215f
C1192 VDD1.n0 VSUBS 0.029909f
C1193 VDD1.n1 VSUBS 0.027537f
C1194 VDD1.n2 VSUBS 0.014797f
C1195 VDD1.n3 VSUBS 0.034975f
C1196 VDD1.n4 VSUBS 0.015668f
C1197 VDD1.n5 VSUBS 0.027537f
C1198 VDD1.n6 VSUBS 0.015232f
C1199 VDD1.n7 VSUBS 0.034975f
C1200 VDD1.n8 VSUBS 0.014797f
C1201 VDD1.n9 VSUBS 0.015668f
C1202 VDD1.n10 VSUBS 0.027537f
C1203 VDD1.n11 VSUBS 0.014797f
C1204 VDD1.n12 VSUBS 0.034975f
C1205 VDD1.n13 VSUBS 0.015668f
C1206 VDD1.n14 VSUBS 0.027537f
C1207 VDD1.n15 VSUBS 0.014797f
C1208 VDD1.n16 VSUBS 0.034975f
C1209 VDD1.n17 VSUBS 0.015668f
C1210 VDD1.n18 VSUBS 0.027537f
C1211 VDD1.n19 VSUBS 0.014797f
C1212 VDD1.n20 VSUBS 0.034975f
C1213 VDD1.n21 VSUBS 0.015668f
C1214 VDD1.n22 VSUBS 0.027537f
C1215 VDD1.n23 VSUBS 0.014797f
C1216 VDD1.n24 VSUBS 0.034975f
C1217 VDD1.n25 VSUBS 0.015668f
C1218 VDD1.n26 VSUBS 0.027537f
C1219 VDD1.n27 VSUBS 0.014797f
C1220 VDD1.n28 VSUBS 0.026231f
C1221 VDD1.n29 VSUBS 0.02225f
C1222 VDD1.t5 VSUBS 0.074956f
C1223 VDD1.n30 VSUBS 0.203697f
C1224 VDD1.n31 VSUBS 1.90581f
C1225 VDD1.n32 VSUBS 0.014797f
C1226 VDD1.n33 VSUBS 0.015668f
C1227 VDD1.n34 VSUBS 0.034975f
C1228 VDD1.n35 VSUBS 0.034975f
C1229 VDD1.n36 VSUBS 0.015668f
C1230 VDD1.n37 VSUBS 0.014797f
C1231 VDD1.n38 VSUBS 0.027537f
C1232 VDD1.n39 VSUBS 0.027537f
C1233 VDD1.n40 VSUBS 0.014797f
C1234 VDD1.n41 VSUBS 0.015668f
C1235 VDD1.n42 VSUBS 0.034975f
C1236 VDD1.n43 VSUBS 0.034975f
C1237 VDD1.n44 VSUBS 0.015668f
C1238 VDD1.n45 VSUBS 0.014797f
C1239 VDD1.n46 VSUBS 0.027537f
C1240 VDD1.n47 VSUBS 0.027537f
C1241 VDD1.n48 VSUBS 0.014797f
C1242 VDD1.n49 VSUBS 0.015668f
C1243 VDD1.n50 VSUBS 0.034975f
C1244 VDD1.n51 VSUBS 0.034975f
C1245 VDD1.n52 VSUBS 0.015668f
C1246 VDD1.n53 VSUBS 0.014797f
C1247 VDD1.n54 VSUBS 0.027537f
C1248 VDD1.n55 VSUBS 0.027537f
C1249 VDD1.n56 VSUBS 0.014797f
C1250 VDD1.n57 VSUBS 0.015668f
C1251 VDD1.n58 VSUBS 0.034975f
C1252 VDD1.n59 VSUBS 0.034975f
C1253 VDD1.n60 VSUBS 0.015668f
C1254 VDD1.n61 VSUBS 0.014797f
C1255 VDD1.n62 VSUBS 0.027537f
C1256 VDD1.n63 VSUBS 0.027537f
C1257 VDD1.n64 VSUBS 0.014797f
C1258 VDD1.n65 VSUBS 0.015668f
C1259 VDD1.n66 VSUBS 0.034975f
C1260 VDD1.n67 VSUBS 0.034975f
C1261 VDD1.n68 VSUBS 0.015668f
C1262 VDD1.n69 VSUBS 0.014797f
C1263 VDD1.n70 VSUBS 0.027537f
C1264 VDD1.n71 VSUBS 0.027537f
C1265 VDD1.n72 VSUBS 0.014797f
C1266 VDD1.n73 VSUBS 0.015668f
C1267 VDD1.n74 VSUBS 0.034975f
C1268 VDD1.n75 VSUBS 0.034975f
C1269 VDD1.n76 VSUBS 0.034975f
C1270 VDD1.n77 VSUBS 0.015232f
C1271 VDD1.n78 VSUBS 0.014797f
C1272 VDD1.n79 VSUBS 0.027537f
C1273 VDD1.n80 VSUBS 0.027537f
C1274 VDD1.n81 VSUBS 0.014797f
C1275 VDD1.n82 VSUBS 0.015668f
C1276 VDD1.n83 VSUBS 0.034975f
C1277 VDD1.n84 VSUBS 0.083484f
C1278 VDD1.n85 VSUBS 0.015668f
C1279 VDD1.n86 VSUBS 0.014797f
C1280 VDD1.n87 VSUBS 0.067413f
C1281 VDD1.n88 VSUBS 0.075f
C1282 VDD1.n89 VSUBS 0.029909f
C1283 VDD1.n90 VSUBS 0.027537f
C1284 VDD1.n91 VSUBS 0.014797f
C1285 VDD1.n92 VSUBS 0.034975f
C1286 VDD1.n93 VSUBS 0.015668f
C1287 VDD1.n94 VSUBS 0.027537f
C1288 VDD1.n95 VSUBS 0.015232f
C1289 VDD1.n96 VSUBS 0.034975f
C1290 VDD1.n97 VSUBS 0.015668f
C1291 VDD1.n98 VSUBS 0.027537f
C1292 VDD1.n99 VSUBS 0.014797f
C1293 VDD1.n100 VSUBS 0.034975f
C1294 VDD1.n101 VSUBS 0.015668f
C1295 VDD1.n102 VSUBS 0.027537f
C1296 VDD1.n103 VSUBS 0.014797f
C1297 VDD1.n104 VSUBS 0.034975f
C1298 VDD1.n105 VSUBS 0.015668f
C1299 VDD1.n106 VSUBS 0.027537f
C1300 VDD1.n107 VSUBS 0.014797f
C1301 VDD1.n108 VSUBS 0.034975f
C1302 VDD1.n109 VSUBS 0.015668f
C1303 VDD1.n110 VSUBS 0.027537f
C1304 VDD1.n111 VSUBS 0.014797f
C1305 VDD1.n112 VSUBS 0.034975f
C1306 VDD1.n113 VSUBS 0.015668f
C1307 VDD1.n114 VSUBS 0.027537f
C1308 VDD1.n115 VSUBS 0.014797f
C1309 VDD1.n116 VSUBS 0.026231f
C1310 VDD1.n117 VSUBS 0.02225f
C1311 VDD1.t1 VSUBS 0.074956f
C1312 VDD1.n118 VSUBS 0.203697f
C1313 VDD1.n119 VSUBS 1.90581f
C1314 VDD1.n120 VSUBS 0.014797f
C1315 VDD1.n121 VSUBS 0.015668f
C1316 VDD1.n122 VSUBS 0.034975f
C1317 VDD1.n123 VSUBS 0.034975f
C1318 VDD1.n124 VSUBS 0.015668f
C1319 VDD1.n125 VSUBS 0.014797f
C1320 VDD1.n126 VSUBS 0.027537f
C1321 VDD1.n127 VSUBS 0.027537f
C1322 VDD1.n128 VSUBS 0.014797f
C1323 VDD1.n129 VSUBS 0.015668f
C1324 VDD1.n130 VSUBS 0.034975f
C1325 VDD1.n131 VSUBS 0.034975f
C1326 VDD1.n132 VSUBS 0.015668f
C1327 VDD1.n133 VSUBS 0.014797f
C1328 VDD1.n134 VSUBS 0.027537f
C1329 VDD1.n135 VSUBS 0.027537f
C1330 VDD1.n136 VSUBS 0.014797f
C1331 VDD1.n137 VSUBS 0.015668f
C1332 VDD1.n138 VSUBS 0.034975f
C1333 VDD1.n139 VSUBS 0.034975f
C1334 VDD1.n140 VSUBS 0.015668f
C1335 VDD1.n141 VSUBS 0.014797f
C1336 VDD1.n142 VSUBS 0.027537f
C1337 VDD1.n143 VSUBS 0.027537f
C1338 VDD1.n144 VSUBS 0.014797f
C1339 VDD1.n145 VSUBS 0.015668f
C1340 VDD1.n146 VSUBS 0.034975f
C1341 VDD1.n147 VSUBS 0.034975f
C1342 VDD1.n148 VSUBS 0.015668f
C1343 VDD1.n149 VSUBS 0.014797f
C1344 VDD1.n150 VSUBS 0.027537f
C1345 VDD1.n151 VSUBS 0.027537f
C1346 VDD1.n152 VSUBS 0.014797f
C1347 VDD1.n153 VSUBS 0.015668f
C1348 VDD1.n154 VSUBS 0.034975f
C1349 VDD1.n155 VSUBS 0.034975f
C1350 VDD1.n156 VSUBS 0.015668f
C1351 VDD1.n157 VSUBS 0.014797f
C1352 VDD1.n158 VSUBS 0.027537f
C1353 VDD1.n159 VSUBS 0.027537f
C1354 VDD1.n160 VSUBS 0.014797f
C1355 VDD1.n161 VSUBS 0.014797f
C1356 VDD1.n162 VSUBS 0.015668f
C1357 VDD1.n163 VSUBS 0.034975f
C1358 VDD1.n164 VSUBS 0.034975f
C1359 VDD1.n165 VSUBS 0.034975f
C1360 VDD1.n166 VSUBS 0.015232f
C1361 VDD1.n167 VSUBS 0.014797f
C1362 VDD1.n168 VSUBS 0.027537f
C1363 VDD1.n169 VSUBS 0.027537f
C1364 VDD1.n170 VSUBS 0.014797f
C1365 VDD1.n171 VSUBS 0.015668f
C1366 VDD1.n172 VSUBS 0.034975f
C1367 VDD1.n173 VSUBS 0.083484f
C1368 VDD1.n174 VSUBS 0.015668f
C1369 VDD1.n175 VSUBS 0.014797f
C1370 VDD1.n176 VSUBS 0.067413f
C1371 VDD1.n177 VSUBS 0.073961f
C1372 VDD1.t2 VSUBS 0.352088f
C1373 VDD1.t4 VSUBS 0.352088f
C1374 VDD1.n178 VSUBS 2.90412f
C1375 VDD1.n179 VSUBS 4.18722f
C1376 VDD1.t3 VSUBS 0.352088f
C1377 VDD1.t0 VSUBS 0.352088f
C1378 VDD1.n180 VSUBS 2.89416f
C1379 VDD1.n181 VSUBS 4.03269f
C1380 VTAIL.t1 VSUBS 0.364908f
C1381 VTAIL.t3 VSUBS 0.364908f
C1382 VTAIL.n0 VSUBS 2.83604f
C1383 VTAIL.n1 VSUBS 0.95277f
C1384 VTAIL.n2 VSUBS 0.030998f
C1385 VTAIL.n3 VSUBS 0.02854f
C1386 VTAIL.n4 VSUBS 0.015336f
C1387 VTAIL.n5 VSUBS 0.036249f
C1388 VTAIL.n6 VSUBS 0.016238f
C1389 VTAIL.n7 VSUBS 0.02854f
C1390 VTAIL.n8 VSUBS 0.015787f
C1391 VTAIL.n9 VSUBS 0.036249f
C1392 VTAIL.n10 VSUBS 0.016238f
C1393 VTAIL.n11 VSUBS 0.02854f
C1394 VTAIL.n12 VSUBS 0.015336f
C1395 VTAIL.n13 VSUBS 0.036249f
C1396 VTAIL.n14 VSUBS 0.016238f
C1397 VTAIL.n15 VSUBS 0.02854f
C1398 VTAIL.n16 VSUBS 0.015336f
C1399 VTAIL.n17 VSUBS 0.036249f
C1400 VTAIL.n18 VSUBS 0.016238f
C1401 VTAIL.n19 VSUBS 0.02854f
C1402 VTAIL.n20 VSUBS 0.015336f
C1403 VTAIL.n21 VSUBS 0.036249f
C1404 VTAIL.n22 VSUBS 0.016238f
C1405 VTAIL.n23 VSUBS 0.02854f
C1406 VTAIL.n24 VSUBS 0.015336f
C1407 VTAIL.n25 VSUBS 0.036249f
C1408 VTAIL.n26 VSUBS 0.016238f
C1409 VTAIL.n27 VSUBS 0.02854f
C1410 VTAIL.n28 VSUBS 0.015336f
C1411 VTAIL.n29 VSUBS 0.027187f
C1412 VTAIL.n30 VSUBS 0.02306f
C1413 VTAIL.t10 VSUBS 0.077685f
C1414 VTAIL.n31 VSUBS 0.211114f
C1415 VTAIL.n32 VSUBS 1.97521f
C1416 VTAIL.n33 VSUBS 0.015336f
C1417 VTAIL.n34 VSUBS 0.016238f
C1418 VTAIL.n35 VSUBS 0.036249f
C1419 VTAIL.n36 VSUBS 0.036249f
C1420 VTAIL.n37 VSUBS 0.016238f
C1421 VTAIL.n38 VSUBS 0.015336f
C1422 VTAIL.n39 VSUBS 0.02854f
C1423 VTAIL.n40 VSUBS 0.02854f
C1424 VTAIL.n41 VSUBS 0.015336f
C1425 VTAIL.n42 VSUBS 0.016238f
C1426 VTAIL.n43 VSUBS 0.036249f
C1427 VTAIL.n44 VSUBS 0.036249f
C1428 VTAIL.n45 VSUBS 0.016238f
C1429 VTAIL.n46 VSUBS 0.015336f
C1430 VTAIL.n47 VSUBS 0.02854f
C1431 VTAIL.n48 VSUBS 0.02854f
C1432 VTAIL.n49 VSUBS 0.015336f
C1433 VTAIL.n50 VSUBS 0.016238f
C1434 VTAIL.n51 VSUBS 0.036249f
C1435 VTAIL.n52 VSUBS 0.036249f
C1436 VTAIL.n53 VSUBS 0.016238f
C1437 VTAIL.n54 VSUBS 0.015336f
C1438 VTAIL.n55 VSUBS 0.02854f
C1439 VTAIL.n56 VSUBS 0.02854f
C1440 VTAIL.n57 VSUBS 0.015336f
C1441 VTAIL.n58 VSUBS 0.016238f
C1442 VTAIL.n59 VSUBS 0.036249f
C1443 VTAIL.n60 VSUBS 0.036249f
C1444 VTAIL.n61 VSUBS 0.016238f
C1445 VTAIL.n62 VSUBS 0.015336f
C1446 VTAIL.n63 VSUBS 0.02854f
C1447 VTAIL.n64 VSUBS 0.02854f
C1448 VTAIL.n65 VSUBS 0.015336f
C1449 VTAIL.n66 VSUBS 0.016238f
C1450 VTAIL.n67 VSUBS 0.036249f
C1451 VTAIL.n68 VSUBS 0.036249f
C1452 VTAIL.n69 VSUBS 0.016238f
C1453 VTAIL.n70 VSUBS 0.015336f
C1454 VTAIL.n71 VSUBS 0.02854f
C1455 VTAIL.n72 VSUBS 0.02854f
C1456 VTAIL.n73 VSUBS 0.015336f
C1457 VTAIL.n74 VSUBS 0.015336f
C1458 VTAIL.n75 VSUBS 0.016238f
C1459 VTAIL.n76 VSUBS 0.036249f
C1460 VTAIL.n77 VSUBS 0.036249f
C1461 VTAIL.n78 VSUBS 0.036249f
C1462 VTAIL.n79 VSUBS 0.015787f
C1463 VTAIL.n80 VSUBS 0.015336f
C1464 VTAIL.n81 VSUBS 0.02854f
C1465 VTAIL.n82 VSUBS 0.02854f
C1466 VTAIL.n83 VSUBS 0.015336f
C1467 VTAIL.n84 VSUBS 0.016238f
C1468 VTAIL.n85 VSUBS 0.036249f
C1469 VTAIL.n86 VSUBS 0.086524f
C1470 VTAIL.n87 VSUBS 0.016238f
C1471 VTAIL.n88 VSUBS 0.015336f
C1472 VTAIL.n89 VSUBS 0.069867f
C1473 VTAIL.n90 VSUBS 0.043574f
C1474 VTAIL.n91 VSUBS 0.538314f
C1475 VTAIL.t7 VSUBS 0.364908f
C1476 VTAIL.t8 VSUBS 0.364908f
C1477 VTAIL.n92 VSUBS 2.83604f
C1478 VTAIL.n93 VSUBS 3.2774f
C1479 VTAIL.t5 VSUBS 0.364908f
C1480 VTAIL.t0 VSUBS 0.364908f
C1481 VTAIL.n94 VSUBS 2.83606f
C1482 VTAIL.n95 VSUBS 3.27738f
C1483 VTAIL.n96 VSUBS 0.030998f
C1484 VTAIL.n97 VSUBS 0.02854f
C1485 VTAIL.n98 VSUBS 0.015336f
C1486 VTAIL.n99 VSUBS 0.036249f
C1487 VTAIL.n100 VSUBS 0.016238f
C1488 VTAIL.n101 VSUBS 0.02854f
C1489 VTAIL.n102 VSUBS 0.015787f
C1490 VTAIL.n103 VSUBS 0.036249f
C1491 VTAIL.n104 VSUBS 0.015336f
C1492 VTAIL.n105 VSUBS 0.016238f
C1493 VTAIL.n106 VSUBS 0.02854f
C1494 VTAIL.n107 VSUBS 0.015336f
C1495 VTAIL.n108 VSUBS 0.036249f
C1496 VTAIL.n109 VSUBS 0.016238f
C1497 VTAIL.n110 VSUBS 0.02854f
C1498 VTAIL.n111 VSUBS 0.015336f
C1499 VTAIL.n112 VSUBS 0.036249f
C1500 VTAIL.n113 VSUBS 0.016238f
C1501 VTAIL.n114 VSUBS 0.02854f
C1502 VTAIL.n115 VSUBS 0.015336f
C1503 VTAIL.n116 VSUBS 0.036249f
C1504 VTAIL.n117 VSUBS 0.016238f
C1505 VTAIL.n118 VSUBS 0.02854f
C1506 VTAIL.n119 VSUBS 0.015336f
C1507 VTAIL.n120 VSUBS 0.036249f
C1508 VTAIL.n121 VSUBS 0.016238f
C1509 VTAIL.n122 VSUBS 0.02854f
C1510 VTAIL.n123 VSUBS 0.015336f
C1511 VTAIL.n124 VSUBS 0.027187f
C1512 VTAIL.n125 VSUBS 0.02306f
C1513 VTAIL.t2 VSUBS 0.077685f
C1514 VTAIL.n126 VSUBS 0.211114f
C1515 VTAIL.n127 VSUBS 1.97521f
C1516 VTAIL.n128 VSUBS 0.015336f
C1517 VTAIL.n129 VSUBS 0.016238f
C1518 VTAIL.n130 VSUBS 0.036249f
C1519 VTAIL.n131 VSUBS 0.036249f
C1520 VTAIL.n132 VSUBS 0.016238f
C1521 VTAIL.n133 VSUBS 0.015336f
C1522 VTAIL.n134 VSUBS 0.02854f
C1523 VTAIL.n135 VSUBS 0.02854f
C1524 VTAIL.n136 VSUBS 0.015336f
C1525 VTAIL.n137 VSUBS 0.016238f
C1526 VTAIL.n138 VSUBS 0.036249f
C1527 VTAIL.n139 VSUBS 0.036249f
C1528 VTAIL.n140 VSUBS 0.016238f
C1529 VTAIL.n141 VSUBS 0.015336f
C1530 VTAIL.n142 VSUBS 0.02854f
C1531 VTAIL.n143 VSUBS 0.02854f
C1532 VTAIL.n144 VSUBS 0.015336f
C1533 VTAIL.n145 VSUBS 0.016238f
C1534 VTAIL.n146 VSUBS 0.036249f
C1535 VTAIL.n147 VSUBS 0.036249f
C1536 VTAIL.n148 VSUBS 0.016238f
C1537 VTAIL.n149 VSUBS 0.015336f
C1538 VTAIL.n150 VSUBS 0.02854f
C1539 VTAIL.n151 VSUBS 0.02854f
C1540 VTAIL.n152 VSUBS 0.015336f
C1541 VTAIL.n153 VSUBS 0.016238f
C1542 VTAIL.n154 VSUBS 0.036249f
C1543 VTAIL.n155 VSUBS 0.036249f
C1544 VTAIL.n156 VSUBS 0.016238f
C1545 VTAIL.n157 VSUBS 0.015336f
C1546 VTAIL.n158 VSUBS 0.02854f
C1547 VTAIL.n159 VSUBS 0.02854f
C1548 VTAIL.n160 VSUBS 0.015336f
C1549 VTAIL.n161 VSUBS 0.016238f
C1550 VTAIL.n162 VSUBS 0.036249f
C1551 VTAIL.n163 VSUBS 0.036249f
C1552 VTAIL.n164 VSUBS 0.016238f
C1553 VTAIL.n165 VSUBS 0.015336f
C1554 VTAIL.n166 VSUBS 0.02854f
C1555 VTAIL.n167 VSUBS 0.02854f
C1556 VTAIL.n168 VSUBS 0.015336f
C1557 VTAIL.n169 VSUBS 0.016238f
C1558 VTAIL.n170 VSUBS 0.036249f
C1559 VTAIL.n171 VSUBS 0.036249f
C1560 VTAIL.n172 VSUBS 0.036249f
C1561 VTAIL.n173 VSUBS 0.015787f
C1562 VTAIL.n174 VSUBS 0.015336f
C1563 VTAIL.n175 VSUBS 0.02854f
C1564 VTAIL.n176 VSUBS 0.02854f
C1565 VTAIL.n177 VSUBS 0.015336f
C1566 VTAIL.n178 VSUBS 0.016238f
C1567 VTAIL.n179 VSUBS 0.036249f
C1568 VTAIL.n180 VSUBS 0.086524f
C1569 VTAIL.n181 VSUBS 0.016238f
C1570 VTAIL.n182 VSUBS 0.015336f
C1571 VTAIL.n183 VSUBS 0.069867f
C1572 VTAIL.n184 VSUBS 0.043574f
C1573 VTAIL.n185 VSUBS 0.538314f
C1574 VTAIL.t11 VSUBS 0.364908f
C1575 VTAIL.t6 VSUBS 0.364908f
C1576 VTAIL.n186 VSUBS 2.83606f
C1577 VTAIL.n187 VSUBS 1.18167f
C1578 VTAIL.n188 VSUBS 0.030998f
C1579 VTAIL.n189 VSUBS 0.02854f
C1580 VTAIL.n190 VSUBS 0.015336f
C1581 VTAIL.n191 VSUBS 0.036249f
C1582 VTAIL.n192 VSUBS 0.016238f
C1583 VTAIL.n193 VSUBS 0.02854f
C1584 VTAIL.n194 VSUBS 0.015787f
C1585 VTAIL.n195 VSUBS 0.036249f
C1586 VTAIL.n196 VSUBS 0.015336f
C1587 VTAIL.n197 VSUBS 0.016238f
C1588 VTAIL.n198 VSUBS 0.02854f
C1589 VTAIL.n199 VSUBS 0.015336f
C1590 VTAIL.n200 VSUBS 0.036249f
C1591 VTAIL.n201 VSUBS 0.016238f
C1592 VTAIL.n202 VSUBS 0.02854f
C1593 VTAIL.n203 VSUBS 0.015336f
C1594 VTAIL.n204 VSUBS 0.036249f
C1595 VTAIL.n205 VSUBS 0.016238f
C1596 VTAIL.n206 VSUBS 0.02854f
C1597 VTAIL.n207 VSUBS 0.015336f
C1598 VTAIL.n208 VSUBS 0.036249f
C1599 VTAIL.n209 VSUBS 0.016238f
C1600 VTAIL.n210 VSUBS 0.02854f
C1601 VTAIL.n211 VSUBS 0.015336f
C1602 VTAIL.n212 VSUBS 0.036249f
C1603 VTAIL.n213 VSUBS 0.016238f
C1604 VTAIL.n214 VSUBS 0.02854f
C1605 VTAIL.n215 VSUBS 0.015336f
C1606 VTAIL.n216 VSUBS 0.027187f
C1607 VTAIL.n217 VSUBS 0.02306f
C1608 VTAIL.t9 VSUBS 0.077685f
C1609 VTAIL.n218 VSUBS 0.211114f
C1610 VTAIL.n219 VSUBS 1.97521f
C1611 VTAIL.n220 VSUBS 0.015336f
C1612 VTAIL.n221 VSUBS 0.016238f
C1613 VTAIL.n222 VSUBS 0.036249f
C1614 VTAIL.n223 VSUBS 0.036249f
C1615 VTAIL.n224 VSUBS 0.016238f
C1616 VTAIL.n225 VSUBS 0.015336f
C1617 VTAIL.n226 VSUBS 0.02854f
C1618 VTAIL.n227 VSUBS 0.02854f
C1619 VTAIL.n228 VSUBS 0.015336f
C1620 VTAIL.n229 VSUBS 0.016238f
C1621 VTAIL.n230 VSUBS 0.036249f
C1622 VTAIL.n231 VSUBS 0.036249f
C1623 VTAIL.n232 VSUBS 0.016238f
C1624 VTAIL.n233 VSUBS 0.015336f
C1625 VTAIL.n234 VSUBS 0.02854f
C1626 VTAIL.n235 VSUBS 0.02854f
C1627 VTAIL.n236 VSUBS 0.015336f
C1628 VTAIL.n237 VSUBS 0.016238f
C1629 VTAIL.n238 VSUBS 0.036249f
C1630 VTAIL.n239 VSUBS 0.036249f
C1631 VTAIL.n240 VSUBS 0.016238f
C1632 VTAIL.n241 VSUBS 0.015336f
C1633 VTAIL.n242 VSUBS 0.02854f
C1634 VTAIL.n243 VSUBS 0.02854f
C1635 VTAIL.n244 VSUBS 0.015336f
C1636 VTAIL.n245 VSUBS 0.016238f
C1637 VTAIL.n246 VSUBS 0.036249f
C1638 VTAIL.n247 VSUBS 0.036249f
C1639 VTAIL.n248 VSUBS 0.016238f
C1640 VTAIL.n249 VSUBS 0.015336f
C1641 VTAIL.n250 VSUBS 0.02854f
C1642 VTAIL.n251 VSUBS 0.02854f
C1643 VTAIL.n252 VSUBS 0.015336f
C1644 VTAIL.n253 VSUBS 0.016238f
C1645 VTAIL.n254 VSUBS 0.036249f
C1646 VTAIL.n255 VSUBS 0.036249f
C1647 VTAIL.n256 VSUBS 0.016238f
C1648 VTAIL.n257 VSUBS 0.015336f
C1649 VTAIL.n258 VSUBS 0.02854f
C1650 VTAIL.n259 VSUBS 0.02854f
C1651 VTAIL.n260 VSUBS 0.015336f
C1652 VTAIL.n261 VSUBS 0.016238f
C1653 VTAIL.n262 VSUBS 0.036249f
C1654 VTAIL.n263 VSUBS 0.036249f
C1655 VTAIL.n264 VSUBS 0.036249f
C1656 VTAIL.n265 VSUBS 0.015787f
C1657 VTAIL.n266 VSUBS 0.015336f
C1658 VTAIL.n267 VSUBS 0.02854f
C1659 VTAIL.n268 VSUBS 0.02854f
C1660 VTAIL.n269 VSUBS 0.015336f
C1661 VTAIL.n270 VSUBS 0.016238f
C1662 VTAIL.n271 VSUBS 0.036249f
C1663 VTAIL.n272 VSUBS 0.086524f
C1664 VTAIL.n273 VSUBS 0.016238f
C1665 VTAIL.n274 VSUBS 0.015336f
C1666 VTAIL.n275 VSUBS 0.069867f
C1667 VTAIL.n276 VSUBS 0.043574f
C1668 VTAIL.n277 VSUBS 2.32167f
C1669 VTAIL.n278 VSUBS 0.030998f
C1670 VTAIL.n279 VSUBS 0.02854f
C1671 VTAIL.n280 VSUBS 0.015336f
C1672 VTAIL.n281 VSUBS 0.036249f
C1673 VTAIL.n282 VSUBS 0.016238f
C1674 VTAIL.n283 VSUBS 0.02854f
C1675 VTAIL.n284 VSUBS 0.015787f
C1676 VTAIL.n285 VSUBS 0.036249f
C1677 VTAIL.n286 VSUBS 0.016238f
C1678 VTAIL.n287 VSUBS 0.02854f
C1679 VTAIL.n288 VSUBS 0.015336f
C1680 VTAIL.n289 VSUBS 0.036249f
C1681 VTAIL.n290 VSUBS 0.016238f
C1682 VTAIL.n291 VSUBS 0.02854f
C1683 VTAIL.n292 VSUBS 0.015336f
C1684 VTAIL.n293 VSUBS 0.036249f
C1685 VTAIL.n294 VSUBS 0.016238f
C1686 VTAIL.n295 VSUBS 0.02854f
C1687 VTAIL.n296 VSUBS 0.015336f
C1688 VTAIL.n297 VSUBS 0.036249f
C1689 VTAIL.n298 VSUBS 0.016238f
C1690 VTAIL.n299 VSUBS 0.02854f
C1691 VTAIL.n300 VSUBS 0.015336f
C1692 VTAIL.n301 VSUBS 0.036249f
C1693 VTAIL.n302 VSUBS 0.016238f
C1694 VTAIL.n303 VSUBS 0.02854f
C1695 VTAIL.n304 VSUBS 0.015336f
C1696 VTAIL.n305 VSUBS 0.027187f
C1697 VTAIL.n306 VSUBS 0.02306f
C1698 VTAIL.t4 VSUBS 0.077685f
C1699 VTAIL.n307 VSUBS 0.211114f
C1700 VTAIL.n308 VSUBS 1.97521f
C1701 VTAIL.n309 VSUBS 0.015336f
C1702 VTAIL.n310 VSUBS 0.016238f
C1703 VTAIL.n311 VSUBS 0.036249f
C1704 VTAIL.n312 VSUBS 0.036249f
C1705 VTAIL.n313 VSUBS 0.016238f
C1706 VTAIL.n314 VSUBS 0.015336f
C1707 VTAIL.n315 VSUBS 0.02854f
C1708 VTAIL.n316 VSUBS 0.02854f
C1709 VTAIL.n317 VSUBS 0.015336f
C1710 VTAIL.n318 VSUBS 0.016238f
C1711 VTAIL.n319 VSUBS 0.036249f
C1712 VTAIL.n320 VSUBS 0.036249f
C1713 VTAIL.n321 VSUBS 0.016238f
C1714 VTAIL.n322 VSUBS 0.015336f
C1715 VTAIL.n323 VSUBS 0.02854f
C1716 VTAIL.n324 VSUBS 0.02854f
C1717 VTAIL.n325 VSUBS 0.015336f
C1718 VTAIL.n326 VSUBS 0.016238f
C1719 VTAIL.n327 VSUBS 0.036249f
C1720 VTAIL.n328 VSUBS 0.036249f
C1721 VTAIL.n329 VSUBS 0.016238f
C1722 VTAIL.n330 VSUBS 0.015336f
C1723 VTAIL.n331 VSUBS 0.02854f
C1724 VTAIL.n332 VSUBS 0.02854f
C1725 VTAIL.n333 VSUBS 0.015336f
C1726 VTAIL.n334 VSUBS 0.016238f
C1727 VTAIL.n335 VSUBS 0.036249f
C1728 VTAIL.n336 VSUBS 0.036249f
C1729 VTAIL.n337 VSUBS 0.016238f
C1730 VTAIL.n338 VSUBS 0.015336f
C1731 VTAIL.n339 VSUBS 0.02854f
C1732 VTAIL.n340 VSUBS 0.02854f
C1733 VTAIL.n341 VSUBS 0.015336f
C1734 VTAIL.n342 VSUBS 0.016238f
C1735 VTAIL.n343 VSUBS 0.036249f
C1736 VTAIL.n344 VSUBS 0.036249f
C1737 VTAIL.n345 VSUBS 0.016238f
C1738 VTAIL.n346 VSUBS 0.015336f
C1739 VTAIL.n347 VSUBS 0.02854f
C1740 VTAIL.n348 VSUBS 0.02854f
C1741 VTAIL.n349 VSUBS 0.015336f
C1742 VTAIL.n350 VSUBS 0.015336f
C1743 VTAIL.n351 VSUBS 0.016238f
C1744 VTAIL.n352 VSUBS 0.036249f
C1745 VTAIL.n353 VSUBS 0.036249f
C1746 VTAIL.n354 VSUBS 0.036249f
C1747 VTAIL.n355 VSUBS 0.015787f
C1748 VTAIL.n356 VSUBS 0.015336f
C1749 VTAIL.n357 VSUBS 0.02854f
C1750 VTAIL.n358 VSUBS 0.02854f
C1751 VTAIL.n359 VSUBS 0.015336f
C1752 VTAIL.n360 VSUBS 0.016238f
C1753 VTAIL.n361 VSUBS 0.036249f
C1754 VTAIL.n362 VSUBS 0.086524f
C1755 VTAIL.n363 VSUBS 0.016238f
C1756 VTAIL.n364 VSUBS 0.015336f
C1757 VTAIL.n365 VSUBS 0.069867f
C1758 VTAIL.n366 VSUBS 0.043574f
C1759 VTAIL.n367 VSUBS 2.23823f
C1760 VP.t1 VSUBS 4.06737f
C1761 VP.n0 VSUBS 1.50652f
C1762 VP.n1 VSUBS 0.02537f
C1763 VP.n2 VSUBS 0.038986f
C1764 VP.n3 VSUBS 0.02537f
C1765 VP.n4 VSUBS 0.035434f
C1766 VP.n5 VSUBS 0.02537f
C1767 VP.n6 VSUBS 0.034774f
C1768 VP.n7 VSUBS 0.02537f
C1769 VP.n8 VSUBS 0.032647f
C1770 VP.t5 VSUBS 4.06737f
C1771 VP.n9 VSUBS 1.50652f
C1772 VP.n10 VSUBS 0.02537f
C1773 VP.n11 VSUBS 0.038986f
C1774 VP.n12 VSUBS 0.02537f
C1775 VP.n13 VSUBS 0.035434f
C1776 VP.t0 VSUBS 4.44485f
C1777 VP.t2 VSUBS 4.06737f
C1778 VP.n14 VSUBS 1.49518f
C1779 VP.n15 VSUBS 1.4227f
C1780 VP.n16 VSUBS 0.316923f
C1781 VP.n17 VSUBS 0.02537f
C1782 VP.n18 VSUBS 0.047047f
C1783 VP.n19 VSUBS 0.047047f
C1784 VP.n20 VSUBS 0.034774f
C1785 VP.n21 VSUBS 0.02537f
C1786 VP.n22 VSUBS 0.02537f
C1787 VP.n23 VSUBS 0.02537f
C1788 VP.n24 VSUBS 0.047047f
C1789 VP.n25 VSUBS 0.047047f
C1790 VP.n26 VSUBS 0.032647f
C1791 VP.n27 VSUBS 0.040941f
C1792 VP.n28 VSUBS 1.69771f
C1793 VP.t4 VSUBS 4.06737f
C1794 VP.n29 VSUBS 1.50652f
C1795 VP.n30 VSUBS 1.71407f
C1796 VP.n31 VSUBS 0.040941f
C1797 VP.n32 VSUBS 0.02537f
C1798 VP.n33 VSUBS 0.047047f
C1799 VP.n34 VSUBS 0.047047f
C1800 VP.n35 VSUBS 0.038986f
C1801 VP.n36 VSUBS 0.02537f
C1802 VP.n37 VSUBS 0.02537f
C1803 VP.n38 VSUBS 0.02537f
C1804 VP.n39 VSUBS 0.047047f
C1805 VP.n40 VSUBS 0.047047f
C1806 VP.t3 VSUBS 4.06737f
C1807 VP.n41 VSUBS 1.40753f
C1808 VP.n42 VSUBS 0.035434f
C1809 VP.n43 VSUBS 0.02537f
C1810 VP.n44 VSUBS 0.02537f
C1811 VP.n45 VSUBS 0.02537f
C1812 VP.n46 VSUBS 0.047047f
C1813 VP.n47 VSUBS 0.047047f
C1814 VP.n48 VSUBS 0.034774f
C1815 VP.n49 VSUBS 0.02537f
C1816 VP.n50 VSUBS 0.02537f
C1817 VP.n51 VSUBS 0.02537f
C1818 VP.n52 VSUBS 0.047047f
C1819 VP.n53 VSUBS 0.047047f
C1820 VP.n54 VSUBS 0.032647f
C1821 VP.n55 VSUBS 0.040941f
C1822 VP.n56 VSUBS 0.070028f
.ends

