* NGSPICE file created from diff_pair_sample_1135.ext - technology: sky130A

.subckt diff_pair_sample_1135 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=6.5325 pd=34.28 as=0 ps=0 w=16.75 l=1.31
X1 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=6.5325 pd=34.28 as=0 ps=0 w=16.75 l=1.31
X2 VDD1.t1 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=6.5325 pd=34.28 as=6.5325 ps=34.28 w=16.75 l=1.31
X3 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=6.5325 pd=34.28 as=0 ps=0 w=16.75 l=1.31
X4 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.5325 pd=34.28 as=0 ps=0 w=16.75 l=1.31
X5 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.5325 pd=34.28 as=6.5325 ps=34.28 w=16.75 l=1.31
X6 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.5325 pd=34.28 as=6.5325 ps=34.28 w=16.75 l=1.31
X7 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=6.5325 pd=34.28 as=6.5325 ps=34.28 w=16.75 l=1.31
R0 B.n758 B.n757 585
R1 B.n759 B.n758 585
R2 B.n340 B.n95 585
R3 B.n339 B.n338 585
R4 B.n337 B.n336 585
R5 B.n335 B.n334 585
R6 B.n333 B.n332 585
R7 B.n331 B.n330 585
R8 B.n329 B.n328 585
R9 B.n327 B.n326 585
R10 B.n325 B.n324 585
R11 B.n323 B.n322 585
R12 B.n321 B.n320 585
R13 B.n319 B.n318 585
R14 B.n317 B.n316 585
R15 B.n315 B.n314 585
R16 B.n313 B.n312 585
R17 B.n311 B.n310 585
R18 B.n309 B.n308 585
R19 B.n307 B.n306 585
R20 B.n305 B.n304 585
R21 B.n303 B.n302 585
R22 B.n301 B.n300 585
R23 B.n299 B.n298 585
R24 B.n297 B.n296 585
R25 B.n295 B.n294 585
R26 B.n293 B.n292 585
R27 B.n291 B.n290 585
R28 B.n289 B.n288 585
R29 B.n287 B.n286 585
R30 B.n285 B.n284 585
R31 B.n283 B.n282 585
R32 B.n281 B.n280 585
R33 B.n279 B.n278 585
R34 B.n277 B.n276 585
R35 B.n275 B.n274 585
R36 B.n273 B.n272 585
R37 B.n271 B.n270 585
R38 B.n269 B.n268 585
R39 B.n267 B.n266 585
R40 B.n265 B.n264 585
R41 B.n263 B.n262 585
R42 B.n261 B.n260 585
R43 B.n259 B.n258 585
R44 B.n257 B.n256 585
R45 B.n255 B.n254 585
R46 B.n253 B.n252 585
R47 B.n251 B.n250 585
R48 B.n249 B.n248 585
R49 B.n247 B.n246 585
R50 B.n245 B.n244 585
R51 B.n243 B.n242 585
R52 B.n241 B.n240 585
R53 B.n239 B.n238 585
R54 B.n237 B.n236 585
R55 B.n235 B.n234 585
R56 B.n233 B.n232 585
R57 B.n230 B.n229 585
R58 B.n228 B.n227 585
R59 B.n226 B.n225 585
R60 B.n224 B.n223 585
R61 B.n222 B.n221 585
R62 B.n220 B.n219 585
R63 B.n218 B.n217 585
R64 B.n216 B.n215 585
R65 B.n214 B.n213 585
R66 B.n212 B.n211 585
R67 B.n210 B.n209 585
R68 B.n208 B.n207 585
R69 B.n206 B.n205 585
R70 B.n204 B.n203 585
R71 B.n202 B.n201 585
R72 B.n200 B.n199 585
R73 B.n198 B.n197 585
R74 B.n196 B.n195 585
R75 B.n194 B.n193 585
R76 B.n192 B.n191 585
R77 B.n190 B.n189 585
R78 B.n188 B.n187 585
R79 B.n186 B.n185 585
R80 B.n184 B.n183 585
R81 B.n182 B.n181 585
R82 B.n180 B.n179 585
R83 B.n178 B.n177 585
R84 B.n176 B.n175 585
R85 B.n174 B.n173 585
R86 B.n172 B.n171 585
R87 B.n170 B.n169 585
R88 B.n168 B.n167 585
R89 B.n166 B.n165 585
R90 B.n164 B.n163 585
R91 B.n162 B.n161 585
R92 B.n160 B.n159 585
R93 B.n158 B.n157 585
R94 B.n156 B.n155 585
R95 B.n154 B.n153 585
R96 B.n152 B.n151 585
R97 B.n150 B.n149 585
R98 B.n148 B.n147 585
R99 B.n146 B.n145 585
R100 B.n144 B.n143 585
R101 B.n142 B.n141 585
R102 B.n140 B.n139 585
R103 B.n138 B.n137 585
R104 B.n136 B.n135 585
R105 B.n134 B.n133 585
R106 B.n132 B.n131 585
R107 B.n130 B.n129 585
R108 B.n128 B.n127 585
R109 B.n126 B.n125 585
R110 B.n124 B.n123 585
R111 B.n122 B.n121 585
R112 B.n120 B.n119 585
R113 B.n118 B.n117 585
R114 B.n116 B.n115 585
R115 B.n114 B.n113 585
R116 B.n112 B.n111 585
R117 B.n110 B.n109 585
R118 B.n108 B.n107 585
R119 B.n106 B.n105 585
R120 B.n104 B.n103 585
R121 B.n102 B.n101 585
R122 B.n756 B.n34 585
R123 B.n760 B.n34 585
R124 B.n755 B.n33 585
R125 B.n761 B.n33 585
R126 B.n754 B.n753 585
R127 B.n753 B.n29 585
R128 B.n752 B.n28 585
R129 B.n767 B.n28 585
R130 B.n751 B.n27 585
R131 B.n768 B.n27 585
R132 B.n750 B.n26 585
R133 B.n769 B.n26 585
R134 B.n749 B.n748 585
R135 B.n748 B.n22 585
R136 B.n747 B.n21 585
R137 B.n775 B.n21 585
R138 B.n746 B.n20 585
R139 B.n776 B.n20 585
R140 B.n745 B.n19 585
R141 B.n777 B.n19 585
R142 B.n744 B.n743 585
R143 B.n743 B.n15 585
R144 B.n742 B.n14 585
R145 B.n783 B.n14 585
R146 B.n741 B.n13 585
R147 B.n784 B.n13 585
R148 B.n740 B.n12 585
R149 B.n785 B.n12 585
R150 B.n739 B.n738 585
R151 B.n738 B.n737 585
R152 B.n736 B.n735 585
R153 B.n736 B.n8 585
R154 B.n734 B.n7 585
R155 B.n792 B.n7 585
R156 B.n733 B.n6 585
R157 B.n793 B.n6 585
R158 B.n732 B.n5 585
R159 B.n794 B.n5 585
R160 B.n731 B.n730 585
R161 B.n730 B.n4 585
R162 B.n729 B.n341 585
R163 B.n729 B.n728 585
R164 B.n719 B.n342 585
R165 B.n343 B.n342 585
R166 B.n721 B.n720 585
R167 B.n722 B.n721 585
R168 B.n718 B.n348 585
R169 B.n348 B.n347 585
R170 B.n717 B.n716 585
R171 B.n716 B.n715 585
R172 B.n350 B.n349 585
R173 B.n351 B.n350 585
R174 B.n708 B.n707 585
R175 B.n709 B.n708 585
R176 B.n706 B.n356 585
R177 B.n356 B.n355 585
R178 B.n705 B.n704 585
R179 B.n704 B.n703 585
R180 B.n358 B.n357 585
R181 B.n359 B.n358 585
R182 B.n696 B.n695 585
R183 B.n697 B.n696 585
R184 B.n694 B.n364 585
R185 B.n364 B.n363 585
R186 B.n693 B.n692 585
R187 B.n692 B.n691 585
R188 B.n366 B.n365 585
R189 B.n367 B.n366 585
R190 B.n684 B.n683 585
R191 B.n685 B.n684 585
R192 B.n682 B.n372 585
R193 B.n372 B.n371 585
R194 B.n676 B.n675 585
R195 B.n674 B.n434 585
R196 B.n673 B.n433 585
R197 B.n678 B.n433 585
R198 B.n672 B.n671 585
R199 B.n670 B.n669 585
R200 B.n668 B.n667 585
R201 B.n666 B.n665 585
R202 B.n664 B.n663 585
R203 B.n662 B.n661 585
R204 B.n660 B.n659 585
R205 B.n658 B.n657 585
R206 B.n656 B.n655 585
R207 B.n654 B.n653 585
R208 B.n652 B.n651 585
R209 B.n650 B.n649 585
R210 B.n648 B.n647 585
R211 B.n646 B.n645 585
R212 B.n644 B.n643 585
R213 B.n642 B.n641 585
R214 B.n640 B.n639 585
R215 B.n638 B.n637 585
R216 B.n636 B.n635 585
R217 B.n634 B.n633 585
R218 B.n632 B.n631 585
R219 B.n630 B.n629 585
R220 B.n628 B.n627 585
R221 B.n626 B.n625 585
R222 B.n624 B.n623 585
R223 B.n622 B.n621 585
R224 B.n620 B.n619 585
R225 B.n618 B.n617 585
R226 B.n616 B.n615 585
R227 B.n614 B.n613 585
R228 B.n612 B.n611 585
R229 B.n610 B.n609 585
R230 B.n608 B.n607 585
R231 B.n606 B.n605 585
R232 B.n604 B.n603 585
R233 B.n602 B.n601 585
R234 B.n600 B.n599 585
R235 B.n598 B.n597 585
R236 B.n596 B.n595 585
R237 B.n594 B.n593 585
R238 B.n592 B.n591 585
R239 B.n590 B.n589 585
R240 B.n588 B.n587 585
R241 B.n586 B.n585 585
R242 B.n584 B.n583 585
R243 B.n582 B.n581 585
R244 B.n580 B.n579 585
R245 B.n578 B.n577 585
R246 B.n576 B.n575 585
R247 B.n574 B.n573 585
R248 B.n572 B.n571 585
R249 B.n570 B.n569 585
R250 B.n568 B.n567 585
R251 B.n565 B.n564 585
R252 B.n563 B.n562 585
R253 B.n561 B.n560 585
R254 B.n559 B.n558 585
R255 B.n557 B.n556 585
R256 B.n555 B.n554 585
R257 B.n553 B.n552 585
R258 B.n551 B.n550 585
R259 B.n549 B.n548 585
R260 B.n547 B.n546 585
R261 B.n545 B.n544 585
R262 B.n543 B.n542 585
R263 B.n541 B.n540 585
R264 B.n539 B.n538 585
R265 B.n537 B.n536 585
R266 B.n535 B.n534 585
R267 B.n533 B.n532 585
R268 B.n531 B.n530 585
R269 B.n529 B.n528 585
R270 B.n527 B.n526 585
R271 B.n525 B.n524 585
R272 B.n523 B.n522 585
R273 B.n521 B.n520 585
R274 B.n519 B.n518 585
R275 B.n517 B.n516 585
R276 B.n515 B.n514 585
R277 B.n513 B.n512 585
R278 B.n511 B.n510 585
R279 B.n509 B.n508 585
R280 B.n507 B.n506 585
R281 B.n505 B.n504 585
R282 B.n503 B.n502 585
R283 B.n501 B.n500 585
R284 B.n499 B.n498 585
R285 B.n497 B.n496 585
R286 B.n495 B.n494 585
R287 B.n493 B.n492 585
R288 B.n491 B.n490 585
R289 B.n489 B.n488 585
R290 B.n487 B.n486 585
R291 B.n485 B.n484 585
R292 B.n483 B.n482 585
R293 B.n481 B.n480 585
R294 B.n479 B.n478 585
R295 B.n477 B.n476 585
R296 B.n475 B.n474 585
R297 B.n473 B.n472 585
R298 B.n471 B.n470 585
R299 B.n469 B.n468 585
R300 B.n467 B.n466 585
R301 B.n465 B.n464 585
R302 B.n463 B.n462 585
R303 B.n461 B.n460 585
R304 B.n459 B.n458 585
R305 B.n457 B.n456 585
R306 B.n455 B.n454 585
R307 B.n453 B.n452 585
R308 B.n451 B.n450 585
R309 B.n449 B.n448 585
R310 B.n447 B.n446 585
R311 B.n445 B.n444 585
R312 B.n443 B.n442 585
R313 B.n441 B.n440 585
R314 B.n374 B.n373 585
R315 B.n681 B.n680 585
R316 B.n370 B.n369 585
R317 B.n371 B.n370 585
R318 B.n687 B.n686 585
R319 B.n686 B.n685 585
R320 B.n688 B.n368 585
R321 B.n368 B.n367 585
R322 B.n690 B.n689 585
R323 B.n691 B.n690 585
R324 B.n362 B.n361 585
R325 B.n363 B.n362 585
R326 B.n699 B.n698 585
R327 B.n698 B.n697 585
R328 B.n700 B.n360 585
R329 B.n360 B.n359 585
R330 B.n702 B.n701 585
R331 B.n703 B.n702 585
R332 B.n354 B.n353 585
R333 B.n355 B.n354 585
R334 B.n711 B.n710 585
R335 B.n710 B.n709 585
R336 B.n712 B.n352 585
R337 B.n352 B.n351 585
R338 B.n714 B.n713 585
R339 B.n715 B.n714 585
R340 B.n346 B.n345 585
R341 B.n347 B.n346 585
R342 B.n724 B.n723 585
R343 B.n723 B.n722 585
R344 B.n725 B.n344 585
R345 B.n344 B.n343 585
R346 B.n727 B.n726 585
R347 B.n728 B.n727 585
R348 B.n3 B.n0 585
R349 B.n4 B.n3 585
R350 B.n791 B.n1 585
R351 B.n792 B.n791 585
R352 B.n790 B.n789 585
R353 B.n790 B.n8 585
R354 B.n788 B.n9 585
R355 B.n737 B.n9 585
R356 B.n787 B.n786 585
R357 B.n786 B.n785 585
R358 B.n11 B.n10 585
R359 B.n784 B.n11 585
R360 B.n782 B.n781 585
R361 B.n783 B.n782 585
R362 B.n780 B.n16 585
R363 B.n16 B.n15 585
R364 B.n779 B.n778 585
R365 B.n778 B.n777 585
R366 B.n18 B.n17 585
R367 B.n776 B.n18 585
R368 B.n774 B.n773 585
R369 B.n775 B.n774 585
R370 B.n772 B.n23 585
R371 B.n23 B.n22 585
R372 B.n771 B.n770 585
R373 B.n770 B.n769 585
R374 B.n25 B.n24 585
R375 B.n768 B.n25 585
R376 B.n766 B.n765 585
R377 B.n767 B.n766 585
R378 B.n764 B.n30 585
R379 B.n30 B.n29 585
R380 B.n763 B.n762 585
R381 B.n762 B.n761 585
R382 B.n32 B.n31 585
R383 B.n760 B.n32 585
R384 B.n795 B.n794 585
R385 B.n793 B.n2 585
R386 B.n101 B.n32 521.33
R387 B.n758 B.n34 521.33
R388 B.n680 B.n372 521.33
R389 B.n676 B.n370 521.33
R390 B.n98 B.t6 512.804
R391 B.n96 B.t2 512.804
R392 B.n437 B.t13 512.804
R393 B.n435 B.t9 512.804
R394 B.n96 B.t4 395.608
R395 B.n437 B.t15 395.608
R396 B.n98 B.t7 395.608
R397 B.n435 B.t12 395.608
R398 B.n97 B.t5 363.801
R399 B.n438 B.t14 363.801
R400 B.n99 B.t8 363.801
R401 B.n436 B.t11 363.801
R402 B.n759 B.n94 256.663
R403 B.n759 B.n93 256.663
R404 B.n759 B.n92 256.663
R405 B.n759 B.n91 256.663
R406 B.n759 B.n90 256.663
R407 B.n759 B.n89 256.663
R408 B.n759 B.n88 256.663
R409 B.n759 B.n87 256.663
R410 B.n759 B.n86 256.663
R411 B.n759 B.n85 256.663
R412 B.n759 B.n84 256.663
R413 B.n759 B.n83 256.663
R414 B.n759 B.n82 256.663
R415 B.n759 B.n81 256.663
R416 B.n759 B.n80 256.663
R417 B.n759 B.n79 256.663
R418 B.n759 B.n78 256.663
R419 B.n759 B.n77 256.663
R420 B.n759 B.n76 256.663
R421 B.n759 B.n75 256.663
R422 B.n759 B.n74 256.663
R423 B.n759 B.n73 256.663
R424 B.n759 B.n72 256.663
R425 B.n759 B.n71 256.663
R426 B.n759 B.n70 256.663
R427 B.n759 B.n69 256.663
R428 B.n759 B.n68 256.663
R429 B.n759 B.n67 256.663
R430 B.n759 B.n66 256.663
R431 B.n759 B.n65 256.663
R432 B.n759 B.n64 256.663
R433 B.n759 B.n63 256.663
R434 B.n759 B.n62 256.663
R435 B.n759 B.n61 256.663
R436 B.n759 B.n60 256.663
R437 B.n759 B.n59 256.663
R438 B.n759 B.n58 256.663
R439 B.n759 B.n57 256.663
R440 B.n759 B.n56 256.663
R441 B.n759 B.n55 256.663
R442 B.n759 B.n54 256.663
R443 B.n759 B.n53 256.663
R444 B.n759 B.n52 256.663
R445 B.n759 B.n51 256.663
R446 B.n759 B.n50 256.663
R447 B.n759 B.n49 256.663
R448 B.n759 B.n48 256.663
R449 B.n759 B.n47 256.663
R450 B.n759 B.n46 256.663
R451 B.n759 B.n45 256.663
R452 B.n759 B.n44 256.663
R453 B.n759 B.n43 256.663
R454 B.n759 B.n42 256.663
R455 B.n759 B.n41 256.663
R456 B.n759 B.n40 256.663
R457 B.n759 B.n39 256.663
R458 B.n759 B.n38 256.663
R459 B.n759 B.n37 256.663
R460 B.n759 B.n36 256.663
R461 B.n759 B.n35 256.663
R462 B.n678 B.n677 256.663
R463 B.n678 B.n375 256.663
R464 B.n678 B.n376 256.663
R465 B.n678 B.n377 256.663
R466 B.n678 B.n378 256.663
R467 B.n678 B.n379 256.663
R468 B.n678 B.n380 256.663
R469 B.n678 B.n381 256.663
R470 B.n678 B.n382 256.663
R471 B.n678 B.n383 256.663
R472 B.n678 B.n384 256.663
R473 B.n678 B.n385 256.663
R474 B.n678 B.n386 256.663
R475 B.n678 B.n387 256.663
R476 B.n678 B.n388 256.663
R477 B.n678 B.n389 256.663
R478 B.n678 B.n390 256.663
R479 B.n678 B.n391 256.663
R480 B.n678 B.n392 256.663
R481 B.n678 B.n393 256.663
R482 B.n678 B.n394 256.663
R483 B.n678 B.n395 256.663
R484 B.n678 B.n396 256.663
R485 B.n678 B.n397 256.663
R486 B.n678 B.n398 256.663
R487 B.n678 B.n399 256.663
R488 B.n678 B.n400 256.663
R489 B.n678 B.n401 256.663
R490 B.n678 B.n402 256.663
R491 B.n678 B.n403 256.663
R492 B.n678 B.n404 256.663
R493 B.n678 B.n405 256.663
R494 B.n678 B.n406 256.663
R495 B.n678 B.n407 256.663
R496 B.n678 B.n408 256.663
R497 B.n678 B.n409 256.663
R498 B.n678 B.n410 256.663
R499 B.n678 B.n411 256.663
R500 B.n678 B.n412 256.663
R501 B.n678 B.n413 256.663
R502 B.n678 B.n414 256.663
R503 B.n678 B.n415 256.663
R504 B.n678 B.n416 256.663
R505 B.n678 B.n417 256.663
R506 B.n678 B.n418 256.663
R507 B.n678 B.n419 256.663
R508 B.n678 B.n420 256.663
R509 B.n678 B.n421 256.663
R510 B.n678 B.n422 256.663
R511 B.n678 B.n423 256.663
R512 B.n678 B.n424 256.663
R513 B.n678 B.n425 256.663
R514 B.n678 B.n426 256.663
R515 B.n678 B.n427 256.663
R516 B.n678 B.n428 256.663
R517 B.n678 B.n429 256.663
R518 B.n678 B.n430 256.663
R519 B.n678 B.n431 256.663
R520 B.n678 B.n432 256.663
R521 B.n679 B.n678 256.663
R522 B.n797 B.n796 256.663
R523 B.n105 B.n104 163.367
R524 B.n109 B.n108 163.367
R525 B.n113 B.n112 163.367
R526 B.n117 B.n116 163.367
R527 B.n121 B.n120 163.367
R528 B.n125 B.n124 163.367
R529 B.n129 B.n128 163.367
R530 B.n133 B.n132 163.367
R531 B.n137 B.n136 163.367
R532 B.n141 B.n140 163.367
R533 B.n145 B.n144 163.367
R534 B.n149 B.n148 163.367
R535 B.n153 B.n152 163.367
R536 B.n157 B.n156 163.367
R537 B.n161 B.n160 163.367
R538 B.n165 B.n164 163.367
R539 B.n169 B.n168 163.367
R540 B.n173 B.n172 163.367
R541 B.n177 B.n176 163.367
R542 B.n181 B.n180 163.367
R543 B.n185 B.n184 163.367
R544 B.n189 B.n188 163.367
R545 B.n193 B.n192 163.367
R546 B.n197 B.n196 163.367
R547 B.n201 B.n200 163.367
R548 B.n205 B.n204 163.367
R549 B.n209 B.n208 163.367
R550 B.n213 B.n212 163.367
R551 B.n217 B.n216 163.367
R552 B.n221 B.n220 163.367
R553 B.n225 B.n224 163.367
R554 B.n229 B.n228 163.367
R555 B.n234 B.n233 163.367
R556 B.n238 B.n237 163.367
R557 B.n242 B.n241 163.367
R558 B.n246 B.n245 163.367
R559 B.n250 B.n249 163.367
R560 B.n254 B.n253 163.367
R561 B.n258 B.n257 163.367
R562 B.n262 B.n261 163.367
R563 B.n266 B.n265 163.367
R564 B.n270 B.n269 163.367
R565 B.n274 B.n273 163.367
R566 B.n278 B.n277 163.367
R567 B.n282 B.n281 163.367
R568 B.n286 B.n285 163.367
R569 B.n290 B.n289 163.367
R570 B.n294 B.n293 163.367
R571 B.n298 B.n297 163.367
R572 B.n302 B.n301 163.367
R573 B.n306 B.n305 163.367
R574 B.n310 B.n309 163.367
R575 B.n314 B.n313 163.367
R576 B.n318 B.n317 163.367
R577 B.n322 B.n321 163.367
R578 B.n326 B.n325 163.367
R579 B.n330 B.n329 163.367
R580 B.n334 B.n333 163.367
R581 B.n338 B.n337 163.367
R582 B.n758 B.n95 163.367
R583 B.n684 B.n372 163.367
R584 B.n684 B.n366 163.367
R585 B.n692 B.n366 163.367
R586 B.n692 B.n364 163.367
R587 B.n696 B.n364 163.367
R588 B.n696 B.n358 163.367
R589 B.n704 B.n358 163.367
R590 B.n704 B.n356 163.367
R591 B.n708 B.n356 163.367
R592 B.n708 B.n350 163.367
R593 B.n716 B.n350 163.367
R594 B.n716 B.n348 163.367
R595 B.n721 B.n348 163.367
R596 B.n721 B.n342 163.367
R597 B.n729 B.n342 163.367
R598 B.n730 B.n729 163.367
R599 B.n730 B.n5 163.367
R600 B.n6 B.n5 163.367
R601 B.n7 B.n6 163.367
R602 B.n736 B.n7 163.367
R603 B.n738 B.n736 163.367
R604 B.n738 B.n12 163.367
R605 B.n13 B.n12 163.367
R606 B.n14 B.n13 163.367
R607 B.n743 B.n14 163.367
R608 B.n743 B.n19 163.367
R609 B.n20 B.n19 163.367
R610 B.n21 B.n20 163.367
R611 B.n748 B.n21 163.367
R612 B.n748 B.n26 163.367
R613 B.n27 B.n26 163.367
R614 B.n28 B.n27 163.367
R615 B.n753 B.n28 163.367
R616 B.n753 B.n33 163.367
R617 B.n34 B.n33 163.367
R618 B.n434 B.n433 163.367
R619 B.n671 B.n433 163.367
R620 B.n669 B.n668 163.367
R621 B.n665 B.n664 163.367
R622 B.n661 B.n660 163.367
R623 B.n657 B.n656 163.367
R624 B.n653 B.n652 163.367
R625 B.n649 B.n648 163.367
R626 B.n645 B.n644 163.367
R627 B.n641 B.n640 163.367
R628 B.n637 B.n636 163.367
R629 B.n633 B.n632 163.367
R630 B.n629 B.n628 163.367
R631 B.n625 B.n624 163.367
R632 B.n621 B.n620 163.367
R633 B.n617 B.n616 163.367
R634 B.n613 B.n612 163.367
R635 B.n609 B.n608 163.367
R636 B.n605 B.n604 163.367
R637 B.n601 B.n600 163.367
R638 B.n597 B.n596 163.367
R639 B.n593 B.n592 163.367
R640 B.n589 B.n588 163.367
R641 B.n585 B.n584 163.367
R642 B.n581 B.n580 163.367
R643 B.n577 B.n576 163.367
R644 B.n573 B.n572 163.367
R645 B.n569 B.n568 163.367
R646 B.n564 B.n563 163.367
R647 B.n560 B.n559 163.367
R648 B.n556 B.n555 163.367
R649 B.n552 B.n551 163.367
R650 B.n548 B.n547 163.367
R651 B.n544 B.n543 163.367
R652 B.n540 B.n539 163.367
R653 B.n536 B.n535 163.367
R654 B.n532 B.n531 163.367
R655 B.n528 B.n527 163.367
R656 B.n524 B.n523 163.367
R657 B.n520 B.n519 163.367
R658 B.n516 B.n515 163.367
R659 B.n512 B.n511 163.367
R660 B.n508 B.n507 163.367
R661 B.n504 B.n503 163.367
R662 B.n500 B.n499 163.367
R663 B.n496 B.n495 163.367
R664 B.n492 B.n491 163.367
R665 B.n488 B.n487 163.367
R666 B.n484 B.n483 163.367
R667 B.n480 B.n479 163.367
R668 B.n476 B.n475 163.367
R669 B.n472 B.n471 163.367
R670 B.n468 B.n467 163.367
R671 B.n464 B.n463 163.367
R672 B.n460 B.n459 163.367
R673 B.n456 B.n455 163.367
R674 B.n452 B.n451 163.367
R675 B.n448 B.n447 163.367
R676 B.n444 B.n443 163.367
R677 B.n440 B.n374 163.367
R678 B.n686 B.n370 163.367
R679 B.n686 B.n368 163.367
R680 B.n690 B.n368 163.367
R681 B.n690 B.n362 163.367
R682 B.n698 B.n362 163.367
R683 B.n698 B.n360 163.367
R684 B.n702 B.n360 163.367
R685 B.n702 B.n354 163.367
R686 B.n710 B.n354 163.367
R687 B.n710 B.n352 163.367
R688 B.n714 B.n352 163.367
R689 B.n714 B.n346 163.367
R690 B.n723 B.n346 163.367
R691 B.n723 B.n344 163.367
R692 B.n727 B.n344 163.367
R693 B.n727 B.n3 163.367
R694 B.n795 B.n3 163.367
R695 B.n791 B.n2 163.367
R696 B.n791 B.n790 163.367
R697 B.n790 B.n9 163.367
R698 B.n786 B.n9 163.367
R699 B.n786 B.n11 163.367
R700 B.n782 B.n11 163.367
R701 B.n782 B.n16 163.367
R702 B.n778 B.n16 163.367
R703 B.n778 B.n18 163.367
R704 B.n774 B.n18 163.367
R705 B.n774 B.n23 163.367
R706 B.n770 B.n23 163.367
R707 B.n770 B.n25 163.367
R708 B.n766 B.n25 163.367
R709 B.n766 B.n30 163.367
R710 B.n762 B.n30 163.367
R711 B.n762 B.n32 163.367
R712 B.n101 B.n35 71.676
R713 B.n105 B.n36 71.676
R714 B.n109 B.n37 71.676
R715 B.n113 B.n38 71.676
R716 B.n117 B.n39 71.676
R717 B.n121 B.n40 71.676
R718 B.n125 B.n41 71.676
R719 B.n129 B.n42 71.676
R720 B.n133 B.n43 71.676
R721 B.n137 B.n44 71.676
R722 B.n141 B.n45 71.676
R723 B.n145 B.n46 71.676
R724 B.n149 B.n47 71.676
R725 B.n153 B.n48 71.676
R726 B.n157 B.n49 71.676
R727 B.n161 B.n50 71.676
R728 B.n165 B.n51 71.676
R729 B.n169 B.n52 71.676
R730 B.n173 B.n53 71.676
R731 B.n177 B.n54 71.676
R732 B.n181 B.n55 71.676
R733 B.n185 B.n56 71.676
R734 B.n189 B.n57 71.676
R735 B.n193 B.n58 71.676
R736 B.n197 B.n59 71.676
R737 B.n201 B.n60 71.676
R738 B.n205 B.n61 71.676
R739 B.n209 B.n62 71.676
R740 B.n213 B.n63 71.676
R741 B.n217 B.n64 71.676
R742 B.n221 B.n65 71.676
R743 B.n225 B.n66 71.676
R744 B.n229 B.n67 71.676
R745 B.n234 B.n68 71.676
R746 B.n238 B.n69 71.676
R747 B.n242 B.n70 71.676
R748 B.n246 B.n71 71.676
R749 B.n250 B.n72 71.676
R750 B.n254 B.n73 71.676
R751 B.n258 B.n74 71.676
R752 B.n262 B.n75 71.676
R753 B.n266 B.n76 71.676
R754 B.n270 B.n77 71.676
R755 B.n274 B.n78 71.676
R756 B.n278 B.n79 71.676
R757 B.n282 B.n80 71.676
R758 B.n286 B.n81 71.676
R759 B.n290 B.n82 71.676
R760 B.n294 B.n83 71.676
R761 B.n298 B.n84 71.676
R762 B.n302 B.n85 71.676
R763 B.n306 B.n86 71.676
R764 B.n310 B.n87 71.676
R765 B.n314 B.n88 71.676
R766 B.n318 B.n89 71.676
R767 B.n322 B.n90 71.676
R768 B.n326 B.n91 71.676
R769 B.n330 B.n92 71.676
R770 B.n334 B.n93 71.676
R771 B.n338 B.n94 71.676
R772 B.n95 B.n94 71.676
R773 B.n337 B.n93 71.676
R774 B.n333 B.n92 71.676
R775 B.n329 B.n91 71.676
R776 B.n325 B.n90 71.676
R777 B.n321 B.n89 71.676
R778 B.n317 B.n88 71.676
R779 B.n313 B.n87 71.676
R780 B.n309 B.n86 71.676
R781 B.n305 B.n85 71.676
R782 B.n301 B.n84 71.676
R783 B.n297 B.n83 71.676
R784 B.n293 B.n82 71.676
R785 B.n289 B.n81 71.676
R786 B.n285 B.n80 71.676
R787 B.n281 B.n79 71.676
R788 B.n277 B.n78 71.676
R789 B.n273 B.n77 71.676
R790 B.n269 B.n76 71.676
R791 B.n265 B.n75 71.676
R792 B.n261 B.n74 71.676
R793 B.n257 B.n73 71.676
R794 B.n253 B.n72 71.676
R795 B.n249 B.n71 71.676
R796 B.n245 B.n70 71.676
R797 B.n241 B.n69 71.676
R798 B.n237 B.n68 71.676
R799 B.n233 B.n67 71.676
R800 B.n228 B.n66 71.676
R801 B.n224 B.n65 71.676
R802 B.n220 B.n64 71.676
R803 B.n216 B.n63 71.676
R804 B.n212 B.n62 71.676
R805 B.n208 B.n61 71.676
R806 B.n204 B.n60 71.676
R807 B.n200 B.n59 71.676
R808 B.n196 B.n58 71.676
R809 B.n192 B.n57 71.676
R810 B.n188 B.n56 71.676
R811 B.n184 B.n55 71.676
R812 B.n180 B.n54 71.676
R813 B.n176 B.n53 71.676
R814 B.n172 B.n52 71.676
R815 B.n168 B.n51 71.676
R816 B.n164 B.n50 71.676
R817 B.n160 B.n49 71.676
R818 B.n156 B.n48 71.676
R819 B.n152 B.n47 71.676
R820 B.n148 B.n46 71.676
R821 B.n144 B.n45 71.676
R822 B.n140 B.n44 71.676
R823 B.n136 B.n43 71.676
R824 B.n132 B.n42 71.676
R825 B.n128 B.n41 71.676
R826 B.n124 B.n40 71.676
R827 B.n120 B.n39 71.676
R828 B.n116 B.n38 71.676
R829 B.n112 B.n37 71.676
R830 B.n108 B.n36 71.676
R831 B.n104 B.n35 71.676
R832 B.n677 B.n676 71.676
R833 B.n671 B.n375 71.676
R834 B.n668 B.n376 71.676
R835 B.n664 B.n377 71.676
R836 B.n660 B.n378 71.676
R837 B.n656 B.n379 71.676
R838 B.n652 B.n380 71.676
R839 B.n648 B.n381 71.676
R840 B.n644 B.n382 71.676
R841 B.n640 B.n383 71.676
R842 B.n636 B.n384 71.676
R843 B.n632 B.n385 71.676
R844 B.n628 B.n386 71.676
R845 B.n624 B.n387 71.676
R846 B.n620 B.n388 71.676
R847 B.n616 B.n389 71.676
R848 B.n612 B.n390 71.676
R849 B.n608 B.n391 71.676
R850 B.n604 B.n392 71.676
R851 B.n600 B.n393 71.676
R852 B.n596 B.n394 71.676
R853 B.n592 B.n395 71.676
R854 B.n588 B.n396 71.676
R855 B.n584 B.n397 71.676
R856 B.n580 B.n398 71.676
R857 B.n576 B.n399 71.676
R858 B.n572 B.n400 71.676
R859 B.n568 B.n401 71.676
R860 B.n563 B.n402 71.676
R861 B.n559 B.n403 71.676
R862 B.n555 B.n404 71.676
R863 B.n551 B.n405 71.676
R864 B.n547 B.n406 71.676
R865 B.n543 B.n407 71.676
R866 B.n539 B.n408 71.676
R867 B.n535 B.n409 71.676
R868 B.n531 B.n410 71.676
R869 B.n527 B.n411 71.676
R870 B.n523 B.n412 71.676
R871 B.n519 B.n413 71.676
R872 B.n515 B.n414 71.676
R873 B.n511 B.n415 71.676
R874 B.n507 B.n416 71.676
R875 B.n503 B.n417 71.676
R876 B.n499 B.n418 71.676
R877 B.n495 B.n419 71.676
R878 B.n491 B.n420 71.676
R879 B.n487 B.n421 71.676
R880 B.n483 B.n422 71.676
R881 B.n479 B.n423 71.676
R882 B.n475 B.n424 71.676
R883 B.n471 B.n425 71.676
R884 B.n467 B.n426 71.676
R885 B.n463 B.n427 71.676
R886 B.n459 B.n428 71.676
R887 B.n455 B.n429 71.676
R888 B.n451 B.n430 71.676
R889 B.n447 B.n431 71.676
R890 B.n443 B.n432 71.676
R891 B.n679 B.n374 71.676
R892 B.n677 B.n434 71.676
R893 B.n669 B.n375 71.676
R894 B.n665 B.n376 71.676
R895 B.n661 B.n377 71.676
R896 B.n657 B.n378 71.676
R897 B.n653 B.n379 71.676
R898 B.n649 B.n380 71.676
R899 B.n645 B.n381 71.676
R900 B.n641 B.n382 71.676
R901 B.n637 B.n383 71.676
R902 B.n633 B.n384 71.676
R903 B.n629 B.n385 71.676
R904 B.n625 B.n386 71.676
R905 B.n621 B.n387 71.676
R906 B.n617 B.n388 71.676
R907 B.n613 B.n389 71.676
R908 B.n609 B.n390 71.676
R909 B.n605 B.n391 71.676
R910 B.n601 B.n392 71.676
R911 B.n597 B.n393 71.676
R912 B.n593 B.n394 71.676
R913 B.n589 B.n395 71.676
R914 B.n585 B.n396 71.676
R915 B.n581 B.n397 71.676
R916 B.n577 B.n398 71.676
R917 B.n573 B.n399 71.676
R918 B.n569 B.n400 71.676
R919 B.n564 B.n401 71.676
R920 B.n560 B.n402 71.676
R921 B.n556 B.n403 71.676
R922 B.n552 B.n404 71.676
R923 B.n548 B.n405 71.676
R924 B.n544 B.n406 71.676
R925 B.n540 B.n407 71.676
R926 B.n536 B.n408 71.676
R927 B.n532 B.n409 71.676
R928 B.n528 B.n410 71.676
R929 B.n524 B.n411 71.676
R930 B.n520 B.n412 71.676
R931 B.n516 B.n413 71.676
R932 B.n512 B.n414 71.676
R933 B.n508 B.n415 71.676
R934 B.n504 B.n416 71.676
R935 B.n500 B.n417 71.676
R936 B.n496 B.n418 71.676
R937 B.n492 B.n419 71.676
R938 B.n488 B.n420 71.676
R939 B.n484 B.n421 71.676
R940 B.n480 B.n422 71.676
R941 B.n476 B.n423 71.676
R942 B.n472 B.n424 71.676
R943 B.n468 B.n425 71.676
R944 B.n464 B.n426 71.676
R945 B.n460 B.n427 71.676
R946 B.n456 B.n428 71.676
R947 B.n452 B.n429 71.676
R948 B.n448 B.n430 71.676
R949 B.n444 B.n431 71.676
R950 B.n440 B.n432 71.676
R951 B.n680 B.n679 71.676
R952 B.n796 B.n795 71.676
R953 B.n796 B.n2 71.676
R954 B.n678 B.n371 70.4205
R955 B.n760 B.n759 70.4205
R956 B.n100 B.n99 59.5399
R957 B.n231 B.n97 59.5399
R958 B.n439 B.n438 59.5399
R959 B.n566 B.n436 59.5399
R960 B.n685 B.n371 33.9619
R961 B.n685 B.n367 33.9619
R962 B.n691 B.n367 33.9619
R963 B.n691 B.n363 33.9619
R964 B.n697 B.n363 33.9619
R965 B.n703 B.n359 33.9619
R966 B.n703 B.n355 33.9619
R967 B.n709 B.n355 33.9619
R968 B.n709 B.n351 33.9619
R969 B.n715 B.n351 33.9619
R970 B.n715 B.n347 33.9619
R971 B.n722 B.n347 33.9619
R972 B.n728 B.n343 33.9619
R973 B.n728 B.n4 33.9619
R974 B.n794 B.n4 33.9619
R975 B.n794 B.n793 33.9619
R976 B.n793 B.n792 33.9619
R977 B.n792 B.n8 33.9619
R978 B.n737 B.n8 33.9619
R979 B.n785 B.n784 33.9619
R980 B.n784 B.n783 33.9619
R981 B.n783 B.n15 33.9619
R982 B.n777 B.n15 33.9619
R983 B.n777 B.n776 33.9619
R984 B.n776 B.n775 33.9619
R985 B.n775 B.n22 33.9619
R986 B.n769 B.n768 33.9619
R987 B.n768 B.n767 33.9619
R988 B.n767 B.n29 33.9619
R989 B.n761 B.n29 33.9619
R990 B.n761 B.n760 33.9619
R991 B.n675 B.n369 33.8737
R992 B.n682 B.n681 33.8737
R993 B.n757 B.n756 33.8737
R994 B.n102 B.n31 33.8737
R995 B.n99 B.n98 31.8066
R996 B.n97 B.n96 31.8066
R997 B.n438 B.n437 31.8066
R998 B.n436 B.n435 31.8066
R999 B.t10 B.n359 18.4795
R1000 B.t3 B.n22 18.4795
R1001 B B.n797 18.0485
R1002 B.t0 B.n343 17.4806
R1003 B.n737 B.t1 17.4806
R1004 B.n722 B.t0 16.4818
R1005 B.n785 B.t1 16.4818
R1006 B.n697 B.t10 15.4829
R1007 B.n769 B.t3 15.4829
R1008 B.n687 B.n369 10.6151
R1009 B.n688 B.n687 10.6151
R1010 B.n689 B.n688 10.6151
R1011 B.n689 B.n361 10.6151
R1012 B.n699 B.n361 10.6151
R1013 B.n700 B.n699 10.6151
R1014 B.n701 B.n700 10.6151
R1015 B.n701 B.n353 10.6151
R1016 B.n711 B.n353 10.6151
R1017 B.n712 B.n711 10.6151
R1018 B.n713 B.n712 10.6151
R1019 B.n713 B.n345 10.6151
R1020 B.n724 B.n345 10.6151
R1021 B.n725 B.n724 10.6151
R1022 B.n726 B.n725 10.6151
R1023 B.n726 B.n0 10.6151
R1024 B.n675 B.n674 10.6151
R1025 B.n674 B.n673 10.6151
R1026 B.n673 B.n672 10.6151
R1027 B.n672 B.n670 10.6151
R1028 B.n670 B.n667 10.6151
R1029 B.n667 B.n666 10.6151
R1030 B.n666 B.n663 10.6151
R1031 B.n663 B.n662 10.6151
R1032 B.n662 B.n659 10.6151
R1033 B.n659 B.n658 10.6151
R1034 B.n658 B.n655 10.6151
R1035 B.n655 B.n654 10.6151
R1036 B.n654 B.n651 10.6151
R1037 B.n651 B.n650 10.6151
R1038 B.n650 B.n647 10.6151
R1039 B.n647 B.n646 10.6151
R1040 B.n646 B.n643 10.6151
R1041 B.n643 B.n642 10.6151
R1042 B.n642 B.n639 10.6151
R1043 B.n639 B.n638 10.6151
R1044 B.n638 B.n635 10.6151
R1045 B.n635 B.n634 10.6151
R1046 B.n634 B.n631 10.6151
R1047 B.n631 B.n630 10.6151
R1048 B.n630 B.n627 10.6151
R1049 B.n627 B.n626 10.6151
R1050 B.n626 B.n623 10.6151
R1051 B.n623 B.n622 10.6151
R1052 B.n622 B.n619 10.6151
R1053 B.n619 B.n618 10.6151
R1054 B.n618 B.n615 10.6151
R1055 B.n615 B.n614 10.6151
R1056 B.n614 B.n611 10.6151
R1057 B.n611 B.n610 10.6151
R1058 B.n610 B.n607 10.6151
R1059 B.n607 B.n606 10.6151
R1060 B.n606 B.n603 10.6151
R1061 B.n603 B.n602 10.6151
R1062 B.n602 B.n599 10.6151
R1063 B.n599 B.n598 10.6151
R1064 B.n598 B.n595 10.6151
R1065 B.n595 B.n594 10.6151
R1066 B.n594 B.n591 10.6151
R1067 B.n591 B.n590 10.6151
R1068 B.n590 B.n587 10.6151
R1069 B.n587 B.n586 10.6151
R1070 B.n586 B.n583 10.6151
R1071 B.n583 B.n582 10.6151
R1072 B.n582 B.n579 10.6151
R1073 B.n579 B.n578 10.6151
R1074 B.n578 B.n575 10.6151
R1075 B.n575 B.n574 10.6151
R1076 B.n574 B.n571 10.6151
R1077 B.n571 B.n570 10.6151
R1078 B.n570 B.n567 10.6151
R1079 B.n565 B.n562 10.6151
R1080 B.n562 B.n561 10.6151
R1081 B.n561 B.n558 10.6151
R1082 B.n558 B.n557 10.6151
R1083 B.n557 B.n554 10.6151
R1084 B.n554 B.n553 10.6151
R1085 B.n553 B.n550 10.6151
R1086 B.n550 B.n549 10.6151
R1087 B.n546 B.n545 10.6151
R1088 B.n545 B.n542 10.6151
R1089 B.n542 B.n541 10.6151
R1090 B.n541 B.n538 10.6151
R1091 B.n538 B.n537 10.6151
R1092 B.n537 B.n534 10.6151
R1093 B.n534 B.n533 10.6151
R1094 B.n533 B.n530 10.6151
R1095 B.n530 B.n529 10.6151
R1096 B.n529 B.n526 10.6151
R1097 B.n526 B.n525 10.6151
R1098 B.n525 B.n522 10.6151
R1099 B.n522 B.n521 10.6151
R1100 B.n521 B.n518 10.6151
R1101 B.n518 B.n517 10.6151
R1102 B.n517 B.n514 10.6151
R1103 B.n514 B.n513 10.6151
R1104 B.n513 B.n510 10.6151
R1105 B.n510 B.n509 10.6151
R1106 B.n509 B.n506 10.6151
R1107 B.n506 B.n505 10.6151
R1108 B.n505 B.n502 10.6151
R1109 B.n502 B.n501 10.6151
R1110 B.n501 B.n498 10.6151
R1111 B.n498 B.n497 10.6151
R1112 B.n497 B.n494 10.6151
R1113 B.n494 B.n493 10.6151
R1114 B.n493 B.n490 10.6151
R1115 B.n490 B.n489 10.6151
R1116 B.n489 B.n486 10.6151
R1117 B.n486 B.n485 10.6151
R1118 B.n485 B.n482 10.6151
R1119 B.n482 B.n481 10.6151
R1120 B.n481 B.n478 10.6151
R1121 B.n478 B.n477 10.6151
R1122 B.n477 B.n474 10.6151
R1123 B.n474 B.n473 10.6151
R1124 B.n473 B.n470 10.6151
R1125 B.n470 B.n469 10.6151
R1126 B.n469 B.n466 10.6151
R1127 B.n466 B.n465 10.6151
R1128 B.n465 B.n462 10.6151
R1129 B.n462 B.n461 10.6151
R1130 B.n461 B.n458 10.6151
R1131 B.n458 B.n457 10.6151
R1132 B.n457 B.n454 10.6151
R1133 B.n454 B.n453 10.6151
R1134 B.n453 B.n450 10.6151
R1135 B.n450 B.n449 10.6151
R1136 B.n449 B.n446 10.6151
R1137 B.n446 B.n445 10.6151
R1138 B.n445 B.n442 10.6151
R1139 B.n442 B.n441 10.6151
R1140 B.n441 B.n373 10.6151
R1141 B.n681 B.n373 10.6151
R1142 B.n683 B.n682 10.6151
R1143 B.n683 B.n365 10.6151
R1144 B.n693 B.n365 10.6151
R1145 B.n694 B.n693 10.6151
R1146 B.n695 B.n694 10.6151
R1147 B.n695 B.n357 10.6151
R1148 B.n705 B.n357 10.6151
R1149 B.n706 B.n705 10.6151
R1150 B.n707 B.n706 10.6151
R1151 B.n707 B.n349 10.6151
R1152 B.n717 B.n349 10.6151
R1153 B.n718 B.n717 10.6151
R1154 B.n720 B.n718 10.6151
R1155 B.n720 B.n719 10.6151
R1156 B.n719 B.n341 10.6151
R1157 B.n731 B.n341 10.6151
R1158 B.n732 B.n731 10.6151
R1159 B.n733 B.n732 10.6151
R1160 B.n734 B.n733 10.6151
R1161 B.n735 B.n734 10.6151
R1162 B.n739 B.n735 10.6151
R1163 B.n740 B.n739 10.6151
R1164 B.n741 B.n740 10.6151
R1165 B.n742 B.n741 10.6151
R1166 B.n744 B.n742 10.6151
R1167 B.n745 B.n744 10.6151
R1168 B.n746 B.n745 10.6151
R1169 B.n747 B.n746 10.6151
R1170 B.n749 B.n747 10.6151
R1171 B.n750 B.n749 10.6151
R1172 B.n751 B.n750 10.6151
R1173 B.n752 B.n751 10.6151
R1174 B.n754 B.n752 10.6151
R1175 B.n755 B.n754 10.6151
R1176 B.n756 B.n755 10.6151
R1177 B.n789 B.n1 10.6151
R1178 B.n789 B.n788 10.6151
R1179 B.n788 B.n787 10.6151
R1180 B.n787 B.n10 10.6151
R1181 B.n781 B.n10 10.6151
R1182 B.n781 B.n780 10.6151
R1183 B.n780 B.n779 10.6151
R1184 B.n779 B.n17 10.6151
R1185 B.n773 B.n17 10.6151
R1186 B.n773 B.n772 10.6151
R1187 B.n772 B.n771 10.6151
R1188 B.n771 B.n24 10.6151
R1189 B.n765 B.n24 10.6151
R1190 B.n765 B.n764 10.6151
R1191 B.n764 B.n763 10.6151
R1192 B.n763 B.n31 10.6151
R1193 B.n103 B.n102 10.6151
R1194 B.n106 B.n103 10.6151
R1195 B.n107 B.n106 10.6151
R1196 B.n110 B.n107 10.6151
R1197 B.n111 B.n110 10.6151
R1198 B.n114 B.n111 10.6151
R1199 B.n115 B.n114 10.6151
R1200 B.n118 B.n115 10.6151
R1201 B.n119 B.n118 10.6151
R1202 B.n122 B.n119 10.6151
R1203 B.n123 B.n122 10.6151
R1204 B.n126 B.n123 10.6151
R1205 B.n127 B.n126 10.6151
R1206 B.n130 B.n127 10.6151
R1207 B.n131 B.n130 10.6151
R1208 B.n134 B.n131 10.6151
R1209 B.n135 B.n134 10.6151
R1210 B.n138 B.n135 10.6151
R1211 B.n139 B.n138 10.6151
R1212 B.n142 B.n139 10.6151
R1213 B.n143 B.n142 10.6151
R1214 B.n146 B.n143 10.6151
R1215 B.n147 B.n146 10.6151
R1216 B.n150 B.n147 10.6151
R1217 B.n151 B.n150 10.6151
R1218 B.n154 B.n151 10.6151
R1219 B.n155 B.n154 10.6151
R1220 B.n158 B.n155 10.6151
R1221 B.n159 B.n158 10.6151
R1222 B.n162 B.n159 10.6151
R1223 B.n163 B.n162 10.6151
R1224 B.n166 B.n163 10.6151
R1225 B.n167 B.n166 10.6151
R1226 B.n170 B.n167 10.6151
R1227 B.n171 B.n170 10.6151
R1228 B.n174 B.n171 10.6151
R1229 B.n175 B.n174 10.6151
R1230 B.n178 B.n175 10.6151
R1231 B.n179 B.n178 10.6151
R1232 B.n182 B.n179 10.6151
R1233 B.n183 B.n182 10.6151
R1234 B.n186 B.n183 10.6151
R1235 B.n187 B.n186 10.6151
R1236 B.n190 B.n187 10.6151
R1237 B.n191 B.n190 10.6151
R1238 B.n194 B.n191 10.6151
R1239 B.n195 B.n194 10.6151
R1240 B.n198 B.n195 10.6151
R1241 B.n199 B.n198 10.6151
R1242 B.n202 B.n199 10.6151
R1243 B.n203 B.n202 10.6151
R1244 B.n206 B.n203 10.6151
R1245 B.n207 B.n206 10.6151
R1246 B.n210 B.n207 10.6151
R1247 B.n211 B.n210 10.6151
R1248 B.n215 B.n214 10.6151
R1249 B.n218 B.n215 10.6151
R1250 B.n219 B.n218 10.6151
R1251 B.n222 B.n219 10.6151
R1252 B.n223 B.n222 10.6151
R1253 B.n226 B.n223 10.6151
R1254 B.n227 B.n226 10.6151
R1255 B.n230 B.n227 10.6151
R1256 B.n235 B.n232 10.6151
R1257 B.n236 B.n235 10.6151
R1258 B.n239 B.n236 10.6151
R1259 B.n240 B.n239 10.6151
R1260 B.n243 B.n240 10.6151
R1261 B.n244 B.n243 10.6151
R1262 B.n247 B.n244 10.6151
R1263 B.n248 B.n247 10.6151
R1264 B.n251 B.n248 10.6151
R1265 B.n252 B.n251 10.6151
R1266 B.n255 B.n252 10.6151
R1267 B.n256 B.n255 10.6151
R1268 B.n259 B.n256 10.6151
R1269 B.n260 B.n259 10.6151
R1270 B.n263 B.n260 10.6151
R1271 B.n264 B.n263 10.6151
R1272 B.n267 B.n264 10.6151
R1273 B.n268 B.n267 10.6151
R1274 B.n271 B.n268 10.6151
R1275 B.n272 B.n271 10.6151
R1276 B.n275 B.n272 10.6151
R1277 B.n276 B.n275 10.6151
R1278 B.n279 B.n276 10.6151
R1279 B.n280 B.n279 10.6151
R1280 B.n283 B.n280 10.6151
R1281 B.n284 B.n283 10.6151
R1282 B.n287 B.n284 10.6151
R1283 B.n288 B.n287 10.6151
R1284 B.n291 B.n288 10.6151
R1285 B.n292 B.n291 10.6151
R1286 B.n295 B.n292 10.6151
R1287 B.n296 B.n295 10.6151
R1288 B.n299 B.n296 10.6151
R1289 B.n300 B.n299 10.6151
R1290 B.n303 B.n300 10.6151
R1291 B.n304 B.n303 10.6151
R1292 B.n307 B.n304 10.6151
R1293 B.n308 B.n307 10.6151
R1294 B.n311 B.n308 10.6151
R1295 B.n312 B.n311 10.6151
R1296 B.n315 B.n312 10.6151
R1297 B.n316 B.n315 10.6151
R1298 B.n319 B.n316 10.6151
R1299 B.n320 B.n319 10.6151
R1300 B.n323 B.n320 10.6151
R1301 B.n324 B.n323 10.6151
R1302 B.n327 B.n324 10.6151
R1303 B.n328 B.n327 10.6151
R1304 B.n331 B.n328 10.6151
R1305 B.n332 B.n331 10.6151
R1306 B.n335 B.n332 10.6151
R1307 B.n336 B.n335 10.6151
R1308 B.n339 B.n336 10.6151
R1309 B.n340 B.n339 10.6151
R1310 B.n757 B.n340 10.6151
R1311 B.n797 B.n0 8.11757
R1312 B.n797 B.n1 8.11757
R1313 B.n566 B.n565 6.5566
R1314 B.n549 B.n439 6.5566
R1315 B.n214 B.n100 6.5566
R1316 B.n231 B.n230 6.5566
R1317 B.n567 B.n566 4.05904
R1318 B.n546 B.n439 4.05904
R1319 B.n211 B.n100 4.05904
R1320 B.n232 B.n231 4.05904
R1321 VP.n0 VP.t1 463.757
R1322 VP.n0 VP.t0 418.923
R1323 VP VP.n0 0.146778
R1324 VTAIL.n370 VTAIL.n282 289.615
R1325 VTAIL.n88 VTAIL.n0 289.615
R1326 VTAIL.n276 VTAIL.n188 289.615
R1327 VTAIL.n182 VTAIL.n94 289.615
R1328 VTAIL.n313 VTAIL.n312 185
R1329 VTAIL.n310 VTAIL.n309 185
R1330 VTAIL.n319 VTAIL.n318 185
R1331 VTAIL.n321 VTAIL.n320 185
R1332 VTAIL.n306 VTAIL.n305 185
R1333 VTAIL.n327 VTAIL.n326 185
R1334 VTAIL.n329 VTAIL.n328 185
R1335 VTAIL.n302 VTAIL.n301 185
R1336 VTAIL.n335 VTAIL.n334 185
R1337 VTAIL.n337 VTAIL.n336 185
R1338 VTAIL.n298 VTAIL.n297 185
R1339 VTAIL.n343 VTAIL.n342 185
R1340 VTAIL.n345 VTAIL.n344 185
R1341 VTAIL.n294 VTAIL.n293 185
R1342 VTAIL.n351 VTAIL.n350 185
R1343 VTAIL.n354 VTAIL.n353 185
R1344 VTAIL.n352 VTAIL.n290 185
R1345 VTAIL.n359 VTAIL.n289 185
R1346 VTAIL.n361 VTAIL.n360 185
R1347 VTAIL.n363 VTAIL.n362 185
R1348 VTAIL.n286 VTAIL.n285 185
R1349 VTAIL.n369 VTAIL.n368 185
R1350 VTAIL.n371 VTAIL.n370 185
R1351 VTAIL.n31 VTAIL.n30 185
R1352 VTAIL.n28 VTAIL.n27 185
R1353 VTAIL.n37 VTAIL.n36 185
R1354 VTAIL.n39 VTAIL.n38 185
R1355 VTAIL.n24 VTAIL.n23 185
R1356 VTAIL.n45 VTAIL.n44 185
R1357 VTAIL.n47 VTAIL.n46 185
R1358 VTAIL.n20 VTAIL.n19 185
R1359 VTAIL.n53 VTAIL.n52 185
R1360 VTAIL.n55 VTAIL.n54 185
R1361 VTAIL.n16 VTAIL.n15 185
R1362 VTAIL.n61 VTAIL.n60 185
R1363 VTAIL.n63 VTAIL.n62 185
R1364 VTAIL.n12 VTAIL.n11 185
R1365 VTAIL.n69 VTAIL.n68 185
R1366 VTAIL.n72 VTAIL.n71 185
R1367 VTAIL.n70 VTAIL.n8 185
R1368 VTAIL.n77 VTAIL.n7 185
R1369 VTAIL.n79 VTAIL.n78 185
R1370 VTAIL.n81 VTAIL.n80 185
R1371 VTAIL.n4 VTAIL.n3 185
R1372 VTAIL.n87 VTAIL.n86 185
R1373 VTAIL.n89 VTAIL.n88 185
R1374 VTAIL.n277 VTAIL.n276 185
R1375 VTAIL.n275 VTAIL.n274 185
R1376 VTAIL.n192 VTAIL.n191 185
R1377 VTAIL.n269 VTAIL.n268 185
R1378 VTAIL.n267 VTAIL.n266 185
R1379 VTAIL.n265 VTAIL.n195 185
R1380 VTAIL.n199 VTAIL.n196 185
R1381 VTAIL.n260 VTAIL.n259 185
R1382 VTAIL.n258 VTAIL.n257 185
R1383 VTAIL.n201 VTAIL.n200 185
R1384 VTAIL.n252 VTAIL.n251 185
R1385 VTAIL.n250 VTAIL.n249 185
R1386 VTAIL.n205 VTAIL.n204 185
R1387 VTAIL.n244 VTAIL.n243 185
R1388 VTAIL.n242 VTAIL.n241 185
R1389 VTAIL.n209 VTAIL.n208 185
R1390 VTAIL.n236 VTAIL.n235 185
R1391 VTAIL.n234 VTAIL.n233 185
R1392 VTAIL.n213 VTAIL.n212 185
R1393 VTAIL.n228 VTAIL.n227 185
R1394 VTAIL.n226 VTAIL.n225 185
R1395 VTAIL.n217 VTAIL.n216 185
R1396 VTAIL.n220 VTAIL.n219 185
R1397 VTAIL.n183 VTAIL.n182 185
R1398 VTAIL.n181 VTAIL.n180 185
R1399 VTAIL.n98 VTAIL.n97 185
R1400 VTAIL.n175 VTAIL.n174 185
R1401 VTAIL.n173 VTAIL.n172 185
R1402 VTAIL.n171 VTAIL.n101 185
R1403 VTAIL.n105 VTAIL.n102 185
R1404 VTAIL.n166 VTAIL.n165 185
R1405 VTAIL.n164 VTAIL.n163 185
R1406 VTAIL.n107 VTAIL.n106 185
R1407 VTAIL.n158 VTAIL.n157 185
R1408 VTAIL.n156 VTAIL.n155 185
R1409 VTAIL.n111 VTAIL.n110 185
R1410 VTAIL.n150 VTAIL.n149 185
R1411 VTAIL.n148 VTAIL.n147 185
R1412 VTAIL.n115 VTAIL.n114 185
R1413 VTAIL.n142 VTAIL.n141 185
R1414 VTAIL.n140 VTAIL.n139 185
R1415 VTAIL.n119 VTAIL.n118 185
R1416 VTAIL.n134 VTAIL.n133 185
R1417 VTAIL.n132 VTAIL.n131 185
R1418 VTAIL.n123 VTAIL.n122 185
R1419 VTAIL.n126 VTAIL.n125 185
R1420 VTAIL.t2 VTAIL.n218 147.659
R1421 VTAIL.t0 VTAIL.n124 147.659
R1422 VTAIL.t1 VTAIL.n311 147.659
R1423 VTAIL.t3 VTAIL.n29 147.659
R1424 VTAIL.n312 VTAIL.n309 104.615
R1425 VTAIL.n319 VTAIL.n309 104.615
R1426 VTAIL.n320 VTAIL.n319 104.615
R1427 VTAIL.n320 VTAIL.n305 104.615
R1428 VTAIL.n327 VTAIL.n305 104.615
R1429 VTAIL.n328 VTAIL.n327 104.615
R1430 VTAIL.n328 VTAIL.n301 104.615
R1431 VTAIL.n335 VTAIL.n301 104.615
R1432 VTAIL.n336 VTAIL.n335 104.615
R1433 VTAIL.n336 VTAIL.n297 104.615
R1434 VTAIL.n343 VTAIL.n297 104.615
R1435 VTAIL.n344 VTAIL.n343 104.615
R1436 VTAIL.n344 VTAIL.n293 104.615
R1437 VTAIL.n351 VTAIL.n293 104.615
R1438 VTAIL.n353 VTAIL.n351 104.615
R1439 VTAIL.n353 VTAIL.n352 104.615
R1440 VTAIL.n352 VTAIL.n289 104.615
R1441 VTAIL.n361 VTAIL.n289 104.615
R1442 VTAIL.n362 VTAIL.n361 104.615
R1443 VTAIL.n362 VTAIL.n285 104.615
R1444 VTAIL.n369 VTAIL.n285 104.615
R1445 VTAIL.n370 VTAIL.n369 104.615
R1446 VTAIL.n30 VTAIL.n27 104.615
R1447 VTAIL.n37 VTAIL.n27 104.615
R1448 VTAIL.n38 VTAIL.n37 104.615
R1449 VTAIL.n38 VTAIL.n23 104.615
R1450 VTAIL.n45 VTAIL.n23 104.615
R1451 VTAIL.n46 VTAIL.n45 104.615
R1452 VTAIL.n46 VTAIL.n19 104.615
R1453 VTAIL.n53 VTAIL.n19 104.615
R1454 VTAIL.n54 VTAIL.n53 104.615
R1455 VTAIL.n54 VTAIL.n15 104.615
R1456 VTAIL.n61 VTAIL.n15 104.615
R1457 VTAIL.n62 VTAIL.n61 104.615
R1458 VTAIL.n62 VTAIL.n11 104.615
R1459 VTAIL.n69 VTAIL.n11 104.615
R1460 VTAIL.n71 VTAIL.n69 104.615
R1461 VTAIL.n71 VTAIL.n70 104.615
R1462 VTAIL.n70 VTAIL.n7 104.615
R1463 VTAIL.n79 VTAIL.n7 104.615
R1464 VTAIL.n80 VTAIL.n79 104.615
R1465 VTAIL.n80 VTAIL.n3 104.615
R1466 VTAIL.n87 VTAIL.n3 104.615
R1467 VTAIL.n88 VTAIL.n87 104.615
R1468 VTAIL.n276 VTAIL.n275 104.615
R1469 VTAIL.n275 VTAIL.n191 104.615
R1470 VTAIL.n268 VTAIL.n191 104.615
R1471 VTAIL.n268 VTAIL.n267 104.615
R1472 VTAIL.n267 VTAIL.n195 104.615
R1473 VTAIL.n199 VTAIL.n195 104.615
R1474 VTAIL.n259 VTAIL.n199 104.615
R1475 VTAIL.n259 VTAIL.n258 104.615
R1476 VTAIL.n258 VTAIL.n200 104.615
R1477 VTAIL.n251 VTAIL.n200 104.615
R1478 VTAIL.n251 VTAIL.n250 104.615
R1479 VTAIL.n250 VTAIL.n204 104.615
R1480 VTAIL.n243 VTAIL.n204 104.615
R1481 VTAIL.n243 VTAIL.n242 104.615
R1482 VTAIL.n242 VTAIL.n208 104.615
R1483 VTAIL.n235 VTAIL.n208 104.615
R1484 VTAIL.n235 VTAIL.n234 104.615
R1485 VTAIL.n234 VTAIL.n212 104.615
R1486 VTAIL.n227 VTAIL.n212 104.615
R1487 VTAIL.n227 VTAIL.n226 104.615
R1488 VTAIL.n226 VTAIL.n216 104.615
R1489 VTAIL.n219 VTAIL.n216 104.615
R1490 VTAIL.n182 VTAIL.n181 104.615
R1491 VTAIL.n181 VTAIL.n97 104.615
R1492 VTAIL.n174 VTAIL.n97 104.615
R1493 VTAIL.n174 VTAIL.n173 104.615
R1494 VTAIL.n173 VTAIL.n101 104.615
R1495 VTAIL.n105 VTAIL.n101 104.615
R1496 VTAIL.n165 VTAIL.n105 104.615
R1497 VTAIL.n165 VTAIL.n164 104.615
R1498 VTAIL.n164 VTAIL.n106 104.615
R1499 VTAIL.n157 VTAIL.n106 104.615
R1500 VTAIL.n157 VTAIL.n156 104.615
R1501 VTAIL.n156 VTAIL.n110 104.615
R1502 VTAIL.n149 VTAIL.n110 104.615
R1503 VTAIL.n149 VTAIL.n148 104.615
R1504 VTAIL.n148 VTAIL.n114 104.615
R1505 VTAIL.n141 VTAIL.n114 104.615
R1506 VTAIL.n141 VTAIL.n140 104.615
R1507 VTAIL.n140 VTAIL.n118 104.615
R1508 VTAIL.n133 VTAIL.n118 104.615
R1509 VTAIL.n133 VTAIL.n132 104.615
R1510 VTAIL.n132 VTAIL.n122 104.615
R1511 VTAIL.n125 VTAIL.n122 104.615
R1512 VTAIL.n312 VTAIL.t1 52.3082
R1513 VTAIL.n30 VTAIL.t3 52.3082
R1514 VTAIL.n219 VTAIL.t2 52.3082
R1515 VTAIL.n125 VTAIL.t0 52.3082
R1516 VTAIL.n375 VTAIL.n374 31.2157
R1517 VTAIL.n93 VTAIL.n92 31.2157
R1518 VTAIL.n281 VTAIL.n280 31.2157
R1519 VTAIL.n187 VTAIL.n186 31.2157
R1520 VTAIL.n187 VTAIL.n93 29.6341
R1521 VTAIL.n375 VTAIL.n281 28.2203
R1522 VTAIL.n313 VTAIL.n311 15.6677
R1523 VTAIL.n31 VTAIL.n29 15.6677
R1524 VTAIL.n220 VTAIL.n218 15.6677
R1525 VTAIL.n126 VTAIL.n124 15.6677
R1526 VTAIL.n360 VTAIL.n359 13.1884
R1527 VTAIL.n78 VTAIL.n77 13.1884
R1528 VTAIL.n266 VTAIL.n265 13.1884
R1529 VTAIL.n172 VTAIL.n171 13.1884
R1530 VTAIL.n314 VTAIL.n310 12.8005
R1531 VTAIL.n358 VTAIL.n290 12.8005
R1532 VTAIL.n363 VTAIL.n288 12.8005
R1533 VTAIL.n32 VTAIL.n28 12.8005
R1534 VTAIL.n76 VTAIL.n8 12.8005
R1535 VTAIL.n81 VTAIL.n6 12.8005
R1536 VTAIL.n269 VTAIL.n194 12.8005
R1537 VTAIL.n264 VTAIL.n196 12.8005
R1538 VTAIL.n221 VTAIL.n217 12.8005
R1539 VTAIL.n175 VTAIL.n100 12.8005
R1540 VTAIL.n170 VTAIL.n102 12.8005
R1541 VTAIL.n127 VTAIL.n123 12.8005
R1542 VTAIL.n318 VTAIL.n317 12.0247
R1543 VTAIL.n355 VTAIL.n354 12.0247
R1544 VTAIL.n364 VTAIL.n286 12.0247
R1545 VTAIL.n36 VTAIL.n35 12.0247
R1546 VTAIL.n73 VTAIL.n72 12.0247
R1547 VTAIL.n82 VTAIL.n4 12.0247
R1548 VTAIL.n270 VTAIL.n192 12.0247
R1549 VTAIL.n261 VTAIL.n260 12.0247
R1550 VTAIL.n225 VTAIL.n224 12.0247
R1551 VTAIL.n176 VTAIL.n98 12.0247
R1552 VTAIL.n167 VTAIL.n166 12.0247
R1553 VTAIL.n131 VTAIL.n130 12.0247
R1554 VTAIL.n321 VTAIL.n308 11.249
R1555 VTAIL.n350 VTAIL.n292 11.249
R1556 VTAIL.n368 VTAIL.n367 11.249
R1557 VTAIL.n39 VTAIL.n26 11.249
R1558 VTAIL.n68 VTAIL.n10 11.249
R1559 VTAIL.n86 VTAIL.n85 11.249
R1560 VTAIL.n274 VTAIL.n273 11.249
R1561 VTAIL.n257 VTAIL.n198 11.249
R1562 VTAIL.n228 VTAIL.n215 11.249
R1563 VTAIL.n180 VTAIL.n179 11.249
R1564 VTAIL.n163 VTAIL.n104 11.249
R1565 VTAIL.n134 VTAIL.n121 11.249
R1566 VTAIL.n322 VTAIL.n306 10.4732
R1567 VTAIL.n349 VTAIL.n294 10.4732
R1568 VTAIL.n371 VTAIL.n284 10.4732
R1569 VTAIL.n40 VTAIL.n24 10.4732
R1570 VTAIL.n67 VTAIL.n12 10.4732
R1571 VTAIL.n89 VTAIL.n2 10.4732
R1572 VTAIL.n277 VTAIL.n190 10.4732
R1573 VTAIL.n256 VTAIL.n201 10.4732
R1574 VTAIL.n229 VTAIL.n213 10.4732
R1575 VTAIL.n183 VTAIL.n96 10.4732
R1576 VTAIL.n162 VTAIL.n107 10.4732
R1577 VTAIL.n135 VTAIL.n119 10.4732
R1578 VTAIL.n326 VTAIL.n325 9.69747
R1579 VTAIL.n346 VTAIL.n345 9.69747
R1580 VTAIL.n372 VTAIL.n282 9.69747
R1581 VTAIL.n44 VTAIL.n43 9.69747
R1582 VTAIL.n64 VTAIL.n63 9.69747
R1583 VTAIL.n90 VTAIL.n0 9.69747
R1584 VTAIL.n278 VTAIL.n188 9.69747
R1585 VTAIL.n253 VTAIL.n252 9.69747
R1586 VTAIL.n233 VTAIL.n232 9.69747
R1587 VTAIL.n184 VTAIL.n94 9.69747
R1588 VTAIL.n159 VTAIL.n158 9.69747
R1589 VTAIL.n139 VTAIL.n138 9.69747
R1590 VTAIL.n374 VTAIL.n373 9.45567
R1591 VTAIL.n92 VTAIL.n91 9.45567
R1592 VTAIL.n280 VTAIL.n279 9.45567
R1593 VTAIL.n186 VTAIL.n185 9.45567
R1594 VTAIL.n373 VTAIL.n372 9.3005
R1595 VTAIL.n284 VTAIL.n283 9.3005
R1596 VTAIL.n367 VTAIL.n366 9.3005
R1597 VTAIL.n365 VTAIL.n364 9.3005
R1598 VTAIL.n288 VTAIL.n287 9.3005
R1599 VTAIL.n333 VTAIL.n332 9.3005
R1600 VTAIL.n331 VTAIL.n330 9.3005
R1601 VTAIL.n304 VTAIL.n303 9.3005
R1602 VTAIL.n325 VTAIL.n324 9.3005
R1603 VTAIL.n323 VTAIL.n322 9.3005
R1604 VTAIL.n308 VTAIL.n307 9.3005
R1605 VTAIL.n317 VTAIL.n316 9.3005
R1606 VTAIL.n315 VTAIL.n314 9.3005
R1607 VTAIL.n300 VTAIL.n299 9.3005
R1608 VTAIL.n339 VTAIL.n338 9.3005
R1609 VTAIL.n341 VTAIL.n340 9.3005
R1610 VTAIL.n296 VTAIL.n295 9.3005
R1611 VTAIL.n347 VTAIL.n346 9.3005
R1612 VTAIL.n349 VTAIL.n348 9.3005
R1613 VTAIL.n292 VTAIL.n291 9.3005
R1614 VTAIL.n356 VTAIL.n355 9.3005
R1615 VTAIL.n358 VTAIL.n357 9.3005
R1616 VTAIL.n91 VTAIL.n90 9.3005
R1617 VTAIL.n2 VTAIL.n1 9.3005
R1618 VTAIL.n85 VTAIL.n84 9.3005
R1619 VTAIL.n83 VTAIL.n82 9.3005
R1620 VTAIL.n6 VTAIL.n5 9.3005
R1621 VTAIL.n51 VTAIL.n50 9.3005
R1622 VTAIL.n49 VTAIL.n48 9.3005
R1623 VTAIL.n22 VTAIL.n21 9.3005
R1624 VTAIL.n43 VTAIL.n42 9.3005
R1625 VTAIL.n41 VTAIL.n40 9.3005
R1626 VTAIL.n26 VTAIL.n25 9.3005
R1627 VTAIL.n35 VTAIL.n34 9.3005
R1628 VTAIL.n33 VTAIL.n32 9.3005
R1629 VTAIL.n18 VTAIL.n17 9.3005
R1630 VTAIL.n57 VTAIL.n56 9.3005
R1631 VTAIL.n59 VTAIL.n58 9.3005
R1632 VTAIL.n14 VTAIL.n13 9.3005
R1633 VTAIL.n65 VTAIL.n64 9.3005
R1634 VTAIL.n67 VTAIL.n66 9.3005
R1635 VTAIL.n10 VTAIL.n9 9.3005
R1636 VTAIL.n74 VTAIL.n73 9.3005
R1637 VTAIL.n76 VTAIL.n75 9.3005
R1638 VTAIL.n246 VTAIL.n245 9.3005
R1639 VTAIL.n248 VTAIL.n247 9.3005
R1640 VTAIL.n203 VTAIL.n202 9.3005
R1641 VTAIL.n254 VTAIL.n253 9.3005
R1642 VTAIL.n256 VTAIL.n255 9.3005
R1643 VTAIL.n198 VTAIL.n197 9.3005
R1644 VTAIL.n262 VTAIL.n261 9.3005
R1645 VTAIL.n264 VTAIL.n263 9.3005
R1646 VTAIL.n279 VTAIL.n278 9.3005
R1647 VTAIL.n190 VTAIL.n189 9.3005
R1648 VTAIL.n273 VTAIL.n272 9.3005
R1649 VTAIL.n271 VTAIL.n270 9.3005
R1650 VTAIL.n194 VTAIL.n193 9.3005
R1651 VTAIL.n207 VTAIL.n206 9.3005
R1652 VTAIL.n240 VTAIL.n239 9.3005
R1653 VTAIL.n238 VTAIL.n237 9.3005
R1654 VTAIL.n211 VTAIL.n210 9.3005
R1655 VTAIL.n232 VTAIL.n231 9.3005
R1656 VTAIL.n230 VTAIL.n229 9.3005
R1657 VTAIL.n215 VTAIL.n214 9.3005
R1658 VTAIL.n224 VTAIL.n223 9.3005
R1659 VTAIL.n222 VTAIL.n221 9.3005
R1660 VTAIL.n152 VTAIL.n151 9.3005
R1661 VTAIL.n154 VTAIL.n153 9.3005
R1662 VTAIL.n109 VTAIL.n108 9.3005
R1663 VTAIL.n160 VTAIL.n159 9.3005
R1664 VTAIL.n162 VTAIL.n161 9.3005
R1665 VTAIL.n104 VTAIL.n103 9.3005
R1666 VTAIL.n168 VTAIL.n167 9.3005
R1667 VTAIL.n170 VTAIL.n169 9.3005
R1668 VTAIL.n185 VTAIL.n184 9.3005
R1669 VTAIL.n96 VTAIL.n95 9.3005
R1670 VTAIL.n179 VTAIL.n178 9.3005
R1671 VTAIL.n177 VTAIL.n176 9.3005
R1672 VTAIL.n100 VTAIL.n99 9.3005
R1673 VTAIL.n113 VTAIL.n112 9.3005
R1674 VTAIL.n146 VTAIL.n145 9.3005
R1675 VTAIL.n144 VTAIL.n143 9.3005
R1676 VTAIL.n117 VTAIL.n116 9.3005
R1677 VTAIL.n138 VTAIL.n137 9.3005
R1678 VTAIL.n136 VTAIL.n135 9.3005
R1679 VTAIL.n121 VTAIL.n120 9.3005
R1680 VTAIL.n130 VTAIL.n129 9.3005
R1681 VTAIL.n128 VTAIL.n127 9.3005
R1682 VTAIL.n329 VTAIL.n304 8.92171
R1683 VTAIL.n342 VTAIL.n296 8.92171
R1684 VTAIL.n47 VTAIL.n22 8.92171
R1685 VTAIL.n60 VTAIL.n14 8.92171
R1686 VTAIL.n249 VTAIL.n203 8.92171
R1687 VTAIL.n236 VTAIL.n211 8.92171
R1688 VTAIL.n155 VTAIL.n109 8.92171
R1689 VTAIL.n142 VTAIL.n117 8.92171
R1690 VTAIL.n330 VTAIL.n302 8.14595
R1691 VTAIL.n341 VTAIL.n298 8.14595
R1692 VTAIL.n48 VTAIL.n20 8.14595
R1693 VTAIL.n59 VTAIL.n16 8.14595
R1694 VTAIL.n248 VTAIL.n205 8.14595
R1695 VTAIL.n237 VTAIL.n209 8.14595
R1696 VTAIL.n154 VTAIL.n111 8.14595
R1697 VTAIL.n143 VTAIL.n115 8.14595
R1698 VTAIL.n334 VTAIL.n333 7.3702
R1699 VTAIL.n338 VTAIL.n337 7.3702
R1700 VTAIL.n52 VTAIL.n51 7.3702
R1701 VTAIL.n56 VTAIL.n55 7.3702
R1702 VTAIL.n245 VTAIL.n244 7.3702
R1703 VTAIL.n241 VTAIL.n240 7.3702
R1704 VTAIL.n151 VTAIL.n150 7.3702
R1705 VTAIL.n147 VTAIL.n146 7.3702
R1706 VTAIL.n334 VTAIL.n300 6.59444
R1707 VTAIL.n337 VTAIL.n300 6.59444
R1708 VTAIL.n52 VTAIL.n18 6.59444
R1709 VTAIL.n55 VTAIL.n18 6.59444
R1710 VTAIL.n244 VTAIL.n207 6.59444
R1711 VTAIL.n241 VTAIL.n207 6.59444
R1712 VTAIL.n150 VTAIL.n113 6.59444
R1713 VTAIL.n147 VTAIL.n113 6.59444
R1714 VTAIL.n333 VTAIL.n302 5.81868
R1715 VTAIL.n338 VTAIL.n298 5.81868
R1716 VTAIL.n51 VTAIL.n20 5.81868
R1717 VTAIL.n56 VTAIL.n16 5.81868
R1718 VTAIL.n245 VTAIL.n205 5.81868
R1719 VTAIL.n240 VTAIL.n209 5.81868
R1720 VTAIL.n151 VTAIL.n111 5.81868
R1721 VTAIL.n146 VTAIL.n115 5.81868
R1722 VTAIL.n330 VTAIL.n329 5.04292
R1723 VTAIL.n342 VTAIL.n341 5.04292
R1724 VTAIL.n48 VTAIL.n47 5.04292
R1725 VTAIL.n60 VTAIL.n59 5.04292
R1726 VTAIL.n249 VTAIL.n248 5.04292
R1727 VTAIL.n237 VTAIL.n236 5.04292
R1728 VTAIL.n155 VTAIL.n154 5.04292
R1729 VTAIL.n143 VTAIL.n142 5.04292
R1730 VTAIL.n222 VTAIL.n218 4.38563
R1731 VTAIL.n128 VTAIL.n124 4.38563
R1732 VTAIL.n315 VTAIL.n311 4.38563
R1733 VTAIL.n33 VTAIL.n29 4.38563
R1734 VTAIL.n326 VTAIL.n304 4.26717
R1735 VTAIL.n345 VTAIL.n296 4.26717
R1736 VTAIL.n374 VTAIL.n282 4.26717
R1737 VTAIL.n44 VTAIL.n22 4.26717
R1738 VTAIL.n63 VTAIL.n14 4.26717
R1739 VTAIL.n92 VTAIL.n0 4.26717
R1740 VTAIL.n280 VTAIL.n188 4.26717
R1741 VTAIL.n252 VTAIL.n203 4.26717
R1742 VTAIL.n233 VTAIL.n211 4.26717
R1743 VTAIL.n186 VTAIL.n94 4.26717
R1744 VTAIL.n158 VTAIL.n109 4.26717
R1745 VTAIL.n139 VTAIL.n117 4.26717
R1746 VTAIL.n325 VTAIL.n306 3.49141
R1747 VTAIL.n346 VTAIL.n294 3.49141
R1748 VTAIL.n372 VTAIL.n371 3.49141
R1749 VTAIL.n43 VTAIL.n24 3.49141
R1750 VTAIL.n64 VTAIL.n12 3.49141
R1751 VTAIL.n90 VTAIL.n89 3.49141
R1752 VTAIL.n278 VTAIL.n277 3.49141
R1753 VTAIL.n253 VTAIL.n201 3.49141
R1754 VTAIL.n232 VTAIL.n213 3.49141
R1755 VTAIL.n184 VTAIL.n183 3.49141
R1756 VTAIL.n159 VTAIL.n107 3.49141
R1757 VTAIL.n138 VTAIL.n119 3.49141
R1758 VTAIL.n322 VTAIL.n321 2.71565
R1759 VTAIL.n350 VTAIL.n349 2.71565
R1760 VTAIL.n368 VTAIL.n284 2.71565
R1761 VTAIL.n40 VTAIL.n39 2.71565
R1762 VTAIL.n68 VTAIL.n67 2.71565
R1763 VTAIL.n86 VTAIL.n2 2.71565
R1764 VTAIL.n274 VTAIL.n190 2.71565
R1765 VTAIL.n257 VTAIL.n256 2.71565
R1766 VTAIL.n229 VTAIL.n228 2.71565
R1767 VTAIL.n180 VTAIL.n96 2.71565
R1768 VTAIL.n163 VTAIL.n162 2.71565
R1769 VTAIL.n135 VTAIL.n134 2.71565
R1770 VTAIL.n318 VTAIL.n308 1.93989
R1771 VTAIL.n354 VTAIL.n292 1.93989
R1772 VTAIL.n367 VTAIL.n286 1.93989
R1773 VTAIL.n36 VTAIL.n26 1.93989
R1774 VTAIL.n72 VTAIL.n10 1.93989
R1775 VTAIL.n85 VTAIL.n4 1.93989
R1776 VTAIL.n273 VTAIL.n192 1.93989
R1777 VTAIL.n260 VTAIL.n198 1.93989
R1778 VTAIL.n225 VTAIL.n215 1.93989
R1779 VTAIL.n179 VTAIL.n98 1.93989
R1780 VTAIL.n166 VTAIL.n104 1.93989
R1781 VTAIL.n131 VTAIL.n121 1.93989
R1782 VTAIL.n281 VTAIL.n187 1.17722
R1783 VTAIL.n317 VTAIL.n310 1.16414
R1784 VTAIL.n355 VTAIL.n290 1.16414
R1785 VTAIL.n364 VTAIL.n363 1.16414
R1786 VTAIL.n35 VTAIL.n28 1.16414
R1787 VTAIL.n73 VTAIL.n8 1.16414
R1788 VTAIL.n82 VTAIL.n81 1.16414
R1789 VTAIL.n270 VTAIL.n269 1.16414
R1790 VTAIL.n261 VTAIL.n196 1.16414
R1791 VTAIL.n224 VTAIL.n217 1.16414
R1792 VTAIL.n176 VTAIL.n175 1.16414
R1793 VTAIL.n167 VTAIL.n102 1.16414
R1794 VTAIL.n130 VTAIL.n123 1.16414
R1795 VTAIL VTAIL.n93 0.881965
R1796 VTAIL.n314 VTAIL.n313 0.388379
R1797 VTAIL.n359 VTAIL.n358 0.388379
R1798 VTAIL.n360 VTAIL.n288 0.388379
R1799 VTAIL.n32 VTAIL.n31 0.388379
R1800 VTAIL.n77 VTAIL.n76 0.388379
R1801 VTAIL.n78 VTAIL.n6 0.388379
R1802 VTAIL.n266 VTAIL.n194 0.388379
R1803 VTAIL.n265 VTAIL.n264 0.388379
R1804 VTAIL.n221 VTAIL.n220 0.388379
R1805 VTAIL.n172 VTAIL.n100 0.388379
R1806 VTAIL.n171 VTAIL.n170 0.388379
R1807 VTAIL.n127 VTAIL.n126 0.388379
R1808 VTAIL VTAIL.n375 0.295759
R1809 VTAIL.n316 VTAIL.n315 0.155672
R1810 VTAIL.n316 VTAIL.n307 0.155672
R1811 VTAIL.n323 VTAIL.n307 0.155672
R1812 VTAIL.n324 VTAIL.n323 0.155672
R1813 VTAIL.n324 VTAIL.n303 0.155672
R1814 VTAIL.n331 VTAIL.n303 0.155672
R1815 VTAIL.n332 VTAIL.n331 0.155672
R1816 VTAIL.n332 VTAIL.n299 0.155672
R1817 VTAIL.n339 VTAIL.n299 0.155672
R1818 VTAIL.n340 VTAIL.n339 0.155672
R1819 VTAIL.n340 VTAIL.n295 0.155672
R1820 VTAIL.n347 VTAIL.n295 0.155672
R1821 VTAIL.n348 VTAIL.n347 0.155672
R1822 VTAIL.n348 VTAIL.n291 0.155672
R1823 VTAIL.n356 VTAIL.n291 0.155672
R1824 VTAIL.n357 VTAIL.n356 0.155672
R1825 VTAIL.n357 VTAIL.n287 0.155672
R1826 VTAIL.n365 VTAIL.n287 0.155672
R1827 VTAIL.n366 VTAIL.n365 0.155672
R1828 VTAIL.n366 VTAIL.n283 0.155672
R1829 VTAIL.n373 VTAIL.n283 0.155672
R1830 VTAIL.n34 VTAIL.n33 0.155672
R1831 VTAIL.n34 VTAIL.n25 0.155672
R1832 VTAIL.n41 VTAIL.n25 0.155672
R1833 VTAIL.n42 VTAIL.n41 0.155672
R1834 VTAIL.n42 VTAIL.n21 0.155672
R1835 VTAIL.n49 VTAIL.n21 0.155672
R1836 VTAIL.n50 VTAIL.n49 0.155672
R1837 VTAIL.n50 VTAIL.n17 0.155672
R1838 VTAIL.n57 VTAIL.n17 0.155672
R1839 VTAIL.n58 VTAIL.n57 0.155672
R1840 VTAIL.n58 VTAIL.n13 0.155672
R1841 VTAIL.n65 VTAIL.n13 0.155672
R1842 VTAIL.n66 VTAIL.n65 0.155672
R1843 VTAIL.n66 VTAIL.n9 0.155672
R1844 VTAIL.n74 VTAIL.n9 0.155672
R1845 VTAIL.n75 VTAIL.n74 0.155672
R1846 VTAIL.n75 VTAIL.n5 0.155672
R1847 VTAIL.n83 VTAIL.n5 0.155672
R1848 VTAIL.n84 VTAIL.n83 0.155672
R1849 VTAIL.n84 VTAIL.n1 0.155672
R1850 VTAIL.n91 VTAIL.n1 0.155672
R1851 VTAIL.n279 VTAIL.n189 0.155672
R1852 VTAIL.n272 VTAIL.n189 0.155672
R1853 VTAIL.n272 VTAIL.n271 0.155672
R1854 VTAIL.n271 VTAIL.n193 0.155672
R1855 VTAIL.n263 VTAIL.n193 0.155672
R1856 VTAIL.n263 VTAIL.n262 0.155672
R1857 VTAIL.n262 VTAIL.n197 0.155672
R1858 VTAIL.n255 VTAIL.n197 0.155672
R1859 VTAIL.n255 VTAIL.n254 0.155672
R1860 VTAIL.n254 VTAIL.n202 0.155672
R1861 VTAIL.n247 VTAIL.n202 0.155672
R1862 VTAIL.n247 VTAIL.n246 0.155672
R1863 VTAIL.n246 VTAIL.n206 0.155672
R1864 VTAIL.n239 VTAIL.n206 0.155672
R1865 VTAIL.n239 VTAIL.n238 0.155672
R1866 VTAIL.n238 VTAIL.n210 0.155672
R1867 VTAIL.n231 VTAIL.n210 0.155672
R1868 VTAIL.n231 VTAIL.n230 0.155672
R1869 VTAIL.n230 VTAIL.n214 0.155672
R1870 VTAIL.n223 VTAIL.n214 0.155672
R1871 VTAIL.n223 VTAIL.n222 0.155672
R1872 VTAIL.n185 VTAIL.n95 0.155672
R1873 VTAIL.n178 VTAIL.n95 0.155672
R1874 VTAIL.n178 VTAIL.n177 0.155672
R1875 VTAIL.n177 VTAIL.n99 0.155672
R1876 VTAIL.n169 VTAIL.n99 0.155672
R1877 VTAIL.n169 VTAIL.n168 0.155672
R1878 VTAIL.n168 VTAIL.n103 0.155672
R1879 VTAIL.n161 VTAIL.n103 0.155672
R1880 VTAIL.n161 VTAIL.n160 0.155672
R1881 VTAIL.n160 VTAIL.n108 0.155672
R1882 VTAIL.n153 VTAIL.n108 0.155672
R1883 VTAIL.n153 VTAIL.n152 0.155672
R1884 VTAIL.n152 VTAIL.n112 0.155672
R1885 VTAIL.n145 VTAIL.n112 0.155672
R1886 VTAIL.n145 VTAIL.n144 0.155672
R1887 VTAIL.n144 VTAIL.n116 0.155672
R1888 VTAIL.n137 VTAIL.n116 0.155672
R1889 VTAIL.n137 VTAIL.n136 0.155672
R1890 VTAIL.n136 VTAIL.n120 0.155672
R1891 VTAIL.n129 VTAIL.n120 0.155672
R1892 VTAIL.n129 VTAIL.n128 0.155672
R1893 VDD1.n88 VDD1.n0 289.615
R1894 VDD1.n181 VDD1.n93 289.615
R1895 VDD1.n89 VDD1.n88 185
R1896 VDD1.n87 VDD1.n86 185
R1897 VDD1.n4 VDD1.n3 185
R1898 VDD1.n81 VDD1.n80 185
R1899 VDD1.n79 VDD1.n78 185
R1900 VDD1.n77 VDD1.n7 185
R1901 VDD1.n11 VDD1.n8 185
R1902 VDD1.n72 VDD1.n71 185
R1903 VDD1.n70 VDD1.n69 185
R1904 VDD1.n13 VDD1.n12 185
R1905 VDD1.n64 VDD1.n63 185
R1906 VDD1.n62 VDD1.n61 185
R1907 VDD1.n17 VDD1.n16 185
R1908 VDD1.n56 VDD1.n55 185
R1909 VDD1.n54 VDD1.n53 185
R1910 VDD1.n21 VDD1.n20 185
R1911 VDD1.n48 VDD1.n47 185
R1912 VDD1.n46 VDD1.n45 185
R1913 VDD1.n25 VDD1.n24 185
R1914 VDD1.n40 VDD1.n39 185
R1915 VDD1.n38 VDD1.n37 185
R1916 VDD1.n29 VDD1.n28 185
R1917 VDD1.n32 VDD1.n31 185
R1918 VDD1.n124 VDD1.n123 185
R1919 VDD1.n121 VDD1.n120 185
R1920 VDD1.n130 VDD1.n129 185
R1921 VDD1.n132 VDD1.n131 185
R1922 VDD1.n117 VDD1.n116 185
R1923 VDD1.n138 VDD1.n137 185
R1924 VDD1.n140 VDD1.n139 185
R1925 VDD1.n113 VDD1.n112 185
R1926 VDD1.n146 VDD1.n145 185
R1927 VDD1.n148 VDD1.n147 185
R1928 VDD1.n109 VDD1.n108 185
R1929 VDD1.n154 VDD1.n153 185
R1930 VDD1.n156 VDD1.n155 185
R1931 VDD1.n105 VDD1.n104 185
R1932 VDD1.n162 VDD1.n161 185
R1933 VDD1.n165 VDD1.n164 185
R1934 VDD1.n163 VDD1.n101 185
R1935 VDD1.n170 VDD1.n100 185
R1936 VDD1.n172 VDD1.n171 185
R1937 VDD1.n174 VDD1.n173 185
R1938 VDD1.n97 VDD1.n96 185
R1939 VDD1.n180 VDD1.n179 185
R1940 VDD1.n182 VDD1.n181 185
R1941 VDD1.t0 VDD1.n30 147.659
R1942 VDD1.t1 VDD1.n122 147.659
R1943 VDD1.n88 VDD1.n87 104.615
R1944 VDD1.n87 VDD1.n3 104.615
R1945 VDD1.n80 VDD1.n3 104.615
R1946 VDD1.n80 VDD1.n79 104.615
R1947 VDD1.n79 VDD1.n7 104.615
R1948 VDD1.n11 VDD1.n7 104.615
R1949 VDD1.n71 VDD1.n11 104.615
R1950 VDD1.n71 VDD1.n70 104.615
R1951 VDD1.n70 VDD1.n12 104.615
R1952 VDD1.n63 VDD1.n12 104.615
R1953 VDD1.n63 VDD1.n62 104.615
R1954 VDD1.n62 VDD1.n16 104.615
R1955 VDD1.n55 VDD1.n16 104.615
R1956 VDD1.n55 VDD1.n54 104.615
R1957 VDD1.n54 VDD1.n20 104.615
R1958 VDD1.n47 VDD1.n20 104.615
R1959 VDD1.n47 VDD1.n46 104.615
R1960 VDD1.n46 VDD1.n24 104.615
R1961 VDD1.n39 VDD1.n24 104.615
R1962 VDD1.n39 VDD1.n38 104.615
R1963 VDD1.n38 VDD1.n28 104.615
R1964 VDD1.n31 VDD1.n28 104.615
R1965 VDD1.n123 VDD1.n120 104.615
R1966 VDD1.n130 VDD1.n120 104.615
R1967 VDD1.n131 VDD1.n130 104.615
R1968 VDD1.n131 VDD1.n116 104.615
R1969 VDD1.n138 VDD1.n116 104.615
R1970 VDD1.n139 VDD1.n138 104.615
R1971 VDD1.n139 VDD1.n112 104.615
R1972 VDD1.n146 VDD1.n112 104.615
R1973 VDD1.n147 VDD1.n146 104.615
R1974 VDD1.n147 VDD1.n108 104.615
R1975 VDD1.n154 VDD1.n108 104.615
R1976 VDD1.n155 VDD1.n154 104.615
R1977 VDD1.n155 VDD1.n104 104.615
R1978 VDD1.n162 VDD1.n104 104.615
R1979 VDD1.n164 VDD1.n162 104.615
R1980 VDD1.n164 VDD1.n163 104.615
R1981 VDD1.n163 VDD1.n100 104.615
R1982 VDD1.n172 VDD1.n100 104.615
R1983 VDD1.n173 VDD1.n172 104.615
R1984 VDD1.n173 VDD1.n96 104.615
R1985 VDD1.n180 VDD1.n96 104.615
R1986 VDD1.n181 VDD1.n180 104.615
R1987 VDD1 VDD1.n185 89.6994
R1988 VDD1.n31 VDD1.t0 52.3082
R1989 VDD1.n123 VDD1.t1 52.3082
R1990 VDD1 VDD1.n92 48.3061
R1991 VDD1.n32 VDD1.n30 15.6677
R1992 VDD1.n124 VDD1.n122 15.6677
R1993 VDD1.n78 VDD1.n77 13.1884
R1994 VDD1.n171 VDD1.n170 13.1884
R1995 VDD1.n81 VDD1.n6 12.8005
R1996 VDD1.n76 VDD1.n8 12.8005
R1997 VDD1.n33 VDD1.n29 12.8005
R1998 VDD1.n125 VDD1.n121 12.8005
R1999 VDD1.n169 VDD1.n101 12.8005
R2000 VDD1.n174 VDD1.n99 12.8005
R2001 VDD1.n82 VDD1.n4 12.0247
R2002 VDD1.n73 VDD1.n72 12.0247
R2003 VDD1.n37 VDD1.n36 12.0247
R2004 VDD1.n129 VDD1.n128 12.0247
R2005 VDD1.n166 VDD1.n165 12.0247
R2006 VDD1.n175 VDD1.n97 12.0247
R2007 VDD1.n86 VDD1.n85 11.249
R2008 VDD1.n69 VDD1.n10 11.249
R2009 VDD1.n40 VDD1.n27 11.249
R2010 VDD1.n132 VDD1.n119 11.249
R2011 VDD1.n161 VDD1.n103 11.249
R2012 VDD1.n179 VDD1.n178 11.249
R2013 VDD1.n89 VDD1.n2 10.4732
R2014 VDD1.n68 VDD1.n13 10.4732
R2015 VDD1.n41 VDD1.n25 10.4732
R2016 VDD1.n133 VDD1.n117 10.4732
R2017 VDD1.n160 VDD1.n105 10.4732
R2018 VDD1.n182 VDD1.n95 10.4732
R2019 VDD1.n90 VDD1.n0 9.69747
R2020 VDD1.n65 VDD1.n64 9.69747
R2021 VDD1.n45 VDD1.n44 9.69747
R2022 VDD1.n137 VDD1.n136 9.69747
R2023 VDD1.n157 VDD1.n156 9.69747
R2024 VDD1.n183 VDD1.n93 9.69747
R2025 VDD1.n92 VDD1.n91 9.45567
R2026 VDD1.n185 VDD1.n184 9.45567
R2027 VDD1.n58 VDD1.n57 9.3005
R2028 VDD1.n60 VDD1.n59 9.3005
R2029 VDD1.n15 VDD1.n14 9.3005
R2030 VDD1.n66 VDD1.n65 9.3005
R2031 VDD1.n68 VDD1.n67 9.3005
R2032 VDD1.n10 VDD1.n9 9.3005
R2033 VDD1.n74 VDD1.n73 9.3005
R2034 VDD1.n76 VDD1.n75 9.3005
R2035 VDD1.n91 VDD1.n90 9.3005
R2036 VDD1.n2 VDD1.n1 9.3005
R2037 VDD1.n85 VDD1.n84 9.3005
R2038 VDD1.n83 VDD1.n82 9.3005
R2039 VDD1.n6 VDD1.n5 9.3005
R2040 VDD1.n19 VDD1.n18 9.3005
R2041 VDD1.n52 VDD1.n51 9.3005
R2042 VDD1.n50 VDD1.n49 9.3005
R2043 VDD1.n23 VDD1.n22 9.3005
R2044 VDD1.n44 VDD1.n43 9.3005
R2045 VDD1.n42 VDD1.n41 9.3005
R2046 VDD1.n27 VDD1.n26 9.3005
R2047 VDD1.n36 VDD1.n35 9.3005
R2048 VDD1.n34 VDD1.n33 9.3005
R2049 VDD1.n184 VDD1.n183 9.3005
R2050 VDD1.n95 VDD1.n94 9.3005
R2051 VDD1.n178 VDD1.n177 9.3005
R2052 VDD1.n176 VDD1.n175 9.3005
R2053 VDD1.n99 VDD1.n98 9.3005
R2054 VDD1.n144 VDD1.n143 9.3005
R2055 VDD1.n142 VDD1.n141 9.3005
R2056 VDD1.n115 VDD1.n114 9.3005
R2057 VDD1.n136 VDD1.n135 9.3005
R2058 VDD1.n134 VDD1.n133 9.3005
R2059 VDD1.n119 VDD1.n118 9.3005
R2060 VDD1.n128 VDD1.n127 9.3005
R2061 VDD1.n126 VDD1.n125 9.3005
R2062 VDD1.n111 VDD1.n110 9.3005
R2063 VDD1.n150 VDD1.n149 9.3005
R2064 VDD1.n152 VDD1.n151 9.3005
R2065 VDD1.n107 VDD1.n106 9.3005
R2066 VDD1.n158 VDD1.n157 9.3005
R2067 VDD1.n160 VDD1.n159 9.3005
R2068 VDD1.n103 VDD1.n102 9.3005
R2069 VDD1.n167 VDD1.n166 9.3005
R2070 VDD1.n169 VDD1.n168 9.3005
R2071 VDD1.n61 VDD1.n15 8.92171
R2072 VDD1.n48 VDD1.n23 8.92171
R2073 VDD1.n140 VDD1.n115 8.92171
R2074 VDD1.n153 VDD1.n107 8.92171
R2075 VDD1.n60 VDD1.n17 8.14595
R2076 VDD1.n49 VDD1.n21 8.14595
R2077 VDD1.n141 VDD1.n113 8.14595
R2078 VDD1.n152 VDD1.n109 8.14595
R2079 VDD1.n57 VDD1.n56 7.3702
R2080 VDD1.n53 VDD1.n52 7.3702
R2081 VDD1.n145 VDD1.n144 7.3702
R2082 VDD1.n149 VDD1.n148 7.3702
R2083 VDD1.n56 VDD1.n19 6.59444
R2084 VDD1.n53 VDD1.n19 6.59444
R2085 VDD1.n145 VDD1.n111 6.59444
R2086 VDD1.n148 VDD1.n111 6.59444
R2087 VDD1.n57 VDD1.n17 5.81868
R2088 VDD1.n52 VDD1.n21 5.81868
R2089 VDD1.n144 VDD1.n113 5.81868
R2090 VDD1.n149 VDD1.n109 5.81868
R2091 VDD1.n61 VDD1.n60 5.04292
R2092 VDD1.n49 VDD1.n48 5.04292
R2093 VDD1.n141 VDD1.n140 5.04292
R2094 VDD1.n153 VDD1.n152 5.04292
R2095 VDD1.n34 VDD1.n30 4.38563
R2096 VDD1.n126 VDD1.n122 4.38563
R2097 VDD1.n92 VDD1.n0 4.26717
R2098 VDD1.n64 VDD1.n15 4.26717
R2099 VDD1.n45 VDD1.n23 4.26717
R2100 VDD1.n137 VDD1.n115 4.26717
R2101 VDD1.n156 VDD1.n107 4.26717
R2102 VDD1.n185 VDD1.n93 4.26717
R2103 VDD1.n90 VDD1.n89 3.49141
R2104 VDD1.n65 VDD1.n13 3.49141
R2105 VDD1.n44 VDD1.n25 3.49141
R2106 VDD1.n136 VDD1.n117 3.49141
R2107 VDD1.n157 VDD1.n105 3.49141
R2108 VDD1.n183 VDD1.n182 3.49141
R2109 VDD1.n86 VDD1.n2 2.71565
R2110 VDD1.n69 VDD1.n68 2.71565
R2111 VDD1.n41 VDD1.n40 2.71565
R2112 VDD1.n133 VDD1.n132 2.71565
R2113 VDD1.n161 VDD1.n160 2.71565
R2114 VDD1.n179 VDD1.n95 2.71565
R2115 VDD1.n85 VDD1.n4 1.93989
R2116 VDD1.n72 VDD1.n10 1.93989
R2117 VDD1.n37 VDD1.n27 1.93989
R2118 VDD1.n129 VDD1.n119 1.93989
R2119 VDD1.n165 VDD1.n103 1.93989
R2120 VDD1.n178 VDD1.n97 1.93989
R2121 VDD1.n82 VDD1.n81 1.16414
R2122 VDD1.n73 VDD1.n8 1.16414
R2123 VDD1.n36 VDD1.n29 1.16414
R2124 VDD1.n128 VDD1.n121 1.16414
R2125 VDD1.n166 VDD1.n101 1.16414
R2126 VDD1.n175 VDD1.n174 1.16414
R2127 VDD1.n78 VDD1.n6 0.388379
R2128 VDD1.n77 VDD1.n76 0.388379
R2129 VDD1.n33 VDD1.n32 0.388379
R2130 VDD1.n125 VDD1.n124 0.388379
R2131 VDD1.n170 VDD1.n169 0.388379
R2132 VDD1.n171 VDD1.n99 0.388379
R2133 VDD1.n91 VDD1.n1 0.155672
R2134 VDD1.n84 VDD1.n1 0.155672
R2135 VDD1.n84 VDD1.n83 0.155672
R2136 VDD1.n83 VDD1.n5 0.155672
R2137 VDD1.n75 VDD1.n5 0.155672
R2138 VDD1.n75 VDD1.n74 0.155672
R2139 VDD1.n74 VDD1.n9 0.155672
R2140 VDD1.n67 VDD1.n9 0.155672
R2141 VDD1.n67 VDD1.n66 0.155672
R2142 VDD1.n66 VDD1.n14 0.155672
R2143 VDD1.n59 VDD1.n14 0.155672
R2144 VDD1.n59 VDD1.n58 0.155672
R2145 VDD1.n58 VDD1.n18 0.155672
R2146 VDD1.n51 VDD1.n18 0.155672
R2147 VDD1.n51 VDD1.n50 0.155672
R2148 VDD1.n50 VDD1.n22 0.155672
R2149 VDD1.n43 VDD1.n22 0.155672
R2150 VDD1.n43 VDD1.n42 0.155672
R2151 VDD1.n42 VDD1.n26 0.155672
R2152 VDD1.n35 VDD1.n26 0.155672
R2153 VDD1.n35 VDD1.n34 0.155672
R2154 VDD1.n127 VDD1.n126 0.155672
R2155 VDD1.n127 VDD1.n118 0.155672
R2156 VDD1.n134 VDD1.n118 0.155672
R2157 VDD1.n135 VDD1.n134 0.155672
R2158 VDD1.n135 VDD1.n114 0.155672
R2159 VDD1.n142 VDD1.n114 0.155672
R2160 VDD1.n143 VDD1.n142 0.155672
R2161 VDD1.n143 VDD1.n110 0.155672
R2162 VDD1.n150 VDD1.n110 0.155672
R2163 VDD1.n151 VDD1.n150 0.155672
R2164 VDD1.n151 VDD1.n106 0.155672
R2165 VDD1.n158 VDD1.n106 0.155672
R2166 VDD1.n159 VDD1.n158 0.155672
R2167 VDD1.n159 VDD1.n102 0.155672
R2168 VDD1.n167 VDD1.n102 0.155672
R2169 VDD1.n168 VDD1.n167 0.155672
R2170 VDD1.n168 VDD1.n98 0.155672
R2171 VDD1.n176 VDD1.n98 0.155672
R2172 VDD1.n177 VDD1.n176 0.155672
R2173 VDD1.n177 VDD1.n94 0.155672
R2174 VDD1.n184 VDD1.n94 0.155672
R2175 VN VN.t0 464.043
R2176 VN VN.t1 419.07
R2177 VDD2.n181 VDD2.n93 289.615
R2178 VDD2.n88 VDD2.n0 289.615
R2179 VDD2.n182 VDD2.n181 185
R2180 VDD2.n180 VDD2.n179 185
R2181 VDD2.n97 VDD2.n96 185
R2182 VDD2.n174 VDD2.n173 185
R2183 VDD2.n172 VDD2.n171 185
R2184 VDD2.n170 VDD2.n100 185
R2185 VDD2.n104 VDD2.n101 185
R2186 VDD2.n165 VDD2.n164 185
R2187 VDD2.n163 VDD2.n162 185
R2188 VDD2.n106 VDD2.n105 185
R2189 VDD2.n157 VDD2.n156 185
R2190 VDD2.n155 VDD2.n154 185
R2191 VDD2.n110 VDD2.n109 185
R2192 VDD2.n149 VDD2.n148 185
R2193 VDD2.n147 VDD2.n146 185
R2194 VDD2.n114 VDD2.n113 185
R2195 VDD2.n141 VDD2.n140 185
R2196 VDD2.n139 VDD2.n138 185
R2197 VDD2.n118 VDD2.n117 185
R2198 VDD2.n133 VDD2.n132 185
R2199 VDD2.n131 VDD2.n130 185
R2200 VDD2.n122 VDD2.n121 185
R2201 VDD2.n125 VDD2.n124 185
R2202 VDD2.n31 VDD2.n30 185
R2203 VDD2.n28 VDD2.n27 185
R2204 VDD2.n37 VDD2.n36 185
R2205 VDD2.n39 VDD2.n38 185
R2206 VDD2.n24 VDD2.n23 185
R2207 VDD2.n45 VDD2.n44 185
R2208 VDD2.n47 VDD2.n46 185
R2209 VDD2.n20 VDD2.n19 185
R2210 VDD2.n53 VDD2.n52 185
R2211 VDD2.n55 VDD2.n54 185
R2212 VDD2.n16 VDD2.n15 185
R2213 VDD2.n61 VDD2.n60 185
R2214 VDD2.n63 VDD2.n62 185
R2215 VDD2.n12 VDD2.n11 185
R2216 VDD2.n69 VDD2.n68 185
R2217 VDD2.n72 VDD2.n71 185
R2218 VDD2.n70 VDD2.n8 185
R2219 VDD2.n77 VDD2.n7 185
R2220 VDD2.n79 VDD2.n78 185
R2221 VDD2.n81 VDD2.n80 185
R2222 VDD2.n4 VDD2.n3 185
R2223 VDD2.n87 VDD2.n86 185
R2224 VDD2.n89 VDD2.n88 185
R2225 VDD2.t1 VDD2.n123 147.659
R2226 VDD2.t0 VDD2.n29 147.659
R2227 VDD2.n181 VDD2.n180 104.615
R2228 VDD2.n180 VDD2.n96 104.615
R2229 VDD2.n173 VDD2.n96 104.615
R2230 VDD2.n173 VDD2.n172 104.615
R2231 VDD2.n172 VDD2.n100 104.615
R2232 VDD2.n104 VDD2.n100 104.615
R2233 VDD2.n164 VDD2.n104 104.615
R2234 VDD2.n164 VDD2.n163 104.615
R2235 VDD2.n163 VDD2.n105 104.615
R2236 VDD2.n156 VDD2.n105 104.615
R2237 VDD2.n156 VDD2.n155 104.615
R2238 VDD2.n155 VDD2.n109 104.615
R2239 VDD2.n148 VDD2.n109 104.615
R2240 VDD2.n148 VDD2.n147 104.615
R2241 VDD2.n147 VDD2.n113 104.615
R2242 VDD2.n140 VDD2.n113 104.615
R2243 VDD2.n140 VDD2.n139 104.615
R2244 VDD2.n139 VDD2.n117 104.615
R2245 VDD2.n132 VDD2.n117 104.615
R2246 VDD2.n132 VDD2.n131 104.615
R2247 VDD2.n131 VDD2.n121 104.615
R2248 VDD2.n124 VDD2.n121 104.615
R2249 VDD2.n30 VDD2.n27 104.615
R2250 VDD2.n37 VDD2.n27 104.615
R2251 VDD2.n38 VDD2.n37 104.615
R2252 VDD2.n38 VDD2.n23 104.615
R2253 VDD2.n45 VDD2.n23 104.615
R2254 VDD2.n46 VDD2.n45 104.615
R2255 VDD2.n46 VDD2.n19 104.615
R2256 VDD2.n53 VDD2.n19 104.615
R2257 VDD2.n54 VDD2.n53 104.615
R2258 VDD2.n54 VDD2.n15 104.615
R2259 VDD2.n61 VDD2.n15 104.615
R2260 VDD2.n62 VDD2.n61 104.615
R2261 VDD2.n62 VDD2.n11 104.615
R2262 VDD2.n69 VDD2.n11 104.615
R2263 VDD2.n71 VDD2.n69 104.615
R2264 VDD2.n71 VDD2.n70 104.615
R2265 VDD2.n70 VDD2.n7 104.615
R2266 VDD2.n79 VDD2.n7 104.615
R2267 VDD2.n80 VDD2.n79 104.615
R2268 VDD2.n80 VDD2.n3 104.615
R2269 VDD2.n87 VDD2.n3 104.615
R2270 VDD2.n88 VDD2.n87 104.615
R2271 VDD2.n186 VDD2.n92 88.8211
R2272 VDD2.n124 VDD2.t1 52.3082
R2273 VDD2.n30 VDD2.t0 52.3082
R2274 VDD2.n186 VDD2.n185 47.8944
R2275 VDD2.n125 VDD2.n123 15.6677
R2276 VDD2.n31 VDD2.n29 15.6677
R2277 VDD2.n171 VDD2.n170 13.1884
R2278 VDD2.n78 VDD2.n77 13.1884
R2279 VDD2.n174 VDD2.n99 12.8005
R2280 VDD2.n169 VDD2.n101 12.8005
R2281 VDD2.n126 VDD2.n122 12.8005
R2282 VDD2.n32 VDD2.n28 12.8005
R2283 VDD2.n76 VDD2.n8 12.8005
R2284 VDD2.n81 VDD2.n6 12.8005
R2285 VDD2.n175 VDD2.n97 12.0247
R2286 VDD2.n166 VDD2.n165 12.0247
R2287 VDD2.n130 VDD2.n129 12.0247
R2288 VDD2.n36 VDD2.n35 12.0247
R2289 VDD2.n73 VDD2.n72 12.0247
R2290 VDD2.n82 VDD2.n4 12.0247
R2291 VDD2.n179 VDD2.n178 11.249
R2292 VDD2.n162 VDD2.n103 11.249
R2293 VDD2.n133 VDD2.n120 11.249
R2294 VDD2.n39 VDD2.n26 11.249
R2295 VDD2.n68 VDD2.n10 11.249
R2296 VDD2.n86 VDD2.n85 11.249
R2297 VDD2.n182 VDD2.n95 10.4732
R2298 VDD2.n161 VDD2.n106 10.4732
R2299 VDD2.n134 VDD2.n118 10.4732
R2300 VDD2.n40 VDD2.n24 10.4732
R2301 VDD2.n67 VDD2.n12 10.4732
R2302 VDD2.n89 VDD2.n2 10.4732
R2303 VDD2.n183 VDD2.n93 9.69747
R2304 VDD2.n158 VDD2.n157 9.69747
R2305 VDD2.n138 VDD2.n137 9.69747
R2306 VDD2.n44 VDD2.n43 9.69747
R2307 VDD2.n64 VDD2.n63 9.69747
R2308 VDD2.n90 VDD2.n0 9.69747
R2309 VDD2.n185 VDD2.n184 9.45567
R2310 VDD2.n92 VDD2.n91 9.45567
R2311 VDD2.n151 VDD2.n150 9.3005
R2312 VDD2.n153 VDD2.n152 9.3005
R2313 VDD2.n108 VDD2.n107 9.3005
R2314 VDD2.n159 VDD2.n158 9.3005
R2315 VDD2.n161 VDD2.n160 9.3005
R2316 VDD2.n103 VDD2.n102 9.3005
R2317 VDD2.n167 VDD2.n166 9.3005
R2318 VDD2.n169 VDD2.n168 9.3005
R2319 VDD2.n184 VDD2.n183 9.3005
R2320 VDD2.n95 VDD2.n94 9.3005
R2321 VDD2.n178 VDD2.n177 9.3005
R2322 VDD2.n176 VDD2.n175 9.3005
R2323 VDD2.n99 VDD2.n98 9.3005
R2324 VDD2.n112 VDD2.n111 9.3005
R2325 VDD2.n145 VDD2.n144 9.3005
R2326 VDD2.n143 VDD2.n142 9.3005
R2327 VDD2.n116 VDD2.n115 9.3005
R2328 VDD2.n137 VDD2.n136 9.3005
R2329 VDD2.n135 VDD2.n134 9.3005
R2330 VDD2.n120 VDD2.n119 9.3005
R2331 VDD2.n129 VDD2.n128 9.3005
R2332 VDD2.n127 VDD2.n126 9.3005
R2333 VDD2.n91 VDD2.n90 9.3005
R2334 VDD2.n2 VDD2.n1 9.3005
R2335 VDD2.n85 VDD2.n84 9.3005
R2336 VDD2.n83 VDD2.n82 9.3005
R2337 VDD2.n6 VDD2.n5 9.3005
R2338 VDD2.n51 VDD2.n50 9.3005
R2339 VDD2.n49 VDD2.n48 9.3005
R2340 VDD2.n22 VDD2.n21 9.3005
R2341 VDD2.n43 VDD2.n42 9.3005
R2342 VDD2.n41 VDD2.n40 9.3005
R2343 VDD2.n26 VDD2.n25 9.3005
R2344 VDD2.n35 VDD2.n34 9.3005
R2345 VDD2.n33 VDD2.n32 9.3005
R2346 VDD2.n18 VDD2.n17 9.3005
R2347 VDD2.n57 VDD2.n56 9.3005
R2348 VDD2.n59 VDD2.n58 9.3005
R2349 VDD2.n14 VDD2.n13 9.3005
R2350 VDD2.n65 VDD2.n64 9.3005
R2351 VDD2.n67 VDD2.n66 9.3005
R2352 VDD2.n10 VDD2.n9 9.3005
R2353 VDD2.n74 VDD2.n73 9.3005
R2354 VDD2.n76 VDD2.n75 9.3005
R2355 VDD2.n154 VDD2.n108 8.92171
R2356 VDD2.n141 VDD2.n116 8.92171
R2357 VDD2.n47 VDD2.n22 8.92171
R2358 VDD2.n60 VDD2.n14 8.92171
R2359 VDD2.n153 VDD2.n110 8.14595
R2360 VDD2.n142 VDD2.n114 8.14595
R2361 VDD2.n48 VDD2.n20 8.14595
R2362 VDD2.n59 VDD2.n16 8.14595
R2363 VDD2.n150 VDD2.n149 7.3702
R2364 VDD2.n146 VDD2.n145 7.3702
R2365 VDD2.n52 VDD2.n51 7.3702
R2366 VDD2.n56 VDD2.n55 7.3702
R2367 VDD2.n149 VDD2.n112 6.59444
R2368 VDD2.n146 VDD2.n112 6.59444
R2369 VDD2.n52 VDD2.n18 6.59444
R2370 VDD2.n55 VDD2.n18 6.59444
R2371 VDD2.n150 VDD2.n110 5.81868
R2372 VDD2.n145 VDD2.n114 5.81868
R2373 VDD2.n51 VDD2.n20 5.81868
R2374 VDD2.n56 VDD2.n16 5.81868
R2375 VDD2.n154 VDD2.n153 5.04292
R2376 VDD2.n142 VDD2.n141 5.04292
R2377 VDD2.n48 VDD2.n47 5.04292
R2378 VDD2.n60 VDD2.n59 5.04292
R2379 VDD2.n127 VDD2.n123 4.38563
R2380 VDD2.n33 VDD2.n29 4.38563
R2381 VDD2.n185 VDD2.n93 4.26717
R2382 VDD2.n157 VDD2.n108 4.26717
R2383 VDD2.n138 VDD2.n116 4.26717
R2384 VDD2.n44 VDD2.n22 4.26717
R2385 VDD2.n63 VDD2.n14 4.26717
R2386 VDD2.n92 VDD2.n0 4.26717
R2387 VDD2.n183 VDD2.n182 3.49141
R2388 VDD2.n158 VDD2.n106 3.49141
R2389 VDD2.n137 VDD2.n118 3.49141
R2390 VDD2.n43 VDD2.n24 3.49141
R2391 VDD2.n64 VDD2.n12 3.49141
R2392 VDD2.n90 VDD2.n89 3.49141
R2393 VDD2.n179 VDD2.n95 2.71565
R2394 VDD2.n162 VDD2.n161 2.71565
R2395 VDD2.n134 VDD2.n133 2.71565
R2396 VDD2.n40 VDD2.n39 2.71565
R2397 VDD2.n68 VDD2.n67 2.71565
R2398 VDD2.n86 VDD2.n2 2.71565
R2399 VDD2.n178 VDD2.n97 1.93989
R2400 VDD2.n165 VDD2.n103 1.93989
R2401 VDD2.n130 VDD2.n120 1.93989
R2402 VDD2.n36 VDD2.n26 1.93989
R2403 VDD2.n72 VDD2.n10 1.93989
R2404 VDD2.n85 VDD2.n4 1.93989
R2405 VDD2.n175 VDD2.n174 1.16414
R2406 VDD2.n166 VDD2.n101 1.16414
R2407 VDD2.n129 VDD2.n122 1.16414
R2408 VDD2.n35 VDD2.n28 1.16414
R2409 VDD2.n73 VDD2.n8 1.16414
R2410 VDD2.n82 VDD2.n81 1.16414
R2411 VDD2 VDD2.n186 0.412138
R2412 VDD2.n171 VDD2.n99 0.388379
R2413 VDD2.n170 VDD2.n169 0.388379
R2414 VDD2.n126 VDD2.n125 0.388379
R2415 VDD2.n32 VDD2.n31 0.388379
R2416 VDD2.n77 VDD2.n76 0.388379
R2417 VDD2.n78 VDD2.n6 0.388379
R2418 VDD2.n184 VDD2.n94 0.155672
R2419 VDD2.n177 VDD2.n94 0.155672
R2420 VDD2.n177 VDD2.n176 0.155672
R2421 VDD2.n176 VDD2.n98 0.155672
R2422 VDD2.n168 VDD2.n98 0.155672
R2423 VDD2.n168 VDD2.n167 0.155672
R2424 VDD2.n167 VDD2.n102 0.155672
R2425 VDD2.n160 VDD2.n102 0.155672
R2426 VDD2.n160 VDD2.n159 0.155672
R2427 VDD2.n159 VDD2.n107 0.155672
R2428 VDD2.n152 VDD2.n107 0.155672
R2429 VDD2.n152 VDD2.n151 0.155672
R2430 VDD2.n151 VDD2.n111 0.155672
R2431 VDD2.n144 VDD2.n111 0.155672
R2432 VDD2.n144 VDD2.n143 0.155672
R2433 VDD2.n143 VDD2.n115 0.155672
R2434 VDD2.n136 VDD2.n115 0.155672
R2435 VDD2.n136 VDD2.n135 0.155672
R2436 VDD2.n135 VDD2.n119 0.155672
R2437 VDD2.n128 VDD2.n119 0.155672
R2438 VDD2.n128 VDD2.n127 0.155672
R2439 VDD2.n34 VDD2.n33 0.155672
R2440 VDD2.n34 VDD2.n25 0.155672
R2441 VDD2.n41 VDD2.n25 0.155672
R2442 VDD2.n42 VDD2.n41 0.155672
R2443 VDD2.n42 VDD2.n21 0.155672
R2444 VDD2.n49 VDD2.n21 0.155672
R2445 VDD2.n50 VDD2.n49 0.155672
R2446 VDD2.n50 VDD2.n17 0.155672
R2447 VDD2.n57 VDD2.n17 0.155672
R2448 VDD2.n58 VDD2.n57 0.155672
R2449 VDD2.n58 VDD2.n13 0.155672
R2450 VDD2.n65 VDD2.n13 0.155672
R2451 VDD2.n66 VDD2.n65 0.155672
R2452 VDD2.n66 VDD2.n9 0.155672
R2453 VDD2.n74 VDD2.n9 0.155672
R2454 VDD2.n75 VDD2.n74 0.155672
R2455 VDD2.n75 VDD2.n5 0.155672
R2456 VDD2.n83 VDD2.n5 0.155672
R2457 VDD2.n84 VDD2.n83 0.155672
R2458 VDD2.n84 VDD2.n1 0.155672
R2459 VDD2.n91 VDD2.n1 0.155672
C0 VDD1 VTAIL 6.58222f
C1 VDD2 VTAIL 6.62015f
C2 VDD1 VN 0.147531f
C3 VDD2 VN 3.27622f
C4 VDD1 VP 3.40352f
C5 VDD2 VP 0.279631f
C6 VN VTAIL 2.64923f
C7 VDD1 VDD2 0.52614f
C8 VTAIL VP 2.66382f
C9 VN VP 5.73044f
C10 VDD2 B 4.830771f
C11 VDD1 B 7.66905f
C12 VTAIL B 8.515133f
C13 VN B 10.69649f
C14 VP B 5.112882f
C15 VDD2.n0 B 0.026518f
C16 VDD2.n1 B 0.020122f
C17 VDD2.n2 B 0.010813f
C18 VDD2.n3 B 0.025557f
C19 VDD2.n4 B 0.011449f
C20 VDD2.n5 B 0.020122f
C21 VDD2.n6 B 0.010813f
C22 VDD2.n7 B 0.025557f
C23 VDD2.n8 B 0.011449f
C24 VDD2.n9 B 0.020122f
C25 VDD2.n10 B 0.010813f
C26 VDD2.n11 B 0.025557f
C27 VDD2.n12 B 0.011449f
C28 VDD2.n13 B 0.020122f
C29 VDD2.n14 B 0.010813f
C30 VDD2.n15 B 0.025557f
C31 VDD2.n16 B 0.011449f
C32 VDD2.n17 B 0.020122f
C33 VDD2.n18 B 0.010813f
C34 VDD2.n19 B 0.025557f
C35 VDD2.n20 B 0.011449f
C36 VDD2.n21 B 0.020122f
C37 VDD2.n22 B 0.010813f
C38 VDD2.n23 B 0.025557f
C39 VDD2.n24 B 0.011449f
C40 VDD2.n25 B 0.020122f
C41 VDD2.n26 B 0.010813f
C42 VDD2.n27 B 0.025557f
C43 VDD2.n28 B 0.011449f
C44 VDD2.n29 B 0.140068f
C45 VDD2.t0 B 0.042261f
C46 VDD2.n30 B 0.019168f
C47 VDD2.n31 B 0.015097f
C48 VDD2.n32 B 0.010813f
C49 VDD2.n33 B 1.47054f
C50 VDD2.n34 B 0.020122f
C51 VDD2.n35 B 0.010813f
C52 VDD2.n36 B 0.011449f
C53 VDD2.n37 B 0.025557f
C54 VDD2.n38 B 0.025557f
C55 VDD2.n39 B 0.011449f
C56 VDD2.n40 B 0.010813f
C57 VDD2.n41 B 0.020122f
C58 VDD2.n42 B 0.020122f
C59 VDD2.n43 B 0.010813f
C60 VDD2.n44 B 0.011449f
C61 VDD2.n45 B 0.025557f
C62 VDD2.n46 B 0.025557f
C63 VDD2.n47 B 0.011449f
C64 VDD2.n48 B 0.010813f
C65 VDD2.n49 B 0.020122f
C66 VDD2.n50 B 0.020122f
C67 VDD2.n51 B 0.010813f
C68 VDD2.n52 B 0.011449f
C69 VDD2.n53 B 0.025557f
C70 VDD2.n54 B 0.025557f
C71 VDD2.n55 B 0.011449f
C72 VDD2.n56 B 0.010813f
C73 VDD2.n57 B 0.020122f
C74 VDD2.n58 B 0.020122f
C75 VDD2.n59 B 0.010813f
C76 VDD2.n60 B 0.011449f
C77 VDD2.n61 B 0.025557f
C78 VDD2.n62 B 0.025557f
C79 VDD2.n63 B 0.011449f
C80 VDD2.n64 B 0.010813f
C81 VDD2.n65 B 0.020122f
C82 VDD2.n66 B 0.020122f
C83 VDD2.n67 B 0.010813f
C84 VDD2.n68 B 0.011449f
C85 VDD2.n69 B 0.025557f
C86 VDD2.n70 B 0.025557f
C87 VDD2.n71 B 0.025557f
C88 VDD2.n72 B 0.011449f
C89 VDD2.n73 B 0.010813f
C90 VDD2.n74 B 0.020122f
C91 VDD2.n75 B 0.020122f
C92 VDD2.n76 B 0.010813f
C93 VDD2.n77 B 0.011131f
C94 VDD2.n78 B 0.011131f
C95 VDD2.n79 B 0.025557f
C96 VDD2.n80 B 0.025557f
C97 VDD2.n81 B 0.011449f
C98 VDD2.n82 B 0.010813f
C99 VDD2.n83 B 0.020122f
C100 VDD2.n84 B 0.020122f
C101 VDD2.n85 B 0.010813f
C102 VDD2.n86 B 0.011449f
C103 VDD2.n87 B 0.025557f
C104 VDD2.n88 B 0.052206f
C105 VDD2.n89 B 0.011449f
C106 VDD2.n90 B 0.010813f
C107 VDD2.n91 B 0.045136f
C108 VDD2.n92 B 0.665351f
C109 VDD2.n93 B 0.026518f
C110 VDD2.n94 B 0.020122f
C111 VDD2.n95 B 0.010813f
C112 VDD2.n96 B 0.025557f
C113 VDD2.n97 B 0.011449f
C114 VDD2.n98 B 0.020122f
C115 VDD2.n99 B 0.010813f
C116 VDD2.n100 B 0.025557f
C117 VDD2.n101 B 0.011449f
C118 VDD2.n102 B 0.020122f
C119 VDD2.n103 B 0.010813f
C120 VDD2.n104 B 0.025557f
C121 VDD2.n105 B 0.025557f
C122 VDD2.n106 B 0.011449f
C123 VDD2.n107 B 0.020122f
C124 VDD2.n108 B 0.010813f
C125 VDD2.n109 B 0.025557f
C126 VDD2.n110 B 0.011449f
C127 VDD2.n111 B 0.020122f
C128 VDD2.n112 B 0.010813f
C129 VDD2.n113 B 0.025557f
C130 VDD2.n114 B 0.011449f
C131 VDD2.n115 B 0.020122f
C132 VDD2.n116 B 0.010813f
C133 VDD2.n117 B 0.025557f
C134 VDD2.n118 B 0.011449f
C135 VDD2.n119 B 0.020122f
C136 VDD2.n120 B 0.010813f
C137 VDD2.n121 B 0.025557f
C138 VDD2.n122 B 0.011449f
C139 VDD2.n123 B 0.140068f
C140 VDD2.t1 B 0.042261f
C141 VDD2.n124 B 0.019168f
C142 VDD2.n125 B 0.015097f
C143 VDD2.n126 B 0.010813f
C144 VDD2.n127 B 1.47054f
C145 VDD2.n128 B 0.020122f
C146 VDD2.n129 B 0.010813f
C147 VDD2.n130 B 0.011449f
C148 VDD2.n131 B 0.025557f
C149 VDD2.n132 B 0.025557f
C150 VDD2.n133 B 0.011449f
C151 VDD2.n134 B 0.010813f
C152 VDD2.n135 B 0.020122f
C153 VDD2.n136 B 0.020122f
C154 VDD2.n137 B 0.010813f
C155 VDD2.n138 B 0.011449f
C156 VDD2.n139 B 0.025557f
C157 VDD2.n140 B 0.025557f
C158 VDD2.n141 B 0.011449f
C159 VDD2.n142 B 0.010813f
C160 VDD2.n143 B 0.020122f
C161 VDD2.n144 B 0.020122f
C162 VDD2.n145 B 0.010813f
C163 VDD2.n146 B 0.011449f
C164 VDD2.n147 B 0.025557f
C165 VDD2.n148 B 0.025557f
C166 VDD2.n149 B 0.011449f
C167 VDD2.n150 B 0.010813f
C168 VDD2.n151 B 0.020122f
C169 VDD2.n152 B 0.020122f
C170 VDD2.n153 B 0.010813f
C171 VDD2.n154 B 0.011449f
C172 VDD2.n155 B 0.025557f
C173 VDD2.n156 B 0.025557f
C174 VDD2.n157 B 0.011449f
C175 VDD2.n158 B 0.010813f
C176 VDD2.n159 B 0.020122f
C177 VDD2.n160 B 0.020122f
C178 VDD2.n161 B 0.010813f
C179 VDD2.n162 B 0.011449f
C180 VDD2.n163 B 0.025557f
C181 VDD2.n164 B 0.025557f
C182 VDD2.n165 B 0.011449f
C183 VDD2.n166 B 0.010813f
C184 VDD2.n167 B 0.020122f
C185 VDD2.n168 B 0.020122f
C186 VDD2.n169 B 0.010813f
C187 VDD2.n170 B 0.011131f
C188 VDD2.n171 B 0.011131f
C189 VDD2.n172 B 0.025557f
C190 VDD2.n173 B 0.025557f
C191 VDD2.n174 B 0.011449f
C192 VDD2.n175 B 0.010813f
C193 VDD2.n176 B 0.020122f
C194 VDD2.n177 B 0.020122f
C195 VDD2.n178 B 0.010813f
C196 VDD2.n179 B 0.011449f
C197 VDD2.n180 B 0.025557f
C198 VDD2.n181 B 0.052206f
C199 VDD2.n182 B 0.011449f
C200 VDD2.n183 B 0.010813f
C201 VDD2.n184 B 0.045136f
C202 VDD2.n185 B 0.042752f
C203 VDD2.n186 B 2.64034f
C204 VN.t1 B 2.90037f
C205 VN.t0 B 3.17971f
C206 VDD1.n0 B 0.026586f
C207 VDD1.n1 B 0.020174f
C208 VDD1.n2 B 0.01084f
C209 VDD1.n3 B 0.025623f
C210 VDD1.n4 B 0.011478f
C211 VDD1.n5 B 0.020174f
C212 VDD1.n6 B 0.01084f
C213 VDD1.n7 B 0.025623f
C214 VDD1.n8 B 0.011478f
C215 VDD1.n9 B 0.020174f
C216 VDD1.n10 B 0.01084f
C217 VDD1.n11 B 0.025623f
C218 VDD1.n12 B 0.025623f
C219 VDD1.n13 B 0.011478f
C220 VDD1.n14 B 0.020174f
C221 VDD1.n15 B 0.01084f
C222 VDD1.n16 B 0.025623f
C223 VDD1.n17 B 0.011478f
C224 VDD1.n18 B 0.020174f
C225 VDD1.n19 B 0.01084f
C226 VDD1.n20 B 0.025623f
C227 VDD1.n21 B 0.011478f
C228 VDD1.n22 B 0.020174f
C229 VDD1.n23 B 0.01084f
C230 VDD1.n24 B 0.025623f
C231 VDD1.n25 B 0.011478f
C232 VDD1.n26 B 0.020174f
C233 VDD1.n27 B 0.01084f
C234 VDD1.n28 B 0.025623f
C235 VDD1.n29 B 0.011478f
C236 VDD1.n30 B 0.140428f
C237 VDD1.t0 B 0.04237f
C238 VDD1.n31 B 0.019217f
C239 VDD1.n32 B 0.015136f
C240 VDD1.n33 B 0.01084f
C241 VDD1.n34 B 1.47432f
C242 VDD1.n35 B 0.020174f
C243 VDD1.n36 B 0.01084f
C244 VDD1.n37 B 0.011478f
C245 VDD1.n38 B 0.025623f
C246 VDD1.n39 B 0.025623f
C247 VDD1.n40 B 0.011478f
C248 VDD1.n41 B 0.01084f
C249 VDD1.n42 B 0.020174f
C250 VDD1.n43 B 0.020174f
C251 VDD1.n44 B 0.01084f
C252 VDD1.n45 B 0.011478f
C253 VDD1.n46 B 0.025623f
C254 VDD1.n47 B 0.025623f
C255 VDD1.n48 B 0.011478f
C256 VDD1.n49 B 0.01084f
C257 VDD1.n50 B 0.020174f
C258 VDD1.n51 B 0.020174f
C259 VDD1.n52 B 0.01084f
C260 VDD1.n53 B 0.011478f
C261 VDD1.n54 B 0.025623f
C262 VDD1.n55 B 0.025623f
C263 VDD1.n56 B 0.011478f
C264 VDD1.n57 B 0.01084f
C265 VDD1.n58 B 0.020174f
C266 VDD1.n59 B 0.020174f
C267 VDD1.n60 B 0.01084f
C268 VDD1.n61 B 0.011478f
C269 VDD1.n62 B 0.025623f
C270 VDD1.n63 B 0.025623f
C271 VDD1.n64 B 0.011478f
C272 VDD1.n65 B 0.01084f
C273 VDD1.n66 B 0.020174f
C274 VDD1.n67 B 0.020174f
C275 VDD1.n68 B 0.01084f
C276 VDD1.n69 B 0.011478f
C277 VDD1.n70 B 0.025623f
C278 VDD1.n71 B 0.025623f
C279 VDD1.n72 B 0.011478f
C280 VDD1.n73 B 0.01084f
C281 VDD1.n74 B 0.020174f
C282 VDD1.n75 B 0.020174f
C283 VDD1.n76 B 0.01084f
C284 VDD1.n77 B 0.011159f
C285 VDD1.n78 B 0.011159f
C286 VDD1.n79 B 0.025623f
C287 VDD1.n80 B 0.025623f
C288 VDD1.n81 B 0.011478f
C289 VDD1.n82 B 0.01084f
C290 VDD1.n83 B 0.020174f
C291 VDD1.n84 B 0.020174f
C292 VDD1.n85 B 0.01084f
C293 VDD1.n86 B 0.011478f
C294 VDD1.n87 B 0.025623f
C295 VDD1.n88 B 0.05234f
C296 VDD1.n89 B 0.011478f
C297 VDD1.n90 B 0.01084f
C298 VDD1.n91 B 0.045252f
C299 VDD1.n92 B 0.043415f
C300 VDD1.n93 B 0.026586f
C301 VDD1.n94 B 0.020174f
C302 VDD1.n95 B 0.01084f
C303 VDD1.n96 B 0.025623f
C304 VDD1.n97 B 0.011478f
C305 VDD1.n98 B 0.020174f
C306 VDD1.n99 B 0.01084f
C307 VDD1.n100 B 0.025623f
C308 VDD1.n101 B 0.011478f
C309 VDD1.n102 B 0.020174f
C310 VDD1.n103 B 0.01084f
C311 VDD1.n104 B 0.025623f
C312 VDD1.n105 B 0.011478f
C313 VDD1.n106 B 0.020174f
C314 VDD1.n107 B 0.01084f
C315 VDD1.n108 B 0.025623f
C316 VDD1.n109 B 0.011478f
C317 VDD1.n110 B 0.020174f
C318 VDD1.n111 B 0.01084f
C319 VDD1.n112 B 0.025623f
C320 VDD1.n113 B 0.011478f
C321 VDD1.n114 B 0.020174f
C322 VDD1.n115 B 0.01084f
C323 VDD1.n116 B 0.025623f
C324 VDD1.n117 B 0.011478f
C325 VDD1.n118 B 0.020174f
C326 VDD1.n119 B 0.01084f
C327 VDD1.n120 B 0.025623f
C328 VDD1.n121 B 0.011478f
C329 VDD1.n122 B 0.140428f
C330 VDD1.t1 B 0.04237f
C331 VDD1.n123 B 0.019217f
C332 VDD1.n124 B 0.015136f
C333 VDD1.n125 B 0.01084f
C334 VDD1.n126 B 1.47432f
C335 VDD1.n127 B 0.020174f
C336 VDD1.n128 B 0.01084f
C337 VDD1.n129 B 0.011478f
C338 VDD1.n130 B 0.025623f
C339 VDD1.n131 B 0.025623f
C340 VDD1.n132 B 0.011478f
C341 VDD1.n133 B 0.01084f
C342 VDD1.n134 B 0.020174f
C343 VDD1.n135 B 0.020174f
C344 VDD1.n136 B 0.01084f
C345 VDD1.n137 B 0.011478f
C346 VDD1.n138 B 0.025623f
C347 VDD1.n139 B 0.025623f
C348 VDD1.n140 B 0.011478f
C349 VDD1.n141 B 0.01084f
C350 VDD1.n142 B 0.020174f
C351 VDD1.n143 B 0.020174f
C352 VDD1.n144 B 0.01084f
C353 VDD1.n145 B 0.011478f
C354 VDD1.n146 B 0.025623f
C355 VDD1.n147 B 0.025623f
C356 VDD1.n148 B 0.011478f
C357 VDD1.n149 B 0.01084f
C358 VDD1.n150 B 0.020174f
C359 VDD1.n151 B 0.020174f
C360 VDD1.n152 B 0.01084f
C361 VDD1.n153 B 0.011478f
C362 VDD1.n154 B 0.025623f
C363 VDD1.n155 B 0.025623f
C364 VDD1.n156 B 0.011478f
C365 VDD1.n157 B 0.01084f
C366 VDD1.n158 B 0.020174f
C367 VDD1.n159 B 0.020174f
C368 VDD1.n160 B 0.01084f
C369 VDD1.n161 B 0.011478f
C370 VDD1.n162 B 0.025623f
C371 VDD1.n163 B 0.025623f
C372 VDD1.n164 B 0.025623f
C373 VDD1.n165 B 0.011478f
C374 VDD1.n166 B 0.01084f
C375 VDD1.n167 B 0.020174f
C376 VDD1.n168 B 0.020174f
C377 VDD1.n169 B 0.01084f
C378 VDD1.n170 B 0.011159f
C379 VDD1.n171 B 0.011159f
C380 VDD1.n172 B 0.025623f
C381 VDD1.n173 B 0.025623f
C382 VDD1.n174 B 0.011478f
C383 VDD1.n175 B 0.01084f
C384 VDD1.n176 B 0.020174f
C385 VDD1.n177 B 0.020174f
C386 VDD1.n178 B 0.01084f
C387 VDD1.n179 B 0.011478f
C388 VDD1.n180 B 0.025623f
C389 VDD1.n181 B 0.05234f
C390 VDD1.n182 B 0.011478f
C391 VDD1.n183 B 0.01084f
C392 VDD1.n184 B 0.045252f
C393 VDD1.n185 B 0.700523f
C394 VTAIL.n0 B 0.026052f
C395 VTAIL.n1 B 0.019768f
C396 VTAIL.n2 B 0.010622f
C397 VTAIL.n3 B 0.025107f
C398 VTAIL.n4 B 0.011247f
C399 VTAIL.n5 B 0.019768f
C400 VTAIL.n6 B 0.010622f
C401 VTAIL.n7 B 0.025107f
C402 VTAIL.n8 B 0.011247f
C403 VTAIL.n9 B 0.019768f
C404 VTAIL.n10 B 0.010622f
C405 VTAIL.n11 B 0.025107f
C406 VTAIL.n12 B 0.011247f
C407 VTAIL.n13 B 0.019768f
C408 VTAIL.n14 B 0.010622f
C409 VTAIL.n15 B 0.025107f
C410 VTAIL.n16 B 0.011247f
C411 VTAIL.n17 B 0.019768f
C412 VTAIL.n18 B 0.010622f
C413 VTAIL.n19 B 0.025107f
C414 VTAIL.n20 B 0.011247f
C415 VTAIL.n21 B 0.019768f
C416 VTAIL.n22 B 0.010622f
C417 VTAIL.n23 B 0.025107f
C418 VTAIL.n24 B 0.011247f
C419 VTAIL.n25 B 0.019768f
C420 VTAIL.n26 B 0.010622f
C421 VTAIL.n27 B 0.025107f
C422 VTAIL.n28 B 0.011247f
C423 VTAIL.n29 B 0.137603f
C424 VTAIL.t3 B 0.041518f
C425 VTAIL.n30 B 0.018831f
C426 VTAIL.n31 B 0.014832f
C427 VTAIL.n32 B 0.010622f
C428 VTAIL.n33 B 1.44466f
C429 VTAIL.n34 B 0.019768f
C430 VTAIL.n35 B 0.010622f
C431 VTAIL.n36 B 0.011247f
C432 VTAIL.n37 B 0.025107f
C433 VTAIL.n38 B 0.025107f
C434 VTAIL.n39 B 0.011247f
C435 VTAIL.n40 B 0.010622f
C436 VTAIL.n41 B 0.019768f
C437 VTAIL.n42 B 0.019768f
C438 VTAIL.n43 B 0.010622f
C439 VTAIL.n44 B 0.011247f
C440 VTAIL.n45 B 0.025107f
C441 VTAIL.n46 B 0.025107f
C442 VTAIL.n47 B 0.011247f
C443 VTAIL.n48 B 0.010622f
C444 VTAIL.n49 B 0.019768f
C445 VTAIL.n50 B 0.019768f
C446 VTAIL.n51 B 0.010622f
C447 VTAIL.n52 B 0.011247f
C448 VTAIL.n53 B 0.025107f
C449 VTAIL.n54 B 0.025107f
C450 VTAIL.n55 B 0.011247f
C451 VTAIL.n56 B 0.010622f
C452 VTAIL.n57 B 0.019768f
C453 VTAIL.n58 B 0.019768f
C454 VTAIL.n59 B 0.010622f
C455 VTAIL.n60 B 0.011247f
C456 VTAIL.n61 B 0.025107f
C457 VTAIL.n62 B 0.025107f
C458 VTAIL.n63 B 0.011247f
C459 VTAIL.n64 B 0.010622f
C460 VTAIL.n65 B 0.019768f
C461 VTAIL.n66 B 0.019768f
C462 VTAIL.n67 B 0.010622f
C463 VTAIL.n68 B 0.011247f
C464 VTAIL.n69 B 0.025107f
C465 VTAIL.n70 B 0.025107f
C466 VTAIL.n71 B 0.025107f
C467 VTAIL.n72 B 0.011247f
C468 VTAIL.n73 B 0.010622f
C469 VTAIL.n74 B 0.019768f
C470 VTAIL.n75 B 0.019768f
C471 VTAIL.n76 B 0.010622f
C472 VTAIL.n77 B 0.010935f
C473 VTAIL.n78 B 0.010935f
C474 VTAIL.n79 B 0.025107f
C475 VTAIL.n80 B 0.025107f
C476 VTAIL.n81 B 0.011247f
C477 VTAIL.n82 B 0.010622f
C478 VTAIL.n83 B 0.019768f
C479 VTAIL.n84 B 0.019768f
C480 VTAIL.n85 B 0.010622f
C481 VTAIL.n86 B 0.011247f
C482 VTAIL.n87 B 0.025107f
C483 VTAIL.n88 B 0.051287f
C484 VTAIL.n89 B 0.011247f
C485 VTAIL.n90 B 0.010622f
C486 VTAIL.n91 B 0.044342f
C487 VTAIL.n92 B 0.02834f
C488 VTAIL.n93 B 1.44064f
C489 VTAIL.n94 B 0.026052f
C490 VTAIL.n95 B 0.019768f
C491 VTAIL.n96 B 0.010622f
C492 VTAIL.n97 B 0.025107f
C493 VTAIL.n98 B 0.011247f
C494 VTAIL.n99 B 0.019768f
C495 VTAIL.n100 B 0.010622f
C496 VTAIL.n101 B 0.025107f
C497 VTAIL.n102 B 0.011247f
C498 VTAIL.n103 B 0.019768f
C499 VTAIL.n104 B 0.010622f
C500 VTAIL.n105 B 0.025107f
C501 VTAIL.n106 B 0.025107f
C502 VTAIL.n107 B 0.011247f
C503 VTAIL.n108 B 0.019768f
C504 VTAIL.n109 B 0.010622f
C505 VTAIL.n110 B 0.025107f
C506 VTAIL.n111 B 0.011247f
C507 VTAIL.n112 B 0.019768f
C508 VTAIL.n113 B 0.010622f
C509 VTAIL.n114 B 0.025107f
C510 VTAIL.n115 B 0.011247f
C511 VTAIL.n116 B 0.019768f
C512 VTAIL.n117 B 0.010622f
C513 VTAIL.n118 B 0.025107f
C514 VTAIL.n119 B 0.011247f
C515 VTAIL.n120 B 0.019768f
C516 VTAIL.n121 B 0.010622f
C517 VTAIL.n122 B 0.025107f
C518 VTAIL.n123 B 0.011247f
C519 VTAIL.n124 B 0.137603f
C520 VTAIL.t0 B 0.041518f
C521 VTAIL.n125 B 0.018831f
C522 VTAIL.n126 B 0.014832f
C523 VTAIL.n127 B 0.010622f
C524 VTAIL.n128 B 1.44466f
C525 VTAIL.n129 B 0.019768f
C526 VTAIL.n130 B 0.010622f
C527 VTAIL.n131 B 0.011247f
C528 VTAIL.n132 B 0.025107f
C529 VTAIL.n133 B 0.025107f
C530 VTAIL.n134 B 0.011247f
C531 VTAIL.n135 B 0.010622f
C532 VTAIL.n136 B 0.019768f
C533 VTAIL.n137 B 0.019768f
C534 VTAIL.n138 B 0.010622f
C535 VTAIL.n139 B 0.011247f
C536 VTAIL.n140 B 0.025107f
C537 VTAIL.n141 B 0.025107f
C538 VTAIL.n142 B 0.011247f
C539 VTAIL.n143 B 0.010622f
C540 VTAIL.n144 B 0.019768f
C541 VTAIL.n145 B 0.019768f
C542 VTAIL.n146 B 0.010622f
C543 VTAIL.n147 B 0.011247f
C544 VTAIL.n148 B 0.025107f
C545 VTAIL.n149 B 0.025107f
C546 VTAIL.n150 B 0.011247f
C547 VTAIL.n151 B 0.010622f
C548 VTAIL.n152 B 0.019768f
C549 VTAIL.n153 B 0.019768f
C550 VTAIL.n154 B 0.010622f
C551 VTAIL.n155 B 0.011247f
C552 VTAIL.n156 B 0.025107f
C553 VTAIL.n157 B 0.025107f
C554 VTAIL.n158 B 0.011247f
C555 VTAIL.n159 B 0.010622f
C556 VTAIL.n160 B 0.019768f
C557 VTAIL.n161 B 0.019768f
C558 VTAIL.n162 B 0.010622f
C559 VTAIL.n163 B 0.011247f
C560 VTAIL.n164 B 0.025107f
C561 VTAIL.n165 B 0.025107f
C562 VTAIL.n166 B 0.011247f
C563 VTAIL.n167 B 0.010622f
C564 VTAIL.n168 B 0.019768f
C565 VTAIL.n169 B 0.019768f
C566 VTAIL.n170 B 0.010622f
C567 VTAIL.n171 B 0.010935f
C568 VTAIL.n172 B 0.010935f
C569 VTAIL.n173 B 0.025107f
C570 VTAIL.n174 B 0.025107f
C571 VTAIL.n175 B 0.011247f
C572 VTAIL.n176 B 0.010622f
C573 VTAIL.n177 B 0.019768f
C574 VTAIL.n178 B 0.019768f
C575 VTAIL.n179 B 0.010622f
C576 VTAIL.n180 B 0.011247f
C577 VTAIL.n181 B 0.025107f
C578 VTAIL.n182 B 0.051287f
C579 VTAIL.n183 B 0.011247f
C580 VTAIL.n184 B 0.010622f
C581 VTAIL.n185 B 0.044342f
C582 VTAIL.n186 B 0.02834f
C583 VTAIL.n187 B 1.45945f
C584 VTAIL.n188 B 0.026052f
C585 VTAIL.n189 B 0.019768f
C586 VTAIL.n190 B 0.010622f
C587 VTAIL.n191 B 0.025107f
C588 VTAIL.n192 B 0.011247f
C589 VTAIL.n193 B 0.019768f
C590 VTAIL.n194 B 0.010622f
C591 VTAIL.n195 B 0.025107f
C592 VTAIL.n196 B 0.011247f
C593 VTAIL.n197 B 0.019768f
C594 VTAIL.n198 B 0.010622f
C595 VTAIL.n199 B 0.025107f
C596 VTAIL.n200 B 0.025107f
C597 VTAIL.n201 B 0.011247f
C598 VTAIL.n202 B 0.019768f
C599 VTAIL.n203 B 0.010622f
C600 VTAIL.n204 B 0.025107f
C601 VTAIL.n205 B 0.011247f
C602 VTAIL.n206 B 0.019768f
C603 VTAIL.n207 B 0.010622f
C604 VTAIL.n208 B 0.025107f
C605 VTAIL.n209 B 0.011247f
C606 VTAIL.n210 B 0.019768f
C607 VTAIL.n211 B 0.010622f
C608 VTAIL.n212 B 0.025107f
C609 VTAIL.n213 B 0.011247f
C610 VTAIL.n214 B 0.019768f
C611 VTAIL.n215 B 0.010622f
C612 VTAIL.n216 B 0.025107f
C613 VTAIL.n217 B 0.011247f
C614 VTAIL.n218 B 0.137603f
C615 VTAIL.t2 B 0.041518f
C616 VTAIL.n219 B 0.018831f
C617 VTAIL.n220 B 0.014832f
C618 VTAIL.n221 B 0.010622f
C619 VTAIL.n222 B 1.44466f
C620 VTAIL.n223 B 0.019768f
C621 VTAIL.n224 B 0.010622f
C622 VTAIL.n225 B 0.011247f
C623 VTAIL.n226 B 0.025107f
C624 VTAIL.n227 B 0.025107f
C625 VTAIL.n228 B 0.011247f
C626 VTAIL.n229 B 0.010622f
C627 VTAIL.n230 B 0.019768f
C628 VTAIL.n231 B 0.019768f
C629 VTAIL.n232 B 0.010622f
C630 VTAIL.n233 B 0.011247f
C631 VTAIL.n234 B 0.025107f
C632 VTAIL.n235 B 0.025107f
C633 VTAIL.n236 B 0.011247f
C634 VTAIL.n237 B 0.010622f
C635 VTAIL.n238 B 0.019768f
C636 VTAIL.n239 B 0.019768f
C637 VTAIL.n240 B 0.010622f
C638 VTAIL.n241 B 0.011247f
C639 VTAIL.n242 B 0.025107f
C640 VTAIL.n243 B 0.025107f
C641 VTAIL.n244 B 0.011247f
C642 VTAIL.n245 B 0.010622f
C643 VTAIL.n246 B 0.019768f
C644 VTAIL.n247 B 0.019768f
C645 VTAIL.n248 B 0.010622f
C646 VTAIL.n249 B 0.011247f
C647 VTAIL.n250 B 0.025107f
C648 VTAIL.n251 B 0.025107f
C649 VTAIL.n252 B 0.011247f
C650 VTAIL.n253 B 0.010622f
C651 VTAIL.n254 B 0.019768f
C652 VTAIL.n255 B 0.019768f
C653 VTAIL.n256 B 0.010622f
C654 VTAIL.n257 B 0.011247f
C655 VTAIL.n258 B 0.025107f
C656 VTAIL.n259 B 0.025107f
C657 VTAIL.n260 B 0.011247f
C658 VTAIL.n261 B 0.010622f
C659 VTAIL.n262 B 0.019768f
C660 VTAIL.n263 B 0.019768f
C661 VTAIL.n264 B 0.010622f
C662 VTAIL.n265 B 0.010935f
C663 VTAIL.n266 B 0.010935f
C664 VTAIL.n267 B 0.025107f
C665 VTAIL.n268 B 0.025107f
C666 VTAIL.n269 B 0.011247f
C667 VTAIL.n270 B 0.010622f
C668 VTAIL.n271 B 0.019768f
C669 VTAIL.n272 B 0.019768f
C670 VTAIL.n273 B 0.010622f
C671 VTAIL.n274 B 0.011247f
C672 VTAIL.n275 B 0.025107f
C673 VTAIL.n276 B 0.051287f
C674 VTAIL.n277 B 0.011247f
C675 VTAIL.n278 B 0.010622f
C676 VTAIL.n279 B 0.044342f
C677 VTAIL.n280 B 0.02834f
C678 VTAIL.n281 B 1.3694f
C679 VTAIL.n282 B 0.026052f
C680 VTAIL.n283 B 0.019768f
C681 VTAIL.n284 B 0.010622f
C682 VTAIL.n285 B 0.025107f
C683 VTAIL.n286 B 0.011247f
C684 VTAIL.n287 B 0.019768f
C685 VTAIL.n288 B 0.010622f
C686 VTAIL.n289 B 0.025107f
C687 VTAIL.n290 B 0.011247f
C688 VTAIL.n291 B 0.019768f
C689 VTAIL.n292 B 0.010622f
C690 VTAIL.n293 B 0.025107f
C691 VTAIL.n294 B 0.011247f
C692 VTAIL.n295 B 0.019768f
C693 VTAIL.n296 B 0.010622f
C694 VTAIL.n297 B 0.025107f
C695 VTAIL.n298 B 0.011247f
C696 VTAIL.n299 B 0.019768f
C697 VTAIL.n300 B 0.010622f
C698 VTAIL.n301 B 0.025107f
C699 VTAIL.n302 B 0.011247f
C700 VTAIL.n303 B 0.019768f
C701 VTAIL.n304 B 0.010622f
C702 VTAIL.n305 B 0.025107f
C703 VTAIL.n306 B 0.011247f
C704 VTAIL.n307 B 0.019768f
C705 VTAIL.n308 B 0.010622f
C706 VTAIL.n309 B 0.025107f
C707 VTAIL.n310 B 0.011247f
C708 VTAIL.n311 B 0.137603f
C709 VTAIL.t1 B 0.041518f
C710 VTAIL.n312 B 0.018831f
C711 VTAIL.n313 B 0.014832f
C712 VTAIL.n314 B 0.010622f
C713 VTAIL.n315 B 1.44466f
C714 VTAIL.n316 B 0.019768f
C715 VTAIL.n317 B 0.010622f
C716 VTAIL.n318 B 0.011247f
C717 VTAIL.n319 B 0.025107f
C718 VTAIL.n320 B 0.025107f
C719 VTAIL.n321 B 0.011247f
C720 VTAIL.n322 B 0.010622f
C721 VTAIL.n323 B 0.019768f
C722 VTAIL.n324 B 0.019768f
C723 VTAIL.n325 B 0.010622f
C724 VTAIL.n326 B 0.011247f
C725 VTAIL.n327 B 0.025107f
C726 VTAIL.n328 B 0.025107f
C727 VTAIL.n329 B 0.011247f
C728 VTAIL.n330 B 0.010622f
C729 VTAIL.n331 B 0.019768f
C730 VTAIL.n332 B 0.019768f
C731 VTAIL.n333 B 0.010622f
C732 VTAIL.n334 B 0.011247f
C733 VTAIL.n335 B 0.025107f
C734 VTAIL.n336 B 0.025107f
C735 VTAIL.n337 B 0.011247f
C736 VTAIL.n338 B 0.010622f
C737 VTAIL.n339 B 0.019768f
C738 VTAIL.n340 B 0.019768f
C739 VTAIL.n341 B 0.010622f
C740 VTAIL.n342 B 0.011247f
C741 VTAIL.n343 B 0.025107f
C742 VTAIL.n344 B 0.025107f
C743 VTAIL.n345 B 0.011247f
C744 VTAIL.n346 B 0.010622f
C745 VTAIL.n347 B 0.019768f
C746 VTAIL.n348 B 0.019768f
C747 VTAIL.n349 B 0.010622f
C748 VTAIL.n350 B 0.011247f
C749 VTAIL.n351 B 0.025107f
C750 VTAIL.n352 B 0.025107f
C751 VTAIL.n353 B 0.025107f
C752 VTAIL.n354 B 0.011247f
C753 VTAIL.n355 B 0.010622f
C754 VTAIL.n356 B 0.019768f
C755 VTAIL.n357 B 0.019768f
C756 VTAIL.n358 B 0.010622f
C757 VTAIL.n359 B 0.010935f
C758 VTAIL.n360 B 0.010935f
C759 VTAIL.n361 B 0.025107f
C760 VTAIL.n362 B 0.025107f
C761 VTAIL.n363 B 0.011247f
C762 VTAIL.n364 B 0.010622f
C763 VTAIL.n365 B 0.019768f
C764 VTAIL.n366 B 0.019768f
C765 VTAIL.n367 B 0.010622f
C766 VTAIL.n368 B 0.011247f
C767 VTAIL.n369 B 0.025107f
C768 VTAIL.n370 B 0.051287f
C769 VTAIL.n371 B 0.011247f
C770 VTAIL.n372 B 0.010622f
C771 VTAIL.n373 B 0.044342f
C772 VTAIL.n374 B 0.02834f
C773 VTAIL.n375 B 1.31325f
C774 VP.t1 B 3.24763f
C775 VP.t0 B 2.96567f
C776 VP.n0 B 5.54582f
.ends

