* NGSPICE file created from diff_pair_sample_0393.ext - technology: sky130A

.subckt diff_pair_sample_0393 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=4.3485 pd=23.08 as=0 ps=0 w=11.15 l=0.49
X1 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=4.3485 pd=23.08 as=0 ps=0 w=11.15 l=0.49
X2 VDD1.t3 VP.t0 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.83975 pd=11.48 as=4.3485 ps=23.08 w=11.15 l=0.49
X3 VTAIL.t0 VN.t0 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=4.3485 pd=23.08 as=1.83975 ps=11.48 w=11.15 l=0.49
X4 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=4.3485 pd=23.08 as=0 ps=0 w=11.15 l=0.49
X5 VDD2.t2 VN.t1 VTAIL.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.83975 pd=11.48 as=4.3485 ps=23.08 w=11.15 l=0.49
X6 VDD2.t1 VN.t2 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.83975 pd=11.48 as=4.3485 ps=23.08 w=11.15 l=0.49
X7 VTAIL.t2 VN.t3 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=4.3485 pd=23.08 as=1.83975 ps=11.48 w=11.15 l=0.49
X8 VTAIL.t6 VP.t1 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=4.3485 pd=23.08 as=1.83975 ps=11.48 w=11.15 l=0.49
X9 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=4.3485 pd=23.08 as=0 ps=0 w=11.15 l=0.49
X10 VTAIL.t5 VP.t2 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=4.3485 pd=23.08 as=1.83975 ps=11.48 w=11.15 l=0.49
X11 VDD1.t0 VP.t3 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.83975 pd=11.48 as=4.3485 ps=23.08 w=11.15 l=0.49
R0 B.n80 B.t8 755.052
R1 B.n78 B.t4 755.052
R2 B.n328 B.t15 755.052
R3 B.n325 B.t11 755.052
R4 B.n573 B.n572 585
R5 B.n252 B.n76 585
R6 B.n251 B.n250 585
R7 B.n249 B.n248 585
R8 B.n247 B.n246 585
R9 B.n245 B.n244 585
R10 B.n243 B.n242 585
R11 B.n241 B.n240 585
R12 B.n239 B.n238 585
R13 B.n237 B.n236 585
R14 B.n235 B.n234 585
R15 B.n233 B.n232 585
R16 B.n231 B.n230 585
R17 B.n229 B.n228 585
R18 B.n227 B.n226 585
R19 B.n225 B.n224 585
R20 B.n223 B.n222 585
R21 B.n221 B.n220 585
R22 B.n219 B.n218 585
R23 B.n217 B.n216 585
R24 B.n215 B.n214 585
R25 B.n213 B.n212 585
R26 B.n211 B.n210 585
R27 B.n209 B.n208 585
R28 B.n207 B.n206 585
R29 B.n205 B.n204 585
R30 B.n203 B.n202 585
R31 B.n201 B.n200 585
R32 B.n199 B.n198 585
R33 B.n197 B.n196 585
R34 B.n195 B.n194 585
R35 B.n193 B.n192 585
R36 B.n191 B.n190 585
R37 B.n189 B.n188 585
R38 B.n187 B.n186 585
R39 B.n185 B.n184 585
R40 B.n183 B.n182 585
R41 B.n181 B.n180 585
R42 B.n179 B.n178 585
R43 B.n176 B.n175 585
R44 B.n174 B.n173 585
R45 B.n172 B.n171 585
R46 B.n170 B.n169 585
R47 B.n168 B.n167 585
R48 B.n166 B.n165 585
R49 B.n164 B.n163 585
R50 B.n162 B.n161 585
R51 B.n160 B.n159 585
R52 B.n158 B.n157 585
R53 B.n155 B.n154 585
R54 B.n153 B.n152 585
R55 B.n151 B.n150 585
R56 B.n149 B.n148 585
R57 B.n147 B.n146 585
R58 B.n145 B.n144 585
R59 B.n143 B.n142 585
R60 B.n141 B.n140 585
R61 B.n139 B.n138 585
R62 B.n137 B.n136 585
R63 B.n135 B.n134 585
R64 B.n133 B.n132 585
R65 B.n131 B.n130 585
R66 B.n129 B.n128 585
R67 B.n127 B.n126 585
R68 B.n125 B.n124 585
R69 B.n123 B.n122 585
R70 B.n121 B.n120 585
R71 B.n119 B.n118 585
R72 B.n117 B.n116 585
R73 B.n115 B.n114 585
R74 B.n113 B.n112 585
R75 B.n111 B.n110 585
R76 B.n109 B.n108 585
R77 B.n107 B.n106 585
R78 B.n105 B.n104 585
R79 B.n103 B.n102 585
R80 B.n101 B.n100 585
R81 B.n99 B.n98 585
R82 B.n97 B.n96 585
R83 B.n95 B.n94 585
R84 B.n93 B.n92 585
R85 B.n91 B.n90 585
R86 B.n89 B.n88 585
R87 B.n87 B.n86 585
R88 B.n85 B.n84 585
R89 B.n83 B.n82 585
R90 B.n33 B.n32 585
R91 B.n578 B.n577 585
R92 B.n571 B.n77 585
R93 B.n77 B.n30 585
R94 B.n570 B.n29 585
R95 B.n582 B.n29 585
R96 B.n569 B.n28 585
R97 B.n583 B.n28 585
R98 B.n568 B.n27 585
R99 B.n584 B.n27 585
R100 B.n567 B.n566 585
R101 B.n566 B.n26 585
R102 B.n565 B.n22 585
R103 B.n590 B.n22 585
R104 B.n564 B.n21 585
R105 B.n591 B.n21 585
R106 B.n563 B.n20 585
R107 B.n592 B.n20 585
R108 B.n562 B.n561 585
R109 B.n561 B.n16 585
R110 B.n560 B.n15 585
R111 B.n598 B.n15 585
R112 B.n559 B.n14 585
R113 B.n599 B.n14 585
R114 B.n558 B.n13 585
R115 B.n600 B.n13 585
R116 B.n557 B.n556 585
R117 B.n556 B.n12 585
R118 B.n555 B.n554 585
R119 B.n555 B.n8 585
R120 B.n553 B.n7 585
R121 B.n607 B.n7 585
R122 B.n552 B.n6 585
R123 B.n608 B.n6 585
R124 B.n551 B.n5 585
R125 B.n609 B.n5 585
R126 B.n550 B.n549 585
R127 B.n549 B.n4 585
R128 B.n548 B.n253 585
R129 B.n548 B.n547 585
R130 B.n537 B.n254 585
R131 B.n540 B.n254 585
R132 B.n539 B.n538 585
R133 B.n541 B.n539 585
R134 B.n536 B.n258 585
R135 B.n262 B.n258 585
R136 B.n535 B.n534 585
R137 B.n534 B.n533 585
R138 B.n260 B.n259 585
R139 B.n261 B.n260 585
R140 B.n526 B.n525 585
R141 B.n527 B.n526 585
R142 B.n524 B.n267 585
R143 B.n267 B.n266 585
R144 B.n523 B.n522 585
R145 B.n522 B.n521 585
R146 B.n269 B.n268 585
R147 B.n514 B.n269 585
R148 B.n513 B.n512 585
R149 B.n515 B.n513 585
R150 B.n511 B.n274 585
R151 B.n274 B.n273 585
R152 B.n510 B.n509 585
R153 B.n509 B.n508 585
R154 B.n276 B.n275 585
R155 B.n277 B.n276 585
R156 B.n504 B.n503 585
R157 B.n280 B.n279 585
R158 B.n500 B.n499 585
R159 B.n501 B.n500 585
R160 B.n498 B.n324 585
R161 B.n497 B.n496 585
R162 B.n495 B.n494 585
R163 B.n493 B.n492 585
R164 B.n491 B.n490 585
R165 B.n489 B.n488 585
R166 B.n487 B.n486 585
R167 B.n485 B.n484 585
R168 B.n483 B.n482 585
R169 B.n481 B.n480 585
R170 B.n479 B.n478 585
R171 B.n477 B.n476 585
R172 B.n475 B.n474 585
R173 B.n473 B.n472 585
R174 B.n471 B.n470 585
R175 B.n469 B.n468 585
R176 B.n467 B.n466 585
R177 B.n465 B.n464 585
R178 B.n463 B.n462 585
R179 B.n461 B.n460 585
R180 B.n459 B.n458 585
R181 B.n457 B.n456 585
R182 B.n455 B.n454 585
R183 B.n453 B.n452 585
R184 B.n451 B.n450 585
R185 B.n449 B.n448 585
R186 B.n447 B.n446 585
R187 B.n445 B.n444 585
R188 B.n443 B.n442 585
R189 B.n441 B.n440 585
R190 B.n439 B.n438 585
R191 B.n437 B.n436 585
R192 B.n435 B.n434 585
R193 B.n433 B.n432 585
R194 B.n431 B.n430 585
R195 B.n429 B.n428 585
R196 B.n427 B.n426 585
R197 B.n425 B.n424 585
R198 B.n423 B.n422 585
R199 B.n421 B.n420 585
R200 B.n419 B.n418 585
R201 B.n417 B.n416 585
R202 B.n415 B.n414 585
R203 B.n413 B.n412 585
R204 B.n411 B.n410 585
R205 B.n409 B.n408 585
R206 B.n407 B.n406 585
R207 B.n405 B.n404 585
R208 B.n403 B.n402 585
R209 B.n401 B.n400 585
R210 B.n399 B.n398 585
R211 B.n397 B.n396 585
R212 B.n395 B.n394 585
R213 B.n393 B.n392 585
R214 B.n391 B.n390 585
R215 B.n389 B.n388 585
R216 B.n387 B.n386 585
R217 B.n385 B.n384 585
R218 B.n383 B.n382 585
R219 B.n381 B.n380 585
R220 B.n379 B.n378 585
R221 B.n377 B.n376 585
R222 B.n375 B.n374 585
R223 B.n373 B.n372 585
R224 B.n371 B.n370 585
R225 B.n369 B.n368 585
R226 B.n367 B.n366 585
R227 B.n365 B.n364 585
R228 B.n363 B.n362 585
R229 B.n361 B.n360 585
R230 B.n359 B.n358 585
R231 B.n357 B.n356 585
R232 B.n355 B.n354 585
R233 B.n353 B.n352 585
R234 B.n351 B.n350 585
R235 B.n349 B.n348 585
R236 B.n347 B.n346 585
R237 B.n345 B.n344 585
R238 B.n343 B.n342 585
R239 B.n341 B.n340 585
R240 B.n339 B.n338 585
R241 B.n337 B.n336 585
R242 B.n335 B.n334 585
R243 B.n333 B.n332 585
R244 B.n331 B.n323 585
R245 B.n501 B.n323 585
R246 B.n505 B.n278 585
R247 B.n278 B.n277 585
R248 B.n507 B.n506 585
R249 B.n508 B.n507 585
R250 B.n272 B.n271 585
R251 B.n273 B.n272 585
R252 B.n517 B.n516 585
R253 B.n516 B.n515 585
R254 B.n518 B.n270 585
R255 B.n514 B.n270 585
R256 B.n520 B.n519 585
R257 B.n521 B.n520 585
R258 B.n265 B.n264 585
R259 B.n266 B.n265 585
R260 B.n529 B.n528 585
R261 B.n528 B.n527 585
R262 B.n530 B.n263 585
R263 B.n263 B.n261 585
R264 B.n532 B.n531 585
R265 B.n533 B.n532 585
R266 B.n257 B.n256 585
R267 B.n262 B.n257 585
R268 B.n543 B.n542 585
R269 B.n542 B.n541 585
R270 B.n544 B.n255 585
R271 B.n540 B.n255 585
R272 B.n546 B.n545 585
R273 B.n547 B.n546 585
R274 B.n3 B.n0 585
R275 B.n4 B.n3 585
R276 B.n606 B.n1 585
R277 B.n607 B.n606 585
R278 B.n605 B.n604 585
R279 B.n605 B.n8 585
R280 B.n603 B.n9 585
R281 B.n12 B.n9 585
R282 B.n602 B.n601 585
R283 B.n601 B.n600 585
R284 B.n11 B.n10 585
R285 B.n599 B.n11 585
R286 B.n597 B.n596 585
R287 B.n598 B.n597 585
R288 B.n595 B.n17 585
R289 B.n17 B.n16 585
R290 B.n594 B.n593 585
R291 B.n593 B.n592 585
R292 B.n19 B.n18 585
R293 B.n591 B.n19 585
R294 B.n589 B.n588 585
R295 B.n590 B.n589 585
R296 B.n587 B.n23 585
R297 B.n26 B.n23 585
R298 B.n586 B.n585 585
R299 B.n585 B.n584 585
R300 B.n25 B.n24 585
R301 B.n583 B.n25 585
R302 B.n581 B.n580 585
R303 B.n582 B.n581 585
R304 B.n579 B.n31 585
R305 B.n31 B.n30 585
R306 B.n610 B.n609 585
R307 B.n608 B.n2 585
R308 B.n577 B.n31 458.866
R309 B.n573 B.n77 458.866
R310 B.n323 B.n276 458.866
R311 B.n503 B.n278 458.866
R312 B.n575 B.n574 256.663
R313 B.n575 B.n75 256.663
R314 B.n575 B.n74 256.663
R315 B.n575 B.n73 256.663
R316 B.n575 B.n72 256.663
R317 B.n575 B.n71 256.663
R318 B.n575 B.n70 256.663
R319 B.n575 B.n69 256.663
R320 B.n575 B.n68 256.663
R321 B.n575 B.n67 256.663
R322 B.n575 B.n66 256.663
R323 B.n575 B.n65 256.663
R324 B.n575 B.n64 256.663
R325 B.n575 B.n63 256.663
R326 B.n575 B.n62 256.663
R327 B.n575 B.n61 256.663
R328 B.n575 B.n60 256.663
R329 B.n575 B.n59 256.663
R330 B.n575 B.n58 256.663
R331 B.n575 B.n57 256.663
R332 B.n575 B.n56 256.663
R333 B.n575 B.n55 256.663
R334 B.n575 B.n54 256.663
R335 B.n575 B.n53 256.663
R336 B.n575 B.n52 256.663
R337 B.n575 B.n51 256.663
R338 B.n575 B.n50 256.663
R339 B.n575 B.n49 256.663
R340 B.n575 B.n48 256.663
R341 B.n575 B.n47 256.663
R342 B.n575 B.n46 256.663
R343 B.n575 B.n45 256.663
R344 B.n575 B.n44 256.663
R345 B.n575 B.n43 256.663
R346 B.n575 B.n42 256.663
R347 B.n575 B.n41 256.663
R348 B.n575 B.n40 256.663
R349 B.n575 B.n39 256.663
R350 B.n575 B.n38 256.663
R351 B.n575 B.n37 256.663
R352 B.n575 B.n36 256.663
R353 B.n575 B.n35 256.663
R354 B.n575 B.n34 256.663
R355 B.n576 B.n575 256.663
R356 B.n502 B.n501 256.663
R357 B.n501 B.n281 256.663
R358 B.n501 B.n282 256.663
R359 B.n501 B.n283 256.663
R360 B.n501 B.n284 256.663
R361 B.n501 B.n285 256.663
R362 B.n501 B.n286 256.663
R363 B.n501 B.n287 256.663
R364 B.n501 B.n288 256.663
R365 B.n501 B.n289 256.663
R366 B.n501 B.n290 256.663
R367 B.n501 B.n291 256.663
R368 B.n501 B.n292 256.663
R369 B.n501 B.n293 256.663
R370 B.n501 B.n294 256.663
R371 B.n501 B.n295 256.663
R372 B.n501 B.n296 256.663
R373 B.n501 B.n297 256.663
R374 B.n501 B.n298 256.663
R375 B.n501 B.n299 256.663
R376 B.n501 B.n300 256.663
R377 B.n501 B.n301 256.663
R378 B.n501 B.n302 256.663
R379 B.n501 B.n303 256.663
R380 B.n501 B.n304 256.663
R381 B.n501 B.n305 256.663
R382 B.n501 B.n306 256.663
R383 B.n501 B.n307 256.663
R384 B.n501 B.n308 256.663
R385 B.n501 B.n309 256.663
R386 B.n501 B.n310 256.663
R387 B.n501 B.n311 256.663
R388 B.n501 B.n312 256.663
R389 B.n501 B.n313 256.663
R390 B.n501 B.n314 256.663
R391 B.n501 B.n315 256.663
R392 B.n501 B.n316 256.663
R393 B.n501 B.n317 256.663
R394 B.n501 B.n318 256.663
R395 B.n501 B.n319 256.663
R396 B.n501 B.n320 256.663
R397 B.n501 B.n321 256.663
R398 B.n501 B.n322 256.663
R399 B.n612 B.n611 256.663
R400 B.n82 B.n33 163.367
R401 B.n86 B.n85 163.367
R402 B.n90 B.n89 163.367
R403 B.n94 B.n93 163.367
R404 B.n98 B.n97 163.367
R405 B.n102 B.n101 163.367
R406 B.n106 B.n105 163.367
R407 B.n110 B.n109 163.367
R408 B.n114 B.n113 163.367
R409 B.n118 B.n117 163.367
R410 B.n122 B.n121 163.367
R411 B.n126 B.n125 163.367
R412 B.n130 B.n129 163.367
R413 B.n134 B.n133 163.367
R414 B.n138 B.n137 163.367
R415 B.n142 B.n141 163.367
R416 B.n146 B.n145 163.367
R417 B.n150 B.n149 163.367
R418 B.n154 B.n153 163.367
R419 B.n159 B.n158 163.367
R420 B.n163 B.n162 163.367
R421 B.n167 B.n166 163.367
R422 B.n171 B.n170 163.367
R423 B.n175 B.n174 163.367
R424 B.n180 B.n179 163.367
R425 B.n184 B.n183 163.367
R426 B.n188 B.n187 163.367
R427 B.n192 B.n191 163.367
R428 B.n196 B.n195 163.367
R429 B.n200 B.n199 163.367
R430 B.n204 B.n203 163.367
R431 B.n208 B.n207 163.367
R432 B.n212 B.n211 163.367
R433 B.n216 B.n215 163.367
R434 B.n220 B.n219 163.367
R435 B.n224 B.n223 163.367
R436 B.n228 B.n227 163.367
R437 B.n232 B.n231 163.367
R438 B.n236 B.n235 163.367
R439 B.n240 B.n239 163.367
R440 B.n244 B.n243 163.367
R441 B.n248 B.n247 163.367
R442 B.n250 B.n76 163.367
R443 B.n509 B.n276 163.367
R444 B.n509 B.n274 163.367
R445 B.n513 B.n274 163.367
R446 B.n513 B.n269 163.367
R447 B.n522 B.n269 163.367
R448 B.n522 B.n267 163.367
R449 B.n526 B.n267 163.367
R450 B.n526 B.n260 163.367
R451 B.n534 B.n260 163.367
R452 B.n534 B.n258 163.367
R453 B.n539 B.n258 163.367
R454 B.n539 B.n254 163.367
R455 B.n548 B.n254 163.367
R456 B.n549 B.n548 163.367
R457 B.n549 B.n5 163.367
R458 B.n6 B.n5 163.367
R459 B.n7 B.n6 163.367
R460 B.n555 B.n7 163.367
R461 B.n556 B.n555 163.367
R462 B.n556 B.n13 163.367
R463 B.n14 B.n13 163.367
R464 B.n15 B.n14 163.367
R465 B.n561 B.n15 163.367
R466 B.n561 B.n20 163.367
R467 B.n21 B.n20 163.367
R468 B.n22 B.n21 163.367
R469 B.n566 B.n22 163.367
R470 B.n566 B.n27 163.367
R471 B.n28 B.n27 163.367
R472 B.n29 B.n28 163.367
R473 B.n77 B.n29 163.367
R474 B.n500 B.n280 163.367
R475 B.n500 B.n324 163.367
R476 B.n496 B.n495 163.367
R477 B.n492 B.n491 163.367
R478 B.n488 B.n487 163.367
R479 B.n484 B.n483 163.367
R480 B.n480 B.n479 163.367
R481 B.n476 B.n475 163.367
R482 B.n472 B.n471 163.367
R483 B.n468 B.n467 163.367
R484 B.n464 B.n463 163.367
R485 B.n460 B.n459 163.367
R486 B.n456 B.n455 163.367
R487 B.n452 B.n451 163.367
R488 B.n448 B.n447 163.367
R489 B.n444 B.n443 163.367
R490 B.n440 B.n439 163.367
R491 B.n436 B.n435 163.367
R492 B.n432 B.n431 163.367
R493 B.n428 B.n427 163.367
R494 B.n424 B.n423 163.367
R495 B.n420 B.n419 163.367
R496 B.n416 B.n415 163.367
R497 B.n412 B.n411 163.367
R498 B.n408 B.n407 163.367
R499 B.n404 B.n403 163.367
R500 B.n400 B.n399 163.367
R501 B.n396 B.n395 163.367
R502 B.n392 B.n391 163.367
R503 B.n388 B.n387 163.367
R504 B.n384 B.n383 163.367
R505 B.n380 B.n379 163.367
R506 B.n376 B.n375 163.367
R507 B.n372 B.n371 163.367
R508 B.n368 B.n367 163.367
R509 B.n364 B.n363 163.367
R510 B.n360 B.n359 163.367
R511 B.n356 B.n355 163.367
R512 B.n352 B.n351 163.367
R513 B.n348 B.n347 163.367
R514 B.n344 B.n343 163.367
R515 B.n340 B.n339 163.367
R516 B.n336 B.n335 163.367
R517 B.n332 B.n323 163.367
R518 B.n507 B.n278 163.367
R519 B.n507 B.n272 163.367
R520 B.n516 B.n272 163.367
R521 B.n516 B.n270 163.367
R522 B.n520 B.n270 163.367
R523 B.n520 B.n265 163.367
R524 B.n528 B.n265 163.367
R525 B.n528 B.n263 163.367
R526 B.n532 B.n263 163.367
R527 B.n532 B.n257 163.367
R528 B.n542 B.n257 163.367
R529 B.n542 B.n255 163.367
R530 B.n546 B.n255 163.367
R531 B.n546 B.n3 163.367
R532 B.n610 B.n3 163.367
R533 B.n606 B.n2 163.367
R534 B.n606 B.n605 163.367
R535 B.n605 B.n9 163.367
R536 B.n601 B.n9 163.367
R537 B.n601 B.n11 163.367
R538 B.n597 B.n11 163.367
R539 B.n597 B.n17 163.367
R540 B.n593 B.n17 163.367
R541 B.n593 B.n19 163.367
R542 B.n589 B.n19 163.367
R543 B.n589 B.n23 163.367
R544 B.n585 B.n23 163.367
R545 B.n585 B.n25 163.367
R546 B.n581 B.n25 163.367
R547 B.n581 B.n31 163.367
R548 B.n78 B.t6 89.0536
R549 B.n328 B.t17 89.0536
R550 B.n80 B.t9 89.0398
R551 B.n325 B.t14 89.0398
R552 B.n501 B.n277 75.6778
R553 B.n575 B.n30 75.6778
R554 B.n79 B.t7 73.1505
R555 B.n329 B.t16 73.1505
R556 B.n81 B.t10 73.1368
R557 B.n326 B.t13 73.1368
R558 B.n577 B.n576 71.676
R559 B.n82 B.n34 71.676
R560 B.n86 B.n35 71.676
R561 B.n90 B.n36 71.676
R562 B.n94 B.n37 71.676
R563 B.n98 B.n38 71.676
R564 B.n102 B.n39 71.676
R565 B.n106 B.n40 71.676
R566 B.n110 B.n41 71.676
R567 B.n114 B.n42 71.676
R568 B.n118 B.n43 71.676
R569 B.n122 B.n44 71.676
R570 B.n126 B.n45 71.676
R571 B.n130 B.n46 71.676
R572 B.n134 B.n47 71.676
R573 B.n138 B.n48 71.676
R574 B.n142 B.n49 71.676
R575 B.n146 B.n50 71.676
R576 B.n150 B.n51 71.676
R577 B.n154 B.n52 71.676
R578 B.n159 B.n53 71.676
R579 B.n163 B.n54 71.676
R580 B.n167 B.n55 71.676
R581 B.n171 B.n56 71.676
R582 B.n175 B.n57 71.676
R583 B.n180 B.n58 71.676
R584 B.n184 B.n59 71.676
R585 B.n188 B.n60 71.676
R586 B.n192 B.n61 71.676
R587 B.n196 B.n62 71.676
R588 B.n200 B.n63 71.676
R589 B.n204 B.n64 71.676
R590 B.n208 B.n65 71.676
R591 B.n212 B.n66 71.676
R592 B.n216 B.n67 71.676
R593 B.n220 B.n68 71.676
R594 B.n224 B.n69 71.676
R595 B.n228 B.n70 71.676
R596 B.n232 B.n71 71.676
R597 B.n236 B.n72 71.676
R598 B.n240 B.n73 71.676
R599 B.n244 B.n74 71.676
R600 B.n248 B.n75 71.676
R601 B.n574 B.n76 71.676
R602 B.n574 B.n573 71.676
R603 B.n250 B.n75 71.676
R604 B.n247 B.n74 71.676
R605 B.n243 B.n73 71.676
R606 B.n239 B.n72 71.676
R607 B.n235 B.n71 71.676
R608 B.n231 B.n70 71.676
R609 B.n227 B.n69 71.676
R610 B.n223 B.n68 71.676
R611 B.n219 B.n67 71.676
R612 B.n215 B.n66 71.676
R613 B.n211 B.n65 71.676
R614 B.n207 B.n64 71.676
R615 B.n203 B.n63 71.676
R616 B.n199 B.n62 71.676
R617 B.n195 B.n61 71.676
R618 B.n191 B.n60 71.676
R619 B.n187 B.n59 71.676
R620 B.n183 B.n58 71.676
R621 B.n179 B.n57 71.676
R622 B.n174 B.n56 71.676
R623 B.n170 B.n55 71.676
R624 B.n166 B.n54 71.676
R625 B.n162 B.n53 71.676
R626 B.n158 B.n52 71.676
R627 B.n153 B.n51 71.676
R628 B.n149 B.n50 71.676
R629 B.n145 B.n49 71.676
R630 B.n141 B.n48 71.676
R631 B.n137 B.n47 71.676
R632 B.n133 B.n46 71.676
R633 B.n129 B.n45 71.676
R634 B.n125 B.n44 71.676
R635 B.n121 B.n43 71.676
R636 B.n117 B.n42 71.676
R637 B.n113 B.n41 71.676
R638 B.n109 B.n40 71.676
R639 B.n105 B.n39 71.676
R640 B.n101 B.n38 71.676
R641 B.n97 B.n37 71.676
R642 B.n93 B.n36 71.676
R643 B.n89 B.n35 71.676
R644 B.n85 B.n34 71.676
R645 B.n576 B.n33 71.676
R646 B.n503 B.n502 71.676
R647 B.n324 B.n281 71.676
R648 B.n495 B.n282 71.676
R649 B.n491 B.n283 71.676
R650 B.n487 B.n284 71.676
R651 B.n483 B.n285 71.676
R652 B.n479 B.n286 71.676
R653 B.n475 B.n287 71.676
R654 B.n471 B.n288 71.676
R655 B.n467 B.n289 71.676
R656 B.n463 B.n290 71.676
R657 B.n459 B.n291 71.676
R658 B.n455 B.n292 71.676
R659 B.n451 B.n293 71.676
R660 B.n447 B.n294 71.676
R661 B.n443 B.n295 71.676
R662 B.n439 B.n296 71.676
R663 B.n435 B.n297 71.676
R664 B.n431 B.n298 71.676
R665 B.n427 B.n299 71.676
R666 B.n423 B.n300 71.676
R667 B.n419 B.n301 71.676
R668 B.n415 B.n302 71.676
R669 B.n411 B.n303 71.676
R670 B.n407 B.n304 71.676
R671 B.n403 B.n305 71.676
R672 B.n399 B.n306 71.676
R673 B.n395 B.n307 71.676
R674 B.n391 B.n308 71.676
R675 B.n387 B.n309 71.676
R676 B.n383 B.n310 71.676
R677 B.n379 B.n311 71.676
R678 B.n375 B.n312 71.676
R679 B.n371 B.n313 71.676
R680 B.n367 B.n314 71.676
R681 B.n363 B.n315 71.676
R682 B.n359 B.n316 71.676
R683 B.n355 B.n317 71.676
R684 B.n351 B.n318 71.676
R685 B.n347 B.n319 71.676
R686 B.n343 B.n320 71.676
R687 B.n339 B.n321 71.676
R688 B.n335 B.n322 71.676
R689 B.n502 B.n280 71.676
R690 B.n496 B.n281 71.676
R691 B.n492 B.n282 71.676
R692 B.n488 B.n283 71.676
R693 B.n484 B.n284 71.676
R694 B.n480 B.n285 71.676
R695 B.n476 B.n286 71.676
R696 B.n472 B.n287 71.676
R697 B.n468 B.n288 71.676
R698 B.n464 B.n289 71.676
R699 B.n460 B.n290 71.676
R700 B.n456 B.n291 71.676
R701 B.n452 B.n292 71.676
R702 B.n448 B.n293 71.676
R703 B.n444 B.n294 71.676
R704 B.n440 B.n295 71.676
R705 B.n436 B.n296 71.676
R706 B.n432 B.n297 71.676
R707 B.n428 B.n298 71.676
R708 B.n424 B.n299 71.676
R709 B.n420 B.n300 71.676
R710 B.n416 B.n301 71.676
R711 B.n412 B.n302 71.676
R712 B.n408 B.n303 71.676
R713 B.n404 B.n304 71.676
R714 B.n400 B.n305 71.676
R715 B.n396 B.n306 71.676
R716 B.n392 B.n307 71.676
R717 B.n388 B.n308 71.676
R718 B.n384 B.n309 71.676
R719 B.n380 B.n310 71.676
R720 B.n376 B.n311 71.676
R721 B.n372 B.n312 71.676
R722 B.n368 B.n313 71.676
R723 B.n364 B.n314 71.676
R724 B.n360 B.n315 71.676
R725 B.n356 B.n316 71.676
R726 B.n352 B.n317 71.676
R727 B.n348 B.n318 71.676
R728 B.n344 B.n319 71.676
R729 B.n340 B.n320 71.676
R730 B.n336 B.n321 71.676
R731 B.n332 B.n322 71.676
R732 B.n611 B.n610 71.676
R733 B.n611 B.n2 71.676
R734 B.n156 B.n81 59.5399
R735 B.n177 B.n79 59.5399
R736 B.n330 B.n329 59.5399
R737 B.n327 B.n326 59.5399
R738 B.n508 B.n277 45.5408
R739 B.n508 B.n273 45.5408
R740 B.n515 B.n273 45.5408
R741 B.n515 B.n514 45.5408
R742 B.n521 B.n266 45.5408
R743 B.n527 B.n266 45.5408
R744 B.n527 B.n261 45.5408
R745 B.n533 B.n261 45.5408
R746 B.n533 B.n262 45.5408
R747 B.n541 B.n540 45.5408
R748 B.n547 B.n4 45.5408
R749 B.n609 B.n4 45.5408
R750 B.n609 B.n608 45.5408
R751 B.n608 B.n607 45.5408
R752 B.n607 B.n8 45.5408
R753 B.n600 B.n12 45.5408
R754 B.n599 B.n598 45.5408
R755 B.n598 B.n16 45.5408
R756 B.n592 B.n16 45.5408
R757 B.n592 B.n591 45.5408
R758 B.n591 B.n590 45.5408
R759 B.n584 B.n26 45.5408
R760 B.n584 B.n583 45.5408
R761 B.n583 B.n582 45.5408
R762 B.n582 B.n30 45.5408
R763 B.n541 B.t2 32.8163
R764 B.n600 B.t1 32.8163
R765 B.n540 B.t3 31.4769
R766 B.n12 B.t0 31.4769
R767 B.n514 B.t12 30.1375
R768 B.n26 B.t5 30.1375
R769 B.n505 B.n504 29.8151
R770 B.n331 B.n275 29.8151
R771 B.n572 B.n571 29.8151
R772 B.n579 B.n578 29.8151
R773 B B.n612 18.0485
R774 B.n81 B.n80 15.9035
R775 B.n79 B.n78 15.9035
R776 B.n329 B.n328 15.9035
R777 B.n326 B.n325 15.9035
R778 B.n521 B.t12 15.4038
R779 B.n590 B.t5 15.4038
R780 B.n547 B.t3 14.0644
R781 B.t0 B.n8 14.0644
R782 B.n262 B.t2 12.725
R783 B.t1 B.n599 12.725
R784 B.n506 B.n505 10.6151
R785 B.n506 B.n271 10.6151
R786 B.n517 B.n271 10.6151
R787 B.n518 B.n517 10.6151
R788 B.n519 B.n518 10.6151
R789 B.n519 B.n264 10.6151
R790 B.n529 B.n264 10.6151
R791 B.n530 B.n529 10.6151
R792 B.n531 B.n530 10.6151
R793 B.n531 B.n256 10.6151
R794 B.n543 B.n256 10.6151
R795 B.n544 B.n543 10.6151
R796 B.n545 B.n544 10.6151
R797 B.n545 B.n0 10.6151
R798 B.n504 B.n279 10.6151
R799 B.n499 B.n279 10.6151
R800 B.n499 B.n498 10.6151
R801 B.n498 B.n497 10.6151
R802 B.n497 B.n494 10.6151
R803 B.n494 B.n493 10.6151
R804 B.n493 B.n490 10.6151
R805 B.n490 B.n489 10.6151
R806 B.n489 B.n486 10.6151
R807 B.n486 B.n485 10.6151
R808 B.n485 B.n482 10.6151
R809 B.n482 B.n481 10.6151
R810 B.n481 B.n478 10.6151
R811 B.n478 B.n477 10.6151
R812 B.n477 B.n474 10.6151
R813 B.n474 B.n473 10.6151
R814 B.n473 B.n470 10.6151
R815 B.n470 B.n469 10.6151
R816 B.n469 B.n466 10.6151
R817 B.n466 B.n465 10.6151
R818 B.n465 B.n462 10.6151
R819 B.n462 B.n461 10.6151
R820 B.n461 B.n458 10.6151
R821 B.n458 B.n457 10.6151
R822 B.n457 B.n454 10.6151
R823 B.n454 B.n453 10.6151
R824 B.n453 B.n450 10.6151
R825 B.n450 B.n449 10.6151
R826 B.n449 B.n446 10.6151
R827 B.n446 B.n445 10.6151
R828 B.n445 B.n442 10.6151
R829 B.n442 B.n441 10.6151
R830 B.n441 B.n438 10.6151
R831 B.n438 B.n437 10.6151
R832 B.n437 B.n434 10.6151
R833 B.n434 B.n433 10.6151
R834 B.n433 B.n430 10.6151
R835 B.n430 B.n429 10.6151
R836 B.n426 B.n425 10.6151
R837 B.n425 B.n422 10.6151
R838 B.n422 B.n421 10.6151
R839 B.n421 B.n418 10.6151
R840 B.n418 B.n417 10.6151
R841 B.n417 B.n414 10.6151
R842 B.n414 B.n413 10.6151
R843 B.n413 B.n410 10.6151
R844 B.n410 B.n409 10.6151
R845 B.n406 B.n405 10.6151
R846 B.n405 B.n402 10.6151
R847 B.n402 B.n401 10.6151
R848 B.n401 B.n398 10.6151
R849 B.n398 B.n397 10.6151
R850 B.n397 B.n394 10.6151
R851 B.n394 B.n393 10.6151
R852 B.n393 B.n390 10.6151
R853 B.n390 B.n389 10.6151
R854 B.n389 B.n386 10.6151
R855 B.n386 B.n385 10.6151
R856 B.n385 B.n382 10.6151
R857 B.n382 B.n381 10.6151
R858 B.n381 B.n378 10.6151
R859 B.n378 B.n377 10.6151
R860 B.n377 B.n374 10.6151
R861 B.n374 B.n373 10.6151
R862 B.n373 B.n370 10.6151
R863 B.n370 B.n369 10.6151
R864 B.n369 B.n366 10.6151
R865 B.n366 B.n365 10.6151
R866 B.n365 B.n362 10.6151
R867 B.n362 B.n361 10.6151
R868 B.n361 B.n358 10.6151
R869 B.n358 B.n357 10.6151
R870 B.n357 B.n354 10.6151
R871 B.n354 B.n353 10.6151
R872 B.n353 B.n350 10.6151
R873 B.n350 B.n349 10.6151
R874 B.n349 B.n346 10.6151
R875 B.n346 B.n345 10.6151
R876 B.n345 B.n342 10.6151
R877 B.n342 B.n341 10.6151
R878 B.n341 B.n338 10.6151
R879 B.n338 B.n337 10.6151
R880 B.n337 B.n334 10.6151
R881 B.n334 B.n333 10.6151
R882 B.n333 B.n331 10.6151
R883 B.n510 B.n275 10.6151
R884 B.n511 B.n510 10.6151
R885 B.n512 B.n511 10.6151
R886 B.n512 B.n268 10.6151
R887 B.n523 B.n268 10.6151
R888 B.n524 B.n523 10.6151
R889 B.n525 B.n524 10.6151
R890 B.n525 B.n259 10.6151
R891 B.n535 B.n259 10.6151
R892 B.n536 B.n535 10.6151
R893 B.n538 B.n536 10.6151
R894 B.n538 B.n537 10.6151
R895 B.n537 B.n253 10.6151
R896 B.n550 B.n253 10.6151
R897 B.n551 B.n550 10.6151
R898 B.n552 B.n551 10.6151
R899 B.n553 B.n552 10.6151
R900 B.n554 B.n553 10.6151
R901 B.n557 B.n554 10.6151
R902 B.n558 B.n557 10.6151
R903 B.n559 B.n558 10.6151
R904 B.n560 B.n559 10.6151
R905 B.n562 B.n560 10.6151
R906 B.n563 B.n562 10.6151
R907 B.n564 B.n563 10.6151
R908 B.n565 B.n564 10.6151
R909 B.n567 B.n565 10.6151
R910 B.n568 B.n567 10.6151
R911 B.n569 B.n568 10.6151
R912 B.n570 B.n569 10.6151
R913 B.n571 B.n570 10.6151
R914 B.n604 B.n1 10.6151
R915 B.n604 B.n603 10.6151
R916 B.n603 B.n602 10.6151
R917 B.n602 B.n10 10.6151
R918 B.n596 B.n10 10.6151
R919 B.n596 B.n595 10.6151
R920 B.n595 B.n594 10.6151
R921 B.n594 B.n18 10.6151
R922 B.n588 B.n18 10.6151
R923 B.n588 B.n587 10.6151
R924 B.n587 B.n586 10.6151
R925 B.n586 B.n24 10.6151
R926 B.n580 B.n24 10.6151
R927 B.n580 B.n579 10.6151
R928 B.n578 B.n32 10.6151
R929 B.n83 B.n32 10.6151
R930 B.n84 B.n83 10.6151
R931 B.n87 B.n84 10.6151
R932 B.n88 B.n87 10.6151
R933 B.n91 B.n88 10.6151
R934 B.n92 B.n91 10.6151
R935 B.n95 B.n92 10.6151
R936 B.n96 B.n95 10.6151
R937 B.n99 B.n96 10.6151
R938 B.n100 B.n99 10.6151
R939 B.n103 B.n100 10.6151
R940 B.n104 B.n103 10.6151
R941 B.n107 B.n104 10.6151
R942 B.n108 B.n107 10.6151
R943 B.n111 B.n108 10.6151
R944 B.n112 B.n111 10.6151
R945 B.n115 B.n112 10.6151
R946 B.n116 B.n115 10.6151
R947 B.n119 B.n116 10.6151
R948 B.n120 B.n119 10.6151
R949 B.n123 B.n120 10.6151
R950 B.n124 B.n123 10.6151
R951 B.n127 B.n124 10.6151
R952 B.n128 B.n127 10.6151
R953 B.n131 B.n128 10.6151
R954 B.n132 B.n131 10.6151
R955 B.n135 B.n132 10.6151
R956 B.n136 B.n135 10.6151
R957 B.n139 B.n136 10.6151
R958 B.n140 B.n139 10.6151
R959 B.n143 B.n140 10.6151
R960 B.n144 B.n143 10.6151
R961 B.n147 B.n144 10.6151
R962 B.n148 B.n147 10.6151
R963 B.n151 B.n148 10.6151
R964 B.n152 B.n151 10.6151
R965 B.n155 B.n152 10.6151
R966 B.n160 B.n157 10.6151
R967 B.n161 B.n160 10.6151
R968 B.n164 B.n161 10.6151
R969 B.n165 B.n164 10.6151
R970 B.n168 B.n165 10.6151
R971 B.n169 B.n168 10.6151
R972 B.n172 B.n169 10.6151
R973 B.n173 B.n172 10.6151
R974 B.n176 B.n173 10.6151
R975 B.n181 B.n178 10.6151
R976 B.n182 B.n181 10.6151
R977 B.n185 B.n182 10.6151
R978 B.n186 B.n185 10.6151
R979 B.n189 B.n186 10.6151
R980 B.n190 B.n189 10.6151
R981 B.n193 B.n190 10.6151
R982 B.n194 B.n193 10.6151
R983 B.n197 B.n194 10.6151
R984 B.n198 B.n197 10.6151
R985 B.n201 B.n198 10.6151
R986 B.n202 B.n201 10.6151
R987 B.n205 B.n202 10.6151
R988 B.n206 B.n205 10.6151
R989 B.n209 B.n206 10.6151
R990 B.n210 B.n209 10.6151
R991 B.n213 B.n210 10.6151
R992 B.n214 B.n213 10.6151
R993 B.n217 B.n214 10.6151
R994 B.n218 B.n217 10.6151
R995 B.n221 B.n218 10.6151
R996 B.n222 B.n221 10.6151
R997 B.n225 B.n222 10.6151
R998 B.n226 B.n225 10.6151
R999 B.n229 B.n226 10.6151
R1000 B.n230 B.n229 10.6151
R1001 B.n233 B.n230 10.6151
R1002 B.n234 B.n233 10.6151
R1003 B.n237 B.n234 10.6151
R1004 B.n238 B.n237 10.6151
R1005 B.n241 B.n238 10.6151
R1006 B.n242 B.n241 10.6151
R1007 B.n245 B.n242 10.6151
R1008 B.n246 B.n245 10.6151
R1009 B.n249 B.n246 10.6151
R1010 B.n251 B.n249 10.6151
R1011 B.n252 B.n251 10.6151
R1012 B.n572 B.n252 10.6151
R1013 B.n429 B.n327 9.36635
R1014 B.n406 B.n330 9.36635
R1015 B.n156 B.n155 9.36635
R1016 B.n178 B.n177 9.36635
R1017 B.n612 B.n0 8.11757
R1018 B.n612 B.n1 8.11757
R1019 B.n426 B.n327 1.24928
R1020 B.n409 B.n330 1.24928
R1021 B.n157 B.n156 1.24928
R1022 B.n177 B.n176 1.24928
R1023 VP.n0 VP.t1 650.042
R1024 VP.n0 VP.t3 650.016
R1025 VP.n2 VP.t2 629.059
R1026 VP.n3 VP.t0 629.059
R1027 VP.n4 VP.n3 161.3
R1028 VP.n2 VP.n1 161.3
R1029 VP.n1 VP.n0 109.373
R1030 VP.n3 VP.n2 48.2005
R1031 VP.n4 VP.n1 0.189894
R1032 VP VP.n4 0.0516364
R1033 VTAIL.n5 VTAIL.t6 49.4394
R1034 VTAIL.n4 VTAIL.t1 49.4394
R1035 VTAIL.n3 VTAIL.t2 49.4394
R1036 VTAIL.n7 VTAIL.t3 49.4393
R1037 VTAIL.n0 VTAIL.t0 49.4393
R1038 VTAIL.n1 VTAIL.t7 49.4393
R1039 VTAIL.n2 VTAIL.t5 49.4393
R1040 VTAIL.n6 VTAIL.t4 49.4393
R1041 VTAIL.n7 VTAIL.n6 22.6858
R1042 VTAIL.n3 VTAIL.n2 22.6858
R1043 VTAIL.n4 VTAIL.n3 0.707397
R1044 VTAIL.n6 VTAIL.n5 0.707397
R1045 VTAIL.n2 VTAIL.n1 0.707397
R1046 VTAIL.n5 VTAIL.n4 0.470328
R1047 VTAIL.n1 VTAIL.n0 0.470328
R1048 VTAIL VTAIL.n0 0.412138
R1049 VTAIL VTAIL.n7 0.295759
R1050 VDD1 VDD1.n1 100.314
R1051 VDD1 VDD1.n0 64.4005
R1052 VDD1.n0 VDD1.t2 1.77628
R1053 VDD1.n0 VDD1.t0 1.77628
R1054 VDD1.n1 VDD1.t1 1.77628
R1055 VDD1.n1 VDD1.t3 1.77628
R1056 VN.n0 VN.t0 650.042
R1057 VN.n1 VN.t1 650.042
R1058 VN.n0 VN.t2 650.016
R1059 VN.n1 VN.t3 650.016
R1060 VN VN.n1 109.754
R1061 VN VN.n0 70.265
R1062 VDD2.n2 VDD2.n0 99.7898
R1063 VDD2.n2 VDD2.n1 64.3423
R1064 VDD2.n1 VDD2.t0 1.77628
R1065 VDD2.n1 VDD2.t2 1.77628
R1066 VDD2.n0 VDD2.t3 1.77628
R1067 VDD2.n0 VDD2.t1 1.77628
R1068 VDD2 VDD2.n2 0.0586897
C0 VDD1 VN 0.147197f
C1 VDD1 VTAIL 7.313519f
C2 VP VDD2 0.260147f
C3 VN VP 4.51387f
C4 VN VDD2 2.4915f
C5 VTAIL VP 2.09031f
C6 VDD1 VP 2.60424f
C7 VTAIL VDD2 7.35358f
C8 VDD1 VDD2 0.521314f
C9 VN VTAIL 2.0762f
C10 VDD2 B 2.520195f
C11 VDD1 B 6.21484f
C12 VTAIL B 8.157932f
C13 VN B 7.984049f
C14 VP B 4.392555f
C15 VDD2.t3 B 0.263533f
C16 VDD2.t1 B 0.263533f
C17 VDD2.n0 B 2.92475f
C18 VDD2.t0 B 0.263533f
C19 VDD2.t2 B 0.263533f
C20 VDD2.n1 B 2.33979f
C21 VDD2.n2 B 3.50676f
C22 VN.t0 B 0.867223f
C23 VN.t2 B 0.867207f
C24 VN.n0 B 0.67785f
C25 VN.t1 B 0.867223f
C26 VN.t3 B 0.867207f
C27 VN.n1 B 1.43801f
C28 VDD1.t2 B 0.260624f
C29 VDD1.t0 B 0.260624f
C30 VDD1.n0 B 2.31427f
C31 VDD1.t1 B 0.260624f
C32 VDD1.t3 B 0.260624f
C33 VDD1.n1 B 2.91957f
C34 VTAIL.t0 B 1.67751f
C35 VTAIL.n0 B 0.273334f
C36 VTAIL.t7 B 1.67751f
C37 VTAIL.n1 B 0.289922f
C38 VTAIL.t5 B 1.67751f
C39 VTAIL.n2 B 1.08006f
C40 VTAIL.t2 B 1.67752f
C41 VTAIL.n3 B 1.08005f
C42 VTAIL.t1 B 1.67752f
C43 VTAIL.n4 B 0.289911f
C44 VTAIL.t6 B 1.67752f
C45 VTAIL.n5 B 0.289911f
C46 VTAIL.t4 B 1.67751f
C47 VTAIL.n6 B 1.08006f
C48 VTAIL.t3 B 1.67751f
C49 VTAIL.n7 B 1.05693f
C50 VP.t3 B 0.884229f
C51 VP.t1 B 0.884245f
C52 VP.n0 B 1.44824f
C53 VP.n1 B 3.4572f
C54 VP.t2 B 0.872719f
C55 VP.n2 B 0.357017f
C56 VP.t0 B 0.872719f
C57 VP.n3 B 0.357017f
C58 VP.n4 B 0.043342f
.ends

