* NGSPICE file created from diff_pair_sample_1468.ext - technology: sky130A

.subckt diff_pair_sample_1468 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=5.1207 pd=27.04 as=0 ps=0 w=13.13 l=0.79
X1 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=5.1207 pd=27.04 as=0 ps=0 w=13.13 l=0.79
X2 VTAIL.t18 VP.t0 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.16645 pd=13.46 as=2.16645 ps=13.46 w=13.13 l=0.79
X3 VTAIL.t19 VN.t0 VDD2.t9 B.t6 sky130_fd_pr__nfet_01v8 ad=2.16645 pd=13.46 as=2.16645 ps=13.46 w=13.13 l=0.79
X4 VDD1.t2 VP.t1 VTAIL.t17 B.t5 sky130_fd_pr__nfet_01v8 ad=5.1207 pd=27.04 as=2.16645 ps=13.46 w=13.13 l=0.79
X5 VTAIL.t16 VP.t2 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.16645 pd=13.46 as=2.16645 ps=13.46 w=13.13 l=0.79
X6 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=5.1207 pd=27.04 as=0 ps=0 w=13.13 l=0.79
X7 VTAIL.t15 VP.t3 VDD1.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=2.16645 pd=13.46 as=2.16645 ps=13.46 w=13.13 l=0.79
X8 VDD1.t5 VP.t4 VTAIL.t14 B.t8 sky130_fd_pr__nfet_01v8 ad=5.1207 pd=27.04 as=2.16645 ps=13.46 w=13.13 l=0.79
X9 VDD2.t8 VN.t1 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.1207 pd=27.04 as=2.16645 ps=13.46 w=13.13 l=0.79
X10 VDD2.t7 VN.t2 VTAIL.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=5.1207 pd=27.04 as=2.16645 ps=13.46 w=13.13 l=0.79
X11 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.1207 pd=27.04 as=0 ps=0 w=13.13 l=0.79
X12 VTAIL.t8 VN.t3 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=2.16645 pd=13.46 as=2.16645 ps=13.46 w=13.13 l=0.79
X13 VTAIL.t7 VN.t4 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.16645 pd=13.46 as=2.16645 ps=13.46 w=13.13 l=0.79
X14 VDD2.t4 VN.t5 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.16645 pd=13.46 as=5.1207 ps=27.04 w=13.13 l=0.79
X15 VTAIL.t3 VN.t6 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=2.16645 pd=13.46 as=2.16645 ps=13.46 w=13.13 l=0.79
X16 VDD2.t2 VN.t7 VTAIL.t4 B.t9 sky130_fd_pr__nfet_01v8 ad=2.16645 pd=13.46 as=5.1207 ps=27.04 w=13.13 l=0.79
X17 VDD2.t1 VN.t8 VTAIL.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.16645 pd=13.46 as=2.16645 ps=13.46 w=13.13 l=0.79
X18 VDD1.t0 VP.t5 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=2.16645 pd=13.46 as=5.1207 ps=27.04 w=13.13 l=0.79
X19 VDD1.t3 VP.t6 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=2.16645 pd=13.46 as=2.16645 ps=13.46 w=13.13 l=0.79
X20 VDD2.t0 VN.t9 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.16645 pd=13.46 as=2.16645 ps=13.46 w=13.13 l=0.79
X21 VDD1.t8 VP.t7 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=2.16645 pd=13.46 as=2.16645 ps=13.46 w=13.13 l=0.79
X22 VDD1.t7 VP.t8 VTAIL.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.16645 pd=13.46 as=5.1207 ps=27.04 w=13.13 l=0.79
X23 VTAIL.t9 VP.t9 VDD1.t9 B.t6 sky130_fd_pr__nfet_01v8 ad=2.16645 pd=13.46 as=2.16645 ps=13.46 w=13.13 l=0.79
R0 B.n380 B.t21 602.533
R1 B.n386 B.t10 602.533
R2 B.n108 B.t14 602.533
R3 B.n105 B.t18 602.533
R4 B.n732 B.n731 585
R5 B.n733 B.n732 585
R6 B.n303 B.n104 585
R7 B.n302 B.n301 585
R8 B.n300 B.n299 585
R9 B.n298 B.n297 585
R10 B.n296 B.n295 585
R11 B.n294 B.n293 585
R12 B.n292 B.n291 585
R13 B.n290 B.n289 585
R14 B.n288 B.n287 585
R15 B.n286 B.n285 585
R16 B.n284 B.n283 585
R17 B.n282 B.n281 585
R18 B.n280 B.n279 585
R19 B.n278 B.n277 585
R20 B.n276 B.n275 585
R21 B.n274 B.n273 585
R22 B.n272 B.n271 585
R23 B.n270 B.n269 585
R24 B.n268 B.n267 585
R25 B.n266 B.n265 585
R26 B.n264 B.n263 585
R27 B.n262 B.n261 585
R28 B.n260 B.n259 585
R29 B.n258 B.n257 585
R30 B.n256 B.n255 585
R31 B.n254 B.n253 585
R32 B.n252 B.n251 585
R33 B.n250 B.n249 585
R34 B.n248 B.n247 585
R35 B.n246 B.n245 585
R36 B.n244 B.n243 585
R37 B.n242 B.n241 585
R38 B.n240 B.n239 585
R39 B.n238 B.n237 585
R40 B.n236 B.n235 585
R41 B.n234 B.n233 585
R42 B.n232 B.n231 585
R43 B.n230 B.n229 585
R44 B.n228 B.n227 585
R45 B.n226 B.n225 585
R46 B.n224 B.n223 585
R47 B.n222 B.n221 585
R48 B.n220 B.n219 585
R49 B.n218 B.n217 585
R50 B.n216 B.n215 585
R51 B.n214 B.n213 585
R52 B.n212 B.n211 585
R53 B.n210 B.n209 585
R54 B.n208 B.n207 585
R55 B.n206 B.n205 585
R56 B.n204 B.n203 585
R57 B.n202 B.n201 585
R58 B.n200 B.n199 585
R59 B.n197 B.n196 585
R60 B.n195 B.n194 585
R61 B.n193 B.n192 585
R62 B.n191 B.n190 585
R63 B.n189 B.n188 585
R64 B.n187 B.n186 585
R65 B.n185 B.n184 585
R66 B.n183 B.n182 585
R67 B.n181 B.n180 585
R68 B.n179 B.n178 585
R69 B.n177 B.n176 585
R70 B.n175 B.n174 585
R71 B.n173 B.n172 585
R72 B.n171 B.n170 585
R73 B.n169 B.n168 585
R74 B.n167 B.n166 585
R75 B.n165 B.n164 585
R76 B.n163 B.n162 585
R77 B.n161 B.n160 585
R78 B.n159 B.n158 585
R79 B.n157 B.n156 585
R80 B.n155 B.n154 585
R81 B.n153 B.n152 585
R82 B.n151 B.n150 585
R83 B.n149 B.n148 585
R84 B.n147 B.n146 585
R85 B.n145 B.n144 585
R86 B.n143 B.n142 585
R87 B.n141 B.n140 585
R88 B.n139 B.n138 585
R89 B.n137 B.n136 585
R90 B.n135 B.n134 585
R91 B.n133 B.n132 585
R92 B.n131 B.n130 585
R93 B.n129 B.n128 585
R94 B.n127 B.n126 585
R95 B.n125 B.n124 585
R96 B.n123 B.n122 585
R97 B.n121 B.n120 585
R98 B.n119 B.n118 585
R99 B.n117 B.n116 585
R100 B.n115 B.n114 585
R101 B.n113 B.n112 585
R102 B.n111 B.n110 585
R103 B.n53 B.n52 585
R104 B.n730 B.n54 585
R105 B.n734 B.n54 585
R106 B.n729 B.n728 585
R107 B.n728 B.n50 585
R108 B.n727 B.n49 585
R109 B.n740 B.n49 585
R110 B.n726 B.n48 585
R111 B.n741 B.n48 585
R112 B.n725 B.n47 585
R113 B.n742 B.n47 585
R114 B.n724 B.n723 585
R115 B.n723 B.n46 585
R116 B.n722 B.n42 585
R117 B.n748 B.n42 585
R118 B.n721 B.n41 585
R119 B.n749 B.n41 585
R120 B.n720 B.n40 585
R121 B.n750 B.n40 585
R122 B.n719 B.n718 585
R123 B.n718 B.n36 585
R124 B.n717 B.n35 585
R125 B.n756 B.n35 585
R126 B.n716 B.n34 585
R127 B.n757 B.n34 585
R128 B.n715 B.n33 585
R129 B.n758 B.n33 585
R130 B.n714 B.n713 585
R131 B.n713 B.n29 585
R132 B.n712 B.n28 585
R133 B.n764 B.n28 585
R134 B.n711 B.n27 585
R135 B.n765 B.n27 585
R136 B.n710 B.n26 585
R137 B.n766 B.n26 585
R138 B.n709 B.n708 585
R139 B.n708 B.n22 585
R140 B.n707 B.n21 585
R141 B.n772 B.n21 585
R142 B.n706 B.n20 585
R143 B.n773 B.n20 585
R144 B.n705 B.n19 585
R145 B.n774 B.n19 585
R146 B.n704 B.n703 585
R147 B.n703 B.n18 585
R148 B.n702 B.n14 585
R149 B.n780 B.n14 585
R150 B.n701 B.n13 585
R151 B.n781 B.n13 585
R152 B.n700 B.n12 585
R153 B.n782 B.n12 585
R154 B.n699 B.n698 585
R155 B.n698 B.n8 585
R156 B.n697 B.n7 585
R157 B.n788 B.n7 585
R158 B.n696 B.n6 585
R159 B.n789 B.n6 585
R160 B.n695 B.n5 585
R161 B.n790 B.n5 585
R162 B.n694 B.n693 585
R163 B.n693 B.n4 585
R164 B.n692 B.n304 585
R165 B.n692 B.n691 585
R166 B.n682 B.n305 585
R167 B.n306 B.n305 585
R168 B.n684 B.n683 585
R169 B.n685 B.n684 585
R170 B.n681 B.n311 585
R171 B.n311 B.n310 585
R172 B.n680 B.n679 585
R173 B.n679 B.n678 585
R174 B.n313 B.n312 585
R175 B.n671 B.n313 585
R176 B.n670 B.n669 585
R177 B.n672 B.n670 585
R178 B.n668 B.n318 585
R179 B.n318 B.n317 585
R180 B.n667 B.n666 585
R181 B.n666 B.n665 585
R182 B.n320 B.n319 585
R183 B.n321 B.n320 585
R184 B.n658 B.n657 585
R185 B.n659 B.n658 585
R186 B.n656 B.n326 585
R187 B.n326 B.n325 585
R188 B.n655 B.n654 585
R189 B.n654 B.n653 585
R190 B.n328 B.n327 585
R191 B.n329 B.n328 585
R192 B.n646 B.n645 585
R193 B.n647 B.n646 585
R194 B.n644 B.n333 585
R195 B.n337 B.n333 585
R196 B.n643 B.n642 585
R197 B.n642 B.n641 585
R198 B.n335 B.n334 585
R199 B.n336 B.n335 585
R200 B.n634 B.n633 585
R201 B.n635 B.n634 585
R202 B.n632 B.n342 585
R203 B.n342 B.n341 585
R204 B.n631 B.n630 585
R205 B.n630 B.n629 585
R206 B.n344 B.n343 585
R207 B.n622 B.n344 585
R208 B.n621 B.n620 585
R209 B.n623 B.n621 585
R210 B.n619 B.n349 585
R211 B.n349 B.n348 585
R212 B.n618 B.n617 585
R213 B.n617 B.n616 585
R214 B.n351 B.n350 585
R215 B.n352 B.n351 585
R216 B.n609 B.n608 585
R217 B.n610 B.n609 585
R218 B.n355 B.n354 585
R219 B.n413 B.n412 585
R220 B.n414 B.n410 585
R221 B.n410 B.n356 585
R222 B.n416 B.n415 585
R223 B.n418 B.n409 585
R224 B.n421 B.n420 585
R225 B.n422 B.n408 585
R226 B.n424 B.n423 585
R227 B.n426 B.n407 585
R228 B.n429 B.n428 585
R229 B.n430 B.n406 585
R230 B.n432 B.n431 585
R231 B.n434 B.n405 585
R232 B.n437 B.n436 585
R233 B.n438 B.n404 585
R234 B.n440 B.n439 585
R235 B.n442 B.n403 585
R236 B.n445 B.n444 585
R237 B.n446 B.n402 585
R238 B.n448 B.n447 585
R239 B.n450 B.n401 585
R240 B.n453 B.n452 585
R241 B.n454 B.n400 585
R242 B.n456 B.n455 585
R243 B.n458 B.n399 585
R244 B.n461 B.n460 585
R245 B.n462 B.n398 585
R246 B.n464 B.n463 585
R247 B.n466 B.n397 585
R248 B.n469 B.n468 585
R249 B.n470 B.n396 585
R250 B.n472 B.n471 585
R251 B.n474 B.n395 585
R252 B.n477 B.n476 585
R253 B.n478 B.n394 585
R254 B.n480 B.n479 585
R255 B.n482 B.n393 585
R256 B.n485 B.n484 585
R257 B.n486 B.n392 585
R258 B.n488 B.n487 585
R259 B.n490 B.n391 585
R260 B.n493 B.n492 585
R261 B.n494 B.n390 585
R262 B.n496 B.n495 585
R263 B.n498 B.n389 585
R264 B.n501 B.n500 585
R265 B.n502 B.n385 585
R266 B.n504 B.n503 585
R267 B.n506 B.n384 585
R268 B.n509 B.n508 585
R269 B.n510 B.n383 585
R270 B.n512 B.n511 585
R271 B.n514 B.n382 585
R272 B.n517 B.n516 585
R273 B.n519 B.n379 585
R274 B.n521 B.n520 585
R275 B.n523 B.n378 585
R276 B.n526 B.n525 585
R277 B.n527 B.n377 585
R278 B.n529 B.n528 585
R279 B.n531 B.n376 585
R280 B.n534 B.n533 585
R281 B.n535 B.n375 585
R282 B.n537 B.n536 585
R283 B.n539 B.n374 585
R284 B.n542 B.n541 585
R285 B.n543 B.n373 585
R286 B.n545 B.n544 585
R287 B.n547 B.n372 585
R288 B.n550 B.n549 585
R289 B.n551 B.n371 585
R290 B.n553 B.n552 585
R291 B.n555 B.n370 585
R292 B.n558 B.n557 585
R293 B.n559 B.n369 585
R294 B.n561 B.n560 585
R295 B.n563 B.n368 585
R296 B.n566 B.n565 585
R297 B.n567 B.n367 585
R298 B.n569 B.n568 585
R299 B.n571 B.n366 585
R300 B.n574 B.n573 585
R301 B.n575 B.n365 585
R302 B.n577 B.n576 585
R303 B.n579 B.n364 585
R304 B.n582 B.n581 585
R305 B.n583 B.n363 585
R306 B.n585 B.n584 585
R307 B.n587 B.n362 585
R308 B.n590 B.n589 585
R309 B.n591 B.n361 585
R310 B.n593 B.n592 585
R311 B.n595 B.n360 585
R312 B.n598 B.n597 585
R313 B.n599 B.n359 585
R314 B.n601 B.n600 585
R315 B.n603 B.n358 585
R316 B.n606 B.n605 585
R317 B.n607 B.n357 585
R318 B.n612 B.n611 585
R319 B.n611 B.n610 585
R320 B.n613 B.n353 585
R321 B.n353 B.n352 585
R322 B.n615 B.n614 585
R323 B.n616 B.n615 585
R324 B.n347 B.n346 585
R325 B.n348 B.n347 585
R326 B.n625 B.n624 585
R327 B.n624 B.n623 585
R328 B.n626 B.n345 585
R329 B.n622 B.n345 585
R330 B.n628 B.n627 585
R331 B.n629 B.n628 585
R332 B.n340 B.n339 585
R333 B.n341 B.n340 585
R334 B.n637 B.n636 585
R335 B.n636 B.n635 585
R336 B.n638 B.n338 585
R337 B.n338 B.n336 585
R338 B.n640 B.n639 585
R339 B.n641 B.n640 585
R340 B.n332 B.n331 585
R341 B.n337 B.n332 585
R342 B.n649 B.n648 585
R343 B.n648 B.n647 585
R344 B.n650 B.n330 585
R345 B.n330 B.n329 585
R346 B.n652 B.n651 585
R347 B.n653 B.n652 585
R348 B.n324 B.n323 585
R349 B.n325 B.n324 585
R350 B.n661 B.n660 585
R351 B.n660 B.n659 585
R352 B.n662 B.n322 585
R353 B.n322 B.n321 585
R354 B.n664 B.n663 585
R355 B.n665 B.n664 585
R356 B.n316 B.n315 585
R357 B.n317 B.n316 585
R358 B.n674 B.n673 585
R359 B.n673 B.n672 585
R360 B.n675 B.n314 585
R361 B.n671 B.n314 585
R362 B.n677 B.n676 585
R363 B.n678 B.n677 585
R364 B.n309 B.n308 585
R365 B.n310 B.n309 585
R366 B.n687 B.n686 585
R367 B.n686 B.n685 585
R368 B.n688 B.n307 585
R369 B.n307 B.n306 585
R370 B.n690 B.n689 585
R371 B.n691 B.n690 585
R372 B.n2 B.n0 585
R373 B.n4 B.n2 585
R374 B.n3 B.n1 585
R375 B.n789 B.n3 585
R376 B.n787 B.n786 585
R377 B.n788 B.n787 585
R378 B.n785 B.n9 585
R379 B.n9 B.n8 585
R380 B.n784 B.n783 585
R381 B.n783 B.n782 585
R382 B.n11 B.n10 585
R383 B.n781 B.n11 585
R384 B.n779 B.n778 585
R385 B.n780 B.n779 585
R386 B.n777 B.n15 585
R387 B.n18 B.n15 585
R388 B.n776 B.n775 585
R389 B.n775 B.n774 585
R390 B.n17 B.n16 585
R391 B.n773 B.n17 585
R392 B.n771 B.n770 585
R393 B.n772 B.n771 585
R394 B.n769 B.n23 585
R395 B.n23 B.n22 585
R396 B.n768 B.n767 585
R397 B.n767 B.n766 585
R398 B.n25 B.n24 585
R399 B.n765 B.n25 585
R400 B.n763 B.n762 585
R401 B.n764 B.n763 585
R402 B.n761 B.n30 585
R403 B.n30 B.n29 585
R404 B.n760 B.n759 585
R405 B.n759 B.n758 585
R406 B.n32 B.n31 585
R407 B.n757 B.n32 585
R408 B.n755 B.n754 585
R409 B.n756 B.n755 585
R410 B.n753 B.n37 585
R411 B.n37 B.n36 585
R412 B.n752 B.n751 585
R413 B.n751 B.n750 585
R414 B.n39 B.n38 585
R415 B.n749 B.n39 585
R416 B.n747 B.n746 585
R417 B.n748 B.n747 585
R418 B.n745 B.n43 585
R419 B.n46 B.n43 585
R420 B.n744 B.n743 585
R421 B.n743 B.n742 585
R422 B.n45 B.n44 585
R423 B.n741 B.n45 585
R424 B.n739 B.n738 585
R425 B.n740 B.n739 585
R426 B.n737 B.n51 585
R427 B.n51 B.n50 585
R428 B.n736 B.n735 585
R429 B.n735 B.n734 585
R430 B.n792 B.n791 585
R431 B.n791 B.n790 585
R432 B.n611 B.n355 516.524
R433 B.n735 B.n53 516.524
R434 B.n609 B.n357 516.524
R435 B.n732 B.n54 516.524
R436 B.n733 B.n103 256.663
R437 B.n733 B.n102 256.663
R438 B.n733 B.n101 256.663
R439 B.n733 B.n100 256.663
R440 B.n733 B.n99 256.663
R441 B.n733 B.n98 256.663
R442 B.n733 B.n97 256.663
R443 B.n733 B.n96 256.663
R444 B.n733 B.n95 256.663
R445 B.n733 B.n94 256.663
R446 B.n733 B.n93 256.663
R447 B.n733 B.n92 256.663
R448 B.n733 B.n91 256.663
R449 B.n733 B.n90 256.663
R450 B.n733 B.n89 256.663
R451 B.n733 B.n88 256.663
R452 B.n733 B.n87 256.663
R453 B.n733 B.n86 256.663
R454 B.n733 B.n85 256.663
R455 B.n733 B.n84 256.663
R456 B.n733 B.n83 256.663
R457 B.n733 B.n82 256.663
R458 B.n733 B.n81 256.663
R459 B.n733 B.n80 256.663
R460 B.n733 B.n79 256.663
R461 B.n733 B.n78 256.663
R462 B.n733 B.n77 256.663
R463 B.n733 B.n76 256.663
R464 B.n733 B.n75 256.663
R465 B.n733 B.n74 256.663
R466 B.n733 B.n73 256.663
R467 B.n733 B.n72 256.663
R468 B.n733 B.n71 256.663
R469 B.n733 B.n70 256.663
R470 B.n733 B.n69 256.663
R471 B.n733 B.n68 256.663
R472 B.n733 B.n67 256.663
R473 B.n733 B.n66 256.663
R474 B.n733 B.n65 256.663
R475 B.n733 B.n64 256.663
R476 B.n733 B.n63 256.663
R477 B.n733 B.n62 256.663
R478 B.n733 B.n61 256.663
R479 B.n733 B.n60 256.663
R480 B.n733 B.n59 256.663
R481 B.n733 B.n58 256.663
R482 B.n733 B.n57 256.663
R483 B.n733 B.n56 256.663
R484 B.n733 B.n55 256.663
R485 B.n411 B.n356 256.663
R486 B.n417 B.n356 256.663
R487 B.n419 B.n356 256.663
R488 B.n425 B.n356 256.663
R489 B.n427 B.n356 256.663
R490 B.n433 B.n356 256.663
R491 B.n435 B.n356 256.663
R492 B.n441 B.n356 256.663
R493 B.n443 B.n356 256.663
R494 B.n449 B.n356 256.663
R495 B.n451 B.n356 256.663
R496 B.n457 B.n356 256.663
R497 B.n459 B.n356 256.663
R498 B.n465 B.n356 256.663
R499 B.n467 B.n356 256.663
R500 B.n473 B.n356 256.663
R501 B.n475 B.n356 256.663
R502 B.n481 B.n356 256.663
R503 B.n483 B.n356 256.663
R504 B.n489 B.n356 256.663
R505 B.n491 B.n356 256.663
R506 B.n497 B.n356 256.663
R507 B.n499 B.n356 256.663
R508 B.n505 B.n356 256.663
R509 B.n507 B.n356 256.663
R510 B.n513 B.n356 256.663
R511 B.n515 B.n356 256.663
R512 B.n522 B.n356 256.663
R513 B.n524 B.n356 256.663
R514 B.n530 B.n356 256.663
R515 B.n532 B.n356 256.663
R516 B.n538 B.n356 256.663
R517 B.n540 B.n356 256.663
R518 B.n546 B.n356 256.663
R519 B.n548 B.n356 256.663
R520 B.n554 B.n356 256.663
R521 B.n556 B.n356 256.663
R522 B.n562 B.n356 256.663
R523 B.n564 B.n356 256.663
R524 B.n570 B.n356 256.663
R525 B.n572 B.n356 256.663
R526 B.n578 B.n356 256.663
R527 B.n580 B.n356 256.663
R528 B.n586 B.n356 256.663
R529 B.n588 B.n356 256.663
R530 B.n594 B.n356 256.663
R531 B.n596 B.n356 256.663
R532 B.n602 B.n356 256.663
R533 B.n604 B.n356 256.663
R534 B.n611 B.n353 163.367
R535 B.n615 B.n353 163.367
R536 B.n615 B.n347 163.367
R537 B.n624 B.n347 163.367
R538 B.n624 B.n345 163.367
R539 B.n628 B.n345 163.367
R540 B.n628 B.n340 163.367
R541 B.n636 B.n340 163.367
R542 B.n636 B.n338 163.367
R543 B.n640 B.n338 163.367
R544 B.n640 B.n332 163.367
R545 B.n648 B.n332 163.367
R546 B.n648 B.n330 163.367
R547 B.n652 B.n330 163.367
R548 B.n652 B.n324 163.367
R549 B.n660 B.n324 163.367
R550 B.n660 B.n322 163.367
R551 B.n664 B.n322 163.367
R552 B.n664 B.n316 163.367
R553 B.n673 B.n316 163.367
R554 B.n673 B.n314 163.367
R555 B.n677 B.n314 163.367
R556 B.n677 B.n309 163.367
R557 B.n686 B.n309 163.367
R558 B.n686 B.n307 163.367
R559 B.n690 B.n307 163.367
R560 B.n690 B.n2 163.367
R561 B.n791 B.n2 163.367
R562 B.n791 B.n3 163.367
R563 B.n787 B.n3 163.367
R564 B.n787 B.n9 163.367
R565 B.n783 B.n9 163.367
R566 B.n783 B.n11 163.367
R567 B.n779 B.n11 163.367
R568 B.n779 B.n15 163.367
R569 B.n775 B.n15 163.367
R570 B.n775 B.n17 163.367
R571 B.n771 B.n17 163.367
R572 B.n771 B.n23 163.367
R573 B.n767 B.n23 163.367
R574 B.n767 B.n25 163.367
R575 B.n763 B.n25 163.367
R576 B.n763 B.n30 163.367
R577 B.n759 B.n30 163.367
R578 B.n759 B.n32 163.367
R579 B.n755 B.n32 163.367
R580 B.n755 B.n37 163.367
R581 B.n751 B.n37 163.367
R582 B.n751 B.n39 163.367
R583 B.n747 B.n39 163.367
R584 B.n747 B.n43 163.367
R585 B.n743 B.n43 163.367
R586 B.n743 B.n45 163.367
R587 B.n739 B.n45 163.367
R588 B.n739 B.n51 163.367
R589 B.n735 B.n51 163.367
R590 B.n412 B.n410 163.367
R591 B.n416 B.n410 163.367
R592 B.n420 B.n418 163.367
R593 B.n424 B.n408 163.367
R594 B.n428 B.n426 163.367
R595 B.n432 B.n406 163.367
R596 B.n436 B.n434 163.367
R597 B.n440 B.n404 163.367
R598 B.n444 B.n442 163.367
R599 B.n448 B.n402 163.367
R600 B.n452 B.n450 163.367
R601 B.n456 B.n400 163.367
R602 B.n460 B.n458 163.367
R603 B.n464 B.n398 163.367
R604 B.n468 B.n466 163.367
R605 B.n472 B.n396 163.367
R606 B.n476 B.n474 163.367
R607 B.n480 B.n394 163.367
R608 B.n484 B.n482 163.367
R609 B.n488 B.n392 163.367
R610 B.n492 B.n490 163.367
R611 B.n496 B.n390 163.367
R612 B.n500 B.n498 163.367
R613 B.n504 B.n385 163.367
R614 B.n508 B.n506 163.367
R615 B.n512 B.n383 163.367
R616 B.n516 B.n514 163.367
R617 B.n521 B.n379 163.367
R618 B.n525 B.n523 163.367
R619 B.n529 B.n377 163.367
R620 B.n533 B.n531 163.367
R621 B.n537 B.n375 163.367
R622 B.n541 B.n539 163.367
R623 B.n545 B.n373 163.367
R624 B.n549 B.n547 163.367
R625 B.n553 B.n371 163.367
R626 B.n557 B.n555 163.367
R627 B.n561 B.n369 163.367
R628 B.n565 B.n563 163.367
R629 B.n569 B.n367 163.367
R630 B.n573 B.n571 163.367
R631 B.n577 B.n365 163.367
R632 B.n581 B.n579 163.367
R633 B.n585 B.n363 163.367
R634 B.n589 B.n587 163.367
R635 B.n593 B.n361 163.367
R636 B.n597 B.n595 163.367
R637 B.n601 B.n359 163.367
R638 B.n605 B.n603 163.367
R639 B.n609 B.n351 163.367
R640 B.n617 B.n351 163.367
R641 B.n617 B.n349 163.367
R642 B.n621 B.n349 163.367
R643 B.n621 B.n344 163.367
R644 B.n630 B.n344 163.367
R645 B.n630 B.n342 163.367
R646 B.n634 B.n342 163.367
R647 B.n634 B.n335 163.367
R648 B.n642 B.n335 163.367
R649 B.n642 B.n333 163.367
R650 B.n646 B.n333 163.367
R651 B.n646 B.n328 163.367
R652 B.n654 B.n328 163.367
R653 B.n654 B.n326 163.367
R654 B.n658 B.n326 163.367
R655 B.n658 B.n320 163.367
R656 B.n666 B.n320 163.367
R657 B.n666 B.n318 163.367
R658 B.n670 B.n318 163.367
R659 B.n670 B.n313 163.367
R660 B.n679 B.n313 163.367
R661 B.n679 B.n311 163.367
R662 B.n684 B.n311 163.367
R663 B.n684 B.n305 163.367
R664 B.n692 B.n305 163.367
R665 B.n693 B.n692 163.367
R666 B.n693 B.n5 163.367
R667 B.n6 B.n5 163.367
R668 B.n7 B.n6 163.367
R669 B.n698 B.n7 163.367
R670 B.n698 B.n12 163.367
R671 B.n13 B.n12 163.367
R672 B.n14 B.n13 163.367
R673 B.n703 B.n14 163.367
R674 B.n703 B.n19 163.367
R675 B.n20 B.n19 163.367
R676 B.n21 B.n20 163.367
R677 B.n708 B.n21 163.367
R678 B.n708 B.n26 163.367
R679 B.n27 B.n26 163.367
R680 B.n28 B.n27 163.367
R681 B.n713 B.n28 163.367
R682 B.n713 B.n33 163.367
R683 B.n34 B.n33 163.367
R684 B.n35 B.n34 163.367
R685 B.n718 B.n35 163.367
R686 B.n718 B.n40 163.367
R687 B.n41 B.n40 163.367
R688 B.n42 B.n41 163.367
R689 B.n723 B.n42 163.367
R690 B.n723 B.n47 163.367
R691 B.n48 B.n47 163.367
R692 B.n49 B.n48 163.367
R693 B.n728 B.n49 163.367
R694 B.n728 B.n54 163.367
R695 B.n112 B.n111 163.367
R696 B.n116 B.n115 163.367
R697 B.n120 B.n119 163.367
R698 B.n124 B.n123 163.367
R699 B.n128 B.n127 163.367
R700 B.n132 B.n131 163.367
R701 B.n136 B.n135 163.367
R702 B.n140 B.n139 163.367
R703 B.n144 B.n143 163.367
R704 B.n148 B.n147 163.367
R705 B.n152 B.n151 163.367
R706 B.n156 B.n155 163.367
R707 B.n160 B.n159 163.367
R708 B.n164 B.n163 163.367
R709 B.n168 B.n167 163.367
R710 B.n172 B.n171 163.367
R711 B.n176 B.n175 163.367
R712 B.n180 B.n179 163.367
R713 B.n184 B.n183 163.367
R714 B.n188 B.n187 163.367
R715 B.n192 B.n191 163.367
R716 B.n196 B.n195 163.367
R717 B.n201 B.n200 163.367
R718 B.n205 B.n204 163.367
R719 B.n209 B.n208 163.367
R720 B.n213 B.n212 163.367
R721 B.n217 B.n216 163.367
R722 B.n221 B.n220 163.367
R723 B.n225 B.n224 163.367
R724 B.n229 B.n228 163.367
R725 B.n233 B.n232 163.367
R726 B.n237 B.n236 163.367
R727 B.n241 B.n240 163.367
R728 B.n245 B.n244 163.367
R729 B.n249 B.n248 163.367
R730 B.n253 B.n252 163.367
R731 B.n257 B.n256 163.367
R732 B.n261 B.n260 163.367
R733 B.n265 B.n264 163.367
R734 B.n269 B.n268 163.367
R735 B.n273 B.n272 163.367
R736 B.n277 B.n276 163.367
R737 B.n281 B.n280 163.367
R738 B.n285 B.n284 163.367
R739 B.n289 B.n288 163.367
R740 B.n293 B.n292 163.367
R741 B.n297 B.n296 163.367
R742 B.n301 B.n300 163.367
R743 B.n732 B.n104 163.367
R744 B.n380 B.t23 93.4433
R745 B.n105 B.t19 93.4433
R746 B.n386 B.t13 93.4266
R747 B.n108 B.t16 93.4266
R748 B.n381 B.t22 71.7221
R749 B.n106 B.t20 71.7221
R750 B.n387 B.t12 71.7054
R751 B.n109 B.t17 71.7054
R752 B.n411 B.n355 71.676
R753 B.n417 B.n416 71.676
R754 B.n420 B.n419 71.676
R755 B.n425 B.n424 71.676
R756 B.n428 B.n427 71.676
R757 B.n433 B.n432 71.676
R758 B.n436 B.n435 71.676
R759 B.n441 B.n440 71.676
R760 B.n444 B.n443 71.676
R761 B.n449 B.n448 71.676
R762 B.n452 B.n451 71.676
R763 B.n457 B.n456 71.676
R764 B.n460 B.n459 71.676
R765 B.n465 B.n464 71.676
R766 B.n468 B.n467 71.676
R767 B.n473 B.n472 71.676
R768 B.n476 B.n475 71.676
R769 B.n481 B.n480 71.676
R770 B.n484 B.n483 71.676
R771 B.n489 B.n488 71.676
R772 B.n492 B.n491 71.676
R773 B.n497 B.n496 71.676
R774 B.n500 B.n499 71.676
R775 B.n505 B.n504 71.676
R776 B.n508 B.n507 71.676
R777 B.n513 B.n512 71.676
R778 B.n516 B.n515 71.676
R779 B.n522 B.n521 71.676
R780 B.n525 B.n524 71.676
R781 B.n530 B.n529 71.676
R782 B.n533 B.n532 71.676
R783 B.n538 B.n537 71.676
R784 B.n541 B.n540 71.676
R785 B.n546 B.n545 71.676
R786 B.n549 B.n548 71.676
R787 B.n554 B.n553 71.676
R788 B.n557 B.n556 71.676
R789 B.n562 B.n561 71.676
R790 B.n565 B.n564 71.676
R791 B.n570 B.n569 71.676
R792 B.n573 B.n572 71.676
R793 B.n578 B.n577 71.676
R794 B.n581 B.n580 71.676
R795 B.n586 B.n585 71.676
R796 B.n589 B.n588 71.676
R797 B.n594 B.n593 71.676
R798 B.n597 B.n596 71.676
R799 B.n602 B.n601 71.676
R800 B.n605 B.n604 71.676
R801 B.n55 B.n53 71.676
R802 B.n112 B.n56 71.676
R803 B.n116 B.n57 71.676
R804 B.n120 B.n58 71.676
R805 B.n124 B.n59 71.676
R806 B.n128 B.n60 71.676
R807 B.n132 B.n61 71.676
R808 B.n136 B.n62 71.676
R809 B.n140 B.n63 71.676
R810 B.n144 B.n64 71.676
R811 B.n148 B.n65 71.676
R812 B.n152 B.n66 71.676
R813 B.n156 B.n67 71.676
R814 B.n160 B.n68 71.676
R815 B.n164 B.n69 71.676
R816 B.n168 B.n70 71.676
R817 B.n172 B.n71 71.676
R818 B.n176 B.n72 71.676
R819 B.n180 B.n73 71.676
R820 B.n184 B.n74 71.676
R821 B.n188 B.n75 71.676
R822 B.n192 B.n76 71.676
R823 B.n196 B.n77 71.676
R824 B.n201 B.n78 71.676
R825 B.n205 B.n79 71.676
R826 B.n209 B.n80 71.676
R827 B.n213 B.n81 71.676
R828 B.n217 B.n82 71.676
R829 B.n221 B.n83 71.676
R830 B.n225 B.n84 71.676
R831 B.n229 B.n85 71.676
R832 B.n233 B.n86 71.676
R833 B.n237 B.n87 71.676
R834 B.n241 B.n88 71.676
R835 B.n245 B.n89 71.676
R836 B.n249 B.n90 71.676
R837 B.n253 B.n91 71.676
R838 B.n257 B.n92 71.676
R839 B.n261 B.n93 71.676
R840 B.n265 B.n94 71.676
R841 B.n269 B.n95 71.676
R842 B.n273 B.n96 71.676
R843 B.n277 B.n97 71.676
R844 B.n281 B.n98 71.676
R845 B.n285 B.n99 71.676
R846 B.n289 B.n100 71.676
R847 B.n293 B.n101 71.676
R848 B.n297 B.n102 71.676
R849 B.n301 B.n103 71.676
R850 B.n104 B.n103 71.676
R851 B.n300 B.n102 71.676
R852 B.n296 B.n101 71.676
R853 B.n292 B.n100 71.676
R854 B.n288 B.n99 71.676
R855 B.n284 B.n98 71.676
R856 B.n280 B.n97 71.676
R857 B.n276 B.n96 71.676
R858 B.n272 B.n95 71.676
R859 B.n268 B.n94 71.676
R860 B.n264 B.n93 71.676
R861 B.n260 B.n92 71.676
R862 B.n256 B.n91 71.676
R863 B.n252 B.n90 71.676
R864 B.n248 B.n89 71.676
R865 B.n244 B.n88 71.676
R866 B.n240 B.n87 71.676
R867 B.n236 B.n86 71.676
R868 B.n232 B.n85 71.676
R869 B.n228 B.n84 71.676
R870 B.n224 B.n83 71.676
R871 B.n220 B.n82 71.676
R872 B.n216 B.n81 71.676
R873 B.n212 B.n80 71.676
R874 B.n208 B.n79 71.676
R875 B.n204 B.n78 71.676
R876 B.n200 B.n77 71.676
R877 B.n195 B.n76 71.676
R878 B.n191 B.n75 71.676
R879 B.n187 B.n74 71.676
R880 B.n183 B.n73 71.676
R881 B.n179 B.n72 71.676
R882 B.n175 B.n71 71.676
R883 B.n171 B.n70 71.676
R884 B.n167 B.n69 71.676
R885 B.n163 B.n68 71.676
R886 B.n159 B.n67 71.676
R887 B.n155 B.n66 71.676
R888 B.n151 B.n65 71.676
R889 B.n147 B.n64 71.676
R890 B.n143 B.n63 71.676
R891 B.n139 B.n62 71.676
R892 B.n135 B.n61 71.676
R893 B.n131 B.n60 71.676
R894 B.n127 B.n59 71.676
R895 B.n123 B.n58 71.676
R896 B.n119 B.n57 71.676
R897 B.n115 B.n56 71.676
R898 B.n111 B.n55 71.676
R899 B.n412 B.n411 71.676
R900 B.n418 B.n417 71.676
R901 B.n419 B.n408 71.676
R902 B.n426 B.n425 71.676
R903 B.n427 B.n406 71.676
R904 B.n434 B.n433 71.676
R905 B.n435 B.n404 71.676
R906 B.n442 B.n441 71.676
R907 B.n443 B.n402 71.676
R908 B.n450 B.n449 71.676
R909 B.n451 B.n400 71.676
R910 B.n458 B.n457 71.676
R911 B.n459 B.n398 71.676
R912 B.n466 B.n465 71.676
R913 B.n467 B.n396 71.676
R914 B.n474 B.n473 71.676
R915 B.n475 B.n394 71.676
R916 B.n482 B.n481 71.676
R917 B.n483 B.n392 71.676
R918 B.n490 B.n489 71.676
R919 B.n491 B.n390 71.676
R920 B.n498 B.n497 71.676
R921 B.n499 B.n385 71.676
R922 B.n506 B.n505 71.676
R923 B.n507 B.n383 71.676
R924 B.n514 B.n513 71.676
R925 B.n515 B.n379 71.676
R926 B.n523 B.n522 71.676
R927 B.n524 B.n377 71.676
R928 B.n531 B.n530 71.676
R929 B.n532 B.n375 71.676
R930 B.n539 B.n538 71.676
R931 B.n540 B.n373 71.676
R932 B.n547 B.n546 71.676
R933 B.n548 B.n371 71.676
R934 B.n555 B.n554 71.676
R935 B.n556 B.n369 71.676
R936 B.n563 B.n562 71.676
R937 B.n564 B.n367 71.676
R938 B.n571 B.n570 71.676
R939 B.n572 B.n365 71.676
R940 B.n579 B.n578 71.676
R941 B.n580 B.n363 71.676
R942 B.n587 B.n586 71.676
R943 B.n588 B.n361 71.676
R944 B.n595 B.n594 71.676
R945 B.n596 B.n359 71.676
R946 B.n603 B.n602 71.676
R947 B.n604 B.n357 71.676
R948 B.n610 B.n356 68.7318
R949 B.n734 B.n733 68.7318
R950 B.n518 B.n381 59.5399
R951 B.n388 B.n387 59.5399
R952 B.n198 B.n109 59.5399
R953 B.n107 B.n106 59.5399
R954 B.n610 B.n352 40.6416
R955 B.n616 B.n352 40.6416
R956 B.n616 B.n348 40.6416
R957 B.n623 B.n348 40.6416
R958 B.n623 B.n622 40.6416
R959 B.n629 B.n341 40.6416
R960 B.n635 B.n341 40.6416
R961 B.n635 B.n336 40.6416
R962 B.n641 B.n336 40.6416
R963 B.n641 B.n337 40.6416
R964 B.n647 B.n329 40.6416
R965 B.n653 B.n329 40.6416
R966 B.n659 B.n325 40.6416
R967 B.n659 B.n321 40.6416
R968 B.n665 B.n321 40.6416
R969 B.n672 B.n317 40.6416
R970 B.n672 B.n671 40.6416
R971 B.n678 B.n310 40.6416
R972 B.n685 B.n310 40.6416
R973 B.n691 B.n306 40.6416
R974 B.n691 B.n4 40.6416
R975 B.n790 B.n4 40.6416
R976 B.n790 B.n789 40.6416
R977 B.n789 B.n788 40.6416
R978 B.n788 B.n8 40.6416
R979 B.n782 B.n781 40.6416
R980 B.n781 B.n780 40.6416
R981 B.n774 B.n18 40.6416
R982 B.n774 B.n773 40.6416
R983 B.n772 B.n22 40.6416
R984 B.n766 B.n22 40.6416
R985 B.n766 B.n765 40.6416
R986 B.n764 B.n29 40.6416
R987 B.n758 B.n29 40.6416
R988 B.n757 B.n756 40.6416
R989 B.n756 B.n36 40.6416
R990 B.n750 B.n36 40.6416
R991 B.n750 B.n749 40.6416
R992 B.n749 B.n748 40.6416
R993 B.n742 B.n46 40.6416
R994 B.n742 B.n741 40.6416
R995 B.n741 B.n740 40.6416
R996 B.n740 B.n50 40.6416
R997 B.n734 B.n50 40.6416
R998 B.n629 B.t11 37.6533
R999 B.n748 B.t15 37.6533
R1000 B.n653 B.t4 35.2627
R1001 B.t7 B.n764 35.2627
R1002 B.t0 B.n317 34.0673
R1003 B.n773 B.t2 34.0673
R1004 B.n736 B.n52 33.5615
R1005 B.n731 B.n730 33.5615
R1006 B.n608 B.n607 33.5615
R1007 B.n612 B.n354 33.5615
R1008 B.n685 B.t3 30.4813
R1009 B.n782 B.t8 30.4813
R1010 B.n337 B.t5 23.3094
R1011 B.t9 B.n757 23.3094
R1012 B.n678 B.t6 22.1141
R1013 B.n780 B.t1 22.1141
R1014 B.n381 B.n380 21.7217
R1015 B.n387 B.n386 21.7217
R1016 B.n109 B.n108 21.7217
R1017 B.n106 B.n105 21.7217
R1018 B.n671 B.t6 18.5281
R1019 B.n18 B.t1 18.5281
R1020 B B.n792 18.0485
R1021 B.n647 B.t5 17.3327
R1022 B.n758 B.t9 17.3327
R1023 B.n110 B.n52 10.6151
R1024 B.n113 B.n110 10.6151
R1025 B.n114 B.n113 10.6151
R1026 B.n117 B.n114 10.6151
R1027 B.n118 B.n117 10.6151
R1028 B.n121 B.n118 10.6151
R1029 B.n122 B.n121 10.6151
R1030 B.n125 B.n122 10.6151
R1031 B.n126 B.n125 10.6151
R1032 B.n129 B.n126 10.6151
R1033 B.n130 B.n129 10.6151
R1034 B.n133 B.n130 10.6151
R1035 B.n134 B.n133 10.6151
R1036 B.n137 B.n134 10.6151
R1037 B.n138 B.n137 10.6151
R1038 B.n141 B.n138 10.6151
R1039 B.n142 B.n141 10.6151
R1040 B.n145 B.n142 10.6151
R1041 B.n146 B.n145 10.6151
R1042 B.n149 B.n146 10.6151
R1043 B.n150 B.n149 10.6151
R1044 B.n153 B.n150 10.6151
R1045 B.n154 B.n153 10.6151
R1046 B.n157 B.n154 10.6151
R1047 B.n158 B.n157 10.6151
R1048 B.n161 B.n158 10.6151
R1049 B.n162 B.n161 10.6151
R1050 B.n165 B.n162 10.6151
R1051 B.n166 B.n165 10.6151
R1052 B.n169 B.n166 10.6151
R1053 B.n170 B.n169 10.6151
R1054 B.n173 B.n170 10.6151
R1055 B.n174 B.n173 10.6151
R1056 B.n177 B.n174 10.6151
R1057 B.n178 B.n177 10.6151
R1058 B.n181 B.n178 10.6151
R1059 B.n182 B.n181 10.6151
R1060 B.n185 B.n182 10.6151
R1061 B.n186 B.n185 10.6151
R1062 B.n189 B.n186 10.6151
R1063 B.n190 B.n189 10.6151
R1064 B.n193 B.n190 10.6151
R1065 B.n194 B.n193 10.6151
R1066 B.n197 B.n194 10.6151
R1067 B.n202 B.n199 10.6151
R1068 B.n203 B.n202 10.6151
R1069 B.n206 B.n203 10.6151
R1070 B.n207 B.n206 10.6151
R1071 B.n210 B.n207 10.6151
R1072 B.n211 B.n210 10.6151
R1073 B.n214 B.n211 10.6151
R1074 B.n215 B.n214 10.6151
R1075 B.n219 B.n218 10.6151
R1076 B.n222 B.n219 10.6151
R1077 B.n223 B.n222 10.6151
R1078 B.n226 B.n223 10.6151
R1079 B.n227 B.n226 10.6151
R1080 B.n230 B.n227 10.6151
R1081 B.n231 B.n230 10.6151
R1082 B.n234 B.n231 10.6151
R1083 B.n235 B.n234 10.6151
R1084 B.n238 B.n235 10.6151
R1085 B.n239 B.n238 10.6151
R1086 B.n242 B.n239 10.6151
R1087 B.n243 B.n242 10.6151
R1088 B.n246 B.n243 10.6151
R1089 B.n247 B.n246 10.6151
R1090 B.n250 B.n247 10.6151
R1091 B.n251 B.n250 10.6151
R1092 B.n254 B.n251 10.6151
R1093 B.n255 B.n254 10.6151
R1094 B.n258 B.n255 10.6151
R1095 B.n259 B.n258 10.6151
R1096 B.n262 B.n259 10.6151
R1097 B.n263 B.n262 10.6151
R1098 B.n266 B.n263 10.6151
R1099 B.n267 B.n266 10.6151
R1100 B.n270 B.n267 10.6151
R1101 B.n271 B.n270 10.6151
R1102 B.n274 B.n271 10.6151
R1103 B.n275 B.n274 10.6151
R1104 B.n278 B.n275 10.6151
R1105 B.n279 B.n278 10.6151
R1106 B.n282 B.n279 10.6151
R1107 B.n283 B.n282 10.6151
R1108 B.n286 B.n283 10.6151
R1109 B.n287 B.n286 10.6151
R1110 B.n290 B.n287 10.6151
R1111 B.n291 B.n290 10.6151
R1112 B.n294 B.n291 10.6151
R1113 B.n295 B.n294 10.6151
R1114 B.n298 B.n295 10.6151
R1115 B.n299 B.n298 10.6151
R1116 B.n302 B.n299 10.6151
R1117 B.n303 B.n302 10.6151
R1118 B.n731 B.n303 10.6151
R1119 B.n608 B.n350 10.6151
R1120 B.n618 B.n350 10.6151
R1121 B.n619 B.n618 10.6151
R1122 B.n620 B.n619 10.6151
R1123 B.n620 B.n343 10.6151
R1124 B.n631 B.n343 10.6151
R1125 B.n632 B.n631 10.6151
R1126 B.n633 B.n632 10.6151
R1127 B.n633 B.n334 10.6151
R1128 B.n643 B.n334 10.6151
R1129 B.n644 B.n643 10.6151
R1130 B.n645 B.n644 10.6151
R1131 B.n645 B.n327 10.6151
R1132 B.n655 B.n327 10.6151
R1133 B.n656 B.n655 10.6151
R1134 B.n657 B.n656 10.6151
R1135 B.n657 B.n319 10.6151
R1136 B.n667 B.n319 10.6151
R1137 B.n668 B.n667 10.6151
R1138 B.n669 B.n668 10.6151
R1139 B.n669 B.n312 10.6151
R1140 B.n680 B.n312 10.6151
R1141 B.n681 B.n680 10.6151
R1142 B.n683 B.n681 10.6151
R1143 B.n683 B.n682 10.6151
R1144 B.n682 B.n304 10.6151
R1145 B.n694 B.n304 10.6151
R1146 B.n695 B.n694 10.6151
R1147 B.n696 B.n695 10.6151
R1148 B.n697 B.n696 10.6151
R1149 B.n699 B.n697 10.6151
R1150 B.n700 B.n699 10.6151
R1151 B.n701 B.n700 10.6151
R1152 B.n702 B.n701 10.6151
R1153 B.n704 B.n702 10.6151
R1154 B.n705 B.n704 10.6151
R1155 B.n706 B.n705 10.6151
R1156 B.n707 B.n706 10.6151
R1157 B.n709 B.n707 10.6151
R1158 B.n710 B.n709 10.6151
R1159 B.n711 B.n710 10.6151
R1160 B.n712 B.n711 10.6151
R1161 B.n714 B.n712 10.6151
R1162 B.n715 B.n714 10.6151
R1163 B.n716 B.n715 10.6151
R1164 B.n717 B.n716 10.6151
R1165 B.n719 B.n717 10.6151
R1166 B.n720 B.n719 10.6151
R1167 B.n721 B.n720 10.6151
R1168 B.n722 B.n721 10.6151
R1169 B.n724 B.n722 10.6151
R1170 B.n725 B.n724 10.6151
R1171 B.n726 B.n725 10.6151
R1172 B.n727 B.n726 10.6151
R1173 B.n729 B.n727 10.6151
R1174 B.n730 B.n729 10.6151
R1175 B.n413 B.n354 10.6151
R1176 B.n414 B.n413 10.6151
R1177 B.n415 B.n414 10.6151
R1178 B.n415 B.n409 10.6151
R1179 B.n421 B.n409 10.6151
R1180 B.n422 B.n421 10.6151
R1181 B.n423 B.n422 10.6151
R1182 B.n423 B.n407 10.6151
R1183 B.n429 B.n407 10.6151
R1184 B.n430 B.n429 10.6151
R1185 B.n431 B.n430 10.6151
R1186 B.n431 B.n405 10.6151
R1187 B.n437 B.n405 10.6151
R1188 B.n438 B.n437 10.6151
R1189 B.n439 B.n438 10.6151
R1190 B.n439 B.n403 10.6151
R1191 B.n445 B.n403 10.6151
R1192 B.n446 B.n445 10.6151
R1193 B.n447 B.n446 10.6151
R1194 B.n447 B.n401 10.6151
R1195 B.n453 B.n401 10.6151
R1196 B.n454 B.n453 10.6151
R1197 B.n455 B.n454 10.6151
R1198 B.n455 B.n399 10.6151
R1199 B.n461 B.n399 10.6151
R1200 B.n462 B.n461 10.6151
R1201 B.n463 B.n462 10.6151
R1202 B.n463 B.n397 10.6151
R1203 B.n469 B.n397 10.6151
R1204 B.n470 B.n469 10.6151
R1205 B.n471 B.n470 10.6151
R1206 B.n471 B.n395 10.6151
R1207 B.n477 B.n395 10.6151
R1208 B.n478 B.n477 10.6151
R1209 B.n479 B.n478 10.6151
R1210 B.n479 B.n393 10.6151
R1211 B.n485 B.n393 10.6151
R1212 B.n486 B.n485 10.6151
R1213 B.n487 B.n486 10.6151
R1214 B.n487 B.n391 10.6151
R1215 B.n493 B.n391 10.6151
R1216 B.n494 B.n493 10.6151
R1217 B.n495 B.n494 10.6151
R1218 B.n495 B.n389 10.6151
R1219 B.n502 B.n501 10.6151
R1220 B.n503 B.n502 10.6151
R1221 B.n503 B.n384 10.6151
R1222 B.n509 B.n384 10.6151
R1223 B.n510 B.n509 10.6151
R1224 B.n511 B.n510 10.6151
R1225 B.n511 B.n382 10.6151
R1226 B.n517 B.n382 10.6151
R1227 B.n520 B.n519 10.6151
R1228 B.n520 B.n378 10.6151
R1229 B.n526 B.n378 10.6151
R1230 B.n527 B.n526 10.6151
R1231 B.n528 B.n527 10.6151
R1232 B.n528 B.n376 10.6151
R1233 B.n534 B.n376 10.6151
R1234 B.n535 B.n534 10.6151
R1235 B.n536 B.n535 10.6151
R1236 B.n536 B.n374 10.6151
R1237 B.n542 B.n374 10.6151
R1238 B.n543 B.n542 10.6151
R1239 B.n544 B.n543 10.6151
R1240 B.n544 B.n372 10.6151
R1241 B.n550 B.n372 10.6151
R1242 B.n551 B.n550 10.6151
R1243 B.n552 B.n551 10.6151
R1244 B.n552 B.n370 10.6151
R1245 B.n558 B.n370 10.6151
R1246 B.n559 B.n558 10.6151
R1247 B.n560 B.n559 10.6151
R1248 B.n560 B.n368 10.6151
R1249 B.n566 B.n368 10.6151
R1250 B.n567 B.n566 10.6151
R1251 B.n568 B.n567 10.6151
R1252 B.n568 B.n366 10.6151
R1253 B.n574 B.n366 10.6151
R1254 B.n575 B.n574 10.6151
R1255 B.n576 B.n575 10.6151
R1256 B.n576 B.n364 10.6151
R1257 B.n582 B.n364 10.6151
R1258 B.n583 B.n582 10.6151
R1259 B.n584 B.n583 10.6151
R1260 B.n584 B.n362 10.6151
R1261 B.n590 B.n362 10.6151
R1262 B.n591 B.n590 10.6151
R1263 B.n592 B.n591 10.6151
R1264 B.n592 B.n360 10.6151
R1265 B.n598 B.n360 10.6151
R1266 B.n599 B.n598 10.6151
R1267 B.n600 B.n599 10.6151
R1268 B.n600 B.n358 10.6151
R1269 B.n606 B.n358 10.6151
R1270 B.n607 B.n606 10.6151
R1271 B.n613 B.n612 10.6151
R1272 B.n614 B.n613 10.6151
R1273 B.n614 B.n346 10.6151
R1274 B.n625 B.n346 10.6151
R1275 B.n626 B.n625 10.6151
R1276 B.n627 B.n626 10.6151
R1277 B.n627 B.n339 10.6151
R1278 B.n637 B.n339 10.6151
R1279 B.n638 B.n637 10.6151
R1280 B.n639 B.n638 10.6151
R1281 B.n639 B.n331 10.6151
R1282 B.n649 B.n331 10.6151
R1283 B.n650 B.n649 10.6151
R1284 B.n651 B.n650 10.6151
R1285 B.n651 B.n323 10.6151
R1286 B.n661 B.n323 10.6151
R1287 B.n662 B.n661 10.6151
R1288 B.n663 B.n662 10.6151
R1289 B.n663 B.n315 10.6151
R1290 B.n674 B.n315 10.6151
R1291 B.n675 B.n674 10.6151
R1292 B.n676 B.n675 10.6151
R1293 B.n676 B.n308 10.6151
R1294 B.n687 B.n308 10.6151
R1295 B.n688 B.n687 10.6151
R1296 B.n689 B.n688 10.6151
R1297 B.n689 B.n0 10.6151
R1298 B.n786 B.n1 10.6151
R1299 B.n786 B.n785 10.6151
R1300 B.n785 B.n784 10.6151
R1301 B.n784 B.n10 10.6151
R1302 B.n778 B.n10 10.6151
R1303 B.n778 B.n777 10.6151
R1304 B.n777 B.n776 10.6151
R1305 B.n776 B.n16 10.6151
R1306 B.n770 B.n16 10.6151
R1307 B.n770 B.n769 10.6151
R1308 B.n769 B.n768 10.6151
R1309 B.n768 B.n24 10.6151
R1310 B.n762 B.n24 10.6151
R1311 B.n762 B.n761 10.6151
R1312 B.n761 B.n760 10.6151
R1313 B.n760 B.n31 10.6151
R1314 B.n754 B.n31 10.6151
R1315 B.n754 B.n753 10.6151
R1316 B.n753 B.n752 10.6151
R1317 B.n752 B.n38 10.6151
R1318 B.n746 B.n38 10.6151
R1319 B.n746 B.n745 10.6151
R1320 B.n745 B.n744 10.6151
R1321 B.n744 B.n44 10.6151
R1322 B.n738 B.n44 10.6151
R1323 B.n738 B.n737 10.6151
R1324 B.n737 B.n736 10.6151
R1325 B.t3 B.n306 10.1608
R1326 B.t8 B.n8 10.1608
R1327 B.n665 B.t0 6.5748
R1328 B.t2 B.n772 6.5748
R1329 B.n199 B.n198 6.5566
R1330 B.n215 B.n107 6.5566
R1331 B.n501 B.n388 6.5566
R1332 B.n518 B.n517 6.5566
R1333 B.t4 B.n325 5.37947
R1334 B.n765 B.t7 5.37947
R1335 B.n198 B.n197 4.05904
R1336 B.n218 B.n107 4.05904
R1337 B.n389 B.n388 4.05904
R1338 B.n519 B.n518 4.05904
R1339 B.n622 B.t11 2.98882
R1340 B.n46 B.t15 2.98882
R1341 B.n792 B.n0 2.81026
R1342 B.n792 B.n1 2.81026
R1343 VP.n6 VP.t4 473.207
R1344 VP.n14 VP.t1 450.579
R1345 VP.n16 VP.t2 450.579
R1346 VP.n1 VP.t7 450.579
R1347 VP.n20 VP.t9 450.579
R1348 VP.n22 VP.t5 450.579
R1349 VP.n11 VP.t8 450.579
R1350 VP.n9 VP.t3 450.579
R1351 VP.n8 VP.t6 450.579
R1352 VP.n7 VP.t0 450.579
R1353 VP.n23 VP.n22 161.3
R1354 VP.n10 VP.n3 161.3
R1355 VP.n12 VP.n11 161.3
R1356 VP.n21 VP.n0 161.3
R1357 VP.n15 VP.n2 161.3
R1358 VP.n14 VP.n13 161.3
R1359 VP.n8 VP.n5 80.6037
R1360 VP.n9 VP.n4 80.6037
R1361 VP.n20 VP.n19 80.6037
R1362 VP.n18 VP.n1 80.6037
R1363 VP.n17 VP.n16 80.6037
R1364 VP.n16 VP.n1 48.2005
R1365 VP.n20 VP.n1 48.2005
R1366 VP.n9 VP.n8 48.2005
R1367 VP.n8 VP.n7 48.2005
R1368 VP.n13 VP.n12 44.099
R1369 VP.n16 VP.n15 34.3247
R1370 VP.n21 VP.n20 34.3247
R1371 VP.n10 VP.n9 34.3247
R1372 VP.n6 VP.n5 31.798
R1373 VP.n7 VP.n6 16.5773
R1374 VP.n15 VP.n14 13.8763
R1375 VP.n22 VP.n21 13.8763
R1376 VP.n11 VP.n10 13.8763
R1377 VP.n5 VP.n4 0.380177
R1378 VP.n18 VP.n17 0.380177
R1379 VP.n19 VP.n18 0.380177
R1380 VP.n4 VP.n3 0.285035
R1381 VP.n17 VP.n2 0.285035
R1382 VP.n19 VP.n0 0.285035
R1383 VP.n12 VP.n3 0.189894
R1384 VP.n13 VP.n2 0.189894
R1385 VP.n23 VP.n0 0.189894
R1386 VP VP.n23 0.0516364
R1387 VDD1.n1 VDD1.t5 62.7412
R1388 VDD1.n3 VDD1.t2 62.741
R1389 VDD1.n5 VDD1.n4 60.9365
R1390 VDD1.n1 VDD1.n0 60.2677
R1391 VDD1.n3 VDD1.n2 60.2677
R1392 VDD1.n7 VDD1.n6 60.2676
R1393 VDD1.n7 VDD1.n5 40.6862
R1394 VDD1.n6 VDD1.t1 1.5085
R1395 VDD1.n6 VDD1.t7 1.5085
R1396 VDD1.n0 VDD1.t6 1.5085
R1397 VDD1.n0 VDD1.t3 1.5085
R1398 VDD1.n4 VDD1.t9 1.5085
R1399 VDD1.n4 VDD1.t0 1.5085
R1400 VDD1.n2 VDD1.t4 1.5085
R1401 VDD1.n2 VDD1.t8 1.5085
R1402 VDD1 VDD1.n7 0.666448
R1403 VDD1 VDD1.n1 0.300069
R1404 VDD1.n5 VDD1.n3 0.186533
R1405 VTAIL.n11 VTAIL.t2 45.0969
R1406 VTAIL.n17 VTAIL.t4 45.0967
R1407 VTAIL.n2 VTAIL.t13 45.0967
R1408 VTAIL.n16 VTAIL.t10 45.0967
R1409 VTAIL.n15 VTAIL.n14 43.5889
R1410 VTAIL.n13 VTAIL.n12 43.5889
R1411 VTAIL.n10 VTAIL.n9 43.5889
R1412 VTAIL.n8 VTAIL.n7 43.5889
R1413 VTAIL.n19 VTAIL.n18 43.5889
R1414 VTAIL.n1 VTAIL.n0 43.5889
R1415 VTAIL.n4 VTAIL.n3 43.5889
R1416 VTAIL.n6 VTAIL.n5 43.5889
R1417 VTAIL.n8 VTAIL.n6 25.6169
R1418 VTAIL.n17 VTAIL.n16 24.6514
R1419 VTAIL.n18 VTAIL.t1 1.5085
R1420 VTAIL.n18 VTAIL.t8 1.5085
R1421 VTAIL.n0 VTAIL.t5 1.5085
R1422 VTAIL.n0 VTAIL.t7 1.5085
R1423 VTAIL.n3 VTAIL.t11 1.5085
R1424 VTAIL.n3 VTAIL.t9 1.5085
R1425 VTAIL.n5 VTAIL.t17 1.5085
R1426 VTAIL.n5 VTAIL.t16 1.5085
R1427 VTAIL.n14 VTAIL.t12 1.5085
R1428 VTAIL.n14 VTAIL.t15 1.5085
R1429 VTAIL.n12 VTAIL.t14 1.5085
R1430 VTAIL.n12 VTAIL.t18 1.5085
R1431 VTAIL.n9 VTAIL.t0 1.5085
R1432 VTAIL.n9 VTAIL.t19 1.5085
R1433 VTAIL.n7 VTAIL.t6 1.5085
R1434 VTAIL.n7 VTAIL.t3 1.5085
R1435 VTAIL.n10 VTAIL.n8 0.966017
R1436 VTAIL.n11 VTAIL.n10 0.966017
R1437 VTAIL.n15 VTAIL.n13 0.966017
R1438 VTAIL.n16 VTAIL.n15 0.966017
R1439 VTAIL.n6 VTAIL.n4 0.966017
R1440 VTAIL.n4 VTAIL.n2 0.966017
R1441 VTAIL.n19 VTAIL.n17 0.966017
R1442 VTAIL.n13 VTAIL.n11 0.953086
R1443 VTAIL.n2 VTAIL.n1 0.953086
R1444 VTAIL VTAIL.n1 0.782828
R1445 VTAIL VTAIL.n19 0.18369
R1446 VN.n3 VN.t2 473.207
R1447 VN.n13 VN.t5 473.207
R1448 VN.n2 VN.t4 450.579
R1449 VN.n1 VN.t8 450.579
R1450 VN.n6 VN.t3 450.579
R1451 VN.n8 VN.t7 450.579
R1452 VN.n12 VN.t0 450.579
R1453 VN.n11 VN.t9 450.579
R1454 VN.n16 VN.t6 450.579
R1455 VN.n18 VN.t1 450.579
R1456 VN.n9 VN.n8 161.3
R1457 VN.n19 VN.n18 161.3
R1458 VN.n17 VN.n10 161.3
R1459 VN.n7 VN.n0 161.3
R1460 VN.n16 VN.n15 80.6037
R1461 VN.n14 VN.n11 80.6037
R1462 VN.n6 VN.n5 80.6037
R1463 VN.n4 VN.n1 80.6037
R1464 VN.n2 VN.n1 48.2005
R1465 VN.n6 VN.n1 48.2005
R1466 VN.n12 VN.n11 48.2005
R1467 VN.n16 VN.n11 48.2005
R1468 VN VN.n19 44.4797
R1469 VN.n7 VN.n6 34.3247
R1470 VN.n17 VN.n16 34.3247
R1471 VN.n14 VN.n13 31.798
R1472 VN.n4 VN.n3 31.798
R1473 VN.n3 VN.n2 16.5773
R1474 VN.n13 VN.n12 16.5773
R1475 VN.n8 VN.n7 13.8763
R1476 VN.n18 VN.n17 13.8763
R1477 VN.n15 VN.n14 0.380177
R1478 VN.n5 VN.n4 0.380177
R1479 VN.n15 VN.n10 0.285035
R1480 VN.n5 VN.n0 0.285035
R1481 VN.n19 VN.n10 0.189894
R1482 VN.n9 VN.n0 0.189894
R1483 VN VN.n9 0.0516364
R1484 VDD2.n1 VDD2.t7 62.741
R1485 VDD2.n4 VDD2.t8 61.7757
R1486 VDD2.n3 VDD2.n2 60.9365
R1487 VDD2 VDD2.n7 60.9335
R1488 VDD2.n6 VDD2.n5 60.2677
R1489 VDD2.n1 VDD2.n0 60.2677
R1490 VDD2.n4 VDD2.n3 39.6205
R1491 VDD2.n7 VDD2.t9 1.5085
R1492 VDD2.n7 VDD2.t4 1.5085
R1493 VDD2.n5 VDD2.t3 1.5085
R1494 VDD2.n5 VDD2.t0 1.5085
R1495 VDD2.n2 VDD2.t6 1.5085
R1496 VDD2.n2 VDD2.t2 1.5085
R1497 VDD2.n0 VDD2.t5 1.5085
R1498 VDD2.n0 VDD2.t1 1.5085
R1499 VDD2.n6 VDD2.n4 0.966017
R1500 VDD2 VDD2.n6 0.300069
R1501 VDD2.n3 VDD2.n1 0.186533
C0 VDD2 VP 0.353136f
C1 VP VN 5.94089f
C2 VP VDD1 7.94522f
C3 VP VTAIL 7.59949f
C4 VDD2 VN 7.74624f
C5 VDD2 VDD1 1.02884f
C6 VDD2 VTAIL 14.5585f
C7 VDD1 VN 0.149175f
C8 VN VTAIL 7.58486f
C9 VDD1 VTAIL 14.523999f
C10 VDD2 B 5.283757f
C11 VDD1 B 5.21204f
C12 VTAIL B 7.018719f
C13 VN B 9.966479f
C14 VP B 8.011223f
C15 VDD2.t7 B 2.84663f
C16 VDD2.t5 B 0.24887f
C17 VDD2.t1 B 0.24887f
C18 VDD2.n0 B 2.22737f
C19 VDD2.n1 B 0.639146f
C20 VDD2.t6 B 0.24887f
C21 VDD2.t2 B 0.24887f
C22 VDD2.n2 B 2.23108f
C23 VDD2.n3 B 1.94251f
C24 VDD2.t8 B 2.84123f
C25 VDD2.n4 B 2.41479f
C26 VDD2.t3 B 0.24887f
C27 VDD2.t0 B 0.24887f
C28 VDD2.n5 B 2.22736f
C29 VDD2.n6 B 0.299477f
C30 VDD2.t9 B 0.24887f
C31 VDD2.t4 B 0.24887f
C32 VDD2.n7 B 2.23104f
C33 VN.n0 B 0.05409f
C34 VN.t8 B 1.19749f
C35 VN.n1 B 0.479984f
C36 VN.t2 B 1.22f
C37 VN.t4 B 1.19749f
C38 VN.n2 B 0.479102f
C39 VN.n3 B 0.452551f
C40 VN.n4 B 0.247526f
C41 VN.n5 B 0.067518f
C42 VN.t3 B 1.19749f
C43 VN.n6 B 0.47761f
C44 VN.n7 B 0.009198f
C45 VN.t7 B 1.19749f
C46 VN.n8 B 0.464912f
C47 VN.n9 B 0.031414f
C48 VN.n10 B 0.05409f
C49 VN.t9 B 1.19749f
C50 VN.n11 B 0.479984f
C51 VN.t6 B 1.19749f
C52 VN.t5 B 1.22f
C53 VN.t0 B 1.19749f
C54 VN.n12 B 0.479102f
C55 VN.n13 B 0.452551f
C56 VN.n14 B 0.247526f
C57 VN.n15 B 0.067518f
C58 VN.n16 B 0.47761f
C59 VN.n17 B 0.009198f
C60 VN.t1 B 1.19749f
C61 VN.n18 B 0.464912f
C62 VN.n19 B 1.83905f
C63 VTAIL.t5 B 0.261297f
C64 VTAIL.t7 B 0.261297f
C65 VTAIL.n0 B 2.25939f
C66 VTAIL.n1 B 0.397523f
C67 VTAIL.t13 B 2.88136f
C68 VTAIL.n2 B 0.503043f
C69 VTAIL.t11 B 0.261297f
C70 VTAIL.t9 B 0.261297f
C71 VTAIL.n3 B 2.25939f
C72 VTAIL.n4 B 0.413438f
C73 VTAIL.t17 B 0.261297f
C74 VTAIL.t16 B 0.261297f
C75 VTAIL.n5 B 2.25939f
C76 VTAIL.n6 B 1.75237f
C77 VTAIL.t6 B 0.261297f
C78 VTAIL.t3 B 0.261297f
C79 VTAIL.n7 B 2.25939f
C80 VTAIL.n8 B 1.75237f
C81 VTAIL.t0 B 0.261297f
C82 VTAIL.t19 B 0.261297f
C83 VTAIL.n9 B 2.25939f
C84 VTAIL.n10 B 0.41344f
C85 VTAIL.t2 B 2.88137f
C86 VTAIL.n11 B 0.503035f
C87 VTAIL.t14 B 0.261297f
C88 VTAIL.t18 B 0.261297f
C89 VTAIL.n12 B 2.25939f
C90 VTAIL.n13 B 0.412391f
C91 VTAIL.t12 B 0.261297f
C92 VTAIL.t15 B 0.261297f
C93 VTAIL.n14 B 2.25939f
C94 VTAIL.n15 B 0.41344f
C95 VTAIL.t10 B 2.88136f
C96 VTAIL.n16 B 1.76468f
C97 VTAIL.t4 B 2.88136f
C98 VTAIL.n17 B 1.76468f
C99 VTAIL.t1 B 0.261297f
C100 VTAIL.t8 B 0.261297f
C101 VTAIL.n18 B 2.25939f
C102 VTAIL.n19 B 0.349954f
C103 VDD1.t5 B 2.84808f
C104 VDD1.t6 B 0.248997f
C105 VDD1.t3 B 0.248997f
C106 VDD1.n0 B 2.2285f
C107 VDD1.n1 B 0.645257f
C108 VDD1.t2 B 2.84808f
C109 VDD1.t4 B 0.248997f
C110 VDD1.t8 B 0.248997f
C111 VDD1.n2 B 2.2285f
C112 VDD1.n3 B 0.639471f
C113 VDD1.t9 B 0.248997f
C114 VDD1.t0 B 0.248997f
C115 VDD1.n4 B 2.23222f
C116 VDD1.n5 B 2.0198f
C117 VDD1.t1 B 0.248997f
C118 VDD1.t7 B 0.248997f
C119 VDD1.n6 B 2.22849f
C120 VDD1.n7 B 2.41497f
C121 VP.n0 B 0.054748f
C122 VP.t7 B 1.21205f
C123 VP.n1 B 0.485818f
C124 VP.n2 B 0.054748f
C125 VP.n3 B 0.054748f
C126 VP.t8 B 1.21205f
C127 VP.t3 B 1.21205f
C128 VP.n4 B 0.068338f
C129 VP.t6 B 1.21205f
C130 VP.n5 B 0.250534f
C131 VP.t0 B 1.21205f
C132 VP.t4 B 1.23483f
C133 VP.n6 B 0.458051f
C134 VP.n7 B 0.484926f
C135 VP.n8 B 0.485818f
C136 VP.n9 B 0.483415f
C137 VP.n10 B 0.00931f
C138 VP.n11 B 0.470563f
C139 VP.n12 B 1.83455f
C140 VP.n13 B 1.86799f
C141 VP.t1 B 1.21205f
C142 VP.n14 B 0.470563f
C143 VP.n15 B 0.00931f
C144 VP.t2 B 1.21205f
C145 VP.n16 B 0.483415f
C146 VP.n17 B 0.068338f
C147 VP.n18 B 0.082057f
C148 VP.n19 B 0.068338f
C149 VP.t9 B 1.21205f
C150 VP.n20 B 0.483415f
C151 VP.n21 B 0.00931f
C152 VP.t5 B 1.21205f
C153 VP.n22 B 0.470563f
C154 VP.n23 B 0.031796f
.ends

