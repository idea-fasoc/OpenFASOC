* NGSPICE file created from diff_pair_sample_0386.ext - technology: sky130A

.subckt diff_pair_sample_0386 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=0.5544 pd=3.69 as=0.5544 ps=3.69 w=3.36 l=2.98
X1 VDD2.t5 VN.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.3104 pd=7.5 as=0.5544 ps=3.69 w=3.36 l=2.98
X2 VDD1.t4 VP.t1 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=1.3104 pd=7.5 as=0.5544 ps=3.69 w=3.36 l=2.98
X3 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=1.3104 pd=7.5 as=0 ps=0 w=3.36 l=2.98
X4 VTAIL.t3 VN.t1 VDD2.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.5544 pd=3.69 as=0.5544 ps=3.69 w=3.36 l=2.98
X5 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=1.3104 pd=7.5 as=0 ps=0 w=3.36 l=2.98
X6 VTAIL.t9 VP.t2 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.5544 pd=3.69 as=0.5544 ps=3.69 w=3.36 l=2.98
X7 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.3104 pd=7.5 as=0 ps=0 w=3.36 l=2.98
X8 VDD2.t3 VN.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5544 pd=3.69 as=1.3104 ps=7.5 w=3.36 l=2.98
X9 VDD1.t1 VP.t3 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=1.3104 pd=7.5 as=0.5544 ps=3.69 w=3.36 l=2.98
X10 VDD2.t2 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5544 pd=3.69 as=1.3104 ps=7.5 w=3.36 l=2.98
X11 VDD1.t3 VP.t4 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5544 pd=3.69 as=1.3104 ps=7.5 w=3.36 l=2.98
X12 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.3104 pd=7.5 as=0 ps=0 w=3.36 l=2.98
X13 VDD2.t1 VN.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.3104 pd=7.5 as=0.5544 ps=3.69 w=3.36 l=2.98
X14 VTAIL.t0 VN.t5 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.5544 pd=3.69 as=0.5544 ps=3.69 w=3.36 l=2.98
X15 VDD1.t0 VP.t5 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5544 pd=3.69 as=1.3104 ps=7.5 w=3.36 l=2.98
R0 VP.n14 VP.n11 161.3
R1 VP.n16 VP.n15 161.3
R2 VP.n17 VP.n10 161.3
R3 VP.n19 VP.n18 161.3
R4 VP.n20 VP.n9 161.3
R5 VP.n22 VP.n21 161.3
R6 VP.n23 VP.n8 161.3
R7 VP.n48 VP.n0 161.3
R8 VP.n47 VP.n46 161.3
R9 VP.n45 VP.n1 161.3
R10 VP.n44 VP.n43 161.3
R11 VP.n42 VP.n2 161.3
R12 VP.n41 VP.n40 161.3
R13 VP.n39 VP.n3 161.3
R14 VP.n38 VP.n37 161.3
R15 VP.n35 VP.n4 161.3
R16 VP.n34 VP.n33 161.3
R17 VP.n32 VP.n5 161.3
R18 VP.n31 VP.n30 161.3
R19 VP.n29 VP.n6 161.3
R20 VP.n28 VP.n27 161.3
R21 VP.n26 VP.n7 107.957
R22 VP.n50 VP.n49 107.957
R23 VP.n25 VP.n24 107.957
R24 VP.n13 VP.n12 61.8105
R25 VP.n13 VP.t1 60.2918
R26 VP.n34 VP.n5 49.7803
R27 VP.n43 VP.n42 49.7803
R28 VP.n18 VP.n17 49.7803
R29 VP.n26 VP.n25 43.6247
R30 VP.n30 VP.n5 31.3737
R31 VP.n43 VP.n1 31.3737
R32 VP.n18 VP.n9 31.3737
R33 VP.n7 VP.t3 27.1737
R34 VP.n36 VP.t2 27.1737
R35 VP.n49 VP.t4 27.1737
R36 VP.n24 VP.t5 27.1737
R37 VP.n12 VP.t0 27.1737
R38 VP.n29 VP.n28 24.5923
R39 VP.n30 VP.n29 24.5923
R40 VP.n35 VP.n34 24.5923
R41 VP.n37 VP.n35 24.5923
R42 VP.n41 VP.n3 24.5923
R43 VP.n42 VP.n41 24.5923
R44 VP.n47 VP.n1 24.5923
R45 VP.n48 VP.n47 24.5923
R46 VP.n22 VP.n9 24.5923
R47 VP.n23 VP.n22 24.5923
R48 VP.n16 VP.n11 24.5923
R49 VP.n17 VP.n16 24.5923
R50 VP.n37 VP.n36 12.2964
R51 VP.n36 VP.n3 12.2964
R52 VP.n12 VP.n11 12.2964
R53 VP.n14 VP.n13 5.06578
R54 VP.n28 VP.n7 2.95152
R55 VP.n49 VP.n48 2.95152
R56 VP.n24 VP.n23 2.95152
R57 VP.n25 VP.n8 0.278335
R58 VP.n27 VP.n26 0.278335
R59 VP.n50 VP.n0 0.278335
R60 VP.n15 VP.n14 0.189894
R61 VP.n15 VP.n10 0.189894
R62 VP.n19 VP.n10 0.189894
R63 VP.n20 VP.n19 0.189894
R64 VP.n21 VP.n20 0.189894
R65 VP.n21 VP.n8 0.189894
R66 VP.n27 VP.n6 0.189894
R67 VP.n31 VP.n6 0.189894
R68 VP.n32 VP.n31 0.189894
R69 VP.n33 VP.n32 0.189894
R70 VP.n33 VP.n4 0.189894
R71 VP.n38 VP.n4 0.189894
R72 VP.n39 VP.n38 0.189894
R73 VP.n40 VP.n39 0.189894
R74 VP.n40 VP.n2 0.189894
R75 VP.n44 VP.n2 0.189894
R76 VP.n45 VP.n44 0.189894
R77 VP.n46 VP.n45 0.189894
R78 VP.n46 VP.n0 0.189894
R79 VP VP.n50 0.153485
R80 VDD1.n10 VDD1.n0 289.615
R81 VDD1.n25 VDD1.n15 289.615
R82 VDD1.n11 VDD1.n10 185
R83 VDD1.n9 VDD1.n8 185
R84 VDD1.n4 VDD1.n3 185
R85 VDD1.n19 VDD1.n18 185
R86 VDD1.n24 VDD1.n23 185
R87 VDD1.n26 VDD1.n25 185
R88 VDD1.n5 VDD1.t4 150.499
R89 VDD1.n20 VDD1.t1 150.499
R90 VDD1.n10 VDD1.n9 104.615
R91 VDD1.n9 VDD1.n3 104.615
R92 VDD1.n24 VDD1.n18 104.615
R93 VDD1.n25 VDD1.n24 104.615
R94 VDD1.n31 VDD1.n30 77.2016
R95 VDD1.n33 VDD1.n32 76.5436
R96 VDD1.t4 VDD1.n3 52.3082
R97 VDD1.t1 VDD1.n18 52.3082
R98 VDD1 VDD1.n14 48.7351
R99 VDD1.n31 VDD1.n29 48.6216
R100 VDD1.n33 VDD1.n31 37.8953
R101 VDD1.n5 VDD1.n4 10.2326
R102 VDD1.n20 VDD1.n19 10.2326
R103 VDD1.n14 VDD1.n0 9.69747
R104 VDD1.n29 VDD1.n15 9.69747
R105 VDD1.n14 VDD1.n13 9.45567
R106 VDD1.n29 VDD1.n28 9.45567
R107 VDD1.n2 VDD1.n1 9.3005
R108 VDD1.n13 VDD1.n12 9.3005
R109 VDD1.n7 VDD1.n6 9.3005
R110 VDD1.n22 VDD1.n21 9.3005
R111 VDD1.n17 VDD1.n16 9.3005
R112 VDD1.n28 VDD1.n27 9.3005
R113 VDD1.n12 VDD1.n11 8.92171
R114 VDD1.n27 VDD1.n26 8.92171
R115 VDD1.n8 VDD1.n2 8.14595
R116 VDD1.n23 VDD1.n17 8.14595
R117 VDD1.n7 VDD1.n4 7.3702
R118 VDD1.n22 VDD1.n19 7.3702
R119 VDD1.n32 VDD1.t5 5.89336
R120 VDD1.n32 VDD1.t0 5.89336
R121 VDD1.n30 VDD1.t2 5.89336
R122 VDD1.n30 VDD1.t3 5.89336
R123 VDD1.n8 VDD1.n7 5.81868
R124 VDD1.n23 VDD1.n22 5.81868
R125 VDD1.n11 VDD1.n2 5.04292
R126 VDD1.n26 VDD1.n17 5.04292
R127 VDD1.n12 VDD1.n0 4.26717
R128 VDD1.n27 VDD1.n15 4.26717
R129 VDD1.n6 VDD1.n5 2.88718
R130 VDD1.n21 VDD1.n20 2.88718
R131 VDD1 VDD1.n33 0.655672
R132 VDD1.n13 VDD1.n1 0.155672
R133 VDD1.n6 VDD1.n1 0.155672
R134 VDD1.n21 VDD1.n16 0.155672
R135 VDD1.n28 VDD1.n16 0.155672
R136 VTAIL.n66 VTAIL.n56 289.615
R137 VTAIL.n12 VTAIL.n2 289.615
R138 VTAIL.n50 VTAIL.n40 289.615
R139 VTAIL.n32 VTAIL.n22 289.615
R140 VTAIL.n60 VTAIL.n59 185
R141 VTAIL.n65 VTAIL.n64 185
R142 VTAIL.n67 VTAIL.n66 185
R143 VTAIL.n6 VTAIL.n5 185
R144 VTAIL.n11 VTAIL.n10 185
R145 VTAIL.n13 VTAIL.n12 185
R146 VTAIL.n51 VTAIL.n50 185
R147 VTAIL.n49 VTAIL.n48 185
R148 VTAIL.n44 VTAIL.n43 185
R149 VTAIL.n33 VTAIL.n32 185
R150 VTAIL.n31 VTAIL.n30 185
R151 VTAIL.n26 VTAIL.n25 185
R152 VTAIL.n61 VTAIL.t5 150.499
R153 VTAIL.n7 VTAIL.t7 150.499
R154 VTAIL.n27 VTAIL.t2 150.499
R155 VTAIL.n45 VTAIL.t6 150.499
R156 VTAIL.n65 VTAIL.n59 104.615
R157 VTAIL.n66 VTAIL.n65 104.615
R158 VTAIL.n11 VTAIL.n5 104.615
R159 VTAIL.n12 VTAIL.n11 104.615
R160 VTAIL.n50 VTAIL.n49 104.615
R161 VTAIL.n49 VTAIL.n43 104.615
R162 VTAIL.n32 VTAIL.n31 104.615
R163 VTAIL.n31 VTAIL.n25 104.615
R164 VTAIL.n39 VTAIL.n38 59.8648
R165 VTAIL.n21 VTAIL.n20 59.8648
R166 VTAIL.n1 VTAIL.n0 59.8648
R167 VTAIL.n19 VTAIL.n18 59.8648
R168 VTAIL.t5 VTAIL.n59 52.3082
R169 VTAIL.t7 VTAIL.n5 52.3082
R170 VTAIL.t6 VTAIL.n43 52.3082
R171 VTAIL.t2 VTAIL.n25 52.3082
R172 VTAIL.n71 VTAIL.n70 29.8581
R173 VTAIL.n17 VTAIL.n16 29.8581
R174 VTAIL.n55 VTAIL.n54 29.8581
R175 VTAIL.n37 VTAIL.n36 29.8581
R176 VTAIL.n21 VTAIL.n19 20.9703
R177 VTAIL.n71 VTAIL.n55 18.1169
R178 VTAIL.n61 VTAIL.n60 10.2326
R179 VTAIL.n7 VTAIL.n6 10.2326
R180 VTAIL.n45 VTAIL.n44 10.2326
R181 VTAIL.n27 VTAIL.n26 10.2326
R182 VTAIL.n70 VTAIL.n56 9.69747
R183 VTAIL.n16 VTAIL.n2 9.69747
R184 VTAIL.n54 VTAIL.n40 9.69747
R185 VTAIL.n36 VTAIL.n22 9.69747
R186 VTAIL.n70 VTAIL.n69 9.45567
R187 VTAIL.n16 VTAIL.n15 9.45567
R188 VTAIL.n54 VTAIL.n53 9.45567
R189 VTAIL.n36 VTAIL.n35 9.45567
R190 VTAIL.n63 VTAIL.n62 9.3005
R191 VTAIL.n58 VTAIL.n57 9.3005
R192 VTAIL.n69 VTAIL.n68 9.3005
R193 VTAIL.n9 VTAIL.n8 9.3005
R194 VTAIL.n4 VTAIL.n3 9.3005
R195 VTAIL.n15 VTAIL.n14 9.3005
R196 VTAIL.n42 VTAIL.n41 9.3005
R197 VTAIL.n47 VTAIL.n46 9.3005
R198 VTAIL.n53 VTAIL.n52 9.3005
R199 VTAIL.n24 VTAIL.n23 9.3005
R200 VTAIL.n35 VTAIL.n34 9.3005
R201 VTAIL.n29 VTAIL.n28 9.3005
R202 VTAIL.n68 VTAIL.n67 8.92171
R203 VTAIL.n14 VTAIL.n13 8.92171
R204 VTAIL.n52 VTAIL.n51 8.92171
R205 VTAIL.n34 VTAIL.n33 8.92171
R206 VTAIL.n64 VTAIL.n58 8.14595
R207 VTAIL.n10 VTAIL.n4 8.14595
R208 VTAIL.n48 VTAIL.n42 8.14595
R209 VTAIL.n30 VTAIL.n24 8.14595
R210 VTAIL.n63 VTAIL.n60 7.3702
R211 VTAIL.n9 VTAIL.n6 7.3702
R212 VTAIL.n47 VTAIL.n44 7.3702
R213 VTAIL.n29 VTAIL.n26 7.3702
R214 VTAIL.n0 VTAIL.t1 5.89336
R215 VTAIL.n0 VTAIL.t3 5.89336
R216 VTAIL.n18 VTAIL.t8 5.89336
R217 VTAIL.n18 VTAIL.t9 5.89336
R218 VTAIL.n38 VTAIL.t10 5.89336
R219 VTAIL.n38 VTAIL.t11 5.89336
R220 VTAIL.n20 VTAIL.t4 5.89336
R221 VTAIL.n20 VTAIL.t0 5.89336
R222 VTAIL.n64 VTAIL.n63 5.81868
R223 VTAIL.n10 VTAIL.n9 5.81868
R224 VTAIL.n48 VTAIL.n47 5.81868
R225 VTAIL.n30 VTAIL.n29 5.81868
R226 VTAIL.n67 VTAIL.n58 5.04292
R227 VTAIL.n13 VTAIL.n4 5.04292
R228 VTAIL.n51 VTAIL.n42 5.04292
R229 VTAIL.n33 VTAIL.n24 5.04292
R230 VTAIL.n68 VTAIL.n56 4.26717
R231 VTAIL.n14 VTAIL.n2 4.26717
R232 VTAIL.n52 VTAIL.n40 4.26717
R233 VTAIL.n34 VTAIL.n22 4.26717
R234 VTAIL.n62 VTAIL.n61 2.88718
R235 VTAIL.n8 VTAIL.n7 2.88718
R236 VTAIL.n46 VTAIL.n45 2.88718
R237 VTAIL.n28 VTAIL.n27 2.88718
R238 VTAIL.n37 VTAIL.n21 2.85395
R239 VTAIL.n55 VTAIL.n39 2.85395
R240 VTAIL.n19 VTAIL.n17 2.85395
R241 VTAIL VTAIL.n71 2.0824
R242 VTAIL.n39 VTAIL.n37 1.89705
R243 VTAIL.n17 VTAIL.n1 1.89705
R244 VTAIL VTAIL.n1 0.772052
R245 VTAIL.n62 VTAIL.n57 0.155672
R246 VTAIL.n69 VTAIL.n57 0.155672
R247 VTAIL.n8 VTAIL.n3 0.155672
R248 VTAIL.n15 VTAIL.n3 0.155672
R249 VTAIL.n53 VTAIL.n41 0.155672
R250 VTAIL.n46 VTAIL.n41 0.155672
R251 VTAIL.n35 VTAIL.n23 0.155672
R252 VTAIL.n28 VTAIL.n23 0.155672
R253 B.n596 B.n595 585
R254 B.n192 B.n108 585
R255 B.n191 B.n190 585
R256 B.n189 B.n188 585
R257 B.n187 B.n186 585
R258 B.n185 B.n184 585
R259 B.n183 B.n182 585
R260 B.n181 B.n180 585
R261 B.n179 B.n178 585
R262 B.n177 B.n176 585
R263 B.n175 B.n174 585
R264 B.n173 B.n172 585
R265 B.n171 B.n170 585
R266 B.n169 B.n168 585
R267 B.n167 B.n166 585
R268 B.n165 B.n164 585
R269 B.n163 B.n162 585
R270 B.n161 B.n160 585
R271 B.n159 B.n158 585
R272 B.n157 B.n156 585
R273 B.n155 B.n154 585
R274 B.n153 B.n152 585
R275 B.n151 B.n150 585
R276 B.n149 B.n148 585
R277 B.n147 B.n146 585
R278 B.n145 B.n144 585
R279 B.n143 B.n142 585
R280 B.n141 B.n140 585
R281 B.n139 B.n138 585
R282 B.n137 B.n136 585
R283 B.n135 B.n134 585
R284 B.n133 B.n132 585
R285 B.n131 B.n130 585
R286 B.n129 B.n128 585
R287 B.n127 B.n126 585
R288 B.n125 B.n124 585
R289 B.n123 B.n122 585
R290 B.n121 B.n120 585
R291 B.n119 B.n118 585
R292 B.n117 B.n116 585
R293 B.n88 B.n87 585
R294 B.n601 B.n600 585
R295 B.n594 B.n109 585
R296 B.n109 B.n85 585
R297 B.n593 B.n84 585
R298 B.n605 B.n84 585
R299 B.n592 B.n83 585
R300 B.n606 B.n83 585
R301 B.n591 B.n82 585
R302 B.n607 B.n82 585
R303 B.n590 B.n589 585
R304 B.n589 B.n78 585
R305 B.n588 B.n77 585
R306 B.n613 B.n77 585
R307 B.n587 B.n76 585
R308 B.n614 B.n76 585
R309 B.n586 B.n75 585
R310 B.n615 B.n75 585
R311 B.n585 B.n584 585
R312 B.n584 B.n74 585
R313 B.n583 B.n70 585
R314 B.n621 B.n70 585
R315 B.n582 B.n69 585
R316 B.n622 B.n69 585
R317 B.n581 B.n68 585
R318 B.n623 B.n68 585
R319 B.n580 B.n579 585
R320 B.n579 B.n64 585
R321 B.n578 B.n63 585
R322 B.n629 B.n63 585
R323 B.n577 B.n62 585
R324 B.n630 B.n62 585
R325 B.n576 B.n61 585
R326 B.n631 B.n61 585
R327 B.n575 B.n574 585
R328 B.n574 B.n57 585
R329 B.n573 B.n56 585
R330 B.n637 B.n56 585
R331 B.n572 B.n55 585
R332 B.n638 B.n55 585
R333 B.n571 B.n54 585
R334 B.n639 B.n54 585
R335 B.n570 B.n569 585
R336 B.n569 B.n50 585
R337 B.n568 B.n49 585
R338 B.n645 B.n49 585
R339 B.n567 B.n48 585
R340 B.n646 B.n48 585
R341 B.n566 B.n47 585
R342 B.n647 B.n47 585
R343 B.n565 B.n564 585
R344 B.n564 B.n43 585
R345 B.n563 B.n42 585
R346 B.n653 B.n42 585
R347 B.n562 B.n41 585
R348 B.n654 B.n41 585
R349 B.n561 B.n40 585
R350 B.n655 B.n40 585
R351 B.n560 B.n559 585
R352 B.n559 B.n36 585
R353 B.n558 B.n35 585
R354 B.n661 B.n35 585
R355 B.n557 B.n34 585
R356 B.n662 B.n34 585
R357 B.n556 B.n33 585
R358 B.n663 B.n33 585
R359 B.n555 B.n554 585
R360 B.n554 B.n29 585
R361 B.n553 B.n28 585
R362 B.n669 B.n28 585
R363 B.n552 B.n27 585
R364 B.n670 B.n27 585
R365 B.n551 B.n26 585
R366 B.n671 B.n26 585
R367 B.n550 B.n549 585
R368 B.n549 B.n22 585
R369 B.n548 B.n21 585
R370 B.n677 B.n21 585
R371 B.n547 B.n20 585
R372 B.n678 B.n20 585
R373 B.n546 B.n19 585
R374 B.n679 B.n19 585
R375 B.n545 B.n544 585
R376 B.n544 B.n18 585
R377 B.n543 B.n14 585
R378 B.n685 B.n14 585
R379 B.n542 B.n13 585
R380 B.n686 B.n13 585
R381 B.n541 B.n12 585
R382 B.n687 B.n12 585
R383 B.n540 B.n539 585
R384 B.n539 B.n8 585
R385 B.n538 B.n7 585
R386 B.n693 B.n7 585
R387 B.n537 B.n6 585
R388 B.n694 B.n6 585
R389 B.n536 B.n5 585
R390 B.n695 B.n5 585
R391 B.n535 B.n534 585
R392 B.n534 B.n4 585
R393 B.n533 B.n193 585
R394 B.n533 B.n532 585
R395 B.n523 B.n194 585
R396 B.n195 B.n194 585
R397 B.n525 B.n524 585
R398 B.n526 B.n525 585
R399 B.n522 B.n200 585
R400 B.n200 B.n199 585
R401 B.n521 B.n520 585
R402 B.n520 B.n519 585
R403 B.n202 B.n201 585
R404 B.n512 B.n202 585
R405 B.n511 B.n510 585
R406 B.n513 B.n511 585
R407 B.n509 B.n207 585
R408 B.n207 B.n206 585
R409 B.n508 B.n507 585
R410 B.n507 B.n506 585
R411 B.n209 B.n208 585
R412 B.n210 B.n209 585
R413 B.n499 B.n498 585
R414 B.n500 B.n499 585
R415 B.n497 B.n215 585
R416 B.n215 B.n214 585
R417 B.n496 B.n495 585
R418 B.n495 B.n494 585
R419 B.n217 B.n216 585
R420 B.n218 B.n217 585
R421 B.n487 B.n486 585
R422 B.n488 B.n487 585
R423 B.n485 B.n222 585
R424 B.n226 B.n222 585
R425 B.n484 B.n483 585
R426 B.n483 B.n482 585
R427 B.n224 B.n223 585
R428 B.n225 B.n224 585
R429 B.n475 B.n474 585
R430 B.n476 B.n475 585
R431 B.n473 B.n231 585
R432 B.n231 B.n230 585
R433 B.n472 B.n471 585
R434 B.n471 B.n470 585
R435 B.n233 B.n232 585
R436 B.n234 B.n233 585
R437 B.n463 B.n462 585
R438 B.n464 B.n463 585
R439 B.n461 B.n239 585
R440 B.n239 B.n238 585
R441 B.n460 B.n459 585
R442 B.n459 B.n458 585
R443 B.n241 B.n240 585
R444 B.n242 B.n241 585
R445 B.n451 B.n450 585
R446 B.n452 B.n451 585
R447 B.n449 B.n247 585
R448 B.n247 B.n246 585
R449 B.n448 B.n447 585
R450 B.n447 B.n446 585
R451 B.n249 B.n248 585
R452 B.n250 B.n249 585
R453 B.n439 B.n438 585
R454 B.n440 B.n439 585
R455 B.n437 B.n255 585
R456 B.n255 B.n254 585
R457 B.n436 B.n435 585
R458 B.n435 B.n434 585
R459 B.n257 B.n256 585
R460 B.n258 B.n257 585
R461 B.n427 B.n426 585
R462 B.n428 B.n427 585
R463 B.n425 B.n263 585
R464 B.n263 B.n262 585
R465 B.n424 B.n423 585
R466 B.n423 B.n422 585
R467 B.n265 B.n264 585
R468 B.n415 B.n265 585
R469 B.n414 B.n413 585
R470 B.n416 B.n414 585
R471 B.n412 B.n270 585
R472 B.n270 B.n269 585
R473 B.n411 B.n410 585
R474 B.n410 B.n409 585
R475 B.n272 B.n271 585
R476 B.n273 B.n272 585
R477 B.n402 B.n401 585
R478 B.n403 B.n402 585
R479 B.n400 B.n278 585
R480 B.n278 B.n277 585
R481 B.n399 B.n398 585
R482 B.n398 B.n397 585
R483 B.n280 B.n279 585
R484 B.n281 B.n280 585
R485 B.n393 B.n392 585
R486 B.n284 B.n283 585
R487 B.n389 B.n388 585
R488 B.n390 B.n389 585
R489 B.n387 B.n305 585
R490 B.n386 B.n385 585
R491 B.n384 B.n383 585
R492 B.n382 B.n381 585
R493 B.n380 B.n379 585
R494 B.n378 B.n377 585
R495 B.n376 B.n375 585
R496 B.n374 B.n373 585
R497 B.n372 B.n371 585
R498 B.n370 B.n369 585
R499 B.n368 B.n367 585
R500 B.n366 B.n365 585
R501 B.n364 B.n363 585
R502 B.n361 B.n360 585
R503 B.n359 B.n358 585
R504 B.n357 B.n356 585
R505 B.n355 B.n354 585
R506 B.n353 B.n352 585
R507 B.n351 B.n350 585
R508 B.n349 B.n348 585
R509 B.n347 B.n346 585
R510 B.n345 B.n344 585
R511 B.n343 B.n342 585
R512 B.n340 B.n339 585
R513 B.n338 B.n337 585
R514 B.n336 B.n335 585
R515 B.n334 B.n333 585
R516 B.n332 B.n331 585
R517 B.n330 B.n329 585
R518 B.n328 B.n327 585
R519 B.n326 B.n325 585
R520 B.n324 B.n323 585
R521 B.n322 B.n321 585
R522 B.n320 B.n319 585
R523 B.n318 B.n317 585
R524 B.n316 B.n315 585
R525 B.n314 B.n313 585
R526 B.n312 B.n311 585
R527 B.n310 B.n304 585
R528 B.n390 B.n304 585
R529 B.n394 B.n282 585
R530 B.n282 B.n281 585
R531 B.n396 B.n395 585
R532 B.n397 B.n396 585
R533 B.n276 B.n275 585
R534 B.n277 B.n276 585
R535 B.n405 B.n404 585
R536 B.n404 B.n403 585
R537 B.n406 B.n274 585
R538 B.n274 B.n273 585
R539 B.n408 B.n407 585
R540 B.n409 B.n408 585
R541 B.n268 B.n267 585
R542 B.n269 B.n268 585
R543 B.n418 B.n417 585
R544 B.n417 B.n416 585
R545 B.n419 B.n266 585
R546 B.n415 B.n266 585
R547 B.n421 B.n420 585
R548 B.n422 B.n421 585
R549 B.n261 B.n260 585
R550 B.n262 B.n261 585
R551 B.n430 B.n429 585
R552 B.n429 B.n428 585
R553 B.n431 B.n259 585
R554 B.n259 B.n258 585
R555 B.n433 B.n432 585
R556 B.n434 B.n433 585
R557 B.n253 B.n252 585
R558 B.n254 B.n253 585
R559 B.n442 B.n441 585
R560 B.n441 B.n440 585
R561 B.n443 B.n251 585
R562 B.n251 B.n250 585
R563 B.n445 B.n444 585
R564 B.n446 B.n445 585
R565 B.n245 B.n244 585
R566 B.n246 B.n245 585
R567 B.n454 B.n453 585
R568 B.n453 B.n452 585
R569 B.n455 B.n243 585
R570 B.n243 B.n242 585
R571 B.n457 B.n456 585
R572 B.n458 B.n457 585
R573 B.n237 B.n236 585
R574 B.n238 B.n237 585
R575 B.n466 B.n465 585
R576 B.n465 B.n464 585
R577 B.n467 B.n235 585
R578 B.n235 B.n234 585
R579 B.n469 B.n468 585
R580 B.n470 B.n469 585
R581 B.n229 B.n228 585
R582 B.n230 B.n229 585
R583 B.n478 B.n477 585
R584 B.n477 B.n476 585
R585 B.n479 B.n227 585
R586 B.n227 B.n225 585
R587 B.n481 B.n480 585
R588 B.n482 B.n481 585
R589 B.n221 B.n220 585
R590 B.n226 B.n221 585
R591 B.n490 B.n489 585
R592 B.n489 B.n488 585
R593 B.n491 B.n219 585
R594 B.n219 B.n218 585
R595 B.n493 B.n492 585
R596 B.n494 B.n493 585
R597 B.n213 B.n212 585
R598 B.n214 B.n213 585
R599 B.n502 B.n501 585
R600 B.n501 B.n500 585
R601 B.n503 B.n211 585
R602 B.n211 B.n210 585
R603 B.n505 B.n504 585
R604 B.n506 B.n505 585
R605 B.n205 B.n204 585
R606 B.n206 B.n205 585
R607 B.n515 B.n514 585
R608 B.n514 B.n513 585
R609 B.n516 B.n203 585
R610 B.n512 B.n203 585
R611 B.n518 B.n517 585
R612 B.n519 B.n518 585
R613 B.n198 B.n197 585
R614 B.n199 B.n198 585
R615 B.n528 B.n527 585
R616 B.n527 B.n526 585
R617 B.n529 B.n196 585
R618 B.n196 B.n195 585
R619 B.n531 B.n530 585
R620 B.n532 B.n531 585
R621 B.n2 B.n0 585
R622 B.n4 B.n2 585
R623 B.n3 B.n1 585
R624 B.n694 B.n3 585
R625 B.n692 B.n691 585
R626 B.n693 B.n692 585
R627 B.n690 B.n9 585
R628 B.n9 B.n8 585
R629 B.n689 B.n688 585
R630 B.n688 B.n687 585
R631 B.n11 B.n10 585
R632 B.n686 B.n11 585
R633 B.n684 B.n683 585
R634 B.n685 B.n684 585
R635 B.n682 B.n15 585
R636 B.n18 B.n15 585
R637 B.n681 B.n680 585
R638 B.n680 B.n679 585
R639 B.n17 B.n16 585
R640 B.n678 B.n17 585
R641 B.n676 B.n675 585
R642 B.n677 B.n676 585
R643 B.n674 B.n23 585
R644 B.n23 B.n22 585
R645 B.n673 B.n672 585
R646 B.n672 B.n671 585
R647 B.n25 B.n24 585
R648 B.n670 B.n25 585
R649 B.n668 B.n667 585
R650 B.n669 B.n668 585
R651 B.n666 B.n30 585
R652 B.n30 B.n29 585
R653 B.n665 B.n664 585
R654 B.n664 B.n663 585
R655 B.n32 B.n31 585
R656 B.n662 B.n32 585
R657 B.n660 B.n659 585
R658 B.n661 B.n660 585
R659 B.n658 B.n37 585
R660 B.n37 B.n36 585
R661 B.n657 B.n656 585
R662 B.n656 B.n655 585
R663 B.n39 B.n38 585
R664 B.n654 B.n39 585
R665 B.n652 B.n651 585
R666 B.n653 B.n652 585
R667 B.n650 B.n44 585
R668 B.n44 B.n43 585
R669 B.n649 B.n648 585
R670 B.n648 B.n647 585
R671 B.n46 B.n45 585
R672 B.n646 B.n46 585
R673 B.n644 B.n643 585
R674 B.n645 B.n644 585
R675 B.n642 B.n51 585
R676 B.n51 B.n50 585
R677 B.n641 B.n640 585
R678 B.n640 B.n639 585
R679 B.n53 B.n52 585
R680 B.n638 B.n53 585
R681 B.n636 B.n635 585
R682 B.n637 B.n636 585
R683 B.n634 B.n58 585
R684 B.n58 B.n57 585
R685 B.n633 B.n632 585
R686 B.n632 B.n631 585
R687 B.n60 B.n59 585
R688 B.n630 B.n60 585
R689 B.n628 B.n627 585
R690 B.n629 B.n628 585
R691 B.n626 B.n65 585
R692 B.n65 B.n64 585
R693 B.n625 B.n624 585
R694 B.n624 B.n623 585
R695 B.n67 B.n66 585
R696 B.n622 B.n67 585
R697 B.n620 B.n619 585
R698 B.n621 B.n620 585
R699 B.n618 B.n71 585
R700 B.n74 B.n71 585
R701 B.n617 B.n616 585
R702 B.n616 B.n615 585
R703 B.n73 B.n72 585
R704 B.n614 B.n73 585
R705 B.n612 B.n611 585
R706 B.n613 B.n612 585
R707 B.n610 B.n79 585
R708 B.n79 B.n78 585
R709 B.n609 B.n608 585
R710 B.n608 B.n607 585
R711 B.n81 B.n80 585
R712 B.n606 B.n81 585
R713 B.n604 B.n603 585
R714 B.n605 B.n604 585
R715 B.n602 B.n86 585
R716 B.n86 B.n85 585
R717 B.n697 B.n696 585
R718 B.n696 B.n695 585
R719 B.n392 B.n282 506.916
R720 B.n600 B.n86 506.916
R721 B.n304 B.n280 506.916
R722 B.n596 B.n109 506.916
R723 B.n598 B.n597 256.663
R724 B.n598 B.n107 256.663
R725 B.n598 B.n106 256.663
R726 B.n598 B.n105 256.663
R727 B.n598 B.n104 256.663
R728 B.n598 B.n103 256.663
R729 B.n598 B.n102 256.663
R730 B.n598 B.n101 256.663
R731 B.n598 B.n100 256.663
R732 B.n598 B.n99 256.663
R733 B.n598 B.n98 256.663
R734 B.n598 B.n97 256.663
R735 B.n598 B.n96 256.663
R736 B.n598 B.n95 256.663
R737 B.n598 B.n94 256.663
R738 B.n598 B.n93 256.663
R739 B.n598 B.n92 256.663
R740 B.n598 B.n91 256.663
R741 B.n598 B.n90 256.663
R742 B.n598 B.n89 256.663
R743 B.n599 B.n598 256.663
R744 B.n391 B.n390 256.663
R745 B.n390 B.n285 256.663
R746 B.n390 B.n286 256.663
R747 B.n390 B.n287 256.663
R748 B.n390 B.n288 256.663
R749 B.n390 B.n289 256.663
R750 B.n390 B.n290 256.663
R751 B.n390 B.n291 256.663
R752 B.n390 B.n292 256.663
R753 B.n390 B.n293 256.663
R754 B.n390 B.n294 256.663
R755 B.n390 B.n295 256.663
R756 B.n390 B.n296 256.663
R757 B.n390 B.n297 256.663
R758 B.n390 B.n298 256.663
R759 B.n390 B.n299 256.663
R760 B.n390 B.n300 256.663
R761 B.n390 B.n301 256.663
R762 B.n390 B.n302 256.663
R763 B.n390 B.n303 256.663
R764 B.n308 B.t17 235.73
R765 B.n306 B.t10 235.73
R766 B.n113 B.t6 235.73
R767 B.n110 B.t14 235.73
R768 B.n308 B.t19 199.476
R769 B.n110 B.t15 199.476
R770 B.n306 B.t13 199.476
R771 B.n113 B.t8 199.476
R772 B.n396 B.n282 163.367
R773 B.n396 B.n276 163.367
R774 B.n404 B.n276 163.367
R775 B.n404 B.n274 163.367
R776 B.n408 B.n274 163.367
R777 B.n408 B.n268 163.367
R778 B.n417 B.n268 163.367
R779 B.n417 B.n266 163.367
R780 B.n421 B.n266 163.367
R781 B.n421 B.n261 163.367
R782 B.n429 B.n261 163.367
R783 B.n429 B.n259 163.367
R784 B.n433 B.n259 163.367
R785 B.n433 B.n253 163.367
R786 B.n441 B.n253 163.367
R787 B.n441 B.n251 163.367
R788 B.n445 B.n251 163.367
R789 B.n445 B.n245 163.367
R790 B.n453 B.n245 163.367
R791 B.n453 B.n243 163.367
R792 B.n457 B.n243 163.367
R793 B.n457 B.n237 163.367
R794 B.n465 B.n237 163.367
R795 B.n465 B.n235 163.367
R796 B.n469 B.n235 163.367
R797 B.n469 B.n229 163.367
R798 B.n477 B.n229 163.367
R799 B.n477 B.n227 163.367
R800 B.n481 B.n227 163.367
R801 B.n481 B.n221 163.367
R802 B.n489 B.n221 163.367
R803 B.n489 B.n219 163.367
R804 B.n493 B.n219 163.367
R805 B.n493 B.n213 163.367
R806 B.n501 B.n213 163.367
R807 B.n501 B.n211 163.367
R808 B.n505 B.n211 163.367
R809 B.n505 B.n205 163.367
R810 B.n514 B.n205 163.367
R811 B.n514 B.n203 163.367
R812 B.n518 B.n203 163.367
R813 B.n518 B.n198 163.367
R814 B.n527 B.n198 163.367
R815 B.n527 B.n196 163.367
R816 B.n531 B.n196 163.367
R817 B.n531 B.n2 163.367
R818 B.n696 B.n2 163.367
R819 B.n696 B.n3 163.367
R820 B.n692 B.n3 163.367
R821 B.n692 B.n9 163.367
R822 B.n688 B.n9 163.367
R823 B.n688 B.n11 163.367
R824 B.n684 B.n11 163.367
R825 B.n684 B.n15 163.367
R826 B.n680 B.n15 163.367
R827 B.n680 B.n17 163.367
R828 B.n676 B.n17 163.367
R829 B.n676 B.n23 163.367
R830 B.n672 B.n23 163.367
R831 B.n672 B.n25 163.367
R832 B.n668 B.n25 163.367
R833 B.n668 B.n30 163.367
R834 B.n664 B.n30 163.367
R835 B.n664 B.n32 163.367
R836 B.n660 B.n32 163.367
R837 B.n660 B.n37 163.367
R838 B.n656 B.n37 163.367
R839 B.n656 B.n39 163.367
R840 B.n652 B.n39 163.367
R841 B.n652 B.n44 163.367
R842 B.n648 B.n44 163.367
R843 B.n648 B.n46 163.367
R844 B.n644 B.n46 163.367
R845 B.n644 B.n51 163.367
R846 B.n640 B.n51 163.367
R847 B.n640 B.n53 163.367
R848 B.n636 B.n53 163.367
R849 B.n636 B.n58 163.367
R850 B.n632 B.n58 163.367
R851 B.n632 B.n60 163.367
R852 B.n628 B.n60 163.367
R853 B.n628 B.n65 163.367
R854 B.n624 B.n65 163.367
R855 B.n624 B.n67 163.367
R856 B.n620 B.n67 163.367
R857 B.n620 B.n71 163.367
R858 B.n616 B.n71 163.367
R859 B.n616 B.n73 163.367
R860 B.n612 B.n73 163.367
R861 B.n612 B.n79 163.367
R862 B.n608 B.n79 163.367
R863 B.n608 B.n81 163.367
R864 B.n604 B.n81 163.367
R865 B.n604 B.n86 163.367
R866 B.n389 B.n284 163.367
R867 B.n389 B.n305 163.367
R868 B.n385 B.n384 163.367
R869 B.n381 B.n380 163.367
R870 B.n377 B.n376 163.367
R871 B.n373 B.n372 163.367
R872 B.n369 B.n368 163.367
R873 B.n365 B.n364 163.367
R874 B.n360 B.n359 163.367
R875 B.n356 B.n355 163.367
R876 B.n352 B.n351 163.367
R877 B.n348 B.n347 163.367
R878 B.n344 B.n343 163.367
R879 B.n339 B.n338 163.367
R880 B.n335 B.n334 163.367
R881 B.n331 B.n330 163.367
R882 B.n327 B.n326 163.367
R883 B.n323 B.n322 163.367
R884 B.n319 B.n318 163.367
R885 B.n315 B.n314 163.367
R886 B.n311 B.n304 163.367
R887 B.n398 B.n280 163.367
R888 B.n398 B.n278 163.367
R889 B.n402 B.n278 163.367
R890 B.n402 B.n272 163.367
R891 B.n410 B.n272 163.367
R892 B.n410 B.n270 163.367
R893 B.n414 B.n270 163.367
R894 B.n414 B.n265 163.367
R895 B.n423 B.n265 163.367
R896 B.n423 B.n263 163.367
R897 B.n427 B.n263 163.367
R898 B.n427 B.n257 163.367
R899 B.n435 B.n257 163.367
R900 B.n435 B.n255 163.367
R901 B.n439 B.n255 163.367
R902 B.n439 B.n249 163.367
R903 B.n447 B.n249 163.367
R904 B.n447 B.n247 163.367
R905 B.n451 B.n247 163.367
R906 B.n451 B.n241 163.367
R907 B.n459 B.n241 163.367
R908 B.n459 B.n239 163.367
R909 B.n463 B.n239 163.367
R910 B.n463 B.n233 163.367
R911 B.n471 B.n233 163.367
R912 B.n471 B.n231 163.367
R913 B.n475 B.n231 163.367
R914 B.n475 B.n224 163.367
R915 B.n483 B.n224 163.367
R916 B.n483 B.n222 163.367
R917 B.n487 B.n222 163.367
R918 B.n487 B.n217 163.367
R919 B.n495 B.n217 163.367
R920 B.n495 B.n215 163.367
R921 B.n499 B.n215 163.367
R922 B.n499 B.n209 163.367
R923 B.n507 B.n209 163.367
R924 B.n507 B.n207 163.367
R925 B.n511 B.n207 163.367
R926 B.n511 B.n202 163.367
R927 B.n520 B.n202 163.367
R928 B.n520 B.n200 163.367
R929 B.n525 B.n200 163.367
R930 B.n525 B.n194 163.367
R931 B.n533 B.n194 163.367
R932 B.n534 B.n533 163.367
R933 B.n534 B.n5 163.367
R934 B.n6 B.n5 163.367
R935 B.n7 B.n6 163.367
R936 B.n539 B.n7 163.367
R937 B.n539 B.n12 163.367
R938 B.n13 B.n12 163.367
R939 B.n14 B.n13 163.367
R940 B.n544 B.n14 163.367
R941 B.n544 B.n19 163.367
R942 B.n20 B.n19 163.367
R943 B.n21 B.n20 163.367
R944 B.n549 B.n21 163.367
R945 B.n549 B.n26 163.367
R946 B.n27 B.n26 163.367
R947 B.n28 B.n27 163.367
R948 B.n554 B.n28 163.367
R949 B.n554 B.n33 163.367
R950 B.n34 B.n33 163.367
R951 B.n35 B.n34 163.367
R952 B.n559 B.n35 163.367
R953 B.n559 B.n40 163.367
R954 B.n41 B.n40 163.367
R955 B.n42 B.n41 163.367
R956 B.n564 B.n42 163.367
R957 B.n564 B.n47 163.367
R958 B.n48 B.n47 163.367
R959 B.n49 B.n48 163.367
R960 B.n569 B.n49 163.367
R961 B.n569 B.n54 163.367
R962 B.n55 B.n54 163.367
R963 B.n56 B.n55 163.367
R964 B.n574 B.n56 163.367
R965 B.n574 B.n61 163.367
R966 B.n62 B.n61 163.367
R967 B.n63 B.n62 163.367
R968 B.n579 B.n63 163.367
R969 B.n579 B.n68 163.367
R970 B.n69 B.n68 163.367
R971 B.n70 B.n69 163.367
R972 B.n584 B.n70 163.367
R973 B.n584 B.n75 163.367
R974 B.n76 B.n75 163.367
R975 B.n77 B.n76 163.367
R976 B.n589 B.n77 163.367
R977 B.n589 B.n82 163.367
R978 B.n83 B.n82 163.367
R979 B.n84 B.n83 163.367
R980 B.n109 B.n84 163.367
R981 B.n116 B.n88 163.367
R982 B.n120 B.n119 163.367
R983 B.n124 B.n123 163.367
R984 B.n128 B.n127 163.367
R985 B.n132 B.n131 163.367
R986 B.n136 B.n135 163.367
R987 B.n140 B.n139 163.367
R988 B.n144 B.n143 163.367
R989 B.n148 B.n147 163.367
R990 B.n152 B.n151 163.367
R991 B.n156 B.n155 163.367
R992 B.n160 B.n159 163.367
R993 B.n164 B.n163 163.367
R994 B.n168 B.n167 163.367
R995 B.n172 B.n171 163.367
R996 B.n176 B.n175 163.367
R997 B.n180 B.n179 163.367
R998 B.n184 B.n183 163.367
R999 B.n188 B.n187 163.367
R1000 B.n190 B.n108 163.367
R1001 B.n390 B.n281 161.784
R1002 B.n598 B.n85 161.784
R1003 B.n309 B.t18 135.282
R1004 B.n111 B.t16 135.282
R1005 B.n307 B.t12 135.282
R1006 B.n114 B.t9 135.282
R1007 B.n397 B.n281 86.6247
R1008 B.n397 B.n277 86.6247
R1009 B.n403 B.n277 86.6247
R1010 B.n403 B.n273 86.6247
R1011 B.n409 B.n273 86.6247
R1012 B.n409 B.n269 86.6247
R1013 B.n416 B.n269 86.6247
R1014 B.n416 B.n415 86.6247
R1015 B.n422 B.n262 86.6247
R1016 B.n428 B.n262 86.6247
R1017 B.n428 B.n258 86.6247
R1018 B.n434 B.n258 86.6247
R1019 B.n434 B.n254 86.6247
R1020 B.n440 B.n254 86.6247
R1021 B.n440 B.n250 86.6247
R1022 B.n446 B.n250 86.6247
R1023 B.n446 B.n246 86.6247
R1024 B.n452 B.n246 86.6247
R1025 B.n452 B.n242 86.6247
R1026 B.n458 B.n242 86.6247
R1027 B.n464 B.n238 86.6247
R1028 B.n464 B.n234 86.6247
R1029 B.n470 B.n234 86.6247
R1030 B.n470 B.n230 86.6247
R1031 B.n476 B.n230 86.6247
R1032 B.n476 B.n225 86.6247
R1033 B.n482 B.n225 86.6247
R1034 B.n482 B.n226 86.6247
R1035 B.n488 B.n218 86.6247
R1036 B.n494 B.n218 86.6247
R1037 B.n494 B.n214 86.6247
R1038 B.n500 B.n214 86.6247
R1039 B.n500 B.n210 86.6247
R1040 B.n506 B.n210 86.6247
R1041 B.n506 B.n206 86.6247
R1042 B.n513 B.n206 86.6247
R1043 B.n513 B.n512 86.6247
R1044 B.n519 B.n199 86.6247
R1045 B.n526 B.n199 86.6247
R1046 B.n526 B.n195 86.6247
R1047 B.n532 B.n195 86.6247
R1048 B.n532 B.n4 86.6247
R1049 B.n695 B.n4 86.6247
R1050 B.n695 B.n694 86.6247
R1051 B.n694 B.n693 86.6247
R1052 B.n693 B.n8 86.6247
R1053 B.n687 B.n8 86.6247
R1054 B.n687 B.n686 86.6247
R1055 B.n686 B.n685 86.6247
R1056 B.n679 B.n18 86.6247
R1057 B.n679 B.n678 86.6247
R1058 B.n678 B.n677 86.6247
R1059 B.n677 B.n22 86.6247
R1060 B.n671 B.n22 86.6247
R1061 B.n671 B.n670 86.6247
R1062 B.n670 B.n669 86.6247
R1063 B.n669 B.n29 86.6247
R1064 B.n663 B.n29 86.6247
R1065 B.n662 B.n661 86.6247
R1066 B.n661 B.n36 86.6247
R1067 B.n655 B.n36 86.6247
R1068 B.n655 B.n654 86.6247
R1069 B.n654 B.n653 86.6247
R1070 B.n653 B.n43 86.6247
R1071 B.n647 B.n43 86.6247
R1072 B.n647 B.n646 86.6247
R1073 B.n645 B.n50 86.6247
R1074 B.n639 B.n50 86.6247
R1075 B.n639 B.n638 86.6247
R1076 B.n638 B.n637 86.6247
R1077 B.n637 B.n57 86.6247
R1078 B.n631 B.n57 86.6247
R1079 B.n631 B.n630 86.6247
R1080 B.n630 B.n629 86.6247
R1081 B.n629 B.n64 86.6247
R1082 B.n623 B.n64 86.6247
R1083 B.n623 B.n622 86.6247
R1084 B.n622 B.n621 86.6247
R1085 B.n615 B.n74 86.6247
R1086 B.n615 B.n614 86.6247
R1087 B.n614 B.n613 86.6247
R1088 B.n613 B.n78 86.6247
R1089 B.n607 B.n78 86.6247
R1090 B.n607 B.n606 86.6247
R1091 B.n606 B.n605 86.6247
R1092 B.n605 B.n85 86.6247
R1093 B.t4 B.n238 81.5292
R1094 B.n646 B.t5 81.5292
R1095 B.n422 B.t11 76.4336
R1096 B.n621 B.t7 76.4336
R1097 B.n392 B.n391 71.676
R1098 B.n305 B.n285 71.676
R1099 B.n384 B.n286 71.676
R1100 B.n380 B.n287 71.676
R1101 B.n376 B.n288 71.676
R1102 B.n372 B.n289 71.676
R1103 B.n368 B.n290 71.676
R1104 B.n364 B.n291 71.676
R1105 B.n359 B.n292 71.676
R1106 B.n355 B.n293 71.676
R1107 B.n351 B.n294 71.676
R1108 B.n347 B.n295 71.676
R1109 B.n343 B.n296 71.676
R1110 B.n338 B.n297 71.676
R1111 B.n334 B.n298 71.676
R1112 B.n330 B.n299 71.676
R1113 B.n326 B.n300 71.676
R1114 B.n322 B.n301 71.676
R1115 B.n318 B.n302 71.676
R1116 B.n314 B.n303 71.676
R1117 B.n600 B.n599 71.676
R1118 B.n116 B.n89 71.676
R1119 B.n120 B.n90 71.676
R1120 B.n124 B.n91 71.676
R1121 B.n128 B.n92 71.676
R1122 B.n132 B.n93 71.676
R1123 B.n136 B.n94 71.676
R1124 B.n140 B.n95 71.676
R1125 B.n144 B.n96 71.676
R1126 B.n148 B.n97 71.676
R1127 B.n152 B.n98 71.676
R1128 B.n156 B.n99 71.676
R1129 B.n160 B.n100 71.676
R1130 B.n164 B.n101 71.676
R1131 B.n168 B.n102 71.676
R1132 B.n172 B.n103 71.676
R1133 B.n176 B.n104 71.676
R1134 B.n180 B.n105 71.676
R1135 B.n184 B.n106 71.676
R1136 B.n188 B.n107 71.676
R1137 B.n597 B.n108 71.676
R1138 B.n597 B.n596 71.676
R1139 B.n190 B.n107 71.676
R1140 B.n187 B.n106 71.676
R1141 B.n183 B.n105 71.676
R1142 B.n179 B.n104 71.676
R1143 B.n175 B.n103 71.676
R1144 B.n171 B.n102 71.676
R1145 B.n167 B.n101 71.676
R1146 B.n163 B.n100 71.676
R1147 B.n159 B.n99 71.676
R1148 B.n155 B.n98 71.676
R1149 B.n151 B.n97 71.676
R1150 B.n147 B.n96 71.676
R1151 B.n143 B.n95 71.676
R1152 B.n139 B.n94 71.676
R1153 B.n135 B.n93 71.676
R1154 B.n131 B.n92 71.676
R1155 B.n127 B.n91 71.676
R1156 B.n123 B.n90 71.676
R1157 B.n119 B.n89 71.676
R1158 B.n599 B.n88 71.676
R1159 B.n391 B.n284 71.676
R1160 B.n385 B.n285 71.676
R1161 B.n381 B.n286 71.676
R1162 B.n377 B.n287 71.676
R1163 B.n373 B.n288 71.676
R1164 B.n369 B.n289 71.676
R1165 B.n365 B.n290 71.676
R1166 B.n360 B.n291 71.676
R1167 B.n356 B.n292 71.676
R1168 B.n352 B.n293 71.676
R1169 B.n348 B.n294 71.676
R1170 B.n344 B.n295 71.676
R1171 B.n339 B.n296 71.676
R1172 B.n335 B.n297 71.676
R1173 B.n331 B.n298 71.676
R1174 B.n327 B.n299 71.676
R1175 B.n323 B.n300 71.676
R1176 B.n319 B.n301 71.676
R1177 B.n315 B.n302 71.676
R1178 B.n311 B.n303 71.676
R1179 B.n226 B.t0 68.7903
R1180 B.t3 B.n662 68.7903
R1181 B.n309 B.n308 64.1944
R1182 B.n307 B.n306 64.1944
R1183 B.n114 B.n113 64.1944
R1184 B.n111 B.n110 64.1944
R1185 B.n341 B.n309 59.5399
R1186 B.n362 B.n307 59.5399
R1187 B.n115 B.n114 59.5399
R1188 B.n112 B.n111 59.5399
R1189 B.n512 B.t2 45.8604
R1190 B.n18 B.t1 45.8604
R1191 B.n519 B.t2 40.7648
R1192 B.n685 B.t1 40.7648
R1193 B.n602 B.n601 32.9371
R1194 B.n595 B.n594 32.9371
R1195 B.n310 B.n279 32.9371
R1196 B.n394 B.n393 32.9371
R1197 B B.n697 18.0485
R1198 B.n488 B.t0 17.8349
R1199 B.n663 B.t3 17.8349
R1200 B.n601 B.n87 10.6151
R1201 B.n117 B.n87 10.6151
R1202 B.n118 B.n117 10.6151
R1203 B.n121 B.n118 10.6151
R1204 B.n122 B.n121 10.6151
R1205 B.n125 B.n122 10.6151
R1206 B.n126 B.n125 10.6151
R1207 B.n129 B.n126 10.6151
R1208 B.n130 B.n129 10.6151
R1209 B.n133 B.n130 10.6151
R1210 B.n134 B.n133 10.6151
R1211 B.n137 B.n134 10.6151
R1212 B.n138 B.n137 10.6151
R1213 B.n141 B.n138 10.6151
R1214 B.n142 B.n141 10.6151
R1215 B.n146 B.n145 10.6151
R1216 B.n149 B.n146 10.6151
R1217 B.n150 B.n149 10.6151
R1218 B.n153 B.n150 10.6151
R1219 B.n154 B.n153 10.6151
R1220 B.n157 B.n154 10.6151
R1221 B.n158 B.n157 10.6151
R1222 B.n161 B.n158 10.6151
R1223 B.n162 B.n161 10.6151
R1224 B.n166 B.n165 10.6151
R1225 B.n169 B.n166 10.6151
R1226 B.n170 B.n169 10.6151
R1227 B.n173 B.n170 10.6151
R1228 B.n174 B.n173 10.6151
R1229 B.n177 B.n174 10.6151
R1230 B.n178 B.n177 10.6151
R1231 B.n181 B.n178 10.6151
R1232 B.n182 B.n181 10.6151
R1233 B.n185 B.n182 10.6151
R1234 B.n186 B.n185 10.6151
R1235 B.n189 B.n186 10.6151
R1236 B.n191 B.n189 10.6151
R1237 B.n192 B.n191 10.6151
R1238 B.n595 B.n192 10.6151
R1239 B.n399 B.n279 10.6151
R1240 B.n400 B.n399 10.6151
R1241 B.n401 B.n400 10.6151
R1242 B.n401 B.n271 10.6151
R1243 B.n411 B.n271 10.6151
R1244 B.n412 B.n411 10.6151
R1245 B.n413 B.n412 10.6151
R1246 B.n413 B.n264 10.6151
R1247 B.n424 B.n264 10.6151
R1248 B.n425 B.n424 10.6151
R1249 B.n426 B.n425 10.6151
R1250 B.n426 B.n256 10.6151
R1251 B.n436 B.n256 10.6151
R1252 B.n437 B.n436 10.6151
R1253 B.n438 B.n437 10.6151
R1254 B.n438 B.n248 10.6151
R1255 B.n448 B.n248 10.6151
R1256 B.n449 B.n448 10.6151
R1257 B.n450 B.n449 10.6151
R1258 B.n450 B.n240 10.6151
R1259 B.n460 B.n240 10.6151
R1260 B.n461 B.n460 10.6151
R1261 B.n462 B.n461 10.6151
R1262 B.n462 B.n232 10.6151
R1263 B.n472 B.n232 10.6151
R1264 B.n473 B.n472 10.6151
R1265 B.n474 B.n473 10.6151
R1266 B.n474 B.n223 10.6151
R1267 B.n484 B.n223 10.6151
R1268 B.n485 B.n484 10.6151
R1269 B.n486 B.n485 10.6151
R1270 B.n486 B.n216 10.6151
R1271 B.n496 B.n216 10.6151
R1272 B.n497 B.n496 10.6151
R1273 B.n498 B.n497 10.6151
R1274 B.n498 B.n208 10.6151
R1275 B.n508 B.n208 10.6151
R1276 B.n509 B.n508 10.6151
R1277 B.n510 B.n509 10.6151
R1278 B.n510 B.n201 10.6151
R1279 B.n521 B.n201 10.6151
R1280 B.n522 B.n521 10.6151
R1281 B.n524 B.n522 10.6151
R1282 B.n524 B.n523 10.6151
R1283 B.n523 B.n193 10.6151
R1284 B.n535 B.n193 10.6151
R1285 B.n536 B.n535 10.6151
R1286 B.n537 B.n536 10.6151
R1287 B.n538 B.n537 10.6151
R1288 B.n540 B.n538 10.6151
R1289 B.n541 B.n540 10.6151
R1290 B.n542 B.n541 10.6151
R1291 B.n543 B.n542 10.6151
R1292 B.n545 B.n543 10.6151
R1293 B.n546 B.n545 10.6151
R1294 B.n547 B.n546 10.6151
R1295 B.n548 B.n547 10.6151
R1296 B.n550 B.n548 10.6151
R1297 B.n551 B.n550 10.6151
R1298 B.n552 B.n551 10.6151
R1299 B.n553 B.n552 10.6151
R1300 B.n555 B.n553 10.6151
R1301 B.n556 B.n555 10.6151
R1302 B.n557 B.n556 10.6151
R1303 B.n558 B.n557 10.6151
R1304 B.n560 B.n558 10.6151
R1305 B.n561 B.n560 10.6151
R1306 B.n562 B.n561 10.6151
R1307 B.n563 B.n562 10.6151
R1308 B.n565 B.n563 10.6151
R1309 B.n566 B.n565 10.6151
R1310 B.n567 B.n566 10.6151
R1311 B.n568 B.n567 10.6151
R1312 B.n570 B.n568 10.6151
R1313 B.n571 B.n570 10.6151
R1314 B.n572 B.n571 10.6151
R1315 B.n573 B.n572 10.6151
R1316 B.n575 B.n573 10.6151
R1317 B.n576 B.n575 10.6151
R1318 B.n577 B.n576 10.6151
R1319 B.n578 B.n577 10.6151
R1320 B.n580 B.n578 10.6151
R1321 B.n581 B.n580 10.6151
R1322 B.n582 B.n581 10.6151
R1323 B.n583 B.n582 10.6151
R1324 B.n585 B.n583 10.6151
R1325 B.n586 B.n585 10.6151
R1326 B.n587 B.n586 10.6151
R1327 B.n588 B.n587 10.6151
R1328 B.n590 B.n588 10.6151
R1329 B.n591 B.n590 10.6151
R1330 B.n592 B.n591 10.6151
R1331 B.n593 B.n592 10.6151
R1332 B.n594 B.n593 10.6151
R1333 B.n393 B.n283 10.6151
R1334 B.n388 B.n283 10.6151
R1335 B.n388 B.n387 10.6151
R1336 B.n387 B.n386 10.6151
R1337 B.n386 B.n383 10.6151
R1338 B.n383 B.n382 10.6151
R1339 B.n382 B.n379 10.6151
R1340 B.n379 B.n378 10.6151
R1341 B.n378 B.n375 10.6151
R1342 B.n375 B.n374 10.6151
R1343 B.n374 B.n371 10.6151
R1344 B.n371 B.n370 10.6151
R1345 B.n370 B.n367 10.6151
R1346 B.n367 B.n366 10.6151
R1347 B.n366 B.n363 10.6151
R1348 B.n361 B.n358 10.6151
R1349 B.n358 B.n357 10.6151
R1350 B.n357 B.n354 10.6151
R1351 B.n354 B.n353 10.6151
R1352 B.n353 B.n350 10.6151
R1353 B.n350 B.n349 10.6151
R1354 B.n349 B.n346 10.6151
R1355 B.n346 B.n345 10.6151
R1356 B.n345 B.n342 10.6151
R1357 B.n340 B.n337 10.6151
R1358 B.n337 B.n336 10.6151
R1359 B.n336 B.n333 10.6151
R1360 B.n333 B.n332 10.6151
R1361 B.n332 B.n329 10.6151
R1362 B.n329 B.n328 10.6151
R1363 B.n328 B.n325 10.6151
R1364 B.n325 B.n324 10.6151
R1365 B.n324 B.n321 10.6151
R1366 B.n321 B.n320 10.6151
R1367 B.n320 B.n317 10.6151
R1368 B.n317 B.n316 10.6151
R1369 B.n316 B.n313 10.6151
R1370 B.n313 B.n312 10.6151
R1371 B.n312 B.n310 10.6151
R1372 B.n395 B.n394 10.6151
R1373 B.n395 B.n275 10.6151
R1374 B.n405 B.n275 10.6151
R1375 B.n406 B.n405 10.6151
R1376 B.n407 B.n406 10.6151
R1377 B.n407 B.n267 10.6151
R1378 B.n418 B.n267 10.6151
R1379 B.n419 B.n418 10.6151
R1380 B.n420 B.n419 10.6151
R1381 B.n420 B.n260 10.6151
R1382 B.n430 B.n260 10.6151
R1383 B.n431 B.n430 10.6151
R1384 B.n432 B.n431 10.6151
R1385 B.n432 B.n252 10.6151
R1386 B.n442 B.n252 10.6151
R1387 B.n443 B.n442 10.6151
R1388 B.n444 B.n443 10.6151
R1389 B.n444 B.n244 10.6151
R1390 B.n454 B.n244 10.6151
R1391 B.n455 B.n454 10.6151
R1392 B.n456 B.n455 10.6151
R1393 B.n456 B.n236 10.6151
R1394 B.n466 B.n236 10.6151
R1395 B.n467 B.n466 10.6151
R1396 B.n468 B.n467 10.6151
R1397 B.n468 B.n228 10.6151
R1398 B.n478 B.n228 10.6151
R1399 B.n479 B.n478 10.6151
R1400 B.n480 B.n479 10.6151
R1401 B.n480 B.n220 10.6151
R1402 B.n490 B.n220 10.6151
R1403 B.n491 B.n490 10.6151
R1404 B.n492 B.n491 10.6151
R1405 B.n492 B.n212 10.6151
R1406 B.n502 B.n212 10.6151
R1407 B.n503 B.n502 10.6151
R1408 B.n504 B.n503 10.6151
R1409 B.n504 B.n204 10.6151
R1410 B.n515 B.n204 10.6151
R1411 B.n516 B.n515 10.6151
R1412 B.n517 B.n516 10.6151
R1413 B.n517 B.n197 10.6151
R1414 B.n528 B.n197 10.6151
R1415 B.n529 B.n528 10.6151
R1416 B.n530 B.n529 10.6151
R1417 B.n530 B.n0 10.6151
R1418 B.n691 B.n1 10.6151
R1419 B.n691 B.n690 10.6151
R1420 B.n690 B.n689 10.6151
R1421 B.n689 B.n10 10.6151
R1422 B.n683 B.n10 10.6151
R1423 B.n683 B.n682 10.6151
R1424 B.n682 B.n681 10.6151
R1425 B.n681 B.n16 10.6151
R1426 B.n675 B.n16 10.6151
R1427 B.n675 B.n674 10.6151
R1428 B.n674 B.n673 10.6151
R1429 B.n673 B.n24 10.6151
R1430 B.n667 B.n24 10.6151
R1431 B.n667 B.n666 10.6151
R1432 B.n666 B.n665 10.6151
R1433 B.n665 B.n31 10.6151
R1434 B.n659 B.n31 10.6151
R1435 B.n659 B.n658 10.6151
R1436 B.n658 B.n657 10.6151
R1437 B.n657 B.n38 10.6151
R1438 B.n651 B.n38 10.6151
R1439 B.n651 B.n650 10.6151
R1440 B.n650 B.n649 10.6151
R1441 B.n649 B.n45 10.6151
R1442 B.n643 B.n45 10.6151
R1443 B.n643 B.n642 10.6151
R1444 B.n642 B.n641 10.6151
R1445 B.n641 B.n52 10.6151
R1446 B.n635 B.n52 10.6151
R1447 B.n635 B.n634 10.6151
R1448 B.n634 B.n633 10.6151
R1449 B.n633 B.n59 10.6151
R1450 B.n627 B.n59 10.6151
R1451 B.n627 B.n626 10.6151
R1452 B.n626 B.n625 10.6151
R1453 B.n625 B.n66 10.6151
R1454 B.n619 B.n66 10.6151
R1455 B.n619 B.n618 10.6151
R1456 B.n618 B.n617 10.6151
R1457 B.n617 B.n72 10.6151
R1458 B.n611 B.n72 10.6151
R1459 B.n611 B.n610 10.6151
R1460 B.n610 B.n609 10.6151
R1461 B.n609 B.n80 10.6151
R1462 B.n603 B.n80 10.6151
R1463 B.n603 B.n602 10.6151
R1464 B.n415 B.t11 10.1916
R1465 B.n74 B.t7 10.1916
R1466 B.n142 B.n115 9.36635
R1467 B.n165 B.n112 9.36635
R1468 B.n363 B.n362 9.36635
R1469 B.n341 B.n340 9.36635
R1470 B.n458 B.t4 5.09604
R1471 B.t5 B.n645 5.09604
R1472 B.n697 B.n0 2.81026
R1473 B.n697 B.n1 2.81026
R1474 B.n145 B.n115 1.24928
R1475 B.n162 B.n112 1.24928
R1476 B.n362 B.n361 1.24928
R1477 B.n342 B.n341 1.24928
R1478 VN.n33 VN.n18 161.3
R1479 VN.n32 VN.n31 161.3
R1480 VN.n30 VN.n19 161.3
R1481 VN.n29 VN.n28 161.3
R1482 VN.n27 VN.n20 161.3
R1483 VN.n26 VN.n25 161.3
R1484 VN.n24 VN.n21 161.3
R1485 VN.n15 VN.n0 161.3
R1486 VN.n14 VN.n13 161.3
R1487 VN.n12 VN.n1 161.3
R1488 VN.n11 VN.n10 161.3
R1489 VN.n9 VN.n2 161.3
R1490 VN.n8 VN.n7 161.3
R1491 VN.n6 VN.n3 161.3
R1492 VN.n17 VN.n16 107.957
R1493 VN.n35 VN.n34 107.957
R1494 VN.n5 VN.n4 61.8105
R1495 VN.n23 VN.n22 61.8105
R1496 VN.n5 VN.t4 60.2918
R1497 VN.n23 VN.t3 60.2918
R1498 VN.n10 VN.n9 49.7803
R1499 VN.n28 VN.n27 49.7803
R1500 VN VN.n35 43.9035
R1501 VN.n10 VN.n1 31.3737
R1502 VN.n28 VN.n19 31.3737
R1503 VN.n4 VN.t1 27.1737
R1504 VN.n16 VN.t2 27.1737
R1505 VN.n22 VN.t5 27.1737
R1506 VN.n34 VN.t0 27.1737
R1507 VN.n8 VN.n3 24.5923
R1508 VN.n9 VN.n8 24.5923
R1509 VN.n14 VN.n1 24.5923
R1510 VN.n15 VN.n14 24.5923
R1511 VN.n27 VN.n26 24.5923
R1512 VN.n26 VN.n21 24.5923
R1513 VN.n33 VN.n32 24.5923
R1514 VN.n32 VN.n19 24.5923
R1515 VN.n4 VN.n3 12.2964
R1516 VN.n22 VN.n21 12.2964
R1517 VN.n24 VN.n23 5.06578
R1518 VN.n6 VN.n5 5.06578
R1519 VN.n16 VN.n15 2.95152
R1520 VN.n34 VN.n33 2.95152
R1521 VN.n35 VN.n18 0.278335
R1522 VN.n17 VN.n0 0.278335
R1523 VN.n31 VN.n18 0.189894
R1524 VN.n31 VN.n30 0.189894
R1525 VN.n30 VN.n29 0.189894
R1526 VN.n29 VN.n20 0.189894
R1527 VN.n25 VN.n20 0.189894
R1528 VN.n25 VN.n24 0.189894
R1529 VN.n7 VN.n6 0.189894
R1530 VN.n7 VN.n2 0.189894
R1531 VN.n11 VN.n2 0.189894
R1532 VN.n12 VN.n11 0.189894
R1533 VN.n13 VN.n12 0.189894
R1534 VN.n13 VN.n0 0.189894
R1535 VN VN.n17 0.153485
R1536 VDD2.n27 VDD2.n17 289.615
R1537 VDD2.n10 VDD2.n0 289.615
R1538 VDD2.n28 VDD2.n27 185
R1539 VDD2.n26 VDD2.n25 185
R1540 VDD2.n21 VDD2.n20 185
R1541 VDD2.n4 VDD2.n3 185
R1542 VDD2.n9 VDD2.n8 185
R1543 VDD2.n11 VDD2.n10 185
R1544 VDD2.n22 VDD2.t5 150.499
R1545 VDD2.n5 VDD2.t1 150.499
R1546 VDD2.n27 VDD2.n26 104.615
R1547 VDD2.n26 VDD2.n20 104.615
R1548 VDD2.n9 VDD2.n3 104.615
R1549 VDD2.n10 VDD2.n9 104.615
R1550 VDD2.n16 VDD2.n15 77.2016
R1551 VDD2 VDD2.n33 77.1988
R1552 VDD2.t5 VDD2.n20 52.3082
R1553 VDD2.t1 VDD2.n3 52.3082
R1554 VDD2.n16 VDD2.n14 48.6216
R1555 VDD2.n32 VDD2.n31 46.5369
R1556 VDD2.n32 VDD2.n16 35.8856
R1557 VDD2.n22 VDD2.n21 10.2326
R1558 VDD2.n5 VDD2.n4 10.2326
R1559 VDD2.n31 VDD2.n17 9.69747
R1560 VDD2.n14 VDD2.n0 9.69747
R1561 VDD2.n31 VDD2.n30 9.45567
R1562 VDD2.n14 VDD2.n13 9.45567
R1563 VDD2.n19 VDD2.n18 9.3005
R1564 VDD2.n30 VDD2.n29 9.3005
R1565 VDD2.n24 VDD2.n23 9.3005
R1566 VDD2.n7 VDD2.n6 9.3005
R1567 VDD2.n2 VDD2.n1 9.3005
R1568 VDD2.n13 VDD2.n12 9.3005
R1569 VDD2.n29 VDD2.n28 8.92171
R1570 VDD2.n12 VDD2.n11 8.92171
R1571 VDD2.n25 VDD2.n19 8.14595
R1572 VDD2.n8 VDD2.n2 8.14595
R1573 VDD2.n24 VDD2.n21 7.3702
R1574 VDD2.n7 VDD2.n4 7.3702
R1575 VDD2.n33 VDD2.t0 5.89336
R1576 VDD2.n33 VDD2.t2 5.89336
R1577 VDD2.n15 VDD2.t4 5.89336
R1578 VDD2.n15 VDD2.t3 5.89336
R1579 VDD2.n25 VDD2.n24 5.81868
R1580 VDD2.n8 VDD2.n7 5.81868
R1581 VDD2.n28 VDD2.n19 5.04292
R1582 VDD2.n11 VDD2.n2 5.04292
R1583 VDD2.n29 VDD2.n17 4.26717
R1584 VDD2.n12 VDD2.n0 4.26717
R1585 VDD2.n23 VDD2.n22 2.88718
R1586 VDD2.n6 VDD2.n5 2.88718
R1587 VDD2 VDD2.n32 2.19878
R1588 VDD2.n30 VDD2.n18 0.155672
R1589 VDD2.n23 VDD2.n18 0.155672
R1590 VDD2.n6 VDD2.n1 0.155672
R1591 VDD2.n13 VDD2.n1 0.155672
C0 VTAIL VP 3.0872f
C1 VTAIL VDD1 4.84137f
C2 VDD2 VN 2.21472f
C3 VP VDD2 0.495661f
C4 VP VN 5.694241f
C5 VDD2 VDD1 1.55396f
C6 VTAIL VDD2 4.89687f
C7 VN VDD1 0.156337f
C8 VTAIL VN 3.07306f
C9 VP VDD1 2.55147f
C10 VDD2 B 4.744983f
C11 VDD1 B 4.886579f
C12 VTAIL B 4.192651f
C13 VN B 13.2206f
C14 VP B 11.832218f
C15 VDD2.n0 B 0.032504f
C16 VDD2.n1 B 0.02227f
C17 VDD2.n2 B 0.011967f
C18 VDD2.n3 B 0.021214f
C19 VDD2.n4 B 0.019804f
C20 VDD2.t1 B 0.049406f
C21 VDD2.n5 B 0.089535f
C22 VDD2.n6 B 0.262335f
C23 VDD2.n7 B 0.011967f
C24 VDD2.n8 B 0.012671f
C25 VDD2.n9 B 0.028285f
C26 VDD2.n10 B 0.063359f
C27 VDD2.n11 B 0.012671f
C28 VDD2.n12 B 0.011967f
C29 VDD2.n13 B 0.047825f
C30 VDD2.n14 B 0.059137f
C31 VDD2.t4 B 0.059131f
C32 VDD2.t3 B 0.059131f
C33 VDD2.n15 B 0.442296f
C34 VDD2.n16 B 2.06417f
C35 VDD2.n17 B 0.032504f
C36 VDD2.n18 B 0.02227f
C37 VDD2.n19 B 0.011967f
C38 VDD2.n20 B 0.021214f
C39 VDD2.n21 B 0.019804f
C40 VDD2.t5 B 0.049406f
C41 VDD2.n22 B 0.089535f
C42 VDD2.n23 B 0.262335f
C43 VDD2.n24 B 0.011967f
C44 VDD2.n25 B 0.012671f
C45 VDD2.n26 B 0.028285f
C46 VDD2.n27 B 0.063359f
C47 VDD2.n28 B 0.012671f
C48 VDD2.n29 B 0.011967f
C49 VDD2.n30 B 0.047825f
C50 VDD2.n31 B 0.050963f
C51 VDD2.n32 B 1.76654f
C52 VDD2.t0 B 0.059131f
C53 VDD2.t2 B 0.059131f
C54 VDD2.n33 B 0.442272f
C55 VN.n0 B 0.036262f
C56 VN.t2 B 0.695268f
C57 VN.n1 B 0.054927f
C58 VN.n2 B 0.027506f
C59 VN.n3 B 0.038417f
C60 VN.t4 B 0.95451f
C61 VN.t1 B 0.695268f
C62 VN.n4 B 0.368965f
C63 VN.n5 B 0.357327f
C64 VN.n6 B 0.294095f
C65 VN.n7 B 0.027506f
C66 VN.n8 B 0.051008f
C67 VN.n9 B 0.050498f
C68 VN.n10 B 0.025552f
C69 VN.n11 B 0.027506f
C70 VN.n12 B 0.027506f
C71 VN.n13 B 0.027506f
C72 VN.n14 B 0.051008f
C73 VN.n15 B 0.028848f
C74 VN.n16 B 0.377179f
C75 VN.n17 B 0.053215f
C76 VN.n18 B 0.036262f
C77 VN.t0 B 0.695268f
C78 VN.n19 B 0.054927f
C79 VN.n20 B 0.027506f
C80 VN.n21 B 0.038417f
C81 VN.t3 B 0.95451f
C82 VN.t5 B 0.695268f
C83 VN.n22 B 0.368965f
C84 VN.n23 B 0.357327f
C85 VN.n24 B 0.294095f
C86 VN.n25 B 0.027506f
C87 VN.n26 B 0.051008f
C88 VN.n27 B 0.050498f
C89 VN.n28 B 0.025552f
C90 VN.n29 B 0.027506f
C91 VN.n30 B 0.027506f
C92 VN.n31 B 0.027506f
C93 VN.n32 B 0.051008f
C94 VN.n33 B 0.028848f
C95 VN.n34 B 0.377179f
C96 VN.n35 B 1.26776f
C97 VTAIL.t1 B 0.083328f
C98 VTAIL.t3 B 0.083328f
C99 VTAIL.n0 B 0.548664f
C100 VTAIL.n1 B 0.551223f
C101 VTAIL.n2 B 0.045806f
C102 VTAIL.n3 B 0.031383f
C103 VTAIL.n4 B 0.016864f
C104 VTAIL.n5 B 0.029895f
C105 VTAIL.n6 B 0.027909f
C106 VTAIL.t7 B 0.069624f
C107 VTAIL.n7 B 0.126174f
C108 VTAIL.n8 B 0.369689f
C109 VTAIL.n9 B 0.016864f
C110 VTAIL.n10 B 0.017856f
C111 VTAIL.n11 B 0.03986f
C112 VTAIL.n12 B 0.089286f
C113 VTAIL.n13 B 0.017856f
C114 VTAIL.n14 B 0.016864f
C115 VTAIL.n15 B 0.067396f
C116 VTAIL.n16 B 0.050103f
C117 VTAIL.n17 B 0.504243f
C118 VTAIL.t8 B 0.083328f
C119 VTAIL.t9 B 0.083328f
C120 VTAIL.n18 B 0.548664f
C121 VTAIL.n19 B 1.86628f
C122 VTAIL.t4 B 0.083328f
C123 VTAIL.t0 B 0.083328f
C124 VTAIL.n20 B 0.548667f
C125 VTAIL.n21 B 1.86628f
C126 VTAIL.n22 B 0.045806f
C127 VTAIL.n23 B 0.031383f
C128 VTAIL.n24 B 0.016864f
C129 VTAIL.n25 B 0.029895f
C130 VTAIL.n26 B 0.027909f
C131 VTAIL.t2 B 0.069624f
C132 VTAIL.n27 B 0.126174f
C133 VTAIL.n28 B 0.369689f
C134 VTAIL.n29 B 0.016864f
C135 VTAIL.n30 B 0.017856f
C136 VTAIL.n31 B 0.03986f
C137 VTAIL.n32 B 0.089286f
C138 VTAIL.n33 B 0.017856f
C139 VTAIL.n34 B 0.016864f
C140 VTAIL.n35 B 0.067396f
C141 VTAIL.n36 B 0.050103f
C142 VTAIL.n37 B 0.504243f
C143 VTAIL.t10 B 0.083328f
C144 VTAIL.t11 B 0.083328f
C145 VTAIL.n38 B 0.548667f
C146 VTAIL.n39 B 0.761749f
C147 VTAIL.n40 B 0.045806f
C148 VTAIL.n41 B 0.031383f
C149 VTAIL.n42 B 0.016864f
C150 VTAIL.n43 B 0.029895f
C151 VTAIL.n44 B 0.027909f
C152 VTAIL.t6 B 0.069624f
C153 VTAIL.n45 B 0.126174f
C154 VTAIL.n46 B 0.369689f
C155 VTAIL.n47 B 0.016864f
C156 VTAIL.n48 B 0.017856f
C157 VTAIL.n49 B 0.03986f
C158 VTAIL.n50 B 0.089286f
C159 VTAIL.n51 B 0.017856f
C160 VTAIL.n52 B 0.016864f
C161 VTAIL.n53 B 0.067396f
C162 VTAIL.n54 B 0.050103f
C163 VTAIL.n55 B 1.32022f
C164 VTAIL.n56 B 0.045806f
C165 VTAIL.n57 B 0.031383f
C166 VTAIL.n58 B 0.016864f
C167 VTAIL.n59 B 0.029895f
C168 VTAIL.n60 B 0.027909f
C169 VTAIL.t5 B 0.069624f
C170 VTAIL.n61 B 0.126174f
C171 VTAIL.n62 B 0.369689f
C172 VTAIL.n63 B 0.016864f
C173 VTAIL.n64 B 0.017856f
C174 VTAIL.n65 B 0.03986f
C175 VTAIL.n66 B 0.089286f
C176 VTAIL.n67 B 0.017856f
C177 VTAIL.n68 B 0.016864f
C178 VTAIL.n69 B 0.067396f
C179 VTAIL.n70 B 0.050103f
C180 VTAIL.n71 B 1.2422f
C181 VDD1.n0 B 0.03349f
C182 VDD1.n1 B 0.022945f
C183 VDD1.n2 B 0.01233f
C184 VDD1.n3 B 0.021857f
C185 VDD1.n4 B 0.020405f
C186 VDD1.t4 B 0.050904f
C187 VDD1.n5 B 0.092249f
C188 VDD1.n6 B 0.270289f
C189 VDD1.n7 B 0.01233f
C190 VDD1.n8 B 0.013055f
C191 VDD1.n9 B 0.029143f
C192 VDD1.n10 B 0.06528f
C193 VDD1.n11 B 0.013055f
C194 VDD1.n12 B 0.01233f
C195 VDD1.n13 B 0.049275f
C196 VDD1.n14 B 0.061735f
C197 VDD1.n15 B 0.03349f
C198 VDD1.n16 B 0.022945f
C199 VDD1.n17 B 0.01233f
C200 VDD1.n18 B 0.021857f
C201 VDD1.n19 B 0.020405f
C202 VDD1.t1 B 0.050904f
C203 VDD1.n20 B 0.092249f
C204 VDD1.n21 B 0.270289f
C205 VDD1.n22 B 0.01233f
C206 VDD1.n23 B 0.013055f
C207 VDD1.n24 B 0.029143f
C208 VDD1.n25 B 0.06528f
C209 VDD1.n26 B 0.013055f
C210 VDD1.n27 B 0.01233f
C211 VDD1.n28 B 0.049275f
C212 VDD1.n29 B 0.06093f
C213 VDD1.t2 B 0.060923f
C214 VDD1.t3 B 0.060923f
C215 VDD1.n30 B 0.455705f
C216 VDD1.n31 B 2.24123f
C217 VDD1.t5 B 0.060923f
C218 VDD1.t0 B 0.060923f
C219 VDD1.n32 B 0.45182f
C220 VDD1.n33 B 2.04072f
C221 VP.n0 B 0.037713f
C222 VP.t4 B 0.723093f
C223 VP.n1 B 0.057125f
C224 VP.n2 B 0.028607f
C225 VP.n3 B 0.039955f
C226 VP.n4 B 0.028607f
C227 VP.n5 B 0.026575f
C228 VP.n6 B 0.028607f
C229 VP.t3 B 0.723093f
C230 VP.n7 B 0.392274f
C231 VP.n8 B 0.037713f
C232 VP.t5 B 0.723093f
C233 VP.n9 B 0.057125f
C234 VP.n10 B 0.028607f
C235 VP.n11 B 0.039955f
C236 VP.t1 B 0.992709f
C237 VP.t0 B 0.723093f
C238 VP.n12 B 0.38373f
C239 VP.n13 B 0.371627f
C240 VP.n14 B 0.305864f
C241 VP.n15 B 0.028607f
C242 VP.n16 B 0.053049f
C243 VP.n17 B 0.052519f
C244 VP.n18 B 0.026575f
C245 VP.n19 B 0.028607f
C246 VP.n20 B 0.028607f
C247 VP.n21 B 0.028607f
C248 VP.n22 B 0.053049f
C249 VP.n23 B 0.030003f
C250 VP.n24 B 0.392274f
C251 VP.n25 B 1.30277f
C252 VP.n26 B 1.32641f
C253 VP.n27 B 0.037713f
C254 VP.n28 B 0.030003f
C255 VP.n29 B 0.053049f
C256 VP.n30 B 0.057125f
C257 VP.n31 B 0.028607f
C258 VP.n32 B 0.028607f
C259 VP.n33 B 0.028607f
C260 VP.n34 B 0.052519f
C261 VP.n35 B 0.053049f
C262 VP.t2 B 0.723093f
C263 VP.n36 B 0.293765f
C264 VP.n37 B 0.039955f
C265 VP.n38 B 0.028607f
C266 VP.n39 B 0.028607f
C267 VP.n40 B 0.028607f
C268 VP.n41 B 0.053049f
C269 VP.n42 B 0.052519f
C270 VP.n43 B 0.026575f
C271 VP.n44 B 0.028607f
C272 VP.n45 B 0.028607f
C273 VP.n46 B 0.028607f
C274 VP.n47 B 0.053049f
C275 VP.n48 B 0.030003f
C276 VP.n49 B 0.392274f
C277 VP.n50 B 0.055344f
.ends

