* NGSPICE file created from diff_pair_sample_0174.ext - technology: sky130A

.subckt diff_pair_sample_0174 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=7.7298 pd=40.42 as=0 ps=0 w=19.82 l=0.84
X1 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=7.7298 pd=40.42 as=0 ps=0 w=19.82 l=0.84
X2 VDD2.t3 VN.t0 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=3.2703 pd=20.15 as=7.7298 ps=40.42 w=19.82 l=0.84
X3 VTAIL.t0 VP.t0 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=7.7298 pd=40.42 as=3.2703 ps=20.15 w=19.82 l=0.84
X4 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.7298 pd=40.42 as=0 ps=0 w=19.82 l=0.84
X5 VTAIL.t6 VN.t1 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=7.7298 pd=40.42 as=3.2703 ps=20.15 w=19.82 l=0.84
X6 VDD2.t1 VN.t2 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=3.2703 pd=20.15 as=7.7298 ps=40.42 w=19.82 l=0.84
X7 VDD1.t2 VP.t1 VTAIL.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=3.2703 pd=20.15 as=7.7298 ps=40.42 w=19.82 l=0.84
X8 VTAIL.t2 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.7298 pd=40.42 as=3.2703 ps=20.15 w=19.82 l=0.84
X9 VDD1.t0 VP.t3 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=3.2703 pd=20.15 as=7.7298 ps=40.42 w=19.82 l=0.84
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.7298 pd=40.42 as=0 ps=0 w=19.82 l=0.84
X11 VTAIL.t7 VN.t3 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=7.7298 pd=40.42 as=3.2703 ps=20.15 w=19.82 l=0.84
R0 B.n71 B.t8 770.347
R1 B.n77 B.t15 770.347
R2 B.n187 B.t4 770.347
R3 B.n179 B.t12 770.347
R4 B.n579 B.n112 585
R5 B.n112 B.n37 585
R6 B.n581 B.n580 585
R7 B.n583 B.n111 585
R8 B.n586 B.n585 585
R9 B.n587 B.n110 585
R10 B.n589 B.n588 585
R11 B.n591 B.n109 585
R12 B.n594 B.n593 585
R13 B.n595 B.n108 585
R14 B.n597 B.n596 585
R15 B.n599 B.n107 585
R16 B.n602 B.n601 585
R17 B.n603 B.n106 585
R18 B.n605 B.n604 585
R19 B.n607 B.n105 585
R20 B.n610 B.n609 585
R21 B.n611 B.n104 585
R22 B.n613 B.n612 585
R23 B.n615 B.n103 585
R24 B.n618 B.n617 585
R25 B.n619 B.n102 585
R26 B.n621 B.n620 585
R27 B.n623 B.n101 585
R28 B.n626 B.n625 585
R29 B.n627 B.n100 585
R30 B.n629 B.n628 585
R31 B.n631 B.n99 585
R32 B.n634 B.n633 585
R33 B.n635 B.n98 585
R34 B.n637 B.n636 585
R35 B.n639 B.n97 585
R36 B.n642 B.n641 585
R37 B.n643 B.n96 585
R38 B.n645 B.n644 585
R39 B.n647 B.n95 585
R40 B.n650 B.n649 585
R41 B.n651 B.n94 585
R42 B.n653 B.n652 585
R43 B.n655 B.n93 585
R44 B.n658 B.n657 585
R45 B.n659 B.n92 585
R46 B.n661 B.n660 585
R47 B.n663 B.n91 585
R48 B.n666 B.n665 585
R49 B.n667 B.n90 585
R50 B.n669 B.n668 585
R51 B.n671 B.n89 585
R52 B.n674 B.n673 585
R53 B.n675 B.n88 585
R54 B.n677 B.n676 585
R55 B.n679 B.n87 585
R56 B.n682 B.n681 585
R57 B.n683 B.n86 585
R58 B.n685 B.n684 585
R59 B.n687 B.n85 585
R60 B.n690 B.n689 585
R61 B.n691 B.n84 585
R62 B.n693 B.n692 585
R63 B.n695 B.n83 585
R64 B.n698 B.n697 585
R65 B.n699 B.n82 585
R66 B.n701 B.n700 585
R67 B.n703 B.n81 585
R68 B.n705 B.n704 585
R69 B.n707 B.n706 585
R70 B.n710 B.n709 585
R71 B.n711 B.n76 585
R72 B.n713 B.n712 585
R73 B.n715 B.n75 585
R74 B.n718 B.n717 585
R75 B.n719 B.n74 585
R76 B.n721 B.n720 585
R77 B.n723 B.n73 585
R78 B.n726 B.n725 585
R79 B.n728 B.n70 585
R80 B.n730 B.n729 585
R81 B.n732 B.n69 585
R82 B.n735 B.n734 585
R83 B.n736 B.n68 585
R84 B.n738 B.n737 585
R85 B.n740 B.n67 585
R86 B.n743 B.n742 585
R87 B.n744 B.n66 585
R88 B.n746 B.n745 585
R89 B.n748 B.n65 585
R90 B.n751 B.n750 585
R91 B.n752 B.n64 585
R92 B.n754 B.n753 585
R93 B.n756 B.n63 585
R94 B.n759 B.n758 585
R95 B.n760 B.n62 585
R96 B.n762 B.n761 585
R97 B.n764 B.n61 585
R98 B.n767 B.n766 585
R99 B.n768 B.n60 585
R100 B.n770 B.n769 585
R101 B.n772 B.n59 585
R102 B.n775 B.n774 585
R103 B.n776 B.n58 585
R104 B.n778 B.n777 585
R105 B.n780 B.n57 585
R106 B.n783 B.n782 585
R107 B.n784 B.n56 585
R108 B.n786 B.n785 585
R109 B.n788 B.n55 585
R110 B.n791 B.n790 585
R111 B.n792 B.n54 585
R112 B.n794 B.n793 585
R113 B.n796 B.n53 585
R114 B.n799 B.n798 585
R115 B.n800 B.n52 585
R116 B.n802 B.n801 585
R117 B.n804 B.n51 585
R118 B.n807 B.n806 585
R119 B.n808 B.n50 585
R120 B.n810 B.n809 585
R121 B.n812 B.n49 585
R122 B.n815 B.n814 585
R123 B.n816 B.n48 585
R124 B.n818 B.n817 585
R125 B.n820 B.n47 585
R126 B.n823 B.n822 585
R127 B.n824 B.n46 585
R128 B.n826 B.n825 585
R129 B.n828 B.n45 585
R130 B.n831 B.n830 585
R131 B.n832 B.n44 585
R132 B.n834 B.n833 585
R133 B.n836 B.n43 585
R134 B.n839 B.n838 585
R135 B.n840 B.n42 585
R136 B.n842 B.n841 585
R137 B.n844 B.n41 585
R138 B.n847 B.n846 585
R139 B.n848 B.n40 585
R140 B.n850 B.n849 585
R141 B.n852 B.n39 585
R142 B.n855 B.n854 585
R143 B.n856 B.n38 585
R144 B.n578 B.n36 585
R145 B.n859 B.n36 585
R146 B.n577 B.n35 585
R147 B.n860 B.n35 585
R148 B.n576 B.n34 585
R149 B.n861 B.n34 585
R150 B.n575 B.n574 585
R151 B.n574 B.n30 585
R152 B.n573 B.n29 585
R153 B.n867 B.n29 585
R154 B.n572 B.n28 585
R155 B.n868 B.n28 585
R156 B.n571 B.n27 585
R157 B.n869 B.n27 585
R158 B.n570 B.n569 585
R159 B.n569 B.n23 585
R160 B.n568 B.n22 585
R161 B.n875 B.n22 585
R162 B.n567 B.n21 585
R163 B.n876 B.n21 585
R164 B.n566 B.n20 585
R165 B.n877 B.n20 585
R166 B.n565 B.n564 585
R167 B.n564 B.n19 585
R168 B.n563 B.n15 585
R169 B.n883 B.n15 585
R170 B.n562 B.n14 585
R171 B.n884 B.n14 585
R172 B.n561 B.n13 585
R173 B.n885 B.n13 585
R174 B.n560 B.n559 585
R175 B.n559 B.n12 585
R176 B.n558 B.n557 585
R177 B.n558 B.n8 585
R178 B.n556 B.n7 585
R179 B.n892 B.n7 585
R180 B.n555 B.n6 585
R181 B.n893 B.n6 585
R182 B.n554 B.n5 585
R183 B.n894 B.n5 585
R184 B.n553 B.n552 585
R185 B.n552 B.n4 585
R186 B.n551 B.n113 585
R187 B.n551 B.n550 585
R188 B.n540 B.n114 585
R189 B.n543 B.n114 585
R190 B.n542 B.n541 585
R191 B.n544 B.n542 585
R192 B.n539 B.n119 585
R193 B.n119 B.n118 585
R194 B.n538 B.n537 585
R195 B.n537 B.n536 585
R196 B.n121 B.n120 585
R197 B.n529 B.n121 585
R198 B.n528 B.n527 585
R199 B.n530 B.n528 585
R200 B.n526 B.n126 585
R201 B.n126 B.n125 585
R202 B.n525 B.n524 585
R203 B.n524 B.n523 585
R204 B.n128 B.n127 585
R205 B.n129 B.n128 585
R206 B.n516 B.n515 585
R207 B.n517 B.n516 585
R208 B.n514 B.n133 585
R209 B.n137 B.n133 585
R210 B.n513 B.n512 585
R211 B.n512 B.n511 585
R212 B.n135 B.n134 585
R213 B.n136 B.n135 585
R214 B.n504 B.n503 585
R215 B.n505 B.n504 585
R216 B.n502 B.n142 585
R217 B.n142 B.n141 585
R218 B.n501 B.n500 585
R219 B.n500 B.n499 585
R220 B.n496 B.n146 585
R221 B.n495 B.n494 585
R222 B.n492 B.n147 585
R223 B.n492 B.n145 585
R224 B.n491 B.n490 585
R225 B.n489 B.n488 585
R226 B.n487 B.n149 585
R227 B.n485 B.n484 585
R228 B.n483 B.n150 585
R229 B.n482 B.n481 585
R230 B.n479 B.n151 585
R231 B.n477 B.n476 585
R232 B.n475 B.n152 585
R233 B.n474 B.n473 585
R234 B.n471 B.n153 585
R235 B.n469 B.n468 585
R236 B.n467 B.n154 585
R237 B.n466 B.n465 585
R238 B.n463 B.n155 585
R239 B.n461 B.n460 585
R240 B.n459 B.n156 585
R241 B.n458 B.n457 585
R242 B.n455 B.n157 585
R243 B.n453 B.n452 585
R244 B.n451 B.n158 585
R245 B.n450 B.n449 585
R246 B.n447 B.n159 585
R247 B.n445 B.n444 585
R248 B.n443 B.n160 585
R249 B.n442 B.n441 585
R250 B.n439 B.n161 585
R251 B.n437 B.n436 585
R252 B.n435 B.n162 585
R253 B.n434 B.n433 585
R254 B.n431 B.n163 585
R255 B.n429 B.n428 585
R256 B.n427 B.n164 585
R257 B.n426 B.n425 585
R258 B.n423 B.n165 585
R259 B.n421 B.n420 585
R260 B.n419 B.n166 585
R261 B.n418 B.n417 585
R262 B.n415 B.n167 585
R263 B.n413 B.n412 585
R264 B.n411 B.n168 585
R265 B.n410 B.n409 585
R266 B.n407 B.n169 585
R267 B.n405 B.n404 585
R268 B.n403 B.n170 585
R269 B.n402 B.n401 585
R270 B.n399 B.n171 585
R271 B.n397 B.n396 585
R272 B.n395 B.n172 585
R273 B.n394 B.n393 585
R274 B.n391 B.n173 585
R275 B.n389 B.n388 585
R276 B.n387 B.n174 585
R277 B.n386 B.n385 585
R278 B.n383 B.n175 585
R279 B.n381 B.n380 585
R280 B.n379 B.n176 585
R281 B.n378 B.n377 585
R282 B.n375 B.n177 585
R283 B.n373 B.n372 585
R284 B.n371 B.n178 585
R285 B.n370 B.n369 585
R286 B.n367 B.n366 585
R287 B.n365 B.n364 585
R288 B.n363 B.n183 585
R289 B.n361 B.n360 585
R290 B.n359 B.n184 585
R291 B.n358 B.n357 585
R292 B.n355 B.n185 585
R293 B.n353 B.n352 585
R294 B.n351 B.n186 585
R295 B.n349 B.n348 585
R296 B.n346 B.n189 585
R297 B.n344 B.n343 585
R298 B.n342 B.n190 585
R299 B.n341 B.n340 585
R300 B.n338 B.n191 585
R301 B.n336 B.n335 585
R302 B.n334 B.n192 585
R303 B.n333 B.n332 585
R304 B.n330 B.n193 585
R305 B.n328 B.n327 585
R306 B.n326 B.n194 585
R307 B.n325 B.n324 585
R308 B.n322 B.n195 585
R309 B.n320 B.n319 585
R310 B.n318 B.n196 585
R311 B.n317 B.n316 585
R312 B.n314 B.n197 585
R313 B.n312 B.n311 585
R314 B.n310 B.n198 585
R315 B.n309 B.n308 585
R316 B.n306 B.n199 585
R317 B.n304 B.n303 585
R318 B.n302 B.n200 585
R319 B.n301 B.n300 585
R320 B.n298 B.n201 585
R321 B.n296 B.n295 585
R322 B.n294 B.n202 585
R323 B.n293 B.n292 585
R324 B.n290 B.n203 585
R325 B.n288 B.n287 585
R326 B.n286 B.n204 585
R327 B.n285 B.n284 585
R328 B.n282 B.n205 585
R329 B.n280 B.n279 585
R330 B.n278 B.n206 585
R331 B.n277 B.n276 585
R332 B.n274 B.n207 585
R333 B.n272 B.n271 585
R334 B.n270 B.n208 585
R335 B.n269 B.n268 585
R336 B.n266 B.n209 585
R337 B.n264 B.n263 585
R338 B.n262 B.n210 585
R339 B.n261 B.n260 585
R340 B.n258 B.n211 585
R341 B.n256 B.n255 585
R342 B.n254 B.n212 585
R343 B.n253 B.n252 585
R344 B.n250 B.n213 585
R345 B.n248 B.n247 585
R346 B.n246 B.n214 585
R347 B.n245 B.n244 585
R348 B.n242 B.n215 585
R349 B.n240 B.n239 585
R350 B.n238 B.n216 585
R351 B.n237 B.n236 585
R352 B.n234 B.n217 585
R353 B.n232 B.n231 585
R354 B.n230 B.n218 585
R355 B.n229 B.n228 585
R356 B.n226 B.n219 585
R357 B.n224 B.n223 585
R358 B.n222 B.n221 585
R359 B.n144 B.n143 585
R360 B.n498 B.n497 585
R361 B.n499 B.n498 585
R362 B.n140 B.n139 585
R363 B.n141 B.n140 585
R364 B.n507 B.n506 585
R365 B.n506 B.n505 585
R366 B.n508 B.n138 585
R367 B.n138 B.n136 585
R368 B.n510 B.n509 585
R369 B.n511 B.n510 585
R370 B.n132 B.n131 585
R371 B.n137 B.n132 585
R372 B.n519 B.n518 585
R373 B.n518 B.n517 585
R374 B.n520 B.n130 585
R375 B.n130 B.n129 585
R376 B.n522 B.n521 585
R377 B.n523 B.n522 585
R378 B.n124 B.n123 585
R379 B.n125 B.n124 585
R380 B.n532 B.n531 585
R381 B.n531 B.n530 585
R382 B.n533 B.n122 585
R383 B.n529 B.n122 585
R384 B.n535 B.n534 585
R385 B.n536 B.n535 585
R386 B.n117 B.n116 585
R387 B.n118 B.n117 585
R388 B.n546 B.n545 585
R389 B.n545 B.n544 585
R390 B.n547 B.n115 585
R391 B.n543 B.n115 585
R392 B.n549 B.n548 585
R393 B.n550 B.n549 585
R394 B.n3 B.n0 585
R395 B.n4 B.n3 585
R396 B.n891 B.n1 585
R397 B.n892 B.n891 585
R398 B.n890 B.n889 585
R399 B.n890 B.n8 585
R400 B.n888 B.n9 585
R401 B.n12 B.n9 585
R402 B.n887 B.n886 585
R403 B.n886 B.n885 585
R404 B.n11 B.n10 585
R405 B.n884 B.n11 585
R406 B.n882 B.n881 585
R407 B.n883 B.n882 585
R408 B.n880 B.n16 585
R409 B.n19 B.n16 585
R410 B.n879 B.n878 585
R411 B.n878 B.n877 585
R412 B.n18 B.n17 585
R413 B.n876 B.n18 585
R414 B.n874 B.n873 585
R415 B.n875 B.n874 585
R416 B.n872 B.n24 585
R417 B.n24 B.n23 585
R418 B.n871 B.n870 585
R419 B.n870 B.n869 585
R420 B.n26 B.n25 585
R421 B.n868 B.n26 585
R422 B.n866 B.n865 585
R423 B.n867 B.n866 585
R424 B.n864 B.n31 585
R425 B.n31 B.n30 585
R426 B.n863 B.n862 585
R427 B.n862 B.n861 585
R428 B.n33 B.n32 585
R429 B.n860 B.n33 585
R430 B.n858 B.n857 585
R431 B.n859 B.n858 585
R432 B.n895 B.n894 585
R433 B.n893 B.n2 585
R434 B.n858 B.n38 473.281
R435 B.n112 B.n36 473.281
R436 B.n500 B.n144 473.281
R437 B.n498 B.n146 473.281
R438 B.n582 B.n37 256.663
R439 B.n584 B.n37 256.663
R440 B.n590 B.n37 256.663
R441 B.n592 B.n37 256.663
R442 B.n598 B.n37 256.663
R443 B.n600 B.n37 256.663
R444 B.n606 B.n37 256.663
R445 B.n608 B.n37 256.663
R446 B.n614 B.n37 256.663
R447 B.n616 B.n37 256.663
R448 B.n622 B.n37 256.663
R449 B.n624 B.n37 256.663
R450 B.n630 B.n37 256.663
R451 B.n632 B.n37 256.663
R452 B.n638 B.n37 256.663
R453 B.n640 B.n37 256.663
R454 B.n646 B.n37 256.663
R455 B.n648 B.n37 256.663
R456 B.n654 B.n37 256.663
R457 B.n656 B.n37 256.663
R458 B.n662 B.n37 256.663
R459 B.n664 B.n37 256.663
R460 B.n670 B.n37 256.663
R461 B.n672 B.n37 256.663
R462 B.n678 B.n37 256.663
R463 B.n680 B.n37 256.663
R464 B.n686 B.n37 256.663
R465 B.n688 B.n37 256.663
R466 B.n694 B.n37 256.663
R467 B.n696 B.n37 256.663
R468 B.n702 B.n37 256.663
R469 B.n80 B.n37 256.663
R470 B.n708 B.n37 256.663
R471 B.n714 B.n37 256.663
R472 B.n716 B.n37 256.663
R473 B.n722 B.n37 256.663
R474 B.n724 B.n37 256.663
R475 B.n731 B.n37 256.663
R476 B.n733 B.n37 256.663
R477 B.n739 B.n37 256.663
R478 B.n741 B.n37 256.663
R479 B.n747 B.n37 256.663
R480 B.n749 B.n37 256.663
R481 B.n755 B.n37 256.663
R482 B.n757 B.n37 256.663
R483 B.n763 B.n37 256.663
R484 B.n765 B.n37 256.663
R485 B.n771 B.n37 256.663
R486 B.n773 B.n37 256.663
R487 B.n779 B.n37 256.663
R488 B.n781 B.n37 256.663
R489 B.n787 B.n37 256.663
R490 B.n789 B.n37 256.663
R491 B.n795 B.n37 256.663
R492 B.n797 B.n37 256.663
R493 B.n803 B.n37 256.663
R494 B.n805 B.n37 256.663
R495 B.n811 B.n37 256.663
R496 B.n813 B.n37 256.663
R497 B.n819 B.n37 256.663
R498 B.n821 B.n37 256.663
R499 B.n827 B.n37 256.663
R500 B.n829 B.n37 256.663
R501 B.n835 B.n37 256.663
R502 B.n837 B.n37 256.663
R503 B.n843 B.n37 256.663
R504 B.n845 B.n37 256.663
R505 B.n851 B.n37 256.663
R506 B.n853 B.n37 256.663
R507 B.n493 B.n145 256.663
R508 B.n148 B.n145 256.663
R509 B.n486 B.n145 256.663
R510 B.n480 B.n145 256.663
R511 B.n478 B.n145 256.663
R512 B.n472 B.n145 256.663
R513 B.n470 B.n145 256.663
R514 B.n464 B.n145 256.663
R515 B.n462 B.n145 256.663
R516 B.n456 B.n145 256.663
R517 B.n454 B.n145 256.663
R518 B.n448 B.n145 256.663
R519 B.n446 B.n145 256.663
R520 B.n440 B.n145 256.663
R521 B.n438 B.n145 256.663
R522 B.n432 B.n145 256.663
R523 B.n430 B.n145 256.663
R524 B.n424 B.n145 256.663
R525 B.n422 B.n145 256.663
R526 B.n416 B.n145 256.663
R527 B.n414 B.n145 256.663
R528 B.n408 B.n145 256.663
R529 B.n406 B.n145 256.663
R530 B.n400 B.n145 256.663
R531 B.n398 B.n145 256.663
R532 B.n392 B.n145 256.663
R533 B.n390 B.n145 256.663
R534 B.n384 B.n145 256.663
R535 B.n382 B.n145 256.663
R536 B.n376 B.n145 256.663
R537 B.n374 B.n145 256.663
R538 B.n368 B.n145 256.663
R539 B.n182 B.n145 256.663
R540 B.n362 B.n145 256.663
R541 B.n356 B.n145 256.663
R542 B.n354 B.n145 256.663
R543 B.n347 B.n145 256.663
R544 B.n345 B.n145 256.663
R545 B.n339 B.n145 256.663
R546 B.n337 B.n145 256.663
R547 B.n331 B.n145 256.663
R548 B.n329 B.n145 256.663
R549 B.n323 B.n145 256.663
R550 B.n321 B.n145 256.663
R551 B.n315 B.n145 256.663
R552 B.n313 B.n145 256.663
R553 B.n307 B.n145 256.663
R554 B.n305 B.n145 256.663
R555 B.n299 B.n145 256.663
R556 B.n297 B.n145 256.663
R557 B.n291 B.n145 256.663
R558 B.n289 B.n145 256.663
R559 B.n283 B.n145 256.663
R560 B.n281 B.n145 256.663
R561 B.n275 B.n145 256.663
R562 B.n273 B.n145 256.663
R563 B.n267 B.n145 256.663
R564 B.n265 B.n145 256.663
R565 B.n259 B.n145 256.663
R566 B.n257 B.n145 256.663
R567 B.n251 B.n145 256.663
R568 B.n249 B.n145 256.663
R569 B.n243 B.n145 256.663
R570 B.n241 B.n145 256.663
R571 B.n235 B.n145 256.663
R572 B.n233 B.n145 256.663
R573 B.n227 B.n145 256.663
R574 B.n225 B.n145 256.663
R575 B.n220 B.n145 256.663
R576 B.n897 B.n896 256.663
R577 B.n854 B.n852 163.367
R578 B.n850 B.n40 163.367
R579 B.n846 B.n844 163.367
R580 B.n842 B.n42 163.367
R581 B.n838 B.n836 163.367
R582 B.n834 B.n44 163.367
R583 B.n830 B.n828 163.367
R584 B.n826 B.n46 163.367
R585 B.n822 B.n820 163.367
R586 B.n818 B.n48 163.367
R587 B.n814 B.n812 163.367
R588 B.n810 B.n50 163.367
R589 B.n806 B.n804 163.367
R590 B.n802 B.n52 163.367
R591 B.n798 B.n796 163.367
R592 B.n794 B.n54 163.367
R593 B.n790 B.n788 163.367
R594 B.n786 B.n56 163.367
R595 B.n782 B.n780 163.367
R596 B.n778 B.n58 163.367
R597 B.n774 B.n772 163.367
R598 B.n770 B.n60 163.367
R599 B.n766 B.n764 163.367
R600 B.n762 B.n62 163.367
R601 B.n758 B.n756 163.367
R602 B.n754 B.n64 163.367
R603 B.n750 B.n748 163.367
R604 B.n746 B.n66 163.367
R605 B.n742 B.n740 163.367
R606 B.n738 B.n68 163.367
R607 B.n734 B.n732 163.367
R608 B.n730 B.n70 163.367
R609 B.n725 B.n723 163.367
R610 B.n721 B.n74 163.367
R611 B.n717 B.n715 163.367
R612 B.n713 B.n76 163.367
R613 B.n709 B.n707 163.367
R614 B.n704 B.n703 163.367
R615 B.n701 B.n82 163.367
R616 B.n697 B.n695 163.367
R617 B.n693 B.n84 163.367
R618 B.n689 B.n687 163.367
R619 B.n685 B.n86 163.367
R620 B.n681 B.n679 163.367
R621 B.n677 B.n88 163.367
R622 B.n673 B.n671 163.367
R623 B.n669 B.n90 163.367
R624 B.n665 B.n663 163.367
R625 B.n661 B.n92 163.367
R626 B.n657 B.n655 163.367
R627 B.n653 B.n94 163.367
R628 B.n649 B.n647 163.367
R629 B.n645 B.n96 163.367
R630 B.n641 B.n639 163.367
R631 B.n637 B.n98 163.367
R632 B.n633 B.n631 163.367
R633 B.n629 B.n100 163.367
R634 B.n625 B.n623 163.367
R635 B.n621 B.n102 163.367
R636 B.n617 B.n615 163.367
R637 B.n613 B.n104 163.367
R638 B.n609 B.n607 163.367
R639 B.n605 B.n106 163.367
R640 B.n601 B.n599 163.367
R641 B.n597 B.n108 163.367
R642 B.n593 B.n591 163.367
R643 B.n589 B.n110 163.367
R644 B.n585 B.n583 163.367
R645 B.n581 B.n112 163.367
R646 B.n500 B.n142 163.367
R647 B.n504 B.n142 163.367
R648 B.n504 B.n135 163.367
R649 B.n512 B.n135 163.367
R650 B.n512 B.n133 163.367
R651 B.n516 B.n133 163.367
R652 B.n516 B.n128 163.367
R653 B.n524 B.n128 163.367
R654 B.n524 B.n126 163.367
R655 B.n528 B.n126 163.367
R656 B.n528 B.n121 163.367
R657 B.n537 B.n121 163.367
R658 B.n537 B.n119 163.367
R659 B.n542 B.n119 163.367
R660 B.n542 B.n114 163.367
R661 B.n551 B.n114 163.367
R662 B.n552 B.n551 163.367
R663 B.n552 B.n5 163.367
R664 B.n6 B.n5 163.367
R665 B.n7 B.n6 163.367
R666 B.n558 B.n7 163.367
R667 B.n559 B.n558 163.367
R668 B.n559 B.n13 163.367
R669 B.n14 B.n13 163.367
R670 B.n15 B.n14 163.367
R671 B.n564 B.n15 163.367
R672 B.n564 B.n20 163.367
R673 B.n21 B.n20 163.367
R674 B.n22 B.n21 163.367
R675 B.n569 B.n22 163.367
R676 B.n569 B.n27 163.367
R677 B.n28 B.n27 163.367
R678 B.n29 B.n28 163.367
R679 B.n574 B.n29 163.367
R680 B.n574 B.n34 163.367
R681 B.n35 B.n34 163.367
R682 B.n36 B.n35 163.367
R683 B.n494 B.n492 163.367
R684 B.n492 B.n491 163.367
R685 B.n488 B.n487 163.367
R686 B.n485 B.n150 163.367
R687 B.n481 B.n479 163.367
R688 B.n477 B.n152 163.367
R689 B.n473 B.n471 163.367
R690 B.n469 B.n154 163.367
R691 B.n465 B.n463 163.367
R692 B.n461 B.n156 163.367
R693 B.n457 B.n455 163.367
R694 B.n453 B.n158 163.367
R695 B.n449 B.n447 163.367
R696 B.n445 B.n160 163.367
R697 B.n441 B.n439 163.367
R698 B.n437 B.n162 163.367
R699 B.n433 B.n431 163.367
R700 B.n429 B.n164 163.367
R701 B.n425 B.n423 163.367
R702 B.n421 B.n166 163.367
R703 B.n417 B.n415 163.367
R704 B.n413 B.n168 163.367
R705 B.n409 B.n407 163.367
R706 B.n405 B.n170 163.367
R707 B.n401 B.n399 163.367
R708 B.n397 B.n172 163.367
R709 B.n393 B.n391 163.367
R710 B.n389 B.n174 163.367
R711 B.n385 B.n383 163.367
R712 B.n381 B.n176 163.367
R713 B.n377 B.n375 163.367
R714 B.n373 B.n178 163.367
R715 B.n369 B.n367 163.367
R716 B.n364 B.n363 163.367
R717 B.n361 B.n184 163.367
R718 B.n357 B.n355 163.367
R719 B.n353 B.n186 163.367
R720 B.n348 B.n346 163.367
R721 B.n344 B.n190 163.367
R722 B.n340 B.n338 163.367
R723 B.n336 B.n192 163.367
R724 B.n332 B.n330 163.367
R725 B.n328 B.n194 163.367
R726 B.n324 B.n322 163.367
R727 B.n320 B.n196 163.367
R728 B.n316 B.n314 163.367
R729 B.n312 B.n198 163.367
R730 B.n308 B.n306 163.367
R731 B.n304 B.n200 163.367
R732 B.n300 B.n298 163.367
R733 B.n296 B.n202 163.367
R734 B.n292 B.n290 163.367
R735 B.n288 B.n204 163.367
R736 B.n284 B.n282 163.367
R737 B.n280 B.n206 163.367
R738 B.n276 B.n274 163.367
R739 B.n272 B.n208 163.367
R740 B.n268 B.n266 163.367
R741 B.n264 B.n210 163.367
R742 B.n260 B.n258 163.367
R743 B.n256 B.n212 163.367
R744 B.n252 B.n250 163.367
R745 B.n248 B.n214 163.367
R746 B.n244 B.n242 163.367
R747 B.n240 B.n216 163.367
R748 B.n236 B.n234 163.367
R749 B.n232 B.n218 163.367
R750 B.n228 B.n226 163.367
R751 B.n224 B.n221 163.367
R752 B.n498 B.n140 163.367
R753 B.n506 B.n140 163.367
R754 B.n506 B.n138 163.367
R755 B.n510 B.n138 163.367
R756 B.n510 B.n132 163.367
R757 B.n518 B.n132 163.367
R758 B.n518 B.n130 163.367
R759 B.n522 B.n130 163.367
R760 B.n522 B.n124 163.367
R761 B.n531 B.n124 163.367
R762 B.n531 B.n122 163.367
R763 B.n535 B.n122 163.367
R764 B.n535 B.n117 163.367
R765 B.n545 B.n117 163.367
R766 B.n545 B.n115 163.367
R767 B.n549 B.n115 163.367
R768 B.n549 B.n3 163.367
R769 B.n895 B.n3 163.367
R770 B.n891 B.n2 163.367
R771 B.n891 B.n890 163.367
R772 B.n890 B.n9 163.367
R773 B.n886 B.n9 163.367
R774 B.n886 B.n11 163.367
R775 B.n882 B.n11 163.367
R776 B.n882 B.n16 163.367
R777 B.n878 B.n16 163.367
R778 B.n878 B.n18 163.367
R779 B.n874 B.n18 163.367
R780 B.n874 B.n24 163.367
R781 B.n870 B.n24 163.367
R782 B.n870 B.n26 163.367
R783 B.n866 B.n26 163.367
R784 B.n866 B.n31 163.367
R785 B.n862 B.n31 163.367
R786 B.n862 B.n33 163.367
R787 B.n858 B.n33 163.367
R788 B.n77 B.t16 91.7807
R789 B.n187 B.t7 91.7807
R790 B.n71 B.t10 91.754
R791 B.n179 B.t14 91.754
R792 B.n853 B.n38 71.676
R793 B.n852 B.n851 71.676
R794 B.n845 B.n40 71.676
R795 B.n844 B.n843 71.676
R796 B.n837 B.n42 71.676
R797 B.n836 B.n835 71.676
R798 B.n829 B.n44 71.676
R799 B.n828 B.n827 71.676
R800 B.n821 B.n46 71.676
R801 B.n820 B.n819 71.676
R802 B.n813 B.n48 71.676
R803 B.n812 B.n811 71.676
R804 B.n805 B.n50 71.676
R805 B.n804 B.n803 71.676
R806 B.n797 B.n52 71.676
R807 B.n796 B.n795 71.676
R808 B.n789 B.n54 71.676
R809 B.n788 B.n787 71.676
R810 B.n781 B.n56 71.676
R811 B.n780 B.n779 71.676
R812 B.n773 B.n58 71.676
R813 B.n772 B.n771 71.676
R814 B.n765 B.n60 71.676
R815 B.n764 B.n763 71.676
R816 B.n757 B.n62 71.676
R817 B.n756 B.n755 71.676
R818 B.n749 B.n64 71.676
R819 B.n748 B.n747 71.676
R820 B.n741 B.n66 71.676
R821 B.n740 B.n739 71.676
R822 B.n733 B.n68 71.676
R823 B.n732 B.n731 71.676
R824 B.n724 B.n70 71.676
R825 B.n723 B.n722 71.676
R826 B.n716 B.n74 71.676
R827 B.n715 B.n714 71.676
R828 B.n708 B.n76 71.676
R829 B.n707 B.n80 71.676
R830 B.n703 B.n702 71.676
R831 B.n696 B.n82 71.676
R832 B.n695 B.n694 71.676
R833 B.n688 B.n84 71.676
R834 B.n687 B.n686 71.676
R835 B.n680 B.n86 71.676
R836 B.n679 B.n678 71.676
R837 B.n672 B.n88 71.676
R838 B.n671 B.n670 71.676
R839 B.n664 B.n90 71.676
R840 B.n663 B.n662 71.676
R841 B.n656 B.n92 71.676
R842 B.n655 B.n654 71.676
R843 B.n648 B.n94 71.676
R844 B.n647 B.n646 71.676
R845 B.n640 B.n96 71.676
R846 B.n639 B.n638 71.676
R847 B.n632 B.n98 71.676
R848 B.n631 B.n630 71.676
R849 B.n624 B.n100 71.676
R850 B.n623 B.n622 71.676
R851 B.n616 B.n102 71.676
R852 B.n615 B.n614 71.676
R853 B.n608 B.n104 71.676
R854 B.n607 B.n606 71.676
R855 B.n600 B.n106 71.676
R856 B.n599 B.n598 71.676
R857 B.n592 B.n108 71.676
R858 B.n591 B.n590 71.676
R859 B.n584 B.n110 71.676
R860 B.n583 B.n582 71.676
R861 B.n582 B.n581 71.676
R862 B.n585 B.n584 71.676
R863 B.n590 B.n589 71.676
R864 B.n593 B.n592 71.676
R865 B.n598 B.n597 71.676
R866 B.n601 B.n600 71.676
R867 B.n606 B.n605 71.676
R868 B.n609 B.n608 71.676
R869 B.n614 B.n613 71.676
R870 B.n617 B.n616 71.676
R871 B.n622 B.n621 71.676
R872 B.n625 B.n624 71.676
R873 B.n630 B.n629 71.676
R874 B.n633 B.n632 71.676
R875 B.n638 B.n637 71.676
R876 B.n641 B.n640 71.676
R877 B.n646 B.n645 71.676
R878 B.n649 B.n648 71.676
R879 B.n654 B.n653 71.676
R880 B.n657 B.n656 71.676
R881 B.n662 B.n661 71.676
R882 B.n665 B.n664 71.676
R883 B.n670 B.n669 71.676
R884 B.n673 B.n672 71.676
R885 B.n678 B.n677 71.676
R886 B.n681 B.n680 71.676
R887 B.n686 B.n685 71.676
R888 B.n689 B.n688 71.676
R889 B.n694 B.n693 71.676
R890 B.n697 B.n696 71.676
R891 B.n702 B.n701 71.676
R892 B.n704 B.n80 71.676
R893 B.n709 B.n708 71.676
R894 B.n714 B.n713 71.676
R895 B.n717 B.n716 71.676
R896 B.n722 B.n721 71.676
R897 B.n725 B.n724 71.676
R898 B.n731 B.n730 71.676
R899 B.n734 B.n733 71.676
R900 B.n739 B.n738 71.676
R901 B.n742 B.n741 71.676
R902 B.n747 B.n746 71.676
R903 B.n750 B.n749 71.676
R904 B.n755 B.n754 71.676
R905 B.n758 B.n757 71.676
R906 B.n763 B.n762 71.676
R907 B.n766 B.n765 71.676
R908 B.n771 B.n770 71.676
R909 B.n774 B.n773 71.676
R910 B.n779 B.n778 71.676
R911 B.n782 B.n781 71.676
R912 B.n787 B.n786 71.676
R913 B.n790 B.n789 71.676
R914 B.n795 B.n794 71.676
R915 B.n798 B.n797 71.676
R916 B.n803 B.n802 71.676
R917 B.n806 B.n805 71.676
R918 B.n811 B.n810 71.676
R919 B.n814 B.n813 71.676
R920 B.n819 B.n818 71.676
R921 B.n822 B.n821 71.676
R922 B.n827 B.n826 71.676
R923 B.n830 B.n829 71.676
R924 B.n835 B.n834 71.676
R925 B.n838 B.n837 71.676
R926 B.n843 B.n842 71.676
R927 B.n846 B.n845 71.676
R928 B.n851 B.n850 71.676
R929 B.n854 B.n853 71.676
R930 B.n493 B.n146 71.676
R931 B.n491 B.n148 71.676
R932 B.n487 B.n486 71.676
R933 B.n480 B.n150 71.676
R934 B.n479 B.n478 71.676
R935 B.n472 B.n152 71.676
R936 B.n471 B.n470 71.676
R937 B.n464 B.n154 71.676
R938 B.n463 B.n462 71.676
R939 B.n456 B.n156 71.676
R940 B.n455 B.n454 71.676
R941 B.n448 B.n158 71.676
R942 B.n447 B.n446 71.676
R943 B.n440 B.n160 71.676
R944 B.n439 B.n438 71.676
R945 B.n432 B.n162 71.676
R946 B.n431 B.n430 71.676
R947 B.n424 B.n164 71.676
R948 B.n423 B.n422 71.676
R949 B.n416 B.n166 71.676
R950 B.n415 B.n414 71.676
R951 B.n408 B.n168 71.676
R952 B.n407 B.n406 71.676
R953 B.n400 B.n170 71.676
R954 B.n399 B.n398 71.676
R955 B.n392 B.n172 71.676
R956 B.n391 B.n390 71.676
R957 B.n384 B.n174 71.676
R958 B.n383 B.n382 71.676
R959 B.n376 B.n176 71.676
R960 B.n375 B.n374 71.676
R961 B.n368 B.n178 71.676
R962 B.n367 B.n182 71.676
R963 B.n363 B.n362 71.676
R964 B.n356 B.n184 71.676
R965 B.n355 B.n354 71.676
R966 B.n347 B.n186 71.676
R967 B.n346 B.n345 71.676
R968 B.n339 B.n190 71.676
R969 B.n338 B.n337 71.676
R970 B.n331 B.n192 71.676
R971 B.n330 B.n329 71.676
R972 B.n323 B.n194 71.676
R973 B.n322 B.n321 71.676
R974 B.n315 B.n196 71.676
R975 B.n314 B.n313 71.676
R976 B.n307 B.n198 71.676
R977 B.n306 B.n305 71.676
R978 B.n299 B.n200 71.676
R979 B.n298 B.n297 71.676
R980 B.n291 B.n202 71.676
R981 B.n290 B.n289 71.676
R982 B.n283 B.n204 71.676
R983 B.n282 B.n281 71.676
R984 B.n275 B.n206 71.676
R985 B.n274 B.n273 71.676
R986 B.n267 B.n208 71.676
R987 B.n266 B.n265 71.676
R988 B.n259 B.n210 71.676
R989 B.n258 B.n257 71.676
R990 B.n251 B.n212 71.676
R991 B.n250 B.n249 71.676
R992 B.n243 B.n214 71.676
R993 B.n242 B.n241 71.676
R994 B.n235 B.n216 71.676
R995 B.n234 B.n233 71.676
R996 B.n227 B.n218 71.676
R997 B.n226 B.n225 71.676
R998 B.n221 B.n220 71.676
R999 B.n494 B.n493 71.676
R1000 B.n488 B.n148 71.676
R1001 B.n486 B.n485 71.676
R1002 B.n481 B.n480 71.676
R1003 B.n478 B.n477 71.676
R1004 B.n473 B.n472 71.676
R1005 B.n470 B.n469 71.676
R1006 B.n465 B.n464 71.676
R1007 B.n462 B.n461 71.676
R1008 B.n457 B.n456 71.676
R1009 B.n454 B.n453 71.676
R1010 B.n449 B.n448 71.676
R1011 B.n446 B.n445 71.676
R1012 B.n441 B.n440 71.676
R1013 B.n438 B.n437 71.676
R1014 B.n433 B.n432 71.676
R1015 B.n430 B.n429 71.676
R1016 B.n425 B.n424 71.676
R1017 B.n422 B.n421 71.676
R1018 B.n417 B.n416 71.676
R1019 B.n414 B.n413 71.676
R1020 B.n409 B.n408 71.676
R1021 B.n406 B.n405 71.676
R1022 B.n401 B.n400 71.676
R1023 B.n398 B.n397 71.676
R1024 B.n393 B.n392 71.676
R1025 B.n390 B.n389 71.676
R1026 B.n385 B.n384 71.676
R1027 B.n382 B.n381 71.676
R1028 B.n377 B.n376 71.676
R1029 B.n374 B.n373 71.676
R1030 B.n369 B.n368 71.676
R1031 B.n364 B.n182 71.676
R1032 B.n362 B.n361 71.676
R1033 B.n357 B.n356 71.676
R1034 B.n354 B.n353 71.676
R1035 B.n348 B.n347 71.676
R1036 B.n345 B.n344 71.676
R1037 B.n340 B.n339 71.676
R1038 B.n337 B.n336 71.676
R1039 B.n332 B.n331 71.676
R1040 B.n329 B.n328 71.676
R1041 B.n324 B.n323 71.676
R1042 B.n321 B.n320 71.676
R1043 B.n316 B.n315 71.676
R1044 B.n313 B.n312 71.676
R1045 B.n308 B.n307 71.676
R1046 B.n305 B.n304 71.676
R1047 B.n300 B.n299 71.676
R1048 B.n297 B.n296 71.676
R1049 B.n292 B.n291 71.676
R1050 B.n289 B.n288 71.676
R1051 B.n284 B.n283 71.676
R1052 B.n281 B.n280 71.676
R1053 B.n276 B.n275 71.676
R1054 B.n273 B.n272 71.676
R1055 B.n268 B.n267 71.676
R1056 B.n265 B.n264 71.676
R1057 B.n260 B.n259 71.676
R1058 B.n257 B.n256 71.676
R1059 B.n252 B.n251 71.676
R1060 B.n249 B.n248 71.676
R1061 B.n244 B.n243 71.676
R1062 B.n241 B.n240 71.676
R1063 B.n236 B.n235 71.676
R1064 B.n233 B.n232 71.676
R1065 B.n228 B.n227 71.676
R1066 B.n225 B.n224 71.676
R1067 B.n220 B.n144 71.676
R1068 B.n896 B.n895 71.676
R1069 B.n896 B.n2 71.676
R1070 B.n78 B.t17 69.0898
R1071 B.n188 B.t6 69.0898
R1072 B.n72 B.t11 69.063
R1073 B.n180 B.t13 69.063
R1074 B.n727 B.n72 59.5399
R1075 B.n79 B.n78 59.5399
R1076 B.n350 B.n188 59.5399
R1077 B.n181 B.n180 59.5399
R1078 B.n499 B.n145 52.1623
R1079 B.n859 B.n37 52.1623
R1080 B.n497 B.n496 30.7517
R1081 B.n501 B.n143 30.7517
R1082 B.n579 B.n578 30.7517
R1083 B.n857 B.n856 30.7517
R1084 B.n499 B.n141 29.8072
R1085 B.n505 B.n141 29.8072
R1086 B.n505 B.n136 29.8072
R1087 B.n511 B.n136 29.8072
R1088 B.n511 B.n137 29.8072
R1089 B.n517 B.n129 29.8072
R1090 B.n523 B.n129 29.8072
R1091 B.n523 B.n125 29.8072
R1092 B.n530 B.n125 29.8072
R1093 B.n530 B.n529 29.8072
R1094 B.n536 B.n118 29.8072
R1095 B.n544 B.n118 29.8072
R1096 B.n544 B.n543 29.8072
R1097 B.n550 B.n4 29.8072
R1098 B.n894 B.n4 29.8072
R1099 B.n894 B.n893 29.8072
R1100 B.n893 B.n892 29.8072
R1101 B.n892 B.n8 29.8072
R1102 B.n885 B.n12 29.8072
R1103 B.n885 B.n884 29.8072
R1104 B.n884 B.n883 29.8072
R1105 B.n877 B.n19 29.8072
R1106 B.n877 B.n876 29.8072
R1107 B.n876 B.n875 29.8072
R1108 B.n875 B.n23 29.8072
R1109 B.n869 B.n23 29.8072
R1110 B.n868 B.n867 29.8072
R1111 B.n867 B.n30 29.8072
R1112 B.n861 B.n30 29.8072
R1113 B.n861 B.n860 29.8072
R1114 B.n860 B.n859 29.8072
R1115 B.n517 B.t5 27.1772
R1116 B.n869 B.t9 27.1772
R1117 B.n550 B.t0 24.5472
R1118 B.t3 B.n8 24.5472
R1119 B.n72 B.n71 22.6914
R1120 B.n78 B.n77 22.6914
R1121 B.n188 B.n187 22.6914
R1122 B.n180 B.n179 22.6914
R1123 B.n529 B.t1 21.9172
R1124 B.n19 B.t2 21.9172
R1125 B B.n897 18.0485
R1126 B.n497 B.n139 10.6151
R1127 B.n507 B.n139 10.6151
R1128 B.n508 B.n507 10.6151
R1129 B.n509 B.n508 10.6151
R1130 B.n509 B.n131 10.6151
R1131 B.n519 B.n131 10.6151
R1132 B.n520 B.n519 10.6151
R1133 B.n521 B.n520 10.6151
R1134 B.n521 B.n123 10.6151
R1135 B.n532 B.n123 10.6151
R1136 B.n533 B.n532 10.6151
R1137 B.n534 B.n533 10.6151
R1138 B.n534 B.n116 10.6151
R1139 B.n546 B.n116 10.6151
R1140 B.n547 B.n546 10.6151
R1141 B.n548 B.n547 10.6151
R1142 B.n548 B.n0 10.6151
R1143 B.n496 B.n495 10.6151
R1144 B.n495 B.n147 10.6151
R1145 B.n490 B.n147 10.6151
R1146 B.n490 B.n489 10.6151
R1147 B.n489 B.n149 10.6151
R1148 B.n484 B.n149 10.6151
R1149 B.n484 B.n483 10.6151
R1150 B.n483 B.n482 10.6151
R1151 B.n482 B.n151 10.6151
R1152 B.n476 B.n151 10.6151
R1153 B.n476 B.n475 10.6151
R1154 B.n475 B.n474 10.6151
R1155 B.n474 B.n153 10.6151
R1156 B.n468 B.n153 10.6151
R1157 B.n468 B.n467 10.6151
R1158 B.n467 B.n466 10.6151
R1159 B.n466 B.n155 10.6151
R1160 B.n460 B.n155 10.6151
R1161 B.n460 B.n459 10.6151
R1162 B.n459 B.n458 10.6151
R1163 B.n458 B.n157 10.6151
R1164 B.n452 B.n157 10.6151
R1165 B.n452 B.n451 10.6151
R1166 B.n451 B.n450 10.6151
R1167 B.n450 B.n159 10.6151
R1168 B.n444 B.n159 10.6151
R1169 B.n444 B.n443 10.6151
R1170 B.n443 B.n442 10.6151
R1171 B.n442 B.n161 10.6151
R1172 B.n436 B.n161 10.6151
R1173 B.n436 B.n435 10.6151
R1174 B.n435 B.n434 10.6151
R1175 B.n434 B.n163 10.6151
R1176 B.n428 B.n163 10.6151
R1177 B.n428 B.n427 10.6151
R1178 B.n427 B.n426 10.6151
R1179 B.n426 B.n165 10.6151
R1180 B.n420 B.n165 10.6151
R1181 B.n420 B.n419 10.6151
R1182 B.n419 B.n418 10.6151
R1183 B.n418 B.n167 10.6151
R1184 B.n412 B.n167 10.6151
R1185 B.n412 B.n411 10.6151
R1186 B.n411 B.n410 10.6151
R1187 B.n410 B.n169 10.6151
R1188 B.n404 B.n169 10.6151
R1189 B.n404 B.n403 10.6151
R1190 B.n403 B.n402 10.6151
R1191 B.n402 B.n171 10.6151
R1192 B.n396 B.n171 10.6151
R1193 B.n396 B.n395 10.6151
R1194 B.n395 B.n394 10.6151
R1195 B.n394 B.n173 10.6151
R1196 B.n388 B.n173 10.6151
R1197 B.n388 B.n387 10.6151
R1198 B.n387 B.n386 10.6151
R1199 B.n386 B.n175 10.6151
R1200 B.n380 B.n175 10.6151
R1201 B.n380 B.n379 10.6151
R1202 B.n379 B.n378 10.6151
R1203 B.n378 B.n177 10.6151
R1204 B.n372 B.n177 10.6151
R1205 B.n372 B.n371 10.6151
R1206 B.n371 B.n370 10.6151
R1207 B.n366 B.n365 10.6151
R1208 B.n365 B.n183 10.6151
R1209 B.n360 B.n183 10.6151
R1210 B.n360 B.n359 10.6151
R1211 B.n359 B.n358 10.6151
R1212 B.n358 B.n185 10.6151
R1213 B.n352 B.n185 10.6151
R1214 B.n352 B.n351 10.6151
R1215 B.n349 B.n189 10.6151
R1216 B.n343 B.n189 10.6151
R1217 B.n343 B.n342 10.6151
R1218 B.n342 B.n341 10.6151
R1219 B.n341 B.n191 10.6151
R1220 B.n335 B.n191 10.6151
R1221 B.n335 B.n334 10.6151
R1222 B.n334 B.n333 10.6151
R1223 B.n333 B.n193 10.6151
R1224 B.n327 B.n193 10.6151
R1225 B.n327 B.n326 10.6151
R1226 B.n326 B.n325 10.6151
R1227 B.n325 B.n195 10.6151
R1228 B.n319 B.n195 10.6151
R1229 B.n319 B.n318 10.6151
R1230 B.n318 B.n317 10.6151
R1231 B.n317 B.n197 10.6151
R1232 B.n311 B.n197 10.6151
R1233 B.n311 B.n310 10.6151
R1234 B.n310 B.n309 10.6151
R1235 B.n309 B.n199 10.6151
R1236 B.n303 B.n199 10.6151
R1237 B.n303 B.n302 10.6151
R1238 B.n302 B.n301 10.6151
R1239 B.n301 B.n201 10.6151
R1240 B.n295 B.n201 10.6151
R1241 B.n295 B.n294 10.6151
R1242 B.n294 B.n293 10.6151
R1243 B.n293 B.n203 10.6151
R1244 B.n287 B.n203 10.6151
R1245 B.n287 B.n286 10.6151
R1246 B.n286 B.n285 10.6151
R1247 B.n285 B.n205 10.6151
R1248 B.n279 B.n205 10.6151
R1249 B.n279 B.n278 10.6151
R1250 B.n278 B.n277 10.6151
R1251 B.n277 B.n207 10.6151
R1252 B.n271 B.n207 10.6151
R1253 B.n271 B.n270 10.6151
R1254 B.n270 B.n269 10.6151
R1255 B.n269 B.n209 10.6151
R1256 B.n263 B.n209 10.6151
R1257 B.n263 B.n262 10.6151
R1258 B.n262 B.n261 10.6151
R1259 B.n261 B.n211 10.6151
R1260 B.n255 B.n211 10.6151
R1261 B.n255 B.n254 10.6151
R1262 B.n254 B.n253 10.6151
R1263 B.n253 B.n213 10.6151
R1264 B.n247 B.n213 10.6151
R1265 B.n247 B.n246 10.6151
R1266 B.n246 B.n245 10.6151
R1267 B.n245 B.n215 10.6151
R1268 B.n239 B.n215 10.6151
R1269 B.n239 B.n238 10.6151
R1270 B.n238 B.n237 10.6151
R1271 B.n237 B.n217 10.6151
R1272 B.n231 B.n217 10.6151
R1273 B.n231 B.n230 10.6151
R1274 B.n230 B.n229 10.6151
R1275 B.n229 B.n219 10.6151
R1276 B.n223 B.n219 10.6151
R1277 B.n223 B.n222 10.6151
R1278 B.n222 B.n143 10.6151
R1279 B.n502 B.n501 10.6151
R1280 B.n503 B.n502 10.6151
R1281 B.n503 B.n134 10.6151
R1282 B.n513 B.n134 10.6151
R1283 B.n514 B.n513 10.6151
R1284 B.n515 B.n514 10.6151
R1285 B.n515 B.n127 10.6151
R1286 B.n525 B.n127 10.6151
R1287 B.n526 B.n525 10.6151
R1288 B.n527 B.n526 10.6151
R1289 B.n527 B.n120 10.6151
R1290 B.n538 B.n120 10.6151
R1291 B.n539 B.n538 10.6151
R1292 B.n541 B.n539 10.6151
R1293 B.n541 B.n540 10.6151
R1294 B.n540 B.n113 10.6151
R1295 B.n553 B.n113 10.6151
R1296 B.n554 B.n553 10.6151
R1297 B.n555 B.n554 10.6151
R1298 B.n556 B.n555 10.6151
R1299 B.n557 B.n556 10.6151
R1300 B.n560 B.n557 10.6151
R1301 B.n561 B.n560 10.6151
R1302 B.n562 B.n561 10.6151
R1303 B.n563 B.n562 10.6151
R1304 B.n565 B.n563 10.6151
R1305 B.n566 B.n565 10.6151
R1306 B.n567 B.n566 10.6151
R1307 B.n568 B.n567 10.6151
R1308 B.n570 B.n568 10.6151
R1309 B.n571 B.n570 10.6151
R1310 B.n572 B.n571 10.6151
R1311 B.n573 B.n572 10.6151
R1312 B.n575 B.n573 10.6151
R1313 B.n576 B.n575 10.6151
R1314 B.n577 B.n576 10.6151
R1315 B.n578 B.n577 10.6151
R1316 B.n889 B.n1 10.6151
R1317 B.n889 B.n888 10.6151
R1318 B.n888 B.n887 10.6151
R1319 B.n887 B.n10 10.6151
R1320 B.n881 B.n10 10.6151
R1321 B.n881 B.n880 10.6151
R1322 B.n880 B.n879 10.6151
R1323 B.n879 B.n17 10.6151
R1324 B.n873 B.n17 10.6151
R1325 B.n873 B.n872 10.6151
R1326 B.n872 B.n871 10.6151
R1327 B.n871 B.n25 10.6151
R1328 B.n865 B.n25 10.6151
R1329 B.n865 B.n864 10.6151
R1330 B.n864 B.n863 10.6151
R1331 B.n863 B.n32 10.6151
R1332 B.n857 B.n32 10.6151
R1333 B.n856 B.n855 10.6151
R1334 B.n855 B.n39 10.6151
R1335 B.n849 B.n39 10.6151
R1336 B.n849 B.n848 10.6151
R1337 B.n848 B.n847 10.6151
R1338 B.n847 B.n41 10.6151
R1339 B.n841 B.n41 10.6151
R1340 B.n841 B.n840 10.6151
R1341 B.n840 B.n839 10.6151
R1342 B.n839 B.n43 10.6151
R1343 B.n833 B.n43 10.6151
R1344 B.n833 B.n832 10.6151
R1345 B.n832 B.n831 10.6151
R1346 B.n831 B.n45 10.6151
R1347 B.n825 B.n45 10.6151
R1348 B.n825 B.n824 10.6151
R1349 B.n824 B.n823 10.6151
R1350 B.n823 B.n47 10.6151
R1351 B.n817 B.n47 10.6151
R1352 B.n817 B.n816 10.6151
R1353 B.n816 B.n815 10.6151
R1354 B.n815 B.n49 10.6151
R1355 B.n809 B.n49 10.6151
R1356 B.n809 B.n808 10.6151
R1357 B.n808 B.n807 10.6151
R1358 B.n807 B.n51 10.6151
R1359 B.n801 B.n51 10.6151
R1360 B.n801 B.n800 10.6151
R1361 B.n800 B.n799 10.6151
R1362 B.n799 B.n53 10.6151
R1363 B.n793 B.n53 10.6151
R1364 B.n793 B.n792 10.6151
R1365 B.n792 B.n791 10.6151
R1366 B.n791 B.n55 10.6151
R1367 B.n785 B.n55 10.6151
R1368 B.n785 B.n784 10.6151
R1369 B.n784 B.n783 10.6151
R1370 B.n783 B.n57 10.6151
R1371 B.n777 B.n57 10.6151
R1372 B.n777 B.n776 10.6151
R1373 B.n776 B.n775 10.6151
R1374 B.n775 B.n59 10.6151
R1375 B.n769 B.n59 10.6151
R1376 B.n769 B.n768 10.6151
R1377 B.n768 B.n767 10.6151
R1378 B.n767 B.n61 10.6151
R1379 B.n761 B.n61 10.6151
R1380 B.n761 B.n760 10.6151
R1381 B.n760 B.n759 10.6151
R1382 B.n759 B.n63 10.6151
R1383 B.n753 B.n63 10.6151
R1384 B.n753 B.n752 10.6151
R1385 B.n752 B.n751 10.6151
R1386 B.n751 B.n65 10.6151
R1387 B.n745 B.n65 10.6151
R1388 B.n745 B.n744 10.6151
R1389 B.n744 B.n743 10.6151
R1390 B.n743 B.n67 10.6151
R1391 B.n737 B.n67 10.6151
R1392 B.n737 B.n736 10.6151
R1393 B.n736 B.n735 10.6151
R1394 B.n735 B.n69 10.6151
R1395 B.n729 B.n69 10.6151
R1396 B.n729 B.n728 10.6151
R1397 B.n726 B.n73 10.6151
R1398 B.n720 B.n73 10.6151
R1399 B.n720 B.n719 10.6151
R1400 B.n719 B.n718 10.6151
R1401 B.n718 B.n75 10.6151
R1402 B.n712 B.n75 10.6151
R1403 B.n712 B.n711 10.6151
R1404 B.n711 B.n710 10.6151
R1405 B.n706 B.n705 10.6151
R1406 B.n705 B.n81 10.6151
R1407 B.n700 B.n81 10.6151
R1408 B.n700 B.n699 10.6151
R1409 B.n699 B.n698 10.6151
R1410 B.n698 B.n83 10.6151
R1411 B.n692 B.n83 10.6151
R1412 B.n692 B.n691 10.6151
R1413 B.n691 B.n690 10.6151
R1414 B.n690 B.n85 10.6151
R1415 B.n684 B.n85 10.6151
R1416 B.n684 B.n683 10.6151
R1417 B.n683 B.n682 10.6151
R1418 B.n682 B.n87 10.6151
R1419 B.n676 B.n87 10.6151
R1420 B.n676 B.n675 10.6151
R1421 B.n675 B.n674 10.6151
R1422 B.n674 B.n89 10.6151
R1423 B.n668 B.n89 10.6151
R1424 B.n668 B.n667 10.6151
R1425 B.n667 B.n666 10.6151
R1426 B.n666 B.n91 10.6151
R1427 B.n660 B.n91 10.6151
R1428 B.n660 B.n659 10.6151
R1429 B.n659 B.n658 10.6151
R1430 B.n658 B.n93 10.6151
R1431 B.n652 B.n93 10.6151
R1432 B.n652 B.n651 10.6151
R1433 B.n651 B.n650 10.6151
R1434 B.n650 B.n95 10.6151
R1435 B.n644 B.n95 10.6151
R1436 B.n644 B.n643 10.6151
R1437 B.n643 B.n642 10.6151
R1438 B.n642 B.n97 10.6151
R1439 B.n636 B.n97 10.6151
R1440 B.n636 B.n635 10.6151
R1441 B.n635 B.n634 10.6151
R1442 B.n634 B.n99 10.6151
R1443 B.n628 B.n99 10.6151
R1444 B.n628 B.n627 10.6151
R1445 B.n627 B.n626 10.6151
R1446 B.n626 B.n101 10.6151
R1447 B.n620 B.n101 10.6151
R1448 B.n620 B.n619 10.6151
R1449 B.n619 B.n618 10.6151
R1450 B.n618 B.n103 10.6151
R1451 B.n612 B.n103 10.6151
R1452 B.n612 B.n611 10.6151
R1453 B.n611 B.n610 10.6151
R1454 B.n610 B.n105 10.6151
R1455 B.n604 B.n105 10.6151
R1456 B.n604 B.n603 10.6151
R1457 B.n603 B.n602 10.6151
R1458 B.n602 B.n107 10.6151
R1459 B.n596 B.n107 10.6151
R1460 B.n596 B.n595 10.6151
R1461 B.n595 B.n594 10.6151
R1462 B.n594 B.n109 10.6151
R1463 B.n588 B.n109 10.6151
R1464 B.n588 B.n587 10.6151
R1465 B.n587 B.n586 10.6151
R1466 B.n586 B.n111 10.6151
R1467 B.n580 B.n111 10.6151
R1468 B.n580 B.n579 10.6151
R1469 B.n897 B.n0 8.11757
R1470 B.n897 B.n1 8.11757
R1471 B.n536 B.t1 7.89052
R1472 B.n883 B.t2 7.89052
R1473 B.n366 B.n181 6.5566
R1474 B.n351 B.n350 6.5566
R1475 B.n727 B.n726 6.5566
R1476 B.n710 B.n79 6.5566
R1477 B.n543 B.t0 5.26051
R1478 B.n12 B.t3 5.26051
R1479 B.n370 B.n181 4.05904
R1480 B.n350 B.n349 4.05904
R1481 B.n728 B.n727 4.05904
R1482 B.n706 B.n79 4.05904
R1483 B.n137 B.t5 2.63051
R1484 B.t9 B.n868 2.63051
R1485 VN.n0 VN.t1 636.408
R1486 VN.n1 VN.t2 636.408
R1487 VN.n0 VN.t0 636.357
R1488 VN.n1 VN.t3 636.357
R1489 VN VN.n1 91.9064
R1490 VN VN.n0 44.7132
R1491 VTAIL.n5 VTAIL.t0 47.2402
R1492 VTAIL.n4 VTAIL.t5 47.2402
R1493 VTAIL.n3 VTAIL.t7 47.2402
R1494 VTAIL.n7 VTAIL.t4 47.24
R1495 VTAIL.n0 VTAIL.t6 47.24
R1496 VTAIL.n1 VTAIL.t1 47.24
R1497 VTAIL.n2 VTAIL.t2 47.24
R1498 VTAIL.n6 VTAIL.t3 47.24
R1499 VTAIL.n7 VTAIL.n6 30.4617
R1500 VTAIL.n3 VTAIL.n2 30.4617
R1501 VTAIL.n4 VTAIL.n3 1.00912
R1502 VTAIL.n6 VTAIL.n5 1.00912
R1503 VTAIL.n2 VTAIL.n1 1.00912
R1504 VTAIL VTAIL.n0 0.563
R1505 VTAIL.n5 VTAIL.n4 0.470328
R1506 VTAIL.n1 VTAIL.n0 0.470328
R1507 VTAIL VTAIL.n7 0.446621
R1508 VDD2.n2 VDD2.n0 106.746
R1509 VDD2.n2 VDD2.n1 62.9198
R1510 VDD2.n1 VDD2.t0 0.999491
R1511 VDD2.n1 VDD2.t1 0.999491
R1512 VDD2.n0 VDD2.t2 0.999491
R1513 VDD2.n0 VDD2.t3 0.999491
R1514 VDD2 VDD2.n2 0.0586897
R1515 VP.n1 VP.t0 636.408
R1516 VP.n1 VP.t1 636.357
R1517 VP.n3 VP.t2 615.412
R1518 VP.n5 VP.t3 615.412
R1519 VP.n6 VP.n5 161.3
R1520 VP.n4 VP.n0 161.3
R1521 VP.n3 VP.n2 161.3
R1522 VP.n2 VP.n1 91.5257
R1523 VP.n4 VP.n3 24.1005
R1524 VP.n5 VP.n4 24.1005
R1525 VP.n2 VP.n0 0.189894
R1526 VP.n6 VP.n0 0.189894
R1527 VP VP.n6 0.0516364
R1528 VDD1 VDD1.n1 107.272
R1529 VDD1 VDD1.n0 62.978
R1530 VDD1.n0 VDD1.t3 0.999491
R1531 VDD1.n0 VDD1.t2 0.999491
R1532 VDD1.n1 VDD1.t1 0.999491
R1533 VDD1.n1 VDD1.t0 0.999491
C0 VTAIL VDD2 9.57446f
C1 VN VDD1 0.147551f
C2 VTAIL VP 4.792871f
C3 VDD2 VDD1 0.598778f
C4 VDD1 VP 5.59677f
C5 VTAIL VDD1 9.53205f
C6 VDD2 VN 5.46216f
C7 VN VP 6.36592f
C8 VTAIL VN 4.77877f
C9 VDD2 VP 0.282455f
C10 VDD2 B 3.389575f
C11 VDD1 B 7.97728f
C12 VTAIL B 13.374765f
C13 VN B 9.39625f
C14 VP B 5.719239f
C15 VDD1.t3 B 0.433543f
C16 VDD1.t2 B 0.433543f
C17 VDD1.n0 B 3.97318f
C18 VDD1.t1 B 0.433543f
C19 VDD1.t0 B 0.433543f
C20 VDD1.n1 B 4.88155f
C21 VP.n0 B 0.046302f
C22 VP.t1 B 2.20999f
C23 VP.t0 B 2.21005f
C24 VP.n1 B 2.79755f
C25 VP.n2 B 3.48002f
C26 VP.t2 B 2.18324f
C27 VP.n3 B 0.809117f
C28 VP.n4 B 0.010507f
C29 VP.t3 B 2.18324f
C30 VP.n5 B 0.809117f
C31 VP.n6 B 0.035882f
C32 VDD2.t2 B 0.436498f
C33 VDD2.t3 B 0.436498f
C34 VDD2.n0 B 4.88567f
C35 VDD2.t0 B 0.436498f
C36 VDD2.t1 B 0.436498f
C37 VDD2.n1 B 3.99996f
C38 VDD2.n2 B 4.37181f
C39 VTAIL.t6 B 2.7707f
C40 VTAIL.n0 B 0.252592f
C41 VTAIL.t1 B 2.7707f
C42 VTAIL.n1 B 0.274736f
C43 VTAIL.t2 B 2.7707f
C44 VTAIL.n2 B 1.35886f
C45 VTAIL.t7 B 2.7707f
C46 VTAIL.n3 B 1.35886f
C47 VTAIL.t5 B 2.7707f
C48 VTAIL.n4 B 0.274736f
C49 VTAIL.t0 B 2.7707f
C50 VTAIL.n5 B 0.274736f
C51 VTAIL.t3 B 2.7707f
C52 VTAIL.n6 B 1.35886f
C53 VTAIL.t4 B 2.7707f
C54 VTAIL.n7 B 1.33093f
C55 VN.t1 B 2.18842f
C56 VN.t0 B 2.18835f
C57 VN.n0 B 1.56027f
C58 VN.t2 B 2.18842f
C59 VN.t3 B 2.18835f
C60 VN.n1 B 2.79032f
.ends

