* NGSPICE file created from diff_pair_sample_0206.ext - technology: sky130A

.subckt diff_pair_sample_0206 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=0.4134 pd=2.9 as=0.1749 ps=1.39 w=1.06 l=2.14
X1 VDD1.t4 VP.t1 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=0.1749 pd=1.39 as=0.4134 ps=2.9 w=1.06 l=2.14
X2 VTAIL.t1 VN.t0 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.1749 pd=1.39 as=0.1749 ps=1.39 w=1.06 l=2.14
X3 VDD2.t4 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.4134 pd=2.9 as=0.1749 ps=1.39 w=1.06 l=2.14
X4 VDD1.t3 VP.t2 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=0.4134 pd=2.9 as=0.1749 ps=1.39 w=1.06 l=2.14
X5 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=0.4134 pd=2.9 as=0 ps=0 w=1.06 l=2.14
X6 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=0.4134 pd=2.9 as=0 ps=0 w=1.06 l=2.14
X7 VTAIL.t3 VN.t2 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.1749 pd=1.39 as=0.1749 ps=1.39 w=1.06 l=2.14
X8 VTAIL.t6 VP.t3 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=0.1749 pd=1.39 as=0.1749 ps=1.39 w=1.06 l=2.14
X9 VDD2.t2 VN.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.4134 pd=2.9 as=0.1749 ps=1.39 w=1.06 l=2.14
X10 VDD2.t1 VN.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.1749 pd=1.39 as=0.4134 ps=2.9 w=1.06 l=2.14
X11 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.4134 pd=2.9 as=0 ps=0 w=1.06 l=2.14
X12 VDD2.t0 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.1749 pd=1.39 as=0.4134 ps=2.9 w=1.06 l=2.14
X13 VDD1.t1 VP.t4 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=0.1749 pd=1.39 as=0.4134 ps=2.9 w=1.06 l=2.14
X14 VTAIL.t9 VP.t5 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.1749 pd=1.39 as=0.1749 ps=1.39 w=1.06 l=2.14
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.4134 pd=2.9 as=0 ps=0 w=1.06 l=2.14
R0 VP.n10 VP.n9 161.3
R1 VP.n11 VP.n6 161.3
R2 VP.n13 VP.n12 161.3
R3 VP.n14 VP.n5 161.3
R4 VP.n31 VP.n0 161.3
R5 VP.n30 VP.n29 161.3
R6 VP.n28 VP.n1 161.3
R7 VP.n27 VP.n26 161.3
R8 VP.n25 VP.n2 161.3
R9 VP.n24 VP.n23 161.3
R10 VP.n22 VP.n3 161.3
R11 VP.n21 VP.n20 161.3
R12 VP.n19 VP.n4 161.3
R13 VP.n18 VP.n17 87.7234
R14 VP.n33 VP.n32 87.7234
R15 VP.n16 VP.n15 87.7234
R16 VP.n20 VP.n3 56.4773
R17 VP.n30 VP.n1 56.4773
R18 VP.n13 VP.n6 56.4773
R19 VP.n7 VP.t2 46.4527
R20 VP.n8 VP.n7 46.2445
R21 VP.n17 VP.n16 38.6927
R22 VP.n20 VP.n19 24.3439
R23 VP.n24 VP.n3 24.3439
R24 VP.n25 VP.n24 24.3439
R25 VP.n26 VP.n25 24.3439
R26 VP.n26 VP.n1 24.3439
R27 VP.n31 VP.n30 24.3439
R28 VP.n14 VP.n13 24.3439
R29 VP.n9 VP.n8 24.3439
R30 VP.n9 VP.n6 24.3439
R31 VP.n19 VP.n18 22.8833
R32 VP.n32 VP.n31 22.8833
R33 VP.n15 VP.n14 22.8833
R34 VP.n25 VP.t5 11.9379
R35 VP.n18 VP.t0 11.9379
R36 VP.n32 VP.t4 11.9379
R37 VP.n8 VP.t3 11.9379
R38 VP.n15 VP.t1 11.9379
R39 VP.n10 VP.n7 8.71313
R40 VP.n16 VP.n5 0.278398
R41 VP.n17 VP.n4 0.278398
R42 VP.n33 VP.n0 0.278398
R43 VP.n11 VP.n10 0.189894
R44 VP.n12 VP.n11 0.189894
R45 VP.n12 VP.n5 0.189894
R46 VP.n21 VP.n4 0.189894
R47 VP.n22 VP.n21 0.189894
R48 VP.n23 VP.n22 0.189894
R49 VP.n23 VP.n2 0.189894
R50 VP.n27 VP.n2 0.189894
R51 VP.n28 VP.n27 0.189894
R52 VP.n29 VP.n28 0.189894
R53 VP.n29 VP.n0 0.189894
R54 VP VP.n33 0.153422
R55 VTAIL.n7 VTAIL.t5 154.946
R56 VTAIL.n11 VTAIL.t0 154.946
R57 VTAIL.n2 VTAIL.t7 154.946
R58 VTAIL.n10 VTAIL.t10 154.946
R59 VTAIL.n1 VTAIL.n0 128.784
R60 VTAIL.n4 VTAIL.n3 128.784
R61 VTAIL.n9 VTAIL.n8 128.782
R62 VTAIL.n6 VTAIL.n5 128.782
R63 VTAIL.n0 VTAIL.t2 18.6797
R64 VTAIL.n0 VTAIL.t3 18.6797
R65 VTAIL.n3 VTAIL.t11 18.6797
R66 VTAIL.n3 VTAIL.t9 18.6797
R67 VTAIL.n8 VTAIL.t8 18.6797
R68 VTAIL.n8 VTAIL.t6 18.6797
R69 VTAIL.n5 VTAIL.t4 18.6797
R70 VTAIL.n5 VTAIL.t1 18.6797
R71 VTAIL.n6 VTAIL.n4 17.5393
R72 VTAIL.n11 VTAIL.n10 15.41
R73 VTAIL.n7 VTAIL.n6 2.12981
R74 VTAIL.n10 VTAIL.n9 2.12981
R75 VTAIL.n4 VTAIL.n2 2.12981
R76 VTAIL VTAIL.n11 1.53929
R77 VTAIL.n9 VTAIL.n7 1.53498
R78 VTAIL.n2 VTAIL.n1 1.53498
R79 VTAIL VTAIL.n1 0.591017
R80 VDD1 VDD1.t3 173.28
R81 VDD1.n1 VDD1.t5 173.167
R82 VDD1.n1 VDD1.n0 145.94
R83 VDD1.n3 VDD1.n2 145.463
R84 VDD1.n3 VDD1.n1 33.197
R85 VDD1.n2 VDD1.t2 18.6797
R86 VDD1.n2 VDD1.t4 18.6797
R87 VDD1.n0 VDD1.t0 18.6797
R88 VDD1.n0 VDD1.t1 18.6797
R89 VDD1 VDD1.n3 0.474638
R90 B.n449 B.n448 585
R91 B.n142 B.n83 585
R92 B.n141 B.n140 585
R93 B.n139 B.n138 585
R94 B.n137 B.n136 585
R95 B.n135 B.n134 585
R96 B.n133 B.n132 585
R97 B.n131 B.n130 585
R98 B.n129 B.n128 585
R99 B.n126 B.n125 585
R100 B.n124 B.n123 585
R101 B.n122 B.n121 585
R102 B.n120 B.n119 585
R103 B.n118 B.n117 585
R104 B.n116 B.n115 585
R105 B.n114 B.n113 585
R106 B.n112 B.n111 585
R107 B.n110 B.n109 585
R108 B.n108 B.n107 585
R109 B.n105 B.n104 585
R110 B.n103 B.n102 585
R111 B.n101 B.n100 585
R112 B.n99 B.n98 585
R113 B.n97 B.n96 585
R114 B.n95 B.n94 585
R115 B.n93 B.n92 585
R116 B.n91 B.n90 585
R117 B.n89 B.n88 585
R118 B.n447 B.n69 585
R119 B.n452 B.n69 585
R120 B.n446 B.n68 585
R121 B.n453 B.n68 585
R122 B.n445 B.n444 585
R123 B.n444 B.n64 585
R124 B.n443 B.n63 585
R125 B.n459 B.n63 585
R126 B.n442 B.n62 585
R127 B.n460 B.n62 585
R128 B.n441 B.n61 585
R129 B.n461 B.n61 585
R130 B.n440 B.n439 585
R131 B.n439 B.n60 585
R132 B.n438 B.n56 585
R133 B.n467 B.n56 585
R134 B.n437 B.n55 585
R135 B.n468 B.n55 585
R136 B.n436 B.n54 585
R137 B.n469 B.n54 585
R138 B.n435 B.n434 585
R139 B.n434 B.n50 585
R140 B.n433 B.n49 585
R141 B.n475 B.n49 585
R142 B.n432 B.n48 585
R143 B.n476 B.n48 585
R144 B.n431 B.n47 585
R145 B.n477 B.n47 585
R146 B.n430 B.n429 585
R147 B.n429 B.n43 585
R148 B.n428 B.n42 585
R149 B.n483 B.n42 585
R150 B.n427 B.n41 585
R151 B.n484 B.n41 585
R152 B.n426 B.n40 585
R153 B.n485 B.n40 585
R154 B.n425 B.n424 585
R155 B.n424 B.n36 585
R156 B.n423 B.n35 585
R157 B.n491 B.n35 585
R158 B.n422 B.n34 585
R159 B.n492 B.n34 585
R160 B.n421 B.n33 585
R161 B.n493 B.n33 585
R162 B.n420 B.n419 585
R163 B.n419 B.n29 585
R164 B.n418 B.n28 585
R165 B.n499 B.n28 585
R166 B.n417 B.n27 585
R167 B.n500 B.n27 585
R168 B.n416 B.n26 585
R169 B.n501 B.n26 585
R170 B.n415 B.n414 585
R171 B.n414 B.n22 585
R172 B.n413 B.n21 585
R173 B.n507 B.n21 585
R174 B.n412 B.n20 585
R175 B.n508 B.n20 585
R176 B.n411 B.n19 585
R177 B.n509 B.n19 585
R178 B.n410 B.n409 585
R179 B.n409 B.n15 585
R180 B.n408 B.n14 585
R181 B.n515 B.n14 585
R182 B.n407 B.n13 585
R183 B.n516 B.n13 585
R184 B.n406 B.n12 585
R185 B.n517 B.n12 585
R186 B.n405 B.n404 585
R187 B.n404 B.n8 585
R188 B.n403 B.n7 585
R189 B.n523 B.n7 585
R190 B.n402 B.n6 585
R191 B.n524 B.n6 585
R192 B.n401 B.n5 585
R193 B.n525 B.n5 585
R194 B.n400 B.n399 585
R195 B.n399 B.n4 585
R196 B.n398 B.n143 585
R197 B.n398 B.n397 585
R198 B.n388 B.n144 585
R199 B.n145 B.n144 585
R200 B.n390 B.n389 585
R201 B.n391 B.n390 585
R202 B.n387 B.n150 585
R203 B.n150 B.n149 585
R204 B.n386 B.n385 585
R205 B.n385 B.n384 585
R206 B.n152 B.n151 585
R207 B.n153 B.n152 585
R208 B.n377 B.n376 585
R209 B.n378 B.n377 585
R210 B.n375 B.n158 585
R211 B.n158 B.n157 585
R212 B.n374 B.n373 585
R213 B.n373 B.n372 585
R214 B.n160 B.n159 585
R215 B.n161 B.n160 585
R216 B.n365 B.n364 585
R217 B.n366 B.n365 585
R218 B.n363 B.n165 585
R219 B.n169 B.n165 585
R220 B.n362 B.n361 585
R221 B.n361 B.n360 585
R222 B.n167 B.n166 585
R223 B.n168 B.n167 585
R224 B.n353 B.n352 585
R225 B.n354 B.n353 585
R226 B.n351 B.n174 585
R227 B.n174 B.n173 585
R228 B.n350 B.n349 585
R229 B.n349 B.n348 585
R230 B.n176 B.n175 585
R231 B.n177 B.n176 585
R232 B.n341 B.n340 585
R233 B.n342 B.n341 585
R234 B.n339 B.n182 585
R235 B.n182 B.n181 585
R236 B.n338 B.n337 585
R237 B.n337 B.n336 585
R238 B.n184 B.n183 585
R239 B.n185 B.n184 585
R240 B.n329 B.n328 585
R241 B.n330 B.n329 585
R242 B.n327 B.n190 585
R243 B.n190 B.n189 585
R244 B.n326 B.n325 585
R245 B.n325 B.n324 585
R246 B.n192 B.n191 585
R247 B.n193 B.n192 585
R248 B.n317 B.n316 585
R249 B.n318 B.n317 585
R250 B.n315 B.n198 585
R251 B.n198 B.n197 585
R252 B.n314 B.n313 585
R253 B.n313 B.n312 585
R254 B.n200 B.n199 585
R255 B.n305 B.n200 585
R256 B.n304 B.n303 585
R257 B.n306 B.n304 585
R258 B.n302 B.n205 585
R259 B.n205 B.n204 585
R260 B.n301 B.n300 585
R261 B.n300 B.n299 585
R262 B.n207 B.n206 585
R263 B.n208 B.n207 585
R264 B.n292 B.n291 585
R265 B.n293 B.n292 585
R266 B.n290 B.n213 585
R267 B.n213 B.n212 585
R268 B.n285 B.n284 585
R269 B.n283 B.n229 585
R270 B.n282 B.n228 585
R271 B.n287 B.n228 585
R272 B.n281 B.n280 585
R273 B.n279 B.n278 585
R274 B.n277 B.n276 585
R275 B.n275 B.n274 585
R276 B.n273 B.n272 585
R277 B.n271 B.n270 585
R278 B.n269 B.n268 585
R279 B.n267 B.n266 585
R280 B.n265 B.n264 585
R281 B.n263 B.n262 585
R282 B.n261 B.n260 585
R283 B.n259 B.n258 585
R284 B.n257 B.n256 585
R285 B.n255 B.n254 585
R286 B.n253 B.n252 585
R287 B.n251 B.n250 585
R288 B.n249 B.n248 585
R289 B.n247 B.n246 585
R290 B.n245 B.n244 585
R291 B.n243 B.n242 585
R292 B.n241 B.n240 585
R293 B.n239 B.n238 585
R294 B.n237 B.n236 585
R295 B.n215 B.n214 585
R296 B.n289 B.n288 585
R297 B.n288 B.n287 585
R298 B.n211 B.n210 585
R299 B.n212 B.n211 585
R300 B.n295 B.n294 585
R301 B.n294 B.n293 585
R302 B.n296 B.n209 585
R303 B.n209 B.n208 585
R304 B.n298 B.n297 585
R305 B.n299 B.n298 585
R306 B.n203 B.n202 585
R307 B.n204 B.n203 585
R308 B.n308 B.n307 585
R309 B.n307 B.n306 585
R310 B.n309 B.n201 585
R311 B.n305 B.n201 585
R312 B.n311 B.n310 585
R313 B.n312 B.n311 585
R314 B.n196 B.n195 585
R315 B.n197 B.n196 585
R316 B.n320 B.n319 585
R317 B.n319 B.n318 585
R318 B.n321 B.n194 585
R319 B.n194 B.n193 585
R320 B.n323 B.n322 585
R321 B.n324 B.n323 585
R322 B.n188 B.n187 585
R323 B.n189 B.n188 585
R324 B.n332 B.n331 585
R325 B.n331 B.n330 585
R326 B.n333 B.n186 585
R327 B.n186 B.n185 585
R328 B.n335 B.n334 585
R329 B.n336 B.n335 585
R330 B.n180 B.n179 585
R331 B.n181 B.n180 585
R332 B.n344 B.n343 585
R333 B.n343 B.n342 585
R334 B.n345 B.n178 585
R335 B.n178 B.n177 585
R336 B.n347 B.n346 585
R337 B.n348 B.n347 585
R338 B.n172 B.n171 585
R339 B.n173 B.n172 585
R340 B.n356 B.n355 585
R341 B.n355 B.n354 585
R342 B.n357 B.n170 585
R343 B.n170 B.n168 585
R344 B.n359 B.n358 585
R345 B.n360 B.n359 585
R346 B.n164 B.n163 585
R347 B.n169 B.n164 585
R348 B.n368 B.n367 585
R349 B.n367 B.n366 585
R350 B.n369 B.n162 585
R351 B.n162 B.n161 585
R352 B.n371 B.n370 585
R353 B.n372 B.n371 585
R354 B.n156 B.n155 585
R355 B.n157 B.n156 585
R356 B.n380 B.n379 585
R357 B.n379 B.n378 585
R358 B.n381 B.n154 585
R359 B.n154 B.n153 585
R360 B.n383 B.n382 585
R361 B.n384 B.n383 585
R362 B.n148 B.n147 585
R363 B.n149 B.n148 585
R364 B.n393 B.n392 585
R365 B.n392 B.n391 585
R366 B.n394 B.n146 585
R367 B.n146 B.n145 585
R368 B.n396 B.n395 585
R369 B.n397 B.n396 585
R370 B.n2 B.n0 585
R371 B.n4 B.n2 585
R372 B.n3 B.n1 585
R373 B.n524 B.n3 585
R374 B.n522 B.n521 585
R375 B.n523 B.n522 585
R376 B.n520 B.n9 585
R377 B.n9 B.n8 585
R378 B.n519 B.n518 585
R379 B.n518 B.n517 585
R380 B.n11 B.n10 585
R381 B.n516 B.n11 585
R382 B.n514 B.n513 585
R383 B.n515 B.n514 585
R384 B.n512 B.n16 585
R385 B.n16 B.n15 585
R386 B.n511 B.n510 585
R387 B.n510 B.n509 585
R388 B.n18 B.n17 585
R389 B.n508 B.n18 585
R390 B.n506 B.n505 585
R391 B.n507 B.n506 585
R392 B.n504 B.n23 585
R393 B.n23 B.n22 585
R394 B.n503 B.n502 585
R395 B.n502 B.n501 585
R396 B.n25 B.n24 585
R397 B.n500 B.n25 585
R398 B.n498 B.n497 585
R399 B.n499 B.n498 585
R400 B.n496 B.n30 585
R401 B.n30 B.n29 585
R402 B.n495 B.n494 585
R403 B.n494 B.n493 585
R404 B.n32 B.n31 585
R405 B.n492 B.n32 585
R406 B.n490 B.n489 585
R407 B.n491 B.n490 585
R408 B.n488 B.n37 585
R409 B.n37 B.n36 585
R410 B.n487 B.n486 585
R411 B.n486 B.n485 585
R412 B.n39 B.n38 585
R413 B.n484 B.n39 585
R414 B.n482 B.n481 585
R415 B.n483 B.n482 585
R416 B.n480 B.n44 585
R417 B.n44 B.n43 585
R418 B.n479 B.n478 585
R419 B.n478 B.n477 585
R420 B.n46 B.n45 585
R421 B.n476 B.n46 585
R422 B.n474 B.n473 585
R423 B.n475 B.n474 585
R424 B.n472 B.n51 585
R425 B.n51 B.n50 585
R426 B.n471 B.n470 585
R427 B.n470 B.n469 585
R428 B.n53 B.n52 585
R429 B.n468 B.n53 585
R430 B.n466 B.n465 585
R431 B.n467 B.n466 585
R432 B.n464 B.n57 585
R433 B.n60 B.n57 585
R434 B.n463 B.n462 585
R435 B.n462 B.n461 585
R436 B.n59 B.n58 585
R437 B.n460 B.n59 585
R438 B.n458 B.n457 585
R439 B.n459 B.n458 585
R440 B.n456 B.n65 585
R441 B.n65 B.n64 585
R442 B.n455 B.n454 585
R443 B.n454 B.n453 585
R444 B.n67 B.n66 585
R445 B.n452 B.n67 585
R446 B.n527 B.n526 585
R447 B.n526 B.n525 585
R448 B.n285 B.n211 564.573
R449 B.n88 B.n67 564.573
R450 B.n288 B.n213 564.573
R451 B.n449 B.n69 564.573
R452 B.n451 B.n450 256.663
R453 B.n451 B.n82 256.663
R454 B.n451 B.n81 256.663
R455 B.n451 B.n80 256.663
R456 B.n451 B.n79 256.663
R457 B.n451 B.n78 256.663
R458 B.n451 B.n77 256.663
R459 B.n451 B.n76 256.663
R460 B.n451 B.n75 256.663
R461 B.n451 B.n74 256.663
R462 B.n451 B.n73 256.663
R463 B.n451 B.n72 256.663
R464 B.n451 B.n71 256.663
R465 B.n451 B.n70 256.663
R466 B.n287 B.n286 256.663
R467 B.n287 B.n216 256.663
R468 B.n287 B.n217 256.663
R469 B.n287 B.n218 256.663
R470 B.n287 B.n219 256.663
R471 B.n287 B.n220 256.663
R472 B.n287 B.n221 256.663
R473 B.n287 B.n222 256.663
R474 B.n287 B.n223 256.663
R475 B.n287 B.n224 256.663
R476 B.n287 B.n225 256.663
R477 B.n287 B.n226 256.663
R478 B.n287 B.n227 256.663
R479 B.n287 B.n212 234.412
R480 B.n452 B.n451 234.412
R481 B.n233 B.t14 208.225
R482 B.n230 B.t10 208.225
R483 B.n86 B.t6 208.225
R484 B.n84 B.t17 208.225
R485 B.n230 B.t13 193.427
R486 B.n86 B.t8 193.427
R487 B.n233 B.t16 193.427
R488 B.n84 B.t18 193.427
R489 B.n294 B.n211 163.367
R490 B.n294 B.n209 163.367
R491 B.n298 B.n209 163.367
R492 B.n298 B.n203 163.367
R493 B.n307 B.n203 163.367
R494 B.n307 B.n201 163.367
R495 B.n311 B.n201 163.367
R496 B.n311 B.n196 163.367
R497 B.n319 B.n196 163.367
R498 B.n319 B.n194 163.367
R499 B.n323 B.n194 163.367
R500 B.n323 B.n188 163.367
R501 B.n331 B.n188 163.367
R502 B.n331 B.n186 163.367
R503 B.n335 B.n186 163.367
R504 B.n335 B.n180 163.367
R505 B.n343 B.n180 163.367
R506 B.n343 B.n178 163.367
R507 B.n347 B.n178 163.367
R508 B.n347 B.n172 163.367
R509 B.n355 B.n172 163.367
R510 B.n355 B.n170 163.367
R511 B.n359 B.n170 163.367
R512 B.n359 B.n164 163.367
R513 B.n367 B.n164 163.367
R514 B.n367 B.n162 163.367
R515 B.n371 B.n162 163.367
R516 B.n371 B.n156 163.367
R517 B.n379 B.n156 163.367
R518 B.n379 B.n154 163.367
R519 B.n383 B.n154 163.367
R520 B.n383 B.n148 163.367
R521 B.n392 B.n148 163.367
R522 B.n392 B.n146 163.367
R523 B.n396 B.n146 163.367
R524 B.n396 B.n2 163.367
R525 B.n526 B.n2 163.367
R526 B.n526 B.n3 163.367
R527 B.n522 B.n3 163.367
R528 B.n522 B.n9 163.367
R529 B.n518 B.n9 163.367
R530 B.n518 B.n11 163.367
R531 B.n514 B.n11 163.367
R532 B.n514 B.n16 163.367
R533 B.n510 B.n16 163.367
R534 B.n510 B.n18 163.367
R535 B.n506 B.n18 163.367
R536 B.n506 B.n23 163.367
R537 B.n502 B.n23 163.367
R538 B.n502 B.n25 163.367
R539 B.n498 B.n25 163.367
R540 B.n498 B.n30 163.367
R541 B.n494 B.n30 163.367
R542 B.n494 B.n32 163.367
R543 B.n490 B.n32 163.367
R544 B.n490 B.n37 163.367
R545 B.n486 B.n37 163.367
R546 B.n486 B.n39 163.367
R547 B.n482 B.n39 163.367
R548 B.n482 B.n44 163.367
R549 B.n478 B.n44 163.367
R550 B.n478 B.n46 163.367
R551 B.n474 B.n46 163.367
R552 B.n474 B.n51 163.367
R553 B.n470 B.n51 163.367
R554 B.n470 B.n53 163.367
R555 B.n466 B.n53 163.367
R556 B.n466 B.n57 163.367
R557 B.n462 B.n57 163.367
R558 B.n462 B.n59 163.367
R559 B.n458 B.n59 163.367
R560 B.n458 B.n65 163.367
R561 B.n454 B.n65 163.367
R562 B.n454 B.n67 163.367
R563 B.n229 B.n228 163.367
R564 B.n280 B.n228 163.367
R565 B.n278 B.n277 163.367
R566 B.n274 B.n273 163.367
R567 B.n270 B.n269 163.367
R568 B.n266 B.n265 163.367
R569 B.n262 B.n261 163.367
R570 B.n258 B.n257 163.367
R571 B.n254 B.n253 163.367
R572 B.n250 B.n249 163.367
R573 B.n246 B.n245 163.367
R574 B.n242 B.n241 163.367
R575 B.n238 B.n237 163.367
R576 B.n288 B.n215 163.367
R577 B.n292 B.n213 163.367
R578 B.n292 B.n207 163.367
R579 B.n300 B.n207 163.367
R580 B.n300 B.n205 163.367
R581 B.n304 B.n205 163.367
R582 B.n304 B.n200 163.367
R583 B.n313 B.n200 163.367
R584 B.n313 B.n198 163.367
R585 B.n317 B.n198 163.367
R586 B.n317 B.n192 163.367
R587 B.n325 B.n192 163.367
R588 B.n325 B.n190 163.367
R589 B.n329 B.n190 163.367
R590 B.n329 B.n184 163.367
R591 B.n337 B.n184 163.367
R592 B.n337 B.n182 163.367
R593 B.n341 B.n182 163.367
R594 B.n341 B.n176 163.367
R595 B.n349 B.n176 163.367
R596 B.n349 B.n174 163.367
R597 B.n353 B.n174 163.367
R598 B.n353 B.n167 163.367
R599 B.n361 B.n167 163.367
R600 B.n361 B.n165 163.367
R601 B.n365 B.n165 163.367
R602 B.n365 B.n160 163.367
R603 B.n373 B.n160 163.367
R604 B.n373 B.n158 163.367
R605 B.n377 B.n158 163.367
R606 B.n377 B.n152 163.367
R607 B.n385 B.n152 163.367
R608 B.n385 B.n150 163.367
R609 B.n390 B.n150 163.367
R610 B.n390 B.n144 163.367
R611 B.n398 B.n144 163.367
R612 B.n399 B.n398 163.367
R613 B.n399 B.n5 163.367
R614 B.n6 B.n5 163.367
R615 B.n7 B.n6 163.367
R616 B.n404 B.n7 163.367
R617 B.n404 B.n12 163.367
R618 B.n13 B.n12 163.367
R619 B.n14 B.n13 163.367
R620 B.n409 B.n14 163.367
R621 B.n409 B.n19 163.367
R622 B.n20 B.n19 163.367
R623 B.n21 B.n20 163.367
R624 B.n414 B.n21 163.367
R625 B.n414 B.n26 163.367
R626 B.n27 B.n26 163.367
R627 B.n28 B.n27 163.367
R628 B.n419 B.n28 163.367
R629 B.n419 B.n33 163.367
R630 B.n34 B.n33 163.367
R631 B.n35 B.n34 163.367
R632 B.n424 B.n35 163.367
R633 B.n424 B.n40 163.367
R634 B.n41 B.n40 163.367
R635 B.n42 B.n41 163.367
R636 B.n429 B.n42 163.367
R637 B.n429 B.n47 163.367
R638 B.n48 B.n47 163.367
R639 B.n49 B.n48 163.367
R640 B.n434 B.n49 163.367
R641 B.n434 B.n54 163.367
R642 B.n55 B.n54 163.367
R643 B.n56 B.n55 163.367
R644 B.n439 B.n56 163.367
R645 B.n439 B.n61 163.367
R646 B.n62 B.n61 163.367
R647 B.n63 B.n62 163.367
R648 B.n444 B.n63 163.367
R649 B.n444 B.n68 163.367
R650 B.n69 B.n68 163.367
R651 B.n92 B.n91 163.367
R652 B.n96 B.n95 163.367
R653 B.n100 B.n99 163.367
R654 B.n104 B.n103 163.367
R655 B.n109 B.n108 163.367
R656 B.n113 B.n112 163.367
R657 B.n117 B.n116 163.367
R658 B.n121 B.n120 163.367
R659 B.n125 B.n124 163.367
R660 B.n130 B.n129 163.367
R661 B.n134 B.n133 163.367
R662 B.n138 B.n137 163.367
R663 B.n140 B.n83 163.367
R664 B.n231 B.t12 145.524
R665 B.n87 B.t9 145.524
R666 B.n234 B.t15 145.524
R667 B.n85 B.t19 145.524
R668 B.n293 B.n212 118.075
R669 B.n293 B.n208 118.075
R670 B.n299 B.n208 118.075
R671 B.n299 B.n204 118.075
R672 B.n306 B.n204 118.075
R673 B.n306 B.n305 118.075
R674 B.n312 B.n197 118.075
R675 B.n318 B.n197 118.075
R676 B.n318 B.n193 118.075
R677 B.n324 B.n193 118.075
R678 B.n324 B.n189 118.075
R679 B.n330 B.n189 118.075
R680 B.n330 B.n185 118.075
R681 B.n336 B.n185 118.075
R682 B.n336 B.n181 118.075
R683 B.n342 B.n181 118.075
R684 B.n348 B.n177 118.075
R685 B.n348 B.n173 118.075
R686 B.n354 B.n173 118.075
R687 B.n354 B.n168 118.075
R688 B.n360 B.n168 118.075
R689 B.n360 B.n169 118.075
R690 B.n366 B.n161 118.075
R691 B.n372 B.n161 118.075
R692 B.n372 B.n157 118.075
R693 B.n378 B.n157 118.075
R694 B.n378 B.n153 118.075
R695 B.n384 B.n153 118.075
R696 B.n391 B.n149 118.075
R697 B.n391 B.n145 118.075
R698 B.n397 B.n145 118.075
R699 B.n397 B.n4 118.075
R700 B.n525 B.n4 118.075
R701 B.n525 B.n524 118.075
R702 B.n524 B.n523 118.075
R703 B.n523 B.n8 118.075
R704 B.n517 B.n8 118.075
R705 B.n517 B.n516 118.075
R706 B.n515 B.n15 118.075
R707 B.n509 B.n15 118.075
R708 B.n509 B.n508 118.075
R709 B.n508 B.n507 118.075
R710 B.n507 B.n22 118.075
R711 B.n501 B.n22 118.075
R712 B.n500 B.n499 118.075
R713 B.n499 B.n29 118.075
R714 B.n493 B.n29 118.075
R715 B.n493 B.n492 118.075
R716 B.n492 B.n491 118.075
R717 B.n491 B.n36 118.075
R718 B.n485 B.n484 118.075
R719 B.n484 B.n483 118.075
R720 B.n483 B.n43 118.075
R721 B.n477 B.n43 118.075
R722 B.n477 B.n476 118.075
R723 B.n476 B.n475 118.075
R724 B.n475 B.n50 118.075
R725 B.n469 B.n50 118.075
R726 B.n469 B.n468 118.075
R727 B.n468 B.n467 118.075
R728 B.n461 B.n60 118.075
R729 B.n461 B.n460 118.075
R730 B.n460 B.n459 118.075
R731 B.n459 B.n64 118.075
R732 B.n453 B.n64 118.075
R733 B.n453 B.n452 118.075
R734 B.n305 B.t11 90.2925
R735 B.t4 B.n177 90.2925
R736 B.n384 B.t5 90.2925
R737 B.t2 B.n515 90.2925
R738 B.t0 B.n36 90.2925
R739 B.n60 B.t7 90.2925
R740 B.n286 B.n285 71.676
R741 B.n280 B.n216 71.676
R742 B.n277 B.n217 71.676
R743 B.n273 B.n218 71.676
R744 B.n269 B.n219 71.676
R745 B.n265 B.n220 71.676
R746 B.n261 B.n221 71.676
R747 B.n257 B.n222 71.676
R748 B.n253 B.n223 71.676
R749 B.n249 B.n224 71.676
R750 B.n245 B.n225 71.676
R751 B.n241 B.n226 71.676
R752 B.n237 B.n227 71.676
R753 B.n88 B.n70 71.676
R754 B.n92 B.n71 71.676
R755 B.n96 B.n72 71.676
R756 B.n100 B.n73 71.676
R757 B.n104 B.n74 71.676
R758 B.n109 B.n75 71.676
R759 B.n113 B.n76 71.676
R760 B.n117 B.n77 71.676
R761 B.n121 B.n78 71.676
R762 B.n125 B.n79 71.676
R763 B.n130 B.n80 71.676
R764 B.n134 B.n81 71.676
R765 B.n138 B.n82 71.676
R766 B.n450 B.n83 71.676
R767 B.n450 B.n449 71.676
R768 B.n140 B.n82 71.676
R769 B.n137 B.n81 71.676
R770 B.n133 B.n80 71.676
R771 B.n129 B.n79 71.676
R772 B.n124 B.n78 71.676
R773 B.n120 B.n77 71.676
R774 B.n116 B.n76 71.676
R775 B.n112 B.n75 71.676
R776 B.n108 B.n74 71.676
R777 B.n103 B.n73 71.676
R778 B.n99 B.n72 71.676
R779 B.n95 B.n71 71.676
R780 B.n91 B.n70 71.676
R781 B.n286 B.n229 71.676
R782 B.n278 B.n216 71.676
R783 B.n274 B.n217 71.676
R784 B.n270 B.n218 71.676
R785 B.n266 B.n219 71.676
R786 B.n262 B.n220 71.676
R787 B.n258 B.n221 71.676
R788 B.n254 B.n222 71.676
R789 B.n250 B.n223 71.676
R790 B.n246 B.n224 71.676
R791 B.n242 B.n225 71.676
R792 B.n238 B.n226 71.676
R793 B.n227 B.n215 71.676
R794 B.n235 B.n234 59.5399
R795 B.n232 B.n231 59.5399
R796 B.n106 B.n87 59.5399
R797 B.n127 B.n85 59.5399
R798 B.n169 B.t1 59.0376
R799 B.n366 B.t1 59.0376
R800 B.n501 B.t3 59.0376
R801 B.t3 B.n500 59.0376
R802 B.n234 B.n233 47.9035
R803 B.n231 B.n230 47.9035
R804 B.n87 B.n86 47.9035
R805 B.n85 B.n84 47.9035
R806 B.n89 B.n66 36.6834
R807 B.n448 B.n447 36.6834
R808 B.n290 B.n289 36.6834
R809 B.n284 B.n210 36.6834
R810 B.n312 B.t11 27.7827
R811 B.n342 B.t4 27.7827
R812 B.t5 B.n149 27.7827
R813 B.n516 B.t2 27.7827
R814 B.n485 B.t0 27.7827
R815 B.n467 B.t7 27.7827
R816 B B.n527 18.0485
R817 B.n90 B.n89 10.6151
R818 B.n93 B.n90 10.6151
R819 B.n94 B.n93 10.6151
R820 B.n97 B.n94 10.6151
R821 B.n98 B.n97 10.6151
R822 B.n101 B.n98 10.6151
R823 B.n102 B.n101 10.6151
R824 B.n105 B.n102 10.6151
R825 B.n110 B.n107 10.6151
R826 B.n111 B.n110 10.6151
R827 B.n114 B.n111 10.6151
R828 B.n115 B.n114 10.6151
R829 B.n118 B.n115 10.6151
R830 B.n119 B.n118 10.6151
R831 B.n122 B.n119 10.6151
R832 B.n123 B.n122 10.6151
R833 B.n126 B.n123 10.6151
R834 B.n131 B.n128 10.6151
R835 B.n132 B.n131 10.6151
R836 B.n135 B.n132 10.6151
R837 B.n136 B.n135 10.6151
R838 B.n139 B.n136 10.6151
R839 B.n141 B.n139 10.6151
R840 B.n142 B.n141 10.6151
R841 B.n448 B.n142 10.6151
R842 B.n291 B.n290 10.6151
R843 B.n291 B.n206 10.6151
R844 B.n301 B.n206 10.6151
R845 B.n302 B.n301 10.6151
R846 B.n303 B.n302 10.6151
R847 B.n303 B.n199 10.6151
R848 B.n314 B.n199 10.6151
R849 B.n315 B.n314 10.6151
R850 B.n316 B.n315 10.6151
R851 B.n316 B.n191 10.6151
R852 B.n326 B.n191 10.6151
R853 B.n327 B.n326 10.6151
R854 B.n328 B.n327 10.6151
R855 B.n328 B.n183 10.6151
R856 B.n338 B.n183 10.6151
R857 B.n339 B.n338 10.6151
R858 B.n340 B.n339 10.6151
R859 B.n340 B.n175 10.6151
R860 B.n350 B.n175 10.6151
R861 B.n351 B.n350 10.6151
R862 B.n352 B.n351 10.6151
R863 B.n352 B.n166 10.6151
R864 B.n362 B.n166 10.6151
R865 B.n363 B.n362 10.6151
R866 B.n364 B.n363 10.6151
R867 B.n364 B.n159 10.6151
R868 B.n374 B.n159 10.6151
R869 B.n375 B.n374 10.6151
R870 B.n376 B.n375 10.6151
R871 B.n376 B.n151 10.6151
R872 B.n386 B.n151 10.6151
R873 B.n387 B.n386 10.6151
R874 B.n389 B.n387 10.6151
R875 B.n389 B.n388 10.6151
R876 B.n388 B.n143 10.6151
R877 B.n400 B.n143 10.6151
R878 B.n401 B.n400 10.6151
R879 B.n402 B.n401 10.6151
R880 B.n403 B.n402 10.6151
R881 B.n405 B.n403 10.6151
R882 B.n406 B.n405 10.6151
R883 B.n407 B.n406 10.6151
R884 B.n408 B.n407 10.6151
R885 B.n410 B.n408 10.6151
R886 B.n411 B.n410 10.6151
R887 B.n412 B.n411 10.6151
R888 B.n413 B.n412 10.6151
R889 B.n415 B.n413 10.6151
R890 B.n416 B.n415 10.6151
R891 B.n417 B.n416 10.6151
R892 B.n418 B.n417 10.6151
R893 B.n420 B.n418 10.6151
R894 B.n421 B.n420 10.6151
R895 B.n422 B.n421 10.6151
R896 B.n423 B.n422 10.6151
R897 B.n425 B.n423 10.6151
R898 B.n426 B.n425 10.6151
R899 B.n427 B.n426 10.6151
R900 B.n428 B.n427 10.6151
R901 B.n430 B.n428 10.6151
R902 B.n431 B.n430 10.6151
R903 B.n432 B.n431 10.6151
R904 B.n433 B.n432 10.6151
R905 B.n435 B.n433 10.6151
R906 B.n436 B.n435 10.6151
R907 B.n437 B.n436 10.6151
R908 B.n438 B.n437 10.6151
R909 B.n440 B.n438 10.6151
R910 B.n441 B.n440 10.6151
R911 B.n442 B.n441 10.6151
R912 B.n443 B.n442 10.6151
R913 B.n445 B.n443 10.6151
R914 B.n446 B.n445 10.6151
R915 B.n447 B.n446 10.6151
R916 B.n284 B.n283 10.6151
R917 B.n283 B.n282 10.6151
R918 B.n282 B.n281 10.6151
R919 B.n281 B.n279 10.6151
R920 B.n279 B.n276 10.6151
R921 B.n276 B.n275 10.6151
R922 B.n275 B.n272 10.6151
R923 B.n272 B.n271 10.6151
R924 B.n268 B.n267 10.6151
R925 B.n267 B.n264 10.6151
R926 B.n264 B.n263 10.6151
R927 B.n263 B.n260 10.6151
R928 B.n260 B.n259 10.6151
R929 B.n259 B.n256 10.6151
R930 B.n256 B.n255 10.6151
R931 B.n255 B.n252 10.6151
R932 B.n252 B.n251 10.6151
R933 B.n248 B.n247 10.6151
R934 B.n247 B.n244 10.6151
R935 B.n244 B.n243 10.6151
R936 B.n243 B.n240 10.6151
R937 B.n240 B.n239 10.6151
R938 B.n239 B.n236 10.6151
R939 B.n236 B.n214 10.6151
R940 B.n289 B.n214 10.6151
R941 B.n295 B.n210 10.6151
R942 B.n296 B.n295 10.6151
R943 B.n297 B.n296 10.6151
R944 B.n297 B.n202 10.6151
R945 B.n308 B.n202 10.6151
R946 B.n309 B.n308 10.6151
R947 B.n310 B.n309 10.6151
R948 B.n310 B.n195 10.6151
R949 B.n320 B.n195 10.6151
R950 B.n321 B.n320 10.6151
R951 B.n322 B.n321 10.6151
R952 B.n322 B.n187 10.6151
R953 B.n332 B.n187 10.6151
R954 B.n333 B.n332 10.6151
R955 B.n334 B.n333 10.6151
R956 B.n334 B.n179 10.6151
R957 B.n344 B.n179 10.6151
R958 B.n345 B.n344 10.6151
R959 B.n346 B.n345 10.6151
R960 B.n346 B.n171 10.6151
R961 B.n356 B.n171 10.6151
R962 B.n357 B.n356 10.6151
R963 B.n358 B.n357 10.6151
R964 B.n358 B.n163 10.6151
R965 B.n368 B.n163 10.6151
R966 B.n369 B.n368 10.6151
R967 B.n370 B.n369 10.6151
R968 B.n370 B.n155 10.6151
R969 B.n380 B.n155 10.6151
R970 B.n381 B.n380 10.6151
R971 B.n382 B.n381 10.6151
R972 B.n382 B.n147 10.6151
R973 B.n393 B.n147 10.6151
R974 B.n394 B.n393 10.6151
R975 B.n395 B.n394 10.6151
R976 B.n395 B.n0 10.6151
R977 B.n521 B.n1 10.6151
R978 B.n521 B.n520 10.6151
R979 B.n520 B.n519 10.6151
R980 B.n519 B.n10 10.6151
R981 B.n513 B.n10 10.6151
R982 B.n513 B.n512 10.6151
R983 B.n512 B.n511 10.6151
R984 B.n511 B.n17 10.6151
R985 B.n505 B.n17 10.6151
R986 B.n505 B.n504 10.6151
R987 B.n504 B.n503 10.6151
R988 B.n503 B.n24 10.6151
R989 B.n497 B.n24 10.6151
R990 B.n497 B.n496 10.6151
R991 B.n496 B.n495 10.6151
R992 B.n495 B.n31 10.6151
R993 B.n489 B.n31 10.6151
R994 B.n489 B.n488 10.6151
R995 B.n488 B.n487 10.6151
R996 B.n487 B.n38 10.6151
R997 B.n481 B.n38 10.6151
R998 B.n481 B.n480 10.6151
R999 B.n480 B.n479 10.6151
R1000 B.n479 B.n45 10.6151
R1001 B.n473 B.n45 10.6151
R1002 B.n473 B.n472 10.6151
R1003 B.n472 B.n471 10.6151
R1004 B.n471 B.n52 10.6151
R1005 B.n465 B.n52 10.6151
R1006 B.n465 B.n464 10.6151
R1007 B.n464 B.n463 10.6151
R1008 B.n463 B.n58 10.6151
R1009 B.n457 B.n58 10.6151
R1010 B.n457 B.n456 10.6151
R1011 B.n456 B.n455 10.6151
R1012 B.n455 B.n66 10.6151
R1013 B.n106 B.n105 9.36635
R1014 B.n128 B.n127 9.36635
R1015 B.n271 B.n232 9.36635
R1016 B.n248 B.n235 9.36635
R1017 B.n527 B.n0 2.81026
R1018 B.n527 B.n1 2.81026
R1019 B.n107 B.n106 1.24928
R1020 B.n127 B.n126 1.24928
R1021 B.n268 B.n232 1.24928
R1022 B.n251 B.n235 1.24928
R1023 VN.n21 VN.n12 161.3
R1024 VN.n20 VN.n19 161.3
R1025 VN.n18 VN.n13 161.3
R1026 VN.n17 VN.n16 161.3
R1027 VN.n9 VN.n0 161.3
R1028 VN.n8 VN.n7 161.3
R1029 VN.n6 VN.n1 161.3
R1030 VN.n5 VN.n4 161.3
R1031 VN.n11 VN.n10 87.7234
R1032 VN.n23 VN.n22 87.7234
R1033 VN.n8 VN.n1 56.4773
R1034 VN.n20 VN.n13 56.4773
R1035 VN.n2 VN.t1 46.4527
R1036 VN.n14 VN.t4 46.4527
R1037 VN.n15 VN.n14 46.2445
R1038 VN.n3 VN.n2 46.2445
R1039 VN VN.n23 38.9716
R1040 VN.n4 VN.n3 24.3439
R1041 VN.n4 VN.n1 24.3439
R1042 VN.n9 VN.n8 24.3439
R1043 VN.n16 VN.n13 24.3439
R1044 VN.n16 VN.n15 24.3439
R1045 VN.n21 VN.n20 24.3439
R1046 VN.n10 VN.n9 22.8833
R1047 VN.n22 VN.n21 22.8833
R1048 VN.n3 VN.t2 11.9379
R1049 VN.n10 VN.t5 11.9379
R1050 VN.n15 VN.t0 11.9379
R1051 VN.n22 VN.t3 11.9379
R1052 VN.n17 VN.n14 8.71313
R1053 VN.n5 VN.n2 8.71313
R1054 VN.n23 VN.n12 0.278398
R1055 VN.n11 VN.n0 0.278398
R1056 VN.n19 VN.n12 0.189894
R1057 VN.n19 VN.n18 0.189894
R1058 VN.n18 VN.n17 0.189894
R1059 VN.n6 VN.n5 0.189894
R1060 VN.n7 VN.n6 0.189894
R1061 VN.n7 VN.n0 0.189894
R1062 VN VN.n11 0.153422
R1063 VDD2.n1 VDD2.t4 173.167
R1064 VDD2.n2 VDD2.t2 171.625
R1065 VDD2.n1 VDD2.n0 145.94
R1066 VDD2 VDD2.n3 145.936
R1067 VDD2.n2 VDD2.n1 31.5493
R1068 VDD2.n3 VDD2.t5 18.6797
R1069 VDD2.n3 VDD2.t1 18.6797
R1070 VDD2.n0 VDD2.t3 18.6797
R1071 VDD2.n0 VDD2.t0 18.6797
R1072 VDD2 VDD2.n2 1.65567
C0 VDD2 VP 0.427313f
C1 VDD2 VDD1 1.22695f
C2 VDD2 VTAIL 3.47011f
C3 VDD1 VP 1.1828f
C4 VTAIL VP 1.74118f
C5 VDD2 VN 0.915939f
C6 VTAIL VDD1 3.41988f
C7 VN VP 4.46446f
C8 VDD1 VN 0.1576f
C9 VTAIL VN 1.72705f
C10 VDD2 B 3.554005f
C11 VDD1 B 3.808528f
C12 VTAIL B 2.694323f
C13 VN B 10.157605f
C14 VP B 9.124391f
C15 VDD2.t4 B 0.106203f
C16 VDD2.t3 B 0.015389f
C17 VDD2.t0 B 0.015389f
C18 VDD2.n0 B 0.079716f
C19 VDD2.n1 B 1.41635f
C20 VDD2.t2 B 0.104156f
C21 VDD2.n2 B 1.25127f
C22 VDD2.t5 B 0.015389f
C23 VDD2.t1 B 0.015389f
C24 VDD2.n3 B 0.079707f
C25 VN.n0 B 0.031779f
C26 VN.t5 B 0.105041f
C27 VN.n1 B 0.034324f
C28 VN.t1 B 0.260423f
C29 VN.n2 B 0.119947f
C30 VN.t2 B 0.105041f
C31 VN.n3 B 0.147186f
C32 VN.n4 B 0.045147f
C33 VN.n5 B 0.203344f
C34 VN.n6 B 0.024103f
C35 VN.n7 B 0.024103f
C36 VN.n8 B 0.036353f
C37 VN.n9 B 0.043809f
C38 VN.n10 B 0.157822f
C39 VN.n11 B 0.027216f
C40 VN.n12 B 0.031779f
C41 VN.t3 B 0.105041f
C42 VN.n13 B 0.034324f
C43 VN.t4 B 0.260423f
C44 VN.n14 B 0.119947f
C45 VN.t0 B 0.105041f
C46 VN.n15 B 0.147186f
C47 VN.n16 B 0.045147f
C48 VN.n17 B 0.203344f
C49 VN.n18 B 0.024103f
C50 VN.n19 B 0.024103f
C51 VN.n20 B 0.036353f
C52 VN.n21 B 0.043809f
C53 VN.n22 B 0.157822f
C54 VN.n23 B 0.897022f
C55 VDD1.t3 B 0.101407f
C56 VDD1.t5 B 0.101207f
C57 VDD1.t0 B 0.014665f
C58 VDD1.t1 B 0.014665f
C59 VDD1.n0 B 0.075966f
C60 VDD1.n1 B 1.42064f
C61 VDD1.t2 B 0.014665f
C62 VDD1.t4 B 0.014665f
C63 VDD1.n2 B 0.075103f
C64 VDD1.n3 B 1.2238f
C65 VTAIL.t2 B 0.021325f
C66 VTAIL.t3 B 0.021325f
C67 VTAIL.n0 B 0.089315f
C68 VTAIL.n1 B 0.318092f
C69 VTAIL.t7 B 0.125316f
C70 VTAIL.n2 B 0.466481f
C71 VTAIL.t11 B 0.021325f
C72 VTAIL.t9 B 0.021325f
C73 VTAIL.n3 B 0.089315f
C74 VTAIL.n4 B 1.08857f
C75 VTAIL.t4 B 0.021325f
C76 VTAIL.t1 B 0.021325f
C77 VTAIL.n5 B 0.089315f
C78 VTAIL.n6 B 1.08857f
C79 VTAIL.t5 B 0.125316f
C80 VTAIL.n7 B 0.466481f
C81 VTAIL.t8 B 0.021325f
C82 VTAIL.t6 B 0.021325f
C83 VTAIL.n8 B 0.089315f
C84 VTAIL.n9 B 0.444323f
C85 VTAIL.t10 B 0.125316f
C86 VTAIL.n10 B 0.936059f
C87 VTAIL.t0 B 0.125316f
C88 VTAIL.n11 B 0.887617f
C89 VP.n0 B 0.03202f
C90 VP.t4 B 0.105838f
C91 VP.n1 B 0.034585f
C92 VP.n2 B 0.024286f
C93 VP.t5 B 0.105838f
C94 VP.n3 B 0.034585f
C95 VP.n4 B 0.03202f
C96 VP.t0 B 0.105838f
C97 VP.n5 B 0.03202f
C98 VP.t1 B 0.105838f
C99 VP.n6 B 0.034585f
C100 VP.t2 B 0.262399f
C101 VP.n7 B 0.120857f
C102 VP.t3 B 0.105838f
C103 VP.n8 B 0.148303f
C104 VP.n9 B 0.045489f
C105 VP.n10 B 0.204887f
C106 VP.n11 B 0.024286f
C107 VP.n12 B 0.024286f
C108 VP.n13 B 0.036629f
C109 VP.n14 B 0.044142f
C110 VP.n15 B 0.15902f
C111 VP.n16 B 0.890174f
C112 VP.n17 B 0.912672f
C113 VP.n18 B 0.15902f
C114 VP.n19 B 0.044142f
C115 VP.n20 B 0.036629f
C116 VP.n21 B 0.024286f
C117 VP.n22 B 0.024286f
C118 VP.n23 B 0.024286f
C119 VP.n24 B 0.045489f
C120 VP.n25 B 0.096952f
C121 VP.n26 B 0.045489f
C122 VP.n27 B 0.024286f
C123 VP.n28 B 0.024286f
C124 VP.n29 B 0.024286f
C125 VP.n30 B 0.036629f
C126 VP.n31 B 0.044142f
C127 VP.n32 B 0.15902f
C128 VP.n33 B 0.027423f
.ends

