* NGSPICE file created from diff_pair_sample_1026.ext - technology: sky130A

.subckt diff_pair_sample_1026 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=5.46 pd=28.78 as=0 ps=0 w=14 l=2.17
X1 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=5.46 pd=28.78 as=0 ps=0 w=14 l=2.17
X2 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.46 pd=28.78 as=0 ps=0 w=14 l=2.17
X3 VDD1.t1 VP.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=5.46 pd=28.78 as=5.46 ps=28.78 w=14 l=2.17
X4 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.46 pd=28.78 as=5.46 ps=28.78 w=14 l=2.17
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=5.46 pd=28.78 as=0 ps=0 w=14 l=2.17
X6 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.46 pd=28.78 as=5.46 ps=28.78 w=14 l=2.17
X7 VDD1.t0 VP.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=5.46 pd=28.78 as=5.46 ps=28.78 w=14 l=2.17
R0 B.n720 B.n719 585
R1 B.n721 B.n720 585
R2 B.n308 B.n98 585
R3 B.n307 B.n306 585
R4 B.n305 B.n304 585
R5 B.n303 B.n302 585
R6 B.n301 B.n300 585
R7 B.n299 B.n298 585
R8 B.n297 B.n296 585
R9 B.n295 B.n294 585
R10 B.n293 B.n292 585
R11 B.n291 B.n290 585
R12 B.n289 B.n288 585
R13 B.n287 B.n286 585
R14 B.n285 B.n284 585
R15 B.n283 B.n282 585
R16 B.n281 B.n280 585
R17 B.n279 B.n278 585
R18 B.n277 B.n276 585
R19 B.n275 B.n274 585
R20 B.n273 B.n272 585
R21 B.n271 B.n270 585
R22 B.n269 B.n268 585
R23 B.n267 B.n266 585
R24 B.n265 B.n264 585
R25 B.n263 B.n262 585
R26 B.n261 B.n260 585
R27 B.n259 B.n258 585
R28 B.n257 B.n256 585
R29 B.n255 B.n254 585
R30 B.n253 B.n252 585
R31 B.n251 B.n250 585
R32 B.n249 B.n248 585
R33 B.n247 B.n246 585
R34 B.n245 B.n244 585
R35 B.n243 B.n242 585
R36 B.n241 B.n240 585
R37 B.n239 B.n238 585
R38 B.n237 B.n236 585
R39 B.n235 B.n234 585
R40 B.n233 B.n232 585
R41 B.n231 B.n230 585
R42 B.n229 B.n228 585
R43 B.n227 B.n226 585
R44 B.n225 B.n224 585
R45 B.n223 B.n222 585
R46 B.n221 B.n220 585
R47 B.n219 B.n218 585
R48 B.n217 B.n216 585
R49 B.n214 B.n213 585
R50 B.n212 B.n211 585
R51 B.n210 B.n209 585
R52 B.n208 B.n207 585
R53 B.n206 B.n205 585
R54 B.n204 B.n203 585
R55 B.n202 B.n201 585
R56 B.n200 B.n199 585
R57 B.n198 B.n197 585
R58 B.n196 B.n195 585
R59 B.n194 B.n193 585
R60 B.n192 B.n191 585
R61 B.n190 B.n189 585
R62 B.n188 B.n187 585
R63 B.n186 B.n185 585
R64 B.n184 B.n183 585
R65 B.n182 B.n181 585
R66 B.n180 B.n179 585
R67 B.n178 B.n177 585
R68 B.n176 B.n175 585
R69 B.n174 B.n173 585
R70 B.n172 B.n171 585
R71 B.n170 B.n169 585
R72 B.n168 B.n167 585
R73 B.n166 B.n165 585
R74 B.n164 B.n163 585
R75 B.n162 B.n161 585
R76 B.n160 B.n159 585
R77 B.n158 B.n157 585
R78 B.n156 B.n155 585
R79 B.n154 B.n153 585
R80 B.n152 B.n151 585
R81 B.n150 B.n149 585
R82 B.n148 B.n147 585
R83 B.n146 B.n145 585
R84 B.n144 B.n143 585
R85 B.n142 B.n141 585
R86 B.n140 B.n139 585
R87 B.n138 B.n137 585
R88 B.n136 B.n135 585
R89 B.n134 B.n133 585
R90 B.n132 B.n131 585
R91 B.n130 B.n129 585
R92 B.n128 B.n127 585
R93 B.n126 B.n125 585
R94 B.n124 B.n123 585
R95 B.n122 B.n121 585
R96 B.n120 B.n119 585
R97 B.n118 B.n117 585
R98 B.n116 B.n115 585
R99 B.n114 B.n113 585
R100 B.n112 B.n111 585
R101 B.n110 B.n109 585
R102 B.n108 B.n107 585
R103 B.n106 B.n105 585
R104 B.n46 B.n45 585
R105 B.n724 B.n723 585
R106 B.n718 B.n99 585
R107 B.n99 B.n43 585
R108 B.n717 B.n42 585
R109 B.n728 B.n42 585
R110 B.n716 B.n41 585
R111 B.n729 B.n41 585
R112 B.n715 B.n40 585
R113 B.n730 B.n40 585
R114 B.n714 B.n713 585
R115 B.n713 B.n36 585
R116 B.n712 B.n35 585
R117 B.n736 B.n35 585
R118 B.n711 B.n34 585
R119 B.n737 B.n34 585
R120 B.n710 B.n33 585
R121 B.n738 B.n33 585
R122 B.n709 B.n708 585
R123 B.n708 B.n29 585
R124 B.n707 B.n28 585
R125 B.n744 B.n28 585
R126 B.n706 B.n27 585
R127 B.n745 B.n27 585
R128 B.n705 B.n26 585
R129 B.n746 B.n26 585
R130 B.n704 B.n703 585
R131 B.n703 B.n22 585
R132 B.n702 B.n21 585
R133 B.n752 B.n21 585
R134 B.n701 B.n20 585
R135 B.n753 B.n20 585
R136 B.n700 B.n19 585
R137 B.n754 B.n19 585
R138 B.n699 B.n698 585
R139 B.n698 B.n15 585
R140 B.n697 B.n14 585
R141 B.n760 B.n14 585
R142 B.n696 B.n13 585
R143 B.n761 B.n13 585
R144 B.n695 B.n12 585
R145 B.n762 B.n12 585
R146 B.n694 B.n693 585
R147 B.n693 B.n8 585
R148 B.n692 B.n7 585
R149 B.n768 B.n7 585
R150 B.n691 B.n6 585
R151 B.n769 B.n6 585
R152 B.n690 B.n5 585
R153 B.n770 B.n5 585
R154 B.n689 B.n688 585
R155 B.n688 B.n4 585
R156 B.n687 B.n309 585
R157 B.n687 B.n686 585
R158 B.n677 B.n310 585
R159 B.n311 B.n310 585
R160 B.n679 B.n678 585
R161 B.n680 B.n679 585
R162 B.n676 B.n316 585
R163 B.n316 B.n315 585
R164 B.n675 B.n674 585
R165 B.n674 B.n673 585
R166 B.n318 B.n317 585
R167 B.n319 B.n318 585
R168 B.n666 B.n665 585
R169 B.n667 B.n666 585
R170 B.n664 B.n324 585
R171 B.n324 B.n323 585
R172 B.n663 B.n662 585
R173 B.n662 B.n661 585
R174 B.n326 B.n325 585
R175 B.n327 B.n326 585
R176 B.n654 B.n653 585
R177 B.n655 B.n654 585
R178 B.n652 B.n332 585
R179 B.n332 B.n331 585
R180 B.n651 B.n650 585
R181 B.n650 B.n649 585
R182 B.n334 B.n333 585
R183 B.n335 B.n334 585
R184 B.n642 B.n641 585
R185 B.n643 B.n642 585
R186 B.n640 B.n340 585
R187 B.n340 B.n339 585
R188 B.n639 B.n638 585
R189 B.n638 B.n637 585
R190 B.n342 B.n341 585
R191 B.n343 B.n342 585
R192 B.n630 B.n629 585
R193 B.n631 B.n630 585
R194 B.n628 B.n348 585
R195 B.n348 B.n347 585
R196 B.n627 B.n626 585
R197 B.n626 B.n625 585
R198 B.n350 B.n349 585
R199 B.n351 B.n350 585
R200 B.n621 B.n620 585
R201 B.n354 B.n353 585
R202 B.n617 B.n616 585
R203 B.n618 B.n617 585
R204 B.n615 B.n406 585
R205 B.n614 B.n613 585
R206 B.n612 B.n611 585
R207 B.n610 B.n609 585
R208 B.n608 B.n607 585
R209 B.n606 B.n605 585
R210 B.n604 B.n603 585
R211 B.n602 B.n601 585
R212 B.n600 B.n599 585
R213 B.n598 B.n597 585
R214 B.n596 B.n595 585
R215 B.n594 B.n593 585
R216 B.n592 B.n591 585
R217 B.n590 B.n589 585
R218 B.n588 B.n587 585
R219 B.n586 B.n585 585
R220 B.n584 B.n583 585
R221 B.n582 B.n581 585
R222 B.n580 B.n579 585
R223 B.n578 B.n577 585
R224 B.n576 B.n575 585
R225 B.n574 B.n573 585
R226 B.n572 B.n571 585
R227 B.n570 B.n569 585
R228 B.n568 B.n567 585
R229 B.n566 B.n565 585
R230 B.n564 B.n563 585
R231 B.n562 B.n561 585
R232 B.n560 B.n559 585
R233 B.n558 B.n557 585
R234 B.n556 B.n555 585
R235 B.n554 B.n553 585
R236 B.n552 B.n551 585
R237 B.n550 B.n549 585
R238 B.n548 B.n547 585
R239 B.n546 B.n545 585
R240 B.n544 B.n543 585
R241 B.n542 B.n541 585
R242 B.n540 B.n539 585
R243 B.n538 B.n537 585
R244 B.n536 B.n535 585
R245 B.n534 B.n533 585
R246 B.n532 B.n531 585
R247 B.n530 B.n529 585
R248 B.n528 B.n527 585
R249 B.n525 B.n524 585
R250 B.n523 B.n522 585
R251 B.n521 B.n520 585
R252 B.n519 B.n518 585
R253 B.n517 B.n516 585
R254 B.n515 B.n514 585
R255 B.n513 B.n512 585
R256 B.n511 B.n510 585
R257 B.n509 B.n508 585
R258 B.n507 B.n506 585
R259 B.n505 B.n504 585
R260 B.n503 B.n502 585
R261 B.n501 B.n500 585
R262 B.n499 B.n498 585
R263 B.n497 B.n496 585
R264 B.n495 B.n494 585
R265 B.n493 B.n492 585
R266 B.n491 B.n490 585
R267 B.n489 B.n488 585
R268 B.n487 B.n486 585
R269 B.n485 B.n484 585
R270 B.n483 B.n482 585
R271 B.n481 B.n480 585
R272 B.n479 B.n478 585
R273 B.n477 B.n476 585
R274 B.n475 B.n474 585
R275 B.n473 B.n472 585
R276 B.n471 B.n470 585
R277 B.n469 B.n468 585
R278 B.n467 B.n466 585
R279 B.n465 B.n464 585
R280 B.n463 B.n462 585
R281 B.n461 B.n460 585
R282 B.n459 B.n458 585
R283 B.n457 B.n456 585
R284 B.n455 B.n454 585
R285 B.n453 B.n452 585
R286 B.n451 B.n450 585
R287 B.n449 B.n448 585
R288 B.n447 B.n446 585
R289 B.n445 B.n444 585
R290 B.n443 B.n442 585
R291 B.n441 B.n440 585
R292 B.n439 B.n438 585
R293 B.n437 B.n436 585
R294 B.n435 B.n434 585
R295 B.n433 B.n432 585
R296 B.n431 B.n430 585
R297 B.n429 B.n428 585
R298 B.n427 B.n426 585
R299 B.n425 B.n424 585
R300 B.n423 B.n422 585
R301 B.n421 B.n420 585
R302 B.n419 B.n418 585
R303 B.n417 B.n416 585
R304 B.n415 B.n414 585
R305 B.n413 B.n412 585
R306 B.n622 B.n352 585
R307 B.n352 B.n351 585
R308 B.n624 B.n623 585
R309 B.n625 B.n624 585
R310 B.n346 B.n345 585
R311 B.n347 B.n346 585
R312 B.n633 B.n632 585
R313 B.n632 B.n631 585
R314 B.n634 B.n344 585
R315 B.n344 B.n343 585
R316 B.n636 B.n635 585
R317 B.n637 B.n636 585
R318 B.n338 B.n337 585
R319 B.n339 B.n338 585
R320 B.n645 B.n644 585
R321 B.n644 B.n643 585
R322 B.n646 B.n336 585
R323 B.n336 B.n335 585
R324 B.n648 B.n647 585
R325 B.n649 B.n648 585
R326 B.n330 B.n329 585
R327 B.n331 B.n330 585
R328 B.n657 B.n656 585
R329 B.n656 B.n655 585
R330 B.n658 B.n328 585
R331 B.n328 B.n327 585
R332 B.n660 B.n659 585
R333 B.n661 B.n660 585
R334 B.n322 B.n321 585
R335 B.n323 B.n322 585
R336 B.n669 B.n668 585
R337 B.n668 B.n667 585
R338 B.n670 B.n320 585
R339 B.n320 B.n319 585
R340 B.n672 B.n671 585
R341 B.n673 B.n672 585
R342 B.n314 B.n313 585
R343 B.n315 B.n314 585
R344 B.n682 B.n681 585
R345 B.n681 B.n680 585
R346 B.n683 B.n312 585
R347 B.n312 B.n311 585
R348 B.n685 B.n684 585
R349 B.n686 B.n685 585
R350 B.n2 B.n0 585
R351 B.n4 B.n2 585
R352 B.n3 B.n1 585
R353 B.n769 B.n3 585
R354 B.n767 B.n766 585
R355 B.n768 B.n767 585
R356 B.n765 B.n9 585
R357 B.n9 B.n8 585
R358 B.n764 B.n763 585
R359 B.n763 B.n762 585
R360 B.n11 B.n10 585
R361 B.n761 B.n11 585
R362 B.n759 B.n758 585
R363 B.n760 B.n759 585
R364 B.n757 B.n16 585
R365 B.n16 B.n15 585
R366 B.n756 B.n755 585
R367 B.n755 B.n754 585
R368 B.n18 B.n17 585
R369 B.n753 B.n18 585
R370 B.n751 B.n750 585
R371 B.n752 B.n751 585
R372 B.n749 B.n23 585
R373 B.n23 B.n22 585
R374 B.n748 B.n747 585
R375 B.n747 B.n746 585
R376 B.n25 B.n24 585
R377 B.n745 B.n25 585
R378 B.n743 B.n742 585
R379 B.n744 B.n743 585
R380 B.n741 B.n30 585
R381 B.n30 B.n29 585
R382 B.n740 B.n739 585
R383 B.n739 B.n738 585
R384 B.n32 B.n31 585
R385 B.n737 B.n32 585
R386 B.n735 B.n734 585
R387 B.n736 B.n735 585
R388 B.n733 B.n37 585
R389 B.n37 B.n36 585
R390 B.n732 B.n731 585
R391 B.n731 B.n730 585
R392 B.n39 B.n38 585
R393 B.n729 B.n39 585
R394 B.n727 B.n726 585
R395 B.n728 B.n727 585
R396 B.n725 B.n44 585
R397 B.n44 B.n43 585
R398 B.n772 B.n771 585
R399 B.n771 B.n770 585
R400 B.n620 B.n352 434.841
R401 B.n723 B.n44 434.841
R402 B.n412 B.n350 434.841
R403 B.n720 B.n99 434.841
R404 B.n409 B.t12 364.854
R405 B.n100 B.t14 364.854
R406 B.n407 B.t5 364.854
R407 B.n102 B.t8 364.854
R408 B.n409 B.t10 362.774
R409 B.n407 B.t2 362.774
R410 B.n102 B.t6 362.774
R411 B.n100 B.t13 362.774
R412 B.n410 B.t11 316.37
R413 B.n101 B.t15 316.37
R414 B.n408 B.t4 316.37
R415 B.n103 B.t9 316.37
R416 B.n721 B.n97 256.663
R417 B.n721 B.n96 256.663
R418 B.n721 B.n95 256.663
R419 B.n721 B.n94 256.663
R420 B.n721 B.n93 256.663
R421 B.n721 B.n92 256.663
R422 B.n721 B.n91 256.663
R423 B.n721 B.n90 256.663
R424 B.n721 B.n89 256.663
R425 B.n721 B.n88 256.663
R426 B.n721 B.n87 256.663
R427 B.n721 B.n86 256.663
R428 B.n721 B.n85 256.663
R429 B.n721 B.n84 256.663
R430 B.n721 B.n83 256.663
R431 B.n721 B.n82 256.663
R432 B.n721 B.n81 256.663
R433 B.n721 B.n80 256.663
R434 B.n721 B.n79 256.663
R435 B.n721 B.n78 256.663
R436 B.n721 B.n77 256.663
R437 B.n721 B.n76 256.663
R438 B.n721 B.n75 256.663
R439 B.n721 B.n74 256.663
R440 B.n721 B.n73 256.663
R441 B.n721 B.n72 256.663
R442 B.n721 B.n71 256.663
R443 B.n721 B.n70 256.663
R444 B.n721 B.n69 256.663
R445 B.n721 B.n68 256.663
R446 B.n721 B.n67 256.663
R447 B.n721 B.n66 256.663
R448 B.n721 B.n65 256.663
R449 B.n721 B.n64 256.663
R450 B.n721 B.n63 256.663
R451 B.n721 B.n62 256.663
R452 B.n721 B.n61 256.663
R453 B.n721 B.n60 256.663
R454 B.n721 B.n59 256.663
R455 B.n721 B.n58 256.663
R456 B.n721 B.n57 256.663
R457 B.n721 B.n56 256.663
R458 B.n721 B.n55 256.663
R459 B.n721 B.n54 256.663
R460 B.n721 B.n53 256.663
R461 B.n721 B.n52 256.663
R462 B.n721 B.n51 256.663
R463 B.n721 B.n50 256.663
R464 B.n721 B.n49 256.663
R465 B.n721 B.n48 256.663
R466 B.n721 B.n47 256.663
R467 B.n722 B.n721 256.663
R468 B.n619 B.n618 256.663
R469 B.n618 B.n355 256.663
R470 B.n618 B.n356 256.663
R471 B.n618 B.n357 256.663
R472 B.n618 B.n358 256.663
R473 B.n618 B.n359 256.663
R474 B.n618 B.n360 256.663
R475 B.n618 B.n361 256.663
R476 B.n618 B.n362 256.663
R477 B.n618 B.n363 256.663
R478 B.n618 B.n364 256.663
R479 B.n618 B.n365 256.663
R480 B.n618 B.n366 256.663
R481 B.n618 B.n367 256.663
R482 B.n618 B.n368 256.663
R483 B.n618 B.n369 256.663
R484 B.n618 B.n370 256.663
R485 B.n618 B.n371 256.663
R486 B.n618 B.n372 256.663
R487 B.n618 B.n373 256.663
R488 B.n618 B.n374 256.663
R489 B.n618 B.n375 256.663
R490 B.n618 B.n376 256.663
R491 B.n618 B.n377 256.663
R492 B.n618 B.n378 256.663
R493 B.n618 B.n379 256.663
R494 B.n618 B.n380 256.663
R495 B.n618 B.n381 256.663
R496 B.n618 B.n382 256.663
R497 B.n618 B.n383 256.663
R498 B.n618 B.n384 256.663
R499 B.n618 B.n385 256.663
R500 B.n618 B.n386 256.663
R501 B.n618 B.n387 256.663
R502 B.n618 B.n388 256.663
R503 B.n618 B.n389 256.663
R504 B.n618 B.n390 256.663
R505 B.n618 B.n391 256.663
R506 B.n618 B.n392 256.663
R507 B.n618 B.n393 256.663
R508 B.n618 B.n394 256.663
R509 B.n618 B.n395 256.663
R510 B.n618 B.n396 256.663
R511 B.n618 B.n397 256.663
R512 B.n618 B.n398 256.663
R513 B.n618 B.n399 256.663
R514 B.n618 B.n400 256.663
R515 B.n618 B.n401 256.663
R516 B.n618 B.n402 256.663
R517 B.n618 B.n403 256.663
R518 B.n618 B.n404 256.663
R519 B.n618 B.n405 256.663
R520 B.n624 B.n352 163.367
R521 B.n624 B.n346 163.367
R522 B.n632 B.n346 163.367
R523 B.n632 B.n344 163.367
R524 B.n636 B.n344 163.367
R525 B.n636 B.n338 163.367
R526 B.n644 B.n338 163.367
R527 B.n644 B.n336 163.367
R528 B.n648 B.n336 163.367
R529 B.n648 B.n330 163.367
R530 B.n656 B.n330 163.367
R531 B.n656 B.n328 163.367
R532 B.n660 B.n328 163.367
R533 B.n660 B.n322 163.367
R534 B.n668 B.n322 163.367
R535 B.n668 B.n320 163.367
R536 B.n672 B.n320 163.367
R537 B.n672 B.n314 163.367
R538 B.n681 B.n314 163.367
R539 B.n681 B.n312 163.367
R540 B.n685 B.n312 163.367
R541 B.n685 B.n2 163.367
R542 B.n771 B.n2 163.367
R543 B.n771 B.n3 163.367
R544 B.n767 B.n3 163.367
R545 B.n767 B.n9 163.367
R546 B.n763 B.n9 163.367
R547 B.n763 B.n11 163.367
R548 B.n759 B.n11 163.367
R549 B.n759 B.n16 163.367
R550 B.n755 B.n16 163.367
R551 B.n755 B.n18 163.367
R552 B.n751 B.n18 163.367
R553 B.n751 B.n23 163.367
R554 B.n747 B.n23 163.367
R555 B.n747 B.n25 163.367
R556 B.n743 B.n25 163.367
R557 B.n743 B.n30 163.367
R558 B.n739 B.n30 163.367
R559 B.n739 B.n32 163.367
R560 B.n735 B.n32 163.367
R561 B.n735 B.n37 163.367
R562 B.n731 B.n37 163.367
R563 B.n731 B.n39 163.367
R564 B.n727 B.n39 163.367
R565 B.n727 B.n44 163.367
R566 B.n617 B.n354 163.367
R567 B.n617 B.n406 163.367
R568 B.n613 B.n612 163.367
R569 B.n609 B.n608 163.367
R570 B.n605 B.n604 163.367
R571 B.n601 B.n600 163.367
R572 B.n597 B.n596 163.367
R573 B.n593 B.n592 163.367
R574 B.n589 B.n588 163.367
R575 B.n585 B.n584 163.367
R576 B.n581 B.n580 163.367
R577 B.n577 B.n576 163.367
R578 B.n573 B.n572 163.367
R579 B.n569 B.n568 163.367
R580 B.n565 B.n564 163.367
R581 B.n561 B.n560 163.367
R582 B.n557 B.n556 163.367
R583 B.n553 B.n552 163.367
R584 B.n549 B.n548 163.367
R585 B.n545 B.n544 163.367
R586 B.n541 B.n540 163.367
R587 B.n537 B.n536 163.367
R588 B.n533 B.n532 163.367
R589 B.n529 B.n528 163.367
R590 B.n524 B.n523 163.367
R591 B.n520 B.n519 163.367
R592 B.n516 B.n515 163.367
R593 B.n512 B.n511 163.367
R594 B.n508 B.n507 163.367
R595 B.n504 B.n503 163.367
R596 B.n500 B.n499 163.367
R597 B.n496 B.n495 163.367
R598 B.n492 B.n491 163.367
R599 B.n488 B.n487 163.367
R600 B.n484 B.n483 163.367
R601 B.n480 B.n479 163.367
R602 B.n476 B.n475 163.367
R603 B.n472 B.n471 163.367
R604 B.n468 B.n467 163.367
R605 B.n464 B.n463 163.367
R606 B.n460 B.n459 163.367
R607 B.n456 B.n455 163.367
R608 B.n452 B.n451 163.367
R609 B.n448 B.n447 163.367
R610 B.n444 B.n443 163.367
R611 B.n440 B.n439 163.367
R612 B.n436 B.n435 163.367
R613 B.n432 B.n431 163.367
R614 B.n428 B.n427 163.367
R615 B.n424 B.n423 163.367
R616 B.n420 B.n419 163.367
R617 B.n416 B.n415 163.367
R618 B.n626 B.n350 163.367
R619 B.n626 B.n348 163.367
R620 B.n630 B.n348 163.367
R621 B.n630 B.n342 163.367
R622 B.n638 B.n342 163.367
R623 B.n638 B.n340 163.367
R624 B.n642 B.n340 163.367
R625 B.n642 B.n334 163.367
R626 B.n650 B.n334 163.367
R627 B.n650 B.n332 163.367
R628 B.n654 B.n332 163.367
R629 B.n654 B.n326 163.367
R630 B.n662 B.n326 163.367
R631 B.n662 B.n324 163.367
R632 B.n666 B.n324 163.367
R633 B.n666 B.n318 163.367
R634 B.n674 B.n318 163.367
R635 B.n674 B.n316 163.367
R636 B.n679 B.n316 163.367
R637 B.n679 B.n310 163.367
R638 B.n687 B.n310 163.367
R639 B.n688 B.n687 163.367
R640 B.n688 B.n5 163.367
R641 B.n6 B.n5 163.367
R642 B.n7 B.n6 163.367
R643 B.n693 B.n7 163.367
R644 B.n693 B.n12 163.367
R645 B.n13 B.n12 163.367
R646 B.n14 B.n13 163.367
R647 B.n698 B.n14 163.367
R648 B.n698 B.n19 163.367
R649 B.n20 B.n19 163.367
R650 B.n21 B.n20 163.367
R651 B.n703 B.n21 163.367
R652 B.n703 B.n26 163.367
R653 B.n27 B.n26 163.367
R654 B.n28 B.n27 163.367
R655 B.n708 B.n28 163.367
R656 B.n708 B.n33 163.367
R657 B.n34 B.n33 163.367
R658 B.n35 B.n34 163.367
R659 B.n713 B.n35 163.367
R660 B.n713 B.n40 163.367
R661 B.n41 B.n40 163.367
R662 B.n42 B.n41 163.367
R663 B.n99 B.n42 163.367
R664 B.n105 B.n46 163.367
R665 B.n109 B.n108 163.367
R666 B.n113 B.n112 163.367
R667 B.n117 B.n116 163.367
R668 B.n121 B.n120 163.367
R669 B.n125 B.n124 163.367
R670 B.n129 B.n128 163.367
R671 B.n133 B.n132 163.367
R672 B.n137 B.n136 163.367
R673 B.n141 B.n140 163.367
R674 B.n145 B.n144 163.367
R675 B.n149 B.n148 163.367
R676 B.n153 B.n152 163.367
R677 B.n157 B.n156 163.367
R678 B.n161 B.n160 163.367
R679 B.n165 B.n164 163.367
R680 B.n169 B.n168 163.367
R681 B.n173 B.n172 163.367
R682 B.n177 B.n176 163.367
R683 B.n181 B.n180 163.367
R684 B.n185 B.n184 163.367
R685 B.n189 B.n188 163.367
R686 B.n193 B.n192 163.367
R687 B.n197 B.n196 163.367
R688 B.n201 B.n200 163.367
R689 B.n205 B.n204 163.367
R690 B.n209 B.n208 163.367
R691 B.n213 B.n212 163.367
R692 B.n218 B.n217 163.367
R693 B.n222 B.n221 163.367
R694 B.n226 B.n225 163.367
R695 B.n230 B.n229 163.367
R696 B.n234 B.n233 163.367
R697 B.n238 B.n237 163.367
R698 B.n242 B.n241 163.367
R699 B.n246 B.n245 163.367
R700 B.n250 B.n249 163.367
R701 B.n254 B.n253 163.367
R702 B.n258 B.n257 163.367
R703 B.n262 B.n261 163.367
R704 B.n266 B.n265 163.367
R705 B.n270 B.n269 163.367
R706 B.n274 B.n273 163.367
R707 B.n278 B.n277 163.367
R708 B.n282 B.n281 163.367
R709 B.n286 B.n285 163.367
R710 B.n290 B.n289 163.367
R711 B.n294 B.n293 163.367
R712 B.n298 B.n297 163.367
R713 B.n302 B.n301 163.367
R714 B.n306 B.n305 163.367
R715 B.n720 B.n98 163.367
R716 B.n620 B.n619 71.676
R717 B.n406 B.n355 71.676
R718 B.n612 B.n356 71.676
R719 B.n608 B.n357 71.676
R720 B.n604 B.n358 71.676
R721 B.n600 B.n359 71.676
R722 B.n596 B.n360 71.676
R723 B.n592 B.n361 71.676
R724 B.n588 B.n362 71.676
R725 B.n584 B.n363 71.676
R726 B.n580 B.n364 71.676
R727 B.n576 B.n365 71.676
R728 B.n572 B.n366 71.676
R729 B.n568 B.n367 71.676
R730 B.n564 B.n368 71.676
R731 B.n560 B.n369 71.676
R732 B.n556 B.n370 71.676
R733 B.n552 B.n371 71.676
R734 B.n548 B.n372 71.676
R735 B.n544 B.n373 71.676
R736 B.n540 B.n374 71.676
R737 B.n536 B.n375 71.676
R738 B.n532 B.n376 71.676
R739 B.n528 B.n377 71.676
R740 B.n523 B.n378 71.676
R741 B.n519 B.n379 71.676
R742 B.n515 B.n380 71.676
R743 B.n511 B.n381 71.676
R744 B.n507 B.n382 71.676
R745 B.n503 B.n383 71.676
R746 B.n499 B.n384 71.676
R747 B.n495 B.n385 71.676
R748 B.n491 B.n386 71.676
R749 B.n487 B.n387 71.676
R750 B.n483 B.n388 71.676
R751 B.n479 B.n389 71.676
R752 B.n475 B.n390 71.676
R753 B.n471 B.n391 71.676
R754 B.n467 B.n392 71.676
R755 B.n463 B.n393 71.676
R756 B.n459 B.n394 71.676
R757 B.n455 B.n395 71.676
R758 B.n451 B.n396 71.676
R759 B.n447 B.n397 71.676
R760 B.n443 B.n398 71.676
R761 B.n439 B.n399 71.676
R762 B.n435 B.n400 71.676
R763 B.n431 B.n401 71.676
R764 B.n427 B.n402 71.676
R765 B.n423 B.n403 71.676
R766 B.n419 B.n404 71.676
R767 B.n415 B.n405 71.676
R768 B.n723 B.n722 71.676
R769 B.n105 B.n47 71.676
R770 B.n109 B.n48 71.676
R771 B.n113 B.n49 71.676
R772 B.n117 B.n50 71.676
R773 B.n121 B.n51 71.676
R774 B.n125 B.n52 71.676
R775 B.n129 B.n53 71.676
R776 B.n133 B.n54 71.676
R777 B.n137 B.n55 71.676
R778 B.n141 B.n56 71.676
R779 B.n145 B.n57 71.676
R780 B.n149 B.n58 71.676
R781 B.n153 B.n59 71.676
R782 B.n157 B.n60 71.676
R783 B.n161 B.n61 71.676
R784 B.n165 B.n62 71.676
R785 B.n169 B.n63 71.676
R786 B.n173 B.n64 71.676
R787 B.n177 B.n65 71.676
R788 B.n181 B.n66 71.676
R789 B.n185 B.n67 71.676
R790 B.n189 B.n68 71.676
R791 B.n193 B.n69 71.676
R792 B.n197 B.n70 71.676
R793 B.n201 B.n71 71.676
R794 B.n205 B.n72 71.676
R795 B.n209 B.n73 71.676
R796 B.n213 B.n74 71.676
R797 B.n218 B.n75 71.676
R798 B.n222 B.n76 71.676
R799 B.n226 B.n77 71.676
R800 B.n230 B.n78 71.676
R801 B.n234 B.n79 71.676
R802 B.n238 B.n80 71.676
R803 B.n242 B.n81 71.676
R804 B.n246 B.n82 71.676
R805 B.n250 B.n83 71.676
R806 B.n254 B.n84 71.676
R807 B.n258 B.n85 71.676
R808 B.n262 B.n86 71.676
R809 B.n266 B.n87 71.676
R810 B.n270 B.n88 71.676
R811 B.n274 B.n89 71.676
R812 B.n278 B.n90 71.676
R813 B.n282 B.n91 71.676
R814 B.n286 B.n92 71.676
R815 B.n290 B.n93 71.676
R816 B.n294 B.n94 71.676
R817 B.n298 B.n95 71.676
R818 B.n302 B.n96 71.676
R819 B.n306 B.n97 71.676
R820 B.n98 B.n97 71.676
R821 B.n305 B.n96 71.676
R822 B.n301 B.n95 71.676
R823 B.n297 B.n94 71.676
R824 B.n293 B.n93 71.676
R825 B.n289 B.n92 71.676
R826 B.n285 B.n91 71.676
R827 B.n281 B.n90 71.676
R828 B.n277 B.n89 71.676
R829 B.n273 B.n88 71.676
R830 B.n269 B.n87 71.676
R831 B.n265 B.n86 71.676
R832 B.n261 B.n85 71.676
R833 B.n257 B.n84 71.676
R834 B.n253 B.n83 71.676
R835 B.n249 B.n82 71.676
R836 B.n245 B.n81 71.676
R837 B.n241 B.n80 71.676
R838 B.n237 B.n79 71.676
R839 B.n233 B.n78 71.676
R840 B.n229 B.n77 71.676
R841 B.n225 B.n76 71.676
R842 B.n221 B.n75 71.676
R843 B.n217 B.n74 71.676
R844 B.n212 B.n73 71.676
R845 B.n208 B.n72 71.676
R846 B.n204 B.n71 71.676
R847 B.n200 B.n70 71.676
R848 B.n196 B.n69 71.676
R849 B.n192 B.n68 71.676
R850 B.n188 B.n67 71.676
R851 B.n184 B.n66 71.676
R852 B.n180 B.n65 71.676
R853 B.n176 B.n64 71.676
R854 B.n172 B.n63 71.676
R855 B.n168 B.n62 71.676
R856 B.n164 B.n61 71.676
R857 B.n160 B.n60 71.676
R858 B.n156 B.n59 71.676
R859 B.n152 B.n58 71.676
R860 B.n148 B.n57 71.676
R861 B.n144 B.n56 71.676
R862 B.n140 B.n55 71.676
R863 B.n136 B.n54 71.676
R864 B.n132 B.n53 71.676
R865 B.n128 B.n52 71.676
R866 B.n124 B.n51 71.676
R867 B.n120 B.n50 71.676
R868 B.n116 B.n49 71.676
R869 B.n112 B.n48 71.676
R870 B.n108 B.n47 71.676
R871 B.n722 B.n46 71.676
R872 B.n619 B.n354 71.676
R873 B.n613 B.n355 71.676
R874 B.n609 B.n356 71.676
R875 B.n605 B.n357 71.676
R876 B.n601 B.n358 71.676
R877 B.n597 B.n359 71.676
R878 B.n593 B.n360 71.676
R879 B.n589 B.n361 71.676
R880 B.n585 B.n362 71.676
R881 B.n581 B.n363 71.676
R882 B.n577 B.n364 71.676
R883 B.n573 B.n365 71.676
R884 B.n569 B.n366 71.676
R885 B.n565 B.n367 71.676
R886 B.n561 B.n368 71.676
R887 B.n557 B.n369 71.676
R888 B.n553 B.n370 71.676
R889 B.n549 B.n371 71.676
R890 B.n545 B.n372 71.676
R891 B.n541 B.n373 71.676
R892 B.n537 B.n374 71.676
R893 B.n533 B.n375 71.676
R894 B.n529 B.n376 71.676
R895 B.n524 B.n377 71.676
R896 B.n520 B.n378 71.676
R897 B.n516 B.n379 71.676
R898 B.n512 B.n380 71.676
R899 B.n508 B.n381 71.676
R900 B.n504 B.n382 71.676
R901 B.n500 B.n383 71.676
R902 B.n496 B.n384 71.676
R903 B.n492 B.n385 71.676
R904 B.n488 B.n386 71.676
R905 B.n484 B.n387 71.676
R906 B.n480 B.n388 71.676
R907 B.n476 B.n389 71.676
R908 B.n472 B.n390 71.676
R909 B.n468 B.n391 71.676
R910 B.n464 B.n392 71.676
R911 B.n460 B.n393 71.676
R912 B.n456 B.n394 71.676
R913 B.n452 B.n395 71.676
R914 B.n448 B.n396 71.676
R915 B.n444 B.n397 71.676
R916 B.n440 B.n398 71.676
R917 B.n436 B.n399 71.676
R918 B.n432 B.n400 71.676
R919 B.n428 B.n401 71.676
R920 B.n424 B.n402 71.676
R921 B.n420 B.n403 71.676
R922 B.n416 B.n404 71.676
R923 B.n412 B.n405 71.676
R924 B.n618 B.n351 63.3468
R925 B.n721 B.n43 63.3468
R926 B.n411 B.n410 59.5399
R927 B.n526 B.n408 59.5399
R928 B.n104 B.n103 59.5399
R929 B.n215 B.n101 59.5399
R930 B.n410 B.n409 48.4853
R931 B.n408 B.n407 48.4853
R932 B.n103 B.n102 48.4853
R933 B.n101 B.n100 48.4853
R934 B.n625 B.n351 38.8072
R935 B.n625 B.n347 38.8072
R936 B.n631 B.n347 38.8072
R937 B.n631 B.n343 38.8072
R938 B.n637 B.n343 38.8072
R939 B.n637 B.n339 38.8072
R940 B.n643 B.n339 38.8072
R941 B.n649 B.n335 38.8072
R942 B.n649 B.n331 38.8072
R943 B.n655 B.n331 38.8072
R944 B.n655 B.n327 38.8072
R945 B.n661 B.n327 38.8072
R946 B.n661 B.n323 38.8072
R947 B.n667 B.n323 38.8072
R948 B.n667 B.n319 38.8072
R949 B.n673 B.n319 38.8072
R950 B.n680 B.n315 38.8072
R951 B.n680 B.n311 38.8072
R952 B.n686 B.n311 38.8072
R953 B.n686 B.n4 38.8072
R954 B.n770 B.n4 38.8072
R955 B.n770 B.n769 38.8072
R956 B.n769 B.n768 38.8072
R957 B.n768 B.n8 38.8072
R958 B.n762 B.n8 38.8072
R959 B.n762 B.n761 38.8072
R960 B.n760 B.n15 38.8072
R961 B.n754 B.n15 38.8072
R962 B.n754 B.n753 38.8072
R963 B.n753 B.n752 38.8072
R964 B.n752 B.n22 38.8072
R965 B.n746 B.n22 38.8072
R966 B.n746 B.n745 38.8072
R967 B.n745 B.n744 38.8072
R968 B.n744 B.n29 38.8072
R969 B.n738 B.n737 38.8072
R970 B.n737 B.n736 38.8072
R971 B.n736 B.n36 38.8072
R972 B.n730 B.n36 38.8072
R973 B.n730 B.n729 38.8072
R974 B.n729 B.n728 38.8072
R975 B.n728 B.n43 38.8072
R976 B.t3 B.n335 32.5297
R977 B.t7 B.n29 32.5297
R978 B.n725 B.n724 28.2542
R979 B.n719 B.n718 28.2542
R980 B.n413 B.n349 28.2542
R981 B.n622 B.n621 28.2542
R982 B.n673 B.t0 27.9642
R983 B.t1 B.n760 27.9642
R984 B B.n772 18.0485
R985 B.t0 B.n315 10.8436
R986 B.n761 B.t1 10.8436
R987 B.n724 B.n45 10.6151
R988 B.n106 B.n45 10.6151
R989 B.n107 B.n106 10.6151
R990 B.n110 B.n107 10.6151
R991 B.n111 B.n110 10.6151
R992 B.n114 B.n111 10.6151
R993 B.n115 B.n114 10.6151
R994 B.n118 B.n115 10.6151
R995 B.n119 B.n118 10.6151
R996 B.n122 B.n119 10.6151
R997 B.n123 B.n122 10.6151
R998 B.n126 B.n123 10.6151
R999 B.n127 B.n126 10.6151
R1000 B.n130 B.n127 10.6151
R1001 B.n131 B.n130 10.6151
R1002 B.n134 B.n131 10.6151
R1003 B.n135 B.n134 10.6151
R1004 B.n138 B.n135 10.6151
R1005 B.n139 B.n138 10.6151
R1006 B.n142 B.n139 10.6151
R1007 B.n143 B.n142 10.6151
R1008 B.n146 B.n143 10.6151
R1009 B.n147 B.n146 10.6151
R1010 B.n150 B.n147 10.6151
R1011 B.n151 B.n150 10.6151
R1012 B.n154 B.n151 10.6151
R1013 B.n155 B.n154 10.6151
R1014 B.n158 B.n155 10.6151
R1015 B.n159 B.n158 10.6151
R1016 B.n162 B.n159 10.6151
R1017 B.n163 B.n162 10.6151
R1018 B.n166 B.n163 10.6151
R1019 B.n167 B.n166 10.6151
R1020 B.n170 B.n167 10.6151
R1021 B.n171 B.n170 10.6151
R1022 B.n174 B.n171 10.6151
R1023 B.n175 B.n174 10.6151
R1024 B.n178 B.n175 10.6151
R1025 B.n179 B.n178 10.6151
R1026 B.n182 B.n179 10.6151
R1027 B.n183 B.n182 10.6151
R1028 B.n186 B.n183 10.6151
R1029 B.n187 B.n186 10.6151
R1030 B.n190 B.n187 10.6151
R1031 B.n191 B.n190 10.6151
R1032 B.n194 B.n191 10.6151
R1033 B.n195 B.n194 10.6151
R1034 B.n199 B.n198 10.6151
R1035 B.n202 B.n199 10.6151
R1036 B.n203 B.n202 10.6151
R1037 B.n206 B.n203 10.6151
R1038 B.n207 B.n206 10.6151
R1039 B.n210 B.n207 10.6151
R1040 B.n211 B.n210 10.6151
R1041 B.n214 B.n211 10.6151
R1042 B.n219 B.n216 10.6151
R1043 B.n220 B.n219 10.6151
R1044 B.n223 B.n220 10.6151
R1045 B.n224 B.n223 10.6151
R1046 B.n227 B.n224 10.6151
R1047 B.n228 B.n227 10.6151
R1048 B.n231 B.n228 10.6151
R1049 B.n232 B.n231 10.6151
R1050 B.n235 B.n232 10.6151
R1051 B.n236 B.n235 10.6151
R1052 B.n239 B.n236 10.6151
R1053 B.n240 B.n239 10.6151
R1054 B.n243 B.n240 10.6151
R1055 B.n244 B.n243 10.6151
R1056 B.n247 B.n244 10.6151
R1057 B.n248 B.n247 10.6151
R1058 B.n251 B.n248 10.6151
R1059 B.n252 B.n251 10.6151
R1060 B.n255 B.n252 10.6151
R1061 B.n256 B.n255 10.6151
R1062 B.n259 B.n256 10.6151
R1063 B.n260 B.n259 10.6151
R1064 B.n263 B.n260 10.6151
R1065 B.n264 B.n263 10.6151
R1066 B.n267 B.n264 10.6151
R1067 B.n268 B.n267 10.6151
R1068 B.n271 B.n268 10.6151
R1069 B.n272 B.n271 10.6151
R1070 B.n275 B.n272 10.6151
R1071 B.n276 B.n275 10.6151
R1072 B.n279 B.n276 10.6151
R1073 B.n280 B.n279 10.6151
R1074 B.n283 B.n280 10.6151
R1075 B.n284 B.n283 10.6151
R1076 B.n287 B.n284 10.6151
R1077 B.n288 B.n287 10.6151
R1078 B.n291 B.n288 10.6151
R1079 B.n292 B.n291 10.6151
R1080 B.n295 B.n292 10.6151
R1081 B.n296 B.n295 10.6151
R1082 B.n299 B.n296 10.6151
R1083 B.n300 B.n299 10.6151
R1084 B.n303 B.n300 10.6151
R1085 B.n304 B.n303 10.6151
R1086 B.n307 B.n304 10.6151
R1087 B.n308 B.n307 10.6151
R1088 B.n719 B.n308 10.6151
R1089 B.n627 B.n349 10.6151
R1090 B.n628 B.n627 10.6151
R1091 B.n629 B.n628 10.6151
R1092 B.n629 B.n341 10.6151
R1093 B.n639 B.n341 10.6151
R1094 B.n640 B.n639 10.6151
R1095 B.n641 B.n640 10.6151
R1096 B.n641 B.n333 10.6151
R1097 B.n651 B.n333 10.6151
R1098 B.n652 B.n651 10.6151
R1099 B.n653 B.n652 10.6151
R1100 B.n653 B.n325 10.6151
R1101 B.n663 B.n325 10.6151
R1102 B.n664 B.n663 10.6151
R1103 B.n665 B.n664 10.6151
R1104 B.n665 B.n317 10.6151
R1105 B.n675 B.n317 10.6151
R1106 B.n676 B.n675 10.6151
R1107 B.n678 B.n676 10.6151
R1108 B.n678 B.n677 10.6151
R1109 B.n677 B.n309 10.6151
R1110 B.n689 B.n309 10.6151
R1111 B.n690 B.n689 10.6151
R1112 B.n691 B.n690 10.6151
R1113 B.n692 B.n691 10.6151
R1114 B.n694 B.n692 10.6151
R1115 B.n695 B.n694 10.6151
R1116 B.n696 B.n695 10.6151
R1117 B.n697 B.n696 10.6151
R1118 B.n699 B.n697 10.6151
R1119 B.n700 B.n699 10.6151
R1120 B.n701 B.n700 10.6151
R1121 B.n702 B.n701 10.6151
R1122 B.n704 B.n702 10.6151
R1123 B.n705 B.n704 10.6151
R1124 B.n706 B.n705 10.6151
R1125 B.n707 B.n706 10.6151
R1126 B.n709 B.n707 10.6151
R1127 B.n710 B.n709 10.6151
R1128 B.n711 B.n710 10.6151
R1129 B.n712 B.n711 10.6151
R1130 B.n714 B.n712 10.6151
R1131 B.n715 B.n714 10.6151
R1132 B.n716 B.n715 10.6151
R1133 B.n717 B.n716 10.6151
R1134 B.n718 B.n717 10.6151
R1135 B.n621 B.n353 10.6151
R1136 B.n616 B.n353 10.6151
R1137 B.n616 B.n615 10.6151
R1138 B.n615 B.n614 10.6151
R1139 B.n614 B.n611 10.6151
R1140 B.n611 B.n610 10.6151
R1141 B.n610 B.n607 10.6151
R1142 B.n607 B.n606 10.6151
R1143 B.n606 B.n603 10.6151
R1144 B.n603 B.n602 10.6151
R1145 B.n602 B.n599 10.6151
R1146 B.n599 B.n598 10.6151
R1147 B.n598 B.n595 10.6151
R1148 B.n595 B.n594 10.6151
R1149 B.n594 B.n591 10.6151
R1150 B.n591 B.n590 10.6151
R1151 B.n590 B.n587 10.6151
R1152 B.n587 B.n586 10.6151
R1153 B.n586 B.n583 10.6151
R1154 B.n583 B.n582 10.6151
R1155 B.n582 B.n579 10.6151
R1156 B.n579 B.n578 10.6151
R1157 B.n578 B.n575 10.6151
R1158 B.n575 B.n574 10.6151
R1159 B.n574 B.n571 10.6151
R1160 B.n571 B.n570 10.6151
R1161 B.n570 B.n567 10.6151
R1162 B.n567 B.n566 10.6151
R1163 B.n566 B.n563 10.6151
R1164 B.n563 B.n562 10.6151
R1165 B.n562 B.n559 10.6151
R1166 B.n559 B.n558 10.6151
R1167 B.n558 B.n555 10.6151
R1168 B.n555 B.n554 10.6151
R1169 B.n554 B.n551 10.6151
R1170 B.n551 B.n550 10.6151
R1171 B.n550 B.n547 10.6151
R1172 B.n547 B.n546 10.6151
R1173 B.n546 B.n543 10.6151
R1174 B.n543 B.n542 10.6151
R1175 B.n542 B.n539 10.6151
R1176 B.n539 B.n538 10.6151
R1177 B.n538 B.n535 10.6151
R1178 B.n535 B.n534 10.6151
R1179 B.n534 B.n531 10.6151
R1180 B.n531 B.n530 10.6151
R1181 B.n530 B.n527 10.6151
R1182 B.n525 B.n522 10.6151
R1183 B.n522 B.n521 10.6151
R1184 B.n521 B.n518 10.6151
R1185 B.n518 B.n517 10.6151
R1186 B.n517 B.n514 10.6151
R1187 B.n514 B.n513 10.6151
R1188 B.n513 B.n510 10.6151
R1189 B.n510 B.n509 10.6151
R1190 B.n506 B.n505 10.6151
R1191 B.n505 B.n502 10.6151
R1192 B.n502 B.n501 10.6151
R1193 B.n501 B.n498 10.6151
R1194 B.n498 B.n497 10.6151
R1195 B.n497 B.n494 10.6151
R1196 B.n494 B.n493 10.6151
R1197 B.n493 B.n490 10.6151
R1198 B.n490 B.n489 10.6151
R1199 B.n489 B.n486 10.6151
R1200 B.n486 B.n485 10.6151
R1201 B.n485 B.n482 10.6151
R1202 B.n482 B.n481 10.6151
R1203 B.n481 B.n478 10.6151
R1204 B.n478 B.n477 10.6151
R1205 B.n477 B.n474 10.6151
R1206 B.n474 B.n473 10.6151
R1207 B.n473 B.n470 10.6151
R1208 B.n470 B.n469 10.6151
R1209 B.n469 B.n466 10.6151
R1210 B.n466 B.n465 10.6151
R1211 B.n465 B.n462 10.6151
R1212 B.n462 B.n461 10.6151
R1213 B.n461 B.n458 10.6151
R1214 B.n458 B.n457 10.6151
R1215 B.n457 B.n454 10.6151
R1216 B.n454 B.n453 10.6151
R1217 B.n453 B.n450 10.6151
R1218 B.n450 B.n449 10.6151
R1219 B.n449 B.n446 10.6151
R1220 B.n446 B.n445 10.6151
R1221 B.n445 B.n442 10.6151
R1222 B.n442 B.n441 10.6151
R1223 B.n441 B.n438 10.6151
R1224 B.n438 B.n437 10.6151
R1225 B.n437 B.n434 10.6151
R1226 B.n434 B.n433 10.6151
R1227 B.n433 B.n430 10.6151
R1228 B.n430 B.n429 10.6151
R1229 B.n429 B.n426 10.6151
R1230 B.n426 B.n425 10.6151
R1231 B.n425 B.n422 10.6151
R1232 B.n422 B.n421 10.6151
R1233 B.n421 B.n418 10.6151
R1234 B.n418 B.n417 10.6151
R1235 B.n417 B.n414 10.6151
R1236 B.n414 B.n413 10.6151
R1237 B.n623 B.n622 10.6151
R1238 B.n623 B.n345 10.6151
R1239 B.n633 B.n345 10.6151
R1240 B.n634 B.n633 10.6151
R1241 B.n635 B.n634 10.6151
R1242 B.n635 B.n337 10.6151
R1243 B.n645 B.n337 10.6151
R1244 B.n646 B.n645 10.6151
R1245 B.n647 B.n646 10.6151
R1246 B.n647 B.n329 10.6151
R1247 B.n657 B.n329 10.6151
R1248 B.n658 B.n657 10.6151
R1249 B.n659 B.n658 10.6151
R1250 B.n659 B.n321 10.6151
R1251 B.n669 B.n321 10.6151
R1252 B.n670 B.n669 10.6151
R1253 B.n671 B.n670 10.6151
R1254 B.n671 B.n313 10.6151
R1255 B.n682 B.n313 10.6151
R1256 B.n683 B.n682 10.6151
R1257 B.n684 B.n683 10.6151
R1258 B.n684 B.n0 10.6151
R1259 B.n766 B.n1 10.6151
R1260 B.n766 B.n765 10.6151
R1261 B.n765 B.n764 10.6151
R1262 B.n764 B.n10 10.6151
R1263 B.n758 B.n10 10.6151
R1264 B.n758 B.n757 10.6151
R1265 B.n757 B.n756 10.6151
R1266 B.n756 B.n17 10.6151
R1267 B.n750 B.n17 10.6151
R1268 B.n750 B.n749 10.6151
R1269 B.n749 B.n748 10.6151
R1270 B.n748 B.n24 10.6151
R1271 B.n742 B.n24 10.6151
R1272 B.n742 B.n741 10.6151
R1273 B.n741 B.n740 10.6151
R1274 B.n740 B.n31 10.6151
R1275 B.n734 B.n31 10.6151
R1276 B.n734 B.n733 10.6151
R1277 B.n733 B.n732 10.6151
R1278 B.n732 B.n38 10.6151
R1279 B.n726 B.n38 10.6151
R1280 B.n726 B.n725 10.6151
R1281 B.n198 B.n104 6.5566
R1282 B.n215 B.n214 6.5566
R1283 B.n526 B.n525 6.5566
R1284 B.n509 B.n411 6.5566
R1285 B.n643 B.t3 6.27806
R1286 B.n738 B.t7 6.27806
R1287 B.n195 B.n104 4.05904
R1288 B.n216 B.n215 4.05904
R1289 B.n527 B.n526 4.05904
R1290 B.n506 B.n411 4.05904
R1291 B.n772 B.n0 2.81026
R1292 B.n772 B.n1 2.81026
R1293 VP.n0 VP.t0 249.731
R1294 VP.n0 VP.t1 204.7
R1295 VP VP.n0 0.336784
R1296 VTAIL.n306 VTAIL.n234 289.615
R1297 VTAIL.n72 VTAIL.n0 289.615
R1298 VTAIL.n228 VTAIL.n156 289.615
R1299 VTAIL.n150 VTAIL.n78 289.615
R1300 VTAIL.n258 VTAIL.n257 185
R1301 VTAIL.n263 VTAIL.n262 185
R1302 VTAIL.n265 VTAIL.n264 185
R1303 VTAIL.n254 VTAIL.n253 185
R1304 VTAIL.n271 VTAIL.n270 185
R1305 VTAIL.n273 VTAIL.n272 185
R1306 VTAIL.n250 VTAIL.n249 185
R1307 VTAIL.n279 VTAIL.n278 185
R1308 VTAIL.n281 VTAIL.n280 185
R1309 VTAIL.n246 VTAIL.n245 185
R1310 VTAIL.n287 VTAIL.n286 185
R1311 VTAIL.n289 VTAIL.n288 185
R1312 VTAIL.n242 VTAIL.n241 185
R1313 VTAIL.n295 VTAIL.n294 185
R1314 VTAIL.n297 VTAIL.n296 185
R1315 VTAIL.n238 VTAIL.n237 185
R1316 VTAIL.n304 VTAIL.n303 185
R1317 VTAIL.n305 VTAIL.n236 185
R1318 VTAIL.n307 VTAIL.n306 185
R1319 VTAIL.n24 VTAIL.n23 185
R1320 VTAIL.n29 VTAIL.n28 185
R1321 VTAIL.n31 VTAIL.n30 185
R1322 VTAIL.n20 VTAIL.n19 185
R1323 VTAIL.n37 VTAIL.n36 185
R1324 VTAIL.n39 VTAIL.n38 185
R1325 VTAIL.n16 VTAIL.n15 185
R1326 VTAIL.n45 VTAIL.n44 185
R1327 VTAIL.n47 VTAIL.n46 185
R1328 VTAIL.n12 VTAIL.n11 185
R1329 VTAIL.n53 VTAIL.n52 185
R1330 VTAIL.n55 VTAIL.n54 185
R1331 VTAIL.n8 VTAIL.n7 185
R1332 VTAIL.n61 VTAIL.n60 185
R1333 VTAIL.n63 VTAIL.n62 185
R1334 VTAIL.n4 VTAIL.n3 185
R1335 VTAIL.n70 VTAIL.n69 185
R1336 VTAIL.n71 VTAIL.n2 185
R1337 VTAIL.n73 VTAIL.n72 185
R1338 VTAIL.n229 VTAIL.n228 185
R1339 VTAIL.n227 VTAIL.n158 185
R1340 VTAIL.n226 VTAIL.n225 185
R1341 VTAIL.n161 VTAIL.n159 185
R1342 VTAIL.n220 VTAIL.n219 185
R1343 VTAIL.n218 VTAIL.n217 185
R1344 VTAIL.n165 VTAIL.n164 185
R1345 VTAIL.n212 VTAIL.n211 185
R1346 VTAIL.n210 VTAIL.n209 185
R1347 VTAIL.n169 VTAIL.n168 185
R1348 VTAIL.n204 VTAIL.n203 185
R1349 VTAIL.n202 VTAIL.n201 185
R1350 VTAIL.n173 VTAIL.n172 185
R1351 VTAIL.n196 VTAIL.n195 185
R1352 VTAIL.n194 VTAIL.n193 185
R1353 VTAIL.n177 VTAIL.n176 185
R1354 VTAIL.n188 VTAIL.n187 185
R1355 VTAIL.n186 VTAIL.n185 185
R1356 VTAIL.n181 VTAIL.n180 185
R1357 VTAIL.n151 VTAIL.n150 185
R1358 VTAIL.n149 VTAIL.n80 185
R1359 VTAIL.n148 VTAIL.n147 185
R1360 VTAIL.n83 VTAIL.n81 185
R1361 VTAIL.n142 VTAIL.n141 185
R1362 VTAIL.n140 VTAIL.n139 185
R1363 VTAIL.n87 VTAIL.n86 185
R1364 VTAIL.n134 VTAIL.n133 185
R1365 VTAIL.n132 VTAIL.n131 185
R1366 VTAIL.n91 VTAIL.n90 185
R1367 VTAIL.n126 VTAIL.n125 185
R1368 VTAIL.n124 VTAIL.n123 185
R1369 VTAIL.n95 VTAIL.n94 185
R1370 VTAIL.n118 VTAIL.n117 185
R1371 VTAIL.n116 VTAIL.n115 185
R1372 VTAIL.n99 VTAIL.n98 185
R1373 VTAIL.n110 VTAIL.n109 185
R1374 VTAIL.n108 VTAIL.n107 185
R1375 VTAIL.n103 VTAIL.n102 185
R1376 VTAIL.n259 VTAIL.t1 147.659
R1377 VTAIL.n25 VTAIL.t3 147.659
R1378 VTAIL.n182 VTAIL.t2 147.659
R1379 VTAIL.n104 VTAIL.t0 147.659
R1380 VTAIL.n263 VTAIL.n257 104.615
R1381 VTAIL.n264 VTAIL.n263 104.615
R1382 VTAIL.n264 VTAIL.n253 104.615
R1383 VTAIL.n271 VTAIL.n253 104.615
R1384 VTAIL.n272 VTAIL.n271 104.615
R1385 VTAIL.n272 VTAIL.n249 104.615
R1386 VTAIL.n279 VTAIL.n249 104.615
R1387 VTAIL.n280 VTAIL.n279 104.615
R1388 VTAIL.n280 VTAIL.n245 104.615
R1389 VTAIL.n287 VTAIL.n245 104.615
R1390 VTAIL.n288 VTAIL.n287 104.615
R1391 VTAIL.n288 VTAIL.n241 104.615
R1392 VTAIL.n295 VTAIL.n241 104.615
R1393 VTAIL.n296 VTAIL.n295 104.615
R1394 VTAIL.n296 VTAIL.n237 104.615
R1395 VTAIL.n304 VTAIL.n237 104.615
R1396 VTAIL.n305 VTAIL.n304 104.615
R1397 VTAIL.n306 VTAIL.n305 104.615
R1398 VTAIL.n29 VTAIL.n23 104.615
R1399 VTAIL.n30 VTAIL.n29 104.615
R1400 VTAIL.n30 VTAIL.n19 104.615
R1401 VTAIL.n37 VTAIL.n19 104.615
R1402 VTAIL.n38 VTAIL.n37 104.615
R1403 VTAIL.n38 VTAIL.n15 104.615
R1404 VTAIL.n45 VTAIL.n15 104.615
R1405 VTAIL.n46 VTAIL.n45 104.615
R1406 VTAIL.n46 VTAIL.n11 104.615
R1407 VTAIL.n53 VTAIL.n11 104.615
R1408 VTAIL.n54 VTAIL.n53 104.615
R1409 VTAIL.n54 VTAIL.n7 104.615
R1410 VTAIL.n61 VTAIL.n7 104.615
R1411 VTAIL.n62 VTAIL.n61 104.615
R1412 VTAIL.n62 VTAIL.n3 104.615
R1413 VTAIL.n70 VTAIL.n3 104.615
R1414 VTAIL.n71 VTAIL.n70 104.615
R1415 VTAIL.n72 VTAIL.n71 104.615
R1416 VTAIL.n228 VTAIL.n227 104.615
R1417 VTAIL.n227 VTAIL.n226 104.615
R1418 VTAIL.n226 VTAIL.n159 104.615
R1419 VTAIL.n219 VTAIL.n159 104.615
R1420 VTAIL.n219 VTAIL.n218 104.615
R1421 VTAIL.n218 VTAIL.n164 104.615
R1422 VTAIL.n211 VTAIL.n164 104.615
R1423 VTAIL.n211 VTAIL.n210 104.615
R1424 VTAIL.n210 VTAIL.n168 104.615
R1425 VTAIL.n203 VTAIL.n168 104.615
R1426 VTAIL.n203 VTAIL.n202 104.615
R1427 VTAIL.n202 VTAIL.n172 104.615
R1428 VTAIL.n195 VTAIL.n172 104.615
R1429 VTAIL.n195 VTAIL.n194 104.615
R1430 VTAIL.n194 VTAIL.n176 104.615
R1431 VTAIL.n187 VTAIL.n176 104.615
R1432 VTAIL.n187 VTAIL.n186 104.615
R1433 VTAIL.n186 VTAIL.n180 104.615
R1434 VTAIL.n150 VTAIL.n149 104.615
R1435 VTAIL.n149 VTAIL.n148 104.615
R1436 VTAIL.n148 VTAIL.n81 104.615
R1437 VTAIL.n141 VTAIL.n81 104.615
R1438 VTAIL.n141 VTAIL.n140 104.615
R1439 VTAIL.n140 VTAIL.n86 104.615
R1440 VTAIL.n133 VTAIL.n86 104.615
R1441 VTAIL.n133 VTAIL.n132 104.615
R1442 VTAIL.n132 VTAIL.n90 104.615
R1443 VTAIL.n125 VTAIL.n90 104.615
R1444 VTAIL.n125 VTAIL.n124 104.615
R1445 VTAIL.n124 VTAIL.n94 104.615
R1446 VTAIL.n117 VTAIL.n94 104.615
R1447 VTAIL.n117 VTAIL.n116 104.615
R1448 VTAIL.n116 VTAIL.n98 104.615
R1449 VTAIL.n109 VTAIL.n98 104.615
R1450 VTAIL.n109 VTAIL.n108 104.615
R1451 VTAIL.n108 VTAIL.n102 104.615
R1452 VTAIL.t1 VTAIL.n257 52.3082
R1453 VTAIL.t3 VTAIL.n23 52.3082
R1454 VTAIL.t2 VTAIL.n180 52.3082
R1455 VTAIL.t0 VTAIL.n102 52.3082
R1456 VTAIL.n311 VTAIL.n310 33.7369
R1457 VTAIL.n77 VTAIL.n76 33.7369
R1458 VTAIL.n233 VTAIL.n232 33.7369
R1459 VTAIL.n155 VTAIL.n154 33.7369
R1460 VTAIL.n155 VTAIL.n77 28.7462
R1461 VTAIL.n311 VTAIL.n233 26.591
R1462 VTAIL.n259 VTAIL.n258 15.6677
R1463 VTAIL.n25 VTAIL.n24 15.6677
R1464 VTAIL.n182 VTAIL.n181 15.6677
R1465 VTAIL.n104 VTAIL.n103 15.6677
R1466 VTAIL.n307 VTAIL.n236 13.1884
R1467 VTAIL.n73 VTAIL.n2 13.1884
R1468 VTAIL.n229 VTAIL.n158 13.1884
R1469 VTAIL.n151 VTAIL.n80 13.1884
R1470 VTAIL.n262 VTAIL.n261 12.8005
R1471 VTAIL.n303 VTAIL.n302 12.8005
R1472 VTAIL.n308 VTAIL.n234 12.8005
R1473 VTAIL.n28 VTAIL.n27 12.8005
R1474 VTAIL.n69 VTAIL.n68 12.8005
R1475 VTAIL.n74 VTAIL.n0 12.8005
R1476 VTAIL.n230 VTAIL.n156 12.8005
R1477 VTAIL.n225 VTAIL.n160 12.8005
R1478 VTAIL.n185 VTAIL.n184 12.8005
R1479 VTAIL.n152 VTAIL.n78 12.8005
R1480 VTAIL.n147 VTAIL.n82 12.8005
R1481 VTAIL.n107 VTAIL.n106 12.8005
R1482 VTAIL.n265 VTAIL.n256 12.0247
R1483 VTAIL.n301 VTAIL.n238 12.0247
R1484 VTAIL.n31 VTAIL.n22 12.0247
R1485 VTAIL.n67 VTAIL.n4 12.0247
R1486 VTAIL.n224 VTAIL.n161 12.0247
R1487 VTAIL.n188 VTAIL.n179 12.0247
R1488 VTAIL.n146 VTAIL.n83 12.0247
R1489 VTAIL.n110 VTAIL.n101 12.0247
R1490 VTAIL.n266 VTAIL.n254 11.249
R1491 VTAIL.n298 VTAIL.n297 11.249
R1492 VTAIL.n32 VTAIL.n20 11.249
R1493 VTAIL.n64 VTAIL.n63 11.249
R1494 VTAIL.n221 VTAIL.n220 11.249
R1495 VTAIL.n189 VTAIL.n177 11.249
R1496 VTAIL.n143 VTAIL.n142 11.249
R1497 VTAIL.n111 VTAIL.n99 11.249
R1498 VTAIL.n270 VTAIL.n269 10.4732
R1499 VTAIL.n294 VTAIL.n240 10.4732
R1500 VTAIL.n36 VTAIL.n35 10.4732
R1501 VTAIL.n60 VTAIL.n6 10.4732
R1502 VTAIL.n217 VTAIL.n163 10.4732
R1503 VTAIL.n193 VTAIL.n192 10.4732
R1504 VTAIL.n139 VTAIL.n85 10.4732
R1505 VTAIL.n115 VTAIL.n114 10.4732
R1506 VTAIL.n273 VTAIL.n252 9.69747
R1507 VTAIL.n293 VTAIL.n242 9.69747
R1508 VTAIL.n39 VTAIL.n18 9.69747
R1509 VTAIL.n59 VTAIL.n8 9.69747
R1510 VTAIL.n216 VTAIL.n165 9.69747
R1511 VTAIL.n196 VTAIL.n175 9.69747
R1512 VTAIL.n138 VTAIL.n87 9.69747
R1513 VTAIL.n118 VTAIL.n97 9.69747
R1514 VTAIL.n310 VTAIL.n309 9.45567
R1515 VTAIL.n76 VTAIL.n75 9.45567
R1516 VTAIL.n232 VTAIL.n231 9.45567
R1517 VTAIL.n154 VTAIL.n153 9.45567
R1518 VTAIL.n309 VTAIL.n308 9.3005
R1519 VTAIL.n248 VTAIL.n247 9.3005
R1520 VTAIL.n277 VTAIL.n276 9.3005
R1521 VTAIL.n275 VTAIL.n274 9.3005
R1522 VTAIL.n252 VTAIL.n251 9.3005
R1523 VTAIL.n269 VTAIL.n268 9.3005
R1524 VTAIL.n267 VTAIL.n266 9.3005
R1525 VTAIL.n256 VTAIL.n255 9.3005
R1526 VTAIL.n261 VTAIL.n260 9.3005
R1527 VTAIL.n283 VTAIL.n282 9.3005
R1528 VTAIL.n285 VTAIL.n284 9.3005
R1529 VTAIL.n244 VTAIL.n243 9.3005
R1530 VTAIL.n291 VTAIL.n290 9.3005
R1531 VTAIL.n293 VTAIL.n292 9.3005
R1532 VTAIL.n240 VTAIL.n239 9.3005
R1533 VTAIL.n299 VTAIL.n298 9.3005
R1534 VTAIL.n301 VTAIL.n300 9.3005
R1535 VTAIL.n302 VTAIL.n235 9.3005
R1536 VTAIL.n75 VTAIL.n74 9.3005
R1537 VTAIL.n14 VTAIL.n13 9.3005
R1538 VTAIL.n43 VTAIL.n42 9.3005
R1539 VTAIL.n41 VTAIL.n40 9.3005
R1540 VTAIL.n18 VTAIL.n17 9.3005
R1541 VTAIL.n35 VTAIL.n34 9.3005
R1542 VTAIL.n33 VTAIL.n32 9.3005
R1543 VTAIL.n22 VTAIL.n21 9.3005
R1544 VTAIL.n27 VTAIL.n26 9.3005
R1545 VTAIL.n49 VTAIL.n48 9.3005
R1546 VTAIL.n51 VTAIL.n50 9.3005
R1547 VTAIL.n10 VTAIL.n9 9.3005
R1548 VTAIL.n57 VTAIL.n56 9.3005
R1549 VTAIL.n59 VTAIL.n58 9.3005
R1550 VTAIL.n6 VTAIL.n5 9.3005
R1551 VTAIL.n65 VTAIL.n64 9.3005
R1552 VTAIL.n67 VTAIL.n66 9.3005
R1553 VTAIL.n68 VTAIL.n1 9.3005
R1554 VTAIL.n208 VTAIL.n207 9.3005
R1555 VTAIL.n167 VTAIL.n166 9.3005
R1556 VTAIL.n214 VTAIL.n213 9.3005
R1557 VTAIL.n216 VTAIL.n215 9.3005
R1558 VTAIL.n163 VTAIL.n162 9.3005
R1559 VTAIL.n222 VTAIL.n221 9.3005
R1560 VTAIL.n224 VTAIL.n223 9.3005
R1561 VTAIL.n160 VTAIL.n157 9.3005
R1562 VTAIL.n231 VTAIL.n230 9.3005
R1563 VTAIL.n206 VTAIL.n205 9.3005
R1564 VTAIL.n171 VTAIL.n170 9.3005
R1565 VTAIL.n200 VTAIL.n199 9.3005
R1566 VTAIL.n198 VTAIL.n197 9.3005
R1567 VTAIL.n175 VTAIL.n174 9.3005
R1568 VTAIL.n192 VTAIL.n191 9.3005
R1569 VTAIL.n190 VTAIL.n189 9.3005
R1570 VTAIL.n179 VTAIL.n178 9.3005
R1571 VTAIL.n184 VTAIL.n183 9.3005
R1572 VTAIL.n130 VTAIL.n129 9.3005
R1573 VTAIL.n89 VTAIL.n88 9.3005
R1574 VTAIL.n136 VTAIL.n135 9.3005
R1575 VTAIL.n138 VTAIL.n137 9.3005
R1576 VTAIL.n85 VTAIL.n84 9.3005
R1577 VTAIL.n144 VTAIL.n143 9.3005
R1578 VTAIL.n146 VTAIL.n145 9.3005
R1579 VTAIL.n82 VTAIL.n79 9.3005
R1580 VTAIL.n153 VTAIL.n152 9.3005
R1581 VTAIL.n128 VTAIL.n127 9.3005
R1582 VTAIL.n93 VTAIL.n92 9.3005
R1583 VTAIL.n122 VTAIL.n121 9.3005
R1584 VTAIL.n120 VTAIL.n119 9.3005
R1585 VTAIL.n97 VTAIL.n96 9.3005
R1586 VTAIL.n114 VTAIL.n113 9.3005
R1587 VTAIL.n112 VTAIL.n111 9.3005
R1588 VTAIL.n101 VTAIL.n100 9.3005
R1589 VTAIL.n106 VTAIL.n105 9.3005
R1590 VTAIL.n274 VTAIL.n250 8.92171
R1591 VTAIL.n290 VTAIL.n289 8.92171
R1592 VTAIL.n40 VTAIL.n16 8.92171
R1593 VTAIL.n56 VTAIL.n55 8.92171
R1594 VTAIL.n213 VTAIL.n212 8.92171
R1595 VTAIL.n197 VTAIL.n173 8.92171
R1596 VTAIL.n135 VTAIL.n134 8.92171
R1597 VTAIL.n119 VTAIL.n95 8.92171
R1598 VTAIL.n278 VTAIL.n277 8.14595
R1599 VTAIL.n286 VTAIL.n244 8.14595
R1600 VTAIL.n44 VTAIL.n43 8.14595
R1601 VTAIL.n52 VTAIL.n10 8.14595
R1602 VTAIL.n209 VTAIL.n167 8.14595
R1603 VTAIL.n201 VTAIL.n200 8.14595
R1604 VTAIL.n131 VTAIL.n89 8.14595
R1605 VTAIL.n123 VTAIL.n122 8.14595
R1606 VTAIL.n281 VTAIL.n248 7.3702
R1607 VTAIL.n285 VTAIL.n246 7.3702
R1608 VTAIL.n47 VTAIL.n14 7.3702
R1609 VTAIL.n51 VTAIL.n12 7.3702
R1610 VTAIL.n208 VTAIL.n169 7.3702
R1611 VTAIL.n204 VTAIL.n171 7.3702
R1612 VTAIL.n130 VTAIL.n91 7.3702
R1613 VTAIL.n126 VTAIL.n93 7.3702
R1614 VTAIL.n282 VTAIL.n281 6.59444
R1615 VTAIL.n282 VTAIL.n246 6.59444
R1616 VTAIL.n48 VTAIL.n47 6.59444
R1617 VTAIL.n48 VTAIL.n12 6.59444
R1618 VTAIL.n205 VTAIL.n169 6.59444
R1619 VTAIL.n205 VTAIL.n204 6.59444
R1620 VTAIL.n127 VTAIL.n91 6.59444
R1621 VTAIL.n127 VTAIL.n126 6.59444
R1622 VTAIL.n278 VTAIL.n248 5.81868
R1623 VTAIL.n286 VTAIL.n285 5.81868
R1624 VTAIL.n44 VTAIL.n14 5.81868
R1625 VTAIL.n52 VTAIL.n51 5.81868
R1626 VTAIL.n209 VTAIL.n208 5.81868
R1627 VTAIL.n201 VTAIL.n171 5.81868
R1628 VTAIL.n131 VTAIL.n130 5.81868
R1629 VTAIL.n123 VTAIL.n93 5.81868
R1630 VTAIL.n277 VTAIL.n250 5.04292
R1631 VTAIL.n289 VTAIL.n244 5.04292
R1632 VTAIL.n43 VTAIL.n16 5.04292
R1633 VTAIL.n55 VTAIL.n10 5.04292
R1634 VTAIL.n212 VTAIL.n167 5.04292
R1635 VTAIL.n200 VTAIL.n173 5.04292
R1636 VTAIL.n134 VTAIL.n89 5.04292
R1637 VTAIL.n122 VTAIL.n95 5.04292
R1638 VTAIL.n260 VTAIL.n259 4.38563
R1639 VTAIL.n26 VTAIL.n25 4.38563
R1640 VTAIL.n183 VTAIL.n182 4.38563
R1641 VTAIL.n105 VTAIL.n104 4.38563
R1642 VTAIL.n274 VTAIL.n273 4.26717
R1643 VTAIL.n290 VTAIL.n242 4.26717
R1644 VTAIL.n40 VTAIL.n39 4.26717
R1645 VTAIL.n56 VTAIL.n8 4.26717
R1646 VTAIL.n213 VTAIL.n165 4.26717
R1647 VTAIL.n197 VTAIL.n196 4.26717
R1648 VTAIL.n135 VTAIL.n87 4.26717
R1649 VTAIL.n119 VTAIL.n118 4.26717
R1650 VTAIL.n270 VTAIL.n252 3.49141
R1651 VTAIL.n294 VTAIL.n293 3.49141
R1652 VTAIL.n36 VTAIL.n18 3.49141
R1653 VTAIL.n60 VTAIL.n59 3.49141
R1654 VTAIL.n217 VTAIL.n216 3.49141
R1655 VTAIL.n193 VTAIL.n175 3.49141
R1656 VTAIL.n139 VTAIL.n138 3.49141
R1657 VTAIL.n115 VTAIL.n97 3.49141
R1658 VTAIL.n269 VTAIL.n254 2.71565
R1659 VTAIL.n297 VTAIL.n240 2.71565
R1660 VTAIL.n35 VTAIL.n20 2.71565
R1661 VTAIL.n63 VTAIL.n6 2.71565
R1662 VTAIL.n220 VTAIL.n163 2.71565
R1663 VTAIL.n192 VTAIL.n177 2.71565
R1664 VTAIL.n142 VTAIL.n85 2.71565
R1665 VTAIL.n114 VTAIL.n99 2.71565
R1666 VTAIL.n266 VTAIL.n265 1.93989
R1667 VTAIL.n298 VTAIL.n238 1.93989
R1668 VTAIL.n32 VTAIL.n31 1.93989
R1669 VTAIL.n64 VTAIL.n4 1.93989
R1670 VTAIL.n221 VTAIL.n161 1.93989
R1671 VTAIL.n189 VTAIL.n188 1.93989
R1672 VTAIL.n143 VTAIL.n83 1.93989
R1673 VTAIL.n111 VTAIL.n110 1.93989
R1674 VTAIL.n233 VTAIL.n155 1.54791
R1675 VTAIL.n262 VTAIL.n256 1.16414
R1676 VTAIL.n303 VTAIL.n301 1.16414
R1677 VTAIL.n310 VTAIL.n234 1.16414
R1678 VTAIL.n28 VTAIL.n22 1.16414
R1679 VTAIL.n69 VTAIL.n67 1.16414
R1680 VTAIL.n76 VTAIL.n0 1.16414
R1681 VTAIL.n232 VTAIL.n156 1.16414
R1682 VTAIL.n225 VTAIL.n224 1.16414
R1683 VTAIL.n185 VTAIL.n179 1.16414
R1684 VTAIL.n154 VTAIL.n78 1.16414
R1685 VTAIL.n147 VTAIL.n146 1.16414
R1686 VTAIL.n107 VTAIL.n101 1.16414
R1687 VTAIL VTAIL.n77 1.06731
R1688 VTAIL VTAIL.n311 0.481103
R1689 VTAIL.n261 VTAIL.n258 0.388379
R1690 VTAIL.n302 VTAIL.n236 0.388379
R1691 VTAIL.n308 VTAIL.n307 0.388379
R1692 VTAIL.n27 VTAIL.n24 0.388379
R1693 VTAIL.n68 VTAIL.n2 0.388379
R1694 VTAIL.n74 VTAIL.n73 0.388379
R1695 VTAIL.n230 VTAIL.n229 0.388379
R1696 VTAIL.n160 VTAIL.n158 0.388379
R1697 VTAIL.n184 VTAIL.n181 0.388379
R1698 VTAIL.n152 VTAIL.n151 0.388379
R1699 VTAIL.n82 VTAIL.n80 0.388379
R1700 VTAIL.n106 VTAIL.n103 0.388379
R1701 VTAIL.n260 VTAIL.n255 0.155672
R1702 VTAIL.n267 VTAIL.n255 0.155672
R1703 VTAIL.n268 VTAIL.n267 0.155672
R1704 VTAIL.n268 VTAIL.n251 0.155672
R1705 VTAIL.n275 VTAIL.n251 0.155672
R1706 VTAIL.n276 VTAIL.n275 0.155672
R1707 VTAIL.n276 VTAIL.n247 0.155672
R1708 VTAIL.n283 VTAIL.n247 0.155672
R1709 VTAIL.n284 VTAIL.n283 0.155672
R1710 VTAIL.n284 VTAIL.n243 0.155672
R1711 VTAIL.n291 VTAIL.n243 0.155672
R1712 VTAIL.n292 VTAIL.n291 0.155672
R1713 VTAIL.n292 VTAIL.n239 0.155672
R1714 VTAIL.n299 VTAIL.n239 0.155672
R1715 VTAIL.n300 VTAIL.n299 0.155672
R1716 VTAIL.n300 VTAIL.n235 0.155672
R1717 VTAIL.n309 VTAIL.n235 0.155672
R1718 VTAIL.n26 VTAIL.n21 0.155672
R1719 VTAIL.n33 VTAIL.n21 0.155672
R1720 VTAIL.n34 VTAIL.n33 0.155672
R1721 VTAIL.n34 VTAIL.n17 0.155672
R1722 VTAIL.n41 VTAIL.n17 0.155672
R1723 VTAIL.n42 VTAIL.n41 0.155672
R1724 VTAIL.n42 VTAIL.n13 0.155672
R1725 VTAIL.n49 VTAIL.n13 0.155672
R1726 VTAIL.n50 VTAIL.n49 0.155672
R1727 VTAIL.n50 VTAIL.n9 0.155672
R1728 VTAIL.n57 VTAIL.n9 0.155672
R1729 VTAIL.n58 VTAIL.n57 0.155672
R1730 VTAIL.n58 VTAIL.n5 0.155672
R1731 VTAIL.n65 VTAIL.n5 0.155672
R1732 VTAIL.n66 VTAIL.n65 0.155672
R1733 VTAIL.n66 VTAIL.n1 0.155672
R1734 VTAIL.n75 VTAIL.n1 0.155672
R1735 VTAIL.n231 VTAIL.n157 0.155672
R1736 VTAIL.n223 VTAIL.n157 0.155672
R1737 VTAIL.n223 VTAIL.n222 0.155672
R1738 VTAIL.n222 VTAIL.n162 0.155672
R1739 VTAIL.n215 VTAIL.n162 0.155672
R1740 VTAIL.n215 VTAIL.n214 0.155672
R1741 VTAIL.n214 VTAIL.n166 0.155672
R1742 VTAIL.n207 VTAIL.n166 0.155672
R1743 VTAIL.n207 VTAIL.n206 0.155672
R1744 VTAIL.n206 VTAIL.n170 0.155672
R1745 VTAIL.n199 VTAIL.n170 0.155672
R1746 VTAIL.n199 VTAIL.n198 0.155672
R1747 VTAIL.n198 VTAIL.n174 0.155672
R1748 VTAIL.n191 VTAIL.n174 0.155672
R1749 VTAIL.n191 VTAIL.n190 0.155672
R1750 VTAIL.n190 VTAIL.n178 0.155672
R1751 VTAIL.n183 VTAIL.n178 0.155672
R1752 VTAIL.n153 VTAIL.n79 0.155672
R1753 VTAIL.n145 VTAIL.n79 0.155672
R1754 VTAIL.n145 VTAIL.n144 0.155672
R1755 VTAIL.n144 VTAIL.n84 0.155672
R1756 VTAIL.n137 VTAIL.n84 0.155672
R1757 VTAIL.n137 VTAIL.n136 0.155672
R1758 VTAIL.n136 VTAIL.n88 0.155672
R1759 VTAIL.n129 VTAIL.n88 0.155672
R1760 VTAIL.n129 VTAIL.n128 0.155672
R1761 VTAIL.n128 VTAIL.n92 0.155672
R1762 VTAIL.n121 VTAIL.n92 0.155672
R1763 VTAIL.n121 VTAIL.n120 0.155672
R1764 VTAIL.n120 VTAIL.n96 0.155672
R1765 VTAIL.n113 VTAIL.n96 0.155672
R1766 VTAIL.n113 VTAIL.n112 0.155672
R1767 VTAIL.n112 VTAIL.n100 0.155672
R1768 VTAIL.n105 VTAIL.n100 0.155672
R1769 VDD1.n72 VDD1.n0 289.615
R1770 VDD1.n149 VDD1.n77 289.615
R1771 VDD1.n73 VDD1.n72 185
R1772 VDD1.n71 VDD1.n2 185
R1773 VDD1.n70 VDD1.n69 185
R1774 VDD1.n5 VDD1.n3 185
R1775 VDD1.n64 VDD1.n63 185
R1776 VDD1.n62 VDD1.n61 185
R1777 VDD1.n9 VDD1.n8 185
R1778 VDD1.n56 VDD1.n55 185
R1779 VDD1.n54 VDD1.n53 185
R1780 VDD1.n13 VDD1.n12 185
R1781 VDD1.n48 VDD1.n47 185
R1782 VDD1.n46 VDD1.n45 185
R1783 VDD1.n17 VDD1.n16 185
R1784 VDD1.n40 VDD1.n39 185
R1785 VDD1.n38 VDD1.n37 185
R1786 VDD1.n21 VDD1.n20 185
R1787 VDD1.n32 VDD1.n31 185
R1788 VDD1.n30 VDD1.n29 185
R1789 VDD1.n25 VDD1.n24 185
R1790 VDD1.n101 VDD1.n100 185
R1791 VDD1.n106 VDD1.n105 185
R1792 VDD1.n108 VDD1.n107 185
R1793 VDD1.n97 VDD1.n96 185
R1794 VDD1.n114 VDD1.n113 185
R1795 VDD1.n116 VDD1.n115 185
R1796 VDD1.n93 VDD1.n92 185
R1797 VDD1.n122 VDD1.n121 185
R1798 VDD1.n124 VDD1.n123 185
R1799 VDD1.n89 VDD1.n88 185
R1800 VDD1.n130 VDD1.n129 185
R1801 VDD1.n132 VDD1.n131 185
R1802 VDD1.n85 VDD1.n84 185
R1803 VDD1.n138 VDD1.n137 185
R1804 VDD1.n140 VDD1.n139 185
R1805 VDD1.n81 VDD1.n80 185
R1806 VDD1.n147 VDD1.n146 185
R1807 VDD1.n148 VDD1.n79 185
R1808 VDD1.n150 VDD1.n149 185
R1809 VDD1.n26 VDD1.t1 147.659
R1810 VDD1.n102 VDD1.t0 147.659
R1811 VDD1.n72 VDD1.n71 104.615
R1812 VDD1.n71 VDD1.n70 104.615
R1813 VDD1.n70 VDD1.n3 104.615
R1814 VDD1.n63 VDD1.n3 104.615
R1815 VDD1.n63 VDD1.n62 104.615
R1816 VDD1.n62 VDD1.n8 104.615
R1817 VDD1.n55 VDD1.n8 104.615
R1818 VDD1.n55 VDD1.n54 104.615
R1819 VDD1.n54 VDD1.n12 104.615
R1820 VDD1.n47 VDD1.n12 104.615
R1821 VDD1.n47 VDD1.n46 104.615
R1822 VDD1.n46 VDD1.n16 104.615
R1823 VDD1.n39 VDD1.n16 104.615
R1824 VDD1.n39 VDD1.n38 104.615
R1825 VDD1.n38 VDD1.n20 104.615
R1826 VDD1.n31 VDD1.n20 104.615
R1827 VDD1.n31 VDD1.n30 104.615
R1828 VDD1.n30 VDD1.n24 104.615
R1829 VDD1.n106 VDD1.n100 104.615
R1830 VDD1.n107 VDD1.n106 104.615
R1831 VDD1.n107 VDD1.n96 104.615
R1832 VDD1.n114 VDD1.n96 104.615
R1833 VDD1.n115 VDD1.n114 104.615
R1834 VDD1.n115 VDD1.n92 104.615
R1835 VDD1.n122 VDD1.n92 104.615
R1836 VDD1.n123 VDD1.n122 104.615
R1837 VDD1.n123 VDD1.n88 104.615
R1838 VDD1.n130 VDD1.n88 104.615
R1839 VDD1.n131 VDD1.n130 104.615
R1840 VDD1.n131 VDD1.n84 104.615
R1841 VDD1.n138 VDD1.n84 104.615
R1842 VDD1.n139 VDD1.n138 104.615
R1843 VDD1.n139 VDD1.n80 104.615
R1844 VDD1.n147 VDD1.n80 104.615
R1845 VDD1.n148 VDD1.n147 104.615
R1846 VDD1.n149 VDD1.n148 104.615
R1847 VDD1 VDD1.n153 91.518
R1848 VDD1.t1 VDD1.n24 52.3082
R1849 VDD1.t0 VDD1.n100 52.3082
R1850 VDD1 VDD1.n76 51.0126
R1851 VDD1.n26 VDD1.n25 15.6677
R1852 VDD1.n102 VDD1.n101 15.6677
R1853 VDD1.n73 VDD1.n2 13.1884
R1854 VDD1.n150 VDD1.n79 13.1884
R1855 VDD1.n74 VDD1.n0 12.8005
R1856 VDD1.n69 VDD1.n4 12.8005
R1857 VDD1.n29 VDD1.n28 12.8005
R1858 VDD1.n105 VDD1.n104 12.8005
R1859 VDD1.n146 VDD1.n145 12.8005
R1860 VDD1.n151 VDD1.n77 12.8005
R1861 VDD1.n68 VDD1.n5 12.0247
R1862 VDD1.n32 VDD1.n23 12.0247
R1863 VDD1.n108 VDD1.n99 12.0247
R1864 VDD1.n144 VDD1.n81 12.0247
R1865 VDD1.n65 VDD1.n64 11.249
R1866 VDD1.n33 VDD1.n21 11.249
R1867 VDD1.n109 VDD1.n97 11.249
R1868 VDD1.n141 VDD1.n140 11.249
R1869 VDD1.n61 VDD1.n7 10.4732
R1870 VDD1.n37 VDD1.n36 10.4732
R1871 VDD1.n113 VDD1.n112 10.4732
R1872 VDD1.n137 VDD1.n83 10.4732
R1873 VDD1.n60 VDD1.n9 9.69747
R1874 VDD1.n40 VDD1.n19 9.69747
R1875 VDD1.n116 VDD1.n95 9.69747
R1876 VDD1.n136 VDD1.n85 9.69747
R1877 VDD1.n76 VDD1.n75 9.45567
R1878 VDD1.n153 VDD1.n152 9.45567
R1879 VDD1.n52 VDD1.n51 9.3005
R1880 VDD1.n11 VDD1.n10 9.3005
R1881 VDD1.n58 VDD1.n57 9.3005
R1882 VDD1.n60 VDD1.n59 9.3005
R1883 VDD1.n7 VDD1.n6 9.3005
R1884 VDD1.n66 VDD1.n65 9.3005
R1885 VDD1.n68 VDD1.n67 9.3005
R1886 VDD1.n4 VDD1.n1 9.3005
R1887 VDD1.n75 VDD1.n74 9.3005
R1888 VDD1.n50 VDD1.n49 9.3005
R1889 VDD1.n15 VDD1.n14 9.3005
R1890 VDD1.n44 VDD1.n43 9.3005
R1891 VDD1.n42 VDD1.n41 9.3005
R1892 VDD1.n19 VDD1.n18 9.3005
R1893 VDD1.n36 VDD1.n35 9.3005
R1894 VDD1.n34 VDD1.n33 9.3005
R1895 VDD1.n23 VDD1.n22 9.3005
R1896 VDD1.n28 VDD1.n27 9.3005
R1897 VDD1.n152 VDD1.n151 9.3005
R1898 VDD1.n91 VDD1.n90 9.3005
R1899 VDD1.n120 VDD1.n119 9.3005
R1900 VDD1.n118 VDD1.n117 9.3005
R1901 VDD1.n95 VDD1.n94 9.3005
R1902 VDD1.n112 VDD1.n111 9.3005
R1903 VDD1.n110 VDD1.n109 9.3005
R1904 VDD1.n99 VDD1.n98 9.3005
R1905 VDD1.n104 VDD1.n103 9.3005
R1906 VDD1.n126 VDD1.n125 9.3005
R1907 VDD1.n128 VDD1.n127 9.3005
R1908 VDD1.n87 VDD1.n86 9.3005
R1909 VDD1.n134 VDD1.n133 9.3005
R1910 VDD1.n136 VDD1.n135 9.3005
R1911 VDD1.n83 VDD1.n82 9.3005
R1912 VDD1.n142 VDD1.n141 9.3005
R1913 VDD1.n144 VDD1.n143 9.3005
R1914 VDD1.n145 VDD1.n78 9.3005
R1915 VDD1.n57 VDD1.n56 8.92171
R1916 VDD1.n41 VDD1.n17 8.92171
R1917 VDD1.n117 VDD1.n93 8.92171
R1918 VDD1.n133 VDD1.n132 8.92171
R1919 VDD1.n53 VDD1.n11 8.14595
R1920 VDD1.n45 VDD1.n44 8.14595
R1921 VDD1.n121 VDD1.n120 8.14595
R1922 VDD1.n129 VDD1.n87 8.14595
R1923 VDD1.n52 VDD1.n13 7.3702
R1924 VDD1.n48 VDD1.n15 7.3702
R1925 VDD1.n124 VDD1.n91 7.3702
R1926 VDD1.n128 VDD1.n89 7.3702
R1927 VDD1.n49 VDD1.n13 6.59444
R1928 VDD1.n49 VDD1.n48 6.59444
R1929 VDD1.n125 VDD1.n124 6.59444
R1930 VDD1.n125 VDD1.n89 6.59444
R1931 VDD1.n53 VDD1.n52 5.81868
R1932 VDD1.n45 VDD1.n15 5.81868
R1933 VDD1.n121 VDD1.n91 5.81868
R1934 VDD1.n129 VDD1.n128 5.81868
R1935 VDD1.n56 VDD1.n11 5.04292
R1936 VDD1.n44 VDD1.n17 5.04292
R1937 VDD1.n120 VDD1.n93 5.04292
R1938 VDD1.n132 VDD1.n87 5.04292
R1939 VDD1.n27 VDD1.n26 4.38563
R1940 VDD1.n103 VDD1.n102 4.38563
R1941 VDD1.n57 VDD1.n9 4.26717
R1942 VDD1.n41 VDD1.n40 4.26717
R1943 VDD1.n117 VDD1.n116 4.26717
R1944 VDD1.n133 VDD1.n85 4.26717
R1945 VDD1.n61 VDD1.n60 3.49141
R1946 VDD1.n37 VDD1.n19 3.49141
R1947 VDD1.n113 VDD1.n95 3.49141
R1948 VDD1.n137 VDD1.n136 3.49141
R1949 VDD1.n64 VDD1.n7 2.71565
R1950 VDD1.n36 VDD1.n21 2.71565
R1951 VDD1.n112 VDD1.n97 2.71565
R1952 VDD1.n140 VDD1.n83 2.71565
R1953 VDD1.n65 VDD1.n5 1.93989
R1954 VDD1.n33 VDD1.n32 1.93989
R1955 VDD1.n109 VDD1.n108 1.93989
R1956 VDD1.n141 VDD1.n81 1.93989
R1957 VDD1.n76 VDD1.n0 1.16414
R1958 VDD1.n69 VDD1.n68 1.16414
R1959 VDD1.n29 VDD1.n23 1.16414
R1960 VDD1.n105 VDD1.n99 1.16414
R1961 VDD1.n146 VDD1.n144 1.16414
R1962 VDD1.n153 VDD1.n77 1.16414
R1963 VDD1.n74 VDD1.n73 0.388379
R1964 VDD1.n4 VDD1.n2 0.388379
R1965 VDD1.n28 VDD1.n25 0.388379
R1966 VDD1.n104 VDD1.n101 0.388379
R1967 VDD1.n145 VDD1.n79 0.388379
R1968 VDD1.n151 VDD1.n150 0.388379
R1969 VDD1.n75 VDD1.n1 0.155672
R1970 VDD1.n67 VDD1.n1 0.155672
R1971 VDD1.n67 VDD1.n66 0.155672
R1972 VDD1.n66 VDD1.n6 0.155672
R1973 VDD1.n59 VDD1.n6 0.155672
R1974 VDD1.n59 VDD1.n58 0.155672
R1975 VDD1.n58 VDD1.n10 0.155672
R1976 VDD1.n51 VDD1.n10 0.155672
R1977 VDD1.n51 VDD1.n50 0.155672
R1978 VDD1.n50 VDD1.n14 0.155672
R1979 VDD1.n43 VDD1.n14 0.155672
R1980 VDD1.n43 VDD1.n42 0.155672
R1981 VDD1.n42 VDD1.n18 0.155672
R1982 VDD1.n35 VDD1.n18 0.155672
R1983 VDD1.n35 VDD1.n34 0.155672
R1984 VDD1.n34 VDD1.n22 0.155672
R1985 VDD1.n27 VDD1.n22 0.155672
R1986 VDD1.n103 VDD1.n98 0.155672
R1987 VDD1.n110 VDD1.n98 0.155672
R1988 VDD1.n111 VDD1.n110 0.155672
R1989 VDD1.n111 VDD1.n94 0.155672
R1990 VDD1.n118 VDD1.n94 0.155672
R1991 VDD1.n119 VDD1.n118 0.155672
R1992 VDD1.n119 VDD1.n90 0.155672
R1993 VDD1.n126 VDD1.n90 0.155672
R1994 VDD1.n127 VDD1.n126 0.155672
R1995 VDD1.n127 VDD1.n86 0.155672
R1996 VDD1.n134 VDD1.n86 0.155672
R1997 VDD1.n135 VDD1.n134 0.155672
R1998 VDD1.n135 VDD1.n82 0.155672
R1999 VDD1.n142 VDD1.n82 0.155672
R2000 VDD1.n143 VDD1.n142 0.155672
R2001 VDD1.n143 VDD1.n78 0.155672
R2002 VDD1.n152 VDD1.n78 0.155672
R2003 VN VN.t0 249.827
R2004 VN VN.t1 205.036
R2005 VDD2.n149 VDD2.n77 289.615
R2006 VDD2.n72 VDD2.n0 289.615
R2007 VDD2.n150 VDD2.n149 185
R2008 VDD2.n148 VDD2.n79 185
R2009 VDD2.n147 VDD2.n146 185
R2010 VDD2.n82 VDD2.n80 185
R2011 VDD2.n141 VDD2.n140 185
R2012 VDD2.n139 VDD2.n138 185
R2013 VDD2.n86 VDD2.n85 185
R2014 VDD2.n133 VDD2.n132 185
R2015 VDD2.n131 VDD2.n130 185
R2016 VDD2.n90 VDD2.n89 185
R2017 VDD2.n125 VDD2.n124 185
R2018 VDD2.n123 VDD2.n122 185
R2019 VDD2.n94 VDD2.n93 185
R2020 VDD2.n117 VDD2.n116 185
R2021 VDD2.n115 VDD2.n114 185
R2022 VDD2.n98 VDD2.n97 185
R2023 VDD2.n109 VDD2.n108 185
R2024 VDD2.n107 VDD2.n106 185
R2025 VDD2.n102 VDD2.n101 185
R2026 VDD2.n24 VDD2.n23 185
R2027 VDD2.n29 VDD2.n28 185
R2028 VDD2.n31 VDD2.n30 185
R2029 VDD2.n20 VDD2.n19 185
R2030 VDD2.n37 VDD2.n36 185
R2031 VDD2.n39 VDD2.n38 185
R2032 VDD2.n16 VDD2.n15 185
R2033 VDD2.n45 VDD2.n44 185
R2034 VDD2.n47 VDD2.n46 185
R2035 VDD2.n12 VDD2.n11 185
R2036 VDD2.n53 VDD2.n52 185
R2037 VDD2.n55 VDD2.n54 185
R2038 VDD2.n8 VDD2.n7 185
R2039 VDD2.n61 VDD2.n60 185
R2040 VDD2.n63 VDD2.n62 185
R2041 VDD2.n4 VDD2.n3 185
R2042 VDD2.n70 VDD2.n69 185
R2043 VDD2.n71 VDD2.n2 185
R2044 VDD2.n73 VDD2.n72 185
R2045 VDD2.n103 VDD2.t1 147.659
R2046 VDD2.n25 VDD2.t0 147.659
R2047 VDD2.n149 VDD2.n148 104.615
R2048 VDD2.n148 VDD2.n147 104.615
R2049 VDD2.n147 VDD2.n80 104.615
R2050 VDD2.n140 VDD2.n80 104.615
R2051 VDD2.n140 VDD2.n139 104.615
R2052 VDD2.n139 VDD2.n85 104.615
R2053 VDD2.n132 VDD2.n85 104.615
R2054 VDD2.n132 VDD2.n131 104.615
R2055 VDD2.n131 VDD2.n89 104.615
R2056 VDD2.n124 VDD2.n89 104.615
R2057 VDD2.n124 VDD2.n123 104.615
R2058 VDD2.n123 VDD2.n93 104.615
R2059 VDD2.n116 VDD2.n93 104.615
R2060 VDD2.n116 VDD2.n115 104.615
R2061 VDD2.n115 VDD2.n97 104.615
R2062 VDD2.n108 VDD2.n97 104.615
R2063 VDD2.n108 VDD2.n107 104.615
R2064 VDD2.n107 VDD2.n101 104.615
R2065 VDD2.n29 VDD2.n23 104.615
R2066 VDD2.n30 VDD2.n29 104.615
R2067 VDD2.n30 VDD2.n19 104.615
R2068 VDD2.n37 VDD2.n19 104.615
R2069 VDD2.n38 VDD2.n37 104.615
R2070 VDD2.n38 VDD2.n15 104.615
R2071 VDD2.n45 VDD2.n15 104.615
R2072 VDD2.n46 VDD2.n45 104.615
R2073 VDD2.n46 VDD2.n11 104.615
R2074 VDD2.n53 VDD2.n11 104.615
R2075 VDD2.n54 VDD2.n53 104.615
R2076 VDD2.n54 VDD2.n7 104.615
R2077 VDD2.n61 VDD2.n7 104.615
R2078 VDD2.n62 VDD2.n61 104.615
R2079 VDD2.n62 VDD2.n3 104.615
R2080 VDD2.n70 VDD2.n3 104.615
R2081 VDD2.n71 VDD2.n70 104.615
R2082 VDD2.n72 VDD2.n71 104.615
R2083 VDD2.n154 VDD2.n76 90.4544
R2084 VDD2.t1 VDD2.n101 52.3082
R2085 VDD2.t0 VDD2.n23 52.3082
R2086 VDD2.n154 VDD2.n153 50.4157
R2087 VDD2.n103 VDD2.n102 15.6677
R2088 VDD2.n25 VDD2.n24 15.6677
R2089 VDD2.n150 VDD2.n79 13.1884
R2090 VDD2.n73 VDD2.n2 13.1884
R2091 VDD2.n151 VDD2.n77 12.8005
R2092 VDD2.n146 VDD2.n81 12.8005
R2093 VDD2.n106 VDD2.n105 12.8005
R2094 VDD2.n28 VDD2.n27 12.8005
R2095 VDD2.n69 VDD2.n68 12.8005
R2096 VDD2.n74 VDD2.n0 12.8005
R2097 VDD2.n145 VDD2.n82 12.0247
R2098 VDD2.n109 VDD2.n100 12.0247
R2099 VDD2.n31 VDD2.n22 12.0247
R2100 VDD2.n67 VDD2.n4 12.0247
R2101 VDD2.n142 VDD2.n141 11.249
R2102 VDD2.n110 VDD2.n98 11.249
R2103 VDD2.n32 VDD2.n20 11.249
R2104 VDD2.n64 VDD2.n63 11.249
R2105 VDD2.n138 VDD2.n84 10.4732
R2106 VDD2.n114 VDD2.n113 10.4732
R2107 VDD2.n36 VDD2.n35 10.4732
R2108 VDD2.n60 VDD2.n6 10.4732
R2109 VDD2.n137 VDD2.n86 9.69747
R2110 VDD2.n117 VDD2.n96 9.69747
R2111 VDD2.n39 VDD2.n18 9.69747
R2112 VDD2.n59 VDD2.n8 9.69747
R2113 VDD2.n153 VDD2.n152 9.45567
R2114 VDD2.n76 VDD2.n75 9.45567
R2115 VDD2.n129 VDD2.n128 9.3005
R2116 VDD2.n88 VDD2.n87 9.3005
R2117 VDD2.n135 VDD2.n134 9.3005
R2118 VDD2.n137 VDD2.n136 9.3005
R2119 VDD2.n84 VDD2.n83 9.3005
R2120 VDD2.n143 VDD2.n142 9.3005
R2121 VDD2.n145 VDD2.n144 9.3005
R2122 VDD2.n81 VDD2.n78 9.3005
R2123 VDD2.n152 VDD2.n151 9.3005
R2124 VDD2.n127 VDD2.n126 9.3005
R2125 VDD2.n92 VDD2.n91 9.3005
R2126 VDD2.n121 VDD2.n120 9.3005
R2127 VDD2.n119 VDD2.n118 9.3005
R2128 VDD2.n96 VDD2.n95 9.3005
R2129 VDD2.n113 VDD2.n112 9.3005
R2130 VDD2.n111 VDD2.n110 9.3005
R2131 VDD2.n100 VDD2.n99 9.3005
R2132 VDD2.n105 VDD2.n104 9.3005
R2133 VDD2.n75 VDD2.n74 9.3005
R2134 VDD2.n14 VDD2.n13 9.3005
R2135 VDD2.n43 VDD2.n42 9.3005
R2136 VDD2.n41 VDD2.n40 9.3005
R2137 VDD2.n18 VDD2.n17 9.3005
R2138 VDD2.n35 VDD2.n34 9.3005
R2139 VDD2.n33 VDD2.n32 9.3005
R2140 VDD2.n22 VDD2.n21 9.3005
R2141 VDD2.n27 VDD2.n26 9.3005
R2142 VDD2.n49 VDD2.n48 9.3005
R2143 VDD2.n51 VDD2.n50 9.3005
R2144 VDD2.n10 VDD2.n9 9.3005
R2145 VDD2.n57 VDD2.n56 9.3005
R2146 VDD2.n59 VDD2.n58 9.3005
R2147 VDD2.n6 VDD2.n5 9.3005
R2148 VDD2.n65 VDD2.n64 9.3005
R2149 VDD2.n67 VDD2.n66 9.3005
R2150 VDD2.n68 VDD2.n1 9.3005
R2151 VDD2.n134 VDD2.n133 8.92171
R2152 VDD2.n118 VDD2.n94 8.92171
R2153 VDD2.n40 VDD2.n16 8.92171
R2154 VDD2.n56 VDD2.n55 8.92171
R2155 VDD2.n130 VDD2.n88 8.14595
R2156 VDD2.n122 VDD2.n121 8.14595
R2157 VDD2.n44 VDD2.n43 8.14595
R2158 VDD2.n52 VDD2.n10 8.14595
R2159 VDD2.n129 VDD2.n90 7.3702
R2160 VDD2.n125 VDD2.n92 7.3702
R2161 VDD2.n47 VDD2.n14 7.3702
R2162 VDD2.n51 VDD2.n12 7.3702
R2163 VDD2.n126 VDD2.n90 6.59444
R2164 VDD2.n126 VDD2.n125 6.59444
R2165 VDD2.n48 VDD2.n47 6.59444
R2166 VDD2.n48 VDD2.n12 6.59444
R2167 VDD2.n130 VDD2.n129 5.81868
R2168 VDD2.n122 VDD2.n92 5.81868
R2169 VDD2.n44 VDD2.n14 5.81868
R2170 VDD2.n52 VDD2.n51 5.81868
R2171 VDD2.n133 VDD2.n88 5.04292
R2172 VDD2.n121 VDD2.n94 5.04292
R2173 VDD2.n43 VDD2.n16 5.04292
R2174 VDD2.n55 VDD2.n10 5.04292
R2175 VDD2.n104 VDD2.n103 4.38563
R2176 VDD2.n26 VDD2.n25 4.38563
R2177 VDD2.n134 VDD2.n86 4.26717
R2178 VDD2.n118 VDD2.n117 4.26717
R2179 VDD2.n40 VDD2.n39 4.26717
R2180 VDD2.n56 VDD2.n8 4.26717
R2181 VDD2.n138 VDD2.n137 3.49141
R2182 VDD2.n114 VDD2.n96 3.49141
R2183 VDD2.n36 VDD2.n18 3.49141
R2184 VDD2.n60 VDD2.n59 3.49141
R2185 VDD2.n141 VDD2.n84 2.71565
R2186 VDD2.n113 VDD2.n98 2.71565
R2187 VDD2.n35 VDD2.n20 2.71565
R2188 VDD2.n63 VDD2.n6 2.71565
R2189 VDD2.n142 VDD2.n82 1.93989
R2190 VDD2.n110 VDD2.n109 1.93989
R2191 VDD2.n32 VDD2.n31 1.93989
R2192 VDD2.n64 VDD2.n4 1.93989
R2193 VDD2.n153 VDD2.n77 1.16414
R2194 VDD2.n146 VDD2.n145 1.16414
R2195 VDD2.n106 VDD2.n100 1.16414
R2196 VDD2.n28 VDD2.n22 1.16414
R2197 VDD2.n69 VDD2.n67 1.16414
R2198 VDD2.n76 VDD2.n0 1.16414
R2199 VDD2 VDD2.n154 0.597483
R2200 VDD2.n151 VDD2.n150 0.388379
R2201 VDD2.n81 VDD2.n79 0.388379
R2202 VDD2.n105 VDD2.n102 0.388379
R2203 VDD2.n27 VDD2.n24 0.388379
R2204 VDD2.n68 VDD2.n2 0.388379
R2205 VDD2.n74 VDD2.n73 0.388379
R2206 VDD2.n152 VDD2.n78 0.155672
R2207 VDD2.n144 VDD2.n78 0.155672
R2208 VDD2.n144 VDD2.n143 0.155672
R2209 VDD2.n143 VDD2.n83 0.155672
R2210 VDD2.n136 VDD2.n83 0.155672
R2211 VDD2.n136 VDD2.n135 0.155672
R2212 VDD2.n135 VDD2.n87 0.155672
R2213 VDD2.n128 VDD2.n87 0.155672
R2214 VDD2.n128 VDD2.n127 0.155672
R2215 VDD2.n127 VDD2.n91 0.155672
R2216 VDD2.n120 VDD2.n91 0.155672
R2217 VDD2.n120 VDD2.n119 0.155672
R2218 VDD2.n119 VDD2.n95 0.155672
R2219 VDD2.n112 VDD2.n95 0.155672
R2220 VDD2.n112 VDD2.n111 0.155672
R2221 VDD2.n111 VDD2.n99 0.155672
R2222 VDD2.n104 VDD2.n99 0.155672
R2223 VDD2.n26 VDD2.n21 0.155672
R2224 VDD2.n33 VDD2.n21 0.155672
R2225 VDD2.n34 VDD2.n33 0.155672
R2226 VDD2.n34 VDD2.n17 0.155672
R2227 VDD2.n41 VDD2.n17 0.155672
R2228 VDD2.n42 VDD2.n41 0.155672
R2229 VDD2.n42 VDD2.n13 0.155672
R2230 VDD2.n49 VDD2.n13 0.155672
R2231 VDD2.n50 VDD2.n49 0.155672
R2232 VDD2.n50 VDD2.n9 0.155672
R2233 VDD2.n57 VDD2.n9 0.155672
R2234 VDD2.n58 VDD2.n57 0.155672
R2235 VDD2.n58 VDD2.n5 0.155672
R2236 VDD2.n65 VDD2.n5 0.155672
R2237 VDD2.n66 VDD2.n65 0.155672
R2238 VDD2.n66 VDD2.n1 0.155672
R2239 VDD2.n75 VDD2.n1 0.155672
C0 VN VP 5.62474f
C1 VDD2 VTAIL 5.61809f
C2 VTAIL VP 2.65877f
C3 VDD2 VDD1 0.623607f
C4 VN VTAIL 2.6444f
C5 VDD1 VP 3.27056f
C6 VN VDD1 0.148259f
C7 VDD2 VP 0.315546f
C8 VTAIL VDD1 5.57144f
C9 VDD2 VN 3.10645f
C10 VDD2 B 4.638935f
C11 VDD1 B 7.46102f
C12 VTAIL B 7.955455f
C13 VN B 10.776061f
C14 VP B 6.013072f
C15 VDD2.n0 B 0.025997f
C16 VDD2.n1 B 0.020034f
C17 VDD2.n2 B 0.011082f
C18 VDD2.n3 B 0.025445f
C19 VDD2.n4 B 0.011398f
C20 VDD2.n5 B 0.020034f
C21 VDD2.n6 B 0.010765f
C22 VDD2.n7 B 0.025445f
C23 VDD2.n8 B 0.011398f
C24 VDD2.n9 B 0.020034f
C25 VDD2.n10 B 0.010765f
C26 VDD2.n11 B 0.025445f
C27 VDD2.n12 B 0.011398f
C28 VDD2.n13 B 0.020034f
C29 VDD2.n14 B 0.010765f
C30 VDD2.n15 B 0.025445f
C31 VDD2.n16 B 0.011398f
C32 VDD2.n17 B 0.020034f
C33 VDD2.n18 B 0.010765f
C34 VDD2.n19 B 0.025445f
C35 VDD2.n20 B 0.011398f
C36 VDD2.n21 B 0.020034f
C37 VDD2.n22 B 0.010765f
C38 VDD2.n23 B 0.019084f
C39 VDD2.n24 B 0.015031f
C40 VDD2.t0 B 0.041887f
C41 VDD2.n25 B 0.125642f
C42 VDD2.n26 B 1.21161f
C43 VDD2.n27 B 0.010765f
C44 VDD2.n28 B 0.011398f
C45 VDD2.n29 B 0.025445f
C46 VDD2.n30 B 0.025445f
C47 VDD2.n31 B 0.011398f
C48 VDD2.n32 B 0.010765f
C49 VDD2.n33 B 0.020034f
C50 VDD2.n34 B 0.020034f
C51 VDD2.n35 B 0.010765f
C52 VDD2.n36 B 0.011398f
C53 VDD2.n37 B 0.025445f
C54 VDD2.n38 B 0.025445f
C55 VDD2.n39 B 0.011398f
C56 VDD2.n40 B 0.010765f
C57 VDD2.n41 B 0.020034f
C58 VDD2.n42 B 0.020034f
C59 VDD2.n43 B 0.010765f
C60 VDD2.n44 B 0.011398f
C61 VDD2.n45 B 0.025445f
C62 VDD2.n46 B 0.025445f
C63 VDD2.n47 B 0.011398f
C64 VDD2.n48 B 0.010765f
C65 VDD2.n49 B 0.020034f
C66 VDD2.n50 B 0.020034f
C67 VDD2.n51 B 0.010765f
C68 VDD2.n52 B 0.011398f
C69 VDD2.n53 B 0.025445f
C70 VDD2.n54 B 0.025445f
C71 VDD2.n55 B 0.011398f
C72 VDD2.n56 B 0.010765f
C73 VDD2.n57 B 0.020034f
C74 VDD2.n58 B 0.020034f
C75 VDD2.n59 B 0.010765f
C76 VDD2.n60 B 0.011398f
C77 VDD2.n61 B 0.025445f
C78 VDD2.n62 B 0.025445f
C79 VDD2.n63 B 0.011398f
C80 VDD2.n64 B 0.010765f
C81 VDD2.n65 B 0.020034f
C82 VDD2.n66 B 0.020034f
C83 VDD2.n67 B 0.010765f
C84 VDD2.n68 B 0.010765f
C85 VDD2.n69 B 0.011398f
C86 VDD2.n70 B 0.025445f
C87 VDD2.n71 B 0.025445f
C88 VDD2.n72 B 0.05126f
C89 VDD2.n73 B 0.011082f
C90 VDD2.n74 B 0.010765f
C91 VDD2.n75 B 0.048497f
C92 VDD2.n76 B 0.61187f
C93 VDD2.n77 B 0.025997f
C94 VDD2.n78 B 0.020034f
C95 VDD2.n79 B 0.011082f
C96 VDD2.n80 B 0.025445f
C97 VDD2.n81 B 0.010765f
C98 VDD2.n82 B 0.011398f
C99 VDD2.n83 B 0.020034f
C100 VDD2.n84 B 0.010765f
C101 VDD2.n85 B 0.025445f
C102 VDD2.n86 B 0.011398f
C103 VDD2.n87 B 0.020034f
C104 VDD2.n88 B 0.010765f
C105 VDD2.n89 B 0.025445f
C106 VDD2.n90 B 0.011398f
C107 VDD2.n91 B 0.020034f
C108 VDD2.n92 B 0.010765f
C109 VDD2.n93 B 0.025445f
C110 VDD2.n94 B 0.011398f
C111 VDD2.n95 B 0.020034f
C112 VDD2.n96 B 0.010765f
C113 VDD2.n97 B 0.025445f
C114 VDD2.n98 B 0.011398f
C115 VDD2.n99 B 0.020034f
C116 VDD2.n100 B 0.010765f
C117 VDD2.n101 B 0.019084f
C118 VDD2.n102 B 0.015031f
C119 VDD2.t1 B 0.041887f
C120 VDD2.n103 B 0.125642f
C121 VDD2.n104 B 1.21161f
C122 VDD2.n105 B 0.010765f
C123 VDD2.n106 B 0.011398f
C124 VDD2.n107 B 0.025445f
C125 VDD2.n108 B 0.025445f
C126 VDD2.n109 B 0.011398f
C127 VDD2.n110 B 0.010765f
C128 VDD2.n111 B 0.020034f
C129 VDD2.n112 B 0.020034f
C130 VDD2.n113 B 0.010765f
C131 VDD2.n114 B 0.011398f
C132 VDD2.n115 B 0.025445f
C133 VDD2.n116 B 0.025445f
C134 VDD2.n117 B 0.011398f
C135 VDD2.n118 B 0.010765f
C136 VDD2.n119 B 0.020034f
C137 VDD2.n120 B 0.020034f
C138 VDD2.n121 B 0.010765f
C139 VDD2.n122 B 0.011398f
C140 VDD2.n123 B 0.025445f
C141 VDD2.n124 B 0.025445f
C142 VDD2.n125 B 0.011398f
C143 VDD2.n126 B 0.010765f
C144 VDD2.n127 B 0.020034f
C145 VDD2.n128 B 0.020034f
C146 VDD2.n129 B 0.010765f
C147 VDD2.n130 B 0.011398f
C148 VDD2.n131 B 0.025445f
C149 VDD2.n132 B 0.025445f
C150 VDD2.n133 B 0.011398f
C151 VDD2.n134 B 0.010765f
C152 VDD2.n135 B 0.020034f
C153 VDD2.n136 B 0.020034f
C154 VDD2.n137 B 0.010765f
C155 VDD2.n138 B 0.011398f
C156 VDD2.n139 B 0.025445f
C157 VDD2.n140 B 0.025445f
C158 VDD2.n141 B 0.011398f
C159 VDD2.n142 B 0.010765f
C160 VDD2.n143 B 0.020034f
C161 VDD2.n144 B 0.020034f
C162 VDD2.n145 B 0.010765f
C163 VDD2.n146 B 0.011398f
C164 VDD2.n147 B 0.025445f
C165 VDD2.n148 B 0.025445f
C166 VDD2.n149 B 0.05126f
C167 VDD2.n150 B 0.011082f
C168 VDD2.n151 B 0.010765f
C169 VDD2.n152 B 0.048497f
C170 VDD2.n153 B 0.042171f
C171 VDD2.n154 B 2.55644f
C172 VN.t1 B 3.06086f
C173 VN.t0 B 3.52266f
C174 VDD1.n0 B 0.02637f
C175 VDD1.n1 B 0.020321f
C176 VDD1.n2 B 0.011241f
C177 VDD1.n3 B 0.025811f
C178 VDD1.n4 B 0.01092f
C179 VDD1.n5 B 0.011562f
C180 VDD1.n6 B 0.020321f
C181 VDD1.n7 B 0.01092f
C182 VDD1.n8 B 0.025811f
C183 VDD1.n9 B 0.011562f
C184 VDD1.n10 B 0.020321f
C185 VDD1.n11 B 0.01092f
C186 VDD1.n12 B 0.025811f
C187 VDD1.n13 B 0.011562f
C188 VDD1.n14 B 0.020321f
C189 VDD1.n15 B 0.01092f
C190 VDD1.n16 B 0.025811f
C191 VDD1.n17 B 0.011562f
C192 VDD1.n18 B 0.020321f
C193 VDD1.n19 B 0.01092f
C194 VDD1.n20 B 0.025811f
C195 VDD1.n21 B 0.011562f
C196 VDD1.n22 B 0.020321f
C197 VDD1.n23 B 0.01092f
C198 VDD1.n24 B 0.019358f
C199 VDD1.n25 B 0.015247f
C200 VDD1.t1 B 0.042489f
C201 VDD1.n26 B 0.127446f
C202 VDD1.n27 B 1.22901f
C203 VDD1.n28 B 0.01092f
C204 VDD1.n29 B 0.011562f
C205 VDD1.n30 B 0.025811f
C206 VDD1.n31 B 0.025811f
C207 VDD1.n32 B 0.011562f
C208 VDD1.n33 B 0.01092f
C209 VDD1.n34 B 0.020321f
C210 VDD1.n35 B 0.020321f
C211 VDD1.n36 B 0.01092f
C212 VDD1.n37 B 0.011562f
C213 VDD1.n38 B 0.025811f
C214 VDD1.n39 B 0.025811f
C215 VDD1.n40 B 0.011562f
C216 VDD1.n41 B 0.01092f
C217 VDD1.n42 B 0.020321f
C218 VDD1.n43 B 0.020321f
C219 VDD1.n44 B 0.01092f
C220 VDD1.n45 B 0.011562f
C221 VDD1.n46 B 0.025811f
C222 VDD1.n47 B 0.025811f
C223 VDD1.n48 B 0.011562f
C224 VDD1.n49 B 0.01092f
C225 VDD1.n50 B 0.020321f
C226 VDD1.n51 B 0.020321f
C227 VDD1.n52 B 0.01092f
C228 VDD1.n53 B 0.011562f
C229 VDD1.n54 B 0.025811f
C230 VDD1.n55 B 0.025811f
C231 VDD1.n56 B 0.011562f
C232 VDD1.n57 B 0.01092f
C233 VDD1.n58 B 0.020321f
C234 VDD1.n59 B 0.020321f
C235 VDD1.n60 B 0.01092f
C236 VDD1.n61 B 0.011562f
C237 VDD1.n62 B 0.025811f
C238 VDD1.n63 B 0.025811f
C239 VDD1.n64 B 0.011562f
C240 VDD1.n65 B 0.01092f
C241 VDD1.n66 B 0.020321f
C242 VDD1.n67 B 0.020321f
C243 VDD1.n68 B 0.01092f
C244 VDD1.n69 B 0.011562f
C245 VDD1.n70 B 0.025811f
C246 VDD1.n71 B 0.025811f
C247 VDD1.n72 B 0.051996f
C248 VDD1.n73 B 0.011241f
C249 VDD1.n74 B 0.01092f
C250 VDD1.n75 B 0.049193f
C251 VDD1.n76 B 0.043707f
C252 VDD1.n77 B 0.02637f
C253 VDD1.n78 B 0.020321f
C254 VDD1.n79 B 0.011241f
C255 VDD1.n80 B 0.025811f
C256 VDD1.n81 B 0.011562f
C257 VDD1.n82 B 0.020321f
C258 VDD1.n83 B 0.01092f
C259 VDD1.n84 B 0.025811f
C260 VDD1.n85 B 0.011562f
C261 VDD1.n86 B 0.020321f
C262 VDD1.n87 B 0.01092f
C263 VDD1.n88 B 0.025811f
C264 VDD1.n89 B 0.011562f
C265 VDD1.n90 B 0.020321f
C266 VDD1.n91 B 0.01092f
C267 VDD1.n92 B 0.025811f
C268 VDD1.n93 B 0.011562f
C269 VDD1.n94 B 0.020321f
C270 VDD1.n95 B 0.01092f
C271 VDD1.n96 B 0.025811f
C272 VDD1.n97 B 0.011562f
C273 VDD1.n98 B 0.020321f
C274 VDD1.n99 B 0.01092f
C275 VDD1.n100 B 0.019358f
C276 VDD1.n101 B 0.015247f
C277 VDD1.t0 B 0.042489f
C278 VDD1.n102 B 0.127446f
C279 VDD1.n103 B 1.22901f
C280 VDD1.n104 B 0.01092f
C281 VDD1.n105 B 0.011562f
C282 VDD1.n106 B 0.025811f
C283 VDD1.n107 B 0.025811f
C284 VDD1.n108 B 0.011562f
C285 VDD1.n109 B 0.01092f
C286 VDD1.n110 B 0.020321f
C287 VDD1.n111 B 0.020321f
C288 VDD1.n112 B 0.01092f
C289 VDD1.n113 B 0.011562f
C290 VDD1.n114 B 0.025811f
C291 VDD1.n115 B 0.025811f
C292 VDD1.n116 B 0.011562f
C293 VDD1.n117 B 0.01092f
C294 VDD1.n118 B 0.020321f
C295 VDD1.n119 B 0.020321f
C296 VDD1.n120 B 0.01092f
C297 VDD1.n121 B 0.011562f
C298 VDD1.n122 B 0.025811f
C299 VDD1.n123 B 0.025811f
C300 VDD1.n124 B 0.011562f
C301 VDD1.n125 B 0.01092f
C302 VDD1.n126 B 0.020321f
C303 VDD1.n127 B 0.020321f
C304 VDD1.n128 B 0.01092f
C305 VDD1.n129 B 0.011562f
C306 VDD1.n130 B 0.025811f
C307 VDD1.n131 B 0.025811f
C308 VDD1.n132 B 0.011562f
C309 VDD1.n133 B 0.01092f
C310 VDD1.n134 B 0.020321f
C311 VDD1.n135 B 0.020321f
C312 VDD1.n136 B 0.01092f
C313 VDD1.n137 B 0.011562f
C314 VDD1.n138 B 0.025811f
C315 VDD1.n139 B 0.025811f
C316 VDD1.n140 B 0.011562f
C317 VDD1.n141 B 0.01092f
C318 VDD1.n142 B 0.020321f
C319 VDD1.n143 B 0.020321f
C320 VDD1.n144 B 0.01092f
C321 VDD1.n145 B 0.01092f
C322 VDD1.n146 B 0.011562f
C323 VDD1.n147 B 0.025811f
C324 VDD1.n148 B 0.025811f
C325 VDD1.n149 B 0.051996f
C326 VDD1.n150 B 0.011241f
C327 VDD1.n151 B 0.01092f
C328 VDD1.n152 B 0.049193f
C329 VDD1.n153 B 0.658228f
C330 VTAIL.n0 B 0.026175f
C331 VTAIL.n1 B 0.020171f
C332 VTAIL.n2 B 0.011158f
C333 VTAIL.n3 B 0.025619f
C334 VTAIL.n4 B 0.011477f
C335 VTAIL.n5 B 0.020171f
C336 VTAIL.n6 B 0.010839f
C337 VTAIL.n7 B 0.025619f
C338 VTAIL.n8 B 0.011477f
C339 VTAIL.n9 B 0.020171f
C340 VTAIL.n10 B 0.010839f
C341 VTAIL.n11 B 0.025619f
C342 VTAIL.n12 B 0.011477f
C343 VTAIL.n13 B 0.020171f
C344 VTAIL.n14 B 0.010839f
C345 VTAIL.n15 B 0.025619f
C346 VTAIL.n16 B 0.011477f
C347 VTAIL.n17 B 0.020171f
C348 VTAIL.n18 B 0.010839f
C349 VTAIL.n19 B 0.025619f
C350 VTAIL.n20 B 0.011477f
C351 VTAIL.n21 B 0.020171f
C352 VTAIL.n22 B 0.010839f
C353 VTAIL.n23 B 0.019215f
C354 VTAIL.n24 B 0.015134f
C355 VTAIL.t3 B 0.042174f
C356 VTAIL.n25 B 0.126502f
C357 VTAIL.n26 B 1.21991f
C358 VTAIL.n27 B 0.010839f
C359 VTAIL.n28 B 0.011477f
C360 VTAIL.n29 B 0.025619f
C361 VTAIL.n30 B 0.025619f
C362 VTAIL.n31 B 0.011477f
C363 VTAIL.n32 B 0.010839f
C364 VTAIL.n33 B 0.020171f
C365 VTAIL.n34 B 0.020171f
C366 VTAIL.n35 B 0.010839f
C367 VTAIL.n36 B 0.011477f
C368 VTAIL.n37 B 0.025619f
C369 VTAIL.n38 B 0.025619f
C370 VTAIL.n39 B 0.011477f
C371 VTAIL.n40 B 0.010839f
C372 VTAIL.n41 B 0.020171f
C373 VTAIL.n42 B 0.020171f
C374 VTAIL.n43 B 0.010839f
C375 VTAIL.n44 B 0.011477f
C376 VTAIL.n45 B 0.025619f
C377 VTAIL.n46 B 0.025619f
C378 VTAIL.n47 B 0.011477f
C379 VTAIL.n48 B 0.010839f
C380 VTAIL.n49 B 0.020171f
C381 VTAIL.n50 B 0.020171f
C382 VTAIL.n51 B 0.010839f
C383 VTAIL.n52 B 0.011477f
C384 VTAIL.n53 B 0.025619f
C385 VTAIL.n54 B 0.025619f
C386 VTAIL.n55 B 0.011477f
C387 VTAIL.n56 B 0.010839f
C388 VTAIL.n57 B 0.020171f
C389 VTAIL.n58 B 0.020171f
C390 VTAIL.n59 B 0.010839f
C391 VTAIL.n60 B 0.011477f
C392 VTAIL.n61 B 0.025619f
C393 VTAIL.n62 B 0.025619f
C394 VTAIL.n63 B 0.011477f
C395 VTAIL.n64 B 0.010839f
C396 VTAIL.n65 B 0.020171f
C397 VTAIL.n66 B 0.020171f
C398 VTAIL.n67 B 0.010839f
C399 VTAIL.n68 B 0.010839f
C400 VTAIL.n69 B 0.011477f
C401 VTAIL.n70 B 0.025619f
C402 VTAIL.n71 B 0.025619f
C403 VTAIL.n72 B 0.051611f
C404 VTAIL.n73 B 0.011158f
C405 VTAIL.n74 B 0.010839f
C406 VTAIL.n75 B 0.048829f
C407 VTAIL.n76 B 0.028549f
C408 VTAIL.n77 B 1.42639f
C409 VTAIL.n78 B 0.026175f
C410 VTAIL.n79 B 0.020171f
C411 VTAIL.n80 B 0.011158f
C412 VTAIL.n81 B 0.025619f
C413 VTAIL.n82 B 0.010839f
C414 VTAIL.n83 B 0.011477f
C415 VTAIL.n84 B 0.020171f
C416 VTAIL.n85 B 0.010839f
C417 VTAIL.n86 B 0.025619f
C418 VTAIL.n87 B 0.011477f
C419 VTAIL.n88 B 0.020171f
C420 VTAIL.n89 B 0.010839f
C421 VTAIL.n90 B 0.025619f
C422 VTAIL.n91 B 0.011477f
C423 VTAIL.n92 B 0.020171f
C424 VTAIL.n93 B 0.010839f
C425 VTAIL.n94 B 0.025619f
C426 VTAIL.n95 B 0.011477f
C427 VTAIL.n96 B 0.020171f
C428 VTAIL.n97 B 0.010839f
C429 VTAIL.n98 B 0.025619f
C430 VTAIL.n99 B 0.011477f
C431 VTAIL.n100 B 0.020171f
C432 VTAIL.n101 B 0.010839f
C433 VTAIL.n102 B 0.019215f
C434 VTAIL.n103 B 0.015134f
C435 VTAIL.t0 B 0.042174f
C436 VTAIL.n104 B 0.126502f
C437 VTAIL.n105 B 1.21991f
C438 VTAIL.n106 B 0.010839f
C439 VTAIL.n107 B 0.011477f
C440 VTAIL.n108 B 0.025619f
C441 VTAIL.n109 B 0.025619f
C442 VTAIL.n110 B 0.011477f
C443 VTAIL.n111 B 0.010839f
C444 VTAIL.n112 B 0.020171f
C445 VTAIL.n113 B 0.020171f
C446 VTAIL.n114 B 0.010839f
C447 VTAIL.n115 B 0.011477f
C448 VTAIL.n116 B 0.025619f
C449 VTAIL.n117 B 0.025619f
C450 VTAIL.n118 B 0.011477f
C451 VTAIL.n119 B 0.010839f
C452 VTAIL.n120 B 0.020171f
C453 VTAIL.n121 B 0.020171f
C454 VTAIL.n122 B 0.010839f
C455 VTAIL.n123 B 0.011477f
C456 VTAIL.n124 B 0.025619f
C457 VTAIL.n125 B 0.025619f
C458 VTAIL.n126 B 0.011477f
C459 VTAIL.n127 B 0.010839f
C460 VTAIL.n128 B 0.020171f
C461 VTAIL.n129 B 0.020171f
C462 VTAIL.n130 B 0.010839f
C463 VTAIL.n131 B 0.011477f
C464 VTAIL.n132 B 0.025619f
C465 VTAIL.n133 B 0.025619f
C466 VTAIL.n134 B 0.011477f
C467 VTAIL.n135 B 0.010839f
C468 VTAIL.n136 B 0.020171f
C469 VTAIL.n137 B 0.020171f
C470 VTAIL.n138 B 0.010839f
C471 VTAIL.n139 B 0.011477f
C472 VTAIL.n140 B 0.025619f
C473 VTAIL.n141 B 0.025619f
C474 VTAIL.n142 B 0.011477f
C475 VTAIL.n143 B 0.010839f
C476 VTAIL.n144 B 0.020171f
C477 VTAIL.n145 B 0.020171f
C478 VTAIL.n146 B 0.010839f
C479 VTAIL.n147 B 0.011477f
C480 VTAIL.n148 B 0.025619f
C481 VTAIL.n149 B 0.025619f
C482 VTAIL.n150 B 0.051611f
C483 VTAIL.n151 B 0.011158f
C484 VTAIL.n152 B 0.010839f
C485 VTAIL.n153 B 0.048829f
C486 VTAIL.n154 B 0.028549f
C487 VTAIL.n155 B 1.45763f
C488 VTAIL.n156 B 0.026175f
C489 VTAIL.n157 B 0.020171f
C490 VTAIL.n158 B 0.011158f
C491 VTAIL.n159 B 0.025619f
C492 VTAIL.n160 B 0.010839f
C493 VTAIL.n161 B 0.011477f
C494 VTAIL.n162 B 0.020171f
C495 VTAIL.n163 B 0.010839f
C496 VTAIL.n164 B 0.025619f
C497 VTAIL.n165 B 0.011477f
C498 VTAIL.n166 B 0.020171f
C499 VTAIL.n167 B 0.010839f
C500 VTAIL.n168 B 0.025619f
C501 VTAIL.n169 B 0.011477f
C502 VTAIL.n170 B 0.020171f
C503 VTAIL.n171 B 0.010839f
C504 VTAIL.n172 B 0.025619f
C505 VTAIL.n173 B 0.011477f
C506 VTAIL.n174 B 0.020171f
C507 VTAIL.n175 B 0.010839f
C508 VTAIL.n176 B 0.025619f
C509 VTAIL.n177 B 0.011477f
C510 VTAIL.n178 B 0.020171f
C511 VTAIL.n179 B 0.010839f
C512 VTAIL.n180 B 0.019215f
C513 VTAIL.n181 B 0.015134f
C514 VTAIL.t2 B 0.042174f
C515 VTAIL.n182 B 0.126502f
C516 VTAIL.n183 B 1.21991f
C517 VTAIL.n184 B 0.010839f
C518 VTAIL.n185 B 0.011477f
C519 VTAIL.n186 B 0.025619f
C520 VTAIL.n187 B 0.025619f
C521 VTAIL.n188 B 0.011477f
C522 VTAIL.n189 B 0.010839f
C523 VTAIL.n190 B 0.020171f
C524 VTAIL.n191 B 0.020171f
C525 VTAIL.n192 B 0.010839f
C526 VTAIL.n193 B 0.011477f
C527 VTAIL.n194 B 0.025619f
C528 VTAIL.n195 B 0.025619f
C529 VTAIL.n196 B 0.011477f
C530 VTAIL.n197 B 0.010839f
C531 VTAIL.n198 B 0.020171f
C532 VTAIL.n199 B 0.020171f
C533 VTAIL.n200 B 0.010839f
C534 VTAIL.n201 B 0.011477f
C535 VTAIL.n202 B 0.025619f
C536 VTAIL.n203 B 0.025619f
C537 VTAIL.n204 B 0.011477f
C538 VTAIL.n205 B 0.010839f
C539 VTAIL.n206 B 0.020171f
C540 VTAIL.n207 B 0.020171f
C541 VTAIL.n208 B 0.010839f
C542 VTAIL.n209 B 0.011477f
C543 VTAIL.n210 B 0.025619f
C544 VTAIL.n211 B 0.025619f
C545 VTAIL.n212 B 0.011477f
C546 VTAIL.n213 B 0.010839f
C547 VTAIL.n214 B 0.020171f
C548 VTAIL.n215 B 0.020171f
C549 VTAIL.n216 B 0.010839f
C550 VTAIL.n217 B 0.011477f
C551 VTAIL.n218 B 0.025619f
C552 VTAIL.n219 B 0.025619f
C553 VTAIL.n220 B 0.011477f
C554 VTAIL.n221 B 0.010839f
C555 VTAIL.n222 B 0.020171f
C556 VTAIL.n223 B 0.020171f
C557 VTAIL.n224 B 0.010839f
C558 VTAIL.n225 B 0.011477f
C559 VTAIL.n226 B 0.025619f
C560 VTAIL.n227 B 0.025619f
C561 VTAIL.n228 B 0.051611f
C562 VTAIL.n229 B 0.011158f
C563 VTAIL.n230 B 0.010839f
C564 VTAIL.n231 B 0.048829f
C565 VTAIL.n232 B 0.028549f
C566 VTAIL.n233 B 1.31755f
C567 VTAIL.n234 B 0.026175f
C568 VTAIL.n235 B 0.020171f
C569 VTAIL.n236 B 0.011158f
C570 VTAIL.n237 B 0.025619f
C571 VTAIL.n238 B 0.011477f
C572 VTAIL.n239 B 0.020171f
C573 VTAIL.n240 B 0.010839f
C574 VTAIL.n241 B 0.025619f
C575 VTAIL.n242 B 0.011477f
C576 VTAIL.n243 B 0.020171f
C577 VTAIL.n244 B 0.010839f
C578 VTAIL.n245 B 0.025619f
C579 VTAIL.n246 B 0.011477f
C580 VTAIL.n247 B 0.020171f
C581 VTAIL.n248 B 0.010839f
C582 VTAIL.n249 B 0.025619f
C583 VTAIL.n250 B 0.011477f
C584 VTAIL.n251 B 0.020171f
C585 VTAIL.n252 B 0.010839f
C586 VTAIL.n253 B 0.025619f
C587 VTAIL.n254 B 0.011477f
C588 VTAIL.n255 B 0.020171f
C589 VTAIL.n256 B 0.010839f
C590 VTAIL.n257 B 0.019215f
C591 VTAIL.n258 B 0.015134f
C592 VTAIL.t1 B 0.042174f
C593 VTAIL.n259 B 0.126502f
C594 VTAIL.n260 B 1.21991f
C595 VTAIL.n261 B 0.010839f
C596 VTAIL.n262 B 0.011477f
C597 VTAIL.n263 B 0.025619f
C598 VTAIL.n264 B 0.025619f
C599 VTAIL.n265 B 0.011477f
C600 VTAIL.n266 B 0.010839f
C601 VTAIL.n267 B 0.020171f
C602 VTAIL.n268 B 0.020171f
C603 VTAIL.n269 B 0.010839f
C604 VTAIL.n270 B 0.011477f
C605 VTAIL.n271 B 0.025619f
C606 VTAIL.n272 B 0.025619f
C607 VTAIL.n273 B 0.011477f
C608 VTAIL.n274 B 0.010839f
C609 VTAIL.n275 B 0.020171f
C610 VTAIL.n276 B 0.020171f
C611 VTAIL.n277 B 0.010839f
C612 VTAIL.n278 B 0.011477f
C613 VTAIL.n279 B 0.025619f
C614 VTAIL.n280 B 0.025619f
C615 VTAIL.n281 B 0.011477f
C616 VTAIL.n282 B 0.010839f
C617 VTAIL.n283 B 0.020171f
C618 VTAIL.n284 B 0.020171f
C619 VTAIL.n285 B 0.010839f
C620 VTAIL.n286 B 0.011477f
C621 VTAIL.n287 B 0.025619f
C622 VTAIL.n288 B 0.025619f
C623 VTAIL.n289 B 0.011477f
C624 VTAIL.n290 B 0.010839f
C625 VTAIL.n291 B 0.020171f
C626 VTAIL.n292 B 0.020171f
C627 VTAIL.n293 B 0.010839f
C628 VTAIL.n294 B 0.011477f
C629 VTAIL.n295 B 0.025619f
C630 VTAIL.n296 B 0.025619f
C631 VTAIL.n297 B 0.011477f
C632 VTAIL.n298 B 0.010839f
C633 VTAIL.n299 B 0.020171f
C634 VTAIL.n300 B 0.020171f
C635 VTAIL.n301 B 0.010839f
C636 VTAIL.n302 B 0.010839f
C637 VTAIL.n303 B 0.011477f
C638 VTAIL.n304 B 0.025619f
C639 VTAIL.n305 B 0.025619f
C640 VTAIL.n306 B 0.051611f
C641 VTAIL.n307 B 0.011158f
C642 VTAIL.n308 B 0.010839f
C643 VTAIL.n309 B 0.048829f
C644 VTAIL.n310 B 0.028549f
C645 VTAIL.n311 B 1.24821f
C646 VP.t0 B 3.62827f
C647 VP.t1 B 3.15354f
C648 VP.n0 B 4.74937f
.ends

