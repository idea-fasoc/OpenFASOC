* NGSPICE file created from diff_pair_sample_1618.ext - technology: sky130A

.subckt diff_pair_sample_1618 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.5054 pd=8.5 as=1.5054 ps=8.5 w=3.86 l=0.37
X1 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.5054 pd=8.5 as=1.5054 ps=8.5 w=3.86 l=0.37
X2 VDD1.t0 VP.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.5054 pd=8.5 as=1.5054 ps=8.5 w=3.86 l=0.37
X3 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=1.5054 pd=8.5 as=0 ps=0 w=3.86 l=0.37
X4 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5054 pd=8.5 as=0 ps=0 w=3.86 l=0.37
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.5054 pd=8.5 as=0 ps=0 w=3.86 l=0.37
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5054 pd=8.5 as=0 ps=0 w=3.86 l=0.37
X7 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.5054 pd=8.5 as=1.5054 ps=8.5 w=3.86 l=0.37
R0 VP.n0 VP.t1 551.484
R1 VP.n0 VP.t0 518.893
R2 VP VP.n0 0.0516364
R3 VTAIL.n74 VTAIL.n60 289.615
R4 VTAIL.n14 VTAIL.n0 289.615
R5 VTAIL.n54 VTAIL.n40 289.615
R6 VTAIL.n34 VTAIL.n20 289.615
R7 VTAIL.n67 VTAIL.n66 185
R8 VTAIL.n64 VTAIL.n63 185
R9 VTAIL.n73 VTAIL.n72 185
R10 VTAIL.n75 VTAIL.n74 185
R11 VTAIL.n7 VTAIL.n6 185
R12 VTAIL.n4 VTAIL.n3 185
R13 VTAIL.n13 VTAIL.n12 185
R14 VTAIL.n15 VTAIL.n14 185
R15 VTAIL.n55 VTAIL.n54 185
R16 VTAIL.n53 VTAIL.n52 185
R17 VTAIL.n44 VTAIL.n43 185
R18 VTAIL.n47 VTAIL.n46 185
R19 VTAIL.n35 VTAIL.n34 185
R20 VTAIL.n33 VTAIL.n32 185
R21 VTAIL.n24 VTAIL.n23 185
R22 VTAIL.n27 VTAIL.n26 185
R23 VTAIL.t0 VTAIL.n65 147.888
R24 VTAIL.t3 VTAIL.n5 147.888
R25 VTAIL.t2 VTAIL.n45 147.888
R26 VTAIL.t1 VTAIL.n25 147.888
R27 VTAIL.n66 VTAIL.n63 104.615
R28 VTAIL.n73 VTAIL.n63 104.615
R29 VTAIL.n74 VTAIL.n73 104.615
R30 VTAIL.n6 VTAIL.n3 104.615
R31 VTAIL.n13 VTAIL.n3 104.615
R32 VTAIL.n14 VTAIL.n13 104.615
R33 VTAIL.n54 VTAIL.n53 104.615
R34 VTAIL.n53 VTAIL.n43 104.615
R35 VTAIL.n46 VTAIL.n43 104.615
R36 VTAIL.n34 VTAIL.n33 104.615
R37 VTAIL.n33 VTAIL.n23 104.615
R38 VTAIL.n26 VTAIL.n23 104.615
R39 VTAIL.n66 VTAIL.t0 52.3082
R40 VTAIL.n6 VTAIL.t3 52.3082
R41 VTAIL.n46 VTAIL.t2 52.3082
R42 VTAIL.n26 VTAIL.t1 52.3082
R43 VTAIL.n79 VTAIL.n78 32.5732
R44 VTAIL.n19 VTAIL.n18 32.5732
R45 VTAIL.n59 VTAIL.n58 32.5732
R46 VTAIL.n39 VTAIL.n38 32.5732
R47 VTAIL.n39 VTAIL.n19 16.9186
R48 VTAIL.n79 VTAIL.n59 16.3152
R49 VTAIL.n67 VTAIL.n65 15.6496
R50 VTAIL.n7 VTAIL.n5 15.6496
R51 VTAIL.n47 VTAIL.n45 15.6496
R52 VTAIL.n27 VTAIL.n25 15.6496
R53 VTAIL.n68 VTAIL.n64 12.8005
R54 VTAIL.n8 VTAIL.n4 12.8005
R55 VTAIL.n48 VTAIL.n44 12.8005
R56 VTAIL.n28 VTAIL.n24 12.8005
R57 VTAIL.n72 VTAIL.n71 12.0247
R58 VTAIL.n12 VTAIL.n11 12.0247
R59 VTAIL.n52 VTAIL.n51 12.0247
R60 VTAIL.n32 VTAIL.n31 12.0247
R61 VTAIL.n75 VTAIL.n62 11.249
R62 VTAIL.n15 VTAIL.n2 11.249
R63 VTAIL.n55 VTAIL.n42 11.249
R64 VTAIL.n35 VTAIL.n22 11.249
R65 VTAIL.n76 VTAIL.n60 10.4732
R66 VTAIL.n16 VTAIL.n0 10.4732
R67 VTAIL.n56 VTAIL.n40 10.4732
R68 VTAIL.n36 VTAIL.n20 10.4732
R69 VTAIL.n78 VTAIL.n77 9.45567
R70 VTAIL.n18 VTAIL.n17 9.45567
R71 VTAIL.n58 VTAIL.n57 9.45567
R72 VTAIL.n38 VTAIL.n37 9.45567
R73 VTAIL.n77 VTAIL.n76 9.3005
R74 VTAIL.n62 VTAIL.n61 9.3005
R75 VTAIL.n71 VTAIL.n70 9.3005
R76 VTAIL.n69 VTAIL.n68 9.3005
R77 VTAIL.n17 VTAIL.n16 9.3005
R78 VTAIL.n2 VTAIL.n1 9.3005
R79 VTAIL.n11 VTAIL.n10 9.3005
R80 VTAIL.n9 VTAIL.n8 9.3005
R81 VTAIL.n57 VTAIL.n56 9.3005
R82 VTAIL.n42 VTAIL.n41 9.3005
R83 VTAIL.n51 VTAIL.n50 9.3005
R84 VTAIL.n49 VTAIL.n48 9.3005
R85 VTAIL.n37 VTAIL.n36 9.3005
R86 VTAIL.n22 VTAIL.n21 9.3005
R87 VTAIL.n31 VTAIL.n30 9.3005
R88 VTAIL.n29 VTAIL.n28 9.3005
R89 VTAIL.n69 VTAIL.n65 4.40546
R90 VTAIL.n9 VTAIL.n5 4.40546
R91 VTAIL.n49 VTAIL.n45 4.40546
R92 VTAIL.n29 VTAIL.n25 4.40546
R93 VTAIL.n78 VTAIL.n60 3.49141
R94 VTAIL.n18 VTAIL.n0 3.49141
R95 VTAIL.n58 VTAIL.n40 3.49141
R96 VTAIL.n38 VTAIL.n20 3.49141
R97 VTAIL.n76 VTAIL.n75 2.71565
R98 VTAIL.n16 VTAIL.n15 2.71565
R99 VTAIL.n56 VTAIL.n55 2.71565
R100 VTAIL.n36 VTAIL.n35 2.71565
R101 VTAIL.n72 VTAIL.n62 1.93989
R102 VTAIL.n12 VTAIL.n2 1.93989
R103 VTAIL.n52 VTAIL.n42 1.93989
R104 VTAIL.n32 VTAIL.n22 1.93989
R105 VTAIL.n71 VTAIL.n64 1.16414
R106 VTAIL.n11 VTAIL.n4 1.16414
R107 VTAIL.n51 VTAIL.n44 1.16414
R108 VTAIL.n31 VTAIL.n24 1.16414
R109 VTAIL.n59 VTAIL.n39 0.772052
R110 VTAIL VTAIL.n19 0.679379
R111 VTAIL.n68 VTAIL.n67 0.388379
R112 VTAIL.n8 VTAIL.n7 0.388379
R113 VTAIL.n48 VTAIL.n47 0.388379
R114 VTAIL.n28 VTAIL.n27 0.388379
R115 VTAIL.n70 VTAIL.n69 0.155672
R116 VTAIL.n70 VTAIL.n61 0.155672
R117 VTAIL.n77 VTAIL.n61 0.155672
R118 VTAIL.n10 VTAIL.n9 0.155672
R119 VTAIL.n10 VTAIL.n1 0.155672
R120 VTAIL.n17 VTAIL.n1 0.155672
R121 VTAIL.n57 VTAIL.n41 0.155672
R122 VTAIL.n50 VTAIL.n41 0.155672
R123 VTAIL.n50 VTAIL.n49 0.155672
R124 VTAIL.n37 VTAIL.n21 0.155672
R125 VTAIL.n30 VTAIL.n21 0.155672
R126 VTAIL.n30 VTAIL.n29 0.155672
R127 VTAIL VTAIL.n79 0.0931724
R128 VDD1.n14 VDD1.n0 289.615
R129 VDD1.n33 VDD1.n19 289.615
R130 VDD1.n15 VDD1.n14 185
R131 VDD1.n13 VDD1.n12 185
R132 VDD1.n4 VDD1.n3 185
R133 VDD1.n7 VDD1.n6 185
R134 VDD1.n26 VDD1.n25 185
R135 VDD1.n23 VDD1.n22 185
R136 VDD1.n32 VDD1.n31 185
R137 VDD1.n34 VDD1.n33 185
R138 VDD1.t0 VDD1.n5 147.888
R139 VDD1.t1 VDD1.n24 147.888
R140 VDD1.n14 VDD1.n13 104.615
R141 VDD1.n13 VDD1.n3 104.615
R142 VDD1.n6 VDD1.n3 104.615
R143 VDD1.n25 VDD1.n22 104.615
R144 VDD1.n32 VDD1.n22 104.615
R145 VDD1.n33 VDD1.n32 104.615
R146 VDD1 VDD1.n37 78.1389
R147 VDD1.n6 VDD1.t0 52.3082
R148 VDD1.n25 VDD1.t1 52.3082
R149 VDD1 VDD1.n18 49.4611
R150 VDD1.n7 VDD1.n5 15.6496
R151 VDD1.n26 VDD1.n24 15.6496
R152 VDD1.n8 VDD1.n4 12.8005
R153 VDD1.n27 VDD1.n23 12.8005
R154 VDD1.n12 VDD1.n11 12.0247
R155 VDD1.n31 VDD1.n30 12.0247
R156 VDD1.n15 VDD1.n2 11.249
R157 VDD1.n34 VDD1.n21 11.249
R158 VDD1.n16 VDD1.n0 10.4732
R159 VDD1.n35 VDD1.n19 10.4732
R160 VDD1.n18 VDD1.n17 9.45567
R161 VDD1.n37 VDD1.n36 9.45567
R162 VDD1.n17 VDD1.n16 9.3005
R163 VDD1.n2 VDD1.n1 9.3005
R164 VDD1.n11 VDD1.n10 9.3005
R165 VDD1.n9 VDD1.n8 9.3005
R166 VDD1.n36 VDD1.n35 9.3005
R167 VDD1.n21 VDD1.n20 9.3005
R168 VDD1.n30 VDD1.n29 9.3005
R169 VDD1.n28 VDD1.n27 9.3005
R170 VDD1.n9 VDD1.n5 4.40546
R171 VDD1.n28 VDD1.n24 4.40546
R172 VDD1.n18 VDD1.n0 3.49141
R173 VDD1.n37 VDD1.n19 3.49141
R174 VDD1.n16 VDD1.n15 2.71565
R175 VDD1.n35 VDD1.n34 2.71565
R176 VDD1.n12 VDD1.n2 1.93989
R177 VDD1.n31 VDD1.n21 1.93989
R178 VDD1.n11 VDD1.n4 1.16414
R179 VDD1.n30 VDD1.n23 1.16414
R180 VDD1.n8 VDD1.n7 0.388379
R181 VDD1.n27 VDD1.n26 0.388379
R182 VDD1.n17 VDD1.n1 0.155672
R183 VDD1.n10 VDD1.n1 0.155672
R184 VDD1.n10 VDD1.n9 0.155672
R185 VDD1.n29 VDD1.n28 0.155672
R186 VDD1.n29 VDD1.n20 0.155672
R187 VDD1.n36 VDD1.n20 0.155672
R188 B.n334 B.n333 585
R189 B.n335 B.n334 585
R190 B.n140 B.n49 585
R191 B.n139 B.n138 585
R192 B.n137 B.n136 585
R193 B.n135 B.n134 585
R194 B.n133 B.n132 585
R195 B.n131 B.n130 585
R196 B.n129 B.n128 585
R197 B.n127 B.n126 585
R198 B.n125 B.n124 585
R199 B.n123 B.n122 585
R200 B.n121 B.n120 585
R201 B.n119 B.n118 585
R202 B.n117 B.n116 585
R203 B.n115 B.n114 585
R204 B.n113 B.n112 585
R205 B.n111 B.n110 585
R206 B.n109 B.n108 585
R207 B.n106 B.n105 585
R208 B.n104 B.n103 585
R209 B.n102 B.n101 585
R210 B.n100 B.n99 585
R211 B.n98 B.n97 585
R212 B.n96 B.n95 585
R213 B.n94 B.n93 585
R214 B.n92 B.n91 585
R215 B.n90 B.n89 585
R216 B.n88 B.n87 585
R217 B.n86 B.n85 585
R218 B.n84 B.n83 585
R219 B.n82 B.n81 585
R220 B.n80 B.n79 585
R221 B.n78 B.n77 585
R222 B.n76 B.n75 585
R223 B.n74 B.n73 585
R224 B.n72 B.n71 585
R225 B.n70 B.n69 585
R226 B.n68 B.n67 585
R227 B.n66 B.n65 585
R228 B.n64 B.n63 585
R229 B.n62 B.n61 585
R230 B.n60 B.n59 585
R231 B.n58 B.n57 585
R232 B.n56 B.n55 585
R233 B.n25 B.n24 585
R234 B.n332 B.n26 585
R235 B.n336 B.n26 585
R236 B.n331 B.n330 585
R237 B.n330 B.n22 585
R238 B.n329 B.n21 585
R239 B.n342 B.n21 585
R240 B.n328 B.n20 585
R241 B.n343 B.n20 585
R242 B.n327 B.n19 585
R243 B.n344 B.n19 585
R244 B.n326 B.n325 585
R245 B.n325 B.n15 585
R246 B.n324 B.n14 585
R247 B.n350 B.n14 585
R248 B.n323 B.n13 585
R249 B.n351 B.n13 585
R250 B.n322 B.n12 585
R251 B.n352 B.n12 585
R252 B.n321 B.n320 585
R253 B.n320 B.n11 585
R254 B.n319 B.n7 585
R255 B.n358 B.n7 585
R256 B.n318 B.n6 585
R257 B.n359 B.n6 585
R258 B.n317 B.n5 585
R259 B.n360 B.n5 585
R260 B.n316 B.n315 585
R261 B.n315 B.n4 585
R262 B.n314 B.n141 585
R263 B.n314 B.n313 585
R264 B.n303 B.n142 585
R265 B.n306 B.n142 585
R266 B.n305 B.n304 585
R267 B.n307 B.n305 585
R268 B.n302 B.n147 585
R269 B.n147 B.n146 585
R270 B.n301 B.n300 585
R271 B.n300 B.n299 585
R272 B.n149 B.n148 585
R273 B.n150 B.n149 585
R274 B.n292 B.n291 585
R275 B.n293 B.n292 585
R276 B.n290 B.n155 585
R277 B.n155 B.n154 585
R278 B.n289 B.n288 585
R279 B.n288 B.n287 585
R280 B.n157 B.n156 585
R281 B.n158 B.n157 585
R282 B.n280 B.n279 585
R283 B.n281 B.n280 585
R284 B.n161 B.n160 585
R285 B.n190 B.n188 585
R286 B.n191 B.n187 585
R287 B.n191 B.n162 585
R288 B.n194 B.n193 585
R289 B.n195 B.n186 585
R290 B.n197 B.n196 585
R291 B.n199 B.n185 585
R292 B.n202 B.n201 585
R293 B.n203 B.n184 585
R294 B.n205 B.n204 585
R295 B.n207 B.n183 585
R296 B.n210 B.n209 585
R297 B.n211 B.n182 585
R298 B.n213 B.n212 585
R299 B.n215 B.n181 585
R300 B.n218 B.n217 585
R301 B.n219 B.n180 585
R302 B.n224 B.n223 585
R303 B.n226 B.n179 585
R304 B.n229 B.n228 585
R305 B.n230 B.n178 585
R306 B.n232 B.n231 585
R307 B.n234 B.n177 585
R308 B.n237 B.n236 585
R309 B.n238 B.n176 585
R310 B.n240 B.n239 585
R311 B.n242 B.n175 585
R312 B.n245 B.n244 585
R313 B.n246 B.n171 585
R314 B.n248 B.n247 585
R315 B.n250 B.n170 585
R316 B.n253 B.n252 585
R317 B.n254 B.n169 585
R318 B.n256 B.n255 585
R319 B.n258 B.n168 585
R320 B.n261 B.n260 585
R321 B.n262 B.n167 585
R322 B.n264 B.n263 585
R323 B.n266 B.n166 585
R324 B.n269 B.n268 585
R325 B.n270 B.n165 585
R326 B.n272 B.n271 585
R327 B.n274 B.n164 585
R328 B.n277 B.n276 585
R329 B.n278 B.n163 585
R330 B.n283 B.n282 585
R331 B.n282 B.n281 585
R332 B.n284 B.n159 585
R333 B.n159 B.n158 585
R334 B.n286 B.n285 585
R335 B.n287 B.n286 585
R336 B.n153 B.n152 585
R337 B.n154 B.n153 585
R338 B.n295 B.n294 585
R339 B.n294 B.n293 585
R340 B.n296 B.n151 585
R341 B.n151 B.n150 585
R342 B.n298 B.n297 585
R343 B.n299 B.n298 585
R344 B.n145 B.n144 585
R345 B.n146 B.n145 585
R346 B.n309 B.n308 585
R347 B.n308 B.n307 585
R348 B.n310 B.n143 585
R349 B.n306 B.n143 585
R350 B.n312 B.n311 585
R351 B.n313 B.n312 585
R352 B.n2 B.n0 585
R353 B.n4 B.n2 585
R354 B.n3 B.n1 585
R355 B.n359 B.n3 585
R356 B.n357 B.n356 585
R357 B.n358 B.n357 585
R358 B.n355 B.n8 585
R359 B.n11 B.n8 585
R360 B.n354 B.n353 585
R361 B.n353 B.n352 585
R362 B.n10 B.n9 585
R363 B.n351 B.n10 585
R364 B.n349 B.n348 585
R365 B.n350 B.n349 585
R366 B.n347 B.n16 585
R367 B.n16 B.n15 585
R368 B.n346 B.n345 585
R369 B.n345 B.n344 585
R370 B.n18 B.n17 585
R371 B.n343 B.n18 585
R372 B.n341 B.n340 585
R373 B.n342 B.n341 585
R374 B.n339 B.n23 585
R375 B.n23 B.n22 585
R376 B.n338 B.n337 585
R377 B.n337 B.n336 585
R378 B.n362 B.n361 585
R379 B.n361 B.n360 585
R380 B.n282 B.n161 540.549
R381 B.n337 B.n25 540.549
R382 B.n280 B.n163 540.549
R383 B.n334 B.n26 540.549
R384 B.n172 B.t13 462.063
R385 B.n220 B.t6 462.063
R386 B.n52 B.t10 462.063
R387 B.n50 B.t2 462.063
R388 B.n335 B.n48 256.663
R389 B.n335 B.n47 256.663
R390 B.n335 B.n46 256.663
R391 B.n335 B.n45 256.663
R392 B.n335 B.n44 256.663
R393 B.n335 B.n43 256.663
R394 B.n335 B.n42 256.663
R395 B.n335 B.n41 256.663
R396 B.n335 B.n40 256.663
R397 B.n335 B.n39 256.663
R398 B.n335 B.n38 256.663
R399 B.n335 B.n37 256.663
R400 B.n335 B.n36 256.663
R401 B.n335 B.n35 256.663
R402 B.n335 B.n34 256.663
R403 B.n335 B.n33 256.663
R404 B.n335 B.n32 256.663
R405 B.n335 B.n31 256.663
R406 B.n335 B.n30 256.663
R407 B.n335 B.n29 256.663
R408 B.n335 B.n28 256.663
R409 B.n335 B.n27 256.663
R410 B.n189 B.n162 256.663
R411 B.n192 B.n162 256.663
R412 B.n198 B.n162 256.663
R413 B.n200 B.n162 256.663
R414 B.n206 B.n162 256.663
R415 B.n208 B.n162 256.663
R416 B.n214 B.n162 256.663
R417 B.n216 B.n162 256.663
R418 B.n225 B.n162 256.663
R419 B.n227 B.n162 256.663
R420 B.n233 B.n162 256.663
R421 B.n235 B.n162 256.663
R422 B.n241 B.n162 256.663
R423 B.n243 B.n162 256.663
R424 B.n249 B.n162 256.663
R425 B.n251 B.n162 256.663
R426 B.n257 B.n162 256.663
R427 B.n259 B.n162 256.663
R428 B.n265 B.n162 256.663
R429 B.n267 B.n162 256.663
R430 B.n273 B.n162 256.663
R431 B.n275 B.n162 256.663
R432 B.n281 B.n162 167.013
R433 B.n336 B.n335 167.013
R434 B.n282 B.n159 163.367
R435 B.n286 B.n159 163.367
R436 B.n286 B.n153 163.367
R437 B.n294 B.n153 163.367
R438 B.n294 B.n151 163.367
R439 B.n298 B.n151 163.367
R440 B.n298 B.n145 163.367
R441 B.n308 B.n145 163.367
R442 B.n308 B.n143 163.367
R443 B.n312 B.n143 163.367
R444 B.n312 B.n2 163.367
R445 B.n361 B.n2 163.367
R446 B.n361 B.n3 163.367
R447 B.n357 B.n3 163.367
R448 B.n357 B.n8 163.367
R449 B.n353 B.n8 163.367
R450 B.n353 B.n10 163.367
R451 B.n349 B.n10 163.367
R452 B.n349 B.n16 163.367
R453 B.n345 B.n16 163.367
R454 B.n345 B.n18 163.367
R455 B.n341 B.n18 163.367
R456 B.n341 B.n23 163.367
R457 B.n337 B.n23 163.367
R458 B.n191 B.n190 163.367
R459 B.n193 B.n191 163.367
R460 B.n197 B.n186 163.367
R461 B.n201 B.n199 163.367
R462 B.n205 B.n184 163.367
R463 B.n209 B.n207 163.367
R464 B.n213 B.n182 163.367
R465 B.n217 B.n215 163.367
R466 B.n224 B.n180 163.367
R467 B.n228 B.n226 163.367
R468 B.n232 B.n178 163.367
R469 B.n236 B.n234 163.367
R470 B.n240 B.n176 163.367
R471 B.n244 B.n242 163.367
R472 B.n248 B.n171 163.367
R473 B.n252 B.n250 163.367
R474 B.n256 B.n169 163.367
R475 B.n260 B.n258 163.367
R476 B.n264 B.n167 163.367
R477 B.n268 B.n266 163.367
R478 B.n272 B.n165 163.367
R479 B.n276 B.n274 163.367
R480 B.n280 B.n157 163.367
R481 B.n288 B.n157 163.367
R482 B.n288 B.n155 163.367
R483 B.n292 B.n155 163.367
R484 B.n292 B.n149 163.367
R485 B.n300 B.n149 163.367
R486 B.n300 B.n147 163.367
R487 B.n305 B.n147 163.367
R488 B.n305 B.n142 163.367
R489 B.n314 B.n142 163.367
R490 B.n315 B.n314 163.367
R491 B.n315 B.n5 163.367
R492 B.n6 B.n5 163.367
R493 B.n7 B.n6 163.367
R494 B.n320 B.n7 163.367
R495 B.n320 B.n12 163.367
R496 B.n13 B.n12 163.367
R497 B.n14 B.n13 163.367
R498 B.n325 B.n14 163.367
R499 B.n325 B.n19 163.367
R500 B.n20 B.n19 163.367
R501 B.n21 B.n20 163.367
R502 B.n330 B.n21 163.367
R503 B.n330 B.n26 163.367
R504 B.n57 B.n56 163.367
R505 B.n61 B.n60 163.367
R506 B.n65 B.n64 163.367
R507 B.n69 B.n68 163.367
R508 B.n73 B.n72 163.367
R509 B.n77 B.n76 163.367
R510 B.n81 B.n80 163.367
R511 B.n85 B.n84 163.367
R512 B.n89 B.n88 163.367
R513 B.n93 B.n92 163.367
R514 B.n97 B.n96 163.367
R515 B.n101 B.n100 163.367
R516 B.n105 B.n104 163.367
R517 B.n110 B.n109 163.367
R518 B.n114 B.n113 163.367
R519 B.n118 B.n117 163.367
R520 B.n122 B.n121 163.367
R521 B.n126 B.n125 163.367
R522 B.n130 B.n129 163.367
R523 B.n134 B.n133 163.367
R524 B.n138 B.n137 163.367
R525 B.n334 B.n49 163.367
R526 B.n172 B.t15 156.12
R527 B.n50 B.t4 156.12
R528 B.n220 B.t9 156.12
R529 B.n52 B.t11 156.12
R530 B.n173 B.t14 142.546
R531 B.n51 B.t5 142.546
R532 B.n221 B.t8 142.544
R533 B.n53 B.t12 142.544
R534 B.n281 B.n158 81.7045
R535 B.n287 B.n158 81.7045
R536 B.n287 B.n154 81.7045
R537 B.n293 B.n154 81.7045
R538 B.n299 B.n150 81.7045
R539 B.n299 B.n146 81.7045
R540 B.n307 B.n146 81.7045
R541 B.n307 B.n306 81.7045
R542 B.n313 B.n4 81.7045
R543 B.n360 B.n4 81.7045
R544 B.n360 B.n359 81.7045
R545 B.n359 B.n358 81.7045
R546 B.n352 B.n11 81.7045
R547 B.n352 B.n351 81.7045
R548 B.n351 B.n350 81.7045
R549 B.n350 B.n15 81.7045
R550 B.n344 B.n343 81.7045
R551 B.n343 B.n342 81.7045
R552 B.n342 B.n22 81.7045
R553 B.n336 B.n22 81.7045
R554 B.t7 B.n150 73.2938
R555 B.t3 B.n15 73.2938
R556 B.n189 B.n161 71.676
R557 B.n193 B.n192 71.676
R558 B.n198 B.n197 71.676
R559 B.n201 B.n200 71.676
R560 B.n206 B.n205 71.676
R561 B.n209 B.n208 71.676
R562 B.n214 B.n213 71.676
R563 B.n217 B.n216 71.676
R564 B.n225 B.n224 71.676
R565 B.n228 B.n227 71.676
R566 B.n233 B.n232 71.676
R567 B.n236 B.n235 71.676
R568 B.n241 B.n240 71.676
R569 B.n244 B.n243 71.676
R570 B.n249 B.n248 71.676
R571 B.n252 B.n251 71.676
R572 B.n257 B.n256 71.676
R573 B.n260 B.n259 71.676
R574 B.n265 B.n264 71.676
R575 B.n268 B.n267 71.676
R576 B.n273 B.n272 71.676
R577 B.n276 B.n275 71.676
R578 B.n27 B.n25 71.676
R579 B.n57 B.n28 71.676
R580 B.n61 B.n29 71.676
R581 B.n65 B.n30 71.676
R582 B.n69 B.n31 71.676
R583 B.n73 B.n32 71.676
R584 B.n77 B.n33 71.676
R585 B.n81 B.n34 71.676
R586 B.n85 B.n35 71.676
R587 B.n89 B.n36 71.676
R588 B.n93 B.n37 71.676
R589 B.n97 B.n38 71.676
R590 B.n101 B.n39 71.676
R591 B.n105 B.n40 71.676
R592 B.n110 B.n41 71.676
R593 B.n114 B.n42 71.676
R594 B.n118 B.n43 71.676
R595 B.n122 B.n44 71.676
R596 B.n126 B.n45 71.676
R597 B.n130 B.n46 71.676
R598 B.n134 B.n47 71.676
R599 B.n138 B.n48 71.676
R600 B.n49 B.n48 71.676
R601 B.n137 B.n47 71.676
R602 B.n133 B.n46 71.676
R603 B.n129 B.n45 71.676
R604 B.n125 B.n44 71.676
R605 B.n121 B.n43 71.676
R606 B.n117 B.n42 71.676
R607 B.n113 B.n41 71.676
R608 B.n109 B.n40 71.676
R609 B.n104 B.n39 71.676
R610 B.n100 B.n38 71.676
R611 B.n96 B.n37 71.676
R612 B.n92 B.n36 71.676
R613 B.n88 B.n35 71.676
R614 B.n84 B.n34 71.676
R615 B.n80 B.n33 71.676
R616 B.n76 B.n32 71.676
R617 B.n72 B.n31 71.676
R618 B.n68 B.n30 71.676
R619 B.n64 B.n29 71.676
R620 B.n60 B.n28 71.676
R621 B.n56 B.n27 71.676
R622 B.n190 B.n189 71.676
R623 B.n192 B.n186 71.676
R624 B.n199 B.n198 71.676
R625 B.n200 B.n184 71.676
R626 B.n207 B.n206 71.676
R627 B.n208 B.n182 71.676
R628 B.n215 B.n214 71.676
R629 B.n216 B.n180 71.676
R630 B.n226 B.n225 71.676
R631 B.n227 B.n178 71.676
R632 B.n234 B.n233 71.676
R633 B.n235 B.n176 71.676
R634 B.n242 B.n241 71.676
R635 B.n243 B.n171 71.676
R636 B.n250 B.n249 71.676
R637 B.n251 B.n169 71.676
R638 B.n258 B.n257 71.676
R639 B.n259 B.n167 71.676
R640 B.n266 B.n265 71.676
R641 B.n267 B.n165 71.676
R642 B.n274 B.n273 71.676
R643 B.n275 B.n163 71.676
R644 B.n174 B.n173 59.5399
R645 B.n222 B.n221 59.5399
R646 B.n54 B.n53 59.5399
R647 B.n107 B.n51 59.5399
R648 B.n313 B.t1 51.6663
R649 B.n358 B.t0 51.6663
R650 B.n338 B.n24 35.1225
R651 B.n333 B.n332 35.1225
R652 B.n279 B.n278 35.1225
R653 B.n283 B.n160 35.1225
R654 B.n306 B.t1 30.0387
R655 B.n11 B.t0 30.0387
R656 B B.n362 18.0485
R657 B.n173 B.n172 13.5763
R658 B.n221 B.n220 13.5763
R659 B.n53 B.n52 13.5763
R660 B.n51 B.n50 13.5763
R661 B.n55 B.n24 10.6151
R662 B.n58 B.n55 10.6151
R663 B.n59 B.n58 10.6151
R664 B.n62 B.n59 10.6151
R665 B.n63 B.n62 10.6151
R666 B.n66 B.n63 10.6151
R667 B.n67 B.n66 10.6151
R668 B.n70 B.n67 10.6151
R669 B.n71 B.n70 10.6151
R670 B.n74 B.n71 10.6151
R671 B.n75 B.n74 10.6151
R672 B.n78 B.n75 10.6151
R673 B.n79 B.n78 10.6151
R674 B.n82 B.n79 10.6151
R675 B.n83 B.n82 10.6151
R676 B.n86 B.n83 10.6151
R677 B.n87 B.n86 10.6151
R678 B.n91 B.n90 10.6151
R679 B.n94 B.n91 10.6151
R680 B.n95 B.n94 10.6151
R681 B.n98 B.n95 10.6151
R682 B.n99 B.n98 10.6151
R683 B.n102 B.n99 10.6151
R684 B.n103 B.n102 10.6151
R685 B.n106 B.n103 10.6151
R686 B.n111 B.n108 10.6151
R687 B.n112 B.n111 10.6151
R688 B.n115 B.n112 10.6151
R689 B.n116 B.n115 10.6151
R690 B.n119 B.n116 10.6151
R691 B.n120 B.n119 10.6151
R692 B.n123 B.n120 10.6151
R693 B.n124 B.n123 10.6151
R694 B.n127 B.n124 10.6151
R695 B.n128 B.n127 10.6151
R696 B.n131 B.n128 10.6151
R697 B.n132 B.n131 10.6151
R698 B.n135 B.n132 10.6151
R699 B.n136 B.n135 10.6151
R700 B.n139 B.n136 10.6151
R701 B.n140 B.n139 10.6151
R702 B.n333 B.n140 10.6151
R703 B.n279 B.n156 10.6151
R704 B.n289 B.n156 10.6151
R705 B.n290 B.n289 10.6151
R706 B.n291 B.n290 10.6151
R707 B.n291 B.n148 10.6151
R708 B.n301 B.n148 10.6151
R709 B.n302 B.n301 10.6151
R710 B.n304 B.n302 10.6151
R711 B.n304 B.n303 10.6151
R712 B.n303 B.n141 10.6151
R713 B.n316 B.n141 10.6151
R714 B.n317 B.n316 10.6151
R715 B.n318 B.n317 10.6151
R716 B.n319 B.n318 10.6151
R717 B.n321 B.n319 10.6151
R718 B.n322 B.n321 10.6151
R719 B.n323 B.n322 10.6151
R720 B.n324 B.n323 10.6151
R721 B.n326 B.n324 10.6151
R722 B.n327 B.n326 10.6151
R723 B.n328 B.n327 10.6151
R724 B.n329 B.n328 10.6151
R725 B.n331 B.n329 10.6151
R726 B.n332 B.n331 10.6151
R727 B.n188 B.n160 10.6151
R728 B.n188 B.n187 10.6151
R729 B.n194 B.n187 10.6151
R730 B.n195 B.n194 10.6151
R731 B.n196 B.n195 10.6151
R732 B.n196 B.n185 10.6151
R733 B.n202 B.n185 10.6151
R734 B.n203 B.n202 10.6151
R735 B.n204 B.n203 10.6151
R736 B.n204 B.n183 10.6151
R737 B.n210 B.n183 10.6151
R738 B.n211 B.n210 10.6151
R739 B.n212 B.n211 10.6151
R740 B.n212 B.n181 10.6151
R741 B.n218 B.n181 10.6151
R742 B.n219 B.n218 10.6151
R743 B.n223 B.n219 10.6151
R744 B.n229 B.n179 10.6151
R745 B.n230 B.n229 10.6151
R746 B.n231 B.n230 10.6151
R747 B.n231 B.n177 10.6151
R748 B.n237 B.n177 10.6151
R749 B.n238 B.n237 10.6151
R750 B.n239 B.n238 10.6151
R751 B.n239 B.n175 10.6151
R752 B.n246 B.n245 10.6151
R753 B.n247 B.n246 10.6151
R754 B.n247 B.n170 10.6151
R755 B.n253 B.n170 10.6151
R756 B.n254 B.n253 10.6151
R757 B.n255 B.n254 10.6151
R758 B.n255 B.n168 10.6151
R759 B.n261 B.n168 10.6151
R760 B.n262 B.n261 10.6151
R761 B.n263 B.n262 10.6151
R762 B.n263 B.n166 10.6151
R763 B.n269 B.n166 10.6151
R764 B.n270 B.n269 10.6151
R765 B.n271 B.n270 10.6151
R766 B.n271 B.n164 10.6151
R767 B.n277 B.n164 10.6151
R768 B.n278 B.n277 10.6151
R769 B.n284 B.n283 10.6151
R770 B.n285 B.n284 10.6151
R771 B.n285 B.n152 10.6151
R772 B.n295 B.n152 10.6151
R773 B.n296 B.n295 10.6151
R774 B.n297 B.n296 10.6151
R775 B.n297 B.n144 10.6151
R776 B.n309 B.n144 10.6151
R777 B.n310 B.n309 10.6151
R778 B.n311 B.n310 10.6151
R779 B.n311 B.n0 10.6151
R780 B.n356 B.n1 10.6151
R781 B.n356 B.n355 10.6151
R782 B.n355 B.n354 10.6151
R783 B.n354 B.n9 10.6151
R784 B.n348 B.n9 10.6151
R785 B.n348 B.n347 10.6151
R786 B.n347 B.n346 10.6151
R787 B.n346 B.n17 10.6151
R788 B.n340 B.n17 10.6151
R789 B.n340 B.n339 10.6151
R790 B.n339 B.n338 10.6151
R791 B.n293 B.t7 8.4112
R792 B.n344 B.t3 8.4112
R793 B.n90 B.n54 7.18099
R794 B.n107 B.n106 7.18099
R795 B.n222 B.n179 7.18099
R796 B.n175 B.n174 7.18099
R797 B.n87 B.n54 3.43465
R798 B.n108 B.n107 3.43465
R799 B.n223 B.n222 3.43465
R800 B.n245 B.n174 3.43465
R801 B.n362 B.n0 2.81026
R802 B.n362 B.n1 2.81026
R803 VN VN.t0 551.864
R804 VN VN.t1 518.943
R805 VDD2.n33 VDD2.n19 289.615
R806 VDD2.n14 VDD2.n0 289.615
R807 VDD2.n34 VDD2.n33 185
R808 VDD2.n32 VDD2.n31 185
R809 VDD2.n23 VDD2.n22 185
R810 VDD2.n26 VDD2.n25 185
R811 VDD2.n7 VDD2.n6 185
R812 VDD2.n4 VDD2.n3 185
R813 VDD2.n13 VDD2.n12 185
R814 VDD2.n15 VDD2.n14 185
R815 VDD2.t1 VDD2.n24 147.888
R816 VDD2.t0 VDD2.n5 147.888
R817 VDD2.n33 VDD2.n32 104.615
R818 VDD2.n32 VDD2.n22 104.615
R819 VDD2.n25 VDD2.n22 104.615
R820 VDD2.n6 VDD2.n3 104.615
R821 VDD2.n13 VDD2.n3 104.615
R822 VDD2.n14 VDD2.n13 104.615
R823 VDD2.n38 VDD2.n18 77.4632
R824 VDD2.n25 VDD2.t1 52.3082
R825 VDD2.n6 VDD2.t0 52.3082
R826 VDD2.n38 VDD2.n37 49.252
R827 VDD2.n26 VDD2.n24 15.6496
R828 VDD2.n7 VDD2.n5 15.6496
R829 VDD2.n27 VDD2.n23 12.8005
R830 VDD2.n8 VDD2.n4 12.8005
R831 VDD2.n31 VDD2.n30 12.0247
R832 VDD2.n12 VDD2.n11 12.0247
R833 VDD2.n34 VDD2.n21 11.249
R834 VDD2.n15 VDD2.n2 11.249
R835 VDD2.n35 VDD2.n19 10.4732
R836 VDD2.n16 VDD2.n0 10.4732
R837 VDD2.n37 VDD2.n36 9.45567
R838 VDD2.n18 VDD2.n17 9.45567
R839 VDD2.n36 VDD2.n35 9.3005
R840 VDD2.n21 VDD2.n20 9.3005
R841 VDD2.n30 VDD2.n29 9.3005
R842 VDD2.n28 VDD2.n27 9.3005
R843 VDD2.n17 VDD2.n16 9.3005
R844 VDD2.n2 VDD2.n1 9.3005
R845 VDD2.n11 VDD2.n10 9.3005
R846 VDD2.n9 VDD2.n8 9.3005
R847 VDD2.n28 VDD2.n24 4.40546
R848 VDD2.n9 VDD2.n5 4.40546
R849 VDD2.n37 VDD2.n19 3.49141
R850 VDD2.n18 VDD2.n0 3.49141
R851 VDD2.n35 VDD2.n34 2.71565
R852 VDD2.n16 VDD2.n15 2.71565
R853 VDD2.n31 VDD2.n21 1.93989
R854 VDD2.n12 VDD2.n2 1.93989
R855 VDD2.n30 VDD2.n23 1.16414
R856 VDD2.n11 VDD2.n4 1.16414
R857 VDD2.n27 VDD2.n26 0.388379
R858 VDD2.n8 VDD2.n7 0.388379
R859 VDD2 VDD2.n38 0.209552
R860 VDD2.n36 VDD2.n20 0.155672
R861 VDD2.n29 VDD2.n20 0.155672
R862 VDD2.n29 VDD2.n28 0.155672
R863 VDD2.n10 VDD2.n9 0.155672
R864 VDD2.n10 VDD2.n1 0.155672
R865 VDD2.n17 VDD2.n1 0.155672
C0 VP VTAIL 0.534535f
C1 VDD1 VTAIL 2.88135f
C2 VP VDD2 0.244915f
C3 VDD2 VDD1 0.429789f
C4 VTAIL VN 0.520229f
C5 VDD2 VN 0.65874f
C6 VP VDD1 0.748559f
C7 VDD2 VTAIL 2.91707f
C8 VP VN 2.9087f
C9 VDD1 VN 0.1531f
C10 VDD2 B 2.149508f
C11 VDD1 B 3.5469f
C12 VTAIL B 2.815876f
C13 VN B 5.49798f
C14 VP B 2.995479f
C15 VDD2.n0 B 0.024353f
C16 VDD2.n1 B 0.018199f
C17 VDD2.n2 B 0.009779f
C18 VDD2.n3 B 0.023115f
C19 VDD2.n4 B 0.010355f
C20 VDD2.n5 B 0.069232f
C21 VDD2.t0 B 0.038206f
C22 VDD2.n6 B 0.017336f
C23 VDD2.n7 B 0.013605f
C24 VDD2.n8 B 0.009779f
C25 VDD2.n9 B 0.252805f
C26 VDD2.n10 B 0.018199f
C27 VDD2.n11 B 0.009779f
C28 VDD2.n12 B 0.010355f
C29 VDD2.n13 B 0.023115f
C30 VDD2.n14 B 0.047868f
C31 VDD2.n15 B 0.010355f
C32 VDD2.n16 B 0.009779f
C33 VDD2.n17 B 0.042563f
C34 VDD2.n18 B 0.254142f
C35 VDD2.n19 B 0.024353f
C36 VDD2.n20 B 0.018199f
C37 VDD2.n21 B 0.009779f
C38 VDD2.n22 B 0.023115f
C39 VDD2.n23 B 0.010355f
C40 VDD2.n24 B 0.069232f
C41 VDD2.t1 B 0.038206f
C42 VDD2.n25 B 0.017336f
C43 VDD2.n26 B 0.013605f
C44 VDD2.n27 B 0.009779f
C45 VDD2.n28 B 0.252805f
C46 VDD2.n29 B 0.018199f
C47 VDD2.n30 B 0.009779f
C48 VDD2.n31 B 0.010355f
C49 VDD2.n32 B 0.023115f
C50 VDD2.n33 B 0.047868f
C51 VDD2.n34 B 0.010355f
C52 VDD2.n35 B 0.009779f
C53 VDD2.n36 B 0.042563f
C54 VDD2.n37 B 0.039138f
C55 VDD2.n38 B 1.2587f
C56 VN.t1 B 0.212335f
C57 VN.t0 B 0.284731f
C58 VDD1.n0 B 0.023801f
C59 VDD1.n1 B 0.017787f
C60 VDD1.n2 B 0.009558f
C61 VDD1.n3 B 0.022591f
C62 VDD1.n4 B 0.01012f
C63 VDD1.n5 B 0.067664f
C64 VDD1.t0 B 0.037341f
C65 VDD1.n6 B 0.016944f
C66 VDD1.n7 B 0.013296f
C67 VDD1.n8 B 0.009558f
C68 VDD1.n9 B 0.247078f
C69 VDD1.n10 B 0.017787f
C70 VDD1.n11 B 0.009558f
C71 VDD1.n12 B 0.01012f
C72 VDD1.n13 B 0.022591f
C73 VDD1.n14 B 0.046784f
C74 VDD1.n15 B 0.01012f
C75 VDD1.n16 B 0.009558f
C76 VDD1.n17 B 0.041599f
C77 VDD1.n18 B 0.038448f
C78 VDD1.n19 B 0.023801f
C79 VDD1.n20 B 0.017787f
C80 VDD1.n21 B 0.009558f
C81 VDD1.n22 B 0.022591f
C82 VDD1.n23 B 0.01012f
C83 VDD1.n24 B 0.067664f
C84 VDD1.t1 B 0.037341f
C85 VDD1.n25 B 0.016944f
C86 VDD1.n26 B 0.013296f
C87 VDD1.n27 B 0.009558f
C88 VDD1.n28 B 0.247078f
C89 VDD1.n29 B 0.017787f
C90 VDD1.n30 B 0.009558f
C91 VDD1.n31 B 0.01012f
C92 VDD1.n32 B 0.022591f
C93 VDD1.n33 B 0.046784f
C94 VDD1.n34 B 0.01012f
C95 VDD1.n35 B 0.009558f
C96 VDD1.n36 B 0.041599f
C97 VDD1.n37 B 0.266828f
C98 VTAIL.n0 B 0.028411f
C99 VTAIL.n1 B 0.021232f
C100 VTAIL.n2 B 0.011409f
C101 VTAIL.n3 B 0.026967f
C102 VTAIL.n4 B 0.01208f
C103 VTAIL.n5 B 0.080771f
C104 VTAIL.t3 B 0.044574f
C105 VTAIL.n6 B 0.020226f
C106 VTAIL.n7 B 0.015872f
C107 VTAIL.n8 B 0.011409f
C108 VTAIL.n9 B 0.294938f
C109 VTAIL.n10 B 0.021232f
C110 VTAIL.n11 B 0.011409f
C111 VTAIL.n12 B 0.01208f
C112 VTAIL.n13 B 0.026967f
C113 VTAIL.n14 B 0.055846f
C114 VTAIL.n15 B 0.01208f
C115 VTAIL.n16 B 0.011409f
C116 VTAIL.n17 B 0.049657f
C117 VTAIL.n18 B 0.031006f
C118 VTAIL.n19 B 0.664725f
C119 VTAIL.n20 B 0.028411f
C120 VTAIL.n21 B 0.021232f
C121 VTAIL.n22 B 0.011409f
C122 VTAIL.n23 B 0.026967f
C123 VTAIL.n24 B 0.01208f
C124 VTAIL.n25 B 0.080771f
C125 VTAIL.t1 B 0.044574f
C126 VTAIL.n26 B 0.020226f
C127 VTAIL.n27 B 0.015872f
C128 VTAIL.n28 B 0.011409f
C129 VTAIL.n29 B 0.294938f
C130 VTAIL.n30 B 0.021232f
C131 VTAIL.n31 B 0.011409f
C132 VTAIL.n32 B 0.01208f
C133 VTAIL.n33 B 0.026967f
C134 VTAIL.n34 B 0.055846f
C135 VTAIL.n35 B 0.01208f
C136 VTAIL.n36 B 0.011409f
C137 VTAIL.n37 B 0.049657f
C138 VTAIL.n38 B 0.031006f
C139 VTAIL.n39 B 0.671066f
C140 VTAIL.n40 B 0.028411f
C141 VTAIL.n41 B 0.021232f
C142 VTAIL.n42 B 0.011409f
C143 VTAIL.n43 B 0.026967f
C144 VTAIL.n44 B 0.01208f
C145 VTAIL.n45 B 0.080771f
C146 VTAIL.t2 B 0.044574f
C147 VTAIL.n46 B 0.020226f
C148 VTAIL.n47 B 0.015872f
C149 VTAIL.n48 B 0.011409f
C150 VTAIL.n49 B 0.294938f
C151 VTAIL.n50 B 0.021232f
C152 VTAIL.n51 B 0.011409f
C153 VTAIL.n52 B 0.01208f
C154 VTAIL.n53 B 0.026967f
C155 VTAIL.n54 B 0.055846f
C156 VTAIL.n55 B 0.01208f
C157 VTAIL.n56 B 0.011409f
C158 VTAIL.n57 B 0.049657f
C159 VTAIL.n58 B 0.031006f
C160 VTAIL.n59 B 0.629781f
C161 VTAIL.n60 B 0.028411f
C162 VTAIL.n61 B 0.021232f
C163 VTAIL.n62 B 0.011409f
C164 VTAIL.n63 B 0.026967f
C165 VTAIL.n64 B 0.01208f
C166 VTAIL.n65 B 0.080771f
C167 VTAIL.t0 B 0.044574f
C168 VTAIL.n66 B 0.020226f
C169 VTAIL.n67 B 0.015872f
C170 VTAIL.n68 B 0.011409f
C171 VTAIL.n69 B 0.294938f
C172 VTAIL.n70 B 0.021232f
C173 VTAIL.n71 B 0.011409f
C174 VTAIL.n72 B 0.01208f
C175 VTAIL.n73 B 0.026967f
C176 VTAIL.n74 B 0.055846f
C177 VTAIL.n75 B 0.01208f
C178 VTAIL.n76 B 0.011409f
C179 VTAIL.n77 B 0.049657f
C180 VTAIL.n78 B 0.031006f
C181 VTAIL.n79 B 0.583336f
C182 VP.t1 B 0.288299f
C183 VP.t0 B 0.216893f
C184 VP.n0 B 2.38838f
.ends

