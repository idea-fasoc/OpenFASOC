* NGSPICE file created from diff_pair_sample_0263.ext - technology: sky130A

.subckt diff_pair_sample_0263 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8315 pd=11.43 as=1.8315 ps=11.43 w=11.1 l=0.9
X1 VDD2.t5 VN.t1 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=4.329 pd=22.98 as=1.8315 ps=11.43 w=11.1 l=0.9
X2 VTAIL.t9 VN.t2 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.8315 pd=11.43 as=1.8315 ps=11.43 w=11.1 l=0.9
X3 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=4.329 pd=22.98 as=0 ps=0 w=11.1 l=0.9
X4 VDD1.t5 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.329 pd=22.98 as=1.8315 ps=11.43 w=11.1 l=0.9
X5 VDD2.t2 VN.t3 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=1.8315 pd=11.43 as=4.329 ps=22.98 w=11.1 l=0.9
X6 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=4.329 pd=22.98 as=0 ps=0 w=11.1 l=0.9
X7 VDD1.t4 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.8315 pd=11.43 as=4.329 ps=22.98 w=11.1 l=0.9
X8 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=4.329 pd=22.98 as=0 ps=0 w=11.1 l=0.9
X9 VDD2.t1 VN.t4 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=1.8315 pd=11.43 as=4.329 ps=22.98 w=11.1 l=0.9
X10 VDD1.t3 VP.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.8315 pd=11.43 as=4.329 ps=22.98 w=11.1 l=0.9
X11 VTAIL.t3 VP.t3 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8315 pd=11.43 as=1.8315 ps=11.43 w=11.1 l=0.9
X12 VDD2.t0 VN.t5 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=4.329 pd=22.98 as=1.8315 ps=11.43 w=11.1 l=0.9
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.329 pd=22.98 as=0 ps=0 w=11.1 l=0.9
X14 VDD1.t1 VP.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=4.329 pd=22.98 as=1.8315 ps=11.43 w=11.1 l=0.9
X15 VTAIL.t4 VP.t5 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=1.8315 pd=11.43 as=1.8315 ps=11.43 w=11.1 l=0.9
R0 VN.n2 VN.t1 358.048
R1 VN.n10 VN.t4 358.048
R2 VN.n6 VN.t3 340.882
R3 VN.n14 VN.t5 340.882
R4 VN.n1 VN.t2 297.233
R5 VN.n9 VN.t0 297.233
R6 VN.n7 VN.n6 161.3
R7 VN.n15 VN.n14 161.3
R8 VN.n13 VN.n8 161.3
R9 VN.n12 VN.n11 161.3
R10 VN.n5 VN.n0 161.3
R11 VN.n4 VN.n3 161.3
R12 VN.n5 VN.n4 53.6554
R13 VN.n13 VN.n12 53.6554
R14 VN.n11 VN.n10 43.5444
R15 VN.n3 VN.n2 43.5444
R16 VN.n2 VN.n1 42.6182
R17 VN.n10 VN.n9 42.6182
R18 VN VN.n15 41.6956
R19 VN.n4 VN.n1 12.2964
R20 VN.n12 VN.n9 12.2964
R21 VN.n6 VN.n5 4.38232
R22 VN.n14 VN.n13 4.38232
R23 VN.n15 VN.n8 0.189894
R24 VN.n11 VN.n8 0.189894
R25 VN.n3 VN.n0 0.189894
R26 VN.n7 VN.n0 0.189894
R27 VN VN.n7 0.0516364
R28 VDD2.n1 VDD2.t5 65.8963
R29 VDD2.n2 VDD2.t0 65.1565
R30 VDD2.n1 VDD2.n0 63.5823
R31 VDD2 VDD2.n3 63.5795
R32 VDD2.n2 VDD2.n1 36.7304
R33 VDD2.n3 VDD2.t3 1.78428
R34 VDD2.n3 VDD2.t1 1.78428
R35 VDD2.n0 VDD2.t4 1.78428
R36 VDD2.n0 VDD2.t2 1.78428
R37 VDD2 VDD2.n2 0.853948
R38 VTAIL.n7 VTAIL.t7 48.4777
R39 VTAIL.n11 VTAIL.t8 48.4776
R40 VTAIL.n2 VTAIL.t0 48.4776
R41 VTAIL.n10 VTAIL.t2 48.4776
R42 VTAIL.n9 VTAIL.n8 46.694
R43 VTAIL.n6 VTAIL.n5 46.694
R44 VTAIL.n1 VTAIL.n0 46.6937
R45 VTAIL.n4 VTAIL.n3 46.6937
R46 VTAIL.n6 VTAIL.n4 24.0565
R47 VTAIL.n11 VTAIL.n10 22.9962
R48 VTAIL.n0 VTAIL.t10 1.78428
R49 VTAIL.n0 VTAIL.t9 1.78428
R50 VTAIL.n3 VTAIL.t5 1.78428
R51 VTAIL.n3 VTAIL.t3 1.78428
R52 VTAIL.n8 VTAIL.t1 1.78428
R53 VTAIL.n8 VTAIL.t4 1.78428
R54 VTAIL.n5 VTAIL.t6 1.78428
R55 VTAIL.n5 VTAIL.t11 1.78428
R56 VTAIL.n7 VTAIL.n6 1.06084
R57 VTAIL.n10 VTAIL.n9 1.06084
R58 VTAIL.n4 VTAIL.n2 1.06084
R59 VTAIL.n9 VTAIL.n7 1.0005
R60 VTAIL.n2 VTAIL.n1 1.0005
R61 VTAIL VTAIL.n11 0.737569
R62 VTAIL VTAIL.n1 0.323776
R63 B.n458 B.n457 585
R64 B.n460 B.n93 585
R65 B.n463 B.n462 585
R66 B.n464 B.n92 585
R67 B.n466 B.n465 585
R68 B.n468 B.n91 585
R69 B.n471 B.n470 585
R70 B.n472 B.n90 585
R71 B.n474 B.n473 585
R72 B.n476 B.n89 585
R73 B.n479 B.n478 585
R74 B.n480 B.n88 585
R75 B.n482 B.n481 585
R76 B.n484 B.n87 585
R77 B.n487 B.n486 585
R78 B.n488 B.n86 585
R79 B.n490 B.n489 585
R80 B.n492 B.n85 585
R81 B.n495 B.n494 585
R82 B.n496 B.n84 585
R83 B.n498 B.n497 585
R84 B.n500 B.n83 585
R85 B.n503 B.n502 585
R86 B.n504 B.n82 585
R87 B.n506 B.n505 585
R88 B.n508 B.n81 585
R89 B.n511 B.n510 585
R90 B.n512 B.n80 585
R91 B.n514 B.n513 585
R92 B.n516 B.n79 585
R93 B.n519 B.n518 585
R94 B.n520 B.n78 585
R95 B.n522 B.n521 585
R96 B.n524 B.n77 585
R97 B.n527 B.n526 585
R98 B.n528 B.n76 585
R99 B.n530 B.n529 585
R100 B.n532 B.n75 585
R101 B.n535 B.n534 585
R102 B.n537 B.n72 585
R103 B.n539 B.n538 585
R104 B.n541 B.n71 585
R105 B.n544 B.n543 585
R106 B.n545 B.n70 585
R107 B.n547 B.n546 585
R108 B.n549 B.n69 585
R109 B.n552 B.n551 585
R110 B.n553 B.n65 585
R111 B.n555 B.n554 585
R112 B.n557 B.n64 585
R113 B.n560 B.n559 585
R114 B.n561 B.n63 585
R115 B.n563 B.n562 585
R116 B.n565 B.n62 585
R117 B.n568 B.n567 585
R118 B.n569 B.n61 585
R119 B.n571 B.n570 585
R120 B.n573 B.n60 585
R121 B.n576 B.n575 585
R122 B.n577 B.n59 585
R123 B.n579 B.n578 585
R124 B.n581 B.n58 585
R125 B.n584 B.n583 585
R126 B.n585 B.n57 585
R127 B.n587 B.n586 585
R128 B.n589 B.n56 585
R129 B.n592 B.n591 585
R130 B.n593 B.n55 585
R131 B.n595 B.n594 585
R132 B.n597 B.n54 585
R133 B.n600 B.n599 585
R134 B.n601 B.n53 585
R135 B.n603 B.n602 585
R136 B.n605 B.n52 585
R137 B.n608 B.n607 585
R138 B.n609 B.n51 585
R139 B.n611 B.n610 585
R140 B.n613 B.n50 585
R141 B.n616 B.n615 585
R142 B.n617 B.n49 585
R143 B.n619 B.n618 585
R144 B.n621 B.n48 585
R145 B.n624 B.n623 585
R146 B.n625 B.n47 585
R147 B.n627 B.n626 585
R148 B.n629 B.n46 585
R149 B.n632 B.n631 585
R150 B.n633 B.n45 585
R151 B.n456 B.n43 585
R152 B.n636 B.n43 585
R153 B.n455 B.n42 585
R154 B.n637 B.n42 585
R155 B.n454 B.n41 585
R156 B.n638 B.n41 585
R157 B.n453 B.n452 585
R158 B.n452 B.n37 585
R159 B.n451 B.n36 585
R160 B.n644 B.n36 585
R161 B.n450 B.n35 585
R162 B.n645 B.n35 585
R163 B.n449 B.n34 585
R164 B.n646 B.n34 585
R165 B.n448 B.n447 585
R166 B.n447 B.n30 585
R167 B.n446 B.n29 585
R168 B.n652 B.n29 585
R169 B.n445 B.n28 585
R170 B.n653 B.n28 585
R171 B.n444 B.n27 585
R172 B.n654 B.n27 585
R173 B.n443 B.n442 585
R174 B.n442 B.n26 585
R175 B.n441 B.n22 585
R176 B.n660 B.n22 585
R177 B.n440 B.n21 585
R178 B.n661 B.n21 585
R179 B.n439 B.n20 585
R180 B.n662 B.n20 585
R181 B.n438 B.n437 585
R182 B.n437 B.n19 585
R183 B.n436 B.n15 585
R184 B.n668 B.n15 585
R185 B.n435 B.n14 585
R186 B.n669 B.n14 585
R187 B.n434 B.n13 585
R188 B.n670 B.n13 585
R189 B.n433 B.n432 585
R190 B.n432 B.n12 585
R191 B.n431 B.n430 585
R192 B.n431 B.n8 585
R193 B.n429 B.n7 585
R194 B.n677 B.n7 585
R195 B.n428 B.n6 585
R196 B.n678 B.n6 585
R197 B.n427 B.n5 585
R198 B.n679 B.n5 585
R199 B.n426 B.n425 585
R200 B.n425 B.n4 585
R201 B.n424 B.n94 585
R202 B.n424 B.n423 585
R203 B.n413 B.n95 585
R204 B.n416 B.n95 585
R205 B.n415 B.n414 585
R206 B.n417 B.n415 585
R207 B.n412 B.n100 585
R208 B.n100 B.n99 585
R209 B.n411 B.n410 585
R210 B.n410 B.n409 585
R211 B.n102 B.n101 585
R212 B.n402 B.n102 585
R213 B.n401 B.n400 585
R214 B.n403 B.n401 585
R215 B.n399 B.n107 585
R216 B.n107 B.n106 585
R217 B.n398 B.n397 585
R218 B.n397 B.n396 585
R219 B.n109 B.n108 585
R220 B.n389 B.n109 585
R221 B.n388 B.n387 585
R222 B.n390 B.n388 585
R223 B.n386 B.n114 585
R224 B.n114 B.n113 585
R225 B.n385 B.n384 585
R226 B.n384 B.n383 585
R227 B.n116 B.n115 585
R228 B.n117 B.n116 585
R229 B.n376 B.n375 585
R230 B.n377 B.n376 585
R231 B.n374 B.n121 585
R232 B.n125 B.n121 585
R233 B.n373 B.n372 585
R234 B.n372 B.n371 585
R235 B.n123 B.n122 585
R236 B.n124 B.n123 585
R237 B.n364 B.n363 585
R238 B.n365 B.n364 585
R239 B.n362 B.n130 585
R240 B.n130 B.n129 585
R241 B.n361 B.n360 585
R242 B.n360 B.n359 585
R243 B.n356 B.n134 585
R244 B.n355 B.n354 585
R245 B.n352 B.n135 585
R246 B.n352 B.n133 585
R247 B.n351 B.n350 585
R248 B.n349 B.n348 585
R249 B.n347 B.n137 585
R250 B.n345 B.n344 585
R251 B.n343 B.n138 585
R252 B.n342 B.n341 585
R253 B.n339 B.n139 585
R254 B.n337 B.n336 585
R255 B.n335 B.n140 585
R256 B.n334 B.n333 585
R257 B.n331 B.n141 585
R258 B.n329 B.n328 585
R259 B.n327 B.n142 585
R260 B.n326 B.n325 585
R261 B.n323 B.n143 585
R262 B.n321 B.n320 585
R263 B.n319 B.n144 585
R264 B.n318 B.n317 585
R265 B.n315 B.n145 585
R266 B.n313 B.n312 585
R267 B.n311 B.n146 585
R268 B.n310 B.n309 585
R269 B.n307 B.n147 585
R270 B.n305 B.n304 585
R271 B.n303 B.n148 585
R272 B.n302 B.n301 585
R273 B.n299 B.n149 585
R274 B.n297 B.n296 585
R275 B.n295 B.n150 585
R276 B.n294 B.n293 585
R277 B.n291 B.n151 585
R278 B.n289 B.n288 585
R279 B.n287 B.n152 585
R280 B.n286 B.n285 585
R281 B.n283 B.n153 585
R282 B.n281 B.n280 585
R283 B.n278 B.n154 585
R284 B.n277 B.n276 585
R285 B.n274 B.n157 585
R286 B.n272 B.n271 585
R287 B.n270 B.n158 585
R288 B.n269 B.n268 585
R289 B.n266 B.n159 585
R290 B.n264 B.n263 585
R291 B.n262 B.n160 585
R292 B.n261 B.n260 585
R293 B.n258 B.n257 585
R294 B.n256 B.n255 585
R295 B.n254 B.n165 585
R296 B.n252 B.n251 585
R297 B.n250 B.n166 585
R298 B.n249 B.n248 585
R299 B.n246 B.n167 585
R300 B.n244 B.n243 585
R301 B.n242 B.n168 585
R302 B.n241 B.n240 585
R303 B.n238 B.n169 585
R304 B.n236 B.n235 585
R305 B.n234 B.n170 585
R306 B.n233 B.n232 585
R307 B.n230 B.n171 585
R308 B.n228 B.n227 585
R309 B.n226 B.n172 585
R310 B.n225 B.n224 585
R311 B.n222 B.n173 585
R312 B.n220 B.n219 585
R313 B.n218 B.n174 585
R314 B.n217 B.n216 585
R315 B.n214 B.n175 585
R316 B.n212 B.n211 585
R317 B.n210 B.n176 585
R318 B.n209 B.n208 585
R319 B.n206 B.n177 585
R320 B.n204 B.n203 585
R321 B.n202 B.n178 585
R322 B.n201 B.n200 585
R323 B.n198 B.n179 585
R324 B.n196 B.n195 585
R325 B.n194 B.n180 585
R326 B.n193 B.n192 585
R327 B.n190 B.n181 585
R328 B.n188 B.n187 585
R329 B.n186 B.n182 585
R330 B.n185 B.n184 585
R331 B.n132 B.n131 585
R332 B.n133 B.n132 585
R333 B.n358 B.n357 585
R334 B.n359 B.n358 585
R335 B.n128 B.n127 585
R336 B.n129 B.n128 585
R337 B.n367 B.n366 585
R338 B.n366 B.n365 585
R339 B.n368 B.n126 585
R340 B.n126 B.n124 585
R341 B.n370 B.n369 585
R342 B.n371 B.n370 585
R343 B.n120 B.n119 585
R344 B.n125 B.n120 585
R345 B.n379 B.n378 585
R346 B.n378 B.n377 585
R347 B.n380 B.n118 585
R348 B.n118 B.n117 585
R349 B.n382 B.n381 585
R350 B.n383 B.n382 585
R351 B.n112 B.n111 585
R352 B.n113 B.n112 585
R353 B.n392 B.n391 585
R354 B.n391 B.n390 585
R355 B.n393 B.n110 585
R356 B.n389 B.n110 585
R357 B.n395 B.n394 585
R358 B.n396 B.n395 585
R359 B.n105 B.n104 585
R360 B.n106 B.n105 585
R361 B.n405 B.n404 585
R362 B.n404 B.n403 585
R363 B.n406 B.n103 585
R364 B.n402 B.n103 585
R365 B.n408 B.n407 585
R366 B.n409 B.n408 585
R367 B.n98 B.n97 585
R368 B.n99 B.n98 585
R369 B.n419 B.n418 585
R370 B.n418 B.n417 585
R371 B.n420 B.n96 585
R372 B.n416 B.n96 585
R373 B.n422 B.n421 585
R374 B.n423 B.n422 585
R375 B.n3 B.n0 585
R376 B.n4 B.n3 585
R377 B.n676 B.n1 585
R378 B.n677 B.n676 585
R379 B.n675 B.n674 585
R380 B.n675 B.n8 585
R381 B.n673 B.n9 585
R382 B.n12 B.n9 585
R383 B.n672 B.n671 585
R384 B.n671 B.n670 585
R385 B.n11 B.n10 585
R386 B.n669 B.n11 585
R387 B.n667 B.n666 585
R388 B.n668 B.n667 585
R389 B.n665 B.n16 585
R390 B.n19 B.n16 585
R391 B.n664 B.n663 585
R392 B.n663 B.n662 585
R393 B.n18 B.n17 585
R394 B.n661 B.n18 585
R395 B.n659 B.n658 585
R396 B.n660 B.n659 585
R397 B.n657 B.n23 585
R398 B.n26 B.n23 585
R399 B.n656 B.n655 585
R400 B.n655 B.n654 585
R401 B.n25 B.n24 585
R402 B.n653 B.n25 585
R403 B.n651 B.n650 585
R404 B.n652 B.n651 585
R405 B.n649 B.n31 585
R406 B.n31 B.n30 585
R407 B.n648 B.n647 585
R408 B.n647 B.n646 585
R409 B.n33 B.n32 585
R410 B.n645 B.n33 585
R411 B.n643 B.n642 585
R412 B.n644 B.n643 585
R413 B.n641 B.n38 585
R414 B.n38 B.n37 585
R415 B.n640 B.n639 585
R416 B.n639 B.n638 585
R417 B.n40 B.n39 585
R418 B.n637 B.n40 585
R419 B.n635 B.n634 585
R420 B.n636 B.n635 585
R421 B.n680 B.n679 585
R422 B.n678 B.n2 585
R423 B.n66 B.t13 499.428
R424 B.n73 B.t17 499.428
R425 B.n161 B.t10 499.428
R426 B.n155 B.t6 499.428
R427 B.n635 B.n45 473.281
R428 B.n458 B.n43 473.281
R429 B.n360 B.n132 473.281
R430 B.n358 B.n134 473.281
R431 B.n459 B.n44 256.663
R432 B.n461 B.n44 256.663
R433 B.n467 B.n44 256.663
R434 B.n469 B.n44 256.663
R435 B.n475 B.n44 256.663
R436 B.n477 B.n44 256.663
R437 B.n483 B.n44 256.663
R438 B.n485 B.n44 256.663
R439 B.n491 B.n44 256.663
R440 B.n493 B.n44 256.663
R441 B.n499 B.n44 256.663
R442 B.n501 B.n44 256.663
R443 B.n507 B.n44 256.663
R444 B.n509 B.n44 256.663
R445 B.n515 B.n44 256.663
R446 B.n517 B.n44 256.663
R447 B.n523 B.n44 256.663
R448 B.n525 B.n44 256.663
R449 B.n531 B.n44 256.663
R450 B.n533 B.n44 256.663
R451 B.n540 B.n44 256.663
R452 B.n542 B.n44 256.663
R453 B.n548 B.n44 256.663
R454 B.n550 B.n44 256.663
R455 B.n556 B.n44 256.663
R456 B.n558 B.n44 256.663
R457 B.n564 B.n44 256.663
R458 B.n566 B.n44 256.663
R459 B.n572 B.n44 256.663
R460 B.n574 B.n44 256.663
R461 B.n580 B.n44 256.663
R462 B.n582 B.n44 256.663
R463 B.n588 B.n44 256.663
R464 B.n590 B.n44 256.663
R465 B.n596 B.n44 256.663
R466 B.n598 B.n44 256.663
R467 B.n604 B.n44 256.663
R468 B.n606 B.n44 256.663
R469 B.n612 B.n44 256.663
R470 B.n614 B.n44 256.663
R471 B.n620 B.n44 256.663
R472 B.n622 B.n44 256.663
R473 B.n628 B.n44 256.663
R474 B.n630 B.n44 256.663
R475 B.n353 B.n133 256.663
R476 B.n136 B.n133 256.663
R477 B.n346 B.n133 256.663
R478 B.n340 B.n133 256.663
R479 B.n338 B.n133 256.663
R480 B.n332 B.n133 256.663
R481 B.n330 B.n133 256.663
R482 B.n324 B.n133 256.663
R483 B.n322 B.n133 256.663
R484 B.n316 B.n133 256.663
R485 B.n314 B.n133 256.663
R486 B.n308 B.n133 256.663
R487 B.n306 B.n133 256.663
R488 B.n300 B.n133 256.663
R489 B.n298 B.n133 256.663
R490 B.n292 B.n133 256.663
R491 B.n290 B.n133 256.663
R492 B.n284 B.n133 256.663
R493 B.n282 B.n133 256.663
R494 B.n275 B.n133 256.663
R495 B.n273 B.n133 256.663
R496 B.n267 B.n133 256.663
R497 B.n265 B.n133 256.663
R498 B.n259 B.n133 256.663
R499 B.n164 B.n133 256.663
R500 B.n253 B.n133 256.663
R501 B.n247 B.n133 256.663
R502 B.n245 B.n133 256.663
R503 B.n239 B.n133 256.663
R504 B.n237 B.n133 256.663
R505 B.n231 B.n133 256.663
R506 B.n229 B.n133 256.663
R507 B.n223 B.n133 256.663
R508 B.n221 B.n133 256.663
R509 B.n215 B.n133 256.663
R510 B.n213 B.n133 256.663
R511 B.n207 B.n133 256.663
R512 B.n205 B.n133 256.663
R513 B.n199 B.n133 256.663
R514 B.n197 B.n133 256.663
R515 B.n191 B.n133 256.663
R516 B.n189 B.n133 256.663
R517 B.n183 B.n133 256.663
R518 B.n682 B.n681 256.663
R519 B.n631 B.n629 163.367
R520 B.n627 B.n47 163.367
R521 B.n623 B.n621 163.367
R522 B.n619 B.n49 163.367
R523 B.n615 B.n613 163.367
R524 B.n611 B.n51 163.367
R525 B.n607 B.n605 163.367
R526 B.n603 B.n53 163.367
R527 B.n599 B.n597 163.367
R528 B.n595 B.n55 163.367
R529 B.n591 B.n589 163.367
R530 B.n587 B.n57 163.367
R531 B.n583 B.n581 163.367
R532 B.n579 B.n59 163.367
R533 B.n575 B.n573 163.367
R534 B.n571 B.n61 163.367
R535 B.n567 B.n565 163.367
R536 B.n563 B.n63 163.367
R537 B.n559 B.n557 163.367
R538 B.n555 B.n65 163.367
R539 B.n551 B.n549 163.367
R540 B.n547 B.n70 163.367
R541 B.n543 B.n541 163.367
R542 B.n539 B.n72 163.367
R543 B.n534 B.n532 163.367
R544 B.n530 B.n76 163.367
R545 B.n526 B.n524 163.367
R546 B.n522 B.n78 163.367
R547 B.n518 B.n516 163.367
R548 B.n514 B.n80 163.367
R549 B.n510 B.n508 163.367
R550 B.n506 B.n82 163.367
R551 B.n502 B.n500 163.367
R552 B.n498 B.n84 163.367
R553 B.n494 B.n492 163.367
R554 B.n490 B.n86 163.367
R555 B.n486 B.n484 163.367
R556 B.n482 B.n88 163.367
R557 B.n478 B.n476 163.367
R558 B.n474 B.n90 163.367
R559 B.n470 B.n468 163.367
R560 B.n466 B.n92 163.367
R561 B.n462 B.n460 163.367
R562 B.n360 B.n130 163.367
R563 B.n364 B.n130 163.367
R564 B.n364 B.n123 163.367
R565 B.n372 B.n123 163.367
R566 B.n372 B.n121 163.367
R567 B.n376 B.n121 163.367
R568 B.n376 B.n116 163.367
R569 B.n384 B.n116 163.367
R570 B.n384 B.n114 163.367
R571 B.n388 B.n114 163.367
R572 B.n388 B.n109 163.367
R573 B.n397 B.n109 163.367
R574 B.n397 B.n107 163.367
R575 B.n401 B.n107 163.367
R576 B.n401 B.n102 163.367
R577 B.n410 B.n102 163.367
R578 B.n410 B.n100 163.367
R579 B.n415 B.n100 163.367
R580 B.n415 B.n95 163.367
R581 B.n424 B.n95 163.367
R582 B.n425 B.n424 163.367
R583 B.n425 B.n5 163.367
R584 B.n6 B.n5 163.367
R585 B.n7 B.n6 163.367
R586 B.n431 B.n7 163.367
R587 B.n432 B.n431 163.367
R588 B.n432 B.n13 163.367
R589 B.n14 B.n13 163.367
R590 B.n15 B.n14 163.367
R591 B.n437 B.n15 163.367
R592 B.n437 B.n20 163.367
R593 B.n21 B.n20 163.367
R594 B.n22 B.n21 163.367
R595 B.n442 B.n22 163.367
R596 B.n442 B.n27 163.367
R597 B.n28 B.n27 163.367
R598 B.n29 B.n28 163.367
R599 B.n447 B.n29 163.367
R600 B.n447 B.n34 163.367
R601 B.n35 B.n34 163.367
R602 B.n36 B.n35 163.367
R603 B.n452 B.n36 163.367
R604 B.n452 B.n41 163.367
R605 B.n42 B.n41 163.367
R606 B.n43 B.n42 163.367
R607 B.n354 B.n352 163.367
R608 B.n352 B.n351 163.367
R609 B.n348 B.n347 163.367
R610 B.n345 B.n138 163.367
R611 B.n341 B.n339 163.367
R612 B.n337 B.n140 163.367
R613 B.n333 B.n331 163.367
R614 B.n329 B.n142 163.367
R615 B.n325 B.n323 163.367
R616 B.n321 B.n144 163.367
R617 B.n317 B.n315 163.367
R618 B.n313 B.n146 163.367
R619 B.n309 B.n307 163.367
R620 B.n305 B.n148 163.367
R621 B.n301 B.n299 163.367
R622 B.n297 B.n150 163.367
R623 B.n293 B.n291 163.367
R624 B.n289 B.n152 163.367
R625 B.n285 B.n283 163.367
R626 B.n281 B.n154 163.367
R627 B.n276 B.n274 163.367
R628 B.n272 B.n158 163.367
R629 B.n268 B.n266 163.367
R630 B.n264 B.n160 163.367
R631 B.n260 B.n258 163.367
R632 B.n255 B.n254 163.367
R633 B.n252 B.n166 163.367
R634 B.n248 B.n246 163.367
R635 B.n244 B.n168 163.367
R636 B.n240 B.n238 163.367
R637 B.n236 B.n170 163.367
R638 B.n232 B.n230 163.367
R639 B.n228 B.n172 163.367
R640 B.n224 B.n222 163.367
R641 B.n220 B.n174 163.367
R642 B.n216 B.n214 163.367
R643 B.n212 B.n176 163.367
R644 B.n208 B.n206 163.367
R645 B.n204 B.n178 163.367
R646 B.n200 B.n198 163.367
R647 B.n196 B.n180 163.367
R648 B.n192 B.n190 163.367
R649 B.n188 B.n182 163.367
R650 B.n184 B.n132 163.367
R651 B.n358 B.n128 163.367
R652 B.n366 B.n128 163.367
R653 B.n366 B.n126 163.367
R654 B.n370 B.n126 163.367
R655 B.n370 B.n120 163.367
R656 B.n378 B.n120 163.367
R657 B.n378 B.n118 163.367
R658 B.n382 B.n118 163.367
R659 B.n382 B.n112 163.367
R660 B.n391 B.n112 163.367
R661 B.n391 B.n110 163.367
R662 B.n395 B.n110 163.367
R663 B.n395 B.n105 163.367
R664 B.n404 B.n105 163.367
R665 B.n404 B.n103 163.367
R666 B.n408 B.n103 163.367
R667 B.n408 B.n98 163.367
R668 B.n418 B.n98 163.367
R669 B.n418 B.n96 163.367
R670 B.n422 B.n96 163.367
R671 B.n422 B.n3 163.367
R672 B.n680 B.n3 163.367
R673 B.n676 B.n2 163.367
R674 B.n676 B.n675 163.367
R675 B.n675 B.n9 163.367
R676 B.n671 B.n9 163.367
R677 B.n671 B.n11 163.367
R678 B.n667 B.n11 163.367
R679 B.n667 B.n16 163.367
R680 B.n663 B.n16 163.367
R681 B.n663 B.n18 163.367
R682 B.n659 B.n18 163.367
R683 B.n659 B.n23 163.367
R684 B.n655 B.n23 163.367
R685 B.n655 B.n25 163.367
R686 B.n651 B.n25 163.367
R687 B.n651 B.n31 163.367
R688 B.n647 B.n31 163.367
R689 B.n647 B.n33 163.367
R690 B.n643 B.n33 163.367
R691 B.n643 B.n38 163.367
R692 B.n639 B.n38 163.367
R693 B.n639 B.n40 163.367
R694 B.n635 B.n40 163.367
R695 B.n73 B.t18 96.0434
R696 B.n161 B.t12 96.0434
R697 B.n66 B.t15 96.0297
R698 B.n155 B.t9 96.0297
R699 B.n359 B.n133 86.657
R700 B.n636 B.n44 86.657
R701 B.n74 B.t19 72.1888
R702 B.n162 B.t11 72.1888
R703 B.n67 B.t16 72.1751
R704 B.n156 B.t8 72.1751
R705 B.n630 B.n45 71.676
R706 B.n629 B.n628 71.676
R707 B.n622 B.n47 71.676
R708 B.n621 B.n620 71.676
R709 B.n614 B.n49 71.676
R710 B.n613 B.n612 71.676
R711 B.n606 B.n51 71.676
R712 B.n605 B.n604 71.676
R713 B.n598 B.n53 71.676
R714 B.n597 B.n596 71.676
R715 B.n590 B.n55 71.676
R716 B.n589 B.n588 71.676
R717 B.n582 B.n57 71.676
R718 B.n581 B.n580 71.676
R719 B.n574 B.n59 71.676
R720 B.n573 B.n572 71.676
R721 B.n566 B.n61 71.676
R722 B.n565 B.n564 71.676
R723 B.n558 B.n63 71.676
R724 B.n557 B.n556 71.676
R725 B.n550 B.n65 71.676
R726 B.n549 B.n548 71.676
R727 B.n542 B.n70 71.676
R728 B.n541 B.n540 71.676
R729 B.n533 B.n72 71.676
R730 B.n532 B.n531 71.676
R731 B.n525 B.n76 71.676
R732 B.n524 B.n523 71.676
R733 B.n517 B.n78 71.676
R734 B.n516 B.n515 71.676
R735 B.n509 B.n80 71.676
R736 B.n508 B.n507 71.676
R737 B.n501 B.n82 71.676
R738 B.n500 B.n499 71.676
R739 B.n493 B.n84 71.676
R740 B.n492 B.n491 71.676
R741 B.n485 B.n86 71.676
R742 B.n484 B.n483 71.676
R743 B.n477 B.n88 71.676
R744 B.n476 B.n475 71.676
R745 B.n469 B.n90 71.676
R746 B.n468 B.n467 71.676
R747 B.n461 B.n92 71.676
R748 B.n460 B.n459 71.676
R749 B.n459 B.n458 71.676
R750 B.n462 B.n461 71.676
R751 B.n467 B.n466 71.676
R752 B.n470 B.n469 71.676
R753 B.n475 B.n474 71.676
R754 B.n478 B.n477 71.676
R755 B.n483 B.n482 71.676
R756 B.n486 B.n485 71.676
R757 B.n491 B.n490 71.676
R758 B.n494 B.n493 71.676
R759 B.n499 B.n498 71.676
R760 B.n502 B.n501 71.676
R761 B.n507 B.n506 71.676
R762 B.n510 B.n509 71.676
R763 B.n515 B.n514 71.676
R764 B.n518 B.n517 71.676
R765 B.n523 B.n522 71.676
R766 B.n526 B.n525 71.676
R767 B.n531 B.n530 71.676
R768 B.n534 B.n533 71.676
R769 B.n540 B.n539 71.676
R770 B.n543 B.n542 71.676
R771 B.n548 B.n547 71.676
R772 B.n551 B.n550 71.676
R773 B.n556 B.n555 71.676
R774 B.n559 B.n558 71.676
R775 B.n564 B.n563 71.676
R776 B.n567 B.n566 71.676
R777 B.n572 B.n571 71.676
R778 B.n575 B.n574 71.676
R779 B.n580 B.n579 71.676
R780 B.n583 B.n582 71.676
R781 B.n588 B.n587 71.676
R782 B.n591 B.n590 71.676
R783 B.n596 B.n595 71.676
R784 B.n599 B.n598 71.676
R785 B.n604 B.n603 71.676
R786 B.n607 B.n606 71.676
R787 B.n612 B.n611 71.676
R788 B.n615 B.n614 71.676
R789 B.n620 B.n619 71.676
R790 B.n623 B.n622 71.676
R791 B.n628 B.n627 71.676
R792 B.n631 B.n630 71.676
R793 B.n353 B.n134 71.676
R794 B.n351 B.n136 71.676
R795 B.n347 B.n346 71.676
R796 B.n340 B.n138 71.676
R797 B.n339 B.n338 71.676
R798 B.n332 B.n140 71.676
R799 B.n331 B.n330 71.676
R800 B.n324 B.n142 71.676
R801 B.n323 B.n322 71.676
R802 B.n316 B.n144 71.676
R803 B.n315 B.n314 71.676
R804 B.n308 B.n146 71.676
R805 B.n307 B.n306 71.676
R806 B.n300 B.n148 71.676
R807 B.n299 B.n298 71.676
R808 B.n292 B.n150 71.676
R809 B.n291 B.n290 71.676
R810 B.n284 B.n152 71.676
R811 B.n283 B.n282 71.676
R812 B.n275 B.n154 71.676
R813 B.n274 B.n273 71.676
R814 B.n267 B.n158 71.676
R815 B.n266 B.n265 71.676
R816 B.n259 B.n160 71.676
R817 B.n258 B.n164 71.676
R818 B.n254 B.n253 71.676
R819 B.n247 B.n166 71.676
R820 B.n246 B.n245 71.676
R821 B.n239 B.n168 71.676
R822 B.n238 B.n237 71.676
R823 B.n231 B.n170 71.676
R824 B.n230 B.n229 71.676
R825 B.n223 B.n172 71.676
R826 B.n222 B.n221 71.676
R827 B.n215 B.n174 71.676
R828 B.n214 B.n213 71.676
R829 B.n207 B.n176 71.676
R830 B.n206 B.n205 71.676
R831 B.n199 B.n178 71.676
R832 B.n198 B.n197 71.676
R833 B.n191 B.n180 71.676
R834 B.n190 B.n189 71.676
R835 B.n183 B.n182 71.676
R836 B.n354 B.n353 71.676
R837 B.n348 B.n136 71.676
R838 B.n346 B.n345 71.676
R839 B.n341 B.n340 71.676
R840 B.n338 B.n337 71.676
R841 B.n333 B.n332 71.676
R842 B.n330 B.n329 71.676
R843 B.n325 B.n324 71.676
R844 B.n322 B.n321 71.676
R845 B.n317 B.n316 71.676
R846 B.n314 B.n313 71.676
R847 B.n309 B.n308 71.676
R848 B.n306 B.n305 71.676
R849 B.n301 B.n300 71.676
R850 B.n298 B.n297 71.676
R851 B.n293 B.n292 71.676
R852 B.n290 B.n289 71.676
R853 B.n285 B.n284 71.676
R854 B.n282 B.n281 71.676
R855 B.n276 B.n275 71.676
R856 B.n273 B.n272 71.676
R857 B.n268 B.n267 71.676
R858 B.n265 B.n264 71.676
R859 B.n260 B.n259 71.676
R860 B.n255 B.n164 71.676
R861 B.n253 B.n252 71.676
R862 B.n248 B.n247 71.676
R863 B.n245 B.n244 71.676
R864 B.n240 B.n239 71.676
R865 B.n237 B.n236 71.676
R866 B.n232 B.n231 71.676
R867 B.n229 B.n228 71.676
R868 B.n224 B.n223 71.676
R869 B.n221 B.n220 71.676
R870 B.n216 B.n215 71.676
R871 B.n213 B.n212 71.676
R872 B.n208 B.n207 71.676
R873 B.n205 B.n204 71.676
R874 B.n200 B.n199 71.676
R875 B.n197 B.n196 71.676
R876 B.n192 B.n191 71.676
R877 B.n189 B.n188 71.676
R878 B.n184 B.n183 71.676
R879 B.n681 B.n680 71.676
R880 B.n681 B.n2 71.676
R881 B.n68 B.n67 59.5399
R882 B.n536 B.n74 59.5399
R883 B.n163 B.n162 59.5399
R884 B.n279 B.n156 59.5399
R885 B.n359 B.n129 45.6799
R886 B.n365 B.n129 45.6799
R887 B.n365 B.n124 45.6799
R888 B.n371 B.n124 45.6799
R889 B.n371 B.n125 45.6799
R890 B.n377 B.n117 45.6799
R891 B.n383 B.n117 45.6799
R892 B.n383 B.n113 45.6799
R893 B.n390 B.n113 45.6799
R894 B.n390 B.n389 45.6799
R895 B.n396 B.n106 45.6799
R896 B.n403 B.n106 45.6799
R897 B.n403 B.n402 45.6799
R898 B.n409 B.n99 45.6799
R899 B.n417 B.n99 45.6799
R900 B.n417 B.n416 45.6799
R901 B.n423 B.n4 45.6799
R902 B.n679 B.n4 45.6799
R903 B.n679 B.n678 45.6799
R904 B.n678 B.n677 45.6799
R905 B.n677 B.n8 45.6799
R906 B.n670 B.n12 45.6799
R907 B.n670 B.n669 45.6799
R908 B.n669 B.n668 45.6799
R909 B.n662 B.n19 45.6799
R910 B.n662 B.n661 45.6799
R911 B.n661 B.n660 45.6799
R912 B.n654 B.n26 45.6799
R913 B.n654 B.n653 45.6799
R914 B.n653 B.n652 45.6799
R915 B.n652 B.n30 45.6799
R916 B.n646 B.n30 45.6799
R917 B.n645 B.n644 45.6799
R918 B.n644 B.n37 45.6799
R919 B.n638 B.n37 45.6799
R920 B.n638 B.n637 45.6799
R921 B.n637 B.n636 45.6799
R922 B.n377 B.t7 44.3364
R923 B.n646 B.t14 44.3364
R924 B.n423 B.t0 41.6494
R925 B.t1 B.n8 41.6494
R926 B.n389 B.t5 38.9623
R927 B.n26 B.t2 38.9623
R928 B.n357 B.n356 30.7517
R929 B.n361 B.n131 30.7517
R930 B.n457 B.n456 30.7517
R931 B.n634 B.n633 30.7517
R932 B.n409 B.t3 24.1837
R933 B.n668 B.t4 24.1837
R934 B.n67 B.n66 23.855
R935 B.n74 B.n73 23.855
R936 B.n162 B.n161 23.855
R937 B.n156 B.n155 23.855
R938 B.n402 B.t3 21.4967
R939 B.n19 B.t4 21.4967
R940 B B.n682 18.0485
R941 B.n357 B.n127 10.6151
R942 B.n367 B.n127 10.6151
R943 B.n368 B.n367 10.6151
R944 B.n369 B.n368 10.6151
R945 B.n369 B.n119 10.6151
R946 B.n379 B.n119 10.6151
R947 B.n380 B.n379 10.6151
R948 B.n381 B.n380 10.6151
R949 B.n381 B.n111 10.6151
R950 B.n392 B.n111 10.6151
R951 B.n393 B.n392 10.6151
R952 B.n394 B.n393 10.6151
R953 B.n394 B.n104 10.6151
R954 B.n405 B.n104 10.6151
R955 B.n406 B.n405 10.6151
R956 B.n407 B.n406 10.6151
R957 B.n407 B.n97 10.6151
R958 B.n419 B.n97 10.6151
R959 B.n420 B.n419 10.6151
R960 B.n421 B.n420 10.6151
R961 B.n421 B.n0 10.6151
R962 B.n356 B.n355 10.6151
R963 B.n355 B.n135 10.6151
R964 B.n350 B.n135 10.6151
R965 B.n350 B.n349 10.6151
R966 B.n349 B.n137 10.6151
R967 B.n344 B.n137 10.6151
R968 B.n344 B.n343 10.6151
R969 B.n343 B.n342 10.6151
R970 B.n342 B.n139 10.6151
R971 B.n336 B.n139 10.6151
R972 B.n336 B.n335 10.6151
R973 B.n335 B.n334 10.6151
R974 B.n334 B.n141 10.6151
R975 B.n328 B.n141 10.6151
R976 B.n328 B.n327 10.6151
R977 B.n327 B.n326 10.6151
R978 B.n326 B.n143 10.6151
R979 B.n320 B.n143 10.6151
R980 B.n320 B.n319 10.6151
R981 B.n319 B.n318 10.6151
R982 B.n318 B.n145 10.6151
R983 B.n312 B.n145 10.6151
R984 B.n312 B.n311 10.6151
R985 B.n311 B.n310 10.6151
R986 B.n310 B.n147 10.6151
R987 B.n304 B.n147 10.6151
R988 B.n304 B.n303 10.6151
R989 B.n303 B.n302 10.6151
R990 B.n302 B.n149 10.6151
R991 B.n296 B.n149 10.6151
R992 B.n296 B.n295 10.6151
R993 B.n295 B.n294 10.6151
R994 B.n294 B.n151 10.6151
R995 B.n288 B.n151 10.6151
R996 B.n288 B.n287 10.6151
R997 B.n287 B.n286 10.6151
R998 B.n286 B.n153 10.6151
R999 B.n280 B.n153 10.6151
R1000 B.n278 B.n277 10.6151
R1001 B.n277 B.n157 10.6151
R1002 B.n271 B.n157 10.6151
R1003 B.n271 B.n270 10.6151
R1004 B.n270 B.n269 10.6151
R1005 B.n269 B.n159 10.6151
R1006 B.n263 B.n159 10.6151
R1007 B.n263 B.n262 10.6151
R1008 B.n262 B.n261 10.6151
R1009 B.n257 B.n256 10.6151
R1010 B.n256 B.n165 10.6151
R1011 B.n251 B.n165 10.6151
R1012 B.n251 B.n250 10.6151
R1013 B.n250 B.n249 10.6151
R1014 B.n249 B.n167 10.6151
R1015 B.n243 B.n167 10.6151
R1016 B.n243 B.n242 10.6151
R1017 B.n242 B.n241 10.6151
R1018 B.n241 B.n169 10.6151
R1019 B.n235 B.n169 10.6151
R1020 B.n235 B.n234 10.6151
R1021 B.n234 B.n233 10.6151
R1022 B.n233 B.n171 10.6151
R1023 B.n227 B.n171 10.6151
R1024 B.n227 B.n226 10.6151
R1025 B.n226 B.n225 10.6151
R1026 B.n225 B.n173 10.6151
R1027 B.n219 B.n173 10.6151
R1028 B.n219 B.n218 10.6151
R1029 B.n218 B.n217 10.6151
R1030 B.n217 B.n175 10.6151
R1031 B.n211 B.n175 10.6151
R1032 B.n211 B.n210 10.6151
R1033 B.n210 B.n209 10.6151
R1034 B.n209 B.n177 10.6151
R1035 B.n203 B.n177 10.6151
R1036 B.n203 B.n202 10.6151
R1037 B.n202 B.n201 10.6151
R1038 B.n201 B.n179 10.6151
R1039 B.n195 B.n179 10.6151
R1040 B.n195 B.n194 10.6151
R1041 B.n194 B.n193 10.6151
R1042 B.n193 B.n181 10.6151
R1043 B.n187 B.n181 10.6151
R1044 B.n187 B.n186 10.6151
R1045 B.n186 B.n185 10.6151
R1046 B.n185 B.n131 10.6151
R1047 B.n362 B.n361 10.6151
R1048 B.n363 B.n362 10.6151
R1049 B.n363 B.n122 10.6151
R1050 B.n373 B.n122 10.6151
R1051 B.n374 B.n373 10.6151
R1052 B.n375 B.n374 10.6151
R1053 B.n375 B.n115 10.6151
R1054 B.n385 B.n115 10.6151
R1055 B.n386 B.n385 10.6151
R1056 B.n387 B.n386 10.6151
R1057 B.n387 B.n108 10.6151
R1058 B.n398 B.n108 10.6151
R1059 B.n399 B.n398 10.6151
R1060 B.n400 B.n399 10.6151
R1061 B.n400 B.n101 10.6151
R1062 B.n411 B.n101 10.6151
R1063 B.n412 B.n411 10.6151
R1064 B.n414 B.n412 10.6151
R1065 B.n414 B.n413 10.6151
R1066 B.n413 B.n94 10.6151
R1067 B.n426 B.n94 10.6151
R1068 B.n427 B.n426 10.6151
R1069 B.n428 B.n427 10.6151
R1070 B.n429 B.n428 10.6151
R1071 B.n430 B.n429 10.6151
R1072 B.n433 B.n430 10.6151
R1073 B.n434 B.n433 10.6151
R1074 B.n435 B.n434 10.6151
R1075 B.n436 B.n435 10.6151
R1076 B.n438 B.n436 10.6151
R1077 B.n439 B.n438 10.6151
R1078 B.n440 B.n439 10.6151
R1079 B.n441 B.n440 10.6151
R1080 B.n443 B.n441 10.6151
R1081 B.n444 B.n443 10.6151
R1082 B.n445 B.n444 10.6151
R1083 B.n446 B.n445 10.6151
R1084 B.n448 B.n446 10.6151
R1085 B.n449 B.n448 10.6151
R1086 B.n450 B.n449 10.6151
R1087 B.n451 B.n450 10.6151
R1088 B.n453 B.n451 10.6151
R1089 B.n454 B.n453 10.6151
R1090 B.n455 B.n454 10.6151
R1091 B.n456 B.n455 10.6151
R1092 B.n674 B.n1 10.6151
R1093 B.n674 B.n673 10.6151
R1094 B.n673 B.n672 10.6151
R1095 B.n672 B.n10 10.6151
R1096 B.n666 B.n10 10.6151
R1097 B.n666 B.n665 10.6151
R1098 B.n665 B.n664 10.6151
R1099 B.n664 B.n17 10.6151
R1100 B.n658 B.n17 10.6151
R1101 B.n658 B.n657 10.6151
R1102 B.n657 B.n656 10.6151
R1103 B.n656 B.n24 10.6151
R1104 B.n650 B.n24 10.6151
R1105 B.n650 B.n649 10.6151
R1106 B.n649 B.n648 10.6151
R1107 B.n648 B.n32 10.6151
R1108 B.n642 B.n32 10.6151
R1109 B.n642 B.n641 10.6151
R1110 B.n641 B.n640 10.6151
R1111 B.n640 B.n39 10.6151
R1112 B.n634 B.n39 10.6151
R1113 B.n633 B.n632 10.6151
R1114 B.n632 B.n46 10.6151
R1115 B.n626 B.n46 10.6151
R1116 B.n626 B.n625 10.6151
R1117 B.n625 B.n624 10.6151
R1118 B.n624 B.n48 10.6151
R1119 B.n618 B.n48 10.6151
R1120 B.n618 B.n617 10.6151
R1121 B.n617 B.n616 10.6151
R1122 B.n616 B.n50 10.6151
R1123 B.n610 B.n50 10.6151
R1124 B.n610 B.n609 10.6151
R1125 B.n609 B.n608 10.6151
R1126 B.n608 B.n52 10.6151
R1127 B.n602 B.n52 10.6151
R1128 B.n602 B.n601 10.6151
R1129 B.n601 B.n600 10.6151
R1130 B.n600 B.n54 10.6151
R1131 B.n594 B.n54 10.6151
R1132 B.n594 B.n593 10.6151
R1133 B.n593 B.n592 10.6151
R1134 B.n592 B.n56 10.6151
R1135 B.n586 B.n56 10.6151
R1136 B.n586 B.n585 10.6151
R1137 B.n585 B.n584 10.6151
R1138 B.n584 B.n58 10.6151
R1139 B.n578 B.n58 10.6151
R1140 B.n578 B.n577 10.6151
R1141 B.n577 B.n576 10.6151
R1142 B.n576 B.n60 10.6151
R1143 B.n570 B.n60 10.6151
R1144 B.n570 B.n569 10.6151
R1145 B.n569 B.n568 10.6151
R1146 B.n568 B.n62 10.6151
R1147 B.n562 B.n62 10.6151
R1148 B.n562 B.n561 10.6151
R1149 B.n561 B.n560 10.6151
R1150 B.n560 B.n64 10.6151
R1151 B.n554 B.n553 10.6151
R1152 B.n553 B.n552 10.6151
R1153 B.n552 B.n69 10.6151
R1154 B.n546 B.n69 10.6151
R1155 B.n546 B.n545 10.6151
R1156 B.n545 B.n544 10.6151
R1157 B.n544 B.n71 10.6151
R1158 B.n538 B.n71 10.6151
R1159 B.n538 B.n537 10.6151
R1160 B.n535 B.n75 10.6151
R1161 B.n529 B.n75 10.6151
R1162 B.n529 B.n528 10.6151
R1163 B.n528 B.n527 10.6151
R1164 B.n527 B.n77 10.6151
R1165 B.n521 B.n77 10.6151
R1166 B.n521 B.n520 10.6151
R1167 B.n520 B.n519 10.6151
R1168 B.n519 B.n79 10.6151
R1169 B.n513 B.n79 10.6151
R1170 B.n513 B.n512 10.6151
R1171 B.n512 B.n511 10.6151
R1172 B.n511 B.n81 10.6151
R1173 B.n505 B.n81 10.6151
R1174 B.n505 B.n504 10.6151
R1175 B.n504 B.n503 10.6151
R1176 B.n503 B.n83 10.6151
R1177 B.n497 B.n83 10.6151
R1178 B.n497 B.n496 10.6151
R1179 B.n496 B.n495 10.6151
R1180 B.n495 B.n85 10.6151
R1181 B.n489 B.n85 10.6151
R1182 B.n489 B.n488 10.6151
R1183 B.n488 B.n487 10.6151
R1184 B.n487 B.n87 10.6151
R1185 B.n481 B.n87 10.6151
R1186 B.n481 B.n480 10.6151
R1187 B.n480 B.n479 10.6151
R1188 B.n479 B.n89 10.6151
R1189 B.n473 B.n89 10.6151
R1190 B.n473 B.n472 10.6151
R1191 B.n472 B.n471 10.6151
R1192 B.n471 B.n91 10.6151
R1193 B.n465 B.n91 10.6151
R1194 B.n465 B.n464 10.6151
R1195 B.n464 B.n463 10.6151
R1196 B.n463 B.n93 10.6151
R1197 B.n457 B.n93 10.6151
R1198 B.n280 B.n279 9.36635
R1199 B.n257 B.n163 9.36635
R1200 B.n68 B.n64 9.36635
R1201 B.n536 B.n535 9.36635
R1202 B.n682 B.n0 8.11757
R1203 B.n682 B.n1 8.11757
R1204 B.n396 B.t5 6.71806
R1205 B.n660 B.t2 6.71806
R1206 B.n416 B.t0 4.03103
R1207 B.n12 B.t1 4.03103
R1208 B.n125 B.t7 1.34401
R1209 B.t14 B.n645 1.34401
R1210 B.n279 B.n278 1.24928
R1211 B.n261 B.n163 1.24928
R1212 B.n554 B.n68 1.24928
R1213 B.n537 B.n536 1.24928
R1214 VP.n5 VP.t0 358.048
R1215 VP.n12 VP.t4 340.882
R1216 VP.n19 VP.t2 340.882
R1217 VP.n9 VP.t1 340.882
R1218 VP.n1 VP.t3 297.233
R1219 VP.n4 VP.t5 297.233
R1220 VP.n20 VP.n19 161.3
R1221 VP.n7 VP.n6 161.3
R1222 VP.n8 VP.n3 161.3
R1223 VP.n10 VP.n9 161.3
R1224 VP.n18 VP.n0 161.3
R1225 VP.n17 VP.n16 161.3
R1226 VP.n15 VP.n14 161.3
R1227 VP.n13 VP.n2 161.3
R1228 VP.n12 VP.n11 161.3
R1229 VP.n14 VP.n13 53.6554
R1230 VP.n18 VP.n17 53.6554
R1231 VP.n8 VP.n7 53.6554
R1232 VP.n6 VP.n5 43.5444
R1233 VP.n5 VP.n4 42.6182
R1234 VP.n11 VP.n10 41.3149
R1235 VP.n14 VP.n1 12.2964
R1236 VP.n17 VP.n1 12.2964
R1237 VP.n7 VP.n4 12.2964
R1238 VP.n13 VP.n12 4.38232
R1239 VP.n19 VP.n18 4.38232
R1240 VP.n9 VP.n8 4.38232
R1241 VP.n6 VP.n3 0.189894
R1242 VP.n10 VP.n3 0.189894
R1243 VP.n11 VP.n2 0.189894
R1244 VP.n15 VP.n2 0.189894
R1245 VP.n16 VP.n15 0.189894
R1246 VP.n16 VP.n0 0.189894
R1247 VP.n20 VP.n0 0.189894
R1248 VP VP.n20 0.0516364
R1249 VDD1 VDD1.t5 66.0099
R1250 VDD1.n1 VDD1.t1 65.8963
R1251 VDD1.n1 VDD1.n0 63.5823
R1252 VDD1.n3 VDD1.n2 63.3726
R1253 VDD1.n3 VDD1.n1 37.8436
R1254 VDD1.n2 VDD1.t0 1.78428
R1255 VDD1.n2 VDD1.t4 1.78428
R1256 VDD1.n0 VDD1.t2 1.78428
R1257 VDD1.n0 VDD1.t3 1.78428
R1258 VDD1 VDD1.n3 0.207397
C0 VTAIL VDD1 8.57002f
C1 VN VP 5.10518f
C2 VP VDD2 0.314699f
C3 VP VTAIL 4.32035f
C4 VP VDD1 4.691451f
C5 VN VDD2 4.52948f
C6 VN VTAIL 4.30583f
C7 VN VDD1 0.148745f
C8 VDD2 VTAIL 8.606599f
C9 VDD2 VDD1 0.783354f
C10 VDD2 B 4.485347f
C11 VDD1 B 4.728139f
C12 VTAIL B 6.233491f
C13 VN B 8.107759f
C14 VP B 6.30345f
C15 VDD1.t5 B 2.26361f
C16 VDD1.t1 B 2.26297f
C17 VDD1.t2 B 0.199795f
C18 VDD1.t3 B 0.199795f
C19 VDD1.n0 B 1.77355f
C20 VDD1.n1 B 1.9984f
C21 VDD1.t0 B 0.199795f
C22 VDD1.t4 B 0.199795f
C23 VDD1.n2 B 1.77259f
C24 VDD1.n3 B 2.03974f
C25 VP.n0 B 0.04244f
C26 VP.t3 B 1.15249f
C27 VP.n1 B 0.43491f
C28 VP.n2 B 0.04244f
C29 VP.n3 B 0.04244f
C30 VP.t1 B 1.21065f
C31 VP.t5 B 1.15249f
C32 VP.n4 B 0.474471f
C33 VP.t0 B 1.23421f
C34 VP.n5 B 0.486284f
C35 VP.n6 B 0.178301f
C36 VP.n7 B 0.055065f
C37 VP.n8 B 0.013919f
C38 VP.n9 B 0.479547f
C39 VP.n10 B 1.7041f
C40 VP.n11 B 1.74113f
C41 VP.t4 B 1.21065f
C42 VP.n12 B 0.479547f
C43 VP.n13 B 0.013919f
C44 VP.n14 B 0.055065f
C45 VP.n15 B 0.04244f
C46 VP.n16 B 0.04244f
C47 VP.n17 B 0.055065f
C48 VP.n18 B 0.013919f
C49 VP.t2 B 1.21065f
C50 VP.n19 B 0.479547f
C51 VP.n20 B 0.032889f
C52 VTAIL.t10 B 0.209264f
C53 VTAIL.t9 B 0.209264f
C54 VTAIL.n0 B 1.78848f
C55 VTAIL.n1 B 0.332707f
C56 VTAIL.t0 B 2.28008f
C57 VTAIL.n2 B 0.468482f
C58 VTAIL.t5 B 0.209264f
C59 VTAIL.t3 B 0.209264f
C60 VTAIL.n3 B 1.78848f
C61 VTAIL.n4 B 1.53518f
C62 VTAIL.t6 B 0.209264f
C63 VTAIL.t11 B 0.209264f
C64 VTAIL.n5 B 1.78848f
C65 VTAIL.n6 B 1.53518f
C66 VTAIL.t7 B 2.2801f
C67 VTAIL.n7 B 0.468467f
C68 VTAIL.t1 B 0.209264f
C69 VTAIL.t4 B 0.209264f
C70 VTAIL.n8 B 1.78848f
C71 VTAIL.n9 B 0.389362f
C72 VTAIL.t2 B 2.28008f
C73 VTAIL.n10 B 1.53279f
C74 VTAIL.t8 B 2.28008f
C75 VTAIL.n11 B 1.50794f
C76 VDD2.t5 B 2.24313f
C77 VDD2.t4 B 0.198043f
C78 VDD2.t2 B 0.198043f
C79 VDD2.n0 B 1.758f
C80 VDD2.n1 B 1.90733f
C81 VDD2.t0 B 2.23971f
C82 VDD2.n2 B 2.03937f
C83 VDD2.t3 B 0.198043f
C84 VDD2.t1 B 0.198043f
C85 VDD2.n3 B 1.75798f
C86 VN.n0 B 0.041661f
C87 VN.t2 B 1.13136f
C88 VN.n1 B 0.46577f
C89 VN.t1 B 1.21158f
C90 VN.n2 B 0.477366f
C91 VN.n3 B 0.175031f
C92 VN.n4 B 0.054056f
C93 VN.n5 B 0.013663f
C94 VN.t3 B 1.18845f
C95 VN.n6 B 0.470753f
C96 VN.n7 B 0.032286f
C97 VN.n8 B 0.041661f
C98 VN.t0 B 1.13136f
C99 VN.n9 B 0.46577f
C100 VN.t4 B 1.21158f
C101 VN.n10 B 0.477366f
C102 VN.n11 B 0.175031f
C103 VN.n12 B 0.054056f
C104 VN.n13 B 0.013663f
C105 VN.t5 B 1.18845f
C106 VN.n14 B 0.470753f
C107 VN.n15 B 1.70023f
.ends

