* NGSPICE file created from diff_pair_sample_0717.ext - technology: sky130A

.subckt diff_pair_sample_0717 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t6 w_n2500_n1926# sky130_fd_pr__pfet_01v8 ad=0.79035 pd=5.12 as=0.79035 ps=5.12 w=4.79 l=1.2
X1 B.t11 B.t9 B.t10 w_n2500_n1926# sky130_fd_pr__pfet_01v8 ad=1.8681 pd=10.36 as=0 ps=0 w=4.79 l=1.2
X2 VDD1.t2 VP.t1 VTAIL.t14 w_n2500_n1926# sky130_fd_pr__pfet_01v8 ad=0.79035 pd=5.12 as=1.8681 ps=10.36 w=4.79 l=1.2
X3 B.t8 B.t6 B.t7 w_n2500_n1926# sky130_fd_pr__pfet_01v8 ad=1.8681 pd=10.36 as=0 ps=0 w=4.79 l=1.2
X4 VDD1.t1 VP.t2 VTAIL.t13 w_n2500_n1926# sky130_fd_pr__pfet_01v8 ad=0.79035 pd=5.12 as=0.79035 ps=5.12 w=4.79 l=1.2
X5 VDD2.t7 VN.t0 VTAIL.t6 w_n2500_n1926# sky130_fd_pr__pfet_01v8 ad=0.79035 pd=5.12 as=1.8681 ps=10.36 w=4.79 l=1.2
X6 VTAIL.t3 VN.t1 VDD2.t6 w_n2500_n1926# sky130_fd_pr__pfet_01v8 ad=0.79035 pd=5.12 as=0.79035 ps=5.12 w=4.79 l=1.2
X7 VDD2.t5 VN.t2 VTAIL.t5 w_n2500_n1926# sky130_fd_pr__pfet_01v8 ad=0.79035 pd=5.12 as=1.8681 ps=10.36 w=4.79 l=1.2
X8 VTAIL.t12 VP.t3 VDD1.t3 w_n2500_n1926# sky130_fd_pr__pfet_01v8 ad=0.79035 pd=5.12 as=0.79035 ps=5.12 w=4.79 l=1.2
X9 B.t5 B.t3 B.t4 w_n2500_n1926# sky130_fd_pr__pfet_01v8 ad=1.8681 pd=10.36 as=0 ps=0 w=4.79 l=1.2
X10 VDD1.t4 VP.t4 VTAIL.t11 w_n2500_n1926# sky130_fd_pr__pfet_01v8 ad=0.79035 pd=5.12 as=1.8681 ps=10.36 w=4.79 l=1.2
X11 VDD2.t4 VN.t3 VTAIL.t4 w_n2500_n1926# sky130_fd_pr__pfet_01v8 ad=0.79035 pd=5.12 as=0.79035 ps=5.12 w=4.79 l=1.2
X12 VTAIL.t7 VN.t4 VDD2.t3 w_n2500_n1926# sky130_fd_pr__pfet_01v8 ad=0.79035 pd=5.12 as=0.79035 ps=5.12 w=4.79 l=1.2
X13 VTAIL.t10 VP.t5 VDD1.t5 w_n2500_n1926# sky130_fd_pr__pfet_01v8 ad=1.8681 pd=10.36 as=0.79035 ps=5.12 w=4.79 l=1.2
X14 VTAIL.t2 VN.t5 VDD2.t2 w_n2500_n1926# sky130_fd_pr__pfet_01v8 ad=1.8681 pd=10.36 as=0.79035 ps=5.12 w=4.79 l=1.2
X15 B.t2 B.t0 B.t1 w_n2500_n1926# sky130_fd_pr__pfet_01v8 ad=1.8681 pd=10.36 as=0 ps=0 w=4.79 l=1.2
X16 VTAIL.t9 VP.t6 VDD1.t0 w_n2500_n1926# sky130_fd_pr__pfet_01v8 ad=1.8681 pd=10.36 as=0.79035 ps=5.12 w=4.79 l=1.2
X17 VDD2.t1 VN.t6 VTAIL.t1 w_n2500_n1926# sky130_fd_pr__pfet_01v8 ad=0.79035 pd=5.12 as=0.79035 ps=5.12 w=4.79 l=1.2
X18 VDD1.t7 VP.t7 VTAIL.t8 w_n2500_n1926# sky130_fd_pr__pfet_01v8 ad=0.79035 pd=5.12 as=0.79035 ps=5.12 w=4.79 l=1.2
X19 VTAIL.t0 VN.t7 VDD2.t0 w_n2500_n1926# sky130_fd_pr__pfet_01v8 ad=1.8681 pd=10.36 as=0.79035 ps=5.12 w=4.79 l=1.2
R0 VP.n11 VP.n10 161.3
R1 VP.n12 VP.n7 161.3
R2 VP.n14 VP.n13 161.3
R3 VP.n16 VP.n15 161.3
R4 VP.n17 VP.n5 161.3
R5 VP.n32 VP.n0 161.3
R6 VP.n31 VP.n30 161.3
R7 VP.n29 VP.n28 161.3
R8 VP.n27 VP.n2 161.3
R9 VP.n26 VP.n25 161.3
R10 VP.n24 VP.n23 161.3
R11 VP.n22 VP.n4 161.3
R12 VP.n9 VP.t6 147.639
R13 VP.n21 VP.t5 129.137
R14 VP.n33 VP.t4 129.137
R15 VP.n18 VP.t1 129.137
R16 VP.n3 VP.t2 96.1997
R17 VP.n1 VP.t3 96.1997
R18 VP.n6 VP.t0 96.1997
R19 VP.n8 VP.t7 96.1997
R20 VP.n19 VP.n18 80.6037
R21 VP.n34 VP.n33 80.6037
R22 VP.n21 VP.n20 80.6037
R23 VP.n9 VP.n8 44.8004
R24 VP.n27 VP.n26 40.4934
R25 VP.n28 VP.n27 40.4934
R26 VP.n13 VP.n12 40.4934
R27 VP.n12 VP.n11 40.4934
R28 VP.n20 VP.n19 38.9938
R29 VP.n23 VP.n22 37.5796
R30 VP.n32 VP.n31 37.5796
R31 VP.n17 VP.n16 37.5796
R32 VP.n10 VP.n9 29.7304
R33 VP.n22 VP.n21 28.4823
R34 VP.n33 VP.n32 28.4823
R35 VP.n18 VP.n17 28.4823
R36 VP.n26 VP.n3 12.968
R37 VP.n28 VP.n1 12.968
R38 VP.n13 VP.n6 12.968
R39 VP.n11 VP.n8 12.968
R40 VP.n23 VP.n3 11.5
R41 VP.n31 VP.n1 11.5
R42 VP.n16 VP.n6 11.5
R43 VP.n19 VP.n5 0.285035
R44 VP.n20 VP.n4 0.285035
R45 VP.n34 VP.n0 0.285035
R46 VP.n10 VP.n7 0.189894
R47 VP.n14 VP.n7 0.189894
R48 VP.n15 VP.n14 0.189894
R49 VP.n15 VP.n5 0.189894
R50 VP.n24 VP.n4 0.189894
R51 VP.n25 VP.n24 0.189894
R52 VP.n25 VP.n2 0.189894
R53 VP.n29 VP.n2 0.189894
R54 VP.n30 VP.n29 0.189894
R55 VP.n30 VP.n0 0.189894
R56 VP VP.n34 0.146778
R57 VDD1 VDD1.n0 104.694
R58 VDD1.n3 VDD1.n2 104.579
R59 VDD1.n3 VDD1.n1 104.579
R60 VDD1.n5 VDD1.n4 103.975
R61 VDD1.n5 VDD1.n3 34.363
R62 VDD1.n4 VDD1.t6 6.78651
R63 VDD1.n4 VDD1.t2 6.78651
R64 VDD1.n0 VDD1.t0 6.78651
R65 VDD1.n0 VDD1.t7 6.78651
R66 VDD1.n2 VDD1.t3 6.78651
R67 VDD1.n2 VDD1.t4 6.78651
R68 VDD1.n1 VDD1.t5 6.78651
R69 VDD1.n1 VDD1.t1 6.78651
R70 VDD1 VDD1.n5 0.601793
R71 VTAIL.n11 VTAIL.t9 94.083
R72 VTAIL.n10 VTAIL.t5 94.083
R73 VTAIL.n7 VTAIL.t0 94.083
R74 VTAIL.n14 VTAIL.t14 94.0821
R75 VTAIL.n15 VTAIL.t6 94.082
R76 VTAIL.n2 VTAIL.t2 94.082
R77 VTAIL.n3 VTAIL.t11 94.082
R78 VTAIL.n6 VTAIL.t10 94.082
R79 VTAIL.n13 VTAIL.n12 87.297
R80 VTAIL.n9 VTAIL.n8 87.297
R81 VTAIL.n1 VTAIL.n0 87.296
R82 VTAIL.n5 VTAIL.n4 87.296
R83 VTAIL.n15 VTAIL.n14 17.8152
R84 VTAIL.n7 VTAIL.n6 17.8152
R85 VTAIL.n0 VTAIL.t4 6.78651
R86 VTAIL.n0 VTAIL.t3 6.78651
R87 VTAIL.n4 VTAIL.t13 6.78651
R88 VTAIL.n4 VTAIL.t12 6.78651
R89 VTAIL.n12 VTAIL.t8 6.78651
R90 VTAIL.n12 VTAIL.t15 6.78651
R91 VTAIL.n8 VTAIL.t1 6.78651
R92 VTAIL.n8 VTAIL.t7 6.78651
R93 VTAIL.n9 VTAIL.n7 1.31947
R94 VTAIL.n10 VTAIL.n9 1.31947
R95 VTAIL.n13 VTAIL.n11 1.31947
R96 VTAIL.n14 VTAIL.n13 1.31947
R97 VTAIL.n6 VTAIL.n5 1.31947
R98 VTAIL.n5 VTAIL.n3 1.31947
R99 VTAIL.n2 VTAIL.n1 1.31947
R100 VTAIL VTAIL.n15 1.26128
R101 VTAIL.n11 VTAIL.n10 0.470328
R102 VTAIL.n3 VTAIL.n2 0.470328
R103 VTAIL VTAIL.n1 0.0586897
R104 B.n241 B.n240 585
R105 B.n239 B.n78 585
R106 B.n238 B.n237 585
R107 B.n236 B.n79 585
R108 B.n235 B.n234 585
R109 B.n233 B.n80 585
R110 B.n232 B.n231 585
R111 B.n230 B.n81 585
R112 B.n229 B.n228 585
R113 B.n227 B.n82 585
R114 B.n226 B.n225 585
R115 B.n224 B.n83 585
R116 B.n223 B.n222 585
R117 B.n221 B.n84 585
R118 B.n220 B.n219 585
R119 B.n218 B.n85 585
R120 B.n217 B.n216 585
R121 B.n215 B.n86 585
R122 B.n214 B.n213 585
R123 B.n212 B.n87 585
R124 B.n210 B.n209 585
R125 B.n208 B.n90 585
R126 B.n207 B.n206 585
R127 B.n205 B.n91 585
R128 B.n204 B.n203 585
R129 B.n202 B.n92 585
R130 B.n201 B.n200 585
R131 B.n199 B.n93 585
R132 B.n198 B.n197 585
R133 B.n196 B.n94 585
R134 B.n195 B.n194 585
R135 B.n190 B.n95 585
R136 B.n189 B.n188 585
R137 B.n187 B.n96 585
R138 B.n186 B.n185 585
R139 B.n184 B.n97 585
R140 B.n183 B.n182 585
R141 B.n181 B.n98 585
R142 B.n180 B.n179 585
R143 B.n178 B.n99 585
R144 B.n177 B.n176 585
R145 B.n175 B.n100 585
R146 B.n174 B.n173 585
R147 B.n172 B.n101 585
R148 B.n171 B.n170 585
R149 B.n169 B.n102 585
R150 B.n168 B.n167 585
R151 B.n166 B.n103 585
R152 B.n165 B.n164 585
R153 B.n163 B.n104 585
R154 B.n242 B.n77 585
R155 B.n244 B.n243 585
R156 B.n245 B.n76 585
R157 B.n247 B.n246 585
R158 B.n248 B.n75 585
R159 B.n250 B.n249 585
R160 B.n251 B.n74 585
R161 B.n253 B.n252 585
R162 B.n254 B.n73 585
R163 B.n256 B.n255 585
R164 B.n257 B.n72 585
R165 B.n259 B.n258 585
R166 B.n260 B.n71 585
R167 B.n262 B.n261 585
R168 B.n263 B.n70 585
R169 B.n265 B.n264 585
R170 B.n266 B.n69 585
R171 B.n268 B.n267 585
R172 B.n269 B.n68 585
R173 B.n271 B.n270 585
R174 B.n272 B.n67 585
R175 B.n274 B.n273 585
R176 B.n275 B.n66 585
R177 B.n277 B.n276 585
R178 B.n278 B.n65 585
R179 B.n280 B.n279 585
R180 B.n281 B.n64 585
R181 B.n283 B.n282 585
R182 B.n284 B.n63 585
R183 B.n286 B.n285 585
R184 B.n287 B.n62 585
R185 B.n289 B.n288 585
R186 B.n290 B.n61 585
R187 B.n292 B.n291 585
R188 B.n293 B.n60 585
R189 B.n295 B.n294 585
R190 B.n296 B.n59 585
R191 B.n298 B.n297 585
R192 B.n299 B.n58 585
R193 B.n301 B.n300 585
R194 B.n302 B.n57 585
R195 B.n304 B.n303 585
R196 B.n305 B.n56 585
R197 B.n307 B.n306 585
R198 B.n308 B.n55 585
R199 B.n310 B.n309 585
R200 B.n311 B.n54 585
R201 B.n313 B.n312 585
R202 B.n314 B.n53 585
R203 B.n316 B.n315 585
R204 B.n317 B.n52 585
R205 B.n319 B.n318 585
R206 B.n320 B.n51 585
R207 B.n322 B.n321 585
R208 B.n323 B.n50 585
R209 B.n325 B.n324 585
R210 B.n326 B.n49 585
R211 B.n328 B.n327 585
R212 B.n329 B.n48 585
R213 B.n331 B.n330 585
R214 B.n332 B.n47 585
R215 B.n334 B.n333 585
R216 B.n410 B.n17 585
R217 B.n409 B.n408 585
R218 B.n407 B.n18 585
R219 B.n406 B.n405 585
R220 B.n404 B.n19 585
R221 B.n403 B.n402 585
R222 B.n401 B.n20 585
R223 B.n400 B.n399 585
R224 B.n398 B.n21 585
R225 B.n397 B.n396 585
R226 B.n395 B.n22 585
R227 B.n394 B.n393 585
R228 B.n392 B.n23 585
R229 B.n391 B.n390 585
R230 B.n389 B.n24 585
R231 B.n388 B.n387 585
R232 B.n386 B.n25 585
R233 B.n385 B.n384 585
R234 B.n383 B.n26 585
R235 B.n382 B.n381 585
R236 B.n379 B.n27 585
R237 B.n378 B.n377 585
R238 B.n376 B.n30 585
R239 B.n375 B.n374 585
R240 B.n373 B.n31 585
R241 B.n372 B.n371 585
R242 B.n370 B.n32 585
R243 B.n369 B.n368 585
R244 B.n367 B.n33 585
R245 B.n366 B.n365 585
R246 B.n364 B.n363 585
R247 B.n362 B.n37 585
R248 B.n361 B.n360 585
R249 B.n359 B.n38 585
R250 B.n358 B.n357 585
R251 B.n356 B.n39 585
R252 B.n355 B.n354 585
R253 B.n353 B.n40 585
R254 B.n352 B.n351 585
R255 B.n350 B.n41 585
R256 B.n349 B.n348 585
R257 B.n347 B.n42 585
R258 B.n346 B.n345 585
R259 B.n344 B.n43 585
R260 B.n343 B.n342 585
R261 B.n341 B.n44 585
R262 B.n340 B.n339 585
R263 B.n338 B.n45 585
R264 B.n337 B.n336 585
R265 B.n335 B.n46 585
R266 B.n412 B.n411 585
R267 B.n413 B.n16 585
R268 B.n415 B.n414 585
R269 B.n416 B.n15 585
R270 B.n418 B.n417 585
R271 B.n419 B.n14 585
R272 B.n421 B.n420 585
R273 B.n422 B.n13 585
R274 B.n424 B.n423 585
R275 B.n425 B.n12 585
R276 B.n427 B.n426 585
R277 B.n428 B.n11 585
R278 B.n430 B.n429 585
R279 B.n431 B.n10 585
R280 B.n433 B.n432 585
R281 B.n434 B.n9 585
R282 B.n436 B.n435 585
R283 B.n437 B.n8 585
R284 B.n439 B.n438 585
R285 B.n440 B.n7 585
R286 B.n442 B.n441 585
R287 B.n443 B.n6 585
R288 B.n445 B.n444 585
R289 B.n446 B.n5 585
R290 B.n448 B.n447 585
R291 B.n449 B.n4 585
R292 B.n451 B.n450 585
R293 B.n452 B.n3 585
R294 B.n454 B.n453 585
R295 B.n455 B.n0 585
R296 B.n2 B.n1 585
R297 B.n120 B.n119 585
R298 B.n121 B.n118 585
R299 B.n123 B.n122 585
R300 B.n124 B.n117 585
R301 B.n126 B.n125 585
R302 B.n127 B.n116 585
R303 B.n129 B.n128 585
R304 B.n130 B.n115 585
R305 B.n132 B.n131 585
R306 B.n133 B.n114 585
R307 B.n135 B.n134 585
R308 B.n136 B.n113 585
R309 B.n138 B.n137 585
R310 B.n139 B.n112 585
R311 B.n141 B.n140 585
R312 B.n142 B.n111 585
R313 B.n144 B.n143 585
R314 B.n145 B.n110 585
R315 B.n147 B.n146 585
R316 B.n148 B.n109 585
R317 B.n150 B.n149 585
R318 B.n151 B.n108 585
R319 B.n153 B.n152 585
R320 B.n154 B.n107 585
R321 B.n156 B.n155 585
R322 B.n157 B.n106 585
R323 B.n159 B.n158 585
R324 B.n160 B.n105 585
R325 B.n162 B.n161 585
R326 B.n163 B.n162 550.159
R327 B.n240 B.n77 550.159
R328 B.n335 B.n334 550.159
R329 B.n412 B.n17 550.159
R330 B.n191 B.t9 300.315
R331 B.n88 B.t6 300.315
R332 B.n34 B.t3 300.315
R333 B.n28 B.t0 300.315
R334 B.n457 B.n456 256.663
R335 B.n456 B.n455 235.042
R336 B.n456 B.n2 235.042
R337 B.n164 B.n163 163.367
R338 B.n164 B.n103 163.367
R339 B.n168 B.n103 163.367
R340 B.n169 B.n168 163.367
R341 B.n170 B.n169 163.367
R342 B.n170 B.n101 163.367
R343 B.n174 B.n101 163.367
R344 B.n175 B.n174 163.367
R345 B.n176 B.n175 163.367
R346 B.n176 B.n99 163.367
R347 B.n180 B.n99 163.367
R348 B.n181 B.n180 163.367
R349 B.n182 B.n181 163.367
R350 B.n182 B.n97 163.367
R351 B.n186 B.n97 163.367
R352 B.n187 B.n186 163.367
R353 B.n188 B.n187 163.367
R354 B.n188 B.n95 163.367
R355 B.n195 B.n95 163.367
R356 B.n196 B.n195 163.367
R357 B.n197 B.n196 163.367
R358 B.n197 B.n93 163.367
R359 B.n201 B.n93 163.367
R360 B.n202 B.n201 163.367
R361 B.n203 B.n202 163.367
R362 B.n203 B.n91 163.367
R363 B.n207 B.n91 163.367
R364 B.n208 B.n207 163.367
R365 B.n209 B.n208 163.367
R366 B.n209 B.n87 163.367
R367 B.n214 B.n87 163.367
R368 B.n215 B.n214 163.367
R369 B.n216 B.n215 163.367
R370 B.n216 B.n85 163.367
R371 B.n220 B.n85 163.367
R372 B.n221 B.n220 163.367
R373 B.n222 B.n221 163.367
R374 B.n222 B.n83 163.367
R375 B.n226 B.n83 163.367
R376 B.n227 B.n226 163.367
R377 B.n228 B.n227 163.367
R378 B.n228 B.n81 163.367
R379 B.n232 B.n81 163.367
R380 B.n233 B.n232 163.367
R381 B.n234 B.n233 163.367
R382 B.n234 B.n79 163.367
R383 B.n238 B.n79 163.367
R384 B.n239 B.n238 163.367
R385 B.n240 B.n239 163.367
R386 B.n334 B.n47 163.367
R387 B.n330 B.n47 163.367
R388 B.n330 B.n329 163.367
R389 B.n329 B.n328 163.367
R390 B.n328 B.n49 163.367
R391 B.n324 B.n49 163.367
R392 B.n324 B.n323 163.367
R393 B.n323 B.n322 163.367
R394 B.n322 B.n51 163.367
R395 B.n318 B.n51 163.367
R396 B.n318 B.n317 163.367
R397 B.n317 B.n316 163.367
R398 B.n316 B.n53 163.367
R399 B.n312 B.n53 163.367
R400 B.n312 B.n311 163.367
R401 B.n311 B.n310 163.367
R402 B.n310 B.n55 163.367
R403 B.n306 B.n55 163.367
R404 B.n306 B.n305 163.367
R405 B.n305 B.n304 163.367
R406 B.n304 B.n57 163.367
R407 B.n300 B.n57 163.367
R408 B.n300 B.n299 163.367
R409 B.n299 B.n298 163.367
R410 B.n298 B.n59 163.367
R411 B.n294 B.n59 163.367
R412 B.n294 B.n293 163.367
R413 B.n293 B.n292 163.367
R414 B.n292 B.n61 163.367
R415 B.n288 B.n61 163.367
R416 B.n288 B.n287 163.367
R417 B.n287 B.n286 163.367
R418 B.n286 B.n63 163.367
R419 B.n282 B.n63 163.367
R420 B.n282 B.n281 163.367
R421 B.n281 B.n280 163.367
R422 B.n280 B.n65 163.367
R423 B.n276 B.n65 163.367
R424 B.n276 B.n275 163.367
R425 B.n275 B.n274 163.367
R426 B.n274 B.n67 163.367
R427 B.n270 B.n67 163.367
R428 B.n270 B.n269 163.367
R429 B.n269 B.n268 163.367
R430 B.n268 B.n69 163.367
R431 B.n264 B.n69 163.367
R432 B.n264 B.n263 163.367
R433 B.n263 B.n262 163.367
R434 B.n262 B.n71 163.367
R435 B.n258 B.n71 163.367
R436 B.n258 B.n257 163.367
R437 B.n257 B.n256 163.367
R438 B.n256 B.n73 163.367
R439 B.n252 B.n73 163.367
R440 B.n252 B.n251 163.367
R441 B.n251 B.n250 163.367
R442 B.n250 B.n75 163.367
R443 B.n246 B.n75 163.367
R444 B.n246 B.n245 163.367
R445 B.n245 B.n244 163.367
R446 B.n244 B.n77 163.367
R447 B.n408 B.n17 163.367
R448 B.n408 B.n407 163.367
R449 B.n407 B.n406 163.367
R450 B.n406 B.n19 163.367
R451 B.n402 B.n19 163.367
R452 B.n402 B.n401 163.367
R453 B.n401 B.n400 163.367
R454 B.n400 B.n21 163.367
R455 B.n396 B.n21 163.367
R456 B.n396 B.n395 163.367
R457 B.n395 B.n394 163.367
R458 B.n394 B.n23 163.367
R459 B.n390 B.n23 163.367
R460 B.n390 B.n389 163.367
R461 B.n389 B.n388 163.367
R462 B.n388 B.n25 163.367
R463 B.n384 B.n25 163.367
R464 B.n384 B.n383 163.367
R465 B.n383 B.n382 163.367
R466 B.n382 B.n27 163.367
R467 B.n377 B.n27 163.367
R468 B.n377 B.n376 163.367
R469 B.n376 B.n375 163.367
R470 B.n375 B.n31 163.367
R471 B.n371 B.n31 163.367
R472 B.n371 B.n370 163.367
R473 B.n370 B.n369 163.367
R474 B.n369 B.n33 163.367
R475 B.n365 B.n33 163.367
R476 B.n365 B.n364 163.367
R477 B.n364 B.n37 163.367
R478 B.n360 B.n37 163.367
R479 B.n360 B.n359 163.367
R480 B.n359 B.n358 163.367
R481 B.n358 B.n39 163.367
R482 B.n354 B.n39 163.367
R483 B.n354 B.n353 163.367
R484 B.n353 B.n352 163.367
R485 B.n352 B.n41 163.367
R486 B.n348 B.n41 163.367
R487 B.n348 B.n347 163.367
R488 B.n347 B.n346 163.367
R489 B.n346 B.n43 163.367
R490 B.n342 B.n43 163.367
R491 B.n342 B.n341 163.367
R492 B.n341 B.n340 163.367
R493 B.n340 B.n45 163.367
R494 B.n336 B.n45 163.367
R495 B.n336 B.n335 163.367
R496 B.n413 B.n412 163.367
R497 B.n414 B.n413 163.367
R498 B.n414 B.n15 163.367
R499 B.n418 B.n15 163.367
R500 B.n419 B.n418 163.367
R501 B.n420 B.n419 163.367
R502 B.n420 B.n13 163.367
R503 B.n424 B.n13 163.367
R504 B.n425 B.n424 163.367
R505 B.n426 B.n425 163.367
R506 B.n426 B.n11 163.367
R507 B.n430 B.n11 163.367
R508 B.n431 B.n430 163.367
R509 B.n432 B.n431 163.367
R510 B.n432 B.n9 163.367
R511 B.n436 B.n9 163.367
R512 B.n437 B.n436 163.367
R513 B.n438 B.n437 163.367
R514 B.n438 B.n7 163.367
R515 B.n442 B.n7 163.367
R516 B.n443 B.n442 163.367
R517 B.n444 B.n443 163.367
R518 B.n444 B.n5 163.367
R519 B.n448 B.n5 163.367
R520 B.n449 B.n448 163.367
R521 B.n450 B.n449 163.367
R522 B.n450 B.n3 163.367
R523 B.n454 B.n3 163.367
R524 B.n455 B.n454 163.367
R525 B.n120 B.n2 163.367
R526 B.n121 B.n120 163.367
R527 B.n122 B.n121 163.367
R528 B.n122 B.n117 163.367
R529 B.n126 B.n117 163.367
R530 B.n127 B.n126 163.367
R531 B.n128 B.n127 163.367
R532 B.n128 B.n115 163.367
R533 B.n132 B.n115 163.367
R534 B.n133 B.n132 163.367
R535 B.n134 B.n133 163.367
R536 B.n134 B.n113 163.367
R537 B.n138 B.n113 163.367
R538 B.n139 B.n138 163.367
R539 B.n140 B.n139 163.367
R540 B.n140 B.n111 163.367
R541 B.n144 B.n111 163.367
R542 B.n145 B.n144 163.367
R543 B.n146 B.n145 163.367
R544 B.n146 B.n109 163.367
R545 B.n150 B.n109 163.367
R546 B.n151 B.n150 163.367
R547 B.n152 B.n151 163.367
R548 B.n152 B.n107 163.367
R549 B.n156 B.n107 163.367
R550 B.n157 B.n156 163.367
R551 B.n158 B.n157 163.367
R552 B.n158 B.n105 163.367
R553 B.n162 B.n105 163.367
R554 B.n88 B.t7 145.06
R555 B.n34 B.t5 145.06
R556 B.n191 B.t10 145.054
R557 B.n28 B.t2 145.054
R558 B.n89 B.t8 115.386
R559 B.n35 B.t4 115.386
R560 B.n192 B.t11 115.382
R561 B.n29 B.t1 115.382
R562 B.n193 B.n192 59.5399
R563 B.n211 B.n89 59.5399
R564 B.n36 B.n35 59.5399
R565 B.n380 B.n29 59.5399
R566 B.n411 B.n410 35.7468
R567 B.n333 B.n46 35.7468
R568 B.n161 B.n104 35.7468
R569 B.n242 B.n241 35.7468
R570 B.n192 B.n191 29.6732
R571 B.n89 B.n88 29.6732
R572 B.n35 B.n34 29.6732
R573 B.n29 B.n28 29.6732
R574 B B.n457 18.0485
R575 B.n411 B.n16 10.6151
R576 B.n415 B.n16 10.6151
R577 B.n416 B.n415 10.6151
R578 B.n417 B.n416 10.6151
R579 B.n417 B.n14 10.6151
R580 B.n421 B.n14 10.6151
R581 B.n422 B.n421 10.6151
R582 B.n423 B.n422 10.6151
R583 B.n423 B.n12 10.6151
R584 B.n427 B.n12 10.6151
R585 B.n428 B.n427 10.6151
R586 B.n429 B.n428 10.6151
R587 B.n429 B.n10 10.6151
R588 B.n433 B.n10 10.6151
R589 B.n434 B.n433 10.6151
R590 B.n435 B.n434 10.6151
R591 B.n435 B.n8 10.6151
R592 B.n439 B.n8 10.6151
R593 B.n440 B.n439 10.6151
R594 B.n441 B.n440 10.6151
R595 B.n441 B.n6 10.6151
R596 B.n445 B.n6 10.6151
R597 B.n446 B.n445 10.6151
R598 B.n447 B.n446 10.6151
R599 B.n447 B.n4 10.6151
R600 B.n451 B.n4 10.6151
R601 B.n452 B.n451 10.6151
R602 B.n453 B.n452 10.6151
R603 B.n453 B.n0 10.6151
R604 B.n410 B.n409 10.6151
R605 B.n409 B.n18 10.6151
R606 B.n405 B.n18 10.6151
R607 B.n405 B.n404 10.6151
R608 B.n404 B.n403 10.6151
R609 B.n403 B.n20 10.6151
R610 B.n399 B.n20 10.6151
R611 B.n399 B.n398 10.6151
R612 B.n398 B.n397 10.6151
R613 B.n397 B.n22 10.6151
R614 B.n393 B.n22 10.6151
R615 B.n393 B.n392 10.6151
R616 B.n392 B.n391 10.6151
R617 B.n391 B.n24 10.6151
R618 B.n387 B.n24 10.6151
R619 B.n387 B.n386 10.6151
R620 B.n386 B.n385 10.6151
R621 B.n385 B.n26 10.6151
R622 B.n381 B.n26 10.6151
R623 B.n379 B.n378 10.6151
R624 B.n378 B.n30 10.6151
R625 B.n374 B.n30 10.6151
R626 B.n374 B.n373 10.6151
R627 B.n373 B.n372 10.6151
R628 B.n372 B.n32 10.6151
R629 B.n368 B.n32 10.6151
R630 B.n368 B.n367 10.6151
R631 B.n367 B.n366 10.6151
R632 B.n363 B.n362 10.6151
R633 B.n362 B.n361 10.6151
R634 B.n361 B.n38 10.6151
R635 B.n357 B.n38 10.6151
R636 B.n357 B.n356 10.6151
R637 B.n356 B.n355 10.6151
R638 B.n355 B.n40 10.6151
R639 B.n351 B.n40 10.6151
R640 B.n351 B.n350 10.6151
R641 B.n350 B.n349 10.6151
R642 B.n349 B.n42 10.6151
R643 B.n345 B.n42 10.6151
R644 B.n345 B.n344 10.6151
R645 B.n344 B.n343 10.6151
R646 B.n343 B.n44 10.6151
R647 B.n339 B.n44 10.6151
R648 B.n339 B.n338 10.6151
R649 B.n338 B.n337 10.6151
R650 B.n337 B.n46 10.6151
R651 B.n333 B.n332 10.6151
R652 B.n332 B.n331 10.6151
R653 B.n331 B.n48 10.6151
R654 B.n327 B.n48 10.6151
R655 B.n327 B.n326 10.6151
R656 B.n326 B.n325 10.6151
R657 B.n325 B.n50 10.6151
R658 B.n321 B.n50 10.6151
R659 B.n321 B.n320 10.6151
R660 B.n320 B.n319 10.6151
R661 B.n319 B.n52 10.6151
R662 B.n315 B.n52 10.6151
R663 B.n315 B.n314 10.6151
R664 B.n314 B.n313 10.6151
R665 B.n313 B.n54 10.6151
R666 B.n309 B.n54 10.6151
R667 B.n309 B.n308 10.6151
R668 B.n308 B.n307 10.6151
R669 B.n307 B.n56 10.6151
R670 B.n303 B.n56 10.6151
R671 B.n303 B.n302 10.6151
R672 B.n302 B.n301 10.6151
R673 B.n301 B.n58 10.6151
R674 B.n297 B.n58 10.6151
R675 B.n297 B.n296 10.6151
R676 B.n296 B.n295 10.6151
R677 B.n295 B.n60 10.6151
R678 B.n291 B.n60 10.6151
R679 B.n291 B.n290 10.6151
R680 B.n290 B.n289 10.6151
R681 B.n289 B.n62 10.6151
R682 B.n285 B.n62 10.6151
R683 B.n285 B.n284 10.6151
R684 B.n284 B.n283 10.6151
R685 B.n283 B.n64 10.6151
R686 B.n279 B.n64 10.6151
R687 B.n279 B.n278 10.6151
R688 B.n278 B.n277 10.6151
R689 B.n277 B.n66 10.6151
R690 B.n273 B.n66 10.6151
R691 B.n273 B.n272 10.6151
R692 B.n272 B.n271 10.6151
R693 B.n271 B.n68 10.6151
R694 B.n267 B.n68 10.6151
R695 B.n267 B.n266 10.6151
R696 B.n266 B.n265 10.6151
R697 B.n265 B.n70 10.6151
R698 B.n261 B.n70 10.6151
R699 B.n261 B.n260 10.6151
R700 B.n260 B.n259 10.6151
R701 B.n259 B.n72 10.6151
R702 B.n255 B.n72 10.6151
R703 B.n255 B.n254 10.6151
R704 B.n254 B.n253 10.6151
R705 B.n253 B.n74 10.6151
R706 B.n249 B.n74 10.6151
R707 B.n249 B.n248 10.6151
R708 B.n248 B.n247 10.6151
R709 B.n247 B.n76 10.6151
R710 B.n243 B.n76 10.6151
R711 B.n243 B.n242 10.6151
R712 B.n119 B.n1 10.6151
R713 B.n119 B.n118 10.6151
R714 B.n123 B.n118 10.6151
R715 B.n124 B.n123 10.6151
R716 B.n125 B.n124 10.6151
R717 B.n125 B.n116 10.6151
R718 B.n129 B.n116 10.6151
R719 B.n130 B.n129 10.6151
R720 B.n131 B.n130 10.6151
R721 B.n131 B.n114 10.6151
R722 B.n135 B.n114 10.6151
R723 B.n136 B.n135 10.6151
R724 B.n137 B.n136 10.6151
R725 B.n137 B.n112 10.6151
R726 B.n141 B.n112 10.6151
R727 B.n142 B.n141 10.6151
R728 B.n143 B.n142 10.6151
R729 B.n143 B.n110 10.6151
R730 B.n147 B.n110 10.6151
R731 B.n148 B.n147 10.6151
R732 B.n149 B.n148 10.6151
R733 B.n149 B.n108 10.6151
R734 B.n153 B.n108 10.6151
R735 B.n154 B.n153 10.6151
R736 B.n155 B.n154 10.6151
R737 B.n155 B.n106 10.6151
R738 B.n159 B.n106 10.6151
R739 B.n160 B.n159 10.6151
R740 B.n161 B.n160 10.6151
R741 B.n165 B.n104 10.6151
R742 B.n166 B.n165 10.6151
R743 B.n167 B.n166 10.6151
R744 B.n167 B.n102 10.6151
R745 B.n171 B.n102 10.6151
R746 B.n172 B.n171 10.6151
R747 B.n173 B.n172 10.6151
R748 B.n173 B.n100 10.6151
R749 B.n177 B.n100 10.6151
R750 B.n178 B.n177 10.6151
R751 B.n179 B.n178 10.6151
R752 B.n179 B.n98 10.6151
R753 B.n183 B.n98 10.6151
R754 B.n184 B.n183 10.6151
R755 B.n185 B.n184 10.6151
R756 B.n185 B.n96 10.6151
R757 B.n189 B.n96 10.6151
R758 B.n190 B.n189 10.6151
R759 B.n194 B.n190 10.6151
R760 B.n198 B.n94 10.6151
R761 B.n199 B.n198 10.6151
R762 B.n200 B.n199 10.6151
R763 B.n200 B.n92 10.6151
R764 B.n204 B.n92 10.6151
R765 B.n205 B.n204 10.6151
R766 B.n206 B.n205 10.6151
R767 B.n206 B.n90 10.6151
R768 B.n210 B.n90 10.6151
R769 B.n213 B.n212 10.6151
R770 B.n213 B.n86 10.6151
R771 B.n217 B.n86 10.6151
R772 B.n218 B.n217 10.6151
R773 B.n219 B.n218 10.6151
R774 B.n219 B.n84 10.6151
R775 B.n223 B.n84 10.6151
R776 B.n224 B.n223 10.6151
R777 B.n225 B.n224 10.6151
R778 B.n225 B.n82 10.6151
R779 B.n229 B.n82 10.6151
R780 B.n230 B.n229 10.6151
R781 B.n231 B.n230 10.6151
R782 B.n231 B.n80 10.6151
R783 B.n235 B.n80 10.6151
R784 B.n236 B.n235 10.6151
R785 B.n237 B.n236 10.6151
R786 B.n237 B.n78 10.6151
R787 B.n241 B.n78 10.6151
R788 B.n381 B.n380 9.36635
R789 B.n363 B.n36 9.36635
R790 B.n194 B.n193 9.36635
R791 B.n212 B.n211 9.36635
R792 B.n457 B.n0 8.11757
R793 B.n457 B.n1 8.11757
R794 B.n380 B.n379 1.24928
R795 B.n366 B.n36 1.24928
R796 B.n193 B.n94 1.24928
R797 B.n211 B.n210 1.24928
R798 VN.n27 VN.n15 161.3
R799 VN.n26 VN.n25 161.3
R800 VN.n24 VN.n23 161.3
R801 VN.n22 VN.n17 161.3
R802 VN.n21 VN.n20 161.3
R803 VN.n12 VN.n0 161.3
R804 VN.n11 VN.n10 161.3
R805 VN.n9 VN.n8 161.3
R806 VN.n7 VN.n2 161.3
R807 VN.n6 VN.n5 161.3
R808 VN.n4 VN.t5 147.639
R809 VN.n19 VN.t2 147.639
R810 VN.n13 VN.t0 129.137
R811 VN.n28 VN.t7 129.137
R812 VN.n3 VN.t3 96.1997
R813 VN.n1 VN.t1 96.1997
R814 VN.n18 VN.t4 96.1997
R815 VN.n16 VN.t6 96.1997
R816 VN.n29 VN.n28 80.6037
R817 VN.n14 VN.n13 80.6037
R818 VN.n4 VN.n3 44.8004
R819 VN.n19 VN.n18 44.8004
R820 VN.n7 VN.n6 40.4934
R821 VN.n8 VN.n7 40.4934
R822 VN.n22 VN.n21 40.4934
R823 VN.n23 VN.n22 40.4934
R824 VN VN.n29 39.2794
R825 VN.n12 VN.n11 37.5796
R826 VN.n27 VN.n26 37.5796
R827 VN.n20 VN.n19 29.7304
R828 VN.n5 VN.n4 29.7304
R829 VN.n13 VN.n12 28.4823
R830 VN.n28 VN.n27 28.4823
R831 VN.n6 VN.n3 12.968
R832 VN.n8 VN.n1 12.968
R833 VN.n21 VN.n18 12.968
R834 VN.n23 VN.n16 12.968
R835 VN.n11 VN.n1 11.5
R836 VN.n26 VN.n16 11.5
R837 VN.n29 VN.n15 0.285035
R838 VN.n14 VN.n0 0.285035
R839 VN.n25 VN.n15 0.189894
R840 VN.n25 VN.n24 0.189894
R841 VN.n24 VN.n17 0.189894
R842 VN.n20 VN.n17 0.189894
R843 VN.n5 VN.n2 0.189894
R844 VN.n9 VN.n2 0.189894
R845 VN.n10 VN.n9 0.189894
R846 VN.n10 VN.n0 0.189894
R847 VN VN.n14 0.146778
R848 VDD2.n2 VDD2.n1 104.579
R849 VDD2.n2 VDD2.n0 104.579
R850 VDD2 VDD2.n5 104.576
R851 VDD2.n4 VDD2.n3 103.975
R852 VDD2.n4 VDD2.n2 33.7799
R853 VDD2.n5 VDD2.t3 6.78651
R854 VDD2.n5 VDD2.t5 6.78651
R855 VDD2.n3 VDD2.t0 6.78651
R856 VDD2.n3 VDD2.t1 6.78651
R857 VDD2.n1 VDD2.t6 6.78651
R858 VDD2.n1 VDD2.t7 6.78651
R859 VDD2.n0 VDD2.t2 6.78651
R860 VDD2.n0 VDD2.t4 6.78651
R861 VDD2 VDD2.n4 0.718172
C0 VDD2 VP 0.374501f
C1 w_n2500_n1926# VDD2 1.34081f
C2 VP VN 4.61669f
C3 w_n2500_n1926# VN 4.5722f
C4 VDD1 B 1.02848f
C5 VDD1 VDD2 1.07356f
C6 B VDD2 1.08068f
C7 VDD1 VN 0.152624f
C8 B VN 0.8256f
C9 VTAIL VP 3.38941f
C10 w_n2500_n1926# VTAIL 2.40775f
C11 VDD2 VN 3.05038f
C12 w_n2500_n1926# VP 4.892529f
C13 VDD1 VTAIL 5.16058f
C14 VTAIL B 2.10076f
C15 VDD1 VP 3.27114f
C16 B VP 1.3552f
C17 VDD1 w_n2500_n1926# 1.28528f
C18 w_n2500_n1926# B 5.95454f
C19 VTAIL VDD2 5.20561f
C20 VTAIL VN 3.3753f
C21 VDD2 VSUBS 1.134527f
C22 VDD1 VSUBS 1.535399f
C23 VTAIL VSUBS 0.530948f
C24 VN VSUBS 4.69432f
C25 VP VSUBS 1.7705f
C26 B VSUBS 2.698106f
C27 w_n2500_n1926# VSUBS 60.39f
C28 VDD2.t2 VSUBS 0.095779f
C29 VDD2.t4 VSUBS 0.095779f
C30 VDD2.n0 VSUBS 0.613467f
C31 VDD2.t6 VSUBS 0.095779f
C32 VDD2.t7 VSUBS 0.095779f
C33 VDD2.n1 VSUBS 0.613467f
C34 VDD2.n2 VSUBS 2.37026f
C35 VDD2.t0 VSUBS 0.095779f
C36 VDD2.t1 VSUBS 0.095779f
C37 VDD2.n3 VSUBS 0.610387f
C38 VDD2.n4 VSUBS 2.07615f
C39 VDD2.t3 VSUBS 0.095779f
C40 VDD2.t5 VSUBS 0.095779f
C41 VDD2.n5 VSUBS 0.613443f
C42 VN.n0 VSUBS 0.070797f
C43 VN.t1 VSUBS 0.795181f
C44 VN.n1 VSUBS 0.3337f
C45 VN.n2 VSUBS 0.053056f
C46 VN.t3 VSUBS 0.795181f
C47 VN.n3 VSUBS 0.400975f
C48 VN.t5 VSUBS 0.948216f
C49 VN.n4 VSUBS 0.422098f
C50 VN.n5 VSUBS 0.272357f
C51 VN.n6 VSUBS 0.082501f
C52 VN.n7 VSUBS 0.042891f
C53 VN.n8 VSUBS 0.082501f
C54 VN.n9 VSUBS 0.053056f
C55 VN.n10 VSUBS 0.053056f
C56 VN.n11 VSUBS 0.080838f
C57 VN.n12 VSUBS 0.031076f
C58 VN.t0 VSUBS 0.89272f
C59 VN.n13 VSUBS 0.430546f
C60 VN.n14 VSUBS 0.049689f
C61 VN.n15 VSUBS 0.070797f
C62 VN.t6 VSUBS 0.795181f
C63 VN.n16 VSUBS 0.3337f
C64 VN.n17 VSUBS 0.053056f
C65 VN.t4 VSUBS 0.795181f
C66 VN.n18 VSUBS 0.400975f
C67 VN.t2 VSUBS 0.948216f
C68 VN.n19 VSUBS 0.422098f
C69 VN.n20 VSUBS 0.272357f
C70 VN.n21 VSUBS 0.082501f
C71 VN.n22 VSUBS 0.042891f
C72 VN.n23 VSUBS 0.082501f
C73 VN.n24 VSUBS 0.053056f
C74 VN.n25 VSUBS 0.053056f
C75 VN.n26 VSUBS 0.080838f
C76 VN.n27 VSUBS 0.031076f
C77 VN.t7 VSUBS 0.89272f
C78 VN.n28 VSUBS 0.430546f
C79 VN.n29 VSUBS 1.97768f
C80 B.n0 VSUBS 0.008169f
C81 B.n1 VSUBS 0.008169f
C82 B.n2 VSUBS 0.012082f
C83 B.n3 VSUBS 0.009259f
C84 B.n4 VSUBS 0.009259f
C85 B.n5 VSUBS 0.009259f
C86 B.n6 VSUBS 0.009259f
C87 B.n7 VSUBS 0.009259f
C88 B.n8 VSUBS 0.009259f
C89 B.n9 VSUBS 0.009259f
C90 B.n10 VSUBS 0.009259f
C91 B.n11 VSUBS 0.009259f
C92 B.n12 VSUBS 0.009259f
C93 B.n13 VSUBS 0.009259f
C94 B.n14 VSUBS 0.009259f
C95 B.n15 VSUBS 0.009259f
C96 B.n16 VSUBS 0.009259f
C97 B.n17 VSUBS 0.023413f
C98 B.n18 VSUBS 0.009259f
C99 B.n19 VSUBS 0.009259f
C100 B.n20 VSUBS 0.009259f
C101 B.n21 VSUBS 0.009259f
C102 B.n22 VSUBS 0.009259f
C103 B.n23 VSUBS 0.009259f
C104 B.n24 VSUBS 0.009259f
C105 B.n25 VSUBS 0.009259f
C106 B.n26 VSUBS 0.009259f
C107 B.n27 VSUBS 0.009259f
C108 B.t1 VSUBS 0.175225f
C109 B.t2 VSUBS 0.189814f
C110 B.t0 VSUBS 0.348285f
C111 B.n28 VSUBS 0.114211f
C112 B.n29 VSUBS 0.084521f
C113 B.n30 VSUBS 0.009259f
C114 B.n31 VSUBS 0.009259f
C115 B.n32 VSUBS 0.009259f
C116 B.n33 VSUBS 0.009259f
C117 B.t4 VSUBS 0.175225f
C118 B.t5 VSUBS 0.189813f
C119 B.t3 VSUBS 0.348285f
C120 B.n34 VSUBS 0.114211f
C121 B.n35 VSUBS 0.084521f
C122 B.n36 VSUBS 0.021451f
C123 B.n37 VSUBS 0.009259f
C124 B.n38 VSUBS 0.009259f
C125 B.n39 VSUBS 0.009259f
C126 B.n40 VSUBS 0.009259f
C127 B.n41 VSUBS 0.009259f
C128 B.n42 VSUBS 0.009259f
C129 B.n43 VSUBS 0.009259f
C130 B.n44 VSUBS 0.009259f
C131 B.n45 VSUBS 0.009259f
C132 B.n46 VSUBS 0.023413f
C133 B.n47 VSUBS 0.009259f
C134 B.n48 VSUBS 0.009259f
C135 B.n49 VSUBS 0.009259f
C136 B.n50 VSUBS 0.009259f
C137 B.n51 VSUBS 0.009259f
C138 B.n52 VSUBS 0.009259f
C139 B.n53 VSUBS 0.009259f
C140 B.n54 VSUBS 0.009259f
C141 B.n55 VSUBS 0.009259f
C142 B.n56 VSUBS 0.009259f
C143 B.n57 VSUBS 0.009259f
C144 B.n58 VSUBS 0.009259f
C145 B.n59 VSUBS 0.009259f
C146 B.n60 VSUBS 0.009259f
C147 B.n61 VSUBS 0.009259f
C148 B.n62 VSUBS 0.009259f
C149 B.n63 VSUBS 0.009259f
C150 B.n64 VSUBS 0.009259f
C151 B.n65 VSUBS 0.009259f
C152 B.n66 VSUBS 0.009259f
C153 B.n67 VSUBS 0.009259f
C154 B.n68 VSUBS 0.009259f
C155 B.n69 VSUBS 0.009259f
C156 B.n70 VSUBS 0.009259f
C157 B.n71 VSUBS 0.009259f
C158 B.n72 VSUBS 0.009259f
C159 B.n73 VSUBS 0.009259f
C160 B.n74 VSUBS 0.009259f
C161 B.n75 VSUBS 0.009259f
C162 B.n76 VSUBS 0.009259f
C163 B.n77 VSUBS 0.022608f
C164 B.n78 VSUBS 0.009259f
C165 B.n79 VSUBS 0.009259f
C166 B.n80 VSUBS 0.009259f
C167 B.n81 VSUBS 0.009259f
C168 B.n82 VSUBS 0.009259f
C169 B.n83 VSUBS 0.009259f
C170 B.n84 VSUBS 0.009259f
C171 B.n85 VSUBS 0.009259f
C172 B.n86 VSUBS 0.009259f
C173 B.n87 VSUBS 0.009259f
C174 B.t8 VSUBS 0.175225f
C175 B.t7 VSUBS 0.189813f
C176 B.t6 VSUBS 0.348285f
C177 B.n88 VSUBS 0.114211f
C178 B.n89 VSUBS 0.084521f
C179 B.n90 VSUBS 0.009259f
C180 B.n91 VSUBS 0.009259f
C181 B.n92 VSUBS 0.009259f
C182 B.n93 VSUBS 0.009259f
C183 B.n94 VSUBS 0.005174f
C184 B.n95 VSUBS 0.009259f
C185 B.n96 VSUBS 0.009259f
C186 B.n97 VSUBS 0.009259f
C187 B.n98 VSUBS 0.009259f
C188 B.n99 VSUBS 0.009259f
C189 B.n100 VSUBS 0.009259f
C190 B.n101 VSUBS 0.009259f
C191 B.n102 VSUBS 0.009259f
C192 B.n103 VSUBS 0.009259f
C193 B.n104 VSUBS 0.023413f
C194 B.n105 VSUBS 0.009259f
C195 B.n106 VSUBS 0.009259f
C196 B.n107 VSUBS 0.009259f
C197 B.n108 VSUBS 0.009259f
C198 B.n109 VSUBS 0.009259f
C199 B.n110 VSUBS 0.009259f
C200 B.n111 VSUBS 0.009259f
C201 B.n112 VSUBS 0.009259f
C202 B.n113 VSUBS 0.009259f
C203 B.n114 VSUBS 0.009259f
C204 B.n115 VSUBS 0.009259f
C205 B.n116 VSUBS 0.009259f
C206 B.n117 VSUBS 0.009259f
C207 B.n118 VSUBS 0.009259f
C208 B.n119 VSUBS 0.009259f
C209 B.n120 VSUBS 0.009259f
C210 B.n121 VSUBS 0.009259f
C211 B.n122 VSUBS 0.009259f
C212 B.n123 VSUBS 0.009259f
C213 B.n124 VSUBS 0.009259f
C214 B.n125 VSUBS 0.009259f
C215 B.n126 VSUBS 0.009259f
C216 B.n127 VSUBS 0.009259f
C217 B.n128 VSUBS 0.009259f
C218 B.n129 VSUBS 0.009259f
C219 B.n130 VSUBS 0.009259f
C220 B.n131 VSUBS 0.009259f
C221 B.n132 VSUBS 0.009259f
C222 B.n133 VSUBS 0.009259f
C223 B.n134 VSUBS 0.009259f
C224 B.n135 VSUBS 0.009259f
C225 B.n136 VSUBS 0.009259f
C226 B.n137 VSUBS 0.009259f
C227 B.n138 VSUBS 0.009259f
C228 B.n139 VSUBS 0.009259f
C229 B.n140 VSUBS 0.009259f
C230 B.n141 VSUBS 0.009259f
C231 B.n142 VSUBS 0.009259f
C232 B.n143 VSUBS 0.009259f
C233 B.n144 VSUBS 0.009259f
C234 B.n145 VSUBS 0.009259f
C235 B.n146 VSUBS 0.009259f
C236 B.n147 VSUBS 0.009259f
C237 B.n148 VSUBS 0.009259f
C238 B.n149 VSUBS 0.009259f
C239 B.n150 VSUBS 0.009259f
C240 B.n151 VSUBS 0.009259f
C241 B.n152 VSUBS 0.009259f
C242 B.n153 VSUBS 0.009259f
C243 B.n154 VSUBS 0.009259f
C244 B.n155 VSUBS 0.009259f
C245 B.n156 VSUBS 0.009259f
C246 B.n157 VSUBS 0.009259f
C247 B.n158 VSUBS 0.009259f
C248 B.n159 VSUBS 0.009259f
C249 B.n160 VSUBS 0.009259f
C250 B.n161 VSUBS 0.022608f
C251 B.n162 VSUBS 0.022608f
C252 B.n163 VSUBS 0.023413f
C253 B.n164 VSUBS 0.009259f
C254 B.n165 VSUBS 0.009259f
C255 B.n166 VSUBS 0.009259f
C256 B.n167 VSUBS 0.009259f
C257 B.n168 VSUBS 0.009259f
C258 B.n169 VSUBS 0.009259f
C259 B.n170 VSUBS 0.009259f
C260 B.n171 VSUBS 0.009259f
C261 B.n172 VSUBS 0.009259f
C262 B.n173 VSUBS 0.009259f
C263 B.n174 VSUBS 0.009259f
C264 B.n175 VSUBS 0.009259f
C265 B.n176 VSUBS 0.009259f
C266 B.n177 VSUBS 0.009259f
C267 B.n178 VSUBS 0.009259f
C268 B.n179 VSUBS 0.009259f
C269 B.n180 VSUBS 0.009259f
C270 B.n181 VSUBS 0.009259f
C271 B.n182 VSUBS 0.009259f
C272 B.n183 VSUBS 0.009259f
C273 B.n184 VSUBS 0.009259f
C274 B.n185 VSUBS 0.009259f
C275 B.n186 VSUBS 0.009259f
C276 B.n187 VSUBS 0.009259f
C277 B.n188 VSUBS 0.009259f
C278 B.n189 VSUBS 0.009259f
C279 B.n190 VSUBS 0.009259f
C280 B.t11 VSUBS 0.175225f
C281 B.t10 VSUBS 0.189814f
C282 B.t9 VSUBS 0.348285f
C283 B.n191 VSUBS 0.114211f
C284 B.n192 VSUBS 0.084521f
C285 B.n193 VSUBS 0.021451f
C286 B.n194 VSUBS 0.008714f
C287 B.n195 VSUBS 0.009259f
C288 B.n196 VSUBS 0.009259f
C289 B.n197 VSUBS 0.009259f
C290 B.n198 VSUBS 0.009259f
C291 B.n199 VSUBS 0.009259f
C292 B.n200 VSUBS 0.009259f
C293 B.n201 VSUBS 0.009259f
C294 B.n202 VSUBS 0.009259f
C295 B.n203 VSUBS 0.009259f
C296 B.n204 VSUBS 0.009259f
C297 B.n205 VSUBS 0.009259f
C298 B.n206 VSUBS 0.009259f
C299 B.n207 VSUBS 0.009259f
C300 B.n208 VSUBS 0.009259f
C301 B.n209 VSUBS 0.009259f
C302 B.n210 VSUBS 0.005174f
C303 B.n211 VSUBS 0.021451f
C304 B.n212 VSUBS 0.008714f
C305 B.n213 VSUBS 0.009259f
C306 B.n214 VSUBS 0.009259f
C307 B.n215 VSUBS 0.009259f
C308 B.n216 VSUBS 0.009259f
C309 B.n217 VSUBS 0.009259f
C310 B.n218 VSUBS 0.009259f
C311 B.n219 VSUBS 0.009259f
C312 B.n220 VSUBS 0.009259f
C313 B.n221 VSUBS 0.009259f
C314 B.n222 VSUBS 0.009259f
C315 B.n223 VSUBS 0.009259f
C316 B.n224 VSUBS 0.009259f
C317 B.n225 VSUBS 0.009259f
C318 B.n226 VSUBS 0.009259f
C319 B.n227 VSUBS 0.009259f
C320 B.n228 VSUBS 0.009259f
C321 B.n229 VSUBS 0.009259f
C322 B.n230 VSUBS 0.009259f
C323 B.n231 VSUBS 0.009259f
C324 B.n232 VSUBS 0.009259f
C325 B.n233 VSUBS 0.009259f
C326 B.n234 VSUBS 0.009259f
C327 B.n235 VSUBS 0.009259f
C328 B.n236 VSUBS 0.009259f
C329 B.n237 VSUBS 0.009259f
C330 B.n238 VSUBS 0.009259f
C331 B.n239 VSUBS 0.009259f
C332 B.n240 VSUBS 0.023413f
C333 B.n241 VSUBS 0.022413f
C334 B.n242 VSUBS 0.023608f
C335 B.n243 VSUBS 0.009259f
C336 B.n244 VSUBS 0.009259f
C337 B.n245 VSUBS 0.009259f
C338 B.n246 VSUBS 0.009259f
C339 B.n247 VSUBS 0.009259f
C340 B.n248 VSUBS 0.009259f
C341 B.n249 VSUBS 0.009259f
C342 B.n250 VSUBS 0.009259f
C343 B.n251 VSUBS 0.009259f
C344 B.n252 VSUBS 0.009259f
C345 B.n253 VSUBS 0.009259f
C346 B.n254 VSUBS 0.009259f
C347 B.n255 VSUBS 0.009259f
C348 B.n256 VSUBS 0.009259f
C349 B.n257 VSUBS 0.009259f
C350 B.n258 VSUBS 0.009259f
C351 B.n259 VSUBS 0.009259f
C352 B.n260 VSUBS 0.009259f
C353 B.n261 VSUBS 0.009259f
C354 B.n262 VSUBS 0.009259f
C355 B.n263 VSUBS 0.009259f
C356 B.n264 VSUBS 0.009259f
C357 B.n265 VSUBS 0.009259f
C358 B.n266 VSUBS 0.009259f
C359 B.n267 VSUBS 0.009259f
C360 B.n268 VSUBS 0.009259f
C361 B.n269 VSUBS 0.009259f
C362 B.n270 VSUBS 0.009259f
C363 B.n271 VSUBS 0.009259f
C364 B.n272 VSUBS 0.009259f
C365 B.n273 VSUBS 0.009259f
C366 B.n274 VSUBS 0.009259f
C367 B.n275 VSUBS 0.009259f
C368 B.n276 VSUBS 0.009259f
C369 B.n277 VSUBS 0.009259f
C370 B.n278 VSUBS 0.009259f
C371 B.n279 VSUBS 0.009259f
C372 B.n280 VSUBS 0.009259f
C373 B.n281 VSUBS 0.009259f
C374 B.n282 VSUBS 0.009259f
C375 B.n283 VSUBS 0.009259f
C376 B.n284 VSUBS 0.009259f
C377 B.n285 VSUBS 0.009259f
C378 B.n286 VSUBS 0.009259f
C379 B.n287 VSUBS 0.009259f
C380 B.n288 VSUBS 0.009259f
C381 B.n289 VSUBS 0.009259f
C382 B.n290 VSUBS 0.009259f
C383 B.n291 VSUBS 0.009259f
C384 B.n292 VSUBS 0.009259f
C385 B.n293 VSUBS 0.009259f
C386 B.n294 VSUBS 0.009259f
C387 B.n295 VSUBS 0.009259f
C388 B.n296 VSUBS 0.009259f
C389 B.n297 VSUBS 0.009259f
C390 B.n298 VSUBS 0.009259f
C391 B.n299 VSUBS 0.009259f
C392 B.n300 VSUBS 0.009259f
C393 B.n301 VSUBS 0.009259f
C394 B.n302 VSUBS 0.009259f
C395 B.n303 VSUBS 0.009259f
C396 B.n304 VSUBS 0.009259f
C397 B.n305 VSUBS 0.009259f
C398 B.n306 VSUBS 0.009259f
C399 B.n307 VSUBS 0.009259f
C400 B.n308 VSUBS 0.009259f
C401 B.n309 VSUBS 0.009259f
C402 B.n310 VSUBS 0.009259f
C403 B.n311 VSUBS 0.009259f
C404 B.n312 VSUBS 0.009259f
C405 B.n313 VSUBS 0.009259f
C406 B.n314 VSUBS 0.009259f
C407 B.n315 VSUBS 0.009259f
C408 B.n316 VSUBS 0.009259f
C409 B.n317 VSUBS 0.009259f
C410 B.n318 VSUBS 0.009259f
C411 B.n319 VSUBS 0.009259f
C412 B.n320 VSUBS 0.009259f
C413 B.n321 VSUBS 0.009259f
C414 B.n322 VSUBS 0.009259f
C415 B.n323 VSUBS 0.009259f
C416 B.n324 VSUBS 0.009259f
C417 B.n325 VSUBS 0.009259f
C418 B.n326 VSUBS 0.009259f
C419 B.n327 VSUBS 0.009259f
C420 B.n328 VSUBS 0.009259f
C421 B.n329 VSUBS 0.009259f
C422 B.n330 VSUBS 0.009259f
C423 B.n331 VSUBS 0.009259f
C424 B.n332 VSUBS 0.009259f
C425 B.n333 VSUBS 0.022608f
C426 B.n334 VSUBS 0.022608f
C427 B.n335 VSUBS 0.023413f
C428 B.n336 VSUBS 0.009259f
C429 B.n337 VSUBS 0.009259f
C430 B.n338 VSUBS 0.009259f
C431 B.n339 VSUBS 0.009259f
C432 B.n340 VSUBS 0.009259f
C433 B.n341 VSUBS 0.009259f
C434 B.n342 VSUBS 0.009259f
C435 B.n343 VSUBS 0.009259f
C436 B.n344 VSUBS 0.009259f
C437 B.n345 VSUBS 0.009259f
C438 B.n346 VSUBS 0.009259f
C439 B.n347 VSUBS 0.009259f
C440 B.n348 VSUBS 0.009259f
C441 B.n349 VSUBS 0.009259f
C442 B.n350 VSUBS 0.009259f
C443 B.n351 VSUBS 0.009259f
C444 B.n352 VSUBS 0.009259f
C445 B.n353 VSUBS 0.009259f
C446 B.n354 VSUBS 0.009259f
C447 B.n355 VSUBS 0.009259f
C448 B.n356 VSUBS 0.009259f
C449 B.n357 VSUBS 0.009259f
C450 B.n358 VSUBS 0.009259f
C451 B.n359 VSUBS 0.009259f
C452 B.n360 VSUBS 0.009259f
C453 B.n361 VSUBS 0.009259f
C454 B.n362 VSUBS 0.009259f
C455 B.n363 VSUBS 0.008714f
C456 B.n364 VSUBS 0.009259f
C457 B.n365 VSUBS 0.009259f
C458 B.n366 VSUBS 0.005174f
C459 B.n367 VSUBS 0.009259f
C460 B.n368 VSUBS 0.009259f
C461 B.n369 VSUBS 0.009259f
C462 B.n370 VSUBS 0.009259f
C463 B.n371 VSUBS 0.009259f
C464 B.n372 VSUBS 0.009259f
C465 B.n373 VSUBS 0.009259f
C466 B.n374 VSUBS 0.009259f
C467 B.n375 VSUBS 0.009259f
C468 B.n376 VSUBS 0.009259f
C469 B.n377 VSUBS 0.009259f
C470 B.n378 VSUBS 0.009259f
C471 B.n379 VSUBS 0.005174f
C472 B.n380 VSUBS 0.021451f
C473 B.n381 VSUBS 0.008714f
C474 B.n382 VSUBS 0.009259f
C475 B.n383 VSUBS 0.009259f
C476 B.n384 VSUBS 0.009259f
C477 B.n385 VSUBS 0.009259f
C478 B.n386 VSUBS 0.009259f
C479 B.n387 VSUBS 0.009259f
C480 B.n388 VSUBS 0.009259f
C481 B.n389 VSUBS 0.009259f
C482 B.n390 VSUBS 0.009259f
C483 B.n391 VSUBS 0.009259f
C484 B.n392 VSUBS 0.009259f
C485 B.n393 VSUBS 0.009259f
C486 B.n394 VSUBS 0.009259f
C487 B.n395 VSUBS 0.009259f
C488 B.n396 VSUBS 0.009259f
C489 B.n397 VSUBS 0.009259f
C490 B.n398 VSUBS 0.009259f
C491 B.n399 VSUBS 0.009259f
C492 B.n400 VSUBS 0.009259f
C493 B.n401 VSUBS 0.009259f
C494 B.n402 VSUBS 0.009259f
C495 B.n403 VSUBS 0.009259f
C496 B.n404 VSUBS 0.009259f
C497 B.n405 VSUBS 0.009259f
C498 B.n406 VSUBS 0.009259f
C499 B.n407 VSUBS 0.009259f
C500 B.n408 VSUBS 0.009259f
C501 B.n409 VSUBS 0.009259f
C502 B.n410 VSUBS 0.023413f
C503 B.n411 VSUBS 0.022608f
C504 B.n412 VSUBS 0.022608f
C505 B.n413 VSUBS 0.009259f
C506 B.n414 VSUBS 0.009259f
C507 B.n415 VSUBS 0.009259f
C508 B.n416 VSUBS 0.009259f
C509 B.n417 VSUBS 0.009259f
C510 B.n418 VSUBS 0.009259f
C511 B.n419 VSUBS 0.009259f
C512 B.n420 VSUBS 0.009259f
C513 B.n421 VSUBS 0.009259f
C514 B.n422 VSUBS 0.009259f
C515 B.n423 VSUBS 0.009259f
C516 B.n424 VSUBS 0.009259f
C517 B.n425 VSUBS 0.009259f
C518 B.n426 VSUBS 0.009259f
C519 B.n427 VSUBS 0.009259f
C520 B.n428 VSUBS 0.009259f
C521 B.n429 VSUBS 0.009259f
C522 B.n430 VSUBS 0.009259f
C523 B.n431 VSUBS 0.009259f
C524 B.n432 VSUBS 0.009259f
C525 B.n433 VSUBS 0.009259f
C526 B.n434 VSUBS 0.009259f
C527 B.n435 VSUBS 0.009259f
C528 B.n436 VSUBS 0.009259f
C529 B.n437 VSUBS 0.009259f
C530 B.n438 VSUBS 0.009259f
C531 B.n439 VSUBS 0.009259f
C532 B.n440 VSUBS 0.009259f
C533 B.n441 VSUBS 0.009259f
C534 B.n442 VSUBS 0.009259f
C535 B.n443 VSUBS 0.009259f
C536 B.n444 VSUBS 0.009259f
C537 B.n445 VSUBS 0.009259f
C538 B.n446 VSUBS 0.009259f
C539 B.n447 VSUBS 0.009259f
C540 B.n448 VSUBS 0.009259f
C541 B.n449 VSUBS 0.009259f
C542 B.n450 VSUBS 0.009259f
C543 B.n451 VSUBS 0.009259f
C544 B.n452 VSUBS 0.009259f
C545 B.n453 VSUBS 0.009259f
C546 B.n454 VSUBS 0.009259f
C547 B.n455 VSUBS 0.012082f
C548 B.n456 VSUBS 0.01287f
C549 B.n457 VSUBS 0.025594f
C550 VTAIL.t4 VSUBS 0.108376f
C551 VTAIL.t3 VSUBS 0.108376f
C552 VTAIL.n0 VSUBS 0.612721f
C553 VTAIL.n1 VSUBS 0.579484f
C554 VTAIL.t2 VSUBS 0.850595f
C555 VTAIL.n2 VSUBS 0.675158f
C556 VTAIL.t11 VSUBS 0.850595f
C557 VTAIL.n3 VSUBS 0.675158f
C558 VTAIL.t13 VSUBS 0.108376f
C559 VTAIL.t12 VSUBS 0.108376f
C560 VTAIL.n4 VSUBS 0.612721f
C561 VTAIL.n5 VSUBS 0.695799f
C562 VTAIL.t10 VSUBS 0.850595f
C563 VTAIL.n6 VSUBS 1.52338f
C564 VTAIL.t0 VSUBS 0.850598f
C565 VTAIL.n7 VSUBS 1.52338f
C566 VTAIL.t1 VSUBS 0.108376f
C567 VTAIL.t7 VSUBS 0.108376f
C568 VTAIL.n8 VSUBS 0.612724f
C569 VTAIL.n9 VSUBS 0.695797f
C570 VTAIL.t5 VSUBS 0.850598f
C571 VTAIL.n10 VSUBS 0.675154f
C572 VTAIL.t9 VSUBS 0.850598f
C573 VTAIL.n11 VSUBS 0.675154f
C574 VTAIL.t8 VSUBS 0.108376f
C575 VTAIL.t15 VSUBS 0.108376f
C576 VTAIL.n12 VSUBS 0.612724f
C577 VTAIL.n13 VSUBS 0.695797f
C578 VTAIL.t14 VSUBS 0.850592f
C579 VTAIL.n14 VSUBS 1.52338f
C580 VTAIL.t6 VSUBS 0.850595f
C581 VTAIL.n15 VSUBS 1.51801f
C582 VDD1.t0 VSUBS 0.096995f
C583 VDD1.t7 VSUBS 0.096995f
C584 VDD1.n0 VSUBS 0.621895f
C585 VDD1.t5 VSUBS 0.096995f
C586 VDD1.t1 VSUBS 0.096995f
C587 VDD1.n1 VSUBS 0.621254f
C588 VDD1.t3 VSUBS 0.096995f
C589 VDD1.t4 VSUBS 0.096995f
C590 VDD1.n2 VSUBS 0.621254f
C591 VDD1.n3 VSUBS 2.45488f
C592 VDD1.t6 VSUBS 0.096995f
C593 VDD1.t2 VSUBS 0.096995f
C594 VDD1.n4 VSUBS 0.618132f
C595 VDD1.n5 VSUBS 2.13301f
C596 VP.n0 VSUBS 0.0734f
C597 VP.t3 VSUBS 0.824422f
C598 VP.n1 VSUBS 0.34597f
C599 VP.n2 VSUBS 0.055007f
C600 VP.t2 VSUBS 0.824422f
C601 VP.n3 VSUBS 0.34597f
C602 VP.n4 VSUBS 0.0734f
C603 VP.n5 VSUBS 0.0734f
C604 VP.t1 VSUBS 0.925548f
C605 VP.t0 VSUBS 0.824422f
C606 VP.n6 VSUBS 0.34597f
C607 VP.n7 VSUBS 0.055007f
C608 VP.t7 VSUBS 0.824422f
C609 VP.n8 VSUBS 0.41572f
C610 VP.t6 VSUBS 0.983084f
C611 VP.n9 VSUBS 0.437619f
C612 VP.n10 VSUBS 0.282372f
C613 VP.n11 VSUBS 0.085534f
C614 VP.n12 VSUBS 0.044468f
C615 VP.n13 VSUBS 0.085534f
C616 VP.n14 VSUBS 0.055007f
C617 VP.n15 VSUBS 0.055007f
C618 VP.n16 VSUBS 0.083811f
C619 VP.n17 VSUBS 0.032218f
C620 VP.n18 VSUBS 0.446378f
C621 VP.n19 VSUBS 2.01912f
C622 VP.n20 VSUBS 2.06983f
C623 VP.t5 VSUBS 0.925548f
C624 VP.n21 VSUBS 0.446378f
C625 VP.n22 VSUBS 0.032218f
C626 VP.n23 VSUBS 0.083811f
C627 VP.n24 VSUBS 0.055007f
C628 VP.n25 VSUBS 0.055007f
C629 VP.n26 VSUBS 0.085534f
C630 VP.n27 VSUBS 0.044468f
C631 VP.n28 VSUBS 0.085534f
C632 VP.n29 VSUBS 0.055007f
C633 VP.n30 VSUBS 0.055007f
C634 VP.n31 VSUBS 0.083811f
C635 VP.n32 VSUBS 0.032218f
C636 VP.t4 VSUBS 0.925548f
C637 VP.n33 VSUBS 0.446378f
C638 VP.n34 VSUBS 0.051516f
.ends

