* NGSPICE file created from diff_pair_sample_1425.ext - technology: sky130A

.subckt diff_pair_sample_1425 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=0.60885 pd=4.02 as=0.60885 ps=4.02 w=3.69 l=2.14
X1 VTAIL.t7 VN.t0 VDD2.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.60885 pd=4.02 as=0.60885 ps=4.02 w=3.69 l=2.14
X2 VTAIL.t6 VN.t1 VDD2.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.4391 pd=8.16 as=0.60885 ps=4.02 w=3.69 l=2.14
X3 VDD2.t5 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.60885 pd=4.02 as=1.4391 ps=8.16 w=3.69 l=2.14
X4 VTAIL.t14 VP.t1 VDD1.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.4391 pd=8.16 as=0.60885 ps=4.02 w=3.69 l=2.14
X5 VTAIL.t13 VP.t2 VDD1.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=1.4391 pd=8.16 as=0.60885 ps=4.02 w=3.69 l=2.14
X6 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=1.4391 pd=8.16 as=0 ps=0 w=3.69 l=2.14
X7 VDD1.t4 VP.t3 VTAIL.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=0.60885 pd=4.02 as=1.4391 ps=8.16 w=3.69 l=2.14
X8 VDD2.t4 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.60885 pd=4.02 as=0.60885 ps=4.02 w=3.69 l=2.14
X9 VTAIL.t11 VP.t4 VDD1.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=0.60885 pd=4.02 as=0.60885 ps=4.02 w=3.69 l=2.14
X10 VDD1.t7 VP.t5 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=0.60885 pd=4.02 as=0.60885 ps=4.02 w=3.69 l=2.14
X11 VDD2.t3 VN.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.60885 pd=4.02 as=0.60885 ps=4.02 w=3.69 l=2.14
X12 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=1.4391 pd=8.16 as=0 ps=0 w=3.69 l=2.14
X13 VDD2.t2 VN.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.60885 pd=4.02 as=1.4391 ps=8.16 w=3.69 l=2.14
X14 VDD1.t2 VP.t6 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=0.60885 pd=4.02 as=0.60885 ps=4.02 w=3.69 l=2.14
X15 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=1.4391 pd=8.16 as=0 ps=0 w=3.69 l=2.14
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.4391 pd=8.16 as=0 ps=0 w=3.69 l=2.14
X17 VTAIL.t3 VN.t6 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=0.60885 pd=4.02 as=0.60885 ps=4.02 w=3.69 l=2.14
X18 VDD1.t5 VP.t7 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=0.60885 pd=4.02 as=1.4391 ps=8.16 w=3.69 l=2.14
X19 VTAIL.t2 VN.t7 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.4391 pd=8.16 as=0.60885 ps=4.02 w=3.69 l=2.14
R0 VP.n15 VP.n12 161.3
R1 VP.n17 VP.n16 161.3
R2 VP.n18 VP.n11 161.3
R3 VP.n20 VP.n19 161.3
R4 VP.n22 VP.n10 161.3
R5 VP.n24 VP.n23 161.3
R6 VP.n25 VP.n9 161.3
R7 VP.n27 VP.n26 161.3
R8 VP.n28 VP.n8 161.3
R9 VP.n54 VP.n0 161.3
R10 VP.n53 VP.n52 161.3
R11 VP.n51 VP.n1 161.3
R12 VP.n50 VP.n49 161.3
R13 VP.n48 VP.n2 161.3
R14 VP.n46 VP.n45 161.3
R15 VP.n44 VP.n3 161.3
R16 VP.n43 VP.n42 161.3
R17 VP.n41 VP.n4 161.3
R18 VP.n39 VP.n38 161.3
R19 VP.n37 VP.n5 161.3
R20 VP.n36 VP.n35 161.3
R21 VP.n34 VP.n6 161.3
R22 VP.n33 VP.n32 161.3
R23 VP.n31 VP.n7 88.4915
R24 VP.n56 VP.n55 88.4915
R25 VP.n30 VP.n29 88.4915
R26 VP.n13 VP.t1 76.0516
R27 VP.n35 VP.n34 56.5193
R28 VP.n42 VP.n3 56.5193
R29 VP.n53 VP.n1 56.5193
R30 VP.n27 VP.n9 56.5193
R31 VP.n16 VP.n11 56.5193
R32 VP.n14 VP.n13 47.0153
R33 VP.n31 VP.n30 42.545
R34 VP.n7 VP.t2 41.5561
R35 VP.n40 VP.t6 41.5561
R36 VP.n47 VP.t4 41.5561
R37 VP.n55 VP.t7 41.5561
R38 VP.n29 VP.t3 41.5561
R39 VP.n21 VP.t0 41.5561
R40 VP.n14 VP.t5 41.5561
R41 VP.n34 VP.n33 24.4675
R42 VP.n35 VP.n5 24.4675
R43 VP.n39 VP.n5 24.4675
R44 VP.n42 VP.n41 24.4675
R45 VP.n46 VP.n3 24.4675
R46 VP.n49 VP.n48 24.4675
R47 VP.n49 VP.n1 24.4675
R48 VP.n54 VP.n53 24.4675
R49 VP.n28 VP.n27 24.4675
R50 VP.n20 VP.n11 24.4675
R51 VP.n23 VP.n22 24.4675
R52 VP.n23 VP.n9 24.4675
R53 VP.n16 VP.n15 24.4675
R54 VP.n41 VP.n40 23.7335
R55 VP.n47 VP.n46 23.7335
R56 VP.n21 VP.n20 23.7335
R57 VP.n15 VP.n14 23.7335
R58 VP.n33 VP.n7 22.2655
R59 VP.n55 VP.n54 22.2655
R60 VP.n29 VP.n28 22.2655
R61 VP.n13 VP.n12 8.75906
R62 VP.n40 VP.n39 0.73451
R63 VP.n48 VP.n47 0.73451
R64 VP.n22 VP.n21 0.73451
R65 VP.n30 VP.n8 0.278367
R66 VP.n32 VP.n31 0.278367
R67 VP.n56 VP.n0 0.278367
R68 VP.n17 VP.n12 0.189894
R69 VP.n18 VP.n17 0.189894
R70 VP.n19 VP.n18 0.189894
R71 VP.n19 VP.n10 0.189894
R72 VP.n24 VP.n10 0.189894
R73 VP.n25 VP.n24 0.189894
R74 VP.n26 VP.n25 0.189894
R75 VP.n26 VP.n8 0.189894
R76 VP.n32 VP.n6 0.189894
R77 VP.n36 VP.n6 0.189894
R78 VP.n37 VP.n36 0.189894
R79 VP.n38 VP.n37 0.189894
R80 VP.n38 VP.n4 0.189894
R81 VP.n43 VP.n4 0.189894
R82 VP.n44 VP.n43 0.189894
R83 VP.n45 VP.n44 0.189894
R84 VP.n45 VP.n2 0.189894
R85 VP.n50 VP.n2 0.189894
R86 VP.n51 VP.n50 0.189894
R87 VP.n52 VP.n51 0.189894
R88 VP.n52 VP.n0 0.189894
R89 VP VP.n56 0.153454
R90 VDD1 VDD1.n0 80.5562
R91 VDD1.n3 VDD1.n2 80.4425
R92 VDD1.n3 VDD1.n1 80.4425
R93 VDD1.n5 VDD1.n4 79.4332
R94 VDD1.n5 VDD1.n3 37.0612
R95 VDD1.n4 VDD1.t1 5.36635
R96 VDD1.n4 VDD1.t4 5.36635
R97 VDD1.n0 VDD1.t6 5.36635
R98 VDD1.n0 VDD1.t7 5.36635
R99 VDD1.n2 VDD1.t0 5.36635
R100 VDD1.n2 VDD1.t5 5.36635
R101 VDD1.n1 VDD1.t3 5.36635
R102 VDD1.n1 VDD1.t2 5.36635
R103 VDD1 VDD1.n5 1.00697
R104 VTAIL.n11 VTAIL.t14 68.1203
R105 VTAIL.n10 VTAIL.t4 68.1203
R106 VTAIL.n7 VTAIL.t6 68.1203
R107 VTAIL.n15 VTAIL.t1 68.1203
R108 VTAIL.n2 VTAIL.t2 68.1203
R109 VTAIL.n3 VTAIL.t8 68.1203
R110 VTAIL.n6 VTAIL.t13 68.1203
R111 VTAIL.n14 VTAIL.t12 68.1203
R112 VTAIL.n13 VTAIL.n12 62.7546
R113 VTAIL.n9 VTAIL.n8 62.7546
R114 VTAIL.n1 VTAIL.n0 62.7544
R115 VTAIL.n5 VTAIL.n4 62.7544
R116 VTAIL.n15 VTAIL.n14 17.6772
R117 VTAIL.n7 VTAIL.n6 17.6772
R118 VTAIL.n0 VTAIL.t0 5.36635
R119 VTAIL.n0 VTAIL.t3 5.36635
R120 VTAIL.n4 VTAIL.t9 5.36635
R121 VTAIL.n4 VTAIL.t11 5.36635
R122 VTAIL.n12 VTAIL.t10 5.36635
R123 VTAIL.n12 VTAIL.t15 5.36635
R124 VTAIL.n8 VTAIL.t5 5.36635
R125 VTAIL.n8 VTAIL.t7 5.36635
R126 VTAIL.n9 VTAIL.n7 2.12981
R127 VTAIL.n10 VTAIL.n9 2.12981
R128 VTAIL.n13 VTAIL.n11 2.12981
R129 VTAIL.n14 VTAIL.n13 2.12981
R130 VTAIL.n6 VTAIL.n5 2.12981
R131 VTAIL.n5 VTAIL.n3 2.12981
R132 VTAIL.n2 VTAIL.n1 2.12981
R133 VTAIL VTAIL.n15 2.07162
R134 VTAIL.n11 VTAIL.n10 0.470328
R135 VTAIL.n3 VTAIL.n2 0.470328
R136 VTAIL VTAIL.n1 0.0586897
R137 B.n585 B.n584 585
R138 B.n194 B.n105 585
R139 B.n193 B.n192 585
R140 B.n191 B.n190 585
R141 B.n189 B.n188 585
R142 B.n187 B.n186 585
R143 B.n185 B.n184 585
R144 B.n183 B.n182 585
R145 B.n181 B.n180 585
R146 B.n179 B.n178 585
R147 B.n177 B.n176 585
R148 B.n175 B.n174 585
R149 B.n173 B.n172 585
R150 B.n171 B.n170 585
R151 B.n169 B.n168 585
R152 B.n167 B.n166 585
R153 B.n165 B.n164 585
R154 B.n162 B.n161 585
R155 B.n160 B.n159 585
R156 B.n158 B.n157 585
R157 B.n156 B.n155 585
R158 B.n154 B.n153 585
R159 B.n152 B.n151 585
R160 B.n150 B.n149 585
R161 B.n148 B.n147 585
R162 B.n146 B.n145 585
R163 B.n144 B.n143 585
R164 B.n141 B.n140 585
R165 B.n139 B.n138 585
R166 B.n137 B.n136 585
R167 B.n135 B.n134 585
R168 B.n133 B.n132 585
R169 B.n131 B.n130 585
R170 B.n129 B.n128 585
R171 B.n127 B.n126 585
R172 B.n125 B.n124 585
R173 B.n123 B.n122 585
R174 B.n121 B.n120 585
R175 B.n119 B.n118 585
R176 B.n117 B.n116 585
R177 B.n115 B.n114 585
R178 B.n113 B.n112 585
R179 B.n111 B.n110 585
R180 B.n82 B.n81 585
R181 B.n583 B.n83 585
R182 B.n588 B.n83 585
R183 B.n582 B.n581 585
R184 B.n581 B.n79 585
R185 B.n580 B.n78 585
R186 B.n594 B.n78 585
R187 B.n579 B.n77 585
R188 B.n595 B.n77 585
R189 B.n578 B.n76 585
R190 B.n596 B.n76 585
R191 B.n577 B.n576 585
R192 B.n576 B.n72 585
R193 B.n575 B.n71 585
R194 B.n602 B.n71 585
R195 B.n574 B.n70 585
R196 B.t16 B.n70 585
R197 B.n573 B.n69 585
R198 B.n603 B.n69 585
R199 B.n572 B.n571 585
R200 B.n571 B.n65 585
R201 B.n570 B.n64 585
R202 B.n609 B.n64 585
R203 B.n569 B.n63 585
R204 B.n610 B.n63 585
R205 B.n568 B.n62 585
R206 B.n611 B.n62 585
R207 B.n567 B.n566 585
R208 B.n566 B.n58 585
R209 B.n565 B.n57 585
R210 B.n617 B.n57 585
R211 B.n564 B.n56 585
R212 B.n618 B.n56 585
R213 B.n563 B.n55 585
R214 B.n619 B.n55 585
R215 B.n562 B.n561 585
R216 B.n561 B.n54 585
R217 B.n560 B.n50 585
R218 B.n625 B.n50 585
R219 B.n559 B.n49 585
R220 B.n626 B.n49 585
R221 B.n558 B.n48 585
R222 B.n627 B.n48 585
R223 B.n557 B.n556 585
R224 B.n556 B.n44 585
R225 B.n555 B.n43 585
R226 B.n633 B.n43 585
R227 B.n554 B.n42 585
R228 B.n634 B.n42 585
R229 B.n553 B.n41 585
R230 B.n635 B.n41 585
R231 B.n552 B.n551 585
R232 B.n551 B.n37 585
R233 B.n550 B.n36 585
R234 B.n641 B.n36 585
R235 B.n549 B.n35 585
R236 B.n642 B.n35 585
R237 B.n548 B.n34 585
R238 B.n643 B.n34 585
R239 B.n547 B.n546 585
R240 B.n546 B.n30 585
R241 B.n545 B.n29 585
R242 B.n649 B.n29 585
R243 B.n544 B.n28 585
R244 B.n650 B.n28 585
R245 B.n543 B.n27 585
R246 B.t0 B.n27 585
R247 B.n542 B.n541 585
R248 B.n541 B.n23 585
R249 B.n540 B.n22 585
R250 B.n656 B.n22 585
R251 B.n539 B.n21 585
R252 B.n657 B.n21 585
R253 B.n538 B.n20 585
R254 B.n658 B.n20 585
R255 B.n537 B.n536 585
R256 B.n536 B.n16 585
R257 B.n535 B.n15 585
R258 B.n664 B.n15 585
R259 B.n534 B.n14 585
R260 B.n665 B.n14 585
R261 B.n533 B.n13 585
R262 B.n666 B.n13 585
R263 B.n532 B.n531 585
R264 B.n531 B.n12 585
R265 B.n530 B.n529 585
R266 B.n530 B.n8 585
R267 B.n528 B.n7 585
R268 B.n673 B.n7 585
R269 B.n527 B.n6 585
R270 B.n674 B.n6 585
R271 B.n526 B.n5 585
R272 B.n675 B.n5 585
R273 B.n525 B.n524 585
R274 B.n524 B.n4 585
R275 B.n523 B.n195 585
R276 B.n523 B.n522 585
R277 B.n513 B.n196 585
R278 B.n197 B.n196 585
R279 B.n515 B.n514 585
R280 B.n516 B.n515 585
R281 B.n512 B.n201 585
R282 B.n205 B.n201 585
R283 B.n511 B.n510 585
R284 B.n510 B.n509 585
R285 B.n203 B.n202 585
R286 B.n204 B.n203 585
R287 B.n502 B.n501 585
R288 B.n503 B.n502 585
R289 B.n500 B.n210 585
R290 B.n210 B.n209 585
R291 B.n499 B.n498 585
R292 B.n498 B.n497 585
R293 B.n212 B.n211 585
R294 B.n213 B.n212 585
R295 B.n491 B.n490 585
R296 B.t7 B.n491 585
R297 B.n489 B.n218 585
R298 B.n218 B.n217 585
R299 B.n488 B.n487 585
R300 B.n487 B.n486 585
R301 B.n220 B.n219 585
R302 B.n221 B.n220 585
R303 B.n479 B.n478 585
R304 B.n480 B.n479 585
R305 B.n477 B.n226 585
R306 B.n226 B.n225 585
R307 B.n476 B.n475 585
R308 B.n475 B.n474 585
R309 B.n228 B.n227 585
R310 B.n229 B.n228 585
R311 B.n467 B.n466 585
R312 B.n468 B.n467 585
R313 B.n465 B.n234 585
R314 B.n234 B.n233 585
R315 B.n464 B.n463 585
R316 B.n463 B.n462 585
R317 B.n236 B.n235 585
R318 B.n237 B.n236 585
R319 B.n455 B.n454 585
R320 B.n456 B.n455 585
R321 B.n453 B.n242 585
R322 B.n242 B.n241 585
R323 B.n452 B.n451 585
R324 B.n451 B.n450 585
R325 B.n244 B.n243 585
R326 B.n443 B.n244 585
R327 B.n442 B.n441 585
R328 B.n444 B.n442 585
R329 B.n440 B.n249 585
R330 B.n249 B.n248 585
R331 B.n439 B.n438 585
R332 B.n438 B.n437 585
R333 B.n251 B.n250 585
R334 B.n252 B.n251 585
R335 B.n430 B.n429 585
R336 B.n431 B.n430 585
R337 B.n428 B.n257 585
R338 B.n257 B.n256 585
R339 B.n427 B.n426 585
R340 B.n426 B.n425 585
R341 B.n259 B.n258 585
R342 B.n260 B.n259 585
R343 B.n418 B.n417 585
R344 B.n419 B.n418 585
R345 B.n416 B.n264 585
R346 B.n264 B.t9 585
R347 B.n415 B.n414 585
R348 B.n414 B.n413 585
R349 B.n266 B.n265 585
R350 B.n267 B.n266 585
R351 B.n406 B.n405 585
R352 B.n407 B.n406 585
R353 B.n404 B.n272 585
R354 B.n272 B.n271 585
R355 B.n403 B.n402 585
R356 B.n402 B.n401 585
R357 B.n274 B.n273 585
R358 B.n275 B.n274 585
R359 B.n394 B.n393 585
R360 B.n395 B.n394 585
R361 B.n278 B.n277 585
R362 B.n309 B.n308 585
R363 B.n310 B.n306 585
R364 B.n306 B.n279 585
R365 B.n312 B.n311 585
R366 B.n314 B.n305 585
R367 B.n317 B.n316 585
R368 B.n318 B.n304 585
R369 B.n320 B.n319 585
R370 B.n322 B.n303 585
R371 B.n325 B.n324 585
R372 B.n326 B.n302 585
R373 B.n328 B.n327 585
R374 B.n330 B.n301 585
R375 B.n333 B.n332 585
R376 B.n334 B.n300 585
R377 B.n336 B.n335 585
R378 B.n338 B.n299 585
R379 B.n341 B.n340 585
R380 B.n342 B.n295 585
R381 B.n344 B.n343 585
R382 B.n346 B.n294 585
R383 B.n349 B.n348 585
R384 B.n350 B.n293 585
R385 B.n352 B.n351 585
R386 B.n354 B.n292 585
R387 B.n357 B.n356 585
R388 B.n358 B.n289 585
R389 B.n361 B.n360 585
R390 B.n363 B.n288 585
R391 B.n366 B.n365 585
R392 B.n367 B.n287 585
R393 B.n369 B.n368 585
R394 B.n371 B.n286 585
R395 B.n374 B.n373 585
R396 B.n375 B.n285 585
R397 B.n377 B.n376 585
R398 B.n379 B.n284 585
R399 B.n382 B.n381 585
R400 B.n383 B.n283 585
R401 B.n385 B.n384 585
R402 B.n387 B.n282 585
R403 B.n388 B.n281 585
R404 B.n391 B.n390 585
R405 B.n392 B.n280 585
R406 B.n280 B.n279 585
R407 B.n397 B.n396 585
R408 B.n396 B.n395 585
R409 B.n398 B.n276 585
R410 B.n276 B.n275 585
R411 B.n400 B.n399 585
R412 B.n401 B.n400 585
R413 B.n270 B.n269 585
R414 B.n271 B.n270 585
R415 B.n409 B.n408 585
R416 B.n408 B.n407 585
R417 B.n410 B.n268 585
R418 B.n268 B.n267 585
R419 B.n412 B.n411 585
R420 B.n413 B.n412 585
R421 B.n263 B.n262 585
R422 B.t9 B.n263 585
R423 B.n421 B.n420 585
R424 B.n420 B.n419 585
R425 B.n422 B.n261 585
R426 B.n261 B.n260 585
R427 B.n424 B.n423 585
R428 B.n425 B.n424 585
R429 B.n255 B.n254 585
R430 B.n256 B.n255 585
R431 B.n433 B.n432 585
R432 B.n432 B.n431 585
R433 B.n434 B.n253 585
R434 B.n253 B.n252 585
R435 B.n436 B.n435 585
R436 B.n437 B.n436 585
R437 B.n247 B.n246 585
R438 B.n248 B.n247 585
R439 B.n446 B.n445 585
R440 B.n445 B.n444 585
R441 B.n447 B.n245 585
R442 B.n443 B.n245 585
R443 B.n449 B.n448 585
R444 B.n450 B.n449 585
R445 B.n240 B.n239 585
R446 B.n241 B.n240 585
R447 B.n458 B.n457 585
R448 B.n457 B.n456 585
R449 B.n459 B.n238 585
R450 B.n238 B.n237 585
R451 B.n461 B.n460 585
R452 B.n462 B.n461 585
R453 B.n232 B.n231 585
R454 B.n233 B.n232 585
R455 B.n470 B.n469 585
R456 B.n469 B.n468 585
R457 B.n471 B.n230 585
R458 B.n230 B.n229 585
R459 B.n473 B.n472 585
R460 B.n474 B.n473 585
R461 B.n224 B.n223 585
R462 B.n225 B.n224 585
R463 B.n482 B.n481 585
R464 B.n481 B.n480 585
R465 B.n483 B.n222 585
R466 B.n222 B.n221 585
R467 B.n485 B.n484 585
R468 B.n486 B.n485 585
R469 B.n216 B.n215 585
R470 B.n217 B.n216 585
R471 B.n493 B.n492 585
R472 B.n492 B.t7 585
R473 B.n494 B.n214 585
R474 B.n214 B.n213 585
R475 B.n496 B.n495 585
R476 B.n497 B.n496 585
R477 B.n208 B.n207 585
R478 B.n209 B.n208 585
R479 B.n505 B.n504 585
R480 B.n504 B.n503 585
R481 B.n506 B.n206 585
R482 B.n206 B.n204 585
R483 B.n508 B.n507 585
R484 B.n509 B.n508 585
R485 B.n200 B.n199 585
R486 B.n205 B.n200 585
R487 B.n518 B.n517 585
R488 B.n517 B.n516 585
R489 B.n519 B.n198 585
R490 B.n198 B.n197 585
R491 B.n521 B.n520 585
R492 B.n522 B.n521 585
R493 B.n3 B.n0 585
R494 B.n4 B.n3 585
R495 B.n672 B.n1 585
R496 B.n673 B.n672 585
R497 B.n671 B.n670 585
R498 B.n671 B.n8 585
R499 B.n669 B.n9 585
R500 B.n12 B.n9 585
R501 B.n668 B.n667 585
R502 B.n667 B.n666 585
R503 B.n11 B.n10 585
R504 B.n665 B.n11 585
R505 B.n663 B.n662 585
R506 B.n664 B.n663 585
R507 B.n661 B.n17 585
R508 B.n17 B.n16 585
R509 B.n660 B.n659 585
R510 B.n659 B.n658 585
R511 B.n19 B.n18 585
R512 B.n657 B.n19 585
R513 B.n655 B.n654 585
R514 B.n656 B.n655 585
R515 B.n653 B.n24 585
R516 B.n24 B.n23 585
R517 B.n652 B.n651 585
R518 B.n651 B.t0 585
R519 B.n26 B.n25 585
R520 B.n650 B.n26 585
R521 B.n648 B.n647 585
R522 B.n649 B.n648 585
R523 B.n646 B.n31 585
R524 B.n31 B.n30 585
R525 B.n645 B.n644 585
R526 B.n644 B.n643 585
R527 B.n33 B.n32 585
R528 B.n642 B.n33 585
R529 B.n640 B.n639 585
R530 B.n641 B.n640 585
R531 B.n638 B.n38 585
R532 B.n38 B.n37 585
R533 B.n637 B.n636 585
R534 B.n636 B.n635 585
R535 B.n40 B.n39 585
R536 B.n634 B.n40 585
R537 B.n632 B.n631 585
R538 B.n633 B.n632 585
R539 B.n630 B.n45 585
R540 B.n45 B.n44 585
R541 B.n629 B.n628 585
R542 B.n628 B.n627 585
R543 B.n47 B.n46 585
R544 B.n626 B.n47 585
R545 B.n624 B.n623 585
R546 B.n625 B.n624 585
R547 B.n622 B.n51 585
R548 B.n54 B.n51 585
R549 B.n621 B.n620 585
R550 B.n620 B.n619 585
R551 B.n53 B.n52 585
R552 B.n618 B.n53 585
R553 B.n616 B.n615 585
R554 B.n617 B.n616 585
R555 B.n614 B.n59 585
R556 B.n59 B.n58 585
R557 B.n613 B.n612 585
R558 B.n612 B.n611 585
R559 B.n61 B.n60 585
R560 B.n610 B.n61 585
R561 B.n608 B.n607 585
R562 B.n609 B.n608 585
R563 B.n606 B.n66 585
R564 B.n66 B.n65 585
R565 B.n605 B.n604 585
R566 B.n604 B.n603 585
R567 B.n68 B.n67 585
R568 B.t16 B.n68 585
R569 B.n601 B.n600 585
R570 B.n602 B.n601 585
R571 B.n599 B.n73 585
R572 B.n73 B.n72 585
R573 B.n598 B.n597 585
R574 B.n597 B.n596 585
R575 B.n75 B.n74 585
R576 B.n595 B.n75 585
R577 B.n593 B.n592 585
R578 B.n594 B.n593 585
R579 B.n591 B.n80 585
R580 B.n80 B.n79 585
R581 B.n590 B.n589 585
R582 B.n589 B.n588 585
R583 B.n676 B.n675 585
R584 B.n674 B.n2 585
R585 B.n589 B.n82 482.89
R586 B.n585 B.n83 482.89
R587 B.n394 B.n280 482.89
R588 B.n396 B.n278 482.89
R589 B.n587 B.n586 256.663
R590 B.n587 B.n104 256.663
R591 B.n587 B.n103 256.663
R592 B.n587 B.n102 256.663
R593 B.n587 B.n101 256.663
R594 B.n587 B.n100 256.663
R595 B.n587 B.n99 256.663
R596 B.n587 B.n98 256.663
R597 B.n587 B.n97 256.663
R598 B.n587 B.n96 256.663
R599 B.n587 B.n95 256.663
R600 B.n587 B.n94 256.663
R601 B.n587 B.n93 256.663
R602 B.n587 B.n92 256.663
R603 B.n587 B.n91 256.663
R604 B.n587 B.n90 256.663
R605 B.n587 B.n89 256.663
R606 B.n587 B.n88 256.663
R607 B.n587 B.n87 256.663
R608 B.n587 B.n86 256.663
R609 B.n587 B.n85 256.663
R610 B.n587 B.n84 256.663
R611 B.n307 B.n279 256.663
R612 B.n313 B.n279 256.663
R613 B.n315 B.n279 256.663
R614 B.n321 B.n279 256.663
R615 B.n323 B.n279 256.663
R616 B.n329 B.n279 256.663
R617 B.n331 B.n279 256.663
R618 B.n337 B.n279 256.663
R619 B.n339 B.n279 256.663
R620 B.n345 B.n279 256.663
R621 B.n347 B.n279 256.663
R622 B.n353 B.n279 256.663
R623 B.n355 B.n279 256.663
R624 B.n362 B.n279 256.663
R625 B.n364 B.n279 256.663
R626 B.n370 B.n279 256.663
R627 B.n372 B.n279 256.663
R628 B.n378 B.n279 256.663
R629 B.n380 B.n279 256.663
R630 B.n386 B.n279 256.663
R631 B.n389 B.n279 256.663
R632 B.n678 B.n677 256.663
R633 B.n108 B.t19 248.785
R634 B.n106 B.t15 248.785
R635 B.n290 B.t12 248.785
R636 B.n296 B.t8 248.785
R637 B.n112 B.n111 163.367
R638 B.n116 B.n115 163.367
R639 B.n120 B.n119 163.367
R640 B.n124 B.n123 163.367
R641 B.n128 B.n127 163.367
R642 B.n132 B.n131 163.367
R643 B.n136 B.n135 163.367
R644 B.n140 B.n139 163.367
R645 B.n145 B.n144 163.367
R646 B.n149 B.n148 163.367
R647 B.n153 B.n152 163.367
R648 B.n157 B.n156 163.367
R649 B.n161 B.n160 163.367
R650 B.n166 B.n165 163.367
R651 B.n170 B.n169 163.367
R652 B.n174 B.n173 163.367
R653 B.n178 B.n177 163.367
R654 B.n182 B.n181 163.367
R655 B.n186 B.n185 163.367
R656 B.n190 B.n189 163.367
R657 B.n192 B.n105 163.367
R658 B.n394 B.n274 163.367
R659 B.n402 B.n274 163.367
R660 B.n402 B.n272 163.367
R661 B.n406 B.n272 163.367
R662 B.n406 B.n266 163.367
R663 B.n414 B.n266 163.367
R664 B.n414 B.n264 163.367
R665 B.n418 B.n264 163.367
R666 B.n418 B.n259 163.367
R667 B.n426 B.n259 163.367
R668 B.n426 B.n257 163.367
R669 B.n430 B.n257 163.367
R670 B.n430 B.n251 163.367
R671 B.n438 B.n251 163.367
R672 B.n438 B.n249 163.367
R673 B.n442 B.n249 163.367
R674 B.n442 B.n244 163.367
R675 B.n451 B.n244 163.367
R676 B.n451 B.n242 163.367
R677 B.n455 B.n242 163.367
R678 B.n455 B.n236 163.367
R679 B.n463 B.n236 163.367
R680 B.n463 B.n234 163.367
R681 B.n467 B.n234 163.367
R682 B.n467 B.n228 163.367
R683 B.n475 B.n228 163.367
R684 B.n475 B.n226 163.367
R685 B.n479 B.n226 163.367
R686 B.n479 B.n220 163.367
R687 B.n487 B.n220 163.367
R688 B.n487 B.n218 163.367
R689 B.n491 B.n218 163.367
R690 B.n491 B.n212 163.367
R691 B.n498 B.n212 163.367
R692 B.n498 B.n210 163.367
R693 B.n502 B.n210 163.367
R694 B.n502 B.n203 163.367
R695 B.n510 B.n203 163.367
R696 B.n510 B.n201 163.367
R697 B.n515 B.n201 163.367
R698 B.n515 B.n196 163.367
R699 B.n523 B.n196 163.367
R700 B.n524 B.n523 163.367
R701 B.n524 B.n5 163.367
R702 B.n6 B.n5 163.367
R703 B.n7 B.n6 163.367
R704 B.n530 B.n7 163.367
R705 B.n531 B.n530 163.367
R706 B.n531 B.n13 163.367
R707 B.n14 B.n13 163.367
R708 B.n15 B.n14 163.367
R709 B.n536 B.n15 163.367
R710 B.n536 B.n20 163.367
R711 B.n21 B.n20 163.367
R712 B.n22 B.n21 163.367
R713 B.n541 B.n22 163.367
R714 B.n541 B.n27 163.367
R715 B.n28 B.n27 163.367
R716 B.n29 B.n28 163.367
R717 B.n546 B.n29 163.367
R718 B.n546 B.n34 163.367
R719 B.n35 B.n34 163.367
R720 B.n36 B.n35 163.367
R721 B.n551 B.n36 163.367
R722 B.n551 B.n41 163.367
R723 B.n42 B.n41 163.367
R724 B.n43 B.n42 163.367
R725 B.n556 B.n43 163.367
R726 B.n556 B.n48 163.367
R727 B.n49 B.n48 163.367
R728 B.n50 B.n49 163.367
R729 B.n561 B.n50 163.367
R730 B.n561 B.n55 163.367
R731 B.n56 B.n55 163.367
R732 B.n57 B.n56 163.367
R733 B.n566 B.n57 163.367
R734 B.n566 B.n62 163.367
R735 B.n63 B.n62 163.367
R736 B.n64 B.n63 163.367
R737 B.n571 B.n64 163.367
R738 B.n571 B.n69 163.367
R739 B.n70 B.n69 163.367
R740 B.n71 B.n70 163.367
R741 B.n576 B.n71 163.367
R742 B.n576 B.n76 163.367
R743 B.n77 B.n76 163.367
R744 B.n78 B.n77 163.367
R745 B.n581 B.n78 163.367
R746 B.n581 B.n83 163.367
R747 B.n308 B.n306 163.367
R748 B.n312 B.n306 163.367
R749 B.n316 B.n314 163.367
R750 B.n320 B.n304 163.367
R751 B.n324 B.n322 163.367
R752 B.n328 B.n302 163.367
R753 B.n332 B.n330 163.367
R754 B.n336 B.n300 163.367
R755 B.n340 B.n338 163.367
R756 B.n344 B.n295 163.367
R757 B.n348 B.n346 163.367
R758 B.n352 B.n293 163.367
R759 B.n356 B.n354 163.367
R760 B.n361 B.n289 163.367
R761 B.n365 B.n363 163.367
R762 B.n369 B.n287 163.367
R763 B.n373 B.n371 163.367
R764 B.n377 B.n285 163.367
R765 B.n381 B.n379 163.367
R766 B.n385 B.n283 163.367
R767 B.n388 B.n387 163.367
R768 B.n390 B.n280 163.367
R769 B.n396 B.n276 163.367
R770 B.n400 B.n276 163.367
R771 B.n400 B.n270 163.367
R772 B.n408 B.n270 163.367
R773 B.n408 B.n268 163.367
R774 B.n412 B.n268 163.367
R775 B.n412 B.n263 163.367
R776 B.n420 B.n263 163.367
R777 B.n420 B.n261 163.367
R778 B.n424 B.n261 163.367
R779 B.n424 B.n255 163.367
R780 B.n432 B.n255 163.367
R781 B.n432 B.n253 163.367
R782 B.n436 B.n253 163.367
R783 B.n436 B.n247 163.367
R784 B.n445 B.n247 163.367
R785 B.n445 B.n245 163.367
R786 B.n449 B.n245 163.367
R787 B.n449 B.n240 163.367
R788 B.n457 B.n240 163.367
R789 B.n457 B.n238 163.367
R790 B.n461 B.n238 163.367
R791 B.n461 B.n232 163.367
R792 B.n469 B.n232 163.367
R793 B.n469 B.n230 163.367
R794 B.n473 B.n230 163.367
R795 B.n473 B.n224 163.367
R796 B.n481 B.n224 163.367
R797 B.n481 B.n222 163.367
R798 B.n485 B.n222 163.367
R799 B.n485 B.n216 163.367
R800 B.n492 B.n216 163.367
R801 B.n492 B.n214 163.367
R802 B.n496 B.n214 163.367
R803 B.n496 B.n208 163.367
R804 B.n504 B.n208 163.367
R805 B.n504 B.n206 163.367
R806 B.n508 B.n206 163.367
R807 B.n508 B.n200 163.367
R808 B.n517 B.n200 163.367
R809 B.n517 B.n198 163.367
R810 B.n521 B.n198 163.367
R811 B.n521 B.n3 163.367
R812 B.n676 B.n3 163.367
R813 B.n672 B.n2 163.367
R814 B.n672 B.n671 163.367
R815 B.n671 B.n9 163.367
R816 B.n667 B.n9 163.367
R817 B.n667 B.n11 163.367
R818 B.n663 B.n11 163.367
R819 B.n663 B.n17 163.367
R820 B.n659 B.n17 163.367
R821 B.n659 B.n19 163.367
R822 B.n655 B.n19 163.367
R823 B.n655 B.n24 163.367
R824 B.n651 B.n24 163.367
R825 B.n651 B.n26 163.367
R826 B.n648 B.n26 163.367
R827 B.n648 B.n31 163.367
R828 B.n644 B.n31 163.367
R829 B.n644 B.n33 163.367
R830 B.n640 B.n33 163.367
R831 B.n640 B.n38 163.367
R832 B.n636 B.n38 163.367
R833 B.n636 B.n40 163.367
R834 B.n632 B.n40 163.367
R835 B.n632 B.n45 163.367
R836 B.n628 B.n45 163.367
R837 B.n628 B.n47 163.367
R838 B.n624 B.n47 163.367
R839 B.n624 B.n51 163.367
R840 B.n620 B.n51 163.367
R841 B.n620 B.n53 163.367
R842 B.n616 B.n53 163.367
R843 B.n616 B.n59 163.367
R844 B.n612 B.n59 163.367
R845 B.n612 B.n61 163.367
R846 B.n608 B.n61 163.367
R847 B.n608 B.n66 163.367
R848 B.n604 B.n66 163.367
R849 B.n604 B.n68 163.367
R850 B.n601 B.n68 163.367
R851 B.n601 B.n73 163.367
R852 B.n597 B.n73 163.367
R853 B.n597 B.n75 163.367
R854 B.n593 B.n75 163.367
R855 B.n593 B.n80 163.367
R856 B.n589 B.n80 163.367
R857 B.n395 B.n279 146.012
R858 B.n588 B.n587 146.012
R859 B.n106 B.t17 125.855
R860 B.n290 B.t14 125.855
R861 B.n108 B.t20 125.852
R862 B.n296 B.t11 125.852
R863 B.n395 B.n275 83.4361
R864 B.n401 B.n275 83.4361
R865 B.n401 B.n271 83.4361
R866 B.n407 B.n271 83.4361
R867 B.n407 B.n267 83.4361
R868 B.n413 B.n267 83.4361
R869 B.n413 B.t9 83.4361
R870 B.n419 B.t9 83.4361
R871 B.n419 B.n260 83.4361
R872 B.n425 B.n260 83.4361
R873 B.n425 B.n256 83.4361
R874 B.n431 B.n256 83.4361
R875 B.n431 B.n252 83.4361
R876 B.n437 B.n252 83.4361
R877 B.n437 B.n248 83.4361
R878 B.n444 B.n248 83.4361
R879 B.n444 B.n443 83.4361
R880 B.n450 B.n241 83.4361
R881 B.n456 B.n241 83.4361
R882 B.n456 B.n237 83.4361
R883 B.n462 B.n237 83.4361
R884 B.n462 B.n233 83.4361
R885 B.n468 B.n233 83.4361
R886 B.n474 B.n229 83.4361
R887 B.n474 B.n225 83.4361
R888 B.n480 B.n225 83.4361
R889 B.n480 B.n221 83.4361
R890 B.n486 B.n221 83.4361
R891 B.n486 B.n217 83.4361
R892 B.t7 B.n217 83.4361
R893 B.t7 B.n213 83.4361
R894 B.n497 B.n213 83.4361
R895 B.n497 B.n209 83.4361
R896 B.n503 B.n209 83.4361
R897 B.n503 B.n204 83.4361
R898 B.n509 B.n204 83.4361
R899 B.n509 B.n205 83.4361
R900 B.n516 B.n197 83.4361
R901 B.n522 B.n197 83.4361
R902 B.n522 B.n4 83.4361
R903 B.n675 B.n4 83.4361
R904 B.n675 B.n674 83.4361
R905 B.n674 B.n673 83.4361
R906 B.n673 B.n8 83.4361
R907 B.n12 B.n8 83.4361
R908 B.n666 B.n12 83.4361
R909 B.n665 B.n664 83.4361
R910 B.n664 B.n16 83.4361
R911 B.n658 B.n16 83.4361
R912 B.n658 B.n657 83.4361
R913 B.n657 B.n656 83.4361
R914 B.n656 B.n23 83.4361
R915 B.t0 B.n23 83.4361
R916 B.t0 B.n650 83.4361
R917 B.n650 B.n649 83.4361
R918 B.n649 B.n30 83.4361
R919 B.n643 B.n30 83.4361
R920 B.n643 B.n642 83.4361
R921 B.n642 B.n641 83.4361
R922 B.n641 B.n37 83.4361
R923 B.n635 B.n634 83.4361
R924 B.n634 B.n633 83.4361
R925 B.n633 B.n44 83.4361
R926 B.n627 B.n44 83.4361
R927 B.n627 B.n626 83.4361
R928 B.n626 B.n625 83.4361
R929 B.n619 B.n54 83.4361
R930 B.n619 B.n618 83.4361
R931 B.n618 B.n617 83.4361
R932 B.n617 B.n58 83.4361
R933 B.n611 B.n58 83.4361
R934 B.n611 B.n610 83.4361
R935 B.n610 B.n609 83.4361
R936 B.n609 B.n65 83.4361
R937 B.n603 B.n65 83.4361
R938 B.n603 B.t16 83.4361
R939 B.t16 B.n602 83.4361
R940 B.n602 B.n72 83.4361
R941 B.n596 B.n72 83.4361
R942 B.n596 B.n595 83.4361
R943 B.n595 B.n594 83.4361
R944 B.n594 B.n79 83.4361
R945 B.n588 B.n79 83.4361
R946 B.n107 B.t18 77.9517
R947 B.n291 B.t13 77.9517
R948 B.n109 B.t21 77.9488
R949 B.n297 B.t10 77.9488
R950 B.n84 B.n82 71.676
R951 B.n112 B.n85 71.676
R952 B.n116 B.n86 71.676
R953 B.n120 B.n87 71.676
R954 B.n124 B.n88 71.676
R955 B.n128 B.n89 71.676
R956 B.n132 B.n90 71.676
R957 B.n136 B.n91 71.676
R958 B.n140 B.n92 71.676
R959 B.n145 B.n93 71.676
R960 B.n149 B.n94 71.676
R961 B.n153 B.n95 71.676
R962 B.n157 B.n96 71.676
R963 B.n161 B.n97 71.676
R964 B.n166 B.n98 71.676
R965 B.n170 B.n99 71.676
R966 B.n174 B.n100 71.676
R967 B.n178 B.n101 71.676
R968 B.n182 B.n102 71.676
R969 B.n186 B.n103 71.676
R970 B.n190 B.n104 71.676
R971 B.n586 B.n105 71.676
R972 B.n586 B.n585 71.676
R973 B.n192 B.n104 71.676
R974 B.n189 B.n103 71.676
R975 B.n185 B.n102 71.676
R976 B.n181 B.n101 71.676
R977 B.n177 B.n100 71.676
R978 B.n173 B.n99 71.676
R979 B.n169 B.n98 71.676
R980 B.n165 B.n97 71.676
R981 B.n160 B.n96 71.676
R982 B.n156 B.n95 71.676
R983 B.n152 B.n94 71.676
R984 B.n148 B.n93 71.676
R985 B.n144 B.n92 71.676
R986 B.n139 B.n91 71.676
R987 B.n135 B.n90 71.676
R988 B.n131 B.n89 71.676
R989 B.n127 B.n88 71.676
R990 B.n123 B.n87 71.676
R991 B.n119 B.n86 71.676
R992 B.n115 B.n85 71.676
R993 B.n111 B.n84 71.676
R994 B.n307 B.n278 71.676
R995 B.n313 B.n312 71.676
R996 B.n316 B.n315 71.676
R997 B.n321 B.n320 71.676
R998 B.n324 B.n323 71.676
R999 B.n329 B.n328 71.676
R1000 B.n332 B.n331 71.676
R1001 B.n337 B.n336 71.676
R1002 B.n340 B.n339 71.676
R1003 B.n345 B.n344 71.676
R1004 B.n348 B.n347 71.676
R1005 B.n353 B.n352 71.676
R1006 B.n356 B.n355 71.676
R1007 B.n362 B.n361 71.676
R1008 B.n365 B.n364 71.676
R1009 B.n370 B.n369 71.676
R1010 B.n373 B.n372 71.676
R1011 B.n378 B.n377 71.676
R1012 B.n381 B.n380 71.676
R1013 B.n386 B.n385 71.676
R1014 B.n389 B.n388 71.676
R1015 B.n308 B.n307 71.676
R1016 B.n314 B.n313 71.676
R1017 B.n315 B.n304 71.676
R1018 B.n322 B.n321 71.676
R1019 B.n323 B.n302 71.676
R1020 B.n330 B.n329 71.676
R1021 B.n331 B.n300 71.676
R1022 B.n338 B.n337 71.676
R1023 B.n339 B.n295 71.676
R1024 B.n346 B.n345 71.676
R1025 B.n347 B.n293 71.676
R1026 B.n354 B.n353 71.676
R1027 B.n355 B.n289 71.676
R1028 B.n363 B.n362 71.676
R1029 B.n364 B.n287 71.676
R1030 B.n371 B.n370 71.676
R1031 B.n372 B.n285 71.676
R1032 B.n379 B.n378 71.676
R1033 B.n380 B.n283 71.676
R1034 B.n387 B.n386 71.676
R1035 B.n390 B.n389 71.676
R1036 B.n677 B.n676 71.676
R1037 B.n677 B.n2 71.676
R1038 B.n468 B.t5 61.3502
R1039 B.n516 B.t4 61.3502
R1040 B.n666 B.t2 61.3502
R1041 B.n635 B.t3 61.3502
R1042 B.n142 B.n109 59.5399
R1043 B.n163 B.n107 59.5399
R1044 B.n359 B.n291 59.5399
R1045 B.n298 B.n297 59.5399
R1046 B.n109 B.n108 47.9035
R1047 B.n107 B.n106 47.9035
R1048 B.n291 B.n290 47.9035
R1049 B.n297 B.n296 47.9035
R1050 B.n450 B.t6 44.1723
R1051 B.n625 B.t1 44.1723
R1052 B.n443 B.t6 39.2643
R1053 B.n54 B.t1 39.2643
R1054 B.n397 B.n277 31.3761
R1055 B.n393 B.n392 31.3761
R1056 B.n584 B.n583 31.3761
R1057 B.n590 B.n81 31.3761
R1058 B.t5 B.n229 22.0864
R1059 B.n205 B.t4 22.0864
R1060 B.t2 B.n665 22.0864
R1061 B.t3 B.n37 22.0864
R1062 B B.n678 18.0485
R1063 B.n398 B.n397 10.6151
R1064 B.n399 B.n398 10.6151
R1065 B.n399 B.n269 10.6151
R1066 B.n409 B.n269 10.6151
R1067 B.n410 B.n409 10.6151
R1068 B.n411 B.n410 10.6151
R1069 B.n411 B.n262 10.6151
R1070 B.n421 B.n262 10.6151
R1071 B.n422 B.n421 10.6151
R1072 B.n423 B.n422 10.6151
R1073 B.n423 B.n254 10.6151
R1074 B.n433 B.n254 10.6151
R1075 B.n434 B.n433 10.6151
R1076 B.n435 B.n434 10.6151
R1077 B.n435 B.n246 10.6151
R1078 B.n446 B.n246 10.6151
R1079 B.n447 B.n446 10.6151
R1080 B.n448 B.n447 10.6151
R1081 B.n448 B.n239 10.6151
R1082 B.n458 B.n239 10.6151
R1083 B.n459 B.n458 10.6151
R1084 B.n460 B.n459 10.6151
R1085 B.n460 B.n231 10.6151
R1086 B.n470 B.n231 10.6151
R1087 B.n471 B.n470 10.6151
R1088 B.n472 B.n471 10.6151
R1089 B.n472 B.n223 10.6151
R1090 B.n482 B.n223 10.6151
R1091 B.n483 B.n482 10.6151
R1092 B.n484 B.n483 10.6151
R1093 B.n484 B.n215 10.6151
R1094 B.n493 B.n215 10.6151
R1095 B.n494 B.n493 10.6151
R1096 B.n495 B.n494 10.6151
R1097 B.n495 B.n207 10.6151
R1098 B.n505 B.n207 10.6151
R1099 B.n506 B.n505 10.6151
R1100 B.n507 B.n506 10.6151
R1101 B.n507 B.n199 10.6151
R1102 B.n518 B.n199 10.6151
R1103 B.n519 B.n518 10.6151
R1104 B.n520 B.n519 10.6151
R1105 B.n520 B.n0 10.6151
R1106 B.n309 B.n277 10.6151
R1107 B.n310 B.n309 10.6151
R1108 B.n311 B.n310 10.6151
R1109 B.n311 B.n305 10.6151
R1110 B.n317 B.n305 10.6151
R1111 B.n318 B.n317 10.6151
R1112 B.n319 B.n318 10.6151
R1113 B.n319 B.n303 10.6151
R1114 B.n325 B.n303 10.6151
R1115 B.n326 B.n325 10.6151
R1116 B.n327 B.n326 10.6151
R1117 B.n327 B.n301 10.6151
R1118 B.n333 B.n301 10.6151
R1119 B.n334 B.n333 10.6151
R1120 B.n335 B.n334 10.6151
R1121 B.n335 B.n299 10.6151
R1122 B.n342 B.n341 10.6151
R1123 B.n343 B.n342 10.6151
R1124 B.n343 B.n294 10.6151
R1125 B.n349 B.n294 10.6151
R1126 B.n350 B.n349 10.6151
R1127 B.n351 B.n350 10.6151
R1128 B.n351 B.n292 10.6151
R1129 B.n357 B.n292 10.6151
R1130 B.n358 B.n357 10.6151
R1131 B.n360 B.n288 10.6151
R1132 B.n366 B.n288 10.6151
R1133 B.n367 B.n366 10.6151
R1134 B.n368 B.n367 10.6151
R1135 B.n368 B.n286 10.6151
R1136 B.n374 B.n286 10.6151
R1137 B.n375 B.n374 10.6151
R1138 B.n376 B.n375 10.6151
R1139 B.n376 B.n284 10.6151
R1140 B.n382 B.n284 10.6151
R1141 B.n383 B.n382 10.6151
R1142 B.n384 B.n383 10.6151
R1143 B.n384 B.n282 10.6151
R1144 B.n282 B.n281 10.6151
R1145 B.n391 B.n281 10.6151
R1146 B.n392 B.n391 10.6151
R1147 B.n393 B.n273 10.6151
R1148 B.n403 B.n273 10.6151
R1149 B.n404 B.n403 10.6151
R1150 B.n405 B.n404 10.6151
R1151 B.n405 B.n265 10.6151
R1152 B.n415 B.n265 10.6151
R1153 B.n416 B.n415 10.6151
R1154 B.n417 B.n416 10.6151
R1155 B.n417 B.n258 10.6151
R1156 B.n427 B.n258 10.6151
R1157 B.n428 B.n427 10.6151
R1158 B.n429 B.n428 10.6151
R1159 B.n429 B.n250 10.6151
R1160 B.n439 B.n250 10.6151
R1161 B.n440 B.n439 10.6151
R1162 B.n441 B.n440 10.6151
R1163 B.n441 B.n243 10.6151
R1164 B.n452 B.n243 10.6151
R1165 B.n453 B.n452 10.6151
R1166 B.n454 B.n453 10.6151
R1167 B.n454 B.n235 10.6151
R1168 B.n464 B.n235 10.6151
R1169 B.n465 B.n464 10.6151
R1170 B.n466 B.n465 10.6151
R1171 B.n466 B.n227 10.6151
R1172 B.n476 B.n227 10.6151
R1173 B.n477 B.n476 10.6151
R1174 B.n478 B.n477 10.6151
R1175 B.n478 B.n219 10.6151
R1176 B.n488 B.n219 10.6151
R1177 B.n489 B.n488 10.6151
R1178 B.n490 B.n489 10.6151
R1179 B.n490 B.n211 10.6151
R1180 B.n499 B.n211 10.6151
R1181 B.n500 B.n499 10.6151
R1182 B.n501 B.n500 10.6151
R1183 B.n501 B.n202 10.6151
R1184 B.n511 B.n202 10.6151
R1185 B.n512 B.n511 10.6151
R1186 B.n514 B.n512 10.6151
R1187 B.n514 B.n513 10.6151
R1188 B.n513 B.n195 10.6151
R1189 B.n525 B.n195 10.6151
R1190 B.n526 B.n525 10.6151
R1191 B.n527 B.n526 10.6151
R1192 B.n528 B.n527 10.6151
R1193 B.n529 B.n528 10.6151
R1194 B.n532 B.n529 10.6151
R1195 B.n533 B.n532 10.6151
R1196 B.n534 B.n533 10.6151
R1197 B.n535 B.n534 10.6151
R1198 B.n537 B.n535 10.6151
R1199 B.n538 B.n537 10.6151
R1200 B.n539 B.n538 10.6151
R1201 B.n540 B.n539 10.6151
R1202 B.n542 B.n540 10.6151
R1203 B.n543 B.n542 10.6151
R1204 B.n544 B.n543 10.6151
R1205 B.n545 B.n544 10.6151
R1206 B.n547 B.n545 10.6151
R1207 B.n548 B.n547 10.6151
R1208 B.n549 B.n548 10.6151
R1209 B.n550 B.n549 10.6151
R1210 B.n552 B.n550 10.6151
R1211 B.n553 B.n552 10.6151
R1212 B.n554 B.n553 10.6151
R1213 B.n555 B.n554 10.6151
R1214 B.n557 B.n555 10.6151
R1215 B.n558 B.n557 10.6151
R1216 B.n559 B.n558 10.6151
R1217 B.n560 B.n559 10.6151
R1218 B.n562 B.n560 10.6151
R1219 B.n563 B.n562 10.6151
R1220 B.n564 B.n563 10.6151
R1221 B.n565 B.n564 10.6151
R1222 B.n567 B.n565 10.6151
R1223 B.n568 B.n567 10.6151
R1224 B.n569 B.n568 10.6151
R1225 B.n570 B.n569 10.6151
R1226 B.n572 B.n570 10.6151
R1227 B.n573 B.n572 10.6151
R1228 B.n574 B.n573 10.6151
R1229 B.n575 B.n574 10.6151
R1230 B.n577 B.n575 10.6151
R1231 B.n578 B.n577 10.6151
R1232 B.n579 B.n578 10.6151
R1233 B.n580 B.n579 10.6151
R1234 B.n582 B.n580 10.6151
R1235 B.n583 B.n582 10.6151
R1236 B.n670 B.n1 10.6151
R1237 B.n670 B.n669 10.6151
R1238 B.n669 B.n668 10.6151
R1239 B.n668 B.n10 10.6151
R1240 B.n662 B.n10 10.6151
R1241 B.n662 B.n661 10.6151
R1242 B.n661 B.n660 10.6151
R1243 B.n660 B.n18 10.6151
R1244 B.n654 B.n18 10.6151
R1245 B.n654 B.n653 10.6151
R1246 B.n653 B.n652 10.6151
R1247 B.n652 B.n25 10.6151
R1248 B.n647 B.n25 10.6151
R1249 B.n647 B.n646 10.6151
R1250 B.n646 B.n645 10.6151
R1251 B.n645 B.n32 10.6151
R1252 B.n639 B.n32 10.6151
R1253 B.n639 B.n638 10.6151
R1254 B.n638 B.n637 10.6151
R1255 B.n637 B.n39 10.6151
R1256 B.n631 B.n39 10.6151
R1257 B.n631 B.n630 10.6151
R1258 B.n630 B.n629 10.6151
R1259 B.n629 B.n46 10.6151
R1260 B.n623 B.n46 10.6151
R1261 B.n623 B.n622 10.6151
R1262 B.n622 B.n621 10.6151
R1263 B.n621 B.n52 10.6151
R1264 B.n615 B.n52 10.6151
R1265 B.n615 B.n614 10.6151
R1266 B.n614 B.n613 10.6151
R1267 B.n613 B.n60 10.6151
R1268 B.n607 B.n60 10.6151
R1269 B.n607 B.n606 10.6151
R1270 B.n606 B.n605 10.6151
R1271 B.n605 B.n67 10.6151
R1272 B.n600 B.n67 10.6151
R1273 B.n600 B.n599 10.6151
R1274 B.n599 B.n598 10.6151
R1275 B.n598 B.n74 10.6151
R1276 B.n592 B.n74 10.6151
R1277 B.n592 B.n591 10.6151
R1278 B.n591 B.n590 10.6151
R1279 B.n110 B.n81 10.6151
R1280 B.n113 B.n110 10.6151
R1281 B.n114 B.n113 10.6151
R1282 B.n117 B.n114 10.6151
R1283 B.n118 B.n117 10.6151
R1284 B.n121 B.n118 10.6151
R1285 B.n122 B.n121 10.6151
R1286 B.n125 B.n122 10.6151
R1287 B.n126 B.n125 10.6151
R1288 B.n129 B.n126 10.6151
R1289 B.n130 B.n129 10.6151
R1290 B.n133 B.n130 10.6151
R1291 B.n134 B.n133 10.6151
R1292 B.n137 B.n134 10.6151
R1293 B.n138 B.n137 10.6151
R1294 B.n141 B.n138 10.6151
R1295 B.n146 B.n143 10.6151
R1296 B.n147 B.n146 10.6151
R1297 B.n150 B.n147 10.6151
R1298 B.n151 B.n150 10.6151
R1299 B.n154 B.n151 10.6151
R1300 B.n155 B.n154 10.6151
R1301 B.n158 B.n155 10.6151
R1302 B.n159 B.n158 10.6151
R1303 B.n162 B.n159 10.6151
R1304 B.n167 B.n164 10.6151
R1305 B.n168 B.n167 10.6151
R1306 B.n171 B.n168 10.6151
R1307 B.n172 B.n171 10.6151
R1308 B.n175 B.n172 10.6151
R1309 B.n176 B.n175 10.6151
R1310 B.n179 B.n176 10.6151
R1311 B.n180 B.n179 10.6151
R1312 B.n183 B.n180 10.6151
R1313 B.n184 B.n183 10.6151
R1314 B.n187 B.n184 10.6151
R1315 B.n188 B.n187 10.6151
R1316 B.n191 B.n188 10.6151
R1317 B.n193 B.n191 10.6151
R1318 B.n194 B.n193 10.6151
R1319 B.n584 B.n194 10.6151
R1320 B.n299 B.n298 9.36635
R1321 B.n360 B.n359 9.36635
R1322 B.n142 B.n141 9.36635
R1323 B.n164 B.n163 9.36635
R1324 B.n678 B.n0 8.11757
R1325 B.n678 B.n1 8.11757
R1326 B.n341 B.n298 1.24928
R1327 B.n359 B.n358 1.24928
R1328 B.n143 B.n142 1.24928
R1329 B.n163 B.n162 1.24928
R1330 VN.n43 VN.n23 161.3
R1331 VN.n42 VN.n41 161.3
R1332 VN.n40 VN.n24 161.3
R1333 VN.n39 VN.n38 161.3
R1334 VN.n37 VN.n25 161.3
R1335 VN.n35 VN.n34 161.3
R1336 VN.n33 VN.n26 161.3
R1337 VN.n32 VN.n31 161.3
R1338 VN.n30 VN.n27 161.3
R1339 VN.n20 VN.n0 161.3
R1340 VN.n19 VN.n18 161.3
R1341 VN.n17 VN.n1 161.3
R1342 VN.n16 VN.n15 161.3
R1343 VN.n14 VN.n2 161.3
R1344 VN.n12 VN.n11 161.3
R1345 VN.n10 VN.n3 161.3
R1346 VN.n9 VN.n8 161.3
R1347 VN.n7 VN.n4 161.3
R1348 VN.n22 VN.n21 88.4915
R1349 VN.n45 VN.n44 88.4915
R1350 VN.n5 VN.t7 76.0516
R1351 VN.n28 VN.t5 76.0516
R1352 VN.n8 VN.n3 56.5193
R1353 VN.n19 VN.n1 56.5193
R1354 VN.n31 VN.n26 56.5193
R1355 VN.n42 VN.n24 56.5193
R1356 VN.n6 VN.n5 47.0153
R1357 VN.n29 VN.n28 47.0153
R1358 VN VN.n45 42.8239
R1359 VN.n6 VN.t3 41.5561
R1360 VN.n13 VN.t6 41.5561
R1361 VN.n21 VN.t2 41.5561
R1362 VN.n29 VN.t0 41.5561
R1363 VN.n36 VN.t4 41.5561
R1364 VN.n44 VN.t1 41.5561
R1365 VN.n8 VN.n7 24.4675
R1366 VN.n12 VN.n3 24.4675
R1367 VN.n15 VN.n14 24.4675
R1368 VN.n15 VN.n1 24.4675
R1369 VN.n20 VN.n19 24.4675
R1370 VN.n31 VN.n30 24.4675
R1371 VN.n38 VN.n24 24.4675
R1372 VN.n38 VN.n37 24.4675
R1373 VN.n35 VN.n26 24.4675
R1374 VN.n43 VN.n42 24.4675
R1375 VN.n7 VN.n6 23.7335
R1376 VN.n13 VN.n12 23.7335
R1377 VN.n30 VN.n29 23.7335
R1378 VN.n36 VN.n35 23.7335
R1379 VN.n21 VN.n20 22.2655
R1380 VN.n44 VN.n43 22.2655
R1381 VN.n28 VN.n27 8.75906
R1382 VN.n5 VN.n4 8.75906
R1383 VN.n14 VN.n13 0.73451
R1384 VN.n37 VN.n36 0.73451
R1385 VN.n45 VN.n23 0.278367
R1386 VN.n22 VN.n0 0.278367
R1387 VN.n41 VN.n23 0.189894
R1388 VN.n41 VN.n40 0.189894
R1389 VN.n40 VN.n39 0.189894
R1390 VN.n39 VN.n25 0.189894
R1391 VN.n34 VN.n25 0.189894
R1392 VN.n34 VN.n33 0.189894
R1393 VN.n33 VN.n32 0.189894
R1394 VN.n32 VN.n27 0.189894
R1395 VN.n9 VN.n4 0.189894
R1396 VN.n10 VN.n9 0.189894
R1397 VN.n11 VN.n10 0.189894
R1398 VN.n11 VN.n2 0.189894
R1399 VN.n16 VN.n2 0.189894
R1400 VN.n17 VN.n16 0.189894
R1401 VN.n18 VN.n17 0.189894
R1402 VN.n18 VN.n0 0.189894
R1403 VN VN.n22 0.153454
R1404 VDD2.n2 VDD2.n1 80.4425
R1405 VDD2.n2 VDD2.n0 80.4425
R1406 VDD2 VDD2.n5 80.4397
R1407 VDD2.n4 VDD2.n3 79.4334
R1408 VDD2.n4 VDD2.n2 36.4782
R1409 VDD2.n5 VDD2.t7 5.36635
R1410 VDD2.n5 VDD2.t2 5.36635
R1411 VDD2.n3 VDD2.t6 5.36635
R1412 VDD2.n3 VDD2.t3 5.36635
R1413 VDD2.n1 VDD2.t1 5.36635
R1414 VDD2.n1 VDD2.t5 5.36635
R1415 VDD2.n0 VDD2.t0 5.36635
R1416 VDD2.n0 VDD2.t4 5.36635
R1417 VDD2 VDD2.n4 1.12334
C0 VDD2 VN 2.86515f
C1 VP VN 5.56483f
C2 VDD2 VP 0.475902f
C3 VDD1 VN 0.155481f
C4 VDD2 VDD1 1.53864f
C5 VTAIL VN 3.65119f
C6 VDD2 VTAIL 5.0038f
C7 VDD1 VP 3.1837f
C8 VTAIL VP 3.66529f
C9 VDD1 VTAIL 4.95247f
C10 VDD2 B 4.244772f
C11 VDD1 B 4.642333f
C12 VTAIL B 4.88318f
C13 VN B 12.95325f
C14 VP B 11.513559f
C15 VDD2.t0 B 0.071177f
C16 VDD2.t4 B 0.071177f
C17 VDD2.n0 B 0.555495f
C18 VDD2.t1 B 0.071177f
C19 VDD2.t5 B 0.071177f
C20 VDD2.n1 B 0.555495f
C21 VDD2.n2 B 2.42688f
C22 VDD2.t6 B 0.071177f
C23 VDD2.t3 B 0.071177f
C24 VDD2.n3 B 0.549892f
C25 VDD2.n4 B 2.07952f
C26 VDD2.t7 B 0.071177f
C27 VDD2.t2 B 0.071177f
C28 VDD2.n5 B 0.555469f
C29 VN.n0 B 0.039523f
C30 VN.t2 B 0.603491f
C31 VN.n1 B 0.041257f
C32 VN.n2 B 0.029978f
C33 VN.t6 B 0.603491f
C34 VN.n3 B 0.043763f
C35 VN.n4 B 0.253045f
C36 VN.t3 B 0.603491f
C37 VN.t7 B 0.792034f
C38 VN.n5 B 0.309931f
C39 VN.n6 B 0.338801f
C40 VN.n7 B 0.055043f
C41 VN.n8 B 0.043763f
C42 VN.n9 B 0.029978f
C43 VN.n10 B 0.029978f
C44 VN.n11 B 0.029978f
C45 VN.n12 B 0.055043f
C46 VN.n13 B 0.248722f
C47 VN.n14 B 0.029114f
C48 VN.n15 B 0.055872f
C49 VN.n16 B 0.029978f
C50 VN.n17 B 0.029978f
C51 VN.n18 B 0.029978f
C52 VN.n19 B 0.046269f
C53 VN.n20 B 0.053388f
C54 VN.n21 B 0.351722f
C55 VN.n22 B 0.034625f
C56 VN.n23 B 0.039523f
C57 VN.t1 B 0.603491f
C58 VN.n24 B 0.041257f
C59 VN.n25 B 0.029978f
C60 VN.t4 B 0.603491f
C61 VN.n26 B 0.043763f
C62 VN.n27 B 0.253045f
C63 VN.t0 B 0.603491f
C64 VN.t5 B 0.792034f
C65 VN.n28 B 0.309931f
C66 VN.n29 B 0.338801f
C67 VN.n30 B 0.055043f
C68 VN.n31 B 0.043763f
C69 VN.n32 B 0.029978f
C70 VN.n33 B 0.029978f
C71 VN.n34 B 0.029978f
C72 VN.n35 B 0.055043f
C73 VN.n36 B 0.248722f
C74 VN.n37 B 0.029114f
C75 VN.n38 B 0.055872f
C76 VN.n39 B 0.029978f
C77 VN.n40 B 0.029978f
C78 VN.n41 B 0.029978f
C79 VN.n42 B 0.046269f
C80 VN.n43 B 0.053388f
C81 VN.n44 B 0.351722f
C82 VN.n45 B 1.30521f
C83 VTAIL.t0 B 0.07542f
C84 VTAIL.t3 B 0.07542f
C85 VTAIL.n0 B 0.53062f
C86 VTAIL.n1 B 0.39998f
C87 VTAIL.t2 B 0.68425f
C88 VTAIL.n2 B 0.486346f
C89 VTAIL.t8 B 0.68425f
C90 VTAIL.n3 B 0.486346f
C91 VTAIL.t9 B 0.07542f
C92 VTAIL.t11 B 0.07542f
C93 VTAIL.n4 B 0.53062f
C94 VTAIL.n5 B 0.572591f
C95 VTAIL.t13 B 0.68425f
C96 VTAIL.n6 B 1.2411f
C97 VTAIL.t6 B 0.684254f
C98 VTAIL.n7 B 1.2411f
C99 VTAIL.t5 B 0.07542f
C100 VTAIL.t7 B 0.07542f
C101 VTAIL.n8 B 0.530622f
C102 VTAIL.n9 B 0.572588f
C103 VTAIL.t4 B 0.684254f
C104 VTAIL.n10 B 0.486342f
C105 VTAIL.t14 B 0.684254f
C106 VTAIL.n11 B 0.486342f
C107 VTAIL.t10 B 0.07542f
C108 VTAIL.t15 B 0.07542f
C109 VTAIL.n12 B 0.530622f
C110 VTAIL.n13 B 0.572588f
C111 VTAIL.t12 B 0.68425f
C112 VTAIL.n14 B 1.2411f
C113 VTAIL.t1 B 0.68425f
C114 VTAIL.n15 B 1.23625f
C115 VDD1.t6 B 0.073046f
C116 VDD1.t7 B 0.073046f
C117 VDD1.n0 B 0.570843f
C118 VDD1.t3 B 0.073046f
C119 VDD1.t2 B 0.073046f
C120 VDD1.n1 B 0.570084f
C121 VDD1.t0 B 0.073046f
C122 VDD1.t5 B 0.073046f
C123 VDD1.n2 B 0.570084f
C124 VDD1.n3 B 2.54328f
C125 VDD1.t1 B 0.073046f
C126 VDD1.t4 B 0.073046f
C127 VDD1.n4 B 0.564331f
C128 VDD1.n5 B 2.16459f
C129 VP.n0 B 0.040636f
C130 VP.t7 B 0.620474f
C131 VP.n1 B 0.042418f
C132 VP.n2 B 0.030822f
C133 VP.t4 B 0.620474f
C134 VP.n3 B 0.044995f
C135 VP.n4 B 0.030822f
C136 VP.t6 B 0.620474f
C137 VP.n5 B 0.057444f
C138 VP.n6 B 0.030822f
C139 VP.t2 B 0.620474f
C140 VP.n7 B 0.36162f
C141 VP.n8 B 0.040636f
C142 VP.t3 B 0.620474f
C143 VP.n9 B 0.042418f
C144 VP.n10 B 0.030822f
C145 VP.t0 B 0.620474f
C146 VP.n11 B 0.044995f
C147 VP.n12 B 0.260166f
C148 VP.t5 B 0.620474f
C149 VP.t1 B 0.814323f
C150 VP.n13 B 0.318653f
C151 VP.n14 B 0.348335f
C152 VP.n15 B 0.056592f
C153 VP.n16 B 0.044995f
C154 VP.n17 B 0.030822f
C155 VP.n18 B 0.030822f
C156 VP.n19 B 0.030822f
C157 VP.n20 B 0.056592f
C158 VP.n21 B 0.255721f
C159 VP.n22 B 0.029933f
C160 VP.n23 B 0.057444f
C161 VP.n24 B 0.030822f
C162 VP.n25 B 0.030822f
C163 VP.n26 B 0.030822f
C164 VP.n27 B 0.047571f
C165 VP.n28 B 0.054891f
C166 VP.n29 B 0.36162f
C167 VP.n30 B 1.32492f
C168 VP.n31 B 1.35096f
C169 VP.n32 B 0.040636f
C170 VP.n33 B 0.054891f
C171 VP.n34 B 0.047571f
C172 VP.n35 B 0.042418f
C173 VP.n36 B 0.030822f
C174 VP.n37 B 0.030822f
C175 VP.n38 B 0.030822f
C176 VP.n39 B 0.029933f
C177 VP.n40 B 0.255721f
C178 VP.n41 B 0.056592f
C179 VP.n42 B 0.044995f
C180 VP.n43 B 0.030822f
C181 VP.n44 B 0.030822f
C182 VP.n45 B 0.030822f
C183 VP.n46 B 0.056592f
C184 VP.n47 B 0.255721f
C185 VP.n48 B 0.029933f
C186 VP.n49 B 0.057444f
C187 VP.n50 B 0.030822f
C188 VP.n51 B 0.030822f
C189 VP.n52 B 0.030822f
C190 VP.n53 B 0.047571f
C191 VP.n54 B 0.054891f
C192 VP.n55 B 0.36162f
C193 VP.n56 B 0.035599f
.ends

