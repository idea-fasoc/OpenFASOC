* NGSPICE file created from diff_pair_sample_0160.ext - technology: sky130A

.subckt diff_pair_sample_0160 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=2.2503 pd=12.32 as=0 ps=0 w=5.77 l=1.33
X1 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=2.2503 pd=12.32 as=0 ps=0 w=5.77 l=1.33
X2 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2503 pd=12.32 as=2.2503 ps=12.32 w=5.77 l=1.33
X3 VDD1.t1 VP.t0 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.2503 pd=12.32 as=2.2503 ps=12.32 w=5.77 l=1.33
X4 VDD1.t0 VP.t1 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2503 pd=12.32 as=2.2503 ps=12.32 w=5.77 l=1.33
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.2503 pd=12.32 as=0 ps=0 w=5.77 l=1.33
X6 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.2503 pd=12.32 as=2.2503 ps=12.32 w=5.77 l=1.33
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.2503 pd=12.32 as=0 ps=0 w=5.77 l=1.33
R0 B.n327 B.n326 585
R1 B.n329 B.n69 585
R2 B.n332 B.n331 585
R3 B.n333 B.n68 585
R4 B.n335 B.n334 585
R5 B.n337 B.n67 585
R6 B.n340 B.n339 585
R7 B.n341 B.n66 585
R8 B.n343 B.n342 585
R9 B.n345 B.n65 585
R10 B.n348 B.n347 585
R11 B.n349 B.n64 585
R12 B.n351 B.n350 585
R13 B.n353 B.n63 585
R14 B.n356 B.n355 585
R15 B.n357 B.n62 585
R16 B.n359 B.n358 585
R17 B.n361 B.n61 585
R18 B.n364 B.n363 585
R19 B.n365 B.n60 585
R20 B.n367 B.n366 585
R21 B.n369 B.n59 585
R22 B.n372 B.n371 585
R23 B.n374 B.n56 585
R24 B.n376 B.n375 585
R25 B.n378 B.n55 585
R26 B.n381 B.n380 585
R27 B.n382 B.n54 585
R28 B.n384 B.n383 585
R29 B.n386 B.n53 585
R30 B.n389 B.n388 585
R31 B.n390 B.n49 585
R32 B.n392 B.n391 585
R33 B.n394 B.n48 585
R34 B.n397 B.n396 585
R35 B.n398 B.n47 585
R36 B.n400 B.n399 585
R37 B.n402 B.n46 585
R38 B.n405 B.n404 585
R39 B.n406 B.n45 585
R40 B.n408 B.n407 585
R41 B.n410 B.n44 585
R42 B.n413 B.n412 585
R43 B.n414 B.n43 585
R44 B.n416 B.n415 585
R45 B.n418 B.n42 585
R46 B.n421 B.n420 585
R47 B.n422 B.n41 585
R48 B.n424 B.n423 585
R49 B.n426 B.n40 585
R50 B.n429 B.n428 585
R51 B.n430 B.n39 585
R52 B.n432 B.n431 585
R53 B.n434 B.n38 585
R54 B.n437 B.n436 585
R55 B.n438 B.n37 585
R56 B.n325 B.n35 585
R57 B.n441 B.n35 585
R58 B.n324 B.n34 585
R59 B.n442 B.n34 585
R60 B.n323 B.n33 585
R61 B.n443 B.n33 585
R62 B.n322 B.n321 585
R63 B.n321 B.n29 585
R64 B.n320 B.n28 585
R65 B.n449 B.n28 585
R66 B.n319 B.n27 585
R67 B.n450 B.n27 585
R68 B.n318 B.n26 585
R69 B.n451 B.n26 585
R70 B.n317 B.n316 585
R71 B.n316 B.n22 585
R72 B.n315 B.n21 585
R73 B.n457 B.n21 585
R74 B.n314 B.n20 585
R75 B.n458 B.n20 585
R76 B.n313 B.n19 585
R77 B.n459 B.n19 585
R78 B.n312 B.n311 585
R79 B.n311 B.n15 585
R80 B.n310 B.n14 585
R81 B.n465 B.n14 585
R82 B.n309 B.n13 585
R83 B.n466 B.n13 585
R84 B.n308 B.n12 585
R85 B.n467 B.n12 585
R86 B.n307 B.n306 585
R87 B.n306 B.n8 585
R88 B.n305 B.n7 585
R89 B.n473 B.n7 585
R90 B.n304 B.n6 585
R91 B.n474 B.n6 585
R92 B.n303 B.n5 585
R93 B.n475 B.n5 585
R94 B.n302 B.n301 585
R95 B.n301 B.n4 585
R96 B.n300 B.n70 585
R97 B.n300 B.n299 585
R98 B.n290 B.n71 585
R99 B.n72 B.n71 585
R100 B.n292 B.n291 585
R101 B.n293 B.n292 585
R102 B.n289 B.n76 585
R103 B.n80 B.n76 585
R104 B.n288 B.n287 585
R105 B.n287 B.n286 585
R106 B.n78 B.n77 585
R107 B.n79 B.n78 585
R108 B.n279 B.n278 585
R109 B.n280 B.n279 585
R110 B.n277 B.n85 585
R111 B.n85 B.n84 585
R112 B.n276 B.n275 585
R113 B.n275 B.n274 585
R114 B.n87 B.n86 585
R115 B.n88 B.n87 585
R116 B.n267 B.n266 585
R117 B.n268 B.n267 585
R118 B.n265 B.n92 585
R119 B.n96 B.n92 585
R120 B.n264 B.n263 585
R121 B.n263 B.n262 585
R122 B.n94 B.n93 585
R123 B.n95 B.n94 585
R124 B.n255 B.n254 585
R125 B.n256 B.n255 585
R126 B.n253 B.n101 585
R127 B.n101 B.n100 585
R128 B.n252 B.n251 585
R129 B.n251 B.n250 585
R130 B.n247 B.n105 585
R131 B.n246 B.n245 585
R132 B.n243 B.n106 585
R133 B.n243 B.n104 585
R134 B.n242 B.n241 585
R135 B.n240 B.n239 585
R136 B.n238 B.n108 585
R137 B.n236 B.n235 585
R138 B.n234 B.n109 585
R139 B.n233 B.n232 585
R140 B.n230 B.n110 585
R141 B.n228 B.n227 585
R142 B.n226 B.n111 585
R143 B.n225 B.n224 585
R144 B.n222 B.n112 585
R145 B.n220 B.n219 585
R146 B.n218 B.n113 585
R147 B.n217 B.n216 585
R148 B.n214 B.n114 585
R149 B.n212 B.n211 585
R150 B.n210 B.n115 585
R151 B.n209 B.n208 585
R152 B.n206 B.n116 585
R153 B.n204 B.n203 585
R154 B.n201 B.n117 585
R155 B.n200 B.n199 585
R156 B.n197 B.n120 585
R157 B.n195 B.n194 585
R158 B.n193 B.n121 585
R159 B.n192 B.n191 585
R160 B.n189 B.n122 585
R161 B.n187 B.n186 585
R162 B.n185 B.n123 585
R163 B.n184 B.n183 585
R164 B.n181 B.n180 585
R165 B.n179 B.n178 585
R166 B.n177 B.n128 585
R167 B.n175 B.n174 585
R168 B.n173 B.n129 585
R169 B.n172 B.n171 585
R170 B.n169 B.n130 585
R171 B.n167 B.n166 585
R172 B.n165 B.n131 585
R173 B.n164 B.n163 585
R174 B.n161 B.n132 585
R175 B.n159 B.n158 585
R176 B.n157 B.n133 585
R177 B.n156 B.n155 585
R178 B.n153 B.n134 585
R179 B.n151 B.n150 585
R180 B.n149 B.n135 585
R181 B.n148 B.n147 585
R182 B.n145 B.n136 585
R183 B.n143 B.n142 585
R184 B.n141 B.n137 585
R185 B.n140 B.n139 585
R186 B.n103 B.n102 585
R187 B.n104 B.n103 585
R188 B.n249 B.n248 585
R189 B.n250 B.n249 585
R190 B.n99 B.n98 585
R191 B.n100 B.n99 585
R192 B.n258 B.n257 585
R193 B.n257 B.n256 585
R194 B.n259 B.n97 585
R195 B.n97 B.n95 585
R196 B.n261 B.n260 585
R197 B.n262 B.n261 585
R198 B.n91 B.n90 585
R199 B.n96 B.n91 585
R200 B.n270 B.n269 585
R201 B.n269 B.n268 585
R202 B.n271 B.n89 585
R203 B.n89 B.n88 585
R204 B.n273 B.n272 585
R205 B.n274 B.n273 585
R206 B.n83 B.n82 585
R207 B.n84 B.n83 585
R208 B.n282 B.n281 585
R209 B.n281 B.n280 585
R210 B.n283 B.n81 585
R211 B.n81 B.n79 585
R212 B.n285 B.n284 585
R213 B.n286 B.n285 585
R214 B.n75 B.n74 585
R215 B.n80 B.n75 585
R216 B.n295 B.n294 585
R217 B.n294 B.n293 585
R218 B.n296 B.n73 585
R219 B.n73 B.n72 585
R220 B.n298 B.n297 585
R221 B.n299 B.n298 585
R222 B.n2 B.n0 585
R223 B.n4 B.n2 585
R224 B.n3 B.n1 585
R225 B.n474 B.n3 585
R226 B.n472 B.n471 585
R227 B.n473 B.n472 585
R228 B.n470 B.n9 585
R229 B.n9 B.n8 585
R230 B.n469 B.n468 585
R231 B.n468 B.n467 585
R232 B.n11 B.n10 585
R233 B.n466 B.n11 585
R234 B.n464 B.n463 585
R235 B.n465 B.n464 585
R236 B.n462 B.n16 585
R237 B.n16 B.n15 585
R238 B.n461 B.n460 585
R239 B.n460 B.n459 585
R240 B.n18 B.n17 585
R241 B.n458 B.n18 585
R242 B.n456 B.n455 585
R243 B.n457 B.n456 585
R244 B.n454 B.n23 585
R245 B.n23 B.n22 585
R246 B.n453 B.n452 585
R247 B.n452 B.n451 585
R248 B.n25 B.n24 585
R249 B.n450 B.n25 585
R250 B.n448 B.n447 585
R251 B.n449 B.n448 585
R252 B.n446 B.n30 585
R253 B.n30 B.n29 585
R254 B.n445 B.n444 585
R255 B.n444 B.n443 585
R256 B.n32 B.n31 585
R257 B.n442 B.n32 585
R258 B.n440 B.n439 585
R259 B.n441 B.n440 585
R260 B.n477 B.n476 585
R261 B.n476 B.n475 585
R262 B.n249 B.n105 492.5
R263 B.n440 B.n37 492.5
R264 B.n251 B.n103 492.5
R265 B.n327 B.n35 492.5
R266 B.n124 B.t13 309.3
R267 B.n118 B.t6 309.3
R268 B.n50 B.t2 309.3
R269 B.n57 B.t10 309.3
R270 B.n328 B.n36 256.663
R271 B.n330 B.n36 256.663
R272 B.n336 B.n36 256.663
R273 B.n338 B.n36 256.663
R274 B.n344 B.n36 256.663
R275 B.n346 B.n36 256.663
R276 B.n352 B.n36 256.663
R277 B.n354 B.n36 256.663
R278 B.n360 B.n36 256.663
R279 B.n362 B.n36 256.663
R280 B.n368 B.n36 256.663
R281 B.n370 B.n36 256.663
R282 B.n377 B.n36 256.663
R283 B.n379 B.n36 256.663
R284 B.n385 B.n36 256.663
R285 B.n387 B.n36 256.663
R286 B.n393 B.n36 256.663
R287 B.n395 B.n36 256.663
R288 B.n401 B.n36 256.663
R289 B.n403 B.n36 256.663
R290 B.n409 B.n36 256.663
R291 B.n411 B.n36 256.663
R292 B.n417 B.n36 256.663
R293 B.n419 B.n36 256.663
R294 B.n425 B.n36 256.663
R295 B.n427 B.n36 256.663
R296 B.n433 B.n36 256.663
R297 B.n435 B.n36 256.663
R298 B.n244 B.n104 256.663
R299 B.n107 B.n104 256.663
R300 B.n237 B.n104 256.663
R301 B.n231 B.n104 256.663
R302 B.n229 B.n104 256.663
R303 B.n223 B.n104 256.663
R304 B.n221 B.n104 256.663
R305 B.n215 B.n104 256.663
R306 B.n213 B.n104 256.663
R307 B.n207 B.n104 256.663
R308 B.n205 B.n104 256.663
R309 B.n198 B.n104 256.663
R310 B.n196 B.n104 256.663
R311 B.n190 B.n104 256.663
R312 B.n188 B.n104 256.663
R313 B.n182 B.n104 256.663
R314 B.n127 B.n104 256.663
R315 B.n176 B.n104 256.663
R316 B.n170 B.n104 256.663
R317 B.n168 B.n104 256.663
R318 B.n162 B.n104 256.663
R319 B.n160 B.n104 256.663
R320 B.n154 B.n104 256.663
R321 B.n152 B.n104 256.663
R322 B.n146 B.n104 256.663
R323 B.n144 B.n104 256.663
R324 B.n138 B.n104 256.663
R325 B.n249 B.n99 163.367
R326 B.n257 B.n99 163.367
R327 B.n257 B.n97 163.367
R328 B.n261 B.n97 163.367
R329 B.n261 B.n91 163.367
R330 B.n269 B.n91 163.367
R331 B.n269 B.n89 163.367
R332 B.n273 B.n89 163.367
R333 B.n273 B.n83 163.367
R334 B.n281 B.n83 163.367
R335 B.n281 B.n81 163.367
R336 B.n285 B.n81 163.367
R337 B.n285 B.n75 163.367
R338 B.n294 B.n75 163.367
R339 B.n294 B.n73 163.367
R340 B.n298 B.n73 163.367
R341 B.n298 B.n2 163.367
R342 B.n476 B.n2 163.367
R343 B.n476 B.n3 163.367
R344 B.n472 B.n3 163.367
R345 B.n472 B.n9 163.367
R346 B.n468 B.n9 163.367
R347 B.n468 B.n11 163.367
R348 B.n464 B.n11 163.367
R349 B.n464 B.n16 163.367
R350 B.n460 B.n16 163.367
R351 B.n460 B.n18 163.367
R352 B.n456 B.n18 163.367
R353 B.n456 B.n23 163.367
R354 B.n452 B.n23 163.367
R355 B.n452 B.n25 163.367
R356 B.n448 B.n25 163.367
R357 B.n448 B.n30 163.367
R358 B.n444 B.n30 163.367
R359 B.n444 B.n32 163.367
R360 B.n440 B.n32 163.367
R361 B.n245 B.n243 163.367
R362 B.n243 B.n242 163.367
R363 B.n239 B.n238 163.367
R364 B.n236 B.n109 163.367
R365 B.n232 B.n230 163.367
R366 B.n228 B.n111 163.367
R367 B.n224 B.n222 163.367
R368 B.n220 B.n113 163.367
R369 B.n216 B.n214 163.367
R370 B.n212 B.n115 163.367
R371 B.n208 B.n206 163.367
R372 B.n204 B.n117 163.367
R373 B.n199 B.n197 163.367
R374 B.n195 B.n121 163.367
R375 B.n191 B.n189 163.367
R376 B.n187 B.n123 163.367
R377 B.n183 B.n181 163.367
R378 B.n178 B.n177 163.367
R379 B.n175 B.n129 163.367
R380 B.n171 B.n169 163.367
R381 B.n167 B.n131 163.367
R382 B.n163 B.n161 163.367
R383 B.n159 B.n133 163.367
R384 B.n155 B.n153 163.367
R385 B.n151 B.n135 163.367
R386 B.n147 B.n145 163.367
R387 B.n143 B.n137 163.367
R388 B.n139 B.n103 163.367
R389 B.n251 B.n101 163.367
R390 B.n255 B.n101 163.367
R391 B.n255 B.n94 163.367
R392 B.n263 B.n94 163.367
R393 B.n263 B.n92 163.367
R394 B.n267 B.n92 163.367
R395 B.n267 B.n87 163.367
R396 B.n275 B.n87 163.367
R397 B.n275 B.n85 163.367
R398 B.n279 B.n85 163.367
R399 B.n279 B.n78 163.367
R400 B.n287 B.n78 163.367
R401 B.n287 B.n76 163.367
R402 B.n292 B.n76 163.367
R403 B.n292 B.n71 163.367
R404 B.n300 B.n71 163.367
R405 B.n301 B.n300 163.367
R406 B.n301 B.n5 163.367
R407 B.n6 B.n5 163.367
R408 B.n7 B.n6 163.367
R409 B.n306 B.n7 163.367
R410 B.n306 B.n12 163.367
R411 B.n13 B.n12 163.367
R412 B.n14 B.n13 163.367
R413 B.n311 B.n14 163.367
R414 B.n311 B.n19 163.367
R415 B.n20 B.n19 163.367
R416 B.n21 B.n20 163.367
R417 B.n316 B.n21 163.367
R418 B.n316 B.n26 163.367
R419 B.n27 B.n26 163.367
R420 B.n28 B.n27 163.367
R421 B.n321 B.n28 163.367
R422 B.n321 B.n33 163.367
R423 B.n34 B.n33 163.367
R424 B.n35 B.n34 163.367
R425 B.n436 B.n434 163.367
R426 B.n432 B.n39 163.367
R427 B.n428 B.n426 163.367
R428 B.n424 B.n41 163.367
R429 B.n420 B.n418 163.367
R430 B.n416 B.n43 163.367
R431 B.n412 B.n410 163.367
R432 B.n408 B.n45 163.367
R433 B.n404 B.n402 163.367
R434 B.n400 B.n47 163.367
R435 B.n396 B.n394 163.367
R436 B.n392 B.n49 163.367
R437 B.n388 B.n386 163.367
R438 B.n384 B.n54 163.367
R439 B.n380 B.n378 163.367
R440 B.n376 B.n56 163.367
R441 B.n371 B.n369 163.367
R442 B.n367 B.n60 163.367
R443 B.n363 B.n361 163.367
R444 B.n359 B.n62 163.367
R445 B.n355 B.n353 163.367
R446 B.n351 B.n64 163.367
R447 B.n347 B.n345 163.367
R448 B.n343 B.n66 163.367
R449 B.n339 B.n337 163.367
R450 B.n335 B.n68 163.367
R451 B.n331 B.n329 163.367
R452 B.n250 B.n104 114.531
R453 B.n441 B.n36 114.531
R454 B.n124 B.t15 108.189
R455 B.n57 B.t11 108.189
R456 B.n118 B.t9 108.184
R457 B.n50 B.t4 108.184
R458 B.n125 B.t14 75.9959
R459 B.n58 B.t12 75.9959
R460 B.n119 B.t8 75.9901
R461 B.n51 B.t5 75.9901
R462 B.n244 B.n105 71.676
R463 B.n242 B.n107 71.676
R464 B.n238 B.n237 71.676
R465 B.n231 B.n109 71.676
R466 B.n230 B.n229 71.676
R467 B.n223 B.n111 71.676
R468 B.n222 B.n221 71.676
R469 B.n215 B.n113 71.676
R470 B.n214 B.n213 71.676
R471 B.n207 B.n115 71.676
R472 B.n206 B.n205 71.676
R473 B.n198 B.n117 71.676
R474 B.n197 B.n196 71.676
R475 B.n190 B.n121 71.676
R476 B.n189 B.n188 71.676
R477 B.n182 B.n123 71.676
R478 B.n181 B.n127 71.676
R479 B.n177 B.n176 71.676
R480 B.n170 B.n129 71.676
R481 B.n169 B.n168 71.676
R482 B.n162 B.n131 71.676
R483 B.n161 B.n160 71.676
R484 B.n154 B.n133 71.676
R485 B.n153 B.n152 71.676
R486 B.n146 B.n135 71.676
R487 B.n145 B.n144 71.676
R488 B.n138 B.n137 71.676
R489 B.n435 B.n37 71.676
R490 B.n434 B.n433 71.676
R491 B.n427 B.n39 71.676
R492 B.n426 B.n425 71.676
R493 B.n419 B.n41 71.676
R494 B.n418 B.n417 71.676
R495 B.n411 B.n43 71.676
R496 B.n410 B.n409 71.676
R497 B.n403 B.n45 71.676
R498 B.n402 B.n401 71.676
R499 B.n395 B.n47 71.676
R500 B.n394 B.n393 71.676
R501 B.n387 B.n49 71.676
R502 B.n386 B.n385 71.676
R503 B.n379 B.n54 71.676
R504 B.n378 B.n377 71.676
R505 B.n370 B.n56 71.676
R506 B.n369 B.n368 71.676
R507 B.n362 B.n60 71.676
R508 B.n361 B.n360 71.676
R509 B.n354 B.n62 71.676
R510 B.n353 B.n352 71.676
R511 B.n346 B.n64 71.676
R512 B.n345 B.n344 71.676
R513 B.n338 B.n66 71.676
R514 B.n337 B.n336 71.676
R515 B.n330 B.n68 71.676
R516 B.n329 B.n328 71.676
R517 B.n328 B.n327 71.676
R518 B.n331 B.n330 71.676
R519 B.n336 B.n335 71.676
R520 B.n339 B.n338 71.676
R521 B.n344 B.n343 71.676
R522 B.n347 B.n346 71.676
R523 B.n352 B.n351 71.676
R524 B.n355 B.n354 71.676
R525 B.n360 B.n359 71.676
R526 B.n363 B.n362 71.676
R527 B.n368 B.n367 71.676
R528 B.n371 B.n370 71.676
R529 B.n377 B.n376 71.676
R530 B.n380 B.n379 71.676
R531 B.n385 B.n384 71.676
R532 B.n388 B.n387 71.676
R533 B.n393 B.n392 71.676
R534 B.n396 B.n395 71.676
R535 B.n401 B.n400 71.676
R536 B.n404 B.n403 71.676
R537 B.n409 B.n408 71.676
R538 B.n412 B.n411 71.676
R539 B.n417 B.n416 71.676
R540 B.n420 B.n419 71.676
R541 B.n425 B.n424 71.676
R542 B.n428 B.n427 71.676
R543 B.n433 B.n432 71.676
R544 B.n436 B.n435 71.676
R545 B.n245 B.n244 71.676
R546 B.n239 B.n107 71.676
R547 B.n237 B.n236 71.676
R548 B.n232 B.n231 71.676
R549 B.n229 B.n228 71.676
R550 B.n224 B.n223 71.676
R551 B.n221 B.n220 71.676
R552 B.n216 B.n215 71.676
R553 B.n213 B.n212 71.676
R554 B.n208 B.n207 71.676
R555 B.n205 B.n204 71.676
R556 B.n199 B.n198 71.676
R557 B.n196 B.n195 71.676
R558 B.n191 B.n190 71.676
R559 B.n188 B.n187 71.676
R560 B.n183 B.n182 71.676
R561 B.n178 B.n127 71.676
R562 B.n176 B.n175 71.676
R563 B.n171 B.n170 71.676
R564 B.n168 B.n167 71.676
R565 B.n163 B.n162 71.676
R566 B.n160 B.n159 71.676
R567 B.n155 B.n154 71.676
R568 B.n152 B.n151 71.676
R569 B.n147 B.n146 71.676
R570 B.n144 B.n143 71.676
R571 B.n139 B.n138 71.676
R572 B.n250 B.n100 67.7235
R573 B.n256 B.n100 67.7235
R574 B.n256 B.n95 67.7235
R575 B.n262 B.n95 67.7235
R576 B.n262 B.n96 67.7235
R577 B.n268 B.n88 67.7235
R578 B.n274 B.n88 67.7235
R579 B.n274 B.n84 67.7235
R580 B.n280 B.n84 67.7235
R581 B.n280 B.n79 67.7235
R582 B.n286 B.n79 67.7235
R583 B.n286 B.n80 67.7235
R584 B.n293 B.n72 67.7235
R585 B.n299 B.n72 67.7235
R586 B.n299 B.n4 67.7235
R587 B.n475 B.n4 67.7235
R588 B.n475 B.n474 67.7235
R589 B.n474 B.n473 67.7235
R590 B.n473 B.n8 67.7235
R591 B.n467 B.n8 67.7235
R592 B.n466 B.n465 67.7235
R593 B.n465 B.n15 67.7235
R594 B.n459 B.n15 67.7235
R595 B.n459 B.n458 67.7235
R596 B.n458 B.n457 67.7235
R597 B.n457 B.n22 67.7235
R598 B.n451 B.n22 67.7235
R599 B.n450 B.n449 67.7235
R600 B.n449 B.n29 67.7235
R601 B.n443 B.n29 67.7235
R602 B.n443 B.n442 67.7235
R603 B.n442 B.n441 67.7235
R604 B.n80 B.t1 64.7357
R605 B.t0 B.n466 64.7357
R606 B.n126 B.n125 59.5399
R607 B.n202 B.n119 59.5399
R608 B.n52 B.n51 59.5399
R609 B.n373 B.n58 59.5399
R610 B.n96 B.t7 58.7601
R611 B.t3 B.n450 58.7601
R612 B.n125 B.n124 32.1944
R613 B.n119 B.n118 32.1944
R614 B.n51 B.n50 32.1944
R615 B.n58 B.n57 32.1944
R616 B.n439 B.n438 32.0005
R617 B.n326 B.n325 32.0005
R618 B.n252 B.n102 32.0005
R619 B.n248 B.n247 32.0005
R620 B B.n477 18.0485
R621 B.n438 B.n437 10.6151
R622 B.n437 B.n38 10.6151
R623 B.n431 B.n38 10.6151
R624 B.n431 B.n430 10.6151
R625 B.n430 B.n429 10.6151
R626 B.n429 B.n40 10.6151
R627 B.n423 B.n40 10.6151
R628 B.n423 B.n422 10.6151
R629 B.n422 B.n421 10.6151
R630 B.n421 B.n42 10.6151
R631 B.n415 B.n42 10.6151
R632 B.n415 B.n414 10.6151
R633 B.n414 B.n413 10.6151
R634 B.n413 B.n44 10.6151
R635 B.n407 B.n44 10.6151
R636 B.n407 B.n406 10.6151
R637 B.n406 B.n405 10.6151
R638 B.n405 B.n46 10.6151
R639 B.n399 B.n46 10.6151
R640 B.n399 B.n398 10.6151
R641 B.n398 B.n397 10.6151
R642 B.n397 B.n48 10.6151
R643 B.n391 B.n390 10.6151
R644 B.n390 B.n389 10.6151
R645 B.n389 B.n53 10.6151
R646 B.n383 B.n53 10.6151
R647 B.n383 B.n382 10.6151
R648 B.n382 B.n381 10.6151
R649 B.n381 B.n55 10.6151
R650 B.n375 B.n55 10.6151
R651 B.n375 B.n374 10.6151
R652 B.n372 B.n59 10.6151
R653 B.n366 B.n59 10.6151
R654 B.n366 B.n365 10.6151
R655 B.n365 B.n364 10.6151
R656 B.n364 B.n61 10.6151
R657 B.n358 B.n61 10.6151
R658 B.n358 B.n357 10.6151
R659 B.n357 B.n356 10.6151
R660 B.n356 B.n63 10.6151
R661 B.n350 B.n63 10.6151
R662 B.n350 B.n349 10.6151
R663 B.n349 B.n348 10.6151
R664 B.n348 B.n65 10.6151
R665 B.n342 B.n65 10.6151
R666 B.n342 B.n341 10.6151
R667 B.n341 B.n340 10.6151
R668 B.n340 B.n67 10.6151
R669 B.n334 B.n67 10.6151
R670 B.n334 B.n333 10.6151
R671 B.n333 B.n332 10.6151
R672 B.n332 B.n69 10.6151
R673 B.n326 B.n69 10.6151
R674 B.n253 B.n252 10.6151
R675 B.n254 B.n253 10.6151
R676 B.n254 B.n93 10.6151
R677 B.n264 B.n93 10.6151
R678 B.n265 B.n264 10.6151
R679 B.n266 B.n265 10.6151
R680 B.n266 B.n86 10.6151
R681 B.n276 B.n86 10.6151
R682 B.n277 B.n276 10.6151
R683 B.n278 B.n277 10.6151
R684 B.n278 B.n77 10.6151
R685 B.n288 B.n77 10.6151
R686 B.n289 B.n288 10.6151
R687 B.n291 B.n289 10.6151
R688 B.n291 B.n290 10.6151
R689 B.n290 B.n70 10.6151
R690 B.n302 B.n70 10.6151
R691 B.n303 B.n302 10.6151
R692 B.n304 B.n303 10.6151
R693 B.n305 B.n304 10.6151
R694 B.n307 B.n305 10.6151
R695 B.n308 B.n307 10.6151
R696 B.n309 B.n308 10.6151
R697 B.n310 B.n309 10.6151
R698 B.n312 B.n310 10.6151
R699 B.n313 B.n312 10.6151
R700 B.n314 B.n313 10.6151
R701 B.n315 B.n314 10.6151
R702 B.n317 B.n315 10.6151
R703 B.n318 B.n317 10.6151
R704 B.n319 B.n318 10.6151
R705 B.n320 B.n319 10.6151
R706 B.n322 B.n320 10.6151
R707 B.n323 B.n322 10.6151
R708 B.n324 B.n323 10.6151
R709 B.n325 B.n324 10.6151
R710 B.n247 B.n246 10.6151
R711 B.n246 B.n106 10.6151
R712 B.n241 B.n106 10.6151
R713 B.n241 B.n240 10.6151
R714 B.n240 B.n108 10.6151
R715 B.n235 B.n108 10.6151
R716 B.n235 B.n234 10.6151
R717 B.n234 B.n233 10.6151
R718 B.n233 B.n110 10.6151
R719 B.n227 B.n110 10.6151
R720 B.n227 B.n226 10.6151
R721 B.n226 B.n225 10.6151
R722 B.n225 B.n112 10.6151
R723 B.n219 B.n112 10.6151
R724 B.n219 B.n218 10.6151
R725 B.n218 B.n217 10.6151
R726 B.n217 B.n114 10.6151
R727 B.n211 B.n114 10.6151
R728 B.n211 B.n210 10.6151
R729 B.n210 B.n209 10.6151
R730 B.n209 B.n116 10.6151
R731 B.n203 B.n116 10.6151
R732 B.n201 B.n200 10.6151
R733 B.n200 B.n120 10.6151
R734 B.n194 B.n120 10.6151
R735 B.n194 B.n193 10.6151
R736 B.n193 B.n192 10.6151
R737 B.n192 B.n122 10.6151
R738 B.n186 B.n122 10.6151
R739 B.n186 B.n185 10.6151
R740 B.n185 B.n184 10.6151
R741 B.n180 B.n179 10.6151
R742 B.n179 B.n128 10.6151
R743 B.n174 B.n128 10.6151
R744 B.n174 B.n173 10.6151
R745 B.n173 B.n172 10.6151
R746 B.n172 B.n130 10.6151
R747 B.n166 B.n130 10.6151
R748 B.n166 B.n165 10.6151
R749 B.n165 B.n164 10.6151
R750 B.n164 B.n132 10.6151
R751 B.n158 B.n132 10.6151
R752 B.n158 B.n157 10.6151
R753 B.n157 B.n156 10.6151
R754 B.n156 B.n134 10.6151
R755 B.n150 B.n134 10.6151
R756 B.n150 B.n149 10.6151
R757 B.n149 B.n148 10.6151
R758 B.n148 B.n136 10.6151
R759 B.n142 B.n136 10.6151
R760 B.n142 B.n141 10.6151
R761 B.n141 B.n140 10.6151
R762 B.n140 B.n102 10.6151
R763 B.n248 B.n98 10.6151
R764 B.n258 B.n98 10.6151
R765 B.n259 B.n258 10.6151
R766 B.n260 B.n259 10.6151
R767 B.n260 B.n90 10.6151
R768 B.n270 B.n90 10.6151
R769 B.n271 B.n270 10.6151
R770 B.n272 B.n271 10.6151
R771 B.n272 B.n82 10.6151
R772 B.n282 B.n82 10.6151
R773 B.n283 B.n282 10.6151
R774 B.n284 B.n283 10.6151
R775 B.n284 B.n74 10.6151
R776 B.n295 B.n74 10.6151
R777 B.n296 B.n295 10.6151
R778 B.n297 B.n296 10.6151
R779 B.n297 B.n0 10.6151
R780 B.n471 B.n1 10.6151
R781 B.n471 B.n470 10.6151
R782 B.n470 B.n469 10.6151
R783 B.n469 B.n10 10.6151
R784 B.n463 B.n10 10.6151
R785 B.n463 B.n462 10.6151
R786 B.n462 B.n461 10.6151
R787 B.n461 B.n17 10.6151
R788 B.n455 B.n17 10.6151
R789 B.n455 B.n454 10.6151
R790 B.n454 B.n453 10.6151
R791 B.n453 B.n24 10.6151
R792 B.n447 B.n24 10.6151
R793 B.n447 B.n446 10.6151
R794 B.n446 B.n445 10.6151
R795 B.n445 B.n31 10.6151
R796 B.n439 B.n31 10.6151
R797 B.n52 B.n48 9.36635
R798 B.n373 B.n372 9.36635
R799 B.n203 B.n202 9.36635
R800 B.n180 B.n126 9.36635
R801 B.n268 B.t7 8.96383
R802 B.n451 B.t3 8.96383
R803 B.n293 B.t1 2.98828
R804 B.n467 B.t0 2.98828
R805 B.n477 B.n0 2.81026
R806 B.n477 B.n1 2.81026
R807 B.n391 B.n52 1.24928
R808 B.n374 B.n373 1.24928
R809 B.n202 B.n201 1.24928
R810 B.n184 B.n126 1.24928
R811 VN VN.t0 251.73
R812 VN VN.t1 215.022
R813 VTAIL.n1 VTAIL.t3 57.144
R814 VTAIL.n3 VTAIL.t2 57.1438
R815 VTAIL.n0 VTAIL.t0 57.1438
R816 VTAIL.n2 VTAIL.t1 57.1438
R817 VTAIL.n1 VTAIL.n0 20.2031
R818 VTAIL.n3 VTAIL.n2 18.7721
R819 VTAIL.n2 VTAIL.n1 1.18584
R820 VTAIL VTAIL.n0 0.886276
R821 VTAIL VTAIL.n3 0.300069
R822 VDD2.n0 VDD2.t0 105.319
R823 VDD2.n0 VDD2.t1 73.8226
R824 VDD2 VDD2.n0 0.416448
R825 VP.n0 VP.t0 251.445
R826 VP.n0 VP.t1 214.875
R827 VP VP.n0 0.146778
R828 VDD1 VDD1.t0 106.201
R829 VDD1 VDD1.t1 74.2385
C0 VTAIL VDD2 3.25323f
C1 VP VN 3.70618f
C2 VDD2 VDD1 0.526126f
C3 VP VTAIL 1.20921f
C4 VTAIL VN 1.19493f
C5 VP VDD1 1.42355f
C6 VP VDD2 0.279145f
C7 VN VDD1 0.14754f
C8 VN VDD2 1.29377f
C9 VTAIL VDD1 3.21071f
C10 VDD2 B 2.836915f
C11 VDD1 B 4.51702f
C12 VTAIL B 4.119613f
C13 VN B 6.4788f
C14 VP B 4.306636f
C15 VDD1.t1 B 0.693845f
C16 VDD1.t0 B 0.921695f
C17 VP.t0 B 0.890505f
C18 VP.t1 B 0.72955f
C19 VP.n0 B 2.05386f
C20 VDD2.t0 B 0.949754f
C21 VDD2.t1 B 0.726598f
C22 VDD2.n0 B 1.56824f
C23 VTAIL.t0 B 0.755437f
C24 VTAIL.n0 B 0.891934f
C25 VTAIL.t3 B 0.75544f
C26 VTAIL.n1 B 0.908043f
C27 VTAIL.t1 B 0.755437f
C28 VTAIL.n2 B 0.831079f
C29 VTAIL.t2 B 0.755437f
C30 VTAIL.n3 B 0.783438f
C31 VN.t1 B 0.722025f
C32 VN.t0 B 0.884535f
.ends

