* NGSPICE file created from diff_pair_sample_1587.ext - technology: sky130A

.subckt diff_pair_sample_1587 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t5 w_n4320_n2126# sky130_fd_pr__pfet_01v8 ad=0.95535 pd=6.12 as=0.95535 ps=6.12 w=5.79 l=3.02
X1 VTAIL.t6 VN.t0 VDD2.t7 w_n4320_n2126# sky130_fd_pr__pfet_01v8 ad=2.2581 pd=12.36 as=0.95535 ps=6.12 w=5.79 l=3.02
X2 VTAIL.t7 VN.t1 VDD2.t6 w_n4320_n2126# sky130_fd_pr__pfet_01v8 ad=0.95535 pd=6.12 as=0.95535 ps=6.12 w=5.79 l=3.02
X3 B.t11 B.t9 B.t10 w_n4320_n2126# sky130_fd_pr__pfet_01v8 ad=2.2581 pd=12.36 as=0 ps=0 w=5.79 l=3.02
X4 VTAIL.t5 VN.t2 VDD2.t5 w_n4320_n2126# sky130_fd_pr__pfet_01v8 ad=0.95535 pd=6.12 as=0.95535 ps=6.12 w=5.79 l=3.02
X5 VTAIL.t14 VP.t1 VDD1.t1 w_n4320_n2126# sky130_fd_pr__pfet_01v8 ad=2.2581 pd=12.36 as=0.95535 ps=6.12 w=5.79 l=3.02
X6 VDD2.t4 VN.t3 VTAIL.t1 w_n4320_n2126# sky130_fd_pr__pfet_01v8 ad=0.95535 pd=6.12 as=2.2581 ps=12.36 w=5.79 l=3.02
X7 VDD2.t3 VN.t4 VTAIL.t2 w_n4320_n2126# sky130_fd_pr__pfet_01v8 ad=0.95535 pd=6.12 as=2.2581 ps=12.36 w=5.79 l=3.02
X8 VTAIL.t0 VN.t5 VDD2.t2 w_n4320_n2126# sky130_fd_pr__pfet_01v8 ad=2.2581 pd=12.36 as=0.95535 ps=6.12 w=5.79 l=3.02
X9 B.t8 B.t6 B.t7 w_n4320_n2126# sky130_fd_pr__pfet_01v8 ad=2.2581 pd=12.36 as=0 ps=0 w=5.79 l=3.02
X10 VDD2.t1 VN.t6 VTAIL.t3 w_n4320_n2126# sky130_fd_pr__pfet_01v8 ad=0.95535 pd=6.12 as=0.95535 ps=6.12 w=5.79 l=3.02
X11 VDD1.t2 VP.t2 VTAIL.t13 w_n4320_n2126# sky130_fd_pr__pfet_01v8 ad=0.95535 pd=6.12 as=0.95535 ps=6.12 w=5.79 l=3.02
X12 VTAIL.t12 VP.t3 VDD1.t0 w_n4320_n2126# sky130_fd_pr__pfet_01v8 ad=2.2581 pd=12.36 as=0.95535 ps=6.12 w=5.79 l=3.02
X13 VDD2.t0 VN.t7 VTAIL.t4 w_n4320_n2126# sky130_fd_pr__pfet_01v8 ad=0.95535 pd=6.12 as=0.95535 ps=6.12 w=5.79 l=3.02
X14 B.t5 B.t3 B.t4 w_n4320_n2126# sky130_fd_pr__pfet_01v8 ad=2.2581 pd=12.36 as=0 ps=0 w=5.79 l=3.02
X15 VDD1.t6 VP.t4 VTAIL.t11 w_n4320_n2126# sky130_fd_pr__pfet_01v8 ad=0.95535 pd=6.12 as=2.2581 ps=12.36 w=5.79 l=3.02
X16 VDD1.t4 VP.t5 VTAIL.t10 w_n4320_n2126# sky130_fd_pr__pfet_01v8 ad=0.95535 pd=6.12 as=0.95535 ps=6.12 w=5.79 l=3.02
X17 VDD1.t3 VP.t6 VTAIL.t9 w_n4320_n2126# sky130_fd_pr__pfet_01v8 ad=0.95535 pd=6.12 as=2.2581 ps=12.36 w=5.79 l=3.02
X18 VTAIL.t8 VP.t7 VDD1.t7 w_n4320_n2126# sky130_fd_pr__pfet_01v8 ad=0.95535 pd=6.12 as=0.95535 ps=6.12 w=5.79 l=3.02
X19 B.t2 B.t0 B.t1 w_n4320_n2126# sky130_fd_pr__pfet_01v8 ad=2.2581 pd=12.36 as=0 ps=0 w=5.79 l=3.02
R0 VP.n22 VP.n21 161.3
R1 VP.n23 VP.n18 161.3
R2 VP.n25 VP.n24 161.3
R3 VP.n26 VP.n17 161.3
R4 VP.n28 VP.n27 161.3
R5 VP.n29 VP.n16 161.3
R6 VP.n32 VP.n31 161.3
R7 VP.n33 VP.n15 161.3
R8 VP.n35 VP.n34 161.3
R9 VP.n36 VP.n14 161.3
R10 VP.n38 VP.n37 161.3
R11 VP.n39 VP.n13 161.3
R12 VP.n41 VP.n40 161.3
R13 VP.n42 VP.n12 161.3
R14 VP.n78 VP.n0 161.3
R15 VP.n77 VP.n76 161.3
R16 VP.n75 VP.n1 161.3
R17 VP.n74 VP.n73 161.3
R18 VP.n72 VP.n2 161.3
R19 VP.n71 VP.n70 161.3
R20 VP.n69 VP.n3 161.3
R21 VP.n68 VP.n67 161.3
R22 VP.n65 VP.n4 161.3
R23 VP.n64 VP.n63 161.3
R24 VP.n62 VP.n5 161.3
R25 VP.n61 VP.n60 161.3
R26 VP.n59 VP.n6 161.3
R27 VP.n58 VP.n57 161.3
R28 VP.n56 VP.n55 161.3
R29 VP.n54 VP.n8 161.3
R30 VP.n53 VP.n52 161.3
R31 VP.n51 VP.n9 161.3
R32 VP.n50 VP.n49 161.3
R33 VP.n48 VP.n10 161.3
R34 VP.n47 VP.n46 161.3
R35 VP.n45 VP.n11 109.534
R36 VP.n80 VP.n79 109.534
R37 VP.n44 VP.n43 109.534
R38 VP.n20 VP.t1 78.4735
R39 VP.n20 VP.n19 65.4202
R40 VP.n53 VP.n9 55.0624
R41 VP.n73 VP.n72 55.0624
R42 VP.n37 VP.n36 55.0624
R43 VP.n45 VP.n44 48.1435
R44 VP.n11 VP.t3 46.2055
R45 VP.n7 VP.t2 46.2055
R46 VP.n66 VP.t7 46.2055
R47 VP.n79 VP.t6 46.2055
R48 VP.n43 VP.t4 46.2055
R49 VP.n30 VP.t0 46.2055
R50 VP.n19 VP.t5 46.2055
R51 VP.n60 VP.n5 40.4934
R52 VP.n64 VP.n5 40.4934
R53 VP.n28 VP.n17 40.4934
R54 VP.n24 VP.n17 40.4934
R55 VP.n49 VP.n9 25.9244
R56 VP.n73 VP.n1 25.9244
R57 VP.n37 VP.n13 25.9244
R58 VP.n48 VP.n47 24.4675
R59 VP.n49 VP.n48 24.4675
R60 VP.n54 VP.n53 24.4675
R61 VP.n55 VP.n54 24.4675
R62 VP.n59 VP.n58 24.4675
R63 VP.n60 VP.n59 24.4675
R64 VP.n65 VP.n64 24.4675
R65 VP.n67 VP.n65 24.4675
R66 VP.n71 VP.n3 24.4675
R67 VP.n72 VP.n71 24.4675
R68 VP.n77 VP.n1 24.4675
R69 VP.n78 VP.n77 24.4675
R70 VP.n41 VP.n13 24.4675
R71 VP.n42 VP.n41 24.4675
R72 VP.n29 VP.n28 24.4675
R73 VP.n31 VP.n29 24.4675
R74 VP.n35 VP.n15 24.4675
R75 VP.n36 VP.n35 24.4675
R76 VP.n23 VP.n22 24.4675
R77 VP.n24 VP.n23 24.4675
R78 VP.n55 VP.n7 15.9041
R79 VP.n66 VP.n3 15.9041
R80 VP.n30 VP.n15 15.9041
R81 VP.n58 VP.n7 8.56395
R82 VP.n67 VP.n66 8.56395
R83 VP.n31 VP.n30 8.56395
R84 VP.n22 VP.n19 8.56395
R85 VP.n21 VP.n20 5.17456
R86 VP.n47 VP.n11 1.22385
R87 VP.n79 VP.n78 1.22385
R88 VP.n43 VP.n42 1.22385
R89 VP.n44 VP.n12 0.278367
R90 VP.n46 VP.n45 0.278367
R91 VP.n80 VP.n0 0.278367
R92 VP.n21 VP.n18 0.189894
R93 VP.n25 VP.n18 0.189894
R94 VP.n26 VP.n25 0.189894
R95 VP.n27 VP.n26 0.189894
R96 VP.n27 VP.n16 0.189894
R97 VP.n32 VP.n16 0.189894
R98 VP.n33 VP.n32 0.189894
R99 VP.n34 VP.n33 0.189894
R100 VP.n34 VP.n14 0.189894
R101 VP.n38 VP.n14 0.189894
R102 VP.n39 VP.n38 0.189894
R103 VP.n40 VP.n39 0.189894
R104 VP.n40 VP.n12 0.189894
R105 VP.n46 VP.n10 0.189894
R106 VP.n50 VP.n10 0.189894
R107 VP.n51 VP.n50 0.189894
R108 VP.n52 VP.n51 0.189894
R109 VP.n52 VP.n8 0.189894
R110 VP.n56 VP.n8 0.189894
R111 VP.n57 VP.n56 0.189894
R112 VP.n57 VP.n6 0.189894
R113 VP.n61 VP.n6 0.189894
R114 VP.n62 VP.n61 0.189894
R115 VP.n63 VP.n62 0.189894
R116 VP.n63 VP.n4 0.189894
R117 VP.n68 VP.n4 0.189894
R118 VP.n69 VP.n68 0.189894
R119 VP.n70 VP.n69 0.189894
R120 VP.n70 VP.n2 0.189894
R121 VP.n74 VP.n2 0.189894
R122 VP.n75 VP.n74 0.189894
R123 VP.n76 VP.n75 0.189894
R124 VP.n76 VP.n0 0.189894
R125 VP VP.n80 0.153454
R126 VDD1 VDD1.n0 96.0333
R127 VDD1.n3 VDD1.n2 95.9187
R128 VDD1.n3 VDD1.n1 95.9187
R129 VDD1.n5 VDD1.n4 94.53
R130 VDD1.n5 VDD1.n3 42.2854
R131 VDD1.n4 VDD1.t5 5.61449
R132 VDD1.n4 VDD1.t6 5.61449
R133 VDD1.n0 VDD1.t1 5.61449
R134 VDD1.n0 VDD1.t4 5.61449
R135 VDD1.n2 VDD1.t7 5.61449
R136 VDD1.n2 VDD1.t3 5.61449
R137 VDD1.n1 VDD1.t0 5.61449
R138 VDD1.n1 VDD1.t2 5.61449
R139 VDD1 VDD1.n5 1.38628
R140 VTAIL.n246 VTAIL.n245 756.745
R141 VTAIL.n30 VTAIL.n29 756.745
R142 VTAIL.n60 VTAIL.n59 756.745
R143 VTAIL.n92 VTAIL.n91 756.745
R144 VTAIL.n216 VTAIL.n215 756.745
R145 VTAIL.n184 VTAIL.n183 756.745
R146 VTAIL.n154 VTAIL.n153 756.745
R147 VTAIL.n122 VTAIL.n121 756.745
R148 VTAIL.n229 VTAIL.n228 585
R149 VTAIL.n231 VTAIL.n230 585
R150 VTAIL.n224 VTAIL.n223 585
R151 VTAIL.n237 VTAIL.n236 585
R152 VTAIL.n239 VTAIL.n238 585
R153 VTAIL.n220 VTAIL.n219 585
R154 VTAIL.n245 VTAIL.n244 585
R155 VTAIL.n13 VTAIL.n12 585
R156 VTAIL.n15 VTAIL.n14 585
R157 VTAIL.n8 VTAIL.n7 585
R158 VTAIL.n21 VTAIL.n20 585
R159 VTAIL.n23 VTAIL.n22 585
R160 VTAIL.n4 VTAIL.n3 585
R161 VTAIL.n29 VTAIL.n28 585
R162 VTAIL.n43 VTAIL.n42 585
R163 VTAIL.n45 VTAIL.n44 585
R164 VTAIL.n38 VTAIL.n37 585
R165 VTAIL.n51 VTAIL.n50 585
R166 VTAIL.n53 VTAIL.n52 585
R167 VTAIL.n34 VTAIL.n33 585
R168 VTAIL.n59 VTAIL.n58 585
R169 VTAIL.n75 VTAIL.n74 585
R170 VTAIL.n77 VTAIL.n76 585
R171 VTAIL.n70 VTAIL.n69 585
R172 VTAIL.n83 VTAIL.n82 585
R173 VTAIL.n85 VTAIL.n84 585
R174 VTAIL.n66 VTAIL.n65 585
R175 VTAIL.n91 VTAIL.n90 585
R176 VTAIL.n215 VTAIL.n214 585
R177 VTAIL.n190 VTAIL.n189 585
R178 VTAIL.n209 VTAIL.n208 585
R179 VTAIL.n207 VTAIL.n206 585
R180 VTAIL.n194 VTAIL.n193 585
R181 VTAIL.n201 VTAIL.n200 585
R182 VTAIL.n199 VTAIL.n198 585
R183 VTAIL.n183 VTAIL.n182 585
R184 VTAIL.n158 VTAIL.n157 585
R185 VTAIL.n177 VTAIL.n176 585
R186 VTAIL.n175 VTAIL.n174 585
R187 VTAIL.n162 VTAIL.n161 585
R188 VTAIL.n169 VTAIL.n168 585
R189 VTAIL.n167 VTAIL.n166 585
R190 VTAIL.n153 VTAIL.n152 585
R191 VTAIL.n128 VTAIL.n127 585
R192 VTAIL.n147 VTAIL.n146 585
R193 VTAIL.n145 VTAIL.n144 585
R194 VTAIL.n132 VTAIL.n131 585
R195 VTAIL.n139 VTAIL.n138 585
R196 VTAIL.n137 VTAIL.n136 585
R197 VTAIL.n121 VTAIL.n120 585
R198 VTAIL.n96 VTAIL.n95 585
R199 VTAIL.n115 VTAIL.n114 585
R200 VTAIL.n113 VTAIL.n112 585
R201 VTAIL.n100 VTAIL.n99 585
R202 VTAIL.n107 VTAIL.n106 585
R203 VTAIL.n105 VTAIL.n104 585
R204 VTAIL.n227 VTAIL.t1 329.175
R205 VTAIL.n11 VTAIL.t0 329.175
R206 VTAIL.n41 VTAIL.t9 329.175
R207 VTAIL.n73 VTAIL.t12 329.175
R208 VTAIL.n197 VTAIL.t11 329.175
R209 VTAIL.n165 VTAIL.t14 329.175
R210 VTAIL.n135 VTAIL.t2 329.175
R211 VTAIL.n103 VTAIL.t6 329.175
R212 VTAIL.n230 VTAIL.n229 171.744
R213 VTAIL.n230 VTAIL.n223 171.744
R214 VTAIL.n237 VTAIL.n223 171.744
R215 VTAIL.n238 VTAIL.n237 171.744
R216 VTAIL.n238 VTAIL.n219 171.744
R217 VTAIL.n245 VTAIL.n219 171.744
R218 VTAIL.n14 VTAIL.n13 171.744
R219 VTAIL.n14 VTAIL.n7 171.744
R220 VTAIL.n21 VTAIL.n7 171.744
R221 VTAIL.n22 VTAIL.n21 171.744
R222 VTAIL.n22 VTAIL.n3 171.744
R223 VTAIL.n29 VTAIL.n3 171.744
R224 VTAIL.n44 VTAIL.n43 171.744
R225 VTAIL.n44 VTAIL.n37 171.744
R226 VTAIL.n51 VTAIL.n37 171.744
R227 VTAIL.n52 VTAIL.n51 171.744
R228 VTAIL.n52 VTAIL.n33 171.744
R229 VTAIL.n59 VTAIL.n33 171.744
R230 VTAIL.n76 VTAIL.n75 171.744
R231 VTAIL.n76 VTAIL.n69 171.744
R232 VTAIL.n83 VTAIL.n69 171.744
R233 VTAIL.n84 VTAIL.n83 171.744
R234 VTAIL.n84 VTAIL.n65 171.744
R235 VTAIL.n91 VTAIL.n65 171.744
R236 VTAIL.n215 VTAIL.n189 171.744
R237 VTAIL.n208 VTAIL.n189 171.744
R238 VTAIL.n208 VTAIL.n207 171.744
R239 VTAIL.n207 VTAIL.n193 171.744
R240 VTAIL.n200 VTAIL.n193 171.744
R241 VTAIL.n200 VTAIL.n199 171.744
R242 VTAIL.n183 VTAIL.n157 171.744
R243 VTAIL.n176 VTAIL.n157 171.744
R244 VTAIL.n176 VTAIL.n175 171.744
R245 VTAIL.n175 VTAIL.n161 171.744
R246 VTAIL.n168 VTAIL.n161 171.744
R247 VTAIL.n168 VTAIL.n167 171.744
R248 VTAIL.n153 VTAIL.n127 171.744
R249 VTAIL.n146 VTAIL.n127 171.744
R250 VTAIL.n146 VTAIL.n145 171.744
R251 VTAIL.n145 VTAIL.n131 171.744
R252 VTAIL.n138 VTAIL.n131 171.744
R253 VTAIL.n138 VTAIL.n137 171.744
R254 VTAIL.n121 VTAIL.n95 171.744
R255 VTAIL.n114 VTAIL.n95 171.744
R256 VTAIL.n114 VTAIL.n113 171.744
R257 VTAIL.n113 VTAIL.n99 171.744
R258 VTAIL.n106 VTAIL.n99 171.744
R259 VTAIL.n106 VTAIL.n105 171.744
R260 VTAIL.n229 VTAIL.t1 85.8723
R261 VTAIL.n13 VTAIL.t0 85.8723
R262 VTAIL.n43 VTAIL.t9 85.8723
R263 VTAIL.n75 VTAIL.t12 85.8723
R264 VTAIL.n199 VTAIL.t11 85.8723
R265 VTAIL.n167 VTAIL.t14 85.8723
R266 VTAIL.n137 VTAIL.t2 85.8723
R267 VTAIL.n105 VTAIL.t6 85.8723
R268 VTAIL.n187 VTAIL.n186 77.8523
R269 VTAIL.n125 VTAIL.n124 77.8523
R270 VTAIL.n1 VTAIL.n0 77.8513
R271 VTAIL.n63 VTAIL.n62 77.8513
R272 VTAIL.n247 VTAIL.n246 33.9308
R273 VTAIL.n31 VTAIL.n30 33.9308
R274 VTAIL.n61 VTAIL.n60 33.9308
R275 VTAIL.n93 VTAIL.n92 33.9308
R276 VTAIL.n217 VTAIL.n216 33.9308
R277 VTAIL.n185 VTAIL.n184 33.9308
R278 VTAIL.n155 VTAIL.n154 33.9308
R279 VTAIL.n123 VTAIL.n122 33.9308
R280 VTAIL.n247 VTAIL.n217 20.2462
R281 VTAIL.n123 VTAIL.n93 20.2462
R282 VTAIL.n244 VTAIL.n218 12.0247
R283 VTAIL.n28 VTAIL.n2 12.0247
R284 VTAIL.n58 VTAIL.n32 12.0247
R285 VTAIL.n90 VTAIL.n64 12.0247
R286 VTAIL.n214 VTAIL.n188 12.0247
R287 VTAIL.n182 VTAIL.n156 12.0247
R288 VTAIL.n152 VTAIL.n126 12.0247
R289 VTAIL.n120 VTAIL.n94 12.0247
R290 VTAIL.n243 VTAIL.n220 11.249
R291 VTAIL.n27 VTAIL.n4 11.249
R292 VTAIL.n57 VTAIL.n34 11.249
R293 VTAIL.n89 VTAIL.n66 11.249
R294 VTAIL.n213 VTAIL.n190 11.249
R295 VTAIL.n181 VTAIL.n158 11.249
R296 VTAIL.n151 VTAIL.n128 11.249
R297 VTAIL.n119 VTAIL.n96 11.249
R298 VTAIL.n228 VTAIL.n227 10.722
R299 VTAIL.n12 VTAIL.n11 10.722
R300 VTAIL.n42 VTAIL.n41 10.722
R301 VTAIL.n74 VTAIL.n73 10.722
R302 VTAIL.n198 VTAIL.n197 10.722
R303 VTAIL.n166 VTAIL.n165 10.722
R304 VTAIL.n136 VTAIL.n135 10.722
R305 VTAIL.n104 VTAIL.n103 10.722
R306 VTAIL.n240 VTAIL.n239 10.4732
R307 VTAIL.n24 VTAIL.n23 10.4732
R308 VTAIL.n54 VTAIL.n53 10.4732
R309 VTAIL.n86 VTAIL.n85 10.4732
R310 VTAIL.n210 VTAIL.n209 10.4732
R311 VTAIL.n178 VTAIL.n177 10.4732
R312 VTAIL.n148 VTAIL.n147 10.4732
R313 VTAIL.n116 VTAIL.n115 10.4732
R314 VTAIL.n236 VTAIL.n222 9.69747
R315 VTAIL.n20 VTAIL.n6 9.69747
R316 VTAIL.n50 VTAIL.n36 9.69747
R317 VTAIL.n82 VTAIL.n68 9.69747
R318 VTAIL.n206 VTAIL.n192 9.69747
R319 VTAIL.n174 VTAIL.n160 9.69747
R320 VTAIL.n144 VTAIL.n130 9.69747
R321 VTAIL.n112 VTAIL.n98 9.69747
R322 VTAIL.n242 VTAIL.n218 9.45567
R323 VTAIL.n26 VTAIL.n2 9.45567
R324 VTAIL.n56 VTAIL.n32 9.45567
R325 VTAIL.n88 VTAIL.n64 9.45567
R326 VTAIL.n212 VTAIL.n188 9.45567
R327 VTAIL.n180 VTAIL.n156 9.45567
R328 VTAIL.n150 VTAIL.n126 9.45567
R329 VTAIL.n118 VTAIL.n94 9.45567
R330 VTAIL.n226 VTAIL.n225 9.3005
R331 VTAIL.n233 VTAIL.n232 9.3005
R332 VTAIL.n235 VTAIL.n234 9.3005
R333 VTAIL.n222 VTAIL.n221 9.3005
R334 VTAIL.n241 VTAIL.n240 9.3005
R335 VTAIL.n243 VTAIL.n242 9.3005
R336 VTAIL.n10 VTAIL.n9 9.3005
R337 VTAIL.n17 VTAIL.n16 9.3005
R338 VTAIL.n19 VTAIL.n18 9.3005
R339 VTAIL.n6 VTAIL.n5 9.3005
R340 VTAIL.n25 VTAIL.n24 9.3005
R341 VTAIL.n27 VTAIL.n26 9.3005
R342 VTAIL.n40 VTAIL.n39 9.3005
R343 VTAIL.n47 VTAIL.n46 9.3005
R344 VTAIL.n49 VTAIL.n48 9.3005
R345 VTAIL.n36 VTAIL.n35 9.3005
R346 VTAIL.n55 VTAIL.n54 9.3005
R347 VTAIL.n57 VTAIL.n56 9.3005
R348 VTAIL.n72 VTAIL.n71 9.3005
R349 VTAIL.n79 VTAIL.n78 9.3005
R350 VTAIL.n81 VTAIL.n80 9.3005
R351 VTAIL.n68 VTAIL.n67 9.3005
R352 VTAIL.n87 VTAIL.n86 9.3005
R353 VTAIL.n89 VTAIL.n88 9.3005
R354 VTAIL.n213 VTAIL.n212 9.3005
R355 VTAIL.n211 VTAIL.n210 9.3005
R356 VTAIL.n192 VTAIL.n191 9.3005
R357 VTAIL.n205 VTAIL.n204 9.3005
R358 VTAIL.n203 VTAIL.n202 9.3005
R359 VTAIL.n196 VTAIL.n195 9.3005
R360 VTAIL.n171 VTAIL.n170 9.3005
R361 VTAIL.n173 VTAIL.n172 9.3005
R362 VTAIL.n160 VTAIL.n159 9.3005
R363 VTAIL.n179 VTAIL.n178 9.3005
R364 VTAIL.n181 VTAIL.n180 9.3005
R365 VTAIL.n164 VTAIL.n163 9.3005
R366 VTAIL.n141 VTAIL.n140 9.3005
R367 VTAIL.n143 VTAIL.n142 9.3005
R368 VTAIL.n130 VTAIL.n129 9.3005
R369 VTAIL.n149 VTAIL.n148 9.3005
R370 VTAIL.n151 VTAIL.n150 9.3005
R371 VTAIL.n134 VTAIL.n133 9.3005
R372 VTAIL.n109 VTAIL.n108 9.3005
R373 VTAIL.n111 VTAIL.n110 9.3005
R374 VTAIL.n98 VTAIL.n97 9.3005
R375 VTAIL.n117 VTAIL.n116 9.3005
R376 VTAIL.n119 VTAIL.n118 9.3005
R377 VTAIL.n102 VTAIL.n101 9.3005
R378 VTAIL.n235 VTAIL.n224 8.92171
R379 VTAIL.n19 VTAIL.n8 8.92171
R380 VTAIL.n49 VTAIL.n38 8.92171
R381 VTAIL.n81 VTAIL.n70 8.92171
R382 VTAIL.n205 VTAIL.n194 8.92171
R383 VTAIL.n173 VTAIL.n162 8.92171
R384 VTAIL.n143 VTAIL.n132 8.92171
R385 VTAIL.n111 VTAIL.n100 8.92171
R386 VTAIL.n232 VTAIL.n231 8.14595
R387 VTAIL.n16 VTAIL.n15 8.14595
R388 VTAIL.n46 VTAIL.n45 8.14595
R389 VTAIL.n78 VTAIL.n77 8.14595
R390 VTAIL.n202 VTAIL.n201 8.14595
R391 VTAIL.n170 VTAIL.n169 8.14595
R392 VTAIL.n140 VTAIL.n139 8.14595
R393 VTAIL.n108 VTAIL.n107 8.14595
R394 VTAIL.n228 VTAIL.n226 7.3702
R395 VTAIL.n12 VTAIL.n10 7.3702
R396 VTAIL.n42 VTAIL.n40 7.3702
R397 VTAIL.n74 VTAIL.n72 7.3702
R398 VTAIL.n198 VTAIL.n196 7.3702
R399 VTAIL.n166 VTAIL.n164 7.3702
R400 VTAIL.n136 VTAIL.n134 7.3702
R401 VTAIL.n104 VTAIL.n102 7.3702
R402 VTAIL.n231 VTAIL.n226 5.81868
R403 VTAIL.n15 VTAIL.n10 5.81868
R404 VTAIL.n45 VTAIL.n40 5.81868
R405 VTAIL.n77 VTAIL.n72 5.81868
R406 VTAIL.n201 VTAIL.n196 5.81868
R407 VTAIL.n169 VTAIL.n164 5.81868
R408 VTAIL.n139 VTAIL.n134 5.81868
R409 VTAIL.n107 VTAIL.n102 5.81868
R410 VTAIL.n0 VTAIL.t3 5.61449
R411 VTAIL.n0 VTAIL.t5 5.61449
R412 VTAIL.n62 VTAIL.t13 5.61449
R413 VTAIL.n62 VTAIL.t8 5.61449
R414 VTAIL.n186 VTAIL.t10 5.61449
R415 VTAIL.n186 VTAIL.t15 5.61449
R416 VTAIL.n124 VTAIL.t4 5.61449
R417 VTAIL.n124 VTAIL.t7 5.61449
R418 VTAIL.n232 VTAIL.n224 5.04292
R419 VTAIL.n16 VTAIL.n8 5.04292
R420 VTAIL.n46 VTAIL.n38 5.04292
R421 VTAIL.n78 VTAIL.n70 5.04292
R422 VTAIL.n202 VTAIL.n194 5.04292
R423 VTAIL.n170 VTAIL.n162 5.04292
R424 VTAIL.n140 VTAIL.n132 5.04292
R425 VTAIL.n108 VTAIL.n100 5.04292
R426 VTAIL.n236 VTAIL.n235 4.26717
R427 VTAIL.n20 VTAIL.n19 4.26717
R428 VTAIL.n50 VTAIL.n49 4.26717
R429 VTAIL.n82 VTAIL.n81 4.26717
R430 VTAIL.n206 VTAIL.n205 4.26717
R431 VTAIL.n174 VTAIL.n173 4.26717
R432 VTAIL.n144 VTAIL.n143 4.26717
R433 VTAIL.n112 VTAIL.n111 4.26717
R434 VTAIL.n239 VTAIL.n222 3.49141
R435 VTAIL.n23 VTAIL.n6 3.49141
R436 VTAIL.n53 VTAIL.n36 3.49141
R437 VTAIL.n85 VTAIL.n68 3.49141
R438 VTAIL.n209 VTAIL.n192 3.49141
R439 VTAIL.n177 VTAIL.n160 3.49141
R440 VTAIL.n147 VTAIL.n130 3.49141
R441 VTAIL.n115 VTAIL.n98 3.49141
R442 VTAIL.n125 VTAIL.n123 2.88843
R443 VTAIL.n155 VTAIL.n125 2.88843
R444 VTAIL.n187 VTAIL.n185 2.88843
R445 VTAIL.n217 VTAIL.n187 2.88843
R446 VTAIL.n93 VTAIL.n63 2.88843
R447 VTAIL.n63 VTAIL.n61 2.88843
R448 VTAIL.n31 VTAIL.n1 2.88843
R449 VTAIL VTAIL.n247 2.83024
R450 VTAIL.n240 VTAIL.n220 2.71565
R451 VTAIL.n24 VTAIL.n4 2.71565
R452 VTAIL.n54 VTAIL.n34 2.71565
R453 VTAIL.n86 VTAIL.n66 2.71565
R454 VTAIL.n210 VTAIL.n190 2.71565
R455 VTAIL.n178 VTAIL.n158 2.71565
R456 VTAIL.n148 VTAIL.n128 2.71565
R457 VTAIL.n116 VTAIL.n96 2.71565
R458 VTAIL.n227 VTAIL.n225 2.4147
R459 VTAIL.n11 VTAIL.n9 2.4147
R460 VTAIL.n41 VTAIL.n39 2.4147
R461 VTAIL.n73 VTAIL.n71 2.4147
R462 VTAIL.n197 VTAIL.n195 2.4147
R463 VTAIL.n165 VTAIL.n163 2.4147
R464 VTAIL.n135 VTAIL.n133 2.4147
R465 VTAIL.n103 VTAIL.n101 2.4147
R466 VTAIL.n244 VTAIL.n243 1.93989
R467 VTAIL.n28 VTAIL.n27 1.93989
R468 VTAIL.n58 VTAIL.n57 1.93989
R469 VTAIL.n90 VTAIL.n89 1.93989
R470 VTAIL.n214 VTAIL.n213 1.93989
R471 VTAIL.n182 VTAIL.n181 1.93989
R472 VTAIL.n152 VTAIL.n151 1.93989
R473 VTAIL.n120 VTAIL.n119 1.93989
R474 VTAIL.n246 VTAIL.n218 1.16414
R475 VTAIL.n30 VTAIL.n2 1.16414
R476 VTAIL.n60 VTAIL.n32 1.16414
R477 VTAIL.n92 VTAIL.n64 1.16414
R478 VTAIL.n216 VTAIL.n188 1.16414
R479 VTAIL.n184 VTAIL.n156 1.16414
R480 VTAIL.n154 VTAIL.n126 1.16414
R481 VTAIL.n122 VTAIL.n94 1.16414
R482 VTAIL.n185 VTAIL.n155 0.470328
R483 VTAIL.n61 VTAIL.n31 0.470328
R484 VTAIL.n233 VTAIL.n225 0.155672
R485 VTAIL.n234 VTAIL.n233 0.155672
R486 VTAIL.n234 VTAIL.n221 0.155672
R487 VTAIL.n241 VTAIL.n221 0.155672
R488 VTAIL.n242 VTAIL.n241 0.155672
R489 VTAIL.n17 VTAIL.n9 0.155672
R490 VTAIL.n18 VTAIL.n17 0.155672
R491 VTAIL.n18 VTAIL.n5 0.155672
R492 VTAIL.n25 VTAIL.n5 0.155672
R493 VTAIL.n26 VTAIL.n25 0.155672
R494 VTAIL.n47 VTAIL.n39 0.155672
R495 VTAIL.n48 VTAIL.n47 0.155672
R496 VTAIL.n48 VTAIL.n35 0.155672
R497 VTAIL.n55 VTAIL.n35 0.155672
R498 VTAIL.n56 VTAIL.n55 0.155672
R499 VTAIL.n79 VTAIL.n71 0.155672
R500 VTAIL.n80 VTAIL.n79 0.155672
R501 VTAIL.n80 VTAIL.n67 0.155672
R502 VTAIL.n87 VTAIL.n67 0.155672
R503 VTAIL.n88 VTAIL.n87 0.155672
R504 VTAIL.n212 VTAIL.n211 0.155672
R505 VTAIL.n211 VTAIL.n191 0.155672
R506 VTAIL.n204 VTAIL.n191 0.155672
R507 VTAIL.n204 VTAIL.n203 0.155672
R508 VTAIL.n203 VTAIL.n195 0.155672
R509 VTAIL.n180 VTAIL.n179 0.155672
R510 VTAIL.n179 VTAIL.n159 0.155672
R511 VTAIL.n172 VTAIL.n159 0.155672
R512 VTAIL.n172 VTAIL.n171 0.155672
R513 VTAIL.n171 VTAIL.n163 0.155672
R514 VTAIL.n150 VTAIL.n149 0.155672
R515 VTAIL.n149 VTAIL.n129 0.155672
R516 VTAIL.n142 VTAIL.n129 0.155672
R517 VTAIL.n142 VTAIL.n141 0.155672
R518 VTAIL.n141 VTAIL.n133 0.155672
R519 VTAIL.n118 VTAIL.n117 0.155672
R520 VTAIL.n117 VTAIL.n97 0.155672
R521 VTAIL.n110 VTAIL.n97 0.155672
R522 VTAIL.n110 VTAIL.n109 0.155672
R523 VTAIL.n109 VTAIL.n101 0.155672
R524 VTAIL VTAIL.n1 0.0586897
R525 VN.n63 VN.n33 161.3
R526 VN.n62 VN.n61 161.3
R527 VN.n60 VN.n34 161.3
R528 VN.n59 VN.n58 161.3
R529 VN.n57 VN.n35 161.3
R530 VN.n56 VN.n55 161.3
R531 VN.n54 VN.n36 161.3
R532 VN.n53 VN.n52 161.3
R533 VN.n51 VN.n37 161.3
R534 VN.n50 VN.n49 161.3
R535 VN.n48 VN.n39 161.3
R536 VN.n47 VN.n46 161.3
R537 VN.n45 VN.n40 161.3
R538 VN.n44 VN.n43 161.3
R539 VN.n30 VN.n0 161.3
R540 VN.n29 VN.n28 161.3
R541 VN.n27 VN.n1 161.3
R542 VN.n26 VN.n25 161.3
R543 VN.n24 VN.n2 161.3
R544 VN.n23 VN.n22 161.3
R545 VN.n21 VN.n3 161.3
R546 VN.n20 VN.n19 161.3
R547 VN.n17 VN.n4 161.3
R548 VN.n16 VN.n15 161.3
R549 VN.n14 VN.n5 161.3
R550 VN.n13 VN.n12 161.3
R551 VN.n11 VN.n6 161.3
R552 VN.n10 VN.n9 161.3
R553 VN.n32 VN.n31 109.534
R554 VN.n65 VN.n64 109.534
R555 VN.n8 VN.t5 78.4735
R556 VN.n42 VN.t4 78.4735
R557 VN.n8 VN.n7 65.4202
R558 VN.n42 VN.n41 65.4202
R559 VN.n25 VN.n24 55.0624
R560 VN.n58 VN.n57 55.0624
R561 VN VN.n65 48.4224
R562 VN.n7 VN.t6 46.2055
R563 VN.n18 VN.t2 46.2055
R564 VN.n31 VN.t3 46.2055
R565 VN.n41 VN.t1 46.2055
R566 VN.n38 VN.t7 46.2055
R567 VN.n64 VN.t0 46.2055
R568 VN.n12 VN.n5 40.4934
R569 VN.n16 VN.n5 40.4934
R570 VN.n46 VN.n39 40.4934
R571 VN.n50 VN.n39 40.4934
R572 VN.n25 VN.n1 25.9244
R573 VN.n58 VN.n34 25.9244
R574 VN.n11 VN.n10 24.4675
R575 VN.n12 VN.n11 24.4675
R576 VN.n17 VN.n16 24.4675
R577 VN.n19 VN.n17 24.4675
R578 VN.n23 VN.n3 24.4675
R579 VN.n24 VN.n23 24.4675
R580 VN.n29 VN.n1 24.4675
R581 VN.n30 VN.n29 24.4675
R582 VN.n46 VN.n45 24.4675
R583 VN.n45 VN.n44 24.4675
R584 VN.n57 VN.n56 24.4675
R585 VN.n56 VN.n36 24.4675
R586 VN.n52 VN.n51 24.4675
R587 VN.n51 VN.n50 24.4675
R588 VN.n63 VN.n62 24.4675
R589 VN.n62 VN.n34 24.4675
R590 VN.n18 VN.n3 15.9041
R591 VN.n38 VN.n36 15.9041
R592 VN.n10 VN.n7 8.56395
R593 VN.n19 VN.n18 8.56395
R594 VN.n44 VN.n41 8.56395
R595 VN.n52 VN.n38 8.56395
R596 VN.n43 VN.n42 5.17456
R597 VN.n9 VN.n8 5.17456
R598 VN.n31 VN.n30 1.22385
R599 VN.n64 VN.n63 1.22385
R600 VN.n65 VN.n33 0.278367
R601 VN.n32 VN.n0 0.278367
R602 VN.n61 VN.n33 0.189894
R603 VN.n61 VN.n60 0.189894
R604 VN.n60 VN.n59 0.189894
R605 VN.n59 VN.n35 0.189894
R606 VN.n55 VN.n35 0.189894
R607 VN.n55 VN.n54 0.189894
R608 VN.n54 VN.n53 0.189894
R609 VN.n53 VN.n37 0.189894
R610 VN.n49 VN.n37 0.189894
R611 VN.n49 VN.n48 0.189894
R612 VN.n48 VN.n47 0.189894
R613 VN.n47 VN.n40 0.189894
R614 VN.n43 VN.n40 0.189894
R615 VN.n9 VN.n6 0.189894
R616 VN.n13 VN.n6 0.189894
R617 VN.n14 VN.n13 0.189894
R618 VN.n15 VN.n14 0.189894
R619 VN.n15 VN.n4 0.189894
R620 VN.n20 VN.n4 0.189894
R621 VN.n21 VN.n20 0.189894
R622 VN.n22 VN.n21 0.189894
R623 VN.n22 VN.n2 0.189894
R624 VN.n26 VN.n2 0.189894
R625 VN.n27 VN.n26 0.189894
R626 VN.n28 VN.n27 0.189894
R627 VN.n28 VN.n0 0.189894
R628 VN VN.n32 0.153454
R629 VDD2.n2 VDD2.n1 95.9187
R630 VDD2.n2 VDD2.n0 95.9187
R631 VDD2 VDD2.n5 95.9157
R632 VDD2.n4 VDD2.n3 94.5311
R633 VDD2.n4 VDD2.n2 41.7024
R634 VDD2.n5 VDD2.t6 5.61449
R635 VDD2.n5 VDD2.t3 5.61449
R636 VDD2.n3 VDD2.t7 5.61449
R637 VDD2.n3 VDD2.t0 5.61449
R638 VDD2.n1 VDD2.t5 5.61449
R639 VDD2.n1 VDD2.t4 5.61449
R640 VDD2.n0 VDD2.t2 5.61449
R641 VDD2.n0 VDD2.t1 5.61449
R642 VDD2 VDD2.n4 1.50266
R643 B.n350 B.n121 585
R644 B.n349 B.n348 585
R645 B.n347 B.n122 585
R646 B.n346 B.n345 585
R647 B.n344 B.n123 585
R648 B.n343 B.n342 585
R649 B.n341 B.n124 585
R650 B.n340 B.n339 585
R651 B.n338 B.n125 585
R652 B.n337 B.n336 585
R653 B.n335 B.n126 585
R654 B.n334 B.n333 585
R655 B.n332 B.n127 585
R656 B.n331 B.n330 585
R657 B.n329 B.n128 585
R658 B.n328 B.n327 585
R659 B.n326 B.n129 585
R660 B.n325 B.n324 585
R661 B.n323 B.n130 585
R662 B.n322 B.n321 585
R663 B.n320 B.n131 585
R664 B.n319 B.n318 585
R665 B.n317 B.n132 585
R666 B.n316 B.n315 585
R667 B.n311 B.n133 585
R668 B.n310 B.n309 585
R669 B.n308 B.n134 585
R670 B.n307 B.n306 585
R671 B.n305 B.n135 585
R672 B.n304 B.n303 585
R673 B.n302 B.n136 585
R674 B.n301 B.n300 585
R675 B.n299 B.n137 585
R676 B.n297 B.n296 585
R677 B.n295 B.n140 585
R678 B.n294 B.n293 585
R679 B.n292 B.n141 585
R680 B.n291 B.n290 585
R681 B.n289 B.n142 585
R682 B.n288 B.n287 585
R683 B.n286 B.n143 585
R684 B.n285 B.n284 585
R685 B.n283 B.n144 585
R686 B.n282 B.n281 585
R687 B.n280 B.n145 585
R688 B.n279 B.n278 585
R689 B.n277 B.n146 585
R690 B.n276 B.n275 585
R691 B.n274 B.n147 585
R692 B.n273 B.n272 585
R693 B.n271 B.n148 585
R694 B.n270 B.n269 585
R695 B.n268 B.n149 585
R696 B.n267 B.n266 585
R697 B.n265 B.n150 585
R698 B.n264 B.n263 585
R699 B.n352 B.n351 585
R700 B.n353 B.n120 585
R701 B.n355 B.n354 585
R702 B.n356 B.n119 585
R703 B.n358 B.n357 585
R704 B.n359 B.n118 585
R705 B.n361 B.n360 585
R706 B.n362 B.n117 585
R707 B.n364 B.n363 585
R708 B.n365 B.n116 585
R709 B.n367 B.n366 585
R710 B.n368 B.n115 585
R711 B.n370 B.n369 585
R712 B.n371 B.n114 585
R713 B.n373 B.n372 585
R714 B.n374 B.n113 585
R715 B.n376 B.n375 585
R716 B.n377 B.n112 585
R717 B.n379 B.n378 585
R718 B.n380 B.n111 585
R719 B.n382 B.n381 585
R720 B.n383 B.n110 585
R721 B.n385 B.n384 585
R722 B.n386 B.n109 585
R723 B.n388 B.n387 585
R724 B.n389 B.n108 585
R725 B.n391 B.n390 585
R726 B.n392 B.n107 585
R727 B.n394 B.n393 585
R728 B.n395 B.n106 585
R729 B.n397 B.n396 585
R730 B.n398 B.n105 585
R731 B.n400 B.n399 585
R732 B.n401 B.n104 585
R733 B.n403 B.n402 585
R734 B.n404 B.n103 585
R735 B.n406 B.n405 585
R736 B.n407 B.n102 585
R737 B.n409 B.n408 585
R738 B.n410 B.n101 585
R739 B.n412 B.n411 585
R740 B.n413 B.n100 585
R741 B.n415 B.n414 585
R742 B.n416 B.n99 585
R743 B.n418 B.n417 585
R744 B.n419 B.n98 585
R745 B.n421 B.n420 585
R746 B.n422 B.n97 585
R747 B.n424 B.n423 585
R748 B.n425 B.n96 585
R749 B.n427 B.n426 585
R750 B.n428 B.n95 585
R751 B.n430 B.n429 585
R752 B.n431 B.n94 585
R753 B.n433 B.n432 585
R754 B.n434 B.n93 585
R755 B.n436 B.n435 585
R756 B.n437 B.n92 585
R757 B.n439 B.n438 585
R758 B.n440 B.n91 585
R759 B.n442 B.n441 585
R760 B.n443 B.n90 585
R761 B.n445 B.n444 585
R762 B.n446 B.n89 585
R763 B.n448 B.n447 585
R764 B.n449 B.n88 585
R765 B.n451 B.n450 585
R766 B.n452 B.n87 585
R767 B.n454 B.n453 585
R768 B.n455 B.n86 585
R769 B.n457 B.n456 585
R770 B.n458 B.n85 585
R771 B.n460 B.n459 585
R772 B.n461 B.n84 585
R773 B.n463 B.n462 585
R774 B.n464 B.n83 585
R775 B.n466 B.n465 585
R776 B.n467 B.n82 585
R777 B.n469 B.n468 585
R778 B.n470 B.n81 585
R779 B.n472 B.n471 585
R780 B.n473 B.n80 585
R781 B.n475 B.n474 585
R782 B.n476 B.n79 585
R783 B.n478 B.n477 585
R784 B.n479 B.n78 585
R785 B.n481 B.n480 585
R786 B.n482 B.n77 585
R787 B.n484 B.n483 585
R788 B.n485 B.n76 585
R789 B.n487 B.n486 585
R790 B.n488 B.n75 585
R791 B.n490 B.n489 585
R792 B.n491 B.n74 585
R793 B.n493 B.n492 585
R794 B.n494 B.n73 585
R795 B.n496 B.n495 585
R796 B.n497 B.n72 585
R797 B.n499 B.n498 585
R798 B.n500 B.n71 585
R799 B.n502 B.n501 585
R800 B.n503 B.n70 585
R801 B.n505 B.n504 585
R802 B.n506 B.n69 585
R803 B.n508 B.n507 585
R804 B.n509 B.n68 585
R805 B.n511 B.n510 585
R806 B.n512 B.n67 585
R807 B.n514 B.n513 585
R808 B.n515 B.n66 585
R809 B.n517 B.n516 585
R810 B.n518 B.n65 585
R811 B.n520 B.n519 585
R812 B.n521 B.n64 585
R813 B.n523 B.n522 585
R814 B.n524 B.n63 585
R815 B.n610 B.n609 585
R816 B.n608 B.n31 585
R817 B.n607 B.n606 585
R818 B.n605 B.n32 585
R819 B.n604 B.n603 585
R820 B.n602 B.n33 585
R821 B.n601 B.n600 585
R822 B.n599 B.n34 585
R823 B.n598 B.n597 585
R824 B.n596 B.n35 585
R825 B.n595 B.n594 585
R826 B.n593 B.n36 585
R827 B.n592 B.n591 585
R828 B.n590 B.n37 585
R829 B.n589 B.n588 585
R830 B.n587 B.n38 585
R831 B.n586 B.n585 585
R832 B.n584 B.n39 585
R833 B.n583 B.n582 585
R834 B.n581 B.n40 585
R835 B.n580 B.n579 585
R836 B.n578 B.n41 585
R837 B.n577 B.n576 585
R838 B.n575 B.n574 585
R839 B.n573 B.n45 585
R840 B.n572 B.n571 585
R841 B.n570 B.n46 585
R842 B.n569 B.n568 585
R843 B.n567 B.n47 585
R844 B.n566 B.n565 585
R845 B.n564 B.n48 585
R846 B.n563 B.n562 585
R847 B.n561 B.n49 585
R848 B.n559 B.n558 585
R849 B.n557 B.n52 585
R850 B.n556 B.n555 585
R851 B.n554 B.n53 585
R852 B.n553 B.n552 585
R853 B.n551 B.n54 585
R854 B.n550 B.n549 585
R855 B.n548 B.n55 585
R856 B.n547 B.n546 585
R857 B.n545 B.n56 585
R858 B.n544 B.n543 585
R859 B.n542 B.n57 585
R860 B.n541 B.n540 585
R861 B.n539 B.n58 585
R862 B.n538 B.n537 585
R863 B.n536 B.n59 585
R864 B.n535 B.n534 585
R865 B.n533 B.n60 585
R866 B.n532 B.n531 585
R867 B.n530 B.n61 585
R868 B.n529 B.n528 585
R869 B.n527 B.n62 585
R870 B.n526 B.n525 585
R871 B.n611 B.n30 585
R872 B.n613 B.n612 585
R873 B.n614 B.n29 585
R874 B.n616 B.n615 585
R875 B.n617 B.n28 585
R876 B.n619 B.n618 585
R877 B.n620 B.n27 585
R878 B.n622 B.n621 585
R879 B.n623 B.n26 585
R880 B.n625 B.n624 585
R881 B.n626 B.n25 585
R882 B.n628 B.n627 585
R883 B.n629 B.n24 585
R884 B.n631 B.n630 585
R885 B.n632 B.n23 585
R886 B.n634 B.n633 585
R887 B.n635 B.n22 585
R888 B.n637 B.n636 585
R889 B.n638 B.n21 585
R890 B.n640 B.n639 585
R891 B.n641 B.n20 585
R892 B.n643 B.n642 585
R893 B.n644 B.n19 585
R894 B.n646 B.n645 585
R895 B.n647 B.n18 585
R896 B.n649 B.n648 585
R897 B.n650 B.n17 585
R898 B.n652 B.n651 585
R899 B.n653 B.n16 585
R900 B.n655 B.n654 585
R901 B.n656 B.n15 585
R902 B.n658 B.n657 585
R903 B.n659 B.n14 585
R904 B.n661 B.n660 585
R905 B.n662 B.n13 585
R906 B.n664 B.n663 585
R907 B.n665 B.n12 585
R908 B.n667 B.n666 585
R909 B.n668 B.n11 585
R910 B.n670 B.n669 585
R911 B.n671 B.n10 585
R912 B.n673 B.n672 585
R913 B.n674 B.n9 585
R914 B.n676 B.n675 585
R915 B.n677 B.n8 585
R916 B.n679 B.n678 585
R917 B.n680 B.n7 585
R918 B.n682 B.n681 585
R919 B.n683 B.n6 585
R920 B.n685 B.n684 585
R921 B.n686 B.n5 585
R922 B.n688 B.n687 585
R923 B.n689 B.n4 585
R924 B.n691 B.n690 585
R925 B.n692 B.n3 585
R926 B.n694 B.n693 585
R927 B.n695 B.n0 585
R928 B.n2 B.n1 585
R929 B.n180 B.n179 585
R930 B.n181 B.n178 585
R931 B.n183 B.n182 585
R932 B.n184 B.n177 585
R933 B.n186 B.n185 585
R934 B.n187 B.n176 585
R935 B.n189 B.n188 585
R936 B.n190 B.n175 585
R937 B.n192 B.n191 585
R938 B.n193 B.n174 585
R939 B.n195 B.n194 585
R940 B.n196 B.n173 585
R941 B.n198 B.n197 585
R942 B.n199 B.n172 585
R943 B.n201 B.n200 585
R944 B.n202 B.n171 585
R945 B.n204 B.n203 585
R946 B.n205 B.n170 585
R947 B.n207 B.n206 585
R948 B.n208 B.n169 585
R949 B.n210 B.n209 585
R950 B.n211 B.n168 585
R951 B.n213 B.n212 585
R952 B.n214 B.n167 585
R953 B.n216 B.n215 585
R954 B.n217 B.n166 585
R955 B.n219 B.n218 585
R956 B.n220 B.n165 585
R957 B.n222 B.n221 585
R958 B.n223 B.n164 585
R959 B.n225 B.n224 585
R960 B.n226 B.n163 585
R961 B.n228 B.n227 585
R962 B.n229 B.n162 585
R963 B.n231 B.n230 585
R964 B.n232 B.n161 585
R965 B.n234 B.n233 585
R966 B.n235 B.n160 585
R967 B.n237 B.n236 585
R968 B.n238 B.n159 585
R969 B.n240 B.n239 585
R970 B.n241 B.n158 585
R971 B.n243 B.n242 585
R972 B.n244 B.n157 585
R973 B.n246 B.n245 585
R974 B.n247 B.n156 585
R975 B.n249 B.n248 585
R976 B.n250 B.n155 585
R977 B.n252 B.n251 585
R978 B.n253 B.n154 585
R979 B.n255 B.n254 585
R980 B.n256 B.n153 585
R981 B.n258 B.n257 585
R982 B.n259 B.n152 585
R983 B.n261 B.n260 585
R984 B.n262 B.n151 585
R985 B.n264 B.n151 502.111
R986 B.n352 B.n121 502.111
R987 B.n526 B.n63 502.111
R988 B.n611 B.n610 502.111
R989 B.n312 B.t10 329.089
R990 B.n50 B.t8 329.089
R991 B.n138 B.t4 329.089
R992 B.n42 B.t2 329.089
R993 B.n313 B.t11 264.12
R994 B.n51 B.t7 264.12
R995 B.n139 B.t5 264.12
R996 B.n43 B.t1 264.12
R997 B.n697 B.n696 256.663
R998 B.n138 B.t3 254.809
R999 B.n312 B.t9 254.809
R1000 B.n50 B.t6 254.809
R1001 B.n42 B.t0 254.809
R1002 B.n696 B.n695 235.042
R1003 B.n696 B.n2 235.042
R1004 B.n265 B.n264 163.367
R1005 B.n266 B.n265 163.367
R1006 B.n266 B.n149 163.367
R1007 B.n270 B.n149 163.367
R1008 B.n271 B.n270 163.367
R1009 B.n272 B.n271 163.367
R1010 B.n272 B.n147 163.367
R1011 B.n276 B.n147 163.367
R1012 B.n277 B.n276 163.367
R1013 B.n278 B.n277 163.367
R1014 B.n278 B.n145 163.367
R1015 B.n282 B.n145 163.367
R1016 B.n283 B.n282 163.367
R1017 B.n284 B.n283 163.367
R1018 B.n284 B.n143 163.367
R1019 B.n288 B.n143 163.367
R1020 B.n289 B.n288 163.367
R1021 B.n290 B.n289 163.367
R1022 B.n290 B.n141 163.367
R1023 B.n294 B.n141 163.367
R1024 B.n295 B.n294 163.367
R1025 B.n296 B.n295 163.367
R1026 B.n296 B.n137 163.367
R1027 B.n301 B.n137 163.367
R1028 B.n302 B.n301 163.367
R1029 B.n303 B.n302 163.367
R1030 B.n303 B.n135 163.367
R1031 B.n307 B.n135 163.367
R1032 B.n308 B.n307 163.367
R1033 B.n309 B.n308 163.367
R1034 B.n309 B.n133 163.367
R1035 B.n316 B.n133 163.367
R1036 B.n317 B.n316 163.367
R1037 B.n318 B.n317 163.367
R1038 B.n318 B.n131 163.367
R1039 B.n322 B.n131 163.367
R1040 B.n323 B.n322 163.367
R1041 B.n324 B.n323 163.367
R1042 B.n324 B.n129 163.367
R1043 B.n328 B.n129 163.367
R1044 B.n329 B.n328 163.367
R1045 B.n330 B.n329 163.367
R1046 B.n330 B.n127 163.367
R1047 B.n334 B.n127 163.367
R1048 B.n335 B.n334 163.367
R1049 B.n336 B.n335 163.367
R1050 B.n336 B.n125 163.367
R1051 B.n340 B.n125 163.367
R1052 B.n341 B.n340 163.367
R1053 B.n342 B.n341 163.367
R1054 B.n342 B.n123 163.367
R1055 B.n346 B.n123 163.367
R1056 B.n347 B.n346 163.367
R1057 B.n348 B.n347 163.367
R1058 B.n348 B.n121 163.367
R1059 B.n522 B.n63 163.367
R1060 B.n522 B.n521 163.367
R1061 B.n521 B.n520 163.367
R1062 B.n520 B.n65 163.367
R1063 B.n516 B.n65 163.367
R1064 B.n516 B.n515 163.367
R1065 B.n515 B.n514 163.367
R1066 B.n514 B.n67 163.367
R1067 B.n510 B.n67 163.367
R1068 B.n510 B.n509 163.367
R1069 B.n509 B.n508 163.367
R1070 B.n508 B.n69 163.367
R1071 B.n504 B.n69 163.367
R1072 B.n504 B.n503 163.367
R1073 B.n503 B.n502 163.367
R1074 B.n502 B.n71 163.367
R1075 B.n498 B.n71 163.367
R1076 B.n498 B.n497 163.367
R1077 B.n497 B.n496 163.367
R1078 B.n496 B.n73 163.367
R1079 B.n492 B.n73 163.367
R1080 B.n492 B.n491 163.367
R1081 B.n491 B.n490 163.367
R1082 B.n490 B.n75 163.367
R1083 B.n486 B.n75 163.367
R1084 B.n486 B.n485 163.367
R1085 B.n485 B.n484 163.367
R1086 B.n484 B.n77 163.367
R1087 B.n480 B.n77 163.367
R1088 B.n480 B.n479 163.367
R1089 B.n479 B.n478 163.367
R1090 B.n478 B.n79 163.367
R1091 B.n474 B.n79 163.367
R1092 B.n474 B.n473 163.367
R1093 B.n473 B.n472 163.367
R1094 B.n472 B.n81 163.367
R1095 B.n468 B.n81 163.367
R1096 B.n468 B.n467 163.367
R1097 B.n467 B.n466 163.367
R1098 B.n466 B.n83 163.367
R1099 B.n462 B.n83 163.367
R1100 B.n462 B.n461 163.367
R1101 B.n461 B.n460 163.367
R1102 B.n460 B.n85 163.367
R1103 B.n456 B.n85 163.367
R1104 B.n456 B.n455 163.367
R1105 B.n455 B.n454 163.367
R1106 B.n454 B.n87 163.367
R1107 B.n450 B.n87 163.367
R1108 B.n450 B.n449 163.367
R1109 B.n449 B.n448 163.367
R1110 B.n448 B.n89 163.367
R1111 B.n444 B.n89 163.367
R1112 B.n444 B.n443 163.367
R1113 B.n443 B.n442 163.367
R1114 B.n442 B.n91 163.367
R1115 B.n438 B.n91 163.367
R1116 B.n438 B.n437 163.367
R1117 B.n437 B.n436 163.367
R1118 B.n436 B.n93 163.367
R1119 B.n432 B.n93 163.367
R1120 B.n432 B.n431 163.367
R1121 B.n431 B.n430 163.367
R1122 B.n430 B.n95 163.367
R1123 B.n426 B.n95 163.367
R1124 B.n426 B.n425 163.367
R1125 B.n425 B.n424 163.367
R1126 B.n424 B.n97 163.367
R1127 B.n420 B.n97 163.367
R1128 B.n420 B.n419 163.367
R1129 B.n419 B.n418 163.367
R1130 B.n418 B.n99 163.367
R1131 B.n414 B.n99 163.367
R1132 B.n414 B.n413 163.367
R1133 B.n413 B.n412 163.367
R1134 B.n412 B.n101 163.367
R1135 B.n408 B.n101 163.367
R1136 B.n408 B.n407 163.367
R1137 B.n407 B.n406 163.367
R1138 B.n406 B.n103 163.367
R1139 B.n402 B.n103 163.367
R1140 B.n402 B.n401 163.367
R1141 B.n401 B.n400 163.367
R1142 B.n400 B.n105 163.367
R1143 B.n396 B.n105 163.367
R1144 B.n396 B.n395 163.367
R1145 B.n395 B.n394 163.367
R1146 B.n394 B.n107 163.367
R1147 B.n390 B.n107 163.367
R1148 B.n390 B.n389 163.367
R1149 B.n389 B.n388 163.367
R1150 B.n388 B.n109 163.367
R1151 B.n384 B.n109 163.367
R1152 B.n384 B.n383 163.367
R1153 B.n383 B.n382 163.367
R1154 B.n382 B.n111 163.367
R1155 B.n378 B.n111 163.367
R1156 B.n378 B.n377 163.367
R1157 B.n377 B.n376 163.367
R1158 B.n376 B.n113 163.367
R1159 B.n372 B.n113 163.367
R1160 B.n372 B.n371 163.367
R1161 B.n371 B.n370 163.367
R1162 B.n370 B.n115 163.367
R1163 B.n366 B.n115 163.367
R1164 B.n366 B.n365 163.367
R1165 B.n365 B.n364 163.367
R1166 B.n364 B.n117 163.367
R1167 B.n360 B.n117 163.367
R1168 B.n360 B.n359 163.367
R1169 B.n359 B.n358 163.367
R1170 B.n358 B.n119 163.367
R1171 B.n354 B.n119 163.367
R1172 B.n354 B.n353 163.367
R1173 B.n353 B.n352 163.367
R1174 B.n610 B.n31 163.367
R1175 B.n606 B.n31 163.367
R1176 B.n606 B.n605 163.367
R1177 B.n605 B.n604 163.367
R1178 B.n604 B.n33 163.367
R1179 B.n600 B.n33 163.367
R1180 B.n600 B.n599 163.367
R1181 B.n599 B.n598 163.367
R1182 B.n598 B.n35 163.367
R1183 B.n594 B.n35 163.367
R1184 B.n594 B.n593 163.367
R1185 B.n593 B.n592 163.367
R1186 B.n592 B.n37 163.367
R1187 B.n588 B.n37 163.367
R1188 B.n588 B.n587 163.367
R1189 B.n587 B.n586 163.367
R1190 B.n586 B.n39 163.367
R1191 B.n582 B.n39 163.367
R1192 B.n582 B.n581 163.367
R1193 B.n581 B.n580 163.367
R1194 B.n580 B.n41 163.367
R1195 B.n576 B.n41 163.367
R1196 B.n576 B.n575 163.367
R1197 B.n575 B.n45 163.367
R1198 B.n571 B.n45 163.367
R1199 B.n571 B.n570 163.367
R1200 B.n570 B.n569 163.367
R1201 B.n569 B.n47 163.367
R1202 B.n565 B.n47 163.367
R1203 B.n565 B.n564 163.367
R1204 B.n564 B.n563 163.367
R1205 B.n563 B.n49 163.367
R1206 B.n558 B.n49 163.367
R1207 B.n558 B.n557 163.367
R1208 B.n557 B.n556 163.367
R1209 B.n556 B.n53 163.367
R1210 B.n552 B.n53 163.367
R1211 B.n552 B.n551 163.367
R1212 B.n551 B.n550 163.367
R1213 B.n550 B.n55 163.367
R1214 B.n546 B.n55 163.367
R1215 B.n546 B.n545 163.367
R1216 B.n545 B.n544 163.367
R1217 B.n544 B.n57 163.367
R1218 B.n540 B.n57 163.367
R1219 B.n540 B.n539 163.367
R1220 B.n539 B.n538 163.367
R1221 B.n538 B.n59 163.367
R1222 B.n534 B.n59 163.367
R1223 B.n534 B.n533 163.367
R1224 B.n533 B.n532 163.367
R1225 B.n532 B.n61 163.367
R1226 B.n528 B.n61 163.367
R1227 B.n528 B.n527 163.367
R1228 B.n527 B.n526 163.367
R1229 B.n612 B.n611 163.367
R1230 B.n612 B.n29 163.367
R1231 B.n616 B.n29 163.367
R1232 B.n617 B.n616 163.367
R1233 B.n618 B.n617 163.367
R1234 B.n618 B.n27 163.367
R1235 B.n622 B.n27 163.367
R1236 B.n623 B.n622 163.367
R1237 B.n624 B.n623 163.367
R1238 B.n624 B.n25 163.367
R1239 B.n628 B.n25 163.367
R1240 B.n629 B.n628 163.367
R1241 B.n630 B.n629 163.367
R1242 B.n630 B.n23 163.367
R1243 B.n634 B.n23 163.367
R1244 B.n635 B.n634 163.367
R1245 B.n636 B.n635 163.367
R1246 B.n636 B.n21 163.367
R1247 B.n640 B.n21 163.367
R1248 B.n641 B.n640 163.367
R1249 B.n642 B.n641 163.367
R1250 B.n642 B.n19 163.367
R1251 B.n646 B.n19 163.367
R1252 B.n647 B.n646 163.367
R1253 B.n648 B.n647 163.367
R1254 B.n648 B.n17 163.367
R1255 B.n652 B.n17 163.367
R1256 B.n653 B.n652 163.367
R1257 B.n654 B.n653 163.367
R1258 B.n654 B.n15 163.367
R1259 B.n658 B.n15 163.367
R1260 B.n659 B.n658 163.367
R1261 B.n660 B.n659 163.367
R1262 B.n660 B.n13 163.367
R1263 B.n664 B.n13 163.367
R1264 B.n665 B.n664 163.367
R1265 B.n666 B.n665 163.367
R1266 B.n666 B.n11 163.367
R1267 B.n670 B.n11 163.367
R1268 B.n671 B.n670 163.367
R1269 B.n672 B.n671 163.367
R1270 B.n672 B.n9 163.367
R1271 B.n676 B.n9 163.367
R1272 B.n677 B.n676 163.367
R1273 B.n678 B.n677 163.367
R1274 B.n678 B.n7 163.367
R1275 B.n682 B.n7 163.367
R1276 B.n683 B.n682 163.367
R1277 B.n684 B.n683 163.367
R1278 B.n684 B.n5 163.367
R1279 B.n688 B.n5 163.367
R1280 B.n689 B.n688 163.367
R1281 B.n690 B.n689 163.367
R1282 B.n690 B.n3 163.367
R1283 B.n694 B.n3 163.367
R1284 B.n695 B.n694 163.367
R1285 B.n180 B.n2 163.367
R1286 B.n181 B.n180 163.367
R1287 B.n182 B.n181 163.367
R1288 B.n182 B.n177 163.367
R1289 B.n186 B.n177 163.367
R1290 B.n187 B.n186 163.367
R1291 B.n188 B.n187 163.367
R1292 B.n188 B.n175 163.367
R1293 B.n192 B.n175 163.367
R1294 B.n193 B.n192 163.367
R1295 B.n194 B.n193 163.367
R1296 B.n194 B.n173 163.367
R1297 B.n198 B.n173 163.367
R1298 B.n199 B.n198 163.367
R1299 B.n200 B.n199 163.367
R1300 B.n200 B.n171 163.367
R1301 B.n204 B.n171 163.367
R1302 B.n205 B.n204 163.367
R1303 B.n206 B.n205 163.367
R1304 B.n206 B.n169 163.367
R1305 B.n210 B.n169 163.367
R1306 B.n211 B.n210 163.367
R1307 B.n212 B.n211 163.367
R1308 B.n212 B.n167 163.367
R1309 B.n216 B.n167 163.367
R1310 B.n217 B.n216 163.367
R1311 B.n218 B.n217 163.367
R1312 B.n218 B.n165 163.367
R1313 B.n222 B.n165 163.367
R1314 B.n223 B.n222 163.367
R1315 B.n224 B.n223 163.367
R1316 B.n224 B.n163 163.367
R1317 B.n228 B.n163 163.367
R1318 B.n229 B.n228 163.367
R1319 B.n230 B.n229 163.367
R1320 B.n230 B.n161 163.367
R1321 B.n234 B.n161 163.367
R1322 B.n235 B.n234 163.367
R1323 B.n236 B.n235 163.367
R1324 B.n236 B.n159 163.367
R1325 B.n240 B.n159 163.367
R1326 B.n241 B.n240 163.367
R1327 B.n242 B.n241 163.367
R1328 B.n242 B.n157 163.367
R1329 B.n246 B.n157 163.367
R1330 B.n247 B.n246 163.367
R1331 B.n248 B.n247 163.367
R1332 B.n248 B.n155 163.367
R1333 B.n252 B.n155 163.367
R1334 B.n253 B.n252 163.367
R1335 B.n254 B.n253 163.367
R1336 B.n254 B.n153 163.367
R1337 B.n258 B.n153 163.367
R1338 B.n259 B.n258 163.367
R1339 B.n260 B.n259 163.367
R1340 B.n260 B.n151 163.367
R1341 B.n139 B.n138 64.9702
R1342 B.n313 B.n312 64.9702
R1343 B.n51 B.n50 64.9702
R1344 B.n43 B.n42 64.9702
R1345 B.n298 B.n139 59.5399
R1346 B.n314 B.n313 59.5399
R1347 B.n560 B.n51 59.5399
R1348 B.n44 B.n43 59.5399
R1349 B.n609 B.n30 32.6249
R1350 B.n525 B.n524 32.6249
R1351 B.n351 B.n350 32.6249
R1352 B.n263 B.n262 32.6249
R1353 B B.n697 18.0485
R1354 B.n613 B.n30 10.6151
R1355 B.n614 B.n613 10.6151
R1356 B.n615 B.n614 10.6151
R1357 B.n615 B.n28 10.6151
R1358 B.n619 B.n28 10.6151
R1359 B.n620 B.n619 10.6151
R1360 B.n621 B.n620 10.6151
R1361 B.n621 B.n26 10.6151
R1362 B.n625 B.n26 10.6151
R1363 B.n626 B.n625 10.6151
R1364 B.n627 B.n626 10.6151
R1365 B.n627 B.n24 10.6151
R1366 B.n631 B.n24 10.6151
R1367 B.n632 B.n631 10.6151
R1368 B.n633 B.n632 10.6151
R1369 B.n633 B.n22 10.6151
R1370 B.n637 B.n22 10.6151
R1371 B.n638 B.n637 10.6151
R1372 B.n639 B.n638 10.6151
R1373 B.n639 B.n20 10.6151
R1374 B.n643 B.n20 10.6151
R1375 B.n644 B.n643 10.6151
R1376 B.n645 B.n644 10.6151
R1377 B.n645 B.n18 10.6151
R1378 B.n649 B.n18 10.6151
R1379 B.n650 B.n649 10.6151
R1380 B.n651 B.n650 10.6151
R1381 B.n651 B.n16 10.6151
R1382 B.n655 B.n16 10.6151
R1383 B.n656 B.n655 10.6151
R1384 B.n657 B.n656 10.6151
R1385 B.n657 B.n14 10.6151
R1386 B.n661 B.n14 10.6151
R1387 B.n662 B.n661 10.6151
R1388 B.n663 B.n662 10.6151
R1389 B.n663 B.n12 10.6151
R1390 B.n667 B.n12 10.6151
R1391 B.n668 B.n667 10.6151
R1392 B.n669 B.n668 10.6151
R1393 B.n669 B.n10 10.6151
R1394 B.n673 B.n10 10.6151
R1395 B.n674 B.n673 10.6151
R1396 B.n675 B.n674 10.6151
R1397 B.n675 B.n8 10.6151
R1398 B.n679 B.n8 10.6151
R1399 B.n680 B.n679 10.6151
R1400 B.n681 B.n680 10.6151
R1401 B.n681 B.n6 10.6151
R1402 B.n685 B.n6 10.6151
R1403 B.n686 B.n685 10.6151
R1404 B.n687 B.n686 10.6151
R1405 B.n687 B.n4 10.6151
R1406 B.n691 B.n4 10.6151
R1407 B.n692 B.n691 10.6151
R1408 B.n693 B.n692 10.6151
R1409 B.n693 B.n0 10.6151
R1410 B.n609 B.n608 10.6151
R1411 B.n608 B.n607 10.6151
R1412 B.n607 B.n32 10.6151
R1413 B.n603 B.n32 10.6151
R1414 B.n603 B.n602 10.6151
R1415 B.n602 B.n601 10.6151
R1416 B.n601 B.n34 10.6151
R1417 B.n597 B.n34 10.6151
R1418 B.n597 B.n596 10.6151
R1419 B.n596 B.n595 10.6151
R1420 B.n595 B.n36 10.6151
R1421 B.n591 B.n36 10.6151
R1422 B.n591 B.n590 10.6151
R1423 B.n590 B.n589 10.6151
R1424 B.n589 B.n38 10.6151
R1425 B.n585 B.n38 10.6151
R1426 B.n585 B.n584 10.6151
R1427 B.n584 B.n583 10.6151
R1428 B.n583 B.n40 10.6151
R1429 B.n579 B.n40 10.6151
R1430 B.n579 B.n578 10.6151
R1431 B.n578 B.n577 10.6151
R1432 B.n574 B.n573 10.6151
R1433 B.n573 B.n572 10.6151
R1434 B.n572 B.n46 10.6151
R1435 B.n568 B.n46 10.6151
R1436 B.n568 B.n567 10.6151
R1437 B.n567 B.n566 10.6151
R1438 B.n566 B.n48 10.6151
R1439 B.n562 B.n48 10.6151
R1440 B.n562 B.n561 10.6151
R1441 B.n559 B.n52 10.6151
R1442 B.n555 B.n52 10.6151
R1443 B.n555 B.n554 10.6151
R1444 B.n554 B.n553 10.6151
R1445 B.n553 B.n54 10.6151
R1446 B.n549 B.n54 10.6151
R1447 B.n549 B.n548 10.6151
R1448 B.n548 B.n547 10.6151
R1449 B.n547 B.n56 10.6151
R1450 B.n543 B.n56 10.6151
R1451 B.n543 B.n542 10.6151
R1452 B.n542 B.n541 10.6151
R1453 B.n541 B.n58 10.6151
R1454 B.n537 B.n58 10.6151
R1455 B.n537 B.n536 10.6151
R1456 B.n536 B.n535 10.6151
R1457 B.n535 B.n60 10.6151
R1458 B.n531 B.n60 10.6151
R1459 B.n531 B.n530 10.6151
R1460 B.n530 B.n529 10.6151
R1461 B.n529 B.n62 10.6151
R1462 B.n525 B.n62 10.6151
R1463 B.n524 B.n523 10.6151
R1464 B.n523 B.n64 10.6151
R1465 B.n519 B.n64 10.6151
R1466 B.n519 B.n518 10.6151
R1467 B.n518 B.n517 10.6151
R1468 B.n517 B.n66 10.6151
R1469 B.n513 B.n66 10.6151
R1470 B.n513 B.n512 10.6151
R1471 B.n512 B.n511 10.6151
R1472 B.n511 B.n68 10.6151
R1473 B.n507 B.n68 10.6151
R1474 B.n507 B.n506 10.6151
R1475 B.n506 B.n505 10.6151
R1476 B.n505 B.n70 10.6151
R1477 B.n501 B.n70 10.6151
R1478 B.n501 B.n500 10.6151
R1479 B.n500 B.n499 10.6151
R1480 B.n499 B.n72 10.6151
R1481 B.n495 B.n72 10.6151
R1482 B.n495 B.n494 10.6151
R1483 B.n494 B.n493 10.6151
R1484 B.n493 B.n74 10.6151
R1485 B.n489 B.n74 10.6151
R1486 B.n489 B.n488 10.6151
R1487 B.n488 B.n487 10.6151
R1488 B.n487 B.n76 10.6151
R1489 B.n483 B.n76 10.6151
R1490 B.n483 B.n482 10.6151
R1491 B.n482 B.n481 10.6151
R1492 B.n481 B.n78 10.6151
R1493 B.n477 B.n78 10.6151
R1494 B.n477 B.n476 10.6151
R1495 B.n476 B.n475 10.6151
R1496 B.n475 B.n80 10.6151
R1497 B.n471 B.n80 10.6151
R1498 B.n471 B.n470 10.6151
R1499 B.n470 B.n469 10.6151
R1500 B.n469 B.n82 10.6151
R1501 B.n465 B.n82 10.6151
R1502 B.n465 B.n464 10.6151
R1503 B.n464 B.n463 10.6151
R1504 B.n463 B.n84 10.6151
R1505 B.n459 B.n84 10.6151
R1506 B.n459 B.n458 10.6151
R1507 B.n458 B.n457 10.6151
R1508 B.n457 B.n86 10.6151
R1509 B.n453 B.n86 10.6151
R1510 B.n453 B.n452 10.6151
R1511 B.n452 B.n451 10.6151
R1512 B.n451 B.n88 10.6151
R1513 B.n447 B.n88 10.6151
R1514 B.n447 B.n446 10.6151
R1515 B.n446 B.n445 10.6151
R1516 B.n445 B.n90 10.6151
R1517 B.n441 B.n90 10.6151
R1518 B.n441 B.n440 10.6151
R1519 B.n440 B.n439 10.6151
R1520 B.n439 B.n92 10.6151
R1521 B.n435 B.n92 10.6151
R1522 B.n435 B.n434 10.6151
R1523 B.n434 B.n433 10.6151
R1524 B.n433 B.n94 10.6151
R1525 B.n429 B.n94 10.6151
R1526 B.n429 B.n428 10.6151
R1527 B.n428 B.n427 10.6151
R1528 B.n427 B.n96 10.6151
R1529 B.n423 B.n96 10.6151
R1530 B.n423 B.n422 10.6151
R1531 B.n422 B.n421 10.6151
R1532 B.n421 B.n98 10.6151
R1533 B.n417 B.n98 10.6151
R1534 B.n417 B.n416 10.6151
R1535 B.n416 B.n415 10.6151
R1536 B.n415 B.n100 10.6151
R1537 B.n411 B.n100 10.6151
R1538 B.n411 B.n410 10.6151
R1539 B.n410 B.n409 10.6151
R1540 B.n409 B.n102 10.6151
R1541 B.n405 B.n102 10.6151
R1542 B.n405 B.n404 10.6151
R1543 B.n404 B.n403 10.6151
R1544 B.n403 B.n104 10.6151
R1545 B.n399 B.n104 10.6151
R1546 B.n399 B.n398 10.6151
R1547 B.n398 B.n397 10.6151
R1548 B.n397 B.n106 10.6151
R1549 B.n393 B.n106 10.6151
R1550 B.n393 B.n392 10.6151
R1551 B.n392 B.n391 10.6151
R1552 B.n391 B.n108 10.6151
R1553 B.n387 B.n108 10.6151
R1554 B.n387 B.n386 10.6151
R1555 B.n386 B.n385 10.6151
R1556 B.n385 B.n110 10.6151
R1557 B.n381 B.n110 10.6151
R1558 B.n381 B.n380 10.6151
R1559 B.n380 B.n379 10.6151
R1560 B.n379 B.n112 10.6151
R1561 B.n375 B.n112 10.6151
R1562 B.n375 B.n374 10.6151
R1563 B.n374 B.n373 10.6151
R1564 B.n373 B.n114 10.6151
R1565 B.n369 B.n114 10.6151
R1566 B.n369 B.n368 10.6151
R1567 B.n368 B.n367 10.6151
R1568 B.n367 B.n116 10.6151
R1569 B.n363 B.n116 10.6151
R1570 B.n363 B.n362 10.6151
R1571 B.n362 B.n361 10.6151
R1572 B.n361 B.n118 10.6151
R1573 B.n357 B.n118 10.6151
R1574 B.n357 B.n356 10.6151
R1575 B.n356 B.n355 10.6151
R1576 B.n355 B.n120 10.6151
R1577 B.n351 B.n120 10.6151
R1578 B.n179 B.n1 10.6151
R1579 B.n179 B.n178 10.6151
R1580 B.n183 B.n178 10.6151
R1581 B.n184 B.n183 10.6151
R1582 B.n185 B.n184 10.6151
R1583 B.n185 B.n176 10.6151
R1584 B.n189 B.n176 10.6151
R1585 B.n190 B.n189 10.6151
R1586 B.n191 B.n190 10.6151
R1587 B.n191 B.n174 10.6151
R1588 B.n195 B.n174 10.6151
R1589 B.n196 B.n195 10.6151
R1590 B.n197 B.n196 10.6151
R1591 B.n197 B.n172 10.6151
R1592 B.n201 B.n172 10.6151
R1593 B.n202 B.n201 10.6151
R1594 B.n203 B.n202 10.6151
R1595 B.n203 B.n170 10.6151
R1596 B.n207 B.n170 10.6151
R1597 B.n208 B.n207 10.6151
R1598 B.n209 B.n208 10.6151
R1599 B.n209 B.n168 10.6151
R1600 B.n213 B.n168 10.6151
R1601 B.n214 B.n213 10.6151
R1602 B.n215 B.n214 10.6151
R1603 B.n215 B.n166 10.6151
R1604 B.n219 B.n166 10.6151
R1605 B.n220 B.n219 10.6151
R1606 B.n221 B.n220 10.6151
R1607 B.n221 B.n164 10.6151
R1608 B.n225 B.n164 10.6151
R1609 B.n226 B.n225 10.6151
R1610 B.n227 B.n226 10.6151
R1611 B.n227 B.n162 10.6151
R1612 B.n231 B.n162 10.6151
R1613 B.n232 B.n231 10.6151
R1614 B.n233 B.n232 10.6151
R1615 B.n233 B.n160 10.6151
R1616 B.n237 B.n160 10.6151
R1617 B.n238 B.n237 10.6151
R1618 B.n239 B.n238 10.6151
R1619 B.n239 B.n158 10.6151
R1620 B.n243 B.n158 10.6151
R1621 B.n244 B.n243 10.6151
R1622 B.n245 B.n244 10.6151
R1623 B.n245 B.n156 10.6151
R1624 B.n249 B.n156 10.6151
R1625 B.n250 B.n249 10.6151
R1626 B.n251 B.n250 10.6151
R1627 B.n251 B.n154 10.6151
R1628 B.n255 B.n154 10.6151
R1629 B.n256 B.n255 10.6151
R1630 B.n257 B.n256 10.6151
R1631 B.n257 B.n152 10.6151
R1632 B.n261 B.n152 10.6151
R1633 B.n262 B.n261 10.6151
R1634 B.n263 B.n150 10.6151
R1635 B.n267 B.n150 10.6151
R1636 B.n268 B.n267 10.6151
R1637 B.n269 B.n268 10.6151
R1638 B.n269 B.n148 10.6151
R1639 B.n273 B.n148 10.6151
R1640 B.n274 B.n273 10.6151
R1641 B.n275 B.n274 10.6151
R1642 B.n275 B.n146 10.6151
R1643 B.n279 B.n146 10.6151
R1644 B.n280 B.n279 10.6151
R1645 B.n281 B.n280 10.6151
R1646 B.n281 B.n144 10.6151
R1647 B.n285 B.n144 10.6151
R1648 B.n286 B.n285 10.6151
R1649 B.n287 B.n286 10.6151
R1650 B.n287 B.n142 10.6151
R1651 B.n291 B.n142 10.6151
R1652 B.n292 B.n291 10.6151
R1653 B.n293 B.n292 10.6151
R1654 B.n293 B.n140 10.6151
R1655 B.n297 B.n140 10.6151
R1656 B.n300 B.n299 10.6151
R1657 B.n300 B.n136 10.6151
R1658 B.n304 B.n136 10.6151
R1659 B.n305 B.n304 10.6151
R1660 B.n306 B.n305 10.6151
R1661 B.n306 B.n134 10.6151
R1662 B.n310 B.n134 10.6151
R1663 B.n311 B.n310 10.6151
R1664 B.n315 B.n311 10.6151
R1665 B.n319 B.n132 10.6151
R1666 B.n320 B.n319 10.6151
R1667 B.n321 B.n320 10.6151
R1668 B.n321 B.n130 10.6151
R1669 B.n325 B.n130 10.6151
R1670 B.n326 B.n325 10.6151
R1671 B.n327 B.n326 10.6151
R1672 B.n327 B.n128 10.6151
R1673 B.n331 B.n128 10.6151
R1674 B.n332 B.n331 10.6151
R1675 B.n333 B.n332 10.6151
R1676 B.n333 B.n126 10.6151
R1677 B.n337 B.n126 10.6151
R1678 B.n338 B.n337 10.6151
R1679 B.n339 B.n338 10.6151
R1680 B.n339 B.n124 10.6151
R1681 B.n343 B.n124 10.6151
R1682 B.n344 B.n343 10.6151
R1683 B.n345 B.n344 10.6151
R1684 B.n345 B.n122 10.6151
R1685 B.n349 B.n122 10.6151
R1686 B.n350 B.n349 10.6151
R1687 B.n577 B.n44 9.36635
R1688 B.n560 B.n559 9.36635
R1689 B.n298 B.n297 9.36635
R1690 B.n314 B.n132 9.36635
R1691 B.n697 B.n0 8.11757
R1692 B.n697 B.n1 8.11757
R1693 B.n574 B.n44 1.24928
R1694 B.n561 B.n560 1.24928
R1695 B.n299 B.n298 1.24928
R1696 B.n315 B.n314 1.24928
C0 VDD2 VDD1 1.99652f
C1 B VTAIL 3.06891f
C2 B w_n4320_n2126# 9.03197f
C3 VDD1 VTAIL 6.27187f
C4 VP B 2.18826f
C5 VDD1 w_n4320_n2126# 1.92496f
C6 VN B 1.24381f
C7 VP VDD1 4.95898f
C8 VDD2 VTAIL 6.3291f
C9 VN VDD1 0.152537f
C10 VDD2 w_n4320_n2126# 2.05724f
C11 VP VDD2 0.564413f
C12 VTAIL w_n4320_n2126# 2.85588f
C13 VN VDD2 4.54872f
C14 VP VTAIL 5.59046f
C15 VP w_n4320_n2126# 9.358191f
C16 VDD1 B 1.60984f
C17 VN VTAIL 5.57636f
C18 VN w_n4320_n2126# 8.796121f
C19 VN VP 7.02431f
C20 VDD2 B 1.71917f
C21 VDD2 VSUBS 1.831995f
C22 VDD1 VSUBS 2.401f
C23 VTAIL VSUBS 0.737381f
C24 VN VSUBS 7.04158f
C25 VP VSUBS 3.570046f
C26 B VSUBS 4.949981f
C27 w_n4320_n2126# VSUBS 0.114722p
C28 B.n0 VSUBS 0.008368f
C29 B.n1 VSUBS 0.008368f
C30 B.n2 VSUBS 0.012376f
C31 B.n3 VSUBS 0.009484f
C32 B.n4 VSUBS 0.009484f
C33 B.n5 VSUBS 0.009484f
C34 B.n6 VSUBS 0.009484f
C35 B.n7 VSUBS 0.009484f
C36 B.n8 VSUBS 0.009484f
C37 B.n9 VSUBS 0.009484f
C38 B.n10 VSUBS 0.009484f
C39 B.n11 VSUBS 0.009484f
C40 B.n12 VSUBS 0.009484f
C41 B.n13 VSUBS 0.009484f
C42 B.n14 VSUBS 0.009484f
C43 B.n15 VSUBS 0.009484f
C44 B.n16 VSUBS 0.009484f
C45 B.n17 VSUBS 0.009484f
C46 B.n18 VSUBS 0.009484f
C47 B.n19 VSUBS 0.009484f
C48 B.n20 VSUBS 0.009484f
C49 B.n21 VSUBS 0.009484f
C50 B.n22 VSUBS 0.009484f
C51 B.n23 VSUBS 0.009484f
C52 B.n24 VSUBS 0.009484f
C53 B.n25 VSUBS 0.009484f
C54 B.n26 VSUBS 0.009484f
C55 B.n27 VSUBS 0.009484f
C56 B.n28 VSUBS 0.009484f
C57 B.n29 VSUBS 0.009484f
C58 B.n30 VSUBS 0.021888f
C59 B.n31 VSUBS 0.009484f
C60 B.n32 VSUBS 0.009484f
C61 B.n33 VSUBS 0.009484f
C62 B.n34 VSUBS 0.009484f
C63 B.n35 VSUBS 0.009484f
C64 B.n36 VSUBS 0.009484f
C65 B.n37 VSUBS 0.009484f
C66 B.n38 VSUBS 0.009484f
C67 B.n39 VSUBS 0.009484f
C68 B.n40 VSUBS 0.009484f
C69 B.n41 VSUBS 0.009484f
C70 B.t1 VSUBS 0.115748f
C71 B.t2 VSUBS 0.154439f
C72 B.t0 VSUBS 1.12996f
C73 B.n42 VSUBS 0.261924f
C74 B.n43 VSUBS 0.209506f
C75 B.n44 VSUBS 0.021972f
C76 B.n45 VSUBS 0.009484f
C77 B.n46 VSUBS 0.009484f
C78 B.n47 VSUBS 0.009484f
C79 B.n48 VSUBS 0.009484f
C80 B.n49 VSUBS 0.009484f
C81 B.t7 VSUBS 0.115751f
C82 B.t8 VSUBS 0.154441f
C83 B.t6 VSUBS 1.12996f
C84 B.n50 VSUBS 0.261922f
C85 B.n51 VSUBS 0.209504f
C86 B.n52 VSUBS 0.009484f
C87 B.n53 VSUBS 0.009484f
C88 B.n54 VSUBS 0.009484f
C89 B.n55 VSUBS 0.009484f
C90 B.n56 VSUBS 0.009484f
C91 B.n57 VSUBS 0.009484f
C92 B.n58 VSUBS 0.009484f
C93 B.n59 VSUBS 0.009484f
C94 B.n60 VSUBS 0.009484f
C95 B.n61 VSUBS 0.009484f
C96 B.n62 VSUBS 0.009484f
C97 B.n63 VSUBS 0.021888f
C98 B.n64 VSUBS 0.009484f
C99 B.n65 VSUBS 0.009484f
C100 B.n66 VSUBS 0.009484f
C101 B.n67 VSUBS 0.009484f
C102 B.n68 VSUBS 0.009484f
C103 B.n69 VSUBS 0.009484f
C104 B.n70 VSUBS 0.009484f
C105 B.n71 VSUBS 0.009484f
C106 B.n72 VSUBS 0.009484f
C107 B.n73 VSUBS 0.009484f
C108 B.n74 VSUBS 0.009484f
C109 B.n75 VSUBS 0.009484f
C110 B.n76 VSUBS 0.009484f
C111 B.n77 VSUBS 0.009484f
C112 B.n78 VSUBS 0.009484f
C113 B.n79 VSUBS 0.009484f
C114 B.n80 VSUBS 0.009484f
C115 B.n81 VSUBS 0.009484f
C116 B.n82 VSUBS 0.009484f
C117 B.n83 VSUBS 0.009484f
C118 B.n84 VSUBS 0.009484f
C119 B.n85 VSUBS 0.009484f
C120 B.n86 VSUBS 0.009484f
C121 B.n87 VSUBS 0.009484f
C122 B.n88 VSUBS 0.009484f
C123 B.n89 VSUBS 0.009484f
C124 B.n90 VSUBS 0.009484f
C125 B.n91 VSUBS 0.009484f
C126 B.n92 VSUBS 0.009484f
C127 B.n93 VSUBS 0.009484f
C128 B.n94 VSUBS 0.009484f
C129 B.n95 VSUBS 0.009484f
C130 B.n96 VSUBS 0.009484f
C131 B.n97 VSUBS 0.009484f
C132 B.n98 VSUBS 0.009484f
C133 B.n99 VSUBS 0.009484f
C134 B.n100 VSUBS 0.009484f
C135 B.n101 VSUBS 0.009484f
C136 B.n102 VSUBS 0.009484f
C137 B.n103 VSUBS 0.009484f
C138 B.n104 VSUBS 0.009484f
C139 B.n105 VSUBS 0.009484f
C140 B.n106 VSUBS 0.009484f
C141 B.n107 VSUBS 0.009484f
C142 B.n108 VSUBS 0.009484f
C143 B.n109 VSUBS 0.009484f
C144 B.n110 VSUBS 0.009484f
C145 B.n111 VSUBS 0.009484f
C146 B.n112 VSUBS 0.009484f
C147 B.n113 VSUBS 0.009484f
C148 B.n114 VSUBS 0.009484f
C149 B.n115 VSUBS 0.009484f
C150 B.n116 VSUBS 0.009484f
C151 B.n117 VSUBS 0.009484f
C152 B.n118 VSUBS 0.009484f
C153 B.n119 VSUBS 0.009484f
C154 B.n120 VSUBS 0.009484f
C155 B.n121 VSUBS 0.022462f
C156 B.n122 VSUBS 0.009484f
C157 B.n123 VSUBS 0.009484f
C158 B.n124 VSUBS 0.009484f
C159 B.n125 VSUBS 0.009484f
C160 B.n126 VSUBS 0.009484f
C161 B.n127 VSUBS 0.009484f
C162 B.n128 VSUBS 0.009484f
C163 B.n129 VSUBS 0.009484f
C164 B.n130 VSUBS 0.009484f
C165 B.n131 VSUBS 0.009484f
C166 B.n132 VSUBS 0.008926f
C167 B.n133 VSUBS 0.009484f
C168 B.n134 VSUBS 0.009484f
C169 B.n135 VSUBS 0.009484f
C170 B.n136 VSUBS 0.009484f
C171 B.n137 VSUBS 0.009484f
C172 B.t5 VSUBS 0.115748f
C173 B.t4 VSUBS 0.154439f
C174 B.t3 VSUBS 1.12996f
C175 B.n138 VSUBS 0.261924f
C176 B.n139 VSUBS 0.209506f
C177 B.n140 VSUBS 0.009484f
C178 B.n141 VSUBS 0.009484f
C179 B.n142 VSUBS 0.009484f
C180 B.n143 VSUBS 0.009484f
C181 B.n144 VSUBS 0.009484f
C182 B.n145 VSUBS 0.009484f
C183 B.n146 VSUBS 0.009484f
C184 B.n147 VSUBS 0.009484f
C185 B.n148 VSUBS 0.009484f
C186 B.n149 VSUBS 0.009484f
C187 B.n150 VSUBS 0.009484f
C188 B.n151 VSUBS 0.021888f
C189 B.n152 VSUBS 0.009484f
C190 B.n153 VSUBS 0.009484f
C191 B.n154 VSUBS 0.009484f
C192 B.n155 VSUBS 0.009484f
C193 B.n156 VSUBS 0.009484f
C194 B.n157 VSUBS 0.009484f
C195 B.n158 VSUBS 0.009484f
C196 B.n159 VSUBS 0.009484f
C197 B.n160 VSUBS 0.009484f
C198 B.n161 VSUBS 0.009484f
C199 B.n162 VSUBS 0.009484f
C200 B.n163 VSUBS 0.009484f
C201 B.n164 VSUBS 0.009484f
C202 B.n165 VSUBS 0.009484f
C203 B.n166 VSUBS 0.009484f
C204 B.n167 VSUBS 0.009484f
C205 B.n168 VSUBS 0.009484f
C206 B.n169 VSUBS 0.009484f
C207 B.n170 VSUBS 0.009484f
C208 B.n171 VSUBS 0.009484f
C209 B.n172 VSUBS 0.009484f
C210 B.n173 VSUBS 0.009484f
C211 B.n174 VSUBS 0.009484f
C212 B.n175 VSUBS 0.009484f
C213 B.n176 VSUBS 0.009484f
C214 B.n177 VSUBS 0.009484f
C215 B.n178 VSUBS 0.009484f
C216 B.n179 VSUBS 0.009484f
C217 B.n180 VSUBS 0.009484f
C218 B.n181 VSUBS 0.009484f
C219 B.n182 VSUBS 0.009484f
C220 B.n183 VSUBS 0.009484f
C221 B.n184 VSUBS 0.009484f
C222 B.n185 VSUBS 0.009484f
C223 B.n186 VSUBS 0.009484f
C224 B.n187 VSUBS 0.009484f
C225 B.n188 VSUBS 0.009484f
C226 B.n189 VSUBS 0.009484f
C227 B.n190 VSUBS 0.009484f
C228 B.n191 VSUBS 0.009484f
C229 B.n192 VSUBS 0.009484f
C230 B.n193 VSUBS 0.009484f
C231 B.n194 VSUBS 0.009484f
C232 B.n195 VSUBS 0.009484f
C233 B.n196 VSUBS 0.009484f
C234 B.n197 VSUBS 0.009484f
C235 B.n198 VSUBS 0.009484f
C236 B.n199 VSUBS 0.009484f
C237 B.n200 VSUBS 0.009484f
C238 B.n201 VSUBS 0.009484f
C239 B.n202 VSUBS 0.009484f
C240 B.n203 VSUBS 0.009484f
C241 B.n204 VSUBS 0.009484f
C242 B.n205 VSUBS 0.009484f
C243 B.n206 VSUBS 0.009484f
C244 B.n207 VSUBS 0.009484f
C245 B.n208 VSUBS 0.009484f
C246 B.n209 VSUBS 0.009484f
C247 B.n210 VSUBS 0.009484f
C248 B.n211 VSUBS 0.009484f
C249 B.n212 VSUBS 0.009484f
C250 B.n213 VSUBS 0.009484f
C251 B.n214 VSUBS 0.009484f
C252 B.n215 VSUBS 0.009484f
C253 B.n216 VSUBS 0.009484f
C254 B.n217 VSUBS 0.009484f
C255 B.n218 VSUBS 0.009484f
C256 B.n219 VSUBS 0.009484f
C257 B.n220 VSUBS 0.009484f
C258 B.n221 VSUBS 0.009484f
C259 B.n222 VSUBS 0.009484f
C260 B.n223 VSUBS 0.009484f
C261 B.n224 VSUBS 0.009484f
C262 B.n225 VSUBS 0.009484f
C263 B.n226 VSUBS 0.009484f
C264 B.n227 VSUBS 0.009484f
C265 B.n228 VSUBS 0.009484f
C266 B.n229 VSUBS 0.009484f
C267 B.n230 VSUBS 0.009484f
C268 B.n231 VSUBS 0.009484f
C269 B.n232 VSUBS 0.009484f
C270 B.n233 VSUBS 0.009484f
C271 B.n234 VSUBS 0.009484f
C272 B.n235 VSUBS 0.009484f
C273 B.n236 VSUBS 0.009484f
C274 B.n237 VSUBS 0.009484f
C275 B.n238 VSUBS 0.009484f
C276 B.n239 VSUBS 0.009484f
C277 B.n240 VSUBS 0.009484f
C278 B.n241 VSUBS 0.009484f
C279 B.n242 VSUBS 0.009484f
C280 B.n243 VSUBS 0.009484f
C281 B.n244 VSUBS 0.009484f
C282 B.n245 VSUBS 0.009484f
C283 B.n246 VSUBS 0.009484f
C284 B.n247 VSUBS 0.009484f
C285 B.n248 VSUBS 0.009484f
C286 B.n249 VSUBS 0.009484f
C287 B.n250 VSUBS 0.009484f
C288 B.n251 VSUBS 0.009484f
C289 B.n252 VSUBS 0.009484f
C290 B.n253 VSUBS 0.009484f
C291 B.n254 VSUBS 0.009484f
C292 B.n255 VSUBS 0.009484f
C293 B.n256 VSUBS 0.009484f
C294 B.n257 VSUBS 0.009484f
C295 B.n258 VSUBS 0.009484f
C296 B.n259 VSUBS 0.009484f
C297 B.n260 VSUBS 0.009484f
C298 B.n261 VSUBS 0.009484f
C299 B.n262 VSUBS 0.021888f
C300 B.n263 VSUBS 0.022462f
C301 B.n264 VSUBS 0.022462f
C302 B.n265 VSUBS 0.009484f
C303 B.n266 VSUBS 0.009484f
C304 B.n267 VSUBS 0.009484f
C305 B.n268 VSUBS 0.009484f
C306 B.n269 VSUBS 0.009484f
C307 B.n270 VSUBS 0.009484f
C308 B.n271 VSUBS 0.009484f
C309 B.n272 VSUBS 0.009484f
C310 B.n273 VSUBS 0.009484f
C311 B.n274 VSUBS 0.009484f
C312 B.n275 VSUBS 0.009484f
C313 B.n276 VSUBS 0.009484f
C314 B.n277 VSUBS 0.009484f
C315 B.n278 VSUBS 0.009484f
C316 B.n279 VSUBS 0.009484f
C317 B.n280 VSUBS 0.009484f
C318 B.n281 VSUBS 0.009484f
C319 B.n282 VSUBS 0.009484f
C320 B.n283 VSUBS 0.009484f
C321 B.n284 VSUBS 0.009484f
C322 B.n285 VSUBS 0.009484f
C323 B.n286 VSUBS 0.009484f
C324 B.n287 VSUBS 0.009484f
C325 B.n288 VSUBS 0.009484f
C326 B.n289 VSUBS 0.009484f
C327 B.n290 VSUBS 0.009484f
C328 B.n291 VSUBS 0.009484f
C329 B.n292 VSUBS 0.009484f
C330 B.n293 VSUBS 0.009484f
C331 B.n294 VSUBS 0.009484f
C332 B.n295 VSUBS 0.009484f
C333 B.n296 VSUBS 0.009484f
C334 B.n297 VSUBS 0.008926f
C335 B.n298 VSUBS 0.021972f
C336 B.n299 VSUBS 0.0053f
C337 B.n300 VSUBS 0.009484f
C338 B.n301 VSUBS 0.009484f
C339 B.n302 VSUBS 0.009484f
C340 B.n303 VSUBS 0.009484f
C341 B.n304 VSUBS 0.009484f
C342 B.n305 VSUBS 0.009484f
C343 B.n306 VSUBS 0.009484f
C344 B.n307 VSUBS 0.009484f
C345 B.n308 VSUBS 0.009484f
C346 B.n309 VSUBS 0.009484f
C347 B.n310 VSUBS 0.009484f
C348 B.n311 VSUBS 0.009484f
C349 B.t11 VSUBS 0.115751f
C350 B.t10 VSUBS 0.154441f
C351 B.t9 VSUBS 1.12996f
C352 B.n312 VSUBS 0.261922f
C353 B.n313 VSUBS 0.209504f
C354 B.n314 VSUBS 0.021972f
C355 B.n315 VSUBS 0.0053f
C356 B.n316 VSUBS 0.009484f
C357 B.n317 VSUBS 0.009484f
C358 B.n318 VSUBS 0.009484f
C359 B.n319 VSUBS 0.009484f
C360 B.n320 VSUBS 0.009484f
C361 B.n321 VSUBS 0.009484f
C362 B.n322 VSUBS 0.009484f
C363 B.n323 VSUBS 0.009484f
C364 B.n324 VSUBS 0.009484f
C365 B.n325 VSUBS 0.009484f
C366 B.n326 VSUBS 0.009484f
C367 B.n327 VSUBS 0.009484f
C368 B.n328 VSUBS 0.009484f
C369 B.n329 VSUBS 0.009484f
C370 B.n330 VSUBS 0.009484f
C371 B.n331 VSUBS 0.009484f
C372 B.n332 VSUBS 0.009484f
C373 B.n333 VSUBS 0.009484f
C374 B.n334 VSUBS 0.009484f
C375 B.n335 VSUBS 0.009484f
C376 B.n336 VSUBS 0.009484f
C377 B.n337 VSUBS 0.009484f
C378 B.n338 VSUBS 0.009484f
C379 B.n339 VSUBS 0.009484f
C380 B.n340 VSUBS 0.009484f
C381 B.n341 VSUBS 0.009484f
C382 B.n342 VSUBS 0.009484f
C383 B.n343 VSUBS 0.009484f
C384 B.n344 VSUBS 0.009484f
C385 B.n345 VSUBS 0.009484f
C386 B.n346 VSUBS 0.009484f
C387 B.n347 VSUBS 0.009484f
C388 B.n348 VSUBS 0.009484f
C389 B.n349 VSUBS 0.009484f
C390 B.n350 VSUBS 0.02134f
C391 B.n351 VSUBS 0.023009f
C392 B.n352 VSUBS 0.021888f
C393 B.n353 VSUBS 0.009484f
C394 B.n354 VSUBS 0.009484f
C395 B.n355 VSUBS 0.009484f
C396 B.n356 VSUBS 0.009484f
C397 B.n357 VSUBS 0.009484f
C398 B.n358 VSUBS 0.009484f
C399 B.n359 VSUBS 0.009484f
C400 B.n360 VSUBS 0.009484f
C401 B.n361 VSUBS 0.009484f
C402 B.n362 VSUBS 0.009484f
C403 B.n363 VSUBS 0.009484f
C404 B.n364 VSUBS 0.009484f
C405 B.n365 VSUBS 0.009484f
C406 B.n366 VSUBS 0.009484f
C407 B.n367 VSUBS 0.009484f
C408 B.n368 VSUBS 0.009484f
C409 B.n369 VSUBS 0.009484f
C410 B.n370 VSUBS 0.009484f
C411 B.n371 VSUBS 0.009484f
C412 B.n372 VSUBS 0.009484f
C413 B.n373 VSUBS 0.009484f
C414 B.n374 VSUBS 0.009484f
C415 B.n375 VSUBS 0.009484f
C416 B.n376 VSUBS 0.009484f
C417 B.n377 VSUBS 0.009484f
C418 B.n378 VSUBS 0.009484f
C419 B.n379 VSUBS 0.009484f
C420 B.n380 VSUBS 0.009484f
C421 B.n381 VSUBS 0.009484f
C422 B.n382 VSUBS 0.009484f
C423 B.n383 VSUBS 0.009484f
C424 B.n384 VSUBS 0.009484f
C425 B.n385 VSUBS 0.009484f
C426 B.n386 VSUBS 0.009484f
C427 B.n387 VSUBS 0.009484f
C428 B.n388 VSUBS 0.009484f
C429 B.n389 VSUBS 0.009484f
C430 B.n390 VSUBS 0.009484f
C431 B.n391 VSUBS 0.009484f
C432 B.n392 VSUBS 0.009484f
C433 B.n393 VSUBS 0.009484f
C434 B.n394 VSUBS 0.009484f
C435 B.n395 VSUBS 0.009484f
C436 B.n396 VSUBS 0.009484f
C437 B.n397 VSUBS 0.009484f
C438 B.n398 VSUBS 0.009484f
C439 B.n399 VSUBS 0.009484f
C440 B.n400 VSUBS 0.009484f
C441 B.n401 VSUBS 0.009484f
C442 B.n402 VSUBS 0.009484f
C443 B.n403 VSUBS 0.009484f
C444 B.n404 VSUBS 0.009484f
C445 B.n405 VSUBS 0.009484f
C446 B.n406 VSUBS 0.009484f
C447 B.n407 VSUBS 0.009484f
C448 B.n408 VSUBS 0.009484f
C449 B.n409 VSUBS 0.009484f
C450 B.n410 VSUBS 0.009484f
C451 B.n411 VSUBS 0.009484f
C452 B.n412 VSUBS 0.009484f
C453 B.n413 VSUBS 0.009484f
C454 B.n414 VSUBS 0.009484f
C455 B.n415 VSUBS 0.009484f
C456 B.n416 VSUBS 0.009484f
C457 B.n417 VSUBS 0.009484f
C458 B.n418 VSUBS 0.009484f
C459 B.n419 VSUBS 0.009484f
C460 B.n420 VSUBS 0.009484f
C461 B.n421 VSUBS 0.009484f
C462 B.n422 VSUBS 0.009484f
C463 B.n423 VSUBS 0.009484f
C464 B.n424 VSUBS 0.009484f
C465 B.n425 VSUBS 0.009484f
C466 B.n426 VSUBS 0.009484f
C467 B.n427 VSUBS 0.009484f
C468 B.n428 VSUBS 0.009484f
C469 B.n429 VSUBS 0.009484f
C470 B.n430 VSUBS 0.009484f
C471 B.n431 VSUBS 0.009484f
C472 B.n432 VSUBS 0.009484f
C473 B.n433 VSUBS 0.009484f
C474 B.n434 VSUBS 0.009484f
C475 B.n435 VSUBS 0.009484f
C476 B.n436 VSUBS 0.009484f
C477 B.n437 VSUBS 0.009484f
C478 B.n438 VSUBS 0.009484f
C479 B.n439 VSUBS 0.009484f
C480 B.n440 VSUBS 0.009484f
C481 B.n441 VSUBS 0.009484f
C482 B.n442 VSUBS 0.009484f
C483 B.n443 VSUBS 0.009484f
C484 B.n444 VSUBS 0.009484f
C485 B.n445 VSUBS 0.009484f
C486 B.n446 VSUBS 0.009484f
C487 B.n447 VSUBS 0.009484f
C488 B.n448 VSUBS 0.009484f
C489 B.n449 VSUBS 0.009484f
C490 B.n450 VSUBS 0.009484f
C491 B.n451 VSUBS 0.009484f
C492 B.n452 VSUBS 0.009484f
C493 B.n453 VSUBS 0.009484f
C494 B.n454 VSUBS 0.009484f
C495 B.n455 VSUBS 0.009484f
C496 B.n456 VSUBS 0.009484f
C497 B.n457 VSUBS 0.009484f
C498 B.n458 VSUBS 0.009484f
C499 B.n459 VSUBS 0.009484f
C500 B.n460 VSUBS 0.009484f
C501 B.n461 VSUBS 0.009484f
C502 B.n462 VSUBS 0.009484f
C503 B.n463 VSUBS 0.009484f
C504 B.n464 VSUBS 0.009484f
C505 B.n465 VSUBS 0.009484f
C506 B.n466 VSUBS 0.009484f
C507 B.n467 VSUBS 0.009484f
C508 B.n468 VSUBS 0.009484f
C509 B.n469 VSUBS 0.009484f
C510 B.n470 VSUBS 0.009484f
C511 B.n471 VSUBS 0.009484f
C512 B.n472 VSUBS 0.009484f
C513 B.n473 VSUBS 0.009484f
C514 B.n474 VSUBS 0.009484f
C515 B.n475 VSUBS 0.009484f
C516 B.n476 VSUBS 0.009484f
C517 B.n477 VSUBS 0.009484f
C518 B.n478 VSUBS 0.009484f
C519 B.n479 VSUBS 0.009484f
C520 B.n480 VSUBS 0.009484f
C521 B.n481 VSUBS 0.009484f
C522 B.n482 VSUBS 0.009484f
C523 B.n483 VSUBS 0.009484f
C524 B.n484 VSUBS 0.009484f
C525 B.n485 VSUBS 0.009484f
C526 B.n486 VSUBS 0.009484f
C527 B.n487 VSUBS 0.009484f
C528 B.n488 VSUBS 0.009484f
C529 B.n489 VSUBS 0.009484f
C530 B.n490 VSUBS 0.009484f
C531 B.n491 VSUBS 0.009484f
C532 B.n492 VSUBS 0.009484f
C533 B.n493 VSUBS 0.009484f
C534 B.n494 VSUBS 0.009484f
C535 B.n495 VSUBS 0.009484f
C536 B.n496 VSUBS 0.009484f
C537 B.n497 VSUBS 0.009484f
C538 B.n498 VSUBS 0.009484f
C539 B.n499 VSUBS 0.009484f
C540 B.n500 VSUBS 0.009484f
C541 B.n501 VSUBS 0.009484f
C542 B.n502 VSUBS 0.009484f
C543 B.n503 VSUBS 0.009484f
C544 B.n504 VSUBS 0.009484f
C545 B.n505 VSUBS 0.009484f
C546 B.n506 VSUBS 0.009484f
C547 B.n507 VSUBS 0.009484f
C548 B.n508 VSUBS 0.009484f
C549 B.n509 VSUBS 0.009484f
C550 B.n510 VSUBS 0.009484f
C551 B.n511 VSUBS 0.009484f
C552 B.n512 VSUBS 0.009484f
C553 B.n513 VSUBS 0.009484f
C554 B.n514 VSUBS 0.009484f
C555 B.n515 VSUBS 0.009484f
C556 B.n516 VSUBS 0.009484f
C557 B.n517 VSUBS 0.009484f
C558 B.n518 VSUBS 0.009484f
C559 B.n519 VSUBS 0.009484f
C560 B.n520 VSUBS 0.009484f
C561 B.n521 VSUBS 0.009484f
C562 B.n522 VSUBS 0.009484f
C563 B.n523 VSUBS 0.009484f
C564 B.n524 VSUBS 0.021888f
C565 B.n525 VSUBS 0.022462f
C566 B.n526 VSUBS 0.022462f
C567 B.n527 VSUBS 0.009484f
C568 B.n528 VSUBS 0.009484f
C569 B.n529 VSUBS 0.009484f
C570 B.n530 VSUBS 0.009484f
C571 B.n531 VSUBS 0.009484f
C572 B.n532 VSUBS 0.009484f
C573 B.n533 VSUBS 0.009484f
C574 B.n534 VSUBS 0.009484f
C575 B.n535 VSUBS 0.009484f
C576 B.n536 VSUBS 0.009484f
C577 B.n537 VSUBS 0.009484f
C578 B.n538 VSUBS 0.009484f
C579 B.n539 VSUBS 0.009484f
C580 B.n540 VSUBS 0.009484f
C581 B.n541 VSUBS 0.009484f
C582 B.n542 VSUBS 0.009484f
C583 B.n543 VSUBS 0.009484f
C584 B.n544 VSUBS 0.009484f
C585 B.n545 VSUBS 0.009484f
C586 B.n546 VSUBS 0.009484f
C587 B.n547 VSUBS 0.009484f
C588 B.n548 VSUBS 0.009484f
C589 B.n549 VSUBS 0.009484f
C590 B.n550 VSUBS 0.009484f
C591 B.n551 VSUBS 0.009484f
C592 B.n552 VSUBS 0.009484f
C593 B.n553 VSUBS 0.009484f
C594 B.n554 VSUBS 0.009484f
C595 B.n555 VSUBS 0.009484f
C596 B.n556 VSUBS 0.009484f
C597 B.n557 VSUBS 0.009484f
C598 B.n558 VSUBS 0.009484f
C599 B.n559 VSUBS 0.008926f
C600 B.n560 VSUBS 0.021972f
C601 B.n561 VSUBS 0.0053f
C602 B.n562 VSUBS 0.009484f
C603 B.n563 VSUBS 0.009484f
C604 B.n564 VSUBS 0.009484f
C605 B.n565 VSUBS 0.009484f
C606 B.n566 VSUBS 0.009484f
C607 B.n567 VSUBS 0.009484f
C608 B.n568 VSUBS 0.009484f
C609 B.n569 VSUBS 0.009484f
C610 B.n570 VSUBS 0.009484f
C611 B.n571 VSUBS 0.009484f
C612 B.n572 VSUBS 0.009484f
C613 B.n573 VSUBS 0.009484f
C614 B.n574 VSUBS 0.0053f
C615 B.n575 VSUBS 0.009484f
C616 B.n576 VSUBS 0.009484f
C617 B.n577 VSUBS 0.008926f
C618 B.n578 VSUBS 0.009484f
C619 B.n579 VSUBS 0.009484f
C620 B.n580 VSUBS 0.009484f
C621 B.n581 VSUBS 0.009484f
C622 B.n582 VSUBS 0.009484f
C623 B.n583 VSUBS 0.009484f
C624 B.n584 VSUBS 0.009484f
C625 B.n585 VSUBS 0.009484f
C626 B.n586 VSUBS 0.009484f
C627 B.n587 VSUBS 0.009484f
C628 B.n588 VSUBS 0.009484f
C629 B.n589 VSUBS 0.009484f
C630 B.n590 VSUBS 0.009484f
C631 B.n591 VSUBS 0.009484f
C632 B.n592 VSUBS 0.009484f
C633 B.n593 VSUBS 0.009484f
C634 B.n594 VSUBS 0.009484f
C635 B.n595 VSUBS 0.009484f
C636 B.n596 VSUBS 0.009484f
C637 B.n597 VSUBS 0.009484f
C638 B.n598 VSUBS 0.009484f
C639 B.n599 VSUBS 0.009484f
C640 B.n600 VSUBS 0.009484f
C641 B.n601 VSUBS 0.009484f
C642 B.n602 VSUBS 0.009484f
C643 B.n603 VSUBS 0.009484f
C644 B.n604 VSUBS 0.009484f
C645 B.n605 VSUBS 0.009484f
C646 B.n606 VSUBS 0.009484f
C647 B.n607 VSUBS 0.009484f
C648 B.n608 VSUBS 0.009484f
C649 B.n609 VSUBS 0.022462f
C650 B.n610 VSUBS 0.022462f
C651 B.n611 VSUBS 0.021888f
C652 B.n612 VSUBS 0.009484f
C653 B.n613 VSUBS 0.009484f
C654 B.n614 VSUBS 0.009484f
C655 B.n615 VSUBS 0.009484f
C656 B.n616 VSUBS 0.009484f
C657 B.n617 VSUBS 0.009484f
C658 B.n618 VSUBS 0.009484f
C659 B.n619 VSUBS 0.009484f
C660 B.n620 VSUBS 0.009484f
C661 B.n621 VSUBS 0.009484f
C662 B.n622 VSUBS 0.009484f
C663 B.n623 VSUBS 0.009484f
C664 B.n624 VSUBS 0.009484f
C665 B.n625 VSUBS 0.009484f
C666 B.n626 VSUBS 0.009484f
C667 B.n627 VSUBS 0.009484f
C668 B.n628 VSUBS 0.009484f
C669 B.n629 VSUBS 0.009484f
C670 B.n630 VSUBS 0.009484f
C671 B.n631 VSUBS 0.009484f
C672 B.n632 VSUBS 0.009484f
C673 B.n633 VSUBS 0.009484f
C674 B.n634 VSUBS 0.009484f
C675 B.n635 VSUBS 0.009484f
C676 B.n636 VSUBS 0.009484f
C677 B.n637 VSUBS 0.009484f
C678 B.n638 VSUBS 0.009484f
C679 B.n639 VSUBS 0.009484f
C680 B.n640 VSUBS 0.009484f
C681 B.n641 VSUBS 0.009484f
C682 B.n642 VSUBS 0.009484f
C683 B.n643 VSUBS 0.009484f
C684 B.n644 VSUBS 0.009484f
C685 B.n645 VSUBS 0.009484f
C686 B.n646 VSUBS 0.009484f
C687 B.n647 VSUBS 0.009484f
C688 B.n648 VSUBS 0.009484f
C689 B.n649 VSUBS 0.009484f
C690 B.n650 VSUBS 0.009484f
C691 B.n651 VSUBS 0.009484f
C692 B.n652 VSUBS 0.009484f
C693 B.n653 VSUBS 0.009484f
C694 B.n654 VSUBS 0.009484f
C695 B.n655 VSUBS 0.009484f
C696 B.n656 VSUBS 0.009484f
C697 B.n657 VSUBS 0.009484f
C698 B.n658 VSUBS 0.009484f
C699 B.n659 VSUBS 0.009484f
C700 B.n660 VSUBS 0.009484f
C701 B.n661 VSUBS 0.009484f
C702 B.n662 VSUBS 0.009484f
C703 B.n663 VSUBS 0.009484f
C704 B.n664 VSUBS 0.009484f
C705 B.n665 VSUBS 0.009484f
C706 B.n666 VSUBS 0.009484f
C707 B.n667 VSUBS 0.009484f
C708 B.n668 VSUBS 0.009484f
C709 B.n669 VSUBS 0.009484f
C710 B.n670 VSUBS 0.009484f
C711 B.n671 VSUBS 0.009484f
C712 B.n672 VSUBS 0.009484f
C713 B.n673 VSUBS 0.009484f
C714 B.n674 VSUBS 0.009484f
C715 B.n675 VSUBS 0.009484f
C716 B.n676 VSUBS 0.009484f
C717 B.n677 VSUBS 0.009484f
C718 B.n678 VSUBS 0.009484f
C719 B.n679 VSUBS 0.009484f
C720 B.n680 VSUBS 0.009484f
C721 B.n681 VSUBS 0.009484f
C722 B.n682 VSUBS 0.009484f
C723 B.n683 VSUBS 0.009484f
C724 B.n684 VSUBS 0.009484f
C725 B.n685 VSUBS 0.009484f
C726 B.n686 VSUBS 0.009484f
C727 B.n687 VSUBS 0.009484f
C728 B.n688 VSUBS 0.009484f
C729 B.n689 VSUBS 0.009484f
C730 B.n690 VSUBS 0.009484f
C731 B.n691 VSUBS 0.009484f
C732 B.n692 VSUBS 0.009484f
C733 B.n693 VSUBS 0.009484f
C734 B.n694 VSUBS 0.009484f
C735 B.n695 VSUBS 0.012376f
C736 B.n696 VSUBS 0.013183f
C737 B.n697 VSUBS 0.026216f
C738 VDD2.t2 VSUBS 0.130912f
C739 VDD2.t1 VSUBS 0.130912f
C740 VDD2.n0 VSUBS 0.890301f
C741 VDD2.t5 VSUBS 0.130912f
C742 VDD2.t4 VSUBS 0.130912f
C743 VDD2.n1 VSUBS 0.890301f
C744 VDD2.n2 VSUBS 4.00294f
C745 VDD2.t7 VSUBS 0.130912f
C746 VDD2.t0 VSUBS 0.130912f
C747 VDD2.n3 VSUBS 0.878045f
C748 VDD2.n4 VSUBS 3.20088f
C749 VDD2.t6 VSUBS 0.130912f
C750 VDD2.t3 VSUBS 0.130912f
C751 VDD2.n5 VSUBS 0.890263f
C752 VN.n0 VSUBS 0.045802f
C753 VN.t3 VSUBS 1.6044f
C754 VN.n1 VSUBS 0.066435f
C755 VN.n2 VSUBS 0.034741f
C756 VN.n3 VSUBS 0.053558f
C757 VN.n4 VSUBS 0.034741f
C758 VN.n5 VSUBS 0.028085f
C759 VN.n6 VSUBS 0.034741f
C760 VN.t6 VSUBS 1.6044f
C761 VN.n7 VSUBS 0.705835f
C762 VN.t5 VSUBS 1.95026f
C763 VN.n8 VSUBS 0.681523f
C764 VN.n9 VSUBS 0.37322f
C765 VN.n10 VSUBS 0.043968f
C766 VN.n11 VSUBS 0.064748f
C767 VN.n12 VSUBS 0.069047f
C768 VN.n13 VSUBS 0.034741f
C769 VN.n14 VSUBS 0.034741f
C770 VN.n15 VSUBS 0.034741f
C771 VN.n16 VSUBS 0.069047f
C772 VN.n17 VSUBS 0.064748f
C773 VN.t2 VSUBS 1.6044f
C774 VN.n18 VSUBS 0.599434f
C775 VN.n19 VSUBS 0.043968f
C776 VN.n20 VSUBS 0.034741f
C777 VN.n21 VSUBS 0.034741f
C778 VN.n22 VSUBS 0.034741f
C779 VN.n23 VSUBS 0.064748f
C780 VN.n24 VSUBS 0.060127f
C781 VN.n25 VSUBS 0.039617f
C782 VN.n26 VSUBS 0.034741f
C783 VN.n27 VSUBS 0.034741f
C784 VN.n28 VSUBS 0.034741f
C785 VN.n29 VSUBS 0.064748f
C786 VN.n30 VSUBS 0.034378f
C787 VN.n31 VSUBS 0.718399f
C788 VN.n32 VSUBS 0.069181f
C789 VN.n33 VSUBS 0.045802f
C790 VN.t0 VSUBS 1.6044f
C791 VN.n34 VSUBS 0.066435f
C792 VN.n35 VSUBS 0.034741f
C793 VN.n36 VSUBS 0.053558f
C794 VN.n37 VSUBS 0.034741f
C795 VN.t7 VSUBS 1.6044f
C796 VN.n38 VSUBS 0.599434f
C797 VN.n39 VSUBS 0.028085f
C798 VN.n40 VSUBS 0.034741f
C799 VN.t1 VSUBS 1.6044f
C800 VN.n41 VSUBS 0.705835f
C801 VN.t4 VSUBS 1.95026f
C802 VN.n42 VSUBS 0.681523f
C803 VN.n43 VSUBS 0.37322f
C804 VN.n44 VSUBS 0.043968f
C805 VN.n45 VSUBS 0.064748f
C806 VN.n46 VSUBS 0.069047f
C807 VN.n47 VSUBS 0.034741f
C808 VN.n48 VSUBS 0.034741f
C809 VN.n49 VSUBS 0.034741f
C810 VN.n50 VSUBS 0.069047f
C811 VN.n51 VSUBS 0.064748f
C812 VN.n52 VSUBS 0.043968f
C813 VN.n53 VSUBS 0.034741f
C814 VN.n54 VSUBS 0.034741f
C815 VN.n55 VSUBS 0.034741f
C816 VN.n56 VSUBS 0.064748f
C817 VN.n57 VSUBS 0.060127f
C818 VN.n58 VSUBS 0.039617f
C819 VN.n59 VSUBS 0.034741f
C820 VN.n60 VSUBS 0.034741f
C821 VN.n61 VSUBS 0.034741f
C822 VN.n62 VSUBS 0.064748f
C823 VN.n63 VSUBS 0.034378f
C824 VN.n64 VSUBS 0.718399f
C825 VN.n65 VSUBS 1.8596f
C826 VTAIL.t3 VSUBS 0.138576f
C827 VTAIL.t5 VSUBS 0.138576f
C828 VTAIL.n0 VSUBS 0.830804f
C829 VTAIL.n1 VSUBS 0.811183f
C830 VTAIL.n2 VSUBS 0.017041f
C831 VTAIL.n3 VSUBS 0.038468f
C832 VTAIL.n4 VSUBS 0.017232f
C833 VTAIL.n5 VSUBS 0.030287f
C834 VTAIL.n6 VSUBS 0.016275f
C835 VTAIL.n7 VSUBS 0.038468f
C836 VTAIL.n8 VSUBS 0.017232f
C837 VTAIL.n9 VSUBS 0.663036f
C838 VTAIL.n10 VSUBS 0.016275f
C839 VTAIL.t0 VSUBS 0.082798f
C840 VTAIL.n11 VSUBS 0.15391f
C841 VTAIL.n12 VSUBS 0.028925f
C842 VTAIL.n13 VSUBS 0.028851f
C843 VTAIL.n14 VSUBS 0.038468f
C844 VTAIL.n15 VSUBS 0.017232f
C845 VTAIL.n16 VSUBS 0.016275f
C846 VTAIL.n17 VSUBS 0.030287f
C847 VTAIL.n18 VSUBS 0.030287f
C848 VTAIL.n19 VSUBS 0.016275f
C849 VTAIL.n20 VSUBS 0.017232f
C850 VTAIL.n21 VSUBS 0.038468f
C851 VTAIL.n22 VSUBS 0.038468f
C852 VTAIL.n23 VSUBS 0.017232f
C853 VTAIL.n24 VSUBS 0.016275f
C854 VTAIL.n25 VSUBS 0.030287f
C855 VTAIL.n26 VSUBS 0.076213f
C856 VTAIL.n27 VSUBS 0.016275f
C857 VTAIL.n28 VSUBS 0.017232f
C858 VTAIL.n29 VSUBS 0.083512f
C859 VTAIL.n30 VSUBS 0.055617f
C860 VTAIL.n31 VSUBS 0.35566f
C861 VTAIL.n32 VSUBS 0.017041f
C862 VTAIL.n33 VSUBS 0.038468f
C863 VTAIL.n34 VSUBS 0.017232f
C864 VTAIL.n35 VSUBS 0.030287f
C865 VTAIL.n36 VSUBS 0.016275f
C866 VTAIL.n37 VSUBS 0.038468f
C867 VTAIL.n38 VSUBS 0.017232f
C868 VTAIL.n39 VSUBS 0.663036f
C869 VTAIL.n40 VSUBS 0.016275f
C870 VTAIL.t9 VSUBS 0.082798f
C871 VTAIL.n41 VSUBS 0.15391f
C872 VTAIL.n42 VSUBS 0.028925f
C873 VTAIL.n43 VSUBS 0.028851f
C874 VTAIL.n44 VSUBS 0.038468f
C875 VTAIL.n45 VSUBS 0.017232f
C876 VTAIL.n46 VSUBS 0.016275f
C877 VTAIL.n47 VSUBS 0.030287f
C878 VTAIL.n48 VSUBS 0.030287f
C879 VTAIL.n49 VSUBS 0.016275f
C880 VTAIL.n50 VSUBS 0.017232f
C881 VTAIL.n51 VSUBS 0.038468f
C882 VTAIL.n52 VSUBS 0.038468f
C883 VTAIL.n53 VSUBS 0.017232f
C884 VTAIL.n54 VSUBS 0.016275f
C885 VTAIL.n55 VSUBS 0.030287f
C886 VTAIL.n56 VSUBS 0.076213f
C887 VTAIL.n57 VSUBS 0.016275f
C888 VTAIL.n58 VSUBS 0.017232f
C889 VTAIL.n59 VSUBS 0.083512f
C890 VTAIL.n60 VSUBS 0.055617f
C891 VTAIL.n61 VSUBS 0.35566f
C892 VTAIL.t13 VSUBS 0.138576f
C893 VTAIL.t8 VSUBS 0.138576f
C894 VTAIL.n62 VSUBS 0.830804f
C895 VTAIL.n63 VSUBS 1.08734f
C896 VTAIL.n64 VSUBS 0.017041f
C897 VTAIL.n65 VSUBS 0.038468f
C898 VTAIL.n66 VSUBS 0.017232f
C899 VTAIL.n67 VSUBS 0.030287f
C900 VTAIL.n68 VSUBS 0.016275f
C901 VTAIL.n69 VSUBS 0.038468f
C902 VTAIL.n70 VSUBS 0.017232f
C903 VTAIL.n71 VSUBS 0.663036f
C904 VTAIL.n72 VSUBS 0.016275f
C905 VTAIL.t12 VSUBS 0.082798f
C906 VTAIL.n73 VSUBS 0.15391f
C907 VTAIL.n74 VSUBS 0.028925f
C908 VTAIL.n75 VSUBS 0.028851f
C909 VTAIL.n76 VSUBS 0.038468f
C910 VTAIL.n77 VSUBS 0.017232f
C911 VTAIL.n78 VSUBS 0.016275f
C912 VTAIL.n79 VSUBS 0.030287f
C913 VTAIL.n80 VSUBS 0.030287f
C914 VTAIL.n81 VSUBS 0.016275f
C915 VTAIL.n82 VSUBS 0.017232f
C916 VTAIL.n83 VSUBS 0.038468f
C917 VTAIL.n84 VSUBS 0.038468f
C918 VTAIL.n85 VSUBS 0.017232f
C919 VTAIL.n86 VSUBS 0.016275f
C920 VTAIL.n87 VSUBS 0.030287f
C921 VTAIL.n88 VSUBS 0.076213f
C922 VTAIL.n89 VSUBS 0.016275f
C923 VTAIL.n90 VSUBS 0.017232f
C924 VTAIL.n91 VSUBS 0.083512f
C925 VTAIL.n92 VSUBS 0.055617f
C926 VTAIL.n93 VSUBS 1.49017f
C927 VTAIL.n94 VSUBS 0.017041f
C928 VTAIL.n95 VSUBS 0.038468f
C929 VTAIL.n96 VSUBS 0.017232f
C930 VTAIL.n97 VSUBS 0.030287f
C931 VTAIL.n98 VSUBS 0.016275f
C932 VTAIL.n99 VSUBS 0.038468f
C933 VTAIL.n100 VSUBS 0.017232f
C934 VTAIL.n101 VSUBS 0.663036f
C935 VTAIL.n102 VSUBS 0.016275f
C936 VTAIL.t6 VSUBS 0.082798f
C937 VTAIL.n103 VSUBS 0.15391f
C938 VTAIL.n104 VSUBS 0.028925f
C939 VTAIL.n105 VSUBS 0.028851f
C940 VTAIL.n106 VSUBS 0.038468f
C941 VTAIL.n107 VSUBS 0.017232f
C942 VTAIL.n108 VSUBS 0.016275f
C943 VTAIL.n109 VSUBS 0.030287f
C944 VTAIL.n110 VSUBS 0.030287f
C945 VTAIL.n111 VSUBS 0.016275f
C946 VTAIL.n112 VSUBS 0.017232f
C947 VTAIL.n113 VSUBS 0.038468f
C948 VTAIL.n114 VSUBS 0.038468f
C949 VTAIL.n115 VSUBS 0.017232f
C950 VTAIL.n116 VSUBS 0.016275f
C951 VTAIL.n117 VSUBS 0.030287f
C952 VTAIL.n118 VSUBS 0.076213f
C953 VTAIL.n119 VSUBS 0.016275f
C954 VTAIL.n120 VSUBS 0.017232f
C955 VTAIL.n121 VSUBS 0.083512f
C956 VTAIL.n122 VSUBS 0.055617f
C957 VTAIL.n123 VSUBS 1.49017f
C958 VTAIL.t4 VSUBS 0.138576f
C959 VTAIL.t7 VSUBS 0.138576f
C960 VTAIL.n124 VSUBS 0.830808f
C961 VTAIL.n125 VSUBS 1.08734f
C962 VTAIL.n126 VSUBS 0.017041f
C963 VTAIL.n127 VSUBS 0.038468f
C964 VTAIL.n128 VSUBS 0.017232f
C965 VTAIL.n129 VSUBS 0.030287f
C966 VTAIL.n130 VSUBS 0.016275f
C967 VTAIL.n131 VSUBS 0.038468f
C968 VTAIL.n132 VSUBS 0.017232f
C969 VTAIL.n133 VSUBS 0.663036f
C970 VTAIL.n134 VSUBS 0.016275f
C971 VTAIL.t2 VSUBS 0.082798f
C972 VTAIL.n135 VSUBS 0.15391f
C973 VTAIL.n136 VSUBS 0.028925f
C974 VTAIL.n137 VSUBS 0.028851f
C975 VTAIL.n138 VSUBS 0.038468f
C976 VTAIL.n139 VSUBS 0.017232f
C977 VTAIL.n140 VSUBS 0.016275f
C978 VTAIL.n141 VSUBS 0.030287f
C979 VTAIL.n142 VSUBS 0.030287f
C980 VTAIL.n143 VSUBS 0.016275f
C981 VTAIL.n144 VSUBS 0.017232f
C982 VTAIL.n145 VSUBS 0.038468f
C983 VTAIL.n146 VSUBS 0.038468f
C984 VTAIL.n147 VSUBS 0.017232f
C985 VTAIL.n148 VSUBS 0.016275f
C986 VTAIL.n149 VSUBS 0.030287f
C987 VTAIL.n150 VSUBS 0.076213f
C988 VTAIL.n151 VSUBS 0.016275f
C989 VTAIL.n152 VSUBS 0.017232f
C990 VTAIL.n153 VSUBS 0.083512f
C991 VTAIL.n154 VSUBS 0.055617f
C992 VTAIL.n155 VSUBS 0.35566f
C993 VTAIL.n156 VSUBS 0.017041f
C994 VTAIL.n157 VSUBS 0.038468f
C995 VTAIL.n158 VSUBS 0.017232f
C996 VTAIL.n159 VSUBS 0.030287f
C997 VTAIL.n160 VSUBS 0.016275f
C998 VTAIL.n161 VSUBS 0.038468f
C999 VTAIL.n162 VSUBS 0.017232f
C1000 VTAIL.n163 VSUBS 0.663036f
C1001 VTAIL.n164 VSUBS 0.016275f
C1002 VTAIL.t14 VSUBS 0.082798f
C1003 VTAIL.n165 VSUBS 0.15391f
C1004 VTAIL.n166 VSUBS 0.028925f
C1005 VTAIL.n167 VSUBS 0.028851f
C1006 VTAIL.n168 VSUBS 0.038468f
C1007 VTAIL.n169 VSUBS 0.017232f
C1008 VTAIL.n170 VSUBS 0.016275f
C1009 VTAIL.n171 VSUBS 0.030287f
C1010 VTAIL.n172 VSUBS 0.030287f
C1011 VTAIL.n173 VSUBS 0.016275f
C1012 VTAIL.n174 VSUBS 0.017232f
C1013 VTAIL.n175 VSUBS 0.038468f
C1014 VTAIL.n176 VSUBS 0.038468f
C1015 VTAIL.n177 VSUBS 0.017232f
C1016 VTAIL.n178 VSUBS 0.016275f
C1017 VTAIL.n179 VSUBS 0.030287f
C1018 VTAIL.n180 VSUBS 0.076213f
C1019 VTAIL.n181 VSUBS 0.016275f
C1020 VTAIL.n182 VSUBS 0.017232f
C1021 VTAIL.n183 VSUBS 0.083512f
C1022 VTAIL.n184 VSUBS 0.055617f
C1023 VTAIL.n185 VSUBS 0.35566f
C1024 VTAIL.t10 VSUBS 0.138576f
C1025 VTAIL.t15 VSUBS 0.138576f
C1026 VTAIL.n186 VSUBS 0.830808f
C1027 VTAIL.n187 VSUBS 1.08734f
C1028 VTAIL.n188 VSUBS 0.017041f
C1029 VTAIL.n189 VSUBS 0.038468f
C1030 VTAIL.n190 VSUBS 0.017232f
C1031 VTAIL.n191 VSUBS 0.030287f
C1032 VTAIL.n192 VSUBS 0.016275f
C1033 VTAIL.n193 VSUBS 0.038468f
C1034 VTAIL.n194 VSUBS 0.017232f
C1035 VTAIL.n195 VSUBS 0.663036f
C1036 VTAIL.n196 VSUBS 0.016275f
C1037 VTAIL.t11 VSUBS 0.082798f
C1038 VTAIL.n197 VSUBS 0.15391f
C1039 VTAIL.n198 VSUBS 0.028925f
C1040 VTAIL.n199 VSUBS 0.028851f
C1041 VTAIL.n200 VSUBS 0.038468f
C1042 VTAIL.n201 VSUBS 0.017232f
C1043 VTAIL.n202 VSUBS 0.016275f
C1044 VTAIL.n203 VSUBS 0.030287f
C1045 VTAIL.n204 VSUBS 0.030287f
C1046 VTAIL.n205 VSUBS 0.016275f
C1047 VTAIL.n206 VSUBS 0.017232f
C1048 VTAIL.n207 VSUBS 0.038468f
C1049 VTAIL.n208 VSUBS 0.038468f
C1050 VTAIL.n209 VSUBS 0.017232f
C1051 VTAIL.n210 VSUBS 0.016275f
C1052 VTAIL.n211 VSUBS 0.030287f
C1053 VTAIL.n212 VSUBS 0.076213f
C1054 VTAIL.n213 VSUBS 0.016275f
C1055 VTAIL.n214 VSUBS 0.017232f
C1056 VTAIL.n215 VSUBS 0.083512f
C1057 VTAIL.n216 VSUBS 0.055617f
C1058 VTAIL.n217 VSUBS 1.49017f
C1059 VTAIL.n218 VSUBS 0.017041f
C1060 VTAIL.n219 VSUBS 0.038468f
C1061 VTAIL.n220 VSUBS 0.017232f
C1062 VTAIL.n221 VSUBS 0.030287f
C1063 VTAIL.n222 VSUBS 0.016275f
C1064 VTAIL.n223 VSUBS 0.038468f
C1065 VTAIL.n224 VSUBS 0.017232f
C1066 VTAIL.n225 VSUBS 0.663036f
C1067 VTAIL.n226 VSUBS 0.016275f
C1068 VTAIL.t1 VSUBS 0.082798f
C1069 VTAIL.n227 VSUBS 0.15391f
C1070 VTAIL.n228 VSUBS 0.028925f
C1071 VTAIL.n229 VSUBS 0.028851f
C1072 VTAIL.n230 VSUBS 0.038468f
C1073 VTAIL.n231 VSUBS 0.017232f
C1074 VTAIL.n232 VSUBS 0.016275f
C1075 VTAIL.n233 VSUBS 0.030287f
C1076 VTAIL.n234 VSUBS 0.030287f
C1077 VTAIL.n235 VSUBS 0.016275f
C1078 VTAIL.n236 VSUBS 0.017232f
C1079 VTAIL.n237 VSUBS 0.038468f
C1080 VTAIL.n238 VSUBS 0.038468f
C1081 VTAIL.n239 VSUBS 0.017232f
C1082 VTAIL.n240 VSUBS 0.016275f
C1083 VTAIL.n241 VSUBS 0.030287f
C1084 VTAIL.n242 VSUBS 0.076213f
C1085 VTAIL.n243 VSUBS 0.016275f
C1086 VTAIL.n244 VSUBS 0.017232f
C1087 VTAIL.n245 VSUBS 0.083512f
C1088 VTAIL.n246 VSUBS 0.055617f
C1089 VTAIL.n247 VSUBS 1.48449f
C1090 VDD1.t1 VSUBS 0.113743f
C1091 VDD1.t4 VSUBS 0.113743f
C1092 VDD1.n0 VSUBS 0.774534f
C1093 VDD1.t0 VSUBS 0.113743f
C1094 VDD1.t2 VSUBS 0.113743f
C1095 VDD1.n1 VSUBS 0.77354f
C1096 VDD1.t7 VSUBS 0.113743f
C1097 VDD1.t3 VSUBS 0.113743f
C1098 VDD1.n2 VSUBS 0.77354f
C1099 VDD1.n3 VSUBS 3.52968f
C1100 VDD1.t5 VSUBS 0.113743f
C1101 VDD1.t6 VSUBS 0.113743f
C1102 VDD1.n4 VSUBS 0.762887f
C1103 VDD1.n5 VSUBS 2.81187f
C1104 VP.n0 VSUBS 0.051736f
C1105 VP.t6 VSUBS 1.81224f
C1106 VP.n1 VSUBS 0.075041f
C1107 VP.n2 VSUBS 0.039241f
C1108 VP.n3 VSUBS 0.060496f
C1109 VP.n4 VSUBS 0.039241f
C1110 VP.n5 VSUBS 0.031723f
C1111 VP.n6 VSUBS 0.039241f
C1112 VP.t2 VSUBS 1.81224f
C1113 VP.n7 VSUBS 0.677087f
C1114 VP.n8 VSUBS 0.039241f
C1115 VP.n9 VSUBS 0.044749f
C1116 VP.n10 VSUBS 0.039241f
C1117 VP.t3 VSUBS 1.81224f
C1118 VP.n11 VSUBS 0.811462f
C1119 VP.n12 VSUBS 0.051736f
C1120 VP.t4 VSUBS 1.81224f
C1121 VP.n13 VSUBS 0.075041f
C1122 VP.n14 VSUBS 0.039241f
C1123 VP.n15 VSUBS 0.060496f
C1124 VP.n16 VSUBS 0.039241f
C1125 VP.n17 VSUBS 0.031723f
C1126 VP.n18 VSUBS 0.039241f
C1127 VP.t5 VSUBS 1.81224f
C1128 VP.n19 VSUBS 0.797271f
C1129 VP.t1 VSUBS 2.2029f
C1130 VP.n20 VSUBS 0.769809f
C1131 VP.n21 VSUBS 0.421568f
C1132 VP.n22 VSUBS 0.049664f
C1133 VP.n23 VSUBS 0.073136f
C1134 VP.n24 VSUBS 0.077991f
C1135 VP.n25 VSUBS 0.039241f
C1136 VP.n26 VSUBS 0.039241f
C1137 VP.n27 VSUBS 0.039241f
C1138 VP.n28 VSUBS 0.077991f
C1139 VP.n29 VSUBS 0.073136f
C1140 VP.t0 VSUBS 1.81224f
C1141 VP.n30 VSUBS 0.677087f
C1142 VP.n31 VSUBS 0.049664f
C1143 VP.n32 VSUBS 0.039241f
C1144 VP.n33 VSUBS 0.039241f
C1145 VP.n34 VSUBS 0.039241f
C1146 VP.n35 VSUBS 0.073136f
C1147 VP.n36 VSUBS 0.067916f
C1148 VP.n37 VSUBS 0.044749f
C1149 VP.n38 VSUBS 0.039241f
C1150 VP.n39 VSUBS 0.039241f
C1151 VP.n40 VSUBS 0.039241f
C1152 VP.n41 VSUBS 0.073136f
C1153 VP.n42 VSUBS 0.038832f
C1154 VP.n43 VSUBS 0.811462f
C1155 VP.n44 VSUBS 2.07928f
C1156 VP.n45 VSUBS 2.10858f
C1157 VP.n46 VSUBS 0.051736f
C1158 VP.n47 VSUBS 0.038832f
C1159 VP.n48 VSUBS 0.073136f
C1160 VP.n49 VSUBS 0.075041f
C1161 VP.n50 VSUBS 0.039241f
C1162 VP.n51 VSUBS 0.039241f
C1163 VP.n52 VSUBS 0.039241f
C1164 VP.n53 VSUBS 0.067916f
C1165 VP.n54 VSUBS 0.073136f
C1166 VP.n55 VSUBS 0.060496f
C1167 VP.n56 VSUBS 0.039241f
C1168 VP.n57 VSUBS 0.039241f
C1169 VP.n58 VSUBS 0.049664f
C1170 VP.n59 VSUBS 0.073136f
C1171 VP.n60 VSUBS 0.077991f
C1172 VP.n61 VSUBS 0.039241f
C1173 VP.n62 VSUBS 0.039241f
C1174 VP.n63 VSUBS 0.039241f
C1175 VP.n64 VSUBS 0.077991f
C1176 VP.n65 VSUBS 0.073136f
C1177 VP.t7 VSUBS 1.81224f
C1178 VP.n66 VSUBS 0.677087f
C1179 VP.n67 VSUBS 0.049664f
C1180 VP.n68 VSUBS 0.039241f
C1181 VP.n69 VSUBS 0.039241f
C1182 VP.n70 VSUBS 0.039241f
C1183 VP.n71 VSUBS 0.073136f
C1184 VP.n72 VSUBS 0.067916f
C1185 VP.n73 VSUBS 0.044749f
C1186 VP.n74 VSUBS 0.039241f
C1187 VP.n75 VSUBS 0.039241f
C1188 VP.n76 VSUBS 0.039241f
C1189 VP.n77 VSUBS 0.073136f
C1190 VP.n78 VSUBS 0.038832f
C1191 VP.n79 VSUBS 0.811462f
C1192 VP.n80 VSUBS 0.078143f
.ends

