* NGSPICE file created from diff_pair_sample_1790.ext - technology: sky130A

.subckt diff_pair_sample_1790 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t1 w_n2220_n1258# sky130_fd_pr__pfet_01v8 ad=0.5655 pd=3.68 as=0.23925 ps=1.78 w=1.45 l=0.92
X1 B.t11 B.t9 B.t10 w_n2220_n1258# sky130_fd_pr__pfet_01v8 ad=0.5655 pd=3.68 as=0 ps=0 w=1.45 l=0.92
X2 VDD1.t7 VP.t0 VTAIL.t3 w_n2220_n1258# sky130_fd_pr__pfet_01v8 ad=0.23925 pd=1.78 as=0.23925 ps=1.78 w=1.45 l=0.92
X3 VDD1.t6 VP.t1 VTAIL.t7 w_n2220_n1258# sky130_fd_pr__pfet_01v8 ad=0.23925 pd=1.78 as=0.23925 ps=1.78 w=1.45 l=0.92
X4 VTAIL.t4 VP.t2 VDD1.t5 w_n2220_n1258# sky130_fd_pr__pfet_01v8 ad=0.5655 pd=3.68 as=0.23925 ps=1.78 w=1.45 l=0.92
X5 B.t8 B.t6 B.t7 w_n2220_n1258# sky130_fd_pr__pfet_01v8 ad=0.5655 pd=3.68 as=0 ps=0 w=1.45 l=0.92
X6 VDD1.t4 VP.t3 VTAIL.t5 w_n2220_n1258# sky130_fd_pr__pfet_01v8 ad=0.23925 pd=1.78 as=0.5655 ps=3.68 w=1.45 l=0.92
X7 VTAIL.t6 VP.t4 VDD1.t3 w_n2220_n1258# sky130_fd_pr__pfet_01v8 ad=0.23925 pd=1.78 as=0.23925 ps=1.78 w=1.45 l=0.92
X8 VTAIL.t14 VN.t1 VDD2.t7 w_n2220_n1258# sky130_fd_pr__pfet_01v8 ad=0.23925 pd=1.78 as=0.23925 ps=1.78 w=1.45 l=0.92
X9 B.t5 B.t3 B.t4 w_n2220_n1258# sky130_fd_pr__pfet_01v8 ad=0.5655 pd=3.68 as=0 ps=0 w=1.45 l=0.92
X10 VDD2.t5 VN.t2 VTAIL.t13 w_n2220_n1258# sky130_fd_pr__pfet_01v8 ad=0.23925 pd=1.78 as=0.5655 ps=3.68 w=1.45 l=0.92
X11 VTAIL.t2 VP.t5 VDD1.t2 w_n2220_n1258# sky130_fd_pr__pfet_01v8 ad=0.23925 pd=1.78 as=0.23925 ps=1.78 w=1.45 l=0.92
X12 VDD2.t4 VN.t3 VTAIL.t12 w_n2220_n1258# sky130_fd_pr__pfet_01v8 ad=0.23925 pd=1.78 as=0.5655 ps=3.68 w=1.45 l=0.92
X13 VDD1.t1 VP.t6 VTAIL.t0 w_n2220_n1258# sky130_fd_pr__pfet_01v8 ad=0.23925 pd=1.78 as=0.5655 ps=3.68 w=1.45 l=0.92
X14 VTAIL.t11 VN.t4 VDD2.t3 w_n2220_n1258# sky130_fd_pr__pfet_01v8 ad=0.23925 pd=1.78 as=0.23925 ps=1.78 w=1.45 l=0.92
X15 VDD2.t2 VN.t5 VTAIL.t10 w_n2220_n1258# sky130_fd_pr__pfet_01v8 ad=0.23925 pd=1.78 as=0.23925 ps=1.78 w=1.45 l=0.92
X16 VTAIL.t9 VN.t6 VDD2.t0 w_n2220_n1258# sky130_fd_pr__pfet_01v8 ad=0.5655 pd=3.68 as=0.23925 ps=1.78 w=1.45 l=0.92
X17 B.t2 B.t0 B.t1 w_n2220_n1258# sky130_fd_pr__pfet_01v8 ad=0.5655 pd=3.68 as=0 ps=0 w=1.45 l=0.92
X18 VTAIL.t1 VP.t7 VDD1.t0 w_n2220_n1258# sky130_fd_pr__pfet_01v8 ad=0.5655 pd=3.68 as=0.23925 ps=1.78 w=1.45 l=0.92
X19 VDD2.t6 VN.t7 VTAIL.t8 w_n2220_n1258# sky130_fd_pr__pfet_01v8 ad=0.23925 pd=1.78 as=0.23925 ps=1.78 w=1.45 l=0.92
R0 VN.n23 VN.n13 161.3
R1 VN.n21 VN.n20 161.3
R2 VN.n19 VN.n14 161.3
R3 VN.n18 VN.n17 161.3
R4 VN.n10 VN.n0 161.3
R5 VN.n8 VN.n7 161.3
R6 VN.n6 VN.n1 161.3
R7 VN.n5 VN.n4 161.3
R8 VN.n2 VN.t6 95.3244
R9 VN.n15 VN.t2 95.3244
R10 VN.n11 VN.t3 80.9451
R11 VN.n24 VN.t0 80.9451
R12 VN.n25 VN.n24 80.6037
R13 VN.n12 VN.n11 80.6037
R14 VN.n11 VN.n10 52.3599
R15 VN.n24 VN.n23 52.3599
R16 VN.n3 VN.n2 47.0243
R17 VN.n16 VN.n15 47.0243
R18 VN.n18 VN.n15 44.4862
R19 VN.n5 VN.n2 44.4862
R20 VN.n4 VN.n1 40.4934
R21 VN.n8 VN.n1 40.4934
R22 VN.n17 VN.n14 40.4934
R23 VN.n21 VN.n14 40.4934
R24 VN.n3 VN.t5 37.9842
R25 VN.n9 VN.t1 37.9842
R26 VN.n16 VN.t4 37.9842
R27 VN.n22 VN.t7 37.9842
R28 VN VN.n25 35.4309
R29 VN.n10 VN.n9 18.3508
R30 VN.n23 VN.n22 18.3508
R31 VN.n4 VN.n3 6.11725
R32 VN.n9 VN.n8 6.11725
R33 VN.n17 VN.n16 6.11725
R34 VN.n22 VN.n21 6.11725
R35 VN.n25 VN.n13 0.285035
R36 VN.n12 VN.n0 0.285035
R37 VN.n20 VN.n13 0.189894
R38 VN.n20 VN.n19 0.189894
R39 VN.n19 VN.n18 0.189894
R40 VN.n6 VN.n5 0.189894
R41 VN.n7 VN.n6 0.189894
R42 VN.n7 VN.n0 0.189894
R43 VN VN.n12 0.146778
R44 VDD2.n2 VDD2.n1 250.466
R45 VDD2.n2 VDD2.n0 250.466
R46 VDD2 VDD2.n5 250.464
R47 VDD2.n4 VDD2.n3 249.982
R48 VDD2.n4 VDD2.n2 29.8144
R49 VDD2.n5 VDD2.t3 22.4177
R50 VDD2.n5 VDD2.t5 22.4177
R51 VDD2.n3 VDD2.t1 22.4177
R52 VDD2.n3 VDD2.t6 22.4177
R53 VDD2.n1 VDD2.t7 22.4177
R54 VDD2.n1 VDD2.t4 22.4177
R55 VDD2.n0 VDD2.t0 22.4177
R56 VDD2.n0 VDD2.t2 22.4177
R57 VDD2 VDD2.n4 0.597483
R58 VTAIL.n11 VTAIL.t1 255.721
R59 VTAIL.n10 VTAIL.t13 255.721
R60 VTAIL.n7 VTAIL.t15 255.721
R61 VTAIL.n15 VTAIL.t12 255.721
R62 VTAIL.n2 VTAIL.t9 255.721
R63 VTAIL.n3 VTAIL.t5 255.721
R64 VTAIL.n6 VTAIL.t4 255.721
R65 VTAIL.n14 VTAIL.t0 255.721
R66 VTAIL.n13 VTAIL.n12 233.304
R67 VTAIL.n9 VTAIL.n8 233.304
R68 VTAIL.n1 VTAIL.n0 233.304
R69 VTAIL.n5 VTAIL.n4 233.304
R70 VTAIL.n0 VTAIL.t10 22.4177
R71 VTAIL.n0 VTAIL.t14 22.4177
R72 VTAIL.n4 VTAIL.t7 22.4177
R73 VTAIL.n4 VTAIL.t6 22.4177
R74 VTAIL.n12 VTAIL.t3 22.4177
R75 VTAIL.n12 VTAIL.t2 22.4177
R76 VTAIL.n8 VTAIL.t8 22.4177
R77 VTAIL.n8 VTAIL.t11 22.4177
R78 VTAIL.n15 VTAIL.n14 14.6945
R79 VTAIL.n7 VTAIL.n6 14.6945
R80 VTAIL.n9 VTAIL.n7 1.07809
R81 VTAIL.n10 VTAIL.n9 1.07809
R82 VTAIL.n13 VTAIL.n11 1.07809
R83 VTAIL.n14 VTAIL.n13 1.07809
R84 VTAIL.n6 VTAIL.n5 1.07809
R85 VTAIL.n5 VTAIL.n3 1.07809
R86 VTAIL.n2 VTAIL.n1 1.07809
R87 VTAIL VTAIL.n15 1.0199
R88 VTAIL.n11 VTAIL.n10 0.470328
R89 VTAIL.n3 VTAIL.n2 0.470328
R90 VTAIL VTAIL.n1 0.0586897
R91 B.n180 B.n179 585
R92 B.n178 B.n63 585
R93 B.n177 B.n176 585
R94 B.n175 B.n64 585
R95 B.n174 B.n173 585
R96 B.n172 B.n65 585
R97 B.n171 B.n170 585
R98 B.n169 B.n66 585
R99 B.n168 B.n167 585
R100 B.n166 B.n67 585
R101 B.n165 B.n164 585
R102 B.n162 B.n68 585
R103 B.n161 B.n160 585
R104 B.n159 B.n71 585
R105 B.n158 B.n157 585
R106 B.n156 B.n72 585
R107 B.n155 B.n154 585
R108 B.n153 B.n73 585
R109 B.n152 B.n151 585
R110 B.n150 B.n74 585
R111 B.n148 B.n147 585
R112 B.n146 B.n77 585
R113 B.n145 B.n144 585
R114 B.n143 B.n78 585
R115 B.n142 B.n141 585
R116 B.n140 B.n79 585
R117 B.n139 B.n138 585
R118 B.n137 B.n80 585
R119 B.n136 B.n135 585
R120 B.n134 B.n81 585
R121 B.n133 B.n132 585
R122 B.n181 B.n62 585
R123 B.n183 B.n182 585
R124 B.n184 B.n61 585
R125 B.n186 B.n185 585
R126 B.n187 B.n60 585
R127 B.n189 B.n188 585
R128 B.n190 B.n59 585
R129 B.n192 B.n191 585
R130 B.n193 B.n58 585
R131 B.n195 B.n194 585
R132 B.n196 B.n57 585
R133 B.n198 B.n197 585
R134 B.n199 B.n56 585
R135 B.n201 B.n200 585
R136 B.n202 B.n55 585
R137 B.n204 B.n203 585
R138 B.n205 B.n54 585
R139 B.n207 B.n206 585
R140 B.n208 B.n53 585
R141 B.n210 B.n209 585
R142 B.n211 B.n52 585
R143 B.n213 B.n212 585
R144 B.n214 B.n51 585
R145 B.n216 B.n215 585
R146 B.n217 B.n50 585
R147 B.n219 B.n218 585
R148 B.n220 B.n49 585
R149 B.n222 B.n221 585
R150 B.n223 B.n48 585
R151 B.n225 B.n224 585
R152 B.n226 B.n47 585
R153 B.n228 B.n227 585
R154 B.n229 B.n46 585
R155 B.n231 B.n230 585
R156 B.n232 B.n45 585
R157 B.n234 B.n233 585
R158 B.n235 B.n44 585
R159 B.n237 B.n236 585
R160 B.n238 B.n43 585
R161 B.n240 B.n239 585
R162 B.n241 B.n42 585
R163 B.n243 B.n242 585
R164 B.n244 B.n41 585
R165 B.n246 B.n245 585
R166 B.n247 B.n40 585
R167 B.n249 B.n248 585
R168 B.n250 B.n39 585
R169 B.n252 B.n251 585
R170 B.n253 B.n38 585
R171 B.n255 B.n254 585
R172 B.n256 B.n37 585
R173 B.n258 B.n257 585
R174 B.n259 B.n36 585
R175 B.n261 B.n260 585
R176 B.n308 B.n15 585
R177 B.n307 B.n306 585
R178 B.n305 B.n16 585
R179 B.n304 B.n303 585
R180 B.n302 B.n17 585
R181 B.n301 B.n300 585
R182 B.n299 B.n18 585
R183 B.n298 B.n297 585
R184 B.n296 B.n19 585
R185 B.n295 B.n294 585
R186 B.n293 B.n20 585
R187 B.n292 B.n291 585
R188 B.n290 B.n21 585
R189 B.n289 B.n288 585
R190 B.n287 B.n25 585
R191 B.n286 B.n285 585
R192 B.n284 B.n26 585
R193 B.n283 B.n282 585
R194 B.n281 B.n27 585
R195 B.n280 B.n279 585
R196 B.n277 B.n28 585
R197 B.n276 B.n275 585
R198 B.n274 B.n31 585
R199 B.n273 B.n272 585
R200 B.n271 B.n32 585
R201 B.n270 B.n269 585
R202 B.n268 B.n33 585
R203 B.n267 B.n266 585
R204 B.n265 B.n34 585
R205 B.n264 B.n263 585
R206 B.n262 B.n35 585
R207 B.n310 B.n309 585
R208 B.n311 B.n14 585
R209 B.n313 B.n312 585
R210 B.n314 B.n13 585
R211 B.n316 B.n315 585
R212 B.n317 B.n12 585
R213 B.n319 B.n318 585
R214 B.n320 B.n11 585
R215 B.n322 B.n321 585
R216 B.n323 B.n10 585
R217 B.n325 B.n324 585
R218 B.n326 B.n9 585
R219 B.n328 B.n327 585
R220 B.n329 B.n8 585
R221 B.n331 B.n330 585
R222 B.n332 B.n7 585
R223 B.n334 B.n333 585
R224 B.n335 B.n6 585
R225 B.n337 B.n336 585
R226 B.n338 B.n5 585
R227 B.n340 B.n339 585
R228 B.n341 B.n4 585
R229 B.n343 B.n342 585
R230 B.n344 B.n3 585
R231 B.n346 B.n345 585
R232 B.n347 B.n0 585
R233 B.n2 B.n1 585
R234 B.n95 B.n94 585
R235 B.n97 B.n96 585
R236 B.n98 B.n93 585
R237 B.n100 B.n99 585
R238 B.n101 B.n92 585
R239 B.n103 B.n102 585
R240 B.n104 B.n91 585
R241 B.n106 B.n105 585
R242 B.n107 B.n90 585
R243 B.n109 B.n108 585
R244 B.n110 B.n89 585
R245 B.n112 B.n111 585
R246 B.n113 B.n88 585
R247 B.n115 B.n114 585
R248 B.n116 B.n87 585
R249 B.n118 B.n117 585
R250 B.n119 B.n86 585
R251 B.n121 B.n120 585
R252 B.n122 B.n85 585
R253 B.n124 B.n123 585
R254 B.n125 B.n84 585
R255 B.n127 B.n126 585
R256 B.n128 B.n83 585
R257 B.n130 B.n129 585
R258 B.n131 B.n82 585
R259 B.n133 B.n82 478.086
R260 B.n179 B.n62 478.086
R261 B.n262 B.n261 478.086
R262 B.n310 B.n15 478.086
R263 B.n69 B.t1 273.467
R264 B.n29 B.t8 273.467
R265 B.n75 B.t4 273.467
R266 B.n22 B.t11 273.467
R267 B.n349 B.n348 256.663
R268 B.n70 B.t2 249.226
R269 B.n30 B.t7 249.226
R270 B.n76 B.t5 249.225
R271 B.n23 B.t10 249.225
R272 B.n75 B.t3 240.334
R273 B.n69 B.t0 240.334
R274 B.n29 B.t6 240.334
R275 B.n22 B.t9 240.334
R276 B.n348 B.n347 235.042
R277 B.n348 B.n2 235.042
R278 B.n134 B.n133 163.367
R279 B.n135 B.n134 163.367
R280 B.n135 B.n80 163.367
R281 B.n139 B.n80 163.367
R282 B.n140 B.n139 163.367
R283 B.n141 B.n140 163.367
R284 B.n141 B.n78 163.367
R285 B.n145 B.n78 163.367
R286 B.n146 B.n145 163.367
R287 B.n147 B.n146 163.367
R288 B.n147 B.n74 163.367
R289 B.n152 B.n74 163.367
R290 B.n153 B.n152 163.367
R291 B.n154 B.n153 163.367
R292 B.n154 B.n72 163.367
R293 B.n158 B.n72 163.367
R294 B.n159 B.n158 163.367
R295 B.n160 B.n159 163.367
R296 B.n160 B.n68 163.367
R297 B.n165 B.n68 163.367
R298 B.n166 B.n165 163.367
R299 B.n167 B.n166 163.367
R300 B.n167 B.n66 163.367
R301 B.n171 B.n66 163.367
R302 B.n172 B.n171 163.367
R303 B.n173 B.n172 163.367
R304 B.n173 B.n64 163.367
R305 B.n177 B.n64 163.367
R306 B.n178 B.n177 163.367
R307 B.n179 B.n178 163.367
R308 B.n261 B.n36 163.367
R309 B.n257 B.n36 163.367
R310 B.n257 B.n256 163.367
R311 B.n256 B.n255 163.367
R312 B.n255 B.n38 163.367
R313 B.n251 B.n38 163.367
R314 B.n251 B.n250 163.367
R315 B.n250 B.n249 163.367
R316 B.n249 B.n40 163.367
R317 B.n245 B.n40 163.367
R318 B.n245 B.n244 163.367
R319 B.n244 B.n243 163.367
R320 B.n243 B.n42 163.367
R321 B.n239 B.n42 163.367
R322 B.n239 B.n238 163.367
R323 B.n238 B.n237 163.367
R324 B.n237 B.n44 163.367
R325 B.n233 B.n44 163.367
R326 B.n233 B.n232 163.367
R327 B.n232 B.n231 163.367
R328 B.n231 B.n46 163.367
R329 B.n227 B.n46 163.367
R330 B.n227 B.n226 163.367
R331 B.n226 B.n225 163.367
R332 B.n225 B.n48 163.367
R333 B.n221 B.n48 163.367
R334 B.n221 B.n220 163.367
R335 B.n220 B.n219 163.367
R336 B.n219 B.n50 163.367
R337 B.n215 B.n50 163.367
R338 B.n215 B.n214 163.367
R339 B.n214 B.n213 163.367
R340 B.n213 B.n52 163.367
R341 B.n209 B.n52 163.367
R342 B.n209 B.n208 163.367
R343 B.n208 B.n207 163.367
R344 B.n207 B.n54 163.367
R345 B.n203 B.n54 163.367
R346 B.n203 B.n202 163.367
R347 B.n202 B.n201 163.367
R348 B.n201 B.n56 163.367
R349 B.n197 B.n56 163.367
R350 B.n197 B.n196 163.367
R351 B.n196 B.n195 163.367
R352 B.n195 B.n58 163.367
R353 B.n191 B.n58 163.367
R354 B.n191 B.n190 163.367
R355 B.n190 B.n189 163.367
R356 B.n189 B.n60 163.367
R357 B.n185 B.n60 163.367
R358 B.n185 B.n184 163.367
R359 B.n184 B.n183 163.367
R360 B.n183 B.n62 163.367
R361 B.n306 B.n15 163.367
R362 B.n306 B.n305 163.367
R363 B.n305 B.n304 163.367
R364 B.n304 B.n17 163.367
R365 B.n300 B.n17 163.367
R366 B.n300 B.n299 163.367
R367 B.n299 B.n298 163.367
R368 B.n298 B.n19 163.367
R369 B.n294 B.n19 163.367
R370 B.n294 B.n293 163.367
R371 B.n293 B.n292 163.367
R372 B.n292 B.n21 163.367
R373 B.n288 B.n21 163.367
R374 B.n288 B.n287 163.367
R375 B.n287 B.n286 163.367
R376 B.n286 B.n26 163.367
R377 B.n282 B.n26 163.367
R378 B.n282 B.n281 163.367
R379 B.n281 B.n280 163.367
R380 B.n280 B.n28 163.367
R381 B.n275 B.n28 163.367
R382 B.n275 B.n274 163.367
R383 B.n274 B.n273 163.367
R384 B.n273 B.n32 163.367
R385 B.n269 B.n32 163.367
R386 B.n269 B.n268 163.367
R387 B.n268 B.n267 163.367
R388 B.n267 B.n34 163.367
R389 B.n263 B.n34 163.367
R390 B.n263 B.n262 163.367
R391 B.n311 B.n310 163.367
R392 B.n312 B.n311 163.367
R393 B.n312 B.n13 163.367
R394 B.n316 B.n13 163.367
R395 B.n317 B.n316 163.367
R396 B.n318 B.n317 163.367
R397 B.n318 B.n11 163.367
R398 B.n322 B.n11 163.367
R399 B.n323 B.n322 163.367
R400 B.n324 B.n323 163.367
R401 B.n324 B.n9 163.367
R402 B.n328 B.n9 163.367
R403 B.n329 B.n328 163.367
R404 B.n330 B.n329 163.367
R405 B.n330 B.n7 163.367
R406 B.n334 B.n7 163.367
R407 B.n335 B.n334 163.367
R408 B.n336 B.n335 163.367
R409 B.n336 B.n5 163.367
R410 B.n340 B.n5 163.367
R411 B.n341 B.n340 163.367
R412 B.n342 B.n341 163.367
R413 B.n342 B.n3 163.367
R414 B.n346 B.n3 163.367
R415 B.n347 B.n346 163.367
R416 B.n94 B.n2 163.367
R417 B.n97 B.n94 163.367
R418 B.n98 B.n97 163.367
R419 B.n99 B.n98 163.367
R420 B.n99 B.n92 163.367
R421 B.n103 B.n92 163.367
R422 B.n104 B.n103 163.367
R423 B.n105 B.n104 163.367
R424 B.n105 B.n90 163.367
R425 B.n109 B.n90 163.367
R426 B.n110 B.n109 163.367
R427 B.n111 B.n110 163.367
R428 B.n111 B.n88 163.367
R429 B.n115 B.n88 163.367
R430 B.n116 B.n115 163.367
R431 B.n117 B.n116 163.367
R432 B.n117 B.n86 163.367
R433 B.n121 B.n86 163.367
R434 B.n122 B.n121 163.367
R435 B.n123 B.n122 163.367
R436 B.n123 B.n84 163.367
R437 B.n127 B.n84 163.367
R438 B.n128 B.n127 163.367
R439 B.n129 B.n128 163.367
R440 B.n129 B.n82 163.367
R441 B.n149 B.n76 59.5399
R442 B.n163 B.n70 59.5399
R443 B.n278 B.n30 59.5399
R444 B.n24 B.n23 59.5399
R445 B.n309 B.n308 31.0639
R446 B.n260 B.n35 31.0639
R447 B.n181 B.n180 31.0639
R448 B.n132 B.n131 31.0639
R449 B.n76 B.n75 24.2429
R450 B.n70 B.n69 24.2429
R451 B.n30 B.n29 24.2429
R452 B.n23 B.n22 24.2429
R453 B B.n349 18.0485
R454 B.n309 B.n14 10.6151
R455 B.n313 B.n14 10.6151
R456 B.n314 B.n313 10.6151
R457 B.n315 B.n314 10.6151
R458 B.n315 B.n12 10.6151
R459 B.n319 B.n12 10.6151
R460 B.n320 B.n319 10.6151
R461 B.n321 B.n320 10.6151
R462 B.n321 B.n10 10.6151
R463 B.n325 B.n10 10.6151
R464 B.n326 B.n325 10.6151
R465 B.n327 B.n326 10.6151
R466 B.n327 B.n8 10.6151
R467 B.n331 B.n8 10.6151
R468 B.n332 B.n331 10.6151
R469 B.n333 B.n332 10.6151
R470 B.n333 B.n6 10.6151
R471 B.n337 B.n6 10.6151
R472 B.n338 B.n337 10.6151
R473 B.n339 B.n338 10.6151
R474 B.n339 B.n4 10.6151
R475 B.n343 B.n4 10.6151
R476 B.n344 B.n343 10.6151
R477 B.n345 B.n344 10.6151
R478 B.n345 B.n0 10.6151
R479 B.n308 B.n307 10.6151
R480 B.n307 B.n16 10.6151
R481 B.n303 B.n16 10.6151
R482 B.n303 B.n302 10.6151
R483 B.n302 B.n301 10.6151
R484 B.n301 B.n18 10.6151
R485 B.n297 B.n18 10.6151
R486 B.n297 B.n296 10.6151
R487 B.n296 B.n295 10.6151
R488 B.n295 B.n20 10.6151
R489 B.n291 B.n290 10.6151
R490 B.n290 B.n289 10.6151
R491 B.n289 B.n25 10.6151
R492 B.n285 B.n25 10.6151
R493 B.n285 B.n284 10.6151
R494 B.n284 B.n283 10.6151
R495 B.n283 B.n27 10.6151
R496 B.n279 B.n27 10.6151
R497 B.n277 B.n276 10.6151
R498 B.n276 B.n31 10.6151
R499 B.n272 B.n31 10.6151
R500 B.n272 B.n271 10.6151
R501 B.n271 B.n270 10.6151
R502 B.n270 B.n33 10.6151
R503 B.n266 B.n33 10.6151
R504 B.n266 B.n265 10.6151
R505 B.n265 B.n264 10.6151
R506 B.n264 B.n35 10.6151
R507 B.n260 B.n259 10.6151
R508 B.n259 B.n258 10.6151
R509 B.n258 B.n37 10.6151
R510 B.n254 B.n37 10.6151
R511 B.n254 B.n253 10.6151
R512 B.n253 B.n252 10.6151
R513 B.n252 B.n39 10.6151
R514 B.n248 B.n39 10.6151
R515 B.n248 B.n247 10.6151
R516 B.n247 B.n246 10.6151
R517 B.n246 B.n41 10.6151
R518 B.n242 B.n41 10.6151
R519 B.n242 B.n241 10.6151
R520 B.n241 B.n240 10.6151
R521 B.n240 B.n43 10.6151
R522 B.n236 B.n43 10.6151
R523 B.n236 B.n235 10.6151
R524 B.n235 B.n234 10.6151
R525 B.n234 B.n45 10.6151
R526 B.n230 B.n45 10.6151
R527 B.n230 B.n229 10.6151
R528 B.n229 B.n228 10.6151
R529 B.n228 B.n47 10.6151
R530 B.n224 B.n47 10.6151
R531 B.n224 B.n223 10.6151
R532 B.n223 B.n222 10.6151
R533 B.n222 B.n49 10.6151
R534 B.n218 B.n49 10.6151
R535 B.n218 B.n217 10.6151
R536 B.n217 B.n216 10.6151
R537 B.n216 B.n51 10.6151
R538 B.n212 B.n51 10.6151
R539 B.n212 B.n211 10.6151
R540 B.n211 B.n210 10.6151
R541 B.n210 B.n53 10.6151
R542 B.n206 B.n53 10.6151
R543 B.n206 B.n205 10.6151
R544 B.n205 B.n204 10.6151
R545 B.n204 B.n55 10.6151
R546 B.n200 B.n55 10.6151
R547 B.n200 B.n199 10.6151
R548 B.n199 B.n198 10.6151
R549 B.n198 B.n57 10.6151
R550 B.n194 B.n57 10.6151
R551 B.n194 B.n193 10.6151
R552 B.n193 B.n192 10.6151
R553 B.n192 B.n59 10.6151
R554 B.n188 B.n59 10.6151
R555 B.n188 B.n187 10.6151
R556 B.n187 B.n186 10.6151
R557 B.n186 B.n61 10.6151
R558 B.n182 B.n61 10.6151
R559 B.n182 B.n181 10.6151
R560 B.n95 B.n1 10.6151
R561 B.n96 B.n95 10.6151
R562 B.n96 B.n93 10.6151
R563 B.n100 B.n93 10.6151
R564 B.n101 B.n100 10.6151
R565 B.n102 B.n101 10.6151
R566 B.n102 B.n91 10.6151
R567 B.n106 B.n91 10.6151
R568 B.n107 B.n106 10.6151
R569 B.n108 B.n107 10.6151
R570 B.n108 B.n89 10.6151
R571 B.n112 B.n89 10.6151
R572 B.n113 B.n112 10.6151
R573 B.n114 B.n113 10.6151
R574 B.n114 B.n87 10.6151
R575 B.n118 B.n87 10.6151
R576 B.n119 B.n118 10.6151
R577 B.n120 B.n119 10.6151
R578 B.n120 B.n85 10.6151
R579 B.n124 B.n85 10.6151
R580 B.n125 B.n124 10.6151
R581 B.n126 B.n125 10.6151
R582 B.n126 B.n83 10.6151
R583 B.n130 B.n83 10.6151
R584 B.n131 B.n130 10.6151
R585 B.n132 B.n81 10.6151
R586 B.n136 B.n81 10.6151
R587 B.n137 B.n136 10.6151
R588 B.n138 B.n137 10.6151
R589 B.n138 B.n79 10.6151
R590 B.n142 B.n79 10.6151
R591 B.n143 B.n142 10.6151
R592 B.n144 B.n143 10.6151
R593 B.n144 B.n77 10.6151
R594 B.n148 B.n77 10.6151
R595 B.n151 B.n150 10.6151
R596 B.n151 B.n73 10.6151
R597 B.n155 B.n73 10.6151
R598 B.n156 B.n155 10.6151
R599 B.n157 B.n156 10.6151
R600 B.n157 B.n71 10.6151
R601 B.n161 B.n71 10.6151
R602 B.n162 B.n161 10.6151
R603 B.n164 B.n67 10.6151
R604 B.n168 B.n67 10.6151
R605 B.n169 B.n168 10.6151
R606 B.n170 B.n169 10.6151
R607 B.n170 B.n65 10.6151
R608 B.n174 B.n65 10.6151
R609 B.n175 B.n174 10.6151
R610 B.n176 B.n175 10.6151
R611 B.n176 B.n63 10.6151
R612 B.n180 B.n63 10.6151
R613 B.n349 B.n0 8.11757
R614 B.n349 B.n1 8.11757
R615 B.n291 B.n24 6.5566
R616 B.n279 B.n278 6.5566
R617 B.n150 B.n149 6.5566
R618 B.n163 B.n162 6.5566
R619 B.n24 B.n20 4.05904
R620 B.n278 B.n277 4.05904
R621 B.n149 B.n148 4.05904
R622 B.n164 B.n163 4.05904
R623 VP.n8 VP.n7 161.3
R624 VP.n9 VP.n4 161.3
R625 VP.n11 VP.n10 161.3
R626 VP.n13 VP.n3 161.3
R627 VP.n26 VP.n0 161.3
R628 VP.n24 VP.n23 161.3
R629 VP.n22 VP.n1 161.3
R630 VP.n21 VP.n20 161.3
R631 VP.n18 VP.n2 161.3
R632 VP.n5 VP.t7 95.3244
R633 VP.n17 VP.t2 80.9451
R634 VP.n27 VP.t3 80.9451
R635 VP.n14 VP.t6 80.9451
R636 VP.n15 VP.n14 80.6037
R637 VP.n28 VP.n27 80.6037
R638 VP.n17 VP.n16 80.6037
R639 VP.n18 VP.n17 52.3599
R640 VP.n27 VP.n26 52.3599
R641 VP.n14 VP.n13 52.3599
R642 VP.n6 VP.n5 47.0243
R643 VP.n8 VP.n5 44.4862
R644 VP.n20 VP.n1 40.4934
R645 VP.n24 VP.n1 40.4934
R646 VP.n11 VP.n4 40.4934
R647 VP.n7 VP.n4 40.4934
R648 VP.n19 VP.t1 37.9842
R649 VP.n25 VP.t4 37.9842
R650 VP.n12 VP.t5 37.9842
R651 VP.n6 VP.t0 37.9842
R652 VP.n16 VP.n15 35.1453
R653 VP.n19 VP.n18 18.3508
R654 VP.n26 VP.n25 18.3508
R655 VP.n13 VP.n12 18.3508
R656 VP.n20 VP.n19 6.11725
R657 VP.n25 VP.n24 6.11725
R658 VP.n12 VP.n11 6.11725
R659 VP.n7 VP.n6 6.11725
R660 VP.n15 VP.n3 0.285035
R661 VP.n16 VP.n2 0.285035
R662 VP.n28 VP.n0 0.285035
R663 VP.n9 VP.n8 0.189894
R664 VP.n10 VP.n9 0.189894
R665 VP.n10 VP.n3 0.189894
R666 VP.n21 VP.n2 0.189894
R667 VP.n22 VP.n21 0.189894
R668 VP.n23 VP.n22 0.189894
R669 VP.n23 VP.n0 0.189894
R670 VP VP.n28 0.146778
R671 VDD1 VDD1.n0 250.579
R672 VDD1.n3 VDD1.n2 250.466
R673 VDD1.n3 VDD1.n1 250.466
R674 VDD1.n5 VDD1.n4 249.982
R675 VDD1.n5 VDD1.n3 30.3974
R676 VDD1.n4 VDD1.t2 22.4177
R677 VDD1.n4 VDD1.t1 22.4177
R678 VDD1.n0 VDD1.t0 22.4177
R679 VDD1.n0 VDD1.t7 22.4177
R680 VDD1.n2 VDD1.t3 22.4177
R681 VDD1.n2 VDD1.t4 22.4177
R682 VDD1.n1 VDD1.t5 22.4177
R683 VDD1.n1 VDD1.t6 22.4177
R684 VDD1 VDD1.n5 0.481103
C0 B VDD2 0.895016f
C1 VN VDD2 1.10672f
C2 VDD2 VDD1 0.936073f
C3 VTAIL w_n2220_n1258# 1.51169f
C4 VTAIL VP 1.546f
C5 VTAIL B 0.998286f
C6 VN VTAIL 1.5319f
C7 VTAIL VDD1 3.24432f
C8 VTAIL VDD2 3.28747f
C9 w_n2220_n1258# VP 4.10807f
C10 w_n2220_n1258# B 4.58038f
C11 VN w_n2220_n1258# 3.83112f
C12 VP B 1.16117f
C13 VN VP 3.66588f
C14 w_n2220_n1258# VDD1 1.09558f
C15 VP VDD1 1.29828f
C16 VN B 0.696294f
C17 B VDD1 0.851308f
C18 VN VDD1 0.155208f
C19 w_n2220_n1258# VDD2 1.13865f
C20 VP VDD2 0.34846f
C21 VDD2 VSUBS 0.73142f
C22 VDD1 VSUBS 1.055482f
C23 VTAIL VSUBS 0.309983f
C24 VN VSUBS 3.8668f
C25 VP VSUBS 1.36414f
C26 B VSUBS 2.120506f
C27 w_n2220_n1258# VSUBS 35.830803f
C28 VDD1.t0 VSUBS 0.020468f
C29 VDD1.t7 VSUBS 0.020468f
C30 VDD1.n0 VSUBS 0.078611f
C31 VDD1.t5 VSUBS 0.020468f
C32 VDD1.t6 VSUBS 0.020468f
C33 VDD1.n1 VSUBS 0.07848f
C34 VDD1.t3 VSUBS 0.020468f
C35 VDD1.t4 VSUBS 0.020468f
C36 VDD1.n2 VSUBS 0.07848f
C37 VDD1.n3 VSUBS 1.27115f
C38 VDD1.t2 VSUBS 0.020468f
C39 VDD1.t1 VSUBS 0.020468f
C40 VDD1.n4 VSUBS 0.077978f
C41 VDD1.n5 VSUBS 1.12435f
C42 VP.n0 VSUBS 0.074536f
C43 VP.t4 VSUBS 0.16082f
C44 VP.n1 VSUBS 0.045156f
C45 VP.n2 VSUBS 0.074536f
C46 VP.t1 VSUBS 0.16082f
C47 VP.n3 VSUBS 0.074536f
C48 VP.t6 VSUBS 0.23955f
C49 VP.t5 VSUBS 0.16082f
C50 VP.n4 VSUBS 0.045156f
C51 VP.t7 VSUBS 0.269109f
C52 VP.n5 VSUBS 0.193313f
C53 VP.t0 VSUBS 0.16082f
C54 VP.n6 VSUBS 0.161913f
C55 VP.n7 VSUBS 0.072467f
C56 VP.n8 VSUBS 0.228204f
C57 VP.n9 VSUBS 0.055858f
C58 VP.n10 VSUBS 0.055858f
C59 VP.n11 VSUBS 0.072467f
C60 VP.n12 VSUBS 0.121001f
C61 VP.n13 VSUBS 0.067094f
C62 VP.n14 VSUBS 0.195605f
C63 VP.n15 VSUBS 1.69766f
C64 VP.n16 VSUBS 1.75479f
C65 VP.t2 VSUBS 0.23955f
C66 VP.n17 VSUBS 0.195605f
C67 VP.n18 VSUBS 0.067094f
C68 VP.n19 VSUBS 0.121001f
C69 VP.n20 VSUBS 0.072467f
C70 VP.n21 VSUBS 0.055858f
C71 VP.n22 VSUBS 0.055858f
C72 VP.n23 VSUBS 0.055858f
C73 VP.n24 VSUBS 0.072467f
C74 VP.n25 VSUBS 0.121001f
C75 VP.n26 VSUBS 0.067094f
C76 VP.t3 VSUBS 0.23955f
C77 VP.n27 VSUBS 0.195605f
C78 VP.n28 VSUBS 0.052314f
C79 B.n0 VSUBS 0.008183f
C80 B.n1 VSUBS 0.008183f
C81 B.n2 VSUBS 0.012102f
C82 B.n3 VSUBS 0.009274f
C83 B.n4 VSUBS 0.009274f
C84 B.n5 VSUBS 0.009274f
C85 B.n6 VSUBS 0.009274f
C86 B.n7 VSUBS 0.009274f
C87 B.n8 VSUBS 0.009274f
C88 B.n9 VSUBS 0.009274f
C89 B.n10 VSUBS 0.009274f
C90 B.n11 VSUBS 0.009274f
C91 B.n12 VSUBS 0.009274f
C92 B.n13 VSUBS 0.009274f
C93 B.n14 VSUBS 0.009274f
C94 B.n15 VSUBS 0.021663f
C95 B.n16 VSUBS 0.009274f
C96 B.n17 VSUBS 0.009274f
C97 B.n18 VSUBS 0.009274f
C98 B.n19 VSUBS 0.009274f
C99 B.n20 VSUBS 0.00641f
C100 B.n21 VSUBS 0.009274f
C101 B.t10 VSUBS 0.038842f
C102 B.t11 VSUBS 0.042971f
C103 B.t9 VSUBS 0.087264f
C104 B.n22 VSUBS 0.064905f
C105 B.n23 VSUBS 0.059812f
C106 B.n24 VSUBS 0.021487f
C107 B.n25 VSUBS 0.009274f
C108 B.n26 VSUBS 0.009274f
C109 B.n27 VSUBS 0.009274f
C110 B.n28 VSUBS 0.009274f
C111 B.t7 VSUBS 0.038842f
C112 B.t8 VSUBS 0.042971f
C113 B.t6 VSUBS 0.087264f
C114 B.n29 VSUBS 0.064905f
C115 B.n30 VSUBS 0.059812f
C116 B.n31 VSUBS 0.009274f
C117 B.n32 VSUBS 0.009274f
C118 B.n33 VSUBS 0.009274f
C119 B.n34 VSUBS 0.009274f
C120 B.n35 VSUBS 0.021663f
C121 B.n36 VSUBS 0.009274f
C122 B.n37 VSUBS 0.009274f
C123 B.n38 VSUBS 0.009274f
C124 B.n39 VSUBS 0.009274f
C125 B.n40 VSUBS 0.009274f
C126 B.n41 VSUBS 0.009274f
C127 B.n42 VSUBS 0.009274f
C128 B.n43 VSUBS 0.009274f
C129 B.n44 VSUBS 0.009274f
C130 B.n45 VSUBS 0.009274f
C131 B.n46 VSUBS 0.009274f
C132 B.n47 VSUBS 0.009274f
C133 B.n48 VSUBS 0.009274f
C134 B.n49 VSUBS 0.009274f
C135 B.n50 VSUBS 0.009274f
C136 B.n51 VSUBS 0.009274f
C137 B.n52 VSUBS 0.009274f
C138 B.n53 VSUBS 0.009274f
C139 B.n54 VSUBS 0.009274f
C140 B.n55 VSUBS 0.009274f
C141 B.n56 VSUBS 0.009274f
C142 B.n57 VSUBS 0.009274f
C143 B.n58 VSUBS 0.009274f
C144 B.n59 VSUBS 0.009274f
C145 B.n60 VSUBS 0.009274f
C146 B.n61 VSUBS 0.009274f
C147 B.n62 VSUBS 0.020342f
C148 B.n63 VSUBS 0.009274f
C149 B.n64 VSUBS 0.009274f
C150 B.n65 VSUBS 0.009274f
C151 B.n66 VSUBS 0.009274f
C152 B.n67 VSUBS 0.009274f
C153 B.n68 VSUBS 0.009274f
C154 B.t2 VSUBS 0.038842f
C155 B.t1 VSUBS 0.042971f
C156 B.t0 VSUBS 0.087264f
C157 B.n69 VSUBS 0.064905f
C158 B.n70 VSUBS 0.059812f
C159 B.n71 VSUBS 0.009274f
C160 B.n72 VSUBS 0.009274f
C161 B.n73 VSUBS 0.009274f
C162 B.n74 VSUBS 0.009274f
C163 B.t5 VSUBS 0.038842f
C164 B.t4 VSUBS 0.042971f
C165 B.t3 VSUBS 0.087264f
C166 B.n75 VSUBS 0.064905f
C167 B.n76 VSUBS 0.059812f
C168 B.n77 VSUBS 0.009274f
C169 B.n78 VSUBS 0.009274f
C170 B.n79 VSUBS 0.009274f
C171 B.n80 VSUBS 0.009274f
C172 B.n81 VSUBS 0.009274f
C173 B.n82 VSUBS 0.020342f
C174 B.n83 VSUBS 0.009274f
C175 B.n84 VSUBS 0.009274f
C176 B.n85 VSUBS 0.009274f
C177 B.n86 VSUBS 0.009274f
C178 B.n87 VSUBS 0.009274f
C179 B.n88 VSUBS 0.009274f
C180 B.n89 VSUBS 0.009274f
C181 B.n90 VSUBS 0.009274f
C182 B.n91 VSUBS 0.009274f
C183 B.n92 VSUBS 0.009274f
C184 B.n93 VSUBS 0.009274f
C185 B.n94 VSUBS 0.009274f
C186 B.n95 VSUBS 0.009274f
C187 B.n96 VSUBS 0.009274f
C188 B.n97 VSUBS 0.009274f
C189 B.n98 VSUBS 0.009274f
C190 B.n99 VSUBS 0.009274f
C191 B.n100 VSUBS 0.009274f
C192 B.n101 VSUBS 0.009274f
C193 B.n102 VSUBS 0.009274f
C194 B.n103 VSUBS 0.009274f
C195 B.n104 VSUBS 0.009274f
C196 B.n105 VSUBS 0.009274f
C197 B.n106 VSUBS 0.009274f
C198 B.n107 VSUBS 0.009274f
C199 B.n108 VSUBS 0.009274f
C200 B.n109 VSUBS 0.009274f
C201 B.n110 VSUBS 0.009274f
C202 B.n111 VSUBS 0.009274f
C203 B.n112 VSUBS 0.009274f
C204 B.n113 VSUBS 0.009274f
C205 B.n114 VSUBS 0.009274f
C206 B.n115 VSUBS 0.009274f
C207 B.n116 VSUBS 0.009274f
C208 B.n117 VSUBS 0.009274f
C209 B.n118 VSUBS 0.009274f
C210 B.n119 VSUBS 0.009274f
C211 B.n120 VSUBS 0.009274f
C212 B.n121 VSUBS 0.009274f
C213 B.n122 VSUBS 0.009274f
C214 B.n123 VSUBS 0.009274f
C215 B.n124 VSUBS 0.009274f
C216 B.n125 VSUBS 0.009274f
C217 B.n126 VSUBS 0.009274f
C218 B.n127 VSUBS 0.009274f
C219 B.n128 VSUBS 0.009274f
C220 B.n129 VSUBS 0.009274f
C221 B.n130 VSUBS 0.009274f
C222 B.n131 VSUBS 0.020342f
C223 B.n132 VSUBS 0.021663f
C224 B.n133 VSUBS 0.021663f
C225 B.n134 VSUBS 0.009274f
C226 B.n135 VSUBS 0.009274f
C227 B.n136 VSUBS 0.009274f
C228 B.n137 VSUBS 0.009274f
C229 B.n138 VSUBS 0.009274f
C230 B.n139 VSUBS 0.009274f
C231 B.n140 VSUBS 0.009274f
C232 B.n141 VSUBS 0.009274f
C233 B.n142 VSUBS 0.009274f
C234 B.n143 VSUBS 0.009274f
C235 B.n144 VSUBS 0.009274f
C236 B.n145 VSUBS 0.009274f
C237 B.n146 VSUBS 0.009274f
C238 B.n147 VSUBS 0.009274f
C239 B.n148 VSUBS 0.00641f
C240 B.n149 VSUBS 0.021487f
C241 B.n150 VSUBS 0.007501f
C242 B.n151 VSUBS 0.009274f
C243 B.n152 VSUBS 0.009274f
C244 B.n153 VSUBS 0.009274f
C245 B.n154 VSUBS 0.009274f
C246 B.n155 VSUBS 0.009274f
C247 B.n156 VSUBS 0.009274f
C248 B.n157 VSUBS 0.009274f
C249 B.n158 VSUBS 0.009274f
C250 B.n159 VSUBS 0.009274f
C251 B.n160 VSUBS 0.009274f
C252 B.n161 VSUBS 0.009274f
C253 B.n162 VSUBS 0.007501f
C254 B.n163 VSUBS 0.021487f
C255 B.n164 VSUBS 0.00641f
C256 B.n165 VSUBS 0.009274f
C257 B.n166 VSUBS 0.009274f
C258 B.n167 VSUBS 0.009274f
C259 B.n168 VSUBS 0.009274f
C260 B.n169 VSUBS 0.009274f
C261 B.n170 VSUBS 0.009274f
C262 B.n171 VSUBS 0.009274f
C263 B.n172 VSUBS 0.009274f
C264 B.n173 VSUBS 0.009274f
C265 B.n174 VSUBS 0.009274f
C266 B.n175 VSUBS 0.009274f
C267 B.n176 VSUBS 0.009274f
C268 B.n177 VSUBS 0.009274f
C269 B.n178 VSUBS 0.009274f
C270 B.n179 VSUBS 0.021663f
C271 B.n180 VSUBS 0.020511f
C272 B.n181 VSUBS 0.021494f
C273 B.n182 VSUBS 0.009274f
C274 B.n183 VSUBS 0.009274f
C275 B.n184 VSUBS 0.009274f
C276 B.n185 VSUBS 0.009274f
C277 B.n186 VSUBS 0.009274f
C278 B.n187 VSUBS 0.009274f
C279 B.n188 VSUBS 0.009274f
C280 B.n189 VSUBS 0.009274f
C281 B.n190 VSUBS 0.009274f
C282 B.n191 VSUBS 0.009274f
C283 B.n192 VSUBS 0.009274f
C284 B.n193 VSUBS 0.009274f
C285 B.n194 VSUBS 0.009274f
C286 B.n195 VSUBS 0.009274f
C287 B.n196 VSUBS 0.009274f
C288 B.n197 VSUBS 0.009274f
C289 B.n198 VSUBS 0.009274f
C290 B.n199 VSUBS 0.009274f
C291 B.n200 VSUBS 0.009274f
C292 B.n201 VSUBS 0.009274f
C293 B.n202 VSUBS 0.009274f
C294 B.n203 VSUBS 0.009274f
C295 B.n204 VSUBS 0.009274f
C296 B.n205 VSUBS 0.009274f
C297 B.n206 VSUBS 0.009274f
C298 B.n207 VSUBS 0.009274f
C299 B.n208 VSUBS 0.009274f
C300 B.n209 VSUBS 0.009274f
C301 B.n210 VSUBS 0.009274f
C302 B.n211 VSUBS 0.009274f
C303 B.n212 VSUBS 0.009274f
C304 B.n213 VSUBS 0.009274f
C305 B.n214 VSUBS 0.009274f
C306 B.n215 VSUBS 0.009274f
C307 B.n216 VSUBS 0.009274f
C308 B.n217 VSUBS 0.009274f
C309 B.n218 VSUBS 0.009274f
C310 B.n219 VSUBS 0.009274f
C311 B.n220 VSUBS 0.009274f
C312 B.n221 VSUBS 0.009274f
C313 B.n222 VSUBS 0.009274f
C314 B.n223 VSUBS 0.009274f
C315 B.n224 VSUBS 0.009274f
C316 B.n225 VSUBS 0.009274f
C317 B.n226 VSUBS 0.009274f
C318 B.n227 VSUBS 0.009274f
C319 B.n228 VSUBS 0.009274f
C320 B.n229 VSUBS 0.009274f
C321 B.n230 VSUBS 0.009274f
C322 B.n231 VSUBS 0.009274f
C323 B.n232 VSUBS 0.009274f
C324 B.n233 VSUBS 0.009274f
C325 B.n234 VSUBS 0.009274f
C326 B.n235 VSUBS 0.009274f
C327 B.n236 VSUBS 0.009274f
C328 B.n237 VSUBS 0.009274f
C329 B.n238 VSUBS 0.009274f
C330 B.n239 VSUBS 0.009274f
C331 B.n240 VSUBS 0.009274f
C332 B.n241 VSUBS 0.009274f
C333 B.n242 VSUBS 0.009274f
C334 B.n243 VSUBS 0.009274f
C335 B.n244 VSUBS 0.009274f
C336 B.n245 VSUBS 0.009274f
C337 B.n246 VSUBS 0.009274f
C338 B.n247 VSUBS 0.009274f
C339 B.n248 VSUBS 0.009274f
C340 B.n249 VSUBS 0.009274f
C341 B.n250 VSUBS 0.009274f
C342 B.n251 VSUBS 0.009274f
C343 B.n252 VSUBS 0.009274f
C344 B.n253 VSUBS 0.009274f
C345 B.n254 VSUBS 0.009274f
C346 B.n255 VSUBS 0.009274f
C347 B.n256 VSUBS 0.009274f
C348 B.n257 VSUBS 0.009274f
C349 B.n258 VSUBS 0.009274f
C350 B.n259 VSUBS 0.009274f
C351 B.n260 VSUBS 0.020342f
C352 B.n261 VSUBS 0.020342f
C353 B.n262 VSUBS 0.021663f
C354 B.n263 VSUBS 0.009274f
C355 B.n264 VSUBS 0.009274f
C356 B.n265 VSUBS 0.009274f
C357 B.n266 VSUBS 0.009274f
C358 B.n267 VSUBS 0.009274f
C359 B.n268 VSUBS 0.009274f
C360 B.n269 VSUBS 0.009274f
C361 B.n270 VSUBS 0.009274f
C362 B.n271 VSUBS 0.009274f
C363 B.n272 VSUBS 0.009274f
C364 B.n273 VSUBS 0.009274f
C365 B.n274 VSUBS 0.009274f
C366 B.n275 VSUBS 0.009274f
C367 B.n276 VSUBS 0.009274f
C368 B.n277 VSUBS 0.00641f
C369 B.n278 VSUBS 0.021487f
C370 B.n279 VSUBS 0.007501f
C371 B.n280 VSUBS 0.009274f
C372 B.n281 VSUBS 0.009274f
C373 B.n282 VSUBS 0.009274f
C374 B.n283 VSUBS 0.009274f
C375 B.n284 VSUBS 0.009274f
C376 B.n285 VSUBS 0.009274f
C377 B.n286 VSUBS 0.009274f
C378 B.n287 VSUBS 0.009274f
C379 B.n288 VSUBS 0.009274f
C380 B.n289 VSUBS 0.009274f
C381 B.n290 VSUBS 0.009274f
C382 B.n291 VSUBS 0.007501f
C383 B.n292 VSUBS 0.009274f
C384 B.n293 VSUBS 0.009274f
C385 B.n294 VSUBS 0.009274f
C386 B.n295 VSUBS 0.009274f
C387 B.n296 VSUBS 0.009274f
C388 B.n297 VSUBS 0.009274f
C389 B.n298 VSUBS 0.009274f
C390 B.n299 VSUBS 0.009274f
C391 B.n300 VSUBS 0.009274f
C392 B.n301 VSUBS 0.009274f
C393 B.n302 VSUBS 0.009274f
C394 B.n303 VSUBS 0.009274f
C395 B.n304 VSUBS 0.009274f
C396 B.n305 VSUBS 0.009274f
C397 B.n306 VSUBS 0.009274f
C398 B.n307 VSUBS 0.009274f
C399 B.n308 VSUBS 0.021663f
C400 B.n309 VSUBS 0.020342f
C401 B.n310 VSUBS 0.020342f
C402 B.n311 VSUBS 0.009274f
C403 B.n312 VSUBS 0.009274f
C404 B.n313 VSUBS 0.009274f
C405 B.n314 VSUBS 0.009274f
C406 B.n315 VSUBS 0.009274f
C407 B.n316 VSUBS 0.009274f
C408 B.n317 VSUBS 0.009274f
C409 B.n318 VSUBS 0.009274f
C410 B.n319 VSUBS 0.009274f
C411 B.n320 VSUBS 0.009274f
C412 B.n321 VSUBS 0.009274f
C413 B.n322 VSUBS 0.009274f
C414 B.n323 VSUBS 0.009274f
C415 B.n324 VSUBS 0.009274f
C416 B.n325 VSUBS 0.009274f
C417 B.n326 VSUBS 0.009274f
C418 B.n327 VSUBS 0.009274f
C419 B.n328 VSUBS 0.009274f
C420 B.n329 VSUBS 0.009274f
C421 B.n330 VSUBS 0.009274f
C422 B.n331 VSUBS 0.009274f
C423 B.n332 VSUBS 0.009274f
C424 B.n333 VSUBS 0.009274f
C425 B.n334 VSUBS 0.009274f
C426 B.n335 VSUBS 0.009274f
C427 B.n336 VSUBS 0.009274f
C428 B.n337 VSUBS 0.009274f
C429 B.n338 VSUBS 0.009274f
C430 B.n339 VSUBS 0.009274f
C431 B.n340 VSUBS 0.009274f
C432 B.n341 VSUBS 0.009274f
C433 B.n342 VSUBS 0.009274f
C434 B.n343 VSUBS 0.009274f
C435 B.n344 VSUBS 0.009274f
C436 B.n345 VSUBS 0.009274f
C437 B.n346 VSUBS 0.009274f
C438 B.n347 VSUBS 0.012102f
C439 B.n348 VSUBS 0.012892f
C440 B.n349 VSUBS 0.025636f
C441 VTAIL.t10 VSUBS 0.022905f
C442 VTAIL.t14 VSUBS 0.022905f
C443 VTAIL.n0 VSUBS 0.074554f
C444 VTAIL.n1 VSUBS 0.240238f
C445 VTAIL.t9 VSUBS 0.127017f
C446 VTAIL.n2 VSUBS 0.276756f
C447 VTAIL.t5 VSUBS 0.127017f
C448 VTAIL.n3 VSUBS 0.276756f
C449 VTAIL.t7 VSUBS 0.022905f
C450 VTAIL.t6 VSUBS 0.022905f
C451 VTAIL.n4 VSUBS 0.074554f
C452 VTAIL.n5 VSUBS 0.305898f
C453 VTAIL.t4 VSUBS 0.127017f
C454 VTAIL.n6 VSUBS 0.667949f
C455 VTAIL.t15 VSUBS 0.127017f
C456 VTAIL.n7 VSUBS 0.667949f
C457 VTAIL.t8 VSUBS 0.022905f
C458 VTAIL.t11 VSUBS 0.022905f
C459 VTAIL.n8 VSUBS 0.074554f
C460 VTAIL.n9 VSUBS 0.305898f
C461 VTAIL.t13 VSUBS 0.127017f
C462 VTAIL.n10 VSUBS 0.276756f
C463 VTAIL.t1 VSUBS 0.127017f
C464 VTAIL.n11 VSUBS 0.276756f
C465 VTAIL.t3 VSUBS 0.022905f
C466 VTAIL.t2 VSUBS 0.022905f
C467 VTAIL.n12 VSUBS 0.074554f
C468 VTAIL.n13 VSUBS 0.305898f
C469 VTAIL.t0 VSUBS 0.127017f
C470 VTAIL.n14 VSUBS 0.667949f
C471 VTAIL.t12 VSUBS 0.127017f
C472 VTAIL.n15 VSUBS 0.664201f
C473 VDD2.t0 VSUBS 0.021552f
C474 VDD2.t2 VSUBS 0.021552f
C475 VDD2.n0 VSUBS 0.082636f
C476 VDD2.t7 VSUBS 0.021552f
C477 VDD2.t4 VSUBS 0.021552f
C478 VDD2.n1 VSUBS 0.082636f
C479 VDD2.n2 VSUBS 1.29831f
C480 VDD2.t1 VSUBS 0.021552f
C481 VDD2.t6 VSUBS 0.021552f
C482 VDD2.n3 VSUBS 0.082108f
C483 VDD2.n4 VSUBS 1.16164f
C484 VDD2.t3 VSUBS 0.021552f
C485 VDD2.t5 VSUBS 0.021552f
C486 VDD2.n5 VSUBS 0.082631f
C487 VN.n0 VSUBS 0.070955f
C488 VN.t1 VSUBS 0.153094f
C489 VN.n1 VSUBS 0.042987f
C490 VN.t6 VSUBS 0.25618f
C491 VN.n2 VSUBS 0.184026f
C492 VN.t5 VSUBS 0.153094f
C493 VN.n3 VSUBS 0.154134f
C494 VN.n4 VSUBS 0.068985f
C495 VN.n5 VSUBS 0.21724f
C496 VN.n6 VSUBS 0.053175f
C497 VN.n7 VSUBS 0.053175f
C498 VN.n8 VSUBS 0.068985f
C499 VN.n9 VSUBS 0.115188f
C500 VN.n10 VSUBS 0.063871f
C501 VN.t3 VSUBS 0.228041f
C502 VN.n11 VSUBS 0.186208f
C503 VN.n12 VSUBS 0.0498f
C504 VN.n13 VSUBS 0.070955f
C505 VN.t7 VSUBS 0.153094f
C506 VN.n14 VSUBS 0.042987f
C507 VN.t2 VSUBS 0.25618f
C508 VN.n15 VSUBS 0.184026f
C509 VN.t4 VSUBS 0.153094f
C510 VN.n16 VSUBS 0.154134f
C511 VN.n17 VSUBS 0.068985f
C512 VN.n18 VSUBS 0.21724f
C513 VN.n19 VSUBS 0.053175f
C514 VN.n20 VSUBS 0.053175f
C515 VN.n21 VSUBS 0.068985f
C516 VN.n22 VSUBS 0.115188f
C517 VN.n23 VSUBS 0.063871f
C518 VN.t0 VSUBS 0.228041f
C519 VN.n24 VSUBS 0.186208f
C520 VN.n25 VSUBS 1.64696f
.ends

