* NGSPICE file created from diff_pair_sample_1616.ext - technology: sky130A

.subckt diff_pair_sample_1616 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=6.9732 pd=36.54 as=0 ps=0 w=17.88 l=1.42
X1 VTAIL.t15 VN.t0 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=2.9502 pd=18.21 as=2.9502 ps=18.21 w=17.88 l=1.42
X2 VTAIL.t2 VP.t0 VDD1.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=6.9732 pd=36.54 as=2.9502 ps=18.21 w=17.88 l=1.42
X3 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=6.9732 pd=36.54 as=0 ps=0 w=17.88 l=1.42
X4 VDD2.t1 VN.t1 VTAIL.t14 B.t2 sky130_fd_pr__nfet_01v8 ad=2.9502 pd=18.21 as=2.9502 ps=18.21 w=17.88 l=1.42
X5 VTAIL.t13 VN.t2 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9502 pd=18.21 as=2.9502 ps=18.21 w=17.88 l=1.42
X6 VTAIL.t12 VN.t3 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=6.9732 pd=36.54 as=2.9502 ps=18.21 w=17.88 l=1.42
X7 VDD1.t6 VP.t1 VTAIL.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=2.9502 pd=18.21 as=6.9732 ps=36.54 w=17.88 l=1.42
X8 VDD1.t5 VP.t2 VTAIL.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=2.9502 pd=18.21 as=6.9732 ps=36.54 w=17.88 l=1.42
X9 VDD2.t3 VN.t4 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=2.9502 pd=18.21 as=2.9502 ps=18.21 w=17.88 l=1.42
X10 VDD2.t7 VN.t5 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=2.9502 pd=18.21 as=6.9732 ps=36.54 w=17.88 l=1.42
X11 VDD2.t6 VN.t6 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=2.9502 pd=18.21 as=6.9732 ps=36.54 w=17.88 l=1.42
X12 VTAIL.t7 VP.t3 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=2.9502 pd=18.21 as=2.9502 ps=18.21 w=17.88 l=1.42
X13 VDD1.t3 VP.t4 VTAIL.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.9502 pd=18.21 as=2.9502 ps=18.21 w=17.88 l=1.42
X14 VTAIL.t8 VN.t7 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=6.9732 pd=36.54 as=2.9502 ps=18.21 w=17.88 l=1.42
X15 VDD1.t2 VP.t5 VTAIL.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=2.9502 pd=18.21 as=2.9502 ps=18.21 w=17.88 l=1.42
X16 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=6.9732 pd=36.54 as=0 ps=0 w=17.88 l=1.42
X17 VTAIL.t4 VP.t6 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=6.9732 pd=36.54 as=2.9502 ps=18.21 w=17.88 l=1.42
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.9732 pd=36.54 as=0 ps=0 w=17.88 l=1.42
X19 VTAIL.t3 VP.t7 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9502 pd=18.21 as=2.9502 ps=18.21 w=17.88 l=1.42
R0 B.n668 B.n667 585
R1 B.n668 B.n64 585
R2 B.n671 B.n670 585
R3 B.n672 B.n132 585
R4 B.n674 B.n673 585
R5 B.n676 B.n131 585
R6 B.n679 B.n678 585
R7 B.n680 B.n130 585
R8 B.n682 B.n681 585
R9 B.n684 B.n129 585
R10 B.n687 B.n686 585
R11 B.n688 B.n128 585
R12 B.n690 B.n689 585
R13 B.n692 B.n127 585
R14 B.n695 B.n694 585
R15 B.n696 B.n126 585
R16 B.n698 B.n697 585
R17 B.n700 B.n125 585
R18 B.n703 B.n702 585
R19 B.n704 B.n124 585
R20 B.n706 B.n705 585
R21 B.n708 B.n123 585
R22 B.n711 B.n710 585
R23 B.n712 B.n122 585
R24 B.n714 B.n713 585
R25 B.n716 B.n121 585
R26 B.n719 B.n718 585
R27 B.n720 B.n120 585
R28 B.n722 B.n721 585
R29 B.n724 B.n119 585
R30 B.n727 B.n726 585
R31 B.n728 B.n118 585
R32 B.n730 B.n729 585
R33 B.n732 B.n117 585
R34 B.n735 B.n734 585
R35 B.n736 B.n116 585
R36 B.n738 B.n737 585
R37 B.n740 B.n115 585
R38 B.n743 B.n742 585
R39 B.n744 B.n114 585
R40 B.n746 B.n745 585
R41 B.n748 B.n113 585
R42 B.n751 B.n750 585
R43 B.n752 B.n112 585
R44 B.n754 B.n753 585
R45 B.n756 B.n111 585
R46 B.n759 B.n758 585
R47 B.n760 B.n110 585
R48 B.n762 B.n761 585
R49 B.n764 B.n109 585
R50 B.n767 B.n766 585
R51 B.n768 B.n108 585
R52 B.n770 B.n769 585
R53 B.n772 B.n107 585
R54 B.n775 B.n774 585
R55 B.n776 B.n106 585
R56 B.n778 B.n777 585
R57 B.n780 B.n105 585
R58 B.n783 B.n782 585
R59 B.n784 B.n102 585
R60 B.n787 B.n786 585
R61 B.n789 B.n101 585
R62 B.n792 B.n791 585
R63 B.n793 B.n100 585
R64 B.n795 B.n794 585
R65 B.n797 B.n99 585
R66 B.n800 B.n799 585
R67 B.n801 B.n95 585
R68 B.n803 B.n802 585
R69 B.n805 B.n94 585
R70 B.n808 B.n807 585
R71 B.n809 B.n93 585
R72 B.n811 B.n810 585
R73 B.n813 B.n92 585
R74 B.n816 B.n815 585
R75 B.n817 B.n91 585
R76 B.n819 B.n818 585
R77 B.n821 B.n90 585
R78 B.n824 B.n823 585
R79 B.n825 B.n89 585
R80 B.n827 B.n826 585
R81 B.n829 B.n88 585
R82 B.n832 B.n831 585
R83 B.n833 B.n87 585
R84 B.n835 B.n834 585
R85 B.n837 B.n86 585
R86 B.n840 B.n839 585
R87 B.n841 B.n85 585
R88 B.n843 B.n842 585
R89 B.n845 B.n84 585
R90 B.n848 B.n847 585
R91 B.n849 B.n83 585
R92 B.n851 B.n850 585
R93 B.n853 B.n82 585
R94 B.n856 B.n855 585
R95 B.n857 B.n81 585
R96 B.n859 B.n858 585
R97 B.n861 B.n80 585
R98 B.n864 B.n863 585
R99 B.n865 B.n79 585
R100 B.n867 B.n866 585
R101 B.n869 B.n78 585
R102 B.n872 B.n871 585
R103 B.n873 B.n77 585
R104 B.n875 B.n874 585
R105 B.n877 B.n76 585
R106 B.n880 B.n879 585
R107 B.n881 B.n75 585
R108 B.n883 B.n882 585
R109 B.n885 B.n74 585
R110 B.n888 B.n887 585
R111 B.n889 B.n73 585
R112 B.n891 B.n890 585
R113 B.n893 B.n72 585
R114 B.n896 B.n895 585
R115 B.n897 B.n71 585
R116 B.n899 B.n898 585
R117 B.n901 B.n70 585
R118 B.n904 B.n903 585
R119 B.n905 B.n69 585
R120 B.n907 B.n906 585
R121 B.n909 B.n68 585
R122 B.n912 B.n911 585
R123 B.n913 B.n67 585
R124 B.n915 B.n914 585
R125 B.n917 B.n66 585
R126 B.n920 B.n919 585
R127 B.n921 B.n65 585
R128 B.n666 B.n63 585
R129 B.n924 B.n63 585
R130 B.n665 B.n62 585
R131 B.n925 B.n62 585
R132 B.n664 B.n61 585
R133 B.n926 B.n61 585
R134 B.n663 B.n662 585
R135 B.n662 B.n57 585
R136 B.n661 B.n56 585
R137 B.n932 B.n56 585
R138 B.n660 B.n55 585
R139 B.n933 B.n55 585
R140 B.n659 B.n54 585
R141 B.n934 B.n54 585
R142 B.n658 B.n657 585
R143 B.n657 B.n50 585
R144 B.n656 B.n49 585
R145 B.n940 B.n49 585
R146 B.n655 B.n48 585
R147 B.n941 B.n48 585
R148 B.n654 B.n47 585
R149 B.n942 B.n47 585
R150 B.n653 B.n652 585
R151 B.n652 B.n43 585
R152 B.n651 B.n42 585
R153 B.n948 B.n42 585
R154 B.n650 B.n41 585
R155 B.n949 B.n41 585
R156 B.n649 B.n40 585
R157 B.n950 B.n40 585
R158 B.n648 B.n647 585
R159 B.n647 B.n36 585
R160 B.n646 B.n35 585
R161 B.n956 B.n35 585
R162 B.n645 B.n34 585
R163 B.n957 B.n34 585
R164 B.n644 B.n33 585
R165 B.n958 B.n33 585
R166 B.n643 B.n642 585
R167 B.n642 B.n32 585
R168 B.n641 B.n28 585
R169 B.n964 B.n28 585
R170 B.n640 B.n27 585
R171 B.n965 B.n27 585
R172 B.n639 B.n26 585
R173 B.n966 B.n26 585
R174 B.n638 B.n637 585
R175 B.n637 B.n22 585
R176 B.n636 B.n21 585
R177 B.n972 B.n21 585
R178 B.n635 B.n20 585
R179 B.n973 B.n20 585
R180 B.n634 B.n19 585
R181 B.n974 B.n19 585
R182 B.n633 B.n632 585
R183 B.n632 B.n15 585
R184 B.n631 B.n14 585
R185 B.n980 B.n14 585
R186 B.n630 B.n13 585
R187 B.n981 B.n13 585
R188 B.n629 B.n12 585
R189 B.n982 B.n12 585
R190 B.n628 B.n627 585
R191 B.n627 B.n8 585
R192 B.n626 B.n7 585
R193 B.n988 B.n7 585
R194 B.n625 B.n6 585
R195 B.n989 B.n6 585
R196 B.n624 B.n5 585
R197 B.n990 B.n5 585
R198 B.n623 B.n622 585
R199 B.n622 B.n4 585
R200 B.n621 B.n133 585
R201 B.n621 B.n620 585
R202 B.n611 B.n134 585
R203 B.n135 B.n134 585
R204 B.n613 B.n612 585
R205 B.n614 B.n613 585
R206 B.n610 B.n139 585
R207 B.n143 B.n139 585
R208 B.n609 B.n608 585
R209 B.n608 B.n607 585
R210 B.n141 B.n140 585
R211 B.n142 B.n141 585
R212 B.n600 B.n599 585
R213 B.n601 B.n600 585
R214 B.n598 B.n148 585
R215 B.n148 B.n147 585
R216 B.n597 B.n596 585
R217 B.n596 B.n595 585
R218 B.n150 B.n149 585
R219 B.n151 B.n150 585
R220 B.n588 B.n587 585
R221 B.n589 B.n588 585
R222 B.n586 B.n156 585
R223 B.n156 B.n155 585
R224 B.n585 B.n584 585
R225 B.n584 B.n583 585
R226 B.n158 B.n157 585
R227 B.n576 B.n158 585
R228 B.n575 B.n574 585
R229 B.n577 B.n575 585
R230 B.n573 B.n163 585
R231 B.n163 B.n162 585
R232 B.n572 B.n571 585
R233 B.n571 B.n570 585
R234 B.n165 B.n164 585
R235 B.n166 B.n165 585
R236 B.n563 B.n562 585
R237 B.n564 B.n563 585
R238 B.n561 B.n171 585
R239 B.n171 B.n170 585
R240 B.n560 B.n559 585
R241 B.n559 B.n558 585
R242 B.n173 B.n172 585
R243 B.n174 B.n173 585
R244 B.n551 B.n550 585
R245 B.n552 B.n551 585
R246 B.n549 B.n179 585
R247 B.n179 B.n178 585
R248 B.n548 B.n547 585
R249 B.n547 B.n546 585
R250 B.n181 B.n180 585
R251 B.n182 B.n181 585
R252 B.n539 B.n538 585
R253 B.n540 B.n539 585
R254 B.n537 B.n187 585
R255 B.n187 B.n186 585
R256 B.n536 B.n535 585
R257 B.n535 B.n534 585
R258 B.n189 B.n188 585
R259 B.n190 B.n189 585
R260 B.n527 B.n526 585
R261 B.n528 B.n527 585
R262 B.n525 B.n195 585
R263 B.n195 B.n194 585
R264 B.n524 B.n523 585
R265 B.n523 B.n522 585
R266 B.n519 B.n199 585
R267 B.n518 B.n517 585
R268 B.n515 B.n200 585
R269 B.n515 B.n198 585
R270 B.n514 B.n513 585
R271 B.n512 B.n511 585
R272 B.n510 B.n202 585
R273 B.n508 B.n507 585
R274 B.n506 B.n203 585
R275 B.n505 B.n504 585
R276 B.n502 B.n204 585
R277 B.n500 B.n499 585
R278 B.n498 B.n205 585
R279 B.n497 B.n496 585
R280 B.n494 B.n206 585
R281 B.n492 B.n491 585
R282 B.n490 B.n207 585
R283 B.n489 B.n488 585
R284 B.n486 B.n208 585
R285 B.n484 B.n483 585
R286 B.n482 B.n209 585
R287 B.n481 B.n480 585
R288 B.n478 B.n210 585
R289 B.n476 B.n475 585
R290 B.n474 B.n211 585
R291 B.n473 B.n472 585
R292 B.n470 B.n212 585
R293 B.n468 B.n467 585
R294 B.n466 B.n213 585
R295 B.n465 B.n464 585
R296 B.n462 B.n214 585
R297 B.n460 B.n459 585
R298 B.n458 B.n215 585
R299 B.n457 B.n456 585
R300 B.n454 B.n216 585
R301 B.n452 B.n451 585
R302 B.n450 B.n217 585
R303 B.n449 B.n448 585
R304 B.n446 B.n218 585
R305 B.n444 B.n443 585
R306 B.n442 B.n219 585
R307 B.n441 B.n440 585
R308 B.n438 B.n220 585
R309 B.n436 B.n435 585
R310 B.n434 B.n221 585
R311 B.n433 B.n432 585
R312 B.n430 B.n222 585
R313 B.n428 B.n427 585
R314 B.n426 B.n223 585
R315 B.n425 B.n424 585
R316 B.n422 B.n224 585
R317 B.n420 B.n419 585
R318 B.n418 B.n225 585
R319 B.n417 B.n416 585
R320 B.n414 B.n226 585
R321 B.n412 B.n411 585
R322 B.n410 B.n227 585
R323 B.n409 B.n408 585
R324 B.n406 B.n228 585
R325 B.n404 B.n403 585
R326 B.n401 B.n229 585
R327 B.n400 B.n399 585
R328 B.n397 B.n232 585
R329 B.n395 B.n394 585
R330 B.n393 B.n233 585
R331 B.n392 B.n391 585
R332 B.n389 B.n234 585
R333 B.n387 B.n386 585
R334 B.n385 B.n235 585
R335 B.n383 B.n382 585
R336 B.n380 B.n238 585
R337 B.n378 B.n377 585
R338 B.n376 B.n239 585
R339 B.n375 B.n374 585
R340 B.n372 B.n240 585
R341 B.n370 B.n369 585
R342 B.n368 B.n241 585
R343 B.n367 B.n366 585
R344 B.n364 B.n242 585
R345 B.n362 B.n361 585
R346 B.n360 B.n243 585
R347 B.n359 B.n358 585
R348 B.n356 B.n244 585
R349 B.n354 B.n353 585
R350 B.n352 B.n245 585
R351 B.n351 B.n350 585
R352 B.n348 B.n246 585
R353 B.n346 B.n345 585
R354 B.n344 B.n247 585
R355 B.n343 B.n342 585
R356 B.n340 B.n248 585
R357 B.n338 B.n337 585
R358 B.n336 B.n249 585
R359 B.n335 B.n334 585
R360 B.n332 B.n250 585
R361 B.n330 B.n329 585
R362 B.n328 B.n251 585
R363 B.n327 B.n326 585
R364 B.n324 B.n252 585
R365 B.n322 B.n321 585
R366 B.n320 B.n253 585
R367 B.n319 B.n318 585
R368 B.n316 B.n254 585
R369 B.n314 B.n313 585
R370 B.n312 B.n255 585
R371 B.n311 B.n310 585
R372 B.n308 B.n256 585
R373 B.n306 B.n305 585
R374 B.n304 B.n257 585
R375 B.n303 B.n302 585
R376 B.n300 B.n258 585
R377 B.n298 B.n297 585
R378 B.n296 B.n259 585
R379 B.n295 B.n294 585
R380 B.n292 B.n260 585
R381 B.n290 B.n289 585
R382 B.n288 B.n261 585
R383 B.n287 B.n286 585
R384 B.n284 B.n262 585
R385 B.n282 B.n281 585
R386 B.n280 B.n263 585
R387 B.n279 B.n278 585
R388 B.n276 B.n264 585
R389 B.n274 B.n273 585
R390 B.n272 B.n265 585
R391 B.n271 B.n270 585
R392 B.n268 B.n266 585
R393 B.n197 B.n196 585
R394 B.n521 B.n520 585
R395 B.n522 B.n521 585
R396 B.n193 B.n192 585
R397 B.n194 B.n193 585
R398 B.n530 B.n529 585
R399 B.n529 B.n528 585
R400 B.n531 B.n191 585
R401 B.n191 B.n190 585
R402 B.n533 B.n532 585
R403 B.n534 B.n533 585
R404 B.n185 B.n184 585
R405 B.n186 B.n185 585
R406 B.n542 B.n541 585
R407 B.n541 B.n540 585
R408 B.n543 B.n183 585
R409 B.n183 B.n182 585
R410 B.n545 B.n544 585
R411 B.n546 B.n545 585
R412 B.n177 B.n176 585
R413 B.n178 B.n177 585
R414 B.n554 B.n553 585
R415 B.n553 B.n552 585
R416 B.n555 B.n175 585
R417 B.n175 B.n174 585
R418 B.n557 B.n556 585
R419 B.n558 B.n557 585
R420 B.n169 B.n168 585
R421 B.n170 B.n169 585
R422 B.n566 B.n565 585
R423 B.n565 B.n564 585
R424 B.n567 B.n167 585
R425 B.n167 B.n166 585
R426 B.n569 B.n568 585
R427 B.n570 B.n569 585
R428 B.n161 B.n160 585
R429 B.n162 B.n161 585
R430 B.n579 B.n578 585
R431 B.n578 B.n577 585
R432 B.n580 B.n159 585
R433 B.n576 B.n159 585
R434 B.n582 B.n581 585
R435 B.n583 B.n582 585
R436 B.n154 B.n153 585
R437 B.n155 B.n154 585
R438 B.n591 B.n590 585
R439 B.n590 B.n589 585
R440 B.n592 B.n152 585
R441 B.n152 B.n151 585
R442 B.n594 B.n593 585
R443 B.n595 B.n594 585
R444 B.n146 B.n145 585
R445 B.n147 B.n146 585
R446 B.n603 B.n602 585
R447 B.n602 B.n601 585
R448 B.n604 B.n144 585
R449 B.n144 B.n142 585
R450 B.n606 B.n605 585
R451 B.n607 B.n606 585
R452 B.n138 B.n137 585
R453 B.n143 B.n138 585
R454 B.n616 B.n615 585
R455 B.n615 B.n614 585
R456 B.n617 B.n136 585
R457 B.n136 B.n135 585
R458 B.n619 B.n618 585
R459 B.n620 B.n619 585
R460 B.n2 B.n0 585
R461 B.n4 B.n2 585
R462 B.n3 B.n1 585
R463 B.n989 B.n3 585
R464 B.n987 B.n986 585
R465 B.n988 B.n987 585
R466 B.n985 B.n9 585
R467 B.n9 B.n8 585
R468 B.n984 B.n983 585
R469 B.n983 B.n982 585
R470 B.n11 B.n10 585
R471 B.n981 B.n11 585
R472 B.n979 B.n978 585
R473 B.n980 B.n979 585
R474 B.n977 B.n16 585
R475 B.n16 B.n15 585
R476 B.n976 B.n975 585
R477 B.n975 B.n974 585
R478 B.n18 B.n17 585
R479 B.n973 B.n18 585
R480 B.n971 B.n970 585
R481 B.n972 B.n971 585
R482 B.n969 B.n23 585
R483 B.n23 B.n22 585
R484 B.n968 B.n967 585
R485 B.n967 B.n966 585
R486 B.n25 B.n24 585
R487 B.n965 B.n25 585
R488 B.n963 B.n962 585
R489 B.n964 B.n963 585
R490 B.n961 B.n29 585
R491 B.n32 B.n29 585
R492 B.n960 B.n959 585
R493 B.n959 B.n958 585
R494 B.n31 B.n30 585
R495 B.n957 B.n31 585
R496 B.n955 B.n954 585
R497 B.n956 B.n955 585
R498 B.n953 B.n37 585
R499 B.n37 B.n36 585
R500 B.n952 B.n951 585
R501 B.n951 B.n950 585
R502 B.n39 B.n38 585
R503 B.n949 B.n39 585
R504 B.n947 B.n946 585
R505 B.n948 B.n947 585
R506 B.n945 B.n44 585
R507 B.n44 B.n43 585
R508 B.n944 B.n943 585
R509 B.n943 B.n942 585
R510 B.n46 B.n45 585
R511 B.n941 B.n46 585
R512 B.n939 B.n938 585
R513 B.n940 B.n939 585
R514 B.n937 B.n51 585
R515 B.n51 B.n50 585
R516 B.n936 B.n935 585
R517 B.n935 B.n934 585
R518 B.n53 B.n52 585
R519 B.n933 B.n53 585
R520 B.n931 B.n930 585
R521 B.n932 B.n931 585
R522 B.n929 B.n58 585
R523 B.n58 B.n57 585
R524 B.n928 B.n927 585
R525 B.n927 B.n926 585
R526 B.n60 B.n59 585
R527 B.n925 B.n60 585
R528 B.n923 B.n922 585
R529 B.n924 B.n923 585
R530 B.n992 B.n991 585
R531 B.n991 B.n990 585
R532 B.n236 B.t8 508.586
R533 B.n230 B.t19 508.586
R534 B.n96 B.t12 508.586
R535 B.n103 B.t16 508.586
R536 B.n521 B.n199 506.916
R537 B.n923 B.n65 506.916
R538 B.n523 B.n197 506.916
R539 B.n668 B.n63 506.916
R540 B.n669 B.n64 256.663
R541 B.n675 B.n64 256.663
R542 B.n677 B.n64 256.663
R543 B.n683 B.n64 256.663
R544 B.n685 B.n64 256.663
R545 B.n691 B.n64 256.663
R546 B.n693 B.n64 256.663
R547 B.n699 B.n64 256.663
R548 B.n701 B.n64 256.663
R549 B.n707 B.n64 256.663
R550 B.n709 B.n64 256.663
R551 B.n715 B.n64 256.663
R552 B.n717 B.n64 256.663
R553 B.n723 B.n64 256.663
R554 B.n725 B.n64 256.663
R555 B.n731 B.n64 256.663
R556 B.n733 B.n64 256.663
R557 B.n739 B.n64 256.663
R558 B.n741 B.n64 256.663
R559 B.n747 B.n64 256.663
R560 B.n749 B.n64 256.663
R561 B.n755 B.n64 256.663
R562 B.n757 B.n64 256.663
R563 B.n763 B.n64 256.663
R564 B.n765 B.n64 256.663
R565 B.n771 B.n64 256.663
R566 B.n773 B.n64 256.663
R567 B.n779 B.n64 256.663
R568 B.n781 B.n64 256.663
R569 B.n788 B.n64 256.663
R570 B.n790 B.n64 256.663
R571 B.n796 B.n64 256.663
R572 B.n798 B.n64 256.663
R573 B.n804 B.n64 256.663
R574 B.n806 B.n64 256.663
R575 B.n812 B.n64 256.663
R576 B.n814 B.n64 256.663
R577 B.n820 B.n64 256.663
R578 B.n822 B.n64 256.663
R579 B.n828 B.n64 256.663
R580 B.n830 B.n64 256.663
R581 B.n836 B.n64 256.663
R582 B.n838 B.n64 256.663
R583 B.n844 B.n64 256.663
R584 B.n846 B.n64 256.663
R585 B.n852 B.n64 256.663
R586 B.n854 B.n64 256.663
R587 B.n860 B.n64 256.663
R588 B.n862 B.n64 256.663
R589 B.n868 B.n64 256.663
R590 B.n870 B.n64 256.663
R591 B.n876 B.n64 256.663
R592 B.n878 B.n64 256.663
R593 B.n884 B.n64 256.663
R594 B.n886 B.n64 256.663
R595 B.n892 B.n64 256.663
R596 B.n894 B.n64 256.663
R597 B.n900 B.n64 256.663
R598 B.n902 B.n64 256.663
R599 B.n908 B.n64 256.663
R600 B.n910 B.n64 256.663
R601 B.n916 B.n64 256.663
R602 B.n918 B.n64 256.663
R603 B.n516 B.n198 256.663
R604 B.n201 B.n198 256.663
R605 B.n509 B.n198 256.663
R606 B.n503 B.n198 256.663
R607 B.n501 B.n198 256.663
R608 B.n495 B.n198 256.663
R609 B.n493 B.n198 256.663
R610 B.n487 B.n198 256.663
R611 B.n485 B.n198 256.663
R612 B.n479 B.n198 256.663
R613 B.n477 B.n198 256.663
R614 B.n471 B.n198 256.663
R615 B.n469 B.n198 256.663
R616 B.n463 B.n198 256.663
R617 B.n461 B.n198 256.663
R618 B.n455 B.n198 256.663
R619 B.n453 B.n198 256.663
R620 B.n447 B.n198 256.663
R621 B.n445 B.n198 256.663
R622 B.n439 B.n198 256.663
R623 B.n437 B.n198 256.663
R624 B.n431 B.n198 256.663
R625 B.n429 B.n198 256.663
R626 B.n423 B.n198 256.663
R627 B.n421 B.n198 256.663
R628 B.n415 B.n198 256.663
R629 B.n413 B.n198 256.663
R630 B.n407 B.n198 256.663
R631 B.n405 B.n198 256.663
R632 B.n398 B.n198 256.663
R633 B.n396 B.n198 256.663
R634 B.n390 B.n198 256.663
R635 B.n388 B.n198 256.663
R636 B.n381 B.n198 256.663
R637 B.n379 B.n198 256.663
R638 B.n373 B.n198 256.663
R639 B.n371 B.n198 256.663
R640 B.n365 B.n198 256.663
R641 B.n363 B.n198 256.663
R642 B.n357 B.n198 256.663
R643 B.n355 B.n198 256.663
R644 B.n349 B.n198 256.663
R645 B.n347 B.n198 256.663
R646 B.n341 B.n198 256.663
R647 B.n339 B.n198 256.663
R648 B.n333 B.n198 256.663
R649 B.n331 B.n198 256.663
R650 B.n325 B.n198 256.663
R651 B.n323 B.n198 256.663
R652 B.n317 B.n198 256.663
R653 B.n315 B.n198 256.663
R654 B.n309 B.n198 256.663
R655 B.n307 B.n198 256.663
R656 B.n301 B.n198 256.663
R657 B.n299 B.n198 256.663
R658 B.n293 B.n198 256.663
R659 B.n291 B.n198 256.663
R660 B.n285 B.n198 256.663
R661 B.n283 B.n198 256.663
R662 B.n277 B.n198 256.663
R663 B.n275 B.n198 256.663
R664 B.n269 B.n198 256.663
R665 B.n267 B.n198 256.663
R666 B.n521 B.n193 163.367
R667 B.n529 B.n193 163.367
R668 B.n529 B.n191 163.367
R669 B.n533 B.n191 163.367
R670 B.n533 B.n185 163.367
R671 B.n541 B.n185 163.367
R672 B.n541 B.n183 163.367
R673 B.n545 B.n183 163.367
R674 B.n545 B.n177 163.367
R675 B.n553 B.n177 163.367
R676 B.n553 B.n175 163.367
R677 B.n557 B.n175 163.367
R678 B.n557 B.n169 163.367
R679 B.n565 B.n169 163.367
R680 B.n565 B.n167 163.367
R681 B.n569 B.n167 163.367
R682 B.n569 B.n161 163.367
R683 B.n578 B.n161 163.367
R684 B.n578 B.n159 163.367
R685 B.n582 B.n159 163.367
R686 B.n582 B.n154 163.367
R687 B.n590 B.n154 163.367
R688 B.n590 B.n152 163.367
R689 B.n594 B.n152 163.367
R690 B.n594 B.n146 163.367
R691 B.n602 B.n146 163.367
R692 B.n602 B.n144 163.367
R693 B.n606 B.n144 163.367
R694 B.n606 B.n138 163.367
R695 B.n615 B.n138 163.367
R696 B.n615 B.n136 163.367
R697 B.n619 B.n136 163.367
R698 B.n619 B.n2 163.367
R699 B.n991 B.n2 163.367
R700 B.n991 B.n3 163.367
R701 B.n987 B.n3 163.367
R702 B.n987 B.n9 163.367
R703 B.n983 B.n9 163.367
R704 B.n983 B.n11 163.367
R705 B.n979 B.n11 163.367
R706 B.n979 B.n16 163.367
R707 B.n975 B.n16 163.367
R708 B.n975 B.n18 163.367
R709 B.n971 B.n18 163.367
R710 B.n971 B.n23 163.367
R711 B.n967 B.n23 163.367
R712 B.n967 B.n25 163.367
R713 B.n963 B.n25 163.367
R714 B.n963 B.n29 163.367
R715 B.n959 B.n29 163.367
R716 B.n959 B.n31 163.367
R717 B.n955 B.n31 163.367
R718 B.n955 B.n37 163.367
R719 B.n951 B.n37 163.367
R720 B.n951 B.n39 163.367
R721 B.n947 B.n39 163.367
R722 B.n947 B.n44 163.367
R723 B.n943 B.n44 163.367
R724 B.n943 B.n46 163.367
R725 B.n939 B.n46 163.367
R726 B.n939 B.n51 163.367
R727 B.n935 B.n51 163.367
R728 B.n935 B.n53 163.367
R729 B.n931 B.n53 163.367
R730 B.n931 B.n58 163.367
R731 B.n927 B.n58 163.367
R732 B.n927 B.n60 163.367
R733 B.n923 B.n60 163.367
R734 B.n517 B.n515 163.367
R735 B.n515 B.n514 163.367
R736 B.n511 B.n510 163.367
R737 B.n508 B.n203 163.367
R738 B.n504 B.n502 163.367
R739 B.n500 B.n205 163.367
R740 B.n496 B.n494 163.367
R741 B.n492 B.n207 163.367
R742 B.n488 B.n486 163.367
R743 B.n484 B.n209 163.367
R744 B.n480 B.n478 163.367
R745 B.n476 B.n211 163.367
R746 B.n472 B.n470 163.367
R747 B.n468 B.n213 163.367
R748 B.n464 B.n462 163.367
R749 B.n460 B.n215 163.367
R750 B.n456 B.n454 163.367
R751 B.n452 B.n217 163.367
R752 B.n448 B.n446 163.367
R753 B.n444 B.n219 163.367
R754 B.n440 B.n438 163.367
R755 B.n436 B.n221 163.367
R756 B.n432 B.n430 163.367
R757 B.n428 B.n223 163.367
R758 B.n424 B.n422 163.367
R759 B.n420 B.n225 163.367
R760 B.n416 B.n414 163.367
R761 B.n412 B.n227 163.367
R762 B.n408 B.n406 163.367
R763 B.n404 B.n229 163.367
R764 B.n399 B.n397 163.367
R765 B.n395 B.n233 163.367
R766 B.n391 B.n389 163.367
R767 B.n387 B.n235 163.367
R768 B.n382 B.n380 163.367
R769 B.n378 B.n239 163.367
R770 B.n374 B.n372 163.367
R771 B.n370 B.n241 163.367
R772 B.n366 B.n364 163.367
R773 B.n362 B.n243 163.367
R774 B.n358 B.n356 163.367
R775 B.n354 B.n245 163.367
R776 B.n350 B.n348 163.367
R777 B.n346 B.n247 163.367
R778 B.n342 B.n340 163.367
R779 B.n338 B.n249 163.367
R780 B.n334 B.n332 163.367
R781 B.n330 B.n251 163.367
R782 B.n326 B.n324 163.367
R783 B.n322 B.n253 163.367
R784 B.n318 B.n316 163.367
R785 B.n314 B.n255 163.367
R786 B.n310 B.n308 163.367
R787 B.n306 B.n257 163.367
R788 B.n302 B.n300 163.367
R789 B.n298 B.n259 163.367
R790 B.n294 B.n292 163.367
R791 B.n290 B.n261 163.367
R792 B.n286 B.n284 163.367
R793 B.n282 B.n263 163.367
R794 B.n278 B.n276 163.367
R795 B.n274 B.n265 163.367
R796 B.n270 B.n268 163.367
R797 B.n523 B.n195 163.367
R798 B.n527 B.n195 163.367
R799 B.n527 B.n189 163.367
R800 B.n535 B.n189 163.367
R801 B.n535 B.n187 163.367
R802 B.n539 B.n187 163.367
R803 B.n539 B.n181 163.367
R804 B.n547 B.n181 163.367
R805 B.n547 B.n179 163.367
R806 B.n551 B.n179 163.367
R807 B.n551 B.n173 163.367
R808 B.n559 B.n173 163.367
R809 B.n559 B.n171 163.367
R810 B.n563 B.n171 163.367
R811 B.n563 B.n165 163.367
R812 B.n571 B.n165 163.367
R813 B.n571 B.n163 163.367
R814 B.n575 B.n163 163.367
R815 B.n575 B.n158 163.367
R816 B.n584 B.n158 163.367
R817 B.n584 B.n156 163.367
R818 B.n588 B.n156 163.367
R819 B.n588 B.n150 163.367
R820 B.n596 B.n150 163.367
R821 B.n596 B.n148 163.367
R822 B.n600 B.n148 163.367
R823 B.n600 B.n141 163.367
R824 B.n608 B.n141 163.367
R825 B.n608 B.n139 163.367
R826 B.n613 B.n139 163.367
R827 B.n613 B.n134 163.367
R828 B.n621 B.n134 163.367
R829 B.n622 B.n621 163.367
R830 B.n622 B.n5 163.367
R831 B.n6 B.n5 163.367
R832 B.n7 B.n6 163.367
R833 B.n627 B.n7 163.367
R834 B.n627 B.n12 163.367
R835 B.n13 B.n12 163.367
R836 B.n14 B.n13 163.367
R837 B.n632 B.n14 163.367
R838 B.n632 B.n19 163.367
R839 B.n20 B.n19 163.367
R840 B.n21 B.n20 163.367
R841 B.n637 B.n21 163.367
R842 B.n637 B.n26 163.367
R843 B.n27 B.n26 163.367
R844 B.n28 B.n27 163.367
R845 B.n642 B.n28 163.367
R846 B.n642 B.n33 163.367
R847 B.n34 B.n33 163.367
R848 B.n35 B.n34 163.367
R849 B.n647 B.n35 163.367
R850 B.n647 B.n40 163.367
R851 B.n41 B.n40 163.367
R852 B.n42 B.n41 163.367
R853 B.n652 B.n42 163.367
R854 B.n652 B.n47 163.367
R855 B.n48 B.n47 163.367
R856 B.n49 B.n48 163.367
R857 B.n657 B.n49 163.367
R858 B.n657 B.n54 163.367
R859 B.n55 B.n54 163.367
R860 B.n56 B.n55 163.367
R861 B.n662 B.n56 163.367
R862 B.n662 B.n61 163.367
R863 B.n62 B.n61 163.367
R864 B.n63 B.n62 163.367
R865 B.n919 B.n917 163.367
R866 B.n915 B.n67 163.367
R867 B.n911 B.n909 163.367
R868 B.n907 B.n69 163.367
R869 B.n903 B.n901 163.367
R870 B.n899 B.n71 163.367
R871 B.n895 B.n893 163.367
R872 B.n891 B.n73 163.367
R873 B.n887 B.n885 163.367
R874 B.n883 B.n75 163.367
R875 B.n879 B.n877 163.367
R876 B.n875 B.n77 163.367
R877 B.n871 B.n869 163.367
R878 B.n867 B.n79 163.367
R879 B.n863 B.n861 163.367
R880 B.n859 B.n81 163.367
R881 B.n855 B.n853 163.367
R882 B.n851 B.n83 163.367
R883 B.n847 B.n845 163.367
R884 B.n843 B.n85 163.367
R885 B.n839 B.n837 163.367
R886 B.n835 B.n87 163.367
R887 B.n831 B.n829 163.367
R888 B.n827 B.n89 163.367
R889 B.n823 B.n821 163.367
R890 B.n819 B.n91 163.367
R891 B.n815 B.n813 163.367
R892 B.n811 B.n93 163.367
R893 B.n807 B.n805 163.367
R894 B.n803 B.n95 163.367
R895 B.n799 B.n797 163.367
R896 B.n795 B.n100 163.367
R897 B.n791 B.n789 163.367
R898 B.n787 B.n102 163.367
R899 B.n782 B.n780 163.367
R900 B.n778 B.n106 163.367
R901 B.n774 B.n772 163.367
R902 B.n770 B.n108 163.367
R903 B.n766 B.n764 163.367
R904 B.n762 B.n110 163.367
R905 B.n758 B.n756 163.367
R906 B.n754 B.n112 163.367
R907 B.n750 B.n748 163.367
R908 B.n746 B.n114 163.367
R909 B.n742 B.n740 163.367
R910 B.n738 B.n116 163.367
R911 B.n734 B.n732 163.367
R912 B.n730 B.n118 163.367
R913 B.n726 B.n724 163.367
R914 B.n722 B.n120 163.367
R915 B.n718 B.n716 163.367
R916 B.n714 B.n122 163.367
R917 B.n710 B.n708 163.367
R918 B.n706 B.n124 163.367
R919 B.n702 B.n700 163.367
R920 B.n698 B.n126 163.367
R921 B.n694 B.n692 163.367
R922 B.n690 B.n128 163.367
R923 B.n686 B.n684 163.367
R924 B.n682 B.n130 163.367
R925 B.n678 B.n676 163.367
R926 B.n674 B.n132 163.367
R927 B.n670 B.n668 163.367
R928 B.n236 B.t11 105.073
R929 B.n103 B.t17 105.073
R930 B.n230 B.t21 105.05
R931 B.n96 B.t14 105.05
R932 B.n516 B.n199 71.676
R933 B.n514 B.n201 71.676
R934 B.n510 B.n509 71.676
R935 B.n503 B.n203 71.676
R936 B.n502 B.n501 71.676
R937 B.n495 B.n205 71.676
R938 B.n494 B.n493 71.676
R939 B.n487 B.n207 71.676
R940 B.n486 B.n485 71.676
R941 B.n479 B.n209 71.676
R942 B.n478 B.n477 71.676
R943 B.n471 B.n211 71.676
R944 B.n470 B.n469 71.676
R945 B.n463 B.n213 71.676
R946 B.n462 B.n461 71.676
R947 B.n455 B.n215 71.676
R948 B.n454 B.n453 71.676
R949 B.n447 B.n217 71.676
R950 B.n446 B.n445 71.676
R951 B.n439 B.n219 71.676
R952 B.n438 B.n437 71.676
R953 B.n431 B.n221 71.676
R954 B.n430 B.n429 71.676
R955 B.n423 B.n223 71.676
R956 B.n422 B.n421 71.676
R957 B.n415 B.n225 71.676
R958 B.n414 B.n413 71.676
R959 B.n407 B.n227 71.676
R960 B.n406 B.n405 71.676
R961 B.n398 B.n229 71.676
R962 B.n397 B.n396 71.676
R963 B.n390 B.n233 71.676
R964 B.n389 B.n388 71.676
R965 B.n381 B.n235 71.676
R966 B.n380 B.n379 71.676
R967 B.n373 B.n239 71.676
R968 B.n372 B.n371 71.676
R969 B.n365 B.n241 71.676
R970 B.n364 B.n363 71.676
R971 B.n357 B.n243 71.676
R972 B.n356 B.n355 71.676
R973 B.n349 B.n245 71.676
R974 B.n348 B.n347 71.676
R975 B.n341 B.n247 71.676
R976 B.n340 B.n339 71.676
R977 B.n333 B.n249 71.676
R978 B.n332 B.n331 71.676
R979 B.n325 B.n251 71.676
R980 B.n324 B.n323 71.676
R981 B.n317 B.n253 71.676
R982 B.n316 B.n315 71.676
R983 B.n309 B.n255 71.676
R984 B.n308 B.n307 71.676
R985 B.n301 B.n257 71.676
R986 B.n300 B.n299 71.676
R987 B.n293 B.n259 71.676
R988 B.n292 B.n291 71.676
R989 B.n285 B.n261 71.676
R990 B.n284 B.n283 71.676
R991 B.n277 B.n263 71.676
R992 B.n276 B.n275 71.676
R993 B.n269 B.n265 71.676
R994 B.n268 B.n267 71.676
R995 B.n918 B.n65 71.676
R996 B.n917 B.n916 71.676
R997 B.n910 B.n67 71.676
R998 B.n909 B.n908 71.676
R999 B.n902 B.n69 71.676
R1000 B.n901 B.n900 71.676
R1001 B.n894 B.n71 71.676
R1002 B.n893 B.n892 71.676
R1003 B.n886 B.n73 71.676
R1004 B.n885 B.n884 71.676
R1005 B.n878 B.n75 71.676
R1006 B.n877 B.n876 71.676
R1007 B.n870 B.n77 71.676
R1008 B.n869 B.n868 71.676
R1009 B.n862 B.n79 71.676
R1010 B.n861 B.n860 71.676
R1011 B.n854 B.n81 71.676
R1012 B.n853 B.n852 71.676
R1013 B.n846 B.n83 71.676
R1014 B.n845 B.n844 71.676
R1015 B.n838 B.n85 71.676
R1016 B.n837 B.n836 71.676
R1017 B.n830 B.n87 71.676
R1018 B.n829 B.n828 71.676
R1019 B.n822 B.n89 71.676
R1020 B.n821 B.n820 71.676
R1021 B.n814 B.n91 71.676
R1022 B.n813 B.n812 71.676
R1023 B.n806 B.n93 71.676
R1024 B.n805 B.n804 71.676
R1025 B.n798 B.n95 71.676
R1026 B.n797 B.n796 71.676
R1027 B.n790 B.n100 71.676
R1028 B.n789 B.n788 71.676
R1029 B.n781 B.n102 71.676
R1030 B.n780 B.n779 71.676
R1031 B.n773 B.n106 71.676
R1032 B.n772 B.n771 71.676
R1033 B.n765 B.n108 71.676
R1034 B.n764 B.n763 71.676
R1035 B.n757 B.n110 71.676
R1036 B.n756 B.n755 71.676
R1037 B.n749 B.n112 71.676
R1038 B.n748 B.n747 71.676
R1039 B.n741 B.n114 71.676
R1040 B.n740 B.n739 71.676
R1041 B.n733 B.n116 71.676
R1042 B.n732 B.n731 71.676
R1043 B.n725 B.n118 71.676
R1044 B.n724 B.n723 71.676
R1045 B.n717 B.n120 71.676
R1046 B.n716 B.n715 71.676
R1047 B.n709 B.n122 71.676
R1048 B.n708 B.n707 71.676
R1049 B.n701 B.n124 71.676
R1050 B.n700 B.n699 71.676
R1051 B.n693 B.n126 71.676
R1052 B.n692 B.n691 71.676
R1053 B.n685 B.n128 71.676
R1054 B.n684 B.n683 71.676
R1055 B.n677 B.n130 71.676
R1056 B.n676 B.n675 71.676
R1057 B.n669 B.n132 71.676
R1058 B.n670 B.n669 71.676
R1059 B.n675 B.n674 71.676
R1060 B.n678 B.n677 71.676
R1061 B.n683 B.n682 71.676
R1062 B.n686 B.n685 71.676
R1063 B.n691 B.n690 71.676
R1064 B.n694 B.n693 71.676
R1065 B.n699 B.n698 71.676
R1066 B.n702 B.n701 71.676
R1067 B.n707 B.n706 71.676
R1068 B.n710 B.n709 71.676
R1069 B.n715 B.n714 71.676
R1070 B.n718 B.n717 71.676
R1071 B.n723 B.n722 71.676
R1072 B.n726 B.n725 71.676
R1073 B.n731 B.n730 71.676
R1074 B.n734 B.n733 71.676
R1075 B.n739 B.n738 71.676
R1076 B.n742 B.n741 71.676
R1077 B.n747 B.n746 71.676
R1078 B.n750 B.n749 71.676
R1079 B.n755 B.n754 71.676
R1080 B.n758 B.n757 71.676
R1081 B.n763 B.n762 71.676
R1082 B.n766 B.n765 71.676
R1083 B.n771 B.n770 71.676
R1084 B.n774 B.n773 71.676
R1085 B.n779 B.n778 71.676
R1086 B.n782 B.n781 71.676
R1087 B.n788 B.n787 71.676
R1088 B.n791 B.n790 71.676
R1089 B.n796 B.n795 71.676
R1090 B.n799 B.n798 71.676
R1091 B.n804 B.n803 71.676
R1092 B.n807 B.n806 71.676
R1093 B.n812 B.n811 71.676
R1094 B.n815 B.n814 71.676
R1095 B.n820 B.n819 71.676
R1096 B.n823 B.n822 71.676
R1097 B.n828 B.n827 71.676
R1098 B.n831 B.n830 71.676
R1099 B.n836 B.n835 71.676
R1100 B.n839 B.n838 71.676
R1101 B.n844 B.n843 71.676
R1102 B.n847 B.n846 71.676
R1103 B.n852 B.n851 71.676
R1104 B.n855 B.n854 71.676
R1105 B.n860 B.n859 71.676
R1106 B.n863 B.n862 71.676
R1107 B.n868 B.n867 71.676
R1108 B.n871 B.n870 71.676
R1109 B.n876 B.n875 71.676
R1110 B.n879 B.n878 71.676
R1111 B.n884 B.n883 71.676
R1112 B.n887 B.n886 71.676
R1113 B.n892 B.n891 71.676
R1114 B.n895 B.n894 71.676
R1115 B.n900 B.n899 71.676
R1116 B.n903 B.n902 71.676
R1117 B.n908 B.n907 71.676
R1118 B.n911 B.n910 71.676
R1119 B.n916 B.n915 71.676
R1120 B.n919 B.n918 71.676
R1121 B.n517 B.n516 71.676
R1122 B.n511 B.n201 71.676
R1123 B.n509 B.n508 71.676
R1124 B.n504 B.n503 71.676
R1125 B.n501 B.n500 71.676
R1126 B.n496 B.n495 71.676
R1127 B.n493 B.n492 71.676
R1128 B.n488 B.n487 71.676
R1129 B.n485 B.n484 71.676
R1130 B.n480 B.n479 71.676
R1131 B.n477 B.n476 71.676
R1132 B.n472 B.n471 71.676
R1133 B.n469 B.n468 71.676
R1134 B.n464 B.n463 71.676
R1135 B.n461 B.n460 71.676
R1136 B.n456 B.n455 71.676
R1137 B.n453 B.n452 71.676
R1138 B.n448 B.n447 71.676
R1139 B.n445 B.n444 71.676
R1140 B.n440 B.n439 71.676
R1141 B.n437 B.n436 71.676
R1142 B.n432 B.n431 71.676
R1143 B.n429 B.n428 71.676
R1144 B.n424 B.n423 71.676
R1145 B.n421 B.n420 71.676
R1146 B.n416 B.n415 71.676
R1147 B.n413 B.n412 71.676
R1148 B.n408 B.n407 71.676
R1149 B.n405 B.n404 71.676
R1150 B.n399 B.n398 71.676
R1151 B.n396 B.n395 71.676
R1152 B.n391 B.n390 71.676
R1153 B.n388 B.n387 71.676
R1154 B.n382 B.n381 71.676
R1155 B.n379 B.n378 71.676
R1156 B.n374 B.n373 71.676
R1157 B.n371 B.n370 71.676
R1158 B.n366 B.n365 71.676
R1159 B.n363 B.n362 71.676
R1160 B.n358 B.n357 71.676
R1161 B.n355 B.n354 71.676
R1162 B.n350 B.n349 71.676
R1163 B.n347 B.n346 71.676
R1164 B.n342 B.n341 71.676
R1165 B.n339 B.n338 71.676
R1166 B.n334 B.n333 71.676
R1167 B.n331 B.n330 71.676
R1168 B.n326 B.n325 71.676
R1169 B.n323 B.n322 71.676
R1170 B.n318 B.n317 71.676
R1171 B.n315 B.n314 71.676
R1172 B.n310 B.n309 71.676
R1173 B.n307 B.n306 71.676
R1174 B.n302 B.n301 71.676
R1175 B.n299 B.n298 71.676
R1176 B.n294 B.n293 71.676
R1177 B.n291 B.n290 71.676
R1178 B.n286 B.n285 71.676
R1179 B.n283 B.n282 71.676
R1180 B.n278 B.n277 71.676
R1181 B.n275 B.n274 71.676
R1182 B.n270 B.n269 71.676
R1183 B.n267 B.n197 71.676
R1184 B.n237 B.t10 71.1345
R1185 B.n104 B.t18 71.1345
R1186 B.n231 B.t20 71.1108
R1187 B.n97 B.t15 71.1108
R1188 B.n384 B.n237 59.5399
R1189 B.n402 B.n231 59.5399
R1190 B.n98 B.n97 59.5399
R1191 B.n785 B.n104 59.5399
R1192 B.n522 B.n198 53.6822
R1193 B.n924 B.n64 53.6822
R1194 B.n237 B.n236 33.9399
R1195 B.n231 B.n230 33.9399
R1196 B.n97 B.n96 33.9399
R1197 B.n104 B.n103 33.9399
R1198 B.n922 B.n921 32.9371
R1199 B.n667 B.n666 32.9371
R1200 B.n524 B.n196 32.9371
R1201 B.n520 B.n519 32.9371
R1202 B.n522 B.n194 32.3045
R1203 B.n528 B.n194 32.3045
R1204 B.n528 B.n190 32.3045
R1205 B.n534 B.n190 32.3045
R1206 B.n534 B.n186 32.3045
R1207 B.n540 B.n186 32.3045
R1208 B.n546 B.n182 32.3045
R1209 B.n546 B.n178 32.3045
R1210 B.n552 B.n178 32.3045
R1211 B.n552 B.n174 32.3045
R1212 B.n558 B.n174 32.3045
R1213 B.n558 B.n170 32.3045
R1214 B.n564 B.n170 32.3045
R1215 B.n570 B.n166 32.3045
R1216 B.n570 B.n162 32.3045
R1217 B.n577 B.n162 32.3045
R1218 B.n577 B.n576 32.3045
R1219 B.n583 B.n155 32.3045
R1220 B.n589 B.n155 32.3045
R1221 B.n589 B.n151 32.3045
R1222 B.n595 B.n151 32.3045
R1223 B.n601 B.n147 32.3045
R1224 B.n601 B.n142 32.3045
R1225 B.n607 B.n142 32.3045
R1226 B.n607 B.n143 32.3045
R1227 B.n614 B.n135 32.3045
R1228 B.n620 B.n135 32.3045
R1229 B.n620 B.n4 32.3045
R1230 B.n990 B.n4 32.3045
R1231 B.n990 B.n989 32.3045
R1232 B.n989 B.n988 32.3045
R1233 B.n988 B.n8 32.3045
R1234 B.n982 B.n8 32.3045
R1235 B.n981 B.n980 32.3045
R1236 B.n980 B.n15 32.3045
R1237 B.n974 B.n15 32.3045
R1238 B.n974 B.n973 32.3045
R1239 B.n972 B.n22 32.3045
R1240 B.n966 B.n22 32.3045
R1241 B.n966 B.n965 32.3045
R1242 B.n965 B.n964 32.3045
R1243 B.n958 B.n32 32.3045
R1244 B.n958 B.n957 32.3045
R1245 B.n957 B.n956 32.3045
R1246 B.n956 B.n36 32.3045
R1247 B.n950 B.n949 32.3045
R1248 B.n949 B.n948 32.3045
R1249 B.n948 B.n43 32.3045
R1250 B.n942 B.n43 32.3045
R1251 B.n942 B.n941 32.3045
R1252 B.n941 B.n940 32.3045
R1253 B.n940 B.n50 32.3045
R1254 B.n934 B.n933 32.3045
R1255 B.n933 B.n932 32.3045
R1256 B.n932 B.n57 32.3045
R1257 B.n926 B.n57 32.3045
R1258 B.n926 B.n925 32.3045
R1259 B.n925 B.n924 32.3045
R1260 B.t9 B.n182 31.3544
R1261 B.t13 B.n50 31.3544
R1262 B.n143 B.t7 26.6038
R1263 B.t4 B.n981 26.6038
R1264 B.n595 B.t1 21.8532
R1265 B.t2 B.n972 21.8532
R1266 B.t0 B.n166 19.953
R1267 B.t3 B.n36 19.953
R1268 B B.n992 18.0485
R1269 B.n576 B.t6 17.1026
R1270 B.n32 B.t5 17.1026
R1271 B.n583 B.t6 15.2024
R1272 B.n964 B.t5 15.2024
R1273 B.n564 B.t0 12.352
R1274 B.n950 B.t3 12.352
R1275 B.n921 B.n920 10.6151
R1276 B.n920 B.n66 10.6151
R1277 B.n914 B.n66 10.6151
R1278 B.n914 B.n913 10.6151
R1279 B.n913 B.n912 10.6151
R1280 B.n912 B.n68 10.6151
R1281 B.n906 B.n68 10.6151
R1282 B.n906 B.n905 10.6151
R1283 B.n905 B.n904 10.6151
R1284 B.n904 B.n70 10.6151
R1285 B.n898 B.n70 10.6151
R1286 B.n898 B.n897 10.6151
R1287 B.n897 B.n896 10.6151
R1288 B.n896 B.n72 10.6151
R1289 B.n890 B.n72 10.6151
R1290 B.n890 B.n889 10.6151
R1291 B.n889 B.n888 10.6151
R1292 B.n888 B.n74 10.6151
R1293 B.n882 B.n74 10.6151
R1294 B.n882 B.n881 10.6151
R1295 B.n881 B.n880 10.6151
R1296 B.n880 B.n76 10.6151
R1297 B.n874 B.n76 10.6151
R1298 B.n874 B.n873 10.6151
R1299 B.n873 B.n872 10.6151
R1300 B.n872 B.n78 10.6151
R1301 B.n866 B.n78 10.6151
R1302 B.n866 B.n865 10.6151
R1303 B.n865 B.n864 10.6151
R1304 B.n864 B.n80 10.6151
R1305 B.n858 B.n80 10.6151
R1306 B.n858 B.n857 10.6151
R1307 B.n857 B.n856 10.6151
R1308 B.n856 B.n82 10.6151
R1309 B.n850 B.n82 10.6151
R1310 B.n850 B.n849 10.6151
R1311 B.n849 B.n848 10.6151
R1312 B.n848 B.n84 10.6151
R1313 B.n842 B.n84 10.6151
R1314 B.n842 B.n841 10.6151
R1315 B.n841 B.n840 10.6151
R1316 B.n840 B.n86 10.6151
R1317 B.n834 B.n86 10.6151
R1318 B.n834 B.n833 10.6151
R1319 B.n833 B.n832 10.6151
R1320 B.n832 B.n88 10.6151
R1321 B.n826 B.n88 10.6151
R1322 B.n826 B.n825 10.6151
R1323 B.n825 B.n824 10.6151
R1324 B.n824 B.n90 10.6151
R1325 B.n818 B.n90 10.6151
R1326 B.n818 B.n817 10.6151
R1327 B.n817 B.n816 10.6151
R1328 B.n816 B.n92 10.6151
R1329 B.n810 B.n92 10.6151
R1330 B.n810 B.n809 10.6151
R1331 B.n809 B.n808 10.6151
R1332 B.n808 B.n94 10.6151
R1333 B.n802 B.n801 10.6151
R1334 B.n801 B.n800 10.6151
R1335 B.n800 B.n99 10.6151
R1336 B.n794 B.n99 10.6151
R1337 B.n794 B.n793 10.6151
R1338 B.n793 B.n792 10.6151
R1339 B.n792 B.n101 10.6151
R1340 B.n786 B.n101 10.6151
R1341 B.n784 B.n783 10.6151
R1342 B.n783 B.n105 10.6151
R1343 B.n777 B.n105 10.6151
R1344 B.n777 B.n776 10.6151
R1345 B.n776 B.n775 10.6151
R1346 B.n775 B.n107 10.6151
R1347 B.n769 B.n107 10.6151
R1348 B.n769 B.n768 10.6151
R1349 B.n768 B.n767 10.6151
R1350 B.n767 B.n109 10.6151
R1351 B.n761 B.n109 10.6151
R1352 B.n761 B.n760 10.6151
R1353 B.n760 B.n759 10.6151
R1354 B.n759 B.n111 10.6151
R1355 B.n753 B.n111 10.6151
R1356 B.n753 B.n752 10.6151
R1357 B.n752 B.n751 10.6151
R1358 B.n751 B.n113 10.6151
R1359 B.n745 B.n113 10.6151
R1360 B.n745 B.n744 10.6151
R1361 B.n744 B.n743 10.6151
R1362 B.n743 B.n115 10.6151
R1363 B.n737 B.n115 10.6151
R1364 B.n737 B.n736 10.6151
R1365 B.n736 B.n735 10.6151
R1366 B.n735 B.n117 10.6151
R1367 B.n729 B.n117 10.6151
R1368 B.n729 B.n728 10.6151
R1369 B.n728 B.n727 10.6151
R1370 B.n727 B.n119 10.6151
R1371 B.n721 B.n119 10.6151
R1372 B.n721 B.n720 10.6151
R1373 B.n720 B.n719 10.6151
R1374 B.n719 B.n121 10.6151
R1375 B.n713 B.n121 10.6151
R1376 B.n713 B.n712 10.6151
R1377 B.n712 B.n711 10.6151
R1378 B.n711 B.n123 10.6151
R1379 B.n705 B.n123 10.6151
R1380 B.n705 B.n704 10.6151
R1381 B.n704 B.n703 10.6151
R1382 B.n703 B.n125 10.6151
R1383 B.n697 B.n125 10.6151
R1384 B.n697 B.n696 10.6151
R1385 B.n696 B.n695 10.6151
R1386 B.n695 B.n127 10.6151
R1387 B.n689 B.n127 10.6151
R1388 B.n689 B.n688 10.6151
R1389 B.n688 B.n687 10.6151
R1390 B.n687 B.n129 10.6151
R1391 B.n681 B.n129 10.6151
R1392 B.n681 B.n680 10.6151
R1393 B.n680 B.n679 10.6151
R1394 B.n679 B.n131 10.6151
R1395 B.n673 B.n131 10.6151
R1396 B.n673 B.n672 10.6151
R1397 B.n672 B.n671 10.6151
R1398 B.n671 B.n667 10.6151
R1399 B.n525 B.n524 10.6151
R1400 B.n526 B.n525 10.6151
R1401 B.n526 B.n188 10.6151
R1402 B.n536 B.n188 10.6151
R1403 B.n537 B.n536 10.6151
R1404 B.n538 B.n537 10.6151
R1405 B.n538 B.n180 10.6151
R1406 B.n548 B.n180 10.6151
R1407 B.n549 B.n548 10.6151
R1408 B.n550 B.n549 10.6151
R1409 B.n550 B.n172 10.6151
R1410 B.n560 B.n172 10.6151
R1411 B.n561 B.n560 10.6151
R1412 B.n562 B.n561 10.6151
R1413 B.n562 B.n164 10.6151
R1414 B.n572 B.n164 10.6151
R1415 B.n573 B.n572 10.6151
R1416 B.n574 B.n573 10.6151
R1417 B.n574 B.n157 10.6151
R1418 B.n585 B.n157 10.6151
R1419 B.n586 B.n585 10.6151
R1420 B.n587 B.n586 10.6151
R1421 B.n587 B.n149 10.6151
R1422 B.n597 B.n149 10.6151
R1423 B.n598 B.n597 10.6151
R1424 B.n599 B.n598 10.6151
R1425 B.n599 B.n140 10.6151
R1426 B.n609 B.n140 10.6151
R1427 B.n610 B.n609 10.6151
R1428 B.n612 B.n610 10.6151
R1429 B.n612 B.n611 10.6151
R1430 B.n611 B.n133 10.6151
R1431 B.n623 B.n133 10.6151
R1432 B.n624 B.n623 10.6151
R1433 B.n625 B.n624 10.6151
R1434 B.n626 B.n625 10.6151
R1435 B.n628 B.n626 10.6151
R1436 B.n629 B.n628 10.6151
R1437 B.n630 B.n629 10.6151
R1438 B.n631 B.n630 10.6151
R1439 B.n633 B.n631 10.6151
R1440 B.n634 B.n633 10.6151
R1441 B.n635 B.n634 10.6151
R1442 B.n636 B.n635 10.6151
R1443 B.n638 B.n636 10.6151
R1444 B.n639 B.n638 10.6151
R1445 B.n640 B.n639 10.6151
R1446 B.n641 B.n640 10.6151
R1447 B.n643 B.n641 10.6151
R1448 B.n644 B.n643 10.6151
R1449 B.n645 B.n644 10.6151
R1450 B.n646 B.n645 10.6151
R1451 B.n648 B.n646 10.6151
R1452 B.n649 B.n648 10.6151
R1453 B.n650 B.n649 10.6151
R1454 B.n651 B.n650 10.6151
R1455 B.n653 B.n651 10.6151
R1456 B.n654 B.n653 10.6151
R1457 B.n655 B.n654 10.6151
R1458 B.n656 B.n655 10.6151
R1459 B.n658 B.n656 10.6151
R1460 B.n659 B.n658 10.6151
R1461 B.n660 B.n659 10.6151
R1462 B.n661 B.n660 10.6151
R1463 B.n663 B.n661 10.6151
R1464 B.n664 B.n663 10.6151
R1465 B.n665 B.n664 10.6151
R1466 B.n666 B.n665 10.6151
R1467 B.n519 B.n518 10.6151
R1468 B.n518 B.n200 10.6151
R1469 B.n513 B.n200 10.6151
R1470 B.n513 B.n512 10.6151
R1471 B.n512 B.n202 10.6151
R1472 B.n507 B.n202 10.6151
R1473 B.n507 B.n506 10.6151
R1474 B.n506 B.n505 10.6151
R1475 B.n505 B.n204 10.6151
R1476 B.n499 B.n204 10.6151
R1477 B.n499 B.n498 10.6151
R1478 B.n498 B.n497 10.6151
R1479 B.n497 B.n206 10.6151
R1480 B.n491 B.n206 10.6151
R1481 B.n491 B.n490 10.6151
R1482 B.n490 B.n489 10.6151
R1483 B.n489 B.n208 10.6151
R1484 B.n483 B.n208 10.6151
R1485 B.n483 B.n482 10.6151
R1486 B.n482 B.n481 10.6151
R1487 B.n481 B.n210 10.6151
R1488 B.n475 B.n210 10.6151
R1489 B.n475 B.n474 10.6151
R1490 B.n474 B.n473 10.6151
R1491 B.n473 B.n212 10.6151
R1492 B.n467 B.n212 10.6151
R1493 B.n467 B.n466 10.6151
R1494 B.n466 B.n465 10.6151
R1495 B.n465 B.n214 10.6151
R1496 B.n459 B.n214 10.6151
R1497 B.n459 B.n458 10.6151
R1498 B.n458 B.n457 10.6151
R1499 B.n457 B.n216 10.6151
R1500 B.n451 B.n216 10.6151
R1501 B.n451 B.n450 10.6151
R1502 B.n450 B.n449 10.6151
R1503 B.n449 B.n218 10.6151
R1504 B.n443 B.n218 10.6151
R1505 B.n443 B.n442 10.6151
R1506 B.n442 B.n441 10.6151
R1507 B.n441 B.n220 10.6151
R1508 B.n435 B.n220 10.6151
R1509 B.n435 B.n434 10.6151
R1510 B.n434 B.n433 10.6151
R1511 B.n433 B.n222 10.6151
R1512 B.n427 B.n222 10.6151
R1513 B.n427 B.n426 10.6151
R1514 B.n426 B.n425 10.6151
R1515 B.n425 B.n224 10.6151
R1516 B.n419 B.n224 10.6151
R1517 B.n419 B.n418 10.6151
R1518 B.n418 B.n417 10.6151
R1519 B.n417 B.n226 10.6151
R1520 B.n411 B.n226 10.6151
R1521 B.n411 B.n410 10.6151
R1522 B.n410 B.n409 10.6151
R1523 B.n409 B.n228 10.6151
R1524 B.n403 B.n228 10.6151
R1525 B.n401 B.n400 10.6151
R1526 B.n400 B.n232 10.6151
R1527 B.n394 B.n232 10.6151
R1528 B.n394 B.n393 10.6151
R1529 B.n393 B.n392 10.6151
R1530 B.n392 B.n234 10.6151
R1531 B.n386 B.n234 10.6151
R1532 B.n386 B.n385 10.6151
R1533 B.n383 B.n238 10.6151
R1534 B.n377 B.n238 10.6151
R1535 B.n377 B.n376 10.6151
R1536 B.n376 B.n375 10.6151
R1537 B.n375 B.n240 10.6151
R1538 B.n369 B.n240 10.6151
R1539 B.n369 B.n368 10.6151
R1540 B.n368 B.n367 10.6151
R1541 B.n367 B.n242 10.6151
R1542 B.n361 B.n242 10.6151
R1543 B.n361 B.n360 10.6151
R1544 B.n360 B.n359 10.6151
R1545 B.n359 B.n244 10.6151
R1546 B.n353 B.n244 10.6151
R1547 B.n353 B.n352 10.6151
R1548 B.n352 B.n351 10.6151
R1549 B.n351 B.n246 10.6151
R1550 B.n345 B.n246 10.6151
R1551 B.n345 B.n344 10.6151
R1552 B.n344 B.n343 10.6151
R1553 B.n343 B.n248 10.6151
R1554 B.n337 B.n248 10.6151
R1555 B.n337 B.n336 10.6151
R1556 B.n336 B.n335 10.6151
R1557 B.n335 B.n250 10.6151
R1558 B.n329 B.n250 10.6151
R1559 B.n329 B.n328 10.6151
R1560 B.n328 B.n327 10.6151
R1561 B.n327 B.n252 10.6151
R1562 B.n321 B.n252 10.6151
R1563 B.n321 B.n320 10.6151
R1564 B.n320 B.n319 10.6151
R1565 B.n319 B.n254 10.6151
R1566 B.n313 B.n254 10.6151
R1567 B.n313 B.n312 10.6151
R1568 B.n312 B.n311 10.6151
R1569 B.n311 B.n256 10.6151
R1570 B.n305 B.n256 10.6151
R1571 B.n305 B.n304 10.6151
R1572 B.n304 B.n303 10.6151
R1573 B.n303 B.n258 10.6151
R1574 B.n297 B.n258 10.6151
R1575 B.n297 B.n296 10.6151
R1576 B.n296 B.n295 10.6151
R1577 B.n295 B.n260 10.6151
R1578 B.n289 B.n260 10.6151
R1579 B.n289 B.n288 10.6151
R1580 B.n288 B.n287 10.6151
R1581 B.n287 B.n262 10.6151
R1582 B.n281 B.n262 10.6151
R1583 B.n281 B.n280 10.6151
R1584 B.n280 B.n279 10.6151
R1585 B.n279 B.n264 10.6151
R1586 B.n273 B.n264 10.6151
R1587 B.n273 B.n272 10.6151
R1588 B.n272 B.n271 10.6151
R1589 B.n271 B.n266 10.6151
R1590 B.n266 B.n196 10.6151
R1591 B.n520 B.n192 10.6151
R1592 B.n530 B.n192 10.6151
R1593 B.n531 B.n530 10.6151
R1594 B.n532 B.n531 10.6151
R1595 B.n532 B.n184 10.6151
R1596 B.n542 B.n184 10.6151
R1597 B.n543 B.n542 10.6151
R1598 B.n544 B.n543 10.6151
R1599 B.n544 B.n176 10.6151
R1600 B.n554 B.n176 10.6151
R1601 B.n555 B.n554 10.6151
R1602 B.n556 B.n555 10.6151
R1603 B.n556 B.n168 10.6151
R1604 B.n566 B.n168 10.6151
R1605 B.n567 B.n566 10.6151
R1606 B.n568 B.n567 10.6151
R1607 B.n568 B.n160 10.6151
R1608 B.n579 B.n160 10.6151
R1609 B.n580 B.n579 10.6151
R1610 B.n581 B.n580 10.6151
R1611 B.n581 B.n153 10.6151
R1612 B.n591 B.n153 10.6151
R1613 B.n592 B.n591 10.6151
R1614 B.n593 B.n592 10.6151
R1615 B.n593 B.n145 10.6151
R1616 B.n603 B.n145 10.6151
R1617 B.n604 B.n603 10.6151
R1618 B.n605 B.n604 10.6151
R1619 B.n605 B.n137 10.6151
R1620 B.n616 B.n137 10.6151
R1621 B.n617 B.n616 10.6151
R1622 B.n618 B.n617 10.6151
R1623 B.n618 B.n0 10.6151
R1624 B.n986 B.n1 10.6151
R1625 B.n986 B.n985 10.6151
R1626 B.n985 B.n984 10.6151
R1627 B.n984 B.n10 10.6151
R1628 B.n978 B.n10 10.6151
R1629 B.n978 B.n977 10.6151
R1630 B.n977 B.n976 10.6151
R1631 B.n976 B.n17 10.6151
R1632 B.n970 B.n17 10.6151
R1633 B.n970 B.n969 10.6151
R1634 B.n969 B.n968 10.6151
R1635 B.n968 B.n24 10.6151
R1636 B.n962 B.n24 10.6151
R1637 B.n962 B.n961 10.6151
R1638 B.n961 B.n960 10.6151
R1639 B.n960 B.n30 10.6151
R1640 B.n954 B.n30 10.6151
R1641 B.n954 B.n953 10.6151
R1642 B.n953 B.n952 10.6151
R1643 B.n952 B.n38 10.6151
R1644 B.n946 B.n38 10.6151
R1645 B.n946 B.n945 10.6151
R1646 B.n945 B.n944 10.6151
R1647 B.n944 B.n45 10.6151
R1648 B.n938 B.n45 10.6151
R1649 B.n938 B.n937 10.6151
R1650 B.n937 B.n936 10.6151
R1651 B.n936 B.n52 10.6151
R1652 B.n930 B.n52 10.6151
R1653 B.n930 B.n929 10.6151
R1654 B.n929 B.n928 10.6151
R1655 B.n928 B.n59 10.6151
R1656 B.n922 B.n59 10.6151
R1657 B.t1 B.n147 10.4518
R1658 B.n973 B.t2 10.4518
R1659 B.n802 B.n98 6.5566
R1660 B.n786 B.n785 6.5566
R1661 B.n402 B.n401 6.5566
R1662 B.n385 B.n384 6.5566
R1663 B.n614 B.t7 5.70121
R1664 B.n982 B.t4 5.70121
R1665 B.n98 B.n94 4.05904
R1666 B.n785 B.n784 4.05904
R1667 B.n403 B.n402 4.05904
R1668 B.n384 B.n383 4.05904
R1669 B.n992 B.n0 2.81026
R1670 B.n992 B.n1 2.81026
R1671 B.n540 B.t9 0.950619
R1672 B.n934 B.t13 0.950619
R1673 VN.n5 VN.t7 335.183
R1674 VN.n24 VN.t5 335.183
R1675 VN.n4 VN.t1 303.457
R1676 VN.n10 VN.t0 303.457
R1677 VN.n17 VN.t6 303.457
R1678 VN.n23 VN.t2 303.457
R1679 VN.n29 VN.t4 303.457
R1680 VN.n36 VN.t3 303.457
R1681 VN.n18 VN.n17 179.744
R1682 VN.n37 VN.n36 179.744
R1683 VN.n35 VN.n19 161.3
R1684 VN.n34 VN.n33 161.3
R1685 VN.n32 VN.n20 161.3
R1686 VN.n31 VN.n30 161.3
R1687 VN.n28 VN.n21 161.3
R1688 VN.n27 VN.n26 161.3
R1689 VN.n25 VN.n22 161.3
R1690 VN.n16 VN.n0 161.3
R1691 VN.n15 VN.n14 161.3
R1692 VN.n13 VN.n1 161.3
R1693 VN.n12 VN.n11 161.3
R1694 VN.n9 VN.n2 161.3
R1695 VN.n8 VN.n7 161.3
R1696 VN.n6 VN.n3 161.3
R1697 VN.n15 VN.n1 56.5617
R1698 VN.n34 VN.n20 56.5617
R1699 VN VN.n37 50.0554
R1700 VN.n5 VN.n4 47.7556
R1701 VN.n24 VN.n23 47.7556
R1702 VN.n8 VN.n3 40.577
R1703 VN.n9 VN.n8 40.577
R1704 VN.n27 VN.n22 40.577
R1705 VN.n28 VN.n27 40.577
R1706 VN.n11 VN.n1 24.5923
R1707 VN.n16 VN.n15 24.5923
R1708 VN.n30 VN.n20 24.5923
R1709 VN.n35 VN.n34 24.5923
R1710 VN.n4 VN.n3 18.4444
R1711 VN.n10 VN.n9 18.4444
R1712 VN.n23 VN.n22 18.4444
R1713 VN.n29 VN.n28 18.4444
R1714 VN.n25 VN.n24 18.1442
R1715 VN.n6 VN.n5 18.1442
R1716 VN.n11 VN.n10 6.14846
R1717 VN.n17 VN.n16 6.14846
R1718 VN.n30 VN.n29 6.14846
R1719 VN.n36 VN.n35 6.14846
R1720 VN.n37 VN.n19 0.189894
R1721 VN.n33 VN.n19 0.189894
R1722 VN.n33 VN.n32 0.189894
R1723 VN.n32 VN.n31 0.189894
R1724 VN.n31 VN.n21 0.189894
R1725 VN.n26 VN.n21 0.189894
R1726 VN.n26 VN.n25 0.189894
R1727 VN.n7 VN.n6 0.189894
R1728 VN.n7 VN.n2 0.189894
R1729 VN.n12 VN.n2 0.189894
R1730 VN.n13 VN.n12 0.189894
R1731 VN.n14 VN.n13 0.189894
R1732 VN.n14 VN.n0 0.189894
R1733 VN.n18 VN.n0 0.189894
R1734 VN VN.n18 0.0516364
R1735 VDD2.n2 VDD2.n1 61.3627
R1736 VDD2.n2 VDD2.n0 61.3627
R1737 VDD2 VDD2.n5 61.3599
R1738 VDD2.n4 VDD2.n3 60.664
R1739 VDD2.n4 VDD2.n2 45.9179
R1740 VDD2.n5 VDD2.t0 1.10788
R1741 VDD2.n5 VDD2.t7 1.10788
R1742 VDD2.n3 VDD2.t4 1.10788
R1743 VDD2.n3 VDD2.t3 1.10788
R1744 VDD2.n1 VDD2.t2 1.10788
R1745 VDD2.n1 VDD2.t6 1.10788
R1746 VDD2.n0 VDD2.t5 1.10788
R1747 VDD2.n0 VDD2.t1 1.10788
R1748 VDD2 VDD2.n4 0.813
R1749 VTAIL.n11 VTAIL.t4 45.0926
R1750 VTAIL.n10 VTAIL.t10 45.0926
R1751 VTAIL.n7 VTAIL.t12 45.0926
R1752 VTAIL.n15 VTAIL.t9 45.0924
R1753 VTAIL.n2 VTAIL.t8 45.0924
R1754 VTAIL.n3 VTAIL.t6 45.0924
R1755 VTAIL.n6 VTAIL.t2 45.0924
R1756 VTAIL.n14 VTAIL.t1 45.0924
R1757 VTAIL.n13 VTAIL.n12 43.9852
R1758 VTAIL.n9 VTAIL.n8 43.9852
R1759 VTAIL.n1 VTAIL.n0 43.985
R1760 VTAIL.n5 VTAIL.n4 43.985
R1761 VTAIL.n15 VTAIL.n14 29.2893
R1762 VTAIL.n7 VTAIL.n6 29.2893
R1763 VTAIL.n9 VTAIL.n7 1.50912
R1764 VTAIL.n10 VTAIL.n9 1.50912
R1765 VTAIL.n13 VTAIL.n11 1.50912
R1766 VTAIL.n14 VTAIL.n13 1.50912
R1767 VTAIL.n6 VTAIL.n5 1.50912
R1768 VTAIL.n5 VTAIL.n3 1.50912
R1769 VTAIL.n2 VTAIL.n1 1.50912
R1770 VTAIL VTAIL.n15 1.45093
R1771 VTAIL.n0 VTAIL.t14 1.10788
R1772 VTAIL.n0 VTAIL.t15 1.10788
R1773 VTAIL.n4 VTAIL.t5 1.10788
R1774 VTAIL.n4 VTAIL.t3 1.10788
R1775 VTAIL.n12 VTAIL.t0 1.10788
R1776 VTAIL.n12 VTAIL.t7 1.10788
R1777 VTAIL.n8 VTAIL.t11 1.10788
R1778 VTAIL.n8 VTAIL.t13 1.10788
R1779 VTAIL.n11 VTAIL.n10 0.470328
R1780 VTAIL.n3 VTAIL.n2 0.470328
R1781 VTAIL VTAIL.n1 0.0586897
R1782 VP.n11 VP.t6 335.183
R1783 VP.n25 VP.t0 303.457
R1784 VP.n31 VP.t5 303.457
R1785 VP.n38 VP.t7 303.457
R1786 VP.n45 VP.t1 303.457
R1787 VP.n23 VP.t2 303.457
R1788 VP.n16 VP.t3 303.457
R1789 VP.n10 VP.t4 303.457
R1790 VP.n26 VP.n25 179.744
R1791 VP.n46 VP.n45 179.744
R1792 VP.n24 VP.n23 179.744
R1793 VP.n12 VP.n9 161.3
R1794 VP.n14 VP.n13 161.3
R1795 VP.n15 VP.n8 161.3
R1796 VP.n18 VP.n17 161.3
R1797 VP.n19 VP.n7 161.3
R1798 VP.n21 VP.n20 161.3
R1799 VP.n22 VP.n6 161.3
R1800 VP.n44 VP.n0 161.3
R1801 VP.n43 VP.n42 161.3
R1802 VP.n41 VP.n1 161.3
R1803 VP.n40 VP.n39 161.3
R1804 VP.n37 VP.n2 161.3
R1805 VP.n36 VP.n35 161.3
R1806 VP.n34 VP.n3 161.3
R1807 VP.n33 VP.n32 161.3
R1808 VP.n30 VP.n4 161.3
R1809 VP.n29 VP.n28 161.3
R1810 VP.n27 VP.n5 161.3
R1811 VP.n30 VP.n29 56.5617
R1812 VP.n43 VP.n1 56.5617
R1813 VP.n21 VP.n7 56.5617
R1814 VP.n26 VP.n24 49.6747
R1815 VP.n11 VP.n10 47.7556
R1816 VP.n36 VP.n3 40.577
R1817 VP.n37 VP.n36 40.577
R1818 VP.n15 VP.n14 40.577
R1819 VP.n14 VP.n9 40.577
R1820 VP.n29 VP.n5 24.5923
R1821 VP.n32 VP.n30 24.5923
R1822 VP.n39 VP.n1 24.5923
R1823 VP.n44 VP.n43 24.5923
R1824 VP.n22 VP.n21 24.5923
R1825 VP.n17 VP.n7 24.5923
R1826 VP.n31 VP.n3 18.4444
R1827 VP.n38 VP.n37 18.4444
R1828 VP.n16 VP.n15 18.4444
R1829 VP.n10 VP.n9 18.4444
R1830 VP.n12 VP.n11 18.1442
R1831 VP.n25 VP.n5 6.14846
R1832 VP.n32 VP.n31 6.14846
R1833 VP.n39 VP.n38 6.14846
R1834 VP.n45 VP.n44 6.14846
R1835 VP.n23 VP.n22 6.14846
R1836 VP.n17 VP.n16 6.14846
R1837 VP.n13 VP.n12 0.189894
R1838 VP.n13 VP.n8 0.189894
R1839 VP.n18 VP.n8 0.189894
R1840 VP.n19 VP.n18 0.189894
R1841 VP.n20 VP.n19 0.189894
R1842 VP.n20 VP.n6 0.189894
R1843 VP.n24 VP.n6 0.189894
R1844 VP.n27 VP.n26 0.189894
R1845 VP.n28 VP.n27 0.189894
R1846 VP.n28 VP.n4 0.189894
R1847 VP.n33 VP.n4 0.189894
R1848 VP.n34 VP.n33 0.189894
R1849 VP.n35 VP.n34 0.189894
R1850 VP.n35 VP.n2 0.189894
R1851 VP.n40 VP.n2 0.189894
R1852 VP.n41 VP.n40 0.189894
R1853 VP.n42 VP.n41 0.189894
R1854 VP.n42 VP.n0 0.189894
R1855 VP.n46 VP.n0 0.189894
R1856 VP VP.n46 0.0516364
R1857 VDD1 VDD1.n0 61.4765
R1858 VDD1.n3 VDD1.n2 61.3627
R1859 VDD1.n3 VDD1.n1 61.3627
R1860 VDD1.n5 VDD1.n4 60.6638
R1861 VDD1.n5 VDD1.n3 46.5009
R1862 VDD1.n4 VDD1.t4 1.10788
R1863 VDD1.n4 VDD1.t5 1.10788
R1864 VDD1.n0 VDD1.t1 1.10788
R1865 VDD1.n0 VDD1.t3 1.10788
R1866 VDD1.n2 VDD1.t0 1.10788
R1867 VDD1.n2 VDD1.t6 1.10788
R1868 VDD1.n1 VDD1.t7 1.10788
R1869 VDD1.n1 VDD1.t2 1.10788
R1870 VDD1 VDD1.n5 0.696621
C0 VDD1 VP 11.1103f
C1 VTAIL VN 10.6582f
C2 VDD1 VN 0.149993f
C3 VDD1 VTAIL 11.3946f
C4 VDD2 VP 0.394505f
C5 VDD2 VN 10.866599f
C6 VDD2 VTAIL 11.441099f
C7 VDD2 VDD1 1.18872f
C8 VN VP 7.30773f
C9 VTAIL VP 10.6723f
C10 VDD2 B 4.643646f
C11 VDD1 B 4.953212f
C12 VTAIL B 12.994035f
C13 VN B 11.68083f
C14 VP B 9.8514f
C15 VDD1.t1 B 0.356934f
C16 VDD1.t3 B 0.356934f
C17 VDD1.n0 B 3.25592f
C18 VDD1.t7 B 0.356934f
C19 VDD1.t2 B 0.356934f
C20 VDD1.n1 B 3.25507f
C21 VDD1.t0 B 0.356934f
C22 VDD1.t6 B 0.356934f
C23 VDD1.n2 B 3.25507f
C24 VDD1.n3 B 3.04827f
C25 VDD1.t4 B 0.356934f
C26 VDD1.t5 B 0.356934f
C27 VDD1.n4 B 3.2505f
C28 VDD1.n5 B 3.05313f
C29 VP.n0 B 0.031439f
C30 VP.t1 B 2.19527f
C31 VP.n1 B 0.045701f
C32 VP.n2 B 0.031439f
C33 VP.t7 B 2.19527f
C34 VP.n3 B 0.05496f
C35 VP.n4 B 0.031439f
C36 VP.n5 B 0.036714f
C37 VP.n6 B 0.031439f
C38 VP.t2 B 2.19527f
C39 VP.n7 B 0.045701f
C40 VP.n8 B 0.031439f
C41 VP.t3 B 2.19527f
C42 VP.n9 B 0.05496f
C43 VP.t6 B 2.27938f
C44 VP.t4 B 2.19527f
C45 VP.n10 B 0.837437f
C46 VP.n11 B 0.850024f
C47 VP.n12 B 0.194952f
C48 VP.n13 B 0.031439f
C49 VP.n14 B 0.025392f
C50 VP.n15 B 0.05496f
C51 VP.n16 B 0.774438f
C52 VP.n17 B 0.036714f
C53 VP.n18 B 0.031439f
C54 VP.n19 B 0.031439f
C55 VP.n20 B 0.031439f
C56 VP.n21 B 0.045701f
C57 VP.n22 B 0.036714f
C58 VP.n23 B 0.82908f
C59 VP.n24 B 1.69871f
C60 VP.t0 B 2.19527f
C61 VP.n25 B 0.82908f
C62 VP.n26 B 1.72153f
C63 VP.n27 B 0.031439f
C64 VP.n28 B 0.031439f
C65 VP.n29 B 0.045701f
C66 VP.n30 B 0.045701f
C67 VP.t5 B 2.19527f
C68 VP.n31 B 0.774438f
C69 VP.n32 B 0.036714f
C70 VP.n33 B 0.031439f
C71 VP.n34 B 0.031439f
C72 VP.n35 B 0.031439f
C73 VP.n36 B 0.025392f
C74 VP.n37 B 0.05496f
C75 VP.n38 B 0.774438f
C76 VP.n39 B 0.036714f
C77 VP.n40 B 0.031439f
C78 VP.n41 B 0.031439f
C79 VP.n42 B 0.031439f
C80 VP.n43 B 0.045701f
C81 VP.n44 B 0.036714f
C82 VP.n45 B 0.82908f
C83 VP.n46 B 0.030612f
C84 VTAIL.t14 B 0.25966f
C85 VTAIL.t15 B 0.25966f
C86 VTAIL.n0 B 2.30804f
C87 VTAIL.n1 B 0.277233f
C88 VTAIL.t8 B 2.94851f
C89 VTAIL.n2 B 0.369305f
C90 VTAIL.t6 B 2.94851f
C91 VTAIL.n3 B 0.369305f
C92 VTAIL.t5 B 0.25966f
C93 VTAIL.t3 B 0.25966f
C94 VTAIL.n4 B 2.30804f
C95 VTAIL.n5 B 0.363122f
C96 VTAIL.t2 B 2.94851f
C97 VTAIL.n6 B 1.5932f
C98 VTAIL.t12 B 2.94851f
C99 VTAIL.n7 B 1.5932f
C100 VTAIL.t11 B 0.25966f
C101 VTAIL.t13 B 0.25966f
C102 VTAIL.n8 B 2.30804f
C103 VTAIL.n9 B 0.363118f
C104 VTAIL.t10 B 2.94851f
C105 VTAIL.n10 B 0.369301f
C106 VTAIL.t4 B 2.94851f
C107 VTAIL.n11 B 0.369301f
C108 VTAIL.t0 B 0.25966f
C109 VTAIL.t7 B 0.25966f
C110 VTAIL.n12 B 2.30804f
C111 VTAIL.n13 B 0.363118f
C112 VTAIL.t1 B 2.94851f
C113 VTAIL.n14 B 1.5932f
C114 VTAIL.t9 B 2.94851f
C115 VTAIL.n15 B 1.58975f
C116 VDD2.t5 B 0.355235f
C117 VDD2.t1 B 0.355235f
C118 VDD2.n0 B 3.23957f
C119 VDD2.t2 B 0.355235f
C120 VDD2.t6 B 0.355235f
C121 VDD2.n1 B 3.23957f
C122 VDD2.n2 B 2.98095f
C123 VDD2.t4 B 0.355235f
C124 VDD2.t3 B 0.355235f
C125 VDD2.n3 B 3.23503f
C126 VDD2.n4 B 3.00796f
C127 VDD2.t0 B 0.355235f
C128 VDD2.t7 B 0.355235f
C129 VDD2.n5 B 3.23953f
C130 VN.n0 B 0.031175f
C131 VN.t6 B 2.17687f
C132 VN.n1 B 0.045318f
C133 VN.n2 B 0.031175f
C134 VN.t0 B 2.17687f
C135 VN.n3 B 0.054499f
C136 VN.t7 B 2.26028f
C137 VN.t1 B 2.17687f
C138 VN.n4 B 0.83042f
C139 VN.n5 B 0.842901f
C140 VN.n6 B 0.193319f
C141 VN.n7 B 0.031175f
C142 VN.n8 B 0.025179f
C143 VN.n9 B 0.054499f
C144 VN.n10 B 0.767949f
C145 VN.n11 B 0.036407f
C146 VN.n12 B 0.031175f
C147 VN.n13 B 0.031175f
C148 VN.n14 B 0.031175f
C149 VN.n15 B 0.045318f
C150 VN.n16 B 0.036407f
C151 VN.n17 B 0.822133f
C152 VN.n18 B 0.030355f
C153 VN.n19 B 0.031175f
C154 VN.t3 B 2.17687f
C155 VN.n20 B 0.045318f
C156 VN.n21 B 0.031175f
C157 VN.t4 B 2.17687f
C158 VN.n22 B 0.054499f
C159 VN.t5 B 2.26028f
C160 VN.t2 B 2.17687f
C161 VN.n23 B 0.83042f
C162 VN.n24 B 0.842901f
C163 VN.n25 B 0.193319f
C164 VN.n26 B 0.031175f
C165 VN.n27 B 0.025179f
C166 VN.n28 B 0.054499f
C167 VN.n29 B 0.767949f
C168 VN.n30 B 0.036407f
C169 VN.n31 B 0.031175f
C170 VN.n32 B 0.031175f
C171 VN.n33 B 0.031175f
C172 VN.n34 B 0.045318f
C173 VN.n35 B 0.036407f
C174 VN.n36 B 0.822133f
C175 VN.n37 B 1.70475f
.ends

