* NGSPICE file created from diff_pair_sample_0038.ext - technology: sky130A

.subckt diff_pair_sample_0038 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1978_n3580# sky130_fd_pr__pfet_01v8 ad=5.0934 pd=26.9 as=0 ps=0 w=13.06 l=0.93
X1 VTAIL.t11 VN.t0 VDD2.t0 w_n1978_n3580# sky130_fd_pr__pfet_01v8 ad=2.1549 pd=13.39 as=2.1549 ps=13.39 w=13.06 l=0.93
X2 VDD2.t3 VN.t1 VTAIL.t10 w_n1978_n3580# sky130_fd_pr__pfet_01v8 ad=5.0934 pd=26.9 as=2.1549 ps=13.39 w=13.06 l=0.93
X3 VDD2.t2 VN.t2 VTAIL.t9 w_n1978_n3580# sky130_fd_pr__pfet_01v8 ad=2.1549 pd=13.39 as=5.0934 ps=26.9 w=13.06 l=0.93
X4 VDD1.t5 VP.t0 VTAIL.t0 w_n1978_n3580# sky130_fd_pr__pfet_01v8 ad=2.1549 pd=13.39 as=5.0934 ps=26.9 w=13.06 l=0.93
X5 VTAIL.t5 VP.t1 VDD1.t4 w_n1978_n3580# sky130_fd_pr__pfet_01v8 ad=2.1549 pd=13.39 as=2.1549 ps=13.39 w=13.06 l=0.93
X6 VDD1.t3 VP.t2 VTAIL.t4 w_n1978_n3580# sky130_fd_pr__pfet_01v8 ad=5.0934 pd=26.9 as=2.1549 ps=13.39 w=13.06 l=0.93
X7 B.t8 B.t6 B.t7 w_n1978_n3580# sky130_fd_pr__pfet_01v8 ad=5.0934 pd=26.9 as=0 ps=0 w=13.06 l=0.93
X8 VDD2.t5 VN.t3 VTAIL.t8 w_n1978_n3580# sky130_fd_pr__pfet_01v8 ad=2.1549 pd=13.39 as=5.0934 ps=26.9 w=13.06 l=0.93
X9 VDD1.t2 VP.t3 VTAIL.t1 w_n1978_n3580# sky130_fd_pr__pfet_01v8 ad=2.1549 pd=13.39 as=5.0934 ps=26.9 w=13.06 l=0.93
X10 VDD1.t1 VP.t4 VTAIL.t2 w_n1978_n3580# sky130_fd_pr__pfet_01v8 ad=5.0934 pd=26.9 as=2.1549 ps=13.39 w=13.06 l=0.93
X11 VDD2.t4 VN.t4 VTAIL.t7 w_n1978_n3580# sky130_fd_pr__pfet_01v8 ad=5.0934 pd=26.9 as=2.1549 ps=13.39 w=13.06 l=0.93
X12 B.t5 B.t3 B.t4 w_n1978_n3580# sky130_fd_pr__pfet_01v8 ad=5.0934 pd=26.9 as=0 ps=0 w=13.06 l=0.93
X13 B.t2 B.t0 B.t1 w_n1978_n3580# sky130_fd_pr__pfet_01v8 ad=5.0934 pd=26.9 as=0 ps=0 w=13.06 l=0.93
X14 VTAIL.t3 VP.t5 VDD1.t0 w_n1978_n3580# sky130_fd_pr__pfet_01v8 ad=2.1549 pd=13.39 as=2.1549 ps=13.39 w=13.06 l=0.93
X15 VTAIL.t6 VN.t5 VDD2.t1 w_n1978_n3580# sky130_fd_pr__pfet_01v8 ad=2.1549 pd=13.39 as=2.1549 ps=13.39 w=13.06 l=0.93
R0 B.n410 B.n67 585
R1 B.n412 B.n411 585
R2 B.n413 B.n66 585
R3 B.n415 B.n414 585
R4 B.n416 B.n65 585
R5 B.n418 B.n417 585
R6 B.n419 B.n64 585
R7 B.n421 B.n420 585
R8 B.n422 B.n63 585
R9 B.n424 B.n423 585
R10 B.n425 B.n62 585
R11 B.n427 B.n426 585
R12 B.n428 B.n61 585
R13 B.n430 B.n429 585
R14 B.n431 B.n60 585
R15 B.n433 B.n432 585
R16 B.n434 B.n59 585
R17 B.n436 B.n435 585
R18 B.n437 B.n58 585
R19 B.n439 B.n438 585
R20 B.n440 B.n57 585
R21 B.n442 B.n441 585
R22 B.n443 B.n56 585
R23 B.n445 B.n444 585
R24 B.n446 B.n55 585
R25 B.n448 B.n447 585
R26 B.n449 B.n54 585
R27 B.n451 B.n450 585
R28 B.n452 B.n53 585
R29 B.n454 B.n453 585
R30 B.n455 B.n52 585
R31 B.n457 B.n456 585
R32 B.n458 B.n51 585
R33 B.n460 B.n459 585
R34 B.n461 B.n50 585
R35 B.n463 B.n462 585
R36 B.n464 B.n49 585
R37 B.n466 B.n465 585
R38 B.n467 B.n48 585
R39 B.n469 B.n468 585
R40 B.n470 B.n47 585
R41 B.n472 B.n471 585
R42 B.n473 B.n46 585
R43 B.n475 B.n474 585
R44 B.n476 B.n43 585
R45 B.n479 B.n478 585
R46 B.n480 B.n42 585
R47 B.n482 B.n481 585
R48 B.n483 B.n41 585
R49 B.n485 B.n484 585
R50 B.n486 B.n40 585
R51 B.n488 B.n487 585
R52 B.n489 B.n39 585
R53 B.n491 B.n490 585
R54 B.n493 B.n492 585
R55 B.n494 B.n35 585
R56 B.n496 B.n495 585
R57 B.n497 B.n34 585
R58 B.n499 B.n498 585
R59 B.n500 B.n33 585
R60 B.n502 B.n501 585
R61 B.n503 B.n32 585
R62 B.n505 B.n504 585
R63 B.n506 B.n31 585
R64 B.n508 B.n507 585
R65 B.n509 B.n30 585
R66 B.n511 B.n510 585
R67 B.n512 B.n29 585
R68 B.n514 B.n513 585
R69 B.n515 B.n28 585
R70 B.n517 B.n516 585
R71 B.n518 B.n27 585
R72 B.n520 B.n519 585
R73 B.n521 B.n26 585
R74 B.n523 B.n522 585
R75 B.n524 B.n25 585
R76 B.n526 B.n525 585
R77 B.n527 B.n24 585
R78 B.n529 B.n528 585
R79 B.n530 B.n23 585
R80 B.n532 B.n531 585
R81 B.n533 B.n22 585
R82 B.n535 B.n534 585
R83 B.n536 B.n21 585
R84 B.n538 B.n537 585
R85 B.n539 B.n20 585
R86 B.n541 B.n540 585
R87 B.n542 B.n19 585
R88 B.n544 B.n543 585
R89 B.n545 B.n18 585
R90 B.n547 B.n546 585
R91 B.n548 B.n17 585
R92 B.n550 B.n549 585
R93 B.n551 B.n16 585
R94 B.n553 B.n552 585
R95 B.n554 B.n15 585
R96 B.n556 B.n555 585
R97 B.n557 B.n14 585
R98 B.n559 B.n558 585
R99 B.n409 B.n408 585
R100 B.n407 B.n68 585
R101 B.n406 B.n405 585
R102 B.n404 B.n69 585
R103 B.n403 B.n402 585
R104 B.n401 B.n70 585
R105 B.n400 B.n399 585
R106 B.n398 B.n71 585
R107 B.n397 B.n396 585
R108 B.n395 B.n72 585
R109 B.n394 B.n393 585
R110 B.n392 B.n73 585
R111 B.n391 B.n390 585
R112 B.n389 B.n74 585
R113 B.n388 B.n387 585
R114 B.n386 B.n75 585
R115 B.n385 B.n384 585
R116 B.n383 B.n76 585
R117 B.n382 B.n381 585
R118 B.n380 B.n77 585
R119 B.n379 B.n378 585
R120 B.n377 B.n78 585
R121 B.n376 B.n375 585
R122 B.n374 B.n79 585
R123 B.n373 B.n372 585
R124 B.n371 B.n80 585
R125 B.n370 B.n369 585
R126 B.n368 B.n81 585
R127 B.n367 B.n366 585
R128 B.n365 B.n82 585
R129 B.n364 B.n363 585
R130 B.n362 B.n83 585
R131 B.n361 B.n360 585
R132 B.n359 B.n84 585
R133 B.n358 B.n357 585
R134 B.n356 B.n85 585
R135 B.n355 B.n354 585
R136 B.n353 B.n86 585
R137 B.n352 B.n351 585
R138 B.n350 B.n87 585
R139 B.n349 B.n348 585
R140 B.n347 B.n88 585
R141 B.n346 B.n345 585
R142 B.n344 B.n89 585
R143 B.n343 B.n342 585
R144 B.n341 B.n90 585
R145 B.n340 B.n339 585
R146 B.n190 B.n189 585
R147 B.n191 B.n144 585
R148 B.n193 B.n192 585
R149 B.n194 B.n143 585
R150 B.n196 B.n195 585
R151 B.n197 B.n142 585
R152 B.n199 B.n198 585
R153 B.n200 B.n141 585
R154 B.n202 B.n201 585
R155 B.n203 B.n140 585
R156 B.n205 B.n204 585
R157 B.n206 B.n139 585
R158 B.n208 B.n207 585
R159 B.n209 B.n138 585
R160 B.n211 B.n210 585
R161 B.n212 B.n137 585
R162 B.n214 B.n213 585
R163 B.n215 B.n136 585
R164 B.n217 B.n216 585
R165 B.n218 B.n135 585
R166 B.n220 B.n219 585
R167 B.n221 B.n134 585
R168 B.n223 B.n222 585
R169 B.n224 B.n133 585
R170 B.n226 B.n225 585
R171 B.n227 B.n132 585
R172 B.n229 B.n228 585
R173 B.n230 B.n131 585
R174 B.n232 B.n231 585
R175 B.n233 B.n130 585
R176 B.n235 B.n234 585
R177 B.n236 B.n129 585
R178 B.n238 B.n237 585
R179 B.n239 B.n128 585
R180 B.n241 B.n240 585
R181 B.n242 B.n127 585
R182 B.n244 B.n243 585
R183 B.n245 B.n126 585
R184 B.n247 B.n246 585
R185 B.n248 B.n125 585
R186 B.n250 B.n249 585
R187 B.n251 B.n124 585
R188 B.n253 B.n252 585
R189 B.n254 B.n123 585
R190 B.n256 B.n255 585
R191 B.n258 B.n257 585
R192 B.n259 B.n119 585
R193 B.n261 B.n260 585
R194 B.n262 B.n118 585
R195 B.n264 B.n263 585
R196 B.n265 B.n117 585
R197 B.n267 B.n266 585
R198 B.n268 B.n116 585
R199 B.n270 B.n269 585
R200 B.n272 B.n113 585
R201 B.n274 B.n273 585
R202 B.n275 B.n112 585
R203 B.n277 B.n276 585
R204 B.n278 B.n111 585
R205 B.n280 B.n279 585
R206 B.n281 B.n110 585
R207 B.n283 B.n282 585
R208 B.n284 B.n109 585
R209 B.n286 B.n285 585
R210 B.n287 B.n108 585
R211 B.n289 B.n288 585
R212 B.n290 B.n107 585
R213 B.n292 B.n291 585
R214 B.n293 B.n106 585
R215 B.n295 B.n294 585
R216 B.n296 B.n105 585
R217 B.n298 B.n297 585
R218 B.n299 B.n104 585
R219 B.n301 B.n300 585
R220 B.n302 B.n103 585
R221 B.n304 B.n303 585
R222 B.n305 B.n102 585
R223 B.n307 B.n306 585
R224 B.n308 B.n101 585
R225 B.n310 B.n309 585
R226 B.n311 B.n100 585
R227 B.n313 B.n312 585
R228 B.n314 B.n99 585
R229 B.n316 B.n315 585
R230 B.n317 B.n98 585
R231 B.n319 B.n318 585
R232 B.n320 B.n97 585
R233 B.n322 B.n321 585
R234 B.n323 B.n96 585
R235 B.n325 B.n324 585
R236 B.n326 B.n95 585
R237 B.n328 B.n327 585
R238 B.n329 B.n94 585
R239 B.n331 B.n330 585
R240 B.n332 B.n93 585
R241 B.n334 B.n333 585
R242 B.n335 B.n92 585
R243 B.n337 B.n336 585
R244 B.n338 B.n91 585
R245 B.n188 B.n145 585
R246 B.n187 B.n186 585
R247 B.n185 B.n146 585
R248 B.n184 B.n183 585
R249 B.n182 B.n147 585
R250 B.n181 B.n180 585
R251 B.n179 B.n148 585
R252 B.n178 B.n177 585
R253 B.n176 B.n149 585
R254 B.n175 B.n174 585
R255 B.n173 B.n150 585
R256 B.n172 B.n171 585
R257 B.n170 B.n151 585
R258 B.n169 B.n168 585
R259 B.n167 B.n152 585
R260 B.n166 B.n165 585
R261 B.n164 B.n153 585
R262 B.n163 B.n162 585
R263 B.n161 B.n154 585
R264 B.n160 B.n159 585
R265 B.n158 B.n155 585
R266 B.n157 B.n156 585
R267 B.n2 B.n0 585
R268 B.n593 B.n1 585
R269 B.n592 B.n591 585
R270 B.n590 B.n3 585
R271 B.n589 B.n588 585
R272 B.n587 B.n4 585
R273 B.n586 B.n585 585
R274 B.n584 B.n5 585
R275 B.n583 B.n582 585
R276 B.n581 B.n6 585
R277 B.n580 B.n579 585
R278 B.n578 B.n7 585
R279 B.n577 B.n576 585
R280 B.n575 B.n8 585
R281 B.n574 B.n573 585
R282 B.n572 B.n9 585
R283 B.n571 B.n570 585
R284 B.n569 B.n10 585
R285 B.n568 B.n567 585
R286 B.n566 B.n11 585
R287 B.n565 B.n564 585
R288 B.n563 B.n12 585
R289 B.n562 B.n561 585
R290 B.n560 B.n13 585
R291 B.n595 B.n594 585
R292 B.n114 B.t0 540.864
R293 B.n120 B.t9 540.864
R294 B.n36 B.t3 540.864
R295 B.n44 B.t6 540.864
R296 B.n190 B.n145 492.5
R297 B.n558 B.n13 492.5
R298 B.n340 B.n91 492.5
R299 B.n408 B.n67 492.5
R300 B.n186 B.n145 163.367
R301 B.n186 B.n185 163.367
R302 B.n185 B.n184 163.367
R303 B.n184 B.n147 163.367
R304 B.n180 B.n147 163.367
R305 B.n180 B.n179 163.367
R306 B.n179 B.n178 163.367
R307 B.n178 B.n149 163.367
R308 B.n174 B.n149 163.367
R309 B.n174 B.n173 163.367
R310 B.n173 B.n172 163.367
R311 B.n172 B.n151 163.367
R312 B.n168 B.n151 163.367
R313 B.n168 B.n167 163.367
R314 B.n167 B.n166 163.367
R315 B.n166 B.n153 163.367
R316 B.n162 B.n153 163.367
R317 B.n162 B.n161 163.367
R318 B.n161 B.n160 163.367
R319 B.n160 B.n155 163.367
R320 B.n156 B.n155 163.367
R321 B.n156 B.n2 163.367
R322 B.n594 B.n2 163.367
R323 B.n594 B.n593 163.367
R324 B.n593 B.n592 163.367
R325 B.n592 B.n3 163.367
R326 B.n588 B.n3 163.367
R327 B.n588 B.n587 163.367
R328 B.n587 B.n586 163.367
R329 B.n586 B.n5 163.367
R330 B.n582 B.n5 163.367
R331 B.n582 B.n581 163.367
R332 B.n581 B.n580 163.367
R333 B.n580 B.n7 163.367
R334 B.n576 B.n7 163.367
R335 B.n576 B.n575 163.367
R336 B.n575 B.n574 163.367
R337 B.n574 B.n9 163.367
R338 B.n570 B.n9 163.367
R339 B.n570 B.n569 163.367
R340 B.n569 B.n568 163.367
R341 B.n568 B.n11 163.367
R342 B.n564 B.n11 163.367
R343 B.n564 B.n563 163.367
R344 B.n563 B.n562 163.367
R345 B.n562 B.n13 163.367
R346 B.n191 B.n190 163.367
R347 B.n192 B.n191 163.367
R348 B.n192 B.n143 163.367
R349 B.n196 B.n143 163.367
R350 B.n197 B.n196 163.367
R351 B.n198 B.n197 163.367
R352 B.n198 B.n141 163.367
R353 B.n202 B.n141 163.367
R354 B.n203 B.n202 163.367
R355 B.n204 B.n203 163.367
R356 B.n204 B.n139 163.367
R357 B.n208 B.n139 163.367
R358 B.n209 B.n208 163.367
R359 B.n210 B.n209 163.367
R360 B.n210 B.n137 163.367
R361 B.n214 B.n137 163.367
R362 B.n215 B.n214 163.367
R363 B.n216 B.n215 163.367
R364 B.n216 B.n135 163.367
R365 B.n220 B.n135 163.367
R366 B.n221 B.n220 163.367
R367 B.n222 B.n221 163.367
R368 B.n222 B.n133 163.367
R369 B.n226 B.n133 163.367
R370 B.n227 B.n226 163.367
R371 B.n228 B.n227 163.367
R372 B.n228 B.n131 163.367
R373 B.n232 B.n131 163.367
R374 B.n233 B.n232 163.367
R375 B.n234 B.n233 163.367
R376 B.n234 B.n129 163.367
R377 B.n238 B.n129 163.367
R378 B.n239 B.n238 163.367
R379 B.n240 B.n239 163.367
R380 B.n240 B.n127 163.367
R381 B.n244 B.n127 163.367
R382 B.n245 B.n244 163.367
R383 B.n246 B.n245 163.367
R384 B.n246 B.n125 163.367
R385 B.n250 B.n125 163.367
R386 B.n251 B.n250 163.367
R387 B.n252 B.n251 163.367
R388 B.n252 B.n123 163.367
R389 B.n256 B.n123 163.367
R390 B.n257 B.n256 163.367
R391 B.n257 B.n119 163.367
R392 B.n261 B.n119 163.367
R393 B.n262 B.n261 163.367
R394 B.n263 B.n262 163.367
R395 B.n263 B.n117 163.367
R396 B.n267 B.n117 163.367
R397 B.n268 B.n267 163.367
R398 B.n269 B.n268 163.367
R399 B.n269 B.n113 163.367
R400 B.n274 B.n113 163.367
R401 B.n275 B.n274 163.367
R402 B.n276 B.n275 163.367
R403 B.n276 B.n111 163.367
R404 B.n280 B.n111 163.367
R405 B.n281 B.n280 163.367
R406 B.n282 B.n281 163.367
R407 B.n282 B.n109 163.367
R408 B.n286 B.n109 163.367
R409 B.n287 B.n286 163.367
R410 B.n288 B.n287 163.367
R411 B.n288 B.n107 163.367
R412 B.n292 B.n107 163.367
R413 B.n293 B.n292 163.367
R414 B.n294 B.n293 163.367
R415 B.n294 B.n105 163.367
R416 B.n298 B.n105 163.367
R417 B.n299 B.n298 163.367
R418 B.n300 B.n299 163.367
R419 B.n300 B.n103 163.367
R420 B.n304 B.n103 163.367
R421 B.n305 B.n304 163.367
R422 B.n306 B.n305 163.367
R423 B.n306 B.n101 163.367
R424 B.n310 B.n101 163.367
R425 B.n311 B.n310 163.367
R426 B.n312 B.n311 163.367
R427 B.n312 B.n99 163.367
R428 B.n316 B.n99 163.367
R429 B.n317 B.n316 163.367
R430 B.n318 B.n317 163.367
R431 B.n318 B.n97 163.367
R432 B.n322 B.n97 163.367
R433 B.n323 B.n322 163.367
R434 B.n324 B.n323 163.367
R435 B.n324 B.n95 163.367
R436 B.n328 B.n95 163.367
R437 B.n329 B.n328 163.367
R438 B.n330 B.n329 163.367
R439 B.n330 B.n93 163.367
R440 B.n334 B.n93 163.367
R441 B.n335 B.n334 163.367
R442 B.n336 B.n335 163.367
R443 B.n336 B.n91 163.367
R444 B.n341 B.n340 163.367
R445 B.n342 B.n341 163.367
R446 B.n342 B.n89 163.367
R447 B.n346 B.n89 163.367
R448 B.n347 B.n346 163.367
R449 B.n348 B.n347 163.367
R450 B.n348 B.n87 163.367
R451 B.n352 B.n87 163.367
R452 B.n353 B.n352 163.367
R453 B.n354 B.n353 163.367
R454 B.n354 B.n85 163.367
R455 B.n358 B.n85 163.367
R456 B.n359 B.n358 163.367
R457 B.n360 B.n359 163.367
R458 B.n360 B.n83 163.367
R459 B.n364 B.n83 163.367
R460 B.n365 B.n364 163.367
R461 B.n366 B.n365 163.367
R462 B.n366 B.n81 163.367
R463 B.n370 B.n81 163.367
R464 B.n371 B.n370 163.367
R465 B.n372 B.n371 163.367
R466 B.n372 B.n79 163.367
R467 B.n376 B.n79 163.367
R468 B.n377 B.n376 163.367
R469 B.n378 B.n377 163.367
R470 B.n378 B.n77 163.367
R471 B.n382 B.n77 163.367
R472 B.n383 B.n382 163.367
R473 B.n384 B.n383 163.367
R474 B.n384 B.n75 163.367
R475 B.n388 B.n75 163.367
R476 B.n389 B.n388 163.367
R477 B.n390 B.n389 163.367
R478 B.n390 B.n73 163.367
R479 B.n394 B.n73 163.367
R480 B.n395 B.n394 163.367
R481 B.n396 B.n395 163.367
R482 B.n396 B.n71 163.367
R483 B.n400 B.n71 163.367
R484 B.n401 B.n400 163.367
R485 B.n402 B.n401 163.367
R486 B.n402 B.n69 163.367
R487 B.n406 B.n69 163.367
R488 B.n407 B.n406 163.367
R489 B.n408 B.n407 163.367
R490 B.n558 B.n557 163.367
R491 B.n557 B.n556 163.367
R492 B.n556 B.n15 163.367
R493 B.n552 B.n15 163.367
R494 B.n552 B.n551 163.367
R495 B.n551 B.n550 163.367
R496 B.n550 B.n17 163.367
R497 B.n546 B.n17 163.367
R498 B.n546 B.n545 163.367
R499 B.n545 B.n544 163.367
R500 B.n544 B.n19 163.367
R501 B.n540 B.n19 163.367
R502 B.n540 B.n539 163.367
R503 B.n539 B.n538 163.367
R504 B.n538 B.n21 163.367
R505 B.n534 B.n21 163.367
R506 B.n534 B.n533 163.367
R507 B.n533 B.n532 163.367
R508 B.n532 B.n23 163.367
R509 B.n528 B.n23 163.367
R510 B.n528 B.n527 163.367
R511 B.n527 B.n526 163.367
R512 B.n526 B.n25 163.367
R513 B.n522 B.n25 163.367
R514 B.n522 B.n521 163.367
R515 B.n521 B.n520 163.367
R516 B.n520 B.n27 163.367
R517 B.n516 B.n27 163.367
R518 B.n516 B.n515 163.367
R519 B.n515 B.n514 163.367
R520 B.n514 B.n29 163.367
R521 B.n510 B.n29 163.367
R522 B.n510 B.n509 163.367
R523 B.n509 B.n508 163.367
R524 B.n508 B.n31 163.367
R525 B.n504 B.n31 163.367
R526 B.n504 B.n503 163.367
R527 B.n503 B.n502 163.367
R528 B.n502 B.n33 163.367
R529 B.n498 B.n33 163.367
R530 B.n498 B.n497 163.367
R531 B.n497 B.n496 163.367
R532 B.n496 B.n35 163.367
R533 B.n492 B.n35 163.367
R534 B.n492 B.n491 163.367
R535 B.n491 B.n39 163.367
R536 B.n487 B.n39 163.367
R537 B.n487 B.n486 163.367
R538 B.n486 B.n485 163.367
R539 B.n485 B.n41 163.367
R540 B.n481 B.n41 163.367
R541 B.n481 B.n480 163.367
R542 B.n480 B.n479 163.367
R543 B.n479 B.n43 163.367
R544 B.n474 B.n43 163.367
R545 B.n474 B.n473 163.367
R546 B.n473 B.n472 163.367
R547 B.n472 B.n47 163.367
R548 B.n468 B.n47 163.367
R549 B.n468 B.n467 163.367
R550 B.n467 B.n466 163.367
R551 B.n466 B.n49 163.367
R552 B.n462 B.n49 163.367
R553 B.n462 B.n461 163.367
R554 B.n461 B.n460 163.367
R555 B.n460 B.n51 163.367
R556 B.n456 B.n51 163.367
R557 B.n456 B.n455 163.367
R558 B.n455 B.n454 163.367
R559 B.n454 B.n53 163.367
R560 B.n450 B.n53 163.367
R561 B.n450 B.n449 163.367
R562 B.n449 B.n448 163.367
R563 B.n448 B.n55 163.367
R564 B.n444 B.n55 163.367
R565 B.n444 B.n443 163.367
R566 B.n443 B.n442 163.367
R567 B.n442 B.n57 163.367
R568 B.n438 B.n57 163.367
R569 B.n438 B.n437 163.367
R570 B.n437 B.n436 163.367
R571 B.n436 B.n59 163.367
R572 B.n432 B.n59 163.367
R573 B.n432 B.n431 163.367
R574 B.n431 B.n430 163.367
R575 B.n430 B.n61 163.367
R576 B.n426 B.n61 163.367
R577 B.n426 B.n425 163.367
R578 B.n425 B.n424 163.367
R579 B.n424 B.n63 163.367
R580 B.n420 B.n63 163.367
R581 B.n420 B.n419 163.367
R582 B.n419 B.n418 163.367
R583 B.n418 B.n65 163.367
R584 B.n414 B.n65 163.367
R585 B.n414 B.n413 163.367
R586 B.n413 B.n412 163.367
R587 B.n412 B.n67 163.367
R588 B.n114 B.t2 134.034
R589 B.n44 B.t7 134.034
R590 B.n120 B.t11 134.018
R591 B.n36 B.t4 134.018
R592 B.n115 B.t1 109.597
R593 B.n45 B.t8 109.597
R594 B.n121 B.t10 109.582
R595 B.n37 B.t5 109.582
R596 B.n271 B.n115 59.5399
R597 B.n122 B.n121 59.5399
R598 B.n38 B.n37 59.5399
R599 B.n477 B.n45 59.5399
R600 B.n560 B.n559 32.0005
R601 B.n410 B.n409 32.0005
R602 B.n339 B.n338 32.0005
R603 B.n189 B.n188 32.0005
R604 B.n115 B.n114 24.4369
R605 B.n121 B.n120 24.4369
R606 B.n37 B.n36 24.4369
R607 B.n45 B.n44 24.4369
R608 B B.n595 18.0485
R609 B.n559 B.n14 10.6151
R610 B.n555 B.n14 10.6151
R611 B.n555 B.n554 10.6151
R612 B.n554 B.n553 10.6151
R613 B.n553 B.n16 10.6151
R614 B.n549 B.n16 10.6151
R615 B.n549 B.n548 10.6151
R616 B.n548 B.n547 10.6151
R617 B.n547 B.n18 10.6151
R618 B.n543 B.n18 10.6151
R619 B.n543 B.n542 10.6151
R620 B.n542 B.n541 10.6151
R621 B.n541 B.n20 10.6151
R622 B.n537 B.n20 10.6151
R623 B.n537 B.n536 10.6151
R624 B.n536 B.n535 10.6151
R625 B.n535 B.n22 10.6151
R626 B.n531 B.n22 10.6151
R627 B.n531 B.n530 10.6151
R628 B.n530 B.n529 10.6151
R629 B.n529 B.n24 10.6151
R630 B.n525 B.n24 10.6151
R631 B.n525 B.n524 10.6151
R632 B.n524 B.n523 10.6151
R633 B.n523 B.n26 10.6151
R634 B.n519 B.n26 10.6151
R635 B.n519 B.n518 10.6151
R636 B.n518 B.n517 10.6151
R637 B.n517 B.n28 10.6151
R638 B.n513 B.n28 10.6151
R639 B.n513 B.n512 10.6151
R640 B.n512 B.n511 10.6151
R641 B.n511 B.n30 10.6151
R642 B.n507 B.n30 10.6151
R643 B.n507 B.n506 10.6151
R644 B.n506 B.n505 10.6151
R645 B.n505 B.n32 10.6151
R646 B.n501 B.n32 10.6151
R647 B.n501 B.n500 10.6151
R648 B.n500 B.n499 10.6151
R649 B.n499 B.n34 10.6151
R650 B.n495 B.n34 10.6151
R651 B.n495 B.n494 10.6151
R652 B.n494 B.n493 10.6151
R653 B.n490 B.n489 10.6151
R654 B.n489 B.n488 10.6151
R655 B.n488 B.n40 10.6151
R656 B.n484 B.n40 10.6151
R657 B.n484 B.n483 10.6151
R658 B.n483 B.n482 10.6151
R659 B.n482 B.n42 10.6151
R660 B.n478 B.n42 10.6151
R661 B.n476 B.n475 10.6151
R662 B.n475 B.n46 10.6151
R663 B.n471 B.n46 10.6151
R664 B.n471 B.n470 10.6151
R665 B.n470 B.n469 10.6151
R666 B.n469 B.n48 10.6151
R667 B.n465 B.n48 10.6151
R668 B.n465 B.n464 10.6151
R669 B.n464 B.n463 10.6151
R670 B.n463 B.n50 10.6151
R671 B.n459 B.n50 10.6151
R672 B.n459 B.n458 10.6151
R673 B.n458 B.n457 10.6151
R674 B.n457 B.n52 10.6151
R675 B.n453 B.n52 10.6151
R676 B.n453 B.n452 10.6151
R677 B.n452 B.n451 10.6151
R678 B.n451 B.n54 10.6151
R679 B.n447 B.n54 10.6151
R680 B.n447 B.n446 10.6151
R681 B.n446 B.n445 10.6151
R682 B.n445 B.n56 10.6151
R683 B.n441 B.n56 10.6151
R684 B.n441 B.n440 10.6151
R685 B.n440 B.n439 10.6151
R686 B.n439 B.n58 10.6151
R687 B.n435 B.n58 10.6151
R688 B.n435 B.n434 10.6151
R689 B.n434 B.n433 10.6151
R690 B.n433 B.n60 10.6151
R691 B.n429 B.n60 10.6151
R692 B.n429 B.n428 10.6151
R693 B.n428 B.n427 10.6151
R694 B.n427 B.n62 10.6151
R695 B.n423 B.n62 10.6151
R696 B.n423 B.n422 10.6151
R697 B.n422 B.n421 10.6151
R698 B.n421 B.n64 10.6151
R699 B.n417 B.n64 10.6151
R700 B.n417 B.n416 10.6151
R701 B.n416 B.n415 10.6151
R702 B.n415 B.n66 10.6151
R703 B.n411 B.n66 10.6151
R704 B.n411 B.n410 10.6151
R705 B.n339 B.n90 10.6151
R706 B.n343 B.n90 10.6151
R707 B.n344 B.n343 10.6151
R708 B.n345 B.n344 10.6151
R709 B.n345 B.n88 10.6151
R710 B.n349 B.n88 10.6151
R711 B.n350 B.n349 10.6151
R712 B.n351 B.n350 10.6151
R713 B.n351 B.n86 10.6151
R714 B.n355 B.n86 10.6151
R715 B.n356 B.n355 10.6151
R716 B.n357 B.n356 10.6151
R717 B.n357 B.n84 10.6151
R718 B.n361 B.n84 10.6151
R719 B.n362 B.n361 10.6151
R720 B.n363 B.n362 10.6151
R721 B.n363 B.n82 10.6151
R722 B.n367 B.n82 10.6151
R723 B.n368 B.n367 10.6151
R724 B.n369 B.n368 10.6151
R725 B.n369 B.n80 10.6151
R726 B.n373 B.n80 10.6151
R727 B.n374 B.n373 10.6151
R728 B.n375 B.n374 10.6151
R729 B.n375 B.n78 10.6151
R730 B.n379 B.n78 10.6151
R731 B.n380 B.n379 10.6151
R732 B.n381 B.n380 10.6151
R733 B.n381 B.n76 10.6151
R734 B.n385 B.n76 10.6151
R735 B.n386 B.n385 10.6151
R736 B.n387 B.n386 10.6151
R737 B.n387 B.n74 10.6151
R738 B.n391 B.n74 10.6151
R739 B.n392 B.n391 10.6151
R740 B.n393 B.n392 10.6151
R741 B.n393 B.n72 10.6151
R742 B.n397 B.n72 10.6151
R743 B.n398 B.n397 10.6151
R744 B.n399 B.n398 10.6151
R745 B.n399 B.n70 10.6151
R746 B.n403 B.n70 10.6151
R747 B.n404 B.n403 10.6151
R748 B.n405 B.n404 10.6151
R749 B.n405 B.n68 10.6151
R750 B.n409 B.n68 10.6151
R751 B.n189 B.n144 10.6151
R752 B.n193 B.n144 10.6151
R753 B.n194 B.n193 10.6151
R754 B.n195 B.n194 10.6151
R755 B.n195 B.n142 10.6151
R756 B.n199 B.n142 10.6151
R757 B.n200 B.n199 10.6151
R758 B.n201 B.n200 10.6151
R759 B.n201 B.n140 10.6151
R760 B.n205 B.n140 10.6151
R761 B.n206 B.n205 10.6151
R762 B.n207 B.n206 10.6151
R763 B.n207 B.n138 10.6151
R764 B.n211 B.n138 10.6151
R765 B.n212 B.n211 10.6151
R766 B.n213 B.n212 10.6151
R767 B.n213 B.n136 10.6151
R768 B.n217 B.n136 10.6151
R769 B.n218 B.n217 10.6151
R770 B.n219 B.n218 10.6151
R771 B.n219 B.n134 10.6151
R772 B.n223 B.n134 10.6151
R773 B.n224 B.n223 10.6151
R774 B.n225 B.n224 10.6151
R775 B.n225 B.n132 10.6151
R776 B.n229 B.n132 10.6151
R777 B.n230 B.n229 10.6151
R778 B.n231 B.n230 10.6151
R779 B.n231 B.n130 10.6151
R780 B.n235 B.n130 10.6151
R781 B.n236 B.n235 10.6151
R782 B.n237 B.n236 10.6151
R783 B.n237 B.n128 10.6151
R784 B.n241 B.n128 10.6151
R785 B.n242 B.n241 10.6151
R786 B.n243 B.n242 10.6151
R787 B.n243 B.n126 10.6151
R788 B.n247 B.n126 10.6151
R789 B.n248 B.n247 10.6151
R790 B.n249 B.n248 10.6151
R791 B.n249 B.n124 10.6151
R792 B.n253 B.n124 10.6151
R793 B.n254 B.n253 10.6151
R794 B.n255 B.n254 10.6151
R795 B.n259 B.n258 10.6151
R796 B.n260 B.n259 10.6151
R797 B.n260 B.n118 10.6151
R798 B.n264 B.n118 10.6151
R799 B.n265 B.n264 10.6151
R800 B.n266 B.n265 10.6151
R801 B.n266 B.n116 10.6151
R802 B.n270 B.n116 10.6151
R803 B.n273 B.n272 10.6151
R804 B.n273 B.n112 10.6151
R805 B.n277 B.n112 10.6151
R806 B.n278 B.n277 10.6151
R807 B.n279 B.n278 10.6151
R808 B.n279 B.n110 10.6151
R809 B.n283 B.n110 10.6151
R810 B.n284 B.n283 10.6151
R811 B.n285 B.n284 10.6151
R812 B.n285 B.n108 10.6151
R813 B.n289 B.n108 10.6151
R814 B.n290 B.n289 10.6151
R815 B.n291 B.n290 10.6151
R816 B.n291 B.n106 10.6151
R817 B.n295 B.n106 10.6151
R818 B.n296 B.n295 10.6151
R819 B.n297 B.n296 10.6151
R820 B.n297 B.n104 10.6151
R821 B.n301 B.n104 10.6151
R822 B.n302 B.n301 10.6151
R823 B.n303 B.n302 10.6151
R824 B.n303 B.n102 10.6151
R825 B.n307 B.n102 10.6151
R826 B.n308 B.n307 10.6151
R827 B.n309 B.n308 10.6151
R828 B.n309 B.n100 10.6151
R829 B.n313 B.n100 10.6151
R830 B.n314 B.n313 10.6151
R831 B.n315 B.n314 10.6151
R832 B.n315 B.n98 10.6151
R833 B.n319 B.n98 10.6151
R834 B.n320 B.n319 10.6151
R835 B.n321 B.n320 10.6151
R836 B.n321 B.n96 10.6151
R837 B.n325 B.n96 10.6151
R838 B.n326 B.n325 10.6151
R839 B.n327 B.n326 10.6151
R840 B.n327 B.n94 10.6151
R841 B.n331 B.n94 10.6151
R842 B.n332 B.n331 10.6151
R843 B.n333 B.n332 10.6151
R844 B.n333 B.n92 10.6151
R845 B.n337 B.n92 10.6151
R846 B.n338 B.n337 10.6151
R847 B.n188 B.n187 10.6151
R848 B.n187 B.n146 10.6151
R849 B.n183 B.n146 10.6151
R850 B.n183 B.n182 10.6151
R851 B.n182 B.n181 10.6151
R852 B.n181 B.n148 10.6151
R853 B.n177 B.n148 10.6151
R854 B.n177 B.n176 10.6151
R855 B.n176 B.n175 10.6151
R856 B.n175 B.n150 10.6151
R857 B.n171 B.n150 10.6151
R858 B.n171 B.n170 10.6151
R859 B.n170 B.n169 10.6151
R860 B.n169 B.n152 10.6151
R861 B.n165 B.n152 10.6151
R862 B.n165 B.n164 10.6151
R863 B.n164 B.n163 10.6151
R864 B.n163 B.n154 10.6151
R865 B.n159 B.n154 10.6151
R866 B.n159 B.n158 10.6151
R867 B.n158 B.n157 10.6151
R868 B.n157 B.n0 10.6151
R869 B.n591 B.n1 10.6151
R870 B.n591 B.n590 10.6151
R871 B.n590 B.n589 10.6151
R872 B.n589 B.n4 10.6151
R873 B.n585 B.n4 10.6151
R874 B.n585 B.n584 10.6151
R875 B.n584 B.n583 10.6151
R876 B.n583 B.n6 10.6151
R877 B.n579 B.n6 10.6151
R878 B.n579 B.n578 10.6151
R879 B.n578 B.n577 10.6151
R880 B.n577 B.n8 10.6151
R881 B.n573 B.n8 10.6151
R882 B.n573 B.n572 10.6151
R883 B.n572 B.n571 10.6151
R884 B.n571 B.n10 10.6151
R885 B.n567 B.n10 10.6151
R886 B.n567 B.n566 10.6151
R887 B.n566 B.n565 10.6151
R888 B.n565 B.n12 10.6151
R889 B.n561 B.n12 10.6151
R890 B.n561 B.n560 10.6151
R891 B.n490 B.n38 6.5566
R892 B.n478 B.n477 6.5566
R893 B.n258 B.n122 6.5566
R894 B.n271 B.n270 6.5566
R895 B.n493 B.n38 4.05904
R896 B.n477 B.n476 4.05904
R897 B.n255 B.n122 4.05904
R898 B.n272 B.n271 4.05904
R899 B.n595 B.n0 2.81026
R900 B.n595 B.n1 2.81026
R901 VN.n2 VN.t1 399.238
R902 VN.n10 VN.t3 399.238
R903 VN.n6 VN.t2 381.195
R904 VN.n14 VN.t4 381.195
R905 VN.n1 VN.t0 338.438
R906 VN.n9 VN.t5 338.438
R907 VN.n7 VN.n6 161.3
R908 VN.n15 VN.n14 161.3
R909 VN.n13 VN.n8 161.3
R910 VN.n12 VN.n11 161.3
R911 VN.n5 VN.n0 161.3
R912 VN.n4 VN.n3 161.3
R913 VN.n5 VN.n4 52.0954
R914 VN.n13 VN.n12 52.0954
R915 VN.n11 VN.n10 43.4068
R916 VN.n3 VN.n2 43.4068
R917 VN VN.n15 43.3282
R918 VN.n2 VN.n1 42.3264
R919 VN.n10 VN.n9 42.3264
R920 VN.n4 VN.n1 12.1722
R921 VN.n12 VN.n9 12.1722
R922 VN.n6 VN.n5 6.57323
R923 VN.n14 VN.n13 6.57323
R924 VN.n15 VN.n8 0.189894
R925 VN.n11 VN.n8 0.189894
R926 VN.n3 VN.n0 0.189894
R927 VN.n7 VN.n0 0.189894
R928 VN VN.n7 0.0516364
R929 VDD2.n1 VDD2.t3 79.8235
R930 VDD2.n2 VDD2.t4 79.0653
R931 VDD2.n1 VDD2.n0 76.7915
R932 VDD2 VDD2.n3 76.7887
R933 VDD2.n2 VDD2.n1 38.5041
R934 VDD2.n3 VDD2.t1 2.4894
R935 VDD2.n3 VDD2.t5 2.4894
R936 VDD2.n0 VDD2.t0 2.4894
R937 VDD2.n0 VDD2.t2 2.4894
R938 VDD2 VDD2.n2 0.873345
R939 VTAIL.n7 VTAIL.t8 62.3865
R940 VTAIL.n11 VTAIL.t9 62.3854
R941 VTAIL.n2 VTAIL.t0 62.3854
R942 VTAIL.n10 VTAIL.t1 62.3854
R943 VTAIL.n9 VTAIL.n8 59.8977
R944 VTAIL.n6 VTAIL.n5 59.8977
R945 VTAIL.n1 VTAIL.n0 59.8965
R946 VTAIL.n4 VTAIL.n3 59.8965
R947 VTAIL.n6 VTAIL.n4 25.7979
R948 VTAIL.n11 VTAIL.n10 24.7117
R949 VTAIL.n0 VTAIL.t10 2.4894
R950 VTAIL.n0 VTAIL.t11 2.4894
R951 VTAIL.n3 VTAIL.t2 2.4894
R952 VTAIL.n3 VTAIL.t5 2.4894
R953 VTAIL.n8 VTAIL.t4 2.4894
R954 VTAIL.n8 VTAIL.t3 2.4894
R955 VTAIL.n5 VTAIL.t7 2.4894
R956 VTAIL.n5 VTAIL.t6 2.4894
R957 VTAIL.n7 VTAIL.n6 1.08671
R958 VTAIL.n10 VTAIL.n9 1.08671
R959 VTAIL.n4 VTAIL.n2 1.08671
R960 VTAIL.n9 VTAIL.n7 1.01343
R961 VTAIL.n2 VTAIL.n1 1.01343
R962 VTAIL VTAIL.n11 0.756965
R963 VTAIL VTAIL.n1 0.330241
R964 VP.n5 VP.t2 399.238
R965 VP.n12 VP.t4 381.195
R966 VP.n19 VP.t0 381.195
R967 VP.n9 VP.t3 381.195
R968 VP.n1 VP.t1 338.438
R969 VP.n4 VP.t5 338.438
R970 VP.n20 VP.n19 161.3
R971 VP.n7 VP.n6 161.3
R972 VP.n8 VP.n3 161.3
R973 VP.n10 VP.n9 161.3
R974 VP.n18 VP.n0 161.3
R975 VP.n17 VP.n16 161.3
R976 VP.n15 VP.n14 161.3
R977 VP.n13 VP.n2 161.3
R978 VP.n12 VP.n11 161.3
R979 VP.n14 VP.n13 52.0954
R980 VP.n18 VP.n17 52.0954
R981 VP.n8 VP.n7 52.0954
R982 VP.n6 VP.n5 43.4068
R983 VP.n11 VP.n10 42.9475
R984 VP.n5 VP.n4 42.3264
R985 VP.n14 VP.n1 12.1722
R986 VP.n17 VP.n1 12.1722
R987 VP.n7 VP.n4 12.1722
R988 VP.n13 VP.n12 6.57323
R989 VP.n19 VP.n18 6.57323
R990 VP.n9 VP.n8 6.57323
R991 VP.n6 VP.n3 0.189894
R992 VP.n10 VP.n3 0.189894
R993 VP.n11 VP.n2 0.189894
R994 VP.n15 VP.n2 0.189894
R995 VP.n16 VP.n15 0.189894
R996 VP.n16 VP.n0 0.189894
R997 VP.n20 VP.n0 0.189894
R998 VP VP.n20 0.0516364
R999 VDD1 VDD1.t3 79.9382
R1000 VDD1.n1 VDD1.t1 79.8235
R1001 VDD1.n1 VDD1.n0 76.7915
R1002 VDD1.n3 VDD1.n2 76.5753
R1003 VDD1.n3 VDD1.n1 39.6302
R1004 VDD1.n2 VDD1.t0 2.4894
R1005 VDD1.n2 VDD1.t2 2.4894
R1006 VDD1.n0 VDD1.t4 2.4894
R1007 VDD1.n0 VDD1.t5 2.4894
R1008 VDD1 VDD1.n3 0.213862
C0 VDD1 w_n1978_n3580# 1.95015f
C1 VN w_n1978_n3580# 3.36287f
C2 VTAIL B 3.05433f
C3 VP VDD2 0.316813f
C4 VP w_n1978_n3580# 3.61395f
C5 w_n1978_n3580# VDD2 1.98161f
C6 VDD1 B 1.70786f
C7 VN B 0.823507f
C8 VTAIL VDD1 9.62012f
C9 VN VTAIL 5.04938f
C10 VP B 1.23429f
C11 B VDD2 1.74223f
C12 VP VTAIL 5.06395f
C13 VTAIL VDD2 9.65604f
C14 w_n1978_n3580# B 7.66765f
C15 VTAIL w_n1978_n3580# 3.09547f
C16 VN VDD1 0.148094f
C17 VP VDD1 5.50889f
C18 VDD1 VDD2 0.794682f
C19 VN VP 5.50189f
C20 VN VDD2 5.34474f
C21 VDD2 VSUBS 1.359157f
C22 VDD1 VSUBS 1.678833f
C23 VTAIL VSUBS 0.856328f
C24 VN VSUBS 4.59482f
C25 VP VSUBS 1.683699f
C26 B VSUBS 3.06921f
C27 w_n1978_n3580# VSUBS 87.0399f
C28 VDD1.t3 VSUBS 2.43378f
C29 VDD1.t1 VSUBS 2.43292f
C30 VDD1.t4 VSUBS 0.232792f
C31 VDD1.t5 VSUBS 0.232792f
C32 VDD1.n0 VSUBS 1.86564f
C33 VDD1.n1 VSUBS 2.55885f
C34 VDD1.t0 VSUBS 0.232792f
C35 VDD1.t2 VSUBS 0.232792f
C36 VDD1.n2 VSUBS 1.86419f
C37 VDD1.n3 VSUBS 2.38843f
C38 VP.n0 VSUBS 0.050945f
C39 VP.t1 VSUBS 1.68981f
C40 VP.n1 VSUBS 0.625138f
C41 VP.n2 VSUBS 0.050945f
C42 VP.n3 VSUBS 0.050945f
C43 VP.t3 VSUBS 1.76284f
C44 VP.t5 VSUBS 1.68981f
C45 VP.n4 VSUBS 0.674557f
C46 VP.t2 VSUBS 1.79432f
C47 VP.n5 VSUBS 0.688828f
C48 VP.n6 VSUBS 0.216833f
C49 VP.n7 VSUBS 0.068353f
C50 VP.n8 VSUBS 0.01743f
C51 VP.n9 VSUBS 0.68287f
C52 VP.n10 VSUBS 2.18195f
C53 VP.n11 VSUBS 2.22447f
C54 VP.t4 VSUBS 1.76284f
C55 VP.n12 VSUBS 0.68287f
C56 VP.n13 VSUBS 0.01743f
C57 VP.n14 VSUBS 0.068353f
C58 VP.n15 VSUBS 0.050945f
C59 VP.n16 VSUBS 0.050945f
C60 VP.n17 VSUBS 0.068353f
C61 VP.n18 VSUBS 0.01743f
C62 VP.t0 VSUBS 1.76284f
C63 VP.n19 VSUBS 0.68287f
C64 VP.n20 VSUBS 0.03948f
C65 VTAIL.t10 VSUBS 0.293518f
C66 VTAIL.t11 VSUBS 0.293518f
C67 VTAIL.n0 VSUBS 2.20866f
C68 VTAIL.n1 VSUBS 0.740963f
C69 VTAIL.t0 VSUBS 2.90081f
C70 VTAIL.n2 VSUBS 0.918631f
C71 VTAIL.t2 VSUBS 0.293518f
C72 VTAIL.t5 VSUBS 0.293518f
C73 VTAIL.n3 VSUBS 2.20866f
C74 VTAIL.n4 VSUBS 2.33463f
C75 VTAIL.t7 VSUBS 0.293518f
C76 VTAIL.t6 VSUBS 0.293518f
C77 VTAIL.n5 VSUBS 2.20868f
C78 VTAIL.n6 VSUBS 2.33461f
C79 VTAIL.t8 VSUBS 2.90084f
C80 VTAIL.n7 VSUBS 0.918608f
C81 VTAIL.t4 VSUBS 0.293518f
C82 VTAIL.t3 VSUBS 0.293518f
C83 VTAIL.n8 VSUBS 2.20868f
C84 VTAIL.n9 VSUBS 0.810268f
C85 VTAIL.t1 VSUBS 2.90081f
C86 VTAIL.n10 VSUBS 2.34344f
C87 VTAIL.t9 VSUBS 2.90081f
C88 VTAIL.n11 VSUBS 2.31322f
C89 VDD2.t3 VSUBS 2.43021f
C90 VDD2.t0 VSUBS 0.232533f
C91 VDD2.t2 VSUBS 0.232533f
C92 VDD2.n0 VSUBS 1.86357f
C93 VDD2.n1 VSUBS 2.48128f
C94 VDD2.t4 VSUBS 2.42505f
C95 VDD2.n2 VSUBS 2.41755f
C96 VDD2.t1 VSUBS 0.232533f
C97 VDD2.t5 VSUBS 0.232533f
C98 VDD2.n3 VSUBS 1.86354f
C99 VN.n0 VSUBS 0.049472f
C100 VN.t0 VSUBS 1.64096f
C101 VN.n1 VSUBS 0.655055f
C102 VN.t1 VSUBS 1.74245f
C103 VN.n2 VSUBS 0.668914f
C104 VN.n3 VSUBS 0.210564f
C105 VN.n4 VSUBS 0.066377f
C106 VN.n5 VSUBS 0.016926f
C107 VN.t2 VSUBS 1.71187f
C108 VN.n6 VSUBS 0.663128f
C109 VN.n7 VSUBS 0.038339f
C110 VN.n8 VSUBS 0.049472f
C111 VN.t5 VSUBS 1.64096f
C112 VN.n9 VSUBS 0.655055f
C113 VN.t3 VSUBS 1.74245f
C114 VN.n10 VSUBS 0.668914f
C115 VN.n11 VSUBS 0.210564f
C116 VN.n12 VSUBS 0.066377f
C117 VN.n13 VSUBS 0.016926f
C118 VN.t4 VSUBS 1.71187f
C119 VN.n14 VSUBS 0.663128f
C120 VN.n15 VSUBS 2.1513f
C121 B.n0 VSUBS 0.004461f
C122 B.n1 VSUBS 0.004461f
C123 B.n2 VSUBS 0.007055f
C124 B.n3 VSUBS 0.007055f
C125 B.n4 VSUBS 0.007055f
C126 B.n5 VSUBS 0.007055f
C127 B.n6 VSUBS 0.007055f
C128 B.n7 VSUBS 0.007055f
C129 B.n8 VSUBS 0.007055f
C130 B.n9 VSUBS 0.007055f
C131 B.n10 VSUBS 0.007055f
C132 B.n11 VSUBS 0.007055f
C133 B.n12 VSUBS 0.007055f
C134 B.n13 VSUBS 0.015947f
C135 B.n14 VSUBS 0.007055f
C136 B.n15 VSUBS 0.007055f
C137 B.n16 VSUBS 0.007055f
C138 B.n17 VSUBS 0.007055f
C139 B.n18 VSUBS 0.007055f
C140 B.n19 VSUBS 0.007055f
C141 B.n20 VSUBS 0.007055f
C142 B.n21 VSUBS 0.007055f
C143 B.n22 VSUBS 0.007055f
C144 B.n23 VSUBS 0.007055f
C145 B.n24 VSUBS 0.007055f
C146 B.n25 VSUBS 0.007055f
C147 B.n26 VSUBS 0.007055f
C148 B.n27 VSUBS 0.007055f
C149 B.n28 VSUBS 0.007055f
C150 B.n29 VSUBS 0.007055f
C151 B.n30 VSUBS 0.007055f
C152 B.n31 VSUBS 0.007055f
C153 B.n32 VSUBS 0.007055f
C154 B.n33 VSUBS 0.007055f
C155 B.n34 VSUBS 0.007055f
C156 B.n35 VSUBS 0.007055f
C157 B.t5 VSUBS 0.432705f
C158 B.t4 VSUBS 0.442806f
C159 B.t3 VSUBS 0.512691f
C160 B.n36 VSUBS 0.163355f
C161 B.n37 VSUBS 0.065459f
C162 B.n38 VSUBS 0.016346f
C163 B.n39 VSUBS 0.007055f
C164 B.n40 VSUBS 0.007055f
C165 B.n41 VSUBS 0.007055f
C166 B.n42 VSUBS 0.007055f
C167 B.n43 VSUBS 0.007055f
C168 B.t8 VSUBS 0.432696f
C169 B.t7 VSUBS 0.442797f
C170 B.t6 VSUBS 0.512691f
C171 B.n44 VSUBS 0.163364f
C172 B.n45 VSUBS 0.065469f
C173 B.n46 VSUBS 0.007055f
C174 B.n47 VSUBS 0.007055f
C175 B.n48 VSUBS 0.007055f
C176 B.n49 VSUBS 0.007055f
C177 B.n50 VSUBS 0.007055f
C178 B.n51 VSUBS 0.007055f
C179 B.n52 VSUBS 0.007055f
C180 B.n53 VSUBS 0.007055f
C181 B.n54 VSUBS 0.007055f
C182 B.n55 VSUBS 0.007055f
C183 B.n56 VSUBS 0.007055f
C184 B.n57 VSUBS 0.007055f
C185 B.n58 VSUBS 0.007055f
C186 B.n59 VSUBS 0.007055f
C187 B.n60 VSUBS 0.007055f
C188 B.n61 VSUBS 0.007055f
C189 B.n62 VSUBS 0.007055f
C190 B.n63 VSUBS 0.007055f
C191 B.n64 VSUBS 0.007055f
C192 B.n65 VSUBS 0.007055f
C193 B.n66 VSUBS 0.007055f
C194 B.n67 VSUBS 0.016632f
C195 B.n68 VSUBS 0.007055f
C196 B.n69 VSUBS 0.007055f
C197 B.n70 VSUBS 0.007055f
C198 B.n71 VSUBS 0.007055f
C199 B.n72 VSUBS 0.007055f
C200 B.n73 VSUBS 0.007055f
C201 B.n74 VSUBS 0.007055f
C202 B.n75 VSUBS 0.007055f
C203 B.n76 VSUBS 0.007055f
C204 B.n77 VSUBS 0.007055f
C205 B.n78 VSUBS 0.007055f
C206 B.n79 VSUBS 0.007055f
C207 B.n80 VSUBS 0.007055f
C208 B.n81 VSUBS 0.007055f
C209 B.n82 VSUBS 0.007055f
C210 B.n83 VSUBS 0.007055f
C211 B.n84 VSUBS 0.007055f
C212 B.n85 VSUBS 0.007055f
C213 B.n86 VSUBS 0.007055f
C214 B.n87 VSUBS 0.007055f
C215 B.n88 VSUBS 0.007055f
C216 B.n89 VSUBS 0.007055f
C217 B.n90 VSUBS 0.007055f
C218 B.n91 VSUBS 0.016632f
C219 B.n92 VSUBS 0.007055f
C220 B.n93 VSUBS 0.007055f
C221 B.n94 VSUBS 0.007055f
C222 B.n95 VSUBS 0.007055f
C223 B.n96 VSUBS 0.007055f
C224 B.n97 VSUBS 0.007055f
C225 B.n98 VSUBS 0.007055f
C226 B.n99 VSUBS 0.007055f
C227 B.n100 VSUBS 0.007055f
C228 B.n101 VSUBS 0.007055f
C229 B.n102 VSUBS 0.007055f
C230 B.n103 VSUBS 0.007055f
C231 B.n104 VSUBS 0.007055f
C232 B.n105 VSUBS 0.007055f
C233 B.n106 VSUBS 0.007055f
C234 B.n107 VSUBS 0.007055f
C235 B.n108 VSUBS 0.007055f
C236 B.n109 VSUBS 0.007055f
C237 B.n110 VSUBS 0.007055f
C238 B.n111 VSUBS 0.007055f
C239 B.n112 VSUBS 0.007055f
C240 B.n113 VSUBS 0.007055f
C241 B.t1 VSUBS 0.432696f
C242 B.t2 VSUBS 0.442797f
C243 B.t0 VSUBS 0.512691f
C244 B.n114 VSUBS 0.163364f
C245 B.n115 VSUBS 0.065469f
C246 B.n116 VSUBS 0.007055f
C247 B.n117 VSUBS 0.007055f
C248 B.n118 VSUBS 0.007055f
C249 B.n119 VSUBS 0.007055f
C250 B.t10 VSUBS 0.432705f
C251 B.t11 VSUBS 0.442806f
C252 B.t9 VSUBS 0.512691f
C253 B.n120 VSUBS 0.163355f
C254 B.n121 VSUBS 0.065459f
C255 B.n122 VSUBS 0.016346f
C256 B.n123 VSUBS 0.007055f
C257 B.n124 VSUBS 0.007055f
C258 B.n125 VSUBS 0.007055f
C259 B.n126 VSUBS 0.007055f
C260 B.n127 VSUBS 0.007055f
C261 B.n128 VSUBS 0.007055f
C262 B.n129 VSUBS 0.007055f
C263 B.n130 VSUBS 0.007055f
C264 B.n131 VSUBS 0.007055f
C265 B.n132 VSUBS 0.007055f
C266 B.n133 VSUBS 0.007055f
C267 B.n134 VSUBS 0.007055f
C268 B.n135 VSUBS 0.007055f
C269 B.n136 VSUBS 0.007055f
C270 B.n137 VSUBS 0.007055f
C271 B.n138 VSUBS 0.007055f
C272 B.n139 VSUBS 0.007055f
C273 B.n140 VSUBS 0.007055f
C274 B.n141 VSUBS 0.007055f
C275 B.n142 VSUBS 0.007055f
C276 B.n143 VSUBS 0.007055f
C277 B.n144 VSUBS 0.007055f
C278 B.n145 VSUBS 0.015947f
C279 B.n146 VSUBS 0.007055f
C280 B.n147 VSUBS 0.007055f
C281 B.n148 VSUBS 0.007055f
C282 B.n149 VSUBS 0.007055f
C283 B.n150 VSUBS 0.007055f
C284 B.n151 VSUBS 0.007055f
C285 B.n152 VSUBS 0.007055f
C286 B.n153 VSUBS 0.007055f
C287 B.n154 VSUBS 0.007055f
C288 B.n155 VSUBS 0.007055f
C289 B.n156 VSUBS 0.007055f
C290 B.n157 VSUBS 0.007055f
C291 B.n158 VSUBS 0.007055f
C292 B.n159 VSUBS 0.007055f
C293 B.n160 VSUBS 0.007055f
C294 B.n161 VSUBS 0.007055f
C295 B.n162 VSUBS 0.007055f
C296 B.n163 VSUBS 0.007055f
C297 B.n164 VSUBS 0.007055f
C298 B.n165 VSUBS 0.007055f
C299 B.n166 VSUBS 0.007055f
C300 B.n167 VSUBS 0.007055f
C301 B.n168 VSUBS 0.007055f
C302 B.n169 VSUBS 0.007055f
C303 B.n170 VSUBS 0.007055f
C304 B.n171 VSUBS 0.007055f
C305 B.n172 VSUBS 0.007055f
C306 B.n173 VSUBS 0.007055f
C307 B.n174 VSUBS 0.007055f
C308 B.n175 VSUBS 0.007055f
C309 B.n176 VSUBS 0.007055f
C310 B.n177 VSUBS 0.007055f
C311 B.n178 VSUBS 0.007055f
C312 B.n179 VSUBS 0.007055f
C313 B.n180 VSUBS 0.007055f
C314 B.n181 VSUBS 0.007055f
C315 B.n182 VSUBS 0.007055f
C316 B.n183 VSUBS 0.007055f
C317 B.n184 VSUBS 0.007055f
C318 B.n185 VSUBS 0.007055f
C319 B.n186 VSUBS 0.007055f
C320 B.n187 VSUBS 0.007055f
C321 B.n188 VSUBS 0.015947f
C322 B.n189 VSUBS 0.016632f
C323 B.n190 VSUBS 0.016632f
C324 B.n191 VSUBS 0.007055f
C325 B.n192 VSUBS 0.007055f
C326 B.n193 VSUBS 0.007055f
C327 B.n194 VSUBS 0.007055f
C328 B.n195 VSUBS 0.007055f
C329 B.n196 VSUBS 0.007055f
C330 B.n197 VSUBS 0.007055f
C331 B.n198 VSUBS 0.007055f
C332 B.n199 VSUBS 0.007055f
C333 B.n200 VSUBS 0.007055f
C334 B.n201 VSUBS 0.007055f
C335 B.n202 VSUBS 0.007055f
C336 B.n203 VSUBS 0.007055f
C337 B.n204 VSUBS 0.007055f
C338 B.n205 VSUBS 0.007055f
C339 B.n206 VSUBS 0.007055f
C340 B.n207 VSUBS 0.007055f
C341 B.n208 VSUBS 0.007055f
C342 B.n209 VSUBS 0.007055f
C343 B.n210 VSUBS 0.007055f
C344 B.n211 VSUBS 0.007055f
C345 B.n212 VSUBS 0.007055f
C346 B.n213 VSUBS 0.007055f
C347 B.n214 VSUBS 0.007055f
C348 B.n215 VSUBS 0.007055f
C349 B.n216 VSUBS 0.007055f
C350 B.n217 VSUBS 0.007055f
C351 B.n218 VSUBS 0.007055f
C352 B.n219 VSUBS 0.007055f
C353 B.n220 VSUBS 0.007055f
C354 B.n221 VSUBS 0.007055f
C355 B.n222 VSUBS 0.007055f
C356 B.n223 VSUBS 0.007055f
C357 B.n224 VSUBS 0.007055f
C358 B.n225 VSUBS 0.007055f
C359 B.n226 VSUBS 0.007055f
C360 B.n227 VSUBS 0.007055f
C361 B.n228 VSUBS 0.007055f
C362 B.n229 VSUBS 0.007055f
C363 B.n230 VSUBS 0.007055f
C364 B.n231 VSUBS 0.007055f
C365 B.n232 VSUBS 0.007055f
C366 B.n233 VSUBS 0.007055f
C367 B.n234 VSUBS 0.007055f
C368 B.n235 VSUBS 0.007055f
C369 B.n236 VSUBS 0.007055f
C370 B.n237 VSUBS 0.007055f
C371 B.n238 VSUBS 0.007055f
C372 B.n239 VSUBS 0.007055f
C373 B.n240 VSUBS 0.007055f
C374 B.n241 VSUBS 0.007055f
C375 B.n242 VSUBS 0.007055f
C376 B.n243 VSUBS 0.007055f
C377 B.n244 VSUBS 0.007055f
C378 B.n245 VSUBS 0.007055f
C379 B.n246 VSUBS 0.007055f
C380 B.n247 VSUBS 0.007055f
C381 B.n248 VSUBS 0.007055f
C382 B.n249 VSUBS 0.007055f
C383 B.n250 VSUBS 0.007055f
C384 B.n251 VSUBS 0.007055f
C385 B.n252 VSUBS 0.007055f
C386 B.n253 VSUBS 0.007055f
C387 B.n254 VSUBS 0.007055f
C388 B.n255 VSUBS 0.004876f
C389 B.n256 VSUBS 0.007055f
C390 B.n257 VSUBS 0.007055f
C391 B.n258 VSUBS 0.005706f
C392 B.n259 VSUBS 0.007055f
C393 B.n260 VSUBS 0.007055f
C394 B.n261 VSUBS 0.007055f
C395 B.n262 VSUBS 0.007055f
C396 B.n263 VSUBS 0.007055f
C397 B.n264 VSUBS 0.007055f
C398 B.n265 VSUBS 0.007055f
C399 B.n266 VSUBS 0.007055f
C400 B.n267 VSUBS 0.007055f
C401 B.n268 VSUBS 0.007055f
C402 B.n269 VSUBS 0.007055f
C403 B.n270 VSUBS 0.005706f
C404 B.n271 VSUBS 0.016346f
C405 B.n272 VSUBS 0.004876f
C406 B.n273 VSUBS 0.007055f
C407 B.n274 VSUBS 0.007055f
C408 B.n275 VSUBS 0.007055f
C409 B.n276 VSUBS 0.007055f
C410 B.n277 VSUBS 0.007055f
C411 B.n278 VSUBS 0.007055f
C412 B.n279 VSUBS 0.007055f
C413 B.n280 VSUBS 0.007055f
C414 B.n281 VSUBS 0.007055f
C415 B.n282 VSUBS 0.007055f
C416 B.n283 VSUBS 0.007055f
C417 B.n284 VSUBS 0.007055f
C418 B.n285 VSUBS 0.007055f
C419 B.n286 VSUBS 0.007055f
C420 B.n287 VSUBS 0.007055f
C421 B.n288 VSUBS 0.007055f
C422 B.n289 VSUBS 0.007055f
C423 B.n290 VSUBS 0.007055f
C424 B.n291 VSUBS 0.007055f
C425 B.n292 VSUBS 0.007055f
C426 B.n293 VSUBS 0.007055f
C427 B.n294 VSUBS 0.007055f
C428 B.n295 VSUBS 0.007055f
C429 B.n296 VSUBS 0.007055f
C430 B.n297 VSUBS 0.007055f
C431 B.n298 VSUBS 0.007055f
C432 B.n299 VSUBS 0.007055f
C433 B.n300 VSUBS 0.007055f
C434 B.n301 VSUBS 0.007055f
C435 B.n302 VSUBS 0.007055f
C436 B.n303 VSUBS 0.007055f
C437 B.n304 VSUBS 0.007055f
C438 B.n305 VSUBS 0.007055f
C439 B.n306 VSUBS 0.007055f
C440 B.n307 VSUBS 0.007055f
C441 B.n308 VSUBS 0.007055f
C442 B.n309 VSUBS 0.007055f
C443 B.n310 VSUBS 0.007055f
C444 B.n311 VSUBS 0.007055f
C445 B.n312 VSUBS 0.007055f
C446 B.n313 VSUBS 0.007055f
C447 B.n314 VSUBS 0.007055f
C448 B.n315 VSUBS 0.007055f
C449 B.n316 VSUBS 0.007055f
C450 B.n317 VSUBS 0.007055f
C451 B.n318 VSUBS 0.007055f
C452 B.n319 VSUBS 0.007055f
C453 B.n320 VSUBS 0.007055f
C454 B.n321 VSUBS 0.007055f
C455 B.n322 VSUBS 0.007055f
C456 B.n323 VSUBS 0.007055f
C457 B.n324 VSUBS 0.007055f
C458 B.n325 VSUBS 0.007055f
C459 B.n326 VSUBS 0.007055f
C460 B.n327 VSUBS 0.007055f
C461 B.n328 VSUBS 0.007055f
C462 B.n329 VSUBS 0.007055f
C463 B.n330 VSUBS 0.007055f
C464 B.n331 VSUBS 0.007055f
C465 B.n332 VSUBS 0.007055f
C466 B.n333 VSUBS 0.007055f
C467 B.n334 VSUBS 0.007055f
C468 B.n335 VSUBS 0.007055f
C469 B.n336 VSUBS 0.007055f
C470 B.n337 VSUBS 0.007055f
C471 B.n338 VSUBS 0.016632f
C472 B.n339 VSUBS 0.015947f
C473 B.n340 VSUBS 0.015947f
C474 B.n341 VSUBS 0.007055f
C475 B.n342 VSUBS 0.007055f
C476 B.n343 VSUBS 0.007055f
C477 B.n344 VSUBS 0.007055f
C478 B.n345 VSUBS 0.007055f
C479 B.n346 VSUBS 0.007055f
C480 B.n347 VSUBS 0.007055f
C481 B.n348 VSUBS 0.007055f
C482 B.n349 VSUBS 0.007055f
C483 B.n350 VSUBS 0.007055f
C484 B.n351 VSUBS 0.007055f
C485 B.n352 VSUBS 0.007055f
C486 B.n353 VSUBS 0.007055f
C487 B.n354 VSUBS 0.007055f
C488 B.n355 VSUBS 0.007055f
C489 B.n356 VSUBS 0.007055f
C490 B.n357 VSUBS 0.007055f
C491 B.n358 VSUBS 0.007055f
C492 B.n359 VSUBS 0.007055f
C493 B.n360 VSUBS 0.007055f
C494 B.n361 VSUBS 0.007055f
C495 B.n362 VSUBS 0.007055f
C496 B.n363 VSUBS 0.007055f
C497 B.n364 VSUBS 0.007055f
C498 B.n365 VSUBS 0.007055f
C499 B.n366 VSUBS 0.007055f
C500 B.n367 VSUBS 0.007055f
C501 B.n368 VSUBS 0.007055f
C502 B.n369 VSUBS 0.007055f
C503 B.n370 VSUBS 0.007055f
C504 B.n371 VSUBS 0.007055f
C505 B.n372 VSUBS 0.007055f
C506 B.n373 VSUBS 0.007055f
C507 B.n374 VSUBS 0.007055f
C508 B.n375 VSUBS 0.007055f
C509 B.n376 VSUBS 0.007055f
C510 B.n377 VSUBS 0.007055f
C511 B.n378 VSUBS 0.007055f
C512 B.n379 VSUBS 0.007055f
C513 B.n380 VSUBS 0.007055f
C514 B.n381 VSUBS 0.007055f
C515 B.n382 VSUBS 0.007055f
C516 B.n383 VSUBS 0.007055f
C517 B.n384 VSUBS 0.007055f
C518 B.n385 VSUBS 0.007055f
C519 B.n386 VSUBS 0.007055f
C520 B.n387 VSUBS 0.007055f
C521 B.n388 VSUBS 0.007055f
C522 B.n389 VSUBS 0.007055f
C523 B.n390 VSUBS 0.007055f
C524 B.n391 VSUBS 0.007055f
C525 B.n392 VSUBS 0.007055f
C526 B.n393 VSUBS 0.007055f
C527 B.n394 VSUBS 0.007055f
C528 B.n395 VSUBS 0.007055f
C529 B.n396 VSUBS 0.007055f
C530 B.n397 VSUBS 0.007055f
C531 B.n398 VSUBS 0.007055f
C532 B.n399 VSUBS 0.007055f
C533 B.n400 VSUBS 0.007055f
C534 B.n401 VSUBS 0.007055f
C535 B.n402 VSUBS 0.007055f
C536 B.n403 VSUBS 0.007055f
C537 B.n404 VSUBS 0.007055f
C538 B.n405 VSUBS 0.007055f
C539 B.n406 VSUBS 0.007055f
C540 B.n407 VSUBS 0.007055f
C541 B.n408 VSUBS 0.015947f
C542 B.n409 VSUBS 0.016798f
C543 B.n410 VSUBS 0.015781f
C544 B.n411 VSUBS 0.007055f
C545 B.n412 VSUBS 0.007055f
C546 B.n413 VSUBS 0.007055f
C547 B.n414 VSUBS 0.007055f
C548 B.n415 VSUBS 0.007055f
C549 B.n416 VSUBS 0.007055f
C550 B.n417 VSUBS 0.007055f
C551 B.n418 VSUBS 0.007055f
C552 B.n419 VSUBS 0.007055f
C553 B.n420 VSUBS 0.007055f
C554 B.n421 VSUBS 0.007055f
C555 B.n422 VSUBS 0.007055f
C556 B.n423 VSUBS 0.007055f
C557 B.n424 VSUBS 0.007055f
C558 B.n425 VSUBS 0.007055f
C559 B.n426 VSUBS 0.007055f
C560 B.n427 VSUBS 0.007055f
C561 B.n428 VSUBS 0.007055f
C562 B.n429 VSUBS 0.007055f
C563 B.n430 VSUBS 0.007055f
C564 B.n431 VSUBS 0.007055f
C565 B.n432 VSUBS 0.007055f
C566 B.n433 VSUBS 0.007055f
C567 B.n434 VSUBS 0.007055f
C568 B.n435 VSUBS 0.007055f
C569 B.n436 VSUBS 0.007055f
C570 B.n437 VSUBS 0.007055f
C571 B.n438 VSUBS 0.007055f
C572 B.n439 VSUBS 0.007055f
C573 B.n440 VSUBS 0.007055f
C574 B.n441 VSUBS 0.007055f
C575 B.n442 VSUBS 0.007055f
C576 B.n443 VSUBS 0.007055f
C577 B.n444 VSUBS 0.007055f
C578 B.n445 VSUBS 0.007055f
C579 B.n446 VSUBS 0.007055f
C580 B.n447 VSUBS 0.007055f
C581 B.n448 VSUBS 0.007055f
C582 B.n449 VSUBS 0.007055f
C583 B.n450 VSUBS 0.007055f
C584 B.n451 VSUBS 0.007055f
C585 B.n452 VSUBS 0.007055f
C586 B.n453 VSUBS 0.007055f
C587 B.n454 VSUBS 0.007055f
C588 B.n455 VSUBS 0.007055f
C589 B.n456 VSUBS 0.007055f
C590 B.n457 VSUBS 0.007055f
C591 B.n458 VSUBS 0.007055f
C592 B.n459 VSUBS 0.007055f
C593 B.n460 VSUBS 0.007055f
C594 B.n461 VSUBS 0.007055f
C595 B.n462 VSUBS 0.007055f
C596 B.n463 VSUBS 0.007055f
C597 B.n464 VSUBS 0.007055f
C598 B.n465 VSUBS 0.007055f
C599 B.n466 VSUBS 0.007055f
C600 B.n467 VSUBS 0.007055f
C601 B.n468 VSUBS 0.007055f
C602 B.n469 VSUBS 0.007055f
C603 B.n470 VSUBS 0.007055f
C604 B.n471 VSUBS 0.007055f
C605 B.n472 VSUBS 0.007055f
C606 B.n473 VSUBS 0.007055f
C607 B.n474 VSUBS 0.007055f
C608 B.n475 VSUBS 0.007055f
C609 B.n476 VSUBS 0.004876f
C610 B.n477 VSUBS 0.016346f
C611 B.n478 VSUBS 0.005706f
C612 B.n479 VSUBS 0.007055f
C613 B.n480 VSUBS 0.007055f
C614 B.n481 VSUBS 0.007055f
C615 B.n482 VSUBS 0.007055f
C616 B.n483 VSUBS 0.007055f
C617 B.n484 VSUBS 0.007055f
C618 B.n485 VSUBS 0.007055f
C619 B.n486 VSUBS 0.007055f
C620 B.n487 VSUBS 0.007055f
C621 B.n488 VSUBS 0.007055f
C622 B.n489 VSUBS 0.007055f
C623 B.n490 VSUBS 0.005706f
C624 B.n491 VSUBS 0.007055f
C625 B.n492 VSUBS 0.007055f
C626 B.n493 VSUBS 0.004876f
C627 B.n494 VSUBS 0.007055f
C628 B.n495 VSUBS 0.007055f
C629 B.n496 VSUBS 0.007055f
C630 B.n497 VSUBS 0.007055f
C631 B.n498 VSUBS 0.007055f
C632 B.n499 VSUBS 0.007055f
C633 B.n500 VSUBS 0.007055f
C634 B.n501 VSUBS 0.007055f
C635 B.n502 VSUBS 0.007055f
C636 B.n503 VSUBS 0.007055f
C637 B.n504 VSUBS 0.007055f
C638 B.n505 VSUBS 0.007055f
C639 B.n506 VSUBS 0.007055f
C640 B.n507 VSUBS 0.007055f
C641 B.n508 VSUBS 0.007055f
C642 B.n509 VSUBS 0.007055f
C643 B.n510 VSUBS 0.007055f
C644 B.n511 VSUBS 0.007055f
C645 B.n512 VSUBS 0.007055f
C646 B.n513 VSUBS 0.007055f
C647 B.n514 VSUBS 0.007055f
C648 B.n515 VSUBS 0.007055f
C649 B.n516 VSUBS 0.007055f
C650 B.n517 VSUBS 0.007055f
C651 B.n518 VSUBS 0.007055f
C652 B.n519 VSUBS 0.007055f
C653 B.n520 VSUBS 0.007055f
C654 B.n521 VSUBS 0.007055f
C655 B.n522 VSUBS 0.007055f
C656 B.n523 VSUBS 0.007055f
C657 B.n524 VSUBS 0.007055f
C658 B.n525 VSUBS 0.007055f
C659 B.n526 VSUBS 0.007055f
C660 B.n527 VSUBS 0.007055f
C661 B.n528 VSUBS 0.007055f
C662 B.n529 VSUBS 0.007055f
C663 B.n530 VSUBS 0.007055f
C664 B.n531 VSUBS 0.007055f
C665 B.n532 VSUBS 0.007055f
C666 B.n533 VSUBS 0.007055f
C667 B.n534 VSUBS 0.007055f
C668 B.n535 VSUBS 0.007055f
C669 B.n536 VSUBS 0.007055f
C670 B.n537 VSUBS 0.007055f
C671 B.n538 VSUBS 0.007055f
C672 B.n539 VSUBS 0.007055f
C673 B.n540 VSUBS 0.007055f
C674 B.n541 VSUBS 0.007055f
C675 B.n542 VSUBS 0.007055f
C676 B.n543 VSUBS 0.007055f
C677 B.n544 VSUBS 0.007055f
C678 B.n545 VSUBS 0.007055f
C679 B.n546 VSUBS 0.007055f
C680 B.n547 VSUBS 0.007055f
C681 B.n548 VSUBS 0.007055f
C682 B.n549 VSUBS 0.007055f
C683 B.n550 VSUBS 0.007055f
C684 B.n551 VSUBS 0.007055f
C685 B.n552 VSUBS 0.007055f
C686 B.n553 VSUBS 0.007055f
C687 B.n554 VSUBS 0.007055f
C688 B.n555 VSUBS 0.007055f
C689 B.n556 VSUBS 0.007055f
C690 B.n557 VSUBS 0.007055f
C691 B.n558 VSUBS 0.016632f
C692 B.n559 VSUBS 0.016632f
C693 B.n560 VSUBS 0.015947f
C694 B.n561 VSUBS 0.007055f
C695 B.n562 VSUBS 0.007055f
C696 B.n563 VSUBS 0.007055f
C697 B.n564 VSUBS 0.007055f
C698 B.n565 VSUBS 0.007055f
C699 B.n566 VSUBS 0.007055f
C700 B.n567 VSUBS 0.007055f
C701 B.n568 VSUBS 0.007055f
C702 B.n569 VSUBS 0.007055f
C703 B.n570 VSUBS 0.007055f
C704 B.n571 VSUBS 0.007055f
C705 B.n572 VSUBS 0.007055f
C706 B.n573 VSUBS 0.007055f
C707 B.n574 VSUBS 0.007055f
C708 B.n575 VSUBS 0.007055f
C709 B.n576 VSUBS 0.007055f
C710 B.n577 VSUBS 0.007055f
C711 B.n578 VSUBS 0.007055f
C712 B.n579 VSUBS 0.007055f
C713 B.n580 VSUBS 0.007055f
C714 B.n581 VSUBS 0.007055f
C715 B.n582 VSUBS 0.007055f
C716 B.n583 VSUBS 0.007055f
C717 B.n584 VSUBS 0.007055f
C718 B.n585 VSUBS 0.007055f
C719 B.n586 VSUBS 0.007055f
C720 B.n587 VSUBS 0.007055f
C721 B.n588 VSUBS 0.007055f
C722 B.n589 VSUBS 0.007055f
C723 B.n590 VSUBS 0.007055f
C724 B.n591 VSUBS 0.007055f
C725 B.n592 VSUBS 0.007055f
C726 B.n593 VSUBS 0.007055f
C727 B.n594 VSUBS 0.007055f
C728 B.n595 VSUBS 0.015975f
.ends

