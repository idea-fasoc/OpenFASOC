* NGSPICE file created from diff_pair_sample_1193.ext - technology: sky130A

.subckt diff_pair_sample_1193 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=3.4359 pd=18.4 as=0 ps=0 w=8.81 l=1.76
X1 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=3.4359 pd=18.4 as=0 ps=0 w=8.81 l=1.76
X2 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.4359 pd=18.4 as=0 ps=0 w=8.81 l=1.76
X3 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.4359 pd=18.4 as=0 ps=0 w=8.81 l=1.76
X4 VDD1.t1 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=3.4359 pd=18.4 as=3.4359 ps=18.4 w=8.81 l=1.76
X5 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.4359 pd=18.4 as=3.4359 ps=18.4 w=8.81 l=1.76
X6 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=3.4359 pd=18.4 as=3.4359 ps=18.4 w=8.81 l=1.76
X7 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.4359 pd=18.4 as=3.4359 ps=18.4 w=8.81 l=1.76
R0 B.n545 B.n544 585
R1 B.n227 B.n78 585
R2 B.n226 B.n225 585
R3 B.n224 B.n223 585
R4 B.n222 B.n221 585
R5 B.n220 B.n219 585
R6 B.n218 B.n217 585
R7 B.n216 B.n215 585
R8 B.n214 B.n213 585
R9 B.n212 B.n211 585
R10 B.n210 B.n209 585
R11 B.n208 B.n207 585
R12 B.n206 B.n205 585
R13 B.n204 B.n203 585
R14 B.n202 B.n201 585
R15 B.n200 B.n199 585
R16 B.n198 B.n197 585
R17 B.n196 B.n195 585
R18 B.n194 B.n193 585
R19 B.n192 B.n191 585
R20 B.n190 B.n189 585
R21 B.n188 B.n187 585
R22 B.n186 B.n185 585
R23 B.n184 B.n183 585
R24 B.n182 B.n181 585
R25 B.n180 B.n179 585
R26 B.n178 B.n177 585
R27 B.n176 B.n175 585
R28 B.n174 B.n173 585
R29 B.n172 B.n171 585
R30 B.n170 B.n169 585
R31 B.n168 B.n167 585
R32 B.n166 B.n165 585
R33 B.n164 B.n163 585
R34 B.n162 B.n161 585
R35 B.n160 B.n159 585
R36 B.n158 B.n157 585
R37 B.n156 B.n155 585
R38 B.n154 B.n153 585
R39 B.n152 B.n151 585
R40 B.n150 B.n149 585
R41 B.n148 B.n147 585
R42 B.n146 B.n145 585
R43 B.n144 B.n143 585
R44 B.n142 B.n141 585
R45 B.n140 B.n139 585
R46 B.n138 B.n137 585
R47 B.n136 B.n135 585
R48 B.n134 B.n133 585
R49 B.n132 B.n131 585
R50 B.n130 B.n129 585
R51 B.n128 B.n127 585
R52 B.n126 B.n125 585
R53 B.n124 B.n123 585
R54 B.n122 B.n121 585
R55 B.n120 B.n119 585
R56 B.n118 B.n117 585
R57 B.n116 B.n115 585
R58 B.n114 B.n113 585
R59 B.n112 B.n111 585
R60 B.n110 B.n109 585
R61 B.n108 B.n107 585
R62 B.n106 B.n105 585
R63 B.n104 B.n103 585
R64 B.n102 B.n101 585
R65 B.n100 B.n99 585
R66 B.n98 B.n97 585
R67 B.n96 B.n95 585
R68 B.n94 B.n93 585
R69 B.n92 B.n91 585
R70 B.n90 B.n89 585
R71 B.n88 B.n87 585
R72 B.n86 B.n85 585
R73 B.n40 B.n39 585
R74 B.n543 B.n41 585
R75 B.n548 B.n41 585
R76 B.n542 B.n541 585
R77 B.n541 B.n37 585
R78 B.n540 B.n36 585
R79 B.n554 B.n36 585
R80 B.n539 B.n35 585
R81 B.n555 B.n35 585
R82 B.n538 B.n34 585
R83 B.n556 B.n34 585
R84 B.n537 B.n536 585
R85 B.n536 B.n30 585
R86 B.n535 B.n29 585
R87 B.n562 B.n29 585
R88 B.n534 B.n28 585
R89 B.n563 B.n28 585
R90 B.n533 B.n27 585
R91 B.n564 B.n27 585
R92 B.n532 B.n531 585
R93 B.n531 B.n23 585
R94 B.n530 B.n22 585
R95 B.n570 B.n22 585
R96 B.n529 B.n21 585
R97 B.n571 B.n21 585
R98 B.n528 B.n20 585
R99 B.n572 B.n20 585
R100 B.n527 B.n526 585
R101 B.n526 B.n16 585
R102 B.n525 B.n15 585
R103 B.n578 B.n15 585
R104 B.n524 B.n14 585
R105 B.n579 B.n14 585
R106 B.n523 B.n13 585
R107 B.n580 B.n13 585
R108 B.n522 B.n521 585
R109 B.n521 B.n12 585
R110 B.n520 B.n519 585
R111 B.n520 B.n8 585
R112 B.n518 B.n7 585
R113 B.n587 B.n7 585
R114 B.n517 B.n6 585
R115 B.n588 B.n6 585
R116 B.n516 B.n5 585
R117 B.n589 B.n5 585
R118 B.n515 B.n514 585
R119 B.n514 B.n4 585
R120 B.n513 B.n228 585
R121 B.n513 B.n512 585
R122 B.n503 B.n229 585
R123 B.n230 B.n229 585
R124 B.n505 B.n504 585
R125 B.n506 B.n505 585
R126 B.n502 B.n234 585
R127 B.n238 B.n234 585
R128 B.n501 B.n500 585
R129 B.n500 B.n499 585
R130 B.n236 B.n235 585
R131 B.n237 B.n236 585
R132 B.n492 B.n491 585
R133 B.n493 B.n492 585
R134 B.n490 B.n243 585
R135 B.n243 B.n242 585
R136 B.n489 B.n488 585
R137 B.n488 B.n487 585
R138 B.n245 B.n244 585
R139 B.n246 B.n245 585
R140 B.n480 B.n479 585
R141 B.n481 B.n480 585
R142 B.n478 B.n251 585
R143 B.n251 B.n250 585
R144 B.n477 B.n476 585
R145 B.n476 B.n475 585
R146 B.n253 B.n252 585
R147 B.n254 B.n253 585
R148 B.n468 B.n467 585
R149 B.n469 B.n468 585
R150 B.n466 B.n259 585
R151 B.n259 B.n258 585
R152 B.n465 B.n464 585
R153 B.n464 B.n463 585
R154 B.n261 B.n260 585
R155 B.n262 B.n261 585
R156 B.n456 B.n455 585
R157 B.n457 B.n456 585
R158 B.n265 B.n264 585
R159 B.n308 B.n306 585
R160 B.n309 B.n305 585
R161 B.n309 B.n266 585
R162 B.n312 B.n311 585
R163 B.n313 B.n304 585
R164 B.n315 B.n314 585
R165 B.n317 B.n303 585
R166 B.n320 B.n319 585
R167 B.n321 B.n302 585
R168 B.n323 B.n322 585
R169 B.n325 B.n301 585
R170 B.n328 B.n327 585
R171 B.n329 B.n300 585
R172 B.n331 B.n330 585
R173 B.n333 B.n299 585
R174 B.n336 B.n335 585
R175 B.n337 B.n298 585
R176 B.n339 B.n338 585
R177 B.n341 B.n297 585
R178 B.n344 B.n343 585
R179 B.n345 B.n296 585
R180 B.n347 B.n346 585
R181 B.n349 B.n295 585
R182 B.n352 B.n351 585
R183 B.n353 B.n294 585
R184 B.n355 B.n354 585
R185 B.n357 B.n293 585
R186 B.n360 B.n359 585
R187 B.n361 B.n292 585
R188 B.n363 B.n362 585
R189 B.n365 B.n291 585
R190 B.n368 B.n367 585
R191 B.n370 B.n288 585
R192 B.n372 B.n371 585
R193 B.n374 B.n287 585
R194 B.n377 B.n376 585
R195 B.n378 B.n286 585
R196 B.n380 B.n379 585
R197 B.n382 B.n285 585
R198 B.n385 B.n384 585
R199 B.n386 B.n284 585
R200 B.n391 B.n390 585
R201 B.n393 B.n283 585
R202 B.n396 B.n395 585
R203 B.n397 B.n282 585
R204 B.n399 B.n398 585
R205 B.n401 B.n281 585
R206 B.n404 B.n403 585
R207 B.n405 B.n280 585
R208 B.n407 B.n406 585
R209 B.n409 B.n279 585
R210 B.n412 B.n411 585
R211 B.n413 B.n278 585
R212 B.n415 B.n414 585
R213 B.n417 B.n277 585
R214 B.n420 B.n419 585
R215 B.n421 B.n276 585
R216 B.n423 B.n422 585
R217 B.n425 B.n275 585
R218 B.n428 B.n427 585
R219 B.n429 B.n274 585
R220 B.n431 B.n430 585
R221 B.n433 B.n273 585
R222 B.n436 B.n435 585
R223 B.n437 B.n272 585
R224 B.n439 B.n438 585
R225 B.n441 B.n271 585
R226 B.n444 B.n443 585
R227 B.n445 B.n270 585
R228 B.n447 B.n446 585
R229 B.n449 B.n269 585
R230 B.n450 B.n268 585
R231 B.n453 B.n452 585
R232 B.n454 B.n267 585
R233 B.n267 B.n266 585
R234 B.n459 B.n458 585
R235 B.n458 B.n457 585
R236 B.n460 B.n263 585
R237 B.n263 B.n262 585
R238 B.n462 B.n461 585
R239 B.n463 B.n462 585
R240 B.n257 B.n256 585
R241 B.n258 B.n257 585
R242 B.n471 B.n470 585
R243 B.n470 B.n469 585
R244 B.n472 B.n255 585
R245 B.n255 B.n254 585
R246 B.n474 B.n473 585
R247 B.n475 B.n474 585
R248 B.n249 B.n248 585
R249 B.n250 B.n249 585
R250 B.n483 B.n482 585
R251 B.n482 B.n481 585
R252 B.n484 B.n247 585
R253 B.n247 B.n246 585
R254 B.n486 B.n485 585
R255 B.n487 B.n486 585
R256 B.n241 B.n240 585
R257 B.n242 B.n241 585
R258 B.n495 B.n494 585
R259 B.n494 B.n493 585
R260 B.n496 B.n239 585
R261 B.n239 B.n237 585
R262 B.n498 B.n497 585
R263 B.n499 B.n498 585
R264 B.n233 B.n232 585
R265 B.n238 B.n233 585
R266 B.n508 B.n507 585
R267 B.n507 B.n506 585
R268 B.n509 B.n231 585
R269 B.n231 B.n230 585
R270 B.n511 B.n510 585
R271 B.n512 B.n511 585
R272 B.n3 B.n0 585
R273 B.n4 B.n3 585
R274 B.n586 B.n1 585
R275 B.n587 B.n586 585
R276 B.n585 B.n584 585
R277 B.n585 B.n8 585
R278 B.n583 B.n9 585
R279 B.n12 B.n9 585
R280 B.n582 B.n581 585
R281 B.n581 B.n580 585
R282 B.n11 B.n10 585
R283 B.n579 B.n11 585
R284 B.n577 B.n576 585
R285 B.n578 B.n577 585
R286 B.n575 B.n17 585
R287 B.n17 B.n16 585
R288 B.n574 B.n573 585
R289 B.n573 B.n572 585
R290 B.n19 B.n18 585
R291 B.n571 B.n19 585
R292 B.n569 B.n568 585
R293 B.n570 B.n569 585
R294 B.n567 B.n24 585
R295 B.n24 B.n23 585
R296 B.n566 B.n565 585
R297 B.n565 B.n564 585
R298 B.n26 B.n25 585
R299 B.n563 B.n26 585
R300 B.n561 B.n560 585
R301 B.n562 B.n561 585
R302 B.n559 B.n31 585
R303 B.n31 B.n30 585
R304 B.n558 B.n557 585
R305 B.n557 B.n556 585
R306 B.n33 B.n32 585
R307 B.n555 B.n33 585
R308 B.n553 B.n552 585
R309 B.n554 B.n553 585
R310 B.n551 B.n38 585
R311 B.n38 B.n37 585
R312 B.n550 B.n549 585
R313 B.n549 B.n548 585
R314 B.n590 B.n589 585
R315 B.n588 B.n2 585
R316 B.n549 B.n40 487.695
R317 B.n545 B.n41 487.695
R318 B.n456 B.n267 487.695
R319 B.n458 B.n265 487.695
R320 B.n82 B.t6 326.93
R321 B.n79 B.t13 326.93
R322 B.n387 B.t2 326.93
R323 B.n289 B.t10 326.93
R324 B.n79 B.t14 268.055
R325 B.n387 B.t5 268.055
R326 B.n82 B.t8 268.055
R327 B.n289 B.t12 268.055
R328 B.n547 B.n546 256.663
R329 B.n547 B.n77 256.663
R330 B.n547 B.n76 256.663
R331 B.n547 B.n75 256.663
R332 B.n547 B.n74 256.663
R333 B.n547 B.n73 256.663
R334 B.n547 B.n72 256.663
R335 B.n547 B.n71 256.663
R336 B.n547 B.n70 256.663
R337 B.n547 B.n69 256.663
R338 B.n547 B.n68 256.663
R339 B.n547 B.n67 256.663
R340 B.n547 B.n66 256.663
R341 B.n547 B.n65 256.663
R342 B.n547 B.n64 256.663
R343 B.n547 B.n63 256.663
R344 B.n547 B.n62 256.663
R345 B.n547 B.n61 256.663
R346 B.n547 B.n60 256.663
R347 B.n547 B.n59 256.663
R348 B.n547 B.n58 256.663
R349 B.n547 B.n57 256.663
R350 B.n547 B.n56 256.663
R351 B.n547 B.n55 256.663
R352 B.n547 B.n54 256.663
R353 B.n547 B.n53 256.663
R354 B.n547 B.n52 256.663
R355 B.n547 B.n51 256.663
R356 B.n547 B.n50 256.663
R357 B.n547 B.n49 256.663
R358 B.n547 B.n48 256.663
R359 B.n547 B.n47 256.663
R360 B.n547 B.n46 256.663
R361 B.n547 B.n45 256.663
R362 B.n547 B.n44 256.663
R363 B.n547 B.n43 256.663
R364 B.n547 B.n42 256.663
R365 B.n307 B.n266 256.663
R366 B.n310 B.n266 256.663
R367 B.n316 B.n266 256.663
R368 B.n318 B.n266 256.663
R369 B.n324 B.n266 256.663
R370 B.n326 B.n266 256.663
R371 B.n332 B.n266 256.663
R372 B.n334 B.n266 256.663
R373 B.n340 B.n266 256.663
R374 B.n342 B.n266 256.663
R375 B.n348 B.n266 256.663
R376 B.n350 B.n266 256.663
R377 B.n356 B.n266 256.663
R378 B.n358 B.n266 256.663
R379 B.n364 B.n266 256.663
R380 B.n366 B.n266 256.663
R381 B.n373 B.n266 256.663
R382 B.n375 B.n266 256.663
R383 B.n381 B.n266 256.663
R384 B.n383 B.n266 256.663
R385 B.n392 B.n266 256.663
R386 B.n394 B.n266 256.663
R387 B.n400 B.n266 256.663
R388 B.n402 B.n266 256.663
R389 B.n408 B.n266 256.663
R390 B.n410 B.n266 256.663
R391 B.n416 B.n266 256.663
R392 B.n418 B.n266 256.663
R393 B.n424 B.n266 256.663
R394 B.n426 B.n266 256.663
R395 B.n432 B.n266 256.663
R396 B.n434 B.n266 256.663
R397 B.n440 B.n266 256.663
R398 B.n442 B.n266 256.663
R399 B.n448 B.n266 256.663
R400 B.n451 B.n266 256.663
R401 B.n592 B.n591 256.663
R402 B.n80 B.t15 227.522
R403 B.n388 B.t4 227.522
R404 B.n83 B.t9 227.522
R405 B.n290 B.t11 227.522
R406 B.n87 B.n86 163.367
R407 B.n91 B.n90 163.367
R408 B.n95 B.n94 163.367
R409 B.n99 B.n98 163.367
R410 B.n103 B.n102 163.367
R411 B.n107 B.n106 163.367
R412 B.n111 B.n110 163.367
R413 B.n115 B.n114 163.367
R414 B.n119 B.n118 163.367
R415 B.n123 B.n122 163.367
R416 B.n127 B.n126 163.367
R417 B.n131 B.n130 163.367
R418 B.n135 B.n134 163.367
R419 B.n139 B.n138 163.367
R420 B.n143 B.n142 163.367
R421 B.n147 B.n146 163.367
R422 B.n151 B.n150 163.367
R423 B.n155 B.n154 163.367
R424 B.n159 B.n158 163.367
R425 B.n163 B.n162 163.367
R426 B.n167 B.n166 163.367
R427 B.n171 B.n170 163.367
R428 B.n175 B.n174 163.367
R429 B.n179 B.n178 163.367
R430 B.n183 B.n182 163.367
R431 B.n187 B.n186 163.367
R432 B.n191 B.n190 163.367
R433 B.n195 B.n194 163.367
R434 B.n199 B.n198 163.367
R435 B.n203 B.n202 163.367
R436 B.n207 B.n206 163.367
R437 B.n211 B.n210 163.367
R438 B.n215 B.n214 163.367
R439 B.n219 B.n218 163.367
R440 B.n223 B.n222 163.367
R441 B.n225 B.n78 163.367
R442 B.n456 B.n261 163.367
R443 B.n464 B.n261 163.367
R444 B.n464 B.n259 163.367
R445 B.n468 B.n259 163.367
R446 B.n468 B.n253 163.367
R447 B.n476 B.n253 163.367
R448 B.n476 B.n251 163.367
R449 B.n480 B.n251 163.367
R450 B.n480 B.n245 163.367
R451 B.n488 B.n245 163.367
R452 B.n488 B.n243 163.367
R453 B.n492 B.n243 163.367
R454 B.n492 B.n236 163.367
R455 B.n500 B.n236 163.367
R456 B.n500 B.n234 163.367
R457 B.n505 B.n234 163.367
R458 B.n505 B.n229 163.367
R459 B.n513 B.n229 163.367
R460 B.n514 B.n513 163.367
R461 B.n514 B.n5 163.367
R462 B.n6 B.n5 163.367
R463 B.n7 B.n6 163.367
R464 B.n520 B.n7 163.367
R465 B.n521 B.n520 163.367
R466 B.n521 B.n13 163.367
R467 B.n14 B.n13 163.367
R468 B.n15 B.n14 163.367
R469 B.n526 B.n15 163.367
R470 B.n526 B.n20 163.367
R471 B.n21 B.n20 163.367
R472 B.n22 B.n21 163.367
R473 B.n531 B.n22 163.367
R474 B.n531 B.n27 163.367
R475 B.n28 B.n27 163.367
R476 B.n29 B.n28 163.367
R477 B.n536 B.n29 163.367
R478 B.n536 B.n34 163.367
R479 B.n35 B.n34 163.367
R480 B.n36 B.n35 163.367
R481 B.n541 B.n36 163.367
R482 B.n541 B.n41 163.367
R483 B.n309 B.n308 163.367
R484 B.n311 B.n309 163.367
R485 B.n315 B.n304 163.367
R486 B.n319 B.n317 163.367
R487 B.n323 B.n302 163.367
R488 B.n327 B.n325 163.367
R489 B.n331 B.n300 163.367
R490 B.n335 B.n333 163.367
R491 B.n339 B.n298 163.367
R492 B.n343 B.n341 163.367
R493 B.n347 B.n296 163.367
R494 B.n351 B.n349 163.367
R495 B.n355 B.n294 163.367
R496 B.n359 B.n357 163.367
R497 B.n363 B.n292 163.367
R498 B.n367 B.n365 163.367
R499 B.n372 B.n288 163.367
R500 B.n376 B.n374 163.367
R501 B.n380 B.n286 163.367
R502 B.n384 B.n382 163.367
R503 B.n391 B.n284 163.367
R504 B.n395 B.n393 163.367
R505 B.n399 B.n282 163.367
R506 B.n403 B.n401 163.367
R507 B.n407 B.n280 163.367
R508 B.n411 B.n409 163.367
R509 B.n415 B.n278 163.367
R510 B.n419 B.n417 163.367
R511 B.n423 B.n276 163.367
R512 B.n427 B.n425 163.367
R513 B.n431 B.n274 163.367
R514 B.n435 B.n433 163.367
R515 B.n439 B.n272 163.367
R516 B.n443 B.n441 163.367
R517 B.n447 B.n270 163.367
R518 B.n450 B.n449 163.367
R519 B.n452 B.n267 163.367
R520 B.n458 B.n263 163.367
R521 B.n462 B.n263 163.367
R522 B.n462 B.n257 163.367
R523 B.n470 B.n257 163.367
R524 B.n470 B.n255 163.367
R525 B.n474 B.n255 163.367
R526 B.n474 B.n249 163.367
R527 B.n482 B.n249 163.367
R528 B.n482 B.n247 163.367
R529 B.n486 B.n247 163.367
R530 B.n486 B.n241 163.367
R531 B.n494 B.n241 163.367
R532 B.n494 B.n239 163.367
R533 B.n498 B.n239 163.367
R534 B.n498 B.n233 163.367
R535 B.n507 B.n233 163.367
R536 B.n507 B.n231 163.367
R537 B.n511 B.n231 163.367
R538 B.n511 B.n3 163.367
R539 B.n590 B.n3 163.367
R540 B.n586 B.n2 163.367
R541 B.n586 B.n585 163.367
R542 B.n585 B.n9 163.367
R543 B.n581 B.n9 163.367
R544 B.n581 B.n11 163.367
R545 B.n577 B.n11 163.367
R546 B.n577 B.n17 163.367
R547 B.n573 B.n17 163.367
R548 B.n573 B.n19 163.367
R549 B.n569 B.n19 163.367
R550 B.n569 B.n24 163.367
R551 B.n565 B.n24 163.367
R552 B.n565 B.n26 163.367
R553 B.n561 B.n26 163.367
R554 B.n561 B.n31 163.367
R555 B.n557 B.n31 163.367
R556 B.n557 B.n33 163.367
R557 B.n553 B.n33 163.367
R558 B.n553 B.n38 163.367
R559 B.n549 B.n38 163.367
R560 B.n457 B.n266 91.3743
R561 B.n548 B.n547 91.3743
R562 B.n42 B.n40 71.676
R563 B.n87 B.n43 71.676
R564 B.n91 B.n44 71.676
R565 B.n95 B.n45 71.676
R566 B.n99 B.n46 71.676
R567 B.n103 B.n47 71.676
R568 B.n107 B.n48 71.676
R569 B.n111 B.n49 71.676
R570 B.n115 B.n50 71.676
R571 B.n119 B.n51 71.676
R572 B.n123 B.n52 71.676
R573 B.n127 B.n53 71.676
R574 B.n131 B.n54 71.676
R575 B.n135 B.n55 71.676
R576 B.n139 B.n56 71.676
R577 B.n143 B.n57 71.676
R578 B.n147 B.n58 71.676
R579 B.n151 B.n59 71.676
R580 B.n155 B.n60 71.676
R581 B.n159 B.n61 71.676
R582 B.n163 B.n62 71.676
R583 B.n167 B.n63 71.676
R584 B.n171 B.n64 71.676
R585 B.n175 B.n65 71.676
R586 B.n179 B.n66 71.676
R587 B.n183 B.n67 71.676
R588 B.n187 B.n68 71.676
R589 B.n191 B.n69 71.676
R590 B.n195 B.n70 71.676
R591 B.n199 B.n71 71.676
R592 B.n203 B.n72 71.676
R593 B.n207 B.n73 71.676
R594 B.n211 B.n74 71.676
R595 B.n215 B.n75 71.676
R596 B.n219 B.n76 71.676
R597 B.n223 B.n77 71.676
R598 B.n546 B.n78 71.676
R599 B.n546 B.n545 71.676
R600 B.n225 B.n77 71.676
R601 B.n222 B.n76 71.676
R602 B.n218 B.n75 71.676
R603 B.n214 B.n74 71.676
R604 B.n210 B.n73 71.676
R605 B.n206 B.n72 71.676
R606 B.n202 B.n71 71.676
R607 B.n198 B.n70 71.676
R608 B.n194 B.n69 71.676
R609 B.n190 B.n68 71.676
R610 B.n186 B.n67 71.676
R611 B.n182 B.n66 71.676
R612 B.n178 B.n65 71.676
R613 B.n174 B.n64 71.676
R614 B.n170 B.n63 71.676
R615 B.n166 B.n62 71.676
R616 B.n162 B.n61 71.676
R617 B.n158 B.n60 71.676
R618 B.n154 B.n59 71.676
R619 B.n150 B.n58 71.676
R620 B.n146 B.n57 71.676
R621 B.n142 B.n56 71.676
R622 B.n138 B.n55 71.676
R623 B.n134 B.n54 71.676
R624 B.n130 B.n53 71.676
R625 B.n126 B.n52 71.676
R626 B.n122 B.n51 71.676
R627 B.n118 B.n50 71.676
R628 B.n114 B.n49 71.676
R629 B.n110 B.n48 71.676
R630 B.n106 B.n47 71.676
R631 B.n102 B.n46 71.676
R632 B.n98 B.n45 71.676
R633 B.n94 B.n44 71.676
R634 B.n90 B.n43 71.676
R635 B.n86 B.n42 71.676
R636 B.n307 B.n265 71.676
R637 B.n311 B.n310 71.676
R638 B.n316 B.n315 71.676
R639 B.n319 B.n318 71.676
R640 B.n324 B.n323 71.676
R641 B.n327 B.n326 71.676
R642 B.n332 B.n331 71.676
R643 B.n335 B.n334 71.676
R644 B.n340 B.n339 71.676
R645 B.n343 B.n342 71.676
R646 B.n348 B.n347 71.676
R647 B.n351 B.n350 71.676
R648 B.n356 B.n355 71.676
R649 B.n359 B.n358 71.676
R650 B.n364 B.n363 71.676
R651 B.n367 B.n366 71.676
R652 B.n373 B.n372 71.676
R653 B.n376 B.n375 71.676
R654 B.n381 B.n380 71.676
R655 B.n384 B.n383 71.676
R656 B.n392 B.n391 71.676
R657 B.n395 B.n394 71.676
R658 B.n400 B.n399 71.676
R659 B.n403 B.n402 71.676
R660 B.n408 B.n407 71.676
R661 B.n411 B.n410 71.676
R662 B.n416 B.n415 71.676
R663 B.n419 B.n418 71.676
R664 B.n424 B.n423 71.676
R665 B.n427 B.n426 71.676
R666 B.n432 B.n431 71.676
R667 B.n435 B.n434 71.676
R668 B.n440 B.n439 71.676
R669 B.n443 B.n442 71.676
R670 B.n448 B.n447 71.676
R671 B.n451 B.n450 71.676
R672 B.n308 B.n307 71.676
R673 B.n310 B.n304 71.676
R674 B.n317 B.n316 71.676
R675 B.n318 B.n302 71.676
R676 B.n325 B.n324 71.676
R677 B.n326 B.n300 71.676
R678 B.n333 B.n332 71.676
R679 B.n334 B.n298 71.676
R680 B.n341 B.n340 71.676
R681 B.n342 B.n296 71.676
R682 B.n349 B.n348 71.676
R683 B.n350 B.n294 71.676
R684 B.n357 B.n356 71.676
R685 B.n358 B.n292 71.676
R686 B.n365 B.n364 71.676
R687 B.n366 B.n288 71.676
R688 B.n374 B.n373 71.676
R689 B.n375 B.n286 71.676
R690 B.n382 B.n381 71.676
R691 B.n383 B.n284 71.676
R692 B.n393 B.n392 71.676
R693 B.n394 B.n282 71.676
R694 B.n401 B.n400 71.676
R695 B.n402 B.n280 71.676
R696 B.n409 B.n408 71.676
R697 B.n410 B.n278 71.676
R698 B.n417 B.n416 71.676
R699 B.n418 B.n276 71.676
R700 B.n425 B.n424 71.676
R701 B.n426 B.n274 71.676
R702 B.n433 B.n432 71.676
R703 B.n434 B.n272 71.676
R704 B.n441 B.n440 71.676
R705 B.n442 B.n270 71.676
R706 B.n449 B.n448 71.676
R707 B.n452 B.n451 71.676
R708 B.n591 B.n590 71.676
R709 B.n591 B.n2 71.676
R710 B.n84 B.n83 59.5399
R711 B.n81 B.n80 59.5399
R712 B.n389 B.n388 59.5399
R713 B.n369 B.n290 59.5399
R714 B.n457 B.n262 53.1066
R715 B.n463 B.n262 53.1066
R716 B.n463 B.n258 53.1066
R717 B.n469 B.n258 53.1066
R718 B.n469 B.n254 53.1066
R719 B.n475 B.n254 53.1066
R720 B.n481 B.n250 53.1066
R721 B.n481 B.n246 53.1066
R722 B.n487 B.n246 53.1066
R723 B.n487 B.n242 53.1066
R724 B.n493 B.n242 53.1066
R725 B.n493 B.n237 53.1066
R726 B.n499 B.n237 53.1066
R727 B.n499 B.n238 53.1066
R728 B.n506 B.n230 53.1066
R729 B.n512 B.n230 53.1066
R730 B.n512 B.n4 53.1066
R731 B.n589 B.n4 53.1066
R732 B.n589 B.n588 53.1066
R733 B.n588 B.n587 53.1066
R734 B.n587 B.n8 53.1066
R735 B.n12 B.n8 53.1066
R736 B.n580 B.n12 53.1066
R737 B.n579 B.n578 53.1066
R738 B.n578 B.n16 53.1066
R739 B.n572 B.n16 53.1066
R740 B.n572 B.n571 53.1066
R741 B.n571 B.n570 53.1066
R742 B.n570 B.n23 53.1066
R743 B.n564 B.n23 53.1066
R744 B.n564 B.n563 53.1066
R745 B.n562 B.n30 53.1066
R746 B.n556 B.n30 53.1066
R747 B.n556 B.n555 53.1066
R748 B.n555 B.n554 53.1066
R749 B.n554 B.n37 53.1066
R750 B.n548 B.n37 53.1066
R751 B.n238 B.t0 43.735
R752 B.t1 B.n579 43.735
R753 B.n83 B.n82 40.5338
R754 B.n80 B.n79 40.5338
R755 B.n388 B.n387 40.5338
R756 B.n290 B.n289 40.5338
R757 B.n459 B.n264 31.6883
R758 B.n455 B.n454 31.6883
R759 B.n544 B.n543 31.6883
R760 B.n550 B.n39 31.6883
R761 B.t3 B.n250 28.1155
R762 B.n563 B.t7 28.1155
R763 B.n475 B.t3 24.9916
R764 B.t7 B.n562 24.9916
R765 B B.n592 18.0485
R766 B.n460 B.n459 10.6151
R767 B.n461 B.n460 10.6151
R768 B.n461 B.n256 10.6151
R769 B.n471 B.n256 10.6151
R770 B.n472 B.n471 10.6151
R771 B.n473 B.n472 10.6151
R772 B.n473 B.n248 10.6151
R773 B.n483 B.n248 10.6151
R774 B.n484 B.n483 10.6151
R775 B.n485 B.n484 10.6151
R776 B.n485 B.n240 10.6151
R777 B.n495 B.n240 10.6151
R778 B.n496 B.n495 10.6151
R779 B.n497 B.n496 10.6151
R780 B.n497 B.n232 10.6151
R781 B.n508 B.n232 10.6151
R782 B.n509 B.n508 10.6151
R783 B.n510 B.n509 10.6151
R784 B.n510 B.n0 10.6151
R785 B.n306 B.n264 10.6151
R786 B.n306 B.n305 10.6151
R787 B.n312 B.n305 10.6151
R788 B.n313 B.n312 10.6151
R789 B.n314 B.n313 10.6151
R790 B.n314 B.n303 10.6151
R791 B.n320 B.n303 10.6151
R792 B.n321 B.n320 10.6151
R793 B.n322 B.n321 10.6151
R794 B.n322 B.n301 10.6151
R795 B.n328 B.n301 10.6151
R796 B.n329 B.n328 10.6151
R797 B.n330 B.n329 10.6151
R798 B.n330 B.n299 10.6151
R799 B.n336 B.n299 10.6151
R800 B.n337 B.n336 10.6151
R801 B.n338 B.n337 10.6151
R802 B.n338 B.n297 10.6151
R803 B.n344 B.n297 10.6151
R804 B.n345 B.n344 10.6151
R805 B.n346 B.n345 10.6151
R806 B.n346 B.n295 10.6151
R807 B.n352 B.n295 10.6151
R808 B.n353 B.n352 10.6151
R809 B.n354 B.n353 10.6151
R810 B.n354 B.n293 10.6151
R811 B.n360 B.n293 10.6151
R812 B.n361 B.n360 10.6151
R813 B.n362 B.n361 10.6151
R814 B.n362 B.n291 10.6151
R815 B.n368 B.n291 10.6151
R816 B.n371 B.n370 10.6151
R817 B.n371 B.n287 10.6151
R818 B.n377 B.n287 10.6151
R819 B.n378 B.n377 10.6151
R820 B.n379 B.n378 10.6151
R821 B.n379 B.n285 10.6151
R822 B.n385 B.n285 10.6151
R823 B.n386 B.n385 10.6151
R824 B.n390 B.n386 10.6151
R825 B.n396 B.n283 10.6151
R826 B.n397 B.n396 10.6151
R827 B.n398 B.n397 10.6151
R828 B.n398 B.n281 10.6151
R829 B.n404 B.n281 10.6151
R830 B.n405 B.n404 10.6151
R831 B.n406 B.n405 10.6151
R832 B.n406 B.n279 10.6151
R833 B.n412 B.n279 10.6151
R834 B.n413 B.n412 10.6151
R835 B.n414 B.n413 10.6151
R836 B.n414 B.n277 10.6151
R837 B.n420 B.n277 10.6151
R838 B.n421 B.n420 10.6151
R839 B.n422 B.n421 10.6151
R840 B.n422 B.n275 10.6151
R841 B.n428 B.n275 10.6151
R842 B.n429 B.n428 10.6151
R843 B.n430 B.n429 10.6151
R844 B.n430 B.n273 10.6151
R845 B.n436 B.n273 10.6151
R846 B.n437 B.n436 10.6151
R847 B.n438 B.n437 10.6151
R848 B.n438 B.n271 10.6151
R849 B.n444 B.n271 10.6151
R850 B.n445 B.n444 10.6151
R851 B.n446 B.n445 10.6151
R852 B.n446 B.n269 10.6151
R853 B.n269 B.n268 10.6151
R854 B.n453 B.n268 10.6151
R855 B.n454 B.n453 10.6151
R856 B.n455 B.n260 10.6151
R857 B.n465 B.n260 10.6151
R858 B.n466 B.n465 10.6151
R859 B.n467 B.n466 10.6151
R860 B.n467 B.n252 10.6151
R861 B.n477 B.n252 10.6151
R862 B.n478 B.n477 10.6151
R863 B.n479 B.n478 10.6151
R864 B.n479 B.n244 10.6151
R865 B.n489 B.n244 10.6151
R866 B.n490 B.n489 10.6151
R867 B.n491 B.n490 10.6151
R868 B.n491 B.n235 10.6151
R869 B.n501 B.n235 10.6151
R870 B.n502 B.n501 10.6151
R871 B.n504 B.n502 10.6151
R872 B.n504 B.n503 10.6151
R873 B.n503 B.n228 10.6151
R874 B.n515 B.n228 10.6151
R875 B.n516 B.n515 10.6151
R876 B.n517 B.n516 10.6151
R877 B.n518 B.n517 10.6151
R878 B.n519 B.n518 10.6151
R879 B.n522 B.n519 10.6151
R880 B.n523 B.n522 10.6151
R881 B.n524 B.n523 10.6151
R882 B.n525 B.n524 10.6151
R883 B.n527 B.n525 10.6151
R884 B.n528 B.n527 10.6151
R885 B.n529 B.n528 10.6151
R886 B.n530 B.n529 10.6151
R887 B.n532 B.n530 10.6151
R888 B.n533 B.n532 10.6151
R889 B.n534 B.n533 10.6151
R890 B.n535 B.n534 10.6151
R891 B.n537 B.n535 10.6151
R892 B.n538 B.n537 10.6151
R893 B.n539 B.n538 10.6151
R894 B.n540 B.n539 10.6151
R895 B.n542 B.n540 10.6151
R896 B.n543 B.n542 10.6151
R897 B.n584 B.n1 10.6151
R898 B.n584 B.n583 10.6151
R899 B.n583 B.n582 10.6151
R900 B.n582 B.n10 10.6151
R901 B.n576 B.n10 10.6151
R902 B.n576 B.n575 10.6151
R903 B.n575 B.n574 10.6151
R904 B.n574 B.n18 10.6151
R905 B.n568 B.n18 10.6151
R906 B.n568 B.n567 10.6151
R907 B.n567 B.n566 10.6151
R908 B.n566 B.n25 10.6151
R909 B.n560 B.n25 10.6151
R910 B.n560 B.n559 10.6151
R911 B.n559 B.n558 10.6151
R912 B.n558 B.n32 10.6151
R913 B.n552 B.n32 10.6151
R914 B.n552 B.n551 10.6151
R915 B.n551 B.n550 10.6151
R916 B.n85 B.n39 10.6151
R917 B.n88 B.n85 10.6151
R918 B.n89 B.n88 10.6151
R919 B.n92 B.n89 10.6151
R920 B.n93 B.n92 10.6151
R921 B.n96 B.n93 10.6151
R922 B.n97 B.n96 10.6151
R923 B.n100 B.n97 10.6151
R924 B.n101 B.n100 10.6151
R925 B.n104 B.n101 10.6151
R926 B.n105 B.n104 10.6151
R927 B.n108 B.n105 10.6151
R928 B.n109 B.n108 10.6151
R929 B.n112 B.n109 10.6151
R930 B.n113 B.n112 10.6151
R931 B.n116 B.n113 10.6151
R932 B.n117 B.n116 10.6151
R933 B.n120 B.n117 10.6151
R934 B.n121 B.n120 10.6151
R935 B.n124 B.n121 10.6151
R936 B.n125 B.n124 10.6151
R937 B.n128 B.n125 10.6151
R938 B.n129 B.n128 10.6151
R939 B.n132 B.n129 10.6151
R940 B.n133 B.n132 10.6151
R941 B.n136 B.n133 10.6151
R942 B.n137 B.n136 10.6151
R943 B.n140 B.n137 10.6151
R944 B.n141 B.n140 10.6151
R945 B.n144 B.n141 10.6151
R946 B.n145 B.n144 10.6151
R947 B.n149 B.n148 10.6151
R948 B.n152 B.n149 10.6151
R949 B.n153 B.n152 10.6151
R950 B.n156 B.n153 10.6151
R951 B.n157 B.n156 10.6151
R952 B.n160 B.n157 10.6151
R953 B.n161 B.n160 10.6151
R954 B.n164 B.n161 10.6151
R955 B.n165 B.n164 10.6151
R956 B.n169 B.n168 10.6151
R957 B.n172 B.n169 10.6151
R958 B.n173 B.n172 10.6151
R959 B.n176 B.n173 10.6151
R960 B.n177 B.n176 10.6151
R961 B.n180 B.n177 10.6151
R962 B.n181 B.n180 10.6151
R963 B.n184 B.n181 10.6151
R964 B.n185 B.n184 10.6151
R965 B.n188 B.n185 10.6151
R966 B.n189 B.n188 10.6151
R967 B.n192 B.n189 10.6151
R968 B.n193 B.n192 10.6151
R969 B.n196 B.n193 10.6151
R970 B.n197 B.n196 10.6151
R971 B.n200 B.n197 10.6151
R972 B.n201 B.n200 10.6151
R973 B.n204 B.n201 10.6151
R974 B.n205 B.n204 10.6151
R975 B.n208 B.n205 10.6151
R976 B.n209 B.n208 10.6151
R977 B.n212 B.n209 10.6151
R978 B.n213 B.n212 10.6151
R979 B.n216 B.n213 10.6151
R980 B.n217 B.n216 10.6151
R981 B.n220 B.n217 10.6151
R982 B.n221 B.n220 10.6151
R983 B.n224 B.n221 10.6151
R984 B.n226 B.n224 10.6151
R985 B.n227 B.n226 10.6151
R986 B.n544 B.n227 10.6151
R987 B.n506 B.t0 9.37217
R988 B.n580 B.t1 9.37217
R989 B.n369 B.n368 9.36635
R990 B.n389 B.n283 9.36635
R991 B.n145 B.n84 9.36635
R992 B.n168 B.n81 9.36635
R993 B.n592 B.n0 8.11757
R994 B.n592 B.n1 8.11757
R995 B.n370 B.n369 1.24928
R996 B.n390 B.n389 1.24928
R997 B.n148 B.n84 1.24928
R998 B.n165 B.n81 1.24928
R999 VP.n0 VP.t1 219.511
R1000 VP.n0 VP.t0 179.499
R1001 VP VP.n0 0.241678
R1002 VTAIL.n186 VTAIL.n144 289.615
R1003 VTAIL.n42 VTAIL.n0 289.615
R1004 VTAIL.n138 VTAIL.n96 289.615
R1005 VTAIL.n90 VTAIL.n48 289.615
R1006 VTAIL.n161 VTAIL.n160 185
R1007 VTAIL.n163 VTAIL.n162 185
R1008 VTAIL.n156 VTAIL.n155 185
R1009 VTAIL.n169 VTAIL.n168 185
R1010 VTAIL.n171 VTAIL.n170 185
R1011 VTAIL.n152 VTAIL.n151 185
R1012 VTAIL.n177 VTAIL.n176 185
R1013 VTAIL.n179 VTAIL.n178 185
R1014 VTAIL.n148 VTAIL.n147 185
R1015 VTAIL.n185 VTAIL.n184 185
R1016 VTAIL.n187 VTAIL.n186 185
R1017 VTAIL.n17 VTAIL.n16 185
R1018 VTAIL.n19 VTAIL.n18 185
R1019 VTAIL.n12 VTAIL.n11 185
R1020 VTAIL.n25 VTAIL.n24 185
R1021 VTAIL.n27 VTAIL.n26 185
R1022 VTAIL.n8 VTAIL.n7 185
R1023 VTAIL.n33 VTAIL.n32 185
R1024 VTAIL.n35 VTAIL.n34 185
R1025 VTAIL.n4 VTAIL.n3 185
R1026 VTAIL.n41 VTAIL.n40 185
R1027 VTAIL.n43 VTAIL.n42 185
R1028 VTAIL.n139 VTAIL.n138 185
R1029 VTAIL.n137 VTAIL.n136 185
R1030 VTAIL.n100 VTAIL.n99 185
R1031 VTAIL.n131 VTAIL.n130 185
R1032 VTAIL.n129 VTAIL.n128 185
R1033 VTAIL.n104 VTAIL.n103 185
R1034 VTAIL.n123 VTAIL.n122 185
R1035 VTAIL.n121 VTAIL.n120 185
R1036 VTAIL.n108 VTAIL.n107 185
R1037 VTAIL.n115 VTAIL.n114 185
R1038 VTAIL.n113 VTAIL.n112 185
R1039 VTAIL.n91 VTAIL.n90 185
R1040 VTAIL.n89 VTAIL.n88 185
R1041 VTAIL.n52 VTAIL.n51 185
R1042 VTAIL.n83 VTAIL.n82 185
R1043 VTAIL.n81 VTAIL.n80 185
R1044 VTAIL.n56 VTAIL.n55 185
R1045 VTAIL.n75 VTAIL.n74 185
R1046 VTAIL.n73 VTAIL.n72 185
R1047 VTAIL.n60 VTAIL.n59 185
R1048 VTAIL.n67 VTAIL.n66 185
R1049 VTAIL.n65 VTAIL.n64 185
R1050 VTAIL.n63 VTAIL.t0 147.659
R1051 VTAIL.n159 VTAIL.t1 147.659
R1052 VTAIL.n15 VTAIL.t3 147.659
R1053 VTAIL.n111 VTAIL.t2 147.659
R1054 VTAIL.n162 VTAIL.n161 104.615
R1055 VTAIL.n162 VTAIL.n155 104.615
R1056 VTAIL.n169 VTAIL.n155 104.615
R1057 VTAIL.n170 VTAIL.n169 104.615
R1058 VTAIL.n170 VTAIL.n151 104.615
R1059 VTAIL.n177 VTAIL.n151 104.615
R1060 VTAIL.n178 VTAIL.n177 104.615
R1061 VTAIL.n178 VTAIL.n147 104.615
R1062 VTAIL.n185 VTAIL.n147 104.615
R1063 VTAIL.n186 VTAIL.n185 104.615
R1064 VTAIL.n18 VTAIL.n17 104.615
R1065 VTAIL.n18 VTAIL.n11 104.615
R1066 VTAIL.n25 VTAIL.n11 104.615
R1067 VTAIL.n26 VTAIL.n25 104.615
R1068 VTAIL.n26 VTAIL.n7 104.615
R1069 VTAIL.n33 VTAIL.n7 104.615
R1070 VTAIL.n34 VTAIL.n33 104.615
R1071 VTAIL.n34 VTAIL.n3 104.615
R1072 VTAIL.n41 VTAIL.n3 104.615
R1073 VTAIL.n42 VTAIL.n41 104.615
R1074 VTAIL.n138 VTAIL.n137 104.615
R1075 VTAIL.n137 VTAIL.n99 104.615
R1076 VTAIL.n130 VTAIL.n99 104.615
R1077 VTAIL.n130 VTAIL.n129 104.615
R1078 VTAIL.n129 VTAIL.n103 104.615
R1079 VTAIL.n122 VTAIL.n103 104.615
R1080 VTAIL.n122 VTAIL.n121 104.615
R1081 VTAIL.n121 VTAIL.n107 104.615
R1082 VTAIL.n114 VTAIL.n107 104.615
R1083 VTAIL.n114 VTAIL.n113 104.615
R1084 VTAIL.n90 VTAIL.n89 104.615
R1085 VTAIL.n89 VTAIL.n51 104.615
R1086 VTAIL.n82 VTAIL.n51 104.615
R1087 VTAIL.n82 VTAIL.n81 104.615
R1088 VTAIL.n81 VTAIL.n55 104.615
R1089 VTAIL.n74 VTAIL.n55 104.615
R1090 VTAIL.n74 VTAIL.n73 104.615
R1091 VTAIL.n73 VTAIL.n59 104.615
R1092 VTAIL.n66 VTAIL.n59 104.615
R1093 VTAIL.n66 VTAIL.n65 104.615
R1094 VTAIL.n161 VTAIL.t1 52.3082
R1095 VTAIL.n17 VTAIL.t3 52.3082
R1096 VTAIL.n113 VTAIL.t2 52.3082
R1097 VTAIL.n65 VTAIL.t0 52.3082
R1098 VTAIL.n191 VTAIL.n190 30.8278
R1099 VTAIL.n47 VTAIL.n46 30.8278
R1100 VTAIL.n143 VTAIL.n142 30.8278
R1101 VTAIL.n95 VTAIL.n94 30.8278
R1102 VTAIL.n95 VTAIL.n47 23.5652
R1103 VTAIL.n191 VTAIL.n143 21.7634
R1104 VTAIL.n160 VTAIL.n159 15.6677
R1105 VTAIL.n16 VTAIL.n15 15.6677
R1106 VTAIL.n112 VTAIL.n111 15.6677
R1107 VTAIL.n64 VTAIL.n63 15.6677
R1108 VTAIL.n163 VTAIL.n158 12.8005
R1109 VTAIL.n19 VTAIL.n14 12.8005
R1110 VTAIL.n115 VTAIL.n110 12.8005
R1111 VTAIL.n67 VTAIL.n62 12.8005
R1112 VTAIL.n164 VTAIL.n156 12.0247
R1113 VTAIL.n20 VTAIL.n12 12.0247
R1114 VTAIL.n116 VTAIL.n108 12.0247
R1115 VTAIL.n68 VTAIL.n60 12.0247
R1116 VTAIL.n168 VTAIL.n167 11.249
R1117 VTAIL.n24 VTAIL.n23 11.249
R1118 VTAIL.n120 VTAIL.n119 11.249
R1119 VTAIL.n72 VTAIL.n71 11.249
R1120 VTAIL.n171 VTAIL.n154 10.4732
R1121 VTAIL.n27 VTAIL.n10 10.4732
R1122 VTAIL.n123 VTAIL.n106 10.4732
R1123 VTAIL.n75 VTAIL.n58 10.4732
R1124 VTAIL.n172 VTAIL.n152 9.69747
R1125 VTAIL.n28 VTAIL.n8 9.69747
R1126 VTAIL.n124 VTAIL.n104 9.69747
R1127 VTAIL.n76 VTAIL.n56 9.69747
R1128 VTAIL.n190 VTAIL.n189 9.45567
R1129 VTAIL.n46 VTAIL.n45 9.45567
R1130 VTAIL.n142 VTAIL.n141 9.45567
R1131 VTAIL.n94 VTAIL.n93 9.45567
R1132 VTAIL.n183 VTAIL.n182 9.3005
R1133 VTAIL.n146 VTAIL.n145 9.3005
R1134 VTAIL.n189 VTAIL.n188 9.3005
R1135 VTAIL.n150 VTAIL.n149 9.3005
R1136 VTAIL.n175 VTAIL.n174 9.3005
R1137 VTAIL.n173 VTAIL.n172 9.3005
R1138 VTAIL.n154 VTAIL.n153 9.3005
R1139 VTAIL.n167 VTAIL.n166 9.3005
R1140 VTAIL.n165 VTAIL.n164 9.3005
R1141 VTAIL.n158 VTAIL.n157 9.3005
R1142 VTAIL.n181 VTAIL.n180 9.3005
R1143 VTAIL.n39 VTAIL.n38 9.3005
R1144 VTAIL.n2 VTAIL.n1 9.3005
R1145 VTAIL.n45 VTAIL.n44 9.3005
R1146 VTAIL.n6 VTAIL.n5 9.3005
R1147 VTAIL.n31 VTAIL.n30 9.3005
R1148 VTAIL.n29 VTAIL.n28 9.3005
R1149 VTAIL.n10 VTAIL.n9 9.3005
R1150 VTAIL.n23 VTAIL.n22 9.3005
R1151 VTAIL.n21 VTAIL.n20 9.3005
R1152 VTAIL.n14 VTAIL.n13 9.3005
R1153 VTAIL.n37 VTAIL.n36 9.3005
R1154 VTAIL.n98 VTAIL.n97 9.3005
R1155 VTAIL.n135 VTAIL.n134 9.3005
R1156 VTAIL.n133 VTAIL.n132 9.3005
R1157 VTAIL.n102 VTAIL.n101 9.3005
R1158 VTAIL.n127 VTAIL.n126 9.3005
R1159 VTAIL.n125 VTAIL.n124 9.3005
R1160 VTAIL.n106 VTAIL.n105 9.3005
R1161 VTAIL.n119 VTAIL.n118 9.3005
R1162 VTAIL.n117 VTAIL.n116 9.3005
R1163 VTAIL.n110 VTAIL.n109 9.3005
R1164 VTAIL.n141 VTAIL.n140 9.3005
R1165 VTAIL.n50 VTAIL.n49 9.3005
R1166 VTAIL.n93 VTAIL.n92 9.3005
R1167 VTAIL.n87 VTAIL.n86 9.3005
R1168 VTAIL.n85 VTAIL.n84 9.3005
R1169 VTAIL.n54 VTAIL.n53 9.3005
R1170 VTAIL.n79 VTAIL.n78 9.3005
R1171 VTAIL.n77 VTAIL.n76 9.3005
R1172 VTAIL.n58 VTAIL.n57 9.3005
R1173 VTAIL.n71 VTAIL.n70 9.3005
R1174 VTAIL.n69 VTAIL.n68 9.3005
R1175 VTAIL.n62 VTAIL.n61 9.3005
R1176 VTAIL.n176 VTAIL.n175 8.92171
R1177 VTAIL.n190 VTAIL.n144 8.92171
R1178 VTAIL.n32 VTAIL.n31 8.92171
R1179 VTAIL.n46 VTAIL.n0 8.92171
R1180 VTAIL.n142 VTAIL.n96 8.92171
R1181 VTAIL.n128 VTAIL.n127 8.92171
R1182 VTAIL.n94 VTAIL.n48 8.92171
R1183 VTAIL.n80 VTAIL.n79 8.92171
R1184 VTAIL.n179 VTAIL.n150 8.14595
R1185 VTAIL.n188 VTAIL.n187 8.14595
R1186 VTAIL.n35 VTAIL.n6 8.14595
R1187 VTAIL.n44 VTAIL.n43 8.14595
R1188 VTAIL.n140 VTAIL.n139 8.14595
R1189 VTAIL.n131 VTAIL.n102 8.14595
R1190 VTAIL.n92 VTAIL.n91 8.14595
R1191 VTAIL.n83 VTAIL.n54 8.14595
R1192 VTAIL.n180 VTAIL.n148 7.3702
R1193 VTAIL.n184 VTAIL.n146 7.3702
R1194 VTAIL.n36 VTAIL.n4 7.3702
R1195 VTAIL.n40 VTAIL.n2 7.3702
R1196 VTAIL.n136 VTAIL.n98 7.3702
R1197 VTAIL.n132 VTAIL.n100 7.3702
R1198 VTAIL.n88 VTAIL.n50 7.3702
R1199 VTAIL.n84 VTAIL.n52 7.3702
R1200 VTAIL.n183 VTAIL.n148 6.59444
R1201 VTAIL.n184 VTAIL.n183 6.59444
R1202 VTAIL.n39 VTAIL.n4 6.59444
R1203 VTAIL.n40 VTAIL.n39 6.59444
R1204 VTAIL.n136 VTAIL.n135 6.59444
R1205 VTAIL.n135 VTAIL.n100 6.59444
R1206 VTAIL.n88 VTAIL.n87 6.59444
R1207 VTAIL.n87 VTAIL.n52 6.59444
R1208 VTAIL.n180 VTAIL.n179 5.81868
R1209 VTAIL.n187 VTAIL.n146 5.81868
R1210 VTAIL.n36 VTAIL.n35 5.81868
R1211 VTAIL.n43 VTAIL.n2 5.81868
R1212 VTAIL.n139 VTAIL.n98 5.81868
R1213 VTAIL.n132 VTAIL.n131 5.81868
R1214 VTAIL.n91 VTAIL.n50 5.81868
R1215 VTAIL.n84 VTAIL.n83 5.81868
R1216 VTAIL.n176 VTAIL.n150 5.04292
R1217 VTAIL.n188 VTAIL.n144 5.04292
R1218 VTAIL.n32 VTAIL.n6 5.04292
R1219 VTAIL.n44 VTAIL.n0 5.04292
R1220 VTAIL.n140 VTAIL.n96 5.04292
R1221 VTAIL.n128 VTAIL.n102 5.04292
R1222 VTAIL.n92 VTAIL.n48 5.04292
R1223 VTAIL.n80 VTAIL.n54 5.04292
R1224 VTAIL.n159 VTAIL.n157 4.38563
R1225 VTAIL.n15 VTAIL.n13 4.38563
R1226 VTAIL.n111 VTAIL.n109 4.38563
R1227 VTAIL.n63 VTAIL.n61 4.38563
R1228 VTAIL.n175 VTAIL.n152 4.26717
R1229 VTAIL.n31 VTAIL.n8 4.26717
R1230 VTAIL.n127 VTAIL.n104 4.26717
R1231 VTAIL.n79 VTAIL.n56 4.26717
R1232 VTAIL.n172 VTAIL.n171 3.49141
R1233 VTAIL.n28 VTAIL.n27 3.49141
R1234 VTAIL.n124 VTAIL.n123 3.49141
R1235 VTAIL.n76 VTAIL.n75 3.49141
R1236 VTAIL.n168 VTAIL.n154 2.71565
R1237 VTAIL.n24 VTAIL.n10 2.71565
R1238 VTAIL.n120 VTAIL.n106 2.71565
R1239 VTAIL.n72 VTAIL.n58 2.71565
R1240 VTAIL.n167 VTAIL.n156 1.93989
R1241 VTAIL.n23 VTAIL.n12 1.93989
R1242 VTAIL.n119 VTAIL.n108 1.93989
R1243 VTAIL.n71 VTAIL.n60 1.93989
R1244 VTAIL.n143 VTAIL.n95 1.37119
R1245 VTAIL.n164 VTAIL.n163 1.16414
R1246 VTAIL.n20 VTAIL.n19 1.16414
R1247 VTAIL.n116 VTAIL.n115 1.16414
R1248 VTAIL.n68 VTAIL.n67 1.16414
R1249 VTAIL VTAIL.n47 0.978948
R1250 VTAIL VTAIL.n191 0.392741
R1251 VTAIL.n160 VTAIL.n158 0.388379
R1252 VTAIL.n16 VTAIL.n14 0.388379
R1253 VTAIL.n112 VTAIL.n110 0.388379
R1254 VTAIL.n64 VTAIL.n62 0.388379
R1255 VTAIL.n165 VTAIL.n157 0.155672
R1256 VTAIL.n166 VTAIL.n165 0.155672
R1257 VTAIL.n166 VTAIL.n153 0.155672
R1258 VTAIL.n173 VTAIL.n153 0.155672
R1259 VTAIL.n174 VTAIL.n173 0.155672
R1260 VTAIL.n174 VTAIL.n149 0.155672
R1261 VTAIL.n181 VTAIL.n149 0.155672
R1262 VTAIL.n182 VTAIL.n181 0.155672
R1263 VTAIL.n182 VTAIL.n145 0.155672
R1264 VTAIL.n189 VTAIL.n145 0.155672
R1265 VTAIL.n21 VTAIL.n13 0.155672
R1266 VTAIL.n22 VTAIL.n21 0.155672
R1267 VTAIL.n22 VTAIL.n9 0.155672
R1268 VTAIL.n29 VTAIL.n9 0.155672
R1269 VTAIL.n30 VTAIL.n29 0.155672
R1270 VTAIL.n30 VTAIL.n5 0.155672
R1271 VTAIL.n37 VTAIL.n5 0.155672
R1272 VTAIL.n38 VTAIL.n37 0.155672
R1273 VTAIL.n38 VTAIL.n1 0.155672
R1274 VTAIL.n45 VTAIL.n1 0.155672
R1275 VTAIL.n141 VTAIL.n97 0.155672
R1276 VTAIL.n134 VTAIL.n97 0.155672
R1277 VTAIL.n134 VTAIL.n133 0.155672
R1278 VTAIL.n133 VTAIL.n101 0.155672
R1279 VTAIL.n126 VTAIL.n101 0.155672
R1280 VTAIL.n126 VTAIL.n125 0.155672
R1281 VTAIL.n125 VTAIL.n105 0.155672
R1282 VTAIL.n118 VTAIL.n105 0.155672
R1283 VTAIL.n118 VTAIL.n117 0.155672
R1284 VTAIL.n117 VTAIL.n109 0.155672
R1285 VTAIL.n93 VTAIL.n49 0.155672
R1286 VTAIL.n86 VTAIL.n49 0.155672
R1287 VTAIL.n86 VTAIL.n85 0.155672
R1288 VTAIL.n85 VTAIL.n53 0.155672
R1289 VTAIL.n78 VTAIL.n53 0.155672
R1290 VTAIL.n78 VTAIL.n77 0.155672
R1291 VTAIL.n77 VTAIL.n57 0.155672
R1292 VTAIL.n70 VTAIL.n57 0.155672
R1293 VTAIL.n70 VTAIL.n69 0.155672
R1294 VTAIL.n69 VTAIL.n61 0.155672
R1295 VDD1.n42 VDD1.n0 289.615
R1296 VDD1.n89 VDD1.n47 289.615
R1297 VDD1.n43 VDD1.n42 185
R1298 VDD1.n41 VDD1.n40 185
R1299 VDD1.n4 VDD1.n3 185
R1300 VDD1.n35 VDD1.n34 185
R1301 VDD1.n33 VDD1.n32 185
R1302 VDD1.n8 VDD1.n7 185
R1303 VDD1.n27 VDD1.n26 185
R1304 VDD1.n25 VDD1.n24 185
R1305 VDD1.n12 VDD1.n11 185
R1306 VDD1.n19 VDD1.n18 185
R1307 VDD1.n17 VDD1.n16 185
R1308 VDD1.n64 VDD1.n63 185
R1309 VDD1.n66 VDD1.n65 185
R1310 VDD1.n59 VDD1.n58 185
R1311 VDD1.n72 VDD1.n71 185
R1312 VDD1.n74 VDD1.n73 185
R1313 VDD1.n55 VDD1.n54 185
R1314 VDD1.n80 VDD1.n79 185
R1315 VDD1.n82 VDD1.n81 185
R1316 VDD1.n51 VDD1.n50 185
R1317 VDD1.n88 VDD1.n87 185
R1318 VDD1.n90 VDD1.n89 185
R1319 VDD1.n15 VDD1.t0 147.659
R1320 VDD1.n62 VDD1.t1 147.659
R1321 VDD1.n42 VDD1.n41 104.615
R1322 VDD1.n41 VDD1.n3 104.615
R1323 VDD1.n34 VDD1.n3 104.615
R1324 VDD1.n34 VDD1.n33 104.615
R1325 VDD1.n33 VDD1.n7 104.615
R1326 VDD1.n26 VDD1.n7 104.615
R1327 VDD1.n26 VDD1.n25 104.615
R1328 VDD1.n25 VDD1.n11 104.615
R1329 VDD1.n18 VDD1.n11 104.615
R1330 VDD1.n18 VDD1.n17 104.615
R1331 VDD1.n65 VDD1.n64 104.615
R1332 VDD1.n65 VDD1.n58 104.615
R1333 VDD1.n72 VDD1.n58 104.615
R1334 VDD1.n73 VDD1.n72 104.615
R1335 VDD1.n73 VDD1.n54 104.615
R1336 VDD1.n80 VDD1.n54 104.615
R1337 VDD1.n81 VDD1.n80 104.615
R1338 VDD1.n81 VDD1.n50 104.615
R1339 VDD1.n88 VDD1.n50 104.615
R1340 VDD1.n89 VDD1.n88 104.615
R1341 VDD1 VDD1.n93 83.3395
R1342 VDD1.n17 VDD1.t0 52.3082
R1343 VDD1.n64 VDD1.t1 52.3082
R1344 VDD1 VDD1.n46 48.0152
R1345 VDD1.n16 VDD1.n15 15.6677
R1346 VDD1.n63 VDD1.n62 15.6677
R1347 VDD1.n19 VDD1.n14 12.8005
R1348 VDD1.n66 VDD1.n61 12.8005
R1349 VDD1.n20 VDD1.n12 12.0247
R1350 VDD1.n67 VDD1.n59 12.0247
R1351 VDD1.n24 VDD1.n23 11.249
R1352 VDD1.n71 VDD1.n70 11.249
R1353 VDD1.n27 VDD1.n10 10.4732
R1354 VDD1.n74 VDD1.n57 10.4732
R1355 VDD1.n28 VDD1.n8 9.69747
R1356 VDD1.n75 VDD1.n55 9.69747
R1357 VDD1.n46 VDD1.n45 9.45567
R1358 VDD1.n93 VDD1.n92 9.45567
R1359 VDD1.n2 VDD1.n1 9.3005
R1360 VDD1.n39 VDD1.n38 9.3005
R1361 VDD1.n37 VDD1.n36 9.3005
R1362 VDD1.n6 VDD1.n5 9.3005
R1363 VDD1.n31 VDD1.n30 9.3005
R1364 VDD1.n29 VDD1.n28 9.3005
R1365 VDD1.n10 VDD1.n9 9.3005
R1366 VDD1.n23 VDD1.n22 9.3005
R1367 VDD1.n21 VDD1.n20 9.3005
R1368 VDD1.n14 VDD1.n13 9.3005
R1369 VDD1.n45 VDD1.n44 9.3005
R1370 VDD1.n86 VDD1.n85 9.3005
R1371 VDD1.n49 VDD1.n48 9.3005
R1372 VDD1.n92 VDD1.n91 9.3005
R1373 VDD1.n53 VDD1.n52 9.3005
R1374 VDD1.n78 VDD1.n77 9.3005
R1375 VDD1.n76 VDD1.n75 9.3005
R1376 VDD1.n57 VDD1.n56 9.3005
R1377 VDD1.n70 VDD1.n69 9.3005
R1378 VDD1.n68 VDD1.n67 9.3005
R1379 VDD1.n61 VDD1.n60 9.3005
R1380 VDD1.n84 VDD1.n83 9.3005
R1381 VDD1.n46 VDD1.n0 8.92171
R1382 VDD1.n32 VDD1.n31 8.92171
R1383 VDD1.n79 VDD1.n78 8.92171
R1384 VDD1.n93 VDD1.n47 8.92171
R1385 VDD1.n44 VDD1.n43 8.14595
R1386 VDD1.n35 VDD1.n6 8.14595
R1387 VDD1.n82 VDD1.n53 8.14595
R1388 VDD1.n91 VDD1.n90 8.14595
R1389 VDD1.n40 VDD1.n2 7.3702
R1390 VDD1.n36 VDD1.n4 7.3702
R1391 VDD1.n83 VDD1.n51 7.3702
R1392 VDD1.n87 VDD1.n49 7.3702
R1393 VDD1.n40 VDD1.n39 6.59444
R1394 VDD1.n39 VDD1.n4 6.59444
R1395 VDD1.n86 VDD1.n51 6.59444
R1396 VDD1.n87 VDD1.n86 6.59444
R1397 VDD1.n43 VDD1.n2 5.81868
R1398 VDD1.n36 VDD1.n35 5.81868
R1399 VDD1.n83 VDD1.n82 5.81868
R1400 VDD1.n90 VDD1.n49 5.81868
R1401 VDD1.n44 VDD1.n0 5.04292
R1402 VDD1.n32 VDD1.n6 5.04292
R1403 VDD1.n79 VDD1.n53 5.04292
R1404 VDD1.n91 VDD1.n47 5.04292
R1405 VDD1.n15 VDD1.n13 4.38563
R1406 VDD1.n62 VDD1.n60 4.38563
R1407 VDD1.n31 VDD1.n8 4.26717
R1408 VDD1.n78 VDD1.n55 4.26717
R1409 VDD1.n28 VDD1.n27 3.49141
R1410 VDD1.n75 VDD1.n74 3.49141
R1411 VDD1.n24 VDD1.n10 2.71565
R1412 VDD1.n71 VDD1.n57 2.71565
R1413 VDD1.n23 VDD1.n12 1.93989
R1414 VDD1.n70 VDD1.n59 1.93989
R1415 VDD1.n20 VDD1.n19 1.16414
R1416 VDD1.n67 VDD1.n66 1.16414
R1417 VDD1.n16 VDD1.n14 0.388379
R1418 VDD1.n63 VDD1.n61 0.388379
R1419 VDD1.n45 VDD1.n1 0.155672
R1420 VDD1.n38 VDD1.n1 0.155672
R1421 VDD1.n38 VDD1.n37 0.155672
R1422 VDD1.n37 VDD1.n5 0.155672
R1423 VDD1.n30 VDD1.n5 0.155672
R1424 VDD1.n30 VDD1.n29 0.155672
R1425 VDD1.n29 VDD1.n9 0.155672
R1426 VDD1.n22 VDD1.n9 0.155672
R1427 VDD1.n22 VDD1.n21 0.155672
R1428 VDD1.n21 VDD1.n13 0.155672
R1429 VDD1.n68 VDD1.n60 0.155672
R1430 VDD1.n69 VDD1.n68 0.155672
R1431 VDD1.n69 VDD1.n56 0.155672
R1432 VDD1.n76 VDD1.n56 0.155672
R1433 VDD1.n77 VDD1.n76 0.155672
R1434 VDD1.n77 VDD1.n52 0.155672
R1435 VDD1.n84 VDD1.n52 0.155672
R1436 VDD1.n85 VDD1.n84 0.155672
R1437 VDD1.n85 VDD1.n48 0.155672
R1438 VDD1.n92 VDD1.n48 0.155672
R1439 VN VN.t0 219.702
R1440 VN VN.t1 179.739
R1441 VDD2.n89 VDD2.n47 289.615
R1442 VDD2.n42 VDD2.n0 289.615
R1443 VDD2.n90 VDD2.n89 185
R1444 VDD2.n88 VDD2.n87 185
R1445 VDD2.n51 VDD2.n50 185
R1446 VDD2.n82 VDD2.n81 185
R1447 VDD2.n80 VDD2.n79 185
R1448 VDD2.n55 VDD2.n54 185
R1449 VDD2.n74 VDD2.n73 185
R1450 VDD2.n72 VDD2.n71 185
R1451 VDD2.n59 VDD2.n58 185
R1452 VDD2.n66 VDD2.n65 185
R1453 VDD2.n64 VDD2.n63 185
R1454 VDD2.n17 VDD2.n16 185
R1455 VDD2.n19 VDD2.n18 185
R1456 VDD2.n12 VDD2.n11 185
R1457 VDD2.n25 VDD2.n24 185
R1458 VDD2.n27 VDD2.n26 185
R1459 VDD2.n8 VDD2.n7 185
R1460 VDD2.n33 VDD2.n32 185
R1461 VDD2.n35 VDD2.n34 185
R1462 VDD2.n4 VDD2.n3 185
R1463 VDD2.n41 VDD2.n40 185
R1464 VDD2.n43 VDD2.n42 185
R1465 VDD2.n62 VDD2.t1 147.659
R1466 VDD2.n15 VDD2.t0 147.659
R1467 VDD2.n89 VDD2.n88 104.615
R1468 VDD2.n88 VDD2.n50 104.615
R1469 VDD2.n81 VDD2.n50 104.615
R1470 VDD2.n81 VDD2.n80 104.615
R1471 VDD2.n80 VDD2.n54 104.615
R1472 VDD2.n73 VDD2.n54 104.615
R1473 VDD2.n73 VDD2.n72 104.615
R1474 VDD2.n72 VDD2.n58 104.615
R1475 VDD2.n65 VDD2.n58 104.615
R1476 VDD2.n65 VDD2.n64 104.615
R1477 VDD2.n18 VDD2.n17 104.615
R1478 VDD2.n18 VDD2.n11 104.615
R1479 VDD2.n25 VDD2.n11 104.615
R1480 VDD2.n26 VDD2.n25 104.615
R1481 VDD2.n26 VDD2.n7 104.615
R1482 VDD2.n33 VDD2.n7 104.615
R1483 VDD2.n34 VDD2.n33 104.615
R1484 VDD2.n34 VDD2.n3 104.615
R1485 VDD2.n41 VDD2.n3 104.615
R1486 VDD2.n42 VDD2.n41 104.615
R1487 VDD2.n94 VDD2.n46 82.3643
R1488 VDD2.n64 VDD2.t1 52.3082
R1489 VDD2.n17 VDD2.t0 52.3082
R1490 VDD2.n94 VDD2.n93 47.5066
R1491 VDD2.n63 VDD2.n62 15.6677
R1492 VDD2.n16 VDD2.n15 15.6677
R1493 VDD2.n66 VDD2.n61 12.8005
R1494 VDD2.n19 VDD2.n14 12.8005
R1495 VDD2.n67 VDD2.n59 12.0247
R1496 VDD2.n20 VDD2.n12 12.0247
R1497 VDD2.n71 VDD2.n70 11.249
R1498 VDD2.n24 VDD2.n23 11.249
R1499 VDD2.n74 VDD2.n57 10.4732
R1500 VDD2.n27 VDD2.n10 10.4732
R1501 VDD2.n75 VDD2.n55 9.69747
R1502 VDD2.n28 VDD2.n8 9.69747
R1503 VDD2.n93 VDD2.n92 9.45567
R1504 VDD2.n46 VDD2.n45 9.45567
R1505 VDD2.n49 VDD2.n48 9.3005
R1506 VDD2.n86 VDD2.n85 9.3005
R1507 VDD2.n84 VDD2.n83 9.3005
R1508 VDD2.n53 VDD2.n52 9.3005
R1509 VDD2.n78 VDD2.n77 9.3005
R1510 VDD2.n76 VDD2.n75 9.3005
R1511 VDD2.n57 VDD2.n56 9.3005
R1512 VDD2.n70 VDD2.n69 9.3005
R1513 VDD2.n68 VDD2.n67 9.3005
R1514 VDD2.n61 VDD2.n60 9.3005
R1515 VDD2.n92 VDD2.n91 9.3005
R1516 VDD2.n39 VDD2.n38 9.3005
R1517 VDD2.n2 VDD2.n1 9.3005
R1518 VDD2.n45 VDD2.n44 9.3005
R1519 VDD2.n6 VDD2.n5 9.3005
R1520 VDD2.n31 VDD2.n30 9.3005
R1521 VDD2.n29 VDD2.n28 9.3005
R1522 VDD2.n10 VDD2.n9 9.3005
R1523 VDD2.n23 VDD2.n22 9.3005
R1524 VDD2.n21 VDD2.n20 9.3005
R1525 VDD2.n14 VDD2.n13 9.3005
R1526 VDD2.n37 VDD2.n36 9.3005
R1527 VDD2.n93 VDD2.n47 8.92171
R1528 VDD2.n79 VDD2.n78 8.92171
R1529 VDD2.n32 VDD2.n31 8.92171
R1530 VDD2.n46 VDD2.n0 8.92171
R1531 VDD2.n91 VDD2.n90 8.14595
R1532 VDD2.n82 VDD2.n53 8.14595
R1533 VDD2.n35 VDD2.n6 8.14595
R1534 VDD2.n44 VDD2.n43 8.14595
R1535 VDD2.n87 VDD2.n49 7.3702
R1536 VDD2.n83 VDD2.n51 7.3702
R1537 VDD2.n36 VDD2.n4 7.3702
R1538 VDD2.n40 VDD2.n2 7.3702
R1539 VDD2.n87 VDD2.n86 6.59444
R1540 VDD2.n86 VDD2.n51 6.59444
R1541 VDD2.n39 VDD2.n4 6.59444
R1542 VDD2.n40 VDD2.n39 6.59444
R1543 VDD2.n90 VDD2.n49 5.81868
R1544 VDD2.n83 VDD2.n82 5.81868
R1545 VDD2.n36 VDD2.n35 5.81868
R1546 VDD2.n43 VDD2.n2 5.81868
R1547 VDD2.n91 VDD2.n47 5.04292
R1548 VDD2.n79 VDD2.n53 5.04292
R1549 VDD2.n32 VDD2.n6 5.04292
R1550 VDD2.n44 VDD2.n0 5.04292
R1551 VDD2.n62 VDD2.n60 4.38563
R1552 VDD2.n15 VDD2.n13 4.38563
R1553 VDD2.n78 VDD2.n55 4.26717
R1554 VDD2.n31 VDD2.n8 4.26717
R1555 VDD2.n75 VDD2.n74 3.49141
R1556 VDD2.n28 VDD2.n27 3.49141
R1557 VDD2.n71 VDD2.n57 2.71565
R1558 VDD2.n24 VDD2.n10 2.71565
R1559 VDD2.n70 VDD2.n59 1.93989
R1560 VDD2.n23 VDD2.n12 1.93989
R1561 VDD2.n67 VDD2.n66 1.16414
R1562 VDD2.n20 VDD2.n19 1.16414
R1563 VDD2 VDD2.n94 0.509121
R1564 VDD2.n63 VDD2.n61 0.388379
R1565 VDD2.n16 VDD2.n14 0.388379
R1566 VDD2.n92 VDD2.n48 0.155672
R1567 VDD2.n85 VDD2.n48 0.155672
R1568 VDD2.n85 VDD2.n84 0.155672
R1569 VDD2.n84 VDD2.n52 0.155672
R1570 VDD2.n77 VDD2.n52 0.155672
R1571 VDD2.n77 VDD2.n76 0.155672
R1572 VDD2.n76 VDD2.n56 0.155672
R1573 VDD2.n69 VDD2.n56 0.155672
R1574 VDD2.n69 VDD2.n68 0.155672
R1575 VDD2.n68 VDD2.n60 0.155672
R1576 VDD2.n21 VDD2.n13 0.155672
R1577 VDD2.n22 VDD2.n21 0.155672
R1578 VDD2.n22 VDD2.n9 0.155672
R1579 VDD2.n29 VDD2.n9 0.155672
R1580 VDD2.n30 VDD2.n29 0.155672
R1581 VDD2.n30 VDD2.n5 0.155672
R1582 VDD2.n37 VDD2.n5 0.155672
R1583 VDD2.n38 VDD2.n37 0.155672
R1584 VDD2.n38 VDD2.n1 0.155672
R1585 VDD2.n45 VDD2.n1 0.155672
C0 VDD1 VTAIL 4.11558f
C1 VN VP 4.47236f
C2 VDD2 VP 0.297531f
C3 VP VDD1 2.11318f
C4 VN VDD2 1.96574f
C5 VP VTAIL 1.72612f
C6 VN VDD1 0.147737f
C7 VDD2 VDD1 0.575098f
C8 VN VTAIL 1.71181f
C9 VDD2 VTAIL 4.16043f
C10 VDD2 B 3.533416f
C11 VDD1 B 5.86027f
C12 VTAIL B 5.653795f
C13 VN B 7.372149f
C14 VP B 5.134114f
C15 VDD2.n0 B 0.020536f
C16 VDD2.n1 B 0.014005f
C17 VDD2.n2 B 0.007526f
C18 VDD2.n3 B 0.017788f
C19 VDD2.n4 B 0.007968f
C20 VDD2.n5 B 0.014005f
C21 VDD2.n6 B 0.007526f
C22 VDD2.n7 B 0.017788f
C23 VDD2.n8 B 0.007968f
C24 VDD2.n9 B 0.014005f
C25 VDD2.n10 B 0.007526f
C26 VDD2.n11 B 0.017788f
C27 VDD2.n12 B 0.007968f
C28 VDD2.n13 B 0.513866f
C29 VDD2.n14 B 0.007526f
C30 VDD2.t0 B 0.02904f
C31 VDD2.n15 B 0.069623f
C32 VDD2.n16 B 0.010508f
C33 VDD2.n17 B 0.013341f
C34 VDD2.n18 B 0.017788f
C35 VDD2.n19 B 0.007968f
C36 VDD2.n20 B 0.007526f
C37 VDD2.n21 B 0.014005f
C38 VDD2.n22 B 0.014005f
C39 VDD2.n23 B 0.007526f
C40 VDD2.n24 B 0.007968f
C41 VDD2.n25 B 0.017788f
C42 VDD2.n26 B 0.017788f
C43 VDD2.n27 B 0.007968f
C44 VDD2.n28 B 0.007526f
C45 VDD2.n29 B 0.014005f
C46 VDD2.n30 B 0.014005f
C47 VDD2.n31 B 0.007526f
C48 VDD2.n32 B 0.007968f
C49 VDD2.n33 B 0.017788f
C50 VDD2.n34 B 0.017788f
C51 VDD2.n35 B 0.007968f
C52 VDD2.n36 B 0.007526f
C53 VDD2.n37 B 0.014005f
C54 VDD2.n38 B 0.014005f
C55 VDD2.n39 B 0.007526f
C56 VDD2.n40 B 0.007968f
C57 VDD2.n41 B 0.017788f
C58 VDD2.n42 B 0.040012f
C59 VDD2.n43 B 0.007968f
C60 VDD2.n44 B 0.007526f
C61 VDD2.n45 B 0.031033f
C62 VDD2.n46 B 0.326993f
C63 VDD2.n47 B 0.020536f
C64 VDD2.n48 B 0.014005f
C65 VDD2.n49 B 0.007526f
C66 VDD2.n50 B 0.017788f
C67 VDD2.n51 B 0.007968f
C68 VDD2.n52 B 0.014005f
C69 VDD2.n53 B 0.007526f
C70 VDD2.n54 B 0.017788f
C71 VDD2.n55 B 0.007968f
C72 VDD2.n56 B 0.014005f
C73 VDD2.n57 B 0.007526f
C74 VDD2.n58 B 0.017788f
C75 VDD2.n59 B 0.007968f
C76 VDD2.n60 B 0.513866f
C77 VDD2.n61 B 0.007526f
C78 VDD2.t1 B 0.02904f
C79 VDD2.n62 B 0.069623f
C80 VDD2.n63 B 0.010508f
C81 VDD2.n64 B 0.013341f
C82 VDD2.n65 B 0.017788f
C83 VDD2.n66 B 0.007968f
C84 VDD2.n67 B 0.007526f
C85 VDD2.n68 B 0.014005f
C86 VDD2.n69 B 0.014005f
C87 VDD2.n70 B 0.007526f
C88 VDD2.n71 B 0.007968f
C89 VDD2.n72 B 0.017788f
C90 VDD2.n73 B 0.017788f
C91 VDD2.n74 B 0.007968f
C92 VDD2.n75 B 0.007526f
C93 VDD2.n76 B 0.014005f
C94 VDD2.n77 B 0.014005f
C95 VDD2.n78 B 0.007526f
C96 VDD2.n79 B 0.007968f
C97 VDD2.n80 B 0.017788f
C98 VDD2.n81 B 0.017788f
C99 VDD2.n82 B 0.007968f
C100 VDD2.n83 B 0.007526f
C101 VDD2.n84 B 0.014005f
C102 VDD2.n85 B 0.014005f
C103 VDD2.n86 B 0.007526f
C104 VDD2.n87 B 0.007968f
C105 VDD2.n88 B 0.017788f
C106 VDD2.n89 B 0.040012f
C107 VDD2.n90 B 0.007968f
C108 VDD2.n91 B 0.007526f
C109 VDD2.n92 B 0.031033f
C110 VDD2.n93 B 0.032183f
C111 VDD2.n94 B 1.42369f
C112 VN.t1 B 1.05433f
C113 VN.t0 B 1.27003f
C114 VDD1.n0 B 0.029946f
C115 VDD1.n1 B 0.020423f
C116 VDD1.n2 B 0.010974f
C117 VDD1.n3 B 0.025939f
C118 VDD1.n4 B 0.01162f
C119 VDD1.n5 B 0.020423f
C120 VDD1.n6 B 0.010974f
C121 VDD1.n7 B 0.025939f
C122 VDD1.n8 B 0.01162f
C123 VDD1.n9 B 0.020423f
C124 VDD1.n10 B 0.010974f
C125 VDD1.n11 B 0.025939f
C126 VDD1.n12 B 0.01162f
C127 VDD1.n13 B 0.749336f
C128 VDD1.n14 B 0.010974f
C129 VDD1.t0 B 0.042347f
C130 VDD1.n15 B 0.101526f
C131 VDD1.n16 B 0.015323f
C132 VDD1.n17 B 0.019454f
C133 VDD1.n18 B 0.025939f
C134 VDD1.n19 B 0.01162f
C135 VDD1.n20 B 0.010974f
C136 VDD1.n21 B 0.020423f
C137 VDD1.n22 B 0.020423f
C138 VDD1.n23 B 0.010974f
C139 VDD1.n24 B 0.01162f
C140 VDD1.n25 B 0.025939f
C141 VDD1.n26 B 0.025939f
C142 VDD1.n27 B 0.01162f
C143 VDD1.n28 B 0.010974f
C144 VDD1.n29 B 0.020423f
C145 VDD1.n30 B 0.020423f
C146 VDD1.n31 B 0.010974f
C147 VDD1.n32 B 0.01162f
C148 VDD1.n33 B 0.025939f
C149 VDD1.n34 B 0.025939f
C150 VDD1.n35 B 0.01162f
C151 VDD1.n36 B 0.010974f
C152 VDD1.n37 B 0.020423f
C153 VDD1.n38 B 0.020423f
C154 VDD1.n39 B 0.010974f
C155 VDD1.n40 B 0.01162f
C156 VDD1.n41 B 0.025939f
C157 VDD1.n42 B 0.058347f
C158 VDD1.n43 B 0.01162f
C159 VDD1.n44 B 0.010974f
C160 VDD1.n45 B 0.045253f
C161 VDD1.n46 B 0.047689f
C162 VDD1.n47 B 0.029946f
C163 VDD1.n48 B 0.020423f
C164 VDD1.n49 B 0.010974f
C165 VDD1.n50 B 0.025939f
C166 VDD1.n51 B 0.01162f
C167 VDD1.n52 B 0.020423f
C168 VDD1.n53 B 0.010974f
C169 VDD1.n54 B 0.025939f
C170 VDD1.n55 B 0.01162f
C171 VDD1.n56 B 0.020423f
C172 VDD1.n57 B 0.010974f
C173 VDD1.n58 B 0.025939f
C174 VDD1.n59 B 0.01162f
C175 VDD1.n60 B 0.749336f
C176 VDD1.n61 B 0.010974f
C177 VDD1.t1 B 0.042347f
C178 VDD1.n62 B 0.101526f
C179 VDD1.n63 B 0.015323f
C180 VDD1.n64 B 0.019454f
C181 VDD1.n65 B 0.025939f
C182 VDD1.n66 B 0.01162f
C183 VDD1.n67 B 0.010974f
C184 VDD1.n68 B 0.020423f
C185 VDD1.n69 B 0.020423f
C186 VDD1.n70 B 0.010974f
C187 VDD1.n71 B 0.01162f
C188 VDD1.n72 B 0.025939f
C189 VDD1.n73 B 0.025939f
C190 VDD1.n74 B 0.01162f
C191 VDD1.n75 B 0.010974f
C192 VDD1.n76 B 0.020423f
C193 VDD1.n77 B 0.020423f
C194 VDD1.n78 B 0.010974f
C195 VDD1.n79 B 0.01162f
C196 VDD1.n80 B 0.025939f
C197 VDD1.n81 B 0.025939f
C198 VDD1.n82 B 0.01162f
C199 VDD1.n83 B 0.010974f
C200 VDD1.n84 B 0.020423f
C201 VDD1.n85 B 0.020423f
C202 VDD1.n86 B 0.010974f
C203 VDD1.n87 B 0.01162f
C204 VDD1.n88 B 0.025939f
C205 VDD1.n89 B 0.058347f
C206 VDD1.n90 B 0.01162f
C207 VDD1.n91 B 0.010974f
C208 VDD1.n92 B 0.045253f
C209 VDD1.n93 B 0.50944f
C210 VTAIL.n0 B 0.022112f
C211 VTAIL.n1 B 0.01508f
C212 VTAIL.n2 B 0.008103f
C213 VTAIL.n3 B 0.019154f
C214 VTAIL.n4 B 0.00858f
C215 VTAIL.n5 B 0.01508f
C216 VTAIL.n6 B 0.008103f
C217 VTAIL.n7 B 0.019154f
C218 VTAIL.n8 B 0.00858f
C219 VTAIL.n9 B 0.01508f
C220 VTAIL.n10 B 0.008103f
C221 VTAIL.n11 B 0.019154f
C222 VTAIL.n12 B 0.00858f
C223 VTAIL.n13 B 0.553311f
C224 VTAIL.n14 B 0.008103f
C225 VTAIL.t3 B 0.031269f
C226 VTAIL.n15 B 0.074967f
C227 VTAIL.n16 B 0.011315f
C228 VTAIL.n17 B 0.014365f
C229 VTAIL.n18 B 0.019154f
C230 VTAIL.n19 B 0.00858f
C231 VTAIL.n20 B 0.008103f
C232 VTAIL.n21 B 0.01508f
C233 VTAIL.n22 B 0.01508f
C234 VTAIL.n23 B 0.008103f
C235 VTAIL.n24 B 0.00858f
C236 VTAIL.n25 B 0.019154f
C237 VTAIL.n26 B 0.019154f
C238 VTAIL.n27 B 0.00858f
C239 VTAIL.n28 B 0.008103f
C240 VTAIL.n29 B 0.01508f
C241 VTAIL.n30 B 0.01508f
C242 VTAIL.n31 B 0.008103f
C243 VTAIL.n32 B 0.00858f
C244 VTAIL.n33 B 0.019154f
C245 VTAIL.n34 B 0.019154f
C246 VTAIL.n35 B 0.00858f
C247 VTAIL.n36 B 0.008103f
C248 VTAIL.n37 B 0.01508f
C249 VTAIL.n38 B 0.01508f
C250 VTAIL.n39 B 0.008103f
C251 VTAIL.n40 B 0.00858f
C252 VTAIL.n41 B 0.019154f
C253 VTAIL.n42 B 0.043084f
C254 VTAIL.n43 B 0.00858f
C255 VTAIL.n44 B 0.008103f
C256 VTAIL.n45 B 0.033415f
C257 VTAIL.n46 B 0.024228f
C258 VTAIL.n47 B 0.808604f
C259 VTAIL.n48 B 0.022112f
C260 VTAIL.n49 B 0.01508f
C261 VTAIL.n50 B 0.008103f
C262 VTAIL.n51 B 0.019154f
C263 VTAIL.n52 B 0.00858f
C264 VTAIL.n53 B 0.01508f
C265 VTAIL.n54 B 0.008103f
C266 VTAIL.n55 B 0.019154f
C267 VTAIL.n56 B 0.00858f
C268 VTAIL.n57 B 0.01508f
C269 VTAIL.n58 B 0.008103f
C270 VTAIL.n59 B 0.019154f
C271 VTAIL.n60 B 0.00858f
C272 VTAIL.n61 B 0.553311f
C273 VTAIL.n62 B 0.008103f
C274 VTAIL.t0 B 0.031269f
C275 VTAIL.n63 B 0.074967f
C276 VTAIL.n64 B 0.011315f
C277 VTAIL.n65 B 0.014365f
C278 VTAIL.n66 B 0.019154f
C279 VTAIL.n67 B 0.00858f
C280 VTAIL.n68 B 0.008103f
C281 VTAIL.n69 B 0.01508f
C282 VTAIL.n70 B 0.01508f
C283 VTAIL.n71 B 0.008103f
C284 VTAIL.n72 B 0.00858f
C285 VTAIL.n73 B 0.019154f
C286 VTAIL.n74 B 0.019154f
C287 VTAIL.n75 B 0.00858f
C288 VTAIL.n76 B 0.008103f
C289 VTAIL.n77 B 0.01508f
C290 VTAIL.n78 B 0.01508f
C291 VTAIL.n79 B 0.008103f
C292 VTAIL.n80 B 0.00858f
C293 VTAIL.n81 B 0.019154f
C294 VTAIL.n82 B 0.019154f
C295 VTAIL.n83 B 0.00858f
C296 VTAIL.n84 B 0.008103f
C297 VTAIL.n85 B 0.01508f
C298 VTAIL.n86 B 0.01508f
C299 VTAIL.n87 B 0.008103f
C300 VTAIL.n88 B 0.00858f
C301 VTAIL.n89 B 0.019154f
C302 VTAIL.n90 B 0.043084f
C303 VTAIL.n91 B 0.00858f
C304 VTAIL.n92 B 0.008103f
C305 VTAIL.n93 B 0.033415f
C306 VTAIL.n94 B 0.024228f
C307 VTAIL.n95 B 0.827664f
C308 VTAIL.n96 B 0.022112f
C309 VTAIL.n97 B 0.01508f
C310 VTAIL.n98 B 0.008103f
C311 VTAIL.n99 B 0.019154f
C312 VTAIL.n100 B 0.00858f
C313 VTAIL.n101 B 0.01508f
C314 VTAIL.n102 B 0.008103f
C315 VTAIL.n103 B 0.019154f
C316 VTAIL.n104 B 0.00858f
C317 VTAIL.n105 B 0.01508f
C318 VTAIL.n106 B 0.008103f
C319 VTAIL.n107 B 0.019154f
C320 VTAIL.n108 B 0.00858f
C321 VTAIL.n109 B 0.553311f
C322 VTAIL.n110 B 0.008103f
C323 VTAIL.t2 B 0.031269f
C324 VTAIL.n111 B 0.074967f
C325 VTAIL.n112 B 0.011315f
C326 VTAIL.n113 B 0.014365f
C327 VTAIL.n114 B 0.019154f
C328 VTAIL.n115 B 0.00858f
C329 VTAIL.n116 B 0.008103f
C330 VTAIL.n117 B 0.01508f
C331 VTAIL.n118 B 0.01508f
C332 VTAIL.n119 B 0.008103f
C333 VTAIL.n120 B 0.00858f
C334 VTAIL.n121 B 0.019154f
C335 VTAIL.n122 B 0.019154f
C336 VTAIL.n123 B 0.00858f
C337 VTAIL.n124 B 0.008103f
C338 VTAIL.n125 B 0.01508f
C339 VTAIL.n126 B 0.01508f
C340 VTAIL.n127 B 0.008103f
C341 VTAIL.n128 B 0.00858f
C342 VTAIL.n129 B 0.019154f
C343 VTAIL.n130 B 0.019154f
C344 VTAIL.n131 B 0.00858f
C345 VTAIL.n132 B 0.008103f
C346 VTAIL.n133 B 0.01508f
C347 VTAIL.n134 B 0.01508f
C348 VTAIL.n135 B 0.008103f
C349 VTAIL.n136 B 0.00858f
C350 VTAIL.n137 B 0.019154f
C351 VTAIL.n138 B 0.043084f
C352 VTAIL.n139 B 0.00858f
C353 VTAIL.n140 B 0.008103f
C354 VTAIL.n141 B 0.033415f
C355 VTAIL.n142 B 0.024228f
C356 VTAIL.n143 B 0.740114f
C357 VTAIL.n144 B 0.022112f
C358 VTAIL.n145 B 0.01508f
C359 VTAIL.n146 B 0.008103f
C360 VTAIL.n147 B 0.019154f
C361 VTAIL.n148 B 0.00858f
C362 VTAIL.n149 B 0.01508f
C363 VTAIL.n150 B 0.008103f
C364 VTAIL.n151 B 0.019154f
C365 VTAIL.n152 B 0.00858f
C366 VTAIL.n153 B 0.01508f
C367 VTAIL.n154 B 0.008103f
C368 VTAIL.n155 B 0.019154f
C369 VTAIL.n156 B 0.00858f
C370 VTAIL.n157 B 0.553311f
C371 VTAIL.n158 B 0.008103f
C372 VTAIL.t1 B 0.031269f
C373 VTAIL.n159 B 0.074967f
C374 VTAIL.n160 B 0.011315f
C375 VTAIL.n161 B 0.014365f
C376 VTAIL.n162 B 0.019154f
C377 VTAIL.n163 B 0.00858f
C378 VTAIL.n164 B 0.008103f
C379 VTAIL.n165 B 0.01508f
C380 VTAIL.n166 B 0.01508f
C381 VTAIL.n167 B 0.008103f
C382 VTAIL.n168 B 0.00858f
C383 VTAIL.n169 B 0.019154f
C384 VTAIL.n170 B 0.019154f
C385 VTAIL.n171 B 0.00858f
C386 VTAIL.n172 B 0.008103f
C387 VTAIL.n173 B 0.01508f
C388 VTAIL.n174 B 0.01508f
C389 VTAIL.n175 B 0.008103f
C390 VTAIL.n176 B 0.00858f
C391 VTAIL.n177 B 0.019154f
C392 VTAIL.n178 B 0.019154f
C393 VTAIL.n179 B 0.00858f
C394 VTAIL.n180 B 0.008103f
C395 VTAIL.n181 B 0.01508f
C396 VTAIL.n182 B 0.01508f
C397 VTAIL.n183 B 0.008103f
C398 VTAIL.n184 B 0.00858f
C399 VTAIL.n185 B 0.019154f
C400 VTAIL.n186 B 0.043084f
C401 VTAIL.n187 B 0.00858f
C402 VTAIL.n188 B 0.008103f
C403 VTAIL.n189 B 0.033415f
C404 VTAIL.n190 B 0.024228f
C405 VTAIL.n191 B 0.69257f
C406 VP.t1 B 1.87145f
C407 VP.t0 B 1.55622f
C408 VP.n0 B 3.12453f
.ends

