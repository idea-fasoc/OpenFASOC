* NGSPICE file created from diff_pair_sample_0246.ext - technology: sky130A

.subckt diff_pair_sample_0246 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2550_n2140# sky130_fd_pr__pfet_01v8 ad=2.2854 pd=12.5 as=0 ps=0 w=5.86 l=3.62
X1 B.t8 B.t6 B.t7 w_n2550_n2140# sky130_fd_pr__pfet_01v8 ad=2.2854 pd=12.5 as=0 ps=0 w=5.86 l=3.62
X2 VDD1.t1 VP.t0 VTAIL.t2 w_n2550_n2140# sky130_fd_pr__pfet_01v8 ad=2.2854 pd=12.5 as=2.2854 ps=12.5 w=5.86 l=3.62
X3 VDD2.t1 VN.t0 VTAIL.t0 w_n2550_n2140# sky130_fd_pr__pfet_01v8 ad=2.2854 pd=12.5 as=2.2854 ps=12.5 w=5.86 l=3.62
X4 B.t5 B.t3 B.t4 w_n2550_n2140# sky130_fd_pr__pfet_01v8 ad=2.2854 pd=12.5 as=0 ps=0 w=5.86 l=3.62
X5 VDD2.t0 VN.t1 VTAIL.t1 w_n2550_n2140# sky130_fd_pr__pfet_01v8 ad=2.2854 pd=12.5 as=2.2854 ps=12.5 w=5.86 l=3.62
X6 B.t2 B.t0 B.t1 w_n2550_n2140# sky130_fd_pr__pfet_01v8 ad=2.2854 pd=12.5 as=0 ps=0 w=5.86 l=3.62
X7 VDD1.t0 VP.t1 VTAIL.t3 w_n2550_n2140# sky130_fd_pr__pfet_01v8 ad=2.2854 pd=12.5 as=2.2854 ps=12.5 w=5.86 l=3.62
R0 B.n262 B.n261 585
R1 B.n260 B.n83 585
R2 B.n259 B.n258 585
R3 B.n257 B.n84 585
R4 B.n256 B.n255 585
R5 B.n254 B.n85 585
R6 B.n253 B.n252 585
R7 B.n251 B.n86 585
R8 B.n250 B.n249 585
R9 B.n248 B.n87 585
R10 B.n247 B.n246 585
R11 B.n245 B.n88 585
R12 B.n244 B.n243 585
R13 B.n242 B.n89 585
R14 B.n241 B.n240 585
R15 B.n239 B.n90 585
R16 B.n238 B.n237 585
R17 B.n236 B.n91 585
R18 B.n235 B.n234 585
R19 B.n233 B.n92 585
R20 B.n232 B.n231 585
R21 B.n230 B.n93 585
R22 B.n229 B.n228 585
R23 B.n227 B.n94 585
R24 B.n226 B.n225 585
R25 B.n221 B.n95 585
R26 B.n220 B.n219 585
R27 B.n218 B.n96 585
R28 B.n217 B.n216 585
R29 B.n215 B.n97 585
R30 B.n214 B.n213 585
R31 B.n212 B.n98 585
R32 B.n211 B.n210 585
R33 B.n208 B.n99 585
R34 B.n207 B.n206 585
R35 B.n205 B.n102 585
R36 B.n204 B.n203 585
R37 B.n202 B.n103 585
R38 B.n201 B.n200 585
R39 B.n199 B.n104 585
R40 B.n198 B.n197 585
R41 B.n196 B.n105 585
R42 B.n195 B.n194 585
R43 B.n193 B.n106 585
R44 B.n192 B.n191 585
R45 B.n190 B.n107 585
R46 B.n189 B.n188 585
R47 B.n187 B.n108 585
R48 B.n186 B.n185 585
R49 B.n184 B.n109 585
R50 B.n183 B.n182 585
R51 B.n181 B.n110 585
R52 B.n180 B.n179 585
R53 B.n178 B.n111 585
R54 B.n177 B.n176 585
R55 B.n175 B.n112 585
R56 B.n174 B.n173 585
R57 B.n263 B.n82 585
R58 B.n265 B.n264 585
R59 B.n266 B.n81 585
R60 B.n268 B.n267 585
R61 B.n269 B.n80 585
R62 B.n271 B.n270 585
R63 B.n272 B.n79 585
R64 B.n274 B.n273 585
R65 B.n275 B.n78 585
R66 B.n277 B.n276 585
R67 B.n278 B.n77 585
R68 B.n280 B.n279 585
R69 B.n281 B.n76 585
R70 B.n283 B.n282 585
R71 B.n284 B.n75 585
R72 B.n286 B.n285 585
R73 B.n287 B.n74 585
R74 B.n289 B.n288 585
R75 B.n290 B.n73 585
R76 B.n292 B.n291 585
R77 B.n293 B.n72 585
R78 B.n295 B.n294 585
R79 B.n296 B.n71 585
R80 B.n298 B.n297 585
R81 B.n299 B.n70 585
R82 B.n301 B.n300 585
R83 B.n302 B.n69 585
R84 B.n304 B.n303 585
R85 B.n305 B.n68 585
R86 B.n307 B.n306 585
R87 B.n308 B.n67 585
R88 B.n310 B.n309 585
R89 B.n311 B.n66 585
R90 B.n313 B.n312 585
R91 B.n314 B.n65 585
R92 B.n316 B.n315 585
R93 B.n317 B.n64 585
R94 B.n319 B.n318 585
R95 B.n320 B.n63 585
R96 B.n322 B.n321 585
R97 B.n323 B.n62 585
R98 B.n325 B.n324 585
R99 B.n326 B.n61 585
R100 B.n328 B.n327 585
R101 B.n329 B.n60 585
R102 B.n331 B.n330 585
R103 B.n332 B.n59 585
R104 B.n334 B.n333 585
R105 B.n335 B.n58 585
R106 B.n337 B.n336 585
R107 B.n338 B.n57 585
R108 B.n340 B.n339 585
R109 B.n341 B.n56 585
R110 B.n343 B.n342 585
R111 B.n344 B.n55 585
R112 B.n346 B.n345 585
R113 B.n347 B.n54 585
R114 B.n349 B.n348 585
R115 B.n350 B.n53 585
R116 B.n352 B.n351 585
R117 B.n353 B.n52 585
R118 B.n355 B.n354 585
R119 B.n356 B.n51 585
R120 B.n358 B.n357 585
R121 B.n445 B.n444 585
R122 B.n443 B.n18 585
R123 B.n442 B.n441 585
R124 B.n440 B.n19 585
R125 B.n439 B.n438 585
R126 B.n437 B.n20 585
R127 B.n436 B.n435 585
R128 B.n434 B.n21 585
R129 B.n433 B.n432 585
R130 B.n431 B.n22 585
R131 B.n430 B.n429 585
R132 B.n428 B.n23 585
R133 B.n427 B.n426 585
R134 B.n425 B.n24 585
R135 B.n424 B.n423 585
R136 B.n422 B.n25 585
R137 B.n421 B.n420 585
R138 B.n419 B.n26 585
R139 B.n418 B.n417 585
R140 B.n416 B.n27 585
R141 B.n415 B.n414 585
R142 B.n413 B.n28 585
R143 B.n412 B.n411 585
R144 B.n410 B.n29 585
R145 B.n408 B.n407 585
R146 B.n406 B.n32 585
R147 B.n405 B.n404 585
R148 B.n403 B.n33 585
R149 B.n402 B.n401 585
R150 B.n400 B.n34 585
R151 B.n399 B.n398 585
R152 B.n397 B.n35 585
R153 B.n396 B.n395 585
R154 B.n394 B.n393 585
R155 B.n392 B.n39 585
R156 B.n391 B.n390 585
R157 B.n389 B.n40 585
R158 B.n388 B.n387 585
R159 B.n386 B.n41 585
R160 B.n385 B.n384 585
R161 B.n383 B.n42 585
R162 B.n382 B.n381 585
R163 B.n380 B.n43 585
R164 B.n379 B.n378 585
R165 B.n377 B.n44 585
R166 B.n376 B.n375 585
R167 B.n374 B.n45 585
R168 B.n373 B.n372 585
R169 B.n371 B.n46 585
R170 B.n370 B.n369 585
R171 B.n368 B.n47 585
R172 B.n367 B.n366 585
R173 B.n365 B.n48 585
R174 B.n364 B.n363 585
R175 B.n362 B.n49 585
R176 B.n361 B.n360 585
R177 B.n359 B.n50 585
R178 B.n446 B.n17 585
R179 B.n448 B.n447 585
R180 B.n449 B.n16 585
R181 B.n451 B.n450 585
R182 B.n452 B.n15 585
R183 B.n454 B.n453 585
R184 B.n455 B.n14 585
R185 B.n457 B.n456 585
R186 B.n458 B.n13 585
R187 B.n460 B.n459 585
R188 B.n461 B.n12 585
R189 B.n463 B.n462 585
R190 B.n464 B.n11 585
R191 B.n466 B.n465 585
R192 B.n467 B.n10 585
R193 B.n469 B.n468 585
R194 B.n470 B.n9 585
R195 B.n472 B.n471 585
R196 B.n473 B.n8 585
R197 B.n475 B.n474 585
R198 B.n476 B.n7 585
R199 B.n478 B.n477 585
R200 B.n479 B.n6 585
R201 B.n481 B.n480 585
R202 B.n482 B.n5 585
R203 B.n484 B.n483 585
R204 B.n485 B.n4 585
R205 B.n487 B.n486 585
R206 B.n488 B.n3 585
R207 B.n490 B.n489 585
R208 B.n491 B.n0 585
R209 B.n2 B.n1 585
R210 B.n129 B.n128 585
R211 B.n130 B.n127 585
R212 B.n132 B.n131 585
R213 B.n133 B.n126 585
R214 B.n135 B.n134 585
R215 B.n136 B.n125 585
R216 B.n138 B.n137 585
R217 B.n139 B.n124 585
R218 B.n141 B.n140 585
R219 B.n142 B.n123 585
R220 B.n144 B.n143 585
R221 B.n145 B.n122 585
R222 B.n147 B.n146 585
R223 B.n148 B.n121 585
R224 B.n150 B.n149 585
R225 B.n151 B.n120 585
R226 B.n153 B.n152 585
R227 B.n154 B.n119 585
R228 B.n156 B.n155 585
R229 B.n157 B.n118 585
R230 B.n159 B.n158 585
R231 B.n160 B.n117 585
R232 B.n162 B.n161 585
R233 B.n163 B.n116 585
R234 B.n165 B.n164 585
R235 B.n166 B.n115 585
R236 B.n168 B.n167 585
R237 B.n169 B.n114 585
R238 B.n171 B.n170 585
R239 B.n172 B.n113 585
R240 B.n174 B.n113 449.257
R241 B.n263 B.n262 449.257
R242 B.n359 B.n358 449.257
R243 B.n444 B.n17 449.257
R244 B.n222 B.t7 342.084
R245 B.n36 B.t11 342.084
R246 B.n100 B.t4 342.084
R247 B.n30 B.t2 342.084
R248 B.n223 B.t8 265.478
R249 B.n37 B.t10 265.478
R250 B.n101 B.t5 265.478
R251 B.n31 B.t1 265.478
R252 B.n493 B.n492 256.663
R253 B.n100 B.t3 248.212
R254 B.n222 B.t6 248.212
R255 B.n36 B.t9 248.212
R256 B.n30 B.t0 248.212
R257 B.n492 B.n491 235.042
R258 B.n492 B.n2 235.042
R259 B.n175 B.n174 163.367
R260 B.n176 B.n175 163.367
R261 B.n176 B.n111 163.367
R262 B.n180 B.n111 163.367
R263 B.n181 B.n180 163.367
R264 B.n182 B.n181 163.367
R265 B.n182 B.n109 163.367
R266 B.n186 B.n109 163.367
R267 B.n187 B.n186 163.367
R268 B.n188 B.n187 163.367
R269 B.n188 B.n107 163.367
R270 B.n192 B.n107 163.367
R271 B.n193 B.n192 163.367
R272 B.n194 B.n193 163.367
R273 B.n194 B.n105 163.367
R274 B.n198 B.n105 163.367
R275 B.n199 B.n198 163.367
R276 B.n200 B.n199 163.367
R277 B.n200 B.n103 163.367
R278 B.n204 B.n103 163.367
R279 B.n205 B.n204 163.367
R280 B.n206 B.n205 163.367
R281 B.n206 B.n99 163.367
R282 B.n211 B.n99 163.367
R283 B.n212 B.n211 163.367
R284 B.n213 B.n212 163.367
R285 B.n213 B.n97 163.367
R286 B.n217 B.n97 163.367
R287 B.n218 B.n217 163.367
R288 B.n219 B.n218 163.367
R289 B.n219 B.n95 163.367
R290 B.n226 B.n95 163.367
R291 B.n227 B.n226 163.367
R292 B.n228 B.n227 163.367
R293 B.n228 B.n93 163.367
R294 B.n232 B.n93 163.367
R295 B.n233 B.n232 163.367
R296 B.n234 B.n233 163.367
R297 B.n234 B.n91 163.367
R298 B.n238 B.n91 163.367
R299 B.n239 B.n238 163.367
R300 B.n240 B.n239 163.367
R301 B.n240 B.n89 163.367
R302 B.n244 B.n89 163.367
R303 B.n245 B.n244 163.367
R304 B.n246 B.n245 163.367
R305 B.n246 B.n87 163.367
R306 B.n250 B.n87 163.367
R307 B.n251 B.n250 163.367
R308 B.n252 B.n251 163.367
R309 B.n252 B.n85 163.367
R310 B.n256 B.n85 163.367
R311 B.n257 B.n256 163.367
R312 B.n258 B.n257 163.367
R313 B.n258 B.n83 163.367
R314 B.n262 B.n83 163.367
R315 B.n358 B.n51 163.367
R316 B.n354 B.n51 163.367
R317 B.n354 B.n353 163.367
R318 B.n353 B.n352 163.367
R319 B.n352 B.n53 163.367
R320 B.n348 B.n53 163.367
R321 B.n348 B.n347 163.367
R322 B.n347 B.n346 163.367
R323 B.n346 B.n55 163.367
R324 B.n342 B.n55 163.367
R325 B.n342 B.n341 163.367
R326 B.n341 B.n340 163.367
R327 B.n340 B.n57 163.367
R328 B.n336 B.n57 163.367
R329 B.n336 B.n335 163.367
R330 B.n335 B.n334 163.367
R331 B.n334 B.n59 163.367
R332 B.n330 B.n59 163.367
R333 B.n330 B.n329 163.367
R334 B.n329 B.n328 163.367
R335 B.n328 B.n61 163.367
R336 B.n324 B.n61 163.367
R337 B.n324 B.n323 163.367
R338 B.n323 B.n322 163.367
R339 B.n322 B.n63 163.367
R340 B.n318 B.n63 163.367
R341 B.n318 B.n317 163.367
R342 B.n317 B.n316 163.367
R343 B.n316 B.n65 163.367
R344 B.n312 B.n65 163.367
R345 B.n312 B.n311 163.367
R346 B.n311 B.n310 163.367
R347 B.n310 B.n67 163.367
R348 B.n306 B.n67 163.367
R349 B.n306 B.n305 163.367
R350 B.n305 B.n304 163.367
R351 B.n304 B.n69 163.367
R352 B.n300 B.n69 163.367
R353 B.n300 B.n299 163.367
R354 B.n299 B.n298 163.367
R355 B.n298 B.n71 163.367
R356 B.n294 B.n71 163.367
R357 B.n294 B.n293 163.367
R358 B.n293 B.n292 163.367
R359 B.n292 B.n73 163.367
R360 B.n288 B.n73 163.367
R361 B.n288 B.n287 163.367
R362 B.n287 B.n286 163.367
R363 B.n286 B.n75 163.367
R364 B.n282 B.n75 163.367
R365 B.n282 B.n281 163.367
R366 B.n281 B.n280 163.367
R367 B.n280 B.n77 163.367
R368 B.n276 B.n77 163.367
R369 B.n276 B.n275 163.367
R370 B.n275 B.n274 163.367
R371 B.n274 B.n79 163.367
R372 B.n270 B.n79 163.367
R373 B.n270 B.n269 163.367
R374 B.n269 B.n268 163.367
R375 B.n268 B.n81 163.367
R376 B.n264 B.n81 163.367
R377 B.n264 B.n263 163.367
R378 B.n444 B.n443 163.367
R379 B.n443 B.n442 163.367
R380 B.n442 B.n19 163.367
R381 B.n438 B.n19 163.367
R382 B.n438 B.n437 163.367
R383 B.n437 B.n436 163.367
R384 B.n436 B.n21 163.367
R385 B.n432 B.n21 163.367
R386 B.n432 B.n431 163.367
R387 B.n431 B.n430 163.367
R388 B.n430 B.n23 163.367
R389 B.n426 B.n23 163.367
R390 B.n426 B.n425 163.367
R391 B.n425 B.n424 163.367
R392 B.n424 B.n25 163.367
R393 B.n420 B.n25 163.367
R394 B.n420 B.n419 163.367
R395 B.n419 B.n418 163.367
R396 B.n418 B.n27 163.367
R397 B.n414 B.n27 163.367
R398 B.n414 B.n413 163.367
R399 B.n413 B.n412 163.367
R400 B.n412 B.n29 163.367
R401 B.n407 B.n29 163.367
R402 B.n407 B.n406 163.367
R403 B.n406 B.n405 163.367
R404 B.n405 B.n33 163.367
R405 B.n401 B.n33 163.367
R406 B.n401 B.n400 163.367
R407 B.n400 B.n399 163.367
R408 B.n399 B.n35 163.367
R409 B.n395 B.n35 163.367
R410 B.n395 B.n394 163.367
R411 B.n394 B.n39 163.367
R412 B.n390 B.n39 163.367
R413 B.n390 B.n389 163.367
R414 B.n389 B.n388 163.367
R415 B.n388 B.n41 163.367
R416 B.n384 B.n41 163.367
R417 B.n384 B.n383 163.367
R418 B.n383 B.n382 163.367
R419 B.n382 B.n43 163.367
R420 B.n378 B.n43 163.367
R421 B.n378 B.n377 163.367
R422 B.n377 B.n376 163.367
R423 B.n376 B.n45 163.367
R424 B.n372 B.n45 163.367
R425 B.n372 B.n371 163.367
R426 B.n371 B.n370 163.367
R427 B.n370 B.n47 163.367
R428 B.n366 B.n47 163.367
R429 B.n366 B.n365 163.367
R430 B.n365 B.n364 163.367
R431 B.n364 B.n49 163.367
R432 B.n360 B.n49 163.367
R433 B.n360 B.n359 163.367
R434 B.n448 B.n17 163.367
R435 B.n449 B.n448 163.367
R436 B.n450 B.n449 163.367
R437 B.n450 B.n15 163.367
R438 B.n454 B.n15 163.367
R439 B.n455 B.n454 163.367
R440 B.n456 B.n455 163.367
R441 B.n456 B.n13 163.367
R442 B.n460 B.n13 163.367
R443 B.n461 B.n460 163.367
R444 B.n462 B.n461 163.367
R445 B.n462 B.n11 163.367
R446 B.n466 B.n11 163.367
R447 B.n467 B.n466 163.367
R448 B.n468 B.n467 163.367
R449 B.n468 B.n9 163.367
R450 B.n472 B.n9 163.367
R451 B.n473 B.n472 163.367
R452 B.n474 B.n473 163.367
R453 B.n474 B.n7 163.367
R454 B.n478 B.n7 163.367
R455 B.n479 B.n478 163.367
R456 B.n480 B.n479 163.367
R457 B.n480 B.n5 163.367
R458 B.n484 B.n5 163.367
R459 B.n485 B.n484 163.367
R460 B.n486 B.n485 163.367
R461 B.n486 B.n3 163.367
R462 B.n490 B.n3 163.367
R463 B.n491 B.n490 163.367
R464 B.n128 B.n2 163.367
R465 B.n128 B.n127 163.367
R466 B.n132 B.n127 163.367
R467 B.n133 B.n132 163.367
R468 B.n134 B.n133 163.367
R469 B.n134 B.n125 163.367
R470 B.n138 B.n125 163.367
R471 B.n139 B.n138 163.367
R472 B.n140 B.n139 163.367
R473 B.n140 B.n123 163.367
R474 B.n144 B.n123 163.367
R475 B.n145 B.n144 163.367
R476 B.n146 B.n145 163.367
R477 B.n146 B.n121 163.367
R478 B.n150 B.n121 163.367
R479 B.n151 B.n150 163.367
R480 B.n152 B.n151 163.367
R481 B.n152 B.n119 163.367
R482 B.n156 B.n119 163.367
R483 B.n157 B.n156 163.367
R484 B.n158 B.n157 163.367
R485 B.n158 B.n117 163.367
R486 B.n162 B.n117 163.367
R487 B.n163 B.n162 163.367
R488 B.n164 B.n163 163.367
R489 B.n164 B.n115 163.367
R490 B.n168 B.n115 163.367
R491 B.n169 B.n168 163.367
R492 B.n170 B.n169 163.367
R493 B.n170 B.n113 163.367
R494 B.n101 B.n100 76.6066
R495 B.n223 B.n222 76.6066
R496 B.n37 B.n36 76.6066
R497 B.n31 B.n30 76.6066
R498 B.n209 B.n101 59.5399
R499 B.n224 B.n223 59.5399
R500 B.n38 B.n37 59.5399
R501 B.n409 B.n31 59.5399
R502 B.n446 B.n445 29.1907
R503 B.n357 B.n50 29.1907
R504 B.n261 B.n82 29.1907
R505 B.n173 B.n172 29.1907
R506 B B.n493 18.0485
R507 B.n447 B.n446 10.6151
R508 B.n447 B.n16 10.6151
R509 B.n451 B.n16 10.6151
R510 B.n452 B.n451 10.6151
R511 B.n453 B.n452 10.6151
R512 B.n453 B.n14 10.6151
R513 B.n457 B.n14 10.6151
R514 B.n458 B.n457 10.6151
R515 B.n459 B.n458 10.6151
R516 B.n459 B.n12 10.6151
R517 B.n463 B.n12 10.6151
R518 B.n464 B.n463 10.6151
R519 B.n465 B.n464 10.6151
R520 B.n465 B.n10 10.6151
R521 B.n469 B.n10 10.6151
R522 B.n470 B.n469 10.6151
R523 B.n471 B.n470 10.6151
R524 B.n471 B.n8 10.6151
R525 B.n475 B.n8 10.6151
R526 B.n476 B.n475 10.6151
R527 B.n477 B.n476 10.6151
R528 B.n477 B.n6 10.6151
R529 B.n481 B.n6 10.6151
R530 B.n482 B.n481 10.6151
R531 B.n483 B.n482 10.6151
R532 B.n483 B.n4 10.6151
R533 B.n487 B.n4 10.6151
R534 B.n488 B.n487 10.6151
R535 B.n489 B.n488 10.6151
R536 B.n489 B.n0 10.6151
R537 B.n445 B.n18 10.6151
R538 B.n441 B.n18 10.6151
R539 B.n441 B.n440 10.6151
R540 B.n440 B.n439 10.6151
R541 B.n439 B.n20 10.6151
R542 B.n435 B.n20 10.6151
R543 B.n435 B.n434 10.6151
R544 B.n434 B.n433 10.6151
R545 B.n433 B.n22 10.6151
R546 B.n429 B.n22 10.6151
R547 B.n429 B.n428 10.6151
R548 B.n428 B.n427 10.6151
R549 B.n427 B.n24 10.6151
R550 B.n423 B.n24 10.6151
R551 B.n423 B.n422 10.6151
R552 B.n422 B.n421 10.6151
R553 B.n421 B.n26 10.6151
R554 B.n417 B.n26 10.6151
R555 B.n417 B.n416 10.6151
R556 B.n416 B.n415 10.6151
R557 B.n415 B.n28 10.6151
R558 B.n411 B.n28 10.6151
R559 B.n411 B.n410 10.6151
R560 B.n408 B.n32 10.6151
R561 B.n404 B.n32 10.6151
R562 B.n404 B.n403 10.6151
R563 B.n403 B.n402 10.6151
R564 B.n402 B.n34 10.6151
R565 B.n398 B.n34 10.6151
R566 B.n398 B.n397 10.6151
R567 B.n397 B.n396 10.6151
R568 B.n393 B.n392 10.6151
R569 B.n392 B.n391 10.6151
R570 B.n391 B.n40 10.6151
R571 B.n387 B.n40 10.6151
R572 B.n387 B.n386 10.6151
R573 B.n386 B.n385 10.6151
R574 B.n385 B.n42 10.6151
R575 B.n381 B.n42 10.6151
R576 B.n381 B.n380 10.6151
R577 B.n380 B.n379 10.6151
R578 B.n379 B.n44 10.6151
R579 B.n375 B.n44 10.6151
R580 B.n375 B.n374 10.6151
R581 B.n374 B.n373 10.6151
R582 B.n373 B.n46 10.6151
R583 B.n369 B.n46 10.6151
R584 B.n369 B.n368 10.6151
R585 B.n368 B.n367 10.6151
R586 B.n367 B.n48 10.6151
R587 B.n363 B.n48 10.6151
R588 B.n363 B.n362 10.6151
R589 B.n362 B.n361 10.6151
R590 B.n361 B.n50 10.6151
R591 B.n357 B.n356 10.6151
R592 B.n356 B.n355 10.6151
R593 B.n355 B.n52 10.6151
R594 B.n351 B.n52 10.6151
R595 B.n351 B.n350 10.6151
R596 B.n350 B.n349 10.6151
R597 B.n349 B.n54 10.6151
R598 B.n345 B.n54 10.6151
R599 B.n345 B.n344 10.6151
R600 B.n344 B.n343 10.6151
R601 B.n343 B.n56 10.6151
R602 B.n339 B.n56 10.6151
R603 B.n339 B.n338 10.6151
R604 B.n338 B.n337 10.6151
R605 B.n337 B.n58 10.6151
R606 B.n333 B.n58 10.6151
R607 B.n333 B.n332 10.6151
R608 B.n332 B.n331 10.6151
R609 B.n331 B.n60 10.6151
R610 B.n327 B.n60 10.6151
R611 B.n327 B.n326 10.6151
R612 B.n326 B.n325 10.6151
R613 B.n325 B.n62 10.6151
R614 B.n321 B.n62 10.6151
R615 B.n321 B.n320 10.6151
R616 B.n320 B.n319 10.6151
R617 B.n319 B.n64 10.6151
R618 B.n315 B.n64 10.6151
R619 B.n315 B.n314 10.6151
R620 B.n314 B.n313 10.6151
R621 B.n313 B.n66 10.6151
R622 B.n309 B.n66 10.6151
R623 B.n309 B.n308 10.6151
R624 B.n308 B.n307 10.6151
R625 B.n307 B.n68 10.6151
R626 B.n303 B.n68 10.6151
R627 B.n303 B.n302 10.6151
R628 B.n302 B.n301 10.6151
R629 B.n301 B.n70 10.6151
R630 B.n297 B.n70 10.6151
R631 B.n297 B.n296 10.6151
R632 B.n296 B.n295 10.6151
R633 B.n295 B.n72 10.6151
R634 B.n291 B.n72 10.6151
R635 B.n291 B.n290 10.6151
R636 B.n290 B.n289 10.6151
R637 B.n289 B.n74 10.6151
R638 B.n285 B.n74 10.6151
R639 B.n285 B.n284 10.6151
R640 B.n284 B.n283 10.6151
R641 B.n283 B.n76 10.6151
R642 B.n279 B.n76 10.6151
R643 B.n279 B.n278 10.6151
R644 B.n278 B.n277 10.6151
R645 B.n277 B.n78 10.6151
R646 B.n273 B.n78 10.6151
R647 B.n273 B.n272 10.6151
R648 B.n272 B.n271 10.6151
R649 B.n271 B.n80 10.6151
R650 B.n267 B.n80 10.6151
R651 B.n267 B.n266 10.6151
R652 B.n266 B.n265 10.6151
R653 B.n265 B.n82 10.6151
R654 B.n129 B.n1 10.6151
R655 B.n130 B.n129 10.6151
R656 B.n131 B.n130 10.6151
R657 B.n131 B.n126 10.6151
R658 B.n135 B.n126 10.6151
R659 B.n136 B.n135 10.6151
R660 B.n137 B.n136 10.6151
R661 B.n137 B.n124 10.6151
R662 B.n141 B.n124 10.6151
R663 B.n142 B.n141 10.6151
R664 B.n143 B.n142 10.6151
R665 B.n143 B.n122 10.6151
R666 B.n147 B.n122 10.6151
R667 B.n148 B.n147 10.6151
R668 B.n149 B.n148 10.6151
R669 B.n149 B.n120 10.6151
R670 B.n153 B.n120 10.6151
R671 B.n154 B.n153 10.6151
R672 B.n155 B.n154 10.6151
R673 B.n155 B.n118 10.6151
R674 B.n159 B.n118 10.6151
R675 B.n160 B.n159 10.6151
R676 B.n161 B.n160 10.6151
R677 B.n161 B.n116 10.6151
R678 B.n165 B.n116 10.6151
R679 B.n166 B.n165 10.6151
R680 B.n167 B.n166 10.6151
R681 B.n167 B.n114 10.6151
R682 B.n171 B.n114 10.6151
R683 B.n172 B.n171 10.6151
R684 B.n173 B.n112 10.6151
R685 B.n177 B.n112 10.6151
R686 B.n178 B.n177 10.6151
R687 B.n179 B.n178 10.6151
R688 B.n179 B.n110 10.6151
R689 B.n183 B.n110 10.6151
R690 B.n184 B.n183 10.6151
R691 B.n185 B.n184 10.6151
R692 B.n185 B.n108 10.6151
R693 B.n189 B.n108 10.6151
R694 B.n190 B.n189 10.6151
R695 B.n191 B.n190 10.6151
R696 B.n191 B.n106 10.6151
R697 B.n195 B.n106 10.6151
R698 B.n196 B.n195 10.6151
R699 B.n197 B.n196 10.6151
R700 B.n197 B.n104 10.6151
R701 B.n201 B.n104 10.6151
R702 B.n202 B.n201 10.6151
R703 B.n203 B.n202 10.6151
R704 B.n203 B.n102 10.6151
R705 B.n207 B.n102 10.6151
R706 B.n208 B.n207 10.6151
R707 B.n210 B.n98 10.6151
R708 B.n214 B.n98 10.6151
R709 B.n215 B.n214 10.6151
R710 B.n216 B.n215 10.6151
R711 B.n216 B.n96 10.6151
R712 B.n220 B.n96 10.6151
R713 B.n221 B.n220 10.6151
R714 B.n225 B.n221 10.6151
R715 B.n229 B.n94 10.6151
R716 B.n230 B.n229 10.6151
R717 B.n231 B.n230 10.6151
R718 B.n231 B.n92 10.6151
R719 B.n235 B.n92 10.6151
R720 B.n236 B.n235 10.6151
R721 B.n237 B.n236 10.6151
R722 B.n237 B.n90 10.6151
R723 B.n241 B.n90 10.6151
R724 B.n242 B.n241 10.6151
R725 B.n243 B.n242 10.6151
R726 B.n243 B.n88 10.6151
R727 B.n247 B.n88 10.6151
R728 B.n248 B.n247 10.6151
R729 B.n249 B.n248 10.6151
R730 B.n249 B.n86 10.6151
R731 B.n253 B.n86 10.6151
R732 B.n254 B.n253 10.6151
R733 B.n255 B.n254 10.6151
R734 B.n255 B.n84 10.6151
R735 B.n259 B.n84 10.6151
R736 B.n260 B.n259 10.6151
R737 B.n261 B.n260 10.6151
R738 B.n493 B.n0 8.11757
R739 B.n493 B.n1 8.11757
R740 B.n409 B.n408 6.5566
R741 B.n396 B.n38 6.5566
R742 B.n210 B.n209 6.5566
R743 B.n225 B.n224 6.5566
R744 B.n410 B.n409 4.05904
R745 B.n393 B.n38 4.05904
R746 B.n209 B.n208 4.05904
R747 B.n224 B.n94 4.05904
R748 VP.n0 VP.t0 116.814
R749 VP.n0 VP.t1 74.1048
R750 VP VP.n0 0.62124
R751 VTAIL.n118 VTAIL.n117 756.745
R752 VTAIL.n28 VTAIL.n27 756.745
R753 VTAIL.n88 VTAIL.n87 756.745
R754 VTAIL.n58 VTAIL.n57 756.745
R755 VTAIL.n101 VTAIL.n100 585
R756 VTAIL.n103 VTAIL.n102 585
R757 VTAIL.n96 VTAIL.n95 585
R758 VTAIL.n109 VTAIL.n108 585
R759 VTAIL.n111 VTAIL.n110 585
R760 VTAIL.n92 VTAIL.n91 585
R761 VTAIL.n117 VTAIL.n116 585
R762 VTAIL.n11 VTAIL.n10 585
R763 VTAIL.n13 VTAIL.n12 585
R764 VTAIL.n6 VTAIL.n5 585
R765 VTAIL.n19 VTAIL.n18 585
R766 VTAIL.n21 VTAIL.n20 585
R767 VTAIL.n2 VTAIL.n1 585
R768 VTAIL.n27 VTAIL.n26 585
R769 VTAIL.n87 VTAIL.n86 585
R770 VTAIL.n62 VTAIL.n61 585
R771 VTAIL.n81 VTAIL.n80 585
R772 VTAIL.n79 VTAIL.n78 585
R773 VTAIL.n66 VTAIL.n65 585
R774 VTAIL.n73 VTAIL.n72 585
R775 VTAIL.n71 VTAIL.n70 585
R776 VTAIL.n57 VTAIL.n56 585
R777 VTAIL.n32 VTAIL.n31 585
R778 VTAIL.n51 VTAIL.n50 585
R779 VTAIL.n49 VTAIL.n48 585
R780 VTAIL.n36 VTAIL.n35 585
R781 VTAIL.n43 VTAIL.n42 585
R782 VTAIL.n41 VTAIL.n40 585
R783 VTAIL.n99 VTAIL.t1 329.175
R784 VTAIL.n9 VTAIL.t3 329.175
R785 VTAIL.n69 VTAIL.t2 329.175
R786 VTAIL.n39 VTAIL.t0 329.175
R787 VTAIL.n102 VTAIL.n101 171.744
R788 VTAIL.n102 VTAIL.n95 171.744
R789 VTAIL.n109 VTAIL.n95 171.744
R790 VTAIL.n110 VTAIL.n109 171.744
R791 VTAIL.n110 VTAIL.n91 171.744
R792 VTAIL.n117 VTAIL.n91 171.744
R793 VTAIL.n12 VTAIL.n11 171.744
R794 VTAIL.n12 VTAIL.n5 171.744
R795 VTAIL.n19 VTAIL.n5 171.744
R796 VTAIL.n20 VTAIL.n19 171.744
R797 VTAIL.n20 VTAIL.n1 171.744
R798 VTAIL.n27 VTAIL.n1 171.744
R799 VTAIL.n87 VTAIL.n61 171.744
R800 VTAIL.n80 VTAIL.n61 171.744
R801 VTAIL.n80 VTAIL.n79 171.744
R802 VTAIL.n79 VTAIL.n65 171.744
R803 VTAIL.n72 VTAIL.n65 171.744
R804 VTAIL.n72 VTAIL.n71 171.744
R805 VTAIL.n57 VTAIL.n31 171.744
R806 VTAIL.n50 VTAIL.n31 171.744
R807 VTAIL.n50 VTAIL.n49 171.744
R808 VTAIL.n49 VTAIL.n35 171.744
R809 VTAIL.n42 VTAIL.n35 171.744
R810 VTAIL.n42 VTAIL.n41 171.744
R811 VTAIL.n101 VTAIL.t1 85.8723
R812 VTAIL.n11 VTAIL.t3 85.8723
R813 VTAIL.n71 VTAIL.t2 85.8723
R814 VTAIL.n41 VTAIL.t0 85.8723
R815 VTAIL.n119 VTAIL.n118 35.2884
R816 VTAIL.n29 VTAIL.n28 35.2884
R817 VTAIL.n89 VTAIL.n88 35.2884
R818 VTAIL.n59 VTAIL.n58 35.2884
R819 VTAIL.n59 VTAIL.n29 24.2289
R820 VTAIL.n119 VTAIL.n89 20.8238
R821 VTAIL.n116 VTAIL.n90 12.0247
R822 VTAIL.n26 VTAIL.n0 12.0247
R823 VTAIL.n86 VTAIL.n60 12.0247
R824 VTAIL.n56 VTAIL.n30 12.0247
R825 VTAIL.n115 VTAIL.n92 11.249
R826 VTAIL.n25 VTAIL.n2 11.249
R827 VTAIL.n85 VTAIL.n62 11.249
R828 VTAIL.n55 VTAIL.n32 11.249
R829 VTAIL.n100 VTAIL.n99 10.722
R830 VTAIL.n10 VTAIL.n9 10.722
R831 VTAIL.n70 VTAIL.n69 10.722
R832 VTAIL.n40 VTAIL.n39 10.722
R833 VTAIL.n112 VTAIL.n111 10.4732
R834 VTAIL.n22 VTAIL.n21 10.4732
R835 VTAIL.n82 VTAIL.n81 10.4732
R836 VTAIL.n52 VTAIL.n51 10.4732
R837 VTAIL.n108 VTAIL.n94 9.69747
R838 VTAIL.n18 VTAIL.n4 9.69747
R839 VTAIL.n78 VTAIL.n64 9.69747
R840 VTAIL.n48 VTAIL.n34 9.69747
R841 VTAIL.n114 VTAIL.n90 9.45567
R842 VTAIL.n24 VTAIL.n0 9.45567
R843 VTAIL.n84 VTAIL.n60 9.45567
R844 VTAIL.n54 VTAIL.n30 9.45567
R845 VTAIL.n98 VTAIL.n97 9.3005
R846 VTAIL.n105 VTAIL.n104 9.3005
R847 VTAIL.n107 VTAIL.n106 9.3005
R848 VTAIL.n94 VTAIL.n93 9.3005
R849 VTAIL.n113 VTAIL.n112 9.3005
R850 VTAIL.n115 VTAIL.n114 9.3005
R851 VTAIL.n8 VTAIL.n7 9.3005
R852 VTAIL.n15 VTAIL.n14 9.3005
R853 VTAIL.n17 VTAIL.n16 9.3005
R854 VTAIL.n4 VTAIL.n3 9.3005
R855 VTAIL.n23 VTAIL.n22 9.3005
R856 VTAIL.n25 VTAIL.n24 9.3005
R857 VTAIL.n85 VTAIL.n84 9.3005
R858 VTAIL.n83 VTAIL.n82 9.3005
R859 VTAIL.n64 VTAIL.n63 9.3005
R860 VTAIL.n77 VTAIL.n76 9.3005
R861 VTAIL.n75 VTAIL.n74 9.3005
R862 VTAIL.n68 VTAIL.n67 9.3005
R863 VTAIL.n45 VTAIL.n44 9.3005
R864 VTAIL.n47 VTAIL.n46 9.3005
R865 VTAIL.n34 VTAIL.n33 9.3005
R866 VTAIL.n53 VTAIL.n52 9.3005
R867 VTAIL.n55 VTAIL.n54 9.3005
R868 VTAIL.n38 VTAIL.n37 9.3005
R869 VTAIL.n107 VTAIL.n96 8.92171
R870 VTAIL.n17 VTAIL.n6 8.92171
R871 VTAIL.n77 VTAIL.n66 8.92171
R872 VTAIL.n47 VTAIL.n36 8.92171
R873 VTAIL.n104 VTAIL.n103 8.14595
R874 VTAIL.n14 VTAIL.n13 8.14595
R875 VTAIL.n74 VTAIL.n73 8.14595
R876 VTAIL.n44 VTAIL.n43 8.14595
R877 VTAIL.n100 VTAIL.n98 7.3702
R878 VTAIL.n10 VTAIL.n8 7.3702
R879 VTAIL.n70 VTAIL.n68 7.3702
R880 VTAIL.n40 VTAIL.n38 7.3702
R881 VTAIL.n103 VTAIL.n98 5.81868
R882 VTAIL.n13 VTAIL.n8 5.81868
R883 VTAIL.n73 VTAIL.n68 5.81868
R884 VTAIL.n43 VTAIL.n38 5.81868
R885 VTAIL.n104 VTAIL.n96 5.04292
R886 VTAIL.n14 VTAIL.n6 5.04292
R887 VTAIL.n74 VTAIL.n66 5.04292
R888 VTAIL.n44 VTAIL.n36 5.04292
R889 VTAIL.n108 VTAIL.n107 4.26717
R890 VTAIL.n18 VTAIL.n17 4.26717
R891 VTAIL.n78 VTAIL.n77 4.26717
R892 VTAIL.n48 VTAIL.n47 4.26717
R893 VTAIL.n111 VTAIL.n94 3.49141
R894 VTAIL.n21 VTAIL.n4 3.49141
R895 VTAIL.n81 VTAIL.n64 3.49141
R896 VTAIL.n51 VTAIL.n34 3.49141
R897 VTAIL.n112 VTAIL.n92 2.71565
R898 VTAIL.n22 VTAIL.n2 2.71565
R899 VTAIL.n82 VTAIL.n62 2.71565
R900 VTAIL.n52 VTAIL.n32 2.71565
R901 VTAIL.n99 VTAIL.n97 2.4147
R902 VTAIL.n9 VTAIL.n7 2.4147
R903 VTAIL.n69 VTAIL.n67 2.4147
R904 VTAIL.n39 VTAIL.n37 2.4147
R905 VTAIL.n89 VTAIL.n59 2.17291
R906 VTAIL.n116 VTAIL.n115 1.93989
R907 VTAIL.n26 VTAIL.n25 1.93989
R908 VTAIL.n86 VTAIL.n85 1.93989
R909 VTAIL.n56 VTAIL.n55 1.93989
R910 VTAIL VTAIL.n29 1.37981
R911 VTAIL.n118 VTAIL.n90 1.16414
R912 VTAIL.n28 VTAIL.n0 1.16414
R913 VTAIL.n88 VTAIL.n60 1.16414
R914 VTAIL.n58 VTAIL.n30 1.16414
R915 VTAIL VTAIL.n119 0.793603
R916 VTAIL.n105 VTAIL.n97 0.155672
R917 VTAIL.n106 VTAIL.n105 0.155672
R918 VTAIL.n106 VTAIL.n93 0.155672
R919 VTAIL.n113 VTAIL.n93 0.155672
R920 VTAIL.n114 VTAIL.n113 0.155672
R921 VTAIL.n15 VTAIL.n7 0.155672
R922 VTAIL.n16 VTAIL.n15 0.155672
R923 VTAIL.n16 VTAIL.n3 0.155672
R924 VTAIL.n23 VTAIL.n3 0.155672
R925 VTAIL.n24 VTAIL.n23 0.155672
R926 VTAIL.n84 VTAIL.n83 0.155672
R927 VTAIL.n83 VTAIL.n63 0.155672
R928 VTAIL.n76 VTAIL.n63 0.155672
R929 VTAIL.n76 VTAIL.n75 0.155672
R930 VTAIL.n75 VTAIL.n67 0.155672
R931 VTAIL.n54 VTAIL.n53 0.155672
R932 VTAIL.n53 VTAIL.n33 0.155672
R933 VTAIL.n46 VTAIL.n33 0.155672
R934 VTAIL.n46 VTAIL.n45 0.155672
R935 VTAIL.n45 VTAIL.n37 0.155672
R936 VDD1.n28 VDD1.n27 756.745
R937 VDD1.n57 VDD1.n56 756.745
R938 VDD1.n27 VDD1.n26 585
R939 VDD1.n2 VDD1.n1 585
R940 VDD1.n21 VDD1.n20 585
R941 VDD1.n19 VDD1.n18 585
R942 VDD1.n6 VDD1.n5 585
R943 VDD1.n13 VDD1.n12 585
R944 VDD1.n11 VDD1.n10 585
R945 VDD1.n40 VDD1.n39 585
R946 VDD1.n42 VDD1.n41 585
R947 VDD1.n35 VDD1.n34 585
R948 VDD1.n48 VDD1.n47 585
R949 VDD1.n50 VDD1.n49 585
R950 VDD1.n31 VDD1.n30 585
R951 VDD1.n56 VDD1.n55 585
R952 VDD1.n38 VDD1.t0 329.175
R953 VDD1.n9 VDD1.t1 329.175
R954 VDD1.n27 VDD1.n1 171.744
R955 VDD1.n20 VDD1.n1 171.744
R956 VDD1.n20 VDD1.n19 171.744
R957 VDD1.n19 VDD1.n5 171.744
R958 VDD1.n12 VDD1.n5 171.744
R959 VDD1.n12 VDD1.n11 171.744
R960 VDD1.n41 VDD1.n40 171.744
R961 VDD1.n41 VDD1.n34 171.744
R962 VDD1.n48 VDD1.n34 171.744
R963 VDD1.n49 VDD1.n48 171.744
R964 VDD1.n49 VDD1.n30 171.744
R965 VDD1.n56 VDD1.n30 171.744
R966 VDD1 VDD1.n57 88.8648
R967 VDD1.n11 VDD1.t1 85.8723
R968 VDD1.n40 VDD1.t0 85.8723
R969 VDD1 VDD1.n28 52.8766
R970 VDD1.n26 VDD1.n0 12.0247
R971 VDD1.n55 VDD1.n29 12.0247
R972 VDD1.n25 VDD1.n2 11.249
R973 VDD1.n54 VDD1.n31 11.249
R974 VDD1.n10 VDD1.n9 10.722
R975 VDD1.n39 VDD1.n38 10.722
R976 VDD1.n22 VDD1.n21 10.4732
R977 VDD1.n51 VDD1.n50 10.4732
R978 VDD1.n18 VDD1.n4 9.69747
R979 VDD1.n47 VDD1.n33 9.69747
R980 VDD1.n24 VDD1.n0 9.45567
R981 VDD1.n53 VDD1.n29 9.45567
R982 VDD1.n25 VDD1.n24 9.3005
R983 VDD1.n23 VDD1.n22 9.3005
R984 VDD1.n4 VDD1.n3 9.3005
R985 VDD1.n17 VDD1.n16 9.3005
R986 VDD1.n15 VDD1.n14 9.3005
R987 VDD1.n8 VDD1.n7 9.3005
R988 VDD1.n37 VDD1.n36 9.3005
R989 VDD1.n44 VDD1.n43 9.3005
R990 VDD1.n46 VDD1.n45 9.3005
R991 VDD1.n33 VDD1.n32 9.3005
R992 VDD1.n52 VDD1.n51 9.3005
R993 VDD1.n54 VDD1.n53 9.3005
R994 VDD1.n17 VDD1.n6 8.92171
R995 VDD1.n46 VDD1.n35 8.92171
R996 VDD1.n14 VDD1.n13 8.14595
R997 VDD1.n43 VDD1.n42 8.14595
R998 VDD1.n10 VDD1.n8 7.3702
R999 VDD1.n39 VDD1.n37 7.3702
R1000 VDD1.n13 VDD1.n8 5.81868
R1001 VDD1.n42 VDD1.n37 5.81868
R1002 VDD1.n14 VDD1.n6 5.04292
R1003 VDD1.n43 VDD1.n35 5.04292
R1004 VDD1.n18 VDD1.n17 4.26717
R1005 VDD1.n47 VDD1.n46 4.26717
R1006 VDD1.n21 VDD1.n4 3.49141
R1007 VDD1.n50 VDD1.n33 3.49141
R1008 VDD1.n22 VDD1.n2 2.71565
R1009 VDD1.n51 VDD1.n31 2.71565
R1010 VDD1.n38 VDD1.n36 2.4147
R1011 VDD1.n9 VDD1.n7 2.4147
R1012 VDD1.n26 VDD1.n25 1.93989
R1013 VDD1.n55 VDD1.n54 1.93989
R1014 VDD1.n28 VDD1.n0 1.16414
R1015 VDD1.n57 VDD1.n29 1.16414
R1016 VDD1.n24 VDD1.n23 0.155672
R1017 VDD1.n23 VDD1.n3 0.155672
R1018 VDD1.n16 VDD1.n3 0.155672
R1019 VDD1.n16 VDD1.n15 0.155672
R1020 VDD1.n15 VDD1.n7 0.155672
R1021 VDD1.n44 VDD1.n36 0.155672
R1022 VDD1.n45 VDD1.n44 0.155672
R1023 VDD1.n45 VDD1.n32 0.155672
R1024 VDD1.n52 VDD1.n32 0.155672
R1025 VDD1.n53 VDD1.n52 0.155672
R1026 VN VN.t0 116.627
R1027 VN VN.t1 74.7255
R1028 VDD2.n57 VDD2.n56 756.745
R1029 VDD2.n28 VDD2.n27 756.745
R1030 VDD2.n56 VDD2.n55 585
R1031 VDD2.n31 VDD2.n30 585
R1032 VDD2.n50 VDD2.n49 585
R1033 VDD2.n48 VDD2.n47 585
R1034 VDD2.n35 VDD2.n34 585
R1035 VDD2.n42 VDD2.n41 585
R1036 VDD2.n40 VDD2.n39 585
R1037 VDD2.n11 VDD2.n10 585
R1038 VDD2.n13 VDD2.n12 585
R1039 VDD2.n6 VDD2.n5 585
R1040 VDD2.n19 VDD2.n18 585
R1041 VDD2.n21 VDD2.n20 585
R1042 VDD2.n2 VDD2.n1 585
R1043 VDD2.n27 VDD2.n26 585
R1044 VDD2.n9 VDD2.t0 329.175
R1045 VDD2.n38 VDD2.t1 329.175
R1046 VDD2.n56 VDD2.n30 171.744
R1047 VDD2.n49 VDD2.n30 171.744
R1048 VDD2.n49 VDD2.n48 171.744
R1049 VDD2.n48 VDD2.n34 171.744
R1050 VDD2.n41 VDD2.n34 171.744
R1051 VDD2.n41 VDD2.n40 171.744
R1052 VDD2.n12 VDD2.n11 171.744
R1053 VDD2.n12 VDD2.n5 171.744
R1054 VDD2.n19 VDD2.n5 171.744
R1055 VDD2.n20 VDD2.n19 171.744
R1056 VDD2.n20 VDD2.n1 171.744
R1057 VDD2.n27 VDD2.n1 171.744
R1058 VDD2.n58 VDD2.n28 87.4887
R1059 VDD2.n40 VDD2.t1 85.8723
R1060 VDD2.n11 VDD2.t0 85.8723
R1061 VDD2.n58 VDD2.n57 51.9672
R1062 VDD2.n55 VDD2.n29 12.0247
R1063 VDD2.n26 VDD2.n0 12.0247
R1064 VDD2.n54 VDD2.n31 11.249
R1065 VDD2.n25 VDD2.n2 11.249
R1066 VDD2.n39 VDD2.n38 10.722
R1067 VDD2.n10 VDD2.n9 10.722
R1068 VDD2.n51 VDD2.n50 10.4732
R1069 VDD2.n22 VDD2.n21 10.4732
R1070 VDD2.n47 VDD2.n33 9.69747
R1071 VDD2.n18 VDD2.n4 9.69747
R1072 VDD2.n53 VDD2.n29 9.45567
R1073 VDD2.n24 VDD2.n0 9.45567
R1074 VDD2.n54 VDD2.n53 9.3005
R1075 VDD2.n52 VDD2.n51 9.3005
R1076 VDD2.n33 VDD2.n32 9.3005
R1077 VDD2.n46 VDD2.n45 9.3005
R1078 VDD2.n44 VDD2.n43 9.3005
R1079 VDD2.n37 VDD2.n36 9.3005
R1080 VDD2.n8 VDD2.n7 9.3005
R1081 VDD2.n15 VDD2.n14 9.3005
R1082 VDD2.n17 VDD2.n16 9.3005
R1083 VDD2.n4 VDD2.n3 9.3005
R1084 VDD2.n23 VDD2.n22 9.3005
R1085 VDD2.n25 VDD2.n24 9.3005
R1086 VDD2.n46 VDD2.n35 8.92171
R1087 VDD2.n17 VDD2.n6 8.92171
R1088 VDD2.n43 VDD2.n42 8.14595
R1089 VDD2.n14 VDD2.n13 8.14595
R1090 VDD2.n39 VDD2.n37 7.3702
R1091 VDD2.n10 VDD2.n8 7.3702
R1092 VDD2.n42 VDD2.n37 5.81868
R1093 VDD2.n13 VDD2.n8 5.81868
R1094 VDD2.n43 VDD2.n35 5.04292
R1095 VDD2.n14 VDD2.n6 5.04292
R1096 VDD2.n47 VDD2.n46 4.26717
R1097 VDD2.n18 VDD2.n17 4.26717
R1098 VDD2.n50 VDD2.n33 3.49141
R1099 VDD2.n21 VDD2.n4 3.49141
R1100 VDD2.n51 VDD2.n31 2.71565
R1101 VDD2.n22 VDD2.n2 2.71565
R1102 VDD2.n9 VDD2.n7 2.4147
R1103 VDD2.n38 VDD2.n36 2.4147
R1104 VDD2.n55 VDD2.n54 1.93989
R1105 VDD2.n26 VDD2.n25 1.93989
R1106 VDD2.n57 VDD2.n29 1.16414
R1107 VDD2.n28 VDD2.n0 1.16414
R1108 VDD2 VDD2.n58 0.909983
R1109 VDD2.n53 VDD2.n52 0.155672
R1110 VDD2.n52 VDD2.n32 0.155672
R1111 VDD2.n45 VDD2.n32 0.155672
R1112 VDD2.n45 VDD2.n44 0.155672
R1113 VDD2.n44 VDD2.n36 0.155672
R1114 VDD2.n15 VDD2.n7 0.155672
R1115 VDD2.n16 VDD2.n15 0.155672
R1116 VDD2.n16 VDD2.n3 0.155672
R1117 VDD2.n23 VDD2.n3 0.155672
R1118 VDD2.n24 VDD2.n23 0.155672
C0 VDD1 VP 1.77825f
C1 B VP 1.68872f
C2 VDD1 VDD2 0.784645f
C3 B VDD2 1.3849f
C4 VN VTAIL 1.68557f
C5 B VDD1 1.34566f
C6 w_n2550_n2140# VTAIL 1.9355f
C7 VP VTAIL 1.6998f
C8 VDD2 VTAIL 3.78866f
C9 VDD1 VTAIL 3.72934f
C10 B VTAIL 2.56052f
C11 VN w_n2550_n2140# 3.51347f
C12 VN VP 4.79877f
C13 VN VDD2 1.55262f
C14 VN VDD1 0.148925f
C15 VN B 1.147f
C16 w_n2550_n2140# VP 3.84048f
C17 w_n2550_n2140# VDD2 1.51406f
C18 VDD2 VP 0.37583f
C19 w_n2550_n2140# VDD1 1.47561f
C20 B w_n2550_n2140# 8.20557f
C21 VDD2 VSUBS 0.755981f
C22 VDD1 VSUBS 2.621899f
C23 VTAIL VSUBS 0.569268f
C24 VN VSUBS 5.85775f
C25 VP VSUBS 1.633079f
C26 B VSUBS 4.139167f
C27 w_n2550_n2140# VSUBS 68.14621f
C28 VDD2.n0 VSUBS 0.008588f
C29 VDD2.n1 VSUBS 0.019331f
C30 VDD2.n2 VSUBS 0.00866f
C31 VDD2.n3 VSUBS 0.01522f
C32 VDD2.n4 VSUBS 0.008179f
C33 VDD2.n5 VSUBS 0.019331f
C34 VDD2.n6 VSUBS 0.00866f
C35 VDD2.n7 VSUBS 0.337753f
C36 VDD2.n8 VSUBS 0.008179f
C37 VDD2.t0 VSUBS 0.04167f
C38 VDD2.n9 VSUBS 0.077876f
C39 VDD2.n10 VSUBS 0.014536f
C40 VDD2.n11 VSUBS 0.014498f
C41 VDD2.n12 VSUBS 0.019331f
C42 VDD2.n13 VSUBS 0.00866f
C43 VDD2.n14 VSUBS 0.008179f
C44 VDD2.n15 VSUBS 0.01522f
C45 VDD2.n16 VSUBS 0.01522f
C46 VDD2.n17 VSUBS 0.008179f
C47 VDD2.n18 VSUBS 0.00866f
C48 VDD2.n19 VSUBS 0.019331f
C49 VDD2.n20 VSUBS 0.019331f
C50 VDD2.n21 VSUBS 0.00866f
C51 VDD2.n22 VSUBS 0.008179f
C52 VDD2.n23 VSUBS 0.01522f
C53 VDD2.n24 VSUBS 0.039755f
C54 VDD2.n25 VSUBS 0.008179f
C55 VDD2.n26 VSUBS 0.00866f
C56 VDD2.n27 VSUBS 0.043505f
C57 VDD2.n28 VSUBS 0.355078f
C58 VDD2.n29 VSUBS 0.008588f
C59 VDD2.n30 VSUBS 0.019331f
C60 VDD2.n31 VSUBS 0.00866f
C61 VDD2.n32 VSUBS 0.01522f
C62 VDD2.n33 VSUBS 0.008179f
C63 VDD2.n34 VSUBS 0.019331f
C64 VDD2.n35 VSUBS 0.00866f
C65 VDD2.n36 VSUBS 0.337753f
C66 VDD2.n37 VSUBS 0.008179f
C67 VDD2.t1 VSUBS 0.04167f
C68 VDD2.n38 VSUBS 0.077876f
C69 VDD2.n39 VSUBS 0.014536f
C70 VDD2.n40 VSUBS 0.014498f
C71 VDD2.n41 VSUBS 0.019331f
C72 VDD2.n42 VSUBS 0.00866f
C73 VDD2.n43 VSUBS 0.008179f
C74 VDD2.n44 VSUBS 0.01522f
C75 VDD2.n45 VSUBS 0.01522f
C76 VDD2.n46 VSUBS 0.008179f
C77 VDD2.n47 VSUBS 0.00866f
C78 VDD2.n48 VSUBS 0.019331f
C79 VDD2.n49 VSUBS 0.019331f
C80 VDD2.n50 VSUBS 0.00866f
C81 VDD2.n51 VSUBS 0.008179f
C82 VDD2.n52 VSUBS 0.01522f
C83 VDD2.n53 VSUBS 0.039755f
C84 VDD2.n54 VSUBS 0.008179f
C85 VDD2.n55 VSUBS 0.00866f
C86 VDD2.n56 VSUBS 0.043505f
C87 VDD2.n57 VSUBS 0.039746f
C88 VDD2.n58 VSUBS 1.60316f
C89 VN.t1 VSUBS 2.11168f
C90 VN.t0 VSUBS 2.83933f
C91 VDD1.n0 VSUBS 0.00824f
C92 VDD1.n1 VSUBS 0.018548f
C93 VDD1.n2 VSUBS 0.008309f
C94 VDD1.n3 VSUBS 0.014604f
C95 VDD1.n4 VSUBS 0.007847f
C96 VDD1.n5 VSUBS 0.018548f
C97 VDD1.n6 VSUBS 0.008309f
C98 VDD1.n7 VSUBS 0.324071f
C99 VDD1.n8 VSUBS 0.007847f
C100 VDD1.t1 VSUBS 0.039982f
C101 VDD1.n9 VSUBS 0.074721f
C102 VDD1.n10 VSUBS 0.013947f
C103 VDD1.n11 VSUBS 0.013911f
C104 VDD1.n12 VSUBS 0.018548f
C105 VDD1.n13 VSUBS 0.008309f
C106 VDD1.n14 VSUBS 0.007847f
C107 VDD1.n15 VSUBS 0.014604f
C108 VDD1.n16 VSUBS 0.014604f
C109 VDD1.n17 VSUBS 0.007847f
C110 VDD1.n18 VSUBS 0.008309f
C111 VDD1.n19 VSUBS 0.018548f
C112 VDD1.n20 VSUBS 0.018548f
C113 VDD1.n21 VSUBS 0.008309f
C114 VDD1.n22 VSUBS 0.007847f
C115 VDD1.n23 VSUBS 0.014604f
C116 VDD1.n24 VSUBS 0.038144f
C117 VDD1.n25 VSUBS 0.007847f
C118 VDD1.n26 VSUBS 0.008309f
C119 VDD1.n27 VSUBS 0.041743f
C120 VDD1.n28 VSUBS 0.039387f
C121 VDD1.n29 VSUBS 0.00824f
C122 VDD1.n30 VSUBS 0.018548f
C123 VDD1.n31 VSUBS 0.008309f
C124 VDD1.n32 VSUBS 0.014604f
C125 VDD1.n33 VSUBS 0.007847f
C126 VDD1.n34 VSUBS 0.018548f
C127 VDD1.n35 VSUBS 0.008309f
C128 VDD1.n36 VSUBS 0.324071f
C129 VDD1.n37 VSUBS 0.007847f
C130 VDD1.t0 VSUBS 0.039982f
C131 VDD1.n38 VSUBS 0.074721f
C132 VDD1.n39 VSUBS 0.013947f
C133 VDD1.n40 VSUBS 0.013911f
C134 VDD1.n41 VSUBS 0.018548f
C135 VDD1.n42 VSUBS 0.008309f
C136 VDD1.n43 VSUBS 0.007847f
C137 VDD1.n44 VSUBS 0.014604f
C138 VDD1.n45 VSUBS 0.014604f
C139 VDD1.n46 VSUBS 0.007847f
C140 VDD1.n47 VSUBS 0.008309f
C141 VDD1.n48 VSUBS 0.018548f
C142 VDD1.n49 VSUBS 0.018548f
C143 VDD1.n50 VSUBS 0.008309f
C144 VDD1.n51 VSUBS 0.007847f
C145 VDD1.n52 VSUBS 0.014604f
C146 VDD1.n53 VSUBS 0.038144f
C147 VDD1.n54 VSUBS 0.007847f
C148 VDD1.n55 VSUBS 0.008309f
C149 VDD1.n56 VSUBS 0.041743f
C150 VDD1.n57 VSUBS 0.370044f
C151 VTAIL.n0 VSUBS 0.012813f
C152 VTAIL.n1 VSUBS 0.028841f
C153 VTAIL.n2 VSUBS 0.01292f
C154 VTAIL.n3 VSUBS 0.022708f
C155 VTAIL.n4 VSUBS 0.012202f
C156 VTAIL.n5 VSUBS 0.028841f
C157 VTAIL.n6 VSUBS 0.01292f
C158 VTAIL.n7 VSUBS 0.50391f
C159 VTAIL.n8 VSUBS 0.012202f
C160 VTAIL.t3 VSUBS 0.06217f
C161 VTAIL.n9 VSUBS 0.116187f
C162 VTAIL.n10 VSUBS 0.021687f
C163 VTAIL.n11 VSUBS 0.021631f
C164 VTAIL.n12 VSUBS 0.028841f
C165 VTAIL.n13 VSUBS 0.01292f
C166 VTAIL.n14 VSUBS 0.012202f
C167 VTAIL.n15 VSUBS 0.022708f
C168 VTAIL.n16 VSUBS 0.022708f
C169 VTAIL.n17 VSUBS 0.012202f
C170 VTAIL.n18 VSUBS 0.01292f
C171 VTAIL.n19 VSUBS 0.028841f
C172 VTAIL.n20 VSUBS 0.028841f
C173 VTAIL.n21 VSUBS 0.01292f
C174 VTAIL.n22 VSUBS 0.012202f
C175 VTAIL.n23 VSUBS 0.022708f
C176 VTAIL.n24 VSUBS 0.059312f
C177 VTAIL.n25 VSUBS 0.012202f
C178 VTAIL.n26 VSUBS 0.01292f
C179 VTAIL.n27 VSUBS 0.064907f
C180 VTAIL.n28 VSUBS 0.043655f
C181 VTAIL.n29 VSUBS 1.29951f
C182 VTAIL.n30 VSUBS 0.012813f
C183 VTAIL.n31 VSUBS 0.028841f
C184 VTAIL.n32 VSUBS 0.01292f
C185 VTAIL.n33 VSUBS 0.022708f
C186 VTAIL.n34 VSUBS 0.012202f
C187 VTAIL.n35 VSUBS 0.028841f
C188 VTAIL.n36 VSUBS 0.01292f
C189 VTAIL.n37 VSUBS 0.50391f
C190 VTAIL.n38 VSUBS 0.012202f
C191 VTAIL.t0 VSUBS 0.06217f
C192 VTAIL.n39 VSUBS 0.116187f
C193 VTAIL.n40 VSUBS 0.021687f
C194 VTAIL.n41 VSUBS 0.021631f
C195 VTAIL.n42 VSUBS 0.028841f
C196 VTAIL.n43 VSUBS 0.01292f
C197 VTAIL.n44 VSUBS 0.012202f
C198 VTAIL.n45 VSUBS 0.022708f
C199 VTAIL.n46 VSUBS 0.022708f
C200 VTAIL.n47 VSUBS 0.012202f
C201 VTAIL.n48 VSUBS 0.01292f
C202 VTAIL.n49 VSUBS 0.028841f
C203 VTAIL.n50 VSUBS 0.028841f
C204 VTAIL.n51 VSUBS 0.01292f
C205 VTAIL.n52 VSUBS 0.012202f
C206 VTAIL.n53 VSUBS 0.022708f
C207 VTAIL.n54 VSUBS 0.059312f
C208 VTAIL.n55 VSUBS 0.012202f
C209 VTAIL.n56 VSUBS 0.01292f
C210 VTAIL.n57 VSUBS 0.064907f
C211 VTAIL.n58 VSUBS 0.043655f
C212 VTAIL.n59 VSUBS 1.35754f
C213 VTAIL.n60 VSUBS 0.012813f
C214 VTAIL.n61 VSUBS 0.028841f
C215 VTAIL.n62 VSUBS 0.01292f
C216 VTAIL.n63 VSUBS 0.022708f
C217 VTAIL.n64 VSUBS 0.012202f
C218 VTAIL.n65 VSUBS 0.028841f
C219 VTAIL.n66 VSUBS 0.01292f
C220 VTAIL.n67 VSUBS 0.50391f
C221 VTAIL.n68 VSUBS 0.012202f
C222 VTAIL.t2 VSUBS 0.06217f
C223 VTAIL.n69 VSUBS 0.116187f
C224 VTAIL.n70 VSUBS 0.021687f
C225 VTAIL.n71 VSUBS 0.021631f
C226 VTAIL.n72 VSUBS 0.028841f
C227 VTAIL.n73 VSUBS 0.01292f
C228 VTAIL.n74 VSUBS 0.012202f
C229 VTAIL.n75 VSUBS 0.022708f
C230 VTAIL.n76 VSUBS 0.022708f
C231 VTAIL.n77 VSUBS 0.012202f
C232 VTAIL.n78 VSUBS 0.01292f
C233 VTAIL.n79 VSUBS 0.028841f
C234 VTAIL.n80 VSUBS 0.028841f
C235 VTAIL.n81 VSUBS 0.01292f
C236 VTAIL.n82 VSUBS 0.012202f
C237 VTAIL.n83 VSUBS 0.022708f
C238 VTAIL.n84 VSUBS 0.059312f
C239 VTAIL.n85 VSUBS 0.012202f
C240 VTAIL.n86 VSUBS 0.01292f
C241 VTAIL.n87 VSUBS 0.064907f
C242 VTAIL.n88 VSUBS 0.043655f
C243 VTAIL.n89 VSUBS 1.10839f
C244 VTAIL.n90 VSUBS 0.012813f
C245 VTAIL.n91 VSUBS 0.028841f
C246 VTAIL.n92 VSUBS 0.01292f
C247 VTAIL.n93 VSUBS 0.022708f
C248 VTAIL.n94 VSUBS 0.012202f
C249 VTAIL.n95 VSUBS 0.028841f
C250 VTAIL.n96 VSUBS 0.01292f
C251 VTAIL.n97 VSUBS 0.50391f
C252 VTAIL.n98 VSUBS 0.012202f
C253 VTAIL.t1 VSUBS 0.06217f
C254 VTAIL.n99 VSUBS 0.116187f
C255 VTAIL.n100 VSUBS 0.021687f
C256 VTAIL.n101 VSUBS 0.021631f
C257 VTAIL.n102 VSUBS 0.028841f
C258 VTAIL.n103 VSUBS 0.01292f
C259 VTAIL.n104 VSUBS 0.012202f
C260 VTAIL.n105 VSUBS 0.022708f
C261 VTAIL.n106 VSUBS 0.022708f
C262 VTAIL.n107 VSUBS 0.012202f
C263 VTAIL.n108 VSUBS 0.01292f
C264 VTAIL.n109 VSUBS 0.028841f
C265 VTAIL.n110 VSUBS 0.028841f
C266 VTAIL.n111 VSUBS 0.01292f
C267 VTAIL.n112 VSUBS 0.012202f
C268 VTAIL.n113 VSUBS 0.022708f
C269 VTAIL.n114 VSUBS 0.059312f
C270 VTAIL.n115 VSUBS 0.012202f
C271 VTAIL.n116 VSUBS 0.01292f
C272 VTAIL.n117 VSUBS 0.064907f
C273 VTAIL.n118 VSUBS 0.043655f
C274 VTAIL.n119 VSUBS 1.00746f
C275 VP.t0 VSUBS 2.95869f
C276 VP.t1 VSUBS 2.1933f
C277 VP.n0 VSUBS 3.32145f
C278 B.n0 VSUBS 0.006726f
C279 B.n1 VSUBS 0.006726f
C280 B.n2 VSUBS 0.009947f
C281 B.n3 VSUBS 0.007623f
C282 B.n4 VSUBS 0.007623f
C283 B.n5 VSUBS 0.007623f
C284 B.n6 VSUBS 0.007623f
C285 B.n7 VSUBS 0.007623f
C286 B.n8 VSUBS 0.007623f
C287 B.n9 VSUBS 0.007623f
C288 B.n10 VSUBS 0.007623f
C289 B.n11 VSUBS 0.007623f
C290 B.n12 VSUBS 0.007623f
C291 B.n13 VSUBS 0.007623f
C292 B.n14 VSUBS 0.007623f
C293 B.n15 VSUBS 0.007623f
C294 B.n16 VSUBS 0.007623f
C295 B.n17 VSUBS 0.016111f
C296 B.n18 VSUBS 0.007623f
C297 B.n19 VSUBS 0.007623f
C298 B.n20 VSUBS 0.007623f
C299 B.n21 VSUBS 0.007623f
C300 B.n22 VSUBS 0.007623f
C301 B.n23 VSUBS 0.007623f
C302 B.n24 VSUBS 0.007623f
C303 B.n25 VSUBS 0.007623f
C304 B.n26 VSUBS 0.007623f
C305 B.n27 VSUBS 0.007623f
C306 B.n28 VSUBS 0.007623f
C307 B.n29 VSUBS 0.007623f
C308 B.t1 VSUBS 0.094501f
C309 B.t2 VSUBS 0.130673f
C310 B.t0 VSUBS 1.10947f
C311 B.n30 VSUBS 0.217472f
C312 B.n31 VSUBS 0.172396f
C313 B.n32 VSUBS 0.007623f
C314 B.n33 VSUBS 0.007623f
C315 B.n34 VSUBS 0.007623f
C316 B.n35 VSUBS 0.007623f
C317 B.t10 VSUBS 0.094503f
C318 B.t11 VSUBS 0.130674f
C319 B.t9 VSUBS 1.10947f
C320 B.n36 VSUBS 0.21747f
C321 B.n37 VSUBS 0.172394f
C322 B.n38 VSUBS 0.017661f
C323 B.n39 VSUBS 0.007623f
C324 B.n40 VSUBS 0.007623f
C325 B.n41 VSUBS 0.007623f
C326 B.n42 VSUBS 0.007623f
C327 B.n43 VSUBS 0.007623f
C328 B.n44 VSUBS 0.007623f
C329 B.n45 VSUBS 0.007623f
C330 B.n46 VSUBS 0.007623f
C331 B.n47 VSUBS 0.007623f
C332 B.n48 VSUBS 0.007623f
C333 B.n49 VSUBS 0.007623f
C334 B.n50 VSUBS 0.01707f
C335 B.n51 VSUBS 0.007623f
C336 B.n52 VSUBS 0.007623f
C337 B.n53 VSUBS 0.007623f
C338 B.n54 VSUBS 0.007623f
C339 B.n55 VSUBS 0.007623f
C340 B.n56 VSUBS 0.007623f
C341 B.n57 VSUBS 0.007623f
C342 B.n58 VSUBS 0.007623f
C343 B.n59 VSUBS 0.007623f
C344 B.n60 VSUBS 0.007623f
C345 B.n61 VSUBS 0.007623f
C346 B.n62 VSUBS 0.007623f
C347 B.n63 VSUBS 0.007623f
C348 B.n64 VSUBS 0.007623f
C349 B.n65 VSUBS 0.007623f
C350 B.n66 VSUBS 0.007623f
C351 B.n67 VSUBS 0.007623f
C352 B.n68 VSUBS 0.007623f
C353 B.n69 VSUBS 0.007623f
C354 B.n70 VSUBS 0.007623f
C355 B.n71 VSUBS 0.007623f
C356 B.n72 VSUBS 0.007623f
C357 B.n73 VSUBS 0.007623f
C358 B.n74 VSUBS 0.007623f
C359 B.n75 VSUBS 0.007623f
C360 B.n76 VSUBS 0.007623f
C361 B.n77 VSUBS 0.007623f
C362 B.n78 VSUBS 0.007623f
C363 B.n79 VSUBS 0.007623f
C364 B.n80 VSUBS 0.007623f
C365 B.n81 VSUBS 0.007623f
C366 B.n82 VSUBS 0.017119f
C367 B.n83 VSUBS 0.007623f
C368 B.n84 VSUBS 0.007623f
C369 B.n85 VSUBS 0.007623f
C370 B.n86 VSUBS 0.007623f
C371 B.n87 VSUBS 0.007623f
C372 B.n88 VSUBS 0.007623f
C373 B.n89 VSUBS 0.007623f
C374 B.n90 VSUBS 0.007623f
C375 B.n91 VSUBS 0.007623f
C376 B.n92 VSUBS 0.007623f
C377 B.n93 VSUBS 0.007623f
C378 B.n94 VSUBS 0.005269f
C379 B.n95 VSUBS 0.007623f
C380 B.n96 VSUBS 0.007623f
C381 B.n97 VSUBS 0.007623f
C382 B.n98 VSUBS 0.007623f
C383 B.n99 VSUBS 0.007623f
C384 B.t5 VSUBS 0.094501f
C385 B.t4 VSUBS 0.130673f
C386 B.t3 VSUBS 1.10947f
C387 B.n100 VSUBS 0.217472f
C388 B.n101 VSUBS 0.172396f
C389 B.n102 VSUBS 0.007623f
C390 B.n103 VSUBS 0.007623f
C391 B.n104 VSUBS 0.007623f
C392 B.n105 VSUBS 0.007623f
C393 B.n106 VSUBS 0.007623f
C394 B.n107 VSUBS 0.007623f
C395 B.n108 VSUBS 0.007623f
C396 B.n109 VSUBS 0.007623f
C397 B.n110 VSUBS 0.007623f
C398 B.n111 VSUBS 0.007623f
C399 B.n112 VSUBS 0.007623f
C400 B.n113 VSUBS 0.016111f
C401 B.n114 VSUBS 0.007623f
C402 B.n115 VSUBS 0.007623f
C403 B.n116 VSUBS 0.007623f
C404 B.n117 VSUBS 0.007623f
C405 B.n118 VSUBS 0.007623f
C406 B.n119 VSUBS 0.007623f
C407 B.n120 VSUBS 0.007623f
C408 B.n121 VSUBS 0.007623f
C409 B.n122 VSUBS 0.007623f
C410 B.n123 VSUBS 0.007623f
C411 B.n124 VSUBS 0.007623f
C412 B.n125 VSUBS 0.007623f
C413 B.n126 VSUBS 0.007623f
C414 B.n127 VSUBS 0.007623f
C415 B.n128 VSUBS 0.007623f
C416 B.n129 VSUBS 0.007623f
C417 B.n130 VSUBS 0.007623f
C418 B.n131 VSUBS 0.007623f
C419 B.n132 VSUBS 0.007623f
C420 B.n133 VSUBS 0.007623f
C421 B.n134 VSUBS 0.007623f
C422 B.n135 VSUBS 0.007623f
C423 B.n136 VSUBS 0.007623f
C424 B.n137 VSUBS 0.007623f
C425 B.n138 VSUBS 0.007623f
C426 B.n139 VSUBS 0.007623f
C427 B.n140 VSUBS 0.007623f
C428 B.n141 VSUBS 0.007623f
C429 B.n142 VSUBS 0.007623f
C430 B.n143 VSUBS 0.007623f
C431 B.n144 VSUBS 0.007623f
C432 B.n145 VSUBS 0.007623f
C433 B.n146 VSUBS 0.007623f
C434 B.n147 VSUBS 0.007623f
C435 B.n148 VSUBS 0.007623f
C436 B.n149 VSUBS 0.007623f
C437 B.n150 VSUBS 0.007623f
C438 B.n151 VSUBS 0.007623f
C439 B.n152 VSUBS 0.007623f
C440 B.n153 VSUBS 0.007623f
C441 B.n154 VSUBS 0.007623f
C442 B.n155 VSUBS 0.007623f
C443 B.n156 VSUBS 0.007623f
C444 B.n157 VSUBS 0.007623f
C445 B.n158 VSUBS 0.007623f
C446 B.n159 VSUBS 0.007623f
C447 B.n160 VSUBS 0.007623f
C448 B.n161 VSUBS 0.007623f
C449 B.n162 VSUBS 0.007623f
C450 B.n163 VSUBS 0.007623f
C451 B.n164 VSUBS 0.007623f
C452 B.n165 VSUBS 0.007623f
C453 B.n166 VSUBS 0.007623f
C454 B.n167 VSUBS 0.007623f
C455 B.n168 VSUBS 0.007623f
C456 B.n169 VSUBS 0.007623f
C457 B.n170 VSUBS 0.007623f
C458 B.n171 VSUBS 0.007623f
C459 B.n172 VSUBS 0.016111f
C460 B.n173 VSUBS 0.01707f
C461 B.n174 VSUBS 0.01707f
C462 B.n175 VSUBS 0.007623f
C463 B.n176 VSUBS 0.007623f
C464 B.n177 VSUBS 0.007623f
C465 B.n178 VSUBS 0.007623f
C466 B.n179 VSUBS 0.007623f
C467 B.n180 VSUBS 0.007623f
C468 B.n181 VSUBS 0.007623f
C469 B.n182 VSUBS 0.007623f
C470 B.n183 VSUBS 0.007623f
C471 B.n184 VSUBS 0.007623f
C472 B.n185 VSUBS 0.007623f
C473 B.n186 VSUBS 0.007623f
C474 B.n187 VSUBS 0.007623f
C475 B.n188 VSUBS 0.007623f
C476 B.n189 VSUBS 0.007623f
C477 B.n190 VSUBS 0.007623f
C478 B.n191 VSUBS 0.007623f
C479 B.n192 VSUBS 0.007623f
C480 B.n193 VSUBS 0.007623f
C481 B.n194 VSUBS 0.007623f
C482 B.n195 VSUBS 0.007623f
C483 B.n196 VSUBS 0.007623f
C484 B.n197 VSUBS 0.007623f
C485 B.n198 VSUBS 0.007623f
C486 B.n199 VSUBS 0.007623f
C487 B.n200 VSUBS 0.007623f
C488 B.n201 VSUBS 0.007623f
C489 B.n202 VSUBS 0.007623f
C490 B.n203 VSUBS 0.007623f
C491 B.n204 VSUBS 0.007623f
C492 B.n205 VSUBS 0.007623f
C493 B.n206 VSUBS 0.007623f
C494 B.n207 VSUBS 0.007623f
C495 B.n208 VSUBS 0.005269f
C496 B.n209 VSUBS 0.017661f
C497 B.n210 VSUBS 0.006165f
C498 B.n211 VSUBS 0.007623f
C499 B.n212 VSUBS 0.007623f
C500 B.n213 VSUBS 0.007623f
C501 B.n214 VSUBS 0.007623f
C502 B.n215 VSUBS 0.007623f
C503 B.n216 VSUBS 0.007623f
C504 B.n217 VSUBS 0.007623f
C505 B.n218 VSUBS 0.007623f
C506 B.n219 VSUBS 0.007623f
C507 B.n220 VSUBS 0.007623f
C508 B.n221 VSUBS 0.007623f
C509 B.t8 VSUBS 0.094503f
C510 B.t7 VSUBS 0.130674f
C511 B.t6 VSUBS 1.10947f
C512 B.n222 VSUBS 0.21747f
C513 B.n223 VSUBS 0.172394f
C514 B.n224 VSUBS 0.017661f
C515 B.n225 VSUBS 0.006165f
C516 B.n226 VSUBS 0.007623f
C517 B.n227 VSUBS 0.007623f
C518 B.n228 VSUBS 0.007623f
C519 B.n229 VSUBS 0.007623f
C520 B.n230 VSUBS 0.007623f
C521 B.n231 VSUBS 0.007623f
C522 B.n232 VSUBS 0.007623f
C523 B.n233 VSUBS 0.007623f
C524 B.n234 VSUBS 0.007623f
C525 B.n235 VSUBS 0.007623f
C526 B.n236 VSUBS 0.007623f
C527 B.n237 VSUBS 0.007623f
C528 B.n238 VSUBS 0.007623f
C529 B.n239 VSUBS 0.007623f
C530 B.n240 VSUBS 0.007623f
C531 B.n241 VSUBS 0.007623f
C532 B.n242 VSUBS 0.007623f
C533 B.n243 VSUBS 0.007623f
C534 B.n244 VSUBS 0.007623f
C535 B.n245 VSUBS 0.007623f
C536 B.n246 VSUBS 0.007623f
C537 B.n247 VSUBS 0.007623f
C538 B.n248 VSUBS 0.007623f
C539 B.n249 VSUBS 0.007623f
C540 B.n250 VSUBS 0.007623f
C541 B.n251 VSUBS 0.007623f
C542 B.n252 VSUBS 0.007623f
C543 B.n253 VSUBS 0.007623f
C544 B.n254 VSUBS 0.007623f
C545 B.n255 VSUBS 0.007623f
C546 B.n256 VSUBS 0.007623f
C547 B.n257 VSUBS 0.007623f
C548 B.n258 VSUBS 0.007623f
C549 B.n259 VSUBS 0.007623f
C550 B.n260 VSUBS 0.007623f
C551 B.n261 VSUBS 0.016062f
C552 B.n262 VSUBS 0.01707f
C553 B.n263 VSUBS 0.016111f
C554 B.n264 VSUBS 0.007623f
C555 B.n265 VSUBS 0.007623f
C556 B.n266 VSUBS 0.007623f
C557 B.n267 VSUBS 0.007623f
C558 B.n268 VSUBS 0.007623f
C559 B.n269 VSUBS 0.007623f
C560 B.n270 VSUBS 0.007623f
C561 B.n271 VSUBS 0.007623f
C562 B.n272 VSUBS 0.007623f
C563 B.n273 VSUBS 0.007623f
C564 B.n274 VSUBS 0.007623f
C565 B.n275 VSUBS 0.007623f
C566 B.n276 VSUBS 0.007623f
C567 B.n277 VSUBS 0.007623f
C568 B.n278 VSUBS 0.007623f
C569 B.n279 VSUBS 0.007623f
C570 B.n280 VSUBS 0.007623f
C571 B.n281 VSUBS 0.007623f
C572 B.n282 VSUBS 0.007623f
C573 B.n283 VSUBS 0.007623f
C574 B.n284 VSUBS 0.007623f
C575 B.n285 VSUBS 0.007623f
C576 B.n286 VSUBS 0.007623f
C577 B.n287 VSUBS 0.007623f
C578 B.n288 VSUBS 0.007623f
C579 B.n289 VSUBS 0.007623f
C580 B.n290 VSUBS 0.007623f
C581 B.n291 VSUBS 0.007623f
C582 B.n292 VSUBS 0.007623f
C583 B.n293 VSUBS 0.007623f
C584 B.n294 VSUBS 0.007623f
C585 B.n295 VSUBS 0.007623f
C586 B.n296 VSUBS 0.007623f
C587 B.n297 VSUBS 0.007623f
C588 B.n298 VSUBS 0.007623f
C589 B.n299 VSUBS 0.007623f
C590 B.n300 VSUBS 0.007623f
C591 B.n301 VSUBS 0.007623f
C592 B.n302 VSUBS 0.007623f
C593 B.n303 VSUBS 0.007623f
C594 B.n304 VSUBS 0.007623f
C595 B.n305 VSUBS 0.007623f
C596 B.n306 VSUBS 0.007623f
C597 B.n307 VSUBS 0.007623f
C598 B.n308 VSUBS 0.007623f
C599 B.n309 VSUBS 0.007623f
C600 B.n310 VSUBS 0.007623f
C601 B.n311 VSUBS 0.007623f
C602 B.n312 VSUBS 0.007623f
C603 B.n313 VSUBS 0.007623f
C604 B.n314 VSUBS 0.007623f
C605 B.n315 VSUBS 0.007623f
C606 B.n316 VSUBS 0.007623f
C607 B.n317 VSUBS 0.007623f
C608 B.n318 VSUBS 0.007623f
C609 B.n319 VSUBS 0.007623f
C610 B.n320 VSUBS 0.007623f
C611 B.n321 VSUBS 0.007623f
C612 B.n322 VSUBS 0.007623f
C613 B.n323 VSUBS 0.007623f
C614 B.n324 VSUBS 0.007623f
C615 B.n325 VSUBS 0.007623f
C616 B.n326 VSUBS 0.007623f
C617 B.n327 VSUBS 0.007623f
C618 B.n328 VSUBS 0.007623f
C619 B.n329 VSUBS 0.007623f
C620 B.n330 VSUBS 0.007623f
C621 B.n331 VSUBS 0.007623f
C622 B.n332 VSUBS 0.007623f
C623 B.n333 VSUBS 0.007623f
C624 B.n334 VSUBS 0.007623f
C625 B.n335 VSUBS 0.007623f
C626 B.n336 VSUBS 0.007623f
C627 B.n337 VSUBS 0.007623f
C628 B.n338 VSUBS 0.007623f
C629 B.n339 VSUBS 0.007623f
C630 B.n340 VSUBS 0.007623f
C631 B.n341 VSUBS 0.007623f
C632 B.n342 VSUBS 0.007623f
C633 B.n343 VSUBS 0.007623f
C634 B.n344 VSUBS 0.007623f
C635 B.n345 VSUBS 0.007623f
C636 B.n346 VSUBS 0.007623f
C637 B.n347 VSUBS 0.007623f
C638 B.n348 VSUBS 0.007623f
C639 B.n349 VSUBS 0.007623f
C640 B.n350 VSUBS 0.007623f
C641 B.n351 VSUBS 0.007623f
C642 B.n352 VSUBS 0.007623f
C643 B.n353 VSUBS 0.007623f
C644 B.n354 VSUBS 0.007623f
C645 B.n355 VSUBS 0.007623f
C646 B.n356 VSUBS 0.007623f
C647 B.n357 VSUBS 0.016111f
C648 B.n358 VSUBS 0.016111f
C649 B.n359 VSUBS 0.01707f
C650 B.n360 VSUBS 0.007623f
C651 B.n361 VSUBS 0.007623f
C652 B.n362 VSUBS 0.007623f
C653 B.n363 VSUBS 0.007623f
C654 B.n364 VSUBS 0.007623f
C655 B.n365 VSUBS 0.007623f
C656 B.n366 VSUBS 0.007623f
C657 B.n367 VSUBS 0.007623f
C658 B.n368 VSUBS 0.007623f
C659 B.n369 VSUBS 0.007623f
C660 B.n370 VSUBS 0.007623f
C661 B.n371 VSUBS 0.007623f
C662 B.n372 VSUBS 0.007623f
C663 B.n373 VSUBS 0.007623f
C664 B.n374 VSUBS 0.007623f
C665 B.n375 VSUBS 0.007623f
C666 B.n376 VSUBS 0.007623f
C667 B.n377 VSUBS 0.007623f
C668 B.n378 VSUBS 0.007623f
C669 B.n379 VSUBS 0.007623f
C670 B.n380 VSUBS 0.007623f
C671 B.n381 VSUBS 0.007623f
C672 B.n382 VSUBS 0.007623f
C673 B.n383 VSUBS 0.007623f
C674 B.n384 VSUBS 0.007623f
C675 B.n385 VSUBS 0.007623f
C676 B.n386 VSUBS 0.007623f
C677 B.n387 VSUBS 0.007623f
C678 B.n388 VSUBS 0.007623f
C679 B.n389 VSUBS 0.007623f
C680 B.n390 VSUBS 0.007623f
C681 B.n391 VSUBS 0.007623f
C682 B.n392 VSUBS 0.007623f
C683 B.n393 VSUBS 0.005269f
C684 B.n394 VSUBS 0.007623f
C685 B.n395 VSUBS 0.007623f
C686 B.n396 VSUBS 0.006165f
C687 B.n397 VSUBS 0.007623f
C688 B.n398 VSUBS 0.007623f
C689 B.n399 VSUBS 0.007623f
C690 B.n400 VSUBS 0.007623f
C691 B.n401 VSUBS 0.007623f
C692 B.n402 VSUBS 0.007623f
C693 B.n403 VSUBS 0.007623f
C694 B.n404 VSUBS 0.007623f
C695 B.n405 VSUBS 0.007623f
C696 B.n406 VSUBS 0.007623f
C697 B.n407 VSUBS 0.007623f
C698 B.n408 VSUBS 0.006165f
C699 B.n409 VSUBS 0.017661f
C700 B.n410 VSUBS 0.005269f
C701 B.n411 VSUBS 0.007623f
C702 B.n412 VSUBS 0.007623f
C703 B.n413 VSUBS 0.007623f
C704 B.n414 VSUBS 0.007623f
C705 B.n415 VSUBS 0.007623f
C706 B.n416 VSUBS 0.007623f
C707 B.n417 VSUBS 0.007623f
C708 B.n418 VSUBS 0.007623f
C709 B.n419 VSUBS 0.007623f
C710 B.n420 VSUBS 0.007623f
C711 B.n421 VSUBS 0.007623f
C712 B.n422 VSUBS 0.007623f
C713 B.n423 VSUBS 0.007623f
C714 B.n424 VSUBS 0.007623f
C715 B.n425 VSUBS 0.007623f
C716 B.n426 VSUBS 0.007623f
C717 B.n427 VSUBS 0.007623f
C718 B.n428 VSUBS 0.007623f
C719 B.n429 VSUBS 0.007623f
C720 B.n430 VSUBS 0.007623f
C721 B.n431 VSUBS 0.007623f
C722 B.n432 VSUBS 0.007623f
C723 B.n433 VSUBS 0.007623f
C724 B.n434 VSUBS 0.007623f
C725 B.n435 VSUBS 0.007623f
C726 B.n436 VSUBS 0.007623f
C727 B.n437 VSUBS 0.007623f
C728 B.n438 VSUBS 0.007623f
C729 B.n439 VSUBS 0.007623f
C730 B.n440 VSUBS 0.007623f
C731 B.n441 VSUBS 0.007623f
C732 B.n442 VSUBS 0.007623f
C733 B.n443 VSUBS 0.007623f
C734 B.n444 VSUBS 0.01707f
C735 B.n445 VSUBS 0.01707f
C736 B.n446 VSUBS 0.016111f
C737 B.n447 VSUBS 0.007623f
C738 B.n448 VSUBS 0.007623f
C739 B.n449 VSUBS 0.007623f
C740 B.n450 VSUBS 0.007623f
C741 B.n451 VSUBS 0.007623f
C742 B.n452 VSUBS 0.007623f
C743 B.n453 VSUBS 0.007623f
C744 B.n454 VSUBS 0.007623f
C745 B.n455 VSUBS 0.007623f
C746 B.n456 VSUBS 0.007623f
C747 B.n457 VSUBS 0.007623f
C748 B.n458 VSUBS 0.007623f
C749 B.n459 VSUBS 0.007623f
C750 B.n460 VSUBS 0.007623f
C751 B.n461 VSUBS 0.007623f
C752 B.n462 VSUBS 0.007623f
C753 B.n463 VSUBS 0.007623f
C754 B.n464 VSUBS 0.007623f
C755 B.n465 VSUBS 0.007623f
C756 B.n466 VSUBS 0.007623f
C757 B.n467 VSUBS 0.007623f
C758 B.n468 VSUBS 0.007623f
C759 B.n469 VSUBS 0.007623f
C760 B.n470 VSUBS 0.007623f
C761 B.n471 VSUBS 0.007623f
C762 B.n472 VSUBS 0.007623f
C763 B.n473 VSUBS 0.007623f
C764 B.n474 VSUBS 0.007623f
C765 B.n475 VSUBS 0.007623f
C766 B.n476 VSUBS 0.007623f
C767 B.n477 VSUBS 0.007623f
C768 B.n478 VSUBS 0.007623f
C769 B.n479 VSUBS 0.007623f
C770 B.n480 VSUBS 0.007623f
C771 B.n481 VSUBS 0.007623f
C772 B.n482 VSUBS 0.007623f
C773 B.n483 VSUBS 0.007623f
C774 B.n484 VSUBS 0.007623f
C775 B.n485 VSUBS 0.007623f
C776 B.n486 VSUBS 0.007623f
C777 B.n487 VSUBS 0.007623f
C778 B.n488 VSUBS 0.007623f
C779 B.n489 VSUBS 0.007623f
C780 B.n490 VSUBS 0.007623f
C781 B.n491 VSUBS 0.009947f
C782 B.n492 VSUBS 0.010596f
C783 B.n493 VSUBS 0.021072f
.ends

