* NGSPICE file created from diff_pair_sample_1733.ext - technology: sky130A

.subckt diff_pair_sample_1733 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t7 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=5.3781 pd=28.36 as=2.27535 ps=14.12 w=13.79 l=2.39
X1 VDD2.t9 VN.t0 VTAIL.t6 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=2.27535 pd=14.12 as=2.27535 ps=14.12 w=13.79 l=2.39
X2 VTAIL.t19 VN.t1 VDD2.t8 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=2.27535 pd=14.12 as=2.27535 ps=14.12 w=13.79 l=2.39
X3 VDD1.t8 VP.t1 VTAIL.t12 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=2.27535 pd=14.12 as=5.3781 ps=28.36 w=13.79 l=2.39
X4 VTAIL.t9 VP.t2 VDD1.t7 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=2.27535 pd=14.12 as=2.27535 ps=14.12 w=13.79 l=2.39
X5 VTAIL.t8 VP.t3 VDD1.t6 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=2.27535 pd=14.12 as=2.27535 ps=14.12 w=13.79 l=2.39
X6 VDD2.t7 VN.t2 VTAIL.t1 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=2.27535 pd=14.12 as=2.27535 ps=14.12 w=13.79 l=2.39
X7 VDD2.t6 VN.t3 VTAIL.t3 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=5.3781 pd=28.36 as=2.27535 ps=14.12 w=13.79 l=2.39
X8 VTAIL.t4 VN.t4 VDD2.t5 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=2.27535 pd=14.12 as=2.27535 ps=14.12 w=13.79 l=2.39
X9 VTAIL.t5 VN.t5 VDD2.t4 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=2.27535 pd=14.12 as=2.27535 ps=14.12 w=13.79 l=2.39
X10 B.t11 B.t9 B.t10 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=5.3781 pd=28.36 as=0 ps=0 w=13.79 l=2.39
X11 VDD2.t3 VN.t6 VTAIL.t17 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=2.27535 pd=14.12 as=5.3781 ps=28.36 w=13.79 l=2.39
X12 VDD2.t2 VN.t7 VTAIL.t18 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=2.27535 pd=14.12 as=5.3781 ps=28.36 w=13.79 l=2.39
X13 VTAIL.t15 VP.t4 VDD1.t5 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=2.27535 pd=14.12 as=2.27535 ps=14.12 w=13.79 l=2.39
X14 VTAIL.t14 VP.t5 VDD1.t4 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=2.27535 pd=14.12 as=2.27535 ps=14.12 w=13.79 l=2.39
X15 VDD2.t1 VN.t8 VTAIL.t2 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=5.3781 pd=28.36 as=2.27535 ps=14.12 w=13.79 l=2.39
X16 VDD1.t3 VP.t6 VTAIL.t13 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=2.27535 pd=14.12 as=2.27535 ps=14.12 w=13.79 l=2.39
X17 B.t8 B.t6 B.t7 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=5.3781 pd=28.36 as=0 ps=0 w=13.79 l=2.39
X18 VDD1.t2 VP.t7 VTAIL.t16 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=2.27535 pd=14.12 as=5.3781 ps=28.36 w=13.79 l=2.39
X19 VTAIL.t0 VN.t9 VDD2.t0 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=2.27535 pd=14.12 as=2.27535 ps=14.12 w=13.79 l=2.39
X20 VDD1.t1 VP.t8 VTAIL.t10 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=5.3781 pd=28.36 as=2.27535 ps=14.12 w=13.79 l=2.39
X21 VDD1.t0 VP.t9 VTAIL.t11 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=2.27535 pd=14.12 as=2.27535 ps=14.12 w=13.79 l=2.39
X22 B.t5 B.t3 B.t4 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=5.3781 pd=28.36 as=0 ps=0 w=13.79 l=2.39
X23 B.t2 B.t0 B.t1 w_n4234_n3726# sky130_fd_pr__pfet_01v8 ad=5.3781 pd=28.36 as=0 ps=0 w=13.79 l=2.39
R0 VP.n21 VP.t0 172.46
R1 VP.n23 VP.n20 161.3
R2 VP.n25 VP.n24 161.3
R3 VP.n26 VP.n19 161.3
R4 VP.n28 VP.n27 161.3
R5 VP.n29 VP.n18 161.3
R6 VP.n32 VP.n31 161.3
R7 VP.n33 VP.n17 161.3
R8 VP.n35 VP.n34 161.3
R9 VP.n36 VP.n16 161.3
R10 VP.n38 VP.n37 161.3
R11 VP.n40 VP.n39 161.3
R12 VP.n41 VP.n14 161.3
R13 VP.n43 VP.n42 161.3
R14 VP.n44 VP.n13 161.3
R15 VP.n46 VP.n45 161.3
R16 VP.n47 VP.n12 161.3
R17 VP.n86 VP.n0 161.3
R18 VP.n85 VP.n84 161.3
R19 VP.n83 VP.n1 161.3
R20 VP.n82 VP.n81 161.3
R21 VP.n80 VP.n2 161.3
R22 VP.n79 VP.n78 161.3
R23 VP.n77 VP.n76 161.3
R24 VP.n75 VP.n4 161.3
R25 VP.n74 VP.n73 161.3
R26 VP.n72 VP.n5 161.3
R27 VP.n71 VP.n70 161.3
R28 VP.n68 VP.n6 161.3
R29 VP.n67 VP.n66 161.3
R30 VP.n65 VP.n7 161.3
R31 VP.n64 VP.n63 161.3
R32 VP.n62 VP.n8 161.3
R33 VP.n60 VP.n59 161.3
R34 VP.n58 VP.n9 161.3
R35 VP.n57 VP.n56 161.3
R36 VP.n55 VP.n10 161.3
R37 VP.n54 VP.n53 161.3
R38 VP.n52 VP.n11 161.3
R39 VP.n50 VP.t8 139.054
R40 VP.n61 VP.t2 139.054
R41 VP.n69 VP.t9 139.054
R42 VP.n3 VP.t4 139.054
R43 VP.n87 VP.t1 139.054
R44 VP.n48 VP.t7 139.054
R45 VP.n15 VP.t5 139.054
R46 VP.n30 VP.t6 139.054
R47 VP.n22 VP.t3 139.054
R48 VP.n51 VP.n50 101.459
R49 VP.n88 VP.n87 101.459
R50 VP.n49 VP.n48 101.459
R51 VP.n56 VP.n55 56.5193
R52 VP.n81 VP.n1 56.5193
R53 VP.n42 VP.n13 56.5193
R54 VP.n51 VP.n49 53.2875
R55 VP.n63 VP.n7 51.1773
R56 VP.n75 VP.n74 51.1773
R57 VP.n36 VP.n35 51.1773
R58 VP.n24 VP.n19 51.1773
R59 VP.n22 VP.n21 49.4099
R60 VP.n67 VP.n7 29.8095
R61 VP.n74 VP.n5 29.8095
R62 VP.n35 VP.n17 29.8095
R63 VP.n28 VP.n19 29.8095
R64 VP.n54 VP.n11 24.4675
R65 VP.n55 VP.n54 24.4675
R66 VP.n56 VP.n9 24.4675
R67 VP.n60 VP.n9 24.4675
R68 VP.n63 VP.n62 24.4675
R69 VP.n68 VP.n67 24.4675
R70 VP.n70 VP.n5 24.4675
R71 VP.n76 VP.n75 24.4675
R72 VP.n80 VP.n79 24.4675
R73 VP.n81 VP.n80 24.4675
R74 VP.n85 VP.n1 24.4675
R75 VP.n86 VP.n85 24.4675
R76 VP.n46 VP.n13 24.4675
R77 VP.n47 VP.n46 24.4675
R78 VP.n37 VP.n36 24.4675
R79 VP.n41 VP.n40 24.4675
R80 VP.n42 VP.n41 24.4675
R81 VP.n29 VP.n28 24.4675
R82 VP.n31 VP.n17 24.4675
R83 VP.n24 VP.n23 24.4675
R84 VP.n62 VP.n61 22.9995
R85 VP.n76 VP.n3 22.9995
R86 VP.n37 VP.n15 22.9995
R87 VP.n23 VP.n22 22.9995
R88 VP.n69 VP.n68 12.234
R89 VP.n70 VP.n69 12.234
R90 VP.n30 VP.n29 12.234
R91 VP.n31 VP.n30 12.234
R92 VP.n50 VP.n11 9.29796
R93 VP.n87 VP.n86 9.29796
R94 VP.n48 VP.n47 9.29796
R95 VP.n21 VP.n20 6.89416
R96 VP.n61 VP.n60 1.46852
R97 VP.n79 VP.n3 1.46852
R98 VP.n40 VP.n15 1.46852
R99 VP.n49 VP.n12 0.278367
R100 VP.n52 VP.n51 0.278367
R101 VP.n88 VP.n0 0.278367
R102 VP.n25 VP.n20 0.189894
R103 VP.n26 VP.n25 0.189894
R104 VP.n27 VP.n26 0.189894
R105 VP.n27 VP.n18 0.189894
R106 VP.n32 VP.n18 0.189894
R107 VP.n33 VP.n32 0.189894
R108 VP.n34 VP.n33 0.189894
R109 VP.n34 VP.n16 0.189894
R110 VP.n38 VP.n16 0.189894
R111 VP.n39 VP.n38 0.189894
R112 VP.n39 VP.n14 0.189894
R113 VP.n43 VP.n14 0.189894
R114 VP.n44 VP.n43 0.189894
R115 VP.n45 VP.n44 0.189894
R116 VP.n45 VP.n12 0.189894
R117 VP.n53 VP.n52 0.189894
R118 VP.n53 VP.n10 0.189894
R119 VP.n57 VP.n10 0.189894
R120 VP.n58 VP.n57 0.189894
R121 VP.n59 VP.n58 0.189894
R122 VP.n59 VP.n8 0.189894
R123 VP.n64 VP.n8 0.189894
R124 VP.n65 VP.n64 0.189894
R125 VP.n66 VP.n65 0.189894
R126 VP.n66 VP.n6 0.189894
R127 VP.n71 VP.n6 0.189894
R128 VP.n72 VP.n71 0.189894
R129 VP.n73 VP.n72 0.189894
R130 VP.n73 VP.n4 0.189894
R131 VP.n77 VP.n4 0.189894
R132 VP.n78 VP.n77 0.189894
R133 VP.n78 VP.n2 0.189894
R134 VP.n82 VP.n2 0.189894
R135 VP.n83 VP.n82 0.189894
R136 VP.n84 VP.n83 0.189894
R137 VP.n84 VP.n0 0.189894
R138 VP VP.n88 0.153454
R139 VTAIL.n11 VTAIL.t17 61.782
R140 VTAIL.n17 VTAIL.t18 61.7818
R141 VTAIL.n2 VTAIL.t12 61.7818
R142 VTAIL.n16 VTAIL.t16 61.7818
R143 VTAIL.n15 VTAIL.n14 59.4248
R144 VTAIL.n13 VTAIL.n12 59.4248
R145 VTAIL.n10 VTAIL.n9 59.4248
R146 VTAIL.n8 VTAIL.n7 59.4248
R147 VTAIL.n19 VTAIL.n18 59.4246
R148 VTAIL.n1 VTAIL.n0 59.4246
R149 VTAIL.n4 VTAIL.n3 59.4246
R150 VTAIL.n6 VTAIL.n5 59.4246
R151 VTAIL.n8 VTAIL.n6 28.9445
R152 VTAIL.n17 VTAIL.n16 26.5996
R153 VTAIL.n18 VTAIL.t6 2.35764
R154 VTAIL.n18 VTAIL.t19 2.35764
R155 VTAIL.n0 VTAIL.t3 2.35764
R156 VTAIL.n0 VTAIL.t4 2.35764
R157 VTAIL.n3 VTAIL.t11 2.35764
R158 VTAIL.n3 VTAIL.t15 2.35764
R159 VTAIL.n5 VTAIL.t10 2.35764
R160 VTAIL.n5 VTAIL.t9 2.35764
R161 VTAIL.n14 VTAIL.t13 2.35764
R162 VTAIL.n14 VTAIL.t14 2.35764
R163 VTAIL.n12 VTAIL.t7 2.35764
R164 VTAIL.n12 VTAIL.t8 2.35764
R165 VTAIL.n9 VTAIL.t1 2.35764
R166 VTAIL.n9 VTAIL.t0 2.35764
R167 VTAIL.n7 VTAIL.t2 2.35764
R168 VTAIL.n7 VTAIL.t5 2.35764
R169 VTAIL.n10 VTAIL.n8 2.34533
R170 VTAIL.n11 VTAIL.n10 2.34533
R171 VTAIL.n15 VTAIL.n13 2.34533
R172 VTAIL.n16 VTAIL.n15 2.34533
R173 VTAIL.n6 VTAIL.n4 2.34533
R174 VTAIL.n4 VTAIL.n2 2.34533
R175 VTAIL.n19 VTAIL.n17 2.34533
R176 VTAIL VTAIL.n1 1.81731
R177 VTAIL.n13 VTAIL.n11 1.64274
R178 VTAIL.n2 VTAIL.n1 1.64274
R179 VTAIL VTAIL.n19 0.528517
R180 VDD1.n1 VDD1.t9 80.8056
R181 VDD1.n3 VDD1.t1 80.8054
R182 VDD1.n5 VDD1.n4 77.8067
R183 VDD1.n1 VDD1.n0 76.1036
R184 VDD1.n7 VDD1.n6 76.1035
R185 VDD1.n3 VDD1.n2 76.1034
R186 VDD1.n7 VDD1.n5 48.4966
R187 VDD1.n6 VDD1.t4 2.35764
R188 VDD1.n6 VDD1.t2 2.35764
R189 VDD1.n0 VDD1.t6 2.35764
R190 VDD1.n0 VDD1.t3 2.35764
R191 VDD1.n4 VDD1.t5 2.35764
R192 VDD1.n4 VDD1.t8 2.35764
R193 VDD1.n2 VDD1.t7 2.35764
R194 VDD1.n2 VDD1.t0 2.35764
R195 VDD1 VDD1.n7 1.70093
R196 VDD1 VDD1.n1 0.644897
R197 VDD1.n5 VDD1.n3 0.531361
R198 VN.n9 VN.t3 172.46
R199 VN.n47 VN.t6 172.46
R200 VN.n73 VN.n38 161.3
R201 VN.n72 VN.n71 161.3
R202 VN.n70 VN.n39 161.3
R203 VN.n69 VN.n68 161.3
R204 VN.n67 VN.n40 161.3
R205 VN.n66 VN.n65 161.3
R206 VN.n64 VN.n63 161.3
R207 VN.n62 VN.n42 161.3
R208 VN.n61 VN.n60 161.3
R209 VN.n59 VN.n43 161.3
R210 VN.n58 VN.n57 161.3
R211 VN.n55 VN.n44 161.3
R212 VN.n54 VN.n53 161.3
R213 VN.n52 VN.n45 161.3
R214 VN.n51 VN.n50 161.3
R215 VN.n49 VN.n46 161.3
R216 VN.n35 VN.n0 161.3
R217 VN.n34 VN.n33 161.3
R218 VN.n32 VN.n1 161.3
R219 VN.n31 VN.n30 161.3
R220 VN.n29 VN.n2 161.3
R221 VN.n28 VN.n27 161.3
R222 VN.n26 VN.n25 161.3
R223 VN.n24 VN.n4 161.3
R224 VN.n23 VN.n22 161.3
R225 VN.n21 VN.n5 161.3
R226 VN.n20 VN.n19 161.3
R227 VN.n17 VN.n6 161.3
R228 VN.n16 VN.n15 161.3
R229 VN.n14 VN.n7 161.3
R230 VN.n13 VN.n12 161.3
R231 VN.n11 VN.n8 161.3
R232 VN.n10 VN.t4 139.054
R233 VN.n18 VN.t0 139.054
R234 VN.n3 VN.t1 139.054
R235 VN.n36 VN.t7 139.054
R236 VN.n48 VN.t9 139.054
R237 VN.n56 VN.t2 139.054
R238 VN.n41 VN.t5 139.054
R239 VN.n74 VN.t8 139.054
R240 VN.n37 VN.n36 101.459
R241 VN.n75 VN.n74 101.459
R242 VN.n30 VN.n1 56.5193
R243 VN.n68 VN.n39 56.5193
R244 VN VN.n75 53.5663
R245 VN.n12 VN.n7 51.1773
R246 VN.n24 VN.n23 51.1773
R247 VN.n50 VN.n45 51.1773
R248 VN.n62 VN.n61 51.1773
R249 VN.n10 VN.n9 49.4099
R250 VN.n48 VN.n47 49.4099
R251 VN.n16 VN.n7 29.8095
R252 VN.n23 VN.n5 29.8095
R253 VN.n54 VN.n45 29.8095
R254 VN.n61 VN.n43 29.8095
R255 VN.n12 VN.n11 24.4675
R256 VN.n17 VN.n16 24.4675
R257 VN.n19 VN.n5 24.4675
R258 VN.n25 VN.n24 24.4675
R259 VN.n29 VN.n28 24.4675
R260 VN.n30 VN.n29 24.4675
R261 VN.n34 VN.n1 24.4675
R262 VN.n35 VN.n34 24.4675
R263 VN.n50 VN.n49 24.4675
R264 VN.n57 VN.n43 24.4675
R265 VN.n55 VN.n54 24.4675
R266 VN.n68 VN.n67 24.4675
R267 VN.n67 VN.n66 24.4675
R268 VN.n63 VN.n62 24.4675
R269 VN.n73 VN.n72 24.4675
R270 VN.n72 VN.n39 24.4675
R271 VN.n11 VN.n10 22.9995
R272 VN.n25 VN.n3 22.9995
R273 VN.n49 VN.n48 22.9995
R274 VN.n63 VN.n41 22.9995
R275 VN.n18 VN.n17 12.234
R276 VN.n19 VN.n18 12.234
R277 VN.n57 VN.n56 12.234
R278 VN.n56 VN.n55 12.234
R279 VN.n36 VN.n35 9.29796
R280 VN.n74 VN.n73 9.29796
R281 VN.n47 VN.n46 6.89416
R282 VN.n9 VN.n8 6.89416
R283 VN.n28 VN.n3 1.46852
R284 VN.n66 VN.n41 1.46852
R285 VN.n75 VN.n38 0.278367
R286 VN.n37 VN.n0 0.278367
R287 VN.n71 VN.n38 0.189894
R288 VN.n71 VN.n70 0.189894
R289 VN.n70 VN.n69 0.189894
R290 VN.n69 VN.n40 0.189894
R291 VN.n65 VN.n40 0.189894
R292 VN.n65 VN.n64 0.189894
R293 VN.n64 VN.n42 0.189894
R294 VN.n60 VN.n42 0.189894
R295 VN.n60 VN.n59 0.189894
R296 VN.n59 VN.n58 0.189894
R297 VN.n58 VN.n44 0.189894
R298 VN.n53 VN.n44 0.189894
R299 VN.n53 VN.n52 0.189894
R300 VN.n52 VN.n51 0.189894
R301 VN.n51 VN.n46 0.189894
R302 VN.n13 VN.n8 0.189894
R303 VN.n14 VN.n13 0.189894
R304 VN.n15 VN.n14 0.189894
R305 VN.n15 VN.n6 0.189894
R306 VN.n20 VN.n6 0.189894
R307 VN.n21 VN.n20 0.189894
R308 VN.n22 VN.n21 0.189894
R309 VN.n22 VN.n4 0.189894
R310 VN.n26 VN.n4 0.189894
R311 VN.n27 VN.n26 0.189894
R312 VN.n27 VN.n2 0.189894
R313 VN.n31 VN.n2 0.189894
R314 VN.n32 VN.n31 0.189894
R315 VN.n33 VN.n32 0.189894
R316 VN.n33 VN.n0 0.189894
R317 VN VN.n37 0.153454
R318 VDD2.n1 VDD2.t6 80.8054
R319 VDD2.n4 VDD2.t1 78.4608
R320 VDD2.n3 VDD2.n2 77.8067
R321 VDD2 VDD2.n7 77.8039
R322 VDD2.n6 VDD2.n5 76.1036
R323 VDD2.n1 VDD2.n0 76.1034
R324 VDD2.n4 VDD2.n3 46.7412
R325 VDD2.n7 VDD2.t0 2.35764
R326 VDD2.n7 VDD2.t3 2.35764
R327 VDD2.n5 VDD2.t4 2.35764
R328 VDD2.n5 VDD2.t7 2.35764
R329 VDD2.n2 VDD2.t8 2.35764
R330 VDD2.n2 VDD2.t2 2.35764
R331 VDD2.n0 VDD2.t5 2.35764
R332 VDD2.n0 VDD2.t9 2.35764
R333 VDD2.n6 VDD2.n4 2.34533
R334 VDD2 VDD2.n6 0.644897
R335 VDD2.n3 VDD2.n1 0.531361
R336 B.n635 B.n634 585
R337 B.n636 B.n85 585
R338 B.n638 B.n637 585
R339 B.n639 B.n84 585
R340 B.n641 B.n640 585
R341 B.n642 B.n83 585
R342 B.n644 B.n643 585
R343 B.n645 B.n82 585
R344 B.n647 B.n646 585
R345 B.n648 B.n81 585
R346 B.n650 B.n649 585
R347 B.n651 B.n80 585
R348 B.n653 B.n652 585
R349 B.n654 B.n79 585
R350 B.n656 B.n655 585
R351 B.n657 B.n78 585
R352 B.n659 B.n658 585
R353 B.n660 B.n77 585
R354 B.n662 B.n661 585
R355 B.n663 B.n76 585
R356 B.n665 B.n664 585
R357 B.n666 B.n75 585
R358 B.n668 B.n667 585
R359 B.n669 B.n74 585
R360 B.n671 B.n670 585
R361 B.n672 B.n73 585
R362 B.n674 B.n673 585
R363 B.n675 B.n72 585
R364 B.n677 B.n676 585
R365 B.n678 B.n71 585
R366 B.n680 B.n679 585
R367 B.n681 B.n70 585
R368 B.n683 B.n682 585
R369 B.n684 B.n69 585
R370 B.n686 B.n685 585
R371 B.n687 B.n68 585
R372 B.n689 B.n688 585
R373 B.n690 B.n67 585
R374 B.n692 B.n691 585
R375 B.n693 B.n66 585
R376 B.n695 B.n694 585
R377 B.n696 B.n65 585
R378 B.n698 B.n697 585
R379 B.n699 B.n64 585
R380 B.n701 B.n700 585
R381 B.n702 B.n63 585
R382 B.n704 B.n703 585
R383 B.n706 B.n705 585
R384 B.n707 B.n59 585
R385 B.n709 B.n708 585
R386 B.n710 B.n58 585
R387 B.n712 B.n711 585
R388 B.n713 B.n57 585
R389 B.n715 B.n714 585
R390 B.n716 B.n56 585
R391 B.n718 B.n717 585
R392 B.n720 B.n53 585
R393 B.n722 B.n721 585
R394 B.n723 B.n52 585
R395 B.n725 B.n724 585
R396 B.n726 B.n51 585
R397 B.n728 B.n727 585
R398 B.n729 B.n50 585
R399 B.n731 B.n730 585
R400 B.n732 B.n49 585
R401 B.n734 B.n733 585
R402 B.n735 B.n48 585
R403 B.n737 B.n736 585
R404 B.n738 B.n47 585
R405 B.n740 B.n739 585
R406 B.n741 B.n46 585
R407 B.n743 B.n742 585
R408 B.n744 B.n45 585
R409 B.n746 B.n745 585
R410 B.n747 B.n44 585
R411 B.n749 B.n748 585
R412 B.n750 B.n43 585
R413 B.n752 B.n751 585
R414 B.n753 B.n42 585
R415 B.n755 B.n754 585
R416 B.n756 B.n41 585
R417 B.n758 B.n757 585
R418 B.n759 B.n40 585
R419 B.n761 B.n760 585
R420 B.n762 B.n39 585
R421 B.n764 B.n763 585
R422 B.n765 B.n38 585
R423 B.n767 B.n766 585
R424 B.n768 B.n37 585
R425 B.n770 B.n769 585
R426 B.n771 B.n36 585
R427 B.n773 B.n772 585
R428 B.n774 B.n35 585
R429 B.n776 B.n775 585
R430 B.n777 B.n34 585
R431 B.n779 B.n778 585
R432 B.n780 B.n33 585
R433 B.n782 B.n781 585
R434 B.n783 B.n32 585
R435 B.n785 B.n784 585
R436 B.n786 B.n31 585
R437 B.n788 B.n787 585
R438 B.n789 B.n30 585
R439 B.n633 B.n86 585
R440 B.n632 B.n631 585
R441 B.n630 B.n87 585
R442 B.n629 B.n628 585
R443 B.n627 B.n88 585
R444 B.n626 B.n625 585
R445 B.n624 B.n89 585
R446 B.n623 B.n622 585
R447 B.n621 B.n90 585
R448 B.n620 B.n619 585
R449 B.n618 B.n91 585
R450 B.n617 B.n616 585
R451 B.n615 B.n92 585
R452 B.n614 B.n613 585
R453 B.n612 B.n93 585
R454 B.n611 B.n610 585
R455 B.n609 B.n94 585
R456 B.n608 B.n607 585
R457 B.n606 B.n95 585
R458 B.n605 B.n604 585
R459 B.n603 B.n96 585
R460 B.n602 B.n601 585
R461 B.n600 B.n97 585
R462 B.n599 B.n598 585
R463 B.n597 B.n98 585
R464 B.n596 B.n595 585
R465 B.n594 B.n99 585
R466 B.n593 B.n592 585
R467 B.n591 B.n100 585
R468 B.n590 B.n589 585
R469 B.n588 B.n101 585
R470 B.n587 B.n586 585
R471 B.n585 B.n102 585
R472 B.n584 B.n583 585
R473 B.n582 B.n103 585
R474 B.n581 B.n580 585
R475 B.n579 B.n104 585
R476 B.n578 B.n577 585
R477 B.n576 B.n105 585
R478 B.n575 B.n574 585
R479 B.n573 B.n106 585
R480 B.n572 B.n571 585
R481 B.n570 B.n107 585
R482 B.n569 B.n568 585
R483 B.n567 B.n108 585
R484 B.n566 B.n565 585
R485 B.n564 B.n109 585
R486 B.n563 B.n562 585
R487 B.n561 B.n110 585
R488 B.n560 B.n559 585
R489 B.n558 B.n111 585
R490 B.n557 B.n556 585
R491 B.n555 B.n112 585
R492 B.n554 B.n553 585
R493 B.n552 B.n113 585
R494 B.n551 B.n550 585
R495 B.n549 B.n114 585
R496 B.n548 B.n547 585
R497 B.n546 B.n115 585
R498 B.n545 B.n544 585
R499 B.n543 B.n116 585
R500 B.n542 B.n541 585
R501 B.n540 B.n117 585
R502 B.n539 B.n538 585
R503 B.n537 B.n118 585
R504 B.n536 B.n535 585
R505 B.n534 B.n119 585
R506 B.n533 B.n532 585
R507 B.n531 B.n120 585
R508 B.n530 B.n529 585
R509 B.n528 B.n121 585
R510 B.n527 B.n526 585
R511 B.n525 B.n122 585
R512 B.n524 B.n523 585
R513 B.n522 B.n123 585
R514 B.n521 B.n520 585
R515 B.n519 B.n124 585
R516 B.n518 B.n517 585
R517 B.n516 B.n125 585
R518 B.n515 B.n514 585
R519 B.n513 B.n126 585
R520 B.n512 B.n511 585
R521 B.n510 B.n127 585
R522 B.n509 B.n508 585
R523 B.n507 B.n128 585
R524 B.n506 B.n505 585
R525 B.n504 B.n129 585
R526 B.n503 B.n502 585
R527 B.n501 B.n130 585
R528 B.n500 B.n499 585
R529 B.n498 B.n131 585
R530 B.n497 B.n496 585
R531 B.n495 B.n132 585
R532 B.n494 B.n493 585
R533 B.n492 B.n133 585
R534 B.n491 B.n490 585
R535 B.n489 B.n134 585
R536 B.n488 B.n487 585
R537 B.n486 B.n135 585
R538 B.n485 B.n484 585
R539 B.n483 B.n136 585
R540 B.n482 B.n481 585
R541 B.n480 B.n137 585
R542 B.n479 B.n478 585
R543 B.n477 B.n138 585
R544 B.n476 B.n475 585
R545 B.n474 B.n139 585
R546 B.n473 B.n472 585
R547 B.n471 B.n140 585
R548 B.n470 B.n469 585
R549 B.n468 B.n141 585
R550 B.n467 B.n466 585
R551 B.n465 B.n142 585
R552 B.n309 B.n198 585
R553 B.n311 B.n310 585
R554 B.n312 B.n197 585
R555 B.n314 B.n313 585
R556 B.n315 B.n196 585
R557 B.n317 B.n316 585
R558 B.n318 B.n195 585
R559 B.n320 B.n319 585
R560 B.n321 B.n194 585
R561 B.n323 B.n322 585
R562 B.n324 B.n193 585
R563 B.n326 B.n325 585
R564 B.n327 B.n192 585
R565 B.n329 B.n328 585
R566 B.n330 B.n191 585
R567 B.n332 B.n331 585
R568 B.n333 B.n190 585
R569 B.n335 B.n334 585
R570 B.n336 B.n189 585
R571 B.n338 B.n337 585
R572 B.n339 B.n188 585
R573 B.n341 B.n340 585
R574 B.n342 B.n187 585
R575 B.n344 B.n343 585
R576 B.n345 B.n186 585
R577 B.n347 B.n346 585
R578 B.n348 B.n185 585
R579 B.n350 B.n349 585
R580 B.n351 B.n184 585
R581 B.n353 B.n352 585
R582 B.n354 B.n183 585
R583 B.n356 B.n355 585
R584 B.n357 B.n182 585
R585 B.n359 B.n358 585
R586 B.n360 B.n181 585
R587 B.n362 B.n361 585
R588 B.n363 B.n180 585
R589 B.n365 B.n364 585
R590 B.n366 B.n179 585
R591 B.n368 B.n367 585
R592 B.n369 B.n178 585
R593 B.n371 B.n370 585
R594 B.n372 B.n177 585
R595 B.n374 B.n373 585
R596 B.n375 B.n176 585
R597 B.n377 B.n376 585
R598 B.n378 B.n173 585
R599 B.n381 B.n380 585
R600 B.n382 B.n172 585
R601 B.n384 B.n383 585
R602 B.n385 B.n171 585
R603 B.n387 B.n386 585
R604 B.n388 B.n170 585
R605 B.n390 B.n389 585
R606 B.n391 B.n169 585
R607 B.n393 B.n392 585
R608 B.n395 B.n394 585
R609 B.n396 B.n165 585
R610 B.n398 B.n397 585
R611 B.n399 B.n164 585
R612 B.n401 B.n400 585
R613 B.n402 B.n163 585
R614 B.n404 B.n403 585
R615 B.n405 B.n162 585
R616 B.n407 B.n406 585
R617 B.n408 B.n161 585
R618 B.n410 B.n409 585
R619 B.n411 B.n160 585
R620 B.n413 B.n412 585
R621 B.n414 B.n159 585
R622 B.n416 B.n415 585
R623 B.n417 B.n158 585
R624 B.n419 B.n418 585
R625 B.n420 B.n157 585
R626 B.n422 B.n421 585
R627 B.n423 B.n156 585
R628 B.n425 B.n424 585
R629 B.n426 B.n155 585
R630 B.n428 B.n427 585
R631 B.n429 B.n154 585
R632 B.n431 B.n430 585
R633 B.n432 B.n153 585
R634 B.n434 B.n433 585
R635 B.n435 B.n152 585
R636 B.n437 B.n436 585
R637 B.n438 B.n151 585
R638 B.n440 B.n439 585
R639 B.n441 B.n150 585
R640 B.n443 B.n442 585
R641 B.n444 B.n149 585
R642 B.n446 B.n445 585
R643 B.n447 B.n148 585
R644 B.n449 B.n448 585
R645 B.n450 B.n147 585
R646 B.n452 B.n451 585
R647 B.n453 B.n146 585
R648 B.n455 B.n454 585
R649 B.n456 B.n145 585
R650 B.n458 B.n457 585
R651 B.n459 B.n144 585
R652 B.n461 B.n460 585
R653 B.n462 B.n143 585
R654 B.n464 B.n463 585
R655 B.n308 B.n307 585
R656 B.n306 B.n199 585
R657 B.n305 B.n304 585
R658 B.n303 B.n200 585
R659 B.n302 B.n301 585
R660 B.n300 B.n201 585
R661 B.n299 B.n298 585
R662 B.n297 B.n202 585
R663 B.n296 B.n295 585
R664 B.n294 B.n203 585
R665 B.n293 B.n292 585
R666 B.n291 B.n204 585
R667 B.n290 B.n289 585
R668 B.n288 B.n205 585
R669 B.n287 B.n286 585
R670 B.n285 B.n206 585
R671 B.n284 B.n283 585
R672 B.n282 B.n207 585
R673 B.n281 B.n280 585
R674 B.n279 B.n208 585
R675 B.n278 B.n277 585
R676 B.n276 B.n209 585
R677 B.n275 B.n274 585
R678 B.n273 B.n210 585
R679 B.n272 B.n271 585
R680 B.n270 B.n211 585
R681 B.n269 B.n268 585
R682 B.n267 B.n212 585
R683 B.n266 B.n265 585
R684 B.n264 B.n213 585
R685 B.n263 B.n262 585
R686 B.n261 B.n214 585
R687 B.n260 B.n259 585
R688 B.n258 B.n215 585
R689 B.n257 B.n256 585
R690 B.n255 B.n216 585
R691 B.n254 B.n253 585
R692 B.n252 B.n217 585
R693 B.n251 B.n250 585
R694 B.n249 B.n218 585
R695 B.n248 B.n247 585
R696 B.n246 B.n219 585
R697 B.n245 B.n244 585
R698 B.n243 B.n220 585
R699 B.n242 B.n241 585
R700 B.n240 B.n221 585
R701 B.n239 B.n238 585
R702 B.n237 B.n222 585
R703 B.n236 B.n235 585
R704 B.n234 B.n223 585
R705 B.n233 B.n232 585
R706 B.n231 B.n224 585
R707 B.n230 B.n229 585
R708 B.n228 B.n225 585
R709 B.n227 B.n226 585
R710 B.n2 B.n0 585
R711 B.n873 B.n1 585
R712 B.n872 B.n871 585
R713 B.n870 B.n3 585
R714 B.n869 B.n868 585
R715 B.n867 B.n4 585
R716 B.n866 B.n865 585
R717 B.n864 B.n5 585
R718 B.n863 B.n862 585
R719 B.n861 B.n6 585
R720 B.n860 B.n859 585
R721 B.n858 B.n7 585
R722 B.n857 B.n856 585
R723 B.n855 B.n8 585
R724 B.n854 B.n853 585
R725 B.n852 B.n9 585
R726 B.n851 B.n850 585
R727 B.n849 B.n10 585
R728 B.n848 B.n847 585
R729 B.n846 B.n11 585
R730 B.n845 B.n844 585
R731 B.n843 B.n12 585
R732 B.n842 B.n841 585
R733 B.n840 B.n13 585
R734 B.n839 B.n838 585
R735 B.n837 B.n14 585
R736 B.n836 B.n835 585
R737 B.n834 B.n15 585
R738 B.n833 B.n832 585
R739 B.n831 B.n16 585
R740 B.n830 B.n829 585
R741 B.n828 B.n17 585
R742 B.n827 B.n826 585
R743 B.n825 B.n18 585
R744 B.n824 B.n823 585
R745 B.n822 B.n19 585
R746 B.n821 B.n820 585
R747 B.n819 B.n20 585
R748 B.n818 B.n817 585
R749 B.n816 B.n21 585
R750 B.n815 B.n814 585
R751 B.n813 B.n22 585
R752 B.n812 B.n811 585
R753 B.n810 B.n23 585
R754 B.n809 B.n808 585
R755 B.n807 B.n24 585
R756 B.n806 B.n805 585
R757 B.n804 B.n25 585
R758 B.n803 B.n802 585
R759 B.n801 B.n26 585
R760 B.n800 B.n799 585
R761 B.n798 B.n27 585
R762 B.n797 B.n796 585
R763 B.n795 B.n28 585
R764 B.n794 B.n793 585
R765 B.n792 B.n29 585
R766 B.n791 B.n790 585
R767 B.n875 B.n874 585
R768 B.n309 B.n308 545.355
R769 B.n790 B.n789 545.355
R770 B.n465 B.n464 545.355
R771 B.n634 B.n633 545.355
R772 B.n166 B.t6 346.76
R773 B.n174 B.t3 346.76
R774 B.n54 B.t9 346.76
R775 B.n60 B.t0 346.76
R776 B.n308 B.n199 163.367
R777 B.n304 B.n199 163.367
R778 B.n304 B.n303 163.367
R779 B.n303 B.n302 163.367
R780 B.n302 B.n201 163.367
R781 B.n298 B.n201 163.367
R782 B.n298 B.n297 163.367
R783 B.n297 B.n296 163.367
R784 B.n296 B.n203 163.367
R785 B.n292 B.n203 163.367
R786 B.n292 B.n291 163.367
R787 B.n291 B.n290 163.367
R788 B.n290 B.n205 163.367
R789 B.n286 B.n205 163.367
R790 B.n286 B.n285 163.367
R791 B.n285 B.n284 163.367
R792 B.n284 B.n207 163.367
R793 B.n280 B.n207 163.367
R794 B.n280 B.n279 163.367
R795 B.n279 B.n278 163.367
R796 B.n278 B.n209 163.367
R797 B.n274 B.n209 163.367
R798 B.n274 B.n273 163.367
R799 B.n273 B.n272 163.367
R800 B.n272 B.n211 163.367
R801 B.n268 B.n211 163.367
R802 B.n268 B.n267 163.367
R803 B.n267 B.n266 163.367
R804 B.n266 B.n213 163.367
R805 B.n262 B.n213 163.367
R806 B.n262 B.n261 163.367
R807 B.n261 B.n260 163.367
R808 B.n260 B.n215 163.367
R809 B.n256 B.n215 163.367
R810 B.n256 B.n255 163.367
R811 B.n255 B.n254 163.367
R812 B.n254 B.n217 163.367
R813 B.n250 B.n217 163.367
R814 B.n250 B.n249 163.367
R815 B.n249 B.n248 163.367
R816 B.n248 B.n219 163.367
R817 B.n244 B.n219 163.367
R818 B.n244 B.n243 163.367
R819 B.n243 B.n242 163.367
R820 B.n242 B.n221 163.367
R821 B.n238 B.n221 163.367
R822 B.n238 B.n237 163.367
R823 B.n237 B.n236 163.367
R824 B.n236 B.n223 163.367
R825 B.n232 B.n223 163.367
R826 B.n232 B.n231 163.367
R827 B.n231 B.n230 163.367
R828 B.n230 B.n225 163.367
R829 B.n226 B.n225 163.367
R830 B.n226 B.n2 163.367
R831 B.n874 B.n2 163.367
R832 B.n874 B.n873 163.367
R833 B.n873 B.n872 163.367
R834 B.n872 B.n3 163.367
R835 B.n868 B.n3 163.367
R836 B.n868 B.n867 163.367
R837 B.n867 B.n866 163.367
R838 B.n866 B.n5 163.367
R839 B.n862 B.n5 163.367
R840 B.n862 B.n861 163.367
R841 B.n861 B.n860 163.367
R842 B.n860 B.n7 163.367
R843 B.n856 B.n7 163.367
R844 B.n856 B.n855 163.367
R845 B.n855 B.n854 163.367
R846 B.n854 B.n9 163.367
R847 B.n850 B.n9 163.367
R848 B.n850 B.n849 163.367
R849 B.n849 B.n848 163.367
R850 B.n848 B.n11 163.367
R851 B.n844 B.n11 163.367
R852 B.n844 B.n843 163.367
R853 B.n843 B.n842 163.367
R854 B.n842 B.n13 163.367
R855 B.n838 B.n13 163.367
R856 B.n838 B.n837 163.367
R857 B.n837 B.n836 163.367
R858 B.n836 B.n15 163.367
R859 B.n832 B.n15 163.367
R860 B.n832 B.n831 163.367
R861 B.n831 B.n830 163.367
R862 B.n830 B.n17 163.367
R863 B.n826 B.n17 163.367
R864 B.n826 B.n825 163.367
R865 B.n825 B.n824 163.367
R866 B.n824 B.n19 163.367
R867 B.n820 B.n19 163.367
R868 B.n820 B.n819 163.367
R869 B.n819 B.n818 163.367
R870 B.n818 B.n21 163.367
R871 B.n814 B.n21 163.367
R872 B.n814 B.n813 163.367
R873 B.n813 B.n812 163.367
R874 B.n812 B.n23 163.367
R875 B.n808 B.n23 163.367
R876 B.n808 B.n807 163.367
R877 B.n807 B.n806 163.367
R878 B.n806 B.n25 163.367
R879 B.n802 B.n25 163.367
R880 B.n802 B.n801 163.367
R881 B.n801 B.n800 163.367
R882 B.n800 B.n27 163.367
R883 B.n796 B.n27 163.367
R884 B.n796 B.n795 163.367
R885 B.n795 B.n794 163.367
R886 B.n794 B.n29 163.367
R887 B.n790 B.n29 163.367
R888 B.n310 B.n309 163.367
R889 B.n310 B.n197 163.367
R890 B.n314 B.n197 163.367
R891 B.n315 B.n314 163.367
R892 B.n316 B.n315 163.367
R893 B.n316 B.n195 163.367
R894 B.n320 B.n195 163.367
R895 B.n321 B.n320 163.367
R896 B.n322 B.n321 163.367
R897 B.n322 B.n193 163.367
R898 B.n326 B.n193 163.367
R899 B.n327 B.n326 163.367
R900 B.n328 B.n327 163.367
R901 B.n328 B.n191 163.367
R902 B.n332 B.n191 163.367
R903 B.n333 B.n332 163.367
R904 B.n334 B.n333 163.367
R905 B.n334 B.n189 163.367
R906 B.n338 B.n189 163.367
R907 B.n339 B.n338 163.367
R908 B.n340 B.n339 163.367
R909 B.n340 B.n187 163.367
R910 B.n344 B.n187 163.367
R911 B.n345 B.n344 163.367
R912 B.n346 B.n345 163.367
R913 B.n346 B.n185 163.367
R914 B.n350 B.n185 163.367
R915 B.n351 B.n350 163.367
R916 B.n352 B.n351 163.367
R917 B.n352 B.n183 163.367
R918 B.n356 B.n183 163.367
R919 B.n357 B.n356 163.367
R920 B.n358 B.n357 163.367
R921 B.n358 B.n181 163.367
R922 B.n362 B.n181 163.367
R923 B.n363 B.n362 163.367
R924 B.n364 B.n363 163.367
R925 B.n364 B.n179 163.367
R926 B.n368 B.n179 163.367
R927 B.n369 B.n368 163.367
R928 B.n370 B.n369 163.367
R929 B.n370 B.n177 163.367
R930 B.n374 B.n177 163.367
R931 B.n375 B.n374 163.367
R932 B.n376 B.n375 163.367
R933 B.n376 B.n173 163.367
R934 B.n381 B.n173 163.367
R935 B.n382 B.n381 163.367
R936 B.n383 B.n382 163.367
R937 B.n383 B.n171 163.367
R938 B.n387 B.n171 163.367
R939 B.n388 B.n387 163.367
R940 B.n389 B.n388 163.367
R941 B.n389 B.n169 163.367
R942 B.n393 B.n169 163.367
R943 B.n394 B.n393 163.367
R944 B.n394 B.n165 163.367
R945 B.n398 B.n165 163.367
R946 B.n399 B.n398 163.367
R947 B.n400 B.n399 163.367
R948 B.n400 B.n163 163.367
R949 B.n404 B.n163 163.367
R950 B.n405 B.n404 163.367
R951 B.n406 B.n405 163.367
R952 B.n406 B.n161 163.367
R953 B.n410 B.n161 163.367
R954 B.n411 B.n410 163.367
R955 B.n412 B.n411 163.367
R956 B.n412 B.n159 163.367
R957 B.n416 B.n159 163.367
R958 B.n417 B.n416 163.367
R959 B.n418 B.n417 163.367
R960 B.n418 B.n157 163.367
R961 B.n422 B.n157 163.367
R962 B.n423 B.n422 163.367
R963 B.n424 B.n423 163.367
R964 B.n424 B.n155 163.367
R965 B.n428 B.n155 163.367
R966 B.n429 B.n428 163.367
R967 B.n430 B.n429 163.367
R968 B.n430 B.n153 163.367
R969 B.n434 B.n153 163.367
R970 B.n435 B.n434 163.367
R971 B.n436 B.n435 163.367
R972 B.n436 B.n151 163.367
R973 B.n440 B.n151 163.367
R974 B.n441 B.n440 163.367
R975 B.n442 B.n441 163.367
R976 B.n442 B.n149 163.367
R977 B.n446 B.n149 163.367
R978 B.n447 B.n446 163.367
R979 B.n448 B.n447 163.367
R980 B.n448 B.n147 163.367
R981 B.n452 B.n147 163.367
R982 B.n453 B.n452 163.367
R983 B.n454 B.n453 163.367
R984 B.n454 B.n145 163.367
R985 B.n458 B.n145 163.367
R986 B.n459 B.n458 163.367
R987 B.n460 B.n459 163.367
R988 B.n460 B.n143 163.367
R989 B.n464 B.n143 163.367
R990 B.n466 B.n465 163.367
R991 B.n466 B.n141 163.367
R992 B.n470 B.n141 163.367
R993 B.n471 B.n470 163.367
R994 B.n472 B.n471 163.367
R995 B.n472 B.n139 163.367
R996 B.n476 B.n139 163.367
R997 B.n477 B.n476 163.367
R998 B.n478 B.n477 163.367
R999 B.n478 B.n137 163.367
R1000 B.n482 B.n137 163.367
R1001 B.n483 B.n482 163.367
R1002 B.n484 B.n483 163.367
R1003 B.n484 B.n135 163.367
R1004 B.n488 B.n135 163.367
R1005 B.n489 B.n488 163.367
R1006 B.n490 B.n489 163.367
R1007 B.n490 B.n133 163.367
R1008 B.n494 B.n133 163.367
R1009 B.n495 B.n494 163.367
R1010 B.n496 B.n495 163.367
R1011 B.n496 B.n131 163.367
R1012 B.n500 B.n131 163.367
R1013 B.n501 B.n500 163.367
R1014 B.n502 B.n501 163.367
R1015 B.n502 B.n129 163.367
R1016 B.n506 B.n129 163.367
R1017 B.n507 B.n506 163.367
R1018 B.n508 B.n507 163.367
R1019 B.n508 B.n127 163.367
R1020 B.n512 B.n127 163.367
R1021 B.n513 B.n512 163.367
R1022 B.n514 B.n513 163.367
R1023 B.n514 B.n125 163.367
R1024 B.n518 B.n125 163.367
R1025 B.n519 B.n518 163.367
R1026 B.n520 B.n519 163.367
R1027 B.n520 B.n123 163.367
R1028 B.n524 B.n123 163.367
R1029 B.n525 B.n524 163.367
R1030 B.n526 B.n525 163.367
R1031 B.n526 B.n121 163.367
R1032 B.n530 B.n121 163.367
R1033 B.n531 B.n530 163.367
R1034 B.n532 B.n531 163.367
R1035 B.n532 B.n119 163.367
R1036 B.n536 B.n119 163.367
R1037 B.n537 B.n536 163.367
R1038 B.n538 B.n537 163.367
R1039 B.n538 B.n117 163.367
R1040 B.n542 B.n117 163.367
R1041 B.n543 B.n542 163.367
R1042 B.n544 B.n543 163.367
R1043 B.n544 B.n115 163.367
R1044 B.n548 B.n115 163.367
R1045 B.n549 B.n548 163.367
R1046 B.n550 B.n549 163.367
R1047 B.n550 B.n113 163.367
R1048 B.n554 B.n113 163.367
R1049 B.n555 B.n554 163.367
R1050 B.n556 B.n555 163.367
R1051 B.n556 B.n111 163.367
R1052 B.n560 B.n111 163.367
R1053 B.n561 B.n560 163.367
R1054 B.n562 B.n561 163.367
R1055 B.n562 B.n109 163.367
R1056 B.n566 B.n109 163.367
R1057 B.n567 B.n566 163.367
R1058 B.n568 B.n567 163.367
R1059 B.n568 B.n107 163.367
R1060 B.n572 B.n107 163.367
R1061 B.n573 B.n572 163.367
R1062 B.n574 B.n573 163.367
R1063 B.n574 B.n105 163.367
R1064 B.n578 B.n105 163.367
R1065 B.n579 B.n578 163.367
R1066 B.n580 B.n579 163.367
R1067 B.n580 B.n103 163.367
R1068 B.n584 B.n103 163.367
R1069 B.n585 B.n584 163.367
R1070 B.n586 B.n585 163.367
R1071 B.n586 B.n101 163.367
R1072 B.n590 B.n101 163.367
R1073 B.n591 B.n590 163.367
R1074 B.n592 B.n591 163.367
R1075 B.n592 B.n99 163.367
R1076 B.n596 B.n99 163.367
R1077 B.n597 B.n596 163.367
R1078 B.n598 B.n597 163.367
R1079 B.n598 B.n97 163.367
R1080 B.n602 B.n97 163.367
R1081 B.n603 B.n602 163.367
R1082 B.n604 B.n603 163.367
R1083 B.n604 B.n95 163.367
R1084 B.n608 B.n95 163.367
R1085 B.n609 B.n608 163.367
R1086 B.n610 B.n609 163.367
R1087 B.n610 B.n93 163.367
R1088 B.n614 B.n93 163.367
R1089 B.n615 B.n614 163.367
R1090 B.n616 B.n615 163.367
R1091 B.n616 B.n91 163.367
R1092 B.n620 B.n91 163.367
R1093 B.n621 B.n620 163.367
R1094 B.n622 B.n621 163.367
R1095 B.n622 B.n89 163.367
R1096 B.n626 B.n89 163.367
R1097 B.n627 B.n626 163.367
R1098 B.n628 B.n627 163.367
R1099 B.n628 B.n87 163.367
R1100 B.n632 B.n87 163.367
R1101 B.n633 B.n632 163.367
R1102 B.n789 B.n788 163.367
R1103 B.n788 B.n31 163.367
R1104 B.n784 B.n31 163.367
R1105 B.n784 B.n783 163.367
R1106 B.n783 B.n782 163.367
R1107 B.n782 B.n33 163.367
R1108 B.n778 B.n33 163.367
R1109 B.n778 B.n777 163.367
R1110 B.n777 B.n776 163.367
R1111 B.n776 B.n35 163.367
R1112 B.n772 B.n35 163.367
R1113 B.n772 B.n771 163.367
R1114 B.n771 B.n770 163.367
R1115 B.n770 B.n37 163.367
R1116 B.n766 B.n37 163.367
R1117 B.n766 B.n765 163.367
R1118 B.n765 B.n764 163.367
R1119 B.n764 B.n39 163.367
R1120 B.n760 B.n39 163.367
R1121 B.n760 B.n759 163.367
R1122 B.n759 B.n758 163.367
R1123 B.n758 B.n41 163.367
R1124 B.n754 B.n41 163.367
R1125 B.n754 B.n753 163.367
R1126 B.n753 B.n752 163.367
R1127 B.n752 B.n43 163.367
R1128 B.n748 B.n43 163.367
R1129 B.n748 B.n747 163.367
R1130 B.n747 B.n746 163.367
R1131 B.n746 B.n45 163.367
R1132 B.n742 B.n45 163.367
R1133 B.n742 B.n741 163.367
R1134 B.n741 B.n740 163.367
R1135 B.n740 B.n47 163.367
R1136 B.n736 B.n47 163.367
R1137 B.n736 B.n735 163.367
R1138 B.n735 B.n734 163.367
R1139 B.n734 B.n49 163.367
R1140 B.n730 B.n49 163.367
R1141 B.n730 B.n729 163.367
R1142 B.n729 B.n728 163.367
R1143 B.n728 B.n51 163.367
R1144 B.n724 B.n51 163.367
R1145 B.n724 B.n723 163.367
R1146 B.n723 B.n722 163.367
R1147 B.n722 B.n53 163.367
R1148 B.n717 B.n53 163.367
R1149 B.n717 B.n716 163.367
R1150 B.n716 B.n715 163.367
R1151 B.n715 B.n57 163.367
R1152 B.n711 B.n57 163.367
R1153 B.n711 B.n710 163.367
R1154 B.n710 B.n709 163.367
R1155 B.n709 B.n59 163.367
R1156 B.n705 B.n59 163.367
R1157 B.n705 B.n704 163.367
R1158 B.n704 B.n63 163.367
R1159 B.n700 B.n63 163.367
R1160 B.n700 B.n699 163.367
R1161 B.n699 B.n698 163.367
R1162 B.n698 B.n65 163.367
R1163 B.n694 B.n65 163.367
R1164 B.n694 B.n693 163.367
R1165 B.n693 B.n692 163.367
R1166 B.n692 B.n67 163.367
R1167 B.n688 B.n67 163.367
R1168 B.n688 B.n687 163.367
R1169 B.n687 B.n686 163.367
R1170 B.n686 B.n69 163.367
R1171 B.n682 B.n69 163.367
R1172 B.n682 B.n681 163.367
R1173 B.n681 B.n680 163.367
R1174 B.n680 B.n71 163.367
R1175 B.n676 B.n71 163.367
R1176 B.n676 B.n675 163.367
R1177 B.n675 B.n674 163.367
R1178 B.n674 B.n73 163.367
R1179 B.n670 B.n73 163.367
R1180 B.n670 B.n669 163.367
R1181 B.n669 B.n668 163.367
R1182 B.n668 B.n75 163.367
R1183 B.n664 B.n75 163.367
R1184 B.n664 B.n663 163.367
R1185 B.n663 B.n662 163.367
R1186 B.n662 B.n77 163.367
R1187 B.n658 B.n77 163.367
R1188 B.n658 B.n657 163.367
R1189 B.n657 B.n656 163.367
R1190 B.n656 B.n79 163.367
R1191 B.n652 B.n79 163.367
R1192 B.n652 B.n651 163.367
R1193 B.n651 B.n650 163.367
R1194 B.n650 B.n81 163.367
R1195 B.n646 B.n81 163.367
R1196 B.n646 B.n645 163.367
R1197 B.n645 B.n644 163.367
R1198 B.n644 B.n83 163.367
R1199 B.n640 B.n83 163.367
R1200 B.n640 B.n639 163.367
R1201 B.n639 B.n638 163.367
R1202 B.n638 B.n85 163.367
R1203 B.n634 B.n85 163.367
R1204 B.n166 B.t8 163.186
R1205 B.n60 B.t1 163.186
R1206 B.n174 B.t5 163.169
R1207 B.n54 B.t10 163.169
R1208 B.n167 B.t7 110.436
R1209 B.n61 B.t2 110.436
R1210 B.n175 B.t4 110.418
R1211 B.n55 B.t11 110.418
R1212 B.n168 B.n167 59.5399
R1213 B.n379 B.n175 59.5399
R1214 B.n719 B.n55 59.5399
R1215 B.n62 B.n61 59.5399
R1216 B.n167 B.n166 52.752
R1217 B.n175 B.n174 52.752
R1218 B.n55 B.n54 52.752
R1219 B.n61 B.n60 52.752
R1220 B.n791 B.n30 35.4346
R1221 B.n463 B.n142 35.4346
R1222 B.n307 B.n198 35.4346
R1223 B.n635 B.n86 35.4346
R1224 B B.n875 18.0485
R1225 B.n787 B.n30 10.6151
R1226 B.n787 B.n786 10.6151
R1227 B.n786 B.n785 10.6151
R1228 B.n785 B.n32 10.6151
R1229 B.n781 B.n32 10.6151
R1230 B.n781 B.n780 10.6151
R1231 B.n780 B.n779 10.6151
R1232 B.n779 B.n34 10.6151
R1233 B.n775 B.n34 10.6151
R1234 B.n775 B.n774 10.6151
R1235 B.n774 B.n773 10.6151
R1236 B.n773 B.n36 10.6151
R1237 B.n769 B.n36 10.6151
R1238 B.n769 B.n768 10.6151
R1239 B.n768 B.n767 10.6151
R1240 B.n767 B.n38 10.6151
R1241 B.n763 B.n38 10.6151
R1242 B.n763 B.n762 10.6151
R1243 B.n762 B.n761 10.6151
R1244 B.n761 B.n40 10.6151
R1245 B.n757 B.n40 10.6151
R1246 B.n757 B.n756 10.6151
R1247 B.n756 B.n755 10.6151
R1248 B.n755 B.n42 10.6151
R1249 B.n751 B.n42 10.6151
R1250 B.n751 B.n750 10.6151
R1251 B.n750 B.n749 10.6151
R1252 B.n749 B.n44 10.6151
R1253 B.n745 B.n44 10.6151
R1254 B.n745 B.n744 10.6151
R1255 B.n744 B.n743 10.6151
R1256 B.n743 B.n46 10.6151
R1257 B.n739 B.n46 10.6151
R1258 B.n739 B.n738 10.6151
R1259 B.n738 B.n737 10.6151
R1260 B.n737 B.n48 10.6151
R1261 B.n733 B.n48 10.6151
R1262 B.n733 B.n732 10.6151
R1263 B.n732 B.n731 10.6151
R1264 B.n731 B.n50 10.6151
R1265 B.n727 B.n50 10.6151
R1266 B.n727 B.n726 10.6151
R1267 B.n726 B.n725 10.6151
R1268 B.n725 B.n52 10.6151
R1269 B.n721 B.n52 10.6151
R1270 B.n721 B.n720 10.6151
R1271 B.n718 B.n56 10.6151
R1272 B.n714 B.n56 10.6151
R1273 B.n714 B.n713 10.6151
R1274 B.n713 B.n712 10.6151
R1275 B.n712 B.n58 10.6151
R1276 B.n708 B.n58 10.6151
R1277 B.n708 B.n707 10.6151
R1278 B.n707 B.n706 10.6151
R1279 B.n703 B.n702 10.6151
R1280 B.n702 B.n701 10.6151
R1281 B.n701 B.n64 10.6151
R1282 B.n697 B.n64 10.6151
R1283 B.n697 B.n696 10.6151
R1284 B.n696 B.n695 10.6151
R1285 B.n695 B.n66 10.6151
R1286 B.n691 B.n66 10.6151
R1287 B.n691 B.n690 10.6151
R1288 B.n690 B.n689 10.6151
R1289 B.n689 B.n68 10.6151
R1290 B.n685 B.n68 10.6151
R1291 B.n685 B.n684 10.6151
R1292 B.n684 B.n683 10.6151
R1293 B.n683 B.n70 10.6151
R1294 B.n679 B.n70 10.6151
R1295 B.n679 B.n678 10.6151
R1296 B.n678 B.n677 10.6151
R1297 B.n677 B.n72 10.6151
R1298 B.n673 B.n72 10.6151
R1299 B.n673 B.n672 10.6151
R1300 B.n672 B.n671 10.6151
R1301 B.n671 B.n74 10.6151
R1302 B.n667 B.n74 10.6151
R1303 B.n667 B.n666 10.6151
R1304 B.n666 B.n665 10.6151
R1305 B.n665 B.n76 10.6151
R1306 B.n661 B.n76 10.6151
R1307 B.n661 B.n660 10.6151
R1308 B.n660 B.n659 10.6151
R1309 B.n659 B.n78 10.6151
R1310 B.n655 B.n78 10.6151
R1311 B.n655 B.n654 10.6151
R1312 B.n654 B.n653 10.6151
R1313 B.n653 B.n80 10.6151
R1314 B.n649 B.n80 10.6151
R1315 B.n649 B.n648 10.6151
R1316 B.n648 B.n647 10.6151
R1317 B.n647 B.n82 10.6151
R1318 B.n643 B.n82 10.6151
R1319 B.n643 B.n642 10.6151
R1320 B.n642 B.n641 10.6151
R1321 B.n641 B.n84 10.6151
R1322 B.n637 B.n84 10.6151
R1323 B.n637 B.n636 10.6151
R1324 B.n636 B.n635 10.6151
R1325 B.n467 B.n142 10.6151
R1326 B.n468 B.n467 10.6151
R1327 B.n469 B.n468 10.6151
R1328 B.n469 B.n140 10.6151
R1329 B.n473 B.n140 10.6151
R1330 B.n474 B.n473 10.6151
R1331 B.n475 B.n474 10.6151
R1332 B.n475 B.n138 10.6151
R1333 B.n479 B.n138 10.6151
R1334 B.n480 B.n479 10.6151
R1335 B.n481 B.n480 10.6151
R1336 B.n481 B.n136 10.6151
R1337 B.n485 B.n136 10.6151
R1338 B.n486 B.n485 10.6151
R1339 B.n487 B.n486 10.6151
R1340 B.n487 B.n134 10.6151
R1341 B.n491 B.n134 10.6151
R1342 B.n492 B.n491 10.6151
R1343 B.n493 B.n492 10.6151
R1344 B.n493 B.n132 10.6151
R1345 B.n497 B.n132 10.6151
R1346 B.n498 B.n497 10.6151
R1347 B.n499 B.n498 10.6151
R1348 B.n499 B.n130 10.6151
R1349 B.n503 B.n130 10.6151
R1350 B.n504 B.n503 10.6151
R1351 B.n505 B.n504 10.6151
R1352 B.n505 B.n128 10.6151
R1353 B.n509 B.n128 10.6151
R1354 B.n510 B.n509 10.6151
R1355 B.n511 B.n510 10.6151
R1356 B.n511 B.n126 10.6151
R1357 B.n515 B.n126 10.6151
R1358 B.n516 B.n515 10.6151
R1359 B.n517 B.n516 10.6151
R1360 B.n517 B.n124 10.6151
R1361 B.n521 B.n124 10.6151
R1362 B.n522 B.n521 10.6151
R1363 B.n523 B.n522 10.6151
R1364 B.n523 B.n122 10.6151
R1365 B.n527 B.n122 10.6151
R1366 B.n528 B.n527 10.6151
R1367 B.n529 B.n528 10.6151
R1368 B.n529 B.n120 10.6151
R1369 B.n533 B.n120 10.6151
R1370 B.n534 B.n533 10.6151
R1371 B.n535 B.n534 10.6151
R1372 B.n535 B.n118 10.6151
R1373 B.n539 B.n118 10.6151
R1374 B.n540 B.n539 10.6151
R1375 B.n541 B.n540 10.6151
R1376 B.n541 B.n116 10.6151
R1377 B.n545 B.n116 10.6151
R1378 B.n546 B.n545 10.6151
R1379 B.n547 B.n546 10.6151
R1380 B.n547 B.n114 10.6151
R1381 B.n551 B.n114 10.6151
R1382 B.n552 B.n551 10.6151
R1383 B.n553 B.n552 10.6151
R1384 B.n553 B.n112 10.6151
R1385 B.n557 B.n112 10.6151
R1386 B.n558 B.n557 10.6151
R1387 B.n559 B.n558 10.6151
R1388 B.n559 B.n110 10.6151
R1389 B.n563 B.n110 10.6151
R1390 B.n564 B.n563 10.6151
R1391 B.n565 B.n564 10.6151
R1392 B.n565 B.n108 10.6151
R1393 B.n569 B.n108 10.6151
R1394 B.n570 B.n569 10.6151
R1395 B.n571 B.n570 10.6151
R1396 B.n571 B.n106 10.6151
R1397 B.n575 B.n106 10.6151
R1398 B.n576 B.n575 10.6151
R1399 B.n577 B.n576 10.6151
R1400 B.n577 B.n104 10.6151
R1401 B.n581 B.n104 10.6151
R1402 B.n582 B.n581 10.6151
R1403 B.n583 B.n582 10.6151
R1404 B.n583 B.n102 10.6151
R1405 B.n587 B.n102 10.6151
R1406 B.n588 B.n587 10.6151
R1407 B.n589 B.n588 10.6151
R1408 B.n589 B.n100 10.6151
R1409 B.n593 B.n100 10.6151
R1410 B.n594 B.n593 10.6151
R1411 B.n595 B.n594 10.6151
R1412 B.n595 B.n98 10.6151
R1413 B.n599 B.n98 10.6151
R1414 B.n600 B.n599 10.6151
R1415 B.n601 B.n600 10.6151
R1416 B.n601 B.n96 10.6151
R1417 B.n605 B.n96 10.6151
R1418 B.n606 B.n605 10.6151
R1419 B.n607 B.n606 10.6151
R1420 B.n607 B.n94 10.6151
R1421 B.n611 B.n94 10.6151
R1422 B.n612 B.n611 10.6151
R1423 B.n613 B.n612 10.6151
R1424 B.n613 B.n92 10.6151
R1425 B.n617 B.n92 10.6151
R1426 B.n618 B.n617 10.6151
R1427 B.n619 B.n618 10.6151
R1428 B.n619 B.n90 10.6151
R1429 B.n623 B.n90 10.6151
R1430 B.n624 B.n623 10.6151
R1431 B.n625 B.n624 10.6151
R1432 B.n625 B.n88 10.6151
R1433 B.n629 B.n88 10.6151
R1434 B.n630 B.n629 10.6151
R1435 B.n631 B.n630 10.6151
R1436 B.n631 B.n86 10.6151
R1437 B.n311 B.n198 10.6151
R1438 B.n312 B.n311 10.6151
R1439 B.n313 B.n312 10.6151
R1440 B.n313 B.n196 10.6151
R1441 B.n317 B.n196 10.6151
R1442 B.n318 B.n317 10.6151
R1443 B.n319 B.n318 10.6151
R1444 B.n319 B.n194 10.6151
R1445 B.n323 B.n194 10.6151
R1446 B.n324 B.n323 10.6151
R1447 B.n325 B.n324 10.6151
R1448 B.n325 B.n192 10.6151
R1449 B.n329 B.n192 10.6151
R1450 B.n330 B.n329 10.6151
R1451 B.n331 B.n330 10.6151
R1452 B.n331 B.n190 10.6151
R1453 B.n335 B.n190 10.6151
R1454 B.n336 B.n335 10.6151
R1455 B.n337 B.n336 10.6151
R1456 B.n337 B.n188 10.6151
R1457 B.n341 B.n188 10.6151
R1458 B.n342 B.n341 10.6151
R1459 B.n343 B.n342 10.6151
R1460 B.n343 B.n186 10.6151
R1461 B.n347 B.n186 10.6151
R1462 B.n348 B.n347 10.6151
R1463 B.n349 B.n348 10.6151
R1464 B.n349 B.n184 10.6151
R1465 B.n353 B.n184 10.6151
R1466 B.n354 B.n353 10.6151
R1467 B.n355 B.n354 10.6151
R1468 B.n355 B.n182 10.6151
R1469 B.n359 B.n182 10.6151
R1470 B.n360 B.n359 10.6151
R1471 B.n361 B.n360 10.6151
R1472 B.n361 B.n180 10.6151
R1473 B.n365 B.n180 10.6151
R1474 B.n366 B.n365 10.6151
R1475 B.n367 B.n366 10.6151
R1476 B.n367 B.n178 10.6151
R1477 B.n371 B.n178 10.6151
R1478 B.n372 B.n371 10.6151
R1479 B.n373 B.n372 10.6151
R1480 B.n373 B.n176 10.6151
R1481 B.n377 B.n176 10.6151
R1482 B.n378 B.n377 10.6151
R1483 B.n380 B.n172 10.6151
R1484 B.n384 B.n172 10.6151
R1485 B.n385 B.n384 10.6151
R1486 B.n386 B.n385 10.6151
R1487 B.n386 B.n170 10.6151
R1488 B.n390 B.n170 10.6151
R1489 B.n391 B.n390 10.6151
R1490 B.n392 B.n391 10.6151
R1491 B.n396 B.n395 10.6151
R1492 B.n397 B.n396 10.6151
R1493 B.n397 B.n164 10.6151
R1494 B.n401 B.n164 10.6151
R1495 B.n402 B.n401 10.6151
R1496 B.n403 B.n402 10.6151
R1497 B.n403 B.n162 10.6151
R1498 B.n407 B.n162 10.6151
R1499 B.n408 B.n407 10.6151
R1500 B.n409 B.n408 10.6151
R1501 B.n409 B.n160 10.6151
R1502 B.n413 B.n160 10.6151
R1503 B.n414 B.n413 10.6151
R1504 B.n415 B.n414 10.6151
R1505 B.n415 B.n158 10.6151
R1506 B.n419 B.n158 10.6151
R1507 B.n420 B.n419 10.6151
R1508 B.n421 B.n420 10.6151
R1509 B.n421 B.n156 10.6151
R1510 B.n425 B.n156 10.6151
R1511 B.n426 B.n425 10.6151
R1512 B.n427 B.n426 10.6151
R1513 B.n427 B.n154 10.6151
R1514 B.n431 B.n154 10.6151
R1515 B.n432 B.n431 10.6151
R1516 B.n433 B.n432 10.6151
R1517 B.n433 B.n152 10.6151
R1518 B.n437 B.n152 10.6151
R1519 B.n438 B.n437 10.6151
R1520 B.n439 B.n438 10.6151
R1521 B.n439 B.n150 10.6151
R1522 B.n443 B.n150 10.6151
R1523 B.n444 B.n443 10.6151
R1524 B.n445 B.n444 10.6151
R1525 B.n445 B.n148 10.6151
R1526 B.n449 B.n148 10.6151
R1527 B.n450 B.n449 10.6151
R1528 B.n451 B.n450 10.6151
R1529 B.n451 B.n146 10.6151
R1530 B.n455 B.n146 10.6151
R1531 B.n456 B.n455 10.6151
R1532 B.n457 B.n456 10.6151
R1533 B.n457 B.n144 10.6151
R1534 B.n461 B.n144 10.6151
R1535 B.n462 B.n461 10.6151
R1536 B.n463 B.n462 10.6151
R1537 B.n307 B.n306 10.6151
R1538 B.n306 B.n305 10.6151
R1539 B.n305 B.n200 10.6151
R1540 B.n301 B.n200 10.6151
R1541 B.n301 B.n300 10.6151
R1542 B.n300 B.n299 10.6151
R1543 B.n299 B.n202 10.6151
R1544 B.n295 B.n202 10.6151
R1545 B.n295 B.n294 10.6151
R1546 B.n294 B.n293 10.6151
R1547 B.n293 B.n204 10.6151
R1548 B.n289 B.n204 10.6151
R1549 B.n289 B.n288 10.6151
R1550 B.n288 B.n287 10.6151
R1551 B.n287 B.n206 10.6151
R1552 B.n283 B.n206 10.6151
R1553 B.n283 B.n282 10.6151
R1554 B.n282 B.n281 10.6151
R1555 B.n281 B.n208 10.6151
R1556 B.n277 B.n208 10.6151
R1557 B.n277 B.n276 10.6151
R1558 B.n276 B.n275 10.6151
R1559 B.n275 B.n210 10.6151
R1560 B.n271 B.n210 10.6151
R1561 B.n271 B.n270 10.6151
R1562 B.n270 B.n269 10.6151
R1563 B.n269 B.n212 10.6151
R1564 B.n265 B.n212 10.6151
R1565 B.n265 B.n264 10.6151
R1566 B.n264 B.n263 10.6151
R1567 B.n263 B.n214 10.6151
R1568 B.n259 B.n214 10.6151
R1569 B.n259 B.n258 10.6151
R1570 B.n258 B.n257 10.6151
R1571 B.n257 B.n216 10.6151
R1572 B.n253 B.n216 10.6151
R1573 B.n253 B.n252 10.6151
R1574 B.n252 B.n251 10.6151
R1575 B.n251 B.n218 10.6151
R1576 B.n247 B.n218 10.6151
R1577 B.n247 B.n246 10.6151
R1578 B.n246 B.n245 10.6151
R1579 B.n245 B.n220 10.6151
R1580 B.n241 B.n220 10.6151
R1581 B.n241 B.n240 10.6151
R1582 B.n240 B.n239 10.6151
R1583 B.n239 B.n222 10.6151
R1584 B.n235 B.n222 10.6151
R1585 B.n235 B.n234 10.6151
R1586 B.n234 B.n233 10.6151
R1587 B.n233 B.n224 10.6151
R1588 B.n229 B.n224 10.6151
R1589 B.n229 B.n228 10.6151
R1590 B.n228 B.n227 10.6151
R1591 B.n227 B.n0 10.6151
R1592 B.n871 B.n1 10.6151
R1593 B.n871 B.n870 10.6151
R1594 B.n870 B.n869 10.6151
R1595 B.n869 B.n4 10.6151
R1596 B.n865 B.n4 10.6151
R1597 B.n865 B.n864 10.6151
R1598 B.n864 B.n863 10.6151
R1599 B.n863 B.n6 10.6151
R1600 B.n859 B.n6 10.6151
R1601 B.n859 B.n858 10.6151
R1602 B.n858 B.n857 10.6151
R1603 B.n857 B.n8 10.6151
R1604 B.n853 B.n8 10.6151
R1605 B.n853 B.n852 10.6151
R1606 B.n852 B.n851 10.6151
R1607 B.n851 B.n10 10.6151
R1608 B.n847 B.n10 10.6151
R1609 B.n847 B.n846 10.6151
R1610 B.n846 B.n845 10.6151
R1611 B.n845 B.n12 10.6151
R1612 B.n841 B.n12 10.6151
R1613 B.n841 B.n840 10.6151
R1614 B.n840 B.n839 10.6151
R1615 B.n839 B.n14 10.6151
R1616 B.n835 B.n14 10.6151
R1617 B.n835 B.n834 10.6151
R1618 B.n834 B.n833 10.6151
R1619 B.n833 B.n16 10.6151
R1620 B.n829 B.n16 10.6151
R1621 B.n829 B.n828 10.6151
R1622 B.n828 B.n827 10.6151
R1623 B.n827 B.n18 10.6151
R1624 B.n823 B.n18 10.6151
R1625 B.n823 B.n822 10.6151
R1626 B.n822 B.n821 10.6151
R1627 B.n821 B.n20 10.6151
R1628 B.n817 B.n20 10.6151
R1629 B.n817 B.n816 10.6151
R1630 B.n816 B.n815 10.6151
R1631 B.n815 B.n22 10.6151
R1632 B.n811 B.n22 10.6151
R1633 B.n811 B.n810 10.6151
R1634 B.n810 B.n809 10.6151
R1635 B.n809 B.n24 10.6151
R1636 B.n805 B.n24 10.6151
R1637 B.n805 B.n804 10.6151
R1638 B.n804 B.n803 10.6151
R1639 B.n803 B.n26 10.6151
R1640 B.n799 B.n26 10.6151
R1641 B.n799 B.n798 10.6151
R1642 B.n798 B.n797 10.6151
R1643 B.n797 B.n28 10.6151
R1644 B.n793 B.n28 10.6151
R1645 B.n793 B.n792 10.6151
R1646 B.n792 B.n791 10.6151
R1647 B.n719 B.n718 6.5566
R1648 B.n706 B.n62 6.5566
R1649 B.n380 B.n379 6.5566
R1650 B.n392 B.n168 6.5566
R1651 B.n720 B.n719 4.05904
R1652 B.n703 B.n62 4.05904
R1653 B.n379 B.n378 4.05904
R1654 B.n395 B.n168 4.05904
R1655 B.n875 B.n0 2.81026
R1656 B.n875 B.n1 2.81026
C0 VP VDD1 12.3685f
C1 VP w_n4234_n3726# 9.58005f
C2 VN VDD1 0.152929f
C3 VP VTAIL 12.4578f
C4 VN w_n4234_n3726# 9.02945f
C5 VN VTAIL 12.443501f
C6 B VDD2 2.64926f
C7 VN VP 8.42298f
C8 VDD1 VDD2 2.03833f
C9 VDD2 w_n4234_n3726# 2.96777f
C10 VTAIL VDD2 11.279099f
C11 B VDD1 2.53952f
C12 B w_n4234_n3726# 10.6958f
C13 VP VDD2 0.556998f
C14 VTAIL B 4.03703f
C15 VN VDD2 11.968599f
C16 VDD1 w_n4234_n3726# 2.83505f
C17 VTAIL VDD1 11.2303f
C18 VP B 2.17566f
C19 VTAIL w_n4234_n3726# 3.43671f
C20 VN B 1.25096f
C21 VDD2 VSUBS 2.11761f
C22 VDD1 VSUBS 1.91966f
C23 VTAIL VSUBS 1.308823f
C24 VN VSUBS 7.3913f
C25 VP VSUBS 4.033945f
C26 B VSUBS 5.255862f
C27 w_n4234_n3726# VSUBS 0.193731p
C28 B.n0 VSUBS 0.005668f
C29 B.n1 VSUBS 0.005668f
C30 B.n2 VSUBS 0.008963f
C31 B.n3 VSUBS 0.008963f
C32 B.n4 VSUBS 0.008963f
C33 B.n5 VSUBS 0.008963f
C34 B.n6 VSUBS 0.008963f
C35 B.n7 VSUBS 0.008963f
C36 B.n8 VSUBS 0.008963f
C37 B.n9 VSUBS 0.008963f
C38 B.n10 VSUBS 0.008963f
C39 B.n11 VSUBS 0.008963f
C40 B.n12 VSUBS 0.008963f
C41 B.n13 VSUBS 0.008963f
C42 B.n14 VSUBS 0.008963f
C43 B.n15 VSUBS 0.008963f
C44 B.n16 VSUBS 0.008963f
C45 B.n17 VSUBS 0.008963f
C46 B.n18 VSUBS 0.008963f
C47 B.n19 VSUBS 0.008963f
C48 B.n20 VSUBS 0.008963f
C49 B.n21 VSUBS 0.008963f
C50 B.n22 VSUBS 0.008963f
C51 B.n23 VSUBS 0.008963f
C52 B.n24 VSUBS 0.008963f
C53 B.n25 VSUBS 0.008963f
C54 B.n26 VSUBS 0.008963f
C55 B.n27 VSUBS 0.008963f
C56 B.n28 VSUBS 0.008963f
C57 B.n29 VSUBS 0.008963f
C58 B.n30 VSUBS 0.02256f
C59 B.n31 VSUBS 0.008963f
C60 B.n32 VSUBS 0.008963f
C61 B.n33 VSUBS 0.008963f
C62 B.n34 VSUBS 0.008963f
C63 B.n35 VSUBS 0.008963f
C64 B.n36 VSUBS 0.008963f
C65 B.n37 VSUBS 0.008963f
C66 B.n38 VSUBS 0.008963f
C67 B.n39 VSUBS 0.008963f
C68 B.n40 VSUBS 0.008963f
C69 B.n41 VSUBS 0.008963f
C70 B.n42 VSUBS 0.008963f
C71 B.n43 VSUBS 0.008963f
C72 B.n44 VSUBS 0.008963f
C73 B.n45 VSUBS 0.008963f
C74 B.n46 VSUBS 0.008963f
C75 B.n47 VSUBS 0.008963f
C76 B.n48 VSUBS 0.008963f
C77 B.n49 VSUBS 0.008963f
C78 B.n50 VSUBS 0.008963f
C79 B.n51 VSUBS 0.008963f
C80 B.n52 VSUBS 0.008963f
C81 B.n53 VSUBS 0.008963f
C82 B.t11 VSUBS 0.583453f
C83 B.t10 VSUBS 0.608724f
C84 B.t9 VSUBS 1.89389f
C85 B.n54 VSUBS 0.313956f
C86 B.n55 VSUBS 0.090952f
C87 B.n56 VSUBS 0.008963f
C88 B.n57 VSUBS 0.008963f
C89 B.n58 VSUBS 0.008963f
C90 B.n59 VSUBS 0.008963f
C91 B.t2 VSUBS 0.583439f
C92 B.t1 VSUBS 0.608712f
C93 B.t0 VSUBS 1.89389f
C94 B.n60 VSUBS 0.313968f
C95 B.n61 VSUBS 0.090966f
C96 B.n62 VSUBS 0.020766f
C97 B.n63 VSUBS 0.008963f
C98 B.n64 VSUBS 0.008963f
C99 B.n65 VSUBS 0.008963f
C100 B.n66 VSUBS 0.008963f
C101 B.n67 VSUBS 0.008963f
C102 B.n68 VSUBS 0.008963f
C103 B.n69 VSUBS 0.008963f
C104 B.n70 VSUBS 0.008963f
C105 B.n71 VSUBS 0.008963f
C106 B.n72 VSUBS 0.008963f
C107 B.n73 VSUBS 0.008963f
C108 B.n74 VSUBS 0.008963f
C109 B.n75 VSUBS 0.008963f
C110 B.n76 VSUBS 0.008963f
C111 B.n77 VSUBS 0.008963f
C112 B.n78 VSUBS 0.008963f
C113 B.n79 VSUBS 0.008963f
C114 B.n80 VSUBS 0.008963f
C115 B.n81 VSUBS 0.008963f
C116 B.n82 VSUBS 0.008963f
C117 B.n83 VSUBS 0.008963f
C118 B.n84 VSUBS 0.008963f
C119 B.n85 VSUBS 0.008963f
C120 B.n86 VSUBS 0.022703f
C121 B.n87 VSUBS 0.008963f
C122 B.n88 VSUBS 0.008963f
C123 B.n89 VSUBS 0.008963f
C124 B.n90 VSUBS 0.008963f
C125 B.n91 VSUBS 0.008963f
C126 B.n92 VSUBS 0.008963f
C127 B.n93 VSUBS 0.008963f
C128 B.n94 VSUBS 0.008963f
C129 B.n95 VSUBS 0.008963f
C130 B.n96 VSUBS 0.008963f
C131 B.n97 VSUBS 0.008963f
C132 B.n98 VSUBS 0.008963f
C133 B.n99 VSUBS 0.008963f
C134 B.n100 VSUBS 0.008963f
C135 B.n101 VSUBS 0.008963f
C136 B.n102 VSUBS 0.008963f
C137 B.n103 VSUBS 0.008963f
C138 B.n104 VSUBS 0.008963f
C139 B.n105 VSUBS 0.008963f
C140 B.n106 VSUBS 0.008963f
C141 B.n107 VSUBS 0.008963f
C142 B.n108 VSUBS 0.008963f
C143 B.n109 VSUBS 0.008963f
C144 B.n110 VSUBS 0.008963f
C145 B.n111 VSUBS 0.008963f
C146 B.n112 VSUBS 0.008963f
C147 B.n113 VSUBS 0.008963f
C148 B.n114 VSUBS 0.008963f
C149 B.n115 VSUBS 0.008963f
C150 B.n116 VSUBS 0.008963f
C151 B.n117 VSUBS 0.008963f
C152 B.n118 VSUBS 0.008963f
C153 B.n119 VSUBS 0.008963f
C154 B.n120 VSUBS 0.008963f
C155 B.n121 VSUBS 0.008963f
C156 B.n122 VSUBS 0.008963f
C157 B.n123 VSUBS 0.008963f
C158 B.n124 VSUBS 0.008963f
C159 B.n125 VSUBS 0.008963f
C160 B.n126 VSUBS 0.008963f
C161 B.n127 VSUBS 0.008963f
C162 B.n128 VSUBS 0.008963f
C163 B.n129 VSUBS 0.008963f
C164 B.n130 VSUBS 0.008963f
C165 B.n131 VSUBS 0.008963f
C166 B.n132 VSUBS 0.008963f
C167 B.n133 VSUBS 0.008963f
C168 B.n134 VSUBS 0.008963f
C169 B.n135 VSUBS 0.008963f
C170 B.n136 VSUBS 0.008963f
C171 B.n137 VSUBS 0.008963f
C172 B.n138 VSUBS 0.008963f
C173 B.n139 VSUBS 0.008963f
C174 B.n140 VSUBS 0.008963f
C175 B.n141 VSUBS 0.008963f
C176 B.n142 VSUBS 0.021727f
C177 B.n143 VSUBS 0.008963f
C178 B.n144 VSUBS 0.008963f
C179 B.n145 VSUBS 0.008963f
C180 B.n146 VSUBS 0.008963f
C181 B.n147 VSUBS 0.008963f
C182 B.n148 VSUBS 0.008963f
C183 B.n149 VSUBS 0.008963f
C184 B.n150 VSUBS 0.008963f
C185 B.n151 VSUBS 0.008963f
C186 B.n152 VSUBS 0.008963f
C187 B.n153 VSUBS 0.008963f
C188 B.n154 VSUBS 0.008963f
C189 B.n155 VSUBS 0.008963f
C190 B.n156 VSUBS 0.008963f
C191 B.n157 VSUBS 0.008963f
C192 B.n158 VSUBS 0.008963f
C193 B.n159 VSUBS 0.008963f
C194 B.n160 VSUBS 0.008963f
C195 B.n161 VSUBS 0.008963f
C196 B.n162 VSUBS 0.008963f
C197 B.n163 VSUBS 0.008963f
C198 B.n164 VSUBS 0.008963f
C199 B.n165 VSUBS 0.008963f
C200 B.t7 VSUBS 0.583439f
C201 B.t8 VSUBS 0.608712f
C202 B.t6 VSUBS 1.89389f
C203 B.n166 VSUBS 0.313968f
C204 B.n167 VSUBS 0.090966f
C205 B.n168 VSUBS 0.020766f
C206 B.n169 VSUBS 0.008963f
C207 B.n170 VSUBS 0.008963f
C208 B.n171 VSUBS 0.008963f
C209 B.n172 VSUBS 0.008963f
C210 B.n173 VSUBS 0.008963f
C211 B.t4 VSUBS 0.583453f
C212 B.t5 VSUBS 0.608724f
C213 B.t3 VSUBS 1.89389f
C214 B.n174 VSUBS 0.313956f
C215 B.n175 VSUBS 0.090952f
C216 B.n176 VSUBS 0.008963f
C217 B.n177 VSUBS 0.008963f
C218 B.n178 VSUBS 0.008963f
C219 B.n179 VSUBS 0.008963f
C220 B.n180 VSUBS 0.008963f
C221 B.n181 VSUBS 0.008963f
C222 B.n182 VSUBS 0.008963f
C223 B.n183 VSUBS 0.008963f
C224 B.n184 VSUBS 0.008963f
C225 B.n185 VSUBS 0.008963f
C226 B.n186 VSUBS 0.008963f
C227 B.n187 VSUBS 0.008963f
C228 B.n188 VSUBS 0.008963f
C229 B.n189 VSUBS 0.008963f
C230 B.n190 VSUBS 0.008963f
C231 B.n191 VSUBS 0.008963f
C232 B.n192 VSUBS 0.008963f
C233 B.n193 VSUBS 0.008963f
C234 B.n194 VSUBS 0.008963f
C235 B.n195 VSUBS 0.008963f
C236 B.n196 VSUBS 0.008963f
C237 B.n197 VSUBS 0.008963f
C238 B.n198 VSUBS 0.02256f
C239 B.n199 VSUBS 0.008963f
C240 B.n200 VSUBS 0.008963f
C241 B.n201 VSUBS 0.008963f
C242 B.n202 VSUBS 0.008963f
C243 B.n203 VSUBS 0.008963f
C244 B.n204 VSUBS 0.008963f
C245 B.n205 VSUBS 0.008963f
C246 B.n206 VSUBS 0.008963f
C247 B.n207 VSUBS 0.008963f
C248 B.n208 VSUBS 0.008963f
C249 B.n209 VSUBS 0.008963f
C250 B.n210 VSUBS 0.008963f
C251 B.n211 VSUBS 0.008963f
C252 B.n212 VSUBS 0.008963f
C253 B.n213 VSUBS 0.008963f
C254 B.n214 VSUBS 0.008963f
C255 B.n215 VSUBS 0.008963f
C256 B.n216 VSUBS 0.008963f
C257 B.n217 VSUBS 0.008963f
C258 B.n218 VSUBS 0.008963f
C259 B.n219 VSUBS 0.008963f
C260 B.n220 VSUBS 0.008963f
C261 B.n221 VSUBS 0.008963f
C262 B.n222 VSUBS 0.008963f
C263 B.n223 VSUBS 0.008963f
C264 B.n224 VSUBS 0.008963f
C265 B.n225 VSUBS 0.008963f
C266 B.n226 VSUBS 0.008963f
C267 B.n227 VSUBS 0.008963f
C268 B.n228 VSUBS 0.008963f
C269 B.n229 VSUBS 0.008963f
C270 B.n230 VSUBS 0.008963f
C271 B.n231 VSUBS 0.008963f
C272 B.n232 VSUBS 0.008963f
C273 B.n233 VSUBS 0.008963f
C274 B.n234 VSUBS 0.008963f
C275 B.n235 VSUBS 0.008963f
C276 B.n236 VSUBS 0.008963f
C277 B.n237 VSUBS 0.008963f
C278 B.n238 VSUBS 0.008963f
C279 B.n239 VSUBS 0.008963f
C280 B.n240 VSUBS 0.008963f
C281 B.n241 VSUBS 0.008963f
C282 B.n242 VSUBS 0.008963f
C283 B.n243 VSUBS 0.008963f
C284 B.n244 VSUBS 0.008963f
C285 B.n245 VSUBS 0.008963f
C286 B.n246 VSUBS 0.008963f
C287 B.n247 VSUBS 0.008963f
C288 B.n248 VSUBS 0.008963f
C289 B.n249 VSUBS 0.008963f
C290 B.n250 VSUBS 0.008963f
C291 B.n251 VSUBS 0.008963f
C292 B.n252 VSUBS 0.008963f
C293 B.n253 VSUBS 0.008963f
C294 B.n254 VSUBS 0.008963f
C295 B.n255 VSUBS 0.008963f
C296 B.n256 VSUBS 0.008963f
C297 B.n257 VSUBS 0.008963f
C298 B.n258 VSUBS 0.008963f
C299 B.n259 VSUBS 0.008963f
C300 B.n260 VSUBS 0.008963f
C301 B.n261 VSUBS 0.008963f
C302 B.n262 VSUBS 0.008963f
C303 B.n263 VSUBS 0.008963f
C304 B.n264 VSUBS 0.008963f
C305 B.n265 VSUBS 0.008963f
C306 B.n266 VSUBS 0.008963f
C307 B.n267 VSUBS 0.008963f
C308 B.n268 VSUBS 0.008963f
C309 B.n269 VSUBS 0.008963f
C310 B.n270 VSUBS 0.008963f
C311 B.n271 VSUBS 0.008963f
C312 B.n272 VSUBS 0.008963f
C313 B.n273 VSUBS 0.008963f
C314 B.n274 VSUBS 0.008963f
C315 B.n275 VSUBS 0.008963f
C316 B.n276 VSUBS 0.008963f
C317 B.n277 VSUBS 0.008963f
C318 B.n278 VSUBS 0.008963f
C319 B.n279 VSUBS 0.008963f
C320 B.n280 VSUBS 0.008963f
C321 B.n281 VSUBS 0.008963f
C322 B.n282 VSUBS 0.008963f
C323 B.n283 VSUBS 0.008963f
C324 B.n284 VSUBS 0.008963f
C325 B.n285 VSUBS 0.008963f
C326 B.n286 VSUBS 0.008963f
C327 B.n287 VSUBS 0.008963f
C328 B.n288 VSUBS 0.008963f
C329 B.n289 VSUBS 0.008963f
C330 B.n290 VSUBS 0.008963f
C331 B.n291 VSUBS 0.008963f
C332 B.n292 VSUBS 0.008963f
C333 B.n293 VSUBS 0.008963f
C334 B.n294 VSUBS 0.008963f
C335 B.n295 VSUBS 0.008963f
C336 B.n296 VSUBS 0.008963f
C337 B.n297 VSUBS 0.008963f
C338 B.n298 VSUBS 0.008963f
C339 B.n299 VSUBS 0.008963f
C340 B.n300 VSUBS 0.008963f
C341 B.n301 VSUBS 0.008963f
C342 B.n302 VSUBS 0.008963f
C343 B.n303 VSUBS 0.008963f
C344 B.n304 VSUBS 0.008963f
C345 B.n305 VSUBS 0.008963f
C346 B.n306 VSUBS 0.008963f
C347 B.n307 VSUBS 0.021727f
C348 B.n308 VSUBS 0.021727f
C349 B.n309 VSUBS 0.02256f
C350 B.n310 VSUBS 0.008963f
C351 B.n311 VSUBS 0.008963f
C352 B.n312 VSUBS 0.008963f
C353 B.n313 VSUBS 0.008963f
C354 B.n314 VSUBS 0.008963f
C355 B.n315 VSUBS 0.008963f
C356 B.n316 VSUBS 0.008963f
C357 B.n317 VSUBS 0.008963f
C358 B.n318 VSUBS 0.008963f
C359 B.n319 VSUBS 0.008963f
C360 B.n320 VSUBS 0.008963f
C361 B.n321 VSUBS 0.008963f
C362 B.n322 VSUBS 0.008963f
C363 B.n323 VSUBS 0.008963f
C364 B.n324 VSUBS 0.008963f
C365 B.n325 VSUBS 0.008963f
C366 B.n326 VSUBS 0.008963f
C367 B.n327 VSUBS 0.008963f
C368 B.n328 VSUBS 0.008963f
C369 B.n329 VSUBS 0.008963f
C370 B.n330 VSUBS 0.008963f
C371 B.n331 VSUBS 0.008963f
C372 B.n332 VSUBS 0.008963f
C373 B.n333 VSUBS 0.008963f
C374 B.n334 VSUBS 0.008963f
C375 B.n335 VSUBS 0.008963f
C376 B.n336 VSUBS 0.008963f
C377 B.n337 VSUBS 0.008963f
C378 B.n338 VSUBS 0.008963f
C379 B.n339 VSUBS 0.008963f
C380 B.n340 VSUBS 0.008963f
C381 B.n341 VSUBS 0.008963f
C382 B.n342 VSUBS 0.008963f
C383 B.n343 VSUBS 0.008963f
C384 B.n344 VSUBS 0.008963f
C385 B.n345 VSUBS 0.008963f
C386 B.n346 VSUBS 0.008963f
C387 B.n347 VSUBS 0.008963f
C388 B.n348 VSUBS 0.008963f
C389 B.n349 VSUBS 0.008963f
C390 B.n350 VSUBS 0.008963f
C391 B.n351 VSUBS 0.008963f
C392 B.n352 VSUBS 0.008963f
C393 B.n353 VSUBS 0.008963f
C394 B.n354 VSUBS 0.008963f
C395 B.n355 VSUBS 0.008963f
C396 B.n356 VSUBS 0.008963f
C397 B.n357 VSUBS 0.008963f
C398 B.n358 VSUBS 0.008963f
C399 B.n359 VSUBS 0.008963f
C400 B.n360 VSUBS 0.008963f
C401 B.n361 VSUBS 0.008963f
C402 B.n362 VSUBS 0.008963f
C403 B.n363 VSUBS 0.008963f
C404 B.n364 VSUBS 0.008963f
C405 B.n365 VSUBS 0.008963f
C406 B.n366 VSUBS 0.008963f
C407 B.n367 VSUBS 0.008963f
C408 B.n368 VSUBS 0.008963f
C409 B.n369 VSUBS 0.008963f
C410 B.n370 VSUBS 0.008963f
C411 B.n371 VSUBS 0.008963f
C412 B.n372 VSUBS 0.008963f
C413 B.n373 VSUBS 0.008963f
C414 B.n374 VSUBS 0.008963f
C415 B.n375 VSUBS 0.008963f
C416 B.n376 VSUBS 0.008963f
C417 B.n377 VSUBS 0.008963f
C418 B.n378 VSUBS 0.006195f
C419 B.n379 VSUBS 0.020766f
C420 B.n380 VSUBS 0.007249f
C421 B.n381 VSUBS 0.008963f
C422 B.n382 VSUBS 0.008963f
C423 B.n383 VSUBS 0.008963f
C424 B.n384 VSUBS 0.008963f
C425 B.n385 VSUBS 0.008963f
C426 B.n386 VSUBS 0.008963f
C427 B.n387 VSUBS 0.008963f
C428 B.n388 VSUBS 0.008963f
C429 B.n389 VSUBS 0.008963f
C430 B.n390 VSUBS 0.008963f
C431 B.n391 VSUBS 0.008963f
C432 B.n392 VSUBS 0.007249f
C433 B.n393 VSUBS 0.008963f
C434 B.n394 VSUBS 0.008963f
C435 B.n395 VSUBS 0.006195f
C436 B.n396 VSUBS 0.008963f
C437 B.n397 VSUBS 0.008963f
C438 B.n398 VSUBS 0.008963f
C439 B.n399 VSUBS 0.008963f
C440 B.n400 VSUBS 0.008963f
C441 B.n401 VSUBS 0.008963f
C442 B.n402 VSUBS 0.008963f
C443 B.n403 VSUBS 0.008963f
C444 B.n404 VSUBS 0.008963f
C445 B.n405 VSUBS 0.008963f
C446 B.n406 VSUBS 0.008963f
C447 B.n407 VSUBS 0.008963f
C448 B.n408 VSUBS 0.008963f
C449 B.n409 VSUBS 0.008963f
C450 B.n410 VSUBS 0.008963f
C451 B.n411 VSUBS 0.008963f
C452 B.n412 VSUBS 0.008963f
C453 B.n413 VSUBS 0.008963f
C454 B.n414 VSUBS 0.008963f
C455 B.n415 VSUBS 0.008963f
C456 B.n416 VSUBS 0.008963f
C457 B.n417 VSUBS 0.008963f
C458 B.n418 VSUBS 0.008963f
C459 B.n419 VSUBS 0.008963f
C460 B.n420 VSUBS 0.008963f
C461 B.n421 VSUBS 0.008963f
C462 B.n422 VSUBS 0.008963f
C463 B.n423 VSUBS 0.008963f
C464 B.n424 VSUBS 0.008963f
C465 B.n425 VSUBS 0.008963f
C466 B.n426 VSUBS 0.008963f
C467 B.n427 VSUBS 0.008963f
C468 B.n428 VSUBS 0.008963f
C469 B.n429 VSUBS 0.008963f
C470 B.n430 VSUBS 0.008963f
C471 B.n431 VSUBS 0.008963f
C472 B.n432 VSUBS 0.008963f
C473 B.n433 VSUBS 0.008963f
C474 B.n434 VSUBS 0.008963f
C475 B.n435 VSUBS 0.008963f
C476 B.n436 VSUBS 0.008963f
C477 B.n437 VSUBS 0.008963f
C478 B.n438 VSUBS 0.008963f
C479 B.n439 VSUBS 0.008963f
C480 B.n440 VSUBS 0.008963f
C481 B.n441 VSUBS 0.008963f
C482 B.n442 VSUBS 0.008963f
C483 B.n443 VSUBS 0.008963f
C484 B.n444 VSUBS 0.008963f
C485 B.n445 VSUBS 0.008963f
C486 B.n446 VSUBS 0.008963f
C487 B.n447 VSUBS 0.008963f
C488 B.n448 VSUBS 0.008963f
C489 B.n449 VSUBS 0.008963f
C490 B.n450 VSUBS 0.008963f
C491 B.n451 VSUBS 0.008963f
C492 B.n452 VSUBS 0.008963f
C493 B.n453 VSUBS 0.008963f
C494 B.n454 VSUBS 0.008963f
C495 B.n455 VSUBS 0.008963f
C496 B.n456 VSUBS 0.008963f
C497 B.n457 VSUBS 0.008963f
C498 B.n458 VSUBS 0.008963f
C499 B.n459 VSUBS 0.008963f
C500 B.n460 VSUBS 0.008963f
C501 B.n461 VSUBS 0.008963f
C502 B.n462 VSUBS 0.008963f
C503 B.n463 VSUBS 0.02256f
C504 B.n464 VSUBS 0.02256f
C505 B.n465 VSUBS 0.021727f
C506 B.n466 VSUBS 0.008963f
C507 B.n467 VSUBS 0.008963f
C508 B.n468 VSUBS 0.008963f
C509 B.n469 VSUBS 0.008963f
C510 B.n470 VSUBS 0.008963f
C511 B.n471 VSUBS 0.008963f
C512 B.n472 VSUBS 0.008963f
C513 B.n473 VSUBS 0.008963f
C514 B.n474 VSUBS 0.008963f
C515 B.n475 VSUBS 0.008963f
C516 B.n476 VSUBS 0.008963f
C517 B.n477 VSUBS 0.008963f
C518 B.n478 VSUBS 0.008963f
C519 B.n479 VSUBS 0.008963f
C520 B.n480 VSUBS 0.008963f
C521 B.n481 VSUBS 0.008963f
C522 B.n482 VSUBS 0.008963f
C523 B.n483 VSUBS 0.008963f
C524 B.n484 VSUBS 0.008963f
C525 B.n485 VSUBS 0.008963f
C526 B.n486 VSUBS 0.008963f
C527 B.n487 VSUBS 0.008963f
C528 B.n488 VSUBS 0.008963f
C529 B.n489 VSUBS 0.008963f
C530 B.n490 VSUBS 0.008963f
C531 B.n491 VSUBS 0.008963f
C532 B.n492 VSUBS 0.008963f
C533 B.n493 VSUBS 0.008963f
C534 B.n494 VSUBS 0.008963f
C535 B.n495 VSUBS 0.008963f
C536 B.n496 VSUBS 0.008963f
C537 B.n497 VSUBS 0.008963f
C538 B.n498 VSUBS 0.008963f
C539 B.n499 VSUBS 0.008963f
C540 B.n500 VSUBS 0.008963f
C541 B.n501 VSUBS 0.008963f
C542 B.n502 VSUBS 0.008963f
C543 B.n503 VSUBS 0.008963f
C544 B.n504 VSUBS 0.008963f
C545 B.n505 VSUBS 0.008963f
C546 B.n506 VSUBS 0.008963f
C547 B.n507 VSUBS 0.008963f
C548 B.n508 VSUBS 0.008963f
C549 B.n509 VSUBS 0.008963f
C550 B.n510 VSUBS 0.008963f
C551 B.n511 VSUBS 0.008963f
C552 B.n512 VSUBS 0.008963f
C553 B.n513 VSUBS 0.008963f
C554 B.n514 VSUBS 0.008963f
C555 B.n515 VSUBS 0.008963f
C556 B.n516 VSUBS 0.008963f
C557 B.n517 VSUBS 0.008963f
C558 B.n518 VSUBS 0.008963f
C559 B.n519 VSUBS 0.008963f
C560 B.n520 VSUBS 0.008963f
C561 B.n521 VSUBS 0.008963f
C562 B.n522 VSUBS 0.008963f
C563 B.n523 VSUBS 0.008963f
C564 B.n524 VSUBS 0.008963f
C565 B.n525 VSUBS 0.008963f
C566 B.n526 VSUBS 0.008963f
C567 B.n527 VSUBS 0.008963f
C568 B.n528 VSUBS 0.008963f
C569 B.n529 VSUBS 0.008963f
C570 B.n530 VSUBS 0.008963f
C571 B.n531 VSUBS 0.008963f
C572 B.n532 VSUBS 0.008963f
C573 B.n533 VSUBS 0.008963f
C574 B.n534 VSUBS 0.008963f
C575 B.n535 VSUBS 0.008963f
C576 B.n536 VSUBS 0.008963f
C577 B.n537 VSUBS 0.008963f
C578 B.n538 VSUBS 0.008963f
C579 B.n539 VSUBS 0.008963f
C580 B.n540 VSUBS 0.008963f
C581 B.n541 VSUBS 0.008963f
C582 B.n542 VSUBS 0.008963f
C583 B.n543 VSUBS 0.008963f
C584 B.n544 VSUBS 0.008963f
C585 B.n545 VSUBS 0.008963f
C586 B.n546 VSUBS 0.008963f
C587 B.n547 VSUBS 0.008963f
C588 B.n548 VSUBS 0.008963f
C589 B.n549 VSUBS 0.008963f
C590 B.n550 VSUBS 0.008963f
C591 B.n551 VSUBS 0.008963f
C592 B.n552 VSUBS 0.008963f
C593 B.n553 VSUBS 0.008963f
C594 B.n554 VSUBS 0.008963f
C595 B.n555 VSUBS 0.008963f
C596 B.n556 VSUBS 0.008963f
C597 B.n557 VSUBS 0.008963f
C598 B.n558 VSUBS 0.008963f
C599 B.n559 VSUBS 0.008963f
C600 B.n560 VSUBS 0.008963f
C601 B.n561 VSUBS 0.008963f
C602 B.n562 VSUBS 0.008963f
C603 B.n563 VSUBS 0.008963f
C604 B.n564 VSUBS 0.008963f
C605 B.n565 VSUBS 0.008963f
C606 B.n566 VSUBS 0.008963f
C607 B.n567 VSUBS 0.008963f
C608 B.n568 VSUBS 0.008963f
C609 B.n569 VSUBS 0.008963f
C610 B.n570 VSUBS 0.008963f
C611 B.n571 VSUBS 0.008963f
C612 B.n572 VSUBS 0.008963f
C613 B.n573 VSUBS 0.008963f
C614 B.n574 VSUBS 0.008963f
C615 B.n575 VSUBS 0.008963f
C616 B.n576 VSUBS 0.008963f
C617 B.n577 VSUBS 0.008963f
C618 B.n578 VSUBS 0.008963f
C619 B.n579 VSUBS 0.008963f
C620 B.n580 VSUBS 0.008963f
C621 B.n581 VSUBS 0.008963f
C622 B.n582 VSUBS 0.008963f
C623 B.n583 VSUBS 0.008963f
C624 B.n584 VSUBS 0.008963f
C625 B.n585 VSUBS 0.008963f
C626 B.n586 VSUBS 0.008963f
C627 B.n587 VSUBS 0.008963f
C628 B.n588 VSUBS 0.008963f
C629 B.n589 VSUBS 0.008963f
C630 B.n590 VSUBS 0.008963f
C631 B.n591 VSUBS 0.008963f
C632 B.n592 VSUBS 0.008963f
C633 B.n593 VSUBS 0.008963f
C634 B.n594 VSUBS 0.008963f
C635 B.n595 VSUBS 0.008963f
C636 B.n596 VSUBS 0.008963f
C637 B.n597 VSUBS 0.008963f
C638 B.n598 VSUBS 0.008963f
C639 B.n599 VSUBS 0.008963f
C640 B.n600 VSUBS 0.008963f
C641 B.n601 VSUBS 0.008963f
C642 B.n602 VSUBS 0.008963f
C643 B.n603 VSUBS 0.008963f
C644 B.n604 VSUBS 0.008963f
C645 B.n605 VSUBS 0.008963f
C646 B.n606 VSUBS 0.008963f
C647 B.n607 VSUBS 0.008963f
C648 B.n608 VSUBS 0.008963f
C649 B.n609 VSUBS 0.008963f
C650 B.n610 VSUBS 0.008963f
C651 B.n611 VSUBS 0.008963f
C652 B.n612 VSUBS 0.008963f
C653 B.n613 VSUBS 0.008963f
C654 B.n614 VSUBS 0.008963f
C655 B.n615 VSUBS 0.008963f
C656 B.n616 VSUBS 0.008963f
C657 B.n617 VSUBS 0.008963f
C658 B.n618 VSUBS 0.008963f
C659 B.n619 VSUBS 0.008963f
C660 B.n620 VSUBS 0.008963f
C661 B.n621 VSUBS 0.008963f
C662 B.n622 VSUBS 0.008963f
C663 B.n623 VSUBS 0.008963f
C664 B.n624 VSUBS 0.008963f
C665 B.n625 VSUBS 0.008963f
C666 B.n626 VSUBS 0.008963f
C667 B.n627 VSUBS 0.008963f
C668 B.n628 VSUBS 0.008963f
C669 B.n629 VSUBS 0.008963f
C670 B.n630 VSUBS 0.008963f
C671 B.n631 VSUBS 0.008963f
C672 B.n632 VSUBS 0.008963f
C673 B.n633 VSUBS 0.021727f
C674 B.n634 VSUBS 0.02256f
C675 B.n635 VSUBS 0.021584f
C676 B.n636 VSUBS 0.008963f
C677 B.n637 VSUBS 0.008963f
C678 B.n638 VSUBS 0.008963f
C679 B.n639 VSUBS 0.008963f
C680 B.n640 VSUBS 0.008963f
C681 B.n641 VSUBS 0.008963f
C682 B.n642 VSUBS 0.008963f
C683 B.n643 VSUBS 0.008963f
C684 B.n644 VSUBS 0.008963f
C685 B.n645 VSUBS 0.008963f
C686 B.n646 VSUBS 0.008963f
C687 B.n647 VSUBS 0.008963f
C688 B.n648 VSUBS 0.008963f
C689 B.n649 VSUBS 0.008963f
C690 B.n650 VSUBS 0.008963f
C691 B.n651 VSUBS 0.008963f
C692 B.n652 VSUBS 0.008963f
C693 B.n653 VSUBS 0.008963f
C694 B.n654 VSUBS 0.008963f
C695 B.n655 VSUBS 0.008963f
C696 B.n656 VSUBS 0.008963f
C697 B.n657 VSUBS 0.008963f
C698 B.n658 VSUBS 0.008963f
C699 B.n659 VSUBS 0.008963f
C700 B.n660 VSUBS 0.008963f
C701 B.n661 VSUBS 0.008963f
C702 B.n662 VSUBS 0.008963f
C703 B.n663 VSUBS 0.008963f
C704 B.n664 VSUBS 0.008963f
C705 B.n665 VSUBS 0.008963f
C706 B.n666 VSUBS 0.008963f
C707 B.n667 VSUBS 0.008963f
C708 B.n668 VSUBS 0.008963f
C709 B.n669 VSUBS 0.008963f
C710 B.n670 VSUBS 0.008963f
C711 B.n671 VSUBS 0.008963f
C712 B.n672 VSUBS 0.008963f
C713 B.n673 VSUBS 0.008963f
C714 B.n674 VSUBS 0.008963f
C715 B.n675 VSUBS 0.008963f
C716 B.n676 VSUBS 0.008963f
C717 B.n677 VSUBS 0.008963f
C718 B.n678 VSUBS 0.008963f
C719 B.n679 VSUBS 0.008963f
C720 B.n680 VSUBS 0.008963f
C721 B.n681 VSUBS 0.008963f
C722 B.n682 VSUBS 0.008963f
C723 B.n683 VSUBS 0.008963f
C724 B.n684 VSUBS 0.008963f
C725 B.n685 VSUBS 0.008963f
C726 B.n686 VSUBS 0.008963f
C727 B.n687 VSUBS 0.008963f
C728 B.n688 VSUBS 0.008963f
C729 B.n689 VSUBS 0.008963f
C730 B.n690 VSUBS 0.008963f
C731 B.n691 VSUBS 0.008963f
C732 B.n692 VSUBS 0.008963f
C733 B.n693 VSUBS 0.008963f
C734 B.n694 VSUBS 0.008963f
C735 B.n695 VSUBS 0.008963f
C736 B.n696 VSUBS 0.008963f
C737 B.n697 VSUBS 0.008963f
C738 B.n698 VSUBS 0.008963f
C739 B.n699 VSUBS 0.008963f
C740 B.n700 VSUBS 0.008963f
C741 B.n701 VSUBS 0.008963f
C742 B.n702 VSUBS 0.008963f
C743 B.n703 VSUBS 0.006195f
C744 B.n704 VSUBS 0.008963f
C745 B.n705 VSUBS 0.008963f
C746 B.n706 VSUBS 0.007249f
C747 B.n707 VSUBS 0.008963f
C748 B.n708 VSUBS 0.008963f
C749 B.n709 VSUBS 0.008963f
C750 B.n710 VSUBS 0.008963f
C751 B.n711 VSUBS 0.008963f
C752 B.n712 VSUBS 0.008963f
C753 B.n713 VSUBS 0.008963f
C754 B.n714 VSUBS 0.008963f
C755 B.n715 VSUBS 0.008963f
C756 B.n716 VSUBS 0.008963f
C757 B.n717 VSUBS 0.008963f
C758 B.n718 VSUBS 0.007249f
C759 B.n719 VSUBS 0.020766f
C760 B.n720 VSUBS 0.006195f
C761 B.n721 VSUBS 0.008963f
C762 B.n722 VSUBS 0.008963f
C763 B.n723 VSUBS 0.008963f
C764 B.n724 VSUBS 0.008963f
C765 B.n725 VSUBS 0.008963f
C766 B.n726 VSUBS 0.008963f
C767 B.n727 VSUBS 0.008963f
C768 B.n728 VSUBS 0.008963f
C769 B.n729 VSUBS 0.008963f
C770 B.n730 VSUBS 0.008963f
C771 B.n731 VSUBS 0.008963f
C772 B.n732 VSUBS 0.008963f
C773 B.n733 VSUBS 0.008963f
C774 B.n734 VSUBS 0.008963f
C775 B.n735 VSUBS 0.008963f
C776 B.n736 VSUBS 0.008963f
C777 B.n737 VSUBS 0.008963f
C778 B.n738 VSUBS 0.008963f
C779 B.n739 VSUBS 0.008963f
C780 B.n740 VSUBS 0.008963f
C781 B.n741 VSUBS 0.008963f
C782 B.n742 VSUBS 0.008963f
C783 B.n743 VSUBS 0.008963f
C784 B.n744 VSUBS 0.008963f
C785 B.n745 VSUBS 0.008963f
C786 B.n746 VSUBS 0.008963f
C787 B.n747 VSUBS 0.008963f
C788 B.n748 VSUBS 0.008963f
C789 B.n749 VSUBS 0.008963f
C790 B.n750 VSUBS 0.008963f
C791 B.n751 VSUBS 0.008963f
C792 B.n752 VSUBS 0.008963f
C793 B.n753 VSUBS 0.008963f
C794 B.n754 VSUBS 0.008963f
C795 B.n755 VSUBS 0.008963f
C796 B.n756 VSUBS 0.008963f
C797 B.n757 VSUBS 0.008963f
C798 B.n758 VSUBS 0.008963f
C799 B.n759 VSUBS 0.008963f
C800 B.n760 VSUBS 0.008963f
C801 B.n761 VSUBS 0.008963f
C802 B.n762 VSUBS 0.008963f
C803 B.n763 VSUBS 0.008963f
C804 B.n764 VSUBS 0.008963f
C805 B.n765 VSUBS 0.008963f
C806 B.n766 VSUBS 0.008963f
C807 B.n767 VSUBS 0.008963f
C808 B.n768 VSUBS 0.008963f
C809 B.n769 VSUBS 0.008963f
C810 B.n770 VSUBS 0.008963f
C811 B.n771 VSUBS 0.008963f
C812 B.n772 VSUBS 0.008963f
C813 B.n773 VSUBS 0.008963f
C814 B.n774 VSUBS 0.008963f
C815 B.n775 VSUBS 0.008963f
C816 B.n776 VSUBS 0.008963f
C817 B.n777 VSUBS 0.008963f
C818 B.n778 VSUBS 0.008963f
C819 B.n779 VSUBS 0.008963f
C820 B.n780 VSUBS 0.008963f
C821 B.n781 VSUBS 0.008963f
C822 B.n782 VSUBS 0.008963f
C823 B.n783 VSUBS 0.008963f
C824 B.n784 VSUBS 0.008963f
C825 B.n785 VSUBS 0.008963f
C826 B.n786 VSUBS 0.008963f
C827 B.n787 VSUBS 0.008963f
C828 B.n788 VSUBS 0.008963f
C829 B.n789 VSUBS 0.02256f
C830 B.n790 VSUBS 0.021727f
C831 B.n791 VSUBS 0.021727f
C832 B.n792 VSUBS 0.008963f
C833 B.n793 VSUBS 0.008963f
C834 B.n794 VSUBS 0.008963f
C835 B.n795 VSUBS 0.008963f
C836 B.n796 VSUBS 0.008963f
C837 B.n797 VSUBS 0.008963f
C838 B.n798 VSUBS 0.008963f
C839 B.n799 VSUBS 0.008963f
C840 B.n800 VSUBS 0.008963f
C841 B.n801 VSUBS 0.008963f
C842 B.n802 VSUBS 0.008963f
C843 B.n803 VSUBS 0.008963f
C844 B.n804 VSUBS 0.008963f
C845 B.n805 VSUBS 0.008963f
C846 B.n806 VSUBS 0.008963f
C847 B.n807 VSUBS 0.008963f
C848 B.n808 VSUBS 0.008963f
C849 B.n809 VSUBS 0.008963f
C850 B.n810 VSUBS 0.008963f
C851 B.n811 VSUBS 0.008963f
C852 B.n812 VSUBS 0.008963f
C853 B.n813 VSUBS 0.008963f
C854 B.n814 VSUBS 0.008963f
C855 B.n815 VSUBS 0.008963f
C856 B.n816 VSUBS 0.008963f
C857 B.n817 VSUBS 0.008963f
C858 B.n818 VSUBS 0.008963f
C859 B.n819 VSUBS 0.008963f
C860 B.n820 VSUBS 0.008963f
C861 B.n821 VSUBS 0.008963f
C862 B.n822 VSUBS 0.008963f
C863 B.n823 VSUBS 0.008963f
C864 B.n824 VSUBS 0.008963f
C865 B.n825 VSUBS 0.008963f
C866 B.n826 VSUBS 0.008963f
C867 B.n827 VSUBS 0.008963f
C868 B.n828 VSUBS 0.008963f
C869 B.n829 VSUBS 0.008963f
C870 B.n830 VSUBS 0.008963f
C871 B.n831 VSUBS 0.008963f
C872 B.n832 VSUBS 0.008963f
C873 B.n833 VSUBS 0.008963f
C874 B.n834 VSUBS 0.008963f
C875 B.n835 VSUBS 0.008963f
C876 B.n836 VSUBS 0.008963f
C877 B.n837 VSUBS 0.008963f
C878 B.n838 VSUBS 0.008963f
C879 B.n839 VSUBS 0.008963f
C880 B.n840 VSUBS 0.008963f
C881 B.n841 VSUBS 0.008963f
C882 B.n842 VSUBS 0.008963f
C883 B.n843 VSUBS 0.008963f
C884 B.n844 VSUBS 0.008963f
C885 B.n845 VSUBS 0.008963f
C886 B.n846 VSUBS 0.008963f
C887 B.n847 VSUBS 0.008963f
C888 B.n848 VSUBS 0.008963f
C889 B.n849 VSUBS 0.008963f
C890 B.n850 VSUBS 0.008963f
C891 B.n851 VSUBS 0.008963f
C892 B.n852 VSUBS 0.008963f
C893 B.n853 VSUBS 0.008963f
C894 B.n854 VSUBS 0.008963f
C895 B.n855 VSUBS 0.008963f
C896 B.n856 VSUBS 0.008963f
C897 B.n857 VSUBS 0.008963f
C898 B.n858 VSUBS 0.008963f
C899 B.n859 VSUBS 0.008963f
C900 B.n860 VSUBS 0.008963f
C901 B.n861 VSUBS 0.008963f
C902 B.n862 VSUBS 0.008963f
C903 B.n863 VSUBS 0.008963f
C904 B.n864 VSUBS 0.008963f
C905 B.n865 VSUBS 0.008963f
C906 B.n866 VSUBS 0.008963f
C907 B.n867 VSUBS 0.008963f
C908 B.n868 VSUBS 0.008963f
C909 B.n869 VSUBS 0.008963f
C910 B.n870 VSUBS 0.008963f
C911 B.n871 VSUBS 0.008963f
C912 B.n872 VSUBS 0.008963f
C913 B.n873 VSUBS 0.008963f
C914 B.n874 VSUBS 0.008963f
C915 B.n875 VSUBS 0.020295f
C916 VDD2.t6 VSUBS 3.37263f
C917 VDD2.t5 VSUBS 0.318614f
C918 VDD2.t9 VSUBS 0.318614f
C919 VDD2.n0 VSUBS 2.57254f
C920 VDD2.n1 VSUBS 1.64078f
C921 VDD2.t8 VSUBS 0.318614f
C922 VDD2.t2 VSUBS 0.318614f
C923 VDD2.n2 VSUBS 2.59284f
C924 VDD2.n3 VSUBS 3.68871f
C925 VDD2.t1 VSUBS 3.34768f
C926 VDD2.n4 VSUBS 4.02837f
C927 VDD2.t4 VSUBS 0.318614f
C928 VDD2.t7 VSUBS 0.318614f
C929 VDD2.n5 VSUBS 2.57255f
C930 VDD2.n6 VSUBS 0.815133f
C931 VDD2.t0 VSUBS 0.318614f
C932 VDD2.t3 VSUBS 0.318614f
C933 VDD2.n7 VSUBS 2.59279f
C934 VN.n0 VSUBS 0.037416f
C935 VN.t7 VSUBS 2.55794f
C936 VN.n1 VSUBS 0.035103f
C937 VN.n2 VSUBS 0.02838f
C938 VN.t1 VSUBS 2.55794f
C939 VN.n3 VSUBS 0.89988f
C940 VN.n4 VSUBS 0.02838f
C941 VN.n5 VSUBS 0.056542f
C942 VN.n6 VSUBS 0.02838f
C943 VN.t0 VSUBS 2.55794f
C944 VN.n7 VSUBS 0.027683f
C945 VN.n8 VSUBS 0.268273f
C946 VN.t4 VSUBS 2.55794f
C947 VN.t3 VSUBS 2.76428f
C948 VN.n9 VSUBS 0.957893f
C949 VN.n10 VSUBS 0.991056f
C950 VN.n11 VSUBS 0.051327f
C951 VN.n12 VSUBS 0.051528f
C952 VN.n13 VSUBS 0.02838f
C953 VN.n14 VSUBS 0.02838f
C954 VN.n15 VSUBS 0.02838f
C955 VN.n16 VSUBS 0.056542f
C956 VN.n17 VSUBS 0.039836f
C957 VN.n18 VSUBS 0.89988f
C958 VN.n19 VSUBS 0.039836f
C959 VN.n20 VSUBS 0.02838f
C960 VN.n21 VSUBS 0.02838f
C961 VN.n22 VSUBS 0.02838f
C962 VN.n23 VSUBS 0.027683f
C963 VN.n24 VSUBS 0.051528f
C964 VN.n25 VSUBS 0.051327f
C965 VN.n26 VSUBS 0.02838f
C966 VN.n27 VSUBS 0.02838f
C967 VN.n28 VSUBS 0.028346f
C968 VN.n29 VSUBS 0.052893f
C969 VN.n30 VSUBS 0.047757f
C970 VN.n31 VSUBS 0.02838f
C971 VN.n32 VSUBS 0.02838f
C972 VN.n33 VSUBS 0.02838f
C973 VN.n34 VSUBS 0.052893f
C974 VN.n35 VSUBS 0.036703f
C975 VN.n36 VSUBS 0.985899f
C976 VN.n37 VSUBS 0.044769f
C977 VN.n38 VSUBS 0.037416f
C978 VN.t8 VSUBS 2.55794f
C979 VN.n39 VSUBS 0.035103f
C980 VN.n40 VSUBS 0.02838f
C981 VN.t5 VSUBS 2.55794f
C982 VN.n41 VSUBS 0.89988f
C983 VN.n42 VSUBS 0.02838f
C984 VN.n43 VSUBS 0.056542f
C985 VN.n44 VSUBS 0.02838f
C986 VN.t2 VSUBS 2.55794f
C987 VN.n45 VSUBS 0.027683f
C988 VN.n46 VSUBS 0.268273f
C989 VN.t9 VSUBS 2.55794f
C990 VN.t6 VSUBS 2.76428f
C991 VN.n47 VSUBS 0.957893f
C992 VN.n48 VSUBS 0.991056f
C993 VN.n49 VSUBS 0.051327f
C994 VN.n50 VSUBS 0.051528f
C995 VN.n51 VSUBS 0.02838f
C996 VN.n52 VSUBS 0.02838f
C997 VN.n53 VSUBS 0.02838f
C998 VN.n54 VSUBS 0.056542f
C999 VN.n55 VSUBS 0.039836f
C1000 VN.n56 VSUBS 0.89988f
C1001 VN.n57 VSUBS 0.039836f
C1002 VN.n58 VSUBS 0.02838f
C1003 VN.n59 VSUBS 0.02838f
C1004 VN.n60 VSUBS 0.02838f
C1005 VN.n61 VSUBS 0.027683f
C1006 VN.n62 VSUBS 0.051528f
C1007 VN.n63 VSUBS 0.051327f
C1008 VN.n64 VSUBS 0.02838f
C1009 VN.n65 VSUBS 0.02838f
C1010 VN.n66 VSUBS 0.028346f
C1011 VN.n67 VSUBS 0.052893f
C1012 VN.n68 VSUBS 0.047757f
C1013 VN.n69 VSUBS 0.02838f
C1014 VN.n70 VSUBS 0.02838f
C1015 VN.n71 VSUBS 0.02838f
C1016 VN.n72 VSUBS 0.052893f
C1017 VN.n73 VSUBS 0.036703f
C1018 VN.n74 VSUBS 0.985899f
C1019 VN.n75 VSUBS 1.74441f
C1020 VDD1.t9 VSUBS 3.36089f
C1021 VDD1.t6 VSUBS 0.317505f
C1022 VDD1.t3 VSUBS 0.317505f
C1023 VDD1.n0 VSUBS 2.56359f
C1024 VDD1.n1 VSUBS 1.64445f
C1025 VDD1.t1 VSUBS 3.36088f
C1026 VDD1.t7 VSUBS 0.317505f
C1027 VDD1.t0 VSUBS 0.317505f
C1028 VDD1.n2 VSUBS 2.56358f
C1029 VDD1.n3 VSUBS 1.63507f
C1030 VDD1.t5 VSUBS 0.317505f
C1031 VDD1.t8 VSUBS 0.317505f
C1032 VDD1.n4 VSUBS 2.58381f
C1033 VDD1.n5 VSUBS 3.8164f
C1034 VDD1.t4 VSUBS 0.317505f
C1035 VDD1.t2 VSUBS 0.317505f
C1036 VDD1.n6 VSUBS 2.56358f
C1037 VDD1.n7 VSUBS 4.04757f
C1038 VTAIL.t3 VSUBS 0.306764f
C1039 VTAIL.t4 VSUBS 0.306764f
C1040 VTAIL.n0 VSUBS 2.33419f
C1041 VTAIL.n1 VSUBS 0.931844f
C1042 VTAIL.t12 VSUBS 3.06155f
C1043 VTAIL.n2 VSUBS 1.08901f
C1044 VTAIL.t11 VSUBS 0.306764f
C1045 VTAIL.t15 VSUBS 0.306764f
C1046 VTAIL.n3 VSUBS 2.33419f
C1047 VTAIL.n4 VSUBS 1.04347f
C1048 VTAIL.t10 VSUBS 0.306764f
C1049 VTAIL.t9 VSUBS 0.306764f
C1050 VTAIL.n5 VSUBS 2.33419f
C1051 VTAIL.n6 VSUBS 2.71688f
C1052 VTAIL.t2 VSUBS 0.306764f
C1053 VTAIL.t5 VSUBS 0.306764f
C1054 VTAIL.n7 VSUBS 2.3342f
C1055 VTAIL.n8 VSUBS 2.71687f
C1056 VTAIL.t1 VSUBS 0.306764f
C1057 VTAIL.t0 VSUBS 0.306764f
C1058 VTAIL.n9 VSUBS 2.3342f
C1059 VTAIL.n10 VSUBS 1.04346f
C1060 VTAIL.t17 VSUBS 3.06155f
C1061 VTAIL.n11 VSUBS 1.08901f
C1062 VTAIL.t7 VSUBS 0.306764f
C1063 VTAIL.t8 VSUBS 0.306764f
C1064 VTAIL.n12 VSUBS 2.3342f
C1065 VTAIL.n13 VSUBS 0.979735f
C1066 VTAIL.t13 VSUBS 0.306764f
C1067 VTAIL.t14 VSUBS 0.306764f
C1068 VTAIL.n14 VSUBS 2.3342f
C1069 VTAIL.n15 VSUBS 1.04346f
C1070 VTAIL.t16 VSUBS 3.06155f
C1071 VTAIL.n16 VSUBS 2.61346f
C1072 VTAIL.t18 VSUBS 3.06155f
C1073 VTAIL.n17 VSUBS 2.61346f
C1074 VTAIL.t6 VSUBS 0.306764f
C1075 VTAIL.t19 VSUBS 0.306764f
C1076 VTAIL.n18 VSUBS 2.33419f
C1077 VTAIL.n19 VSUBS 0.878671f
C1078 VP.n0 VSUBS 0.040409f
C1079 VP.t1 VSUBS 2.76252f
C1080 VP.n1 VSUBS 0.03791f
C1081 VP.n2 VSUBS 0.03065f
C1082 VP.t4 VSUBS 2.76252f
C1083 VP.n3 VSUBS 0.971851f
C1084 VP.n4 VSUBS 0.03065f
C1085 VP.n5 VSUBS 0.061064f
C1086 VP.n6 VSUBS 0.03065f
C1087 VP.t9 VSUBS 2.76252f
C1088 VP.n7 VSUBS 0.029897f
C1089 VP.n8 VSUBS 0.03065f
C1090 VP.t2 VSUBS 2.76252f
C1091 VP.n9 VSUBS 0.057124f
C1092 VP.n10 VSUBS 0.03065f
C1093 VP.n11 VSUBS 0.039638f
C1094 VP.n12 VSUBS 0.040409f
C1095 VP.t7 VSUBS 2.76252f
C1096 VP.n13 VSUBS 0.03791f
C1097 VP.n14 VSUBS 0.03065f
C1098 VP.t5 VSUBS 2.76252f
C1099 VP.n15 VSUBS 0.971851f
C1100 VP.n16 VSUBS 0.03065f
C1101 VP.n17 VSUBS 0.061064f
C1102 VP.n18 VSUBS 0.03065f
C1103 VP.t6 VSUBS 2.76252f
C1104 VP.n19 VSUBS 0.029897f
C1105 VP.n20 VSUBS 0.289729f
C1106 VP.t3 VSUBS 2.76252f
C1107 VP.t0 VSUBS 2.98536f
C1108 VP.n21 VSUBS 1.0345f
C1109 VP.n22 VSUBS 1.07032f
C1110 VP.n23 VSUBS 0.055432f
C1111 VP.n24 VSUBS 0.055649f
C1112 VP.n25 VSUBS 0.03065f
C1113 VP.n26 VSUBS 0.03065f
C1114 VP.n27 VSUBS 0.03065f
C1115 VP.n28 VSUBS 0.061064f
C1116 VP.n29 VSUBS 0.043022f
C1117 VP.n30 VSUBS 0.971851f
C1118 VP.n31 VSUBS 0.043022f
C1119 VP.n32 VSUBS 0.03065f
C1120 VP.n33 VSUBS 0.03065f
C1121 VP.n34 VSUBS 0.03065f
C1122 VP.n35 VSUBS 0.029897f
C1123 VP.n36 VSUBS 0.055649f
C1124 VP.n37 VSUBS 0.055432f
C1125 VP.n38 VSUBS 0.03065f
C1126 VP.n39 VSUBS 0.03065f
C1127 VP.n40 VSUBS 0.030614f
C1128 VP.n41 VSUBS 0.057124f
C1129 VP.n42 VSUBS 0.051576f
C1130 VP.n43 VSUBS 0.03065f
C1131 VP.n44 VSUBS 0.03065f
C1132 VP.n45 VSUBS 0.03065f
C1133 VP.n46 VSUBS 0.057124f
C1134 VP.n47 VSUBS 0.039638f
C1135 VP.n48 VSUBS 1.06475f
C1136 VP.n49 VSUBS 1.86761f
C1137 VP.t8 VSUBS 2.76252f
C1138 VP.n50 VSUBS 1.06475f
C1139 VP.n51 VSUBS 1.88829f
C1140 VP.n52 VSUBS 0.040409f
C1141 VP.n53 VSUBS 0.03065f
C1142 VP.n54 VSUBS 0.057124f
C1143 VP.n55 VSUBS 0.03791f
C1144 VP.n56 VSUBS 0.051576f
C1145 VP.n57 VSUBS 0.03065f
C1146 VP.n58 VSUBS 0.03065f
C1147 VP.n59 VSUBS 0.03065f
C1148 VP.n60 VSUBS 0.030614f
C1149 VP.n61 VSUBS 0.971851f
C1150 VP.n62 VSUBS 0.055432f
C1151 VP.n63 VSUBS 0.055649f
C1152 VP.n64 VSUBS 0.03065f
C1153 VP.n65 VSUBS 0.03065f
C1154 VP.n66 VSUBS 0.03065f
C1155 VP.n67 VSUBS 0.061064f
C1156 VP.n68 VSUBS 0.043022f
C1157 VP.n69 VSUBS 0.971851f
C1158 VP.n70 VSUBS 0.043022f
C1159 VP.n71 VSUBS 0.03065f
C1160 VP.n72 VSUBS 0.03065f
C1161 VP.n73 VSUBS 0.03065f
C1162 VP.n74 VSUBS 0.029897f
C1163 VP.n75 VSUBS 0.055649f
C1164 VP.n76 VSUBS 0.055432f
C1165 VP.n77 VSUBS 0.03065f
C1166 VP.n78 VSUBS 0.03065f
C1167 VP.n79 VSUBS 0.030614f
C1168 VP.n80 VSUBS 0.057124f
C1169 VP.n81 VSUBS 0.051576f
C1170 VP.n82 VSUBS 0.03065f
C1171 VP.n83 VSUBS 0.03065f
C1172 VP.n84 VSUBS 0.03065f
C1173 VP.n85 VSUBS 0.057124f
C1174 VP.n86 VSUBS 0.039638f
C1175 VP.n87 VSUBS 1.06475f
C1176 VP.n88 VSUBS 0.048349f
.ends

