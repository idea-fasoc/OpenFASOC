* NGSPICE file created from diff_pair_sample_0618.ext - technology: sky130A

.subckt diff_pair_sample_0618 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.49325 pd=9.38 as=3.5295 ps=18.88 w=9.05 l=2.58
X1 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=3.5295 pd=18.88 as=0 ps=0 w=9.05 l=2.58
X2 VDD2.t3 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.49325 pd=9.38 as=3.5295 ps=18.88 w=9.05 l=2.58
X3 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=3.5295 pd=18.88 as=0 ps=0 w=9.05 l=2.58
X4 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.5295 pd=18.88 as=0 ps=0 w=9.05 l=2.58
X5 VTAIL.t2 VP.t1 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=3.5295 pd=18.88 as=1.49325 ps=9.38 w=9.05 l=2.58
X6 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.5295 pd=18.88 as=0 ps=0 w=9.05 l=2.58
X7 VDD2.t2 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.49325 pd=9.38 as=3.5295 ps=18.88 w=9.05 l=2.58
X8 VTAIL.t7 VN.t2 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=3.5295 pd=18.88 as=1.49325 ps=9.38 w=9.05 l=2.58
X9 VDD1.t1 VP.t2 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.49325 pd=9.38 as=3.5295 ps=18.88 w=9.05 l=2.58
X10 VTAIL.t5 VP.t3 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=3.5295 pd=18.88 as=1.49325 ps=9.38 w=9.05 l=2.58
X11 VTAIL.t6 VN.t3 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=3.5295 pd=18.88 as=1.49325 ps=9.38 w=9.05 l=2.58
R0 VP.n14 VP.n0 161.3
R1 VP.n13 VP.n12 161.3
R2 VP.n11 VP.n1 161.3
R3 VP.n10 VP.n9 161.3
R4 VP.n8 VP.n2 161.3
R5 VP.n7 VP.n6 161.3
R6 VP.n4 VP.t3 120.582
R7 VP.n4 VP.t2 119.811
R8 VP.n5 VP.n3 100.725
R9 VP.n16 VP.n15 100.725
R10 VP.n3 VP.t1 84.5373
R11 VP.n15 VP.t0 84.5373
R12 VP.n9 VP.n1 56.5193
R13 VP.n5 VP.n4 48.391
R14 VP.n8 VP.n7 24.4675
R15 VP.n9 VP.n8 24.4675
R16 VP.n13 VP.n1 24.4675
R17 VP.n14 VP.n13 24.4675
R18 VP.n7 VP.n3 10.032
R19 VP.n15 VP.n14 10.032
R20 VP.n6 VP.n5 0.278367
R21 VP.n16 VP.n0 0.278367
R22 VP.n6 VP.n2 0.189894
R23 VP.n10 VP.n2 0.189894
R24 VP.n11 VP.n10 0.189894
R25 VP.n12 VP.n11 0.189894
R26 VP.n12 VP.n0 0.189894
R27 VP VP.n16 0.153454
R28 VTAIL.n5 VTAIL.t5 52.0163
R29 VTAIL.n4 VTAIL.t1 52.0163
R30 VTAIL.n3 VTAIL.t7 52.0163
R31 VTAIL.n7 VTAIL.t0 52.0161
R32 VTAIL.n0 VTAIL.t6 52.0161
R33 VTAIL.n1 VTAIL.t3 52.0161
R34 VTAIL.n2 VTAIL.t2 52.0161
R35 VTAIL.n6 VTAIL.t4 52.0161
R36 VTAIL.n7 VTAIL.n6 22.6772
R37 VTAIL.n3 VTAIL.n2 22.6772
R38 VTAIL.n4 VTAIL.n3 2.50912
R39 VTAIL.n6 VTAIL.n5 2.50912
R40 VTAIL.n2 VTAIL.n1 2.50912
R41 VTAIL VTAIL.n0 1.313
R42 VTAIL VTAIL.n7 1.19662
R43 VTAIL.n5 VTAIL.n4 0.470328
R44 VTAIL.n1 VTAIL.n0 0.470328
R45 VDD1 VDD1.n1 106.075
R46 VDD1 VDD1.n0 66.5653
R47 VDD1.n0 VDD1.t0 2.18835
R48 VDD1.n0 VDD1.t1 2.18835
R49 VDD1.n1 VDD1.t2 2.18835
R50 VDD1.n1 VDD1.t3 2.18835
R51 B.n512 B.n107 585
R52 B.n107 B.n64 585
R53 B.n514 B.n513 585
R54 B.n516 B.n106 585
R55 B.n519 B.n518 585
R56 B.n520 B.n105 585
R57 B.n522 B.n521 585
R58 B.n524 B.n104 585
R59 B.n527 B.n526 585
R60 B.n528 B.n103 585
R61 B.n530 B.n529 585
R62 B.n532 B.n102 585
R63 B.n535 B.n534 585
R64 B.n536 B.n101 585
R65 B.n538 B.n537 585
R66 B.n540 B.n100 585
R67 B.n543 B.n542 585
R68 B.n544 B.n99 585
R69 B.n546 B.n545 585
R70 B.n548 B.n98 585
R71 B.n551 B.n550 585
R72 B.n552 B.n97 585
R73 B.n554 B.n553 585
R74 B.n556 B.n96 585
R75 B.n559 B.n558 585
R76 B.n560 B.n95 585
R77 B.n562 B.n561 585
R78 B.n564 B.n94 585
R79 B.n567 B.n566 585
R80 B.n568 B.n93 585
R81 B.n570 B.n569 585
R82 B.n572 B.n92 585
R83 B.n574 B.n573 585
R84 B.n576 B.n575 585
R85 B.n579 B.n578 585
R86 B.n580 B.n87 585
R87 B.n582 B.n581 585
R88 B.n584 B.n86 585
R89 B.n587 B.n586 585
R90 B.n588 B.n85 585
R91 B.n590 B.n589 585
R92 B.n592 B.n84 585
R93 B.n595 B.n594 585
R94 B.n597 B.n81 585
R95 B.n599 B.n598 585
R96 B.n601 B.n80 585
R97 B.n604 B.n603 585
R98 B.n605 B.n79 585
R99 B.n607 B.n606 585
R100 B.n609 B.n78 585
R101 B.n612 B.n611 585
R102 B.n613 B.n77 585
R103 B.n615 B.n614 585
R104 B.n617 B.n76 585
R105 B.n620 B.n619 585
R106 B.n621 B.n75 585
R107 B.n623 B.n622 585
R108 B.n625 B.n74 585
R109 B.n628 B.n627 585
R110 B.n629 B.n73 585
R111 B.n631 B.n630 585
R112 B.n633 B.n72 585
R113 B.n636 B.n635 585
R114 B.n637 B.n71 585
R115 B.n639 B.n638 585
R116 B.n641 B.n70 585
R117 B.n644 B.n643 585
R118 B.n645 B.n69 585
R119 B.n647 B.n646 585
R120 B.n649 B.n68 585
R121 B.n652 B.n651 585
R122 B.n653 B.n67 585
R123 B.n655 B.n654 585
R124 B.n657 B.n66 585
R125 B.n660 B.n659 585
R126 B.n661 B.n65 585
R127 B.n511 B.n63 585
R128 B.n664 B.n63 585
R129 B.n510 B.n62 585
R130 B.n665 B.n62 585
R131 B.n509 B.n61 585
R132 B.n666 B.n61 585
R133 B.n508 B.n507 585
R134 B.n507 B.n57 585
R135 B.n506 B.n56 585
R136 B.n672 B.n56 585
R137 B.n505 B.n55 585
R138 B.n673 B.n55 585
R139 B.n504 B.n54 585
R140 B.n674 B.n54 585
R141 B.n503 B.n502 585
R142 B.n502 B.n53 585
R143 B.n501 B.n49 585
R144 B.n680 B.n49 585
R145 B.n500 B.n48 585
R146 B.n681 B.n48 585
R147 B.n499 B.n47 585
R148 B.n682 B.n47 585
R149 B.n498 B.n497 585
R150 B.n497 B.n43 585
R151 B.n496 B.n42 585
R152 B.n688 B.n42 585
R153 B.n495 B.n41 585
R154 B.n689 B.n41 585
R155 B.n494 B.n40 585
R156 B.n690 B.n40 585
R157 B.n493 B.n492 585
R158 B.n492 B.n36 585
R159 B.n491 B.n35 585
R160 B.n696 B.n35 585
R161 B.n490 B.n34 585
R162 B.n697 B.n34 585
R163 B.n489 B.n33 585
R164 B.n698 B.n33 585
R165 B.n488 B.n487 585
R166 B.n487 B.n32 585
R167 B.n486 B.n28 585
R168 B.n704 B.n28 585
R169 B.n485 B.n27 585
R170 B.n705 B.n27 585
R171 B.n484 B.n26 585
R172 B.n706 B.n26 585
R173 B.n483 B.n482 585
R174 B.n482 B.n22 585
R175 B.n481 B.n21 585
R176 B.n712 B.n21 585
R177 B.n480 B.n20 585
R178 B.n713 B.n20 585
R179 B.n479 B.n19 585
R180 B.n714 B.n19 585
R181 B.n478 B.n477 585
R182 B.n477 B.n15 585
R183 B.n476 B.n14 585
R184 B.n720 B.n14 585
R185 B.n475 B.n13 585
R186 B.n721 B.n13 585
R187 B.n474 B.n12 585
R188 B.n722 B.n12 585
R189 B.n473 B.n472 585
R190 B.n472 B.n8 585
R191 B.n471 B.n7 585
R192 B.n728 B.n7 585
R193 B.n470 B.n6 585
R194 B.n729 B.n6 585
R195 B.n469 B.n5 585
R196 B.n730 B.n5 585
R197 B.n468 B.n467 585
R198 B.n467 B.n4 585
R199 B.n466 B.n108 585
R200 B.n466 B.n465 585
R201 B.n456 B.n109 585
R202 B.n110 B.n109 585
R203 B.n458 B.n457 585
R204 B.n459 B.n458 585
R205 B.n455 B.n115 585
R206 B.n115 B.n114 585
R207 B.n454 B.n453 585
R208 B.n453 B.n452 585
R209 B.n117 B.n116 585
R210 B.n118 B.n117 585
R211 B.n445 B.n444 585
R212 B.n446 B.n445 585
R213 B.n443 B.n123 585
R214 B.n123 B.n122 585
R215 B.n442 B.n441 585
R216 B.n441 B.n440 585
R217 B.n125 B.n124 585
R218 B.n126 B.n125 585
R219 B.n433 B.n432 585
R220 B.n434 B.n433 585
R221 B.n431 B.n131 585
R222 B.n131 B.n130 585
R223 B.n430 B.n429 585
R224 B.n429 B.n428 585
R225 B.n133 B.n132 585
R226 B.n421 B.n133 585
R227 B.n420 B.n419 585
R228 B.n422 B.n420 585
R229 B.n418 B.n138 585
R230 B.n138 B.n137 585
R231 B.n417 B.n416 585
R232 B.n416 B.n415 585
R233 B.n140 B.n139 585
R234 B.n141 B.n140 585
R235 B.n408 B.n407 585
R236 B.n409 B.n408 585
R237 B.n406 B.n146 585
R238 B.n146 B.n145 585
R239 B.n405 B.n404 585
R240 B.n404 B.n403 585
R241 B.n148 B.n147 585
R242 B.n149 B.n148 585
R243 B.n396 B.n395 585
R244 B.n397 B.n396 585
R245 B.n394 B.n154 585
R246 B.n154 B.n153 585
R247 B.n393 B.n392 585
R248 B.n392 B.n391 585
R249 B.n156 B.n155 585
R250 B.n384 B.n156 585
R251 B.n383 B.n382 585
R252 B.n385 B.n383 585
R253 B.n381 B.n161 585
R254 B.n161 B.n160 585
R255 B.n380 B.n379 585
R256 B.n379 B.n378 585
R257 B.n163 B.n162 585
R258 B.n164 B.n163 585
R259 B.n371 B.n370 585
R260 B.n372 B.n371 585
R261 B.n369 B.n169 585
R262 B.n169 B.n168 585
R263 B.n368 B.n367 585
R264 B.n367 B.n366 585
R265 B.n363 B.n173 585
R266 B.n362 B.n361 585
R267 B.n359 B.n174 585
R268 B.n359 B.n172 585
R269 B.n358 B.n357 585
R270 B.n356 B.n355 585
R271 B.n354 B.n176 585
R272 B.n352 B.n351 585
R273 B.n350 B.n177 585
R274 B.n349 B.n348 585
R275 B.n346 B.n178 585
R276 B.n344 B.n343 585
R277 B.n342 B.n179 585
R278 B.n341 B.n340 585
R279 B.n338 B.n180 585
R280 B.n336 B.n335 585
R281 B.n334 B.n181 585
R282 B.n333 B.n332 585
R283 B.n330 B.n182 585
R284 B.n328 B.n327 585
R285 B.n326 B.n183 585
R286 B.n325 B.n324 585
R287 B.n322 B.n184 585
R288 B.n320 B.n319 585
R289 B.n318 B.n185 585
R290 B.n317 B.n316 585
R291 B.n314 B.n186 585
R292 B.n312 B.n311 585
R293 B.n310 B.n187 585
R294 B.n309 B.n308 585
R295 B.n306 B.n188 585
R296 B.n304 B.n303 585
R297 B.n302 B.n189 585
R298 B.n301 B.n300 585
R299 B.n298 B.n297 585
R300 B.n296 B.n295 585
R301 B.n294 B.n194 585
R302 B.n292 B.n291 585
R303 B.n290 B.n195 585
R304 B.n289 B.n288 585
R305 B.n286 B.n196 585
R306 B.n284 B.n283 585
R307 B.n282 B.n197 585
R308 B.n280 B.n279 585
R309 B.n277 B.n200 585
R310 B.n275 B.n274 585
R311 B.n273 B.n201 585
R312 B.n272 B.n271 585
R313 B.n269 B.n202 585
R314 B.n267 B.n266 585
R315 B.n265 B.n203 585
R316 B.n264 B.n263 585
R317 B.n261 B.n204 585
R318 B.n259 B.n258 585
R319 B.n257 B.n205 585
R320 B.n256 B.n255 585
R321 B.n253 B.n206 585
R322 B.n251 B.n250 585
R323 B.n249 B.n207 585
R324 B.n248 B.n247 585
R325 B.n245 B.n208 585
R326 B.n243 B.n242 585
R327 B.n241 B.n209 585
R328 B.n240 B.n239 585
R329 B.n237 B.n210 585
R330 B.n235 B.n234 585
R331 B.n233 B.n211 585
R332 B.n232 B.n231 585
R333 B.n229 B.n212 585
R334 B.n227 B.n226 585
R335 B.n225 B.n213 585
R336 B.n224 B.n223 585
R337 B.n221 B.n214 585
R338 B.n219 B.n218 585
R339 B.n217 B.n216 585
R340 B.n171 B.n170 585
R341 B.n365 B.n364 585
R342 B.n366 B.n365 585
R343 B.n167 B.n166 585
R344 B.n168 B.n167 585
R345 B.n374 B.n373 585
R346 B.n373 B.n372 585
R347 B.n375 B.n165 585
R348 B.n165 B.n164 585
R349 B.n377 B.n376 585
R350 B.n378 B.n377 585
R351 B.n159 B.n158 585
R352 B.n160 B.n159 585
R353 B.n387 B.n386 585
R354 B.n386 B.n385 585
R355 B.n388 B.n157 585
R356 B.n384 B.n157 585
R357 B.n390 B.n389 585
R358 B.n391 B.n390 585
R359 B.n152 B.n151 585
R360 B.n153 B.n152 585
R361 B.n399 B.n398 585
R362 B.n398 B.n397 585
R363 B.n400 B.n150 585
R364 B.n150 B.n149 585
R365 B.n402 B.n401 585
R366 B.n403 B.n402 585
R367 B.n144 B.n143 585
R368 B.n145 B.n144 585
R369 B.n411 B.n410 585
R370 B.n410 B.n409 585
R371 B.n412 B.n142 585
R372 B.n142 B.n141 585
R373 B.n414 B.n413 585
R374 B.n415 B.n414 585
R375 B.n136 B.n135 585
R376 B.n137 B.n136 585
R377 B.n424 B.n423 585
R378 B.n423 B.n422 585
R379 B.n425 B.n134 585
R380 B.n421 B.n134 585
R381 B.n427 B.n426 585
R382 B.n428 B.n427 585
R383 B.n129 B.n128 585
R384 B.n130 B.n129 585
R385 B.n436 B.n435 585
R386 B.n435 B.n434 585
R387 B.n437 B.n127 585
R388 B.n127 B.n126 585
R389 B.n439 B.n438 585
R390 B.n440 B.n439 585
R391 B.n121 B.n120 585
R392 B.n122 B.n121 585
R393 B.n448 B.n447 585
R394 B.n447 B.n446 585
R395 B.n449 B.n119 585
R396 B.n119 B.n118 585
R397 B.n451 B.n450 585
R398 B.n452 B.n451 585
R399 B.n113 B.n112 585
R400 B.n114 B.n113 585
R401 B.n461 B.n460 585
R402 B.n460 B.n459 585
R403 B.n462 B.n111 585
R404 B.n111 B.n110 585
R405 B.n464 B.n463 585
R406 B.n465 B.n464 585
R407 B.n2 B.n0 585
R408 B.n4 B.n2 585
R409 B.n3 B.n1 585
R410 B.n729 B.n3 585
R411 B.n727 B.n726 585
R412 B.n728 B.n727 585
R413 B.n725 B.n9 585
R414 B.n9 B.n8 585
R415 B.n724 B.n723 585
R416 B.n723 B.n722 585
R417 B.n11 B.n10 585
R418 B.n721 B.n11 585
R419 B.n719 B.n718 585
R420 B.n720 B.n719 585
R421 B.n717 B.n16 585
R422 B.n16 B.n15 585
R423 B.n716 B.n715 585
R424 B.n715 B.n714 585
R425 B.n18 B.n17 585
R426 B.n713 B.n18 585
R427 B.n711 B.n710 585
R428 B.n712 B.n711 585
R429 B.n709 B.n23 585
R430 B.n23 B.n22 585
R431 B.n708 B.n707 585
R432 B.n707 B.n706 585
R433 B.n25 B.n24 585
R434 B.n705 B.n25 585
R435 B.n703 B.n702 585
R436 B.n704 B.n703 585
R437 B.n701 B.n29 585
R438 B.n32 B.n29 585
R439 B.n700 B.n699 585
R440 B.n699 B.n698 585
R441 B.n31 B.n30 585
R442 B.n697 B.n31 585
R443 B.n695 B.n694 585
R444 B.n696 B.n695 585
R445 B.n693 B.n37 585
R446 B.n37 B.n36 585
R447 B.n692 B.n691 585
R448 B.n691 B.n690 585
R449 B.n39 B.n38 585
R450 B.n689 B.n39 585
R451 B.n687 B.n686 585
R452 B.n688 B.n687 585
R453 B.n685 B.n44 585
R454 B.n44 B.n43 585
R455 B.n684 B.n683 585
R456 B.n683 B.n682 585
R457 B.n46 B.n45 585
R458 B.n681 B.n46 585
R459 B.n679 B.n678 585
R460 B.n680 B.n679 585
R461 B.n677 B.n50 585
R462 B.n53 B.n50 585
R463 B.n676 B.n675 585
R464 B.n675 B.n674 585
R465 B.n52 B.n51 585
R466 B.n673 B.n52 585
R467 B.n671 B.n670 585
R468 B.n672 B.n671 585
R469 B.n669 B.n58 585
R470 B.n58 B.n57 585
R471 B.n668 B.n667 585
R472 B.n667 B.n666 585
R473 B.n60 B.n59 585
R474 B.n665 B.n60 585
R475 B.n663 B.n662 585
R476 B.n664 B.n663 585
R477 B.n732 B.n731 585
R478 B.n731 B.n730 585
R479 B.n365 B.n173 502.111
R480 B.n663 B.n65 502.111
R481 B.n367 B.n171 502.111
R482 B.n107 B.n63 502.111
R483 B.n198 B.t4 292.553
R484 B.n190 B.t12 292.553
R485 B.n82 B.t15 292.553
R486 B.n88 B.t8 292.553
R487 B.n515 B.n64 256.663
R488 B.n517 B.n64 256.663
R489 B.n523 B.n64 256.663
R490 B.n525 B.n64 256.663
R491 B.n531 B.n64 256.663
R492 B.n533 B.n64 256.663
R493 B.n539 B.n64 256.663
R494 B.n541 B.n64 256.663
R495 B.n547 B.n64 256.663
R496 B.n549 B.n64 256.663
R497 B.n555 B.n64 256.663
R498 B.n557 B.n64 256.663
R499 B.n563 B.n64 256.663
R500 B.n565 B.n64 256.663
R501 B.n571 B.n64 256.663
R502 B.n91 B.n64 256.663
R503 B.n577 B.n64 256.663
R504 B.n583 B.n64 256.663
R505 B.n585 B.n64 256.663
R506 B.n591 B.n64 256.663
R507 B.n593 B.n64 256.663
R508 B.n600 B.n64 256.663
R509 B.n602 B.n64 256.663
R510 B.n608 B.n64 256.663
R511 B.n610 B.n64 256.663
R512 B.n616 B.n64 256.663
R513 B.n618 B.n64 256.663
R514 B.n624 B.n64 256.663
R515 B.n626 B.n64 256.663
R516 B.n632 B.n64 256.663
R517 B.n634 B.n64 256.663
R518 B.n640 B.n64 256.663
R519 B.n642 B.n64 256.663
R520 B.n648 B.n64 256.663
R521 B.n650 B.n64 256.663
R522 B.n656 B.n64 256.663
R523 B.n658 B.n64 256.663
R524 B.n360 B.n172 256.663
R525 B.n175 B.n172 256.663
R526 B.n353 B.n172 256.663
R527 B.n347 B.n172 256.663
R528 B.n345 B.n172 256.663
R529 B.n339 B.n172 256.663
R530 B.n337 B.n172 256.663
R531 B.n331 B.n172 256.663
R532 B.n329 B.n172 256.663
R533 B.n323 B.n172 256.663
R534 B.n321 B.n172 256.663
R535 B.n315 B.n172 256.663
R536 B.n313 B.n172 256.663
R537 B.n307 B.n172 256.663
R538 B.n305 B.n172 256.663
R539 B.n299 B.n172 256.663
R540 B.n193 B.n172 256.663
R541 B.n293 B.n172 256.663
R542 B.n287 B.n172 256.663
R543 B.n285 B.n172 256.663
R544 B.n278 B.n172 256.663
R545 B.n276 B.n172 256.663
R546 B.n270 B.n172 256.663
R547 B.n268 B.n172 256.663
R548 B.n262 B.n172 256.663
R549 B.n260 B.n172 256.663
R550 B.n254 B.n172 256.663
R551 B.n252 B.n172 256.663
R552 B.n246 B.n172 256.663
R553 B.n244 B.n172 256.663
R554 B.n238 B.n172 256.663
R555 B.n236 B.n172 256.663
R556 B.n230 B.n172 256.663
R557 B.n228 B.n172 256.663
R558 B.n222 B.n172 256.663
R559 B.n220 B.n172 256.663
R560 B.n215 B.n172 256.663
R561 B.n365 B.n167 163.367
R562 B.n373 B.n167 163.367
R563 B.n373 B.n165 163.367
R564 B.n377 B.n165 163.367
R565 B.n377 B.n159 163.367
R566 B.n386 B.n159 163.367
R567 B.n386 B.n157 163.367
R568 B.n390 B.n157 163.367
R569 B.n390 B.n152 163.367
R570 B.n398 B.n152 163.367
R571 B.n398 B.n150 163.367
R572 B.n402 B.n150 163.367
R573 B.n402 B.n144 163.367
R574 B.n410 B.n144 163.367
R575 B.n410 B.n142 163.367
R576 B.n414 B.n142 163.367
R577 B.n414 B.n136 163.367
R578 B.n423 B.n136 163.367
R579 B.n423 B.n134 163.367
R580 B.n427 B.n134 163.367
R581 B.n427 B.n129 163.367
R582 B.n435 B.n129 163.367
R583 B.n435 B.n127 163.367
R584 B.n439 B.n127 163.367
R585 B.n439 B.n121 163.367
R586 B.n447 B.n121 163.367
R587 B.n447 B.n119 163.367
R588 B.n451 B.n119 163.367
R589 B.n451 B.n113 163.367
R590 B.n460 B.n113 163.367
R591 B.n460 B.n111 163.367
R592 B.n464 B.n111 163.367
R593 B.n464 B.n2 163.367
R594 B.n731 B.n2 163.367
R595 B.n731 B.n3 163.367
R596 B.n727 B.n3 163.367
R597 B.n727 B.n9 163.367
R598 B.n723 B.n9 163.367
R599 B.n723 B.n11 163.367
R600 B.n719 B.n11 163.367
R601 B.n719 B.n16 163.367
R602 B.n715 B.n16 163.367
R603 B.n715 B.n18 163.367
R604 B.n711 B.n18 163.367
R605 B.n711 B.n23 163.367
R606 B.n707 B.n23 163.367
R607 B.n707 B.n25 163.367
R608 B.n703 B.n25 163.367
R609 B.n703 B.n29 163.367
R610 B.n699 B.n29 163.367
R611 B.n699 B.n31 163.367
R612 B.n695 B.n31 163.367
R613 B.n695 B.n37 163.367
R614 B.n691 B.n37 163.367
R615 B.n691 B.n39 163.367
R616 B.n687 B.n39 163.367
R617 B.n687 B.n44 163.367
R618 B.n683 B.n44 163.367
R619 B.n683 B.n46 163.367
R620 B.n679 B.n46 163.367
R621 B.n679 B.n50 163.367
R622 B.n675 B.n50 163.367
R623 B.n675 B.n52 163.367
R624 B.n671 B.n52 163.367
R625 B.n671 B.n58 163.367
R626 B.n667 B.n58 163.367
R627 B.n667 B.n60 163.367
R628 B.n663 B.n60 163.367
R629 B.n361 B.n359 163.367
R630 B.n359 B.n358 163.367
R631 B.n355 B.n354 163.367
R632 B.n352 B.n177 163.367
R633 B.n348 B.n346 163.367
R634 B.n344 B.n179 163.367
R635 B.n340 B.n338 163.367
R636 B.n336 B.n181 163.367
R637 B.n332 B.n330 163.367
R638 B.n328 B.n183 163.367
R639 B.n324 B.n322 163.367
R640 B.n320 B.n185 163.367
R641 B.n316 B.n314 163.367
R642 B.n312 B.n187 163.367
R643 B.n308 B.n306 163.367
R644 B.n304 B.n189 163.367
R645 B.n300 B.n298 163.367
R646 B.n295 B.n294 163.367
R647 B.n292 B.n195 163.367
R648 B.n288 B.n286 163.367
R649 B.n284 B.n197 163.367
R650 B.n279 B.n277 163.367
R651 B.n275 B.n201 163.367
R652 B.n271 B.n269 163.367
R653 B.n267 B.n203 163.367
R654 B.n263 B.n261 163.367
R655 B.n259 B.n205 163.367
R656 B.n255 B.n253 163.367
R657 B.n251 B.n207 163.367
R658 B.n247 B.n245 163.367
R659 B.n243 B.n209 163.367
R660 B.n239 B.n237 163.367
R661 B.n235 B.n211 163.367
R662 B.n231 B.n229 163.367
R663 B.n227 B.n213 163.367
R664 B.n223 B.n221 163.367
R665 B.n219 B.n216 163.367
R666 B.n367 B.n169 163.367
R667 B.n371 B.n169 163.367
R668 B.n371 B.n163 163.367
R669 B.n379 B.n163 163.367
R670 B.n379 B.n161 163.367
R671 B.n383 B.n161 163.367
R672 B.n383 B.n156 163.367
R673 B.n392 B.n156 163.367
R674 B.n392 B.n154 163.367
R675 B.n396 B.n154 163.367
R676 B.n396 B.n148 163.367
R677 B.n404 B.n148 163.367
R678 B.n404 B.n146 163.367
R679 B.n408 B.n146 163.367
R680 B.n408 B.n140 163.367
R681 B.n416 B.n140 163.367
R682 B.n416 B.n138 163.367
R683 B.n420 B.n138 163.367
R684 B.n420 B.n133 163.367
R685 B.n429 B.n133 163.367
R686 B.n429 B.n131 163.367
R687 B.n433 B.n131 163.367
R688 B.n433 B.n125 163.367
R689 B.n441 B.n125 163.367
R690 B.n441 B.n123 163.367
R691 B.n445 B.n123 163.367
R692 B.n445 B.n117 163.367
R693 B.n453 B.n117 163.367
R694 B.n453 B.n115 163.367
R695 B.n458 B.n115 163.367
R696 B.n458 B.n109 163.367
R697 B.n466 B.n109 163.367
R698 B.n467 B.n466 163.367
R699 B.n467 B.n5 163.367
R700 B.n6 B.n5 163.367
R701 B.n7 B.n6 163.367
R702 B.n472 B.n7 163.367
R703 B.n472 B.n12 163.367
R704 B.n13 B.n12 163.367
R705 B.n14 B.n13 163.367
R706 B.n477 B.n14 163.367
R707 B.n477 B.n19 163.367
R708 B.n20 B.n19 163.367
R709 B.n21 B.n20 163.367
R710 B.n482 B.n21 163.367
R711 B.n482 B.n26 163.367
R712 B.n27 B.n26 163.367
R713 B.n28 B.n27 163.367
R714 B.n487 B.n28 163.367
R715 B.n487 B.n33 163.367
R716 B.n34 B.n33 163.367
R717 B.n35 B.n34 163.367
R718 B.n492 B.n35 163.367
R719 B.n492 B.n40 163.367
R720 B.n41 B.n40 163.367
R721 B.n42 B.n41 163.367
R722 B.n497 B.n42 163.367
R723 B.n497 B.n47 163.367
R724 B.n48 B.n47 163.367
R725 B.n49 B.n48 163.367
R726 B.n502 B.n49 163.367
R727 B.n502 B.n54 163.367
R728 B.n55 B.n54 163.367
R729 B.n56 B.n55 163.367
R730 B.n507 B.n56 163.367
R731 B.n507 B.n61 163.367
R732 B.n62 B.n61 163.367
R733 B.n63 B.n62 163.367
R734 B.n659 B.n657 163.367
R735 B.n655 B.n67 163.367
R736 B.n651 B.n649 163.367
R737 B.n647 B.n69 163.367
R738 B.n643 B.n641 163.367
R739 B.n639 B.n71 163.367
R740 B.n635 B.n633 163.367
R741 B.n631 B.n73 163.367
R742 B.n627 B.n625 163.367
R743 B.n623 B.n75 163.367
R744 B.n619 B.n617 163.367
R745 B.n615 B.n77 163.367
R746 B.n611 B.n609 163.367
R747 B.n607 B.n79 163.367
R748 B.n603 B.n601 163.367
R749 B.n599 B.n81 163.367
R750 B.n594 B.n592 163.367
R751 B.n590 B.n85 163.367
R752 B.n586 B.n584 163.367
R753 B.n582 B.n87 163.367
R754 B.n578 B.n576 163.367
R755 B.n573 B.n572 163.367
R756 B.n570 B.n93 163.367
R757 B.n566 B.n564 163.367
R758 B.n562 B.n95 163.367
R759 B.n558 B.n556 163.367
R760 B.n554 B.n97 163.367
R761 B.n550 B.n548 163.367
R762 B.n546 B.n99 163.367
R763 B.n542 B.n540 163.367
R764 B.n538 B.n101 163.367
R765 B.n534 B.n532 163.367
R766 B.n530 B.n103 163.367
R767 B.n526 B.n524 163.367
R768 B.n522 B.n105 163.367
R769 B.n518 B.n516 163.367
R770 B.n514 B.n107 163.367
R771 B.n198 B.t7 128.833
R772 B.n88 B.t10 128.833
R773 B.n190 B.t14 128.821
R774 B.n82 B.t16 128.821
R775 B.n366 B.n172 83.7003
R776 B.n664 B.n64 83.7003
R777 B.n199 B.t6 72.3961
R778 B.n89 B.t11 72.3961
R779 B.n191 B.t13 72.3854
R780 B.n83 B.t17 72.3854
R781 B.n360 B.n173 71.676
R782 B.n358 B.n175 71.676
R783 B.n354 B.n353 71.676
R784 B.n347 B.n177 71.676
R785 B.n346 B.n345 71.676
R786 B.n339 B.n179 71.676
R787 B.n338 B.n337 71.676
R788 B.n331 B.n181 71.676
R789 B.n330 B.n329 71.676
R790 B.n323 B.n183 71.676
R791 B.n322 B.n321 71.676
R792 B.n315 B.n185 71.676
R793 B.n314 B.n313 71.676
R794 B.n307 B.n187 71.676
R795 B.n306 B.n305 71.676
R796 B.n299 B.n189 71.676
R797 B.n298 B.n193 71.676
R798 B.n294 B.n293 71.676
R799 B.n287 B.n195 71.676
R800 B.n286 B.n285 71.676
R801 B.n278 B.n197 71.676
R802 B.n277 B.n276 71.676
R803 B.n270 B.n201 71.676
R804 B.n269 B.n268 71.676
R805 B.n262 B.n203 71.676
R806 B.n261 B.n260 71.676
R807 B.n254 B.n205 71.676
R808 B.n253 B.n252 71.676
R809 B.n246 B.n207 71.676
R810 B.n245 B.n244 71.676
R811 B.n238 B.n209 71.676
R812 B.n237 B.n236 71.676
R813 B.n230 B.n211 71.676
R814 B.n229 B.n228 71.676
R815 B.n222 B.n213 71.676
R816 B.n221 B.n220 71.676
R817 B.n216 B.n215 71.676
R818 B.n658 B.n65 71.676
R819 B.n657 B.n656 71.676
R820 B.n650 B.n67 71.676
R821 B.n649 B.n648 71.676
R822 B.n642 B.n69 71.676
R823 B.n641 B.n640 71.676
R824 B.n634 B.n71 71.676
R825 B.n633 B.n632 71.676
R826 B.n626 B.n73 71.676
R827 B.n625 B.n624 71.676
R828 B.n618 B.n75 71.676
R829 B.n617 B.n616 71.676
R830 B.n610 B.n77 71.676
R831 B.n609 B.n608 71.676
R832 B.n602 B.n79 71.676
R833 B.n601 B.n600 71.676
R834 B.n593 B.n81 71.676
R835 B.n592 B.n591 71.676
R836 B.n585 B.n85 71.676
R837 B.n584 B.n583 71.676
R838 B.n577 B.n87 71.676
R839 B.n576 B.n91 71.676
R840 B.n572 B.n571 71.676
R841 B.n565 B.n93 71.676
R842 B.n564 B.n563 71.676
R843 B.n557 B.n95 71.676
R844 B.n556 B.n555 71.676
R845 B.n549 B.n97 71.676
R846 B.n548 B.n547 71.676
R847 B.n541 B.n99 71.676
R848 B.n540 B.n539 71.676
R849 B.n533 B.n101 71.676
R850 B.n532 B.n531 71.676
R851 B.n525 B.n103 71.676
R852 B.n524 B.n523 71.676
R853 B.n517 B.n105 71.676
R854 B.n516 B.n515 71.676
R855 B.n515 B.n514 71.676
R856 B.n518 B.n517 71.676
R857 B.n523 B.n522 71.676
R858 B.n526 B.n525 71.676
R859 B.n531 B.n530 71.676
R860 B.n534 B.n533 71.676
R861 B.n539 B.n538 71.676
R862 B.n542 B.n541 71.676
R863 B.n547 B.n546 71.676
R864 B.n550 B.n549 71.676
R865 B.n555 B.n554 71.676
R866 B.n558 B.n557 71.676
R867 B.n563 B.n562 71.676
R868 B.n566 B.n565 71.676
R869 B.n571 B.n570 71.676
R870 B.n573 B.n91 71.676
R871 B.n578 B.n577 71.676
R872 B.n583 B.n582 71.676
R873 B.n586 B.n585 71.676
R874 B.n591 B.n590 71.676
R875 B.n594 B.n593 71.676
R876 B.n600 B.n599 71.676
R877 B.n603 B.n602 71.676
R878 B.n608 B.n607 71.676
R879 B.n611 B.n610 71.676
R880 B.n616 B.n615 71.676
R881 B.n619 B.n618 71.676
R882 B.n624 B.n623 71.676
R883 B.n627 B.n626 71.676
R884 B.n632 B.n631 71.676
R885 B.n635 B.n634 71.676
R886 B.n640 B.n639 71.676
R887 B.n643 B.n642 71.676
R888 B.n648 B.n647 71.676
R889 B.n651 B.n650 71.676
R890 B.n656 B.n655 71.676
R891 B.n659 B.n658 71.676
R892 B.n361 B.n360 71.676
R893 B.n355 B.n175 71.676
R894 B.n353 B.n352 71.676
R895 B.n348 B.n347 71.676
R896 B.n345 B.n344 71.676
R897 B.n340 B.n339 71.676
R898 B.n337 B.n336 71.676
R899 B.n332 B.n331 71.676
R900 B.n329 B.n328 71.676
R901 B.n324 B.n323 71.676
R902 B.n321 B.n320 71.676
R903 B.n316 B.n315 71.676
R904 B.n313 B.n312 71.676
R905 B.n308 B.n307 71.676
R906 B.n305 B.n304 71.676
R907 B.n300 B.n299 71.676
R908 B.n295 B.n193 71.676
R909 B.n293 B.n292 71.676
R910 B.n288 B.n287 71.676
R911 B.n285 B.n284 71.676
R912 B.n279 B.n278 71.676
R913 B.n276 B.n275 71.676
R914 B.n271 B.n270 71.676
R915 B.n268 B.n267 71.676
R916 B.n263 B.n262 71.676
R917 B.n260 B.n259 71.676
R918 B.n255 B.n254 71.676
R919 B.n252 B.n251 71.676
R920 B.n247 B.n246 71.676
R921 B.n244 B.n243 71.676
R922 B.n239 B.n238 71.676
R923 B.n236 B.n235 71.676
R924 B.n231 B.n230 71.676
R925 B.n228 B.n227 71.676
R926 B.n223 B.n222 71.676
R927 B.n220 B.n219 71.676
R928 B.n215 B.n171 71.676
R929 B.n281 B.n199 59.5399
R930 B.n192 B.n191 59.5399
R931 B.n596 B.n83 59.5399
R932 B.n90 B.n89 59.5399
R933 B.n199 B.n198 56.4369
R934 B.n191 B.n190 56.4369
R935 B.n83 B.n82 56.4369
R936 B.n89 B.n88 56.4369
R937 B.n366 B.n168 52.2169
R938 B.n372 B.n168 52.2169
R939 B.n372 B.n164 52.2169
R940 B.n378 B.n164 52.2169
R941 B.n378 B.n160 52.2169
R942 B.n385 B.n160 52.2169
R943 B.n385 B.n384 52.2169
R944 B.n391 B.n153 52.2169
R945 B.n397 B.n153 52.2169
R946 B.n397 B.n149 52.2169
R947 B.n403 B.n149 52.2169
R948 B.n403 B.n145 52.2169
R949 B.n409 B.n145 52.2169
R950 B.n409 B.n141 52.2169
R951 B.n415 B.n141 52.2169
R952 B.n415 B.n137 52.2169
R953 B.n422 B.n137 52.2169
R954 B.n422 B.n421 52.2169
R955 B.n428 B.n130 52.2169
R956 B.n434 B.n130 52.2169
R957 B.n434 B.n126 52.2169
R958 B.n440 B.n126 52.2169
R959 B.n440 B.n122 52.2169
R960 B.n446 B.n122 52.2169
R961 B.n446 B.n118 52.2169
R962 B.n452 B.n118 52.2169
R963 B.n459 B.n114 52.2169
R964 B.n459 B.n110 52.2169
R965 B.n465 B.n110 52.2169
R966 B.n465 B.n4 52.2169
R967 B.n730 B.n4 52.2169
R968 B.n730 B.n729 52.2169
R969 B.n729 B.n728 52.2169
R970 B.n728 B.n8 52.2169
R971 B.n722 B.n8 52.2169
R972 B.n722 B.n721 52.2169
R973 B.n720 B.n15 52.2169
R974 B.n714 B.n15 52.2169
R975 B.n714 B.n713 52.2169
R976 B.n713 B.n712 52.2169
R977 B.n712 B.n22 52.2169
R978 B.n706 B.n22 52.2169
R979 B.n706 B.n705 52.2169
R980 B.n705 B.n704 52.2169
R981 B.n698 B.n32 52.2169
R982 B.n698 B.n697 52.2169
R983 B.n697 B.n696 52.2169
R984 B.n696 B.n36 52.2169
R985 B.n690 B.n36 52.2169
R986 B.n690 B.n689 52.2169
R987 B.n689 B.n688 52.2169
R988 B.n688 B.n43 52.2169
R989 B.n682 B.n43 52.2169
R990 B.n682 B.n681 52.2169
R991 B.n681 B.n680 52.2169
R992 B.n674 B.n53 52.2169
R993 B.n674 B.n673 52.2169
R994 B.n673 B.n672 52.2169
R995 B.n672 B.n57 52.2169
R996 B.n666 B.n57 52.2169
R997 B.n666 B.n665 52.2169
R998 B.n665 B.n664 52.2169
R999 B.t1 B.n114 46.0738
R1000 B.n721 B.t2 46.0738
R1001 B.n384 B.t5 41.4665
R1002 B.n53 B.t9 41.4665
R1003 B.n662 B.n661 32.6249
R1004 B.n512 B.n511 32.6249
R1005 B.n368 B.n170 32.6249
R1006 B.n364 B.n363 32.6249
R1007 B.n421 B.t3 29.1803
R1008 B.n32 B.t0 29.1803
R1009 B.n428 B.t3 23.0371
R1010 B.n704 B.t0 23.0371
R1011 B B.n732 18.0485
R1012 B.n391 B.t5 10.7509
R1013 B.n680 B.t9 10.7509
R1014 B.n661 B.n660 10.6151
R1015 B.n660 B.n66 10.6151
R1016 B.n654 B.n66 10.6151
R1017 B.n654 B.n653 10.6151
R1018 B.n653 B.n652 10.6151
R1019 B.n652 B.n68 10.6151
R1020 B.n646 B.n68 10.6151
R1021 B.n646 B.n645 10.6151
R1022 B.n645 B.n644 10.6151
R1023 B.n644 B.n70 10.6151
R1024 B.n638 B.n70 10.6151
R1025 B.n638 B.n637 10.6151
R1026 B.n637 B.n636 10.6151
R1027 B.n636 B.n72 10.6151
R1028 B.n630 B.n72 10.6151
R1029 B.n630 B.n629 10.6151
R1030 B.n629 B.n628 10.6151
R1031 B.n628 B.n74 10.6151
R1032 B.n622 B.n74 10.6151
R1033 B.n622 B.n621 10.6151
R1034 B.n621 B.n620 10.6151
R1035 B.n620 B.n76 10.6151
R1036 B.n614 B.n76 10.6151
R1037 B.n614 B.n613 10.6151
R1038 B.n613 B.n612 10.6151
R1039 B.n612 B.n78 10.6151
R1040 B.n606 B.n78 10.6151
R1041 B.n606 B.n605 10.6151
R1042 B.n605 B.n604 10.6151
R1043 B.n604 B.n80 10.6151
R1044 B.n598 B.n80 10.6151
R1045 B.n598 B.n597 10.6151
R1046 B.n595 B.n84 10.6151
R1047 B.n589 B.n84 10.6151
R1048 B.n589 B.n588 10.6151
R1049 B.n588 B.n587 10.6151
R1050 B.n587 B.n86 10.6151
R1051 B.n581 B.n86 10.6151
R1052 B.n581 B.n580 10.6151
R1053 B.n580 B.n579 10.6151
R1054 B.n575 B.n574 10.6151
R1055 B.n574 B.n92 10.6151
R1056 B.n569 B.n92 10.6151
R1057 B.n569 B.n568 10.6151
R1058 B.n568 B.n567 10.6151
R1059 B.n567 B.n94 10.6151
R1060 B.n561 B.n94 10.6151
R1061 B.n561 B.n560 10.6151
R1062 B.n560 B.n559 10.6151
R1063 B.n559 B.n96 10.6151
R1064 B.n553 B.n96 10.6151
R1065 B.n553 B.n552 10.6151
R1066 B.n552 B.n551 10.6151
R1067 B.n551 B.n98 10.6151
R1068 B.n545 B.n98 10.6151
R1069 B.n545 B.n544 10.6151
R1070 B.n544 B.n543 10.6151
R1071 B.n543 B.n100 10.6151
R1072 B.n537 B.n100 10.6151
R1073 B.n537 B.n536 10.6151
R1074 B.n536 B.n535 10.6151
R1075 B.n535 B.n102 10.6151
R1076 B.n529 B.n102 10.6151
R1077 B.n529 B.n528 10.6151
R1078 B.n528 B.n527 10.6151
R1079 B.n527 B.n104 10.6151
R1080 B.n521 B.n104 10.6151
R1081 B.n521 B.n520 10.6151
R1082 B.n520 B.n519 10.6151
R1083 B.n519 B.n106 10.6151
R1084 B.n513 B.n106 10.6151
R1085 B.n513 B.n512 10.6151
R1086 B.n369 B.n368 10.6151
R1087 B.n370 B.n369 10.6151
R1088 B.n370 B.n162 10.6151
R1089 B.n380 B.n162 10.6151
R1090 B.n381 B.n380 10.6151
R1091 B.n382 B.n381 10.6151
R1092 B.n382 B.n155 10.6151
R1093 B.n393 B.n155 10.6151
R1094 B.n394 B.n393 10.6151
R1095 B.n395 B.n394 10.6151
R1096 B.n395 B.n147 10.6151
R1097 B.n405 B.n147 10.6151
R1098 B.n406 B.n405 10.6151
R1099 B.n407 B.n406 10.6151
R1100 B.n407 B.n139 10.6151
R1101 B.n417 B.n139 10.6151
R1102 B.n418 B.n417 10.6151
R1103 B.n419 B.n418 10.6151
R1104 B.n419 B.n132 10.6151
R1105 B.n430 B.n132 10.6151
R1106 B.n431 B.n430 10.6151
R1107 B.n432 B.n431 10.6151
R1108 B.n432 B.n124 10.6151
R1109 B.n442 B.n124 10.6151
R1110 B.n443 B.n442 10.6151
R1111 B.n444 B.n443 10.6151
R1112 B.n444 B.n116 10.6151
R1113 B.n454 B.n116 10.6151
R1114 B.n455 B.n454 10.6151
R1115 B.n457 B.n455 10.6151
R1116 B.n457 B.n456 10.6151
R1117 B.n456 B.n108 10.6151
R1118 B.n468 B.n108 10.6151
R1119 B.n469 B.n468 10.6151
R1120 B.n470 B.n469 10.6151
R1121 B.n471 B.n470 10.6151
R1122 B.n473 B.n471 10.6151
R1123 B.n474 B.n473 10.6151
R1124 B.n475 B.n474 10.6151
R1125 B.n476 B.n475 10.6151
R1126 B.n478 B.n476 10.6151
R1127 B.n479 B.n478 10.6151
R1128 B.n480 B.n479 10.6151
R1129 B.n481 B.n480 10.6151
R1130 B.n483 B.n481 10.6151
R1131 B.n484 B.n483 10.6151
R1132 B.n485 B.n484 10.6151
R1133 B.n486 B.n485 10.6151
R1134 B.n488 B.n486 10.6151
R1135 B.n489 B.n488 10.6151
R1136 B.n490 B.n489 10.6151
R1137 B.n491 B.n490 10.6151
R1138 B.n493 B.n491 10.6151
R1139 B.n494 B.n493 10.6151
R1140 B.n495 B.n494 10.6151
R1141 B.n496 B.n495 10.6151
R1142 B.n498 B.n496 10.6151
R1143 B.n499 B.n498 10.6151
R1144 B.n500 B.n499 10.6151
R1145 B.n501 B.n500 10.6151
R1146 B.n503 B.n501 10.6151
R1147 B.n504 B.n503 10.6151
R1148 B.n505 B.n504 10.6151
R1149 B.n506 B.n505 10.6151
R1150 B.n508 B.n506 10.6151
R1151 B.n509 B.n508 10.6151
R1152 B.n510 B.n509 10.6151
R1153 B.n511 B.n510 10.6151
R1154 B.n363 B.n362 10.6151
R1155 B.n362 B.n174 10.6151
R1156 B.n357 B.n174 10.6151
R1157 B.n357 B.n356 10.6151
R1158 B.n356 B.n176 10.6151
R1159 B.n351 B.n176 10.6151
R1160 B.n351 B.n350 10.6151
R1161 B.n350 B.n349 10.6151
R1162 B.n349 B.n178 10.6151
R1163 B.n343 B.n178 10.6151
R1164 B.n343 B.n342 10.6151
R1165 B.n342 B.n341 10.6151
R1166 B.n341 B.n180 10.6151
R1167 B.n335 B.n180 10.6151
R1168 B.n335 B.n334 10.6151
R1169 B.n334 B.n333 10.6151
R1170 B.n333 B.n182 10.6151
R1171 B.n327 B.n182 10.6151
R1172 B.n327 B.n326 10.6151
R1173 B.n326 B.n325 10.6151
R1174 B.n325 B.n184 10.6151
R1175 B.n319 B.n184 10.6151
R1176 B.n319 B.n318 10.6151
R1177 B.n318 B.n317 10.6151
R1178 B.n317 B.n186 10.6151
R1179 B.n311 B.n186 10.6151
R1180 B.n311 B.n310 10.6151
R1181 B.n310 B.n309 10.6151
R1182 B.n309 B.n188 10.6151
R1183 B.n303 B.n188 10.6151
R1184 B.n303 B.n302 10.6151
R1185 B.n302 B.n301 10.6151
R1186 B.n297 B.n296 10.6151
R1187 B.n296 B.n194 10.6151
R1188 B.n291 B.n194 10.6151
R1189 B.n291 B.n290 10.6151
R1190 B.n290 B.n289 10.6151
R1191 B.n289 B.n196 10.6151
R1192 B.n283 B.n196 10.6151
R1193 B.n283 B.n282 10.6151
R1194 B.n280 B.n200 10.6151
R1195 B.n274 B.n200 10.6151
R1196 B.n274 B.n273 10.6151
R1197 B.n273 B.n272 10.6151
R1198 B.n272 B.n202 10.6151
R1199 B.n266 B.n202 10.6151
R1200 B.n266 B.n265 10.6151
R1201 B.n265 B.n264 10.6151
R1202 B.n264 B.n204 10.6151
R1203 B.n258 B.n204 10.6151
R1204 B.n258 B.n257 10.6151
R1205 B.n257 B.n256 10.6151
R1206 B.n256 B.n206 10.6151
R1207 B.n250 B.n206 10.6151
R1208 B.n250 B.n249 10.6151
R1209 B.n249 B.n248 10.6151
R1210 B.n248 B.n208 10.6151
R1211 B.n242 B.n208 10.6151
R1212 B.n242 B.n241 10.6151
R1213 B.n241 B.n240 10.6151
R1214 B.n240 B.n210 10.6151
R1215 B.n234 B.n210 10.6151
R1216 B.n234 B.n233 10.6151
R1217 B.n233 B.n232 10.6151
R1218 B.n232 B.n212 10.6151
R1219 B.n226 B.n212 10.6151
R1220 B.n226 B.n225 10.6151
R1221 B.n225 B.n224 10.6151
R1222 B.n224 B.n214 10.6151
R1223 B.n218 B.n214 10.6151
R1224 B.n218 B.n217 10.6151
R1225 B.n217 B.n170 10.6151
R1226 B.n364 B.n166 10.6151
R1227 B.n374 B.n166 10.6151
R1228 B.n375 B.n374 10.6151
R1229 B.n376 B.n375 10.6151
R1230 B.n376 B.n158 10.6151
R1231 B.n387 B.n158 10.6151
R1232 B.n388 B.n387 10.6151
R1233 B.n389 B.n388 10.6151
R1234 B.n389 B.n151 10.6151
R1235 B.n399 B.n151 10.6151
R1236 B.n400 B.n399 10.6151
R1237 B.n401 B.n400 10.6151
R1238 B.n401 B.n143 10.6151
R1239 B.n411 B.n143 10.6151
R1240 B.n412 B.n411 10.6151
R1241 B.n413 B.n412 10.6151
R1242 B.n413 B.n135 10.6151
R1243 B.n424 B.n135 10.6151
R1244 B.n425 B.n424 10.6151
R1245 B.n426 B.n425 10.6151
R1246 B.n426 B.n128 10.6151
R1247 B.n436 B.n128 10.6151
R1248 B.n437 B.n436 10.6151
R1249 B.n438 B.n437 10.6151
R1250 B.n438 B.n120 10.6151
R1251 B.n448 B.n120 10.6151
R1252 B.n449 B.n448 10.6151
R1253 B.n450 B.n449 10.6151
R1254 B.n450 B.n112 10.6151
R1255 B.n461 B.n112 10.6151
R1256 B.n462 B.n461 10.6151
R1257 B.n463 B.n462 10.6151
R1258 B.n463 B.n0 10.6151
R1259 B.n726 B.n1 10.6151
R1260 B.n726 B.n725 10.6151
R1261 B.n725 B.n724 10.6151
R1262 B.n724 B.n10 10.6151
R1263 B.n718 B.n10 10.6151
R1264 B.n718 B.n717 10.6151
R1265 B.n717 B.n716 10.6151
R1266 B.n716 B.n17 10.6151
R1267 B.n710 B.n17 10.6151
R1268 B.n710 B.n709 10.6151
R1269 B.n709 B.n708 10.6151
R1270 B.n708 B.n24 10.6151
R1271 B.n702 B.n24 10.6151
R1272 B.n702 B.n701 10.6151
R1273 B.n701 B.n700 10.6151
R1274 B.n700 B.n30 10.6151
R1275 B.n694 B.n30 10.6151
R1276 B.n694 B.n693 10.6151
R1277 B.n693 B.n692 10.6151
R1278 B.n692 B.n38 10.6151
R1279 B.n686 B.n38 10.6151
R1280 B.n686 B.n685 10.6151
R1281 B.n685 B.n684 10.6151
R1282 B.n684 B.n45 10.6151
R1283 B.n678 B.n45 10.6151
R1284 B.n678 B.n677 10.6151
R1285 B.n677 B.n676 10.6151
R1286 B.n676 B.n51 10.6151
R1287 B.n670 B.n51 10.6151
R1288 B.n670 B.n669 10.6151
R1289 B.n669 B.n668 10.6151
R1290 B.n668 B.n59 10.6151
R1291 B.n662 B.n59 10.6151
R1292 B.n596 B.n595 6.5566
R1293 B.n579 B.n90 6.5566
R1294 B.n297 B.n192 6.5566
R1295 B.n282 B.n281 6.5566
R1296 B.n452 B.t1 6.14361
R1297 B.t2 B.n720 6.14361
R1298 B.n597 B.n596 4.05904
R1299 B.n575 B.n90 4.05904
R1300 B.n301 B.n192 4.05904
R1301 B.n281 B.n280 4.05904
R1302 B.n732 B.n0 2.81026
R1303 B.n732 B.n1 2.81026
R1304 VN.n0 VN.t3 120.582
R1305 VN.n1 VN.t1 120.582
R1306 VN.n0 VN.t0 119.811
R1307 VN.n1 VN.t2 119.811
R1308 VN VN.n1 48.6699
R1309 VN VN.n0 4.37066
R1310 VDD2.n2 VDD2.n0 105.549
R1311 VDD2.n2 VDD2.n1 66.5071
R1312 VDD2.n1 VDD2.t1 2.18835
R1313 VDD2.n1 VDD2.t2 2.18835
R1314 VDD2.n0 VDD2.t0 2.18835
R1315 VDD2.n0 VDD2.t3 2.18835
R1316 VDD2 VDD2.n2 0.0586897
C0 VDD2 VDD1 1.01786f
C1 VDD2 VP 0.393168f
C2 VDD2 VN 3.65117f
C3 VDD2 VTAIL 4.7546f
C4 VP VDD1 3.89448f
C5 VDD1 VN 0.149117f
C6 VP VN 5.62921f
C7 VTAIL VDD1 4.70052f
C8 VTAIL VP 3.70553f
C9 VTAIL VN 3.69142f
C10 VDD2 B 3.539727f
C11 VDD1 B 7.39061f
C12 VTAIL B 8.296496f
C13 VN B 10.41855f
C14 VP B 8.689119f
C15 VDD2.t0 B 0.196001f
C16 VDD2.t3 B 0.196001f
C17 VDD2.n0 B 2.27068f
C18 VDD2.t1 B 0.196001f
C19 VDD2.t2 B 0.196001f
C20 VDD2.n1 B 1.71576f
C21 VDD2.n2 B 3.50212f
C22 VN.t3 B 1.90961f
C23 VN.t0 B 1.90478f
C24 VN.n0 B 1.20332f
C25 VN.t1 B 1.90961f
C26 VN.t2 B 1.90478f
C27 VN.n1 B 2.54268f
C28 VDD1.t0 B 0.195973f
C29 VDD1.t1 B 0.195973f
C30 VDD1.n0 B 1.71592f
C31 VDD1.t2 B 0.195973f
C32 VDD1.t3 B 0.195973f
C33 VDD1.n1 B 2.29549f
C34 VTAIL.t6 B 1.33501f
C35 VTAIL.n0 B 0.314759f
C36 VTAIL.t3 B 1.33501f
C37 VTAIL.n1 B 0.382058f
C38 VTAIL.t2 B 1.33501f
C39 VTAIL.n2 B 1.17292f
C40 VTAIL.t7 B 1.33501f
C41 VTAIL.n3 B 1.17292f
C42 VTAIL.t1 B 1.33501f
C43 VTAIL.n4 B 0.382055f
C44 VTAIL.t5 B 1.33501f
C45 VTAIL.n5 B 0.382055f
C46 VTAIL.t4 B 1.33501f
C47 VTAIL.n6 B 1.17292f
C48 VTAIL.t0 B 1.33501f
C49 VTAIL.n7 B 1.09907f
C50 VP.n0 B 0.035732f
C51 VP.t0 B 1.70813f
C52 VP.n1 B 0.039565f
C53 VP.n2 B 0.027103f
C54 VP.t1 B 1.70813f
C55 VP.n3 B 0.706353f
C56 VP.t2 B 1.93967f
C57 VP.t3 B 1.94459f
C58 VP.n4 B 2.57493f
C59 VP.n5 B 1.40149f
C60 VP.n6 B 0.035732f
C61 VP.n7 B 0.035798f
C62 VP.n8 B 0.050512f
C63 VP.n9 B 0.039565f
C64 VP.n10 B 0.027103f
C65 VP.n11 B 0.027103f
C66 VP.n12 B 0.027103f
C67 VP.n13 B 0.050512f
C68 VP.n14 B 0.035798f
C69 VP.n15 B 0.706353f
C70 VP.n16 B 0.043896f
.ends

