* NGSPICE file created from diff_pair_sample_0025.ext - technology: sky130A

.subckt diff_pair_sample_0025 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t8 B.t19 sky130_fd_pr__nfet_01v8 ad=2.0241 pd=11.16 as=0.85635 ps=5.52 w=5.19 l=0.99
X1 VTAIL.t5 VN.t1 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.85635 pd=5.52 as=0.85635 ps=5.52 w=5.19 l=0.99
X2 B.t18 B.t16 B.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=2.0241 pd=11.16 as=0 ps=0 w=5.19 l=0.99
X3 VDD2.t3 VN.t2 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=0.85635 pd=5.52 as=2.0241 ps=11.16 w=5.19 l=0.99
X4 VTAIL.t1 VP.t0 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.85635 pd=5.52 as=0.85635 ps=5.52 w=5.19 l=0.99
X5 VDD1.t4 VP.t1 VTAIL.t11 B.t19 sky130_fd_pr__nfet_01v8 ad=2.0241 pd=11.16 as=0.85635 ps=5.52 w=5.19 l=0.99
X6 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=2.0241 pd=11.16 as=0 ps=0 w=5.19 l=0.99
X7 VTAIL.t7 VN.t3 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=0.85635 pd=5.52 as=0.85635 ps=5.52 w=5.19 l=0.99
X8 VTAIL.t3 VP.t2 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.85635 pd=5.52 as=0.85635 ps=5.52 w=5.19 l=0.99
X9 VDD1.t2 VP.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.0241 pd=11.16 as=0.85635 ps=5.52 w=5.19 l=0.99
X10 VDD2.t1 VN.t4 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.85635 pd=5.52 as=2.0241 ps=11.16 w=5.19 l=0.99
X11 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=2.0241 pd=11.16 as=0 ps=0 w=5.19 l=0.99
X12 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=2.0241 pd=11.16 as=0 ps=0 w=5.19 l=0.99
X13 VDD2.t0 VN.t5 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=2.0241 pd=11.16 as=0.85635 ps=5.52 w=5.19 l=0.99
X14 VDD1.t1 VP.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.85635 pd=5.52 as=2.0241 ps=11.16 w=5.19 l=0.99
X15 VDD1.t0 VP.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.85635 pd=5.52 as=2.0241 ps=11.16 w=5.19 l=0.99
R0 VN.n1 VN.t5 188.536
R1 VN.n7 VN.t4 188.536
R2 VN.n4 VN.t2 166.267
R3 VN.n10 VN.t0 166.267
R4 VN.n9 VN.n6 161.3
R5 VN.n3 VN.n0 161.3
R6 VN.n2 VN.t1 126.343
R7 VN.n8 VN.t3 126.343
R8 VN.n11 VN.n10 80.6037
R9 VN.n5 VN.n4 80.6037
R10 VN.n4 VN.n3 47.4702
R11 VN.n10 VN.n9 47.4702
R12 VN VN.n11 37.5672
R13 VN.n2 VN.n1 32.1379
R14 VN.n8 VN.n7 32.1379
R15 VN.n7 VN.n6 28.4787
R16 VN.n1 VN.n0 28.4787
R17 VN.n3 VN.n2 24.9531
R18 VN.n9 VN.n8 24.9531
R19 VN.n11 VN.n6 0.285035
R20 VN.n5 VN.n0 0.285035
R21 VN VN.n5 0.146778
R22 VTAIL.n114 VTAIL.n92 289.615
R23 VTAIL.n24 VTAIL.n2 289.615
R24 VTAIL.n86 VTAIL.n64 289.615
R25 VTAIL.n56 VTAIL.n34 289.615
R26 VTAIL.n100 VTAIL.n99 185
R27 VTAIL.n105 VTAIL.n104 185
R28 VTAIL.n107 VTAIL.n106 185
R29 VTAIL.n96 VTAIL.n95 185
R30 VTAIL.n113 VTAIL.n112 185
R31 VTAIL.n115 VTAIL.n114 185
R32 VTAIL.n10 VTAIL.n9 185
R33 VTAIL.n15 VTAIL.n14 185
R34 VTAIL.n17 VTAIL.n16 185
R35 VTAIL.n6 VTAIL.n5 185
R36 VTAIL.n23 VTAIL.n22 185
R37 VTAIL.n25 VTAIL.n24 185
R38 VTAIL.n87 VTAIL.n86 185
R39 VTAIL.n85 VTAIL.n84 185
R40 VTAIL.n68 VTAIL.n67 185
R41 VTAIL.n79 VTAIL.n78 185
R42 VTAIL.n77 VTAIL.n76 185
R43 VTAIL.n72 VTAIL.n71 185
R44 VTAIL.n57 VTAIL.n56 185
R45 VTAIL.n55 VTAIL.n54 185
R46 VTAIL.n38 VTAIL.n37 185
R47 VTAIL.n49 VTAIL.n48 185
R48 VTAIL.n47 VTAIL.n46 185
R49 VTAIL.n42 VTAIL.n41 185
R50 VTAIL.n101 VTAIL.t10 147.672
R51 VTAIL.n11 VTAIL.t0 147.672
R52 VTAIL.n73 VTAIL.t2 147.672
R53 VTAIL.n43 VTAIL.t6 147.672
R54 VTAIL.n105 VTAIL.n99 104.615
R55 VTAIL.n106 VTAIL.n105 104.615
R56 VTAIL.n106 VTAIL.n95 104.615
R57 VTAIL.n113 VTAIL.n95 104.615
R58 VTAIL.n114 VTAIL.n113 104.615
R59 VTAIL.n15 VTAIL.n9 104.615
R60 VTAIL.n16 VTAIL.n15 104.615
R61 VTAIL.n16 VTAIL.n5 104.615
R62 VTAIL.n23 VTAIL.n5 104.615
R63 VTAIL.n24 VTAIL.n23 104.615
R64 VTAIL.n86 VTAIL.n85 104.615
R65 VTAIL.n85 VTAIL.n67 104.615
R66 VTAIL.n78 VTAIL.n67 104.615
R67 VTAIL.n78 VTAIL.n77 104.615
R68 VTAIL.n77 VTAIL.n71 104.615
R69 VTAIL.n56 VTAIL.n55 104.615
R70 VTAIL.n55 VTAIL.n37 104.615
R71 VTAIL.n48 VTAIL.n37 104.615
R72 VTAIL.n48 VTAIL.n47 104.615
R73 VTAIL.n47 VTAIL.n41 104.615
R74 VTAIL.t10 VTAIL.n99 52.3082
R75 VTAIL.t0 VTAIL.n9 52.3082
R76 VTAIL.t2 VTAIL.n71 52.3082
R77 VTAIL.t6 VTAIL.n41 52.3082
R78 VTAIL.n63 VTAIL.n62 50.231
R79 VTAIL.n33 VTAIL.n32 50.231
R80 VTAIL.n1 VTAIL.n0 50.2309
R81 VTAIL.n31 VTAIL.n30 50.2309
R82 VTAIL.n119 VTAIL.n118 30.4399
R83 VTAIL.n29 VTAIL.n28 30.4399
R84 VTAIL.n91 VTAIL.n90 30.4399
R85 VTAIL.n61 VTAIL.n60 30.4399
R86 VTAIL.n33 VTAIL.n31 19.1169
R87 VTAIL.n119 VTAIL.n91 17.9789
R88 VTAIL.n101 VTAIL.n100 15.6666
R89 VTAIL.n11 VTAIL.n10 15.6666
R90 VTAIL.n73 VTAIL.n72 15.6666
R91 VTAIL.n43 VTAIL.n42 15.6666
R92 VTAIL.n104 VTAIL.n103 12.8005
R93 VTAIL.n14 VTAIL.n13 12.8005
R94 VTAIL.n76 VTAIL.n75 12.8005
R95 VTAIL.n46 VTAIL.n45 12.8005
R96 VTAIL.n107 VTAIL.n98 12.0247
R97 VTAIL.n17 VTAIL.n8 12.0247
R98 VTAIL.n79 VTAIL.n70 12.0247
R99 VTAIL.n49 VTAIL.n40 12.0247
R100 VTAIL.n108 VTAIL.n96 11.249
R101 VTAIL.n18 VTAIL.n6 11.249
R102 VTAIL.n80 VTAIL.n68 11.249
R103 VTAIL.n50 VTAIL.n38 11.249
R104 VTAIL.n112 VTAIL.n111 10.4732
R105 VTAIL.n22 VTAIL.n21 10.4732
R106 VTAIL.n84 VTAIL.n83 10.4732
R107 VTAIL.n54 VTAIL.n53 10.4732
R108 VTAIL.n115 VTAIL.n94 9.69747
R109 VTAIL.n25 VTAIL.n4 9.69747
R110 VTAIL.n87 VTAIL.n66 9.69747
R111 VTAIL.n57 VTAIL.n36 9.69747
R112 VTAIL.n118 VTAIL.n117 9.45567
R113 VTAIL.n28 VTAIL.n27 9.45567
R114 VTAIL.n90 VTAIL.n89 9.45567
R115 VTAIL.n60 VTAIL.n59 9.45567
R116 VTAIL.n117 VTAIL.n116 9.3005
R117 VTAIL.n94 VTAIL.n93 9.3005
R118 VTAIL.n111 VTAIL.n110 9.3005
R119 VTAIL.n109 VTAIL.n108 9.3005
R120 VTAIL.n98 VTAIL.n97 9.3005
R121 VTAIL.n103 VTAIL.n102 9.3005
R122 VTAIL.n27 VTAIL.n26 9.3005
R123 VTAIL.n4 VTAIL.n3 9.3005
R124 VTAIL.n21 VTAIL.n20 9.3005
R125 VTAIL.n19 VTAIL.n18 9.3005
R126 VTAIL.n8 VTAIL.n7 9.3005
R127 VTAIL.n13 VTAIL.n12 9.3005
R128 VTAIL.n89 VTAIL.n88 9.3005
R129 VTAIL.n66 VTAIL.n65 9.3005
R130 VTAIL.n83 VTAIL.n82 9.3005
R131 VTAIL.n81 VTAIL.n80 9.3005
R132 VTAIL.n70 VTAIL.n69 9.3005
R133 VTAIL.n75 VTAIL.n74 9.3005
R134 VTAIL.n59 VTAIL.n58 9.3005
R135 VTAIL.n36 VTAIL.n35 9.3005
R136 VTAIL.n53 VTAIL.n52 9.3005
R137 VTAIL.n51 VTAIL.n50 9.3005
R138 VTAIL.n40 VTAIL.n39 9.3005
R139 VTAIL.n45 VTAIL.n44 9.3005
R140 VTAIL.n116 VTAIL.n92 8.92171
R141 VTAIL.n26 VTAIL.n2 8.92171
R142 VTAIL.n88 VTAIL.n64 8.92171
R143 VTAIL.n58 VTAIL.n34 8.92171
R144 VTAIL.n118 VTAIL.n92 5.04292
R145 VTAIL.n28 VTAIL.n2 5.04292
R146 VTAIL.n90 VTAIL.n64 5.04292
R147 VTAIL.n60 VTAIL.n34 5.04292
R148 VTAIL.n102 VTAIL.n101 4.38687
R149 VTAIL.n12 VTAIL.n11 4.38687
R150 VTAIL.n74 VTAIL.n73 4.38687
R151 VTAIL.n44 VTAIL.n43 4.38687
R152 VTAIL.n116 VTAIL.n115 4.26717
R153 VTAIL.n26 VTAIL.n25 4.26717
R154 VTAIL.n88 VTAIL.n87 4.26717
R155 VTAIL.n58 VTAIL.n57 4.26717
R156 VTAIL.n0 VTAIL.t9 3.81553
R157 VTAIL.n0 VTAIL.t5 3.81553
R158 VTAIL.n30 VTAIL.t11 3.81553
R159 VTAIL.n30 VTAIL.t3 3.81553
R160 VTAIL.n62 VTAIL.t4 3.81553
R161 VTAIL.n62 VTAIL.t1 3.81553
R162 VTAIL.n32 VTAIL.t8 3.81553
R163 VTAIL.n32 VTAIL.t7 3.81553
R164 VTAIL.n112 VTAIL.n94 3.49141
R165 VTAIL.n22 VTAIL.n4 3.49141
R166 VTAIL.n84 VTAIL.n66 3.49141
R167 VTAIL.n54 VTAIL.n36 3.49141
R168 VTAIL.n111 VTAIL.n96 2.71565
R169 VTAIL.n21 VTAIL.n6 2.71565
R170 VTAIL.n83 VTAIL.n68 2.71565
R171 VTAIL.n53 VTAIL.n38 2.71565
R172 VTAIL.n108 VTAIL.n107 1.93989
R173 VTAIL.n18 VTAIL.n17 1.93989
R174 VTAIL.n80 VTAIL.n79 1.93989
R175 VTAIL.n50 VTAIL.n49 1.93989
R176 VTAIL.n104 VTAIL.n98 1.16414
R177 VTAIL.n14 VTAIL.n8 1.16414
R178 VTAIL.n76 VTAIL.n70 1.16414
R179 VTAIL.n46 VTAIL.n40 1.16414
R180 VTAIL.n61 VTAIL.n33 1.13843
R181 VTAIL.n91 VTAIL.n63 1.13843
R182 VTAIL.n31 VTAIL.n29 1.13843
R183 VTAIL.n63 VTAIL.n61 1.03929
R184 VTAIL.n29 VTAIL.n1 1.03929
R185 VTAIL VTAIL.n119 0.795759
R186 VTAIL.n103 VTAIL.n100 0.388379
R187 VTAIL.n13 VTAIL.n10 0.388379
R188 VTAIL.n75 VTAIL.n72 0.388379
R189 VTAIL.n45 VTAIL.n42 0.388379
R190 VTAIL VTAIL.n1 0.343172
R191 VTAIL.n102 VTAIL.n97 0.155672
R192 VTAIL.n109 VTAIL.n97 0.155672
R193 VTAIL.n110 VTAIL.n109 0.155672
R194 VTAIL.n110 VTAIL.n93 0.155672
R195 VTAIL.n117 VTAIL.n93 0.155672
R196 VTAIL.n12 VTAIL.n7 0.155672
R197 VTAIL.n19 VTAIL.n7 0.155672
R198 VTAIL.n20 VTAIL.n19 0.155672
R199 VTAIL.n20 VTAIL.n3 0.155672
R200 VTAIL.n27 VTAIL.n3 0.155672
R201 VTAIL.n89 VTAIL.n65 0.155672
R202 VTAIL.n82 VTAIL.n65 0.155672
R203 VTAIL.n82 VTAIL.n81 0.155672
R204 VTAIL.n81 VTAIL.n69 0.155672
R205 VTAIL.n74 VTAIL.n69 0.155672
R206 VTAIL.n59 VTAIL.n35 0.155672
R207 VTAIL.n52 VTAIL.n35 0.155672
R208 VTAIL.n52 VTAIL.n51 0.155672
R209 VTAIL.n51 VTAIL.n39 0.155672
R210 VTAIL.n44 VTAIL.n39 0.155672
R211 VDD2.n51 VDD2.n29 289.615
R212 VDD2.n22 VDD2.n0 289.615
R213 VDD2.n52 VDD2.n51 185
R214 VDD2.n50 VDD2.n49 185
R215 VDD2.n33 VDD2.n32 185
R216 VDD2.n44 VDD2.n43 185
R217 VDD2.n42 VDD2.n41 185
R218 VDD2.n37 VDD2.n36 185
R219 VDD2.n8 VDD2.n7 185
R220 VDD2.n13 VDD2.n12 185
R221 VDD2.n15 VDD2.n14 185
R222 VDD2.n4 VDD2.n3 185
R223 VDD2.n21 VDD2.n20 185
R224 VDD2.n23 VDD2.n22 185
R225 VDD2.n38 VDD2.t5 147.672
R226 VDD2.n9 VDD2.t0 147.672
R227 VDD2.n51 VDD2.n50 104.615
R228 VDD2.n50 VDD2.n32 104.615
R229 VDD2.n43 VDD2.n32 104.615
R230 VDD2.n43 VDD2.n42 104.615
R231 VDD2.n42 VDD2.n36 104.615
R232 VDD2.n13 VDD2.n7 104.615
R233 VDD2.n14 VDD2.n13 104.615
R234 VDD2.n14 VDD2.n3 104.615
R235 VDD2.n21 VDD2.n3 104.615
R236 VDD2.n22 VDD2.n21 104.615
R237 VDD2.n28 VDD2.n27 67.1388
R238 VDD2 VDD2.n57 67.1359
R239 VDD2.t5 VDD2.n36 52.3082
R240 VDD2.t0 VDD2.n7 52.3082
R241 VDD2.n28 VDD2.n26 47.9168
R242 VDD2.n56 VDD2.n55 47.1187
R243 VDD2.n56 VDD2.n28 31.8877
R244 VDD2.n38 VDD2.n37 15.6666
R245 VDD2.n9 VDD2.n8 15.6666
R246 VDD2.n41 VDD2.n40 12.8005
R247 VDD2.n12 VDD2.n11 12.8005
R248 VDD2.n44 VDD2.n35 12.0247
R249 VDD2.n15 VDD2.n6 12.0247
R250 VDD2.n45 VDD2.n33 11.249
R251 VDD2.n16 VDD2.n4 11.249
R252 VDD2.n49 VDD2.n48 10.4732
R253 VDD2.n20 VDD2.n19 10.4732
R254 VDD2.n52 VDD2.n31 9.69747
R255 VDD2.n23 VDD2.n2 9.69747
R256 VDD2.n55 VDD2.n54 9.45567
R257 VDD2.n26 VDD2.n25 9.45567
R258 VDD2.n54 VDD2.n53 9.3005
R259 VDD2.n31 VDD2.n30 9.3005
R260 VDD2.n48 VDD2.n47 9.3005
R261 VDD2.n46 VDD2.n45 9.3005
R262 VDD2.n35 VDD2.n34 9.3005
R263 VDD2.n40 VDD2.n39 9.3005
R264 VDD2.n25 VDD2.n24 9.3005
R265 VDD2.n2 VDD2.n1 9.3005
R266 VDD2.n19 VDD2.n18 9.3005
R267 VDD2.n17 VDD2.n16 9.3005
R268 VDD2.n6 VDD2.n5 9.3005
R269 VDD2.n11 VDD2.n10 9.3005
R270 VDD2.n53 VDD2.n29 8.92171
R271 VDD2.n24 VDD2.n0 8.92171
R272 VDD2.n55 VDD2.n29 5.04292
R273 VDD2.n26 VDD2.n0 5.04292
R274 VDD2.n39 VDD2.n38 4.38687
R275 VDD2.n10 VDD2.n9 4.38687
R276 VDD2.n53 VDD2.n52 4.26717
R277 VDD2.n24 VDD2.n23 4.26717
R278 VDD2.n57 VDD2.t2 3.81553
R279 VDD2.n57 VDD2.t1 3.81553
R280 VDD2.n27 VDD2.t4 3.81553
R281 VDD2.n27 VDD2.t3 3.81553
R282 VDD2.n49 VDD2.n31 3.49141
R283 VDD2.n20 VDD2.n2 3.49141
R284 VDD2.n48 VDD2.n33 2.71565
R285 VDD2.n19 VDD2.n4 2.71565
R286 VDD2.n45 VDD2.n44 1.93989
R287 VDD2.n16 VDD2.n15 1.93989
R288 VDD2.n41 VDD2.n35 1.16414
R289 VDD2.n12 VDD2.n6 1.16414
R290 VDD2 VDD2.n56 0.912138
R291 VDD2.n40 VDD2.n37 0.388379
R292 VDD2.n11 VDD2.n8 0.388379
R293 VDD2.n54 VDD2.n30 0.155672
R294 VDD2.n47 VDD2.n30 0.155672
R295 VDD2.n47 VDD2.n46 0.155672
R296 VDD2.n46 VDD2.n34 0.155672
R297 VDD2.n39 VDD2.n34 0.155672
R298 VDD2.n10 VDD2.n5 0.155672
R299 VDD2.n17 VDD2.n5 0.155672
R300 VDD2.n18 VDD2.n17 0.155672
R301 VDD2.n18 VDD2.n1 0.155672
R302 VDD2.n25 VDD2.n1 0.155672
R303 B.n463 B.n462 585
R304 B.n464 B.n463 585
R305 B.n178 B.n72 585
R306 B.n177 B.n176 585
R307 B.n175 B.n174 585
R308 B.n173 B.n172 585
R309 B.n171 B.n170 585
R310 B.n169 B.n168 585
R311 B.n167 B.n166 585
R312 B.n165 B.n164 585
R313 B.n163 B.n162 585
R314 B.n161 B.n160 585
R315 B.n159 B.n158 585
R316 B.n157 B.n156 585
R317 B.n155 B.n154 585
R318 B.n153 B.n152 585
R319 B.n151 B.n150 585
R320 B.n149 B.n148 585
R321 B.n147 B.n146 585
R322 B.n145 B.n144 585
R323 B.n143 B.n142 585
R324 B.n141 B.n140 585
R325 B.n139 B.n138 585
R326 B.n136 B.n135 585
R327 B.n134 B.n133 585
R328 B.n132 B.n131 585
R329 B.n130 B.n129 585
R330 B.n128 B.n127 585
R331 B.n126 B.n125 585
R332 B.n124 B.n123 585
R333 B.n122 B.n121 585
R334 B.n120 B.n119 585
R335 B.n118 B.n117 585
R336 B.n116 B.n115 585
R337 B.n114 B.n113 585
R338 B.n112 B.n111 585
R339 B.n110 B.n109 585
R340 B.n108 B.n107 585
R341 B.n106 B.n105 585
R342 B.n104 B.n103 585
R343 B.n102 B.n101 585
R344 B.n100 B.n99 585
R345 B.n98 B.n97 585
R346 B.n96 B.n95 585
R347 B.n94 B.n93 585
R348 B.n92 B.n91 585
R349 B.n90 B.n89 585
R350 B.n88 B.n87 585
R351 B.n86 B.n85 585
R352 B.n84 B.n83 585
R353 B.n82 B.n81 585
R354 B.n80 B.n79 585
R355 B.n46 B.n45 585
R356 B.n467 B.n466 585
R357 B.n461 B.n73 585
R358 B.n73 B.n43 585
R359 B.n460 B.n42 585
R360 B.n471 B.n42 585
R361 B.n459 B.n41 585
R362 B.n472 B.n41 585
R363 B.n458 B.n40 585
R364 B.n473 B.n40 585
R365 B.n457 B.n456 585
R366 B.n456 B.n36 585
R367 B.n455 B.n35 585
R368 B.n479 B.n35 585
R369 B.n454 B.n34 585
R370 B.n480 B.n34 585
R371 B.n453 B.n33 585
R372 B.n481 B.n33 585
R373 B.n452 B.n451 585
R374 B.n451 B.n29 585
R375 B.n450 B.n28 585
R376 B.n487 B.n28 585
R377 B.n449 B.n27 585
R378 B.n488 B.n27 585
R379 B.n448 B.n26 585
R380 B.n489 B.n26 585
R381 B.n447 B.n446 585
R382 B.n446 B.n25 585
R383 B.n445 B.n21 585
R384 B.n495 B.n21 585
R385 B.n444 B.n20 585
R386 B.n496 B.n20 585
R387 B.n443 B.n19 585
R388 B.n497 B.n19 585
R389 B.n442 B.n441 585
R390 B.n441 B.n18 585
R391 B.n440 B.n14 585
R392 B.n503 B.n14 585
R393 B.n439 B.n13 585
R394 B.n504 B.n13 585
R395 B.n438 B.n12 585
R396 B.n505 B.n12 585
R397 B.n437 B.n436 585
R398 B.n436 B.n435 585
R399 B.n434 B.n433 585
R400 B.n434 B.n8 585
R401 B.n432 B.n7 585
R402 B.n512 B.n7 585
R403 B.n431 B.n6 585
R404 B.n513 B.n6 585
R405 B.n430 B.n5 585
R406 B.n514 B.n5 585
R407 B.n429 B.n428 585
R408 B.n428 B.n4 585
R409 B.n427 B.n179 585
R410 B.n427 B.n426 585
R411 B.n417 B.n180 585
R412 B.n181 B.n180 585
R413 B.n419 B.n418 585
R414 B.n420 B.n419 585
R415 B.n416 B.n186 585
R416 B.n186 B.n185 585
R417 B.n415 B.n414 585
R418 B.n414 B.n413 585
R419 B.n188 B.n187 585
R420 B.n406 B.n188 585
R421 B.n405 B.n404 585
R422 B.n407 B.n405 585
R423 B.n403 B.n193 585
R424 B.n193 B.n192 585
R425 B.n402 B.n401 585
R426 B.n401 B.n400 585
R427 B.n195 B.n194 585
R428 B.n393 B.n195 585
R429 B.n392 B.n391 585
R430 B.n394 B.n392 585
R431 B.n390 B.n200 585
R432 B.n200 B.n199 585
R433 B.n389 B.n388 585
R434 B.n388 B.n387 585
R435 B.n202 B.n201 585
R436 B.n203 B.n202 585
R437 B.n380 B.n379 585
R438 B.n381 B.n380 585
R439 B.n378 B.n208 585
R440 B.n208 B.n207 585
R441 B.n377 B.n376 585
R442 B.n376 B.n375 585
R443 B.n210 B.n209 585
R444 B.n211 B.n210 585
R445 B.n368 B.n367 585
R446 B.n369 B.n368 585
R447 B.n366 B.n216 585
R448 B.n216 B.n215 585
R449 B.n365 B.n364 585
R450 B.n364 B.n363 585
R451 B.n218 B.n217 585
R452 B.n219 B.n218 585
R453 B.n359 B.n358 585
R454 B.n222 B.n221 585
R455 B.n355 B.n354 585
R456 B.n356 B.n355 585
R457 B.n353 B.n248 585
R458 B.n352 B.n351 585
R459 B.n350 B.n349 585
R460 B.n348 B.n347 585
R461 B.n346 B.n345 585
R462 B.n344 B.n343 585
R463 B.n342 B.n341 585
R464 B.n340 B.n339 585
R465 B.n338 B.n337 585
R466 B.n336 B.n335 585
R467 B.n334 B.n333 585
R468 B.n332 B.n331 585
R469 B.n330 B.n329 585
R470 B.n328 B.n327 585
R471 B.n326 B.n325 585
R472 B.n324 B.n323 585
R473 B.n322 B.n321 585
R474 B.n320 B.n319 585
R475 B.n318 B.n317 585
R476 B.n315 B.n314 585
R477 B.n313 B.n312 585
R478 B.n311 B.n310 585
R479 B.n309 B.n308 585
R480 B.n307 B.n306 585
R481 B.n305 B.n304 585
R482 B.n303 B.n302 585
R483 B.n301 B.n300 585
R484 B.n299 B.n298 585
R485 B.n297 B.n296 585
R486 B.n295 B.n294 585
R487 B.n293 B.n292 585
R488 B.n291 B.n290 585
R489 B.n289 B.n288 585
R490 B.n287 B.n286 585
R491 B.n285 B.n284 585
R492 B.n283 B.n282 585
R493 B.n281 B.n280 585
R494 B.n279 B.n278 585
R495 B.n277 B.n276 585
R496 B.n275 B.n274 585
R497 B.n273 B.n272 585
R498 B.n271 B.n270 585
R499 B.n269 B.n268 585
R500 B.n267 B.n266 585
R501 B.n265 B.n264 585
R502 B.n263 B.n262 585
R503 B.n261 B.n260 585
R504 B.n259 B.n258 585
R505 B.n257 B.n256 585
R506 B.n255 B.n254 585
R507 B.n360 B.n220 585
R508 B.n220 B.n219 585
R509 B.n362 B.n361 585
R510 B.n363 B.n362 585
R511 B.n214 B.n213 585
R512 B.n215 B.n214 585
R513 B.n371 B.n370 585
R514 B.n370 B.n369 585
R515 B.n372 B.n212 585
R516 B.n212 B.n211 585
R517 B.n374 B.n373 585
R518 B.n375 B.n374 585
R519 B.n206 B.n205 585
R520 B.n207 B.n206 585
R521 B.n383 B.n382 585
R522 B.n382 B.n381 585
R523 B.n384 B.n204 585
R524 B.n204 B.n203 585
R525 B.n386 B.n385 585
R526 B.n387 B.n386 585
R527 B.n198 B.n197 585
R528 B.n199 B.n198 585
R529 B.n396 B.n395 585
R530 B.n395 B.n394 585
R531 B.n397 B.n196 585
R532 B.n393 B.n196 585
R533 B.n399 B.n398 585
R534 B.n400 B.n399 585
R535 B.n191 B.n190 585
R536 B.n192 B.n191 585
R537 B.n409 B.n408 585
R538 B.n408 B.n407 585
R539 B.n410 B.n189 585
R540 B.n406 B.n189 585
R541 B.n412 B.n411 585
R542 B.n413 B.n412 585
R543 B.n184 B.n183 585
R544 B.n185 B.n184 585
R545 B.n422 B.n421 585
R546 B.n421 B.n420 585
R547 B.n423 B.n182 585
R548 B.n182 B.n181 585
R549 B.n425 B.n424 585
R550 B.n426 B.n425 585
R551 B.n3 B.n0 585
R552 B.n4 B.n3 585
R553 B.n511 B.n1 585
R554 B.n512 B.n511 585
R555 B.n510 B.n509 585
R556 B.n510 B.n8 585
R557 B.n508 B.n9 585
R558 B.n435 B.n9 585
R559 B.n507 B.n506 585
R560 B.n506 B.n505 585
R561 B.n11 B.n10 585
R562 B.n504 B.n11 585
R563 B.n502 B.n501 585
R564 B.n503 B.n502 585
R565 B.n500 B.n15 585
R566 B.n18 B.n15 585
R567 B.n499 B.n498 585
R568 B.n498 B.n497 585
R569 B.n17 B.n16 585
R570 B.n496 B.n17 585
R571 B.n494 B.n493 585
R572 B.n495 B.n494 585
R573 B.n492 B.n22 585
R574 B.n25 B.n22 585
R575 B.n491 B.n490 585
R576 B.n490 B.n489 585
R577 B.n24 B.n23 585
R578 B.n488 B.n24 585
R579 B.n486 B.n485 585
R580 B.n487 B.n486 585
R581 B.n484 B.n30 585
R582 B.n30 B.n29 585
R583 B.n483 B.n482 585
R584 B.n482 B.n481 585
R585 B.n32 B.n31 585
R586 B.n480 B.n32 585
R587 B.n478 B.n477 585
R588 B.n479 B.n478 585
R589 B.n476 B.n37 585
R590 B.n37 B.n36 585
R591 B.n475 B.n474 585
R592 B.n474 B.n473 585
R593 B.n39 B.n38 585
R594 B.n472 B.n39 585
R595 B.n470 B.n469 585
R596 B.n471 B.n470 585
R597 B.n468 B.n44 585
R598 B.n44 B.n43 585
R599 B.n515 B.n514 585
R600 B.n513 B.n2 585
R601 B.n466 B.n44 502.111
R602 B.n463 B.n73 502.111
R603 B.n254 B.n218 502.111
R604 B.n358 B.n220 502.111
R605 B.n76 B.t16 329.2
R606 B.n74 B.t5 329.2
R607 B.n251 B.t9 329.2
R608 B.n249 B.t13 329.2
R609 B.n464 B.n71 256.663
R610 B.n464 B.n70 256.663
R611 B.n464 B.n69 256.663
R612 B.n464 B.n68 256.663
R613 B.n464 B.n67 256.663
R614 B.n464 B.n66 256.663
R615 B.n464 B.n65 256.663
R616 B.n464 B.n64 256.663
R617 B.n464 B.n63 256.663
R618 B.n464 B.n62 256.663
R619 B.n464 B.n61 256.663
R620 B.n464 B.n60 256.663
R621 B.n464 B.n59 256.663
R622 B.n464 B.n58 256.663
R623 B.n464 B.n57 256.663
R624 B.n464 B.n56 256.663
R625 B.n464 B.n55 256.663
R626 B.n464 B.n54 256.663
R627 B.n464 B.n53 256.663
R628 B.n464 B.n52 256.663
R629 B.n464 B.n51 256.663
R630 B.n464 B.n50 256.663
R631 B.n464 B.n49 256.663
R632 B.n464 B.n48 256.663
R633 B.n464 B.n47 256.663
R634 B.n465 B.n464 256.663
R635 B.n357 B.n356 256.663
R636 B.n356 B.n223 256.663
R637 B.n356 B.n224 256.663
R638 B.n356 B.n225 256.663
R639 B.n356 B.n226 256.663
R640 B.n356 B.n227 256.663
R641 B.n356 B.n228 256.663
R642 B.n356 B.n229 256.663
R643 B.n356 B.n230 256.663
R644 B.n356 B.n231 256.663
R645 B.n356 B.n232 256.663
R646 B.n356 B.n233 256.663
R647 B.n356 B.n234 256.663
R648 B.n356 B.n235 256.663
R649 B.n356 B.n236 256.663
R650 B.n356 B.n237 256.663
R651 B.n356 B.n238 256.663
R652 B.n356 B.n239 256.663
R653 B.n356 B.n240 256.663
R654 B.n356 B.n241 256.663
R655 B.n356 B.n242 256.663
R656 B.n356 B.n243 256.663
R657 B.n356 B.n244 256.663
R658 B.n356 B.n245 256.663
R659 B.n356 B.n246 256.663
R660 B.n356 B.n247 256.663
R661 B.n517 B.n516 256.663
R662 B.n74 B.t7 190.429
R663 B.n251 B.t12 190.429
R664 B.n76 B.t17 190.429
R665 B.n249 B.t15 190.429
R666 B.n75 B.t8 164.828
R667 B.n252 B.t11 164.828
R668 B.n77 B.t18 164.828
R669 B.n250 B.t14 164.828
R670 B.n79 B.n46 163.367
R671 B.n83 B.n82 163.367
R672 B.n87 B.n86 163.367
R673 B.n91 B.n90 163.367
R674 B.n95 B.n94 163.367
R675 B.n99 B.n98 163.367
R676 B.n103 B.n102 163.367
R677 B.n107 B.n106 163.367
R678 B.n111 B.n110 163.367
R679 B.n115 B.n114 163.367
R680 B.n119 B.n118 163.367
R681 B.n123 B.n122 163.367
R682 B.n127 B.n126 163.367
R683 B.n131 B.n130 163.367
R684 B.n135 B.n134 163.367
R685 B.n140 B.n139 163.367
R686 B.n144 B.n143 163.367
R687 B.n148 B.n147 163.367
R688 B.n152 B.n151 163.367
R689 B.n156 B.n155 163.367
R690 B.n160 B.n159 163.367
R691 B.n164 B.n163 163.367
R692 B.n168 B.n167 163.367
R693 B.n172 B.n171 163.367
R694 B.n176 B.n175 163.367
R695 B.n463 B.n72 163.367
R696 B.n364 B.n218 163.367
R697 B.n364 B.n216 163.367
R698 B.n368 B.n216 163.367
R699 B.n368 B.n210 163.367
R700 B.n376 B.n210 163.367
R701 B.n376 B.n208 163.367
R702 B.n380 B.n208 163.367
R703 B.n380 B.n202 163.367
R704 B.n388 B.n202 163.367
R705 B.n388 B.n200 163.367
R706 B.n392 B.n200 163.367
R707 B.n392 B.n195 163.367
R708 B.n401 B.n195 163.367
R709 B.n401 B.n193 163.367
R710 B.n405 B.n193 163.367
R711 B.n405 B.n188 163.367
R712 B.n414 B.n188 163.367
R713 B.n414 B.n186 163.367
R714 B.n419 B.n186 163.367
R715 B.n419 B.n180 163.367
R716 B.n427 B.n180 163.367
R717 B.n428 B.n427 163.367
R718 B.n428 B.n5 163.367
R719 B.n6 B.n5 163.367
R720 B.n7 B.n6 163.367
R721 B.n434 B.n7 163.367
R722 B.n436 B.n434 163.367
R723 B.n436 B.n12 163.367
R724 B.n13 B.n12 163.367
R725 B.n14 B.n13 163.367
R726 B.n441 B.n14 163.367
R727 B.n441 B.n19 163.367
R728 B.n20 B.n19 163.367
R729 B.n21 B.n20 163.367
R730 B.n446 B.n21 163.367
R731 B.n446 B.n26 163.367
R732 B.n27 B.n26 163.367
R733 B.n28 B.n27 163.367
R734 B.n451 B.n28 163.367
R735 B.n451 B.n33 163.367
R736 B.n34 B.n33 163.367
R737 B.n35 B.n34 163.367
R738 B.n456 B.n35 163.367
R739 B.n456 B.n40 163.367
R740 B.n41 B.n40 163.367
R741 B.n42 B.n41 163.367
R742 B.n73 B.n42 163.367
R743 B.n355 B.n222 163.367
R744 B.n355 B.n248 163.367
R745 B.n351 B.n350 163.367
R746 B.n347 B.n346 163.367
R747 B.n343 B.n342 163.367
R748 B.n339 B.n338 163.367
R749 B.n335 B.n334 163.367
R750 B.n331 B.n330 163.367
R751 B.n327 B.n326 163.367
R752 B.n323 B.n322 163.367
R753 B.n319 B.n318 163.367
R754 B.n314 B.n313 163.367
R755 B.n310 B.n309 163.367
R756 B.n306 B.n305 163.367
R757 B.n302 B.n301 163.367
R758 B.n298 B.n297 163.367
R759 B.n294 B.n293 163.367
R760 B.n290 B.n289 163.367
R761 B.n286 B.n285 163.367
R762 B.n282 B.n281 163.367
R763 B.n278 B.n277 163.367
R764 B.n274 B.n273 163.367
R765 B.n270 B.n269 163.367
R766 B.n266 B.n265 163.367
R767 B.n262 B.n261 163.367
R768 B.n258 B.n257 163.367
R769 B.n362 B.n220 163.367
R770 B.n362 B.n214 163.367
R771 B.n370 B.n214 163.367
R772 B.n370 B.n212 163.367
R773 B.n374 B.n212 163.367
R774 B.n374 B.n206 163.367
R775 B.n382 B.n206 163.367
R776 B.n382 B.n204 163.367
R777 B.n386 B.n204 163.367
R778 B.n386 B.n198 163.367
R779 B.n395 B.n198 163.367
R780 B.n395 B.n196 163.367
R781 B.n399 B.n196 163.367
R782 B.n399 B.n191 163.367
R783 B.n408 B.n191 163.367
R784 B.n408 B.n189 163.367
R785 B.n412 B.n189 163.367
R786 B.n412 B.n184 163.367
R787 B.n421 B.n184 163.367
R788 B.n421 B.n182 163.367
R789 B.n425 B.n182 163.367
R790 B.n425 B.n3 163.367
R791 B.n515 B.n3 163.367
R792 B.n511 B.n2 163.367
R793 B.n511 B.n510 163.367
R794 B.n510 B.n9 163.367
R795 B.n506 B.n9 163.367
R796 B.n506 B.n11 163.367
R797 B.n502 B.n11 163.367
R798 B.n502 B.n15 163.367
R799 B.n498 B.n15 163.367
R800 B.n498 B.n17 163.367
R801 B.n494 B.n17 163.367
R802 B.n494 B.n22 163.367
R803 B.n490 B.n22 163.367
R804 B.n490 B.n24 163.367
R805 B.n486 B.n24 163.367
R806 B.n486 B.n30 163.367
R807 B.n482 B.n30 163.367
R808 B.n482 B.n32 163.367
R809 B.n478 B.n32 163.367
R810 B.n478 B.n37 163.367
R811 B.n474 B.n37 163.367
R812 B.n474 B.n39 163.367
R813 B.n470 B.n39 163.367
R814 B.n470 B.n44 163.367
R815 B.n356 B.n219 139.799
R816 B.n464 B.n43 139.799
R817 B.n466 B.n465 71.676
R818 B.n79 B.n47 71.676
R819 B.n83 B.n48 71.676
R820 B.n87 B.n49 71.676
R821 B.n91 B.n50 71.676
R822 B.n95 B.n51 71.676
R823 B.n99 B.n52 71.676
R824 B.n103 B.n53 71.676
R825 B.n107 B.n54 71.676
R826 B.n111 B.n55 71.676
R827 B.n115 B.n56 71.676
R828 B.n119 B.n57 71.676
R829 B.n123 B.n58 71.676
R830 B.n127 B.n59 71.676
R831 B.n131 B.n60 71.676
R832 B.n135 B.n61 71.676
R833 B.n140 B.n62 71.676
R834 B.n144 B.n63 71.676
R835 B.n148 B.n64 71.676
R836 B.n152 B.n65 71.676
R837 B.n156 B.n66 71.676
R838 B.n160 B.n67 71.676
R839 B.n164 B.n68 71.676
R840 B.n168 B.n69 71.676
R841 B.n172 B.n70 71.676
R842 B.n176 B.n71 71.676
R843 B.n72 B.n71 71.676
R844 B.n175 B.n70 71.676
R845 B.n171 B.n69 71.676
R846 B.n167 B.n68 71.676
R847 B.n163 B.n67 71.676
R848 B.n159 B.n66 71.676
R849 B.n155 B.n65 71.676
R850 B.n151 B.n64 71.676
R851 B.n147 B.n63 71.676
R852 B.n143 B.n62 71.676
R853 B.n139 B.n61 71.676
R854 B.n134 B.n60 71.676
R855 B.n130 B.n59 71.676
R856 B.n126 B.n58 71.676
R857 B.n122 B.n57 71.676
R858 B.n118 B.n56 71.676
R859 B.n114 B.n55 71.676
R860 B.n110 B.n54 71.676
R861 B.n106 B.n53 71.676
R862 B.n102 B.n52 71.676
R863 B.n98 B.n51 71.676
R864 B.n94 B.n50 71.676
R865 B.n90 B.n49 71.676
R866 B.n86 B.n48 71.676
R867 B.n82 B.n47 71.676
R868 B.n465 B.n46 71.676
R869 B.n358 B.n357 71.676
R870 B.n248 B.n223 71.676
R871 B.n350 B.n224 71.676
R872 B.n346 B.n225 71.676
R873 B.n342 B.n226 71.676
R874 B.n338 B.n227 71.676
R875 B.n334 B.n228 71.676
R876 B.n330 B.n229 71.676
R877 B.n326 B.n230 71.676
R878 B.n322 B.n231 71.676
R879 B.n318 B.n232 71.676
R880 B.n313 B.n233 71.676
R881 B.n309 B.n234 71.676
R882 B.n305 B.n235 71.676
R883 B.n301 B.n236 71.676
R884 B.n297 B.n237 71.676
R885 B.n293 B.n238 71.676
R886 B.n289 B.n239 71.676
R887 B.n285 B.n240 71.676
R888 B.n281 B.n241 71.676
R889 B.n277 B.n242 71.676
R890 B.n273 B.n243 71.676
R891 B.n269 B.n244 71.676
R892 B.n265 B.n245 71.676
R893 B.n261 B.n246 71.676
R894 B.n257 B.n247 71.676
R895 B.n357 B.n222 71.676
R896 B.n351 B.n223 71.676
R897 B.n347 B.n224 71.676
R898 B.n343 B.n225 71.676
R899 B.n339 B.n226 71.676
R900 B.n335 B.n227 71.676
R901 B.n331 B.n228 71.676
R902 B.n327 B.n229 71.676
R903 B.n323 B.n230 71.676
R904 B.n319 B.n231 71.676
R905 B.n314 B.n232 71.676
R906 B.n310 B.n233 71.676
R907 B.n306 B.n234 71.676
R908 B.n302 B.n235 71.676
R909 B.n298 B.n236 71.676
R910 B.n294 B.n237 71.676
R911 B.n290 B.n238 71.676
R912 B.n286 B.n239 71.676
R913 B.n282 B.n240 71.676
R914 B.n278 B.n241 71.676
R915 B.n274 B.n242 71.676
R916 B.n270 B.n243 71.676
R917 B.n266 B.n244 71.676
R918 B.n262 B.n245 71.676
R919 B.n258 B.n246 71.676
R920 B.n254 B.n247 71.676
R921 B.n516 B.n515 71.676
R922 B.n516 B.n2 71.676
R923 B.n363 B.n219 71.4768
R924 B.n363 B.n215 71.4768
R925 B.n369 B.n215 71.4768
R926 B.n369 B.n211 71.4768
R927 B.n375 B.n211 71.4768
R928 B.n381 B.n207 71.4768
R929 B.n381 B.n203 71.4768
R930 B.n387 B.n203 71.4768
R931 B.n387 B.n199 71.4768
R932 B.n394 B.n199 71.4768
R933 B.n394 B.n393 71.4768
R934 B.n400 B.n192 71.4768
R935 B.n407 B.n192 71.4768
R936 B.n407 B.n406 71.4768
R937 B.n413 B.n185 71.4768
R938 B.n420 B.n185 71.4768
R939 B.n426 B.n181 71.4768
R940 B.n426 B.n4 71.4768
R941 B.n514 B.n4 71.4768
R942 B.n514 B.n513 71.4768
R943 B.n513 B.n512 71.4768
R944 B.n512 B.n8 71.4768
R945 B.n435 B.n8 71.4768
R946 B.n505 B.n504 71.4768
R947 B.n504 B.n503 71.4768
R948 B.n497 B.n18 71.4768
R949 B.n497 B.n496 71.4768
R950 B.n496 B.n495 71.4768
R951 B.n489 B.n25 71.4768
R952 B.n489 B.n488 71.4768
R953 B.n488 B.n487 71.4768
R954 B.n487 B.n29 71.4768
R955 B.n481 B.n29 71.4768
R956 B.n481 B.n480 71.4768
R957 B.n479 B.n36 71.4768
R958 B.n473 B.n36 71.4768
R959 B.n473 B.n472 71.4768
R960 B.n472 B.n471 71.4768
R961 B.n471 B.n43 71.4768
R962 B.n420 B.t0 68.3235
R963 B.n505 B.t4 68.3235
R964 B.n413 B.t3 66.2212
R965 B.n503 B.t1 66.2212
R966 B.t10 B.n207 64.119
R967 B.n480 B.t6 64.119
R968 B.n78 B.n77 59.5399
R969 B.n137 B.n75 59.5399
R970 B.n253 B.n252 59.5399
R971 B.n316 B.n250 59.5399
R972 B.n400 B.t19 57.8123
R973 B.n495 B.t2 57.8123
R974 B.n360 B.n359 32.6249
R975 B.n255 B.n217 32.6249
R976 B.n462 B.n461 32.6249
R977 B.n468 B.n467 32.6249
R978 B.n77 B.n76 25.6005
R979 B.n75 B.n74 25.6005
R980 B.n252 B.n251 25.6005
R981 B.n250 B.n249 25.6005
R982 B B.n517 18.0485
R983 B.n393 B.t19 13.6651
R984 B.n25 B.t2 13.6651
R985 B.n361 B.n360 10.6151
R986 B.n361 B.n213 10.6151
R987 B.n371 B.n213 10.6151
R988 B.n372 B.n371 10.6151
R989 B.n373 B.n372 10.6151
R990 B.n373 B.n205 10.6151
R991 B.n383 B.n205 10.6151
R992 B.n384 B.n383 10.6151
R993 B.n385 B.n384 10.6151
R994 B.n385 B.n197 10.6151
R995 B.n396 B.n197 10.6151
R996 B.n397 B.n396 10.6151
R997 B.n398 B.n397 10.6151
R998 B.n398 B.n190 10.6151
R999 B.n409 B.n190 10.6151
R1000 B.n410 B.n409 10.6151
R1001 B.n411 B.n410 10.6151
R1002 B.n411 B.n183 10.6151
R1003 B.n422 B.n183 10.6151
R1004 B.n423 B.n422 10.6151
R1005 B.n424 B.n423 10.6151
R1006 B.n424 B.n0 10.6151
R1007 B.n359 B.n221 10.6151
R1008 B.n354 B.n221 10.6151
R1009 B.n354 B.n353 10.6151
R1010 B.n353 B.n352 10.6151
R1011 B.n352 B.n349 10.6151
R1012 B.n349 B.n348 10.6151
R1013 B.n348 B.n345 10.6151
R1014 B.n345 B.n344 10.6151
R1015 B.n344 B.n341 10.6151
R1016 B.n341 B.n340 10.6151
R1017 B.n340 B.n337 10.6151
R1018 B.n337 B.n336 10.6151
R1019 B.n336 B.n333 10.6151
R1020 B.n333 B.n332 10.6151
R1021 B.n332 B.n329 10.6151
R1022 B.n329 B.n328 10.6151
R1023 B.n328 B.n325 10.6151
R1024 B.n325 B.n324 10.6151
R1025 B.n324 B.n321 10.6151
R1026 B.n321 B.n320 10.6151
R1027 B.n320 B.n317 10.6151
R1028 B.n315 B.n312 10.6151
R1029 B.n312 B.n311 10.6151
R1030 B.n311 B.n308 10.6151
R1031 B.n308 B.n307 10.6151
R1032 B.n307 B.n304 10.6151
R1033 B.n304 B.n303 10.6151
R1034 B.n303 B.n300 10.6151
R1035 B.n300 B.n299 10.6151
R1036 B.n296 B.n295 10.6151
R1037 B.n295 B.n292 10.6151
R1038 B.n292 B.n291 10.6151
R1039 B.n291 B.n288 10.6151
R1040 B.n288 B.n287 10.6151
R1041 B.n287 B.n284 10.6151
R1042 B.n284 B.n283 10.6151
R1043 B.n283 B.n280 10.6151
R1044 B.n280 B.n279 10.6151
R1045 B.n279 B.n276 10.6151
R1046 B.n276 B.n275 10.6151
R1047 B.n275 B.n272 10.6151
R1048 B.n272 B.n271 10.6151
R1049 B.n271 B.n268 10.6151
R1050 B.n268 B.n267 10.6151
R1051 B.n267 B.n264 10.6151
R1052 B.n264 B.n263 10.6151
R1053 B.n263 B.n260 10.6151
R1054 B.n260 B.n259 10.6151
R1055 B.n259 B.n256 10.6151
R1056 B.n256 B.n255 10.6151
R1057 B.n365 B.n217 10.6151
R1058 B.n366 B.n365 10.6151
R1059 B.n367 B.n366 10.6151
R1060 B.n367 B.n209 10.6151
R1061 B.n377 B.n209 10.6151
R1062 B.n378 B.n377 10.6151
R1063 B.n379 B.n378 10.6151
R1064 B.n379 B.n201 10.6151
R1065 B.n389 B.n201 10.6151
R1066 B.n390 B.n389 10.6151
R1067 B.n391 B.n390 10.6151
R1068 B.n391 B.n194 10.6151
R1069 B.n402 B.n194 10.6151
R1070 B.n403 B.n402 10.6151
R1071 B.n404 B.n403 10.6151
R1072 B.n404 B.n187 10.6151
R1073 B.n415 B.n187 10.6151
R1074 B.n416 B.n415 10.6151
R1075 B.n418 B.n416 10.6151
R1076 B.n418 B.n417 10.6151
R1077 B.n417 B.n179 10.6151
R1078 B.n429 B.n179 10.6151
R1079 B.n430 B.n429 10.6151
R1080 B.n431 B.n430 10.6151
R1081 B.n432 B.n431 10.6151
R1082 B.n433 B.n432 10.6151
R1083 B.n437 B.n433 10.6151
R1084 B.n438 B.n437 10.6151
R1085 B.n439 B.n438 10.6151
R1086 B.n440 B.n439 10.6151
R1087 B.n442 B.n440 10.6151
R1088 B.n443 B.n442 10.6151
R1089 B.n444 B.n443 10.6151
R1090 B.n445 B.n444 10.6151
R1091 B.n447 B.n445 10.6151
R1092 B.n448 B.n447 10.6151
R1093 B.n449 B.n448 10.6151
R1094 B.n450 B.n449 10.6151
R1095 B.n452 B.n450 10.6151
R1096 B.n453 B.n452 10.6151
R1097 B.n454 B.n453 10.6151
R1098 B.n455 B.n454 10.6151
R1099 B.n457 B.n455 10.6151
R1100 B.n458 B.n457 10.6151
R1101 B.n459 B.n458 10.6151
R1102 B.n460 B.n459 10.6151
R1103 B.n461 B.n460 10.6151
R1104 B.n509 B.n1 10.6151
R1105 B.n509 B.n508 10.6151
R1106 B.n508 B.n507 10.6151
R1107 B.n507 B.n10 10.6151
R1108 B.n501 B.n10 10.6151
R1109 B.n501 B.n500 10.6151
R1110 B.n500 B.n499 10.6151
R1111 B.n499 B.n16 10.6151
R1112 B.n493 B.n16 10.6151
R1113 B.n493 B.n492 10.6151
R1114 B.n492 B.n491 10.6151
R1115 B.n491 B.n23 10.6151
R1116 B.n485 B.n23 10.6151
R1117 B.n485 B.n484 10.6151
R1118 B.n484 B.n483 10.6151
R1119 B.n483 B.n31 10.6151
R1120 B.n477 B.n31 10.6151
R1121 B.n477 B.n476 10.6151
R1122 B.n476 B.n475 10.6151
R1123 B.n475 B.n38 10.6151
R1124 B.n469 B.n38 10.6151
R1125 B.n469 B.n468 10.6151
R1126 B.n467 B.n45 10.6151
R1127 B.n80 B.n45 10.6151
R1128 B.n81 B.n80 10.6151
R1129 B.n84 B.n81 10.6151
R1130 B.n85 B.n84 10.6151
R1131 B.n88 B.n85 10.6151
R1132 B.n89 B.n88 10.6151
R1133 B.n92 B.n89 10.6151
R1134 B.n93 B.n92 10.6151
R1135 B.n96 B.n93 10.6151
R1136 B.n97 B.n96 10.6151
R1137 B.n100 B.n97 10.6151
R1138 B.n101 B.n100 10.6151
R1139 B.n104 B.n101 10.6151
R1140 B.n105 B.n104 10.6151
R1141 B.n108 B.n105 10.6151
R1142 B.n109 B.n108 10.6151
R1143 B.n112 B.n109 10.6151
R1144 B.n113 B.n112 10.6151
R1145 B.n116 B.n113 10.6151
R1146 B.n117 B.n116 10.6151
R1147 B.n121 B.n120 10.6151
R1148 B.n124 B.n121 10.6151
R1149 B.n125 B.n124 10.6151
R1150 B.n128 B.n125 10.6151
R1151 B.n129 B.n128 10.6151
R1152 B.n132 B.n129 10.6151
R1153 B.n133 B.n132 10.6151
R1154 B.n136 B.n133 10.6151
R1155 B.n141 B.n138 10.6151
R1156 B.n142 B.n141 10.6151
R1157 B.n145 B.n142 10.6151
R1158 B.n146 B.n145 10.6151
R1159 B.n149 B.n146 10.6151
R1160 B.n150 B.n149 10.6151
R1161 B.n153 B.n150 10.6151
R1162 B.n154 B.n153 10.6151
R1163 B.n157 B.n154 10.6151
R1164 B.n158 B.n157 10.6151
R1165 B.n161 B.n158 10.6151
R1166 B.n162 B.n161 10.6151
R1167 B.n165 B.n162 10.6151
R1168 B.n166 B.n165 10.6151
R1169 B.n169 B.n166 10.6151
R1170 B.n170 B.n169 10.6151
R1171 B.n173 B.n170 10.6151
R1172 B.n174 B.n173 10.6151
R1173 B.n177 B.n174 10.6151
R1174 B.n178 B.n177 10.6151
R1175 B.n462 B.n178 10.6151
R1176 B.n517 B.n0 8.11757
R1177 B.n517 B.n1 8.11757
R1178 B.n375 B.t10 7.35836
R1179 B.t6 B.n479 7.35836
R1180 B.n316 B.n315 6.5566
R1181 B.n299 B.n253 6.5566
R1182 B.n120 B.n78 6.5566
R1183 B.n137 B.n136 6.5566
R1184 B.n406 B.t3 5.25611
R1185 B.n18 B.t1 5.25611
R1186 B.n317 B.n316 4.05904
R1187 B.n296 B.n253 4.05904
R1188 B.n117 B.n78 4.05904
R1189 B.n138 B.n137 4.05904
R1190 B.t0 B.n181 3.15387
R1191 B.n435 B.t4 3.15387
R1192 VP.n3 VP.t3 188.536
R1193 VP.n8 VP.t1 166.267
R1194 VP.n14 VP.t5 166.267
R1195 VP.n6 VP.t4 166.267
R1196 VP.n5 VP.n2 161.3
R1197 VP.n13 VP.n0 161.3
R1198 VP.n12 VP.n11 161.3
R1199 VP.n10 VP.n1 161.3
R1200 VP.n12 VP.t2 126.343
R1201 VP.n4 VP.t0 126.343
R1202 VP.n7 VP.n6 80.6037
R1203 VP.n15 VP.n14 80.6037
R1204 VP.n9 VP.n8 80.6037
R1205 VP.n8 VP.n1 47.4702
R1206 VP.n14 VP.n13 47.4702
R1207 VP.n6 VP.n5 47.4702
R1208 VP.n9 VP.n7 37.2817
R1209 VP.n4 VP.n3 32.1379
R1210 VP.n3 VP.n2 28.4787
R1211 VP.n12 VP.n1 24.9531
R1212 VP.n13 VP.n12 24.9531
R1213 VP.n5 VP.n4 24.9531
R1214 VP.n7 VP.n2 0.285035
R1215 VP.n10 VP.n9 0.285035
R1216 VP.n15 VP.n0 0.285035
R1217 VP.n11 VP.n10 0.189894
R1218 VP.n11 VP.n0 0.189894
R1219 VP VP.n15 0.146778
R1220 VDD1.n22 VDD1.n0 289.615
R1221 VDD1.n49 VDD1.n27 289.615
R1222 VDD1.n23 VDD1.n22 185
R1223 VDD1.n21 VDD1.n20 185
R1224 VDD1.n4 VDD1.n3 185
R1225 VDD1.n15 VDD1.n14 185
R1226 VDD1.n13 VDD1.n12 185
R1227 VDD1.n8 VDD1.n7 185
R1228 VDD1.n35 VDD1.n34 185
R1229 VDD1.n40 VDD1.n39 185
R1230 VDD1.n42 VDD1.n41 185
R1231 VDD1.n31 VDD1.n30 185
R1232 VDD1.n48 VDD1.n47 185
R1233 VDD1.n50 VDD1.n49 185
R1234 VDD1.n9 VDD1.t2 147.672
R1235 VDD1.n36 VDD1.t4 147.672
R1236 VDD1.n22 VDD1.n21 104.615
R1237 VDD1.n21 VDD1.n3 104.615
R1238 VDD1.n14 VDD1.n3 104.615
R1239 VDD1.n14 VDD1.n13 104.615
R1240 VDD1.n13 VDD1.n7 104.615
R1241 VDD1.n40 VDD1.n34 104.615
R1242 VDD1.n41 VDD1.n40 104.615
R1243 VDD1.n41 VDD1.n30 104.615
R1244 VDD1.n48 VDD1.n30 104.615
R1245 VDD1.n49 VDD1.n48 104.615
R1246 VDD1.n55 VDD1.n54 67.1388
R1247 VDD1.n57 VDD1.n56 66.9097
R1248 VDD1.t2 VDD1.n7 52.3082
R1249 VDD1.t4 VDD1.n34 52.3082
R1250 VDD1 VDD1.n26 48.0303
R1251 VDD1.n55 VDD1.n53 47.9168
R1252 VDD1.n57 VDD1.n55 33.0397
R1253 VDD1.n9 VDD1.n8 15.6666
R1254 VDD1.n36 VDD1.n35 15.6666
R1255 VDD1.n12 VDD1.n11 12.8005
R1256 VDD1.n39 VDD1.n38 12.8005
R1257 VDD1.n15 VDD1.n6 12.0247
R1258 VDD1.n42 VDD1.n33 12.0247
R1259 VDD1.n16 VDD1.n4 11.249
R1260 VDD1.n43 VDD1.n31 11.249
R1261 VDD1.n20 VDD1.n19 10.4732
R1262 VDD1.n47 VDD1.n46 10.4732
R1263 VDD1.n23 VDD1.n2 9.69747
R1264 VDD1.n50 VDD1.n29 9.69747
R1265 VDD1.n26 VDD1.n25 9.45567
R1266 VDD1.n53 VDD1.n52 9.45567
R1267 VDD1.n25 VDD1.n24 9.3005
R1268 VDD1.n2 VDD1.n1 9.3005
R1269 VDD1.n19 VDD1.n18 9.3005
R1270 VDD1.n17 VDD1.n16 9.3005
R1271 VDD1.n6 VDD1.n5 9.3005
R1272 VDD1.n11 VDD1.n10 9.3005
R1273 VDD1.n52 VDD1.n51 9.3005
R1274 VDD1.n29 VDD1.n28 9.3005
R1275 VDD1.n46 VDD1.n45 9.3005
R1276 VDD1.n44 VDD1.n43 9.3005
R1277 VDD1.n33 VDD1.n32 9.3005
R1278 VDD1.n38 VDD1.n37 9.3005
R1279 VDD1.n24 VDD1.n0 8.92171
R1280 VDD1.n51 VDD1.n27 8.92171
R1281 VDD1.n26 VDD1.n0 5.04292
R1282 VDD1.n53 VDD1.n27 5.04292
R1283 VDD1.n10 VDD1.n9 4.38687
R1284 VDD1.n37 VDD1.n36 4.38687
R1285 VDD1.n24 VDD1.n23 4.26717
R1286 VDD1.n51 VDD1.n50 4.26717
R1287 VDD1.n56 VDD1.t5 3.81553
R1288 VDD1.n56 VDD1.t1 3.81553
R1289 VDD1.n54 VDD1.t3 3.81553
R1290 VDD1.n54 VDD1.t0 3.81553
R1291 VDD1.n20 VDD1.n2 3.49141
R1292 VDD1.n47 VDD1.n29 3.49141
R1293 VDD1.n19 VDD1.n4 2.71565
R1294 VDD1.n46 VDD1.n31 2.71565
R1295 VDD1.n16 VDD1.n15 1.93989
R1296 VDD1.n43 VDD1.n42 1.93989
R1297 VDD1.n12 VDD1.n6 1.16414
R1298 VDD1.n39 VDD1.n33 1.16414
R1299 VDD1.n11 VDD1.n8 0.388379
R1300 VDD1.n38 VDD1.n35 0.388379
R1301 VDD1 VDD1.n57 0.226793
R1302 VDD1.n25 VDD1.n1 0.155672
R1303 VDD1.n18 VDD1.n1 0.155672
R1304 VDD1.n18 VDD1.n17 0.155672
R1305 VDD1.n17 VDD1.n5 0.155672
R1306 VDD1.n10 VDD1.n5 0.155672
R1307 VDD1.n37 VDD1.n32 0.155672
R1308 VDD1.n44 VDD1.n32 0.155672
R1309 VDD1.n45 VDD1.n44 0.155672
R1310 VDD1.n45 VDD1.n28 0.155672
R1311 VDD1.n52 VDD1.n28 0.155672
C0 VN VP 4.10501f
C1 VDD2 VDD1 0.815425f
C2 VDD2 VTAIL 5.04988f
C3 VDD1 VP 2.55924f
C4 VDD1 VN 0.148581f
C5 VTAIL VP 2.51809f
C6 VN VTAIL 2.50381f
C7 VDD1 VTAIL 5.00961f
C8 VDD2 VP 0.325217f
C9 VDD2 VN 2.38872f
C10 VDD2 B 3.486715f
C11 VDD1 B 3.534708f
C12 VTAIL B 3.927194f
C13 VN B 7.65202f
C14 VP B 6.106374f
C15 VDD1.n0 B 0.030142f
C16 VDD1.n1 B 0.022871f
C17 VDD1.n2 B 0.01229f
C18 VDD1.n3 B 0.029049f
C19 VDD1.n4 B 0.013013f
C20 VDD1.n5 B 0.022871f
C21 VDD1.n6 B 0.01229f
C22 VDD1.n7 B 0.021787f
C23 VDD1.n8 B 0.017156f
C24 VDD1.t2 B 0.047363f
C25 VDD1.n9 B 0.09337f
C26 VDD1.n10 B 0.459083f
C27 VDD1.n11 B 0.01229f
C28 VDD1.n12 B 0.013013f
C29 VDD1.n13 B 0.029049f
C30 VDD1.n14 B 0.029049f
C31 VDD1.n15 B 0.013013f
C32 VDD1.n16 B 0.01229f
C33 VDD1.n17 B 0.022871f
C34 VDD1.n18 B 0.022871f
C35 VDD1.n19 B 0.01229f
C36 VDD1.n20 B 0.013013f
C37 VDD1.n21 B 0.029049f
C38 VDD1.n22 B 0.05934f
C39 VDD1.n23 B 0.013013f
C40 VDD1.n24 B 0.01229f
C41 VDD1.n25 B 0.050054f
C42 VDD1.n26 B 0.050646f
C43 VDD1.n27 B 0.030142f
C44 VDD1.n28 B 0.022871f
C45 VDD1.n29 B 0.01229f
C46 VDD1.n30 B 0.029049f
C47 VDD1.n31 B 0.013013f
C48 VDD1.n32 B 0.022871f
C49 VDD1.n33 B 0.01229f
C50 VDD1.n34 B 0.021787f
C51 VDD1.n35 B 0.017156f
C52 VDD1.t4 B 0.047363f
C53 VDD1.n36 B 0.09337f
C54 VDD1.n37 B 0.459083f
C55 VDD1.n38 B 0.01229f
C56 VDD1.n39 B 0.013013f
C57 VDD1.n40 B 0.029049f
C58 VDD1.n41 B 0.029049f
C59 VDD1.n42 B 0.013013f
C60 VDD1.n43 B 0.01229f
C61 VDD1.n44 B 0.022871f
C62 VDD1.n45 B 0.022871f
C63 VDD1.n46 B 0.01229f
C64 VDD1.n47 B 0.013013f
C65 VDD1.n48 B 0.029049f
C66 VDD1.n49 B 0.05934f
C67 VDD1.n50 B 0.013013f
C68 VDD1.n51 B 0.01229f
C69 VDD1.n52 B 0.050054f
C70 VDD1.n53 B 0.050263f
C71 VDD1.t3 B 0.093803f
C72 VDD1.t0 B 0.093803f
C73 VDD1.n54 B 0.768497f
C74 VDD1.n55 B 1.50761f
C75 VDD1.t5 B 0.093803f
C76 VDD1.t1 B 0.093803f
C77 VDD1.n56 B 0.767488f
C78 VDD1.n57 B 1.63932f
C79 VP.n0 B 0.05762f
C80 VP.t2 B 0.581848f
C81 VP.n1 B 0.04811f
C82 VP.n2 B 0.231819f
C83 VP.t4 B 0.647341f
C84 VP.t0 B 0.581848f
C85 VP.t3 B 0.685107f
C86 VP.n3 B 0.297372f
C87 VP.n4 B 0.314001f
C88 VP.n5 B 0.04811f
C89 VP.n6 B 0.309789f
C90 VP.n7 B 1.46379f
C91 VP.t1 B 0.647341f
C92 VP.n8 B 0.309789f
C93 VP.n9 B 1.50543f
C94 VP.n10 B 0.05762f
C95 VP.n11 B 0.043181f
C96 VP.n12 B 0.289252f
C97 VP.n13 B 0.04811f
C98 VP.t5 B 0.647341f
C99 VP.n14 B 0.309789f
C100 VP.n15 B 0.040441f
C101 VDD2.n0 B 0.029678f
C102 VDD2.n1 B 0.02252f
C103 VDD2.n2 B 0.012101f
C104 VDD2.n3 B 0.028603f
C105 VDD2.n4 B 0.012813f
C106 VDD2.n5 B 0.02252f
C107 VDD2.n6 B 0.012101f
C108 VDD2.n7 B 0.021452f
C109 VDD2.n8 B 0.016892f
C110 VDD2.t0 B 0.046635f
C111 VDD2.n9 B 0.091935f
C112 VDD2.n10 B 0.452026f
C113 VDD2.n11 B 0.012101f
C114 VDD2.n12 B 0.012813f
C115 VDD2.n13 B 0.028603f
C116 VDD2.n14 B 0.028603f
C117 VDD2.n15 B 0.012813f
C118 VDD2.n16 B 0.012101f
C119 VDD2.n17 B 0.02252f
C120 VDD2.n18 B 0.02252f
C121 VDD2.n19 B 0.012101f
C122 VDD2.n20 B 0.012813f
C123 VDD2.n21 B 0.028603f
C124 VDD2.n22 B 0.058427f
C125 VDD2.n23 B 0.012813f
C126 VDD2.n24 B 0.012101f
C127 VDD2.n25 B 0.049285f
C128 VDD2.n26 B 0.049491f
C129 VDD2.t4 B 0.092361f
C130 VDD2.t3 B 0.092361f
C131 VDD2.n27 B 0.756684f
C132 VDD2.n28 B 1.41216f
C133 VDD2.n29 B 0.029678f
C134 VDD2.n30 B 0.02252f
C135 VDD2.n31 B 0.012101f
C136 VDD2.n32 B 0.028603f
C137 VDD2.n33 B 0.012813f
C138 VDD2.n34 B 0.02252f
C139 VDD2.n35 B 0.012101f
C140 VDD2.n36 B 0.021452f
C141 VDD2.n37 B 0.016892f
C142 VDD2.t5 B 0.046635f
C143 VDD2.n38 B 0.091935f
C144 VDD2.n39 B 0.452026f
C145 VDD2.n40 B 0.012101f
C146 VDD2.n41 B 0.012813f
C147 VDD2.n42 B 0.028603f
C148 VDD2.n43 B 0.028603f
C149 VDD2.n44 B 0.012813f
C150 VDD2.n45 B 0.012101f
C151 VDD2.n46 B 0.02252f
C152 VDD2.n47 B 0.02252f
C153 VDD2.n48 B 0.012101f
C154 VDD2.n49 B 0.012813f
C155 VDD2.n50 B 0.028603f
C156 VDD2.n51 B 0.058427f
C157 VDD2.n52 B 0.012813f
C158 VDD2.n53 B 0.012101f
C159 VDD2.n54 B 0.049285f
C160 VDD2.n55 B 0.047819f
C161 VDD2.n56 B 1.42264f
C162 VDD2.t2 B 0.092361f
C163 VDD2.t1 B 0.092361f
C164 VDD2.n57 B 0.756663f
C165 VTAIL.t9 B 0.106813f
C166 VTAIL.t5 B 0.106813f
C167 VTAIL.n0 B 0.806295f
C168 VTAIL.n1 B 0.356849f
C169 VTAIL.n2 B 0.034323f
C170 VTAIL.n3 B 0.026044f
C171 VTAIL.n4 B 0.013995f
C172 VTAIL.n5 B 0.033078f
C173 VTAIL.n6 B 0.014818f
C174 VTAIL.n7 B 0.026044f
C175 VTAIL.n8 B 0.013995f
C176 VTAIL.n9 B 0.024809f
C177 VTAIL.n10 B 0.019535f
C178 VTAIL.t0 B 0.053932f
C179 VTAIL.n11 B 0.106321f
C180 VTAIL.n12 B 0.522757f
C181 VTAIL.n13 B 0.013995f
C182 VTAIL.n14 B 0.014818f
C183 VTAIL.n15 B 0.033078f
C184 VTAIL.n16 B 0.033078f
C185 VTAIL.n17 B 0.014818f
C186 VTAIL.n18 B 0.013995f
C187 VTAIL.n19 B 0.026044f
C188 VTAIL.n20 B 0.026044f
C189 VTAIL.n21 B 0.013995f
C190 VTAIL.n22 B 0.014818f
C191 VTAIL.n23 B 0.033078f
C192 VTAIL.n24 B 0.06757f
C193 VTAIL.n25 B 0.014818f
C194 VTAIL.n26 B 0.013995f
C195 VTAIL.n27 B 0.056997f
C196 VTAIL.n28 B 0.037292f
C197 VTAIL.n29 B 0.203106f
C198 VTAIL.t11 B 0.106813f
C199 VTAIL.t3 B 0.106813f
C200 VTAIL.n30 B 0.806295f
C201 VTAIL.n31 B 1.25664f
C202 VTAIL.t8 B 0.106813f
C203 VTAIL.t7 B 0.106813f
C204 VTAIL.n32 B 0.806301f
C205 VTAIL.n33 B 1.25663f
C206 VTAIL.n34 B 0.034323f
C207 VTAIL.n35 B 0.026044f
C208 VTAIL.n36 B 0.013995f
C209 VTAIL.n37 B 0.033078f
C210 VTAIL.n38 B 0.014818f
C211 VTAIL.n39 B 0.026044f
C212 VTAIL.n40 B 0.013995f
C213 VTAIL.n41 B 0.024809f
C214 VTAIL.n42 B 0.019535f
C215 VTAIL.t6 B 0.053932f
C216 VTAIL.n43 B 0.106321f
C217 VTAIL.n44 B 0.522757f
C218 VTAIL.n45 B 0.013995f
C219 VTAIL.n46 B 0.014818f
C220 VTAIL.n47 B 0.033078f
C221 VTAIL.n48 B 0.033078f
C222 VTAIL.n49 B 0.014818f
C223 VTAIL.n50 B 0.013995f
C224 VTAIL.n51 B 0.026044f
C225 VTAIL.n52 B 0.026044f
C226 VTAIL.n53 B 0.013995f
C227 VTAIL.n54 B 0.014818f
C228 VTAIL.n55 B 0.033078f
C229 VTAIL.n56 B 0.06757f
C230 VTAIL.n57 B 0.014818f
C231 VTAIL.n58 B 0.013995f
C232 VTAIL.n59 B 0.056997f
C233 VTAIL.n60 B 0.037292f
C234 VTAIL.n61 B 0.203106f
C235 VTAIL.t4 B 0.106813f
C236 VTAIL.t1 B 0.106813f
C237 VTAIL.n62 B 0.806301f
C238 VTAIL.n63 B 0.42358f
C239 VTAIL.n64 B 0.034323f
C240 VTAIL.n65 B 0.026044f
C241 VTAIL.n66 B 0.013995f
C242 VTAIL.n67 B 0.033078f
C243 VTAIL.n68 B 0.014818f
C244 VTAIL.n69 B 0.026044f
C245 VTAIL.n70 B 0.013995f
C246 VTAIL.n71 B 0.024809f
C247 VTAIL.n72 B 0.019535f
C248 VTAIL.t2 B 0.053932f
C249 VTAIL.n73 B 0.106321f
C250 VTAIL.n74 B 0.522757f
C251 VTAIL.n75 B 0.013995f
C252 VTAIL.n76 B 0.014818f
C253 VTAIL.n77 B 0.033078f
C254 VTAIL.n78 B 0.033078f
C255 VTAIL.n79 B 0.014818f
C256 VTAIL.n80 B 0.013995f
C257 VTAIL.n81 B 0.026044f
C258 VTAIL.n82 B 0.026044f
C259 VTAIL.n83 B 0.013995f
C260 VTAIL.n84 B 0.014818f
C261 VTAIL.n85 B 0.033078f
C262 VTAIL.n86 B 0.06757f
C263 VTAIL.n87 B 0.014818f
C264 VTAIL.n88 B 0.013995f
C265 VTAIL.n89 B 0.056997f
C266 VTAIL.n90 B 0.037292f
C267 VTAIL.n91 B 0.940663f
C268 VTAIL.n92 B 0.034323f
C269 VTAIL.n93 B 0.026044f
C270 VTAIL.n94 B 0.013995f
C271 VTAIL.n95 B 0.033078f
C272 VTAIL.n96 B 0.014818f
C273 VTAIL.n97 B 0.026044f
C274 VTAIL.n98 B 0.013995f
C275 VTAIL.n99 B 0.024809f
C276 VTAIL.n100 B 0.019535f
C277 VTAIL.t10 B 0.053932f
C278 VTAIL.n101 B 0.106321f
C279 VTAIL.n102 B 0.522757f
C280 VTAIL.n103 B 0.013995f
C281 VTAIL.n104 B 0.014818f
C282 VTAIL.n105 B 0.033078f
C283 VTAIL.n106 B 0.033078f
C284 VTAIL.n107 B 0.014818f
C285 VTAIL.n108 B 0.013995f
C286 VTAIL.n109 B 0.026044f
C287 VTAIL.n110 B 0.026044f
C288 VTAIL.n111 B 0.013995f
C289 VTAIL.n112 B 0.014818f
C290 VTAIL.n113 B 0.033078f
C291 VTAIL.n114 B 0.06757f
C292 VTAIL.n115 B 0.014818f
C293 VTAIL.n116 B 0.013995f
C294 VTAIL.n117 B 0.056997f
C295 VTAIL.n118 B 0.037292f
C296 VTAIL.n119 B 0.911907f
C297 VN.n0 B 0.225293f
C298 VN.t1 B 0.565469f
C299 VN.t5 B 0.665821f
C300 VN.n1 B 0.289001f
C301 VN.n2 B 0.305161f
C302 VN.n3 B 0.046756f
C303 VN.t2 B 0.629118f
C304 VN.n4 B 0.301069f
C305 VN.n5 B 0.039303f
C306 VN.n6 B 0.225293f
C307 VN.t3 B 0.565469f
C308 VN.t4 B 0.665821f
C309 VN.n7 B 0.289001f
C310 VN.n8 B 0.305161f
C311 VN.n9 B 0.046756f
C312 VN.t0 B 0.629118f
C313 VN.n10 B 0.301069f
C314 VN.n11 B 1.44666f
.ends

