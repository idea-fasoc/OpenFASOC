* NGSPICE file created from diff_pair_sample_1219.ext - technology: sky130A

.subckt diff_pair_sample_1219 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=3.9156 pd=20.86 as=0 ps=0 w=10.04 l=1.11
X1 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=3.9156 pd=20.86 as=0 ps=0 w=10.04 l=1.11
X2 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.9156 pd=20.86 as=0 ps=0 w=10.04 l=1.11
X3 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.9156 pd=20.86 as=0 ps=0 w=10.04 l=1.11
X4 VDD2.t3 VN.t0 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6566 pd=10.37 as=3.9156 ps=20.86 w=10.04 l=1.11
X5 VTAIL.t2 VP.t0 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=3.9156 pd=20.86 as=1.6566 ps=10.37 w=10.04 l=1.11
X6 VDD2.t2 VN.t1 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6566 pd=10.37 as=3.9156 ps=20.86 w=10.04 l=1.11
X7 VTAIL.t7 VN.t2 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=3.9156 pd=20.86 as=1.6566 ps=10.37 w=10.04 l=1.11
X8 VDD1.t2 VP.t1 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6566 pd=10.37 as=3.9156 ps=20.86 w=10.04 l=1.11
X9 VTAIL.t3 VP.t2 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=3.9156 pd=20.86 as=1.6566 ps=10.37 w=10.04 l=1.11
X10 VDD1.t0 VP.t3 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6566 pd=10.37 as=3.9156 ps=20.86 w=10.04 l=1.11
X11 VTAIL.t4 VN.t3 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=3.9156 pd=20.86 as=1.6566 ps=10.37 w=10.04 l=1.11
R0 B.n587 B.n586 585
R1 B.n588 B.n587 585
R2 B.n247 B.n82 585
R3 B.n246 B.n245 585
R4 B.n244 B.n243 585
R5 B.n242 B.n241 585
R6 B.n240 B.n239 585
R7 B.n238 B.n237 585
R8 B.n236 B.n235 585
R9 B.n234 B.n233 585
R10 B.n232 B.n231 585
R11 B.n230 B.n229 585
R12 B.n228 B.n227 585
R13 B.n226 B.n225 585
R14 B.n224 B.n223 585
R15 B.n222 B.n221 585
R16 B.n220 B.n219 585
R17 B.n218 B.n217 585
R18 B.n216 B.n215 585
R19 B.n214 B.n213 585
R20 B.n212 B.n211 585
R21 B.n210 B.n209 585
R22 B.n208 B.n207 585
R23 B.n206 B.n205 585
R24 B.n204 B.n203 585
R25 B.n202 B.n201 585
R26 B.n200 B.n199 585
R27 B.n198 B.n197 585
R28 B.n196 B.n195 585
R29 B.n194 B.n193 585
R30 B.n192 B.n191 585
R31 B.n190 B.n189 585
R32 B.n188 B.n187 585
R33 B.n186 B.n185 585
R34 B.n184 B.n183 585
R35 B.n182 B.n181 585
R36 B.n180 B.n179 585
R37 B.n177 B.n176 585
R38 B.n175 B.n174 585
R39 B.n173 B.n172 585
R40 B.n171 B.n170 585
R41 B.n169 B.n168 585
R42 B.n167 B.n166 585
R43 B.n165 B.n164 585
R44 B.n163 B.n162 585
R45 B.n161 B.n160 585
R46 B.n159 B.n158 585
R47 B.n157 B.n156 585
R48 B.n155 B.n154 585
R49 B.n153 B.n152 585
R50 B.n151 B.n150 585
R51 B.n149 B.n148 585
R52 B.n147 B.n146 585
R53 B.n145 B.n144 585
R54 B.n143 B.n142 585
R55 B.n141 B.n140 585
R56 B.n139 B.n138 585
R57 B.n137 B.n136 585
R58 B.n135 B.n134 585
R59 B.n133 B.n132 585
R60 B.n131 B.n130 585
R61 B.n129 B.n128 585
R62 B.n127 B.n126 585
R63 B.n125 B.n124 585
R64 B.n123 B.n122 585
R65 B.n121 B.n120 585
R66 B.n119 B.n118 585
R67 B.n117 B.n116 585
R68 B.n115 B.n114 585
R69 B.n113 B.n112 585
R70 B.n111 B.n110 585
R71 B.n109 B.n108 585
R72 B.n107 B.n106 585
R73 B.n105 B.n104 585
R74 B.n103 B.n102 585
R75 B.n101 B.n100 585
R76 B.n99 B.n98 585
R77 B.n97 B.n96 585
R78 B.n95 B.n94 585
R79 B.n93 B.n92 585
R80 B.n91 B.n90 585
R81 B.n89 B.n88 585
R82 B.n585 B.n41 585
R83 B.n589 B.n41 585
R84 B.n584 B.n40 585
R85 B.n590 B.n40 585
R86 B.n583 B.n582 585
R87 B.n582 B.n36 585
R88 B.n581 B.n35 585
R89 B.n596 B.n35 585
R90 B.n580 B.n34 585
R91 B.n597 B.n34 585
R92 B.n579 B.n33 585
R93 B.n598 B.n33 585
R94 B.n578 B.n577 585
R95 B.n577 B.n29 585
R96 B.n576 B.n28 585
R97 B.n604 B.n28 585
R98 B.n575 B.n27 585
R99 B.n605 B.n27 585
R100 B.n574 B.n26 585
R101 B.n606 B.n26 585
R102 B.n573 B.n572 585
R103 B.n572 B.n22 585
R104 B.n571 B.n21 585
R105 B.n612 B.n21 585
R106 B.n570 B.n20 585
R107 B.n613 B.n20 585
R108 B.n569 B.n19 585
R109 B.n614 B.n19 585
R110 B.n568 B.n567 585
R111 B.n567 B.n15 585
R112 B.n566 B.n14 585
R113 B.n620 B.n14 585
R114 B.n565 B.n13 585
R115 B.n621 B.n13 585
R116 B.n564 B.n12 585
R117 B.n622 B.n12 585
R118 B.n563 B.n562 585
R119 B.n562 B.n8 585
R120 B.n561 B.n7 585
R121 B.n628 B.n7 585
R122 B.n560 B.n6 585
R123 B.n629 B.n6 585
R124 B.n559 B.n5 585
R125 B.n630 B.n5 585
R126 B.n558 B.n557 585
R127 B.n557 B.n4 585
R128 B.n556 B.n248 585
R129 B.n556 B.n555 585
R130 B.n546 B.n249 585
R131 B.n250 B.n249 585
R132 B.n548 B.n547 585
R133 B.n549 B.n548 585
R134 B.n545 B.n255 585
R135 B.n255 B.n254 585
R136 B.n544 B.n543 585
R137 B.n543 B.n542 585
R138 B.n257 B.n256 585
R139 B.n258 B.n257 585
R140 B.n535 B.n534 585
R141 B.n536 B.n535 585
R142 B.n533 B.n263 585
R143 B.n263 B.n262 585
R144 B.n532 B.n531 585
R145 B.n531 B.n530 585
R146 B.n265 B.n264 585
R147 B.n266 B.n265 585
R148 B.n523 B.n522 585
R149 B.n524 B.n523 585
R150 B.n521 B.n271 585
R151 B.n271 B.n270 585
R152 B.n520 B.n519 585
R153 B.n519 B.n518 585
R154 B.n273 B.n272 585
R155 B.n274 B.n273 585
R156 B.n511 B.n510 585
R157 B.n512 B.n511 585
R158 B.n509 B.n279 585
R159 B.n279 B.n278 585
R160 B.n508 B.n507 585
R161 B.n507 B.n506 585
R162 B.n281 B.n280 585
R163 B.n282 B.n281 585
R164 B.n499 B.n498 585
R165 B.n500 B.n499 585
R166 B.n497 B.n287 585
R167 B.n287 B.n286 585
R168 B.n491 B.n490 585
R169 B.n489 B.n329 585
R170 B.n488 B.n328 585
R171 B.n493 B.n328 585
R172 B.n487 B.n486 585
R173 B.n485 B.n484 585
R174 B.n483 B.n482 585
R175 B.n481 B.n480 585
R176 B.n479 B.n478 585
R177 B.n477 B.n476 585
R178 B.n475 B.n474 585
R179 B.n473 B.n472 585
R180 B.n471 B.n470 585
R181 B.n469 B.n468 585
R182 B.n467 B.n466 585
R183 B.n465 B.n464 585
R184 B.n463 B.n462 585
R185 B.n461 B.n460 585
R186 B.n459 B.n458 585
R187 B.n457 B.n456 585
R188 B.n455 B.n454 585
R189 B.n453 B.n452 585
R190 B.n451 B.n450 585
R191 B.n449 B.n448 585
R192 B.n447 B.n446 585
R193 B.n445 B.n444 585
R194 B.n443 B.n442 585
R195 B.n441 B.n440 585
R196 B.n439 B.n438 585
R197 B.n437 B.n436 585
R198 B.n435 B.n434 585
R199 B.n433 B.n432 585
R200 B.n431 B.n430 585
R201 B.n429 B.n428 585
R202 B.n427 B.n426 585
R203 B.n425 B.n424 585
R204 B.n423 B.n422 585
R205 B.n420 B.n419 585
R206 B.n418 B.n417 585
R207 B.n416 B.n415 585
R208 B.n414 B.n413 585
R209 B.n412 B.n411 585
R210 B.n410 B.n409 585
R211 B.n408 B.n407 585
R212 B.n406 B.n405 585
R213 B.n404 B.n403 585
R214 B.n402 B.n401 585
R215 B.n400 B.n399 585
R216 B.n398 B.n397 585
R217 B.n396 B.n395 585
R218 B.n394 B.n393 585
R219 B.n392 B.n391 585
R220 B.n390 B.n389 585
R221 B.n388 B.n387 585
R222 B.n386 B.n385 585
R223 B.n384 B.n383 585
R224 B.n382 B.n381 585
R225 B.n380 B.n379 585
R226 B.n378 B.n377 585
R227 B.n376 B.n375 585
R228 B.n374 B.n373 585
R229 B.n372 B.n371 585
R230 B.n370 B.n369 585
R231 B.n368 B.n367 585
R232 B.n366 B.n365 585
R233 B.n364 B.n363 585
R234 B.n362 B.n361 585
R235 B.n360 B.n359 585
R236 B.n358 B.n357 585
R237 B.n356 B.n355 585
R238 B.n354 B.n353 585
R239 B.n352 B.n351 585
R240 B.n350 B.n349 585
R241 B.n348 B.n347 585
R242 B.n346 B.n345 585
R243 B.n344 B.n343 585
R244 B.n342 B.n341 585
R245 B.n340 B.n339 585
R246 B.n338 B.n337 585
R247 B.n336 B.n335 585
R248 B.n289 B.n288 585
R249 B.n496 B.n495 585
R250 B.n285 B.n284 585
R251 B.n286 B.n285 585
R252 B.n502 B.n501 585
R253 B.n501 B.n500 585
R254 B.n503 B.n283 585
R255 B.n283 B.n282 585
R256 B.n505 B.n504 585
R257 B.n506 B.n505 585
R258 B.n277 B.n276 585
R259 B.n278 B.n277 585
R260 B.n514 B.n513 585
R261 B.n513 B.n512 585
R262 B.n515 B.n275 585
R263 B.n275 B.n274 585
R264 B.n517 B.n516 585
R265 B.n518 B.n517 585
R266 B.n269 B.n268 585
R267 B.n270 B.n269 585
R268 B.n526 B.n525 585
R269 B.n525 B.n524 585
R270 B.n527 B.n267 585
R271 B.n267 B.n266 585
R272 B.n529 B.n528 585
R273 B.n530 B.n529 585
R274 B.n261 B.n260 585
R275 B.n262 B.n261 585
R276 B.n538 B.n537 585
R277 B.n537 B.n536 585
R278 B.n539 B.n259 585
R279 B.n259 B.n258 585
R280 B.n541 B.n540 585
R281 B.n542 B.n541 585
R282 B.n253 B.n252 585
R283 B.n254 B.n253 585
R284 B.n551 B.n550 585
R285 B.n550 B.n549 585
R286 B.n552 B.n251 585
R287 B.n251 B.n250 585
R288 B.n554 B.n553 585
R289 B.n555 B.n554 585
R290 B.n2 B.n0 585
R291 B.n4 B.n2 585
R292 B.n3 B.n1 585
R293 B.n629 B.n3 585
R294 B.n627 B.n626 585
R295 B.n628 B.n627 585
R296 B.n625 B.n9 585
R297 B.n9 B.n8 585
R298 B.n624 B.n623 585
R299 B.n623 B.n622 585
R300 B.n11 B.n10 585
R301 B.n621 B.n11 585
R302 B.n619 B.n618 585
R303 B.n620 B.n619 585
R304 B.n617 B.n16 585
R305 B.n16 B.n15 585
R306 B.n616 B.n615 585
R307 B.n615 B.n614 585
R308 B.n18 B.n17 585
R309 B.n613 B.n18 585
R310 B.n611 B.n610 585
R311 B.n612 B.n611 585
R312 B.n609 B.n23 585
R313 B.n23 B.n22 585
R314 B.n608 B.n607 585
R315 B.n607 B.n606 585
R316 B.n25 B.n24 585
R317 B.n605 B.n25 585
R318 B.n603 B.n602 585
R319 B.n604 B.n603 585
R320 B.n601 B.n30 585
R321 B.n30 B.n29 585
R322 B.n600 B.n599 585
R323 B.n599 B.n598 585
R324 B.n32 B.n31 585
R325 B.n597 B.n32 585
R326 B.n595 B.n594 585
R327 B.n596 B.n595 585
R328 B.n593 B.n37 585
R329 B.n37 B.n36 585
R330 B.n592 B.n591 585
R331 B.n591 B.n590 585
R332 B.n39 B.n38 585
R333 B.n589 B.n39 585
R334 B.n632 B.n631 585
R335 B.n631 B.n630 585
R336 B.n491 B.n285 492.5
R337 B.n88 B.n39 492.5
R338 B.n495 B.n287 492.5
R339 B.n587 B.n41 492.5
R340 B.n332 B.t8 421.606
R341 B.n330 B.t15 421.606
R342 B.n85 B.t4 421.606
R343 B.n83 B.t12 421.606
R344 B.n332 B.t11 276.351
R345 B.n83 B.t13 276.351
R346 B.n330 B.t17 276.351
R347 B.n85 B.t6 276.351
R348 B.n588 B.n81 256.663
R349 B.n588 B.n80 256.663
R350 B.n588 B.n79 256.663
R351 B.n588 B.n78 256.663
R352 B.n588 B.n77 256.663
R353 B.n588 B.n76 256.663
R354 B.n588 B.n75 256.663
R355 B.n588 B.n74 256.663
R356 B.n588 B.n73 256.663
R357 B.n588 B.n72 256.663
R358 B.n588 B.n71 256.663
R359 B.n588 B.n70 256.663
R360 B.n588 B.n69 256.663
R361 B.n588 B.n68 256.663
R362 B.n588 B.n67 256.663
R363 B.n588 B.n66 256.663
R364 B.n588 B.n65 256.663
R365 B.n588 B.n64 256.663
R366 B.n588 B.n63 256.663
R367 B.n588 B.n62 256.663
R368 B.n588 B.n61 256.663
R369 B.n588 B.n60 256.663
R370 B.n588 B.n59 256.663
R371 B.n588 B.n58 256.663
R372 B.n588 B.n57 256.663
R373 B.n588 B.n56 256.663
R374 B.n588 B.n55 256.663
R375 B.n588 B.n54 256.663
R376 B.n588 B.n53 256.663
R377 B.n588 B.n52 256.663
R378 B.n588 B.n51 256.663
R379 B.n588 B.n50 256.663
R380 B.n588 B.n49 256.663
R381 B.n588 B.n48 256.663
R382 B.n588 B.n47 256.663
R383 B.n588 B.n46 256.663
R384 B.n588 B.n45 256.663
R385 B.n588 B.n44 256.663
R386 B.n588 B.n43 256.663
R387 B.n588 B.n42 256.663
R388 B.n493 B.n492 256.663
R389 B.n493 B.n290 256.663
R390 B.n493 B.n291 256.663
R391 B.n493 B.n292 256.663
R392 B.n493 B.n293 256.663
R393 B.n493 B.n294 256.663
R394 B.n493 B.n295 256.663
R395 B.n493 B.n296 256.663
R396 B.n493 B.n297 256.663
R397 B.n493 B.n298 256.663
R398 B.n493 B.n299 256.663
R399 B.n493 B.n300 256.663
R400 B.n493 B.n301 256.663
R401 B.n493 B.n302 256.663
R402 B.n493 B.n303 256.663
R403 B.n493 B.n304 256.663
R404 B.n493 B.n305 256.663
R405 B.n493 B.n306 256.663
R406 B.n493 B.n307 256.663
R407 B.n493 B.n308 256.663
R408 B.n493 B.n309 256.663
R409 B.n493 B.n310 256.663
R410 B.n493 B.n311 256.663
R411 B.n493 B.n312 256.663
R412 B.n493 B.n313 256.663
R413 B.n493 B.n314 256.663
R414 B.n493 B.n315 256.663
R415 B.n493 B.n316 256.663
R416 B.n493 B.n317 256.663
R417 B.n493 B.n318 256.663
R418 B.n493 B.n319 256.663
R419 B.n493 B.n320 256.663
R420 B.n493 B.n321 256.663
R421 B.n493 B.n322 256.663
R422 B.n493 B.n323 256.663
R423 B.n493 B.n324 256.663
R424 B.n493 B.n325 256.663
R425 B.n493 B.n326 256.663
R426 B.n493 B.n327 256.663
R427 B.n494 B.n493 256.663
R428 B.n333 B.t10 248.423
R429 B.n84 B.t14 248.423
R430 B.n331 B.t16 248.423
R431 B.n86 B.t7 248.423
R432 B.n501 B.n285 163.367
R433 B.n501 B.n283 163.367
R434 B.n505 B.n283 163.367
R435 B.n505 B.n277 163.367
R436 B.n513 B.n277 163.367
R437 B.n513 B.n275 163.367
R438 B.n517 B.n275 163.367
R439 B.n517 B.n269 163.367
R440 B.n525 B.n269 163.367
R441 B.n525 B.n267 163.367
R442 B.n529 B.n267 163.367
R443 B.n529 B.n261 163.367
R444 B.n537 B.n261 163.367
R445 B.n537 B.n259 163.367
R446 B.n541 B.n259 163.367
R447 B.n541 B.n253 163.367
R448 B.n550 B.n253 163.367
R449 B.n550 B.n251 163.367
R450 B.n554 B.n251 163.367
R451 B.n554 B.n2 163.367
R452 B.n631 B.n2 163.367
R453 B.n631 B.n3 163.367
R454 B.n627 B.n3 163.367
R455 B.n627 B.n9 163.367
R456 B.n623 B.n9 163.367
R457 B.n623 B.n11 163.367
R458 B.n619 B.n11 163.367
R459 B.n619 B.n16 163.367
R460 B.n615 B.n16 163.367
R461 B.n615 B.n18 163.367
R462 B.n611 B.n18 163.367
R463 B.n611 B.n23 163.367
R464 B.n607 B.n23 163.367
R465 B.n607 B.n25 163.367
R466 B.n603 B.n25 163.367
R467 B.n603 B.n30 163.367
R468 B.n599 B.n30 163.367
R469 B.n599 B.n32 163.367
R470 B.n595 B.n32 163.367
R471 B.n595 B.n37 163.367
R472 B.n591 B.n37 163.367
R473 B.n591 B.n39 163.367
R474 B.n329 B.n328 163.367
R475 B.n486 B.n328 163.367
R476 B.n484 B.n483 163.367
R477 B.n480 B.n479 163.367
R478 B.n476 B.n475 163.367
R479 B.n472 B.n471 163.367
R480 B.n468 B.n467 163.367
R481 B.n464 B.n463 163.367
R482 B.n460 B.n459 163.367
R483 B.n456 B.n455 163.367
R484 B.n452 B.n451 163.367
R485 B.n448 B.n447 163.367
R486 B.n444 B.n443 163.367
R487 B.n440 B.n439 163.367
R488 B.n436 B.n435 163.367
R489 B.n432 B.n431 163.367
R490 B.n428 B.n427 163.367
R491 B.n424 B.n423 163.367
R492 B.n419 B.n418 163.367
R493 B.n415 B.n414 163.367
R494 B.n411 B.n410 163.367
R495 B.n407 B.n406 163.367
R496 B.n403 B.n402 163.367
R497 B.n399 B.n398 163.367
R498 B.n395 B.n394 163.367
R499 B.n391 B.n390 163.367
R500 B.n387 B.n386 163.367
R501 B.n383 B.n382 163.367
R502 B.n379 B.n378 163.367
R503 B.n375 B.n374 163.367
R504 B.n371 B.n370 163.367
R505 B.n367 B.n366 163.367
R506 B.n363 B.n362 163.367
R507 B.n359 B.n358 163.367
R508 B.n355 B.n354 163.367
R509 B.n351 B.n350 163.367
R510 B.n347 B.n346 163.367
R511 B.n343 B.n342 163.367
R512 B.n339 B.n338 163.367
R513 B.n335 B.n289 163.367
R514 B.n499 B.n287 163.367
R515 B.n499 B.n281 163.367
R516 B.n507 B.n281 163.367
R517 B.n507 B.n279 163.367
R518 B.n511 B.n279 163.367
R519 B.n511 B.n273 163.367
R520 B.n519 B.n273 163.367
R521 B.n519 B.n271 163.367
R522 B.n523 B.n271 163.367
R523 B.n523 B.n265 163.367
R524 B.n531 B.n265 163.367
R525 B.n531 B.n263 163.367
R526 B.n535 B.n263 163.367
R527 B.n535 B.n257 163.367
R528 B.n543 B.n257 163.367
R529 B.n543 B.n255 163.367
R530 B.n548 B.n255 163.367
R531 B.n548 B.n249 163.367
R532 B.n556 B.n249 163.367
R533 B.n557 B.n556 163.367
R534 B.n557 B.n5 163.367
R535 B.n6 B.n5 163.367
R536 B.n7 B.n6 163.367
R537 B.n562 B.n7 163.367
R538 B.n562 B.n12 163.367
R539 B.n13 B.n12 163.367
R540 B.n14 B.n13 163.367
R541 B.n567 B.n14 163.367
R542 B.n567 B.n19 163.367
R543 B.n20 B.n19 163.367
R544 B.n21 B.n20 163.367
R545 B.n572 B.n21 163.367
R546 B.n572 B.n26 163.367
R547 B.n27 B.n26 163.367
R548 B.n28 B.n27 163.367
R549 B.n577 B.n28 163.367
R550 B.n577 B.n33 163.367
R551 B.n34 B.n33 163.367
R552 B.n35 B.n34 163.367
R553 B.n582 B.n35 163.367
R554 B.n582 B.n40 163.367
R555 B.n41 B.n40 163.367
R556 B.n92 B.n91 163.367
R557 B.n96 B.n95 163.367
R558 B.n100 B.n99 163.367
R559 B.n104 B.n103 163.367
R560 B.n108 B.n107 163.367
R561 B.n112 B.n111 163.367
R562 B.n116 B.n115 163.367
R563 B.n120 B.n119 163.367
R564 B.n124 B.n123 163.367
R565 B.n128 B.n127 163.367
R566 B.n132 B.n131 163.367
R567 B.n136 B.n135 163.367
R568 B.n140 B.n139 163.367
R569 B.n144 B.n143 163.367
R570 B.n148 B.n147 163.367
R571 B.n152 B.n151 163.367
R572 B.n156 B.n155 163.367
R573 B.n160 B.n159 163.367
R574 B.n164 B.n163 163.367
R575 B.n168 B.n167 163.367
R576 B.n172 B.n171 163.367
R577 B.n176 B.n175 163.367
R578 B.n181 B.n180 163.367
R579 B.n185 B.n184 163.367
R580 B.n189 B.n188 163.367
R581 B.n193 B.n192 163.367
R582 B.n197 B.n196 163.367
R583 B.n201 B.n200 163.367
R584 B.n205 B.n204 163.367
R585 B.n209 B.n208 163.367
R586 B.n213 B.n212 163.367
R587 B.n217 B.n216 163.367
R588 B.n221 B.n220 163.367
R589 B.n225 B.n224 163.367
R590 B.n229 B.n228 163.367
R591 B.n233 B.n232 163.367
R592 B.n237 B.n236 163.367
R593 B.n241 B.n240 163.367
R594 B.n245 B.n244 163.367
R595 B.n587 B.n82 163.367
R596 B.n493 B.n286 79.7263
R597 B.n589 B.n588 79.7263
R598 B.n492 B.n491 71.676
R599 B.n486 B.n290 71.676
R600 B.n483 B.n291 71.676
R601 B.n479 B.n292 71.676
R602 B.n475 B.n293 71.676
R603 B.n471 B.n294 71.676
R604 B.n467 B.n295 71.676
R605 B.n463 B.n296 71.676
R606 B.n459 B.n297 71.676
R607 B.n455 B.n298 71.676
R608 B.n451 B.n299 71.676
R609 B.n447 B.n300 71.676
R610 B.n443 B.n301 71.676
R611 B.n439 B.n302 71.676
R612 B.n435 B.n303 71.676
R613 B.n431 B.n304 71.676
R614 B.n427 B.n305 71.676
R615 B.n423 B.n306 71.676
R616 B.n418 B.n307 71.676
R617 B.n414 B.n308 71.676
R618 B.n410 B.n309 71.676
R619 B.n406 B.n310 71.676
R620 B.n402 B.n311 71.676
R621 B.n398 B.n312 71.676
R622 B.n394 B.n313 71.676
R623 B.n390 B.n314 71.676
R624 B.n386 B.n315 71.676
R625 B.n382 B.n316 71.676
R626 B.n378 B.n317 71.676
R627 B.n374 B.n318 71.676
R628 B.n370 B.n319 71.676
R629 B.n366 B.n320 71.676
R630 B.n362 B.n321 71.676
R631 B.n358 B.n322 71.676
R632 B.n354 B.n323 71.676
R633 B.n350 B.n324 71.676
R634 B.n346 B.n325 71.676
R635 B.n342 B.n326 71.676
R636 B.n338 B.n327 71.676
R637 B.n494 B.n289 71.676
R638 B.n88 B.n42 71.676
R639 B.n92 B.n43 71.676
R640 B.n96 B.n44 71.676
R641 B.n100 B.n45 71.676
R642 B.n104 B.n46 71.676
R643 B.n108 B.n47 71.676
R644 B.n112 B.n48 71.676
R645 B.n116 B.n49 71.676
R646 B.n120 B.n50 71.676
R647 B.n124 B.n51 71.676
R648 B.n128 B.n52 71.676
R649 B.n132 B.n53 71.676
R650 B.n136 B.n54 71.676
R651 B.n140 B.n55 71.676
R652 B.n144 B.n56 71.676
R653 B.n148 B.n57 71.676
R654 B.n152 B.n58 71.676
R655 B.n156 B.n59 71.676
R656 B.n160 B.n60 71.676
R657 B.n164 B.n61 71.676
R658 B.n168 B.n62 71.676
R659 B.n172 B.n63 71.676
R660 B.n176 B.n64 71.676
R661 B.n181 B.n65 71.676
R662 B.n185 B.n66 71.676
R663 B.n189 B.n67 71.676
R664 B.n193 B.n68 71.676
R665 B.n197 B.n69 71.676
R666 B.n201 B.n70 71.676
R667 B.n205 B.n71 71.676
R668 B.n209 B.n72 71.676
R669 B.n213 B.n73 71.676
R670 B.n217 B.n74 71.676
R671 B.n221 B.n75 71.676
R672 B.n225 B.n76 71.676
R673 B.n229 B.n77 71.676
R674 B.n233 B.n78 71.676
R675 B.n237 B.n79 71.676
R676 B.n241 B.n80 71.676
R677 B.n245 B.n81 71.676
R678 B.n82 B.n81 71.676
R679 B.n244 B.n80 71.676
R680 B.n240 B.n79 71.676
R681 B.n236 B.n78 71.676
R682 B.n232 B.n77 71.676
R683 B.n228 B.n76 71.676
R684 B.n224 B.n75 71.676
R685 B.n220 B.n74 71.676
R686 B.n216 B.n73 71.676
R687 B.n212 B.n72 71.676
R688 B.n208 B.n71 71.676
R689 B.n204 B.n70 71.676
R690 B.n200 B.n69 71.676
R691 B.n196 B.n68 71.676
R692 B.n192 B.n67 71.676
R693 B.n188 B.n66 71.676
R694 B.n184 B.n65 71.676
R695 B.n180 B.n64 71.676
R696 B.n175 B.n63 71.676
R697 B.n171 B.n62 71.676
R698 B.n167 B.n61 71.676
R699 B.n163 B.n60 71.676
R700 B.n159 B.n59 71.676
R701 B.n155 B.n58 71.676
R702 B.n151 B.n57 71.676
R703 B.n147 B.n56 71.676
R704 B.n143 B.n55 71.676
R705 B.n139 B.n54 71.676
R706 B.n135 B.n53 71.676
R707 B.n131 B.n52 71.676
R708 B.n127 B.n51 71.676
R709 B.n123 B.n50 71.676
R710 B.n119 B.n49 71.676
R711 B.n115 B.n48 71.676
R712 B.n111 B.n47 71.676
R713 B.n107 B.n46 71.676
R714 B.n103 B.n45 71.676
R715 B.n99 B.n44 71.676
R716 B.n95 B.n43 71.676
R717 B.n91 B.n42 71.676
R718 B.n492 B.n329 71.676
R719 B.n484 B.n290 71.676
R720 B.n480 B.n291 71.676
R721 B.n476 B.n292 71.676
R722 B.n472 B.n293 71.676
R723 B.n468 B.n294 71.676
R724 B.n464 B.n295 71.676
R725 B.n460 B.n296 71.676
R726 B.n456 B.n297 71.676
R727 B.n452 B.n298 71.676
R728 B.n448 B.n299 71.676
R729 B.n444 B.n300 71.676
R730 B.n440 B.n301 71.676
R731 B.n436 B.n302 71.676
R732 B.n432 B.n303 71.676
R733 B.n428 B.n304 71.676
R734 B.n424 B.n305 71.676
R735 B.n419 B.n306 71.676
R736 B.n415 B.n307 71.676
R737 B.n411 B.n308 71.676
R738 B.n407 B.n309 71.676
R739 B.n403 B.n310 71.676
R740 B.n399 B.n311 71.676
R741 B.n395 B.n312 71.676
R742 B.n391 B.n313 71.676
R743 B.n387 B.n314 71.676
R744 B.n383 B.n315 71.676
R745 B.n379 B.n316 71.676
R746 B.n375 B.n317 71.676
R747 B.n371 B.n318 71.676
R748 B.n367 B.n319 71.676
R749 B.n363 B.n320 71.676
R750 B.n359 B.n321 71.676
R751 B.n355 B.n322 71.676
R752 B.n351 B.n323 71.676
R753 B.n347 B.n324 71.676
R754 B.n343 B.n325 71.676
R755 B.n339 B.n326 71.676
R756 B.n335 B.n327 71.676
R757 B.n495 B.n494 71.676
R758 B.n334 B.n333 59.5399
R759 B.n421 B.n331 59.5399
R760 B.n87 B.n86 59.5399
R761 B.n178 B.n84 59.5399
R762 B.n500 B.n286 48.8415
R763 B.n500 B.n282 48.8415
R764 B.n506 B.n282 48.8415
R765 B.n506 B.n278 48.8415
R766 B.n512 B.n278 48.8415
R767 B.n518 B.n274 48.8415
R768 B.n518 B.n270 48.8415
R769 B.n524 B.n270 48.8415
R770 B.n524 B.n266 48.8415
R771 B.n530 B.n266 48.8415
R772 B.n530 B.n262 48.8415
R773 B.n536 B.n262 48.8415
R774 B.n542 B.n258 48.8415
R775 B.n542 B.n254 48.8415
R776 B.n549 B.n254 48.8415
R777 B.n555 B.n250 48.8415
R778 B.n555 B.n4 48.8415
R779 B.n630 B.n4 48.8415
R780 B.n630 B.n629 48.8415
R781 B.n629 B.n628 48.8415
R782 B.n628 B.n8 48.8415
R783 B.n622 B.n621 48.8415
R784 B.n621 B.n620 48.8415
R785 B.n620 B.n15 48.8415
R786 B.n614 B.n613 48.8415
R787 B.n613 B.n612 48.8415
R788 B.n612 B.n22 48.8415
R789 B.n606 B.n22 48.8415
R790 B.n606 B.n605 48.8415
R791 B.n605 B.n604 48.8415
R792 B.n604 B.n29 48.8415
R793 B.n598 B.n597 48.8415
R794 B.n597 B.n596 48.8415
R795 B.n596 B.n36 48.8415
R796 B.n590 B.n36 48.8415
R797 B.n590 B.n589 48.8415
R798 B.t2 B.n258 46.6868
R799 B.t0 B.n15 46.6868
R800 B.t1 B.n250 35.1948
R801 B.t3 B.n8 35.1948
R802 B.n89 B.n38 32.0005
R803 B.n586 B.n585 32.0005
R804 B.n497 B.n496 32.0005
R805 B.n490 B.n284 32.0005
R806 B.n512 B.t9 29.4488
R807 B.n598 B.t5 29.4488
R808 B.n333 B.n332 27.9278
R809 B.n331 B.n330 27.9278
R810 B.n86 B.n85 27.9278
R811 B.n84 B.n83 27.9278
R812 B.t9 B.n274 19.3933
R813 B.t5 B.n29 19.3933
R814 B B.n632 18.0485
R815 B.n549 B.t1 13.6473
R816 B.n622 B.t3 13.6473
R817 B.n90 B.n89 10.6151
R818 B.n93 B.n90 10.6151
R819 B.n94 B.n93 10.6151
R820 B.n97 B.n94 10.6151
R821 B.n98 B.n97 10.6151
R822 B.n101 B.n98 10.6151
R823 B.n102 B.n101 10.6151
R824 B.n105 B.n102 10.6151
R825 B.n106 B.n105 10.6151
R826 B.n109 B.n106 10.6151
R827 B.n110 B.n109 10.6151
R828 B.n113 B.n110 10.6151
R829 B.n114 B.n113 10.6151
R830 B.n117 B.n114 10.6151
R831 B.n118 B.n117 10.6151
R832 B.n121 B.n118 10.6151
R833 B.n122 B.n121 10.6151
R834 B.n125 B.n122 10.6151
R835 B.n126 B.n125 10.6151
R836 B.n129 B.n126 10.6151
R837 B.n130 B.n129 10.6151
R838 B.n133 B.n130 10.6151
R839 B.n134 B.n133 10.6151
R840 B.n137 B.n134 10.6151
R841 B.n138 B.n137 10.6151
R842 B.n141 B.n138 10.6151
R843 B.n142 B.n141 10.6151
R844 B.n145 B.n142 10.6151
R845 B.n146 B.n145 10.6151
R846 B.n149 B.n146 10.6151
R847 B.n150 B.n149 10.6151
R848 B.n153 B.n150 10.6151
R849 B.n154 B.n153 10.6151
R850 B.n157 B.n154 10.6151
R851 B.n158 B.n157 10.6151
R852 B.n162 B.n161 10.6151
R853 B.n165 B.n162 10.6151
R854 B.n166 B.n165 10.6151
R855 B.n169 B.n166 10.6151
R856 B.n170 B.n169 10.6151
R857 B.n173 B.n170 10.6151
R858 B.n174 B.n173 10.6151
R859 B.n177 B.n174 10.6151
R860 B.n182 B.n179 10.6151
R861 B.n183 B.n182 10.6151
R862 B.n186 B.n183 10.6151
R863 B.n187 B.n186 10.6151
R864 B.n190 B.n187 10.6151
R865 B.n191 B.n190 10.6151
R866 B.n194 B.n191 10.6151
R867 B.n195 B.n194 10.6151
R868 B.n198 B.n195 10.6151
R869 B.n199 B.n198 10.6151
R870 B.n202 B.n199 10.6151
R871 B.n203 B.n202 10.6151
R872 B.n206 B.n203 10.6151
R873 B.n207 B.n206 10.6151
R874 B.n210 B.n207 10.6151
R875 B.n211 B.n210 10.6151
R876 B.n214 B.n211 10.6151
R877 B.n215 B.n214 10.6151
R878 B.n218 B.n215 10.6151
R879 B.n219 B.n218 10.6151
R880 B.n222 B.n219 10.6151
R881 B.n223 B.n222 10.6151
R882 B.n226 B.n223 10.6151
R883 B.n227 B.n226 10.6151
R884 B.n230 B.n227 10.6151
R885 B.n231 B.n230 10.6151
R886 B.n234 B.n231 10.6151
R887 B.n235 B.n234 10.6151
R888 B.n238 B.n235 10.6151
R889 B.n239 B.n238 10.6151
R890 B.n242 B.n239 10.6151
R891 B.n243 B.n242 10.6151
R892 B.n246 B.n243 10.6151
R893 B.n247 B.n246 10.6151
R894 B.n586 B.n247 10.6151
R895 B.n498 B.n497 10.6151
R896 B.n498 B.n280 10.6151
R897 B.n508 B.n280 10.6151
R898 B.n509 B.n508 10.6151
R899 B.n510 B.n509 10.6151
R900 B.n510 B.n272 10.6151
R901 B.n520 B.n272 10.6151
R902 B.n521 B.n520 10.6151
R903 B.n522 B.n521 10.6151
R904 B.n522 B.n264 10.6151
R905 B.n532 B.n264 10.6151
R906 B.n533 B.n532 10.6151
R907 B.n534 B.n533 10.6151
R908 B.n534 B.n256 10.6151
R909 B.n544 B.n256 10.6151
R910 B.n545 B.n544 10.6151
R911 B.n547 B.n545 10.6151
R912 B.n547 B.n546 10.6151
R913 B.n546 B.n248 10.6151
R914 B.n558 B.n248 10.6151
R915 B.n559 B.n558 10.6151
R916 B.n560 B.n559 10.6151
R917 B.n561 B.n560 10.6151
R918 B.n563 B.n561 10.6151
R919 B.n564 B.n563 10.6151
R920 B.n565 B.n564 10.6151
R921 B.n566 B.n565 10.6151
R922 B.n568 B.n566 10.6151
R923 B.n569 B.n568 10.6151
R924 B.n570 B.n569 10.6151
R925 B.n571 B.n570 10.6151
R926 B.n573 B.n571 10.6151
R927 B.n574 B.n573 10.6151
R928 B.n575 B.n574 10.6151
R929 B.n576 B.n575 10.6151
R930 B.n578 B.n576 10.6151
R931 B.n579 B.n578 10.6151
R932 B.n580 B.n579 10.6151
R933 B.n581 B.n580 10.6151
R934 B.n583 B.n581 10.6151
R935 B.n584 B.n583 10.6151
R936 B.n585 B.n584 10.6151
R937 B.n490 B.n489 10.6151
R938 B.n489 B.n488 10.6151
R939 B.n488 B.n487 10.6151
R940 B.n487 B.n485 10.6151
R941 B.n485 B.n482 10.6151
R942 B.n482 B.n481 10.6151
R943 B.n481 B.n478 10.6151
R944 B.n478 B.n477 10.6151
R945 B.n477 B.n474 10.6151
R946 B.n474 B.n473 10.6151
R947 B.n473 B.n470 10.6151
R948 B.n470 B.n469 10.6151
R949 B.n469 B.n466 10.6151
R950 B.n466 B.n465 10.6151
R951 B.n465 B.n462 10.6151
R952 B.n462 B.n461 10.6151
R953 B.n461 B.n458 10.6151
R954 B.n458 B.n457 10.6151
R955 B.n457 B.n454 10.6151
R956 B.n454 B.n453 10.6151
R957 B.n453 B.n450 10.6151
R958 B.n450 B.n449 10.6151
R959 B.n449 B.n446 10.6151
R960 B.n446 B.n445 10.6151
R961 B.n445 B.n442 10.6151
R962 B.n442 B.n441 10.6151
R963 B.n441 B.n438 10.6151
R964 B.n438 B.n437 10.6151
R965 B.n437 B.n434 10.6151
R966 B.n434 B.n433 10.6151
R967 B.n433 B.n430 10.6151
R968 B.n430 B.n429 10.6151
R969 B.n429 B.n426 10.6151
R970 B.n426 B.n425 10.6151
R971 B.n425 B.n422 10.6151
R972 B.n420 B.n417 10.6151
R973 B.n417 B.n416 10.6151
R974 B.n416 B.n413 10.6151
R975 B.n413 B.n412 10.6151
R976 B.n412 B.n409 10.6151
R977 B.n409 B.n408 10.6151
R978 B.n408 B.n405 10.6151
R979 B.n405 B.n404 10.6151
R980 B.n401 B.n400 10.6151
R981 B.n400 B.n397 10.6151
R982 B.n397 B.n396 10.6151
R983 B.n396 B.n393 10.6151
R984 B.n393 B.n392 10.6151
R985 B.n392 B.n389 10.6151
R986 B.n389 B.n388 10.6151
R987 B.n388 B.n385 10.6151
R988 B.n385 B.n384 10.6151
R989 B.n384 B.n381 10.6151
R990 B.n381 B.n380 10.6151
R991 B.n380 B.n377 10.6151
R992 B.n377 B.n376 10.6151
R993 B.n376 B.n373 10.6151
R994 B.n373 B.n372 10.6151
R995 B.n372 B.n369 10.6151
R996 B.n369 B.n368 10.6151
R997 B.n368 B.n365 10.6151
R998 B.n365 B.n364 10.6151
R999 B.n364 B.n361 10.6151
R1000 B.n361 B.n360 10.6151
R1001 B.n360 B.n357 10.6151
R1002 B.n357 B.n356 10.6151
R1003 B.n356 B.n353 10.6151
R1004 B.n353 B.n352 10.6151
R1005 B.n352 B.n349 10.6151
R1006 B.n349 B.n348 10.6151
R1007 B.n348 B.n345 10.6151
R1008 B.n345 B.n344 10.6151
R1009 B.n344 B.n341 10.6151
R1010 B.n341 B.n340 10.6151
R1011 B.n340 B.n337 10.6151
R1012 B.n337 B.n336 10.6151
R1013 B.n336 B.n288 10.6151
R1014 B.n496 B.n288 10.6151
R1015 B.n502 B.n284 10.6151
R1016 B.n503 B.n502 10.6151
R1017 B.n504 B.n503 10.6151
R1018 B.n504 B.n276 10.6151
R1019 B.n514 B.n276 10.6151
R1020 B.n515 B.n514 10.6151
R1021 B.n516 B.n515 10.6151
R1022 B.n516 B.n268 10.6151
R1023 B.n526 B.n268 10.6151
R1024 B.n527 B.n526 10.6151
R1025 B.n528 B.n527 10.6151
R1026 B.n528 B.n260 10.6151
R1027 B.n538 B.n260 10.6151
R1028 B.n539 B.n538 10.6151
R1029 B.n540 B.n539 10.6151
R1030 B.n540 B.n252 10.6151
R1031 B.n551 B.n252 10.6151
R1032 B.n552 B.n551 10.6151
R1033 B.n553 B.n552 10.6151
R1034 B.n553 B.n0 10.6151
R1035 B.n626 B.n1 10.6151
R1036 B.n626 B.n625 10.6151
R1037 B.n625 B.n624 10.6151
R1038 B.n624 B.n10 10.6151
R1039 B.n618 B.n10 10.6151
R1040 B.n618 B.n617 10.6151
R1041 B.n617 B.n616 10.6151
R1042 B.n616 B.n17 10.6151
R1043 B.n610 B.n17 10.6151
R1044 B.n610 B.n609 10.6151
R1045 B.n609 B.n608 10.6151
R1046 B.n608 B.n24 10.6151
R1047 B.n602 B.n24 10.6151
R1048 B.n602 B.n601 10.6151
R1049 B.n601 B.n600 10.6151
R1050 B.n600 B.n31 10.6151
R1051 B.n594 B.n31 10.6151
R1052 B.n594 B.n593 10.6151
R1053 B.n593 B.n592 10.6151
R1054 B.n592 B.n38 10.6151
R1055 B.n161 B.n87 6.5566
R1056 B.n178 B.n177 6.5566
R1057 B.n421 B.n420 6.5566
R1058 B.n404 B.n334 6.5566
R1059 B.n158 B.n87 4.05904
R1060 B.n179 B.n178 4.05904
R1061 B.n422 B.n421 4.05904
R1062 B.n401 B.n334 4.05904
R1063 B.n632 B.n0 2.81026
R1064 B.n632 B.n1 2.81026
R1065 B.n536 B.t2 2.15525
R1066 B.n614 B.t0 2.15525
R1067 VN.n0 VN.t3 271.983
R1068 VN.n1 VN.t1 271.983
R1069 VN.n1 VN.t2 271.896
R1070 VN.n0 VN.t0 271.896
R1071 VN VN.n1 71.8796
R1072 VN VN.n0 31.2622
R1073 VTAIL.n426 VTAIL.n378 289.615
R1074 VTAIL.n48 VTAIL.n0 289.615
R1075 VTAIL.n102 VTAIL.n54 289.615
R1076 VTAIL.n156 VTAIL.n108 289.615
R1077 VTAIL.n372 VTAIL.n324 289.615
R1078 VTAIL.n318 VTAIL.n270 289.615
R1079 VTAIL.n264 VTAIL.n216 289.615
R1080 VTAIL.n210 VTAIL.n162 289.615
R1081 VTAIL.n394 VTAIL.n393 185
R1082 VTAIL.n399 VTAIL.n398 185
R1083 VTAIL.n401 VTAIL.n400 185
R1084 VTAIL.n390 VTAIL.n389 185
R1085 VTAIL.n407 VTAIL.n406 185
R1086 VTAIL.n409 VTAIL.n408 185
R1087 VTAIL.n386 VTAIL.n385 185
R1088 VTAIL.n416 VTAIL.n415 185
R1089 VTAIL.n417 VTAIL.n384 185
R1090 VTAIL.n419 VTAIL.n418 185
R1091 VTAIL.n382 VTAIL.n381 185
R1092 VTAIL.n425 VTAIL.n424 185
R1093 VTAIL.n427 VTAIL.n426 185
R1094 VTAIL.n16 VTAIL.n15 185
R1095 VTAIL.n21 VTAIL.n20 185
R1096 VTAIL.n23 VTAIL.n22 185
R1097 VTAIL.n12 VTAIL.n11 185
R1098 VTAIL.n29 VTAIL.n28 185
R1099 VTAIL.n31 VTAIL.n30 185
R1100 VTAIL.n8 VTAIL.n7 185
R1101 VTAIL.n38 VTAIL.n37 185
R1102 VTAIL.n39 VTAIL.n6 185
R1103 VTAIL.n41 VTAIL.n40 185
R1104 VTAIL.n4 VTAIL.n3 185
R1105 VTAIL.n47 VTAIL.n46 185
R1106 VTAIL.n49 VTAIL.n48 185
R1107 VTAIL.n70 VTAIL.n69 185
R1108 VTAIL.n75 VTAIL.n74 185
R1109 VTAIL.n77 VTAIL.n76 185
R1110 VTAIL.n66 VTAIL.n65 185
R1111 VTAIL.n83 VTAIL.n82 185
R1112 VTAIL.n85 VTAIL.n84 185
R1113 VTAIL.n62 VTAIL.n61 185
R1114 VTAIL.n92 VTAIL.n91 185
R1115 VTAIL.n93 VTAIL.n60 185
R1116 VTAIL.n95 VTAIL.n94 185
R1117 VTAIL.n58 VTAIL.n57 185
R1118 VTAIL.n101 VTAIL.n100 185
R1119 VTAIL.n103 VTAIL.n102 185
R1120 VTAIL.n124 VTAIL.n123 185
R1121 VTAIL.n129 VTAIL.n128 185
R1122 VTAIL.n131 VTAIL.n130 185
R1123 VTAIL.n120 VTAIL.n119 185
R1124 VTAIL.n137 VTAIL.n136 185
R1125 VTAIL.n139 VTAIL.n138 185
R1126 VTAIL.n116 VTAIL.n115 185
R1127 VTAIL.n146 VTAIL.n145 185
R1128 VTAIL.n147 VTAIL.n114 185
R1129 VTAIL.n149 VTAIL.n148 185
R1130 VTAIL.n112 VTAIL.n111 185
R1131 VTAIL.n155 VTAIL.n154 185
R1132 VTAIL.n157 VTAIL.n156 185
R1133 VTAIL.n373 VTAIL.n372 185
R1134 VTAIL.n371 VTAIL.n370 185
R1135 VTAIL.n328 VTAIL.n327 185
R1136 VTAIL.n365 VTAIL.n364 185
R1137 VTAIL.n363 VTAIL.n330 185
R1138 VTAIL.n362 VTAIL.n361 185
R1139 VTAIL.n333 VTAIL.n331 185
R1140 VTAIL.n356 VTAIL.n355 185
R1141 VTAIL.n354 VTAIL.n353 185
R1142 VTAIL.n337 VTAIL.n336 185
R1143 VTAIL.n348 VTAIL.n347 185
R1144 VTAIL.n346 VTAIL.n345 185
R1145 VTAIL.n341 VTAIL.n340 185
R1146 VTAIL.n319 VTAIL.n318 185
R1147 VTAIL.n317 VTAIL.n316 185
R1148 VTAIL.n274 VTAIL.n273 185
R1149 VTAIL.n311 VTAIL.n310 185
R1150 VTAIL.n309 VTAIL.n276 185
R1151 VTAIL.n308 VTAIL.n307 185
R1152 VTAIL.n279 VTAIL.n277 185
R1153 VTAIL.n302 VTAIL.n301 185
R1154 VTAIL.n300 VTAIL.n299 185
R1155 VTAIL.n283 VTAIL.n282 185
R1156 VTAIL.n294 VTAIL.n293 185
R1157 VTAIL.n292 VTAIL.n291 185
R1158 VTAIL.n287 VTAIL.n286 185
R1159 VTAIL.n265 VTAIL.n264 185
R1160 VTAIL.n263 VTAIL.n262 185
R1161 VTAIL.n220 VTAIL.n219 185
R1162 VTAIL.n257 VTAIL.n256 185
R1163 VTAIL.n255 VTAIL.n222 185
R1164 VTAIL.n254 VTAIL.n253 185
R1165 VTAIL.n225 VTAIL.n223 185
R1166 VTAIL.n248 VTAIL.n247 185
R1167 VTAIL.n246 VTAIL.n245 185
R1168 VTAIL.n229 VTAIL.n228 185
R1169 VTAIL.n240 VTAIL.n239 185
R1170 VTAIL.n238 VTAIL.n237 185
R1171 VTAIL.n233 VTAIL.n232 185
R1172 VTAIL.n211 VTAIL.n210 185
R1173 VTAIL.n209 VTAIL.n208 185
R1174 VTAIL.n166 VTAIL.n165 185
R1175 VTAIL.n203 VTAIL.n202 185
R1176 VTAIL.n201 VTAIL.n168 185
R1177 VTAIL.n200 VTAIL.n199 185
R1178 VTAIL.n171 VTAIL.n169 185
R1179 VTAIL.n194 VTAIL.n193 185
R1180 VTAIL.n192 VTAIL.n191 185
R1181 VTAIL.n175 VTAIL.n174 185
R1182 VTAIL.n186 VTAIL.n185 185
R1183 VTAIL.n184 VTAIL.n183 185
R1184 VTAIL.n179 VTAIL.n178 185
R1185 VTAIL.n395 VTAIL.t6 149.524
R1186 VTAIL.n17 VTAIL.t4 149.524
R1187 VTAIL.n71 VTAIL.t0 149.524
R1188 VTAIL.n125 VTAIL.t2 149.524
R1189 VTAIL.n342 VTAIL.t1 149.524
R1190 VTAIL.n288 VTAIL.t3 149.524
R1191 VTAIL.n234 VTAIL.t5 149.524
R1192 VTAIL.n180 VTAIL.t7 149.524
R1193 VTAIL.n399 VTAIL.n393 104.615
R1194 VTAIL.n400 VTAIL.n399 104.615
R1195 VTAIL.n400 VTAIL.n389 104.615
R1196 VTAIL.n407 VTAIL.n389 104.615
R1197 VTAIL.n408 VTAIL.n407 104.615
R1198 VTAIL.n408 VTAIL.n385 104.615
R1199 VTAIL.n416 VTAIL.n385 104.615
R1200 VTAIL.n417 VTAIL.n416 104.615
R1201 VTAIL.n418 VTAIL.n417 104.615
R1202 VTAIL.n418 VTAIL.n381 104.615
R1203 VTAIL.n425 VTAIL.n381 104.615
R1204 VTAIL.n426 VTAIL.n425 104.615
R1205 VTAIL.n21 VTAIL.n15 104.615
R1206 VTAIL.n22 VTAIL.n21 104.615
R1207 VTAIL.n22 VTAIL.n11 104.615
R1208 VTAIL.n29 VTAIL.n11 104.615
R1209 VTAIL.n30 VTAIL.n29 104.615
R1210 VTAIL.n30 VTAIL.n7 104.615
R1211 VTAIL.n38 VTAIL.n7 104.615
R1212 VTAIL.n39 VTAIL.n38 104.615
R1213 VTAIL.n40 VTAIL.n39 104.615
R1214 VTAIL.n40 VTAIL.n3 104.615
R1215 VTAIL.n47 VTAIL.n3 104.615
R1216 VTAIL.n48 VTAIL.n47 104.615
R1217 VTAIL.n75 VTAIL.n69 104.615
R1218 VTAIL.n76 VTAIL.n75 104.615
R1219 VTAIL.n76 VTAIL.n65 104.615
R1220 VTAIL.n83 VTAIL.n65 104.615
R1221 VTAIL.n84 VTAIL.n83 104.615
R1222 VTAIL.n84 VTAIL.n61 104.615
R1223 VTAIL.n92 VTAIL.n61 104.615
R1224 VTAIL.n93 VTAIL.n92 104.615
R1225 VTAIL.n94 VTAIL.n93 104.615
R1226 VTAIL.n94 VTAIL.n57 104.615
R1227 VTAIL.n101 VTAIL.n57 104.615
R1228 VTAIL.n102 VTAIL.n101 104.615
R1229 VTAIL.n129 VTAIL.n123 104.615
R1230 VTAIL.n130 VTAIL.n129 104.615
R1231 VTAIL.n130 VTAIL.n119 104.615
R1232 VTAIL.n137 VTAIL.n119 104.615
R1233 VTAIL.n138 VTAIL.n137 104.615
R1234 VTAIL.n138 VTAIL.n115 104.615
R1235 VTAIL.n146 VTAIL.n115 104.615
R1236 VTAIL.n147 VTAIL.n146 104.615
R1237 VTAIL.n148 VTAIL.n147 104.615
R1238 VTAIL.n148 VTAIL.n111 104.615
R1239 VTAIL.n155 VTAIL.n111 104.615
R1240 VTAIL.n156 VTAIL.n155 104.615
R1241 VTAIL.n372 VTAIL.n371 104.615
R1242 VTAIL.n371 VTAIL.n327 104.615
R1243 VTAIL.n364 VTAIL.n327 104.615
R1244 VTAIL.n364 VTAIL.n363 104.615
R1245 VTAIL.n363 VTAIL.n362 104.615
R1246 VTAIL.n362 VTAIL.n331 104.615
R1247 VTAIL.n355 VTAIL.n331 104.615
R1248 VTAIL.n355 VTAIL.n354 104.615
R1249 VTAIL.n354 VTAIL.n336 104.615
R1250 VTAIL.n347 VTAIL.n336 104.615
R1251 VTAIL.n347 VTAIL.n346 104.615
R1252 VTAIL.n346 VTAIL.n340 104.615
R1253 VTAIL.n318 VTAIL.n317 104.615
R1254 VTAIL.n317 VTAIL.n273 104.615
R1255 VTAIL.n310 VTAIL.n273 104.615
R1256 VTAIL.n310 VTAIL.n309 104.615
R1257 VTAIL.n309 VTAIL.n308 104.615
R1258 VTAIL.n308 VTAIL.n277 104.615
R1259 VTAIL.n301 VTAIL.n277 104.615
R1260 VTAIL.n301 VTAIL.n300 104.615
R1261 VTAIL.n300 VTAIL.n282 104.615
R1262 VTAIL.n293 VTAIL.n282 104.615
R1263 VTAIL.n293 VTAIL.n292 104.615
R1264 VTAIL.n292 VTAIL.n286 104.615
R1265 VTAIL.n264 VTAIL.n263 104.615
R1266 VTAIL.n263 VTAIL.n219 104.615
R1267 VTAIL.n256 VTAIL.n219 104.615
R1268 VTAIL.n256 VTAIL.n255 104.615
R1269 VTAIL.n255 VTAIL.n254 104.615
R1270 VTAIL.n254 VTAIL.n223 104.615
R1271 VTAIL.n247 VTAIL.n223 104.615
R1272 VTAIL.n247 VTAIL.n246 104.615
R1273 VTAIL.n246 VTAIL.n228 104.615
R1274 VTAIL.n239 VTAIL.n228 104.615
R1275 VTAIL.n239 VTAIL.n238 104.615
R1276 VTAIL.n238 VTAIL.n232 104.615
R1277 VTAIL.n210 VTAIL.n209 104.615
R1278 VTAIL.n209 VTAIL.n165 104.615
R1279 VTAIL.n202 VTAIL.n165 104.615
R1280 VTAIL.n202 VTAIL.n201 104.615
R1281 VTAIL.n201 VTAIL.n200 104.615
R1282 VTAIL.n200 VTAIL.n169 104.615
R1283 VTAIL.n193 VTAIL.n169 104.615
R1284 VTAIL.n193 VTAIL.n192 104.615
R1285 VTAIL.n192 VTAIL.n174 104.615
R1286 VTAIL.n185 VTAIL.n174 104.615
R1287 VTAIL.n185 VTAIL.n184 104.615
R1288 VTAIL.n184 VTAIL.n178 104.615
R1289 VTAIL.t6 VTAIL.n393 52.3082
R1290 VTAIL.t4 VTAIL.n15 52.3082
R1291 VTAIL.t0 VTAIL.n69 52.3082
R1292 VTAIL.t2 VTAIL.n123 52.3082
R1293 VTAIL.t1 VTAIL.n340 52.3082
R1294 VTAIL.t3 VTAIL.n286 52.3082
R1295 VTAIL.t5 VTAIL.n232 52.3082
R1296 VTAIL.t7 VTAIL.n178 52.3082
R1297 VTAIL.n431 VTAIL.n430 33.7369
R1298 VTAIL.n53 VTAIL.n52 33.7369
R1299 VTAIL.n107 VTAIL.n106 33.7369
R1300 VTAIL.n161 VTAIL.n160 33.7369
R1301 VTAIL.n377 VTAIL.n376 33.7369
R1302 VTAIL.n323 VTAIL.n322 33.7369
R1303 VTAIL.n269 VTAIL.n268 33.7369
R1304 VTAIL.n215 VTAIL.n214 33.7369
R1305 VTAIL.n431 VTAIL.n377 22.2634
R1306 VTAIL.n215 VTAIL.n161 22.2634
R1307 VTAIL.n419 VTAIL.n384 13.1884
R1308 VTAIL.n41 VTAIL.n6 13.1884
R1309 VTAIL.n95 VTAIL.n60 13.1884
R1310 VTAIL.n149 VTAIL.n114 13.1884
R1311 VTAIL.n365 VTAIL.n330 13.1884
R1312 VTAIL.n311 VTAIL.n276 13.1884
R1313 VTAIL.n257 VTAIL.n222 13.1884
R1314 VTAIL.n203 VTAIL.n168 13.1884
R1315 VTAIL.n415 VTAIL.n414 12.8005
R1316 VTAIL.n420 VTAIL.n382 12.8005
R1317 VTAIL.n37 VTAIL.n36 12.8005
R1318 VTAIL.n42 VTAIL.n4 12.8005
R1319 VTAIL.n91 VTAIL.n90 12.8005
R1320 VTAIL.n96 VTAIL.n58 12.8005
R1321 VTAIL.n145 VTAIL.n144 12.8005
R1322 VTAIL.n150 VTAIL.n112 12.8005
R1323 VTAIL.n366 VTAIL.n328 12.8005
R1324 VTAIL.n361 VTAIL.n332 12.8005
R1325 VTAIL.n312 VTAIL.n274 12.8005
R1326 VTAIL.n307 VTAIL.n278 12.8005
R1327 VTAIL.n258 VTAIL.n220 12.8005
R1328 VTAIL.n253 VTAIL.n224 12.8005
R1329 VTAIL.n204 VTAIL.n166 12.8005
R1330 VTAIL.n199 VTAIL.n170 12.8005
R1331 VTAIL.n413 VTAIL.n386 12.0247
R1332 VTAIL.n424 VTAIL.n423 12.0247
R1333 VTAIL.n35 VTAIL.n8 12.0247
R1334 VTAIL.n46 VTAIL.n45 12.0247
R1335 VTAIL.n89 VTAIL.n62 12.0247
R1336 VTAIL.n100 VTAIL.n99 12.0247
R1337 VTAIL.n143 VTAIL.n116 12.0247
R1338 VTAIL.n154 VTAIL.n153 12.0247
R1339 VTAIL.n370 VTAIL.n369 12.0247
R1340 VTAIL.n360 VTAIL.n333 12.0247
R1341 VTAIL.n316 VTAIL.n315 12.0247
R1342 VTAIL.n306 VTAIL.n279 12.0247
R1343 VTAIL.n262 VTAIL.n261 12.0247
R1344 VTAIL.n252 VTAIL.n225 12.0247
R1345 VTAIL.n208 VTAIL.n207 12.0247
R1346 VTAIL.n198 VTAIL.n171 12.0247
R1347 VTAIL.n410 VTAIL.n409 11.249
R1348 VTAIL.n427 VTAIL.n380 11.249
R1349 VTAIL.n32 VTAIL.n31 11.249
R1350 VTAIL.n49 VTAIL.n2 11.249
R1351 VTAIL.n86 VTAIL.n85 11.249
R1352 VTAIL.n103 VTAIL.n56 11.249
R1353 VTAIL.n140 VTAIL.n139 11.249
R1354 VTAIL.n157 VTAIL.n110 11.249
R1355 VTAIL.n373 VTAIL.n326 11.249
R1356 VTAIL.n357 VTAIL.n356 11.249
R1357 VTAIL.n319 VTAIL.n272 11.249
R1358 VTAIL.n303 VTAIL.n302 11.249
R1359 VTAIL.n265 VTAIL.n218 11.249
R1360 VTAIL.n249 VTAIL.n248 11.249
R1361 VTAIL.n211 VTAIL.n164 11.249
R1362 VTAIL.n195 VTAIL.n194 11.249
R1363 VTAIL.n406 VTAIL.n388 10.4732
R1364 VTAIL.n428 VTAIL.n378 10.4732
R1365 VTAIL.n28 VTAIL.n10 10.4732
R1366 VTAIL.n50 VTAIL.n0 10.4732
R1367 VTAIL.n82 VTAIL.n64 10.4732
R1368 VTAIL.n104 VTAIL.n54 10.4732
R1369 VTAIL.n136 VTAIL.n118 10.4732
R1370 VTAIL.n158 VTAIL.n108 10.4732
R1371 VTAIL.n374 VTAIL.n324 10.4732
R1372 VTAIL.n353 VTAIL.n335 10.4732
R1373 VTAIL.n320 VTAIL.n270 10.4732
R1374 VTAIL.n299 VTAIL.n281 10.4732
R1375 VTAIL.n266 VTAIL.n216 10.4732
R1376 VTAIL.n245 VTAIL.n227 10.4732
R1377 VTAIL.n212 VTAIL.n162 10.4732
R1378 VTAIL.n191 VTAIL.n173 10.4732
R1379 VTAIL.n395 VTAIL.n394 10.2747
R1380 VTAIL.n17 VTAIL.n16 10.2747
R1381 VTAIL.n71 VTAIL.n70 10.2747
R1382 VTAIL.n125 VTAIL.n124 10.2747
R1383 VTAIL.n342 VTAIL.n341 10.2747
R1384 VTAIL.n288 VTAIL.n287 10.2747
R1385 VTAIL.n234 VTAIL.n233 10.2747
R1386 VTAIL.n180 VTAIL.n179 10.2747
R1387 VTAIL.n405 VTAIL.n390 9.69747
R1388 VTAIL.n27 VTAIL.n12 9.69747
R1389 VTAIL.n81 VTAIL.n66 9.69747
R1390 VTAIL.n135 VTAIL.n120 9.69747
R1391 VTAIL.n352 VTAIL.n337 9.69747
R1392 VTAIL.n298 VTAIL.n283 9.69747
R1393 VTAIL.n244 VTAIL.n229 9.69747
R1394 VTAIL.n190 VTAIL.n175 9.69747
R1395 VTAIL.n430 VTAIL.n429 9.45567
R1396 VTAIL.n52 VTAIL.n51 9.45567
R1397 VTAIL.n106 VTAIL.n105 9.45567
R1398 VTAIL.n160 VTAIL.n159 9.45567
R1399 VTAIL.n376 VTAIL.n375 9.45567
R1400 VTAIL.n322 VTAIL.n321 9.45567
R1401 VTAIL.n268 VTAIL.n267 9.45567
R1402 VTAIL.n214 VTAIL.n213 9.45567
R1403 VTAIL.n429 VTAIL.n428 9.3005
R1404 VTAIL.n380 VTAIL.n379 9.3005
R1405 VTAIL.n423 VTAIL.n422 9.3005
R1406 VTAIL.n421 VTAIL.n420 9.3005
R1407 VTAIL.n397 VTAIL.n396 9.3005
R1408 VTAIL.n392 VTAIL.n391 9.3005
R1409 VTAIL.n403 VTAIL.n402 9.3005
R1410 VTAIL.n405 VTAIL.n404 9.3005
R1411 VTAIL.n388 VTAIL.n387 9.3005
R1412 VTAIL.n411 VTAIL.n410 9.3005
R1413 VTAIL.n413 VTAIL.n412 9.3005
R1414 VTAIL.n414 VTAIL.n383 9.3005
R1415 VTAIL.n51 VTAIL.n50 9.3005
R1416 VTAIL.n2 VTAIL.n1 9.3005
R1417 VTAIL.n45 VTAIL.n44 9.3005
R1418 VTAIL.n43 VTAIL.n42 9.3005
R1419 VTAIL.n19 VTAIL.n18 9.3005
R1420 VTAIL.n14 VTAIL.n13 9.3005
R1421 VTAIL.n25 VTAIL.n24 9.3005
R1422 VTAIL.n27 VTAIL.n26 9.3005
R1423 VTAIL.n10 VTAIL.n9 9.3005
R1424 VTAIL.n33 VTAIL.n32 9.3005
R1425 VTAIL.n35 VTAIL.n34 9.3005
R1426 VTAIL.n36 VTAIL.n5 9.3005
R1427 VTAIL.n105 VTAIL.n104 9.3005
R1428 VTAIL.n56 VTAIL.n55 9.3005
R1429 VTAIL.n99 VTAIL.n98 9.3005
R1430 VTAIL.n97 VTAIL.n96 9.3005
R1431 VTAIL.n73 VTAIL.n72 9.3005
R1432 VTAIL.n68 VTAIL.n67 9.3005
R1433 VTAIL.n79 VTAIL.n78 9.3005
R1434 VTAIL.n81 VTAIL.n80 9.3005
R1435 VTAIL.n64 VTAIL.n63 9.3005
R1436 VTAIL.n87 VTAIL.n86 9.3005
R1437 VTAIL.n89 VTAIL.n88 9.3005
R1438 VTAIL.n90 VTAIL.n59 9.3005
R1439 VTAIL.n159 VTAIL.n158 9.3005
R1440 VTAIL.n110 VTAIL.n109 9.3005
R1441 VTAIL.n153 VTAIL.n152 9.3005
R1442 VTAIL.n151 VTAIL.n150 9.3005
R1443 VTAIL.n127 VTAIL.n126 9.3005
R1444 VTAIL.n122 VTAIL.n121 9.3005
R1445 VTAIL.n133 VTAIL.n132 9.3005
R1446 VTAIL.n135 VTAIL.n134 9.3005
R1447 VTAIL.n118 VTAIL.n117 9.3005
R1448 VTAIL.n141 VTAIL.n140 9.3005
R1449 VTAIL.n143 VTAIL.n142 9.3005
R1450 VTAIL.n144 VTAIL.n113 9.3005
R1451 VTAIL.n344 VTAIL.n343 9.3005
R1452 VTAIL.n339 VTAIL.n338 9.3005
R1453 VTAIL.n350 VTAIL.n349 9.3005
R1454 VTAIL.n352 VTAIL.n351 9.3005
R1455 VTAIL.n335 VTAIL.n334 9.3005
R1456 VTAIL.n358 VTAIL.n357 9.3005
R1457 VTAIL.n360 VTAIL.n359 9.3005
R1458 VTAIL.n332 VTAIL.n329 9.3005
R1459 VTAIL.n375 VTAIL.n374 9.3005
R1460 VTAIL.n326 VTAIL.n325 9.3005
R1461 VTAIL.n369 VTAIL.n368 9.3005
R1462 VTAIL.n367 VTAIL.n366 9.3005
R1463 VTAIL.n290 VTAIL.n289 9.3005
R1464 VTAIL.n285 VTAIL.n284 9.3005
R1465 VTAIL.n296 VTAIL.n295 9.3005
R1466 VTAIL.n298 VTAIL.n297 9.3005
R1467 VTAIL.n281 VTAIL.n280 9.3005
R1468 VTAIL.n304 VTAIL.n303 9.3005
R1469 VTAIL.n306 VTAIL.n305 9.3005
R1470 VTAIL.n278 VTAIL.n275 9.3005
R1471 VTAIL.n321 VTAIL.n320 9.3005
R1472 VTAIL.n272 VTAIL.n271 9.3005
R1473 VTAIL.n315 VTAIL.n314 9.3005
R1474 VTAIL.n313 VTAIL.n312 9.3005
R1475 VTAIL.n236 VTAIL.n235 9.3005
R1476 VTAIL.n231 VTAIL.n230 9.3005
R1477 VTAIL.n242 VTAIL.n241 9.3005
R1478 VTAIL.n244 VTAIL.n243 9.3005
R1479 VTAIL.n227 VTAIL.n226 9.3005
R1480 VTAIL.n250 VTAIL.n249 9.3005
R1481 VTAIL.n252 VTAIL.n251 9.3005
R1482 VTAIL.n224 VTAIL.n221 9.3005
R1483 VTAIL.n267 VTAIL.n266 9.3005
R1484 VTAIL.n218 VTAIL.n217 9.3005
R1485 VTAIL.n261 VTAIL.n260 9.3005
R1486 VTAIL.n259 VTAIL.n258 9.3005
R1487 VTAIL.n182 VTAIL.n181 9.3005
R1488 VTAIL.n177 VTAIL.n176 9.3005
R1489 VTAIL.n188 VTAIL.n187 9.3005
R1490 VTAIL.n190 VTAIL.n189 9.3005
R1491 VTAIL.n173 VTAIL.n172 9.3005
R1492 VTAIL.n196 VTAIL.n195 9.3005
R1493 VTAIL.n198 VTAIL.n197 9.3005
R1494 VTAIL.n170 VTAIL.n167 9.3005
R1495 VTAIL.n213 VTAIL.n212 9.3005
R1496 VTAIL.n164 VTAIL.n163 9.3005
R1497 VTAIL.n207 VTAIL.n206 9.3005
R1498 VTAIL.n205 VTAIL.n204 9.3005
R1499 VTAIL.n402 VTAIL.n401 8.92171
R1500 VTAIL.n24 VTAIL.n23 8.92171
R1501 VTAIL.n78 VTAIL.n77 8.92171
R1502 VTAIL.n132 VTAIL.n131 8.92171
R1503 VTAIL.n349 VTAIL.n348 8.92171
R1504 VTAIL.n295 VTAIL.n294 8.92171
R1505 VTAIL.n241 VTAIL.n240 8.92171
R1506 VTAIL.n187 VTAIL.n186 8.92171
R1507 VTAIL.n398 VTAIL.n392 8.14595
R1508 VTAIL.n20 VTAIL.n14 8.14595
R1509 VTAIL.n74 VTAIL.n68 8.14595
R1510 VTAIL.n128 VTAIL.n122 8.14595
R1511 VTAIL.n345 VTAIL.n339 8.14595
R1512 VTAIL.n291 VTAIL.n285 8.14595
R1513 VTAIL.n237 VTAIL.n231 8.14595
R1514 VTAIL.n183 VTAIL.n177 8.14595
R1515 VTAIL.n397 VTAIL.n394 7.3702
R1516 VTAIL.n19 VTAIL.n16 7.3702
R1517 VTAIL.n73 VTAIL.n70 7.3702
R1518 VTAIL.n127 VTAIL.n124 7.3702
R1519 VTAIL.n344 VTAIL.n341 7.3702
R1520 VTAIL.n290 VTAIL.n287 7.3702
R1521 VTAIL.n236 VTAIL.n233 7.3702
R1522 VTAIL.n182 VTAIL.n179 7.3702
R1523 VTAIL.n398 VTAIL.n397 5.81868
R1524 VTAIL.n20 VTAIL.n19 5.81868
R1525 VTAIL.n74 VTAIL.n73 5.81868
R1526 VTAIL.n128 VTAIL.n127 5.81868
R1527 VTAIL.n345 VTAIL.n344 5.81868
R1528 VTAIL.n291 VTAIL.n290 5.81868
R1529 VTAIL.n237 VTAIL.n236 5.81868
R1530 VTAIL.n183 VTAIL.n182 5.81868
R1531 VTAIL.n401 VTAIL.n392 5.04292
R1532 VTAIL.n23 VTAIL.n14 5.04292
R1533 VTAIL.n77 VTAIL.n68 5.04292
R1534 VTAIL.n131 VTAIL.n122 5.04292
R1535 VTAIL.n348 VTAIL.n339 5.04292
R1536 VTAIL.n294 VTAIL.n285 5.04292
R1537 VTAIL.n240 VTAIL.n231 5.04292
R1538 VTAIL.n186 VTAIL.n177 5.04292
R1539 VTAIL.n402 VTAIL.n390 4.26717
R1540 VTAIL.n24 VTAIL.n12 4.26717
R1541 VTAIL.n78 VTAIL.n66 4.26717
R1542 VTAIL.n132 VTAIL.n120 4.26717
R1543 VTAIL.n349 VTAIL.n337 4.26717
R1544 VTAIL.n295 VTAIL.n283 4.26717
R1545 VTAIL.n241 VTAIL.n229 4.26717
R1546 VTAIL.n187 VTAIL.n175 4.26717
R1547 VTAIL.n406 VTAIL.n405 3.49141
R1548 VTAIL.n430 VTAIL.n378 3.49141
R1549 VTAIL.n28 VTAIL.n27 3.49141
R1550 VTAIL.n52 VTAIL.n0 3.49141
R1551 VTAIL.n82 VTAIL.n81 3.49141
R1552 VTAIL.n106 VTAIL.n54 3.49141
R1553 VTAIL.n136 VTAIL.n135 3.49141
R1554 VTAIL.n160 VTAIL.n108 3.49141
R1555 VTAIL.n376 VTAIL.n324 3.49141
R1556 VTAIL.n353 VTAIL.n352 3.49141
R1557 VTAIL.n322 VTAIL.n270 3.49141
R1558 VTAIL.n299 VTAIL.n298 3.49141
R1559 VTAIL.n268 VTAIL.n216 3.49141
R1560 VTAIL.n245 VTAIL.n244 3.49141
R1561 VTAIL.n214 VTAIL.n162 3.49141
R1562 VTAIL.n191 VTAIL.n190 3.49141
R1563 VTAIL.n396 VTAIL.n395 2.84303
R1564 VTAIL.n18 VTAIL.n17 2.84303
R1565 VTAIL.n72 VTAIL.n71 2.84303
R1566 VTAIL.n126 VTAIL.n125 2.84303
R1567 VTAIL.n343 VTAIL.n342 2.84303
R1568 VTAIL.n289 VTAIL.n288 2.84303
R1569 VTAIL.n235 VTAIL.n234 2.84303
R1570 VTAIL.n181 VTAIL.n180 2.84303
R1571 VTAIL.n409 VTAIL.n388 2.71565
R1572 VTAIL.n428 VTAIL.n427 2.71565
R1573 VTAIL.n31 VTAIL.n10 2.71565
R1574 VTAIL.n50 VTAIL.n49 2.71565
R1575 VTAIL.n85 VTAIL.n64 2.71565
R1576 VTAIL.n104 VTAIL.n103 2.71565
R1577 VTAIL.n139 VTAIL.n118 2.71565
R1578 VTAIL.n158 VTAIL.n157 2.71565
R1579 VTAIL.n374 VTAIL.n373 2.71565
R1580 VTAIL.n356 VTAIL.n335 2.71565
R1581 VTAIL.n320 VTAIL.n319 2.71565
R1582 VTAIL.n302 VTAIL.n281 2.71565
R1583 VTAIL.n266 VTAIL.n265 2.71565
R1584 VTAIL.n248 VTAIL.n227 2.71565
R1585 VTAIL.n212 VTAIL.n211 2.71565
R1586 VTAIL.n194 VTAIL.n173 2.71565
R1587 VTAIL.n410 VTAIL.n386 1.93989
R1588 VTAIL.n424 VTAIL.n380 1.93989
R1589 VTAIL.n32 VTAIL.n8 1.93989
R1590 VTAIL.n46 VTAIL.n2 1.93989
R1591 VTAIL.n86 VTAIL.n62 1.93989
R1592 VTAIL.n100 VTAIL.n56 1.93989
R1593 VTAIL.n140 VTAIL.n116 1.93989
R1594 VTAIL.n154 VTAIL.n110 1.93989
R1595 VTAIL.n370 VTAIL.n326 1.93989
R1596 VTAIL.n357 VTAIL.n333 1.93989
R1597 VTAIL.n316 VTAIL.n272 1.93989
R1598 VTAIL.n303 VTAIL.n279 1.93989
R1599 VTAIL.n262 VTAIL.n218 1.93989
R1600 VTAIL.n249 VTAIL.n225 1.93989
R1601 VTAIL.n208 VTAIL.n164 1.93989
R1602 VTAIL.n195 VTAIL.n171 1.93989
R1603 VTAIL.n269 VTAIL.n215 1.24188
R1604 VTAIL.n377 VTAIL.n323 1.24188
R1605 VTAIL.n161 VTAIL.n107 1.24188
R1606 VTAIL.n415 VTAIL.n413 1.16414
R1607 VTAIL.n423 VTAIL.n382 1.16414
R1608 VTAIL.n37 VTAIL.n35 1.16414
R1609 VTAIL.n45 VTAIL.n4 1.16414
R1610 VTAIL.n91 VTAIL.n89 1.16414
R1611 VTAIL.n99 VTAIL.n58 1.16414
R1612 VTAIL.n145 VTAIL.n143 1.16414
R1613 VTAIL.n153 VTAIL.n112 1.16414
R1614 VTAIL.n369 VTAIL.n328 1.16414
R1615 VTAIL.n361 VTAIL.n360 1.16414
R1616 VTAIL.n315 VTAIL.n274 1.16414
R1617 VTAIL.n307 VTAIL.n306 1.16414
R1618 VTAIL.n261 VTAIL.n220 1.16414
R1619 VTAIL.n253 VTAIL.n252 1.16414
R1620 VTAIL.n207 VTAIL.n166 1.16414
R1621 VTAIL.n199 VTAIL.n198 1.16414
R1622 VTAIL VTAIL.n53 0.679379
R1623 VTAIL VTAIL.n431 0.563
R1624 VTAIL.n323 VTAIL.n269 0.470328
R1625 VTAIL.n107 VTAIL.n53 0.470328
R1626 VTAIL.n414 VTAIL.n384 0.388379
R1627 VTAIL.n420 VTAIL.n419 0.388379
R1628 VTAIL.n36 VTAIL.n6 0.388379
R1629 VTAIL.n42 VTAIL.n41 0.388379
R1630 VTAIL.n90 VTAIL.n60 0.388379
R1631 VTAIL.n96 VTAIL.n95 0.388379
R1632 VTAIL.n144 VTAIL.n114 0.388379
R1633 VTAIL.n150 VTAIL.n149 0.388379
R1634 VTAIL.n366 VTAIL.n365 0.388379
R1635 VTAIL.n332 VTAIL.n330 0.388379
R1636 VTAIL.n312 VTAIL.n311 0.388379
R1637 VTAIL.n278 VTAIL.n276 0.388379
R1638 VTAIL.n258 VTAIL.n257 0.388379
R1639 VTAIL.n224 VTAIL.n222 0.388379
R1640 VTAIL.n204 VTAIL.n203 0.388379
R1641 VTAIL.n170 VTAIL.n168 0.388379
R1642 VTAIL.n396 VTAIL.n391 0.155672
R1643 VTAIL.n403 VTAIL.n391 0.155672
R1644 VTAIL.n404 VTAIL.n403 0.155672
R1645 VTAIL.n404 VTAIL.n387 0.155672
R1646 VTAIL.n411 VTAIL.n387 0.155672
R1647 VTAIL.n412 VTAIL.n411 0.155672
R1648 VTAIL.n412 VTAIL.n383 0.155672
R1649 VTAIL.n421 VTAIL.n383 0.155672
R1650 VTAIL.n422 VTAIL.n421 0.155672
R1651 VTAIL.n422 VTAIL.n379 0.155672
R1652 VTAIL.n429 VTAIL.n379 0.155672
R1653 VTAIL.n18 VTAIL.n13 0.155672
R1654 VTAIL.n25 VTAIL.n13 0.155672
R1655 VTAIL.n26 VTAIL.n25 0.155672
R1656 VTAIL.n26 VTAIL.n9 0.155672
R1657 VTAIL.n33 VTAIL.n9 0.155672
R1658 VTAIL.n34 VTAIL.n33 0.155672
R1659 VTAIL.n34 VTAIL.n5 0.155672
R1660 VTAIL.n43 VTAIL.n5 0.155672
R1661 VTAIL.n44 VTAIL.n43 0.155672
R1662 VTAIL.n44 VTAIL.n1 0.155672
R1663 VTAIL.n51 VTAIL.n1 0.155672
R1664 VTAIL.n72 VTAIL.n67 0.155672
R1665 VTAIL.n79 VTAIL.n67 0.155672
R1666 VTAIL.n80 VTAIL.n79 0.155672
R1667 VTAIL.n80 VTAIL.n63 0.155672
R1668 VTAIL.n87 VTAIL.n63 0.155672
R1669 VTAIL.n88 VTAIL.n87 0.155672
R1670 VTAIL.n88 VTAIL.n59 0.155672
R1671 VTAIL.n97 VTAIL.n59 0.155672
R1672 VTAIL.n98 VTAIL.n97 0.155672
R1673 VTAIL.n98 VTAIL.n55 0.155672
R1674 VTAIL.n105 VTAIL.n55 0.155672
R1675 VTAIL.n126 VTAIL.n121 0.155672
R1676 VTAIL.n133 VTAIL.n121 0.155672
R1677 VTAIL.n134 VTAIL.n133 0.155672
R1678 VTAIL.n134 VTAIL.n117 0.155672
R1679 VTAIL.n141 VTAIL.n117 0.155672
R1680 VTAIL.n142 VTAIL.n141 0.155672
R1681 VTAIL.n142 VTAIL.n113 0.155672
R1682 VTAIL.n151 VTAIL.n113 0.155672
R1683 VTAIL.n152 VTAIL.n151 0.155672
R1684 VTAIL.n152 VTAIL.n109 0.155672
R1685 VTAIL.n159 VTAIL.n109 0.155672
R1686 VTAIL.n375 VTAIL.n325 0.155672
R1687 VTAIL.n368 VTAIL.n325 0.155672
R1688 VTAIL.n368 VTAIL.n367 0.155672
R1689 VTAIL.n367 VTAIL.n329 0.155672
R1690 VTAIL.n359 VTAIL.n329 0.155672
R1691 VTAIL.n359 VTAIL.n358 0.155672
R1692 VTAIL.n358 VTAIL.n334 0.155672
R1693 VTAIL.n351 VTAIL.n334 0.155672
R1694 VTAIL.n351 VTAIL.n350 0.155672
R1695 VTAIL.n350 VTAIL.n338 0.155672
R1696 VTAIL.n343 VTAIL.n338 0.155672
R1697 VTAIL.n321 VTAIL.n271 0.155672
R1698 VTAIL.n314 VTAIL.n271 0.155672
R1699 VTAIL.n314 VTAIL.n313 0.155672
R1700 VTAIL.n313 VTAIL.n275 0.155672
R1701 VTAIL.n305 VTAIL.n275 0.155672
R1702 VTAIL.n305 VTAIL.n304 0.155672
R1703 VTAIL.n304 VTAIL.n280 0.155672
R1704 VTAIL.n297 VTAIL.n280 0.155672
R1705 VTAIL.n297 VTAIL.n296 0.155672
R1706 VTAIL.n296 VTAIL.n284 0.155672
R1707 VTAIL.n289 VTAIL.n284 0.155672
R1708 VTAIL.n267 VTAIL.n217 0.155672
R1709 VTAIL.n260 VTAIL.n217 0.155672
R1710 VTAIL.n260 VTAIL.n259 0.155672
R1711 VTAIL.n259 VTAIL.n221 0.155672
R1712 VTAIL.n251 VTAIL.n221 0.155672
R1713 VTAIL.n251 VTAIL.n250 0.155672
R1714 VTAIL.n250 VTAIL.n226 0.155672
R1715 VTAIL.n243 VTAIL.n226 0.155672
R1716 VTAIL.n243 VTAIL.n242 0.155672
R1717 VTAIL.n242 VTAIL.n230 0.155672
R1718 VTAIL.n235 VTAIL.n230 0.155672
R1719 VTAIL.n213 VTAIL.n163 0.155672
R1720 VTAIL.n206 VTAIL.n163 0.155672
R1721 VTAIL.n206 VTAIL.n205 0.155672
R1722 VTAIL.n205 VTAIL.n167 0.155672
R1723 VTAIL.n197 VTAIL.n167 0.155672
R1724 VTAIL.n197 VTAIL.n196 0.155672
R1725 VTAIL.n196 VTAIL.n172 0.155672
R1726 VTAIL.n189 VTAIL.n172 0.155672
R1727 VTAIL.n189 VTAIL.n188 0.155672
R1728 VTAIL.n188 VTAIL.n176 0.155672
R1729 VTAIL.n181 VTAIL.n176 0.155672
R1730 VDD2.n2 VDD2.n0 100.285
R1731 VDD2.n2 VDD2.n1 64.1917
R1732 VDD2.n1 VDD2.t1 1.97261
R1733 VDD2.n1 VDD2.t2 1.97261
R1734 VDD2.n0 VDD2.t0 1.97261
R1735 VDD2.n0 VDD2.t3 1.97261
R1736 VDD2 VDD2.n2 0.0586897
R1737 VP.n0 VP.t2 271.983
R1738 VP.n0 VP.t1 271.896
R1739 VP.n2 VP.t0 253.376
R1740 VP.n3 VP.t3 253.376
R1741 VP.n4 VP.n3 80.6037
R1742 VP.n2 VP.n1 80.6037
R1743 VP.n1 VP.n0 71.5941
R1744 VP.n3 VP.n2 48.2005
R1745 VP.n4 VP.n1 0.380177
R1746 VP VP.n4 0.146778
R1747 VDD1 VDD1.n1 100.811
R1748 VDD1 VDD1.n0 64.2499
R1749 VDD1.n0 VDD1.t1 1.97261
R1750 VDD1.n0 VDD1.t2 1.97261
R1751 VDD1.n1 VDD1.t3 1.97261
R1752 VDD1.n1 VDD1.t0 1.97261
C0 VDD1 VTAIL 5.19995f
C1 VDD1 VP 3.37683f
C2 VTAIL VN 2.9901f
C3 VP VN 4.74863f
C4 VDD1 VDD2 0.664848f
C5 VDD2 VN 3.22535f
C6 VTAIL VP 3.00421f
C7 VTAIL VDD2 5.24416f
C8 VP VDD2 0.29994f
C9 VDD1 VN 0.148099f
C10 VDD2 B 2.780117f
C11 VDD1 B 6.25601f
C12 VTAIL B 7.979419f
C13 VN B 8.250331f
C14 VP B 5.645488f
C15 VDD1.t1 B 0.215284f
C16 VDD1.t2 B 0.215284f
C17 VDD1.n0 B 1.89787f
C18 VDD1.t3 B 0.215284f
C19 VDD1.t0 B 0.215284f
C20 VDD1.n1 B 2.4476f
C21 VP.t1 B 1.37692f
C22 VP.t2 B 1.37712f
C23 VP.n0 B 2.01397f
C24 VP.n1 B 2.45915f
C25 VP.t0 B 1.33962f
C26 VP.n2 B 0.547673f
C27 VP.t3 B 1.33962f
C28 VP.n3 B 0.547673f
C29 VP.n4 B 0.053396f
C30 VDD2.t0 B 0.212757f
C31 VDD2.t3 B 0.212757f
C32 VDD2.n0 B 2.39431f
C33 VDD2.t1 B 0.212757f
C34 VDD2.t2 B 0.212757f
C35 VDD2.n1 B 1.87528f
C36 VDD2.n2 B 3.16635f
C37 VTAIL.n0 B 0.022464f
C38 VTAIL.n1 B 0.016295f
C39 VTAIL.n2 B 0.008756f
C40 VTAIL.n3 B 0.020696f
C41 VTAIL.n4 B 0.009271f
C42 VTAIL.n5 B 0.016295f
C43 VTAIL.n6 B 0.009014f
C44 VTAIL.n7 B 0.020696f
C45 VTAIL.n8 B 0.009271f
C46 VTAIL.n9 B 0.016295f
C47 VTAIL.n10 B 0.008756f
C48 VTAIL.n11 B 0.020696f
C49 VTAIL.n12 B 0.009271f
C50 VTAIL.n13 B 0.016295f
C51 VTAIL.n14 B 0.008756f
C52 VTAIL.n15 B 0.015522f
C53 VTAIL.n16 B 0.01463f
C54 VTAIL.t4 B 0.034784f
C55 VTAIL.n17 B 0.105223f
C56 VTAIL.n18 B 0.679975f
C57 VTAIL.n19 B 0.008756f
C58 VTAIL.n20 B 0.009271f
C59 VTAIL.n21 B 0.020696f
C60 VTAIL.n22 B 0.020696f
C61 VTAIL.n23 B 0.009271f
C62 VTAIL.n24 B 0.008756f
C63 VTAIL.n25 B 0.016295f
C64 VTAIL.n26 B 0.016295f
C65 VTAIL.n27 B 0.008756f
C66 VTAIL.n28 B 0.009271f
C67 VTAIL.n29 B 0.020696f
C68 VTAIL.n30 B 0.020696f
C69 VTAIL.n31 B 0.009271f
C70 VTAIL.n32 B 0.008756f
C71 VTAIL.n33 B 0.016295f
C72 VTAIL.n34 B 0.016295f
C73 VTAIL.n35 B 0.008756f
C74 VTAIL.n36 B 0.008756f
C75 VTAIL.n37 B 0.009271f
C76 VTAIL.n38 B 0.020696f
C77 VTAIL.n39 B 0.020696f
C78 VTAIL.n40 B 0.020696f
C79 VTAIL.n41 B 0.009014f
C80 VTAIL.n42 B 0.008756f
C81 VTAIL.n43 B 0.016295f
C82 VTAIL.n44 B 0.016295f
C83 VTAIL.n45 B 0.008756f
C84 VTAIL.n46 B 0.009271f
C85 VTAIL.n47 B 0.020696f
C86 VTAIL.n48 B 0.044026f
C87 VTAIL.n49 B 0.009271f
C88 VTAIL.n50 B 0.008756f
C89 VTAIL.n51 B 0.039445f
C90 VTAIL.n52 B 0.024608f
C91 VTAIL.n53 B 0.075235f
C92 VTAIL.n54 B 0.022464f
C93 VTAIL.n55 B 0.016295f
C94 VTAIL.n56 B 0.008756f
C95 VTAIL.n57 B 0.020696f
C96 VTAIL.n58 B 0.009271f
C97 VTAIL.n59 B 0.016295f
C98 VTAIL.n60 B 0.009014f
C99 VTAIL.n61 B 0.020696f
C100 VTAIL.n62 B 0.009271f
C101 VTAIL.n63 B 0.016295f
C102 VTAIL.n64 B 0.008756f
C103 VTAIL.n65 B 0.020696f
C104 VTAIL.n66 B 0.009271f
C105 VTAIL.n67 B 0.016295f
C106 VTAIL.n68 B 0.008756f
C107 VTAIL.n69 B 0.015522f
C108 VTAIL.n70 B 0.01463f
C109 VTAIL.t0 B 0.034784f
C110 VTAIL.n71 B 0.105223f
C111 VTAIL.n72 B 0.679975f
C112 VTAIL.n73 B 0.008756f
C113 VTAIL.n74 B 0.009271f
C114 VTAIL.n75 B 0.020696f
C115 VTAIL.n76 B 0.020696f
C116 VTAIL.n77 B 0.009271f
C117 VTAIL.n78 B 0.008756f
C118 VTAIL.n79 B 0.016295f
C119 VTAIL.n80 B 0.016295f
C120 VTAIL.n81 B 0.008756f
C121 VTAIL.n82 B 0.009271f
C122 VTAIL.n83 B 0.020696f
C123 VTAIL.n84 B 0.020696f
C124 VTAIL.n85 B 0.009271f
C125 VTAIL.n86 B 0.008756f
C126 VTAIL.n87 B 0.016295f
C127 VTAIL.n88 B 0.016295f
C128 VTAIL.n89 B 0.008756f
C129 VTAIL.n90 B 0.008756f
C130 VTAIL.n91 B 0.009271f
C131 VTAIL.n92 B 0.020696f
C132 VTAIL.n93 B 0.020696f
C133 VTAIL.n94 B 0.020696f
C134 VTAIL.n95 B 0.009014f
C135 VTAIL.n96 B 0.008756f
C136 VTAIL.n97 B 0.016295f
C137 VTAIL.n98 B 0.016295f
C138 VTAIL.n99 B 0.008756f
C139 VTAIL.n100 B 0.009271f
C140 VTAIL.n101 B 0.020696f
C141 VTAIL.n102 B 0.044026f
C142 VTAIL.n103 B 0.009271f
C143 VTAIL.n104 B 0.008756f
C144 VTAIL.n105 B 0.039445f
C145 VTAIL.n106 B 0.024608f
C146 VTAIL.n107 B 0.104769f
C147 VTAIL.n108 B 0.022464f
C148 VTAIL.n109 B 0.016295f
C149 VTAIL.n110 B 0.008756f
C150 VTAIL.n111 B 0.020696f
C151 VTAIL.n112 B 0.009271f
C152 VTAIL.n113 B 0.016295f
C153 VTAIL.n114 B 0.009014f
C154 VTAIL.n115 B 0.020696f
C155 VTAIL.n116 B 0.009271f
C156 VTAIL.n117 B 0.016295f
C157 VTAIL.n118 B 0.008756f
C158 VTAIL.n119 B 0.020696f
C159 VTAIL.n120 B 0.009271f
C160 VTAIL.n121 B 0.016295f
C161 VTAIL.n122 B 0.008756f
C162 VTAIL.n123 B 0.015522f
C163 VTAIL.n124 B 0.01463f
C164 VTAIL.t2 B 0.034784f
C165 VTAIL.n125 B 0.105223f
C166 VTAIL.n126 B 0.679975f
C167 VTAIL.n127 B 0.008756f
C168 VTAIL.n128 B 0.009271f
C169 VTAIL.n129 B 0.020696f
C170 VTAIL.n130 B 0.020696f
C171 VTAIL.n131 B 0.009271f
C172 VTAIL.n132 B 0.008756f
C173 VTAIL.n133 B 0.016295f
C174 VTAIL.n134 B 0.016295f
C175 VTAIL.n135 B 0.008756f
C176 VTAIL.n136 B 0.009271f
C177 VTAIL.n137 B 0.020696f
C178 VTAIL.n138 B 0.020696f
C179 VTAIL.n139 B 0.009271f
C180 VTAIL.n140 B 0.008756f
C181 VTAIL.n141 B 0.016295f
C182 VTAIL.n142 B 0.016295f
C183 VTAIL.n143 B 0.008756f
C184 VTAIL.n144 B 0.008756f
C185 VTAIL.n145 B 0.009271f
C186 VTAIL.n146 B 0.020696f
C187 VTAIL.n147 B 0.020696f
C188 VTAIL.n148 B 0.020696f
C189 VTAIL.n149 B 0.009014f
C190 VTAIL.n150 B 0.008756f
C191 VTAIL.n151 B 0.016295f
C192 VTAIL.n152 B 0.016295f
C193 VTAIL.n153 B 0.008756f
C194 VTAIL.n154 B 0.009271f
C195 VTAIL.n155 B 0.020696f
C196 VTAIL.n156 B 0.044026f
C197 VTAIL.n157 B 0.009271f
C198 VTAIL.n158 B 0.008756f
C199 VTAIL.n159 B 0.039445f
C200 VTAIL.n160 B 0.024608f
C201 VTAIL.n161 B 0.821059f
C202 VTAIL.n162 B 0.022464f
C203 VTAIL.n163 B 0.016295f
C204 VTAIL.n164 B 0.008756f
C205 VTAIL.n165 B 0.020696f
C206 VTAIL.n166 B 0.009271f
C207 VTAIL.n167 B 0.016295f
C208 VTAIL.n168 B 0.009014f
C209 VTAIL.n169 B 0.020696f
C210 VTAIL.n170 B 0.008756f
C211 VTAIL.n171 B 0.009271f
C212 VTAIL.n172 B 0.016295f
C213 VTAIL.n173 B 0.008756f
C214 VTAIL.n174 B 0.020696f
C215 VTAIL.n175 B 0.009271f
C216 VTAIL.n176 B 0.016295f
C217 VTAIL.n177 B 0.008756f
C218 VTAIL.n178 B 0.015522f
C219 VTAIL.n179 B 0.01463f
C220 VTAIL.t7 B 0.034784f
C221 VTAIL.n180 B 0.105223f
C222 VTAIL.n181 B 0.679975f
C223 VTAIL.n182 B 0.008756f
C224 VTAIL.n183 B 0.009271f
C225 VTAIL.n184 B 0.020696f
C226 VTAIL.n185 B 0.020696f
C227 VTAIL.n186 B 0.009271f
C228 VTAIL.n187 B 0.008756f
C229 VTAIL.n188 B 0.016295f
C230 VTAIL.n189 B 0.016295f
C231 VTAIL.n190 B 0.008756f
C232 VTAIL.n191 B 0.009271f
C233 VTAIL.n192 B 0.020696f
C234 VTAIL.n193 B 0.020696f
C235 VTAIL.n194 B 0.009271f
C236 VTAIL.n195 B 0.008756f
C237 VTAIL.n196 B 0.016295f
C238 VTAIL.n197 B 0.016295f
C239 VTAIL.n198 B 0.008756f
C240 VTAIL.n199 B 0.009271f
C241 VTAIL.n200 B 0.020696f
C242 VTAIL.n201 B 0.020696f
C243 VTAIL.n202 B 0.020696f
C244 VTAIL.n203 B 0.009014f
C245 VTAIL.n204 B 0.008756f
C246 VTAIL.n205 B 0.016295f
C247 VTAIL.n206 B 0.016295f
C248 VTAIL.n207 B 0.008756f
C249 VTAIL.n208 B 0.009271f
C250 VTAIL.n209 B 0.020696f
C251 VTAIL.n210 B 0.044026f
C252 VTAIL.n211 B 0.009271f
C253 VTAIL.n212 B 0.008756f
C254 VTAIL.n213 B 0.039445f
C255 VTAIL.n214 B 0.024608f
C256 VTAIL.n215 B 0.821059f
C257 VTAIL.n216 B 0.022464f
C258 VTAIL.n217 B 0.016295f
C259 VTAIL.n218 B 0.008756f
C260 VTAIL.n219 B 0.020696f
C261 VTAIL.n220 B 0.009271f
C262 VTAIL.n221 B 0.016295f
C263 VTAIL.n222 B 0.009014f
C264 VTAIL.n223 B 0.020696f
C265 VTAIL.n224 B 0.008756f
C266 VTAIL.n225 B 0.009271f
C267 VTAIL.n226 B 0.016295f
C268 VTAIL.n227 B 0.008756f
C269 VTAIL.n228 B 0.020696f
C270 VTAIL.n229 B 0.009271f
C271 VTAIL.n230 B 0.016295f
C272 VTAIL.n231 B 0.008756f
C273 VTAIL.n232 B 0.015522f
C274 VTAIL.n233 B 0.01463f
C275 VTAIL.t5 B 0.034784f
C276 VTAIL.n234 B 0.105223f
C277 VTAIL.n235 B 0.679975f
C278 VTAIL.n236 B 0.008756f
C279 VTAIL.n237 B 0.009271f
C280 VTAIL.n238 B 0.020696f
C281 VTAIL.n239 B 0.020696f
C282 VTAIL.n240 B 0.009271f
C283 VTAIL.n241 B 0.008756f
C284 VTAIL.n242 B 0.016295f
C285 VTAIL.n243 B 0.016295f
C286 VTAIL.n244 B 0.008756f
C287 VTAIL.n245 B 0.009271f
C288 VTAIL.n246 B 0.020696f
C289 VTAIL.n247 B 0.020696f
C290 VTAIL.n248 B 0.009271f
C291 VTAIL.n249 B 0.008756f
C292 VTAIL.n250 B 0.016295f
C293 VTAIL.n251 B 0.016295f
C294 VTAIL.n252 B 0.008756f
C295 VTAIL.n253 B 0.009271f
C296 VTAIL.n254 B 0.020696f
C297 VTAIL.n255 B 0.020696f
C298 VTAIL.n256 B 0.020696f
C299 VTAIL.n257 B 0.009014f
C300 VTAIL.n258 B 0.008756f
C301 VTAIL.n259 B 0.016295f
C302 VTAIL.n260 B 0.016295f
C303 VTAIL.n261 B 0.008756f
C304 VTAIL.n262 B 0.009271f
C305 VTAIL.n263 B 0.020696f
C306 VTAIL.n264 B 0.044026f
C307 VTAIL.n265 B 0.009271f
C308 VTAIL.n266 B 0.008756f
C309 VTAIL.n267 B 0.039445f
C310 VTAIL.n268 B 0.024608f
C311 VTAIL.n269 B 0.104769f
C312 VTAIL.n270 B 0.022464f
C313 VTAIL.n271 B 0.016295f
C314 VTAIL.n272 B 0.008756f
C315 VTAIL.n273 B 0.020696f
C316 VTAIL.n274 B 0.009271f
C317 VTAIL.n275 B 0.016295f
C318 VTAIL.n276 B 0.009014f
C319 VTAIL.n277 B 0.020696f
C320 VTAIL.n278 B 0.008756f
C321 VTAIL.n279 B 0.009271f
C322 VTAIL.n280 B 0.016295f
C323 VTAIL.n281 B 0.008756f
C324 VTAIL.n282 B 0.020696f
C325 VTAIL.n283 B 0.009271f
C326 VTAIL.n284 B 0.016295f
C327 VTAIL.n285 B 0.008756f
C328 VTAIL.n286 B 0.015522f
C329 VTAIL.n287 B 0.01463f
C330 VTAIL.t3 B 0.034784f
C331 VTAIL.n288 B 0.105223f
C332 VTAIL.n289 B 0.679975f
C333 VTAIL.n290 B 0.008756f
C334 VTAIL.n291 B 0.009271f
C335 VTAIL.n292 B 0.020696f
C336 VTAIL.n293 B 0.020696f
C337 VTAIL.n294 B 0.009271f
C338 VTAIL.n295 B 0.008756f
C339 VTAIL.n296 B 0.016295f
C340 VTAIL.n297 B 0.016295f
C341 VTAIL.n298 B 0.008756f
C342 VTAIL.n299 B 0.009271f
C343 VTAIL.n300 B 0.020696f
C344 VTAIL.n301 B 0.020696f
C345 VTAIL.n302 B 0.009271f
C346 VTAIL.n303 B 0.008756f
C347 VTAIL.n304 B 0.016295f
C348 VTAIL.n305 B 0.016295f
C349 VTAIL.n306 B 0.008756f
C350 VTAIL.n307 B 0.009271f
C351 VTAIL.n308 B 0.020696f
C352 VTAIL.n309 B 0.020696f
C353 VTAIL.n310 B 0.020696f
C354 VTAIL.n311 B 0.009014f
C355 VTAIL.n312 B 0.008756f
C356 VTAIL.n313 B 0.016295f
C357 VTAIL.n314 B 0.016295f
C358 VTAIL.n315 B 0.008756f
C359 VTAIL.n316 B 0.009271f
C360 VTAIL.n317 B 0.020696f
C361 VTAIL.n318 B 0.044026f
C362 VTAIL.n319 B 0.009271f
C363 VTAIL.n320 B 0.008756f
C364 VTAIL.n321 B 0.039445f
C365 VTAIL.n322 B 0.024608f
C366 VTAIL.n323 B 0.104769f
C367 VTAIL.n324 B 0.022464f
C368 VTAIL.n325 B 0.016295f
C369 VTAIL.n326 B 0.008756f
C370 VTAIL.n327 B 0.020696f
C371 VTAIL.n328 B 0.009271f
C372 VTAIL.n329 B 0.016295f
C373 VTAIL.n330 B 0.009014f
C374 VTAIL.n331 B 0.020696f
C375 VTAIL.n332 B 0.008756f
C376 VTAIL.n333 B 0.009271f
C377 VTAIL.n334 B 0.016295f
C378 VTAIL.n335 B 0.008756f
C379 VTAIL.n336 B 0.020696f
C380 VTAIL.n337 B 0.009271f
C381 VTAIL.n338 B 0.016295f
C382 VTAIL.n339 B 0.008756f
C383 VTAIL.n340 B 0.015522f
C384 VTAIL.n341 B 0.01463f
C385 VTAIL.t1 B 0.034784f
C386 VTAIL.n342 B 0.105223f
C387 VTAIL.n343 B 0.679975f
C388 VTAIL.n344 B 0.008756f
C389 VTAIL.n345 B 0.009271f
C390 VTAIL.n346 B 0.020696f
C391 VTAIL.n347 B 0.020696f
C392 VTAIL.n348 B 0.009271f
C393 VTAIL.n349 B 0.008756f
C394 VTAIL.n350 B 0.016295f
C395 VTAIL.n351 B 0.016295f
C396 VTAIL.n352 B 0.008756f
C397 VTAIL.n353 B 0.009271f
C398 VTAIL.n354 B 0.020696f
C399 VTAIL.n355 B 0.020696f
C400 VTAIL.n356 B 0.009271f
C401 VTAIL.n357 B 0.008756f
C402 VTAIL.n358 B 0.016295f
C403 VTAIL.n359 B 0.016295f
C404 VTAIL.n360 B 0.008756f
C405 VTAIL.n361 B 0.009271f
C406 VTAIL.n362 B 0.020696f
C407 VTAIL.n363 B 0.020696f
C408 VTAIL.n364 B 0.020696f
C409 VTAIL.n365 B 0.009014f
C410 VTAIL.n366 B 0.008756f
C411 VTAIL.n367 B 0.016295f
C412 VTAIL.n368 B 0.016295f
C413 VTAIL.n369 B 0.008756f
C414 VTAIL.n370 B 0.009271f
C415 VTAIL.n371 B 0.020696f
C416 VTAIL.n372 B 0.044026f
C417 VTAIL.n373 B 0.009271f
C418 VTAIL.n374 B 0.008756f
C419 VTAIL.n375 B 0.039445f
C420 VTAIL.n376 B 0.024608f
C421 VTAIL.n377 B 0.821059f
C422 VTAIL.n378 B 0.022464f
C423 VTAIL.n379 B 0.016295f
C424 VTAIL.n380 B 0.008756f
C425 VTAIL.n381 B 0.020696f
C426 VTAIL.n382 B 0.009271f
C427 VTAIL.n383 B 0.016295f
C428 VTAIL.n384 B 0.009014f
C429 VTAIL.n385 B 0.020696f
C430 VTAIL.n386 B 0.009271f
C431 VTAIL.n387 B 0.016295f
C432 VTAIL.n388 B 0.008756f
C433 VTAIL.n389 B 0.020696f
C434 VTAIL.n390 B 0.009271f
C435 VTAIL.n391 B 0.016295f
C436 VTAIL.n392 B 0.008756f
C437 VTAIL.n393 B 0.015522f
C438 VTAIL.n394 B 0.01463f
C439 VTAIL.t6 B 0.034784f
C440 VTAIL.n395 B 0.105223f
C441 VTAIL.n396 B 0.679975f
C442 VTAIL.n397 B 0.008756f
C443 VTAIL.n398 B 0.009271f
C444 VTAIL.n399 B 0.020696f
C445 VTAIL.n400 B 0.020696f
C446 VTAIL.n401 B 0.009271f
C447 VTAIL.n402 B 0.008756f
C448 VTAIL.n403 B 0.016295f
C449 VTAIL.n404 B 0.016295f
C450 VTAIL.n405 B 0.008756f
C451 VTAIL.n406 B 0.009271f
C452 VTAIL.n407 B 0.020696f
C453 VTAIL.n408 B 0.020696f
C454 VTAIL.n409 B 0.009271f
C455 VTAIL.n410 B 0.008756f
C456 VTAIL.n411 B 0.016295f
C457 VTAIL.n412 B 0.016295f
C458 VTAIL.n413 B 0.008756f
C459 VTAIL.n414 B 0.008756f
C460 VTAIL.n415 B 0.009271f
C461 VTAIL.n416 B 0.020696f
C462 VTAIL.n417 B 0.020696f
C463 VTAIL.n418 B 0.020696f
C464 VTAIL.n419 B 0.009014f
C465 VTAIL.n420 B 0.008756f
C466 VTAIL.n421 B 0.016295f
C467 VTAIL.n422 B 0.016295f
C468 VTAIL.n423 B 0.008756f
C469 VTAIL.n424 B 0.009271f
C470 VTAIL.n425 B 0.020696f
C471 VTAIL.n426 B 0.044026f
C472 VTAIL.n427 B 0.009271f
C473 VTAIL.n428 B 0.008756f
C474 VTAIL.n429 B 0.039445f
C475 VTAIL.n430 B 0.024608f
C476 VTAIL.n431 B 0.785414f
C477 VN.t3 B 1.34515f
C478 VN.t0 B 1.34495f
C479 VN.n0 B 0.997992f
C480 VN.t1 B 1.34515f
C481 VN.t2 B 1.34495f
C482 VN.n1 B 1.98332f
.ends

