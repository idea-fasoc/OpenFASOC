* NGSPICE file created from diff_pair_sample_0776.ext - technology: sky130A

.subckt diff_pair_sample_0776 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 w_n2458_n1362# sky130_fd_pr__pfet_01v8 ad=0.7683 pd=4.72 as=0.7683 ps=4.72 w=1.97 l=3.39
X1 VDD1.t1 VP.t0 VTAIL.t0 w_n2458_n1362# sky130_fd_pr__pfet_01v8 ad=0.7683 pd=4.72 as=0.7683 ps=4.72 w=1.97 l=3.39
X2 VDD2.t0 VN.t1 VTAIL.t1 w_n2458_n1362# sky130_fd_pr__pfet_01v8 ad=0.7683 pd=4.72 as=0.7683 ps=4.72 w=1.97 l=3.39
X3 B.t11 B.t9 B.t10 w_n2458_n1362# sky130_fd_pr__pfet_01v8 ad=0.7683 pd=4.72 as=0 ps=0 w=1.97 l=3.39
X4 VDD1.t0 VP.t1 VTAIL.t3 w_n2458_n1362# sky130_fd_pr__pfet_01v8 ad=0.7683 pd=4.72 as=0.7683 ps=4.72 w=1.97 l=3.39
X5 B.t8 B.t6 B.t7 w_n2458_n1362# sky130_fd_pr__pfet_01v8 ad=0.7683 pd=4.72 as=0 ps=0 w=1.97 l=3.39
X6 B.t5 B.t3 B.t4 w_n2458_n1362# sky130_fd_pr__pfet_01v8 ad=0.7683 pd=4.72 as=0 ps=0 w=1.97 l=3.39
X7 B.t2 B.t0 B.t1 w_n2458_n1362# sky130_fd_pr__pfet_01v8 ad=0.7683 pd=4.72 as=0 ps=0 w=1.97 l=3.39
R0 VN VN.t1 91.8532
R1 VN VN.t0 53.3191
R2 VTAIL.n26 VTAIL.n24 756.745
R3 VTAIL.n2 VTAIL.n0 756.745
R4 VTAIL.n18 VTAIL.n16 756.745
R5 VTAIL.n10 VTAIL.n8 756.745
R6 VTAIL.n27 VTAIL.n26 585
R7 VTAIL.n3 VTAIL.n2 585
R8 VTAIL.n19 VTAIL.n18 585
R9 VTAIL.n11 VTAIL.n10 585
R10 VTAIL.t2 VTAIL.n25 417.779
R11 VTAIL.t3 VTAIL.n1 417.779
R12 VTAIL.t0 VTAIL.n17 417.779
R13 VTAIL.t1 VTAIL.n9 417.779
R14 VTAIL.n26 VTAIL.t2 85.8723
R15 VTAIL.n2 VTAIL.t3 85.8723
R16 VTAIL.n18 VTAIL.t0 85.8723
R17 VTAIL.n10 VTAIL.t1 85.8723
R18 VTAIL.n31 VTAIL.n30 30.8278
R19 VTAIL.n7 VTAIL.n6 30.8278
R20 VTAIL.n23 VTAIL.n22 30.8278
R21 VTAIL.n15 VTAIL.n14 30.8278
R22 VTAIL.n15 VTAIL.n7 20.4789
R23 VTAIL.n31 VTAIL.n23 17.2721
R24 VTAIL.n27 VTAIL.n25 9.84608
R25 VTAIL.n3 VTAIL.n1 9.84608
R26 VTAIL.n19 VTAIL.n17 9.84608
R27 VTAIL.n11 VTAIL.n9 9.84608
R28 VTAIL.n30 VTAIL.n29 9.45567
R29 VTAIL.n6 VTAIL.n5 9.45567
R30 VTAIL.n22 VTAIL.n21 9.45567
R31 VTAIL.n14 VTAIL.n13 9.45567
R32 VTAIL.n29 VTAIL.n28 9.3005
R33 VTAIL.n5 VTAIL.n4 9.3005
R34 VTAIL.n21 VTAIL.n20 9.3005
R35 VTAIL.n13 VTAIL.n12 9.3005
R36 VTAIL.n30 VTAIL.n24 8.14595
R37 VTAIL.n6 VTAIL.n0 8.14595
R38 VTAIL.n22 VTAIL.n16 8.14595
R39 VTAIL.n14 VTAIL.n8 8.14595
R40 VTAIL.n28 VTAIL.n27 7.3702
R41 VTAIL.n4 VTAIL.n3 7.3702
R42 VTAIL.n20 VTAIL.n19 7.3702
R43 VTAIL.n12 VTAIL.n11 7.3702
R44 VTAIL.n28 VTAIL.n24 5.81868
R45 VTAIL.n4 VTAIL.n0 5.81868
R46 VTAIL.n20 VTAIL.n16 5.81868
R47 VTAIL.n12 VTAIL.n8 5.81868
R48 VTAIL.n13 VTAIL.n9 3.32369
R49 VTAIL.n29 VTAIL.n25 3.32369
R50 VTAIL.n5 VTAIL.n1 3.32369
R51 VTAIL.n21 VTAIL.n17 3.32369
R52 VTAIL.n23 VTAIL.n15 2.07378
R53 VTAIL VTAIL.n7 1.33024
R54 VTAIL VTAIL.n31 0.744035
R55 VDD2.n9 VDD2.n7 756.745
R56 VDD2.n2 VDD2.n0 756.745
R57 VDD2.n10 VDD2.n9 585
R58 VDD2.n3 VDD2.n2 585
R59 VDD2.t1 VDD2.n1 417.779
R60 VDD2.t0 VDD2.n8 417.779
R61 VDD2.n9 VDD2.t0 85.8723
R62 VDD2.n2 VDD2.t1 85.8723
R63 VDD2.n14 VDD2.n6 79.2781
R64 VDD2.n14 VDD2.n13 47.5066
R65 VDD2.n10 VDD2.n8 9.84608
R66 VDD2.n3 VDD2.n1 9.84608
R67 VDD2.n13 VDD2.n12 9.45567
R68 VDD2.n6 VDD2.n5 9.45567
R69 VDD2.n12 VDD2.n11 9.3005
R70 VDD2.n5 VDD2.n4 9.3005
R71 VDD2.n13 VDD2.n7 8.14595
R72 VDD2.n6 VDD2.n0 8.14595
R73 VDD2.n11 VDD2.n10 7.3702
R74 VDD2.n4 VDD2.n3 7.3702
R75 VDD2.n11 VDD2.n7 5.81868
R76 VDD2.n4 VDD2.n0 5.81868
R77 VDD2.n12 VDD2.n8 3.32369
R78 VDD2.n5 VDD2.n1 3.32369
R79 VDD2 VDD2.n14 0.860414
R80 VP.n0 VP.t0 91.9461
R81 VP.n0 VP.t1 52.7933
R82 VP VP.n0 0.52637
R83 VDD1.n2 VDD1.n0 756.745
R84 VDD1.n9 VDD1.n7 756.745
R85 VDD1.n3 VDD1.n2 585
R86 VDD1.n10 VDD1.n9 585
R87 VDD1.t0 VDD1.n8 417.779
R88 VDD1.t1 VDD1.n1 417.779
R89 VDD1.n2 VDD1.t1 85.8723
R90 VDD1.n9 VDD1.t0 85.8723
R91 VDD1 VDD1.n13 80.6046
R92 VDD1 VDD1.n6 48.3665
R93 VDD1.n3 VDD1.n1 9.84608
R94 VDD1.n10 VDD1.n8 9.84608
R95 VDD1.n6 VDD1.n5 9.45567
R96 VDD1.n13 VDD1.n12 9.45567
R97 VDD1.n5 VDD1.n4 9.3005
R98 VDD1.n12 VDD1.n11 9.3005
R99 VDD1.n6 VDD1.n0 8.14595
R100 VDD1.n13 VDD1.n7 8.14595
R101 VDD1.n4 VDD1.n3 7.3702
R102 VDD1.n11 VDD1.n10 7.3702
R103 VDD1.n4 VDD1.n0 5.81868
R104 VDD1.n11 VDD1.n7 5.81868
R105 VDD1.n5 VDD1.n1 3.32369
R106 VDD1.n12 VDD1.n8 3.32369
R107 B.n293 B.n38 585
R108 B.n295 B.n294 585
R109 B.n296 B.n37 585
R110 B.n298 B.n297 585
R111 B.n299 B.n36 585
R112 B.n301 B.n300 585
R113 B.n302 B.n35 585
R114 B.n304 B.n303 585
R115 B.n305 B.n34 585
R116 B.n307 B.n306 585
R117 B.n308 B.n33 585
R118 B.n310 B.n309 585
R119 B.n312 B.n311 585
R120 B.n313 B.n29 585
R121 B.n315 B.n314 585
R122 B.n316 B.n28 585
R123 B.n318 B.n317 585
R124 B.n319 B.n27 585
R125 B.n321 B.n320 585
R126 B.n322 B.n26 585
R127 B.n324 B.n323 585
R128 B.n325 B.n23 585
R129 B.n328 B.n327 585
R130 B.n329 B.n22 585
R131 B.n331 B.n330 585
R132 B.n332 B.n21 585
R133 B.n334 B.n333 585
R134 B.n335 B.n20 585
R135 B.n337 B.n336 585
R136 B.n338 B.n19 585
R137 B.n340 B.n339 585
R138 B.n341 B.n18 585
R139 B.n343 B.n342 585
R140 B.n344 B.n17 585
R141 B.n292 B.n291 585
R142 B.n290 B.n39 585
R143 B.n289 B.n288 585
R144 B.n287 B.n40 585
R145 B.n286 B.n285 585
R146 B.n284 B.n41 585
R147 B.n283 B.n282 585
R148 B.n281 B.n42 585
R149 B.n280 B.n279 585
R150 B.n278 B.n43 585
R151 B.n277 B.n276 585
R152 B.n275 B.n44 585
R153 B.n274 B.n273 585
R154 B.n272 B.n45 585
R155 B.n271 B.n270 585
R156 B.n269 B.n46 585
R157 B.n268 B.n267 585
R158 B.n266 B.n47 585
R159 B.n265 B.n264 585
R160 B.n263 B.n48 585
R161 B.n262 B.n261 585
R162 B.n260 B.n49 585
R163 B.n259 B.n258 585
R164 B.n257 B.n50 585
R165 B.n256 B.n255 585
R166 B.n254 B.n51 585
R167 B.n253 B.n252 585
R168 B.n251 B.n52 585
R169 B.n250 B.n249 585
R170 B.n248 B.n53 585
R171 B.n247 B.n246 585
R172 B.n245 B.n54 585
R173 B.n244 B.n243 585
R174 B.n242 B.n55 585
R175 B.n241 B.n240 585
R176 B.n239 B.n56 585
R177 B.n238 B.n237 585
R178 B.n236 B.n57 585
R179 B.n235 B.n234 585
R180 B.n233 B.n58 585
R181 B.n232 B.n231 585
R182 B.n230 B.n59 585
R183 B.n229 B.n228 585
R184 B.n227 B.n60 585
R185 B.n226 B.n225 585
R186 B.n224 B.n61 585
R187 B.n223 B.n222 585
R188 B.n221 B.n62 585
R189 B.n220 B.n219 585
R190 B.n218 B.n63 585
R191 B.n217 B.n216 585
R192 B.n215 B.n64 585
R193 B.n214 B.n213 585
R194 B.n212 B.n65 585
R195 B.n211 B.n210 585
R196 B.n209 B.n66 585
R197 B.n208 B.n207 585
R198 B.n206 B.n67 585
R199 B.n205 B.n204 585
R200 B.n203 B.n68 585
R201 B.n202 B.n201 585
R202 B.n149 B.n90 585
R203 B.n151 B.n150 585
R204 B.n152 B.n89 585
R205 B.n154 B.n153 585
R206 B.n155 B.n88 585
R207 B.n157 B.n156 585
R208 B.n158 B.n87 585
R209 B.n160 B.n159 585
R210 B.n161 B.n86 585
R211 B.n163 B.n162 585
R212 B.n164 B.n85 585
R213 B.n166 B.n165 585
R214 B.n168 B.n167 585
R215 B.n169 B.n81 585
R216 B.n171 B.n170 585
R217 B.n172 B.n80 585
R218 B.n174 B.n173 585
R219 B.n175 B.n79 585
R220 B.n177 B.n176 585
R221 B.n178 B.n78 585
R222 B.n180 B.n179 585
R223 B.n181 B.n75 585
R224 B.n184 B.n183 585
R225 B.n185 B.n74 585
R226 B.n187 B.n186 585
R227 B.n188 B.n73 585
R228 B.n190 B.n189 585
R229 B.n191 B.n72 585
R230 B.n193 B.n192 585
R231 B.n194 B.n71 585
R232 B.n196 B.n195 585
R233 B.n197 B.n70 585
R234 B.n199 B.n198 585
R235 B.n200 B.n69 585
R236 B.n148 B.n147 585
R237 B.n146 B.n91 585
R238 B.n145 B.n144 585
R239 B.n143 B.n92 585
R240 B.n142 B.n141 585
R241 B.n140 B.n93 585
R242 B.n139 B.n138 585
R243 B.n137 B.n94 585
R244 B.n136 B.n135 585
R245 B.n134 B.n95 585
R246 B.n133 B.n132 585
R247 B.n131 B.n96 585
R248 B.n130 B.n129 585
R249 B.n128 B.n97 585
R250 B.n127 B.n126 585
R251 B.n125 B.n98 585
R252 B.n124 B.n123 585
R253 B.n122 B.n99 585
R254 B.n121 B.n120 585
R255 B.n119 B.n100 585
R256 B.n118 B.n117 585
R257 B.n116 B.n101 585
R258 B.n115 B.n114 585
R259 B.n113 B.n102 585
R260 B.n112 B.n111 585
R261 B.n110 B.n103 585
R262 B.n109 B.n108 585
R263 B.n107 B.n104 585
R264 B.n106 B.n105 585
R265 B.n2 B.n0 585
R266 B.n389 B.n1 585
R267 B.n388 B.n387 585
R268 B.n386 B.n3 585
R269 B.n385 B.n384 585
R270 B.n383 B.n4 585
R271 B.n382 B.n381 585
R272 B.n380 B.n5 585
R273 B.n379 B.n378 585
R274 B.n377 B.n6 585
R275 B.n376 B.n375 585
R276 B.n374 B.n7 585
R277 B.n373 B.n372 585
R278 B.n371 B.n8 585
R279 B.n370 B.n369 585
R280 B.n368 B.n9 585
R281 B.n367 B.n366 585
R282 B.n365 B.n10 585
R283 B.n364 B.n363 585
R284 B.n362 B.n11 585
R285 B.n361 B.n360 585
R286 B.n359 B.n12 585
R287 B.n358 B.n357 585
R288 B.n356 B.n13 585
R289 B.n355 B.n354 585
R290 B.n353 B.n14 585
R291 B.n352 B.n351 585
R292 B.n350 B.n15 585
R293 B.n349 B.n348 585
R294 B.n347 B.n16 585
R295 B.n346 B.n345 585
R296 B.n391 B.n390 585
R297 B.n149 B.n148 482.89
R298 B.n346 B.n17 482.89
R299 B.n202 B.n69 482.89
R300 B.n293 B.n292 482.89
R301 B.n76 B.t2 319.901
R302 B.n30 B.t7 319.901
R303 B.n82 B.t5 319.901
R304 B.n24 B.t10 319.901
R305 B.n77 B.t1 247.756
R306 B.n31 B.t8 247.756
R307 B.n83 B.t4 247.756
R308 B.n25 B.t11 247.756
R309 B.n76 B.t0 222.998
R310 B.n82 B.t3 222.998
R311 B.n24 B.t9 222.998
R312 B.n30 B.t6 222.998
R313 B.n148 B.n91 163.367
R314 B.n144 B.n91 163.367
R315 B.n144 B.n143 163.367
R316 B.n143 B.n142 163.367
R317 B.n142 B.n93 163.367
R318 B.n138 B.n93 163.367
R319 B.n138 B.n137 163.367
R320 B.n137 B.n136 163.367
R321 B.n136 B.n95 163.367
R322 B.n132 B.n95 163.367
R323 B.n132 B.n131 163.367
R324 B.n131 B.n130 163.367
R325 B.n130 B.n97 163.367
R326 B.n126 B.n97 163.367
R327 B.n126 B.n125 163.367
R328 B.n125 B.n124 163.367
R329 B.n124 B.n99 163.367
R330 B.n120 B.n99 163.367
R331 B.n120 B.n119 163.367
R332 B.n119 B.n118 163.367
R333 B.n118 B.n101 163.367
R334 B.n114 B.n101 163.367
R335 B.n114 B.n113 163.367
R336 B.n113 B.n112 163.367
R337 B.n112 B.n103 163.367
R338 B.n108 B.n103 163.367
R339 B.n108 B.n107 163.367
R340 B.n107 B.n106 163.367
R341 B.n106 B.n2 163.367
R342 B.n390 B.n2 163.367
R343 B.n390 B.n389 163.367
R344 B.n389 B.n388 163.367
R345 B.n388 B.n3 163.367
R346 B.n384 B.n3 163.367
R347 B.n384 B.n383 163.367
R348 B.n383 B.n382 163.367
R349 B.n382 B.n5 163.367
R350 B.n378 B.n5 163.367
R351 B.n378 B.n377 163.367
R352 B.n377 B.n376 163.367
R353 B.n376 B.n7 163.367
R354 B.n372 B.n7 163.367
R355 B.n372 B.n371 163.367
R356 B.n371 B.n370 163.367
R357 B.n370 B.n9 163.367
R358 B.n366 B.n9 163.367
R359 B.n366 B.n365 163.367
R360 B.n365 B.n364 163.367
R361 B.n364 B.n11 163.367
R362 B.n360 B.n11 163.367
R363 B.n360 B.n359 163.367
R364 B.n359 B.n358 163.367
R365 B.n358 B.n13 163.367
R366 B.n354 B.n13 163.367
R367 B.n354 B.n353 163.367
R368 B.n353 B.n352 163.367
R369 B.n352 B.n15 163.367
R370 B.n348 B.n15 163.367
R371 B.n348 B.n347 163.367
R372 B.n347 B.n346 163.367
R373 B.n150 B.n149 163.367
R374 B.n150 B.n89 163.367
R375 B.n154 B.n89 163.367
R376 B.n155 B.n154 163.367
R377 B.n156 B.n155 163.367
R378 B.n156 B.n87 163.367
R379 B.n160 B.n87 163.367
R380 B.n161 B.n160 163.367
R381 B.n162 B.n161 163.367
R382 B.n162 B.n85 163.367
R383 B.n166 B.n85 163.367
R384 B.n167 B.n166 163.367
R385 B.n167 B.n81 163.367
R386 B.n171 B.n81 163.367
R387 B.n172 B.n171 163.367
R388 B.n173 B.n172 163.367
R389 B.n173 B.n79 163.367
R390 B.n177 B.n79 163.367
R391 B.n178 B.n177 163.367
R392 B.n179 B.n178 163.367
R393 B.n179 B.n75 163.367
R394 B.n184 B.n75 163.367
R395 B.n185 B.n184 163.367
R396 B.n186 B.n185 163.367
R397 B.n186 B.n73 163.367
R398 B.n190 B.n73 163.367
R399 B.n191 B.n190 163.367
R400 B.n192 B.n191 163.367
R401 B.n192 B.n71 163.367
R402 B.n196 B.n71 163.367
R403 B.n197 B.n196 163.367
R404 B.n198 B.n197 163.367
R405 B.n198 B.n69 163.367
R406 B.n203 B.n202 163.367
R407 B.n204 B.n203 163.367
R408 B.n204 B.n67 163.367
R409 B.n208 B.n67 163.367
R410 B.n209 B.n208 163.367
R411 B.n210 B.n209 163.367
R412 B.n210 B.n65 163.367
R413 B.n214 B.n65 163.367
R414 B.n215 B.n214 163.367
R415 B.n216 B.n215 163.367
R416 B.n216 B.n63 163.367
R417 B.n220 B.n63 163.367
R418 B.n221 B.n220 163.367
R419 B.n222 B.n221 163.367
R420 B.n222 B.n61 163.367
R421 B.n226 B.n61 163.367
R422 B.n227 B.n226 163.367
R423 B.n228 B.n227 163.367
R424 B.n228 B.n59 163.367
R425 B.n232 B.n59 163.367
R426 B.n233 B.n232 163.367
R427 B.n234 B.n233 163.367
R428 B.n234 B.n57 163.367
R429 B.n238 B.n57 163.367
R430 B.n239 B.n238 163.367
R431 B.n240 B.n239 163.367
R432 B.n240 B.n55 163.367
R433 B.n244 B.n55 163.367
R434 B.n245 B.n244 163.367
R435 B.n246 B.n245 163.367
R436 B.n246 B.n53 163.367
R437 B.n250 B.n53 163.367
R438 B.n251 B.n250 163.367
R439 B.n252 B.n251 163.367
R440 B.n252 B.n51 163.367
R441 B.n256 B.n51 163.367
R442 B.n257 B.n256 163.367
R443 B.n258 B.n257 163.367
R444 B.n258 B.n49 163.367
R445 B.n262 B.n49 163.367
R446 B.n263 B.n262 163.367
R447 B.n264 B.n263 163.367
R448 B.n264 B.n47 163.367
R449 B.n268 B.n47 163.367
R450 B.n269 B.n268 163.367
R451 B.n270 B.n269 163.367
R452 B.n270 B.n45 163.367
R453 B.n274 B.n45 163.367
R454 B.n275 B.n274 163.367
R455 B.n276 B.n275 163.367
R456 B.n276 B.n43 163.367
R457 B.n280 B.n43 163.367
R458 B.n281 B.n280 163.367
R459 B.n282 B.n281 163.367
R460 B.n282 B.n41 163.367
R461 B.n286 B.n41 163.367
R462 B.n287 B.n286 163.367
R463 B.n288 B.n287 163.367
R464 B.n288 B.n39 163.367
R465 B.n292 B.n39 163.367
R466 B.n342 B.n17 163.367
R467 B.n342 B.n341 163.367
R468 B.n341 B.n340 163.367
R469 B.n340 B.n19 163.367
R470 B.n336 B.n19 163.367
R471 B.n336 B.n335 163.367
R472 B.n335 B.n334 163.367
R473 B.n334 B.n21 163.367
R474 B.n330 B.n21 163.367
R475 B.n330 B.n329 163.367
R476 B.n329 B.n328 163.367
R477 B.n328 B.n23 163.367
R478 B.n323 B.n23 163.367
R479 B.n323 B.n322 163.367
R480 B.n322 B.n321 163.367
R481 B.n321 B.n27 163.367
R482 B.n317 B.n27 163.367
R483 B.n317 B.n316 163.367
R484 B.n316 B.n315 163.367
R485 B.n315 B.n29 163.367
R486 B.n311 B.n29 163.367
R487 B.n311 B.n310 163.367
R488 B.n310 B.n33 163.367
R489 B.n306 B.n33 163.367
R490 B.n306 B.n305 163.367
R491 B.n305 B.n304 163.367
R492 B.n304 B.n35 163.367
R493 B.n300 B.n35 163.367
R494 B.n300 B.n299 163.367
R495 B.n299 B.n298 163.367
R496 B.n298 B.n37 163.367
R497 B.n294 B.n37 163.367
R498 B.n294 B.n293 163.367
R499 B.n77 B.n76 72.146
R500 B.n83 B.n82 72.146
R501 B.n25 B.n24 72.146
R502 B.n31 B.n30 72.146
R503 B.n182 B.n77 59.5399
R504 B.n84 B.n83 59.5399
R505 B.n326 B.n25 59.5399
R506 B.n32 B.n31 59.5399
R507 B.n345 B.n344 31.3761
R508 B.n291 B.n38 31.3761
R509 B.n201 B.n200 31.3761
R510 B.n147 B.n90 31.3761
R511 B B.n391 18.0485
R512 B.n344 B.n343 10.6151
R513 B.n343 B.n18 10.6151
R514 B.n339 B.n18 10.6151
R515 B.n339 B.n338 10.6151
R516 B.n338 B.n337 10.6151
R517 B.n337 B.n20 10.6151
R518 B.n333 B.n20 10.6151
R519 B.n333 B.n332 10.6151
R520 B.n332 B.n331 10.6151
R521 B.n331 B.n22 10.6151
R522 B.n327 B.n22 10.6151
R523 B.n325 B.n324 10.6151
R524 B.n324 B.n26 10.6151
R525 B.n320 B.n26 10.6151
R526 B.n320 B.n319 10.6151
R527 B.n319 B.n318 10.6151
R528 B.n318 B.n28 10.6151
R529 B.n314 B.n28 10.6151
R530 B.n314 B.n313 10.6151
R531 B.n313 B.n312 10.6151
R532 B.n309 B.n308 10.6151
R533 B.n308 B.n307 10.6151
R534 B.n307 B.n34 10.6151
R535 B.n303 B.n34 10.6151
R536 B.n303 B.n302 10.6151
R537 B.n302 B.n301 10.6151
R538 B.n301 B.n36 10.6151
R539 B.n297 B.n36 10.6151
R540 B.n297 B.n296 10.6151
R541 B.n296 B.n295 10.6151
R542 B.n295 B.n38 10.6151
R543 B.n201 B.n68 10.6151
R544 B.n205 B.n68 10.6151
R545 B.n206 B.n205 10.6151
R546 B.n207 B.n206 10.6151
R547 B.n207 B.n66 10.6151
R548 B.n211 B.n66 10.6151
R549 B.n212 B.n211 10.6151
R550 B.n213 B.n212 10.6151
R551 B.n213 B.n64 10.6151
R552 B.n217 B.n64 10.6151
R553 B.n218 B.n217 10.6151
R554 B.n219 B.n218 10.6151
R555 B.n219 B.n62 10.6151
R556 B.n223 B.n62 10.6151
R557 B.n224 B.n223 10.6151
R558 B.n225 B.n224 10.6151
R559 B.n225 B.n60 10.6151
R560 B.n229 B.n60 10.6151
R561 B.n230 B.n229 10.6151
R562 B.n231 B.n230 10.6151
R563 B.n231 B.n58 10.6151
R564 B.n235 B.n58 10.6151
R565 B.n236 B.n235 10.6151
R566 B.n237 B.n236 10.6151
R567 B.n237 B.n56 10.6151
R568 B.n241 B.n56 10.6151
R569 B.n242 B.n241 10.6151
R570 B.n243 B.n242 10.6151
R571 B.n243 B.n54 10.6151
R572 B.n247 B.n54 10.6151
R573 B.n248 B.n247 10.6151
R574 B.n249 B.n248 10.6151
R575 B.n249 B.n52 10.6151
R576 B.n253 B.n52 10.6151
R577 B.n254 B.n253 10.6151
R578 B.n255 B.n254 10.6151
R579 B.n255 B.n50 10.6151
R580 B.n259 B.n50 10.6151
R581 B.n260 B.n259 10.6151
R582 B.n261 B.n260 10.6151
R583 B.n261 B.n48 10.6151
R584 B.n265 B.n48 10.6151
R585 B.n266 B.n265 10.6151
R586 B.n267 B.n266 10.6151
R587 B.n267 B.n46 10.6151
R588 B.n271 B.n46 10.6151
R589 B.n272 B.n271 10.6151
R590 B.n273 B.n272 10.6151
R591 B.n273 B.n44 10.6151
R592 B.n277 B.n44 10.6151
R593 B.n278 B.n277 10.6151
R594 B.n279 B.n278 10.6151
R595 B.n279 B.n42 10.6151
R596 B.n283 B.n42 10.6151
R597 B.n284 B.n283 10.6151
R598 B.n285 B.n284 10.6151
R599 B.n285 B.n40 10.6151
R600 B.n289 B.n40 10.6151
R601 B.n290 B.n289 10.6151
R602 B.n291 B.n290 10.6151
R603 B.n151 B.n90 10.6151
R604 B.n152 B.n151 10.6151
R605 B.n153 B.n152 10.6151
R606 B.n153 B.n88 10.6151
R607 B.n157 B.n88 10.6151
R608 B.n158 B.n157 10.6151
R609 B.n159 B.n158 10.6151
R610 B.n159 B.n86 10.6151
R611 B.n163 B.n86 10.6151
R612 B.n164 B.n163 10.6151
R613 B.n165 B.n164 10.6151
R614 B.n169 B.n168 10.6151
R615 B.n170 B.n169 10.6151
R616 B.n170 B.n80 10.6151
R617 B.n174 B.n80 10.6151
R618 B.n175 B.n174 10.6151
R619 B.n176 B.n175 10.6151
R620 B.n176 B.n78 10.6151
R621 B.n180 B.n78 10.6151
R622 B.n181 B.n180 10.6151
R623 B.n183 B.n74 10.6151
R624 B.n187 B.n74 10.6151
R625 B.n188 B.n187 10.6151
R626 B.n189 B.n188 10.6151
R627 B.n189 B.n72 10.6151
R628 B.n193 B.n72 10.6151
R629 B.n194 B.n193 10.6151
R630 B.n195 B.n194 10.6151
R631 B.n195 B.n70 10.6151
R632 B.n199 B.n70 10.6151
R633 B.n200 B.n199 10.6151
R634 B.n147 B.n146 10.6151
R635 B.n146 B.n145 10.6151
R636 B.n145 B.n92 10.6151
R637 B.n141 B.n92 10.6151
R638 B.n141 B.n140 10.6151
R639 B.n140 B.n139 10.6151
R640 B.n139 B.n94 10.6151
R641 B.n135 B.n94 10.6151
R642 B.n135 B.n134 10.6151
R643 B.n134 B.n133 10.6151
R644 B.n133 B.n96 10.6151
R645 B.n129 B.n96 10.6151
R646 B.n129 B.n128 10.6151
R647 B.n128 B.n127 10.6151
R648 B.n127 B.n98 10.6151
R649 B.n123 B.n98 10.6151
R650 B.n123 B.n122 10.6151
R651 B.n122 B.n121 10.6151
R652 B.n121 B.n100 10.6151
R653 B.n117 B.n100 10.6151
R654 B.n117 B.n116 10.6151
R655 B.n116 B.n115 10.6151
R656 B.n115 B.n102 10.6151
R657 B.n111 B.n102 10.6151
R658 B.n111 B.n110 10.6151
R659 B.n110 B.n109 10.6151
R660 B.n109 B.n104 10.6151
R661 B.n105 B.n104 10.6151
R662 B.n105 B.n0 10.6151
R663 B.n387 B.n1 10.6151
R664 B.n387 B.n386 10.6151
R665 B.n386 B.n385 10.6151
R666 B.n385 B.n4 10.6151
R667 B.n381 B.n4 10.6151
R668 B.n381 B.n380 10.6151
R669 B.n380 B.n379 10.6151
R670 B.n379 B.n6 10.6151
R671 B.n375 B.n6 10.6151
R672 B.n375 B.n374 10.6151
R673 B.n374 B.n373 10.6151
R674 B.n373 B.n8 10.6151
R675 B.n369 B.n8 10.6151
R676 B.n369 B.n368 10.6151
R677 B.n368 B.n367 10.6151
R678 B.n367 B.n10 10.6151
R679 B.n363 B.n10 10.6151
R680 B.n363 B.n362 10.6151
R681 B.n362 B.n361 10.6151
R682 B.n361 B.n12 10.6151
R683 B.n357 B.n12 10.6151
R684 B.n357 B.n356 10.6151
R685 B.n356 B.n355 10.6151
R686 B.n355 B.n14 10.6151
R687 B.n351 B.n14 10.6151
R688 B.n351 B.n350 10.6151
R689 B.n350 B.n349 10.6151
R690 B.n349 B.n16 10.6151
R691 B.n345 B.n16 10.6151
R692 B.n327 B.n326 9.36635
R693 B.n309 B.n32 9.36635
R694 B.n165 B.n84 9.36635
R695 B.n183 B.n182 9.36635
R696 B.n391 B.n0 2.81026
R697 B.n391 B.n1 2.81026
R698 B.n326 B.n325 1.24928
R699 B.n312 B.n32 1.24928
R700 B.n168 B.n84 1.24928
R701 B.n182 B.n181 1.24928
C0 B VP 1.53972f
C1 w_n2458_n1362# VTAIL 1.3491f
C2 w_n2458_n1362# B 6.89573f
C3 VDD1 VN 0.154825f
C4 VTAIL B 1.47572f
C5 VDD2 VDD1 0.770134f
C6 VDD1 VP 0.907396f
C7 w_n2458_n1362# VDD1 1.17631f
C8 VDD2 VN 0.691176f
C9 VDD1 VTAIL 2.67512f
C10 VDD1 B 1.0042f
C11 VN VP 3.97692f
C12 w_n2458_n1362# VN 3.26056f
C13 VDD2 VP 0.372759f
C14 w_n2458_n1362# VDD2 1.21127f
C15 VTAIL VN 1.08521f
C16 VN B 1.01975f
C17 w_n2458_n1362# VP 3.57068f
C18 VDD2 VTAIL 2.7335f
C19 VDD2 B 1.04175f
C20 VTAIL VP 1.09934f
C21 VDD2 VSUBS 0.617466f
C22 VDD1 VSUBS 2.442585f
C23 VTAIL VSUBS 0.394519f
C24 VN VSUBS 6.00233f
C25 VP VSUBS 1.443155f
C26 B VSUBS 3.443938f
C27 w_n2458_n1362# VSUBS 42.7397f
C28 B.n0 VSUBS 0.005941f
C29 B.n1 VSUBS 0.005941f
C30 B.n2 VSUBS 0.009394f
C31 B.n3 VSUBS 0.009394f
C32 B.n4 VSUBS 0.009394f
C33 B.n5 VSUBS 0.009394f
C34 B.n6 VSUBS 0.009394f
C35 B.n7 VSUBS 0.009394f
C36 B.n8 VSUBS 0.009394f
C37 B.n9 VSUBS 0.009394f
C38 B.n10 VSUBS 0.009394f
C39 B.n11 VSUBS 0.009394f
C40 B.n12 VSUBS 0.009394f
C41 B.n13 VSUBS 0.009394f
C42 B.n14 VSUBS 0.009394f
C43 B.n15 VSUBS 0.009394f
C44 B.n16 VSUBS 0.009394f
C45 B.n17 VSUBS 0.022048f
C46 B.n18 VSUBS 0.009394f
C47 B.n19 VSUBS 0.009394f
C48 B.n20 VSUBS 0.009394f
C49 B.n21 VSUBS 0.009394f
C50 B.n22 VSUBS 0.009394f
C51 B.n23 VSUBS 0.009394f
C52 B.t11 VSUBS 0.04501f
C53 B.t10 VSUBS 0.063163f
C54 B.t9 VSUBS 0.443378f
C55 B.n24 VSUBS 0.117728f
C56 B.n25 VSUBS 0.09389f
C57 B.n26 VSUBS 0.009394f
C58 B.n27 VSUBS 0.009394f
C59 B.n28 VSUBS 0.009394f
C60 B.n29 VSUBS 0.009394f
C61 B.t8 VSUBS 0.04501f
C62 B.t7 VSUBS 0.063163f
C63 B.t6 VSUBS 0.443378f
C64 B.n30 VSUBS 0.117728f
C65 B.n31 VSUBS 0.09389f
C66 B.n32 VSUBS 0.021766f
C67 B.n33 VSUBS 0.009394f
C68 B.n34 VSUBS 0.009394f
C69 B.n35 VSUBS 0.009394f
C70 B.n36 VSUBS 0.009394f
C71 B.n37 VSUBS 0.009394f
C72 B.n38 VSUBS 0.020892f
C73 B.n39 VSUBS 0.009394f
C74 B.n40 VSUBS 0.009394f
C75 B.n41 VSUBS 0.009394f
C76 B.n42 VSUBS 0.009394f
C77 B.n43 VSUBS 0.009394f
C78 B.n44 VSUBS 0.009394f
C79 B.n45 VSUBS 0.009394f
C80 B.n46 VSUBS 0.009394f
C81 B.n47 VSUBS 0.009394f
C82 B.n48 VSUBS 0.009394f
C83 B.n49 VSUBS 0.009394f
C84 B.n50 VSUBS 0.009394f
C85 B.n51 VSUBS 0.009394f
C86 B.n52 VSUBS 0.009394f
C87 B.n53 VSUBS 0.009394f
C88 B.n54 VSUBS 0.009394f
C89 B.n55 VSUBS 0.009394f
C90 B.n56 VSUBS 0.009394f
C91 B.n57 VSUBS 0.009394f
C92 B.n58 VSUBS 0.009394f
C93 B.n59 VSUBS 0.009394f
C94 B.n60 VSUBS 0.009394f
C95 B.n61 VSUBS 0.009394f
C96 B.n62 VSUBS 0.009394f
C97 B.n63 VSUBS 0.009394f
C98 B.n64 VSUBS 0.009394f
C99 B.n65 VSUBS 0.009394f
C100 B.n66 VSUBS 0.009394f
C101 B.n67 VSUBS 0.009394f
C102 B.n68 VSUBS 0.009394f
C103 B.n69 VSUBS 0.022048f
C104 B.n70 VSUBS 0.009394f
C105 B.n71 VSUBS 0.009394f
C106 B.n72 VSUBS 0.009394f
C107 B.n73 VSUBS 0.009394f
C108 B.n74 VSUBS 0.009394f
C109 B.n75 VSUBS 0.009394f
C110 B.t1 VSUBS 0.04501f
C111 B.t2 VSUBS 0.063163f
C112 B.t0 VSUBS 0.443378f
C113 B.n76 VSUBS 0.117728f
C114 B.n77 VSUBS 0.09389f
C115 B.n78 VSUBS 0.009394f
C116 B.n79 VSUBS 0.009394f
C117 B.n80 VSUBS 0.009394f
C118 B.n81 VSUBS 0.009394f
C119 B.t4 VSUBS 0.04501f
C120 B.t5 VSUBS 0.063163f
C121 B.t3 VSUBS 0.443378f
C122 B.n82 VSUBS 0.117728f
C123 B.n83 VSUBS 0.09389f
C124 B.n84 VSUBS 0.021766f
C125 B.n85 VSUBS 0.009394f
C126 B.n86 VSUBS 0.009394f
C127 B.n87 VSUBS 0.009394f
C128 B.n88 VSUBS 0.009394f
C129 B.n89 VSUBS 0.009394f
C130 B.n90 VSUBS 0.022048f
C131 B.n91 VSUBS 0.009394f
C132 B.n92 VSUBS 0.009394f
C133 B.n93 VSUBS 0.009394f
C134 B.n94 VSUBS 0.009394f
C135 B.n95 VSUBS 0.009394f
C136 B.n96 VSUBS 0.009394f
C137 B.n97 VSUBS 0.009394f
C138 B.n98 VSUBS 0.009394f
C139 B.n99 VSUBS 0.009394f
C140 B.n100 VSUBS 0.009394f
C141 B.n101 VSUBS 0.009394f
C142 B.n102 VSUBS 0.009394f
C143 B.n103 VSUBS 0.009394f
C144 B.n104 VSUBS 0.009394f
C145 B.n105 VSUBS 0.009394f
C146 B.n106 VSUBS 0.009394f
C147 B.n107 VSUBS 0.009394f
C148 B.n108 VSUBS 0.009394f
C149 B.n109 VSUBS 0.009394f
C150 B.n110 VSUBS 0.009394f
C151 B.n111 VSUBS 0.009394f
C152 B.n112 VSUBS 0.009394f
C153 B.n113 VSUBS 0.009394f
C154 B.n114 VSUBS 0.009394f
C155 B.n115 VSUBS 0.009394f
C156 B.n116 VSUBS 0.009394f
C157 B.n117 VSUBS 0.009394f
C158 B.n118 VSUBS 0.009394f
C159 B.n119 VSUBS 0.009394f
C160 B.n120 VSUBS 0.009394f
C161 B.n121 VSUBS 0.009394f
C162 B.n122 VSUBS 0.009394f
C163 B.n123 VSUBS 0.009394f
C164 B.n124 VSUBS 0.009394f
C165 B.n125 VSUBS 0.009394f
C166 B.n126 VSUBS 0.009394f
C167 B.n127 VSUBS 0.009394f
C168 B.n128 VSUBS 0.009394f
C169 B.n129 VSUBS 0.009394f
C170 B.n130 VSUBS 0.009394f
C171 B.n131 VSUBS 0.009394f
C172 B.n132 VSUBS 0.009394f
C173 B.n133 VSUBS 0.009394f
C174 B.n134 VSUBS 0.009394f
C175 B.n135 VSUBS 0.009394f
C176 B.n136 VSUBS 0.009394f
C177 B.n137 VSUBS 0.009394f
C178 B.n138 VSUBS 0.009394f
C179 B.n139 VSUBS 0.009394f
C180 B.n140 VSUBS 0.009394f
C181 B.n141 VSUBS 0.009394f
C182 B.n142 VSUBS 0.009394f
C183 B.n143 VSUBS 0.009394f
C184 B.n144 VSUBS 0.009394f
C185 B.n145 VSUBS 0.009394f
C186 B.n146 VSUBS 0.009394f
C187 B.n147 VSUBS 0.02078f
C188 B.n148 VSUBS 0.02078f
C189 B.n149 VSUBS 0.022048f
C190 B.n150 VSUBS 0.009394f
C191 B.n151 VSUBS 0.009394f
C192 B.n152 VSUBS 0.009394f
C193 B.n153 VSUBS 0.009394f
C194 B.n154 VSUBS 0.009394f
C195 B.n155 VSUBS 0.009394f
C196 B.n156 VSUBS 0.009394f
C197 B.n157 VSUBS 0.009394f
C198 B.n158 VSUBS 0.009394f
C199 B.n159 VSUBS 0.009394f
C200 B.n160 VSUBS 0.009394f
C201 B.n161 VSUBS 0.009394f
C202 B.n162 VSUBS 0.009394f
C203 B.n163 VSUBS 0.009394f
C204 B.n164 VSUBS 0.009394f
C205 B.n165 VSUBS 0.008842f
C206 B.n166 VSUBS 0.009394f
C207 B.n167 VSUBS 0.009394f
C208 B.n168 VSUBS 0.00525f
C209 B.n169 VSUBS 0.009394f
C210 B.n170 VSUBS 0.009394f
C211 B.n171 VSUBS 0.009394f
C212 B.n172 VSUBS 0.009394f
C213 B.n173 VSUBS 0.009394f
C214 B.n174 VSUBS 0.009394f
C215 B.n175 VSUBS 0.009394f
C216 B.n176 VSUBS 0.009394f
C217 B.n177 VSUBS 0.009394f
C218 B.n178 VSUBS 0.009394f
C219 B.n179 VSUBS 0.009394f
C220 B.n180 VSUBS 0.009394f
C221 B.n181 VSUBS 0.00525f
C222 B.n182 VSUBS 0.021766f
C223 B.n183 VSUBS 0.008842f
C224 B.n184 VSUBS 0.009394f
C225 B.n185 VSUBS 0.009394f
C226 B.n186 VSUBS 0.009394f
C227 B.n187 VSUBS 0.009394f
C228 B.n188 VSUBS 0.009394f
C229 B.n189 VSUBS 0.009394f
C230 B.n190 VSUBS 0.009394f
C231 B.n191 VSUBS 0.009394f
C232 B.n192 VSUBS 0.009394f
C233 B.n193 VSUBS 0.009394f
C234 B.n194 VSUBS 0.009394f
C235 B.n195 VSUBS 0.009394f
C236 B.n196 VSUBS 0.009394f
C237 B.n197 VSUBS 0.009394f
C238 B.n198 VSUBS 0.009394f
C239 B.n199 VSUBS 0.009394f
C240 B.n200 VSUBS 0.022048f
C241 B.n201 VSUBS 0.02078f
C242 B.n202 VSUBS 0.02078f
C243 B.n203 VSUBS 0.009394f
C244 B.n204 VSUBS 0.009394f
C245 B.n205 VSUBS 0.009394f
C246 B.n206 VSUBS 0.009394f
C247 B.n207 VSUBS 0.009394f
C248 B.n208 VSUBS 0.009394f
C249 B.n209 VSUBS 0.009394f
C250 B.n210 VSUBS 0.009394f
C251 B.n211 VSUBS 0.009394f
C252 B.n212 VSUBS 0.009394f
C253 B.n213 VSUBS 0.009394f
C254 B.n214 VSUBS 0.009394f
C255 B.n215 VSUBS 0.009394f
C256 B.n216 VSUBS 0.009394f
C257 B.n217 VSUBS 0.009394f
C258 B.n218 VSUBS 0.009394f
C259 B.n219 VSUBS 0.009394f
C260 B.n220 VSUBS 0.009394f
C261 B.n221 VSUBS 0.009394f
C262 B.n222 VSUBS 0.009394f
C263 B.n223 VSUBS 0.009394f
C264 B.n224 VSUBS 0.009394f
C265 B.n225 VSUBS 0.009394f
C266 B.n226 VSUBS 0.009394f
C267 B.n227 VSUBS 0.009394f
C268 B.n228 VSUBS 0.009394f
C269 B.n229 VSUBS 0.009394f
C270 B.n230 VSUBS 0.009394f
C271 B.n231 VSUBS 0.009394f
C272 B.n232 VSUBS 0.009394f
C273 B.n233 VSUBS 0.009394f
C274 B.n234 VSUBS 0.009394f
C275 B.n235 VSUBS 0.009394f
C276 B.n236 VSUBS 0.009394f
C277 B.n237 VSUBS 0.009394f
C278 B.n238 VSUBS 0.009394f
C279 B.n239 VSUBS 0.009394f
C280 B.n240 VSUBS 0.009394f
C281 B.n241 VSUBS 0.009394f
C282 B.n242 VSUBS 0.009394f
C283 B.n243 VSUBS 0.009394f
C284 B.n244 VSUBS 0.009394f
C285 B.n245 VSUBS 0.009394f
C286 B.n246 VSUBS 0.009394f
C287 B.n247 VSUBS 0.009394f
C288 B.n248 VSUBS 0.009394f
C289 B.n249 VSUBS 0.009394f
C290 B.n250 VSUBS 0.009394f
C291 B.n251 VSUBS 0.009394f
C292 B.n252 VSUBS 0.009394f
C293 B.n253 VSUBS 0.009394f
C294 B.n254 VSUBS 0.009394f
C295 B.n255 VSUBS 0.009394f
C296 B.n256 VSUBS 0.009394f
C297 B.n257 VSUBS 0.009394f
C298 B.n258 VSUBS 0.009394f
C299 B.n259 VSUBS 0.009394f
C300 B.n260 VSUBS 0.009394f
C301 B.n261 VSUBS 0.009394f
C302 B.n262 VSUBS 0.009394f
C303 B.n263 VSUBS 0.009394f
C304 B.n264 VSUBS 0.009394f
C305 B.n265 VSUBS 0.009394f
C306 B.n266 VSUBS 0.009394f
C307 B.n267 VSUBS 0.009394f
C308 B.n268 VSUBS 0.009394f
C309 B.n269 VSUBS 0.009394f
C310 B.n270 VSUBS 0.009394f
C311 B.n271 VSUBS 0.009394f
C312 B.n272 VSUBS 0.009394f
C313 B.n273 VSUBS 0.009394f
C314 B.n274 VSUBS 0.009394f
C315 B.n275 VSUBS 0.009394f
C316 B.n276 VSUBS 0.009394f
C317 B.n277 VSUBS 0.009394f
C318 B.n278 VSUBS 0.009394f
C319 B.n279 VSUBS 0.009394f
C320 B.n280 VSUBS 0.009394f
C321 B.n281 VSUBS 0.009394f
C322 B.n282 VSUBS 0.009394f
C323 B.n283 VSUBS 0.009394f
C324 B.n284 VSUBS 0.009394f
C325 B.n285 VSUBS 0.009394f
C326 B.n286 VSUBS 0.009394f
C327 B.n287 VSUBS 0.009394f
C328 B.n288 VSUBS 0.009394f
C329 B.n289 VSUBS 0.009394f
C330 B.n290 VSUBS 0.009394f
C331 B.n291 VSUBS 0.021935f
C332 B.n292 VSUBS 0.02078f
C333 B.n293 VSUBS 0.022048f
C334 B.n294 VSUBS 0.009394f
C335 B.n295 VSUBS 0.009394f
C336 B.n296 VSUBS 0.009394f
C337 B.n297 VSUBS 0.009394f
C338 B.n298 VSUBS 0.009394f
C339 B.n299 VSUBS 0.009394f
C340 B.n300 VSUBS 0.009394f
C341 B.n301 VSUBS 0.009394f
C342 B.n302 VSUBS 0.009394f
C343 B.n303 VSUBS 0.009394f
C344 B.n304 VSUBS 0.009394f
C345 B.n305 VSUBS 0.009394f
C346 B.n306 VSUBS 0.009394f
C347 B.n307 VSUBS 0.009394f
C348 B.n308 VSUBS 0.009394f
C349 B.n309 VSUBS 0.008842f
C350 B.n310 VSUBS 0.009394f
C351 B.n311 VSUBS 0.009394f
C352 B.n312 VSUBS 0.00525f
C353 B.n313 VSUBS 0.009394f
C354 B.n314 VSUBS 0.009394f
C355 B.n315 VSUBS 0.009394f
C356 B.n316 VSUBS 0.009394f
C357 B.n317 VSUBS 0.009394f
C358 B.n318 VSUBS 0.009394f
C359 B.n319 VSUBS 0.009394f
C360 B.n320 VSUBS 0.009394f
C361 B.n321 VSUBS 0.009394f
C362 B.n322 VSUBS 0.009394f
C363 B.n323 VSUBS 0.009394f
C364 B.n324 VSUBS 0.009394f
C365 B.n325 VSUBS 0.00525f
C366 B.n326 VSUBS 0.021766f
C367 B.n327 VSUBS 0.008842f
C368 B.n328 VSUBS 0.009394f
C369 B.n329 VSUBS 0.009394f
C370 B.n330 VSUBS 0.009394f
C371 B.n331 VSUBS 0.009394f
C372 B.n332 VSUBS 0.009394f
C373 B.n333 VSUBS 0.009394f
C374 B.n334 VSUBS 0.009394f
C375 B.n335 VSUBS 0.009394f
C376 B.n336 VSUBS 0.009394f
C377 B.n337 VSUBS 0.009394f
C378 B.n338 VSUBS 0.009394f
C379 B.n339 VSUBS 0.009394f
C380 B.n340 VSUBS 0.009394f
C381 B.n341 VSUBS 0.009394f
C382 B.n342 VSUBS 0.009394f
C383 B.n343 VSUBS 0.009394f
C384 B.n344 VSUBS 0.022048f
C385 B.n345 VSUBS 0.02078f
C386 B.n346 VSUBS 0.02078f
C387 B.n347 VSUBS 0.009394f
C388 B.n348 VSUBS 0.009394f
C389 B.n349 VSUBS 0.009394f
C390 B.n350 VSUBS 0.009394f
C391 B.n351 VSUBS 0.009394f
C392 B.n352 VSUBS 0.009394f
C393 B.n353 VSUBS 0.009394f
C394 B.n354 VSUBS 0.009394f
C395 B.n355 VSUBS 0.009394f
C396 B.n356 VSUBS 0.009394f
C397 B.n357 VSUBS 0.009394f
C398 B.n358 VSUBS 0.009394f
C399 B.n359 VSUBS 0.009394f
C400 B.n360 VSUBS 0.009394f
C401 B.n361 VSUBS 0.009394f
C402 B.n362 VSUBS 0.009394f
C403 B.n363 VSUBS 0.009394f
C404 B.n364 VSUBS 0.009394f
C405 B.n365 VSUBS 0.009394f
C406 B.n366 VSUBS 0.009394f
C407 B.n367 VSUBS 0.009394f
C408 B.n368 VSUBS 0.009394f
C409 B.n369 VSUBS 0.009394f
C410 B.n370 VSUBS 0.009394f
C411 B.n371 VSUBS 0.009394f
C412 B.n372 VSUBS 0.009394f
C413 B.n373 VSUBS 0.009394f
C414 B.n374 VSUBS 0.009394f
C415 B.n375 VSUBS 0.009394f
C416 B.n376 VSUBS 0.009394f
C417 B.n377 VSUBS 0.009394f
C418 B.n378 VSUBS 0.009394f
C419 B.n379 VSUBS 0.009394f
C420 B.n380 VSUBS 0.009394f
C421 B.n381 VSUBS 0.009394f
C422 B.n382 VSUBS 0.009394f
C423 B.n383 VSUBS 0.009394f
C424 B.n384 VSUBS 0.009394f
C425 B.n385 VSUBS 0.009394f
C426 B.n386 VSUBS 0.009394f
C427 B.n387 VSUBS 0.009394f
C428 B.n388 VSUBS 0.009394f
C429 B.n389 VSUBS 0.009394f
C430 B.n390 VSUBS 0.009394f
C431 B.n391 VSUBS 0.021272f
C432 VDD1.n0 VSUBS 0.019612f
C433 VDD1.n1 VSUBS 0.050655f
C434 VDD1.t1 VSUBS 0.05081f
C435 VDD1.n2 VSUBS 0.049483f
C436 VDD1.n3 VSUBS 0.01456f
C437 VDD1.n4 VSUBS 0.009445f
C438 VDD1.n5 VSUBS 0.119507f
C439 VDD1.n6 VSUBS 0.041285f
C440 VDD1.n7 VSUBS 0.019612f
C441 VDD1.n8 VSUBS 0.050655f
C442 VDD1.t0 VSUBS 0.05081f
C443 VDD1.n9 VSUBS 0.049483f
C444 VDD1.n10 VSUBS 0.01456f
C445 VDD1.n11 VSUBS 0.009445f
C446 VDD1.n12 VSUBS 0.119507f
C447 VDD1.n13 VSUBS 0.360189f
C448 VP.t0 VSUBS 2.37766f
C449 VP.t1 VSUBS 1.33997f
C450 VP.n0 VSUBS 3.70011f
C451 VDD2.n0 VSUBS 0.020095f
C452 VDD2.n1 VSUBS 0.051903f
C453 VDD2.t1 VSUBS 0.052062f
C454 VDD2.n2 VSUBS 0.050702f
C455 VDD2.n3 VSUBS 0.014919f
C456 VDD2.n4 VSUBS 0.009678f
C457 VDD2.n5 VSUBS 0.122451f
C458 VDD2.n6 VSUBS 0.336157f
C459 VDD2.n7 VSUBS 0.020095f
C460 VDD2.n8 VSUBS 0.051903f
C461 VDD2.t0 VSUBS 0.052062f
C462 VDD2.n9 VSUBS 0.050702f
C463 VDD2.n10 VSUBS 0.014919f
C464 VDD2.n11 VSUBS 0.009678f
C465 VDD2.n12 VSUBS 0.122451f
C466 VDD2.n13 VSUBS 0.040815f
C467 VDD2.n14 VSUBS 1.53596f
C468 VTAIL.n0 VSUBS 0.024501f
C469 VTAIL.n1 VSUBS 0.063283f
C470 VTAIL.t3 VSUBS 0.063476f
C471 VTAIL.n2 VSUBS 0.061818f
C472 VTAIL.n3 VSUBS 0.018189f
C473 VTAIL.n4 VSUBS 0.011799f
C474 VTAIL.n5 VSUBS 0.149297f
C475 VTAIL.n6 VSUBS 0.034584f
C476 VTAIL.n7 VSUBS 0.983895f
C477 VTAIL.n8 VSUBS 0.024501f
C478 VTAIL.n9 VSUBS 0.063283f
C479 VTAIL.t1 VSUBS 0.063476f
C480 VTAIL.n10 VSUBS 0.061818f
C481 VTAIL.n11 VSUBS 0.018189f
C482 VTAIL.n12 VSUBS 0.011799f
C483 VTAIL.n13 VSUBS 0.149297f
C484 VTAIL.n14 VSUBS 0.034584f
C485 VTAIL.n15 VSUBS 1.0365f
C486 VTAIL.n16 VSUBS 0.024501f
C487 VTAIL.n17 VSUBS 0.063283f
C488 VTAIL.t0 VSUBS 0.063476f
C489 VTAIL.n18 VSUBS 0.061818f
C490 VTAIL.n19 VSUBS 0.018189f
C491 VTAIL.n20 VSUBS 0.011799f
C492 VTAIL.n21 VSUBS 0.149297f
C493 VTAIL.n22 VSUBS 0.034584f
C494 VTAIL.n23 VSUBS 0.809602f
C495 VTAIL.n24 VSUBS 0.024501f
C496 VTAIL.n25 VSUBS 0.063283f
C497 VTAIL.t2 VSUBS 0.063476f
C498 VTAIL.n26 VSUBS 0.061818f
C499 VTAIL.n27 VSUBS 0.018189f
C500 VTAIL.n28 VSUBS 0.011799f
C501 VTAIL.n29 VSUBS 0.149297f
C502 VTAIL.n30 VSUBS 0.034584f
C503 VTAIL.n31 VSUBS 0.715517f
C504 VN.t0 VSUBS 1.28026f
C505 VN.t1 VSUBS 2.265f
.ends

