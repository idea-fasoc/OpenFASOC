* NGSPICE file created from diff_pair_sample_0687.ext - technology: sky130A

.subckt diff_pair_sample_0687 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VN.t0 VDD2.t1 B.t8 sky130_fd_pr__nfet_01v8 ad=1.03785 pd=6.62 as=1.03785 ps=6.62 w=6.29 l=3.29
X1 VTAIL.t3 VP.t0 VDD1.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=1.03785 pd=6.62 as=1.03785 ps=6.62 w=6.29 l=3.29
X2 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=2.4531 pd=13.36 as=0 ps=0 w=6.29 l=3.29
X3 VTAIL.t6 VP.t1 VDD1.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=1.03785 pd=6.62 as=1.03785 ps=6.62 w=6.29 l=3.29
X4 VDD1.t7 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.4531 pd=13.36 as=1.03785 ps=6.62 w=6.29 l=3.29
X5 VDD2.t2 VN.t1 VTAIL.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=1.03785 pd=6.62 as=2.4531 ps=13.36 w=6.29 l=3.29
X6 VDD2.t5 VN.t2 VTAIL.t16 B.t0 sky130_fd_pr__nfet_01v8 ad=1.03785 pd=6.62 as=1.03785 ps=6.62 w=6.29 l=3.29
X7 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=2.4531 pd=13.36 as=0 ps=0 w=6.29 l=3.29
X8 VTAIL.t4 VP.t3 VDD1.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=1.03785 pd=6.62 as=1.03785 ps=6.62 w=6.29 l=3.29
X9 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=2.4531 pd=13.36 as=0 ps=0 w=6.29 l=3.29
X10 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.4531 pd=13.36 as=0 ps=0 w=6.29 l=3.29
X11 VTAIL.t8 VP.t4 VDD1.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=1.03785 pd=6.62 as=1.03785 ps=6.62 w=6.29 l=3.29
X12 VDD2.t3 VN.t3 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=1.03785 pd=6.62 as=2.4531 ps=13.36 w=6.29 l=3.29
X13 VTAIL.t14 VN.t4 VDD2.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.03785 pd=6.62 as=1.03785 ps=6.62 w=6.29 l=3.29
X14 VTAIL.t13 VN.t5 VDD2.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=1.03785 pd=6.62 as=1.03785 ps=6.62 w=6.29 l=3.29
X15 VDD1.t4 VP.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.03785 pd=6.62 as=1.03785 ps=6.62 w=6.29 l=3.29
X16 VTAIL.t12 VN.t6 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=1.03785 pd=6.62 as=1.03785 ps=6.62 w=6.29 l=3.29
X17 VDD1.t3 VP.t6 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.03785 pd=6.62 as=2.4531 ps=13.36 w=6.29 l=3.29
X18 VDD1.t2 VP.t7 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.4531 pd=13.36 as=1.03785 ps=6.62 w=6.29 l=3.29
X19 VDD2.t9 VN.t7 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=2.4531 pd=13.36 as=1.03785 ps=6.62 w=6.29 l=3.29
X20 VDD1.t1 VP.t8 VTAIL.t19 B.t9 sky130_fd_pr__nfet_01v8 ad=1.03785 pd=6.62 as=2.4531 ps=13.36 w=6.29 l=3.29
X21 VDD2.t8 VN.t8 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=1.03785 pd=6.62 as=1.03785 ps=6.62 w=6.29 l=3.29
X22 VDD2.t6 VN.t9 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.4531 pd=13.36 as=1.03785 ps=6.62 w=6.29 l=3.29
X23 VDD1.t0 VP.t9 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.03785 pd=6.62 as=1.03785 ps=6.62 w=6.29 l=3.29
R0 VN.n96 VN.n95 161.3
R1 VN.n94 VN.n50 161.3
R2 VN.n93 VN.n92 161.3
R3 VN.n91 VN.n51 161.3
R4 VN.n90 VN.n89 161.3
R5 VN.n88 VN.n52 161.3
R6 VN.n87 VN.n86 161.3
R7 VN.n85 VN.n84 161.3
R8 VN.n83 VN.n54 161.3
R9 VN.n82 VN.n81 161.3
R10 VN.n80 VN.n55 161.3
R11 VN.n79 VN.n78 161.3
R12 VN.n77 VN.n56 161.3
R13 VN.n76 VN.n75 161.3
R14 VN.n74 VN.n57 161.3
R15 VN.n73 VN.n72 161.3
R16 VN.n71 VN.n58 161.3
R17 VN.n70 VN.n69 161.3
R18 VN.n68 VN.n59 161.3
R19 VN.n67 VN.n66 161.3
R20 VN.n65 VN.n60 161.3
R21 VN.n64 VN.n63 161.3
R22 VN.n47 VN.n46 161.3
R23 VN.n45 VN.n1 161.3
R24 VN.n44 VN.n43 161.3
R25 VN.n42 VN.n2 161.3
R26 VN.n41 VN.n40 161.3
R27 VN.n39 VN.n3 161.3
R28 VN.n38 VN.n37 161.3
R29 VN.n36 VN.n35 161.3
R30 VN.n34 VN.n5 161.3
R31 VN.n33 VN.n32 161.3
R32 VN.n31 VN.n6 161.3
R33 VN.n30 VN.n29 161.3
R34 VN.n28 VN.n7 161.3
R35 VN.n27 VN.n26 161.3
R36 VN.n25 VN.n8 161.3
R37 VN.n24 VN.n23 161.3
R38 VN.n22 VN.n9 161.3
R39 VN.n21 VN.n20 161.3
R40 VN.n19 VN.n10 161.3
R41 VN.n18 VN.n17 161.3
R42 VN.n16 VN.n11 161.3
R43 VN.n15 VN.n14 161.3
R44 VN.n62 VN.t3 78.5415
R45 VN.n13 VN.t9 78.5415
R46 VN.n48 VN.n0 78.3232
R47 VN.n97 VN.n49 78.3232
R48 VN.n13 VN.n12 68.6407
R49 VN.n62 VN.n61 68.6407
R50 VN.n21 VN.n10 56.5193
R51 VN.n29 VN.n6 56.5193
R52 VN.n70 VN.n59 56.5193
R53 VN.n78 VN.n55 56.5193
R54 VN VN.n97 52.7707
R55 VN.n40 VN.n2 47.2923
R56 VN.n89 VN.n51 47.2923
R57 VN.n8 VN.t2 46.0762
R58 VN.n12 VN.t5 46.0762
R59 VN.n4 VN.t4 46.0762
R60 VN.n0 VN.t1 46.0762
R61 VN.n57 VN.t8 46.0762
R62 VN.n61 VN.t6 46.0762
R63 VN.n53 VN.t0 46.0762
R64 VN.n49 VN.t7 46.0762
R65 VN.n44 VN.n2 33.6945
R66 VN.n93 VN.n51 33.6945
R67 VN.n16 VN.n15 24.4675
R68 VN.n17 VN.n16 24.4675
R69 VN.n17 VN.n10 24.4675
R70 VN.n22 VN.n21 24.4675
R71 VN.n23 VN.n22 24.4675
R72 VN.n23 VN.n8 24.4675
R73 VN.n27 VN.n8 24.4675
R74 VN.n28 VN.n27 24.4675
R75 VN.n29 VN.n28 24.4675
R76 VN.n33 VN.n6 24.4675
R77 VN.n34 VN.n33 24.4675
R78 VN.n35 VN.n34 24.4675
R79 VN.n39 VN.n38 24.4675
R80 VN.n40 VN.n39 24.4675
R81 VN.n45 VN.n44 24.4675
R82 VN.n46 VN.n45 24.4675
R83 VN.n66 VN.n59 24.4675
R84 VN.n66 VN.n65 24.4675
R85 VN.n65 VN.n64 24.4675
R86 VN.n78 VN.n77 24.4675
R87 VN.n77 VN.n76 24.4675
R88 VN.n76 VN.n57 24.4675
R89 VN.n72 VN.n57 24.4675
R90 VN.n72 VN.n71 24.4675
R91 VN.n71 VN.n70 24.4675
R92 VN.n89 VN.n88 24.4675
R93 VN.n88 VN.n87 24.4675
R94 VN.n84 VN.n83 24.4675
R95 VN.n83 VN.n82 24.4675
R96 VN.n82 VN.n55 24.4675
R97 VN.n95 VN.n94 24.4675
R98 VN.n94 VN.n93 24.4675
R99 VN.n38 VN.n4 18.5954
R100 VN.n87 VN.n53 18.5954
R101 VN.n46 VN.n0 11.7447
R102 VN.n95 VN.n49 11.7447
R103 VN.n15 VN.n12 5.87258
R104 VN.n35 VN.n4 5.87258
R105 VN.n64 VN.n61 5.87258
R106 VN.n84 VN.n53 5.87258
R107 VN.n14 VN.n13 4.31092
R108 VN.n63 VN.n62 4.31092
R109 VN.n97 VN.n96 0.354971
R110 VN.n48 VN.n47 0.354971
R111 VN VN.n48 0.26696
R112 VN.n96 VN.n50 0.189894
R113 VN.n92 VN.n50 0.189894
R114 VN.n92 VN.n91 0.189894
R115 VN.n91 VN.n90 0.189894
R116 VN.n90 VN.n52 0.189894
R117 VN.n86 VN.n52 0.189894
R118 VN.n86 VN.n85 0.189894
R119 VN.n85 VN.n54 0.189894
R120 VN.n81 VN.n54 0.189894
R121 VN.n81 VN.n80 0.189894
R122 VN.n80 VN.n79 0.189894
R123 VN.n79 VN.n56 0.189894
R124 VN.n75 VN.n56 0.189894
R125 VN.n75 VN.n74 0.189894
R126 VN.n74 VN.n73 0.189894
R127 VN.n73 VN.n58 0.189894
R128 VN.n69 VN.n58 0.189894
R129 VN.n69 VN.n68 0.189894
R130 VN.n68 VN.n67 0.189894
R131 VN.n67 VN.n60 0.189894
R132 VN.n63 VN.n60 0.189894
R133 VN.n14 VN.n11 0.189894
R134 VN.n18 VN.n11 0.189894
R135 VN.n19 VN.n18 0.189894
R136 VN.n20 VN.n19 0.189894
R137 VN.n20 VN.n9 0.189894
R138 VN.n24 VN.n9 0.189894
R139 VN.n25 VN.n24 0.189894
R140 VN.n26 VN.n25 0.189894
R141 VN.n26 VN.n7 0.189894
R142 VN.n30 VN.n7 0.189894
R143 VN.n31 VN.n30 0.189894
R144 VN.n32 VN.n31 0.189894
R145 VN.n32 VN.n5 0.189894
R146 VN.n36 VN.n5 0.189894
R147 VN.n37 VN.n36 0.189894
R148 VN.n37 VN.n3 0.189894
R149 VN.n41 VN.n3 0.189894
R150 VN.n42 VN.n41 0.189894
R151 VN.n43 VN.n42 0.189894
R152 VN.n43 VN.n1 0.189894
R153 VN.n47 VN.n1 0.189894
R154 VDD2.n1 VDD2.t6 71.5069
R155 VDD2.n4 VDD2.t9 68.3863
R156 VDD2.n3 VDD2.n2 67.5234
R157 VDD2 VDD2.n7 67.5206
R158 VDD2.n6 VDD2.n5 65.2385
R159 VDD2.n1 VDD2.n0 65.2383
R160 VDD2.n4 VDD2.n3 43.961
R161 VDD2.n7 VDD2.t0 3.14835
R162 VDD2.n7 VDD2.t3 3.14835
R163 VDD2.n5 VDD2.t1 3.14835
R164 VDD2.n5 VDD2.t8 3.14835
R165 VDD2.n2 VDD2.t7 3.14835
R166 VDD2.n2 VDD2.t2 3.14835
R167 VDD2.n0 VDD2.t4 3.14835
R168 VDD2.n0 VDD2.t5 3.14835
R169 VDD2.n6 VDD2.n4 3.12119
R170 VDD2 VDD2.n6 0.838862
R171 VDD2.n3 VDD2.n1 0.725326
R172 VTAIL.n11 VTAIL.t15 51.7075
R173 VTAIL.n16 VTAIL.t19 51.7074
R174 VTAIL.n17 VTAIL.t17 51.7074
R175 VTAIL.n2 VTAIL.t7 51.7074
R176 VTAIL.n15 VTAIL.n14 48.5597
R177 VTAIL.n13 VTAIL.n12 48.5597
R178 VTAIL.n10 VTAIL.n9 48.5597
R179 VTAIL.n8 VTAIL.n7 48.5597
R180 VTAIL.n19 VTAIL.n18 48.5595
R181 VTAIL.n1 VTAIL.n0 48.5595
R182 VTAIL.n4 VTAIL.n3 48.5595
R183 VTAIL.n6 VTAIL.n5 48.5595
R184 VTAIL.n8 VTAIL.n6 24.0307
R185 VTAIL.n17 VTAIL.n16 20.91
R186 VTAIL.n18 VTAIL.t16 3.14835
R187 VTAIL.n18 VTAIL.t14 3.14835
R188 VTAIL.n0 VTAIL.t9 3.14835
R189 VTAIL.n0 VTAIL.t13 3.14835
R190 VTAIL.n3 VTAIL.t2 3.14835
R191 VTAIL.n3 VTAIL.t4 3.14835
R192 VTAIL.n5 VTAIL.t1 3.14835
R193 VTAIL.n5 VTAIL.t8 3.14835
R194 VTAIL.n14 VTAIL.t0 3.14835
R195 VTAIL.n14 VTAIL.t3 3.14835
R196 VTAIL.n12 VTAIL.t5 3.14835
R197 VTAIL.n12 VTAIL.t6 3.14835
R198 VTAIL.n9 VTAIL.t10 3.14835
R199 VTAIL.n9 VTAIL.t12 3.14835
R200 VTAIL.n7 VTAIL.t11 3.14835
R201 VTAIL.n7 VTAIL.t18 3.14835
R202 VTAIL.n10 VTAIL.n8 3.12119
R203 VTAIL.n11 VTAIL.n10 3.12119
R204 VTAIL.n15 VTAIL.n13 3.12119
R205 VTAIL.n16 VTAIL.n15 3.12119
R206 VTAIL.n6 VTAIL.n4 3.12119
R207 VTAIL.n4 VTAIL.n2 3.12119
R208 VTAIL.n19 VTAIL.n17 3.12119
R209 VTAIL VTAIL.n1 2.39921
R210 VTAIL.n13 VTAIL.n11 2.03067
R211 VTAIL.n2 VTAIL.n1 2.03067
R212 VTAIL VTAIL.n19 0.722483
R213 B.n884 B.n883 585
R214 B.n885 B.n884 585
R215 B.n280 B.n161 585
R216 B.n279 B.n278 585
R217 B.n277 B.n276 585
R218 B.n275 B.n274 585
R219 B.n273 B.n272 585
R220 B.n271 B.n270 585
R221 B.n269 B.n268 585
R222 B.n267 B.n266 585
R223 B.n265 B.n264 585
R224 B.n263 B.n262 585
R225 B.n261 B.n260 585
R226 B.n259 B.n258 585
R227 B.n257 B.n256 585
R228 B.n255 B.n254 585
R229 B.n253 B.n252 585
R230 B.n251 B.n250 585
R231 B.n249 B.n248 585
R232 B.n247 B.n246 585
R233 B.n245 B.n244 585
R234 B.n243 B.n242 585
R235 B.n241 B.n240 585
R236 B.n239 B.n238 585
R237 B.n237 B.n236 585
R238 B.n235 B.n234 585
R239 B.n233 B.n232 585
R240 B.n231 B.n230 585
R241 B.n229 B.n228 585
R242 B.n227 B.n226 585
R243 B.n225 B.n224 585
R244 B.n223 B.n222 585
R245 B.n221 B.n220 585
R246 B.n219 B.n218 585
R247 B.n217 B.n216 585
R248 B.n214 B.n213 585
R249 B.n212 B.n211 585
R250 B.n210 B.n209 585
R251 B.n208 B.n207 585
R252 B.n206 B.n205 585
R253 B.n204 B.n203 585
R254 B.n202 B.n201 585
R255 B.n200 B.n199 585
R256 B.n198 B.n197 585
R257 B.n196 B.n195 585
R258 B.n194 B.n193 585
R259 B.n192 B.n191 585
R260 B.n190 B.n189 585
R261 B.n188 B.n187 585
R262 B.n186 B.n185 585
R263 B.n184 B.n183 585
R264 B.n182 B.n181 585
R265 B.n180 B.n179 585
R266 B.n178 B.n177 585
R267 B.n176 B.n175 585
R268 B.n174 B.n173 585
R269 B.n172 B.n171 585
R270 B.n170 B.n169 585
R271 B.n168 B.n167 585
R272 B.n130 B.n129 585
R273 B.n882 B.n131 585
R274 B.n886 B.n131 585
R275 B.n881 B.n880 585
R276 B.n880 B.n127 585
R277 B.n879 B.n126 585
R278 B.n892 B.n126 585
R279 B.n878 B.n125 585
R280 B.n893 B.n125 585
R281 B.n877 B.n124 585
R282 B.n894 B.n124 585
R283 B.n876 B.n875 585
R284 B.n875 B.n120 585
R285 B.n874 B.n119 585
R286 B.n900 B.n119 585
R287 B.n873 B.n118 585
R288 B.n901 B.n118 585
R289 B.n872 B.n117 585
R290 B.n902 B.n117 585
R291 B.n871 B.n870 585
R292 B.n870 B.n113 585
R293 B.n869 B.n112 585
R294 B.n908 B.n112 585
R295 B.n868 B.n111 585
R296 B.n909 B.n111 585
R297 B.n867 B.n110 585
R298 B.n910 B.n110 585
R299 B.n866 B.n865 585
R300 B.n865 B.n106 585
R301 B.n864 B.n105 585
R302 B.n916 B.n105 585
R303 B.n863 B.n104 585
R304 B.n917 B.n104 585
R305 B.n862 B.n103 585
R306 B.n918 B.n103 585
R307 B.n861 B.n860 585
R308 B.n860 B.n99 585
R309 B.n859 B.n98 585
R310 B.n924 B.n98 585
R311 B.n858 B.n97 585
R312 B.n925 B.n97 585
R313 B.n857 B.n96 585
R314 B.n926 B.n96 585
R315 B.n856 B.n855 585
R316 B.n855 B.n92 585
R317 B.n854 B.n91 585
R318 B.n932 B.n91 585
R319 B.n853 B.n90 585
R320 B.n933 B.n90 585
R321 B.n852 B.n89 585
R322 B.n934 B.n89 585
R323 B.n851 B.n850 585
R324 B.n850 B.n85 585
R325 B.n849 B.n84 585
R326 B.n940 B.n84 585
R327 B.n848 B.n83 585
R328 B.n941 B.n83 585
R329 B.n847 B.n82 585
R330 B.n942 B.n82 585
R331 B.n846 B.n845 585
R332 B.n845 B.n78 585
R333 B.n844 B.n77 585
R334 B.n948 B.n77 585
R335 B.n843 B.n76 585
R336 B.n949 B.n76 585
R337 B.n842 B.n75 585
R338 B.n950 B.n75 585
R339 B.n841 B.n840 585
R340 B.n840 B.n74 585
R341 B.n839 B.n70 585
R342 B.n956 B.n70 585
R343 B.n838 B.n69 585
R344 B.n957 B.n69 585
R345 B.n837 B.n68 585
R346 B.n958 B.n68 585
R347 B.n836 B.n835 585
R348 B.n835 B.n64 585
R349 B.n834 B.n63 585
R350 B.n964 B.n63 585
R351 B.n833 B.n62 585
R352 B.n965 B.n62 585
R353 B.n832 B.n61 585
R354 B.n966 B.n61 585
R355 B.n831 B.n830 585
R356 B.n830 B.n57 585
R357 B.n829 B.n56 585
R358 B.n972 B.n56 585
R359 B.n828 B.n55 585
R360 B.n973 B.n55 585
R361 B.n827 B.n54 585
R362 B.n974 B.n54 585
R363 B.n826 B.n825 585
R364 B.n825 B.n50 585
R365 B.n824 B.n49 585
R366 B.n980 B.n49 585
R367 B.n823 B.n48 585
R368 B.n981 B.n48 585
R369 B.n822 B.n47 585
R370 B.n982 B.n47 585
R371 B.n821 B.n820 585
R372 B.n820 B.n43 585
R373 B.n819 B.n42 585
R374 B.n988 B.n42 585
R375 B.n818 B.n41 585
R376 B.n989 B.n41 585
R377 B.n817 B.n40 585
R378 B.n990 B.n40 585
R379 B.n816 B.n815 585
R380 B.n815 B.n36 585
R381 B.n814 B.n35 585
R382 B.n996 B.n35 585
R383 B.n813 B.n34 585
R384 B.n997 B.n34 585
R385 B.n812 B.n33 585
R386 B.n998 B.n33 585
R387 B.n811 B.n810 585
R388 B.n810 B.n29 585
R389 B.n809 B.n28 585
R390 B.n1004 B.n28 585
R391 B.n808 B.n27 585
R392 B.n1005 B.n27 585
R393 B.n807 B.n26 585
R394 B.n1006 B.n26 585
R395 B.n806 B.n805 585
R396 B.n805 B.n22 585
R397 B.n804 B.n21 585
R398 B.n1012 B.n21 585
R399 B.n803 B.n20 585
R400 B.n1013 B.n20 585
R401 B.n802 B.n19 585
R402 B.n1014 B.n19 585
R403 B.n801 B.n800 585
R404 B.n800 B.n18 585
R405 B.n799 B.n14 585
R406 B.n1020 B.n14 585
R407 B.n798 B.n13 585
R408 B.n1021 B.n13 585
R409 B.n797 B.n12 585
R410 B.n1022 B.n12 585
R411 B.n796 B.n795 585
R412 B.n795 B.n8 585
R413 B.n794 B.n7 585
R414 B.n1028 B.n7 585
R415 B.n793 B.n6 585
R416 B.n1029 B.n6 585
R417 B.n792 B.n5 585
R418 B.n1030 B.n5 585
R419 B.n791 B.n790 585
R420 B.n790 B.n4 585
R421 B.n789 B.n281 585
R422 B.n789 B.n788 585
R423 B.n779 B.n282 585
R424 B.n283 B.n282 585
R425 B.n781 B.n780 585
R426 B.n782 B.n781 585
R427 B.n778 B.n288 585
R428 B.n288 B.n287 585
R429 B.n777 B.n776 585
R430 B.n776 B.n775 585
R431 B.n290 B.n289 585
R432 B.n768 B.n290 585
R433 B.n767 B.n766 585
R434 B.n769 B.n767 585
R435 B.n765 B.n295 585
R436 B.n295 B.n294 585
R437 B.n764 B.n763 585
R438 B.n763 B.n762 585
R439 B.n297 B.n296 585
R440 B.n298 B.n297 585
R441 B.n755 B.n754 585
R442 B.n756 B.n755 585
R443 B.n753 B.n303 585
R444 B.n303 B.n302 585
R445 B.n752 B.n751 585
R446 B.n751 B.n750 585
R447 B.n305 B.n304 585
R448 B.n306 B.n305 585
R449 B.n743 B.n742 585
R450 B.n744 B.n743 585
R451 B.n741 B.n311 585
R452 B.n311 B.n310 585
R453 B.n740 B.n739 585
R454 B.n739 B.n738 585
R455 B.n313 B.n312 585
R456 B.n314 B.n313 585
R457 B.n731 B.n730 585
R458 B.n732 B.n731 585
R459 B.n729 B.n319 585
R460 B.n319 B.n318 585
R461 B.n728 B.n727 585
R462 B.n727 B.n726 585
R463 B.n321 B.n320 585
R464 B.n322 B.n321 585
R465 B.n719 B.n718 585
R466 B.n720 B.n719 585
R467 B.n717 B.n327 585
R468 B.n327 B.n326 585
R469 B.n716 B.n715 585
R470 B.n715 B.n714 585
R471 B.n329 B.n328 585
R472 B.n330 B.n329 585
R473 B.n707 B.n706 585
R474 B.n708 B.n707 585
R475 B.n705 B.n334 585
R476 B.n338 B.n334 585
R477 B.n704 B.n703 585
R478 B.n703 B.n702 585
R479 B.n336 B.n335 585
R480 B.n337 B.n336 585
R481 B.n695 B.n694 585
R482 B.n696 B.n695 585
R483 B.n693 B.n343 585
R484 B.n343 B.n342 585
R485 B.n692 B.n691 585
R486 B.n691 B.n690 585
R487 B.n345 B.n344 585
R488 B.n346 B.n345 585
R489 B.n683 B.n682 585
R490 B.n684 B.n683 585
R491 B.n681 B.n351 585
R492 B.n351 B.n350 585
R493 B.n680 B.n679 585
R494 B.n679 B.n678 585
R495 B.n353 B.n352 585
R496 B.n671 B.n353 585
R497 B.n670 B.n669 585
R498 B.n672 B.n670 585
R499 B.n668 B.n358 585
R500 B.n358 B.n357 585
R501 B.n667 B.n666 585
R502 B.n666 B.n665 585
R503 B.n360 B.n359 585
R504 B.n361 B.n360 585
R505 B.n658 B.n657 585
R506 B.n659 B.n658 585
R507 B.n656 B.n366 585
R508 B.n366 B.n365 585
R509 B.n655 B.n654 585
R510 B.n654 B.n653 585
R511 B.n368 B.n367 585
R512 B.n369 B.n368 585
R513 B.n646 B.n645 585
R514 B.n647 B.n646 585
R515 B.n644 B.n374 585
R516 B.n374 B.n373 585
R517 B.n643 B.n642 585
R518 B.n642 B.n641 585
R519 B.n376 B.n375 585
R520 B.n377 B.n376 585
R521 B.n634 B.n633 585
R522 B.n635 B.n634 585
R523 B.n632 B.n382 585
R524 B.n382 B.n381 585
R525 B.n631 B.n630 585
R526 B.n630 B.n629 585
R527 B.n384 B.n383 585
R528 B.n385 B.n384 585
R529 B.n622 B.n621 585
R530 B.n623 B.n622 585
R531 B.n620 B.n390 585
R532 B.n390 B.n389 585
R533 B.n619 B.n618 585
R534 B.n618 B.n617 585
R535 B.n392 B.n391 585
R536 B.n393 B.n392 585
R537 B.n610 B.n609 585
R538 B.n611 B.n610 585
R539 B.n608 B.n398 585
R540 B.n398 B.n397 585
R541 B.n607 B.n606 585
R542 B.n606 B.n605 585
R543 B.n400 B.n399 585
R544 B.n401 B.n400 585
R545 B.n598 B.n597 585
R546 B.n599 B.n598 585
R547 B.n596 B.n406 585
R548 B.n406 B.n405 585
R549 B.n595 B.n594 585
R550 B.n594 B.n593 585
R551 B.n408 B.n407 585
R552 B.n409 B.n408 585
R553 B.n586 B.n585 585
R554 B.n587 B.n586 585
R555 B.n584 B.n414 585
R556 B.n414 B.n413 585
R557 B.n583 B.n582 585
R558 B.n582 B.n581 585
R559 B.n416 B.n415 585
R560 B.n417 B.n416 585
R561 B.n574 B.n573 585
R562 B.n575 B.n574 585
R563 B.n420 B.n419 585
R564 B.n458 B.n457 585
R565 B.n459 B.n455 585
R566 B.n455 B.n421 585
R567 B.n461 B.n460 585
R568 B.n463 B.n454 585
R569 B.n466 B.n465 585
R570 B.n467 B.n453 585
R571 B.n469 B.n468 585
R572 B.n471 B.n452 585
R573 B.n474 B.n473 585
R574 B.n475 B.n451 585
R575 B.n477 B.n476 585
R576 B.n479 B.n450 585
R577 B.n482 B.n481 585
R578 B.n483 B.n449 585
R579 B.n485 B.n484 585
R580 B.n487 B.n448 585
R581 B.n490 B.n489 585
R582 B.n491 B.n447 585
R583 B.n493 B.n492 585
R584 B.n495 B.n446 585
R585 B.n498 B.n497 585
R586 B.n499 B.n445 585
R587 B.n501 B.n500 585
R588 B.n503 B.n444 585
R589 B.n506 B.n505 585
R590 B.n507 B.n440 585
R591 B.n509 B.n508 585
R592 B.n511 B.n439 585
R593 B.n514 B.n513 585
R594 B.n515 B.n438 585
R595 B.n517 B.n516 585
R596 B.n519 B.n437 585
R597 B.n522 B.n521 585
R598 B.n524 B.n434 585
R599 B.n526 B.n525 585
R600 B.n528 B.n433 585
R601 B.n531 B.n530 585
R602 B.n532 B.n432 585
R603 B.n534 B.n533 585
R604 B.n536 B.n431 585
R605 B.n539 B.n538 585
R606 B.n540 B.n430 585
R607 B.n542 B.n541 585
R608 B.n544 B.n429 585
R609 B.n547 B.n546 585
R610 B.n548 B.n428 585
R611 B.n550 B.n549 585
R612 B.n552 B.n427 585
R613 B.n555 B.n554 585
R614 B.n556 B.n426 585
R615 B.n558 B.n557 585
R616 B.n560 B.n425 585
R617 B.n563 B.n562 585
R618 B.n564 B.n424 585
R619 B.n566 B.n565 585
R620 B.n568 B.n423 585
R621 B.n571 B.n570 585
R622 B.n572 B.n422 585
R623 B.n577 B.n576 585
R624 B.n576 B.n575 585
R625 B.n578 B.n418 585
R626 B.n418 B.n417 585
R627 B.n580 B.n579 585
R628 B.n581 B.n580 585
R629 B.n412 B.n411 585
R630 B.n413 B.n412 585
R631 B.n589 B.n588 585
R632 B.n588 B.n587 585
R633 B.n590 B.n410 585
R634 B.n410 B.n409 585
R635 B.n592 B.n591 585
R636 B.n593 B.n592 585
R637 B.n404 B.n403 585
R638 B.n405 B.n404 585
R639 B.n601 B.n600 585
R640 B.n600 B.n599 585
R641 B.n602 B.n402 585
R642 B.n402 B.n401 585
R643 B.n604 B.n603 585
R644 B.n605 B.n604 585
R645 B.n396 B.n395 585
R646 B.n397 B.n396 585
R647 B.n613 B.n612 585
R648 B.n612 B.n611 585
R649 B.n614 B.n394 585
R650 B.n394 B.n393 585
R651 B.n616 B.n615 585
R652 B.n617 B.n616 585
R653 B.n388 B.n387 585
R654 B.n389 B.n388 585
R655 B.n625 B.n624 585
R656 B.n624 B.n623 585
R657 B.n626 B.n386 585
R658 B.n386 B.n385 585
R659 B.n628 B.n627 585
R660 B.n629 B.n628 585
R661 B.n380 B.n379 585
R662 B.n381 B.n380 585
R663 B.n637 B.n636 585
R664 B.n636 B.n635 585
R665 B.n638 B.n378 585
R666 B.n378 B.n377 585
R667 B.n640 B.n639 585
R668 B.n641 B.n640 585
R669 B.n372 B.n371 585
R670 B.n373 B.n372 585
R671 B.n649 B.n648 585
R672 B.n648 B.n647 585
R673 B.n650 B.n370 585
R674 B.n370 B.n369 585
R675 B.n652 B.n651 585
R676 B.n653 B.n652 585
R677 B.n364 B.n363 585
R678 B.n365 B.n364 585
R679 B.n661 B.n660 585
R680 B.n660 B.n659 585
R681 B.n662 B.n362 585
R682 B.n362 B.n361 585
R683 B.n664 B.n663 585
R684 B.n665 B.n664 585
R685 B.n356 B.n355 585
R686 B.n357 B.n356 585
R687 B.n674 B.n673 585
R688 B.n673 B.n672 585
R689 B.n675 B.n354 585
R690 B.n671 B.n354 585
R691 B.n677 B.n676 585
R692 B.n678 B.n677 585
R693 B.n349 B.n348 585
R694 B.n350 B.n349 585
R695 B.n686 B.n685 585
R696 B.n685 B.n684 585
R697 B.n687 B.n347 585
R698 B.n347 B.n346 585
R699 B.n689 B.n688 585
R700 B.n690 B.n689 585
R701 B.n341 B.n340 585
R702 B.n342 B.n341 585
R703 B.n698 B.n697 585
R704 B.n697 B.n696 585
R705 B.n699 B.n339 585
R706 B.n339 B.n337 585
R707 B.n701 B.n700 585
R708 B.n702 B.n701 585
R709 B.n333 B.n332 585
R710 B.n338 B.n333 585
R711 B.n710 B.n709 585
R712 B.n709 B.n708 585
R713 B.n711 B.n331 585
R714 B.n331 B.n330 585
R715 B.n713 B.n712 585
R716 B.n714 B.n713 585
R717 B.n325 B.n324 585
R718 B.n326 B.n325 585
R719 B.n722 B.n721 585
R720 B.n721 B.n720 585
R721 B.n723 B.n323 585
R722 B.n323 B.n322 585
R723 B.n725 B.n724 585
R724 B.n726 B.n725 585
R725 B.n317 B.n316 585
R726 B.n318 B.n317 585
R727 B.n734 B.n733 585
R728 B.n733 B.n732 585
R729 B.n735 B.n315 585
R730 B.n315 B.n314 585
R731 B.n737 B.n736 585
R732 B.n738 B.n737 585
R733 B.n309 B.n308 585
R734 B.n310 B.n309 585
R735 B.n746 B.n745 585
R736 B.n745 B.n744 585
R737 B.n747 B.n307 585
R738 B.n307 B.n306 585
R739 B.n749 B.n748 585
R740 B.n750 B.n749 585
R741 B.n301 B.n300 585
R742 B.n302 B.n301 585
R743 B.n758 B.n757 585
R744 B.n757 B.n756 585
R745 B.n759 B.n299 585
R746 B.n299 B.n298 585
R747 B.n761 B.n760 585
R748 B.n762 B.n761 585
R749 B.n293 B.n292 585
R750 B.n294 B.n293 585
R751 B.n771 B.n770 585
R752 B.n770 B.n769 585
R753 B.n772 B.n291 585
R754 B.n768 B.n291 585
R755 B.n774 B.n773 585
R756 B.n775 B.n774 585
R757 B.n286 B.n285 585
R758 B.n287 B.n286 585
R759 B.n784 B.n783 585
R760 B.n783 B.n782 585
R761 B.n785 B.n284 585
R762 B.n284 B.n283 585
R763 B.n787 B.n786 585
R764 B.n788 B.n787 585
R765 B.n2 B.n0 585
R766 B.n4 B.n2 585
R767 B.n3 B.n1 585
R768 B.n1029 B.n3 585
R769 B.n1027 B.n1026 585
R770 B.n1028 B.n1027 585
R771 B.n1025 B.n9 585
R772 B.n9 B.n8 585
R773 B.n1024 B.n1023 585
R774 B.n1023 B.n1022 585
R775 B.n11 B.n10 585
R776 B.n1021 B.n11 585
R777 B.n1019 B.n1018 585
R778 B.n1020 B.n1019 585
R779 B.n1017 B.n15 585
R780 B.n18 B.n15 585
R781 B.n1016 B.n1015 585
R782 B.n1015 B.n1014 585
R783 B.n17 B.n16 585
R784 B.n1013 B.n17 585
R785 B.n1011 B.n1010 585
R786 B.n1012 B.n1011 585
R787 B.n1009 B.n23 585
R788 B.n23 B.n22 585
R789 B.n1008 B.n1007 585
R790 B.n1007 B.n1006 585
R791 B.n25 B.n24 585
R792 B.n1005 B.n25 585
R793 B.n1003 B.n1002 585
R794 B.n1004 B.n1003 585
R795 B.n1001 B.n30 585
R796 B.n30 B.n29 585
R797 B.n1000 B.n999 585
R798 B.n999 B.n998 585
R799 B.n32 B.n31 585
R800 B.n997 B.n32 585
R801 B.n995 B.n994 585
R802 B.n996 B.n995 585
R803 B.n993 B.n37 585
R804 B.n37 B.n36 585
R805 B.n992 B.n991 585
R806 B.n991 B.n990 585
R807 B.n39 B.n38 585
R808 B.n989 B.n39 585
R809 B.n987 B.n986 585
R810 B.n988 B.n987 585
R811 B.n985 B.n44 585
R812 B.n44 B.n43 585
R813 B.n984 B.n983 585
R814 B.n983 B.n982 585
R815 B.n46 B.n45 585
R816 B.n981 B.n46 585
R817 B.n979 B.n978 585
R818 B.n980 B.n979 585
R819 B.n977 B.n51 585
R820 B.n51 B.n50 585
R821 B.n976 B.n975 585
R822 B.n975 B.n974 585
R823 B.n53 B.n52 585
R824 B.n973 B.n53 585
R825 B.n971 B.n970 585
R826 B.n972 B.n971 585
R827 B.n969 B.n58 585
R828 B.n58 B.n57 585
R829 B.n968 B.n967 585
R830 B.n967 B.n966 585
R831 B.n60 B.n59 585
R832 B.n965 B.n60 585
R833 B.n963 B.n962 585
R834 B.n964 B.n963 585
R835 B.n961 B.n65 585
R836 B.n65 B.n64 585
R837 B.n960 B.n959 585
R838 B.n959 B.n958 585
R839 B.n67 B.n66 585
R840 B.n957 B.n67 585
R841 B.n955 B.n954 585
R842 B.n956 B.n955 585
R843 B.n953 B.n71 585
R844 B.n74 B.n71 585
R845 B.n952 B.n951 585
R846 B.n951 B.n950 585
R847 B.n73 B.n72 585
R848 B.n949 B.n73 585
R849 B.n947 B.n946 585
R850 B.n948 B.n947 585
R851 B.n945 B.n79 585
R852 B.n79 B.n78 585
R853 B.n944 B.n943 585
R854 B.n943 B.n942 585
R855 B.n81 B.n80 585
R856 B.n941 B.n81 585
R857 B.n939 B.n938 585
R858 B.n940 B.n939 585
R859 B.n937 B.n86 585
R860 B.n86 B.n85 585
R861 B.n936 B.n935 585
R862 B.n935 B.n934 585
R863 B.n88 B.n87 585
R864 B.n933 B.n88 585
R865 B.n931 B.n930 585
R866 B.n932 B.n931 585
R867 B.n929 B.n93 585
R868 B.n93 B.n92 585
R869 B.n928 B.n927 585
R870 B.n927 B.n926 585
R871 B.n95 B.n94 585
R872 B.n925 B.n95 585
R873 B.n923 B.n922 585
R874 B.n924 B.n923 585
R875 B.n921 B.n100 585
R876 B.n100 B.n99 585
R877 B.n920 B.n919 585
R878 B.n919 B.n918 585
R879 B.n102 B.n101 585
R880 B.n917 B.n102 585
R881 B.n915 B.n914 585
R882 B.n916 B.n915 585
R883 B.n913 B.n107 585
R884 B.n107 B.n106 585
R885 B.n912 B.n911 585
R886 B.n911 B.n910 585
R887 B.n109 B.n108 585
R888 B.n909 B.n109 585
R889 B.n907 B.n906 585
R890 B.n908 B.n907 585
R891 B.n905 B.n114 585
R892 B.n114 B.n113 585
R893 B.n904 B.n903 585
R894 B.n903 B.n902 585
R895 B.n116 B.n115 585
R896 B.n901 B.n116 585
R897 B.n899 B.n898 585
R898 B.n900 B.n899 585
R899 B.n897 B.n121 585
R900 B.n121 B.n120 585
R901 B.n896 B.n895 585
R902 B.n895 B.n894 585
R903 B.n123 B.n122 585
R904 B.n893 B.n123 585
R905 B.n891 B.n890 585
R906 B.n892 B.n891 585
R907 B.n889 B.n128 585
R908 B.n128 B.n127 585
R909 B.n888 B.n887 585
R910 B.n887 B.n886 585
R911 B.n1032 B.n1031 585
R912 B.n1031 B.n1030 585
R913 B.n576 B.n420 516.524
R914 B.n887 B.n130 516.524
R915 B.n574 B.n422 516.524
R916 B.n884 B.n131 516.524
R917 B.n885 B.n160 256.663
R918 B.n885 B.n159 256.663
R919 B.n885 B.n158 256.663
R920 B.n885 B.n157 256.663
R921 B.n885 B.n156 256.663
R922 B.n885 B.n155 256.663
R923 B.n885 B.n154 256.663
R924 B.n885 B.n153 256.663
R925 B.n885 B.n152 256.663
R926 B.n885 B.n151 256.663
R927 B.n885 B.n150 256.663
R928 B.n885 B.n149 256.663
R929 B.n885 B.n148 256.663
R930 B.n885 B.n147 256.663
R931 B.n885 B.n146 256.663
R932 B.n885 B.n145 256.663
R933 B.n885 B.n144 256.663
R934 B.n885 B.n143 256.663
R935 B.n885 B.n142 256.663
R936 B.n885 B.n141 256.663
R937 B.n885 B.n140 256.663
R938 B.n885 B.n139 256.663
R939 B.n885 B.n138 256.663
R940 B.n885 B.n137 256.663
R941 B.n885 B.n136 256.663
R942 B.n885 B.n135 256.663
R943 B.n885 B.n134 256.663
R944 B.n885 B.n133 256.663
R945 B.n885 B.n132 256.663
R946 B.n456 B.n421 256.663
R947 B.n462 B.n421 256.663
R948 B.n464 B.n421 256.663
R949 B.n470 B.n421 256.663
R950 B.n472 B.n421 256.663
R951 B.n478 B.n421 256.663
R952 B.n480 B.n421 256.663
R953 B.n486 B.n421 256.663
R954 B.n488 B.n421 256.663
R955 B.n494 B.n421 256.663
R956 B.n496 B.n421 256.663
R957 B.n502 B.n421 256.663
R958 B.n504 B.n421 256.663
R959 B.n510 B.n421 256.663
R960 B.n512 B.n421 256.663
R961 B.n518 B.n421 256.663
R962 B.n520 B.n421 256.663
R963 B.n527 B.n421 256.663
R964 B.n529 B.n421 256.663
R965 B.n535 B.n421 256.663
R966 B.n537 B.n421 256.663
R967 B.n543 B.n421 256.663
R968 B.n545 B.n421 256.663
R969 B.n551 B.n421 256.663
R970 B.n553 B.n421 256.663
R971 B.n559 B.n421 256.663
R972 B.n561 B.n421 256.663
R973 B.n567 B.n421 256.663
R974 B.n569 B.n421 256.663
R975 B.n435 B.t14 254.97
R976 B.n441 B.t18 254.97
R977 B.n165 B.t10 254.97
R978 B.n162 B.t21 254.97
R979 B.n576 B.n418 163.367
R980 B.n580 B.n418 163.367
R981 B.n580 B.n412 163.367
R982 B.n588 B.n412 163.367
R983 B.n588 B.n410 163.367
R984 B.n592 B.n410 163.367
R985 B.n592 B.n404 163.367
R986 B.n600 B.n404 163.367
R987 B.n600 B.n402 163.367
R988 B.n604 B.n402 163.367
R989 B.n604 B.n396 163.367
R990 B.n612 B.n396 163.367
R991 B.n612 B.n394 163.367
R992 B.n616 B.n394 163.367
R993 B.n616 B.n388 163.367
R994 B.n624 B.n388 163.367
R995 B.n624 B.n386 163.367
R996 B.n628 B.n386 163.367
R997 B.n628 B.n380 163.367
R998 B.n636 B.n380 163.367
R999 B.n636 B.n378 163.367
R1000 B.n640 B.n378 163.367
R1001 B.n640 B.n372 163.367
R1002 B.n648 B.n372 163.367
R1003 B.n648 B.n370 163.367
R1004 B.n652 B.n370 163.367
R1005 B.n652 B.n364 163.367
R1006 B.n660 B.n364 163.367
R1007 B.n660 B.n362 163.367
R1008 B.n664 B.n362 163.367
R1009 B.n664 B.n356 163.367
R1010 B.n673 B.n356 163.367
R1011 B.n673 B.n354 163.367
R1012 B.n677 B.n354 163.367
R1013 B.n677 B.n349 163.367
R1014 B.n685 B.n349 163.367
R1015 B.n685 B.n347 163.367
R1016 B.n689 B.n347 163.367
R1017 B.n689 B.n341 163.367
R1018 B.n697 B.n341 163.367
R1019 B.n697 B.n339 163.367
R1020 B.n701 B.n339 163.367
R1021 B.n701 B.n333 163.367
R1022 B.n709 B.n333 163.367
R1023 B.n709 B.n331 163.367
R1024 B.n713 B.n331 163.367
R1025 B.n713 B.n325 163.367
R1026 B.n721 B.n325 163.367
R1027 B.n721 B.n323 163.367
R1028 B.n725 B.n323 163.367
R1029 B.n725 B.n317 163.367
R1030 B.n733 B.n317 163.367
R1031 B.n733 B.n315 163.367
R1032 B.n737 B.n315 163.367
R1033 B.n737 B.n309 163.367
R1034 B.n745 B.n309 163.367
R1035 B.n745 B.n307 163.367
R1036 B.n749 B.n307 163.367
R1037 B.n749 B.n301 163.367
R1038 B.n757 B.n301 163.367
R1039 B.n757 B.n299 163.367
R1040 B.n761 B.n299 163.367
R1041 B.n761 B.n293 163.367
R1042 B.n770 B.n293 163.367
R1043 B.n770 B.n291 163.367
R1044 B.n774 B.n291 163.367
R1045 B.n774 B.n286 163.367
R1046 B.n783 B.n286 163.367
R1047 B.n783 B.n284 163.367
R1048 B.n787 B.n284 163.367
R1049 B.n787 B.n2 163.367
R1050 B.n1031 B.n2 163.367
R1051 B.n1031 B.n3 163.367
R1052 B.n1027 B.n3 163.367
R1053 B.n1027 B.n9 163.367
R1054 B.n1023 B.n9 163.367
R1055 B.n1023 B.n11 163.367
R1056 B.n1019 B.n11 163.367
R1057 B.n1019 B.n15 163.367
R1058 B.n1015 B.n15 163.367
R1059 B.n1015 B.n17 163.367
R1060 B.n1011 B.n17 163.367
R1061 B.n1011 B.n23 163.367
R1062 B.n1007 B.n23 163.367
R1063 B.n1007 B.n25 163.367
R1064 B.n1003 B.n25 163.367
R1065 B.n1003 B.n30 163.367
R1066 B.n999 B.n30 163.367
R1067 B.n999 B.n32 163.367
R1068 B.n995 B.n32 163.367
R1069 B.n995 B.n37 163.367
R1070 B.n991 B.n37 163.367
R1071 B.n991 B.n39 163.367
R1072 B.n987 B.n39 163.367
R1073 B.n987 B.n44 163.367
R1074 B.n983 B.n44 163.367
R1075 B.n983 B.n46 163.367
R1076 B.n979 B.n46 163.367
R1077 B.n979 B.n51 163.367
R1078 B.n975 B.n51 163.367
R1079 B.n975 B.n53 163.367
R1080 B.n971 B.n53 163.367
R1081 B.n971 B.n58 163.367
R1082 B.n967 B.n58 163.367
R1083 B.n967 B.n60 163.367
R1084 B.n963 B.n60 163.367
R1085 B.n963 B.n65 163.367
R1086 B.n959 B.n65 163.367
R1087 B.n959 B.n67 163.367
R1088 B.n955 B.n67 163.367
R1089 B.n955 B.n71 163.367
R1090 B.n951 B.n71 163.367
R1091 B.n951 B.n73 163.367
R1092 B.n947 B.n73 163.367
R1093 B.n947 B.n79 163.367
R1094 B.n943 B.n79 163.367
R1095 B.n943 B.n81 163.367
R1096 B.n939 B.n81 163.367
R1097 B.n939 B.n86 163.367
R1098 B.n935 B.n86 163.367
R1099 B.n935 B.n88 163.367
R1100 B.n931 B.n88 163.367
R1101 B.n931 B.n93 163.367
R1102 B.n927 B.n93 163.367
R1103 B.n927 B.n95 163.367
R1104 B.n923 B.n95 163.367
R1105 B.n923 B.n100 163.367
R1106 B.n919 B.n100 163.367
R1107 B.n919 B.n102 163.367
R1108 B.n915 B.n102 163.367
R1109 B.n915 B.n107 163.367
R1110 B.n911 B.n107 163.367
R1111 B.n911 B.n109 163.367
R1112 B.n907 B.n109 163.367
R1113 B.n907 B.n114 163.367
R1114 B.n903 B.n114 163.367
R1115 B.n903 B.n116 163.367
R1116 B.n899 B.n116 163.367
R1117 B.n899 B.n121 163.367
R1118 B.n895 B.n121 163.367
R1119 B.n895 B.n123 163.367
R1120 B.n891 B.n123 163.367
R1121 B.n891 B.n128 163.367
R1122 B.n887 B.n128 163.367
R1123 B.n457 B.n455 163.367
R1124 B.n461 B.n455 163.367
R1125 B.n465 B.n463 163.367
R1126 B.n469 B.n453 163.367
R1127 B.n473 B.n471 163.367
R1128 B.n477 B.n451 163.367
R1129 B.n481 B.n479 163.367
R1130 B.n485 B.n449 163.367
R1131 B.n489 B.n487 163.367
R1132 B.n493 B.n447 163.367
R1133 B.n497 B.n495 163.367
R1134 B.n501 B.n445 163.367
R1135 B.n505 B.n503 163.367
R1136 B.n509 B.n440 163.367
R1137 B.n513 B.n511 163.367
R1138 B.n517 B.n438 163.367
R1139 B.n521 B.n519 163.367
R1140 B.n526 B.n434 163.367
R1141 B.n530 B.n528 163.367
R1142 B.n534 B.n432 163.367
R1143 B.n538 B.n536 163.367
R1144 B.n542 B.n430 163.367
R1145 B.n546 B.n544 163.367
R1146 B.n550 B.n428 163.367
R1147 B.n554 B.n552 163.367
R1148 B.n558 B.n426 163.367
R1149 B.n562 B.n560 163.367
R1150 B.n566 B.n424 163.367
R1151 B.n570 B.n568 163.367
R1152 B.n574 B.n416 163.367
R1153 B.n582 B.n416 163.367
R1154 B.n582 B.n414 163.367
R1155 B.n586 B.n414 163.367
R1156 B.n586 B.n408 163.367
R1157 B.n594 B.n408 163.367
R1158 B.n594 B.n406 163.367
R1159 B.n598 B.n406 163.367
R1160 B.n598 B.n400 163.367
R1161 B.n606 B.n400 163.367
R1162 B.n606 B.n398 163.367
R1163 B.n610 B.n398 163.367
R1164 B.n610 B.n392 163.367
R1165 B.n618 B.n392 163.367
R1166 B.n618 B.n390 163.367
R1167 B.n622 B.n390 163.367
R1168 B.n622 B.n384 163.367
R1169 B.n630 B.n384 163.367
R1170 B.n630 B.n382 163.367
R1171 B.n634 B.n382 163.367
R1172 B.n634 B.n376 163.367
R1173 B.n642 B.n376 163.367
R1174 B.n642 B.n374 163.367
R1175 B.n646 B.n374 163.367
R1176 B.n646 B.n368 163.367
R1177 B.n654 B.n368 163.367
R1178 B.n654 B.n366 163.367
R1179 B.n658 B.n366 163.367
R1180 B.n658 B.n360 163.367
R1181 B.n666 B.n360 163.367
R1182 B.n666 B.n358 163.367
R1183 B.n670 B.n358 163.367
R1184 B.n670 B.n353 163.367
R1185 B.n679 B.n353 163.367
R1186 B.n679 B.n351 163.367
R1187 B.n683 B.n351 163.367
R1188 B.n683 B.n345 163.367
R1189 B.n691 B.n345 163.367
R1190 B.n691 B.n343 163.367
R1191 B.n695 B.n343 163.367
R1192 B.n695 B.n336 163.367
R1193 B.n703 B.n336 163.367
R1194 B.n703 B.n334 163.367
R1195 B.n707 B.n334 163.367
R1196 B.n707 B.n329 163.367
R1197 B.n715 B.n329 163.367
R1198 B.n715 B.n327 163.367
R1199 B.n719 B.n327 163.367
R1200 B.n719 B.n321 163.367
R1201 B.n727 B.n321 163.367
R1202 B.n727 B.n319 163.367
R1203 B.n731 B.n319 163.367
R1204 B.n731 B.n313 163.367
R1205 B.n739 B.n313 163.367
R1206 B.n739 B.n311 163.367
R1207 B.n743 B.n311 163.367
R1208 B.n743 B.n305 163.367
R1209 B.n751 B.n305 163.367
R1210 B.n751 B.n303 163.367
R1211 B.n755 B.n303 163.367
R1212 B.n755 B.n297 163.367
R1213 B.n763 B.n297 163.367
R1214 B.n763 B.n295 163.367
R1215 B.n767 B.n295 163.367
R1216 B.n767 B.n290 163.367
R1217 B.n776 B.n290 163.367
R1218 B.n776 B.n288 163.367
R1219 B.n781 B.n288 163.367
R1220 B.n781 B.n282 163.367
R1221 B.n789 B.n282 163.367
R1222 B.n790 B.n789 163.367
R1223 B.n790 B.n5 163.367
R1224 B.n6 B.n5 163.367
R1225 B.n7 B.n6 163.367
R1226 B.n795 B.n7 163.367
R1227 B.n795 B.n12 163.367
R1228 B.n13 B.n12 163.367
R1229 B.n14 B.n13 163.367
R1230 B.n800 B.n14 163.367
R1231 B.n800 B.n19 163.367
R1232 B.n20 B.n19 163.367
R1233 B.n21 B.n20 163.367
R1234 B.n805 B.n21 163.367
R1235 B.n805 B.n26 163.367
R1236 B.n27 B.n26 163.367
R1237 B.n28 B.n27 163.367
R1238 B.n810 B.n28 163.367
R1239 B.n810 B.n33 163.367
R1240 B.n34 B.n33 163.367
R1241 B.n35 B.n34 163.367
R1242 B.n815 B.n35 163.367
R1243 B.n815 B.n40 163.367
R1244 B.n41 B.n40 163.367
R1245 B.n42 B.n41 163.367
R1246 B.n820 B.n42 163.367
R1247 B.n820 B.n47 163.367
R1248 B.n48 B.n47 163.367
R1249 B.n49 B.n48 163.367
R1250 B.n825 B.n49 163.367
R1251 B.n825 B.n54 163.367
R1252 B.n55 B.n54 163.367
R1253 B.n56 B.n55 163.367
R1254 B.n830 B.n56 163.367
R1255 B.n830 B.n61 163.367
R1256 B.n62 B.n61 163.367
R1257 B.n63 B.n62 163.367
R1258 B.n835 B.n63 163.367
R1259 B.n835 B.n68 163.367
R1260 B.n69 B.n68 163.367
R1261 B.n70 B.n69 163.367
R1262 B.n840 B.n70 163.367
R1263 B.n840 B.n75 163.367
R1264 B.n76 B.n75 163.367
R1265 B.n77 B.n76 163.367
R1266 B.n845 B.n77 163.367
R1267 B.n845 B.n82 163.367
R1268 B.n83 B.n82 163.367
R1269 B.n84 B.n83 163.367
R1270 B.n850 B.n84 163.367
R1271 B.n850 B.n89 163.367
R1272 B.n90 B.n89 163.367
R1273 B.n91 B.n90 163.367
R1274 B.n855 B.n91 163.367
R1275 B.n855 B.n96 163.367
R1276 B.n97 B.n96 163.367
R1277 B.n98 B.n97 163.367
R1278 B.n860 B.n98 163.367
R1279 B.n860 B.n103 163.367
R1280 B.n104 B.n103 163.367
R1281 B.n105 B.n104 163.367
R1282 B.n865 B.n105 163.367
R1283 B.n865 B.n110 163.367
R1284 B.n111 B.n110 163.367
R1285 B.n112 B.n111 163.367
R1286 B.n870 B.n112 163.367
R1287 B.n870 B.n117 163.367
R1288 B.n118 B.n117 163.367
R1289 B.n119 B.n118 163.367
R1290 B.n875 B.n119 163.367
R1291 B.n875 B.n124 163.367
R1292 B.n125 B.n124 163.367
R1293 B.n126 B.n125 163.367
R1294 B.n880 B.n126 163.367
R1295 B.n880 B.n131 163.367
R1296 B.n169 B.n168 163.367
R1297 B.n173 B.n172 163.367
R1298 B.n177 B.n176 163.367
R1299 B.n181 B.n180 163.367
R1300 B.n185 B.n184 163.367
R1301 B.n189 B.n188 163.367
R1302 B.n193 B.n192 163.367
R1303 B.n197 B.n196 163.367
R1304 B.n201 B.n200 163.367
R1305 B.n205 B.n204 163.367
R1306 B.n209 B.n208 163.367
R1307 B.n213 B.n212 163.367
R1308 B.n218 B.n217 163.367
R1309 B.n222 B.n221 163.367
R1310 B.n226 B.n225 163.367
R1311 B.n230 B.n229 163.367
R1312 B.n234 B.n233 163.367
R1313 B.n238 B.n237 163.367
R1314 B.n242 B.n241 163.367
R1315 B.n246 B.n245 163.367
R1316 B.n250 B.n249 163.367
R1317 B.n254 B.n253 163.367
R1318 B.n258 B.n257 163.367
R1319 B.n262 B.n261 163.367
R1320 B.n266 B.n265 163.367
R1321 B.n270 B.n269 163.367
R1322 B.n274 B.n273 163.367
R1323 B.n278 B.n277 163.367
R1324 B.n884 B.n161 163.367
R1325 B.n435 B.t17 142.794
R1326 B.n162 B.t22 142.794
R1327 B.n441 B.t20 142.787
R1328 B.n165 B.t12 142.787
R1329 B.n575 B.n421 116.992
R1330 B.n886 B.n885 116.992
R1331 B.n436 B.t16 72.5879
R1332 B.n163 B.t23 72.5879
R1333 B.n442 B.t19 72.5812
R1334 B.n166 B.t13 72.5812
R1335 B.n456 B.n420 71.676
R1336 B.n462 B.n461 71.676
R1337 B.n465 B.n464 71.676
R1338 B.n470 B.n469 71.676
R1339 B.n473 B.n472 71.676
R1340 B.n478 B.n477 71.676
R1341 B.n481 B.n480 71.676
R1342 B.n486 B.n485 71.676
R1343 B.n489 B.n488 71.676
R1344 B.n494 B.n493 71.676
R1345 B.n497 B.n496 71.676
R1346 B.n502 B.n501 71.676
R1347 B.n505 B.n504 71.676
R1348 B.n510 B.n509 71.676
R1349 B.n513 B.n512 71.676
R1350 B.n518 B.n517 71.676
R1351 B.n521 B.n520 71.676
R1352 B.n527 B.n526 71.676
R1353 B.n530 B.n529 71.676
R1354 B.n535 B.n534 71.676
R1355 B.n538 B.n537 71.676
R1356 B.n543 B.n542 71.676
R1357 B.n546 B.n545 71.676
R1358 B.n551 B.n550 71.676
R1359 B.n554 B.n553 71.676
R1360 B.n559 B.n558 71.676
R1361 B.n562 B.n561 71.676
R1362 B.n567 B.n566 71.676
R1363 B.n570 B.n569 71.676
R1364 B.n132 B.n130 71.676
R1365 B.n169 B.n133 71.676
R1366 B.n173 B.n134 71.676
R1367 B.n177 B.n135 71.676
R1368 B.n181 B.n136 71.676
R1369 B.n185 B.n137 71.676
R1370 B.n189 B.n138 71.676
R1371 B.n193 B.n139 71.676
R1372 B.n197 B.n140 71.676
R1373 B.n201 B.n141 71.676
R1374 B.n205 B.n142 71.676
R1375 B.n209 B.n143 71.676
R1376 B.n213 B.n144 71.676
R1377 B.n218 B.n145 71.676
R1378 B.n222 B.n146 71.676
R1379 B.n226 B.n147 71.676
R1380 B.n230 B.n148 71.676
R1381 B.n234 B.n149 71.676
R1382 B.n238 B.n150 71.676
R1383 B.n242 B.n151 71.676
R1384 B.n246 B.n152 71.676
R1385 B.n250 B.n153 71.676
R1386 B.n254 B.n154 71.676
R1387 B.n258 B.n155 71.676
R1388 B.n262 B.n156 71.676
R1389 B.n266 B.n157 71.676
R1390 B.n270 B.n158 71.676
R1391 B.n274 B.n159 71.676
R1392 B.n278 B.n160 71.676
R1393 B.n161 B.n160 71.676
R1394 B.n277 B.n159 71.676
R1395 B.n273 B.n158 71.676
R1396 B.n269 B.n157 71.676
R1397 B.n265 B.n156 71.676
R1398 B.n261 B.n155 71.676
R1399 B.n257 B.n154 71.676
R1400 B.n253 B.n153 71.676
R1401 B.n249 B.n152 71.676
R1402 B.n245 B.n151 71.676
R1403 B.n241 B.n150 71.676
R1404 B.n237 B.n149 71.676
R1405 B.n233 B.n148 71.676
R1406 B.n229 B.n147 71.676
R1407 B.n225 B.n146 71.676
R1408 B.n221 B.n145 71.676
R1409 B.n217 B.n144 71.676
R1410 B.n212 B.n143 71.676
R1411 B.n208 B.n142 71.676
R1412 B.n204 B.n141 71.676
R1413 B.n200 B.n140 71.676
R1414 B.n196 B.n139 71.676
R1415 B.n192 B.n138 71.676
R1416 B.n188 B.n137 71.676
R1417 B.n184 B.n136 71.676
R1418 B.n180 B.n135 71.676
R1419 B.n176 B.n134 71.676
R1420 B.n172 B.n133 71.676
R1421 B.n168 B.n132 71.676
R1422 B.n457 B.n456 71.676
R1423 B.n463 B.n462 71.676
R1424 B.n464 B.n453 71.676
R1425 B.n471 B.n470 71.676
R1426 B.n472 B.n451 71.676
R1427 B.n479 B.n478 71.676
R1428 B.n480 B.n449 71.676
R1429 B.n487 B.n486 71.676
R1430 B.n488 B.n447 71.676
R1431 B.n495 B.n494 71.676
R1432 B.n496 B.n445 71.676
R1433 B.n503 B.n502 71.676
R1434 B.n504 B.n440 71.676
R1435 B.n511 B.n510 71.676
R1436 B.n512 B.n438 71.676
R1437 B.n519 B.n518 71.676
R1438 B.n520 B.n434 71.676
R1439 B.n528 B.n527 71.676
R1440 B.n529 B.n432 71.676
R1441 B.n536 B.n535 71.676
R1442 B.n537 B.n430 71.676
R1443 B.n544 B.n543 71.676
R1444 B.n545 B.n428 71.676
R1445 B.n552 B.n551 71.676
R1446 B.n553 B.n426 71.676
R1447 B.n560 B.n559 71.676
R1448 B.n561 B.n424 71.676
R1449 B.n568 B.n567 71.676
R1450 B.n569 B.n422 71.676
R1451 B.n436 B.n435 70.2066
R1452 B.n442 B.n441 70.2066
R1453 B.n166 B.n165 70.2066
R1454 B.n163 B.n162 70.2066
R1455 B.n575 B.n417 64.6784
R1456 B.n581 B.n417 64.6784
R1457 B.n581 B.n413 64.6784
R1458 B.n587 B.n413 64.6784
R1459 B.n587 B.n409 64.6784
R1460 B.n593 B.n409 64.6784
R1461 B.n593 B.n405 64.6784
R1462 B.n599 B.n405 64.6784
R1463 B.n605 B.n401 64.6784
R1464 B.n605 B.n397 64.6784
R1465 B.n611 B.n397 64.6784
R1466 B.n611 B.n393 64.6784
R1467 B.n617 B.n393 64.6784
R1468 B.n617 B.n389 64.6784
R1469 B.n623 B.n389 64.6784
R1470 B.n623 B.n385 64.6784
R1471 B.n629 B.n385 64.6784
R1472 B.n629 B.n381 64.6784
R1473 B.n635 B.n381 64.6784
R1474 B.n635 B.n377 64.6784
R1475 B.n641 B.n377 64.6784
R1476 B.n647 B.n373 64.6784
R1477 B.n647 B.n369 64.6784
R1478 B.n653 B.n369 64.6784
R1479 B.n653 B.n365 64.6784
R1480 B.n659 B.n365 64.6784
R1481 B.n659 B.n361 64.6784
R1482 B.n665 B.n361 64.6784
R1483 B.n665 B.n357 64.6784
R1484 B.n672 B.n357 64.6784
R1485 B.n672 B.n671 64.6784
R1486 B.n678 B.n350 64.6784
R1487 B.n684 B.n350 64.6784
R1488 B.n684 B.n346 64.6784
R1489 B.n690 B.n346 64.6784
R1490 B.n690 B.n342 64.6784
R1491 B.n696 B.n342 64.6784
R1492 B.n696 B.n337 64.6784
R1493 B.n702 B.n337 64.6784
R1494 B.n702 B.n338 64.6784
R1495 B.n708 B.n330 64.6784
R1496 B.n714 B.n330 64.6784
R1497 B.n714 B.n326 64.6784
R1498 B.n720 B.n326 64.6784
R1499 B.n720 B.n322 64.6784
R1500 B.n726 B.n322 64.6784
R1501 B.n726 B.n318 64.6784
R1502 B.n732 B.n318 64.6784
R1503 B.n732 B.n314 64.6784
R1504 B.n738 B.n314 64.6784
R1505 B.n744 B.n310 64.6784
R1506 B.n744 B.n306 64.6784
R1507 B.n750 B.n306 64.6784
R1508 B.n750 B.n302 64.6784
R1509 B.n756 B.n302 64.6784
R1510 B.n756 B.n298 64.6784
R1511 B.n762 B.n298 64.6784
R1512 B.n762 B.n294 64.6784
R1513 B.n769 B.n294 64.6784
R1514 B.n769 B.n768 64.6784
R1515 B.n775 B.n287 64.6784
R1516 B.n782 B.n287 64.6784
R1517 B.n782 B.n283 64.6784
R1518 B.n788 B.n283 64.6784
R1519 B.n788 B.n4 64.6784
R1520 B.n1030 B.n4 64.6784
R1521 B.n1030 B.n1029 64.6784
R1522 B.n1029 B.n1028 64.6784
R1523 B.n1028 B.n8 64.6784
R1524 B.n1022 B.n8 64.6784
R1525 B.n1022 B.n1021 64.6784
R1526 B.n1021 B.n1020 64.6784
R1527 B.n1014 B.n18 64.6784
R1528 B.n1014 B.n1013 64.6784
R1529 B.n1013 B.n1012 64.6784
R1530 B.n1012 B.n22 64.6784
R1531 B.n1006 B.n22 64.6784
R1532 B.n1006 B.n1005 64.6784
R1533 B.n1005 B.n1004 64.6784
R1534 B.n1004 B.n29 64.6784
R1535 B.n998 B.n29 64.6784
R1536 B.n998 B.n997 64.6784
R1537 B.n996 B.n36 64.6784
R1538 B.n990 B.n36 64.6784
R1539 B.n990 B.n989 64.6784
R1540 B.n989 B.n988 64.6784
R1541 B.n988 B.n43 64.6784
R1542 B.n982 B.n43 64.6784
R1543 B.n982 B.n981 64.6784
R1544 B.n981 B.n980 64.6784
R1545 B.n980 B.n50 64.6784
R1546 B.n974 B.n50 64.6784
R1547 B.n973 B.n972 64.6784
R1548 B.n972 B.n57 64.6784
R1549 B.n966 B.n57 64.6784
R1550 B.n966 B.n965 64.6784
R1551 B.n965 B.n964 64.6784
R1552 B.n964 B.n64 64.6784
R1553 B.n958 B.n64 64.6784
R1554 B.n958 B.n957 64.6784
R1555 B.n957 B.n956 64.6784
R1556 B.n950 B.n74 64.6784
R1557 B.n950 B.n949 64.6784
R1558 B.n949 B.n948 64.6784
R1559 B.n948 B.n78 64.6784
R1560 B.n942 B.n78 64.6784
R1561 B.n942 B.n941 64.6784
R1562 B.n941 B.n940 64.6784
R1563 B.n940 B.n85 64.6784
R1564 B.n934 B.n85 64.6784
R1565 B.n934 B.n933 64.6784
R1566 B.n932 B.n92 64.6784
R1567 B.n926 B.n92 64.6784
R1568 B.n926 B.n925 64.6784
R1569 B.n925 B.n924 64.6784
R1570 B.n924 B.n99 64.6784
R1571 B.n918 B.n99 64.6784
R1572 B.n918 B.n917 64.6784
R1573 B.n917 B.n916 64.6784
R1574 B.n916 B.n106 64.6784
R1575 B.n910 B.n106 64.6784
R1576 B.n910 B.n909 64.6784
R1577 B.n909 B.n908 64.6784
R1578 B.n908 B.n113 64.6784
R1579 B.n902 B.n901 64.6784
R1580 B.n901 B.n900 64.6784
R1581 B.n900 B.n120 64.6784
R1582 B.n894 B.n120 64.6784
R1583 B.n894 B.n893 64.6784
R1584 B.n893 B.n892 64.6784
R1585 B.n892 B.n127 64.6784
R1586 B.n886 B.n127 64.6784
R1587 B.n775 B.t7 59.9227
R1588 B.n1020 B.t5 59.9227
R1589 B.n523 B.n436 59.5399
R1590 B.n443 B.n442 59.5399
R1591 B.n215 B.n166 59.5399
R1592 B.n164 B.n163 59.5399
R1593 B.n678 B.t8 56.1181
R1594 B.n956 B.t3 56.1181
R1595 B.n338 B.t2 50.4112
R1596 B.t0 B.n973 50.4112
R1597 B.n599 B.t15 40.8998
R1598 B.n902 B.t11 40.8998
R1599 B.t4 B.n310 37.0952
R1600 B.n997 B.t6 37.0952
R1601 B.n888 B.n129 33.5615
R1602 B.n883 B.n882 33.5615
R1603 B.n573 B.n572 33.5615
R1604 B.n577 B.n419 33.5615
R1605 B.t1 B.n373 33.2906
R1606 B.n933 B.t9 33.2906
R1607 B.n641 B.t1 31.3883
R1608 B.t9 B.n932 31.3883
R1609 B.n738 B.t4 27.5837
R1610 B.t6 B.n996 27.5837
R1611 B.t15 B.n401 23.7791
R1612 B.t11 B.n113 23.7791
R1613 B B.n1032 18.0485
R1614 B.n708 B.t2 14.2677
R1615 B.n974 B.t0 14.2677
R1616 B.n167 B.n129 10.6151
R1617 B.n170 B.n167 10.6151
R1618 B.n171 B.n170 10.6151
R1619 B.n174 B.n171 10.6151
R1620 B.n175 B.n174 10.6151
R1621 B.n178 B.n175 10.6151
R1622 B.n179 B.n178 10.6151
R1623 B.n182 B.n179 10.6151
R1624 B.n183 B.n182 10.6151
R1625 B.n186 B.n183 10.6151
R1626 B.n187 B.n186 10.6151
R1627 B.n190 B.n187 10.6151
R1628 B.n191 B.n190 10.6151
R1629 B.n194 B.n191 10.6151
R1630 B.n195 B.n194 10.6151
R1631 B.n198 B.n195 10.6151
R1632 B.n199 B.n198 10.6151
R1633 B.n202 B.n199 10.6151
R1634 B.n203 B.n202 10.6151
R1635 B.n206 B.n203 10.6151
R1636 B.n207 B.n206 10.6151
R1637 B.n210 B.n207 10.6151
R1638 B.n211 B.n210 10.6151
R1639 B.n214 B.n211 10.6151
R1640 B.n219 B.n216 10.6151
R1641 B.n220 B.n219 10.6151
R1642 B.n223 B.n220 10.6151
R1643 B.n224 B.n223 10.6151
R1644 B.n227 B.n224 10.6151
R1645 B.n228 B.n227 10.6151
R1646 B.n231 B.n228 10.6151
R1647 B.n232 B.n231 10.6151
R1648 B.n236 B.n235 10.6151
R1649 B.n239 B.n236 10.6151
R1650 B.n240 B.n239 10.6151
R1651 B.n243 B.n240 10.6151
R1652 B.n244 B.n243 10.6151
R1653 B.n247 B.n244 10.6151
R1654 B.n248 B.n247 10.6151
R1655 B.n251 B.n248 10.6151
R1656 B.n252 B.n251 10.6151
R1657 B.n255 B.n252 10.6151
R1658 B.n256 B.n255 10.6151
R1659 B.n259 B.n256 10.6151
R1660 B.n260 B.n259 10.6151
R1661 B.n263 B.n260 10.6151
R1662 B.n264 B.n263 10.6151
R1663 B.n267 B.n264 10.6151
R1664 B.n268 B.n267 10.6151
R1665 B.n271 B.n268 10.6151
R1666 B.n272 B.n271 10.6151
R1667 B.n275 B.n272 10.6151
R1668 B.n276 B.n275 10.6151
R1669 B.n279 B.n276 10.6151
R1670 B.n280 B.n279 10.6151
R1671 B.n883 B.n280 10.6151
R1672 B.n573 B.n415 10.6151
R1673 B.n583 B.n415 10.6151
R1674 B.n584 B.n583 10.6151
R1675 B.n585 B.n584 10.6151
R1676 B.n585 B.n407 10.6151
R1677 B.n595 B.n407 10.6151
R1678 B.n596 B.n595 10.6151
R1679 B.n597 B.n596 10.6151
R1680 B.n597 B.n399 10.6151
R1681 B.n607 B.n399 10.6151
R1682 B.n608 B.n607 10.6151
R1683 B.n609 B.n608 10.6151
R1684 B.n609 B.n391 10.6151
R1685 B.n619 B.n391 10.6151
R1686 B.n620 B.n619 10.6151
R1687 B.n621 B.n620 10.6151
R1688 B.n621 B.n383 10.6151
R1689 B.n631 B.n383 10.6151
R1690 B.n632 B.n631 10.6151
R1691 B.n633 B.n632 10.6151
R1692 B.n633 B.n375 10.6151
R1693 B.n643 B.n375 10.6151
R1694 B.n644 B.n643 10.6151
R1695 B.n645 B.n644 10.6151
R1696 B.n645 B.n367 10.6151
R1697 B.n655 B.n367 10.6151
R1698 B.n656 B.n655 10.6151
R1699 B.n657 B.n656 10.6151
R1700 B.n657 B.n359 10.6151
R1701 B.n667 B.n359 10.6151
R1702 B.n668 B.n667 10.6151
R1703 B.n669 B.n668 10.6151
R1704 B.n669 B.n352 10.6151
R1705 B.n680 B.n352 10.6151
R1706 B.n681 B.n680 10.6151
R1707 B.n682 B.n681 10.6151
R1708 B.n682 B.n344 10.6151
R1709 B.n692 B.n344 10.6151
R1710 B.n693 B.n692 10.6151
R1711 B.n694 B.n693 10.6151
R1712 B.n694 B.n335 10.6151
R1713 B.n704 B.n335 10.6151
R1714 B.n705 B.n704 10.6151
R1715 B.n706 B.n705 10.6151
R1716 B.n706 B.n328 10.6151
R1717 B.n716 B.n328 10.6151
R1718 B.n717 B.n716 10.6151
R1719 B.n718 B.n717 10.6151
R1720 B.n718 B.n320 10.6151
R1721 B.n728 B.n320 10.6151
R1722 B.n729 B.n728 10.6151
R1723 B.n730 B.n729 10.6151
R1724 B.n730 B.n312 10.6151
R1725 B.n740 B.n312 10.6151
R1726 B.n741 B.n740 10.6151
R1727 B.n742 B.n741 10.6151
R1728 B.n742 B.n304 10.6151
R1729 B.n752 B.n304 10.6151
R1730 B.n753 B.n752 10.6151
R1731 B.n754 B.n753 10.6151
R1732 B.n754 B.n296 10.6151
R1733 B.n764 B.n296 10.6151
R1734 B.n765 B.n764 10.6151
R1735 B.n766 B.n765 10.6151
R1736 B.n766 B.n289 10.6151
R1737 B.n777 B.n289 10.6151
R1738 B.n778 B.n777 10.6151
R1739 B.n780 B.n778 10.6151
R1740 B.n780 B.n779 10.6151
R1741 B.n779 B.n281 10.6151
R1742 B.n791 B.n281 10.6151
R1743 B.n792 B.n791 10.6151
R1744 B.n793 B.n792 10.6151
R1745 B.n794 B.n793 10.6151
R1746 B.n796 B.n794 10.6151
R1747 B.n797 B.n796 10.6151
R1748 B.n798 B.n797 10.6151
R1749 B.n799 B.n798 10.6151
R1750 B.n801 B.n799 10.6151
R1751 B.n802 B.n801 10.6151
R1752 B.n803 B.n802 10.6151
R1753 B.n804 B.n803 10.6151
R1754 B.n806 B.n804 10.6151
R1755 B.n807 B.n806 10.6151
R1756 B.n808 B.n807 10.6151
R1757 B.n809 B.n808 10.6151
R1758 B.n811 B.n809 10.6151
R1759 B.n812 B.n811 10.6151
R1760 B.n813 B.n812 10.6151
R1761 B.n814 B.n813 10.6151
R1762 B.n816 B.n814 10.6151
R1763 B.n817 B.n816 10.6151
R1764 B.n818 B.n817 10.6151
R1765 B.n819 B.n818 10.6151
R1766 B.n821 B.n819 10.6151
R1767 B.n822 B.n821 10.6151
R1768 B.n823 B.n822 10.6151
R1769 B.n824 B.n823 10.6151
R1770 B.n826 B.n824 10.6151
R1771 B.n827 B.n826 10.6151
R1772 B.n828 B.n827 10.6151
R1773 B.n829 B.n828 10.6151
R1774 B.n831 B.n829 10.6151
R1775 B.n832 B.n831 10.6151
R1776 B.n833 B.n832 10.6151
R1777 B.n834 B.n833 10.6151
R1778 B.n836 B.n834 10.6151
R1779 B.n837 B.n836 10.6151
R1780 B.n838 B.n837 10.6151
R1781 B.n839 B.n838 10.6151
R1782 B.n841 B.n839 10.6151
R1783 B.n842 B.n841 10.6151
R1784 B.n843 B.n842 10.6151
R1785 B.n844 B.n843 10.6151
R1786 B.n846 B.n844 10.6151
R1787 B.n847 B.n846 10.6151
R1788 B.n848 B.n847 10.6151
R1789 B.n849 B.n848 10.6151
R1790 B.n851 B.n849 10.6151
R1791 B.n852 B.n851 10.6151
R1792 B.n853 B.n852 10.6151
R1793 B.n854 B.n853 10.6151
R1794 B.n856 B.n854 10.6151
R1795 B.n857 B.n856 10.6151
R1796 B.n858 B.n857 10.6151
R1797 B.n859 B.n858 10.6151
R1798 B.n861 B.n859 10.6151
R1799 B.n862 B.n861 10.6151
R1800 B.n863 B.n862 10.6151
R1801 B.n864 B.n863 10.6151
R1802 B.n866 B.n864 10.6151
R1803 B.n867 B.n866 10.6151
R1804 B.n868 B.n867 10.6151
R1805 B.n869 B.n868 10.6151
R1806 B.n871 B.n869 10.6151
R1807 B.n872 B.n871 10.6151
R1808 B.n873 B.n872 10.6151
R1809 B.n874 B.n873 10.6151
R1810 B.n876 B.n874 10.6151
R1811 B.n877 B.n876 10.6151
R1812 B.n878 B.n877 10.6151
R1813 B.n879 B.n878 10.6151
R1814 B.n881 B.n879 10.6151
R1815 B.n882 B.n881 10.6151
R1816 B.n458 B.n419 10.6151
R1817 B.n459 B.n458 10.6151
R1818 B.n460 B.n459 10.6151
R1819 B.n460 B.n454 10.6151
R1820 B.n466 B.n454 10.6151
R1821 B.n467 B.n466 10.6151
R1822 B.n468 B.n467 10.6151
R1823 B.n468 B.n452 10.6151
R1824 B.n474 B.n452 10.6151
R1825 B.n475 B.n474 10.6151
R1826 B.n476 B.n475 10.6151
R1827 B.n476 B.n450 10.6151
R1828 B.n482 B.n450 10.6151
R1829 B.n483 B.n482 10.6151
R1830 B.n484 B.n483 10.6151
R1831 B.n484 B.n448 10.6151
R1832 B.n490 B.n448 10.6151
R1833 B.n491 B.n490 10.6151
R1834 B.n492 B.n491 10.6151
R1835 B.n492 B.n446 10.6151
R1836 B.n498 B.n446 10.6151
R1837 B.n499 B.n498 10.6151
R1838 B.n500 B.n499 10.6151
R1839 B.n500 B.n444 10.6151
R1840 B.n507 B.n506 10.6151
R1841 B.n508 B.n507 10.6151
R1842 B.n508 B.n439 10.6151
R1843 B.n514 B.n439 10.6151
R1844 B.n515 B.n514 10.6151
R1845 B.n516 B.n515 10.6151
R1846 B.n516 B.n437 10.6151
R1847 B.n522 B.n437 10.6151
R1848 B.n525 B.n524 10.6151
R1849 B.n525 B.n433 10.6151
R1850 B.n531 B.n433 10.6151
R1851 B.n532 B.n531 10.6151
R1852 B.n533 B.n532 10.6151
R1853 B.n533 B.n431 10.6151
R1854 B.n539 B.n431 10.6151
R1855 B.n540 B.n539 10.6151
R1856 B.n541 B.n540 10.6151
R1857 B.n541 B.n429 10.6151
R1858 B.n547 B.n429 10.6151
R1859 B.n548 B.n547 10.6151
R1860 B.n549 B.n548 10.6151
R1861 B.n549 B.n427 10.6151
R1862 B.n555 B.n427 10.6151
R1863 B.n556 B.n555 10.6151
R1864 B.n557 B.n556 10.6151
R1865 B.n557 B.n425 10.6151
R1866 B.n563 B.n425 10.6151
R1867 B.n564 B.n563 10.6151
R1868 B.n565 B.n564 10.6151
R1869 B.n565 B.n423 10.6151
R1870 B.n571 B.n423 10.6151
R1871 B.n572 B.n571 10.6151
R1872 B.n578 B.n577 10.6151
R1873 B.n579 B.n578 10.6151
R1874 B.n579 B.n411 10.6151
R1875 B.n589 B.n411 10.6151
R1876 B.n590 B.n589 10.6151
R1877 B.n591 B.n590 10.6151
R1878 B.n591 B.n403 10.6151
R1879 B.n601 B.n403 10.6151
R1880 B.n602 B.n601 10.6151
R1881 B.n603 B.n602 10.6151
R1882 B.n603 B.n395 10.6151
R1883 B.n613 B.n395 10.6151
R1884 B.n614 B.n613 10.6151
R1885 B.n615 B.n614 10.6151
R1886 B.n615 B.n387 10.6151
R1887 B.n625 B.n387 10.6151
R1888 B.n626 B.n625 10.6151
R1889 B.n627 B.n626 10.6151
R1890 B.n627 B.n379 10.6151
R1891 B.n637 B.n379 10.6151
R1892 B.n638 B.n637 10.6151
R1893 B.n639 B.n638 10.6151
R1894 B.n639 B.n371 10.6151
R1895 B.n649 B.n371 10.6151
R1896 B.n650 B.n649 10.6151
R1897 B.n651 B.n650 10.6151
R1898 B.n651 B.n363 10.6151
R1899 B.n661 B.n363 10.6151
R1900 B.n662 B.n661 10.6151
R1901 B.n663 B.n662 10.6151
R1902 B.n663 B.n355 10.6151
R1903 B.n674 B.n355 10.6151
R1904 B.n675 B.n674 10.6151
R1905 B.n676 B.n675 10.6151
R1906 B.n676 B.n348 10.6151
R1907 B.n686 B.n348 10.6151
R1908 B.n687 B.n686 10.6151
R1909 B.n688 B.n687 10.6151
R1910 B.n688 B.n340 10.6151
R1911 B.n698 B.n340 10.6151
R1912 B.n699 B.n698 10.6151
R1913 B.n700 B.n699 10.6151
R1914 B.n700 B.n332 10.6151
R1915 B.n710 B.n332 10.6151
R1916 B.n711 B.n710 10.6151
R1917 B.n712 B.n711 10.6151
R1918 B.n712 B.n324 10.6151
R1919 B.n722 B.n324 10.6151
R1920 B.n723 B.n722 10.6151
R1921 B.n724 B.n723 10.6151
R1922 B.n724 B.n316 10.6151
R1923 B.n734 B.n316 10.6151
R1924 B.n735 B.n734 10.6151
R1925 B.n736 B.n735 10.6151
R1926 B.n736 B.n308 10.6151
R1927 B.n746 B.n308 10.6151
R1928 B.n747 B.n746 10.6151
R1929 B.n748 B.n747 10.6151
R1930 B.n748 B.n300 10.6151
R1931 B.n758 B.n300 10.6151
R1932 B.n759 B.n758 10.6151
R1933 B.n760 B.n759 10.6151
R1934 B.n760 B.n292 10.6151
R1935 B.n771 B.n292 10.6151
R1936 B.n772 B.n771 10.6151
R1937 B.n773 B.n772 10.6151
R1938 B.n773 B.n285 10.6151
R1939 B.n784 B.n285 10.6151
R1940 B.n785 B.n784 10.6151
R1941 B.n786 B.n785 10.6151
R1942 B.n786 B.n0 10.6151
R1943 B.n1026 B.n1 10.6151
R1944 B.n1026 B.n1025 10.6151
R1945 B.n1025 B.n1024 10.6151
R1946 B.n1024 B.n10 10.6151
R1947 B.n1018 B.n10 10.6151
R1948 B.n1018 B.n1017 10.6151
R1949 B.n1017 B.n1016 10.6151
R1950 B.n1016 B.n16 10.6151
R1951 B.n1010 B.n16 10.6151
R1952 B.n1010 B.n1009 10.6151
R1953 B.n1009 B.n1008 10.6151
R1954 B.n1008 B.n24 10.6151
R1955 B.n1002 B.n24 10.6151
R1956 B.n1002 B.n1001 10.6151
R1957 B.n1001 B.n1000 10.6151
R1958 B.n1000 B.n31 10.6151
R1959 B.n994 B.n31 10.6151
R1960 B.n994 B.n993 10.6151
R1961 B.n993 B.n992 10.6151
R1962 B.n992 B.n38 10.6151
R1963 B.n986 B.n38 10.6151
R1964 B.n986 B.n985 10.6151
R1965 B.n985 B.n984 10.6151
R1966 B.n984 B.n45 10.6151
R1967 B.n978 B.n45 10.6151
R1968 B.n978 B.n977 10.6151
R1969 B.n977 B.n976 10.6151
R1970 B.n976 B.n52 10.6151
R1971 B.n970 B.n52 10.6151
R1972 B.n970 B.n969 10.6151
R1973 B.n969 B.n968 10.6151
R1974 B.n968 B.n59 10.6151
R1975 B.n962 B.n59 10.6151
R1976 B.n962 B.n961 10.6151
R1977 B.n961 B.n960 10.6151
R1978 B.n960 B.n66 10.6151
R1979 B.n954 B.n66 10.6151
R1980 B.n954 B.n953 10.6151
R1981 B.n953 B.n952 10.6151
R1982 B.n952 B.n72 10.6151
R1983 B.n946 B.n72 10.6151
R1984 B.n946 B.n945 10.6151
R1985 B.n945 B.n944 10.6151
R1986 B.n944 B.n80 10.6151
R1987 B.n938 B.n80 10.6151
R1988 B.n938 B.n937 10.6151
R1989 B.n937 B.n936 10.6151
R1990 B.n936 B.n87 10.6151
R1991 B.n930 B.n87 10.6151
R1992 B.n930 B.n929 10.6151
R1993 B.n929 B.n928 10.6151
R1994 B.n928 B.n94 10.6151
R1995 B.n922 B.n94 10.6151
R1996 B.n922 B.n921 10.6151
R1997 B.n921 B.n920 10.6151
R1998 B.n920 B.n101 10.6151
R1999 B.n914 B.n101 10.6151
R2000 B.n914 B.n913 10.6151
R2001 B.n913 B.n912 10.6151
R2002 B.n912 B.n108 10.6151
R2003 B.n906 B.n108 10.6151
R2004 B.n906 B.n905 10.6151
R2005 B.n905 B.n904 10.6151
R2006 B.n904 B.n115 10.6151
R2007 B.n898 B.n115 10.6151
R2008 B.n898 B.n897 10.6151
R2009 B.n897 B.n896 10.6151
R2010 B.n896 B.n122 10.6151
R2011 B.n890 B.n122 10.6151
R2012 B.n890 B.n889 10.6151
R2013 B.n889 B.n888 10.6151
R2014 B.n671 B.t8 8.56081
R2015 B.n74 B.t3 8.56081
R2016 B.n216 B.n215 6.5566
R2017 B.n232 B.n164 6.5566
R2018 B.n506 B.n443 6.5566
R2019 B.n523 B.n522 6.5566
R2020 B.n768 B.t7 4.75623
R2021 B.n18 B.t5 4.75623
R2022 B.n215 B.n214 4.05904
R2023 B.n235 B.n164 4.05904
R2024 B.n444 B.n443 4.05904
R2025 B.n524 B.n523 4.05904
R2026 B.n1032 B.n0 2.81026
R2027 B.n1032 B.n1 2.81026
R2028 VP.n32 VP.n31 161.3
R2029 VP.n33 VP.n28 161.3
R2030 VP.n35 VP.n34 161.3
R2031 VP.n36 VP.n27 161.3
R2032 VP.n38 VP.n37 161.3
R2033 VP.n39 VP.n26 161.3
R2034 VP.n41 VP.n40 161.3
R2035 VP.n42 VP.n25 161.3
R2036 VP.n44 VP.n43 161.3
R2037 VP.n45 VP.n24 161.3
R2038 VP.n47 VP.n46 161.3
R2039 VP.n48 VP.n23 161.3
R2040 VP.n50 VP.n49 161.3
R2041 VP.n51 VP.n22 161.3
R2042 VP.n53 VP.n52 161.3
R2043 VP.n55 VP.n54 161.3
R2044 VP.n56 VP.n20 161.3
R2045 VP.n58 VP.n57 161.3
R2046 VP.n59 VP.n19 161.3
R2047 VP.n61 VP.n60 161.3
R2048 VP.n62 VP.n18 161.3
R2049 VP.n64 VP.n63 161.3
R2050 VP.n111 VP.n110 161.3
R2051 VP.n109 VP.n1 161.3
R2052 VP.n108 VP.n107 161.3
R2053 VP.n106 VP.n2 161.3
R2054 VP.n105 VP.n104 161.3
R2055 VP.n103 VP.n3 161.3
R2056 VP.n102 VP.n101 161.3
R2057 VP.n100 VP.n99 161.3
R2058 VP.n98 VP.n5 161.3
R2059 VP.n97 VP.n96 161.3
R2060 VP.n95 VP.n6 161.3
R2061 VP.n94 VP.n93 161.3
R2062 VP.n92 VP.n7 161.3
R2063 VP.n91 VP.n90 161.3
R2064 VP.n89 VP.n8 161.3
R2065 VP.n88 VP.n87 161.3
R2066 VP.n86 VP.n9 161.3
R2067 VP.n85 VP.n84 161.3
R2068 VP.n83 VP.n10 161.3
R2069 VP.n82 VP.n81 161.3
R2070 VP.n80 VP.n11 161.3
R2071 VP.n79 VP.n78 161.3
R2072 VP.n77 VP.n76 161.3
R2073 VP.n75 VP.n13 161.3
R2074 VP.n74 VP.n73 161.3
R2075 VP.n72 VP.n14 161.3
R2076 VP.n71 VP.n70 161.3
R2077 VP.n69 VP.n15 161.3
R2078 VP.n68 VP.n67 161.3
R2079 VP.n30 VP.t7 78.5414
R2080 VP.n66 VP.n16 78.3232
R2081 VP.n112 VP.n0 78.3232
R2082 VP.n65 VP.n17 78.3232
R2083 VP.n30 VP.n29 68.6407
R2084 VP.n85 VP.n10 56.5193
R2085 VP.n93 VP.n6 56.5193
R2086 VP.n46 VP.n23 56.5193
R2087 VP.n38 VP.n27 56.5193
R2088 VP.n66 VP.n65 52.6054
R2089 VP.n74 VP.n14 47.2923
R2090 VP.n104 VP.n2 47.2923
R2091 VP.n57 VP.n19 47.2923
R2092 VP.n8 VP.t5 46.0762
R2093 VP.n16 VP.t2 46.0762
R2094 VP.n12 VP.t4 46.0762
R2095 VP.n4 VP.t3 46.0762
R2096 VP.n0 VP.t6 46.0762
R2097 VP.n25 VP.t9 46.0762
R2098 VP.n17 VP.t8 46.0762
R2099 VP.n21 VP.t0 46.0762
R2100 VP.n29 VP.t1 46.0762
R2101 VP.n70 VP.n14 33.6945
R2102 VP.n108 VP.n2 33.6945
R2103 VP.n61 VP.n19 33.6945
R2104 VP.n69 VP.n68 24.4675
R2105 VP.n70 VP.n69 24.4675
R2106 VP.n75 VP.n74 24.4675
R2107 VP.n76 VP.n75 24.4675
R2108 VP.n80 VP.n79 24.4675
R2109 VP.n81 VP.n80 24.4675
R2110 VP.n81 VP.n10 24.4675
R2111 VP.n86 VP.n85 24.4675
R2112 VP.n87 VP.n86 24.4675
R2113 VP.n87 VP.n8 24.4675
R2114 VP.n91 VP.n8 24.4675
R2115 VP.n92 VP.n91 24.4675
R2116 VP.n93 VP.n92 24.4675
R2117 VP.n97 VP.n6 24.4675
R2118 VP.n98 VP.n97 24.4675
R2119 VP.n99 VP.n98 24.4675
R2120 VP.n103 VP.n102 24.4675
R2121 VP.n104 VP.n103 24.4675
R2122 VP.n109 VP.n108 24.4675
R2123 VP.n110 VP.n109 24.4675
R2124 VP.n62 VP.n61 24.4675
R2125 VP.n63 VP.n62 24.4675
R2126 VP.n50 VP.n23 24.4675
R2127 VP.n51 VP.n50 24.4675
R2128 VP.n52 VP.n51 24.4675
R2129 VP.n56 VP.n55 24.4675
R2130 VP.n57 VP.n56 24.4675
R2131 VP.n39 VP.n38 24.4675
R2132 VP.n40 VP.n39 24.4675
R2133 VP.n40 VP.n25 24.4675
R2134 VP.n44 VP.n25 24.4675
R2135 VP.n45 VP.n44 24.4675
R2136 VP.n46 VP.n45 24.4675
R2137 VP.n33 VP.n32 24.4675
R2138 VP.n34 VP.n33 24.4675
R2139 VP.n34 VP.n27 24.4675
R2140 VP.n76 VP.n12 18.5954
R2141 VP.n102 VP.n4 18.5954
R2142 VP.n55 VP.n21 18.5954
R2143 VP.n68 VP.n16 11.7447
R2144 VP.n110 VP.n0 11.7447
R2145 VP.n63 VP.n17 11.7447
R2146 VP.n79 VP.n12 5.87258
R2147 VP.n99 VP.n4 5.87258
R2148 VP.n52 VP.n21 5.87258
R2149 VP.n32 VP.n29 5.87258
R2150 VP.n31 VP.n30 4.31089
R2151 VP.n65 VP.n64 0.354971
R2152 VP.n67 VP.n66 0.354971
R2153 VP.n112 VP.n111 0.354971
R2154 VP VP.n112 0.26696
R2155 VP.n31 VP.n28 0.189894
R2156 VP.n35 VP.n28 0.189894
R2157 VP.n36 VP.n35 0.189894
R2158 VP.n37 VP.n36 0.189894
R2159 VP.n37 VP.n26 0.189894
R2160 VP.n41 VP.n26 0.189894
R2161 VP.n42 VP.n41 0.189894
R2162 VP.n43 VP.n42 0.189894
R2163 VP.n43 VP.n24 0.189894
R2164 VP.n47 VP.n24 0.189894
R2165 VP.n48 VP.n47 0.189894
R2166 VP.n49 VP.n48 0.189894
R2167 VP.n49 VP.n22 0.189894
R2168 VP.n53 VP.n22 0.189894
R2169 VP.n54 VP.n53 0.189894
R2170 VP.n54 VP.n20 0.189894
R2171 VP.n58 VP.n20 0.189894
R2172 VP.n59 VP.n58 0.189894
R2173 VP.n60 VP.n59 0.189894
R2174 VP.n60 VP.n18 0.189894
R2175 VP.n64 VP.n18 0.189894
R2176 VP.n67 VP.n15 0.189894
R2177 VP.n71 VP.n15 0.189894
R2178 VP.n72 VP.n71 0.189894
R2179 VP.n73 VP.n72 0.189894
R2180 VP.n73 VP.n13 0.189894
R2181 VP.n77 VP.n13 0.189894
R2182 VP.n78 VP.n77 0.189894
R2183 VP.n78 VP.n11 0.189894
R2184 VP.n82 VP.n11 0.189894
R2185 VP.n83 VP.n82 0.189894
R2186 VP.n84 VP.n83 0.189894
R2187 VP.n84 VP.n9 0.189894
R2188 VP.n88 VP.n9 0.189894
R2189 VP.n89 VP.n88 0.189894
R2190 VP.n90 VP.n89 0.189894
R2191 VP.n90 VP.n7 0.189894
R2192 VP.n94 VP.n7 0.189894
R2193 VP.n95 VP.n94 0.189894
R2194 VP.n96 VP.n95 0.189894
R2195 VP.n96 VP.n5 0.189894
R2196 VP.n100 VP.n5 0.189894
R2197 VP.n101 VP.n100 0.189894
R2198 VP.n101 VP.n3 0.189894
R2199 VP.n105 VP.n3 0.189894
R2200 VP.n106 VP.n105 0.189894
R2201 VP.n107 VP.n106 0.189894
R2202 VP.n107 VP.n1 0.189894
R2203 VP.n111 VP.n1 0.189894
R2204 VDD1.n1 VDD1.t2 71.507
R2205 VDD1.n3 VDD1.t7 71.5069
R2206 VDD1.n5 VDD1.n4 67.5234
R2207 VDD1.n1 VDD1.n0 65.2385
R2208 VDD1.n7 VDD1.n6 65.2383
R2209 VDD1.n3 VDD1.n2 65.2383
R2210 VDD1.n7 VDD1.n5 46.1043
R2211 VDD1.n6 VDD1.t9 3.14835
R2212 VDD1.n6 VDD1.t1 3.14835
R2213 VDD1.n0 VDD1.t8 3.14835
R2214 VDD1.n0 VDD1.t0 3.14835
R2215 VDD1.n4 VDD1.t6 3.14835
R2216 VDD1.n4 VDD1.t3 3.14835
R2217 VDD1.n2 VDD1.t5 3.14835
R2218 VDD1.n2 VDD1.t4 3.14835
R2219 VDD1 VDD1.n7 2.28283
R2220 VDD1 VDD1.n1 0.838862
R2221 VDD1.n5 VDD1.n3 0.725326
C0 VTAIL VP 7.55393f
C1 VTAIL VDD2 8.375401f
C2 VDD1 VP 6.60462f
C3 VDD1 VDD2 2.62327f
C4 VP VDD2 0.671231f
C5 VTAIL VN 7.53975f
C6 VDD1 VN 0.154932f
C7 VP VN 8.36153f
C8 VDD2 VN 6.09141f
C9 VDD1 VTAIL 8.31816f
C10 VDD2 B 7.067836f
C11 VDD1 B 6.989308f
C12 VTAIL B 5.896627f
C13 VN B 20.796198f
C14 VP B 19.356356f
C15 VDD1.t2 B 1.45008f
C16 VDD1.t8 B 0.133922f
C17 VDD1.t0 B 0.133922f
C18 VDD1.n0 B 1.12252f
C19 VDD1.n1 B 1.10382f
C20 VDD1.t7 B 1.45007f
C21 VDD1.t5 B 0.133922f
C22 VDD1.t4 B 0.133922f
C23 VDD1.n2 B 1.12252f
C24 VDD1.n3 B 1.09483f
C25 VDD1.t6 B 0.133922f
C26 VDD1.t3 B 0.133922f
C27 VDD1.n4 B 1.14624f
C28 VDD1.n5 B 3.29008f
C29 VDD1.t9 B 0.133922f
C30 VDD1.t1 B 0.133922f
C31 VDD1.n6 B 1.12252f
C32 VDD1.n7 B 3.25502f
C33 VP.t6 B 1.17832f
C34 VP.n0 B 0.514837f
C35 VP.n1 B 0.021455f
C36 VP.n2 B 0.018733f
C37 VP.n3 B 0.021455f
C38 VP.t3 B 1.17832f
C39 VP.n4 B 0.434495f
C40 VP.n5 B 0.021455f
C41 VP.n6 B 0.027733f
C42 VP.n7 B 0.021455f
C43 VP.t5 B 1.17832f
C44 VP.n8 B 0.454739f
C45 VP.n9 B 0.021455f
C46 VP.n10 B 0.027733f
C47 VP.n11 B 0.021455f
C48 VP.t4 B 1.17832f
C49 VP.n12 B 0.434495f
C50 VP.n13 B 0.021455f
C51 VP.n14 B 0.018733f
C52 VP.n15 B 0.021455f
C53 VP.t2 B 1.17832f
C54 VP.n16 B 0.514837f
C55 VP.t8 B 1.17832f
C56 VP.n17 B 0.514837f
C57 VP.n18 B 0.021455f
C58 VP.n19 B 0.018733f
C59 VP.n20 B 0.021455f
C60 VP.t0 B 1.17832f
C61 VP.n21 B 0.434495f
C62 VP.n22 B 0.021455f
C63 VP.n23 B 0.027733f
C64 VP.n24 B 0.021455f
C65 VP.t9 B 1.17832f
C66 VP.n25 B 0.454739f
C67 VP.n26 B 0.021455f
C68 VP.n27 B 0.027733f
C69 VP.n28 B 0.021455f
C70 VP.t1 B 1.17832f
C71 VP.n29 B 0.501539f
C72 VP.t7 B 1.42027f
C73 VP.n30 B 0.480899f
C74 VP.n31 B 0.252891f
C75 VP.n32 B 0.024983f
C76 VP.n33 B 0.039986f
C77 VP.n34 B 0.039986f
C78 VP.n35 B 0.021455f
C79 VP.n36 B 0.021455f
C80 VP.n37 B 0.021455f
C81 VP.n38 B 0.034907f
C82 VP.n39 B 0.039986f
C83 VP.n40 B 0.039986f
C84 VP.n41 B 0.021455f
C85 VP.n42 B 0.021455f
C86 VP.n43 B 0.021455f
C87 VP.n44 B 0.039986f
C88 VP.n45 B 0.039986f
C89 VP.n46 B 0.034907f
C90 VP.n47 B 0.021455f
C91 VP.n48 B 0.021455f
C92 VP.n49 B 0.021455f
C93 VP.n50 B 0.039986f
C94 VP.n51 B 0.039986f
C95 VP.n52 B 0.024983f
C96 VP.n53 B 0.021455f
C97 VP.n54 B 0.021455f
C98 VP.n55 B 0.035248f
C99 VP.n56 B 0.039986f
C100 VP.n57 B 0.040556f
C101 VP.n58 B 0.021455f
C102 VP.n59 B 0.021455f
C103 VP.n60 B 0.021455f
C104 VP.n61 B 0.043337f
C105 VP.n62 B 0.039986f
C106 VP.n63 B 0.029721f
C107 VP.n64 B 0.034627f
C108 VP.n65 B 1.31329f
C109 VP.n66 B 1.32795f
C110 VP.n67 B 0.034627f
C111 VP.n68 B 0.029721f
C112 VP.n69 B 0.039986f
C113 VP.n70 B 0.043337f
C114 VP.n71 B 0.021455f
C115 VP.n72 B 0.021455f
C116 VP.n73 B 0.021455f
C117 VP.n74 B 0.040556f
C118 VP.n75 B 0.039986f
C119 VP.n76 B 0.035248f
C120 VP.n77 B 0.021455f
C121 VP.n78 B 0.021455f
C122 VP.n79 B 0.024983f
C123 VP.n80 B 0.039986f
C124 VP.n81 B 0.039986f
C125 VP.n82 B 0.021455f
C126 VP.n83 B 0.021455f
C127 VP.n84 B 0.021455f
C128 VP.n85 B 0.034907f
C129 VP.n86 B 0.039986f
C130 VP.n87 B 0.039986f
C131 VP.n88 B 0.021455f
C132 VP.n89 B 0.021455f
C133 VP.n90 B 0.021455f
C134 VP.n91 B 0.039986f
C135 VP.n92 B 0.039986f
C136 VP.n93 B 0.034907f
C137 VP.n94 B 0.021455f
C138 VP.n95 B 0.021455f
C139 VP.n96 B 0.021455f
C140 VP.n97 B 0.039986f
C141 VP.n98 B 0.039986f
C142 VP.n99 B 0.024983f
C143 VP.n100 B 0.021455f
C144 VP.n101 B 0.021455f
C145 VP.n102 B 0.035248f
C146 VP.n103 B 0.039986f
C147 VP.n104 B 0.040556f
C148 VP.n105 B 0.021455f
C149 VP.n106 B 0.021455f
C150 VP.n107 B 0.021455f
C151 VP.n108 B 0.043337f
C152 VP.n109 B 0.039986f
C153 VP.n110 B 0.029721f
C154 VP.n111 B 0.034627f
C155 VP.n112 B 0.054208f
C156 VTAIL.t9 B 0.145394f
C157 VTAIL.t13 B 0.145394f
C158 VTAIL.n0 B 1.13843f
C159 VTAIL.n1 B 0.697126f
C160 VTAIL.t7 B 1.45037f
C161 VTAIL.n2 B 0.849773f
C162 VTAIL.t2 B 0.145394f
C163 VTAIL.t4 B 0.145394f
C164 VTAIL.n3 B 1.13843f
C165 VTAIL.n4 B 0.867961f
C166 VTAIL.t1 B 0.145394f
C167 VTAIL.t8 B 0.145394f
C168 VTAIL.n5 B 1.13843f
C169 VTAIL.n6 B 2.07052f
C170 VTAIL.t11 B 0.145394f
C171 VTAIL.t18 B 0.145394f
C172 VTAIL.n7 B 1.13844f
C173 VTAIL.n8 B 2.07052f
C174 VTAIL.t10 B 0.145394f
C175 VTAIL.t12 B 0.145394f
C176 VTAIL.n9 B 1.13844f
C177 VTAIL.n10 B 0.867955f
C178 VTAIL.t15 B 1.45038f
C179 VTAIL.n11 B 0.849763f
C180 VTAIL.t5 B 0.145394f
C181 VTAIL.t6 B 0.145394f
C182 VTAIL.n12 B 1.13844f
C183 VTAIL.n13 B 0.765169f
C184 VTAIL.t0 B 0.145394f
C185 VTAIL.t3 B 0.145394f
C186 VTAIL.n14 B 1.13844f
C187 VTAIL.n15 B 0.867955f
C188 VTAIL.t19 B 1.45037f
C189 VTAIL.n16 B 1.86098f
C190 VTAIL.t17 B 1.45037f
C191 VTAIL.n17 B 1.86098f
C192 VTAIL.t16 B 0.145394f
C193 VTAIL.t14 B 0.145394f
C194 VTAIL.n18 B 1.13843f
C195 VTAIL.n19 B 0.641874f
C196 VDD2.t6 B 1.42503f
C197 VDD2.t4 B 0.131609f
C198 VDD2.t5 B 0.131609f
C199 VDD2.n0 B 1.10313f
C200 VDD2.n1 B 1.07593f
C201 VDD2.t7 B 0.131609f
C202 VDD2.t2 B 0.131609f
C203 VDD2.n2 B 1.12644f
C204 VDD2.n3 B 3.08618f
C205 VDD2.t9 B 1.40083f
C206 VDD2.n4 B 3.11461f
C207 VDD2.t1 B 0.131609f
C208 VDD2.t8 B 0.131609f
C209 VDD2.n5 B 1.10314f
C210 VDD2.n6 B 0.554292f
C211 VDD2.t0 B 0.131609f
C212 VDD2.t3 B 0.131609f
C213 VDD2.n7 B 1.12639f
C214 VN.t1 B 1.14551f
C215 VN.n0 B 0.500501f
C216 VN.n1 B 0.020857f
C217 VN.n2 B 0.018212f
C218 VN.n3 B 0.020857f
C219 VN.t4 B 1.14551f
C220 VN.n4 B 0.422396f
C221 VN.n5 B 0.020857f
C222 VN.n6 B 0.026961f
C223 VN.n7 B 0.020857f
C224 VN.t2 B 1.14551f
C225 VN.n8 B 0.442077f
C226 VN.n9 B 0.020857f
C227 VN.n10 B 0.026961f
C228 VN.n11 B 0.020857f
C229 VN.t5 B 1.14551f
C230 VN.n12 B 0.487573f
C231 VN.t9 B 1.38072f
C232 VN.n13 B 0.467508f
C233 VN.n14 B 0.245849f
C234 VN.n15 B 0.024287f
C235 VN.n16 B 0.038873f
C236 VN.n17 B 0.038873f
C237 VN.n18 B 0.020857f
C238 VN.n19 B 0.020857f
C239 VN.n20 B 0.020857f
C240 VN.n21 B 0.033935f
C241 VN.n22 B 0.038873f
C242 VN.n23 B 0.038873f
C243 VN.n24 B 0.020857f
C244 VN.n25 B 0.020857f
C245 VN.n26 B 0.020857f
C246 VN.n27 B 0.038873f
C247 VN.n28 B 0.038873f
C248 VN.n29 B 0.033935f
C249 VN.n30 B 0.020857f
C250 VN.n31 B 0.020857f
C251 VN.n32 B 0.020857f
C252 VN.n33 B 0.038873f
C253 VN.n34 B 0.038873f
C254 VN.n35 B 0.024287f
C255 VN.n36 B 0.020857f
C256 VN.n37 B 0.020857f
C257 VN.n38 B 0.034267f
C258 VN.n39 B 0.038873f
C259 VN.n40 B 0.039427f
C260 VN.n41 B 0.020857f
C261 VN.n42 B 0.020857f
C262 VN.n43 B 0.020857f
C263 VN.n44 B 0.04213f
C264 VN.n45 B 0.038873f
C265 VN.n46 B 0.028893f
C266 VN.n47 B 0.033663f
C267 VN.n48 B 0.052698f
C268 VN.t7 B 1.14551f
C269 VN.n49 B 0.500501f
C270 VN.n50 B 0.020857f
C271 VN.n51 B 0.018212f
C272 VN.n52 B 0.020857f
C273 VN.t0 B 1.14551f
C274 VN.n53 B 0.422396f
C275 VN.n54 B 0.020857f
C276 VN.n55 B 0.026961f
C277 VN.n56 B 0.020857f
C278 VN.t8 B 1.14551f
C279 VN.n57 B 0.442077f
C280 VN.n58 B 0.020857f
C281 VN.n59 B 0.026961f
C282 VN.n60 B 0.020857f
C283 VN.t6 B 1.14551f
C284 VN.n61 B 0.487573f
C285 VN.t3 B 1.38072f
C286 VN.n62 B 0.467508f
C287 VN.n63 B 0.245849f
C288 VN.n64 B 0.024287f
C289 VN.n65 B 0.038873f
C290 VN.n66 B 0.038873f
C291 VN.n67 B 0.020857f
C292 VN.n68 B 0.020857f
C293 VN.n69 B 0.020857f
C294 VN.n70 B 0.033935f
C295 VN.n71 B 0.038873f
C296 VN.n72 B 0.038873f
C297 VN.n73 B 0.020857f
C298 VN.n74 B 0.020857f
C299 VN.n75 B 0.020857f
C300 VN.n76 B 0.038873f
C301 VN.n77 B 0.038873f
C302 VN.n78 B 0.033935f
C303 VN.n79 B 0.020857f
C304 VN.n80 B 0.020857f
C305 VN.n81 B 0.020857f
C306 VN.n82 B 0.038873f
C307 VN.n83 B 0.038873f
C308 VN.n84 B 0.024287f
C309 VN.n85 B 0.020857f
C310 VN.n86 B 0.020857f
C311 VN.n87 B 0.034267f
C312 VN.n88 B 0.038873f
C313 VN.n89 B 0.039427f
C314 VN.n90 B 0.020857f
C315 VN.n91 B 0.020857f
C316 VN.n92 B 0.020857f
C317 VN.n93 B 0.04213f
C318 VN.n94 B 0.038873f
C319 VN.n95 B 0.028893f
C320 VN.n96 B 0.033663f
C321 VN.n97 B 1.28511f
.ends

