* NGSPICE file created from diff_pair_sample_0674.ext - technology: sky130A

.subckt diff_pair_sample_0674 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=6.1737 pd=32.44 as=0 ps=0 w=15.83 l=1.84
X1 VDD1.t3 VP.t0 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.61195 pd=16.16 as=6.1737 ps=32.44 w=15.83 l=1.84
X2 VTAIL.t0 VN.t0 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=6.1737 pd=32.44 as=2.61195 ps=16.16 w=15.83 l=1.84
X3 VDD1.t2 VP.t1 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.61195 pd=16.16 as=6.1737 ps=32.44 w=15.83 l=1.84
X4 VTAIL.t1 VN.t1 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=6.1737 pd=32.44 as=2.61195 ps=16.16 w=15.83 l=1.84
X5 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=6.1737 pd=32.44 as=0 ps=0 w=15.83 l=1.84
X6 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=6.1737 pd=32.44 as=0 ps=0 w=15.83 l=1.84
X7 VDD2.t1 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.61195 pd=16.16 as=6.1737 ps=32.44 w=15.83 l=1.84
X8 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.1737 pd=32.44 as=0 ps=0 w=15.83 l=1.84
X9 VTAIL.t4 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=6.1737 pd=32.44 as=2.61195 ps=16.16 w=15.83 l=1.84
X10 VTAIL.t7 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=6.1737 pd=32.44 as=2.61195 ps=16.16 w=15.83 l=1.84
X11 VDD2.t0 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.61195 pd=16.16 as=6.1737 ps=32.44 w=15.83 l=1.84
R0 B.n802 B.n801 585
R1 B.n803 B.n802 585
R2 B.n340 B.n110 585
R3 B.n339 B.n338 585
R4 B.n337 B.n336 585
R5 B.n335 B.n334 585
R6 B.n333 B.n332 585
R7 B.n331 B.n330 585
R8 B.n329 B.n328 585
R9 B.n327 B.n326 585
R10 B.n325 B.n324 585
R11 B.n323 B.n322 585
R12 B.n321 B.n320 585
R13 B.n319 B.n318 585
R14 B.n317 B.n316 585
R15 B.n315 B.n314 585
R16 B.n313 B.n312 585
R17 B.n311 B.n310 585
R18 B.n309 B.n308 585
R19 B.n307 B.n306 585
R20 B.n305 B.n304 585
R21 B.n303 B.n302 585
R22 B.n301 B.n300 585
R23 B.n299 B.n298 585
R24 B.n297 B.n296 585
R25 B.n295 B.n294 585
R26 B.n293 B.n292 585
R27 B.n291 B.n290 585
R28 B.n289 B.n288 585
R29 B.n287 B.n286 585
R30 B.n285 B.n284 585
R31 B.n283 B.n282 585
R32 B.n281 B.n280 585
R33 B.n279 B.n278 585
R34 B.n277 B.n276 585
R35 B.n275 B.n274 585
R36 B.n273 B.n272 585
R37 B.n271 B.n270 585
R38 B.n269 B.n268 585
R39 B.n267 B.n266 585
R40 B.n265 B.n264 585
R41 B.n263 B.n262 585
R42 B.n261 B.n260 585
R43 B.n259 B.n258 585
R44 B.n257 B.n256 585
R45 B.n255 B.n254 585
R46 B.n253 B.n252 585
R47 B.n251 B.n250 585
R48 B.n249 B.n248 585
R49 B.n247 B.n246 585
R50 B.n245 B.n244 585
R51 B.n243 B.n242 585
R52 B.n241 B.n240 585
R53 B.n239 B.n238 585
R54 B.n237 B.n236 585
R55 B.n235 B.n234 585
R56 B.n233 B.n232 585
R57 B.n231 B.n230 585
R58 B.n229 B.n228 585
R59 B.n227 B.n226 585
R60 B.n225 B.n224 585
R61 B.n223 B.n222 585
R62 B.n221 B.n220 585
R63 B.n218 B.n217 585
R64 B.n216 B.n215 585
R65 B.n214 B.n213 585
R66 B.n212 B.n211 585
R67 B.n210 B.n209 585
R68 B.n208 B.n207 585
R69 B.n206 B.n205 585
R70 B.n204 B.n203 585
R71 B.n202 B.n201 585
R72 B.n200 B.n199 585
R73 B.n198 B.n197 585
R74 B.n196 B.n195 585
R75 B.n194 B.n193 585
R76 B.n192 B.n191 585
R77 B.n190 B.n189 585
R78 B.n188 B.n187 585
R79 B.n186 B.n185 585
R80 B.n184 B.n183 585
R81 B.n182 B.n181 585
R82 B.n180 B.n179 585
R83 B.n178 B.n177 585
R84 B.n176 B.n175 585
R85 B.n174 B.n173 585
R86 B.n172 B.n171 585
R87 B.n170 B.n169 585
R88 B.n168 B.n167 585
R89 B.n166 B.n165 585
R90 B.n164 B.n163 585
R91 B.n162 B.n161 585
R92 B.n160 B.n159 585
R93 B.n158 B.n157 585
R94 B.n156 B.n155 585
R95 B.n154 B.n153 585
R96 B.n152 B.n151 585
R97 B.n150 B.n149 585
R98 B.n148 B.n147 585
R99 B.n146 B.n145 585
R100 B.n144 B.n143 585
R101 B.n142 B.n141 585
R102 B.n140 B.n139 585
R103 B.n138 B.n137 585
R104 B.n136 B.n135 585
R105 B.n134 B.n133 585
R106 B.n132 B.n131 585
R107 B.n130 B.n129 585
R108 B.n128 B.n127 585
R109 B.n126 B.n125 585
R110 B.n124 B.n123 585
R111 B.n122 B.n121 585
R112 B.n120 B.n119 585
R113 B.n118 B.n117 585
R114 B.n53 B.n52 585
R115 B.n806 B.n805 585
R116 B.n800 B.n111 585
R117 B.n111 B.n50 585
R118 B.n799 B.n49 585
R119 B.n810 B.n49 585
R120 B.n798 B.n48 585
R121 B.n811 B.n48 585
R122 B.n797 B.n47 585
R123 B.n812 B.n47 585
R124 B.n796 B.n795 585
R125 B.n795 B.n43 585
R126 B.n794 B.n42 585
R127 B.n818 B.n42 585
R128 B.n793 B.n41 585
R129 B.n819 B.n41 585
R130 B.n792 B.n40 585
R131 B.n820 B.n40 585
R132 B.n791 B.n790 585
R133 B.n790 B.n36 585
R134 B.n789 B.n35 585
R135 B.n826 B.n35 585
R136 B.n788 B.n34 585
R137 B.n827 B.n34 585
R138 B.n787 B.n33 585
R139 B.n828 B.n33 585
R140 B.n786 B.n785 585
R141 B.n785 B.n29 585
R142 B.n784 B.n28 585
R143 B.n834 B.n28 585
R144 B.n783 B.n27 585
R145 B.n835 B.n27 585
R146 B.n782 B.n26 585
R147 B.n836 B.n26 585
R148 B.n781 B.n780 585
R149 B.n780 B.n22 585
R150 B.n779 B.n21 585
R151 B.n842 B.n21 585
R152 B.n778 B.n20 585
R153 B.n843 B.n20 585
R154 B.n777 B.n19 585
R155 B.n844 B.n19 585
R156 B.n776 B.n775 585
R157 B.n775 B.n15 585
R158 B.n774 B.n14 585
R159 B.n850 B.n14 585
R160 B.n773 B.n13 585
R161 B.n851 B.n13 585
R162 B.n772 B.n12 585
R163 B.n852 B.n12 585
R164 B.n771 B.n770 585
R165 B.n770 B.n8 585
R166 B.n769 B.n7 585
R167 B.n858 B.n7 585
R168 B.n768 B.n6 585
R169 B.n859 B.n6 585
R170 B.n767 B.n5 585
R171 B.n860 B.n5 585
R172 B.n766 B.n765 585
R173 B.n765 B.n4 585
R174 B.n764 B.n341 585
R175 B.n764 B.n763 585
R176 B.n754 B.n342 585
R177 B.n343 B.n342 585
R178 B.n756 B.n755 585
R179 B.n757 B.n756 585
R180 B.n753 B.n347 585
R181 B.n351 B.n347 585
R182 B.n752 B.n751 585
R183 B.n751 B.n750 585
R184 B.n349 B.n348 585
R185 B.n350 B.n349 585
R186 B.n743 B.n742 585
R187 B.n744 B.n743 585
R188 B.n741 B.n356 585
R189 B.n356 B.n355 585
R190 B.n740 B.n739 585
R191 B.n739 B.n738 585
R192 B.n358 B.n357 585
R193 B.n359 B.n358 585
R194 B.n731 B.n730 585
R195 B.n732 B.n731 585
R196 B.n729 B.n364 585
R197 B.n364 B.n363 585
R198 B.n728 B.n727 585
R199 B.n727 B.n726 585
R200 B.n366 B.n365 585
R201 B.n367 B.n366 585
R202 B.n719 B.n718 585
R203 B.n720 B.n719 585
R204 B.n717 B.n372 585
R205 B.n372 B.n371 585
R206 B.n716 B.n715 585
R207 B.n715 B.n714 585
R208 B.n374 B.n373 585
R209 B.n375 B.n374 585
R210 B.n707 B.n706 585
R211 B.n708 B.n707 585
R212 B.n705 B.n379 585
R213 B.n383 B.n379 585
R214 B.n704 B.n703 585
R215 B.n703 B.n702 585
R216 B.n381 B.n380 585
R217 B.n382 B.n381 585
R218 B.n695 B.n694 585
R219 B.n696 B.n695 585
R220 B.n693 B.n388 585
R221 B.n388 B.n387 585
R222 B.n692 B.n691 585
R223 B.n691 B.n690 585
R224 B.n390 B.n389 585
R225 B.n391 B.n390 585
R226 B.n686 B.n685 585
R227 B.n394 B.n393 585
R228 B.n682 B.n681 585
R229 B.n683 B.n682 585
R230 B.n680 B.n451 585
R231 B.n679 B.n678 585
R232 B.n677 B.n676 585
R233 B.n675 B.n674 585
R234 B.n673 B.n672 585
R235 B.n671 B.n670 585
R236 B.n669 B.n668 585
R237 B.n667 B.n666 585
R238 B.n665 B.n664 585
R239 B.n663 B.n662 585
R240 B.n661 B.n660 585
R241 B.n659 B.n658 585
R242 B.n657 B.n656 585
R243 B.n655 B.n654 585
R244 B.n653 B.n652 585
R245 B.n651 B.n650 585
R246 B.n649 B.n648 585
R247 B.n647 B.n646 585
R248 B.n645 B.n644 585
R249 B.n643 B.n642 585
R250 B.n641 B.n640 585
R251 B.n639 B.n638 585
R252 B.n637 B.n636 585
R253 B.n635 B.n634 585
R254 B.n633 B.n632 585
R255 B.n631 B.n630 585
R256 B.n629 B.n628 585
R257 B.n627 B.n626 585
R258 B.n625 B.n624 585
R259 B.n623 B.n622 585
R260 B.n621 B.n620 585
R261 B.n619 B.n618 585
R262 B.n617 B.n616 585
R263 B.n615 B.n614 585
R264 B.n613 B.n612 585
R265 B.n611 B.n610 585
R266 B.n609 B.n608 585
R267 B.n607 B.n606 585
R268 B.n605 B.n604 585
R269 B.n603 B.n602 585
R270 B.n601 B.n600 585
R271 B.n599 B.n598 585
R272 B.n597 B.n596 585
R273 B.n595 B.n594 585
R274 B.n593 B.n592 585
R275 B.n591 B.n590 585
R276 B.n589 B.n588 585
R277 B.n587 B.n586 585
R278 B.n585 B.n584 585
R279 B.n583 B.n582 585
R280 B.n581 B.n580 585
R281 B.n579 B.n578 585
R282 B.n577 B.n576 585
R283 B.n575 B.n574 585
R284 B.n573 B.n572 585
R285 B.n571 B.n570 585
R286 B.n569 B.n568 585
R287 B.n567 B.n566 585
R288 B.n565 B.n564 585
R289 B.n562 B.n561 585
R290 B.n560 B.n559 585
R291 B.n558 B.n557 585
R292 B.n556 B.n555 585
R293 B.n554 B.n553 585
R294 B.n552 B.n551 585
R295 B.n550 B.n549 585
R296 B.n548 B.n547 585
R297 B.n546 B.n545 585
R298 B.n544 B.n543 585
R299 B.n542 B.n541 585
R300 B.n540 B.n539 585
R301 B.n538 B.n537 585
R302 B.n536 B.n535 585
R303 B.n534 B.n533 585
R304 B.n532 B.n531 585
R305 B.n530 B.n529 585
R306 B.n528 B.n527 585
R307 B.n526 B.n525 585
R308 B.n524 B.n523 585
R309 B.n522 B.n521 585
R310 B.n520 B.n519 585
R311 B.n518 B.n517 585
R312 B.n516 B.n515 585
R313 B.n514 B.n513 585
R314 B.n512 B.n511 585
R315 B.n510 B.n509 585
R316 B.n508 B.n507 585
R317 B.n506 B.n505 585
R318 B.n504 B.n503 585
R319 B.n502 B.n501 585
R320 B.n500 B.n499 585
R321 B.n498 B.n497 585
R322 B.n496 B.n495 585
R323 B.n494 B.n493 585
R324 B.n492 B.n491 585
R325 B.n490 B.n489 585
R326 B.n488 B.n487 585
R327 B.n486 B.n485 585
R328 B.n484 B.n483 585
R329 B.n482 B.n481 585
R330 B.n480 B.n479 585
R331 B.n478 B.n477 585
R332 B.n476 B.n475 585
R333 B.n474 B.n473 585
R334 B.n472 B.n471 585
R335 B.n470 B.n469 585
R336 B.n468 B.n467 585
R337 B.n466 B.n465 585
R338 B.n464 B.n463 585
R339 B.n462 B.n461 585
R340 B.n460 B.n459 585
R341 B.n458 B.n457 585
R342 B.n687 B.n392 585
R343 B.n392 B.n391 585
R344 B.n689 B.n688 585
R345 B.n690 B.n689 585
R346 B.n386 B.n385 585
R347 B.n387 B.n386 585
R348 B.n698 B.n697 585
R349 B.n697 B.n696 585
R350 B.n699 B.n384 585
R351 B.n384 B.n382 585
R352 B.n701 B.n700 585
R353 B.n702 B.n701 585
R354 B.n378 B.n377 585
R355 B.n383 B.n378 585
R356 B.n710 B.n709 585
R357 B.n709 B.n708 585
R358 B.n711 B.n376 585
R359 B.n376 B.n375 585
R360 B.n713 B.n712 585
R361 B.n714 B.n713 585
R362 B.n370 B.n369 585
R363 B.n371 B.n370 585
R364 B.n722 B.n721 585
R365 B.n721 B.n720 585
R366 B.n723 B.n368 585
R367 B.n368 B.n367 585
R368 B.n725 B.n724 585
R369 B.n726 B.n725 585
R370 B.n362 B.n361 585
R371 B.n363 B.n362 585
R372 B.n734 B.n733 585
R373 B.n733 B.n732 585
R374 B.n735 B.n360 585
R375 B.n360 B.n359 585
R376 B.n737 B.n736 585
R377 B.n738 B.n737 585
R378 B.n354 B.n353 585
R379 B.n355 B.n354 585
R380 B.n746 B.n745 585
R381 B.n745 B.n744 585
R382 B.n747 B.n352 585
R383 B.n352 B.n350 585
R384 B.n749 B.n748 585
R385 B.n750 B.n749 585
R386 B.n346 B.n345 585
R387 B.n351 B.n346 585
R388 B.n759 B.n758 585
R389 B.n758 B.n757 585
R390 B.n760 B.n344 585
R391 B.n344 B.n343 585
R392 B.n762 B.n761 585
R393 B.n763 B.n762 585
R394 B.n2 B.n0 585
R395 B.n4 B.n2 585
R396 B.n3 B.n1 585
R397 B.n859 B.n3 585
R398 B.n857 B.n856 585
R399 B.n858 B.n857 585
R400 B.n855 B.n9 585
R401 B.n9 B.n8 585
R402 B.n854 B.n853 585
R403 B.n853 B.n852 585
R404 B.n11 B.n10 585
R405 B.n851 B.n11 585
R406 B.n849 B.n848 585
R407 B.n850 B.n849 585
R408 B.n847 B.n16 585
R409 B.n16 B.n15 585
R410 B.n846 B.n845 585
R411 B.n845 B.n844 585
R412 B.n18 B.n17 585
R413 B.n843 B.n18 585
R414 B.n841 B.n840 585
R415 B.n842 B.n841 585
R416 B.n839 B.n23 585
R417 B.n23 B.n22 585
R418 B.n838 B.n837 585
R419 B.n837 B.n836 585
R420 B.n25 B.n24 585
R421 B.n835 B.n25 585
R422 B.n833 B.n832 585
R423 B.n834 B.n833 585
R424 B.n831 B.n30 585
R425 B.n30 B.n29 585
R426 B.n830 B.n829 585
R427 B.n829 B.n828 585
R428 B.n32 B.n31 585
R429 B.n827 B.n32 585
R430 B.n825 B.n824 585
R431 B.n826 B.n825 585
R432 B.n823 B.n37 585
R433 B.n37 B.n36 585
R434 B.n822 B.n821 585
R435 B.n821 B.n820 585
R436 B.n39 B.n38 585
R437 B.n819 B.n39 585
R438 B.n817 B.n816 585
R439 B.n818 B.n817 585
R440 B.n815 B.n44 585
R441 B.n44 B.n43 585
R442 B.n814 B.n813 585
R443 B.n813 B.n812 585
R444 B.n46 B.n45 585
R445 B.n811 B.n46 585
R446 B.n809 B.n808 585
R447 B.n810 B.n809 585
R448 B.n807 B.n51 585
R449 B.n51 B.n50 585
R450 B.n862 B.n861 585
R451 B.n861 B.n860 585
R452 B.n685 B.n392 569.379
R453 B.n805 B.n51 569.379
R454 B.n457 B.n390 569.379
R455 B.n802 B.n111 569.379
R456 B.n455 B.t11 413.854
R457 B.n452 B.t15 413.854
R458 B.n115 B.t4 413.854
R459 B.n112 B.t8 413.854
R460 B.n803 B.n109 256.663
R461 B.n803 B.n108 256.663
R462 B.n803 B.n107 256.663
R463 B.n803 B.n106 256.663
R464 B.n803 B.n105 256.663
R465 B.n803 B.n104 256.663
R466 B.n803 B.n103 256.663
R467 B.n803 B.n102 256.663
R468 B.n803 B.n101 256.663
R469 B.n803 B.n100 256.663
R470 B.n803 B.n99 256.663
R471 B.n803 B.n98 256.663
R472 B.n803 B.n97 256.663
R473 B.n803 B.n96 256.663
R474 B.n803 B.n95 256.663
R475 B.n803 B.n94 256.663
R476 B.n803 B.n93 256.663
R477 B.n803 B.n92 256.663
R478 B.n803 B.n91 256.663
R479 B.n803 B.n90 256.663
R480 B.n803 B.n89 256.663
R481 B.n803 B.n88 256.663
R482 B.n803 B.n87 256.663
R483 B.n803 B.n86 256.663
R484 B.n803 B.n85 256.663
R485 B.n803 B.n84 256.663
R486 B.n803 B.n83 256.663
R487 B.n803 B.n82 256.663
R488 B.n803 B.n81 256.663
R489 B.n803 B.n80 256.663
R490 B.n803 B.n79 256.663
R491 B.n803 B.n78 256.663
R492 B.n803 B.n77 256.663
R493 B.n803 B.n76 256.663
R494 B.n803 B.n75 256.663
R495 B.n803 B.n74 256.663
R496 B.n803 B.n73 256.663
R497 B.n803 B.n72 256.663
R498 B.n803 B.n71 256.663
R499 B.n803 B.n70 256.663
R500 B.n803 B.n69 256.663
R501 B.n803 B.n68 256.663
R502 B.n803 B.n67 256.663
R503 B.n803 B.n66 256.663
R504 B.n803 B.n65 256.663
R505 B.n803 B.n64 256.663
R506 B.n803 B.n63 256.663
R507 B.n803 B.n62 256.663
R508 B.n803 B.n61 256.663
R509 B.n803 B.n60 256.663
R510 B.n803 B.n59 256.663
R511 B.n803 B.n58 256.663
R512 B.n803 B.n57 256.663
R513 B.n803 B.n56 256.663
R514 B.n803 B.n55 256.663
R515 B.n803 B.n54 256.663
R516 B.n804 B.n803 256.663
R517 B.n684 B.n683 256.663
R518 B.n683 B.n395 256.663
R519 B.n683 B.n396 256.663
R520 B.n683 B.n397 256.663
R521 B.n683 B.n398 256.663
R522 B.n683 B.n399 256.663
R523 B.n683 B.n400 256.663
R524 B.n683 B.n401 256.663
R525 B.n683 B.n402 256.663
R526 B.n683 B.n403 256.663
R527 B.n683 B.n404 256.663
R528 B.n683 B.n405 256.663
R529 B.n683 B.n406 256.663
R530 B.n683 B.n407 256.663
R531 B.n683 B.n408 256.663
R532 B.n683 B.n409 256.663
R533 B.n683 B.n410 256.663
R534 B.n683 B.n411 256.663
R535 B.n683 B.n412 256.663
R536 B.n683 B.n413 256.663
R537 B.n683 B.n414 256.663
R538 B.n683 B.n415 256.663
R539 B.n683 B.n416 256.663
R540 B.n683 B.n417 256.663
R541 B.n683 B.n418 256.663
R542 B.n683 B.n419 256.663
R543 B.n683 B.n420 256.663
R544 B.n683 B.n421 256.663
R545 B.n683 B.n422 256.663
R546 B.n683 B.n423 256.663
R547 B.n683 B.n424 256.663
R548 B.n683 B.n425 256.663
R549 B.n683 B.n426 256.663
R550 B.n683 B.n427 256.663
R551 B.n683 B.n428 256.663
R552 B.n683 B.n429 256.663
R553 B.n683 B.n430 256.663
R554 B.n683 B.n431 256.663
R555 B.n683 B.n432 256.663
R556 B.n683 B.n433 256.663
R557 B.n683 B.n434 256.663
R558 B.n683 B.n435 256.663
R559 B.n683 B.n436 256.663
R560 B.n683 B.n437 256.663
R561 B.n683 B.n438 256.663
R562 B.n683 B.n439 256.663
R563 B.n683 B.n440 256.663
R564 B.n683 B.n441 256.663
R565 B.n683 B.n442 256.663
R566 B.n683 B.n443 256.663
R567 B.n683 B.n444 256.663
R568 B.n683 B.n445 256.663
R569 B.n683 B.n446 256.663
R570 B.n683 B.n447 256.663
R571 B.n683 B.n448 256.663
R572 B.n683 B.n449 256.663
R573 B.n683 B.n450 256.663
R574 B.n689 B.n392 163.367
R575 B.n689 B.n386 163.367
R576 B.n697 B.n386 163.367
R577 B.n697 B.n384 163.367
R578 B.n701 B.n384 163.367
R579 B.n701 B.n378 163.367
R580 B.n709 B.n378 163.367
R581 B.n709 B.n376 163.367
R582 B.n713 B.n376 163.367
R583 B.n713 B.n370 163.367
R584 B.n721 B.n370 163.367
R585 B.n721 B.n368 163.367
R586 B.n725 B.n368 163.367
R587 B.n725 B.n362 163.367
R588 B.n733 B.n362 163.367
R589 B.n733 B.n360 163.367
R590 B.n737 B.n360 163.367
R591 B.n737 B.n354 163.367
R592 B.n745 B.n354 163.367
R593 B.n745 B.n352 163.367
R594 B.n749 B.n352 163.367
R595 B.n749 B.n346 163.367
R596 B.n758 B.n346 163.367
R597 B.n758 B.n344 163.367
R598 B.n762 B.n344 163.367
R599 B.n762 B.n2 163.367
R600 B.n861 B.n2 163.367
R601 B.n861 B.n3 163.367
R602 B.n857 B.n3 163.367
R603 B.n857 B.n9 163.367
R604 B.n853 B.n9 163.367
R605 B.n853 B.n11 163.367
R606 B.n849 B.n11 163.367
R607 B.n849 B.n16 163.367
R608 B.n845 B.n16 163.367
R609 B.n845 B.n18 163.367
R610 B.n841 B.n18 163.367
R611 B.n841 B.n23 163.367
R612 B.n837 B.n23 163.367
R613 B.n837 B.n25 163.367
R614 B.n833 B.n25 163.367
R615 B.n833 B.n30 163.367
R616 B.n829 B.n30 163.367
R617 B.n829 B.n32 163.367
R618 B.n825 B.n32 163.367
R619 B.n825 B.n37 163.367
R620 B.n821 B.n37 163.367
R621 B.n821 B.n39 163.367
R622 B.n817 B.n39 163.367
R623 B.n817 B.n44 163.367
R624 B.n813 B.n44 163.367
R625 B.n813 B.n46 163.367
R626 B.n809 B.n46 163.367
R627 B.n809 B.n51 163.367
R628 B.n682 B.n394 163.367
R629 B.n682 B.n451 163.367
R630 B.n678 B.n677 163.367
R631 B.n674 B.n673 163.367
R632 B.n670 B.n669 163.367
R633 B.n666 B.n665 163.367
R634 B.n662 B.n661 163.367
R635 B.n658 B.n657 163.367
R636 B.n654 B.n653 163.367
R637 B.n650 B.n649 163.367
R638 B.n646 B.n645 163.367
R639 B.n642 B.n641 163.367
R640 B.n638 B.n637 163.367
R641 B.n634 B.n633 163.367
R642 B.n630 B.n629 163.367
R643 B.n626 B.n625 163.367
R644 B.n622 B.n621 163.367
R645 B.n618 B.n617 163.367
R646 B.n614 B.n613 163.367
R647 B.n610 B.n609 163.367
R648 B.n606 B.n605 163.367
R649 B.n602 B.n601 163.367
R650 B.n598 B.n597 163.367
R651 B.n594 B.n593 163.367
R652 B.n590 B.n589 163.367
R653 B.n586 B.n585 163.367
R654 B.n582 B.n581 163.367
R655 B.n578 B.n577 163.367
R656 B.n574 B.n573 163.367
R657 B.n570 B.n569 163.367
R658 B.n566 B.n565 163.367
R659 B.n561 B.n560 163.367
R660 B.n557 B.n556 163.367
R661 B.n553 B.n552 163.367
R662 B.n549 B.n548 163.367
R663 B.n545 B.n544 163.367
R664 B.n541 B.n540 163.367
R665 B.n537 B.n536 163.367
R666 B.n533 B.n532 163.367
R667 B.n529 B.n528 163.367
R668 B.n525 B.n524 163.367
R669 B.n521 B.n520 163.367
R670 B.n517 B.n516 163.367
R671 B.n513 B.n512 163.367
R672 B.n509 B.n508 163.367
R673 B.n505 B.n504 163.367
R674 B.n501 B.n500 163.367
R675 B.n497 B.n496 163.367
R676 B.n493 B.n492 163.367
R677 B.n489 B.n488 163.367
R678 B.n485 B.n484 163.367
R679 B.n481 B.n480 163.367
R680 B.n477 B.n476 163.367
R681 B.n473 B.n472 163.367
R682 B.n469 B.n468 163.367
R683 B.n465 B.n464 163.367
R684 B.n461 B.n460 163.367
R685 B.n691 B.n390 163.367
R686 B.n691 B.n388 163.367
R687 B.n695 B.n388 163.367
R688 B.n695 B.n381 163.367
R689 B.n703 B.n381 163.367
R690 B.n703 B.n379 163.367
R691 B.n707 B.n379 163.367
R692 B.n707 B.n374 163.367
R693 B.n715 B.n374 163.367
R694 B.n715 B.n372 163.367
R695 B.n719 B.n372 163.367
R696 B.n719 B.n366 163.367
R697 B.n727 B.n366 163.367
R698 B.n727 B.n364 163.367
R699 B.n731 B.n364 163.367
R700 B.n731 B.n358 163.367
R701 B.n739 B.n358 163.367
R702 B.n739 B.n356 163.367
R703 B.n743 B.n356 163.367
R704 B.n743 B.n349 163.367
R705 B.n751 B.n349 163.367
R706 B.n751 B.n347 163.367
R707 B.n756 B.n347 163.367
R708 B.n756 B.n342 163.367
R709 B.n764 B.n342 163.367
R710 B.n765 B.n764 163.367
R711 B.n765 B.n5 163.367
R712 B.n6 B.n5 163.367
R713 B.n7 B.n6 163.367
R714 B.n770 B.n7 163.367
R715 B.n770 B.n12 163.367
R716 B.n13 B.n12 163.367
R717 B.n14 B.n13 163.367
R718 B.n775 B.n14 163.367
R719 B.n775 B.n19 163.367
R720 B.n20 B.n19 163.367
R721 B.n21 B.n20 163.367
R722 B.n780 B.n21 163.367
R723 B.n780 B.n26 163.367
R724 B.n27 B.n26 163.367
R725 B.n28 B.n27 163.367
R726 B.n785 B.n28 163.367
R727 B.n785 B.n33 163.367
R728 B.n34 B.n33 163.367
R729 B.n35 B.n34 163.367
R730 B.n790 B.n35 163.367
R731 B.n790 B.n40 163.367
R732 B.n41 B.n40 163.367
R733 B.n42 B.n41 163.367
R734 B.n795 B.n42 163.367
R735 B.n795 B.n47 163.367
R736 B.n48 B.n47 163.367
R737 B.n49 B.n48 163.367
R738 B.n111 B.n49 163.367
R739 B.n117 B.n53 163.367
R740 B.n121 B.n120 163.367
R741 B.n125 B.n124 163.367
R742 B.n129 B.n128 163.367
R743 B.n133 B.n132 163.367
R744 B.n137 B.n136 163.367
R745 B.n141 B.n140 163.367
R746 B.n145 B.n144 163.367
R747 B.n149 B.n148 163.367
R748 B.n153 B.n152 163.367
R749 B.n157 B.n156 163.367
R750 B.n161 B.n160 163.367
R751 B.n165 B.n164 163.367
R752 B.n169 B.n168 163.367
R753 B.n173 B.n172 163.367
R754 B.n177 B.n176 163.367
R755 B.n181 B.n180 163.367
R756 B.n185 B.n184 163.367
R757 B.n189 B.n188 163.367
R758 B.n193 B.n192 163.367
R759 B.n197 B.n196 163.367
R760 B.n201 B.n200 163.367
R761 B.n205 B.n204 163.367
R762 B.n209 B.n208 163.367
R763 B.n213 B.n212 163.367
R764 B.n217 B.n216 163.367
R765 B.n222 B.n221 163.367
R766 B.n226 B.n225 163.367
R767 B.n230 B.n229 163.367
R768 B.n234 B.n233 163.367
R769 B.n238 B.n237 163.367
R770 B.n242 B.n241 163.367
R771 B.n246 B.n245 163.367
R772 B.n250 B.n249 163.367
R773 B.n254 B.n253 163.367
R774 B.n258 B.n257 163.367
R775 B.n262 B.n261 163.367
R776 B.n266 B.n265 163.367
R777 B.n270 B.n269 163.367
R778 B.n274 B.n273 163.367
R779 B.n278 B.n277 163.367
R780 B.n282 B.n281 163.367
R781 B.n286 B.n285 163.367
R782 B.n290 B.n289 163.367
R783 B.n294 B.n293 163.367
R784 B.n298 B.n297 163.367
R785 B.n302 B.n301 163.367
R786 B.n306 B.n305 163.367
R787 B.n310 B.n309 163.367
R788 B.n314 B.n313 163.367
R789 B.n318 B.n317 163.367
R790 B.n322 B.n321 163.367
R791 B.n326 B.n325 163.367
R792 B.n330 B.n329 163.367
R793 B.n334 B.n333 163.367
R794 B.n338 B.n337 163.367
R795 B.n802 B.n110 163.367
R796 B.n455 B.t14 113.165
R797 B.n112 B.t9 113.165
R798 B.n452 B.t17 113.145
R799 B.n115 B.t6 113.145
R800 B.n683 B.n391 73.4902
R801 B.n803 B.n50 73.4902
R802 B.n685 B.n684 71.676
R803 B.n451 B.n395 71.676
R804 B.n677 B.n396 71.676
R805 B.n673 B.n397 71.676
R806 B.n669 B.n398 71.676
R807 B.n665 B.n399 71.676
R808 B.n661 B.n400 71.676
R809 B.n657 B.n401 71.676
R810 B.n653 B.n402 71.676
R811 B.n649 B.n403 71.676
R812 B.n645 B.n404 71.676
R813 B.n641 B.n405 71.676
R814 B.n637 B.n406 71.676
R815 B.n633 B.n407 71.676
R816 B.n629 B.n408 71.676
R817 B.n625 B.n409 71.676
R818 B.n621 B.n410 71.676
R819 B.n617 B.n411 71.676
R820 B.n613 B.n412 71.676
R821 B.n609 B.n413 71.676
R822 B.n605 B.n414 71.676
R823 B.n601 B.n415 71.676
R824 B.n597 B.n416 71.676
R825 B.n593 B.n417 71.676
R826 B.n589 B.n418 71.676
R827 B.n585 B.n419 71.676
R828 B.n581 B.n420 71.676
R829 B.n577 B.n421 71.676
R830 B.n573 B.n422 71.676
R831 B.n569 B.n423 71.676
R832 B.n565 B.n424 71.676
R833 B.n560 B.n425 71.676
R834 B.n556 B.n426 71.676
R835 B.n552 B.n427 71.676
R836 B.n548 B.n428 71.676
R837 B.n544 B.n429 71.676
R838 B.n540 B.n430 71.676
R839 B.n536 B.n431 71.676
R840 B.n532 B.n432 71.676
R841 B.n528 B.n433 71.676
R842 B.n524 B.n434 71.676
R843 B.n520 B.n435 71.676
R844 B.n516 B.n436 71.676
R845 B.n512 B.n437 71.676
R846 B.n508 B.n438 71.676
R847 B.n504 B.n439 71.676
R848 B.n500 B.n440 71.676
R849 B.n496 B.n441 71.676
R850 B.n492 B.n442 71.676
R851 B.n488 B.n443 71.676
R852 B.n484 B.n444 71.676
R853 B.n480 B.n445 71.676
R854 B.n476 B.n446 71.676
R855 B.n472 B.n447 71.676
R856 B.n468 B.n448 71.676
R857 B.n464 B.n449 71.676
R858 B.n460 B.n450 71.676
R859 B.n805 B.n804 71.676
R860 B.n117 B.n54 71.676
R861 B.n121 B.n55 71.676
R862 B.n125 B.n56 71.676
R863 B.n129 B.n57 71.676
R864 B.n133 B.n58 71.676
R865 B.n137 B.n59 71.676
R866 B.n141 B.n60 71.676
R867 B.n145 B.n61 71.676
R868 B.n149 B.n62 71.676
R869 B.n153 B.n63 71.676
R870 B.n157 B.n64 71.676
R871 B.n161 B.n65 71.676
R872 B.n165 B.n66 71.676
R873 B.n169 B.n67 71.676
R874 B.n173 B.n68 71.676
R875 B.n177 B.n69 71.676
R876 B.n181 B.n70 71.676
R877 B.n185 B.n71 71.676
R878 B.n189 B.n72 71.676
R879 B.n193 B.n73 71.676
R880 B.n197 B.n74 71.676
R881 B.n201 B.n75 71.676
R882 B.n205 B.n76 71.676
R883 B.n209 B.n77 71.676
R884 B.n213 B.n78 71.676
R885 B.n217 B.n79 71.676
R886 B.n222 B.n80 71.676
R887 B.n226 B.n81 71.676
R888 B.n230 B.n82 71.676
R889 B.n234 B.n83 71.676
R890 B.n238 B.n84 71.676
R891 B.n242 B.n85 71.676
R892 B.n246 B.n86 71.676
R893 B.n250 B.n87 71.676
R894 B.n254 B.n88 71.676
R895 B.n258 B.n89 71.676
R896 B.n262 B.n90 71.676
R897 B.n266 B.n91 71.676
R898 B.n270 B.n92 71.676
R899 B.n274 B.n93 71.676
R900 B.n278 B.n94 71.676
R901 B.n282 B.n95 71.676
R902 B.n286 B.n96 71.676
R903 B.n290 B.n97 71.676
R904 B.n294 B.n98 71.676
R905 B.n298 B.n99 71.676
R906 B.n302 B.n100 71.676
R907 B.n306 B.n101 71.676
R908 B.n310 B.n102 71.676
R909 B.n314 B.n103 71.676
R910 B.n318 B.n104 71.676
R911 B.n322 B.n105 71.676
R912 B.n326 B.n106 71.676
R913 B.n330 B.n107 71.676
R914 B.n334 B.n108 71.676
R915 B.n338 B.n109 71.676
R916 B.n110 B.n109 71.676
R917 B.n337 B.n108 71.676
R918 B.n333 B.n107 71.676
R919 B.n329 B.n106 71.676
R920 B.n325 B.n105 71.676
R921 B.n321 B.n104 71.676
R922 B.n317 B.n103 71.676
R923 B.n313 B.n102 71.676
R924 B.n309 B.n101 71.676
R925 B.n305 B.n100 71.676
R926 B.n301 B.n99 71.676
R927 B.n297 B.n98 71.676
R928 B.n293 B.n97 71.676
R929 B.n289 B.n96 71.676
R930 B.n285 B.n95 71.676
R931 B.n281 B.n94 71.676
R932 B.n277 B.n93 71.676
R933 B.n273 B.n92 71.676
R934 B.n269 B.n91 71.676
R935 B.n265 B.n90 71.676
R936 B.n261 B.n89 71.676
R937 B.n257 B.n88 71.676
R938 B.n253 B.n87 71.676
R939 B.n249 B.n86 71.676
R940 B.n245 B.n85 71.676
R941 B.n241 B.n84 71.676
R942 B.n237 B.n83 71.676
R943 B.n233 B.n82 71.676
R944 B.n229 B.n81 71.676
R945 B.n225 B.n80 71.676
R946 B.n221 B.n79 71.676
R947 B.n216 B.n78 71.676
R948 B.n212 B.n77 71.676
R949 B.n208 B.n76 71.676
R950 B.n204 B.n75 71.676
R951 B.n200 B.n74 71.676
R952 B.n196 B.n73 71.676
R953 B.n192 B.n72 71.676
R954 B.n188 B.n71 71.676
R955 B.n184 B.n70 71.676
R956 B.n180 B.n69 71.676
R957 B.n176 B.n68 71.676
R958 B.n172 B.n67 71.676
R959 B.n168 B.n66 71.676
R960 B.n164 B.n65 71.676
R961 B.n160 B.n64 71.676
R962 B.n156 B.n63 71.676
R963 B.n152 B.n62 71.676
R964 B.n148 B.n61 71.676
R965 B.n144 B.n60 71.676
R966 B.n140 B.n59 71.676
R967 B.n136 B.n58 71.676
R968 B.n132 B.n57 71.676
R969 B.n128 B.n56 71.676
R970 B.n124 B.n55 71.676
R971 B.n120 B.n54 71.676
R972 B.n804 B.n53 71.676
R973 B.n684 B.n394 71.676
R974 B.n678 B.n395 71.676
R975 B.n674 B.n396 71.676
R976 B.n670 B.n397 71.676
R977 B.n666 B.n398 71.676
R978 B.n662 B.n399 71.676
R979 B.n658 B.n400 71.676
R980 B.n654 B.n401 71.676
R981 B.n650 B.n402 71.676
R982 B.n646 B.n403 71.676
R983 B.n642 B.n404 71.676
R984 B.n638 B.n405 71.676
R985 B.n634 B.n406 71.676
R986 B.n630 B.n407 71.676
R987 B.n626 B.n408 71.676
R988 B.n622 B.n409 71.676
R989 B.n618 B.n410 71.676
R990 B.n614 B.n411 71.676
R991 B.n610 B.n412 71.676
R992 B.n606 B.n413 71.676
R993 B.n602 B.n414 71.676
R994 B.n598 B.n415 71.676
R995 B.n594 B.n416 71.676
R996 B.n590 B.n417 71.676
R997 B.n586 B.n418 71.676
R998 B.n582 B.n419 71.676
R999 B.n578 B.n420 71.676
R1000 B.n574 B.n421 71.676
R1001 B.n570 B.n422 71.676
R1002 B.n566 B.n423 71.676
R1003 B.n561 B.n424 71.676
R1004 B.n557 B.n425 71.676
R1005 B.n553 B.n426 71.676
R1006 B.n549 B.n427 71.676
R1007 B.n545 B.n428 71.676
R1008 B.n541 B.n429 71.676
R1009 B.n537 B.n430 71.676
R1010 B.n533 B.n431 71.676
R1011 B.n529 B.n432 71.676
R1012 B.n525 B.n433 71.676
R1013 B.n521 B.n434 71.676
R1014 B.n517 B.n435 71.676
R1015 B.n513 B.n436 71.676
R1016 B.n509 B.n437 71.676
R1017 B.n505 B.n438 71.676
R1018 B.n501 B.n439 71.676
R1019 B.n497 B.n440 71.676
R1020 B.n493 B.n441 71.676
R1021 B.n489 B.n442 71.676
R1022 B.n485 B.n443 71.676
R1023 B.n481 B.n444 71.676
R1024 B.n477 B.n445 71.676
R1025 B.n473 B.n446 71.676
R1026 B.n469 B.n447 71.676
R1027 B.n465 B.n448 71.676
R1028 B.n461 B.n449 71.676
R1029 B.n457 B.n450 71.676
R1030 B.n456 B.t13 71.081
R1031 B.n113 B.t10 71.081
R1032 B.n453 B.t16 71.0603
R1033 B.n116 B.t7 71.0603
R1034 B.n563 B.n456 59.5399
R1035 B.n454 B.n453 59.5399
R1036 B.n219 B.n116 59.5399
R1037 B.n114 B.n113 59.5399
R1038 B.n456 B.n455 42.0853
R1039 B.n453 B.n452 42.0853
R1040 B.n116 B.n115 42.0853
R1041 B.n113 B.n112 42.0853
R1042 B.n807 B.n806 36.9956
R1043 B.n801 B.n800 36.9956
R1044 B.n458 B.n389 36.9956
R1045 B.n687 B.n686 36.9956
R1046 B.n690 B.n391 35.4423
R1047 B.n690 B.n387 35.4423
R1048 B.n696 B.n387 35.4423
R1049 B.n696 B.n382 35.4423
R1050 B.n702 B.n382 35.4423
R1051 B.n702 B.n383 35.4423
R1052 B.n708 B.n375 35.4423
R1053 B.n714 B.n375 35.4423
R1054 B.n714 B.n371 35.4423
R1055 B.n720 B.n371 35.4423
R1056 B.n720 B.n367 35.4423
R1057 B.n726 B.n367 35.4423
R1058 B.n726 B.n363 35.4423
R1059 B.n732 B.n363 35.4423
R1060 B.n738 B.n359 35.4423
R1061 B.n738 B.n355 35.4423
R1062 B.n744 B.n355 35.4423
R1063 B.n744 B.n350 35.4423
R1064 B.n750 B.n350 35.4423
R1065 B.n750 B.n351 35.4423
R1066 B.n757 B.n343 35.4423
R1067 B.n763 B.n343 35.4423
R1068 B.n763 B.n4 35.4423
R1069 B.n860 B.n4 35.4423
R1070 B.n860 B.n859 35.4423
R1071 B.n859 B.n858 35.4423
R1072 B.n858 B.n8 35.4423
R1073 B.n852 B.n8 35.4423
R1074 B.n851 B.n850 35.4423
R1075 B.n850 B.n15 35.4423
R1076 B.n844 B.n15 35.4423
R1077 B.n844 B.n843 35.4423
R1078 B.n843 B.n842 35.4423
R1079 B.n842 B.n22 35.4423
R1080 B.n836 B.n835 35.4423
R1081 B.n835 B.n834 35.4423
R1082 B.n834 B.n29 35.4423
R1083 B.n828 B.n29 35.4423
R1084 B.n828 B.n827 35.4423
R1085 B.n827 B.n826 35.4423
R1086 B.n826 B.n36 35.4423
R1087 B.n820 B.n36 35.4423
R1088 B.n819 B.n818 35.4423
R1089 B.n818 B.n43 35.4423
R1090 B.n812 B.n43 35.4423
R1091 B.n812 B.n811 35.4423
R1092 B.n811 B.n810 35.4423
R1093 B.n810 B.n50 35.4423
R1094 B.n732 B.t0 29.1879
R1095 B.n836 B.t3 29.1879
R1096 B.n757 B.t2 28.1455
R1097 B.n852 B.t1 28.1455
R1098 B.n708 B.t12 27.1031
R1099 B.n820 B.t5 27.1031
R1100 B B.n862 18.0485
R1101 B.n806 B.n52 10.6151
R1102 B.n118 B.n52 10.6151
R1103 B.n119 B.n118 10.6151
R1104 B.n122 B.n119 10.6151
R1105 B.n123 B.n122 10.6151
R1106 B.n126 B.n123 10.6151
R1107 B.n127 B.n126 10.6151
R1108 B.n130 B.n127 10.6151
R1109 B.n131 B.n130 10.6151
R1110 B.n134 B.n131 10.6151
R1111 B.n135 B.n134 10.6151
R1112 B.n138 B.n135 10.6151
R1113 B.n139 B.n138 10.6151
R1114 B.n142 B.n139 10.6151
R1115 B.n143 B.n142 10.6151
R1116 B.n146 B.n143 10.6151
R1117 B.n147 B.n146 10.6151
R1118 B.n150 B.n147 10.6151
R1119 B.n151 B.n150 10.6151
R1120 B.n154 B.n151 10.6151
R1121 B.n155 B.n154 10.6151
R1122 B.n158 B.n155 10.6151
R1123 B.n159 B.n158 10.6151
R1124 B.n162 B.n159 10.6151
R1125 B.n163 B.n162 10.6151
R1126 B.n166 B.n163 10.6151
R1127 B.n167 B.n166 10.6151
R1128 B.n170 B.n167 10.6151
R1129 B.n171 B.n170 10.6151
R1130 B.n174 B.n171 10.6151
R1131 B.n175 B.n174 10.6151
R1132 B.n178 B.n175 10.6151
R1133 B.n179 B.n178 10.6151
R1134 B.n182 B.n179 10.6151
R1135 B.n183 B.n182 10.6151
R1136 B.n186 B.n183 10.6151
R1137 B.n187 B.n186 10.6151
R1138 B.n190 B.n187 10.6151
R1139 B.n191 B.n190 10.6151
R1140 B.n194 B.n191 10.6151
R1141 B.n195 B.n194 10.6151
R1142 B.n198 B.n195 10.6151
R1143 B.n199 B.n198 10.6151
R1144 B.n202 B.n199 10.6151
R1145 B.n203 B.n202 10.6151
R1146 B.n206 B.n203 10.6151
R1147 B.n207 B.n206 10.6151
R1148 B.n210 B.n207 10.6151
R1149 B.n211 B.n210 10.6151
R1150 B.n214 B.n211 10.6151
R1151 B.n215 B.n214 10.6151
R1152 B.n218 B.n215 10.6151
R1153 B.n223 B.n220 10.6151
R1154 B.n224 B.n223 10.6151
R1155 B.n227 B.n224 10.6151
R1156 B.n228 B.n227 10.6151
R1157 B.n231 B.n228 10.6151
R1158 B.n232 B.n231 10.6151
R1159 B.n235 B.n232 10.6151
R1160 B.n236 B.n235 10.6151
R1161 B.n240 B.n239 10.6151
R1162 B.n243 B.n240 10.6151
R1163 B.n244 B.n243 10.6151
R1164 B.n247 B.n244 10.6151
R1165 B.n248 B.n247 10.6151
R1166 B.n251 B.n248 10.6151
R1167 B.n252 B.n251 10.6151
R1168 B.n255 B.n252 10.6151
R1169 B.n256 B.n255 10.6151
R1170 B.n259 B.n256 10.6151
R1171 B.n260 B.n259 10.6151
R1172 B.n263 B.n260 10.6151
R1173 B.n264 B.n263 10.6151
R1174 B.n267 B.n264 10.6151
R1175 B.n268 B.n267 10.6151
R1176 B.n271 B.n268 10.6151
R1177 B.n272 B.n271 10.6151
R1178 B.n275 B.n272 10.6151
R1179 B.n276 B.n275 10.6151
R1180 B.n279 B.n276 10.6151
R1181 B.n280 B.n279 10.6151
R1182 B.n283 B.n280 10.6151
R1183 B.n284 B.n283 10.6151
R1184 B.n287 B.n284 10.6151
R1185 B.n288 B.n287 10.6151
R1186 B.n291 B.n288 10.6151
R1187 B.n292 B.n291 10.6151
R1188 B.n295 B.n292 10.6151
R1189 B.n296 B.n295 10.6151
R1190 B.n299 B.n296 10.6151
R1191 B.n300 B.n299 10.6151
R1192 B.n303 B.n300 10.6151
R1193 B.n304 B.n303 10.6151
R1194 B.n307 B.n304 10.6151
R1195 B.n308 B.n307 10.6151
R1196 B.n311 B.n308 10.6151
R1197 B.n312 B.n311 10.6151
R1198 B.n315 B.n312 10.6151
R1199 B.n316 B.n315 10.6151
R1200 B.n319 B.n316 10.6151
R1201 B.n320 B.n319 10.6151
R1202 B.n323 B.n320 10.6151
R1203 B.n324 B.n323 10.6151
R1204 B.n327 B.n324 10.6151
R1205 B.n328 B.n327 10.6151
R1206 B.n331 B.n328 10.6151
R1207 B.n332 B.n331 10.6151
R1208 B.n335 B.n332 10.6151
R1209 B.n336 B.n335 10.6151
R1210 B.n339 B.n336 10.6151
R1211 B.n340 B.n339 10.6151
R1212 B.n801 B.n340 10.6151
R1213 B.n692 B.n389 10.6151
R1214 B.n693 B.n692 10.6151
R1215 B.n694 B.n693 10.6151
R1216 B.n694 B.n380 10.6151
R1217 B.n704 B.n380 10.6151
R1218 B.n705 B.n704 10.6151
R1219 B.n706 B.n705 10.6151
R1220 B.n706 B.n373 10.6151
R1221 B.n716 B.n373 10.6151
R1222 B.n717 B.n716 10.6151
R1223 B.n718 B.n717 10.6151
R1224 B.n718 B.n365 10.6151
R1225 B.n728 B.n365 10.6151
R1226 B.n729 B.n728 10.6151
R1227 B.n730 B.n729 10.6151
R1228 B.n730 B.n357 10.6151
R1229 B.n740 B.n357 10.6151
R1230 B.n741 B.n740 10.6151
R1231 B.n742 B.n741 10.6151
R1232 B.n742 B.n348 10.6151
R1233 B.n752 B.n348 10.6151
R1234 B.n753 B.n752 10.6151
R1235 B.n755 B.n753 10.6151
R1236 B.n755 B.n754 10.6151
R1237 B.n754 B.n341 10.6151
R1238 B.n766 B.n341 10.6151
R1239 B.n767 B.n766 10.6151
R1240 B.n768 B.n767 10.6151
R1241 B.n769 B.n768 10.6151
R1242 B.n771 B.n769 10.6151
R1243 B.n772 B.n771 10.6151
R1244 B.n773 B.n772 10.6151
R1245 B.n774 B.n773 10.6151
R1246 B.n776 B.n774 10.6151
R1247 B.n777 B.n776 10.6151
R1248 B.n778 B.n777 10.6151
R1249 B.n779 B.n778 10.6151
R1250 B.n781 B.n779 10.6151
R1251 B.n782 B.n781 10.6151
R1252 B.n783 B.n782 10.6151
R1253 B.n784 B.n783 10.6151
R1254 B.n786 B.n784 10.6151
R1255 B.n787 B.n786 10.6151
R1256 B.n788 B.n787 10.6151
R1257 B.n789 B.n788 10.6151
R1258 B.n791 B.n789 10.6151
R1259 B.n792 B.n791 10.6151
R1260 B.n793 B.n792 10.6151
R1261 B.n794 B.n793 10.6151
R1262 B.n796 B.n794 10.6151
R1263 B.n797 B.n796 10.6151
R1264 B.n798 B.n797 10.6151
R1265 B.n799 B.n798 10.6151
R1266 B.n800 B.n799 10.6151
R1267 B.n686 B.n393 10.6151
R1268 B.n681 B.n393 10.6151
R1269 B.n681 B.n680 10.6151
R1270 B.n680 B.n679 10.6151
R1271 B.n679 B.n676 10.6151
R1272 B.n676 B.n675 10.6151
R1273 B.n675 B.n672 10.6151
R1274 B.n672 B.n671 10.6151
R1275 B.n671 B.n668 10.6151
R1276 B.n668 B.n667 10.6151
R1277 B.n667 B.n664 10.6151
R1278 B.n664 B.n663 10.6151
R1279 B.n663 B.n660 10.6151
R1280 B.n660 B.n659 10.6151
R1281 B.n659 B.n656 10.6151
R1282 B.n656 B.n655 10.6151
R1283 B.n655 B.n652 10.6151
R1284 B.n652 B.n651 10.6151
R1285 B.n651 B.n648 10.6151
R1286 B.n648 B.n647 10.6151
R1287 B.n647 B.n644 10.6151
R1288 B.n644 B.n643 10.6151
R1289 B.n643 B.n640 10.6151
R1290 B.n640 B.n639 10.6151
R1291 B.n639 B.n636 10.6151
R1292 B.n636 B.n635 10.6151
R1293 B.n635 B.n632 10.6151
R1294 B.n632 B.n631 10.6151
R1295 B.n631 B.n628 10.6151
R1296 B.n628 B.n627 10.6151
R1297 B.n627 B.n624 10.6151
R1298 B.n624 B.n623 10.6151
R1299 B.n623 B.n620 10.6151
R1300 B.n620 B.n619 10.6151
R1301 B.n619 B.n616 10.6151
R1302 B.n616 B.n615 10.6151
R1303 B.n615 B.n612 10.6151
R1304 B.n612 B.n611 10.6151
R1305 B.n611 B.n608 10.6151
R1306 B.n608 B.n607 10.6151
R1307 B.n607 B.n604 10.6151
R1308 B.n604 B.n603 10.6151
R1309 B.n603 B.n600 10.6151
R1310 B.n600 B.n599 10.6151
R1311 B.n599 B.n596 10.6151
R1312 B.n596 B.n595 10.6151
R1313 B.n595 B.n592 10.6151
R1314 B.n592 B.n591 10.6151
R1315 B.n591 B.n588 10.6151
R1316 B.n588 B.n587 10.6151
R1317 B.n587 B.n584 10.6151
R1318 B.n584 B.n583 10.6151
R1319 B.n580 B.n579 10.6151
R1320 B.n579 B.n576 10.6151
R1321 B.n576 B.n575 10.6151
R1322 B.n575 B.n572 10.6151
R1323 B.n572 B.n571 10.6151
R1324 B.n571 B.n568 10.6151
R1325 B.n568 B.n567 10.6151
R1326 B.n567 B.n564 10.6151
R1327 B.n562 B.n559 10.6151
R1328 B.n559 B.n558 10.6151
R1329 B.n558 B.n555 10.6151
R1330 B.n555 B.n554 10.6151
R1331 B.n554 B.n551 10.6151
R1332 B.n551 B.n550 10.6151
R1333 B.n550 B.n547 10.6151
R1334 B.n547 B.n546 10.6151
R1335 B.n546 B.n543 10.6151
R1336 B.n543 B.n542 10.6151
R1337 B.n542 B.n539 10.6151
R1338 B.n539 B.n538 10.6151
R1339 B.n538 B.n535 10.6151
R1340 B.n535 B.n534 10.6151
R1341 B.n534 B.n531 10.6151
R1342 B.n531 B.n530 10.6151
R1343 B.n530 B.n527 10.6151
R1344 B.n527 B.n526 10.6151
R1345 B.n526 B.n523 10.6151
R1346 B.n523 B.n522 10.6151
R1347 B.n522 B.n519 10.6151
R1348 B.n519 B.n518 10.6151
R1349 B.n518 B.n515 10.6151
R1350 B.n515 B.n514 10.6151
R1351 B.n514 B.n511 10.6151
R1352 B.n511 B.n510 10.6151
R1353 B.n510 B.n507 10.6151
R1354 B.n507 B.n506 10.6151
R1355 B.n506 B.n503 10.6151
R1356 B.n503 B.n502 10.6151
R1357 B.n502 B.n499 10.6151
R1358 B.n499 B.n498 10.6151
R1359 B.n498 B.n495 10.6151
R1360 B.n495 B.n494 10.6151
R1361 B.n494 B.n491 10.6151
R1362 B.n491 B.n490 10.6151
R1363 B.n490 B.n487 10.6151
R1364 B.n487 B.n486 10.6151
R1365 B.n486 B.n483 10.6151
R1366 B.n483 B.n482 10.6151
R1367 B.n482 B.n479 10.6151
R1368 B.n479 B.n478 10.6151
R1369 B.n478 B.n475 10.6151
R1370 B.n475 B.n474 10.6151
R1371 B.n474 B.n471 10.6151
R1372 B.n471 B.n470 10.6151
R1373 B.n470 B.n467 10.6151
R1374 B.n467 B.n466 10.6151
R1375 B.n466 B.n463 10.6151
R1376 B.n463 B.n462 10.6151
R1377 B.n462 B.n459 10.6151
R1378 B.n459 B.n458 10.6151
R1379 B.n688 B.n687 10.6151
R1380 B.n688 B.n385 10.6151
R1381 B.n698 B.n385 10.6151
R1382 B.n699 B.n698 10.6151
R1383 B.n700 B.n699 10.6151
R1384 B.n700 B.n377 10.6151
R1385 B.n710 B.n377 10.6151
R1386 B.n711 B.n710 10.6151
R1387 B.n712 B.n711 10.6151
R1388 B.n712 B.n369 10.6151
R1389 B.n722 B.n369 10.6151
R1390 B.n723 B.n722 10.6151
R1391 B.n724 B.n723 10.6151
R1392 B.n724 B.n361 10.6151
R1393 B.n734 B.n361 10.6151
R1394 B.n735 B.n734 10.6151
R1395 B.n736 B.n735 10.6151
R1396 B.n736 B.n353 10.6151
R1397 B.n746 B.n353 10.6151
R1398 B.n747 B.n746 10.6151
R1399 B.n748 B.n747 10.6151
R1400 B.n748 B.n345 10.6151
R1401 B.n759 B.n345 10.6151
R1402 B.n760 B.n759 10.6151
R1403 B.n761 B.n760 10.6151
R1404 B.n761 B.n0 10.6151
R1405 B.n856 B.n1 10.6151
R1406 B.n856 B.n855 10.6151
R1407 B.n855 B.n854 10.6151
R1408 B.n854 B.n10 10.6151
R1409 B.n848 B.n10 10.6151
R1410 B.n848 B.n847 10.6151
R1411 B.n847 B.n846 10.6151
R1412 B.n846 B.n17 10.6151
R1413 B.n840 B.n17 10.6151
R1414 B.n840 B.n839 10.6151
R1415 B.n839 B.n838 10.6151
R1416 B.n838 B.n24 10.6151
R1417 B.n832 B.n24 10.6151
R1418 B.n832 B.n831 10.6151
R1419 B.n831 B.n830 10.6151
R1420 B.n830 B.n31 10.6151
R1421 B.n824 B.n31 10.6151
R1422 B.n824 B.n823 10.6151
R1423 B.n823 B.n822 10.6151
R1424 B.n822 B.n38 10.6151
R1425 B.n816 B.n38 10.6151
R1426 B.n816 B.n815 10.6151
R1427 B.n815 B.n814 10.6151
R1428 B.n814 B.n45 10.6151
R1429 B.n808 B.n45 10.6151
R1430 B.n808 B.n807 10.6151
R1431 B.n383 B.t12 8.33976
R1432 B.t5 B.n819 8.33976
R1433 B.n351 B.t2 7.29735
R1434 B.t1 B.n851 7.29735
R1435 B.n220 B.n219 6.5566
R1436 B.n236 B.n114 6.5566
R1437 B.n580 B.n454 6.5566
R1438 B.n564 B.n563 6.5566
R1439 B.t0 B.n359 6.25494
R1440 B.t3 B.n22 6.25494
R1441 B.n219 B.n218 4.05904
R1442 B.n239 B.n114 4.05904
R1443 B.n583 B.n454 4.05904
R1444 B.n563 B.n562 4.05904
R1445 B.n862 B.n0 2.81026
R1446 B.n862 B.n1 2.81026
R1447 VP.n3 VP.t3 244.472
R1448 VP.n3 VP.t1 244.038
R1449 VP.n5 VP.t2 207.339
R1450 VP.n13 VP.t0 207.339
R1451 VP.n5 VP.n4 181.608
R1452 VP.n14 VP.n13 181.608
R1453 VP.n12 VP.n0 161.3
R1454 VP.n11 VP.n10 161.3
R1455 VP.n9 VP.n1 161.3
R1456 VP.n8 VP.n7 161.3
R1457 VP.n6 VP.n2 161.3
R1458 VP.n4 VP.n3 56.0406
R1459 VP.n7 VP.n1 40.4934
R1460 VP.n11 VP.n1 40.4934
R1461 VP.n7 VP.n6 24.4675
R1462 VP.n12 VP.n11 24.4675
R1463 VP.n6 VP.n5 4.15989
R1464 VP.n13 VP.n12 4.15989
R1465 VP.n4 VP.n2 0.189894
R1466 VP.n8 VP.n2 0.189894
R1467 VP.n9 VP.n8 0.189894
R1468 VP.n10 VP.n9 0.189894
R1469 VP.n10 VP.n0 0.189894
R1470 VP.n14 VP.n0 0.189894
R1471 VP VP.n14 0.0516364
R1472 VTAIL.n5 VTAIL.t7 47.5136
R1473 VTAIL.n4 VTAIL.t2 47.5136
R1474 VTAIL.n3 VTAIL.t0 47.5136
R1475 VTAIL.n7 VTAIL.t3 47.5135
R1476 VTAIL.n0 VTAIL.t1 47.5135
R1477 VTAIL.n1 VTAIL.t6 47.5135
R1478 VTAIL.n2 VTAIL.t4 47.5135
R1479 VTAIL.n6 VTAIL.t5 47.5135
R1480 VTAIL.n7 VTAIL.n6 27.8841
R1481 VTAIL.n3 VTAIL.n2 27.8841
R1482 VTAIL.n4 VTAIL.n3 1.87119
R1483 VTAIL.n6 VTAIL.n5 1.87119
R1484 VTAIL.n2 VTAIL.n1 1.87119
R1485 VTAIL VTAIL.n0 0.994035
R1486 VTAIL VTAIL.n7 0.877655
R1487 VTAIL.n5 VTAIL.n4 0.470328
R1488 VTAIL.n1 VTAIL.n0 0.470328
R1489 VDD1 VDD1.n1 106.439
R1490 VDD1 VDD1.n0 62.9996
R1491 VDD1.n0 VDD1.t0 1.25129
R1492 VDD1.n0 VDD1.t2 1.25129
R1493 VDD1.n1 VDD1.t1 1.25129
R1494 VDD1.n1 VDD1.t3 1.25129
R1495 VN.n0 VN.t1 244.472
R1496 VN.n1 VN.t2 244.472
R1497 VN.n0 VN.t3 244.038
R1498 VN.n1 VN.t0 244.038
R1499 VN VN.n1 56.4212
R1500 VN VN.n0 9.22048
R1501 VDD2.n2 VDD2.n0 105.915
R1502 VDD2.n2 VDD2.n1 62.9415
R1503 VDD2.n1 VDD2.t3 1.25129
R1504 VDD2.n1 VDD2.t1 1.25129
R1505 VDD2.n0 VDD2.t2 1.25129
R1506 VDD2.n0 VDD2.t0 1.25129
R1507 VDD2 VDD2.n2 0.0586897
C0 VP VTAIL 5.3954f
C1 VDD1 VN 0.148135f
C2 VDD2 VDD1 0.84174f
C3 VP VN 6.35075f
C4 VP VDD2 0.345768f
C5 VN VTAIL 5.3813f
C6 VDD2 VTAIL 6.50658f
C7 VP VDD1 5.93185f
C8 VDD2 VN 5.73476f
C9 VDD1 VTAIL 6.45746f
C10 VDD2 B 3.632475f
C11 VDD1 B 7.92594f
C12 VTAIL B 11.894259f
C13 VN B 9.71694f
C14 VP B 7.563123f
C15 VDD2.t2 B 0.331105f
C16 VDD2.t0 B 0.331105f
C17 VDD2.n0 B 3.75384f
C18 VDD2.t3 B 0.331105f
C19 VDD2.t1 B 0.331105f
C20 VDD2.n1 B 3.00264f
C21 VDD2.n2 B 3.95385f
C22 VN.t1 B 2.60766f
C23 VN.t3 B 2.60586f
C24 VN.n0 B 1.78664f
C25 VN.t2 B 2.60766f
C26 VN.t0 B 2.60586f
C27 VN.n1 B 3.24075f
C28 VDD1.t0 B 0.333857f
C29 VDD1.t2 B 0.333857f
C30 VDD1.n0 B 3.02797f
C31 VDD1.t1 B 0.333857f
C32 VDD1.t3 B 0.333857f
C33 VDD1.n1 B 3.8122f
C34 VTAIL.t1 B 2.17782f
C35 VTAIL.n0 B 0.274971f
C36 VTAIL.t6 B 2.17782f
C37 VTAIL.n1 B 0.31856f
C38 VTAIL.t4 B 2.17782f
C39 VTAIL.n2 B 1.2758f
C40 VTAIL.t0 B 2.17783f
C41 VTAIL.n3 B 1.27579f
C42 VTAIL.t2 B 2.17783f
C43 VTAIL.n4 B 0.318546f
C44 VTAIL.t7 B 2.17783f
C45 VTAIL.n5 B 0.318546f
C46 VTAIL.t5 B 2.17782f
C47 VTAIL.n6 B 1.2758f
C48 VTAIL.t3 B 2.17782f
C49 VTAIL.n7 B 1.22643f
C50 VP.n0 B 0.031129f
C51 VP.t0 B 2.48749f
C52 VP.n1 B 0.025165f
C53 VP.n2 B 0.031129f
C54 VP.t2 B 2.48749f
C55 VP.t3 B 2.64398f
C56 VP.t1 B 2.64215f
C57 VP.n3 B 3.26696f
C58 VP.n4 B 1.85118f
C59 VP.n5 B 0.948791f
C60 VP.n6 B 0.034241f
C61 VP.n7 B 0.061868f
C62 VP.n8 B 0.031129f
C63 VP.n9 B 0.031129f
C64 VP.n10 B 0.031129f
C65 VP.n11 B 0.061868f
C66 VP.n12 B 0.034241f
C67 VP.n13 B 0.948791f
C68 VP.n14 B 0.033334f
.ends

