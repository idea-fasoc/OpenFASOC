* NGSPICE file created from diff_pair_sample_0011.ext - technology: sky130A

.subckt diff_pair_sample_0011 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t3 w_n2274_n1264# sky130_fd_pr__pfet_01v8 ad=0.2442 pd=1.81 as=0.2442 ps=1.81 w=1.48 l=1.3
X1 VTAIL.t5 VN.t0 VDD2.t5 w_n2274_n1264# sky130_fd_pr__pfet_01v8 ad=0.2442 pd=1.81 as=0.2442 ps=1.81 w=1.48 l=1.3
X2 VDD1.t5 VP.t1 VTAIL.t10 w_n2274_n1264# sky130_fd_pr__pfet_01v8 ad=0.5772 pd=3.74 as=0.2442 ps=1.81 w=1.48 l=1.3
X3 B.t11 B.t9 B.t10 w_n2274_n1264# sky130_fd_pr__pfet_01v8 ad=0.5772 pd=3.74 as=0 ps=0 w=1.48 l=1.3
X4 VDD2.t4 VN.t1 VTAIL.t2 w_n2274_n1264# sky130_fd_pr__pfet_01v8 ad=0.5772 pd=3.74 as=0.2442 ps=1.81 w=1.48 l=1.3
X5 VDD2.t3 VN.t2 VTAIL.t0 w_n2274_n1264# sky130_fd_pr__pfet_01v8 ad=0.2442 pd=1.81 as=0.5772 ps=3.74 w=1.48 l=1.3
X6 VDD1.t0 VP.t2 VTAIL.t9 w_n2274_n1264# sky130_fd_pr__pfet_01v8 ad=0.5772 pd=3.74 as=0.2442 ps=1.81 w=1.48 l=1.3
X7 B.t8 B.t6 B.t7 w_n2274_n1264# sky130_fd_pr__pfet_01v8 ad=0.5772 pd=3.74 as=0 ps=0 w=1.48 l=1.3
X8 VTAIL.t4 VN.t3 VDD2.t2 w_n2274_n1264# sky130_fd_pr__pfet_01v8 ad=0.2442 pd=1.81 as=0.2442 ps=1.81 w=1.48 l=1.3
X9 B.t5 B.t3 B.t4 w_n2274_n1264# sky130_fd_pr__pfet_01v8 ad=0.5772 pd=3.74 as=0 ps=0 w=1.48 l=1.3
X10 VDD1.t1 VP.t3 VTAIL.t8 w_n2274_n1264# sky130_fd_pr__pfet_01v8 ad=0.2442 pd=1.81 as=0.5772 ps=3.74 w=1.48 l=1.3
X11 VDD1.t2 VP.t4 VTAIL.t7 w_n2274_n1264# sky130_fd_pr__pfet_01v8 ad=0.2442 pd=1.81 as=0.5772 ps=3.74 w=1.48 l=1.3
X12 VDD2.t1 VN.t4 VTAIL.t3 w_n2274_n1264# sky130_fd_pr__pfet_01v8 ad=0.5772 pd=3.74 as=0.2442 ps=1.81 w=1.48 l=1.3
X13 VTAIL.t6 VP.t5 VDD1.t4 w_n2274_n1264# sky130_fd_pr__pfet_01v8 ad=0.2442 pd=1.81 as=0.2442 ps=1.81 w=1.48 l=1.3
X14 B.t2 B.t0 B.t1 w_n2274_n1264# sky130_fd_pr__pfet_01v8 ad=0.5772 pd=3.74 as=0 ps=0 w=1.48 l=1.3
X15 VDD2.t0 VN.t5 VTAIL.t1 w_n2274_n1264# sky130_fd_pr__pfet_01v8 ad=0.2442 pd=1.81 as=0.5772 ps=3.74 w=1.48 l=1.3
R0 VP.n7 VP.n6 161.3
R1 VP.n8 VP.n3 161.3
R2 VP.n18 VP.n0 161.3
R3 VP.n17 VP.n16 161.3
R4 VP.n15 VP.n14 161.3
R5 VP.n13 VP.n2 161.3
R6 VP.n10 VP.n9 80.6037
R7 VP.n20 VP.n19 80.6037
R8 VP.n12 VP.n11 80.6037
R9 VP.n5 VP.t2 77.6015
R10 VP.n12 VP.t1 58.0259
R11 VP.n19 VP.t4 58.0259
R12 VP.n9 VP.t3 58.0259
R13 VP.n5 VP.n4 45.1847
R14 VP.n11 VP.n10 35.8082
R15 VP.n14 VP.n13 34.0813
R16 VP.n18 VP.n17 34.0813
R17 VP.n8 VP.n7 34.0813
R18 VP.n13 VP.n12 33.5944
R19 VP.n19 VP.n18 33.5944
R20 VP.n9 VP.n8 33.5944
R21 VP.n6 VP.n5 29.3746
R22 VP.n1 VP.t5 27.4374
R23 VP.n4 VP.t0 27.4374
R24 VP.n14 VP.n1 12.1722
R25 VP.n17 VP.n1 12.1722
R26 VP.n7 VP.n4 12.1722
R27 VP.n10 VP.n3 0.285035
R28 VP.n11 VP.n2 0.285035
R29 VP.n20 VP.n0 0.285035
R30 VP.n6 VP.n3 0.189894
R31 VP.n15 VP.n2 0.189894
R32 VP.n16 VP.n15 0.189894
R33 VP.n16 VP.n0 0.189894
R34 VP VP.n20 0.146778
R35 VDD1 VDD1.t0 273.639
R36 VDD1.n1 VDD1.t5 273.526
R37 VDD1.n1 VDD1.n0 250.861
R38 VDD1.n3 VDD1.n2 250.565
R39 VDD1.n3 VDD1.n1 30.8436
R40 VDD1.n2 VDD1.t3 21.9633
R41 VDD1.n2 VDD1.t1 21.9633
R42 VDD1.n0 VDD1.t4 21.9633
R43 VDD1.n0 VDD1.t2 21.9633
R44 VDD1 VDD1.n3 0.293603
R45 VTAIL.n7 VTAIL.t0 255.849
R46 VTAIL.n11 VTAIL.t1 255.849
R47 VTAIL.n2 VTAIL.t7 255.849
R48 VTAIL.n10 VTAIL.t8 255.849
R49 VTAIL.n9 VTAIL.n8 233.886
R50 VTAIL.n6 VTAIL.n5 233.886
R51 VTAIL.n1 VTAIL.n0 233.886
R52 VTAIL.n4 VTAIL.n3 233.886
R53 VTAIL.n0 VTAIL.t2 21.9633
R54 VTAIL.n0 VTAIL.t4 21.9633
R55 VTAIL.n3 VTAIL.t10 21.9633
R56 VTAIL.n3 VTAIL.t6 21.9633
R57 VTAIL.n8 VTAIL.t9 21.9633
R58 VTAIL.n8 VTAIL.t11 21.9633
R59 VTAIL.n5 VTAIL.t3 21.9633
R60 VTAIL.n5 VTAIL.t5 21.9633
R61 VTAIL.n6 VTAIL.n4 16.4531
R62 VTAIL.n11 VTAIL.n10 15.0479
R63 VTAIL.n7 VTAIL.n6 1.40567
R64 VTAIL.n10 VTAIL.n9 1.40567
R65 VTAIL.n4 VTAIL.n2 1.40567
R66 VTAIL.n9 VTAIL.n7 1.17291
R67 VTAIL.n2 VTAIL.n1 1.17291
R68 VTAIL VTAIL.n11 0.99619
R69 VTAIL VTAIL.n1 0.409983
R70 VN.n13 VN.n8 161.3
R71 VN.n12 VN.n11 161.3
R72 VN.n5 VN.n0 161.3
R73 VN.n4 VN.n3 161.3
R74 VN.n15 VN.n14 80.6037
R75 VN.n7 VN.n6 80.6037
R76 VN.n2 VN.t1 77.6015
R77 VN.n10 VN.t2 77.6015
R78 VN.n6 VN.t5 58.0259
R79 VN.n14 VN.t4 58.0259
R80 VN.n2 VN.n1 45.1847
R81 VN.n10 VN.n9 45.1847
R82 VN VN.n15 36.0937
R83 VN.n5 VN.n4 34.0813
R84 VN.n13 VN.n12 34.0813
R85 VN.n6 VN.n5 33.5944
R86 VN.n14 VN.n13 33.5944
R87 VN.n11 VN.n10 29.3746
R88 VN.n3 VN.n2 29.3746
R89 VN.n1 VN.t3 27.4374
R90 VN.n9 VN.t0 27.4374
R91 VN.n4 VN.n1 12.1722
R92 VN.n12 VN.n9 12.1722
R93 VN.n15 VN.n8 0.285035
R94 VN.n7 VN.n0 0.285035
R95 VN.n11 VN.n8 0.189894
R96 VN.n3 VN.n0 0.189894
R97 VN VN.n7 0.146778
R98 VDD2.n1 VDD2.t4 273.526
R99 VDD2.n2 VDD2.t1 272.527
R100 VDD2.n1 VDD2.n0 250.861
R101 VDD2 VDD2.n3 250.857
R102 VDD2.n2 VDD2.n1 29.558
R103 VDD2.n3 VDD2.t5 21.9633
R104 VDD2.n3 VDD2.t3 21.9633
R105 VDD2.n0 VDD2.t2 21.9633
R106 VDD2.n0 VDD2.t0 21.9633
R107 VDD2 VDD2.n2 1.11257
R108 B.n266 B.n265 585
R109 B.n267 B.n34 585
R110 B.n269 B.n268 585
R111 B.n270 B.n33 585
R112 B.n272 B.n271 585
R113 B.n273 B.n32 585
R114 B.n275 B.n274 585
R115 B.n276 B.n31 585
R116 B.n278 B.n277 585
R117 B.n279 B.n30 585
R118 B.n281 B.n280 585
R119 B.n283 B.n27 585
R120 B.n285 B.n284 585
R121 B.n286 B.n26 585
R122 B.n288 B.n287 585
R123 B.n289 B.n25 585
R124 B.n291 B.n290 585
R125 B.n292 B.n24 585
R126 B.n294 B.n293 585
R127 B.n295 B.n21 585
R128 B.n298 B.n297 585
R129 B.n299 B.n20 585
R130 B.n301 B.n300 585
R131 B.n302 B.n19 585
R132 B.n304 B.n303 585
R133 B.n305 B.n18 585
R134 B.n307 B.n306 585
R135 B.n308 B.n17 585
R136 B.n310 B.n309 585
R137 B.n311 B.n16 585
R138 B.n313 B.n312 585
R139 B.n264 B.n35 585
R140 B.n263 B.n262 585
R141 B.n261 B.n36 585
R142 B.n260 B.n259 585
R143 B.n258 B.n37 585
R144 B.n257 B.n256 585
R145 B.n255 B.n38 585
R146 B.n254 B.n253 585
R147 B.n252 B.n39 585
R148 B.n251 B.n250 585
R149 B.n249 B.n40 585
R150 B.n248 B.n247 585
R151 B.n246 B.n41 585
R152 B.n245 B.n244 585
R153 B.n243 B.n42 585
R154 B.n242 B.n241 585
R155 B.n240 B.n43 585
R156 B.n239 B.n238 585
R157 B.n237 B.n44 585
R158 B.n236 B.n235 585
R159 B.n234 B.n45 585
R160 B.n233 B.n232 585
R161 B.n231 B.n46 585
R162 B.n230 B.n229 585
R163 B.n228 B.n47 585
R164 B.n227 B.n226 585
R165 B.n225 B.n48 585
R166 B.n224 B.n223 585
R167 B.n222 B.n49 585
R168 B.n221 B.n220 585
R169 B.n219 B.n50 585
R170 B.n218 B.n217 585
R171 B.n216 B.n51 585
R172 B.n215 B.n214 585
R173 B.n213 B.n52 585
R174 B.n212 B.n211 585
R175 B.n210 B.n53 585
R176 B.n209 B.n208 585
R177 B.n207 B.n54 585
R178 B.n206 B.n205 585
R179 B.n204 B.n55 585
R180 B.n203 B.n202 585
R181 B.n201 B.n56 585
R182 B.n200 B.n199 585
R183 B.n198 B.n57 585
R184 B.n197 B.n196 585
R185 B.n195 B.n58 585
R186 B.n194 B.n193 585
R187 B.n192 B.n59 585
R188 B.n191 B.n190 585
R189 B.n189 B.n60 585
R190 B.n188 B.n187 585
R191 B.n186 B.n61 585
R192 B.n185 B.n184 585
R193 B.n183 B.n62 585
R194 B.n135 B.n82 585
R195 B.n137 B.n136 585
R196 B.n138 B.n81 585
R197 B.n140 B.n139 585
R198 B.n141 B.n80 585
R199 B.n143 B.n142 585
R200 B.n144 B.n79 585
R201 B.n146 B.n145 585
R202 B.n147 B.n78 585
R203 B.n149 B.n148 585
R204 B.n150 B.n75 585
R205 B.n153 B.n152 585
R206 B.n154 B.n74 585
R207 B.n156 B.n155 585
R208 B.n157 B.n73 585
R209 B.n159 B.n158 585
R210 B.n160 B.n72 585
R211 B.n162 B.n161 585
R212 B.n163 B.n71 585
R213 B.n165 B.n164 585
R214 B.n167 B.n166 585
R215 B.n168 B.n67 585
R216 B.n170 B.n169 585
R217 B.n171 B.n66 585
R218 B.n173 B.n172 585
R219 B.n174 B.n65 585
R220 B.n176 B.n175 585
R221 B.n177 B.n64 585
R222 B.n179 B.n178 585
R223 B.n180 B.n63 585
R224 B.n182 B.n181 585
R225 B.n134 B.n133 585
R226 B.n132 B.n83 585
R227 B.n131 B.n130 585
R228 B.n129 B.n84 585
R229 B.n128 B.n127 585
R230 B.n126 B.n85 585
R231 B.n125 B.n124 585
R232 B.n123 B.n86 585
R233 B.n122 B.n121 585
R234 B.n120 B.n87 585
R235 B.n119 B.n118 585
R236 B.n117 B.n88 585
R237 B.n116 B.n115 585
R238 B.n114 B.n89 585
R239 B.n113 B.n112 585
R240 B.n111 B.n90 585
R241 B.n110 B.n109 585
R242 B.n108 B.n91 585
R243 B.n107 B.n106 585
R244 B.n105 B.n92 585
R245 B.n104 B.n103 585
R246 B.n102 B.n93 585
R247 B.n101 B.n100 585
R248 B.n99 B.n94 585
R249 B.n98 B.n97 585
R250 B.n96 B.n95 585
R251 B.n2 B.n0 585
R252 B.n353 B.n1 585
R253 B.n352 B.n351 585
R254 B.n350 B.n3 585
R255 B.n349 B.n348 585
R256 B.n347 B.n4 585
R257 B.n346 B.n345 585
R258 B.n344 B.n5 585
R259 B.n343 B.n342 585
R260 B.n341 B.n6 585
R261 B.n340 B.n339 585
R262 B.n338 B.n7 585
R263 B.n337 B.n336 585
R264 B.n335 B.n8 585
R265 B.n334 B.n333 585
R266 B.n332 B.n9 585
R267 B.n331 B.n330 585
R268 B.n329 B.n10 585
R269 B.n328 B.n327 585
R270 B.n326 B.n11 585
R271 B.n325 B.n324 585
R272 B.n323 B.n12 585
R273 B.n322 B.n321 585
R274 B.n320 B.n13 585
R275 B.n319 B.n318 585
R276 B.n317 B.n14 585
R277 B.n316 B.n315 585
R278 B.n314 B.n15 585
R279 B.n355 B.n354 585
R280 B.n135 B.n134 540.549
R281 B.n312 B.n15 540.549
R282 B.n183 B.n182 540.549
R283 B.n266 B.n35 540.549
R284 B.n68 B.t5 280.964
R285 B.n28 B.t7 280.964
R286 B.n76 B.t11 280.964
R287 B.n22 B.t1 280.964
R288 B.n69 B.t4 249.352
R289 B.n29 B.t8 249.352
R290 B.n77 B.t10 249.352
R291 B.n23 B.t2 249.352
R292 B.n68 B.t3 232.046
R293 B.n76 B.t9 232.046
R294 B.n22 B.t0 232.046
R295 B.n28 B.t6 232.046
R296 B.n134 B.n83 163.367
R297 B.n130 B.n83 163.367
R298 B.n130 B.n129 163.367
R299 B.n129 B.n128 163.367
R300 B.n128 B.n85 163.367
R301 B.n124 B.n85 163.367
R302 B.n124 B.n123 163.367
R303 B.n123 B.n122 163.367
R304 B.n122 B.n87 163.367
R305 B.n118 B.n87 163.367
R306 B.n118 B.n117 163.367
R307 B.n117 B.n116 163.367
R308 B.n116 B.n89 163.367
R309 B.n112 B.n89 163.367
R310 B.n112 B.n111 163.367
R311 B.n111 B.n110 163.367
R312 B.n110 B.n91 163.367
R313 B.n106 B.n91 163.367
R314 B.n106 B.n105 163.367
R315 B.n105 B.n104 163.367
R316 B.n104 B.n93 163.367
R317 B.n100 B.n93 163.367
R318 B.n100 B.n99 163.367
R319 B.n99 B.n98 163.367
R320 B.n98 B.n95 163.367
R321 B.n95 B.n2 163.367
R322 B.n354 B.n2 163.367
R323 B.n354 B.n353 163.367
R324 B.n353 B.n352 163.367
R325 B.n352 B.n3 163.367
R326 B.n348 B.n3 163.367
R327 B.n348 B.n347 163.367
R328 B.n347 B.n346 163.367
R329 B.n346 B.n5 163.367
R330 B.n342 B.n5 163.367
R331 B.n342 B.n341 163.367
R332 B.n341 B.n340 163.367
R333 B.n340 B.n7 163.367
R334 B.n336 B.n7 163.367
R335 B.n336 B.n335 163.367
R336 B.n335 B.n334 163.367
R337 B.n334 B.n9 163.367
R338 B.n330 B.n9 163.367
R339 B.n330 B.n329 163.367
R340 B.n329 B.n328 163.367
R341 B.n328 B.n11 163.367
R342 B.n324 B.n11 163.367
R343 B.n324 B.n323 163.367
R344 B.n323 B.n322 163.367
R345 B.n322 B.n13 163.367
R346 B.n318 B.n13 163.367
R347 B.n318 B.n317 163.367
R348 B.n317 B.n316 163.367
R349 B.n316 B.n15 163.367
R350 B.n136 B.n135 163.367
R351 B.n136 B.n81 163.367
R352 B.n140 B.n81 163.367
R353 B.n141 B.n140 163.367
R354 B.n142 B.n141 163.367
R355 B.n142 B.n79 163.367
R356 B.n146 B.n79 163.367
R357 B.n147 B.n146 163.367
R358 B.n148 B.n147 163.367
R359 B.n148 B.n75 163.367
R360 B.n153 B.n75 163.367
R361 B.n154 B.n153 163.367
R362 B.n155 B.n154 163.367
R363 B.n155 B.n73 163.367
R364 B.n159 B.n73 163.367
R365 B.n160 B.n159 163.367
R366 B.n161 B.n160 163.367
R367 B.n161 B.n71 163.367
R368 B.n165 B.n71 163.367
R369 B.n166 B.n165 163.367
R370 B.n166 B.n67 163.367
R371 B.n170 B.n67 163.367
R372 B.n171 B.n170 163.367
R373 B.n172 B.n171 163.367
R374 B.n172 B.n65 163.367
R375 B.n176 B.n65 163.367
R376 B.n177 B.n176 163.367
R377 B.n178 B.n177 163.367
R378 B.n178 B.n63 163.367
R379 B.n182 B.n63 163.367
R380 B.n184 B.n183 163.367
R381 B.n184 B.n61 163.367
R382 B.n188 B.n61 163.367
R383 B.n189 B.n188 163.367
R384 B.n190 B.n189 163.367
R385 B.n190 B.n59 163.367
R386 B.n194 B.n59 163.367
R387 B.n195 B.n194 163.367
R388 B.n196 B.n195 163.367
R389 B.n196 B.n57 163.367
R390 B.n200 B.n57 163.367
R391 B.n201 B.n200 163.367
R392 B.n202 B.n201 163.367
R393 B.n202 B.n55 163.367
R394 B.n206 B.n55 163.367
R395 B.n207 B.n206 163.367
R396 B.n208 B.n207 163.367
R397 B.n208 B.n53 163.367
R398 B.n212 B.n53 163.367
R399 B.n213 B.n212 163.367
R400 B.n214 B.n213 163.367
R401 B.n214 B.n51 163.367
R402 B.n218 B.n51 163.367
R403 B.n219 B.n218 163.367
R404 B.n220 B.n219 163.367
R405 B.n220 B.n49 163.367
R406 B.n224 B.n49 163.367
R407 B.n225 B.n224 163.367
R408 B.n226 B.n225 163.367
R409 B.n226 B.n47 163.367
R410 B.n230 B.n47 163.367
R411 B.n231 B.n230 163.367
R412 B.n232 B.n231 163.367
R413 B.n232 B.n45 163.367
R414 B.n236 B.n45 163.367
R415 B.n237 B.n236 163.367
R416 B.n238 B.n237 163.367
R417 B.n238 B.n43 163.367
R418 B.n242 B.n43 163.367
R419 B.n243 B.n242 163.367
R420 B.n244 B.n243 163.367
R421 B.n244 B.n41 163.367
R422 B.n248 B.n41 163.367
R423 B.n249 B.n248 163.367
R424 B.n250 B.n249 163.367
R425 B.n250 B.n39 163.367
R426 B.n254 B.n39 163.367
R427 B.n255 B.n254 163.367
R428 B.n256 B.n255 163.367
R429 B.n256 B.n37 163.367
R430 B.n260 B.n37 163.367
R431 B.n261 B.n260 163.367
R432 B.n262 B.n261 163.367
R433 B.n262 B.n35 163.367
R434 B.n312 B.n311 163.367
R435 B.n311 B.n310 163.367
R436 B.n310 B.n17 163.367
R437 B.n306 B.n17 163.367
R438 B.n306 B.n305 163.367
R439 B.n305 B.n304 163.367
R440 B.n304 B.n19 163.367
R441 B.n300 B.n19 163.367
R442 B.n300 B.n299 163.367
R443 B.n299 B.n298 163.367
R444 B.n298 B.n21 163.367
R445 B.n293 B.n21 163.367
R446 B.n293 B.n292 163.367
R447 B.n292 B.n291 163.367
R448 B.n291 B.n25 163.367
R449 B.n287 B.n25 163.367
R450 B.n287 B.n286 163.367
R451 B.n286 B.n285 163.367
R452 B.n285 B.n27 163.367
R453 B.n280 B.n27 163.367
R454 B.n280 B.n279 163.367
R455 B.n279 B.n278 163.367
R456 B.n278 B.n31 163.367
R457 B.n274 B.n31 163.367
R458 B.n274 B.n273 163.367
R459 B.n273 B.n272 163.367
R460 B.n272 B.n33 163.367
R461 B.n268 B.n33 163.367
R462 B.n268 B.n267 163.367
R463 B.n267 B.n266 163.367
R464 B.n70 B.n69 59.5399
R465 B.n151 B.n77 59.5399
R466 B.n296 B.n23 59.5399
R467 B.n282 B.n29 59.5399
R468 B.n314 B.n313 35.1225
R469 B.n265 B.n264 35.1225
R470 B.n181 B.n62 35.1225
R471 B.n133 B.n82 35.1225
R472 B.n69 B.n68 31.6126
R473 B.n77 B.n76 31.6126
R474 B.n23 B.n22 31.6126
R475 B.n29 B.n28 31.6126
R476 B B.n355 18.0485
R477 B.n313 B.n16 10.6151
R478 B.n309 B.n16 10.6151
R479 B.n309 B.n308 10.6151
R480 B.n308 B.n307 10.6151
R481 B.n307 B.n18 10.6151
R482 B.n303 B.n18 10.6151
R483 B.n303 B.n302 10.6151
R484 B.n302 B.n301 10.6151
R485 B.n301 B.n20 10.6151
R486 B.n297 B.n20 10.6151
R487 B.n295 B.n294 10.6151
R488 B.n294 B.n24 10.6151
R489 B.n290 B.n24 10.6151
R490 B.n290 B.n289 10.6151
R491 B.n289 B.n288 10.6151
R492 B.n288 B.n26 10.6151
R493 B.n284 B.n26 10.6151
R494 B.n284 B.n283 10.6151
R495 B.n281 B.n30 10.6151
R496 B.n277 B.n30 10.6151
R497 B.n277 B.n276 10.6151
R498 B.n276 B.n275 10.6151
R499 B.n275 B.n32 10.6151
R500 B.n271 B.n32 10.6151
R501 B.n271 B.n270 10.6151
R502 B.n270 B.n269 10.6151
R503 B.n269 B.n34 10.6151
R504 B.n265 B.n34 10.6151
R505 B.n185 B.n62 10.6151
R506 B.n186 B.n185 10.6151
R507 B.n187 B.n186 10.6151
R508 B.n187 B.n60 10.6151
R509 B.n191 B.n60 10.6151
R510 B.n192 B.n191 10.6151
R511 B.n193 B.n192 10.6151
R512 B.n193 B.n58 10.6151
R513 B.n197 B.n58 10.6151
R514 B.n198 B.n197 10.6151
R515 B.n199 B.n198 10.6151
R516 B.n199 B.n56 10.6151
R517 B.n203 B.n56 10.6151
R518 B.n204 B.n203 10.6151
R519 B.n205 B.n204 10.6151
R520 B.n205 B.n54 10.6151
R521 B.n209 B.n54 10.6151
R522 B.n210 B.n209 10.6151
R523 B.n211 B.n210 10.6151
R524 B.n211 B.n52 10.6151
R525 B.n215 B.n52 10.6151
R526 B.n216 B.n215 10.6151
R527 B.n217 B.n216 10.6151
R528 B.n217 B.n50 10.6151
R529 B.n221 B.n50 10.6151
R530 B.n222 B.n221 10.6151
R531 B.n223 B.n222 10.6151
R532 B.n223 B.n48 10.6151
R533 B.n227 B.n48 10.6151
R534 B.n228 B.n227 10.6151
R535 B.n229 B.n228 10.6151
R536 B.n229 B.n46 10.6151
R537 B.n233 B.n46 10.6151
R538 B.n234 B.n233 10.6151
R539 B.n235 B.n234 10.6151
R540 B.n235 B.n44 10.6151
R541 B.n239 B.n44 10.6151
R542 B.n240 B.n239 10.6151
R543 B.n241 B.n240 10.6151
R544 B.n241 B.n42 10.6151
R545 B.n245 B.n42 10.6151
R546 B.n246 B.n245 10.6151
R547 B.n247 B.n246 10.6151
R548 B.n247 B.n40 10.6151
R549 B.n251 B.n40 10.6151
R550 B.n252 B.n251 10.6151
R551 B.n253 B.n252 10.6151
R552 B.n253 B.n38 10.6151
R553 B.n257 B.n38 10.6151
R554 B.n258 B.n257 10.6151
R555 B.n259 B.n258 10.6151
R556 B.n259 B.n36 10.6151
R557 B.n263 B.n36 10.6151
R558 B.n264 B.n263 10.6151
R559 B.n137 B.n82 10.6151
R560 B.n138 B.n137 10.6151
R561 B.n139 B.n138 10.6151
R562 B.n139 B.n80 10.6151
R563 B.n143 B.n80 10.6151
R564 B.n144 B.n143 10.6151
R565 B.n145 B.n144 10.6151
R566 B.n145 B.n78 10.6151
R567 B.n149 B.n78 10.6151
R568 B.n150 B.n149 10.6151
R569 B.n152 B.n74 10.6151
R570 B.n156 B.n74 10.6151
R571 B.n157 B.n156 10.6151
R572 B.n158 B.n157 10.6151
R573 B.n158 B.n72 10.6151
R574 B.n162 B.n72 10.6151
R575 B.n163 B.n162 10.6151
R576 B.n164 B.n163 10.6151
R577 B.n168 B.n167 10.6151
R578 B.n169 B.n168 10.6151
R579 B.n169 B.n66 10.6151
R580 B.n173 B.n66 10.6151
R581 B.n174 B.n173 10.6151
R582 B.n175 B.n174 10.6151
R583 B.n175 B.n64 10.6151
R584 B.n179 B.n64 10.6151
R585 B.n180 B.n179 10.6151
R586 B.n181 B.n180 10.6151
R587 B.n133 B.n132 10.6151
R588 B.n132 B.n131 10.6151
R589 B.n131 B.n84 10.6151
R590 B.n127 B.n84 10.6151
R591 B.n127 B.n126 10.6151
R592 B.n126 B.n125 10.6151
R593 B.n125 B.n86 10.6151
R594 B.n121 B.n86 10.6151
R595 B.n121 B.n120 10.6151
R596 B.n120 B.n119 10.6151
R597 B.n119 B.n88 10.6151
R598 B.n115 B.n88 10.6151
R599 B.n115 B.n114 10.6151
R600 B.n114 B.n113 10.6151
R601 B.n113 B.n90 10.6151
R602 B.n109 B.n90 10.6151
R603 B.n109 B.n108 10.6151
R604 B.n108 B.n107 10.6151
R605 B.n107 B.n92 10.6151
R606 B.n103 B.n92 10.6151
R607 B.n103 B.n102 10.6151
R608 B.n102 B.n101 10.6151
R609 B.n101 B.n94 10.6151
R610 B.n97 B.n94 10.6151
R611 B.n97 B.n96 10.6151
R612 B.n96 B.n0 10.6151
R613 B.n351 B.n1 10.6151
R614 B.n351 B.n350 10.6151
R615 B.n350 B.n349 10.6151
R616 B.n349 B.n4 10.6151
R617 B.n345 B.n4 10.6151
R618 B.n345 B.n344 10.6151
R619 B.n344 B.n343 10.6151
R620 B.n343 B.n6 10.6151
R621 B.n339 B.n6 10.6151
R622 B.n339 B.n338 10.6151
R623 B.n338 B.n337 10.6151
R624 B.n337 B.n8 10.6151
R625 B.n333 B.n8 10.6151
R626 B.n333 B.n332 10.6151
R627 B.n332 B.n331 10.6151
R628 B.n331 B.n10 10.6151
R629 B.n327 B.n10 10.6151
R630 B.n327 B.n326 10.6151
R631 B.n326 B.n325 10.6151
R632 B.n325 B.n12 10.6151
R633 B.n321 B.n12 10.6151
R634 B.n321 B.n320 10.6151
R635 B.n320 B.n319 10.6151
R636 B.n319 B.n14 10.6151
R637 B.n315 B.n14 10.6151
R638 B.n315 B.n314 10.6151
R639 B.n296 B.n295 6.5566
R640 B.n283 B.n282 6.5566
R641 B.n152 B.n151 6.5566
R642 B.n164 B.n70 6.5566
R643 B.n297 B.n296 4.05904
R644 B.n282 B.n281 4.05904
R645 B.n151 B.n150 4.05904
R646 B.n167 B.n70 4.05904
R647 B.n355 B.n0 2.81026
R648 B.n355 B.n1 2.81026
C0 VN VDD2 1.0092f
C1 VDD1 VP 1.20611f
C2 B VTAIL 0.927251f
C3 w_n2274_n1264# VP 4.05038f
C4 VDD1 VTAIL 3.06186f
C5 w_n2274_n1264# VTAIL 1.27125f
C6 B VN 0.743702f
C7 VDD1 VN 0.155696f
C8 VP VTAIL 1.47832f
C9 VN w_n2274_n1264# 3.76622f
C10 B VDD2 0.984857f
C11 VDD1 VDD2 0.929008f
C12 VN VP 3.72406f
C13 w_n2274_n1264# VDD2 1.24556f
C14 VN VTAIL 1.46417f
C15 VP VDD2 0.354737f
C16 B VDD1 0.941463f
C17 VDD2 VTAIL 3.1061f
C18 B w_n2274_n1264# 4.93942f
C19 VDD1 w_n2274_n1264# 1.2033f
C20 B VP 1.22099f
C21 VDD2 VSUBS 0.755371f
C22 VDD1 VSUBS 1.05747f
C23 VTAIL VSUBS 0.324743f
C24 VN VSUBS 3.94259f
C25 VP VSUBS 1.425422f
C26 B VSUBS 2.336084f
C27 w_n2274_n1264# VSUBS 36.866104f
C28 B.n0 VSUBS 0.005904f
C29 B.n1 VSUBS 0.005904f
C30 B.n2 VSUBS 0.009336f
C31 B.n3 VSUBS 0.009336f
C32 B.n4 VSUBS 0.009336f
C33 B.n5 VSUBS 0.009336f
C34 B.n6 VSUBS 0.009336f
C35 B.n7 VSUBS 0.009336f
C36 B.n8 VSUBS 0.009336f
C37 B.n9 VSUBS 0.009336f
C38 B.n10 VSUBS 0.009336f
C39 B.n11 VSUBS 0.009336f
C40 B.n12 VSUBS 0.009336f
C41 B.n13 VSUBS 0.009336f
C42 B.n14 VSUBS 0.009336f
C43 B.n15 VSUBS 0.022166f
C44 B.n16 VSUBS 0.009336f
C45 B.n17 VSUBS 0.009336f
C46 B.n18 VSUBS 0.009336f
C47 B.n19 VSUBS 0.009336f
C48 B.n20 VSUBS 0.009336f
C49 B.n21 VSUBS 0.009336f
C50 B.t2 VSUBS 0.040024f
C51 B.t1 VSUBS 0.045596f
C52 B.t0 VSUBS 0.126971f
C53 B.n22 VSUBS 0.071143f
C54 B.n23 VSUBS 0.062838f
C55 B.n24 VSUBS 0.009336f
C56 B.n25 VSUBS 0.009336f
C57 B.n26 VSUBS 0.009336f
C58 B.n27 VSUBS 0.009336f
C59 B.t8 VSUBS 0.040024f
C60 B.t7 VSUBS 0.045596f
C61 B.t6 VSUBS 0.126971f
C62 B.n28 VSUBS 0.071143f
C63 B.n29 VSUBS 0.062838f
C64 B.n30 VSUBS 0.009336f
C65 B.n31 VSUBS 0.009336f
C66 B.n32 VSUBS 0.009336f
C67 B.n33 VSUBS 0.009336f
C68 B.n34 VSUBS 0.009336f
C69 B.n35 VSUBS 0.022166f
C70 B.n36 VSUBS 0.009336f
C71 B.n37 VSUBS 0.009336f
C72 B.n38 VSUBS 0.009336f
C73 B.n39 VSUBS 0.009336f
C74 B.n40 VSUBS 0.009336f
C75 B.n41 VSUBS 0.009336f
C76 B.n42 VSUBS 0.009336f
C77 B.n43 VSUBS 0.009336f
C78 B.n44 VSUBS 0.009336f
C79 B.n45 VSUBS 0.009336f
C80 B.n46 VSUBS 0.009336f
C81 B.n47 VSUBS 0.009336f
C82 B.n48 VSUBS 0.009336f
C83 B.n49 VSUBS 0.009336f
C84 B.n50 VSUBS 0.009336f
C85 B.n51 VSUBS 0.009336f
C86 B.n52 VSUBS 0.009336f
C87 B.n53 VSUBS 0.009336f
C88 B.n54 VSUBS 0.009336f
C89 B.n55 VSUBS 0.009336f
C90 B.n56 VSUBS 0.009336f
C91 B.n57 VSUBS 0.009336f
C92 B.n58 VSUBS 0.009336f
C93 B.n59 VSUBS 0.009336f
C94 B.n60 VSUBS 0.009336f
C95 B.n61 VSUBS 0.009336f
C96 B.n62 VSUBS 0.022166f
C97 B.n63 VSUBS 0.009336f
C98 B.n64 VSUBS 0.009336f
C99 B.n65 VSUBS 0.009336f
C100 B.n66 VSUBS 0.009336f
C101 B.n67 VSUBS 0.009336f
C102 B.t4 VSUBS 0.040024f
C103 B.t5 VSUBS 0.045596f
C104 B.t3 VSUBS 0.126971f
C105 B.n68 VSUBS 0.071143f
C106 B.n69 VSUBS 0.062838f
C107 B.n70 VSUBS 0.021631f
C108 B.n71 VSUBS 0.009336f
C109 B.n72 VSUBS 0.009336f
C110 B.n73 VSUBS 0.009336f
C111 B.n74 VSUBS 0.009336f
C112 B.n75 VSUBS 0.009336f
C113 B.t10 VSUBS 0.040024f
C114 B.t11 VSUBS 0.045596f
C115 B.t9 VSUBS 0.126971f
C116 B.n76 VSUBS 0.071143f
C117 B.n77 VSUBS 0.062838f
C118 B.n78 VSUBS 0.009336f
C119 B.n79 VSUBS 0.009336f
C120 B.n80 VSUBS 0.009336f
C121 B.n81 VSUBS 0.009336f
C122 B.n82 VSUBS 0.023692f
C123 B.n83 VSUBS 0.009336f
C124 B.n84 VSUBS 0.009336f
C125 B.n85 VSUBS 0.009336f
C126 B.n86 VSUBS 0.009336f
C127 B.n87 VSUBS 0.009336f
C128 B.n88 VSUBS 0.009336f
C129 B.n89 VSUBS 0.009336f
C130 B.n90 VSUBS 0.009336f
C131 B.n91 VSUBS 0.009336f
C132 B.n92 VSUBS 0.009336f
C133 B.n93 VSUBS 0.009336f
C134 B.n94 VSUBS 0.009336f
C135 B.n95 VSUBS 0.009336f
C136 B.n96 VSUBS 0.009336f
C137 B.n97 VSUBS 0.009336f
C138 B.n98 VSUBS 0.009336f
C139 B.n99 VSUBS 0.009336f
C140 B.n100 VSUBS 0.009336f
C141 B.n101 VSUBS 0.009336f
C142 B.n102 VSUBS 0.009336f
C143 B.n103 VSUBS 0.009336f
C144 B.n104 VSUBS 0.009336f
C145 B.n105 VSUBS 0.009336f
C146 B.n106 VSUBS 0.009336f
C147 B.n107 VSUBS 0.009336f
C148 B.n108 VSUBS 0.009336f
C149 B.n109 VSUBS 0.009336f
C150 B.n110 VSUBS 0.009336f
C151 B.n111 VSUBS 0.009336f
C152 B.n112 VSUBS 0.009336f
C153 B.n113 VSUBS 0.009336f
C154 B.n114 VSUBS 0.009336f
C155 B.n115 VSUBS 0.009336f
C156 B.n116 VSUBS 0.009336f
C157 B.n117 VSUBS 0.009336f
C158 B.n118 VSUBS 0.009336f
C159 B.n119 VSUBS 0.009336f
C160 B.n120 VSUBS 0.009336f
C161 B.n121 VSUBS 0.009336f
C162 B.n122 VSUBS 0.009336f
C163 B.n123 VSUBS 0.009336f
C164 B.n124 VSUBS 0.009336f
C165 B.n125 VSUBS 0.009336f
C166 B.n126 VSUBS 0.009336f
C167 B.n127 VSUBS 0.009336f
C168 B.n128 VSUBS 0.009336f
C169 B.n129 VSUBS 0.009336f
C170 B.n130 VSUBS 0.009336f
C171 B.n131 VSUBS 0.009336f
C172 B.n132 VSUBS 0.009336f
C173 B.n133 VSUBS 0.022166f
C174 B.n134 VSUBS 0.022166f
C175 B.n135 VSUBS 0.023692f
C176 B.n136 VSUBS 0.009336f
C177 B.n137 VSUBS 0.009336f
C178 B.n138 VSUBS 0.009336f
C179 B.n139 VSUBS 0.009336f
C180 B.n140 VSUBS 0.009336f
C181 B.n141 VSUBS 0.009336f
C182 B.n142 VSUBS 0.009336f
C183 B.n143 VSUBS 0.009336f
C184 B.n144 VSUBS 0.009336f
C185 B.n145 VSUBS 0.009336f
C186 B.n146 VSUBS 0.009336f
C187 B.n147 VSUBS 0.009336f
C188 B.n148 VSUBS 0.009336f
C189 B.n149 VSUBS 0.009336f
C190 B.n150 VSUBS 0.006453f
C191 B.n151 VSUBS 0.021631f
C192 B.n152 VSUBS 0.007551f
C193 B.n153 VSUBS 0.009336f
C194 B.n154 VSUBS 0.009336f
C195 B.n155 VSUBS 0.009336f
C196 B.n156 VSUBS 0.009336f
C197 B.n157 VSUBS 0.009336f
C198 B.n158 VSUBS 0.009336f
C199 B.n159 VSUBS 0.009336f
C200 B.n160 VSUBS 0.009336f
C201 B.n161 VSUBS 0.009336f
C202 B.n162 VSUBS 0.009336f
C203 B.n163 VSUBS 0.009336f
C204 B.n164 VSUBS 0.007551f
C205 B.n165 VSUBS 0.009336f
C206 B.n166 VSUBS 0.009336f
C207 B.n167 VSUBS 0.006453f
C208 B.n168 VSUBS 0.009336f
C209 B.n169 VSUBS 0.009336f
C210 B.n170 VSUBS 0.009336f
C211 B.n171 VSUBS 0.009336f
C212 B.n172 VSUBS 0.009336f
C213 B.n173 VSUBS 0.009336f
C214 B.n174 VSUBS 0.009336f
C215 B.n175 VSUBS 0.009336f
C216 B.n176 VSUBS 0.009336f
C217 B.n177 VSUBS 0.009336f
C218 B.n178 VSUBS 0.009336f
C219 B.n179 VSUBS 0.009336f
C220 B.n180 VSUBS 0.009336f
C221 B.n181 VSUBS 0.023692f
C222 B.n182 VSUBS 0.023692f
C223 B.n183 VSUBS 0.022166f
C224 B.n184 VSUBS 0.009336f
C225 B.n185 VSUBS 0.009336f
C226 B.n186 VSUBS 0.009336f
C227 B.n187 VSUBS 0.009336f
C228 B.n188 VSUBS 0.009336f
C229 B.n189 VSUBS 0.009336f
C230 B.n190 VSUBS 0.009336f
C231 B.n191 VSUBS 0.009336f
C232 B.n192 VSUBS 0.009336f
C233 B.n193 VSUBS 0.009336f
C234 B.n194 VSUBS 0.009336f
C235 B.n195 VSUBS 0.009336f
C236 B.n196 VSUBS 0.009336f
C237 B.n197 VSUBS 0.009336f
C238 B.n198 VSUBS 0.009336f
C239 B.n199 VSUBS 0.009336f
C240 B.n200 VSUBS 0.009336f
C241 B.n201 VSUBS 0.009336f
C242 B.n202 VSUBS 0.009336f
C243 B.n203 VSUBS 0.009336f
C244 B.n204 VSUBS 0.009336f
C245 B.n205 VSUBS 0.009336f
C246 B.n206 VSUBS 0.009336f
C247 B.n207 VSUBS 0.009336f
C248 B.n208 VSUBS 0.009336f
C249 B.n209 VSUBS 0.009336f
C250 B.n210 VSUBS 0.009336f
C251 B.n211 VSUBS 0.009336f
C252 B.n212 VSUBS 0.009336f
C253 B.n213 VSUBS 0.009336f
C254 B.n214 VSUBS 0.009336f
C255 B.n215 VSUBS 0.009336f
C256 B.n216 VSUBS 0.009336f
C257 B.n217 VSUBS 0.009336f
C258 B.n218 VSUBS 0.009336f
C259 B.n219 VSUBS 0.009336f
C260 B.n220 VSUBS 0.009336f
C261 B.n221 VSUBS 0.009336f
C262 B.n222 VSUBS 0.009336f
C263 B.n223 VSUBS 0.009336f
C264 B.n224 VSUBS 0.009336f
C265 B.n225 VSUBS 0.009336f
C266 B.n226 VSUBS 0.009336f
C267 B.n227 VSUBS 0.009336f
C268 B.n228 VSUBS 0.009336f
C269 B.n229 VSUBS 0.009336f
C270 B.n230 VSUBS 0.009336f
C271 B.n231 VSUBS 0.009336f
C272 B.n232 VSUBS 0.009336f
C273 B.n233 VSUBS 0.009336f
C274 B.n234 VSUBS 0.009336f
C275 B.n235 VSUBS 0.009336f
C276 B.n236 VSUBS 0.009336f
C277 B.n237 VSUBS 0.009336f
C278 B.n238 VSUBS 0.009336f
C279 B.n239 VSUBS 0.009336f
C280 B.n240 VSUBS 0.009336f
C281 B.n241 VSUBS 0.009336f
C282 B.n242 VSUBS 0.009336f
C283 B.n243 VSUBS 0.009336f
C284 B.n244 VSUBS 0.009336f
C285 B.n245 VSUBS 0.009336f
C286 B.n246 VSUBS 0.009336f
C287 B.n247 VSUBS 0.009336f
C288 B.n248 VSUBS 0.009336f
C289 B.n249 VSUBS 0.009336f
C290 B.n250 VSUBS 0.009336f
C291 B.n251 VSUBS 0.009336f
C292 B.n252 VSUBS 0.009336f
C293 B.n253 VSUBS 0.009336f
C294 B.n254 VSUBS 0.009336f
C295 B.n255 VSUBS 0.009336f
C296 B.n256 VSUBS 0.009336f
C297 B.n257 VSUBS 0.009336f
C298 B.n258 VSUBS 0.009336f
C299 B.n259 VSUBS 0.009336f
C300 B.n260 VSUBS 0.009336f
C301 B.n261 VSUBS 0.009336f
C302 B.n262 VSUBS 0.009336f
C303 B.n263 VSUBS 0.009336f
C304 B.n264 VSUBS 0.023191f
C305 B.n265 VSUBS 0.022666f
C306 B.n266 VSUBS 0.023692f
C307 B.n267 VSUBS 0.009336f
C308 B.n268 VSUBS 0.009336f
C309 B.n269 VSUBS 0.009336f
C310 B.n270 VSUBS 0.009336f
C311 B.n271 VSUBS 0.009336f
C312 B.n272 VSUBS 0.009336f
C313 B.n273 VSUBS 0.009336f
C314 B.n274 VSUBS 0.009336f
C315 B.n275 VSUBS 0.009336f
C316 B.n276 VSUBS 0.009336f
C317 B.n277 VSUBS 0.009336f
C318 B.n278 VSUBS 0.009336f
C319 B.n279 VSUBS 0.009336f
C320 B.n280 VSUBS 0.009336f
C321 B.n281 VSUBS 0.006453f
C322 B.n282 VSUBS 0.021631f
C323 B.n283 VSUBS 0.007551f
C324 B.n284 VSUBS 0.009336f
C325 B.n285 VSUBS 0.009336f
C326 B.n286 VSUBS 0.009336f
C327 B.n287 VSUBS 0.009336f
C328 B.n288 VSUBS 0.009336f
C329 B.n289 VSUBS 0.009336f
C330 B.n290 VSUBS 0.009336f
C331 B.n291 VSUBS 0.009336f
C332 B.n292 VSUBS 0.009336f
C333 B.n293 VSUBS 0.009336f
C334 B.n294 VSUBS 0.009336f
C335 B.n295 VSUBS 0.007551f
C336 B.n296 VSUBS 0.021631f
C337 B.n297 VSUBS 0.006453f
C338 B.n298 VSUBS 0.009336f
C339 B.n299 VSUBS 0.009336f
C340 B.n300 VSUBS 0.009336f
C341 B.n301 VSUBS 0.009336f
C342 B.n302 VSUBS 0.009336f
C343 B.n303 VSUBS 0.009336f
C344 B.n304 VSUBS 0.009336f
C345 B.n305 VSUBS 0.009336f
C346 B.n306 VSUBS 0.009336f
C347 B.n307 VSUBS 0.009336f
C348 B.n308 VSUBS 0.009336f
C349 B.n309 VSUBS 0.009336f
C350 B.n310 VSUBS 0.009336f
C351 B.n311 VSUBS 0.009336f
C352 B.n312 VSUBS 0.023692f
C353 B.n313 VSUBS 0.023692f
C354 B.n314 VSUBS 0.022166f
C355 B.n315 VSUBS 0.009336f
C356 B.n316 VSUBS 0.009336f
C357 B.n317 VSUBS 0.009336f
C358 B.n318 VSUBS 0.009336f
C359 B.n319 VSUBS 0.009336f
C360 B.n320 VSUBS 0.009336f
C361 B.n321 VSUBS 0.009336f
C362 B.n322 VSUBS 0.009336f
C363 B.n323 VSUBS 0.009336f
C364 B.n324 VSUBS 0.009336f
C365 B.n325 VSUBS 0.009336f
C366 B.n326 VSUBS 0.009336f
C367 B.n327 VSUBS 0.009336f
C368 B.n328 VSUBS 0.009336f
C369 B.n329 VSUBS 0.009336f
C370 B.n330 VSUBS 0.009336f
C371 B.n331 VSUBS 0.009336f
C372 B.n332 VSUBS 0.009336f
C373 B.n333 VSUBS 0.009336f
C374 B.n334 VSUBS 0.009336f
C375 B.n335 VSUBS 0.009336f
C376 B.n336 VSUBS 0.009336f
C377 B.n337 VSUBS 0.009336f
C378 B.n338 VSUBS 0.009336f
C379 B.n339 VSUBS 0.009336f
C380 B.n340 VSUBS 0.009336f
C381 B.n341 VSUBS 0.009336f
C382 B.n342 VSUBS 0.009336f
C383 B.n343 VSUBS 0.009336f
C384 B.n344 VSUBS 0.009336f
C385 B.n345 VSUBS 0.009336f
C386 B.n346 VSUBS 0.009336f
C387 B.n347 VSUBS 0.009336f
C388 B.n348 VSUBS 0.009336f
C389 B.n349 VSUBS 0.009336f
C390 B.n350 VSUBS 0.009336f
C391 B.n351 VSUBS 0.009336f
C392 B.n352 VSUBS 0.009336f
C393 B.n353 VSUBS 0.009336f
C394 B.n354 VSUBS 0.009336f
C395 B.n355 VSUBS 0.02114f
C396 VDD2.t4 VSUBS 0.124039f
C397 VDD2.t2 VSUBS 0.020204f
C398 VDD2.t0 VSUBS 0.020204f
C399 VDD2.n0 VSUBS 0.077431f
C400 VDD2.n1 VSUBS 1.19613f
C401 VDD2.t1 VSUBS 0.123196f
C402 VDD2.n2 VSUBS 1.08248f
C403 VDD2.t5 VSUBS 0.020204f
C404 VDD2.t3 VSUBS 0.020204f
C405 VDD2.n3 VSUBS 0.077426f
C406 VN.n0 VSUBS 0.068812f
C407 VN.t3 VSUBS 0.215431f
C408 VN.n1 VSUBS 0.208939f
C409 VN.t1 VSUBS 0.384077f
C410 VN.n2 VSUBS 0.231941f
C411 VN.n3 VSUBS 0.27316f
C412 VN.n4 VSUBS 0.080923f
C413 VN.n5 VSUBS 0.035321f
C414 VN.t5 VSUBS 0.318763f
C415 VN.n6 VSUBS 0.247083f
C416 VN.n7 VSUBS 0.048296f
C417 VN.n8 VSUBS 0.068812f
C418 VN.t0 VSUBS 0.215431f
C419 VN.n9 VSUBS 0.208939f
C420 VN.t2 VSUBS 0.384077f
C421 VN.n10 VSUBS 0.231941f
C422 VN.n11 VSUBS 0.27316f
C423 VN.n12 VSUBS 0.080923f
C424 VN.n13 VSUBS 0.035321f
C425 VN.t4 VSUBS 0.318763f
C426 VN.n14 VSUBS 0.247083f
C427 VN.n15 VSUBS 1.65331f
C428 VTAIL.t2 VSUBS 0.026866f
C429 VTAIL.t4 VSUBS 0.026866f
C430 VTAIL.n0 VSUBS 0.087777f
C431 VTAIL.n1 VSUBS 0.312171f
C432 VTAIL.t7 VSUBS 0.149528f
C433 VTAIL.n2 VSUBS 0.397389f
C434 VTAIL.t10 VSUBS 0.026866f
C435 VTAIL.t6 VSUBS 0.026866f
C436 VTAIL.n3 VSUBS 0.087777f
C437 VTAIL.n4 VSUBS 0.913579f
C438 VTAIL.t3 VSUBS 0.026866f
C439 VTAIL.t5 VSUBS 0.026866f
C440 VTAIL.n5 VSUBS 0.087777f
C441 VTAIL.n6 VSUBS 0.913579f
C442 VTAIL.t0 VSUBS 0.149528f
C443 VTAIL.n7 VSUBS 0.397389f
C444 VTAIL.t9 VSUBS 0.026866f
C445 VTAIL.t11 VSUBS 0.026866f
C446 VTAIL.n8 VSUBS 0.087777f
C447 VTAIL.n9 VSUBS 0.38587f
C448 VTAIL.t8 VSUBS 0.149528f
C449 VTAIL.n10 VSUBS 0.821089f
C450 VTAIL.t1 VSUBS 0.149528f
C451 VTAIL.n11 VSUBS 0.79078f
C452 VDD1.t0 VSUBS 0.121655f
C453 VDD1.t5 VSUBS 0.121538f
C454 VDD1.t4 VSUBS 0.019797f
C455 VDD1.t2 VSUBS 0.019797f
C456 VDD1.n0 VSUBS 0.075869f
C457 VDD1.n1 VSUBS 1.2285f
C458 VDD1.t3 VSUBS 0.019797f
C459 VDD1.t1 VSUBS 0.019797f
C460 VDD1.n2 VSUBS 0.075566f
C461 VDD1.n3 VSUBS 1.08979f
C462 VP.n0 VSUBS 0.072263f
C463 VP.t5 VSUBS 0.226235f
C464 VP.n1 VSUBS 0.147417f
C465 VP.n2 VSUBS 0.072263f
C466 VP.n3 VSUBS 0.072263f
C467 VP.t3 VSUBS 0.334749f
C468 VP.t0 VSUBS 0.226235f
C469 VP.n4 VSUBS 0.219417f
C470 VP.t2 VSUBS 0.403339f
C471 VP.n5 VSUBS 0.243572f
C472 VP.n6 VSUBS 0.286859f
C473 VP.n7 VSUBS 0.084981f
C474 VP.n8 VSUBS 0.037092f
C475 VP.n9 VSUBS 0.259474f
C476 VP.n10 VSUBS 1.70491f
C477 VP.n11 VSUBS 1.75912f
C478 VP.t1 VSUBS 0.334749f
C479 VP.n12 VSUBS 0.259474f
C480 VP.n13 VSUBS 0.037092f
C481 VP.n14 VSUBS 0.084981f
C482 VP.n15 VSUBS 0.054155f
C483 VP.n16 VSUBS 0.054155f
C484 VP.n17 VSUBS 0.084981f
C485 VP.n18 VSUBS 0.037092f
C486 VP.t4 VSUBS 0.334749f
C487 VP.n19 VSUBS 0.259474f
C488 VP.n20 VSUBS 0.050718f
.ends

