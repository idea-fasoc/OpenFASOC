* NGSPICE file created from diff_pair_sample_1253.ext - technology: sky130A

.subckt diff_pair_sample_1253 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t13 w_n1510_n2050# sky130_fd_pr__pfet_01v8 ad=0.89265 pd=5.74 as=2.1099 ps=11.6 w=5.41 l=0.21
X1 B.t11 B.t9 B.t10 w_n1510_n2050# sky130_fd_pr__pfet_01v8 ad=2.1099 pd=11.6 as=0 ps=0 w=5.41 l=0.21
X2 VTAIL.t2 VP.t0 VDD1.t7 w_n1510_n2050# sky130_fd_pr__pfet_01v8 ad=0.89265 pd=5.74 as=0.89265 ps=5.74 w=5.41 l=0.21
X3 VDD1.t6 VP.t1 VTAIL.t4 w_n1510_n2050# sky130_fd_pr__pfet_01v8 ad=0.89265 pd=5.74 as=2.1099 ps=11.6 w=5.41 l=0.21
X4 B.t8 B.t6 B.t7 w_n1510_n2050# sky130_fd_pr__pfet_01v8 ad=2.1099 pd=11.6 as=0 ps=0 w=5.41 l=0.21
X5 B.t5 B.t3 B.t4 w_n1510_n2050# sky130_fd_pr__pfet_01v8 ad=2.1099 pd=11.6 as=0 ps=0 w=5.41 l=0.21
X6 VDD2.t6 VN.t1 VTAIL.t15 w_n1510_n2050# sky130_fd_pr__pfet_01v8 ad=0.89265 pd=5.74 as=2.1099 ps=11.6 w=5.41 l=0.21
X7 VTAIL.t14 VN.t2 VDD2.t5 w_n1510_n2050# sky130_fd_pr__pfet_01v8 ad=0.89265 pd=5.74 as=0.89265 ps=5.74 w=5.41 l=0.21
X8 VTAIL.t12 VN.t3 VDD2.t4 w_n1510_n2050# sky130_fd_pr__pfet_01v8 ad=0.89265 pd=5.74 as=0.89265 ps=5.74 w=5.41 l=0.21
X9 VDD2.t3 VN.t4 VTAIL.t10 w_n1510_n2050# sky130_fd_pr__pfet_01v8 ad=0.89265 pd=5.74 as=0.89265 ps=5.74 w=5.41 l=0.21
X10 VTAIL.t9 VN.t5 VDD2.t2 w_n1510_n2050# sky130_fd_pr__pfet_01v8 ad=2.1099 pd=11.6 as=0.89265 ps=5.74 w=5.41 l=0.21
X11 VTAIL.t1 VP.t2 VDD1.t5 w_n1510_n2050# sky130_fd_pr__pfet_01v8 ad=2.1099 pd=11.6 as=0.89265 ps=5.74 w=5.41 l=0.21
X12 VDD1.t4 VP.t3 VTAIL.t7 w_n1510_n2050# sky130_fd_pr__pfet_01v8 ad=0.89265 pd=5.74 as=0.89265 ps=5.74 w=5.41 l=0.21
X13 VDD1.t3 VP.t4 VTAIL.t3 w_n1510_n2050# sky130_fd_pr__pfet_01v8 ad=0.89265 pd=5.74 as=0.89265 ps=5.74 w=5.41 l=0.21
X14 VTAIL.t8 VN.t6 VDD2.t1 w_n1510_n2050# sky130_fd_pr__pfet_01v8 ad=2.1099 pd=11.6 as=0.89265 ps=5.74 w=5.41 l=0.21
X15 B.t2 B.t0 B.t1 w_n1510_n2050# sky130_fd_pr__pfet_01v8 ad=2.1099 pd=11.6 as=0 ps=0 w=5.41 l=0.21
X16 VTAIL.t0 VP.t5 VDD1.t2 w_n1510_n2050# sky130_fd_pr__pfet_01v8 ad=0.89265 pd=5.74 as=0.89265 ps=5.74 w=5.41 l=0.21
X17 VDD2.t0 VN.t7 VTAIL.t11 w_n1510_n2050# sky130_fd_pr__pfet_01v8 ad=0.89265 pd=5.74 as=0.89265 ps=5.74 w=5.41 l=0.21
X18 VDD1.t1 VP.t6 VTAIL.t5 w_n1510_n2050# sky130_fd_pr__pfet_01v8 ad=0.89265 pd=5.74 as=2.1099 ps=11.6 w=5.41 l=0.21
X19 VTAIL.t6 VP.t7 VDD1.t0 w_n1510_n2050# sky130_fd_pr__pfet_01v8 ad=2.1099 pd=11.6 as=0.89265 ps=5.74 w=5.41 l=0.21
R0 VN.n5 VN.t0 816.48
R1 VN.n1 VN.t5 816.48
R2 VN.n12 VN.t6 816.48
R3 VN.n8 VN.t1 816.48
R4 VN.n4 VN.t2 771.201
R5 VN.n2 VN.t7 771.201
R6 VN.n11 VN.t4 771.201
R7 VN.n9 VN.t3 771.201
R8 VN.n8 VN.n7 161.489
R9 VN.n1 VN.n0 161.489
R10 VN.n6 VN.n5 161.3
R11 VN.n13 VN.n12 161.3
R12 VN.n10 VN.n7 161.3
R13 VN.n3 VN.n0 161.3
R14 VN.n3 VN.n2 39.4369
R15 VN.n4 VN.n3 39.4369
R16 VN.n11 VN.n10 39.4369
R17 VN.n10 VN.n9 39.4369
R18 VN VN.n13 35.1691
R19 VN.n2 VN.n1 33.5944
R20 VN.n5 VN.n4 33.5944
R21 VN.n12 VN.n11 33.5944
R22 VN.n9 VN.n8 33.5944
R23 VN.n13 VN.n7 0.189894
R24 VN.n6 VN.n0 0.189894
R25 VN VN.n6 0.0516364
R26 VTAIL.n226 VTAIL.n204 756.745
R27 VTAIL.n24 VTAIL.n2 756.745
R28 VTAIL.n52 VTAIL.n30 756.745
R29 VTAIL.n82 VTAIL.n60 756.745
R30 VTAIL.n198 VTAIL.n176 756.745
R31 VTAIL.n168 VTAIL.n146 756.745
R32 VTAIL.n140 VTAIL.n118 756.745
R33 VTAIL.n110 VTAIL.n88 756.745
R34 VTAIL.n212 VTAIL.n211 585
R35 VTAIL.n217 VTAIL.n216 585
R36 VTAIL.n219 VTAIL.n218 585
R37 VTAIL.n208 VTAIL.n207 585
R38 VTAIL.n225 VTAIL.n224 585
R39 VTAIL.n227 VTAIL.n226 585
R40 VTAIL.n10 VTAIL.n9 585
R41 VTAIL.n15 VTAIL.n14 585
R42 VTAIL.n17 VTAIL.n16 585
R43 VTAIL.n6 VTAIL.n5 585
R44 VTAIL.n23 VTAIL.n22 585
R45 VTAIL.n25 VTAIL.n24 585
R46 VTAIL.n38 VTAIL.n37 585
R47 VTAIL.n43 VTAIL.n42 585
R48 VTAIL.n45 VTAIL.n44 585
R49 VTAIL.n34 VTAIL.n33 585
R50 VTAIL.n51 VTAIL.n50 585
R51 VTAIL.n53 VTAIL.n52 585
R52 VTAIL.n68 VTAIL.n67 585
R53 VTAIL.n73 VTAIL.n72 585
R54 VTAIL.n75 VTAIL.n74 585
R55 VTAIL.n64 VTAIL.n63 585
R56 VTAIL.n81 VTAIL.n80 585
R57 VTAIL.n83 VTAIL.n82 585
R58 VTAIL.n199 VTAIL.n198 585
R59 VTAIL.n197 VTAIL.n196 585
R60 VTAIL.n180 VTAIL.n179 585
R61 VTAIL.n191 VTAIL.n190 585
R62 VTAIL.n189 VTAIL.n188 585
R63 VTAIL.n184 VTAIL.n183 585
R64 VTAIL.n169 VTAIL.n168 585
R65 VTAIL.n167 VTAIL.n166 585
R66 VTAIL.n150 VTAIL.n149 585
R67 VTAIL.n161 VTAIL.n160 585
R68 VTAIL.n159 VTAIL.n158 585
R69 VTAIL.n154 VTAIL.n153 585
R70 VTAIL.n141 VTAIL.n140 585
R71 VTAIL.n139 VTAIL.n138 585
R72 VTAIL.n122 VTAIL.n121 585
R73 VTAIL.n133 VTAIL.n132 585
R74 VTAIL.n131 VTAIL.n130 585
R75 VTAIL.n126 VTAIL.n125 585
R76 VTAIL.n111 VTAIL.n110 585
R77 VTAIL.n109 VTAIL.n108 585
R78 VTAIL.n92 VTAIL.n91 585
R79 VTAIL.n103 VTAIL.n102 585
R80 VTAIL.n101 VTAIL.n100 585
R81 VTAIL.n96 VTAIL.n95 585
R82 VTAIL.n213 VTAIL.t13 327.856
R83 VTAIL.n11 VTAIL.t9 327.856
R84 VTAIL.n39 VTAIL.t5 327.856
R85 VTAIL.n69 VTAIL.t6 327.856
R86 VTAIL.n185 VTAIL.t4 327.856
R87 VTAIL.n155 VTAIL.t1 327.856
R88 VTAIL.n127 VTAIL.t15 327.856
R89 VTAIL.n97 VTAIL.t8 327.856
R90 VTAIL.n217 VTAIL.n211 171.744
R91 VTAIL.n218 VTAIL.n217 171.744
R92 VTAIL.n218 VTAIL.n207 171.744
R93 VTAIL.n225 VTAIL.n207 171.744
R94 VTAIL.n226 VTAIL.n225 171.744
R95 VTAIL.n15 VTAIL.n9 171.744
R96 VTAIL.n16 VTAIL.n15 171.744
R97 VTAIL.n16 VTAIL.n5 171.744
R98 VTAIL.n23 VTAIL.n5 171.744
R99 VTAIL.n24 VTAIL.n23 171.744
R100 VTAIL.n43 VTAIL.n37 171.744
R101 VTAIL.n44 VTAIL.n43 171.744
R102 VTAIL.n44 VTAIL.n33 171.744
R103 VTAIL.n51 VTAIL.n33 171.744
R104 VTAIL.n52 VTAIL.n51 171.744
R105 VTAIL.n73 VTAIL.n67 171.744
R106 VTAIL.n74 VTAIL.n73 171.744
R107 VTAIL.n74 VTAIL.n63 171.744
R108 VTAIL.n81 VTAIL.n63 171.744
R109 VTAIL.n82 VTAIL.n81 171.744
R110 VTAIL.n198 VTAIL.n197 171.744
R111 VTAIL.n197 VTAIL.n179 171.744
R112 VTAIL.n190 VTAIL.n179 171.744
R113 VTAIL.n190 VTAIL.n189 171.744
R114 VTAIL.n189 VTAIL.n183 171.744
R115 VTAIL.n168 VTAIL.n167 171.744
R116 VTAIL.n167 VTAIL.n149 171.744
R117 VTAIL.n160 VTAIL.n149 171.744
R118 VTAIL.n160 VTAIL.n159 171.744
R119 VTAIL.n159 VTAIL.n153 171.744
R120 VTAIL.n140 VTAIL.n139 171.744
R121 VTAIL.n139 VTAIL.n121 171.744
R122 VTAIL.n132 VTAIL.n121 171.744
R123 VTAIL.n132 VTAIL.n131 171.744
R124 VTAIL.n131 VTAIL.n125 171.744
R125 VTAIL.n110 VTAIL.n109 171.744
R126 VTAIL.n109 VTAIL.n91 171.744
R127 VTAIL.n102 VTAIL.n91 171.744
R128 VTAIL.n102 VTAIL.n101 171.744
R129 VTAIL.n101 VTAIL.n95 171.744
R130 VTAIL.t13 VTAIL.n211 85.8723
R131 VTAIL.t9 VTAIL.n9 85.8723
R132 VTAIL.t5 VTAIL.n37 85.8723
R133 VTAIL.t6 VTAIL.n67 85.8723
R134 VTAIL.t4 VTAIL.n183 85.8723
R135 VTAIL.t1 VTAIL.n153 85.8723
R136 VTAIL.t15 VTAIL.n125 85.8723
R137 VTAIL.t8 VTAIL.n95 85.8723
R138 VTAIL.n175 VTAIL.n174 83.1733
R139 VTAIL.n117 VTAIL.n116 83.1733
R140 VTAIL.n1 VTAIL.n0 83.1732
R141 VTAIL.n59 VTAIL.n58 83.1732
R142 VTAIL.n231 VTAIL.n230 34.7066
R143 VTAIL.n29 VTAIL.n28 34.7066
R144 VTAIL.n57 VTAIL.n56 34.7066
R145 VTAIL.n87 VTAIL.n86 34.7066
R146 VTAIL.n203 VTAIL.n202 34.7066
R147 VTAIL.n173 VTAIL.n172 34.7066
R148 VTAIL.n145 VTAIL.n144 34.7066
R149 VTAIL.n115 VTAIL.n114 34.7066
R150 VTAIL.n231 VTAIL.n203 17.4962
R151 VTAIL.n115 VTAIL.n87 17.4962
R152 VTAIL.n213 VTAIL.n212 16.381
R153 VTAIL.n11 VTAIL.n10 16.381
R154 VTAIL.n39 VTAIL.n38 16.381
R155 VTAIL.n69 VTAIL.n68 16.381
R156 VTAIL.n185 VTAIL.n184 16.381
R157 VTAIL.n155 VTAIL.n154 16.381
R158 VTAIL.n127 VTAIL.n126 16.381
R159 VTAIL.n97 VTAIL.n96 16.381
R160 VTAIL.n216 VTAIL.n215 12.8005
R161 VTAIL.n14 VTAIL.n13 12.8005
R162 VTAIL.n42 VTAIL.n41 12.8005
R163 VTAIL.n72 VTAIL.n71 12.8005
R164 VTAIL.n188 VTAIL.n187 12.8005
R165 VTAIL.n158 VTAIL.n157 12.8005
R166 VTAIL.n130 VTAIL.n129 12.8005
R167 VTAIL.n100 VTAIL.n99 12.8005
R168 VTAIL.n219 VTAIL.n210 12.0247
R169 VTAIL.n17 VTAIL.n8 12.0247
R170 VTAIL.n45 VTAIL.n36 12.0247
R171 VTAIL.n75 VTAIL.n66 12.0247
R172 VTAIL.n191 VTAIL.n182 12.0247
R173 VTAIL.n161 VTAIL.n152 12.0247
R174 VTAIL.n133 VTAIL.n124 12.0247
R175 VTAIL.n103 VTAIL.n94 12.0247
R176 VTAIL.n220 VTAIL.n208 11.249
R177 VTAIL.n18 VTAIL.n6 11.249
R178 VTAIL.n46 VTAIL.n34 11.249
R179 VTAIL.n76 VTAIL.n64 11.249
R180 VTAIL.n192 VTAIL.n180 11.249
R181 VTAIL.n162 VTAIL.n150 11.249
R182 VTAIL.n134 VTAIL.n122 11.249
R183 VTAIL.n104 VTAIL.n92 11.249
R184 VTAIL.n224 VTAIL.n223 10.4732
R185 VTAIL.n22 VTAIL.n21 10.4732
R186 VTAIL.n50 VTAIL.n49 10.4732
R187 VTAIL.n80 VTAIL.n79 10.4732
R188 VTAIL.n196 VTAIL.n195 10.4732
R189 VTAIL.n166 VTAIL.n165 10.4732
R190 VTAIL.n138 VTAIL.n137 10.4732
R191 VTAIL.n108 VTAIL.n107 10.4732
R192 VTAIL.n227 VTAIL.n206 9.69747
R193 VTAIL.n25 VTAIL.n4 9.69747
R194 VTAIL.n53 VTAIL.n32 9.69747
R195 VTAIL.n83 VTAIL.n62 9.69747
R196 VTAIL.n199 VTAIL.n178 9.69747
R197 VTAIL.n169 VTAIL.n148 9.69747
R198 VTAIL.n141 VTAIL.n120 9.69747
R199 VTAIL.n111 VTAIL.n90 9.69747
R200 VTAIL.n230 VTAIL.n229 9.45567
R201 VTAIL.n28 VTAIL.n27 9.45567
R202 VTAIL.n56 VTAIL.n55 9.45567
R203 VTAIL.n86 VTAIL.n85 9.45567
R204 VTAIL.n202 VTAIL.n201 9.45567
R205 VTAIL.n172 VTAIL.n171 9.45567
R206 VTAIL.n144 VTAIL.n143 9.45567
R207 VTAIL.n114 VTAIL.n113 9.45567
R208 VTAIL.n229 VTAIL.n228 9.3005
R209 VTAIL.n206 VTAIL.n205 9.3005
R210 VTAIL.n223 VTAIL.n222 9.3005
R211 VTAIL.n221 VTAIL.n220 9.3005
R212 VTAIL.n210 VTAIL.n209 9.3005
R213 VTAIL.n215 VTAIL.n214 9.3005
R214 VTAIL.n27 VTAIL.n26 9.3005
R215 VTAIL.n4 VTAIL.n3 9.3005
R216 VTAIL.n21 VTAIL.n20 9.3005
R217 VTAIL.n19 VTAIL.n18 9.3005
R218 VTAIL.n8 VTAIL.n7 9.3005
R219 VTAIL.n13 VTAIL.n12 9.3005
R220 VTAIL.n55 VTAIL.n54 9.3005
R221 VTAIL.n32 VTAIL.n31 9.3005
R222 VTAIL.n49 VTAIL.n48 9.3005
R223 VTAIL.n47 VTAIL.n46 9.3005
R224 VTAIL.n36 VTAIL.n35 9.3005
R225 VTAIL.n41 VTAIL.n40 9.3005
R226 VTAIL.n85 VTAIL.n84 9.3005
R227 VTAIL.n62 VTAIL.n61 9.3005
R228 VTAIL.n79 VTAIL.n78 9.3005
R229 VTAIL.n77 VTAIL.n76 9.3005
R230 VTAIL.n66 VTAIL.n65 9.3005
R231 VTAIL.n71 VTAIL.n70 9.3005
R232 VTAIL.n201 VTAIL.n200 9.3005
R233 VTAIL.n178 VTAIL.n177 9.3005
R234 VTAIL.n195 VTAIL.n194 9.3005
R235 VTAIL.n193 VTAIL.n192 9.3005
R236 VTAIL.n182 VTAIL.n181 9.3005
R237 VTAIL.n187 VTAIL.n186 9.3005
R238 VTAIL.n171 VTAIL.n170 9.3005
R239 VTAIL.n148 VTAIL.n147 9.3005
R240 VTAIL.n165 VTAIL.n164 9.3005
R241 VTAIL.n163 VTAIL.n162 9.3005
R242 VTAIL.n152 VTAIL.n151 9.3005
R243 VTAIL.n157 VTAIL.n156 9.3005
R244 VTAIL.n143 VTAIL.n142 9.3005
R245 VTAIL.n120 VTAIL.n119 9.3005
R246 VTAIL.n137 VTAIL.n136 9.3005
R247 VTAIL.n135 VTAIL.n134 9.3005
R248 VTAIL.n124 VTAIL.n123 9.3005
R249 VTAIL.n129 VTAIL.n128 9.3005
R250 VTAIL.n113 VTAIL.n112 9.3005
R251 VTAIL.n90 VTAIL.n89 9.3005
R252 VTAIL.n107 VTAIL.n106 9.3005
R253 VTAIL.n105 VTAIL.n104 9.3005
R254 VTAIL.n94 VTAIL.n93 9.3005
R255 VTAIL.n99 VTAIL.n98 9.3005
R256 VTAIL.n228 VTAIL.n204 8.92171
R257 VTAIL.n26 VTAIL.n2 8.92171
R258 VTAIL.n54 VTAIL.n30 8.92171
R259 VTAIL.n84 VTAIL.n60 8.92171
R260 VTAIL.n200 VTAIL.n176 8.92171
R261 VTAIL.n170 VTAIL.n146 8.92171
R262 VTAIL.n142 VTAIL.n118 8.92171
R263 VTAIL.n112 VTAIL.n88 8.92171
R264 VTAIL.n0 VTAIL.t11 6.00882
R265 VTAIL.n0 VTAIL.t14 6.00882
R266 VTAIL.n58 VTAIL.t7 6.00882
R267 VTAIL.n58 VTAIL.t2 6.00882
R268 VTAIL.n174 VTAIL.t3 6.00882
R269 VTAIL.n174 VTAIL.t0 6.00882
R270 VTAIL.n116 VTAIL.t10 6.00882
R271 VTAIL.n116 VTAIL.t12 6.00882
R272 VTAIL.n230 VTAIL.n204 5.04292
R273 VTAIL.n28 VTAIL.n2 5.04292
R274 VTAIL.n56 VTAIL.n30 5.04292
R275 VTAIL.n86 VTAIL.n60 5.04292
R276 VTAIL.n202 VTAIL.n176 5.04292
R277 VTAIL.n172 VTAIL.n146 5.04292
R278 VTAIL.n144 VTAIL.n118 5.04292
R279 VTAIL.n114 VTAIL.n88 5.04292
R280 VTAIL.n228 VTAIL.n227 4.26717
R281 VTAIL.n26 VTAIL.n25 4.26717
R282 VTAIL.n54 VTAIL.n53 4.26717
R283 VTAIL.n84 VTAIL.n83 4.26717
R284 VTAIL.n200 VTAIL.n199 4.26717
R285 VTAIL.n170 VTAIL.n169 4.26717
R286 VTAIL.n142 VTAIL.n141 4.26717
R287 VTAIL.n112 VTAIL.n111 4.26717
R288 VTAIL.n186 VTAIL.n185 3.71853
R289 VTAIL.n156 VTAIL.n155 3.71853
R290 VTAIL.n128 VTAIL.n127 3.71853
R291 VTAIL.n98 VTAIL.n97 3.71853
R292 VTAIL.n214 VTAIL.n213 3.71853
R293 VTAIL.n12 VTAIL.n11 3.71853
R294 VTAIL.n40 VTAIL.n39 3.71853
R295 VTAIL.n70 VTAIL.n69 3.71853
R296 VTAIL.n224 VTAIL.n206 3.49141
R297 VTAIL.n22 VTAIL.n4 3.49141
R298 VTAIL.n50 VTAIL.n32 3.49141
R299 VTAIL.n80 VTAIL.n62 3.49141
R300 VTAIL.n196 VTAIL.n178 3.49141
R301 VTAIL.n166 VTAIL.n148 3.49141
R302 VTAIL.n138 VTAIL.n120 3.49141
R303 VTAIL.n108 VTAIL.n90 3.49141
R304 VTAIL.n223 VTAIL.n208 2.71565
R305 VTAIL.n21 VTAIL.n6 2.71565
R306 VTAIL.n49 VTAIL.n34 2.71565
R307 VTAIL.n79 VTAIL.n64 2.71565
R308 VTAIL.n195 VTAIL.n180 2.71565
R309 VTAIL.n165 VTAIL.n150 2.71565
R310 VTAIL.n137 VTAIL.n122 2.71565
R311 VTAIL.n107 VTAIL.n92 2.71565
R312 VTAIL.n220 VTAIL.n219 1.93989
R313 VTAIL.n18 VTAIL.n17 1.93989
R314 VTAIL.n46 VTAIL.n45 1.93989
R315 VTAIL.n76 VTAIL.n75 1.93989
R316 VTAIL.n192 VTAIL.n191 1.93989
R317 VTAIL.n162 VTAIL.n161 1.93989
R318 VTAIL.n134 VTAIL.n133 1.93989
R319 VTAIL.n104 VTAIL.n103 1.93989
R320 VTAIL.n216 VTAIL.n210 1.16414
R321 VTAIL.n14 VTAIL.n8 1.16414
R322 VTAIL.n42 VTAIL.n36 1.16414
R323 VTAIL.n72 VTAIL.n66 1.16414
R324 VTAIL.n188 VTAIL.n182 1.16414
R325 VTAIL.n158 VTAIL.n152 1.16414
R326 VTAIL.n130 VTAIL.n124 1.16414
R327 VTAIL.n100 VTAIL.n94 1.16414
R328 VTAIL.n173 VTAIL.n145 0.470328
R329 VTAIL.n57 VTAIL.n29 0.470328
R330 VTAIL.n117 VTAIL.n115 0.466017
R331 VTAIL.n145 VTAIL.n117 0.466017
R332 VTAIL.n175 VTAIL.n173 0.466017
R333 VTAIL.n203 VTAIL.n175 0.466017
R334 VTAIL.n87 VTAIL.n59 0.466017
R335 VTAIL.n59 VTAIL.n57 0.466017
R336 VTAIL.n29 VTAIL.n1 0.466017
R337 VTAIL VTAIL.n231 0.407828
R338 VTAIL.n215 VTAIL.n212 0.388379
R339 VTAIL.n13 VTAIL.n10 0.388379
R340 VTAIL.n41 VTAIL.n38 0.388379
R341 VTAIL.n71 VTAIL.n68 0.388379
R342 VTAIL.n187 VTAIL.n184 0.388379
R343 VTAIL.n157 VTAIL.n154 0.388379
R344 VTAIL.n129 VTAIL.n126 0.388379
R345 VTAIL.n99 VTAIL.n96 0.388379
R346 VTAIL.n214 VTAIL.n209 0.155672
R347 VTAIL.n221 VTAIL.n209 0.155672
R348 VTAIL.n222 VTAIL.n221 0.155672
R349 VTAIL.n222 VTAIL.n205 0.155672
R350 VTAIL.n229 VTAIL.n205 0.155672
R351 VTAIL.n12 VTAIL.n7 0.155672
R352 VTAIL.n19 VTAIL.n7 0.155672
R353 VTAIL.n20 VTAIL.n19 0.155672
R354 VTAIL.n20 VTAIL.n3 0.155672
R355 VTAIL.n27 VTAIL.n3 0.155672
R356 VTAIL.n40 VTAIL.n35 0.155672
R357 VTAIL.n47 VTAIL.n35 0.155672
R358 VTAIL.n48 VTAIL.n47 0.155672
R359 VTAIL.n48 VTAIL.n31 0.155672
R360 VTAIL.n55 VTAIL.n31 0.155672
R361 VTAIL.n70 VTAIL.n65 0.155672
R362 VTAIL.n77 VTAIL.n65 0.155672
R363 VTAIL.n78 VTAIL.n77 0.155672
R364 VTAIL.n78 VTAIL.n61 0.155672
R365 VTAIL.n85 VTAIL.n61 0.155672
R366 VTAIL.n201 VTAIL.n177 0.155672
R367 VTAIL.n194 VTAIL.n177 0.155672
R368 VTAIL.n194 VTAIL.n193 0.155672
R369 VTAIL.n193 VTAIL.n181 0.155672
R370 VTAIL.n186 VTAIL.n181 0.155672
R371 VTAIL.n171 VTAIL.n147 0.155672
R372 VTAIL.n164 VTAIL.n147 0.155672
R373 VTAIL.n164 VTAIL.n163 0.155672
R374 VTAIL.n163 VTAIL.n151 0.155672
R375 VTAIL.n156 VTAIL.n151 0.155672
R376 VTAIL.n143 VTAIL.n119 0.155672
R377 VTAIL.n136 VTAIL.n119 0.155672
R378 VTAIL.n136 VTAIL.n135 0.155672
R379 VTAIL.n135 VTAIL.n123 0.155672
R380 VTAIL.n128 VTAIL.n123 0.155672
R381 VTAIL.n113 VTAIL.n89 0.155672
R382 VTAIL.n106 VTAIL.n89 0.155672
R383 VTAIL.n106 VTAIL.n105 0.155672
R384 VTAIL.n105 VTAIL.n93 0.155672
R385 VTAIL.n98 VTAIL.n93 0.155672
R386 VTAIL VTAIL.n1 0.0586897
R387 VDD2.n2 VDD2.n1 100.029
R388 VDD2.n2 VDD2.n0 100.029
R389 VDD2 VDD2.n5 100.026
R390 VDD2.n4 VDD2.n3 99.8521
R391 VDD2.n4 VDD2.n2 30.4739
R392 VDD2.n5 VDD2.t4 6.00882
R393 VDD2.n5 VDD2.t6 6.00882
R394 VDD2.n3 VDD2.t1 6.00882
R395 VDD2.n3 VDD2.t3 6.00882
R396 VDD2.n1 VDD2.t5 6.00882
R397 VDD2.n1 VDD2.t7 6.00882
R398 VDD2.n0 VDD2.t2 6.00882
R399 VDD2.n0 VDD2.t0 6.00882
R400 VDD2 VDD2.n4 0.291448
R401 B.n70 B.t9 854.343
R402 B.n76 B.t3 854.343
R403 B.n22 B.t0 854.343
R404 B.n28 B.t6 854.343
R405 B.n252 B.n41 585
R406 B.n254 B.n253 585
R407 B.n255 B.n40 585
R408 B.n257 B.n256 585
R409 B.n258 B.n39 585
R410 B.n260 B.n259 585
R411 B.n261 B.n38 585
R412 B.n263 B.n262 585
R413 B.n264 B.n37 585
R414 B.n266 B.n265 585
R415 B.n267 B.n36 585
R416 B.n269 B.n268 585
R417 B.n270 B.n35 585
R418 B.n272 B.n271 585
R419 B.n273 B.n34 585
R420 B.n275 B.n274 585
R421 B.n276 B.n33 585
R422 B.n278 B.n277 585
R423 B.n279 B.n32 585
R424 B.n281 B.n280 585
R425 B.n282 B.n31 585
R426 B.n284 B.n283 585
R427 B.n286 B.n285 585
R428 B.n287 B.n27 585
R429 B.n289 B.n288 585
R430 B.n290 B.n26 585
R431 B.n292 B.n291 585
R432 B.n293 B.n25 585
R433 B.n295 B.n294 585
R434 B.n296 B.n24 585
R435 B.n298 B.n297 585
R436 B.n299 B.n21 585
R437 B.n302 B.n301 585
R438 B.n303 B.n20 585
R439 B.n305 B.n304 585
R440 B.n306 B.n19 585
R441 B.n308 B.n307 585
R442 B.n309 B.n18 585
R443 B.n311 B.n310 585
R444 B.n312 B.n17 585
R445 B.n314 B.n313 585
R446 B.n315 B.n16 585
R447 B.n317 B.n316 585
R448 B.n318 B.n15 585
R449 B.n320 B.n319 585
R450 B.n321 B.n14 585
R451 B.n323 B.n322 585
R452 B.n324 B.n13 585
R453 B.n326 B.n325 585
R454 B.n327 B.n12 585
R455 B.n329 B.n328 585
R456 B.n330 B.n11 585
R457 B.n332 B.n331 585
R458 B.n333 B.n10 585
R459 B.n251 B.n250 585
R460 B.n249 B.n42 585
R461 B.n248 B.n247 585
R462 B.n246 B.n43 585
R463 B.n245 B.n244 585
R464 B.n243 B.n44 585
R465 B.n242 B.n241 585
R466 B.n240 B.n45 585
R467 B.n239 B.n238 585
R468 B.n237 B.n46 585
R469 B.n236 B.n235 585
R470 B.n234 B.n47 585
R471 B.n233 B.n232 585
R472 B.n231 B.n48 585
R473 B.n230 B.n229 585
R474 B.n228 B.n49 585
R475 B.n227 B.n226 585
R476 B.n225 B.n50 585
R477 B.n224 B.n223 585
R478 B.n222 B.n51 585
R479 B.n221 B.n220 585
R480 B.n219 B.n52 585
R481 B.n218 B.n217 585
R482 B.n216 B.n53 585
R483 B.n215 B.n214 585
R484 B.n213 B.n54 585
R485 B.n212 B.n211 585
R486 B.n210 B.n55 585
R487 B.n209 B.n208 585
R488 B.n207 B.n56 585
R489 B.n206 B.n205 585
R490 B.n204 B.n57 585
R491 B.n203 B.n202 585
R492 B.n120 B.n89 585
R493 B.n122 B.n121 585
R494 B.n123 B.n88 585
R495 B.n125 B.n124 585
R496 B.n126 B.n87 585
R497 B.n128 B.n127 585
R498 B.n129 B.n86 585
R499 B.n131 B.n130 585
R500 B.n132 B.n85 585
R501 B.n134 B.n133 585
R502 B.n135 B.n84 585
R503 B.n137 B.n136 585
R504 B.n138 B.n83 585
R505 B.n140 B.n139 585
R506 B.n141 B.n82 585
R507 B.n143 B.n142 585
R508 B.n144 B.n81 585
R509 B.n146 B.n145 585
R510 B.n147 B.n80 585
R511 B.n149 B.n148 585
R512 B.n150 B.n79 585
R513 B.n152 B.n151 585
R514 B.n154 B.n153 585
R515 B.n155 B.n75 585
R516 B.n157 B.n156 585
R517 B.n158 B.n74 585
R518 B.n160 B.n159 585
R519 B.n161 B.n73 585
R520 B.n163 B.n162 585
R521 B.n164 B.n72 585
R522 B.n166 B.n165 585
R523 B.n167 B.n69 585
R524 B.n170 B.n169 585
R525 B.n171 B.n68 585
R526 B.n173 B.n172 585
R527 B.n174 B.n67 585
R528 B.n176 B.n175 585
R529 B.n177 B.n66 585
R530 B.n179 B.n178 585
R531 B.n180 B.n65 585
R532 B.n182 B.n181 585
R533 B.n183 B.n64 585
R534 B.n185 B.n184 585
R535 B.n186 B.n63 585
R536 B.n188 B.n187 585
R537 B.n189 B.n62 585
R538 B.n191 B.n190 585
R539 B.n192 B.n61 585
R540 B.n194 B.n193 585
R541 B.n195 B.n60 585
R542 B.n197 B.n196 585
R543 B.n198 B.n59 585
R544 B.n200 B.n199 585
R545 B.n201 B.n58 585
R546 B.n119 B.n118 585
R547 B.n117 B.n90 585
R548 B.n116 B.n115 585
R549 B.n114 B.n91 585
R550 B.n113 B.n112 585
R551 B.n111 B.n92 585
R552 B.n110 B.n109 585
R553 B.n108 B.n93 585
R554 B.n107 B.n106 585
R555 B.n105 B.n94 585
R556 B.n104 B.n103 585
R557 B.n102 B.n95 585
R558 B.n101 B.n100 585
R559 B.n99 B.n96 585
R560 B.n98 B.n97 585
R561 B.n2 B.n0 585
R562 B.n357 B.n1 585
R563 B.n356 B.n355 585
R564 B.n354 B.n3 585
R565 B.n353 B.n352 585
R566 B.n351 B.n4 585
R567 B.n350 B.n349 585
R568 B.n348 B.n5 585
R569 B.n347 B.n346 585
R570 B.n345 B.n6 585
R571 B.n344 B.n343 585
R572 B.n342 B.n7 585
R573 B.n341 B.n340 585
R574 B.n339 B.n8 585
R575 B.n338 B.n337 585
R576 B.n336 B.n9 585
R577 B.n335 B.n334 585
R578 B.n359 B.n358 585
R579 B.n118 B.n89 511.721
R580 B.n334 B.n333 511.721
R581 B.n202 B.n201 511.721
R582 B.n250 B.n41 511.721
R583 B.n70 B.t11 268.642
R584 B.n28 B.t7 268.642
R585 B.n76 B.t5 268.642
R586 B.n22 B.t1 268.642
R587 B.n71 B.t10 258.17
R588 B.n29 B.t8 258.17
R589 B.n77 B.t4 258.17
R590 B.n23 B.t2 258.17
R591 B.n118 B.n117 163.367
R592 B.n117 B.n116 163.367
R593 B.n116 B.n91 163.367
R594 B.n112 B.n91 163.367
R595 B.n112 B.n111 163.367
R596 B.n111 B.n110 163.367
R597 B.n110 B.n93 163.367
R598 B.n106 B.n93 163.367
R599 B.n106 B.n105 163.367
R600 B.n105 B.n104 163.367
R601 B.n104 B.n95 163.367
R602 B.n100 B.n95 163.367
R603 B.n100 B.n99 163.367
R604 B.n99 B.n98 163.367
R605 B.n98 B.n2 163.367
R606 B.n358 B.n2 163.367
R607 B.n358 B.n357 163.367
R608 B.n357 B.n356 163.367
R609 B.n356 B.n3 163.367
R610 B.n352 B.n3 163.367
R611 B.n352 B.n351 163.367
R612 B.n351 B.n350 163.367
R613 B.n350 B.n5 163.367
R614 B.n346 B.n5 163.367
R615 B.n346 B.n345 163.367
R616 B.n345 B.n344 163.367
R617 B.n344 B.n7 163.367
R618 B.n340 B.n7 163.367
R619 B.n340 B.n339 163.367
R620 B.n339 B.n338 163.367
R621 B.n338 B.n9 163.367
R622 B.n334 B.n9 163.367
R623 B.n122 B.n89 163.367
R624 B.n123 B.n122 163.367
R625 B.n124 B.n123 163.367
R626 B.n124 B.n87 163.367
R627 B.n128 B.n87 163.367
R628 B.n129 B.n128 163.367
R629 B.n130 B.n129 163.367
R630 B.n130 B.n85 163.367
R631 B.n134 B.n85 163.367
R632 B.n135 B.n134 163.367
R633 B.n136 B.n135 163.367
R634 B.n136 B.n83 163.367
R635 B.n140 B.n83 163.367
R636 B.n141 B.n140 163.367
R637 B.n142 B.n141 163.367
R638 B.n142 B.n81 163.367
R639 B.n146 B.n81 163.367
R640 B.n147 B.n146 163.367
R641 B.n148 B.n147 163.367
R642 B.n148 B.n79 163.367
R643 B.n152 B.n79 163.367
R644 B.n153 B.n152 163.367
R645 B.n153 B.n75 163.367
R646 B.n157 B.n75 163.367
R647 B.n158 B.n157 163.367
R648 B.n159 B.n158 163.367
R649 B.n159 B.n73 163.367
R650 B.n163 B.n73 163.367
R651 B.n164 B.n163 163.367
R652 B.n165 B.n164 163.367
R653 B.n165 B.n69 163.367
R654 B.n170 B.n69 163.367
R655 B.n171 B.n170 163.367
R656 B.n172 B.n171 163.367
R657 B.n172 B.n67 163.367
R658 B.n176 B.n67 163.367
R659 B.n177 B.n176 163.367
R660 B.n178 B.n177 163.367
R661 B.n178 B.n65 163.367
R662 B.n182 B.n65 163.367
R663 B.n183 B.n182 163.367
R664 B.n184 B.n183 163.367
R665 B.n184 B.n63 163.367
R666 B.n188 B.n63 163.367
R667 B.n189 B.n188 163.367
R668 B.n190 B.n189 163.367
R669 B.n190 B.n61 163.367
R670 B.n194 B.n61 163.367
R671 B.n195 B.n194 163.367
R672 B.n196 B.n195 163.367
R673 B.n196 B.n59 163.367
R674 B.n200 B.n59 163.367
R675 B.n201 B.n200 163.367
R676 B.n202 B.n57 163.367
R677 B.n206 B.n57 163.367
R678 B.n207 B.n206 163.367
R679 B.n208 B.n207 163.367
R680 B.n208 B.n55 163.367
R681 B.n212 B.n55 163.367
R682 B.n213 B.n212 163.367
R683 B.n214 B.n213 163.367
R684 B.n214 B.n53 163.367
R685 B.n218 B.n53 163.367
R686 B.n219 B.n218 163.367
R687 B.n220 B.n219 163.367
R688 B.n220 B.n51 163.367
R689 B.n224 B.n51 163.367
R690 B.n225 B.n224 163.367
R691 B.n226 B.n225 163.367
R692 B.n226 B.n49 163.367
R693 B.n230 B.n49 163.367
R694 B.n231 B.n230 163.367
R695 B.n232 B.n231 163.367
R696 B.n232 B.n47 163.367
R697 B.n236 B.n47 163.367
R698 B.n237 B.n236 163.367
R699 B.n238 B.n237 163.367
R700 B.n238 B.n45 163.367
R701 B.n242 B.n45 163.367
R702 B.n243 B.n242 163.367
R703 B.n244 B.n243 163.367
R704 B.n244 B.n43 163.367
R705 B.n248 B.n43 163.367
R706 B.n249 B.n248 163.367
R707 B.n250 B.n249 163.367
R708 B.n333 B.n332 163.367
R709 B.n332 B.n11 163.367
R710 B.n328 B.n11 163.367
R711 B.n328 B.n327 163.367
R712 B.n327 B.n326 163.367
R713 B.n326 B.n13 163.367
R714 B.n322 B.n13 163.367
R715 B.n322 B.n321 163.367
R716 B.n321 B.n320 163.367
R717 B.n320 B.n15 163.367
R718 B.n316 B.n15 163.367
R719 B.n316 B.n315 163.367
R720 B.n315 B.n314 163.367
R721 B.n314 B.n17 163.367
R722 B.n310 B.n17 163.367
R723 B.n310 B.n309 163.367
R724 B.n309 B.n308 163.367
R725 B.n308 B.n19 163.367
R726 B.n304 B.n19 163.367
R727 B.n304 B.n303 163.367
R728 B.n303 B.n302 163.367
R729 B.n302 B.n21 163.367
R730 B.n297 B.n21 163.367
R731 B.n297 B.n296 163.367
R732 B.n296 B.n295 163.367
R733 B.n295 B.n25 163.367
R734 B.n291 B.n25 163.367
R735 B.n291 B.n290 163.367
R736 B.n290 B.n289 163.367
R737 B.n289 B.n27 163.367
R738 B.n285 B.n27 163.367
R739 B.n285 B.n284 163.367
R740 B.n284 B.n31 163.367
R741 B.n280 B.n31 163.367
R742 B.n280 B.n279 163.367
R743 B.n279 B.n278 163.367
R744 B.n278 B.n33 163.367
R745 B.n274 B.n33 163.367
R746 B.n274 B.n273 163.367
R747 B.n273 B.n272 163.367
R748 B.n272 B.n35 163.367
R749 B.n268 B.n35 163.367
R750 B.n268 B.n267 163.367
R751 B.n267 B.n266 163.367
R752 B.n266 B.n37 163.367
R753 B.n262 B.n37 163.367
R754 B.n262 B.n261 163.367
R755 B.n261 B.n260 163.367
R756 B.n260 B.n39 163.367
R757 B.n256 B.n39 163.367
R758 B.n256 B.n255 163.367
R759 B.n255 B.n254 163.367
R760 B.n254 B.n41 163.367
R761 B.n168 B.n71 59.5399
R762 B.n78 B.n77 59.5399
R763 B.n300 B.n23 59.5399
R764 B.n30 B.n29 59.5399
R765 B.n335 B.n10 33.2493
R766 B.n252 B.n251 33.2493
R767 B.n203 B.n58 33.2493
R768 B.n120 B.n119 33.2493
R769 B B.n359 18.0485
R770 B.n331 B.n10 10.6151
R771 B.n331 B.n330 10.6151
R772 B.n330 B.n329 10.6151
R773 B.n329 B.n12 10.6151
R774 B.n325 B.n12 10.6151
R775 B.n325 B.n324 10.6151
R776 B.n324 B.n323 10.6151
R777 B.n323 B.n14 10.6151
R778 B.n319 B.n14 10.6151
R779 B.n319 B.n318 10.6151
R780 B.n318 B.n317 10.6151
R781 B.n317 B.n16 10.6151
R782 B.n313 B.n16 10.6151
R783 B.n313 B.n312 10.6151
R784 B.n312 B.n311 10.6151
R785 B.n311 B.n18 10.6151
R786 B.n307 B.n18 10.6151
R787 B.n307 B.n306 10.6151
R788 B.n306 B.n305 10.6151
R789 B.n305 B.n20 10.6151
R790 B.n301 B.n20 10.6151
R791 B.n299 B.n298 10.6151
R792 B.n298 B.n24 10.6151
R793 B.n294 B.n24 10.6151
R794 B.n294 B.n293 10.6151
R795 B.n293 B.n292 10.6151
R796 B.n292 B.n26 10.6151
R797 B.n288 B.n26 10.6151
R798 B.n288 B.n287 10.6151
R799 B.n287 B.n286 10.6151
R800 B.n283 B.n282 10.6151
R801 B.n282 B.n281 10.6151
R802 B.n281 B.n32 10.6151
R803 B.n277 B.n32 10.6151
R804 B.n277 B.n276 10.6151
R805 B.n276 B.n275 10.6151
R806 B.n275 B.n34 10.6151
R807 B.n271 B.n34 10.6151
R808 B.n271 B.n270 10.6151
R809 B.n270 B.n269 10.6151
R810 B.n269 B.n36 10.6151
R811 B.n265 B.n36 10.6151
R812 B.n265 B.n264 10.6151
R813 B.n264 B.n263 10.6151
R814 B.n263 B.n38 10.6151
R815 B.n259 B.n38 10.6151
R816 B.n259 B.n258 10.6151
R817 B.n258 B.n257 10.6151
R818 B.n257 B.n40 10.6151
R819 B.n253 B.n40 10.6151
R820 B.n253 B.n252 10.6151
R821 B.n204 B.n203 10.6151
R822 B.n205 B.n204 10.6151
R823 B.n205 B.n56 10.6151
R824 B.n209 B.n56 10.6151
R825 B.n210 B.n209 10.6151
R826 B.n211 B.n210 10.6151
R827 B.n211 B.n54 10.6151
R828 B.n215 B.n54 10.6151
R829 B.n216 B.n215 10.6151
R830 B.n217 B.n216 10.6151
R831 B.n217 B.n52 10.6151
R832 B.n221 B.n52 10.6151
R833 B.n222 B.n221 10.6151
R834 B.n223 B.n222 10.6151
R835 B.n223 B.n50 10.6151
R836 B.n227 B.n50 10.6151
R837 B.n228 B.n227 10.6151
R838 B.n229 B.n228 10.6151
R839 B.n229 B.n48 10.6151
R840 B.n233 B.n48 10.6151
R841 B.n234 B.n233 10.6151
R842 B.n235 B.n234 10.6151
R843 B.n235 B.n46 10.6151
R844 B.n239 B.n46 10.6151
R845 B.n240 B.n239 10.6151
R846 B.n241 B.n240 10.6151
R847 B.n241 B.n44 10.6151
R848 B.n245 B.n44 10.6151
R849 B.n246 B.n245 10.6151
R850 B.n247 B.n246 10.6151
R851 B.n247 B.n42 10.6151
R852 B.n251 B.n42 10.6151
R853 B.n121 B.n120 10.6151
R854 B.n121 B.n88 10.6151
R855 B.n125 B.n88 10.6151
R856 B.n126 B.n125 10.6151
R857 B.n127 B.n126 10.6151
R858 B.n127 B.n86 10.6151
R859 B.n131 B.n86 10.6151
R860 B.n132 B.n131 10.6151
R861 B.n133 B.n132 10.6151
R862 B.n133 B.n84 10.6151
R863 B.n137 B.n84 10.6151
R864 B.n138 B.n137 10.6151
R865 B.n139 B.n138 10.6151
R866 B.n139 B.n82 10.6151
R867 B.n143 B.n82 10.6151
R868 B.n144 B.n143 10.6151
R869 B.n145 B.n144 10.6151
R870 B.n145 B.n80 10.6151
R871 B.n149 B.n80 10.6151
R872 B.n150 B.n149 10.6151
R873 B.n151 B.n150 10.6151
R874 B.n155 B.n154 10.6151
R875 B.n156 B.n155 10.6151
R876 B.n156 B.n74 10.6151
R877 B.n160 B.n74 10.6151
R878 B.n161 B.n160 10.6151
R879 B.n162 B.n161 10.6151
R880 B.n162 B.n72 10.6151
R881 B.n166 B.n72 10.6151
R882 B.n167 B.n166 10.6151
R883 B.n169 B.n68 10.6151
R884 B.n173 B.n68 10.6151
R885 B.n174 B.n173 10.6151
R886 B.n175 B.n174 10.6151
R887 B.n175 B.n66 10.6151
R888 B.n179 B.n66 10.6151
R889 B.n180 B.n179 10.6151
R890 B.n181 B.n180 10.6151
R891 B.n181 B.n64 10.6151
R892 B.n185 B.n64 10.6151
R893 B.n186 B.n185 10.6151
R894 B.n187 B.n186 10.6151
R895 B.n187 B.n62 10.6151
R896 B.n191 B.n62 10.6151
R897 B.n192 B.n191 10.6151
R898 B.n193 B.n192 10.6151
R899 B.n193 B.n60 10.6151
R900 B.n197 B.n60 10.6151
R901 B.n198 B.n197 10.6151
R902 B.n199 B.n198 10.6151
R903 B.n199 B.n58 10.6151
R904 B.n119 B.n90 10.6151
R905 B.n115 B.n90 10.6151
R906 B.n115 B.n114 10.6151
R907 B.n114 B.n113 10.6151
R908 B.n113 B.n92 10.6151
R909 B.n109 B.n92 10.6151
R910 B.n109 B.n108 10.6151
R911 B.n108 B.n107 10.6151
R912 B.n107 B.n94 10.6151
R913 B.n103 B.n94 10.6151
R914 B.n103 B.n102 10.6151
R915 B.n102 B.n101 10.6151
R916 B.n101 B.n96 10.6151
R917 B.n97 B.n96 10.6151
R918 B.n97 B.n0 10.6151
R919 B.n355 B.n1 10.6151
R920 B.n355 B.n354 10.6151
R921 B.n354 B.n353 10.6151
R922 B.n353 B.n4 10.6151
R923 B.n349 B.n4 10.6151
R924 B.n349 B.n348 10.6151
R925 B.n348 B.n347 10.6151
R926 B.n347 B.n6 10.6151
R927 B.n343 B.n6 10.6151
R928 B.n343 B.n342 10.6151
R929 B.n342 B.n341 10.6151
R930 B.n341 B.n8 10.6151
R931 B.n337 B.n8 10.6151
R932 B.n337 B.n336 10.6151
R933 B.n336 B.n335 10.6151
R934 B.n71 B.n70 10.4732
R935 B.n77 B.n76 10.4732
R936 B.n23 B.n22 10.4732
R937 B.n29 B.n28 10.4732
R938 B.n301 B.n300 9.36635
R939 B.n283 B.n30 9.36635
R940 B.n151 B.n78 9.36635
R941 B.n169 B.n168 9.36635
R942 B.n359 B.n0 2.81026
R943 B.n359 B.n1 2.81026
R944 B.n300 B.n299 1.24928
R945 B.n286 B.n30 1.24928
R946 B.n154 B.n78 1.24928
R947 B.n168 B.n167 1.24928
R948 VP.n13 VP.t6 816.48
R949 VP.n9 VP.t7 816.48
R950 VP.n2 VP.t2 816.48
R951 VP.n6 VP.t1 816.48
R952 VP.n12 VP.t0 771.201
R953 VP.n10 VP.t3 771.201
R954 VP.n3 VP.t4 771.201
R955 VP.n5 VP.t5 771.201
R956 VP.n2 VP.n1 161.489
R957 VP.n14 VP.n13 161.3
R958 VP.n4 VP.n1 161.3
R959 VP.n7 VP.n6 161.3
R960 VP.n11 VP.n0 161.3
R961 VP.n9 VP.n8 161.3
R962 VP.n11 VP.n10 39.4369
R963 VP.n12 VP.n11 39.4369
R964 VP.n4 VP.n3 39.4369
R965 VP.n5 VP.n4 39.4369
R966 VP.n8 VP.n7 34.7884
R967 VP.n10 VP.n9 33.5944
R968 VP.n13 VP.n12 33.5944
R969 VP.n3 VP.n2 33.5944
R970 VP.n6 VP.n5 33.5944
R971 VP.n7 VP.n1 0.189894
R972 VP.n8 VP.n0 0.189894
R973 VP.n14 VP.n0 0.189894
R974 VP VP.n14 0.0516364
R975 VDD1 VDD1.n0 100.144
R976 VDD1.n3 VDD1.n2 100.029
R977 VDD1.n3 VDD1.n1 100.029
R978 VDD1.n5 VDD1.n4 99.852
R979 VDD1.n5 VDD1.n3 31.0569
R980 VDD1.n4 VDD1.t2 6.00882
R981 VDD1.n4 VDD1.t6 6.00882
R982 VDD1.n0 VDD1.t5 6.00882
R983 VDD1.n0 VDD1.t3 6.00882
R984 VDD1.n2 VDD1.t7 6.00882
R985 VDD1.n2 VDD1.t1 6.00882
R986 VDD1.n1 VDD1.t0 6.00882
R987 VDD1.n1 VDD1.t4 6.00882
R988 VDD1 VDD1.n5 0.175069
C0 VN VDD2 1.40138f
C1 VTAIL VDD2 9.604731f
C2 VP VDD1 1.51913f
C3 B VDD2 0.764704f
C4 VDD1 VTAIL 9.56634f
C5 VN VDD1 0.146975f
C6 VP w_n1510_n2050# 2.47201f
C7 VDD1 B 0.742616f
C8 VDD1 VDD2 0.587463f
C9 VN w_n1510_n2050# 2.28306f
C10 VTAIL w_n1510_n2050# 2.53914f
C11 w_n1510_n2050# B 4.66605f
C12 w_n1510_n2050# VDD2 0.927313f
C13 VDD1 w_n1510_n2050# 0.912571f
C14 VN VP 3.51944f
C15 VP VTAIL 1.25574f
C16 VP B 0.88868f
C17 VN VTAIL 1.24163f
C18 VP VDD2 0.268756f
C19 VN B 0.584623f
C20 VTAIL B 1.79458f
C21 VDD2 VSUBS 1.02724f
C22 VDD1 VSUBS 1.229835f
C23 VTAIL VSUBS 0.372824f
C24 VN VSUBS 3.07616f
C25 VP VSUBS 0.850014f
C26 B VSUBS 1.710946f
C27 w_n1510_n2050# VSUBS 38.7224f
C28 VDD1.t5 VSUBS 0.130821f
C29 VDD1.t3 VSUBS 0.130821f
C30 VDD1.n0 VSUBS 0.845665f
C31 VDD1.t0 VSUBS 0.130821f
C32 VDD1.t4 VSUBS 0.130821f
C33 VDD1.n1 VSUBS 0.845008f
C34 VDD1.t7 VSUBS 0.130821f
C35 VDD1.t1 VSUBS 0.130821f
C36 VDD1.n2 VSUBS 0.845008f
C37 VDD1.n3 VSUBS 2.35013f
C38 VDD1.t2 VSUBS 0.130821f
C39 VDD1.t6 VSUBS 0.130821f
C40 VDD1.n4 VSUBS 0.844017f
C41 VDD1.n5 VSUBS 2.21381f
C42 VP.n0 VSUBS 0.056873f
C43 VP.t0 VSUBS 0.184536f
C44 VP.t3 VSUBS 0.184536f
C45 VP.t7 VSUBS 0.189705f
C46 VP.n1 VSUBS 0.125237f
C47 VP.t5 VSUBS 0.184536f
C48 VP.t4 VSUBS 0.184536f
C49 VP.t2 VSUBS 0.189705f
C50 VP.n2 VSUBS 0.108389f
C51 VP.n3 VSUBS 0.092507f
C52 VP.n4 VSUBS 0.020269f
C53 VP.n5 VSUBS 0.092507f
C54 VP.t1 VSUBS 0.189705f
C55 VP.n6 VSUBS 0.108309f
C56 VP.n7 VSUBS 1.67492f
C57 VP.n8 VSUBS 1.73368f
C58 VP.n9 VSUBS 0.108309f
C59 VP.n10 VSUBS 0.092507f
C60 VP.n11 VSUBS 0.020269f
C61 VP.n12 VSUBS 0.092507f
C62 VP.t6 VSUBS 0.189705f
C63 VP.n13 VSUBS 0.108309f
C64 VP.n14 VSUBS 0.044075f
C65 B.n0 VSUBS 0.004524f
C66 B.n1 VSUBS 0.004524f
C67 B.n2 VSUBS 0.007155f
C68 B.n3 VSUBS 0.007155f
C69 B.n4 VSUBS 0.007155f
C70 B.n5 VSUBS 0.007155f
C71 B.n6 VSUBS 0.007155f
C72 B.n7 VSUBS 0.007155f
C73 B.n8 VSUBS 0.007155f
C74 B.n9 VSUBS 0.007155f
C75 B.n10 VSUBS 0.017356f
C76 B.n11 VSUBS 0.007155f
C77 B.n12 VSUBS 0.007155f
C78 B.n13 VSUBS 0.007155f
C79 B.n14 VSUBS 0.007155f
C80 B.n15 VSUBS 0.007155f
C81 B.n16 VSUBS 0.007155f
C82 B.n17 VSUBS 0.007155f
C83 B.n18 VSUBS 0.007155f
C84 B.n19 VSUBS 0.007155f
C85 B.n20 VSUBS 0.007155f
C86 B.n21 VSUBS 0.007155f
C87 B.t2 VSUBS 0.081463f
C88 B.t1 VSUBS 0.086445f
C89 B.t0 VSUBS 0.046703f
C90 B.n22 VSUBS 0.144571f
C91 B.n23 VSUBS 0.137986f
C92 B.n24 VSUBS 0.007155f
C93 B.n25 VSUBS 0.007155f
C94 B.n26 VSUBS 0.007155f
C95 B.n27 VSUBS 0.007155f
C96 B.t8 VSUBS 0.081465f
C97 B.t7 VSUBS 0.086446f
C98 B.t6 VSUBS 0.046703f
C99 B.n28 VSUBS 0.14457f
C100 B.n29 VSUBS 0.137984f
C101 B.n30 VSUBS 0.016577f
C102 B.n31 VSUBS 0.007155f
C103 B.n32 VSUBS 0.007155f
C104 B.n33 VSUBS 0.007155f
C105 B.n34 VSUBS 0.007155f
C106 B.n35 VSUBS 0.007155f
C107 B.n36 VSUBS 0.007155f
C108 B.n37 VSUBS 0.007155f
C109 B.n38 VSUBS 0.007155f
C110 B.n39 VSUBS 0.007155f
C111 B.n40 VSUBS 0.007155f
C112 B.n41 VSUBS 0.017356f
C113 B.n42 VSUBS 0.007155f
C114 B.n43 VSUBS 0.007155f
C115 B.n44 VSUBS 0.007155f
C116 B.n45 VSUBS 0.007155f
C117 B.n46 VSUBS 0.007155f
C118 B.n47 VSUBS 0.007155f
C119 B.n48 VSUBS 0.007155f
C120 B.n49 VSUBS 0.007155f
C121 B.n50 VSUBS 0.007155f
C122 B.n51 VSUBS 0.007155f
C123 B.n52 VSUBS 0.007155f
C124 B.n53 VSUBS 0.007155f
C125 B.n54 VSUBS 0.007155f
C126 B.n55 VSUBS 0.007155f
C127 B.n56 VSUBS 0.007155f
C128 B.n57 VSUBS 0.007155f
C129 B.n58 VSUBS 0.017356f
C130 B.n59 VSUBS 0.007155f
C131 B.n60 VSUBS 0.007155f
C132 B.n61 VSUBS 0.007155f
C133 B.n62 VSUBS 0.007155f
C134 B.n63 VSUBS 0.007155f
C135 B.n64 VSUBS 0.007155f
C136 B.n65 VSUBS 0.007155f
C137 B.n66 VSUBS 0.007155f
C138 B.n67 VSUBS 0.007155f
C139 B.n68 VSUBS 0.007155f
C140 B.n69 VSUBS 0.007155f
C141 B.t10 VSUBS 0.081465f
C142 B.t11 VSUBS 0.086446f
C143 B.t9 VSUBS 0.046703f
C144 B.n70 VSUBS 0.14457f
C145 B.n71 VSUBS 0.137984f
C146 B.n72 VSUBS 0.007155f
C147 B.n73 VSUBS 0.007155f
C148 B.n74 VSUBS 0.007155f
C149 B.n75 VSUBS 0.007155f
C150 B.t4 VSUBS 0.081463f
C151 B.t5 VSUBS 0.086445f
C152 B.t3 VSUBS 0.046703f
C153 B.n76 VSUBS 0.144571f
C154 B.n77 VSUBS 0.137986f
C155 B.n78 VSUBS 0.016577f
C156 B.n79 VSUBS 0.007155f
C157 B.n80 VSUBS 0.007155f
C158 B.n81 VSUBS 0.007155f
C159 B.n82 VSUBS 0.007155f
C160 B.n83 VSUBS 0.007155f
C161 B.n84 VSUBS 0.007155f
C162 B.n85 VSUBS 0.007155f
C163 B.n86 VSUBS 0.007155f
C164 B.n87 VSUBS 0.007155f
C165 B.n88 VSUBS 0.007155f
C166 B.n89 VSUBS 0.017356f
C167 B.n90 VSUBS 0.007155f
C168 B.n91 VSUBS 0.007155f
C169 B.n92 VSUBS 0.007155f
C170 B.n93 VSUBS 0.007155f
C171 B.n94 VSUBS 0.007155f
C172 B.n95 VSUBS 0.007155f
C173 B.n96 VSUBS 0.007155f
C174 B.n97 VSUBS 0.007155f
C175 B.n98 VSUBS 0.007155f
C176 B.n99 VSUBS 0.007155f
C177 B.n100 VSUBS 0.007155f
C178 B.n101 VSUBS 0.007155f
C179 B.n102 VSUBS 0.007155f
C180 B.n103 VSUBS 0.007155f
C181 B.n104 VSUBS 0.007155f
C182 B.n105 VSUBS 0.007155f
C183 B.n106 VSUBS 0.007155f
C184 B.n107 VSUBS 0.007155f
C185 B.n108 VSUBS 0.007155f
C186 B.n109 VSUBS 0.007155f
C187 B.n110 VSUBS 0.007155f
C188 B.n111 VSUBS 0.007155f
C189 B.n112 VSUBS 0.007155f
C190 B.n113 VSUBS 0.007155f
C191 B.n114 VSUBS 0.007155f
C192 B.n115 VSUBS 0.007155f
C193 B.n116 VSUBS 0.007155f
C194 B.n117 VSUBS 0.007155f
C195 B.n118 VSUBS 0.016525f
C196 B.n119 VSUBS 0.016525f
C197 B.n120 VSUBS 0.017356f
C198 B.n121 VSUBS 0.007155f
C199 B.n122 VSUBS 0.007155f
C200 B.n123 VSUBS 0.007155f
C201 B.n124 VSUBS 0.007155f
C202 B.n125 VSUBS 0.007155f
C203 B.n126 VSUBS 0.007155f
C204 B.n127 VSUBS 0.007155f
C205 B.n128 VSUBS 0.007155f
C206 B.n129 VSUBS 0.007155f
C207 B.n130 VSUBS 0.007155f
C208 B.n131 VSUBS 0.007155f
C209 B.n132 VSUBS 0.007155f
C210 B.n133 VSUBS 0.007155f
C211 B.n134 VSUBS 0.007155f
C212 B.n135 VSUBS 0.007155f
C213 B.n136 VSUBS 0.007155f
C214 B.n137 VSUBS 0.007155f
C215 B.n138 VSUBS 0.007155f
C216 B.n139 VSUBS 0.007155f
C217 B.n140 VSUBS 0.007155f
C218 B.n141 VSUBS 0.007155f
C219 B.n142 VSUBS 0.007155f
C220 B.n143 VSUBS 0.007155f
C221 B.n144 VSUBS 0.007155f
C222 B.n145 VSUBS 0.007155f
C223 B.n146 VSUBS 0.007155f
C224 B.n147 VSUBS 0.007155f
C225 B.n148 VSUBS 0.007155f
C226 B.n149 VSUBS 0.007155f
C227 B.n150 VSUBS 0.007155f
C228 B.n151 VSUBS 0.006734f
C229 B.n152 VSUBS 0.007155f
C230 B.n153 VSUBS 0.007155f
C231 B.n154 VSUBS 0.003998f
C232 B.n155 VSUBS 0.007155f
C233 B.n156 VSUBS 0.007155f
C234 B.n157 VSUBS 0.007155f
C235 B.n158 VSUBS 0.007155f
C236 B.n159 VSUBS 0.007155f
C237 B.n160 VSUBS 0.007155f
C238 B.n161 VSUBS 0.007155f
C239 B.n162 VSUBS 0.007155f
C240 B.n163 VSUBS 0.007155f
C241 B.n164 VSUBS 0.007155f
C242 B.n165 VSUBS 0.007155f
C243 B.n166 VSUBS 0.007155f
C244 B.n167 VSUBS 0.003998f
C245 B.n168 VSUBS 0.016577f
C246 B.n169 VSUBS 0.006734f
C247 B.n170 VSUBS 0.007155f
C248 B.n171 VSUBS 0.007155f
C249 B.n172 VSUBS 0.007155f
C250 B.n173 VSUBS 0.007155f
C251 B.n174 VSUBS 0.007155f
C252 B.n175 VSUBS 0.007155f
C253 B.n176 VSUBS 0.007155f
C254 B.n177 VSUBS 0.007155f
C255 B.n178 VSUBS 0.007155f
C256 B.n179 VSUBS 0.007155f
C257 B.n180 VSUBS 0.007155f
C258 B.n181 VSUBS 0.007155f
C259 B.n182 VSUBS 0.007155f
C260 B.n183 VSUBS 0.007155f
C261 B.n184 VSUBS 0.007155f
C262 B.n185 VSUBS 0.007155f
C263 B.n186 VSUBS 0.007155f
C264 B.n187 VSUBS 0.007155f
C265 B.n188 VSUBS 0.007155f
C266 B.n189 VSUBS 0.007155f
C267 B.n190 VSUBS 0.007155f
C268 B.n191 VSUBS 0.007155f
C269 B.n192 VSUBS 0.007155f
C270 B.n193 VSUBS 0.007155f
C271 B.n194 VSUBS 0.007155f
C272 B.n195 VSUBS 0.007155f
C273 B.n196 VSUBS 0.007155f
C274 B.n197 VSUBS 0.007155f
C275 B.n198 VSUBS 0.007155f
C276 B.n199 VSUBS 0.007155f
C277 B.n200 VSUBS 0.007155f
C278 B.n201 VSUBS 0.017356f
C279 B.n202 VSUBS 0.016525f
C280 B.n203 VSUBS 0.016525f
C281 B.n204 VSUBS 0.007155f
C282 B.n205 VSUBS 0.007155f
C283 B.n206 VSUBS 0.007155f
C284 B.n207 VSUBS 0.007155f
C285 B.n208 VSUBS 0.007155f
C286 B.n209 VSUBS 0.007155f
C287 B.n210 VSUBS 0.007155f
C288 B.n211 VSUBS 0.007155f
C289 B.n212 VSUBS 0.007155f
C290 B.n213 VSUBS 0.007155f
C291 B.n214 VSUBS 0.007155f
C292 B.n215 VSUBS 0.007155f
C293 B.n216 VSUBS 0.007155f
C294 B.n217 VSUBS 0.007155f
C295 B.n218 VSUBS 0.007155f
C296 B.n219 VSUBS 0.007155f
C297 B.n220 VSUBS 0.007155f
C298 B.n221 VSUBS 0.007155f
C299 B.n222 VSUBS 0.007155f
C300 B.n223 VSUBS 0.007155f
C301 B.n224 VSUBS 0.007155f
C302 B.n225 VSUBS 0.007155f
C303 B.n226 VSUBS 0.007155f
C304 B.n227 VSUBS 0.007155f
C305 B.n228 VSUBS 0.007155f
C306 B.n229 VSUBS 0.007155f
C307 B.n230 VSUBS 0.007155f
C308 B.n231 VSUBS 0.007155f
C309 B.n232 VSUBS 0.007155f
C310 B.n233 VSUBS 0.007155f
C311 B.n234 VSUBS 0.007155f
C312 B.n235 VSUBS 0.007155f
C313 B.n236 VSUBS 0.007155f
C314 B.n237 VSUBS 0.007155f
C315 B.n238 VSUBS 0.007155f
C316 B.n239 VSUBS 0.007155f
C317 B.n240 VSUBS 0.007155f
C318 B.n241 VSUBS 0.007155f
C319 B.n242 VSUBS 0.007155f
C320 B.n243 VSUBS 0.007155f
C321 B.n244 VSUBS 0.007155f
C322 B.n245 VSUBS 0.007155f
C323 B.n246 VSUBS 0.007155f
C324 B.n247 VSUBS 0.007155f
C325 B.n248 VSUBS 0.007155f
C326 B.n249 VSUBS 0.007155f
C327 B.n250 VSUBS 0.016525f
C328 B.n251 VSUBS 0.017356f
C329 B.n252 VSUBS 0.016525f
C330 B.n253 VSUBS 0.007155f
C331 B.n254 VSUBS 0.007155f
C332 B.n255 VSUBS 0.007155f
C333 B.n256 VSUBS 0.007155f
C334 B.n257 VSUBS 0.007155f
C335 B.n258 VSUBS 0.007155f
C336 B.n259 VSUBS 0.007155f
C337 B.n260 VSUBS 0.007155f
C338 B.n261 VSUBS 0.007155f
C339 B.n262 VSUBS 0.007155f
C340 B.n263 VSUBS 0.007155f
C341 B.n264 VSUBS 0.007155f
C342 B.n265 VSUBS 0.007155f
C343 B.n266 VSUBS 0.007155f
C344 B.n267 VSUBS 0.007155f
C345 B.n268 VSUBS 0.007155f
C346 B.n269 VSUBS 0.007155f
C347 B.n270 VSUBS 0.007155f
C348 B.n271 VSUBS 0.007155f
C349 B.n272 VSUBS 0.007155f
C350 B.n273 VSUBS 0.007155f
C351 B.n274 VSUBS 0.007155f
C352 B.n275 VSUBS 0.007155f
C353 B.n276 VSUBS 0.007155f
C354 B.n277 VSUBS 0.007155f
C355 B.n278 VSUBS 0.007155f
C356 B.n279 VSUBS 0.007155f
C357 B.n280 VSUBS 0.007155f
C358 B.n281 VSUBS 0.007155f
C359 B.n282 VSUBS 0.007155f
C360 B.n283 VSUBS 0.006734f
C361 B.n284 VSUBS 0.007155f
C362 B.n285 VSUBS 0.007155f
C363 B.n286 VSUBS 0.003998f
C364 B.n287 VSUBS 0.007155f
C365 B.n288 VSUBS 0.007155f
C366 B.n289 VSUBS 0.007155f
C367 B.n290 VSUBS 0.007155f
C368 B.n291 VSUBS 0.007155f
C369 B.n292 VSUBS 0.007155f
C370 B.n293 VSUBS 0.007155f
C371 B.n294 VSUBS 0.007155f
C372 B.n295 VSUBS 0.007155f
C373 B.n296 VSUBS 0.007155f
C374 B.n297 VSUBS 0.007155f
C375 B.n298 VSUBS 0.007155f
C376 B.n299 VSUBS 0.003998f
C377 B.n300 VSUBS 0.016577f
C378 B.n301 VSUBS 0.006734f
C379 B.n302 VSUBS 0.007155f
C380 B.n303 VSUBS 0.007155f
C381 B.n304 VSUBS 0.007155f
C382 B.n305 VSUBS 0.007155f
C383 B.n306 VSUBS 0.007155f
C384 B.n307 VSUBS 0.007155f
C385 B.n308 VSUBS 0.007155f
C386 B.n309 VSUBS 0.007155f
C387 B.n310 VSUBS 0.007155f
C388 B.n311 VSUBS 0.007155f
C389 B.n312 VSUBS 0.007155f
C390 B.n313 VSUBS 0.007155f
C391 B.n314 VSUBS 0.007155f
C392 B.n315 VSUBS 0.007155f
C393 B.n316 VSUBS 0.007155f
C394 B.n317 VSUBS 0.007155f
C395 B.n318 VSUBS 0.007155f
C396 B.n319 VSUBS 0.007155f
C397 B.n320 VSUBS 0.007155f
C398 B.n321 VSUBS 0.007155f
C399 B.n322 VSUBS 0.007155f
C400 B.n323 VSUBS 0.007155f
C401 B.n324 VSUBS 0.007155f
C402 B.n325 VSUBS 0.007155f
C403 B.n326 VSUBS 0.007155f
C404 B.n327 VSUBS 0.007155f
C405 B.n328 VSUBS 0.007155f
C406 B.n329 VSUBS 0.007155f
C407 B.n330 VSUBS 0.007155f
C408 B.n331 VSUBS 0.007155f
C409 B.n332 VSUBS 0.007155f
C410 B.n333 VSUBS 0.017356f
C411 B.n334 VSUBS 0.016525f
C412 B.n335 VSUBS 0.016525f
C413 B.n336 VSUBS 0.007155f
C414 B.n337 VSUBS 0.007155f
C415 B.n338 VSUBS 0.007155f
C416 B.n339 VSUBS 0.007155f
C417 B.n340 VSUBS 0.007155f
C418 B.n341 VSUBS 0.007155f
C419 B.n342 VSUBS 0.007155f
C420 B.n343 VSUBS 0.007155f
C421 B.n344 VSUBS 0.007155f
C422 B.n345 VSUBS 0.007155f
C423 B.n346 VSUBS 0.007155f
C424 B.n347 VSUBS 0.007155f
C425 B.n348 VSUBS 0.007155f
C426 B.n349 VSUBS 0.007155f
C427 B.n350 VSUBS 0.007155f
C428 B.n351 VSUBS 0.007155f
C429 B.n352 VSUBS 0.007155f
C430 B.n353 VSUBS 0.007155f
C431 B.n354 VSUBS 0.007155f
C432 B.n355 VSUBS 0.007155f
C433 B.n356 VSUBS 0.007155f
C434 B.n357 VSUBS 0.007155f
C435 B.n358 VSUBS 0.007155f
C436 B.n359 VSUBS 0.016201f
C437 VDD2.t2 VSUBS 0.132379f
C438 VDD2.t0 VSUBS 0.132379f
C439 VDD2.n0 VSUBS 0.855075f
C440 VDD2.t5 VSUBS 0.132379f
C441 VDD2.t7 VSUBS 0.132379f
C442 VDD2.n1 VSUBS 0.855075f
C443 VDD2.n2 VSUBS 2.31123f
C444 VDD2.t1 VSUBS 0.132379f
C445 VDD2.t3 VSUBS 0.132379f
C446 VDD2.n3 VSUBS 0.854077f
C447 VDD2.n4 VSUBS 2.20433f
C448 VDD2.t4 VSUBS 0.132379f
C449 VDD2.t6 VSUBS 0.132379f
C450 VDD2.n5 VSUBS 0.855051f
C451 VTAIL.t11 VSUBS 0.118884f
C452 VTAIL.t14 VSUBS 0.118884f
C453 VTAIL.n0 VSUBS 0.680844f
C454 VTAIL.n1 VSUBS 0.530243f
C455 VTAIL.n2 VSUBS 0.0315f
C456 VTAIL.n3 VSUBS 0.027808f
C457 VTAIL.n4 VSUBS 0.014943f
C458 VTAIL.n5 VSUBS 0.03532f
C459 VTAIL.n6 VSUBS 0.015822f
C460 VTAIL.n7 VSUBS 0.027808f
C461 VTAIL.n8 VSUBS 0.014943f
C462 VTAIL.n9 VSUBS 0.02649f
C463 VTAIL.n10 VSUBS 0.022435f
C464 VTAIL.t9 VSUBS 0.076499f
C465 VTAIL.n11 VSUBS 0.11879f
C466 VTAIL.n12 VSUBS 0.56201f
C467 VTAIL.n13 VSUBS 0.014943f
C468 VTAIL.n14 VSUBS 0.015822f
C469 VTAIL.n15 VSUBS 0.03532f
C470 VTAIL.n16 VSUBS 0.03532f
C471 VTAIL.n17 VSUBS 0.015822f
C472 VTAIL.n18 VSUBS 0.014943f
C473 VTAIL.n19 VSUBS 0.027808f
C474 VTAIL.n20 VSUBS 0.027808f
C475 VTAIL.n21 VSUBS 0.014943f
C476 VTAIL.n22 VSUBS 0.015822f
C477 VTAIL.n23 VSUBS 0.03532f
C478 VTAIL.n24 VSUBS 0.088723f
C479 VTAIL.n25 VSUBS 0.015822f
C480 VTAIL.n26 VSUBS 0.014943f
C481 VTAIL.n27 VSUBS 0.069216f
C482 VTAIL.n28 VSUBS 0.044907f
C483 VTAIL.n29 VSUBS 0.110353f
C484 VTAIL.n30 VSUBS 0.0315f
C485 VTAIL.n31 VSUBS 0.027808f
C486 VTAIL.n32 VSUBS 0.014943f
C487 VTAIL.n33 VSUBS 0.03532f
C488 VTAIL.n34 VSUBS 0.015822f
C489 VTAIL.n35 VSUBS 0.027808f
C490 VTAIL.n36 VSUBS 0.014943f
C491 VTAIL.n37 VSUBS 0.02649f
C492 VTAIL.n38 VSUBS 0.022435f
C493 VTAIL.t5 VSUBS 0.076499f
C494 VTAIL.n39 VSUBS 0.11879f
C495 VTAIL.n40 VSUBS 0.56201f
C496 VTAIL.n41 VSUBS 0.014943f
C497 VTAIL.n42 VSUBS 0.015822f
C498 VTAIL.n43 VSUBS 0.03532f
C499 VTAIL.n44 VSUBS 0.03532f
C500 VTAIL.n45 VSUBS 0.015822f
C501 VTAIL.n46 VSUBS 0.014943f
C502 VTAIL.n47 VSUBS 0.027808f
C503 VTAIL.n48 VSUBS 0.027808f
C504 VTAIL.n49 VSUBS 0.014943f
C505 VTAIL.n50 VSUBS 0.015822f
C506 VTAIL.n51 VSUBS 0.03532f
C507 VTAIL.n52 VSUBS 0.088723f
C508 VTAIL.n53 VSUBS 0.015822f
C509 VTAIL.n54 VSUBS 0.014943f
C510 VTAIL.n55 VSUBS 0.069216f
C511 VTAIL.n56 VSUBS 0.044907f
C512 VTAIL.n57 VSUBS 0.110353f
C513 VTAIL.t7 VSUBS 0.118884f
C514 VTAIL.t2 VSUBS 0.118884f
C515 VTAIL.n58 VSUBS 0.680844f
C516 VTAIL.n59 VSUBS 0.566741f
C517 VTAIL.n60 VSUBS 0.0315f
C518 VTAIL.n61 VSUBS 0.027808f
C519 VTAIL.n62 VSUBS 0.014943f
C520 VTAIL.n63 VSUBS 0.03532f
C521 VTAIL.n64 VSUBS 0.015822f
C522 VTAIL.n65 VSUBS 0.027808f
C523 VTAIL.n66 VSUBS 0.014943f
C524 VTAIL.n67 VSUBS 0.02649f
C525 VTAIL.n68 VSUBS 0.022435f
C526 VTAIL.t6 VSUBS 0.076499f
C527 VTAIL.n69 VSUBS 0.11879f
C528 VTAIL.n70 VSUBS 0.56201f
C529 VTAIL.n71 VSUBS 0.014943f
C530 VTAIL.n72 VSUBS 0.015822f
C531 VTAIL.n73 VSUBS 0.03532f
C532 VTAIL.n74 VSUBS 0.03532f
C533 VTAIL.n75 VSUBS 0.015822f
C534 VTAIL.n76 VSUBS 0.014943f
C535 VTAIL.n77 VSUBS 0.027808f
C536 VTAIL.n78 VSUBS 0.027808f
C537 VTAIL.n79 VSUBS 0.014943f
C538 VTAIL.n80 VSUBS 0.015822f
C539 VTAIL.n81 VSUBS 0.03532f
C540 VTAIL.n82 VSUBS 0.088723f
C541 VTAIL.n83 VSUBS 0.015822f
C542 VTAIL.n84 VSUBS 0.014943f
C543 VTAIL.n85 VSUBS 0.069216f
C544 VTAIL.n86 VSUBS 0.044907f
C545 VTAIL.n87 VSUBS 0.905603f
C546 VTAIL.n88 VSUBS 0.0315f
C547 VTAIL.n89 VSUBS 0.027808f
C548 VTAIL.n90 VSUBS 0.014943f
C549 VTAIL.n91 VSUBS 0.03532f
C550 VTAIL.n92 VSUBS 0.015822f
C551 VTAIL.n93 VSUBS 0.027808f
C552 VTAIL.n94 VSUBS 0.014943f
C553 VTAIL.n95 VSUBS 0.02649f
C554 VTAIL.n96 VSUBS 0.022435f
C555 VTAIL.t8 VSUBS 0.076499f
C556 VTAIL.n97 VSUBS 0.11879f
C557 VTAIL.n98 VSUBS 0.56201f
C558 VTAIL.n99 VSUBS 0.014943f
C559 VTAIL.n100 VSUBS 0.015822f
C560 VTAIL.n101 VSUBS 0.03532f
C561 VTAIL.n102 VSUBS 0.03532f
C562 VTAIL.n103 VSUBS 0.015822f
C563 VTAIL.n104 VSUBS 0.014943f
C564 VTAIL.n105 VSUBS 0.027808f
C565 VTAIL.n106 VSUBS 0.027808f
C566 VTAIL.n107 VSUBS 0.014943f
C567 VTAIL.n108 VSUBS 0.015822f
C568 VTAIL.n109 VSUBS 0.03532f
C569 VTAIL.n110 VSUBS 0.088723f
C570 VTAIL.n111 VSUBS 0.015822f
C571 VTAIL.n112 VSUBS 0.014943f
C572 VTAIL.n113 VSUBS 0.069216f
C573 VTAIL.n114 VSUBS 0.044907f
C574 VTAIL.n115 VSUBS 0.905603f
C575 VTAIL.t10 VSUBS 0.118884f
C576 VTAIL.t12 VSUBS 0.118884f
C577 VTAIL.n116 VSUBS 0.680849f
C578 VTAIL.n117 VSUBS 0.566736f
C579 VTAIL.n118 VSUBS 0.0315f
C580 VTAIL.n119 VSUBS 0.027808f
C581 VTAIL.n120 VSUBS 0.014943f
C582 VTAIL.n121 VSUBS 0.03532f
C583 VTAIL.n122 VSUBS 0.015822f
C584 VTAIL.n123 VSUBS 0.027808f
C585 VTAIL.n124 VSUBS 0.014943f
C586 VTAIL.n125 VSUBS 0.02649f
C587 VTAIL.n126 VSUBS 0.022435f
C588 VTAIL.t15 VSUBS 0.076499f
C589 VTAIL.n127 VSUBS 0.11879f
C590 VTAIL.n128 VSUBS 0.56201f
C591 VTAIL.n129 VSUBS 0.014943f
C592 VTAIL.n130 VSUBS 0.015822f
C593 VTAIL.n131 VSUBS 0.03532f
C594 VTAIL.n132 VSUBS 0.03532f
C595 VTAIL.n133 VSUBS 0.015822f
C596 VTAIL.n134 VSUBS 0.014943f
C597 VTAIL.n135 VSUBS 0.027808f
C598 VTAIL.n136 VSUBS 0.027808f
C599 VTAIL.n137 VSUBS 0.014943f
C600 VTAIL.n138 VSUBS 0.015822f
C601 VTAIL.n139 VSUBS 0.03532f
C602 VTAIL.n140 VSUBS 0.088723f
C603 VTAIL.n141 VSUBS 0.015822f
C604 VTAIL.n142 VSUBS 0.014943f
C605 VTAIL.n143 VSUBS 0.069216f
C606 VTAIL.n144 VSUBS 0.044907f
C607 VTAIL.n145 VSUBS 0.110353f
C608 VTAIL.n146 VSUBS 0.0315f
C609 VTAIL.n147 VSUBS 0.027808f
C610 VTAIL.n148 VSUBS 0.014943f
C611 VTAIL.n149 VSUBS 0.03532f
C612 VTAIL.n150 VSUBS 0.015822f
C613 VTAIL.n151 VSUBS 0.027808f
C614 VTAIL.n152 VSUBS 0.014943f
C615 VTAIL.n153 VSUBS 0.02649f
C616 VTAIL.n154 VSUBS 0.022435f
C617 VTAIL.t1 VSUBS 0.076499f
C618 VTAIL.n155 VSUBS 0.11879f
C619 VTAIL.n156 VSUBS 0.56201f
C620 VTAIL.n157 VSUBS 0.014943f
C621 VTAIL.n158 VSUBS 0.015822f
C622 VTAIL.n159 VSUBS 0.03532f
C623 VTAIL.n160 VSUBS 0.03532f
C624 VTAIL.n161 VSUBS 0.015822f
C625 VTAIL.n162 VSUBS 0.014943f
C626 VTAIL.n163 VSUBS 0.027808f
C627 VTAIL.n164 VSUBS 0.027808f
C628 VTAIL.n165 VSUBS 0.014943f
C629 VTAIL.n166 VSUBS 0.015822f
C630 VTAIL.n167 VSUBS 0.03532f
C631 VTAIL.n168 VSUBS 0.088723f
C632 VTAIL.n169 VSUBS 0.015822f
C633 VTAIL.n170 VSUBS 0.014943f
C634 VTAIL.n171 VSUBS 0.069216f
C635 VTAIL.n172 VSUBS 0.044907f
C636 VTAIL.n173 VSUBS 0.110353f
C637 VTAIL.t3 VSUBS 0.118884f
C638 VTAIL.t0 VSUBS 0.118884f
C639 VTAIL.n174 VSUBS 0.680849f
C640 VTAIL.n175 VSUBS 0.566736f
C641 VTAIL.n176 VSUBS 0.0315f
C642 VTAIL.n177 VSUBS 0.027808f
C643 VTAIL.n178 VSUBS 0.014943f
C644 VTAIL.n179 VSUBS 0.03532f
C645 VTAIL.n180 VSUBS 0.015822f
C646 VTAIL.n181 VSUBS 0.027808f
C647 VTAIL.n182 VSUBS 0.014943f
C648 VTAIL.n183 VSUBS 0.02649f
C649 VTAIL.n184 VSUBS 0.022435f
C650 VTAIL.t4 VSUBS 0.076499f
C651 VTAIL.n185 VSUBS 0.11879f
C652 VTAIL.n186 VSUBS 0.56201f
C653 VTAIL.n187 VSUBS 0.014943f
C654 VTAIL.n188 VSUBS 0.015822f
C655 VTAIL.n189 VSUBS 0.03532f
C656 VTAIL.n190 VSUBS 0.03532f
C657 VTAIL.n191 VSUBS 0.015822f
C658 VTAIL.n192 VSUBS 0.014943f
C659 VTAIL.n193 VSUBS 0.027808f
C660 VTAIL.n194 VSUBS 0.027808f
C661 VTAIL.n195 VSUBS 0.014943f
C662 VTAIL.n196 VSUBS 0.015822f
C663 VTAIL.n197 VSUBS 0.03532f
C664 VTAIL.n198 VSUBS 0.088723f
C665 VTAIL.n199 VSUBS 0.015822f
C666 VTAIL.n200 VSUBS 0.014943f
C667 VTAIL.n201 VSUBS 0.069216f
C668 VTAIL.n202 VSUBS 0.044907f
C669 VTAIL.n203 VSUBS 0.905602f
C670 VTAIL.n204 VSUBS 0.0315f
C671 VTAIL.n205 VSUBS 0.027808f
C672 VTAIL.n206 VSUBS 0.014943f
C673 VTAIL.n207 VSUBS 0.03532f
C674 VTAIL.n208 VSUBS 0.015822f
C675 VTAIL.n209 VSUBS 0.027808f
C676 VTAIL.n210 VSUBS 0.014943f
C677 VTAIL.n211 VSUBS 0.02649f
C678 VTAIL.n212 VSUBS 0.022435f
C679 VTAIL.t13 VSUBS 0.076499f
C680 VTAIL.n213 VSUBS 0.11879f
C681 VTAIL.n214 VSUBS 0.56201f
C682 VTAIL.n215 VSUBS 0.014943f
C683 VTAIL.n216 VSUBS 0.015822f
C684 VTAIL.n217 VSUBS 0.03532f
C685 VTAIL.n218 VSUBS 0.03532f
C686 VTAIL.n219 VSUBS 0.015822f
C687 VTAIL.n220 VSUBS 0.014943f
C688 VTAIL.n221 VSUBS 0.027808f
C689 VTAIL.n222 VSUBS 0.027808f
C690 VTAIL.n223 VSUBS 0.014943f
C691 VTAIL.n224 VSUBS 0.015822f
C692 VTAIL.n225 VSUBS 0.03532f
C693 VTAIL.n226 VSUBS 0.088723f
C694 VTAIL.n227 VSUBS 0.015822f
C695 VTAIL.n228 VSUBS 0.014943f
C696 VTAIL.n229 VSUBS 0.069216f
C697 VTAIL.n230 VSUBS 0.044907f
C698 VTAIL.n231 VSUBS 0.900389f
C699 VN.n0 VSUBS 0.119471f
C700 VN.t2 VSUBS 0.176039f
C701 VN.t7 VSUBS 0.176039f
C702 VN.t5 VSUBS 0.18097f
C703 VN.n1 VSUBS 0.103398f
C704 VN.n2 VSUBS 0.088248f
C705 VN.n3 VSUBS 0.019336f
C706 VN.n4 VSUBS 0.088248f
C707 VN.t0 VSUBS 0.18097f
C708 VN.n5 VSUBS 0.103322f
C709 VN.n6 VSUBS 0.042045f
C710 VN.n7 VSUBS 0.119471f
C711 VN.t6 VSUBS 0.18097f
C712 VN.t4 VSUBS 0.176039f
C713 VN.t3 VSUBS 0.176039f
C714 VN.t1 VSUBS 0.18097f
C715 VN.n8 VSUBS 0.103398f
C716 VN.n9 VSUBS 0.088248f
C717 VN.n10 VSUBS 0.019336f
C718 VN.n11 VSUBS 0.088248f
C719 VN.n12 VSUBS 0.103322f
C720 VN.n13 VSUBS 1.63387f
.ends

