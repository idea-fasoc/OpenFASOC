* NGSPICE file created from diff_pair_sample_1392.ext - technology: sky130A

.subckt diff_pair_sample_1392 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=2.4552 pd=15.21 as=2.4552 ps=15.21 w=14.88 l=0.58
X1 VDD1.t5 VP.t1 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=5.8032 pd=30.54 as=2.4552 ps=15.21 w=14.88 l=0.58
X2 VDD2.t5 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=5.8032 pd=30.54 as=2.4552 ps=15.21 w=14.88 l=0.58
X3 VTAIL.t1 VN.t1 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.4552 pd=15.21 as=2.4552 ps=15.21 w=14.88 l=0.58
X4 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=5.8032 pd=30.54 as=0 ps=0 w=14.88 l=0.58
X5 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=5.8032 pd=30.54 as=0 ps=0 w=14.88 l=0.58
X6 VTAIL.t9 VP.t2 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.4552 pd=15.21 as=2.4552 ps=15.21 w=14.88 l=0.58
X7 VDD1.t1 VP.t3 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=2.4552 pd=15.21 as=5.8032 ps=30.54 w=14.88 l=0.58
X8 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=5.8032 pd=30.54 as=0 ps=0 w=14.88 l=0.58
X9 VDD2.t3 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=5.8032 pd=30.54 as=2.4552 ps=15.21 w=14.88 l=0.58
X10 VDD1.t2 VP.t4 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=2.4552 pd=15.21 as=5.8032 ps=30.54 w=14.88 l=0.58
X11 VDD2.t2 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.4552 pd=15.21 as=5.8032 ps=30.54 w=14.88 l=0.58
X12 VDD2.t1 VN.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.4552 pd=15.21 as=5.8032 ps=30.54 w=14.88 l=0.58
X13 VDD1.t4 VP.t5 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=5.8032 pd=30.54 as=2.4552 ps=15.21 w=14.88 l=0.58
X14 VTAIL.t4 VN.t5 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=2.4552 pd=15.21 as=2.4552 ps=15.21 w=14.88 l=0.58
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.8032 pd=30.54 as=0 ps=0 w=14.88 l=0.58
R0 VP.n1 VP.t1 712.841
R1 VP.n6 VP.t5 686.019
R2 VP.n7 VP.t0 686.019
R3 VP.n8 VP.t3 686.019
R4 VP.n3 VP.t4 686.019
R5 VP.n2 VP.t2 686.019
R6 VP.n9 VP.n8 161.3
R7 VP.n4 VP.n3 161.3
R8 VP.n6 VP.n5 161.3
R9 VP.n7 VP.n0 80.6037
R10 VP.n7 VP.n6 48.2005
R11 VP.n8 VP.n7 48.2005
R12 VP.n3 VP.n2 48.2005
R13 VP.n4 VP.n1 45.1367
R14 VP.n5 VP.n4 42.9816
R15 VP.n2 VP.n1 13.3799
R16 VP.n5 VP.n0 0.285035
R17 VP.n9 VP.n0 0.285035
R18 VP VP.n9 0.0516364
R19 VDD1.n76 VDD1.n0 289.615
R20 VDD1.n157 VDD1.n81 289.615
R21 VDD1.n77 VDD1.n76 185
R22 VDD1.n75 VDD1.n74 185
R23 VDD1.n4 VDD1.n3 185
R24 VDD1.n69 VDD1.n68 185
R25 VDD1.n67 VDD1.n66 185
R26 VDD1.n8 VDD1.n7 185
R27 VDD1.n61 VDD1.n60 185
R28 VDD1.n59 VDD1.n58 185
R29 VDD1.n12 VDD1.n11 185
R30 VDD1.n53 VDD1.n52 185
R31 VDD1.n51 VDD1.n50 185
R32 VDD1.n49 VDD1.n15 185
R33 VDD1.n19 VDD1.n16 185
R34 VDD1.n44 VDD1.n43 185
R35 VDD1.n42 VDD1.n41 185
R36 VDD1.n21 VDD1.n20 185
R37 VDD1.n36 VDD1.n35 185
R38 VDD1.n34 VDD1.n33 185
R39 VDD1.n25 VDD1.n24 185
R40 VDD1.n28 VDD1.n27 185
R41 VDD1.n108 VDD1.n107 185
R42 VDD1.n105 VDD1.n104 185
R43 VDD1.n114 VDD1.n113 185
R44 VDD1.n116 VDD1.n115 185
R45 VDD1.n101 VDD1.n100 185
R46 VDD1.n122 VDD1.n121 185
R47 VDD1.n125 VDD1.n124 185
R48 VDD1.n123 VDD1.n97 185
R49 VDD1.n130 VDD1.n96 185
R50 VDD1.n132 VDD1.n131 185
R51 VDD1.n134 VDD1.n133 185
R52 VDD1.n93 VDD1.n92 185
R53 VDD1.n140 VDD1.n139 185
R54 VDD1.n142 VDD1.n141 185
R55 VDD1.n89 VDD1.n88 185
R56 VDD1.n148 VDD1.n147 185
R57 VDD1.n150 VDD1.n149 185
R58 VDD1.n85 VDD1.n84 185
R59 VDD1.n156 VDD1.n155 185
R60 VDD1.n158 VDD1.n157 185
R61 VDD1.t5 VDD1.n26 149.524
R62 VDD1.t4 VDD1.n106 149.524
R63 VDD1.n76 VDD1.n75 104.615
R64 VDD1.n75 VDD1.n3 104.615
R65 VDD1.n68 VDD1.n3 104.615
R66 VDD1.n68 VDD1.n67 104.615
R67 VDD1.n67 VDD1.n7 104.615
R68 VDD1.n60 VDD1.n7 104.615
R69 VDD1.n60 VDD1.n59 104.615
R70 VDD1.n59 VDD1.n11 104.615
R71 VDD1.n52 VDD1.n11 104.615
R72 VDD1.n52 VDD1.n51 104.615
R73 VDD1.n51 VDD1.n15 104.615
R74 VDD1.n19 VDD1.n15 104.615
R75 VDD1.n43 VDD1.n19 104.615
R76 VDD1.n43 VDD1.n42 104.615
R77 VDD1.n42 VDD1.n20 104.615
R78 VDD1.n35 VDD1.n20 104.615
R79 VDD1.n35 VDD1.n34 104.615
R80 VDD1.n34 VDD1.n24 104.615
R81 VDD1.n27 VDD1.n24 104.615
R82 VDD1.n107 VDD1.n104 104.615
R83 VDD1.n114 VDD1.n104 104.615
R84 VDD1.n115 VDD1.n114 104.615
R85 VDD1.n115 VDD1.n100 104.615
R86 VDD1.n122 VDD1.n100 104.615
R87 VDD1.n124 VDD1.n122 104.615
R88 VDD1.n124 VDD1.n123 104.615
R89 VDD1.n123 VDD1.n96 104.615
R90 VDD1.n132 VDD1.n96 104.615
R91 VDD1.n133 VDD1.n132 104.615
R92 VDD1.n133 VDD1.n92 104.615
R93 VDD1.n140 VDD1.n92 104.615
R94 VDD1.n141 VDD1.n140 104.615
R95 VDD1.n141 VDD1.n88 104.615
R96 VDD1.n148 VDD1.n88 104.615
R97 VDD1.n149 VDD1.n148 104.615
R98 VDD1.n149 VDD1.n84 104.615
R99 VDD1.n156 VDD1.n84 104.615
R100 VDD1.n157 VDD1.n156 104.615
R101 VDD1.n163 VDD1.n162 59.135
R102 VDD1.n165 VDD1.n164 58.9944
R103 VDD1.n27 VDD1.t5 52.3082
R104 VDD1.n107 VDD1.t4 52.3082
R105 VDD1 VDD1.n80 47.1834
R106 VDD1.n163 VDD1.n161 47.0699
R107 VDD1.n165 VDD1.n163 40.0677
R108 VDD1.n50 VDD1.n49 13.1884
R109 VDD1.n131 VDD1.n130 13.1884
R110 VDD1.n53 VDD1.n14 12.8005
R111 VDD1.n48 VDD1.n16 12.8005
R112 VDD1.n129 VDD1.n97 12.8005
R113 VDD1.n134 VDD1.n95 12.8005
R114 VDD1.n54 VDD1.n12 12.0247
R115 VDD1.n45 VDD1.n44 12.0247
R116 VDD1.n126 VDD1.n125 12.0247
R117 VDD1.n135 VDD1.n93 12.0247
R118 VDD1.n58 VDD1.n57 11.249
R119 VDD1.n41 VDD1.n18 11.249
R120 VDD1.n121 VDD1.n99 11.249
R121 VDD1.n139 VDD1.n138 11.249
R122 VDD1.n61 VDD1.n10 10.4732
R123 VDD1.n40 VDD1.n21 10.4732
R124 VDD1.n120 VDD1.n101 10.4732
R125 VDD1.n142 VDD1.n91 10.4732
R126 VDD1.n28 VDD1.n26 10.2747
R127 VDD1.n108 VDD1.n106 10.2747
R128 VDD1.n62 VDD1.n8 9.69747
R129 VDD1.n37 VDD1.n36 9.69747
R130 VDD1.n117 VDD1.n116 9.69747
R131 VDD1.n143 VDD1.n89 9.69747
R132 VDD1.n80 VDD1.n79 9.45567
R133 VDD1.n161 VDD1.n160 9.45567
R134 VDD1.n30 VDD1.n29 9.3005
R135 VDD1.n32 VDD1.n31 9.3005
R136 VDD1.n23 VDD1.n22 9.3005
R137 VDD1.n38 VDD1.n37 9.3005
R138 VDD1.n40 VDD1.n39 9.3005
R139 VDD1.n18 VDD1.n17 9.3005
R140 VDD1.n46 VDD1.n45 9.3005
R141 VDD1.n48 VDD1.n47 9.3005
R142 VDD1.n2 VDD1.n1 9.3005
R143 VDD1.n79 VDD1.n78 9.3005
R144 VDD1.n73 VDD1.n72 9.3005
R145 VDD1.n71 VDD1.n70 9.3005
R146 VDD1.n6 VDD1.n5 9.3005
R147 VDD1.n65 VDD1.n64 9.3005
R148 VDD1.n63 VDD1.n62 9.3005
R149 VDD1.n10 VDD1.n9 9.3005
R150 VDD1.n57 VDD1.n56 9.3005
R151 VDD1.n55 VDD1.n54 9.3005
R152 VDD1.n14 VDD1.n13 9.3005
R153 VDD1.n154 VDD1.n153 9.3005
R154 VDD1.n83 VDD1.n82 9.3005
R155 VDD1.n160 VDD1.n159 9.3005
R156 VDD1.n87 VDD1.n86 9.3005
R157 VDD1.n146 VDD1.n145 9.3005
R158 VDD1.n144 VDD1.n143 9.3005
R159 VDD1.n91 VDD1.n90 9.3005
R160 VDD1.n138 VDD1.n137 9.3005
R161 VDD1.n136 VDD1.n135 9.3005
R162 VDD1.n95 VDD1.n94 9.3005
R163 VDD1.n110 VDD1.n109 9.3005
R164 VDD1.n112 VDD1.n111 9.3005
R165 VDD1.n103 VDD1.n102 9.3005
R166 VDD1.n118 VDD1.n117 9.3005
R167 VDD1.n120 VDD1.n119 9.3005
R168 VDD1.n99 VDD1.n98 9.3005
R169 VDD1.n127 VDD1.n126 9.3005
R170 VDD1.n129 VDD1.n128 9.3005
R171 VDD1.n152 VDD1.n151 9.3005
R172 VDD1.n80 VDD1.n0 8.92171
R173 VDD1.n66 VDD1.n65 8.92171
R174 VDD1.n33 VDD1.n23 8.92171
R175 VDD1.n113 VDD1.n103 8.92171
R176 VDD1.n147 VDD1.n146 8.92171
R177 VDD1.n161 VDD1.n81 8.92171
R178 VDD1.n78 VDD1.n77 8.14595
R179 VDD1.n69 VDD1.n6 8.14595
R180 VDD1.n32 VDD1.n25 8.14595
R181 VDD1.n112 VDD1.n105 8.14595
R182 VDD1.n150 VDD1.n87 8.14595
R183 VDD1.n159 VDD1.n158 8.14595
R184 VDD1.n74 VDD1.n2 7.3702
R185 VDD1.n70 VDD1.n4 7.3702
R186 VDD1.n29 VDD1.n28 7.3702
R187 VDD1.n109 VDD1.n108 7.3702
R188 VDD1.n151 VDD1.n85 7.3702
R189 VDD1.n155 VDD1.n83 7.3702
R190 VDD1.n74 VDD1.n73 6.59444
R191 VDD1.n73 VDD1.n4 6.59444
R192 VDD1.n154 VDD1.n85 6.59444
R193 VDD1.n155 VDD1.n154 6.59444
R194 VDD1.n77 VDD1.n2 5.81868
R195 VDD1.n70 VDD1.n69 5.81868
R196 VDD1.n29 VDD1.n25 5.81868
R197 VDD1.n109 VDD1.n105 5.81868
R198 VDD1.n151 VDD1.n150 5.81868
R199 VDD1.n158 VDD1.n83 5.81868
R200 VDD1.n78 VDD1.n0 5.04292
R201 VDD1.n66 VDD1.n6 5.04292
R202 VDD1.n33 VDD1.n32 5.04292
R203 VDD1.n113 VDD1.n112 5.04292
R204 VDD1.n147 VDD1.n87 5.04292
R205 VDD1.n159 VDD1.n81 5.04292
R206 VDD1.n65 VDD1.n8 4.26717
R207 VDD1.n36 VDD1.n23 4.26717
R208 VDD1.n116 VDD1.n103 4.26717
R209 VDD1.n146 VDD1.n89 4.26717
R210 VDD1.n62 VDD1.n61 3.49141
R211 VDD1.n37 VDD1.n21 3.49141
R212 VDD1.n117 VDD1.n101 3.49141
R213 VDD1.n143 VDD1.n142 3.49141
R214 VDD1.n110 VDD1.n106 2.84303
R215 VDD1.n30 VDD1.n26 2.84303
R216 VDD1.n58 VDD1.n10 2.71565
R217 VDD1.n41 VDD1.n40 2.71565
R218 VDD1.n121 VDD1.n120 2.71565
R219 VDD1.n139 VDD1.n91 2.71565
R220 VDD1.n57 VDD1.n12 1.93989
R221 VDD1.n44 VDD1.n18 1.93989
R222 VDD1.n125 VDD1.n99 1.93989
R223 VDD1.n138 VDD1.n93 1.93989
R224 VDD1.n164 VDD1.t0 1.33115
R225 VDD1.n164 VDD1.t2 1.33115
R226 VDD1.n162 VDD1.t3 1.33115
R227 VDD1.n162 VDD1.t1 1.33115
R228 VDD1.n54 VDD1.n53 1.16414
R229 VDD1.n45 VDD1.n16 1.16414
R230 VDD1.n126 VDD1.n97 1.16414
R231 VDD1.n135 VDD1.n134 1.16414
R232 VDD1.n50 VDD1.n14 0.388379
R233 VDD1.n49 VDD1.n48 0.388379
R234 VDD1.n130 VDD1.n129 0.388379
R235 VDD1.n131 VDD1.n95 0.388379
R236 VDD1.n79 VDD1.n1 0.155672
R237 VDD1.n72 VDD1.n1 0.155672
R238 VDD1.n72 VDD1.n71 0.155672
R239 VDD1.n71 VDD1.n5 0.155672
R240 VDD1.n64 VDD1.n5 0.155672
R241 VDD1.n64 VDD1.n63 0.155672
R242 VDD1.n63 VDD1.n9 0.155672
R243 VDD1.n56 VDD1.n9 0.155672
R244 VDD1.n56 VDD1.n55 0.155672
R245 VDD1.n55 VDD1.n13 0.155672
R246 VDD1.n47 VDD1.n13 0.155672
R247 VDD1.n47 VDD1.n46 0.155672
R248 VDD1.n46 VDD1.n17 0.155672
R249 VDD1.n39 VDD1.n17 0.155672
R250 VDD1.n39 VDD1.n38 0.155672
R251 VDD1.n38 VDD1.n22 0.155672
R252 VDD1.n31 VDD1.n22 0.155672
R253 VDD1.n31 VDD1.n30 0.155672
R254 VDD1.n111 VDD1.n110 0.155672
R255 VDD1.n111 VDD1.n102 0.155672
R256 VDD1.n118 VDD1.n102 0.155672
R257 VDD1.n119 VDD1.n118 0.155672
R258 VDD1.n119 VDD1.n98 0.155672
R259 VDD1.n127 VDD1.n98 0.155672
R260 VDD1.n128 VDD1.n127 0.155672
R261 VDD1.n128 VDD1.n94 0.155672
R262 VDD1.n136 VDD1.n94 0.155672
R263 VDD1.n137 VDD1.n136 0.155672
R264 VDD1.n137 VDD1.n90 0.155672
R265 VDD1.n144 VDD1.n90 0.155672
R266 VDD1.n145 VDD1.n144 0.155672
R267 VDD1.n145 VDD1.n86 0.155672
R268 VDD1.n152 VDD1.n86 0.155672
R269 VDD1.n153 VDD1.n152 0.155672
R270 VDD1.n153 VDD1.n82 0.155672
R271 VDD1.n160 VDD1.n82 0.155672
R272 VDD1 VDD1.n165 0.138431
R273 VTAIL.n330 VTAIL.n254 289.615
R274 VTAIL.n78 VTAIL.n2 289.615
R275 VTAIL.n248 VTAIL.n172 289.615
R276 VTAIL.n164 VTAIL.n88 289.615
R277 VTAIL.n281 VTAIL.n280 185
R278 VTAIL.n278 VTAIL.n277 185
R279 VTAIL.n287 VTAIL.n286 185
R280 VTAIL.n289 VTAIL.n288 185
R281 VTAIL.n274 VTAIL.n273 185
R282 VTAIL.n295 VTAIL.n294 185
R283 VTAIL.n298 VTAIL.n297 185
R284 VTAIL.n296 VTAIL.n270 185
R285 VTAIL.n303 VTAIL.n269 185
R286 VTAIL.n305 VTAIL.n304 185
R287 VTAIL.n307 VTAIL.n306 185
R288 VTAIL.n266 VTAIL.n265 185
R289 VTAIL.n313 VTAIL.n312 185
R290 VTAIL.n315 VTAIL.n314 185
R291 VTAIL.n262 VTAIL.n261 185
R292 VTAIL.n321 VTAIL.n320 185
R293 VTAIL.n323 VTAIL.n322 185
R294 VTAIL.n258 VTAIL.n257 185
R295 VTAIL.n329 VTAIL.n328 185
R296 VTAIL.n331 VTAIL.n330 185
R297 VTAIL.n29 VTAIL.n28 185
R298 VTAIL.n26 VTAIL.n25 185
R299 VTAIL.n35 VTAIL.n34 185
R300 VTAIL.n37 VTAIL.n36 185
R301 VTAIL.n22 VTAIL.n21 185
R302 VTAIL.n43 VTAIL.n42 185
R303 VTAIL.n46 VTAIL.n45 185
R304 VTAIL.n44 VTAIL.n18 185
R305 VTAIL.n51 VTAIL.n17 185
R306 VTAIL.n53 VTAIL.n52 185
R307 VTAIL.n55 VTAIL.n54 185
R308 VTAIL.n14 VTAIL.n13 185
R309 VTAIL.n61 VTAIL.n60 185
R310 VTAIL.n63 VTAIL.n62 185
R311 VTAIL.n10 VTAIL.n9 185
R312 VTAIL.n69 VTAIL.n68 185
R313 VTAIL.n71 VTAIL.n70 185
R314 VTAIL.n6 VTAIL.n5 185
R315 VTAIL.n77 VTAIL.n76 185
R316 VTAIL.n79 VTAIL.n78 185
R317 VTAIL.n249 VTAIL.n248 185
R318 VTAIL.n247 VTAIL.n246 185
R319 VTAIL.n176 VTAIL.n175 185
R320 VTAIL.n241 VTAIL.n240 185
R321 VTAIL.n239 VTAIL.n238 185
R322 VTAIL.n180 VTAIL.n179 185
R323 VTAIL.n233 VTAIL.n232 185
R324 VTAIL.n231 VTAIL.n230 185
R325 VTAIL.n184 VTAIL.n183 185
R326 VTAIL.n225 VTAIL.n224 185
R327 VTAIL.n223 VTAIL.n222 185
R328 VTAIL.n221 VTAIL.n187 185
R329 VTAIL.n191 VTAIL.n188 185
R330 VTAIL.n216 VTAIL.n215 185
R331 VTAIL.n214 VTAIL.n213 185
R332 VTAIL.n193 VTAIL.n192 185
R333 VTAIL.n208 VTAIL.n207 185
R334 VTAIL.n206 VTAIL.n205 185
R335 VTAIL.n197 VTAIL.n196 185
R336 VTAIL.n200 VTAIL.n199 185
R337 VTAIL.n165 VTAIL.n164 185
R338 VTAIL.n163 VTAIL.n162 185
R339 VTAIL.n92 VTAIL.n91 185
R340 VTAIL.n157 VTAIL.n156 185
R341 VTAIL.n155 VTAIL.n154 185
R342 VTAIL.n96 VTAIL.n95 185
R343 VTAIL.n149 VTAIL.n148 185
R344 VTAIL.n147 VTAIL.n146 185
R345 VTAIL.n100 VTAIL.n99 185
R346 VTAIL.n141 VTAIL.n140 185
R347 VTAIL.n139 VTAIL.n138 185
R348 VTAIL.n137 VTAIL.n103 185
R349 VTAIL.n107 VTAIL.n104 185
R350 VTAIL.n132 VTAIL.n131 185
R351 VTAIL.n130 VTAIL.n129 185
R352 VTAIL.n109 VTAIL.n108 185
R353 VTAIL.n124 VTAIL.n123 185
R354 VTAIL.n122 VTAIL.n121 185
R355 VTAIL.n113 VTAIL.n112 185
R356 VTAIL.n116 VTAIL.n115 185
R357 VTAIL.t5 VTAIL.n279 149.524
R358 VTAIL.t8 VTAIL.n27 149.524
R359 VTAIL.t7 VTAIL.n198 149.524
R360 VTAIL.t0 VTAIL.n114 149.524
R361 VTAIL.n280 VTAIL.n277 104.615
R362 VTAIL.n287 VTAIL.n277 104.615
R363 VTAIL.n288 VTAIL.n287 104.615
R364 VTAIL.n288 VTAIL.n273 104.615
R365 VTAIL.n295 VTAIL.n273 104.615
R366 VTAIL.n297 VTAIL.n295 104.615
R367 VTAIL.n297 VTAIL.n296 104.615
R368 VTAIL.n296 VTAIL.n269 104.615
R369 VTAIL.n305 VTAIL.n269 104.615
R370 VTAIL.n306 VTAIL.n305 104.615
R371 VTAIL.n306 VTAIL.n265 104.615
R372 VTAIL.n313 VTAIL.n265 104.615
R373 VTAIL.n314 VTAIL.n313 104.615
R374 VTAIL.n314 VTAIL.n261 104.615
R375 VTAIL.n321 VTAIL.n261 104.615
R376 VTAIL.n322 VTAIL.n321 104.615
R377 VTAIL.n322 VTAIL.n257 104.615
R378 VTAIL.n329 VTAIL.n257 104.615
R379 VTAIL.n330 VTAIL.n329 104.615
R380 VTAIL.n28 VTAIL.n25 104.615
R381 VTAIL.n35 VTAIL.n25 104.615
R382 VTAIL.n36 VTAIL.n35 104.615
R383 VTAIL.n36 VTAIL.n21 104.615
R384 VTAIL.n43 VTAIL.n21 104.615
R385 VTAIL.n45 VTAIL.n43 104.615
R386 VTAIL.n45 VTAIL.n44 104.615
R387 VTAIL.n44 VTAIL.n17 104.615
R388 VTAIL.n53 VTAIL.n17 104.615
R389 VTAIL.n54 VTAIL.n53 104.615
R390 VTAIL.n54 VTAIL.n13 104.615
R391 VTAIL.n61 VTAIL.n13 104.615
R392 VTAIL.n62 VTAIL.n61 104.615
R393 VTAIL.n62 VTAIL.n9 104.615
R394 VTAIL.n69 VTAIL.n9 104.615
R395 VTAIL.n70 VTAIL.n69 104.615
R396 VTAIL.n70 VTAIL.n5 104.615
R397 VTAIL.n77 VTAIL.n5 104.615
R398 VTAIL.n78 VTAIL.n77 104.615
R399 VTAIL.n248 VTAIL.n247 104.615
R400 VTAIL.n247 VTAIL.n175 104.615
R401 VTAIL.n240 VTAIL.n175 104.615
R402 VTAIL.n240 VTAIL.n239 104.615
R403 VTAIL.n239 VTAIL.n179 104.615
R404 VTAIL.n232 VTAIL.n179 104.615
R405 VTAIL.n232 VTAIL.n231 104.615
R406 VTAIL.n231 VTAIL.n183 104.615
R407 VTAIL.n224 VTAIL.n183 104.615
R408 VTAIL.n224 VTAIL.n223 104.615
R409 VTAIL.n223 VTAIL.n187 104.615
R410 VTAIL.n191 VTAIL.n187 104.615
R411 VTAIL.n215 VTAIL.n191 104.615
R412 VTAIL.n215 VTAIL.n214 104.615
R413 VTAIL.n214 VTAIL.n192 104.615
R414 VTAIL.n207 VTAIL.n192 104.615
R415 VTAIL.n207 VTAIL.n206 104.615
R416 VTAIL.n206 VTAIL.n196 104.615
R417 VTAIL.n199 VTAIL.n196 104.615
R418 VTAIL.n164 VTAIL.n163 104.615
R419 VTAIL.n163 VTAIL.n91 104.615
R420 VTAIL.n156 VTAIL.n91 104.615
R421 VTAIL.n156 VTAIL.n155 104.615
R422 VTAIL.n155 VTAIL.n95 104.615
R423 VTAIL.n148 VTAIL.n95 104.615
R424 VTAIL.n148 VTAIL.n147 104.615
R425 VTAIL.n147 VTAIL.n99 104.615
R426 VTAIL.n140 VTAIL.n99 104.615
R427 VTAIL.n140 VTAIL.n139 104.615
R428 VTAIL.n139 VTAIL.n103 104.615
R429 VTAIL.n107 VTAIL.n103 104.615
R430 VTAIL.n131 VTAIL.n107 104.615
R431 VTAIL.n131 VTAIL.n130 104.615
R432 VTAIL.n130 VTAIL.n108 104.615
R433 VTAIL.n123 VTAIL.n108 104.615
R434 VTAIL.n123 VTAIL.n122 104.615
R435 VTAIL.n122 VTAIL.n112 104.615
R436 VTAIL.n115 VTAIL.n112 104.615
R437 VTAIL.n280 VTAIL.t5 52.3082
R438 VTAIL.n28 VTAIL.t8 52.3082
R439 VTAIL.n199 VTAIL.t7 52.3082
R440 VTAIL.n115 VTAIL.t0 52.3082
R441 VTAIL.n171 VTAIL.n170 42.3156
R442 VTAIL.n87 VTAIL.n86 42.3156
R443 VTAIL.n1 VTAIL.n0 42.3154
R444 VTAIL.n85 VTAIL.n84 42.3154
R445 VTAIL.n335 VTAIL.n334 29.8581
R446 VTAIL.n83 VTAIL.n82 29.8581
R447 VTAIL.n253 VTAIL.n252 29.8581
R448 VTAIL.n169 VTAIL.n168 29.8581
R449 VTAIL.n87 VTAIL.n85 26.7634
R450 VTAIL.n335 VTAIL.n253 25.9789
R451 VTAIL.n304 VTAIL.n303 13.1884
R452 VTAIL.n52 VTAIL.n51 13.1884
R453 VTAIL.n222 VTAIL.n221 13.1884
R454 VTAIL.n138 VTAIL.n137 13.1884
R455 VTAIL.n302 VTAIL.n270 12.8005
R456 VTAIL.n307 VTAIL.n268 12.8005
R457 VTAIL.n50 VTAIL.n18 12.8005
R458 VTAIL.n55 VTAIL.n16 12.8005
R459 VTAIL.n225 VTAIL.n186 12.8005
R460 VTAIL.n220 VTAIL.n188 12.8005
R461 VTAIL.n141 VTAIL.n102 12.8005
R462 VTAIL.n136 VTAIL.n104 12.8005
R463 VTAIL.n299 VTAIL.n298 12.0247
R464 VTAIL.n308 VTAIL.n266 12.0247
R465 VTAIL.n47 VTAIL.n46 12.0247
R466 VTAIL.n56 VTAIL.n14 12.0247
R467 VTAIL.n226 VTAIL.n184 12.0247
R468 VTAIL.n217 VTAIL.n216 12.0247
R469 VTAIL.n142 VTAIL.n100 12.0247
R470 VTAIL.n133 VTAIL.n132 12.0247
R471 VTAIL.n294 VTAIL.n272 11.249
R472 VTAIL.n312 VTAIL.n311 11.249
R473 VTAIL.n42 VTAIL.n20 11.249
R474 VTAIL.n60 VTAIL.n59 11.249
R475 VTAIL.n230 VTAIL.n229 11.249
R476 VTAIL.n213 VTAIL.n190 11.249
R477 VTAIL.n146 VTAIL.n145 11.249
R478 VTAIL.n129 VTAIL.n106 11.249
R479 VTAIL.n293 VTAIL.n274 10.4732
R480 VTAIL.n315 VTAIL.n264 10.4732
R481 VTAIL.n41 VTAIL.n22 10.4732
R482 VTAIL.n63 VTAIL.n12 10.4732
R483 VTAIL.n233 VTAIL.n182 10.4732
R484 VTAIL.n212 VTAIL.n193 10.4732
R485 VTAIL.n149 VTAIL.n98 10.4732
R486 VTAIL.n128 VTAIL.n109 10.4732
R487 VTAIL.n281 VTAIL.n279 10.2747
R488 VTAIL.n29 VTAIL.n27 10.2747
R489 VTAIL.n200 VTAIL.n198 10.2747
R490 VTAIL.n116 VTAIL.n114 10.2747
R491 VTAIL.n290 VTAIL.n289 9.69747
R492 VTAIL.n316 VTAIL.n262 9.69747
R493 VTAIL.n38 VTAIL.n37 9.69747
R494 VTAIL.n64 VTAIL.n10 9.69747
R495 VTAIL.n234 VTAIL.n180 9.69747
R496 VTAIL.n209 VTAIL.n208 9.69747
R497 VTAIL.n150 VTAIL.n96 9.69747
R498 VTAIL.n125 VTAIL.n124 9.69747
R499 VTAIL.n334 VTAIL.n333 9.45567
R500 VTAIL.n82 VTAIL.n81 9.45567
R501 VTAIL.n252 VTAIL.n251 9.45567
R502 VTAIL.n168 VTAIL.n167 9.45567
R503 VTAIL.n327 VTAIL.n326 9.3005
R504 VTAIL.n256 VTAIL.n255 9.3005
R505 VTAIL.n333 VTAIL.n332 9.3005
R506 VTAIL.n260 VTAIL.n259 9.3005
R507 VTAIL.n319 VTAIL.n318 9.3005
R508 VTAIL.n317 VTAIL.n316 9.3005
R509 VTAIL.n264 VTAIL.n263 9.3005
R510 VTAIL.n311 VTAIL.n310 9.3005
R511 VTAIL.n309 VTAIL.n308 9.3005
R512 VTAIL.n268 VTAIL.n267 9.3005
R513 VTAIL.n283 VTAIL.n282 9.3005
R514 VTAIL.n285 VTAIL.n284 9.3005
R515 VTAIL.n276 VTAIL.n275 9.3005
R516 VTAIL.n291 VTAIL.n290 9.3005
R517 VTAIL.n293 VTAIL.n292 9.3005
R518 VTAIL.n272 VTAIL.n271 9.3005
R519 VTAIL.n300 VTAIL.n299 9.3005
R520 VTAIL.n302 VTAIL.n301 9.3005
R521 VTAIL.n325 VTAIL.n324 9.3005
R522 VTAIL.n75 VTAIL.n74 9.3005
R523 VTAIL.n4 VTAIL.n3 9.3005
R524 VTAIL.n81 VTAIL.n80 9.3005
R525 VTAIL.n8 VTAIL.n7 9.3005
R526 VTAIL.n67 VTAIL.n66 9.3005
R527 VTAIL.n65 VTAIL.n64 9.3005
R528 VTAIL.n12 VTAIL.n11 9.3005
R529 VTAIL.n59 VTAIL.n58 9.3005
R530 VTAIL.n57 VTAIL.n56 9.3005
R531 VTAIL.n16 VTAIL.n15 9.3005
R532 VTAIL.n31 VTAIL.n30 9.3005
R533 VTAIL.n33 VTAIL.n32 9.3005
R534 VTAIL.n24 VTAIL.n23 9.3005
R535 VTAIL.n39 VTAIL.n38 9.3005
R536 VTAIL.n41 VTAIL.n40 9.3005
R537 VTAIL.n20 VTAIL.n19 9.3005
R538 VTAIL.n48 VTAIL.n47 9.3005
R539 VTAIL.n50 VTAIL.n49 9.3005
R540 VTAIL.n73 VTAIL.n72 9.3005
R541 VTAIL.n174 VTAIL.n173 9.3005
R542 VTAIL.n245 VTAIL.n244 9.3005
R543 VTAIL.n243 VTAIL.n242 9.3005
R544 VTAIL.n178 VTAIL.n177 9.3005
R545 VTAIL.n237 VTAIL.n236 9.3005
R546 VTAIL.n235 VTAIL.n234 9.3005
R547 VTAIL.n182 VTAIL.n181 9.3005
R548 VTAIL.n229 VTAIL.n228 9.3005
R549 VTAIL.n227 VTAIL.n226 9.3005
R550 VTAIL.n186 VTAIL.n185 9.3005
R551 VTAIL.n220 VTAIL.n219 9.3005
R552 VTAIL.n218 VTAIL.n217 9.3005
R553 VTAIL.n190 VTAIL.n189 9.3005
R554 VTAIL.n212 VTAIL.n211 9.3005
R555 VTAIL.n210 VTAIL.n209 9.3005
R556 VTAIL.n195 VTAIL.n194 9.3005
R557 VTAIL.n204 VTAIL.n203 9.3005
R558 VTAIL.n202 VTAIL.n201 9.3005
R559 VTAIL.n251 VTAIL.n250 9.3005
R560 VTAIL.n118 VTAIL.n117 9.3005
R561 VTAIL.n120 VTAIL.n119 9.3005
R562 VTAIL.n111 VTAIL.n110 9.3005
R563 VTAIL.n126 VTAIL.n125 9.3005
R564 VTAIL.n128 VTAIL.n127 9.3005
R565 VTAIL.n106 VTAIL.n105 9.3005
R566 VTAIL.n134 VTAIL.n133 9.3005
R567 VTAIL.n136 VTAIL.n135 9.3005
R568 VTAIL.n90 VTAIL.n89 9.3005
R569 VTAIL.n167 VTAIL.n166 9.3005
R570 VTAIL.n161 VTAIL.n160 9.3005
R571 VTAIL.n159 VTAIL.n158 9.3005
R572 VTAIL.n94 VTAIL.n93 9.3005
R573 VTAIL.n153 VTAIL.n152 9.3005
R574 VTAIL.n151 VTAIL.n150 9.3005
R575 VTAIL.n98 VTAIL.n97 9.3005
R576 VTAIL.n145 VTAIL.n144 9.3005
R577 VTAIL.n143 VTAIL.n142 9.3005
R578 VTAIL.n102 VTAIL.n101 9.3005
R579 VTAIL.n286 VTAIL.n276 8.92171
R580 VTAIL.n320 VTAIL.n319 8.92171
R581 VTAIL.n334 VTAIL.n254 8.92171
R582 VTAIL.n34 VTAIL.n24 8.92171
R583 VTAIL.n68 VTAIL.n67 8.92171
R584 VTAIL.n82 VTAIL.n2 8.92171
R585 VTAIL.n252 VTAIL.n172 8.92171
R586 VTAIL.n238 VTAIL.n237 8.92171
R587 VTAIL.n205 VTAIL.n195 8.92171
R588 VTAIL.n168 VTAIL.n88 8.92171
R589 VTAIL.n154 VTAIL.n153 8.92171
R590 VTAIL.n121 VTAIL.n111 8.92171
R591 VTAIL.n285 VTAIL.n278 8.14595
R592 VTAIL.n323 VTAIL.n260 8.14595
R593 VTAIL.n332 VTAIL.n331 8.14595
R594 VTAIL.n33 VTAIL.n26 8.14595
R595 VTAIL.n71 VTAIL.n8 8.14595
R596 VTAIL.n80 VTAIL.n79 8.14595
R597 VTAIL.n250 VTAIL.n249 8.14595
R598 VTAIL.n241 VTAIL.n178 8.14595
R599 VTAIL.n204 VTAIL.n197 8.14595
R600 VTAIL.n166 VTAIL.n165 8.14595
R601 VTAIL.n157 VTAIL.n94 8.14595
R602 VTAIL.n120 VTAIL.n113 8.14595
R603 VTAIL.n282 VTAIL.n281 7.3702
R604 VTAIL.n324 VTAIL.n258 7.3702
R605 VTAIL.n328 VTAIL.n256 7.3702
R606 VTAIL.n30 VTAIL.n29 7.3702
R607 VTAIL.n72 VTAIL.n6 7.3702
R608 VTAIL.n76 VTAIL.n4 7.3702
R609 VTAIL.n246 VTAIL.n174 7.3702
R610 VTAIL.n242 VTAIL.n176 7.3702
R611 VTAIL.n201 VTAIL.n200 7.3702
R612 VTAIL.n162 VTAIL.n90 7.3702
R613 VTAIL.n158 VTAIL.n92 7.3702
R614 VTAIL.n117 VTAIL.n116 7.3702
R615 VTAIL.n327 VTAIL.n258 6.59444
R616 VTAIL.n328 VTAIL.n327 6.59444
R617 VTAIL.n75 VTAIL.n6 6.59444
R618 VTAIL.n76 VTAIL.n75 6.59444
R619 VTAIL.n246 VTAIL.n245 6.59444
R620 VTAIL.n245 VTAIL.n176 6.59444
R621 VTAIL.n162 VTAIL.n161 6.59444
R622 VTAIL.n161 VTAIL.n92 6.59444
R623 VTAIL.n282 VTAIL.n278 5.81868
R624 VTAIL.n324 VTAIL.n323 5.81868
R625 VTAIL.n331 VTAIL.n256 5.81868
R626 VTAIL.n30 VTAIL.n26 5.81868
R627 VTAIL.n72 VTAIL.n71 5.81868
R628 VTAIL.n79 VTAIL.n4 5.81868
R629 VTAIL.n249 VTAIL.n174 5.81868
R630 VTAIL.n242 VTAIL.n241 5.81868
R631 VTAIL.n201 VTAIL.n197 5.81868
R632 VTAIL.n165 VTAIL.n90 5.81868
R633 VTAIL.n158 VTAIL.n157 5.81868
R634 VTAIL.n117 VTAIL.n113 5.81868
R635 VTAIL.n286 VTAIL.n285 5.04292
R636 VTAIL.n320 VTAIL.n260 5.04292
R637 VTAIL.n332 VTAIL.n254 5.04292
R638 VTAIL.n34 VTAIL.n33 5.04292
R639 VTAIL.n68 VTAIL.n8 5.04292
R640 VTAIL.n80 VTAIL.n2 5.04292
R641 VTAIL.n250 VTAIL.n172 5.04292
R642 VTAIL.n238 VTAIL.n178 5.04292
R643 VTAIL.n205 VTAIL.n204 5.04292
R644 VTAIL.n166 VTAIL.n88 5.04292
R645 VTAIL.n154 VTAIL.n94 5.04292
R646 VTAIL.n121 VTAIL.n120 5.04292
R647 VTAIL.n289 VTAIL.n276 4.26717
R648 VTAIL.n319 VTAIL.n262 4.26717
R649 VTAIL.n37 VTAIL.n24 4.26717
R650 VTAIL.n67 VTAIL.n10 4.26717
R651 VTAIL.n237 VTAIL.n180 4.26717
R652 VTAIL.n208 VTAIL.n195 4.26717
R653 VTAIL.n153 VTAIL.n96 4.26717
R654 VTAIL.n124 VTAIL.n111 4.26717
R655 VTAIL.n290 VTAIL.n274 3.49141
R656 VTAIL.n316 VTAIL.n315 3.49141
R657 VTAIL.n38 VTAIL.n22 3.49141
R658 VTAIL.n64 VTAIL.n63 3.49141
R659 VTAIL.n234 VTAIL.n233 3.49141
R660 VTAIL.n209 VTAIL.n193 3.49141
R661 VTAIL.n150 VTAIL.n149 3.49141
R662 VTAIL.n125 VTAIL.n109 3.49141
R663 VTAIL.n283 VTAIL.n279 2.84303
R664 VTAIL.n31 VTAIL.n27 2.84303
R665 VTAIL.n202 VTAIL.n198 2.84303
R666 VTAIL.n118 VTAIL.n114 2.84303
R667 VTAIL.n294 VTAIL.n293 2.71565
R668 VTAIL.n312 VTAIL.n264 2.71565
R669 VTAIL.n42 VTAIL.n41 2.71565
R670 VTAIL.n60 VTAIL.n12 2.71565
R671 VTAIL.n230 VTAIL.n182 2.71565
R672 VTAIL.n213 VTAIL.n212 2.71565
R673 VTAIL.n146 VTAIL.n98 2.71565
R674 VTAIL.n129 VTAIL.n128 2.71565
R675 VTAIL.n298 VTAIL.n272 1.93989
R676 VTAIL.n311 VTAIL.n266 1.93989
R677 VTAIL.n46 VTAIL.n20 1.93989
R678 VTAIL.n59 VTAIL.n14 1.93989
R679 VTAIL.n229 VTAIL.n184 1.93989
R680 VTAIL.n216 VTAIL.n190 1.93989
R681 VTAIL.n145 VTAIL.n100 1.93989
R682 VTAIL.n132 VTAIL.n106 1.93989
R683 VTAIL.n0 VTAIL.t2 1.33115
R684 VTAIL.n0 VTAIL.t1 1.33115
R685 VTAIL.n84 VTAIL.t6 1.33115
R686 VTAIL.n84 VTAIL.t11 1.33115
R687 VTAIL.n170 VTAIL.t10 1.33115
R688 VTAIL.n170 VTAIL.t9 1.33115
R689 VTAIL.n86 VTAIL.t3 1.33115
R690 VTAIL.n86 VTAIL.t4 1.33115
R691 VTAIL.n299 VTAIL.n270 1.16414
R692 VTAIL.n308 VTAIL.n307 1.16414
R693 VTAIL.n47 VTAIL.n18 1.16414
R694 VTAIL.n56 VTAIL.n55 1.16414
R695 VTAIL.n226 VTAIL.n225 1.16414
R696 VTAIL.n217 VTAIL.n188 1.16414
R697 VTAIL.n142 VTAIL.n141 1.16414
R698 VTAIL.n133 VTAIL.n104 1.16414
R699 VTAIL.n171 VTAIL.n169 0.862569
R700 VTAIL.n83 VTAIL.n1 0.862569
R701 VTAIL.n169 VTAIL.n87 0.784983
R702 VTAIL.n253 VTAIL.n171 0.784983
R703 VTAIL.n85 VTAIL.n83 0.784983
R704 VTAIL VTAIL.n335 0.530672
R705 VTAIL.n303 VTAIL.n302 0.388379
R706 VTAIL.n304 VTAIL.n268 0.388379
R707 VTAIL.n51 VTAIL.n50 0.388379
R708 VTAIL.n52 VTAIL.n16 0.388379
R709 VTAIL.n222 VTAIL.n186 0.388379
R710 VTAIL.n221 VTAIL.n220 0.388379
R711 VTAIL.n138 VTAIL.n102 0.388379
R712 VTAIL.n137 VTAIL.n136 0.388379
R713 VTAIL VTAIL.n1 0.25481
R714 VTAIL.n284 VTAIL.n283 0.155672
R715 VTAIL.n284 VTAIL.n275 0.155672
R716 VTAIL.n291 VTAIL.n275 0.155672
R717 VTAIL.n292 VTAIL.n291 0.155672
R718 VTAIL.n292 VTAIL.n271 0.155672
R719 VTAIL.n300 VTAIL.n271 0.155672
R720 VTAIL.n301 VTAIL.n300 0.155672
R721 VTAIL.n301 VTAIL.n267 0.155672
R722 VTAIL.n309 VTAIL.n267 0.155672
R723 VTAIL.n310 VTAIL.n309 0.155672
R724 VTAIL.n310 VTAIL.n263 0.155672
R725 VTAIL.n317 VTAIL.n263 0.155672
R726 VTAIL.n318 VTAIL.n317 0.155672
R727 VTAIL.n318 VTAIL.n259 0.155672
R728 VTAIL.n325 VTAIL.n259 0.155672
R729 VTAIL.n326 VTAIL.n325 0.155672
R730 VTAIL.n326 VTAIL.n255 0.155672
R731 VTAIL.n333 VTAIL.n255 0.155672
R732 VTAIL.n32 VTAIL.n31 0.155672
R733 VTAIL.n32 VTAIL.n23 0.155672
R734 VTAIL.n39 VTAIL.n23 0.155672
R735 VTAIL.n40 VTAIL.n39 0.155672
R736 VTAIL.n40 VTAIL.n19 0.155672
R737 VTAIL.n48 VTAIL.n19 0.155672
R738 VTAIL.n49 VTAIL.n48 0.155672
R739 VTAIL.n49 VTAIL.n15 0.155672
R740 VTAIL.n57 VTAIL.n15 0.155672
R741 VTAIL.n58 VTAIL.n57 0.155672
R742 VTAIL.n58 VTAIL.n11 0.155672
R743 VTAIL.n65 VTAIL.n11 0.155672
R744 VTAIL.n66 VTAIL.n65 0.155672
R745 VTAIL.n66 VTAIL.n7 0.155672
R746 VTAIL.n73 VTAIL.n7 0.155672
R747 VTAIL.n74 VTAIL.n73 0.155672
R748 VTAIL.n74 VTAIL.n3 0.155672
R749 VTAIL.n81 VTAIL.n3 0.155672
R750 VTAIL.n251 VTAIL.n173 0.155672
R751 VTAIL.n244 VTAIL.n173 0.155672
R752 VTAIL.n244 VTAIL.n243 0.155672
R753 VTAIL.n243 VTAIL.n177 0.155672
R754 VTAIL.n236 VTAIL.n177 0.155672
R755 VTAIL.n236 VTAIL.n235 0.155672
R756 VTAIL.n235 VTAIL.n181 0.155672
R757 VTAIL.n228 VTAIL.n181 0.155672
R758 VTAIL.n228 VTAIL.n227 0.155672
R759 VTAIL.n227 VTAIL.n185 0.155672
R760 VTAIL.n219 VTAIL.n185 0.155672
R761 VTAIL.n219 VTAIL.n218 0.155672
R762 VTAIL.n218 VTAIL.n189 0.155672
R763 VTAIL.n211 VTAIL.n189 0.155672
R764 VTAIL.n211 VTAIL.n210 0.155672
R765 VTAIL.n210 VTAIL.n194 0.155672
R766 VTAIL.n203 VTAIL.n194 0.155672
R767 VTAIL.n203 VTAIL.n202 0.155672
R768 VTAIL.n167 VTAIL.n89 0.155672
R769 VTAIL.n160 VTAIL.n89 0.155672
R770 VTAIL.n160 VTAIL.n159 0.155672
R771 VTAIL.n159 VTAIL.n93 0.155672
R772 VTAIL.n152 VTAIL.n93 0.155672
R773 VTAIL.n152 VTAIL.n151 0.155672
R774 VTAIL.n151 VTAIL.n97 0.155672
R775 VTAIL.n144 VTAIL.n97 0.155672
R776 VTAIL.n144 VTAIL.n143 0.155672
R777 VTAIL.n143 VTAIL.n101 0.155672
R778 VTAIL.n135 VTAIL.n101 0.155672
R779 VTAIL.n135 VTAIL.n134 0.155672
R780 VTAIL.n134 VTAIL.n105 0.155672
R781 VTAIL.n127 VTAIL.n105 0.155672
R782 VTAIL.n127 VTAIL.n126 0.155672
R783 VTAIL.n126 VTAIL.n110 0.155672
R784 VTAIL.n119 VTAIL.n110 0.155672
R785 VTAIL.n119 VTAIL.n118 0.155672
R786 B.n407 B.t10 823.035
R787 B.n405 B.t6 823.035
R788 B.n98 B.t17 823.035
R789 B.n95 B.t13 823.035
R790 B.n712 B.n711 585
R791 B.n313 B.n93 585
R792 B.n312 B.n311 585
R793 B.n310 B.n309 585
R794 B.n308 B.n307 585
R795 B.n306 B.n305 585
R796 B.n304 B.n303 585
R797 B.n302 B.n301 585
R798 B.n300 B.n299 585
R799 B.n298 B.n297 585
R800 B.n296 B.n295 585
R801 B.n294 B.n293 585
R802 B.n292 B.n291 585
R803 B.n290 B.n289 585
R804 B.n288 B.n287 585
R805 B.n286 B.n285 585
R806 B.n284 B.n283 585
R807 B.n282 B.n281 585
R808 B.n280 B.n279 585
R809 B.n278 B.n277 585
R810 B.n276 B.n275 585
R811 B.n274 B.n273 585
R812 B.n272 B.n271 585
R813 B.n270 B.n269 585
R814 B.n268 B.n267 585
R815 B.n266 B.n265 585
R816 B.n264 B.n263 585
R817 B.n262 B.n261 585
R818 B.n260 B.n259 585
R819 B.n258 B.n257 585
R820 B.n256 B.n255 585
R821 B.n254 B.n253 585
R822 B.n252 B.n251 585
R823 B.n250 B.n249 585
R824 B.n248 B.n247 585
R825 B.n246 B.n245 585
R826 B.n244 B.n243 585
R827 B.n242 B.n241 585
R828 B.n240 B.n239 585
R829 B.n238 B.n237 585
R830 B.n236 B.n235 585
R831 B.n234 B.n233 585
R832 B.n232 B.n231 585
R833 B.n230 B.n229 585
R834 B.n228 B.n227 585
R835 B.n226 B.n225 585
R836 B.n224 B.n223 585
R837 B.n222 B.n221 585
R838 B.n220 B.n219 585
R839 B.n218 B.n217 585
R840 B.n216 B.n215 585
R841 B.n214 B.n213 585
R842 B.n212 B.n211 585
R843 B.n210 B.n209 585
R844 B.n208 B.n207 585
R845 B.n206 B.n205 585
R846 B.n204 B.n203 585
R847 B.n202 B.n201 585
R848 B.n200 B.n199 585
R849 B.n198 B.n197 585
R850 B.n196 B.n195 585
R851 B.n194 B.n193 585
R852 B.n192 B.n191 585
R853 B.n190 B.n189 585
R854 B.n188 B.n187 585
R855 B.n186 B.n185 585
R856 B.n184 B.n183 585
R857 B.n182 B.n181 585
R858 B.n180 B.n179 585
R859 B.n178 B.n177 585
R860 B.n176 B.n175 585
R861 B.n174 B.n173 585
R862 B.n172 B.n171 585
R863 B.n170 B.n169 585
R864 B.n168 B.n167 585
R865 B.n166 B.n165 585
R866 B.n164 B.n163 585
R867 B.n162 B.n161 585
R868 B.n160 B.n159 585
R869 B.n158 B.n157 585
R870 B.n156 B.n155 585
R871 B.n154 B.n153 585
R872 B.n152 B.n151 585
R873 B.n150 B.n149 585
R874 B.n148 B.n147 585
R875 B.n146 B.n145 585
R876 B.n144 B.n143 585
R877 B.n142 B.n141 585
R878 B.n140 B.n139 585
R879 B.n138 B.n137 585
R880 B.n136 B.n135 585
R881 B.n134 B.n133 585
R882 B.n132 B.n131 585
R883 B.n130 B.n129 585
R884 B.n128 B.n127 585
R885 B.n126 B.n125 585
R886 B.n124 B.n123 585
R887 B.n122 B.n121 585
R888 B.n120 B.n119 585
R889 B.n118 B.n117 585
R890 B.n116 B.n115 585
R891 B.n114 B.n113 585
R892 B.n112 B.n111 585
R893 B.n110 B.n109 585
R894 B.n108 B.n107 585
R895 B.n106 B.n105 585
R896 B.n104 B.n103 585
R897 B.n102 B.n101 585
R898 B.n39 B.n38 585
R899 B.n717 B.n716 585
R900 B.n710 B.n94 585
R901 B.n94 B.n36 585
R902 B.n709 B.n35 585
R903 B.n721 B.n35 585
R904 B.n708 B.n34 585
R905 B.n722 B.n34 585
R906 B.n707 B.n33 585
R907 B.n723 B.n33 585
R908 B.n706 B.n705 585
R909 B.n705 B.n32 585
R910 B.n704 B.n28 585
R911 B.n729 B.n28 585
R912 B.n703 B.n27 585
R913 B.n730 B.n27 585
R914 B.n702 B.n26 585
R915 B.n731 B.n26 585
R916 B.n701 B.n700 585
R917 B.n700 B.n22 585
R918 B.n699 B.n21 585
R919 B.n737 B.n21 585
R920 B.n698 B.n20 585
R921 B.n738 B.n20 585
R922 B.n697 B.n19 585
R923 B.n739 B.n19 585
R924 B.n696 B.n695 585
R925 B.n695 B.n15 585
R926 B.n694 B.n14 585
R927 B.n745 B.n14 585
R928 B.n693 B.n13 585
R929 B.n746 B.n13 585
R930 B.n692 B.n12 585
R931 B.n747 B.n12 585
R932 B.n691 B.n690 585
R933 B.n690 B.n11 585
R934 B.n689 B.n7 585
R935 B.n753 B.n7 585
R936 B.n688 B.n6 585
R937 B.n754 B.n6 585
R938 B.n687 B.n5 585
R939 B.n755 B.n5 585
R940 B.n686 B.n685 585
R941 B.n685 B.n4 585
R942 B.n684 B.n314 585
R943 B.n684 B.n683 585
R944 B.n673 B.n315 585
R945 B.n676 B.n315 585
R946 B.n675 B.n674 585
R947 B.n677 B.n675 585
R948 B.n672 B.n320 585
R949 B.n320 B.n319 585
R950 B.n671 B.n670 585
R951 B.n670 B.n669 585
R952 B.n322 B.n321 585
R953 B.n323 B.n322 585
R954 B.n662 B.n661 585
R955 B.n663 B.n662 585
R956 B.n660 B.n327 585
R957 B.n331 B.n327 585
R958 B.n659 B.n658 585
R959 B.n658 B.n657 585
R960 B.n329 B.n328 585
R961 B.n330 B.n329 585
R962 B.n650 B.n649 585
R963 B.n651 B.n650 585
R964 B.n648 B.n336 585
R965 B.n336 B.n335 585
R966 B.n647 B.n646 585
R967 B.n646 B.n645 585
R968 B.n338 B.n337 585
R969 B.n638 B.n338 585
R970 B.n637 B.n636 585
R971 B.n639 B.n637 585
R972 B.n635 B.n343 585
R973 B.n343 B.n342 585
R974 B.n634 B.n633 585
R975 B.n633 B.n632 585
R976 B.n345 B.n344 585
R977 B.n346 B.n345 585
R978 B.n628 B.n627 585
R979 B.n349 B.n348 585
R980 B.n624 B.n623 585
R981 B.n625 B.n624 585
R982 B.n622 B.n404 585
R983 B.n621 B.n620 585
R984 B.n619 B.n618 585
R985 B.n617 B.n616 585
R986 B.n615 B.n614 585
R987 B.n613 B.n612 585
R988 B.n611 B.n610 585
R989 B.n609 B.n608 585
R990 B.n607 B.n606 585
R991 B.n605 B.n604 585
R992 B.n603 B.n602 585
R993 B.n601 B.n600 585
R994 B.n599 B.n598 585
R995 B.n597 B.n596 585
R996 B.n595 B.n594 585
R997 B.n593 B.n592 585
R998 B.n591 B.n590 585
R999 B.n589 B.n588 585
R1000 B.n587 B.n586 585
R1001 B.n585 B.n584 585
R1002 B.n583 B.n582 585
R1003 B.n581 B.n580 585
R1004 B.n579 B.n578 585
R1005 B.n577 B.n576 585
R1006 B.n575 B.n574 585
R1007 B.n573 B.n572 585
R1008 B.n571 B.n570 585
R1009 B.n569 B.n568 585
R1010 B.n567 B.n566 585
R1011 B.n565 B.n564 585
R1012 B.n563 B.n562 585
R1013 B.n561 B.n560 585
R1014 B.n559 B.n558 585
R1015 B.n557 B.n556 585
R1016 B.n555 B.n554 585
R1017 B.n553 B.n552 585
R1018 B.n551 B.n550 585
R1019 B.n549 B.n548 585
R1020 B.n547 B.n546 585
R1021 B.n545 B.n544 585
R1022 B.n543 B.n542 585
R1023 B.n541 B.n540 585
R1024 B.n539 B.n538 585
R1025 B.n537 B.n536 585
R1026 B.n535 B.n534 585
R1027 B.n533 B.n532 585
R1028 B.n531 B.n530 585
R1029 B.n528 B.n527 585
R1030 B.n526 B.n525 585
R1031 B.n524 B.n523 585
R1032 B.n522 B.n521 585
R1033 B.n520 B.n519 585
R1034 B.n518 B.n517 585
R1035 B.n516 B.n515 585
R1036 B.n514 B.n513 585
R1037 B.n512 B.n511 585
R1038 B.n510 B.n509 585
R1039 B.n507 B.n506 585
R1040 B.n505 B.n504 585
R1041 B.n503 B.n502 585
R1042 B.n501 B.n500 585
R1043 B.n499 B.n498 585
R1044 B.n497 B.n496 585
R1045 B.n495 B.n494 585
R1046 B.n493 B.n492 585
R1047 B.n491 B.n490 585
R1048 B.n489 B.n488 585
R1049 B.n487 B.n486 585
R1050 B.n485 B.n484 585
R1051 B.n483 B.n482 585
R1052 B.n481 B.n480 585
R1053 B.n479 B.n478 585
R1054 B.n477 B.n476 585
R1055 B.n475 B.n474 585
R1056 B.n473 B.n472 585
R1057 B.n471 B.n470 585
R1058 B.n469 B.n468 585
R1059 B.n467 B.n466 585
R1060 B.n465 B.n464 585
R1061 B.n463 B.n462 585
R1062 B.n461 B.n460 585
R1063 B.n459 B.n458 585
R1064 B.n457 B.n456 585
R1065 B.n455 B.n454 585
R1066 B.n453 B.n452 585
R1067 B.n451 B.n450 585
R1068 B.n449 B.n448 585
R1069 B.n447 B.n446 585
R1070 B.n445 B.n444 585
R1071 B.n443 B.n442 585
R1072 B.n441 B.n440 585
R1073 B.n439 B.n438 585
R1074 B.n437 B.n436 585
R1075 B.n435 B.n434 585
R1076 B.n433 B.n432 585
R1077 B.n431 B.n430 585
R1078 B.n429 B.n428 585
R1079 B.n427 B.n426 585
R1080 B.n425 B.n424 585
R1081 B.n423 B.n422 585
R1082 B.n421 B.n420 585
R1083 B.n419 B.n418 585
R1084 B.n417 B.n416 585
R1085 B.n415 B.n414 585
R1086 B.n413 B.n412 585
R1087 B.n411 B.n410 585
R1088 B.n409 B.n403 585
R1089 B.n625 B.n403 585
R1090 B.n629 B.n347 585
R1091 B.n347 B.n346 585
R1092 B.n631 B.n630 585
R1093 B.n632 B.n631 585
R1094 B.n341 B.n340 585
R1095 B.n342 B.n341 585
R1096 B.n641 B.n640 585
R1097 B.n640 B.n639 585
R1098 B.n642 B.n339 585
R1099 B.n638 B.n339 585
R1100 B.n644 B.n643 585
R1101 B.n645 B.n644 585
R1102 B.n334 B.n333 585
R1103 B.n335 B.n334 585
R1104 B.n653 B.n652 585
R1105 B.n652 B.n651 585
R1106 B.n654 B.n332 585
R1107 B.n332 B.n330 585
R1108 B.n656 B.n655 585
R1109 B.n657 B.n656 585
R1110 B.n326 B.n325 585
R1111 B.n331 B.n326 585
R1112 B.n665 B.n664 585
R1113 B.n664 B.n663 585
R1114 B.n666 B.n324 585
R1115 B.n324 B.n323 585
R1116 B.n668 B.n667 585
R1117 B.n669 B.n668 585
R1118 B.n318 B.n317 585
R1119 B.n319 B.n318 585
R1120 B.n679 B.n678 585
R1121 B.n678 B.n677 585
R1122 B.n680 B.n316 585
R1123 B.n676 B.n316 585
R1124 B.n682 B.n681 585
R1125 B.n683 B.n682 585
R1126 B.n2 B.n0 585
R1127 B.n4 B.n2 585
R1128 B.n3 B.n1 585
R1129 B.n754 B.n3 585
R1130 B.n752 B.n751 585
R1131 B.n753 B.n752 585
R1132 B.n750 B.n8 585
R1133 B.n11 B.n8 585
R1134 B.n749 B.n748 585
R1135 B.n748 B.n747 585
R1136 B.n10 B.n9 585
R1137 B.n746 B.n10 585
R1138 B.n744 B.n743 585
R1139 B.n745 B.n744 585
R1140 B.n742 B.n16 585
R1141 B.n16 B.n15 585
R1142 B.n741 B.n740 585
R1143 B.n740 B.n739 585
R1144 B.n18 B.n17 585
R1145 B.n738 B.n18 585
R1146 B.n736 B.n735 585
R1147 B.n737 B.n736 585
R1148 B.n734 B.n23 585
R1149 B.n23 B.n22 585
R1150 B.n733 B.n732 585
R1151 B.n732 B.n731 585
R1152 B.n25 B.n24 585
R1153 B.n730 B.n25 585
R1154 B.n728 B.n727 585
R1155 B.n729 B.n728 585
R1156 B.n726 B.n29 585
R1157 B.n32 B.n29 585
R1158 B.n725 B.n724 585
R1159 B.n724 B.n723 585
R1160 B.n31 B.n30 585
R1161 B.n722 B.n31 585
R1162 B.n720 B.n719 585
R1163 B.n721 B.n720 585
R1164 B.n718 B.n37 585
R1165 B.n37 B.n36 585
R1166 B.n757 B.n756 585
R1167 B.n756 B.n755 585
R1168 B.n627 B.n347 449.257
R1169 B.n716 B.n37 449.257
R1170 B.n403 B.n345 449.257
R1171 B.n712 B.n94 449.257
R1172 B.n407 B.t12 349.61
R1173 B.n95 B.t15 349.61
R1174 B.n405 B.t9 349.61
R1175 B.n98 B.t18 349.61
R1176 B.n408 B.t11 331.961
R1177 B.n96 B.t16 331.961
R1178 B.n406 B.t8 331.961
R1179 B.n99 B.t19 331.961
R1180 B.n714 B.n713 256.663
R1181 B.n714 B.n92 256.663
R1182 B.n714 B.n91 256.663
R1183 B.n714 B.n90 256.663
R1184 B.n714 B.n89 256.663
R1185 B.n714 B.n88 256.663
R1186 B.n714 B.n87 256.663
R1187 B.n714 B.n86 256.663
R1188 B.n714 B.n85 256.663
R1189 B.n714 B.n84 256.663
R1190 B.n714 B.n83 256.663
R1191 B.n714 B.n82 256.663
R1192 B.n714 B.n81 256.663
R1193 B.n714 B.n80 256.663
R1194 B.n714 B.n79 256.663
R1195 B.n714 B.n78 256.663
R1196 B.n714 B.n77 256.663
R1197 B.n714 B.n76 256.663
R1198 B.n714 B.n75 256.663
R1199 B.n714 B.n74 256.663
R1200 B.n714 B.n73 256.663
R1201 B.n714 B.n72 256.663
R1202 B.n714 B.n71 256.663
R1203 B.n714 B.n70 256.663
R1204 B.n714 B.n69 256.663
R1205 B.n714 B.n68 256.663
R1206 B.n714 B.n67 256.663
R1207 B.n714 B.n66 256.663
R1208 B.n714 B.n65 256.663
R1209 B.n714 B.n64 256.663
R1210 B.n714 B.n63 256.663
R1211 B.n714 B.n62 256.663
R1212 B.n714 B.n61 256.663
R1213 B.n714 B.n60 256.663
R1214 B.n714 B.n59 256.663
R1215 B.n714 B.n58 256.663
R1216 B.n714 B.n57 256.663
R1217 B.n714 B.n56 256.663
R1218 B.n714 B.n55 256.663
R1219 B.n714 B.n54 256.663
R1220 B.n714 B.n53 256.663
R1221 B.n714 B.n52 256.663
R1222 B.n714 B.n51 256.663
R1223 B.n714 B.n50 256.663
R1224 B.n714 B.n49 256.663
R1225 B.n714 B.n48 256.663
R1226 B.n714 B.n47 256.663
R1227 B.n714 B.n46 256.663
R1228 B.n714 B.n45 256.663
R1229 B.n714 B.n44 256.663
R1230 B.n714 B.n43 256.663
R1231 B.n714 B.n42 256.663
R1232 B.n714 B.n41 256.663
R1233 B.n714 B.n40 256.663
R1234 B.n715 B.n714 256.663
R1235 B.n626 B.n625 256.663
R1236 B.n625 B.n350 256.663
R1237 B.n625 B.n351 256.663
R1238 B.n625 B.n352 256.663
R1239 B.n625 B.n353 256.663
R1240 B.n625 B.n354 256.663
R1241 B.n625 B.n355 256.663
R1242 B.n625 B.n356 256.663
R1243 B.n625 B.n357 256.663
R1244 B.n625 B.n358 256.663
R1245 B.n625 B.n359 256.663
R1246 B.n625 B.n360 256.663
R1247 B.n625 B.n361 256.663
R1248 B.n625 B.n362 256.663
R1249 B.n625 B.n363 256.663
R1250 B.n625 B.n364 256.663
R1251 B.n625 B.n365 256.663
R1252 B.n625 B.n366 256.663
R1253 B.n625 B.n367 256.663
R1254 B.n625 B.n368 256.663
R1255 B.n625 B.n369 256.663
R1256 B.n625 B.n370 256.663
R1257 B.n625 B.n371 256.663
R1258 B.n625 B.n372 256.663
R1259 B.n625 B.n373 256.663
R1260 B.n625 B.n374 256.663
R1261 B.n625 B.n375 256.663
R1262 B.n625 B.n376 256.663
R1263 B.n625 B.n377 256.663
R1264 B.n625 B.n378 256.663
R1265 B.n625 B.n379 256.663
R1266 B.n625 B.n380 256.663
R1267 B.n625 B.n381 256.663
R1268 B.n625 B.n382 256.663
R1269 B.n625 B.n383 256.663
R1270 B.n625 B.n384 256.663
R1271 B.n625 B.n385 256.663
R1272 B.n625 B.n386 256.663
R1273 B.n625 B.n387 256.663
R1274 B.n625 B.n388 256.663
R1275 B.n625 B.n389 256.663
R1276 B.n625 B.n390 256.663
R1277 B.n625 B.n391 256.663
R1278 B.n625 B.n392 256.663
R1279 B.n625 B.n393 256.663
R1280 B.n625 B.n394 256.663
R1281 B.n625 B.n395 256.663
R1282 B.n625 B.n396 256.663
R1283 B.n625 B.n397 256.663
R1284 B.n625 B.n398 256.663
R1285 B.n625 B.n399 256.663
R1286 B.n625 B.n400 256.663
R1287 B.n625 B.n401 256.663
R1288 B.n625 B.n402 256.663
R1289 B.n631 B.n347 163.367
R1290 B.n631 B.n341 163.367
R1291 B.n640 B.n341 163.367
R1292 B.n640 B.n339 163.367
R1293 B.n644 B.n339 163.367
R1294 B.n644 B.n334 163.367
R1295 B.n652 B.n334 163.367
R1296 B.n652 B.n332 163.367
R1297 B.n656 B.n332 163.367
R1298 B.n656 B.n326 163.367
R1299 B.n664 B.n326 163.367
R1300 B.n664 B.n324 163.367
R1301 B.n668 B.n324 163.367
R1302 B.n668 B.n318 163.367
R1303 B.n678 B.n318 163.367
R1304 B.n678 B.n316 163.367
R1305 B.n682 B.n316 163.367
R1306 B.n682 B.n2 163.367
R1307 B.n756 B.n2 163.367
R1308 B.n756 B.n3 163.367
R1309 B.n752 B.n3 163.367
R1310 B.n752 B.n8 163.367
R1311 B.n748 B.n8 163.367
R1312 B.n748 B.n10 163.367
R1313 B.n744 B.n10 163.367
R1314 B.n744 B.n16 163.367
R1315 B.n740 B.n16 163.367
R1316 B.n740 B.n18 163.367
R1317 B.n736 B.n18 163.367
R1318 B.n736 B.n23 163.367
R1319 B.n732 B.n23 163.367
R1320 B.n732 B.n25 163.367
R1321 B.n728 B.n25 163.367
R1322 B.n728 B.n29 163.367
R1323 B.n724 B.n29 163.367
R1324 B.n724 B.n31 163.367
R1325 B.n720 B.n31 163.367
R1326 B.n720 B.n37 163.367
R1327 B.n624 B.n349 163.367
R1328 B.n624 B.n404 163.367
R1329 B.n620 B.n619 163.367
R1330 B.n616 B.n615 163.367
R1331 B.n612 B.n611 163.367
R1332 B.n608 B.n607 163.367
R1333 B.n604 B.n603 163.367
R1334 B.n600 B.n599 163.367
R1335 B.n596 B.n595 163.367
R1336 B.n592 B.n591 163.367
R1337 B.n588 B.n587 163.367
R1338 B.n584 B.n583 163.367
R1339 B.n580 B.n579 163.367
R1340 B.n576 B.n575 163.367
R1341 B.n572 B.n571 163.367
R1342 B.n568 B.n567 163.367
R1343 B.n564 B.n563 163.367
R1344 B.n560 B.n559 163.367
R1345 B.n556 B.n555 163.367
R1346 B.n552 B.n551 163.367
R1347 B.n548 B.n547 163.367
R1348 B.n544 B.n543 163.367
R1349 B.n540 B.n539 163.367
R1350 B.n536 B.n535 163.367
R1351 B.n532 B.n531 163.367
R1352 B.n527 B.n526 163.367
R1353 B.n523 B.n522 163.367
R1354 B.n519 B.n518 163.367
R1355 B.n515 B.n514 163.367
R1356 B.n511 B.n510 163.367
R1357 B.n506 B.n505 163.367
R1358 B.n502 B.n501 163.367
R1359 B.n498 B.n497 163.367
R1360 B.n494 B.n493 163.367
R1361 B.n490 B.n489 163.367
R1362 B.n486 B.n485 163.367
R1363 B.n482 B.n481 163.367
R1364 B.n478 B.n477 163.367
R1365 B.n474 B.n473 163.367
R1366 B.n470 B.n469 163.367
R1367 B.n466 B.n465 163.367
R1368 B.n462 B.n461 163.367
R1369 B.n458 B.n457 163.367
R1370 B.n454 B.n453 163.367
R1371 B.n450 B.n449 163.367
R1372 B.n446 B.n445 163.367
R1373 B.n442 B.n441 163.367
R1374 B.n438 B.n437 163.367
R1375 B.n434 B.n433 163.367
R1376 B.n430 B.n429 163.367
R1377 B.n426 B.n425 163.367
R1378 B.n422 B.n421 163.367
R1379 B.n418 B.n417 163.367
R1380 B.n414 B.n413 163.367
R1381 B.n410 B.n403 163.367
R1382 B.n633 B.n345 163.367
R1383 B.n633 B.n343 163.367
R1384 B.n637 B.n343 163.367
R1385 B.n637 B.n338 163.367
R1386 B.n646 B.n338 163.367
R1387 B.n646 B.n336 163.367
R1388 B.n650 B.n336 163.367
R1389 B.n650 B.n329 163.367
R1390 B.n658 B.n329 163.367
R1391 B.n658 B.n327 163.367
R1392 B.n662 B.n327 163.367
R1393 B.n662 B.n322 163.367
R1394 B.n670 B.n322 163.367
R1395 B.n670 B.n320 163.367
R1396 B.n675 B.n320 163.367
R1397 B.n675 B.n315 163.367
R1398 B.n684 B.n315 163.367
R1399 B.n685 B.n684 163.367
R1400 B.n685 B.n5 163.367
R1401 B.n6 B.n5 163.367
R1402 B.n7 B.n6 163.367
R1403 B.n690 B.n7 163.367
R1404 B.n690 B.n12 163.367
R1405 B.n13 B.n12 163.367
R1406 B.n14 B.n13 163.367
R1407 B.n695 B.n14 163.367
R1408 B.n695 B.n19 163.367
R1409 B.n20 B.n19 163.367
R1410 B.n21 B.n20 163.367
R1411 B.n700 B.n21 163.367
R1412 B.n700 B.n26 163.367
R1413 B.n27 B.n26 163.367
R1414 B.n28 B.n27 163.367
R1415 B.n705 B.n28 163.367
R1416 B.n705 B.n33 163.367
R1417 B.n34 B.n33 163.367
R1418 B.n35 B.n34 163.367
R1419 B.n94 B.n35 163.367
R1420 B.n101 B.n39 163.367
R1421 B.n105 B.n104 163.367
R1422 B.n109 B.n108 163.367
R1423 B.n113 B.n112 163.367
R1424 B.n117 B.n116 163.367
R1425 B.n121 B.n120 163.367
R1426 B.n125 B.n124 163.367
R1427 B.n129 B.n128 163.367
R1428 B.n133 B.n132 163.367
R1429 B.n137 B.n136 163.367
R1430 B.n141 B.n140 163.367
R1431 B.n145 B.n144 163.367
R1432 B.n149 B.n148 163.367
R1433 B.n153 B.n152 163.367
R1434 B.n157 B.n156 163.367
R1435 B.n161 B.n160 163.367
R1436 B.n165 B.n164 163.367
R1437 B.n169 B.n168 163.367
R1438 B.n173 B.n172 163.367
R1439 B.n177 B.n176 163.367
R1440 B.n181 B.n180 163.367
R1441 B.n185 B.n184 163.367
R1442 B.n189 B.n188 163.367
R1443 B.n193 B.n192 163.367
R1444 B.n197 B.n196 163.367
R1445 B.n201 B.n200 163.367
R1446 B.n205 B.n204 163.367
R1447 B.n209 B.n208 163.367
R1448 B.n213 B.n212 163.367
R1449 B.n217 B.n216 163.367
R1450 B.n221 B.n220 163.367
R1451 B.n225 B.n224 163.367
R1452 B.n229 B.n228 163.367
R1453 B.n233 B.n232 163.367
R1454 B.n237 B.n236 163.367
R1455 B.n241 B.n240 163.367
R1456 B.n245 B.n244 163.367
R1457 B.n249 B.n248 163.367
R1458 B.n253 B.n252 163.367
R1459 B.n257 B.n256 163.367
R1460 B.n261 B.n260 163.367
R1461 B.n265 B.n264 163.367
R1462 B.n269 B.n268 163.367
R1463 B.n273 B.n272 163.367
R1464 B.n277 B.n276 163.367
R1465 B.n281 B.n280 163.367
R1466 B.n285 B.n284 163.367
R1467 B.n289 B.n288 163.367
R1468 B.n293 B.n292 163.367
R1469 B.n297 B.n296 163.367
R1470 B.n301 B.n300 163.367
R1471 B.n305 B.n304 163.367
R1472 B.n309 B.n308 163.367
R1473 B.n311 B.n93 163.367
R1474 B.n627 B.n626 71.676
R1475 B.n404 B.n350 71.676
R1476 B.n619 B.n351 71.676
R1477 B.n615 B.n352 71.676
R1478 B.n611 B.n353 71.676
R1479 B.n607 B.n354 71.676
R1480 B.n603 B.n355 71.676
R1481 B.n599 B.n356 71.676
R1482 B.n595 B.n357 71.676
R1483 B.n591 B.n358 71.676
R1484 B.n587 B.n359 71.676
R1485 B.n583 B.n360 71.676
R1486 B.n579 B.n361 71.676
R1487 B.n575 B.n362 71.676
R1488 B.n571 B.n363 71.676
R1489 B.n567 B.n364 71.676
R1490 B.n563 B.n365 71.676
R1491 B.n559 B.n366 71.676
R1492 B.n555 B.n367 71.676
R1493 B.n551 B.n368 71.676
R1494 B.n547 B.n369 71.676
R1495 B.n543 B.n370 71.676
R1496 B.n539 B.n371 71.676
R1497 B.n535 B.n372 71.676
R1498 B.n531 B.n373 71.676
R1499 B.n526 B.n374 71.676
R1500 B.n522 B.n375 71.676
R1501 B.n518 B.n376 71.676
R1502 B.n514 B.n377 71.676
R1503 B.n510 B.n378 71.676
R1504 B.n505 B.n379 71.676
R1505 B.n501 B.n380 71.676
R1506 B.n497 B.n381 71.676
R1507 B.n493 B.n382 71.676
R1508 B.n489 B.n383 71.676
R1509 B.n485 B.n384 71.676
R1510 B.n481 B.n385 71.676
R1511 B.n477 B.n386 71.676
R1512 B.n473 B.n387 71.676
R1513 B.n469 B.n388 71.676
R1514 B.n465 B.n389 71.676
R1515 B.n461 B.n390 71.676
R1516 B.n457 B.n391 71.676
R1517 B.n453 B.n392 71.676
R1518 B.n449 B.n393 71.676
R1519 B.n445 B.n394 71.676
R1520 B.n441 B.n395 71.676
R1521 B.n437 B.n396 71.676
R1522 B.n433 B.n397 71.676
R1523 B.n429 B.n398 71.676
R1524 B.n425 B.n399 71.676
R1525 B.n421 B.n400 71.676
R1526 B.n417 B.n401 71.676
R1527 B.n413 B.n402 71.676
R1528 B.n716 B.n715 71.676
R1529 B.n101 B.n40 71.676
R1530 B.n105 B.n41 71.676
R1531 B.n109 B.n42 71.676
R1532 B.n113 B.n43 71.676
R1533 B.n117 B.n44 71.676
R1534 B.n121 B.n45 71.676
R1535 B.n125 B.n46 71.676
R1536 B.n129 B.n47 71.676
R1537 B.n133 B.n48 71.676
R1538 B.n137 B.n49 71.676
R1539 B.n141 B.n50 71.676
R1540 B.n145 B.n51 71.676
R1541 B.n149 B.n52 71.676
R1542 B.n153 B.n53 71.676
R1543 B.n157 B.n54 71.676
R1544 B.n161 B.n55 71.676
R1545 B.n165 B.n56 71.676
R1546 B.n169 B.n57 71.676
R1547 B.n173 B.n58 71.676
R1548 B.n177 B.n59 71.676
R1549 B.n181 B.n60 71.676
R1550 B.n185 B.n61 71.676
R1551 B.n189 B.n62 71.676
R1552 B.n193 B.n63 71.676
R1553 B.n197 B.n64 71.676
R1554 B.n201 B.n65 71.676
R1555 B.n205 B.n66 71.676
R1556 B.n209 B.n67 71.676
R1557 B.n213 B.n68 71.676
R1558 B.n217 B.n69 71.676
R1559 B.n221 B.n70 71.676
R1560 B.n225 B.n71 71.676
R1561 B.n229 B.n72 71.676
R1562 B.n233 B.n73 71.676
R1563 B.n237 B.n74 71.676
R1564 B.n241 B.n75 71.676
R1565 B.n245 B.n76 71.676
R1566 B.n249 B.n77 71.676
R1567 B.n253 B.n78 71.676
R1568 B.n257 B.n79 71.676
R1569 B.n261 B.n80 71.676
R1570 B.n265 B.n81 71.676
R1571 B.n269 B.n82 71.676
R1572 B.n273 B.n83 71.676
R1573 B.n277 B.n84 71.676
R1574 B.n281 B.n85 71.676
R1575 B.n285 B.n86 71.676
R1576 B.n289 B.n87 71.676
R1577 B.n293 B.n88 71.676
R1578 B.n297 B.n89 71.676
R1579 B.n301 B.n90 71.676
R1580 B.n305 B.n91 71.676
R1581 B.n309 B.n92 71.676
R1582 B.n713 B.n93 71.676
R1583 B.n713 B.n712 71.676
R1584 B.n311 B.n92 71.676
R1585 B.n308 B.n91 71.676
R1586 B.n304 B.n90 71.676
R1587 B.n300 B.n89 71.676
R1588 B.n296 B.n88 71.676
R1589 B.n292 B.n87 71.676
R1590 B.n288 B.n86 71.676
R1591 B.n284 B.n85 71.676
R1592 B.n280 B.n84 71.676
R1593 B.n276 B.n83 71.676
R1594 B.n272 B.n82 71.676
R1595 B.n268 B.n81 71.676
R1596 B.n264 B.n80 71.676
R1597 B.n260 B.n79 71.676
R1598 B.n256 B.n78 71.676
R1599 B.n252 B.n77 71.676
R1600 B.n248 B.n76 71.676
R1601 B.n244 B.n75 71.676
R1602 B.n240 B.n74 71.676
R1603 B.n236 B.n73 71.676
R1604 B.n232 B.n72 71.676
R1605 B.n228 B.n71 71.676
R1606 B.n224 B.n70 71.676
R1607 B.n220 B.n69 71.676
R1608 B.n216 B.n68 71.676
R1609 B.n212 B.n67 71.676
R1610 B.n208 B.n66 71.676
R1611 B.n204 B.n65 71.676
R1612 B.n200 B.n64 71.676
R1613 B.n196 B.n63 71.676
R1614 B.n192 B.n62 71.676
R1615 B.n188 B.n61 71.676
R1616 B.n184 B.n60 71.676
R1617 B.n180 B.n59 71.676
R1618 B.n176 B.n58 71.676
R1619 B.n172 B.n57 71.676
R1620 B.n168 B.n56 71.676
R1621 B.n164 B.n55 71.676
R1622 B.n160 B.n54 71.676
R1623 B.n156 B.n53 71.676
R1624 B.n152 B.n52 71.676
R1625 B.n148 B.n51 71.676
R1626 B.n144 B.n50 71.676
R1627 B.n140 B.n49 71.676
R1628 B.n136 B.n48 71.676
R1629 B.n132 B.n47 71.676
R1630 B.n128 B.n46 71.676
R1631 B.n124 B.n45 71.676
R1632 B.n120 B.n44 71.676
R1633 B.n116 B.n43 71.676
R1634 B.n112 B.n42 71.676
R1635 B.n108 B.n41 71.676
R1636 B.n104 B.n40 71.676
R1637 B.n715 B.n39 71.676
R1638 B.n626 B.n349 71.676
R1639 B.n620 B.n350 71.676
R1640 B.n616 B.n351 71.676
R1641 B.n612 B.n352 71.676
R1642 B.n608 B.n353 71.676
R1643 B.n604 B.n354 71.676
R1644 B.n600 B.n355 71.676
R1645 B.n596 B.n356 71.676
R1646 B.n592 B.n357 71.676
R1647 B.n588 B.n358 71.676
R1648 B.n584 B.n359 71.676
R1649 B.n580 B.n360 71.676
R1650 B.n576 B.n361 71.676
R1651 B.n572 B.n362 71.676
R1652 B.n568 B.n363 71.676
R1653 B.n564 B.n364 71.676
R1654 B.n560 B.n365 71.676
R1655 B.n556 B.n366 71.676
R1656 B.n552 B.n367 71.676
R1657 B.n548 B.n368 71.676
R1658 B.n544 B.n369 71.676
R1659 B.n540 B.n370 71.676
R1660 B.n536 B.n371 71.676
R1661 B.n532 B.n372 71.676
R1662 B.n527 B.n373 71.676
R1663 B.n523 B.n374 71.676
R1664 B.n519 B.n375 71.676
R1665 B.n515 B.n376 71.676
R1666 B.n511 B.n377 71.676
R1667 B.n506 B.n378 71.676
R1668 B.n502 B.n379 71.676
R1669 B.n498 B.n380 71.676
R1670 B.n494 B.n381 71.676
R1671 B.n490 B.n382 71.676
R1672 B.n486 B.n383 71.676
R1673 B.n482 B.n384 71.676
R1674 B.n478 B.n385 71.676
R1675 B.n474 B.n386 71.676
R1676 B.n470 B.n387 71.676
R1677 B.n466 B.n388 71.676
R1678 B.n462 B.n389 71.676
R1679 B.n458 B.n390 71.676
R1680 B.n454 B.n391 71.676
R1681 B.n450 B.n392 71.676
R1682 B.n446 B.n393 71.676
R1683 B.n442 B.n394 71.676
R1684 B.n438 B.n395 71.676
R1685 B.n434 B.n396 71.676
R1686 B.n430 B.n397 71.676
R1687 B.n426 B.n398 71.676
R1688 B.n422 B.n399 71.676
R1689 B.n418 B.n400 71.676
R1690 B.n414 B.n401 71.676
R1691 B.n410 B.n402 71.676
R1692 B.n625 B.n346 60.581
R1693 B.n714 B.n36 60.581
R1694 B.n508 B.n408 59.5399
R1695 B.n529 B.n406 59.5399
R1696 B.n100 B.n99 59.5399
R1697 B.n97 B.n96 59.5399
R1698 B.n632 B.n346 37.1129
R1699 B.n632 B.n342 37.1129
R1700 B.n639 B.n342 37.1129
R1701 B.n639 B.n638 37.1129
R1702 B.n645 B.n335 37.1129
R1703 B.n651 B.n335 37.1129
R1704 B.n651 B.n330 37.1129
R1705 B.n657 B.n330 37.1129
R1706 B.n657 B.n331 37.1129
R1707 B.n663 B.n323 37.1129
R1708 B.n669 B.n323 37.1129
R1709 B.n677 B.n319 37.1129
R1710 B.n677 B.n676 37.1129
R1711 B.n683 B.n4 37.1129
R1712 B.n755 B.n4 37.1129
R1713 B.n755 B.n754 37.1129
R1714 B.n754 B.n753 37.1129
R1715 B.n747 B.n11 37.1129
R1716 B.n747 B.n746 37.1129
R1717 B.n745 B.n15 37.1129
R1718 B.n739 B.n15 37.1129
R1719 B.n738 B.n737 37.1129
R1720 B.n737 B.n22 37.1129
R1721 B.n731 B.n22 37.1129
R1722 B.n731 B.n730 37.1129
R1723 B.n730 B.n729 37.1129
R1724 B.n723 B.n32 37.1129
R1725 B.n723 B.n722 37.1129
R1726 B.n722 B.n721 37.1129
R1727 B.n721 B.n36 37.1129
R1728 B.n683 B.t0 34.9298
R1729 B.n753 B.t2 34.9298
R1730 B.n638 B.t7 30.5636
R1731 B.n32 B.t14 30.5636
R1732 B.n718 B.n717 29.1907
R1733 B.n409 B.n344 29.1907
R1734 B.n629 B.n628 29.1907
R1735 B.n711 B.n710 29.1907
R1736 B.n331 B.t3 26.1975
R1737 B.t5 B.n738 26.1975
R1738 B.t4 B.n319 22.9229
R1739 B.n746 B.t1 22.9229
R1740 B B.n757 18.0485
R1741 B.n408 B.n407 17.649
R1742 B.n406 B.n405 17.649
R1743 B.n99 B.n98 17.649
R1744 B.n96 B.n95 17.649
R1745 B.n669 B.t4 14.1905
R1746 B.t1 B.n745 14.1905
R1747 B.n663 B.t3 10.9159
R1748 B.n739 B.t5 10.9159
R1749 B.n717 B.n38 10.6151
R1750 B.n102 B.n38 10.6151
R1751 B.n103 B.n102 10.6151
R1752 B.n106 B.n103 10.6151
R1753 B.n107 B.n106 10.6151
R1754 B.n110 B.n107 10.6151
R1755 B.n111 B.n110 10.6151
R1756 B.n114 B.n111 10.6151
R1757 B.n115 B.n114 10.6151
R1758 B.n118 B.n115 10.6151
R1759 B.n119 B.n118 10.6151
R1760 B.n122 B.n119 10.6151
R1761 B.n123 B.n122 10.6151
R1762 B.n126 B.n123 10.6151
R1763 B.n127 B.n126 10.6151
R1764 B.n130 B.n127 10.6151
R1765 B.n131 B.n130 10.6151
R1766 B.n134 B.n131 10.6151
R1767 B.n135 B.n134 10.6151
R1768 B.n138 B.n135 10.6151
R1769 B.n139 B.n138 10.6151
R1770 B.n142 B.n139 10.6151
R1771 B.n143 B.n142 10.6151
R1772 B.n146 B.n143 10.6151
R1773 B.n147 B.n146 10.6151
R1774 B.n150 B.n147 10.6151
R1775 B.n151 B.n150 10.6151
R1776 B.n154 B.n151 10.6151
R1777 B.n155 B.n154 10.6151
R1778 B.n158 B.n155 10.6151
R1779 B.n159 B.n158 10.6151
R1780 B.n162 B.n159 10.6151
R1781 B.n163 B.n162 10.6151
R1782 B.n166 B.n163 10.6151
R1783 B.n167 B.n166 10.6151
R1784 B.n170 B.n167 10.6151
R1785 B.n171 B.n170 10.6151
R1786 B.n174 B.n171 10.6151
R1787 B.n175 B.n174 10.6151
R1788 B.n178 B.n175 10.6151
R1789 B.n179 B.n178 10.6151
R1790 B.n182 B.n179 10.6151
R1791 B.n183 B.n182 10.6151
R1792 B.n186 B.n183 10.6151
R1793 B.n187 B.n186 10.6151
R1794 B.n190 B.n187 10.6151
R1795 B.n191 B.n190 10.6151
R1796 B.n194 B.n191 10.6151
R1797 B.n195 B.n194 10.6151
R1798 B.n199 B.n198 10.6151
R1799 B.n202 B.n199 10.6151
R1800 B.n203 B.n202 10.6151
R1801 B.n206 B.n203 10.6151
R1802 B.n207 B.n206 10.6151
R1803 B.n210 B.n207 10.6151
R1804 B.n211 B.n210 10.6151
R1805 B.n214 B.n211 10.6151
R1806 B.n215 B.n214 10.6151
R1807 B.n219 B.n218 10.6151
R1808 B.n222 B.n219 10.6151
R1809 B.n223 B.n222 10.6151
R1810 B.n226 B.n223 10.6151
R1811 B.n227 B.n226 10.6151
R1812 B.n230 B.n227 10.6151
R1813 B.n231 B.n230 10.6151
R1814 B.n234 B.n231 10.6151
R1815 B.n235 B.n234 10.6151
R1816 B.n238 B.n235 10.6151
R1817 B.n239 B.n238 10.6151
R1818 B.n242 B.n239 10.6151
R1819 B.n243 B.n242 10.6151
R1820 B.n246 B.n243 10.6151
R1821 B.n247 B.n246 10.6151
R1822 B.n250 B.n247 10.6151
R1823 B.n251 B.n250 10.6151
R1824 B.n254 B.n251 10.6151
R1825 B.n255 B.n254 10.6151
R1826 B.n258 B.n255 10.6151
R1827 B.n259 B.n258 10.6151
R1828 B.n262 B.n259 10.6151
R1829 B.n263 B.n262 10.6151
R1830 B.n266 B.n263 10.6151
R1831 B.n267 B.n266 10.6151
R1832 B.n270 B.n267 10.6151
R1833 B.n271 B.n270 10.6151
R1834 B.n274 B.n271 10.6151
R1835 B.n275 B.n274 10.6151
R1836 B.n278 B.n275 10.6151
R1837 B.n279 B.n278 10.6151
R1838 B.n282 B.n279 10.6151
R1839 B.n283 B.n282 10.6151
R1840 B.n286 B.n283 10.6151
R1841 B.n287 B.n286 10.6151
R1842 B.n290 B.n287 10.6151
R1843 B.n291 B.n290 10.6151
R1844 B.n294 B.n291 10.6151
R1845 B.n295 B.n294 10.6151
R1846 B.n298 B.n295 10.6151
R1847 B.n299 B.n298 10.6151
R1848 B.n302 B.n299 10.6151
R1849 B.n303 B.n302 10.6151
R1850 B.n306 B.n303 10.6151
R1851 B.n307 B.n306 10.6151
R1852 B.n310 B.n307 10.6151
R1853 B.n312 B.n310 10.6151
R1854 B.n313 B.n312 10.6151
R1855 B.n711 B.n313 10.6151
R1856 B.n634 B.n344 10.6151
R1857 B.n635 B.n634 10.6151
R1858 B.n636 B.n635 10.6151
R1859 B.n636 B.n337 10.6151
R1860 B.n647 B.n337 10.6151
R1861 B.n648 B.n647 10.6151
R1862 B.n649 B.n648 10.6151
R1863 B.n649 B.n328 10.6151
R1864 B.n659 B.n328 10.6151
R1865 B.n660 B.n659 10.6151
R1866 B.n661 B.n660 10.6151
R1867 B.n661 B.n321 10.6151
R1868 B.n671 B.n321 10.6151
R1869 B.n672 B.n671 10.6151
R1870 B.n674 B.n672 10.6151
R1871 B.n674 B.n673 10.6151
R1872 B.n673 B.n314 10.6151
R1873 B.n686 B.n314 10.6151
R1874 B.n687 B.n686 10.6151
R1875 B.n688 B.n687 10.6151
R1876 B.n689 B.n688 10.6151
R1877 B.n691 B.n689 10.6151
R1878 B.n692 B.n691 10.6151
R1879 B.n693 B.n692 10.6151
R1880 B.n694 B.n693 10.6151
R1881 B.n696 B.n694 10.6151
R1882 B.n697 B.n696 10.6151
R1883 B.n698 B.n697 10.6151
R1884 B.n699 B.n698 10.6151
R1885 B.n701 B.n699 10.6151
R1886 B.n702 B.n701 10.6151
R1887 B.n703 B.n702 10.6151
R1888 B.n704 B.n703 10.6151
R1889 B.n706 B.n704 10.6151
R1890 B.n707 B.n706 10.6151
R1891 B.n708 B.n707 10.6151
R1892 B.n709 B.n708 10.6151
R1893 B.n710 B.n709 10.6151
R1894 B.n628 B.n348 10.6151
R1895 B.n623 B.n348 10.6151
R1896 B.n623 B.n622 10.6151
R1897 B.n622 B.n621 10.6151
R1898 B.n621 B.n618 10.6151
R1899 B.n618 B.n617 10.6151
R1900 B.n617 B.n614 10.6151
R1901 B.n614 B.n613 10.6151
R1902 B.n613 B.n610 10.6151
R1903 B.n610 B.n609 10.6151
R1904 B.n609 B.n606 10.6151
R1905 B.n606 B.n605 10.6151
R1906 B.n605 B.n602 10.6151
R1907 B.n602 B.n601 10.6151
R1908 B.n601 B.n598 10.6151
R1909 B.n598 B.n597 10.6151
R1910 B.n597 B.n594 10.6151
R1911 B.n594 B.n593 10.6151
R1912 B.n593 B.n590 10.6151
R1913 B.n590 B.n589 10.6151
R1914 B.n589 B.n586 10.6151
R1915 B.n586 B.n585 10.6151
R1916 B.n585 B.n582 10.6151
R1917 B.n582 B.n581 10.6151
R1918 B.n581 B.n578 10.6151
R1919 B.n578 B.n577 10.6151
R1920 B.n577 B.n574 10.6151
R1921 B.n574 B.n573 10.6151
R1922 B.n573 B.n570 10.6151
R1923 B.n570 B.n569 10.6151
R1924 B.n569 B.n566 10.6151
R1925 B.n566 B.n565 10.6151
R1926 B.n565 B.n562 10.6151
R1927 B.n562 B.n561 10.6151
R1928 B.n561 B.n558 10.6151
R1929 B.n558 B.n557 10.6151
R1930 B.n557 B.n554 10.6151
R1931 B.n554 B.n553 10.6151
R1932 B.n553 B.n550 10.6151
R1933 B.n550 B.n549 10.6151
R1934 B.n549 B.n546 10.6151
R1935 B.n546 B.n545 10.6151
R1936 B.n545 B.n542 10.6151
R1937 B.n542 B.n541 10.6151
R1938 B.n541 B.n538 10.6151
R1939 B.n538 B.n537 10.6151
R1940 B.n537 B.n534 10.6151
R1941 B.n534 B.n533 10.6151
R1942 B.n533 B.n530 10.6151
R1943 B.n528 B.n525 10.6151
R1944 B.n525 B.n524 10.6151
R1945 B.n524 B.n521 10.6151
R1946 B.n521 B.n520 10.6151
R1947 B.n520 B.n517 10.6151
R1948 B.n517 B.n516 10.6151
R1949 B.n516 B.n513 10.6151
R1950 B.n513 B.n512 10.6151
R1951 B.n512 B.n509 10.6151
R1952 B.n507 B.n504 10.6151
R1953 B.n504 B.n503 10.6151
R1954 B.n503 B.n500 10.6151
R1955 B.n500 B.n499 10.6151
R1956 B.n499 B.n496 10.6151
R1957 B.n496 B.n495 10.6151
R1958 B.n495 B.n492 10.6151
R1959 B.n492 B.n491 10.6151
R1960 B.n491 B.n488 10.6151
R1961 B.n488 B.n487 10.6151
R1962 B.n487 B.n484 10.6151
R1963 B.n484 B.n483 10.6151
R1964 B.n483 B.n480 10.6151
R1965 B.n480 B.n479 10.6151
R1966 B.n479 B.n476 10.6151
R1967 B.n476 B.n475 10.6151
R1968 B.n475 B.n472 10.6151
R1969 B.n472 B.n471 10.6151
R1970 B.n471 B.n468 10.6151
R1971 B.n468 B.n467 10.6151
R1972 B.n467 B.n464 10.6151
R1973 B.n464 B.n463 10.6151
R1974 B.n463 B.n460 10.6151
R1975 B.n460 B.n459 10.6151
R1976 B.n459 B.n456 10.6151
R1977 B.n456 B.n455 10.6151
R1978 B.n455 B.n452 10.6151
R1979 B.n452 B.n451 10.6151
R1980 B.n451 B.n448 10.6151
R1981 B.n448 B.n447 10.6151
R1982 B.n447 B.n444 10.6151
R1983 B.n444 B.n443 10.6151
R1984 B.n443 B.n440 10.6151
R1985 B.n440 B.n439 10.6151
R1986 B.n439 B.n436 10.6151
R1987 B.n436 B.n435 10.6151
R1988 B.n435 B.n432 10.6151
R1989 B.n432 B.n431 10.6151
R1990 B.n431 B.n428 10.6151
R1991 B.n428 B.n427 10.6151
R1992 B.n427 B.n424 10.6151
R1993 B.n424 B.n423 10.6151
R1994 B.n423 B.n420 10.6151
R1995 B.n420 B.n419 10.6151
R1996 B.n419 B.n416 10.6151
R1997 B.n416 B.n415 10.6151
R1998 B.n415 B.n412 10.6151
R1999 B.n412 B.n411 10.6151
R2000 B.n411 B.n409 10.6151
R2001 B.n630 B.n629 10.6151
R2002 B.n630 B.n340 10.6151
R2003 B.n641 B.n340 10.6151
R2004 B.n642 B.n641 10.6151
R2005 B.n643 B.n642 10.6151
R2006 B.n643 B.n333 10.6151
R2007 B.n653 B.n333 10.6151
R2008 B.n654 B.n653 10.6151
R2009 B.n655 B.n654 10.6151
R2010 B.n655 B.n325 10.6151
R2011 B.n665 B.n325 10.6151
R2012 B.n666 B.n665 10.6151
R2013 B.n667 B.n666 10.6151
R2014 B.n667 B.n317 10.6151
R2015 B.n679 B.n317 10.6151
R2016 B.n680 B.n679 10.6151
R2017 B.n681 B.n680 10.6151
R2018 B.n681 B.n0 10.6151
R2019 B.n751 B.n1 10.6151
R2020 B.n751 B.n750 10.6151
R2021 B.n750 B.n749 10.6151
R2022 B.n749 B.n9 10.6151
R2023 B.n743 B.n9 10.6151
R2024 B.n743 B.n742 10.6151
R2025 B.n742 B.n741 10.6151
R2026 B.n741 B.n17 10.6151
R2027 B.n735 B.n17 10.6151
R2028 B.n735 B.n734 10.6151
R2029 B.n734 B.n733 10.6151
R2030 B.n733 B.n24 10.6151
R2031 B.n727 B.n24 10.6151
R2032 B.n727 B.n726 10.6151
R2033 B.n726 B.n725 10.6151
R2034 B.n725 B.n30 10.6151
R2035 B.n719 B.n30 10.6151
R2036 B.n719 B.n718 10.6151
R2037 B.n195 B.n100 9.36635
R2038 B.n218 B.n97 9.36635
R2039 B.n530 B.n529 9.36635
R2040 B.n508 B.n507 9.36635
R2041 B.n645 B.t7 6.54974
R2042 B.n729 B.t14 6.54974
R2043 B.n757 B.n0 2.81026
R2044 B.n757 B.n1 2.81026
R2045 B.n676 B.t0 2.18358
R2046 B.n11 B.t2 2.18358
R2047 B.n198 B.n100 1.24928
R2048 B.n215 B.n97 1.24928
R2049 B.n529 B.n528 1.24928
R2050 B.n509 B.n508 1.24928
R2051 VN.n0 VN.t2 712.841
R2052 VN.n4 VN.t3 712.841
R2053 VN.n1 VN.t1 686.019
R2054 VN.n2 VN.t4 686.019
R2055 VN.n5 VN.t5 686.019
R2056 VN.n6 VN.t0 686.019
R2057 VN.n3 VN.n2 161.3
R2058 VN.n7 VN.n6 161.3
R2059 VN.n2 VN.n1 48.2005
R2060 VN.n6 VN.n5 48.2005
R2061 VN.n7 VN.n4 45.1367
R2062 VN.n3 VN.n0 45.1367
R2063 VN VN.n7 43.3622
R2064 VN.n5 VN.n4 13.3799
R2065 VN.n1 VN.n0 13.3799
R2066 VN VN.n3 0.0516364
R2067 VDD2.n159 VDD2.n83 289.615
R2068 VDD2.n76 VDD2.n0 289.615
R2069 VDD2.n160 VDD2.n159 185
R2070 VDD2.n158 VDD2.n157 185
R2071 VDD2.n87 VDD2.n86 185
R2072 VDD2.n152 VDD2.n151 185
R2073 VDD2.n150 VDD2.n149 185
R2074 VDD2.n91 VDD2.n90 185
R2075 VDD2.n144 VDD2.n143 185
R2076 VDD2.n142 VDD2.n141 185
R2077 VDD2.n95 VDD2.n94 185
R2078 VDD2.n136 VDD2.n135 185
R2079 VDD2.n134 VDD2.n133 185
R2080 VDD2.n132 VDD2.n98 185
R2081 VDD2.n102 VDD2.n99 185
R2082 VDD2.n127 VDD2.n126 185
R2083 VDD2.n125 VDD2.n124 185
R2084 VDD2.n104 VDD2.n103 185
R2085 VDD2.n119 VDD2.n118 185
R2086 VDD2.n117 VDD2.n116 185
R2087 VDD2.n108 VDD2.n107 185
R2088 VDD2.n111 VDD2.n110 185
R2089 VDD2.n27 VDD2.n26 185
R2090 VDD2.n24 VDD2.n23 185
R2091 VDD2.n33 VDD2.n32 185
R2092 VDD2.n35 VDD2.n34 185
R2093 VDD2.n20 VDD2.n19 185
R2094 VDD2.n41 VDD2.n40 185
R2095 VDD2.n44 VDD2.n43 185
R2096 VDD2.n42 VDD2.n16 185
R2097 VDD2.n49 VDD2.n15 185
R2098 VDD2.n51 VDD2.n50 185
R2099 VDD2.n53 VDD2.n52 185
R2100 VDD2.n12 VDD2.n11 185
R2101 VDD2.n59 VDD2.n58 185
R2102 VDD2.n61 VDD2.n60 185
R2103 VDD2.n8 VDD2.n7 185
R2104 VDD2.n67 VDD2.n66 185
R2105 VDD2.n69 VDD2.n68 185
R2106 VDD2.n4 VDD2.n3 185
R2107 VDD2.n75 VDD2.n74 185
R2108 VDD2.n77 VDD2.n76 185
R2109 VDD2.t5 VDD2.n109 149.524
R2110 VDD2.t3 VDD2.n25 149.524
R2111 VDD2.n159 VDD2.n158 104.615
R2112 VDD2.n158 VDD2.n86 104.615
R2113 VDD2.n151 VDD2.n86 104.615
R2114 VDD2.n151 VDD2.n150 104.615
R2115 VDD2.n150 VDD2.n90 104.615
R2116 VDD2.n143 VDD2.n90 104.615
R2117 VDD2.n143 VDD2.n142 104.615
R2118 VDD2.n142 VDD2.n94 104.615
R2119 VDD2.n135 VDD2.n94 104.615
R2120 VDD2.n135 VDD2.n134 104.615
R2121 VDD2.n134 VDD2.n98 104.615
R2122 VDD2.n102 VDD2.n98 104.615
R2123 VDD2.n126 VDD2.n102 104.615
R2124 VDD2.n126 VDD2.n125 104.615
R2125 VDD2.n125 VDD2.n103 104.615
R2126 VDD2.n118 VDD2.n103 104.615
R2127 VDD2.n118 VDD2.n117 104.615
R2128 VDD2.n117 VDD2.n107 104.615
R2129 VDD2.n110 VDD2.n107 104.615
R2130 VDD2.n26 VDD2.n23 104.615
R2131 VDD2.n33 VDD2.n23 104.615
R2132 VDD2.n34 VDD2.n33 104.615
R2133 VDD2.n34 VDD2.n19 104.615
R2134 VDD2.n41 VDD2.n19 104.615
R2135 VDD2.n43 VDD2.n41 104.615
R2136 VDD2.n43 VDD2.n42 104.615
R2137 VDD2.n42 VDD2.n15 104.615
R2138 VDD2.n51 VDD2.n15 104.615
R2139 VDD2.n52 VDD2.n51 104.615
R2140 VDD2.n52 VDD2.n11 104.615
R2141 VDD2.n59 VDD2.n11 104.615
R2142 VDD2.n60 VDD2.n59 104.615
R2143 VDD2.n60 VDD2.n7 104.615
R2144 VDD2.n67 VDD2.n7 104.615
R2145 VDD2.n68 VDD2.n67 104.615
R2146 VDD2.n68 VDD2.n3 104.615
R2147 VDD2.n75 VDD2.n3 104.615
R2148 VDD2.n76 VDD2.n75 104.615
R2149 VDD2.n82 VDD2.n81 59.135
R2150 VDD2 VDD2.n165 59.1323
R2151 VDD2.n110 VDD2.t5 52.3082
R2152 VDD2.n26 VDD2.t3 52.3082
R2153 VDD2.n82 VDD2.n80 47.0699
R2154 VDD2.n164 VDD2.n163 46.5369
R2155 VDD2.n164 VDD2.n82 39.0924
R2156 VDD2.n133 VDD2.n132 13.1884
R2157 VDD2.n50 VDD2.n49 13.1884
R2158 VDD2.n136 VDD2.n97 12.8005
R2159 VDD2.n131 VDD2.n99 12.8005
R2160 VDD2.n48 VDD2.n16 12.8005
R2161 VDD2.n53 VDD2.n14 12.8005
R2162 VDD2.n137 VDD2.n95 12.0247
R2163 VDD2.n128 VDD2.n127 12.0247
R2164 VDD2.n45 VDD2.n44 12.0247
R2165 VDD2.n54 VDD2.n12 12.0247
R2166 VDD2.n141 VDD2.n140 11.249
R2167 VDD2.n124 VDD2.n101 11.249
R2168 VDD2.n40 VDD2.n18 11.249
R2169 VDD2.n58 VDD2.n57 11.249
R2170 VDD2.n144 VDD2.n93 10.4732
R2171 VDD2.n123 VDD2.n104 10.4732
R2172 VDD2.n39 VDD2.n20 10.4732
R2173 VDD2.n61 VDD2.n10 10.4732
R2174 VDD2.n111 VDD2.n109 10.2747
R2175 VDD2.n27 VDD2.n25 10.2747
R2176 VDD2.n145 VDD2.n91 9.69747
R2177 VDD2.n120 VDD2.n119 9.69747
R2178 VDD2.n36 VDD2.n35 9.69747
R2179 VDD2.n62 VDD2.n8 9.69747
R2180 VDD2.n163 VDD2.n162 9.45567
R2181 VDD2.n80 VDD2.n79 9.45567
R2182 VDD2.n113 VDD2.n112 9.3005
R2183 VDD2.n115 VDD2.n114 9.3005
R2184 VDD2.n106 VDD2.n105 9.3005
R2185 VDD2.n121 VDD2.n120 9.3005
R2186 VDD2.n123 VDD2.n122 9.3005
R2187 VDD2.n101 VDD2.n100 9.3005
R2188 VDD2.n129 VDD2.n128 9.3005
R2189 VDD2.n131 VDD2.n130 9.3005
R2190 VDD2.n85 VDD2.n84 9.3005
R2191 VDD2.n162 VDD2.n161 9.3005
R2192 VDD2.n156 VDD2.n155 9.3005
R2193 VDD2.n154 VDD2.n153 9.3005
R2194 VDD2.n89 VDD2.n88 9.3005
R2195 VDD2.n148 VDD2.n147 9.3005
R2196 VDD2.n146 VDD2.n145 9.3005
R2197 VDD2.n93 VDD2.n92 9.3005
R2198 VDD2.n140 VDD2.n139 9.3005
R2199 VDD2.n138 VDD2.n137 9.3005
R2200 VDD2.n97 VDD2.n96 9.3005
R2201 VDD2.n73 VDD2.n72 9.3005
R2202 VDD2.n2 VDD2.n1 9.3005
R2203 VDD2.n79 VDD2.n78 9.3005
R2204 VDD2.n6 VDD2.n5 9.3005
R2205 VDD2.n65 VDD2.n64 9.3005
R2206 VDD2.n63 VDD2.n62 9.3005
R2207 VDD2.n10 VDD2.n9 9.3005
R2208 VDD2.n57 VDD2.n56 9.3005
R2209 VDD2.n55 VDD2.n54 9.3005
R2210 VDD2.n14 VDD2.n13 9.3005
R2211 VDD2.n29 VDD2.n28 9.3005
R2212 VDD2.n31 VDD2.n30 9.3005
R2213 VDD2.n22 VDD2.n21 9.3005
R2214 VDD2.n37 VDD2.n36 9.3005
R2215 VDD2.n39 VDD2.n38 9.3005
R2216 VDD2.n18 VDD2.n17 9.3005
R2217 VDD2.n46 VDD2.n45 9.3005
R2218 VDD2.n48 VDD2.n47 9.3005
R2219 VDD2.n71 VDD2.n70 9.3005
R2220 VDD2.n163 VDD2.n83 8.92171
R2221 VDD2.n149 VDD2.n148 8.92171
R2222 VDD2.n116 VDD2.n106 8.92171
R2223 VDD2.n32 VDD2.n22 8.92171
R2224 VDD2.n66 VDD2.n65 8.92171
R2225 VDD2.n80 VDD2.n0 8.92171
R2226 VDD2.n161 VDD2.n160 8.14595
R2227 VDD2.n152 VDD2.n89 8.14595
R2228 VDD2.n115 VDD2.n108 8.14595
R2229 VDD2.n31 VDD2.n24 8.14595
R2230 VDD2.n69 VDD2.n6 8.14595
R2231 VDD2.n78 VDD2.n77 8.14595
R2232 VDD2.n157 VDD2.n85 7.3702
R2233 VDD2.n153 VDD2.n87 7.3702
R2234 VDD2.n112 VDD2.n111 7.3702
R2235 VDD2.n28 VDD2.n27 7.3702
R2236 VDD2.n70 VDD2.n4 7.3702
R2237 VDD2.n74 VDD2.n2 7.3702
R2238 VDD2.n157 VDD2.n156 6.59444
R2239 VDD2.n156 VDD2.n87 6.59444
R2240 VDD2.n73 VDD2.n4 6.59444
R2241 VDD2.n74 VDD2.n73 6.59444
R2242 VDD2.n160 VDD2.n85 5.81868
R2243 VDD2.n153 VDD2.n152 5.81868
R2244 VDD2.n112 VDD2.n108 5.81868
R2245 VDD2.n28 VDD2.n24 5.81868
R2246 VDD2.n70 VDD2.n69 5.81868
R2247 VDD2.n77 VDD2.n2 5.81868
R2248 VDD2.n161 VDD2.n83 5.04292
R2249 VDD2.n149 VDD2.n89 5.04292
R2250 VDD2.n116 VDD2.n115 5.04292
R2251 VDD2.n32 VDD2.n31 5.04292
R2252 VDD2.n66 VDD2.n6 5.04292
R2253 VDD2.n78 VDD2.n0 5.04292
R2254 VDD2.n148 VDD2.n91 4.26717
R2255 VDD2.n119 VDD2.n106 4.26717
R2256 VDD2.n35 VDD2.n22 4.26717
R2257 VDD2.n65 VDD2.n8 4.26717
R2258 VDD2.n145 VDD2.n144 3.49141
R2259 VDD2.n120 VDD2.n104 3.49141
R2260 VDD2.n36 VDD2.n20 3.49141
R2261 VDD2.n62 VDD2.n61 3.49141
R2262 VDD2.n29 VDD2.n25 2.84303
R2263 VDD2.n113 VDD2.n109 2.84303
R2264 VDD2.n141 VDD2.n93 2.71565
R2265 VDD2.n124 VDD2.n123 2.71565
R2266 VDD2.n40 VDD2.n39 2.71565
R2267 VDD2.n58 VDD2.n10 2.71565
R2268 VDD2.n140 VDD2.n95 1.93989
R2269 VDD2.n127 VDD2.n101 1.93989
R2270 VDD2.n44 VDD2.n18 1.93989
R2271 VDD2.n57 VDD2.n12 1.93989
R2272 VDD2.n165 VDD2.t0 1.33115
R2273 VDD2.n165 VDD2.t2 1.33115
R2274 VDD2.n81 VDD2.t4 1.33115
R2275 VDD2.n81 VDD2.t1 1.33115
R2276 VDD2.n137 VDD2.n136 1.16414
R2277 VDD2.n128 VDD2.n99 1.16414
R2278 VDD2.n45 VDD2.n16 1.16414
R2279 VDD2.n54 VDD2.n53 1.16414
R2280 VDD2 VDD2.n164 0.647052
R2281 VDD2.n133 VDD2.n97 0.388379
R2282 VDD2.n132 VDD2.n131 0.388379
R2283 VDD2.n49 VDD2.n48 0.388379
R2284 VDD2.n50 VDD2.n14 0.388379
R2285 VDD2.n162 VDD2.n84 0.155672
R2286 VDD2.n155 VDD2.n84 0.155672
R2287 VDD2.n155 VDD2.n154 0.155672
R2288 VDD2.n154 VDD2.n88 0.155672
R2289 VDD2.n147 VDD2.n88 0.155672
R2290 VDD2.n147 VDD2.n146 0.155672
R2291 VDD2.n146 VDD2.n92 0.155672
R2292 VDD2.n139 VDD2.n92 0.155672
R2293 VDD2.n139 VDD2.n138 0.155672
R2294 VDD2.n138 VDD2.n96 0.155672
R2295 VDD2.n130 VDD2.n96 0.155672
R2296 VDD2.n130 VDD2.n129 0.155672
R2297 VDD2.n129 VDD2.n100 0.155672
R2298 VDD2.n122 VDD2.n100 0.155672
R2299 VDD2.n122 VDD2.n121 0.155672
R2300 VDD2.n121 VDD2.n105 0.155672
R2301 VDD2.n114 VDD2.n105 0.155672
R2302 VDD2.n114 VDD2.n113 0.155672
R2303 VDD2.n30 VDD2.n29 0.155672
R2304 VDD2.n30 VDD2.n21 0.155672
R2305 VDD2.n37 VDD2.n21 0.155672
R2306 VDD2.n38 VDD2.n37 0.155672
R2307 VDD2.n38 VDD2.n17 0.155672
R2308 VDD2.n46 VDD2.n17 0.155672
R2309 VDD2.n47 VDD2.n46 0.155672
R2310 VDD2.n47 VDD2.n13 0.155672
R2311 VDD2.n55 VDD2.n13 0.155672
R2312 VDD2.n56 VDD2.n55 0.155672
R2313 VDD2.n56 VDD2.n9 0.155672
R2314 VDD2.n63 VDD2.n9 0.155672
R2315 VDD2.n64 VDD2.n63 0.155672
R2316 VDD2.n64 VDD2.n5 0.155672
R2317 VDD2.n71 VDD2.n5 0.155672
R2318 VDD2.n72 VDD2.n71 0.155672
R2319 VDD2.n72 VDD2.n1 0.155672
R2320 VDD2.n79 VDD2.n1 0.155672
C0 VDD2 VTAIL 12.838401f
C1 VTAIL VDD1 12.8073f
C2 VDD2 VDD1 0.669141f
C3 VN VTAIL 4.34075f
C4 VDD2 VN 4.80607f
C5 VN VDD1 0.148366f
C6 VP VTAIL 4.35553f
C7 VDD2 VP 0.288362f
C8 VP VDD1 4.94031f
C9 VP VN 5.49371f
C10 VDD2 B 4.926055f
C11 VDD1 B 4.923352f
C12 VTAIL B 7.326048f
C13 VN B 7.8083f
C14 VP B 5.593132f
C15 VDD2.n0 B 0.034443f
C16 VDD2.n1 B 0.024043f
C17 VDD2.n2 B 0.012919f
C18 VDD2.n3 B 0.030537f
C19 VDD2.n4 B 0.013679f
C20 VDD2.n5 B 0.024043f
C21 VDD2.n6 B 0.012919f
C22 VDD2.n7 B 0.030537f
C23 VDD2.n8 B 0.013679f
C24 VDD2.n9 B 0.024043f
C25 VDD2.n10 B 0.012919f
C26 VDD2.n11 B 0.030537f
C27 VDD2.n12 B 0.013679f
C28 VDD2.n13 B 0.024043f
C29 VDD2.n14 B 0.012919f
C30 VDD2.n15 B 0.030537f
C31 VDD2.n16 B 0.013679f
C32 VDD2.n17 B 0.024043f
C33 VDD2.n18 B 0.012919f
C34 VDD2.n19 B 0.030537f
C35 VDD2.n20 B 0.013679f
C36 VDD2.n21 B 0.024043f
C37 VDD2.n22 B 0.012919f
C38 VDD2.n23 B 0.030537f
C39 VDD2.n24 B 0.013679f
C40 VDD2.n25 B 0.199928f
C41 VDD2.t3 B 0.051947f
C42 VDD2.n26 B 0.022903f
C43 VDD2.n27 B 0.021587f
C44 VDD2.n28 B 0.012919f
C45 VDD2.n29 B 1.52089f
C46 VDD2.n30 B 0.024043f
C47 VDD2.n31 B 0.012919f
C48 VDD2.n32 B 0.013679f
C49 VDD2.n33 B 0.030537f
C50 VDD2.n34 B 0.030537f
C51 VDD2.n35 B 0.013679f
C52 VDD2.n36 B 0.012919f
C53 VDD2.n37 B 0.024043f
C54 VDD2.n38 B 0.024043f
C55 VDD2.n39 B 0.012919f
C56 VDD2.n40 B 0.013679f
C57 VDD2.n41 B 0.030537f
C58 VDD2.n42 B 0.030537f
C59 VDD2.n43 B 0.030537f
C60 VDD2.n44 B 0.013679f
C61 VDD2.n45 B 0.012919f
C62 VDD2.n46 B 0.024043f
C63 VDD2.n47 B 0.024043f
C64 VDD2.n48 B 0.012919f
C65 VDD2.n49 B 0.013299f
C66 VDD2.n50 B 0.013299f
C67 VDD2.n51 B 0.030537f
C68 VDD2.n52 B 0.030537f
C69 VDD2.n53 B 0.013679f
C70 VDD2.n54 B 0.012919f
C71 VDD2.n55 B 0.024043f
C72 VDD2.n56 B 0.024043f
C73 VDD2.n57 B 0.012919f
C74 VDD2.n58 B 0.013679f
C75 VDD2.n59 B 0.030537f
C76 VDD2.n60 B 0.030537f
C77 VDD2.n61 B 0.013679f
C78 VDD2.n62 B 0.012919f
C79 VDD2.n63 B 0.024043f
C80 VDD2.n64 B 0.024043f
C81 VDD2.n65 B 0.012919f
C82 VDD2.n66 B 0.013679f
C83 VDD2.n67 B 0.030537f
C84 VDD2.n68 B 0.030537f
C85 VDD2.n69 B 0.013679f
C86 VDD2.n70 B 0.012919f
C87 VDD2.n71 B 0.024043f
C88 VDD2.n72 B 0.024043f
C89 VDD2.n73 B 0.012919f
C90 VDD2.n74 B 0.013679f
C91 VDD2.n75 B 0.030537f
C92 VDD2.n76 B 0.067255f
C93 VDD2.n77 B 0.013679f
C94 VDD2.n78 B 0.012919f
C95 VDD2.n79 B 0.051632f
C96 VDD2.n80 B 0.055238f
C97 VDD2.t4 B 0.282708f
C98 VDD2.t1 B 0.282708f
C99 VDD2.n81 B 2.54632f
C100 VDD2.n82 B 1.90589f
C101 VDD2.n83 B 0.034443f
C102 VDD2.n84 B 0.024043f
C103 VDD2.n85 B 0.012919f
C104 VDD2.n86 B 0.030537f
C105 VDD2.n87 B 0.013679f
C106 VDD2.n88 B 0.024043f
C107 VDD2.n89 B 0.012919f
C108 VDD2.n90 B 0.030537f
C109 VDD2.n91 B 0.013679f
C110 VDD2.n92 B 0.024043f
C111 VDD2.n93 B 0.012919f
C112 VDD2.n94 B 0.030537f
C113 VDD2.n95 B 0.013679f
C114 VDD2.n96 B 0.024043f
C115 VDD2.n97 B 0.012919f
C116 VDD2.n98 B 0.030537f
C117 VDD2.n99 B 0.013679f
C118 VDD2.n100 B 0.024043f
C119 VDD2.n101 B 0.012919f
C120 VDD2.n102 B 0.030537f
C121 VDD2.n103 B 0.030537f
C122 VDD2.n104 B 0.013679f
C123 VDD2.n105 B 0.024043f
C124 VDD2.n106 B 0.012919f
C125 VDD2.n107 B 0.030537f
C126 VDD2.n108 B 0.013679f
C127 VDD2.n109 B 0.199928f
C128 VDD2.t5 B 0.051947f
C129 VDD2.n110 B 0.022903f
C130 VDD2.n111 B 0.021587f
C131 VDD2.n112 B 0.012919f
C132 VDD2.n113 B 1.52089f
C133 VDD2.n114 B 0.024043f
C134 VDD2.n115 B 0.012919f
C135 VDD2.n116 B 0.013679f
C136 VDD2.n117 B 0.030537f
C137 VDD2.n118 B 0.030537f
C138 VDD2.n119 B 0.013679f
C139 VDD2.n120 B 0.012919f
C140 VDD2.n121 B 0.024043f
C141 VDD2.n122 B 0.024043f
C142 VDD2.n123 B 0.012919f
C143 VDD2.n124 B 0.013679f
C144 VDD2.n125 B 0.030537f
C145 VDD2.n126 B 0.030537f
C146 VDD2.n127 B 0.013679f
C147 VDD2.n128 B 0.012919f
C148 VDD2.n129 B 0.024043f
C149 VDD2.n130 B 0.024043f
C150 VDD2.n131 B 0.012919f
C151 VDD2.n132 B 0.013299f
C152 VDD2.n133 B 0.013299f
C153 VDD2.n134 B 0.030537f
C154 VDD2.n135 B 0.030537f
C155 VDD2.n136 B 0.013679f
C156 VDD2.n137 B 0.012919f
C157 VDD2.n138 B 0.024043f
C158 VDD2.n139 B 0.024043f
C159 VDD2.n140 B 0.012919f
C160 VDD2.n141 B 0.013679f
C161 VDD2.n142 B 0.030537f
C162 VDD2.n143 B 0.030537f
C163 VDD2.n144 B 0.013679f
C164 VDD2.n145 B 0.012919f
C165 VDD2.n146 B 0.024043f
C166 VDD2.n147 B 0.024043f
C167 VDD2.n148 B 0.012919f
C168 VDD2.n149 B 0.013679f
C169 VDD2.n150 B 0.030537f
C170 VDD2.n151 B 0.030537f
C171 VDD2.n152 B 0.013679f
C172 VDD2.n153 B 0.012919f
C173 VDD2.n154 B 0.024043f
C174 VDD2.n155 B 0.024043f
C175 VDD2.n156 B 0.012919f
C176 VDD2.n157 B 0.013679f
C177 VDD2.n158 B 0.030537f
C178 VDD2.n159 B 0.067255f
C179 VDD2.n160 B 0.013679f
C180 VDD2.n161 B 0.012919f
C181 VDD2.n162 B 0.051632f
C182 VDD2.n163 B 0.054259f
C183 VDD2.n164 B 2.14717f
C184 VDD2.t0 B 0.282708f
C185 VDD2.t2 B 0.282708f
C186 VDD2.n165 B 2.54631f
C187 VN.t2 B 1.21396f
C188 VN.n0 B 0.448398f
C189 VN.t1 B 1.19646f
C190 VN.n1 B 0.475933f
C191 VN.t4 B 1.19646f
C192 VN.n2 B 0.464864f
C193 VN.n3 B 0.195142f
C194 VN.t3 B 1.21396f
C195 VN.n4 B 0.448398f
C196 VN.t5 B 1.19646f
C197 VN.n5 B 0.475933f
C198 VN.t0 B 1.19646f
C199 VN.n6 B 0.464864f
C200 VN.n7 B 2.28116f
C201 VTAIL.t2 B 0.289518f
C202 VTAIL.t1 B 0.289518f
C203 VTAIL.n0 B 2.52583f
C204 VTAIL.n1 B 0.346737f
C205 VTAIL.n2 B 0.035273f
C206 VTAIL.n3 B 0.024622f
C207 VTAIL.n4 B 0.013231f
C208 VTAIL.n5 B 0.031273f
C209 VTAIL.n6 B 0.014009f
C210 VTAIL.n7 B 0.024622f
C211 VTAIL.n8 B 0.013231f
C212 VTAIL.n9 B 0.031273f
C213 VTAIL.n10 B 0.014009f
C214 VTAIL.n11 B 0.024622f
C215 VTAIL.n12 B 0.013231f
C216 VTAIL.n13 B 0.031273f
C217 VTAIL.n14 B 0.014009f
C218 VTAIL.n15 B 0.024622f
C219 VTAIL.n16 B 0.013231f
C220 VTAIL.n17 B 0.031273f
C221 VTAIL.n18 B 0.014009f
C222 VTAIL.n19 B 0.024622f
C223 VTAIL.n20 B 0.013231f
C224 VTAIL.n21 B 0.031273f
C225 VTAIL.n22 B 0.014009f
C226 VTAIL.n23 B 0.024622f
C227 VTAIL.n24 B 0.013231f
C228 VTAIL.n25 B 0.031273f
C229 VTAIL.n26 B 0.014009f
C230 VTAIL.n27 B 0.204744f
C231 VTAIL.t8 B 0.053199f
C232 VTAIL.n28 B 0.023454f
C233 VTAIL.n29 B 0.022107f
C234 VTAIL.n30 B 0.013231f
C235 VTAIL.n31 B 1.55753f
C236 VTAIL.n32 B 0.024622f
C237 VTAIL.n33 B 0.013231f
C238 VTAIL.n34 B 0.014009f
C239 VTAIL.n35 B 0.031273f
C240 VTAIL.n36 B 0.031273f
C241 VTAIL.n37 B 0.014009f
C242 VTAIL.n38 B 0.013231f
C243 VTAIL.n39 B 0.024622f
C244 VTAIL.n40 B 0.024622f
C245 VTAIL.n41 B 0.013231f
C246 VTAIL.n42 B 0.014009f
C247 VTAIL.n43 B 0.031273f
C248 VTAIL.n44 B 0.031273f
C249 VTAIL.n45 B 0.031273f
C250 VTAIL.n46 B 0.014009f
C251 VTAIL.n47 B 0.013231f
C252 VTAIL.n48 B 0.024622f
C253 VTAIL.n49 B 0.024622f
C254 VTAIL.n50 B 0.013231f
C255 VTAIL.n51 B 0.01362f
C256 VTAIL.n52 B 0.01362f
C257 VTAIL.n53 B 0.031273f
C258 VTAIL.n54 B 0.031273f
C259 VTAIL.n55 B 0.014009f
C260 VTAIL.n56 B 0.013231f
C261 VTAIL.n57 B 0.024622f
C262 VTAIL.n58 B 0.024622f
C263 VTAIL.n59 B 0.013231f
C264 VTAIL.n60 B 0.014009f
C265 VTAIL.n61 B 0.031273f
C266 VTAIL.n62 B 0.031273f
C267 VTAIL.n63 B 0.014009f
C268 VTAIL.n64 B 0.013231f
C269 VTAIL.n65 B 0.024622f
C270 VTAIL.n66 B 0.024622f
C271 VTAIL.n67 B 0.013231f
C272 VTAIL.n68 B 0.014009f
C273 VTAIL.n69 B 0.031273f
C274 VTAIL.n70 B 0.031273f
C275 VTAIL.n71 B 0.014009f
C276 VTAIL.n72 B 0.013231f
C277 VTAIL.n73 B 0.024622f
C278 VTAIL.n74 B 0.024622f
C279 VTAIL.n75 B 0.013231f
C280 VTAIL.n76 B 0.014009f
C281 VTAIL.n77 B 0.031273f
C282 VTAIL.n78 B 0.068875f
C283 VTAIL.n79 B 0.014009f
C284 VTAIL.n80 B 0.013231f
C285 VTAIL.n81 B 0.052876f
C286 VTAIL.n82 B 0.03853f
C287 VTAIL.n83 B 0.149387f
C288 VTAIL.t6 B 0.289518f
C289 VTAIL.t11 B 0.289518f
C290 VTAIL.n84 B 2.52583f
C291 VTAIL.n85 B 1.79704f
C292 VTAIL.t3 B 0.289518f
C293 VTAIL.t4 B 0.289518f
C294 VTAIL.n86 B 2.52584f
C295 VTAIL.n87 B 1.79703f
C296 VTAIL.n88 B 0.035273f
C297 VTAIL.n89 B 0.024622f
C298 VTAIL.n90 B 0.013231f
C299 VTAIL.n91 B 0.031273f
C300 VTAIL.n92 B 0.014009f
C301 VTAIL.n93 B 0.024622f
C302 VTAIL.n94 B 0.013231f
C303 VTAIL.n95 B 0.031273f
C304 VTAIL.n96 B 0.014009f
C305 VTAIL.n97 B 0.024622f
C306 VTAIL.n98 B 0.013231f
C307 VTAIL.n99 B 0.031273f
C308 VTAIL.n100 B 0.014009f
C309 VTAIL.n101 B 0.024622f
C310 VTAIL.n102 B 0.013231f
C311 VTAIL.n103 B 0.031273f
C312 VTAIL.n104 B 0.014009f
C313 VTAIL.n105 B 0.024622f
C314 VTAIL.n106 B 0.013231f
C315 VTAIL.n107 B 0.031273f
C316 VTAIL.n108 B 0.031273f
C317 VTAIL.n109 B 0.014009f
C318 VTAIL.n110 B 0.024622f
C319 VTAIL.n111 B 0.013231f
C320 VTAIL.n112 B 0.031273f
C321 VTAIL.n113 B 0.014009f
C322 VTAIL.n114 B 0.204744f
C323 VTAIL.t0 B 0.053199f
C324 VTAIL.n115 B 0.023454f
C325 VTAIL.n116 B 0.022107f
C326 VTAIL.n117 B 0.013231f
C327 VTAIL.n118 B 1.55753f
C328 VTAIL.n119 B 0.024622f
C329 VTAIL.n120 B 0.013231f
C330 VTAIL.n121 B 0.014009f
C331 VTAIL.n122 B 0.031273f
C332 VTAIL.n123 B 0.031273f
C333 VTAIL.n124 B 0.014009f
C334 VTAIL.n125 B 0.013231f
C335 VTAIL.n126 B 0.024622f
C336 VTAIL.n127 B 0.024622f
C337 VTAIL.n128 B 0.013231f
C338 VTAIL.n129 B 0.014009f
C339 VTAIL.n130 B 0.031273f
C340 VTAIL.n131 B 0.031273f
C341 VTAIL.n132 B 0.014009f
C342 VTAIL.n133 B 0.013231f
C343 VTAIL.n134 B 0.024622f
C344 VTAIL.n135 B 0.024622f
C345 VTAIL.n136 B 0.013231f
C346 VTAIL.n137 B 0.01362f
C347 VTAIL.n138 B 0.01362f
C348 VTAIL.n139 B 0.031273f
C349 VTAIL.n140 B 0.031273f
C350 VTAIL.n141 B 0.014009f
C351 VTAIL.n142 B 0.013231f
C352 VTAIL.n143 B 0.024622f
C353 VTAIL.n144 B 0.024622f
C354 VTAIL.n145 B 0.013231f
C355 VTAIL.n146 B 0.014009f
C356 VTAIL.n147 B 0.031273f
C357 VTAIL.n148 B 0.031273f
C358 VTAIL.n149 B 0.014009f
C359 VTAIL.n150 B 0.013231f
C360 VTAIL.n151 B 0.024622f
C361 VTAIL.n152 B 0.024622f
C362 VTAIL.n153 B 0.013231f
C363 VTAIL.n154 B 0.014009f
C364 VTAIL.n155 B 0.031273f
C365 VTAIL.n156 B 0.031273f
C366 VTAIL.n157 B 0.014009f
C367 VTAIL.n158 B 0.013231f
C368 VTAIL.n159 B 0.024622f
C369 VTAIL.n160 B 0.024622f
C370 VTAIL.n161 B 0.013231f
C371 VTAIL.n162 B 0.014009f
C372 VTAIL.n163 B 0.031273f
C373 VTAIL.n164 B 0.068875f
C374 VTAIL.n165 B 0.014009f
C375 VTAIL.n166 B 0.013231f
C376 VTAIL.n167 B 0.052876f
C377 VTAIL.n168 B 0.03853f
C378 VTAIL.n169 B 0.149387f
C379 VTAIL.t10 B 0.289518f
C380 VTAIL.t9 B 0.289518f
C381 VTAIL.n170 B 2.52584f
C382 VTAIL.n171 B 0.388786f
C383 VTAIL.n172 B 0.035273f
C384 VTAIL.n173 B 0.024622f
C385 VTAIL.n174 B 0.013231f
C386 VTAIL.n175 B 0.031273f
C387 VTAIL.n176 B 0.014009f
C388 VTAIL.n177 B 0.024622f
C389 VTAIL.n178 B 0.013231f
C390 VTAIL.n179 B 0.031273f
C391 VTAIL.n180 B 0.014009f
C392 VTAIL.n181 B 0.024622f
C393 VTAIL.n182 B 0.013231f
C394 VTAIL.n183 B 0.031273f
C395 VTAIL.n184 B 0.014009f
C396 VTAIL.n185 B 0.024622f
C397 VTAIL.n186 B 0.013231f
C398 VTAIL.n187 B 0.031273f
C399 VTAIL.n188 B 0.014009f
C400 VTAIL.n189 B 0.024622f
C401 VTAIL.n190 B 0.013231f
C402 VTAIL.n191 B 0.031273f
C403 VTAIL.n192 B 0.031273f
C404 VTAIL.n193 B 0.014009f
C405 VTAIL.n194 B 0.024622f
C406 VTAIL.n195 B 0.013231f
C407 VTAIL.n196 B 0.031273f
C408 VTAIL.n197 B 0.014009f
C409 VTAIL.n198 B 0.204744f
C410 VTAIL.t7 B 0.053199f
C411 VTAIL.n199 B 0.023454f
C412 VTAIL.n200 B 0.022107f
C413 VTAIL.n201 B 0.013231f
C414 VTAIL.n202 B 1.55753f
C415 VTAIL.n203 B 0.024622f
C416 VTAIL.n204 B 0.013231f
C417 VTAIL.n205 B 0.014009f
C418 VTAIL.n206 B 0.031273f
C419 VTAIL.n207 B 0.031273f
C420 VTAIL.n208 B 0.014009f
C421 VTAIL.n209 B 0.013231f
C422 VTAIL.n210 B 0.024622f
C423 VTAIL.n211 B 0.024622f
C424 VTAIL.n212 B 0.013231f
C425 VTAIL.n213 B 0.014009f
C426 VTAIL.n214 B 0.031273f
C427 VTAIL.n215 B 0.031273f
C428 VTAIL.n216 B 0.014009f
C429 VTAIL.n217 B 0.013231f
C430 VTAIL.n218 B 0.024622f
C431 VTAIL.n219 B 0.024622f
C432 VTAIL.n220 B 0.013231f
C433 VTAIL.n221 B 0.01362f
C434 VTAIL.n222 B 0.01362f
C435 VTAIL.n223 B 0.031273f
C436 VTAIL.n224 B 0.031273f
C437 VTAIL.n225 B 0.014009f
C438 VTAIL.n226 B 0.013231f
C439 VTAIL.n227 B 0.024622f
C440 VTAIL.n228 B 0.024622f
C441 VTAIL.n229 B 0.013231f
C442 VTAIL.n230 B 0.014009f
C443 VTAIL.n231 B 0.031273f
C444 VTAIL.n232 B 0.031273f
C445 VTAIL.n233 B 0.014009f
C446 VTAIL.n234 B 0.013231f
C447 VTAIL.n235 B 0.024622f
C448 VTAIL.n236 B 0.024622f
C449 VTAIL.n237 B 0.013231f
C450 VTAIL.n238 B 0.014009f
C451 VTAIL.n239 B 0.031273f
C452 VTAIL.n240 B 0.031273f
C453 VTAIL.n241 B 0.014009f
C454 VTAIL.n242 B 0.013231f
C455 VTAIL.n243 B 0.024622f
C456 VTAIL.n244 B 0.024622f
C457 VTAIL.n245 B 0.013231f
C458 VTAIL.n246 B 0.014009f
C459 VTAIL.n247 B 0.031273f
C460 VTAIL.n248 B 0.068875f
C461 VTAIL.n249 B 0.014009f
C462 VTAIL.n250 B 0.013231f
C463 VTAIL.n251 B 0.052876f
C464 VTAIL.n252 B 0.03853f
C465 VTAIL.n253 B 1.49539f
C466 VTAIL.n254 B 0.035273f
C467 VTAIL.n255 B 0.024622f
C468 VTAIL.n256 B 0.013231f
C469 VTAIL.n257 B 0.031273f
C470 VTAIL.n258 B 0.014009f
C471 VTAIL.n259 B 0.024622f
C472 VTAIL.n260 B 0.013231f
C473 VTAIL.n261 B 0.031273f
C474 VTAIL.n262 B 0.014009f
C475 VTAIL.n263 B 0.024622f
C476 VTAIL.n264 B 0.013231f
C477 VTAIL.n265 B 0.031273f
C478 VTAIL.n266 B 0.014009f
C479 VTAIL.n267 B 0.024622f
C480 VTAIL.n268 B 0.013231f
C481 VTAIL.n269 B 0.031273f
C482 VTAIL.n270 B 0.014009f
C483 VTAIL.n271 B 0.024622f
C484 VTAIL.n272 B 0.013231f
C485 VTAIL.n273 B 0.031273f
C486 VTAIL.n274 B 0.014009f
C487 VTAIL.n275 B 0.024622f
C488 VTAIL.n276 B 0.013231f
C489 VTAIL.n277 B 0.031273f
C490 VTAIL.n278 B 0.014009f
C491 VTAIL.n279 B 0.204744f
C492 VTAIL.t5 B 0.053199f
C493 VTAIL.n280 B 0.023454f
C494 VTAIL.n281 B 0.022107f
C495 VTAIL.n282 B 0.013231f
C496 VTAIL.n283 B 1.55753f
C497 VTAIL.n284 B 0.024622f
C498 VTAIL.n285 B 0.013231f
C499 VTAIL.n286 B 0.014009f
C500 VTAIL.n287 B 0.031273f
C501 VTAIL.n288 B 0.031273f
C502 VTAIL.n289 B 0.014009f
C503 VTAIL.n290 B 0.013231f
C504 VTAIL.n291 B 0.024622f
C505 VTAIL.n292 B 0.024622f
C506 VTAIL.n293 B 0.013231f
C507 VTAIL.n294 B 0.014009f
C508 VTAIL.n295 B 0.031273f
C509 VTAIL.n296 B 0.031273f
C510 VTAIL.n297 B 0.031273f
C511 VTAIL.n298 B 0.014009f
C512 VTAIL.n299 B 0.013231f
C513 VTAIL.n300 B 0.024622f
C514 VTAIL.n301 B 0.024622f
C515 VTAIL.n302 B 0.013231f
C516 VTAIL.n303 B 0.01362f
C517 VTAIL.n304 B 0.01362f
C518 VTAIL.n305 B 0.031273f
C519 VTAIL.n306 B 0.031273f
C520 VTAIL.n307 B 0.014009f
C521 VTAIL.n308 B 0.013231f
C522 VTAIL.n309 B 0.024622f
C523 VTAIL.n310 B 0.024622f
C524 VTAIL.n311 B 0.013231f
C525 VTAIL.n312 B 0.014009f
C526 VTAIL.n313 B 0.031273f
C527 VTAIL.n314 B 0.031273f
C528 VTAIL.n315 B 0.014009f
C529 VTAIL.n316 B 0.013231f
C530 VTAIL.n317 B 0.024622f
C531 VTAIL.n318 B 0.024622f
C532 VTAIL.n319 B 0.013231f
C533 VTAIL.n320 B 0.014009f
C534 VTAIL.n321 B 0.031273f
C535 VTAIL.n322 B 0.031273f
C536 VTAIL.n323 B 0.014009f
C537 VTAIL.n324 B 0.013231f
C538 VTAIL.n325 B 0.024622f
C539 VTAIL.n326 B 0.024622f
C540 VTAIL.n327 B 0.013231f
C541 VTAIL.n328 B 0.014009f
C542 VTAIL.n329 B 0.031273f
C543 VTAIL.n330 B 0.068875f
C544 VTAIL.n331 B 0.014009f
C545 VTAIL.n332 B 0.013231f
C546 VTAIL.n333 B 0.052876f
C547 VTAIL.n334 B 0.03853f
C548 VTAIL.n335 B 1.47521f
C549 VDD1.n0 B 0.034465f
C550 VDD1.n1 B 0.024058f
C551 VDD1.n2 B 0.012928f
C552 VDD1.n3 B 0.030556f
C553 VDD1.n4 B 0.013688f
C554 VDD1.n5 B 0.024058f
C555 VDD1.n6 B 0.012928f
C556 VDD1.n7 B 0.030556f
C557 VDD1.n8 B 0.013688f
C558 VDD1.n9 B 0.024058f
C559 VDD1.n10 B 0.012928f
C560 VDD1.n11 B 0.030556f
C561 VDD1.n12 B 0.013688f
C562 VDD1.n13 B 0.024058f
C563 VDD1.n14 B 0.012928f
C564 VDD1.n15 B 0.030556f
C565 VDD1.n16 B 0.013688f
C566 VDD1.n17 B 0.024058f
C567 VDD1.n18 B 0.012928f
C568 VDD1.n19 B 0.030556f
C569 VDD1.n20 B 0.030556f
C570 VDD1.n21 B 0.013688f
C571 VDD1.n22 B 0.024058f
C572 VDD1.n23 B 0.012928f
C573 VDD1.n24 B 0.030556f
C574 VDD1.n25 B 0.013688f
C575 VDD1.n26 B 0.200054f
C576 VDD1.t5 B 0.05198f
C577 VDD1.n27 B 0.022917f
C578 VDD1.n28 B 0.021601f
C579 VDD1.n29 B 0.012928f
C580 VDD1.n30 B 1.52185f
C581 VDD1.n31 B 0.024058f
C582 VDD1.n32 B 0.012928f
C583 VDD1.n33 B 0.013688f
C584 VDD1.n34 B 0.030556f
C585 VDD1.n35 B 0.030556f
C586 VDD1.n36 B 0.013688f
C587 VDD1.n37 B 0.012928f
C588 VDD1.n38 B 0.024058f
C589 VDD1.n39 B 0.024058f
C590 VDD1.n40 B 0.012928f
C591 VDD1.n41 B 0.013688f
C592 VDD1.n42 B 0.030556f
C593 VDD1.n43 B 0.030556f
C594 VDD1.n44 B 0.013688f
C595 VDD1.n45 B 0.012928f
C596 VDD1.n46 B 0.024058f
C597 VDD1.n47 B 0.024058f
C598 VDD1.n48 B 0.012928f
C599 VDD1.n49 B 0.013308f
C600 VDD1.n50 B 0.013308f
C601 VDD1.n51 B 0.030556f
C602 VDD1.n52 B 0.030556f
C603 VDD1.n53 B 0.013688f
C604 VDD1.n54 B 0.012928f
C605 VDD1.n55 B 0.024058f
C606 VDD1.n56 B 0.024058f
C607 VDD1.n57 B 0.012928f
C608 VDD1.n58 B 0.013688f
C609 VDD1.n59 B 0.030556f
C610 VDD1.n60 B 0.030556f
C611 VDD1.n61 B 0.013688f
C612 VDD1.n62 B 0.012928f
C613 VDD1.n63 B 0.024058f
C614 VDD1.n64 B 0.024058f
C615 VDD1.n65 B 0.012928f
C616 VDD1.n66 B 0.013688f
C617 VDD1.n67 B 0.030556f
C618 VDD1.n68 B 0.030556f
C619 VDD1.n69 B 0.013688f
C620 VDD1.n70 B 0.012928f
C621 VDD1.n71 B 0.024058f
C622 VDD1.n72 B 0.024058f
C623 VDD1.n73 B 0.012928f
C624 VDD1.n74 B 0.013688f
C625 VDD1.n75 B 0.030556f
C626 VDD1.n76 B 0.067297f
C627 VDD1.n77 B 0.013688f
C628 VDD1.n78 B 0.012928f
C629 VDD1.n79 B 0.051665f
C630 VDD1.n80 B 0.055584f
C631 VDD1.n81 B 0.034465f
C632 VDD1.n82 B 0.024058f
C633 VDD1.n83 B 0.012928f
C634 VDD1.n84 B 0.030556f
C635 VDD1.n85 B 0.013688f
C636 VDD1.n86 B 0.024058f
C637 VDD1.n87 B 0.012928f
C638 VDD1.n88 B 0.030556f
C639 VDD1.n89 B 0.013688f
C640 VDD1.n90 B 0.024058f
C641 VDD1.n91 B 0.012928f
C642 VDD1.n92 B 0.030556f
C643 VDD1.n93 B 0.013688f
C644 VDD1.n94 B 0.024058f
C645 VDD1.n95 B 0.012928f
C646 VDD1.n96 B 0.030556f
C647 VDD1.n97 B 0.013688f
C648 VDD1.n98 B 0.024058f
C649 VDD1.n99 B 0.012928f
C650 VDD1.n100 B 0.030556f
C651 VDD1.n101 B 0.013688f
C652 VDD1.n102 B 0.024058f
C653 VDD1.n103 B 0.012928f
C654 VDD1.n104 B 0.030556f
C655 VDD1.n105 B 0.013688f
C656 VDD1.n106 B 0.200054f
C657 VDD1.t4 B 0.05198f
C658 VDD1.n107 B 0.022917f
C659 VDD1.n108 B 0.021601f
C660 VDD1.n109 B 0.012928f
C661 VDD1.n110 B 1.52185f
C662 VDD1.n111 B 0.024058f
C663 VDD1.n112 B 0.012928f
C664 VDD1.n113 B 0.013688f
C665 VDD1.n114 B 0.030556f
C666 VDD1.n115 B 0.030556f
C667 VDD1.n116 B 0.013688f
C668 VDD1.n117 B 0.012928f
C669 VDD1.n118 B 0.024058f
C670 VDD1.n119 B 0.024058f
C671 VDD1.n120 B 0.012928f
C672 VDD1.n121 B 0.013688f
C673 VDD1.n122 B 0.030556f
C674 VDD1.n123 B 0.030556f
C675 VDD1.n124 B 0.030556f
C676 VDD1.n125 B 0.013688f
C677 VDD1.n126 B 0.012928f
C678 VDD1.n127 B 0.024058f
C679 VDD1.n128 B 0.024058f
C680 VDD1.n129 B 0.012928f
C681 VDD1.n130 B 0.013308f
C682 VDD1.n131 B 0.013308f
C683 VDD1.n132 B 0.030556f
C684 VDD1.n133 B 0.030556f
C685 VDD1.n134 B 0.013688f
C686 VDD1.n135 B 0.012928f
C687 VDD1.n136 B 0.024058f
C688 VDD1.n137 B 0.024058f
C689 VDD1.n138 B 0.012928f
C690 VDD1.n139 B 0.013688f
C691 VDD1.n140 B 0.030556f
C692 VDD1.n141 B 0.030556f
C693 VDD1.n142 B 0.013688f
C694 VDD1.n143 B 0.012928f
C695 VDD1.n144 B 0.024058f
C696 VDD1.n145 B 0.024058f
C697 VDD1.n146 B 0.012928f
C698 VDD1.n147 B 0.013688f
C699 VDD1.n148 B 0.030556f
C700 VDD1.n149 B 0.030556f
C701 VDD1.n150 B 0.013688f
C702 VDD1.n151 B 0.012928f
C703 VDD1.n152 B 0.024058f
C704 VDD1.n153 B 0.024058f
C705 VDD1.n154 B 0.012928f
C706 VDD1.n155 B 0.013688f
C707 VDD1.n156 B 0.030556f
C708 VDD1.n157 B 0.067297f
C709 VDD1.n158 B 0.013688f
C710 VDD1.n159 B 0.012928f
C711 VDD1.n160 B 0.051665f
C712 VDD1.n161 B 0.055273f
C713 VDD1.t3 B 0.282887f
C714 VDD1.t1 B 0.282887f
C715 VDD1.n162 B 2.54793f
C716 VDD1.n163 B 1.97935f
C717 VDD1.t0 B 0.282887f
C718 VDD1.t2 B 0.282887f
C719 VDD1.n164 B 2.54725f
C720 VDD1.n165 B 2.35782f
C721 VP.n0 B 0.066138f
C722 VP.t1 B 1.2364f
C723 VP.n1 B 0.456685f
C724 VP.t4 B 1.21858f
C725 VP.t2 B 1.21858f
C726 VP.n2 B 0.484729f
C727 VP.n3 B 0.473455f
C728 VP.n4 B 2.29075f
C729 VP.n5 B 2.18878f
C730 VP.t5 B 1.21858f
C731 VP.n6 B 0.473455f
C732 VP.t0 B 1.21858f
C733 VP.n7 B 0.484729f
C734 VP.t3 B 1.21858f
C735 VP.n8 B 0.473455f
C736 VP.n9 B 0.055113f
.ends

