* NGSPICE file created from diff_pair_sample_0397.ext - technology: sky130A

.subckt diff_pair_sample_0397 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=5.2221 pd=27.56 as=5.2221 ps=27.56 w=13.39 l=3.05
X1 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.2221 pd=27.56 as=5.2221 ps=27.56 w=13.39 l=3.05
X2 VDD2.t0 VN.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=5.2221 pd=27.56 as=5.2221 ps=27.56 w=13.39 l=3.05
X3 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=5.2221 pd=27.56 as=0 ps=0 w=13.39 l=3.05
X4 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=5.2221 pd=27.56 as=0 ps=0 w=13.39 l=3.05
X5 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.2221 pd=27.56 as=5.2221 ps=27.56 w=13.39 l=3.05
X6 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=5.2221 pd=27.56 as=0 ps=0 w=13.39 l=3.05
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=5.2221 pd=27.56 as=0 ps=0 w=13.39 l=3.05
R0 VN VN.t1 193.804
R1 VN VN.t0 147.331
R2 VTAIL.n282 VTAIL.n216 214.453
R3 VTAIL.n66 VTAIL.n0 214.453
R4 VTAIL.n210 VTAIL.n144 214.453
R5 VTAIL.n138 VTAIL.n72 214.453
R6 VTAIL.n241 VTAIL.n240 185
R7 VTAIL.n243 VTAIL.n242 185
R8 VTAIL.n236 VTAIL.n235 185
R9 VTAIL.n249 VTAIL.n248 185
R10 VTAIL.n251 VTAIL.n250 185
R11 VTAIL.n232 VTAIL.n231 185
R12 VTAIL.n257 VTAIL.n256 185
R13 VTAIL.n259 VTAIL.n258 185
R14 VTAIL.n228 VTAIL.n227 185
R15 VTAIL.n265 VTAIL.n264 185
R16 VTAIL.n267 VTAIL.n266 185
R17 VTAIL.n224 VTAIL.n223 185
R18 VTAIL.n273 VTAIL.n272 185
R19 VTAIL.n275 VTAIL.n274 185
R20 VTAIL.n220 VTAIL.n219 185
R21 VTAIL.n281 VTAIL.n280 185
R22 VTAIL.n283 VTAIL.n282 185
R23 VTAIL.n25 VTAIL.n24 185
R24 VTAIL.n27 VTAIL.n26 185
R25 VTAIL.n20 VTAIL.n19 185
R26 VTAIL.n33 VTAIL.n32 185
R27 VTAIL.n35 VTAIL.n34 185
R28 VTAIL.n16 VTAIL.n15 185
R29 VTAIL.n41 VTAIL.n40 185
R30 VTAIL.n43 VTAIL.n42 185
R31 VTAIL.n12 VTAIL.n11 185
R32 VTAIL.n49 VTAIL.n48 185
R33 VTAIL.n51 VTAIL.n50 185
R34 VTAIL.n8 VTAIL.n7 185
R35 VTAIL.n57 VTAIL.n56 185
R36 VTAIL.n59 VTAIL.n58 185
R37 VTAIL.n4 VTAIL.n3 185
R38 VTAIL.n65 VTAIL.n64 185
R39 VTAIL.n67 VTAIL.n66 185
R40 VTAIL.n211 VTAIL.n210 185
R41 VTAIL.n209 VTAIL.n208 185
R42 VTAIL.n148 VTAIL.n147 185
R43 VTAIL.n203 VTAIL.n202 185
R44 VTAIL.n201 VTAIL.n200 185
R45 VTAIL.n152 VTAIL.n151 185
R46 VTAIL.n195 VTAIL.n194 185
R47 VTAIL.n193 VTAIL.n192 185
R48 VTAIL.n156 VTAIL.n155 185
R49 VTAIL.n187 VTAIL.n186 185
R50 VTAIL.n185 VTAIL.n184 185
R51 VTAIL.n160 VTAIL.n159 185
R52 VTAIL.n179 VTAIL.n178 185
R53 VTAIL.n177 VTAIL.n176 185
R54 VTAIL.n164 VTAIL.n163 185
R55 VTAIL.n171 VTAIL.n170 185
R56 VTAIL.n169 VTAIL.n168 185
R57 VTAIL.n139 VTAIL.n138 185
R58 VTAIL.n137 VTAIL.n136 185
R59 VTAIL.n76 VTAIL.n75 185
R60 VTAIL.n131 VTAIL.n130 185
R61 VTAIL.n129 VTAIL.n128 185
R62 VTAIL.n80 VTAIL.n79 185
R63 VTAIL.n123 VTAIL.n122 185
R64 VTAIL.n121 VTAIL.n120 185
R65 VTAIL.n84 VTAIL.n83 185
R66 VTAIL.n115 VTAIL.n114 185
R67 VTAIL.n113 VTAIL.n112 185
R68 VTAIL.n88 VTAIL.n87 185
R69 VTAIL.n107 VTAIL.n106 185
R70 VTAIL.n105 VTAIL.n104 185
R71 VTAIL.n92 VTAIL.n91 185
R72 VTAIL.n99 VTAIL.n98 185
R73 VTAIL.n97 VTAIL.n96 185
R74 VTAIL.n239 VTAIL.t3 147.659
R75 VTAIL.n23 VTAIL.t1 147.659
R76 VTAIL.n167 VTAIL.t0 147.659
R77 VTAIL.n95 VTAIL.t2 147.659
R78 VTAIL.n242 VTAIL.n241 104.615
R79 VTAIL.n242 VTAIL.n235 104.615
R80 VTAIL.n249 VTAIL.n235 104.615
R81 VTAIL.n250 VTAIL.n249 104.615
R82 VTAIL.n250 VTAIL.n231 104.615
R83 VTAIL.n257 VTAIL.n231 104.615
R84 VTAIL.n258 VTAIL.n257 104.615
R85 VTAIL.n258 VTAIL.n227 104.615
R86 VTAIL.n265 VTAIL.n227 104.615
R87 VTAIL.n266 VTAIL.n265 104.615
R88 VTAIL.n266 VTAIL.n223 104.615
R89 VTAIL.n273 VTAIL.n223 104.615
R90 VTAIL.n274 VTAIL.n273 104.615
R91 VTAIL.n274 VTAIL.n219 104.615
R92 VTAIL.n281 VTAIL.n219 104.615
R93 VTAIL.n282 VTAIL.n281 104.615
R94 VTAIL.n26 VTAIL.n25 104.615
R95 VTAIL.n26 VTAIL.n19 104.615
R96 VTAIL.n33 VTAIL.n19 104.615
R97 VTAIL.n34 VTAIL.n33 104.615
R98 VTAIL.n34 VTAIL.n15 104.615
R99 VTAIL.n41 VTAIL.n15 104.615
R100 VTAIL.n42 VTAIL.n41 104.615
R101 VTAIL.n42 VTAIL.n11 104.615
R102 VTAIL.n49 VTAIL.n11 104.615
R103 VTAIL.n50 VTAIL.n49 104.615
R104 VTAIL.n50 VTAIL.n7 104.615
R105 VTAIL.n57 VTAIL.n7 104.615
R106 VTAIL.n58 VTAIL.n57 104.615
R107 VTAIL.n58 VTAIL.n3 104.615
R108 VTAIL.n65 VTAIL.n3 104.615
R109 VTAIL.n66 VTAIL.n65 104.615
R110 VTAIL.n210 VTAIL.n209 104.615
R111 VTAIL.n209 VTAIL.n147 104.615
R112 VTAIL.n202 VTAIL.n147 104.615
R113 VTAIL.n202 VTAIL.n201 104.615
R114 VTAIL.n201 VTAIL.n151 104.615
R115 VTAIL.n194 VTAIL.n151 104.615
R116 VTAIL.n194 VTAIL.n193 104.615
R117 VTAIL.n193 VTAIL.n155 104.615
R118 VTAIL.n186 VTAIL.n155 104.615
R119 VTAIL.n186 VTAIL.n185 104.615
R120 VTAIL.n185 VTAIL.n159 104.615
R121 VTAIL.n178 VTAIL.n159 104.615
R122 VTAIL.n178 VTAIL.n177 104.615
R123 VTAIL.n177 VTAIL.n163 104.615
R124 VTAIL.n170 VTAIL.n163 104.615
R125 VTAIL.n170 VTAIL.n169 104.615
R126 VTAIL.n138 VTAIL.n137 104.615
R127 VTAIL.n137 VTAIL.n75 104.615
R128 VTAIL.n130 VTAIL.n75 104.615
R129 VTAIL.n130 VTAIL.n129 104.615
R130 VTAIL.n129 VTAIL.n79 104.615
R131 VTAIL.n122 VTAIL.n79 104.615
R132 VTAIL.n122 VTAIL.n121 104.615
R133 VTAIL.n121 VTAIL.n83 104.615
R134 VTAIL.n114 VTAIL.n83 104.615
R135 VTAIL.n114 VTAIL.n113 104.615
R136 VTAIL.n113 VTAIL.n87 104.615
R137 VTAIL.n106 VTAIL.n87 104.615
R138 VTAIL.n106 VTAIL.n105 104.615
R139 VTAIL.n105 VTAIL.n91 104.615
R140 VTAIL.n98 VTAIL.n91 104.615
R141 VTAIL.n98 VTAIL.n97 104.615
R142 VTAIL.n241 VTAIL.t3 52.3082
R143 VTAIL.n25 VTAIL.t1 52.3082
R144 VTAIL.n169 VTAIL.t0 52.3082
R145 VTAIL.n97 VTAIL.t2 52.3082
R146 VTAIL.n287 VTAIL.n286 35.8702
R147 VTAIL.n71 VTAIL.n70 35.8702
R148 VTAIL.n215 VTAIL.n214 35.8702
R149 VTAIL.n143 VTAIL.n142 35.8702
R150 VTAIL.n143 VTAIL.n71 29.7376
R151 VTAIL.n287 VTAIL.n215 26.8238
R152 VTAIL.n240 VTAIL.n239 15.6677
R153 VTAIL.n24 VTAIL.n23 15.6677
R154 VTAIL.n168 VTAIL.n167 15.6677
R155 VTAIL.n96 VTAIL.n95 15.6677
R156 VTAIL.n243 VTAIL.n238 12.8005
R157 VTAIL.n284 VTAIL.n283 12.8005
R158 VTAIL.n27 VTAIL.n22 12.8005
R159 VTAIL.n68 VTAIL.n67 12.8005
R160 VTAIL.n212 VTAIL.n211 12.8005
R161 VTAIL.n171 VTAIL.n166 12.8005
R162 VTAIL.n140 VTAIL.n139 12.8005
R163 VTAIL.n99 VTAIL.n94 12.8005
R164 VTAIL.n244 VTAIL.n236 12.0247
R165 VTAIL.n280 VTAIL.n218 12.0247
R166 VTAIL.n28 VTAIL.n20 12.0247
R167 VTAIL.n64 VTAIL.n2 12.0247
R168 VTAIL.n208 VTAIL.n146 12.0247
R169 VTAIL.n172 VTAIL.n164 12.0247
R170 VTAIL.n136 VTAIL.n74 12.0247
R171 VTAIL.n100 VTAIL.n92 12.0247
R172 VTAIL.n248 VTAIL.n247 11.249
R173 VTAIL.n279 VTAIL.n220 11.249
R174 VTAIL.n32 VTAIL.n31 11.249
R175 VTAIL.n63 VTAIL.n4 11.249
R176 VTAIL.n207 VTAIL.n148 11.249
R177 VTAIL.n176 VTAIL.n175 11.249
R178 VTAIL.n135 VTAIL.n76 11.249
R179 VTAIL.n104 VTAIL.n103 11.249
R180 VTAIL.n251 VTAIL.n234 10.4732
R181 VTAIL.n276 VTAIL.n275 10.4732
R182 VTAIL.n35 VTAIL.n18 10.4732
R183 VTAIL.n60 VTAIL.n59 10.4732
R184 VTAIL.n204 VTAIL.n203 10.4732
R185 VTAIL.n179 VTAIL.n162 10.4732
R186 VTAIL.n132 VTAIL.n131 10.4732
R187 VTAIL.n107 VTAIL.n90 10.4732
R188 VTAIL.n252 VTAIL.n232 9.69747
R189 VTAIL.n272 VTAIL.n222 9.69747
R190 VTAIL.n36 VTAIL.n16 9.69747
R191 VTAIL.n56 VTAIL.n6 9.69747
R192 VTAIL.n200 VTAIL.n150 9.69747
R193 VTAIL.n180 VTAIL.n160 9.69747
R194 VTAIL.n128 VTAIL.n78 9.69747
R195 VTAIL.n108 VTAIL.n88 9.69747
R196 VTAIL.n286 VTAIL.n285 9.45567
R197 VTAIL.n70 VTAIL.n69 9.45567
R198 VTAIL.n214 VTAIL.n213 9.45567
R199 VTAIL.n142 VTAIL.n141 9.45567
R200 VTAIL.n261 VTAIL.n260 9.3005
R201 VTAIL.n230 VTAIL.n229 9.3005
R202 VTAIL.n255 VTAIL.n254 9.3005
R203 VTAIL.n253 VTAIL.n252 9.3005
R204 VTAIL.n234 VTAIL.n233 9.3005
R205 VTAIL.n247 VTAIL.n246 9.3005
R206 VTAIL.n245 VTAIL.n244 9.3005
R207 VTAIL.n238 VTAIL.n237 9.3005
R208 VTAIL.n263 VTAIL.n262 9.3005
R209 VTAIL.n226 VTAIL.n225 9.3005
R210 VTAIL.n269 VTAIL.n268 9.3005
R211 VTAIL.n271 VTAIL.n270 9.3005
R212 VTAIL.n222 VTAIL.n221 9.3005
R213 VTAIL.n277 VTAIL.n276 9.3005
R214 VTAIL.n279 VTAIL.n278 9.3005
R215 VTAIL.n218 VTAIL.n217 9.3005
R216 VTAIL.n285 VTAIL.n284 9.3005
R217 VTAIL.n45 VTAIL.n44 9.3005
R218 VTAIL.n14 VTAIL.n13 9.3005
R219 VTAIL.n39 VTAIL.n38 9.3005
R220 VTAIL.n37 VTAIL.n36 9.3005
R221 VTAIL.n18 VTAIL.n17 9.3005
R222 VTAIL.n31 VTAIL.n30 9.3005
R223 VTAIL.n29 VTAIL.n28 9.3005
R224 VTAIL.n22 VTAIL.n21 9.3005
R225 VTAIL.n47 VTAIL.n46 9.3005
R226 VTAIL.n10 VTAIL.n9 9.3005
R227 VTAIL.n53 VTAIL.n52 9.3005
R228 VTAIL.n55 VTAIL.n54 9.3005
R229 VTAIL.n6 VTAIL.n5 9.3005
R230 VTAIL.n61 VTAIL.n60 9.3005
R231 VTAIL.n63 VTAIL.n62 9.3005
R232 VTAIL.n2 VTAIL.n1 9.3005
R233 VTAIL.n69 VTAIL.n68 9.3005
R234 VTAIL.n154 VTAIL.n153 9.3005
R235 VTAIL.n197 VTAIL.n196 9.3005
R236 VTAIL.n199 VTAIL.n198 9.3005
R237 VTAIL.n150 VTAIL.n149 9.3005
R238 VTAIL.n205 VTAIL.n204 9.3005
R239 VTAIL.n207 VTAIL.n206 9.3005
R240 VTAIL.n146 VTAIL.n145 9.3005
R241 VTAIL.n213 VTAIL.n212 9.3005
R242 VTAIL.n191 VTAIL.n190 9.3005
R243 VTAIL.n189 VTAIL.n188 9.3005
R244 VTAIL.n158 VTAIL.n157 9.3005
R245 VTAIL.n183 VTAIL.n182 9.3005
R246 VTAIL.n181 VTAIL.n180 9.3005
R247 VTAIL.n162 VTAIL.n161 9.3005
R248 VTAIL.n175 VTAIL.n174 9.3005
R249 VTAIL.n173 VTAIL.n172 9.3005
R250 VTAIL.n166 VTAIL.n165 9.3005
R251 VTAIL.n82 VTAIL.n81 9.3005
R252 VTAIL.n125 VTAIL.n124 9.3005
R253 VTAIL.n127 VTAIL.n126 9.3005
R254 VTAIL.n78 VTAIL.n77 9.3005
R255 VTAIL.n133 VTAIL.n132 9.3005
R256 VTAIL.n135 VTAIL.n134 9.3005
R257 VTAIL.n74 VTAIL.n73 9.3005
R258 VTAIL.n141 VTAIL.n140 9.3005
R259 VTAIL.n119 VTAIL.n118 9.3005
R260 VTAIL.n117 VTAIL.n116 9.3005
R261 VTAIL.n86 VTAIL.n85 9.3005
R262 VTAIL.n111 VTAIL.n110 9.3005
R263 VTAIL.n109 VTAIL.n108 9.3005
R264 VTAIL.n90 VTAIL.n89 9.3005
R265 VTAIL.n103 VTAIL.n102 9.3005
R266 VTAIL.n101 VTAIL.n100 9.3005
R267 VTAIL.n94 VTAIL.n93 9.3005
R268 VTAIL.n256 VTAIL.n255 8.92171
R269 VTAIL.n271 VTAIL.n224 8.92171
R270 VTAIL.n40 VTAIL.n39 8.92171
R271 VTAIL.n55 VTAIL.n8 8.92171
R272 VTAIL.n199 VTAIL.n152 8.92171
R273 VTAIL.n184 VTAIL.n183 8.92171
R274 VTAIL.n127 VTAIL.n80 8.92171
R275 VTAIL.n112 VTAIL.n111 8.92171
R276 VTAIL.n286 VTAIL.n216 8.2187
R277 VTAIL.n70 VTAIL.n0 8.2187
R278 VTAIL.n214 VTAIL.n144 8.2187
R279 VTAIL.n142 VTAIL.n72 8.2187
R280 VTAIL.n259 VTAIL.n230 8.14595
R281 VTAIL.n268 VTAIL.n267 8.14595
R282 VTAIL.n43 VTAIL.n14 8.14595
R283 VTAIL.n52 VTAIL.n51 8.14595
R284 VTAIL.n196 VTAIL.n195 8.14595
R285 VTAIL.n187 VTAIL.n158 8.14595
R286 VTAIL.n124 VTAIL.n123 8.14595
R287 VTAIL.n115 VTAIL.n86 8.14595
R288 VTAIL.n260 VTAIL.n228 7.3702
R289 VTAIL.n264 VTAIL.n226 7.3702
R290 VTAIL.n44 VTAIL.n12 7.3702
R291 VTAIL.n48 VTAIL.n10 7.3702
R292 VTAIL.n192 VTAIL.n154 7.3702
R293 VTAIL.n188 VTAIL.n156 7.3702
R294 VTAIL.n120 VTAIL.n82 7.3702
R295 VTAIL.n116 VTAIL.n84 7.3702
R296 VTAIL.n263 VTAIL.n228 6.59444
R297 VTAIL.n264 VTAIL.n263 6.59444
R298 VTAIL.n47 VTAIL.n12 6.59444
R299 VTAIL.n48 VTAIL.n47 6.59444
R300 VTAIL.n192 VTAIL.n191 6.59444
R301 VTAIL.n191 VTAIL.n156 6.59444
R302 VTAIL.n120 VTAIL.n119 6.59444
R303 VTAIL.n119 VTAIL.n84 6.59444
R304 VTAIL.n260 VTAIL.n259 5.81868
R305 VTAIL.n267 VTAIL.n226 5.81868
R306 VTAIL.n44 VTAIL.n43 5.81868
R307 VTAIL.n51 VTAIL.n10 5.81868
R308 VTAIL.n195 VTAIL.n154 5.81868
R309 VTAIL.n188 VTAIL.n187 5.81868
R310 VTAIL.n123 VTAIL.n82 5.81868
R311 VTAIL.n116 VTAIL.n115 5.81868
R312 VTAIL.n284 VTAIL.n216 5.3904
R313 VTAIL.n68 VTAIL.n0 5.3904
R314 VTAIL.n212 VTAIL.n144 5.3904
R315 VTAIL.n140 VTAIL.n72 5.3904
R316 VTAIL.n256 VTAIL.n230 5.04292
R317 VTAIL.n268 VTAIL.n224 5.04292
R318 VTAIL.n40 VTAIL.n14 5.04292
R319 VTAIL.n52 VTAIL.n8 5.04292
R320 VTAIL.n196 VTAIL.n152 5.04292
R321 VTAIL.n184 VTAIL.n158 5.04292
R322 VTAIL.n124 VTAIL.n80 5.04292
R323 VTAIL.n112 VTAIL.n86 5.04292
R324 VTAIL.n239 VTAIL.n237 4.38563
R325 VTAIL.n23 VTAIL.n21 4.38563
R326 VTAIL.n167 VTAIL.n165 4.38563
R327 VTAIL.n95 VTAIL.n93 4.38563
R328 VTAIL.n255 VTAIL.n232 4.26717
R329 VTAIL.n272 VTAIL.n271 4.26717
R330 VTAIL.n39 VTAIL.n16 4.26717
R331 VTAIL.n56 VTAIL.n55 4.26717
R332 VTAIL.n200 VTAIL.n199 4.26717
R333 VTAIL.n183 VTAIL.n160 4.26717
R334 VTAIL.n128 VTAIL.n127 4.26717
R335 VTAIL.n111 VTAIL.n88 4.26717
R336 VTAIL.n252 VTAIL.n251 3.49141
R337 VTAIL.n275 VTAIL.n222 3.49141
R338 VTAIL.n36 VTAIL.n35 3.49141
R339 VTAIL.n59 VTAIL.n6 3.49141
R340 VTAIL.n203 VTAIL.n150 3.49141
R341 VTAIL.n180 VTAIL.n179 3.49141
R342 VTAIL.n131 VTAIL.n78 3.49141
R343 VTAIL.n108 VTAIL.n107 3.49141
R344 VTAIL.n248 VTAIL.n234 2.71565
R345 VTAIL.n276 VTAIL.n220 2.71565
R346 VTAIL.n32 VTAIL.n18 2.71565
R347 VTAIL.n60 VTAIL.n4 2.71565
R348 VTAIL.n204 VTAIL.n148 2.71565
R349 VTAIL.n176 VTAIL.n162 2.71565
R350 VTAIL.n132 VTAIL.n76 2.71565
R351 VTAIL.n104 VTAIL.n90 2.71565
R352 VTAIL.n247 VTAIL.n236 1.93989
R353 VTAIL.n280 VTAIL.n279 1.93989
R354 VTAIL.n31 VTAIL.n20 1.93989
R355 VTAIL.n64 VTAIL.n63 1.93989
R356 VTAIL.n208 VTAIL.n207 1.93989
R357 VTAIL.n175 VTAIL.n164 1.93989
R358 VTAIL.n136 VTAIL.n135 1.93989
R359 VTAIL.n103 VTAIL.n92 1.93989
R360 VTAIL.n215 VTAIL.n143 1.92722
R361 VTAIL VTAIL.n71 1.25697
R362 VTAIL.n244 VTAIL.n243 1.16414
R363 VTAIL.n283 VTAIL.n218 1.16414
R364 VTAIL.n28 VTAIL.n27 1.16414
R365 VTAIL.n67 VTAIL.n2 1.16414
R366 VTAIL.n211 VTAIL.n146 1.16414
R367 VTAIL.n172 VTAIL.n171 1.16414
R368 VTAIL.n139 VTAIL.n74 1.16414
R369 VTAIL.n100 VTAIL.n99 1.16414
R370 VTAIL VTAIL.n287 0.670759
R371 VTAIL.n240 VTAIL.n238 0.388379
R372 VTAIL.n24 VTAIL.n22 0.388379
R373 VTAIL.n168 VTAIL.n166 0.388379
R374 VTAIL.n96 VTAIL.n94 0.388379
R375 VTAIL.n245 VTAIL.n237 0.155672
R376 VTAIL.n246 VTAIL.n245 0.155672
R377 VTAIL.n246 VTAIL.n233 0.155672
R378 VTAIL.n253 VTAIL.n233 0.155672
R379 VTAIL.n254 VTAIL.n253 0.155672
R380 VTAIL.n254 VTAIL.n229 0.155672
R381 VTAIL.n261 VTAIL.n229 0.155672
R382 VTAIL.n262 VTAIL.n261 0.155672
R383 VTAIL.n262 VTAIL.n225 0.155672
R384 VTAIL.n269 VTAIL.n225 0.155672
R385 VTAIL.n270 VTAIL.n269 0.155672
R386 VTAIL.n270 VTAIL.n221 0.155672
R387 VTAIL.n277 VTAIL.n221 0.155672
R388 VTAIL.n278 VTAIL.n277 0.155672
R389 VTAIL.n278 VTAIL.n217 0.155672
R390 VTAIL.n285 VTAIL.n217 0.155672
R391 VTAIL.n29 VTAIL.n21 0.155672
R392 VTAIL.n30 VTAIL.n29 0.155672
R393 VTAIL.n30 VTAIL.n17 0.155672
R394 VTAIL.n37 VTAIL.n17 0.155672
R395 VTAIL.n38 VTAIL.n37 0.155672
R396 VTAIL.n38 VTAIL.n13 0.155672
R397 VTAIL.n45 VTAIL.n13 0.155672
R398 VTAIL.n46 VTAIL.n45 0.155672
R399 VTAIL.n46 VTAIL.n9 0.155672
R400 VTAIL.n53 VTAIL.n9 0.155672
R401 VTAIL.n54 VTAIL.n53 0.155672
R402 VTAIL.n54 VTAIL.n5 0.155672
R403 VTAIL.n61 VTAIL.n5 0.155672
R404 VTAIL.n62 VTAIL.n61 0.155672
R405 VTAIL.n62 VTAIL.n1 0.155672
R406 VTAIL.n69 VTAIL.n1 0.155672
R407 VTAIL.n213 VTAIL.n145 0.155672
R408 VTAIL.n206 VTAIL.n145 0.155672
R409 VTAIL.n206 VTAIL.n205 0.155672
R410 VTAIL.n205 VTAIL.n149 0.155672
R411 VTAIL.n198 VTAIL.n149 0.155672
R412 VTAIL.n198 VTAIL.n197 0.155672
R413 VTAIL.n197 VTAIL.n153 0.155672
R414 VTAIL.n190 VTAIL.n153 0.155672
R415 VTAIL.n190 VTAIL.n189 0.155672
R416 VTAIL.n189 VTAIL.n157 0.155672
R417 VTAIL.n182 VTAIL.n157 0.155672
R418 VTAIL.n182 VTAIL.n181 0.155672
R419 VTAIL.n181 VTAIL.n161 0.155672
R420 VTAIL.n174 VTAIL.n161 0.155672
R421 VTAIL.n174 VTAIL.n173 0.155672
R422 VTAIL.n173 VTAIL.n165 0.155672
R423 VTAIL.n141 VTAIL.n73 0.155672
R424 VTAIL.n134 VTAIL.n73 0.155672
R425 VTAIL.n134 VTAIL.n133 0.155672
R426 VTAIL.n133 VTAIL.n77 0.155672
R427 VTAIL.n126 VTAIL.n77 0.155672
R428 VTAIL.n126 VTAIL.n125 0.155672
R429 VTAIL.n125 VTAIL.n81 0.155672
R430 VTAIL.n118 VTAIL.n81 0.155672
R431 VTAIL.n118 VTAIL.n117 0.155672
R432 VTAIL.n117 VTAIL.n85 0.155672
R433 VTAIL.n110 VTAIL.n85 0.155672
R434 VTAIL.n110 VTAIL.n109 0.155672
R435 VTAIL.n109 VTAIL.n89 0.155672
R436 VTAIL.n102 VTAIL.n89 0.155672
R437 VTAIL.n102 VTAIL.n101 0.155672
R438 VTAIL.n101 VTAIL.n93 0.155672
R439 VDD2.n137 VDD2.n71 214.453
R440 VDD2.n66 VDD2.n0 214.453
R441 VDD2.n138 VDD2.n137 185
R442 VDD2.n136 VDD2.n135 185
R443 VDD2.n75 VDD2.n74 185
R444 VDD2.n130 VDD2.n129 185
R445 VDD2.n128 VDD2.n127 185
R446 VDD2.n79 VDD2.n78 185
R447 VDD2.n122 VDD2.n121 185
R448 VDD2.n120 VDD2.n119 185
R449 VDD2.n83 VDD2.n82 185
R450 VDD2.n114 VDD2.n113 185
R451 VDD2.n112 VDD2.n111 185
R452 VDD2.n87 VDD2.n86 185
R453 VDD2.n106 VDD2.n105 185
R454 VDD2.n104 VDD2.n103 185
R455 VDD2.n91 VDD2.n90 185
R456 VDD2.n98 VDD2.n97 185
R457 VDD2.n96 VDD2.n95 185
R458 VDD2.n25 VDD2.n24 185
R459 VDD2.n27 VDD2.n26 185
R460 VDD2.n20 VDD2.n19 185
R461 VDD2.n33 VDD2.n32 185
R462 VDD2.n35 VDD2.n34 185
R463 VDD2.n16 VDD2.n15 185
R464 VDD2.n41 VDD2.n40 185
R465 VDD2.n43 VDD2.n42 185
R466 VDD2.n12 VDD2.n11 185
R467 VDD2.n49 VDD2.n48 185
R468 VDD2.n51 VDD2.n50 185
R469 VDD2.n8 VDD2.n7 185
R470 VDD2.n57 VDD2.n56 185
R471 VDD2.n59 VDD2.n58 185
R472 VDD2.n4 VDD2.n3 185
R473 VDD2.n65 VDD2.n64 185
R474 VDD2.n67 VDD2.n66 185
R475 VDD2.n23 VDD2.t1 147.659
R476 VDD2.n94 VDD2.t0 147.659
R477 VDD2.n137 VDD2.n136 104.615
R478 VDD2.n136 VDD2.n74 104.615
R479 VDD2.n129 VDD2.n74 104.615
R480 VDD2.n129 VDD2.n128 104.615
R481 VDD2.n128 VDD2.n78 104.615
R482 VDD2.n121 VDD2.n78 104.615
R483 VDD2.n121 VDD2.n120 104.615
R484 VDD2.n120 VDD2.n82 104.615
R485 VDD2.n113 VDD2.n82 104.615
R486 VDD2.n113 VDD2.n112 104.615
R487 VDD2.n112 VDD2.n86 104.615
R488 VDD2.n105 VDD2.n86 104.615
R489 VDD2.n105 VDD2.n104 104.615
R490 VDD2.n104 VDD2.n90 104.615
R491 VDD2.n97 VDD2.n90 104.615
R492 VDD2.n97 VDD2.n96 104.615
R493 VDD2.n26 VDD2.n25 104.615
R494 VDD2.n26 VDD2.n19 104.615
R495 VDD2.n33 VDD2.n19 104.615
R496 VDD2.n34 VDD2.n33 104.615
R497 VDD2.n34 VDD2.n15 104.615
R498 VDD2.n41 VDD2.n15 104.615
R499 VDD2.n42 VDD2.n41 104.615
R500 VDD2.n42 VDD2.n11 104.615
R501 VDD2.n49 VDD2.n11 104.615
R502 VDD2.n50 VDD2.n49 104.615
R503 VDD2.n50 VDD2.n7 104.615
R504 VDD2.n57 VDD2.n7 104.615
R505 VDD2.n58 VDD2.n57 104.615
R506 VDD2.n58 VDD2.n3 104.615
R507 VDD2.n65 VDD2.n3 104.615
R508 VDD2.n66 VDD2.n65 104.615
R509 VDD2.n142 VDD2.n70 93.5791
R510 VDD2.n142 VDD2.n141 52.549
R511 VDD2.n96 VDD2.t0 52.3082
R512 VDD2.n25 VDD2.t1 52.3082
R513 VDD2.n95 VDD2.n94 15.6677
R514 VDD2.n24 VDD2.n23 15.6677
R515 VDD2.n139 VDD2.n138 12.8005
R516 VDD2.n98 VDD2.n93 12.8005
R517 VDD2.n27 VDD2.n22 12.8005
R518 VDD2.n68 VDD2.n67 12.8005
R519 VDD2.n135 VDD2.n73 12.0247
R520 VDD2.n99 VDD2.n91 12.0247
R521 VDD2.n28 VDD2.n20 12.0247
R522 VDD2.n64 VDD2.n2 12.0247
R523 VDD2.n134 VDD2.n75 11.249
R524 VDD2.n103 VDD2.n102 11.249
R525 VDD2.n32 VDD2.n31 11.249
R526 VDD2.n63 VDD2.n4 11.249
R527 VDD2.n131 VDD2.n130 10.4732
R528 VDD2.n106 VDD2.n89 10.4732
R529 VDD2.n35 VDD2.n18 10.4732
R530 VDD2.n60 VDD2.n59 10.4732
R531 VDD2.n127 VDD2.n77 9.69747
R532 VDD2.n107 VDD2.n87 9.69747
R533 VDD2.n36 VDD2.n16 9.69747
R534 VDD2.n56 VDD2.n6 9.69747
R535 VDD2.n141 VDD2.n140 9.45567
R536 VDD2.n70 VDD2.n69 9.45567
R537 VDD2.n81 VDD2.n80 9.3005
R538 VDD2.n124 VDD2.n123 9.3005
R539 VDD2.n126 VDD2.n125 9.3005
R540 VDD2.n77 VDD2.n76 9.3005
R541 VDD2.n132 VDD2.n131 9.3005
R542 VDD2.n134 VDD2.n133 9.3005
R543 VDD2.n73 VDD2.n72 9.3005
R544 VDD2.n140 VDD2.n139 9.3005
R545 VDD2.n118 VDD2.n117 9.3005
R546 VDD2.n116 VDD2.n115 9.3005
R547 VDD2.n85 VDD2.n84 9.3005
R548 VDD2.n110 VDD2.n109 9.3005
R549 VDD2.n108 VDD2.n107 9.3005
R550 VDD2.n89 VDD2.n88 9.3005
R551 VDD2.n102 VDD2.n101 9.3005
R552 VDD2.n100 VDD2.n99 9.3005
R553 VDD2.n93 VDD2.n92 9.3005
R554 VDD2.n45 VDD2.n44 9.3005
R555 VDD2.n14 VDD2.n13 9.3005
R556 VDD2.n39 VDD2.n38 9.3005
R557 VDD2.n37 VDD2.n36 9.3005
R558 VDD2.n18 VDD2.n17 9.3005
R559 VDD2.n31 VDD2.n30 9.3005
R560 VDD2.n29 VDD2.n28 9.3005
R561 VDD2.n22 VDD2.n21 9.3005
R562 VDD2.n47 VDD2.n46 9.3005
R563 VDD2.n10 VDD2.n9 9.3005
R564 VDD2.n53 VDD2.n52 9.3005
R565 VDD2.n55 VDD2.n54 9.3005
R566 VDD2.n6 VDD2.n5 9.3005
R567 VDD2.n61 VDD2.n60 9.3005
R568 VDD2.n63 VDD2.n62 9.3005
R569 VDD2.n2 VDD2.n1 9.3005
R570 VDD2.n69 VDD2.n68 9.3005
R571 VDD2.n126 VDD2.n79 8.92171
R572 VDD2.n111 VDD2.n110 8.92171
R573 VDD2.n40 VDD2.n39 8.92171
R574 VDD2.n55 VDD2.n8 8.92171
R575 VDD2.n141 VDD2.n71 8.2187
R576 VDD2.n70 VDD2.n0 8.2187
R577 VDD2.n123 VDD2.n122 8.14595
R578 VDD2.n114 VDD2.n85 8.14595
R579 VDD2.n43 VDD2.n14 8.14595
R580 VDD2.n52 VDD2.n51 8.14595
R581 VDD2.n119 VDD2.n81 7.3702
R582 VDD2.n115 VDD2.n83 7.3702
R583 VDD2.n44 VDD2.n12 7.3702
R584 VDD2.n48 VDD2.n10 7.3702
R585 VDD2.n119 VDD2.n118 6.59444
R586 VDD2.n118 VDD2.n83 6.59444
R587 VDD2.n47 VDD2.n12 6.59444
R588 VDD2.n48 VDD2.n47 6.59444
R589 VDD2.n122 VDD2.n81 5.81868
R590 VDD2.n115 VDD2.n114 5.81868
R591 VDD2.n44 VDD2.n43 5.81868
R592 VDD2.n51 VDD2.n10 5.81868
R593 VDD2.n139 VDD2.n71 5.3904
R594 VDD2.n68 VDD2.n0 5.3904
R595 VDD2.n123 VDD2.n79 5.04292
R596 VDD2.n111 VDD2.n85 5.04292
R597 VDD2.n40 VDD2.n14 5.04292
R598 VDD2.n52 VDD2.n8 5.04292
R599 VDD2.n23 VDD2.n21 4.38563
R600 VDD2.n94 VDD2.n92 4.38563
R601 VDD2.n127 VDD2.n126 4.26717
R602 VDD2.n110 VDD2.n87 4.26717
R603 VDD2.n39 VDD2.n16 4.26717
R604 VDD2.n56 VDD2.n55 4.26717
R605 VDD2.n130 VDD2.n77 3.49141
R606 VDD2.n107 VDD2.n106 3.49141
R607 VDD2.n36 VDD2.n35 3.49141
R608 VDD2.n59 VDD2.n6 3.49141
R609 VDD2.n131 VDD2.n75 2.71565
R610 VDD2.n103 VDD2.n89 2.71565
R611 VDD2.n32 VDD2.n18 2.71565
R612 VDD2.n60 VDD2.n4 2.71565
R613 VDD2.n135 VDD2.n134 1.93989
R614 VDD2.n102 VDD2.n91 1.93989
R615 VDD2.n31 VDD2.n20 1.93989
R616 VDD2.n64 VDD2.n63 1.93989
R617 VDD2.n138 VDD2.n73 1.16414
R618 VDD2.n99 VDD2.n98 1.16414
R619 VDD2.n28 VDD2.n27 1.16414
R620 VDD2.n67 VDD2.n2 1.16414
R621 VDD2 VDD2.n142 0.787138
R622 VDD2.n95 VDD2.n93 0.388379
R623 VDD2.n24 VDD2.n22 0.388379
R624 VDD2.n140 VDD2.n72 0.155672
R625 VDD2.n133 VDD2.n72 0.155672
R626 VDD2.n133 VDD2.n132 0.155672
R627 VDD2.n132 VDD2.n76 0.155672
R628 VDD2.n125 VDD2.n76 0.155672
R629 VDD2.n125 VDD2.n124 0.155672
R630 VDD2.n124 VDD2.n80 0.155672
R631 VDD2.n117 VDD2.n80 0.155672
R632 VDD2.n117 VDD2.n116 0.155672
R633 VDD2.n116 VDD2.n84 0.155672
R634 VDD2.n109 VDD2.n84 0.155672
R635 VDD2.n109 VDD2.n108 0.155672
R636 VDD2.n108 VDD2.n88 0.155672
R637 VDD2.n101 VDD2.n88 0.155672
R638 VDD2.n101 VDD2.n100 0.155672
R639 VDD2.n100 VDD2.n92 0.155672
R640 VDD2.n29 VDD2.n21 0.155672
R641 VDD2.n30 VDD2.n29 0.155672
R642 VDD2.n30 VDD2.n17 0.155672
R643 VDD2.n37 VDD2.n17 0.155672
R644 VDD2.n38 VDD2.n37 0.155672
R645 VDD2.n38 VDD2.n13 0.155672
R646 VDD2.n45 VDD2.n13 0.155672
R647 VDD2.n46 VDD2.n45 0.155672
R648 VDD2.n46 VDD2.n9 0.155672
R649 VDD2.n53 VDD2.n9 0.155672
R650 VDD2.n54 VDD2.n53 0.155672
R651 VDD2.n54 VDD2.n5 0.155672
R652 VDD2.n61 VDD2.n5 0.155672
R653 VDD2.n62 VDD2.n61 0.155672
R654 VDD2.n62 VDD2.n1 0.155672
R655 VDD2.n69 VDD2.n1 0.155672
R656 B.n742 B.n741 585
R657 B.n743 B.n742 585
R658 B.n308 B.n105 585
R659 B.n307 B.n306 585
R660 B.n305 B.n304 585
R661 B.n303 B.n302 585
R662 B.n301 B.n300 585
R663 B.n299 B.n298 585
R664 B.n297 B.n296 585
R665 B.n295 B.n294 585
R666 B.n293 B.n292 585
R667 B.n291 B.n290 585
R668 B.n289 B.n288 585
R669 B.n287 B.n286 585
R670 B.n285 B.n284 585
R671 B.n283 B.n282 585
R672 B.n281 B.n280 585
R673 B.n279 B.n278 585
R674 B.n277 B.n276 585
R675 B.n275 B.n274 585
R676 B.n273 B.n272 585
R677 B.n271 B.n270 585
R678 B.n269 B.n268 585
R679 B.n267 B.n266 585
R680 B.n265 B.n264 585
R681 B.n263 B.n262 585
R682 B.n261 B.n260 585
R683 B.n259 B.n258 585
R684 B.n257 B.n256 585
R685 B.n255 B.n254 585
R686 B.n253 B.n252 585
R687 B.n251 B.n250 585
R688 B.n249 B.n248 585
R689 B.n247 B.n246 585
R690 B.n245 B.n244 585
R691 B.n243 B.n242 585
R692 B.n241 B.n240 585
R693 B.n239 B.n238 585
R694 B.n237 B.n236 585
R695 B.n235 B.n234 585
R696 B.n233 B.n232 585
R697 B.n231 B.n230 585
R698 B.n229 B.n228 585
R699 B.n227 B.n226 585
R700 B.n225 B.n224 585
R701 B.n223 B.n222 585
R702 B.n221 B.n220 585
R703 B.n218 B.n217 585
R704 B.n216 B.n215 585
R705 B.n214 B.n213 585
R706 B.n212 B.n211 585
R707 B.n210 B.n209 585
R708 B.n208 B.n207 585
R709 B.n206 B.n205 585
R710 B.n204 B.n203 585
R711 B.n202 B.n201 585
R712 B.n200 B.n199 585
R713 B.n198 B.n197 585
R714 B.n196 B.n195 585
R715 B.n194 B.n193 585
R716 B.n192 B.n191 585
R717 B.n190 B.n189 585
R718 B.n188 B.n187 585
R719 B.n186 B.n185 585
R720 B.n184 B.n183 585
R721 B.n182 B.n181 585
R722 B.n180 B.n179 585
R723 B.n178 B.n177 585
R724 B.n176 B.n175 585
R725 B.n174 B.n173 585
R726 B.n172 B.n171 585
R727 B.n170 B.n169 585
R728 B.n168 B.n167 585
R729 B.n166 B.n165 585
R730 B.n164 B.n163 585
R731 B.n162 B.n161 585
R732 B.n160 B.n159 585
R733 B.n158 B.n157 585
R734 B.n156 B.n155 585
R735 B.n154 B.n153 585
R736 B.n152 B.n151 585
R737 B.n150 B.n149 585
R738 B.n148 B.n147 585
R739 B.n146 B.n145 585
R740 B.n144 B.n143 585
R741 B.n142 B.n141 585
R742 B.n140 B.n139 585
R743 B.n138 B.n137 585
R744 B.n136 B.n135 585
R745 B.n134 B.n133 585
R746 B.n132 B.n131 585
R747 B.n130 B.n129 585
R748 B.n128 B.n127 585
R749 B.n126 B.n125 585
R750 B.n124 B.n123 585
R751 B.n122 B.n121 585
R752 B.n120 B.n119 585
R753 B.n118 B.n117 585
R754 B.n116 B.n115 585
R755 B.n114 B.n113 585
R756 B.n112 B.n111 585
R757 B.n53 B.n52 585
R758 B.n740 B.n54 585
R759 B.n744 B.n54 585
R760 B.n739 B.n738 585
R761 B.n738 B.n50 585
R762 B.n737 B.n49 585
R763 B.n750 B.n49 585
R764 B.n736 B.n48 585
R765 B.n751 B.n48 585
R766 B.n735 B.n47 585
R767 B.n752 B.n47 585
R768 B.n734 B.n733 585
R769 B.n733 B.n43 585
R770 B.n732 B.n42 585
R771 B.n758 B.n42 585
R772 B.n731 B.n41 585
R773 B.n759 B.n41 585
R774 B.n730 B.n40 585
R775 B.n760 B.n40 585
R776 B.n729 B.n728 585
R777 B.n728 B.n36 585
R778 B.n727 B.n35 585
R779 B.n766 B.n35 585
R780 B.n726 B.n34 585
R781 B.n767 B.n34 585
R782 B.n725 B.n33 585
R783 B.n768 B.n33 585
R784 B.n724 B.n723 585
R785 B.n723 B.n29 585
R786 B.n722 B.n28 585
R787 B.n774 B.n28 585
R788 B.n721 B.n27 585
R789 B.n775 B.n27 585
R790 B.n720 B.n26 585
R791 B.n776 B.n26 585
R792 B.n719 B.n718 585
R793 B.n718 B.n22 585
R794 B.n717 B.n21 585
R795 B.n782 B.n21 585
R796 B.n716 B.n20 585
R797 B.n783 B.n20 585
R798 B.n715 B.n19 585
R799 B.n784 B.n19 585
R800 B.n714 B.n713 585
R801 B.n713 B.n18 585
R802 B.n712 B.n14 585
R803 B.n790 B.n14 585
R804 B.n711 B.n13 585
R805 B.n791 B.n13 585
R806 B.n710 B.n12 585
R807 B.n792 B.n12 585
R808 B.n709 B.n708 585
R809 B.n708 B.n8 585
R810 B.n707 B.n7 585
R811 B.n798 B.n7 585
R812 B.n706 B.n6 585
R813 B.n799 B.n6 585
R814 B.n705 B.n5 585
R815 B.n800 B.n5 585
R816 B.n704 B.n703 585
R817 B.n703 B.n4 585
R818 B.n702 B.n309 585
R819 B.n702 B.n701 585
R820 B.n692 B.n310 585
R821 B.n311 B.n310 585
R822 B.n694 B.n693 585
R823 B.n695 B.n694 585
R824 B.n691 B.n316 585
R825 B.n316 B.n315 585
R826 B.n690 B.n689 585
R827 B.n689 B.n688 585
R828 B.n318 B.n317 585
R829 B.n681 B.n318 585
R830 B.n680 B.n679 585
R831 B.n682 B.n680 585
R832 B.n678 B.n323 585
R833 B.n323 B.n322 585
R834 B.n677 B.n676 585
R835 B.n676 B.n675 585
R836 B.n325 B.n324 585
R837 B.n326 B.n325 585
R838 B.n668 B.n667 585
R839 B.n669 B.n668 585
R840 B.n666 B.n331 585
R841 B.n331 B.n330 585
R842 B.n665 B.n664 585
R843 B.n664 B.n663 585
R844 B.n333 B.n332 585
R845 B.n334 B.n333 585
R846 B.n656 B.n655 585
R847 B.n657 B.n656 585
R848 B.n654 B.n339 585
R849 B.n339 B.n338 585
R850 B.n653 B.n652 585
R851 B.n652 B.n651 585
R852 B.n341 B.n340 585
R853 B.n342 B.n341 585
R854 B.n644 B.n643 585
R855 B.n645 B.n644 585
R856 B.n642 B.n347 585
R857 B.n347 B.n346 585
R858 B.n641 B.n640 585
R859 B.n640 B.n639 585
R860 B.n349 B.n348 585
R861 B.n350 B.n349 585
R862 B.n632 B.n631 585
R863 B.n633 B.n632 585
R864 B.n630 B.n355 585
R865 B.n355 B.n354 585
R866 B.n629 B.n628 585
R867 B.n628 B.n627 585
R868 B.n357 B.n356 585
R869 B.n358 B.n357 585
R870 B.n620 B.n619 585
R871 B.n621 B.n620 585
R872 B.n361 B.n360 585
R873 B.n418 B.n416 585
R874 B.n419 B.n415 585
R875 B.n419 B.n362 585
R876 B.n422 B.n421 585
R877 B.n423 B.n414 585
R878 B.n425 B.n424 585
R879 B.n427 B.n413 585
R880 B.n430 B.n429 585
R881 B.n431 B.n412 585
R882 B.n433 B.n432 585
R883 B.n435 B.n411 585
R884 B.n438 B.n437 585
R885 B.n439 B.n410 585
R886 B.n441 B.n440 585
R887 B.n443 B.n409 585
R888 B.n446 B.n445 585
R889 B.n447 B.n408 585
R890 B.n449 B.n448 585
R891 B.n451 B.n407 585
R892 B.n454 B.n453 585
R893 B.n455 B.n406 585
R894 B.n457 B.n456 585
R895 B.n459 B.n405 585
R896 B.n462 B.n461 585
R897 B.n463 B.n404 585
R898 B.n465 B.n464 585
R899 B.n467 B.n403 585
R900 B.n470 B.n469 585
R901 B.n471 B.n402 585
R902 B.n473 B.n472 585
R903 B.n475 B.n401 585
R904 B.n478 B.n477 585
R905 B.n479 B.n400 585
R906 B.n481 B.n480 585
R907 B.n483 B.n399 585
R908 B.n486 B.n485 585
R909 B.n487 B.n398 585
R910 B.n489 B.n488 585
R911 B.n491 B.n397 585
R912 B.n494 B.n493 585
R913 B.n495 B.n396 585
R914 B.n497 B.n496 585
R915 B.n499 B.n395 585
R916 B.n502 B.n501 585
R917 B.n503 B.n394 585
R918 B.n508 B.n507 585
R919 B.n510 B.n393 585
R920 B.n513 B.n512 585
R921 B.n514 B.n392 585
R922 B.n516 B.n515 585
R923 B.n518 B.n391 585
R924 B.n521 B.n520 585
R925 B.n522 B.n390 585
R926 B.n524 B.n523 585
R927 B.n526 B.n389 585
R928 B.n529 B.n528 585
R929 B.n530 B.n385 585
R930 B.n532 B.n531 585
R931 B.n534 B.n384 585
R932 B.n537 B.n536 585
R933 B.n538 B.n383 585
R934 B.n540 B.n539 585
R935 B.n542 B.n382 585
R936 B.n545 B.n544 585
R937 B.n546 B.n381 585
R938 B.n548 B.n547 585
R939 B.n550 B.n380 585
R940 B.n553 B.n552 585
R941 B.n554 B.n379 585
R942 B.n556 B.n555 585
R943 B.n558 B.n378 585
R944 B.n561 B.n560 585
R945 B.n562 B.n377 585
R946 B.n564 B.n563 585
R947 B.n566 B.n376 585
R948 B.n569 B.n568 585
R949 B.n570 B.n375 585
R950 B.n572 B.n571 585
R951 B.n574 B.n374 585
R952 B.n577 B.n576 585
R953 B.n578 B.n373 585
R954 B.n580 B.n579 585
R955 B.n582 B.n372 585
R956 B.n585 B.n584 585
R957 B.n586 B.n371 585
R958 B.n588 B.n587 585
R959 B.n590 B.n370 585
R960 B.n593 B.n592 585
R961 B.n594 B.n369 585
R962 B.n596 B.n595 585
R963 B.n598 B.n368 585
R964 B.n601 B.n600 585
R965 B.n602 B.n367 585
R966 B.n604 B.n603 585
R967 B.n606 B.n366 585
R968 B.n609 B.n608 585
R969 B.n610 B.n365 585
R970 B.n612 B.n611 585
R971 B.n614 B.n364 585
R972 B.n617 B.n616 585
R973 B.n618 B.n363 585
R974 B.n623 B.n622 585
R975 B.n622 B.n621 585
R976 B.n624 B.n359 585
R977 B.n359 B.n358 585
R978 B.n626 B.n625 585
R979 B.n627 B.n626 585
R980 B.n353 B.n352 585
R981 B.n354 B.n353 585
R982 B.n635 B.n634 585
R983 B.n634 B.n633 585
R984 B.n636 B.n351 585
R985 B.n351 B.n350 585
R986 B.n638 B.n637 585
R987 B.n639 B.n638 585
R988 B.n345 B.n344 585
R989 B.n346 B.n345 585
R990 B.n647 B.n646 585
R991 B.n646 B.n645 585
R992 B.n648 B.n343 585
R993 B.n343 B.n342 585
R994 B.n650 B.n649 585
R995 B.n651 B.n650 585
R996 B.n337 B.n336 585
R997 B.n338 B.n337 585
R998 B.n659 B.n658 585
R999 B.n658 B.n657 585
R1000 B.n660 B.n335 585
R1001 B.n335 B.n334 585
R1002 B.n662 B.n661 585
R1003 B.n663 B.n662 585
R1004 B.n329 B.n328 585
R1005 B.n330 B.n329 585
R1006 B.n671 B.n670 585
R1007 B.n670 B.n669 585
R1008 B.n672 B.n327 585
R1009 B.n327 B.n326 585
R1010 B.n674 B.n673 585
R1011 B.n675 B.n674 585
R1012 B.n321 B.n320 585
R1013 B.n322 B.n321 585
R1014 B.n684 B.n683 585
R1015 B.n683 B.n682 585
R1016 B.n685 B.n319 585
R1017 B.n681 B.n319 585
R1018 B.n687 B.n686 585
R1019 B.n688 B.n687 585
R1020 B.n314 B.n313 585
R1021 B.n315 B.n314 585
R1022 B.n697 B.n696 585
R1023 B.n696 B.n695 585
R1024 B.n698 B.n312 585
R1025 B.n312 B.n311 585
R1026 B.n700 B.n699 585
R1027 B.n701 B.n700 585
R1028 B.n2 B.n0 585
R1029 B.n4 B.n2 585
R1030 B.n3 B.n1 585
R1031 B.n799 B.n3 585
R1032 B.n797 B.n796 585
R1033 B.n798 B.n797 585
R1034 B.n795 B.n9 585
R1035 B.n9 B.n8 585
R1036 B.n794 B.n793 585
R1037 B.n793 B.n792 585
R1038 B.n11 B.n10 585
R1039 B.n791 B.n11 585
R1040 B.n789 B.n788 585
R1041 B.n790 B.n789 585
R1042 B.n787 B.n15 585
R1043 B.n18 B.n15 585
R1044 B.n786 B.n785 585
R1045 B.n785 B.n784 585
R1046 B.n17 B.n16 585
R1047 B.n783 B.n17 585
R1048 B.n781 B.n780 585
R1049 B.n782 B.n781 585
R1050 B.n779 B.n23 585
R1051 B.n23 B.n22 585
R1052 B.n778 B.n777 585
R1053 B.n777 B.n776 585
R1054 B.n25 B.n24 585
R1055 B.n775 B.n25 585
R1056 B.n773 B.n772 585
R1057 B.n774 B.n773 585
R1058 B.n771 B.n30 585
R1059 B.n30 B.n29 585
R1060 B.n770 B.n769 585
R1061 B.n769 B.n768 585
R1062 B.n32 B.n31 585
R1063 B.n767 B.n32 585
R1064 B.n765 B.n764 585
R1065 B.n766 B.n765 585
R1066 B.n763 B.n37 585
R1067 B.n37 B.n36 585
R1068 B.n762 B.n761 585
R1069 B.n761 B.n760 585
R1070 B.n39 B.n38 585
R1071 B.n759 B.n39 585
R1072 B.n757 B.n756 585
R1073 B.n758 B.n757 585
R1074 B.n755 B.n44 585
R1075 B.n44 B.n43 585
R1076 B.n754 B.n753 585
R1077 B.n753 B.n752 585
R1078 B.n46 B.n45 585
R1079 B.n751 B.n46 585
R1080 B.n749 B.n748 585
R1081 B.n750 B.n749 585
R1082 B.n747 B.n51 585
R1083 B.n51 B.n50 585
R1084 B.n746 B.n745 585
R1085 B.n745 B.n744 585
R1086 B.n802 B.n801 585
R1087 B.n801 B.n800 585
R1088 B.n622 B.n361 497.305
R1089 B.n745 B.n53 497.305
R1090 B.n620 B.n363 497.305
R1091 B.n742 B.n54 497.305
R1092 B.n386 B.t8 371.567
R1093 B.n106 B.t14 371.567
R1094 B.n504 B.t5 371.567
R1095 B.n108 B.t11 371.567
R1096 B.n386 B.t6 314.442
R1097 B.n504 B.t2 314.442
R1098 B.n108 B.t9 314.442
R1099 B.n106 B.t13 314.442
R1100 B.n387 B.t7 306.014
R1101 B.n107 B.t15 306.014
R1102 B.n505 B.t4 306.014
R1103 B.n109 B.t12 306.014
R1104 B.n743 B.n104 256.663
R1105 B.n743 B.n103 256.663
R1106 B.n743 B.n102 256.663
R1107 B.n743 B.n101 256.663
R1108 B.n743 B.n100 256.663
R1109 B.n743 B.n99 256.663
R1110 B.n743 B.n98 256.663
R1111 B.n743 B.n97 256.663
R1112 B.n743 B.n96 256.663
R1113 B.n743 B.n95 256.663
R1114 B.n743 B.n94 256.663
R1115 B.n743 B.n93 256.663
R1116 B.n743 B.n92 256.663
R1117 B.n743 B.n91 256.663
R1118 B.n743 B.n90 256.663
R1119 B.n743 B.n89 256.663
R1120 B.n743 B.n88 256.663
R1121 B.n743 B.n87 256.663
R1122 B.n743 B.n86 256.663
R1123 B.n743 B.n85 256.663
R1124 B.n743 B.n84 256.663
R1125 B.n743 B.n83 256.663
R1126 B.n743 B.n82 256.663
R1127 B.n743 B.n81 256.663
R1128 B.n743 B.n80 256.663
R1129 B.n743 B.n79 256.663
R1130 B.n743 B.n78 256.663
R1131 B.n743 B.n77 256.663
R1132 B.n743 B.n76 256.663
R1133 B.n743 B.n75 256.663
R1134 B.n743 B.n74 256.663
R1135 B.n743 B.n73 256.663
R1136 B.n743 B.n72 256.663
R1137 B.n743 B.n71 256.663
R1138 B.n743 B.n70 256.663
R1139 B.n743 B.n69 256.663
R1140 B.n743 B.n68 256.663
R1141 B.n743 B.n67 256.663
R1142 B.n743 B.n66 256.663
R1143 B.n743 B.n65 256.663
R1144 B.n743 B.n64 256.663
R1145 B.n743 B.n63 256.663
R1146 B.n743 B.n62 256.663
R1147 B.n743 B.n61 256.663
R1148 B.n743 B.n60 256.663
R1149 B.n743 B.n59 256.663
R1150 B.n743 B.n58 256.663
R1151 B.n743 B.n57 256.663
R1152 B.n743 B.n56 256.663
R1153 B.n743 B.n55 256.663
R1154 B.n417 B.n362 256.663
R1155 B.n420 B.n362 256.663
R1156 B.n426 B.n362 256.663
R1157 B.n428 B.n362 256.663
R1158 B.n434 B.n362 256.663
R1159 B.n436 B.n362 256.663
R1160 B.n442 B.n362 256.663
R1161 B.n444 B.n362 256.663
R1162 B.n450 B.n362 256.663
R1163 B.n452 B.n362 256.663
R1164 B.n458 B.n362 256.663
R1165 B.n460 B.n362 256.663
R1166 B.n466 B.n362 256.663
R1167 B.n468 B.n362 256.663
R1168 B.n474 B.n362 256.663
R1169 B.n476 B.n362 256.663
R1170 B.n482 B.n362 256.663
R1171 B.n484 B.n362 256.663
R1172 B.n490 B.n362 256.663
R1173 B.n492 B.n362 256.663
R1174 B.n498 B.n362 256.663
R1175 B.n500 B.n362 256.663
R1176 B.n509 B.n362 256.663
R1177 B.n511 B.n362 256.663
R1178 B.n517 B.n362 256.663
R1179 B.n519 B.n362 256.663
R1180 B.n525 B.n362 256.663
R1181 B.n527 B.n362 256.663
R1182 B.n533 B.n362 256.663
R1183 B.n535 B.n362 256.663
R1184 B.n541 B.n362 256.663
R1185 B.n543 B.n362 256.663
R1186 B.n549 B.n362 256.663
R1187 B.n551 B.n362 256.663
R1188 B.n557 B.n362 256.663
R1189 B.n559 B.n362 256.663
R1190 B.n565 B.n362 256.663
R1191 B.n567 B.n362 256.663
R1192 B.n573 B.n362 256.663
R1193 B.n575 B.n362 256.663
R1194 B.n581 B.n362 256.663
R1195 B.n583 B.n362 256.663
R1196 B.n589 B.n362 256.663
R1197 B.n591 B.n362 256.663
R1198 B.n597 B.n362 256.663
R1199 B.n599 B.n362 256.663
R1200 B.n605 B.n362 256.663
R1201 B.n607 B.n362 256.663
R1202 B.n613 B.n362 256.663
R1203 B.n615 B.n362 256.663
R1204 B.n622 B.n359 163.367
R1205 B.n626 B.n359 163.367
R1206 B.n626 B.n353 163.367
R1207 B.n634 B.n353 163.367
R1208 B.n634 B.n351 163.367
R1209 B.n638 B.n351 163.367
R1210 B.n638 B.n345 163.367
R1211 B.n646 B.n345 163.367
R1212 B.n646 B.n343 163.367
R1213 B.n650 B.n343 163.367
R1214 B.n650 B.n337 163.367
R1215 B.n658 B.n337 163.367
R1216 B.n658 B.n335 163.367
R1217 B.n662 B.n335 163.367
R1218 B.n662 B.n329 163.367
R1219 B.n670 B.n329 163.367
R1220 B.n670 B.n327 163.367
R1221 B.n674 B.n327 163.367
R1222 B.n674 B.n321 163.367
R1223 B.n683 B.n321 163.367
R1224 B.n683 B.n319 163.367
R1225 B.n687 B.n319 163.367
R1226 B.n687 B.n314 163.367
R1227 B.n696 B.n314 163.367
R1228 B.n696 B.n312 163.367
R1229 B.n700 B.n312 163.367
R1230 B.n700 B.n2 163.367
R1231 B.n801 B.n2 163.367
R1232 B.n801 B.n3 163.367
R1233 B.n797 B.n3 163.367
R1234 B.n797 B.n9 163.367
R1235 B.n793 B.n9 163.367
R1236 B.n793 B.n11 163.367
R1237 B.n789 B.n11 163.367
R1238 B.n789 B.n15 163.367
R1239 B.n785 B.n15 163.367
R1240 B.n785 B.n17 163.367
R1241 B.n781 B.n17 163.367
R1242 B.n781 B.n23 163.367
R1243 B.n777 B.n23 163.367
R1244 B.n777 B.n25 163.367
R1245 B.n773 B.n25 163.367
R1246 B.n773 B.n30 163.367
R1247 B.n769 B.n30 163.367
R1248 B.n769 B.n32 163.367
R1249 B.n765 B.n32 163.367
R1250 B.n765 B.n37 163.367
R1251 B.n761 B.n37 163.367
R1252 B.n761 B.n39 163.367
R1253 B.n757 B.n39 163.367
R1254 B.n757 B.n44 163.367
R1255 B.n753 B.n44 163.367
R1256 B.n753 B.n46 163.367
R1257 B.n749 B.n46 163.367
R1258 B.n749 B.n51 163.367
R1259 B.n745 B.n51 163.367
R1260 B.n419 B.n418 163.367
R1261 B.n421 B.n419 163.367
R1262 B.n425 B.n414 163.367
R1263 B.n429 B.n427 163.367
R1264 B.n433 B.n412 163.367
R1265 B.n437 B.n435 163.367
R1266 B.n441 B.n410 163.367
R1267 B.n445 B.n443 163.367
R1268 B.n449 B.n408 163.367
R1269 B.n453 B.n451 163.367
R1270 B.n457 B.n406 163.367
R1271 B.n461 B.n459 163.367
R1272 B.n465 B.n404 163.367
R1273 B.n469 B.n467 163.367
R1274 B.n473 B.n402 163.367
R1275 B.n477 B.n475 163.367
R1276 B.n481 B.n400 163.367
R1277 B.n485 B.n483 163.367
R1278 B.n489 B.n398 163.367
R1279 B.n493 B.n491 163.367
R1280 B.n497 B.n396 163.367
R1281 B.n501 B.n499 163.367
R1282 B.n508 B.n394 163.367
R1283 B.n512 B.n510 163.367
R1284 B.n516 B.n392 163.367
R1285 B.n520 B.n518 163.367
R1286 B.n524 B.n390 163.367
R1287 B.n528 B.n526 163.367
R1288 B.n532 B.n385 163.367
R1289 B.n536 B.n534 163.367
R1290 B.n540 B.n383 163.367
R1291 B.n544 B.n542 163.367
R1292 B.n548 B.n381 163.367
R1293 B.n552 B.n550 163.367
R1294 B.n556 B.n379 163.367
R1295 B.n560 B.n558 163.367
R1296 B.n564 B.n377 163.367
R1297 B.n568 B.n566 163.367
R1298 B.n572 B.n375 163.367
R1299 B.n576 B.n574 163.367
R1300 B.n580 B.n373 163.367
R1301 B.n584 B.n582 163.367
R1302 B.n588 B.n371 163.367
R1303 B.n592 B.n590 163.367
R1304 B.n596 B.n369 163.367
R1305 B.n600 B.n598 163.367
R1306 B.n604 B.n367 163.367
R1307 B.n608 B.n606 163.367
R1308 B.n612 B.n365 163.367
R1309 B.n616 B.n614 163.367
R1310 B.n620 B.n357 163.367
R1311 B.n628 B.n357 163.367
R1312 B.n628 B.n355 163.367
R1313 B.n632 B.n355 163.367
R1314 B.n632 B.n349 163.367
R1315 B.n640 B.n349 163.367
R1316 B.n640 B.n347 163.367
R1317 B.n644 B.n347 163.367
R1318 B.n644 B.n341 163.367
R1319 B.n652 B.n341 163.367
R1320 B.n652 B.n339 163.367
R1321 B.n656 B.n339 163.367
R1322 B.n656 B.n333 163.367
R1323 B.n664 B.n333 163.367
R1324 B.n664 B.n331 163.367
R1325 B.n668 B.n331 163.367
R1326 B.n668 B.n325 163.367
R1327 B.n676 B.n325 163.367
R1328 B.n676 B.n323 163.367
R1329 B.n680 B.n323 163.367
R1330 B.n680 B.n318 163.367
R1331 B.n689 B.n318 163.367
R1332 B.n689 B.n316 163.367
R1333 B.n694 B.n316 163.367
R1334 B.n694 B.n310 163.367
R1335 B.n702 B.n310 163.367
R1336 B.n703 B.n702 163.367
R1337 B.n703 B.n5 163.367
R1338 B.n6 B.n5 163.367
R1339 B.n7 B.n6 163.367
R1340 B.n708 B.n7 163.367
R1341 B.n708 B.n12 163.367
R1342 B.n13 B.n12 163.367
R1343 B.n14 B.n13 163.367
R1344 B.n713 B.n14 163.367
R1345 B.n713 B.n19 163.367
R1346 B.n20 B.n19 163.367
R1347 B.n21 B.n20 163.367
R1348 B.n718 B.n21 163.367
R1349 B.n718 B.n26 163.367
R1350 B.n27 B.n26 163.367
R1351 B.n28 B.n27 163.367
R1352 B.n723 B.n28 163.367
R1353 B.n723 B.n33 163.367
R1354 B.n34 B.n33 163.367
R1355 B.n35 B.n34 163.367
R1356 B.n728 B.n35 163.367
R1357 B.n728 B.n40 163.367
R1358 B.n41 B.n40 163.367
R1359 B.n42 B.n41 163.367
R1360 B.n733 B.n42 163.367
R1361 B.n733 B.n47 163.367
R1362 B.n48 B.n47 163.367
R1363 B.n49 B.n48 163.367
R1364 B.n738 B.n49 163.367
R1365 B.n738 B.n54 163.367
R1366 B.n113 B.n112 163.367
R1367 B.n117 B.n116 163.367
R1368 B.n121 B.n120 163.367
R1369 B.n125 B.n124 163.367
R1370 B.n129 B.n128 163.367
R1371 B.n133 B.n132 163.367
R1372 B.n137 B.n136 163.367
R1373 B.n141 B.n140 163.367
R1374 B.n145 B.n144 163.367
R1375 B.n149 B.n148 163.367
R1376 B.n153 B.n152 163.367
R1377 B.n157 B.n156 163.367
R1378 B.n161 B.n160 163.367
R1379 B.n165 B.n164 163.367
R1380 B.n169 B.n168 163.367
R1381 B.n173 B.n172 163.367
R1382 B.n177 B.n176 163.367
R1383 B.n181 B.n180 163.367
R1384 B.n185 B.n184 163.367
R1385 B.n189 B.n188 163.367
R1386 B.n193 B.n192 163.367
R1387 B.n197 B.n196 163.367
R1388 B.n201 B.n200 163.367
R1389 B.n205 B.n204 163.367
R1390 B.n209 B.n208 163.367
R1391 B.n213 B.n212 163.367
R1392 B.n217 B.n216 163.367
R1393 B.n222 B.n221 163.367
R1394 B.n226 B.n225 163.367
R1395 B.n230 B.n229 163.367
R1396 B.n234 B.n233 163.367
R1397 B.n238 B.n237 163.367
R1398 B.n242 B.n241 163.367
R1399 B.n246 B.n245 163.367
R1400 B.n250 B.n249 163.367
R1401 B.n254 B.n253 163.367
R1402 B.n258 B.n257 163.367
R1403 B.n262 B.n261 163.367
R1404 B.n266 B.n265 163.367
R1405 B.n270 B.n269 163.367
R1406 B.n274 B.n273 163.367
R1407 B.n278 B.n277 163.367
R1408 B.n282 B.n281 163.367
R1409 B.n286 B.n285 163.367
R1410 B.n290 B.n289 163.367
R1411 B.n294 B.n293 163.367
R1412 B.n298 B.n297 163.367
R1413 B.n302 B.n301 163.367
R1414 B.n306 B.n305 163.367
R1415 B.n742 B.n105 163.367
R1416 B.n621 B.n362 72.4891
R1417 B.n744 B.n743 72.4891
R1418 B.n417 B.n361 71.676
R1419 B.n421 B.n420 71.676
R1420 B.n426 B.n425 71.676
R1421 B.n429 B.n428 71.676
R1422 B.n434 B.n433 71.676
R1423 B.n437 B.n436 71.676
R1424 B.n442 B.n441 71.676
R1425 B.n445 B.n444 71.676
R1426 B.n450 B.n449 71.676
R1427 B.n453 B.n452 71.676
R1428 B.n458 B.n457 71.676
R1429 B.n461 B.n460 71.676
R1430 B.n466 B.n465 71.676
R1431 B.n469 B.n468 71.676
R1432 B.n474 B.n473 71.676
R1433 B.n477 B.n476 71.676
R1434 B.n482 B.n481 71.676
R1435 B.n485 B.n484 71.676
R1436 B.n490 B.n489 71.676
R1437 B.n493 B.n492 71.676
R1438 B.n498 B.n497 71.676
R1439 B.n501 B.n500 71.676
R1440 B.n509 B.n508 71.676
R1441 B.n512 B.n511 71.676
R1442 B.n517 B.n516 71.676
R1443 B.n520 B.n519 71.676
R1444 B.n525 B.n524 71.676
R1445 B.n528 B.n527 71.676
R1446 B.n533 B.n532 71.676
R1447 B.n536 B.n535 71.676
R1448 B.n541 B.n540 71.676
R1449 B.n544 B.n543 71.676
R1450 B.n549 B.n548 71.676
R1451 B.n552 B.n551 71.676
R1452 B.n557 B.n556 71.676
R1453 B.n560 B.n559 71.676
R1454 B.n565 B.n564 71.676
R1455 B.n568 B.n567 71.676
R1456 B.n573 B.n572 71.676
R1457 B.n576 B.n575 71.676
R1458 B.n581 B.n580 71.676
R1459 B.n584 B.n583 71.676
R1460 B.n589 B.n588 71.676
R1461 B.n592 B.n591 71.676
R1462 B.n597 B.n596 71.676
R1463 B.n600 B.n599 71.676
R1464 B.n605 B.n604 71.676
R1465 B.n608 B.n607 71.676
R1466 B.n613 B.n612 71.676
R1467 B.n616 B.n615 71.676
R1468 B.n55 B.n53 71.676
R1469 B.n113 B.n56 71.676
R1470 B.n117 B.n57 71.676
R1471 B.n121 B.n58 71.676
R1472 B.n125 B.n59 71.676
R1473 B.n129 B.n60 71.676
R1474 B.n133 B.n61 71.676
R1475 B.n137 B.n62 71.676
R1476 B.n141 B.n63 71.676
R1477 B.n145 B.n64 71.676
R1478 B.n149 B.n65 71.676
R1479 B.n153 B.n66 71.676
R1480 B.n157 B.n67 71.676
R1481 B.n161 B.n68 71.676
R1482 B.n165 B.n69 71.676
R1483 B.n169 B.n70 71.676
R1484 B.n173 B.n71 71.676
R1485 B.n177 B.n72 71.676
R1486 B.n181 B.n73 71.676
R1487 B.n185 B.n74 71.676
R1488 B.n189 B.n75 71.676
R1489 B.n193 B.n76 71.676
R1490 B.n197 B.n77 71.676
R1491 B.n201 B.n78 71.676
R1492 B.n205 B.n79 71.676
R1493 B.n209 B.n80 71.676
R1494 B.n213 B.n81 71.676
R1495 B.n217 B.n82 71.676
R1496 B.n222 B.n83 71.676
R1497 B.n226 B.n84 71.676
R1498 B.n230 B.n85 71.676
R1499 B.n234 B.n86 71.676
R1500 B.n238 B.n87 71.676
R1501 B.n242 B.n88 71.676
R1502 B.n246 B.n89 71.676
R1503 B.n250 B.n90 71.676
R1504 B.n254 B.n91 71.676
R1505 B.n258 B.n92 71.676
R1506 B.n262 B.n93 71.676
R1507 B.n266 B.n94 71.676
R1508 B.n270 B.n95 71.676
R1509 B.n274 B.n96 71.676
R1510 B.n278 B.n97 71.676
R1511 B.n282 B.n98 71.676
R1512 B.n286 B.n99 71.676
R1513 B.n290 B.n100 71.676
R1514 B.n294 B.n101 71.676
R1515 B.n298 B.n102 71.676
R1516 B.n302 B.n103 71.676
R1517 B.n306 B.n104 71.676
R1518 B.n105 B.n104 71.676
R1519 B.n305 B.n103 71.676
R1520 B.n301 B.n102 71.676
R1521 B.n297 B.n101 71.676
R1522 B.n293 B.n100 71.676
R1523 B.n289 B.n99 71.676
R1524 B.n285 B.n98 71.676
R1525 B.n281 B.n97 71.676
R1526 B.n277 B.n96 71.676
R1527 B.n273 B.n95 71.676
R1528 B.n269 B.n94 71.676
R1529 B.n265 B.n93 71.676
R1530 B.n261 B.n92 71.676
R1531 B.n257 B.n91 71.676
R1532 B.n253 B.n90 71.676
R1533 B.n249 B.n89 71.676
R1534 B.n245 B.n88 71.676
R1535 B.n241 B.n87 71.676
R1536 B.n237 B.n86 71.676
R1537 B.n233 B.n85 71.676
R1538 B.n229 B.n84 71.676
R1539 B.n225 B.n83 71.676
R1540 B.n221 B.n82 71.676
R1541 B.n216 B.n81 71.676
R1542 B.n212 B.n80 71.676
R1543 B.n208 B.n79 71.676
R1544 B.n204 B.n78 71.676
R1545 B.n200 B.n77 71.676
R1546 B.n196 B.n76 71.676
R1547 B.n192 B.n75 71.676
R1548 B.n188 B.n74 71.676
R1549 B.n184 B.n73 71.676
R1550 B.n180 B.n72 71.676
R1551 B.n176 B.n71 71.676
R1552 B.n172 B.n70 71.676
R1553 B.n168 B.n69 71.676
R1554 B.n164 B.n68 71.676
R1555 B.n160 B.n67 71.676
R1556 B.n156 B.n66 71.676
R1557 B.n152 B.n65 71.676
R1558 B.n148 B.n64 71.676
R1559 B.n144 B.n63 71.676
R1560 B.n140 B.n62 71.676
R1561 B.n136 B.n61 71.676
R1562 B.n132 B.n60 71.676
R1563 B.n128 B.n59 71.676
R1564 B.n124 B.n58 71.676
R1565 B.n120 B.n57 71.676
R1566 B.n116 B.n56 71.676
R1567 B.n112 B.n55 71.676
R1568 B.n418 B.n417 71.676
R1569 B.n420 B.n414 71.676
R1570 B.n427 B.n426 71.676
R1571 B.n428 B.n412 71.676
R1572 B.n435 B.n434 71.676
R1573 B.n436 B.n410 71.676
R1574 B.n443 B.n442 71.676
R1575 B.n444 B.n408 71.676
R1576 B.n451 B.n450 71.676
R1577 B.n452 B.n406 71.676
R1578 B.n459 B.n458 71.676
R1579 B.n460 B.n404 71.676
R1580 B.n467 B.n466 71.676
R1581 B.n468 B.n402 71.676
R1582 B.n475 B.n474 71.676
R1583 B.n476 B.n400 71.676
R1584 B.n483 B.n482 71.676
R1585 B.n484 B.n398 71.676
R1586 B.n491 B.n490 71.676
R1587 B.n492 B.n396 71.676
R1588 B.n499 B.n498 71.676
R1589 B.n500 B.n394 71.676
R1590 B.n510 B.n509 71.676
R1591 B.n511 B.n392 71.676
R1592 B.n518 B.n517 71.676
R1593 B.n519 B.n390 71.676
R1594 B.n526 B.n525 71.676
R1595 B.n527 B.n385 71.676
R1596 B.n534 B.n533 71.676
R1597 B.n535 B.n383 71.676
R1598 B.n542 B.n541 71.676
R1599 B.n543 B.n381 71.676
R1600 B.n550 B.n549 71.676
R1601 B.n551 B.n379 71.676
R1602 B.n558 B.n557 71.676
R1603 B.n559 B.n377 71.676
R1604 B.n566 B.n565 71.676
R1605 B.n567 B.n375 71.676
R1606 B.n574 B.n573 71.676
R1607 B.n575 B.n373 71.676
R1608 B.n582 B.n581 71.676
R1609 B.n583 B.n371 71.676
R1610 B.n590 B.n589 71.676
R1611 B.n591 B.n369 71.676
R1612 B.n598 B.n597 71.676
R1613 B.n599 B.n367 71.676
R1614 B.n606 B.n605 71.676
R1615 B.n607 B.n365 71.676
R1616 B.n614 B.n613 71.676
R1617 B.n615 B.n363 71.676
R1618 B.n387 B.n386 65.552
R1619 B.n505 B.n504 65.552
R1620 B.n109 B.n108 65.552
R1621 B.n107 B.n106 65.552
R1622 B.n388 B.n387 59.5399
R1623 B.n506 B.n505 59.5399
R1624 B.n110 B.n109 59.5399
R1625 B.n219 B.n107 59.5399
R1626 B.n621 B.n358 40.0755
R1627 B.n627 B.n358 40.0755
R1628 B.n627 B.n354 40.0755
R1629 B.n633 B.n354 40.0755
R1630 B.n633 B.n350 40.0755
R1631 B.n639 B.n350 40.0755
R1632 B.n639 B.n346 40.0755
R1633 B.n645 B.n346 40.0755
R1634 B.n651 B.n342 40.0755
R1635 B.n651 B.n338 40.0755
R1636 B.n657 B.n338 40.0755
R1637 B.n657 B.n334 40.0755
R1638 B.n663 B.n334 40.0755
R1639 B.n663 B.n330 40.0755
R1640 B.n669 B.n330 40.0755
R1641 B.n669 B.n326 40.0755
R1642 B.n675 B.n326 40.0755
R1643 B.n675 B.n322 40.0755
R1644 B.n682 B.n322 40.0755
R1645 B.n682 B.n681 40.0755
R1646 B.n688 B.n315 40.0755
R1647 B.n695 B.n315 40.0755
R1648 B.n695 B.n311 40.0755
R1649 B.n701 B.n311 40.0755
R1650 B.n701 B.n4 40.0755
R1651 B.n800 B.n4 40.0755
R1652 B.n800 B.n799 40.0755
R1653 B.n799 B.n798 40.0755
R1654 B.n798 B.n8 40.0755
R1655 B.n792 B.n8 40.0755
R1656 B.n792 B.n791 40.0755
R1657 B.n791 B.n790 40.0755
R1658 B.n784 B.n18 40.0755
R1659 B.n784 B.n783 40.0755
R1660 B.n783 B.n782 40.0755
R1661 B.n782 B.n22 40.0755
R1662 B.n776 B.n22 40.0755
R1663 B.n776 B.n775 40.0755
R1664 B.n775 B.n774 40.0755
R1665 B.n774 B.n29 40.0755
R1666 B.n768 B.n29 40.0755
R1667 B.n768 B.n767 40.0755
R1668 B.n767 B.n766 40.0755
R1669 B.n766 B.n36 40.0755
R1670 B.n760 B.n759 40.0755
R1671 B.n759 B.n758 40.0755
R1672 B.n758 B.n43 40.0755
R1673 B.n752 B.n43 40.0755
R1674 B.n752 B.n751 40.0755
R1675 B.n751 B.n750 40.0755
R1676 B.n750 B.n50 40.0755
R1677 B.n744 B.n50 40.0755
R1678 B.n746 B.n52 32.3127
R1679 B.n741 B.n740 32.3127
R1680 B.n619 B.n618 32.3127
R1681 B.n623 B.n360 32.3127
R1682 B.t3 B.n342 28.8781
R1683 B.t10 B.n36 28.8781
R1684 B.n688 B.t1 22.9847
R1685 B.n790 B.t0 22.9847
R1686 B B.n802 18.0485
R1687 B.n681 B.t1 17.0913
R1688 B.n18 B.t0 17.0913
R1689 B.n645 B.t3 11.1979
R1690 B.n760 B.t10 11.1979
R1691 B.n111 B.n52 10.6151
R1692 B.n114 B.n111 10.6151
R1693 B.n115 B.n114 10.6151
R1694 B.n118 B.n115 10.6151
R1695 B.n119 B.n118 10.6151
R1696 B.n122 B.n119 10.6151
R1697 B.n123 B.n122 10.6151
R1698 B.n126 B.n123 10.6151
R1699 B.n127 B.n126 10.6151
R1700 B.n130 B.n127 10.6151
R1701 B.n131 B.n130 10.6151
R1702 B.n134 B.n131 10.6151
R1703 B.n135 B.n134 10.6151
R1704 B.n138 B.n135 10.6151
R1705 B.n139 B.n138 10.6151
R1706 B.n142 B.n139 10.6151
R1707 B.n143 B.n142 10.6151
R1708 B.n146 B.n143 10.6151
R1709 B.n147 B.n146 10.6151
R1710 B.n150 B.n147 10.6151
R1711 B.n151 B.n150 10.6151
R1712 B.n154 B.n151 10.6151
R1713 B.n155 B.n154 10.6151
R1714 B.n158 B.n155 10.6151
R1715 B.n159 B.n158 10.6151
R1716 B.n162 B.n159 10.6151
R1717 B.n163 B.n162 10.6151
R1718 B.n166 B.n163 10.6151
R1719 B.n167 B.n166 10.6151
R1720 B.n170 B.n167 10.6151
R1721 B.n171 B.n170 10.6151
R1722 B.n174 B.n171 10.6151
R1723 B.n175 B.n174 10.6151
R1724 B.n178 B.n175 10.6151
R1725 B.n179 B.n178 10.6151
R1726 B.n182 B.n179 10.6151
R1727 B.n183 B.n182 10.6151
R1728 B.n186 B.n183 10.6151
R1729 B.n187 B.n186 10.6151
R1730 B.n190 B.n187 10.6151
R1731 B.n191 B.n190 10.6151
R1732 B.n194 B.n191 10.6151
R1733 B.n195 B.n194 10.6151
R1734 B.n198 B.n195 10.6151
R1735 B.n199 B.n198 10.6151
R1736 B.n203 B.n202 10.6151
R1737 B.n206 B.n203 10.6151
R1738 B.n207 B.n206 10.6151
R1739 B.n210 B.n207 10.6151
R1740 B.n211 B.n210 10.6151
R1741 B.n214 B.n211 10.6151
R1742 B.n215 B.n214 10.6151
R1743 B.n218 B.n215 10.6151
R1744 B.n223 B.n220 10.6151
R1745 B.n224 B.n223 10.6151
R1746 B.n227 B.n224 10.6151
R1747 B.n228 B.n227 10.6151
R1748 B.n231 B.n228 10.6151
R1749 B.n232 B.n231 10.6151
R1750 B.n235 B.n232 10.6151
R1751 B.n236 B.n235 10.6151
R1752 B.n239 B.n236 10.6151
R1753 B.n240 B.n239 10.6151
R1754 B.n243 B.n240 10.6151
R1755 B.n244 B.n243 10.6151
R1756 B.n247 B.n244 10.6151
R1757 B.n248 B.n247 10.6151
R1758 B.n251 B.n248 10.6151
R1759 B.n252 B.n251 10.6151
R1760 B.n255 B.n252 10.6151
R1761 B.n256 B.n255 10.6151
R1762 B.n259 B.n256 10.6151
R1763 B.n260 B.n259 10.6151
R1764 B.n263 B.n260 10.6151
R1765 B.n264 B.n263 10.6151
R1766 B.n267 B.n264 10.6151
R1767 B.n268 B.n267 10.6151
R1768 B.n271 B.n268 10.6151
R1769 B.n272 B.n271 10.6151
R1770 B.n275 B.n272 10.6151
R1771 B.n276 B.n275 10.6151
R1772 B.n279 B.n276 10.6151
R1773 B.n280 B.n279 10.6151
R1774 B.n283 B.n280 10.6151
R1775 B.n284 B.n283 10.6151
R1776 B.n287 B.n284 10.6151
R1777 B.n288 B.n287 10.6151
R1778 B.n291 B.n288 10.6151
R1779 B.n292 B.n291 10.6151
R1780 B.n295 B.n292 10.6151
R1781 B.n296 B.n295 10.6151
R1782 B.n299 B.n296 10.6151
R1783 B.n300 B.n299 10.6151
R1784 B.n303 B.n300 10.6151
R1785 B.n304 B.n303 10.6151
R1786 B.n307 B.n304 10.6151
R1787 B.n308 B.n307 10.6151
R1788 B.n741 B.n308 10.6151
R1789 B.n619 B.n356 10.6151
R1790 B.n629 B.n356 10.6151
R1791 B.n630 B.n629 10.6151
R1792 B.n631 B.n630 10.6151
R1793 B.n631 B.n348 10.6151
R1794 B.n641 B.n348 10.6151
R1795 B.n642 B.n641 10.6151
R1796 B.n643 B.n642 10.6151
R1797 B.n643 B.n340 10.6151
R1798 B.n653 B.n340 10.6151
R1799 B.n654 B.n653 10.6151
R1800 B.n655 B.n654 10.6151
R1801 B.n655 B.n332 10.6151
R1802 B.n665 B.n332 10.6151
R1803 B.n666 B.n665 10.6151
R1804 B.n667 B.n666 10.6151
R1805 B.n667 B.n324 10.6151
R1806 B.n677 B.n324 10.6151
R1807 B.n678 B.n677 10.6151
R1808 B.n679 B.n678 10.6151
R1809 B.n679 B.n317 10.6151
R1810 B.n690 B.n317 10.6151
R1811 B.n691 B.n690 10.6151
R1812 B.n693 B.n691 10.6151
R1813 B.n693 B.n692 10.6151
R1814 B.n692 B.n309 10.6151
R1815 B.n704 B.n309 10.6151
R1816 B.n705 B.n704 10.6151
R1817 B.n706 B.n705 10.6151
R1818 B.n707 B.n706 10.6151
R1819 B.n709 B.n707 10.6151
R1820 B.n710 B.n709 10.6151
R1821 B.n711 B.n710 10.6151
R1822 B.n712 B.n711 10.6151
R1823 B.n714 B.n712 10.6151
R1824 B.n715 B.n714 10.6151
R1825 B.n716 B.n715 10.6151
R1826 B.n717 B.n716 10.6151
R1827 B.n719 B.n717 10.6151
R1828 B.n720 B.n719 10.6151
R1829 B.n721 B.n720 10.6151
R1830 B.n722 B.n721 10.6151
R1831 B.n724 B.n722 10.6151
R1832 B.n725 B.n724 10.6151
R1833 B.n726 B.n725 10.6151
R1834 B.n727 B.n726 10.6151
R1835 B.n729 B.n727 10.6151
R1836 B.n730 B.n729 10.6151
R1837 B.n731 B.n730 10.6151
R1838 B.n732 B.n731 10.6151
R1839 B.n734 B.n732 10.6151
R1840 B.n735 B.n734 10.6151
R1841 B.n736 B.n735 10.6151
R1842 B.n737 B.n736 10.6151
R1843 B.n739 B.n737 10.6151
R1844 B.n740 B.n739 10.6151
R1845 B.n416 B.n360 10.6151
R1846 B.n416 B.n415 10.6151
R1847 B.n422 B.n415 10.6151
R1848 B.n423 B.n422 10.6151
R1849 B.n424 B.n423 10.6151
R1850 B.n424 B.n413 10.6151
R1851 B.n430 B.n413 10.6151
R1852 B.n431 B.n430 10.6151
R1853 B.n432 B.n431 10.6151
R1854 B.n432 B.n411 10.6151
R1855 B.n438 B.n411 10.6151
R1856 B.n439 B.n438 10.6151
R1857 B.n440 B.n439 10.6151
R1858 B.n440 B.n409 10.6151
R1859 B.n446 B.n409 10.6151
R1860 B.n447 B.n446 10.6151
R1861 B.n448 B.n447 10.6151
R1862 B.n448 B.n407 10.6151
R1863 B.n454 B.n407 10.6151
R1864 B.n455 B.n454 10.6151
R1865 B.n456 B.n455 10.6151
R1866 B.n456 B.n405 10.6151
R1867 B.n462 B.n405 10.6151
R1868 B.n463 B.n462 10.6151
R1869 B.n464 B.n463 10.6151
R1870 B.n464 B.n403 10.6151
R1871 B.n470 B.n403 10.6151
R1872 B.n471 B.n470 10.6151
R1873 B.n472 B.n471 10.6151
R1874 B.n472 B.n401 10.6151
R1875 B.n478 B.n401 10.6151
R1876 B.n479 B.n478 10.6151
R1877 B.n480 B.n479 10.6151
R1878 B.n480 B.n399 10.6151
R1879 B.n486 B.n399 10.6151
R1880 B.n487 B.n486 10.6151
R1881 B.n488 B.n487 10.6151
R1882 B.n488 B.n397 10.6151
R1883 B.n494 B.n397 10.6151
R1884 B.n495 B.n494 10.6151
R1885 B.n496 B.n495 10.6151
R1886 B.n496 B.n395 10.6151
R1887 B.n502 B.n395 10.6151
R1888 B.n503 B.n502 10.6151
R1889 B.n507 B.n503 10.6151
R1890 B.n513 B.n393 10.6151
R1891 B.n514 B.n513 10.6151
R1892 B.n515 B.n514 10.6151
R1893 B.n515 B.n391 10.6151
R1894 B.n521 B.n391 10.6151
R1895 B.n522 B.n521 10.6151
R1896 B.n523 B.n522 10.6151
R1897 B.n523 B.n389 10.6151
R1898 B.n530 B.n529 10.6151
R1899 B.n531 B.n530 10.6151
R1900 B.n531 B.n384 10.6151
R1901 B.n537 B.n384 10.6151
R1902 B.n538 B.n537 10.6151
R1903 B.n539 B.n538 10.6151
R1904 B.n539 B.n382 10.6151
R1905 B.n545 B.n382 10.6151
R1906 B.n546 B.n545 10.6151
R1907 B.n547 B.n546 10.6151
R1908 B.n547 B.n380 10.6151
R1909 B.n553 B.n380 10.6151
R1910 B.n554 B.n553 10.6151
R1911 B.n555 B.n554 10.6151
R1912 B.n555 B.n378 10.6151
R1913 B.n561 B.n378 10.6151
R1914 B.n562 B.n561 10.6151
R1915 B.n563 B.n562 10.6151
R1916 B.n563 B.n376 10.6151
R1917 B.n569 B.n376 10.6151
R1918 B.n570 B.n569 10.6151
R1919 B.n571 B.n570 10.6151
R1920 B.n571 B.n374 10.6151
R1921 B.n577 B.n374 10.6151
R1922 B.n578 B.n577 10.6151
R1923 B.n579 B.n578 10.6151
R1924 B.n579 B.n372 10.6151
R1925 B.n585 B.n372 10.6151
R1926 B.n586 B.n585 10.6151
R1927 B.n587 B.n586 10.6151
R1928 B.n587 B.n370 10.6151
R1929 B.n593 B.n370 10.6151
R1930 B.n594 B.n593 10.6151
R1931 B.n595 B.n594 10.6151
R1932 B.n595 B.n368 10.6151
R1933 B.n601 B.n368 10.6151
R1934 B.n602 B.n601 10.6151
R1935 B.n603 B.n602 10.6151
R1936 B.n603 B.n366 10.6151
R1937 B.n609 B.n366 10.6151
R1938 B.n610 B.n609 10.6151
R1939 B.n611 B.n610 10.6151
R1940 B.n611 B.n364 10.6151
R1941 B.n617 B.n364 10.6151
R1942 B.n618 B.n617 10.6151
R1943 B.n624 B.n623 10.6151
R1944 B.n625 B.n624 10.6151
R1945 B.n625 B.n352 10.6151
R1946 B.n635 B.n352 10.6151
R1947 B.n636 B.n635 10.6151
R1948 B.n637 B.n636 10.6151
R1949 B.n637 B.n344 10.6151
R1950 B.n647 B.n344 10.6151
R1951 B.n648 B.n647 10.6151
R1952 B.n649 B.n648 10.6151
R1953 B.n649 B.n336 10.6151
R1954 B.n659 B.n336 10.6151
R1955 B.n660 B.n659 10.6151
R1956 B.n661 B.n660 10.6151
R1957 B.n661 B.n328 10.6151
R1958 B.n671 B.n328 10.6151
R1959 B.n672 B.n671 10.6151
R1960 B.n673 B.n672 10.6151
R1961 B.n673 B.n320 10.6151
R1962 B.n684 B.n320 10.6151
R1963 B.n685 B.n684 10.6151
R1964 B.n686 B.n685 10.6151
R1965 B.n686 B.n313 10.6151
R1966 B.n697 B.n313 10.6151
R1967 B.n698 B.n697 10.6151
R1968 B.n699 B.n698 10.6151
R1969 B.n699 B.n0 10.6151
R1970 B.n796 B.n1 10.6151
R1971 B.n796 B.n795 10.6151
R1972 B.n795 B.n794 10.6151
R1973 B.n794 B.n10 10.6151
R1974 B.n788 B.n10 10.6151
R1975 B.n788 B.n787 10.6151
R1976 B.n787 B.n786 10.6151
R1977 B.n786 B.n16 10.6151
R1978 B.n780 B.n16 10.6151
R1979 B.n780 B.n779 10.6151
R1980 B.n779 B.n778 10.6151
R1981 B.n778 B.n24 10.6151
R1982 B.n772 B.n24 10.6151
R1983 B.n772 B.n771 10.6151
R1984 B.n771 B.n770 10.6151
R1985 B.n770 B.n31 10.6151
R1986 B.n764 B.n31 10.6151
R1987 B.n764 B.n763 10.6151
R1988 B.n763 B.n762 10.6151
R1989 B.n762 B.n38 10.6151
R1990 B.n756 B.n38 10.6151
R1991 B.n756 B.n755 10.6151
R1992 B.n755 B.n754 10.6151
R1993 B.n754 B.n45 10.6151
R1994 B.n748 B.n45 10.6151
R1995 B.n748 B.n747 10.6151
R1996 B.n747 B.n746 10.6151
R1997 B.n202 B.n110 6.5566
R1998 B.n219 B.n218 6.5566
R1999 B.n506 B.n393 6.5566
R2000 B.n389 B.n388 6.5566
R2001 B.n199 B.n110 4.05904
R2002 B.n220 B.n219 4.05904
R2003 B.n507 B.n506 4.05904
R2004 B.n529 B.n388 4.05904
R2005 B.n802 B.n0 2.81026
R2006 B.n802 B.n1 2.81026
R2007 VP.n0 VP.t0 193.803
R2008 VP.n0 VP.t1 146.899
R2009 VP VP.n0 0.431811
R2010 VDD1.n66 VDD1.n0 214.453
R2011 VDD1.n137 VDD1.n71 214.453
R2012 VDD1.n67 VDD1.n66 185
R2013 VDD1.n65 VDD1.n64 185
R2014 VDD1.n4 VDD1.n3 185
R2015 VDD1.n59 VDD1.n58 185
R2016 VDD1.n57 VDD1.n56 185
R2017 VDD1.n8 VDD1.n7 185
R2018 VDD1.n51 VDD1.n50 185
R2019 VDD1.n49 VDD1.n48 185
R2020 VDD1.n12 VDD1.n11 185
R2021 VDD1.n43 VDD1.n42 185
R2022 VDD1.n41 VDD1.n40 185
R2023 VDD1.n16 VDD1.n15 185
R2024 VDD1.n35 VDD1.n34 185
R2025 VDD1.n33 VDD1.n32 185
R2026 VDD1.n20 VDD1.n19 185
R2027 VDD1.n27 VDD1.n26 185
R2028 VDD1.n25 VDD1.n24 185
R2029 VDD1.n96 VDD1.n95 185
R2030 VDD1.n98 VDD1.n97 185
R2031 VDD1.n91 VDD1.n90 185
R2032 VDD1.n104 VDD1.n103 185
R2033 VDD1.n106 VDD1.n105 185
R2034 VDD1.n87 VDD1.n86 185
R2035 VDD1.n112 VDD1.n111 185
R2036 VDD1.n114 VDD1.n113 185
R2037 VDD1.n83 VDD1.n82 185
R2038 VDD1.n120 VDD1.n119 185
R2039 VDD1.n122 VDD1.n121 185
R2040 VDD1.n79 VDD1.n78 185
R2041 VDD1.n128 VDD1.n127 185
R2042 VDD1.n130 VDD1.n129 185
R2043 VDD1.n75 VDD1.n74 185
R2044 VDD1.n136 VDD1.n135 185
R2045 VDD1.n138 VDD1.n137 185
R2046 VDD1.n94 VDD1.t0 147.659
R2047 VDD1.n23 VDD1.t1 147.659
R2048 VDD1.n66 VDD1.n65 104.615
R2049 VDD1.n65 VDD1.n3 104.615
R2050 VDD1.n58 VDD1.n3 104.615
R2051 VDD1.n58 VDD1.n57 104.615
R2052 VDD1.n57 VDD1.n7 104.615
R2053 VDD1.n50 VDD1.n7 104.615
R2054 VDD1.n50 VDD1.n49 104.615
R2055 VDD1.n49 VDD1.n11 104.615
R2056 VDD1.n42 VDD1.n11 104.615
R2057 VDD1.n42 VDD1.n41 104.615
R2058 VDD1.n41 VDD1.n15 104.615
R2059 VDD1.n34 VDD1.n15 104.615
R2060 VDD1.n34 VDD1.n33 104.615
R2061 VDD1.n33 VDD1.n19 104.615
R2062 VDD1.n26 VDD1.n19 104.615
R2063 VDD1.n26 VDD1.n25 104.615
R2064 VDD1.n97 VDD1.n96 104.615
R2065 VDD1.n97 VDD1.n90 104.615
R2066 VDD1.n104 VDD1.n90 104.615
R2067 VDD1.n105 VDD1.n104 104.615
R2068 VDD1.n105 VDD1.n86 104.615
R2069 VDD1.n112 VDD1.n86 104.615
R2070 VDD1.n113 VDD1.n112 104.615
R2071 VDD1.n113 VDD1.n82 104.615
R2072 VDD1.n120 VDD1.n82 104.615
R2073 VDD1.n121 VDD1.n120 104.615
R2074 VDD1.n121 VDD1.n78 104.615
R2075 VDD1.n128 VDD1.n78 104.615
R2076 VDD1.n129 VDD1.n128 104.615
R2077 VDD1.n129 VDD1.n74 104.615
R2078 VDD1.n136 VDD1.n74 104.615
R2079 VDD1.n137 VDD1.n136 104.615
R2080 VDD1 VDD1.n141 94.8324
R2081 VDD1 VDD1.n70 53.3356
R2082 VDD1.n25 VDD1.t1 52.3082
R2083 VDD1.n96 VDD1.t0 52.3082
R2084 VDD1.n24 VDD1.n23 15.6677
R2085 VDD1.n95 VDD1.n94 15.6677
R2086 VDD1.n68 VDD1.n67 12.8005
R2087 VDD1.n27 VDD1.n22 12.8005
R2088 VDD1.n98 VDD1.n93 12.8005
R2089 VDD1.n139 VDD1.n138 12.8005
R2090 VDD1.n64 VDD1.n2 12.0247
R2091 VDD1.n28 VDD1.n20 12.0247
R2092 VDD1.n99 VDD1.n91 12.0247
R2093 VDD1.n135 VDD1.n73 12.0247
R2094 VDD1.n63 VDD1.n4 11.249
R2095 VDD1.n32 VDD1.n31 11.249
R2096 VDD1.n103 VDD1.n102 11.249
R2097 VDD1.n134 VDD1.n75 11.249
R2098 VDD1.n60 VDD1.n59 10.4732
R2099 VDD1.n35 VDD1.n18 10.4732
R2100 VDD1.n106 VDD1.n89 10.4732
R2101 VDD1.n131 VDD1.n130 10.4732
R2102 VDD1.n56 VDD1.n6 9.69747
R2103 VDD1.n36 VDD1.n16 9.69747
R2104 VDD1.n107 VDD1.n87 9.69747
R2105 VDD1.n127 VDD1.n77 9.69747
R2106 VDD1.n70 VDD1.n69 9.45567
R2107 VDD1.n141 VDD1.n140 9.45567
R2108 VDD1.n10 VDD1.n9 9.3005
R2109 VDD1.n53 VDD1.n52 9.3005
R2110 VDD1.n55 VDD1.n54 9.3005
R2111 VDD1.n6 VDD1.n5 9.3005
R2112 VDD1.n61 VDD1.n60 9.3005
R2113 VDD1.n63 VDD1.n62 9.3005
R2114 VDD1.n2 VDD1.n1 9.3005
R2115 VDD1.n69 VDD1.n68 9.3005
R2116 VDD1.n47 VDD1.n46 9.3005
R2117 VDD1.n45 VDD1.n44 9.3005
R2118 VDD1.n14 VDD1.n13 9.3005
R2119 VDD1.n39 VDD1.n38 9.3005
R2120 VDD1.n37 VDD1.n36 9.3005
R2121 VDD1.n18 VDD1.n17 9.3005
R2122 VDD1.n31 VDD1.n30 9.3005
R2123 VDD1.n29 VDD1.n28 9.3005
R2124 VDD1.n22 VDD1.n21 9.3005
R2125 VDD1.n116 VDD1.n115 9.3005
R2126 VDD1.n85 VDD1.n84 9.3005
R2127 VDD1.n110 VDD1.n109 9.3005
R2128 VDD1.n108 VDD1.n107 9.3005
R2129 VDD1.n89 VDD1.n88 9.3005
R2130 VDD1.n102 VDD1.n101 9.3005
R2131 VDD1.n100 VDD1.n99 9.3005
R2132 VDD1.n93 VDD1.n92 9.3005
R2133 VDD1.n118 VDD1.n117 9.3005
R2134 VDD1.n81 VDD1.n80 9.3005
R2135 VDD1.n124 VDD1.n123 9.3005
R2136 VDD1.n126 VDD1.n125 9.3005
R2137 VDD1.n77 VDD1.n76 9.3005
R2138 VDD1.n132 VDD1.n131 9.3005
R2139 VDD1.n134 VDD1.n133 9.3005
R2140 VDD1.n73 VDD1.n72 9.3005
R2141 VDD1.n140 VDD1.n139 9.3005
R2142 VDD1.n55 VDD1.n8 8.92171
R2143 VDD1.n40 VDD1.n39 8.92171
R2144 VDD1.n111 VDD1.n110 8.92171
R2145 VDD1.n126 VDD1.n79 8.92171
R2146 VDD1.n70 VDD1.n0 8.2187
R2147 VDD1.n141 VDD1.n71 8.2187
R2148 VDD1.n52 VDD1.n51 8.14595
R2149 VDD1.n43 VDD1.n14 8.14595
R2150 VDD1.n114 VDD1.n85 8.14595
R2151 VDD1.n123 VDD1.n122 8.14595
R2152 VDD1.n48 VDD1.n10 7.3702
R2153 VDD1.n44 VDD1.n12 7.3702
R2154 VDD1.n115 VDD1.n83 7.3702
R2155 VDD1.n119 VDD1.n81 7.3702
R2156 VDD1.n48 VDD1.n47 6.59444
R2157 VDD1.n47 VDD1.n12 6.59444
R2158 VDD1.n118 VDD1.n83 6.59444
R2159 VDD1.n119 VDD1.n118 6.59444
R2160 VDD1.n51 VDD1.n10 5.81868
R2161 VDD1.n44 VDD1.n43 5.81868
R2162 VDD1.n115 VDD1.n114 5.81868
R2163 VDD1.n122 VDD1.n81 5.81868
R2164 VDD1.n68 VDD1.n0 5.3904
R2165 VDD1.n139 VDD1.n71 5.3904
R2166 VDD1.n52 VDD1.n8 5.04292
R2167 VDD1.n40 VDD1.n14 5.04292
R2168 VDD1.n111 VDD1.n85 5.04292
R2169 VDD1.n123 VDD1.n79 5.04292
R2170 VDD1.n94 VDD1.n92 4.38563
R2171 VDD1.n23 VDD1.n21 4.38563
R2172 VDD1.n56 VDD1.n55 4.26717
R2173 VDD1.n39 VDD1.n16 4.26717
R2174 VDD1.n110 VDD1.n87 4.26717
R2175 VDD1.n127 VDD1.n126 4.26717
R2176 VDD1.n59 VDD1.n6 3.49141
R2177 VDD1.n36 VDD1.n35 3.49141
R2178 VDD1.n107 VDD1.n106 3.49141
R2179 VDD1.n130 VDD1.n77 3.49141
R2180 VDD1.n60 VDD1.n4 2.71565
R2181 VDD1.n32 VDD1.n18 2.71565
R2182 VDD1.n103 VDD1.n89 2.71565
R2183 VDD1.n131 VDD1.n75 2.71565
R2184 VDD1.n64 VDD1.n63 1.93989
R2185 VDD1.n31 VDD1.n20 1.93989
R2186 VDD1.n102 VDD1.n91 1.93989
R2187 VDD1.n135 VDD1.n134 1.93989
R2188 VDD1.n67 VDD1.n2 1.16414
R2189 VDD1.n28 VDD1.n27 1.16414
R2190 VDD1.n99 VDD1.n98 1.16414
R2191 VDD1.n138 VDD1.n73 1.16414
R2192 VDD1.n24 VDD1.n22 0.388379
R2193 VDD1.n95 VDD1.n93 0.388379
R2194 VDD1.n69 VDD1.n1 0.155672
R2195 VDD1.n62 VDD1.n1 0.155672
R2196 VDD1.n62 VDD1.n61 0.155672
R2197 VDD1.n61 VDD1.n5 0.155672
R2198 VDD1.n54 VDD1.n5 0.155672
R2199 VDD1.n54 VDD1.n53 0.155672
R2200 VDD1.n53 VDD1.n9 0.155672
R2201 VDD1.n46 VDD1.n9 0.155672
R2202 VDD1.n46 VDD1.n45 0.155672
R2203 VDD1.n45 VDD1.n13 0.155672
R2204 VDD1.n38 VDD1.n13 0.155672
R2205 VDD1.n38 VDD1.n37 0.155672
R2206 VDD1.n37 VDD1.n17 0.155672
R2207 VDD1.n30 VDD1.n17 0.155672
R2208 VDD1.n30 VDD1.n29 0.155672
R2209 VDD1.n29 VDD1.n21 0.155672
R2210 VDD1.n100 VDD1.n92 0.155672
R2211 VDD1.n101 VDD1.n100 0.155672
R2212 VDD1.n101 VDD1.n88 0.155672
R2213 VDD1.n108 VDD1.n88 0.155672
R2214 VDD1.n109 VDD1.n108 0.155672
R2215 VDD1.n109 VDD1.n84 0.155672
R2216 VDD1.n116 VDD1.n84 0.155672
R2217 VDD1.n117 VDD1.n116 0.155672
R2218 VDD1.n117 VDD1.n80 0.155672
R2219 VDD1.n124 VDD1.n80 0.155672
R2220 VDD1.n125 VDD1.n124 0.155672
R2221 VDD1.n125 VDD1.n76 0.155672
R2222 VDD1.n132 VDD1.n76 0.155672
R2223 VDD1.n133 VDD1.n132 0.155672
R2224 VDD1.n133 VDD1.n72 0.155672
R2225 VDD1.n140 VDD1.n72 0.155672
C0 VN VTAIL 2.78084f
C1 VP VDD2 0.352063f
C2 VDD2 VDD1 0.72939f
C3 VP VDD1 3.34566f
C4 VDD2 VTAIL 5.55371f
C5 VP VTAIL 2.79512f
C6 VDD1 VTAIL 5.49993f
C7 VN VDD2 3.14447f
C8 VN VP 5.92191f
C9 VN VDD1 0.148329f
C10 VDD2 B 4.836471f
C11 VDD1 B 7.77659f
C12 VTAIL B 8.149636f
C13 VN B 11.430599f
C14 VP B 7.042014f
C15 VDD1.n0 B 0.028229f
C16 VDD1.n1 B 0.020287f
C17 VDD1.n2 B 0.010902f
C18 VDD1.n3 B 0.025767f
C19 VDD1.n4 B 0.011543f
C20 VDD1.n5 B 0.020287f
C21 VDD1.n6 B 0.010902f
C22 VDD1.n7 B 0.025767f
C23 VDD1.n8 B 0.011543f
C24 VDD1.n9 B 0.020287f
C25 VDD1.n10 B 0.010902f
C26 VDD1.n11 B 0.025767f
C27 VDD1.n12 B 0.011543f
C28 VDD1.n13 B 0.020287f
C29 VDD1.n14 B 0.010902f
C30 VDD1.n15 B 0.025767f
C31 VDD1.n16 B 0.011543f
C32 VDD1.n17 B 0.020287f
C33 VDD1.n18 B 0.010902f
C34 VDD1.n19 B 0.025767f
C35 VDD1.n20 B 0.011543f
C36 VDD1.n21 B 1.17023f
C37 VDD1.n22 B 0.010902f
C38 VDD1.t1 B 0.042375f
C39 VDD1.n23 B 0.124129f
C40 VDD1.n24 B 0.015221f
C41 VDD1.n25 B 0.019325f
C42 VDD1.n26 B 0.025767f
C43 VDD1.n27 B 0.011543f
C44 VDD1.n28 B 0.010902f
C45 VDD1.n29 B 0.020287f
C46 VDD1.n30 B 0.020287f
C47 VDD1.n31 B 0.010902f
C48 VDD1.n32 B 0.011543f
C49 VDD1.n33 B 0.025767f
C50 VDD1.n34 B 0.025767f
C51 VDD1.n35 B 0.011543f
C52 VDD1.n36 B 0.010902f
C53 VDD1.n37 B 0.020287f
C54 VDD1.n38 B 0.020287f
C55 VDD1.n39 B 0.010902f
C56 VDD1.n40 B 0.011543f
C57 VDD1.n41 B 0.025767f
C58 VDD1.n42 B 0.025767f
C59 VDD1.n43 B 0.011543f
C60 VDD1.n44 B 0.010902f
C61 VDD1.n45 B 0.020287f
C62 VDD1.n46 B 0.020287f
C63 VDD1.n47 B 0.010902f
C64 VDD1.n48 B 0.011543f
C65 VDD1.n49 B 0.025767f
C66 VDD1.n50 B 0.025767f
C67 VDD1.n51 B 0.011543f
C68 VDD1.n52 B 0.010902f
C69 VDD1.n53 B 0.020287f
C70 VDD1.n54 B 0.020287f
C71 VDD1.n55 B 0.010902f
C72 VDD1.n56 B 0.011543f
C73 VDD1.n57 B 0.025767f
C74 VDD1.n58 B 0.025767f
C75 VDD1.n59 B 0.011543f
C76 VDD1.n60 B 0.010902f
C77 VDD1.n61 B 0.020287f
C78 VDD1.n62 B 0.020287f
C79 VDD1.n63 B 0.010902f
C80 VDD1.n64 B 0.011543f
C81 VDD1.n65 B 0.025767f
C82 VDD1.n66 B 0.053221f
C83 VDD1.n67 B 0.011543f
C84 VDD1.n68 B 0.021316f
C85 VDD1.n69 B 0.052159f
C86 VDD1.n70 B 0.070964f
C87 VDD1.n71 B 0.028229f
C88 VDD1.n72 B 0.020287f
C89 VDD1.n73 B 0.010902f
C90 VDD1.n74 B 0.025767f
C91 VDD1.n75 B 0.011543f
C92 VDD1.n76 B 0.020287f
C93 VDD1.n77 B 0.010902f
C94 VDD1.n78 B 0.025767f
C95 VDD1.n79 B 0.011543f
C96 VDD1.n80 B 0.020287f
C97 VDD1.n81 B 0.010902f
C98 VDD1.n82 B 0.025767f
C99 VDD1.n83 B 0.011543f
C100 VDD1.n84 B 0.020287f
C101 VDD1.n85 B 0.010902f
C102 VDD1.n86 B 0.025767f
C103 VDD1.n87 B 0.011543f
C104 VDD1.n88 B 0.020287f
C105 VDD1.n89 B 0.010902f
C106 VDD1.n90 B 0.025767f
C107 VDD1.n91 B 0.011543f
C108 VDD1.n92 B 1.17023f
C109 VDD1.n93 B 0.010902f
C110 VDD1.t0 B 0.042375f
C111 VDD1.n94 B 0.124129f
C112 VDD1.n95 B 0.015221f
C113 VDD1.n96 B 0.019325f
C114 VDD1.n97 B 0.025767f
C115 VDD1.n98 B 0.011543f
C116 VDD1.n99 B 0.010902f
C117 VDD1.n100 B 0.020287f
C118 VDD1.n101 B 0.020287f
C119 VDD1.n102 B 0.010902f
C120 VDD1.n103 B 0.011543f
C121 VDD1.n104 B 0.025767f
C122 VDD1.n105 B 0.025767f
C123 VDD1.n106 B 0.011543f
C124 VDD1.n107 B 0.010902f
C125 VDD1.n108 B 0.020287f
C126 VDD1.n109 B 0.020287f
C127 VDD1.n110 B 0.010902f
C128 VDD1.n111 B 0.011543f
C129 VDD1.n112 B 0.025767f
C130 VDD1.n113 B 0.025767f
C131 VDD1.n114 B 0.011543f
C132 VDD1.n115 B 0.010902f
C133 VDD1.n116 B 0.020287f
C134 VDD1.n117 B 0.020287f
C135 VDD1.n118 B 0.010902f
C136 VDD1.n119 B 0.011543f
C137 VDD1.n120 B 0.025767f
C138 VDD1.n121 B 0.025767f
C139 VDD1.n122 B 0.011543f
C140 VDD1.n123 B 0.010902f
C141 VDD1.n124 B 0.020287f
C142 VDD1.n125 B 0.020287f
C143 VDD1.n126 B 0.010902f
C144 VDD1.n127 B 0.011543f
C145 VDD1.n128 B 0.025767f
C146 VDD1.n129 B 0.025767f
C147 VDD1.n130 B 0.011543f
C148 VDD1.n131 B 0.010902f
C149 VDD1.n132 B 0.020287f
C150 VDD1.n133 B 0.020287f
C151 VDD1.n134 B 0.010902f
C152 VDD1.n135 B 0.011543f
C153 VDD1.n136 B 0.025767f
C154 VDD1.n137 B 0.053221f
C155 VDD1.n138 B 0.011543f
C156 VDD1.n139 B 0.021316f
C157 VDD1.n140 B 0.052159f
C158 VDD1.n141 B 0.705708f
C159 VP.t1 B 3.49806f
C160 VP.t0 B 4.10097f
C161 VP.n0 B 4.31583f
C162 VDD2.n0 B 0.028148f
C163 VDD2.n1 B 0.020229f
C164 VDD2.n2 B 0.01087f
C165 VDD2.n3 B 0.025693f
C166 VDD2.n4 B 0.01151f
C167 VDD2.n5 B 0.020229f
C168 VDD2.n6 B 0.01087f
C169 VDD2.n7 B 0.025693f
C170 VDD2.n8 B 0.01151f
C171 VDD2.n9 B 0.020229f
C172 VDD2.n10 B 0.01087f
C173 VDD2.n11 B 0.025693f
C174 VDD2.n12 B 0.01151f
C175 VDD2.n13 B 0.020229f
C176 VDD2.n14 B 0.01087f
C177 VDD2.n15 B 0.025693f
C178 VDD2.n16 B 0.01151f
C179 VDD2.n17 B 0.020229f
C180 VDD2.n18 B 0.01087f
C181 VDD2.n19 B 0.025693f
C182 VDD2.n20 B 0.01151f
C183 VDD2.n21 B 1.16687f
C184 VDD2.n22 B 0.01087f
C185 VDD2.t1 B 0.042253f
C186 VDD2.n23 B 0.123772f
C187 VDD2.n24 B 0.015178f
C188 VDD2.n25 B 0.01927f
C189 VDD2.n26 B 0.025693f
C190 VDD2.n27 B 0.01151f
C191 VDD2.n28 B 0.01087f
C192 VDD2.n29 B 0.020229f
C193 VDD2.n30 B 0.020229f
C194 VDD2.n31 B 0.01087f
C195 VDD2.n32 B 0.01151f
C196 VDD2.n33 B 0.025693f
C197 VDD2.n34 B 0.025693f
C198 VDD2.n35 B 0.01151f
C199 VDD2.n36 B 0.01087f
C200 VDD2.n37 B 0.020229f
C201 VDD2.n38 B 0.020229f
C202 VDD2.n39 B 0.01087f
C203 VDD2.n40 B 0.01151f
C204 VDD2.n41 B 0.025693f
C205 VDD2.n42 B 0.025693f
C206 VDD2.n43 B 0.01151f
C207 VDD2.n44 B 0.01087f
C208 VDD2.n45 B 0.020229f
C209 VDD2.n46 B 0.020229f
C210 VDD2.n47 B 0.01087f
C211 VDD2.n48 B 0.01151f
C212 VDD2.n49 B 0.025693f
C213 VDD2.n50 B 0.025693f
C214 VDD2.n51 B 0.01151f
C215 VDD2.n52 B 0.01087f
C216 VDD2.n53 B 0.020229f
C217 VDD2.n54 B 0.020229f
C218 VDD2.n55 B 0.01087f
C219 VDD2.n56 B 0.01151f
C220 VDD2.n57 B 0.025693f
C221 VDD2.n58 B 0.025693f
C222 VDD2.n59 B 0.01151f
C223 VDD2.n60 B 0.01087f
C224 VDD2.n61 B 0.020229f
C225 VDD2.n62 B 0.020229f
C226 VDD2.n63 B 0.01087f
C227 VDD2.n64 B 0.01151f
C228 VDD2.n65 B 0.025693f
C229 VDD2.n66 B 0.053069f
C230 VDD2.n67 B 0.01151f
C231 VDD2.n68 B 0.021255f
C232 VDD2.n69 B 0.052009f
C233 VDD2.n70 B 0.661092f
C234 VDD2.n71 B 0.028148f
C235 VDD2.n72 B 0.020229f
C236 VDD2.n73 B 0.01087f
C237 VDD2.n74 B 0.025693f
C238 VDD2.n75 B 0.01151f
C239 VDD2.n76 B 0.020229f
C240 VDD2.n77 B 0.01087f
C241 VDD2.n78 B 0.025693f
C242 VDD2.n79 B 0.01151f
C243 VDD2.n80 B 0.020229f
C244 VDD2.n81 B 0.01087f
C245 VDD2.n82 B 0.025693f
C246 VDD2.n83 B 0.01151f
C247 VDD2.n84 B 0.020229f
C248 VDD2.n85 B 0.01087f
C249 VDD2.n86 B 0.025693f
C250 VDD2.n87 B 0.01151f
C251 VDD2.n88 B 0.020229f
C252 VDD2.n89 B 0.01087f
C253 VDD2.n90 B 0.025693f
C254 VDD2.n91 B 0.01151f
C255 VDD2.n92 B 1.16687f
C256 VDD2.n93 B 0.01087f
C257 VDD2.t0 B 0.042253f
C258 VDD2.n94 B 0.123772f
C259 VDD2.n95 B 0.015178f
C260 VDD2.n96 B 0.01927f
C261 VDD2.n97 B 0.025693f
C262 VDD2.n98 B 0.01151f
C263 VDD2.n99 B 0.01087f
C264 VDD2.n100 B 0.020229f
C265 VDD2.n101 B 0.020229f
C266 VDD2.n102 B 0.01087f
C267 VDD2.n103 B 0.01151f
C268 VDD2.n104 B 0.025693f
C269 VDD2.n105 B 0.025693f
C270 VDD2.n106 B 0.01151f
C271 VDD2.n107 B 0.01087f
C272 VDD2.n108 B 0.020229f
C273 VDD2.n109 B 0.020229f
C274 VDD2.n110 B 0.01087f
C275 VDD2.n111 B 0.01151f
C276 VDD2.n112 B 0.025693f
C277 VDD2.n113 B 0.025693f
C278 VDD2.n114 B 0.01151f
C279 VDD2.n115 B 0.01087f
C280 VDD2.n116 B 0.020229f
C281 VDD2.n117 B 0.020229f
C282 VDD2.n118 B 0.01087f
C283 VDD2.n119 B 0.01151f
C284 VDD2.n120 B 0.025693f
C285 VDD2.n121 B 0.025693f
C286 VDD2.n122 B 0.01151f
C287 VDD2.n123 B 0.01087f
C288 VDD2.n124 B 0.020229f
C289 VDD2.n125 B 0.020229f
C290 VDD2.n126 B 0.01087f
C291 VDD2.n127 B 0.01151f
C292 VDD2.n128 B 0.025693f
C293 VDD2.n129 B 0.025693f
C294 VDD2.n130 B 0.01151f
C295 VDD2.n131 B 0.01087f
C296 VDD2.n132 B 0.020229f
C297 VDD2.n133 B 0.020229f
C298 VDD2.n134 B 0.01087f
C299 VDD2.n135 B 0.01151f
C300 VDD2.n136 B 0.025693f
C301 VDD2.n137 B 0.053069f
C302 VDD2.n138 B 0.01151f
C303 VDD2.n139 B 0.021255f
C304 VDD2.n140 B 0.052009f
C305 VDD2.n141 B 0.069385f
C306 VDD2.n142 B 2.68526f
C307 VTAIL.n0 B 0.028789f
C308 VTAIL.n1 B 0.020689f
C309 VTAIL.n2 B 0.011118f
C310 VTAIL.n3 B 0.026278f
C311 VTAIL.n4 B 0.011772f
C312 VTAIL.n5 B 0.020689f
C313 VTAIL.n6 B 0.011118f
C314 VTAIL.n7 B 0.026278f
C315 VTAIL.n8 B 0.011772f
C316 VTAIL.n9 B 0.020689f
C317 VTAIL.n10 B 0.011118f
C318 VTAIL.n11 B 0.026278f
C319 VTAIL.n12 B 0.011772f
C320 VTAIL.n13 B 0.020689f
C321 VTAIL.n14 B 0.011118f
C322 VTAIL.n15 B 0.026278f
C323 VTAIL.n16 B 0.011772f
C324 VTAIL.n17 B 0.020689f
C325 VTAIL.n18 B 0.011118f
C326 VTAIL.n19 B 0.026278f
C327 VTAIL.n20 B 0.011772f
C328 VTAIL.n21 B 1.19342f
C329 VTAIL.n22 B 0.011118f
C330 VTAIL.t1 B 0.043215f
C331 VTAIL.n23 B 0.126589f
C332 VTAIL.n24 B 0.015523f
C333 VTAIL.n25 B 0.019708f
C334 VTAIL.n26 B 0.026278f
C335 VTAIL.n27 B 0.011772f
C336 VTAIL.n28 B 0.011118f
C337 VTAIL.n29 B 0.020689f
C338 VTAIL.n30 B 0.020689f
C339 VTAIL.n31 B 0.011118f
C340 VTAIL.n32 B 0.011772f
C341 VTAIL.n33 B 0.026278f
C342 VTAIL.n34 B 0.026278f
C343 VTAIL.n35 B 0.011772f
C344 VTAIL.n36 B 0.011118f
C345 VTAIL.n37 B 0.020689f
C346 VTAIL.n38 B 0.020689f
C347 VTAIL.n39 B 0.011118f
C348 VTAIL.n40 B 0.011772f
C349 VTAIL.n41 B 0.026278f
C350 VTAIL.n42 B 0.026278f
C351 VTAIL.n43 B 0.011772f
C352 VTAIL.n44 B 0.011118f
C353 VTAIL.n45 B 0.020689f
C354 VTAIL.n46 B 0.020689f
C355 VTAIL.n47 B 0.011118f
C356 VTAIL.n48 B 0.011772f
C357 VTAIL.n49 B 0.026278f
C358 VTAIL.n50 B 0.026278f
C359 VTAIL.n51 B 0.011772f
C360 VTAIL.n52 B 0.011118f
C361 VTAIL.n53 B 0.020689f
C362 VTAIL.n54 B 0.020689f
C363 VTAIL.n55 B 0.011118f
C364 VTAIL.n56 B 0.011772f
C365 VTAIL.n57 B 0.026278f
C366 VTAIL.n58 B 0.026278f
C367 VTAIL.n59 B 0.011772f
C368 VTAIL.n60 B 0.011118f
C369 VTAIL.n61 B 0.020689f
C370 VTAIL.n62 B 0.020689f
C371 VTAIL.n63 B 0.011118f
C372 VTAIL.n64 B 0.011772f
C373 VTAIL.n65 B 0.026278f
C374 VTAIL.n66 B 0.054276f
C375 VTAIL.n67 B 0.011772f
C376 VTAIL.n68 B 0.021738f
C377 VTAIL.n69 B 0.053193f
C378 VTAIL.n70 B 0.056716f
C379 VTAIL.n71 B 1.54354f
C380 VTAIL.n72 B 0.028789f
C381 VTAIL.n73 B 0.020689f
C382 VTAIL.n74 B 0.011118f
C383 VTAIL.n75 B 0.026278f
C384 VTAIL.n76 B 0.011772f
C385 VTAIL.n77 B 0.020689f
C386 VTAIL.n78 B 0.011118f
C387 VTAIL.n79 B 0.026278f
C388 VTAIL.n80 B 0.011772f
C389 VTAIL.n81 B 0.020689f
C390 VTAIL.n82 B 0.011118f
C391 VTAIL.n83 B 0.026278f
C392 VTAIL.n84 B 0.011772f
C393 VTAIL.n85 B 0.020689f
C394 VTAIL.n86 B 0.011118f
C395 VTAIL.n87 B 0.026278f
C396 VTAIL.n88 B 0.011772f
C397 VTAIL.n89 B 0.020689f
C398 VTAIL.n90 B 0.011118f
C399 VTAIL.n91 B 0.026278f
C400 VTAIL.n92 B 0.011772f
C401 VTAIL.n93 B 1.19342f
C402 VTAIL.n94 B 0.011118f
C403 VTAIL.t2 B 0.043215f
C404 VTAIL.n95 B 0.126589f
C405 VTAIL.n96 B 0.015523f
C406 VTAIL.n97 B 0.019708f
C407 VTAIL.n98 B 0.026278f
C408 VTAIL.n99 B 0.011772f
C409 VTAIL.n100 B 0.011118f
C410 VTAIL.n101 B 0.020689f
C411 VTAIL.n102 B 0.020689f
C412 VTAIL.n103 B 0.011118f
C413 VTAIL.n104 B 0.011772f
C414 VTAIL.n105 B 0.026278f
C415 VTAIL.n106 B 0.026278f
C416 VTAIL.n107 B 0.011772f
C417 VTAIL.n108 B 0.011118f
C418 VTAIL.n109 B 0.020689f
C419 VTAIL.n110 B 0.020689f
C420 VTAIL.n111 B 0.011118f
C421 VTAIL.n112 B 0.011772f
C422 VTAIL.n113 B 0.026278f
C423 VTAIL.n114 B 0.026278f
C424 VTAIL.n115 B 0.011772f
C425 VTAIL.n116 B 0.011118f
C426 VTAIL.n117 B 0.020689f
C427 VTAIL.n118 B 0.020689f
C428 VTAIL.n119 B 0.011118f
C429 VTAIL.n120 B 0.011772f
C430 VTAIL.n121 B 0.026278f
C431 VTAIL.n122 B 0.026278f
C432 VTAIL.n123 B 0.011772f
C433 VTAIL.n124 B 0.011118f
C434 VTAIL.n125 B 0.020689f
C435 VTAIL.n126 B 0.020689f
C436 VTAIL.n127 B 0.011118f
C437 VTAIL.n128 B 0.011772f
C438 VTAIL.n129 B 0.026278f
C439 VTAIL.n130 B 0.026278f
C440 VTAIL.n131 B 0.011772f
C441 VTAIL.n132 B 0.011118f
C442 VTAIL.n133 B 0.020689f
C443 VTAIL.n134 B 0.020689f
C444 VTAIL.n135 B 0.011118f
C445 VTAIL.n136 B 0.011772f
C446 VTAIL.n137 B 0.026278f
C447 VTAIL.n138 B 0.054276f
C448 VTAIL.n139 B 0.011772f
C449 VTAIL.n140 B 0.021738f
C450 VTAIL.n141 B 0.053193f
C451 VTAIL.n142 B 0.056716f
C452 VTAIL.n143 B 1.58823f
C453 VTAIL.n144 B 0.028789f
C454 VTAIL.n145 B 0.020689f
C455 VTAIL.n146 B 0.011118f
C456 VTAIL.n147 B 0.026278f
C457 VTAIL.n148 B 0.011772f
C458 VTAIL.n149 B 0.020689f
C459 VTAIL.n150 B 0.011118f
C460 VTAIL.n151 B 0.026278f
C461 VTAIL.n152 B 0.011772f
C462 VTAIL.n153 B 0.020689f
C463 VTAIL.n154 B 0.011118f
C464 VTAIL.n155 B 0.026278f
C465 VTAIL.n156 B 0.011772f
C466 VTAIL.n157 B 0.020689f
C467 VTAIL.n158 B 0.011118f
C468 VTAIL.n159 B 0.026278f
C469 VTAIL.n160 B 0.011772f
C470 VTAIL.n161 B 0.020689f
C471 VTAIL.n162 B 0.011118f
C472 VTAIL.n163 B 0.026278f
C473 VTAIL.n164 B 0.011772f
C474 VTAIL.n165 B 1.19342f
C475 VTAIL.n166 B 0.011118f
C476 VTAIL.t0 B 0.043215f
C477 VTAIL.n167 B 0.126589f
C478 VTAIL.n168 B 0.015523f
C479 VTAIL.n169 B 0.019708f
C480 VTAIL.n170 B 0.026278f
C481 VTAIL.n171 B 0.011772f
C482 VTAIL.n172 B 0.011118f
C483 VTAIL.n173 B 0.020689f
C484 VTAIL.n174 B 0.020689f
C485 VTAIL.n175 B 0.011118f
C486 VTAIL.n176 B 0.011772f
C487 VTAIL.n177 B 0.026278f
C488 VTAIL.n178 B 0.026278f
C489 VTAIL.n179 B 0.011772f
C490 VTAIL.n180 B 0.011118f
C491 VTAIL.n181 B 0.020689f
C492 VTAIL.n182 B 0.020689f
C493 VTAIL.n183 B 0.011118f
C494 VTAIL.n184 B 0.011772f
C495 VTAIL.n185 B 0.026278f
C496 VTAIL.n186 B 0.026278f
C497 VTAIL.n187 B 0.011772f
C498 VTAIL.n188 B 0.011118f
C499 VTAIL.n189 B 0.020689f
C500 VTAIL.n190 B 0.020689f
C501 VTAIL.n191 B 0.011118f
C502 VTAIL.n192 B 0.011772f
C503 VTAIL.n193 B 0.026278f
C504 VTAIL.n194 B 0.026278f
C505 VTAIL.n195 B 0.011772f
C506 VTAIL.n196 B 0.011118f
C507 VTAIL.n197 B 0.020689f
C508 VTAIL.n198 B 0.020689f
C509 VTAIL.n199 B 0.011118f
C510 VTAIL.n200 B 0.011772f
C511 VTAIL.n201 B 0.026278f
C512 VTAIL.n202 B 0.026278f
C513 VTAIL.n203 B 0.011772f
C514 VTAIL.n204 B 0.011118f
C515 VTAIL.n205 B 0.020689f
C516 VTAIL.n206 B 0.020689f
C517 VTAIL.n207 B 0.011118f
C518 VTAIL.n208 B 0.011772f
C519 VTAIL.n209 B 0.026278f
C520 VTAIL.n210 B 0.054276f
C521 VTAIL.n211 B 0.011772f
C522 VTAIL.n212 B 0.021738f
C523 VTAIL.n213 B 0.053193f
C524 VTAIL.n214 B 0.056716f
C525 VTAIL.n215 B 1.39397f
C526 VTAIL.n216 B 0.028789f
C527 VTAIL.n217 B 0.020689f
C528 VTAIL.n218 B 0.011118f
C529 VTAIL.n219 B 0.026278f
C530 VTAIL.n220 B 0.011772f
C531 VTAIL.n221 B 0.020689f
C532 VTAIL.n222 B 0.011118f
C533 VTAIL.n223 B 0.026278f
C534 VTAIL.n224 B 0.011772f
C535 VTAIL.n225 B 0.020689f
C536 VTAIL.n226 B 0.011118f
C537 VTAIL.n227 B 0.026278f
C538 VTAIL.n228 B 0.011772f
C539 VTAIL.n229 B 0.020689f
C540 VTAIL.n230 B 0.011118f
C541 VTAIL.n231 B 0.026278f
C542 VTAIL.n232 B 0.011772f
C543 VTAIL.n233 B 0.020689f
C544 VTAIL.n234 B 0.011118f
C545 VTAIL.n235 B 0.026278f
C546 VTAIL.n236 B 0.011772f
C547 VTAIL.n237 B 1.19342f
C548 VTAIL.n238 B 0.011118f
C549 VTAIL.t3 B 0.043215f
C550 VTAIL.n239 B 0.126589f
C551 VTAIL.n240 B 0.015523f
C552 VTAIL.n241 B 0.019708f
C553 VTAIL.n242 B 0.026278f
C554 VTAIL.n243 B 0.011772f
C555 VTAIL.n244 B 0.011118f
C556 VTAIL.n245 B 0.020689f
C557 VTAIL.n246 B 0.020689f
C558 VTAIL.n247 B 0.011118f
C559 VTAIL.n248 B 0.011772f
C560 VTAIL.n249 B 0.026278f
C561 VTAIL.n250 B 0.026278f
C562 VTAIL.n251 B 0.011772f
C563 VTAIL.n252 B 0.011118f
C564 VTAIL.n253 B 0.020689f
C565 VTAIL.n254 B 0.020689f
C566 VTAIL.n255 B 0.011118f
C567 VTAIL.n256 B 0.011772f
C568 VTAIL.n257 B 0.026278f
C569 VTAIL.n258 B 0.026278f
C570 VTAIL.n259 B 0.011772f
C571 VTAIL.n260 B 0.011118f
C572 VTAIL.n261 B 0.020689f
C573 VTAIL.n262 B 0.020689f
C574 VTAIL.n263 B 0.011118f
C575 VTAIL.n264 B 0.011772f
C576 VTAIL.n265 B 0.026278f
C577 VTAIL.n266 B 0.026278f
C578 VTAIL.n267 B 0.011772f
C579 VTAIL.n268 B 0.011118f
C580 VTAIL.n269 B 0.020689f
C581 VTAIL.n270 B 0.020689f
C582 VTAIL.n271 B 0.011118f
C583 VTAIL.n272 B 0.011772f
C584 VTAIL.n273 B 0.026278f
C585 VTAIL.n274 B 0.026278f
C586 VTAIL.n275 B 0.011772f
C587 VTAIL.n276 B 0.011118f
C588 VTAIL.n277 B 0.020689f
C589 VTAIL.n278 B 0.020689f
C590 VTAIL.n279 B 0.011118f
C591 VTAIL.n280 B 0.011772f
C592 VTAIL.n281 B 0.026278f
C593 VTAIL.n282 B 0.054276f
C594 VTAIL.n283 B 0.011772f
C595 VTAIL.n284 B 0.021738f
C596 VTAIL.n285 B 0.053193f
C597 VTAIL.n286 B 0.056716f
C598 VTAIL.n287 B 1.31021f
C599 VN.t0 B 3.43163f
C600 VN.t1 B 4.02099f
.ends

