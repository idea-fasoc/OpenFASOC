* NGSPICE file created from diff_pair_sample_1423.ext - technology: sky130A

.subckt diff_pair_sample_1423 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t9 VN.t0 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=1.2441 pd=7.87 as=1.2441 ps=7.87 w=7.54 l=1.63
X1 VDD2.t4 VN.t1 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=2.9406 pd=15.86 as=1.2441 ps=7.87 w=7.54 l=1.63
X2 VDD1.t5 VP.t0 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=2.9406 pd=15.86 as=1.2441 ps=7.87 w=7.54 l=1.63
X3 VDD1.t4 VP.t1 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=1.2441 pd=7.87 as=2.9406 ps=15.86 w=7.54 l=1.63
X4 VDD2.t2 VN.t2 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2441 pd=7.87 as=2.9406 ps=15.86 w=7.54 l=1.63
X5 VTAIL.t6 VN.t3 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2441 pd=7.87 as=1.2441 ps=7.87 w=7.54 l=1.63
X6 VDD2.t0 VN.t4 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9406 pd=15.86 as=1.2441 ps=7.87 w=7.54 l=1.63
X7 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=2.9406 pd=15.86 as=0 ps=0 w=7.54 l=1.63
X8 VTAIL.t3 VP.t2 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2441 pd=7.87 as=1.2441 ps=7.87 w=7.54 l=1.63
X9 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=2.9406 pd=15.86 as=0 ps=0 w=7.54 l=1.63
X10 VDD2.t5 VN.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.2441 pd=7.87 as=2.9406 ps=15.86 w=7.54 l=1.63
X11 VTAIL.t2 VP.t3 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.2441 pd=7.87 as=1.2441 ps=7.87 w=7.54 l=1.63
X12 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.9406 pd=15.86 as=0 ps=0 w=7.54 l=1.63
X13 VDD1.t1 VP.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2441 pd=7.87 as=2.9406 ps=15.86 w=7.54 l=1.63
X14 VDD1.t0 VP.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9406 pd=15.86 as=1.2441 ps=7.87 w=7.54 l=1.63
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.9406 pd=15.86 as=0 ps=0 w=7.54 l=1.63
R0 VN.n11 VN.n10 175.564
R1 VN.n23 VN.n22 175.564
R2 VN.n21 VN.n12 161.3
R3 VN.n20 VN.n19 161.3
R4 VN.n18 VN.n13 161.3
R5 VN.n17 VN.n16 161.3
R6 VN.n9 VN.n0 161.3
R7 VN.n8 VN.n7 161.3
R8 VN.n6 VN.n1 161.3
R9 VN.n5 VN.n4 161.3
R10 VN.n2 VN.t1 145.44
R11 VN.n14 VN.t5 145.44
R12 VN.n3 VN.t3 111.481
R13 VN.n10 VN.t2 111.481
R14 VN.n15 VN.t0 111.481
R15 VN.n22 VN.t4 111.481
R16 VN.n8 VN.n1 56.5617
R17 VN.n20 VN.n13 56.5617
R18 VN.n3 VN.n2 54.3154
R19 VN.n15 VN.n14 54.3154
R20 VN VN.n23 41.8357
R21 VN.n4 VN.n1 24.5923
R22 VN.n9 VN.n8 24.5923
R23 VN.n16 VN.n13 24.5923
R24 VN.n21 VN.n20 24.5923
R25 VN.n17 VN.n14 17.7323
R26 VN.n5 VN.n2 17.7323
R27 VN.n4 VN.n3 12.2964
R28 VN.n16 VN.n15 12.2964
R29 VN.n10 VN.n9 10.3291
R30 VN.n22 VN.n21 10.3291
R31 VN.n23 VN.n12 0.189894
R32 VN.n19 VN.n12 0.189894
R33 VN.n19 VN.n18 0.189894
R34 VN.n18 VN.n17 0.189894
R35 VN.n6 VN.n5 0.189894
R36 VN.n7 VN.n6 0.189894
R37 VN.n7 VN.n0 0.189894
R38 VN.n11 VN.n0 0.189894
R39 VN VN.n11 0.0516364
R40 VDD2.n1 VDD2.t4 70.0684
R41 VDD2.n2 VDD2.t0 68.8567
R42 VDD2.n1 VDD2.n0 66.5975
R43 VDD2 VDD2.n3 66.5947
R44 VDD2.n2 VDD2.n1 35.7067
R45 VDD2.n3 VDD2.t3 2.62649
R46 VDD2.n3 VDD2.t5 2.62649
R47 VDD2.n0 VDD2.t1 2.62649
R48 VDD2.n0 VDD2.t2 2.62649
R49 VDD2 VDD2.n2 1.32593
R50 VTAIL.n7 VTAIL.t4 52.1779
R51 VTAIL.n11 VTAIL.t7 52.1777
R52 VTAIL.n2 VTAIL.t10 52.1777
R53 VTAIL.n10 VTAIL.t0 52.1777
R54 VTAIL.n9 VTAIL.n8 49.5519
R55 VTAIL.n6 VTAIL.n5 49.5519
R56 VTAIL.n1 VTAIL.n0 49.5517
R57 VTAIL.n4 VTAIL.n3 49.5517
R58 VTAIL.n6 VTAIL.n4 22.2462
R59 VTAIL.n11 VTAIL.n10 20.5565
R60 VTAIL.n0 VTAIL.t8 2.62649
R61 VTAIL.n0 VTAIL.t6 2.62649
R62 VTAIL.n3 VTAIL.t1 2.62649
R63 VTAIL.n3 VTAIL.t2 2.62649
R64 VTAIL.n8 VTAIL.t11 2.62649
R65 VTAIL.n8 VTAIL.t3 2.62649
R66 VTAIL.n5 VTAIL.t5 2.62649
R67 VTAIL.n5 VTAIL.t9 2.62649
R68 VTAIL.n7 VTAIL.n6 1.69016
R69 VTAIL.n10 VTAIL.n9 1.69016
R70 VTAIL.n4 VTAIL.n2 1.69016
R71 VTAIL.n9 VTAIL.n7 1.31516
R72 VTAIL.n2 VTAIL.n1 1.31516
R73 VTAIL VTAIL.n11 1.20955
R74 VTAIL VTAIL.n1 0.481103
R75 B.n594 B.n593 585
R76 B.n595 B.n594 585
R77 B.n227 B.n93 585
R78 B.n226 B.n225 585
R79 B.n224 B.n223 585
R80 B.n222 B.n221 585
R81 B.n220 B.n219 585
R82 B.n218 B.n217 585
R83 B.n216 B.n215 585
R84 B.n214 B.n213 585
R85 B.n212 B.n211 585
R86 B.n210 B.n209 585
R87 B.n208 B.n207 585
R88 B.n206 B.n205 585
R89 B.n204 B.n203 585
R90 B.n202 B.n201 585
R91 B.n200 B.n199 585
R92 B.n198 B.n197 585
R93 B.n196 B.n195 585
R94 B.n194 B.n193 585
R95 B.n192 B.n191 585
R96 B.n190 B.n189 585
R97 B.n188 B.n187 585
R98 B.n186 B.n185 585
R99 B.n184 B.n183 585
R100 B.n182 B.n181 585
R101 B.n180 B.n179 585
R102 B.n178 B.n177 585
R103 B.n176 B.n175 585
R104 B.n174 B.n173 585
R105 B.n172 B.n171 585
R106 B.n170 B.n169 585
R107 B.n168 B.n167 585
R108 B.n166 B.n165 585
R109 B.n164 B.n163 585
R110 B.n162 B.n161 585
R111 B.n160 B.n159 585
R112 B.n158 B.n157 585
R113 B.n156 B.n155 585
R114 B.n153 B.n152 585
R115 B.n151 B.n150 585
R116 B.n149 B.n148 585
R117 B.n147 B.n146 585
R118 B.n145 B.n144 585
R119 B.n143 B.n142 585
R120 B.n141 B.n140 585
R121 B.n139 B.n138 585
R122 B.n137 B.n136 585
R123 B.n135 B.n134 585
R124 B.n133 B.n132 585
R125 B.n131 B.n130 585
R126 B.n129 B.n128 585
R127 B.n127 B.n126 585
R128 B.n125 B.n124 585
R129 B.n123 B.n122 585
R130 B.n121 B.n120 585
R131 B.n119 B.n118 585
R132 B.n117 B.n116 585
R133 B.n115 B.n114 585
R134 B.n113 B.n112 585
R135 B.n111 B.n110 585
R136 B.n109 B.n108 585
R137 B.n107 B.n106 585
R138 B.n105 B.n104 585
R139 B.n103 B.n102 585
R140 B.n101 B.n100 585
R141 B.n60 B.n59 585
R142 B.n598 B.n597 585
R143 B.n592 B.n94 585
R144 B.n94 B.n57 585
R145 B.n591 B.n56 585
R146 B.n602 B.n56 585
R147 B.n590 B.n55 585
R148 B.n603 B.n55 585
R149 B.n589 B.n54 585
R150 B.n604 B.n54 585
R151 B.n588 B.n587 585
R152 B.n587 B.n50 585
R153 B.n586 B.n49 585
R154 B.n610 B.n49 585
R155 B.n585 B.n48 585
R156 B.n611 B.n48 585
R157 B.n584 B.n47 585
R158 B.n612 B.n47 585
R159 B.n583 B.n582 585
R160 B.n582 B.n43 585
R161 B.n581 B.n42 585
R162 B.n618 B.n42 585
R163 B.n580 B.n41 585
R164 B.n619 B.n41 585
R165 B.n579 B.n40 585
R166 B.n620 B.n40 585
R167 B.n578 B.n577 585
R168 B.n577 B.n36 585
R169 B.n576 B.n35 585
R170 B.n626 B.n35 585
R171 B.n575 B.n34 585
R172 B.n627 B.n34 585
R173 B.n574 B.n33 585
R174 B.n628 B.n33 585
R175 B.n573 B.n572 585
R176 B.n572 B.n29 585
R177 B.n571 B.n28 585
R178 B.n634 B.n28 585
R179 B.n570 B.n27 585
R180 B.n635 B.n27 585
R181 B.n569 B.n26 585
R182 B.n636 B.n26 585
R183 B.n568 B.n567 585
R184 B.n567 B.n25 585
R185 B.n566 B.n21 585
R186 B.n642 B.n21 585
R187 B.n565 B.n20 585
R188 B.n643 B.n20 585
R189 B.n564 B.n19 585
R190 B.n644 B.n19 585
R191 B.n563 B.n562 585
R192 B.n562 B.n15 585
R193 B.n561 B.n14 585
R194 B.n650 B.n14 585
R195 B.n560 B.n13 585
R196 B.n651 B.n13 585
R197 B.n559 B.n12 585
R198 B.n652 B.n12 585
R199 B.n558 B.n557 585
R200 B.n557 B.n8 585
R201 B.n556 B.n7 585
R202 B.n658 B.n7 585
R203 B.n555 B.n6 585
R204 B.n659 B.n6 585
R205 B.n554 B.n5 585
R206 B.n660 B.n5 585
R207 B.n553 B.n552 585
R208 B.n552 B.n4 585
R209 B.n551 B.n228 585
R210 B.n551 B.n550 585
R211 B.n541 B.n229 585
R212 B.n230 B.n229 585
R213 B.n543 B.n542 585
R214 B.n544 B.n543 585
R215 B.n540 B.n234 585
R216 B.n238 B.n234 585
R217 B.n539 B.n538 585
R218 B.n538 B.n537 585
R219 B.n236 B.n235 585
R220 B.n237 B.n236 585
R221 B.n530 B.n529 585
R222 B.n531 B.n530 585
R223 B.n528 B.n243 585
R224 B.n243 B.n242 585
R225 B.n527 B.n526 585
R226 B.n526 B.n525 585
R227 B.n245 B.n244 585
R228 B.n518 B.n245 585
R229 B.n517 B.n516 585
R230 B.n519 B.n517 585
R231 B.n515 B.n250 585
R232 B.n250 B.n249 585
R233 B.n514 B.n513 585
R234 B.n513 B.n512 585
R235 B.n252 B.n251 585
R236 B.n253 B.n252 585
R237 B.n505 B.n504 585
R238 B.n506 B.n505 585
R239 B.n503 B.n257 585
R240 B.n261 B.n257 585
R241 B.n502 B.n501 585
R242 B.n501 B.n500 585
R243 B.n259 B.n258 585
R244 B.n260 B.n259 585
R245 B.n493 B.n492 585
R246 B.n494 B.n493 585
R247 B.n491 B.n266 585
R248 B.n266 B.n265 585
R249 B.n490 B.n489 585
R250 B.n489 B.n488 585
R251 B.n268 B.n267 585
R252 B.n269 B.n268 585
R253 B.n481 B.n480 585
R254 B.n482 B.n481 585
R255 B.n479 B.n273 585
R256 B.n277 B.n273 585
R257 B.n478 B.n477 585
R258 B.n477 B.n476 585
R259 B.n275 B.n274 585
R260 B.n276 B.n275 585
R261 B.n469 B.n468 585
R262 B.n470 B.n469 585
R263 B.n467 B.n282 585
R264 B.n282 B.n281 585
R265 B.n466 B.n465 585
R266 B.n465 B.n464 585
R267 B.n284 B.n283 585
R268 B.n285 B.n284 585
R269 B.n460 B.n459 585
R270 B.n288 B.n287 585
R271 B.n456 B.n455 585
R272 B.n457 B.n456 585
R273 B.n454 B.n321 585
R274 B.n453 B.n452 585
R275 B.n451 B.n450 585
R276 B.n449 B.n448 585
R277 B.n447 B.n446 585
R278 B.n445 B.n444 585
R279 B.n443 B.n442 585
R280 B.n441 B.n440 585
R281 B.n439 B.n438 585
R282 B.n437 B.n436 585
R283 B.n435 B.n434 585
R284 B.n433 B.n432 585
R285 B.n431 B.n430 585
R286 B.n429 B.n428 585
R287 B.n427 B.n426 585
R288 B.n425 B.n424 585
R289 B.n423 B.n422 585
R290 B.n421 B.n420 585
R291 B.n419 B.n418 585
R292 B.n417 B.n416 585
R293 B.n415 B.n414 585
R294 B.n413 B.n412 585
R295 B.n411 B.n410 585
R296 B.n409 B.n408 585
R297 B.n407 B.n406 585
R298 B.n405 B.n404 585
R299 B.n403 B.n402 585
R300 B.n401 B.n400 585
R301 B.n399 B.n398 585
R302 B.n397 B.n396 585
R303 B.n395 B.n394 585
R304 B.n393 B.n392 585
R305 B.n391 B.n390 585
R306 B.n389 B.n388 585
R307 B.n387 B.n386 585
R308 B.n384 B.n383 585
R309 B.n382 B.n381 585
R310 B.n380 B.n379 585
R311 B.n378 B.n377 585
R312 B.n376 B.n375 585
R313 B.n374 B.n373 585
R314 B.n372 B.n371 585
R315 B.n370 B.n369 585
R316 B.n368 B.n367 585
R317 B.n366 B.n365 585
R318 B.n364 B.n363 585
R319 B.n362 B.n361 585
R320 B.n360 B.n359 585
R321 B.n358 B.n357 585
R322 B.n356 B.n355 585
R323 B.n354 B.n353 585
R324 B.n352 B.n351 585
R325 B.n350 B.n349 585
R326 B.n348 B.n347 585
R327 B.n346 B.n345 585
R328 B.n344 B.n343 585
R329 B.n342 B.n341 585
R330 B.n340 B.n339 585
R331 B.n338 B.n337 585
R332 B.n336 B.n335 585
R333 B.n334 B.n333 585
R334 B.n332 B.n331 585
R335 B.n330 B.n329 585
R336 B.n328 B.n327 585
R337 B.n461 B.n286 585
R338 B.n286 B.n285 585
R339 B.n463 B.n462 585
R340 B.n464 B.n463 585
R341 B.n280 B.n279 585
R342 B.n281 B.n280 585
R343 B.n472 B.n471 585
R344 B.n471 B.n470 585
R345 B.n473 B.n278 585
R346 B.n278 B.n276 585
R347 B.n475 B.n474 585
R348 B.n476 B.n475 585
R349 B.n272 B.n271 585
R350 B.n277 B.n272 585
R351 B.n484 B.n483 585
R352 B.n483 B.n482 585
R353 B.n485 B.n270 585
R354 B.n270 B.n269 585
R355 B.n487 B.n486 585
R356 B.n488 B.n487 585
R357 B.n264 B.n263 585
R358 B.n265 B.n264 585
R359 B.n496 B.n495 585
R360 B.n495 B.n494 585
R361 B.n497 B.n262 585
R362 B.n262 B.n260 585
R363 B.n499 B.n498 585
R364 B.n500 B.n499 585
R365 B.n256 B.n255 585
R366 B.n261 B.n256 585
R367 B.n508 B.n507 585
R368 B.n507 B.n506 585
R369 B.n509 B.n254 585
R370 B.n254 B.n253 585
R371 B.n511 B.n510 585
R372 B.n512 B.n511 585
R373 B.n248 B.n247 585
R374 B.n249 B.n248 585
R375 B.n521 B.n520 585
R376 B.n520 B.n519 585
R377 B.n522 B.n246 585
R378 B.n518 B.n246 585
R379 B.n524 B.n523 585
R380 B.n525 B.n524 585
R381 B.n241 B.n240 585
R382 B.n242 B.n241 585
R383 B.n533 B.n532 585
R384 B.n532 B.n531 585
R385 B.n534 B.n239 585
R386 B.n239 B.n237 585
R387 B.n536 B.n535 585
R388 B.n537 B.n536 585
R389 B.n233 B.n232 585
R390 B.n238 B.n233 585
R391 B.n546 B.n545 585
R392 B.n545 B.n544 585
R393 B.n547 B.n231 585
R394 B.n231 B.n230 585
R395 B.n549 B.n548 585
R396 B.n550 B.n549 585
R397 B.n2 B.n0 585
R398 B.n4 B.n2 585
R399 B.n3 B.n1 585
R400 B.n659 B.n3 585
R401 B.n657 B.n656 585
R402 B.n658 B.n657 585
R403 B.n655 B.n9 585
R404 B.n9 B.n8 585
R405 B.n654 B.n653 585
R406 B.n653 B.n652 585
R407 B.n11 B.n10 585
R408 B.n651 B.n11 585
R409 B.n649 B.n648 585
R410 B.n650 B.n649 585
R411 B.n647 B.n16 585
R412 B.n16 B.n15 585
R413 B.n646 B.n645 585
R414 B.n645 B.n644 585
R415 B.n18 B.n17 585
R416 B.n643 B.n18 585
R417 B.n641 B.n640 585
R418 B.n642 B.n641 585
R419 B.n639 B.n22 585
R420 B.n25 B.n22 585
R421 B.n638 B.n637 585
R422 B.n637 B.n636 585
R423 B.n24 B.n23 585
R424 B.n635 B.n24 585
R425 B.n633 B.n632 585
R426 B.n634 B.n633 585
R427 B.n631 B.n30 585
R428 B.n30 B.n29 585
R429 B.n630 B.n629 585
R430 B.n629 B.n628 585
R431 B.n32 B.n31 585
R432 B.n627 B.n32 585
R433 B.n625 B.n624 585
R434 B.n626 B.n625 585
R435 B.n623 B.n37 585
R436 B.n37 B.n36 585
R437 B.n622 B.n621 585
R438 B.n621 B.n620 585
R439 B.n39 B.n38 585
R440 B.n619 B.n39 585
R441 B.n617 B.n616 585
R442 B.n618 B.n617 585
R443 B.n615 B.n44 585
R444 B.n44 B.n43 585
R445 B.n614 B.n613 585
R446 B.n613 B.n612 585
R447 B.n46 B.n45 585
R448 B.n611 B.n46 585
R449 B.n609 B.n608 585
R450 B.n610 B.n609 585
R451 B.n607 B.n51 585
R452 B.n51 B.n50 585
R453 B.n606 B.n605 585
R454 B.n605 B.n604 585
R455 B.n53 B.n52 585
R456 B.n603 B.n53 585
R457 B.n601 B.n600 585
R458 B.n602 B.n601 585
R459 B.n599 B.n58 585
R460 B.n58 B.n57 585
R461 B.n662 B.n661 585
R462 B.n661 B.n660 585
R463 B.n459 B.n286 492.5
R464 B.n597 B.n58 492.5
R465 B.n327 B.n284 492.5
R466 B.n594 B.n94 492.5
R467 B.n325 B.t6 317.375
R468 B.n322 B.t17 317.375
R469 B.n98 B.t10 317.375
R470 B.n95 B.t14 317.375
R471 B.n595 B.n92 256.663
R472 B.n595 B.n91 256.663
R473 B.n595 B.n90 256.663
R474 B.n595 B.n89 256.663
R475 B.n595 B.n88 256.663
R476 B.n595 B.n87 256.663
R477 B.n595 B.n86 256.663
R478 B.n595 B.n85 256.663
R479 B.n595 B.n84 256.663
R480 B.n595 B.n83 256.663
R481 B.n595 B.n82 256.663
R482 B.n595 B.n81 256.663
R483 B.n595 B.n80 256.663
R484 B.n595 B.n79 256.663
R485 B.n595 B.n78 256.663
R486 B.n595 B.n77 256.663
R487 B.n595 B.n76 256.663
R488 B.n595 B.n75 256.663
R489 B.n595 B.n74 256.663
R490 B.n595 B.n73 256.663
R491 B.n595 B.n72 256.663
R492 B.n595 B.n71 256.663
R493 B.n595 B.n70 256.663
R494 B.n595 B.n69 256.663
R495 B.n595 B.n68 256.663
R496 B.n595 B.n67 256.663
R497 B.n595 B.n66 256.663
R498 B.n595 B.n65 256.663
R499 B.n595 B.n64 256.663
R500 B.n595 B.n63 256.663
R501 B.n595 B.n62 256.663
R502 B.n595 B.n61 256.663
R503 B.n596 B.n595 256.663
R504 B.n458 B.n457 256.663
R505 B.n457 B.n289 256.663
R506 B.n457 B.n290 256.663
R507 B.n457 B.n291 256.663
R508 B.n457 B.n292 256.663
R509 B.n457 B.n293 256.663
R510 B.n457 B.n294 256.663
R511 B.n457 B.n295 256.663
R512 B.n457 B.n296 256.663
R513 B.n457 B.n297 256.663
R514 B.n457 B.n298 256.663
R515 B.n457 B.n299 256.663
R516 B.n457 B.n300 256.663
R517 B.n457 B.n301 256.663
R518 B.n457 B.n302 256.663
R519 B.n457 B.n303 256.663
R520 B.n457 B.n304 256.663
R521 B.n457 B.n305 256.663
R522 B.n457 B.n306 256.663
R523 B.n457 B.n307 256.663
R524 B.n457 B.n308 256.663
R525 B.n457 B.n309 256.663
R526 B.n457 B.n310 256.663
R527 B.n457 B.n311 256.663
R528 B.n457 B.n312 256.663
R529 B.n457 B.n313 256.663
R530 B.n457 B.n314 256.663
R531 B.n457 B.n315 256.663
R532 B.n457 B.n316 256.663
R533 B.n457 B.n317 256.663
R534 B.n457 B.n318 256.663
R535 B.n457 B.n319 256.663
R536 B.n457 B.n320 256.663
R537 B.n463 B.n286 163.367
R538 B.n463 B.n280 163.367
R539 B.n471 B.n280 163.367
R540 B.n471 B.n278 163.367
R541 B.n475 B.n278 163.367
R542 B.n475 B.n272 163.367
R543 B.n483 B.n272 163.367
R544 B.n483 B.n270 163.367
R545 B.n487 B.n270 163.367
R546 B.n487 B.n264 163.367
R547 B.n495 B.n264 163.367
R548 B.n495 B.n262 163.367
R549 B.n499 B.n262 163.367
R550 B.n499 B.n256 163.367
R551 B.n507 B.n256 163.367
R552 B.n507 B.n254 163.367
R553 B.n511 B.n254 163.367
R554 B.n511 B.n248 163.367
R555 B.n520 B.n248 163.367
R556 B.n520 B.n246 163.367
R557 B.n524 B.n246 163.367
R558 B.n524 B.n241 163.367
R559 B.n532 B.n241 163.367
R560 B.n532 B.n239 163.367
R561 B.n536 B.n239 163.367
R562 B.n536 B.n233 163.367
R563 B.n545 B.n233 163.367
R564 B.n545 B.n231 163.367
R565 B.n549 B.n231 163.367
R566 B.n549 B.n2 163.367
R567 B.n661 B.n2 163.367
R568 B.n661 B.n3 163.367
R569 B.n657 B.n3 163.367
R570 B.n657 B.n9 163.367
R571 B.n653 B.n9 163.367
R572 B.n653 B.n11 163.367
R573 B.n649 B.n11 163.367
R574 B.n649 B.n16 163.367
R575 B.n645 B.n16 163.367
R576 B.n645 B.n18 163.367
R577 B.n641 B.n18 163.367
R578 B.n641 B.n22 163.367
R579 B.n637 B.n22 163.367
R580 B.n637 B.n24 163.367
R581 B.n633 B.n24 163.367
R582 B.n633 B.n30 163.367
R583 B.n629 B.n30 163.367
R584 B.n629 B.n32 163.367
R585 B.n625 B.n32 163.367
R586 B.n625 B.n37 163.367
R587 B.n621 B.n37 163.367
R588 B.n621 B.n39 163.367
R589 B.n617 B.n39 163.367
R590 B.n617 B.n44 163.367
R591 B.n613 B.n44 163.367
R592 B.n613 B.n46 163.367
R593 B.n609 B.n46 163.367
R594 B.n609 B.n51 163.367
R595 B.n605 B.n51 163.367
R596 B.n605 B.n53 163.367
R597 B.n601 B.n53 163.367
R598 B.n601 B.n58 163.367
R599 B.n456 B.n288 163.367
R600 B.n456 B.n321 163.367
R601 B.n452 B.n451 163.367
R602 B.n448 B.n447 163.367
R603 B.n444 B.n443 163.367
R604 B.n440 B.n439 163.367
R605 B.n436 B.n435 163.367
R606 B.n432 B.n431 163.367
R607 B.n428 B.n427 163.367
R608 B.n424 B.n423 163.367
R609 B.n420 B.n419 163.367
R610 B.n416 B.n415 163.367
R611 B.n412 B.n411 163.367
R612 B.n408 B.n407 163.367
R613 B.n404 B.n403 163.367
R614 B.n400 B.n399 163.367
R615 B.n396 B.n395 163.367
R616 B.n392 B.n391 163.367
R617 B.n388 B.n387 163.367
R618 B.n383 B.n382 163.367
R619 B.n379 B.n378 163.367
R620 B.n375 B.n374 163.367
R621 B.n371 B.n370 163.367
R622 B.n367 B.n366 163.367
R623 B.n363 B.n362 163.367
R624 B.n359 B.n358 163.367
R625 B.n355 B.n354 163.367
R626 B.n351 B.n350 163.367
R627 B.n347 B.n346 163.367
R628 B.n343 B.n342 163.367
R629 B.n339 B.n338 163.367
R630 B.n335 B.n334 163.367
R631 B.n331 B.n330 163.367
R632 B.n465 B.n284 163.367
R633 B.n465 B.n282 163.367
R634 B.n469 B.n282 163.367
R635 B.n469 B.n275 163.367
R636 B.n477 B.n275 163.367
R637 B.n477 B.n273 163.367
R638 B.n481 B.n273 163.367
R639 B.n481 B.n268 163.367
R640 B.n489 B.n268 163.367
R641 B.n489 B.n266 163.367
R642 B.n493 B.n266 163.367
R643 B.n493 B.n259 163.367
R644 B.n501 B.n259 163.367
R645 B.n501 B.n257 163.367
R646 B.n505 B.n257 163.367
R647 B.n505 B.n252 163.367
R648 B.n513 B.n252 163.367
R649 B.n513 B.n250 163.367
R650 B.n517 B.n250 163.367
R651 B.n517 B.n245 163.367
R652 B.n526 B.n245 163.367
R653 B.n526 B.n243 163.367
R654 B.n530 B.n243 163.367
R655 B.n530 B.n236 163.367
R656 B.n538 B.n236 163.367
R657 B.n538 B.n234 163.367
R658 B.n543 B.n234 163.367
R659 B.n543 B.n229 163.367
R660 B.n551 B.n229 163.367
R661 B.n552 B.n551 163.367
R662 B.n552 B.n5 163.367
R663 B.n6 B.n5 163.367
R664 B.n7 B.n6 163.367
R665 B.n557 B.n7 163.367
R666 B.n557 B.n12 163.367
R667 B.n13 B.n12 163.367
R668 B.n14 B.n13 163.367
R669 B.n562 B.n14 163.367
R670 B.n562 B.n19 163.367
R671 B.n20 B.n19 163.367
R672 B.n21 B.n20 163.367
R673 B.n567 B.n21 163.367
R674 B.n567 B.n26 163.367
R675 B.n27 B.n26 163.367
R676 B.n28 B.n27 163.367
R677 B.n572 B.n28 163.367
R678 B.n572 B.n33 163.367
R679 B.n34 B.n33 163.367
R680 B.n35 B.n34 163.367
R681 B.n577 B.n35 163.367
R682 B.n577 B.n40 163.367
R683 B.n41 B.n40 163.367
R684 B.n42 B.n41 163.367
R685 B.n582 B.n42 163.367
R686 B.n582 B.n47 163.367
R687 B.n48 B.n47 163.367
R688 B.n49 B.n48 163.367
R689 B.n587 B.n49 163.367
R690 B.n587 B.n54 163.367
R691 B.n55 B.n54 163.367
R692 B.n56 B.n55 163.367
R693 B.n94 B.n56 163.367
R694 B.n100 B.n60 163.367
R695 B.n104 B.n103 163.367
R696 B.n108 B.n107 163.367
R697 B.n112 B.n111 163.367
R698 B.n116 B.n115 163.367
R699 B.n120 B.n119 163.367
R700 B.n124 B.n123 163.367
R701 B.n128 B.n127 163.367
R702 B.n132 B.n131 163.367
R703 B.n136 B.n135 163.367
R704 B.n140 B.n139 163.367
R705 B.n144 B.n143 163.367
R706 B.n148 B.n147 163.367
R707 B.n152 B.n151 163.367
R708 B.n157 B.n156 163.367
R709 B.n161 B.n160 163.367
R710 B.n165 B.n164 163.367
R711 B.n169 B.n168 163.367
R712 B.n173 B.n172 163.367
R713 B.n177 B.n176 163.367
R714 B.n181 B.n180 163.367
R715 B.n185 B.n184 163.367
R716 B.n189 B.n188 163.367
R717 B.n193 B.n192 163.367
R718 B.n197 B.n196 163.367
R719 B.n201 B.n200 163.367
R720 B.n205 B.n204 163.367
R721 B.n209 B.n208 163.367
R722 B.n213 B.n212 163.367
R723 B.n217 B.n216 163.367
R724 B.n221 B.n220 163.367
R725 B.n225 B.n224 163.367
R726 B.n594 B.n93 163.367
R727 B.n457 B.n285 115.88
R728 B.n595 B.n57 115.88
R729 B.n325 B.t9 107.936
R730 B.n95 B.t15 107.936
R731 B.n322 B.t19 107.927
R732 B.n98 B.t12 107.927
R733 B.n459 B.n458 71.676
R734 B.n321 B.n289 71.676
R735 B.n451 B.n290 71.676
R736 B.n447 B.n291 71.676
R737 B.n443 B.n292 71.676
R738 B.n439 B.n293 71.676
R739 B.n435 B.n294 71.676
R740 B.n431 B.n295 71.676
R741 B.n427 B.n296 71.676
R742 B.n423 B.n297 71.676
R743 B.n419 B.n298 71.676
R744 B.n415 B.n299 71.676
R745 B.n411 B.n300 71.676
R746 B.n407 B.n301 71.676
R747 B.n403 B.n302 71.676
R748 B.n399 B.n303 71.676
R749 B.n395 B.n304 71.676
R750 B.n391 B.n305 71.676
R751 B.n387 B.n306 71.676
R752 B.n382 B.n307 71.676
R753 B.n378 B.n308 71.676
R754 B.n374 B.n309 71.676
R755 B.n370 B.n310 71.676
R756 B.n366 B.n311 71.676
R757 B.n362 B.n312 71.676
R758 B.n358 B.n313 71.676
R759 B.n354 B.n314 71.676
R760 B.n350 B.n315 71.676
R761 B.n346 B.n316 71.676
R762 B.n342 B.n317 71.676
R763 B.n338 B.n318 71.676
R764 B.n334 B.n319 71.676
R765 B.n330 B.n320 71.676
R766 B.n597 B.n596 71.676
R767 B.n100 B.n61 71.676
R768 B.n104 B.n62 71.676
R769 B.n108 B.n63 71.676
R770 B.n112 B.n64 71.676
R771 B.n116 B.n65 71.676
R772 B.n120 B.n66 71.676
R773 B.n124 B.n67 71.676
R774 B.n128 B.n68 71.676
R775 B.n132 B.n69 71.676
R776 B.n136 B.n70 71.676
R777 B.n140 B.n71 71.676
R778 B.n144 B.n72 71.676
R779 B.n148 B.n73 71.676
R780 B.n152 B.n74 71.676
R781 B.n157 B.n75 71.676
R782 B.n161 B.n76 71.676
R783 B.n165 B.n77 71.676
R784 B.n169 B.n78 71.676
R785 B.n173 B.n79 71.676
R786 B.n177 B.n80 71.676
R787 B.n181 B.n81 71.676
R788 B.n185 B.n82 71.676
R789 B.n189 B.n83 71.676
R790 B.n193 B.n84 71.676
R791 B.n197 B.n85 71.676
R792 B.n201 B.n86 71.676
R793 B.n205 B.n87 71.676
R794 B.n209 B.n88 71.676
R795 B.n213 B.n89 71.676
R796 B.n217 B.n90 71.676
R797 B.n221 B.n91 71.676
R798 B.n225 B.n92 71.676
R799 B.n93 B.n92 71.676
R800 B.n224 B.n91 71.676
R801 B.n220 B.n90 71.676
R802 B.n216 B.n89 71.676
R803 B.n212 B.n88 71.676
R804 B.n208 B.n87 71.676
R805 B.n204 B.n86 71.676
R806 B.n200 B.n85 71.676
R807 B.n196 B.n84 71.676
R808 B.n192 B.n83 71.676
R809 B.n188 B.n82 71.676
R810 B.n184 B.n81 71.676
R811 B.n180 B.n80 71.676
R812 B.n176 B.n79 71.676
R813 B.n172 B.n78 71.676
R814 B.n168 B.n77 71.676
R815 B.n164 B.n76 71.676
R816 B.n160 B.n75 71.676
R817 B.n156 B.n74 71.676
R818 B.n151 B.n73 71.676
R819 B.n147 B.n72 71.676
R820 B.n143 B.n71 71.676
R821 B.n139 B.n70 71.676
R822 B.n135 B.n69 71.676
R823 B.n131 B.n68 71.676
R824 B.n127 B.n67 71.676
R825 B.n123 B.n66 71.676
R826 B.n119 B.n65 71.676
R827 B.n115 B.n64 71.676
R828 B.n111 B.n63 71.676
R829 B.n107 B.n62 71.676
R830 B.n103 B.n61 71.676
R831 B.n596 B.n60 71.676
R832 B.n458 B.n288 71.676
R833 B.n452 B.n289 71.676
R834 B.n448 B.n290 71.676
R835 B.n444 B.n291 71.676
R836 B.n440 B.n292 71.676
R837 B.n436 B.n293 71.676
R838 B.n432 B.n294 71.676
R839 B.n428 B.n295 71.676
R840 B.n424 B.n296 71.676
R841 B.n420 B.n297 71.676
R842 B.n416 B.n298 71.676
R843 B.n412 B.n299 71.676
R844 B.n408 B.n300 71.676
R845 B.n404 B.n301 71.676
R846 B.n400 B.n302 71.676
R847 B.n396 B.n303 71.676
R848 B.n392 B.n304 71.676
R849 B.n388 B.n305 71.676
R850 B.n383 B.n306 71.676
R851 B.n379 B.n307 71.676
R852 B.n375 B.n308 71.676
R853 B.n371 B.n309 71.676
R854 B.n367 B.n310 71.676
R855 B.n363 B.n311 71.676
R856 B.n359 B.n312 71.676
R857 B.n355 B.n313 71.676
R858 B.n351 B.n314 71.676
R859 B.n347 B.n315 71.676
R860 B.n343 B.n316 71.676
R861 B.n339 B.n317 71.676
R862 B.n335 B.n318 71.676
R863 B.n331 B.n319 71.676
R864 B.n327 B.n320 71.676
R865 B.n326 B.t8 69.9244
R866 B.n96 B.t16 69.9244
R867 B.n323 B.t18 69.9157
R868 B.n99 B.t13 69.9157
R869 B.n385 B.n326 59.5399
R870 B.n324 B.n323 59.5399
R871 B.n154 B.n99 59.5399
R872 B.n97 B.n96 59.5399
R873 B.n464 B.n285 58.3696
R874 B.n464 B.n281 58.3696
R875 B.n470 B.n281 58.3696
R876 B.n470 B.n276 58.3696
R877 B.n476 B.n276 58.3696
R878 B.n476 B.n277 58.3696
R879 B.n482 B.n269 58.3696
R880 B.n488 B.n269 58.3696
R881 B.n488 B.n265 58.3696
R882 B.n494 B.n265 58.3696
R883 B.n494 B.n260 58.3696
R884 B.n500 B.n260 58.3696
R885 B.n500 B.n261 58.3696
R886 B.n506 B.n253 58.3696
R887 B.n512 B.n253 58.3696
R888 B.n512 B.n249 58.3696
R889 B.n519 B.n249 58.3696
R890 B.n519 B.n518 58.3696
R891 B.n525 B.n242 58.3696
R892 B.n531 B.n242 58.3696
R893 B.n531 B.n237 58.3696
R894 B.n537 B.n237 58.3696
R895 B.n537 B.n238 58.3696
R896 B.n544 B.n230 58.3696
R897 B.n550 B.n230 58.3696
R898 B.n550 B.n4 58.3696
R899 B.n660 B.n4 58.3696
R900 B.n660 B.n659 58.3696
R901 B.n659 B.n658 58.3696
R902 B.n658 B.n8 58.3696
R903 B.n652 B.n8 58.3696
R904 B.n651 B.n650 58.3696
R905 B.n650 B.n15 58.3696
R906 B.n644 B.n15 58.3696
R907 B.n644 B.n643 58.3696
R908 B.n643 B.n642 58.3696
R909 B.n636 B.n25 58.3696
R910 B.n636 B.n635 58.3696
R911 B.n635 B.n634 58.3696
R912 B.n634 B.n29 58.3696
R913 B.n628 B.n29 58.3696
R914 B.n627 B.n626 58.3696
R915 B.n626 B.n36 58.3696
R916 B.n620 B.n36 58.3696
R917 B.n620 B.n619 58.3696
R918 B.n619 B.n618 58.3696
R919 B.n618 B.n43 58.3696
R920 B.n612 B.n43 58.3696
R921 B.n611 B.n610 58.3696
R922 B.n610 B.n50 58.3696
R923 B.n604 B.n50 58.3696
R924 B.n604 B.n603 58.3696
R925 B.n603 B.n602 58.3696
R926 B.n602 B.n57 58.3696
R927 B.n482 B.t7 57.5112
R928 B.n261 B.t1 57.5112
R929 B.t0 B.n627 57.5112
R930 B.n612 B.t11 57.5112
R931 B.n518 B.t2 43.7773
R932 B.n25 B.t3 43.7773
R933 B.n326 B.n325 38.0126
R934 B.n323 B.n322 38.0126
R935 B.n99 B.n98 38.0126
R936 B.n96 B.n95 38.0126
R937 B.n599 B.n598 32.0005
R938 B.n593 B.n592 32.0005
R939 B.n328 B.n283 32.0005
R940 B.n461 B.n460 32.0005
R941 B.n238 B.t4 30.0434
R942 B.t5 B.n651 30.0434
R943 B.n544 B.t4 28.3267
R944 B.n652 B.t5 28.3267
R945 B B.n662 18.0485
R946 B.n525 B.t2 14.5928
R947 B.n642 B.t3 14.5928
R948 B.n598 B.n59 10.6151
R949 B.n101 B.n59 10.6151
R950 B.n102 B.n101 10.6151
R951 B.n105 B.n102 10.6151
R952 B.n106 B.n105 10.6151
R953 B.n109 B.n106 10.6151
R954 B.n110 B.n109 10.6151
R955 B.n113 B.n110 10.6151
R956 B.n114 B.n113 10.6151
R957 B.n117 B.n114 10.6151
R958 B.n118 B.n117 10.6151
R959 B.n121 B.n118 10.6151
R960 B.n122 B.n121 10.6151
R961 B.n125 B.n122 10.6151
R962 B.n126 B.n125 10.6151
R963 B.n129 B.n126 10.6151
R964 B.n130 B.n129 10.6151
R965 B.n133 B.n130 10.6151
R966 B.n134 B.n133 10.6151
R967 B.n137 B.n134 10.6151
R968 B.n138 B.n137 10.6151
R969 B.n141 B.n138 10.6151
R970 B.n142 B.n141 10.6151
R971 B.n145 B.n142 10.6151
R972 B.n146 B.n145 10.6151
R973 B.n149 B.n146 10.6151
R974 B.n150 B.n149 10.6151
R975 B.n153 B.n150 10.6151
R976 B.n158 B.n155 10.6151
R977 B.n159 B.n158 10.6151
R978 B.n162 B.n159 10.6151
R979 B.n163 B.n162 10.6151
R980 B.n166 B.n163 10.6151
R981 B.n167 B.n166 10.6151
R982 B.n170 B.n167 10.6151
R983 B.n171 B.n170 10.6151
R984 B.n175 B.n174 10.6151
R985 B.n178 B.n175 10.6151
R986 B.n179 B.n178 10.6151
R987 B.n182 B.n179 10.6151
R988 B.n183 B.n182 10.6151
R989 B.n186 B.n183 10.6151
R990 B.n187 B.n186 10.6151
R991 B.n190 B.n187 10.6151
R992 B.n191 B.n190 10.6151
R993 B.n194 B.n191 10.6151
R994 B.n195 B.n194 10.6151
R995 B.n198 B.n195 10.6151
R996 B.n199 B.n198 10.6151
R997 B.n202 B.n199 10.6151
R998 B.n203 B.n202 10.6151
R999 B.n206 B.n203 10.6151
R1000 B.n207 B.n206 10.6151
R1001 B.n210 B.n207 10.6151
R1002 B.n211 B.n210 10.6151
R1003 B.n214 B.n211 10.6151
R1004 B.n215 B.n214 10.6151
R1005 B.n218 B.n215 10.6151
R1006 B.n219 B.n218 10.6151
R1007 B.n222 B.n219 10.6151
R1008 B.n223 B.n222 10.6151
R1009 B.n226 B.n223 10.6151
R1010 B.n227 B.n226 10.6151
R1011 B.n593 B.n227 10.6151
R1012 B.n466 B.n283 10.6151
R1013 B.n467 B.n466 10.6151
R1014 B.n468 B.n467 10.6151
R1015 B.n468 B.n274 10.6151
R1016 B.n478 B.n274 10.6151
R1017 B.n479 B.n478 10.6151
R1018 B.n480 B.n479 10.6151
R1019 B.n480 B.n267 10.6151
R1020 B.n490 B.n267 10.6151
R1021 B.n491 B.n490 10.6151
R1022 B.n492 B.n491 10.6151
R1023 B.n492 B.n258 10.6151
R1024 B.n502 B.n258 10.6151
R1025 B.n503 B.n502 10.6151
R1026 B.n504 B.n503 10.6151
R1027 B.n504 B.n251 10.6151
R1028 B.n514 B.n251 10.6151
R1029 B.n515 B.n514 10.6151
R1030 B.n516 B.n515 10.6151
R1031 B.n516 B.n244 10.6151
R1032 B.n527 B.n244 10.6151
R1033 B.n528 B.n527 10.6151
R1034 B.n529 B.n528 10.6151
R1035 B.n529 B.n235 10.6151
R1036 B.n539 B.n235 10.6151
R1037 B.n540 B.n539 10.6151
R1038 B.n542 B.n540 10.6151
R1039 B.n542 B.n541 10.6151
R1040 B.n541 B.n228 10.6151
R1041 B.n553 B.n228 10.6151
R1042 B.n554 B.n553 10.6151
R1043 B.n555 B.n554 10.6151
R1044 B.n556 B.n555 10.6151
R1045 B.n558 B.n556 10.6151
R1046 B.n559 B.n558 10.6151
R1047 B.n560 B.n559 10.6151
R1048 B.n561 B.n560 10.6151
R1049 B.n563 B.n561 10.6151
R1050 B.n564 B.n563 10.6151
R1051 B.n565 B.n564 10.6151
R1052 B.n566 B.n565 10.6151
R1053 B.n568 B.n566 10.6151
R1054 B.n569 B.n568 10.6151
R1055 B.n570 B.n569 10.6151
R1056 B.n571 B.n570 10.6151
R1057 B.n573 B.n571 10.6151
R1058 B.n574 B.n573 10.6151
R1059 B.n575 B.n574 10.6151
R1060 B.n576 B.n575 10.6151
R1061 B.n578 B.n576 10.6151
R1062 B.n579 B.n578 10.6151
R1063 B.n580 B.n579 10.6151
R1064 B.n581 B.n580 10.6151
R1065 B.n583 B.n581 10.6151
R1066 B.n584 B.n583 10.6151
R1067 B.n585 B.n584 10.6151
R1068 B.n586 B.n585 10.6151
R1069 B.n588 B.n586 10.6151
R1070 B.n589 B.n588 10.6151
R1071 B.n590 B.n589 10.6151
R1072 B.n591 B.n590 10.6151
R1073 B.n592 B.n591 10.6151
R1074 B.n460 B.n287 10.6151
R1075 B.n455 B.n287 10.6151
R1076 B.n455 B.n454 10.6151
R1077 B.n454 B.n453 10.6151
R1078 B.n453 B.n450 10.6151
R1079 B.n450 B.n449 10.6151
R1080 B.n449 B.n446 10.6151
R1081 B.n446 B.n445 10.6151
R1082 B.n445 B.n442 10.6151
R1083 B.n442 B.n441 10.6151
R1084 B.n441 B.n438 10.6151
R1085 B.n438 B.n437 10.6151
R1086 B.n437 B.n434 10.6151
R1087 B.n434 B.n433 10.6151
R1088 B.n433 B.n430 10.6151
R1089 B.n430 B.n429 10.6151
R1090 B.n429 B.n426 10.6151
R1091 B.n426 B.n425 10.6151
R1092 B.n425 B.n422 10.6151
R1093 B.n422 B.n421 10.6151
R1094 B.n421 B.n418 10.6151
R1095 B.n418 B.n417 10.6151
R1096 B.n417 B.n414 10.6151
R1097 B.n414 B.n413 10.6151
R1098 B.n413 B.n410 10.6151
R1099 B.n410 B.n409 10.6151
R1100 B.n409 B.n406 10.6151
R1101 B.n406 B.n405 10.6151
R1102 B.n402 B.n401 10.6151
R1103 B.n401 B.n398 10.6151
R1104 B.n398 B.n397 10.6151
R1105 B.n397 B.n394 10.6151
R1106 B.n394 B.n393 10.6151
R1107 B.n393 B.n390 10.6151
R1108 B.n390 B.n389 10.6151
R1109 B.n389 B.n386 10.6151
R1110 B.n384 B.n381 10.6151
R1111 B.n381 B.n380 10.6151
R1112 B.n380 B.n377 10.6151
R1113 B.n377 B.n376 10.6151
R1114 B.n376 B.n373 10.6151
R1115 B.n373 B.n372 10.6151
R1116 B.n372 B.n369 10.6151
R1117 B.n369 B.n368 10.6151
R1118 B.n368 B.n365 10.6151
R1119 B.n365 B.n364 10.6151
R1120 B.n364 B.n361 10.6151
R1121 B.n361 B.n360 10.6151
R1122 B.n360 B.n357 10.6151
R1123 B.n357 B.n356 10.6151
R1124 B.n356 B.n353 10.6151
R1125 B.n353 B.n352 10.6151
R1126 B.n352 B.n349 10.6151
R1127 B.n349 B.n348 10.6151
R1128 B.n348 B.n345 10.6151
R1129 B.n345 B.n344 10.6151
R1130 B.n344 B.n341 10.6151
R1131 B.n341 B.n340 10.6151
R1132 B.n340 B.n337 10.6151
R1133 B.n337 B.n336 10.6151
R1134 B.n336 B.n333 10.6151
R1135 B.n333 B.n332 10.6151
R1136 B.n332 B.n329 10.6151
R1137 B.n329 B.n328 10.6151
R1138 B.n462 B.n461 10.6151
R1139 B.n462 B.n279 10.6151
R1140 B.n472 B.n279 10.6151
R1141 B.n473 B.n472 10.6151
R1142 B.n474 B.n473 10.6151
R1143 B.n474 B.n271 10.6151
R1144 B.n484 B.n271 10.6151
R1145 B.n485 B.n484 10.6151
R1146 B.n486 B.n485 10.6151
R1147 B.n486 B.n263 10.6151
R1148 B.n496 B.n263 10.6151
R1149 B.n497 B.n496 10.6151
R1150 B.n498 B.n497 10.6151
R1151 B.n498 B.n255 10.6151
R1152 B.n508 B.n255 10.6151
R1153 B.n509 B.n508 10.6151
R1154 B.n510 B.n509 10.6151
R1155 B.n510 B.n247 10.6151
R1156 B.n521 B.n247 10.6151
R1157 B.n522 B.n521 10.6151
R1158 B.n523 B.n522 10.6151
R1159 B.n523 B.n240 10.6151
R1160 B.n533 B.n240 10.6151
R1161 B.n534 B.n533 10.6151
R1162 B.n535 B.n534 10.6151
R1163 B.n535 B.n232 10.6151
R1164 B.n546 B.n232 10.6151
R1165 B.n547 B.n546 10.6151
R1166 B.n548 B.n547 10.6151
R1167 B.n548 B.n0 10.6151
R1168 B.n656 B.n1 10.6151
R1169 B.n656 B.n655 10.6151
R1170 B.n655 B.n654 10.6151
R1171 B.n654 B.n10 10.6151
R1172 B.n648 B.n10 10.6151
R1173 B.n648 B.n647 10.6151
R1174 B.n647 B.n646 10.6151
R1175 B.n646 B.n17 10.6151
R1176 B.n640 B.n17 10.6151
R1177 B.n640 B.n639 10.6151
R1178 B.n639 B.n638 10.6151
R1179 B.n638 B.n23 10.6151
R1180 B.n632 B.n23 10.6151
R1181 B.n632 B.n631 10.6151
R1182 B.n631 B.n630 10.6151
R1183 B.n630 B.n31 10.6151
R1184 B.n624 B.n31 10.6151
R1185 B.n624 B.n623 10.6151
R1186 B.n623 B.n622 10.6151
R1187 B.n622 B.n38 10.6151
R1188 B.n616 B.n38 10.6151
R1189 B.n616 B.n615 10.6151
R1190 B.n615 B.n614 10.6151
R1191 B.n614 B.n45 10.6151
R1192 B.n608 B.n45 10.6151
R1193 B.n608 B.n607 10.6151
R1194 B.n607 B.n606 10.6151
R1195 B.n606 B.n52 10.6151
R1196 B.n600 B.n52 10.6151
R1197 B.n600 B.n599 10.6151
R1198 B.n155 B.n154 6.5566
R1199 B.n171 B.n97 6.5566
R1200 B.n402 B.n324 6.5566
R1201 B.n386 B.n385 6.5566
R1202 B.n154 B.n153 4.05904
R1203 B.n174 B.n97 4.05904
R1204 B.n405 B.n324 4.05904
R1205 B.n385 B.n384 4.05904
R1206 B.n662 B.n0 2.81026
R1207 B.n662 B.n1 2.81026
R1208 B.n277 B.t7 0.858869
R1209 B.n506 B.t1 0.858869
R1210 B.n628 B.t0 0.858869
R1211 B.t11 B.n611 0.858869
R1212 VP.n17 VP.n16 175.564
R1213 VP.n32 VP.n31 175.564
R1214 VP.n15 VP.n14 175.564
R1215 VP.n9 VP.n8 161.3
R1216 VP.n10 VP.n5 161.3
R1217 VP.n12 VP.n11 161.3
R1218 VP.n13 VP.n4 161.3
R1219 VP.n30 VP.n0 161.3
R1220 VP.n29 VP.n28 161.3
R1221 VP.n27 VP.n1 161.3
R1222 VP.n26 VP.n25 161.3
R1223 VP.n23 VP.n2 161.3
R1224 VP.n22 VP.n21 161.3
R1225 VP.n20 VP.n3 161.3
R1226 VP.n19 VP.n18 161.3
R1227 VP.n6 VP.t0 145.44
R1228 VP.n17 VP.t5 111.481
R1229 VP.n24 VP.t3 111.481
R1230 VP.n31 VP.t1 111.481
R1231 VP.n14 VP.t4 111.481
R1232 VP.n7 VP.t2 111.481
R1233 VP.n22 VP.n3 56.5617
R1234 VP.n29 VP.n1 56.5617
R1235 VP.n12 VP.n5 56.5617
R1236 VP.n7 VP.n6 54.3154
R1237 VP.n16 VP.n15 41.455
R1238 VP.n18 VP.n3 24.5923
R1239 VP.n23 VP.n22 24.5923
R1240 VP.n25 VP.n1 24.5923
R1241 VP.n30 VP.n29 24.5923
R1242 VP.n13 VP.n12 24.5923
R1243 VP.n8 VP.n5 24.5923
R1244 VP.n9 VP.n6 17.7323
R1245 VP.n24 VP.n23 12.2964
R1246 VP.n25 VP.n24 12.2964
R1247 VP.n8 VP.n7 12.2964
R1248 VP.n18 VP.n17 10.3291
R1249 VP.n31 VP.n30 10.3291
R1250 VP.n14 VP.n13 10.3291
R1251 VP.n10 VP.n9 0.189894
R1252 VP.n11 VP.n10 0.189894
R1253 VP.n11 VP.n4 0.189894
R1254 VP.n15 VP.n4 0.189894
R1255 VP.n19 VP.n16 0.189894
R1256 VP.n20 VP.n19 0.189894
R1257 VP.n21 VP.n20 0.189894
R1258 VP.n21 VP.n2 0.189894
R1259 VP.n26 VP.n2 0.189894
R1260 VP.n27 VP.n26 0.189894
R1261 VP.n28 VP.n27 0.189894
R1262 VP.n28 VP.n0 0.189894
R1263 VP.n32 VP.n0 0.189894
R1264 VP VP.n32 0.0516364
R1265 VDD1 VDD1.t5 70.1821
R1266 VDD1.n1 VDD1.t0 70.0684
R1267 VDD1.n1 VDD1.n0 66.5975
R1268 VDD1.n3 VDD1.n2 66.2305
R1269 VDD1.n3 VDD1.n1 37.1345
R1270 VDD1.n2 VDD1.t3 2.62649
R1271 VDD1.n2 VDD1.t1 2.62649
R1272 VDD1.n0 VDD1.t2 2.62649
R1273 VDD1.n0 VDD1.t4 2.62649
R1274 VDD1 VDD1.n3 0.364724
C0 VP VDD2 0.376098f
C1 VP VTAIL 4.04585f
C2 VP VDD1 4.14005f
C3 VN VDD2 3.9163f
C4 VN VTAIL 4.03156f
C5 VN VDD1 0.149814f
C6 VDD2 VTAIL 5.96927f
C7 VDD2 VDD1 1.05594f
C8 VTAIL VDD1 5.92481f
C9 VN VP 5.15179f
C10 VDD2 B 4.415565f
C11 VDD1 B 4.684105f
C12 VTAIL B 5.411818f
C13 VN B 9.702109f
C14 VP B 8.256904f
C15 VDD1.t5 B 1.43755f
C16 VDD1.t0 B 1.43689f
C17 VDD1.t2 B 0.130721f
C18 VDD1.t4 B 0.130721f
C19 VDD1.n0 B 1.12824f
C20 VDD1.n1 B 2.01148f
C21 VDD1.t3 B 0.130721f
C22 VDD1.t1 B 0.130721f
C23 VDD1.n2 B 1.12642f
C24 VDD1.n3 B 1.89594f
C25 VP.n0 B 0.032869f
C26 VP.t1 B 1.08207f
C27 VP.n1 B 0.045962f
C28 VP.n2 B 0.032869f
C29 VP.t3 B 1.08207f
C30 VP.n3 B 0.0496f
C31 VP.n4 B 0.032869f
C32 VP.t4 B 1.08207f
C33 VP.n5 B 0.045962f
C34 VP.t0 B 1.20906f
C35 VP.n6 B 0.479431f
C36 VP.t2 B 1.08207f
C37 VP.n7 B 0.471919f
C38 VP.n8 B 0.045908f
C39 VP.n9 B 0.211338f
C40 VP.n10 B 0.032869f
C41 VP.n11 B 0.032869f
C42 VP.n12 B 0.0496f
C43 VP.n13 B 0.0435f
C44 VP.n14 B 0.482265f
C45 VP.n15 B 1.33398f
C46 VP.n16 B 1.36257f
C47 VP.t5 B 1.08207f
C48 VP.n17 B 0.482265f
C49 VP.n18 B 0.0435f
C50 VP.n19 B 0.032869f
C51 VP.n20 B 0.032869f
C52 VP.n21 B 0.032869f
C53 VP.n22 B 0.045962f
C54 VP.n23 B 0.045908f
C55 VP.n24 B 0.407464f
C56 VP.n25 B 0.045908f
C57 VP.n26 B 0.032869f
C58 VP.n27 B 0.032869f
C59 VP.n28 B 0.032869f
C60 VP.n29 B 0.0496f
C61 VP.n30 B 0.0435f
C62 VP.n31 B 0.482265f
C63 VP.n32 B 0.032087f
C64 VTAIL.t8 B 0.146931f
C65 VTAIL.t6 B 0.146931f
C66 VTAIL.n0 B 1.20215f
C67 VTAIL.n1 B 0.367799f
C68 VTAIL.t10 B 1.52959f
C69 VTAIL.n2 B 0.537144f
C70 VTAIL.t1 B 0.146931f
C71 VTAIL.t2 B 0.146931f
C72 VTAIL.n3 B 1.20215f
C73 VTAIL.n4 B 1.47938f
C74 VTAIL.t5 B 0.146931f
C75 VTAIL.t9 B 0.146931f
C76 VTAIL.n5 B 1.20215f
C77 VTAIL.n6 B 1.47938f
C78 VTAIL.t4 B 1.5296f
C79 VTAIL.n7 B 0.537141f
C80 VTAIL.t11 B 0.146931f
C81 VTAIL.t3 B 0.146931f
C82 VTAIL.n8 B 1.20215f
C83 VTAIL.n9 B 0.463866f
C84 VTAIL.t0 B 1.52959f
C85 VTAIL.n10 B 1.4184f
C86 VTAIL.t7 B 1.52959f
C87 VTAIL.n11 B 1.38021f
C88 VDD2.t4 B 1.43415f
C89 VDD2.t1 B 0.130471f
C90 VDD2.t2 B 0.130471f
C91 VDD2.n0 B 1.12608f
C92 VDD2.n1 B 1.92316f
C93 VDD2.t0 B 1.42863f
C94 VDD2.n2 B 1.89598f
C95 VDD2.t3 B 0.130471f
C96 VDD2.t5 B 0.130471f
C97 VDD2.n3 B 1.12606f
C98 VN.n0 B 0.032263f
C99 VN.t2 B 1.06211f
C100 VN.n1 B 0.045114f
C101 VN.t1 B 1.18675f
C102 VN.n2 B 0.470587f
C103 VN.t3 B 1.06211f
C104 VN.n3 B 0.463213f
C105 VN.n4 B 0.045061f
C106 VN.n5 B 0.20744f
C107 VN.n6 B 0.032263f
C108 VN.n7 B 0.032263f
C109 VN.n8 B 0.048685f
C110 VN.n9 B 0.042698f
C111 VN.n10 B 0.473368f
C112 VN.n11 B 0.031495f
C113 VN.n12 B 0.032263f
C114 VN.t4 B 1.06211f
C115 VN.n13 B 0.045114f
C116 VN.t5 B 1.18675f
C117 VN.n14 B 0.470587f
C118 VN.t0 B 1.06211f
C119 VN.n15 B 0.463213f
C120 VN.n16 B 0.045061f
C121 VN.n17 B 0.20744f
C122 VN.n18 B 0.032263f
C123 VN.n19 B 0.032263f
C124 VN.n20 B 0.048685f
C125 VN.n21 B 0.042698f
C126 VN.n22 B 0.473368f
C127 VN.n23 B 1.33057f
.ends

