* NGSPICE file created from diff_pair_sample_0708.ext - technology: sky130A

.subckt diff_pair_sample_0708 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t16 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=6.9498 pd=36.42 as=2.9403 ps=18.15 w=17.82 l=1.94
X1 VDD1.t8 VP.t1 VTAIL.t15 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=6.9498 pd=36.42 as=2.9403 ps=18.15 w=17.82 l=1.94
X2 VDD1.t7 VP.t2 VTAIL.t11 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=2.9403 pd=18.15 as=6.9498 ps=36.42 w=17.82 l=1.94
X3 VTAIL.t10 VP.t3 VDD1.t6 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=2.9403 pd=18.15 as=2.9403 ps=18.15 w=17.82 l=1.94
X4 B.t11 B.t9 B.t10 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=6.9498 pd=36.42 as=0 ps=0 w=17.82 l=1.94
X5 VDD2.t9 VN.t0 VTAIL.t4 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=2.9403 pd=18.15 as=2.9403 ps=18.15 w=17.82 l=1.94
X6 B.t8 B.t6 B.t7 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=6.9498 pd=36.42 as=0 ps=0 w=17.82 l=1.94
X7 VTAIL.t14 VP.t4 VDD1.t5 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=2.9403 pd=18.15 as=2.9403 ps=18.15 w=17.82 l=1.94
X8 VDD1.t4 VP.t5 VTAIL.t13 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=2.9403 pd=18.15 as=2.9403 ps=18.15 w=17.82 l=1.94
X9 VDD2.t8 VN.t1 VTAIL.t19 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=2.9403 pd=18.15 as=6.9498 ps=36.42 w=17.82 l=1.94
X10 VTAIL.t18 VN.t2 VDD2.t7 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=2.9403 pd=18.15 as=2.9403 ps=18.15 w=17.82 l=1.94
X11 VDD2.t6 VN.t3 VTAIL.t5 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=2.9403 pd=18.15 as=2.9403 ps=18.15 w=17.82 l=1.94
X12 VDD1.t3 VP.t6 VTAIL.t12 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=2.9403 pd=18.15 as=2.9403 ps=18.15 w=17.82 l=1.94
X13 VTAIL.t6 VN.t4 VDD2.t5 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=2.9403 pd=18.15 as=2.9403 ps=18.15 w=17.82 l=1.94
X14 VTAIL.t17 VN.t5 VDD2.t4 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=2.9403 pd=18.15 as=2.9403 ps=18.15 w=17.82 l=1.94
X15 B.t5 B.t3 B.t4 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=6.9498 pd=36.42 as=0 ps=0 w=17.82 l=1.94
X16 VTAIL.t7 VP.t7 VDD1.t2 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=2.9403 pd=18.15 as=2.9403 ps=18.15 w=17.82 l=1.94
X17 VDD2.t3 VN.t6 VTAIL.t3 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=2.9403 pd=18.15 as=6.9498 ps=36.42 w=17.82 l=1.94
X18 VTAIL.t9 VP.t8 VDD1.t1 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=2.9403 pd=18.15 as=2.9403 ps=18.15 w=17.82 l=1.94
X19 VTAIL.t1 VN.t7 VDD2.t2 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=2.9403 pd=18.15 as=2.9403 ps=18.15 w=17.82 l=1.94
X20 VDD1.t0 VP.t9 VTAIL.t8 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=2.9403 pd=18.15 as=6.9498 ps=36.42 w=17.82 l=1.94
X21 B.t2 B.t0 B.t1 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=6.9498 pd=36.42 as=0 ps=0 w=17.82 l=1.94
X22 VDD2.t1 VN.t8 VTAIL.t0 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=6.9498 pd=36.42 as=2.9403 ps=18.15 w=17.82 l=1.94
X23 VDD2.t0 VN.t9 VTAIL.t2 w_n3694_n4532# sky130_fd_pr__pfet_01v8 ad=6.9498 pd=36.42 as=2.9403 ps=18.15 w=17.82 l=1.94
R0 VP.n18 VP.t1 254.249
R1 VP.n60 VP.t5 221.373
R2 VP.n44 VP.t0 221.373
R3 VP.n7 VP.t7 221.373
R4 VP.n67 VP.t3 221.373
R5 VP.n75 VP.t9 221.373
R6 VP.n26 VP.t6 221.373
R7 VP.n41 VP.t2 221.373
R8 VP.n33 VP.t8 221.373
R9 VP.n17 VP.t4 221.373
R10 VP.n44 VP.n43 183.924
R11 VP.n76 VP.n75 183.924
R12 VP.n42 VP.n41 183.924
R13 VP.n20 VP.n19 161.3
R14 VP.n21 VP.n16 161.3
R15 VP.n23 VP.n22 161.3
R16 VP.n24 VP.n15 161.3
R17 VP.n26 VP.n25 161.3
R18 VP.n27 VP.n14 161.3
R19 VP.n29 VP.n28 161.3
R20 VP.n30 VP.n13 161.3
R21 VP.n32 VP.n31 161.3
R22 VP.n34 VP.n12 161.3
R23 VP.n36 VP.n35 161.3
R24 VP.n37 VP.n11 161.3
R25 VP.n39 VP.n38 161.3
R26 VP.n40 VP.n10 161.3
R27 VP.n74 VP.n0 161.3
R28 VP.n73 VP.n72 161.3
R29 VP.n71 VP.n1 161.3
R30 VP.n70 VP.n69 161.3
R31 VP.n68 VP.n2 161.3
R32 VP.n66 VP.n65 161.3
R33 VP.n64 VP.n3 161.3
R34 VP.n63 VP.n62 161.3
R35 VP.n61 VP.n4 161.3
R36 VP.n60 VP.n59 161.3
R37 VP.n58 VP.n5 161.3
R38 VP.n57 VP.n56 161.3
R39 VP.n55 VP.n6 161.3
R40 VP.n54 VP.n53 161.3
R41 VP.n52 VP.n51 161.3
R42 VP.n50 VP.n8 161.3
R43 VP.n49 VP.n48 161.3
R44 VP.n47 VP.n9 161.3
R45 VP.n46 VP.n45 161.3
R46 VP.n18 VP.n17 56.9995
R47 VP.n43 VP.n42 53.8452
R48 VP.n56 VP.n55 53.6554
R49 VP.n62 VP.n3 53.6554
R50 VP.n28 VP.n13 53.6554
R51 VP.n22 VP.n21 53.6554
R52 VP.n50 VP.n49 49.7803
R53 VP.n69 VP.n1 49.7803
R54 VP.n35 VP.n11 49.7803
R55 VP.n49 VP.n9 31.3737
R56 VP.n73 VP.n1 31.3737
R57 VP.n39 VP.n11 31.3737
R58 VP.n56 VP.n5 27.4986
R59 VP.n62 VP.n61 27.4986
R60 VP.n28 VP.n27 27.4986
R61 VP.n22 VP.n15 27.4986
R62 VP.n45 VP.n9 24.5923
R63 VP.n51 VP.n50 24.5923
R64 VP.n55 VP.n54 24.5923
R65 VP.n60 VP.n5 24.5923
R66 VP.n61 VP.n60 24.5923
R67 VP.n66 VP.n3 24.5923
R68 VP.n69 VP.n68 24.5923
R69 VP.n74 VP.n73 24.5923
R70 VP.n40 VP.n39 24.5923
R71 VP.n32 VP.n13 24.5923
R72 VP.n35 VP.n34 24.5923
R73 VP.n26 VP.n15 24.5923
R74 VP.n27 VP.n26 24.5923
R75 VP.n21 VP.n20 24.5923
R76 VP.n54 VP.n7 13.2801
R77 VP.n67 VP.n66 13.2801
R78 VP.n33 VP.n32 13.2801
R79 VP.n20 VP.n17 13.2801
R80 VP.n19 VP.n18 12.447
R81 VP.n51 VP.n7 11.3127
R82 VP.n68 VP.n67 11.3127
R83 VP.n34 VP.n33 11.3127
R84 VP.n45 VP.n44 1.96785
R85 VP.n75 VP.n74 1.96785
R86 VP.n41 VP.n40 1.96785
R87 VP.n19 VP.n16 0.189894
R88 VP.n23 VP.n16 0.189894
R89 VP.n24 VP.n23 0.189894
R90 VP.n25 VP.n24 0.189894
R91 VP.n25 VP.n14 0.189894
R92 VP.n29 VP.n14 0.189894
R93 VP.n30 VP.n29 0.189894
R94 VP.n31 VP.n30 0.189894
R95 VP.n31 VP.n12 0.189894
R96 VP.n36 VP.n12 0.189894
R97 VP.n37 VP.n36 0.189894
R98 VP.n38 VP.n37 0.189894
R99 VP.n38 VP.n10 0.189894
R100 VP.n42 VP.n10 0.189894
R101 VP.n46 VP.n43 0.189894
R102 VP.n47 VP.n46 0.189894
R103 VP.n48 VP.n47 0.189894
R104 VP.n48 VP.n8 0.189894
R105 VP.n52 VP.n8 0.189894
R106 VP.n53 VP.n52 0.189894
R107 VP.n53 VP.n6 0.189894
R108 VP.n57 VP.n6 0.189894
R109 VP.n58 VP.n57 0.189894
R110 VP.n59 VP.n58 0.189894
R111 VP.n59 VP.n4 0.189894
R112 VP.n63 VP.n4 0.189894
R113 VP.n64 VP.n63 0.189894
R114 VP.n65 VP.n64 0.189894
R115 VP.n65 VP.n2 0.189894
R116 VP.n70 VP.n2 0.189894
R117 VP.n71 VP.n70 0.189894
R118 VP.n72 VP.n71 0.189894
R119 VP.n72 VP.n0 0.189894
R120 VP.n76 VP.n0 0.189894
R121 VP VP.n76 0.0516364
R122 VTAIL.n11 VTAIL.t19 52.8323
R123 VTAIL.n17 VTAIL.t3 52.8321
R124 VTAIL.n2 VTAIL.t8 52.8321
R125 VTAIL.n16 VTAIL.t11 52.8321
R126 VTAIL.n15 VTAIL.n14 51.0083
R127 VTAIL.n13 VTAIL.n12 51.0083
R128 VTAIL.n10 VTAIL.n9 51.0083
R129 VTAIL.n8 VTAIL.n7 51.0083
R130 VTAIL.n19 VTAIL.n18 51.008
R131 VTAIL.n1 VTAIL.n0 51.008
R132 VTAIL.n4 VTAIL.n3 51.008
R133 VTAIL.n6 VTAIL.n5 51.008
R134 VTAIL.n8 VTAIL.n6 31.6427
R135 VTAIL.n17 VTAIL.n16 29.6858
R136 VTAIL.n10 VTAIL.n8 1.9574
R137 VTAIL.n11 VTAIL.n10 1.9574
R138 VTAIL.n15 VTAIL.n13 1.9574
R139 VTAIL.n16 VTAIL.n15 1.9574
R140 VTAIL.n6 VTAIL.n4 1.9574
R141 VTAIL.n4 VTAIL.n2 1.9574
R142 VTAIL.n19 VTAIL.n17 1.9574
R143 VTAIL.n18 VTAIL.t5 1.82457
R144 VTAIL.n18 VTAIL.t18 1.82457
R145 VTAIL.n0 VTAIL.t0 1.82457
R146 VTAIL.n0 VTAIL.t1 1.82457
R147 VTAIL.n3 VTAIL.t13 1.82457
R148 VTAIL.n3 VTAIL.t10 1.82457
R149 VTAIL.n5 VTAIL.t16 1.82457
R150 VTAIL.n5 VTAIL.t7 1.82457
R151 VTAIL.n14 VTAIL.t12 1.82457
R152 VTAIL.n14 VTAIL.t9 1.82457
R153 VTAIL.n12 VTAIL.t15 1.82457
R154 VTAIL.n12 VTAIL.t14 1.82457
R155 VTAIL.n9 VTAIL.t4 1.82457
R156 VTAIL.n9 VTAIL.t6 1.82457
R157 VTAIL.n7 VTAIL.t2 1.82457
R158 VTAIL.n7 VTAIL.t17 1.82457
R159 VTAIL VTAIL.n1 1.52636
R160 VTAIL.n13 VTAIL.n11 1.44878
R161 VTAIL.n2 VTAIL.n1 1.44878
R162 VTAIL VTAIL.n19 0.431534
R163 VDD1.n1 VDD1.t8 71.468
R164 VDD1.n3 VDD1.t9 71.4678
R165 VDD1.n5 VDD1.n4 69.0991
R166 VDD1.n1 VDD1.n0 67.6871
R167 VDD1.n7 VDD1.n6 67.6869
R168 VDD1.n3 VDD1.n2 67.6868
R169 VDD1.n7 VDD1.n5 49.9341
R170 VDD1.n6 VDD1.t1 1.82457
R171 VDD1.n6 VDD1.t7 1.82457
R172 VDD1.n0 VDD1.t5 1.82457
R173 VDD1.n0 VDD1.t3 1.82457
R174 VDD1.n4 VDD1.t6 1.82457
R175 VDD1.n4 VDD1.t0 1.82457
R176 VDD1.n2 VDD1.t2 1.82457
R177 VDD1.n2 VDD1.t4 1.82457
R178 VDD1 VDD1.n7 1.40998
R179 VDD1 VDD1.n1 0.547914
R180 VDD1.n5 VDD1.n3 0.434378
R181 B.n643 B.n642 585
R182 B.n644 B.n93 585
R183 B.n646 B.n645 585
R184 B.n647 B.n92 585
R185 B.n649 B.n648 585
R186 B.n650 B.n91 585
R187 B.n652 B.n651 585
R188 B.n653 B.n90 585
R189 B.n655 B.n654 585
R190 B.n656 B.n89 585
R191 B.n658 B.n657 585
R192 B.n659 B.n88 585
R193 B.n661 B.n660 585
R194 B.n662 B.n87 585
R195 B.n664 B.n663 585
R196 B.n665 B.n86 585
R197 B.n667 B.n666 585
R198 B.n668 B.n85 585
R199 B.n670 B.n669 585
R200 B.n671 B.n84 585
R201 B.n673 B.n672 585
R202 B.n674 B.n83 585
R203 B.n676 B.n675 585
R204 B.n677 B.n82 585
R205 B.n679 B.n678 585
R206 B.n680 B.n81 585
R207 B.n682 B.n681 585
R208 B.n683 B.n80 585
R209 B.n685 B.n684 585
R210 B.n686 B.n79 585
R211 B.n688 B.n687 585
R212 B.n689 B.n78 585
R213 B.n691 B.n690 585
R214 B.n692 B.n77 585
R215 B.n694 B.n693 585
R216 B.n695 B.n76 585
R217 B.n697 B.n696 585
R218 B.n698 B.n75 585
R219 B.n700 B.n699 585
R220 B.n701 B.n74 585
R221 B.n703 B.n702 585
R222 B.n704 B.n73 585
R223 B.n706 B.n705 585
R224 B.n707 B.n72 585
R225 B.n709 B.n708 585
R226 B.n710 B.n71 585
R227 B.n712 B.n711 585
R228 B.n713 B.n70 585
R229 B.n715 B.n714 585
R230 B.n716 B.n69 585
R231 B.n718 B.n717 585
R232 B.n719 B.n68 585
R233 B.n721 B.n720 585
R234 B.n722 B.n67 585
R235 B.n724 B.n723 585
R236 B.n725 B.n66 585
R237 B.n727 B.n726 585
R238 B.n728 B.n65 585
R239 B.n730 B.n729 585
R240 B.n732 B.n731 585
R241 B.n733 B.n61 585
R242 B.n735 B.n734 585
R243 B.n736 B.n60 585
R244 B.n738 B.n737 585
R245 B.n739 B.n59 585
R246 B.n741 B.n740 585
R247 B.n742 B.n58 585
R248 B.n744 B.n743 585
R249 B.n746 B.n55 585
R250 B.n748 B.n747 585
R251 B.n749 B.n54 585
R252 B.n751 B.n750 585
R253 B.n752 B.n53 585
R254 B.n754 B.n753 585
R255 B.n755 B.n52 585
R256 B.n757 B.n756 585
R257 B.n758 B.n51 585
R258 B.n760 B.n759 585
R259 B.n761 B.n50 585
R260 B.n763 B.n762 585
R261 B.n764 B.n49 585
R262 B.n766 B.n765 585
R263 B.n767 B.n48 585
R264 B.n769 B.n768 585
R265 B.n770 B.n47 585
R266 B.n772 B.n771 585
R267 B.n773 B.n46 585
R268 B.n775 B.n774 585
R269 B.n776 B.n45 585
R270 B.n778 B.n777 585
R271 B.n779 B.n44 585
R272 B.n781 B.n780 585
R273 B.n782 B.n43 585
R274 B.n784 B.n783 585
R275 B.n785 B.n42 585
R276 B.n787 B.n786 585
R277 B.n788 B.n41 585
R278 B.n790 B.n789 585
R279 B.n791 B.n40 585
R280 B.n793 B.n792 585
R281 B.n794 B.n39 585
R282 B.n796 B.n795 585
R283 B.n797 B.n38 585
R284 B.n799 B.n798 585
R285 B.n800 B.n37 585
R286 B.n802 B.n801 585
R287 B.n803 B.n36 585
R288 B.n805 B.n804 585
R289 B.n806 B.n35 585
R290 B.n808 B.n807 585
R291 B.n809 B.n34 585
R292 B.n811 B.n810 585
R293 B.n812 B.n33 585
R294 B.n814 B.n813 585
R295 B.n815 B.n32 585
R296 B.n817 B.n816 585
R297 B.n818 B.n31 585
R298 B.n820 B.n819 585
R299 B.n821 B.n30 585
R300 B.n823 B.n822 585
R301 B.n824 B.n29 585
R302 B.n826 B.n825 585
R303 B.n827 B.n28 585
R304 B.n829 B.n828 585
R305 B.n830 B.n27 585
R306 B.n832 B.n831 585
R307 B.n833 B.n26 585
R308 B.n641 B.n94 585
R309 B.n640 B.n639 585
R310 B.n638 B.n95 585
R311 B.n637 B.n636 585
R312 B.n635 B.n96 585
R313 B.n634 B.n633 585
R314 B.n632 B.n97 585
R315 B.n631 B.n630 585
R316 B.n629 B.n98 585
R317 B.n628 B.n627 585
R318 B.n626 B.n99 585
R319 B.n625 B.n624 585
R320 B.n623 B.n100 585
R321 B.n622 B.n621 585
R322 B.n620 B.n101 585
R323 B.n619 B.n618 585
R324 B.n617 B.n102 585
R325 B.n616 B.n615 585
R326 B.n614 B.n103 585
R327 B.n613 B.n612 585
R328 B.n611 B.n104 585
R329 B.n610 B.n609 585
R330 B.n608 B.n105 585
R331 B.n607 B.n606 585
R332 B.n605 B.n106 585
R333 B.n604 B.n603 585
R334 B.n602 B.n107 585
R335 B.n601 B.n600 585
R336 B.n599 B.n108 585
R337 B.n598 B.n597 585
R338 B.n596 B.n109 585
R339 B.n595 B.n594 585
R340 B.n593 B.n110 585
R341 B.n592 B.n591 585
R342 B.n590 B.n111 585
R343 B.n589 B.n588 585
R344 B.n587 B.n112 585
R345 B.n586 B.n585 585
R346 B.n584 B.n113 585
R347 B.n583 B.n582 585
R348 B.n581 B.n114 585
R349 B.n580 B.n579 585
R350 B.n578 B.n115 585
R351 B.n577 B.n576 585
R352 B.n575 B.n116 585
R353 B.n574 B.n573 585
R354 B.n572 B.n117 585
R355 B.n571 B.n570 585
R356 B.n569 B.n118 585
R357 B.n568 B.n567 585
R358 B.n566 B.n119 585
R359 B.n565 B.n564 585
R360 B.n563 B.n120 585
R361 B.n562 B.n561 585
R362 B.n560 B.n121 585
R363 B.n559 B.n558 585
R364 B.n557 B.n122 585
R365 B.n556 B.n555 585
R366 B.n554 B.n123 585
R367 B.n553 B.n552 585
R368 B.n551 B.n124 585
R369 B.n550 B.n549 585
R370 B.n548 B.n125 585
R371 B.n547 B.n546 585
R372 B.n545 B.n126 585
R373 B.n544 B.n543 585
R374 B.n542 B.n127 585
R375 B.n541 B.n540 585
R376 B.n539 B.n128 585
R377 B.n538 B.n537 585
R378 B.n536 B.n129 585
R379 B.n535 B.n534 585
R380 B.n533 B.n130 585
R381 B.n532 B.n531 585
R382 B.n530 B.n131 585
R383 B.n529 B.n528 585
R384 B.n527 B.n132 585
R385 B.n526 B.n525 585
R386 B.n524 B.n133 585
R387 B.n523 B.n522 585
R388 B.n521 B.n134 585
R389 B.n520 B.n519 585
R390 B.n518 B.n135 585
R391 B.n517 B.n516 585
R392 B.n515 B.n136 585
R393 B.n514 B.n513 585
R394 B.n512 B.n137 585
R395 B.n511 B.n510 585
R396 B.n509 B.n138 585
R397 B.n508 B.n507 585
R398 B.n506 B.n139 585
R399 B.n505 B.n504 585
R400 B.n503 B.n140 585
R401 B.n502 B.n501 585
R402 B.n500 B.n141 585
R403 B.n499 B.n498 585
R404 B.n497 B.n142 585
R405 B.n305 B.n210 585
R406 B.n307 B.n306 585
R407 B.n308 B.n209 585
R408 B.n310 B.n309 585
R409 B.n311 B.n208 585
R410 B.n313 B.n312 585
R411 B.n314 B.n207 585
R412 B.n316 B.n315 585
R413 B.n317 B.n206 585
R414 B.n319 B.n318 585
R415 B.n320 B.n205 585
R416 B.n322 B.n321 585
R417 B.n323 B.n204 585
R418 B.n325 B.n324 585
R419 B.n326 B.n203 585
R420 B.n328 B.n327 585
R421 B.n329 B.n202 585
R422 B.n331 B.n330 585
R423 B.n332 B.n201 585
R424 B.n334 B.n333 585
R425 B.n335 B.n200 585
R426 B.n337 B.n336 585
R427 B.n338 B.n199 585
R428 B.n340 B.n339 585
R429 B.n341 B.n198 585
R430 B.n343 B.n342 585
R431 B.n344 B.n197 585
R432 B.n346 B.n345 585
R433 B.n347 B.n196 585
R434 B.n349 B.n348 585
R435 B.n350 B.n195 585
R436 B.n352 B.n351 585
R437 B.n353 B.n194 585
R438 B.n355 B.n354 585
R439 B.n356 B.n193 585
R440 B.n358 B.n357 585
R441 B.n359 B.n192 585
R442 B.n361 B.n360 585
R443 B.n362 B.n191 585
R444 B.n364 B.n363 585
R445 B.n365 B.n190 585
R446 B.n367 B.n366 585
R447 B.n368 B.n189 585
R448 B.n370 B.n369 585
R449 B.n371 B.n188 585
R450 B.n373 B.n372 585
R451 B.n374 B.n187 585
R452 B.n376 B.n375 585
R453 B.n377 B.n186 585
R454 B.n379 B.n378 585
R455 B.n380 B.n185 585
R456 B.n382 B.n381 585
R457 B.n383 B.n184 585
R458 B.n385 B.n384 585
R459 B.n386 B.n183 585
R460 B.n388 B.n387 585
R461 B.n389 B.n182 585
R462 B.n391 B.n390 585
R463 B.n392 B.n179 585
R464 B.n395 B.n394 585
R465 B.n396 B.n178 585
R466 B.n398 B.n397 585
R467 B.n399 B.n177 585
R468 B.n401 B.n400 585
R469 B.n402 B.n176 585
R470 B.n404 B.n403 585
R471 B.n405 B.n175 585
R472 B.n407 B.n406 585
R473 B.n409 B.n408 585
R474 B.n410 B.n171 585
R475 B.n412 B.n411 585
R476 B.n413 B.n170 585
R477 B.n415 B.n414 585
R478 B.n416 B.n169 585
R479 B.n418 B.n417 585
R480 B.n419 B.n168 585
R481 B.n421 B.n420 585
R482 B.n422 B.n167 585
R483 B.n424 B.n423 585
R484 B.n425 B.n166 585
R485 B.n427 B.n426 585
R486 B.n428 B.n165 585
R487 B.n430 B.n429 585
R488 B.n431 B.n164 585
R489 B.n433 B.n432 585
R490 B.n434 B.n163 585
R491 B.n436 B.n435 585
R492 B.n437 B.n162 585
R493 B.n439 B.n438 585
R494 B.n440 B.n161 585
R495 B.n442 B.n441 585
R496 B.n443 B.n160 585
R497 B.n445 B.n444 585
R498 B.n446 B.n159 585
R499 B.n448 B.n447 585
R500 B.n449 B.n158 585
R501 B.n451 B.n450 585
R502 B.n452 B.n157 585
R503 B.n454 B.n453 585
R504 B.n455 B.n156 585
R505 B.n457 B.n456 585
R506 B.n458 B.n155 585
R507 B.n460 B.n459 585
R508 B.n461 B.n154 585
R509 B.n463 B.n462 585
R510 B.n464 B.n153 585
R511 B.n466 B.n465 585
R512 B.n467 B.n152 585
R513 B.n469 B.n468 585
R514 B.n470 B.n151 585
R515 B.n472 B.n471 585
R516 B.n473 B.n150 585
R517 B.n475 B.n474 585
R518 B.n476 B.n149 585
R519 B.n478 B.n477 585
R520 B.n479 B.n148 585
R521 B.n481 B.n480 585
R522 B.n482 B.n147 585
R523 B.n484 B.n483 585
R524 B.n485 B.n146 585
R525 B.n487 B.n486 585
R526 B.n488 B.n145 585
R527 B.n490 B.n489 585
R528 B.n491 B.n144 585
R529 B.n493 B.n492 585
R530 B.n494 B.n143 585
R531 B.n496 B.n495 585
R532 B.n304 B.n303 585
R533 B.n302 B.n211 585
R534 B.n301 B.n300 585
R535 B.n299 B.n212 585
R536 B.n298 B.n297 585
R537 B.n296 B.n213 585
R538 B.n295 B.n294 585
R539 B.n293 B.n214 585
R540 B.n292 B.n291 585
R541 B.n290 B.n215 585
R542 B.n289 B.n288 585
R543 B.n287 B.n216 585
R544 B.n286 B.n285 585
R545 B.n284 B.n217 585
R546 B.n283 B.n282 585
R547 B.n281 B.n218 585
R548 B.n280 B.n279 585
R549 B.n278 B.n219 585
R550 B.n277 B.n276 585
R551 B.n275 B.n220 585
R552 B.n274 B.n273 585
R553 B.n272 B.n221 585
R554 B.n271 B.n270 585
R555 B.n269 B.n222 585
R556 B.n268 B.n267 585
R557 B.n266 B.n223 585
R558 B.n265 B.n264 585
R559 B.n263 B.n224 585
R560 B.n262 B.n261 585
R561 B.n260 B.n225 585
R562 B.n259 B.n258 585
R563 B.n257 B.n226 585
R564 B.n256 B.n255 585
R565 B.n254 B.n227 585
R566 B.n253 B.n252 585
R567 B.n251 B.n228 585
R568 B.n250 B.n249 585
R569 B.n248 B.n229 585
R570 B.n247 B.n246 585
R571 B.n245 B.n230 585
R572 B.n244 B.n243 585
R573 B.n242 B.n231 585
R574 B.n241 B.n240 585
R575 B.n239 B.n232 585
R576 B.n238 B.n237 585
R577 B.n236 B.n233 585
R578 B.n235 B.n234 585
R579 B.n2 B.n0 585
R580 B.n905 B.n1 585
R581 B.n904 B.n903 585
R582 B.n902 B.n3 585
R583 B.n901 B.n900 585
R584 B.n899 B.n4 585
R585 B.n898 B.n897 585
R586 B.n896 B.n5 585
R587 B.n895 B.n894 585
R588 B.n893 B.n6 585
R589 B.n892 B.n891 585
R590 B.n890 B.n7 585
R591 B.n889 B.n888 585
R592 B.n887 B.n8 585
R593 B.n886 B.n885 585
R594 B.n884 B.n9 585
R595 B.n883 B.n882 585
R596 B.n881 B.n10 585
R597 B.n880 B.n879 585
R598 B.n878 B.n11 585
R599 B.n877 B.n876 585
R600 B.n875 B.n12 585
R601 B.n874 B.n873 585
R602 B.n872 B.n13 585
R603 B.n871 B.n870 585
R604 B.n869 B.n14 585
R605 B.n868 B.n867 585
R606 B.n866 B.n15 585
R607 B.n865 B.n864 585
R608 B.n863 B.n16 585
R609 B.n862 B.n861 585
R610 B.n860 B.n17 585
R611 B.n859 B.n858 585
R612 B.n857 B.n18 585
R613 B.n856 B.n855 585
R614 B.n854 B.n19 585
R615 B.n853 B.n852 585
R616 B.n851 B.n20 585
R617 B.n850 B.n849 585
R618 B.n848 B.n21 585
R619 B.n847 B.n846 585
R620 B.n845 B.n22 585
R621 B.n844 B.n843 585
R622 B.n842 B.n23 585
R623 B.n841 B.n840 585
R624 B.n839 B.n24 585
R625 B.n838 B.n837 585
R626 B.n836 B.n25 585
R627 B.n835 B.n834 585
R628 B.n907 B.n906 585
R629 B.n305 B.n304 530.939
R630 B.n834 B.n833 530.939
R631 B.n497 B.n496 530.939
R632 B.n642 B.n641 530.939
R633 B.n172 B.t9 428.146
R634 B.n180 B.t3 428.146
R635 B.n56 B.t0 428.146
R636 B.n62 B.t6 428.146
R637 B.n304 B.n211 163.367
R638 B.n300 B.n211 163.367
R639 B.n300 B.n299 163.367
R640 B.n299 B.n298 163.367
R641 B.n298 B.n213 163.367
R642 B.n294 B.n213 163.367
R643 B.n294 B.n293 163.367
R644 B.n293 B.n292 163.367
R645 B.n292 B.n215 163.367
R646 B.n288 B.n215 163.367
R647 B.n288 B.n287 163.367
R648 B.n287 B.n286 163.367
R649 B.n286 B.n217 163.367
R650 B.n282 B.n217 163.367
R651 B.n282 B.n281 163.367
R652 B.n281 B.n280 163.367
R653 B.n280 B.n219 163.367
R654 B.n276 B.n219 163.367
R655 B.n276 B.n275 163.367
R656 B.n275 B.n274 163.367
R657 B.n274 B.n221 163.367
R658 B.n270 B.n221 163.367
R659 B.n270 B.n269 163.367
R660 B.n269 B.n268 163.367
R661 B.n268 B.n223 163.367
R662 B.n264 B.n223 163.367
R663 B.n264 B.n263 163.367
R664 B.n263 B.n262 163.367
R665 B.n262 B.n225 163.367
R666 B.n258 B.n225 163.367
R667 B.n258 B.n257 163.367
R668 B.n257 B.n256 163.367
R669 B.n256 B.n227 163.367
R670 B.n252 B.n227 163.367
R671 B.n252 B.n251 163.367
R672 B.n251 B.n250 163.367
R673 B.n250 B.n229 163.367
R674 B.n246 B.n229 163.367
R675 B.n246 B.n245 163.367
R676 B.n245 B.n244 163.367
R677 B.n244 B.n231 163.367
R678 B.n240 B.n231 163.367
R679 B.n240 B.n239 163.367
R680 B.n239 B.n238 163.367
R681 B.n238 B.n233 163.367
R682 B.n234 B.n233 163.367
R683 B.n234 B.n2 163.367
R684 B.n906 B.n2 163.367
R685 B.n906 B.n905 163.367
R686 B.n905 B.n904 163.367
R687 B.n904 B.n3 163.367
R688 B.n900 B.n3 163.367
R689 B.n900 B.n899 163.367
R690 B.n899 B.n898 163.367
R691 B.n898 B.n5 163.367
R692 B.n894 B.n5 163.367
R693 B.n894 B.n893 163.367
R694 B.n893 B.n892 163.367
R695 B.n892 B.n7 163.367
R696 B.n888 B.n7 163.367
R697 B.n888 B.n887 163.367
R698 B.n887 B.n886 163.367
R699 B.n886 B.n9 163.367
R700 B.n882 B.n9 163.367
R701 B.n882 B.n881 163.367
R702 B.n881 B.n880 163.367
R703 B.n880 B.n11 163.367
R704 B.n876 B.n11 163.367
R705 B.n876 B.n875 163.367
R706 B.n875 B.n874 163.367
R707 B.n874 B.n13 163.367
R708 B.n870 B.n13 163.367
R709 B.n870 B.n869 163.367
R710 B.n869 B.n868 163.367
R711 B.n868 B.n15 163.367
R712 B.n864 B.n15 163.367
R713 B.n864 B.n863 163.367
R714 B.n863 B.n862 163.367
R715 B.n862 B.n17 163.367
R716 B.n858 B.n17 163.367
R717 B.n858 B.n857 163.367
R718 B.n857 B.n856 163.367
R719 B.n856 B.n19 163.367
R720 B.n852 B.n19 163.367
R721 B.n852 B.n851 163.367
R722 B.n851 B.n850 163.367
R723 B.n850 B.n21 163.367
R724 B.n846 B.n21 163.367
R725 B.n846 B.n845 163.367
R726 B.n845 B.n844 163.367
R727 B.n844 B.n23 163.367
R728 B.n840 B.n23 163.367
R729 B.n840 B.n839 163.367
R730 B.n839 B.n838 163.367
R731 B.n838 B.n25 163.367
R732 B.n834 B.n25 163.367
R733 B.n306 B.n305 163.367
R734 B.n306 B.n209 163.367
R735 B.n310 B.n209 163.367
R736 B.n311 B.n310 163.367
R737 B.n312 B.n311 163.367
R738 B.n312 B.n207 163.367
R739 B.n316 B.n207 163.367
R740 B.n317 B.n316 163.367
R741 B.n318 B.n317 163.367
R742 B.n318 B.n205 163.367
R743 B.n322 B.n205 163.367
R744 B.n323 B.n322 163.367
R745 B.n324 B.n323 163.367
R746 B.n324 B.n203 163.367
R747 B.n328 B.n203 163.367
R748 B.n329 B.n328 163.367
R749 B.n330 B.n329 163.367
R750 B.n330 B.n201 163.367
R751 B.n334 B.n201 163.367
R752 B.n335 B.n334 163.367
R753 B.n336 B.n335 163.367
R754 B.n336 B.n199 163.367
R755 B.n340 B.n199 163.367
R756 B.n341 B.n340 163.367
R757 B.n342 B.n341 163.367
R758 B.n342 B.n197 163.367
R759 B.n346 B.n197 163.367
R760 B.n347 B.n346 163.367
R761 B.n348 B.n347 163.367
R762 B.n348 B.n195 163.367
R763 B.n352 B.n195 163.367
R764 B.n353 B.n352 163.367
R765 B.n354 B.n353 163.367
R766 B.n354 B.n193 163.367
R767 B.n358 B.n193 163.367
R768 B.n359 B.n358 163.367
R769 B.n360 B.n359 163.367
R770 B.n360 B.n191 163.367
R771 B.n364 B.n191 163.367
R772 B.n365 B.n364 163.367
R773 B.n366 B.n365 163.367
R774 B.n366 B.n189 163.367
R775 B.n370 B.n189 163.367
R776 B.n371 B.n370 163.367
R777 B.n372 B.n371 163.367
R778 B.n372 B.n187 163.367
R779 B.n376 B.n187 163.367
R780 B.n377 B.n376 163.367
R781 B.n378 B.n377 163.367
R782 B.n378 B.n185 163.367
R783 B.n382 B.n185 163.367
R784 B.n383 B.n382 163.367
R785 B.n384 B.n383 163.367
R786 B.n384 B.n183 163.367
R787 B.n388 B.n183 163.367
R788 B.n389 B.n388 163.367
R789 B.n390 B.n389 163.367
R790 B.n390 B.n179 163.367
R791 B.n395 B.n179 163.367
R792 B.n396 B.n395 163.367
R793 B.n397 B.n396 163.367
R794 B.n397 B.n177 163.367
R795 B.n401 B.n177 163.367
R796 B.n402 B.n401 163.367
R797 B.n403 B.n402 163.367
R798 B.n403 B.n175 163.367
R799 B.n407 B.n175 163.367
R800 B.n408 B.n407 163.367
R801 B.n408 B.n171 163.367
R802 B.n412 B.n171 163.367
R803 B.n413 B.n412 163.367
R804 B.n414 B.n413 163.367
R805 B.n414 B.n169 163.367
R806 B.n418 B.n169 163.367
R807 B.n419 B.n418 163.367
R808 B.n420 B.n419 163.367
R809 B.n420 B.n167 163.367
R810 B.n424 B.n167 163.367
R811 B.n425 B.n424 163.367
R812 B.n426 B.n425 163.367
R813 B.n426 B.n165 163.367
R814 B.n430 B.n165 163.367
R815 B.n431 B.n430 163.367
R816 B.n432 B.n431 163.367
R817 B.n432 B.n163 163.367
R818 B.n436 B.n163 163.367
R819 B.n437 B.n436 163.367
R820 B.n438 B.n437 163.367
R821 B.n438 B.n161 163.367
R822 B.n442 B.n161 163.367
R823 B.n443 B.n442 163.367
R824 B.n444 B.n443 163.367
R825 B.n444 B.n159 163.367
R826 B.n448 B.n159 163.367
R827 B.n449 B.n448 163.367
R828 B.n450 B.n449 163.367
R829 B.n450 B.n157 163.367
R830 B.n454 B.n157 163.367
R831 B.n455 B.n454 163.367
R832 B.n456 B.n455 163.367
R833 B.n456 B.n155 163.367
R834 B.n460 B.n155 163.367
R835 B.n461 B.n460 163.367
R836 B.n462 B.n461 163.367
R837 B.n462 B.n153 163.367
R838 B.n466 B.n153 163.367
R839 B.n467 B.n466 163.367
R840 B.n468 B.n467 163.367
R841 B.n468 B.n151 163.367
R842 B.n472 B.n151 163.367
R843 B.n473 B.n472 163.367
R844 B.n474 B.n473 163.367
R845 B.n474 B.n149 163.367
R846 B.n478 B.n149 163.367
R847 B.n479 B.n478 163.367
R848 B.n480 B.n479 163.367
R849 B.n480 B.n147 163.367
R850 B.n484 B.n147 163.367
R851 B.n485 B.n484 163.367
R852 B.n486 B.n485 163.367
R853 B.n486 B.n145 163.367
R854 B.n490 B.n145 163.367
R855 B.n491 B.n490 163.367
R856 B.n492 B.n491 163.367
R857 B.n492 B.n143 163.367
R858 B.n496 B.n143 163.367
R859 B.n498 B.n497 163.367
R860 B.n498 B.n141 163.367
R861 B.n502 B.n141 163.367
R862 B.n503 B.n502 163.367
R863 B.n504 B.n503 163.367
R864 B.n504 B.n139 163.367
R865 B.n508 B.n139 163.367
R866 B.n509 B.n508 163.367
R867 B.n510 B.n509 163.367
R868 B.n510 B.n137 163.367
R869 B.n514 B.n137 163.367
R870 B.n515 B.n514 163.367
R871 B.n516 B.n515 163.367
R872 B.n516 B.n135 163.367
R873 B.n520 B.n135 163.367
R874 B.n521 B.n520 163.367
R875 B.n522 B.n521 163.367
R876 B.n522 B.n133 163.367
R877 B.n526 B.n133 163.367
R878 B.n527 B.n526 163.367
R879 B.n528 B.n527 163.367
R880 B.n528 B.n131 163.367
R881 B.n532 B.n131 163.367
R882 B.n533 B.n532 163.367
R883 B.n534 B.n533 163.367
R884 B.n534 B.n129 163.367
R885 B.n538 B.n129 163.367
R886 B.n539 B.n538 163.367
R887 B.n540 B.n539 163.367
R888 B.n540 B.n127 163.367
R889 B.n544 B.n127 163.367
R890 B.n545 B.n544 163.367
R891 B.n546 B.n545 163.367
R892 B.n546 B.n125 163.367
R893 B.n550 B.n125 163.367
R894 B.n551 B.n550 163.367
R895 B.n552 B.n551 163.367
R896 B.n552 B.n123 163.367
R897 B.n556 B.n123 163.367
R898 B.n557 B.n556 163.367
R899 B.n558 B.n557 163.367
R900 B.n558 B.n121 163.367
R901 B.n562 B.n121 163.367
R902 B.n563 B.n562 163.367
R903 B.n564 B.n563 163.367
R904 B.n564 B.n119 163.367
R905 B.n568 B.n119 163.367
R906 B.n569 B.n568 163.367
R907 B.n570 B.n569 163.367
R908 B.n570 B.n117 163.367
R909 B.n574 B.n117 163.367
R910 B.n575 B.n574 163.367
R911 B.n576 B.n575 163.367
R912 B.n576 B.n115 163.367
R913 B.n580 B.n115 163.367
R914 B.n581 B.n580 163.367
R915 B.n582 B.n581 163.367
R916 B.n582 B.n113 163.367
R917 B.n586 B.n113 163.367
R918 B.n587 B.n586 163.367
R919 B.n588 B.n587 163.367
R920 B.n588 B.n111 163.367
R921 B.n592 B.n111 163.367
R922 B.n593 B.n592 163.367
R923 B.n594 B.n593 163.367
R924 B.n594 B.n109 163.367
R925 B.n598 B.n109 163.367
R926 B.n599 B.n598 163.367
R927 B.n600 B.n599 163.367
R928 B.n600 B.n107 163.367
R929 B.n604 B.n107 163.367
R930 B.n605 B.n604 163.367
R931 B.n606 B.n605 163.367
R932 B.n606 B.n105 163.367
R933 B.n610 B.n105 163.367
R934 B.n611 B.n610 163.367
R935 B.n612 B.n611 163.367
R936 B.n612 B.n103 163.367
R937 B.n616 B.n103 163.367
R938 B.n617 B.n616 163.367
R939 B.n618 B.n617 163.367
R940 B.n618 B.n101 163.367
R941 B.n622 B.n101 163.367
R942 B.n623 B.n622 163.367
R943 B.n624 B.n623 163.367
R944 B.n624 B.n99 163.367
R945 B.n628 B.n99 163.367
R946 B.n629 B.n628 163.367
R947 B.n630 B.n629 163.367
R948 B.n630 B.n97 163.367
R949 B.n634 B.n97 163.367
R950 B.n635 B.n634 163.367
R951 B.n636 B.n635 163.367
R952 B.n636 B.n95 163.367
R953 B.n640 B.n95 163.367
R954 B.n641 B.n640 163.367
R955 B.n833 B.n832 163.367
R956 B.n832 B.n27 163.367
R957 B.n828 B.n27 163.367
R958 B.n828 B.n827 163.367
R959 B.n827 B.n826 163.367
R960 B.n826 B.n29 163.367
R961 B.n822 B.n29 163.367
R962 B.n822 B.n821 163.367
R963 B.n821 B.n820 163.367
R964 B.n820 B.n31 163.367
R965 B.n816 B.n31 163.367
R966 B.n816 B.n815 163.367
R967 B.n815 B.n814 163.367
R968 B.n814 B.n33 163.367
R969 B.n810 B.n33 163.367
R970 B.n810 B.n809 163.367
R971 B.n809 B.n808 163.367
R972 B.n808 B.n35 163.367
R973 B.n804 B.n35 163.367
R974 B.n804 B.n803 163.367
R975 B.n803 B.n802 163.367
R976 B.n802 B.n37 163.367
R977 B.n798 B.n37 163.367
R978 B.n798 B.n797 163.367
R979 B.n797 B.n796 163.367
R980 B.n796 B.n39 163.367
R981 B.n792 B.n39 163.367
R982 B.n792 B.n791 163.367
R983 B.n791 B.n790 163.367
R984 B.n790 B.n41 163.367
R985 B.n786 B.n41 163.367
R986 B.n786 B.n785 163.367
R987 B.n785 B.n784 163.367
R988 B.n784 B.n43 163.367
R989 B.n780 B.n43 163.367
R990 B.n780 B.n779 163.367
R991 B.n779 B.n778 163.367
R992 B.n778 B.n45 163.367
R993 B.n774 B.n45 163.367
R994 B.n774 B.n773 163.367
R995 B.n773 B.n772 163.367
R996 B.n772 B.n47 163.367
R997 B.n768 B.n47 163.367
R998 B.n768 B.n767 163.367
R999 B.n767 B.n766 163.367
R1000 B.n766 B.n49 163.367
R1001 B.n762 B.n49 163.367
R1002 B.n762 B.n761 163.367
R1003 B.n761 B.n760 163.367
R1004 B.n760 B.n51 163.367
R1005 B.n756 B.n51 163.367
R1006 B.n756 B.n755 163.367
R1007 B.n755 B.n754 163.367
R1008 B.n754 B.n53 163.367
R1009 B.n750 B.n53 163.367
R1010 B.n750 B.n749 163.367
R1011 B.n749 B.n748 163.367
R1012 B.n748 B.n55 163.367
R1013 B.n743 B.n55 163.367
R1014 B.n743 B.n742 163.367
R1015 B.n742 B.n741 163.367
R1016 B.n741 B.n59 163.367
R1017 B.n737 B.n59 163.367
R1018 B.n737 B.n736 163.367
R1019 B.n736 B.n735 163.367
R1020 B.n735 B.n61 163.367
R1021 B.n731 B.n61 163.367
R1022 B.n731 B.n730 163.367
R1023 B.n730 B.n65 163.367
R1024 B.n726 B.n65 163.367
R1025 B.n726 B.n725 163.367
R1026 B.n725 B.n724 163.367
R1027 B.n724 B.n67 163.367
R1028 B.n720 B.n67 163.367
R1029 B.n720 B.n719 163.367
R1030 B.n719 B.n718 163.367
R1031 B.n718 B.n69 163.367
R1032 B.n714 B.n69 163.367
R1033 B.n714 B.n713 163.367
R1034 B.n713 B.n712 163.367
R1035 B.n712 B.n71 163.367
R1036 B.n708 B.n71 163.367
R1037 B.n708 B.n707 163.367
R1038 B.n707 B.n706 163.367
R1039 B.n706 B.n73 163.367
R1040 B.n702 B.n73 163.367
R1041 B.n702 B.n701 163.367
R1042 B.n701 B.n700 163.367
R1043 B.n700 B.n75 163.367
R1044 B.n696 B.n75 163.367
R1045 B.n696 B.n695 163.367
R1046 B.n695 B.n694 163.367
R1047 B.n694 B.n77 163.367
R1048 B.n690 B.n77 163.367
R1049 B.n690 B.n689 163.367
R1050 B.n689 B.n688 163.367
R1051 B.n688 B.n79 163.367
R1052 B.n684 B.n79 163.367
R1053 B.n684 B.n683 163.367
R1054 B.n683 B.n682 163.367
R1055 B.n682 B.n81 163.367
R1056 B.n678 B.n81 163.367
R1057 B.n678 B.n677 163.367
R1058 B.n677 B.n676 163.367
R1059 B.n676 B.n83 163.367
R1060 B.n672 B.n83 163.367
R1061 B.n672 B.n671 163.367
R1062 B.n671 B.n670 163.367
R1063 B.n670 B.n85 163.367
R1064 B.n666 B.n85 163.367
R1065 B.n666 B.n665 163.367
R1066 B.n665 B.n664 163.367
R1067 B.n664 B.n87 163.367
R1068 B.n660 B.n87 163.367
R1069 B.n660 B.n659 163.367
R1070 B.n659 B.n658 163.367
R1071 B.n658 B.n89 163.367
R1072 B.n654 B.n89 163.367
R1073 B.n654 B.n653 163.367
R1074 B.n653 B.n652 163.367
R1075 B.n652 B.n91 163.367
R1076 B.n648 B.n91 163.367
R1077 B.n648 B.n647 163.367
R1078 B.n647 B.n646 163.367
R1079 B.n646 B.n93 163.367
R1080 B.n642 B.n93 163.367
R1081 B.n172 B.t11 152.962
R1082 B.n62 B.t7 152.962
R1083 B.n180 B.t5 152.939
R1084 B.n56 B.t1 152.939
R1085 B.n173 B.t10 108.938
R1086 B.n63 B.t8 108.938
R1087 B.n181 B.t4 108.915
R1088 B.n57 B.t2 108.915
R1089 B.n174 B.n173 59.5399
R1090 B.n393 B.n181 59.5399
R1091 B.n745 B.n57 59.5399
R1092 B.n64 B.n63 59.5399
R1093 B.n173 B.n172 44.0247
R1094 B.n181 B.n180 44.0247
R1095 B.n57 B.n56 44.0247
R1096 B.n63 B.n62 44.0247
R1097 B.n835 B.n26 34.4981
R1098 B.n643 B.n94 34.4981
R1099 B.n495 B.n142 34.4981
R1100 B.n303 B.n210 34.4981
R1101 B B.n907 18.0485
R1102 B.n831 B.n26 10.6151
R1103 B.n831 B.n830 10.6151
R1104 B.n830 B.n829 10.6151
R1105 B.n829 B.n28 10.6151
R1106 B.n825 B.n28 10.6151
R1107 B.n825 B.n824 10.6151
R1108 B.n824 B.n823 10.6151
R1109 B.n823 B.n30 10.6151
R1110 B.n819 B.n30 10.6151
R1111 B.n819 B.n818 10.6151
R1112 B.n818 B.n817 10.6151
R1113 B.n817 B.n32 10.6151
R1114 B.n813 B.n32 10.6151
R1115 B.n813 B.n812 10.6151
R1116 B.n812 B.n811 10.6151
R1117 B.n811 B.n34 10.6151
R1118 B.n807 B.n34 10.6151
R1119 B.n807 B.n806 10.6151
R1120 B.n806 B.n805 10.6151
R1121 B.n805 B.n36 10.6151
R1122 B.n801 B.n36 10.6151
R1123 B.n801 B.n800 10.6151
R1124 B.n800 B.n799 10.6151
R1125 B.n799 B.n38 10.6151
R1126 B.n795 B.n38 10.6151
R1127 B.n795 B.n794 10.6151
R1128 B.n794 B.n793 10.6151
R1129 B.n793 B.n40 10.6151
R1130 B.n789 B.n40 10.6151
R1131 B.n789 B.n788 10.6151
R1132 B.n788 B.n787 10.6151
R1133 B.n787 B.n42 10.6151
R1134 B.n783 B.n42 10.6151
R1135 B.n783 B.n782 10.6151
R1136 B.n782 B.n781 10.6151
R1137 B.n781 B.n44 10.6151
R1138 B.n777 B.n44 10.6151
R1139 B.n777 B.n776 10.6151
R1140 B.n776 B.n775 10.6151
R1141 B.n775 B.n46 10.6151
R1142 B.n771 B.n46 10.6151
R1143 B.n771 B.n770 10.6151
R1144 B.n770 B.n769 10.6151
R1145 B.n769 B.n48 10.6151
R1146 B.n765 B.n48 10.6151
R1147 B.n765 B.n764 10.6151
R1148 B.n764 B.n763 10.6151
R1149 B.n763 B.n50 10.6151
R1150 B.n759 B.n50 10.6151
R1151 B.n759 B.n758 10.6151
R1152 B.n758 B.n757 10.6151
R1153 B.n757 B.n52 10.6151
R1154 B.n753 B.n52 10.6151
R1155 B.n753 B.n752 10.6151
R1156 B.n752 B.n751 10.6151
R1157 B.n751 B.n54 10.6151
R1158 B.n747 B.n54 10.6151
R1159 B.n747 B.n746 10.6151
R1160 B.n744 B.n58 10.6151
R1161 B.n740 B.n58 10.6151
R1162 B.n740 B.n739 10.6151
R1163 B.n739 B.n738 10.6151
R1164 B.n738 B.n60 10.6151
R1165 B.n734 B.n60 10.6151
R1166 B.n734 B.n733 10.6151
R1167 B.n733 B.n732 10.6151
R1168 B.n729 B.n728 10.6151
R1169 B.n728 B.n727 10.6151
R1170 B.n727 B.n66 10.6151
R1171 B.n723 B.n66 10.6151
R1172 B.n723 B.n722 10.6151
R1173 B.n722 B.n721 10.6151
R1174 B.n721 B.n68 10.6151
R1175 B.n717 B.n68 10.6151
R1176 B.n717 B.n716 10.6151
R1177 B.n716 B.n715 10.6151
R1178 B.n715 B.n70 10.6151
R1179 B.n711 B.n70 10.6151
R1180 B.n711 B.n710 10.6151
R1181 B.n710 B.n709 10.6151
R1182 B.n709 B.n72 10.6151
R1183 B.n705 B.n72 10.6151
R1184 B.n705 B.n704 10.6151
R1185 B.n704 B.n703 10.6151
R1186 B.n703 B.n74 10.6151
R1187 B.n699 B.n74 10.6151
R1188 B.n699 B.n698 10.6151
R1189 B.n698 B.n697 10.6151
R1190 B.n697 B.n76 10.6151
R1191 B.n693 B.n76 10.6151
R1192 B.n693 B.n692 10.6151
R1193 B.n692 B.n691 10.6151
R1194 B.n691 B.n78 10.6151
R1195 B.n687 B.n78 10.6151
R1196 B.n687 B.n686 10.6151
R1197 B.n686 B.n685 10.6151
R1198 B.n685 B.n80 10.6151
R1199 B.n681 B.n80 10.6151
R1200 B.n681 B.n680 10.6151
R1201 B.n680 B.n679 10.6151
R1202 B.n679 B.n82 10.6151
R1203 B.n675 B.n82 10.6151
R1204 B.n675 B.n674 10.6151
R1205 B.n674 B.n673 10.6151
R1206 B.n673 B.n84 10.6151
R1207 B.n669 B.n84 10.6151
R1208 B.n669 B.n668 10.6151
R1209 B.n668 B.n667 10.6151
R1210 B.n667 B.n86 10.6151
R1211 B.n663 B.n86 10.6151
R1212 B.n663 B.n662 10.6151
R1213 B.n662 B.n661 10.6151
R1214 B.n661 B.n88 10.6151
R1215 B.n657 B.n88 10.6151
R1216 B.n657 B.n656 10.6151
R1217 B.n656 B.n655 10.6151
R1218 B.n655 B.n90 10.6151
R1219 B.n651 B.n90 10.6151
R1220 B.n651 B.n650 10.6151
R1221 B.n650 B.n649 10.6151
R1222 B.n649 B.n92 10.6151
R1223 B.n645 B.n92 10.6151
R1224 B.n645 B.n644 10.6151
R1225 B.n644 B.n643 10.6151
R1226 B.n499 B.n142 10.6151
R1227 B.n500 B.n499 10.6151
R1228 B.n501 B.n500 10.6151
R1229 B.n501 B.n140 10.6151
R1230 B.n505 B.n140 10.6151
R1231 B.n506 B.n505 10.6151
R1232 B.n507 B.n506 10.6151
R1233 B.n507 B.n138 10.6151
R1234 B.n511 B.n138 10.6151
R1235 B.n512 B.n511 10.6151
R1236 B.n513 B.n512 10.6151
R1237 B.n513 B.n136 10.6151
R1238 B.n517 B.n136 10.6151
R1239 B.n518 B.n517 10.6151
R1240 B.n519 B.n518 10.6151
R1241 B.n519 B.n134 10.6151
R1242 B.n523 B.n134 10.6151
R1243 B.n524 B.n523 10.6151
R1244 B.n525 B.n524 10.6151
R1245 B.n525 B.n132 10.6151
R1246 B.n529 B.n132 10.6151
R1247 B.n530 B.n529 10.6151
R1248 B.n531 B.n530 10.6151
R1249 B.n531 B.n130 10.6151
R1250 B.n535 B.n130 10.6151
R1251 B.n536 B.n535 10.6151
R1252 B.n537 B.n536 10.6151
R1253 B.n537 B.n128 10.6151
R1254 B.n541 B.n128 10.6151
R1255 B.n542 B.n541 10.6151
R1256 B.n543 B.n542 10.6151
R1257 B.n543 B.n126 10.6151
R1258 B.n547 B.n126 10.6151
R1259 B.n548 B.n547 10.6151
R1260 B.n549 B.n548 10.6151
R1261 B.n549 B.n124 10.6151
R1262 B.n553 B.n124 10.6151
R1263 B.n554 B.n553 10.6151
R1264 B.n555 B.n554 10.6151
R1265 B.n555 B.n122 10.6151
R1266 B.n559 B.n122 10.6151
R1267 B.n560 B.n559 10.6151
R1268 B.n561 B.n560 10.6151
R1269 B.n561 B.n120 10.6151
R1270 B.n565 B.n120 10.6151
R1271 B.n566 B.n565 10.6151
R1272 B.n567 B.n566 10.6151
R1273 B.n567 B.n118 10.6151
R1274 B.n571 B.n118 10.6151
R1275 B.n572 B.n571 10.6151
R1276 B.n573 B.n572 10.6151
R1277 B.n573 B.n116 10.6151
R1278 B.n577 B.n116 10.6151
R1279 B.n578 B.n577 10.6151
R1280 B.n579 B.n578 10.6151
R1281 B.n579 B.n114 10.6151
R1282 B.n583 B.n114 10.6151
R1283 B.n584 B.n583 10.6151
R1284 B.n585 B.n584 10.6151
R1285 B.n585 B.n112 10.6151
R1286 B.n589 B.n112 10.6151
R1287 B.n590 B.n589 10.6151
R1288 B.n591 B.n590 10.6151
R1289 B.n591 B.n110 10.6151
R1290 B.n595 B.n110 10.6151
R1291 B.n596 B.n595 10.6151
R1292 B.n597 B.n596 10.6151
R1293 B.n597 B.n108 10.6151
R1294 B.n601 B.n108 10.6151
R1295 B.n602 B.n601 10.6151
R1296 B.n603 B.n602 10.6151
R1297 B.n603 B.n106 10.6151
R1298 B.n607 B.n106 10.6151
R1299 B.n608 B.n607 10.6151
R1300 B.n609 B.n608 10.6151
R1301 B.n609 B.n104 10.6151
R1302 B.n613 B.n104 10.6151
R1303 B.n614 B.n613 10.6151
R1304 B.n615 B.n614 10.6151
R1305 B.n615 B.n102 10.6151
R1306 B.n619 B.n102 10.6151
R1307 B.n620 B.n619 10.6151
R1308 B.n621 B.n620 10.6151
R1309 B.n621 B.n100 10.6151
R1310 B.n625 B.n100 10.6151
R1311 B.n626 B.n625 10.6151
R1312 B.n627 B.n626 10.6151
R1313 B.n627 B.n98 10.6151
R1314 B.n631 B.n98 10.6151
R1315 B.n632 B.n631 10.6151
R1316 B.n633 B.n632 10.6151
R1317 B.n633 B.n96 10.6151
R1318 B.n637 B.n96 10.6151
R1319 B.n638 B.n637 10.6151
R1320 B.n639 B.n638 10.6151
R1321 B.n639 B.n94 10.6151
R1322 B.n307 B.n210 10.6151
R1323 B.n308 B.n307 10.6151
R1324 B.n309 B.n308 10.6151
R1325 B.n309 B.n208 10.6151
R1326 B.n313 B.n208 10.6151
R1327 B.n314 B.n313 10.6151
R1328 B.n315 B.n314 10.6151
R1329 B.n315 B.n206 10.6151
R1330 B.n319 B.n206 10.6151
R1331 B.n320 B.n319 10.6151
R1332 B.n321 B.n320 10.6151
R1333 B.n321 B.n204 10.6151
R1334 B.n325 B.n204 10.6151
R1335 B.n326 B.n325 10.6151
R1336 B.n327 B.n326 10.6151
R1337 B.n327 B.n202 10.6151
R1338 B.n331 B.n202 10.6151
R1339 B.n332 B.n331 10.6151
R1340 B.n333 B.n332 10.6151
R1341 B.n333 B.n200 10.6151
R1342 B.n337 B.n200 10.6151
R1343 B.n338 B.n337 10.6151
R1344 B.n339 B.n338 10.6151
R1345 B.n339 B.n198 10.6151
R1346 B.n343 B.n198 10.6151
R1347 B.n344 B.n343 10.6151
R1348 B.n345 B.n344 10.6151
R1349 B.n345 B.n196 10.6151
R1350 B.n349 B.n196 10.6151
R1351 B.n350 B.n349 10.6151
R1352 B.n351 B.n350 10.6151
R1353 B.n351 B.n194 10.6151
R1354 B.n355 B.n194 10.6151
R1355 B.n356 B.n355 10.6151
R1356 B.n357 B.n356 10.6151
R1357 B.n357 B.n192 10.6151
R1358 B.n361 B.n192 10.6151
R1359 B.n362 B.n361 10.6151
R1360 B.n363 B.n362 10.6151
R1361 B.n363 B.n190 10.6151
R1362 B.n367 B.n190 10.6151
R1363 B.n368 B.n367 10.6151
R1364 B.n369 B.n368 10.6151
R1365 B.n369 B.n188 10.6151
R1366 B.n373 B.n188 10.6151
R1367 B.n374 B.n373 10.6151
R1368 B.n375 B.n374 10.6151
R1369 B.n375 B.n186 10.6151
R1370 B.n379 B.n186 10.6151
R1371 B.n380 B.n379 10.6151
R1372 B.n381 B.n380 10.6151
R1373 B.n381 B.n184 10.6151
R1374 B.n385 B.n184 10.6151
R1375 B.n386 B.n385 10.6151
R1376 B.n387 B.n386 10.6151
R1377 B.n387 B.n182 10.6151
R1378 B.n391 B.n182 10.6151
R1379 B.n392 B.n391 10.6151
R1380 B.n394 B.n178 10.6151
R1381 B.n398 B.n178 10.6151
R1382 B.n399 B.n398 10.6151
R1383 B.n400 B.n399 10.6151
R1384 B.n400 B.n176 10.6151
R1385 B.n404 B.n176 10.6151
R1386 B.n405 B.n404 10.6151
R1387 B.n406 B.n405 10.6151
R1388 B.n410 B.n409 10.6151
R1389 B.n411 B.n410 10.6151
R1390 B.n411 B.n170 10.6151
R1391 B.n415 B.n170 10.6151
R1392 B.n416 B.n415 10.6151
R1393 B.n417 B.n416 10.6151
R1394 B.n417 B.n168 10.6151
R1395 B.n421 B.n168 10.6151
R1396 B.n422 B.n421 10.6151
R1397 B.n423 B.n422 10.6151
R1398 B.n423 B.n166 10.6151
R1399 B.n427 B.n166 10.6151
R1400 B.n428 B.n427 10.6151
R1401 B.n429 B.n428 10.6151
R1402 B.n429 B.n164 10.6151
R1403 B.n433 B.n164 10.6151
R1404 B.n434 B.n433 10.6151
R1405 B.n435 B.n434 10.6151
R1406 B.n435 B.n162 10.6151
R1407 B.n439 B.n162 10.6151
R1408 B.n440 B.n439 10.6151
R1409 B.n441 B.n440 10.6151
R1410 B.n441 B.n160 10.6151
R1411 B.n445 B.n160 10.6151
R1412 B.n446 B.n445 10.6151
R1413 B.n447 B.n446 10.6151
R1414 B.n447 B.n158 10.6151
R1415 B.n451 B.n158 10.6151
R1416 B.n452 B.n451 10.6151
R1417 B.n453 B.n452 10.6151
R1418 B.n453 B.n156 10.6151
R1419 B.n457 B.n156 10.6151
R1420 B.n458 B.n457 10.6151
R1421 B.n459 B.n458 10.6151
R1422 B.n459 B.n154 10.6151
R1423 B.n463 B.n154 10.6151
R1424 B.n464 B.n463 10.6151
R1425 B.n465 B.n464 10.6151
R1426 B.n465 B.n152 10.6151
R1427 B.n469 B.n152 10.6151
R1428 B.n470 B.n469 10.6151
R1429 B.n471 B.n470 10.6151
R1430 B.n471 B.n150 10.6151
R1431 B.n475 B.n150 10.6151
R1432 B.n476 B.n475 10.6151
R1433 B.n477 B.n476 10.6151
R1434 B.n477 B.n148 10.6151
R1435 B.n481 B.n148 10.6151
R1436 B.n482 B.n481 10.6151
R1437 B.n483 B.n482 10.6151
R1438 B.n483 B.n146 10.6151
R1439 B.n487 B.n146 10.6151
R1440 B.n488 B.n487 10.6151
R1441 B.n489 B.n488 10.6151
R1442 B.n489 B.n144 10.6151
R1443 B.n493 B.n144 10.6151
R1444 B.n494 B.n493 10.6151
R1445 B.n495 B.n494 10.6151
R1446 B.n303 B.n302 10.6151
R1447 B.n302 B.n301 10.6151
R1448 B.n301 B.n212 10.6151
R1449 B.n297 B.n212 10.6151
R1450 B.n297 B.n296 10.6151
R1451 B.n296 B.n295 10.6151
R1452 B.n295 B.n214 10.6151
R1453 B.n291 B.n214 10.6151
R1454 B.n291 B.n290 10.6151
R1455 B.n290 B.n289 10.6151
R1456 B.n289 B.n216 10.6151
R1457 B.n285 B.n216 10.6151
R1458 B.n285 B.n284 10.6151
R1459 B.n284 B.n283 10.6151
R1460 B.n283 B.n218 10.6151
R1461 B.n279 B.n218 10.6151
R1462 B.n279 B.n278 10.6151
R1463 B.n278 B.n277 10.6151
R1464 B.n277 B.n220 10.6151
R1465 B.n273 B.n220 10.6151
R1466 B.n273 B.n272 10.6151
R1467 B.n272 B.n271 10.6151
R1468 B.n271 B.n222 10.6151
R1469 B.n267 B.n222 10.6151
R1470 B.n267 B.n266 10.6151
R1471 B.n266 B.n265 10.6151
R1472 B.n265 B.n224 10.6151
R1473 B.n261 B.n224 10.6151
R1474 B.n261 B.n260 10.6151
R1475 B.n260 B.n259 10.6151
R1476 B.n259 B.n226 10.6151
R1477 B.n255 B.n226 10.6151
R1478 B.n255 B.n254 10.6151
R1479 B.n254 B.n253 10.6151
R1480 B.n253 B.n228 10.6151
R1481 B.n249 B.n228 10.6151
R1482 B.n249 B.n248 10.6151
R1483 B.n248 B.n247 10.6151
R1484 B.n247 B.n230 10.6151
R1485 B.n243 B.n230 10.6151
R1486 B.n243 B.n242 10.6151
R1487 B.n242 B.n241 10.6151
R1488 B.n241 B.n232 10.6151
R1489 B.n237 B.n232 10.6151
R1490 B.n237 B.n236 10.6151
R1491 B.n236 B.n235 10.6151
R1492 B.n235 B.n0 10.6151
R1493 B.n903 B.n1 10.6151
R1494 B.n903 B.n902 10.6151
R1495 B.n902 B.n901 10.6151
R1496 B.n901 B.n4 10.6151
R1497 B.n897 B.n4 10.6151
R1498 B.n897 B.n896 10.6151
R1499 B.n896 B.n895 10.6151
R1500 B.n895 B.n6 10.6151
R1501 B.n891 B.n6 10.6151
R1502 B.n891 B.n890 10.6151
R1503 B.n890 B.n889 10.6151
R1504 B.n889 B.n8 10.6151
R1505 B.n885 B.n8 10.6151
R1506 B.n885 B.n884 10.6151
R1507 B.n884 B.n883 10.6151
R1508 B.n883 B.n10 10.6151
R1509 B.n879 B.n10 10.6151
R1510 B.n879 B.n878 10.6151
R1511 B.n878 B.n877 10.6151
R1512 B.n877 B.n12 10.6151
R1513 B.n873 B.n12 10.6151
R1514 B.n873 B.n872 10.6151
R1515 B.n872 B.n871 10.6151
R1516 B.n871 B.n14 10.6151
R1517 B.n867 B.n14 10.6151
R1518 B.n867 B.n866 10.6151
R1519 B.n866 B.n865 10.6151
R1520 B.n865 B.n16 10.6151
R1521 B.n861 B.n16 10.6151
R1522 B.n861 B.n860 10.6151
R1523 B.n860 B.n859 10.6151
R1524 B.n859 B.n18 10.6151
R1525 B.n855 B.n18 10.6151
R1526 B.n855 B.n854 10.6151
R1527 B.n854 B.n853 10.6151
R1528 B.n853 B.n20 10.6151
R1529 B.n849 B.n20 10.6151
R1530 B.n849 B.n848 10.6151
R1531 B.n848 B.n847 10.6151
R1532 B.n847 B.n22 10.6151
R1533 B.n843 B.n22 10.6151
R1534 B.n843 B.n842 10.6151
R1535 B.n842 B.n841 10.6151
R1536 B.n841 B.n24 10.6151
R1537 B.n837 B.n24 10.6151
R1538 B.n837 B.n836 10.6151
R1539 B.n836 B.n835 10.6151
R1540 B.n745 B.n744 6.5566
R1541 B.n732 B.n64 6.5566
R1542 B.n394 B.n393 6.5566
R1543 B.n406 B.n174 6.5566
R1544 B.n746 B.n745 4.05904
R1545 B.n729 B.n64 4.05904
R1546 B.n393 B.n392 4.05904
R1547 B.n409 B.n174 4.05904
R1548 B.n907 B.n0 2.81026
R1549 B.n907 B.n1 2.81026
R1550 VN.n8 VN.t8 254.249
R1551 VN.n41 VN.t1 254.249
R1552 VN.n16 VN.t3 221.373
R1553 VN.n7 VN.t7 221.373
R1554 VN.n23 VN.t2 221.373
R1555 VN.n31 VN.t6 221.373
R1556 VN.n49 VN.t0 221.373
R1557 VN.n40 VN.t4 221.373
R1558 VN.n56 VN.t5 221.373
R1559 VN.n64 VN.t9 221.373
R1560 VN.n32 VN.n31 183.924
R1561 VN.n65 VN.n64 183.924
R1562 VN.n63 VN.n33 161.3
R1563 VN.n62 VN.n61 161.3
R1564 VN.n60 VN.n34 161.3
R1565 VN.n59 VN.n58 161.3
R1566 VN.n57 VN.n35 161.3
R1567 VN.n55 VN.n54 161.3
R1568 VN.n53 VN.n36 161.3
R1569 VN.n52 VN.n51 161.3
R1570 VN.n50 VN.n37 161.3
R1571 VN.n49 VN.n48 161.3
R1572 VN.n47 VN.n38 161.3
R1573 VN.n46 VN.n45 161.3
R1574 VN.n44 VN.n39 161.3
R1575 VN.n43 VN.n42 161.3
R1576 VN.n30 VN.n0 161.3
R1577 VN.n29 VN.n28 161.3
R1578 VN.n27 VN.n1 161.3
R1579 VN.n26 VN.n25 161.3
R1580 VN.n24 VN.n2 161.3
R1581 VN.n22 VN.n21 161.3
R1582 VN.n20 VN.n3 161.3
R1583 VN.n19 VN.n18 161.3
R1584 VN.n17 VN.n4 161.3
R1585 VN.n16 VN.n15 161.3
R1586 VN.n14 VN.n5 161.3
R1587 VN.n13 VN.n12 161.3
R1588 VN.n11 VN.n6 161.3
R1589 VN.n10 VN.n9 161.3
R1590 VN.n8 VN.n7 56.9995
R1591 VN.n41 VN.n40 56.9995
R1592 VN VN.n65 54.2259
R1593 VN.n12 VN.n11 53.6554
R1594 VN.n18 VN.n3 53.6554
R1595 VN.n45 VN.n44 53.6554
R1596 VN.n51 VN.n36 53.6554
R1597 VN.n25 VN.n1 49.7803
R1598 VN.n58 VN.n34 49.7803
R1599 VN.n29 VN.n1 31.3737
R1600 VN.n62 VN.n34 31.3737
R1601 VN.n12 VN.n5 27.4986
R1602 VN.n18 VN.n17 27.4986
R1603 VN.n45 VN.n38 27.4986
R1604 VN.n51 VN.n50 27.4986
R1605 VN.n11 VN.n10 24.5923
R1606 VN.n16 VN.n5 24.5923
R1607 VN.n17 VN.n16 24.5923
R1608 VN.n22 VN.n3 24.5923
R1609 VN.n25 VN.n24 24.5923
R1610 VN.n30 VN.n29 24.5923
R1611 VN.n44 VN.n43 24.5923
R1612 VN.n50 VN.n49 24.5923
R1613 VN.n49 VN.n38 24.5923
R1614 VN.n58 VN.n57 24.5923
R1615 VN.n55 VN.n36 24.5923
R1616 VN.n63 VN.n62 24.5923
R1617 VN.n10 VN.n7 13.2801
R1618 VN.n23 VN.n22 13.2801
R1619 VN.n43 VN.n40 13.2801
R1620 VN.n56 VN.n55 13.2801
R1621 VN.n42 VN.n41 12.447
R1622 VN.n9 VN.n8 12.447
R1623 VN.n24 VN.n23 11.3127
R1624 VN.n57 VN.n56 11.3127
R1625 VN.n31 VN.n30 1.96785
R1626 VN.n64 VN.n63 1.96785
R1627 VN.n65 VN.n33 0.189894
R1628 VN.n61 VN.n33 0.189894
R1629 VN.n61 VN.n60 0.189894
R1630 VN.n60 VN.n59 0.189894
R1631 VN.n59 VN.n35 0.189894
R1632 VN.n54 VN.n35 0.189894
R1633 VN.n54 VN.n53 0.189894
R1634 VN.n53 VN.n52 0.189894
R1635 VN.n52 VN.n37 0.189894
R1636 VN.n48 VN.n37 0.189894
R1637 VN.n48 VN.n47 0.189894
R1638 VN.n47 VN.n46 0.189894
R1639 VN.n46 VN.n39 0.189894
R1640 VN.n42 VN.n39 0.189894
R1641 VN.n9 VN.n6 0.189894
R1642 VN.n13 VN.n6 0.189894
R1643 VN.n14 VN.n13 0.189894
R1644 VN.n15 VN.n14 0.189894
R1645 VN.n15 VN.n4 0.189894
R1646 VN.n19 VN.n4 0.189894
R1647 VN.n20 VN.n19 0.189894
R1648 VN.n21 VN.n20 0.189894
R1649 VN.n21 VN.n2 0.189894
R1650 VN.n26 VN.n2 0.189894
R1651 VN.n27 VN.n26 0.189894
R1652 VN.n28 VN.n27 0.189894
R1653 VN.n28 VN.n0 0.189894
R1654 VN.n32 VN.n0 0.189894
R1655 VN VN.n32 0.0516364
R1656 VDD2.n1 VDD2.t1 71.4678
R1657 VDD2.n4 VDD2.t0 69.5111
R1658 VDD2.n3 VDD2.n2 69.0991
R1659 VDD2 VDD2.n7 69.0963
R1660 VDD2.n6 VDD2.n5 67.6871
R1661 VDD2.n1 VDD2.n0 67.6868
R1662 VDD2.n4 VDD2.n3 48.3726
R1663 VDD2.n6 VDD2.n4 1.9574
R1664 VDD2.n7 VDD2.t5 1.82457
R1665 VDD2.n7 VDD2.t8 1.82457
R1666 VDD2.n5 VDD2.t4 1.82457
R1667 VDD2.n5 VDD2.t9 1.82457
R1668 VDD2.n2 VDD2.t7 1.82457
R1669 VDD2.n2 VDD2.t3 1.82457
R1670 VDD2.n0 VDD2.t2 1.82457
R1671 VDD2.n0 VDD2.t6 1.82457
R1672 VDD2 VDD2.n6 0.547914
R1673 VDD2.n3 VDD2.n1 0.434378
C0 VP VDD2 0.500282f
C1 VN VDD2 14.5766f
C2 VP VN 8.495741f
C3 w_n3694_n4532# B 11.0688f
C4 w_n3694_n4532# VTAIL 3.9592f
C5 B VTAIL 4.67253f
C6 w_n3694_n4532# VDD1 2.94696f
C7 B VDD1 2.67096f
C8 w_n3694_n4532# VDD2 3.05631f
C9 B VDD2 2.76318f
C10 VP w_n3694_n4532# 8.27308f
C11 w_n3694_n4532# VN 7.79417f
C12 VDD1 VTAIL 13.5999f
C13 VP B 1.98863f
C14 VN B 1.18696f
C15 VTAIL VDD2 13.6438f
C16 VP VTAIL 14.7154f
C17 VN VTAIL 14.701f
C18 VDD1 VDD2 1.74561f
C19 VP VDD1 14.919499f
C20 VN VDD1 0.152137f
C21 VDD2 VSUBS 2.049889f
C22 VDD1 VSUBS 1.845563f
C23 VTAIL VSUBS 1.348117f
C24 VN VSUBS 6.8787f
C25 VP VSUBS 3.59667f
C26 B VSUBS 5.038505f
C27 w_n3694_n4532# VSUBS 0.204751p
C28 VDD2.t1 VSUBS 4.05438f
C29 VDD2.t2 VSUBS 0.375292f
C30 VDD2.t6 VSUBS 0.375292f
C31 VDD2.n0 VSUBS 3.10726f
C32 VDD2.n1 VSUBS 1.52494f
C33 VDD2.t7 VSUBS 0.375292f
C34 VDD2.t3 VSUBS 0.375292f
C35 VDD2.n2 VSUBS 3.12427f
C36 VDD2.n3 VSUBS 3.42216f
C37 VDD2.t0 VSUBS 4.03224f
C38 VDD2.n4 VSUBS 3.87197f
C39 VDD2.t4 VSUBS 0.375292f
C40 VDD2.t9 VSUBS 0.375292f
C41 VDD2.n5 VSUBS 3.10726f
C42 VDD2.n6 VSUBS 0.746563f
C43 VDD2.t5 VSUBS 0.375292f
C44 VDD2.t8 VSUBS 0.375292f
C45 VDD2.n7 VSUBS 3.12421f
C46 VN.n0 VSUBS 0.03014f
C47 VN.t6 VSUBS 2.86542f
C48 VN.n1 VSUBS 0.027998f
C49 VN.n2 VSUBS 0.03014f
C50 VN.t2 VSUBS 2.86542f
C51 VN.n3 VSUBS 0.052902f
C52 VN.n4 VSUBS 0.03014f
C53 VN.t3 VSUBS 2.86542f
C54 VN.n5 VSUBS 0.058458f
C55 VN.n6 VSUBS 0.03014f
C56 VN.t7 VSUBS 2.86542f
C57 VN.n7 VSUBS 1.0721f
C58 VN.t8 VSUBS 3.01418f
C59 VN.n8 VSUBS 1.07442f
C60 VN.n9 VSUBS 0.224629f
C61 VN.n10 VSUBS 0.043199f
C62 VN.n11 VSUBS 0.052902f
C63 VN.n12 VSUBS 0.032157f
C64 VN.n13 VSUBS 0.03014f
C65 VN.n14 VSUBS 0.03014f
C66 VN.n15 VSUBS 0.03014f
C67 VN.n16 VSUBS 1.02924f
C68 VN.n17 VSUBS 0.058458f
C69 VN.n18 VSUBS 0.032157f
C70 VN.n19 VSUBS 0.03014f
C71 VN.n20 VSUBS 0.03014f
C72 VN.n21 VSUBS 0.03014f
C73 VN.n22 VSUBS 0.043199f
C74 VN.n23 VSUBS 1.00094f
C75 VN.n24 VSUBS 0.040992f
C76 VN.n25 VSUBS 0.055333f
C77 VN.n26 VSUBS 0.03014f
C78 VN.n27 VSUBS 0.03014f
C79 VN.n28 VSUBS 0.03014f
C80 VN.n29 VSUBS 0.060185f
C81 VN.n30 VSUBS 0.030507f
C82 VN.n31 VSUBS 1.07318f
C83 VN.n32 VSUBS 0.033491f
C84 VN.n33 VSUBS 0.03014f
C85 VN.t9 VSUBS 2.86542f
C86 VN.n34 VSUBS 0.027998f
C87 VN.n35 VSUBS 0.03014f
C88 VN.t5 VSUBS 2.86542f
C89 VN.n36 VSUBS 0.052902f
C90 VN.n37 VSUBS 0.03014f
C91 VN.t0 VSUBS 2.86542f
C92 VN.n38 VSUBS 0.058458f
C93 VN.n39 VSUBS 0.03014f
C94 VN.t4 VSUBS 2.86542f
C95 VN.n40 VSUBS 1.0721f
C96 VN.t1 VSUBS 3.01418f
C97 VN.n41 VSUBS 1.07442f
C98 VN.n42 VSUBS 0.224629f
C99 VN.n43 VSUBS 0.043199f
C100 VN.n44 VSUBS 0.052902f
C101 VN.n45 VSUBS 0.032157f
C102 VN.n46 VSUBS 0.03014f
C103 VN.n47 VSUBS 0.03014f
C104 VN.n48 VSUBS 0.03014f
C105 VN.n49 VSUBS 1.02924f
C106 VN.n50 VSUBS 0.058458f
C107 VN.n51 VSUBS 0.032157f
C108 VN.n52 VSUBS 0.03014f
C109 VN.n53 VSUBS 0.03014f
C110 VN.n54 VSUBS 0.03014f
C111 VN.n55 VSUBS 0.043199f
C112 VN.n56 VSUBS 1.00094f
C113 VN.n57 VSUBS 0.040992f
C114 VN.n58 VSUBS 0.055333f
C115 VN.n59 VSUBS 0.03014f
C116 VN.n60 VSUBS 0.03014f
C117 VN.n61 VSUBS 0.03014f
C118 VN.n62 VSUBS 0.060185f
C119 VN.n63 VSUBS 0.030507f
C120 VN.n64 VSUBS 1.07318f
C121 VN.n65 VSUBS 1.85763f
C122 B.n0 VSUBS 0.004999f
C123 B.n1 VSUBS 0.004999f
C124 B.n2 VSUBS 0.007905f
C125 B.n3 VSUBS 0.007905f
C126 B.n4 VSUBS 0.007905f
C127 B.n5 VSUBS 0.007905f
C128 B.n6 VSUBS 0.007905f
C129 B.n7 VSUBS 0.007905f
C130 B.n8 VSUBS 0.007905f
C131 B.n9 VSUBS 0.007905f
C132 B.n10 VSUBS 0.007905f
C133 B.n11 VSUBS 0.007905f
C134 B.n12 VSUBS 0.007905f
C135 B.n13 VSUBS 0.007905f
C136 B.n14 VSUBS 0.007905f
C137 B.n15 VSUBS 0.007905f
C138 B.n16 VSUBS 0.007905f
C139 B.n17 VSUBS 0.007905f
C140 B.n18 VSUBS 0.007905f
C141 B.n19 VSUBS 0.007905f
C142 B.n20 VSUBS 0.007905f
C143 B.n21 VSUBS 0.007905f
C144 B.n22 VSUBS 0.007905f
C145 B.n23 VSUBS 0.007905f
C146 B.n24 VSUBS 0.007905f
C147 B.n25 VSUBS 0.007905f
C148 B.n26 VSUBS 0.019711f
C149 B.n27 VSUBS 0.007905f
C150 B.n28 VSUBS 0.007905f
C151 B.n29 VSUBS 0.007905f
C152 B.n30 VSUBS 0.007905f
C153 B.n31 VSUBS 0.007905f
C154 B.n32 VSUBS 0.007905f
C155 B.n33 VSUBS 0.007905f
C156 B.n34 VSUBS 0.007905f
C157 B.n35 VSUBS 0.007905f
C158 B.n36 VSUBS 0.007905f
C159 B.n37 VSUBS 0.007905f
C160 B.n38 VSUBS 0.007905f
C161 B.n39 VSUBS 0.007905f
C162 B.n40 VSUBS 0.007905f
C163 B.n41 VSUBS 0.007905f
C164 B.n42 VSUBS 0.007905f
C165 B.n43 VSUBS 0.007905f
C166 B.n44 VSUBS 0.007905f
C167 B.n45 VSUBS 0.007905f
C168 B.n46 VSUBS 0.007905f
C169 B.n47 VSUBS 0.007905f
C170 B.n48 VSUBS 0.007905f
C171 B.n49 VSUBS 0.007905f
C172 B.n50 VSUBS 0.007905f
C173 B.n51 VSUBS 0.007905f
C174 B.n52 VSUBS 0.007905f
C175 B.n53 VSUBS 0.007905f
C176 B.n54 VSUBS 0.007905f
C177 B.n55 VSUBS 0.007905f
C178 B.t2 VSUBS 0.678928f
C179 B.t1 VSUBS 0.698234f
C180 B.t0 VSUBS 1.69483f
C181 B.n56 VSUBS 0.340857f
C182 B.n57 VSUBS 0.078344f
C183 B.n58 VSUBS 0.007905f
C184 B.n59 VSUBS 0.007905f
C185 B.n60 VSUBS 0.007905f
C186 B.n61 VSUBS 0.007905f
C187 B.t8 VSUBS 0.678903f
C188 B.t7 VSUBS 0.698213f
C189 B.t6 VSUBS 1.69483f
C190 B.n62 VSUBS 0.340877f
C191 B.n63 VSUBS 0.078369f
C192 B.n64 VSUBS 0.018316f
C193 B.n65 VSUBS 0.007905f
C194 B.n66 VSUBS 0.007905f
C195 B.n67 VSUBS 0.007905f
C196 B.n68 VSUBS 0.007905f
C197 B.n69 VSUBS 0.007905f
C198 B.n70 VSUBS 0.007905f
C199 B.n71 VSUBS 0.007905f
C200 B.n72 VSUBS 0.007905f
C201 B.n73 VSUBS 0.007905f
C202 B.n74 VSUBS 0.007905f
C203 B.n75 VSUBS 0.007905f
C204 B.n76 VSUBS 0.007905f
C205 B.n77 VSUBS 0.007905f
C206 B.n78 VSUBS 0.007905f
C207 B.n79 VSUBS 0.007905f
C208 B.n80 VSUBS 0.007905f
C209 B.n81 VSUBS 0.007905f
C210 B.n82 VSUBS 0.007905f
C211 B.n83 VSUBS 0.007905f
C212 B.n84 VSUBS 0.007905f
C213 B.n85 VSUBS 0.007905f
C214 B.n86 VSUBS 0.007905f
C215 B.n87 VSUBS 0.007905f
C216 B.n88 VSUBS 0.007905f
C217 B.n89 VSUBS 0.007905f
C218 B.n90 VSUBS 0.007905f
C219 B.n91 VSUBS 0.007905f
C220 B.n92 VSUBS 0.007905f
C221 B.n93 VSUBS 0.007905f
C222 B.n94 VSUBS 0.019538f
C223 B.n95 VSUBS 0.007905f
C224 B.n96 VSUBS 0.007905f
C225 B.n97 VSUBS 0.007905f
C226 B.n98 VSUBS 0.007905f
C227 B.n99 VSUBS 0.007905f
C228 B.n100 VSUBS 0.007905f
C229 B.n101 VSUBS 0.007905f
C230 B.n102 VSUBS 0.007905f
C231 B.n103 VSUBS 0.007905f
C232 B.n104 VSUBS 0.007905f
C233 B.n105 VSUBS 0.007905f
C234 B.n106 VSUBS 0.007905f
C235 B.n107 VSUBS 0.007905f
C236 B.n108 VSUBS 0.007905f
C237 B.n109 VSUBS 0.007905f
C238 B.n110 VSUBS 0.007905f
C239 B.n111 VSUBS 0.007905f
C240 B.n112 VSUBS 0.007905f
C241 B.n113 VSUBS 0.007905f
C242 B.n114 VSUBS 0.007905f
C243 B.n115 VSUBS 0.007905f
C244 B.n116 VSUBS 0.007905f
C245 B.n117 VSUBS 0.007905f
C246 B.n118 VSUBS 0.007905f
C247 B.n119 VSUBS 0.007905f
C248 B.n120 VSUBS 0.007905f
C249 B.n121 VSUBS 0.007905f
C250 B.n122 VSUBS 0.007905f
C251 B.n123 VSUBS 0.007905f
C252 B.n124 VSUBS 0.007905f
C253 B.n125 VSUBS 0.007905f
C254 B.n126 VSUBS 0.007905f
C255 B.n127 VSUBS 0.007905f
C256 B.n128 VSUBS 0.007905f
C257 B.n129 VSUBS 0.007905f
C258 B.n130 VSUBS 0.007905f
C259 B.n131 VSUBS 0.007905f
C260 B.n132 VSUBS 0.007905f
C261 B.n133 VSUBS 0.007905f
C262 B.n134 VSUBS 0.007905f
C263 B.n135 VSUBS 0.007905f
C264 B.n136 VSUBS 0.007905f
C265 B.n137 VSUBS 0.007905f
C266 B.n138 VSUBS 0.007905f
C267 B.n139 VSUBS 0.007905f
C268 B.n140 VSUBS 0.007905f
C269 B.n141 VSUBS 0.007905f
C270 B.n142 VSUBS 0.018654f
C271 B.n143 VSUBS 0.007905f
C272 B.n144 VSUBS 0.007905f
C273 B.n145 VSUBS 0.007905f
C274 B.n146 VSUBS 0.007905f
C275 B.n147 VSUBS 0.007905f
C276 B.n148 VSUBS 0.007905f
C277 B.n149 VSUBS 0.007905f
C278 B.n150 VSUBS 0.007905f
C279 B.n151 VSUBS 0.007905f
C280 B.n152 VSUBS 0.007905f
C281 B.n153 VSUBS 0.007905f
C282 B.n154 VSUBS 0.007905f
C283 B.n155 VSUBS 0.007905f
C284 B.n156 VSUBS 0.007905f
C285 B.n157 VSUBS 0.007905f
C286 B.n158 VSUBS 0.007905f
C287 B.n159 VSUBS 0.007905f
C288 B.n160 VSUBS 0.007905f
C289 B.n161 VSUBS 0.007905f
C290 B.n162 VSUBS 0.007905f
C291 B.n163 VSUBS 0.007905f
C292 B.n164 VSUBS 0.007905f
C293 B.n165 VSUBS 0.007905f
C294 B.n166 VSUBS 0.007905f
C295 B.n167 VSUBS 0.007905f
C296 B.n168 VSUBS 0.007905f
C297 B.n169 VSUBS 0.007905f
C298 B.n170 VSUBS 0.007905f
C299 B.n171 VSUBS 0.007905f
C300 B.t10 VSUBS 0.678903f
C301 B.t11 VSUBS 0.698213f
C302 B.t9 VSUBS 1.69483f
C303 B.n172 VSUBS 0.340877f
C304 B.n173 VSUBS 0.078369f
C305 B.n174 VSUBS 0.018316f
C306 B.n175 VSUBS 0.007905f
C307 B.n176 VSUBS 0.007905f
C308 B.n177 VSUBS 0.007905f
C309 B.n178 VSUBS 0.007905f
C310 B.n179 VSUBS 0.007905f
C311 B.t4 VSUBS 0.678928f
C312 B.t5 VSUBS 0.698234f
C313 B.t3 VSUBS 1.69483f
C314 B.n180 VSUBS 0.340857f
C315 B.n181 VSUBS 0.078344f
C316 B.n182 VSUBS 0.007905f
C317 B.n183 VSUBS 0.007905f
C318 B.n184 VSUBS 0.007905f
C319 B.n185 VSUBS 0.007905f
C320 B.n186 VSUBS 0.007905f
C321 B.n187 VSUBS 0.007905f
C322 B.n188 VSUBS 0.007905f
C323 B.n189 VSUBS 0.007905f
C324 B.n190 VSUBS 0.007905f
C325 B.n191 VSUBS 0.007905f
C326 B.n192 VSUBS 0.007905f
C327 B.n193 VSUBS 0.007905f
C328 B.n194 VSUBS 0.007905f
C329 B.n195 VSUBS 0.007905f
C330 B.n196 VSUBS 0.007905f
C331 B.n197 VSUBS 0.007905f
C332 B.n198 VSUBS 0.007905f
C333 B.n199 VSUBS 0.007905f
C334 B.n200 VSUBS 0.007905f
C335 B.n201 VSUBS 0.007905f
C336 B.n202 VSUBS 0.007905f
C337 B.n203 VSUBS 0.007905f
C338 B.n204 VSUBS 0.007905f
C339 B.n205 VSUBS 0.007905f
C340 B.n206 VSUBS 0.007905f
C341 B.n207 VSUBS 0.007905f
C342 B.n208 VSUBS 0.007905f
C343 B.n209 VSUBS 0.007905f
C344 B.n210 VSUBS 0.019711f
C345 B.n211 VSUBS 0.007905f
C346 B.n212 VSUBS 0.007905f
C347 B.n213 VSUBS 0.007905f
C348 B.n214 VSUBS 0.007905f
C349 B.n215 VSUBS 0.007905f
C350 B.n216 VSUBS 0.007905f
C351 B.n217 VSUBS 0.007905f
C352 B.n218 VSUBS 0.007905f
C353 B.n219 VSUBS 0.007905f
C354 B.n220 VSUBS 0.007905f
C355 B.n221 VSUBS 0.007905f
C356 B.n222 VSUBS 0.007905f
C357 B.n223 VSUBS 0.007905f
C358 B.n224 VSUBS 0.007905f
C359 B.n225 VSUBS 0.007905f
C360 B.n226 VSUBS 0.007905f
C361 B.n227 VSUBS 0.007905f
C362 B.n228 VSUBS 0.007905f
C363 B.n229 VSUBS 0.007905f
C364 B.n230 VSUBS 0.007905f
C365 B.n231 VSUBS 0.007905f
C366 B.n232 VSUBS 0.007905f
C367 B.n233 VSUBS 0.007905f
C368 B.n234 VSUBS 0.007905f
C369 B.n235 VSUBS 0.007905f
C370 B.n236 VSUBS 0.007905f
C371 B.n237 VSUBS 0.007905f
C372 B.n238 VSUBS 0.007905f
C373 B.n239 VSUBS 0.007905f
C374 B.n240 VSUBS 0.007905f
C375 B.n241 VSUBS 0.007905f
C376 B.n242 VSUBS 0.007905f
C377 B.n243 VSUBS 0.007905f
C378 B.n244 VSUBS 0.007905f
C379 B.n245 VSUBS 0.007905f
C380 B.n246 VSUBS 0.007905f
C381 B.n247 VSUBS 0.007905f
C382 B.n248 VSUBS 0.007905f
C383 B.n249 VSUBS 0.007905f
C384 B.n250 VSUBS 0.007905f
C385 B.n251 VSUBS 0.007905f
C386 B.n252 VSUBS 0.007905f
C387 B.n253 VSUBS 0.007905f
C388 B.n254 VSUBS 0.007905f
C389 B.n255 VSUBS 0.007905f
C390 B.n256 VSUBS 0.007905f
C391 B.n257 VSUBS 0.007905f
C392 B.n258 VSUBS 0.007905f
C393 B.n259 VSUBS 0.007905f
C394 B.n260 VSUBS 0.007905f
C395 B.n261 VSUBS 0.007905f
C396 B.n262 VSUBS 0.007905f
C397 B.n263 VSUBS 0.007905f
C398 B.n264 VSUBS 0.007905f
C399 B.n265 VSUBS 0.007905f
C400 B.n266 VSUBS 0.007905f
C401 B.n267 VSUBS 0.007905f
C402 B.n268 VSUBS 0.007905f
C403 B.n269 VSUBS 0.007905f
C404 B.n270 VSUBS 0.007905f
C405 B.n271 VSUBS 0.007905f
C406 B.n272 VSUBS 0.007905f
C407 B.n273 VSUBS 0.007905f
C408 B.n274 VSUBS 0.007905f
C409 B.n275 VSUBS 0.007905f
C410 B.n276 VSUBS 0.007905f
C411 B.n277 VSUBS 0.007905f
C412 B.n278 VSUBS 0.007905f
C413 B.n279 VSUBS 0.007905f
C414 B.n280 VSUBS 0.007905f
C415 B.n281 VSUBS 0.007905f
C416 B.n282 VSUBS 0.007905f
C417 B.n283 VSUBS 0.007905f
C418 B.n284 VSUBS 0.007905f
C419 B.n285 VSUBS 0.007905f
C420 B.n286 VSUBS 0.007905f
C421 B.n287 VSUBS 0.007905f
C422 B.n288 VSUBS 0.007905f
C423 B.n289 VSUBS 0.007905f
C424 B.n290 VSUBS 0.007905f
C425 B.n291 VSUBS 0.007905f
C426 B.n292 VSUBS 0.007905f
C427 B.n293 VSUBS 0.007905f
C428 B.n294 VSUBS 0.007905f
C429 B.n295 VSUBS 0.007905f
C430 B.n296 VSUBS 0.007905f
C431 B.n297 VSUBS 0.007905f
C432 B.n298 VSUBS 0.007905f
C433 B.n299 VSUBS 0.007905f
C434 B.n300 VSUBS 0.007905f
C435 B.n301 VSUBS 0.007905f
C436 B.n302 VSUBS 0.007905f
C437 B.n303 VSUBS 0.018654f
C438 B.n304 VSUBS 0.018654f
C439 B.n305 VSUBS 0.019711f
C440 B.n306 VSUBS 0.007905f
C441 B.n307 VSUBS 0.007905f
C442 B.n308 VSUBS 0.007905f
C443 B.n309 VSUBS 0.007905f
C444 B.n310 VSUBS 0.007905f
C445 B.n311 VSUBS 0.007905f
C446 B.n312 VSUBS 0.007905f
C447 B.n313 VSUBS 0.007905f
C448 B.n314 VSUBS 0.007905f
C449 B.n315 VSUBS 0.007905f
C450 B.n316 VSUBS 0.007905f
C451 B.n317 VSUBS 0.007905f
C452 B.n318 VSUBS 0.007905f
C453 B.n319 VSUBS 0.007905f
C454 B.n320 VSUBS 0.007905f
C455 B.n321 VSUBS 0.007905f
C456 B.n322 VSUBS 0.007905f
C457 B.n323 VSUBS 0.007905f
C458 B.n324 VSUBS 0.007905f
C459 B.n325 VSUBS 0.007905f
C460 B.n326 VSUBS 0.007905f
C461 B.n327 VSUBS 0.007905f
C462 B.n328 VSUBS 0.007905f
C463 B.n329 VSUBS 0.007905f
C464 B.n330 VSUBS 0.007905f
C465 B.n331 VSUBS 0.007905f
C466 B.n332 VSUBS 0.007905f
C467 B.n333 VSUBS 0.007905f
C468 B.n334 VSUBS 0.007905f
C469 B.n335 VSUBS 0.007905f
C470 B.n336 VSUBS 0.007905f
C471 B.n337 VSUBS 0.007905f
C472 B.n338 VSUBS 0.007905f
C473 B.n339 VSUBS 0.007905f
C474 B.n340 VSUBS 0.007905f
C475 B.n341 VSUBS 0.007905f
C476 B.n342 VSUBS 0.007905f
C477 B.n343 VSUBS 0.007905f
C478 B.n344 VSUBS 0.007905f
C479 B.n345 VSUBS 0.007905f
C480 B.n346 VSUBS 0.007905f
C481 B.n347 VSUBS 0.007905f
C482 B.n348 VSUBS 0.007905f
C483 B.n349 VSUBS 0.007905f
C484 B.n350 VSUBS 0.007905f
C485 B.n351 VSUBS 0.007905f
C486 B.n352 VSUBS 0.007905f
C487 B.n353 VSUBS 0.007905f
C488 B.n354 VSUBS 0.007905f
C489 B.n355 VSUBS 0.007905f
C490 B.n356 VSUBS 0.007905f
C491 B.n357 VSUBS 0.007905f
C492 B.n358 VSUBS 0.007905f
C493 B.n359 VSUBS 0.007905f
C494 B.n360 VSUBS 0.007905f
C495 B.n361 VSUBS 0.007905f
C496 B.n362 VSUBS 0.007905f
C497 B.n363 VSUBS 0.007905f
C498 B.n364 VSUBS 0.007905f
C499 B.n365 VSUBS 0.007905f
C500 B.n366 VSUBS 0.007905f
C501 B.n367 VSUBS 0.007905f
C502 B.n368 VSUBS 0.007905f
C503 B.n369 VSUBS 0.007905f
C504 B.n370 VSUBS 0.007905f
C505 B.n371 VSUBS 0.007905f
C506 B.n372 VSUBS 0.007905f
C507 B.n373 VSUBS 0.007905f
C508 B.n374 VSUBS 0.007905f
C509 B.n375 VSUBS 0.007905f
C510 B.n376 VSUBS 0.007905f
C511 B.n377 VSUBS 0.007905f
C512 B.n378 VSUBS 0.007905f
C513 B.n379 VSUBS 0.007905f
C514 B.n380 VSUBS 0.007905f
C515 B.n381 VSUBS 0.007905f
C516 B.n382 VSUBS 0.007905f
C517 B.n383 VSUBS 0.007905f
C518 B.n384 VSUBS 0.007905f
C519 B.n385 VSUBS 0.007905f
C520 B.n386 VSUBS 0.007905f
C521 B.n387 VSUBS 0.007905f
C522 B.n388 VSUBS 0.007905f
C523 B.n389 VSUBS 0.007905f
C524 B.n390 VSUBS 0.007905f
C525 B.n391 VSUBS 0.007905f
C526 B.n392 VSUBS 0.005464f
C527 B.n393 VSUBS 0.018316f
C528 B.n394 VSUBS 0.006394f
C529 B.n395 VSUBS 0.007905f
C530 B.n396 VSUBS 0.007905f
C531 B.n397 VSUBS 0.007905f
C532 B.n398 VSUBS 0.007905f
C533 B.n399 VSUBS 0.007905f
C534 B.n400 VSUBS 0.007905f
C535 B.n401 VSUBS 0.007905f
C536 B.n402 VSUBS 0.007905f
C537 B.n403 VSUBS 0.007905f
C538 B.n404 VSUBS 0.007905f
C539 B.n405 VSUBS 0.007905f
C540 B.n406 VSUBS 0.006394f
C541 B.n407 VSUBS 0.007905f
C542 B.n408 VSUBS 0.007905f
C543 B.n409 VSUBS 0.005464f
C544 B.n410 VSUBS 0.007905f
C545 B.n411 VSUBS 0.007905f
C546 B.n412 VSUBS 0.007905f
C547 B.n413 VSUBS 0.007905f
C548 B.n414 VSUBS 0.007905f
C549 B.n415 VSUBS 0.007905f
C550 B.n416 VSUBS 0.007905f
C551 B.n417 VSUBS 0.007905f
C552 B.n418 VSUBS 0.007905f
C553 B.n419 VSUBS 0.007905f
C554 B.n420 VSUBS 0.007905f
C555 B.n421 VSUBS 0.007905f
C556 B.n422 VSUBS 0.007905f
C557 B.n423 VSUBS 0.007905f
C558 B.n424 VSUBS 0.007905f
C559 B.n425 VSUBS 0.007905f
C560 B.n426 VSUBS 0.007905f
C561 B.n427 VSUBS 0.007905f
C562 B.n428 VSUBS 0.007905f
C563 B.n429 VSUBS 0.007905f
C564 B.n430 VSUBS 0.007905f
C565 B.n431 VSUBS 0.007905f
C566 B.n432 VSUBS 0.007905f
C567 B.n433 VSUBS 0.007905f
C568 B.n434 VSUBS 0.007905f
C569 B.n435 VSUBS 0.007905f
C570 B.n436 VSUBS 0.007905f
C571 B.n437 VSUBS 0.007905f
C572 B.n438 VSUBS 0.007905f
C573 B.n439 VSUBS 0.007905f
C574 B.n440 VSUBS 0.007905f
C575 B.n441 VSUBS 0.007905f
C576 B.n442 VSUBS 0.007905f
C577 B.n443 VSUBS 0.007905f
C578 B.n444 VSUBS 0.007905f
C579 B.n445 VSUBS 0.007905f
C580 B.n446 VSUBS 0.007905f
C581 B.n447 VSUBS 0.007905f
C582 B.n448 VSUBS 0.007905f
C583 B.n449 VSUBS 0.007905f
C584 B.n450 VSUBS 0.007905f
C585 B.n451 VSUBS 0.007905f
C586 B.n452 VSUBS 0.007905f
C587 B.n453 VSUBS 0.007905f
C588 B.n454 VSUBS 0.007905f
C589 B.n455 VSUBS 0.007905f
C590 B.n456 VSUBS 0.007905f
C591 B.n457 VSUBS 0.007905f
C592 B.n458 VSUBS 0.007905f
C593 B.n459 VSUBS 0.007905f
C594 B.n460 VSUBS 0.007905f
C595 B.n461 VSUBS 0.007905f
C596 B.n462 VSUBS 0.007905f
C597 B.n463 VSUBS 0.007905f
C598 B.n464 VSUBS 0.007905f
C599 B.n465 VSUBS 0.007905f
C600 B.n466 VSUBS 0.007905f
C601 B.n467 VSUBS 0.007905f
C602 B.n468 VSUBS 0.007905f
C603 B.n469 VSUBS 0.007905f
C604 B.n470 VSUBS 0.007905f
C605 B.n471 VSUBS 0.007905f
C606 B.n472 VSUBS 0.007905f
C607 B.n473 VSUBS 0.007905f
C608 B.n474 VSUBS 0.007905f
C609 B.n475 VSUBS 0.007905f
C610 B.n476 VSUBS 0.007905f
C611 B.n477 VSUBS 0.007905f
C612 B.n478 VSUBS 0.007905f
C613 B.n479 VSUBS 0.007905f
C614 B.n480 VSUBS 0.007905f
C615 B.n481 VSUBS 0.007905f
C616 B.n482 VSUBS 0.007905f
C617 B.n483 VSUBS 0.007905f
C618 B.n484 VSUBS 0.007905f
C619 B.n485 VSUBS 0.007905f
C620 B.n486 VSUBS 0.007905f
C621 B.n487 VSUBS 0.007905f
C622 B.n488 VSUBS 0.007905f
C623 B.n489 VSUBS 0.007905f
C624 B.n490 VSUBS 0.007905f
C625 B.n491 VSUBS 0.007905f
C626 B.n492 VSUBS 0.007905f
C627 B.n493 VSUBS 0.007905f
C628 B.n494 VSUBS 0.007905f
C629 B.n495 VSUBS 0.019711f
C630 B.n496 VSUBS 0.019711f
C631 B.n497 VSUBS 0.018654f
C632 B.n498 VSUBS 0.007905f
C633 B.n499 VSUBS 0.007905f
C634 B.n500 VSUBS 0.007905f
C635 B.n501 VSUBS 0.007905f
C636 B.n502 VSUBS 0.007905f
C637 B.n503 VSUBS 0.007905f
C638 B.n504 VSUBS 0.007905f
C639 B.n505 VSUBS 0.007905f
C640 B.n506 VSUBS 0.007905f
C641 B.n507 VSUBS 0.007905f
C642 B.n508 VSUBS 0.007905f
C643 B.n509 VSUBS 0.007905f
C644 B.n510 VSUBS 0.007905f
C645 B.n511 VSUBS 0.007905f
C646 B.n512 VSUBS 0.007905f
C647 B.n513 VSUBS 0.007905f
C648 B.n514 VSUBS 0.007905f
C649 B.n515 VSUBS 0.007905f
C650 B.n516 VSUBS 0.007905f
C651 B.n517 VSUBS 0.007905f
C652 B.n518 VSUBS 0.007905f
C653 B.n519 VSUBS 0.007905f
C654 B.n520 VSUBS 0.007905f
C655 B.n521 VSUBS 0.007905f
C656 B.n522 VSUBS 0.007905f
C657 B.n523 VSUBS 0.007905f
C658 B.n524 VSUBS 0.007905f
C659 B.n525 VSUBS 0.007905f
C660 B.n526 VSUBS 0.007905f
C661 B.n527 VSUBS 0.007905f
C662 B.n528 VSUBS 0.007905f
C663 B.n529 VSUBS 0.007905f
C664 B.n530 VSUBS 0.007905f
C665 B.n531 VSUBS 0.007905f
C666 B.n532 VSUBS 0.007905f
C667 B.n533 VSUBS 0.007905f
C668 B.n534 VSUBS 0.007905f
C669 B.n535 VSUBS 0.007905f
C670 B.n536 VSUBS 0.007905f
C671 B.n537 VSUBS 0.007905f
C672 B.n538 VSUBS 0.007905f
C673 B.n539 VSUBS 0.007905f
C674 B.n540 VSUBS 0.007905f
C675 B.n541 VSUBS 0.007905f
C676 B.n542 VSUBS 0.007905f
C677 B.n543 VSUBS 0.007905f
C678 B.n544 VSUBS 0.007905f
C679 B.n545 VSUBS 0.007905f
C680 B.n546 VSUBS 0.007905f
C681 B.n547 VSUBS 0.007905f
C682 B.n548 VSUBS 0.007905f
C683 B.n549 VSUBS 0.007905f
C684 B.n550 VSUBS 0.007905f
C685 B.n551 VSUBS 0.007905f
C686 B.n552 VSUBS 0.007905f
C687 B.n553 VSUBS 0.007905f
C688 B.n554 VSUBS 0.007905f
C689 B.n555 VSUBS 0.007905f
C690 B.n556 VSUBS 0.007905f
C691 B.n557 VSUBS 0.007905f
C692 B.n558 VSUBS 0.007905f
C693 B.n559 VSUBS 0.007905f
C694 B.n560 VSUBS 0.007905f
C695 B.n561 VSUBS 0.007905f
C696 B.n562 VSUBS 0.007905f
C697 B.n563 VSUBS 0.007905f
C698 B.n564 VSUBS 0.007905f
C699 B.n565 VSUBS 0.007905f
C700 B.n566 VSUBS 0.007905f
C701 B.n567 VSUBS 0.007905f
C702 B.n568 VSUBS 0.007905f
C703 B.n569 VSUBS 0.007905f
C704 B.n570 VSUBS 0.007905f
C705 B.n571 VSUBS 0.007905f
C706 B.n572 VSUBS 0.007905f
C707 B.n573 VSUBS 0.007905f
C708 B.n574 VSUBS 0.007905f
C709 B.n575 VSUBS 0.007905f
C710 B.n576 VSUBS 0.007905f
C711 B.n577 VSUBS 0.007905f
C712 B.n578 VSUBS 0.007905f
C713 B.n579 VSUBS 0.007905f
C714 B.n580 VSUBS 0.007905f
C715 B.n581 VSUBS 0.007905f
C716 B.n582 VSUBS 0.007905f
C717 B.n583 VSUBS 0.007905f
C718 B.n584 VSUBS 0.007905f
C719 B.n585 VSUBS 0.007905f
C720 B.n586 VSUBS 0.007905f
C721 B.n587 VSUBS 0.007905f
C722 B.n588 VSUBS 0.007905f
C723 B.n589 VSUBS 0.007905f
C724 B.n590 VSUBS 0.007905f
C725 B.n591 VSUBS 0.007905f
C726 B.n592 VSUBS 0.007905f
C727 B.n593 VSUBS 0.007905f
C728 B.n594 VSUBS 0.007905f
C729 B.n595 VSUBS 0.007905f
C730 B.n596 VSUBS 0.007905f
C731 B.n597 VSUBS 0.007905f
C732 B.n598 VSUBS 0.007905f
C733 B.n599 VSUBS 0.007905f
C734 B.n600 VSUBS 0.007905f
C735 B.n601 VSUBS 0.007905f
C736 B.n602 VSUBS 0.007905f
C737 B.n603 VSUBS 0.007905f
C738 B.n604 VSUBS 0.007905f
C739 B.n605 VSUBS 0.007905f
C740 B.n606 VSUBS 0.007905f
C741 B.n607 VSUBS 0.007905f
C742 B.n608 VSUBS 0.007905f
C743 B.n609 VSUBS 0.007905f
C744 B.n610 VSUBS 0.007905f
C745 B.n611 VSUBS 0.007905f
C746 B.n612 VSUBS 0.007905f
C747 B.n613 VSUBS 0.007905f
C748 B.n614 VSUBS 0.007905f
C749 B.n615 VSUBS 0.007905f
C750 B.n616 VSUBS 0.007905f
C751 B.n617 VSUBS 0.007905f
C752 B.n618 VSUBS 0.007905f
C753 B.n619 VSUBS 0.007905f
C754 B.n620 VSUBS 0.007905f
C755 B.n621 VSUBS 0.007905f
C756 B.n622 VSUBS 0.007905f
C757 B.n623 VSUBS 0.007905f
C758 B.n624 VSUBS 0.007905f
C759 B.n625 VSUBS 0.007905f
C760 B.n626 VSUBS 0.007905f
C761 B.n627 VSUBS 0.007905f
C762 B.n628 VSUBS 0.007905f
C763 B.n629 VSUBS 0.007905f
C764 B.n630 VSUBS 0.007905f
C765 B.n631 VSUBS 0.007905f
C766 B.n632 VSUBS 0.007905f
C767 B.n633 VSUBS 0.007905f
C768 B.n634 VSUBS 0.007905f
C769 B.n635 VSUBS 0.007905f
C770 B.n636 VSUBS 0.007905f
C771 B.n637 VSUBS 0.007905f
C772 B.n638 VSUBS 0.007905f
C773 B.n639 VSUBS 0.007905f
C774 B.n640 VSUBS 0.007905f
C775 B.n641 VSUBS 0.018654f
C776 B.n642 VSUBS 0.019711f
C777 B.n643 VSUBS 0.018826f
C778 B.n644 VSUBS 0.007905f
C779 B.n645 VSUBS 0.007905f
C780 B.n646 VSUBS 0.007905f
C781 B.n647 VSUBS 0.007905f
C782 B.n648 VSUBS 0.007905f
C783 B.n649 VSUBS 0.007905f
C784 B.n650 VSUBS 0.007905f
C785 B.n651 VSUBS 0.007905f
C786 B.n652 VSUBS 0.007905f
C787 B.n653 VSUBS 0.007905f
C788 B.n654 VSUBS 0.007905f
C789 B.n655 VSUBS 0.007905f
C790 B.n656 VSUBS 0.007905f
C791 B.n657 VSUBS 0.007905f
C792 B.n658 VSUBS 0.007905f
C793 B.n659 VSUBS 0.007905f
C794 B.n660 VSUBS 0.007905f
C795 B.n661 VSUBS 0.007905f
C796 B.n662 VSUBS 0.007905f
C797 B.n663 VSUBS 0.007905f
C798 B.n664 VSUBS 0.007905f
C799 B.n665 VSUBS 0.007905f
C800 B.n666 VSUBS 0.007905f
C801 B.n667 VSUBS 0.007905f
C802 B.n668 VSUBS 0.007905f
C803 B.n669 VSUBS 0.007905f
C804 B.n670 VSUBS 0.007905f
C805 B.n671 VSUBS 0.007905f
C806 B.n672 VSUBS 0.007905f
C807 B.n673 VSUBS 0.007905f
C808 B.n674 VSUBS 0.007905f
C809 B.n675 VSUBS 0.007905f
C810 B.n676 VSUBS 0.007905f
C811 B.n677 VSUBS 0.007905f
C812 B.n678 VSUBS 0.007905f
C813 B.n679 VSUBS 0.007905f
C814 B.n680 VSUBS 0.007905f
C815 B.n681 VSUBS 0.007905f
C816 B.n682 VSUBS 0.007905f
C817 B.n683 VSUBS 0.007905f
C818 B.n684 VSUBS 0.007905f
C819 B.n685 VSUBS 0.007905f
C820 B.n686 VSUBS 0.007905f
C821 B.n687 VSUBS 0.007905f
C822 B.n688 VSUBS 0.007905f
C823 B.n689 VSUBS 0.007905f
C824 B.n690 VSUBS 0.007905f
C825 B.n691 VSUBS 0.007905f
C826 B.n692 VSUBS 0.007905f
C827 B.n693 VSUBS 0.007905f
C828 B.n694 VSUBS 0.007905f
C829 B.n695 VSUBS 0.007905f
C830 B.n696 VSUBS 0.007905f
C831 B.n697 VSUBS 0.007905f
C832 B.n698 VSUBS 0.007905f
C833 B.n699 VSUBS 0.007905f
C834 B.n700 VSUBS 0.007905f
C835 B.n701 VSUBS 0.007905f
C836 B.n702 VSUBS 0.007905f
C837 B.n703 VSUBS 0.007905f
C838 B.n704 VSUBS 0.007905f
C839 B.n705 VSUBS 0.007905f
C840 B.n706 VSUBS 0.007905f
C841 B.n707 VSUBS 0.007905f
C842 B.n708 VSUBS 0.007905f
C843 B.n709 VSUBS 0.007905f
C844 B.n710 VSUBS 0.007905f
C845 B.n711 VSUBS 0.007905f
C846 B.n712 VSUBS 0.007905f
C847 B.n713 VSUBS 0.007905f
C848 B.n714 VSUBS 0.007905f
C849 B.n715 VSUBS 0.007905f
C850 B.n716 VSUBS 0.007905f
C851 B.n717 VSUBS 0.007905f
C852 B.n718 VSUBS 0.007905f
C853 B.n719 VSUBS 0.007905f
C854 B.n720 VSUBS 0.007905f
C855 B.n721 VSUBS 0.007905f
C856 B.n722 VSUBS 0.007905f
C857 B.n723 VSUBS 0.007905f
C858 B.n724 VSUBS 0.007905f
C859 B.n725 VSUBS 0.007905f
C860 B.n726 VSUBS 0.007905f
C861 B.n727 VSUBS 0.007905f
C862 B.n728 VSUBS 0.007905f
C863 B.n729 VSUBS 0.005464f
C864 B.n730 VSUBS 0.007905f
C865 B.n731 VSUBS 0.007905f
C866 B.n732 VSUBS 0.006394f
C867 B.n733 VSUBS 0.007905f
C868 B.n734 VSUBS 0.007905f
C869 B.n735 VSUBS 0.007905f
C870 B.n736 VSUBS 0.007905f
C871 B.n737 VSUBS 0.007905f
C872 B.n738 VSUBS 0.007905f
C873 B.n739 VSUBS 0.007905f
C874 B.n740 VSUBS 0.007905f
C875 B.n741 VSUBS 0.007905f
C876 B.n742 VSUBS 0.007905f
C877 B.n743 VSUBS 0.007905f
C878 B.n744 VSUBS 0.006394f
C879 B.n745 VSUBS 0.018316f
C880 B.n746 VSUBS 0.005464f
C881 B.n747 VSUBS 0.007905f
C882 B.n748 VSUBS 0.007905f
C883 B.n749 VSUBS 0.007905f
C884 B.n750 VSUBS 0.007905f
C885 B.n751 VSUBS 0.007905f
C886 B.n752 VSUBS 0.007905f
C887 B.n753 VSUBS 0.007905f
C888 B.n754 VSUBS 0.007905f
C889 B.n755 VSUBS 0.007905f
C890 B.n756 VSUBS 0.007905f
C891 B.n757 VSUBS 0.007905f
C892 B.n758 VSUBS 0.007905f
C893 B.n759 VSUBS 0.007905f
C894 B.n760 VSUBS 0.007905f
C895 B.n761 VSUBS 0.007905f
C896 B.n762 VSUBS 0.007905f
C897 B.n763 VSUBS 0.007905f
C898 B.n764 VSUBS 0.007905f
C899 B.n765 VSUBS 0.007905f
C900 B.n766 VSUBS 0.007905f
C901 B.n767 VSUBS 0.007905f
C902 B.n768 VSUBS 0.007905f
C903 B.n769 VSUBS 0.007905f
C904 B.n770 VSUBS 0.007905f
C905 B.n771 VSUBS 0.007905f
C906 B.n772 VSUBS 0.007905f
C907 B.n773 VSUBS 0.007905f
C908 B.n774 VSUBS 0.007905f
C909 B.n775 VSUBS 0.007905f
C910 B.n776 VSUBS 0.007905f
C911 B.n777 VSUBS 0.007905f
C912 B.n778 VSUBS 0.007905f
C913 B.n779 VSUBS 0.007905f
C914 B.n780 VSUBS 0.007905f
C915 B.n781 VSUBS 0.007905f
C916 B.n782 VSUBS 0.007905f
C917 B.n783 VSUBS 0.007905f
C918 B.n784 VSUBS 0.007905f
C919 B.n785 VSUBS 0.007905f
C920 B.n786 VSUBS 0.007905f
C921 B.n787 VSUBS 0.007905f
C922 B.n788 VSUBS 0.007905f
C923 B.n789 VSUBS 0.007905f
C924 B.n790 VSUBS 0.007905f
C925 B.n791 VSUBS 0.007905f
C926 B.n792 VSUBS 0.007905f
C927 B.n793 VSUBS 0.007905f
C928 B.n794 VSUBS 0.007905f
C929 B.n795 VSUBS 0.007905f
C930 B.n796 VSUBS 0.007905f
C931 B.n797 VSUBS 0.007905f
C932 B.n798 VSUBS 0.007905f
C933 B.n799 VSUBS 0.007905f
C934 B.n800 VSUBS 0.007905f
C935 B.n801 VSUBS 0.007905f
C936 B.n802 VSUBS 0.007905f
C937 B.n803 VSUBS 0.007905f
C938 B.n804 VSUBS 0.007905f
C939 B.n805 VSUBS 0.007905f
C940 B.n806 VSUBS 0.007905f
C941 B.n807 VSUBS 0.007905f
C942 B.n808 VSUBS 0.007905f
C943 B.n809 VSUBS 0.007905f
C944 B.n810 VSUBS 0.007905f
C945 B.n811 VSUBS 0.007905f
C946 B.n812 VSUBS 0.007905f
C947 B.n813 VSUBS 0.007905f
C948 B.n814 VSUBS 0.007905f
C949 B.n815 VSUBS 0.007905f
C950 B.n816 VSUBS 0.007905f
C951 B.n817 VSUBS 0.007905f
C952 B.n818 VSUBS 0.007905f
C953 B.n819 VSUBS 0.007905f
C954 B.n820 VSUBS 0.007905f
C955 B.n821 VSUBS 0.007905f
C956 B.n822 VSUBS 0.007905f
C957 B.n823 VSUBS 0.007905f
C958 B.n824 VSUBS 0.007905f
C959 B.n825 VSUBS 0.007905f
C960 B.n826 VSUBS 0.007905f
C961 B.n827 VSUBS 0.007905f
C962 B.n828 VSUBS 0.007905f
C963 B.n829 VSUBS 0.007905f
C964 B.n830 VSUBS 0.007905f
C965 B.n831 VSUBS 0.007905f
C966 B.n832 VSUBS 0.007905f
C967 B.n833 VSUBS 0.019711f
C968 B.n834 VSUBS 0.018654f
C969 B.n835 VSUBS 0.018654f
C970 B.n836 VSUBS 0.007905f
C971 B.n837 VSUBS 0.007905f
C972 B.n838 VSUBS 0.007905f
C973 B.n839 VSUBS 0.007905f
C974 B.n840 VSUBS 0.007905f
C975 B.n841 VSUBS 0.007905f
C976 B.n842 VSUBS 0.007905f
C977 B.n843 VSUBS 0.007905f
C978 B.n844 VSUBS 0.007905f
C979 B.n845 VSUBS 0.007905f
C980 B.n846 VSUBS 0.007905f
C981 B.n847 VSUBS 0.007905f
C982 B.n848 VSUBS 0.007905f
C983 B.n849 VSUBS 0.007905f
C984 B.n850 VSUBS 0.007905f
C985 B.n851 VSUBS 0.007905f
C986 B.n852 VSUBS 0.007905f
C987 B.n853 VSUBS 0.007905f
C988 B.n854 VSUBS 0.007905f
C989 B.n855 VSUBS 0.007905f
C990 B.n856 VSUBS 0.007905f
C991 B.n857 VSUBS 0.007905f
C992 B.n858 VSUBS 0.007905f
C993 B.n859 VSUBS 0.007905f
C994 B.n860 VSUBS 0.007905f
C995 B.n861 VSUBS 0.007905f
C996 B.n862 VSUBS 0.007905f
C997 B.n863 VSUBS 0.007905f
C998 B.n864 VSUBS 0.007905f
C999 B.n865 VSUBS 0.007905f
C1000 B.n866 VSUBS 0.007905f
C1001 B.n867 VSUBS 0.007905f
C1002 B.n868 VSUBS 0.007905f
C1003 B.n869 VSUBS 0.007905f
C1004 B.n870 VSUBS 0.007905f
C1005 B.n871 VSUBS 0.007905f
C1006 B.n872 VSUBS 0.007905f
C1007 B.n873 VSUBS 0.007905f
C1008 B.n874 VSUBS 0.007905f
C1009 B.n875 VSUBS 0.007905f
C1010 B.n876 VSUBS 0.007905f
C1011 B.n877 VSUBS 0.007905f
C1012 B.n878 VSUBS 0.007905f
C1013 B.n879 VSUBS 0.007905f
C1014 B.n880 VSUBS 0.007905f
C1015 B.n881 VSUBS 0.007905f
C1016 B.n882 VSUBS 0.007905f
C1017 B.n883 VSUBS 0.007905f
C1018 B.n884 VSUBS 0.007905f
C1019 B.n885 VSUBS 0.007905f
C1020 B.n886 VSUBS 0.007905f
C1021 B.n887 VSUBS 0.007905f
C1022 B.n888 VSUBS 0.007905f
C1023 B.n889 VSUBS 0.007905f
C1024 B.n890 VSUBS 0.007905f
C1025 B.n891 VSUBS 0.007905f
C1026 B.n892 VSUBS 0.007905f
C1027 B.n893 VSUBS 0.007905f
C1028 B.n894 VSUBS 0.007905f
C1029 B.n895 VSUBS 0.007905f
C1030 B.n896 VSUBS 0.007905f
C1031 B.n897 VSUBS 0.007905f
C1032 B.n898 VSUBS 0.007905f
C1033 B.n899 VSUBS 0.007905f
C1034 B.n900 VSUBS 0.007905f
C1035 B.n901 VSUBS 0.007905f
C1036 B.n902 VSUBS 0.007905f
C1037 B.n903 VSUBS 0.007905f
C1038 B.n904 VSUBS 0.007905f
C1039 B.n905 VSUBS 0.007905f
C1040 B.n906 VSUBS 0.007905f
C1041 B.n907 VSUBS 0.0179f
C1042 VDD1.t8 VSUBS 4.04271f
C1043 VDD1.t5 VSUBS 0.374211f
C1044 VDD1.t3 VSUBS 0.374211f
C1045 VDD1.n0 VSUBS 3.09832f
C1046 VDD1.n1 VSUBS 1.52884f
C1047 VDD1.t9 VSUBS 4.04271f
C1048 VDD1.t2 VSUBS 0.374211f
C1049 VDD1.t4 VSUBS 0.374211f
C1050 VDD1.n2 VSUBS 3.09832f
C1051 VDD1.n3 VSUBS 1.52055f
C1052 VDD1.t6 VSUBS 0.374211f
C1053 VDD1.t0 VSUBS 0.374211f
C1054 VDD1.n4 VSUBS 3.11527f
C1055 VDD1.n5 VSUBS 3.52988f
C1056 VDD1.t1 VSUBS 0.374211f
C1057 VDD1.t7 VSUBS 0.374211f
C1058 VDD1.n6 VSUBS 3.09831f
C1059 VDD1.n7 VSUBS 3.86384f
C1060 VTAIL.t0 VSUBS 0.381432f
C1061 VTAIL.t1 VSUBS 0.381432f
C1062 VTAIL.n0 VSUBS 2.98315f
C1063 VTAIL.n1 VSUBS 0.937927f
C1064 VTAIL.t8 VSUBS 3.89767f
C1065 VTAIL.n2 VSUBS 1.10129f
C1066 VTAIL.t13 VSUBS 0.381432f
C1067 VTAIL.t10 VSUBS 0.381432f
C1068 VTAIL.n3 VSUBS 2.98315f
C1069 VTAIL.n4 VSUBS 1.01994f
C1070 VTAIL.t16 VSUBS 0.381432f
C1071 VTAIL.t7 VSUBS 0.381432f
C1072 VTAIL.n5 VSUBS 2.98315f
C1073 VTAIL.n6 VSUBS 2.89947f
C1074 VTAIL.t2 VSUBS 0.381432f
C1075 VTAIL.t17 VSUBS 0.381432f
C1076 VTAIL.n7 VSUBS 2.98315f
C1077 VTAIL.n8 VSUBS 2.89946f
C1078 VTAIL.t4 VSUBS 0.381432f
C1079 VTAIL.t6 VSUBS 0.381432f
C1080 VTAIL.n9 VSUBS 2.98315f
C1081 VTAIL.n10 VSUBS 1.01993f
C1082 VTAIL.t19 VSUBS 3.89768f
C1083 VTAIL.n11 VSUBS 1.10128f
C1084 VTAIL.t15 VSUBS 0.381432f
C1085 VTAIL.t14 VSUBS 0.381432f
C1086 VTAIL.n12 VSUBS 2.98315f
C1087 VTAIL.n13 VSUBS 0.975541f
C1088 VTAIL.t12 VSUBS 0.381432f
C1089 VTAIL.t9 VSUBS 0.381432f
C1090 VTAIL.n14 VSUBS 2.98315f
C1091 VTAIL.n15 VSUBS 1.01993f
C1092 VTAIL.t11 VSUBS 3.89767f
C1093 VTAIL.n16 VSUBS 2.85442f
C1094 VTAIL.t3 VSUBS 3.89767f
C1095 VTAIL.n17 VSUBS 2.85442f
C1096 VTAIL.t5 VSUBS 0.381432f
C1097 VTAIL.t18 VSUBS 0.381432f
C1098 VTAIL.n18 VSUBS 2.98315f
C1099 VTAIL.n19 VSUBS 0.886764f
C1100 VP.n0 VSUBS 0.030697f
C1101 VP.t9 VSUBS 2.9184f
C1102 VP.n1 VSUBS 0.028516f
C1103 VP.n2 VSUBS 0.030697f
C1104 VP.t3 VSUBS 2.9184f
C1105 VP.n3 VSUBS 0.05388f
C1106 VP.n4 VSUBS 0.030697f
C1107 VP.t5 VSUBS 2.9184f
C1108 VP.n5 VSUBS 0.059538f
C1109 VP.n6 VSUBS 0.030697f
C1110 VP.t7 VSUBS 2.9184f
C1111 VP.n7 VSUBS 1.01945f
C1112 VP.n8 VSUBS 0.030697f
C1113 VP.n9 VSUBS 0.061298f
C1114 VP.n10 VSUBS 0.030697f
C1115 VP.t2 VSUBS 2.9184f
C1116 VP.n11 VSUBS 0.028516f
C1117 VP.n12 VSUBS 0.030697f
C1118 VP.t8 VSUBS 2.9184f
C1119 VP.n13 VSUBS 0.05388f
C1120 VP.n14 VSUBS 0.030697f
C1121 VP.t6 VSUBS 2.9184f
C1122 VP.n15 VSUBS 0.059538f
C1123 VP.n16 VSUBS 0.030697f
C1124 VP.t4 VSUBS 2.9184f
C1125 VP.n17 VSUBS 1.09193f
C1126 VP.t1 VSUBS 3.06991f
C1127 VP.n18 VSUBS 1.09429f
C1128 VP.n19 VSUBS 0.228782f
C1129 VP.n20 VSUBS 0.043998f
C1130 VP.n21 VSUBS 0.05388f
C1131 VP.n22 VSUBS 0.032751f
C1132 VP.n23 VSUBS 0.030697f
C1133 VP.n24 VSUBS 0.030697f
C1134 VP.n25 VSUBS 0.030697f
C1135 VP.n26 VSUBS 1.04827f
C1136 VP.n27 VSUBS 0.059538f
C1137 VP.n28 VSUBS 0.032751f
C1138 VP.n29 VSUBS 0.030697f
C1139 VP.n30 VSUBS 0.030697f
C1140 VP.n31 VSUBS 0.030697f
C1141 VP.n32 VSUBS 0.043998f
C1142 VP.n33 VSUBS 1.01945f
C1143 VP.n34 VSUBS 0.041749f
C1144 VP.n35 VSUBS 0.056356f
C1145 VP.n36 VSUBS 0.030697f
C1146 VP.n37 VSUBS 0.030697f
C1147 VP.n38 VSUBS 0.030697f
C1148 VP.n39 VSUBS 0.061298f
C1149 VP.n40 VSUBS 0.031071f
C1150 VP.n41 VSUBS 1.09303f
C1151 VP.n42 VSUBS 1.8721f
C1152 VP.n43 VSUBS 1.89265f
C1153 VP.t0 VSUBS 2.9184f
C1154 VP.n44 VSUBS 1.09303f
C1155 VP.n45 VSUBS 0.031071f
C1156 VP.n46 VSUBS 0.030697f
C1157 VP.n47 VSUBS 0.030697f
C1158 VP.n48 VSUBS 0.030697f
C1159 VP.n49 VSUBS 0.028516f
C1160 VP.n50 VSUBS 0.056356f
C1161 VP.n51 VSUBS 0.041749f
C1162 VP.n52 VSUBS 0.030697f
C1163 VP.n53 VSUBS 0.030697f
C1164 VP.n54 VSUBS 0.043998f
C1165 VP.n55 VSUBS 0.05388f
C1166 VP.n56 VSUBS 0.032751f
C1167 VP.n57 VSUBS 0.030697f
C1168 VP.n58 VSUBS 0.030697f
C1169 VP.n59 VSUBS 0.030697f
C1170 VP.n60 VSUBS 1.04827f
C1171 VP.n61 VSUBS 0.059538f
C1172 VP.n62 VSUBS 0.032751f
C1173 VP.n63 VSUBS 0.030697f
C1174 VP.n64 VSUBS 0.030697f
C1175 VP.n65 VSUBS 0.030697f
C1176 VP.n66 VSUBS 0.043998f
C1177 VP.n67 VSUBS 1.01945f
C1178 VP.n68 VSUBS 0.041749f
C1179 VP.n69 VSUBS 0.056356f
C1180 VP.n70 VSUBS 0.030697f
C1181 VP.n71 VSUBS 0.030697f
C1182 VP.n72 VSUBS 0.030697f
C1183 VP.n73 VSUBS 0.061298f
C1184 VP.n74 VSUBS 0.031071f
C1185 VP.n75 VSUBS 1.09303f
C1186 VP.n76 VSUBS 0.03411f
.ends

