* NGSPICE file created from diff_pair_sample_1046.ext - technology: sky130A

.subckt diff_pair_sample_1046 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.3861 pd=2.76 as=0.16335 ps=1.32 w=0.99 l=3.81
X1 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=0.3861 pd=2.76 as=0 ps=0 w=0.99 l=3.81
X2 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=0.3861 pd=2.76 as=0 ps=0 w=0.99 l=3.81
X3 VDD2.t0 VN.t1 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.16335 pd=1.32 as=0.3861 ps=2.76 w=0.99 l=3.81
X4 VTAIL.t1 VP.t0 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3861 pd=2.76 as=0.16335 ps=1.32 w=0.99 l=3.81
X5 VTAIL.t2 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.3861 pd=2.76 as=0.16335 ps=1.32 w=0.99 l=3.81
X6 VDD2.t2 VN.t2 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=0.16335 pd=1.32 as=0.3861 ps=2.76 w=0.99 l=3.81
X7 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=0.3861 pd=2.76 as=0 ps=0 w=0.99 l=3.81
X8 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.3861 pd=2.76 as=0 ps=0 w=0.99 l=3.81
X9 VTAIL.t4 VN.t3 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3861 pd=2.76 as=0.16335 ps=1.32 w=0.99 l=3.81
X10 VDD1.t1 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.16335 pd=1.32 as=0.3861 ps=2.76 w=0.99 l=3.81
X11 VDD1.t0 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.16335 pd=1.32 as=0.3861 ps=2.76 w=0.99 l=3.81
R0 VN VN.n1 43.7552
R1 VN.n1 VN.t2 40.2664
R2 VN.n0 VN.t3 40.2664
R3 VN.n1 VN.t0 38.9138
R4 VN.n0 VN.t1 38.9138
R5 VN VN.n0 1.84986
R6 VDD2.n2 VDD2.n0 275.214
R7 VDD2.n2 VDD2.n1 239.939
R8 VDD2.n1 VDD2.t3 20.0005
R9 VDD2.n1 VDD2.t2 20.0005
R10 VDD2.n0 VDD2.t1 20.0005
R11 VDD2.n0 VDD2.t0 20.0005
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n6 VTAIL.t0 243.261
R14 VTAIL.n5 VTAIL.t1 243.261
R15 VTAIL.n4 VTAIL.t5 243.261
R16 VTAIL.n3 VTAIL.t7 243.261
R17 VTAIL.n7 VTAIL.t6 243.26
R18 VTAIL.n0 VTAIL.t4 243.26
R19 VTAIL.n1 VTAIL.t3 243.26
R20 VTAIL.n2 VTAIL.t2 243.26
R21 VTAIL.n7 VTAIL.n6 16.7893
R22 VTAIL.n3 VTAIL.n2 16.7893
R23 VTAIL.n4 VTAIL.n3 3.56947
R24 VTAIL.n6 VTAIL.n5 3.56947
R25 VTAIL.n2 VTAIL.n1 3.56947
R26 VTAIL VTAIL.n0 1.84317
R27 VTAIL VTAIL.n7 1.72679
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 B.n507 B.n506 585
R31 B.n154 B.n97 585
R32 B.n153 B.n152 585
R33 B.n151 B.n150 585
R34 B.n149 B.n148 585
R35 B.n147 B.n146 585
R36 B.n145 B.n144 585
R37 B.n143 B.n142 585
R38 B.n141 B.n140 585
R39 B.n138 B.n137 585
R40 B.n136 B.n135 585
R41 B.n134 B.n133 585
R42 B.n132 B.n131 585
R43 B.n130 B.n129 585
R44 B.n128 B.n127 585
R45 B.n126 B.n125 585
R46 B.n124 B.n123 585
R47 B.n122 B.n121 585
R48 B.n120 B.n119 585
R49 B.n117 B.n116 585
R50 B.n115 B.n114 585
R51 B.n113 B.n112 585
R52 B.n111 B.n110 585
R53 B.n109 B.n108 585
R54 B.n107 B.n106 585
R55 B.n105 B.n104 585
R56 B.n103 B.n102 585
R57 B.n82 B.n81 585
R58 B.n505 B.n83 585
R59 B.n510 B.n83 585
R60 B.n504 B.n503 585
R61 B.n503 B.n79 585
R62 B.n502 B.n78 585
R63 B.n516 B.n78 585
R64 B.n501 B.n77 585
R65 B.n517 B.n77 585
R66 B.n500 B.n76 585
R67 B.n518 B.n76 585
R68 B.n499 B.n498 585
R69 B.n498 B.n72 585
R70 B.n497 B.n71 585
R71 B.n524 B.n71 585
R72 B.n496 B.n70 585
R73 B.n525 B.n70 585
R74 B.n495 B.n69 585
R75 B.n526 B.n69 585
R76 B.n494 B.n493 585
R77 B.n493 B.n68 585
R78 B.n492 B.n64 585
R79 B.n532 B.n64 585
R80 B.n491 B.n63 585
R81 B.n533 B.n63 585
R82 B.n490 B.n62 585
R83 B.n534 B.n62 585
R84 B.n489 B.n488 585
R85 B.n488 B.n58 585
R86 B.n487 B.n57 585
R87 B.n540 B.n57 585
R88 B.n486 B.n56 585
R89 B.n541 B.n56 585
R90 B.n485 B.n55 585
R91 B.n542 B.n55 585
R92 B.n484 B.n483 585
R93 B.n483 B.n51 585
R94 B.n482 B.n50 585
R95 B.n548 B.n50 585
R96 B.n481 B.n49 585
R97 B.n549 B.n49 585
R98 B.n480 B.n48 585
R99 B.n550 B.n48 585
R100 B.n479 B.n478 585
R101 B.n478 B.n44 585
R102 B.n477 B.n43 585
R103 B.n556 B.n43 585
R104 B.n476 B.n42 585
R105 B.n557 B.n42 585
R106 B.n475 B.n41 585
R107 B.n558 B.n41 585
R108 B.n474 B.n473 585
R109 B.n473 B.n37 585
R110 B.n472 B.n36 585
R111 B.n564 B.n36 585
R112 B.n471 B.n35 585
R113 B.n565 B.n35 585
R114 B.n470 B.n34 585
R115 B.n566 B.n34 585
R116 B.n469 B.n468 585
R117 B.n468 B.n30 585
R118 B.n467 B.n29 585
R119 B.n572 B.n29 585
R120 B.n466 B.n28 585
R121 B.n573 B.n28 585
R122 B.n465 B.n27 585
R123 B.n574 B.n27 585
R124 B.n464 B.n463 585
R125 B.n463 B.n23 585
R126 B.n462 B.n22 585
R127 B.n580 B.n22 585
R128 B.n461 B.n21 585
R129 B.n581 B.n21 585
R130 B.n460 B.n20 585
R131 B.n582 B.n20 585
R132 B.n459 B.n458 585
R133 B.n458 B.n16 585
R134 B.n457 B.n15 585
R135 B.n588 B.n15 585
R136 B.n456 B.n14 585
R137 B.n589 B.n14 585
R138 B.n455 B.n13 585
R139 B.n590 B.n13 585
R140 B.n454 B.n453 585
R141 B.n453 B.n12 585
R142 B.n452 B.n451 585
R143 B.n452 B.n8 585
R144 B.n450 B.n7 585
R145 B.n597 B.n7 585
R146 B.n449 B.n6 585
R147 B.n598 B.n6 585
R148 B.n448 B.n5 585
R149 B.n599 B.n5 585
R150 B.n447 B.n446 585
R151 B.n446 B.n4 585
R152 B.n445 B.n155 585
R153 B.n445 B.n444 585
R154 B.n435 B.n156 585
R155 B.n157 B.n156 585
R156 B.n437 B.n436 585
R157 B.n438 B.n437 585
R158 B.n434 B.n162 585
R159 B.n162 B.n161 585
R160 B.n433 B.n432 585
R161 B.n432 B.n431 585
R162 B.n164 B.n163 585
R163 B.n165 B.n164 585
R164 B.n424 B.n423 585
R165 B.n425 B.n424 585
R166 B.n422 B.n170 585
R167 B.n170 B.n169 585
R168 B.n421 B.n420 585
R169 B.n420 B.n419 585
R170 B.n172 B.n171 585
R171 B.n173 B.n172 585
R172 B.n412 B.n411 585
R173 B.n413 B.n412 585
R174 B.n410 B.n178 585
R175 B.n178 B.n177 585
R176 B.n409 B.n408 585
R177 B.n408 B.n407 585
R178 B.n180 B.n179 585
R179 B.n181 B.n180 585
R180 B.n400 B.n399 585
R181 B.n401 B.n400 585
R182 B.n398 B.n186 585
R183 B.n186 B.n185 585
R184 B.n397 B.n396 585
R185 B.n396 B.n395 585
R186 B.n188 B.n187 585
R187 B.n189 B.n188 585
R188 B.n388 B.n387 585
R189 B.n389 B.n388 585
R190 B.n386 B.n194 585
R191 B.n194 B.n193 585
R192 B.n385 B.n384 585
R193 B.n384 B.n383 585
R194 B.n196 B.n195 585
R195 B.n197 B.n196 585
R196 B.n376 B.n375 585
R197 B.n377 B.n376 585
R198 B.n374 B.n202 585
R199 B.n202 B.n201 585
R200 B.n373 B.n372 585
R201 B.n372 B.n371 585
R202 B.n204 B.n203 585
R203 B.n205 B.n204 585
R204 B.n364 B.n363 585
R205 B.n365 B.n364 585
R206 B.n362 B.n210 585
R207 B.n210 B.n209 585
R208 B.n361 B.n360 585
R209 B.n360 B.n359 585
R210 B.n212 B.n211 585
R211 B.n213 B.n212 585
R212 B.n352 B.n351 585
R213 B.n353 B.n352 585
R214 B.n350 B.n218 585
R215 B.n218 B.n217 585
R216 B.n349 B.n348 585
R217 B.n348 B.n347 585
R218 B.n220 B.n219 585
R219 B.n340 B.n220 585
R220 B.n339 B.n338 585
R221 B.n341 B.n339 585
R222 B.n337 B.n225 585
R223 B.n225 B.n224 585
R224 B.n336 B.n335 585
R225 B.n335 B.n334 585
R226 B.n227 B.n226 585
R227 B.n228 B.n227 585
R228 B.n327 B.n326 585
R229 B.n328 B.n327 585
R230 B.n325 B.n233 585
R231 B.n233 B.n232 585
R232 B.n324 B.n323 585
R233 B.n323 B.n322 585
R234 B.n235 B.n234 585
R235 B.n236 B.n235 585
R236 B.n315 B.n314 585
R237 B.n316 B.n315 585
R238 B.n239 B.n238 585
R239 B.n262 B.n261 585
R240 B.n263 B.n259 585
R241 B.n259 B.n240 585
R242 B.n265 B.n264 585
R243 B.n267 B.n258 585
R244 B.n270 B.n269 585
R245 B.n271 B.n257 585
R246 B.n273 B.n272 585
R247 B.n275 B.n256 585
R248 B.n278 B.n277 585
R249 B.n279 B.n252 585
R250 B.n281 B.n280 585
R251 B.n283 B.n251 585
R252 B.n286 B.n285 585
R253 B.n287 B.n250 585
R254 B.n289 B.n288 585
R255 B.n291 B.n249 585
R256 B.n294 B.n293 585
R257 B.n295 B.n246 585
R258 B.n298 B.n297 585
R259 B.n300 B.n245 585
R260 B.n303 B.n302 585
R261 B.n304 B.n244 585
R262 B.n306 B.n305 585
R263 B.n308 B.n243 585
R264 B.n309 B.n242 585
R265 B.n312 B.n311 585
R266 B.n313 B.n241 585
R267 B.n241 B.n240 585
R268 B.n318 B.n317 585
R269 B.n317 B.n316 585
R270 B.n319 B.n237 585
R271 B.n237 B.n236 585
R272 B.n321 B.n320 585
R273 B.n322 B.n321 585
R274 B.n231 B.n230 585
R275 B.n232 B.n231 585
R276 B.n330 B.n329 585
R277 B.n329 B.n328 585
R278 B.n331 B.n229 585
R279 B.n229 B.n228 585
R280 B.n333 B.n332 585
R281 B.n334 B.n333 585
R282 B.n223 B.n222 585
R283 B.n224 B.n223 585
R284 B.n343 B.n342 585
R285 B.n342 B.n341 585
R286 B.n344 B.n221 585
R287 B.n340 B.n221 585
R288 B.n346 B.n345 585
R289 B.n347 B.n346 585
R290 B.n216 B.n215 585
R291 B.n217 B.n216 585
R292 B.n355 B.n354 585
R293 B.n354 B.n353 585
R294 B.n356 B.n214 585
R295 B.n214 B.n213 585
R296 B.n358 B.n357 585
R297 B.n359 B.n358 585
R298 B.n208 B.n207 585
R299 B.n209 B.n208 585
R300 B.n367 B.n366 585
R301 B.n366 B.n365 585
R302 B.n368 B.n206 585
R303 B.n206 B.n205 585
R304 B.n370 B.n369 585
R305 B.n371 B.n370 585
R306 B.n200 B.n199 585
R307 B.n201 B.n200 585
R308 B.n379 B.n378 585
R309 B.n378 B.n377 585
R310 B.n380 B.n198 585
R311 B.n198 B.n197 585
R312 B.n382 B.n381 585
R313 B.n383 B.n382 585
R314 B.n192 B.n191 585
R315 B.n193 B.n192 585
R316 B.n391 B.n390 585
R317 B.n390 B.n389 585
R318 B.n392 B.n190 585
R319 B.n190 B.n189 585
R320 B.n394 B.n393 585
R321 B.n395 B.n394 585
R322 B.n184 B.n183 585
R323 B.n185 B.n184 585
R324 B.n403 B.n402 585
R325 B.n402 B.n401 585
R326 B.n404 B.n182 585
R327 B.n182 B.n181 585
R328 B.n406 B.n405 585
R329 B.n407 B.n406 585
R330 B.n176 B.n175 585
R331 B.n177 B.n176 585
R332 B.n415 B.n414 585
R333 B.n414 B.n413 585
R334 B.n416 B.n174 585
R335 B.n174 B.n173 585
R336 B.n418 B.n417 585
R337 B.n419 B.n418 585
R338 B.n168 B.n167 585
R339 B.n169 B.n168 585
R340 B.n427 B.n426 585
R341 B.n426 B.n425 585
R342 B.n428 B.n166 585
R343 B.n166 B.n165 585
R344 B.n430 B.n429 585
R345 B.n431 B.n430 585
R346 B.n160 B.n159 585
R347 B.n161 B.n160 585
R348 B.n440 B.n439 585
R349 B.n439 B.n438 585
R350 B.n441 B.n158 585
R351 B.n158 B.n157 585
R352 B.n443 B.n442 585
R353 B.n444 B.n443 585
R354 B.n3 B.n0 585
R355 B.n4 B.n3 585
R356 B.n596 B.n1 585
R357 B.n597 B.n596 585
R358 B.n595 B.n594 585
R359 B.n595 B.n8 585
R360 B.n593 B.n9 585
R361 B.n12 B.n9 585
R362 B.n592 B.n591 585
R363 B.n591 B.n590 585
R364 B.n11 B.n10 585
R365 B.n589 B.n11 585
R366 B.n587 B.n586 585
R367 B.n588 B.n587 585
R368 B.n585 B.n17 585
R369 B.n17 B.n16 585
R370 B.n584 B.n583 585
R371 B.n583 B.n582 585
R372 B.n19 B.n18 585
R373 B.n581 B.n19 585
R374 B.n579 B.n578 585
R375 B.n580 B.n579 585
R376 B.n577 B.n24 585
R377 B.n24 B.n23 585
R378 B.n576 B.n575 585
R379 B.n575 B.n574 585
R380 B.n26 B.n25 585
R381 B.n573 B.n26 585
R382 B.n571 B.n570 585
R383 B.n572 B.n571 585
R384 B.n569 B.n31 585
R385 B.n31 B.n30 585
R386 B.n568 B.n567 585
R387 B.n567 B.n566 585
R388 B.n33 B.n32 585
R389 B.n565 B.n33 585
R390 B.n563 B.n562 585
R391 B.n564 B.n563 585
R392 B.n561 B.n38 585
R393 B.n38 B.n37 585
R394 B.n560 B.n559 585
R395 B.n559 B.n558 585
R396 B.n40 B.n39 585
R397 B.n557 B.n40 585
R398 B.n555 B.n554 585
R399 B.n556 B.n555 585
R400 B.n553 B.n45 585
R401 B.n45 B.n44 585
R402 B.n552 B.n551 585
R403 B.n551 B.n550 585
R404 B.n47 B.n46 585
R405 B.n549 B.n47 585
R406 B.n547 B.n546 585
R407 B.n548 B.n547 585
R408 B.n545 B.n52 585
R409 B.n52 B.n51 585
R410 B.n544 B.n543 585
R411 B.n543 B.n542 585
R412 B.n54 B.n53 585
R413 B.n541 B.n54 585
R414 B.n539 B.n538 585
R415 B.n540 B.n539 585
R416 B.n537 B.n59 585
R417 B.n59 B.n58 585
R418 B.n536 B.n535 585
R419 B.n535 B.n534 585
R420 B.n61 B.n60 585
R421 B.n533 B.n61 585
R422 B.n531 B.n530 585
R423 B.n532 B.n531 585
R424 B.n529 B.n65 585
R425 B.n68 B.n65 585
R426 B.n528 B.n527 585
R427 B.n527 B.n526 585
R428 B.n67 B.n66 585
R429 B.n525 B.n67 585
R430 B.n523 B.n522 585
R431 B.n524 B.n523 585
R432 B.n521 B.n73 585
R433 B.n73 B.n72 585
R434 B.n520 B.n519 585
R435 B.n519 B.n518 585
R436 B.n75 B.n74 585
R437 B.n517 B.n75 585
R438 B.n515 B.n514 585
R439 B.n516 B.n515 585
R440 B.n513 B.n80 585
R441 B.n80 B.n79 585
R442 B.n512 B.n511 585
R443 B.n511 B.n510 585
R444 B.n600 B.n599 585
R445 B.n598 B.n2 585
R446 B.n511 B.n82 526.135
R447 B.n507 B.n83 526.135
R448 B.n315 B.n241 526.135
R449 B.n317 B.n239 526.135
R450 B.n100 B.t6 314.188
R451 B.n98 B.t9 314.188
R452 B.n247 B.t14 314.188
R453 B.n253 B.t17 314.188
R454 B.n509 B.n508 256.663
R455 B.n509 B.n96 256.663
R456 B.n509 B.n95 256.663
R457 B.n509 B.n94 256.663
R458 B.n509 B.n93 256.663
R459 B.n509 B.n92 256.663
R460 B.n509 B.n91 256.663
R461 B.n509 B.n90 256.663
R462 B.n509 B.n89 256.663
R463 B.n509 B.n88 256.663
R464 B.n509 B.n87 256.663
R465 B.n509 B.n86 256.663
R466 B.n509 B.n85 256.663
R467 B.n509 B.n84 256.663
R468 B.n260 B.n240 256.663
R469 B.n266 B.n240 256.663
R470 B.n268 B.n240 256.663
R471 B.n274 B.n240 256.663
R472 B.n276 B.n240 256.663
R473 B.n282 B.n240 256.663
R474 B.n284 B.n240 256.663
R475 B.n290 B.n240 256.663
R476 B.n292 B.n240 256.663
R477 B.n299 B.n240 256.663
R478 B.n301 B.n240 256.663
R479 B.n307 B.n240 256.663
R480 B.n310 B.n240 256.663
R481 B.n602 B.n601 256.663
R482 B.n101 B.t7 233.898
R483 B.n99 B.t10 233.898
R484 B.n248 B.t13 233.898
R485 B.n254 B.t16 233.898
R486 B.n316 B.n240 233.52
R487 B.n510 B.n509 233.52
R488 B.n100 B.t4 209.998
R489 B.n98 B.t8 209.998
R490 B.n247 B.t11 209.998
R491 B.n253 B.t15 209.998
R492 B.n104 B.n103 163.367
R493 B.n108 B.n107 163.367
R494 B.n112 B.n111 163.367
R495 B.n116 B.n115 163.367
R496 B.n121 B.n120 163.367
R497 B.n125 B.n124 163.367
R498 B.n129 B.n128 163.367
R499 B.n133 B.n132 163.367
R500 B.n137 B.n136 163.367
R501 B.n142 B.n141 163.367
R502 B.n146 B.n145 163.367
R503 B.n150 B.n149 163.367
R504 B.n152 B.n97 163.367
R505 B.n315 B.n235 163.367
R506 B.n323 B.n235 163.367
R507 B.n323 B.n233 163.367
R508 B.n327 B.n233 163.367
R509 B.n327 B.n227 163.367
R510 B.n335 B.n227 163.367
R511 B.n335 B.n225 163.367
R512 B.n339 B.n225 163.367
R513 B.n339 B.n220 163.367
R514 B.n348 B.n220 163.367
R515 B.n348 B.n218 163.367
R516 B.n352 B.n218 163.367
R517 B.n352 B.n212 163.367
R518 B.n360 B.n212 163.367
R519 B.n360 B.n210 163.367
R520 B.n364 B.n210 163.367
R521 B.n364 B.n204 163.367
R522 B.n372 B.n204 163.367
R523 B.n372 B.n202 163.367
R524 B.n376 B.n202 163.367
R525 B.n376 B.n196 163.367
R526 B.n384 B.n196 163.367
R527 B.n384 B.n194 163.367
R528 B.n388 B.n194 163.367
R529 B.n388 B.n188 163.367
R530 B.n396 B.n188 163.367
R531 B.n396 B.n186 163.367
R532 B.n400 B.n186 163.367
R533 B.n400 B.n180 163.367
R534 B.n408 B.n180 163.367
R535 B.n408 B.n178 163.367
R536 B.n412 B.n178 163.367
R537 B.n412 B.n172 163.367
R538 B.n420 B.n172 163.367
R539 B.n420 B.n170 163.367
R540 B.n424 B.n170 163.367
R541 B.n424 B.n164 163.367
R542 B.n432 B.n164 163.367
R543 B.n432 B.n162 163.367
R544 B.n437 B.n162 163.367
R545 B.n437 B.n156 163.367
R546 B.n445 B.n156 163.367
R547 B.n446 B.n445 163.367
R548 B.n446 B.n5 163.367
R549 B.n6 B.n5 163.367
R550 B.n7 B.n6 163.367
R551 B.n452 B.n7 163.367
R552 B.n453 B.n452 163.367
R553 B.n453 B.n13 163.367
R554 B.n14 B.n13 163.367
R555 B.n15 B.n14 163.367
R556 B.n458 B.n15 163.367
R557 B.n458 B.n20 163.367
R558 B.n21 B.n20 163.367
R559 B.n22 B.n21 163.367
R560 B.n463 B.n22 163.367
R561 B.n463 B.n27 163.367
R562 B.n28 B.n27 163.367
R563 B.n29 B.n28 163.367
R564 B.n468 B.n29 163.367
R565 B.n468 B.n34 163.367
R566 B.n35 B.n34 163.367
R567 B.n36 B.n35 163.367
R568 B.n473 B.n36 163.367
R569 B.n473 B.n41 163.367
R570 B.n42 B.n41 163.367
R571 B.n43 B.n42 163.367
R572 B.n478 B.n43 163.367
R573 B.n478 B.n48 163.367
R574 B.n49 B.n48 163.367
R575 B.n50 B.n49 163.367
R576 B.n483 B.n50 163.367
R577 B.n483 B.n55 163.367
R578 B.n56 B.n55 163.367
R579 B.n57 B.n56 163.367
R580 B.n488 B.n57 163.367
R581 B.n488 B.n62 163.367
R582 B.n63 B.n62 163.367
R583 B.n64 B.n63 163.367
R584 B.n493 B.n64 163.367
R585 B.n493 B.n69 163.367
R586 B.n70 B.n69 163.367
R587 B.n71 B.n70 163.367
R588 B.n498 B.n71 163.367
R589 B.n498 B.n76 163.367
R590 B.n77 B.n76 163.367
R591 B.n78 B.n77 163.367
R592 B.n503 B.n78 163.367
R593 B.n503 B.n83 163.367
R594 B.n261 B.n259 163.367
R595 B.n265 B.n259 163.367
R596 B.n269 B.n267 163.367
R597 B.n273 B.n257 163.367
R598 B.n277 B.n275 163.367
R599 B.n281 B.n252 163.367
R600 B.n285 B.n283 163.367
R601 B.n289 B.n250 163.367
R602 B.n293 B.n291 163.367
R603 B.n298 B.n246 163.367
R604 B.n302 B.n300 163.367
R605 B.n306 B.n244 163.367
R606 B.n309 B.n308 163.367
R607 B.n311 B.n241 163.367
R608 B.n317 B.n237 163.367
R609 B.n321 B.n237 163.367
R610 B.n321 B.n231 163.367
R611 B.n329 B.n231 163.367
R612 B.n329 B.n229 163.367
R613 B.n333 B.n229 163.367
R614 B.n333 B.n223 163.367
R615 B.n342 B.n223 163.367
R616 B.n342 B.n221 163.367
R617 B.n346 B.n221 163.367
R618 B.n346 B.n216 163.367
R619 B.n354 B.n216 163.367
R620 B.n354 B.n214 163.367
R621 B.n358 B.n214 163.367
R622 B.n358 B.n208 163.367
R623 B.n366 B.n208 163.367
R624 B.n366 B.n206 163.367
R625 B.n370 B.n206 163.367
R626 B.n370 B.n200 163.367
R627 B.n378 B.n200 163.367
R628 B.n378 B.n198 163.367
R629 B.n382 B.n198 163.367
R630 B.n382 B.n192 163.367
R631 B.n390 B.n192 163.367
R632 B.n390 B.n190 163.367
R633 B.n394 B.n190 163.367
R634 B.n394 B.n184 163.367
R635 B.n402 B.n184 163.367
R636 B.n402 B.n182 163.367
R637 B.n406 B.n182 163.367
R638 B.n406 B.n176 163.367
R639 B.n414 B.n176 163.367
R640 B.n414 B.n174 163.367
R641 B.n418 B.n174 163.367
R642 B.n418 B.n168 163.367
R643 B.n426 B.n168 163.367
R644 B.n426 B.n166 163.367
R645 B.n430 B.n166 163.367
R646 B.n430 B.n160 163.367
R647 B.n439 B.n160 163.367
R648 B.n439 B.n158 163.367
R649 B.n443 B.n158 163.367
R650 B.n443 B.n3 163.367
R651 B.n600 B.n3 163.367
R652 B.n596 B.n2 163.367
R653 B.n596 B.n595 163.367
R654 B.n595 B.n9 163.367
R655 B.n591 B.n9 163.367
R656 B.n591 B.n11 163.367
R657 B.n587 B.n11 163.367
R658 B.n587 B.n17 163.367
R659 B.n583 B.n17 163.367
R660 B.n583 B.n19 163.367
R661 B.n579 B.n19 163.367
R662 B.n579 B.n24 163.367
R663 B.n575 B.n24 163.367
R664 B.n575 B.n26 163.367
R665 B.n571 B.n26 163.367
R666 B.n571 B.n31 163.367
R667 B.n567 B.n31 163.367
R668 B.n567 B.n33 163.367
R669 B.n563 B.n33 163.367
R670 B.n563 B.n38 163.367
R671 B.n559 B.n38 163.367
R672 B.n559 B.n40 163.367
R673 B.n555 B.n40 163.367
R674 B.n555 B.n45 163.367
R675 B.n551 B.n45 163.367
R676 B.n551 B.n47 163.367
R677 B.n547 B.n47 163.367
R678 B.n547 B.n52 163.367
R679 B.n543 B.n52 163.367
R680 B.n543 B.n54 163.367
R681 B.n539 B.n54 163.367
R682 B.n539 B.n59 163.367
R683 B.n535 B.n59 163.367
R684 B.n535 B.n61 163.367
R685 B.n531 B.n61 163.367
R686 B.n531 B.n65 163.367
R687 B.n527 B.n65 163.367
R688 B.n527 B.n67 163.367
R689 B.n523 B.n67 163.367
R690 B.n523 B.n73 163.367
R691 B.n519 B.n73 163.367
R692 B.n519 B.n75 163.367
R693 B.n515 B.n75 163.367
R694 B.n515 B.n80 163.367
R695 B.n511 B.n80 163.367
R696 B.n316 B.n236 119.394
R697 B.n322 B.n236 119.394
R698 B.n322 B.n232 119.394
R699 B.n328 B.n232 119.394
R700 B.n328 B.n228 119.394
R701 B.n334 B.n228 119.394
R702 B.n334 B.n224 119.394
R703 B.n341 B.n224 119.394
R704 B.n341 B.n340 119.394
R705 B.n347 B.n217 119.394
R706 B.n353 B.n217 119.394
R707 B.n353 B.n213 119.394
R708 B.n359 B.n213 119.394
R709 B.n359 B.n209 119.394
R710 B.n365 B.n209 119.394
R711 B.n365 B.n205 119.394
R712 B.n371 B.n205 119.394
R713 B.n371 B.n201 119.394
R714 B.n377 B.n201 119.394
R715 B.n377 B.n197 119.394
R716 B.n383 B.n197 119.394
R717 B.n383 B.n193 119.394
R718 B.n389 B.n193 119.394
R719 B.n395 B.n189 119.394
R720 B.n395 B.n185 119.394
R721 B.n401 B.n185 119.394
R722 B.n401 B.n181 119.394
R723 B.n407 B.n181 119.394
R724 B.n407 B.n177 119.394
R725 B.n413 B.n177 119.394
R726 B.n413 B.n173 119.394
R727 B.n419 B.n173 119.394
R728 B.n419 B.n169 119.394
R729 B.n425 B.n169 119.394
R730 B.n431 B.n165 119.394
R731 B.n431 B.n161 119.394
R732 B.n438 B.n161 119.394
R733 B.n438 B.n157 119.394
R734 B.n444 B.n157 119.394
R735 B.n444 B.n4 119.394
R736 B.n599 B.n4 119.394
R737 B.n599 B.n598 119.394
R738 B.n598 B.n597 119.394
R739 B.n597 B.n8 119.394
R740 B.n12 B.n8 119.394
R741 B.n590 B.n12 119.394
R742 B.n590 B.n589 119.394
R743 B.n589 B.n588 119.394
R744 B.n588 B.n16 119.394
R745 B.n582 B.n581 119.394
R746 B.n581 B.n580 119.394
R747 B.n580 B.n23 119.394
R748 B.n574 B.n23 119.394
R749 B.n574 B.n573 119.394
R750 B.n573 B.n572 119.394
R751 B.n572 B.n30 119.394
R752 B.n566 B.n30 119.394
R753 B.n566 B.n565 119.394
R754 B.n565 B.n564 119.394
R755 B.n564 B.n37 119.394
R756 B.n558 B.n557 119.394
R757 B.n557 B.n556 119.394
R758 B.n556 B.n44 119.394
R759 B.n550 B.n44 119.394
R760 B.n550 B.n549 119.394
R761 B.n549 B.n548 119.394
R762 B.n548 B.n51 119.394
R763 B.n542 B.n51 119.394
R764 B.n542 B.n541 119.394
R765 B.n541 B.n540 119.394
R766 B.n540 B.n58 119.394
R767 B.n534 B.n58 119.394
R768 B.n534 B.n533 119.394
R769 B.n533 B.n532 119.394
R770 B.n526 B.n68 119.394
R771 B.n526 B.n525 119.394
R772 B.n525 B.n524 119.394
R773 B.n524 B.n72 119.394
R774 B.n518 B.n72 119.394
R775 B.n518 B.n517 119.394
R776 B.n517 B.n516 119.394
R777 B.n516 B.n79 119.394
R778 B.n510 B.n79 119.394
R779 B.n425 B.t3 96.5687
R780 B.n582 B.t1 96.5687
R781 B.n347 B.t12 89.5456
R782 B.n532 B.t5 89.5456
R783 B.n101 B.n100 80.2914
R784 B.n99 B.n98 80.2914
R785 B.n248 B.n247 80.2914
R786 B.n254 B.n253 80.2914
R787 B.n389 B.t2 75.4993
R788 B.n558 B.t0 75.4993
R789 B.n84 B.n82 71.676
R790 B.n104 B.n85 71.676
R791 B.n108 B.n86 71.676
R792 B.n112 B.n87 71.676
R793 B.n116 B.n88 71.676
R794 B.n121 B.n89 71.676
R795 B.n125 B.n90 71.676
R796 B.n129 B.n91 71.676
R797 B.n133 B.n92 71.676
R798 B.n137 B.n93 71.676
R799 B.n142 B.n94 71.676
R800 B.n146 B.n95 71.676
R801 B.n150 B.n96 71.676
R802 B.n508 B.n97 71.676
R803 B.n508 B.n507 71.676
R804 B.n152 B.n96 71.676
R805 B.n149 B.n95 71.676
R806 B.n145 B.n94 71.676
R807 B.n141 B.n93 71.676
R808 B.n136 B.n92 71.676
R809 B.n132 B.n91 71.676
R810 B.n128 B.n90 71.676
R811 B.n124 B.n89 71.676
R812 B.n120 B.n88 71.676
R813 B.n115 B.n87 71.676
R814 B.n111 B.n86 71.676
R815 B.n107 B.n85 71.676
R816 B.n103 B.n84 71.676
R817 B.n260 B.n239 71.676
R818 B.n266 B.n265 71.676
R819 B.n269 B.n268 71.676
R820 B.n274 B.n273 71.676
R821 B.n277 B.n276 71.676
R822 B.n282 B.n281 71.676
R823 B.n285 B.n284 71.676
R824 B.n290 B.n289 71.676
R825 B.n293 B.n292 71.676
R826 B.n299 B.n298 71.676
R827 B.n302 B.n301 71.676
R828 B.n307 B.n306 71.676
R829 B.n310 B.n309 71.676
R830 B.n261 B.n260 71.676
R831 B.n267 B.n266 71.676
R832 B.n268 B.n257 71.676
R833 B.n275 B.n274 71.676
R834 B.n276 B.n252 71.676
R835 B.n283 B.n282 71.676
R836 B.n284 B.n250 71.676
R837 B.n291 B.n290 71.676
R838 B.n292 B.n246 71.676
R839 B.n300 B.n299 71.676
R840 B.n301 B.n244 71.676
R841 B.n308 B.n307 71.676
R842 B.n311 B.n310 71.676
R843 B.n601 B.n600 71.676
R844 B.n601 B.n2 71.676
R845 B.n118 B.n101 59.5399
R846 B.n139 B.n99 59.5399
R847 B.n296 B.n248 59.5399
R848 B.n255 B.n254 59.5399
R849 B.t2 B.n189 43.8952
R850 B.t0 B.n37 43.8952
R851 B.n318 B.n238 34.1859
R852 B.n314 B.n313 34.1859
R853 B.n506 B.n505 34.1859
R854 B.n512 B.n81 34.1859
R855 B.n340 B.t12 29.8489
R856 B.n68 B.t5 29.8489
R857 B.t3 B.n165 22.8257
R858 B.t1 B.n16 22.8257
R859 B B.n602 18.0485
R860 B.n319 B.n318 10.6151
R861 B.n320 B.n319 10.6151
R862 B.n320 B.n230 10.6151
R863 B.n330 B.n230 10.6151
R864 B.n331 B.n330 10.6151
R865 B.n332 B.n331 10.6151
R866 B.n332 B.n222 10.6151
R867 B.n343 B.n222 10.6151
R868 B.n344 B.n343 10.6151
R869 B.n345 B.n344 10.6151
R870 B.n345 B.n215 10.6151
R871 B.n355 B.n215 10.6151
R872 B.n356 B.n355 10.6151
R873 B.n357 B.n356 10.6151
R874 B.n357 B.n207 10.6151
R875 B.n367 B.n207 10.6151
R876 B.n368 B.n367 10.6151
R877 B.n369 B.n368 10.6151
R878 B.n369 B.n199 10.6151
R879 B.n379 B.n199 10.6151
R880 B.n380 B.n379 10.6151
R881 B.n381 B.n380 10.6151
R882 B.n381 B.n191 10.6151
R883 B.n391 B.n191 10.6151
R884 B.n392 B.n391 10.6151
R885 B.n393 B.n392 10.6151
R886 B.n393 B.n183 10.6151
R887 B.n403 B.n183 10.6151
R888 B.n404 B.n403 10.6151
R889 B.n405 B.n404 10.6151
R890 B.n405 B.n175 10.6151
R891 B.n415 B.n175 10.6151
R892 B.n416 B.n415 10.6151
R893 B.n417 B.n416 10.6151
R894 B.n417 B.n167 10.6151
R895 B.n427 B.n167 10.6151
R896 B.n428 B.n427 10.6151
R897 B.n429 B.n428 10.6151
R898 B.n429 B.n159 10.6151
R899 B.n440 B.n159 10.6151
R900 B.n441 B.n440 10.6151
R901 B.n442 B.n441 10.6151
R902 B.n442 B.n0 10.6151
R903 B.n262 B.n238 10.6151
R904 B.n263 B.n262 10.6151
R905 B.n264 B.n263 10.6151
R906 B.n264 B.n258 10.6151
R907 B.n270 B.n258 10.6151
R908 B.n271 B.n270 10.6151
R909 B.n272 B.n271 10.6151
R910 B.n272 B.n256 10.6151
R911 B.n279 B.n278 10.6151
R912 B.n280 B.n279 10.6151
R913 B.n280 B.n251 10.6151
R914 B.n286 B.n251 10.6151
R915 B.n287 B.n286 10.6151
R916 B.n288 B.n287 10.6151
R917 B.n288 B.n249 10.6151
R918 B.n294 B.n249 10.6151
R919 B.n295 B.n294 10.6151
R920 B.n297 B.n245 10.6151
R921 B.n303 B.n245 10.6151
R922 B.n304 B.n303 10.6151
R923 B.n305 B.n304 10.6151
R924 B.n305 B.n243 10.6151
R925 B.n243 B.n242 10.6151
R926 B.n312 B.n242 10.6151
R927 B.n313 B.n312 10.6151
R928 B.n314 B.n234 10.6151
R929 B.n324 B.n234 10.6151
R930 B.n325 B.n324 10.6151
R931 B.n326 B.n325 10.6151
R932 B.n326 B.n226 10.6151
R933 B.n336 B.n226 10.6151
R934 B.n337 B.n336 10.6151
R935 B.n338 B.n337 10.6151
R936 B.n338 B.n219 10.6151
R937 B.n349 B.n219 10.6151
R938 B.n350 B.n349 10.6151
R939 B.n351 B.n350 10.6151
R940 B.n351 B.n211 10.6151
R941 B.n361 B.n211 10.6151
R942 B.n362 B.n361 10.6151
R943 B.n363 B.n362 10.6151
R944 B.n363 B.n203 10.6151
R945 B.n373 B.n203 10.6151
R946 B.n374 B.n373 10.6151
R947 B.n375 B.n374 10.6151
R948 B.n375 B.n195 10.6151
R949 B.n385 B.n195 10.6151
R950 B.n386 B.n385 10.6151
R951 B.n387 B.n386 10.6151
R952 B.n387 B.n187 10.6151
R953 B.n397 B.n187 10.6151
R954 B.n398 B.n397 10.6151
R955 B.n399 B.n398 10.6151
R956 B.n399 B.n179 10.6151
R957 B.n409 B.n179 10.6151
R958 B.n410 B.n409 10.6151
R959 B.n411 B.n410 10.6151
R960 B.n411 B.n171 10.6151
R961 B.n421 B.n171 10.6151
R962 B.n422 B.n421 10.6151
R963 B.n423 B.n422 10.6151
R964 B.n423 B.n163 10.6151
R965 B.n433 B.n163 10.6151
R966 B.n434 B.n433 10.6151
R967 B.n436 B.n434 10.6151
R968 B.n436 B.n435 10.6151
R969 B.n435 B.n155 10.6151
R970 B.n447 B.n155 10.6151
R971 B.n448 B.n447 10.6151
R972 B.n449 B.n448 10.6151
R973 B.n450 B.n449 10.6151
R974 B.n451 B.n450 10.6151
R975 B.n454 B.n451 10.6151
R976 B.n455 B.n454 10.6151
R977 B.n456 B.n455 10.6151
R978 B.n457 B.n456 10.6151
R979 B.n459 B.n457 10.6151
R980 B.n460 B.n459 10.6151
R981 B.n461 B.n460 10.6151
R982 B.n462 B.n461 10.6151
R983 B.n464 B.n462 10.6151
R984 B.n465 B.n464 10.6151
R985 B.n466 B.n465 10.6151
R986 B.n467 B.n466 10.6151
R987 B.n469 B.n467 10.6151
R988 B.n470 B.n469 10.6151
R989 B.n471 B.n470 10.6151
R990 B.n472 B.n471 10.6151
R991 B.n474 B.n472 10.6151
R992 B.n475 B.n474 10.6151
R993 B.n476 B.n475 10.6151
R994 B.n477 B.n476 10.6151
R995 B.n479 B.n477 10.6151
R996 B.n480 B.n479 10.6151
R997 B.n481 B.n480 10.6151
R998 B.n482 B.n481 10.6151
R999 B.n484 B.n482 10.6151
R1000 B.n485 B.n484 10.6151
R1001 B.n486 B.n485 10.6151
R1002 B.n487 B.n486 10.6151
R1003 B.n489 B.n487 10.6151
R1004 B.n490 B.n489 10.6151
R1005 B.n491 B.n490 10.6151
R1006 B.n492 B.n491 10.6151
R1007 B.n494 B.n492 10.6151
R1008 B.n495 B.n494 10.6151
R1009 B.n496 B.n495 10.6151
R1010 B.n497 B.n496 10.6151
R1011 B.n499 B.n497 10.6151
R1012 B.n500 B.n499 10.6151
R1013 B.n501 B.n500 10.6151
R1014 B.n502 B.n501 10.6151
R1015 B.n504 B.n502 10.6151
R1016 B.n505 B.n504 10.6151
R1017 B.n594 B.n1 10.6151
R1018 B.n594 B.n593 10.6151
R1019 B.n593 B.n592 10.6151
R1020 B.n592 B.n10 10.6151
R1021 B.n586 B.n10 10.6151
R1022 B.n586 B.n585 10.6151
R1023 B.n585 B.n584 10.6151
R1024 B.n584 B.n18 10.6151
R1025 B.n578 B.n18 10.6151
R1026 B.n578 B.n577 10.6151
R1027 B.n577 B.n576 10.6151
R1028 B.n576 B.n25 10.6151
R1029 B.n570 B.n25 10.6151
R1030 B.n570 B.n569 10.6151
R1031 B.n569 B.n568 10.6151
R1032 B.n568 B.n32 10.6151
R1033 B.n562 B.n32 10.6151
R1034 B.n562 B.n561 10.6151
R1035 B.n561 B.n560 10.6151
R1036 B.n560 B.n39 10.6151
R1037 B.n554 B.n39 10.6151
R1038 B.n554 B.n553 10.6151
R1039 B.n553 B.n552 10.6151
R1040 B.n552 B.n46 10.6151
R1041 B.n546 B.n46 10.6151
R1042 B.n546 B.n545 10.6151
R1043 B.n545 B.n544 10.6151
R1044 B.n544 B.n53 10.6151
R1045 B.n538 B.n53 10.6151
R1046 B.n538 B.n537 10.6151
R1047 B.n537 B.n536 10.6151
R1048 B.n536 B.n60 10.6151
R1049 B.n530 B.n60 10.6151
R1050 B.n530 B.n529 10.6151
R1051 B.n529 B.n528 10.6151
R1052 B.n528 B.n66 10.6151
R1053 B.n522 B.n66 10.6151
R1054 B.n522 B.n521 10.6151
R1055 B.n521 B.n520 10.6151
R1056 B.n520 B.n74 10.6151
R1057 B.n514 B.n74 10.6151
R1058 B.n514 B.n513 10.6151
R1059 B.n513 B.n512 10.6151
R1060 B.n102 B.n81 10.6151
R1061 B.n105 B.n102 10.6151
R1062 B.n106 B.n105 10.6151
R1063 B.n109 B.n106 10.6151
R1064 B.n110 B.n109 10.6151
R1065 B.n113 B.n110 10.6151
R1066 B.n114 B.n113 10.6151
R1067 B.n117 B.n114 10.6151
R1068 B.n122 B.n119 10.6151
R1069 B.n123 B.n122 10.6151
R1070 B.n126 B.n123 10.6151
R1071 B.n127 B.n126 10.6151
R1072 B.n130 B.n127 10.6151
R1073 B.n131 B.n130 10.6151
R1074 B.n134 B.n131 10.6151
R1075 B.n135 B.n134 10.6151
R1076 B.n138 B.n135 10.6151
R1077 B.n143 B.n140 10.6151
R1078 B.n144 B.n143 10.6151
R1079 B.n147 B.n144 10.6151
R1080 B.n148 B.n147 10.6151
R1081 B.n151 B.n148 10.6151
R1082 B.n153 B.n151 10.6151
R1083 B.n154 B.n153 10.6151
R1084 B.n506 B.n154 10.6151
R1085 B.n256 B.n255 9.36635
R1086 B.n297 B.n296 9.36635
R1087 B.n118 B.n117 9.36635
R1088 B.n140 B.n139 9.36635
R1089 B.n602 B.n0 8.11757
R1090 B.n602 B.n1 8.11757
R1091 B.n278 B.n255 1.24928
R1092 B.n296 B.n295 1.24928
R1093 B.n119 B.n118 1.24928
R1094 B.n139 B.n138 1.24928
R1095 VP.n21 VP.n20 161.3
R1096 VP.n19 VP.n1 161.3
R1097 VP.n18 VP.n17 161.3
R1098 VP.n16 VP.n2 161.3
R1099 VP.n15 VP.n14 161.3
R1100 VP.n13 VP.n3 161.3
R1101 VP.n12 VP.n11 161.3
R1102 VP.n10 VP.n4 161.3
R1103 VP.n9 VP.n8 161.3
R1104 VP.n7 VP.n6 86.642
R1105 VP.n22 VP.n0 86.642
R1106 VP.n6 VP.n5 43.5898
R1107 VP.n14 VP.n13 40.4934
R1108 VP.n14 VP.n2 40.4934
R1109 VP.n5 VP.t0 40.2662
R1110 VP.n5 VP.t3 38.9138
R1111 VP.n8 VP.n4 24.4675
R1112 VP.n12 VP.n4 24.4675
R1113 VP.n13 VP.n12 24.4675
R1114 VP.n18 VP.n2 24.4675
R1115 VP.n19 VP.n18 24.4675
R1116 VP.n20 VP.n19 24.4675
R1117 VP.n7 VP.t1 6.2627
R1118 VP.n0 VP.t2 6.2627
R1119 VP.n8 VP.n7 3.42588
R1120 VP.n20 VP.n0 3.42588
R1121 VP.n9 VP.n6 0.354971
R1122 VP.n22 VP.n21 0.354971
R1123 VP VP.n22 0.26696
R1124 VP.n10 VP.n9 0.189894
R1125 VP.n11 VP.n10 0.189894
R1126 VP.n11 VP.n3 0.189894
R1127 VP.n15 VP.n3 0.189894
R1128 VP.n16 VP.n15 0.189894
R1129 VP.n17 VP.n16 0.189894
R1130 VP.n17 VP.n1 0.189894
R1131 VP.n21 VP.n1 0.189894
R1132 VDD1 VDD1.n1 275.738
R1133 VDD1 VDD1.n0 239.998
R1134 VDD1.n0 VDD1.t3 20.0005
R1135 VDD1.n0 VDD1.t0 20.0005
R1136 VDD1.n1 VDD1.t2 20.0005
R1137 VDD1.n1 VDD1.t1 20.0005
C0 VTAIL VDD2 3.52362f
C1 VDD1 VDD2 1.32077f
C2 VDD1 VTAIL 3.4613f
C3 VDD2 VP 0.47981f
C4 VTAIL VP 1.75264f
C5 VDD2 VN 0.735278f
C6 VDD1 VP 1.05514f
C7 VTAIL VN 1.73854f
C8 VDD1 VN 0.156975f
C9 VP VN 5.03327f
C10 VDD2 B 3.563102f
C11 VDD1 B 6.7419f
C12 VTAIL B 3.424185f
C13 VN B 11.94529f
C14 VP B 10.445541f
C15 VDD1.t3 B 0.019634f
C16 VDD1.t0 B 0.019634f
C17 VDD1.n0 B 0.076394f
C18 VDD1.t2 B 0.019634f
C19 VDD1.t1 B 0.019634f
C20 VDD1.n1 B 0.203559f
C21 VP.t2 B 0.166675f
C22 VP.n0 B 0.195769f
C23 VP.n1 B 0.023772f
C24 VP.n2 B 0.047246f
C25 VP.n3 B 0.023772f
C26 VP.n4 B 0.044304f
C27 VP.t0 B 0.42218f
C28 VP.t3 B 0.409873f
C29 VP.n5 B 1.60934f
C30 VP.n6 B 1.12595f
C31 VP.t1 B 0.166675f
C32 VP.n7 B 0.195769f
C33 VP.n8 B 0.025493f
C34 VP.n9 B 0.038367f
C35 VP.n10 B 0.023772f
C36 VP.n11 B 0.023772f
C37 VP.n12 B 0.044304f
C38 VP.n13 B 0.047246f
C39 VP.n14 B 0.019217f
C40 VP.n15 B 0.023772f
C41 VP.n16 B 0.023772f
C42 VP.n17 B 0.023772f
C43 VP.n18 B 0.044304f
C44 VP.n19 B 0.044304f
C45 VP.n20 B 0.025493f
C46 VP.n21 B 0.038367f
C47 VP.n22 B 0.072774f
C48 VTAIL.t4 B 0.103012f
C49 VTAIL.n0 B 0.328469f
C50 VTAIL.t3 B 0.103012f
C51 VTAIL.n1 B 0.46024f
C52 VTAIL.t2 B 0.103012f
C53 VTAIL.n2 B 1.08374f
C54 VTAIL.t7 B 0.103012f
C55 VTAIL.n3 B 1.08374f
C56 VTAIL.t5 B 0.103012f
C57 VTAIL.n4 B 0.46024f
C58 VTAIL.t1 B 0.103012f
C59 VTAIL.n5 B 0.46024f
C60 VTAIL.t0 B 0.103012f
C61 VTAIL.n6 B 1.08374f
C62 VTAIL.t6 B 0.103012f
C63 VTAIL.n7 B 0.943081f
C64 VDD2.t1 B 0.020169f
C65 VDD2.t0 B 0.020169f
C66 VDD2.n0 B 0.200796f
C67 VDD2.t3 B 0.020169f
C68 VDD2.t2 B 0.020169f
C69 VDD2.n1 B 0.078353f
C70 VDD2.n2 B 2.83816f
C71 VN.t1 B 0.407152f
C72 VN.t3 B 0.419378f
C73 VN.n0 B 0.371798f
C74 VN.t0 B 0.407152f
C75 VN.t2 B 0.419378f
C76 VN.n1 B 1.60875f
.ends

