* NGSPICE file created from diff_pair_sample_1696.ext - technology: sky130A

.subckt diff_pair_sample_1696 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=1.6926 pd=9.46 as=0 ps=0 w=4.34 l=2.86
X1 VTAIL.t11 VP.t0 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6926 pd=9.46 as=0.7161 ps=4.67 w=4.34 l=2.86
X2 VTAIL.t15 VN.t0 VDD2.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6926 pd=9.46 as=0.7161 ps=4.67 w=4.34 l=2.86
X3 VDD1.t6 VP.t1 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=0.7161 pd=4.67 as=0.7161 ps=4.67 w=4.34 l=2.86
X4 VDD2.t6 VN.t1 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7161 pd=4.67 as=1.6926 ps=9.46 w=4.34 l=2.86
X5 VDD1.t5 VP.t2 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7161 pd=4.67 as=1.6926 ps=9.46 w=4.34 l=2.86
X6 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=1.6926 pd=9.46 as=0 ps=0 w=4.34 l=2.86
X7 VTAIL.t8 VP.t3 VDD1.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=0.7161 pd=4.67 as=0.7161 ps=4.67 w=4.34 l=2.86
X8 VTAIL.t0 VN.t2 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=0.7161 pd=4.67 as=0.7161 ps=4.67 w=4.34 l=2.86
X9 VTAIL.t3 VN.t3 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6926 pd=9.46 as=0.7161 ps=4.67 w=4.34 l=2.86
X10 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=1.6926 pd=9.46 as=0 ps=0 w=4.34 l=2.86
X11 VDD1.t7 VP.t4 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7161 pd=4.67 as=0.7161 ps=4.67 w=4.34 l=2.86
X12 VDD2.t3 VN.t4 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7161 pd=4.67 as=0.7161 ps=4.67 w=4.34 l=2.86
X13 VDD2.t2 VN.t5 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=0.7161 pd=4.67 as=1.6926 ps=9.46 w=4.34 l=2.86
X14 VDD2.t1 VN.t6 VTAIL.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=0.7161 pd=4.67 as=0.7161 ps=4.67 w=4.34 l=2.86
X15 VDD1.t2 VP.t5 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.7161 pd=4.67 as=1.6926 ps=9.46 w=4.34 l=2.86
X16 VTAIL.t5 VP.t6 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=0.7161 pd=4.67 as=0.7161 ps=4.67 w=4.34 l=2.86
X17 VTAIL.t4 VP.t7 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6926 pd=9.46 as=0.7161 ps=4.67 w=4.34 l=2.86
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.6926 pd=9.46 as=0 ps=0 w=4.34 l=2.86
X19 VTAIL.t1 VN.t7 VDD2.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=0.7161 pd=4.67 as=0.7161 ps=4.67 w=4.34 l=2.86
R0 B.n690 B.n689 585
R1 B.n221 B.n125 585
R2 B.n220 B.n219 585
R3 B.n218 B.n217 585
R4 B.n216 B.n215 585
R5 B.n214 B.n213 585
R6 B.n212 B.n211 585
R7 B.n210 B.n209 585
R8 B.n208 B.n207 585
R9 B.n206 B.n205 585
R10 B.n204 B.n203 585
R11 B.n202 B.n201 585
R12 B.n200 B.n199 585
R13 B.n198 B.n197 585
R14 B.n196 B.n195 585
R15 B.n194 B.n193 585
R16 B.n192 B.n191 585
R17 B.n190 B.n189 585
R18 B.n188 B.n187 585
R19 B.n185 B.n184 585
R20 B.n183 B.n182 585
R21 B.n181 B.n180 585
R22 B.n179 B.n178 585
R23 B.n177 B.n176 585
R24 B.n175 B.n174 585
R25 B.n173 B.n172 585
R26 B.n171 B.n170 585
R27 B.n169 B.n168 585
R28 B.n167 B.n166 585
R29 B.n164 B.n163 585
R30 B.n162 B.n161 585
R31 B.n160 B.n159 585
R32 B.n158 B.n157 585
R33 B.n156 B.n155 585
R34 B.n154 B.n153 585
R35 B.n152 B.n151 585
R36 B.n150 B.n149 585
R37 B.n148 B.n147 585
R38 B.n146 B.n145 585
R39 B.n144 B.n143 585
R40 B.n142 B.n141 585
R41 B.n140 B.n139 585
R42 B.n138 B.n137 585
R43 B.n136 B.n135 585
R44 B.n134 B.n133 585
R45 B.n132 B.n131 585
R46 B.n102 B.n101 585
R47 B.n695 B.n694 585
R48 B.n688 B.n126 585
R49 B.n126 B.n99 585
R50 B.n687 B.n98 585
R51 B.n699 B.n98 585
R52 B.n686 B.n97 585
R53 B.n700 B.n97 585
R54 B.n685 B.n96 585
R55 B.n701 B.n96 585
R56 B.n684 B.n683 585
R57 B.n683 B.n92 585
R58 B.n682 B.n91 585
R59 B.n707 B.n91 585
R60 B.n681 B.n90 585
R61 B.n708 B.n90 585
R62 B.n680 B.n89 585
R63 B.n709 B.n89 585
R64 B.n679 B.n678 585
R65 B.n678 B.n85 585
R66 B.n677 B.n84 585
R67 B.n715 B.n84 585
R68 B.n676 B.n83 585
R69 B.n716 B.n83 585
R70 B.n675 B.n82 585
R71 B.n717 B.n82 585
R72 B.n674 B.n673 585
R73 B.n673 B.n78 585
R74 B.n672 B.n77 585
R75 B.n723 B.n77 585
R76 B.n671 B.n76 585
R77 B.n724 B.n76 585
R78 B.n670 B.n75 585
R79 B.n725 B.n75 585
R80 B.n669 B.n668 585
R81 B.n668 B.n71 585
R82 B.n667 B.n70 585
R83 B.n731 B.n70 585
R84 B.n666 B.n69 585
R85 B.n732 B.n69 585
R86 B.n665 B.n68 585
R87 B.n733 B.n68 585
R88 B.n664 B.n663 585
R89 B.n663 B.n67 585
R90 B.n662 B.n63 585
R91 B.n739 B.n63 585
R92 B.n661 B.n62 585
R93 B.n740 B.n62 585
R94 B.n660 B.n61 585
R95 B.n741 B.n61 585
R96 B.n659 B.n658 585
R97 B.n658 B.n57 585
R98 B.n657 B.n56 585
R99 B.n747 B.n56 585
R100 B.n656 B.n55 585
R101 B.n748 B.n55 585
R102 B.n655 B.n54 585
R103 B.n749 B.n54 585
R104 B.n654 B.n653 585
R105 B.n653 B.n50 585
R106 B.n652 B.n49 585
R107 B.n755 B.n49 585
R108 B.n651 B.n48 585
R109 B.n756 B.n48 585
R110 B.n650 B.n47 585
R111 B.n757 B.n47 585
R112 B.n649 B.n648 585
R113 B.n648 B.n43 585
R114 B.n647 B.n42 585
R115 B.n763 B.n42 585
R116 B.n646 B.n41 585
R117 B.n764 B.n41 585
R118 B.n645 B.n40 585
R119 B.n765 B.n40 585
R120 B.n644 B.n643 585
R121 B.n643 B.n36 585
R122 B.n642 B.n35 585
R123 B.n771 B.n35 585
R124 B.n641 B.n34 585
R125 B.n772 B.n34 585
R126 B.n640 B.n33 585
R127 B.n773 B.n33 585
R128 B.n639 B.n638 585
R129 B.n638 B.n29 585
R130 B.n637 B.n28 585
R131 B.n779 B.n28 585
R132 B.n636 B.n27 585
R133 B.n780 B.n27 585
R134 B.n635 B.n26 585
R135 B.n781 B.n26 585
R136 B.n634 B.n633 585
R137 B.n633 B.n22 585
R138 B.n632 B.n21 585
R139 B.n787 B.n21 585
R140 B.n631 B.n20 585
R141 B.n788 B.n20 585
R142 B.n630 B.n19 585
R143 B.n789 B.n19 585
R144 B.n629 B.n628 585
R145 B.n628 B.n18 585
R146 B.n627 B.n14 585
R147 B.n795 B.n14 585
R148 B.n626 B.n13 585
R149 B.n796 B.n13 585
R150 B.n625 B.n12 585
R151 B.n797 B.n12 585
R152 B.n624 B.n623 585
R153 B.n623 B.n8 585
R154 B.n622 B.n7 585
R155 B.n803 B.n7 585
R156 B.n621 B.n6 585
R157 B.n804 B.n6 585
R158 B.n620 B.n5 585
R159 B.n805 B.n5 585
R160 B.n619 B.n618 585
R161 B.n618 B.n4 585
R162 B.n617 B.n222 585
R163 B.n617 B.n616 585
R164 B.n607 B.n223 585
R165 B.n224 B.n223 585
R166 B.n609 B.n608 585
R167 B.n610 B.n609 585
R168 B.n606 B.n229 585
R169 B.n229 B.n228 585
R170 B.n605 B.n604 585
R171 B.n604 B.n603 585
R172 B.n231 B.n230 585
R173 B.n596 B.n231 585
R174 B.n595 B.n594 585
R175 B.n597 B.n595 585
R176 B.n593 B.n236 585
R177 B.n236 B.n235 585
R178 B.n592 B.n591 585
R179 B.n591 B.n590 585
R180 B.n238 B.n237 585
R181 B.n239 B.n238 585
R182 B.n583 B.n582 585
R183 B.n584 B.n583 585
R184 B.n581 B.n244 585
R185 B.n244 B.n243 585
R186 B.n580 B.n579 585
R187 B.n579 B.n578 585
R188 B.n246 B.n245 585
R189 B.n247 B.n246 585
R190 B.n571 B.n570 585
R191 B.n572 B.n571 585
R192 B.n569 B.n252 585
R193 B.n252 B.n251 585
R194 B.n568 B.n567 585
R195 B.n567 B.n566 585
R196 B.n254 B.n253 585
R197 B.n255 B.n254 585
R198 B.n559 B.n558 585
R199 B.n560 B.n559 585
R200 B.n557 B.n260 585
R201 B.n260 B.n259 585
R202 B.n556 B.n555 585
R203 B.n555 B.n554 585
R204 B.n262 B.n261 585
R205 B.n263 B.n262 585
R206 B.n547 B.n546 585
R207 B.n548 B.n547 585
R208 B.n545 B.n268 585
R209 B.n268 B.n267 585
R210 B.n544 B.n543 585
R211 B.n543 B.n542 585
R212 B.n270 B.n269 585
R213 B.n271 B.n270 585
R214 B.n535 B.n534 585
R215 B.n536 B.n535 585
R216 B.n533 B.n276 585
R217 B.n276 B.n275 585
R218 B.n532 B.n531 585
R219 B.n531 B.n530 585
R220 B.n278 B.n277 585
R221 B.n279 B.n278 585
R222 B.n523 B.n522 585
R223 B.n524 B.n523 585
R224 B.n521 B.n284 585
R225 B.n284 B.n283 585
R226 B.n520 B.n519 585
R227 B.n519 B.n518 585
R228 B.n286 B.n285 585
R229 B.n511 B.n286 585
R230 B.n510 B.n509 585
R231 B.n512 B.n510 585
R232 B.n508 B.n291 585
R233 B.n291 B.n290 585
R234 B.n507 B.n506 585
R235 B.n506 B.n505 585
R236 B.n293 B.n292 585
R237 B.n294 B.n293 585
R238 B.n498 B.n497 585
R239 B.n499 B.n498 585
R240 B.n496 B.n299 585
R241 B.n299 B.n298 585
R242 B.n495 B.n494 585
R243 B.n494 B.n493 585
R244 B.n301 B.n300 585
R245 B.n302 B.n301 585
R246 B.n486 B.n485 585
R247 B.n487 B.n486 585
R248 B.n484 B.n307 585
R249 B.n307 B.n306 585
R250 B.n483 B.n482 585
R251 B.n482 B.n481 585
R252 B.n309 B.n308 585
R253 B.n310 B.n309 585
R254 B.n474 B.n473 585
R255 B.n475 B.n474 585
R256 B.n472 B.n315 585
R257 B.n315 B.n314 585
R258 B.n471 B.n470 585
R259 B.n470 B.n469 585
R260 B.n317 B.n316 585
R261 B.n318 B.n317 585
R262 B.n462 B.n461 585
R263 B.n463 B.n462 585
R264 B.n460 B.n323 585
R265 B.n323 B.n322 585
R266 B.n459 B.n458 585
R267 B.n458 B.n457 585
R268 B.n325 B.n324 585
R269 B.n326 B.n325 585
R270 B.n453 B.n452 585
R271 B.n329 B.n328 585
R272 B.n449 B.n448 585
R273 B.n450 B.n449 585
R274 B.n447 B.n353 585
R275 B.n446 B.n445 585
R276 B.n444 B.n443 585
R277 B.n442 B.n441 585
R278 B.n440 B.n439 585
R279 B.n438 B.n437 585
R280 B.n436 B.n435 585
R281 B.n434 B.n433 585
R282 B.n432 B.n431 585
R283 B.n430 B.n429 585
R284 B.n428 B.n427 585
R285 B.n426 B.n425 585
R286 B.n424 B.n423 585
R287 B.n422 B.n421 585
R288 B.n420 B.n419 585
R289 B.n418 B.n417 585
R290 B.n416 B.n415 585
R291 B.n414 B.n413 585
R292 B.n412 B.n411 585
R293 B.n410 B.n409 585
R294 B.n408 B.n407 585
R295 B.n406 B.n405 585
R296 B.n404 B.n403 585
R297 B.n402 B.n401 585
R298 B.n400 B.n399 585
R299 B.n398 B.n397 585
R300 B.n396 B.n395 585
R301 B.n394 B.n393 585
R302 B.n392 B.n391 585
R303 B.n390 B.n389 585
R304 B.n388 B.n387 585
R305 B.n386 B.n385 585
R306 B.n384 B.n383 585
R307 B.n382 B.n381 585
R308 B.n380 B.n379 585
R309 B.n378 B.n377 585
R310 B.n376 B.n375 585
R311 B.n374 B.n373 585
R312 B.n372 B.n371 585
R313 B.n370 B.n369 585
R314 B.n368 B.n367 585
R315 B.n366 B.n365 585
R316 B.n364 B.n363 585
R317 B.n362 B.n361 585
R318 B.n360 B.n352 585
R319 B.n450 B.n352 585
R320 B.n454 B.n327 585
R321 B.n327 B.n326 585
R322 B.n456 B.n455 585
R323 B.n457 B.n456 585
R324 B.n321 B.n320 585
R325 B.n322 B.n321 585
R326 B.n465 B.n464 585
R327 B.n464 B.n463 585
R328 B.n466 B.n319 585
R329 B.n319 B.n318 585
R330 B.n468 B.n467 585
R331 B.n469 B.n468 585
R332 B.n313 B.n312 585
R333 B.n314 B.n313 585
R334 B.n477 B.n476 585
R335 B.n476 B.n475 585
R336 B.n478 B.n311 585
R337 B.n311 B.n310 585
R338 B.n480 B.n479 585
R339 B.n481 B.n480 585
R340 B.n305 B.n304 585
R341 B.n306 B.n305 585
R342 B.n489 B.n488 585
R343 B.n488 B.n487 585
R344 B.n490 B.n303 585
R345 B.n303 B.n302 585
R346 B.n492 B.n491 585
R347 B.n493 B.n492 585
R348 B.n297 B.n296 585
R349 B.n298 B.n297 585
R350 B.n501 B.n500 585
R351 B.n500 B.n499 585
R352 B.n502 B.n295 585
R353 B.n295 B.n294 585
R354 B.n504 B.n503 585
R355 B.n505 B.n504 585
R356 B.n289 B.n288 585
R357 B.n290 B.n289 585
R358 B.n514 B.n513 585
R359 B.n513 B.n512 585
R360 B.n515 B.n287 585
R361 B.n511 B.n287 585
R362 B.n517 B.n516 585
R363 B.n518 B.n517 585
R364 B.n282 B.n281 585
R365 B.n283 B.n282 585
R366 B.n526 B.n525 585
R367 B.n525 B.n524 585
R368 B.n527 B.n280 585
R369 B.n280 B.n279 585
R370 B.n529 B.n528 585
R371 B.n530 B.n529 585
R372 B.n274 B.n273 585
R373 B.n275 B.n274 585
R374 B.n538 B.n537 585
R375 B.n537 B.n536 585
R376 B.n539 B.n272 585
R377 B.n272 B.n271 585
R378 B.n541 B.n540 585
R379 B.n542 B.n541 585
R380 B.n266 B.n265 585
R381 B.n267 B.n266 585
R382 B.n550 B.n549 585
R383 B.n549 B.n548 585
R384 B.n551 B.n264 585
R385 B.n264 B.n263 585
R386 B.n553 B.n552 585
R387 B.n554 B.n553 585
R388 B.n258 B.n257 585
R389 B.n259 B.n258 585
R390 B.n562 B.n561 585
R391 B.n561 B.n560 585
R392 B.n563 B.n256 585
R393 B.n256 B.n255 585
R394 B.n565 B.n564 585
R395 B.n566 B.n565 585
R396 B.n250 B.n249 585
R397 B.n251 B.n250 585
R398 B.n574 B.n573 585
R399 B.n573 B.n572 585
R400 B.n575 B.n248 585
R401 B.n248 B.n247 585
R402 B.n577 B.n576 585
R403 B.n578 B.n577 585
R404 B.n242 B.n241 585
R405 B.n243 B.n242 585
R406 B.n586 B.n585 585
R407 B.n585 B.n584 585
R408 B.n587 B.n240 585
R409 B.n240 B.n239 585
R410 B.n589 B.n588 585
R411 B.n590 B.n589 585
R412 B.n234 B.n233 585
R413 B.n235 B.n234 585
R414 B.n599 B.n598 585
R415 B.n598 B.n597 585
R416 B.n600 B.n232 585
R417 B.n596 B.n232 585
R418 B.n602 B.n601 585
R419 B.n603 B.n602 585
R420 B.n227 B.n226 585
R421 B.n228 B.n227 585
R422 B.n612 B.n611 585
R423 B.n611 B.n610 585
R424 B.n613 B.n225 585
R425 B.n225 B.n224 585
R426 B.n615 B.n614 585
R427 B.n616 B.n615 585
R428 B.n2 B.n0 585
R429 B.n4 B.n2 585
R430 B.n3 B.n1 585
R431 B.n804 B.n3 585
R432 B.n802 B.n801 585
R433 B.n803 B.n802 585
R434 B.n800 B.n9 585
R435 B.n9 B.n8 585
R436 B.n799 B.n798 585
R437 B.n798 B.n797 585
R438 B.n11 B.n10 585
R439 B.n796 B.n11 585
R440 B.n794 B.n793 585
R441 B.n795 B.n794 585
R442 B.n792 B.n15 585
R443 B.n18 B.n15 585
R444 B.n791 B.n790 585
R445 B.n790 B.n789 585
R446 B.n17 B.n16 585
R447 B.n788 B.n17 585
R448 B.n786 B.n785 585
R449 B.n787 B.n786 585
R450 B.n784 B.n23 585
R451 B.n23 B.n22 585
R452 B.n783 B.n782 585
R453 B.n782 B.n781 585
R454 B.n25 B.n24 585
R455 B.n780 B.n25 585
R456 B.n778 B.n777 585
R457 B.n779 B.n778 585
R458 B.n776 B.n30 585
R459 B.n30 B.n29 585
R460 B.n775 B.n774 585
R461 B.n774 B.n773 585
R462 B.n32 B.n31 585
R463 B.n772 B.n32 585
R464 B.n770 B.n769 585
R465 B.n771 B.n770 585
R466 B.n768 B.n37 585
R467 B.n37 B.n36 585
R468 B.n767 B.n766 585
R469 B.n766 B.n765 585
R470 B.n39 B.n38 585
R471 B.n764 B.n39 585
R472 B.n762 B.n761 585
R473 B.n763 B.n762 585
R474 B.n760 B.n44 585
R475 B.n44 B.n43 585
R476 B.n759 B.n758 585
R477 B.n758 B.n757 585
R478 B.n46 B.n45 585
R479 B.n756 B.n46 585
R480 B.n754 B.n753 585
R481 B.n755 B.n754 585
R482 B.n752 B.n51 585
R483 B.n51 B.n50 585
R484 B.n751 B.n750 585
R485 B.n750 B.n749 585
R486 B.n53 B.n52 585
R487 B.n748 B.n53 585
R488 B.n746 B.n745 585
R489 B.n747 B.n746 585
R490 B.n744 B.n58 585
R491 B.n58 B.n57 585
R492 B.n743 B.n742 585
R493 B.n742 B.n741 585
R494 B.n60 B.n59 585
R495 B.n740 B.n60 585
R496 B.n738 B.n737 585
R497 B.n739 B.n738 585
R498 B.n736 B.n64 585
R499 B.n67 B.n64 585
R500 B.n735 B.n734 585
R501 B.n734 B.n733 585
R502 B.n66 B.n65 585
R503 B.n732 B.n66 585
R504 B.n730 B.n729 585
R505 B.n731 B.n730 585
R506 B.n728 B.n72 585
R507 B.n72 B.n71 585
R508 B.n727 B.n726 585
R509 B.n726 B.n725 585
R510 B.n74 B.n73 585
R511 B.n724 B.n74 585
R512 B.n722 B.n721 585
R513 B.n723 B.n722 585
R514 B.n720 B.n79 585
R515 B.n79 B.n78 585
R516 B.n719 B.n718 585
R517 B.n718 B.n717 585
R518 B.n81 B.n80 585
R519 B.n716 B.n81 585
R520 B.n714 B.n713 585
R521 B.n715 B.n714 585
R522 B.n712 B.n86 585
R523 B.n86 B.n85 585
R524 B.n711 B.n710 585
R525 B.n710 B.n709 585
R526 B.n88 B.n87 585
R527 B.n708 B.n88 585
R528 B.n706 B.n705 585
R529 B.n707 B.n706 585
R530 B.n704 B.n93 585
R531 B.n93 B.n92 585
R532 B.n703 B.n702 585
R533 B.n702 B.n701 585
R534 B.n95 B.n94 585
R535 B.n700 B.n95 585
R536 B.n698 B.n697 585
R537 B.n699 B.n698 585
R538 B.n696 B.n100 585
R539 B.n100 B.n99 585
R540 B.n807 B.n806 585
R541 B.n806 B.n805 585
R542 B.n452 B.n327 482.89
R543 B.n694 B.n100 482.89
R544 B.n352 B.n325 482.89
R545 B.n690 B.n126 482.89
R546 B.n692 B.n691 256.663
R547 B.n692 B.n124 256.663
R548 B.n692 B.n123 256.663
R549 B.n692 B.n122 256.663
R550 B.n692 B.n121 256.663
R551 B.n692 B.n120 256.663
R552 B.n692 B.n119 256.663
R553 B.n692 B.n118 256.663
R554 B.n692 B.n117 256.663
R555 B.n692 B.n116 256.663
R556 B.n692 B.n115 256.663
R557 B.n692 B.n114 256.663
R558 B.n692 B.n113 256.663
R559 B.n692 B.n112 256.663
R560 B.n692 B.n111 256.663
R561 B.n692 B.n110 256.663
R562 B.n692 B.n109 256.663
R563 B.n692 B.n108 256.663
R564 B.n692 B.n107 256.663
R565 B.n692 B.n106 256.663
R566 B.n692 B.n105 256.663
R567 B.n692 B.n104 256.663
R568 B.n692 B.n103 256.663
R569 B.n693 B.n692 256.663
R570 B.n451 B.n450 256.663
R571 B.n450 B.n330 256.663
R572 B.n450 B.n331 256.663
R573 B.n450 B.n332 256.663
R574 B.n450 B.n333 256.663
R575 B.n450 B.n334 256.663
R576 B.n450 B.n335 256.663
R577 B.n450 B.n336 256.663
R578 B.n450 B.n337 256.663
R579 B.n450 B.n338 256.663
R580 B.n450 B.n339 256.663
R581 B.n450 B.n340 256.663
R582 B.n450 B.n341 256.663
R583 B.n450 B.n342 256.663
R584 B.n450 B.n343 256.663
R585 B.n450 B.n344 256.663
R586 B.n450 B.n345 256.663
R587 B.n450 B.n346 256.663
R588 B.n450 B.n347 256.663
R589 B.n450 B.n348 256.663
R590 B.n450 B.n349 256.663
R591 B.n450 B.n350 256.663
R592 B.n450 B.n351 256.663
R593 B.n357 B.t12 244.98
R594 B.n354 B.t8 244.98
R595 B.n129 B.t15 244.98
R596 B.n127 B.t19 244.98
R597 B.n456 B.n327 163.367
R598 B.n456 B.n321 163.367
R599 B.n464 B.n321 163.367
R600 B.n464 B.n319 163.367
R601 B.n468 B.n319 163.367
R602 B.n468 B.n313 163.367
R603 B.n476 B.n313 163.367
R604 B.n476 B.n311 163.367
R605 B.n480 B.n311 163.367
R606 B.n480 B.n305 163.367
R607 B.n488 B.n305 163.367
R608 B.n488 B.n303 163.367
R609 B.n492 B.n303 163.367
R610 B.n492 B.n297 163.367
R611 B.n500 B.n297 163.367
R612 B.n500 B.n295 163.367
R613 B.n504 B.n295 163.367
R614 B.n504 B.n289 163.367
R615 B.n513 B.n289 163.367
R616 B.n513 B.n287 163.367
R617 B.n517 B.n287 163.367
R618 B.n517 B.n282 163.367
R619 B.n525 B.n282 163.367
R620 B.n525 B.n280 163.367
R621 B.n529 B.n280 163.367
R622 B.n529 B.n274 163.367
R623 B.n537 B.n274 163.367
R624 B.n537 B.n272 163.367
R625 B.n541 B.n272 163.367
R626 B.n541 B.n266 163.367
R627 B.n549 B.n266 163.367
R628 B.n549 B.n264 163.367
R629 B.n553 B.n264 163.367
R630 B.n553 B.n258 163.367
R631 B.n561 B.n258 163.367
R632 B.n561 B.n256 163.367
R633 B.n565 B.n256 163.367
R634 B.n565 B.n250 163.367
R635 B.n573 B.n250 163.367
R636 B.n573 B.n248 163.367
R637 B.n577 B.n248 163.367
R638 B.n577 B.n242 163.367
R639 B.n585 B.n242 163.367
R640 B.n585 B.n240 163.367
R641 B.n589 B.n240 163.367
R642 B.n589 B.n234 163.367
R643 B.n598 B.n234 163.367
R644 B.n598 B.n232 163.367
R645 B.n602 B.n232 163.367
R646 B.n602 B.n227 163.367
R647 B.n611 B.n227 163.367
R648 B.n611 B.n225 163.367
R649 B.n615 B.n225 163.367
R650 B.n615 B.n2 163.367
R651 B.n806 B.n2 163.367
R652 B.n806 B.n3 163.367
R653 B.n802 B.n3 163.367
R654 B.n802 B.n9 163.367
R655 B.n798 B.n9 163.367
R656 B.n798 B.n11 163.367
R657 B.n794 B.n11 163.367
R658 B.n794 B.n15 163.367
R659 B.n790 B.n15 163.367
R660 B.n790 B.n17 163.367
R661 B.n786 B.n17 163.367
R662 B.n786 B.n23 163.367
R663 B.n782 B.n23 163.367
R664 B.n782 B.n25 163.367
R665 B.n778 B.n25 163.367
R666 B.n778 B.n30 163.367
R667 B.n774 B.n30 163.367
R668 B.n774 B.n32 163.367
R669 B.n770 B.n32 163.367
R670 B.n770 B.n37 163.367
R671 B.n766 B.n37 163.367
R672 B.n766 B.n39 163.367
R673 B.n762 B.n39 163.367
R674 B.n762 B.n44 163.367
R675 B.n758 B.n44 163.367
R676 B.n758 B.n46 163.367
R677 B.n754 B.n46 163.367
R678 B.n754 B.n51 163.367
R679 B.n750 B.n51 163.367
R680 B.n750 B.n53 163.367
R681 B.n746 B.n53 163.367
R682 B.n746 B.n58 163.367
R683 B.n742 B.n58 163.367
R684 B.n742 B.n60 163.367
R685 B.n738 B.n60 163.367
R686 B.n738 B.n64 163.367
R687 B.n734 B.n64 163.367
R688 B.n734 B.n66 163.367
R689 B.n730 B.n66 163.367
R690 B.n730 B.n72 163.367
R691 B.n726 B.n72 163.367
R692 B.n726 B.n74 163.367
R693 B.n722 B.n74 163.367
R694 B.n722 B.n79 163.367
R695 B.n718 B.n79 163.367
R696 B.n718 B.n81 163.367
R697 B.n714 B.n81 163.367
R698 B.n714 B.n86 163.367
R699 B.n710 B.n86 163.367
R700 B.n710 B.n88 163.367
R701 B.n706 B.n88 163.367
R702 B.n706 B.n93 163.367
R703 B.n702 B.n93 163.367
R704 B.n702 B.n95 163.367
R705 B.n698 B.n95 163.367
R706 B.n698 B.n100 163.367
R707 B.n449 B.n329 163.367
R708 B.n449 B.n353 163.367
R709 B.n445 B.n444 163.367
R710 B.n441 B.n440 163.367
R711 B.n437 B.n436 163.367
R712 B.n433 B.n432 163.367
R713 B.n429 B.n428 163.367
R714 B.n425 B.n424 163.367
R715 B.n421 B.n420 163.367
R716 B.n417 B.n416 163.367
R717 B.n413 B.n412 163.367
R718 B.n409 B.n408 163.367
R719 B.n405 B.n404 163.367
R720 B.n401 B.n400 163.367
R721 B.n397 B.n396 163.367
R722 B.n393 B.n392 163.367
R723 B.n389 B.n388 163.367
R724 B.n385 B.n384 163.367
R725 B.n381 B.n380 163.367
R726 B.n377 B.n376 163.367
R727 B.n373 B.n372 163.367
R728 B.n369 B.n368 163.367
R729 B.n365 B.n364 163.367
R730 B.n361 B.n352 163.367
R731 B.n458 B.n325 163.367
R732 B.n458 B.n323 163.367
R733 B.n462 B.n323 163.367
R734 B.n462 B.n317 163.367
R735 B.n470 B.n317 163.367
R736 B.n470 B.n315 163.367
R737 B.n474 B.n315 163.367
R738 B.n474 B.n309 163.367
R739 B.n482 B.n309 163.367
R740 B.n482 B.n307 163.367
R741 B.n486 B.n307 163.367
R742 B.n486 B.n301 163.367
R743 B.n494 B.n301 163.367
R744 B.n494 B.n299 163.367
R745 B.n498 B.n299 163.367
R746 B.n498 B.n293 163.367
R747 B.n506 B.n293 163.367
R748 B.n506 B.n291 163.367
R749 B.n510 B.n291 163.367
R750 B.n510 B.n286 163.367
R751 B.n519 B.n286 163.367
R752 B.n519 B.n284 163.367
R753 B.n523 B.n284 163.367
R754 B.n523 B.n278 163.367
R755 B.n531 B.n278 163.367
R756 B.n531 B.n276 163.367
R757 B.n535 B.n276 163.367
R758 B.n535 B.n270 163.367
R759 B.n543 B.n270 163.367
R760 B.n543 B.n268 163.367
R761 B.n547 B.n268 163.367
R762 B.n547 B.n262 163.367
R763 B.n555 B.n262 163.367
R764 B.n555 B.n260 163.367
R765 B.n559 B.n260 163.367
R766 B.n559 B.n254 163.367
R767 B.n567 B.n254 163.367
R768 B.n567 B.n252 163.367
R769 B.n571 B.n252 163.367
R770 B.n571 B.n246 163.367
R771 B.n579 B.n246 163.367
R772 B.n579 B.n244 163.367
R773 B.n583 B.n244 163.367
R774 B.n583 B.n238 163.367
R775 B.n591 B.n238 163.367
R776 B.n591 B.n236 163.367
R777 B.n595 B.n236 163.367
R778 B.n595 B.n231 163.367
R779 B.n604 B.n231 163.367
R780 B.n604 B.n229 163.367
R781 B.n609 B.n229 163.367
R782 B.n609 B.n223 163.367
R783 B.n617 B.n223 163.367
R784 B.n618 B.n617 163.367
R785 B.n618 B.n5 163.367
R786 B.n6 B.n5 163.367
R787 B.n7 B.n6 163.367
R788 B.n623 B.n7 163.367
R789 B.n623 B.n12 163.367
R790 B.n13 B.n12 163.367
R791 B.n14 B.n13 163.367
R792 B.n628 B.n14 163.367
R793 B.n628 B.n19 163.367
R794 B.n20 B.n19 163.367
R795 B.n21 B.n20 163.367
R796 B.n633 B.n21 163.367
R797 B.n633 B.n26 163.367
R798 B.n27 B.n26 163.367
R799 B.n28 B.n27 163.367
R800 B.n638 B.n28 163.367
R801 B.n638 B.n33 163.367
R802 B.n34 B.n33 163.367
R803 B.n35 B.n34 163.367
R804 B.n643 B.n35 163.367
R805 B.n643 B.n40 163.367
R806 B.n41 B.n40 163.367
R807 B.n42 B.n41 163.367
R808 B.n648 B.n42 163.367
R809 B.n648 B.n47 163.367
R810 B.n48 B.n47 163.367
R811 B.n49 B.n48 163.367
R812 B.n653 B.n49 163.367
R813 B.n653 B.n54 163.367
R814 B.n55 B.n54 163.367
R815 B.n56 B.n55 163.367
R816 B.n658 B.n56 163.367
R817 B.n658 B.n61 163.367
R818 B.n62 B.n61 163.367
R819 B.n63 B.n62 163.367
R820 B.n663 B.n63 163.367
R821 B.n663 B.n68 163.367
R822 B.n69 B.n68 163.367
R823 B.n70 B.n69 163.367
R824 B.n668 B.n70 163.367
R825 B.n668 B.n75 163.367
R826 B.n76 B.n75 163.367
R827 B.n77 B.n76 163.367
R828 B.n673 B.n77 163.367
R829 B.n673 B.n82 163.367
R830 B.n83 B.n82 163.367
R831 B.n84 B.n83 163.367
R832 B.n678 B.n84 163.367
R833 B.n678 B.n89 163.367
R834 B.n90 B.n89 163.367
R835 B.n91 B.n90 163.367
R836 B.n683 B.n91 163.367
R837 B.n683 B.n96 163.367
R838 B.n97 B.n96 163.367
R839 B.n98 B.n97 163.367
R840 B.n126 B.n98 163.367
R841 B.n131 B.n102 163.367
R842 B.n135 B.n134 163.367
R843 B.n139 B.n138 163.367
R844 B.n143 B.n142 163.367
R845 B.n147 B.n146 163.367
R846 B.n151 B.n150 163.367
R847 B.n155 B.n154 163.367
R848 B.n159 B.n158 163.367
R849 B.n163 B.n162 163.367
R850 B.n168 B.n167 163.367
R851 B.n172 B.n171 163.367
R852 B.n176 B.n175 163.367
R853 B.n180 B.n179 163.367
R854 B.n184 B.n183 163.367
R855 B.n189 B.n188 163.367
R856 B.n193 B.n192 163.367
R857 B.n197 B.n196 163.367
R858 B.n201 B.n200 163.367
R859 B.n205 B.n204 163.367
R860 B.n209 B.n208 163.367
R861 B.n213 B.n212 163.367
R862 B.n217 B.n216 163.367
R863 B.n219 B.n125 163.367
R864 B.n450 B.n326 143.006
R865 B.n692 B.n99 143.006
R866 B.n357 B.t14 137.886
R867 B.n127 B.t20 137.886
R868 B.n354 B.t11 137.881
R869 B.n129 B.t17 137.881
R870 B.n457 B.n326 77.7956
R871 B.n457 B.n322 77.7956
R872 B.n463 B.n322 77.7956
R873 B.n463 B.n318 77.7956
R874 B.n469 B.n318 77.7956
R875 B.n469 B.n314 77.7956
R876 B.n475 B.n314 77.7956
R877 B.n481 B.n310 77.7956
R878 B.n481 B.n306 77.7956
R879 B.n487 B.n306 77.7956
R880 B.n487 B.n302 77.7956
R881 B.n493 B.n302 77.7956
R882 B.n493 B.n298 77.7956
R883 B.n499 B.n298 77.7956
R884 B.n499 B.n294 77.7956
R885 B.n505 B.n294 77.7956
R886 B.n505 B.n290 77.7956
R887 B.n512 B.n290 77.7956
R888 B.n512 B.n511 77.7956
R889 B.n518 B.n283 77.7956
R890 B.n524 B.n283 77.7956
R891 B.n524 B.n279 77.7956
R892 B.n530 B.n279 77.7956
R893 B.n530 B.n275 77.7956
R894 B.n536 B.n275 77.7956
R895 B.n536 B.n271 77.7956
R896 B.n542 B.n271 77.7956
R897 B.n548 B.n267 77.7956
R898 B.n548 B.n263 77.7956
R899 B.n554 B.n263 77.7956
R900 B.n554 B.n259 77.7956
R901 B.n560 B.n259 77.7956
R902 B.n560 B.n255 77.7956
R903 B.n566 B.n255 77.7956
R904 B.n566 B.n251 77.7956
R905 B.n572 B.n251 77.7956
R906 B.n578 B.n247 77.7956
R907 B.n578 B.n243 77.7956
R908 B.n584 B.n243 77.7956
R909 B.n584 B.n239 77.7956
R910 B.n590 B.n239 77.7956
R911 B.n590 B.n235 77.7956
R912 B.n597 B.n235 77.7956
R913 B.n597 B.n596 77.7956
R914 B.n603 B.n228 77.7956
R915 B.n610 B.n228 77.7956
R916 B.n610 B.n224 77.7956
R917 B.n616 B.n224 77.7956
R918 B.n616 B.n4 77.7956
R919 B.n805 B.n4 77.7956
R920 B.n805 B.n804 77.7956
R921 B.n804 B.n803 77.7956
R922 B.n803 B.n8 77.7956
R923 B.n797 B.n8 77.7956
R924 B.n797 B.n796 77.7956
R925 B.n796 B.n795 77.7956
R926 B.n789 B.n18 77.7956
R927 B.n789 B.n788 77.7956
R928 B.n788 B.n787 77.7956
R929 B.n787 B.n22 77.7956
R930 B.n781 B.n22 77.7956
R931 B.n781 B.n780 77.7956
R932 B.n780 B.n779 77.7956
R933 B.n779 B.n29 77.7956
R934 B.n773 B.n772 77.7956
R935 B.n772 B.n771 77.7956
R936 B.n771 B.n36 77.7956
R937 B.n765 B.n36 77.7956
R938 B.n765 B.n764 77.7956
R939 B.n764 B.n763 77.7956
R940 B.n763 B.n43 77.7956
R941 B.n757 B.n43 77.7956
R942 B.n757 B.n756 77.7956
R943 B.n755 B.n50 77.7956
R944 B.n749 B.n50 77.7956
R945 B.n749 B.n748 77.7956
R946 B.n748 B.n747 77.7956
R947 B.n747 B.n57 77.7956
R948 B.n741 B.n57 77.7956
R949 B.n741 B.n740 77.7956
R950 B.n740 B.n739 77.7956
R951 B.n733 B.n67 77.7956
R952 B.n733 B.n732 77.7956
R953 B.n732 B.n731 77.7956
R954 B.n731 B.n71 77.7956
R955 B.n725 B.n71 77.7956
R956 B.n725 B.n724 77.7956
R957 B.n724 B.n723 77.7956
R958 B.n723 B.n78 77.7956
R959 B.n717 B.n78 77.7956
R960 B.n717 B.n716 77.7956
R961 B.n716 B.n715 77.7956
R962 B.n715 B.n85 77.7956
R963 B.n709 B.n708 77.7956
R964 B.n708 B.n707 77.7956
R965 B.n707 B.n92 77.7956
R966 B.n701 B.n92 77.7956
R967 B.n701 B.n700 77.7956
R968 B.n700 B.n699 77.7956
R969 B.n699 B.n99 77.7956
R970 B.n358 B.t13 76.0192
R971 B.n128 B.t21 76.0192
R972 B.n355 B.t10 76.0153
R973 B.n130 B.t18 76.0153
R974 B.n475 B.t9 75.5075
R975 B.n709 B.t16 75.5075
R976 B.n542 B.t5 73.2194
R977 B.t7 B.n755 73.2194
R978 B.n452 B.n451 71.676
R979 B.n353 B.n330 71.676
R980 B.n444 B.n331 71.676
R981 B.n440 B.n332 71.676
R982 B.n436 B.n333 71.676
R983 B.n432 B.n334 71.676
R984 B.n428 B.n335 71.676
R985 B.n424 B.n336 71.676
R986 B.n420 B.n337 71.676
R987 B.n416 B.n338 71.676
R988 B.n412 B.n339 71.676
R989 B.n408 B.n340 71.676
R990 B.n404 B.n341 71.676
R991 B.n400 B.n342 71.676
R992 B.n396 B.n343 71.676
R993 B.n392 B.n344 71.676
R994 B.n388 B.n345 71.676
R995 B.n384 B.n346 71.676
R996 B.n380 B.n347 71.676
R997 B.n376 B.n348 71.676
R998 B.n372 B.n349 71.676
R999 B.n368 B.n350 71.676
R1000 B.n364 B.n351 71.676
R1001 B.n694 B.n693 71.676
R1002 B.n131 B.n103 71.676
R1003 B.n135 B.n104 71.676
R1004 B.n139 B.n105 71.676
R1005 B.n143 B.n106 71.676
R1006 B.n147 B.n107 71.676
R1007 B.n151 B.n108 71.676
R1008 B.n155 B.n109 71.676
R1009 B.n159 B.n110 71.676
R1010 B.n163 B.n111 71.676
R1011 B.n168 B.n112 71.676
R1012 B.n172 B.n113 71.676
R1013 B.n176 B.n114 71.676
R1014 B.n180 B.n115 71.676
R1015 B.n184 B.n116 71.676
R1016 B.n189 B.n117 71.676
R1017 B.n193 B.n118 71.676
R1018 B.n197 B.n119 71.676
R1019 B.n201 B.n120 71.676
R1020 B.n205 B.n121 71.676
R1021 B.n209 B.n122 71.676
R1022 B.n213 B.n123 71.676
R1023 B.n217 B.n124 71.676
R1024 B.n691 B.n125 71.676
R1025 B.n691 B.n690 71.676
R1026 B.n219 B.n124 71.676
R1027 B.n216 B.n123 71.676
R1028 B.n212 B.n122 71.676
R1029 B.n208 B.n121 71.676
R1030 B.n204 B.n120 71.676
R1031 B.n200 B.n119 71.676
R1032 B.n196 B.n118 71.676
R1033 B.n192 B.n117 71.676
R1034 B.n188 B.n116 71.676
R1035 B.n183 B.n115 71.676
R1036 B.n179 B.n114 71.676
R1037 B.n175 B.n113 71.676
R1038 B.n171 B.n112 71.676
R1039 B.n167 B.n111 71.676
R1040 B.n162 B.n110 71.676
R1041 B.n158 B.n109 71.676
R1042 B.n154 B.n108 71.676
R1043 B.n150 B.n107 71.676
R1044 B.n146 B.n106 71.676
R1045 B.n142 B.n105 71.676
R1046 B.n138 B.n104 71.676
R1047 B.n134 B.n103 71.676
R1048 B.n693 B.n102 71.676
R1049 B.n451 B.n329 71.676
R1050 B.n445 B.n330 71.676
R1051 B.n441 B.n331 71.676
R1052 B.n437 B.n332 71.676
R1053 B.n433 B.n333 71.676
R1054 B.n429 B.n334 71.676
R1055 B.n425 B.n335 71.676
R1056 B.n421 B.n336 71.676
R1057 B.n417 B.n337 71.676
R1058 B.n413 B.n338 71.676
R1059 B.n409 B.n339 71.676
R1060 B.n405 B.n340 71.676
R1061 B.n401 B.n341 71.676
R1062 B.n397 B.n342 71.676
R1063 B.n393 B.n343 71.676
R1064 B.n389 B.n344 71.676
R1065 B.n385 B.n345 71.676
R1066 B.n381 B.n346 71.676
R1067 B.n377 B.n347 71.676
R1068 B.n373 B.n348 71.676
R1069 B.n369 B.n349 71.676
R1070 B.n365 B.n350 71.676
R1071 B.n361 B.n351 71.676
R1072 B.n358 B.n357 61.8672
R1073 B.n355 B.n354 61.8672
R1074 B.n130 B.n129 61.8672
R1075 B.n128 B.n127 61.8672
R1076 B.n359 B.n358 59.5399
R1077 B.n356 B.n355 59.5399
R1078 B.n165 B.n130 59.5399
R1079 B.n186 B.n128 59.5399
R1080 B.n596 B.t6 54.9147
R1081 B.n18 B.t2 54.9147
R1082 B.t4 B.n247 52.6266
R1083 B.t1 B.n29 52.6266
R1084 B.n511 B.t0 43.4742
R1085 B.n67 B.t3 43.4742
R1086 B.n518 B.t0 34.3219
R1087 B.n739 B.t3 34.3219
R1088 B.n696 B.n695 31.3761
R1089 B.n689 B.n688 31.3761
R1090 B.n360 B.n324 31.3761
R1091 B.n454 B.n453 31.3761
R1092 B.n572 B.t4 25.1695
R1093 B.n773 B.t1 25.1695
R1094 B.n603 B.t6 22.8814
R1095 B.n795 B.t2 22.8814
R1096 B B.n807 18.0485
R1097 B.n695 B.n101 10.6151
R1098 B.n132 B.n101 10.6151
R1099 B.n133 B.n132 10.6151
R1100 B.n136 B.n133 10.6151
R1101 B.n137 B.n136 10.6151
R1102 B.n140 B.n137 10.6151
R1103 B.n141 B.n140 10.6151
R1104 B.n144 B.n141 10.6151
R1105 B.n145 B.n144 10.6151
R1106 B.n148 B.n145 10.6151
R1107 B.n149 B.n148 10.6151
R1108 B.n152 B.n149 10.6151
R1109 B.n153 B.n152 10.6151
R1110 B.n156 B.n153 10.6151
R1111 B.n157 B.n156 10.6151
R1112 B.n160 B.n157 10.6151
R1113 B.n161 B.n160 10.6151
R1114 B.n164 B.n161 10.6151
R1115 B.n169 B.n166 10.6151
R1116 B.n170 B.n169 10.6151
R1117 B.n173 B.n170 10.6151
R1118 B.n174 B.n173 10.6151
R1119 B.n177 B.n174 10.6151
R1120 B.n178 B.n177 10.6151
R1121 B.n181 B.n178 10.6151
R1122 B.n182 B.n181 10.6151
R1123 B.n185 B.n182 10.6151
R1124 B.n190 B.n187 10.6151
R1125 B.n191 B.n190 10.6151
R1126 B.n194 B.n191 10.6151
R1127 B.n195 B.n194 10.6151
R1128 B.n198 B.n195 10.6151
R1129 B.n199 B.n198 10.6151
R1130 B.n202 B.n199 10.6151
R1131 B.n203 B.n202 10.6151
R1132 B.n206 B.n203 10.6151
R1133 B.n207 B.n206 10.6151
R1134 B.n210 B.n207 10.6151
R1135 B.n211 B.n210 10.6151
R1136 B.n214 B.n211 10.6151
R1137 B.n215 B.n214 10.6151
R1138 B.n218 B.n215 10.6151
R1139 B.n220 B.n218 10.6151
R1140 B.n221 B.n220 10.6151
R1141 B.n689 B.n221 10.6151
R1142 B.n459 B.n324 10.6151
R1143 B.n460 B.n459 10.6151
R1144 B.n461 B.n460 10.6151
R1145 B.n461 B.n316 10.6151
R1146 B.n471 B.n316 10.6151
R1147 B.n472 B.n471 10.6151
R1148 B.n473 B.n472 10.6151
R1149 B.n473 B.n308 10.6151
R1150 B.n483 B.n308 10.6151
R1151 B.n484 B.n483 10.6151
R1152 B.n485 B.n484 10.6151
R1153 B.n485 B.n300 10.6151
R1154 B.n495 B.n300 10.6151
R1155 B.n496 B.n495 10.6151
R1156 B.n497 B.n496 10.6151
R1157 B.n497 B.n292 10.6151
R1158 B.n507 B.n292 10.6151
R1159 B.n508 B.n507 10.6151
R1160 B.n509 B.n508 10.6151
R1161 B.n509 B.n285 10.6151
R1162 B.n520 B.n285 10.6151
R1163 B.n521 B.n520 10.6151
R1164 B.n522 B.n521 10.6151
R1165 B.n522 B.n277 10.6151
R1166 B.n532 B.n277 10.6151
R1167 B.n533 B.n532 10.6151
R1168 B.n534 B.n533 10.6151
R1169 B.n534 B.n269 10.6151
R1170 B.n544 B.n269 10.6151
R1171 B.n545 B.n544 10.6151
R1172 B.n546 B.n545 10.6151
R1173 B.n546 B.n261 10.6151
R1174 B.n556 B.n261 10.6151
R1175 B.n557 B.n556 10.6151
R1176 B.n558 B.n557 10.6151
R1177 B.n558 B.n253 10.6151
R1178 B.n568 B.n253 10.6151
R1179 B.n569 B.n568 10.6151
R1180 B.n570 B.n569 10.6151
R1181 B.n570 B.n245 10.6151
R1182 B.n580 B.n245 10.6151
R1183 B.n581 B.n580 10.6151
R1184 B.n582 B.n581 10.6151
R1185 B.n582 B.n237 10.6151
R1186 B.n592 B.n237 10.6151
R1187 B.n593 B.n592 10.6151
R1188 B.n594 B.n593 10.6151
R1189 B.n594 B.n230 10.6151
R1190 B.n605 B.n230 10.6151
R1191 B.n606 B.n605 10.6151
R1192 B.n608 B.n606 10.6151
R1193 B.n608 B.n607 10.6151
R1194 B.n607 B.n222 10.6151
R1195 B.n619 B.n222 10.6151
R1196 B.n620 B.n619 10.6151
R1197 B.n621 B.n620 10.6151
R1198 B.n622 B.n621 10.6151
R1199 B.n624 B.n622 10.6151
R1200 B.n625 B.n624 10.6151
R1201 B.n626 B.n625 10.6151
R1202 B.n627 B.n626 10.6151
R1203 B.n629 B.n627 10.6151
R1204 B.n630 B.n629 10.6151
R1205 B.n631 B.n630 10.6151
R1206 B.n632 B.n631 10.6151
R1207 B.n634 B.n632 10.6151
R1208 B.n635 B.n634 10.6151
R1209 B.n636 B.n635 10.6151
R1210 B.n637 B.n636 10.6151
R1211 B.n639 B.n637 10.6151
R1212 B.n640 B.n639 10.6151
R1213 B.n641 B.n640 10.6151
R1214 B.n642 B.n641 10.6151
R1215 B.n644 B.n642 10.6151
R1216 B.n645 B.n644 10.6151
R1217 B.n646 B.n645 10.6151
R1218 B.n647 B.n646 10.6151
R1219 B.n649 B.n647 10.6151
R1220 B.n650 B.n649 10.6151
R1221 B.n651 B.n650 10.6151
R1222 B.n652 B.n651 10.6151
R1223 B.n654 B.n652 10.6151
R1224 B.n655 B.n654 10.6151
R1225 B.n656 B.n655 10.6151
R1226 B.n657 B.n656 10.6151
R1227 B.n659 B.n657 10.6151
R1228 B.n660 B.n659 10.6151
R1229 B.n661 B.n660 10.6151
R1230 B.n662 B.n661 10.6151
R1231 B.n664 B.n662 10.6151
R1232 B.n665 B.n664 10.6151
R1233 B.n666 B.n665 10.6151
R1234 B.n667 B.n666 10.6151
R1235 B.n669 B.n667 10.6151
R1236 B.n670 B.n669 10.6151
R1237 B.n671 B.n670 10.6151
R1238 B.n672 B.n671 10.6151
R1239 B.n674 B.n672 10.6151
R1240 B.n675 B.n674 10.6151
R1241 B.n676 B.n675 10.6151
R1242 B.n677 B.n676 10.6151
R1243 B.n679 B.n677 10.6151
R1244 B.n680 B.n679 10.6151
R1245 B.n681 B.n680 10.6151
R1246 B.n682 B.n681 10.6151
R1247 B.n684 B.n682 10.6151
R1248 B.n685 B.n684 10.6151
R1249 B.n686 B.n685 10.6151
R1250 B.n687 B.n686 10.6151
R1251 B.n688 B.n687 10.6151
R1252 B.n453 B.n328 10.6151
R1253 B.n448 B.n328 10.6151
R1254 B.n448 B.n447 10.6151
R1255 B.n447 B.n446 10.6151
R1256 B.n446 B.n443 10.6151
R1257 B.n443 B.n442 10.6151
R1258 B.n442 B.n439 10.6151
R1259 B.n439 B.n438 10.6151
R1260 B.n438 B.n435 10.6151
R1261 B.n435 B.n434 10.6151
R1262 B.n434 B.n431 10.6151
R1263 B.n431 B.n430 10.6151
R1264 B.n430 B.n427 10.6151
R1265 B.n427 B.n426 10.6151
R1266 B.n426 B.n423 10.6151
R1267 B.n423 B.n422 10.6151
R1268 B.n422 B.n419 10.6151
R1269 B.n419 B.n418 10.6151
R1270 B.n415 B.n414 10.6151
R1271 B.n414 B.n411 10.6151
R1272 B.n411 B.n410 10.6151
R1273 B.n410 B.n407 10.6151
R1274 B.n407 B.n406 10.6151
R1275 B.n406 B.n403 10.6151
R1276 B.n403 B.n402 10.6151
R1277 B.n402 B.n399 10.6151
R1278 B.n399 B.n398 10.6151
R1279 B.n395 B.n394 10.6151
R1280 B.n394 B.n391 10.6151
R1281 B.n391 B.n390 10.6151
R1282 B.n390 B.n387 10.6151
R1283 B.n387 B.n386 10.6151
R1284 B.n386 B.n383 10.6151
R1285 B.n383 B.n382 10.6151
R1286 B.n382 B.n379 10.6151
R1287 B.n379 B.n378 10.6151
R1288 B.n378 B.n375 10.6151
R1289 B.n375 B.n374 10.6151
R1290 B.n374 B.n371 10.6151
R1291 B.n371 B.n370 10.6151
R1292 B.n370 B.n367 10.6151
R1293 B.n367 B.n366 10.6151
R1294 B.n366 B.n363 10.6151
R1295 B.n363 B.n362 10.6151
R1296 B.n362 B.n360 10.6151
R1297 B.n455 B.n454 10.6151
R1298 B.n455 B.n320 10.6151
R1299 B.n465 B.n320 10.6151
R1300 B.n466 B.n465 10.6151
R1301 B.n467 B.n466 10.6151
R1302 B.n467 B.n312 10.6151
R1303 B.n477 B.n312 10.6151
R1304 B.n478 B.n477 10.6151
R1305 B.n479 B.n478 10.6151
R1306 B.n479 B.n304 10.6151
R1307 B.n489 B.n304 10.6151
R1308 B.n490 B.n489 10.6151
R1309 B.n491 B.n490 10.6151
R1310 B.n491 B.n296 10.6151
R1311 B.n501 B.n296 10.6151
R1312 B.n502 B.n501 10.6151
R1313 B.n503 B.n502 10.6151
R1314 B.n503 B.n288 10.6151
R1315 B.n514 B.n288 10.6151
R1316 B.n515 B.n514 10.6151
R1317 B.n516 B.n515 10.6151
R1318 B.n516 B.n281 10.6151
R1319 B.n526 B.n281 10.6151
R1320 B.n527 B.n526 10.6151
R1321 B.n528 B.n527 10.6151
R1322 B.n528 B.n273 10.6151
R1323 B.n538 B.n273 10.6151
R1324 B.n539 B.n538 10.6151
R1325 B.n540 B.n539 10.6151
R1326 B.n540 B.n265 10.6151
R1327 B.n550 B.n265 10.6151
R1328 B.n551 B.n550 10.6151
R1329 B.n552 B.n551 10.6151
R1330 B.n552 B.n257 10.6151
R1331 B.n562 B.n257 10.6151
R1332 B.n563 B.n562 10.6151
R1333 B.n564 B.n563 10.6151
R1334 B.n564 B.n249 10.6151
R1335 B.n574 B.n249 10.6151
R1336 B.n575 B.n574 10.6151
R1337 B.n576 B.n575 10.6151
R1338 B.n576 B.n241 10.6151
R1339 B.n586 B.n241 10.6151
R1340 B.n587 B.n586 10.6151
R1341 B.n588 B.n587 10.6151
R1342 B.n588 B.n233 10.6151
R1343 B.n599 B.n233 10.6151
R1344 B.n600 B.n599 10.6151
R1345 B.n601 B.n600 10.6151
R1346 B.n601 B.n226 10.6151
R1347 B.n612 B.n226 10.6151
R1348 B.n613 B.n612 10.6151
R1349 B.n614 B.n613 10.6151
R1350 B.n614 B.n0 10.6151
R1351 B.n801 B.n1 10.6151
R1352 B.n801 B.n800 10.6151
R1353 B.n800 B.n799 10.6151
R1354 B.n799 B.n10 10.6151
R1355 B.n793 B.n10 10.6151
R1356 B.n793 B.n792 10.6151
R1357 B.n792 B.n791 10.6151
R1358 B.n791 B.n16 10.6151
R1359 B.n785 B.n16 10.6151
R1360 B.n785 B.n784 10.6151
R1361 B.n784 B.n783 10.6151
R1362 B.n783 B.n24 10.6151
R1363 B.n777 B.n24 10.6151
R1364 B.n777 B.n776 10.6151
R1365 B.n776 B.n775 10.6151
R1366 B.n775 B.n31 10.6151
R1367 B.n769 B.n31 10.6151
R1368 B.n769 B.n768 10.6151
R1369 B.n768 B.n767 10.6151
R1370 B.n767 B.n38 10.6151
R1371 B.n761 B.n38 10.6151
R1372 B.n761 B.n760 10.6151
R1373 B.n760 B.n759 10.6151
R1374 B.n759 B.n45 10.6151
R1375 B.n753 B.n45 10.6151
R1376 B.n753 B.n752 10.6151
R1377 B.n752 B.n751 10.6151
R1378 B.n751 B.n52 10.6151
R1379 B.n745 B.n52 10.6151
R1380 B.n745 B.n744 10.6151
R1381 B.n744 B.n743 10.6151
R1382 B.n743 B.n59 10.6151
R1383 B.n737 B.n59 10.6151
R1384 B.n737 B.n736 10.6151
R1385 B.n736 B.n735 10.6151
R1386 B.n735 B.n65 10.6151
R1387 B.n729 B.n65 10.6151
R1388 B.n729 B.n728 10.6151
R1389 B.n728 B.n727 10.6151
R1390 B.n727 B.n73 10.6151
R1391 B.n721 B.n73 10.6151
R1392 B.n721 B.n720 10.6151
R1393 B.n720 B.n719 10.6151
R1394 B.n719 B.n80 10.6151
R1395 B.n713 B.n80 10.6151
R1396 B.n713 B.n712 10.6151
R1397 B.n712 B.n711 10.6151
R1398 B.n711 B.n87 10.6151
R1399 B.n705 B.n87 10.6151
R1400 B.n705 B.n704 10.6151
R1401 B.n704 B.n703 10.6151
R1402 B.n703 B.n94 10.6151
R1403 B.n697 B.n94 10.6151
R1404 B.n697 B.n696 10.6151
R1405 B.n165 B.n164 9.36635
R1406 B.n187 B.n186 9.36635
R1407 B.n418 B.n356 9.36635
R1408 B.n395 B.n359 9.36635
R1409 B.t5 B.n267 4.57668
R1410 B.n756 B.t7 4.57668
R1411 B.n807 B.n0 2.81026
R1412 B.n807 B.n1 2.81026
R1413 B.t9 B.n310 2.28859
R1414 B.t16 B.n85 2.28859
R1415 B.n166 B.n165 1.24928
R1416 B.n186 B.n185 1.24928
R1417 B.n415 B.n356 1.24928
R1418 B.n398 B.n359 1.24928
R1419 VP.n19 VP.n16 161.3
R1420 VP.n21 VP.n20 161.3
R1421 VP.n22 VP.n15 161.3
R1422 VP.n24 VP.n23 161.3
R1423 VP.n25 VP.n14 161.3
R1424 VP.n28 VP.n27 161.3
R1425 VP.n29 VP.n13 161.3
R1426 VP.n31 VP.n30 161.3
R1427 VP.n32 VP.n12 161.3
R1428 VP.n34 VP.n33 161.3
R1429 VP.n35 VP.n11 161.3
R1430 VP.n37 VP.n36 161.3
R1431 VP.n38 VP.n10 161.3
R1432 VP.n74 VP.n0 161.3
R1433 VP.n73 VP.n72 161.3
R1434 VP.n71 VP.n1 161.3
R1435 VP.n70 VP.n69 161.3
R1436 VP.n68 VP.n2 161.3
R1437 VP.n67 VP.n66 161.3
R1438 VP.n65 VP.n3 161.3
R1439 VP.n64 VP.n63 161.3
R1440 VP.n61 VP.n4 161.3
R1441 VP.n60 VP.n59 161.3
R1442 VP.n58 VP.n5 161.3
R1443 VP.n57 VP.n56 161.3
R1444 VP.n55 VP.n6 161.3
R1445 VP.n53 VP.n52 161.3
R1446 VP.n51 VP.n7 161.3
R1447 VP.n50 VP.n49 161.3
R1448 VP.n48 VP.n8 161.3
R1449 VP.n47 VP.n46 161.3
R1450 VP.n45 VP.n9 161.3
R1451 VP.n44 VP.n43 161.3
R1452 VP.n42 VP.n41 109.186
R1453 VP.n76 VP.n75 109.186
R1454 VP.n40 VP.n39 109.186
R1455 VP.n17 VP.t7 69.3223
R1456 VP.n18 VP.n17 56.9625
R1457 VP.n60 VP.n5 56.5617
R1458 VP.n24 VP.n15 56.5617
R1459 VP.n49 VP.n48 46.3896
R1460 VP.n69 VP.n68 46.3896
R1461 VP.n33 VP.n32 46.3896
R1462 VP.n41 VP.n40 46.2648
R1463 VP.n42 VP.t0 36.5718
R1464 VP.n54 VP.t1 36.5718
R1465 VP.n62 VP.t6 36.5718
R1466 VP.n75 VP.t5 36.5718
R1467 VP.n39 VP.t2 36.5718
R1468 VP.n26 VP.t3 36.5718
R1469 VP.n18 VP.t4 36.5718
R1470 VP.n48 VP.n47 34.7644
R1471 VP.n69 VP.n1 34.7644
R1472 VP.n33 VP.n11 34.7644
R1473 VP.n43 VP.n9 24.5923
R1474 VP.n47 VP.n9 24.5923
R1475 VP.n49 VP.n7 24.5923
R1476 VP.n53 VP.n7 24.5923
R1477 VP.n56 VP.n55 24.5923
R1478 VP.n56 VP.n5 24.5923
R1479 VP.n61 VP.n60 24.5923
R1480 VP.n63 VP.n61 24.5923
R1481 VP.n67 VP.n3 24.5923
R1482 VP.n68 VP.n67 24.5923
R1483 VP.n73 VP.n1 24.5923
R1484 VP.n74 VP.n73 24.5923
R1485 VP.n37 VP.n11 24.5923
R1486 VP.n38 VP.n37 24.5923
R1487 VP.n25 VP.n24 24.5923
R1488 VP.n27 VP.n25 24.5923
R1489 VP.n31 VP.n13 24.5923
R1490 VP.n32 VP.n31 24.5923
R1491 VP.n20 VP.n19 24.5923
R1492 VP.n20 VP.n15 24.5923
R1493 VP.n55 VP.n54 16.9689
R1494 VP.n63 VP.n62 16.9689
R1495 VP.n27 VP.n26 16.9689
R1496 VP.n19 VP.n18 16.9689
R1497 VP.n54 VP.n53 7.62397
R1498 VP.n62 VP.n3 7.62397
R1499 VP.n26 VP.n13 7.62397
R1500 VP.n17 VP.n16 5.10887
R1501 VP.n43 VP.n42 1.72193
R1502 VP.n75 VP.n74 1.72193
R1503 VP.n39 VP.n38 1.72193
R1504 VP.n40 VP.n10 0.278335
R1505 VP.n44 VP.n41 0.278335
R1506 VP.n76 VP.n0 0.278335
R1507 VP.n21 VP.n16 0.189894
R1508 VP.n22 VP.n21 0.189894
R1509 VP.n23 VP.n22 0.189894
R1510 VP.n23 VP.n14 0.189894
R1511 VP.n28 VP.n14 0.189894
R1512 VP.n29 VP.n28 0.189894
R1513 VP.n30 VP.n29 0.189894
R1514 VP.n30 VP.n12 0.189894
R1515 VP.n34 VP.n12 0.189894
R1516 VP.n35 VP.n34 0.189894
R1517 VP.n36 VP.n35 0.189894
R1518 VP.n36 VP.n10 0.189894
R1519 VP.n45 VP.n44 0.189894
R1520 VP.n46 VP.n45 0.189894
R1521 VP.n46 VP.n8 0.189894
R1522 VP.n50 VP.n8 0.189894
R1523 VP.n51 VP.n50 0.189894
R1524 VP.n52 VP.n51 0.189894
R1525 VP.n52 VP.n6 0.189894
R1526 VP.n57 VP.n6 0.189894
R1527 VP.n58 VP.n57 0.189894
R1528 VP.n59 VP.n58 0.189894
R1529 VP.n59 VP.n4 0.189894
R1530 VP.n64 VP.n4 0.189894
R1531 VP.n65 VP.n64 0.189894
R1532 VP.n66 VP.n65 0.189894
R1533 VP.n66 VP.n2 0.189894
R1534 VP.n70 VP.n2 0.189894
R1535 VP.n71 VP.n70 0.189894
R1536 VP.n72 VP.n71 0.189894
R1537 VP.n72 VP.n0 0.189894
R1538 VP VP.n76 0.153485
R1539 VDD1 VDD1.n0 76.0668
R1540 VDD1.n3 VDD1.n2 75.953
R1541 VDD1.n3 VDD1.n1 75.953
R1542 VDD1.n5 VDD1.n4 74.6334
R1543 VDD1.n5 VDD1.n3 40.4147
R1544 VDD1.n4 VDD1.t0 4.56271
R1545 VDD1.n4 VDD1.t5 4.56271
R1546 VDD1.n0 VDD1.t4 4.56271
R1547 VDD1.n0 VDD1.t7 4.56271
R1548 VDD1.n2 VDD1.t1 4.56271
R1549 VDD1.n2 VDD1.t2 4.56271
R1550 VDD1.n1 VDD1.t3 4.56271
R1551 VDD1.n1 VDD1.t6 4.56271
R1552 VDD1 VDD1.n5 1.31731
R1553 VTAIL.n11 VTAIL.t4 62.517
R1554 VTAIL.n10 VTAIL.t12 62.517
R1555 VTAIL.n7 VTAIL.t15 62.517
R1556 VTAIL.n14 VTAIL.t9 62.5168
R1557 VTAIL.n15 VTAIL.t13 62.5168
R1558 VTAIL.n2 VTAIL.t3 62.5168
R1559 VTAIL.n3 VTAIL.t6 62.5168
R1560 VTAIL.n6 VTAIL.t11 62.5168
R1561 VTAIL.n13 VTAIL.n12 57.9548
R1562 VTAIL.n9 VTAIL.n8 57.9548
R1563 VTAIL.n1 VTAIL.n0 57.9546
R1564 VTAIL.n5 VTAIL.n4 57.9546
R1565 VTAIL.n15 VTAIL.n14 18.8583
R1566 VTAIL.n7 VTAIL.n6 18.8583
R1567 VTAIL.n0 VTAIL.t14 4.56271
R1568 VTAIL.n0 VTAIL.t1 4.56271
R1569 VTAIL.n4 VTAIL.t10 4.56271
R1570 VTAIL.n4 VTAIL.t5 4.56271
R1571 VTAIL.n12 VTAIL.t7 4.56271
R1572 VTAIL.n12 VTAIL.t8 4.56271
R1573 VTAIL.n8 VTAIL.t2 4.56271
R1574 VTAIL.n8 VTAIL.t0 4.56271
R1575 VTAIL.n9 VTAIL.n7 2.7505
R1576 VTAIL.n10 VTAIL.n9 2.7505
R1577 VTAIL.n13 VTAIL.n11 2.7505
R1578 VTAIL.n14 VTAIL.n13 2.7505
R1579 VTAIL.n6 VTAIL.n5 2.7505
R1580 VTAIL.n5 VTAIL.n3 2.7505
R1581 VTAIL.n2 VTAIL.n1 2.7505
R1582 VTAIL VTAIL.n15 2.69231
R1583 VTAIL.n11 VTAIL.n10 0.470328
R1584 VTAIL.n3 VTAIL.n2 0.470328
R1585 VTAIL VTAIL.n1 0.0586897
R1586 VN.n59 VN.n31 161.3
R1587 VN.n58 VN.n57 161.3
R1588 VN.n56 VN.n32 161.3
R1589 VN.n55 VN.n54 161.3
R1590 VN.n53 VN.n33 161.3
R1591 VN.n52 VN.n51 161.3
R1592 VN.n50 VN.n34 161.3
R1593 VN.n49 VN.n48 161.3
R1594 VN.n47 VN.n35 161.3
R1595 VN.n46 VN.n45 161.3
R1596 VN.n44 VN.n37 161.3
R1597 VN.n43 VN.n42 161.3
R1598 VN.n41 VN.n38 161.3
R1599 VN.n28 VN.n0 161.3
R1600 VN.n27 VN.n26 161.3
R1601 VN.n25 VN.n1 161.3
R1602 VN.n24 VN.n23 161.3
R1603 VN.n22 VN.n2 161.3
R1604 VN.n21 VN.n20 161.3
R1605 VN.n19 VN.n3 161.3
R1606 VN.n18 VN.n17 161.3
R1607 VN.n15 VN.n4 161.3
R1608 VN.n14 VN.n13 161.3
R1609 VN.n12 VN.n5 161.3
R1610 VN.n11 VN.n10 161.3
R1611 VN.n9 VN.n6 161.3
R1612 VN.n30 VN.n29 109.186
R1613 VN.n61 VN.n60 109.186
R1614 VN.n7 VN.t3 69.3223
R1615 VN.n39 VN.t5 69.3223
R1616 VN.n8 VN.n7 56.9625
R1617 VN.n40 VN.n39 56.9625
R1618 VN.n14 VN.n5 56.5617
R1619 VN.n46 VN.n37 56.5617
R1620 VN VN.n61 46.5436
R1621 VN.n23 VN.n22 46.3896
R1622 VN.n54 VN.n53 46.3896
R1623 VN.n8 VN.t4 36.5718
R1624 VN.n16 VN.t7 36.5718
R1625 VN.n29 VN.t1 36.5718
R1626 VN.n40 VN.t2 36.5718
R1627 VN.n36 VN.t6 36.5718
R1628 VN.n60 VN.t0 36.5718
R1629 VN.n23 VN.n1 34.7644
R1630 VN.n54 VN.n32 34.7644
R1631 VN.n10 VN.n9 24.5923
R1632 VN.n10 VN.n5 24.5923
R1633 VN.n15 VN.n14 24.5923
R1634 VN.n17 VN.n15 24.5923
R1635 VN.n21 VN.n3 24.5923
R1636 VN.n22 VN.n21 24.5923
R1637 VN.n27 VN.n1 24.5923
R1638 VN.n28 VN.n27 24.5923
R1639 VN.n42 VN.n37 24.5923
R1640 VN.n42 VN.n41 24.5923
R1641 VN.n53 VN.n52 24.5923
R1642 VN.n52 VN.n34 24.5923
R1643 VN.n48 VN.n47 24.5923
R1644 VN.n47 VN.n46 24.5923
R1645 VN.n59 VN.n58 24.5923
R1646 VN.n58 VN.n32 24.5923
R1647 VN.n9 VN.n8 16.9689
R1648 VN.n17 VN.n16 16.9689
R1649 VN.n41 VN.n40 16.9689
R1650 VN.n48 VN.n36 16.9689
R1651 VN.n16 VN.n3 7.62397
R1652 VN.n36 VN.n34 7.62397
R1653 VN.n39 VN.n38 5.10887
R1654 VN.n7 VN.n6 5.10887
R1655 VN.n29 VN.n28 1.72193
R1656 VN.n60 VN.n59 1.72193
R1657 VN.n61 VN.n31 0.278335
R1658 VN.n30 VN.n0 0.278335
R1659 VN.n57 VN.n31 0.189894
R1660 VN.n57 VN.n56 0.189894
R1661 VN.n56 VN.n55 0.189894
R1662 VN.n55 VN.n33 0.189894
R1663 VN.n51 VN.n33 0.189894
R1664 VN.n51 VN.n50 0.189894
R1665 VN.n50 VN.n49 0.189894
R1666 VN.n49 VN.n35 0.189894
R1667 VN.n45 VN.n35 0.189894
R1668 VN.n45 VN.n44 0.189894
R1669 VN.n44 VN.n43 0.189894
R1670 VN.n43 VN.n38 0.189894
R1671 VN.n11 VN.n6 0.189894
R1672 VN.n12 VN.n11 0.189894
R1673 VN.n13 VN.n12 0.189894
R1674 VN.n13 VN.n4 0.189894
R1675 VN.n18 VN.n4 0.189894
R1676 VN.n19 VN.n18 0.189894
R1677 VN.n20 VN.n19 0.189894
R1678 VN.n20 VN.n2 0.189894
R1679 VN.n24 VN.n2 0.189894
R1680 VN.n25 VN.n24 0.189894
R1681 VN.n26 VN.n25 0.189894
R1682 VN.n26 VN.n0 0.189894
R1683 VN VN.n30 0.153485
R1684 VDD2.n2 VDD2.n1 75.953
R1685 VDD2.n2 VDD2.n0 75.953
R1686 VDD2 VDD2.n5 75.9503
R1687 VDD2.n4 VDD2.n3 74.6336
R1688 VDD2.n4 VDD2.n2 39.8317
R1689 VDD2.n5 VDD2.t5 4.56271
R1690 VDD2.n5 VDD2.t2 4.56271
R1691 VDD2.n3 VDD2.t7 4.56271
R1692 VDD2.n3 VDD2.t1 4.56271
R1693 VDD2.n1 VDD2.t0 4.56271
R1694 VDD2.n1 VDD2.t6 4.56271
R1695 VDD2.n0 VDD2.t4 4.56271
R1696 VDD2.n0 VDD2.t3 4.56271
R1697 VDD2 VDD2.n4 1.43369
C0 VN VTAIL 4.53738f
C1 VTAIL VDD2 5.75169f
C2 VN VDD1 0.156369f
C3 VDD1 VDD2 1.91088f
C4 VTAIL VP 4.55149f
C5 VP VDD1 3.89388f
C6 VN VDD2 3.50039f
C7 VN VP 6.56144f
C8 VP VDD2 0.552068f
C9 VTAIL VDD1 5.695529f
C10 VDD2 B 4.983034f
C11 VDD1 B 5.454711f
C12 VTAIL B 5.647181f
C13 VN B 15.74533f
C14 VP B 14.33454f
C15 VDD2.t4 B 0.083296f
C16 VDD2.t3 B 0.083296f
C17 VDD2.n0 B 0.67249f
C18 VDD2.t0 B 0.083296f
C19 VDD2.t6 B 0.083296f
C20 VDD2.n1 B 0.67249f
C21 VDD2.n2 B 2.85848f
C22 VDD2.t7 B 0.083296f
C23 VDD2.t1 B 0.083296f
C24 VDD2.n3 B 0.663464f
C25 VDD2.n4 B 2.36908f
C26 VDD2.t5 B 0.083296f
C27 VDD2.t2 B 0.083296f
C28 VDD2.n5 B 0.672458f
C29 VN.n0 B 0.033095f
C30 VN.t1 B 0.806172f
C31 VN.n1 B 0.050453f
C32 VN.n2 B 0.025104f
C33 VN.n3 B 0.030695f
C34 VN.n4 B 0.025104f
C35 VN.n5 B 0.036492f
C36 VN.n6 B 0.265092f
C37 VN.t4 B 0.806172f
C38 VN.t3 B 1.03401f
C39 VN.n7 B 0.376798f
C40 VN.n8 B 0.395859f
C41 VN.n9 B 0.039428f
C42 VN.n10 B 0.046553f
C43 VN.n11 B 0.025104f
C44 VN.n12 B 0.025104f
C45 VN.n13 B 0.025104f
C46 VN.n14 B 0.036492f
C47 VN.n15 B 0.046553f
C48 VN.t7 B 0.806172f
C49 VN.n16 B 0.314062f
C50 VN.n17 B 0.039428f
C51 VN.n18 B 0.025104f
C52 VN.n19 B 0.025104f
C53 VN.n20 B 0.025104f
C54 VN.n21 B 0.046553f
C55 VN.n22 B 0.047632f
C56 VN.n23 B 0.021452f
C57 VN.n24 B 0.025104f
C58 VN.n25 B 0.025104f
C59 VN.n26 B 0.025104f
C60 VN.n27 B 0.046553f
C61 VN.n28 B 0.025179f
C62 VN.n29 B 0.395082f
C63 VN.n30 B 0.048015f
C64 VN.n31 B 0.033095f
C65 VN.t0 B 0.806172f
C66 VN.n32 B 0.050453f
C67 VN.n33 B 0.025104f
C68 VN.n34 B 0.030695f
C69 VN.n35 B 0.025104f
C70 VN.t6 B 0.806172f
C71 VN.n36 B 0.314062f
C72 VN.n37 B 0.036492f
C73 VN.n38 B 0.265092f
C74 VN.t2 B 0.806172f
C75 VN.t5 B 1.03401f
C76 VN.n39 B 0.376798f
C77 VN.n40 B 0.395859f
C78 VN.n41 B 0.039428f
C79 VN.n42 B 0.046553f
C80 VN.n43 B 0.025104f
C81 VN.n44 B 0.025104f
C82 VN.n45 B 0.025104f
C83 VN.n46 B 0.036492f
C84 VN.n47 B 0.046553f
C85 VN.n48 B 0.039428f
C86 VN.n49 B 0.025104f
C87 VN.n50 B 0.025104f
C88 VN.n51 B 0.025104f
C89 VN.n52 B 0.046553f
C90 VN.n53 B 0.047632f
C91 VN.n54 B 0.021452f
C92 VN.n55 B 0.025104f
C93 VN.n56 B 0.025104f
C94 VN.n57 B 0.025104f
C95 VN.n58 B 0.046553f
C96 VN.n59 B 0.025179f
C97 VN.n60 B 0.395082f
C98 VN.n61 B 1.26412f
C99 VTAIL.t14 B 0.088988f
C100 VTAIL.t1 B 0.088988f
C101 VTAIL.n0 B 0.651527f
C102 VTAIL.n1 B 0.460751f
C103 VTAIL.t3 B 0.83546f
C104 VTAIL.n2 B 0.553931f
C105 VTAIL.t6 B 0.83546f
C106 VTAIL.n3 B 0.553931f
C107 VTAIL.t10 B 0.088988f
C108 VTAIL.t5 B 0.088988f
C109 VTAIL.n4 B 0.651527f
C110 VTAIL.n5 B 0.685807f
C111 VTAIL.t11 B 0.83546f
C112 VTAIL.n6 B 1.40984f
C113 VTAIL.t15 B 0.835463f
C114 VTAIL.n7 B 1.40984f
C115 VTAIL.t2 B 0.088988f
C116 VTAIL.t0 B 0.088988f
C117 VTAIL.n8 B 0.651531f
C118 VTAIL.n9 B 0.685804f
C119 VTAIL.t12 B 0.835463f
C120 VTAIL.n10 B 0.553927f
C121 VTAIL.t4 B 0.835463f
C122 VTAIL.n11 B 0.553927f
C123 VTAIL.t7 B 0.088988f
C124 VTAIL.t8 B 0.088988f
C125 VTAIL.n12 B 0.651531f
C126 VTAIL.n13 B 0.685804f
C127 VTAIL.t9 B 0.83546f
C128 VTAIL.n14 B 1.40984f
C129 VTAIL.t13 B 0.83546f
C130 VTAIL.n15 B 1.40497f
C131 VDD1.t4 B 0.085161f
C132 VDD1.t7 B 0.085161f
C133 VDD1.n0 B 0.688495f
C134 VDD1.t3 B 0.085161f
C135 VDD1.t6 B 0.085161f
C136 VDD1.n1 B 0.687551f
C137 VDD1.t1 B 0.085161f
C138 VDD1.t2 B 0.085161f
C139 VDD1.n2 B 0.687551f
C140 VDD1.n3 B 2.97427f
C141 VDD1.t0 B 0.085161f
C142 VDD1.t5 B 0.085161f
C143 VDD1.n4 B 0.67832f
C144 VDD1.n5 B 2.45277f
C145 VP.n0 B 0.034311f
C146 VP.t5 B 0.8358f
C147 VP.n1 B 0.052307f
C148 VP.n2 B 0.026026f
C149 VP.n3 B 0.031823f
C150 VP.n4 B 0.026026f
C151 VP.n5 B 0.037833f
C152 VP.n6 B 0.026026f
C153 VP.t1 B 0.8358f
C154 VP.n7 B 0.048263f
C155 VP.n8 B 0.026026f
C156 VP.n9 B 0.048263f
C157 VP.n10 B 0.034311f
C158 VP.t2 B 0.8358f
C159 VP.n11 B 0.052307f
C160 VP.n12 B 0.026026f
C161 VP.n13 B 0.031823f
C162 VP.n14 B 0.026026f
C163 VP.n15 B 0.037833f
C164 VP.n16 B 0.274835f
C165 VP.t4 B 0.8358f
C166 VP.t7 B 1.07202f
C167 VP.n17 B 0.390647f
C168 VP.n18 B 0.410408f
C169 VP.n19 B 0.040877f
C170 VP.n20 B 0.048263f
C171 VP.n21 B 0.026026f
C172 VP.n22 B 0.026026f
C173 VP.n23 B 0.026026f
C174 VP.n24 B 0.037833f
C175 VP.n25 B 0.048263f
C176 VP.t3 B 0.8358f
C177 VP.n26 B 0.325604f
C178 VP.n27 B 0.040877f
C179 VP.n28 B 0.026026f
C180 VP.n29 B 0.026026f
C181 VP.n30 B 0.026026f
C182 VP.n31 B 0.048263f
C183 VP.n32 B 0.049383f
C184 VP.n33 B 0.02224f
C185 VP.n34 B 0.026026f
C186 VP.n35 B 0.026026f
C187 VP.n36 B 0.026026f
C188 VP.n37 B 0.048263f
C189 VP.n38 B 0.026105f
C190 VP.n39 B 0.409602f
C191 VP.n40 B 1.29641f
C192 VP.n41 B 1.31669f
C193 VP.t0 B 0.8358f
C194 VP.n42 B 0.409602f
C195 VP.n43 B 0.026105f
C196 VP.n44 B 0.034311f
C197 VP.n45 B 0.026026f
C198 VP.n46 B 0.026026f
C199 VP.n47 B 0.052307f
C200 VP.n48 B 0.02224f
C201 VP.n49 B 0.049383f
C202 VP.n50 B 0.026026f
C203 VP.n51 B 0.026026f
C204 VP.n52 B 0.026026f
C205 VP.n53 B 0.031823f
C206 VP.n54 B 0.325604f
C207 VP.n55 B 0.040877f
C208 VP.n56 B 0.048263f
C209 VP.n57 B 0.026026f
C210 VP.n58 B 0.026026f
C211 VP.n59 B 0.026026f
C212 VP.n60 B 0.037833f
C213 VP.n61 B 0.048263f
C214 VP.t6 B 0.8358f
C215 VP.n62 B 0.325604f
C216 VP.n63 B 0.040877f
C217 VP.n64 B 0.026026f
C218 VP.n65 B 0.026026f
C219 VP.n66 B 0.026026f
C220 VP.n67 B 0.048263f
C221 VP.n68 B 0.049383f
C222 VP.n69 B 0.02224f
C223 VP.n70 B 0.026026f
C224 VP.n71 B 0.026026f
C225 VP.n72 B 0.026026f
C226 VP.n73 B 0.048263f
C227 VP.n74 B 0.026105f
C228 VP.n75 B 0.409602f
C229 VP.n76 B 0.04978f
.ends

