* NGSPICE file created from diff_pair_sample_0154.ext - technology: sky130A

.subckt diff_pair_sample_0154 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t1 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=3.26865 pd=20.14 as=3.26865 ps=20.14 w=19.81 l=1.22
X1 VTAIL.t7 VN.t0 VDD2.t9 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=3.26865 pd=20.14 as=3.26865 ps=20.14 w=19.81 l=1.22
X2 B.t11 B.t9 B.t10 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=7.7259 pd=40.4 as=0 ps=0 w=19.81 l=1.22
X3 VTAIL.t18 VP.t1 VDD1.t0 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=3.26865 pd=20.14 as=3.26865 ps=20.14 w=19.81 l=1.22
X4 VDD2.t8 VN.t1 VTAIL.t1 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=3.26865 pd=20.14 as=3.26865 ps=20.14 w=19.81 l=1.22
X5 VTAIL.t9 VN.t2 VDD2.t7 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=3.26865 pd=20.14 as=3.26865 ps=20.14 w=19.81 l=1.22
X6 B.t8 B.t6 B.t7 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=7.7259 pd=40.4 as=0 ps=0 w=19.81 l=1.22
X7 VTAIL.t17 VP.t2 VDD1.t5 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=3.26865 pd=20.14 as=3.26865 ps=20.14 w=19.81 l=1.22
X8 B.t5 B.t3 B.t4 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=7.7259 pd=40.4 as=0 ps=0 w=19.81 l=1.22
X9 VTAIL.t16 VP.t3 VDD1.t4 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=3.26865 pd=20.14 as=3.26865 ps=20.14 w=19.81 l=1.22
X10 VDD1.t3 VP.t4 VTAIL.t15 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=3.26865 pd=20.14 as=3.26865 ps=20.14 w=19.81 l=1.22
X11 VTAIL.t0 VN.t3 VDD2.t6 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=3.26865 pd=20.14 as=3.26865 ps=20.14 w=19.81 l=1.22
X12 VDD1.t2 VP.t5 VTAIL.t14 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=7.7259 pd=40.4 as=3.26865 ps=20.14 w=19.81 l=1.22
X13 VDD2.t5 VN.t4 VTAIL.t3 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=3.26865 pd=20.14 as=7.7259 ps=40.4 w=19.81 l=1.22
X14 VTAIL.t4 VN.t5 VDD2.t4 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=3.26865 pd=20.14 as=3.26865 ps=20.14 w=19.81 l=1.22
X15 VDD1.t7 VP.t6 VTAIL.t13 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=7.7259 pd=40.4 as=3.26865 ps=20.14 w=19.81 l=1.22
X16 B.t2 B.t0 B.t1 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=7.7259 pd=40.4 as=0 ps=0 w=19.81 l=1.22
X17 VDD2.t3 VN.t6 VTAIL.t8 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=7.7259 pd=40.4 as=3.26865 ps=20.14 w=19.81 l=1.22
X18 VDD1.t6 VP.t7 VTAIL.t12 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=3.26865 pd=20.14 as=3.26865 ps=20.14 w=19.81 l=1.22
X19 VDD1.t9 VP.t8 VTAIL.t11 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=3.26865 pd=20.14 as=7.7259 ps=40.4 w=19.81 l=1.22
X20 VDD2.t2 VN.t7 VTAIL.t2 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=7.7259 pd=40.4 as=3.26865 ps=20.14 w=19.81 l=1.22
X21 VDD2.t1 VN.t8 VTAIL.t5 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=3.26865 pd=20.14 as=7.7259 ps=40.4 w=19.81 l=1.22
X22 VDD2.t0 VN.t9 VTAIL.t6 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=3.26865 pd=20.14 as=3.26865 ps=20.14 w=19.81 l=1.22
X23 VDD1.t8 VP.t9 VTAIL.t10 w_n2830_n4930# sky130_fd_pr__pfet_01v8 ad=3.26865 pd=20.14 as=7.7259 ps=40.4 w=19.81 l=1.22
R0 VP.n13 VP.t5 443.615
R1 VP.n30 VP.t6 423.726
R2 VP.n47 VP.t8 423.726
R3 VP.n27 VP.t9 423.726
R4 VP.n5 VP.t0 391.329
R5 VP.n3 VP.t7 391.329
R6 VP.n1 VP.t2 391.329
R7 VP.n8 VP.t1 391.329
R8 VP.n10 VP.t4 391.329
R9 VP.n12 VP.t3 391.329
R10 VP.n15 VP.n14 161.3
R11 VP.n16 VP.n11 161.3
R12 VP.n18 VP.n17 161.3
R13 VP.n20 VP.n19 161.3
R14 VP.n21 VP.n9 161.3
R15 VP.n23 VP.n22 161.3
R16 VP.n25 VP.n24 161.3
R17 VP.n26 VP.n7 161.3
R18 VP.n46 VP.n0 161.3
R19 VP.n45 VP.n44 161.3
R20 VP.n43 VP.n42 161.3
R21 VP.n41 VP.n2 161.3
R22 VP.n40 VP.n39 161.3
R23 VP.n38 VP.n37 161.3
R24 VP.n36 VP.n4 161.3
R25 VP.n35 VP.n34 161.3
R26 VP.n33 VP.n32 161.3
R27 VP.n31 VP.n6 161.3
R28 VP.n28 VP.n27 80.6037
R29 VP.n48 VP.n47 80.6037
R30 VP.n30 VP.n29 80.6037
R31 VP.n29 VP.n28 51.687
R32 VP.n36 VP.n35 42.9216
R33 VP.n42 VP.n41 42.9216
R34 VP.n22 VP.n21 42.9216
R35 VP.n16 VP.n15 42.9216
R36 VP.n13 VP.n12 42.7694
R37 VP.n37 VP.n36 38.0652
R38 VP.n41 VP.n40 38.0652
R39 VP.n21 VP.n20 38.0652
R40 VP.n17 VP.n16 38.0652
R41 VP.n31 VP.n30 35.055
R42 VP.n47 VP.n46 35.055
R43 VP.n27 VP.n26 35.055
R44 VP.n32 VP.n31 33.2089
R45 VP.n46 VP.n45 33.2089
R46 VP.n26 VP.n25 33.2089
R47 VP.n14 VP.n13 29.263
R48 VP.n35 VP.n5 14.6807
R49 VP.n42 VP.n1 14.6807
R50 VP.n22 VP.n8 14.6807
R51 VP.n15 VP.n12 14.6807
R52 VP.n37 VP.n3 12.234
R53 VP.n40 VP.n3 12.234
R54 VP.n17 VP.n10 12.234
R55 VP.n20 VP.n10 12.234
R56 VP.n32 VP.n5 9.7873
R57 VP.n45 VP.n1 9.7873
R58 VP.n25 VP.n8 9.7873
R59 VP.n28 VP.n7 0.285035
R60 VP.n29 VP.n6 0.285035
R61 VP.n48 VP.n0 0.285035
R62 VP.n14 VP.n11 0.189894
R63 VP.n18 VP.n11 0.189894
R64 VP.n19 VP.n18 0.189894
R65 VP.n19 VP.n9 0.189894
R66 VP.n23 VP.n9 0.189894
R67 VP.n24 VP.n23 0.189894
R68 VP.n24 VP.n7 0.189894
R69 VP.n33 VP.n6 0.189894
R70 VP.n34 VP.n33 0.189894
R71 VP.n34 VP.n4 0.189894
R72 VP.n38 VP.n4 0.189894
R73 VP.n39 VP.n38 0.189894
R74 VP.n39 VP.n2 0.189894
R75 VP.n43 VP.n2 0.189894
R76 VP.n44 VP.n43 0.189894
R77 VP.n44 VP.n0 0.189894
R78 VP VP.n48 0.146778
R79 VDD1.n1 VDD1.t2 73.2204
R80 VDD1.n3 VDD1.t7 73.2202
R81 VDD1.n5 VDD1.n4 71.19
R82 VDD1.n1 VDD1.n0 70.2434
R83 VDD1.n7 VDD1.n6 70.2433
R84 VDD1.n3 VDD1.n2 70.2432
R85 VDD1.n7 VDD1.n5 48.391
R86 VDD1.n6 VDD1.t0 1.64134
R87 VDD1.n6 VDD1.t8 1.64134
R88 VDD1.n0 VDD1.t4 1.64134
R89 VDD1.n0 VDD1.t3 1.64134
R90 VDD1.n4 VDD1.t5 1.64134
R91 VDD1.n4 VDD1.t9 1.64134
R92 VDD1.n2 VDD1.t1 1.64134
R93 VDD1.n2 VDD1.t6 1.64134
R94 VDD1 VDD1.n7 0.944465
R95 VDD1 VDD1.n1 0.392741
R96 VDD1.n5 VDD1.n3 0.279206
R97 VTAIL.n11 VTAIL.t3 55.2055
R98 VTAIL.n17 VTAIL.t5 55.2053
R99 VTAIL.n2 VTAIL.t11 55.2053
R100 VTAIL.n16 VTAIL.t10 55.2053
R101 VTAIL.n15 VTAIL.n14 53.5646
R102 VTAIL.n13 VTAIL.n12 53.5646
R103 VTAIL.n10 VTAIL.n9 53.5646
R104 VTAIL.n8 VTAIL.n7 53.5646
R105 VTAIL.n19 VTAIL.n18 53.5644
R106 VTAIL.n1 VTAIL.n0 53.5644
R107 VTAIL.n4 VTAIL.n3 53.5644
R108 VTAIL.n6 VTAIL.n5 53.5644
R109 VTAIL.n8 VTAIL.n6 32.1169
R110 VTAIL.n17 VTAIL.n16 30.7807
R111 VTAIL.n18 VTAIL.t6 1.64134
R112 VTAIL.n18 VTAIL.t4 1.64134
R113 VTAIL.n0 VTAIL.t8 1.64134
R114 VTAIL.n0 VTAIL.t9 1.64134
R115 VTAIL.n3 VTAIL.t12 1.64134
R116 VTAIL.n3 VTAIL.t17 1.64134
R117 VTAIL.n5 VTAIL.t13 1.64134
R118 VTAIL.n5 VTAIL.t19 1.64134
R119 VTAIL.n14 VTAIL.t15 1.64134
R120 VTAIL.n14 VTAIL.t18 1.64134
R121 VTAIL.n12 VTAIL.t14 1.64134
R122 VTAIL.n12 VTAIL.t16 1.64134
R123 VTAIL.n9 VTAIL.t1 1.64134
R124 VTAIL.n9 VTAIL.t0 1.64134
R125 VTAIL.n7 VTAIL.t2 1.64134
R126 VTAIL.n7 VTAIL.t7 1.64134
R127 VTAIL.n10 VTAIL.n8 1.33671
R128 VTAIL.n11 VTAIL.n10 1.33671
R129 VTAIL.n15 VTAIL.n13 1.33671
R130 VTAIL.n16 VTAIL.n15 1.33671
R131 VTAIL.n6 VTAIL.n4 1.33671
R132 VTAIL.n4 VTAIL.n2 1.33671
R133 VTAIL.n19 VTAIL.n17 1.33671
R134 VTAIL.n13 VTAIL.n11 1.13843
R135 VTAIL.n2 VTAIL.n1 1.13843
R136 VTAIL VTAIL.n1 1.06084
R137 VTAIL VTAIL.n19 0.276362
R138 VN.n6 VN.t6 443.615
R139 VN.n28 VN.t4 443.615
R140 VN.n20 VN.t8 423.726
R141 VN.n42 VN.t7 423.726
R142 VN.n5 VN.t2 391.329
R143 VN.n3 VN.t9 391.329
R144 VN.n1 VN.t5 391.329
R145 VN.n27 VN.t3 391.329
R146 VN.n25 VN.t1 391.329
R147 VN.n23 VN.t0 391.329
R148 VN.n41 VN.n22 161.3
R149 VN.n40 VN.n39 161.3
R150 VN.n38 VN.n37 161.3
R151 VN.n36 VN.n24 161.3
R152 VN.n35 VN.n34 161.3
R153 VN.n33 VN.n32 161.3
R154 VN.n31 VN.n26 161.3
R155 VN.n30 VN.n29 161.3
R156 VN.n19 VN.n0 161.3
R157 VN.n18 VN.n17 161.3
R158 VN.n16 VN.n15 161.3
R159 VN.n14 VN.n2 161.3
R160 VN.n13 VN.n12 161.3
R161 VN.n11 VN.n10 161.3
R162 VN.n9 VN.n4 161.3
R163 VN.n8 VN.n7 161.3
R164 VN.n43 VN.n42 80.6037
R165 VN.n21 VN.n20 80.6037
R166 VN VN.n43 51.9725
R167 VN.n9 VN.n8 42.9216
R168 VN.n15 VN.n14 42.9216
R169 VN.n31 VN.n30 42.9216
R170 VN.n37 VN.n36 42.9216
R171 VN.n6 VN.n5 42.7694
R172 VN.n28 VN.n27 42.7694
R173 VN.n10 VN.n9 38.0652
R174 VN.n14 VN.n13 38.0652
R175 VN.n32 VN.n31 38.0652
R176 VN.n36 VN.n35 38.0652
R177 VN.n20 VN.n19 35.055
R178 VN.n42 VN.n41 35.055
R179 VN.n19 VN.n18 33.2089
R180 VN.n41 VN.n40 33.2089
R181 VN.n29 VN.n28 29.263
R182 VN.n7 VN.n6 29.263
R183 VN.n8 VN.n5 14.6807
R184 VN.n15 VN.n1 14.6807
R185 VN.n30 VN.n27 14.6807
R186 VN.n37 VN.n23 14.6807
R187 VN.n10 VN.n3 12.234
R188 VN.n13 VN.n3 12.234
R189 VN.n35 VN.n25 12.234
R190 VN.n32 VN.n25 12.234
R191 VN.n18 VN.n1 9.7873
R192 VN.n40 VN.n23 9.7873
R193 VN.n43 VN.n22 0.285035
R194 VN.n21 VN.n0 0.285035
R195 VN.n39 VN.n22 0.189894
R196 VN.n39 VN.n38 0.189894
R197 VN.n38 VN.n24 0.189894
R198 VN.n34 VN.n24 0.189894
R199 VN.n34 VN.n33 0.189894
R200 VN.n33 VN.n26 0.189894
R201 VN.n29 VN.n26 0.189894
R202 VN.n7 VN.n4 0.189894
R203 VN.n11 VN.n4 0.189894
R204 VN.n12 VN.n11 0.189894
R205 VN.n12 VN.n2 0.189894
R206 VN.n16 VN.n2 0.189894
R207 VN.n17 VN.n16 0.189894
R208 VN.n17 VN.n0 0.189894
R209 VN VN.n21 0.146778
R210 VDD2.n1 VDD2.t3 73.2202
R211 VDD2.n4 VDD2.t2 71.8842
R212 VDD2.n3 VDD2.n2 71.19
R213 VDD2 VDD2.n7 71.1872
R214 VDD2.n6 VDD2.n5 70.2434
R215 VDD2.n1 VDD2.n0 70.2432
R216 VDD2.n4 VDD2.n3 47.1399
R217 VDD2.n7 VDD2.t6 1.64134
R218 VDD2.n7 VDD2.t5 1.64134
R219 VDD2.n5 VDD2.t9 1.64134
R220 VDD2.n5 VDD2.t8 1.64134
R221 VDD2.n2 VDD2.t4 1.64134
R222 VDD2.n2 VDD2.t1 1.64134
R223 VDD2.n0 VDD2.t7 1.64134
R224 VDD2.n0 VDD2.t0 1.64134
R225 VDD2.n6 VDD2.n4 1.33671
R226 VDD2 VDD2.n6 0.392741
R227 VDD2.n3 VDD2.n1 0.279206
R228 B.n170 B.t9 595.548
R229 B.n162 B.t6 595.548
R230 B.n60 B.t3 595.548
R231 B.n52 B.t0 595.548
R232 B.n481 B.n480 585
R233 B.n479 B.n130 585
R234 B.n478 B.n477 585
R235 B.n476 B.n131 585
R236 B.n475 B.n474 585
R237 B.n473 B.n132 585
R238 B.n472 B.n471 585
R239 B.n470 B.n133 585
R240 B.n469 B.n468 585
R241 B.n467 B.n134 585
R242 B.n466 B.n465 585
R243 B.n464 B.n135 585
R244 B.n463 B.n462 585
R245 B.n461 B.n136 585
R246 B.n460 B.n459 585
R247 B.n458 B.n137 585
R248 B.n457 B.n456 585
R249 B.n455 B.n138 585
R250 B.n454 B.n453 585
R251 B.n452 B.n139 585
R252 B.n451 B.n450 585
R253 B.n449 B.n140 585
R254 B.n448 B.n447 585
R255 B.n446 B.n141 585
R256 B.n445 B.n444 585
R257 B.n443 B.n142 585
R258 B.n442 B.n441 585
R259 B.n440 B.n143 585
R260 B.n439 B.n438 585
R261 B.n437 B.n144 585
R262 B.n436 B.n435 585
R263 B.n434 B.n145 585
R264 B.n433 B.n432 585
R265 B.n431 B.n146 585
R266 B.n430 B.n429 585
R267 B.n428 B.n147 585
R268 B.n427 B.n426 585
R269 B.n425 B.n148 585
R270 B.n424 B.n423 585
R271 B.n422 B.n149 585
R272 B.n421 B.n420 585
R273 B.n419 B.n150 585
R274 B.n418 B.n417 585
R275 B.n416 B.n151 585
R276 B.n415 B.n414 585
R277 B.n413 B.n152 585
R278 B.n412 B.n411 585
R279 B.n410 B.n153 585
R280 B.n409 B.n408 585
R281 B.n407 B.n154 585
R282 B.n406 B.n405 585
R283 B.n404 B.n155 585
R284 B.n403 B.n402 585
R285 B.n401 B.n156 585
R286 B.n400 B.n399 585
R287 B.n398 B.n157 585
R288 B.n397 B.n396 585
R289 B.n395 B.n158 585
R290 B.n394 B.n393 585
R291 B.n392 B.n159 585
R292 B.n391 B.n390 585
R293 B.n389 B.n160 585
R294 B.n388 B.n387 585
R295 B.n386 B.n161 585
R296 B.n385 B.n384 585
R297 B.n383 B.n382 585
R298 B.n381 B.n165 585
R299 B.n380 B.n379 585
R300 B.n378 B.n166 585
R301 B.n377 B.n376 585
R302 B.n375 B.n167 585
R303 B.n374 B.n373 585
R304 B.n372 B.n168 585
R305 B.n371 B.n370 585
R306 B.n368 B.n169 585
R307 B.n367 B.n366 585
R308 B.n365 B.n172 585
R309 B.n364 B.n363 585
R310 B.n362 B.n173 585
R311 B.n361 B.n360 585
R312 B.n359 B.n174 585
R313 B.n358 B.n357 585
R314 B.n356 B.n175 585
R315 B.n355 B.n354 585
R316 B.n353 B.n176 585
R317 B.n352 B.n351 585
R318 B.n350 B.n177 585
R319 B.n349 B.n348 585
R320 B.n347 B.n178 585
R321 B.n346 B.n345 585
R322 B.n344 B.n179 585
R323 B.n343 B.n342 585
R324 B.n341 B.n180 585
R325 B.n340 B.n339 585
R326 B.n338 B.n181 585
R327 B.n337 B.n336 585
R328 B.n335 B.n182 585
R329 B.n334 B.n333 585
R330 B.n332 B.n183 585
R331 B.n331 B.n330 585
R332 B.n329 B.n184 585
R333 B.n328 B.n327 585
R334 B.n326 B.n185 585
R335 B.n325 B.n324 585
R336 B.n323 B.n186 585
R337 B.n322 B.n321 585
R338 B.n320 B.n187 585
R339 B.n319 B.n318 585
R340 B.n317 B.n188 585
R341 B.n316 B.n315 585
R342 B.n314 B.n189 585
R343 B.n313 B.n312 585
R344 B.n311 B.n190 585
R345 B.n310 B.n309 585
R346 B.n308 B.n191 585
R347 B.n307 B.n306 585
R348 B.n305 B.n192 585
R349 B.n304 B.n303 585
R350 B.n302 B.n193 585
R351 B.n301 B.n300 585
R352 B.n299 B.n194 585
R353 B.n298 B.n297 585
R354 B.n296 B.n195 585
R355 B.n295 B.n294 585
R356 B.n293 B.n196 585
R357 B.n292 B.n291 585
R358 B.n290 B.n197 585
R359 B.n289 B.n288 585
R360 B.n287 B.n198 585
R361 B.n286 B.n285 585
R362 B.n284 B.n199 585
R363 B.n283 B.n282 585
R364 B.n281 B.n200 585
R365 B.n280 B.n279 585
R366 B.n278 B.n201 585
R367 B.n277 B.n276 585
R368 B.n275 B.n202 585
R369 B.n274 B.n273 585
R370 B.n272 B.n203 585
R371 B.n482 B.n129 585
R372 B.n484 B.n483 585
R373 B.n485 B.n128 585
R374 B.n487 B.n486 585
R375 B.n488 B.n127 585
R376 B.n490 B.n489 585
R377 B.n491 B.n126 585
R378 B.n493 B.n492 585
R379 B.n494 B.n125 585
R380 B.n496 B.n495 585
R381 B.n497 B.n124 585
R382 B.n499 B.n498 585
R383 B.n500 B.n123 585
R384 B.n502 B.n501 585
R385 B.n503 B.n122 585
R386 B.n505 B.n504 585
R387 B.n506 B.n121 585
R388 B.n508 B.n507 585
R389 B.n509 B.n120 585
R390 B.n511 B.n510 585
R391 B.n512 B.n119 585
R392 B.n514 B.n513 585
R393 B.n515 B.n118 585
R394 B.n517 B.n516 585
R395 B.n518 B.n117 585
R396 B.n520 B.n519 585
R397 B.n521 B.n116 585
R398 B.n523 B.n522 585
R399 B.n524 B.n115 585
R400 B.n526 B.n525 585
R401 B.n527 B.n114 585
R402 B.n529 B.n528 585
R403 B.n530 B.n113 585
R404 B.n532 B.n531 585
R405 B.n533 B.n112 585
R406 B.n535 B.n534 585
R407 B.n536 B.n111 585
R408 B.n538 B.n537 585
R409 B.n539 B.n110 585
R410 B.n541 B.n540 585
R411 B.n542 B.n109 585
R412 B.n544 B.n543 585
R413 B.n545 B.n108 585
R414 B.n547 B.n546 585
R415 B.n548 B.n107 585
R416 B.n550 B.n549 585
R417 B.n551 B.n106 585
R418 B.n553 B.n552 585
R419 B.n554 B.n105 585
R420 B.n556 B.n555 585
R421 B.n557 B.n104 585
R422 B.n559 B.n558 585
R423 B.n560 B.n103 585
R424 B.n562 B.n561 585
R425 B.n563 B.n102 585
R426 B.n565 B.n564 585
R427 B.n566 B.n101 585
R428 B.n568 B.n567 585
R429 B.n569 B.n100 585
R430 B.n571 B.n570 585
R431 B.n572 B.n99 585
R432 B.n574 B.n573 585
R433 B.n575 B.n98 585
R434 B.n577 B.n576 585
R435 B.n578 B.n97 585
R436 B.n580 B.n579 585
R437 B.n581 B.n96 585
R438 B.n583 B.n582 585
R439 B.n584 B.n95 585
R440 B.n586 B.n585 585
R441 B.n587 B.n94 585
R442 B.n589 B.n588 585
R443 B.n799 B.n798 585
R444 B.n797 B.n20 585
R445 B.n796 B.n795 585
R446 B.n794 B.n21 585
R447 B.n793 B.n792 585
R448 B.n791 B.n22 585
R449 B.n790 B.n789 585
R450 B.n788 B.n23 585
R451 B.n787 B.n786 585
R452 B.n785 B.n24 585
R453 B.n784 B.n783 585
R454 B.n782 B.n25 585
R455 B.n781 B.n780 585
R456 B.n779 B.n26 585
R457 B.n778 B.n777 585
R458 B.n776 B.n27 585
R459 B.n775 B.n774 585
R460 B.n773 B.n28 585
R461 B.n772 B.n771 585
R462 B.n770 B.n29 585
R463 B.n769 B.n768 585
R464 B.n767 B.n30 585
R465 B.n766 B.n765 585
R466 B.n764 B.n31 585
R467 B.n763 B.n762 585
R468 B.n761 B.n32 585
R469 B.n760 B.n759 585
R470 B.n758 B.n33 585
R471 B.n757 B.n756 585
R472 B.n755 B.n34 585
R473 B.n754 B.n753 585
R474 B.n752 B.n35 585
R475 B.n751 B.n750 585
R476 B.n749 B.n36 585
R477 B.n748 B.n747 585
R478 B.n746 B.n37 585
R479 B.n745 B.n744 585
R480 B.n743 B.n38 585
R481 B.n742 B.n741 585
R482 B.n740 B.n39 585
R483 B.n739 B.n738 585
R484 B.n737 B.n40 585
R485 B.n736 B.n735 585
R486 B.n734 B.n41 585
R487 B.n733 B.n732 585
R488 B.n731 B.n42 585
R489 B.n730 B.n729 585
R490 B.n728 B.n43 585
R491 B.n727 B.n726 585
R492 B.n725 B.n44 585
R493 B.n724 B.n723 585
R494 B.n722 B.n45 585
R495 B.n721 B.n720 585
R496 B.n719 B.n46 585
R497 B.n718 B.n717 585
R498 B.n716 B.n47 585
R499 B.n715 B.n714 585
R500 B.n713 B.n48 585
R501 B.n712 B.n711 585
R502 B.n710 B.n49 585
R503 B.n709 B.n708 585
R504 B.n707 B.n50 585
R505 B.n706 B.n705 585
R506 B.n704 B.n51 585
R507 B.n703 B.n702 585
R508 B.n701 B.n700 585
R509 B.n699 B.n55 585
R510 B.n698 B.n697 585
R511 B.n696 B.n56 585
R512 B.n695 B.n694 585
R513 B.n693 B.n57 585
R514 B.n692 B.n691 585
R515 B.n690 B.n58 585
R516 B.n689 B.n688 585
R517 B.n686 B.n59 585
R518 B.n685 B.n684 585
R519 B.n683 B.n62 585
R520 B.n682 B.n681 585
R521 B.n680 B.n63 585
R522 B.n679 B.n678 585
R523 B.n677 B.n64 585
R524 B.n676 B.n675 585
R525 B.n674 B.n65 585
R526 B.n673 B.n672 585
R527 B.n671 B.n66 585
R528 B.n670 B.n669 585
R529 B.n668 B.n67 585
R530 B.n667 B.n666 585
R531 B.n665 B.n68 585
R532 B.n664 B.n663 585
R533 B.n662 B.n69 585
R534 B.n661 B.n660 585
R535 B.n659 B.n70 585
R536 B.n658 B.n657 585
R537 B.n656 B.n71 585
R538 B.n655 B.n654 585
R539 B.n653 B.n72 585
R540 B.n652 B.n651 585
R541 B.n650 B.n73 585
R542 B.n649 B.n648 585
R543 B.n647 B.n74 585
R544 B.n646 B.n645 585
R545 B.n644 B.n75 585
R546 B.n643 B.n642 585
R547 B.n641 B.n76 585
R548 B.n640 B.n639 585
R549 B.n638 B.n77 585
R550 B.n637 B.n636 585
R551 B.n635 B.n78 585
R552 B.n634 B.n633 585
R553 B.n632 B.n79 585
R554 B.n631 B.n630 585
R555 B.n629 B.n80 585
R556 B.n628 B.n627 585
R557 B.n626 B.n81 585
R558 B.n625 B.n624 585
R559 B.n623 B.n82 585
R560 B.n622 B.n621 585
R561 B.n620 B.n83 585
R562 B.n619 B.n618 585
R563 B.n617 B.n84 585
R564 B.n616 B.n615 585
R565 B.n614 B.n85 585
R566 B.n613 B.n612 585
R567 B.n611 B.n86 585
R568 B.n610 B.n609 585
R569 B.n608 B.n87 585
R570 B.n607 B.n606 585
R571 B.n605 B.n88 585
R572 B.n604 B.n603 585
R573 B.n602 B.n89 585
R574 B.n601 B.n600 585
R575 B.n599 B.n90 585
R576 B.n598 B.n597 585
R577 B.n596 B.n91 585
R578 B.n595 B.n594 585
R579 B.n593 B.n92 585
R580 B.n592 B.n591 585
R581 B.n590 B.n93 585
R582 B.n800 B.n19 585
R583 B.n802 B.n801 585
R584 B.n803 B.n18 585
R585 B.n805 B.n804 585
R586 B.n806 B.n17 585
R587 B.n808 B.n807 585
R588 B.n809 B.n16 585
R589 B.n811 B.n810 585
R590 B.n812 B.n15 585
R591 B.n814 B.n813 585
R592 B.n815 B.n14 585
R593 B.n817 B.n816 585
R594 B.n818 B.n13 585
R595 B.n820 B.n819 585
R596 B.n821 B.n12 585
R597 B.n823 B.n822 585
R598 B.n824 B.n11 585
R599 B.n826 B.n825 585
R600 B.n827 B.n10 585
R601 B.n829 B.n828 585
R602 B.n830 B.n9 585
R603 B.n832 B.n831 585
R604 B.n833 B.n8 585
R605 B.n835 B.n834 585
R606 B.n836 B.n7 585
R607 B.n838 B.n837 585
R608 B.n839 B.n6 585
R609 B.n841 B.n840 585
R610 B.n842 B.n5 585
R611 B.n844 B.n843 585
R612 B.n845 B.n4 585
R613 B.n847 B.n846 585
R614 B.n848 B.n3 585
R615 B.n850 B.n849 585
R616 B.n851 B.n0 585
R617 B.n2 B.n1 585
R618 B.n221 B.n220 585
R619 B.n223 B.n222 585
R620 B.n224 B.n219 585
R621 B.n226 B.n225 585
R622 B.n227 B.n218 585
R623 B.n229 B.n228 585
R624 B.n230 B.n217 585
R625 B.n232 B.n231 585
R626 B.n233 B.n216 585
R627 B.n235 B.n234 585
R628 B.n236 B.n215 585
R629 B.n238 B.n237 585
R630 B.n239 B.n214 585
R631 B.n241 B.n240 585
R632 B.n242 B.n213 585
R633 B.n244 B.n243 585
R634 B.n245 B.n212 585
R635 B.n247 B.n246 585
R636 B.n248 B.n211 585
R637 B.n250 B.n249 585
R638 B.n251 B.n210 585
R639 B.n253 B.n252 585
R640 B.n254 B.n209 585
R641 B.n256 B.n255 585
R642 B.n257 B.n208 585
R643 B.n259 B.n258 585
R644 B.n260 B.n207 585
R645 B.n262 B.n261 585
R646 B.n263 B.n206 585
R647 B.n265 B.n264 585
R648 B.n266 B.n205 585
R649 B.n268 B.n267 585
R650 B.n269 B.n204 585
R651 B.n271 B.n270 585
R652 B.n270 B.n203 473.281
R653 B.n480 B.n129 473.281
R654 B.n588 B.n93 473.281
R655 B.n798 B.n19 473.281
R656 B.n853 B.n852 256.663
R657 B.n852 B.n851 235.042
R658 B.n852 B.n2 235.042
R659 B.n274 B.n203 163.367
R660 B.n275 B.n274 163.367
R661 B.n276 B.n275 163.367
R662 B.n276 B.n201 163.367
R663 B.n280 B.n201 163.367
R664 B.n281 B.n280 163.367
R665 B.n282 B.n281 163.367
R666 B.n282 B.n199 163.367
R667 B.n286 B.n199 163.367
R668 B.n287 B.n286 163.367
R669 B.n288 B.n287 163.367
R670 B.n288 B.n197 163.367
R671 B.n292 B.n197 163.367
R672 B.n293 B.n292 163.367
R673 B.n294 B.n293 163.367
R674 B.n294 B.n195 163.367
R675 B.n298 B.n195 163.367
R676 B.n299 B.n298 163.367
R677 B.n300 B.n299 163.367
R678 B.n300 B.n193 163.367
R679 B.n304 B.n193 163.367
R680 B.n305 B.n304 163.367
R681 B.n306 B.n305 163.367
R682 B.n306 B.n191 163.367
R683 B.n310 B.n191 163.367
R684 B.n311 B.n310 163.367
R685 B.n312 B.n311 163.367
R686 B.n312 B.n189 163.367
R687 B.n316 B.n189 163.367
R688 B.n317 B.n316 163.367
R689 B.n318 B.n317 163.367
R690 B.n318 B.n187 163.367
R691 B.n322 B.n187 163.367
R692 B.n323 B.n322 163.367
R693 B.n324 B.n323 163.367
R694 B.n324 B.n185 163.367
R695 B.n328 B.n185 163.367
R696 B.n329 B.n328 163.367
R697 B.n330 B.n329 163.367
R698 B.n330 B.n183 163.367
R699 B.n334 B.n183 163.367
R700 B.n335 B.n334 163.367
R701 B.n336 B.n335 163.367
R702 B.n336 B.n181 163.367
R703 B.n340 B.n181 163.367
R704 B.n341 B.n340 163.367
R705 B.n342 B.n341 163.367
R706 B.n342 B.n179 163.367
R707 B.n346 B.n179 163.367
R708 B.n347 B.n346 163.367
R709 B.n348 B.n347 163.367
R710 B.n348 B.n177 163.367
R711 B.n352 B.n177 163.367
R712 B.n353 B.n352 163.367
R713 B.n354 B.n353 163.367
R714 B.n354 B.n175 163.367
R715 B.n358 B.n175 163.367
R716 B.n359 B.n358 163.367
R717 B.n360 B.n359 163.367
R718 B.n360 B.n173 163.367
R719 B.n364 B.n173 163.367
R720 B.n365 B.n364 163.367
R721 B.n366 B.n365 163.367
R722 B.n366 B.n169 163.367
R723 B.n371 B.n169 163.367
R724 B.n372 B.n371 163.367
R725 B.n373 B.n372 163.367
R726 B.n373 B.n167 163.367
R727 B.n377 B.n167 163.367
R728 B.n378 B.n377 163.367
R729 B.n379 B.n378 163.367
R730 B.n379 B.n165 163.367
R731 B.n383 B.n165 163.367
R732 B.n384 B.n383 163.367
R733 B.n384 B.n161 163.367
R734 B.n388 B.n161 163.367
R735 B.n389 B.n388 163.367
R736 B.n390 B.n389 163.367
R737 B.n390 B.n159 163.367
R738 B.n394 B.n159 163.367
R739 B.n395 B.n394 163.367
R740 B.n396 B.n395 163.367
R741 B.n396 B.n157 163.367
R742 B.n400 B.n157 163.367
R743 B.n401 B.n400 163.367
R744 B.n402 B.n401 163.367
R745 B.n402 B.n155 163.367
R746 B.n406 B.n155 163.367
R747 B.n407 B.n406 163.367
R748 B.n408 B.n407 163.367
R749 B.n408 B.n153 163.367
R750 B.n412 B.n153 163.367
R751 B.n413 B.n412 163.367
R752 B.n414 B.n413 163.367
R753 B.n414 B.n151 163.367
R754 B.n418 B.n151 163.367
R755 B.n419 B.n418 163.367
R756 B.n420 B.n419 163.367
R757 B.n420 B.n149 163.367
R758 B.n424 B.n149 163.367
R759 B.n425 B.n424 163.367
R760 B.n426 B.n425 163.367
R761 B.n426 B.n147 163.367
R762 B.n430 B.n147 163.367
R763 B.n431 B.n430 163.367
R764 B.n432 B.n431 163.367
R765 B.n432 B.n145 163.367
R766 B.n436 B.n145 163.367
R767 B.n437 B.n436 163.367
R768 B.n438 B.n437 163.367
R769 B.n438 B.n143 163.367
R770 B.n442 B.n143 163.367
R771 B.n443 B.n442 163.367
R772 B.n444 B.n443 163.367
R773 B.n444 B.n141 163.367
R774 B.n448 B.n141 163.367
R775 B.n449 B.n448 163.367
R776 B.n450 B.n449 163.367
R777 B.n450 B.n139 163.367
R778 B.n454 B.n139 163.367
R779 B.n455 B.n454 163.367
R780 B.n456 B.n455 163.367
R781 B.n456 B.n137 163.367
R782 B.n460 B.n137 163.367
R783 B.n461 B.n460 163.367
R784 B.n462 B.n461 163.367
R785 B.n462 B.n135 163.367
R786 B.n466 B.n135 163.367
R787 B.n467 B.n466 163.367
R788 B.n468 B.n467 163.367
R789 B.n468 B.n133 163.367
R790 B.n472 B.n133 163.367
R791 B.n473 B.n472 163.367
R792 B.n474 B.n473 163.367
R793 B.n474 B.n131 163.367
R794 B.n478 B.n131 163.367
R795 B.n479 B.n478 163.367
R796 B.n480 B.n479 163.367
R797 B.n588 B.n587 163.367
R798 B.n587 B.n586 163.367
R799 B.n586 B.n95 163.367
R800 B.n582 B.n95 163.367
R801 B.n582 B.n581 163.367
R802 B.n581 B.n580 163.367
R803 B.n580 B.n97 163.367
R804 B.n576 B.n97 163.367
R805 B.n576 B.n575 163.367
R806 B.n575 B.n574 163.367
R807 B.n574 B.n99 163.367
R808 B.n570 B.n99 163.367
R809 B.n570 B.n569 163.367
R810 B.n569 B.n568 163.367
R811 B.n568 B.n101 163.367
R812 B.n564 B.n101 163.367
R813 B.n564 B.n563 163.367
R814 B.n563 B.n562 163.367
R815 B.n562 B.n103 163.367
R816 B.n558 B.n103 163.367
R817 B.n558 B.n557 163.367
R818 B.n557 B.n556 163.367
R819 B.n556 B.n105 163.367
R820 B.n552 B.n105 163.367
R821 B.n552 B.n551 163.367
R822 B.n551 B.n550 163.367
R823 B.n550 B.n107 163.367
R824 B.n546 B.n107 163.367
R825 B.n546 B.n545 163.367
R826 B.n545 B.n544 163.367
R827 B.n544 B.n109 163.367
R828 B.n540 B.n109 163.367
R829 B.n540 B.n539 163.367
R830 B.n539 B.n538 163.367
R831 B.n538 B.n111 163.367
R832 B.n534 B.n111 163.367
R833 B.n534 B.n533 163.367
R834 B.n533 B.n532 163.367
R835 B.n532 B.n113 163.367
R836 B.n528 B.n113 163.367
R837 B.n528 B.n527 163.367
R838 B.n527 B.n526 163.367
R839 B.n526 B.n115 163.367
R840 B.n522 B.n115 163.367
R841 B.n522 B.n521 163.367
R842 B.n521 B.n520 163.367
R843 B.n520 B.n117 163.367
R844 B.n516 B.n117 163.367
R845 B.n516 B.n515 163.367
R846 B.n515 B.n514 163.367
R847 B.n514 B.n119 163.367
R848 B.n510 B.n119 163.367
R849 B.n510 B.n509 163.367
R850 B.n509 B.n508 163.367
R851 B.n508 B.n121 163.367
R852 B.n504 B.n121 163.367
R853 B.n504 B.n503 163.367
R854 B.n503 B.n502 163.367
R855 B.n502 B.n123 163.367
R856 B.n498 B.n123 163.367
R857 B.n498 B.n497 163.367
R858 B.n497 B.n496 163.367
R859 B.n496 B.n125 163.367
R860 B.n492 B.n125 163.367
R861 B.n492 B.n491 163.367
R862 B.n491 B.n490 163.367
R863 B.n490 B.n127 163.367
R864 B.n486 B.n127 163.367
R865 B.n486 B.n485 163.367
R866 B.n485 B.n484 163.367
R867 B.n484 B.n129 163.367
R868 B.n798 B.n797 163.367
R869 B.n797 B.n796 163.367
R870 B.n796 B.n21 163.367
R871 B.n792 B.n21 163.367
R872 B.n792 B.n791 163.367
R873 B.n791 B.n790 163.367
R874 B.n790 B.n23 163.367
R875 B.n786 B.n23 163.367
R876 B.n786 B.n785 163.367
R877 B.n785 B.n784 163.367
R878 B.n784 B.n25 163.367
R879 B.n780 B.n25 163.367
R880 B.n780 B.n779 163.367
R881 B.n779 B.n778 163.367
R882 B.n778 B.n27 163.367
R883 B.n774 B.n27 163.367
R884 B.n774 B.n773 163.367
R885 B.n773 B.n772 163.367
R886 B.n772 B.n29 163.367
R887 B.n768 B.n29 163.367
R888 B.n768 B.n767 163.367
R889 B.n767 B.n766 163.367
R890 B.n766 B.n31 163.367
R891 B.n762 B.n31 163.367
R892 B.n762 B.n761 163.367
R893 B.n761 B.n760 163.367
R894 B.n760 B.n33 163.367
R895 B.n756 B.n33 163.367
R896 B.n756 B.n755 163.367
R897 B.n755 B.n754 163.367
R898 B.n754 B.n35 163.367
R899 B.n750 B.n35 163.367
R900 B.n750 B.n749 163.367
R901 B.n749 B.n748 163.367
R902 B.n748 B.n37 163.367
R903 B.n744 B.n37 163.367
R904 B.n744 B.n743 163.367
R905 B.n743 B.n742 163.367
R906 B.n742 B.n39 163.367
R907 B.n738 B.n39 163.367
R908 B.n738 B.n737 163.367
R909 B.n737 B.n736 163.367
R910 B.n736 B.n41 163.367
R911 B.n732 B.n41 163.367
R912 B.n732 B.n731 163.367
R913 B.n731 B.n730 163.367
R914 B.n730 B.n43 163.367
R915 B.n726 B.n43 163.367
R916 B.n726 B.n725 163.367
R917 B.n725 B.n724 163.367
R918 B.n724 B.n45 163.367
R919 B.n720 B.n45 163.367
R920 B.n720 B.n719 163.367
R921 B.n719 B.n718 163.367
R922 B.n718 B.n47 163.367
R923 B.n714 B.n47 163.367
R924 B.n714 B.n713 163.367
R925 B.n713 B.n712 163.367
R926 B.n712 B.n49 163.367
R927 B.n708 B.n49 163.367
R928 B.n708 B.n707 163.367
R929 B.n707 B.n706 163.367
R930 B.n706 B.n51 163.367
R931 B.n702 B.n51 163.367
R932 B.n702 B.n701 163.367
R933 B.n701 B.n55 163.367
R934 B.n697 B.n55 163.367
R935 B.n697 B.n696 163.367
R936 B.n696 B.n695 163.367
R937 B.n695 B.n57 163.367
R938 B.n691 B.n57 163.367
R939 B.n691 B.n690 163.367
R940 B.n690 B.n689 163.367
R941 B.n689 B.n59 163.367
R942 B.n684 B.n59 163.367
R943 B.n684 B.n683 163.367
R944 B.n683 B.n682 163.367
R945 B.n682 B.n63 163.367
R946 B.n678 B.n63 163.367
R947 B.n678 B.n677 163.367
R948 B.n677 B.n676 163.367
R949 B.n676 B.n65 163.367
R950 B.n672 B.n65 163.367
R951 B.n672 B.n671 163.367
R952 B.n671 B.n670 163.367
R953 B.n670 B.n67 163.367
R954 B.n666 B.n67 163.367
R955 B.n666 B.n665 163.367
R956 B.n665 B.n664 163.367
R957 B.n664 B.n69 163.367
R958 B.n660 B.n69 163.367
R959 B.n660 B.n659 163.367
R960 B.n659 B.n658 163.367
R961 B.n658 B.n71 163.367
R962 B.n654 B.n71 163.367
R963 B.n654 B.n653 163.367
R964 B.n653 B.n652 163.367
R965 B.n652 B.n73 163.367
R966 B.n648 B.n73 163.367
R967 B.n648 B.n647 163.367
R968 B.n647 B.n646 163.367
R969 B.n646 B.n75 163.367
R970 B.n642 B.n75 163.367
R971 B.n642 B.n641 163.367
R972 B.n641 B.n640 163.367
R973 B.n640 B.n77 163.367
R974 B.n636 B.n77 163.367
R975 B.n636 B.n635 163.367
R976 B.n635 B.n634 163.367
R977 B.n634 B.n79 163.367
R978 B.n630 B.n79 163.367
R979 B.n630 B.n629 163.367
R980 B.n629 B.n628 163.367
R981 B.n628 B.n81 163.367
R982 B.n624 B.n81 163.367
R983 B.n624 B.n623 163.367
R984 B.n623 B.n622 163.367
R985 B.n622 B.n83 163.367
R986 B.n618 B.n83 163.367
R987 B.n618 B.n617 163.367
R988 B.n617 B.n616 163.367
R989 B.n616 B.n85 163.367
R990 B.n612 B.n85 163.367
R991 B.n612 B.n611 163.367
R992 B.n611 B.n610 163.367
R993 B.n610 B.n87 163.367
R994 B.n606 B.n87 163.367
R995 B.n606 B.n605 163.367
R996 B.n605 B.n604 163.367
R997 B.n604 B.n89 163.367
R998 B.n600 B.n89 163.367
R999 B.n600 B.n599 163.367
R1000 B.n599 B.n598 163.367
R1001 B.n598 B.n91 163.367
R1002 B.n594 B.n91 163.367
R1003 B.n594 B.n593 163.367
R1004 B.n593 B.n592 163.367
R1005 B.n592 B.n93 163.367
R1006 B.n802 B.n19 163.367
R1007 B.n803 B.n802 163.367
R1008 B.n804 B.n803 163.367
R1009 B.n804 B.n17 163.367
R1010 B.n808 B.n17 163.367
R1011 B.n809 B.n808 163.367
R1012 B.n810 B.n809 163.367
R1013 B.n810 B.n15 163.367
R1014 B.n814 B.n15 163.367
R1015 B.n815 B.n814 163.367
R1016 B.n816 B.n815 163.367
R1017 B.n816 B.n13 163.367
R1018 B.n820 B.n13 163.367
R1019 B.n821 B.n820 163.367
R1020 B.n822 B.n821 163.367
R1021 B.n822 B.n11 163.367
R1022 B.n826 B.n11 163.367
R1023 B.n827 B.n826 163.367
R1024 B.n828 B.n827 163.367
R1025 B.n828 B.n9 163.367
R1026 B.n832 B.n9 163.367
R1027 B.n833 B.n832 163.367
R1028 B.n834 B.n833 163.367
R1029 B.n834 B.n7 163.367
R1030 B.n838 B.n7 163.367
R1031 B.n839 B.n838 163.367
R1032 B.n840 B.n839 163.367
R1033 B.n840 B.n5 163.367
R1034 B.n844 B.n5 163.367
R1035 B.n845 B.n844 163.367
R1036 B.n846 B.n845 163.367
R1037 B.n846 B.n3 163.367
R1038 B.n850 B.n3 163.367
R1039 B.n851 B.n850 163.367
R1040 B.n221 B.n2 163.367
R1041 B.n222 B.n221 163.367
R1042 B.n222 B.n219 163.367
R1043 B.n226 B.n219 163.367
R1044 B.n227 B.n226 163.367
R1045 B.n228 B.n227 163.367
R1046 B.n228 B.n217 163.367
R1047 B.n232 B.n217 163.367
R1048 B.n233 B.n232 163.367
R1049 B.n234 B.n233 163.367
R1050 B.n234 B.n215 163.367
R1051 B.n238 B.n215 163.367
R1052 B.n239 B.n238 163.367
R1053 B.n240 B.n239 163.367
R1054 B.n240 B.n213 163.367
R1055 B.n244 B.n213 163.367
R1056 B.n245 B.n244 163.367
R1057 B.n246 B.n245 163.367
R1058 B.n246 B.n211 163.367
R1059 B.n250 B.n211 163.367
R1060 B.n251 B.n250 163.367
R1061 B.n252 B.n251 163.367
R1062 B.n252 B.n209 163.367
R1063 B.n256 B.n209 163.367
R1064 B.n257 B.n256 163.367
R1065 B.n258 B.n257 163.367
R1066 B.n258 B.n207 163.367
R1067 B.n262 B.n207 163.367
R1068 B.n263 B.n262 163.367
R1069 B.n264 B.n263 163.367
R1070 B.n264 B.n205 163.367
R1071 B.n268 B.n205 163.367
R1072 B.n269 B.n268 163.367
R1073 B.n270 B.n269 163.367
R1074 B.n162 B.t7 137.847
R1075 B.n60 B.t5 137.847
R1076 B.n170 B.t10 137.821
R1077 B.n52 B.t2 137.821
R1078 B.n163 B.t8 107.787
R1079 B.n61 B.t4 107.787
R1080 B.n171 B.t11 107.761
R1081 B.n53 B.t1 107.761
R1082 B.n369 B.n171 59.5399
R1083 B.n164 B.n163 59.5399
R1084 B.n687 B.n61 59.5399
R1085 B.n54 B.n53 59.5399
R1086 B.n800 B.n799 30.7517
R1087 B.n590 B.n589 30.7517
R1088 B.n482 B.n481 30.7517
R1089 B.n272 B.n271 30.7517
R1090 B.n171 B.n170 30.0611
R1091 B.n163 B.n162 30.0611
R1092 B.n61 B.n60 30.0611
R1093 B.n53 B.n52 30.0611
R1094 B B.n853 18.0485
R1095 B.n801 B.n800 10.6151
R1096 B.n801 B.n18 10.6151
R1097 B.n805 B.n18 10.6151
R1098 B.n806 B.n805 10.6151
R1099 B.n807 B.n806 10.6151
R1100 B.n807 B.n16 10.6151
R1101 B.n811 B.n16 10.6151
R1102 B.n812 B.n811 10.6151
R1103 B.n813 B.n812 10.6151
R1104 B.n813 B.n14 10.6151
R1105 B.n817 B.n14 10.6151
R1106 B.n818 B.n817 10.6151
R1107 B.n819 B.n818 10.6151
R1108 B.n819 B.n12 10.6151
R1109 B.n823 B.n12 10.6151
R1110 B.n824 B.n823 10.6151
R1111 B.n825 B.n824 10.6151
R1112 B.n825 B.n10 10.6151
R1113 B.n829 B.n10 10.6151
R1114 B.n830 B.n829 10.6151
R1115 B.n831 B.n830 10.6151
R1116 B.n831 B.n8 10.6151
R1117 B.n835 B.n8 10.6151
R1118 B.n836 B.n835 10.6151
R1119 B.n837 B.n836 10.6151
R1120 B.n837 B.n6 10.6151
R1121 B.n841 B.n6 10.6151
R1122 B.n842 B.n841 10.6151
R1123 B.n843 B.n842 10.6151
R1124 B.n843 B.n4 10.6151
R1125 B.n847 B.n4 10.6151
R1126 B.n848 B.n847 10.6151
R1127 B.n849 B.n848 10.6151
R1128 B.n849 B.n0 10.6151
R1129 B.n799 B.n20 10.6151
R1130 B.n795 B.n20 10.6151
R1131 B.n795 B.n794 10.6151
R1132 B.n794 B.n793 10.6151
R1133 B.n793 B.n22 10.6151
R1134 B.n789 B.n22 10.6151
R1135 B.n789 B.n788 10.6151
R1136 B.n788 B.n787 10.6151
R1137 B.n787 B.n24 10.6151
R1138 B.n783 B.n24 10.6151
R1139 B.n783 B.n782 10.6151
R1140 B.n782 B.n781 10.6151
R1141 B.n781 B.n26 10.6151
R1142 B.n777 B.n26 10.6151
R1143 B.n777 B.n776 10.6151
R1144 B.n776 B.n775 10.6151
R1145 B.n775 B.n28 10.6151
R1146 B.n771 B.n28 10.6151
R1147 B.n771 B.n770 10.6151
R1148 B.n770 B.n769 10.6151
R1149 B.n769 B.n30 10.6151
R1150 B.n765 B.n30 10.6151
R1151 B.n765 B.n764 10.6151
R1152 B.n764 B.n763 10.6151
R1153 B.n763 B.n32 10.6151
R1154 B.n759 B.n32 10.6151
R1155 B.n759 B.n758 10.6151
R1156 B.n758 B.n757 10.6151
R1157 B.n757 B.n34 10.6151
R1158 B.n753 B.n34 10.6151
R1159 B.n753 B.n752 10.6151
R1160 B.n752 B.n751 10.6151
R1161 B.n751 B.n36 10.6151
R1162 B.n747 B.n36 10.6151
R1163 B.n747 B.n746 10.6151
R1164 B.n746 B.n745 10.6151
R1165 B.n745 B.n38 10.6151
R1166 B.n741 B.n38 10.6151
R1167 B.n741 B.n740 10.6151
R1168 B.n740 B.n739 10.6151
R1169 B.n739 B.n40 10.6151
R1170 B.n735 B.n40 10.6151
R1171 B.n735 B.n734 10.6151
R1172 B.n734 B.n733 10.6151
R1173 B.n733 B.n42 10.6151
R1174 B.n729 B.n42 10.6151
R1175 B.n729 B.n728 10.6151
R1176 B.n728 B.n727 10.6151
R1177 B.n727 B.n44 10.6151
R1178 B.n723 B.n44 10.6151
R1179 B.n723 B.n722 10.6151
R1180 B.n722 B.n721 10.6151
R1181 B.n721 B.n46 10.6151
R1182 B.n717 B.n46 10.6151
R1183 B.n717 B.n716 10.6151
R1184 B.n716 B.n715 10.6151
R1185 B.n715 B.n48 10.6151
R1186 B.n711 B.n48 10.6151
R1187 B.n711 B.n710 10.6151
R1188 B.n710 B.n709 10.6151
R1189 B.n709 B.n50 10.6151
R1190 B.n705 B.n50 10.6151
R1191 B.n705 B.n704 10.6151
R1192 B.n704 B.n703 10.6151
R1193 B.n700 B.n699 10.6151
R1194 B.n699 B.n698 10.6151
R1195 B.n698 B.n56 10.6151
R1196 B.n694 B.n56 10.6151
R1197 B.n694 B.n693 10.6151
R1198 B.n693 B.n692 10.6151
R1199 B.n692 B.n58 10.6151
R1200 B.n688 B.n58 10.6151
R1201 B.n686 B.n685 10.6151
R1202 B.n685 B.n62 10.6151
R1203 B.n681 B.n62 10.6151
R1204 B.n681 B.n680 10.6151
R1205 B.n680 B.n679 10.6151
R1206 B.n679 B.n64 10.6151
R1207 B.n675 B.n64 10.6151
R1208 B.n675 B.n674 10.6151
R1209 B.n674 B.n673 10.6151
R1210 B.n673 B.n66 10.6151
R1211 B.n669 B.n66 10.6151
R1212 B.n669 B.n668 10.6151
R1213 B.n668 B.n667 10.6151
R1214 B.n667 B.n68 10.6151
R1215 B.n663 B.n68 10.6151
R1216 B.n663 B.n662 10.6151
R1217 B.n662 B.n661 10.6151
R1218 B.n661 B.n70 10.6151
R1219 B.n657 B.n70 10.6151
R1220 B.n657 B.n656 10.6151
R1221 B.n656 B.n655 10.6151
R1222 B.n655 B.n72 10.6151
R1223 B.n651 B.n72 10.6151
R1224 B.n651 B.n650 10.6151
R1225 B.n650 B.n649 10.6151
R1226 B.n649 B.n74 10.6151
R1227 B.n645 B.n74 10.6151
R1228 B.n645 B.n644 10.6151
R1229 B.n644 B.n643 10.6151
R1230 B.n643 B.n76 10.6151
R1231 B.n639 B.n76 10.6151
R1232 B.n639 B.n638 10.6151
R1233 B.n638 B.n637 10.6151
R1234 B.n637 B.n78 10.6151
R1235 B.n633 B.n78 10.6151
R1236 B.n633 B.n632 10.6151
R1237 B.n632 B.n631 10.6151
R1238 B.n631 B.n80 10.6151
R1239 B.n627 B.n80 10.6151
R1240 B.n627 B.n626 10.6151
R1241 B.n626 B.n625 10.6151
R1242 B.n625 B.n82 10.6151
R1243 B.n621 B.n82 10.6151
R1244 B.n621 B.n620 10.6151
R1245 B.n620 B.n619 10.6151
R1246 B.n619 B.n84 10.6151
R1247 B.n615 B.n84 10.6151
R1248 B.n615 B.n614 10.6151
R1249 B.n614 B.n613 10.6151
R1250 B.n613 B.n86 10.6151
R1251 B.n609 B.n86 10.6151
R1252 B.n609 B.n608 10.6151
R1253 B.n608 B.n607 10.6151
R1254 B.n607 B.n88 10.6151
R1255 B.n603 B.n88 10.6151
R1256 B.n603 B.n602 10.6151
R1257 B.n602 B.n601 10.6151
R1258 B.n601 B.n90 10.6151
R1259 B.n597 B.n90 10.6151
R1260 B.n597 B.n596 10.6151
R1261 B.n596 B.n595 10.6151
R1262 B.n595 B.n92 10.6151
R1263 B.n591 B.n92 10.6151
R1264 B.n591 B.n590 10.6151
R1265 B.n589 B.n94 10.6151
R1266 B.n585 B.n94 10.6151
R1267 B.n585 B.n584 10.6151
R1268 B.n584 B.n583 10.6151
R1269 B.n583 B.n96 10.6151
R1270 B.n579 B.n96 10.6151
R1271 B.n579 B.n578 10.6151
R1272 B.n578 B.n577 10.6151
R1273 B.n577 B.n98 10.6151
R1274 B.n573 B.n98 10.6151
R1275 B.n573 B.n572 10.6151
R1276 B.n572 B.n571 10.6151
R1277 B.n571 B.n100 10.6151
R1278 B.n567 B.n100 10.6151
R1279 B.n567 B.n566 10.6151
R1280 B.n566 B.n565 10.6151
R1281 B.n565 B.n102 10.6151
R1282 B.n561 B.n102 10.6151
R1283 B.n561 B.n560 10.6151
R1284 B.n560 B.n559 10.6151
R1285 B.n559 B.n104 10.6151
R1286 B.n555 B.n104 10.6151
R1287 B.n555 B.n554 10.6151
R1288 B.n554 B.n553 10.6151
R1289 B.n553 B.n106 10.6151
R1290 B.n549 B.n106 10.6151
R1291 B.n549 B.n548 10.6151
R1292 B.n548 B.n547 10.6151
R1293 B.n547 B.n108 10.6151
R1294 B.n543 B.n108 10.6151
R1295 B.n543 B.n542 10.6151
R1296 B.n542 B.n541 10.6151
R1297 B.n541 B.n110 10.6151
R1298 B.n537 B.n110 10.6151
R1299 B.n537 B.n536 10.6151
R1300 B.n536 B.n535 10.6151
R1301 B.n535 B.n112 10.6151
R1302 B.n531 B.n112 10.6151
R1303 B.n531 B.n530 10.6151
R1304 B.n530 B.n529 10.6151
R1305 B.n529 B.n114 10.6151
R1306 B.n525 B.n114 10.6151
R1307 B.n525 B.n524 10.6151
R1308 B.n524 B.n523 10.6151
R1309 B.n523 B.n116 10.6151
R1310 B.n519 B.n116 10.6151
R1311 B.n519 B.n518 10.6151
R1312 B.n518 B.n517 10.6151
R1313 B.n517 B.n118 10.6151
R1314 B.n513 B.n118 10.6151
R1315 B.n513 B.n512 10.6151
R1316 B.n512 B.n511 10.6151
R1317 B.n511 B.n120 10.6151
R1318 B.n507 B.n120 10.6151
R1319 B.n507 B.n506 10.6151
R1320 B.n506 B.n505 10.6151
R1321 B.n505 B.n122 10.6151
R1322 B.n501 B.n122 10.6151
R1323 B.n501 B.n500 10.6151
R1324 B.n500 B.n499 10.6151
R1325 B.n499 B.n124 10.6151
R1326 B.n495 B.n124 10.6151
R1327 B.n495 B.n494 10.6151
R1328 B.n494 B.n493 10.6151
R1329 B.n493 B.n126 10.6151
R1330 B.n489 B.n126 10.6151
R1331 B.n489 B.n488 10.6151
R1332 B.n488 B.n487 10.6151
R1333 B.n487 B.n128 10.6151
R1334 B.n483 B.n128 10.6151
R1335 B.n483 B.n482 10.6151
R1336 B.n220 B.n1 10.6151
R1337 B.n223 B.n220 10.6151
R1338 B.n224 B.n223 10.6151
R1339 B.n225 B.n224 10.6151
R1340 B.n225 B.n218 10.6151
R1341 B.n229 B.n218 10.6151
R1342 B.n230 B.n229 10.6151
R1343 B.n231 B.n230 10.6151
R1344 B.n231 B.n216 10.6151
R1345 B.n235 B.n216 10.6151
R1346 B.n236 B.n235 10.6151
R1347 B.n237 B.n236 10.6151
R1348 B.n237 B.n214 10.6151
R1349 B.n241 B.n214 10.6151
R1350 B.n242 B.n241 10.6151
R1351 B.n243 B.n242 10.6151
R1352 B.n243 B.n212 10.6151
R1353 B.n247 B.n212 10.6151
R1354 B.n248 B.n247 10.6151
R1355 B.n249 B.n248 10.6151
R1356 B.n249 B.n210 10.6151
R1357 B.n253 B.n210 10.6151
R1358 B.n254 B.n253 10.6151
R1359 B.n255 B.n254 10.6151
R1360 B.n255 B.n208 10.6151
R1361 B.n259 B.n208 10.6151
R1362 B.n260 B.n259 10.6151
R1363 B.n261 B.n260 10.6151
R1364 B.n261 B.n206 10.6151
R1365 B.n265 B.n206 10.6151
R1366 B.n266 B.n265 10.6151
R1367 B.n267 B.n266 10.6151
R1368 B.n267 B.n204 10.6151
R1369 B.n271 B.n204 10.6151
R1370 B.n273 B.n272 10.6151
R1371 B.n273 B.n202 10.6151
R1372 B.n277 B.n202 10.6151
R1373 B.n278 B.n277 10.6151
R1374 B.n279 B.n278 10.6151
R1375 B.n279 B.n200 10.6151
R1376 B.n283 B.n200 10.6151
R1377 B.n284 B.n283 10.6151
R1378 B.n285 B.n284 10.6151
R1379 B.n285 B.n198 10.6151
R1380 B.n289 B.n198 10.6151
R1381 B.n290 B.n289 10.6151
R1382 B.n291 B.n290 10.6151
R1383 B.n291 B.n196 10.6151
R1384 B.n295 B.n196 10.6151
R1385 B.n296 B.n295 10.6151
R1386 B.n297 B.n296 10.6151
R1387 B.n297 B.n194 10.6151
R1388 B.n301 B.n194 10.6151
R1389 B.n302 B.n301 10.6151
R1390 B.n303 B.n302 10.6151
R1391 B.n303 B.n192 10.6151
R1392 B.n307 B.n192 10.6151
R1393 B.n308 B.n307 10.6151
R1394 B.n309 B.n308 10.6151
R1395 B.n309 B.n190 10.6151
R1396 B.n313 B.n190 10.6151
R1397 B.n314 B.n313 10.6151
R1398 B.n315 B.n314 10.6151
R1399 B.n315 B.n188 10.6151
R1400 B.n319 B.n188 10.6151
R1401 B.n320 B.n319 10.6151
R1402 B.n321 B.n320 10.6151
R1403 B.n321 B.n186 10.6151
R1404 B.n325 B.n186 10.6151
R1405 B.n326 B.n325 10.6151
R1406 B.n327 B.n326 10.6151
R1407 B.n327 B.n184 10.6151
R1408 B.n331 B.n184 10.6151
R1409 B.n332 B.n331 10.6151
R1410 B.n333 B.n332 10.6151
R1411 B.n333 B.n182 10.6151
R1412 B.n337 B.n182 10.6151
R1413 B.n338 B.n337 10.6151
R1414 B.n339 B.n338 10.6151
R1415 B.n339 B.n180 10.6151
R1416 B.n343 B.n180 10.6151
R1417 B.n344 B.n343 10.6151
R1418 B.n345 B.n344 10.6151
R1419 B.n345 B.n178 10.6151
R1420 B.n349 B.n178 10.6151
R1421 B.n350 B.n349 10.6151
R1422 B.n351 B.n350 10.6151
R1423 B.n351 B.n176 10.6151
R1424 B.n355 B.n176 10.6151
R1425 B.n356 B.n355 10.6151
R1426 B.n357 B.n356 10.6151
R1427 B.n357 B.n174 10.6151
R1428 B.n361 B.n174 10.6151
R1429 B.n362 B.n361 10.6151
R1430 B.n363 B.n362 10.6151
R1431 B.n363 B.n172 10.6151
R1432 B.n367 B.n172 10.6151
R1433 B.n368 B.n367 10.6151
R1434 B.n370 B.n168 10.6151
R1435 B.n374 B.n168 10.6151
R1436 B.n375 B.n374 10.6151
R1437 B.n376 B.n375 10.6151
R1438 B.n376 B.n166 10.6151
R1439 B.n380 B.n166 10.6151
R1440 B.n381 B.n380 10.6151
R1441 B.n382 B.n381 10.6151
R1442 B.n386 B.n385 10.6151
R1443 B.n387 B.n386 10.6151
R1444 B.n387 B.n160 10.6151
R1445 B.n391 B.n160 10.6151
R1446 B.n392 B.n391 10.6151
R1447 B.n393 B.n392 10.6151
R1448 B.n393 B.n158 10.6151
R1449 B.n397 B.n158 10.6151
R1450 B.n398 B.n397 10.6151
R1451 B.n399 B.n398 10.6151
R1452 B.n399 B.n156 10.6151
R1453 B.n403 B.n156 10.6151
R1454 B.n404 B.n403 10.6151
R1455 B.n405 B.n404 10.6151
R1456 B.n405 B.n154 10.6151
R1457 B.n409 B.n154 10.6151
R1458 B.n410 B.n409 10.6151
R1459 B.n411 B.n410 10.6151
R1460 B.n411 B.n152 10.6151
R1461 B.n415 B.n152 10.6151
R1462 B.n416 B.n415 10.6151
R1463 B.n417 B.n416 10.6151
R1464 B.n417 B.n150 10.6151
R1465 B.n421 B.n150 10.6151
R1466 B.n422 B.n421 10.6151
R1467 B.n423 B.n422 10.6151
R1468 B.n423 B.n148 10.6151
R1469 B.n427 B.n148 10.6151
R1470 B.n428 B.n427 10.6151
R1471 B.n429 B.n428 10.6151
R1472 B.n429 B.n146 10.6151
R1473 B.n433 B.n146 10.6151
R1474 B.n434 B.n433 10.6151
R1475 B.n435 B.n434 10.6151
R1476 B.n435 B.n144 10.6151
R1477 B.n439 B.n144 10.6151
R1478 B.n440 B.n439 10.6151
R1479 B.n441 B.n440 10.6151
R1480 B.n441 B.n142 10.6151
R1481 B.n445 B.n142 10.6151
R1482 B.n446 B.n445 10.6151
R1483 B.n447 B.n446 10.6151
R1484 B.n447 B.n140 10.6151
R1485 B.n451 B.n140 10.6151
R1486 B.n452 B.n451 10.6151
R1487 B.n453 B.n452 10.6151
R1488 B.n453 B.n138 10.6151
R1489 B.n457 B.n138 10.6151
R1490 B.n458 B.n457 10.6151
R1491 B.n459 B.n458 10.6151
R1492 B.n459 B.n136 10.6151
R1493 B.n463 B.n136 10.6151
R1494 B.n464 B.n463 10.6151
R1495 B.n465 B.n464 10.6151
R1496 B.n465 B.n134 10.6151
R1497 B.n469 B.n134 10.6151
R1498 B.n470 B.n469 10.6151
R1499 B.n471 B.n470 10.6151
R1500 B.n471 B.n132 10.6151
R1501 B.n475 B.n132 10.6151
R1502 B.n476 B.n475 10.6151
R1503 B.n477 B.n476 10.6151
R1504 B.n477 B.n130 10.6151
R1505 B.n481 B.n130 10.6151
R1506 B.n853 B.n0 8.11757
R1507 B.n853 B.n1 8.11757
R1508 B.n700 B.n54 6.5566
R1509 B.n688 B.n687 6.5566
R1510 B.n370 B.n369 6.5566
R1511 B.n382 B.n164 6.5566
R1512 B.n703 B.n54 4.05904
R1513 B.n687 B.n686 4.05904
R1514 B.n369 B.n368 4.05904
R1515 B.n385 B.n164 4.05904
C0 VN VTAIL 13.677401f
C1 VP VDD1 14.1727f
C2 VDD2 w_n2830_n4930# 2.88875f
C3 VTAIL VP 13.6921f
C4 VN VP 7.80966f
C5 VDD2 B 2.57698f
C6 VDD2 VDD1 1.29253f
C7 B w_n2830_n4930# 10.4155f
C8 VTAIL VDD2 17.0219f
C9 VN VDD2 13.920599f
C10 VDD1 w_n2830_n4930# 2.81692f
C11 VDD2 VP 0.408405f
C12 VTAIL w_n2830_n4930# 4.20626f
C13 B VDD1 2.51275f
C14 VN w_n2830_n4930# 5.78347f
C15 VTAIL B 4.57959f
C16 VN B 1.02372f
C17 VP w_n2830_n4930# 6.14766f
C18 VTAIL VDD1 16.9858f
C19 VP B 1.62852f
C20 VN VDD1 0.149917f
C21 VDD2 VSUBS 1.871758f
C22 VDD1 VSUBS 1.613539f
C23 VTAIL VSUBS 1.201139f
C24 VN VSUBS 6.06628f
C25 VP VSUBS 2.781483f
C26 B VSUBS 4.316177f
C27 w_n2830_n4930# VSUBS 0.170377p
C28 B.n0 VSUBS 0.007339f
C29 B.n1 VSUBS 0.007339f
C30 B.n2 VSUBS 0.010854f
C31 B.n3 VSUBS 0.008318f
C32 B.n4 VSUBS 0.008318f
C33 B.n5 VSUBS 0.008318f
C34 B.n6 VSUBS 0.008318f
C35 B.n7 VSUBS 0.008318f
C36 B.n8 VSUBS 0.008318f
C37 B.n9 VSUBS 0.008318f
C38 B.n10 VSUBS 0.008318f
C39 B.n11 VSUBS 0.008318f
C40 B.n12 VSUBS 0.008318f
C41 B.n13 VSUBS 0.008318f
C42 B.n14 VSUBS 0.008318f
C43 B.n15 VSUBS 0.008318f
C44 B.n16 VSUBS 0.008318f
C45 B.n17 VSUBS 0.008318f
C46 B.n18 VSUBS 0.008318f
C47 B.n19 VSUBS 0.018142f
C48 B.n20 VSUBS 0.008318f
C49 B.n21 VSUBS 0.008318f
C50 B.n22 VSUBS 0.008318f
C51 B.n23 VSUBS 0.008318f
C52 B.n24 VSUBS 0.008318f
C53 B.n25 VSUBS 0.008318f
C54 B.n26 VSUBS 0.008318f
C55 B.n27 VSUBS 0.008318f
C56 B.n28 VSUBS 0.008318f
C57 B.n29 VSUBS 0.008318f
C58 B.n30 VSUBS 0.008318f
C59 B.n31 VSUBS 0.008318f
C60 B.n32 VSUBS 0.008318f
C61 B.n33 VSUBS 0.008318f
C62 B.n34 VSUBS 0.008318f
C63 B.n35 VSUBS 0.008318f
C64 B.n36 VSUBS 0.008318f
C65 B.n37 VSUBS 0.008318f
C66 B.n38 VSUBS 0.008318f
C67 B.n39 VSUBS 0.008318f
C68 B.n40 VSUBS 0.008318f
C69 B.n41 VSUBS 0.008318f
C70 B.n42 VSUBS 0.008318f
C71 B.n43 VSUBS 0.008318f
C72 B.n44 VSUBS 0.008318f
C73 B.n45 VSUBS 0.008318f
C74 B.n46 VSUBS 0.008318f
C75 B.n47 VSUBS 0.008318f
C76 B.n48 VSUBS 0.008318f
C77 B.n49 VSUBS 0.008318f
C78 B.n50 VSUBS 0.008318f
C79 B.n51 VSUBS 0.008318f
C80 B.t1 VSUBS 0.799752f
C81 B.t2 VSUBS 0.814394f
C82 B.t0 VSUBS 1.19482f
C83 B.n52 VSUBS 0.321531f
C84 B.n53 VSUBS 0.078991f
C85 B.n54 VSUBS 0.019272f
C86 B.n55 VSUBS 0.008318f
C87 B.n56 VSUBS 0.008318f
C88 B.n57 VSUBS 0.008318f
C89 B.n58 VSUBS 0.008318f
C90 B.n59 VSUBS 0.008318f
C91 B.t4 VSUBS 0.799718f
C92 B.t5 VSUBS 0.814364f
C93 B.t3 VSUBS 1.19482f
C94 B.n60 VSUBS 0.321561f
C95 B.n61 VSUBS 0.079026f
C96 B.n62 VSUBS 0.008318f
C97 B.n63 VSUBS 0.008318f
C98 B.n64 VSUBS 0.008318f
C99 B.n65 VSUBS 0.008318f
C100 B.n66 VSUBS 0.008318f
C101 B.n67 VSUBS 0.008318f
C102 B.n68 VSUBS 0.008318f
C103 B.n69 VSUBS 0.008318f
C104 B.n70 VSUBS 0.008318f
C105 B.n71 VSUBS 0.008318f
C106 B.n72 VSUBS 0.008318f
C107 B.n73 VSUBS 0.008318f
C108 B.n74 VSUBS 0.008318f
C109 B.n75 VSUBS 0.008318f
C110 B.n76 VSUBS 0.008318f
C111 B.n77 VSUBS 0.008318f
C112 B.n78 VSUBS 0.008318f
C113 B.n79 VSUBS 0.008318f
C114 B.n80 VSUBS 0.008318f
C115 B.n81 VSUBS 0.008318f
C116 B.n82 VSUBS 0.008318f
C117 B.n83 VSUBS 0.008318f
C118 B.n84 VSUBS 0.008318f
C119 B.n85 VSUBS 0.008318f
C120 B.n86 VSUBS 0.008318f
C121 B.n87 VSUBS 0.008318f
C122 B.n88 VSUBS 0.008318f
C123 B.n89 VSUBS 0.008318f
C124 B.n90 VSUBS 0.008318f
C125 B.n91 VSUBS 0.008318f
C126 B.n92 VSUBS 0.008318f
C127 B.n93 VSUBS 0.019288f
C128 B.n94 VSUBS 0.008318f
C129 B.n95 VSUBS 0.008318f
C130 B.n96 VSUBS 0.008318f
C131 B.n97 VSUBS 0.008318f
C132 B.n98 VSUBS 0.008318f
C133 B.n99 VSUBS 0.008318f
C134 B.n100 VSUBS 0.008318f
C135 B.n101 VSUBS 0.008318f
C136 B.n102 VSUBS 0.008318f
C137 B.n103 VSUBS 0.008318f
C138 B.n104 VSUBS 0.008318f
C139 B.n105 VSUBS 0.008318f
C140 B.n106 VSUBS 0.008318f
C141 B.n107 VSUBS 0.008318f
C142 B.n108 VSUBS 0.008318f
C143 B.n109 VSUBS 0.008318f
C144 B.n110 VSUBS 0.008318f
C145 B.n111 VSUBS 0.008318f
C146 B.n112 VSUBS 0.008318f
C147 B.n113 VSUBS 0.008318f
C148 B.n114 VSUBS 0.008318f
C149 B.n115 VSUBS 0.008318f
C150 B.n116 VSUBS 0.008318f
C151 B.n117 VSUBS 0.008318f
C152 B.n118 VSUBS 0.008318f
C153 B.n119 VSUBS 0.008318f
C154 B.n120 VSUBS 0.008318f
C155 B.n121 VSUBS 0.008318f
C156 B.n122 VSUBS 0.008318f
C157 B.n123 VSUBS 0.008318f
C158 B.n124 VSUBS 0.008318f
C159 B.n125 VSUBS 0.008318f
C160 B.n126 VSUBS 0.008318f
C161 B.n127 VSUBS 0.008318f
C162 B.n128 VSUBS 0.008318f
C163 B.n129 VSUBS 0.018142f
C164 B.n130 VSUBS 0.008318f
C165 B.n131 VSUBS 0.008318f
C166 B.n132 VSUBS 0.008318f
C167 B.n133 VSUBS 0.008318f
C168 B.n134 VSUBS 0.008318f
C169 B.n135 VSUBS 0.008318f
C170 B.n136 VSUBS 0.008318f
C171 B.n137 VSUBS 0.008318f
C172 B.n138 VSUBS 0.008318f
C173 B.n139 VSUBS 0.008318f
C174 B.n140 VSUBS 0.008318f
C175 B.n141 VSUBS 0.008318f
C176 B.n142 VSUBS 0.008318f
C177 B.n143 VSUBS 0.008318f
C178 B.n144 VSUBS 0.008318f
C179 B.n145 VSUBS 0.008318f
C180 B.n146 VSUBS 0.008318f
C181 B.n147 VSUBS 0.008318f
C182 B.n148 VSUBS 0.008318f
C183 B.n149 VSUBS 0.008318f
C184 B.n150 VSUBS 0.008318f
C185 B.n151 VSUBS 0.008318f
C186 B.n152 VSUBS 0.008318f
C187 B.n153 VSUBS 0.008318f
C188 B.n154 VSUBS 0.008318f
C189 B.n155 VSUBS 0.008318f
C190 B.n156 VSUBS 0.008318f
C191 B.n157 VSUBS 0.008318f
C192 B.n158 VSUBS 0.008318f
C193 B.n159 VSUBS 0.008318f
C194 B.n160 VSUBS 0.008318f
C195 B.n161 VSUBS 0.008318f
C196 B.t8 VSUBS 0.799718f
C197 B.t7 VSUBS 0.814364f
C198 B.t6 VSUBS 1.19482f
C199 B.n162 VSUBS 0.321561f
C200 B.n163 VSUBS 0.079026f
C201 B.n164 VSUBS 0.019272f
C202 B.n165 VSUBS 0.008318f
C203 B.n166 VSUBS 0.008318f
C204 B.n167 VSUBS 0.008318f
C205 B.n168 VSUBS 0.008318f
C206 B.n169 VSUBS 0.008318f
C207 B.t11 VSUBS 0.799752f
C208 B.t10 VSUBS 0.814394f
C209 B.t9 VSUBS 1.19482f
C210 B.n170 VSUBS 0.321531f
C211 B.n171 VSUBS 0.078991f
C212 B.n172 VSUBS 0.008318f
C213 B.n173 VSUBS 0.008318f
C214 B.n174 VSUBS 0.008318f
C215 B.n175 VSUBS 0.008318f
C216 B.n176 VSUBS 0.008318f
C217 B.n177 VSUBS 0.008318f
C218 B.n178 VSUBS 0.008318f
C219 B.n179 VSUBS 0.008318f
C220 B.n180 VSUBS 0.008318f
C221 B.n181 VSUBS 0.008318f
C222 B.n182 VSUBS 0.008318f
C223 B.n183 VSUBS 0.008318f
C224 B.n184 VSUBS 0.008318f
C225 B.n185 VSUBS 0.008318f
C226 B.n186 VSUBS 0.008318f
C227 B.n187 VSUBS 0.008318f
C228 B.n188 VSUBS 0.008318f
C229 B.n189 VSUBS 0.008318f
C230 B.n190 VSUBS 0.008318f
C231 B.n191 VSUBS 0.008318f
C232 B.n192 VSUBS 0.008318f
C233 B.n193 VSUBS 0.008318f
C234 B.n194 VSUBS 0.008318f
C235 B.n195 VSUBS 0.008318f
C236 B.n196 VSUBS 0.008318f
C237 B.n197 VSUBS 0.008318f
C238 B.n198 VSUBS 0.008318f
C239 B.n199 VSUBS 0.008318f
C240 B.n200 VSUBS 0.008318f
C241 B.n201 VSUBS 0.008318f
C242 B.n202 VSUBS 0.008318f
C243 B.n203 VSUBS 0.019288f
C244 B.n204 VSUBS 0.008318f
C245 B.n205 VSUBS 0.008318f
C246 B.n206 VSUBS 0.008318f
C247 B.n207 VSUBS 0.008318f
C248 B.n208 VSUBS 0.008318f
C249 B.n209 VSUBS 0.008318f
C250 B.n210 VSUBS 0.008318f
C251 B.n211 VSUBS 0.008318f
C252 B.n212 VSUBS 0.008318f
C253 B.n213 VSUBS 0.008318f
C254 B.n214 VSUBS 0.008318f
C255 B.n215 VSUBS 0.008318f
C256 B.n216 VSUBS 0.008318f
C257 B.n217 VSUBS 0.008318f
C258 B.n218 VSUBS 0.008318f
C259 B.n219 VSUBS 0.008318f
C260 B.n220 VSUBS 0.008318f
C261 B.n221 VSUBS 0.008318f
C262 B.n222 VSUBS 0.008318f
C263 B.n223 VSUBS 0.008318f
C264 B.n224 VSUBS 0.008318f
C265 B.n225 VSUBS 0.008318f
C266 B.n226 VSUBS 0.008318f
C267 B.n227 VSUBS 0.008318f
C268 B.n228 VSUBS 0.008318f
C269 B.n229 VSUBS 0.008318f
C270 B.n230 VSUBS 0.008318f
C271 B.n231 VSUBS 0.008318f
C272 B.n232 VSUBS 0.008318f
C273 B.n233 VSUBS 0.008318f
C274 B.n234 VSUBS 0.008318f
C275 B.n235 VSUBS 0.008318f
C276 B.n236 VSUBS 0.008318f
C277 B.n237 VSUBS 0.008318f
C278 B.n238 VSUBS 0.008318f
C279 B.n239 VSUBS 0.008318f
C280 B.n240 VSUBS 0.008318f
C281 B.n241 VSUBS 0.008318f
C282 B.n242 VSUBS 0.008318f
C283 B.n243 VSUBS 0.008318f
C284 B.n244 VSUBS 0.008318f
C285 B.n245 VSUBS 0.008318f
C286 B.n246 VSUBS 0.008318f
C287 B.n247 VSUBS 0.008318f
C288 B.n248 VSUBS 0.008318f
C289 B.n249 VSUBS 0.008318f
C290 B.n250 VSUBS 0.008318f
C291 B.n251 VSUBS 0.008318f
C292 B.n252 VSUBS 0.008318f
C293 B.n253 VSUBS 0.008318f
C294 B.n254 VSUBS 0.008318f
C295 B.n255 VSUBS 0.008318f
C296 B.n256 VSUBS 0.008318f
C297 B.n257 VSUBS 0.008318f
C298 B.n258 VSUBS 0.008318f
C299 B.n259 VSUBS 0.008318f
C300 B.n260 VSUBS 0.008318f
C301 B.n261 VSUBS 0.008318f
C302 B.n262 VSUBS 0.008318f
C303 B.n263 VSUBS 0.008318f
C304 B.n264 VSUBS 0.008318f
C305 B.n265 VSUBS 0.008318f
C306 B.n266 VSUBS 0.008318f
C307 B.n267 VSUBS 0.008318f
C308 B.n268 VSUBS 0.008318f
C309 B.n269 VSUBS 0.008318f
C310 B.n270 VSUBS 0.018142f
C311 B.n271 VSUBS 0.018142f
C312 B.n272 VSUBS 0.019288f
C313 B.n273 VSUBS 0.008318f
C314 B.n274 VSUBS 0.008318f
C315 B.n275 VSUBS 0.008318f
C316 B.n276 VSUBS 0.008318f
C317 B.n277 VSUBS 0.008318f
C318 B.n278 VSUBS 0.008318f
C319 B.n279 VSUBS 0.008318f
C320 B.n280 VSUBS 0.008318f
C321 B.n281 VSUBS 0.008318f
C322 B.n282 VSUBS 0.008318f
C323 B.n283 VSUBS 0.008318f
C324 B.n284 VSUBS 0.008318f
C325 B.n285 VSUBS 0.008318f
C326 B.n286 VSUBS 0.008318f
C327 B.n287 VSUBS 0.008318f
C328 B.n288 VSUBS 0.008318f
C329 B.n289 VSUBS 0.008318f
C330 B.n290 VSUBS 0.008318f
C331 B.n291 VSUBS 0.008318f
C332 B.n292 VSUBS 0.008318f
C333 B.n293 VSUBS 0.008318f
C334 B.n294 VSUBS 0.008318f
C335 B.n295 VSUBS 0.008318f
C336 B.n296 VSUBS 0.008318f
C337 B.n297 VSUBS 0.008318f
C338 B.n298 VSUBS 0.008318f
C339 B.n299 VSUBS 0.008318f
C340 B.n300 VSUBS 0.008318f
C341 B.n301 VSUBS 0.008318f
C342 B.n302 VSUBS 0.008318f
C343 B.n303 VSUBS 0.008318f
C344 B.n304 VSUBS 0.008318f
C345 B.n305 VSUBS 0.008318f
C346 B.n306 VSUBS 0.008318f
C347 B.n307 VSUBS 0.008318f
C348 B.n308 VSUBS 0.008318f
C349 B.n309 VSUBS 0.008318f
C350 B.n310 VSUBS 0.008318f
C351 B.n311 VSUBS 0.008318f
C352 B.n312 VSUBS 0.008318f
C353 B.n313 VSUBS 0.008318f
C354 B.n314 VSUBS 0.008318f
C355 B.n315 VSUBS 0.008318f
C356 B.n316 VSUBS 0.008318f
C357 B.n317 VSUBS 0.008318f
C358 B.n318 VSUBS 0.008318f
C359 B.n319 VSUBS 0.008318f
C360 B.n320 VSUBS 0.008318f
C361 B.n321 VSUBS 0.008318f
C362 B.n322 VSUBS 0.008318f
C363 B.n323 VSUBS 0.008318f
C364 B.n324 VSUBS 0.008318f
C365 B.n325 VSUBS 0.008318f
C366 B.n326 VSUBS 0.008318f
C367 B.n327 VSUBS 0.008318f
C368 B.n328 VSUBS 0.008318f
C369 B.n329 VSUBS 0.008318f
C370 B.n330 VSUBS 0.008318f
C371 B.n331 VSUBS 0.008318f
C372 B.n332 VSUBS 0.008318f
C373 B.n333 VSUBS 0.008318f
C374 B.n334 VSUBS 0.008318f
C375 B.n335 VSUBS 0.008318f
C376 B.n336 VSUBS 0.008318f
C377 B.n337 VSUBS 0.008318f
C378 B.n338 VSUBS 0.008318f
C379 B.n339 VSUBS 0.008318f
C380 B.n340 VSUBS 0.008318f
C381 B.n341 VSUBS 0.008318f
C382 B.n342 VSUBS 0.008318f
C383 B.n343 VSUBS 0.008318f
C384 B.n344 VSUBS 0.008318f
C385 B.n345 VSUBS 0.008318f
C386 B.n346 VSUBS 0.008318f
C387 B.n347 VSUBS 0.008318f
C388 B.n348 VSUBS 0.008318f
C389 B.n349 VSUBS 0.008318f
C390 B.n350 VSUBS 0.008318f
C391 B.n351 VSUBS 0.008318f
C392 B.n352 VSUBS 0.008318f
C393 B.n353 VSUBS 0.008318f
C394 B.n354 VSUBS 0.008318f
C395 B.n355 VSUBS 0.008318f
C396 B.n356 VSUBS 0.008318f
C397 B.n357 VSUBS 0.008318f
C398 B.n358 VSUBS 0.008318f
C399 B.n359 VSUBS 0.008318f
C400 B.n360 VSUBS 0.008318f
C401 B.n361 VSUBS 0.008318f
C402 B.n362 VSUBS 0.008318f
C403 B.n363 VSUBS 0.008318f
C404 B.n364 VSUBS 0.008318f
C405 B.n365 VSUBS 0.008318f
C406 B.n366 VSUBS 0.008318f
C407 B.n367 VSUBS 0.008318f
C408 B.n368 VSUBS 0.005749f
C409 B.n369 VSUBS 0.019272f
C410 B.n370 VSUBS 0.006728f
C411 B.n371 VSUBS 0.008318f
C412 B.n372 VSUBS 0.008318f
C413 B.n373 VSUBS 0.008318f
C414 B.n374 VSUBS 0.008318f
C415 B.n375 VSUBS 0.008318f
C416 B.n376 VSUBS 0.008318f
C417 B.n377 VSUBS 0.008318f
C418 B.n378 VSUBS 0.008318f
C419 B.n379 VSUBS 0.008318f
C420 B.n380 VSUBS 0.008318f
C421 B.n381 VSUBS 0.008318f
C422 B.n382 VSUBS 0.006728f
C423 B.n383 VSUBS 0.008318f
C424 B.n384 VSUBS 0.008318f
C425 B.n385 VSUBS 0.005749f
C426 B.n386 VSUBS 0.008318f
C427 B.n387 VSUBS 0.008318f
C428 B.n388 VSUBS 0.008318f
C429 B.n389 VSUBS 0.008318f
C430 B.n390 VSUBS 0.008318f
C431 B.n391 VSUBS 0.008318f
C432 B.n392 VSUBS 0.008318f
C433 B.n393 VSUBS 0.008318f
C434 B.n394 VSUBS 0.008318f
C435 B.n395 VSUBS 0.008318f
C436 B.n396 VSUBS 0.008318f
C437 B.n397 VSUBS 0.008318f
C438 B.n398 VSUBS 0.008318f
C439 B.n399 VSUBS 0.008318f
C440 B.n400 VSUBS 0.008318f
C441 B.n401 VSUBS 0.008318f
C442 B.n402 VSUBS 0.008318f
C443 B.n403 VSUBS 0.008318f
C444 B.n404 VSUBS 0.008318f
C445 B.n405 VSUBS 0.008318f
C446 B.n406 VSUBS 0.008318f
C447 B.n407 VSUBS 0.008318f
C448 B.n408 VSUBS 0.008318f
C449 B.n409 VSUBS 0.008318f
C450 B.n410 VSUBS 0.008318f
C451 B.n411 VSUBS 0.008318f
C452 B.n412 VSUBS 0.008318f
C453 B.n413 VSUBS 0.008318f
C454 B.n414 VSUBS 0.008318f
C455 B.n415 VSUBS 0.008318f
C456 B.n416 VSUBS 0.008318f
C457 B.n417 VSUBS 0.008318f
C458 B.n418 VSUBS 0.008318f
C459 B.n419 VSUBS 0.008318f
C460 B.n420 VSUBS 0.008318f
C461 B.n421 VSUBS 0.008318f
C462 B.n422 VSUBS 0.008318f
C463 B.n423 VSUBS 0.008318f
C464 B.n424 VSUBS 0.008318f
C465 B.n425 VSUBS 0.008318f
C466 B.n426 VSUBS 0.008318f
C467 B.n427 VSUBS 0.008318f
C468 B.n428 VSUBS 0.008318f
C469 B.n429 VSUBS 0.008318f
C470 B.n430 VSUBS 0.008318f
C471 B.n431 VSUBS 0.008318f
C472 B.n432 VSUBS 0.008318f
C473 B.n433 VSUBS 0.008318f
C474 B.n434 VSUBS 0.008318f
C475 B.n435 VSUBS 0.008318f
C476 B.n436 VSUBS 0.008318f
C477 B.n437 VSUBS 0.008318f
C478 B.n438 VSUBS 0.008318f
C479 B.n439 VSUBS 0.008318f
C480 B.n440 VSUBS 0.008318f
C481 B.n441 VSUBS 0.008318f
C482 B.n442 VSUBS 0.008318f
C483 B.n443 VSUBS 0.008318f
C484 B.n444 VSUBS 0.008318f
C485 B.n445 VSUBS 0.008318f
C486 B.n446 VSUBS 0.008318f
C487 B.n447 VSUBS 0.008318f
C488 B.n448 VSUBS 0.008318f
C489 B.n449 VSUBS 0.008318f
C490 B.n450 VSUBS 0.008318f
C491 B.n451 VSUBS 0.008318f
C492 B.n452 VSUBS 0.008318f
C493 B.n453 VSUBS 0.008318f
C494 B.n454 VSUBS 0.008318f
C495 B.n455 VSUBS 0.008318f
C496 B.n456 VSUBS 0.008318f
C497 B.n457 VSUBS 0.008318f
C498 B.n458 VSUBS 0.008318f
C499 B.n459 VSUBS 0.008318f
C500 B.n460 VSUBS 0.008318f
C501 B.n461 VSUBS 0.008318f
C502 B.n462 VSUBS 0.008318f
C503 B.n463 VSUBS 0.008318f
C504 B.n464 VSUBS 0.008318f
C505 B.n465 VSUBS 0.008318f
C506 B.n466 VSUBS 0.008318f
C507 B.n467 VSUBS 0.008318f
C508 B.n468 VSUBS 0.008318f
C509 B.n469 VSUBS 0.008318f
C510 B.n470 VSUBS 0.008318f
C511 B.n471 VSUBS 0.008318f
C512 B.n472 VSUBS 0.008318f
C513 B.n473 VSUBS 0.008318f
C514 B.n474 VSUBS 0.008318f
C515 B.n475 VSUBS 0.008318f
C516 B.n476 VSUBS 0.008318f
C517 B.n477 VSUBS 0.008318f
C518 B.n478 VSUBS 0.008318f
C519 B.n479 VSUBS 0.008318f
C520 B.n480 VSUBS 0.019288f
C521 B.n481 VSUBS 0.018244f
C522 B.n482 VSUBS 0.019186f
C523 B.n483 VSUBS 0.008318f
C524 B.n484 VSUBS 0.008318f
C525 B.n485 VSUBS 0.008318f
C526 B.n486 VSUBS 0.008318f
C527 B.n487 VSUBS 0.008318f
C528 B.n488 VSUBS 0.008318f
C529 B.n489 VSUBS 0.008318f
C530 B.n490 VSUBS 0.008318f
C531 B.n491 VSUBS 0.008318f
C532 B.n492 VSUBS 0.008318f
C533 B.n493 VSUBS 0.008318f
C534 B.n494 VSUBS 0.008318f
C535 B.n495 VSUBS 0.008318f
C536 B.n496 VSUBS 0.008318f
C537 B.n497 VSUBS 0.008318f
C538 B.n498 VSUBS 0.008318f
C539 B.n499 VSUBS 0.008318f
C540 B.n500 VSUBS 0.008318f
C541 B.n501 VSUBS 0.008318f
C542 B.n502 VSUBS 0.008318f
C543 B.n503 VSUBS 0.008318f
C544 B.n504 VSUBS 0.008318f
C545 B.n505 VSUBS 0.008318f
C546 B.n506 VSUBS 0.008318f
C547 B.n507 VSUBS 0.008318f
C548 B.n508 VSUBS 0.008318f
C549 B.n509 VSUBS 0.008318f
C550 B.n510 VSUBS 0.008318f
C551 B.n511 VSUBS 0.008318f
C552 B.n512 VSUBS 0.008318f
C553 B.n513 VSUBS 0.008318f
C554 B.n514 VSUBS 0.008318f
C555 B.n515 VSUBS 0.008318f
C556 B.n516 VSUBS 0.008318f
C557 B.n517 VSUBS 0.008318f
C558 B.n518 VSUBS 0.008318f
C559 B.n519 VSUBS 0.008318f
C560 B.n520 VSUBS 0.008318f
C561 B.n521 VSUBS 0.008318f
C562 B.n522 VSUBS 0.008318f
C563 B.n523 VSUBS 0.008318f
C564 B.n524 VSUBS 0.008318f
C565 B.n525 VSUBS 0.008318f
C566 B.n526 VSUBS 0.008318f
C567 B.n527 VSUBS 0.008318f
C568 B.n528 VSUBS 0.008318f
C569 B.n529 VSUBS 0.008318f
C570 B.n530 VSUBS 0.008318f
C571 B.n531 VSUBS 0.008318f
C572 B.n532 VSUBS 0.008318f
C573 B.n533 VSUBS 0.008318f
C574 B.n534 VSUBS 0.008318f
C575 B.n535 VSUBS 0.008318f
C576 B.n536 VSUBS 0.008318f
C577 B.n537 VSUBS 0.008318f
C578 B.n538 VSUBS 0.008318f
C579 B.n539 VSUBS 0.008318f
C580 B.n540 VSUBS 0.008318f
C581 B.n541 VSUBS 0.008318f
C582 B.n542 VSUBS 0.008318f
C583 B.n543 VSUBS 0.008318f
C584 B.n544 VSUBS 0.008318f
C585 B.n545 VSUBS 0.008318f
C586 B.n546 VSUBS 0.008318f
C587 B.n547 VSUBS 0.008318f
C588 B.n548 VSUBS 0.008318f
C589 B.n549 VSUBS 0.008318f
C590 B.n550 VSUBS 0.008318f
C591 B.n551 VSUBS 0.008318f
C592 B.n552 VSUBS 0.008318f
C593 B.n553 VSUBS 0.008318f
C594 B.n554 VSUBS 0.008318f
C595 B.n555 VSUBS 0.008318f
C596 B.n556 VSUBS 0.008318f
C597 B.n557 VSUBS 0.008318f
C598 B.n558 VSUBS 0.008318f
C599 B.n559 VSUBS 0.008318f
C600 B.n560 VSUBS 0.008318f
C601 B.n561 VSUBS 0.008318f
C602 B.n562 VSUBS 0.008318f
C603 B.n563 VSUBS 0.008318f
C604 B.n564 VSUBS 0.008318f
C605 B.n565 VSUBS 0.008318f
C606 B.n566 VSUBS 0.008318f
C607 B.n567 VSUBS 0.008318f
C608 B.n568 VSUBS 0.008318f
C609 B.n569 VSUBS 0.008318f
C610 B.n570 VSUBS 0.008318f
C611 B.n571 VSUBS 0.008318f
C612 B.n572 VSUBS 0.008318f
C613 B.n573 VSUBS 0.008318f
C614 B.n574 VSUBS 0.008318f
C615 B.n575 VSUBS 0.008318f
C616 B.n576 VSUBS 0.008318f
C617 B.n577 VSUBS 0.008318f
C618 B.n578 VSUBS 0.008318f
C619 B.n579 VSUBS 0.008318f
C620 B.n580 VSUBS 0.008318f
C621 B.n581 VSUBS 0.008318f
C622 B.n582 VSUBS 0.008318f
C623 B.n583 VSUBS 0.008318f
C624 B.n584 VSUBS 0.008318f
C625 B.n585 VSUBS 0.008318f
C626 B.n586 VSUBS 0.008318f
C627 B.n587 VSUBS 0.008318f
C628 B.n588 VSUBS 0.018142f
C629 B.n589 VSUBS 0.018142f
C630 B.n590 VSUBS 0.019288f
C631 B.n591 VSUBS 0.008318f
C632 B.n592 VSUBS 0.008318f
C633 B.n593 VSUBS 0.008318f
C634 B.n594 VSUBS 0.008318f
C635 B.n595 VSUBS 0.008318f
C636 B.n596 VSUBS 0.008318f
C637 B.n597 VSUBS 0.008318f
C638 B.n598 VSUBS 0.008318f
C639 B.n599 VSUBS 0.008318f
C640 B.n600 VSUBS 0.008318f
C641 B.n601 VSUBS 0.008318f
C642 B.n602 VSUBS 0.008318f
C643 B.n603 VSUBS 0.008318f
C644 B.n604 VSUBS 0.008318f
C645 B.n605 VSUBS 0.008318f
C646 B.n606 VSUBS 0.008318f
C647 B.n607 VSUBS 0.008318f
C648 B.n608 VSUBS 0.008318f
C649 B.n609 VSUBS 0.008318f
C650 B.n610 VSUBS 0.008318f
C651 B.n611 VSUBS 0.008318f
C652 B.n612 VSUBS 0.008318f
C653 B.n613 VSUBS 0.008318f
C654 B.n614 VSUBS 0.008318f
C655 B.n615 VSUBS 0.008318f
C656 B.n616 VSUBS 0.008318f
C657 B.n617 VSUBS 0.008318f
C658 B.n618 VSUBS 0.008318f
C659 B.n619 VSUBS 0.008318f
C660 B.n620 VSUBS 0.008318f
C661 B.n621 VSUBS 0.008318f
C662 B.n622 VSUBS 0.008318f
C663 B.n623 VSUBS 0.008318f
C664 B.n624 VSUBS 0.008318f
C665 B.n625 VSUBS 0.008318f
C666 B.n626 VSUBS 0.008318f
C667 B.n627 VSUBS 0.008318f
C668 B.n628 VSUBS 0.008318f
C669 B.n629 VSUBS 0.008318f
C670 B.n630 VSUBS 0.008318f
C671 B.n631 VSUBS 0.008318f
C672 B.n632 VSUBS 0.008318f
C673 B.n633 VSUBS 0.008318f
C674 B.n634 VSUBS 0.008318f
C675 B.n635 VSUBS 0.008318f
C676 B.n636 VSUBS 0.008318f
C677 B.n637 VSUBS 0.008318f
C678 B.n638 VSUBS 0.008318f
C679 B.n639 VSUBS 0.008318f
C680 B.n640 VSUBS 0.008318f
C681 B.n641 VSUBS 0.008318f
C682 B.n642 VSUBS 0.008318f
C683 B.n643 VSUBS 0.008318f
C684 B.n644 VSUBS 0.008318f
C685 B.n645 VSUBS 0.008318f
C686 B.n646 VSUBS 0.008318f
C687 B.n647 VSUBS 0.008318f
C688 B.n648 VSUBS 0.008318f
C689 B.n649 VSUBS 0.008318f
C690 B.n650 VSUBS 0.008318f
C691 B.n651 VSUBS 0.008318f
C692 B.n652 VSUBS 0.008318f
C693 B.n653 VSUBS 0.008318f
C694 B.n654 VSUBS 0.008318f
C695 B.n655 VSUBS 0.008318f
C696 B.n656 VSUBS 0.008318f
C697 B.n657 VSUBS 0.008318f
C698 B.n658 VSUBS 0.008318f
C699 B.n659 VSUBS 0.008318f
C700 B.n660 VSUBS 0.008318f
C701 B.n661 VSUBS 0.008318f
C702 B.n662 VSUBS 0.008318f
C703 B.n663 VSUBS 0.008318f
C704 B.n664 VSUBS 0.008318f
C705 B.n665 VSUBS 0.008318f
C706 B.n666 VSUBS 0.008318f
C707 B.n667 VSUBS 0.008318f
C708 B.n668 VSUBS 0.008318f
C709 B.n669 VSUBS 0.008318f
C710 B.n670 VSUBS 0.008318f
C711 B.n671 VSUBS 0.008318f
C712 B.n672 VSUBS 0.008318f
C713 B.n673 VSUBS 0.008318f
C714 B.n674 VSUBS 0.008318f
C715 B.n675 VSUBS 0.008318f
C716 B.n676 VSUBS 0.008318f
C717 B.n677 VSUBS 0.008318f
C718 B.n678 VSUBS 0.008318f
C719 B.n679 VSUBS 0.008318f
C720 B.n680 VSUBS 0.008318f
C721 B.n681 VSUBS 0.008318f
C722 B.n682 VSUBS 0.008318f
C723 B.n683 VSUBS 0.008318f
C724 B.n684 VSUBS 0.008318f
C725 B.n685 VSUBS 0.008318f
C726 B.n686 VSUBS 0.005749f
C727 B.n687 VSUBS 0.019272f
C728 B.n688 VSUBS 0.006728f
C729 B.n689 VSUBS 0.008318f
C730 B.n690 VSUBS 0.008318f
C731 B.n691 VSUBS 0.008318f
C732 B.n692 VSUBS 0.008318f
C733 B.n693 VSUBS 0.008318f
C734 B.n694 VSUBS 0.008318f
C735 B.n695 VSUBS 0.008318f
C736 B.n696 VSUBS 0.008318f
C737 B.n697 VSUBS 0.008318f
C738 B.n698 VSUBS 0.008318f
C739 B.n699 VSUBS 0.008318f
C740 B.n700 VSUBS 0.006728f
C741 B.n701 VSUBS 0.008318f
C742 B.n702 VSUBS 0.008318f
C743 B.n703 VSUBS 0.005749f
C744 B.n704 VSUBS 0.008318f
C745 B.n705 VSUBS 0.008318f
C746 B.n706 VSUBS 0.008318f
C747 B.n707 VSUBS 0.008318f
C748 B.n708 VSUBS 0.008318f
C749 B.n709 VSUBS 0.008318f
C750 B.n710 VSUBS 0.008318f
C751 B.n711 VSUBS 0.008318f
C752 B.n712 VSUBS 0.008318f
C753 B.n713 VSUBS 0.008318f
C754 B.n714 VSUBS 0.008318f
C755 B.n715 VSUBS 0.008318f
C756 B.n716 VSUBS 0.008318f
C757 B.n717 VSUBS 0.008318f
C758 B.n718 VSUBS 0.008318f
C759 B.n719 VSUBS 0.008318f
C760 B.n720 VSUBS 0.008318f
C761 B.n721 VSUBS 0.008318f
C762 B.n722 VSUBS 0.008318f
C763 B.n723 VSUBS 0.008318f
C764 B.n724 VSUBS 0.008318f
C765 B.n725 VSUBS 0.008318f
C766 B.n726 VSUBS 0.008318f
C767 B.n727 VSUBS 0.008318f
C768 B.n728 VSUBS 0.008318f
C769 B.n729 VSUBS 0.008318f
C770 B.n730 VSUBS 0.008318f
C771 B.n731 VSUBS 0.008318f
C772 B.n732 VSUBS 0.008318f
C773 B.n733 VSUBS 0.008318f
C774 B.n734 VSUBS 0.008318f
C775 B.n735 VSUBS 0.008318f
C776 B.n736 VSUBS 0.008318f
C777 B.n737 VSUBS 0.008318f
C778 B.n738 VSUBS 0.008318f
C779 B.n739 VSUBS 0.008318f
C780 B.n740 VSUBS 0.008318f
C781 B.n741 VSUBS 0.008318f
C782 B.n742 VSUBS 0.008318f
C783 B.n743 VSUBS 0.008318f
C784 B.n744 VSUBS 0.008318f
C785 B.n745 VSUBS 0.008318f
C786 B.n746 VSUBS 0.008318f
C787 B.n747 VSUBS 0.008318f
C788 B.n748 VSUBS 0.008318f
C789 B.n749 VSUBS 0.008318f
C790 B.n750 VSUBS 0.008318f
C791 B.n751 VSUBS 0.008318f
C792 B.n752 VSUBS 0.008318f
C793 B.n753 VSUBS 0.008318f
C794 B.n754 VSUBS 0.008318f
C795 B.n755 VSUBS 0.008318f
C796 B.n756 VSUBS 0.008318f
C797 B.n757 VSUBS 0.008318f
C798 B.n758 VSUBS 0.008318f
C799 B.n759 VSUBS 0.008318f
C800 B.n760 VSUBS 0.008318f
C801 B.n761 VSUBS 0.008318f
C802 B.n762 VSUBS 0.008318f
C803 B.n763 VSUBS 0.008318f
C804 B.n764 VSUBS 0.008318f
C805 B.n765 VSUBS 0.008318f
C806 B.n766 VSUBS 0.008318f
C807 B.n767 VSUBS 0.008318f
C808 B.n768 VSUBS 0.008318f
C809 B.n769 VSUBS 0.008318f
C810 B.n770 VSUBS 0.008318f
C811 B.n771 VSUBS 0.008318f
C812 B.n772 VSUBS 0.008318f
C813 B.n773 VSUBS 0.008318f
C814 B.n774 VSUBS 0.008318f
C815 B.n775 VSUBS 0.008318f
C816 B.n776 VSUBS 0.008318f
C817 B.n777 VSUBS 0.008318f
C818 B.n778 VSUBS 0.008318f
C819 B.n779 VSUBS 0.008318f
C820 B.n780 VSUBS 0.008318f
C821 B.n781 VSUBS 0.008318f
C822 B.n782 VSUBS 0.008318f
C823 B.n783 VSUBS 0.008318f
C824 B.n784 VSUBS 0.008318f
C825 B.n785 VSUBS 0.008318f
C826 B.n786 VSUBS 0.008318f
C827 B.n787 VSUBS 0.008318f
C828 B.n788 VSUBS 0.008318f
C829 B.n789 VSUBS 0.008318f
C830 B.n790 VSUBS 0.008318f
C831 B.n791 VSUBS 0.008318f
C832 B.n792 VSUBS 0.008318f
C833 B.n793 VSUBS 0.008318f
C834 B.n794 VSUBS 0.008318f
C835 B.n795 VSUBS 0.008318f
C836 B.n796 VSUBS 0.008318f
C837 B.n797 VSUBS 0.008318f
C838 B.n798 VSUBS 0.019288f
C839 B.n799 VSUBS 0.019288f
C840 B.n800 VSUBS 0.018142f
C841 B.n801 VSUBS 0.008318f
C842 B.n802 VSUBS 0.008318f
C843 B.n803 VSUBS 0.008318f
C844 B.n804 VSUBS 0.008318f
C845 B.n805 VSUBS 0.008318f
C846 B.n806 VSUBS 0.008318f
C847 B.n807 VSUBS 0.008318f
C848 B.n808 VSUBS 0.008318f
C849 B.n809 VSUBS 0.008318f
C850 B.n810 VSUBS 0.008318f
C851 B.n811 VSUBS 0.008318f
C852 B.n812 VSUBS 0.008318f
C853 B.n813 VSUBS 0.008318f
C854 B.n814 VSUBS 0.008318f
C855 B.n815 VSUBS 0.008318f
C856 B.n816 VSUBS 0.008318f
C857 B.n817 VSUBS 0.008318f
C858 B.n818 VSUBS 0.008318f
C859 B.n819 VSUBS 0.008318f
C860 B.n820 VSUBS 0.008318f
C861 B.n821 VSUBS 0.008318f
C862 B.n822 VSUBS 0.008318f
C863 B.n823 VSUBS 0.008318f
C864 B.n824 VSUBS 0.008318f
C865 B.n825 VSUBS 0.008318f
C866 B.n826 VSUBS 0.008318f
C867 B.n827 VSUBS 0.008318f
C868 B.n828 VSUBS 0.008318f
C869 B.n829 VSUBS 0.008318f
C870 B.n830 VSUBS 0.008318f
C871 B.n831 VSUBS 0.008318f
C872 B.n832 VSUBS 0.008318f
C873 B.n833 VSUBS 0.008318f
C874 B.n834 VSUBS 0.008318f
C875 B.n835 VSUBS 0.008318f
C876 B.n836 VSUBS 0.008318f
C877 B.n837 VSUBS 0.008318f
C878 B.n838 VSUBS 0.008318f
C879 B.n839 VSUBS 0.008318f
C880 B.n840 VSUBS 0.008318f
C881 B.n841 VSUBS 0.008318f
C882 B.n842 VSUBS 0.008318f
C883 B.n843 VSUBS 0.008318f
C884 B.n844 VSUBS 0.008318f
C885 B.n845 VSUBS 0.008318f
C886 B.n846 VSUBS 0.008318f
C887 B.n847 VSUBS 0.008318f
C888 B.n848 VSUBS 0.008318f
C889 B.n849 VSUBS 0.008318f
C890 B.n850 VSUBS 0.008318f
C891 B.n851 VSUBS 0.010854f
C892 B.n852 VSUBS 0.011563f
C893 B.n853 VSUBS 0.022994f
C894 VDD2.t3 VSUBS 4.59037f
C895 VDD2.t7 VSUBS 0.418215f
C896 VDD2.t0 VSUBS 0.418215f
C897 VDD2.n0 VSUBS 3.53348f
C898 VDD2.n1 VSUBS 1.37847f
C899 VDD2.t4 VSUBS 0.418215f
C900 VDD2.t1 VSUBS 0.418215f
C901 VDD2.n2 VSUBS 3.54308f
C902 VDD2.n3 VSUBS 3.14046f
C903 VDD2.t2 VSUBS 4.57692f
C904 VDD2.n4 VSUBS 3.72593f
C905 VDD2.t9 VSUBS 0.418215f
C906 VDD2.t8 VSUBS 0.418215f
C907 VDD2.n5 VSUBS 3.53348f
C908 VDD2.n6 VSUBS 0.662664f
C909 VDD2.t6 VSUBS 0.418215f
C910 VDD2.t5 VSUBS 0.418215f
C911 VDD2.n7 VSUBS 3.54303f
C912 VN.n0 VSUBS 0.050775f
C913 VN.t5 VSUBS 2.53389f
C914 VN.n1 VSUBS 0.894097f
C915 VN.n2 VSUBS 0.038052f
C916 VN.t9 VSUBS 2.53389f
C917 VN.n3 VSUBS 0.894097f
C918 VN.n4 VSUBS 0.038052f
C919 VN.t2 VSUBS 2.53389f
C920 VN.n5 VSUBS 0.945133f
C921 VN.t6 VSUBS 2.64872f
C922 VN.n6 VSUBS 0.956357f
C923 VN.n7 VSUBS 0.198313f
C924 VN.n8 VSUBS 0.060526f
C925 VN.n9 VSUBS 0.031069f
C926 VN.n10 VSUBS 0.058915f
C927 VN.n11 VSUBS 0.038052f
C928 VN.n12 VSUBS 0.038052f
C929 VN.n13 VSUBS 0.058915f
C930 VN.n14 VSUBS 0.031069f
C931 VN.n15 VSUBS 0.060526f
C932 VN.n16 VSUBS 0.038052f
C933 VN.n17 VSUBS 0.038052f
C934 VN.n18 VSUBS 0.055809f
C935 VN.n19 VSUBS 0.027256f
C936 VN.t8 VSUBS 2.60501f
C937 VN.n20 VSUBS 0.966243f
C938 VN.n21 VSUBS 0.035637f
C939 VN.n22 VSUBS 0.050775f
C940 VN.t0 VSUBS 2.53389f
C941 VN.n23 VSUBS 0.894097f
C942 VN.n24 VSUBS 0.038052f
C943 VN.t1 VSUBS 2.53389f
C944 VN.n25 VSUBS 0.894097f
C945 VN.n26 VSUBS 0.038052f
C946 VN.t3 VSUBS 2.53389f
C947 VN.n27 VSUBS 0.945133f
C948 VN.t4 VSUBS 2.64872f
C949 VN.n28 VSUBS 0.956357f
C950 VN.n29 VSUBS 0.198313f
C951 VN.n30 VSUBS 0.060526f
C952 VN.n31 VSUBS 0.031069f
C953 VN.n32 VSUBS 0.058915f
C954 VN.n33 VSUBS 0.038052f
C955 VN.n34 VSUBS 0.038052f
C956 VN.n35 VSUBS 0.058915f
C957 VN.n36 VSUBS 0.031069f
C958 VN.n37 VSUBS 0.060526f
C959 VN.n38 VSUBS 0.038052f
C960 VN.n39 VSUBS 0.038052f
C961 VN.n40 VSUBS 0.055809f
C962 VN.n41 VSUBS 0.027256f
C963 VN.t7 VSUBS 2.60501f
C964 VN.n42 VSUBS 0.966243f
C965 VN.n43 VSUBS 2.20786f
C966 VTAIL.t8 VSUBS 0.421574f
C967 VTAIL.t9 VSUBS 0.421574f
C968 VTAIL.n0 VSUBS 3.40217f
C969 VTAIL.n1 VSUBS 0.831852f
C970 VTAIL.t11 VSUBS 4.42915f
C971 VTAIL.n2 VSUBS 0.978554f
C972 VTAIL.t12 VSUBS 0.421574f
C973 VTAIL.t17 VSUBS 0.421574f
C974 VTAIL.n3 VSUBS 3.40217f
C975 VTAIL.n4 VSUBS 0.872995f
C976 VTAIL.t13 VSUBS 0.421574f
C977 VTAIL.t19 VSUBS 0.421574f
C978 VTAIL.n5 VSUBS 3.40217f
C979 VTAIL.n6 VSUBS 2.83665f
C980 VTAIL.t2 VSUBS 0.421574f
C981 VTAIL.t7 VSUBS 0.421574f
C982 VTAIL.n7 VSUBS 3.40216f
C983 VTAIL.n8 VSUBS 2.83665f
C984 VTAIL.t1 VSUBS 0.421574f
C985 VTAIL.t0 VSUBS 0.421574f
C986 VTAIL.n9 VSUBS 3.40216f
C987 VTAIL.n10 VSUBS 0.872994f
C988 VTAIL.t3 VSUBS 4.42915f
C989 VTAIL.n11 VSUBS 0.978553f
C990 VTAIL.t14 VSUBS 0.421574f
C991 VTAIL.t16 VSUBS 0.421574f
C992 VTAIL.n12 VSUBS 3.40216f
C993 VTAIL.n13 VSUBS 0.855789f
C994 VTAIL.t15 VSUBS 0.421574f
C995 VTAIL.t18 VSUBS 0.421574f
C996 VTAIL.n14 VSUBS 3.40216f
C997 VTAIL.n15 VSUBS 0.872994f
C998 VTAIL.t10 VSUBS 4.42915f
C999 VTAIL.n16 VSUBS 2.84347f
C1000 VTAIL.t5 VSUBS 4.42915f
C1001 VTAIL.n17 VSUBS 2.84347f
C1002 VTAIL.t6 VSUBS 0.421574f
C1003 VTAIL.t4 VSUBS 0.421574f
C1004 VTAIL.n18 VSUBS 3.40217f
C1005 VTAIL.n19 VSUBS 0.780984f
C1006 VDD1.t2 VSUBS 4.59053f
C1007 VDD1.t4 VSUBS 0.41823f
C1008 VDD1.t3 VSUBS 0.41823f
C1009 VDD1.n0 VSUBS 3.53361f
C1010 VDD1.n1 VSUBS 1.38607f
C1011 VDD1.t7 VSUBS 4.59053f
C1012 VDD1.t1 VSUBS 0.41823f
C1013 VDD1.t6 VSUBS 0.41823f
C1014 VDD1.n2 VSUBS 3.53361f
C1015 VDD1.n3 VSUBS 1.37852f
C1016 VDD1.t5 VSUBS 0.41823f
C1017 VDD1.t9 VSUBS 0.41823f
C1018 VDD1.n4 VSUBS 3.54321f
C1019 VDD1.n5 VSUBS 3.23918f
C1020 VDD1.t0 VSUBS 0.41823f
C1021 VDD1.t8 VSUBS 0.41823f
C1022 VDD1.n6 VSUBS 3.5336f
C1023 VDD1.n7 VSUBS 3.71026f
C1024 VP.n0 VSUBS 0.051581f
C1025 VP.t2 VSUBS 2.57413f
C1026 VP.n1 VSUBS 0.908298f
C1027 VP.n2 VSUBS 0.038656f
C1028 VP.t7 VSUBS 2.57413f
C1029 VP.n3 VSUBS 0.908298f
C1030 VP.n4 VSUBS 0.038656f
C1031 VP.t0 VSUBS 2.57413f
C1032 VP.n5 VSUBS 0.908298f
C1033 VP.n6 VSUBS 0.051581f
C1034 VP.n7 VSUBS 0.051581f
C1035 VP.t9 VSUBS 2.64638f
C1036 VP.t1 VSUBS 2.57413f
C1037 VP.n8 VSUBS 0.908298f
C1038 VP.n9 VSUBS 0.038656f
C1039 VP.t4 VSUBS 2.57413f
C1040 VP.n10 VSUBS 0.908298f
C1041 VP.n11 VSUBS 0.038656f
C1042 VP.t3 VSUBS 2.57413f
C1043 VP.n12 VSUBS 0.960144f
C1044 VP.t5 VSUBS 2.69079f
C1045 VP.n13 VSUBS 0.971546f
C1046 VP.n14 VSUBS 0.201463f
C1047 VP.n15 VSUBS 0.061488f
C1048 VP.n16 VSUBS 0.031563f
C1049 VP.n17 VSUBS 0.059851f
C1050 VP.n18 VSUBS 0.038656f
C1051 VP.n19 VSUBS 0.038656f
C1052 VP.n20 VSUBS 0.059851f
C1053 VP.n21 VSUBS 0.031563f
C1054 VP.n22 VSUBS 0.061488f
C1055 VP.n23 VSUBS 0.038656f
C1056 VP.n24 VSUBS 0.038656f
C1057 VP.n25 VSUBS 0.056696f
C1058 VP.n26 VSUBS 0.027689f
C1059 VP.n27 VSUBS 0.981589f
C1060 VP.n28 VSUBS 2.22195f
C1061 VP.n29 VSUBS 2.24884f
C1062 VP.t6 VSUBS 2.64638f
C1063 VP.n30 VSUBS 0.981589f
C1064 VP.n31 VSUBS 0.027689f
C1065 VP.n32 VSUBS 0.056696f
C1066 VP.n33 VSUBS 0.038656f
C1067 VP.n34 VSUBS 0.038656f
C1068 VP.n35 VSUBS 0.061488f
C1069 VP.n36 VSUBS 0.031563f
C1070 VP.n37 VSUBS 0.059851f
C1071 VP.n38 VSUBS 0.038656f
C1072 VP.n39 VSUBS 0.038656f
C1073 VP.n40 VSUBS 0.059851f
C1074 VP.n41 VSUBS 0.031563f
C1075 VP.n42 VSUBS 0.061488f
C1076 VP.n43 VSUBS 0.038656f
C1077 VP.n44 VSUBS 0.038656f
C1078 VP.n45 VSUBS 0.056696f
C1079 VP.n46 VSUBS 0.027689f
C1080 VP.t8 VSUBS 2.64638f
C1081 VP.n47 VSUBS 0.981589f
C1082 VP.n48 VSUBS 0.036203f
.ends

