* NGSPICE file created from diff_pair_sample_0456.ext - technology: sky130A

.subckt diff_pair_sample_0456 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.2893 pd=12.52 as=0.96855 ps=6.2 w=5.87 l=3.78
X1 VDD1.t3 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.96855 pd=6.2 as=2.2893 ps=12.52 w=5.87 l=3.78
X2 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=2.2893 pd=12.52 as=0 ps=0 w=5.87 l=3.78
X3 VTAIL.t1 VP.t1 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2893 pd=12.52 as=0.96855 ps=6.2 w=5.87 l=3.78
X4 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=2.2893 pd=12.52 as=0 ps=0 w=5.87 l=3.78
X5 VDD2.t3 VN.t1 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=0.96855 pd=6.2 as=2.2893 ps=12.52 w=5.87 l=3.78
X6 VTAIL.t2 VP.t2 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.2893 pd=12.52 as=0.96855 ps=6.2 w=5.87 l=3.78
X7 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.2893 pd=12.52 as=0 ps=0 w=5.87 l=3.78
X8 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.2893 pd=12.52 as=0 ps=0 w=5.87 l=3.78
X9 VDD2.t2 VN.t2 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=0.96855 pd=6.2 as=2.2893 ps=12.52 w=5.87 l=3.78
X10 VTAIL.t4 VN.t3 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2893 pd=12.52 as=0.96855 ps=6.2 w=5.87 l=3.78
X11 VDD1.t0 VP.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.96855 pd=6.2 as=2.2893 ps=12.52 w=5.87 l=3.78
R0 VN.n1 VN.t2 71.241
R1 VN.n0 VN.t3 71.241
R2 VN.n1 VN.t0 69.8958
R3 VN.n0 VN.t1 69.8958
R4 VN VN.n1 47.3617
R5 VN VN.n0 1.87307
R6 VDD2.n2 VDD2.n0 110.24
R7 VDD2.n2 VDD2.n1 70.8347
R8 VDD2.n1 VDD2.t0 3.37358
R9 VDD2.n1 VDD2.t2 3.37358
R10 VDD2.n0 VDD2.t1 3.37358
R11 VDD2.n0 VDD2.t3 3.37358
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n238 VTAIL.n237 289.615
R14 VTAIL.n28 VTAIL.n27 289.615
R15 VTAIL.n58 VTAIL.n57 289.615
R16 VTAIL.n88 VTAIL.n87 289.615
R17 VTAIL.n208 VTAIL.n207 289.615
R18 VTAIL.n178 VTAIL.n177 289.615
R19 VTAIL.n148 VTAIL.n147 289.615
R20 VTAIL.n118 VTAIL.n117 289.615
R21 VTAIL.n221 VTAIL.n220 185
R22 VTAIL.n223 VTAIL.n222 185
R23 VTAIL.n216 VTAIL.n215 185
R24 VTAIL.n229 VTAIL.n228 185
R25 VTAIL.n231 VTAIL.n230 185
R26 VTAIL.n212 VTAIL.n211 185
R27 VTAIL.n237 VTAIL.n236 185
R28 VTAIL.n11 VTAIL.n10 185
R29 VTAIL.n13 VTAIL.n12 185
R30 VTAIL.n6 VTAIL.n5 185
R31 VTAIL.n19 VTAIL.n18 185
R32 VTAIL.n21 VTAIL.n20 185
R33 VTAIL.n2 VTAIL.n1 185
R34 VTAIL.n27 VTAIL.n26 185
R35 VTAIL.n41 VTAIL.n40 185
R36 VTAIL.n43 VTAIL.n42 185
R37 VTAIL.n36 VTAIL.n35 185
R38 VTAIL.n49 VTAIL.n48 185
R39 VTAIL.n51 VTAIL.n50 185
R40 VTAIL.n32 VTAIL.n31 185
R41 VTAIL.n57 VTAIL.n56 185
R42 VTAIL.n71 VTAIL.n70 185
R43 VTAIL.n73 VTAIL.n72 185
R44 VTAIL.n66 VTAIL.n65 185
R45 VTAIL.n79 VTAIL.n78 185
R46 VTAIL.n81 VTAIL.n80 185
R47 VTAIL.n62 VTAIL.n61 185
R48 VTAIL.n87 VTAIL.n86 185
R49 VTAIL.n207 VTAIL.n206 185
R50 VTAIL.n182 VTAIL.n181 185
R51 VTAIL.n201 VTAIL.n200 185
R52 VTAIL.n199 VTAIL.n198 185
R53 VTAIL.n186 VTAIL.n185 185
R54 VTAIL.n193 VTAIL.n192 185
R55 VTAIL.n191 VTAIL.n190 185
R56 VTAIL.n177 VTAIL.n176 185
R57 VTAIL.n152 VTAIL.n151 185
R58 VTAIL.n171 VTAIL.n170 185
R59 VTAIL.n169 VTAIL.n168 185
R60 VTAIL.n156 VTAIL.n155 185
R61 VTAIL.n163 VTAIL.n162 185
R62 VTAIL.n161 VTAIL.n160 185
R63 VTAIL.n147 VTAIL.n146 185
R64 VTAIL.n122 VTAIL.n121 185
R65 VTAIL.n141 VTAIL.n140 185
R66 VTAIL.n139 VTAIL.n138 185
R67 VTAIL.n126 VTAIL.n125 185
R68 VTAIL.n133 VTAIL.n132 185
R69 VTAIL.n131 VTAIL.n130 185
R70 VTAIL.n117 VTAIL.n116 185
R71 VTAIL.n92 VTAIL.n91 185
R72 VTAIL.n111 VTAIL.n110 185
R73 VTAIL.n109 VTAIL.n108 185
R74 VTAIL.n96 VTAIL.n95 185
R75 VTAIL.n103 VTAIL.n102 185
R76 VTAIL.n101 VTAIL.n100 185
R77 VTAIL.n219 VTAIL.t6 149.528
R78 VTAIL.n9 VTAIL.t4 149.528
R79 VTAIL.n39 VTAIL.t0 149.528
R80 VTAIL.n69 VTAIL.t2 149.528
R81 VTAIL.n189 VTAIL.t3 149.528
R82 VTAIL.n159 VTAIL.t1 149.528
R83 VTAIL.n129 VTAIL.t5 149.528
R84 VTAIL.n99 VTAIL.t7 149.528
R85 VTAIL.n222 VTAIL.n221 104.615
R86 VTAIL.n222 VTAIL.n215 104.615
R87 VTAIL.n229 VTAIL.n215 104.615
R88 VTAIL.n230 VTAIL.n229 104.615
R89 VTAIL.n230 VTAIL.n211 104.615
R90 VTAIL.n237 VTAIL.n211 104.615
R91 VTAIL.n12 VTAIL.n11 104.615
R92 VTAIL.n12 VTAIL.n5 104.615
R93 VTAIL.n19 VTAIL.n5 104.615
R94 VTAIL.n20 VTAIL.n19 104.615
R95 VTAIL.n20 VTAIL.n1 104.615
R96 VTAIL.n27 VTAIL.n1 104.615
R97 VTAIL.n42 VTAIL.n41 104.615
R98 VTAIL.n42 VTAIL.n35 104.615
R99 VTAIL.n49 VTAIL.n35 104.615
R100 VTAIL.n50 VTAIL.n49 104.615
R101 VTAIL.n50 VTAIL.n31 104.615
R102 VTAIL.n57 VTAIL.n31 104.615
R103 VTAIL.n72 VTAIL.n71 104.615
R104 VTAIL.n72 VTAIL.n65 104.615
R105 VTAIL.n79 VTAIL.n65 104.615
R106 VTAIL.n80 VTAIL.n79 104.615
R107 VTAIL.n80 VTAIL.n61 104.615
R108 VTAIL.n87 VTAIL.n61 104.615
R109 VTAIL.n207 VTAIL.n181 104.615
R110 VTAIL.n200 VTAIL.n181 104.615
R111 VTAIL.n200 VTAIL.n199 104.615
R112 VTAIL.n199 VTAIL.n185 104.615
R113 VTAIL.n192 VTAIL.n185 104.615
R114 VTAIL.n192 VTAIL.n191 104.615
R115 VTAIL.n177 VTAIL.n151 104.615
R116 VTAIL.n170 VTAIL.n151 104.615
R117 VTAIL.n170 VTAIL.n169 104.615
R118 VTAIL.n169 VTAIL.n155 104.615
R119 VTAIL.n162 VTAIL.n155 104.615
R120 VTAIL.n162 VTAIL.n161 104.615
R121 VTAIL.n147 VTAIL.n121 104.615
R122 VTAIL.n140 VTAIL.n121 104.615
R123 VTAIL.n140 VTAIL.n139 104.615
R124 VTAIL.n139 VTAIL.n125 104.615
R125 VTAIL.n132 VTAIL.n125 104.615
R126 VTAIL.n132 VTAIL.n131 104.615
R127 VTAIL.n117 VTAIL.n91 104.615
R128 VTAIL.n110 VTAIL.n91 104.615
R129 VTAIL.n110 VTAIL.n109 104.615
R130 VTAIL.n109 VTAIL.n95 104.615
R131 VTAIL.n102 VTAIL.n95 104.615
R132 VTAIL.n102 VTAIL.n101 104.615
R133 VTAIL.n221 VTAIL.t6 52.3082
R134 VTAIL.n11 VTAIL.t4 52.3082
R135 VTAIL.n41 VTAIL.t0 52.3082
R136 VTAIL.n71 VTAIL.t2 52.3082
R137 VTAIL.n191 VTAIL.t3 52.3082
R138 VTAIL.n161 VTAIL.t1 52.3082
R139 VTAIL.n131 VTAIL.t5 52.3082
R140 VTAIL.n101 VTAIL.t7 52.3082
R141 VTAIL.n239 VTAIL.n238 35.4823
R142 VTAIL.n29 VTAIL.n28 35.4823
R143 VTAIL.n59 VTAIL.n58 35.4823
R144 VTAIL.n89 VTAIL.n88 35.4823
R145 VTAIL.n209 VTAIL.n208 35.4823
R146 VTAIL.n179 VTAIL.n178 35.4823
R147 VTAIL.n149 VTAIL.n148 35.4823
R148 VTAIL.n119 VTAIL.n118 35.4823
R149 VTAIL.n239 VTAIL.n209 20.9703
R150 VTAIL.n119 VTAIL.n89 20.9703
R151 VTAIL.n236 VTAIL.n210 12.0247
R152 VTAIL.n26 VTAIL.n0 12.0247
R153 VTAIL.n56 VTAIL.n30 12.0247
R154 VTAIL.n86 VTAIL.n60 12.0247
R155 VTAIL.n206 VTAIL.n180 12.0247
R156 VTAIL.n176 VTAIL.n150 12.0247
R157 VTAIL.n146 VTAIL.n120 12.0247
R158 VTAIL.n116 VTAIL.n90 12.0247
R159 VTAIL.n235 VTAIL.n212 11.249
R160 VTAIL.n25 VTAIL.n2 11.249
R161 VTAIL.n55 VTAIL.n32 11.249
R162 VTAIL.n85 VTAIL.n62 11.249
R163 VTAIL.n205 VTAIL.n182 11.249
R164 VTAIL.n175 VTAIL.n152 11.249
R165 VTAIL.n145 VTAIL.n122 11.249
R166 VTAIL.n115 VTAIL.n92 11.249
R167 VTAIL.n232 VTAIL.n231 10.4732
R168 VTAIL.n22 VTAIL.n21 10.4732
R169 VTAIL.n52 VTAIL.n51 10.4732
R170 VTAIL.n82 VTAIL.n81 10.4732
R171 VTAIL.n202 VTAIL.n201 10.4732
R172 VTAIL.n172 VTAIL.n171 10.4732
R173 VTAIL.n142 VTAIL.n141 10.4732
R174 VTAIL.n112 VTAIL.n111 10.4732
R175 VTAIL.n220 VTAIL.n219 10.2745
R176 VTAIL.n10 VTAIL.n9 10.2745
R177 VTAIL.n40 VTAIL.n39 10.2745
R178 VTAIL.n70 VTAIL.n69 10.2745
R179 VTAIL.n190 VTAIL.n189 10.2745
R180 VTAIL.n160 VTAIL.n159 10.2745
R181 VTAIL.n130 VTAIL.n129 10.2745
R182 VTAIL.n100 VTAIL.n99 10.2745
R183 VTAIL.n228 VTAIL.n214 9.69747
R184 VTAIL.n18 VTAIL.n4 9.69747
R185 VTAIL.n48 VTAIL.n34 9.69747
R186 VTAIL.n78 VTAIL.n64 9.69747
R187 VTAIL.n198 VTAIL.n184 9.69747
R188 VTAIL.n168 VTAIL.n154 9.69747
R189 VTAIL.n138 VTAIL.n124 9.69747
R190 VTAIL.n108 VTAIL.n94 9.69747
R191 VTAIL.n234 VTAIL.n210 9.45567
R192 VTAIL.n24 VTAIL.n0 9.45567
R193 VTAIL.n54 VTAIL.n30 9.45567
R194 VTAIL.n84 VTAIL.n60 9.45567
R195 VTAIL.n204 VTAIL.n180 9.45567
R196 VTAIL.n174 VTAIL.n150 9.45567
R197 VTAIL.n144 VTAIL.n120 9.45567
R198 VTAIL.n114 VTAIL.n90 9.45567
R199 VTAIL.n218 VTAIL.n217 9.3005
R200 VTAIL.n225 VTAIL.n224 9.3005
R201 VTAIL.n227 VTAIL.n226 9.3005
R202 VTAIL.n214 VTAIL.n213 9.3005
R203 VTAIL.n233 VTAIL.n232 9.3005
R204 VTAIL.n235 VTAIL.n234 9.3005
R205 VTAIL.n8 VTAIL.n7 9.3005
R206 VTAIL.n15 VTAIL.n14 9.3005
R207 VTAIL.n17 VTAIL.n16 9.3005
R208 VTAIL.n4 VTAIL.n3 9.3005
R209 VTAIL.n23 VTAIL.n22 9.3005
R210 VTAIL.n25 VTAIL.n24 9.3005
R211 VTAIL.n38 VTAIL.n37 9.3005
R212 VTAIL.n45 VTAIL.n44 9.3005
R213 VTAIL.n47 VTAIL.n46 9.3005
R214 VTAIL.n34 VTAIL.n33 9.3005
R215 VTAIL.n53 VTAIL.n52 9.3005
R216 VTAIL.n55 VTAIL.n54 9.3005
R217 VTAIL.n68 VTAIL.n67 9.3005
R218 VTAIL.n75 VTAIL.n74 9.3005
R219 VTAIL.n77 VTAIL.n76 9.3005
R220 VTAIL.n64 VTAIL.n63 9.3005
R221 VTAIL.n83 VTAIL.n82 9.3005
R222 VTAIL.n85 VTAIL.n84 9.3005
R223 VTAIL.n205 VTAIL.n204 9.3005
R224 VTAIL.n203 VTAIL.n202 9.3005
R225 VTAIL.n184 VTAIL.n183 9.3005
R226 VTAIL.n197 VTAIL.n196 9.3005
R227 VTAIL.n195 VTAIL.n194 9.3005
R228 VTAIL.n188 VTAIL.n187 9.3005
R229 VTAIL.n165 VTAIL.n164 9.3005
R230 VTAIL.n167 VTAIL.n166 9.3005
R231 VTAIL.n154 VTAIL.n153 9.3005
R232 VTAIL.n173 VTAIL.n172 9.3005
R233 VTAIL.n175 VTAIL.n174 9.3005
R234 VTAIL.n158 VTAIL.n157 9.3005
R235 VTAIL.n135 VTAIL.n134 9.3005
R236 VTAIL.n137 VTAIL.n136 9.3005
R237 VTAIL.n124 VTAIL.n123 9.3005
R238 VTAIL.n143 VTAIL.n142 9.3005
R239 VTAIL.n145 VTAIL.n144 9.3005
R240 VTAIL.n128 VTAIL.n127 9.3005
R241 VTAIL.n105 VTAIL.n104 9.3005
R242 VTAIL.n107 VTAIL.n106 9.3005
R243 VTAIL.n94 VTAIL.n93 9.3005
R244 VTAIL.n113 VTAIL.n112 9.3005
R245 VTAIL.n115 VTAIL.n114 9.3005
R246 VTAIL.n98 VTAIL.n97 9.3005
R247 VTAIL.n227 VTAIL.n216 8.92171
R248 VTAIL.n17 VTAIL.n6 8.92171
R249 VTAIL.n47 VTAIL.n36 8.92171
R250 VTAIL.n77 VTAIL.n66 8.92171
R251 VTAIL.n197 VTAIL.n186 8.92171
R252 VTAIL.n167 VTAIL.n156 8.92171
R253 VTAIL.n137 VTAIL.n126 8.92171
R254 VTAIL.n107 VTAIL.n96 8.92171
R255 VTAIL.n224 VTAIL.n223 8.14595
R256 VTAIL.n14 VTAIL.n13 8.14595
R257 VTAIL.n44 VTAIL.n43 8.14595
R258 VTAIL.n74 VTAIL.n73 8.14595
R259 VTAIL.n194 VTAIL.n193 8.14595
R260 VTAIL.n164 VTAIL.n163 8.14595
R261 VTAIL.n134 VTAIL.n133 8.14595
R262 VTAIL.n104 VTAIL.n103 8.14595
R263 VTAIL.n220 VTAIL.n218 7.3702
R264 VTAIL.n10 VTAIL.n8 7.3702
R265 VTAIL.n40 VTAIL.n38 7.3702
R266 VTAIL.n70 VTAIL.n68 7.3702
R267 VTAIL.n190 VTAIL.n188 7.3702
R268 VTAIL.n160 VTAIL.n158 7.3702
R269 VTAIL.n130 VTAIL.n128 7.3702
R270 VTAIL.n100 VTAIL.n98 7.3702
R271 VTAIL.n223 VTAIL.n218 5.81868
R272 VTAIL.n13 VTAIL.n8 5.81868
R273 VTAIL.n43 VTAIL.n38 5.81868
R274 VTAIL.n73 VTAIL.n68 5.81868
R275 VTAIL.n193 VTAIL.n188 5.81868
R276 VTAIL.n163 VTAIL.n158 5.81868
R277 VTAIL.n133 VTAIL.n128 5.81868
R278 VTAIL.n103 VTAIL.n98 5.81868
R279 VTAIL.n224 VTAIL.n216 5.04292
R280 VTAIL.n14 VTAIL.n6 5.04292
R281 VTAIL.n44 VTAIL.n36 5.04292
R282 VTAIL.n74 VTAIL.n66 5.04292
R283 VTAIL.n194 VTAIL.n186 5.04292
R284 VTAIL.n164 VTAIL.n156 5.04292
R285 VTAIL.n134 VTAIL.n126 5.04292
R286 VTAIL.n104 VTAIL.n96 5.04292
R287 VTAIL.n228 VTAIL.n227 4.26717
R288 VTAIL.n18 VTAIL.n17 4.26717
R289 VTAIL.n48 VTAIL.n47 4.26717
R290 VTAIL.n78 VTAIL.n77 4.26717
R291 VTAIL.n198 VTAIL.n197 4.26717
R292 VTAIL.n168 VTAIL.n167 4.26717
R293 VTAIL.n138 VTAIL.n137 4.26717
R294 VTAIL.n108 VTAIL.n107 4.26717
R295 VTAIL.n149 VTAIL.n119 3.5436
R296 VTAIL.n209 VTAIL.n179 3.5436
R297 VTAIL.n89 VTAIL.n59 3.5436
R298 VTAIL.n231 VTAIL.n214 3.49141
R299 VTAIL.n21 VTAIL.n4 3.49141
R300 VTAIL.n51 VTAIL.n34 3.49141
R301 VTAIL.n81 VTAIL.n64 3.49141
R302 VTAIL.n201 VTAIL.n184 3.49141
R303 VTAIL.n171 VTAIL.n154 3.49141
R304 VTAIL.n141 VTAIL.n124 3.49141
R305 VTAIL.n111 VTAIL.n94 3.49141
R306 VTAIL.n189 VTAIL.n187 2.84323
R307 VTAIL.n159 VTAIL.n157 2.84323
R308 VTAIL.n129 VTAIL.n127 2.84323
R309 VTAIL.n99 VTAIL.n97 2.84323
R310 VTAIL.n219 VTAIL.n217 2.84323
R311 VTAIL.n9 VTAIL.n7 2.84323
R312 VTAIL.n39 VTAIL.n37 2.84323
R313 VTAIL.n69 VTAIL.n67 2.84323
R314 VTAIL.n232 VTAIL.n212 2.71565
R315 VTAIL.n22 VTAIL.n2 2.71565
R316 VTAIL.n52 VTAIL.n32 2.71565
R317 VTAIL.n82 VTAIL.n62 2.71565
R318 VTAIL.n202 VTAIL.n182 2.71565
R319 VTAIL.n172 VTAIL.n152 2.71565
R320 VTAIL.n142 VTAIL.n122 2.71565
R321 VTAIL.n112 VTAIL.n92 2.71565
R322 VTAIL.n236 VTAIL.n235 1.93989
R323 VTAIL.n26 VTAIL.n25 1.93989
R324 VTAIL.n56 VTAIL.n55 1.93989
R325 VTAIL.n86 VTAIL.n85 1.93989
R326 VTAIL.n206 VTAIL.n205 1.93989
R327 VTAIL.n176 VTAIL.n175 1.93989
R328 VTAIL.n146 VTAIL.n145 1.93989
R329 VTAIL.n116 VTAIL.n115 1.93989
R330 VTAIL VTAIL.n29 1.83024
R331 VTAIL VTAIL.n239 1.71386
R332 VTAIL.n238 VTAIL.n210 1.16414
R333 VTAIL.n28 VTAIL.n0 1.16414
R334 VTAIL.n58 VTAIL.n30 1.16414
R335 VTAIL.n88 VTAIL.n60 1.16414
R336 VTAIL.n208 VTAIL.n180 1.16414
R337 VTAIL.n178 VTAIL.n150 1.16414
R338 VTAIL.n148 VTAIL.n120 1.16414
R339 VTAIL.n118 VTAIL.n90 1.16414
R340 VTAIL.n179 VTAIL.n149 0.470328
R341 VTAIL.n59 VTAIL.n29 0.470328
R342 VTAIL.n225 VTAIL.n217 0.155672
R343 VTAIL.n226 VTAIL.n225 0.155672
R344 VTAIL.n226 VTAIL.n213 0.155672
R345 VTAIL.n233 VTAIL.n213 0.155672
R346 VTAIL.n234 VTAIL.n233 0.155672
R347 VTAIL.n15 VTAIL.n7 0.155672
R348 VTAIL.n16 VTAIL.n15 0.155672
R349 VTAIL.n16 VTAIL.n3 0.155672
R350 VTAIL.n23 VTAIL.n3 0.155672
R351 VTAIL.n24 VTAIL.n23 0.155672
R352 VTAIL.n45 VTAIL.n37 0.155672
R353 VTAIL.n46 VTAIL.n45 0.155672
R354 VTAIL.n46 VTAIL.n33 0.155672
R355 VTAIL.n53 VTAIL.n33 0.155672
R356 VTAIL.n54 VTAIL.n53 0.155672
R357 VTAIL.n75 VTAIL.n67 0.155672
R358 VTAIL.n76 VTAIL.n75 0.155672
R359 VTAIL.n76 VTAIL.n63 0.155672
R360 VTAIL.n83 VTAIL.n63 0.155672
R361 VTAIL.n84 VTAIL.n83 0.155672
R362 VTAIL.n204 VTAIL.n203 0.155672
R363 VTAIL.n203 VTAIL.n183 0.155672
R364 VTAIL.n196 VTAIL.n183 0.155672
R365 VTAIL.n196 VTAIL.n195 0.155672
R366 VTAIL.n195 VTAIL.n187 0.155672
R367 VTAIL.n174 VTAIL.n173 0.155672
R368 VTAIL.n173 VTAIL.n153 0.155672
R369 VTAIL.n166 VTAIL.n153 0.155672
R370 VTAIL.n166 VTAIL.n165 0.155672
R371 VTAIL.n165 VTAIL.n157 0.155672
R372 VTAIL.n144 VTAIL.n143 0.155672
R373 VTAIL.n143 VTAIL.n123 0.155672
R374 VTAIL.n136 VTAIL.n123 0.155672
R375 VTAIL.n136 VTAIL.n135 0.155672
R376 VTAIL.n135 VTAIL.n127 0.155672
R377 VTAIL.n114 VTAIL.n113 0.155672
R378 VTAIL.n113 VTAIL.n93 0.155672
R379 VTAIL.n106 VTAIL.n93 0.155672
R380 VTAIL.n106 VTAIL.n105 0.155672
R381 VTAIL.n105 VTAIL.n97 0.155672
R382 B.n653 B.n652 585
R383 B.n654 B.n653 585
R384 B.n227 B.n112 585
R385 B.n226 B.n225 585
R386 B.n224 B.n223 585
R387 B.n222 B.n221 585
R388 B.n220 B.n219 585
R389 B.n218 B.n217 585
R390 B.n216 B.n215 585
R391 B.n214 B.n213 585
R392 B.n212 B.n211 585
R393 B.n210 B.n209 585
R394 B.n208 B.n207 585
R395 B.n206 B.n205 585
R396 B.n204 B.n203 585
R397 B.n202 B.n201 585
R398 B.n200 B.n199 585
R399 B.n198 B.n197 585
R400 B.n196 B.n195 585
R401 B.n194 B.n193 585
R402 B.n192 B.n191 585
R403 B.n190 B.n189 585
R404 B.n188 B.n187 585
R405 B.n186 B.n185 585
R406 B.n184 B.n183 585
R407 B.n181 B.n180 585
R408 B.n179 B.n178 585
R409 B.n177 B.n176 585
R410 B.n175 B.n174 585
R411 B.n173 B.n172 585
R412 B.n171 B.n170 585
R413 B.n169 B.n168 585
R414 B.n167 B.n166 585
R415 B.n165 B.n164 585
R416 B.n163 B.n162 585
R417 B.n161 B.n160 585
R418 B.n159 B.n158 585
R419 B.n157 B.n156 585
R420 B.n155 B.n154 585
R421 B.n153 B.n152 585
R422 B.n151 B.n150 585
R423 B.n149 B.n148 585
R424 B.n147 B.n146 585
R425 B.n145 B.n144 585
R426 B.n143 B.n142 585
R427 B.n141 B.n140 585
R428 B.n139 B.n138 585
R429 B.n137 B.n136 585
R430 B.n135 B.n134 585
R431 B.n133 B.n132 585
R432 B.n131 B.n130 585
R433 B.n129 B.n128 585
R434 B.n127 B.n126 585
R435 B.n125 B.n124 585
R436 B.n123 B.n122 585
R437 B.n121 B.n120 585
R438 B.n119 B.n118 585
R439 B.n82 B.n81 585
R440 B.n651 B.n83 585
R441 B.n655 B.n83 585
R442 B.n650 B.n649 585
R443 B.n649 B.n79 585
R444 B.n648 B.n78 585
R445 B.n661 B.n78 585
R446 B.n647 B.n77 585
R447 B.n662 B.n77 585
R448 B.n646 B.n76 585
R449 B.n663 B.n76 585
R450 B.n645 B.n644 585
R451 B.n644 B.n72 585
R452 B.n643 B.n71 585
R453 B.n669 B.n71 585
R454 B.n642 B.n70 585
R455 B.n670 B.n70 585
R456 B.n641 B.n69 585
R457 B.n671 B.n69 585
R458 B.n640 B.n639 585
R459 B.n639 B.n68 585
R460 B.n638 B.n64 585
R461 B.n677 B.n64 585
R462 B.n637 B.n63 585
R463 B.n678 B.n63 585
R464 B.n636 B.n62 585
R465 B.n679 B.n62 585
R466 B.n635 B.n634 585
R467 B.n634 B.n58 585
R468 B.n633 B.n57 585
R469 B.n685 B.n57 585
R470 B.n632 B.n56 585
R471 B.n686 B.n56 585
R472 B.n631 B.n55 585
R473 B.n687 B.n55 585
R474 B.n630 B.n629 585
R475 B.n629 B.n51 585
R476 B.n628 B.n50 585
R477 B.n693 B.n50 585
R478 B.n627 B.n49 585
R479 B.n694 B.n49 585
R480 B.n626 B.n48 585
R481 B.n695 B.n48 585
R482 B.n625 B.n624 585
R483 B.n624 B.n44 585
R484 B.n623 B.n43 585
R485 B.n701 B.n43 585
R486 B.n622 B.n42 585
R487 B.n702 B.n42 585
R488 B.n621 B.n41 585
R489 B.n703 B.n41 585
R490 B.n620 B.n619 585
R491 B.n619 B.n37 585
R492 B.n618 B.n36 585
R493 B.n709 B.n36 585
R494 B.n617 B.n35 585
R495 B.n710 B.n35 585
R496 B.n616 B.n34 585
R497 B.n711 B.n34 585
R498 B.n615 B.n614 585
R499 B.n614 B.n30 585
R500 B.n613 B.n29 585
R501 B.n717 B.n29 585
R502 B.n612 B.n28 585
R503 B.n718 B.n28 585
R504 B.n611 B.n27 585
R505 B.n719 B.n27 585
R506 B.n610 B.n609 585
R507 B.n609 B.n23 585
R508 B.n608 B.n22 585
R509 B.n725 B.n22 585
R510 B.n607 B.n21 585
R511 B.n726 B.n21 585
R512 B.n606 B.n20 585
R513 B.n727 B.n20 585
R514 B.n605 B.n604 585
R515 B.n604 B.n16 585
R516 B.n603 B.n15 585
R517 B.n733 B.n15 585
R518 B.n602 B.n14 585
R519 B.n734 B.n14 585
R520 B.n601 B.n13 585
R521 B.n735 B.n13 585
R522 B.n600 B.n599 585
R523 B.n599 B.n12 585
R524 B.n598 B.n597 585
R525 B.n598 B.n8 585
R526 B.n596 B.n7 585
R527 B.n742 B.n7 585
R528 B.n595 B.n6 585
R529 B.n743 B.n6 585
R530 B.n594 B.n5 585
R531 B.n744 B.n5 585
R532 B.n593 B.n592 585
R533 B.n592 B.n4 585
R534 B.n591 B.n228 585
R535 B.n591 B.n590 585
R536 B.n581 B.n229 585
R537 B.n230 B.n229 585
R538 B.n583 B.n582 585
R539 B.n584 B.n583 585
R540 B.n580 B.n235 585
R541 B.n235 B.n234 585
R542 B.n579 B.n578 585
R543 B.n578 B.n577 585
R544 B.n237 B.n236 585
R545 B.n238 B.n237 585
R546 B.n570 B.n569 585
R547 B.n571 B.n570 585
R548 B.n568 B.n243 585
R549 B.n243 B.n242 585
R550 B.n567 B.n566 585
R551 B.n566 B.n565 585
R552 B.n245 B.n244 585
R553 B.n246 B.n245 585
R554 B.n558 B.n557 585
R555 B.n559 B.n558 585
R556 B.n556 B.n251 585
R557 B.n251 B.n250 585
R558 B.n555 B.n554 585
R559 B.n554 B.n553 585
R560 B.n253 B.n252 585
R561 B.n254 B.n253 585
R562 B.n546 B.n545 585
R563 B.n547 B.n546 585
R564 B.n544 B.n259 585
R565 B.n259 B.n258 585
R566 B.n543 B.n542 585
R567 B.n542 B.n541 585
R568 B.n261 B.n260 585
R569 B.n262 B.n261 585
R570 B.n534 B.n533 585
R571 B.n535 B.n534 585
R572 B.n532 B.n267 585
R573 B.n267 B.n266 585
R574 B.n531 B.n530 585
R575 B.n530 B.n529 585
R576 B.n269 B.n268 585
R577 B.n270 B.n269 585
R578 B.n522 B.n521 585
R579 B.n523 B.n522 585
R580 B.n520 B.n275 585
R581 B.n275 B.n274 585
R582 B.n519 B.n518 585
R583 B.n518 B.n517 585
R584 B.n277 B.n276 585
R585 B.n278 B.n277 585
R586 B.n510 B.n509 585
R587 B.n511 B.n510 585
R588 B.n508 B.n283 585
R589 B.n283 B.n282 585
R590 B.n507 B.n506 585
R591 B.n506 B.n505 585
R592 B.n285 B.n284 585
R593 B.n286 B.n285 585
R594 B.n498 B.n497 585
R595 B.n499 B.n498 585
R596 B.n496 B.n291 585
R597 B.n291 B.n290 585
R598 B.n495 B.n494 585
R599 B.n494 B.n493 585
R600 B.n293 B.n292 585
R601 B.n486 B.n293 585
R602 B.n485 B.n484 585
R603 B.n487 B.n485 585
R604 B.n483 B.n298 585
R605 B.n298 B.n297 585
R606 B.n482 B.n481 585
R607 B.n481 B.n480 585
R608 B.n300 B.n299 585
R609 B.n301 B.n300 585
R610 B.n473 B.n472 585
R611 B.n474 B.n473 585
R612 B.n471 B.n306 585
R613 B.n306 B.n305 585
R614 B.n470 B.n469 585
R615 B.n469 B.n468 585
R616 B.n308 B.n307 585
R617 B.n309 B.n308 585
R618 B.n461 B.n460 585
R619 B.n462 B.n461 585
R620 B.n312 B.n311 585
R621 B.n348 B.n346 585
R622 B.n349 B.n345 585
R623 B.n349 B.n313 585
R624 B.n352 B.n351 585
R625 B.n353 B.n344 585
R626 B.n355 B.n354 585
R627 B.n357 B.n343 585
R628 B.n360 B.n359 585
R629 B.n361 B.n342 585
R630 B.n363 B.n362 585
R631 B.n365 B.n341 585
R632 B.n368 B.n367 585
R633 B.n369 B.n340 585
R634 B.n371 B.n370 585
R635 B.n373 B.n339 585
R636 B.n376 B.n375 585
R637 B.n377 B.n338 585
R638 B.n379 B.n378 585
R639 B.n381 B.n337 585
R640 B.n384 B.n383 585
R641 B.n385 B.n336 585
R642 B.n387 B.n386 585
R643 B.n389 B.n335 585
R644 B.n392 B.n391 585
R645 B.n394 B.n332 585
R646 B.n396 B.n395 585
R647 B.n398 B.n331 585
R648 B.n401 B.n400 585
R649 B.n402 B.n330 585
R650 B.n404 B.n403 585
R651 B.n406 B.n329 585
R652 B.n409 B.n408 585
R653 B.n410 B.n326 585
R654 B.n413 B.n412 585
R655 B.n415 B.n325 585
R656 B.n418 B.n417 585
R657 B.n419 B.n324 585
R658 B.n421 B.n420 585
R659 B.n423 B.n323 585
R660 B.n426 B.n425 585
R661 B.n427 B.n322 585
R662 B.n429 B.n428 585
R663 B.n431 B.n321 585
R664 B.n434 B.n433 585
R665 B.n435 B.n320 585
R666 B.n437 B.n436 585
R667 B.n439 B.n319 585
R668 B.n442 B.n441 585
R669 B.n443 B.n318 585
R670 B.n445 B.n444 585
R671 B.n447 B.n317 585
R672 B.n450 B.n449 585
R673 B.n451 B.n316 585
R674 B.n453 B.n452 585
R675 B.n455 B.n315 585
R676 B.n458 B.n457 585
R677 B.n459 B.n314 585
R678 B.n464 B.n463 585
R679 B.n463 B.n462 585
R680 B.n465 B.n310 585
R681 B.n310 B.n309 585
R682 B.n467 B.n466 585
R683 B.n468 B.n467 585
R684 B.n304 B.n303 585
R685 B.n305 B.n304 585
R686 B.n476 B.n475 585
R687 B.n475 B.n474 585
R688 B.n477 B.n302 585
R689 B.n302 B.n301 585
R690 B.n479 B.n478 585
R691 B.n480 B.n479 585
R692 B.n296 B.n295 585
R693 B.n297 B.n296 585
R694 B.n489 B.n488 585
R695 B.n488 B.n487 585
R696 B.n490 B.n294 585
R697 B.n486 B.n294 585
R698 B.n492 B.n491 585
R699 B.n493 B.n492 585
R700 B.n289 B.n288 585
R701 B.n290 B.n289 585
R702 B.n501 B.n500 585
R703 B.n500 B.n499 585
R704 B.n502 B.n287 585
R705 B.n287 B.n286 585
R706 B.n504 B.n503 585
R707 B.n505 B.n504 585
R708 B.n281 B.n280 585
R709 B.n282 B.n281 585
R710 B.n513 B.n512 585
R711 B.n512 B.n511 585
R712 B.n514 B.n279 585
R713 B.n279 B.n278 585
R714 B.n516 B.n515 585
R715 B.n517 B.n516 585
R716 B.n273 B.n272 585
R717 B.n274 B.n273 585
R718 B.n525 B.n524 585
R719 B.n524 B.n523 585
R720 B.n526 B.n271 585
R721 B.n271 B.n270 585
R722 B.n528 B.n527 585
R723 B.n529 B.n528 585
R724 B.n265 B.n264 585
R725 B.n266 B.n265 585
R726 B.n537 B.n536 585
R727 B.n536 B.n535 585
R728 B.n538 B.n263 585
R729 B.n263 B.n262 585
R730 B.n540 B.n539 585
R731 B.n541 B.n540 585
R732 B.n257 B.n256 585
R733 B.n258 B.n257 585
R734 B.n549 B.n548 585
R735 B.n548 B.n547 585
R736 B.n550 B.n255 585
R737 B.n255 B.n254 585
R738 B.n552 B.n551 585
R739 B.n553 B.n552 585
R740 B.n249 B.n248 585
R741 B.n250 B.n249 585
R742 B.n561 B.n560 585
R743 B.n560 B.n559 585
R744 B.n562 B.n247 585
R745 B.n247 B.n246 585
R746 B.n564 B.n563 585
R747 B.n565 B.n564 585
R748 B.n241 B.n240 585
R749 B.n242 B.n241 585
R750 B.n573 B.n572 585
R751 B.n572 B.n571 585
R752 B.n574 B.n239 585
R753 B.n239 B.n238 585
R754 B.n576 B.n575 585
R755 B.n577 B.n576 585
R756 B.n233 B.n232 585
R757 B.n234 B.n233 585
R758 B.n586 B.n585 585
R759 B.n585 B.n584 585
R760 B.n587 B.n231 585
R761 B.n231 B.n230 585
R762 B.n589 B.n588 585
R763 B.n590 B.n589 585
R764 B.n3 B.n0 585
R765 B.n4 B.n3 585
R766 B.n741 B.n1 585
R767 B.n742 B.n741 585
R768 B.n740 B.n739 585
R769 B.n740 B.n8 585
R770 B.n738 B.n9 585
R771 B.n12 B.n9 585
R772 B.n737 B.n736 585
R773 B.n736 B.n735 585
R774 B.n11 B.n10 585
R775 B.n734 B.n11 585
R776 B.n732 B.n731 585
R777 B.n733 B.n732 585
R778 B.n730 B.n17 585
R779 B.n17 B.n16 585
R780 B.n729 B.n728 585
R781 B.n728 B.n727 585
R782 B.n19 B.n18 585
R783 B.n726 B.n19 585
R784 B.n724 B.n723 585
R785 B.n725 B.n724 585
R786 B.n722 B.n24 585
R787 B.n24 B.n23 585
R788 B.n721 B.n720 585
R789 B.n720 B.n719 585
R790 B.n26 B.n25 585
R791 B.n718 B.n26 585
R792 B.n716 B.n715 585
R793 B.n717 B.n716 585
R794 B.n714 B.n31 585
R795 B.n31 B.n30 585
R796 B.n713 B.n712 585
R797 B.n712 B.n711 585
R798 B.n33 B.n32 585
R799 B.n710 B.n33 585
R800 B.n708 B.n707 585
R801 B.n709 B.n708 585
R802 B.n706 B.n38 585
R803 B.n38 B.n37 585
R804 B.n705 B.n704 585
R805 B.n704 B.n703 585
R806 B.n40 B.n39 585
R807 B.n702 B.n40 585
R808 B.n700 B.n699 585
R809 B.n701 B.n700 585
R810 B.n698 B.n45 585
R811 B.n45 B.n44 585
R812 B.n697 B.n696 585
R813 B.n696 B.n695 585
R814 B.n47 B.n46 585
R815 B.n694 B.n47 585
R816 B.n692 B.n691 585
R817 B.n693 B.n692 585
R818 B.n690 B.n52 585
R819 B.n52 B.n51 585
R820 B.n689 B.n688 585
R821 B.n688 B.n687 585
R822 B.n54 B.n53 585
R823 B.n686 B.n54 585
R824 B.n684 B.n683 585
R825 B.n685 B.n684 585
R826 B.n682 B.n59 585
R827 B.n59 B.n58 585
R828 B.n681 B.n680 585
R829 B.n680 B.n679 585
R830 B.n61 B.n60 585
R831 B.n678 B.n61 585
R832 B.n676 B.n675 585
R833 B.n677 B.n676 585
R834 B.n674 B.n65 585
R835 B.n68 B.n65 585
R836 B.n673 B.n672 585
R837 B.n672 B.n671 585
R838 B.n67 B.n66 585
R839 B.n670 B.n67 585
R840 B.n668 B.n667 585
R841 B.n669 B.n668 585
R842 B.n666 B.n73 585
R843 B.n73 B.n72 585
R844 B.n665 B.n664 585
R845 B.n664 B.n663 585
R846 B.n75 B.n74 585
R847 B.n662 B.n75 585
R848 B.n660 B.n659 585
R849 B.n661 B.n660 585
R850 B.n658 B.n80 585
R851 B.n80 B.n79 585
R852 B.n657 B.n656 585
R853 B.n656 B.n655 585
R854 B.n745 B.n744 585
R855 B.n743 B.n2 585
R856 B.n656 B.n82 458.866
R857 B.n653 B.n83 458.866
R858 B.n461 B.n314 458.866
R859 B.n463 B.n312 458.866
R860 B.n654 B.n111 256.663
R861 B.n654 B.n110 256.663
R862 B.n654 B.n109 256.663
R863 B.n654 B.n108 256.663
R864 B.n654 B.n107 256.663
R865 B.n654 B.n106 256.663
R866 B.n654 B.n105 256.663
R867 B.n654 B.n104 256.663
R868 B.n654 B.n103 256.663
R869 B.n654 B.n102 256.663
R870 B.n654 B.n101 256.663
R871 B.n654 B.n100 256.663
R872 B.n654 B.n99 256.663
R873 B.n654 B.n98 256.663
R874 B.n654 B.n97 256.663
R875 B.n654 B.n96 256.663
R876 B.n654 B.n95 256.663
R877 B.n654 B.n94 256.663
R878 B.n654 B.n93 256.663
R879 B.n654 B.n92 256.663
R880 B.n654 B.n91 256.663
R881 B.n654 B.n90 256.663
R882 B.n654 B.n89 256.663
R883 B.n654 B.n88 256.663
R884 B.n654 B.n87 256.663
R885 B.n654 B.n86 256.663
R886 B.n654 B.n85 256.663
R887 B.n654 B.n84 256.663
R888 B.n347 B.n313 256.663
R889 B.n350 B.n313 256.663
R890 B.n356 B.n313 256.663
R891 B.n358 B.n313 256.663
R892 B.n364 B.n313 256.663
R893 B.n366 B.n313 256.663
R894 B.n372 B.n313 256.663
R895 B.n374 B.n313 256.663
R896 B.n380 B.n313 256.663
R897 B.n382 B.n313 256.663
R898 B.n388 B.n313 256.663
R899 B.n390 B.n313 256.663
R900 B.n397 B.n313 256.663
R901 B.n399 B.n313 256.663
R902 B.n405 B.n313 256.663
R903 B.n407 B.n313 256.663
R904 B.n414 B.n313 256.663
R905 B.n416 B.n313 256.663
R906 B.n422 B.n313 256.663
R907 B.n424 B.n313 256.663
R908 B.n430 B.n313 256.663
R909 B.n432 B.n313 256.663
R910 B.n438 B.n313 256.663
R911 B.n440 B.n313 256.663
R912 B.n446 B.n313 256.663
R913 B.n448 B.n313 256.663
R914 B.n454 B.n313 256.663
R915 B.n456 B.n313 256.663
R916 B.n747 B.n746 256.663
R917 B.n113 B.t13 256.175
R918 B.n327 B.t11 256.175
R919 B.n115 B.t6 256.175
R920 B.n333 B.t17 256.175
R921 B.n115 B.t4 246.754
R922 B.n113 B.t12 246.754
R923 B.n327 B.t8 246.754
R924 B.n333 B.t15 246.754
R925 B.n114 B.t14 176.465
R926 B.n328 B.t10 176.465
R927 B.n116 B.t7 176.465
R928 B.n334 B.t16 176.465
R929 B.n120 B.n119 163.367
R930 B.n124 B.n123 163.367
R931 B.n128 B.n127 163.367
R932 B.n132 B.n131 163.367
R933 B.n136 B.n135 163.367
R934 B.n140 B.n139 163.367
R935 B.n144 B.n143 163.367
R936 B.n148 B.n147 163.367
R937 B.n152 B.n151 163.367
R938 B.n156 B.n155 163.367
R939 B.n160 B.n159 163.367
R940 B.n164 B.n163 163.367
R941 B.n168 B.n167 163.367
R942 B.n172 B.n171 163.367
R943 B.n176 B.n175 163.367
R944 B.n180 B.n179 163.367
R945 B.n185 B.n184 163.367
R946 B.n189 B.n188 163.367
R947 B.n193 B.n192 163.367
R948 B.n197 B.n196 163.367
R949 B.n201 B.n200 163.367
R950 B.n205 B.n204 163.367
R951 B.n209 B.n208 163.367
R952 B.n213 B.n212 163.367
R953 B.n217 B.n216 163.367
R954 B.n221 B.n220 163.367
R955 B.n225 B.n224 163.367
R956 B.n653 B.n112 163.367
R957 B.n461 B.n308 163.367
R958 B.n469 B.n308 163.367
R959 B.n469 B.n306 163.367
R960 B.n473 B.n306 163.367
R961 B.n473 B.n300 163.367
R962 B.n481 B.n300 163.367
R963 B.n481 B.n298 163.367
R964 B.n485 B.n298 163.367
R965 B.n485 B.n293 163.367
R966 B.n494 B.n293 163.367
R967 B.n494 B.n291 163.367
R968 B.n498 B.n291 163.367
R969 B.n498 B.n285 163.367
R970 B.n506 B.n285 163.367
R971 B.n506 B.n283 163.367
R972 B.n510 B.n283 163.367
R973 B.n510 B.n277 163.367
R974 B.n518 B.n277 163.367
R975 B.n518 B.n275 163.367
R976 B.n522 B.n275 163.367
R977 B.n522 B.n269 163.367
R978 B.n530 B.n269 163.367
R979 B.n530 B.n267 163.367
R980 B.n534 B.n267 163.367
R981 B.n534 B.n261 163.367
R982 B.n542 B.n261 163.367
R983 B.n542 B.n259 163.367
R984 B.n546 B.n259 163.367
R985 B.n546 B.n253 163.367
R986 B.n554 B.n253 163.367
R987 B.n554 B.n251 163.367
R988 B.n558 B.n251 163.367
R989 B.n558 B.n245 163.367
R990 B.n566 B.n245 163.367
R991 B.n566 B.n243 163.367
R992 B.n570 B.n243 163.367
R993 B.n570 B.n237 163.367
R994 B.n578 B.n237 163.367
R995 B.n578 B.n235 163.367
R996 B.n583 B.n235 163.367
R997 B.n583 B.n229 163.367
R998 B.n591 B.n229 163.367
R999 B.n592 B.n591 163.367
R1000 B.n592 B.n5 163.367
R1001 B.n6 B.n5 163.367
R1002 B.n7 B.n6 163.367
R1003 B.n598 B.n7 163.367
R1004 B.n599 B.n598 163.367
R1005 B.n599 B.n13 163.367
R1006 B.n14 B.n13 163.367
R1007 B.n15 B.n14 163.367
R1008 B.n604 B.n15 163.367
R1009 B.n604 B.n20 163.367
R1010 B.n21 B.n20 163.367
R1011 B.n22 B.n21 163.367
R1012 B.n609 B.n22 163.367
R1013 B.n609 B.n27 163.367
R1014 B.n28 B.n27 163.367
R1015 B.n29 B.n28 163.367
R1016 B.n614 B.n29 163.367
R1017 B.n614 B.n34 163.367
R1018 B.n35 B.n34 163.367
R1019 B.n36 B.n35 163.367
R1020 B.n619 B.n36 163.367
R1021 B.n619 B.n41 163.367
R1022 B.n42 B.n41 163.367
R1023 B.n43 B.n42 163.367
R1024 B.n624 B.n43 163.367
R1025 B.n624 B.n48 163.367
R1026 B.n49 B.n48 163.367
R1027 B.n50 B.n49 163.367
R1028 B.n629 B.n50 163.367
R1029 B.n629 B.n55 163.367
R1030 B.n56 B.n55 163.367
R1031 B.n57 B.n56 163.367
R1032 B.n634 B.n57 163.367
R1033 B.n634 B.n62 163.367
R1034 B.n63 B.n62 163.367
R1035 B.n64 B.n63 163.367
R1036 B.n639 B.n64 163.367
R1037 B.n639 B.n69 163.367
R1038 B.n70 B.n69 163.367
R1039 B.n71 B.n70 163.367
R1040 B.n644 B.n71 163.367
R1041 B.n644 B.n76 163.367
R1042 B.n77 B.n76 163.367
R1043 B.n78 B.n77 163.367
R1044 B.n649 B.n78 163.367
R1045 B.n649 B.n83 163.367
R1046 B.n349 B.n348 163.367
R1047 B.n351 B.n349 163.367
R1048 B.n355 B.n344 163.367
R1049 B.n359 B.n357 163.367
R1050 B.n363 B.n342 163.367
R1051 B.n367 B.n365 163.367
R1052 B.n371 B.n340 163.367
R1053 B.n375 B.n373 163.367
R1054 B.n379 B.n338 163.367
R1055 B.n383 B.n381 163.367
R1056 B.n387 B.n336 163.367
R1057 B.n391 B.n389 163.367
R1058 B.n396 B.n332 163.367
R1059 B.n400 B.n398 163.367
R1060 B.n404 B.n330 163.367
R1061 B.n408 B.n406 163.367
R1062 B.n413 B.n326 163.367
R1063 B.n417 B.n415 163.367
R1064 B.n421 B.n324 163.367
R1065 B.n425 B.n423 163.367
R1066 B.n429 B.n322 163.367
R1067 B.n433 B.n431 163.367
R1068 B.n437 B.n320 163.367
R1069 B.n441 B.n439 163.367
R1070 B.n445 B.n318 163.367
R1071 B.n449 B.n447 163.367
R1072 B.n453 B.n316 163.367
R1073 B.n457 B.n455 163.367
R1074 B.n463 B.n310 163.367
R1075 B.n467 B.n310 163.367
R1076 B.n467 B.n304 163.367
R1077 B.n475 B.n304 163.367
R1078 B.n475 B.n302 163.367
R1079 B.n479 B.n302 163.367
R1080 B.n479 B.n296 163.367
R1081 B.n488 B.n296 163.367
R1082 B.n488 B.n294 163.367
R1083 B.n492 B.n294 163.367
R1084 B.n492 B.n289 163.367
R1085 B.n500 B.n289 163.367
R1086 B.n500 B.n287 163.367
R1087 B.n504 B.n287 163.367
R1088 B.n504 B.n281 163.367
R1089 B.n512 B.n281 163.367
R1090 B.n512 B.n279 163.367
R1091 B.n516 B.n279 163.367
R1092 B.n516 B.n273 163.367
R1093 B.n524 B.n273 163.367
R1094 B.n524 B.n271 163.367
R1095 B.n528 B.n271 163.367
R1096 B.n528 B.n265 163.367
R1097 B.n536 B.n265 163.367
R1098 B.n536 B.n263 163.367
R1099 B.n540 B.n263 163.367
R1100 B.n540 B.n257 163.367
R1101 B.n548 B.n257 163.367
R1102 B.n548 B.n255 163.367
R1103 B.n552 B.n255 163.367
R1104 B.n552 B.n249 163.367
R1105 B.n560 B.n249 163.367
R1106 B.n560 B.n247 163.367
R1107 B.n564 B.n247 163.367
R1108 B.n564 B.n241 163.367
R1109 B.n572 B.n241 163.367
R1110 B.n572 B.n239 163.367
R1111 B.n576 B.n239 163.367
R1112 B.n576 B.n233 163.367
R1113 B.n585 B.n233 163.367
R1114 B.n585 B.n231 163.367
R1115 B.n589 B.n231 163.367
R1116 B.n589 B.n3 163.367
R1117 B.n745 B.n3 163.367
R1118 B.n741 B.n2 163.367
R1119 B.n741 B.n740 163.367
R1120 B.n740 B.n9 163.367
R1121 B.n736 B.n9 163.367
R1122 B.n736 B.n11 163.367
R1123 B.n732 B.n11 163.367
R1124 B.n732 B.n17 163.367
R1125 B.n728 B.n17 163.367
R1126 B.n728 B.n19 163.367
R1127 B.n724 B.n19 163.367
R1128 B.n724 B.n24 163.367
R1129 B.n720 B.n24 163.367
R1130 B.n720 B.n26 163.367
R1131 B.n716 B.n26 163.367
R1132 B.n716 B.n31 163.367
R1133 B.n712 B.n31 163.367
R1134 B.n712 B.n33 163.367
R1135 B.n708 B.n33 163.367
R1136 B.n708 B.n38 163.367
R1137 B.n704 B.n38 163.367
R1138 B.n704 B.n40 163.367
R1139 B.n700 B.n40 163.367
R1140 B.n700 B.n45 163.367
R1141 B.n696 B.n45 163.367
R1142 B.n696 B.n47 163.367
R1143 B.n692 B.n47 163.367
R1144 B.n692 B.n52 163.367
R1145 B.n688 B.n52 163.367
R1146 B.n688 B.n54 163.367
R1147 B.n684 B.n54 163.367
R1148 B.n684 B.n59 163.367
R1149 B.n680 B.n59 163.367
R1150 B.n680 B.n61 163.367
R1151 B.n676 B.n61 163.367
R1152 B.n676 B.n65 163.367
R1153 B.n672 B.n65 163.367
R1154 B.n672 B.n67 163.367
R1155 B.n668 B.n67 163.367
R1156 B.n668 B.n73 163.367
R1157 B.n664 B.n73 163.367
R1158 B.n664 B.n75 163.367
R1159 B.n660 B.n75 163.367
R1160 B.n660 B.n80 163.367
R1161 B.n656 B.n80 163.367
R1162 B.n462 B.n313 113.504
R1163 B.n655 B.n654 113.504
R1164 B.n116 B.n115 79.7096
R1165 B.n114 B.n113 79.7096
R1166 B.n328 B.n327 79.7096
R1167 B.n334 B.n333 79.7096
R1168 B.n84 B.n82 71.676
R1169 B.n120 B.n85 71.676
R1170 B.n124 B.n86 71.676
R1171 B.n128 B.n87 71.676
R1172 B.n132 B.n88 71.676
R1173 B.n136 B.n89 71.676
R1174 B.n140 B.n90 71.676
R1175 B.n144 B.n91 71.676
R1176 B.n148 B.n92 71.676
R1177 B.n152 B.n93 71.676
R1178 B.n156 B.n94 71.676
R1179 B.n160 B.n95 71.676
R1180 B.n164 B.n96 71.676
R1181 B.n168 B.n97 71.676
R1182 B.n172 B.n98 71.676
R1183 B.n176 B.n99 71.676
R1184 B.n180 B.n100 71.676
R1185 B.n185 B.n101 71.676
R1186 B.n189 B.n102 71.676
R1187 B.n193 B.n103 71.676
R1188 B.n197 B.n104 71.676
R1189 B.n201 B.n105 71.676
R1190 B.n205 B.n106 71.676
R1191 B.n209 B.n107 71.676
R1192 B.n213 B.n108 71.676
R1193 B.n217 B.n109 71.676
R1194 B.n221 B.n110 71.676
R1195 B.n225 B.n111 71.676
R1196 B.n112 B.n111 71.676
R1197 B.n224 B.n110 71.676
R1198 B.n220 B.n109 71.676
R1199 B.n216 B.n108 71.676
R1200 B.n212 B.n107 71.676
R1201 B.n208 B.n106 71.676
R1202 B.n204 B.n105 71.676
R1203 B.n200 B.n104 71.676
R1204 B.n196 B.n103 71.676
R1205 B.n192 B.n102 71.676
R1206 B.n188 B.n101 71.676
R1207 B.n184 B.n100 71.676
R1208 B.n179 B.n99 71.676
R1209 B.n175 B.n98 71.676
R1210 B.n171 B.n97 71.676
R1211 B.n167 B.n96 71.676
R1212 B.n163 B.n95 71.676
R1213 B.n159 B.n94 71.676
R1214 B.n155 B.n93 71.676
R1215 B.n151 B.n92 71.676
R1216 B.n147 B.n91 71.676
R1217 B.n143 B.n90 71.676
R1218 B.n139 B.n89 71.676
R1219 B.n135 B.n88 71.676
R1220 B.n131 B.n87 71.676
R1221 B.n127 B.n86 71.676
R1222 B.n123 B.n85 71.676
R1223 B.n119 B.n84 71.676
R1224 B.n347 B.n312 71.676
R1225 B.n351 B.n350 71.676
R1226 B.n356 B.n355 71.676
R1227 B.n359 B.n358 71.676
R1228 B.n364 B.n363 71.676
R1229 B.n367 B.n366 71.676
R1230 B.n372 B.n371 71.676
R1231 B.n375 B.n374 71.676
R1232 B.n380 B.n379 71.676
R1233 B.n383 B.n382 71.676
R1234 B.n388 B.n387 71.676
R1235 B.n391 B.n390 71.676
R1236 B.n397 B.n396 71.676
R1237 B.n400 B.n399 71.676
R1238 B.n405 B.n404 71.676
R1239 B.n408 B.n407 71.676
R1240 B.n414 B.n413 71.676
R1241 B.n417 B.n416 71.676
R1242 B.n422 B.n421 71.676
R1243 B.n425 B.n424 71.676
R1244 B.n430 B.n429 71.676
R1245 B.n433 B.n432 71.676
R1246 B.n438 B.n437 71.676
R1247 B.n441 B.n440 71.676
R1248 B.n446 B.n445 71.676
R1249 B.n449 B.n448 71.676
R1250 B.n454 B.n453 71.676
R1251 B.n457 B.n456 71.676
R1252 B.n348 B.n347 71.676
R1253 B.n350 B.n344 71.676
R1254 B.n357 B.n356 71.676
R1255 B.n358 B.n342 71.676
R1256 B.n365 B.n364 71.676
R1257 B.n366 B.n340 71.676
R1258 B.n373 B.n372 71.676
R1259 B.n374 B.n338 71.676
R1260 B.n381 B.n380 71.676
R1261 B.n382 B.n336 71.676
R1262 B.n389 B.n388 71.676
R1263 B.n390 B.n332 71.676
R1264 B.n398 B.n397 71.676
R1265 B.n399 B.n330 71.676
R1266 B.n406 B.n405 71.676
R1267 B.n407 B.n326 71.676
R1268 B.n415 B.n414 71.676
R1269 B.n416 B.n324 71.676
R1270 B.n423 B.n422 71.676
R1271 B.n424 B.n322 71.676
R1272 B.n431 B.n430 71.676
R1273 B.n432 B.n320 71.676
R1274 B.n439 B.n438 71.676
R1275 B.n440 B.n318 71.676
R1276 B.n447 B.n446 71.676
R1277 B.n448 B.n316 71.676
R1278 B.n455 B.n454 71.676
R1279 B.n456 B.n314 71.676
R1280 B.n746 B.n745 71.676
R1281 B.n746 B.n2 71.676
R1282 B.n462 B.n309 67.1158
R1283 B.n468 B.n309 67.1158
R1284 B.n468 B.n305 67.1158
R1285 B.n474 B.n305 67.1158
R1286 B.n474 B.n301 67.1158
R1287 B.n480 B.n301 67.1158
R1288 B.n480 B.n297 67.1158
R1289 B.n487 B.n297 67.1158
R1290 B.n487 B.n486 67.1158
R1291 B.n493 B.n290 67.1158
R1292 B.n499 B.n290 67.1158
R1293 B.n499 B.n286 67.1158
R1294 B.n505 B.n286 67.1158
R1295 B.n505 B.n282 67.1158
R1296 B.n511 B.n282 67.1158
R1297 B.n511 B.n278 67.1158
R1298 B.n517 B.n278 67.1158
R1299 B.n517 B.n274 67.1158
R1300 B.n523 B.n274 67.1158
R1301 B.n523 B.n270 67.1158
R1302 B.n529 B.n270 67.1158
R1303 B.n529 B.n266 67.1158
R1304 B.n535 B.n266 67.1158
R1305 B.n541 B.n262 67.1158
R1306 B.n541 B.n258 67.1158
R1307 B.n547 B.n258 67.1158
R1308 B.n547 B.n254 67.1158
R1309 B.n553 B.n254 67.1158
R1310 B.n553 B.n250 67.1158
R1311 B.n559 B.n250 67.1158
R1312 B.n559 B.n246 67.1158
R1313 B.n565 B.n246 67.1158
R1314 B.n565 B.n242 67.1158
R1315 B.n571 B.n242 67.1158
R1316 B.n577 B.n238 67.1158
R1317 B.n577 B.n234 67.1158
R1318 B.n584 B.n234 67.1158
R1319 B.n584 B.n230 67.1158
R1320 B.n590 B.n230 67.1158
R1321 B.n590 B.n4 67.1158
R1322 B.n744 B.n4 67.1158
R1323 B.n744 B.n743 67.1158
R1324 B.n743 B.n742 67.1158
R1325 B.n742 B.n8 67.1158
R1326 B.n12 B.n8 67.1158
R1327 B.n735 B.n12 67.1158
R1328 B.n735 B.n734 67.1158
R1329 B.n734 B.n733 67.1158
R1330 B.n733 B.n16 67.1158
R1331 B.n727 B.n726 67.1158
R1332 B.n726 B.n725 67.1158
R1333 B.n725 B.n23 67.1158
R1334 B.n719 B.n23 67.1158
R1335 B.n719 B.n718 67.1158
R1336 B.n718 B.n717 67.1158
R1337 B.n717 B.n30 67.1158
R1338 B.n711 B.n30 67.1158
R1339 B.n711 B.n710 67.1158
R1340 B.n710 B.n709 67.1158
R1341 B.n709 B.n37 67.1158
R1342 B.n703 B.n702 67.1158
R1343 B.n702 B.n701 67.1158
R1344 B.n701 B.n44 67.1158
R1345 B.n695 B.n44 67.1158
R1346 B.n695 B.n694 67.1158
R1347 B.n694 B.n693 67.1158
R1348 B.n693 B.n51 67.1158
R1349 B.n687 B.n51 67.1158
R1350 B.n687 B.n686 67.1158
R1351 B.n686 B.n685 67.1158
R1352 B.n685 B.n58 67.1158
R1353 B.n679 B.n58 67.1158
R1354 B.n679 B.n678 67.1158
R1355 B.n678 B.n677 67.1158
R1356 B.n671 B.n68 67.1158
R1357 B.n671 B.n670 67.1158
R1358 B.n670 B.n669 67.1158
R1359 B.n669 B.n72 67.1158
R1360 B.n663 B.n72 67.1158
R1361 B.n663 B.n662 67.1158
R1362 B.n662 B.n661 67.1158
R1363 B.n661 B.n79 67.1158
R1364 B.n655 B.n79 67.1158
R1365 B.n117 B.n116 59.5399
R1366 B.n182 B.n114 59.5399
R1367 B.n411 B.n328 59.5399
R1368 B.n393 B.n334 59.5399
R1369 B.n571 B.t0 57.2459
R1370 B.n727 B.t1 57.2459
R1371 B.n535 B.t2 51.324
R1372 B.n703 B.t3 51.324
R1373 B.n493 B.t9 35.5321
R1374 B.n677 B.t5 35.5321
R1375 B.n486 B.t9 31.5842
R1376 B.n68 B.t5 31.5842
R1377 B.n464 B.n311 29.8151
R1378 B.n460 B.n459 29.8151
R1379 B.n652 B.n651 29.8151
R1380 B.n657 B.n81 29.8151
R1381 B B.n747 18.0485
R1382 B.t2 B.n262 15.7923
R1383 B.t3 B.n37 15.7923
R1384 B.n465 B.n464 10.6151
R1385 B.n466 B.n465 10.6151
R1386 B.n466 B.n303 10.6151
R1387 B.n476 B.n303 10.6151
R1388 B.n477 B.n476 10.6151
R1389 B.n478 B.n477 10.6151
R1390 B.n478 B.n295 10.6151
R1391 B.n489 B.n295 10.6151
R1392 B.n490 B.n489 10.6151
R1393 B.n491 B.n490 10.6151
R1394 B.n491 B.n288 10.6151
R1395 B.n501 B.n288 10.6151
R1396 B.n502 B.n501 10.6151
R1397 B.n503 B.n502 10.6151
R1398 B.n503 B.n280 10.6151
R1399 B.n513 B.n280 10.6151
R1400 B.n514 B.n513 10.6151
R1401 B.n515 B.n514 10.6151
R1402 B.n515 B.n272 10.6151
R1403 B.n525 B.n272 10.6151
R1404 B.n526 B.n525 10.6151
R1405 B.n527 B.n526 10.6151
R1406 B.n527 B.n264 10.6151
R1407 B.n537 B.n264 10.6151
R1408 B.n538 B.n537 10.6151
R1409 B.n539 B.n538 10.6151
R1410 B.n539 B.n256 10.6151
R1411 B.n549 B.n256 10.6151
R1412 B.n550 B.n549 10.6151
R1413 B.n551 B.n550 10.6151
R1414 B.n551 B.n248 10.6151
R1415 B.n561 B.n248 10.6151
R1416 B.n562 B.n561 10.6151
R1417 B.n563 B.n562 10.6151
R1418 B.n563 B.n240 10.6151
R1419 B.n573 B.n240 10.6151
R1420 B.n574 B.n573 10.6151
R1421 B.n575 B.n574 10.6151
R1422 B.n575 B.n232 10.6151
R1423 B.n586 B.n232 10.6151
R1424 B.n587 B.n586 10.6151
R1425 B.n588 B.n587 10.6151
R1426 B.n588 B.n0 10.6151
R1427 B.n346 B.n311 10.6151
R1428 B.n346 B.n345 10.6151
R1429 B.n352 B.n345 10.6151
R1430 B.n353 B.n352 10.6151
R1431 B.n354 B.n353 10.6151
R1432 B.n354 B.n343 10.6151
R1433 B.n360 B.n343 10.6151
R1434 B.n361 B.n360 10.6151
R1435 B.n362 B.n361 10.6151
R1436 B.n362 B.n341 10.6151
R1437 B.n368 B.n341 10.6151
R1438 B.n369 B.n368 10.6151
R1439 B.n370 B.n369 10.6151
R1440 B.n370 B.n339 10.6151
R1441 B.n376 B.n339 10.6151
R1442 B.n377 B.n376 10.6151
R1443 B.n378 B.n377 10.6151
R1444 B.n378 B.n337 10.6151
R1445 B.n384 B.n337 10.6151
R1446 B.n385 B.n384 10.6151
R1447 B.n386 B.n385 10.6151
R1448 B.n386 B.n335 10.6151
R1449 B.n392 B.n335 10.6151
R1450 B.n395 B.n394 10.6151
R1451 B.n395 B.n331 10.6151
R1452 B.n401 B.n331 10.6151
R1453 B.n402 B.n401 10.6151
R1454 B.n403 B.n402 10.6151
R1455 B.n403 B.n329 10.6151
R1456 B.n409 B.n329 10.6151
R1457 B.n410 B.n409 10.6151
R1458 B.n412 B.n325 10.6151
R1459 B.n418 B.n325 10.6151
R1460 B.n419 B.n418 10.6151
R1461 B.n420 B.n419 10.6151
R1462 B.n420 B.n323 10.6151
R1463 B.n426 B.n323 10.6151
R1464 B.n427 B.n426 10.6151
R1465 B.n428 B.n427 10.6151
R1466 B.n428 B.n321 10.6151
R1467 B.n434 B.n321 10.6151
R1468 B.n435 B.n434 10.6151
R1469 B.n436 B.n435 10.6151
R1470 B.n436 B.n319 10.6151
R1471 B.n442 B.n319 10.6151
R1472 B.n443 B.n442 10.6151
R1473 B.n444 B.n443 10.6151
R1474 B.n444 B.n317 10.6151
R1475 B.n450 B.n317 10.6151
R1476 B.n451 B.n450 10.6151
R1477 B.n452 B.n451 10.6151
R1478 B.n452 B.n315 10.6151
R1479 B.n458 B.n315 10.6151
R1480 B.n459 B.n458 10.6151
R1481 B.n460 B.n307 10.6151
R1482 B.n470 B.n307 10.6151
R1483 B.n471 B.n470 10.6151
R1484 B.n472 B.n471 10.6151
R1485 B.n472 B.n299 10.6151
R1486 B.n482 B.n299 10.6151
R1487 B.n483 B.n482 10.6151
R1488 B.n484 B.n483 10.6151
R1489 B.n484 B.n292 10.6151
R1490 B.n495 B.n292 10.6151
R1491 B.n496 B.n495 10.6151
R1492 B.n497 B.n496 10.6151
R1493 B.n497 B.n284 10.6151
R1494 B.n507 B.n284 10.6151
R1495 B.n508 B.n507 10.6151
R1496 B.n509 B.n508 10.6151
R1497 B.n509 B.n276 10.6151
R1498 B.n519 B.n276 10.6151
R1499 B.n520 B.n519 10.6151
R1500 B.n521 B.n520 10.6151
R1501 B.n521 B.n268 10.6151
R1502 B.n531 B.n268 10.6151
R1503 B.n532 B.n531 10.6151
R1504 B.n533 B.n532 10.6151
R1505 B.n533 B.n260 10.6151
R1506 B.n543 B.n260 10.6151
R1507 B.n544 B.n543 10.6151
R1508 B.n545 B.n544 10.6151
R1509 B.n545 B.n252 10.6151
R1510 B.n555 B.n252 10.6151
R1511 B.n556 B.n555 10.6151
R1512 B.n557 B.n556 10.6151
R1513 B.n557 B.n244 10.6151
R1514 B.n567 B.n244 10.6151
R1515 B.n568 B.n567 10.6151
R1516 B.n569 B.n568 10.6151
R1517 B.n569 B.n236 10.6151
R1518 B.n579 B.n236 10.6151
R1519 B.n580 B.n579 10.6151
R1520 B.n582 B.n580 10.6151
R1521 B.n582 B.n581 10.6151
R1522 B.n581 B.n228 10.6151
R1523 B.n593 B.n228 10.6151
R1524 B.n594 B.n593 10.6151
R1525 B.n595 B.n594 10.6151
R1526 B.n596 B.n595 10.6151
R1527 B.n597 B.n596 10.6151
R1528 B.n600 B.n597 10.6151
R1529 B.n601 B.n600 10.6151
R1530 B.n602 B.n601 10.6151
R1531 B.n603 B.n602 10.6151
R1532 B.n605 B.n603 10.6151
R1533 B.n606 B.n605 10.6151
R1534 B.n607 B.n606 10.6151
R1535 B.n608 B.n607 10.6151
R1536 B.n610 B.n608 10.6151
R1537 B.n611 B.n610 10.6151
R1538 B.n612 B.n611 10.6151
R1539 B.n613 B.n612 10.6151
R1540 B.n615 B.n613 10.6151
R1541 B.n616 B.n615 10.6151
R1542 B.n617 B.n616 10.6151
R1543 B.n618 B.n617 10.6151
R1544 B.n620 B.n618 10.6151
R1545 B.n621 B.n620 10.6151
R1546 B.n622 B.n621 10.6151
R1547 B.n623 B.n622 10.6151
R1548 B.n625 B.n623 10.6151
R1549 B.n626 B.n625 10.6151
R1550 B.n627 B.n626 10.6151
R1551 B.n628 B.n627 10.6151
R1552 B.n630 B.n628 10.6151
R1553 B.n631 B.n630 10.6151
R1554 B.n632 B.n631 10.6151
R1555 B.n633 B.n632 10.6151
R1556 B.n635 B.n633 10.6151
R1557 B.n636 B.n635 10.6151
R1558 B.n637 B.n636 10.6151
R1559 B.n638 B.n637 10.6151
R1560 B.n640 B.n638 10.6151
R1561 B.n641 B.n640 10.6151
R1562 B.n642 B.n641 10.6151
R1563 B.n643 B.n642 10.6151
R1564 B.n645 B.n643 10.6151
R1565 B.n646 B.n645 10.6151
R1566 B.n647 B.n646 10.6151
R1567 B.n648 B.n647 10.6151
R1568 B.n650 B.n648 10.6151
R1569 B.n651 B.n650 10.6151
R1570 B.n739 B.n1 10.6151
R1571 B.n739 B.n738 10.6151
R1572 B.n738 B.n737 10.6151
R1573 B.n737 B.n10 10.6151
R1574 B.n731 B.n10 10.6151
R1575 B.n731 B.n730 10.6151
R1576 B.n730 B.n729 10.6151
R1577 B.n729 B.n18 10.6151
R1578 B.n723 B.n18 10.6151
R1579 B.n723 B.n722 10.6151
R1580 B.n722 B.n721 10.6151
R1581 B.n721 B.n25 10.6151
R1582 B.n715 B.n25 10.6151
R1583 B.n715 B.n714 10.6151
R1584 B.n714 B.n713 10.6151
R1585 B.n713 B.n32 10.6151
R1586 B.n707 B.n32 10.6151
R1587 B.n707 B.n706 10.6151
R1588 B.n706 B.n705 10.6151
R1589 B.n705 B.n39 10.6151
R1590 B.n699 B.n39 10.6151
R1591 B.n699 B.n698 10.6151
R1592 B.n698 B.n697 10.6151
R1593 B.n697 B.n46 10.6151
R1594 B.n691 B.n46 10.6151
R1595 B.n691 B.n690 10.6151
R1596 B.n690 B.n689 10.6151
R1597 B.n689 B.n53 10.6151
R1598 B.n683 B.n53 10.6151
R1599 B.n683 B.n682 10.6151
R1600 B.n682 B.n681 10.6151
R1601 B.n681 B.n60 10.6151
R1602 B.n675 B.n60 10.6151
R1603 B.n675 B.n674 10.6151
R1604 B.n674 B.n673 10.6151
R1605 B.n673 B.n66 10.6151
R1606 B.n667 B.n66 10.6151
R1607 B.n667 B.n666 10.6151
R1608 B.n666 B.n665 10.6151
R1609 B.n665 B.n74 10.6151
R1610 B.n659 B.n74 10.6151
R1611 B.n659 B.n658 10.6151
R1612 B.n658 B.n657 10.6151
R1613 B.n118 B.n81 10.6151
R1614 B.n121 B.n118 10.6151
R1615 B.n122 B.n121 10.6151
R1616 B.n125 B.n122 10.6151
R1617 B.n126 B.n125 10.6151
R1618 B.n129 B.n126 10.6151
R1619 B.n130 B.n129 10.6151
R1620 B.n133 B.n130 10.6151
R1621 B.n134 B.n133 10.6151
R1622 B.n137 B.n134 10.6151
R1623 B.n138 B.n137 10.6151
R1624 B.n141 B.n138 10.6151
R1625 B.n142 B.n141 10.6151
R1626 B.n145 B.n142 10.6151
R1627 B.n146 B.n145 10.6151
R1628 B.n149 B.n146 10.6151
R1629 B.n150 B.n149 10.6151
R1630 B.n153 B.n150 10.6151
R1631 B.n154 B.n153 10.6151
R1632 B.n157 B.n154 10.6151
R1633 B.n158 B.n157 10.6151
R1634 B.n161 B.n158 10.6151
R1635 B.n162 B.n161 10.6151
R1636 B.n166 B.n165 10.6151
R1637 B.n169 B.n166 10.6151
R1638 B.n170 B.n169 10.6151
R1639 B.n173 B.n170 10.6151
R1640 B.n174 B.n173 10.6151
R1641 B.n177 B.n174 10.6151
R1642 B.n178 B.n177 10.6151
R1643 B.n181 B.n178 10.6151
R1644 B.n186 B.n183 10.6151
R1645 B.n187 B.n186 10.6151
R1646 B.n190 B.n187 10.6151
R1647 B.n191 B.n190 10.6151
R1648 B.n194 B.n191 10.6151
R1649 B.n195 B.n194 10.6151
R1650 B.n198 B.n195 10.6151
R1651 B.n199 B.n198 10.6151
R1652 B.n202 B.n199 10.6151
R1653 B.n203 B.n202 10.6151
R1654 B.n206 B.n203 10.6151
R1655 B.n207 B.n206 10.6151
R1656 B.n210 B.n207 10.6151
R1657 B.n211 B.n210 10.6151
R1658 B.n214 B.n211 10.6151
R1659 B.n215 B.n214 10.6151
R1660 B.n218 B.n215 10.6151
R1661 B.n219 B.n218 10.6151
R1662 B.n222 B.n219 10.6151
R1663 B.n223 B.n222 10.6151
R1664 B.n226 B.n223 10.6151
R1665 B.n227 B.n226 10.6151
R1666 B.n652 B.n227 10.6151
R1667 B.t0 B.n238 9.8704
R1668 B.t1 B.n16 9.8704
R1669 B.n747 B.n0 8.11757
R1670 B.n747 B.n1 8.11757
R1671 B.n394 B.n393 6.5566
R1672 B.n411 B.n410 6.5566
R1673 B.n165 B.n117 6.5566
R1674 B.n182 B.n181 6.5566
R1675 B.n393 B.n392 4.05904
R1676 B.n412 B.n411 4.05904
R1677 B.n162 B.n117 4.05904
R1678 B.n183 B.n182 4.05904
R1679 VP.n21 VP.n20 161.3
R1680 VP.n19 VP.n1 161.3
R1681 VP.n18 VP.n17 161.3
R1682 VP.n16 VP.n2 161.3
R1683 VP.n15 VP.n14 161.3
R1684 VP.n13 VP.n3 161.3
R1685 VP.n12 VP.n11 161.3
R1686 VP.n10 VP.n4 161.3
R1687 VP.n9 VP.n8 161.3
R1688 VP.n7 VP.n6 87.376
R1689 VP.n22 VP.n0 87.376
R1690 VP.n5 VP.t1 71.2408
R1691 VP.n5 VP.t3 69.8958
R1692 VP.n6 VP.n5 47.1964
R1693 VP.n14 VP.n13 40.4934
R1694 VP.n14 VP.n2 40.4934
R1695 VP.n7 VP.t2 37.4256
R1696 VP.n0 VP.t0 37.4256
R1697 VP.n8 VP.n4 24.4675
R1698 VP.n12 VP.n4 24.4675
R1699 VP.n13 VP.n12 24.4675
R1700 VP.n18 VP.n2 24.4675
R1701 VP.n19 VP.n18 24.4675
R1702 VP.n20 VP.n19 24.4675
R1703 VP.n8 VP.n7 2.69187
R1704 VP.n20 VP.n0 2.69187
R1705 VP.n9 VP.n6 0.354971
R1706 VP.n22 VP.n21 0.354971
R1707 VP VP.n22 0.26696
R1708 VP.n10 VP.n9 0.189894
R1709 VP.n11 VP.n10 0.189894
R1710 VP.n11 VP.n3 0.189894
R1711 VP.n15 VP.n3 0.189894
R1712 VP.n16 VP.n15 0.189894
R1713 VP.n17 VP.n16 0.189894
R1714 VP.n17 VP.n1 0.189894
R1715 VP.n21 VP.n1 0.189894
R1716 VDD1 VDD1.n1 110.764
R1717 VDD1 VDD1.n0 70.8928
R1718 VDD1.n0 VDD1.t2 3.37358
R1719 VDD1.n0 VDD1.t0 3.37358
R1720 VDD1.n1 VDD1.t1 3.37358
R1721 VDD1.n1 VDD1.t3 3.37358
C0 VDD1 VDD2 1.31245f
C1 VP VN 5.90735f
C2 VN VTAIL 3.16725f
C3 VP VTAIL 3.18135f
C4 VDD1 VN 0.149921f
C5 VN VDD2 2.63613f
C6 VDD1 VTAIL 4.46265f
C7 VP VDD1 2.95442f
C8 VP VDD2 0.469245f
C9 VTAIL VDD2 4.52477f
C10 VDD2 B 3.961437f
C11 VDD1 B 8.08287f
C12 VTAIL B 6.660898f
C13 VN B 12.47305f
C14 VP B 10.864256f
C15 VDD1.t2 B 0.13645f
C16 VDD1.t0 B 0.13645f
C17 VDD1.n0 B 1.14815f
C18 VDD1.t1 B 0.13645f
C19 VDD1.t3 B 0.13645f
C20 VDD1.n1 B 1.6934f
C21 VP.t0 B 1.42834f
C22 VP.n0 B 0.617886f
C23 VP.n1 B 0.024353f
C24 VP.n2 B 0.048401f
C25 VP.n3 B 0.024353f
C26 VP.n4 B 0.045388f
C27 VP.t1 B 1.7738f
C28 VP.t3 B 1.76044f
C29 VP.n5 B 2.45482f
C30 VP.n6 B 1.29604f
C31 VP.t2 B 1.42834f
C32 VP.n7 B 0.617886f
C33 VP.n8 B 0.025443f
C34 VP.n9 B 0.039305f
C35 VP.n10 B 0.024353f
C36 VP.n11 B 0.024353f
C37 VP.n12 B 0.045388f
C38 VP.n13 B 0.048401f
C39 VP.n14 B 0.019687f
C40 VP.n15 B 0.024353f
C41 VP.n16 B 0.024353f
C42 VP.n17 B 0.024353f
C43 VP.n18 B 0.045388f
C44 VP.n19 B 0.045388f
C45 VP.n20 B 0.025443f
C46 VP.n21 B 0.039305f
C47 VP.n22 B 0.074679f
C48 VTAIL.n0 B 0.011967f
C49 VTAIL.n1 B 0.026927f
C50 VTAIL.n2 B 0.012062f
C51 VTAIL.n3 B 0.0212f
C52 VTAIL.n4 B 0.011392f
C53 VTAIL.n5 B 0.026927f
C54 VTAIL.n6 B 0.012062f
C55 VTAIL.n7 B 0.491138f
C56 VTAIL.n8 B 0.011392f
C57 VTAIL.t4 B 0.044903f
C58 VTAIL.n9 B 0.103182f
C59 VTAIL.n10 B 0.019034f
C60 VTAIL.n11 B 0.020195f
C61 VTAIL.n12 B 0.026927f
C62 VTAIL.n13 B 0.012062f
C63 VTAIL.n14 B 0.011392f
C64 VTAIL.n15 B 0.0212f
C65 VTAIL.n16 B 0.0212f
C66 VTAIL.n17 B 0.011392f
C67 VTAIL.n18 B 0.012062f
C68 VTAIL.n19 B 0.026927f
C69 VTAIL.n20 B 0.026927f
C70 VTAIL.n21 B 0.012062f
C71 VTAIL.n22 B 0.011392f
C72 VTAIL.n23 B 0.0212f
C73 VTAIL.n24 B 0.055665f
C74 VTAIL.n25 B 0.011392f
C75 VTAIL.n26 B 0.012062f
C76 VTAIL.n27 B 0.055004f
C77 VTAIL.n28 B 0.04692f
C78 VTAIL.n29 B 0.177981f
C79 VTAIL.n30 B 0.011967f
C80 VTAIL.n31 B 0.026927f
C81 VTAIL.n32 B 0.012062f
C82 VTAIL.n33 B 0.0212f
C83 VTAIL.n34 B 0.011392f
C84 VTAIL.n35 B 0.026927f
C85 VTAIL.n36 B 0.012062f
C86 VTAIL.n37 B 0.491138f
C87 VTAIL.n38 B 0.011392f
C88 VTAIL.t0 B 0.044903f
C89 VTAIL.n39 B 0.103182f
C90 VTAIL.n40 B 0.019034f
C91 VTAIL.n41 B 0.020195f
C92 VTAIL.n42 B 0.026927f
C93 VTAIL.n43 B 0.012062f
C94 VTAIL.n44 B 0.011392f
C95 VTAIL.n45 B 0.0212f
C96 VTAIL.n46 B 0.0212f
C97 VTAIL.n47 B 0.011392f
C98 VTAIL.n48 B 0.012062f
C99 VTAIL.n49 B 0.026927f
C100 VTAIL.n50 B 0.026927f
C101 VTAIL.n51 B 0.012062f
C102 VTAIL.n52 B 0.011392f
C103 VTAIL.n53 B 0.0212f
C104 VTAIL.n54 B 0.055665f
C105 VTAIL.n55 B 0.011392f
C106 VTAIL.n56 B 0.012062f
C107 VTAIL.n57 B 0.055004f
C108 VTAIL.n58 B 0.04692f
C109 VTAIL.n59 B 0.295024f
C110 VTAIL.n60 B 0.011967f
C111 VTAIL.n61 B 0.026927f
C112 VTAIL.n62 B 0.012062f
C113 VTAIL.n63 B 0.0212f
C114 VTAIL.n64 B 0.011392f
C115 VTAIL.n65 B 0.026927f
C116 VTAIL.n66 B 0.012062f
C117 VTAIL.n67 B 0.491138f
C118 VTAIL.n68 B 0.011392f
C119 VTAIL.t2 B 0.044903f
C120 VTAIL.n69 B 0.103182f
C121 VTAIL.n70 B 0.019034f
C122 VTAIL.n71 B 0.020195f
C123 VTAIL.n72 B 0.026927f
C124 VTAIL.n73 B 0.012062f
C125 VTAIL.n74 B 0.011392f
C126 VTAIL.n75 B 0.0212f
C127 VTAIL.n76 B 0.0212f
C128 VTAIL.n77 B 0.011392f
C129 VTAIL.n78 B 0.012062f
C130 VTAIL.n79 B 0.026927f
C131 VTAIL.n80 B 0.026927f
C132 VTAIL.n81 B 0.012062f
C133 VTAIL.n82 B 0.011392f
C134 VTAIL.n83 B 0.0212f
C135 VTAIL.n84 B 0.055665f
C136 VTAIL.n85 B 0.011392f
C137 VTAIL.n86 B 0.012062f
C138 VTAIL.n87 B 0.055004f
C139 VTAIL.n88 B 0.04692f
C140 VTAIL.n89 B 1.13863f
C141 VTAIL.n90 B 0.011967f
C142 VTAIL.n91 B 0.026927f
C143 VTAIL.n92 B 0.012062f
C144 VTAIL.n93 B 0.0212f
C145 VTAIL.n94 B 0.011392f
C146 VTAIL.n95 B 0.026927f
C147 VTAIL.n96 B 0.012062f
C148 VTAIL.n97 B 0.491138f
C149 VTAIL.n98 B 0.011392f
C150 VTAIL.t7 B 0.044903f
C151 VTAIL.n99 B 0.103182f
C152 VTAIL.n100 B 0.019034f
C153 VTAIL.n101 B 0.020195f
C154 VTAIL.n102 B 0.026927f
C155 VTAIL.n103 B 0.012062f
C156 VTAIL.n104 B 0.011392f
C157 VTAIL.n105 B 0.0212f
C158 VTAIL.n106 B 0.0212f
C159 VTAIL.n107 B 0.011392f
C160 VTAIL.n108 B 0.012062f
C161 VTAIL.n109 B 0.026927f
C162 VTAIL.n110 B 0.026927f
C163 VTAIL.n111 B 0.012062f
C164 VTAIL.n112 B 0.011392f
C165 VTAIL.n113 B 0.0212f
C166 VTAIL.n114 B 0.055665f
C167 VTAIL.n115 B 0.011392f
C168 VTAIL.n116 B 0.012062f
C169 VTAIL.n117 B 0.055004f
C170 VTAIL.n118 B 0.04692f
C171 VTAIL.n119 B 1.13863f
C172 VTAIL.n120 B 0.011967f
C173 VTAIL.n121 B 0.026927f
C174 VTAIL.n122 B 0.012062f
C175 VTAIL.n123 B 0.0212f
C176 VTAIL.n124 B 0.011392f
C177 VTAIL.n125 B 0.026927f
C178 VTAIL.n126 B 0.012062f
C179 VTAIL.n127 B 0.491138f
C180 VTAIL.n128 B 0.011392f
C181 VTAIL.t5 B 0.044903f
C182 VTAIL.n129 B 0.103182f
C183 VTAIL.n130 B 0.019034f
C184 VTAIL.n131 B 0.020195f
C185 VTAIL.n132 B 0.026927f
C186 VTAIL.n133 B 0.012062f
C187 VTAIL.n134 B 0.011392f
C188 VTAIL.n135 B 0.0212f
C189 VTAIL.n136 B 0.0212f
C190 VTAIL.n137 B 0.011392f
C191 VTAIL.n138 B 0.012062f
C192 VTAIL.n139 B 0.026927f
C193 VTAIL.n140 B 0.026927f
C194 VTAIL.n141 B 0.012062f
C195 VTAIL.n142 B 0.011392f
C196 VTAIL.n143 B 0.0212f
C197 VTAIL.n144 B 0.055665f
C198 VTAIL.n145 B 0.011392f
C199 VTAIL.n146 B 0.012062f
C200 VTAIL.n147 B 0.055004f
C201 VTAIL.n148 B 0.04692f
C202 VTAIL.n149 B 0.295024f
C203 VTAIL.n150 B 0.011967f
C204 VTAIL.n151 B 0.026927f
C205 VTAIL.n152 B 0.012062f
C206 VTAIL.n153 B 0.0212f
C207 VTAIL.n154 B 0.011392f
C208 VTAIL.n155 B 0.026927f
C209 VTAIL.n156 B 0.012062f
C210 VTAIL.n157 B 0.491138f
C211 VTAIL.n158 B 0.011392f
C212 VTAIL.t1 B 0.044903f
C213 VTAIL.n159 B 0.103182f
C214 VTAIL.n160 B 0.019034f
C215 VTAIL.n161 B 0.020195f
C216 VTAIL.n162 B 0.026927f
C217 VTAIL.n163 B 0.012062f
C218 VTAIL.n164 B 0.011392f
C219 VTAIL.n165 B 0.0212f
C220 VTAIL.n166 B 0.0212f
C221 VTAIL.n167 B 0.011392f
C222 VTAIL.n168 B 0.012062f
C223 VTAIL.n169 B 0.026927f
C224 VTAIL.n170 B 0.026927f
C225 VTAIL.n171 B 0.012062f
C226 VTAIL.n172 B 0.011392f
C227 VTAIL.n173 B 0.0212f
C228 VTAIL.n174 B 0.055665f
C229 VTAIL.n175 B 0.011392f
C230 VTAIL.n176 B 0.012062f
C231 VTAIL.n177 B 0.055004f
C232 VTAIL.n178 B 0.04692f
C233 VTAIL.n179 B 0.295024f
C234 VTAIL.n180 B 0.011967f
C235 VTAIL.n181 B 0.026927f
C236 VTAIL.n182 B 0.012062f
C237 VTAIL.n183 B 0.0212f
C238 VTAIL.n184 B 0.011392f
C239 VTAIL.n185 B 0.026927f
C240 VTAIL.n186 B 0.012062f
C241 VTAIL.n187 B 0.491138f
C242 VTAIL.n188 B 0.011392f
C243 VTAIL.t3 B 0.044903f
C244 VTAIL.n189 B 0.103182f
C245 VTAIL.n190 B 0.019034f
C246 VTAIL.n191 B 0.020195f
C247 VTAIL.n192 B 0.026927f
C248 VTAIL.n193 B 0.012062f
C249 VTAIL.n194 B 0.011392f
C250 VTAIL.n195 B 0.0212f
C251 VTAIL.n196 B 0.0212f
C252 VTAIL.n197 B 0.011392f
C253 VTAIL.n198 B 0.012062f
C254 VTAIL.n199 B 0.026927f
C255 VTAIL.n200 B 0.026927f
C256 VTAIL.n201 B 0.012062f
C257 VTAIL.n202 B 0.011392f
C258 VTAIL.n203 B 0.0212f
C259 VTAIL.n204 B 0.055665f
C260 VTAIL.n205 B 0.011392f
C261 VTAIL.n206 B 0.012062f
C262 VTAIL.n207 B 0.055004f
C263 VTAIL.n208 B 0.04692f
C264 VTAIL.n209 B 1.13863f
C265 VTAIL.n210 B 0.011967f
C266 VTAIL.n211 B 0.026927f
C267 VTAIL.n212 B 0.012062f
C268 VTAIL.n213 B 0.0212f
C269 VTAIL.n214 B 0.011392f
C270 VTAIL.n215 B 0.026927f
C271 VTAIL.n216 B 0.012062f
C272 VTAIL.n217 B 0.491138f
C273 VTAIL.n218 B 0.011392f
C274 VTAIL.t6 B 0.044903f
C275 VTAIL.n219 B 0.103182f
C276 VTAIL.n220 B 0.019034f
C277 VTAIL.n221 B 0.020195f
C278 VTAIL.n222 B 0.026927f
C279 VTAIL.n223 B 0.012062f
C280 VTAIL.n224 B 0.011392f
C281 VTAIL.n225 B 0.0212f
C282 VTAIL.n226 B 0.0212f
C283 VTAIL.n227 B 0.011392f
C284 VTAIL.n228 B 0.012062f
C285 VTAIL.n229 B 0.026927f
C286 VTAIL.n230 B 0.026927f
C287 VTAIL.n231 B 0.012062f
C288 VTAIL.n232 B 0.011392f
C289 VTAIL.n233 B 0.0212f
C290 VTAIL.n234 B 0.055665f
C291 VTAIL.n235 B 0.011392f
C292 VTAIL.n236 B 0.012062f
C293 VTAIL.n237 B 0.055004f
C294 VTAIL.n238 B 0.04692f
C295 VTAIL.n239 B 1.01364f
C296 VDD2.t1 B 0.131072f
C297 VDD2.t3 B 0.131072f
C298 VDD2.n0 B 1.60211f
C299 VDD2.t0 B 0.131072f
C300 VDD2.t2 B 0.131072f
C301 VDD2.n1 B 1.10244f
C302 VDD2.n2 B 3.54248f
C303 VN.t1 B 1.69744f
C304 VN.t3 B 1.71032f
C305 VN.n0 B 1.01098f
C306 VN.t0 B 1.69744f
C307 VN.t2 B 1.71032f
C308 VN.n1 B 2.37674f
.ends

