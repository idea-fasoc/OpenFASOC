* NGSPICE file created from diff_pair_sample_0914.ext - technology: sky130A

.subckt diff_pair_sample_0914 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=3.07395 pd=18.96 as=7.2657 ps=38.04 w=18.63 l=3.51
X1 VTAIL.t10 VP.t1 VDD1.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=3.07395 pd=18.96 as=3.07395 ps=18.96 w=18.63 l=3.51
X2 VTAIL.t15 VP.t2 VDD1.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=3.07395 pd=18.96 as=3.07395 ps=18.96 w=18.63 l=3.51
X3 VDD2.t9 VN.t0 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=7.2657 pd=38.04 as=3.07395 ps=18.96 w=18.63 l=3.51
X4 VTAIL.t8 VN.t1 VDD2.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=3.07395 pd=18.96 as=3.07395 ps=18.96 w=18.63 l=3.51
X5 VDD1.t6 VP.t3 VTAIL.t16 B.t6 sky130_fd_pr__nfet_01v8 ad=3.07395 pd=18.96 as=3.07395 ps=18.96 w=18.63 l=3.51
X6 VTAIL.t7 VN.t2 VDD2.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=3.07395 pd=18.96 as=3.07395 ps=18.96 w=18.63 l=3.51
X7 VDD1.t5 VP.t4 VTAIL.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=7.2657 pd=38.04 as=3.07395 ps=18.96 w=18.63 l=3.51
X8 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=7.2657 pd=38.04 as=0 ps=0 w=18.63 l=3.51
X9 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=7.2657 pd=38.04 as=0 ps=0 w=18.63 l=3.51
X10 VDD1.t4 VP.t5 VTAIL.t17 B.t4 sky130_fd_pr__nfet_01v8 ad=3.07395 pd=18.96 as=3.07395 ps=18.96 w=18.63 l=3.51
X11 VDD1.t3 VP.t6 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=3.07395 pd=18.96 as=7.2657 ps=38.04 w=18.63 l=3.51
X12 VDD2.t6 VN.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=3.07395 pd=18.96 as=3.07395 ps=18.96 w=18.63 l=3.51
X13 VDD2.t5 VN.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=7.2657 pd=38.04 as=3.07395 ps=18.96 w=18.63 l=3.51
X14 VDD2.t4 VN.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.07395 pd=18.96 as=3.07395 ps=18.96 w=18.63 l=3.51
X15 VDD2.t3 VN.t6 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.07395 pd=18.96 as=7.2657 ps=38.04 w=18.63 l=3.51
X16 VDD2.t2 VN.t7 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.07395 pd=18.96 as=7.2657 ps=38.04 w=18.63 l=3.51
X17 VTAIL.t1 VN.t8 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.07395 pd=18.96 as=3.07395 ps=18.96 w=18.63 l=3.51
X18 VTAIL.t19 VP.t7 VDD1.t2 B.t8 sky130_fd_pr__nfet_01v8 ad=3.07395 pd=18.96 as=3.07395 ps=18.96 w=18.63 l=3.51
X19 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=7.2657 pd=38.04 as=0 ps=0 w=18.63 l=3.51
X20 VDD1.t1 VP.t8 VTAIL.t18 B.t5 sky130_fd_pr__nfet_01v8 ad=7.2657 pd=38.04 as=3.07395 ps=18.96 w=18.63 l=3.51
X21 VTAIL.t12 VP.t9 VDD1.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=3.07395 pd=18.96 as=3.07395 ps=18.96 w=18.63 l=3.51
X22 VTAIL.t0 VN.t9 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.07395 pd=18.96 as=3.07395 ps=18.96 w=18.63 l=3.51
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.2657 pd=38.04 as=0 ps=0 w=18.63 l=3.51
R0 VP.n32 VP.n31 161.3
R1 VP.n33 VP.n28 161.3
R2 VP.n35 VP.n34 161.3
R3 VP.n36 VP.n27 161.3
R4 VP.n38 VP.n37 161.3
R5 VP.n39 VP.n26 161.3
R6 VP.n41 VP.n40 161.3
R7 VP.n42 VP.n25 161.3
R8 VP.n44 VP.n43 161.3
R9 VP.n45 VP.n24 161.3
R10 VP.n47 VP.n46 161.3
R11 VP.n48 VP.n23 161.3
R12 VP.n50 VP.n49 161.3
R13 VP.n51 VP.n22 161.3
R14 VP.n54 VP.n53 161.3
R15 VP.n55 VP.n21 161.3
R16 VP.n57 VP.n56 161.3
R17 VP.n58 VP.n20 161.3
R18 VP.n60 VP.n59 161.3
R19 VP.n61 VP.n19 161.3
R20 VP.n63 VP.n62 161.3
R21 VP.n64 VP.n18 161.3
R22 VP.n66 VP.n65 161.3
R23 VP.n117 VP.n116 161.3
R24 VP.n115 VP.n1 161.3
R25 VP.n114 VP.n113 161.3
R26 VP.n112 VP.n2 161.3
R27 VP.n111 VP.n110 161.3
R28 VP.n109 VP.n3 161.3
R29 VP.n108 VP.n107 161.3
R30 VP.n106 VP.n4 161.3
R31 VP.n105 VP.n104 161.3
R32 VP.n102 VP.n5 161.3
R33 VP.n101 VP.n100 161.3
R34 VP.n99 VP.n6 161.3
R35 VP.n98 VP.n97 161.3
R36 VP.n96 VP.n7 161.3
R37 VP.n95 VP.n94 161.3
R38 VP.n93 VP.n8 161.3
R39 VP.n92 VP.n91 161.3
R40 VP.n90 VP.n9 161.3
R41 VP.n89 VP.n88 161.3
R42 VP.n87 VP.n10 161.3
R43 VP.n86 VP.n85 161.3
R44 VP.n84 VP.n11 161.3
R45 VP.n83 VP.n82 161.3
R46 VP.n81 VP.n80 161.3
R47 VP.n79 VP.n13 161.3
R48 VP.n78 VP.n77 161.3
R49 VP.n76 VP.n14 161.3
R50 VP.n75 VP.n74 161.3
R51 VP.n73 VP.n15 161.3
R52 VP.n72 VP.n71 161.3
R53 VP.n70 VP.n16 161.3
R54 VP.n30 VP.t8 161.114
R55 VP.n8 VP.t5 127.915
R56 VP.n68 VP.t4 127.915
R57 VP.n12 VP.t9 127.915
R58 VP.n103 VP.t2 127.915
R59 VP.n0 VP.t6 127.915
R60 VP.n25 VP.t3 127.915
R61 VP.n17 VP.t0 127.915
R62 VP.n52 VP.t1 127.915
R63 VP.n29 VP.t7 127.915
R64 VP.n69 VP.n68 81.2593
R65 VP.n118 VP.n0 81.2593
R66 VP.n67 VP.n17 81.2593
R67 VP.n69 VP.n67 63.1584
R68 VP.n30 VP.n29 57.9282
R69 VP.n74 VP.n14 56.5193
R70 VP.n110 VP.n2 56.5193
R71 VP.n59 VP.n19 56.5193
R72 VP.n89 VP.n10 48.2635
R73 VP.n97 VP.n6 48.2635
R74 VP.n46 VP.n23 48.2635
R75 VP.n38 VP.n27 48.2635
R76 VP.n85 VP.n10 32.7233
R77 VP.n101 VP.n6 32.7233
R78 VP.n50 VP.n23 32.7233
R79 VP.n34 VP.n27 32.7233
R80 VP.n72 VP.n16 24.4675
R81 VP.n73 VP.n72 24.4675
R82 VP.n74 VP.n73 24.4675
R83 VP.n78 VP.n14 24.4675
R84 VP.n79 VP.n78 24.4675
R85 VP.n80 VP.n79 24.4675
R86 VP.n84 VP.n83 24.4675
R87 VP.n85 VP.n84 24.4675
R88 VP.n90 VP.n89 24.4675
R89 VP.n91 VP.n90 24.4675
R90 VP.n91 VP.n8 24.4675
R91 VP.n95 VP.n8 24.4675
R92 VP.n96 VP.n95 24.4675
R93 VP.n97 VP.n96 24.4675
R94 VP.n102 VP.n101 24.4675
R95 VP.n104 VP.n102 24.4675
R96 VP.n108 VP.n4 24.4675
R97 VP.n109 VP.n108 24.4675
R98 VP.n110 VP.n109 24.4675
R99 VP.n114 VP.n2 24.4675
R100 VP.n115 VP.n114 24.4675
R101 VP.n116 VP.n115 24.4675
R102 VP.n63 VP.n19 24.4675
R103 VP.n64 VP.n63 24.4675
R104 VP.n65 VP.n64 24.4675
R105 VP.n51 VP.n50 24.4675
R106 VP.n53 VP.n51 24.4675
R107 VP.n57 VP.n21 24.4675
R108 VP.n58 VP.n57 24.4675
R109 VP.n59 VP.n58 24.4675
R110 VP.n39 VP.n38 24.4675
R111 VP.n40 VP.n39 24.4675
R112 VP.n40 VP.n25 24.4675
R113 VP.n44 VP.n25 24.4675
R114 VP.n45 VP.n44 24.4675
R115 VP.n46 VP.n45 24.4675
R116 VP.n33 VP.n32 24.4675
R117 VP.n34 VP.n33 24.4675
R118 VP.n83 VP.n12 16.6381
R119 VP.n104 VP.n103 16.6381
R120 VP.n53 VP.n52 16.6381
R121 VP.n32 VP.n29 16.6381
R122 VP.n68 VP.n16 8.80862
R123 VP.n116 VP.n0 8.80862
R124 VP.n65 VP.n17 8.80862
R125 VP.n80 VP.n12 7.82994
R126 VP.n103 VP.n4 7.82994
R127 VP.n52 VP.n21 7.82994
R128 VP.n31 VP.n30 3.19587
R129 VP.n67 VP.n66 0.354971
R130 VP.n70 VP.n69 0.354971
R131 VP.n118 VP.n117 0.354971
R132 VP VP.n118 0.26696
R133 VP.n31 VP.n28 0.189894
R134 VP.n35 VP.n28 0.189894
R135 VP.n36 VP.n35 0.189894
R136 VP.n37 VP.n36 0.189894
R137 VP.n37 VP.n26 0.189894
R138 VP.n41 VP.n26 0.189894
R139 VP.n42 VP.n41 0.189894
R140 VP.n43 VP.n42 0.189894
R141 VP.n43 VP.n24 0.189894
R142 VP.n47 VP.n24 0.189894
R143 VP.n48 VP.n47 0.189894
R144 VP.n49 VP.n48 0.189894
R145 VP.n49 VP.n22 0.189894
R146 VP.n54 VP.n22 0.189894
R147 VP.n55 VP.n54 0.189894
R148 VP.n56 VP.n55 0.189894
R149 VP.n56 VP.n20 0.189894
R150 VP.n60 VP.n20 0.189894
R151 VP.n61 VP.n60 0.189894
R152 VP.n62 VP.n61 0.189894
R153 VP.n62 VP.n18 0.189894
R154 VP.n66 VP.n18 0.189894
R155 VP.n71 VP.n70 0.189894
R156 VP.n71 VP.n15 0.189894
R157 VP.n75 VP.n15 0.189894
R158 VP.n76 VP.n75 0.189894
R159 VP.n77 VP.n76 0.189894
R160 VP.n77 VP.n13 0.189894
R161 VP.n81 VP.n13 0.189894
R162 VP.n82 VP.n81 0.189894
R163 VP.n82 VP.n11 0.189894
R164 VP.n86 VP.n11 0.189894
R165 VP.n87 VP.n86 0.189894
R166 VP.n88 VP.n87 0.189894
R167 VP.n88 VP.n9 0.189894
R168 VP.n92 VP.n9 0.189894
R169 VP.n93 VP.n92 0.189894
R170 VP.n94 VP.n93 0.189894
R171 VP.n94 VP.n7 0.189894
R172 VP.n98 VP.n7 0.189894
R173 VP.n99 VP.n98 0.189894
R174 VP.n100 VP.n99 0.189894
R175 VP.n100 VP.n5 0.189894
R176 VP.n105 VP.n5 0.189894
R177 VP.n106 VP.n105 0.189894
R178 VP.n107 VP.n106 0.189894
R179 VP.n107 VP.n3 0.189894
R180 VP.n111 VP.n3 0.189894
R181 VP.n112 VP.n111 0.189894
R182 VP.n113 VP.n112 0.189894
R183 VP.n113 VP.n1 0.189894
R184 VP.n117 VP.n1 0.189894
R185 VTAIL.n11 VTAIL.t2 45.5998
R186 VTAIL.n17 VTAIL.t3 45.5997
R187 VTAIL.n2 VTAIL.t11 45.5997
R188 VTAIL.n16 VTAIL.t14 45.5997
R189 VTAIL.n15 VTAIL.n14 44.5371
R190 VTAIL.n13 VTAIL.n12 44.5371
R191 VTAIL.n10 VTAIL.n9 44.5371
R192 VTAIL.n8 VTAIL.n7 44.5371
R193 VTAIL.n19 VTAIL.n18 44.5369
R194 VTAIL.n1 VTAIL.n0 44.5369
R195 VTAIL.n4 VTAIL.n3 44.5369
R196 VTAIL.n6 VTAIL.n5 44.5369
R197 VTAIL.n8 VTAIL.n6 35.0479
R198 VTAIL.n17 VTAIL.n16 31.7376
R199 VTAIL.n10 VTAIL.n8 3.31084
R200 VTAIL.n11 VTAIL.n10 3.31084
R201 VTAIL.n15 VTAIL.n13 3.31084
R202 VTAIL.n16 VTAIL.n15 3.31084
R203 VTAIL.n6 VTAIL.n4 3.31084
R204 VTAIL.n4 VTAIL.n2 3.31084
R205 VTAIL.n19 VTAIL.n17 3.31084
R206 VTAIL VTAIL.n1 2.54145
R207 VTAIL.n13 VTAIL.n11 2.1255
R208 VTAIL.n2 VTAIL.n1 2.1255
R209 VTAIL.n18 VTAIL.t6 1.0633
R210 VTAIL.n18 VTAIL.t0 1.0633
R211 VTAIL.n0 VTAIL.t5 1.0633
R212 VTAIL.n0 VTAIL.t8 1.0633
R213 VTAIL.n3 VTAIL.t17 1.0633
R214 VTAIL.n3 VTAIL.t15 1.0633
R215 VTAIL.n5 VTAIL.t13 1.0633
R216 VTAIL.n5 VTAIL.t12 1.0633
R217 VTAIL.n14 VTAIL.t16 1.0633
R218 VTAIL.n14 VTAIL.t10 1.0633
R219 VTAIL.n12 VTAIL.t18 1.0633
R220 VTAIL.n12 VTAIL.t19 1.0633
R221 VTAIL.n9 VTAIL.t4 1.0633
R222 VTAIL.n9 VTAIL.t1 1.0633
R223 VTAIL.n7 VTAIL.t9 1.0633
R224 VTAIL.n7 VTAIL.t7 1.0633
R225 VTAIL VTAIL.n19 0.769897
R226 VDD1.n1 VDD1.t1 65.589
R227 VDD1.n3 VDD1.t5 65.5888
R228 VDD1.n5 VDD1.n4 63.6431
R229 VDD1.n1 VDD1.n0 61.2159
R230 VDD1.n7 VDD1.n6 61.2157
R231 VDD1.n3 VDD1.n2 61.2157
R232 VDD1.n7 VDD1.n5 57.738
R233 VDD1 VDD1.n7 2.42507
R234 VDD1.n6 VDD1.t8 1.0633
R235 VDD1.n6 VDD1.t9 1.0633
R236 VDD1.n0 VDD1.t2 1.0633
R237 VDD1.n0 VDD1.t6 1.0633
R238 VDD1.n4 VDD1.t7 1.0633
R239 VDD1.n4 VDD1.t3 1.0633
R240 VDD1.n2 VDD1.t0 1.0633
R241 VDD1.n2 VDD1.t4 1.0633
R242 VDD1 VDD1.n1 0.886276
R243 VDD1.n5 VDD1.n3 0.77274
R244 B.n1280 B.n1279 585
R245 B.n469 B.n204 585
R246 B.n468 B.n467 585
R247 B.n466 B.n465 585
R248 B.n464 B.n463 585
R249 B.n462 B.n461 585
R250 B.n460 B.n459 585
R251 B.n458 B.n457 585
R252 B.n456 B.n455 585
R253 B.n454 B.n453 585
R254 B.n452 B.n451 585
R255 B.n450 B.n449 585
R256 B.n448 B.n447 585
R257 B.n446 B.n445 585
R258 B.n444 B.n443 585
R259 B.n442 B.n441 585
R260 B.n440 B.n439 585
R261 B.n438 B.n437 585
R262 B.n436 B.n435 585
R263 B.n434 B.n433 585
R264 B.n432 B.n431 585
R265 B.n430 B.n429 585
R266 B.n428 B.n427 585
R267 B.n426 B.n425 585
R268 B.n424 B.n423 585
R269 B.n422 B.n421 585
R270 B.n420 B.n419 585
R271 B.n418 B.n417 585
R272 B.n416 B.n415 585
R273 B.n414 B.n413 585
R274 B.n412 B.n411 585
R275 B.n410 B.n409 585
R276 B.n408 B.n407 585
R277 B.n406 B.n405 585
R278 B.n404 B.n403 585
R279 B.n402 B.n401 585
R280 B.n400 B.n399 585
R281 B.n398 B.n397 585
R282 B.n396 B.n395 585
R283 B.n394 B.n393 585
R284 B.n392 B.n391 585
R285 B.n390 B.n389 585
R286 B.n388 B.n387 585
R287 B.n386 B.n385 585
R288 B.n384 B.n383 585
R289 B.n382 B.n381 585
R290 B.n380 B.n379 585
R291 B.n378 B.n377 585
R292 B.n376 B.n375 585
R293 B.n374 B.n373 585
R294 B.n372 B.n371 585
R295 B.n370 B.n369 585
R296 B.n368 B.n367 585
R297 B.n366 B.n365 585
R298 B.n364 B.n363 585
R299 B.n362 B.n361 585
R300 B.n360 B.n359 585
R301 B.n358 B.n357 585
R302 B.n356 B.n355 585
R303 B.n354 B.n353 585
R304 B.n352 B.n351 585
R305 B.n349 B.n348 585
R306 B.n347 B.n346 585
R307 B.n345 B.n344 585
R308 B.n343 B.n342 585
R309 B.n341 B.n340 585
R310 B.n339 B.n338 585
R311 B.n337 B.n336 585
R312 B.n335 B.n334 585
R313 B.n333 B.n332 585
R314 B.n331 B.n330 585
R315 B.n328 B.n327 585
R316 B.n326 B.n325 585
R317 B.n324 B.n323 585
R318 B.n322 B.n321 585
R319 B.n320 B.n319 585
R320 B.n318 B.n317 585
R321 B.n316 B.n315 585
R322 B.n314 B.n313 585
R323 B.n312 B.n311 585
R324 B.n310 B.n309 585
R325 B.n308 B.n307 585
R326 B.n306 B.n305 585
R327 B.n304 B.n303 585
R328 B.n302 B.n301 585
R329 B.n300 B.n299 585
R330 B.n298 B.n297 585
R331 B.n296 B.n295 585
R332 B.n294 B.n293 585
R333 B.n292 B.n291 585
R334 B.n290 B.n289 585
R335 B.n288 B.n287 585
R336 B.n286 B.n285 585
R337 B.n284 B.n283 585
R338 B.n282 B.n281 585
R339 B.n280 B.n279 585
R340 B.n278 B.n277 585
R341 B.n276 B.n275 585
R342 B.n274 B.n273 585
R343 B.n272 B.n271 585
R344 B.n270 B.n269 585
R345 B.n268 B.n267 585
R346 B.n266 B.n265 585
R347 B.n264 B.n263 585
R348 B.n262 B.n261 585
R349 B.n260 B.n259 585
R350 B.n258 B.n257 585
R351 B.n256 B.n255 585
R352 B.n254 B.n253 585
R353 B.n252 B.n251 585
R354 B.n250 B.n249 585
R355 B.n248 B.n247 585
R356 B.n246 B.n245 585
R357 B.n244 B.n243 585
R358 B.n242 B.n241 585
R359 B.n240 B.n239 585
R360 B.n238 B.n237 585
R361 B.n236 B.n235 585
R362 B.n234 B.n233 585
R363 B.n232 B.n231 585
R364 B.n230 B.n229 585
R365 B.n228 B.n227 585
R366 B.n226 B.n225 585
R367 B.n224 B.n223 585
R368 B.n222 B.n221 585
R369 B.n220 B.n219 585
R370 B.n218 B.n217 585
R371 B.n216 B.n215 585
R372 B.n214 B.n213 585
R373 B.n212 B.n211 585
R374 B.n210 B.n209 585
R375 B.n137 B.n136 585
R376 B.n1278 B.n138 585
R377 B.n1283 B.n138 585
R378 B.n1277 B.n1276 585
R379 B.n1276 B.n134 585
R380 B.n1275 B.n133 585
R381 B.n1289 B.n133 585
R382 B.n1274 B.n132 585
R383 B.n1290 B.n132 585
R384 B.n1273 B.n131 585
R385 B.n1291 B.n131 585
R386 B.n1272 B.n1271 585
R387 B.n1271 B.n127 585
R388 B.n1270 B.n126 585
R389 B.n1297 B.n126 585
R390 B.n1269 B.n125 585
R391 B.n1298 B.n125 585
R392 B.n1268 B.n124 585
R393 B.n1299 B.n124 585
R394 B.n1267 B.n1266 585
R395 B.n1266 B.n123 585
R396 B.n1265 B.n119 585
R397 B.n1305 B.n119 585
R398 B.n1264 B.n118 585
R399 B.n1306 B.n118 585
R400 B.n1263 B.n117 585
R401 B.n1307 B.n117 585
R402 B.n1262 B.n1261 585
R403 B.n1261 B.n113 585
R404 B.n1260 B.n112 585
R405 B.n1313 B.n112 585
R406 B.n1259 B.n111 585
R407 B.n1314 B.n111 585
R408 B.n1258 B.n110 585
R409 B.n1315 B.n110 585
R410 B.n1257 B.n1256 585
R411 B.n1256 B.n106 585
R412 B.n1255 B.n105 585
R413 B.n1321 B.n105 585
R414 B.n1254 B.n104 585
R415 B.n1322 B.n104 585
R416 B.n1253 B.n103 585
R417 B.n1323 B.n103 585
R418 B.n1252 B.n1251 585
R419 B.n1251 B.n99 585
R420 B.n1250 B.n98 585
R421 B.n1329 B.n98 585
R422 B.n1249 B.n97 585
R423 B.n1330 B.n97 585
R424 B.n1248 B.n96 585
R425 B.n1331 B.n96 585
R426 B.n1247 B.n1246 585
R427 B.n1246 B.n92 585
R428 B.n1245 B.n91 585
R429 B.n1337 B.n91 585
R430 B.n1244 B.n90 585
R431 B.n1338 B.n90 585
R432 B.n1243 B.n89 585
R433 B.n1339 B.n89 585
R434 B.n1242 B.n1241 585
R435 B.n1241 B.n85 585
R436 B.n1240 B.n84 585
R437 B.n1345 B.n84 585
R438 B.n1239 B.n83 585
R439 B.n1346 B.n83 585
R440 B.n1238 B.n82 585
R441 B.n1347 B.n82 585
R442 B.n1237 B.n1236 585
R443 B.n1236 B.n78 585
R444 B.n1235 B.n77 585
R445 B.n1353 B.n77 585
R446 B.n1234 B.n76 585
R447 B.n1354 B.n76 585
R448 B.n1233 B.n75 585
R449 B.n1355 B.n75 585
R450 B.n1232 B.n1231 585
R451 B.n1231 B.n71 585
R452 B.n1230 B.n70 585
R453 B.n1361 B.n70 585
R454 B.n1229 B.n69 585
R455 B.n1362 B.n69 585
R456 B.n1228 B.n68 585
R457 B.n1363 B.n68 585
R458 B.n1227 B.n1226 585
R459 B.n1226 B.n64 585
R460 B.n1225 B.n63 585
R461 B.n1369 B.n63 585
R462 B.n1224 B.n62 585
R463 B.n1370 B.n62 585
R464 B.n1223 B.n61 585
R465 B.n1371 B.n61 585
R466 B.n1222 B.n1221 585
R467 B.n1221 B.n57 585
R468 B.n1220 B.n56 585
R469 B.n1377 B.n56 585
R470 B.n1219 B.n55 585
R471 B.n1378 B.n55 585
R472 B.n1218 B.n54 585
R473 B.n1379 B.n54 585
R474 B.n1217 B.n1216 585
R475 B.n1216 B.n50 585
R476 B.n1215 B.n49 585
R477 B.n1385 B.n49 585
R478 B.n1214 B.n48 585
R479 B.n1386 B.n48 585
R480 B.n1213 B.n47 585
R481 B.n1387 B.n47 585
R482 B.n1212 B.n1211 585
R483 B.n1211 B.n43 585
R484 B.n1210 B.n42 585
R485 B.n1393 B.n42 585
R486 B.n1209 B.n41 585
R487 B.n1394 B.n41 585
R488 B.n1208 B.n40 585
R489 B.n1395 B.n40 585
R490 B.n1207 B.n1206 585
R491 B.n1206 B.n39 585
R492 B.n1205 B.n35 585
R493 B.n1401 B.n35 585
R494 B.n1204 B.n34 585
R495 B.n1402 B.n34 585
R496 B.n1203 B.n33 585
R497 B.n1403 B.n33 585
R498 B.n1202 B.n1201 585
R499 B.n1201 B.n29 585
R500 B.n1200 B.n28 585
R501 B.n1409 B.n28 585
R502 B.n1199 B.n27 585
R503 B.n1410 B.n27 585
R504 B.n1198 B.n26 585
R505 B.n1411 B.n26 585
R506 B.n1197 B.n1196 585
R507 B.n1196 B.n22 585
R508 B.n1195 B.n21 585
R509 B.n1417 B.n21 585
R510 B.n1194 B.n20 585
R511 B.n1418 B.n20 585
R512 B.n1193 B.n19 585
R513 B.n1419 B.n19 585
R514 B.n1192 B.n1191 585
R515 B.n1191 B.n15 585
R516 B.n1190 B.n14 585
R517 B.n1425 B.n14 585
R518 B.n1189 B.n13 585
R519 B.n1426 B.n13 585
R520 B.n1188 B.n12 585
R521 B.n1427 B.n12 585
R522 B.n1187 B.n1186 585
R523 B.n1186 B.n8 585
R524 B.n1185 B.n7 585
R525 B.n1433 B.n7 585
R526 B.n1184 B.n6 585
R527 B.n1434 B.n6 585
R528 B.n1183 B.n5 585
R529 B.n1435 B.n5 585
R530 B.n1182 B.n1181 585
R531 B.n1181 B.n4 585
R532 B.n1180 B.n470 585
R533 B.n1180 B.n1179 585
R534 B.n1170 B.n471 585
R535 B.n472 B.n471 585
R536 B.n1172 B.n1171 585
R537 B.n1173 B.n1172 585
R538 B.n1169 B.n477 585
R539 B.n477 B.n476 585
R540 B.n1168 B.n1167 585
R541 B.n1167 B.n1166 585
R542 B.n479 B.n478 585
R543 B.n480 B.n479 585
R544 B.n1159 B.n1158 585
R545 B.n1160 B.n1159 585
R546 B.n1157 B.n485 585
R547 B.n485 B.n484 585
R548 B.n1156 B.n1155 585
R549 B.n1155 B.n1154 585
R550 B.n487 B.n486 585
R551 B.n488 B.n487 585
R552 B.n1147 B.n1146 585
R553 B.n1148 B.n1147 585
R554 B.n1145 B.n493 585
R555 B.n493 B.n492 585
R556 B.n1144 B.n1143 585
R557 B.n1143 B.n1142 585
R558 B.n495 B.n494 585
R559 B.n496 B.n495 585
R560 B.n1135 B.n1134 585
R561 B.n1136 B.n1135 585
R562 B.n1133 B.n501 585
R563 B.n501 B.n500 585
R564 B.n1132 B.n1131 585
R565 B.n1131 B.n1130 585
R566 B.n503 B.n502 585
R567 B.n1123 B.n503 585
R568 B.n1122 B.n1121 585
R569 B.n1124 B.n1122 585
R570 B.n1120 B.n508 585
R571 B.n508 B.n507 585
R572 B.n1119 B.n1118 585
R573 B.n1118 B.n1117 585
R574 B.n510 B.n509 585
R575 B.n511 B.n510 585
R576 B.n1110 B.n1109 585
R577 B.n1111 B.n1110 585
R578 B.n1108 B.n516 585
R579 B.n516 B.n515 585
R580 B.n1107 B.n1106 585
R581 B.n1106 B.n1105 585
R582 B.n518 B.n517 585
R583 B.n519 B.n518 585
R584 B.n1098 B.n1097 585
R585 B.n1099 B.n1098 585
R586 B.n1096 B.n524 585
R587 B.n524 B.n523 585
R588 B.n1095 B.n1094 585
R589 B.n1094 B.n1093 585
R590 B.n526 B.n525 585
R591 B.n527 B.n526 585
R592 B.n1086 B.n1085 585
R593 B.n1087 B.n1086 585
R594 B.n1084 B.n532 585
R595 B.n532 B.n531 585
R596 B.n1083 B.n1082 585
R597 B.n1082 B.n1081 585
R598 B.n534 B.n533 585
R599 B.n535 B.n534 585
R600 B.n1074 B.n1073 585
R601 B.n1075 B.n1074 585
R602 B.n1072 B.n540 585
R603 B.n540 B.n539 585
R604 B.n1071 B.n1070 585
R605 B.n1070 B.n1069 585
R606 B.n542 B.n541 585
R607 B.n543 B.n542 585
R608 B.n1062 B.n1061 585
R609 B.n1063 B.n1062 585
R610 B.n1060 B.n548 585
R611 B.n548 B.n547 585
R612 B.n1059 B.n1058 585
R613 B.n1058 B.n1057 585
R614 B.n550 B.n549 585
R615 B.n551 B.n550 585
R616 B.n1050 B.n1049 585
R617 B.n1051 B.n1050 585
R618 B.n1048 B.n556 585
R619 B.n556 B.n555 585
R620 B.n1047 B.n1046 585
R621 B.n1046 B.n1045 585
R622 B.n558 B.n557 585
R623 B.n559 B.n558 585
R624 B.n1038 B.n1037 585
R625 B.n1039 B.n1038 585
R626 B.n1036 B.n564 585
R627 B.n564 B.n563 585
R628 B.n1035 B.n1034 585
R629 B.n1034 B.n1033 585
R630 B.n566 B.n565 585
R631 B.n567 B.n566 585
R632 B.n1026 B.n1025 585
R633 B.n1027 B.n1026 585
R634 B.n1024 B.n571 585
R635 B.n575 B.n571 585
R636 B.n1023 B.n1022 585
R637 B.n1022 B.n1021 585
R638 B.n573 B.n572 585
R639 B.n574 B.n573 585
R640 B.n1014 B.n1013 585
R641 B.n1015 B.n1014 585
R642 B.n1012 B.n580 585
R643 B.n580 B.n579 585
R644 B.n1011 B.n1010 585
R645 B.n1010 B.n1009 585
R646 B.n582 B.n581 585
R647 B.n583 B.n582 585
R648 B.n1002 B.n1001 585
R649 B.n1003 B.n1002 585
R650 B.n1000 B.n588 585
R651 B.n588 B.n587 585
R652 B.n999 B.n998 585
R653 B.n998 B.n997 585
R654 B.n590 B.n589 585
R655 B.n591 B.n590 585
R656 B.n990 B.n989 585
R657 B.n991 B.n990 585
R658 B.n988 B.n596 585
R659 B.n596 B.n595 585
R660 B.n987 B.n986 585
R661 B.n986 B.n985 585
R662 B.n598 B.n597 585
R663 B.n978 B.n598 585
R664 B.n977 B.n976 585
R665 B.n979 B.n977 585
R666 B.n975 B.n603 585
R667 B.n603 B.n602 585
R668 B.n974 B.n973 585
R669 B.n973 B.n972 585
R670 B.n605 B.n604 585
R671 B.n606 B.n605 585
R672 B.n965 B.n964 585
R673 B.n966 B.n965 585
R674 B.n963 B.n611 585
R675 B.n611 B.n610 585
R676 B.n962 B.n961 585
R677 B.n961 B.n960 585
R678 B.n613 B.n612 585
R679 B.n614 B.n613 585
R680 B.n953 B.n952 585
R681 B.n954 B.n953 585
R682 B.n617 B.n616 585
R683 B.n692 B.n691 585
R684 B.n693 B.n689 585
R685 B.n689 B.n618 585
R686 B.n695 B.n694 585
R687 B.n697 B.n688 585
R688 B.n700 B.n699 585
R689 B.n701 B.n687 585
R690 B.n703 B.n702 585
R691 B.n705 B.n686 585
R692 B.n708 B.n707 585
R693 B.n709 B.n685 585
R694 B.n711 B.n710 585
R695 B.n713 B.n684 585
R696 B.n716 B.n715 585
R697 B.n717 B.n683 585
R698 B.n719 B.n718 585
R699 B.n721 B.n682 585
R700 B.n724 B.n723 585
R701 B.n725 B.n681 585
R702 B.n727 B.n726 585
R703 B.n729 B.n680 585
R704 B.n732 B.n731 585
R705 B.n733 B.n679 585
R706 B.n735 B.n734 585
R707 B.n737 B.n678 585
R708 B.n740 B.n739 585
R709 B.n741 B.n677 585
R710 B.n743 B.n742 585
R711 B.n745 B.n676 585
R712 B.n748 B.n747 585
R713 B.n749 B.n675 585
R714 B.n751 B.n750 585
R715 B.n753 B.n674 585
R716 B.n756 B.n755 585
R717 B.n757 B.n673 585
R718 B.n759 B.n758 585
R719 B.n761 B.n672 585
R720 B.n764 B.n763 585
R721 B.n765 B.n671 585
R722 B.n767 B.n766 585
R723 B.n769 B.n670 585
R724 B.n772 B.n771 585
R725 B.n773 B.n669 585
R726 B.n775 B.n774 585
R727 B.n777 B.n668 585
R728 B.n780 B.n779 585
R729 B.n781 B.n667 585
R730 B.n783 B.n782 585
R731 B.n785 B.n666 585
R732 B.n788 B.n787 585
R733 B.n789 B.n665 585
R734 B.n791 B.n790 585
R735 B.n793 B.n664 585
R736 B.n796 B.n795 585
R737 B.n797 B.n663 585
R738 B.n799 B.n798 585
R739 B.n801 B.n662 585
R740 B.n804 B.n803 585
R741 B.n805 B.n661 585
R742 B.n807 B.n806 585
R743 B.n809 B.n660 585
R744 B.n812 B.n811 585
R745 B.n813 B.n656 585
R746 B.n815 B.n814 585
R747 B.n817 B.n655 585
R748 B.n820 B.n819 585
R749 B.n821 B.n654 585
R750 B.n823 B.n822 585
R751 B.n825 B.n653 585
R752 B.n828 B.n827 585
R753 B.n829 B.n650 585
R754 B.n832 B.n831 585
R755 B.n834 B.n649 585
R756 B.n837 B.n836 585
R757 B.n838 B.n648 585
R758 B.n840 B.n839 585
R759 B.n842 B.n647 585
R760 B.n845 B.n844 585
R761 B.n846 B.n646 585
R762 B.n848 B.n847 585
R763 B.n850 B.n645 585
R764 B.n853 B.n852 585
R765 B.n854 B.n644 585
R766 B.n856 B.n855 585
R767 B.n858 B.n643 585
R768 B.n861 B.n860 585
R769 B.n862 B.n642 585
R770 B.n864 B.n863 585
R771 B.n866 B.n641 585
R772 B.n869 B.n868 585
R773 B.n870 B.n640 585
R774 B.n872 B.n871 585
R775 B.n874 B.n639 585
R776 B.n877 B.n876 585
R777 B.n878 B.n638 585
R778 B.n880 B.n879 585
R779 B.n882 B.n637 585
R780 B.n885 B.n884 585
R781 B.n886 B.n636 585
R782 B.n888 B.n887 585
R783 B.n890 B.n635 585
R784 B.n893 B.n892 585
R785 B.n894 B.n634 585
R786 B.n896 B.n895 585
R787 B.n898 B.n633 585
R788 B.n901 B.n900 585
R789 B.n902 B.n632 585
R790 B.n904 B.n903 585
R791 B.n906 B.n631 585
R792 B.n909 B.n908 585
R793 B.n910 B.n630 585
R794 B.n912 B.n911 585
R795 B.n914 B.n629 585
R796 B.n917 B.n916 585
R797 B.n918 B.n628 585
R798 B.n920 B.n919 585
R799 B.n922 B.n627 585
R800 B.n925 B.n924 585
R801 B.n926 B.n626 585
R802 B.n928 B.n927 585
R803 B.n930 B.n625 585
R804 B.n933 B.n932 585
R805 B.n934 B.n624 585
R806 B.n936 B.n935 585
R807 B.n938 B.n623 585
R808 B.n941 B.n940 585
R809 B.n942 B.n622 585
R810 B.n944 B.n943 585
R811 B.n946 B.n621 585
R812 B.n947 B.n620 585
R813 B.n950 B.n949 585
R814 B.n951 B.n619 585
R815 B.n619 B.n618 585
R816 B.n956 B.n955 585
R817 B.n955 B.n954 585
R818 B.n957 B.n615 585
R819 B.n615 B.n614 585
R820 B.n959 B.n958 585
R821 B.n960 B.n959 585
R822 B.n609 B.n608 585
R823 B.n610 B.n609 585
R824 B.n968 B.n967 585
R825 B.n967 B.n966 585
R826 B.n969 B.n607 585
R827 B.n607 B.n606 585
R828 B.n971 B.n970 585
R829 B.n972 B.n971 585
R830 B.n601 B.n600 585
R831 B.n602 B.n601 585
R832 B.n981 B.n980 585
R833 B.n980 B.n979 585
R834 B.n982 B.n599 585
R835 B.n978 B.n599 585
R836 B.n984 B.n983 585
R837 B.n985 B.n984 585
R838 B.n594 B.n593 585
R839 B.n595 B.n594 585
R840 B.n993 B.n992 585
R841 B.n992 B.n991 585
R842 B.n994 B.n592 585
R843 B.n592 B.n591 585
R844 B.n996 B.n995 585
R845 B.n997 B.n996 585
R846 B.n586 B.n585 585
R847 B.n587 B.n586 585
R848 B.n1005 B.n1004 585
R849 B.n1004 B.n1003 585
R850 B.n1006 B.n584 585
R851 B.n584 B.n583 585
R852 B.n1008 B.n1007 585
R853 B.n1009 B.n1008 585
R854 B.n578 B.n577 585
R855 B.n579 B.n578 585
R856 B.n1017 B.n1016 585
R857 B.n1016 B.n1015 585
R858 B.n1018 B.n576 585
R859 B.n576 B.n574 585
R860 B.n1020 B.n1019 585
R861 B.n1021 B.n1020 585
R862 B.n570 B.n569 585
R863 B.n575 B.n570 585
R864 B.n1029 B.n1028 585
R865 B.n1028 B.n1027 585
R866 B.n1030 B.n568 585
R867 B.n568 B.n567 585
R868 B.n1032 B.n1031 585
R869 B.n1033 B.n1032 585
R870 B.n562 B.n561 585
R871 B.n563 B.n562 585
R872 B.n1041 B.n1040 585
R873 B.n1040 B.n1039 585
R874 B.n1042 B.n560 585
R875 B.n560 B.n559 585
R876 B.n1044 B.n1043 585
R877 B.n1045 B.n1044 585
R878 B.n554 B.n553 585
R879 B.n555 B.n554 585
R880 B.n1053 B.n1052 585
R881 B.n1052 B.n1051 585
R882 B.n1054 B.n552 585
R883 B.n552 B.n551 585
R884 B.n1056 B.n1055 585
R885 B.n1057 B.n1056 585
R886 B.n546 B.n545 585
R887 B.n547 B.n546 585
R888 B.n1065 B.n1064 585
R889 B.n1064 B.n1063 585
R890 B.n1066 B.n544 585
R891 B.n544 B.n543 585
R892 B.n1068 B.n1067 585
R893 B.n1069 B.n1068 585
R894 B.n538 B.n537 585
R895 B.n539 B.n538 585
R896 B.n1077 B.n1076 585
R897 B.n1076 B.n1075 585
R898 B.n1078 B.n536 585
R899 B.n536 B.n535 585
R900 B.n1080 B.n1079 585
R901 B.n1081 B.n1080 585
R902 B.n530 B.n529 585
R903 B.n531 B.n530 585
R904 B.n1089 B.n1088 585
R905 B.n1088 B.n1087 585
R906 B.n1090 B.n528 585
R907 B.n528 B.n527 585
R908 B.n1092 B.n1091 585
R909 B.n1093 B.n1092 585
R910 B.n522 B.n521 585
R911 B.n523 B.n522 585
R912 B.n1101 B.n1100 585
R913 B.n1100 B.n1099 585
R914 B.n1102 B.n520 585
R915 B.n520 B.n519 585
R916 B.n1104 B.n1103 585
R917 B.n1105 B.n1104 585
R918 B.n514 B.n513 585
R919 B.n515 B.n514 585
R920 B.n1113 B.n1112 585
R921 B.n1112 B.n1111 585
R922 B.n1114 B.n512 585
R923 B.n512 B.n511 585
R924 B.n1116 B.n1115 585
R925 B.n1117 B.n1116 585
R926 B.n506 B.n505 585
R927 B.n507 B.n506 585
R928 B.n1126 B.n1125 585
R929 B.n1125 B.n1124 585
R930 B.n1127 B.n504 585
R931 B.n1123 B.n504 585
R932 B.n1129 B.n1128 585
R933 B.n1130 B.n1129 585
R934 B.n499 B.n498 585
R935 B.n500 B.n499 585
R936 B.n1138 B.n1137 585
R937 B.n1137 B.n1136 585
R938 B.n1139 B.n497 585
R939 B.n497 B.n496 585
R940 B.n1141 B.n1140 585
R941 B.n1142 B.n1141 585
R942 B.n491 B.n490 585
R943 B.n492 B.n491 585
R944 B.n1150 B.n1149 585
R945 B.n1149 B.n1148 585
R946 B.n1151 B.n489 585
R947 B.n489 B.n488 585
R948 B.n1153 B.n1152 585
R949 B.n1154 B.n1153 585
R950 B.n483 B.n482 585
R951 B.n484 B.n483 585
R952 B.n1162 B.n1161 585
R953 B.n1161 B.n1160 585
R954 B.n1163 B.n481 585
R955 B.n481 B.n480 585
R956 B.n1165 B.n1164 585
R957 B.n1166 B.n1165 585
R958 B.n475 B.n474 585
R959 B.n476 B.n475 585
R960 B.n1175 B.n1174 585
R961 B.n1174 B.n1173 585
R962 B.n1176 B.n473 585
R963 B.n473 B.n472 585
R964 B.n1178 B.n1177 585
R965 B.n1179 B.n1178 585
R966 B.n2 B.n0 585
R967 B.n4 B.n2 585
R968 B.n3 B.n1 585
R969 B.n1434 B.n3 585
R970 B.n1432 B.n1431 585
R971 B.n1433 B.n1432 585
R972 B.n1430 B.n9 585
R973 B.n9 B.n8 585
R974 B.n1429 B.n1428 585
R975 B.n1428 B.n1427 585
R976 B.n11 B.n10 585
R977 B.n1426 B.n11 585
R978 B.n1424 B.n1423 585
R979 B.n1425 B.n1424 585
R980 B.n1422 B.n16 585
R981 B.n16 B.n15 585
R982 B.n1421 B.n1420 585
R983 B.n1420 B.n1419 585
R984 B.n18 B.n17 585
R985 B.n1418 B.n18 585
R986 B.n1416 B.n1415 585
R987 B.n1417 B.n1416 585
R988 B.n1414 B.n23 585
R989 B.n23 B.n22 585
R990 B.n1413 B.n1412 585
R991 B.n1412 B.n1411 585
R992 B.n25 B.n24 585
R993 B.n1410 B.n25 585
R994 B.n1408 B.n1407 585
R995 B.n1409 B.n1408 585
R996 B.n1406 B.n30 585
R997 B.n30 B.n29 585
R998 B.n1405 B.n1404 585
R999 B.n1404 B.n1403 585
R1000 B.n32 B.n31 585
R1001 B.n1402 B.n32 585
R1002 B.n1400 B.n1399 585
R1003 B.n1401 B.n1400 585
R1004 B.n1398 B.n36 585
R1005 B.n39 B.n36 585
R1006 B.n1397 B.n1396 585
R1007 B.n1396 B.n1395 585
R1008 B.n38 B.n37 585
R1009 B.n1394 B.n38 585
R1010 B.n1392 B.n1391 585
R1011 B.n1393 B.n1392 585
R1012 B.n1390 B.n44 585
R1013 B.n44 B.n43 585
R1014 B.n1389 B.n1388 585
R1015 B.n1388 B.n1387 585
R1016 B.n46 B.n45 585
R1017 B.n1386 B.n46 585
R1018 B.n1384 B.n1383 585
R1019 B.n1385 B.n1384 585
R1020 B.n1382 B.n51 585
R1021 B.n51 B.n50 585
R1022 B.n1381 B.n1380 585
R1023 B.n1380 B.n1379 585
R1024 B.n53 B.n52 585
R1025 B.n1378 B.n53 585
R1026 B.n1376 B.n1375 585
R1027 B.n1377 B.n1376 585
R1028 B.n1374 B.n58 585
R1029 B.n58 B.n57 585
R1030 B.n1373 B.n1372 585
R1031 B.n1372 B.n1371 585
R1032 B.n60 B.n59 585
R1033 B.n1370 B.n60 585
R1034 B.n1368 B.n1367 585
R1035 B.n1369 B.n1368 585
R1036 B.n1366 B.n65 585
R1037 B.n65 B.n64 585
R1038 B.n1365 B.n1364 585
R1039 B.n1364 B.n1363 585
R1040 B.n67 B.n66 585
R1041 B.n1362 B.n67 585
R1042 B.n1360 B.n1359 585
R1043 B.n1361 B.n1360 585
R1044 B.n1358 B.n72 585
R1045 B.n72 B.n71 585
R1046 B.n1357 B.n1356 585
R1047 B.n1356 B.n1355 585
R1048 B.n74 B.n73 585
R1049 B.n1354 B.n74 585
R1050 B.n1352 B.n1351 585
R1051 B.n1353 B.n1352 585
R1052 B.n1350 B.n79 585
R1053 B.n79 B.n78 585
R1054 B.n1349 B.n1348 585
R1055 B.n1348 B.n1347 585
R1056 B.n81 B.n80 585
R1057 B.n1346 B.n81 585
R1058 B.n1344 B.n1343 585
R1059 B.n1345 B.n1344 585
R1060 B.n1342 B.n86 585
R1061 B.n86 B.n85 585
R1062 B.n1341 B.n1340 585
R1063 B.n1340 B.n1339 585
R1064 B.n88 B.n87 585
R1065 B.n1338 B.n88 585
R1066 B.n1336 B.n1335 585
R1067 B.n1337 B.n1336 585
R1068 B.n1334 B.n93 585
R1069 B.n93 B.n92 585
R1070 B.n1333 B.n1332 585
R1071 B.n1332 B.n1331 585
R1072 B.n95 B.n94 585
R1073 B.n1330 B.n95 585
R1074 B.n1328 B.n1327 585
R1075 B.n1329 B.n1328 585
R1076 B.n1326 B.n100 585
R1077 B.n100 B.n99 585
R1078 B.n1325 B.n1324 585
R1079 B.n1324 B.n1323 585
R1080 B.n102 B.n101 585
R1081 B.n1322 B.n102 585
R1082 B.n1320 B.n1319 585
R1083 B.n1321 B.n1320 585
R1084 B.n1318 B.n107 585
R1085 B.n107 B.n106 585
R1086 B.n1317 B.n1316 585
R1087 B.n1316 B.n1315 585
R1088 B.n109 B.n108 585
R1089 B.n1314 B.n109 585
R1090 B.n1312 B.n1311 585
R1091 B.n1313 B.n1312 585
R1092 B.n1310 B.n114 585
R1093 B.n114 B.n113 585
R1094 B.n1309 B.n1308 585
R1095 B.n1308 B.n1307 585
R1096 B.n116 B.n115 585
R1097 B.n1306 B.n116 585
R1098 B.n1304 B.n1303 585
R1099 B.n1305 B.n1304 585
R1100 B.n1302 B.n120 585
R1101 B.n123 B.n120 585
R1102 B.n1301 B.n1300 585
R1103 B.n1300 B.n1299 585
R1104 B.n122 B.n121 585
R1105 B.n1298 B.n122 585
R1106 B.n1296 B.n1295 585
R1107 B.n1297 B.n1296 585
R1108 B.n1294 B.n128 585
R1109 B.n128 B.n127 585
R1110 B.n1293 B.n1292 585
R1111 B.n1292 B.n1291 585
R1112 B.n130 B.n129 585
R1113 B.n1290 B.n130 585
R1114 B.n1288 B.n1287 585
R1115 B.n1289 B.n1288 585
R1116 B.n1286 B.n135 585
R1117 B.n135 B.n134 585
R1118 B.n1285 B.n1284 585
R1119 B.n1284 B.n1283 585
R1120 B.n1437 B.n1436 585
R1121 B.n1436 B.n1435 585
R1122 B.n955 B.n617 463.671
R1123 B.n1284 B.n137 463.671
R1124 B.n953 B.n619 463.671
R1125 B.n1280 B.n138 463.671
R1126 B.n651 B.t14 337.019
R1127 B.n657 B.t18 337.019
R1128 B.n207 B.t21 337.019
R1129 B.n205 B.t10 337.019
R1130 B.n1282 B.n1281 256.663
R1131 B.n1282 B.n203 256.663
R1132 B.n1282 B.n202 256.663
R1133 B.n1282 B.n201 256.663
R1134 B.n1282 B.n200 256.663
R1135 B.n1282 B.n199 256.663
R1136 B.n1282 B.n198 256.663
R1137 B.n1282 B.n197 256.663
R1138 B.n1282 B.n196 256.663
R1139 B.n1282 B.n195 256.663
R1140 B.n1282 B.n194 256.663
R1141 B.n1282 B.n193 256.663
R1142 B.n1282 B.n192 256.663
R1143 B.n1282 B.n191 256.663
R1144 B.n1282 B.n190 256.663
R1145 B.n1282 B.n189 256.663
R1146 B.n1282 B.n188 256.663
R1147 B.n1282 B.n187 256.663
R1148 B.n1282 B.n186 256.663
R1149 B.n1282 B.n185 256.663
R1150 B.n1282 B.n184 256.663
R1151 B.n1282 B.n183 256.663
R1152 B.n1282 B.n182 256.663
R1153 B.n1282 B.n181 256.663
R1154 B.n1282 B.n180 256.663
R1155 B.n1282 B.n179 256.663
R1156 B.n1282 B.n178 256.663
R1157 B.n1282 B.n177 256.663
R1158 B.n1282 B.n176 256.663
R1159 B.n1282 B.n175 256.663
R1160 B.n1282 B.n174 256.663
R1161 B.n1282 B.n173 256.663
R1162 B.n1282 B.n172 256.663
R1163 B.n1282 B.n171 256.663
R1164 B.n1282 B.n170 256.663
R1165 B.n1282 B.n169 256.663
R1166 B.n1282 B.n168 256.663
R1167 B.n1282 B.n167 256.663
R1168 B.n1282 B.n166 256.663
R1169 B.n1282 B.n165 256.663
R1170 B.n1282 B.n164 256.663
R1171 B.n1282 B.n163 256.663
R1172 B.n1282 B.n162 256.663
R1173 B.n1282 B.n161 256.663
R1174 B.n1282 B.n160 256.663
R1175 B.n1282 B.n159 256.663
R1176 B.n1282 B.n158 256.663
R1177 B.n1282 B.n157 256.663
R1178 B.n1282 B.n156 256.663
R1179 B.n1282 B.n155 256.663
R1180 B.n1282 B.n154 256.663
R1181 B.n1282 B.n153 256.663
R1182 B.n1282 B.n152 256.663
R1183 B.n1282 B.n151 256.663
R1184 B.n1282 B.n150 256.663
R1185 B.n1282 B.n149 256.663
R1186 B.n1282 B.n148 256.663
R1187 B.n1282 B.n147 256.663
R1188 B.n1282 B.n146 256.663
R1189 B.n1282 B.n145 256.663
R1190 B.n1282 B.n144 256.663
R1191 B.n1282 B.n143 256.663
R1192 B.n1282 B.n142 256.663
R1193 B.n1282 B.n141 256.663
R1194 B.n1282 B.n140 256.663
R1195 B.n1282 B.n139 256.663
R1196 B.n690 B.n618 256.663
R1197 B.n696 B.n618 256.663
R1198 B.n698 B.n618 256.663
R1199 B.n704 B.n618 256.663
R1200 B.n706 B.n618 256.663
R1201 B.n712 B.n618 256.663
R1202 B.n714 B.n618 256.663
R1203 B.n720 B.n618 256.663
R1204 B.n722 B.n618 256.663
R1205 B.n728 B.n618 256.663
R1206 B.n730 B.n618 256.663
R1207 B.n736 B.n618 256.663
R1208 B.n738 B.n618 256.663
R1209 B.n744 B.n618 256.663
R1210 B.n746 B.n618 256.663
R1211 B.n752 B.n618 256.663
R1212 B.n754 B.n618 256.663
R1213 B.n760 B.n618 256.663
R1214 B.n762 B.n618 256.663
R1215 B.n768 B.n618 256.663
R1216 B.n770 B.n618 256.663
R1217 B.n776 B.n618 256.663
R1218 B.n778 B.n618 256.663
R1219 B.n784 B.n618 256.663
R1220 B.n786 B.n618 256.663
R1221 B.n792 B.n618 256.663
R1222 B.n794 B.n618 256.663
R1223 B.n800 B.n618 256.663
R1224 B.n802 B.n618 256.663
R1225 B.n808 B.n618 256.663
R1226 B.n810 B.n618 256.663
R1227 B.n816 B.n618 256.663
R1228 B.n818 B.n618 256.663
R1229 B.n824 B.n618 256.663
R1230 B.n826 B.n618 256.663
R1231 B.n833 B.n618 256.663
R1232 B.n835 B.n618 256.663
R1233 B.n841 B.n618 256.663
R1234 B.n843 B.n618 256.663
R1235 B.n849 B.n618 256.663
R1236 B.n851 B.n618 256.663
R1237 B.n857 B.n618 256.663
R1238 B.n859 B.n618 256.663
R1239 B.n865 B.n618 256.663
R1240 B.n867 B.n618 256.663
R1241 B.n873 B.n618 256.663
R1242 B.n875 B.n618 256.663
R1243 B.n881 B.n618 256.663
R1244 B.n883 B.n618 256.663
R1245 B.n889 B.n618 256.663
R1246 B.n891 B.n618 256.663
R1247 B.n897 B.n618 256.663
R1248 B.n899 B.n618 256.663
R1249 B.n905 B.n618 256.663
R1250 B.n907 B.n618 256.663
R1251 B.n913 B.n618 256.663
R1252 B.n915 B.n618 256.663
R1253 B.n921 B.n618 256.663
R1254 B.n923 B.n618 256.663
R1255 B.n929 B.n618 256.663
R1256 B.n931 B.n618 256.663
R1257 B.n937 B.n618 256.663
R1258 B.n939 B.n618 256.663
R1259 B.n945 B.n618 256.663
R1260 B.n948 B.n618 256.663
R1261 B.n955 B.n615 163.367
R1262 B.n959 B.n615 163.367
R1263 B.n959 B.n609 163.367
R1264 B.n967 B.n609 163.367
R1265 B.n967 B.n607 163.367
R1266 B.n971 B.n607 163.367
R1267 B.n971 B.n601 163.367
R1268 B.n980 B.n601 163.367
R1269 B.n980 B.n599 163.367
R1270 B.n984 B.n599 163.367
R1271 B.n984 B.n594 163.367
R1272 B.n992 B.n594 163.367
R1273 B.n992 B.n592 163.367
R1274 B.n996 B.n592 163.367
R1275 B.n996 B.n586 163.367
R1276 B.n1004 B.n586 163.367
R1277 B.n1004 B.n584 163.367
R1278 B.n1008 B.n584 163.367
R1279 B.n1008 B.n578 163.367
R1280 B.n1016 B.n578 163.367
R1281 B.n1016 B.n576 163.367
R1282 B.n1020 B.n576 163.367
R1283 B.n1020 B.n570 163.367
R1284 B.n1028 B.n570 163.367
R1285 B.n1028 B.n568 163.367
R1286 B.n1032 B.n568 163.367
R1287 B.n1032 B.n562 163.367
R1288 B.n1040 B.n562 163.367
R1289 B.n1040 B.n560 163.367
R1290 B.n1044 B.n560 163.367
R1291 B.n1044 B.n554 163.367
R1292 B.n1052 B.n554 163.367
R1293 B.n1052 B.n552 163.367
R1294 B.n1056 B.n552 163.367
R1295 B.n1056 B.n546 163.367
R1296 B.n1064 B.n546 163.367
R1297 B.n1064 B.n544 163.367
R1298 B.n1068 B.n544 163.367
R1299 B.n1068 B.n538 163.367
R1300 B.n1076 B.n538 163.367
R1301 B.n1076 B.n536 163.367
R1302 B.n1080 B.n536 163.367
R1303 B.n1080 B.n530 163.367
R1304 B.n1088 B.n530 163.367
R1305 B.n1088 B.n528 163.367
R1306 B.n1092 B.n528 163.367
R1307 B.n1092 B.n522 163.367
R1308 B.n1100 B.n522 163.367
R1309 B.n1100 B.n520 163.367
R1310 B.n1104 B.n520 163.367
R1311 B.n1104 B.n514 163.367
R1312 B.n1112 B.n514 163.367
R1313 B.n1112 B.n512 163.367
R1314 B.n1116 B.n512 163.367
R1315 B.n1116 B.n506 163.367
R1316 B.n1125 B.n506 163.367
R1317 B.n1125 B.n504 163.367
R1318 B.n1129 B.n504 163.367
R1319 B.n1129 B.n499 163.367
R1320 B.n1137 B.n499 163.367
R1321 B.n1137 B.n497 163.367
R1322 B.n1141 B.n497 163.367
R1323 B.n1141 B.n491 163.367
R1324 B.n1149 B.n491 163.367
R1325 B.n1149 B.n489 163.367
R1326 B.n1153 B.n489 163.367
R1327 B.n1153 B.n483 163.367
R1328 B.n1161 B.n483 163.367
R1329 B.n1161 B.n481 163.367
R1330 B.n1165 B.n481 163.367
R1331 B.n1165 B.n475 163.367
R1332 B.n1174 B.n475 163.367
R1333 B.n1174 B.n473 163.367
R1334 B.n1178 B.n473 163.367
R1335 B.n1178 B.n2 163.367
R1336 B.n1436 B.n2 163.367
R1337 B.n1436 B.n3 163.367
R1338 B.n1432 B.n3 163.367
R1339 B.n1432 B.n9 163.367
R1340 B.n1428 B.n9 163.367
R1341 B.n1428 B.n11 163.367
R1342 B.n1424 B.n11 163.367
R1343 B.n1424 B.n16 163.367
R1344 B.n1420 B.n16 163.367
R1345 B.n1420 B.n18 163.367
R1346 B.n1416 B.n18 163.367
R1347 B.n1416 B.n23 163.367
R1348 B.n1412 B.n23 163.367
R1349 B.n1412 B.n25 163.367
R1350 B.n1408 B.n25 163.367
R1351 B.n1408 B.n30 163.367
R1352 B.n1404 B.n30 163.367
R1353 B.n1404 B.n32 163.367
R1354 B.n1400 B.n32 163.367
R1355 B.n1400 B.n36 163.367
R1356 B.n1396 B.n36 163.367
R1357 B.n1396 B.n38 163.367
R1358 B.n1392 B.n38 163.367
R1359 B.n1392 B.n44 163.367
R1360 B.n1388 B.n44 163.367
R1361 B.n1388 B.n46 163.367
R1362 B.n1384 B.n46 163.367
R1363 B.n1384 B.n51 163.367
R1364 B.n1380 B.n51 163.367
R1365 B.n1380 B.n53 163.367
R1366 B.n1376 B.n53 163.367
R1367 B.n1376 B.n58 163.367
R1368 B.n1372 B.n58 163.367
R1369 B.n1372 B.n60 163.367
R1370 B.n1368 B.n60 163.367
R1371 B.n1368 B.n65 163.367
R1372 B.n1364 B.n65 163.367
R1373 B.n1364 B.n67 163.367
R1374 B.n1360 B.n67 163.367
R1375 B.n1360 B.n72 163.367
R1376 B.n1356 B.n72 163.367
R1377 B.n1356 B.n74 163.367
R1378 B.n1352 B.n74 163.367
R1379 B.n1352 B.n79 163.367
R1380 B.n1348 B.n79 163.367
R1381 B.n1348 B.n81 163.367
R1382 B.n1344 B.n81 163.367
R1383 B.n1344 B.n86 163.367
R1384 B.n1340 B.n86 163.367
R1385 B.n1340 B.n88 163.367
R1386 B.n1336 B.n88 163.367
R1387 B.n1336 B.n93 163.367
R1388 B.n1332 B.n93 163.367
R1389 B.n1332 B.n95 163.367
R1390 B.n1328 B.n95 163.367
R1391 B.n1328 B.n100 163.367
R1392 B.n1324 B.n100 163.367
R1393 B.n1324 B.n102 163.367
R1394 B.n1320 B.n102 163.367
R1395 B.n1320 B.n107 163.367
R1396 B.n1316 B.n107 163.367
R1397 B.n1316 B.n109 163.367
R1398 B.n1312 B.n109 163.367
R1399 B.n1312 B.n114 163.367
R1400 B.n1308 B.n114 163.367
R1401 B.n1308 B.n116 163.367
R1402 B.n1304 B.n116 163.367
R1403 B.n1304 B.n120 163.367
R1404 B.n1300 B.n120 163.367
R1405 B.n1300 B.n122 163.367
R1406 B.n1296 B.n122 163.367
R1407 B.n1296 B.n128 163.367
R1408 B.n1292 B.n128 163.367
R1409 B.n1292 B.n130 163.367
R1410 B.n1288 B.n130 163.367
R1411 B.n1288 B.n135 163.367
R1412 B.n1284 B.n135 163.367
R1413 B.n691 B.n689 163.367
R1414 B.n695 B.n689 163.367
R1415 B.n699 B.n697 163.367
R1416 B.n703 B.n687 163.367
R1417 B.n707 B.n705 163.367
R1418 B.n711 B.n685 163.367
R1419 B.n715 B.n713 163.367
R1420 B.n719 B.n683 163.367
R1421 B.n723 B.n721 163.367
R1422 B.n727 B.n681 163.367
R1423 B.n731 B.n729 163.367
R1424 B.n735 B.n679 163.367
R1425 B.n739 B.n737 163.367
R1426 B.n743 B.n677 163.367
R1427 B.n747 B.n745 163.367
R1428 B.n751 B.n675 163.367
R1429 B.n755 B.n753 163.367
R1430 B.n759 B.n673 163.367
R1431 B.n763 B.n761 163.367
R1432 B.n767 B.n671 163.367
R1433 B.n771 B.n769 163.367
R1434 B.n775 B.n669 163.367
R1435 B.n779 B.n777 163.367
R1436 B.n783 B.n667 163.367
R1437 B.n787 B.n785 163.367
R1438 B.n791 B.n665 163.367
R1439 B.n795 B.n793 163.367
R1440 B.n799 B.n663 163.367
R1441 B.n803 B.n801 163.367
R1442 B.n807 B.n661 163.367
R1443 B.n811 B.n809 163.367
R1444 B.n815 B.n656 163.367
R1445 B.n819 B.n817 163.367
R1446 B.n823 B.n654 163.367
R1447 B.n827 B.n825 163.367
R1448 B.n832 B.n650 163.367
R1449 B.n836 B.n834 163.367
R1450 B.n840 B.n648 163.367
R1451 B.n844 B.n842 163.367
R1452 B.n848 B.n646 163.367
R1453 B.n852 B.n850 163.367
R1454 B.n856 B.n644 163.367
R1455 B.n860 B.n858 163.367
R1456 B.n864 B.n642 163.367
R1457 B.n868 B.n866 163.367
R1458 B.n872 B.n640 163.367
R1459 B.n876 B.n874 163.367
R1460 B.n880 B.n638 163.367
R1461 B.n884 B.n882 163.367
R1462 B.n888 B.n636 163.367
R1463 B.n892 B.n890 163.367
R1464 B.n896 B.n634 163.367
R1465 B.n900 B.n898 163.367
R1466 B.n904 B.n632 163.367
R1467 B.n908 B.n906 163.367
R1468 B.n912 B.n630 163.367
R1469 B.n916 B.n914 163.367
R1470 B.n920 B.n628 163.367
R1471 B.n924 B.n922 163.367
R1472 B.n928 B.n626 163.367
R1473 B.n932 B.n930 163.367
R1474 B.n936 B.n624 163.367
R1475 B.n940 B.n938 163.367
R1476 B.n944 B.n622 163.367
R1477 B.n947 B.n946 163.367
R1478 B.n949 B.n619 163.367
R1479 B.n953 B.n613 163.367
R1480 B.n961 B.n613 163.367
R1481 B.n961 B.n611 163.367
R1482 B.n965 B.n611 163.367
R1483 B.n965 B.n605 163.367
R1484 B.n973 B.n605 163.367
R1485 B.n973 B.n603 163.367
R1486 B.n977 B.n603 163.367
R1487 B.n977 B.n598 163.367
R1488 B.n986 B.n598 163.367
R1489 B.n986 B.n596 163.367
R1490 B.n990 B.n596 163.367
R1491 B.n990 B.n590 163.367
R1492 B.n998 B.n590 163.367
R1493 B.n998 B.n588 163.367
R1494 B.n1002 B.n588 163.367
R1495 B.n1002 B.n582 163.367
R1496 B.n1010 B.n582 163.367
R1497 B.n1010 B.n580 163.367
R1498 B.n1014 B.n580 163.367
R1499 B.n1014 B.n573 163.367
R1500 B.n1022 B.n573 163.367
R1501 B.n1022 B.n571 163.367
R1502 B.n1026 B.n571 163.367
R1503 B.n1026 B.n566 163.367
R1504 B.n1034 B.n566 163.367
R1505 B.n1034 B.n564 163.367
R1506 B.n1038 B.n564 163.367
R1507 B.n1038 B.n558 163.367
R1508 B.n1046 B.n558 163.367
R1509 B.n1046 B.n556 163.367
R1510 B.n1050 B.n556 163.367
R1511 B.n1050 B.n550 163.367
R1512 B.n1058 B.n550 163.367
R1513 B.n1058 B.n548 163.367
R1514 B.n1062 B.n548 163.367
R1515 B.n1062 B.n542 163.367
R1516 B.n1070 B.n542 163.367
R1517 B.n1070 B.n540 163.367
R1518 B.n1074 B.n540 163.367
R1519 B.n1074 B.n534 163.367
R1520 B.n1082 B.n534 163.367
R1521 B.n1082 B.n532 163.367
R1522 B.n1086 B.n532 163.367
R1523 B.n1086 B.n526 163.367
R1524 B.n1094 B.n526 163.367
R1525 B.n1094 B.n524 163.367
R1526 B.n1098 B.n524 163.367
R1527 B.n1098 B.n518 163.367
R1528 B.n1106 B.n518 163.367
R1529 B.n1106 B.n516 163.367
R1530 B.n1110 B.n516 163.367
R1531 B.n1110 B.n510 163.367
R1532 B.n1118 B.n510 163.367
R1533 B.n1118 B.n508 163.367
R1534 B.n1122 B.n508 163.367
R1535 B.n1122 B.n503 163.367
R1536 B.n1131 B.n503 163.367
R1537 B.n1131 B.n501 163.367
R1538 B.n1135 B.n501 163.367
R1539 B.n1135 B.n495 163.367
R1540 B.n1143 B.n495 163.367
R1541 B.n1143 B.n493 163.367
R1542 B.n1147 B.n493 163.367
R1543 B.n1147 B.n487 163.367
R1544 B.n1155 B.n487 163.367
R1545 B.n1155 B.n485 163.367
R1546 B.n1159 B.n485 163.367
R1547 B.n1159 B.n479 163.367
R1548 B.n1167 B.n479 163.367
R1549 B.n1167 B.n477 163.367
R1550 B.n1172 B.n477 163.367
R1551 B.n1172 B.n471 163.367
R1552 B.n1180 B.n471 163.367
R1553 B.n1181 B.n1180 163.367
R1554 B.n1181 B.n5 163.367
R1555 B.n6 B.n5 163.367
R1556 B.n7 B.n6 163.367
R1557 B.n1186 B.n7 163.367
R1558 B.n1186 B.n12 163.367
R1559 B.n13 B.n12 163.367
R1560 B.n14 B.n13 163.367
R1561 B.n1191 B.n14 163.367
R1562 B.n1191 B.n19 163.367
R1563 B.n20 B.n19 163.367
R1564 B.n21 B.n20 163.367
R1565 B.n1196 B.n21 163.367
R1566 B.n1196 B.n26 163.367
R1567 B.n27 B.n26 163.367
R1568 B.n28 B.n27 163.367
R1569 B.n1201 B.n28 163.367
R1570 B.n1201 B.n33 163.367
R1571 B.n34 B.n33 163.367
R1572 B.n35 B.n34 163.367
R1573 B.n1206 B.n35 163.367
R1574 B.n1206 B.n40 163.367
R1575 B.n41 B.n40 163.367
R1576 B.n42 B.n41 163.367
R1577 B.n1211 B.n42 163.367
R1578 B.n1211 B.n47 163.367
R1579 B.n48 B.n47 163.367
R1580 B.n49 B.n48 163.367
R1581 B.n1216 B.n49 163.367
R1582 B.n1216 B.n54 163.367
R1583 B.n55 B.n54 163.367
R1584 B.n56 B.n55 163.367
R1585 B.n1221 B.n56 163.367
R1586 B.n1221 B.n61 163.367
R1587 B.n62 B.n61 163.367
R1588 B.n63 B.n62 163.367
R1589 B.n1226 B.n63 163.367
R1590 B.n1226 B.n68 163.367
R1591 B.n69 B.n68 163.367
R1592 B.n70 B.n69 163.367
R1593 B.n1231 B.n70 163.367
R1594 B.n1231 B.n75 163.367
R1595 B.n76 B.n75 163.367
R1596 B.n77 B.n76 163.367
R1597 B.n1236 B.n77 163.367
R1598 B.n1236 B.n82 163.367
R1599 B.n83 B.n82 163.367
R1600 B.n84 B.n83 163.367
R1601 B.n1241 B.n84 163.367
R1602 B.n1241 B.n89 163.367
R1603 B.n90 B.n89 163.367
R1604 B.n91 B.n90 163.367
R1605 B.n1246 B.n91 163.367
R1606 B.n1246 B.n96 163.367
R1607 B.n97 B.n96 163.367
R1608 B.n98 B.n97 163.367
R1609 B.n1251 B.n98 163.367
R1610 B.n1251 B.n103 163.367
R1611 B.n104 B.n103 163.367
R1612 B.n105 B.n104 163.367
R1613 B.n1256 B.n105 163.367
R1614 B.n1256 B.n110 163.367
R1615 B.n111 B.n110 163.367
R1616 B.n112 B.n111 163.367
R1617 B.n1261 B.n112 163.367
R1618 B.n1261 B.n117 163.367
R1619 B.n118 B.n117 163.367
R1620 B.n119 B.n118 163.367
R1621 B.n1266 B.n119 163.367
R1622 B.n1266 B.n124 163.367
R1623 B.n125 B.n124 163.367
R1624 B.n126 B.n125 163.367
R1625 B.n1271 B.n126 163.367
R1626 B.n1271 B.n131 163.367
R1627 B.n132 B.n131 163.367
R1628 B.n133 B.n132 163.367
R1629 B.n1276 B.n133 163.367
R1630 B.n1276 B.n138 163.367
R1631 B.n211 B.n210 163.367
R1632 B.n215 B.n214 163.367
R1633 B.n219 B.n218 163.367
R1634 B.n223 B.n222 163.367
R1635 B.n227 B.n226 163.367
R1636 B.n231 B.n230 163.367
R1637 B.n235 B.n234 163.367
R1638 B.n239 B.n238 163.367
R1639 B.n243 B.n242 163.367
R1640 B.n247 B.n246 163.367
R1641 B.n251 B.n250 163.367
R1642 B.n255 B.n254 163.367
R1643 B.n259 B.n258 163.367
R1644 B.n263 B.n262 163.367
R1645 B.n267 B.n266 163.367
R1646 B.n271 B.n270 163.367
R1647 B.n275 B.n274 163.367
R1648 B.n279 B.n278 163.367
R1649 B.n283 B.n282 163.367
R1650 B.n287 B.n286 163.367
R1651 B.n291 B.n290 163.367
R1652 B.n295 B.n294 163.367
R1653 B.n299 B.n298 163.367
R1654 B.n303 B.n302 163.367
R1655 B.n307 B.n306 163.367
R1656 B.n311 B.n310 163.367
R1657 B.n315 B.n314 163.367
R1658 B.n319 B.n318 163.367
R1659 B.n323 B.n322 163.367
R1660 B.n327 B.n326 163.367
R1661 B.n332 B.n331 163.367
R1662 B.n336 B.n335 163.367
R1663 B.n340 B.n339 163.367
R1664 B.n344 B.n343 163.367
R1665 B.n348 B.n347 163.367
R1666 B.n353 B.n352 163.367
R1667 B.n357 B.n356 163.367
R1668 B.n361 B.n360 163.367
R1669 B.n365 B.n364 163.367
R1670 B.n369 B.n368 163.367
R1671 B.n373 B.n372 163.367
R1672 B.n377 B.n376 163.367
R1673 B.n381 B.n380 163.367
R1674 B.n385 B.n384 163.367
R1675 B.n389 B.n388 163.367
R1676 B.n393 B.n392 163.367
R1677 B.n397 B.n396 163.367
R1678 B.n401 B.n400 163.367
R1679 B.n405 B.n404 163.367
R1680 B.n409 B.n408 163.367
R1681 B.n413 B.n412 163.367
R1682 B.n417 B.n416 163.367
R1683 B.n421 B.n420 163.367
R1684 B.n425 B.n424 163.367
R1685 B.n429 B.n428 163.367
R1686 B.n433 B.n432 163.367
R1687 B.n437 B.n436 163.367
R1688 B.n441 B.n440 163.367
R1689 B.n445 B.n444 163.367
R1690 B.n449 B.n448 163.367
R1691 B.n453 B.n452 163.367
R1692 B.n457 B.n456 163.367
R1693 B.n461 B.n460 163.367
R1694 B.n465 B.n464 163.367
R1695 B.n467 B.n204 163.367
R1696 B.n651 B.t17 146.922
R1697 B.n205 B.t12 146.922
R1698 B.n657 B.t20 146.897
R1699 B.n207 B.t22 146.897
R1700 B.n652 B.n651 74.4732
R1701 B.n658 B.n657 74.4732
R1702 B.n208 B.n207 74.4732
R1703 B.n206 B.n205 74.4732
R1704 B.n652 B.t16 72.4485
R1705 B.n206 B.t13 72.4485
R1706 B.n658 B.t19 72.4238
R1707 B.n208 B.t23 72.4238
R1708 B.n690 B.n617 71.676
R1709 B.n696 B.n695 71.676
R1710 B.n699 B.n698 71.676
R1711 B.n704 B.n703 71.676
R1712 B.n707 B.n706 71.676
R1713 B.n712 B.n711 71.676
R1714 B.n715 B.n714 71.676
R1715 B.n720 B.n719 71.676
R1716 B.n723 B.n722 71.676
R1717 B.n728 B.n727 71.676
R1718 B.n731 B.n730 71.676
R1719 B.n736 B.n735 71.676
R1720 B.n739 B.n738 71.676
R1721 B.n744 B.n743 71.676
R1722 B.n747 B.n746 71.676
R1723 B.n752 B.n751 71.676
R1724 B.n755 B.n754 71.676
R1725 B.n760 B.n759 71.676
R1726 B.n763 B.n762 71.676
R1727 B.n768 B.n767 71.676
R1728 B.n771 B.n770 71.676
R1729 B.n776 B.n775 71.676
R1730 B.n779 B.n778 71.676
R1731 B.n784 B.n783 71.676
R1732 B.n787 B.n786 71.676
R1733 B.n792 B.n791 71.676
R1734 B.n795 B.n794 71.676
R1735 B.n800 B.n799 71.676
R1736 B.n803 B.n802 71.676
R1737 B.n808 B.n807 71.676
R1738 B.n811 B.n810 71.676
R1739 B.n816 B.n815 71.676
R1740 B.n819 B.n818 71.676
R1741 B.n824 B.n823 71.676
R1742 B.n827 B.n826 71.676
R1743 B.n833 B.n832 71.676
R1744 B.n836 B.n835 71.676
R1745 B.n841 B.n840 71.676
R1746 B.n844 B.n843 71.676
R1747 B.n849 B.n848 71.676
R1748 B.n852 B.n851 71.676
R1749 B.n857 B.n856 71.676
R1750 B.n860 B.n859 71.676
R1751 B.n865 B.n864 71.676
R1752 B.n868 B.n867 71.676
R1753 B.n873 B.n872 71.676
R1754 B.n876 B.n875 71.676
R1755 B.n881 B.n880 71.676
R1756 B.n884 B.n883 71.676
R1757 B.n889 B.n888 71.676
R1758 B.n892 B.n891 71.676
R1759 B.n897 B.n896 71.676
R1760 B.n900 B.n899 71.676
R1761 B.n905 B.n904 71.676
R1762 B.n908 B.n907 71.676
R1763 B.n913 B.n912 71.676
R1764 B.n916 B.n915 71.676
R1765 B.n921 B.n920 71.676
R1766 B.n924 B.n923 71.676
R1767 B.n929 B.n928 71.676
R1768 B.n932 B.n931 71.676
R1769 B.n937 B.n936 71.676
R1770 B.n940 B.n939 71.676
R1771 B.n945 B.n944 71.676
R1772 B.n948 B.n947 71.676
R1773 B.n139 B.n137 71.676
R1774 B.n211 B.n140 71.676
R1775 B.n215 B.n141 71.676
R1776 B.n219 B.n142 71.676
R1777 B.n223 B.n143 71.676
R1778 B.n227 B.n144 71.676
R1779 B.n231 B.n145 71.676
R1780 B.n235 B.n146 71.676
R1781 B.n239 B.n147 71.676
R1782 B.n243 B.n148 71.676
R1783 B.n247 B.n149 71.676
R1784 B.n251 B.n150 71.676
R1785 B.n255 B.n151 71.676
R1786 B.n259 B.n152 71.676
R1787 B.n263 B.n153 71.676
R1788 B.n267 B.n154 71.676
R1789 B.n271 B.n155 71.676
R1790 B.n275 B.n156 71.676
R1791 B.n279 B.n157 71.676
R1792 B.n283 B.n158 71.676
R1793 B.n287 B.n159 71.676
R1794 B.n291 B.n160 71.676
R1795 B.n295 B.n161 71.676
R1796 B.n299 B.n162 71.676
R1797 B.n303 B.n163 71.676
R1798 B.n307 B.n164 71.676
R1799 B.n311 B.n165 71.676
R1800 B.n315 B.n166 71.676
R1801 B.n319 B.n167 71.676
R1802 B.n323 B.n168 71.676
R1803 B.n327 B.n169 71.676
R1804 B.n332 B.n170 71.676
R1805 B.n336 B.n171 71.676
R1806 B.n340 B.n172 71.676
R1807 B.n344 B.n173 71.676
R1808 B.n348 B.n174 71.676
R1809 B.n353 B.n175 71.676
R1810 B.n357 B.n176 71.676
R1811 B.n361 B.n177 71.676
R1812 B.n365 B.n178 71.676
R1813 B.n369 B.n179 71.676
R1814 B.n373 B.n180 71.676
R1815 B.n377 B.n181 71.676
R1816 B.n381 B.n182 71.676
R1817 B.n385 B.n183 71.676
R1818 B.n389 B.n184 71.676
R1819 B.n393 B.n185 71.676
R1820 B.n397 B.n186 71.676
R1821 B.n401 B.n187 71.676
R1822 B.n405 B.n188 71.676
R1823 B.n409 B.n189 71.676
R1824 B.n413 B.n190 71.676
R1825 B.n417 B.n191 71.676
R1826 B.n421 B.n192 71.676
R1827 B.n425 B.n193 71.676
R1828 B.n429 B.n194 71.676
R1829 B.n433 B.n195 71.676
R1830 B.n437 B.n196 71.676
R1831 B.n441 B.n197 71.676
R1832 B.n445 B.n198 71.676
R1833 B.n449 B.n199 71.676
R1834 B.n453 B.n200 71.676
R1835 B.n457 B.n201 71.676
R1836 B.n461 B.n202 71.676
R1837 B.n465 B.n203 71.676
R1838 B.n1281 B.n204 71.676
R1839 B.n1281 B.n1280 71.676
R1840 B.n467 B.n203 71.676
R1841 B.n464 B.n202 71.676
R1842 B.n460 B.n201 71.676
R1843 B.n456 B.n200 71.676
R1844 B.n452 B.n199 71.676
R1845 B.n448 B.n198 71.676
R1846 B.n444 B.n197 71.676
R1847 B.n440 B.n196 71.676
R1848 B.n436 B.n195 71.676
R1849 B.n432 B.n194 71.676
R1850 B.n428 B.n193 71.676
R1851 B.n424 B.n192 71.676
R1852 B.n420 B.n191 71.676
R1853 B.n416 B.n190 71.676
R1854 B.n412 B.n189 71.676
R1855 B.n408 B.n188 71.676
R1856 B.n404 B.n187 71.676
R1857 B.n400 B.n186 71.676
R1858 B.n396 B.n185 71.676
R1859 B.n392 B.n184 71.676
R1860 B.n388 B.n183 71.676
R1861 B.n384 B.n182 71.676
R1862 B.n380 B.n181 71.676
R1863 B.n376 B.n180 71.676
R1864 B.n372 B.n179 71.676
R1865 B.n368 B.n178 71.676
R1866 B.n364 B.n177 71.676
R1867 B.n360 B.n176 71.676
R1868 B.n356 B.n175 71.676
R1869 B.n352 B.n174 71.676
R1870 B.n347 B.n173 71.676
R1871 B.n343 B.n172 71.676
R1872 B.n339 B.n171 71.676
R1873 B.n335 B.n170 71.676
R1874 B.n331 B.n169 71.676
R1875 B.n326 B.n168 71.676
R1876 B.n322 B.n167 71.676
R1877 B.n318 B.n166 71.676
R1878 B.n314 B.n165 71.676
R1879 B.n310 B.n164 71.676
R1880 B.n306 B.n163 71.676
R1881 B.n302 B.n162 71.676
R1882 B.n298 B.n161 71.676
R1883 B.n294 B.n160 71.676
R1884 B.n290 B.n159 71.676
R1885 B.n286 B.n158 71.676
R1886 B.n282 B.n157 71.676
R1887 B.n278 B.n156 71.676
R1888 B.n274 B.n155 71.676
R1889 B.n270 B.n154 71.676
R1890 B.n266 B.n153 71.676
R1891 B.n262 B.n152 71.676
R1892 B.n258 B.n151 71.676
R1893 B.n254 B.n150 71.676
R1894 B.n250 B.n149 71.676
R1895 B.n246 B.n148 71.676
R1896 B.n242 B.n147 71.676
R1897 B.n238 B.n146 71.676
R1898 B.n234 B.n145 71.676
R1899 B.n230 B.n144 71.676
R1900 B.n226 B.n143 71.676
R1901 B.n222 B.n142 71.676
R1902 B.n218 B.n141 71.676
R1903 B.n214 B.n140 71.676
R1904 B.n210 B.n139 71.676
R1905 B.n691 B.n690 71.676
R1906 B.n697 B.n696 71.676
R1907 B.n698 B.n687 71.676
R1908 B.n705 B.n704 71.676
R1909 B.n706 B.n685 71.676
R1910 B.n713 B.n712 71.676
R1911 B.n714 B.n683 71.676
R1912 B.n721 B.n720 71.676
R1913 B.n722 B.n681 71.676
R1914 B.n729 B.n728 71.676
R1915 B.n730 B.n679 71.676
R1916 B.n737 B.n736 71.676
R1917 B.n738 B.n677 71.676
R1918 B.n745 B.n744 71.676
R1919 B.n746 B.n675 71.676
R1920 B.n753 B.n752 71.676
R1921 B.n754 B.n673 71.676
R1922 B.n761 B.n760 71.676
R1923 B.n762 B.n671 71.676
R1924 B.n769 B.n768 71.676
R1925 B.n770 B.n669 71.676
R1926 B.n777 B.n776 71.676
R1927 B.n778 B.n667 71.676
R1928 B.n785 B.n784 71.676
R1929 B.n786 B.n665 71.676
R1930 B.n793 B.n792 71.676
R1931 B.n794 B.n663 71.676
R1932 B.n801 B.n800 71.676
R1933 B.n802 B.n661 71.676
R1934 B.n809 B.n808 71.676
R1935 B.n810 B.n656 71.676
R1936 B.n817 B.n816 71.676
R1937 B.n818 B.n654 71.676
R1938 B.n825 B.n824 71.676
R1939 B.n826 B.n650 71.676
R1940 B.n834 B.n833 71.676
R1941 B.n835 B.n648 71.676
R1942 B.n842 B.n841 71.676
R1943 B.n843 B.n646 71.676
R1944 B.n850 B.n849 71.676
R1945 B.n851 B.n644 71.676
R1946 B.n858 B.n857 71.676
R1947 B.n859 B.n642 71.676
R1948 B.n866 B.n865 71.676
R1949 B.n867 B.n640 71.676
R1950 B.n874 B.n873 71.676
R1951 B.n875 B.n638 71.676
R1952 B.n882 B.n881 71.676
R1953 B.n883 B.n636 71.676
R1954 B.n890 B.n889 71.676
R1955 B.n891 B.n634 71.676
R1956 B.n898 B.n897 71.676
R1957 B.n899 B.n632 71.676
R1958 B.n906 B.n905 71.676
R1959 B.n907 B.n630 71.676
R1960 B.n914 B.n913 71.676
R1961 B.n915 B.n628 71.676
R1962 B.n922 B.n921 71.676
R1963 B.n923 B.n626 71.676
R1964 B.n930 B.n929 71.676
R1965 B.n931 B.n624 71.676
R1966 B.n938 B.n937 71.676
R1967 B.n939 B.n622 71.676
R1968 B.n946 B.n945 71.676
R1969 B.n949 B.n948 71.676
R1970 B.n830 B.n652 59.5399
R1971 B.n659 B.n658 59.5399
R1972 B.n329 B.n208 59.5399
R1973 B.n350 B.n206 59.5399
R1974 B.n954 B.n618 52.9183
R1975 B.n1283 B.n1282 52.9183
R1976 B.n954 B.n614 31.291
R1977 B.n960 B.n614 31.291
R1978 B.n960 B.n610 31.291
R1979 B.n966 B.n610 31.291
R1980 B.n966 B.n606 31.291
R1981 B.n972 B.n606 31.291
R1982 B.n972 B.n602 31.291
R1983 B.n979 B.n602 31.291
R1984 B.n979 B.n978 31.291
R1985 B.n985 B.n595 31.291
R1986 B.n991 B.n595 31.291
R1987 B.n991 B.n591 31.291
R1988 B.n997 B.n591 31.291
R1989 B.n997 B.n587 31.291
R1990 B.n1003 B.n587 31.291
R1991 B.n1003 B.n583 31.291
R1992 B.n1009 B.n583 31.291
R1993 B.n1009 B.n579 31.291
R1994 B.n1015 B.n579 31.291
R1995 B.n1015 B.n574 31.291
R1996 B.n1021 B.n574 31.291
R1997 B.n1021 B.n575 31.291
R1998 B.n1027 B.n567 31.291
R1999 B.n1033 B.n567 31.291
R2000 B.n1033 B.n563 31.291
R2001 B.n1039 B.n563 31.291
R2002 B.n1039 B.n559 31.291
R2003 B.n1045 B.n559 31.291
R2004 B.n1045 B.n555 31.291
R2005 B.n1051 B.n555 31.291
R2006 B.n1051 B.n551 31.291
R2007 B.n1057 B.n551 31.291
R2008 B.n1063 B.n547 31.291
R2009 B.n1063 B.n543 31.291
R2010 B.n1069 B.n543 31.291
R2011 B.n1069 B.n539 31.291
R2012 B.n1075 B.n539 31.291
R2013 B.n1075 B.n535 31.291
R2014 B.n1081 B.n535 31.291
R2015 B.n1081 B.n531 31.291
R2016 B.n1087 B.n531 31.291
R2017 B.n1087 B.n527 31.291
R2018 B.n1093 B.n527 31.291
R2019 B.n1099 B.n523 31.291
R2020 B.n1099 B.n519 31.291
R2021 B.n1105 B.n519 31.291
R2022 B.n1105 B.n515 31.291
R2023 B.n1111 B.n515 31.291
R2024 B.n1111 B.n511 31.291
R2025 B.n1117 B.n511 31.291
R2026 B.n1117 B.n507 31.291
R2027 B.n1124 B.n507 31.291
R2028 B.n1124 B.n1123 31.291
R2029 B.n1130 B.n500 31.291
R2030 B.n1136 B.n500 31.291
R2031 B.n1136 B.n496 31.291
R2032 B.n1142 B.n496 31.291
R2033 B.n1142 B.n492 31.291
R2034 B.n1148 B.n492 31.291
R2035 B.n1148 B.n488 31.291
R2036 B.n1154 B.n488 31.291
R2037 B.n1154 B.n484 31.291
R2038 B.n1160 B.n484 31.291
R2039 B.n1166 B.n480 31.291
R2040 B.n1166 B.n476 31.291
R2041 B.n1173 B.n476 31.291
R2042 B.n1173 B.n472 31.291
R2043 B.n1179 B.n472 31.291
R2044 B.n1179 B.n4 31.291
R2045 B.n1435 B.n4 31.291
R2046 B.n1435 B.n1434 31.291
R2047 B.n1434 B.n1433 31.291
R2048 B.n1433 B.n8 31.291
R2049 B.n1427 B.n8 31.291
R2050 B.n1427 B.n1426 31.291
R2051 B.n1426 B.n1425 31.291
R2052 B.n1425 B.n15 31.291
R2053 B.n1419 B.n1418 31.291
R2054 B.n1418 B.n1417 31.291
R2055 B.n1417 B.n22 31.291
R2056 B.n1411 B.n22 31.291
R2057 B.n1411 B.n1410 31.291
R2058 B.n1410 B.n1409 31.291
R2059 B.n1409 B.n29 31.291
R2060 B.n1403 B.n29 31.291
R2061 B.n1403 B.n1402 31.291
R2062 B.n1402 B.n1401 31.291
R2063 B.n1395 B.n39 31.291
R2064 B.n1395 B.n1394 31.291
R2065 B.n1394 B.n1393 31.291
R2066 B.n1393 B.n43 31.291
R2067 B.n1387 B.n43 31.291
R2068 B.n1387 B.n1386 31.291
R2069 B.n1386 B.n1385 31.291
R2070 B.n1385 B.n50 31.291
R2071 B.n1379 B.n50 31.291
R2072 B.n1379 B.n1378 31.291
R2073 B.n1377 B.n57 31.291
R2074 B.n1371 B.n57 31.291
R2075 B.n1371 B.n1370 31.291
R2076 B.n1370 B.n1369 31.291
R2077 B.n1369 B.n64 31.291
R2078 B.n1363 B.n64 31.291
R2079 B.n1363 B.n1362 31.291
R2080 B.n1362 B.n1361 31.291
R2081 B.n1361 B.n71 31.291
R2082 B.n1355 B.n71 31.291
R2083 B.n1355 B.n1354 31.291
R2084 B.n1353 B.n78 31.291
R2085 B.n1347 B.n78 31.291
R2086 B.n1347 B.n1346 31.291
R2087 B.n1346 B.n1345 31.291
R2088 B.n1345 B.n85 31.291
R2089 B.n1339 B.n85 31.291
R2090 B.n1339 B.n1338 31.291
R2091 B.n1338 B.n1337 31.291
R2092 B.n1337 B.n92 31.291
R2093 B.n1331 B.n92 31.291
R2094 B.n1330 B.n1329 31.291
R2095 B.n1329 B.n99 31.291
R2096 B.n1323 B.n99 31.291
R2097 B.n1323 B.n1322 31.291
R2098 B.n1322 B.n1321 31.291
R2099 B.n1321 B.n106 31.291
R2100 B.n1315 B.n106 31.291
R2101 B.n1315 B.n1314 31.291
R2102 B.n1314 B.n1313 31.291
R2103 B.n1313 B.n113 31.291
R2104 B.n1307 B.n113 31.291
R2105 B.n1307 B.n1306 31.291
R2106 B.n1306 B.n1305 31.291
R2107 B.n1299 B.n123 31.291
R2108 B.n1299 B.n1298 31.291
R2109 B.n1298 B.n1297 31.291
R2110 B.n1297 B.n127 31.291
R2111 B.n1291 B.n127 31.291
R2112 B.n1291 B.n1290 31.291
R2113 B.n1290 B.n1289 31.291
R2114 B.n1289 B.n134 31.291
R2115 B.n1283 B.n134 31.291
R2116 B.n1285 B.n136 30.1273
R2117 B.n1279 B.n1278 30.1273
R2118 B.n952 B.n951 30.1273
R2119 B.n956 B.n616 30.1273
R2120 B.n985 B.t15 28.9903
R2121 B.n1305 B.t11 28.9903
R2122 B.n1057 B.t7 27.1496
R2123 B.t0 B.n1353 27.1496
R2124 B.t4 B.n523 26.2293
R2125 B.n1378 B.t6 26.2293
R2126 B.n1160 B.t2 23.4684
R2127 B.n1419 B.t5 23.4684
R2128 B B.n1437 18.0485
R2129 B.n575 B.t9 17.9465
R2130 B.t3 B.n1330 17.9465
R2131 B.n1130 B.t1 17.0262
R2132 B.n1401 B.t8 17.0262
R2133 B.n1123 B.t1 14.2653
R2134 B.n39 B.t8 14.2653
R2135 B.n1027 B.t9 13.345
R2136 B.n1331 B.t3 13.345
R2137 B.n209 B.n136 10.6151
R2138 B.n212 B.n209 10.6151
R2139 B.n213 B.n212 10.6151
R2140 B.n216 B.n213 10.6151
R2141 B.n217 B.n216 10.6151
R2142 B.n220 B.n217 10.6151
R2143 B.n221 B.n220 10.6151
R2144 B.n224 B.n221 10.6151
R2145 B.n225 B.n224 10.6151
R2146 B.n228 B.n225 10.6151
R2147 B.n229 B.n228 10.6151
R2148 B.n232 B.n229 10.6151
R2149 B.n233 B.n232 10.6151
R2150 B.n236 B.n233 10.6151
R2151 B.n237 B.n236 10.6151
R2152 B.n240 B.n237 10.6151
R2153 B.n241 B.n240 10.6151
R2154 B.n244 B.n241 10.6151
R2155 B.n245 B.n244 10.6151
R2156 B.n248 B.n245 10.6151
R2157 B.n249 B.n248 10.6151
R2158 B.n252 B.n249 10.6151
R2159 B.n253 B.n252 10.6151
R2160 B.n256 B.n253 10.6151
R2161 B.n257 B.n256 10.6151
R2162 B.n260 B.n257 10.6151
R2163 B.n261 B.n260 10.6151
R2164 B.n264 B.n261 10.6151
R2165 B.n265 B.n264 10.6151
R2166 B.n268 B.n265 10.6151
R2167 B.n269 B.n268 10.6151
R2168 B.n272 B.n269 10.6151
R2169 B.n273 B.n272 10.6151
R2170 B.n276 B.n273 10.6151
R2171 B.n277 B.n276 10.6151
R2172 B.n280 B.n277 10.6151
R2173 B.n281 B.n280 10.6151
R2174 B.n284 B.n281 10.6151
R2175 B.n285 B.n284 10.6151
R2176 B.n288 B.n285 10.6151
R2177 B.n289 B.n288 10.6151
R2178 B.n292 B.n289 10.6151
R2179 B.n293 B.n292 10.6151
R2180 B.n296 B.n293 10.6151
R2181 B.n297 B.n296 10.6151
R2182 B.n300 B.n297 10.6151
R2183 B.n301 B.n300 10.6151
R2184 B.n304 B.n301 10.6151
R2185 B.n305 B.n304 10.6151
R2186 B.n308 B.n305 10.6151
R2187 B.n309 B.n308 10.6151
R2188 B.n312 B.n309 10.6151
R2189 B.n313 B.n312 10.6151
R2190 B.n316 B.n313 10.6151
R2191 B.n317 B.n316 10.6151
R2192 B.n320 B.n317 10.6151
R2193 B.n321 B.n320 10.6151
R2194 B.n324 B.n321 10.6151
R2195 B.n325 B.n324 10.6151
R2196 B.n328 B.n325 10.6151
R2197 B.n333 B.n330 10.6151
R2198 B.n334 B.n333 10.6151
R2199 B.n337 B.n334 10.6151
R2200 B.n338 B.n337 10.6151
R2201 B.n341 B.n338 10.6151
R2202 B.n342 B.n341 10.6151
R2203 B.n345 B.n342 10.6151
R2204 B.n346 B.n345 10.6151
R2205 B.n349 B.n346 10.6151
R2206 B.n354 B.n351 10.6151
R2207 B.n355 B.n354 10.6151
R2208 B.n358 B.n355 10.6151
R2209 B.n359 B.n358 10.6151
R2210 B.n362 B.n359 10.6151
R2211 B.n363 B.n362 10.6151
R2212 B.n366 B.n363 10.6151
R2213 B.n367 B.n366 10.6151
R2214 B.n370 B.n367 10.6151
R2215 B.n371 B.n370 10.6151
R2216 B.n374 B.n371 10.6151
R2217 B.n375 B.n374 10.6151
R2218 B.n378 B.n375 10.6151
R2219 B.n379 B.n378 10.6151
R2220 B.n382 B.n379 10.6151
R2221 B.n383 B.n382 10.6151
R2222 B.n386 B.n383 10.6151
R2223 B.n387 B.n386 10.6151
R2224 B.n390 B.n387 10.6151
R2225 B.n391 B.n390 10.6151
R2226 B.n394 B.n391 10.6151
R2227 B.n395 B.n394 10.6151
R2228 B.n398 B.n395 10.6151
R2229 B.n399 B.n398 10.6151
R2230 B.n402 B.n399 10.6151
R2231 B.n403 B.n402 10.6151
R2232 B.n406 B.n403 10.6151
R2233 B.n407 B.n406 10.6151
R2234 B.n410 B.n407 10.6151
R2235 B.n411 B.n410 10.6151
R2236 B.n414 B.n411 10.6151
R2237 B.n415 B.n414 10.6151
R2238 B.n418 B.n415 10.6151
R2239 B.n419 B.n418 10.6151
R2240 B.n422 B.n419 10.6151
R2241 B.n423 B.n422 10.6151
R2242 B.n426 B.n423 10.6151
R2243 B.n427 B.n426 10.6151
R2244 B.n430 B.n427 10.6151
R2245 B.n431 B.n430 10.6151
R2246 B.n434 B.n431 10.6151
R2247 B.n435 B.n434 10.6151
R2248 B.n438 B.n435 10.6151
R2249 B.n439 B.n438 10.6151
R2250 B.n442 B.n439 10.6151
R2251 B.n443 B.n442 10.6151
R2252 B.n446 B.n443 10.6151
R2253 B.n447 B.n446 10.6151
R2254 B.n450 B.n447 10.6151
R2255 B.n451 B.n450 10.6151
R2256 B.n454 B.n451 10.6151
R2257 B.n455 B.n454 10.6151
R2258 B.n458 B.n455 10.6151
R2259 B.n459 B.n458 10.6151
R2260 B.n462 B.n459 10.6151
R2261 B.n463 B.n462 10.6151
R2262 B.n466 B.n463 10.6151
R2263 B.n468 B.n466 10.6151
R2264 B.n469 B.n468 10.6151
R2265 B.n1279 B.n469 10.6151
R2266 B.n952 B.n612 10.6151
R2267 B.n962 B.n612 10.6151
R2268 B.n963 B.n962 10.6151
R2269 B.n964 B.n963 10.6151
R2270 B.n964 B.n604 10.6151
R2271 B.n974 B.n604 10.6151
R2272 B.n975 B.n974 10.6151
R2273 B.n976 B.n975 10.6151
R2274 B.n976 B.n597 10.6151
R2275 B.n987 B.n597 10.6151
R2276 B.n988 B.n987 10.6151
R2277 B.n989 B.n988 10.6151
R2278 B.n989 B.n589 10.6151
R2279 B.n999 B.n589 10.6151
R2280 B.n1000 B.n999 10.6151
R2281 B.n1001 B.n1000 10.6151
R2282 B.n1001 B.n581 10.6151
R2283 B.n1011 B.n581 10.6151
R2284 B.n1012 B.n1011 10.6151
R2285 B.n1013 B.n1012 10.6151
R2286 B.n1013 B.n572 10.6151
R2287 B.n1023 B.n572 10.6151
R2288 B.n1024 B.n1023 10.6151
R2289 B.n1025 B.n1024 10.6151
R2290 B.n1025 B.n565 10.6151
R2291 B.n1035 B.n565 10.6151
R2292 B.n1036 B.n1035 10.6151
R2293 B.n1037 B.n1036 10.6151
R2294 B.n1037 B.n557 10.6151
R2295 B.n1047 B.n557 10.6151
R2296 B.n1048 B.n1047 10.6151
R2297 B.n1049 B.n1048 10.6151
R2298 B.n1049 B.n549 10.6151
R2299 B.n1059 B.n549 10.6151
R2300 B.n1060 B.n1059 10.6151
R2301 B.n1061 B.n1060 10.6151
R2302 B.n1061 B.n541 10.6151
R2303 B.n1071 B.n541 10.6151
R2304 B.n1072 B.n1071 10.6151
R2305 B.n1073 B.n1072 10.6151
R2306 B.n1073 B.n533 10.6151
R2307 B.n1083 B.n533 10.6151
R2308 B.n1084 B.n1083 10.6151
R2309 B.n1085 B.n1084 10.6151
R2310 B.n1085 B.n525 10.6151
R2311 B.n1095 B.n525 10.6151
R2312 B.n1096 B.n1095 10.6151
R2313 B.n1097 B.n1096 10.6151
R2314 B.n1097 B.n517 10.6151
R2315 B.n1107 B.n517 10.6151
R2316 B.n1108 B.n1107 10.6151
R2317 B.n1109 B.n1108 10.6151
R2318 B.n1109 B.n509 10.6151
R2319 B.n1119 B.n509 10.6151
R2320 B.n1120 B.n1119 10.6151
R2321 B.n1121 B.n1120 10.6151
R2322 B.n1121 B.n502 10.6151
R2323 B.n1132 B.n502 10.6151
R2324 B.n1133 B.n1132 10.6151
R2325 B.n1134 B.n1133 10.6151
R2326 B.n1134 B.n494 10.6151
R2327 B.n1144 B.n494 10.6151
R2328 B.n1145 B.n1144 10.6151
R2329 B.n1146 B.n1145 10.6151
R2330 B.n1146 B.n486 10.6151
R2331 B.n1156 B.n486 10.6151
R2332 B.n1157 B.n1156 10.6151
R2333 B.n1158 B.n1157 10.6151
R2334 B.n1158 B.n478 10.6151
R2335 B.n1168 B.n478 10.6151
R2336 B.n1169 B.n1168 10.6151
R2337 B.n1171 B.n1169 10.6151
R2338 B.n1171 B.n1170 10.6151
R2339 B.n1170 B.n470 10.6151
R2340 B.n1182 B.n470 10.6151
R2341 B.n1183 B.n1182 10.6151
R2342 B.n1184 B.n1183 10.6151
R2343 B.n1185 B.n1184 10.6151
R2344 B.n1187 B.n1185 10.6151
R2345 B.n1188 B.n1187 10.6151
R2346 B.n1189 B.n1188 10.6151
R2347 B.n1190 B.n1189 10.6151
R2348 B.n1192 B.n1190 10.6151
R2349 B.n1193 B.n1192 10.6151
R2350 B.n1194 B.n1193 10.6151
R2351 B.n1195 B.n1194 10.6151
R2352 B.n1197 B.n1195 10.6151
R2353 B.n1198 B.n1197 10.6151
R2354 B.n1199 B.n1198 10.6151
R2355 B.n1200 B.n1199 10.6151
R2356 B.n1202 B.n1200 10.6151
R2357 B.n1203 B.n1202 10.6151
R2358 B.n1204 B.n1203 10.6151
R2359 B.n1205 B.n1204 10.6151
R2360 B.n1207 B.n1205 10.6151
R2361 B.n1208 B.n1207 10.6151
R2362 B.n1209 B.n1208 10.6151
R2363 B.n1210 B.n1209 10.6151
R2364 B.n1212 B.n1210 10.6151
R2365 B.n1213 B.n1212 10.6151
R2366 B.n1214 B.n1213 10.6151
R2367 B.n1215 B.n1214 10.6151
R2368 B.n1217 B.n1215 10.6151
R2369 B.n1218 B.n1217 10.6151
R2370 B.n1219 B.n1218 10.6151
R2371 B.n1220 B.n1219 10.6151
R2372 B.n1222 B.n1220 10.6151
R2373 B.n1223 B.n1222 10.6151
R2374 B.n1224 B.n1223 10.6151
R2375 B.n1225 B.n1224 10.6151
R2376 B.n1227 B.n1225 10.6151
R2377 B.n1228 B.n1227 10.6151
R2378 B.n1229 B.n1228 10.6151
R2379 B.n1230 B.n1229 10.6151
R2380 B.n1232 B.n1230 10.6151
R2381 B.n1233 B.n1232 10.6151
R2382 B.n1234 B.n1233 10.6151
R2383 B.n1235 B.n1234 10.6151
R2384 B.n1237 B.n1235 10.6151
R2385 B.n1238 B.n1237 10.6151
R2386 B.n1239 B.n1238 10.6151
R2387 B.n1240 B.n1239 10.6151
R2388 B.n1242 B.n1240 10.6151
R2389 B.n1243 B.n1242 10.6151
R2390 B.n1244 B.n1243 10.6151
R2391 B.n1245 B.n1244 10.6151
R2392 B.n1247 B.n1245 10.6151
R2393 B.n1248 B.n1247 10.6151
R2394 B.n1249 B.n1248 10.6151
R2395 B.n1250 B.n1249 10.6151
R2396 B.n1252 B.n1250 10.6151
R2397 B.n1253 B.n1252 10.6151
R2398 B.n1254 B.n1253 10.6151
R2399 B.n1255 B.n1254 10.6151
R2400 B.n1257 B.n1255 10.6151
R2401 B.n1258 B.n1257 10.6151
R2402 B.n1259 B.n1258 10.6151
R2403 B.n1260 B.n1259 10.6151
R2404 B.n1262 B.n1260 10.6151
R2405 B.n1263 B.n1262 10.6151
R2406 B.n1264 B.n1263 10.6151
R2407 B.n1265 B.n1264 10.6151
R2408 B.n1267 B.n1265 10.6151
R2409 B.n1268 B.n1267 10.6151
R2410 B.n1269 B.n1268 10.6151
R2411 B.n1270 B.n1269 10.6151
R2412 B.n1272 B.n1270 10.6151
R2413 B.n1273 B.n1272 10.6151
R2414 B.n1274 B.n1273 10.6151
R2415 B.n1275 B.n1274 10.6151
R2416 B.n1277 B.n1275 10.6151
R2417 B.n1278 B.n1277 10.6151
R2418 B.n692 B.n616 10.6151
R2419 B.n693 B.n692 10.6151
R2420 B.n694 B.n693 10.6151
R2421 B.n694 B.n688 10.6151
R2422 B.n700 B.n688 10.6151
R2423 B.n701 B.n700 10.6151
R2424 B.n702 B.n701 10.6151
R2425 B.n702 B.n686 10.6151
R2426 B.n708 B.n686 10.6151
R2427 B.n709 B.n708 10.6151
R2428 B.n710 B.n709 10.6151
R2429 B.n710 B.n684 10.6151
R2430 B.n716 B.n684 10.6151
R2431 B.n717 B.n716 10.6151
R2432 B.n718 B.n717 10.6151
R2433 B.n718 B.n682 10.6151
R2434 B.n724 B.n682 10.6151
R2435 B.n725 B.n724 10.6151
R2436 B.n726 B.n725 10.6151
R2437 B.n726 B.n680 10.6151
R2438 B.n732 B.n680 10.6151
R2439 B.n733 B.n732 10.6151
R2440 B.n734 B.n733 10.6151
R2441 B.n734 B.n678 10.6151
R2442 B.n740 B.n678 10.6151
R2443 B.n741 B.n740 10.6151
R2444 B.n742 B.n741 10.6151
R2445 B.n742 B.n676 10.6151
R2446 B.n748 B.n676 10.6151
R2447 B.n749 B.n748 10.6151
R2448 B.n750 B.n749 10.6151
R2449 B.n750 B.n674 10.6151
R2450 B.n756 B.n674 10.6151
R2451 B.n757 B.n756 10.6151
R2452 B.n758 B.n757 10.6151
R2453 B.n758 B.n672 10.6151
R2454 B.n764 B.n672 10.6151
R2455 B.n765 B.n764 10.6151
R2456 B.n766 B.n765 10.6151
R2457 B.n766 B.n670 10.6151
R2458 B.n772 B.n670 10.6151
R2459 B.n773 B.n772 10.6151
R2460 B.n774 B.n773 10.6151
R2461 B.n774 B.n668 10.6151
R2462 B.n780 B.n668 10.6151
R2463 B.n781 B.n780 10.6151
R2464 B.n782 B.n781 10.6151
R2465 B.n782 B.n666 10.6151
R2466 B.n788 B.n666 10.6151
R2467 B.n789 B.n788 10.6151
R2468 B.n790 B.n789 10.6151
R2469 B.n790 B.n664 10.6151
R2470 B.n796 B.n664 10.6151
R2471 B.n797 B.n796 10.6151
R2472 B.n798 B.n797 10.6151
R2473 B.n798 B.n662 10.6151
R2474 B.n804 B.n662 10.6151
R2475 B.n805 B.n804 10.6151
R2476 B.n806 B.n805 10.6151
R2477 B.n806 B.n660 10.6151
R2478 B.n813 B.n812 10.6151
R2479 B.n814 B.n813 10.6151
R2480 B.n814 B.n655 10.6151
R2481 B.n820 B.n655 10.6151
R2482 B.n821 B.n820 10.6151
R2483 B.n822 B.n821 10.6151
R2484 B.n822 B.n653 10.6151
R2485 B.n828 B.n653 10.6151
R2486 B.n829 B.n828 10.6151
R2487 B.n831 B.n649 10.6151
R2488 B.n837 B.n649 10.6151
R2489 B.n838 B.n837 10.6151
R2490 B.n839 B.n838 10.6151
R2491 B.n839 B.n647 10.6151
R2492 B.n845 B.n647 10.6151
R2493 B.n846 B.n845 10.6151
R2494 B.n847 B.n846 10.6151
R2495 B.n847 B.n645 10.6151
R2496 B.n853 B.n645 10.6151
R2497 B.n854 B.n853 10.6151
R2498 B.n855 B.n854 10.6151
R2499 B.n855 B.n643 10.6151
R2500 B.n861 B.n643 10.6151
R2501 B.n862 B.n861 10.6151
R2502 B.n863 B.n862 10.6151
R2503 B.n863 B.n641 10.6151
R2504 B.n869 B.n641 10.6151
R2505 B.n870 B.n869 10.6151
R2506 B.n871 B.n870 10.6151
R2507 B.n871 B.n639 10.6151
R2508 B.n877 B.n639 10.6151
R2509 B.n878 B.n877 10.6151
R2510 B.n879 B.n878 10.6151
R2511 B.n879 B.n637 10.6151
R2512 B.n885 B.n637 10.6151
R2513 B.n886 B.n885 10.6151
R2514 B.n887 B.n886 10.6151
R2515 B.n887 B.n635 10.6151
R2516 B.n893 B.n635 10.6151
R2517 B.n894 B.n893 10.6151
R2518 B.n895 B.n894 10.6151
R2519 B.n895 B.n633 10.6151
R2520 B.n901 B.n633 10.6151
R2521 B.n902 B.n901 10.6151
R2522 B.n903 B.n902 10.6151
R2523 B.n903 B.n631 10.6151
R2524 B.n909 B.n631 10.6151
R2525 B.n910 B.n909 10.6151
R2526 B.n911 B.n910 10.6151
R2527 B.n911 B.n629 10.6151
R2528 B.n917 B.n629 10.6151
R2529 B.n918 B.n917 10.6151
R2530 B.n919 B.n918 10.6151
R2531 B.n919 B.n627 10.6151
R2532 B.n925 B.n627 10.6151
R2533 B.n926 B.n925 10.6151
R2534 B.n927 B.n926 10.6151
R2535 B.n927 B.n625 10.6151
R2536 B.n933 B.n625 10.6151
R2537 B.n934 B.n933 10.6151
R2538 B.n935 B.n934 10.6151
R2539 B.n935 B.n623 10.6151
R2540 B.n941 B.n623 10.6151
R2541 B.n942 B.n941 10.6151
R2542 B.n943 B.n942 10.6151
R2543 B.n943 B.n621 10.6151
R2544 B.n621 B.n620 10.6151
R2545 B.n950 B.n620 10.6151
R2546 B.n951 B.n950 10.6151
R2547 B.n957 B.n956 10.6151
R2548 B.n958 B.n957 10.6151
R2549 B.n958 B.n608 10.6151
R2550 B.n968 B.n608 10.6151
R2551 B.n969 B.n968 10.6151
R2552 B.n970 B.n969 10.6151
R2553 B.n970 B.n600 10.6151
R2554 B.n981 B.n600 10.6151
R2555 B.n982 B.n981 10.6151
R2556 B.n983 B.n982 10.6151
R2557 B.n983 B.n593 10.6151
R2558 B.n993 B.n593 10.6151
R2559 B.n994 B.n993 10.6151
R2560 B.n995 B.n994 10.6151
R2561 B.n995 B.n585 10.6151
R2562 B.n1005 B.n585 10.6151
R2563 B.n1006 B.n1005 10.6151
R2564 B.n1007 B.n1006 10.6151
R2565 B.n1007 B.n577 10.6151
R2566 B.n1017 B.n577 10.6151
R2567 B.n1018 B.n1017 10.6151
R2568 B.n1019 B.n1018 10.6151
R2569 B.n1019 B.n569 10.6151
R2570 B.n1029 B.n569 10.6151
R2571 B.n1030 B.n1029 10.6151
R2572 B.n1031 B.n1030 10.6151
R2573 B.n1031 B.n561 10.6151
R2574 B.n1041 B.n561 10.6151
R2575 B.n1042 B.n1041 10.6151
R2576 B.n1043 B.n1042 10.6151
R2577 B.n1043 B.n553 10.6151
R2578 B.n1053 B.n553 10.6151
R2579 B.n1054 B.n1053 10.6151
R2580 B.n1055 B.n1054 10.6151
R2581 B.n1055 B.n545 10.6151
R2582 B.n1065 B.n545 10.6151
R2583 B.n1066 B.n1065 10.6151
R2584 B.n1067 B.n1066 10.6151
R2585 B.n1067 B.n537 10.6151
R2586 B.n1077 B.n537 10.6151
R2587 B.n1078 B.n1077 10.6151
R2588 B.n1079 B.n1078 10.6151
R2589 B.n1079 B.n529 10.6151
R2590 B.n1089 B.n529 10.6151
R2591 B.n1090 B.n1089 10.6151
R2592 B.n1091 B.n1090 10.6151
R2593 B.n1091 B.n521 10.6151
R2594 B.n1101 B.n521 10.6151
R2595 B.n1102 B.n1101 10.6151
R2596 B.n1103 B.n1102 10.6151
R2597 B.n1103 B.n513 10.6151
R2598 B.n1113 B.n513 10.6151
R2599 B.n1114 B.n1113 10.6151
R2600 B.n1115 B.n1114 10.6151
R2601 B.n1115 B.n505 10.6151
R2602 B.n1126 B.n505 10.6151
R2603 B.n1127 B.n1126 10.6151
R2604 B.n1128 B.n1127 10.6151
R2605 B.n1128 B.n498 10.6151
R2606 B.n1138 B.n498 10.6151
R2607 B.n1139 B.n1138 10.6151
R2608 B.n1140 B.n1139 10.6151
R2609 B.n1140 B.n490 10.6151
R2610 B.n1150 B.n490 10.6151
R2611 B.n1151 B.n1150 10.6151
R2612 B.n1152 B.n1151 10.6151
R2613 B.n1152 B.n482 10.6151
R2614 B.n1162 B.n482 10.6151
R2615 B.n1163 B.n1162 10.6151
R2616 B.n1164 B.n1163 10.6151
R2617 B.n1164 B.n474 10.6151
R2618 B.n1175 B.n474 10.6151
R2619 B.n1176 B.n1175 10.6151
R2620 B.n1177 B.n1176 10.6151
R2621 B.n1177 B.n0 10.6151
R2622 B.n1431 B.n1 10.6151
R2623 B.n1431 B.n1430 10.6151
R2624 B.n1430 B.n1429 10.6151
R2625 B.n1429 B.n10 10.6151
R2626 B.n1423 B.n10 10.6151
R2627 B.n1423 B.n1422 10.6151
R2628 B.n1422 B.n1421 10.6151
R2629 B.n1421 B.n17 10.6151
R2630 B.n1415 B.n17 10.6151
R2631 B.n1415 B.n1414 10.6151
R2632 B.n1414 B.n1413 10.6151
R2633 B.n1413 B.n24 10.6151
R2634 B.n1407 B.n24 10.6151
R2635 B.n1407 B.n1406 10.6151
R2636 B.n1406 B.n1405 10.6151
R2637 B.n1405 B.n31 10.6151
R2638 B.n1399 B.n31 10.6151
R2639 B.n1399 B.n1398 10.6151
R2640 B.n1398 B.n1397 10.6151
R2641 B.n1397 B.n37 10.6151
R2642 B.n1391 B.n37 10.6151
R2643 B.n1391 B.n1390 10.6151
R2644 B.n1390 B.n1389 10.6151
R2645 B.n1389 B.n45 10.6151
R2646 B.n1383 B.n45 10.6151
R2647 B.n1383 B.n1382 10.6151
R2648 B.n1382 B.n1381 10.6151
R2649 B.n1381 B.n52 10.6151
R2650 B.n1375 B.n52 10.6151
R2651 B.n1375 B.n1374 10.6151
R2652 B.n1374 B.n1373 10.6151
R2653 B.n1373 B.n59 10.6151
R2654 B.n1367 B.n59 10.6151
R2655 B.n1367 B.n1366 10.6151
R2656 B.n1366 B.n1365 10.6151
R2657 B.n1365 B.n66 10.6151
R2658 B.n1359 B.n66 10.6151
R2659 B.n1359 B.n1358 10.6151
R2660 B.n1358 B.n1357 10.6151
R2661 B.n1357 B.n73 10.6151
R2662 B.n1351 B.n73 10.6151
R2663 B.n1351 B.n1350 10.6151
R2664 B.n1350 B.n1349 10.6151
R2665 B.n1349 B.n80 10.6151
R2666 B.n1343 B.n80 10.6151
R2667 B.n1343 B.n1342 10.6151
R2668 B.n1342 B.n1341 10.6151
R2669 B.n1341 B.n87 10.6151
R2670 B.n1335 B.n87 10.6151
R2671 B.n1335 B.n1334 10.6151
R2672 B.n1334 B.n1333 10.6151
R2673 B.n1333 B.n94 10.6151
R2674 B.n1327 B.n94 10.6151
R2675 B.n1327 B.n1326 10.6151
R2676 B.n1326 B.n1325 10.6151
R2677 B.n1325 B.n101 10.6151
R2678 B.n1319 B.n101 10.6151
R2679 B.n1319 B.n1318 10.6151
R2680 B.n1318 B.n1317 10.6151
R2681 B.n1317 B.n108 10.6151
R2682 B.n1311 B.n108 10.6151
R2683 B.n1311 B.n1310 10.6151
R2684 B.n1310 B.n1309 10.6151
R2685 B.n1309 B.n115 10.6151
R2686 B.n1303 B.n115 10.6151
R2687 B.n1303 B.n1302 10.6151
R2688 B.n1302 B.n1301 10.6151
R2689 B.n1301 B.n121 10.6151
R2690 B.n1295 B.n121 10.6151
R2691 B.n1295 B.n1294 10.6151
R2692 B.n1294 B.n1293 10.6151
R2693 B.n1293 B.n129 10.6151
R2694 B.n1287 B.n129 10.6151
R2695 B.n1287 B.n1286 10.6151
R2696 B.n1286 B.n1285 10.6151
R2697 B.n329 B.n328 9.36635
R2698 B.n351 B.n350 9.36635
R2699 B.n660 B.n659 9.36635
R2700 B.n831 B.n830 9.36635
R2701 B.t2 B.n480 7.82313
R2702 B.t5 B.n15 7.82313
R2703 B.n1093 B.t4 5.0622
R2704 B.t6 B.n1377 5.0622
R2705 B.t7 B.n547 4.14189
R2706 B.n1354 B.t0 4.14189
R2707 B.n1437 B.n0 2.81026
R2708 B.n1437 B.n1 2.81026
R2709 B.n978 B.t15 2.30127
R2710 B.n123 B.t11 2.30127
R2711 B.n330 B.n329 1.24928
R2712 B.n350 B.n349 1.24928
R2713 B.n812 B.n659 1.24928
R2714 B.n830 B.n829 1.24928
R2715 VN.n100 VN.n99 161.3
R2716 VN.n98 VN.n52 161.3
R2717 VN.n97 VN.n96 161.3
R2718 VN.n95 VN.n53 161.3
R2719 VN.n94 VN.n93 161.3
R2720 VN.n92 VN.n54 161.3
R2721 VN.n91 VN.n90 161.3
R2722 VN.n89 VN.n55 161.3
R2723 VN.n88 VN.n87 161.3
R2724 VN.n86 VN.n56 161.3
R2725 VN.n85 VN.n84 161.3
R2726 VN.n83 VN.n58 161.3
R2727 VN.n82 VN.n81 161.3
R2728 VN.n80 VN.n59 161.3
R2729 VN.n79 VN.n78 161.3
R2730 VN.n77 VN.n60 161.3
R2731 VN.n76 VN.n75 161.3
R2732 VN.n74 VN.n61 161.3
R2733 VN.n73 VN.n72 161.3
R2734 VN.n71 VN.n62 161.3
R2735 VN.n70 VN.n69 161.3
R2736 VN.n68 VN.n63 161.3
R2737 VN.n67 VN.n66 161.3
R2738 VN.n49 VN.n48 161.3
R2739 VN.n47 VN.n1 161.3
R2740 VN.n46 VN.n45 161.3
R2741 VN.n44 VN.n2 161.3
R2742 VN.n43 VN.n42 161.3
R2743 VN.n41 VN.n3 161.3
R2744 VN.n40 VN.n39 161.3
R2745 VN.n38 VN.n4 161.3
R2746 VN.n37 VN.n36 161.3
R2747 VN.n34 VN.n5 161.3
R2748 VN.n33 VN.n32 161.3
R2749 VN.n31 VN.n6 161.3
R2750 VN.n30 VN.n29 161.3
R2751 VN.n28 VN.n7 161.3
R2752 VN.n27 VN.n26 161.3
R2753 VN.n25 VN.n8 161.3
R2754 VN.n24 VN.n23 161.3
R2755 VN.n22 VN.n9 161.3
R2756 VN.n21 VN.n20 161.3
R2757 VN.n19 VN.n10 161.3
R2758 VN.n18 VN.n17 161.3
R2759 VN.n16 VN.n11 161.3
R2760 VN.n15 VN.n14 161.3
R2761 VN.n65 VN.t7 161.114
R2762 VN.n13 VN.t4 161.114
R2763 VN.n8 VN.t3 127.915
R2764 VN.n12 VN.t1 127.915
R2765 VN.n35 VN.t9 127.915
R2766 VN.n0 VN.t6 127.915
R2767 VN.n60 VN.t5 127.915
R2768 VN.n64 VN.t8 127.915
R2769 VN.n57 VN.t2 127.915
R2770 VN.n51 VN.t0 127.915
R2771 VN.n50 VN.n0 81.2593
R2772 VN.n101 VN.n51 81.2593
R2773 VN VN.n101 63.3238
R2774 VN.n13 VN.n12 57.9281
R2775 VN.n65 VN.n64 57.9281
R2776 VN.n42 VN.n2 56.5193
R2777 VN.n93 VN.n53 56.5193
R2778 VN.n21 VN.n10 48.2635
R2779 VN.n29 VN.n6 48.2635
R2780 VN.n73 VN.n62 48.2635
R2781 VN.n81 VN.n58 48.2635
R2782 VN.n17 VN.n10 32.7233
R2783 VN.n33 VN.n6 32.7233
R2784 VN.n69 VN.n62 32.7233
R2785 VN.n85 VN.n58 32.7233
R2786 VN.n16 VN.n15 24.4675
R2787 VN.n17 VN.n16 24.4675
R2788 VN.n22 VN.n21 24.4675
R2789 VN.n23 VN.n22 24.4675
R2790 VN.n23 VN.n8 24.4675
R2791 VN.n27 VN.n8 24.4675
R2792 VN.n28 VN.n27 24.4675
R2793 VN.n29 VN.n28 24.4675
R2794 VN.n34 VN.n33 24.4675
R2795 VN.n36 VN.n34 24.4675
R2796 VN.n40 VN.n4 24.4675
R2797 VN.n41 VN.n40 24.4675
R2798 VN.n42 VN.n41 24.4675
R2799 VN.n46 VN.n2 24.4675
R2800 VN.n47 VN.n46 24.4675
R2801 VN.n48 VN.n47 24.4675
R2802 VN.n69 VN.n68 24.4675
R2803 VN.n68 VN.n67 24.4675
R2804 VN.n81 VN.n80 24.4675
R2805 VN.n80 VN.n79 24.4675
R2806 VN.n79 VN.n60 24.4675
R2807 VN.n75 VN.n60 24.4675
R2808 VN.n75 VN.n74 24.4675
R2809 VN.n74 VN.n73 24.4675
R2810 VN.n93 VN.n92 24.4675
R2811 VN.n92 VN.n91 24.4675
R2812 VN.n91 VN.n55 24.4675
R2813 VN.n87 VN.n86 24.4675
R2814 VN.n86 VN.n85 24.4675
R2815 VN.n99 VN.n98 24.4675
R2816 VN.n98 VN.n97 24.4675
R2817 VN.n97 VN.n53 24.4675
R2818 VN.n15 VN.n12 16.6381
R2819 VN.n36 VN.n35 16.6381
R2820 VN.n67 VN.n64 16.6381
R2821 VN.n87 VN.n57 16.6381
R2822 VN.n48 VN.n0 8.80862
R2823 VN.n99 VN.n51 8.80862
R2824 VN.n35 VN.n4 7.82994
R2825 VN.n57 VN.n55 7.82994
R2826 VN.n66 VN.n65 3.19588
R2827 VN.n14 VN.n13 3.19588
R2828 VN.n101 VN.n100 0.354971
R2829 VN.n50 VN.n49 0.354971
R2830 VN VN.n50 0.26696
R2831 VN.n100 VN.n52 0.189894
R2832 VN.n96 VN.n52 0.189894
R2833 VN.n96 VN.n95 0.189894
R2834 VN.n95 VN.n94 0.189894
R2835 VN.n94 VN.n54 0.189894
R2836 VN.n90 VN.n54 0.189894
R2837 VN.n90 VN.n89 0.189894
R2838 VN.n89 VN.n88 0.189894
R2839 VN.n88 VN.n56 0.189894
R2840 VN.n84 VN.n56 0.189894
R2841 VN.n84 VN.n83 0.189894
R2842 VN.n83 VN.n82 0.189894
R2843 VN.n82 VN.n59 0.189894
R2844 VN.n78 VN.n59 0.189894
R2845 VN.n78 VN.n77 0.189894
R2846 VN.n77 VN.n76 0.189894
R2847 VN.n76 VN.n61 0.189894
R2848 VN.n72 VN.n61 0.189894
R2849 VN.n72 VN.n71 0.189894
R2850 VN.n71 VN.n70 0.189894
R2851 VN.n70 VN.n63 0.189894
R2852 VN.n66 VN.n63 0.189894
R2853 VN.n14 VN.n11 0.189894
R2854 VN.n18 VN.n11 0.189894
R2855 VN.n19 VN.n18 0.189894
R2856 VN.n20 VN.n19 0.189894
R2857 VN.n20 VN.n9 0.189894
R2858 VN.n24 VN.n9 0.189894
R2859 VN.n25 VN.n24 0.189894
R2860 VN.n26 VN.n25 0.189894
R2861 VN.n26 VN.n7 0.189894
R2862 VN.n30 VN.n7 0.189894
R2863 VN.n31 VN.n30 0.189894
R2864 VN.n32 VN.n31 0.189894
R2865 VN.n32 VN.n5 0.189894
R2866 VN.n37 VN.n5 0.189894
R2867 VN.n38 VN.n37 0.189894
R2868 VN.n39 VN.n38 0.189894
R2869 VN.n39 VN.n3 0.189894
R2870 VN.n43 VN.n3 0.189894
R2871 VN.n44 VN.n43 0.189894
R2872 VN.n45 VN.n44 0.189894
R2873 VN.n45 VN.n1 0.189894
R2874 VN.n49 VN.n1 0.189894
R2875 VDD2.n1 VDD2.t5 65.5888
R2876 VDD2.n3 VDD2.n2 63.6431
R2877 VDD2 VDD2.n7 63.6403
R2878 VDD2.n4 VDD2.t9 62.2786
R2879 VDD2.n6 VDD2.n5 61.2159
R2880 VDD2.n1 VDD2.n0 61.2157
R2881 VDD2.n4 VDD2.n3 55.4998
R2882 VDD2.n6 VDD2.n4 3.31084
R2883 VDD2.n7 VDD2.t1 1.0633
R2884 VDD2.n7 VDD2.t2 1.0633
R2885 VDD2.n5 VDD2.t7 1.0633
R2886 VDD2.n5 VDD2.t4 1.0633
R2887 VDD2.n2 VDD2.t0 1.0633
R2888 VDD2.n2 VDD2.t3 1.0633
R2889 VDD2.n0 VDD2.t8 1.0633
R2890 VDD2.n0 VDD2.t6 1.0633
R2891 VDD2 VDD2.n6 0.886276
R2892 VDD2.n3 VDD2.n1 0.77274
C0 VP VN 10.969501f
C1 VDD1 VDD2 2.76788f
C2 VTAIL VDD1 13.465799f
C3 VTAIL VDD2 13.5225f
C4 VDD1 VP 17.6938f
C5 VDD1 VN 0.155457f
C6 VP VDD2 0.70012f
C7 VTAIL VP 17.887901f
C8 VN VDD2 17.154f
C9 VTAIL VN 17.8736f
C10 VDD2 B 9.412612f
C11 VDD1 B 9.405836f
C12 VTAIL B 11.588287f
C13 VN B 23.00062f
C14 VP B 21.51337f
C15 VDD2.t5 B 4.09454f
C16 VDD2.t8 B 0.348735f
C17 VDD2.t6 B 0.348735f
C18 VDD2.n0 B 3.18159f
C19 VDD2.n1 B 1.00659f
C20 VDD2.t0 B 0.348735f
C21 VDD2.t3 B 0.348735f
C22 VDD2.n2 B 3.20618f
C23 VDD2.n3 B 3.59894f
C24 VDD2.t9 B 4.06812f
C25 VDD2.n4 B 3.77684f
C26 VDD2.t7 B 0.348735f
C27 VDD2.t4 B 0.348735f
C28 VDD2.n5 B 3.18159f
C29 VDD2.n6 B 0.51723f
C30 VDD2.t1 B 0.348735f
C31 VDD2.t2 B 0.348735f
C32 VDD2.n7 B 3.20613f
C33 VN.t6 B 2.99577f
C34 VN.n0 B 1.09534f
C35 VN.n1 B 0.016645f
C36 VN.n2 B 0.023835f
C37 VN.n3 B 0.016645f
C38 VN.n4 B 0.020608f
C39 VN.n5 B 0.016645f
C40 VN.n6 B 0.014877f
C41 VN.n7 B 0.016645f
C42 VN.t3 B 2.99577f
C43 VN.n8 B 1.04781f
C44 VN.n9 B 0.016645f
C45 VN.n10 B 0.014877f
C46 VN.n11 B 0.016645f
C47 VN.t1 B 2.99577f
C48 VN.n12 B 1.09227f
C49 VN.t4 B 3.2341f
C50 VN.n13 B 1.04433f
C51 VN.n14 B 0.206222f
C52 VN.n15 B 0.026121f
C53 VN.n16 B 0.031022f
C54 VN.n17 B 0.033572f
C55 VN.n18 B 0.016645f
C56 VN.n19 B 0.016645f
C57 VN.n20 B 0.016645f
C58 VN.n21 B 0.031172f
C59 VN.n22 B 0.031022f
C60 VN.n23 B 0.031022f
C61 VN.n24 B 0.016645f
C62 VN.n25 B 0.016645f
C63 VN.n26 B 0.016645f
C64 VN.n27 B 0.031022f
C65 VN.n28 B 0.031022f
C66 VN.n29 B 0.031172f
C67 VN.n30 B 0.016645f
C68 VN.n31 B 0.016645f
C69 VN.n32 B 0.016645f
C70 VN.n33 B 0.033572f
C71 VN.n34 B 0.031022f
C72 VN.t9 B 2.99577f
C73 VN.n35 B 1.0321f
C74 VN.n36 B 0.026121f
C75 VN.n37 B 0.016645f
C76 VN.n38 B 0.016645f
C77 VN.n39 B 0.016645f
C78 VN.n40 B 0.031022f
C79 VN.n41 B 0.031022f
C80 VN.n42 B 0.024763f
C81 VN.n43 B 0.016645f
C82 VN.n44 B 0.016645f
C83 VN.n45 B 0.016645f
C84 VN.n46 B 0.031022f
C85 VN.n47 B 0.031022f
C86 VN.n48 B 0.02122f
C87 VN.n49 B 0.026865f
C88 VN.n50 B 0.045476f
C89 VN.t0 B 2.99577f
C90 VN.n51 B 1.09534f
C91 VN.n52 B 0.016645f
C92 VN.n53 B 0.023835f
C93 VN.n54 B 0.016645f
C94 VN.n55 B 0.020608f
C95 VN.n56 B 0.016645f
C96 VN.t2 B 2.99577f
C97 VN.n57 B 1.0321f
C98 VN.n58 B 0.014877f
C99 VN.n59 B 0.016645f
C100 VN.t5 B 2.99577f
C101 VN.n60 B 1.04781f
C102 VN.n61 B 0.016645f
C103 VN.n62 B 0.014877f
C104 VN.n63 B 0.016645f
C105 VN.t8 B 2.99577f
C106 VN.n64 B 1.09227f
C107 VN.t7 B 3.2341f
C108 VN.n65 B 1.04433f
C109 VN.n66 B 0.206222f
C110 VN.n67 B 0.026121f
C111 VN.n68 B 0.031022f
C112 VN.n69 B 0.033572f
C113 VN.n70 B 0.016645f
C114 VN.n71 B 0.016645f
C115 VN.n72 B 0.016645f
C116 VN.n73 B 0.031172f
C117 VN.n74 B 0.031022f
C118 VN.n75 B 0.031022f
C119 VN.n76 B 0.016645f
C120 VN.n77 B 0.016645f
C121 VN.n78 B 0.016645f
C122 VN.n79 B 0.031022f
C123 VN.n80 B 0.031022f
C124 VN.n81 B 0.031172f
C125 VN.n82 B 0.016645f
C126 VN.n83 B 0.016645f
C127 VN.n84 B 0.016645f
C128 VN.n85 B 0.033572f
C129 VN.n86 B 0.031022f
C130 VN.n87 B 0.026121f
C131 VN.n88 B 0.016645f
C132 VN.n89 B 0.016645f
C133 VN.n90 B 0.016645f
C134 VN.n91 B 0.031022f
C135 VN.n92 B 0.031022f
C136 VN.n93 B 0.024763f
C137 VN.n94 B 0.016645f
C138 VN.n95 B 0.016645f
C139 VN.n96 B 0.016645f
C140 VN.n97 B 0.031022f
C141 VN.n98 B 0.031022f
C142 VN.n99 B 0.02122f
C143 VN.n100 B 0.026865f
C144 VN.n101 B 1.31607f
C145 VDD1.t1 B 4.14484f
C146 VDD1.t2 B 0.353018f
C147 VDD1.t6 B 0.353018f
C148 VDD1.n0 B 3.22067f
C149 VDD1.n1 B 1.02699f
C150 VDD1.t5 B 4.14483f
C151 VDD1.t0 B 0.353018f
C152 VDD1.t4 B 0.353018f
C153 VDD1.n2 B 3.22067f
C154 VDD1.n3 B 1.01895f
C155 VDD1.t7 B 0.353018f
C156 VDD1.t3 B 0.353018f
C157 VDD1.n4 B 3.24556f
C158 VDD1.n5 B 3.79136f
C159 VDD1.t8 B 0.353018f
C160 VDD1.t9 B 0.353018f
C161 VDD1.n6 B 3.22066f
C162 VDD1.n7 B 3.88556f
C163 VTAIL.t5 B 0.353586f
C164 VTAIL.t8 B 0.353586f
C165 VTAIL.n0 B 3.15278f
C166 VTAIL.n1 B 0.601214f
C167 VTAIL.t11 B 4.02938f
C168 VTAIL.n2 B 0.748485f
C169 VTAIL.t17 B 0.353586f
C170 VTAIL.t15 B 0.353586f
C171 VTAIL.n3 B 3.15278f
C172 VTAIL.n4 B 0.752491f
C173 VTAIL.t13 B 0.353586f
C174 VTAIL.t12 B 0.353586f
C175 VTAIL.n5 B 3.15278f
C176 VTAIL.n6 B 2.57784f
C177 VTAIL.t9 B 0.353586f
C178 VTAIL.t7 B 0.353586f
C179 VTAIL.n7 B 3.15278f
C180 VTAIL.n8 B 2.57783f
C181 VTAIL.t4 B 0.353586f
C182 VTAIL.t1 B 0.353586f
C183 VTAIL.n9 B 3.15278f
C184 VTAIL.n10 B 0.752487f
C185 VTAIL.t2 B 4.0294f
C186 VTAIL.n11 B 0.748462f
C187 VTAIL.t18 B 0.353586f
C188 VTAIL.t19 B 0.353586f
C189 VTAIL.n12 B 3.15278f
C190 VTAIL.n13 B 0.660753f
C191 VTAIL.t16 B 0.353586f
C192 VTAIL.t10 B 0.353586f
C193 VTAIL.n14 B 3.15278f
C194 VTAIL.n15 B 0.752487f
C195 VTAIL.t14 B 4.02938f
C196 VTAIL.n16 B 2.40938f
C197 VTAIL.t3 B 4.02938f
C198 VTAIL.n17 B 2.40938f
C199 VTAIL.t6 B 0.353586f
C200 VTAIL.t0 B 0.353586f
C201 VTAIL.n18 B 3.15278f
C202 VTAIL.n19 B 0.555848f
C203 VP.t6 B 3.0298f
C204 VP.n0 B 1.10778f
C205 VP.n1 B 0.016834f
C206 VP.n2 B 0.024106f
C207 VP.n3 B 0.016834f
C208 VP.n4 B 0.020842f
C209 VP.n5 B 0.016834f
C210 VP.n6 B 0.015046f
C211 VP.n7 B 0.016834f
C212 VP.t5 B 3.0298f
C213 VP.n8 B 1.05971f
C214 VP.n9 B 0.016834f
C215 VP.n10 B 0.015046f
C216 VP.n11 B 0.016834f
C217 VP.t9 B 3.0298f
C218 VP.n12 B 1.04382f
C219 VP.n13 B 0.016834f
C220 VP.n14 B 0.025044f
C221 VP.n15 B 0.016834f
C222 VP.n16 B 0.021461f
C223 VP.t0 B 3.0298f
C224 VP.n17 B 1.10778f
C225 VP.n18 B 0.016834f
C226 VP.n19 B 0.024106f
C227 VP.n20 B 0.016834f
C228 VP.n21 B 0.020842f
C229 VP.n22 B 0.016834f
C230 VP.n23 B 0.015046f
C231 VP.n24 B 0.016834f
C232 VP.t3 B 3.0298f
C233 VP.n25 B 1.05971f
C234 VP.n26 B 0.016834f
C235 VP.n27 B 0.015046f
C236 VP.n28 B 0.016834f
C237 VP.t7 B 3.0298f
C238 VP.n29 B 1.10468f
C239 VP.t8 B 3.27083f
C240 VP.n30 B 1.05619f
C241 VP.n31 B 0.208565f
C242 VP.n32 B 0.026418f
C243 VP.n33 B 0.031375f
C244 VP.n34 B 0.033953f
C245 VP.n35 B 0.016834f
C246 VP.n36 B 0.016834f
C247 VP.n37 B 0.016834f
C248 VP.n38 B 0.031526f
C249 VP.n39 B 0.031375f
C250 VP.n40 B 0.031375f
C251 VP.n41 B 0.016834f
C252 VP.n42 B 0.016834f
C253 VP.n43 B 0.016834f
C254 VP.n44 B 0.031375f
C255 VP.n45 B 0.031375f
C256 VP.n46 B 0.031526f
C257 VP.n47 B 0.016834f
C258 VP.n48 B 0.016834f
C259 VP.n49 B 0.016834f
C260 VP.n50 B 0.033953f
C261 VP.n51 B 0.031375f
C262 VP.t1 B 3.0298f
C263 VP.n52 B 1.04382f
C264 VP.n53 B 0.026418f
C265 VP.n54 B 0.016834f
C266 VP.n55 B 0.016834f
C267 VP.n56 B 0.016834f
C268 VP.n57 B 0.031375f
C269 VP.n58 B 0.031375f
C270 VP.n59 B 0.025044f
C271 VP.n60 B 0.016834f
C272 VP.n61 B 0.016834f
C273 VP.n62 B 0.016834f
C274 VP.n63 B 0.031375f
C275 VP.n64 B 0.031375f
C276 VP.n65 B 0.021461f
C277 VP.n66 B 0.02717f
C278 VP.n67 B 1.32463f
C279 VP.t4 B 3.0298f
C280 VP.n68 B 1.10778f
C281 VP.n69 B 1.33421f
C282 VP.n70 B 0.02717f
C283 VP.n71 B 0.016834f
C284 VP.n72 B 0.031375f
C285 VP.n73 B 0.031375f
C286 VP.n74 B 0.024106f
C287 VP.n75 B 0.016834f
C288 VP.n76 B 0.016834f
C289 VP.n77 B 0.016834f
C290 VP.n78 B 0.031375f
C291 VP.n79 B 0.031375f
C292 VP.n80 B 0.020842f
C293 VP.n81 B 0.016834f
C294 VP.n82 B 0.016834f
C295 VP.n83 B 0.026418f
C296 VP.n84 B 0.031375f
C297 VP.n85 B 0.033953f
C298 VP.n86 B 0.016834f
C299 VP.n87 B 0.016834f
C300 VP.n88 B 0.016834f
C301 VP.n89 B 0.031526f
C302 VP.n90 B 0.031375f
C303 VP.n91 B 0.031375f
C304 VP.n92 B 0.016834f
C305 VP.n93 B 0.016834f
C306 VP.n94 B 0.016834f
C307 VP.n95 B 0.031375f
C308 VP.n96 B 0.031375f
C309 VP.n97 B 0.031526f
C310 VP.n98 B 0.016834f
C311 VP.n99 B 0.016834f
C312 VP.n100 B 0.016834f
C313 VP.n101 B 0.033953f
C314 VP.n102 B 0.031375f
C315 VP.t2 B 3.0298f
C316 VP.n103 B 1.04382f
C317 VP.n104 B 0.026418f
C318 VP.n105 B 0.016834f
C319 VP.n106 B 0.016834f
C320 VP.n107 B 0.016834f
C321 VP.n108 B 0.031375f
C322 VP.n109 B 0.031375f
C323 VP.n110 B 0.025044f
C324 VP.n111 B 0.016834f
C325 VP.n112 B 0.016834f
C326 VP.n113 B 0.016834f
C327 VP.n114 B 0.031375f
C328 VP.n115 B 0.031375f
C329 VP.n116 B 0.021461f
C330 VP.n117 B 0.02717f
C331 VP.n118 B 0.045993f
.ends

