* NGSPICE file created from diff_pair_sample_0711.ext - technology: sky130A

.subckt diff_pair_sample_0711 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 w_n1906_n2668# sky130_fd_pr__pfet_01v8 ad=3.315 pd=17.78 as=3.315 ps=17.78 w=8.5 l=2.01
X1 B.t11 B.t9 B.t10 w_n1906_n2668# sky130_fd_pr__pfet_01v8 ad=3.315 pd=17.78 as=0 ps=0 w=8.5 l=2.01
X2 VDD2.t0 VN.t1 VTAIL.t2 w_n1906_n2668# sky130_fd_pr__pfet_01v8 ad=3.315 pd=17.78 as=3.315 ps=17.78 w=8.5 l=2.01
X3 VDD1.t1 VP.t0 VTAIL.t0 w_n1906_n2668# sky130_fd_pr__pfet_01v8 ad=3.315 pd=17.78 as=3.315 ps=17.78 w=8.5 l=2.01
X4 VDD1.t0 VP.t1 VTAIL.t1 w_n1906_n2668# sky130_fd_pr__pfet_01v8 ad=3.315 pd=17.78 as=3.315 ps=17.78 w=8.5 l=2.01
X5 B.t8 B.t6 B.t7 w_n1906_n2668# sky130_fd_pr__pfet_01v8 ad=3.315 pd=17.78 as=0 ps=0 w=8.5 l=2.01
X6 B.t5 B.t3 B.t4 w_n1906_n2668# sky130_fd_pr__pfet_01v8 ad=3.315 pd=17.78 as=0 ps=0 w=8.5 l=2.01
X7 B.t2 B.t0 B.t1 w_n1906_n2668# sky130_fd_pr__pfet_01v8 ad=3.315 pd=17.78 as=0 ps=0 w=8.5 l=2.01
R0 VN VN.t1 201.434
R1 VN VN.t0 161.042
R2 VTAIL.n1 VTAIL.t2 68.4567
R3 VTAIL.n2 VTAIL.t0 68.4566
R4 VTAIL.n3 VTAIL.t3 68.4565
R5 VTAIL.n0 VTAIL.t1 68.4565
R6 VTAIL.n1 VTAIL.n0 23.7289
R7 VTAIL.n3 VTAIL.n2 21.7117
R8 VTAIL.n2 VTAIL.n1 1.47895
R9 VTAIL VTAIL.n0 1.03283
R10 VTAIL VTAIL.n3 0.446621
R11 VDD2.n0 VDD2.t1 120.156
R12 VDD2.n0 VDD2.t0 85.1354
R13 VDD2 VDD2.n0 0.563
R14 B.n337 B.n336 585
R15 B.n338 B.n53 585
R16 B.n340 B.n339 585
R17 B.n341 B.n52 585
R18 B.n343 B.n342 585
R19 B.n344 B.n51 585
R20 B.n346 B.n345 585
R21 B.n347 B.n50 585
R22 B.n349 B.n348 585
R23 B.n350 B.n49 585
R24 B.n352 B.n351 585
R25 B.n353 B.n48 585
R26 B.n355 B.n354 585
R27 B.n356 B.n47 585
R28 B.n358 B.n357 585
R29 B.n359 B.n46 585
R30 B.n361 B.n360 585
R31 B.n362 B.n45 585
R32 B.n364 B.n363 585
R33 B.n365 B.n44 585
R34 B.n367 B.n366 585
R35 B.n368 B.n43 585
R36 B.n370 B.n369 585
R37 B.n371 B.n42 585
R38 B.n373 B.n372 585
R39 B.n374 B.n41 585
R40 B.n376 B.n375 585
R41 B.n377 B.n40 585
R42 B.n379 B.n378 585
R43 B.n380 B.n39 585
R44 B.n382 B.n381 585
R45 B.n384 B.n36 585
R46 B.n386 B.n385 585
R47 B.n387 B.n35 585
R48 B.n389 B.n388 585
R49 B.n390 B.n34 585
R50 B.n392 B.n391 585
R51 B.n393 B.n33 585
R52 B.n395 B.n394 585
R53 B.n396 B.n29 585
R54 B.n398 B.n397 585
R55 B.n399 B.n28 585
R56 B.n401 B.n400 585
R57 B.n402 B.n27 585
R58 B.n404 B.n403 585
R59 B.n405 B.n26 585
R60 B.n407 B.n406 585
R61 B.n408 B.n25 585
R62 B.n410 B.n409 585
R63 B.n411 B.n24 585
R64 B.n413 B.n412 585
R65 B.n414 B.n23 585
R66 B.n416 B.n415 585
R67 B.n417 B.n22 585
R68 B.n419 B.n418 585
R69 B.n420 B.n21 585
R70 B.n422 B.n421 585
R71 B.n423 B.n20 585
R72 B.n425 B.n424 585
R73 B.n426 B.n19 585
R74 B.n428 B.n427 585
R75 B.n429 B.n18 585
R76 B.n431 B.n430 585
R77 B.n432 B.n17 585
R78 B.n434 B.n433 585
R79 B.n435 B.n16 585
R80 B.n437 B.n436 585
R81 B.n438 B.n15 585
R82 B.n440 B.n439 585
R83 B.n441 B.n14 585
R84 B.n443 B.n442 585
R85 B.n444 B.n13 585
R86 B.n335 B.n54 585
R87 B.n334 B.n333 585
R88 B.n332 B.n55 585
R89 B.n331 B.n330 585
R90 B.n329 B.n56 585
R91 B.n328 B.n327 585
R92 B.n326 B.n57 585
R93 B.n325 B.n324 585
R94 B.n323 B.n58 585
R95 B.n322 B.n321 585
R96 B.n320 B.n59 585
R97 B.n319 B.n318 585
R98 B.n317 B.n60 585
R99 B.n316 B.n315 585
R100 B.n314 B.n61 585
R101 B.n313 B.n312 585
R102 B.n311 B.n62 585
R103 B.n310 B.n309 585
R104 B.n308 B.n63 585
R105 B.n307 B.n306 585
R106 B.n305 B.n64 585
R107 B.n304 B.n303 585
R108 B.n302 B.n65 585
R109 B.n301 B.n300 585
R110 B.n299 B.n66 585
R111 B.n298 B.n297 585
R112 B.n296 B.n67 585
R113 B.n295 B.n294 585
R114 B.n293 B.n68 585
R115 B.n292 B.n291 585
R116 B.n290 B.n69 585
R117 B.n289 B.n288 585
R118 B.n287 B.n70 585
R119 B.n286 B.n285 585
R120 B.n284 B.n71 585
R121 B.n283 B.n282 585
R122 B.n281 B.n72 585
R123 B.n280 B.n279 585
R124 B.n278 B.n73 585
R125 B.n277 B.n276 585
R126 B.n275 B.n74 585
R127 B.n274 B.n273 585
R128 B.n272 B.n75 585
R129 B.n271 B.n270 585
R130 B.n269 B.n76 585
R131 B.n160 B.n159 585
R132 B.n161 B.n116 585
R133 B.n163 B.n162 585
R134 B.n164 B.n115 585
R135 B.n166 B.n165 585
R136 B.n167 B.n114 585
R137 B.n169 B.n168 585
R138 B.n170 B.n113 585
R139 B.n172 B.n171 585
R140 B.n173 B.n112 585
R141 B.n175 B.n174 585
R142 B.n176 B.n111 585
R143 B.n178 B.n177 585
R144 B.n179 B.n110 585
R145 B.n181 B.n180 585
R146 B.n182 B.n109 585
R147 B.n184 B.n183 585
R148 B.n185 B.n108 585
R149 B.n187 B.n186 585
R150 B.n188 B.n107 585
R151 B.n190 B.n189 585
R152 B.n191 B.n106 585
R153 B.n193 B.n192 585
R154 B.n194 B.n105 585
R155 B.n196 B.n195 585
R156 B.n197 B.n104 585
R157 B.n199 B.n198 585
R158 B.n200 B.n103 585
R159 B.n202 B.n201 585
R160 B.n203 B.n102 585
R161 B.n205 B.n204 585
R162 B.n207 B.n206 585
R163 B.n208 B.n98 585
R164 B.n210 B.n209 585
R165 B.n211 B.n97 585
R166 B.n213 B.n212 585
R167 B.n214 B.n96 585
R168 B.n216 B.n215 585
R169 B.n217 B.n95 585
R170 B.n219 B.n218 585
R171 B.n220 B.n92 585
R172 B.n223 B.n222 585
R173 B.n224 B.n91 585
R174 B.n226 B.n225 585
R175 B.n227 B.n90 585
R176 B.n229 B.n228 585
R177 B.n230 B.n89 585
R178 B.n232 B.n231 585
R179 B.n233 B.n88 585
R180 B.n235 B.n234 585
R181 B.n236 B.n87 585
R182 B.n238 B.n237 585
R183 B.n239 B.n86 585
R184 B.n241 B.n240 585
R185 B.n242 B.n85 585
R186 B.n244 B.n243 585
R187 B.n245 B.n84 585
R188 B.n247 B.n246 585
R189 B.n248 B.n83 585
R190 B.n250 B.n249 585
R191 B.n251 B.n82 585
R192 B.n253 B.n252 585
R193 B.n254 B.n81 585
R194 B.n256 B.n255 585
R195 B.n257 B.n80 585
R196 B.n259 B.n258 585
R197 B.n260 B.n79 585
R198 B.n262 B.n261 585
R199 B.n263 B.n78 585
R200 B.n265 B.n264 585
R201 B.n266 B.n77 585
R202 B.n268 B.n267 585
R203 B.n158 B.n117 585
R204 B.n157 B.n156 585
R205 B.n155 B.n118 585
R206 B.n154 B.n153 585
R207 B.n152 B.n119 585
R208 B.n151 B.n150 585
R209 B.n149 B.n120 585
R210 B.n148 B.n147 585
R211 B.n146 B.n121 585
R212 B.n145 B.n144 585
R213 B.n143 B.n122 585
R214 B.n142 B.n141 585
R215 B.n140 B.n123 585
R216 B.n139 B.n138 585
R217 B.n137 B.n124 585
R218 B.n136 B.n135 585
R219 B.n134 B.n125 585
R220 B.n133 B.n132 585
R221 B.n131 B.n126 585
R222 B.n130 B.n129 585
R223 B.n128 B.n127 585
R224 B.n2 B.n0 585
R225 B.n477 B.n1 585
R226 B.n476 B.n475 585
R227 B.n474 B.n3 585
R228 B.n473 B.n472 585
R229 B.n471 B.n4 585
R230 B.n470 B.n469 585
R231 B.n468 B.n5 585
R232 B.n467 B.n466 585
R233 B.n465 B.n6 585
R234 B.n464 B.n463 585
R235 B.n462 B.n7 585
R236 B.n461 B.n460 585
R237 B.n459 B.n8 585
R238 B.n458 B.n457 585
R239 B.n456 B.n9 585
R240 B.n455 B.n454 585
R241 B.n453 B.n10 585
R242 B.n452 B.n451 585
R243 B.n450 B.n11 585
R244 B.n449 B.n448 585
R245 B.n447 B.n12 585
R246 B.n446 B.n445 585
R247 B.n479 B.n478 585
R248 B.n159 B.n158 497.305
R249 B.n446 B.n13 497.305
R250 B.n267 B.n76 497.305
R251 B.n337 B.n54 497.305
R252 B.n93 B.t3 308.856
R253 B.n99 B.t0 308.856
R254 B.n30 B.t6 308.856
R255 B.n37 B.t9 308.856
R256 B.n158 B.n157 163.367
R257 B.n157 B.n118 163.367
R258 B.n153 B.n118 163.367
R259 B.n153 B.n152 163.367
R260 B.n152 B.n151 163.367
R261 B.n151 B.n120 163.367
R262 B.n147 B.n120 163.367
R263 B.n147 B.n146 163.367
R264 B.n146 B.n145 163.367
R265 B.n145 B.n122 163.367
R266 B.n141 B.n122 163.367
R267 B.n141 B.n140 163.367
R268 B.n140 B.n139 163.367
R269 B.n139 B.n124 163.367
R270 B.n135 B.n124 163.367
R271 B.n135 B.n134 163.367
R272 B.n134 B.n133 163.367
R273 B.n133 B.n126 163.367
R274 B.n129 B.n126 163.367
R275 B.n129 B.n128 163.367
R276 B.n128 B.n2 163.367
R277 B.n478 B.n2 163.367
R278 B.n478 B.n477 163.367
R279 B.n477 B.n476 163.367
R280 B.n476 B.n3 163.367
R281 B.n472 B.n3 163.367
R282 B.n472 B.n471 163.367
R283 B.n471 B.n470 163.367
R284 B.n470 B.n5 163.367
R285 B.n466 B.n5 163.367
R286 B.n466 B.n465 163.367
R287 B.n465 B.n464 163.367
R288 B.n464 B.n7 163.367
R289 B.n460 B.n7 163.367
R290 B.n460 B.n459 163.367
R291 B.n459 B.n458 163.367
R292 B.n458 B.n9 163.367
R293 B.n454 B.n9 163.367
R294 B.n454 B.n453 163.367
R295 B.n453 B.n452 163.367
R296 B.n452 B.n11 163.367
R297 B.n448 B.n11 163.367
R298 B.n448 B.n447 163.367
R299 B.n447 B.n446 163.367
R300 B.n159 B.n116 163.367
R301 B.n163 B.n116 163.367
R302 B.n164 B.n163 163.367
R303 B.n165 B.n164 163.367
R304 B.n165 B.n114 163.367
R305 B.n169 B.n114 163.367
R306 B.n170 B.n169 163.367
R307 B.n171 B.n170 163.367
R308 B.n171 B.n112 163.367
R309 B.n175 B.n112 163.367
R310 B.n176 B.n175 163.367
R311 B.n177 B.n176 163.367
R312 B.n177 B.n110 163.367
R313 B.n181 B.n110 163.367
R314 B.n182 B.n181 163.367
R315 B.n183 B.n182 163.367
R316 B.n183 B.n108 163.367
R317 B.n187 B.n108 163.367
R318 B.n188 B.n187 163.367
R319 B.n189 B.n188 163.367
R320 B.n189 B.n106 163.367
R321 B.n193 B.n106 163.367
R322 B.n194 B.n193 163.367
R323 B.n195 B.n194 163.367
R324 B.n195 B.n104 163.367
R325 B.n199 B.n104 163.367
R326 B.n200 B.n199 163.367
R327 B.n201 B.n200 163.367
R328 B.n201 B.n102 163.367
R329 B.n205 B.n102 163.367
R330 B.n206 B.n205 163.367
R331 B.n206 B.n98 163.367
R332 B.n210 B.n98 163.367
R333 B.n211 B.n210 163.367
R334 B.n212 B.n211 163.367
R335 B.n212 B.n96 163.367
R336 B.n216 B.n96 163.367
R337 B.n217 B.n216 163.367
R338 B.n218 B.n217 163.367
R339 B.n218 B.n92 163.367
R340 B.n223 B.n92 163.367
R341 B.n224 B.n223 163.367
R342 B.n225 B.n224 163.367
R343 B.n225 B.n90 163.367
R344 B.n229 B.n90 163.367
R345 B.n230 B.n229 163.367
R346 B.n231 B.n230 163.367
R347 B.n231 B.n88 163.367
R348 B.n235 B.n88 163.367
R349 B.n236 B.n235 163.367
R350 B.n237 B.n236 163.367
R351 B.n237 B.n86 163.367
R352 B.n241 B.n86 163.367
R353 B.n242 B.n241 163.367
R354 B.n243 B.n242 163.367
R355 B.n243 B.n84 163.367
R356 B.n247 B.n84 163.367
R357 B.n248 B.n247 163.367
R358 B.n249 B.n248 163.367
R359 B.n249 B.n82 163.367
R360 B.n253 B.n82 163.367
R361 B.n254 B.n253 163.367
R362 B.n255 B.n254 163.367
R363 B.n255 B.n80 163.367
R364 B.n259 B.n80 163.367
R365 B.n260 B.n259 163.367
R366 B.n261 B.n260 163.367
R367 B.n261 B.n78 163.367
R368 B.n265 B.n78 163.367
R369 B.n266 B.n265 163.367
R370 B.n267 B.n266 163.367
R371 B.n271 B.n76 163.367
R372 B.n272 B.n271 163.367
R373 B.n273 B.n272 163.367
R374 B.n273 B.n74 163.367
R375 B.n277 B.n74 163.367
R376 B.n278 B.n277 163.367
R377 B.n279 B.n278 163.367
R378 B.n279 B.n72 163.367
R379 B.n283 B.n72 163.367
R380 B.n284 B.n283 163.367
R381 B.n285 B.n284 163.367
R382 B.n285 B.n70 163.367
R383 B.n289 B.n70 163.367
R384 B.n290 B.n289 163.367
R385 B.n291 B.n290 163.367
R386 B.n291 B.n68 163.367
R387 B.n295 B.n68 163.367
R388 B.n296 B.n295 163.367
R389 B.n297 B.n296 163.367
R390 B.n297 B.n66 163.367
R391 B.n301 B.n66 163.367
R392 B.n302 B.n301 163.367
R393 B.n303 B.n302 163.367
R394 B.n303 B.n64 163.367
R395 B.n307 B.n64 163.367
R396 B.n308 B.n307 163.367
R397 B.n309 B.n308 163.367
R398 B.n309 B.n62 163.367
R399 B.n313 B.n62 163.367
R400 B.n314 B.n313 163.367
R401 B.n315 B.n314 163.367
R402 B.n315 B.n60 163.367
R403 B.n319 B.n60 163.367
R404 B.n320 B.n319 163.367
R405 B.n321 B.n320 163.367
R406 B.n321 B.n58 163.367
R407 B.n325 B.n58 163.367
R408 B.n326 B.n325 163.367
R409 B.n327 B.n326 163.367
R410 B.n327 B.n56 163.367
R411 B.n331 B.n56 163.367
R412 B.n332 B.n331 163.367
R413 B.n333 B.n332 163.367
R414 B.n333 B.n54 163.367
R415 B.n442 B.n13 163.367
R416 B.n442 B.n441 163.367
R417 B.n441 B.n440 163.367
R418 B.n440 B.n15 163.367
R419 B.n436 B.n15 163.367
R420 B.n436 B.n435 163.367
R421 B.n435 B.n434 163.367
R422 B.n434 B.n17 163.367
R423 B.n430 B.n17 163.367
R424 B.n430 B.n429 163.367
R425 B.n429 B.n428 163.367
R426 B.n428 B.n19 163.367
R427 B.n424 B.n19 163.367
R428 B.n424 B.n423 163.367
R429 B.n423 B.n422 163.367
R430 B.n422 B.n21 163.367
R431 B.n418 B.n21 163.367
R432 B.n418 B.n417 163.367
R433 B.n417 B.n416 163.367
R434 B.n416 B.n23 163.367
R435 B.n412 B.n23 163.367
R436 B.n412 B.n411 163.367
R437 B.n411 B.n410 163.367
R438 B.n410 B.n25 163.367
R439 B.n406 B.n25 163.367
R440 B.n406 B.n405 163.367
R441 B.n405 B.n404 163.367
R442 B.n404 B.n27 163.367
R443 B.n400 B.n27 163.367
R444 B.n400 B.n399 163.367
R445 B.n399 B.n398 163.367
R446 B.n398 B.n29 163.367
R447 B.n394 B.n29 163.367
R448 B.n394 B.n393 163.367
R449 B.n393 B.n392 163.367
R450 B.n392 B.n34 163.367
R451 B.n388 B.n34 163.367
R452 B.n388 B.n387 163.367
R453 B.n387 B.n386 163.367
R454 B.n386 B.n36 163.367
R455 B.n381 B.n36 163.367
R456 B.n381 B.n380 163.367
R457 B.n380 B.n379 163.367
R458 B.n379 B.n40 163.367
R459 B.n375 B.n40 163.367
R460 B.n375 B.n374 163.367
R461 B.n374 B.n373 163.367
R462 B.n373 B.n42 163.367
R463 B.n369 B.n42 163.367
R464 B.n369 B.n368 163.367
R465 B.n368 B.n367 163.367
R466 B.n367 B.n44 163.367
R467 B.n363 B.n44 163.367
R468 B.n363 B.n362 163.367
R469 B.n362 B.n361 163.367
R470 B.n361 B.n46 163.367
R471 B.n357 B.n46 163.367
R472 B.n357 B.n356 163.367
R473 B.n356 B.n355 163.367
R474 B.n355 B.n48 163.367
R475 B.n351 B.n48 163.367
R476 B.n351 B.n350 163.367
R477 B.n350 B.n349 163.367
R478 B.n349 B.n50 163.367
R479 B.n345 B.n50 163.367
R480 B.n345 B.n344 163.367
R481 B.n344 B.n343 163.367
R482 B.n343 B.n52 163.367
R483 B.n339 B.n52 163.367
R484 B.n339 B.n338 163.367
R485 B.n338 B.n337 163.367
R486 B.n93 B.t5 160.362
R487 B.n37 B.t10 160.362
R488 B.n99 B.t2 160.352
R489 B.n30 B.t7 160.352
R490 B.n94 B.t4 114.98
R491 B.n38 B.t11 114.98
R492 B.n100 B.t1 114.971
R493 B.n31 B.t8 114.971
R494 B.n221 B.n94 59.5399
R495 B.n101 B.n100 59.5399
R496 B.n32 B.n31 59.5399
R497 B.n383 B.n38 59.5399
R498 B.n94 B.n93 45.3823
R499 B.n100 B.n99 45.3823
R500 B.n31 B.n30 45.3823
R501 B.n38 B.n37 45.3823
R502 B.n445 B.n444 32.3127
R503 B.n336 B.n335 32.3127
R504 B.n269 B.n268 32.3127
R505 B.n160 B.n117 32.3127
R506 B B.n479 18.0485
R507 B.n444 B.n443 10.6151
R508 B.n443 B.n14 10.6151
R509 B.n439 B.n14 10.6151
R510 B.n439 B.n438 10.6151
R511 B.n438 B.n437 10.6151
R512 B.n437 B.n16 10.6151
R513 B.n433 B.n16 10.6151
R514 B.n433 B.n432 10.6151
R515 B.n432 B.n431 10.6151
R516 B.n431 B.n18 10.6151
R517 B.n427 B.n18 10.6151
R518 B.n427 B.n426 10.6151
R519 B.n426 B.n425 10.6151
R520 B.n425 B.n20 10.6151
R521 B.n421 B.n20 10.6151
R522 B.n421 B.n420 10.6151
R523 B.n420 B.n419 10.6151
R524 B.n419 B.n22 10.6151
R525 B.n415 B.n22 10.6151
R526 B.n415 B.n414 10.6151
R527 B.n414 B.n413 10.6151
R528 B.n413 B.n24 10.6151
R529 B.n409 B.n24 10.6151
R530 B.n409 B.n408 10.6151
R531 B.n408 B.n407 10.6151
R532 B.n407 B.n26 10.6151
R533 B.n403 B.n26 10.6151
R534 B.n403 B.n402 10.6151
R535 B.n402 B.n401 10.6151
R536 B.n401 B.n28 10.6151
R537 B.n397 B.n396 10.6151
R538 B.n396 B.n395 10.6151
R539 B.n395 B.n33 10.6151
R540 B.n391 B.n33 10.6151
R541 B.n391 B.n390 10.6151
R542 B.n390 B.n389 10.6151
R543 B.n389 B.n35 10.6151
R544 B.n385 B.n35 10.6151
R545 B.n385 B.n384 10.6151
R546 B.n382 B.n39 10.6151
R547 B.n378 B.n39 10.6151
R548 B.n378 B.n377 10.6151
R549 B.n377 B.n376 10.6151
R550 B.n376 B.n41 10.6151
R551 B.n372 B.n41 10.6151
R552 B.n372 B.n371 10.6151
R553 B.n371 B.n370 10.6151
R554 B.n370 B.n43 10.6151
R555 B.n366 B.n43 10.6151
R556 B.n366 B.n365 10.6151
R557 B.n365 B.n364 10.6151
R558 B.n364 B.n45 10.6151
R559 B.n360 B.n45 10.6151
R560 B.n360 B.n359 10.6151
R561 B.n359 B.n358 10.6151
R562 B.n358 B.n47 10.6151
R563 B.n354 B.n47 10.6151
R564 B.n354 B.n353 10.6151
R565 B.n353 B.n352 10.6151
R566 B.n352 B.n49 10.6151
R567 B.n348 B.n49 10.6151
R568 B.n348 B.n347 10.6151
R569 B.n347 B.n346 10.6151
R570 B.n346 B.n51 10.6151
R571 B.n342 B.n51 10.6151
R572 B.n342 B.n341 10.6151
R573 B.n341 B.n340 10.6151
R574 B.n340 B.n53 10.6151
R575 B.n336 B.n53 10.6151
R576 B.n270 B.n269 10.6151
R577 B.n270 B.n75 10.6151
R578 B.n274 B.n75 10.6151
R579 B.n275 B.n274 10.6151
R580 B.n276 B.n275 10.6151
R581 B.n276 B.n73 10.6151
R582 B.n280 B.n73 10.6151
R583 B.n281 B.n280 10.6151
R584 B.n282 B.n281 10.6151
R585 B.n282 B.n71 10.6151
R586 B.n286 B.n71 10.6151
R587 B.n287 B.n286 10.6151
R588 B.n288 B.n287 10.6151
R589 B.n288 B.n69 10.6151
R590 B.n292 B.n69 10.6151
R591 B.n293 B.n292 10.6151
R592 B.n294 B.n293 10.6151
R593 B.n294 B.n67 10.6151
R594 B.n298 B.n67 10.6151
R595 B.n299 B.n298 10.6151
R596 B.n300 B.n299 10.6151
R597 B.n300 B.n65 10.6151
R598 B.n304 B.n65 10.6151
R599 B.n305 B.n304 10.6151
R600 B.n306 B.n305 10.6151
R601 B.n306 B.n63 10.6151
R602 B.n310 B.n63 10.6151
R603 B.n311 B.n310 10.6151
R604 B.n312 B.n311 10.6151
R605 B.n312 B.n61 10.6151
R606 B.n316 B.n61 10.6151
R607 B.n317 B.n316 10.6151
R608 B.n318 B.n317 10.6151
R609 B.n318 B.n59 10.6151
R610 B.n322 B.n59 10.6151
R611 B.n323 B.n322 10.6151
R612 B.n324 B.n323 10.6151
R613 B.n324 B.n57 10.6151
R614 B.n328 B.n57 10.6151
R615 B.n329 B.n328 10.6151
R616 B.n330 B.n329 10.6151
R617 B.n330 B.n55 10.6151
R618 B.n334 B.n55 10.6151
R619 B.n335 B.n334 10.6151
R620 B.n161 B.n160 10.6151
R621 B.n162 B.n161 10.6151
R622 B.n162 B.n115 10.6151
R623 B.n166 B.n115 10.6151
R624 B.n167 B.n166 10.6151
R625 B.n168 B.n167 10.6151
R626 B.n168 B.n113 10.6151
R627 B.n172 B.n113 10.6151
R628 B.n173 B.n172 10.6151
R629 B.n174 B.n173 10.6151
R630 B.n174 B.n111 10.6151
R631 B.n178 B.n111 10.6151
R632 B.n179 B.n178 10.6151
R633 B.n180 B.n179 10.6151
R634 B.n180 B.n109 10.6151
R635 B.n184 B.n109 10.6151
R636 B.n185 B.n184 10.6151
R637 B.n186 B.n185 10.6151
R638 B.n186 B.n107 10.6151
R639 B.n190 B.n107 10.6151
R640 B.n191 B.n190 10.6151
R641 B.n192 B.n191 10.6151
R642 B.n192 B.n105 10.6151
R643 B.n196 B.n105 10.6151
R644 B.n197 B.n196 10.6151
R645 B.n198 B.n197 10.6151
R646 B.n198 B.n103 10.6151
R647 B.n202 B.n103 10.6151
R648 B.n203 B.n202 10.6151
R649 B.n204 B.n203 10.6151
R650 B.n208 B.n207 10.6151
R651 B.n209 B.n208 10.6151
R652 B.n209 B.n97 10.6151
R653 B.n213 B.n97 10.6151
R654 B.n214 B.n213 10.6151
R655 B.n215 B.n214 10.6151
R656 B.n215 B.n95 10.6151
R657 B.n219 B.n95 10.6151
R658 B.n220 B.n219 10.6151
R659 B.n222 B.n91 10.6151
R660 B.n226 B.n91 10.6151
R661 B.n227 B.n226 10.6151
R662 B.n228 B.n227 10.6151
R663 B.n228 B.n89 10.6151
R664 B.n232 B.n89 10.6151
R665 B.n233 B.n232 10.6151
R666 B.n234 B.n233 10.6151
R667 B.n234 B.n87 10.6151
R668 B.n238 B.n87 10.6151
R669 B.n239 B.n238 10.6151
R670 B.n240 B.n239 10.6151
R671 B.n240 B.n85 10.6151
R672 B.n244 B.n85 10.6151
R673 B.n245 B.n244 10.6151
R674 B.n246 B.n245 10.6151
R675 B.n246 B.n83 10.6151
R676 B.n250 B.n83 10.6151
R677 B.n251 B.n250 10.6151
R678 B.n252 B.n251 10.6151
R679 B.n252 B.n81 10.6151
R680 B.n256 B.n81 10.6151
R681 B.n257 B.n256 10.6151
R682 B.n258 B.n257 10.6151
R683 B.n258 B.n79 10.6151
R684 B.n262 B.n79 10.6151
R685 B.n263 B.n262 10.6151
R686 B.n264 B.n263 10.6151
R687 B.n264 B.n77 10.6151
R688 B.n268 B.n77 10.6151
R689 B.n156 B.n117 10.6151
R690 B.n156 B.n155 10.6151
R691 B.n155 B.n154 10.6151
R692 B.n154 B.n119 10.6151
R693 B.n150 B.n119 10.6151
R694 B.n150 B.n149 10.6151
R695 B.n149 B.n148 10.6151
R696 B.n148 B.n121 10.6151
R697 B.n144 B.n121 10.6151
R698 B.n144 B.n143 10.6151
R699 B.n143 B.n142 10.6151
R700 B.n142 B.n123 10.6151
R701 B.n138 B.n123 10.6151
R702 B.n138 B.n137 10.6151
R703 B.n137 B.n136 10.6151
R704 B.n136 B.n125 10.6151
R705 B.n132 B.n125 10.6151
R706 B.n132 B.n131 10.6151
R707 B.n131 B.n130 10.6151
R708 B.n130 B.n127 10.6151
R709 B.n127 B.n0 10.6151
R710 B.n475 B.n1 10.6151
R711 B.n475 B.n474 10.6151
R712 B.n474 B.n473 10.6151
R713 B.n473 B.n4 10.6151
R714 B.n469 B.n4 10.6151
R715 B.n469 B.n468 10.6151
R716 B.n468 B.n467 10.6151
R717 B.n467 B.n6 10.6151
R718 B.n463 B.n6 10.6151
R719 B.n463 B.n462 10.6151
R720 B.n462 B.n461 10.6151
R721 B.n461 B.n8 10.6151
R722 B.n457 B.n8 10.6151
R723 B.n457 B.n456 10.6151
R724 B.n456 B.n455 10.6151
R725 B.n455 B.n10 10.6151
R726 B.n451 B.n10 10.6151
R727 B.n451 B.n450 10.6151
R728 B.n450 B.n449 10.6151
R729 B.n449 B.n12 10.6151
R730 B.n445 B.n12 10.6151
R731 B.n32 B.n28 9.36635
R732 B.n383 B.n382 9.36635
R733 B.n204 B.n101 9.36635
R734 B.n222 B.n221 9.36635
R735 B.n479 B.n0 2.81026
R736 B.n479 B.n1 2.81026
R737 B.n397 B.n32 1.24928
R738 B.n384 B.n383 1.24928
R739 B.n207 B.n101 1.24928
R740 B.n221 B.n220 1.24928
R741 VP.n0 VP.t0 201.242
R742 VP.n0 VP.t1 160.802
R743 VP VP.n0 0.241678
R744 VDD1 VDD1.t0 121.186
R745 VDD1 VDD1.t1 85.6979
C0 VDD2 w_n1906_n2668# 1.48789f
C1 w_n1906_n2668# VN 2.50934f
C2 w_n1906_n2668# VDD1 1.46907f
C3 w_n1906_n2668# VP 2.75086f
C4 VDD2 VN 1.95516f
C5 w_n1906_n2668# VTAIL 2.26466f
C6 w_n1906_n2668# B 7.19079f
C7 VDD2 VDD1 0.604003f
C8 VDD2 VP 0.308327f
C9 VDD2 VTAIL 4.09407f
C10 VDD2 B 1.37706f
C11 VN VDD1 0.148185f
C12 VP VN 4.52554f
C13 VN VTAIL 1.7303f
C14 B VN 0.91241f
C15 VP VDD1 2.11315f
C16 VTAIL VDD1 4.04714f
C17 VP VTAIL 1.74457f
C18 B VDD1 1.3522f
C19 B VP 1.30711f
C20 B VTAIL 2.6572f
C21 VDD2 VSUBS 0.697274f
C22 VDD1 VSUBS 3.896922f
C23 VTAIL VSUBS 0.772713f
C24 VN VSUBS 5.26884f
C25 VP VSUBS 1.373859f
C26 B VSUBS 3.15879f
C27 w_n1906_n2668# VSUBS 63.0124f
C28 VDD1.t1 VSUBS 1.312f
C29 VDD1.t0 VSUBS 1.74765f
C30 VP.t0 VSUBS 2.79015f
C31 VP.t1 VSUBS 2.31461f
C32 VP.n0 VSUBS 4.22313f
C33 B.n0 VSUBS 0.004541f
C34 B.n1 VSUBS 0.004541f
C35 B.n2 VSUBS 0.007181f
C36 B.n3 VSUBS 0.007181f
C37 B.n4 VSUBS 0.007181f
C38 B.n5 VSUBS 0.007181f
C39 B.n6 VSUBS 0.007181f
C40 B.n7 VSUBS 0.007181f
C41 B.n8 VSUBS 0.007181f
C42 B.n9 VSUBS 0.007181f
C43 B.n10 VSUBS 0.007181f
C44 B.n11 VSUBS 0.007181f
C45 B.n12 VSUBS 0.007181f
C46 B.n13 VSUBS 0.016927f
C47 B.n14 VSUBS 0.007181f
C48 B.n15 VSUBS 0.007181f
C49 B.n16 VSUBS 0.007181f
C50 B.n17 VSUBS 0.007181f
C51 B.n18 VSUBS 0.007181f
C52 B.n19 VSUBS 0.007181f
C53 B.n20 VSUBS 0.007181f
C54 B.n21 VSUBS 0.007181f
C55 B.n22 VSUBS 0.007181f
C56 B.n23 VSUBS 0.007181f
C57 B.n24 VSUBS 0.007181f
C58 B.n25 VSUBS 0.007181f
C59 B.n26 VSUBS 0.007181f
C60 B.n27 VSUBS 0.007181f
C61 B.n28 VSUBS 0.006759f
C62 B.n29 VSUBS 0.007181f
C63 B.t8 VSUBS 0.271633f
C64 B.t7 VSUBS 0.288798f
C65 B.t6 VSUBS 0.801474f
C66 B.n30 VSUBS 0.147681f
C67 B.n31 VSUBS 0.070894f
C68 B.n32 VSUBS 0.016639f
C69 B.n33 VSUBS 0.007181f
C70 B.n34 VSUBS 0.007181f
C71 B.n35 VSUBS 0.007181f
C72 B.n36 VSUBS 0.007181f
C73 B.t11 VSUBS 0.271631f
C74 B.t10 VSUBS 0.288796f
C75 B.t9 VSUBS 0.801474f
C76 B.n37 VSUBS 0.147683f
C77 B.n38 VSUBS 0.070896f
C78 B.n39 VSUBS 0.007181f
C79 B.n40 VSUBS 0.007181f
C80 B.n41 VSUBS 0.007181f
C81 B.n42 VSUBS 0.007181f
C82 B.n43 VSUBS 0.007181f
C83 B.n44 VSUBS 0.007181f
C84 B.n45 VSUBS 0.007181f
C85 B.n46 VSUBS 0.007181f
C86 B.n47 VSUBS 0.007181f
C87 B.n48 VSUBS 0.007181f
C88 B.n49 VSUBS 0.007181f
C89 B.n50 VSUBS 0.007181f
C90 B.n51 VSUBS 0.007181f
C91 B.n52 VSUBS 0.007181f
C92 B.n53 VSUBS 0.007181f
C93 B.n54 VSUBS 0.016446f
C94 B.n55 VSUBS 0.007181f
C95 B.n56 VSUBS 0.007181f
C96 B.n57 VSUBS 0.007181f
C97 B.n58 VSUBS 0.007181f
C98 B.n59 VSUBS 0.007181f
C99 B.n60 VSUBS 0.007181f
C100 B.n61 VSUBS 0.007181f
C101 B.n62 VSUBS 0.007181f
C102 B.n63 VSUBS 0.007181f
C103 B.n64 VSUBS 0.007181f
C104 B.n65 VSUBS 0.007181f
C105 B.n66 VSUBS 0.007181f
C106 B.n67 VSUBS 0.007181f
C107 B.n68 VSUBS 0.007181f
C108 B.n69 VSUBS 0.007181f
C109 B.n70 VSUBS 0.007181f
C110 B.n71 VSUBS 0.007181f
C111 B.n72 VSUBS 0.007181f
C112 B.n73 VSUBS 0.007181f
C113 B.n74 VSUBS 0.007181f
C114 B.n75 VSUBS 0.007181f
C115 B.n76 VSUBS 0.016446f
C116 B.n77 VSUBS 0.007181f
C117 B.n78 VSUBS 0.007181f
C118 B.n79 VSUBS 0.007181f
C119 B.n80 VSUBS 0.007181f
C120 B.n81 VSUBS 0.007181f
C121 B.n82 VSUBS 0.007181f
C122 B.n83 VSUBS 0.007181f
C123 B.n84 VSUBS 0.007181f
C124 B.n85 VSUBS 0.007181f
C125 B.n86 VSUBS 0.007181f
C126 B.n87 VSUBS 0.007181f
C127 B.n88 VSUBS 0.007181f
C128 B.n89 VSUBS 0.007181f
C129 B.n90 VSUBS 0.007181f
C130 B.n91 VSUBS 0.007181f
C131 B.n92 VSUBS 0.007181f
C132 B.t4 VSUBS 0.271631f
C133 B.t5 VSUBS 0.288796f
C134 B.t3 VSUBS 0.801474f
C135 B.n93 VSUBS 0.147683f
C136 B.n94 VSUBS 0.070896f
C137 B.n95 VSUBS 0.007181f
C138 B.n96 VSUBS 0.007181f
C139 B.n97 VSUBS 0.007181f
C140 B.n98 VSUBS 0.007181f
C141 B.t1 VSUBS 0.271633f
C142 B.t2 VSUBS 0.288798f
C143 B.t0 VSUBS 0.801474f
C144 B.n99 VSUBS 0.147681f
C145 B.n100 VSUBS 0.070894f
C146 B.n101 VSUBS 0.016639f
C147 B.n102 VSUBS 0.007181f
C148 B.n103 VSUBS 0.007181f
C149 B.n104 VSUBS 0.007181f
C150 B.n105 VSUBS 0.007181f
C151 B.n106 VSUBS 0.007181f
C152 B.n107 VSUBS 0.007181f
C153 B.n108 VSUBS 0.007181f
C154 B.n109 VSUBS 0.007181f
C155 B.n110 VSUBS 0.007181f
C156 B.n111 VSUBS 0.007181f
C157 B.n112 VSUBS 0.007181f
C158 B.n113 VSUBS 0.007181f
C159 B.n114 VSUBS 0.007181f
C160 B.n115 VSUBS 0.007181f
C161 B.n116 VSUBS 0.007181f
C162 B.n117 VSUBS 0.016446f
C163 B.n118 VSUBS 0.007181f
C164 B.n119 VSUBS 0.007181f
C165 B.n120 VSUBS 0.007181f
C166 B.n121 VSUBS 0.007181f
C167 B.n122 VSUBS 0.007181f
C168 B.n123 VSUBS 0.007181f
C169 B.n124 VSUBS 0.007181f
C170 B.n125 VSUBS 0.007181f
C171 B.n126 VSUBS 0.007181f
C172 B.n127 VSUBS 0.007181f
C173 B.n128 VSUBS 0.007181f
C174 B.n129 VSUBS 0.007181f
C175 B.n130 VSUBS 0.007181f
C176 B.n131 VSUBS 0.007181f
C177 B.n132 VSUBS 0.007181f
C178 B.n133 VSUBS 0.007181f
C179 B.n134 VSUBS 0.007181f
C180 B.n135 VSUBS 0.007181f
C181 B.n136 VSUBS 0.007181f
C182 B.n137 VSUBS 0.007181f
C183 B.n138 VSUBS 0.007181f
C184 B.n139 VSUBS 0.007181f
C185 B.n140 VSUBS 0.007181f
C186 B.n141 VSUBS 0.007181f
C187 B.n142 VSUBS 0.007181f
C188 B.n143 VSUBS 0.007181f
C189 B.n144 VSUBS 0.007181f
C190 B.n145 VSUBS 0.007181f
C191 B.n146 VSUBS 0.007181f
C192 B.n147 VSUBS 0.007181f
C193 B.n148 VSUBS 0.007181f
C194 B.n149 VSUBS 0.007181f
C195 B.n150 VSUBS 0.007181f
C196 B.n151 VSUBS 0.007181f
C197 B.n152 VSUBS 0.007181f
C198 B.n153 VSUBS 0.007181f
C199 B.n154 VSUBS 0.007181f
C200 B.n155 VSUBS 0.007181f
C201 B.n156 VSUBS 0.007181f
C202 B.n157 VSUBS 0.007181f
C203 B.n158 VSUBS 0.016446f
C204 B.n159 VSUBS 0.016927f
C205 B.n160 VSUBS 0.016927f
C206 B.n161 VSUBS 0.007181f
C207 B.n162 VSUBS 0.007181f
C208 B.n163 VSUBS 0.007181f
C209 B.n164 VSUBS 0.007181f
C210 B.n165 VSUBS 0.007181f
C211 B.n166 VSUBS 0.007181f
C212 B.n167 VSUBS 0.007181f
C213 B.n168 VSUBS 0.007181f
C214 B.n169 VSUBS 0.007181f
C215 B.n170 VSUBS 0.007181f
C216 B.n171 VSUBS 0.007181f
C217 B.n172 VSUBS 0.007181f
C218 B.n173 VSUBS 0.007181f
C219 B.n174 VSUBS 0.007181f
C220 B.n175 VSUBS 0.007181f
C221 B.n176 VSUBS 0.007181f
C222 B.n177 VSUBS 0.007181f
C223 B.n178 VSUBS 0.007181f
C224 B.n179 VSUBS 0.007181f
C225 B.n180 VSUBS 0.007181f
C226 B.n181 VSUBS 0.007181f
C227 B.n182 VSUBS 0.007181f
C228 B.n183 VSUBS 0.007181f
C229 B.n184 VSUBS 0.007181f
C230 B.n185 VSUBS 0.007181f
C231 B.n186 VSUBS 0.007181f
C232 B.n187 VSUBS 0.007181f
C233 B.n188 VSUBS 0.007181f
C234 B.n189 VSUBS 0.007181f
C235 B.n190 VSUBS 0.007181f
C236 B.n191 VSUBS 0.007181f
C237 B.n192 VSUBS 0.007181f
C238 B.n193 VSUBS 0.007181f
C239 B.n194 VSUBS 0.007181f
C240 B.n195 VSUBS 0.007181f
C241 B.n196 VSUBS 0.007181f
C242 B.n197 VSUBS 0.007181f
C243 B.n198 VSUBS 0.007181f
C244 B.n199 VSUBS 0.007181f
C245 B.n200 VSUBS 0.007181f
C246 B.n201 VSUBS 0.007181f
C247 B.n202 VSUBS 0.007181f
C248 B.n203 VSUBS 0.007181f
C249 B.n204 VSUBS 0.006759f
C250 B.n205 VSUBS 0.007181f
C251 B.n206 VSUBS 0.007181f
C252 B.n207 VSUBS 0.004013f
C253 B.n208 VSUBS 0.007181f
C254 B.n209 VSUBS 0.007181f
C255 B.n210 VSUBS 0.007181f
C256 B.n211 VSUBS 0.007181f
C257 B.n212 VSUBS 0.007181f
C258 B.n213 VSUBS 0.007181f
C259 B.n214 VSUBS 0.007181f
C260 B.n215 VSUBS 0.007181f
C261 B.n216 VSUBS 0.007181f
C262 B.n217 VSUBS 0.007181f
C263 B.n218 VSUBS 0.007181f
C264 B.n219 VSUBS 0.007181f
C265 B.n220 VSUBS 0.004013f
C266 B.n221 VSUBS 0.016639f
C267 B.n222 VSUBS 0.006759f
C268 B.n223 VSUBS 0.007181f
C269 B.n224 VSUBS 0.007181f
C270 B.n225 VSUBS 0.007181f
C271 B.n226 VSUBS 0.007181f
C272 B.n227 VSUBS 0.007181f
C273 B.n228 VSUBS 0.007181f
C274 B.n229 VSUBS 0.007181f
C275 B.n230 VSUBS 0.007181f
C276 B.n231 VSUBS 0.007181f
C277 B.n232 VSUBS 0.007181f
C278 B.n233 VSUBS 0.007181f
C279 B.n234 VSUBS 0.007181f
C280 B.n235 VSUBS 0.007181f
C281 B.n236 VSUBS 0.007181f
C282 B.n237 VSUBS 0.007181f
C283 B.n238 VSUBS 0.007181f
C284 B.n239 VSUBS 0.007181f
C285 B.n240 VSUBS 0.007181f
C286 B.n241 VSUBS 0.007181f
C287 B.n242 VSUBS 0.007181f
C288 B.n243 VSUBS 0.007181f
C289 B.n244 VSUBS 0.007181f
C290 B.n245 VSUBS 0.007181f
C291 B.n246 VSUBS 0.007181f
C292 B.n247 VSUBS 0.007181f
C293 B.n248 VSUBS 0.007181f
C294 B.n249 VSUBS 0.007181f
C295 B.n250 VSUBS 0.007181f
C296 B.n251 VSUBS 0.007181f
C297 B.n252 VSUBS 0.007181f
C298 B.n253 VSUBS 0.007181f
C299 B.n254 VSUBS 0.007181f
C300 B.n255 VSUBS 0.007181f
C301 B.n256 VSUBS 0.007181f
C302 B.n257 VSUBS 0.007181f
C303 B.n258 VSUBS 0.007181f
C304 B.n259 VSUBS 0.007181f
C305 B.n260 VSUBS 0.007181f
C306 B.n261 VSUBS 0.007181f
C307 B.n262 VSUBS 0.007181f
C308 B.n263 VSUBS 0.007181f
C309 B.n264 VSUBS 0.007181f
C310 B.n265 VSUBS 0.007181f
C311 B.n266 VSUBS 0.007181f
C312 B.n267 VSUBS 0.016927f
C313 B.n268 VSUBS 0.016927f
C314 B.n269 VSUBS 0.016446f
C315 B.n270 VSUBS 0.007181f
C316 B.n271 VSUBS 0.007181f
C317 B.n272 VSUBS 0.007181f
C318 B.n273 VSUBS 0.007181f
C319 B.n274 VSUBS 0.007181f
C320 B.n275 VSUBS 0.007181f
C321 B.n276 VSUBS 0.007181f
C322 B.n277 VSUBS 0.007181f
C323 B.n278 VSUBS 0.007181f
C324 B.n279 VSUBS 0.007181f
C325 B.n280 VSUBS 0.007181f
C326 B.n281 VSUBS 0.007181f
C327 B.n282 VSUBS 0.007181f
C328 B.n283 VSUBS 0.007181f
C329 B.n284 VSUBS 0.007181f
C330 B.n285 VSUBS 0.007181f
C331 B.n286 VSUBS 0.007181f
C332 B.n287 VSUBS 0.007181f
C333 B.n288 VSUBS 0.007181f
C334 B.n289 VSUBS 0.007181f
C335 B.n290 VSUBS 0.007181f
C336 B.n291 VSUBS 0.007181f
C337 B.n292 VSUBS 0.007181f
C338 B.n293 VSUBS 0.007181f
C339 B.n294 VSUBS 0.007181f
C340 B.n295 VSUBS 0.007181f
C341 B.n296 VSUBS 0.007181f
C342 B.n297 VSUBS 0.007181f
C343 B.n298 VSUBS 0.007181f
C344 B.n299 VSUBS 0.007181f
C345 B.n300 VSUBS 0.007181f
C346 B.n301 VSUBS 0.007181f
C347 B.n302 VSUBS 0.007181f
C348 B.n303 VSUBS 0.007181f
C349 B.n304 VSUBS 0.007181f
C350 B.n305 VSUBS 0.007181f
C351 B.n306 VSUBS 0.007181f
C352 B.n307 VSUBS 0.007181f
C353 B.n308 VSUBS 0.007181f
C354 B.n309 VSUBS 0.007181f
C355 B.n310 VSUBS 0.007181f
C356 B.n311 VSUBS 0.007181f
C357 B.n312 VSUBS 0.007181f
C358 B.n313 VSUBS 0.007181f
C359 B.n314 VSUBS 0.007181f
C360 B.n315 VSUBS 0.007181f
C361 B.n316 VSUBS 0.007181f
C362 B.n317 VSUBS 0.007181f
C363 B.n318 VSUBS 0.007181f
C364 B.n319 VSUBS 0.007181f
C365 B.n320 VSUBS 0.007181f
C366 B.n321 VSUBS 0.007181f
C367 B.n322 VSUBS 0.007181f
C368 B.n323 VSUBS 0.007181f
C369 B.n324 VSUBS 0.007181f
C370 B.n325 VSUBS 0.007181f
C371 B.n326 VSUBS 0.007181f
C372 B.n327 VSUBS 0.007181f
C373 B.n328 VSUBS 0.007181f
C374 B.n329 VSUBS 0.007181f
C375 B.n330 VSUBS 0.007181f
C376 B.n331 VSUBS 0.007181f
C377 B.n332 VSUBS 0.007181f
C378 B.n333 VSUBS 0.007181f
C379 B.n334 VSUBS 0.007181f
C380 B.n335 VSUBS 0.017303f
C381 B.n336 VSUBS 0.016069f
C382 B.n337 VSUBS 0.016927f
C383 B.n338 VSUBS 0.007181f
C384 B.n339 VSUBS 0.007181f
C385 B.n340 VSUBS 0.007181f
C386 B.n341 VSUBS 0.007181f
C387 B.n342 VSUBS 0.007181f
C388 B.n343 VSUBS 0.007181f
C389 B.n344 VSUBS 0.007181f
C390 B.n345 VSUBS 0.007181f
C391 B.n346 VSUBS 0.007181f
C392 B.n347 VSUBS 0.007181f
C393 B.n348 VSUBS 0.007181f
C394 B.n349 VSUBS 0.007181f
C395 B.n350 VSUBS 0.007181f
C396 B.n351 VSUBS 0.007181f
C397 B.n352 VSUBS 0.007181f
C398 B.n353 VSUBS 0.007181f
C399 B.n354 VSUBS 0.007181f
C400 B.n355 VSUBS 0.007181f
C401 B.n356 VSUBS 0.007181f
C402 B.n357 VSUBS 0.007181f
C403 B.n358 VSUBS 0.007181f
C404 B.n359 VSUBS 0.007181f
C405 B.n360 VSUBS 0.007181f
C406 B.n361 VSUBS 0.007181f
C407 B.n362 VSUBS 0.007181f
C408 B.n363 VSUBS 0.007181f
C409 B.n364 VSUBS 0.007181f
C410 B.n365 VSUBS 0.007181f
C411 B.n366 VSUBS 0.007181f
C412 B.n367 VSUBS 0.007181f
C413 B.n368 VSUBS 0.007181f
C414 B.n369 VSUBS 0.007181f
C415 B.n370 VSUBS 0.007181f
C416 B.n371 VSUBS 0.007181f
C417 B.n372 VSUBS 0.007181f
C418 B.n373 VSUBS 0.007181f
C419 B.n374 VSUBS 0.007181f
C420 B.n375 VSUBS 0.007181f
C421 B.n376 VSUBS 0.007181f
C422 B.n377 VSUBS 0.007181f
C423 B.n378 VSUBS 0.007181f
C424 B.n379 VSUBS 0.007181f
C425 B.n380 VSUBS 0.007181f
C426 B.n381 VSUBS 0.007181f
C427 B.n382 VSUBS 0.006759f
C428 B.n383 VSUBS 0.016639f
C429 B.n384 VSUBS 0.004013f
C430 B.n385 VSUBS 0.007181f
C431 B.n386 VSUBS 0.007181f
C432 B.n387 VSUBS 0.007181f
C433 B.n388 VSUBS 0.007181f
C434 B.n389 VSUBS 0.007181f
C435 B.n390 VSUBS 0.007181f
C436 B.n391 VSUBS 0.007181f
C437 B.n392 VSUBS 0.007181f
C438 B.n393 VSUBS 0.007181f
C439 B.n394 VSUBS 0.007181f
C440 B.n395 VSUBS 0.007181f
C441 B.n396 VSUBS 0.007181f
C442 B.n397 VSUBS 0.004013f
C443 B.n398 VSUBS 0.007181f
C444 B.n399 VSUBS 0.007181f
C445 B.n400 VSUBS 0.007181f
C446 B.n401 VSUBS 0.007181f
C447 B.n402 VSUBS 0.007181f
C448 B.n403 VSUBS 0.007181f
C449 B.n404 VSUBS 0.007181f
C450 B.n405 VSUBS 0.007181f
C451 B.n406 VSUBS 0.007181f
C452 B.n407 VSUBS 0.007181f
C453 B.n408 VSUBS 0.007181f
C454 B.n409 VSUBS 0.007181f
C455 B.n410 VSUBS 0.007181f
C456 B.n411 VSUBS 0.007181f
C457 B.n412 VSUBS 0.007181f
C458 B.n413 VSUBS 0.007181f
C459 B.n414 VSUBS 0.007181f
C460 B.n415 VSUBS 0.007181f
C461 B.n416 VSUBS 0.007181f
C462 B.n417 VSUBS 0.007181f
C463 B.n418 VSUBS 0.007181f
C464 B.n419 VSUBS 0.007181f
C465 B.n420 VSUBS 0.007181f
C466 B.n421 VSUBS 0.007181f
C467 B.n422 VSUBS 0.007181f
C468 B.n423 VSUBS 0.007181f
C469 B.n424 VSUBS 0.007181f
C470 B.n425 VSUBS 0.007181f
C471 B.n426 VSUBS 0.007181f
C472 B.n427 VSUBS 0.007181f
C473 B.n428 VSUBS 0.007181f
C474 B.n429 VSUBS 0.007181f
C475 B.n430 VSUBS 0.007181f
C476 B.n431 VSUBS 0.007181f
C477 B.n432 VSUBS 0.007181f
C478 B.n433 VSUBS 0.007181f
C479 B.n434 VSUBS 0.007181f
C480 B.n435 VSUBS 0.007181f
C481 B.n436 VSUBS 0.007181f
C482 B.n437 VSUBS 0.007181f
C483 B.n438 VSUBS 0.007181f
C484 B.n439 VSUBS 0.007181f
C485 B.n440 VSUBS 0.007181f
C486 B.n441 VSUBS 0.007181f
C487 B.n442 VSUBS 0.007181f
C488 B.n443 VSUBS 0.007181f
C489 B.n444 VSUBS 0.016927f
C490 B.n445 VSUBS 0.016446f
C491 B.n446 VSUBS 0.016446f
C492 B.n447 VSUBS 0.007181f
C493 B.n448 VSUBS 0.007181f
C494 B.n449 VSUBS 0.007181f
C495 B.n450 VSUBS 0.007181f
C496 B.n451 VSUBS 0.007181f
C497 B.n452 VSUBS 0.007181f
C498 B.n453 VSUBS 0.007181f
C499 B.n454 VSUBS 0.007181f
C500 B.n455 VSUBS 0.007181f
C501 B.n456 VSUBS 0.007181f
C502 B.n457 VSUBS 0.007181f
C503 B.n458 VSUBS 0.007181f
C504 B.n459 VSUBS 0.007181f
C505 B.n460 VSUBS 0.007181f
C506 B.n461 VSUBS 0.007181f
C507 B.n462 VSUBS 0.007181f
C508 B.n463 VSUBS 0.007181f
C509 B.n464 VSUBS 0.007181f
C510 B.n465 VSUBS 0.007181f
C511 B.n466 VSUBS 0.007181f
C512 B.n467 VSUBS 0.007181f
C513 B.n468 VSUBS 0.007181f
C514 B.n469 VSUBS 0.007181f
C515 B.n470 VSUBS 0.007181f
C516 B.n471 VSUBS 0.007181f
C517 B.n472 VSUBS 0.007181f
C518 B.n473 VSUBS 0.007181f
C519 B.n474 VSUBS 0.007181f
C520 B.n475 VSUBS 0.007181f
C521 B.n476 VSUBS 0.007181f
C522 B.n477 VSUBS 0.007181f
C523 B.n478 VSUBS 0.007181f
C524 B.n479 VSUBS 0.016261f
C525 VDD2.t1 VSUBS 1.17101f
C526 VDD2.t0 VSUBS 0.890785f
C527 VDD2.n0 VSUBS 1.96753f
C528 VTAIL.t1 VSUBS 1.4343f
C529 VTAIL.n0 VSUBS 1.88463f
C530 VTAIL.t2 VSUBS 1.43431f
C531 VTAIL.n1 VSUBS 1.91946f
C532 VTAIL.t0 VSUBS 1.43431f
C533 VTAIL.n2 VSUBS 1.76192f
C534 VTAIL.t3 VSUBS 1.4343f
C535 VTAIL.n3 VSUBS 1.68131f
C536 VN.t0 VSUBS 1.71353f
C537 VN.t1 VSUBS 2.06892f
.ends

