* NGSPICE file created from diff_pair_sample_1430.ext - technology: sky130A

.subckt diff_pair_sample_1430 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3938_n3902# sky130_fd_pr__pfet_01v8 ad=5.7213 pd=30.12 as=0 ps=0 w=14.67 l=3.38
X1 VTAIL.t11 VN.t0 VDD2.t2 w_n3938_n3902# sky130_fd_pr__pfet_01v8 ad=2.42055 pd=15 as=2.42055 ps=15 w=14.67 l=3.38
X2 VDD1.t5 VP.t0 VTAIL.t3 w_n3938_n3902# sky130_fd_pr__pfet_01v8 ad=5.7213 pd=30.12 as=2.42055 ps=15 w=14.67 l=3.38
X3 VTAIL.t4 VP.t1 VDD1.t4 w_n3938_n3902# sky130_fd_pr__pfet_01v8 ad=2.42055 pd=15 as=2.42055 ps=15 w=14.67 l=3.38
X4 VDD2.t3 VN.t1 VTAIL.t10 w_n3938_n3902# sky130_fd_pr__pfet_01v8 ad=5.7213 pd=30.12 as=2.42055 ps=15 w=14.67 l=3.38
X5 VDD2.t4 VN.t2 VTAIL.t9 w_n3938_n3902# sky130_fd_pr__pfet_01v8 ad=5.7213 pd=30.12 as=2.42055 ps=15 w=14.67 l=3.38
X6 VDD2.t5 VN.t3 VTAIL.t8 w_n3938_n3902# sky130_fd_pr__pfet_01v8 ad=2.42055 pd=15 as=5.7213 ps=30.12 w=14.67 l=3.38
X7 B.t8 B.t6 B.t7 w_n3938_n3902# sky130_fd_pr__pfet_01v8 ad=5.7213 pd=30.12 as=0 ps=0 w=14.67 l=3.38
X8 VDD1.t3 VP.t2 VTAIL.t2 w_n3938_n3902# sky130_fd_pr__pfet_01v8 ad=5.7213 pd=30.12 as=2.42055 ps=15 w=14.67 l=3.38
X9 VDD1.t2 VP.t3 VTAIL.t1 w_n3938_n3902# sky130_fd_pr__pfet_01v8 ad=2.42055 pd=15 as=5.7213 ps=30.12 w=14.67 l=3.38
X10 VTAIL.t5 VP.t4 VDD1.t1 w_n3938_n3902# sky130_fd_pr__pfet_01v8 ad=2.42055 pd=15 as=2.42055 ps=15 w=14.67 l=3.38
X11 VTAIL.t7 VN.t4 VDD2.t1 w_n3938_n3902# sky130_fd_pr__pfet_01v8 ad=2.42055 pd=15 as=2.42055 ps=15 w=14.67 l=3.38
X12 VDD1.t0 VP.t5 VTAIL.t0 w_n3938_n3902# sky130_fd_pr__pfet_01v8 ad=2.42055 pd=15 as=5.7213 ps=30.12 w=14.67 l=3.38
X13 B.t5 B.t3 B.t4 w_n3938_n3902# sky130_fd_pr__pfet_01v8 ad=5.7213 pd=30.12 as=0 ps=0 w=14.67 l=3.38
X14 VDD2.t0 VN.t5 VTAIL.t6 w_n3938_n3902# sky130_fd_pr__pfet_01v8 ad=2.42055 pd=15 as=5.7213 ps=30.12 w=14.67 l=3.38
X15 B.t2 B.t0 B.t1 w_n3938_n3902# sky130_fd_pr__pfet_01v8 ad=5.7213 pd=30.12 as=0 ps=0 w=14.67 l=3.38
R0 B.n459 B.n138 585
R1 B.n458 B.n457 585
R2 B.n456 B.n139 585
R3 B.n455 B.n454 585
R4 B.n453 B.n140 585
R5 B.n452 B.n451 585
R6 B.n450 B.n141 585
R7 B.n449 B.n448 585
R8 B.n447 B.n142 585
R9 B.n446 B.n445 585
R10 B.n444 B.n143 585
R11 B.n443 B.n442 585
R12 B.n441 B.n144 585
R13 B.n440 B.n439 585
R14 B.n438 B.n145 585
R15 B.n437 B.n436 585
R16 B.n435 B.n146 585
R17 B.n434 B.n433 585
R18 B.n432 B.n147 585
R19 B.n431 B.n430 585
R20 B.n429 B.n148 585
R21 B.n428 B.n427 585
R22 B.n426 B.n149 585
R23 B.n425 B.n424 585
R24 B.n423 B.n150 585
R25 B.n422 B.n421 585
R26 B.n420 B.n151 585
R27 B.n419 B.n418 585
R28 B.n417 B.n152 585
R29 B.n416 B.n415 585
R30 B.n414 B.n153 585
R31 B.n413 B.n412 585
R32 B.n411 B.n154 585
R33 B.n410 B.n409 585
R34 B.n408 B.n155 585
R35 B.n407 B.n406 585
R36 B.n405 B.n156 585
R37 B.n404 B.n403 585
R38 B.n402 B.n157 585
R39 B.n401 B.n400 585
R40 B.n399 B.n158 585
R41 B.n398 B.n397 585
R42 B.n396 B.n159 585
R43 B.n395 B.n394 585
R44 B.n393 B.n160 585
R45 B.n392 B.n391 585
R46 B.n390 B.n161 585
R47 B.n389 B.n388 585
R48 B.n387 B.n162 585
R49 B.n386 B.n385 585
R50 B.n381 B.n163 585
R51 B.n380 B.n379 585
R52 B.n378 B.n164 585
R53 B.n377 B.n376 585
R54 B.n375 B.n165 585
R55 B.n374 B.n373 585
R56 B.n372 B.n166 585
R57 B.n371 B.n370 585
R58 B.n369 B.n167 585
R59 B.n367 B.n366 585
R60 B.n365 B.n170 585
R61 B.n364 B.n363 585
R62 B.n362 B.n171 585
R63 B.n361 B.n360 585
R64 B.n359 B.n172 585
R65 B.n358 B.n357 585
R66 B.n356 B.n173 585
R67 B.n355 B.n354 585
R68 B.n353 B.n174 585
R69 B.n352 B.n351 585
R70 B.n350 B.n175 585
R71 B.n349 B.n348 585
R72 B.n347 B.n176 585
R73 B.n346 B.n345 585
R74 B.n344 B.n177 585
R75 B.n343 B.n342 585
R76 B.n341 B.n178 585
R77 B.n340 B.n339 585
R78 B.n338 B.n179 585
R79 B.n337 B.n336 585
R80 B.n335 B.n180 585
R81 B.n334 B.n333 585
R82 B.n332 B.n181 585
R83 B.n331 B.n330 585
R84 B.n329 B.n182 585
R85 B.n328 B.n327 585
R86 B.n326 B.n183 585
R87 B.n325 B.n324 585
R88 B.n323 B.n184 585
R89 B.n322 B.n321 585
R90 B.n320 B.n185 585
R91 B.n319 B.n318 585
R92 B.n317 B.n186 585
R93 B.n316 B.n315 585
R94 B.n314 B.n187 585
R95 B.n313 B.n312 585
R96 B.n311 B.n188 585
R97 B.n310 B.n309 585
R98 B.n308 B.n189 585
R99 B.n307 B.n306 585
R100 B.n305 B.n190 585
R101 B.n304 B.n303 585
R102 B.n302 B.n191 585
R103 B.n301 B.n300 585
R104 B.n299 B.n192 585
R105 B.n298 B.n297 585
R106 B.n296 B.n193 585
R107 B.n295 B.n294 585
R108 B.n461 B.n460 585
R109 B.n462 B.n137 585
R110 B.n464 B.n463 585
R111 B.n465 B.n136 585
R112 B.n467 B.n466 585
R113 B.n468 B.n135 585
R114 B.n470 B.n469 585
R115 B.n471 B.n134 585
R116 B.n473 B.n472 585
R117 B.n474 B.n133 585
R118 B.n476 B.n475 585
R119 B.n477 B.n132 585
R120 B.n479 B.n478 585
R121 B.n480 B.n131 585
R122 B.n482 B.n481 585
R123 B.n483 B.n130 585
R124 B.n485 B.n484 585
R125 B.n486 B.n129 585
R126 B.n488 B.n487 585
R127 B.n489 B.n128 585
R128 B.n491 B.n490 585
R129 B.n492 B.n127 585
R130 B.n494 B.n493 585
R131 B.n495 B.n126 585
R132 B.n497 B.n496 585
R133 B.n498 B.n125 585
R134 B.n500 B.n499 585
R135 B.n501 B.n124 585
R136 B.n503 B.n502 585
R137 B.n504 B.n123 585
R138 B.n506 B.n505 585
R139 B.n507 B.n122 585
R140 B.n509 B.n508 585
R141 B.n510 B.n121 585
R142 B.n512 B.n511 585
R143 B.n513 B.n120 585
R144 B.n515 B.n514 585
R145 B.n516 B.n119 585
R146 B.n518 B.n517 585
R147 B.n519 B.n118 585
R148 B.n521 B.n520 585
R149 B.n522 B.n117 585
R150 B.n524 B.n523 585
R151 B.n525 B.n116 585
R152 B.n527 B.n526 585
R153 B.n528 B.n115 585
R154 B.n530 B.n529 585
R155 B.n531 B.n114 585
R156 B.n533 B.n532 585
R157 B.n534 B.n113 585
R158 B.n536 B.n535 585
R159 B.n537 B.n112 585
R160 B.n539 B.n538 585
R161 B.n540 B.n111 585
R162 B.n542 B.n541 585
R163 B.n543 B.n110 585
R164 B.n545 B.n544 585
R165 B.n546 B.n109 585
R166 B.n548 B.n547 585
R167 B.n549 B.n108 585
R168 B.n551 B.n550 585
R169 B.n552 B.n107 585
R170 B.n554 B.n553 585
R171 B.n555 B.n106 585
R172 B.n557 B.n556 585
R173 B.n558 B.n105 585
R174 B.n560 B.n559 585
R175 B.n561 B.n104 585
R176 B.n563 B.n562 585
R177 B.n564 B.n103 585
R178 B.n566 B.n565 585
R179 B.n567 B.n102 585
R180 B.n569 B.n568 585
R181 B.n570 B.n101 585
R182 B.n572 B.n571 585
R183 B.n573 B.n100 585
R184 B.n575 B.n574 585
R185 B.n576 B.n99 585
R186 B.n578 B.n577 585
R187 B.n579 B.n98 585
R188 B.n581 B.n580 585
R189 B.n582 B.n97 585
R190 B.n584 B.n583 585
R191 B.n585 B.n96 585
R192 B.n587 B.n586 585
R193 B.n588 B.n95 585
R194 B.n590 B.n589 585
R195 B.n591 B.n94 585
R196 B.n593 B.n592 585
R197 B.n594 B.n93 585
R198 B.n596 B.n595 585
R199 B.n597 B.n92 585
R200 B.n599 B.n598 585
R201 B.n600 B.n91 585
R202 B.n602 B.n601 585
R203 B.n603 B.n90 585
R204 B.n605 B.n604 585
R205 B.n606 B.n89 585
R206 B.n608 B.n607 585
R207 B.n609 B.n88 585
R208 B.n611 B.n610 585
R209 B.n612 B.n87 585
R210 B.n614 B.n613 585
R211 B.n615 B.n86 585
R212 B.n779 B.n778 585
R213 B.n777 B.n28 585
R214 B.n776 B.n775 585
R215 B.n774 B.n29 585
R216 B.n773 B.n772 585
R217 B.n771 B.n30 585
R218 B.n770 B.n769 585
R219 B.n768 B.n31 585
R220 B.n767 B.n766 585
R221 B.n765 B.n32 585
R222 B.n764 B.n763 585
R223 B.n762 B.n33 585
R224 B.n761 B.n760 585
R225 B.n759 B.n34 585
R226 B.n758 B.n757 585
R227 B.n756 B.n35 585
R228 B.n755 B.n754 585
R229 B.n753 B.n36 585
R230 B.n752 B.n751 585
R231 B.n750 B.n37 585
R232 B.n749 B.n748 585
R233 B.n747 B.n38 585
R234 B.n746 B.n745 585
R235 B.n744 B.n39 585
R236 B.n743 B.n742 585
R237 B.n741 B.n40 585
R238 B.n740 B.n739 585
R239 B.n738 B.n41 585
R240 B.n737 B.n736 585
R241 B.n735 B.n42 585
R242 B.n734 B.n733 585
R243 B.n732 B.n43 585
R244 B.n731 B.n730 585
R245 B.n729 B.n44 585
R246 B.n728 B.n727 585
R247 B.n726 B.n45 585
R248 B.n725 B.n724 585
R249 B.n723 B.n46 585
R250 B.n722 B.n721 585
R251 B.n720 B.n47 585
R252 B.n719 B.n718 585
R253 B.n717 B.n48 585
R254 B.n716 B.n715 585
R255 B.n714 B.n49 585
R256 B.n713 B.n712 585
R257 B.n711 B.n50 585
R258 B.n710 B.n709 585
R259 B.n708 B.n51 585
R260 B.n707 B.n706 585
R261 B.n705 B.n704 585
R262 B.n703 B.n55 585
R263 B.n702 B.n701 585
R264 B.n700 B.n56 585
R265 B.n699 B.n698 585
R266 B.n697 B.n57 585
R267 B.n696 B.n695 585
R268 B.n694 B.n58 585
R269 B.n693 B.n692 585
R270 B.n691 B.n59 585
R271 B.n689 B.n688 585
R272 B.n687 B.n62 585
R273 B.n686 B.n685 585
R274 B.n684 B.n63 585
R275 B.n683 B.n682 585
R276 B.n681 B.n64 585
R277 B.n680 B.n679 585
R278 B.n678 B.n65 585
R279 B.n677 B.n676 585
R280 B.n675 B.n66 585
R281 B.n674 B.n673 585
R282 B.n672 B.n67 585
R283 B.n671 B.n670 585
R284 B.n669 B.n68 585
R285 B.n668 B.n667 585
R286 B.n666 B.n69 585
R287 B.n665 B.n664 585
R288 B.n663 B.n70 585
R289 B.n662 B.n661 585
R290 B.n660 B.n71 585
R291 B.n659 B.n658 585
R292 B.n657 B.n72 585
R293 B.n656 B.n655 585
R294 B.n654 B.n73 585
R295 B.n653 B.n652 585
R296 B.n651 B.n74 585
R297 B.n650 B.n649 585
R298 B.n648 B.n75 585
R299 B.n647 B.n646 585
R300 B.n645 B.n76 585
R301 B.n644 B.n643 585
R302 B.n642 B.n77 585
R303 B.n641 B.n640 585
R304 B.n639 B.n78 585
R305 B.n638 B.n637 585
R306 B.n636 B.n79 585
R307 B.n635 B.n634 585
R308 B.n633 B.n80 585
R309 B.n632 B.n631 585
R310 B.n630 B.n81 585
R311 B.n629 B.n628 585
R312 B.n627 B.n82 585
R313 B.n626 B.n625 585
R314 B.n624 B.n83 585
R315 B.n623 B.n622 585
R316 B.n621 B.n84 585
R317 B.n620 B.n619 585
R318 B.n618 B.n85 585
R319 B.n617 B.n616 585
R320 B.n780 B.n27 585
R321 B.n782 B.n781 585
R322 B.n783 B.n26 585
R323 B.n785 B.n784 585
R324 B.n786 B.n25 585
R325 B.n788 B.n787 585
R326 B.n789 B.n24 585
R327 B.n791 B.n790 585
R328 B.n792 B.n23 585
R329 B.n794 B.n793 585
R330 B.n795 B.n22 585
R331 B.n797 B.n796 585
R332 B.n798 B.n21 585
R333 B.n800 B.n799 585
R334 B.n801 B.n20 585
R335 B.n803 B.n802 585
R336 B.n804 B.n19 585
R337 B.n806 B.n805 585
R338 B.n807 B.n18 585
R339 B.n809 B.n808 585
R340 B.n810 B.n17 585
R341 B.n812 B.n811 585
R342 B.n813 B.n16 585
R343 B.n815 B.n814 585
R344 B.n816 B.n15 585
R345 B.n818 B.n817 585
R346 B.n819 B.n14 585
R347 B.n821 B.n820 585
R348 B.n822 B.n13 585
R349 B.n824 B.n823 585
R350 B.n825 B.n12 585
R351 B.n827 B.n826 585
R352 B.n828 B.n11 585
R353 B.n830 B.n829 585
R354 B.n831 B.n10 585
R355 B.n833 B.n832 585
R356 B.n834 B.n9 585
R357 B.n836 B.n835 585
R358 B.n837 B.n8 585
R359 B.n839 B.n838 585
R360 B.n840 B.n7 585
R361 B.n842 B.n841 585
R362 B.n843 B.n6 585
R363 B.n845 B.n844 585
R364 B.n846 B.n5 585
R365 B.n848 B.n847 585
R366 B.n849 B.n4 585
R367 B.n851 B.n850 585
R368 B.n852 B.n3 585
R369 B.n854 B.n853 585
R370 B.n855 B.n0 585
R371 B.n2 B.n1 585
R372 B.n220 B.n219 585
R373 B.n221 B.n218 585
R374 B.n223 B.n222 585
R375 B.n224 B.n217 585
R376 B.n226 B.n225 585
R377 B.n227 B.n216 585
R378 B.n229 B.n228 585
R379 B.n230 B.n215 585
R380 B.n232 B.n231 585
R381 B.n233 B.n214 585
R382 B.n235 B.n234 585
R383 B.n236 B.n213 585
R384 B.n238 B.n237 585
R385 B.n239 B.n212 585
R386 B.n241 B.n240 585
R387 B.n242 B.n211 585
R388 B.n244 B.n243 585
R389 B.n245 B.n210 585
R390 B.n247 B.n246 585
R391 B.n248 B.n209 585
R392 B.n250 B.n249 585
R393 B.n251 B.n208 585
R394 B.n253 B.n252 585
R395 B.n254 B.n207 585
R396 B.n256 B.n255 585
R397 B.n257 B.n206 585
R398 B.n259 B.n258 585
R399 B.n260 B.n205 585
R400 B.n262 B.n261 585
R401 B.n263 B.n204 585
R402 B.n265 B.n264 585
R403 B.n266 B.n203 585
R404 B.n268 B.n267 585
R405 B.n269 B.n202 585
R406 B.n271 B.n270 585
R407 B.n272 B.n201 585
R408 B.n274 B.n273 585
R409 B.n275 B.n200 585
R410 B.n277 B.n276 585
R411 B.n278 B.n199 585
R412 B.n280 B.n279 585
R413 B.n281 B.n198 585
R414 B.n283 B.n282 585
R415 B.n284 B.n197 585
R416 B.n286 B.n285 585
R417 B.n287 B.n196 585
R418 B.n289 B.n288 585
R419 B.n290 B.n195 585
R420 B.n292 B.n291 585
R421 B.n293 B.n194 585
R422 B.n294 B.n293 583.793
R423 B.n460 B.n459 583.793
R424 B.n616 B.n615 583.793
R425 B.n778 B.n27 583.793
R426 B.n382 B.t7 495.502
R427 B.n60 B.t11 495.502
R428 B.n168 B.t1 495.502
R429 B.n52 B.t5 495.502
R430 B.n383 B.t8 423.55
R431 B.n61 B.t10 423.55
R432 B.n169 B.t2 423.55
R433 B.n53 B.t4 423.55
R434 B.n168 B.t0 313.582
R435 B.n382 B.t6 313.582
R436 B.n60 B.t9 313.582
R437 B.n52 B.t3 313.582
R438 B.n857 B.n856 256.663
R439 B.n856 B.n855 235.042
R440 B.n856 B.n2 235.042
R441 B.n294 B.n193 163.367
R442 B.n298 B.n193 163.367
R443 B.n299 B.n298 163.367
R444 B.n300 B.n299 163.367
R445 B.n300 B.n191 163.367
R446 B.n304 B.n191 163.367
R447 B.n305 B.n304 163.367
R448 B.n306 B.n305 163.367
R449 B.n306 B.n189 163.367
R450 B.n310 B.n189 163.367
R451 B.n311 B.n310 163.367
R452 B.n312 B.n311 163.367
R453 B.n312 B.n187 163.367
R454 B.n316 B.n187 163.367
R455 B.n317 B.n316 163.367
R456 B.n318 B.n317 163.367
R457 B.n318 B.n185 163.367
R458 B.n322 B.n185 163.367
R459 B.n323 B.n322 163.367
R460 B.n324 B.n323 163.367
R461 B.n324 B.n183 163.367
R462 B.n328 B.n183 163.367
R463 B.n329 B.n328 163.367
R464 B.n330 B.n329 163.367
R465 B.n330 B.n181 163.367
R466 B.n334 B.n181 163.367
R467 B.n335 B.n334 163.367
R468 B.n336 B.n335 163.367
R469 B.n336 B.n179 163.367
R470 B.n340 B.n179 163.367
R471 B.n341 B.n340 163.367
R472 B.n342 B.n341 163.367
R473 B.n342 B.n177 163.367
R474 B.n346 B.n177 163.367
R475 B.n347 B.n346 163.367
R476 B.n348 B.n347 163.367
R477 B.n348 B.n175 163.367
R478 B.n352 B.n175 163.367
R479 B.n353 B.n352 163.367
R480 B.n354 B.n353 163.367
R481 B.n354 B.n173 163.367
R482 B.n358 B.n173 163.367
R483 B.n359 B.n358 163.367
R484 B.n360 B.n359 163.367
R485 B.n360 B.n171 163.367
R486 B.n364 B.n171 163.367
R487 B.n365 B.n364 163.367
R488 B.n366 B.n365 163.367
R489 B.n366 B.n167 163.367
R490 B.n371 B.n167 163.367
R491 B.n372 B.n371 163.367
R492 B.n373 B.n372 163.367
R493 B.n373 B.n165 163.367
R494 B.n377 B.n165 163.367
R495 B.n378 B.n377 163.367
R496 B.n379 B.n378 163.367
R497 B.n379 B.n163 163.367
R498 B.n386 B.n163 163.367
R499 B.n387 B.n386 163.367
R500 B.n388 B.n387 163.367
R501 B.n388 B.n161 163.367
R502 B.n392 B.n161 163.367
R503 B.n393 B.n392 163.367
R504 B.n394 B.n393 163.367
R505 B.n394 B.n159 163.367
R506 B.n398 B.n159 163.367
R507 B.n399 B.n398 163.367
R508 B.n400 B.n399 163.367
R509 B.n400 B.n157 163.367
R510 B.n404 B.n157 163.367
R511 B.n405 B.n404 163.367
R512 B.n406 B.n405 163.367
R513 B.n406 B.n155 163.367
R514 B.n410 B.n155 163.367
R515 B.n411 B.n410 163.367
R516 B.n412 B.n411 163.367
R517 B.n412 B.n153 163.367
R518 B.n416 B.n153 163.367
R519 B.n417 B.n416 163.367
R520 B.n418 B.n417 163.367
R521 B.n418 B.n151 163.367
R522 B.n422 B.n151 163.367
R523 B.n423 B.n422 163.367
R524 B.n424 B.n423 163.367
R525 B.n424 B.n149 163.367
R526 B.n428 B.n149 163.367
R527 B.n429 B.n428 163.367
R528 B.n430 B.n429 163.367
R529 B.n430 B.n147 163.367
R530 B.n434 B.n147 163.367
R531 B.n435 B.n434 163.367
R532 B.n436 B.n435 163.367
R533 B.n436 B.n145 163.367
R534 B.n440 B.n145 163.367
R535 B.n441 B.n440 163.367
R536 B.n442 B.n441 163.367
R537 B.n442 B.n143 163.367
R538 B.n446 B.n143 163.367
R539 B.n447 B.n446 163.367
R540 B.n448 B.n447 163.367
R541 B.n448 B.n141 163.367
R542 B.n452 B.n141 163.367
R543 B.n453 B.n452 163.367
R544 B.n454 B.n453 163.367
R545 B.n454 B.n139 163.367
R546 B.n458 B.n139 163.367
R547 B.n459 B.n458 163.367
R548 B.n615 B.n614 163.367
R549 B.n614 B.n87 163.367
R550 B.n610 B.n87 163.367
R551 B.n610 B.n609 163.367
R552 B.n609 B.n608 163.367
R553 B.n608 B.n89 163.367
R554 B.n604 B.n89 163.367
R555 B.n604 B.n603 163.367
R556 B.n603 B.n602 163.367
R557 B.n602 B.n91 163.367
R558 B.n598 B.n91 163.367
R559 B.n598 B.n597 163.367
R560 B.n597 B.n596 163.367
R561 B.n596 B.n93 163.367
R562 B.n592 B.n93 163.367
R563 B.n592 B.n591 163.367
R564 B.n591 B.n590 163.367
R565 B.n590 B.n95 163.367
R566 B.n586 B.n95 163.367
R567 B.n586 B.n585 163.367
R568 B.n585 B.n584 163.367
R569 B.n584 B.n97 163.367
R570 B.n580 B.n97 163.367
R571 B.n580 B.n579 163.367
R572 B.n579 B.n578 163.367
R573 B.n578 B.n99 163.367
R574 B.n574 B.n99 163.367
R575 B.n574 B.n573 163.367
R576 B.n573 B.n572 163.367
R577 B.n572 B.n101 163.367
R578 B.n568 B.n101 163.367
R579 B.n568 B.n567 163.367
R580 B.n567 B.n566 163.367
R581 B.n566 B.n103 163.367
R582 B.n562 B.n103 163.367
R583 B.n562 B.n561 163.367
R584 B.n561 B.n560 163.367
R585 B.n560 B.n105 163.367
R586 B.n556 B.n105 163.367
R587 B.n556 B.n555 163.367
R588 B.n555 B.n554 163.367
R589 B.n554 B.n107 163.367
R590 B.n550 B.n107 163.367
R591 B.n550 B.n549 163.367
R592 B.n549 B.n548 163.367
R593 B.n548 B.n109 163.367
R594 B.n544 B.n109 163.367
R595 B.n544 B.n543 163.367
R596 B.n543 B.n542 163.367
R597 B.n542 B.n111 163.367
R598 B.n538 B.n111 163.367
R599 B.n538 B.n537 163.367
R600 B.n537 B.n536 163.367
R601 B.n536 B.n113 163.367
R602 B.n532 B.n113 163.367
R603 B.n532 B.n531 163.367
R604 B.n531 B.n530 163.367
R605 B.n530 B.n115 163.367
R606 B.n526 B.n115 163.367
R607 B.n526 B.n525 163.367
R608 B.n525 B.n524 163.367
R609 B.n524 B.n117 163.367
R610 B.n520 B.n117 163.367
R611 B.n520 B.n519 163.367
R612 B.n519 B.n518 163.367
R613 B.n518 B.n119 163.367
R614 B.n514 B.n119 163.367
R615 B.n514 B.n513 163.367
R616 B.n513 B.n512 163.367
R617 B.n512 B.n121 163.367
R618 B.n508 B.n121 163.367
R619 B.n508 B.n507 163.367
R620 B.n507 B.n506 163.367
R621 B.n506 B.n123 163.367
R622 B.n502 B.n123 163.367
R623 B.n502 B.n501 163.367
R624 B.n501 B.n500 163.367
R625 B.n500 B.n125 163.367
R626 B.n496 B.n125 163.367
R627 B.n496 B.n495 163.367
R628 B.n495 B.n494 163.367
R629 B.n494 B.n127 163.367
R630 B.n490 B.n127 163.367
R631 B.n490 B.n489 163.367
R632 B.n489 B.n488 163.367
R633 B.n488 B.n129 163.367
R634 B.n484 B.n129 163.367
R635 B.n484 B.n483 163.367
R636 B.n483 B.n482 163.367
R637 B.n482 B.n131 163.367
R638 B.n478 B.n131 163.367
R639 B.n478 B.n477 163.367
R640 B.n477 B.n476 163.367
R641 B.n476 B.n133 163.367
R642 B.n472 B.n133 163.367
R643 B.n472 B.n471 163.367
R644 B.n471 B.n470 163.367
R645 B.n470 B.n135 163.367
R646 B.n466 B.n135 163.367
R647 B.n466 B.n465 163.367
R648 B.n465 B.n464 163.367
R649 B.n464 B.n137 163.367
R650 B.n460 B.n137 163.367
R651 B.n778 B.n777 163.367
R652 B.n777 B.n776 163.367
R653 B.n776 B.n29 163.367
R654 B.n772 B.n29 163.367
R655 B.n772 B.n771 163.367
R656 B.n771 B.n770 163.367
R657 B.n770 B.n31 163.367
R658 B.n766 B.n31 163.367
R659 B.n766 B.n765 163.367
R660 B.n765 B.n764 163.367
R661 B.n764 B.n33 163.367
R662 B.n760 B.n33 163.367
R663 B.n760 B.n759 163.367
R664 B.n759 B.n758 163.367
R665 B.n758 B.n35 163.367
R666 B.n754 B.n35 163.367
R667 B.n754 B.n753 163.367
R668 B.n753 B.n752 163.367
R669 B.n752 B.n37 163.367
R670 B.n748 B.n37 163.367
R671 B.n748 B.n747 163.367
R672 B.n747 B.n746 163.367
R673 B.n746 B.n39 163.367
R674 B.n742 B.n39 163.367
R675 B.n742 B.n741 163.367
R676 B.n741 B.n740 163.367
R677 B.n740 B.n41 163.367
R678 B.n736 B.n41 163.367
R679 B.n736 B.n735 163.367
R680 B.n735 B.n734 163.367
R681 B.n734 B.n43 163.367
R682 B.n730 B.n43 163.367
R683 B.n730 B.n729 163.367
R684 B.n729 B.n728 163.367
R685 B.n728 B.n45 163.367
R686 B.n724 B.n45 163.367
R687 B.n724 B.n723 163.367
R688 B.n723 B.n722 163.367
R689 B.n722 B.n47 163.367
R690 B.n718 B.n47 163.367
R691 B.n718 B.n717 163.367
R692 B.n717 B.n716 163.367
R693 B.n716 B.n49 163.367
R694 B.n712 B.n49 163.367
R695 B.n712 B.n711 163.367
R696 B.n711 B.n710 163.367
R697 B.n710 B.n51 163.367
R698 B.n706 B.n51 163.367
R699 B.n706 B.n705 163.367
R700 B.n705 B.n55 163.367
R701 B.n701 B.n55 163.367
R702 B.n701 B.n700 163.367
R703 B.n700 B.n699 163.367
R704 B.n699 B.n57 163.367
R705 B.n695 B.n57 163.367
R706 B.n695 B.n694 163.367
R707 B.n694 B.n693 163.367
R708 B.n693 B.n59 163.367
R709 B.n688 B.n59 163.367
R710 B.n688 B.n687 163.367
R711 B.n687 B.n686 163.367
R712 B.n686 B.n63 163.367
R713 B.n682 B.n63 163.367
R714 B.n682 B.n681 163.367
R715 B.n681 B.n680 163.367
R716 B.n680 B.n65 163.367
R717 B.n676 B.n65 163.367
R718 B.n676 B.n675 163.367
R719 B.n675 B.n674 163.367
R720 B.n674 B.n67 163.367
R721 B.n670 B.n67 163.367
R722 B.n670 B.n669 163.367
R723 B.n669 B.n668 163.367
R724 B.n668 B.n69 163.367
R725 B.n664 B.n69 163.367
R726 B.n664 B.n663 163.367
R727 B.n663 B.n662 163.367
R728 B.n662 B.n71 163.367
R729 B.n658 B.n71 163.367
R730 B.n658 B.n657 163.367
R731 B.n657 B.n656 163.367
R732 B.n656 B.n73 163.367
R733 B.n652 B.n73 163.367
R734 B.n652 B.n651 163.367
R735 B.n651 B.n650 163.367
R736 B.n650 B.n75 163.367
R737 B.n646 B.n75 163.367
R738 B.n646 B.n645 163.367
R739 B.n645 B.n644 163.367
R740 B.n644 B.n77 163.367
R741 B.n640 B.n77 163.367
R742 B.n640 B.n639 163.367
R743 B.n639 B.n638 163.367
R744 B.n638 B.n79 163.367
R745 B.n634 B.n79 163.367
R746 B.n634 B.n633 163.367
R747 B.n633 B.n632 163.367
R748 B.n632 B.n81 163.367
R749 B.n628 B.n81 163.367
R750 B.n628 B.n627 163.367
R751 B.n627 B.n626 163.367
R752 B.n626 B.n83 163.367
R753 B.n622 B.n83 163.367
R754 B.n622 B.n621 163.367
R755 B.n621 B.n620 163.367
R756 B.n620 B.n85 163.367
R757 B.n616 B.n85 163.367
R758 B.n782 B.n27 163.367
R759 B.n783 B.n782 163.367
R760 B.n784 B.n783 163.367
R761 B.n784 B.n25 163.367
R762 B.n788 B.n25 163.367
R763 B.n789 B.n788 163.367
R764 B.n790 B.n789 163.367
R765 B.n790 B.n23 163.367
R766 B.n794 B.n23 163.367
R767 B.n795 B.n794 163.367
R768 B.n796 B.n795 163.367
R769 B.n796 B.n21 163.367
R770 B.n800 B.n21 163.367
R771 B.n801 B.n800 163.367
R772 B.n802 B.n801 163.367
R773 B.n802 B.n19 163.367
R774 B.n806 B.n19 163.367
R775 B.n807 B.n806 163.367
R776 B.n808 B.n807 163.367
R777 B.n808 B.n17 163.367
R778 B.n812 B.n17 163.367
R779 B.n813 B.n812 163.367
R780 B.n814 B.n813 163.367
R781 B.n814 B.n15 163.367
R782 B.n818 B.n15 163.367
R783 B.n819 B.n818 163.367
R784 B.n820 B.n819 163.367
R785 B.n820 B.n13 163.367
R786 B.n824 B.n13 163.367
R787 B.n825 B.n824 163.367
R788 B.n826 B.n825 163.367
R789 B.n826 B.n11 163.367
R790 B.n830 B.n11 163.367
R791 B.n831 B.n830 163.367
R792 B.n832 B.n831 163.367
R793 B.n832 B.n9 163.367
R794 B.n836 B.n9 163.367
R795 B.n837 B.n836 163.367
R796 B.n838 B.n837 163.367
R797 B.n838 B.n7 163.367
R798 B.n842 B.n7 163.367
R799 B.n843 B.n842 163.367
R800 B.n844 B.n843 163.367
R801 B.n844 B.n5 163.367
R802 B.n848 B.n5 163.367
R803 B.n849 B.n848 163.367
R804 B.n850 B.n849 163.367
R805 B.n850 B.n3 163.367
R806 B.n854 B.n3 163.367
R807 B.n855 B.n854 163.367
R808 B.n220 B.n2 163.367
R809 B.n221 B.n220 163.367
R810 B.n222 B.n221 163.367
R811 B.n222 B.n217 163.367
R812 B.n226 B.n217 163.367
R813 B.n227 B.n226 163.367
R814 B.n228 B.n227 163.367
R815 B.n228 B.n215 163.367
R816 B.n232 B.n215 163.367
R817 B.n233 B.n232 163.367
R818 B.n234 B.n233 163.367
R819 B.n234 B.n213 163.367
R820 B.n238 B.n213 163.367
R821 B.n239 B.n238 163.367
R822 B.n240 B.n239 163.367
R823 B.n240 B.n211 163.367
R824 B.n244 B.n211 163.367
R825 B.n245 B.n244 163.367
R826 B.n246 B.n245 163.367
R827 B.n246 B.n209 163.367
R828 B.n250 B.n209 163.367
R829 B.n251 B.n250 163.367
R830 B.n252 B.n251 163.367
R831 B.n252 B.n207 163.367
R832 B.n256 B.n207 163.367
R833 B.n257 B.n256 163.367
R834 B.n258 B.n257 163.367
R835 B.n258 B.n205 163.367
R836 B.n262 B.n205 163.367
R837 B.n263 B.n262 163.367
R838 B.n264 B.n263 163.367
R839 B.n264 B.n203 163.367
R840 B.n268 B.n203 163.367
R841 B.n269 B.n268 163.367
R842 B.n270 B.n269 163.367
R843 B.n270 B.n201 163.367
R844 B.n274 B.n201 163.367
R845 B.n275 B.n274 163.367
R846 B.n276 B.n275 163.367
R847 B.n276 B.n199 163.367
R848 B.n280 B.n199 163.367
R849 B.n281 B.n280 163.367
R850 B.n282 B.n281 163.367
R851 B.n282 B.n197 163.367
R852 B.n286 B.n197 163.367
R853 B.n287 B.n286 163.367
R854 B.n288 B.n287 163.367
R855 B.n288 B.n195 163.367
R856 B.n292 B.n195 163.367
R857 B.n293 B.n292 163.367
R858 B.n169 B.n168 71.952
R859 B.n383 B.n382 71.952
R860 B.n61 B.n60 71.952
R861 B.n53 B.n52 71.952
R862 B.n368 B.n169 59.5399
R863 B.n384 B.n383 59.5399
R864 B.n690 B.n61 59.5399
R865 B.n54 B.n53 59.5399
R866 B.n780 B.n779 37.9322
R867 B.n617 B.n86 37.9322
R868 B.n461 B.n138 37.9322
R869 B.n295 B.n194 37.9322
R870 B B.n857 18.0485
R871 B.n781 B.n780 10.6151
R872 B.n781 B.n26 10.6151
R873 B.n785 B.n26 10.6151
R874 B.n786 B.n785 10.6151
R875 B.n787 B.n786 10.6151
R876 B.n787 B.n24 10.6151
R877 B.n791 B.n24 10.6151
R878 B.n792 B.n791 10.6151
R879 B.n793 B.n792 10.6151
R880 B.n793 B.n22 10.6151
R881 B.n797 B.n22 10.6151
R882 B.n798 B.n797 10.6151
R883 B.n799 B.n798 10.6151
R884 B.n799 B.n20 10.6151
R885 B.n803 B.n20 10.6151
R886 B.n804 B.n803 10.6151
R887 B.n805 B.n804 10.6151
R888 B.n805 B.n18 10.6151
R889 B.n809 B.n18 10.6151
R890 B.n810 B.n809 10.6151
R891 B.n811 B.n810 10.6151
R892 B.n811 B.n16 10.6151
R893 B.n815 B.n16 10.6151
R894 B.n816 B.n815 10.6151
R895 B.n817 B.n816 10.6151
R896 B.n817 B.n14 10.6151
R897 B.n821 B.n14 10.6151
R898 B.n822 B.n821 10.6151
R899 B.n823 B.n822 10.6151
R900 B.n823 B.n12 10.6151
R901 B.n827 B.n12 10.6151
R902 B.n828 B.n827 10.6151
R903 B.n829 B.n828 10.6151
R904 B.n829 B.n10 10.6151
R905 B.n833 B.n10 10.6151
R906 B.n834 B.n833 10.6151
R907 B.n835 B.n834 10.6151
R908 B.n835 B.n8 10.6151
R909 B.n839 B.n8 10.6151
R910 B.n840 B.n839 10.6151
R911 B.n841 B.n840 10.6151
R912 B.n841 B.n6 10.6151
R913 B.n845 B.n6 10.6151
R914 B.n846 B.n845 10.6151
R915 B.n847 B.n846 10.6151
R916 B.n847 B.n4 10.6151
R917 B.n851 B.n4 10.6151
R918 B.n852 B.n851 10.6151
R919 B.n853 B.n852 10.6151
R920 B.n853 B.n0 10.6151
R921 B.n779 B.n28 10.6151
R922 B.n775 B.n28 10.6151
R923 B.n775 B.n774 10.6151
R924 B.n774 B.n773 10.6151
R925 B.n773 B.n30 10.6151
R926 B.n769 B.n30 10.6151
R927 B.n769 B.n768 10.6151
R928 B.n768 B.n767 10.6151
R929 B.n767 B.n32 10.6151
R930 B.n763 B.n32 10.6151
R931 B.n763 B.n762 10.6151
R932 B.n762 B.n761 10.6151
R933 B.n761 B.n34 10.6151
R934 B.n757 B.n34 10.6151
R935 B.n757 B.n756 10.6151
R936 B.n756 B.n755 10.6151
R937 B.n755 B.n36 10.6151
R938 B.n751 B.n36 10.6151
R939 B.n751 B.n750 10.6151
R940 B.n750 B.n749 10.6151
R941 B.n749 B.n38 10.6151
R942 B.n745 B.n38 10.6151
R943 B.n745 B.n744 10.6151
R944 B.n744 B.n743 10.6151
R945 B.n743 B.n40 10.6151
R946 B.n739 B.n40 10.6151
R947 B.n739 B.n738 10.6151
R948 B.n738 B.n737 10.6151
R949 B.n737 B.n42 10.6151
R950 B.n733 B.n42 10.6151
R951 B.n733 B.n732 10.6151
R952 B.n732 B.n731 10.6151
R953 B.n731 B.n44 10.6151
R954 B.n727 B.n44 10.6151
R955 B.n727 B.n726 10.6151
R956 B.n726 B.n725 10.6151
R957 B.n725 B.n46 10.6151
R958 B.n721 B.n46 10.6151
R959 B.n721 B.n720 10.6151
R960 B.n720 B.n719 10.6151
R961 B.n719 B.n48 10.6151
R962 B.n715 B.n48 10.6151
R963 B.n715 B.n714 10.6151
R964 B.n714 B.n713 10.6151
R965 B.n713 B.n50 10.6151
R966 B.n709 B.n50 10.6151
R967 B.n709 B.n708 10.6151
R968 B.n708 B.n707 10.6151
R969 B.n704 B.n703 10.6151
R970 B.n703 B.n702 10.6151
R971 B.n702 B.n56 10.6151
R972 B.n698 B.n56 10.6151
R973 B.n698 B.n697 10.6151
R974 B.n697 B.n696 10.6151
R975 B.n696 B.n58 10.6151
R976 B.n692 B.n58 10.6151
R977 B.n692 B.n691 10.6151
R978 B.n689 B.n62 10.6151
R979 B.n685 B.n62 10.6151
R980 B.n685 B.n684 10.6151
R981 B.n684 B.n683 10.6151
R982 B.n683 B.n64 10.6151
R983 B.n679 B.n64 10.6151
R984 B.n679 B.n678 10.6151
R985 B.n678 B.n677 10.6151
R986 B.n677 B.n66 10.6151
R987 B.n673 B.n66 10.6151
R988 B.n673 B.n672 10.6151
R989 B.n672 B.n671 10.6151
R990 B.n671 B.n68 10.6151
R991 B.n667 B.n68 10.6151
R992 B.n667 B.n666 10.6151
R993 B.n666 B.n665 10.6151
R994 B.n665 B.n70 10.6151
R995 B.n661 B.n70 10.6151
R996 B.n661 B.n660 10.6151
R997 B.n660 B.n659 10.6151
R998 B.n659 B.n72 10.6151
R999 B.n655 B.n72 10.6151
R1000 B.n655 B.n654 10.6151
R1001 B.n654 B.n653 10.6151
R1002 B.n653 B.n74 10.6151
R1003 B.n649 B.n74 10.6151
R1004 B.n649 B.n648 10.6151
R1005 B.n648 B.n647 10.6151
R1006 B.n647 B.n76 10.6151
R1007 B.n643 B.n76 10.6151
R1008 B.n643 B.n642 10.6151
R1009 B.n642 B.n641 10.6151
R1010 B.n641 B.n78 10.6151
R1011 B.n637 B.n78 10.6151
R1012 B.n637 B.n636 10.6151
R1013 B.n636 B.n635 10.6151
R1014 B.n635 B.n80 10.6151
R1015 B.n631 B.n80 10.6151
R1016 B.n631 B.n630 10.6151
R1017 B.n630 B.n629 10.6151
R1018 B.n629 B.n82 10.6151
R1019 B.n625 B.n82 10.6151
R1020 B.n625 B.n624 10.6151
R1021 B.n624 B.n623 10.6151
R1022 B.n623 B.n84 10.6151
R1023 B.n619 B.n84 10.6151
R1024 B.n619 B.n618 10.6151
R1025 B.n618 B.n617 10.6151
R1026 B.n613 B.n86 10.6151
R1027 B.n613 B.n612 10.6151
R1028 B.n612 B.n611 10.6151
R1029 B.n611 B.n88 10.6151
R1030 B.n607 B.n88 10.6151
R1031 B.n607 B.n606 10.6151
R1032 B.n606 B.n605 10.6151
R1033 B.n605 B.n90 10.6151
R1034 B.n601 B.n90 10.6151
R1035 B.n601 B.n600 10.6151
R1036 B.n600 B.n599 10.6151
R1037 B.n599 B.n92 10.6151
R1038 B.n595 B.n92 10.6151
R1039 B.n595 B.n594 10.6151
R1040 B.n594 B.n593 10.6151
R1041 B.n593 B.n94 10.6151
R1042 B.n589 B.n94 10.6151
R1043 B.n589 B.n588 10.6151
R1044 B.n588 B.n587 10.6151
R1045 B.n587 B.n96 10.6151
R1046 B.n583 B.n96 10.6151
R1047 B.n583 B.n582 10.6151
R1048 B.n582 B.n581 10.6151
R1049 B.n581 B.n98 10.6151
R1050 B.n577 B.n98 10.6151
R1051 B.n577 B.n576 10.6151
R1052 B.n576 B.n575 10.6151
R1053 B.n575 B.n100 10.6151
R1054 B.n571 B.n100 10.6151
R1055 B.n571 B.n570 10.6151
R1056 B.n570 B.n569 10.6151
R1057 B.n569 B.n102 10.6151
R1058 B.n565 B.n102 10.6151
R1059 B.n565 B.n564 10.6151
R1060 B.n564 B.n563 10.6151
R1061 B.n563 B.n104 10.6151
R1062 B.n559 B.n104 10.6151
R1063 B.n559 B.n558 10.6151
R1064 B.n558 B.n557 10.6151
R1065 B.n557 B.n106 10.6151
R1066 B.n553 B.n106 10.6151
R1067 B.n553 B.n552 10.6151
R1068 B.n552 B.n551 10.6151
R1069 B.n551 B.n108 10.6151
R1070 B.n547 B.n108 10.6151
R1071 B.n547 B.n546 10.6151
R1072 B.n546 B.n545 10.6151
R1073 B.n545 B.n110 10.6151
R1074 B.n541 B.n110 10.6151
R1075 B.n541 B.n540 10.6151
R1076 B.n540 B.n539 10.6151
R1077 B.n539 B.n112 10.6151
R1078 B.n535 B.n112 10.6151
R1079 B.n535 B.n534 10.6151
R1080 B.n534 B.n533 10.6151
R1081 B.n533 B.n114 10.6151
R1082 B.n529 B.n114 10.6151
R1083 B.n529 B.n528 10.6151
R1084 B.n528 B.n527 10.6151
R1085 B.n527 B.n116 10.6151
R1086 B.n523 B.n116 10.6151
R1087 B.n523 B.n522 10.6151
R1088 B.n522 B.n521 10.6151
R1089 B.n521 B.n118 10.6151
R1090 B.n517 B.n118 10.6151
R1091 B.n517 B.n516 10.6151
R1092 B.n516 B.n515 10.6151
R1093 B.n515 B.n120 10.6151
R1094 B.n511 B.n120 10.6151
R1095 B.n511 B.n510 10.6151
R1096 B.n510 B.n509 10.6151
R1097 B.n509 B.n122 10.6151
R1098 B.n505 B.n122 10.6151
R1099 B.n505 B.n504 10.6151
R1100 B.n504 B.n503 10.6151
R1101 B.n503 B.n124 10.6151
R1102 B.n499 B.n124 10.6151
R1103 B.n499 B.n498 10.6151
R1104 B.n498 B.n497 10.6151
R1105 B.n497 B.n126 10.6151
R1106 B.n493 B.n126 10.6151
R1107 B.n493 B.n492 10.6151
R1108 B.n492 B.n491 10.6151
R1109 B.n491 B.n128 10.6151
R1110 B.n487 B.n128 10.6151
R1111 B.n487 B.n486 10.6151
R1112 B.n486 B.n485 10.6151
R1113 B.n485 B.n130 10.6151
R1114 B.n481 B.n130 10.6151
R1115 B.n481 B.n480 10.6151
R1116 B.n480 B.n479 10.6151
R1117 B.n479 B.n132 10.6151
R1118 B.n475 B.n132 10.6151
R1119 B.n475 B.n474 10.6151
R1120 B.n474 B.n473 10.6151
R1121 B.n473 B.n134 10.6151
R1122 B.n469 B.n134 10.6151
R1123 B.n469 B.n468 10.6151
R1124 B.n468 B.n467 10.6151
R1125 B.n467 B.n136 10.6151
R1126 B.n463 B.n136 10.6151
R1127 B.n463 B.n462 10.6151
R1128 B.n462 B.n461 10.6151
R1129 B.n219 B.n1 10.6151
R1130 B.n219 B.n218 10.6151
R1131 B.n223 B.n218 10.6151
R1132 B.n224 B.n223 10.6151
R1133 B.n225 B.n224 10.6151
R1134 B.n225 B.n216 10.6151
R1135 B.n229 B.n216 10.6151
R1136 B.n230 B.n229 10.6151
R1137 B.n231 B.n230 10.6151
R1138 B.n231 B.n214 10.6151
R1139 B.n235 B.n214 10.6151
R1140 B.n236 B.n235 10.6151
R1141 B.n237 B.n236 10.6151
R1142 B.n237 B.n212 10.6151
R1143 B.n241 B.n212 10.6151
R1144 B.n242 B.n241 10.6151
R1145 B.n243 B.n242 10.6151
R1146 B.n243 B.n210 10.6151
R1147 B.n247 B.n210 10.6151
R1148 B.n248 B.n247 10.6151
R1149 B.n249 B.n248 10.6151
R1150 B.n249 B.n208 10.6151
R1151 B.n253 B.n208 10.6151
R1152 B.n254 B.n253 10.6151
R1153 B.n255 B.n254 10.6151
R1154 B.n255 B.n206 10.6151
R1155 B.n259 B.n206 10.6151
R1156 B.n260 B.n259 10.6151
R1157 B.n261 B.n260 10.6151
R1158 B.n261 B.n204 10.6151
R1159 B.n265 B.n204 10.6151
R1160 B.n266 B.n265 10.6151
R1161 B.n267 B.n266 10.6151
R1162 B.n267 B.n202 10.6151
R1163 B.n271 B.n202 10.6151
R1164 B.n272 B.n271 10.6151
R1165 B.n273 B.n272 10.6151
R1166 B.n273 B.n200 10.6151
R1167 B.n277 B.n200 10.6151
R1168 B.n278 B.n277 10.6151
R1169 B.n279 B.n278 10.6151
R1170 B.n279 B.n198 10.6151
R1171 B.n283 B.n198 10.6151
R1172 B.n284 B.n283 10.6151
R1173 B.n285 B.n284 10.6151
R1174 B.n285 B.n196 10.6151
R1175 B.n289 B.n196 10.6151
R1176 B.n290 B.n289 10.6151
R1177 B.n291 B.n290 10.6151
R1178 B.n291 B.n194 10.6151
R1179 B.n296 B.n295 10.6151
R1180 B.n297 B.n296 10.6151
R1181 B.n297 B.n192 10.6151
R1182 B.n301 B.n192 10.6151
R1183 B.n302 B.n301 10.6151
R1184 B.n303 B.n302 10.6151
R1185 B.n303 B.n190 10.6151
R1186 B.n307 B.n190 10.6151
R1187 B.n308 B.n307 10.6151
R1188 B.n309 B.n308 10.6151
R1189 B.n309 B.n188 10.6151
R1190 B.n313 B.n188 10.6151
R1191 B.n314 B.n313 10.6151
R1192 B.n315 B.n314 10.6151
R1193 B.n315 B.n186 10.6151
R1194 B.n319 B.n186 10.6151
R1195 B.n320 B.n319 10.6151
R1196 B.n321 B.n320 10.6151
R1197 B.n321 B.n184 10.6151
R1198 B.n325 B.n184 10.6151
R1199 B.n326 B.n325 10.6151
R1200 B.n327 B.n326 10.6151
R1201 B.n327 B.n182 10.6151
R1202 B.n331 B.n182 10.6151
R1203 B.n332 B.n331 10.6151
R1204 B.n333 B.n332 10.6151
R1205 B.n333 B.n180 10.6151
R1206 B.n337 B.n180 10.6151
R1207 B.n338 B.n337 10.6151
R1208 B.n339 B.n338 10.6151
R1209 B.n339 B.n178 10.6151
R1210 B.n343 B.n178 10.6151
R1211 B.n344 B.n343 10.6151
R1212 B.n345 B.n344 10.6151
R1213 B.n345 B.n176 10.6151
R1214 B.n349 B.n176 10.6151
R1215 B.n350 B.n349 10.6151
R1216 B.n351 B.n350 10.6151
R1217 B.n351 B.n174 10.6151
R1218 B.n355 B.n174 10.6151
R1219 B.n356 B.n355 10.6151
R1220 B.n357 B.n356 10.6151
R1221 B.n357 B.n172 10.6151
R1222 B.n361 B.n172 10.6151
R1223 B.n362 B.n361 10.6151
R1224 B.n363 B.n362 10.6151
R1225 B.n363 B.n170 10.6151
R1226 B.n367 B.n170 10.6151
R1227 B.n370 B.n369 10.6151
R1228 B.n370 B.n166 10.6151
R1229 B.n374 B.n166 10.6151
R1230 B.n375 B.n374 10.6151
R1231 B.n376 B.n375 10.6151
R1232 B.n376 B.n164 10.6151
R1233 B.n380 B.n164 10.6151
R1234 B.n381 B.n380 10.6151
R1235 B.n385 B.n381 10.6151
R1236 B.n389 B.n162 10.6151
R1237 B.n390 B.n389 10.6151
R1238 B.n391 B.n390 10.6151
R1239 B.n391 B.n160 10.6151
R1240 B.n395 B.n160 10.6151
R1241 B.n396 B.n395 10.6151
R1242 B.n397 B.n396 10.6151
R1243 B.n397 B.n158 10.6151
R1244 B.n401 B.n158 10.6151
R1245 B.n402 B.n401 10.6151
R1246 B.n403 B.n402 10.6151
R1247 B.n403 B.n156 10.6151
R1248 B.n407 B.n156 10.6151
R1249 B.n408 B.n407 10.6151
R1250 B.n409 B.n408 10.6151
R1251 B.n409 B.n154 10.6151
R1252 B.n413 B.n154 10.6151
R1253 B.n414 B.n413 10.6151
R1254 B.n415 B.n414 10.6151
R1255 B.n415 B.n152 10.6151
R1256 B.n419 B.n152 10.6151
R1257 B.n420 B.n419 10.6151
R1258 B.n421 B.n420 10.6151
R1259 B.n421 B.n150 10.6151
R1260 B.n425 B.n150 10.6151
R1261 B.n426 B.n425 10.6151
R1262 B.n427 B.n426 10.6151
R1263 B.n427 B.n148 10.6151
R1264 B.n431 B.n148 10.6151
R1265 B.n432 B.n431 10.6151
R1266 B.n433 B.n432 10.6151
R1267 B.n433 B.n146 10.6151
R1268 B.n437 B.n146 10.6151
R1269 B.n438 B.n437 10.6151
R1270 B.n439 B.n438 10.6151
R1271 B.n439 B.n144 10.6151
R1272 B.n443 B.n144 10.6151
R1273 B.n444 B.n443 10.6151
R1274 B.n445 B.n444 10.6151
R1275 B.n445 B.n142 10.6151
R1276 B.n449 B.n142 10.6151
R1277 B.n450 B.n449 10.6151
R1278 B.n451 B.n450 10.6151
R1279 B.n451 B.n140 10.6151
R1280 B.n455 B.n140 10.6151
R1281 B.n456 B.n455 10.6151
R1282 B.n457 B.n456 10.6151
R1283 B.n457 B.n138 10.6151
R1284 B.n707 B.n54 9.36635
R1285 B.n690 B.n689 9.36635
R1286 B.n368 B.n367 9.36635
R1287 B.n384 B.n162 9.36635
R1288 B.n857 B.n0 8.11757
R1289 B.n857 B.n1 8.11757
R1290 B.n704 B.n54 1.24928
R1291 B.n691 B.n690 1.24928
R1292 B.n369 B.n368 1.24928
R1293 B.n385 B.n384 1.24928
R1294 VN.n34 VN.n33 161.3
R1295 VN.n32 VN.n19 161.3
R1296 VN.n31 VN.n30 161.3
R1297 VN.n29 VN.n20 161.3
R1298 VN.n28 VN.n27 161.3
R1299 VN.n26 VN.n21 161.3
R1300 VN.n25 VN.n24 161.3
R1301 VN.n16 VN.n15 161.3
R1302 VN.n14 VN.n1 161.3
R1303 VN.n13 VN.n12 161.3
R1304 VN.n11 VN.n2 161.3
R1305 VN.n10 VN.n9 161.3
R1306 VN.n8 VN.n3 161.3
R1307 VN.n7 VN.n6 161.3
R1308 VN.n23 VN.t3 138.075
R1309 VN.n5 VN.t2 138.075
R1310 VN.n4 VN.t0 104.6
R1311 VN.n0 VN.t5 104.6
R1312 VN.n22 VN.t4 104.6
R1313 VN.n18 VN.t1 104.6
R1314 VN.n17 VN.n0 79.7913
R1315 VN.n35 VN.n18 79.7913
R1316 VN.n9 VN.n2 54.5767
R1317 VN.n27 VN.n20 54.5767
R1318 VN VN.n35 53.9867
R1319 VN.n5 VN.n4 50.1196
R1320 VN.n23 VN.n22 50.1196
R1321 VN.n13 VN.n2 26.41
R1322 VN.n31 VN.n20 26.41
R1323 VN.n7 VN.n4 24.4675
R1324 VN.n8 VN.n7 24.4675
R1325 VN.n9 VN.n8 24.4675
R1326 VN.n14 VN.n13 24.4675
R1327 VN.n15 VN.n14 24.4675
R1328 VN.n27 VN.n26 24.4675
R1329 VN.n26 VN.n25 24.4675
R1330 VN.n25 VN.n22 24.4675
R1331 VN.n33 VN.n32 24.4675
R1332 VN.n32 VN.n31 24.4675
R1333 VN.n15 VN.n0 10.2766
R1334 VN.n33 VN.n18 10.2766
R1335 VN.n24 VN.n23 3.14396
R1336 VN.n6 VN.n5 3.14396
R1337 VN.n35 VN.n34 0.354971
R1338 VN.n17 VN.n16 0.354971
R1339 VN VN.n17 0.26696
R1340 VN.n34 VN.n19 0.189894
R1341 VN.n30 VN.n19 0.189894
R1342 VN.n30 VN.n29 0.189894
R1343 VN.n29 VN.n28 0.189894
R1344 VN.n28 VN.n21 0.189894
R1345 VN.n24 VN.n21 0.189894
R1346 VN.n6 VN.n3 0.189894
R1347 VN.n10 VN.n3 0.189894
R1348 VN.n11 VN.n10 0.189894
R1349 VN.n12 VN.n11 0.189894
R1350 VN.n12 VN.n1 0.189894
R1351 VN.n16 VN.n1 0.189894
R1352 VDD2.n159 VDD2.n83 756.745
R1353 VDD2.n76 VDD2.n0 756.745
R1354 VDD2.n160 VDD2.n159 585
R1355 VDD2.n158 VDD2.n157 585
R1356 VDD2.n156 VDD2.n86 585
R1357 VDD2.n90 VDD2.n87 585
R1358 VDD2.n151 VDD2.n150 585
R1359 VDD2.n149 VDD2.n148 585
R1360 VDD2.n92 VDD2.n91 585
R1361 VDD2.n143 VDD2.n142 585
R1362 VDD2.n141 VDD2.n140 585
R1363 VDD2.n96 VDD2.n95 585
R1364 VDD2.n135 VDD2.n134 585
R1365 VDD2.n133 VDD2.n132 585
R1366 VDD2.n100 VDD2.n99 585
R1367 VDD2.n127 VDD2.n126 585
R1368 VDD2.n125 VDD2.n124 585
R1369 VDD2.n104 VDD2.n103 585
R1370 VDD2.n119 VDD2.n118 585
R1371 VDD2.n117 VDD2.n116 585
R1372 VDD2.n108 VDD2.n107 585
R1373 VDD2.n111 VDD2.n110 585
R1374 VDD2.n27 VDD2.n26 585
R1375 VDD2.n24 VDD2.n23 585
R1376 VDD2.n33 VDD2.n32 585
R1377 VDD2.n35 VDD2.n34 585
R1378 VDD2.n20 VDD2.n19 585
R1379 VDD2.n41 VDD2.n40 585
R1380 VDD2.n43 VDD2.n42 585
R1381 VDD2.n16 VDD2.n15 585
R1382 VDD2.n49 VDD2.n48 585
R1383 VDD2.n51 VDD2.n50 585
R1384 VDD2.n12 VDD2.n11 585
R1385 VDD2.n57 VDD2.n56 585
R1386 VDD2.n59 VDD2.n58 585
R1387 VDD2.n8 VDD2.n7 585
R1388 VDD2.n65 VDD2.n64 585
R1389 VDD2.n68 VDD2.n67 585
R1390 VDD2.n66 VDD2.n4 585
R1391 VDD2.n73 VDD2.n3 585
R1392 VDD2.n75 VDD2.n74 585
R1393 VDD2.n77 VDD2.n76 585
R1394 VDD2.t3 VDD2.n109 327.466
R1395 VDD2.t4 VDD2.n25 327.466
R1396 VDD2.n159 VDD2.n158 171.744
R1397 VDD2.n158 VDD2.n86 171.744
R1398 VDD2.n90 VDD2.n86 171.744
R1399 VDD2.n150 VDD2.n90 171.744
R1400 VDD2.n150 VDD2.n149 171.744
R1401 VDD2.n149 VDD2.n91 171.744
R1402 VDD2.n142 VDD2.n91 171.744
R1403 VDD2.n142 VDD2.n141 171.744
R1404 VDD2.n141 VDD2.n95 171.744
R1405 VDD2.n134 VDD2.n95 171.744
R1406 VDD2.n134 VDD2.n133 171.744
R1407 VDD2.n133 VDD2.n99 171.744
R1408 VDD2.n126 VDD2.n99 171.744
R1409 VDD2.n126 VDD2.n125 171.744
R1410 VDD2.n125 VDD2.n103 171.744
R1411 VDD2.n118 VDD2.n103 171.744
R1412 VDD2.n118 VDD2.n117 171.744
R1413 VDD2.n117 VDD2.n107 171.744
R1414 VDD2.n110 VDD2.n107 171.744
R1415 VDD2.n26 VDD2.n23 171.744
R1416 VDD2.n33 VDD2.n23 171.744
R1417 VDD2.n34 VDD2.n33 171.744
R1418 VDD2.n34 VDD2.n19 171.744
R1419 VDD2.n41 VDD2.n19 171.744
R1420 VDD2.n42 VDD2.n41 171.744
R1421 VDD2.n42 VDD2.n15 171.744
R1422 VDD2.n49 VDD2.n15 171.744
R1423 VDD2.n50 VDD2.n49 171.744
R1424 VDD2.n50 VDD2.n11 171.744
R1425 VDD2.n57 VDD2.n11 171.744
R1426 VDD2.n58 VDD2.n57 171.744
R1427 VDD2.n58 VDD2.n7 171.744
R1428 VDD2.n65 VDD2.n7 171.744
R1429 VDD2.n67 VDD2.n65 171.744
R1430 VDD2.n67 VDD2.n66 171.744
R1431 VDD2.n66 VDD2.n3 171.744
R1432 VDD2.n75 VDD2.n3 171.744
R1433 VDD2.n76 VDD2.n75 171.744
R1434 VDD2.n110 VDD2.t3 85.8723
R1435 VDD2.n26 VDD2.t4 85.8723
R1436 VDD2.n82 VDD2.n81 72.0924
R1437 VDD2 VDD2.n165 72.0896
R1438 VDD2.n82 VDD2.n80 51.7893
R1439 VDD2.n164 VDD2.n163 49.446
R1440 VDD2.n164 VDD2.n82 46.7562
R1441 VDD2.n111 VDD2.n109 16.3895
R1442 VDD2.n27 VDD2.n25 16.3895
R1443 VDD2.n157 VDD2.n156 13.1884
R1444 VDD2.n74 VDD2.n73 13.1884
R1445 VDD2.n160 VDD2.n85 12.8005
R1446 VDD2.n155 VDD2.n87 12.8005
R1447 VDD2.n112 VDD2.n108 12.8005
R1448 VDD2.n28 VDD2.n24 12.8005
R1449 VDD2.n72 VDD2.n4 12.8005
R1450 VDD2.n77 VDD2.n2 12.8005
R1451 VDD2.n161 VDD2.n83 12.0247
R1452 VDD2.n152 VDD2.n151 12.0247
R1453 VDD2.n116 VDD2.n115 12.0247
R1454 VDD2.n32 VDD2.n31 12.0247
R1455 VDD2.n69 VDD2.n68 12.0247
R1456 VDD2.n78 VDD2.n0 12.0247
R1457 VDD2.n148 VDD2.n89 11.249
R1458 VDD2.n119 VDD2.n106 11.249
R1459 VDD2.n35 VDD2.n22 11.249
R1460 VDD2.n64 VDD2.n6 11.249
R1461 VDD2.n147 VDD2.n92 10.4732
R1462 VDD2.n120 VDD2.n104 10.4732
R1463 VDD2.n36 VDD2.n20 10.4732
R1464 VDD2.n63 VDD2.n8 10.4732
R1465 VDD2.n144 VDD2.n143 9.69747
R1466 VDD2.n124 VDD2.n123 9.69747
R1467 VDD2.n40 VDD2.n39 9.69747
R1468 VDD2.n60 VDD2.n59 9.69747
R1469 VDD2.n163 VDD2.n162 9.45567
R1470 VDD2.n80 VDD2.n79 9.45567
R1471 VDD2.n137 VDD2.n136 9.3005
R1472 VDD2.n139 VDD2.n138 9.3005
R1473 VDD2.n94 VDD2.n93 9.3005
R1474 VDD2.n145 VDD2.n144 9.3005
R1475 VDD2.n147 VDD2.n146 9.3005
R1476 VDD2.n89 VDD2.n88 9.3005
R1477 VDD2.n153 VDD2.n152 9.3005
R1478 VDD2.n155 VDD2.n154 9.3005
R1479 VDD2.n162 VDD2.n161 9.3005
R1480 VDD2.n85 VDD2.n84 9.3005
R1481 VDD2.n98 VDD2.n97 9.3005
R1482 VDD2.n131 VDD2.n130 9.3005
R1483 VDD2.n129 VDD2.n128 9.3005
R1484 VDD2.n102 VDD2.n101 9.3005
R1485 VDD2.n123 VDD2.n122 9.3005
R1486 VDD2.n121 VDD2.n120 9.3005
R1487 VDD2.n106 VDD2.n105 9.3005
R1488 VDD2.n115 VDD2.n114 9.3005
R1489 VDD2.n113 VDD2.n112 9.3005
R1490 VDD2.n79 VDD2.n78 9.3005
R1491 VDD2.n2 VDD2.n1 9.3005
R1492 VDD2.n47 VDD2.n46 9.3005
R1493 VDD2.n45 VDD2.n44 9.3005
R1494 VDD2.n18 VDD2.n17 9.3005
R1495 VDD2.n39 VDD2.n38 9.3005
R1496 VDD2.n37 VDD2.n36 9.3005
R1497 VDD2.n22 VDD2.n21 9.3005
R1498 VDD2.n31 VDD2.n30 9.3005
R1499 VDD2.n29 VDD2.n28 9.3005
R1500 VDD2.n14 VDD2.n13 9.3005
R1501 VDD2.n53 VDD2.n52 9.3005
R1502 VDD2.n55 VDD2.n54 9.3005
R1503 VDD2.n10 VDD2.n9 9.3005
R1504 VDD2.n61 VDD2.n60 9.3005
R1505 VDD2.n63 VDD2.n62 9.3005
R1506 VDD2.n6 VDD2.n5 9.3005
R1507 VDD2.n70 VDD2.n69 9.3005
R1508 VDD2.n72 VDD2.n71 9.3005
R1509 VDD2.n140 VDD2.n94 8.92171
R1510 VDD2.n127 VDD2.n102 8.92171
R1511 VDD2.n43 VDD2.n18 8.92171
R1512 VDD2.n56 VDD2.n10 8.92171
R1513 VDD2.n139 VDD2.n96 8.14595
R1514 VDD2.n128 VDD2.n100 8.14595
R1515 VDD2.n44 VDD2.n16 8.14595
R1516 VDD2.n55 VDD2.n12 8.14595
R1517 VDD2.n136 VDD2.n135 7.3702
R1518 VDD2.n132 VDD2.n131 7.3702
R1519 VDD2.n48 VDD2.n47 7.3702
R1520 VDD2.n52 VDD2.n51 7.3702
R1521 VDD2.n135 VDD2.n98 6.59444
R1522 VDD2.n132 VDD2.n98 6.59444
R1523 VDD2.n48 VDD2.n14 6.59444
R1524 VDD2.n51 VDD2.n14 6.59444
R1525 VDD2.n136 VDD2.n96 5.81868
R1526 VDD2.n131 VDD2.n100 5.81868
R1527 VDD2.n47 VDD2.n16 5.81868
R1528 VDD2.n52 VDD2.n12 5.81868
R1529 VDD2.n140 VDD2.n139 5.04292
R1530 VDD2.n128 VDD2.n127 5.04292
R1531 VDD2.n44 VDD2.n43 5.04292
R1532 VDD2.n56 VDD2.n55 5.04292
R1533 VDD2.n143 VDD2.n94 4.26717
R1534 VDD2.n124 VDD2.n102 4.26717
R1535 VDD2.n40 VDD2.n18 4.26717
R1536 VDD2.n59 VDD2.n10 4.26717
R1537 VDD2.n113 VDD2.n109 3.70982
R1538 VDD2.n29 VDD2.n25 3.70982
R1539 VDD2.n144 VDD2.n92 3.49141
R1540 VDD2.n123 VDD2.n104 3.49141
R1541 VDD2.n39 VDD2.n20 3.49141
R1542 VDD2.n60 VDD2.n8 3.49141
R1543 VDD2.n148 VDD2.n147 2.71565
R1544 VDD2.n120 VDD2.n119 2.71565
R1545 VDD2.n36 VDD2.n35 2.71565
R1546 VDD2.n64 VDD2.n63 2.71565
R1547 VDD2 VDD2.n164 2.4574
R1548 VDD2.n165 VDD2.t1 2.21625
R1549 VDD2.n165 VDD2.t5 2.21625
R1550 VDD2.n81 VDD2.t2 2.21625
R1551 VDD2.n81 VDD2.t0 2.21625
R1552 VDD2.n163 VDD2.n83 1.93989
R1553 VDD2.n151 VDD2.n89 1.93989
R1554 VDD2.n116 VDD2.n106 1.93989
R1555 VDD2.n32 VDD2.n22 1.93989
R1556 VDD2.n68 VDD2.n6 1.93989
R1557 VDD2.n80 VDD2.n0 1.93989
R1558 VDD2.n161 VDD2.n160 1.16414
R1559 VDD2.n152 VDD2.n87 1.16414
R1560 VDD2.n115 VDD2.n108 1.16414
R1561 VDD2.n31 VDD2.n24 1.16414
R1562 VDD2.n69 VDD2.n4 1.16414
R1563 VDD2.n78 VDD2.n77 1.16414
R1564 VDD2.n157 VDD2.n85 0.388379
R1565 VDD2.n156 VDD2.n155 0.388379
R1566 VDD2.n112 VDD2.n111 0.388379
R1567 VDD2.n28 VDD2.n27 0.388379
R1568 VDD2.n73 VDD2.n72 0.388379
R1569 VDD2.n74 VDD2.n2 0.388379
R1570 VDD2.n162 VDD2.n84 0.155672
R1571 VDD2.n154 VDD2.n84 0.155672
R1572 VDD2.n154 VDD2.n153 0.155672
R1573 VDD2.n153 VDD2.n88 0.155672
R1574 VDD2.n146 VDD2.n88 0.155672
R1575 VDD2.n146 VDD2.n145 0.155672
R1576 VDD2.n145 VDD2.n93 0.155672
R1577 VDD2.n138 VDD2.n93 0.155672
R1578 VDD2.n138 VDD2.n137 0.155672
R1579 VDD2.n137 VDD2.n97 0.155672
R1580 VDD2.n130 VDD2.n97 0.155672
R1581 VDD2.n130 VDD2.n129 0.155672
R1582 VDD2.n129 VDD2.n101 0.155672
R1583 VDD2.n122 VDD2.n101 0.155672
R1584 VDD2.n122 VDD2.n121 0.155672
R1585 VDD2.n121 VDD2.n105 0.155672
R1586 VDD2.n114 VDD2.n105 0.155672
R1587 VDD2.n114 VDD2.n113 0.155672
R1588 VDD2.n30 VDD2.n29 0.155672
R1589 VDD2.n30 VDD2.n21 0.155672
R1590 VDD2.n37 VDD2.n21 0.155672
R1591 VDD2.n38 VDD2.n37 0.155672
R1592 VDD2.n38 VDD2.n17 0.155672
R1593 VDD2.n45 VDD2.n17 0.155672
R1594 VDD2.n46 VDD2.n45 0.155672
R1595 VDD2.n46 VDD2.n13 0.155672
R1596 VDD2.n53 VDD2.n13 0.155672
R1597 VDD2.n54 VDD2.n53 0.155672
R1598 VDD2.n54 VDD2.n9 0.155672
R1599 VDD2.n61 VDD2.n9 0.155672
R1600 VDD2.n62 VDD2.n61 0.155672
R1601 VDD2.n62 VDD2.n5 0.155672
R1602 VDD2.n70 VDD2.n5 0.155672
R1603 VDD2.n71 VDD2.n70 0.155672
R1604 VDD2.n71 VDD2.n1 0.155672
R1605 VDD2.n79 VDD2.n1 0.155672
R1606 VTAIL.n330 VTAIL.n254 756.745
R1607 VTAIL.n78 VTAIL.n2 756.745
R1608 VTAIL.n248 VTAIL.n172 756.745
R1609 VTAIL.n164 VTAIL.n88 756.745
R1610 VTAIL.n281 VTAIL.n280 585
R1611 VTAIL.n278 VTAIL.n277 585
R1612 VTAIL.n287 VTAIL.n286 585
R1613 VTAIL.n289 VTAIL.n288 585
R1614 VTAIL.n274 VTAIL.n273 585
R1615 VTAIL.n295 VTAIL.n294 585
R1616 VTAIL.n297 VTAIL.n296 585
R1617 VTAIL.n270 VTAIL.n269 585
R1618 VTAIL.n303 VTAIL.n302 585
R1619 VTAIL.n305 VTAIL.n304 585
R1620 VTAIL.n266 VTAIL.n265 585
R1621 VTAIL.n311 VTAIL.n310 585
R1622 VTAIL.n313 VTAIL.n312 585
R1623 VTAIL.n262 VTAIL.n261 585
R1624 VTAIL.n319 VTAIL.n318 585
R1625 VTAIL.n322 VTAIL.n321 585
R1626 VTAIL.n320 VTAIL.n258 585
R1627 VTAIL.n327 VTAIL.n257 585
R1628 VTAIL.n329 VTAIL.n328 585
R1629 VTAIL.n331 VTAIL.n330 585
R1630 VTAIL.n29 VTAIL.n28 585
R1631 VTAIL.n26 VTAIL.n25 585
R1632 VTAIL.n35 VTAIL.n34 585
R1633 VTAIL.n37 VTAIL.n36 585
R1634 VTAIL.n22 VTAIL.n21 585
R1635 VTAIL.n43 VTAIL.n42 585
R1636 VTAIL.n45 VTAIL.n44 585
R1637 VTAIL.n18 VTAIL.n17 585
R1638 VTAIL.n51 VTAIL.n50 585
R1639 VTAIL.n53 VTAIL.n52 585
R1640 VTAIL.n14 VTAIL.n13 585
R1641 VTAIL.n59 VTAIL.n58 585
R1642 VTAIL.n61 VTAIL.n60 585
R1643 VTAIL.n10 VTAIL.n9 585
R1644 VTAIL.n67 VTAIL.n66 585
R1645 VTAIL.n70 VTAIL.n69 585
R1646 VTAIL.n68 VTAIL.n6 585
R1647 VTAIL.n75 VTAIL.n5 585
R1648 VTAIL.n77 VTAIL.n76 585
R1649 VTAIL.n79 VTAIL.n78 585
R1650 VTAIL.n249 VTAIL.n248 585
R1651 VTAIL.n247 VTAIL.n246 585
R1652 VTAIL.n245 VTAIL.n175 585
R1653 VTAIL.n179 VTAIL.n176 585
R1654 VTAIL.n240 VTAIL.n239 585
R1655 VTAIL.n238 VTAIL.n237 585
R1656 VTAIL.n181 VTAIL.n180 585
R1657 VTAIL.n232 VTAIL.n231 585
R1658 VTAIL.n230 VTAIL.n229 585
R1659 VTAIL.n185 VTAIL.n184 585
R1660 VTAIL.n224 VTAIL.n223 585
R1661 VTAIL.n222 VTAIL.n221 585
R1662 VTAIL.n189 VTAIL.n188 585
R1663 VTAIL.n216 VTAIL.n215 585
R1664 VTAIL.n214 VTAIL.n213 585
R1665 VTAIL.n193 VTAIL.n192 585
R1666 VTAIL.n208 VTAIL.n207 585
R1667 VTAIL.n206 VTAIL.n205 585
R1668 VTAIL.n197 VTAIL.n196 585
R1669 VTAIL.n200 VTAIL.n199 585
R1670 VTAIL.n165 VTAIL.n164 585
R1671 VTAIL.n163 VTAIL.n162 585
R1672 VTAIL.n161 VTAIL.n91 585
R1673 VTAIL.n95 VTAIL.n92 585
R1674 VTAIL.n156 VTAIL.n155 585
R1675 VTAIL.n154 VTAIL.n153 585
R1676 VTAIL.n97 VTAIL.n96 585
R1677 VTAIL.n148 VTAIL.n147 585
R1678 VTAIL.n146 VTAIL.n145 585
R1679 VTAIL.n101 VTAIL.n100 585
R1680 VTAIL.n140 VTAIL.n139 585
R1681 VTAIL.n138 VTAIL.n137 585
R1682 VTAIL.n105 VTAIL.n104 585
R1683 VTAIL.n132 VTAIL.n131 585
R1684 VTAIL.n130 VTAIL.n129 585
R1685 VTAIL.n109 VTAIL.n108 585
R1686 VTAIL.n124 VTAIL.n123 585
R1687 VTAIL.n122 VTAIL.n121 585
R1688 VTAIL.n113 VTAIL.n112 585
R1689 VTAIL.n116 VTAIL.n115 585
R1690 VTAIL.t1 VTAIL.n198 327.466
R1691 VTAIL.t8 VTAIL.n114 327.466
R1692 VTAIL.t6 VTAIL.n279 327.466
R1693 VTAIL.t0 VTAIL.n27 327.466
R1694 VTAIL.n280 VTAIL.n277 171.744
R1695 VTAIL.n287 VTAIL.n277 171.744
R1696 VTAIL.n288 VTAIL.n287 171.744
R1697 VTAIL.n288 VTAIL.n273 171.744
R1698 VTAIL.n295 VTAIL.n273 171.744
R1699 VTAIL.n296 VTAIL.n295 171.744
R1700 VTAIL.n296 VTAIL.n269 171.744
R1701 VTAIL.n303 VTAIL.n269 171.744
R1702 VTAIL.n304 VTAIL.n303 171.744
R1703 VTAIL.n304 VTAIL.n265 171.744
R1704 VTAIL.n311 VTAIL.n265 171.744
R1705 VTAIL.n312 VTAIL.n311 171.744
R1706 VTAIL.n312 VTAIL.n261 171.744
R1707 VTAIL.n319 VTAIL.n261 171.744
R1708 VTAIL.n321 VTAIL.n319 171.744
R1709 VTAIL.n321 VTAIL.n320 171.744
R1710 VTAIL.n320 VTAIL.n257 171.744
R1711 VTAIL.n329 VTAIL.n257 171.744
R1712 VTAIL.n330 VTAIL.n329 171.744
R1713 VTAIL.n28 VTAIL.n25 171.744
R1714 VTAIL.n35 VTAIL.n25 171.744
R1715 VTAIL.n36 VTAIL.n35 171.744
R1716 VTAIL.n36 VTAIL.n21 171.744
R1717 VTAIL.n43 VTAIL.n21 171.744
R1718 VTAIL.n44 VTAIL.n43 171.744
R1719 VTAIL.n44 VTAIL.n17 171.744
R1720 VTAIL.n51 VTAIL.n17 171.744
R1721 VTAIL.n52 VTAIL.n51 171.744
R1722 VTAIL.n52 VTAIL.n13 171.744
R1723 VTAIL.n59 VTAIL.n13 171.744
R1724 VTAIL.n60 VTAIL.n59 171.744
R1725 VTAIL.n60 VTAIL.n9 171.744
R1726 VTAIL.n67 VTAIL.n9 171.744
R1727 VTAIL.n69 VTAIL.n67 171.744
R1728 VTAIL.n69 VTAIL.n68 171.744
R1729 VTAIL.n68 VTAIL.n5 171.744
R1730 VTAIL.n77 VTAIL.n5 171.744
R1731 VTAIL.n78 VTAIL.n77 171.744
R1732 VTAIL.n248 VTAIL.n247 171.744
R1733 VTAIL.n247 VTAIL.n175 171.744
R1734 VTAIL.n179 VTAIL.n175 171.744
R1735 VTAIL.n239 VTAIL.n179 171.744
R1736 VTAIL.n239 VTAIL.n238 171.744
R1737 VTAIL.n238 VTAIL.n180 171.744
R1738 VTAIL.n231 VTAIL.n180 171.744
R1739 VTAIL.n231 VTAIL.n230 171.744
R1740 VTAIL.n230 VTAIL.n184 171.744
R1741 VTAIL.n223 VTAIL.n184 171.744
R1742 VTAIL.n223 VTAIL.n222 171.744
R1743 VTAIL.n222 VTAIL.n188 171.744
R1744 VTAIL.n215 VTAIL.n188 171.744
R1745 VTAIL.n215 VTAIL.n214 171.744
R1746 VTAIL.n214 VTAIL.n192 171.744
R1747 VTAIL.n207 VTAIL.n192 171.744
R1748 VTAIL.n207 VTAIL.n206 171.744
R1749 VTAIL.n206 VTAIL.n196 171.744
R1750 VTAIL.n199 VTAIL.n196 171.744
R1751 VTAIL.n164 VTAIL.n163 171.744
R1752 VTAIL.n163 VTAIL.n91 171.744
R1753 VTAIL.n95 VTAIL.n91 171.744
R1754 VTAIL.n155 VTAIL.n95 171.744
R1755 VTAIL.n155 VTAIL.n154 171.744
R1756 VTAIL.n154 VTAIL.n96 171.744
R1757 VTAIL.n147 VTAIL.n96 171.744
R1758 VTAIL.n147 VTAIL.n146 171.744
R1759 VTAIL.n146 VTAIL.n100 171.744
R1760 VTAIL.n139 VTAIL.n100 171.744
R1761 VTAIL.n139 VTAIL.n138 171.744
R1762 VTAIL.n138 VTAIL.n104 171.744
R1763 VTAIL.n131 VTAIL.n104 171.744
R1764 VTAIL.n131 VTAIL.n130 171.744
R1765 VTAIL.n130 VTAIL.n108 171.744
R1766 VTAIL.n123 VTAIL.n108 171.744
R1767 VTAIL.n123 VTAIL.n122 171.744
R1768 VTAIL.n122 VTAIL.n112 171.744
R1769 VTAIL.n115 VTAIL.n112 171.744
R1770 VTAIL.n280 VTAIL.t6 85.8723
R1771 VTAIL.n28 VTAIL.t0 85.8723
R1772 VTAIL.n199 VTAIL.t1 85.8723
R1773 VTAIL.n115 VTAIL.t8 85.8723
R1774 VTAIL.n171 VTAIL.n170 54.6696
R1775 VTAIL.n87 VTAIL.n86 54.6696
R1776 VTAIL.n1 VTAIL.n0 54.6694
R1777 VTAIL.n85 VTAIL.n84 54.6694
R1778 VTAIL.n335 VTAIL.n334 32.7672
R1779 VTAIL.n83 VTAIL.n82 32.7672
R1780 VTAIL.n253 VTAIL.n252 32.7672
R1781 VTAIL.n169 VTAIL.n168 32.7672
R1782 VTAIL.n87 VTAIL.n85 31.41
R1783 VTAIL.n335 VTAIL.n253 28.2117
R1784 VTAIL.n281 VTAIL.n279 16.3895
R1785 VTAIL.n29 VTAIL.n27 16.3895
R1786 VTAIL.n200 VTAIL.n198 16.3895
R1787 VTAIL.n116 VTAIL.n114 16.3895
R1788 VTAIL.n328 VTAIL.n327 13.1884
R1789 VTAIL.n76 VTAIL.n75 13.1884
R1790 VTAIL.n246 VTAIL.n245 13.1884
R1791 VTAIL.n162 VTAIL.n161 13.1884
R1792 VTAIL.n282 VTAIL.n278 12.8005
R1793 VTAIL.n326 VTAIL.n258 12.8005
R1794 VTAIL.n331 VTAIL.n256 12.8005
R1795 VTAIL.n30 VTAIL.n26 12.8005
R1796 VTAIL.n74 VTAIL.n6 12.8005
R1797 VTAIL.n79 VTAIL.n4 12.8005
R1798 VTAIL.n249 VTAIL.n174 12.8005
R1799 VTAIL.n244 VTAIL.n176 12.8005
R1800 VTAIL.n201 VTAIL.n197 12.8005
R1801 VTAIL.n165 VTAIL.n90 12.8005
R1802 VTAIL.n160 VTAIL.n92 12.8005
R1803 VTAIL.n117 VTAIL.n113 12.8005
R1804 VTAIL.n286 VTAIL.n285 12.0247
R1805 VTAIL.n323 VTAIL.n322 12.0247
R1806 VTAIL.n332 VTAIL.n254 12.0247
R1807 VTAIL.n34 VTAIL.n33 12.0247
R1808 VTAIL.n71 VTAIL.n70 12.0247
R1809 VTAIL.n80 VTAIL.n2 12.0247
R1810 VTAIL.n250 VTAIL.n172 12.0247
R1811 VTAIL.n241 VTAIL.n240 12.0247
R1812 VTAIL.n205 VTAIL.n204 12.0247
R1813 VTAIL.n166 VTAIL.n88 12.0247
R1814 VTAIL.n157 VTAIL.n156 12.0247
R1815 VTAIL.n121 VTAIL.n120 12.0247
R1816 VTAIL.n289 VTAIL.n276 11.249
R1817 VTAIL.n318 VTAIL.n260 11.249
R1818 VTAIL.n37 VTAIL.n24 11.249
R1819 VTAIL.n66 VTAIL.n8 11.249
R1820 VTAIL.n237 VTAIL.n178 11.249
R1821 VTAIL.n208 VTAIL.n195 11.249
R1822 VTAIL.n153 VTAIL.n94 11.249
R1823 VTAIL.n124 VTAIL.n111 11.249
R1824 VTAIL.n290 VTAIL.n274 10.4732
R1825 VTAIL.n317 VTAIL.n262 10.4732
R1826 VTAIL.n38 VTAIL.n22 10.4732
R1827 VTAIL.n65 VTAIL.n10 10.4732
R1828 VTAIL.n236 VTAIL.n181 10.4732
R1829 VTAIL.n209 VTAIL.n193 10.4732
R1830 VTAIL.n152 VTAIL.n97 10.4732
R1831 VTAIL.n125 VTAIL.n109 10.4732
R1832 VTAIL.n294 VTAIL.n293 9.69747
R1833 VTAIL.n314 VTAIL.n313 9.69747
R1834 VTAIL.n42 VTAIL.n41 9.69747
R1835 VTAIL.n62 VTAIL.n61 9.69747
R1836 VTAIL.n233 VTAIL.n232 9.69747
R1837 VTAIL.n213 VTAIL.n212 9.69747
R1838 VTAIL.n149 VTAIL.n148 9.69747
R1839 VTAIL.n129 VTAIL.n128 9.69747
R1840 VTAIL.n334 VTAIL.n333 9.45567
R1841 VTAIL.n82 VTAIL.n81 9.45567
R1842 VTAIL.n252 VTAIL.n251 9.45567
R1843 VTAIL.n168 VTAIL.n167 9.45567
R1844 VTAIL.n333 VTAIL.n332 9.3005
R1845 VTAIL.n256 VTAIL.n255 9.3005
R1846 VTAIL.n301 VTAIL.n300 9.3005
R1847 VTAIL.n299 VTAIL.n298 9.3005
R1848 VTAIL.n272 VTAIL.n271 9.3005
R1849 VTAIL.n293 VTAIL.n292 9.3005
R1850 VTAIL.n291 VTAIL.n290 9.3005
R1851 VTAIL.n276 VTAIL.n275 9.3005
R1852 VTAIL.n285 VTAIL.n284 9.3005
R1853 VTAIL.n283 VTAIL.n282 9.3005
R1854 VTAIL.n268 VTAIL.n267 9.3005
R1855 VTAIL.n307 VTAIL.n306 9.3005
R1856 VTAIL.n309 VTAIL.n308 9.3005
R1857 VTAIL.n264 VTAIL.n263 9.3005
R1858 VTAIL.n315 VTAIL.n314 9.3005
R1859 VTAIL.n317 VTAIL.n316 9.3005
R1860 VTAIL.n260 VTAIL.n259 9.3005
R1861 VTAIL.n324 VTAIL.n323 9.3005
R1862 VTAIL.n326 VTAIL.n325 9.3005
R1863 VTAIL.n81 VTAIL.n80 9.3005
R1864 VTAIL.n4 VTAIL.n3 9.3005
R1865 VTAIL.n49 VTAIL.n48 9.3005
R1866 VTAIL.n47 VTAIL.n46 9.3005
R1867 VTAIL.n20 VTAIL.n19 9.3005
R1868 VTAIL.n41 VTAIL.n40 9.3005
R1869 VTAIL.n39 VTAIL.n38 9.3005
R1870 VTAIL.n24 VTAIL.n23 9.3005
R1871 VTAIL.n33 VTAIL.n32 9.3005
R1872 VTAIL.n31 VTAIL.n30 9.3005
R1873 VTAIL.n16 VTAIL.n15 9.3005
R1874 VTAIL.n55 VTAIL.n54 9.3005
R1875 VTAIL.n57 VTAIL.n56 9.3005
R1876 VTAIL.n12 VTAIL.n11 9.3005
R1877 VTAIL.n63 VTAIL.n62 9.3005
R1878 VTAIL.n65 VTAIL.n64 9.3005
R1879 VTAIL.n8 VTAIL.n7 9.3005
R1880 VTAIL.n72 VTAIL.n71 9.3005
R1881 VTAIL.n74 VTAIL.n73 9.3005
R1882 VTAIL.n226 VTAIL.n225 9.3005
R1883 VTAIL.n228 VTAIL.n227 9.3005
R1884 VTAIL.n183 VTAIL.n182 9.3005
R1885 VTAIL.n234 VTAIL.n233 9.3005
R1886 VTAIL.n236 VTAIL.n235 9.3005
R1887 VTAIL.n178 VTAIL.n177 9.3005
R1888 VTAIL.n242 VTAIL.n241 9.3005
R1889 VTAIL.n244 VTAIL.n243 9.3005
R1890 VTAIL.n251 VTAIL.n250 9.3005
R1891 VTAIL.n174 VTAIL.n173 9.3005
R1892 VTAIL.n187 VTAIL.n186 9.3005
R1893 VTAIL.n220 VTAIL.n219 9.3005
R1894 VTAIL.n218 VTAIL.n217 9.3005
R1895 VTAIL.n191 VTAIL.n190 9.3005
R1896 VTAIL.n212 VTAIL.n211 9.3005
R1897 VTAIL.n210 VTAIL.n209 9.3005
R1898 VTAIL.n195 VTAIL.n194 9.3005
R1899 VTAIL.n204 VTAIL.n203 9.3005
R1900 VTAIL.n202 VTAIL.n201 9.3005
R1901 VTAIL.n142 VTAIL.n141 9.3005
R1902 VTAIL.n144 VTAIL.n143 9.3005
R1903 VTAIL.n99 VTAIL.n98 9.3005
R1904 VTAIL.n150 VTAIL.n149 9.3005
R1905 VTAIL.n152 VTAIL.n151 9.3005
R1906 VTAIL.n94 VTAIL.n93 9.3005
R1907 VTAIL.n158 VTAIL.n157 9.3005
R1908 VTAIL.n160 VTAIL.n159 9.3005
R1909 VTAIL.n167 VTAIL.n166 9.3005
R1910 VTAIL.n90 VTAIL.n89 9.3005
R1911 VTAIL.n103 VTAIL.n102 9.3005
R1912 VTAIL.n136 VTAIL.n135 9.3005
R1913 VTAIL.n134 VTAIL.n133 9.3005
R1914 VTAIL.n107 VTAIL.n106 9.3005
R1915 VTAIL.n128 VTAIL.n127 9.3005
R1916 VTAIL.n126 VTAIL.n125 9.3005
R1917 VTAIL.n111 VTAIL.n110 9.3005
R1918 VTAIL.n120 VTAIL.n119 9.3005
R1919 VTAIL.n118 VTAIL.n117 9.3005
R1920 VTAIL.n297 VTAIL.n272 8.92171
R1921 VTAIL.n310 VTAIL.n264 8.92171
R1922 VTAIL.n45 VTAIL.n20 8.92171
R1923 VTAIL.n58 VTAIL.n12 8.92171
R1924 VTAIL.n229 VTAIL.n183 8.92171
R1925 VTAIL.n216 VTAIL.n191 8.92171
R1926 VTAIL.n145 VTAIL.n99 8.92171
R1927 VTAIL.n132 VTAIL.n107 8.92171
R1928 VTAIL.n298 VTAIL.n270 8.14595
R1929 VTAIL.n309 VTAIL.n266 8.14595
R1930 VTAIL.n46 VTAIL.n18 8.14595
R1931 VTAIL.n57 VTAIL.n14 8.14595
R1932 VTAIL.n228 VTAIL.n185 8.14595
R1933 VTAIL.n217 VTAIL.n189 8.14595
R1934 VTAIL.n144 VTAIL.n101 8.14595
R1935 VTAIL.n133 VTAIL.n105 8.14595
R1936 VTAIL.n302 VTAIL.n301 7.3702
R1937 VTAIL.n306 VTAIL.n305 7.3702
R1938 VTAIL.n50 VTAIL.n49 7.3702
R1939 VTAIL.n54 VTAIL.n53 7.3702
R1940 VTAIL.n225 VTAIL.n224 7.3702
R1941 VTAIL.n221 VTAIL.n220 7.3702
R1942 VTAIL.n141 VTAIL.n140 7.3702
R1943 VTAIL.n137 VTAIL.n136 7.3702
R1944 VTAIL.n302 VTAIL.n268 6.59444
R1945 VTAIL.n305 VTAIL.n268 6.59444
R1946 VTAIL.n50 VTAIL.n16 6.59444
R1947 VTAIL.n53 VTAIL.n16 6.59444
R1948 VTAIL.n224 VTAIL.n187 6.59444
R1949 VTAIL.n221 VTAIL.n187 6.59444
R1950 VTAIL.n140 VTAIL.n103 6.59444
R1951 VTAIL.n137 VTAIL.n103 6.59444
R1952 VTAIL.n301 VTAIL.n270 5.81868
R1953 VTAIL.n306 VTAIL.n266 5.81868
R1954 VTAIL.n49 VTAIL.n18 5.81868
R1955 VTAIL.n54 VTAIL.n14 5.81868
R1956 VTAIL.n225 VTAIL.n185 5.81868
R1957 VTAIL.n220 VTAIL.n189 5.81868
R1958 VTAIL.n141 VTAIL.n101 5.81868
R1959 VTAIL.n136 VTAIL.n105 5.81868
R1960 VTAIL.n298 VTAIL.n297 5.04292
R1961 VTAIL.n310 VTAIL.n309 5.04292
R1962 VTAIL.n46 VTAIL.n45 5.04292
R1963 VTAIL.n58 VTAIL.n57 5.04292
R1964 VTAIL.n229 VTAIL.n228 5.04292
R1965 VTAIL.n217 VTAIL.n216 5.04292
R1966 VTAIL.n145 VTAIL.n144 5.04292
R1967 VTAIL.n133 VTAIL.n132 5.04292
R1968 VTAIL.n294 VTAIL.n272 4.26717
R1969 VTAIL.n313 VTAIL.n264 4.26717
R1970 VTAIL.n42 VTAIL.n20 4.26717
R1971 VTAIL.n61 VTAIL.n12 4.26717
R1972 VTAIL.n232 VTAIL.n183 4.26717
R1973 VTAIL.n213 VTAIL.n191 4.26717
R1974 VTAIL.n148 VTAIL.n99 4.26717
R1975 VTAIL.n129 VTAIL.n107 4.26717
R1976 VTAIL.n283 VTAIL.n279 3.70982
R1977 VTAIL.n31 VTAIL.n27 3.70982
R1978 VTAIL.n202 VTAIL.n198 3.70982
R1979 VTAIL.n118 VTAIL.n114 3.70982
R1980 VTAIL.n293 VTAIL.n274 3.49141
R1981 VTAIL.n314 VTAIL.n262 3.49141
R1982 VTAIL.n41 VTAIL.n22 3.49141
R1983 VTAIL.n62 VTAIL.n10 3.49141
R1984 VTAIL.n233 VTAIL.n181 3.49141
R1985 VTAIL.n212 VTAIL.n193 3.49141
R1986 VTAIL.n149 VTAIL.n97 3.49141
R1987 VTAIL.n128 VTAIL.n109 3.49141
R1988 VTAIL.n169 VTAIL.n87 3.19878
R1989 VTAIL.n253 VTAIL.n171 3.19878
R1990 VTAIL.n85 VTAIL.n83 3.19878
R1991 VTAIL.n290 VTAIL.n289 2.71565
R1992 VTAIL.n318 VTAIL.n317 2.71565
R1993 VTAIL.n38 VTAIL.n37 2.71565
R1994 VTAIL.n66 VTAIL.n65 2.71565
R1995 VTAIL.n237 VTAIL.n236 2.71565
R1996 VTAIL.n209 VTAIL.n208 2.71565
R1997 VTAIL.n153 VTAIL.n152 2.71565
R1998 VTAIL.n125 VTAIL.n124 2.71565
R1999 VTAIL VTAIL.n335 2.34102
R2000 VTAIL.n0 VTAIL.t9 2.21625
R2001 VTAIL.n0 VTAIL.t11 2.21625
R2002 VTAIL.n84 VTAIL.t2 2.21625
R2003 VTAIL.n84 VTAIL.t5 2.21625
R2004 VTAIL.n170 VTAIL.t3 2.21625
R2005 VTAIL.n170 VTAIL.t4 2.21625
R2006 VTAIL.n86 VTAIL.t10 2.21625
R2007 VTAIL.n86 VTAIL.t7 2.21625
R2008 VTAIL.n171 VTAIL.n169 2.06947
R2009 VTAIL.n83 VTAIL.n1 2.06947
R2010 VTAIL.n286 VTAIL.n276 1.93989
R2011 VTAIL.n322 VTAIL.n260 1.93989
R2012 VTAIL.n334 VTAIL.n254 1.93989
R2013 VTAIL.n34 VTAIL.n24 1.93989
R2014 VTAIL.n70 VTAIL.n8 1.93989
R2015 VTAIL.n82 VTAIL.n2 1.93989
R2016 VTAIL.n252 VTAIL.n172 1.93989
R2017 VTAIL.n240 VTAIL.n178 1.93989
R2018 VTAIL.n205 VTAIL.n195 1.93989
R2019 VTAIL.n168 VTAIL.n88 1.93989
R2020 VTAIL.n156 VTAIL.n94 1.93989
R2021 VTAIL.n121 VTAIL.n111 1.93989
R2022 VTAIL.n285 VTAIL.n278 1.16414
R2023 VTAIL.n323 VTAIL.n258 1.16414
R2024 VTAIL.n332 VTAIL.n331 1.16414
R2025 VTAIL.n33 VTAIL.n26 1.16414
R2026 VTAIL.n71 VTAIL.n6 1.16414
R2027 VTAIL.n80 VTAIL.n79 1.16414
R2028 VTAIL.n250 VTAIL.n249 1.16414
R2029 VTAIL.n241 VTAIL.n176 1.16414
R2030 VTAIL.n204 VTAIL.n197 1.16414
R2031 VTAIL.n166 VTAIL.n165 1.16414
R2032 VTAIL.n157 VTAIL.n92 1.16414
R2033 VTAIL.n120 VTAIL.n113 1.16414
R2034 VTAIL VTAIL.n1 0.858259
R2035 VTAIL.n282 VTAIL.n281 0.388379
R2036 VTAIL.n327 VTAIL.n326 0.388379
R2037 VTAIL.n328 VTAIL.n256 0.388379
R2038 VTAIL.n30 VTAIL.n29 0.388379
R2039 VTAIL.n75 VTAIL.n74 0.388379
R2040 VTAIL.n76 VTAIL.n4 0.388379
R2041 VTAIL.n246 VTAIL.n174 0.388379
R2042 VTAIL.n245 VTAIL.n244 0.388379
R2043 VTAIL.n201 VTAIL.n200 0.388379
R2044 VTAIL.n162 VTAIL.n90 0.388379
R2045 VTAIL.n161 VTAIL.n160 0.388379
R2046 VTAIL.n117 VTAIL.n116 0.388379
R2047 VTAIL.n284 VTAIL.n283 0.155672
R2048 VTAIL.n284 VTAIL.n275 0.155672
R2049 VTAIL.n291 VTAIL.n275 0.155672
R2050 VTAIL.n292 VTAIL.n291 0.155672
R2051 VTAIL.n292 VTAIL.n271 0.155672
R2052 VTAIL.n299 VTAIL.n271 0.155672
R2053 VTAIL.n300 VTAIL.n299 0.155672
R2054 VTAIL.n300 VTAIL.n267 0.155672
R2055 VTAIL.n307 VTAIL.n267 0.155672
R2056 VTAIL.n308 VTAIL.n307 0.155672
R2057 VTAIL.n308 VTAIL.n263 0.155672
R2058 VTAIL.n315 VTAIL.n263 0.155672
R2059 VTAIL.n316 VTAIL.n315 0.155672
R2060 VTAIL.n316 VTAIL.n259 0.155672
R2061 VTAIL.n324 VTAIL.n259 0.155672
R2062 VTAIL.n325 VTAIL.n324 0.155672
R2063 VTAIL.n325 VTAIL.n255 0.155672
R2064 VTAIL.n333 VTAIL.n255 0.155672
R2065 VTAIL.n32 VTAIL.n31 0.155672
R2066 VTAIL.n32 VTAIL.n23 0.155672
R2067 VTAIL.n39 VTAIL.n23 0.155672
R2068 VTAIL.n40 VTAIL.n39 0.155672
R2069 VTAIL.n40 VTAIL.n19 0.155672
R2070 VTAIL.n47 VTAIL.n19 0.155672
R2071 VTAIL.n48 VTAIL.n47 0.155672
R2072 VTAIL.n48 VTAIL.n15 0.155672
R2073 VTAIL.n55 VTAIL.n15 0.155672
R2074 VTAIL.n56 VTAIL.n55 0.155672
R2075 VTAIL.n56 VTAIL.n11 0.155672
R2076 VTAIL.n63 VTAIL.n11 0.155672
R2077 VTAIL.n64 VTAIL.n63 0.155672
R2078 VTAIL.n64 VTAIL.n7 0.155672
R2079 VTAIL.n72 VTAIL.n7 0.155672
R2080 VTAIL.n73 VTAIL.n72 0.155672
R2081 VTAIL.n73 VTAIL.n3 0.155672
R2082 VTAIL.n81 VTAIL.n3 0.155672
R2083 VTAIL.n251 VTAIL.n173 0.155672
R2084 VTAIL.n243 VTAIL.n173 0.155672
R2085 VTAIL.n243 VTAIL.n242 0.155672
R2086 VTAIL.n242 VTAIL.n177 0.155672
R2087 VTAIL.n235 VTAIL.n177 0.155672
R2088 VTAIL.n235 VTAIL.n234 0.155672
R2089 VTAIL.n234 VTAIL.n182 0.155672
R2090 VTAIL.n227 VTAIL.n182 0.155672
R2091 VTAIL.n227 VTAIL.n226 0.155672
R2092 VTAIL.n226 VTAIL.n186 0.155672
R2093 VTAIL.n219 VTAIL.n186 0.155672
R2094 VTAIL.n219 VTAIL.n218 0.155672
R2095 VTAIL.n218 VTAIL.n190 0.155672
R2096 VTAIL.n211 VTAIL.n190 0.155672
R2097 VTAIL.n211 VTAIL.n210 0.155672
R2098 VTAIL.n210 VTAIL.n194 0.155672
R2099 VTAIL.n203 VTAIL.n194 0.155672
R2100 VTAIL.n203 VTAIL.n202 0.155672
R2101 VTAIL.n167 VTAIL.n89 0.155672
R2102 VTAIL.n159 VTAIL.n89 0.155672
R2103 VTAIL.n159 VTAIL.n158 0.155672
R2104 VTAIL.n158 VTAIL.n93 0.155672
R2105 VTAIL.n151 VTAIL.n93 0.155672
R2106 VTAIL.n151 VTAIL.n150 0.155672
R2107 VTAIL.n150 VTAIL.n98 0.155672
R2108 VTAIL.n143 VTAIL.n98 0.155672
R2109 VTAIL.n143 VTAIL.n142 0.155672
R2110 VTAIL.n142 VTAIL.n102 0.155672
R2111 VTAIL.n135 VTAIL.n102 0.155672
R2112 VTAIL.n135 VTAIL.n134 0.155672
R2113 VTAIL.n134 VTAIL.n106 0.155672
R2114 VTAIL.n127 VTAIL.n106 0.155672
R2115 VTAIL.n127 VTAIL.n126 0.155672
R2116 VTAIL.n126 VTAIL.n110 0.155672
R2117 VTAIL.n119 VTAIL.n110 0.155672
R2118 VTAIL.n119 VTAIL.n118 0.155672
R2119 VP.n16 VP.n15 161.3
R2120 VP.n17 VP.n12 161.3
R2121 VP.n19 VP.n18 161.3
R2122 VP.n20 VP.n11 161.3
R2123 VP.n22 VP.n21 161.3
R2124 VP.n23 VP.n10 161.3
R2125 VP.n25 VP.n24 161.3
R2126 VP.n50 VP.n49 161.3
R2127 VP.n48 VP.n1 161.3
R2128 VP.n47 VP.n46 161.3
R2129 VP.n45 VP.n2 161.3
R2130 VP.n44 VP.n43 161.3
R2131 VP.n42 VP.n3 161.3
R2132 VP.n41 VP.n40 161.3
R2133 VP.n39 VP.n4 161.3
R2134 VP.n38 VP.n37 161.3
R2135 VP.n36 VP.n5 161.3
R2136 VP.n35 VP.n34 161.3
R2137 VP.n33 VP.n6 161.3
R2138 VP.n32 VP.n31 161.3
R2139 VP.n30 VP.n7 161.3
R2140 VP.n29 VP.n28 161.3
R2141 VP.n14 VP.t0 138.075
R2142 VP.n4 VP.t4 104.6
R2143 VP.n8 VP.t2 104.6
R2144 VP.n0 VP.t5 104.6
R2145 VP.n13 VP.t1 104.6
R2146 VP.n9 VP.t3 104.6
R2147 VP.n27 VP.n8 79.7913
R2148 VP.n51 VP.n0 79.7913
R2149 VP.n26 VP.n9 79.7913
R2150 VP.n35 VP.n6 54.5767
R2151 VP.n43 VP.n2 54.5767
R2152 VP.n18 VP.n11 54.5767
R2153 VP.n27 VP.n26 53.8213
R2154 VP.n14 VP.n13 50.1196
R2155 VP.n31 VP.n6 26.41
R2156 VP.n47 VP.n2 26.41
R2157 VP.n22 VP.n11 26.41
R2158 VP.n30 VP.n29 24.4675
R2159 VP.n31 VP.n30 24.4675
R2160 VP.n36 VP.n35 24.4675
R2161 VP.n37 VP.n36 24.4675
R2162 VP.n37 VP.n4 24.4675
R2163 VP.n41 VP.n4 24.4675
R2164 VP.n42 VP.n41 24.4675
R2165 VP.n43 VP.n42 24.4675
R2166 VP.n48 VP.n47 24.4675
R2167 VP.n49 VP.n48 24.4675
R2168 VP.n23 VP.n22 24.4675
R2169 VP.n24 VP.n23 24.4675
R2170 VP.n16 VP.n13 24.4675
R2171 VP.n17 VP.n16 24.4675
R2172 VP.n18 VP.n17 24.4675
R2173 VP.n29 VP.n8 10.2766
R2174 VP.n49 VP.n0 10.2766
R2175 VP.n24 VP.n9 10.2766
R2176 VP.n15 VP.n14 3.14395
R2177 VP.n26 VP.n25 0.354971
R2178 VP.n28 VP.n27 0.354971
R2179 VP.n51 VP.n50 0.354971
R2180 VP VP.n51 0.26696
R2181 VP.n15 VP.n12 0.189894
R2182 VP.n19 VP.n12 0.189894
R2183 VP.n20 VP.n19 0.189894
R2184 VP.n21 VP.n20 0.189894
R2185 VP.n21 VP.n10 0.189894
R2186 VP.n25 VP.n10 0.189894
R2187 VP.n28 VP.n7 0.189894
R2188 VP.n32 VP.n7 0.189894
R2189 VP.n33 VP.n32 0.189894
R2190 VP.n34 VP.n33 0.189894
R2191 VP.n34 VP.n5 0.189894
R2192 VP.n38 VP.n5 0.189894
R2193 VP.n39 VP.n38 0.189894
R2194 VP.n40 VP.n39 0.189894
R2195 VP.n40 VP.n3 0.189894
R2196 VP.n44 VP.n3 0.189894
R2197 VP.n45 VP.n44 0.189894
R2198 VP.n46 VP.n45 0.189894
R2199 VP.n46 VP.n1 0.189894
R2200 VP.n50 VP.n1 0.189894
R2201 VDD1.n76 VDD1.n0 756.745
R2202 VDD1.n157 VDD1.n81 756.745
R2203 VDD1.n77 VDD1.n76 585
R2204 VDD1.n75 VDD1.n74 585
R2205 VDD1.n73 VDD1.n3 585
R2206 VDD1.n7 VDD1.n4 585
R2207 VDD1.n68 VDD1.n67 585
R2208 VDD1.n66 VDD1.n65 585
R2209 VDD1.n9 VDD1.n8 585
R2210 VDD1.n60 VDD1.n59 585
R2211 VDD1.n58 VDD1.n57 585
R2212 VDD1.n13 VDD1.n12 585
R2213 VDD1.n52 VDD1.n51 585
R2214 VDD1.n50 VDD1.n49 585
R2215 VDD1.n17 VDD1.n16 585
R2216 VDD1.n44 VDD1.n43 585
R2217 VDD1.n42 VDD1.n41 585
R2218 VDD1.n21 VDD1.n20 585
R2219 VDD1.n36 VDD1.n35 585
R2220 VDD1.n34 VDD1.n33 585
R2221 VDD1.n25 VDD1.n24 585
R2222 VDD1.n28 VDD1.n27 585
R2223 VDD1.n108 VDD1.n107 585
R2224 VDD1.n105 VDD1.n104 585
R2225 VDD1.n114 VDD1.n113 585
R2226 VDD1.n116 VDD1.n115 585
R2227 VDD1.n101 VDD1.n100 585
R2228 VDD1.n122 VDD1.n121 585
R2229 VDD1.n124 VDD1.n123 585
R2230 VDD1.n97 VDD1.n96 585
R2231 VDD1.n130 VDD1.n129 585
R2232 VDD1.n132 VDD1.n131 585
R2233 VDD1.n93 VDD1.n92 585
R2234 VDD1.n138 VDD1.n137 585
R2235 VDD1.n140 VDD1.n139 585
R2236 VDD1.n89 VDD1.n88 585
R2237 VDD1.n146 VDD1.n145 585
R2238 VDD1.n149 VDD1.n148 585
R2239 VDD1.n147 VDD1.n85 585
R2240 VDD1.n154 VDD1.n84 585
R2241 VDD1.n156 VDD1.n155 585
R2242 VDD1.n158 VDD1.n157 585
R2243 VDD1.t5 VDD1.n26 327.466
R2244 VDD1.t3 VDD1.n106 327.466
R2245 VDD1.n76 VDD1.n75 171.744
R2246 VDD1.n75 VDD1.n3 171.744
R2247 VDD1.n7 VDD1.n3 171.744
R2248 VDD1.n67 VDD1.n7 171.744
R2249 VDD1.n67 VDD1.n66 171.744
R2250 VDD1.n66 VDD1.n8 171.744
R2251 VDD1.n59 VDD1.n8 171.744
R2252 VDD1.n59 VDD1.n58 171.744
R2253 VDD1.n58 VDD1.n12 171.744
R2254 VDD1.n51 VDD1.n12 171.744
R2255 VDD1.n51 VDD1.n50 171.744
R2256 VDD1.n50 VDD1.n16 171.744
R2257 VDD1.n43 VDD1.n16 171.744
R2258 VDD1.n43 VDD1.n42 171.744
R2259 VDD1.n42 VDD1.n20 171.744
R2260 VDD1.n35 VDD1.n20 171.744
R2261 VDD1.n35 VDD1.n34 171.744
R2262 VDD1.n34 VDD1.n24 171.744
R2263 VDD1.n27 VDD1.n24 171.744
R2264 VDD1.n107 VDD1.n104 171.744
R2265 VDD1.n114 VDD1.n104 171.744
R2266 VDD1.n115 VDD1.n114 171.744
R2267 VDD1.n115 VDD1.n100 171.744
R2268 VDD1.n122 VDD1.n100 171.744
R2269 VDD1.n123 VDD1.n122 171.744
R2270 VDD1.n123 VDD1.n96 171.744
R2271 VDD1.n130 VDD1.n96 171.744
R2272 VDD1.n131 VDD1.n130 171.744
R2273 VDD1.n131 VDD1.n92 171.744
R2274 VDD1.n138 VDD1.n92 171.744
R2275 VDD1.n139 VDD1.n138 171.744
R2276 VDD1.n139 VDD1.n88 171.744
R2277 VDD1.n146 VDD1.n88 171.744
R2278 VDD1.n148 VDD1.n146 171.744
R2279 VDD1.n148 VDD1.n147 171.744
R2280 VDD1.n147 VDD1.n84 171.744
R2281 VDD1.n156 VDD1.n84 171.744
R2282 VDD1.n157 VDD1.n156 171.744
R2283 VDD1.n27 VDD1.t5 85.8723
R2284 VDD1.n107 VDD1.t3 85.8723
R2285 VDD1.n163 VDD1.n162 72.0924
R2286 VDD1.n165 VDD1.n164 71.3482
R2287 VDD1 VDD1.n80 51.9029
R2288 VDD1.n163 VDD1.n161 51.7893
R2289 VDD1.n165 VDD1.n163 48.9384
R2290 VDD1.n28 VDD1.n26 16.3895
R2291 VDD1.n108 VDD1.n106 16.3895
R2292 VDD1.n74 VDD1.n73 13.1884
R2293 VDD1.n155 VDD1.n154 13.1884
R2294 VDD1.n77 VDD1.n2 12.8005
R2295 VDD1.n72 VDD1.n4 12.8005
R2296 VDD1.n29 VDD1.n25 12.8005
R2297 VDD1.n109 VDD1.n105 12.8005
R2298 VDD1.n153 VDD1.n85 12.8005
R2299 VDD1.n158 VDD1.n83 12.8005
R2300 VDD1.n78 VDD1.n0 12.0247
R2301 VDD1.n69 VDD1.n68 12.0247
R2302 VDD1.n33 VDD1.n32 12.0247
R2303 VDD1.n113 VDD1.n112 12.0247
R2304 VDD1.n150 VDD1.n149 12.0247
R2305 VDD1.n159 VDD1.n81 12.0247
R2306 VDD1.n65 VDD1.n6 11.249
R2307 VDD1.n36 VDD1.n23 11.249
R2308 VDD1.n116 VDD1.n103 11.249
R2309 VDD1.n145 VDD1.n87 11.249
R2310 VDD1.n64 VDD1.n9 10.4732
R2311 VDD1.n37 VDD1.n21 10.4732
R2312 VDD1.n117 VDD1.n101 10.4732
R2313 VDD1.n144 VDD1.n89 10.4732
R2314 VDD1.n61 VDD1.n60 9.69747
R2315 VDD1.n41 VDD1.n40 9.69747
R2316 VDD1.n121 VDD1.n120 9.69747
R2317 VDD1.n141 VDD1.n140 9.69747
R2318 VDD1.n80 VDD1.n79 9.45567
R2319 VDD1.n161 VDD1.n160 9.45567
R2320 VDD1.n54 VDD1.n53 9.3005
R2321 VDD1.n56 VDD1.n55 9.3005
R2322 VDD1.n11 VDD1.n10 9.3005
R2323 VDD1.n62 VDD1.n61 9.3005
R2324 VDD1.n64 VDD1.n63 9.3005
R2325 VDD1.n6 VDD1.n5 9.3005
R2326 VDD1.n70 VDD1.n69 9.3005
R2327 VDD1.n72 VDD1.n71 9.3005
R2328 VDD1.n79 VDD1.n78 9.3005
R2329 VDD1.n2 VDD1.n1 9.3005
R2330 VDD1.n15 VDD1.n14 9.3005
R2331 VDD1.n48 VDD1.n47 9.3005
R2332 VDD1.n46 VDD1.n45 9.3005
R2333 VDD1.n19 VDD1.n18 9.3005
R2334 VDD1.n40 VDD1.n39 9.3005
R2335 VDD1.n38 VDD1.n37 9.3005
R2336 VDD1.n23 VDD1.n22 9.3005
R2337 VDD1.n32 VDD1.n31 9.3005
R2338 VDD1.n30 VDD1.n29 9.3005
R2339 VDD1.n160 VDD1.n159 9.3005
R2340 VDD1.n83 VDD1.n82 9.3005
R2341 VDD1.n128 VDD1.n127 9.3005
R2342 VDD1.n126 VDD1.n125 9.3005
R2343 VDD1.n99 VDD1.n98 9.3005
R2344 VDD1.n120 VDD1.n119 9.3005
R2345 VDD1.n118 VDD1.n117 9.3005
R2346 VDD1.n103 VDD1.n102 9.3005
R2347 VDD1.n112 VDD1.n111 9.3005
R2348 VDD1.n110 VDD1.n109 9.3005
R2349 VDD1.n95 VDD1.n94 9.3005
R2350 VDD1.n134 VDD1.n133 9.3005
R2351 VDD1.n136 VDD1.n135 9.3005
R2352 VDD1.n91 VDD1.n90 9.3005
R2353 VDD1.n142 VDD1.n141 9.3005
R2354 VDD1.n144 VDD1.n143 9.3005
R2355 VDD1.n87 VDD1.n86 9.3005
R2356 VDD1.n151 VDD1.n150 9.3005
R2357 VDD1.n153 VDD1.n152 9.3005
R2358 VDD1.n57 VDD1.n11 8.92171
R2359 VDD1.n44 VDD1.n19 8.92171
R2360 VDD1.n124 VDD1.n99 8.92171
R2361 VDD1.n137 VDD1.n91 8.92171
R2362 VDD1.n56 VDD1.n13 8.14595
R2363 VDD1.n45 VDD1.n17 8.14595
R2364 VDD1.n125 VDD1.n97 8.14595
R2365 VDD1.n136 VDD1.n93 8.14595
R2366 VDD1.n53 VDD1.n52 7.3702
R2367 VDD1.n49 VDD1.n48 7.3702
R2368 VDD1.n129 VDD1.n128 7.3702
R2369 VDD1.n133 VDD1.n132 7.3702
R2370 VDD1.n52 VDD1.n15 6.59444
R2371 VDD1.n49 VDD1.n15 6.59444
R2372 VDD1.n129 VDD1.n95 6.59444
R2373 VDD1.n132 VDD1.n95 6.59444
R2374 VDD1.n53 VDD1.n13 5.81868
R2375 VDD1.n48 VDD1.n17 5.81868
R2376 VDD1.n128 VDD1.n97 5.81868
R2377 VDD1.n133 VDD1.n93 5.81868
R2378 VDD1.n57 VDD1.n56 5.04292
R2379 VDD1.n45 VDD1.n44 5.04292
R2380 VDD1.n125 VDD1.n124 5.04292
R2381 VDD1.n137 VDD1.n136 5.04292
R2382 VDD1.n60 VDD1.n11 4.26717
R2383 VDD1.n41 VDD1.n19 4.26717
R2384 VDD1.n121 VDD1.n99 4.26717
R2385 VDD1.n140 VDD1.n91 4.26717
R2386 VDD1.n30 VDD1.n26 3.70982
R2387 VDD1.n110 VDD1.n106 3.70982
R2388 VDD1.n61 VDD1.n9 3.49141
R2389 VDD1.n40 VDD1.n21 3.49141
R2390 VDD1.n120 VDD1.n101 3.49141
R2391 VDD1.n141 VDD1.n89 3.49141
R2392 VDD1.n65 VDD1.n64 2.71565
R2393 VDD1.n37 VDD1.n36 2.71565
R2394 VDD1.n117 VDD1.n116 2.71565
R2395 VDD1.n145 VDD1.n144 2.71565
R2396 VDD1.n164 VDD1.t4 2.21625
R2397 VDD1.n164 VDD1.t2 2.21625
R2398 VDD1.n162 VDD1.t1 2.21625
R2399 VDD1.n162 VDD1.t0 2.21625
R2400 VDD1.n80 VDD1.n0 1.93989
R2401 VDD1.n68 VDD1.n6 1.93989
R2402 VDD1.n33 VDD1.n23 1.93989
R2403 VDD1.n113 VDD1.n103 1.93989
R2404 VDD1.n149 VDD1.n87 1.93989
R2405 VDD1.n161 VDD1.n81 1.93989
R2406 VDD1.n78 VDD1.n77 1.16414
R2407 VDD1.n69 VDD1.n4 1.16414
R2408 VDD1.n32 VDD1.n25 1.16414
R2409 VDD1.n112 VDD1.n105 1.16414
R2410 VDD1.n150 VDD1.n85 1.16414
R2411 VDD1.n159 VDD1.n158 1.16414
R2412 VDD1 VDD1.n165 0.741879
R2413 VDD1.n74 VDD1.n2 0.388379
R2414 VDD1.n73 VDD1.n72 0.388379
R2415 VDD1.n29 VDD1.n28 0.388379
R2416 VDD1.n109 VDD1.n108 0.388379
R2417 VDD1.n154 VDD1.n153 0.388379
R2418 VDD1.n155 VDD1.n83 0.388379
R2419 VDD1.n79 VDD1.n1 0.155672
R2420 VDD1.n71 VDD1.n1 0.155672
R2421 VDD1.n71 VDD1.n70 0.155672
R2422 VDD1.n70 VDD1.n5 0.155672
R2423 VDD1.n63 VDD1.n5 0.155672
R2424 VDD1.n63 VDD1.n62 0.155672
R2425 VDD1.n62 VDD1.n10 0.155672
R2426 VDD1.n55 VDD1.n10 0.155672
R2427 VDD1.n55 VDD1.n54 0.155672
R2428 VDD1.n54 VDD1.n14 0.155672
R2429 VDD1.n47 VDD1.n14 0.155672
R2430 VDD1.n47 VDD1.n46 0.155672
R2431 VDD1.n46 VDD1.n18 0.155672
R2432 VDD1.n39 VDD1.n18 0.155672
R2433 VDD1.n39 VDD1.n38 0.155672
R2434 VDD1.n38 VDD1.n22 0.155672
R2435 VDD1.n31 VDD1.n22 0.155672
R2436 VDD1.n31 VDD1.n30 0.155672
R2437 VDD1.n111 VDD1.n110 0.155672
R2438 VDD1.n111 VDD1.n102 0.155672
R2439 VDD1.n118 VDD1.n102 0.155672
R2440 VDD1.n119 VDD1.n118 0.155672
R2441 VDD1.n119 VDD1.n98 0.155672
R2442 VDD1.n126 VDD1.n98 0.155672
R2443 VDD1.n127 VDD1.n126 0.155672
R2444 VDD1.n127 VDD1.n94 0.155672
R2445 VDD1.n134 VDD1.n94 0.155672
R2446 VDD1.n135 VDD1.n134 0.155672
R2447 VDD1.n135 VDD1.n90 0.155672
R2448 VDD1.n142 VDD1.n90 0.155672
R2449 VDD1.n143 VDD1.n142 0.155672
R2450 VDD1.n143 VDD1.n86 0.155672
R2451 VDD1.n151 VDD1.n86 0.155672
R2452 VDD1.n152 VDD1.n151 0.155672
R2453 VDD1.n152 VDD1.n82 0.155672
R2454 VDD1.n160 VDD1.n82 0.155672
C0 VN VDD1 0.151854f
C1 VP VDD2 0.524682f
C2 VN VDD2 8.503941f
C3 VDD1 VDD2 1.71184f
C4 w_n3938_n3902# B 11.501901f
C5 w_n3938_n3902# VTAIL 3.40782f
C6 B VTAIL 4.61724f
C7 w_n3938_n3902# VP 8.21431f
C8 B VP 2.22075f
C9 w_n3938_n3902# VN 7.70301f
C10 VP VTAIL 8.740219f
C11 B VN 1.36315f
C12 VN VTAIL 8.72595f
C13 w_n3938_n3902# VDD1 2.66464f
C14 VP VN 8.18189f
C15 B VDD1 2.51084f
C16 VTAIL VDD1 8.851691f
C17 w_n3938_n3902# VDD2 2.77465f
C18 VP VDD1 8.87333f
C19 B VDD2 2.60364f
C20 VTAIL VDD2 8.907969f
C21 VDD2 VSUBS 2.17817f
C22 VDD1 VSUBS 2.170015f
C23 VTAIL VSUBS 1.434805f
C24 VN VSUBS 6.68375f
C25 VP VSUBS 3.640818f
C26 B VSUBS 5.633744f
C27 w_n3938_n3902# VSUBS 0.188504p
C28 VDD1.n0 VSUBS 0.028545f
C29 VDD1.n1 VSUBS 0.027916f
C30 VDD1.n2 VSUBS 0.015001f
C31 VDD1.n3 VSUBS 0.035457f
C32 VDD1.n4 VSUBS 0.015883f
C33 VDD1.n5 VSUBS 0.027916f
C34 VDD1.n6 VSUBS 0.015001f
C35 VDD1.n7 VSUBS 0.035457f
C36 VDD1.n8 VSUBS 0.035457f
C37 VDD1.n9 VSUBS 0.015883f
C38 VDD1.n10 VSUBS 0.027916f
C39 VDD1.n11 VSUBS 0.015001f
C40 VDD1.n12 VSUBS 0.035457f
C41 VDD1.n13 VSUBS 0.015883f
C42 VDD1.n14 VSUBS 0.027916f
C43 VDD1.n15 VSUBS 0.015001f
C44 VDD1.n16 VSUBS 0.035457f
C45 VDD1.n17 VSUBS 0.015883f
C46 VDD1.n18 VSUBS 0.027916f
C47 VDD1.n19 VSUBS 0.015001f
C48 VDD1.n20 VSUBS 0.035457f
C49 VDD1.n21 VSUBS 0.015883f
C50 VDD1.n22 VSUBS 0.027916f
C51 VDD1.n23 VSUBS 0.015001f
C52 VDD1.n24 VSUBS 0.035457f
C53 VDD1.n25 VSUBS 0.015883f
C54 VDD1.n26 VSUBS 0.194067f
C55 VDD1.t5 VSUBS 0.075883f
C56 VDD1.n27 VSUBS 0.026593f
C57 VDD1.n28 VSUBS 0.022556f
C58 VDD1.n29 VSUBS 0.015001f
C59 VDD1.n30 VSUBS 1.74068f
C60 VDD1.n31 VSUBS 0.027916f
C61 VDD1.n32 VSUBS 0.015001f
C62 VDD1.n33 VSUBS 0.015883f
C63 VDD1.n34 VSUBS 0.035457f
C64 VDD1.n35 VSUBS 0.035457f
C65 VDD1.n36 VSUBS 0.015883f
C66 VDD1.n37 VSUBS 0.015001f
C67 VDD1.n38 VSUBS 0.027916f
C68 VDD1.n39 VSUBS 0.027916f
C69 VDD1.n40 VSUBS 0.015001f
C70 VDD1.n41 VSUBS 0.015883f
C71 VDD1.n42 VSUBS 0.035457f
C72 VDD1.n43 VSUBS 0.035457f
C73 VDD1.n44 VSUBS 0.015883f
C74 VDD1.n45 VSUBS 0.015001f
C75 VDD1.n46 VSUBS 0.027916f
C76 VDD1.n47 VSUBS 0.027916f
C77 VDD1.n48 VSUBS 0.015001f
C78 VDD1.n49 VSUBS 0.015883f
C79 VDD1.n50 VSUBS 0.035457f
C80 VDD1.n51 VSUBS 0.035457f
C81 VDD1.n52 VSUBS 0.015883f
C82 VDD1.n53 VSUBS 0.015001f
C83 VDD1.n54 VSUBS 0.027916f
C84 VDD1.n55 VSUBS 0.027916f
C85 VDD1.n56 VSUBS 0.015001f
C86 VDD1.n57 VSUBS 0.015883f
C87 VDD1.n58 VSUBS 0.035457f
C88 VDD1.n59 VSUBS 0.035457f
C89 VDD1.n60 VSUBS 0.015883f
C90 VDD1.n61 VSUBS 0.015001f
C91 VDD1.n62 VSUBS 0.027916f
C92 VDD1.n63 VSUBS 0.027916f
C93 VDD1.n64 VSUBS 0.015001f
C94 VDD1.n65 VSUBS 0.015883f
C95 VDD1.n66 VSUBS 0.035457f
C96 VDD1.n67 VSUBS 0.035457f
C97 VDD1.n68 VSUBS 0.015883f
C98 VDD1.n69 VSUBS 0.015001f
C99 VDD1.n70 VSUBS 0.027916f
C100 VDD1.n71 VSUBS 0.027916f
C101 VDD1.n72 VSUBS 0.015001f
C102 VDD1.n73 VSUBS 0.015442f
C103 VDD1.n74 VSUBS 0.015442f
C104 VDD1.n75 VSUBS 0.035457f
C105 VDD1.n76 VSUBS 0.078587f
C106 VDD1.n77 VSUBS 0.015883f
C107 VDD1.n78 VSUBS 0.015001f
C108 VDD1.n79 VSUBS 0.065671f
C109 VDD1.n80 VSUBS 0.071537f
C110 VDD1.n81 VSUBS 0.028545f
C111 VDD1.n82 VSUBS 0.027916f
C112 VDD1.n83 VSUBS 0.015001f
C113 VDD1.n84 VSUBS 0.035457f
C114 VDD1.n85 VSUBS 0.015883f
C115 VDD1.n86 VSUBS 0.027916f
C116 VDD1.n87 VSUBS 0.015001f
C117 VDD1.n88 VSUBS 0.035457f
C118 VDD1.n89 VSUBS 0.015883f
C119 VDD1.n90 VSUBS 0.027916f
C120 VDD1.n91 VSUBS 0.015001f
C121 VDD1.n92 VSUBS 0.035457f
C122 VDD1.n93 VSUBS 0.015883f
C123 VDD1.n94 VSUBS 0.027916f
C124 VDD1.n95 VSUBS 0.015001f
C125 VDD1.n96 VSUBS 0.035457f
C126 VDD1.n97 VSUBS 0.015883f
C127 VDD1.n98 VSUBS 0.027916f
C128 VDD1.n99 VSUBS 0.015001f
C129 VDD1.n100 VSUBS 0.035457f
C130 VDD1.n101 VSUBS 0.015883f
C131 VDD1.n102 VSUBS 0.027916f
C132 VDD1.n103 VSUBS 0.015001f
C133 VDD1.n104 VSUBS 0.035457f
C134 VDD1.n105 VSUBS 0.015883f
C135 VDD1.n106 VSUBS 0.194067f
C136 VDD1.t3 VSUBS 0.075883f
C137 VDD1.n107 VSUBS 0.026593f
C138 VDD1.n108 VSUBS 0.022556f
C139 VDD1.n109 VSUBS 0.015001f
C140 VDD1.n110 VSUBS 1.74068f
C141 VDD1.n111 VSUBS 0.027916f
C142 VDD1.n112 VSUBS 0.015001f
C143 VDD1.n113 VSUBS 0.015883f
C144 VDD1.n114 VSUBS 0.035457f
C145 VDD1.n115 VSUBS 0.035457f
C146 VDD1.n116 VSUBS 0.015883f
C147 VDD1.n117 VSUBS 0.015001f
C148 VDD1.n118 VSUBS 0.027916f
C149 VDD1.n119 VSUBS 0.027916f
C150 VDD1.n120 VSUBS 0.015001f
C151 VDD1.n121 VSUBS 0.015883f
C152 VDD1.n122 VSUBS 0.035457f
C153 VDD1.n123 VSUBS 0.035457f
C154 VDD1.n124 VSUBS 0.015883f
C155 VDD1.n125 VSUBS 0.015001f
C156 VDD1.n126 VSUBS 0.027916f
C157 VDD1.n127 VSUBS 0.027916f
C158 VDD1.n128 VSUBS 0.015001f
C159 VDD1.n129 VSUBS 0.015883f
C160 VDD1.n130 VSUBS 0.035457f
C161 VDD1.n131 VSUBS 0.035457f
C162 VDD1.n132 VSUBS 0.015883f
C163 VDD1.n133 VSUBS 0.015001f
C164 VDD1.n134 VSUBS 0.027916f
C165 VDD1.n135 VSUBS 0.027916f
C166 VDD1.n136 VSUBS 0.015001f
C167 VDD1.n137 VSUBS 0.015883f
C168 VDD1.n138 VSUBS 0.035457f
C169 VDD1.n139 VSUBS 0.035457f
C170 VDD1.n140 VSUBS 0.015883f
C171 VDD1.n141 VSUBS 0.015001f
C172 VDD1.n142 VSUBS 0.027916f
C173 VDD1.n143 VSUBS 0.027916f
C174 VDD1.n144 VSUBS 0.015001f
C175 VDD1.n145 VSUBS 0.015883f
C176 VDD1.n146 VSUBS 0.035457f
C177 VDD1.n147 VSUBS 0.035457f
C178 VDD1.n148 VSUBS 0.035457f
C179 VDD1.n149 VSUBS 0.015883f
C180 VDD1.n150 VSUBS 0.015001f
C181 VDD1.n151 VSUBS 0.027916f
C182 VDD1.n152 VSUBS 0.027916f
C183 VDD1.n153 VSUBS 0.015001f
C184 VDD1.n154 VSUBS 0.015442f
C185 VDD1.n155 VSUBS 0.015442f
C186 VDD1.n156 VSUBS 0.035457f
C187 VDD1.n157 VSUBS 0.078587f
C188 VDD1.n158 VSUBS 0.015883f
C189 VDD1.n159 VSUBS 0.015001f
C190 VDD1.n160 VSUBS 0.065671f
C191 VDD1.n161 VSUBS 0.070512f
C192 VDD1.t1 VSUBS 0.323622f
C193 VDD1.t0 VSUBS 0.323622f
C194 VDD1.n162 VSUBS 2.62887f
C195 VDD1.n163 VSUBS 4.01541f
C196 VDD1.t4 VSUBS 0.323622f
C197 VDD1.t2 VSUBS 0.323622f
C198 VDD1.n164 VSUBS 2.61961f
C199 VDD1.n165 VSUBS 3.88694f
C200 VP.t5 VSUBS 3.69391f
C201 VP.n0 VSUBS 1.38702f
C202 VP.n1 VSUBS 0.027201f
C203 VP.n2 VSUBS 0.030346f
C204 VP.n3 VSUBS 0.027201f
C205 VP.t4 VSUBS 3.69391f
C206 VP.n4 VSUBS 1.31063f
C207 VP.n5 VSUBS 0.027201f
C208 VP.n6 VSUBS 0.030346f
C209 VP.n7 VSUBS 0.027201f
C210 VP.t2 VSUBS 3.69391f
C211 VP.n8 VSUBS 1.38702f
C212 VP.t3 VSUBS 3.69391f
C213 VP.n9 VSUBS 1.38702f
C214 VP.n10 VSUBS 0.027201f
C215 VP.n11 VSUBS 0.030346f
C216 VP.n12 VSUBS 0.027201f
C217 VP.t1 VSUBS 3.69391f
C218 VP.n13 VSUBS 1.39215f
C219 VP.t0 VSUBS 4.05392f
C220 VP.n14 VSUBS 1.31782f
C221 VP.n15 VSUBS 0.332025f
C222 VP.n16 VSUBS 0.050695f
C223 VP.n17 VSUBS 0.050695f
C224 VP.n18 VSUBS 0.047382f
C225 VP.n19 VSUBS 0.027201f
C226 VP.n20 VSUBS 0.027201f
C227 VP.n21 VSUBS 0.027201f
C228 VP.n22 VSUBS 0.052389f
C229 VP.n23 VSUBS 0.050695f
C230 VP.n24 VSUBS 0.036179f
C231 VP.n25 VSUBS 0.043901f
C232 VP.n26 VSUBS 1.72187f
C233 VP.n27 VSUBS 1.74003f
C234 VP.n28 VSUBS 0.043901f
C235 VP.n29 VSUBS 0.036179f
C236 VP.n30 VSUBS 0.050695f
C237 VP.n31 VSUBS 0.052389f
C238 VP.n32 VSUBS 0.027201f
C239 VP.n33 VSUBS 0.027201f
C240 VP.n34 VSUBS 0.027201f
C241 VP.n35 VSUBS 0.047382f
C242 VP.n36 VSUBS 0.050695f
C243 VP.n37 VSUBS 0.050695f
C244 VP.n38 VSUBS 0.027201f
C245 VP.n39 VSUBS 0.027201f
C246 VP.n40 VSUBS 0.027201f
C247 VP.n41 VSUBS 0.050695f
C248 VP.n42 VSUBS 0.050695f
C249 VP.n43 VSUBS 0.047382f
C250 VP.n44 VSUBS 0.027201f
C251 VP.n45 VSUBS 0.027201f
C252 VP.n46 VSUBS 0.027201f
C253 VP.n47 VSUBS 0.052389f
C254 VP.n48 VSUBS 0.050695f
C255 VP.n49 VSUBS 0.036179f
C256 VP.n50 VSUBS 0.043901f
C257 VP.n51 VSUBS 0.07125f
C258 VTAIL.t9 VSUBS 0.333999f
C259 VTAIL.t11 VSUBS 0.333999f
C260 VTAIL.n0 VSUBS 2.53817f
C261 VTAIL.n1 VSUBS 0.945739f
C262 VTAIL.n2 VSUBS 0.029461f
C263 VTAIL.n3 VSUBS 0.028811f
C264 VTAIL.n4 VSUBS 0.015482f
C265 VTAIL.n5 VSUBS 0.036593f
C266 VTAIL.n6 VSUBS 0.016393f
C267 VTAIL.n7 VSUBS 0.028811f
C268 VTAIL.n8 VSUBS 0.015482f
C269 VTAIL.n9 VSUBS 0.036593f
C270 VTAIL.n10 VSUBS 0.016393f
C271 VTAIL.n11 VSUBS 0.028811f
C272 VTAIL.n12 VSUBS 0.015482f
C273 VTAIL.n13 VSUBS 0.036593f
C274 VTAIL.n14 VSUBS 0.016393f
C275 VTAIL.n15 VSUBS 0.028811f
C276 VTAIL.n16 VSUBS 0.015482f
C277 VTAIL.n17 VSUBS 0.036593f
C278 VTAIL.n18 VSUBS 0.016393f
C279 VTAIL.n19 VSUBS 0.028811f
C280 VTAIL.n20 VSUBS 0.015482f
C281 VTAIL.n21 VSUBS 0.036593f
C282 VTAIL.n22 VSUBS 0.016393f
C283 VTAIL.n23 VSUBS 0.028811f
C284 VTAIL.n24 VSUBS 0.015482f
C285 VTAIL.n25 VSUBS 0.036593f
C286 VTAIL.n26 VSUBS 0.016393f
C287 VTAIL.n27 VSUBS 0.200289f
C288 VTAIL.t0 VSUBS 0.078316f
C289 VTAIL.n28 VSUBS 0.027445f
C290 VTAIL.n29 VSUBS 0.023279f
C291 VTAIL.n30 VSUBS 0.015482f
C292 VTAIL.n31 VSUBS 1.79649f
C293 VTAIL.n32 VSUBS 0.028811f
C294 VTAIL.n33 VSUBS 0.015482f
C295 VTAIL.n34 VSUBS 0.016393f
C296 VTAIL.n35 VSUBS 0.036593f
C297 VTAIL.n36 VSUBS 0.036593f
C298 VTAIL.n37 VSUBS 0.016393f
C299 VTAIL.n38 VSUBS 0.015482f
C300 VTAIL.n39 VSUBS 0.028811f
C301 VTAIL.n40 VSUBS 0.028811f
C302 VTAIL.n41 VSUBS 0.015482f
C303 VTAIL.n42 VSUBS 0.016393f
C304 VTAIL.n43 VSUBS 0.036593f
C305 VTAIL.n44 VSUBS 0.036593f
C306 VTAIL.n45 VSUBS 0.016393f
C307 VTAIL.n46 VSUBS 0.015482f
C308 VTAIL.n47 VSUBS 0.028811f
C309 VTAIL.n48 VSUBS 0.028811f
C310 VTAIL.n49 VSUBS 0.015482f
C311 VTAIL.n50 VSUBS 0.016393f
C312 VTAIL.n51 VSUBS 0.036593f
C313 VTAIL.n52 VSUBS 0.036593f
C314 VTAIL.n53 VSUBS 0.016393f
C315 VTAIL.n54 VSUBS 0.015482f
C316 VTAIL.n55 VSUBS 0.028811f
C317 VTAIL.n56 VSUBS 0.028811f
C318 VTAIL.n57 VSUBS 0.015482f
C319 VTAIL.n58 VSUBS 0.016393f
C320 VTAIL.n59 VSUBS 0.036593f
C321 VTAIL.n60 VSUBS 0.036593f
C322 VTAIL.n61 VSUBS 0.016393f
C323 VTAIL.n62 VSUBS 0.015482f
C324 VTAIL.n63 VSUBS 0.028811f
C325 VTAIL.n64 VSUBS 0.028811f
C326 VTAIL.n65 VSUBS 0.015482f
C327 VTAIL.n66 VSUBS 0.016393f
C328 VTAIL.n67 VSUBS 0.036593f
C329 VTAIL.n68 VSUBS 0.036593f
C330 VTAIL.n69 VSUBS 0.036593f
C331 VTAIL.n70 VSUBS 0.016393f
C332 VTAIL.n71 VSUBS 0.015482f
C333 VTAIL.n72 VSUBS 0.028811f
C334 VTAIL.n73 VSUBS 0.028811f
C335 VTAIL.n74 VSUBS 0.015482f
C336 VTAIL.n75 VSUBS 0.015937f
C337 VTAIL.n76 VSUBS 0.015937f
C338 VTAIL.n77 VSUBS 0.036593f
C339 VTAIL.n78 VSUBS 0.081106f
C340 VTAIL.n79 VSUBS 0.016393f
C341 VTAIL.n80 VSUBS 0.015482f
C342 VTAIL.n81 VSUBS 0.067776f
C343 VTAIL.n82 VSUBS 0.040492f
C344 VTAIL.n83 VSUBS 0.514263f
C345 VTAIL.t2 VSUBS 0.333999f
C346 VTAIL.t5 VSUBS 0.333999f
C347 VTAIL.n84 VSUBS 2.53817f
C348 VTAIL.n85 VSUBS 3.1302f
C349 VTAIL.t10 VSUBS 0.333999f
C350 VTAIL.t7 VSUBS 0.333999f
C351 VTAIL.n86 VSUBS 2.53818f
C352 VTAIL.n87 VSUBS 3.13018f
C353 VTAIL.n88 VSUBS 0.029461f
C354 VTAIL.n89 VSUBS 0.028811f
C355 VTAIL.n90 VSUBS 0.015482f
C356 VTAIL.n91 VSUBS 0.036593f
C357 VTAIL.n92 VSUBS 0.016393f
C358 VTAIL.n93 VSUBS 0.028811f
C359 VTAIL.n94 VSUBS 0.015482f
C360 VTAIL.n95 VSUBS 0.036593f
C361 VTAIL.n96 VSUBS 0.036593f
C362 VTAIL.n97 VSUBS 0.016393f
C363 VTAIL.n98 VSUBS 0.028811f
C364 VTAIL.n99 VSUBS 0.015482f
C365 VTAIL.n100 VSUBS 0.036593f
C366 VTAIL.n101 VSUBS 0.016393f
C367 VTAIL.n102 VSUBS 0.028811f
C368 VTAIL.n103 VSUBS 0.015482f
C369 VTAIL.n104 VSUBS 0.036593f
C370 VTAIL.n105 VSUBS 0.016393f
C371 VTAIL.n106 VSUBS 0.028811f
C372 VTAIL.n107 VSUBS 0.015482f
C373 VTAIL.n108 VSUBS 0.036593f
C374 VTAIL.n109 VSUBS 0.016393f
C375 VTAIL.n110 VSUBS 0.028811f
C376 VTAIL.n111 VSUBS 0.015482f
C377 VTAIL.n112 VSUBS 0.036593f
C378 VTAIL.n113 VSUBS 0.016393f
C379 VTAIL.n114 VSUBS 0.200289f
C380 VTAIL.t8 VSUBS 0.078316f
C381 VTAIL.n115 VSUBS 0.027445f
C382 VTAIL.n116 VSUBS 0.023279f
C383 VTAIL.n117 VSUBS 0.015482f
C384 VTAIL.n118 VSUBS 1.79649f
C385 VTAIL.n119 VSUBS 0.028811f
C386 VTAIL.n120 VSUBS 0.015482f
C387 VTAIL.n121 VSUBS 0.016393f
C388 VTAIL.n122 VSUBS 0.036593f
C389 VTAIL.n123 VSUBS 0.036593f
C390 VTAIL.n124 VSUBS 0.016393f
C391 VTAIL.n125 VSUBS 0.015482f
C392 VTAIL.n126 VSUBS 0.028811f
C393 VTAIL.n127 VSUBS 0.028811f
C394 VTAIL.n128 VSUBS 0.015482f
C395 VTAIL.n129 VSUBS 0.016393f
C396 VTAIL.n130 VSUBS 0.036593f
C397 VTAIL.n131 VSUBS 0.036593f
C398 VTAIL.n132 VSUBS 0.016393f
C399 VTAIL.n133 VSUBS 0.015482f
C400 VTAIL.n134 VSUBS 0.028811f
C401 VTAIL.n135 VSUBS 0.028811f
C402 VTAIL.n136 VSUBS 0.015482f
C403 VTAIL.n137 VSUBS 0.016393f
C404 VTAIL.n138 VSUBS 0.036593f
C405 VTAIL.n139 VSUBS 0.036593f
C406 VTAIL.n140 VSUBS 0.016393f
C407 VTAIL.n141 VSUBS 0.015482f
C408 VTAIL.n142 VSUBS 0.028811f
C409 VTAIL.n143 VSUBS 0.028811f
C410 VTAIL.n144 VSUBS 0.015482f
C411 VTAIL.n145 VSUBS 0.016393f
C412 VTAIL.n146 VSUBS 0.036593f
C413 VTAIL.n147 VSUBS 0.036593f
C414 VTAIL.n148 VSUBS 0.016393f
C415 VTAIL.n149 VSUBS 0.015482f
C416 VTAIL.n150 VSUBS 0.028811f
C417 VTAIL.n151 VSUBS 0.028811f
C418 VTAIL.n152 VSUBS 0.015482f
C419 VTAIL.n153 VSUBS 0.016393f
C420 VTAIL.n154 VSUBS 0.036593f
C421 VTAIL.n155 VSUBS 0.036593f
C422 VTAIL.n156 VSUBS 0.016393f
C423 VTAIL.n157 VSUBS 0.015482f
C424 VTAIL.n158 VSUBS 0.028811f
C425 VTAIL.n159 VSUBS 0.028811f
C426 VTAIL.n160 VSUBS 0.015482f
C427 VTAIL.n161 VSUBS 0.015937f
C428 VTAIL.n162 VSUBS 0.015937f
C429 VTAIL.n163 VSUBS 0.036593f
C430 VTAIL.n164 VSUBS 0.081106f
C431 VTAIL.n165 VSUBS 0.016393f
C432 VTAIL.n166 VSUBS 0.015482f
C433 VTAIL.n167 VSUBS 0.067776f
C434 VTAIL.n168 VSUBS 0.040492f
C435 VTAIL.n169 VSUBS 0.514263f
C436 VTAIL.t3 VSUBS 0.333999f
C437 VTAIL.t4 VSUBS 0.333999f
C438 VTAIL.n170 VSUBS 2.53818f
C439 VTAIL.n171 VSUBS 1.16301f
C440 VTAIL.n172 VSUBS 0.029461f
C441 VTAIL.n173 VSUBS 0.028811f
C442 VTAIL.n174 VSUBS 0.015482f
C443 VTAIL.n175 VSUBS 0.036593f
C444 VTAIL.n176 VSUBS 0.016393f
C445 VTAIL.n177 VSUBS 0.028811f
C446 VTAIL.n178 VSUBS 0.015482f
C447 VTAIL.n179 VSUBS 0.036593f
C448 VTAIL.n180 VSUBS 0.036593f
C449 VTAIL.n181 VSUBS 0.016393f
C450 VTAIL.n182 VSUBS 0.028811f
C451 VTAIL.n183 VSUBS 0.015482f
C452 VTAIL.n184 VSUBS 0.036593f
C453 VTAIL.n185 VSUBS 0.016393f
C454 VTAIL.n186 VSUBS 0.028811f
C455 VTAIL.n187 VSUBS 0.015482f
C456 VTAIL.n188 VSUBS 0.036593f
C457 VTAIL.n189 VSUBS 0.016393f
C458 VTAIL.n190 VSUBS 0.028811f
C459 VTAIL.n191 VSUBS 0.015482f
C460 VTAIL.n192 VSUBS 0.036593f
C461 VTAIL.n193 VSUBS 0.016393f
C462 VTAIL.n194 VSUBS 0.028811f
C463 VTAIL.n195 VSUBS 0.015482f
C464 VTAIL.n196 VSUBS 0.036593f
C465 VTAIL.n197 VSUBS 0.016393f
C466 VTAIL.n198 VSUBS 0.200289f
C467 VTAIL.t1 VSUBS 0.078316f
C468 VTAIL.n199 VSUBS 0.027445f
C469 VTAIL.n200 VSUBS 0.023279f
C470 VTAIL.n201 VSUBS 0.015482f
C471 VTAIL.n202 VSUBS 1.79649f
C472 VTAIL.n203 VSUBS 0.028811f
C473 VTAIL.n204 VSUBS 0.015482f
C474 VTAIL.n205 VSUBS 0.016393f
C475 VTAIL.n206 VSUBS 0.036593f
C476 VTAIL.n207 VSUBS 0.036593f
C477 VTAIL.n208 VSUBS 0.016393f
C478 VTAIL.n209 VSUBS 0.015482f
C479 VTAIL.n210 VSUBS 0.028811f
C480 VTAIL.n211 VSUBS 0.028811f
C481 VTAIL.n212 VSUBS 0.015482f
C482 VTAIL.n213 VSUBS 0.016393f
C483 VTAIL.n214 VSUBS 0.036593f
C484 VTAIL.n215 VSUBS 0.036593f
C485 VTAIL.n216 VSUBS 0.016393f
C486 VTAIL.n217 VSUBS 0.015482f
C487 VTAIL.n218 VSUBS 0.028811f
C488 VTAIL.n219 VSUBS 0.028811f
C489 VTAIL.n220 VSUBS 0.015482f
C490 VTAIL.n221 VSUBS 0.016393f
C491 VTAIL.n222 VSUBS 0.036593f
C492 VTAIL.n223 VSUBS 0.036593f
C493 VTAIL.n224 VSUBS 0.016393f
C494 VTAIL.n225 VSUBS 0.015482f
C495 VTAIL.n226 VSUBS 0.028811f
C496 VTAIL.n227 VSUBS 0.028811f
C497 VTAIL.n228 VSUBS 0.015482f
C498 VTAIL.n229 VSUBS 0.016393f
C499 VTAIL.n230 VSUBS 0.036593f
C500 VTAIL.n231 VSUBS 0.036593f
C501 VTAIL.n232 VSUBS 0.016393f
C502 VTAIL.n233 VSUBS 0.015482f
C503 VTAIL.n234 VSUBS 0.028811f
C504 VTAIL.n235 VSUBS 0.028811f
C505 VTAIL.n236 VSUBS 0.015482f
C506 VTAIL.n237 VSUBS 0.016393f
C507 VTAIL.n238 VSUBS 0.036593f
C508 VTAIL.n239 VSUBS 0.036593f
C509 VTAIL.n240 VSUBS 0.016393f
C510 VTAIL.n241 VSUBS 0.015482f
C511 VTAIL.n242 VSUBS 0.028811f
C512 VTAIL.n243 VSUBS 0.028811f
C513 VTAIL.n244 VSUBS 0.015482f
C514 VTAIL.n245 VSUBS 0.015937f
C515 VTAIL.n246 VSUBS 0.015937f
C516 VTAIL.n247 VSUBS 0.036593f
C517 VTAIL.n248 VSUBS 0.081106f
C518 VTAIL.n249 VSUBS 0.016393f
C519 VTAIL.n250 VSUBS 0.015482f
C520 VTAIL.n251 VSUBS 0.067776f
C521 VTAIL.n252 VSUBS 0.040492f
C522 VTAIL.n253 VSUBS 2.18453f
C523 VTAIL.n254 VSUBS 0.029461f
C524 VTAIL.n255 VSUBS 0.028811f
C525 VTAIL.n256 VSUBS 0.015482f
C526 VTAIL.n257 VSUBS 0.036593f
C527 VTAIL.n258 VSUBS 0.016393f
C528 VTAIL.n259 VSUBS 0.028811f
C529 VTAIL.n260 VSUBS 0.015482f
C530 VTAIL.n261 VSUBS 0.036593f
C531 VTAIL.n262 VSUBS 0.016393f
C532 VTAIL.n263 VSUBS 0.028811f
C533 VTAIL.n264 VSUBS 0.015482f
C534 VTAIL.n265 VSUBS 0.036593f
C535 VTAIL.n266 VSUBS 0.016393f
C536 VTAIL.n267 VSUBS 0.028811f
C537 VTAIL.n268 VSUBS 0.015482f
C538 VTAIL.n269 VSUBS 0.036593f
C539 VTAIL.n270 VSUBS 0.016393f
C540 VTAIL.n271 VSUBS 0.028811f
C541 VTAIL.n272 VSUBS 0.015482f
C542 VTAIL.n273 VSUBS 0.036593f
C543 VTAIL.n274 VSUBS 0.016393f
C544 VTAIL.n275 VSUBS 0.028811f
C545 VTAIL.n276 VSUBS 0.015482f
C546 VTAIL.n277 VSUBS 0.036593f
C547 VTAIL.n278 VSUBS 0.016393f
C548 VTAIL.n279 VSUBS 0.200289f
C549 VTAIL.t6 VSUBS 0.078316f
C550 VTAIL.n280 VSUBS 0.027445f
C551 VTAIL.n281 VSUBS 0.023279f
C552 VTAIL.n282 VSUBS 0.015482f
C553 VTAIL.n283 VSUBS 1.79649f
C554 VTAIL.n284 VSUBS 0.028811f
C555 VTAIL.n285 VSUBS 0.015482f
C556 VTAIL.n286 VSUBS 0.016393f
C557 VTAIL.n287 VSUBS 0.036593f
C558 VTAIL.n288 VSUBS 0.036593f
C559 VTAIL.n289 VSUBS 0.016393f
C560 VTAIL.n290 VSUBS 0.015482f
C561 VTAIL.n291 VSUBS 0.028811f
C562 VTAIL.n292 VSUBS 0.028811f
C563 VTAIL.n293 VSUBS 0.015482f
C564 VTAIL.n294 VSUBS 0.016393f
C565 VTAIL.n295 VSUBS 0.036593f
C566 VTAIL.n296 VSUBS 0.036593f
C567 VTAIL.n297 VSUBS 0.016393f
C568 VTAIL.n298 VSUBS 0.015482f
C569 VTAIL.n299 VSUBS 0.028811f
C570 VTAIL.n300 VSUBS 0.028811f
C571 VTAIL.n301 VSUBS 0.015482f
C572 VTAIL.n302 VSUBS 0.016393f
C573 VTAIL.n303 VSUBS 0.036593f
C574 VTAIL.n304 VSUBS 0.036593f
C575 VTAIL.n305 VSUBS 0.016393f
C576 VTAIL.n306 VSUBS 0.015482f
C577 VTAIL.n307 VSUBS 0.028811f
C578 VTAIL.n308 VSUBS 0.028811f
C579 VTAIL.n309 VSUBS 0.015482f
C580 VTAIL.n310 VSUBS 0.016393f
C581 VTAIL.n311 VSUBS 0.036593f
C582 VTAIL.n312 VSUBS 0.036593f
C583 VTAIL.n313 VSUBS 0.016393f
C584 VTAIL.n314 VSUBS 0.015482f
C585 VTAIL.n315 VSUBS 0.028811f
C586 VTAIL.n316 VSUBS 0.028811f
C587 VTAIL.n317 VSUBS 0.015482f
C588 VTAIL.n318 VSUBS 0.016393f
C589 VTAIL.n319 VSUBS 0.036593f
C590 VTAIL.n320 VSUBS 0.036593f
C591 VTAIL.n321 VSUBS 0.036593f
C592 VTAIL.n322 VSUBS 0.016393f
C593 VTAIL.n323 VSUBS 0.015482f
C594 VTAIL.n324 VSUBS 0.028811f
C595 VTAIL.n325 VSUBS 0.028811f
C596 VTAIL.n326 VSUBS 0.015482f
C597 VTAIL.n327 VSUBS 0.015937f
C598 VTAIL.n328 VSUBS 0.015937f
C599 VTAIL.n329 VSUBS 0.036593f
C600 VTAIL.n330 VSUBS 0.081106f
C601 VTAIL.n331 VSUBS 0.016393f
C602 VTAIL.n332 VSUBS 0.015482f
C603 VTAIL.n333 VSUBS 0.067776f
C604 VTAIL.n334 VSUBS 0.040492f
C605 VTAIL.n335 VSUBS 2.10489f
C606 VDD2.n0 VSUBS 0.028424f
C607 VDD2.n1 VSUBS 0.027798f
C608 VDD2.n2 VSUBS 0.014937f
C609 VDD2.n3 VSUBS 0.035307f
C610 VDD2.n4 VSUBS 0.015816f
C611 VDD2.n5 VSUBS 0.027798f
C612 VDD2.n6 VSUBS 0.014937f
C613 VDD2.n7 VSUBS 0.035307f
C614 VDD2.n8 VSUBS 0.015816f
C615 VDD2.n9 VSUBS 0.027798f
C616 VDD2.n10 VSUBS 0.014937f
C617 VDD2.n11 VSUBS 0.035307f
C618 VDD2.n12 VSUBS 0.015816f
C619 VDD2.n13 VSUBS 0.027798f
C620 VDD2.n14 VSUBS 0.014937f
C621 VDD2.n15 VSUBS 0.035307f
C622 VDD2.n16 VSUBS 0.015816f
C623 VDD2.n17 VSUBS 0.027798f
C624 VDD2.n18 VSUBS 0.014937f
C625 VDD2.n19 VSUBS 0.035307f
C626 VDD2.n20 VSUBS 0.015816f
C627 VDD2.n21 VSUBS 0.027798f
C628 VDD2.n22 VSUBS 0.014937f
C629 VDD2.n23 VSUBS 0.035307f
C630 VDD2.n24 VSUBS 0.015816f
C631 VDD2.n25 VSUBS 0.193246f
C632 VDD2.t4 VSUBS 0.075562f
C633 VDD2.n26 VSUBS 0.02648f
C634 VDD2.n27 VSUBS 0.02246f
C635 VDD2.n28 VSUBS 0.014937f
C636 VDD2.n29 VSUBS 1.73331f
C637 VDD2.n30 VSUBS 0.027798f
C638 VDD2.n31 VSUBS 0.014937f
C639 VDD2.n32 VSUBS 0.015816f
C640 VDD2.n33 VSUBS 0.035307f
C641 VDD2.n34 VSUBS 0.035307f
C642 VDD2.n35 VSUBS 0.015816f
C643 VDD2.n36 VSUBS 0.014937f
C644 VDD2.n37 VSUBS 0.027798f
C645 VDD2.n38 VSUBS 0.027798f
C646 VDD2.n39 VSUBS 0.014937f
C647 VDD2.n40 VSUBS 0.015816f
C648 VDD2.n41 VSUBS 0.035307f
C649 VDD2.n42 VSUBS 0.035307f
C650 VDD2.n43 VSUBS 0.015816f
C651 VDD2.n44 VSUBS 0.014937f
C652 VDD2.n45 VSUBS 0.027798f
C653 VDD2.n46 VSUBS 0.027798f
C654 VDD2.n47 VSUBS 0.014937f
C655 VDD2.n48 VSUBS 0.015816f
C656 VDD2.n49 VSUBS 0.035307f
C657 VDD2.n50 VSUBS 0.035307f
C658 VDD2.n51 VSUBS 0.015816f
C659 VDD2.n52 VSUBS 0.014937f
C660 VDD2.n53 VSUBS 0.027798f
C661 VDD2.n54 VSUBS 0.027798f
C662 VDD2.n55 VSUBS 0.014937f
C663 VDD2.n56 VSUBS 0.015816f
C664 VDD2.n57 VSUBS 0.035307f
C665 VDD2.n58 VSUBS 0.035307f
C666 VDD2.n59 VSUBS 0.015816f
C667 VDD2.n60 VSUBS 0.014937f
C668 VDD2.n61 VSUBS 0.027798f
C669 VDD2.n62 VSUBS 0.027798f
C670 VDD2.n63 VSUBS 0.014937f
C671 VDD2.n64 VSUBS 0.015816f
C672 VDD2.n65 VSUBS 0.035307f
C673 VDD2.n66 VSUBS 0.035307f
C674 VDD2.n67 VSUBS 0.035307f
C675 VDD2.n68 VSUBS 0.015816f
C676 VDD2.n69 VSUBS 0.014937f
C677 VDD2.n70 VSUBS 0.027798f
C678 VDD2.n71 VSUBS 0.027798f
C679 VDD2.n72 VSUBS 0.014937f
C680 VDD2.n73 VSUBS 0.015377f
C681 VDD2.n74 VSUBS 0.015377f
C682 VDD2.n75 VSUBS 0.035307f
C683 VDD2.n76 VSUBS 0.078254f
C684 VDD2.n77 VSUBS 0.015816f
C685 VDD2.n78 VSUBS 0.014937f
C686 VDD2.n79 VSUBS 0.065393f
C687 VDD2.n80 VSUBS 0.070214f
C688 VDD2.t2 VSUBS 0.322252f
C689 VDD2.t0 VSUBS 0.322252f
C690 VDD2.n81 VSUBS 2.61775f
C691 VDD2.n82 VSUBS 3.83494f
C692 VDD2.n83 VSUBS 0.028424f
C693 VDD2.n84 VSUBS 0.027798f
C694 VDD2.n85 VSUBS 0.014937f
C695 VDD2.n86 VSUBS 0.035307f
C696 VDD2.n87 VSUBS 0.015816f
C697 VDD2.n88 VSUBS 0.027798f
C698 VDD2.n89 VSUBS 0.014937f
C699 VDD2.n90 VSUBS 0.035307f
C700 VDD2.n91 VSUBS 0.035307f
C701 VDD2.n92 VSUBS 0.015816f
C702 VDD2.n93 VSUBS 0.027798f
C703 VDD2.n94 VSUBS 0.014937f
C704 VDD2.n95 VSUBS 0.035307f
C705 VDD2.n96 VSUBS 0.015816f
C706 VDD2.n97 VSUBS 0.027798f
C707 VDD2.n98 VSUBS 0.014937f
C708 VDD2.n99 VSUBS 0.035307f
C709 VDD2.n100 VSUBS 0.015816f
C710 VDD2.n101 VSUBS 0.027798f
C711 VDD2.n102 VSUBS 0.014937f
C712 VDD2.n103 VSUBS 0.035307f
C713 VDD2.n104 VSUBS 0.015816f
C714 VDD2.n105 VSUBS 0.027798f
C715 VDD2.n106 VSUBS 0.014937f
C716 VDD2.n107 VSUBS 0.035307f
C717 VDD2.n108 VSUBS 0.015816f
C718 VDD2.n109 VSUBS 0.193246f
C719 VDD2.t3 VSUBS 0.075562f
C720 VDD2.n110 VSUBS 0.02648f
C721 VDD2.n111 VSUBS 0.02246f
C722 VDD2.n112 VSUBS 0.014937f
C723 VDD2.n113 VSUBS 1.73331f
C724 VDD2.n114 VSUBS 0.027798f
C725 VDD2.n115 VSUBS 0.014937f
C726 VDD2.n116 VSUBS 0.015816f
C727 VDD2.n117 VSUBS 0.035307f
C728 VDD2.n118 VSUBS 0.035307f
C729 VDD2.n119 VSUBS 0.015816f
C730 VDD2.n120 VSUBS 0.014937f
C731 VDD2.n121 VSUBS 0.027798f
C732 VDD2.n122 VSUBS 0.027798f
C733 VDD2.n123 VSUBS 0.014937f
C734 VDD2.n124 VSUBS 0.015816f
C735 VDD2.n125 VSUBS 0.035307f
C736 VDD2.n126 VSUBS 0.035307f
C737 VDD2.n127 VSUBS 0.015816f
C738 VDD2.n128 VSUBS 0.014937f
C739 VDD2.n129 VSUBS 0.027798f
C740 VDD2.n130 VSUBS 0.027798f
C741 VDD2.n131 VSUBS 0.014937f
C742 VDD2.n132 VSUBS 0.015816f
C743 VDD2.n133 VSUBS 0.035307f
C744 VDD2.n134 VSUBS 0.035307f
C745 VDD2.n135 VSUBS 0.015816f
C746 VDD2.n136 VSUBS 0.014937f
C747 VDD2.n137 VSUBS 0.027798f
C748 VDD2.n138 VSUBS 0.027798f
C749 VDD2.n139 VSUBS 0.014937f
C750 VDD2.n140 VSUBS 0.015816f
C751 VDD2.n141 VSUBS 0.035307f
C752 VDD2.n142 VSUBS 0.035307f
C753 VDD2.n143 VSUBS 0.015816f
C754 VDD2.n144 VSUBS 0.014937f
C755 VDD2.n145 VSUBS 0.027798f
C756 VDD2.n146 VSUBS 0.027798f
C757 VDD2.n147 VSUBS 0.014937f
C758 VDD2.n148 VSUBS 0.015816f
C759 VDD2.n149 VSUBS 0.035307f
C760 VDD2.n150 VSUBS 0.035307f
C761 VDD2.n151 VSUBS 0.015816f
C762 VDD2.n152 VSUBS 0.014937f
C763 VDD2.n153 VSUBS 0.027798f
C764 VDD2.n154 VSUBS 0.027798f
C765 VDD2.n155 VSUBS 0.014937f
C766 VDD2.n156 VSUBS 0.015377f
C767 VDD2.n157 VSUBS 0.015377f
C768 VDD2.n158 VSUBS 0.035307f
C769 VDD2.n159 VSUBS 0.078254f
C770 VDD2.n160 VSUBS 0.015816f
C771 VDD2.n161 VSUBS 0.014937f
C772 VDD2.n162 VSUBS 0.065393f
C773 VDD2.n163 VSUBS 0.058252f
C774 VDD2.n164 VSUBS 3.31297f
C775 VDD2.t1 VSUBS 0.322252f
C776 VDD2.t5 VSUBS 0.322252f
C777 VDD2.n165 VSUBS 2.6177f
C778 VN.t5 VSUBS 3.37402f
C779 VN.n0 VSUBS 1.2669f
C780 VN.n1 VSUBS 0.024845f
C781 VN.n2 VSUBS 0.027718f
C782 VN.n3 VSUBS 0.024845f
C783 VN.t0 VSUBS 3.37402f
C784 VN.n4 VSUBS 1.27159f
C785 VN.t2 VSUBS 3.70286f
C786 VN.n5 VSUBS 1.2037f
C787 VN.n6 VSUBS 0.303271f
C788 VN.n7 VSUBS 0.046305f
C789 VN.n8 VSUBS 0.046305f
C790 VN.n9 VSUBS 0.043278f
C791 VN.n10 VSUBS 0.024845f
C792 VN.n11 VSUBS 0.024845f
C793 VN.n12 VSUBS 0.024845f
C794 VN.n13 VSUBS 0.047852f
C795 VN.n14 VSUBS 0.046305f
C796 VN.n15 VSUBS 0.033046f
C797 VN.n16 VSUBS 0.0401f
C798 VN.n17 VSUBS 0.06508f
C799 VN.t1 VSUBS 3.37402f
C800 VN.n18 VSUBS 1.2669f
C801 VN.n19 VSUBS 0.024845f
C802 VN.n20 VSUBS 0.027718f
C803 VN.n21 VSUBS 0.024845f
C804 VN.t4 VSUBS 3.37402f
C805 VN.n22 VSUBS 1.27159f
C806 VN.t3 VSUBS 3.70286f
C807 VN.n23 VSUBS 1.2037f
C808 VN.n24 VSUBS 0.303271f
C809 VN.n25 VSUBS 0.046305f
C810 VN.n26 VSUBS 0.046305f
C811 VN.n27 VSUBS 0.043278f
C812 VN.n28 VSUBS 0.024845f
C813 VN.n29 VSUBS 0.024845f
C814 VN.n30 VSUBS 0.024845f
C815 VN.n31 VSUBS 0.047852f
C816 VN.n32 VSUBS 0.046305f
C817 VN.n33 VSUBS 0.033046f
C818 VN.n34 VSUBS 0.0401f
C819 VN.n35 VSUBS 1.58267f
C820 B.n0 VSUBS 0.006968f
C821 B.n1 VSUBS 0.006968f
C822 B.n2 VSUBS 0.010305f
C823 B.n3 VSUBS 0.007897f
C824 B.n4 VSUBS 0.007897f
C825 B.n5 VSUBS 0.007897f
C826 B.n6 VSUBS 0.007897f
C827 B.n7 VSUBS 0.007897f
C828 B.n8 VSUBS 0.007897f
C829 B.n9 VSUBS 0.007897f
C830 B.n10 VSUBS 0.007897f
C831 B.n11 VSUBS 0.007897f
C832 B.n12 VSUBS 0.007897f
C833 B.n13 VSUBS 0.007897f
C834 B.n14 VSUBS 0.007897f
C835 B.n15 VSUBS 0.007897f
C836 B.n16 VSUBS 0.007897f
C837 B.n17 VSUBS 0.007897f
C838 B.n18 VSUBS 0.007897f
C839 B.n19 VSUBS 0.007897f
C840 B.n20 VSUBS 0.007897f
C841 B.n21 VSUBS 0.007897f
C842 B.n22 VSUBS 0.007897f
C843 B.n23 VSUBS 0.007897f
C844 B.n24 VSUBS 0.007897f
C845 B.n25 VSUBS 0.007897f
C846 B.n26 VSUBS 0.007897f
C847 B.n27 VSUBS 0.020056f
C848 B.n28 VSUBS 0.007897f
C849 B.n29 VSUBS 0.007897f
C850 B.n30 VSUBS 0.007897f
C851 B.n31 VSUBS 0.007897f
C852 B.n32 VSUBS 0.007897f
C853 B.n33 VSUBS 0.007897f
C854 B.n34 VSUBS 0.007897f
C855 B.n35 VSUBS 0.007897f
C856 B.n36 VSUBS 0.007897f
C857 B.n37 VSUBS 0.007897f
C858 B.n38 VSUBS 0.007897f
C859 B.n39 VSUBS 0.007897f
C860 B.n40 VSUBS 0.007897f
C861 B.n41 VSUBS 0.007897f
C862 B.n42 VSUBS 0.007897f
C863 B.n43 VSUBS 0.007897f
C864 B.n44 VSUBS 0.007897f
C865 B.n45 VSUBS 0.007897f
C866 B.n46 VSUBS 0.007897f
C867 B.n47 VSUBS 0.007897f
C868 B.n48 VSUBS 0.007897f
C869 B.n49 VSUBS 0.007897f
C870 B.n50 VSUBS 0.007897f
C871 B.n51 VSUBS 0.007897f
C872 B.t4 VSUBS 0.306542f
C873 B.t5 VSUBS 0.352557f
C874 B.t3 VSUBS 2.56104f
C875 B.n52 VSUBS 0.55955f
C876 B.n53 VSUBS 0.328155f
C877 B.n54 VSUBS 0.018296f
C878 B.n55 VSUBS 0.007897f
C879 B.n56 VSUBS 0.007897f
C880 B.n57 VSUBS 0.007897f
C881 B.n58 VSUBS 0.007897f
C882 B.n59 VSUBS 0.007897f
C883 B.t10 VSUBS 0.306545f
C884 B.t11 VSUBS 0.352561f
C885 B.t9 VSUBS 2.56104f
C886 B.n60 VSUBS 0.559547f
C887 B.n61 VSUBS 0.328152f
C888 B.n62 VSUBS 0.007897f
C889 B.n63 VSUBS 0.007897f
C890 B.n64 VSUBS 0.007897f
C891 B.n65 VSUBS 0.007897f
C892 B.n66 VSUBS 0.007897f
C893 B.n67 VSUBS 0.007897f
C894 B.n68 VSUBS 0.007897f
C895 B.n69 VSUBS 0.007897f
C896 B.n70 VSUBS 0.007897f
C897 B.n71 VSUBS 0.007897f
C898 B.n72 VSUBS 0.007897f
C899 B.n73 VSUBS 0.007897f
C900 B.n74 VSUBS 0.007897f
C901 B.n75 VSUBS 0.007897f
C902 B.n76 VSUBS 0.007897f
C903 B.n77 VSUBS 0.007897f
C904 B.n78 VSUBS 0.007897f
C905 B.n79 VSUBS 0.007897f
C906 B.n80 VSUBS 0.007897f
C907 B.n81 VSUBS 0.007897f
C908 B.n82 VSUBS 0.007897f
C909 B.n83 VSUBS 0.007897f
C910 B.n84 VSUBS 0.007897f
C911 B.n85 VSUBS 0.007897f
C912 B.n86 VSUBS 0.020056f
C913 B.n87 VSUBS 0.007897f
C914 B.n88 VSUBS 0.007897f
C915 B.n89 VSUBS 0.007897f
C916 B.n90 VSUBS 0.007897f
C917 B.n91 VSUBS 0.007897f
C918 B.n92 VSUBS 0.007897f
C919 B.n93 VSUBS 0.007897f
C920 B.n94 VSUBS 0.007897f
C921 B.n95 VSUBS 0.007897f
C922 B.n96 VSUBS 0.007897f
C923 B.n97 VSUBS 0.007897f
C924 B.n98 VSUBS 0.007897f
C925 B.n99 VSUBS 0.007897f
C926 B.n100 VSUBS 0.007897f
C927 B.n101 VSUBS 0.007897f
C928 B.n102 VSUBS 0.007897f
C929 B.n103 VSUBS 0.007897f
C930 B.n104 VSUBS 0.007897f
C931 B.n105 VSUBS 0.007897f
C932 B.n106 VSUBS 0.007897f
C933 B.n107 VSUBS 0.007897f
C934 B.n108 VSUBS 0.007897f
C935 B.n109 VSUBS 0.007897f
C936 B.n110 VSUBS 0.007897f
C937 B.n111 VSUBS 0.007897f
C938 B.n112 VSUBS 0.007897f
C939 B.n113 VSUBS 0.007897f
C940 B.n114 VSUBS 0.007897f
C941 B.n115 VSUBS 0.007897f
C942 B.n116 VSUBS 0.007897f
C943 B.n117 VSUBS 0.007897f
C944 B.n118 VSUBS 0.007897f
C945 B.n119 VSUBS 0.007897f
C946 B.n120 VSUBS 0.007897f
C947 B.n121 VSUBS 0.007897f
C948 B.n122 VSUBS 0.007897f
C949 B.n123 VSUBS 0.007897f
C950 B.n124 VSUBS 0.007897f
C951 B.n125 VSUBS 0.007897f
C952 B.n126 VSUBS 0.007897f
C953 B.n127 VSUBS 0.007897f
C954 B.n128 VSUBS 0.007897f
C955 B.n129 VSUBS 0.007897f
C956 B.n130 VSUBS 0.007897f
C957 B.n131 VSUBS 0.007897f
C958 B.n132 VSUBS 0.007897f
C959 B.n133 VSUBS 0.007897f
C960 B.n134 VSUBS 0.007897f
C961 B.n135 VSUBS 0.007897f
C962 B.n136 VSUBS 0.007897f
C963 B.n137 VSUBS 0.007897f
C964 B.n138 VSUBS 0.020017f
C965 B.n139 VSUBS 0.007897f
C966 B.n140 VSUBS 0.007897f
C967 B.n141 VSUBS 0.007897f
C968 B.n142 VSUBS 0.007897f
C969 B.n143 VSUBS 0.007897f
C970 B.n144 VSUBS 0.007897f
C971 B.n145 VSUBS 0.007897f
C972 B.n146 VSUBS 0.007897f
C973 B.n147 VSUBS 0.007897f
C974 B.n148 VSUBS 0.007897f
C975 B.n149 VSUBS 0.007897f
C976 B.n150 VSUBS 0.007897f
C977 B.n151 VSUBS 0.007897f
C978 B.n152 VSUBS 0.007897f
C979 B.n153 VSUBS 0.007897f
C980 B.n154 VSUBS 0.007897f
C981 B.n155 VSUBS 0.007897f
C982 B.n156 VSUBS 0.007897f
C983 B.n157 VSUBS 0.007897f
C984 B.n158 VSUBS 0.007897f
C985 B.n159 VSUBS 0.007897f
C986 B.n160 VSUBS 0.007897f
C987 B.n161 VSUBS 0.007897f
C988 B.n162 VSUBS 0.007432f
C989 B.n163 VSUBS 0.007897f
C990 B.n164 VSUBS 0.007897f
C991 B.n165 VSUBS 0.007897f
C992 B.n166 VSUBS 0.007897f
C993 B.n167 VSUBS 0.007897f
C994 B.t2 VSUBS 0.306542f
C995 B.t1 VSUBS 0.352557f
C996 B.t0 VSUBS 2.56104f
C997 B.n168 VSUBS 0.55955f
C998 B.n169 VSUBS 0.328155f
C999 B.n170 VSUBS 0.007897f
C1000 B.n171 VSUBS 0.007897f
C1001 B.n172 VSUBS 0.007897f
C1002 B.n173 VSUBS 0.007897f
C1003 B.n174 VSUBS 0.007897f
C1004 B.n175 VSUBS 0.007897f
C1005 B.n176 VSUBS 0.007897f
C1006 B.n177 VSUBS 0.007897f
C1007 B.n178 VSUBS 0.007897f
C1008 B.n179 VSUBS 0.007897f
C1009 B.n180 VSUBS 0.007897f
C1010 B.n181 VSUBS 0.007897f
C1011 B.n182 VSUBS 0.007897f
C1012 B.n183 VSUBS 0.007897f
C1013 B.n184 VSUBS 0.007897f
C1014 B.n185 VSUBS 0.007897f
C1015 B.n186 VSUBS 0.007897f
C1016 B.n187 VSUBS 0.007897f
C1017 B.n188 VSUBS 0.007897f
C1018 B.n189 VSUBS 0.007897f
C1019 B.n190 VSUBS 0.007897f
C1020 B.n191 VSUBS 0.007897f
C1021 B.n192 VSUBS 0.007897f
C1022 B.n193 VSUBS 0.007897f
C1023 B.n194 VSUBS 0.020056f
C1024 B.n195 VSUBS 0.007897f
C1025 B.n196 VSUBS 0.007897f
C1026 B.n197 VSUBS 0.007897f
C1027 B.n198 VSUBS 0.007897f
C1028 B.n199 VSUBS 0.007897f
C1029 B.n200 VSUBS 0.007897f
C1030 B.n201 VSUBS 0.007897f
C1031 B.n202 VSUBS 0.007897f
C1032 B.n203 VSUBS 0.007897f
C1033 B.n204 VSUBS 0.007897f
C1034 B.n205 VSUBS 0.007897f
C1035 B.n206 VSUBS 0.007897f
C1036 B.n207 VSUBS 0.007897f
C1037 B.n208 VSUBS 0.007897f
C1038 B.n209 VSUBS 0.007897f
C1039 B.n210 VSUBS 0.007897f
C1040 B.n211 VSUBS 0.007897f
C1041 B.n212 VSUBS 0.007897f
C1042 B.n213 VSUBS 0.007897f
C1043 B.n214 VSUBS 0.007897f
C1044 B.n215 VSUBS 0.007897f
C1045 B.n216 VSUBS 0.007897f
C1046 B.n217 VSUBS 0.007897f
C1047 B.n218 VSUBS 0.007897f
C1048 B.n219 VSUBS 0.007897f
C1049 B.n220 VSUBS 0.007897f
C1050 B.n221 VSUBS 0.007897f
C1051 B.n222 VSUBS 0.007897f
C1052 B.n223 VSUBS 0.007897f
C1053 B.n224 VSUBS 0.007897f
C1054 B.n225 VSUBS 0.007897f
C1055 B.n226 VSUBS 0.007897f
C1056 B.n227 VSUBS 0.007897f
C1057 B.n228 VSUBS 0.007897f
C1058 B.n229 VSUBS 0.007897f
C1059 B.n230 VSUBS 0.007897f
C1060 B.n231 VSUBS 0.007897f
C1061 B.n232 VSUBS 0.007897f
C1062 B.n233 VSUBS 0.007897f
C1063 B.n234 VSUBS 0.007897f
C1064 B.n235 VSUBS 0.007897f
C1065 B.n236 VSUBS 0.007897f
C1066 B.n237 VSUBS 0.007897f
C1067 B.n238 VSUBS 0.007897f
C1068 B.n239 VSUBS 0.007897f
C1069 B.n240 VSUBS 0.007897f
C1070 B.n241 VSUBS 0.007897f
C1071 B.n242 VSUBS 0.007897f
C1072 B.n243 VSUBS 0.007897f
C1073 B.n244 VSUBS 0.007897f
C1074 B.n245 VSUBS 0.007897f
C1075 B.n246 VSUBS 0.007897f
C1076 B.n247 VSUBS 0.007897f
C1077 B.n248 VSUBS 0.007897f
C1078 B.n249 VSUBS 0.007897f
C1079 B.n250 VSUBS 0.007897f
C1080 B.n251 VSUBS 0.007897f
C1081 B.n252 VSUBS 0.007897f
C1082 B.n253 VSUBS 0.007897f
C1083 B.n254 VSUBS 0.007897f
C1084 B.n255 VSUBS 0.007897f
C1085 B.n256 VSUBS 0.007897f
C1086 B.n257 VSUBS 0.007897f
C1087 B.n258 VSUBS 0.007897f
C1088 B.n259 VSUBS 0.007897f
C1089 B.n260 VSUBS 0.007897f
C1090 B.n261 VSUBS 0.007897f
C1091 B.n262 VSUBS 0.007897f
C1092 B.n263 VSUBS 0.007897f
C1093 B.n264 VSUBS 0.007897f
C1094 B.n265 VSUBS 0.007897f
C1095 B.n266 VSUBS 0.007897f
C1096 B.n267 VSUBS 0.007897f
C1097 B.n268 VSUBS 0.007897f
C1098 B.n269 VSUBS 0.007897f
C1099 B.n270 VSUBS 0.007897f
C1100 B.n271 VSUBS 0.007897f
C1101 B.n272 VSUBS 0.007897f
C1102 B.n273 VSUBS 0.007897f
C1103 B.n274 VSUBS 0.007897f
C1104 B.n275 VSUBS 0.007897f
C1105 B.n276 VSUBS 0.007897f
C1106 B.n277 VSUBS 0.007897f
C1107 B.n278 VSUBS 0.007897f
C1108 B.n279 VSUBS 0.007897f
C1109 B.n280 VSUBS 0.007897f
C1110 B.n281 VSUBS 0.007897f
C1111 B.n282 VSUBS 0.007897f
C1112 B.n283 VSUBS 0.007897f
C1113 B.n284 VSUBS 0.007897f
C1114 B.n285 VSUBS 0.007897f
C1115 B.n286 VSUBS 0.007897f
C1116 B.n287 VSUBS 0.007897f
C1117 B.n288 VSUBS 0.007897f
C1118 B.n289 VSUBS 0.007897f
C1119 B.n290 VSUBS 0.007897f
C1120 B.n291 VSUBS 0.007897f
C1121 B.n292 VSUBS 0.007897f
C1122 B.n293 VSUBS 0.020056f
C1123 B.n294 VSUBS 0.020821f
C1124 B.n295 VSUBS 0.020821f
C1125 B.n296 VSUBS 0.007897f
C1126 B.n297 VSUBS 0.007897f
C1127 B.n298 VSUBS 0.007897f
C1128 B.n299 VSUBS 0.007897f
C1129 B.n300 VSUBS 0.007897f
C1130 B.n301 VSUBS 0.007897f
C1131 B.n302 VSUBS 0.007897f
C1132 B.n303 VSUBS 0.007897f
C1133 B.n304 VSUBS 0.007897f
C1134 B.n305 VSUBS 0.007897f
C1135 B.n306 VSUBS 0.007897f
C1136 B.n307 VSUBS 0.007897f
C1137 B.n308 VSUBS 0.007897f
C1138 B.n309 VSUBS 0.007897f
C1139 B.n310 VSUBS 0.007897f
C1140 B.n311 VSUBS 0.007897f
C1141 B.n312 VSUBS 0.007897f
C1142 B.n313 VSUBS 0.007897f
C1143 B.n314 VSUBS 0.007897f
C1144 B.n315 VSUBS 0.007897f
C1145 B.n316 VSUBS 0.007897f
C1146 B.n317 VSUBS 0.007897f
C1147 B.n318 VSUBS 0.007897f
C1148 B.n319 VSUBS 0.007897f
C1149 B.n320 VSUBS 0.007897f
C1150 B.n321 VSUBS 0.007897f
C1151 B.n322 VSUBS 0.007897f
C1152 B.n323 VSUBS 0.007897f
C1153 B.n324 VSUBS 0.007897f
C1154 B.n325 VSUBS 0.007897f
C1155 B.n326 VSUBS 0.007897f
C1156 B.n327 VSUBS 0.007897f
C1157 B.n328 VSUBS 0.007897f
C1158 B.n329 VSUBS 0.007897f
C1159 B.n330 VSUBS 0.007897f
C1160 B.n331 VSUBS 0.007897f
C1161 B.n332 VSUBS 0.007897f
C1162 B.n333 VSUBS 0.007897f
C1163 B.n334 VSUBS 0.007897f
C1164 B.n335 VSUBS 0.007897f
C1165 B.n336 VSUBS 0.007897f
C1166 B.n337 VSUBS 0.007897f
C1167 B.n338 VSUBS 0.007897f
C1168 B.n339 VSUBS 0.007897f
C1169 B.n340 VSUBS 0.007897f
C1170 B.n341 VSUBS 0.007897f
C1171 B.n342 VSUBS 0.007897f
C1172 B.n343 VSUBS 0.007897f
C1173 B.n344 VSUBS 0.007897f
C1174 B.n345 VSUBS 0.007897f
C1175 B.n346 VSUBS 0.007897f
C1176 B.n347 VSUBS 0.007897f
C1177 B.n348 VSUBS 0.007897f
C1178 B.n349 VSUBS 0.007897f
C1179 B.n350 VSUBS 0.007897f
C1180 B.n351 VSUBS 0.007897f
C1181 B.n352 VSUBS 0.007897f
C1182 B.n353 VSUBS 0.007897f
C1183 B.n354 VSUBS 0.007897f
C1184 B.n355 VSUBS 0.007897f
C1185 B.n356 VSUBS 0.007897f
C1186 B.n357 VSUBS 0.007897f
C1187 B.n358 VSUBS 0.007897f
C1188 B.n359 VSUBS 0.007897f
C1189 B.n360 VSUBS 0.007897f
C1190 B.n361 VSUBS 0.007897f
C1191 B.n362 VSUBS 0.007897f
C1192 B.n363 VSUBS 0.007897f
C1193 B.n364 VSUBS 0.007897f
C1194 B.n365 VSUBS 0.007897f
C1195 B.n366 VSUBS 0.007897f
C1196 B.n367 VSUBS 0.007432f
C1197 B.n368 VSUBS 0.018296f
C1198 B.n369 VSUBS 0.004413f
C1199 B.n370 VSUBS 0.007897f
C1200 B.n371 VSUBS 0.007897f
C1201 B.n372 VSUBS 0.007897f
C1202 B.n373 VSUBS 0.007897f
C1203 B.n374 VSUBS 0.007897f
C1204 B.n375 VSUBS 0.007897f
C1205 B.n376 VSUBS 0.007897f
C1206 B.n377 VSUBS 0.007897f
C1207 B.n378 VSUBS 0.007897f
C1208 B.n379 VSUBS 0.007897f
C1209 B.n380 VSUBS 0.007897f
C1210 B.n381 VSUBS 0.007897f
C1211 B.t8 VSUBS 0.306545f
C1212 B.t7 VSUBS 0.352561f
C1213 B.t6 VSUBS 2.56104f
C1214 B.n382 VSUBS 0.559547f
C1215 B.n383 VSUBS 0.328152f
C1216 B.n384 VSUBS 0.018296f
C1217 B.n385 VSUBS 0.004413f
C1218 B.n386 VSUBS 0.007897f
C1219 B.n387 VSUBS 0.007897f
C1220 B.n388 VSUBS 0.007897f
C1221 B.n389 VSUBS 0.007897f
C1222 B.n390 VSUBS 0.007897f
C1223 B.n391 VSUBS 0.007897f
C1224 B.n392 VSUBS 0.007897f
C1225 B.n393 VSUBS 0.007897f
C1226 B.n394 VSUBS 0.007897f
C1227 B.n395 VSUBS 0.007897f
C1228 B.n396 VSUBS 0.007897f
C1229 B.n397 VSUBS 0.007897f
C1230 B.n398 VSUBS 0.007897f
C1231 B.n399 VSUBS 0.007897f
C1232 B.n400 VSUBS 0.007897f
C1233 B.n401 VSUBS 0.007897f
C1234 B.n402 VSUBS 0.007897f
C1235 B.n403 VSUBS 0.007897f
C1236 B.n404 VSUBS 0.007897f
C1237 B.n405 VSUBS 0.007897f
C1238 B.n406 VSUBS 0.007897f
C1239 B.n407 VSUBS 0.007897f
C1240 B.n408 VSUBS 0.007897f
C1241 B.n409 VSUBS 0.007897f
C1242 B.n410 VSUBS 0.007897f
C1243 B.n411 VSUBS 0.007897f
C1244 B.n412 VSUBS 0.007897f
C1245 B.n413 VSUBS 0.007897f
C1246 B.n414 VSUBS 0.007897f
C1247 B.n415 VSUBS 0.007897f
C1248 B.n416 VSUBS 0.007897f
C1249 B.n417 VSUBS 0.007897f
C1250 B.n418 VSUBS 0.007897f
C1251 B.n419 VSUBS 0.007897f
C1252 B.n420 VSUBS 0.007897f
C1253 B.n421 VSUBS 0.007897f
C1254 B.n422 VSUBS 0.007897f
C1255 B.n423 VSUBS 0.007897f
C1256 B.n424 VSUBS 0.007897f
C1257 B.n425 VSUBS 0.007897f
C1258 B.n426 VSUBS 0.007897f
C1259 B.n427 VSUBS 0.007897f
C1260 B.n428 VSUBS 0.007897f
C1261 B.n429 VSUBS 0.007897f
C1262 B.n430 VSUBS 0.007897f
C1263 B.n431 VSUBS 0.007897f
C1264 B.n432 VSUBS 0.007897f
C1265 B.n433 VSUBS 0.007897f
C1266 B.n434 VSUBS 0.007897f
C1267 B.n435 VSUBS 0.007897f
C1268 B.n436 VSUBS 0.007897f
C1269 B.n437 VSUBS 0.007897f
C1270 B.n438 VSUBS 0.007897f
C1271 B.n439 VSUBS 0.007897f
C1272 B.n440 VSUBS 0.007897f
C1273 B.n441 VSUBS 0.007897f
C1274 B.n442 VSUBS 0.007897f
C1275 B.n443 VSUBS 0.007897f
C1276 B.n444 VSUBS 0.007897f
C1277 B.n445 VSUBS 0.007897f
C1278 B.n446 VSUBS 0.007897f
C1279 B.n447 VSUBS 0.007897f
C1280 B.n448 VSUBS 0.007897f
C1281 B.n449 VSUBS 0.007897f
C1282 B.n450 VSUBS 0.007897f
C1283 B.n451 VSUBS 0.007897f
C1284 B.n452 VSUBS 0.007897f
C1285 B.n453 VSUBS 0.007897f
C1286 B.n454 VSUBS 0.007897f
C1287 B.n455 VSUBS 0.007897f
C1288 B.n456 VSUBS 0.007897f
C1289 B.n457 VSUBS 0.007897f
C1290 B.n458 VSUBS 0.007897f
C1291 B.n459 VSUBS 0.020821f
C1292 B.n460 VSUBS 0.020056f
C1293 B.n461 VSUBS 0.02086f
C1294 B.n462 VSUBS 0.007897f
C1295 B.n463 VSUBS 0.007897f
C1296 B.n464 VSUBS 0.007897f
C1297 B.n465 VSUBS 0.007897f
C1298 B.n466 VSUBS 0.007897f
C1299 B.n467 VSUBS 0.007897f
C1300 B.n468 VSUBS 0.007897f
C1301 B.n469 VSUBS 0.007897f
C1302 B.n470 VSUBS 0.007897f
C1303 B.n471 VSUBS 0.007897f
C1304 B.n472 VSUBS 0.007897f
C1305 B.n473 VSUBS 0.007897f
C1306 B.n474 VSUBS 0.007897f
C1307 B.n475 VSUBS 0.007897f
C1308 B.n476 VSUBS 0.007897f
C1309 B.n477 VSUBS 0.007897f
C1310 B.n478 VSUBS 0.007897f
C1311 B.n479 VSUBS 0.007897f
C1312 B.n480 VSUBS 0.007897f
C1313 B.n481 VSUBS 0.007897f
C1314 B.n482 VSUBS 0.007897f
C1315 B.n483 VSUBS 0.007897f
C1316 B.n484 VSUBS 0.007897f
C1317 B.n485 VSUBS 0.007897f
C1318 B.n486 VSUBS 0.007897f
C1319 B.n487 VSUBS 0.007897f
C1320 B.n488 VSUBS 0.007897f
C1321 B.n489 VSUBS 0.007897f
C1322 B.n490 VSUBS 0.007897f
C1323 B.n491 VSUBS 0.007897f
C1324 B.n492 VSUBS 0.007897f
C1325 B.n493 VSUBS 0.007897f
C1326 B.n494 VSUBS 0.007897f
C1327 B.n495 VSUBS 0.007897f
C1328 B.n496 VSUBS 0.007897f
C1329 B.n497 VSUBS 0.007897f
C1330 B.n498 VSUBS 0.007897f
C1331 B.n499 VSUBS 0.007897f
C1332 B.n500 VSUBS 0.007897f
C1333 B.n501 VSUBS 0.007897f
C1334 B.n502 VSUBS 0.007897f
C1335 B.n503 VSUBS 0.007897f
C1336 B.n504 VSUBS 0.007897f
C1337 B.n505 VSUBS 0.007897f
C1338 B.n506 VSUBS 0.007897f
C1339 B.n507 VSUBS 0.007897f
C1340 B.n508 VSUBS 0.007897f
C1341 B.n509 VSUBS 0.007897f
C1342 B.n510 VSUBS 0.007897f
C1343 B.n511 VSUBS 0.007897f
C1344 B.n512 VSUBS 0.007897f
C1345 B.n513 VSUBS 0.007897f
C1346 B.n514 VSUBS 0.007897f
C1347 B.n515 VSUBS 0.007897f
C1348 B.n516 VSUBS 0.007897f
C1349 B.n517 VSUBS 0.007897f
C1350 B.n518 VSUBS 0.007897f
C1351 B.n519 VSUBS 0.007897f
C1352 B.n520 VSUBS 0.007897f
C1353 B.n521 VSUBS 0.007897f
C1354 B.n522 VSUBS 0.007897f
C1355 B.n523 VSUBS 0.007897f
C1356 B.n524 VSUBS 0.007897f
C1357 B.n525 VSUBS 0.007897f
C1358 B.n526 VSUBS 0.007897f
C1359 B.n527 VSUBS 0.007897f
C1360 B.n528 VSUBS 0.007897f
C1361 B.n529 VSUBS 0.007897f
C1362 B.n530 VSUBS 0.007897f
C1363 B.n531 VSUBS 0.007897f
C1364 B.n532 VSUBS 0.007897f
C1365 B.n533 VSUBS 0.007897f
C1366 B.n534 VSUBS 0.007897f
C1367 B.n535 VSUBS 0.007897f
C1368 B.n536 VSUBS 0.007897f
C1369 B.n537 VSUBS 0.007897f
C1370 B.n538 VSUBS 0.007897f
C1371 B.n539 VSUBS 0.007897f
C1372 B.n540 VSUBS 0.007897f
C1373 B.n541 VSUBS 0.007897f
C1374 B.n542 VSUBS 0.007897f
C1375 B.n543 VSUBS 0.007897f
C1376 B.n544 VSUBS 0.007897f
C1377 B.n545 VSUBS 0.007897f
C1378 B.n546 VSUBS 0.007897f
C1379 B.n547 VSUBS 0.007897f
C1380 B.n548 VSUBS 0.007897f
C1381 B.n549 VSUBS 0.007897f
C1382 B.n550 VSUBS 0.007897f
C1383 B.n551 VSUBS 0.007897f
C1384 B.n552 VSUBS 0.007897f
C1385 B.n553 VSUBS 0.007897f
C1386 B.n554 VSUBS 0.007897f
C1387 B.n555 VSUBS 0.007897f
C1388 B.n556 VSUBS 0.007897f
C1389 B.n557 VSUBS 0.007897f
C1390 B.n558 VSUBS 0.007897f
C1391 B.n559 VSUBS 0.007897f
C1392 B.n560 VSUBS 0.007897f
C1393 B.n561 VSUBS 0.007897f
C1394 B.n562 VSUBS 0.007897f
C1395 B.n563 VSUBS 0.007897f
C1396 B.n564 VSUBS 0.007897f
C1397 B.n565 VSUBS 0.007897f
C1398 B.n566 VSUBS 0.007897f
C1399 B.n567 VSUBS 0.007897f
C1400 B.n568 VSUBS 0.007897f
C1401 B.n569 VSUBS 0.007897f
C1402 B.n570 VSUBS 0.007897f
C1403 B.n571 VSUBS 0.007897f
C1404 B.n572 VSUBS 0.007897f
C1405 B.n573 VSUBS 0.007897f
C1406 B.n574 VSUBS 0.007897f
C1407 B.n575 VSUBS 0.007897f
C1408 B.n576 VSUBS 0.007897f
C1409 B.n577 VSUBS 0.007897f
C1410 B.n578 VSUBS 0.007897f
C1411 B.n579 VSUBS 0.007897f
C1412 B.n580 VSUBS 0.007897f
C1413 B.n581 VSUBS 0.007897f
C1414 B.n582 VSUBS 0.007897f
C1415 B.n583 VSUBS 0.007897f
C1416 B.n584 VSUBS 0.007897f
C1417 B.n585 VSUBS 0.007897f
C1418 B.n586 VSUBS 0.007897f
C1419 B.n587 VSUBS 0.007897f
C1420 B.n588 VSUBS 0.007897f
C1421 B.n589 VSUBS 0.007897f
C1422 B.n590 VSUBS 0.007897f
C1423 B.n591 VSUBS 0.007897f
C1424 B.n592 VSUBS 0.007897f
C1425 B.n593 VSUBS 0.007897f
C1426 B.n594 VSUBS 0.007897f
C1427 B.n595 VSUBS 0.007897f
C1428 B.n596 VSUBS 0.007897f
C1429 B.n597 VSUBS 0.007897f
C1430 B.n598 VSUBS 0.007897f
C1431 B.n599 VSUBS 0.007897f
C1432 B.n600 VSUBS 0.007897f
C1433 B.n601 VSUBS 0.007897f
C1434 B.n602 VSUBS 0.007897f
C1435 B.n603 VSUBS 0.007897f
C1436 B.n604 VSUBS 0.007897f
C1437 B.n605 VSUBS 0.007897f
C1438 B.n606 VSUBS 0.007897f
C1439 B.n607 VSUBS 0.007897f
C1440 B.n608 VSUBS 0.007897f
C1441 B.n609 VSUBS 0.007897f
C1442 B.n610 VSUBS 0.007897f
C1443 B.n611 VSUBS 0.007897f
C1444 B.n612 VSUBS 0.007897f
C1445 B.n613 VSUBS 0.007897f
C1446 B.n614 VSUBS 0.007897f
C1447 B.n615 VSUBS 0.020056f
C1448 B.n616 VSUBS 0.020821f
C1449 B.n617 VSUBS 0.020821f
C1450 B.n618 VSUBS 0.007897f
C1451 B.n619 VSUBS 0.007897f
C1452 B.n620 VSUBS 0.007897f
C1453 B.n621 VSUBS 0.007897f
C1454 B.n622 VSUBS 0.007897f
C1455 B.n623 VSUBS 0.007897f
C1456 B.n624 VSUBS 0.007897f
C1457 B.n625 VSUBS 0.007897f
C1458 B.n626 VSUBS 0.007897f
C1459 B.n627 VSUBS 0.007897f
C1460 B.n628 VSUBS 0.007897f
C1461 B.n629 VSUBS 0.007897f
C1462 B.n630 VSUBS 0.007897f
C1463 B.n631 VSUBS 0.007897f
C1464 B.n632 VSUBS 0.007897f
C1465 B.n633 VSUBS 0.007897f
C1466 B.n634 VSUBS 0.007897f
C1467 B.n635 VSUBS 0.007897f
C1468 B.n636 VSUBS 0.007897f
C1469 B.n637 VSUBS 0.007897f
C1470 B.n638 VSUBS 0.007897f
C1471 B.n639 VSUBS 0.007897f
C1472 B.n640 VSUBS 0.007897f
C1473 B.n641 VSUBS 0.007897f
C1474 B.n642 VSUBS 0.007897f
C1475 B.n643 VSUBS 0.007897f
C1476 B.n644 VSUBS 0.007897f
C1477 B.n645 VSUBS 0.007897f
C1478 B.n646 VSUBS 0.007897f
C1479 B.n647 VSUBS 0.007897f
C1480 B.n648 VSUBS 0.007897f
C1481 B.n649 VSUBS 0.007897f
C1482 B.n650 VSUBS 0.007897f
C1483 B.n651 VSUBS 0.007897f
C1484 B.n652 VSUBS 0.007897f
C1485 B.n653 VSUBS 0.007897f
C1486 B.n654 VSUBS 0.007897f
C1487 B.n655 VSUBS 0.007897f
C1488 B.n656 VSUBS 0.007897f
C1489 B.n657 VSUBS 0.007897f
C1490 B.n658 VSUBS 0.007897f
C1491 B.n659 VSUBS 0.007897f
C1492 B.n660 VSUBS 0.007897f
C1493 B.n661 VSUBS 0.007897f
C1494 B.n662 VSUBS 0.007897f
C1495 B.n663 VSUBS 0.007897f
C1496 B.n664 VSUBS 0.007897f
C1497 B.n665 VSUBS 0.007897f
C1498 B.n666 VSUBS 0.007897f
C1499 B.n667 VSUBS 0.007897f
C1500 B.n668 VSUBS 0.007897f
C1501 B.n669 VSUBS 0.007897f
C1502 B.n670 VSUBS 0.007897f
C1503 B.n671 VSUBS 0.007897f
C1504 B.n672 VSUBS 0.007897f
C1505 B.n673 VSUBS 0.007897f
C1506 B.n674 VSUBS 0.007897f
C1507 B.n675 VSUBS 0.007897f
C1508 B.n676 VSUBS 0.007897f
C1509 B.n677 VSUBS 0.007897f
C1510 B.n678 VSUBS 0.007897f
C1511 B.n679 VSUBS 0.007897f
C1512 B.n680 VSUBS 0.007897f
C1513 B.n681 VSUBS 0.007897f
C1514 B.n682 VSUBS 0.007897f
C1515 B.n683 VSUBS 0.007897f
C1516 B.n684 VSUBS 0.007897f
C1517 B.n685 VSUBS 0.007897f
C1518 B.n686 VSUBS 0.007897f
C1519 B.n687 VSUBS 0.007897f
C1520 B.n688 VSUBS 0.007897f
C1521 B.n689 VSUBS 0.007432f
C1522 B.n690 VSUBS 0.018296f
C1523 B.n691 VSUBS 0.004413f
C1524 B.n692 VSUBS 0.007897f
C1525 B.n693 VSUBS 0.007897f
C1526 B.n694 VSUBS 0.007897f
C1527 B.n695 VSUBS 0.007897f
C1528 B.n696 VSUBS 0.007897f
C1529 B.n697 VSUBS 0.007897f
C1530 B.n698 VSUBS 0.007897f
C1531 B.n699 VSUBS 0.007897f
C1532 B.n700 VSUBS 0.007897f
C1533 B.n701 VSUBS 0.007897f
C1534 B.n702 VSUBS 0.007897f
C1535 B.n703 VSUBS 0.007897f
C1536 B.n704 VSUBS 0.004413f
C1537 B.n705 VSUBS 0.007897f
C1538 B.n706 VSUBS 0.007897f
C1539 B.n707 VSUBS 0.007432f
C1540 B.n708 VSUBS 0.007897f
C1541 B.n709 VSUBS 0.007897f
C1542 B.n710 VSUBS 0.007897f
C1543 B.n711 VSUBS 0.007897f
C1544 B.n712 VSUBS 0.007897f
C1545 B.n713 VSUBS 0.007897f
C1546 B.n714 VSUBS 0.007897f
C1547 B.n715 VSUBS 0.007897f
C1548 B.n716 VSUBS 0.007897f
C1549 B.n717 VSUBS 0.007897f
C1550 B.n718 VSUBS 0.007897f
C1551 B.n719 VSUBS 0.007897f
C1552 B.n720 VSUBS 0.007897f
C1553 B.n721 VSUBS 0.007897f
C1554 B.n722 VSUBS 0.007897f
C1555 B.n723 VSUBS 0.007897f
C1556 B.n724 VSUBS 0.007897f
C1557 B.n725 VSUBS 0.007897f
C1558 B.n726 VSUBS 0.007897f
C1559 B.n727 VSUBS 0.007897f
C1560 B.n728 VSUBS 0.007897f
C1561 B.n729 VSUBS 0.007897f
C1562 B.n730 VSUBS 0.007897f
C1563 B.n731 VSUBS 0.007897f
C1564 B.n732 VSUBS 0.007897f
C1565 B.n733 VSUBS 0.007897f
C1566 B.n734 VSUBS 0.007897f
C1567 B.n735 VSUBS 0.007897f
C1568 B.n736 VSUBS 0.007897f
C1569 B.n737 VSUBS 0.007897f
C1570 B.n738 VSUBS 0.007897f
C1571 B.n739 VSUBS 0.007897f
C1572 B.n740 VSUBS 0.007897f
C1573 B.n741 VSUBS 0.007897f
C1574 B.n742 VSUBS 0.007897f
C1575 B.n743 VSUBS 0.007897f
C1576 B.n744 VSUBS 0.007897f
C1577 B.n745 VSUBS 0.007897f
C1578 B.n746 VSUBS 0.007897f
C1579 B.n747 VSUBS 0.007897f
C1580 B.n748 VSUBS 0.007897f
C1581 B.n749 VSUBS 0.007897f
C1582 B.n750 VSUBS 0.007897f
C1583 B.n751 VSUBS 0.007897f
C1584 B.n752 VSUBS 0.007897f
C1585 B.n753 VSUBS 0.007897f
C1586 B.n754 VSUBS 0.007897f
C1587 B.n755 VSUBS 0.007897f
C1588 B.n756 VSUBS 0.007897f
C1589 B.n757 VSUBS 0.007897f
C1590 B.n758 VSUBS 0.007897f
C1591 B.n759 VSUBS 0.007897f
C1592 B.n760 VSUBS 0.007897f
C1593 B.n761 VSUBS 0.007897f
C1594 B.n762 VSUBS 0.007897f
C1595 B.n763 VSUBS 0.007897f
C1596 B.n764 VSUBS 0.007897f
C1597 B.n765 VSUBS 0.007897f
C1598 B.n766 VSUBS 0.007897f
C1599 B.n767 VSUBS 0.007897f
C1600 B.n768 VSUBS 0.007897f
C1601 B.n769 VSUBS 0.007897f
C1602 B.n770 VSUBS 0.007897f
C1603 B.n771 VSUBS 0.007897f
C1604 B.n772 VSUBS 0.007897f
C1605 B.n773 VSUBS 0.007897f
C1606 B.n774 VSUBS 0.007897f
C1607 B.n775 VSUBS 0.007897f
C1608 B.n776 VSUBS 0.007897f
C1609 B.n777 VSUBS 0.007897f
C1610 B.n778 VSUBS 0.020821f
C1611 B.n779 VSUBS 0.020821f
C1612 B.n780 VSUBS 0.020056f
C1613 B.n781 VSUBS 0.007897f
C1614 B.n782 VSUBS 0.007897f
C1615 B.n783 VSUBS 0.007897f
C1616 B.n784 VSUBS 0.007897f
C1617 B.n785 VSUBS 0.007897f
C1618 B.n786 VSUBS 0.007897f
C1619 B.n787 VSUBS 0.007897f
C1620 B.n788 VSUBS 0.007897f
C1621 B.n789 VSUBS 0.007897f
C1622 B.n790 VSUBS 0.007897f
C1623 B.n791 VSUBS 0.007897f
C1624 B.n792 VSUBS 0.007897f
C1625 B.n793 VSUBS 0.007897f
C1626 B.n794 VSUBS 0.007897f
C1627 B.n795 VSUBS 0.007897f
C1628 B.n796 VSUBS 0.007897f
C1629 B.n797 VSUBS 0.007897f
C1630 B.n798 VSUBS 0.007897f
C1631 B.n799 VSUBS 0.007897f
C1632 B.n800 VSUBS 0.007897f
C1633 B.n801 VSUBS 0.007897f
C1634 B.n802 VSUBS 0.007897f
C1635 B.n803 VSUBS 0.007897f
C1636 B.n804 VSUBS 0.007897f
C1637 B.n805 VSUBS 0.007897f
C1638 B.n806 VSUBS 0.007897f
C1639 B.n807 VSUBS 0.007897f
C1640 B.n808 VSUBS 0.007897f
C1641 B.n809 VSUBS 0.007897f
C1642 B.n810 VSUBS 0.007897f
C1643 B.n811 VSUBS 0.007897f
C1644 B.n812 VSUBS 0.007897f
C1645 B.n813 VSUBS 0.007897f
C1646 B.n814 VSUBS 0.007897f
C1647 B.n815 VSUBS 0.007897f
C1648 B.n816 VSUBS 0.007897f
C1649 B.n817 VSUBS 0.007897f
C1650 B.n818 VSUBS 0.007897f
C1651 B.n819 VSUBS 0.007897f
C1652 B.n820 VSUBS 0.007897f
C1653 B.n821 VSUBS 0.007897f
C1654 B.n822 VSUBS 0.007897f
C1655 B.n823 VSUBS 0.007897f
C1656 B.n824 VSUBS 0.007897f
C1657 B.n825 VSUBS 0.007897f
C1658 B.n826 VSUBS 0.007897f
C1659 B.n827 VSUBS 0.007897f
C1660 B.n828 VSUBS 0.007897f
C1661 B.n829 VSUBS 0.007897f
C1662 B.n830 VSUBS 0.007897f
C1663 B.n831 VSUBS 0.007897f
C1664 B.n832 VSUBS 0.007897f
C1665 B.n833 VSUBS 0.007897f
C1666 B.n834 VSUBS 0.007897f
C1667 B.n835 VSUBS 0.007897f
C1668 B.n836 VSUBS 0.007897f
C1669 B.n837 VSUBS 0.007897f
C1670 B.n838 VSUBS 0.007897f
C1671 B.n839 VSUBS 0.007897f
C1672 B.n840 VSUBS 0.007897f
C1673 B.n841 VSUBS 0.007897f
C1674 B.n842 VSUBS 0.007897f
C1675 B.n843 VSUBS 0.007897f
C1676 B.n844 VSUBS 0.007897f
C1677 B.n845 VSUBS 0.007897f
C1678 B.n846 VSUBS 0.007897f
C1679 B.n847 VSUBS 0.007897f
C1680 B.n848 VSUBS 0.007897f
C1681 B.n849 VSUBS 0.007897f
C1682 B.n850 VSUBS 0.007897f
C1683 B.n851 VSUBS 0.007897f
C1684 B.n852 VSUBS 0.007897f
C1685 B.n853 VSUBS 0.007897f
C1686 B.n854 VSUBS 0.007897f
C1687 B.n855 VSUBS 0.010305f
C1688 B.n856 VSUBS 0.010977f
C1689 B.n857 VSUBS 0.021829f
.ends

