* NGSPICE file created from diff_pair_sample_0954.ext - technology: sky130A

.subckt diff_pair_sample_0954 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t4 w_n4700_n3166# sky130_fd_pr__pfet_01v8 ad=1.81335 pd=11.32 as=1.81335 ps=11.32 w=10.99 l=3.4
X1 VDD1.t6 VP.t1 VTAIL.t14 w_n4700_n3166# sky130_fd_pr__pfet_01v8 ad=1.81335 pd=11.32 as=4.2861 ps=22.76 w=10.99 l=3.4
X2 VTAIL.t0 VN.t0 VDD2.t7 w_n4700_n3166# sky130_fd_pr__pfet_01v8 ad=4.2861 pd=22.76 as=1.81335 ps=11.32 w=10.99 l=3.4
X3 VDD2.t6 VN.t1 VTAIL.t3 w_n4700_n3166# sky130_fd_pr__pfet_01v8 ad=1.81335 pd=11.32 as=1.81335 ps=11.32 w=10.99 l=3.4
X4 VTAIL.t1 VN.t2 VDD2.t5 w_n4700_n3166# sky130_fd_pr__pfet_01v8 ad=1.81335 pd=11.32 as=1.81335 ps=11.32 w=10.99 l=3.4
X5 VDD2.t4 VN.t3 VTAIL.t5 w_n4700_n3166# sky130_fd_pr__pfet_01v8 ad=1.81335 pd=11.32 as=4.2861 ps=22.76 w=10.99 l=3.4
X6 VDD2.t3 VN.t4 VTAIL.t7 w_n4700_n3166# sky130_fd_pr__pfet_01v8 ad=1.81335 pd=11.32 as=4.2861 ps=22.76 w=10.99 l=3.4
X7 VTAIL.t13 VP.t2 VDD1.t1 w_n4700_n3166# sky130_fd_pr__pfet_01v8 ad=1.81335 pd=11.32 as=1.81335 ps=11.32 w=10.99 l=3.4
X8 VDD1.t5 VP.t3 VTAIL.t12 w_n4700_n3166# sky130_fd_pr__pfet_01v8 ad=1.81335 pd=11.32 as=1.81335 ps=11.32 w=10.99 l=3.4
X9 VDD1.t0 VP.t4 VTAIL.t11 w_n4700_n3166# sky130_fd_pr__pfet_01v8 ad=1.81335 pd=11.32 as=4.2861 ps=22.76 w=10.99 l=3.4
X10 VDD2.t2 VN.t5 VTAIL.t6 w_n4700_n3166# sky130_fd_pr__pfet_01v8 ad=1.81335 pd=11.32 as=1.81335 ps=11.32 w=10.99 l=3.4
X11 B.t11 B.t9 B.t10 w_n4700_n3166# sky130_fd_pr__pfet_01v8 ad=4.2861 pd=22.76 as=0 ps=0 w=10.99 l=3.4
X12 B.t8 B.t6 B.t7 w_n4700_n3166# sky130_fd_pr__pfet_01v8 ad=4.2861 pd=22.76 as=0 ps=0 w=10.99 l=3.4
X13 VDD1.t7 VP.t5 VTAIL.t10 w_n4700_n3166# sky130_fd_pr__pfet_01v8 ad=1.81335 pd=11.32 as=1.81335 ps=11.32 w=10.99 l=3.4
X14 VTAIL.t9 VP.t6 VDD1.t2 w_n4700_n3166# sky130_fd_pr__pfet_01v8 ad=4.2861 pd=22.76 as=1.81335 ps=11.32 w=10.99 l=3.4
X15 VTAIL.t2 VN.t6 VDD2.t1 w_n4700_n3166# sky130_fd_pr__pfet_01v8 ad=4.2861 pd=22.76 as=1.81335 ps=11.32 w=10.99 l=3.4
X16 B.t5 B.t3 B.t4 w_n4700_n3166# sky130_fd_pr__pfet_01v8 ad=4.2861 pd=22.76 as=0 ps=0 w=10.99 l=3.4
X17 B.t2 B.t0 B.t1 w_n4700_n3166# sky130_fd_pr__pfet_01v8 ad=4.2861 pd=22.76 as=0 ps=0 w=10.99 l=3.4
X18 VTAIL.t4 VN.t7 VDD2.t0 w_n4700_n3166# sky130_fd_pr__pfet_01v8 ad=1.81335 pd=11.32 as=1.81335 ps=11.32 w=10.99 l=3.4
X19 VTAIL.t8 VP.t7 VDD1.t3 w_n4700_n3166# sky130_fd_pr__pfet_01v8 ad=4.2861 pd=22.76 as=1.81335 ps=11.32 w=10.99 l=3.4
R0 VP.n24 VP.n21 161.3
R1 VP.n26 VP.n25 161.3
R2 VP.n27 VP.n20 161.3
R3 VP.n29 VP.n28 161.3
R4 VP.n30 VP.n19 161.3
R5 VP.n32 VP.n31 161.3
R6 VP.n33 VP.n18 161.3
R7 VP.n35 VP.n34 161.3
R8 VP.n37 VP.n36 161.3
R9 VP.n38 VP.n16 161.3
R10 VP.n40 VP.n39 161.3
R11 VP.n41 VP.n15 161.3
R12 VP.n43 VP.n42 161.3
R13 VP.n44 VP.n14 161.3
R14 VP.n46 VP.n45 161.3
R15 VP.n83 VP.n82 161.3
R16 VP.n81 VP.n1 161.3
R17 VP.n80 VP.n79 161.3
R18 VP.n78 VP.n2 161.3
R19 VP.n77 VP.n76 161.3
R20 VP.n75 VP.n3 161.3
R21 VP.n74 VP.n73 161.3
R22 VP.n72 VP.n71 161.3
R23 VP.n70 VP.n5 161.3
R24 VP.n69 VP.n68 161.3
R25 VP.n67 VP.n6 161.3
R26 VP.n66 VP.n65 161.3
R27 VP.n64 VP.n7 161.3
R28 VP.n63 VP.n62 161.3
R29 VP.n61 VP.n8 161.3
R30 VP.n60 VP.n59 161.3
R31 VP.n57 VP.n9 161.3
R32 VP.n56 VP.n55 161.3
R33 VP.n54 VP.n10 161.3
R34 VP.n53 VP.n52 161.3
R35 VP.n51 VP.n11 161.3
R36 VP.n50 VP.n49 161.3
R37 VP.n23 VP.t6 110.983
R38 VP.n12 VP.t7 77.9002
R39 VP.n58 VP.t5 77.9002
R40 VP.n4 VP.t0 77.9002
R41 VP.n0 VP.t4 77.9002
R42 VP.n13 VP.t1 77.9002
R43 VP.n17 VP.t2 77.9002
R44 VP.n22 VP.t3 77.9002
R45 VP.n48 VP.n12 73.1852
R46 VP.n84 VP.n0 73.1852
R47 VP.n47 VP.n13 73.1852
R48 VP.n23 VP.n22 68.9427
R49 VP.n65 VP.n6 56.5193
R50 VP.n28 VP.n19 56.5193
R51 VP.n48 VP.n47 54.0448
R52 VP.n56 VP.n10 42.4359
R53 VP.n76 VP.n2 42.4359
R54 VP.n39 VP.n15 42.4359
R55 VP.n52 VP.n10 38.5509
R56 VP.n80 VP.n2 38.5509
R57 VP.n43 VP.n15 38.5509
R58 VP.n51 VP.n50 24.4675
R59 VP.n52 VP.n51 24.4675
R60 VP.n57 VP.n56 24.4675
R61 VP.n59 VP.n57 24.4675
R62 VP.n63 VP.n8 24.4675
R63 VP.n64 VP.n63 24.4675
R64 VP.n65 VP.n64 24.4675
R65 VP.n69 VP.n6 24.4675
R66 VP.n70 VP.n69 24.4675
R67 VP.n71 VP.n70 24.4675
R68 VP.n75 VP.n74 24.4675
R69 VP.n76 VP.n75 24.4675
R70 VP.n81 VP.n80 24.4675
R71 VP.n82 VP.n81 24.4675
R72 VP.n44 VP.n43 24.4675
R73 VP.n45 VP.n44 24.4675
R74 VP.n32 VP.n19 24.4675
R75 VP.n33 VP.n32 24.4675
R76 VP.n34 VP.n33 24.4675
R77 VP.n38 VP.n37 24.4675
R78 VP.n39 VP.n38 24.4675
R79 VP.n26 VP.n21 24.4675
R80 VP.n27 VP.n26 24.4675
R81 VP.n28 VP.n27 24.4675
R82 VP.n59 VP.n58 18.8401
R83 VP.n74 VP.n4 18.8401
R84 VP.n37 VP.n17 18.8401
R85 VP.n50 VP.n12 16.8827
R86 VP.n82 VP.n0 16.8827
R87 VP.n45 VP.n13 16.8827
R88 VP.n58 VP.n8 5.62791
R89 VP.n71 VP.n4 5.62791
R90 VP.n34 VP.n17 5.62791
R91 VP.n22 VP.n21 5.62791
R92 VP.n24 VP.n23 4.05577
R93 VP.n47 VP.n46 0.354971
R94 VP.n49 VP.n48 0.354971
R95 VP.n84 VP.n83 0.354971
R96 VP VP.n84 0.26696
R97 VP.n25 VP.n24 0.189894
R98 VP.n25 VP.n20 0.189894
R99 VP.n29 VP.n20 0.189894
R100 VP.n30 VP.n29 0.189894
R101 VP.n31 VP.n30 0.189894
R102 VP.n31 VP.n18 0.189894
R103 VP.n35 VP.n18 0.189894
R104 VP.n36 VP.n35 0.189894
R105 VP.n36 VP.n16 0.189894
R106 VP.n40 VP.n16 0.189894
R107 VP.n41 VP.n40 0.189894
R108 VP.n42 VP.n41 0.189894
R109 VP.n42 VP.n14 0.189894
R110 VP.n46 VP.n14 0.189894
R111 VP.n49 VP.n11 0.189894
R112 VP.n53 VP.n11 0.189894
R113 VP.n54 VP.n53 0.189894
R114 VP.n55 VP.n54 0.189894
R115 VP.n55 VP.n9 0.189894
R116 VP.n60 VP.n9 0.189894
R117 VP.n61 VP.n60 0.189894
R118 VP.n62 VP.n61 0.189894
R119 VP.n62 VP.n7 0.189894
R120 VP.n66 VP.n7 0.189894
R121 VP.n67 VP.n66 0.189894
R122 VP.n68 VP.n67 0.189894
R123 VP.n68 VP.n5 0.189894
R124 VP.n72 VP.n5 0.189894
R125 VP.n73 VP.n72 0.189894
R126 VP.n73 VP.n3 0.189894
R127 VP.n77 VP.n3 0.189894
R128 VP.n78 VP.n77 0.189894
R129 VP.n79 VP.n78 0.189894
R130 VP.n79 VP.n1 0.189894
R131 VP.n83 VP.n1 0.189894
R132 VDD1 VDD1.n0 76.0013
R133 VDD1.n3 VDD1.n2 75.8875
R134 VDD1.n3 VDD1.n1 75.8875
R135 VDD1.n5 VDD1.n4 74.3352
R136 VDD1.n5 VDD1.n3 48.2423
R137 VDD1.n4 VDD1.t1 2.95819
R138 VDD1.n4 VDD1.t6 2.95819
R139 VDD1.n0 VDD1.t2 2.95819
R140 VDD1.n0 VDD1.t5 2.95819
R141 VDD1.n2 VDD1.t4 2.95819
R142 VDD1.n2 VDD1.t0 2.95819
R143 VDD1.n1 VDD1.t3 2.95819
R144 VDD1.n1 VDD1.t7 2.95819
R145 VDD1 VDD1.n5 1.55007
R146 VTAIL.n11 VTAIL.t9 60.6142
R147 VTAIL.n10 VTAIL.t7 60.6142
R148 VTAIL.n7 VTAIL.t0 60.6142
R149 VTAIL.n15 VTAIL.t5 60.6141
R150 VTAIL.n2 VTAIL.t2 60.6141
R151 VTAIL.n3 VTAIL.t11 60.6141
R152 VTAIL.n6 VTAIL.t8 60.6141
R153 VTAIL.n14 VTAIL.t14 60.6141
R154 VTAIL.n13 VTAIL.n12 57.6566
R155 VTAIL.n9 VTAIL.n8 57.6566
R156 VTAIL.n1 VTAIL.n0 57.6563
R157 VTAIL.n5 VTAIL.n4 57.6563
R158 VTAIL.n15 VTAIL.n14 25.0565
R159 VTAIL.n7 VTAIL.n6 25.0565
R160 VTAIL.n9 VTAIL.n7 3.21602
R161 VTAIL.n10 VTAIL.n9 3.21602
R162 VTAIL.n13 VTAIL.n11 3.21602
R163 VTAIL.n14 VTAIL.n13 3.21602
R164 VTAIL.n6 VTAIL.n5 3.21602
R165 VTAIL.n5 VTAIL.n3 3.21602
R166 VTAIL.n2 VTAIL.n1 3.21602
R167 VTAIL VTAIL.n15 3.15783
R168 VTAIL.n0 VTAIL.t3 2.95819
R169 VTAIL.n0 VTAIL.t4 2.95819
R170 VTAIL.n4 VTAIL.t10 2.95819
R171 VTAIL.n4 VTAIL.t15 2.95819
R172 VTAIL.n12 VTAIL.t12 2.95819
R173 VTAIL.n12 VTAIL.t13 2.95819
R174 VTAIL.n8 VTAIL.t6 2.95819
R175 VTAIL.n8 VTAIL.t1 2.95819
R176 VTAIL.n11 VTAIL.n10 0.470328
R177 VTAIL.n3 VTAIL.n2 0.470328
R178 VTAIL VTAIL.n1 0.0586897
R179 VN.n68 VN.n67 161.3
R180 VN.n66 VN.n36 161.3
R181 VN.n65 VN.n64 161.3
R182 VN.n63 VN.n37 161.3
R183 VN.n62 VN.n61 161.3
R184 VN.n60 VN.n38 161.3
R185 VN.n59 VN.n58 161.3
R186 VN.n57 VN.n56 161.3
R187 VN.n55 VN.n40 161.3
R188 VN.n54 VN.n53 161.3
R189 VN.n52 VN.n41 161.3
R190 VN.n51 VN.n50 161.3
R191 VN.n49 VN.n42 161.3
R192 VN.n48 VN.n47 161.3
R193 VN.n46 VN.n43 161.3
R194 VN.n33 VN.n32 161.3
R195 VN.n31 VN.n1 161.3
R196 VN.n30 VN.n29 161.3
R197 VN.n28 VN.n2 161.3
R198 VN.n27 VN.n26 161.3
R199 VN.n25 VN.n3 161.3
R200 VN.n24 VN.n23 161.3
R201 VN.n22 VN.n21 161.3
R202 VN.n20 VN.n5 161.3
R203 VN.n19 VN.n18 161.3
R204 VN.n17 VN.n6 161.3
R205 VN.n16 VN.n15 161.3
R206 VN.n14 VN.n7 161.3
R207 VN.n13 VN.n12 161.3
R208 VN.n11 VN.n8 161.3
R209 VN.n45 VN.t4 110.984
R210 VN.n10 VN.t6 110.984
R211 VN.n9 VN.t1 77.9002
R212 VN.n4 VN.t7 77.9002
R213 VN.n0 VN.t3 77.9002
R214 VN.n44 VN.t2 77.9002
R215 VN.n39 VN.t5 77.9002
R216 VN.n35 VN.t0 77.9002
R217 VN.n34 VN.n0 73.1852
R218 VN.n69 VN.n35 73.1852
R219 VN.n10 VN.n9 68.9426
R220 VN.n45 VN.n44 68.9426
R221 VN.n15 VN.n6 56.5193
R222 VN.n50 VN.n41 56.5193
R223 VN VN.n69 54.2101
R224 VN.n26 VN.n2 42.4359
R225 VN.n61 VN.n37 42.4359
R226 VN.n30 VN.n2 38.5509
R227 VN.n65 VN.n37 38.5509
R228 VN.n13 VN.n8 24.4675
R229 VN.n14 VN.n13 24.4675
R230 VN.n15 VN.n14 24.4675
R231 VN.n19 VN.n6 24.4675
R232 VN.n20 VN.n19 24.4675
R233 VN.n21 VN.n20 24.4675
R234 VN.n25 VN.n24 24.4675
R235 VN.n26 VN.n25 24.4675
R236 VN.n31 VN.n30 24.4675
R237 VN.n32 VN.n31 24.4675
R238 VN.n50 VN.n49 24.4675
R239 VN.n49 VN.n48 24.4675
R240 VN.n48 VN.n43 24.4675
R241 VN.n61 VN.n60 24.4675
R242 VN.n60 VN.n59 24.4675
R243 VN.n56 VN.n55 24.4675
R244 VN.n55 VN.n54 24.4675
R245 VN.n54 VN.n41 24.4675
R246 VN.n67 VN.n66 24.4675
R247 VN.n66 VN.n65 24.4675
R248 VN.n24 VN.n4 18.8401
R249 VN.n59 VN.n39 18.8401
R250 VN.n32 VN.n0 16.8827
R251 VN.n67 VN.n35 16.8827
R252 VN.n9 VN.n8 5.62791
R253 VN.n21 VN.n4 5.62791
R254 VN.n44 VN.n43 5.62791
R255 VN.n56 VN.n39 5.62791
R256 VN.n11 VN.n10 4.0558
R257 VN.n46 VN.n45 4.05579
R258 VN.n69 VN.n68 0.354971
R259 VN.n34 VN.n33 0.354971
R260 VN VN.n34 0.26696
R261 VN.n68 VN.n36 0.189894
R262 VN.n64 VN.n36 0.189894
R263 VN.n64 VN.n63 0.189894
R264 VN.n63 VN.n62 0.189894
R265 VN.n62 VN.n38 0.189894
R266 VN.n58 VN.n38 0.189894
R267 VN.n58 VN.n57 0.189894
R268 VN.n57 VN.n40 0.189894
R269 VN.n53 VN.n40 0.189894
R270 VN.n53 VN.n52 0.189894
R271 VN.n52 VN.n51 0.189894
R272 VN.n51 VN.n42 0.189894
R273 VN.n47 VN.n42 0.189894
R274 VN.n47 VN.n46 0.189894
R275 VN.n12 VN.n11 0.189894
R276 VN.n12 VN.n7 0.189894
R277 VN.n16 VN.n7 0.189894
R278 VN.n17 VN.n16 0.189894
R279 VN.n18 VN.n17 0.189894
R280 VN.n18 VN.n5 0.189894
R281 VN.n22 VN.n5 0.189894
R282 VN.n23 VN.n22 0.189894
R283 VN.n23 VN.n3 0.189894
R284 VN.n27 VN.n3 0.189894
R285 VN.n28 VN.n27 0.189894
R286 VN.n29 VN.n28 0.189894
R287 VN.n29 VN.n1 0.189894
R288 VN.n33 VN.n1 0.189894
R289 VDD2.n2 VDD2.n1 75.8875
R290 VDD2.n2 VDD2.n0 75.8875
R291 VDD2 VDD2.n5 75.8847
R292 VDD2.n4 VDD2.n3 74.3354
R293 VDD2.n4 VDD2.n2 47.6593
R294 VDD2.n5 VDD2.t5 2.95819
R295 VDD2.n5 VDD2.t3 2.95819
R296 VDD2.n3 VDD2.t7 2.95819
R297 VDD2.n3 VDD2.t2 2.95819
R298 VDD2.n1 VDD2.t0 2.95819
R299 VDD2.n1 VDD2.t4 2.95819
R300 VDD2.n0 VDD2.t1 2.95819
R301 VDD2.n0 VDD2.t6 2.95819
R302 VDD2 VDD2.n4 1.66645
R303 B.n640 B.n639 585
R304 B.n641 B.n80 585
R305 B.n643 B.n642 585
R306 B.n644 B.n79 585
R307 B.n646 B.n645 585
R308 B.n647 B.n78 585
R309 B.n649 B.n648 585
R310 B.n650 B.n77 585
R311 B.n652 B.n651 585
R312 B.n653 B.n76 585
R313 B.n655 B.n654 585
R314 B.n656 B.n75 585
R315 B.n658 B.n657 585
R316 B.n659 B.n74 585
R317 B.n661 B.n660 585
R318 B.n662 B.n73 585
R319 B.n664 B.n663 585
R320 B.n665 B.n72 585
R321 B.n667 B.n666 585
R322 B.n668 B.n71 585
R323 B.n670 B.n669 585
R324 B.n671 B.n70 585
R325 B.n673 B.n672 585
R326 B.n674 B.n69 585
R327 B.n676 B.n675 585
R328 B.n677 B.n68 585
R329 B.n679 B.n678 585
R330 B.n680 B.n67 585
R331 B.n682 B.n681 585
R332 B.n683 B.n66 585
R333 B.n685 B.n684 585
R334 B.n686 B.n65 585
R335 B.n688 B.n687 585
R336 B.n689 B.n64 585
R337 B.n691 B.n690 585
R338 B.n692 B.n63 585
R339 B.n694 B.n693 585
R340 B.n695 B.n62 585
R341 B.n697 B.n696 585
R342 B.n699 B.n59 585
R343 B.n701 B.n700 585
R344 B.n702 B.n58 585
R345 B.n704 B.n703 585
R346 B.n705 B.n57 585
R347 B.n707 B.n706 585
R348 B.n708 B.n56 585
R349 B.n710 B.n709 585
R350 B.n711 B.n53 585
R351 B.n714 B.n713 585
R352 B.n715 B.n52 585
R353 B.n717 B.n716 585
R354 B.n718 B.n51 585
R355 B.n720 B.n719 585
R356 B.n721 B.n50 585
R357 B.n723 B.n722 585
R358 B.n724 B.n49 585
R359 B.n726 B.n725 585
R360 B.n727 B.n48 585
R361 B.n729 B.n728 585
R362 B.n730 B.n47 585
R363 B.n732 B.n731 585
R364 B.n733 B.n46 585
R365 B.n735 B.n734 585
R366 B.n736 B.n45 585
R367 B.n738 B.n737 585
R368 B.n739 B.n44 585
R369 B.n741 B.n740 585
R370 B.n742 B.n43 585
R371 B.n744 B.n743 585
R372 B.n745 B.n42 585
R373 B.n747 B.n746 585
R374 B.n748 B.n41 585
R375 B.n750 B.n749 585
R376 B.n751 B.n40 585
R377 B.n753 B.n752 585
R378 B.n754 B.n39 585
R379 B.n756 B.n755 585
R380 B.n757 B.n38 585
R381 B.n759 B.n758 585
R382 B.n760 B.n37 585
R383 B.n762 B.n761 585
R384 B.n763 B.n36 585
R385 B.n765 B.n764 585
R386 B.n766 B.n35 585
R387 B.n768 B.n767 585
R388 B.n769 B.n34 585
R389 B.n771 B.n770 585
R390 B.n638 B.n81 585
R391 B.n637 B.n636 585
R392 B.n635 B.n82 585
R393 B.n634 B.n633 585
R394 B.n632 B.n83 585
R395 B.n631 B.n630 585
R396 B.n629 B.n84 585
R397 B.n628 B.n627 585
R398 B.n626 B.n85 585
R399 B.n625 B.n624 585
R400 B.n623 B.n86 585
R401 B.n622 B.n621 585
R402 B.n620 B.n87 585
R403 B.n619 B.n618 585
R404 B.n617 B.n88 585
R405 B.n616 B.n615 585
R406 B.n614 B.n89 585
R407 B.n613 B.n612 585
R408 B.n611 B.n90 585
R409 B.n610 B.n609 585
R410 B.n608 B.n91 585
R411 B.n607 B.n606 585
R412 B.n605 B.n92 585
R413 B.n604 B.n603 585
R414 B.n602 B.n93 585
R415 B.n601 B.n600 585
R416 B.n599 B.n94 585
R417 B.n598 B.n597 585
R418 B.n596 B.n95 585
R419 B.n595 B.n594 585
R420 B.n593 B.n96 585
R421 B.n592 B.n591 585
R422 B.n590 B.n97 585
R423 B.n589 B.n588 585
R424 B.n587 B.n98 585
R425 B.n586 B.n585 585
R426 B.n584 B.n99 585
R427 B.n583 B.n582 585
R428 B.n581 B.n100 585
R429 B.n580 B.n579 585
R430 B.n578 B.n101 585
R431 B.n577 B.n576 585
R432 B.n575 B.n102 585
R433 B.n574 B.n573 585
R434 B.n572 B.n103 585
R435 B.n571 B.n570 585
R436 B.n569 B.n104 585
R437 B.n568 B.n567 585
R438 B.n566 B.n105 585
R439 B.n565 B.n564 585
R440 B.n563 B.n106 585
R441 B.n562 B.n561 585
R442 B.n560 B.n107 585
R443 B.n559 B.n558 585
R444 B.n557 B.n108 585
R445 B.n556 B.n555 585
R446 B.n554 B.n109 585
R447 B.n553 B.n552 585
R448 B.n551 B.n110 585
R449 B.n550 B.n549 585
R450 B.n548 B.n111 585
R451 B.n547 B.n546 585
R452 B.n545 B.n112 585
R453 B.n544 B.n543 585
R454 B.n542 B.n113 585
R455 B.n541 B.n540 585
R456 B.n539 B.n114 585
R457 B.n538 B.n537 585
R458 B.n536 B.n115 585
R459 B.n535 B.n534 585
R460 B.n533 B.n116 585
R461 B.n532 B.n531 585
R462 B.n530 B.n117 585
R463 B.n529 B.n528 585
R464 B.n527 B.n118 585
R465 B.n526 B.n525 585
R466 B.n524 B.n119 585
R467 B.n523 B.n522 585
R468 B.n521 B.n120 585
R469 B.n520 B.n519 585
R470 B.n518 B.n121 585
R471 B.n517 B.n516 585
R472 B.n515 B.n122 585
R473 B.n514 B.n513 585
R474 B.n512 B.n123 585
R475 B.n511 B.n510 585
R476 B.n509 B.n124 585
R477 B.n508 B.n507 585
R478 B.n506 B.n125 585
R479 B.n505 B.n504 585
R480 B.n503 B.n126 585
R481 B.n502 B.n501 585
R482 B.n500 B.n127 585
R483 B.n499 B.n498 585
R484 B.n497 B.n128 585
R485 B.n496 B.n495 585
R486 B.n494 B.n129 585
R487 B.n493 B.n492 585
R488 B.n491 B.n130 585
R489 B.n490 B.n489 585
R490 B.n488 B.n131 585
R491 B.n487 B.n486 585
R492 B.n485 B.n132 585
R493 B.n484 B.n483 585
R494 B.n482 B.n133 585
R495 B.n481 B.n480 585
R496 B.n479 B.n134 585
R497 B.n478 B.n477 585
R498 B.n476 B.n135 585
R499 B.n475 B.n474 585
R500 B.n473 B.n136 585
R501 B.n472 B.n471 585
R502 B.n470 B.n137 585
R503 B.n469 B.n468 585
R504 B.n467 B.n138 585
R505 B.n466 B.n465 585
R506 B.n464 B.n139 585
R507 B.n463 B.n462 585
R508 B.n461 B.n140 585
R509 B.n460 B.n459 585
R510 B.n458 B.n141 585
R511 B.n457 B.n456 585
R512 B.n455 B.n142 585
R513 B.n454 B.n453 585
R514 B.n452 B.n143 585
R515 B.n451 B.n450 585
R516 B.n449 B.n144 585
R517 B.n317 B.n192 585
R518 B.n319 B.n318 585
R519 B.n320 B.n191 585
R520 B.n322 B.n321 585
R521 B.n323 B.n190 585
R522 B.n325 B.n324 585
R523 B.n326 B.n189 585
R524 B.n328 B.n327 585
R525 B.n329 B.n188 585
R526 B.n331 B.n330 585
R527 B.n332 B.n187 585
R528 B.n334 B.n333 585
R529 B.n335 B.n186 585
R530 B.n337 B.n336 585
R531 B.n338 B.n185 585
R532 B.n340 B.n339 585
R533 B.n341 B.n184 585
R534 B.n343 B.n342 585
R535 B.n344 B.n183 585
R536 B.n346 B.n345 585
R537 B.n347 B.n182 585
R538 B.n349 B.n348 585
R539 B.n350 B.n181 585
R540 B.n352 B.n351 585
R541 B.n353 B.n180 585
R542 B.n355 B.n354 585
R543 B.n356 B.n179 585
R544 B.n358 B.n357 585
R545 B.n359 B.n178 585
R546 B.n361 B.n360 585
R547 B.n362 B.n177 585
R548 B.n364 B.n363 585
R549 B.n365 B.n176 585
R550 B.n367 B.n366 585
R551 B.n368 B.n175 585
R552 B.n370 B.n369 585
R553 B.n371 B.n174 585
R554 B.n373 B.n372 585
R555 B.n374 B.n171 585
R556 B.n377 B.n376 585
R557 B.n378 B.n170 585
R558 B.n380 B.n379 585
R559 B.n381 B.n169 585
R560 B.n383 B.n382 585
R561 B.n384 B.n168 585
R562 B.n386 B.n385 585
R563 B.n387 B.n167 585
R564 B.n389 B.n388 585
R565 B.n391 B.n390 585
R566 B.n392 B.n163 585
R567 B.n394 B.n393 585
R568 B.n395 B.n162 585
R569 B.n397 B.n396 585
R570 B.n398 B.n161 585
R571 B.n400 B.n399 585
R572 B.n401 B.n160 585
R573 B.n403 B.n402 585
R574 B.n404 B.n159 585
R575 B.n406 B.n405 585
R576 B.n407 B.n158 585
R577 B.n409 B.n408 585
R578 B.n410 B.n157 585
R579 B.n412 B.n411 585
R580 B.n413 B.n156 585
R581 B.n415 B.n414 585
R582 B.n416 B.n155 585
R583 B.n418 B.n417 585
R584 B.n419 B.n154 585
R585 B.n421 B.n420 585
R586 B.n422 B.n153 585
R587 B.n424 B.n423 585
R588 B.n425 B.n152 585
R589 B.n427 B.n426 585
R590 B.n428 B.n151 585
R591 B.n430 B.n429 585
R592 B.n431 B.n150 585
R593 B.n433 B.n432 585
R594 B.n434 B.n149 585
R595 B.n436 B.n435 585
R596 B.n437 B.n148 585
R597 B.n439 B.n438 585
R598 B.n440 B.n147 585
R599 B.n442 B.n441 585
R600 B.n443 B.n146 585
R601 B.n445 B.n444 585
R602 B.n446 B.n145 585
R603 B.n448 B.n447 585
R604 B.n316 B.n315 585
R605 B.n314 B.n193 585
R606 B.n313 B.n312 585
R607 B.n311 B.n194 585
R608 B.n310 B.n309 585
R609 B.n308 B.n195 585
R610 B.n307 B.n306 585
R611 B.n305 B.n196 585
R612 B.n304 B.n303 585
R613 B.n302 B.n197 585
R614 B.n301 B.n300 585
R615 B.n299 B.n198 585
R616 B.n298 B.n297 585
R617 B.n296 B.n199 585
R618 B.n295 B.n294 585
R619 B.n293 B.n200 585
R620 B.n292 B.n291 585
R621 B.n290 B.n201 585
R622 B.n289 B.n288 585
R623 B.n287 B.n202 585
R624 B.n286 B.n285 585
R625 B.n284 B.n203 585
R626 B.n283 B.n282 585
R627 B.n281 B.n204 585
R628 B.n280 B.n279 585
R629 B.n278 B.n205 585
R630 B.n277 B.n276 585
R631 B.n275 B.n206 585
R632 B.n274 B.n273 585
R633 B.n272 B.n207 585
R634 B.n271 B.n270 585
R635 B.n269 B.n208 585
R636 B.n268 B.n267 585
R637 B.n266 B.n209 585
R638 B.n265 B.n264 585
R639 B.n263 B.n210 585
R640 B.n262 B.n261 585
R641 B.n260 B.n211 585
R642 B.n259 B.n258 585
R643 B.n257 B.n212 585
R644 B.n256 B.n255 585
R645 B.n254 B.n213 585
R646 B.n253 B.n252 585
R647 B.n251 B.n214 585
R648 B.n250 B.n249 585
R649 B.n248 B.n215 585
R650 B.n247 B.n246 585
R651 B.n245 B.n216 585
R652 B.n244 B.n243 585
R653 B.n242 B.n217 585
R654 B.n241 B.n240 585
R655 B.n239 B.n218 585
R656 B.n238 B.n237 585
R657 B.n236 B.n219 585
R658 B.n235 B.n234 585
R659 B.n233 B.n220 585
R660 B.n232 B.n231 585
R661 B.n230 B.n221 585
R662 B.n229 B.n228 585
R663 B.n227 B.n222 585
R664 B.n226 B.n225 585
R665 B.n224 B.n223 585
R666 B.n2 B.n0 585
R667 B.n865 B.n1 585
R668 B.n864 B.n863 585
R669 B.n862 B.n3 585
R670 B.n861 B.n860 585
R671 B.n859 B.n4 585
R672 B.n858 B.n857 585
R673 B.n856 B.n5 585
R674 B.n855 B.n854 585
R675 B.n853 B.n6 585
R676 B.n852 B.n851 585
R677 B.n850 B.n7 585
R678 B.n849 B.n848 585
R679 B.n847 B.n8 585
R680 B.n846 B.n845 585
R681 B.n844 B.n9 585
R682 B.n843 B.n842 585
R683 B.n841 B.n10 585
R684 B.n840 B.n839 585
R685 B.n838 B.n11 585
R686 B.n837 B.n836 585
R687 B.n835 B.n12 585
R688 B.n834 B.n833 585
R689 B.n832 B.n13 585
R690 B.n831 B.n830 585
R691 B.n829 B.n14 585
R692 B.n828 B.n827 585
R693 B.n826 B.n15 585
R694 B.n825 B.n824 585
R695 B.n823 B.n16 585
R696 B.n822 B.n821 585
R697 B.n820 B.n17 585
R698 B.n819 B.n818 585
R699 B.n817 B.n18 585
R700 B.n816 B.n815 585
R701 B.n814 B.n19 585
R702 B.n813 B.n812 585
R703 B.n811 B.n20 585
R704 B.n810 B.n809 585
R705 B.n808 B.n21 585
R706 B.n807 B.n806 585
R707 B.n805 B.n22 585
R708 B.n804 B.n803 585
R709 B.n802 B.n23 585
R710 B.n801 B.n800 585
R711 B.n799 B.n24 585
R712 B.n798 B.n797 585
R713 B.n796 B.n25 585
R714 B.n795 B.n794 585
R715 B.n793 B.n26 585
R716 B.n792 B.n791 585
R717 B.n790 B.n27 585
R718 B.n789 B.n788 585
R719 B.n787 B.n28 585
R720 B.n786 B.n785 585
R721 B.n784 B.n29 585
R722 B.n783 B.n782 585
R723 B.n781 B.n30 585
R724 B.n780 B.n779 585
R725 B.n778 B.n31 585
R726 B.n777 B.n776 585
R727 B.n775 B.n32 585
R728 B.n774 B.n773 585
R729 B.n772 B.n33 585
R730 B.n867 B.n866 585
R731 B.n317 B.n316 482.89
R732 B.n770 B.n33 482.89
R733 B.n449 B.n448 482.89
R734 B.n640 B.n81 482.89
R735 B.n164 B.t9 286.901
R736 B.n172 B.t3 286.901
R737 B.n54 B.t6 286.901
R738 B.n60 B.t0 286.901
R739 B.n164 B.t11 181.834
R740 B.n60 B.t1 181.834
R741 B.n172 B.t5 181.821
R742 B.n54 B.t7 181.821
R743 B.n316 B.n193 163.367
R744 B.n312 B.n193 163.367
R745 B.n312 B.n311 163.367
R746 B.n311 B.n310 163.367
R747 B.n310 B.n195 163.367
R748 B.n306 B.n195 163.367
R749 B.n306 B.n305 163.367
R750 B.n305 B.n304 163.367
R751 B.n304 B.n197 163.367
R752 B.n300 B.n197 163.367
R753 B.n300 B.n299 163.367
R754 B.n299 B.n298 163.367
R755 B.n298 B.n199 163.367
R756 B.n294 B.n199 163.367
R757 B.n294 B.n293 163.367
R758 B.n293 B.n292 163.367
R759 B.n292 B.n201 163.367
R760 B.n288 B.n201 163.367
R761 B.n288 B.n287 163.367
R762 B.n287 B.n286 163.367
R763 B.n286 B.n203 163.367
R764 B.n282 B.n203 163.367
R765 B.n282 B.n281 163.367
R766 B.n281 B.n280 163.367
R767 B.n280 B.n205 163.367
R768 B.n276 B.n205 163.367
R769 B.n276 B.n275 163.367
R770 B.n275 B.n274 163.367
R771 B.n274 B.n207 163.367
R772 B.n270 B.n207 163.367
R773 B.n270 B.n269 163.367
R774 B.n269 B.n268 163.367
R775 B.n268 B.n209 163.367
R776 B.n264 B.n209 163.367
R777 B.n264 B.n263 163.367
R778 B.n263 B.n262 163.367
R779 B.n262 B.n211 163.367
R780 B.n258 B.n211 163.367
R781 B.n258 B.n257 163.367
R782 B.n257 B.n256 163.367
R783 B.n256 B.n213 163.367
R784 B.n252 B.n213 163.367
R785 B.n252 B.n251 163.367
R786 B.n251 B.n250 163.367
R787 B.n250 B.n215 163.367
R788 B.n246 B.n215 163.367
R789 B.n246 B.n245 163.367
R790 B.n245 B.n244 163.367
R791 B.n244 B.n217 163.367
R792 B.n240 B.n217 163.367
R793 B.n240 B.n239 163.367
R794 B.n239 B.n238 163.367
R795 B.n238 B.n219 163.367
R796 B.n234 B.n219 163.367
R797 B.n234 B.n233 163.367
R798 B.n233 B.n232 163.367
R799 B.n232 B.n221 163.367
R800 B.n228 B.n221 163.367
R801 B.n228 B.n227 163.367
R802 B.n227 B.n226 163.367
R803 B.n226 B.n223 163.367
R804 B.n223 B.n2 163.367
R805 B.n866 B.n2 163.367
R806 B.n866 B.n865 163.367
R807 B.n865 B.n864 163.367
R808 B.n864 B.n3 163.367
R809 B.n860 B.n3 163.367
R810 B.n860 B.n859 163.367
R811 B.n859 B.n858 163.367
R812 B.n858 B.n5 163.367
R813 B.n854 B.n5 163.367
R814 B.n854 B.n853 163.367
R815 B.n853 B.n852 163.367
R816 B.n852 B.n7 163.367
R817 B.n848 B.n7 163.367
R818 B.n848 B.n847 163.367
R819 B.n847 B.n846 163.367
R820 B.n846 B.n9 163.367
R821 B.n842 B.n9 163.367
R822 B.n842 B.n841 163.367
R823 B.n841 B.n840 163.367
R824 B.n840 B.n11 163.367
R825 B.n836 B.n11 163.367
R826 B.n836 B.n835 163.367
R827 B.n835 B.n834 163.367
R828 B.n834 B.n13 163.367
R829 B.n830 B.n13 163.367
R830 B.n830 B.n829 163.367
R831 B.n829 B.n828 163.367
R832 B.n828 B.n15 163.367
R833 B.n824 B.n15 163.367
R834 B.n824 B.n823 163.367
R835 B.n823 B.n822 163.367
R836 B.n822 B.n17 163.367
R837 B.n818 B.n17 163.367
R838 B.n818 B.n817 163.367
R839 B.n817 B.n816 163.367
R840 B.n816 B.n19 163.367
R841 B.n812 B.n19 163.367
R842 B.n812 B.n811 163.367
R843 B.n811 B.n810 163.367
R844 B.n810 B.n21 163.367
R845 B.n806 B.n21 163.367
R846 B.n806 B.n805 163.367
R847 B.n805 B.n804 163.367
R848 B.n804 B.n23 163.367
R849 B.n800 B.n23 163.367
R850 B.n800 B.n799 163.367
R851 B.n799 B.n798 163.367
R852 B.n798 B.n25 163.367
R853 B.n794 B.n25 163.367
R854 B.n794 B.n793 163.367
R855 B.n793 B.n792 163.367
R856 B.n792 B.n27 163.367
R857 B.n788 B.n27 163.367
R858 B.n788 B.n787 163.367
R859 B.n787 B.n786 163.367
R860 B.n786 B.n29 163.367
R861 B.n782 B.n29 163.367
R862 B.n782 B.n781 163.367
R863 B.n781 B.n780 163.367
R864 B.n780 B.n31 163.367
R865 B.n776 B.n31 163.367
R866 B.n776 B.n775 163.367
R867 B.n775 B.n774 163.367
R868 B.n774 B.n33 163.367
R869 B.n318 B.n317 163.367
R870 B.n318 B.n191 163.367
R871 B.n322 B.n191 163.367
R872 B.n323 B.n322 163.367
R873 B.n324 B.n323 163.367
R874 B.n324 B.n189 163.367
R875 B.n328 B.n189 163.367
R876 B.n329 B.n328 163.367
R877 B.n330 B.n329 163.367
R878 B.n330 B.n187 163.367
R879 B.n334 B.n187 163.367
R880 B.n335 B.n334 163.367
R881 B.n336 B.n335 163.367
R882 B.n336 B.n185 163.367
R883 B.n340 B.n185 163.367
R884 B.n341 B.n340 163.367
R885 B.n342 B.n341 163.367
R886 B.n342 B.n183 163.367
R887 B.n346 B.n183 163.367
R888 B.n347 B.n346 163.367
R889 B.n348 B.n347 163.367
R890 B.n348 B.n181 163.367
R891 B.n352 B.n181 163.367
R892 B.n353 B.n352 163.367
R893 B.n354 B.n353 163.367
R894 B.n354 B.n179 163.367
R895 B.n358 B.n179 163.367
R896 B.n359 B.n358 163.367
R897 B.n360 B.n359 163.367
R898 B.n360 B.n177 163.367
R899 B.n364 B.n177 163.367
R900 B.n365 B.n364 163.367
R901 B.n366 B.n365 163.367
R902 B.n366 B.n175 163.367
R903 B.n370 B.n175 163.367
R904 B.n371 B.n370 163.367
R905 B.n372 B.n371 163.367
R906 B.n372 B.n171 163.367
R907 B.n377 B.n171 163.367
R908 B.n378 B.n377 163.367
R909 B.n379 B.n378 163.367
R910 B.n379 B.n169 163.367
R911 B.n383 B.n169 163.367
R912 B.n384 B.n383 163.367
R913 B.n385 B.n384 163.367
R914 B.n385 B.n167 163.367
R915 B.n389 B.n167 163.367
R916 B.n390 B.n389 163.367
R917 B.n390 B.n163 163.367
R918 B.n394 B.n163 163.367
R919 B.n395 B.n394 163.367
R920 B.n396 B.n395 163.367
R921 B.n396 B.n161 163.367
R922 B.n400 B.n161 163.367
R923 B.n401 B.n400 163.367
R924 B.n402 B.n401 163.367
R925 B.n402 B.n159 163.367
R926 B.n406 B.n159 163.367
R927 B.n407 B.n406 163.367
R928 B.n408 B.n407 163.367
R929 B.n408 B.n157 163.367
R930 B.n412 B.n157 163.367
R931 B.n413 B.n412 163.367
R932 B.n414 B.n413 163.367
R933 B.n414 B.n155 163.367
R934 B.n418 B.n155 163.367
R935 B.n419 B.n418 163.367
R936 B.n420 B.n419 163.367
R937 B.n420 B.n153 163.367
R938 B.n424 B.n153 163.367
R939 B.n425 B.n424 163.367
R940 B.n426 B.n425 163.367
R941 B.n426 B.n151 163.367
R942 B.n430 B.n151 163.367
R943 B.n431 B.n430 163.367
R944 B.n432 B.n431 163.367
R945 B.n432 B.n149 163.367
R946 B.n436 B.n149 163.367
R947 B.n437 B.n436 163.367
R948 B.n438 B.n437 163.367
R949 B.n438 B.n147 163.367
R950 B.n442 B.n147 163.367
R951 B.n443 B.n442 163.367
R952 B.n444 B.n443 163.367
R953 B.n444 B.n145 163.367
R954 B.n448 B.n145 163.367
R955 B.n450 B.n449 163.367
R956 B.n450 B.n143 163.367
R957 B.n454 B.n143 163.367
R958 B.n455 B.n454 163.367
R959 B.n456 B.n455 163.367
R960 B.n456 B.n141 163.367
R961 B.n460 B.n141 163.367
R962 B.n461 B.n460 163.367
R963 B.n462 B.n461 163.367
R964 B.n462 B.n139 163.367
R965 B.n466 B.n139 163.367
R966 B.n467 B.n466 163.367
R967 B.n468 B.n467 163.367
R968 B.n468 B.n137 163.367
R969 B.n472 B.n137 163.367
R970 B.n473 B.n472 163.367
R971 B.n474 B.n473 163.367
R972 B.n474 B.n135 163.367
R973 B.n478 B.n135 163.367
R974 B.n479 B.n478 163.367
R975 B.n480 B.n479 163.367
R976 B.n480 B.n133 163.367
R977 B.n484 B.n133 163.367
R978 B.n485 B.n484 163.367
R979 B.n486 B.n485 163.367
R980 B.n486 B.n131 163.367
R981 B.n490 B.n131 163.367
R982 B.n491 B.n490 163.367
R983 B.n492 B.n491 163.367
R984 B.n492 B.n129 163.367
R985 B.n496 B.n129 163.367
R986 B.n497 B.n496 163.367
R987 B.n498 B.n497 163.367
R988 B.n498 B.n127 163.367
R989 B.n502 B.n127 163.367
R990 B.n503 B.n502 163.367
R991 B.n504 B.n503 163.367
R992 B.n504 B.n125 163.367
R993 B.n508 B.n125 163.367
R994 B.n509 B.n508 163.367
R995 B.n510 B.n509 163.367
R996 B.n510 B.n123 163.367
R997 B.n514 B.n123 163.367
R998 B.n515 B.n514 163.367
R999 B.n516 B.n515 163.367
R1000 B.n516 B.n121 163.367
R1001 B.n520 B.n121 163.367
R1002 B.n521 B.n520 163.367
R1003 B.n522 B.n521 163.367
R1004 B.n522 B.n119 163.367
R1005 B.n526 B.n119 163.367
R1006 B.n527 B.n526 163.367
R1007 B.n528 B.n527 163.367
R1008 B.n528 B.n117 163.367
R1009 B.n532 B.n117 163.367
R1010 B.n533 B.n532 163.367
R1011 B.n534 B.n533 163.367
R1012 B.n534 B.n115 163.367
R1013 B.n538 B.n115 163.367
R1014 B.n539 B.n538 163.367
R1015 B.n540 B.n539 163.367
R1016 B.n540 B.n113 163.367
R1017 B.n544 B.n113 163.367
R1018 B.n545 B.n544 163.367
R1019 B.n546 B.n545 163.367
R1020 B.n546 B.n111 163.367
R1021 B.n550 B.n111 163.367
R1022 B.n551 B.n550 163.367
R1023 B.n552 B.n551 163.367
R1024 B.n552 B.n109 163.367
R1025 B.n556 B.n109 163.367
R1026 B.n557 B.n556 163.367
R1027 B.n558 B.n557 163.367
R1028 B.n558 B.n107 163.367
R1029 B.n562 B.n107 163.367
R1030 B.n563 B.n562 163.367
R1031 B.n564 B.n563 163.367
R1032 B.n564 B.n105 163.367
R1033 B.n568 B.n105 163.367
R1034 B.n569 B.n568 163.367
R1035 B.n570 B.n569 163.367
R1036 B.n570 B.n103 163.367
R1037 B.n574 B.n103 163.367
R1038 B.n575 B.n574 163.367
R1039 B.n576 B.n575 163.367
R1040 B.n576 B.n101 163.367
R1041 B.n580 B.n101 163.367
R1042 B.n581 B.n580 163.367
R1043 B.n582 B.n581 163.367
R1044 B.n582 B.n99 163.367
R1045 B.n586 B.n99 163.367
R1046 B.n587 B.n586 163.367
R1047 B.n588 B.n587 163.367
R1048 B.n588 B.n97 163.367
R1049 B.n592 B.n97 163.367
R1050 B.n593 B.n592 163.367
R1051 B.n594 B.n593 163.367
R1052 B.n594 B.n95 163.367
R1053 B.n598 B.n95 163.367
R1054 B.n599 B.n598 163.367
R1055 B.n600 B.n599 163.367
R1056 B.n600 B.n93 163.367
R1057 B.n604 B.n93 163.367
R1058 B.n605 B.n604 163.367
R1059 B.n606 B.n605 163.367
R1060 B.n606 B.n91 163.367
R1061 B.n610 B.n91 163.367
R1062 B.n611 B.n610 163.367
R1063 B.n612 B.n611 163.367
R1064 B.n612 B.n89 163.367
R1065 B.n616 B.n89 163.367
R1066 B.n617 B.n616 163.367
R1067 B.n618 B.n617 163.367
R1068 B.n618 B.n87 163.367
R1069 B.n622 B.n87 163.367
R1070 B.n623 B.n622 163.367
R1071 B.n624 B.n623 163.367
R1072 B.n624 B.n85 163.367
R1073 B.n628 B.n85 163.367
R1074 B.n629 B.n628 163.367
R1075 B.n630 B.n629 163.367
R1076 B.n630 B.n83 163.367
R1077 B.n634 B.n83 163.367
R1078 B.n635 B.n634 163.367
R1079 B.n636 B.n635 163.367
R1080 B.n636 B.n81 163.367
R1081 B.n770 B.n769 163.367
R1082 B.n769 B.n768 163.367
R1083 B.n768 B.n35 163.367
R1084 B.n764 B.n35 163.367
R1085 B.n764 B.n763 163.367
R1086 B.n763 B.n762 163.367
R1087 B.n762 B.n37 163.367
R1088 B.n758 B.n37 163.367
R1089 B.n758 B.n757 163.367
R1090 B.n757 B.n756 163.367
R1091 B.n756 B.n39 163.367
R1092 B.n752 B.n39 163.367
R1093 B.n752 B.n751 163.367
R1094 B.n751 B.n750 163.367
R1095 B.n750 B.n41 163.367
R1096 B.n746 B.n41 163.367
R1097 B.n746 B.n745 163.367
R1098 B.n745 B.n744 163.367
R1099 B.n744 B.n43 163.367
R1100 B.n740 B.n43 163.367
R1101 B.n740 B.n739 163.367
R1102 B.n739 B.n738 163.367
R1103 B.n738 B.n45 163.367
R1104 B.n734 B.n45 163.367
R1105 B.n734 B.n733 163.367
R1106 B.n733 B.n732 163.367
R1107 B.n732 B.n47 163.367
R1108 B.n728 B.n47 163.367
R1109 B.n728 B.n727 163.367
R1110 B.n727 B.n726 163.367
R1111 B.n726 B.n49 163.367
R1112 B.n722 B.n49 163.367
R1113 B.n722 B.n721 163.367
R1114 B.n721 B.n720 163.367
R1115 B.n720 B.n51 163.367
R1116 B.n716 B.n51 163.367
R1117 B.n716 B.n715 163.367
R1118 B.n715 B.n714 163.367
R1119 B.n714 B.n53 163.367
R1120 B.n709 B.n53 163.367
R1121 B.n709 B.n708 163.367
R1122 B.n708 B.n707 163.367
R1123 B.n707 B.n57 163.367
R1124 B.n703 B.n57 163.367
R1125 B.n703 B.n702 163.367
R1126 B.n702 B.n701 163.367
R1127 B.n701 B.n59 163.367
R1128 B.n696 B.n59 163.367
R1129 B.n696 B.n695 163.367
R1130 B.n695 B.n694 163.367
R1131 B.n694 B.n63 163.367
R1132 B.n690 B.n63 163.367
R1133 B.n690 B.n689 163.367
R1134 B.n689 B.n688 163.367
R1135 B.n688 B.n65 163.367
R1136 B.n684 B.n65 163.367
R1137 B.n684 B.n683 163.367
R1138 B.n683 B.n682 163.367
R1139 B.n682 B.n67 163.367
R1140 B.n678 B.n67 163.367
R1141 B.n678 B.n677 163.367
R1142 B.n677 B.n676 163.367
R1143 B.n676 B.n69 163.367
R1144 B.n672 B.n69 163.367
R1145 B.n672 B.n671 163.367
R1146 B.n671 B.n670 163.367
R1147 B.n670 B.n71 163.367
R1148 B.n666 B.n71 163.367
R1149 B.n666 B.n665 163.367
R1150 B.n665 B.n664 163.367
R1151 B.n664 B.n73 163.367
R1152 B.n660 B.n73 163.367
R1153 B.n660 B.n659 163.367
R1154 B.n659 B.n658 163.367
R1155 B.n658 B.n75 163.367
R1156 B.n654 B.n75 163.367
R1157 B.n654 B.n653 163.367
R1158 B.n653 B.n652 163.367
R1159 B.n652 B.n77 163.367
R1160 B.n648 B.n77 163.367
R1161 B.n648 B.n647 163.367
R1162 B.n647 B.n646 163.367
R1163 B.n646 B.n79 163.367
R1164 B.n642 B.n79 163.367
R1165 B.n642 B.n641 163.367
R1166 B.n641 B.n640 163.367
R1167 B.n165 B.t10 109.496
R1168 B.n61 B.t2 109.496
R1169 B.n173 B.t4 109.483
R1170 B.n55 B.t8 109.483
R1171 B.n165 B.n164 72.3399
R1172 B.n173 B.n172 72.3399
R1173 B.n55 B.n54 72.3399
R1174 B.n61 B.n60 72.3399
R1175 B.n166 B.n165 59.5399
R1176 B.n375 B.n173 59.5399
R1177 B.n712 B.n55 59.5399
R1178 B.n698 B.n61 59.5399
R1179 B.n772 B.n771 31.3761
R1180 B.n639 B.n638 31.3761
R1181 B.n447 B.n144 31.3761
R1182 B.n315 B.n192 31.3761
R1183 B B.n867 18.0485
R1184 B.n771 B.n34 10.6151
R1185 B.n767 B.n34 10.6151
R1186 B.n767 B.n766 10.6151
R1187 B.n766 B.n765 10.6151
R1188 B.n765 B.n36 10.6151
R1189 B.n761 B.n36 10.6151
R1190 B.n761 B.n760 10.6151
R1191 B.n760 B.n759 10.6151
R1192 B.n759 B.n38 10.6151
R1193 B.n755 B.n38 10.6151
R1194 B.n755 B.n754 10.6151
R1195 B.n754 B.n753 10.6151
R1196 B.n753 B.n40 10.6151
R1197 B.n749 B.n40 10.6151
R1198 B.n749 B.n748 10.6151
R1199 B.n748 B.n747 10.6151
R1200 B.n747 B.n42 10.6151
R1201 B.n743 B.n42 10.6151
R1202 B.n743 B.n742 10.6151
R1203 B.n742 B.n741 10.6151
R1204 B.n741 B.n44 10.6151
R1205 B.n737 B.n44 10.6151
R1206 B.n737 B.n736 10.6151
R1207 B.n736 B.n735 10.6151
R1208 B.n735 B.n46 10.6151
R1209 B.n731 B.n46 10.6151
R1210 B.n731 B.n730 10.6151
R1211 B.n730 B.n729 10.6151
R1212 B.n729 B.n48 10.6151
R1213 B.n725 B.n48 10.6151
R1214 B.n725 B.n724 10.6151
R1215 B.n724 B.n723 10.6151
R1216 B.n723 B.n50 10.6151
R1217 B.n719 B.n50 10.6151
R1218 B.n719 B.n718 10.6151
R1219 B.n718 B.n717 10.6151
R1220 B.n717 B.n52 10.6151
R1221 B.n713 B.n52 10.6151
R1222 B.n711 B.n710 10.6151
R1223 B.n710 B.n56 10.6151
R1224 B.n706 B.n56 10.6151
R1225 B.n706 B.n705 10.6151
R1226 B.n705 B.n704 10.6151
R1227 B.n704 B.n58 10.6151
R1228 B.n700 B.n58 10.6151
R1229 B.n700 B.n699 10.6151
R1230 B.n697 B.n62 10.6151
R1231 B.n693 B.n62 10.6151
R1232 B.n693 B.n692 10.6151
R1233 B.n692 B.n691 10.6151
R1234 B.n691 B.n64 10.6151
R1235 B.n687 B.n64 10.6151
R1236 B.n687 B.n686 10.6151
R1237 B.n686 B.n685 10.6151
R1238 B.n685 B.n66 10.6151
R1239 B.n681 B.n66 10.6151
R1240 B.n681 B.n680 10.6151
R1241 B.n680 B.n679 10.6151
R1242 B.n679 B.n68 10.6151
R1243 B.n675 B.n68 10.6151
R1244 B.n675 B.n674 10.6151
R1245 B.n674 B.n673 10.6151
R1246 B.n673 B.n70 10.6151
R1247 B.n669 B.n70 10.6151
R1248 B.n669 B.n668 10.6151
R1249 B.n668 B.n667 10.6151
R1250 B.n667 B.n72 10.6151
R1251 B.n663 B.n72 10.6151
R1252 B.n663 B.n662 10.6151
R1253 B.n662 B.n661 10.6151
R1254 B.n661 B.n74 10.6151
R1255 B.n657 B.n74 10.6151
R1256 B.n657 B.n656 10.6151
R1257 B.n656 B.n655 10.6151
R1258 B.n655 B.n76 10.6151
R1259 B.n651 B.n76 10.6151
R1260 B.n651 B.n650 10.6151
R1261 B.n650 B.n649 10.6151
R1262 B.n649 B.n78 10.6151
R1263 B.n645 B.n78 10.6151
R1264 B.n645 B.n644 10.6151
R1265 B.n644 B.n643 10.6151
R1266 B.n643 B.n80 10.6151
R1267 B.n639 B.n80 10.6151
R1268 B.n451 B.n144 10.6151
R1269 B.n452 B.n451 10.6151
R1270 B.n453 B.n452 10.6151
R1271 B.n453 B.n142 10.6151
R1272 B.n457 B.n142 10.6151
R1273 B.n458 B.n457 10.6151
R1274 B.n459 B.n458 10.6151
R1275 B.n459 B.n140 10.6151
R1276 B.n463 B.n140 10.6151
R1277 B.n464 B.n463 10.6151
R1278 B.n465 B.n464 10.6151
R1279 B.n465 B.n138 10.6151
R1280 B.n469 B.n138 10.6151
R1281 B.n470 B.n469 10.6151
R1282 B.n471 B.n470 10.6151
R1283 B.n471 B.n136 10.6151
R1284 B.n475 B.n136 10.6151
R1285 B.n476 B.n475 10.6151
R1286 B.n477 B.n476 10.6151
R1287 B.n477 B.n134 10.6151
R1288 B.n481 B.n134 10.6151
R1289 B.n482 B.n481 10.6151
R1290 B.n483 B.n482 10.6151
R1291 B.n483 B.n132 10.6151
R1292 B.n487 B.n132 10.6151
R1293 B.n488 B.n487 10.6151
R1294 B.n489 B.n488 10.6151
R1295 B.n489 B.n130 10.6151
R1296 B.n493 B.n130 10.6151
R1297 B.n494 B.n493 10.6151
R1298 B.n495 B.n494 10.6151
R1299 B.n495 B.n128 10.6151
R1300 B.n499 B.n128 10.6151
R1301 B.n500 B.n499 10.6151
R1302 B.n501 B.n500 10.6151
R1303 B.n501 B.n126 10.6151
R1304 B.n505 B.n126 10.6151
R1305 B.n506 B.n505 10.6151
R1306 B.n507 B.n506 10.6151
R1307 B.n507 B.n124 10.6151
R1308 B.n511 B.n124 10.6151
R1309 B.n512 B.n511 10.6151
R1310 B.n513 B.n512 10.6151
R1311 B.n513 B.n122 10.6151
R1312 B.n517 B.n122 10.6151
R1313 B.n518 B.n517 10.6151
R1314 B.n519 B.n518 10.6151
R1315 B.n519 B.n120 10.6151
R1316 B.n523 B.n120 10.6151
R1317 B.n524 B.n523 10.6151
R1318 B.n525 B.n524 10.6151
R1319 B.n525 B.n118 10.6151
R1320 B.n529 B.n118 10.6151
R1321 B.n530 B.n529 10.6151
R1322 B.n531 B.n530 10.6151
R1323 B.n531 B.n116 10.6151
R1324 B.n535 B.n116 10.6151
R1325 B.n536 B.n535 10.6151
R1326 B.n537 B.n536 10.6151
R1327 B.n537 B.n114 10.6151
R1328 B.n541 B.n114 10.6151
R1329 B.n542 B.n541 10.6151
R1330 B.n543 B.n542 10.6151
R1331 B.n543 B.n112 10.6151
R1332 B.n547 B.n112 10.6151
R1333 B.n548 B.n547 10.6151
R1334 B.n549 B.n548 10.6151
R1335 B.n549 B.n110 10.6151
R1336 B.n553 B.n110 10.6151
R1337 B.n554 B.n553 10.6151
R1338 B.n555 B.n554 10.6151
R1339 B.n555 B.n108 10.6151
R1340 B.n559 B.n108 10.6151
R1341 B.n560 B.n559 10.6151
R1342 B.n561 B.n560 10.6151
R1343 B.n561 B.n106 10.6151
R1344 B.n565 B.n106 10.6151
R1345 B.n566 B.n565 10.6151
R1346 B.n567 B.n566 10.6151
R1347 B.n567 B.n104 10.6151
R1348 B.n571 B.n104 10.6151
R1349 B.n572 B.n571 10.6151
R1350 B.n573 B.n572 10.6151
R1351 B.n573 B.n102 10.6151
R1352 B.n577 B.n102 10.6151
R1353 B.n578 B.n577 10.6151
R1354 B.n579 B.n578 10.6151
R1355 B.n579 B.n100 10.6151
R1356 B.n583 B.n100 10.6151
R1357 B.n584 B.n583 10.6151
R1358 B.n585 B.n584 10.6151
R1359 B.n585 B.n98 10.6151
R1360 B.n589 B.n98 10.6151
R1361 B.n590 B.n589 10.6151
R1362 B.n591 B.n590 10.6151
R1363 B.n591 B.n96 10.6151
R1364 B.n595 B.n96 10.6151
R1365 B.n596 B.n595 10.6151
R1366 B.n597 B.n596 10.6151
R1367 B.n597 B.n94 10.6151
R1368 B.n601 B.n94 10.6151
R1369 B.n602 B.n601 10.6151
R1370 B.n603 B.n602 10.6151
R1371 B.n603 B.n92 10.6151
R1372 B.n607 B.n92 10.6151
R1373 B.n608 B.n607 10.6151
R1374 B.n609 B.n608 10.6151
R1375 B.n609 B.n90 10.6151
R1376 B.n613 B.n90 10.6151
R1377 B.n614 B.n613 10.6151
R1378 B.n615 B.n614 10.6151
R1379 B.n615 B.n88 10.6151
R1380 B.n619 B.n88 10.6151
R1381 B.n620 B.n619 10.6151
R1382 B.n621 B.n620 10.6151
R1383 B.n621 B.n86 10.6151
R1384 B.n625 B.n86 10.6151
R1385 B.n626 B.n625 10.6151
R1386 B.n627 B.n626 10.6151
R1387 B.n627 B.n84 10.6151
R1388 B.n631 B.n84 10.6151
R1389 B.n632 B.n631 10.6151
R1390 B.n633 B.n632 10.6151
R1391 B.n633 B.n82 10.6151
R1392 B.n637 B.n82 10.6151
R1393 B.n638 B.n637 10.6151
R1394 B.n319 B.n192 10.6151
R1395 B.n320 B.n319 10.6151
R1396 B.n321 B.n320 10.6151
R1397 B.n321 B.n190 10.6151
R1398 B.n325 B.n190 10.6151
R1399 B.n326 B.n325 10.6151
R1400 B.n327 B.n326 10.6151
R1401 B.n327 B.n188 10.6151
R1402 B.n331 B.n188 10.6151
R1403 B.n332 B.n331 10.6151
R1404 B.n333 B.n332 10.6151
R1405 B.n333 B.n186 10.6151
R1406 B.n337 B.n186 10.6151
R1407 B.n338 B.n337 10.6151
R1408 B.n339 B.n338 10.6151
R1409 B.n339 B.n184 10.6151
R1410 B.n343 B.n184 10.6151
R1411 B.n344 B.n343 10.6151
R1412 B.n345 B.n344 10.6151
R1413 B.n345 B.n182 10.6151
R1414 B.n349 B.n182 10.6151
R1415 B.n350 B.n349 10.6151
R1416 B.n351 B.n350 10.6151
R1417 B.n351 B.n180 10.6151
R1418 B.n355 B.n180 10.6151
R1419 B.n356 B.n355 10.6151
R1420 B.n357 B.n356 10.6151
R1421 B.n357 B.n178 10.6151
R1422 B.n361 B.n178 10.6151
R1423 B.n362 B.n361 10.6151
R1424 B.n363 B.n362 10.6151
R1425 B.n363 B.n176 10.6151
R1426 B.n367 B.n176 10.6151
R1427 B.n368 B.n367 10.6151
R1428 B.n369 B.n368 10.6151
R1429 B.n369 B.n174 10.6151
R1430 B.n373 B.n174 10.6151
R1431 B.n374 B.n373 10.6151
R1432 B.n376 B.n170 10.6151
R1433 B.n380 B.n170 10.6151
R1434 B.n381 B.n380 10.6151
R1435 B.n382 B.n381 10.6151
R1436 B.n382 B.n168 10.6151
R1437 B.n386 B.n168 10.6151
R1438 B.n387 B.n386 10.6151
R1439 B.n388 B.n387 10.6151
R1440 B.n392 B.n391 10.6151
R1441 B.n393 B.n392 10.6151
R1442 B.n393 B.n162 10.6151
R1443 B.n397 B.n162 10.6151
R1444 B.n398 B.n397 10.6151
R1445 B.n399 B.n398 10.6151
R1446 B.n399 B.n160 10.6151
R1447 B.n403 B.n160 10.6151
R1448 B.n404 B.n403 10.6151
R1449 B.n405 B.n404 10.6151
R1450 B.n405 B.n158 10.6151
R1451 B.n409 B.n158 10.6151
R1452 B.n410 B.n409 10.6151
R1453 B.n411 B.n410 10.6151
R1454 B.n411 B.n156 10.6151
R1455 B.n415 B.n156 10.6151
R1456 B.n416 B.n415 10.6151
R1457 B.n417 B.n416 10.6151
R1458 B.n417 B.n154 10.6151
R1459 B.n421 B.n154 10.6151
R1460 B.n422 B.n421 10.6151
R1461 B.n423 B.n422 10.6151
R1462 B.n423 B.n152 10.6151
R1463 B.n427 B.n152 10.6151
R1464 B.n428 B.n427 10.6151
R1465 B.n429 B.n428 10.6151
R1466 B.n429 B.n150 10.6151
R1467 B.n433 B.n150 10.6151
R1468 B.n434 B.n433 10.6151
R1469 B.n435 B.n434 10.6151
R1470 B.n435 B.n148 10.6151
R1471 B.n439 B.n148 10.6151
R1472 B.n440 B.n439 10.6151
R1473 B.n441 B.n440 10.6151
R1474 B.n441 B.n146 10.6151
R1475 B.n445 B.n146 10.6151
R1476 B.n446 B.n445 10.6151
R1477 B.n447 B.n446 10.6151
R1478 B.n315 B.n314 10.6151
R1479 B.n314 B.n313 10.6151
R1480 B.n313 B.n194 10.6151
R1481 B.n309 B.n194 10.6151
R1482 B.n309 B.n308 10.6151
R1483 B.n308 B.n307 10.6151
R1484 B.n307 B.n196 10.6151
R1485 B.n303 B.n196 10.6151
R1486 B.n303 B.n302 10.6151
R1487 B.n302 B.n301 10.6151
R1488 B.n301 B.n198 10.6151
R1489 B.n297 B.n198 10.6151
R1490 B.n297 B.n296 10.6151
R1491 B.n296 B.n295 10.6151
R1492 B.n295 B.n200 10.6151
R1493 B.n291 B.n200 10.6151
R1494 B.n291 B.n290 10.6151
R1495 B.n290 B.n289 10.6151
R1496 B.n289 B.n202 10.6151
R1497 B.n285 B.n202 10.6151
R1498 B.n285 B.n284 10.6151
R1499 B.n284 B.n283 10.6151
R1500 B.n283 B.n204 10.6151
R1501 B.n279 B.n204 10.6151
R1502 B.n279 B.n278 10.6151
R1503 B.n278 B.n277 10.6151
R1504 B.n277 B.n206 10.6151
R1505 B.n273 B.n206 10.6151
R1506 B.n273 B.n272 10.6151
R1507 B.n272 B.n271 10.6151
R1508 B.n271 B.n208 10.6151
R1509 B.n267 B.n208 10.6151
R1510 B.n267 B.n266 10.6151
R1511 B.n266 B.n265 10.6151
R1512 B.n265 B.n210 10.6151
R1513 B.n261 B.n210 10.6151
R1514 B.n261 B.n260 10.6151
R1515 B.n260 B.n259 10.6151
R1516 B.n259 B.n212 10.6151
R1517 B.n255 B.n212 10.6151
R1518 B.n255 B.n254 10.6151
R1519 B.n254 B.n253 10.6151
R1520 B.n253 B.n214 10.6151
R1521 B.n249 B.n214 10.6151
R1522 B.n249 B.n248 10.6151
R1523 B.n248 B.n247 10.6151
R1524 B.n247 B.n216 10.6151
R1525 B.n243 B.n216 10.6151
R1526 B.n243 B.n242 10.6151
R1527 B.n242 B.n241 10.6151
R1528 B.n241 B.n218 10.6151
R1529 B.n237 B.n218 10.6151
R1530 B.n237 B.n236 10.6151
R1531 B.n236 B.n235 10.6151
R1532 B.n235 B.n220 10.6151
R1533 B.n231 B.n220 10.6151
R1534 B.n231 B.n230 10.6151
R1535 B.n230 B.n229 10.6151
R1536 B.n229 B.n222 10.6151
R1537 B.n225 B.n222 10.6151
R1538 B.n225 B.n224 10.6151
R1539 B.n224 B.n0 10.6151
R1540 B.n863 B.n1 10.6151
R1541 B.n863 B.n862 10.6151
R1542 B.n862 B.n861 10.6151
R1543 B.n861 B.n4 10.6151
R1544 B.n857 B.n4 10.6151
R1545 B.n857 B.n856 10.6151
R1546 B.n856 B.n855 10.6151
R1547 B.n855 B.n6 10.6151
R1548 B.n851 B.n6 10.6151
R1549 B.n851 B.n850 10.6151
R1550 B.n850 B.n849 10.6151
R1551 B.n849 B.n8 10.6151
R1552 B.n845 B.n8 10.6151
R1553 B.n845 B.n844 10.6151
R1554 B.n844 B.n843 10.6151
R1555 B.n843 B.n10 10.6151
R1556 B.n839 B.n10 10.6151
R1557 B.n839 B.n838 10.6151
R1558 B.n838 B.n837 10.6151
R1559 B.n837 B.n12 10.6151
R1560 B.n833 B.n12 10.6151
R1561 B.n833 B.n832 10.6151
R1562 B.n832 B.n831 10.6151
R1563 B.n831 B.n14 10.6151
R1564 B.n827 B.n14 10.6151
R1565 B.n827 B.n826 10.6151
R1566 B.n826 B.n825 10.6151
R1567 B.n825 B.n16 10.6151
R1568 B.n821 B.n16 10.6151
R1569 B.n821 B.n820 10.6151
R1570 B.n820 B.n819 10.6151
R1571 B.n819 B.n18 10.6151
R1572 B.n815 B.n18 10.6151
R1573 B.n815 B.n814 10.6151
R1574 B.n814 B.n813 10.6151
R1575 B.n813 B.n20 10.6151
R1576 B.n809 B.n20 10.6151
R1577 B.n809 B.n808 10.6151
R1578 B.n808 B.n807 10.6151
R1579 B.n807 B.n22 10.6151
R1580 B.n803 B.n22 10.6151
R1581 B.n803 B.n802 10.6151
R1582 B.n802 B.n801 10.6151
R1583 B.n801 B.n24 10.6151
R1584 B.n797 B.n24 10.6151
R1585 B.n797 B.n796 10.6151
R1586 B.n796 B.n795 10.6151
R1587 B.n795 B.n26 10.6151
R1588 B.n791 B.n26 10.6151
R1589 B.n791 B.n790 10.6151
R1590 B.n790 B.n789 10.6151
R1591 B.n789 B.n28 10.6151
R1592 B.n785 B.n28 10.6151
R1593 B.n785 B.n784 10.6151
R1594 B.n784 B.n783 10.6151
R1595 B.n783 B.n30 10.6151
R1596 B.n779 B.n30 10.6151
R1597 B.n779 B.n778 10.6151
R1598 B.n778 B.n777 10.6151
R1599 B.n777 B.n32 10.6151
R1600 B.n773 B.n32 10.6151
R1601 B.n773 B.n772 10.6151
R1602 B.n712 B.n711 6.5566
R1603 B.n699 B.n698 6.5566
R1604 B.n376 B.n375 6.5566
R1605 B.n388 B.n166 6.5566
R1606 B.n713 B.n712 4.05904
R1607 B.n698 B.n697 4.05904
R1608 B.n375 B.n374 4.05904
R1609 B.n391 B.n166 4.05904
R1610 B.n867 B.n0 2.81026
R1611 B.n867 B.n1 2.81026
C0 w_n4700_n3166# VTAIL 4.06394f
C1 VDD2 B 1.98739f
C2 VN w_n4700_n3166# 9.76532f
C3 w_n4700_n3166# VP 10.377799f
C4 VN VTAIL 9.08948f
C5 VTAIL VP 9.10358f
C6 VN VP 8.45191f
C7 VDD1 w_n4700_n3166# 2.17894f
C8 VDD1 VTAIL 8.08034f
C9 VDD1 VN 0.152777f
C10 VDD1 VP 8.83934f
C11 VDD2 w_n4700_n3166# 2.3272f
C12 w_n4700_n3166# B 11.0568f
C13 VDD2 VTAIL 8.140121f
C14 VDD2 VN 8.389519f
C15 VDD2 VP 0.604402f
C16 B VTAIL 4.97609f
C17 VN B 1.39959f
C18 B VP 2.43065f
C19 VDD1 VDD2 2.1888f
C20 VDD1 B 1.8662f
C21 VDD2 VSUBS 2.244349f
C22 VDD1 VSUBS 3.03802f
C23 VTAIL VSUBS 1.438938f
C24 VN VSUBS 7.79858f
C25 VP VSUBS 4.378336f
C26 B VSUBS 5.810103f
C27 w_n4700_n3166# VSUBS 0.183469p
C28 B.n0 VSUBS 0.004748f
C29 B.n1 VSUBS 0.004748f
C30 B.n2 VSUBS 0.007509f
C31 B.n3 VSUBS 0.007509f
C32 B.n4 VSUBS 0.007509f
C33 B.n5 VSUBS 0.007509f
C34 B.n6 VSUBS 0.007509f
C35 B.n7 VSUBS 0.007509f
C36 B.n8 VSUBS 0.007509f
C37 B.n9 VSUBS 0.007509f
C38 B.n10 VSUBS 0.007509f
C39 B.n11 VSUBS 0.007509f
C40 B.n12 VSUBS 0.007509f
C41 B.n13 VSUBS 0.007509f
C42 B.n14 VSUBS 0.007509f
C43 B.n15 VSUBS 0.007509f
C44 B.n16 VSUBS 0.007509f
C45 B.n17 VSUBS 0.007509f
C46 B.n18 VSUBS 0.007509f
C47 B.n19 VSUBS 0.007509f
C48 B.n20 VSUBS 0.007509f
C49 B.n21 VSUBS 0.007509f
C50 B.n22 VSUBS 0.007509f
C51 B.n23 VSUBS 0.007509f
C52 B.n24 VSUBS 0.007509f
C53 B.n25 VSUBS 0.007509f
C54 B.n26 VSUBS 0.007509f
C55 B.n27 VSUBS 0.007509f
C56 B.n28 VSUBS 0.007509f
C57 B.n29 VSUBS 0.007509f
C58 B.n30 VSUBS 0.007509f
C59 B.n31 VSUBS 0.007509f
C60 B.n32 VSUBS 0.007509f
C61 B.n33 VSUBS 0.016654f
C62 B.n34 VSUBS 0.007509f
C63 B.n35 VSUBS 0.007509f
C64 B.n36 VSUBS 0.007509f
C65 B.n37 VSUBS 0.007509f
C66 B.n38 VSUBS 0.007509f
C67 B.n39 VSUBS 0.007509f
C68 B.n40 VSUBS 0.007509f
C69 B.n41 VSUBS 0.007509f
C70 B.n42 VSUBS 0.007509f
C71 B.n43 VSUBS 0.007509f
C72 B.n44 VSUBS 0.007509f
C73 B.n45 VSUBS 0.007509f
C74 B.n46 VSUBS 0.007509f
C75 B.n47 VSUBS 0.007509f
C76 B.n48 VSUBS 0.007509f
C77 B.n49 VSUBS 0.007509f
C78 B.n50 VSUBS 0.007509f
C79 B.n51 VSUBS 0.007509f
C80 B.n52 VSUBS 0.007509f
C81 B.n53 VSUBS 0.007509f
C82 B.t8 VSUBS 0.380391f
C83 B.t7 VSUBS 0.408151f
C84 B.t6 VSUBS 1.86608f
C85 B.n54 VSUBS 0.227619f
C86 B.n55 VSUBS 0.080482f
C87 B.n56 VSUBS 0.007509f
C88 B.n57 VSUBS 0.007509f
C89 B.n58 VSUBS 0.007509f
C90 B.n59 VSUBS 0.007509f
C91 B.t2 VSUBS 0.380385f
C92 B.t1 VSUBS 0.408146f
C93 B.t0 VSUBS 1.86608f
C94 B.n60 VSUBS 0.227624f
C95 B.n61 VSUBS 0.080489f
C96 B.n62 VSUBS 0.007509f
C97 B.n63 VSUBS 0.007509f
C98 B.n64 VSUBS 0.007509f
C99 B.n65 VSUBS 0.007509f
C100 B.n66 VSUBS 0.007509f
C101 B.n67 VSUBS 0.007509f
C102 B.n68 VSUBS 0.007509f
C103 B.n69 VSUBS 0.007509f
C104 B.n70 VSUBS 0.007509f
C105 B.n71 VSUBS 0.007509f
C106 B.n72 VSUBS 0.007509f
C107 B.n73 VSUBS 0.007509f
C108 B.n74 VSUBS 0.007509f
C109 B.n75 VSUBS 0.007509f
C110 B.n76 VSUBS 0.007509f
C111 B.n77 VSUBS 0.007509f
C112 B.n78 VSUBS 0.007509f
C113 B.n79 VSUBS 0.007509f
C114 B.n80 VSUBS 0.007509f
C115 B.n81 VSUBS 0.016654f
C116 B.n82 VSUBS 0.007509f
C117 B.n83 VSUBS 0.007509f
C118 B.n84 VSUBS 0.007509f
C119 B.n85 VSUBS 0.007509f
C120 B.n86 VSUBS 0.007509f
C121 B.n87 VSUBS 0.007509f
C122 B.n88 VSUBS 0.007509f
C123 B.n89 VSUBS 0.007509f
C124 B.n90 VSUBS 0.007509f
C125 B.n91 VSUBS 0.007509f
C126 B.n92 VSUBS 0.007509f
C127 B.n93 VSUBS 0.007509f
C128 B.n94 VSUBS 0.007509f
C129 B.n95 VSUBS 0.007509f
C130 B.n96 VSUBS 0.007509f
C131 B.n97 VSUBS 0.007509f
C132 B.n98 VSUBS 0.007509f
C133 B.n99 VSUBS 0.007509f
C134 B.n100 VSUBS 0.007509f
C135 B.n101 VSUBS 0.007509f
C136 B.n102 VSUBS 0.007509f
C137 B.n103 VSUBS 0.007509f
C138 B.n104 VSUBS 0.007509f
C139 B.n105 VSUBS 0.007509f
C140 B.n106 VSUBS 0.007509f
C141 B.n107 VSUBS 0.007509f
C142 B.n108 VSUBS 0.007509f
C143 B.n109 VSUBS 0.007509f
C144 B.n110 VSUBS 0.007509f
C145 B.n111 VSUBS 0.007509f
C146 B.n112 VSUBS 0.007509f
C147 B.n113 VSUBS 0.007509f
C148 B.n114 VSUBS 0.007509f
C149 B.n115 VSUBS 0.007509f
C150 B.n116 VSUBS 0.007509f
C151 B.n117 VSUBS 0.007509f
C152 B.n118 VSUBS 0.007509f
C153 B.n119 VSUBS 0.007509f
C154 B.n120 VSUBS 0.007509f
C155 B.n121 VSUBS 0.007509f
C156 B.n122 VSUBS 0.007509f
C157 B.n123 VSUBS 0.007509f
C158 B.n124 VSUBS 0.007509f
C159 B.n125 VSUBS 0.007509f
C160 B.n126 VSUBS 0.007509f
C161 B.n127 VSUBS 0.007509f
C162 B.n128 VSUBS 0.007509f
C163 B.n129 VSUBS 0.007509f
C164 B.n130 VSUBS 0.007509f
C165 B.n131 VSUBS 0.007509f
C166 B.n132 VSUBS 0.007509f
C167 B.n133 VSUBS 0.007509f
C168 B.n134 VSUBS 0.007509f
C169 B.n135 VSUBS 0.007509f
C170 B.n136 VSUBS 0.007509f
C171 B.n137 VSUBS 0.007509f
C172 B.n138 VSUBS 0.007509f
C173 B.n139 VSUBS 0.007509f
C174 B.n140 VSUBS 0.007509f
C175 B.n141 VSUBS 0.007509f
C176 B.n142 VSUBS 0.007509f
C177 B.n143 VSUBS 0.007509f
C178 B.n144 VSUBS 0.016654f
C179 B.n145 VSUBS 0.007509f
C180 B.n146 VSUBS 0.007509f
C181 B.n147 VSUBS 0.007509f
C182 B.n148 VSUBS 0.007509f
C183 B.n149 VSUBS 0.007509f
C184 B.n150 VSUBS 0.007509f
C185 B.n151 VSUBS 0.007509f
C186 B.n152 VSUBS 0.007509f
C187 B.n153 VSUBS 0.007509f
C188 B.n154 VSUBS 0.007509f
C189 B.n155 VSUBS 0.007509f
C190 B.n156 VSUBS 0.007509f
C191 B.n157 VSUBS 0.007509f
C192 B.n158 VSUBS 0.007509f
C193 B.n159 VSUBS 0.007509f
C194 B.n160 VSUBS 0.007509f
C195 B.n161 VSUBS 0.007509f
C196 B.n162 VSUBS 0.007509f
C197 B.n163 VSUBS 0.007509f
C198 B.t10 VSUBS 0.380385f
C199 B.t11 VSUBS 0.408146f
C200 B.t9 VSUBS 1.86608f
C201 B.n164 VSUBS 0.227624f
C202 B.n165 VSUBS 0.080489f
C203 B.n166 VSUBS 0.017397f
C204 B.n167 VSUBS 0.007509f
C205 B.n168 VSUBS 0.007509f
C206 B.n169 VSUBS 0.007509f
C207 B.n170 VSUBS 0.007509f
C208 B.n171 VSUBS 0.007509f
C209 B.t4 VSUBS 0.380391f
C210 B.t5 VSUBS 0.408151f
C211 B.t3 VSUBS 1.86608f
C212 B.n172 VSUBS 0.227619f
C213 B.n173 VSUBS 0.080482f
C214 B.n174 VSUBS 0.007509f
C215 B.n175 VSUBS 0.007509f
C216 B.n176 VSUBS 0.007509f
C217 B.n177 VSUBS 0.007509f
C218 B.n178 VSUBS 0.007509f
C219 B.n179 VSUBS 0.007509f
C220 B.n180 VSUBS 0.007509f
C221 B.n181 VSUBS 0.007509f
C222 B.n182 VSUBS 0.007509f
C223 B.n183 VSUBS 0.007509f
C224 B.n184 VSUBS 0.007509f
C225 B.n185 VSUBS 0.007509f
C226 B.n186 VSUBS 0.007509f
C227 B.n187 VSUBS 0.007509f
C228 B.n188 VSUBS 0.007509f
C229 B.n189 VSUBS 0.007509f
C230 B.n190 VSUBS 0.007509f
C231 B.n191 VSUBS 0.007509f
C232 B.n192 VSUBS 0.017577f
C233 B.n193 VSUBS 0.007509f
C234 B.n194 VSUBS 0.007509f
C235 B.n195 VSUBS 0.007509f
C236 B.n196 VSUBS 0.007509f
C237 B.n197 VSUBS 0.007509f
C238 B.n198 VSUBS 0.007509f
C239 B.n199 VSUBS 0.007509f
C240 B.n200 VSUBS 0.007509f
C241 B.n201 VSUBS 0.007509f
C242 B.n202 VSUBS 0.007509f
C243 B.n203 VSUBS 0.007509f
C244 B.n204 VSUBS 0.007509f
C245 B.n205 VSUBS 0.007509f
C246 B.n206 VSUBS 0.007509f
C247 B.n207 VSUBS 0.007509f
C248 B.n208 VSUBS 0.007509f
C249 B.n209 VSUBS 0.007509f
C250 B.n210 VSUBS 0.007509f
C251 B.n211 VSUBS 0.007509f
C252 B.n212 VSUBS 0.007509f
C253 B.n213 VSUBS 0.007509f
C254 B.n214 VSUBS 0.007509f
C255 B.n215 VSUBS 0.007509f
C256 B.n216 VSUBS 0.007509f
C257 B.n217 VSUBS 0.007509f
C258 B.n218 VSUBS 0.007509f
C259 B.n219 VSUBS 0.007509f
C260 B.n220 VSUBS 0.007509f
C261 B.n221 VSUBS 0.007509f
C262 B.n222 VSUBS 0.007509f
C263 B.n223 VSUBS 0.007509f
C264 B.n224 VSUBS 0.007509f
C265 B.n225 VSUBS 0.007509f
C266 B.n226 VSUBS 0.007509f
C267 B.n227 VSUBS 0.007509f
C268 B.n228 VSUBS 0.007509f
C269 B.n229 VSUBS 0.007509f
C270 B.n230 VSUBS 0.007509f
C271 B.n231 VSUBS 0.007509f
C272 B.n232 VSUBS 0.007509f
C273 B.n233 VSUBS 0.007509f
C274 B.n234 VSUBS 0.007509f
C275 B.n235 VSUBS 0.007509f
C276 B.n236 VSUBS 0.007509f
C277 B.n237 VSUBS 0.007509f
C278 B.n238 VSUBS 0.007509f
C279 B.n239 VSUBS 0.007509f
C280 B.n240 VSUBS 0.007509f
C281 B.n241 VSUBS 0.007509f
C282 B.n242 VSUBS 0.007509f
C283 B.n243 VSUBS 0.007509f
C284 B.n244 VSUBS 0.007509f
C285 B.n245 VSUBS 0.007509f
C286 B.n246 VSUBS 0.007509f
C287 B.n247 VSUBS 0.007509f
C288 B.n248 VSUBS 0.007509f
C289 B.n249 VSUBS 0.007509f
C290 B.n250 VSUBS 0.007509f
C291 B.n251 VSUBS 0.007509f
C292 B.n252 VSUBS 0.007509f
C293 B.n253 VSUBS 0.007509f
C294 B.n254 VSUBS 0.007509f
C295 B.n255 VSUBS 0.007509f
C296 B.n256 VSUBS 0.007509f
C297 B.n257 VSUBS 0.007509f
C298 B.n258 VSUBS 0.007509f
C299 B.n259 VSUBS 0.007509f
C300 B.n260 VSUBS 0.007509f
C301 B.n261 VSUBS 0.007509f
C302 B.n262 VSUBS 0.007509f
C303 B.n263 VSUBS 0.007509f
C304 B.n264 VSUBS 0.007509f
C305 B.n265 VSUBS 0.007509f
C306 B.n266 VSUBS 0.007509f
C307 B.n267 VSUBS 0.007509f
C308 B.n268 VSUBS 0.007509f
C309 B.n269 VSUBS 0.007509f
C310 B.n270 VSUBS 0.007509f
C311 B.n271 VSUBS 0.007509f
C312 B.n272 VSUBS 0.007509f
C313 B.n273 VSUBS 0.007509f
C314 B.n274 VSUBS 0.007509f
C315 B.n275 VSUBS 0.007509f
C316 B.n276 VSUBS 0.007509f
C317 B.n277 VSUBS 0.007509f
C318 B.n278 VSUBS 0.007509f
C319 B.n279 VSUBS 0.007509f
C320 B.n280 VSUBS 0.007509f
C321 B.n281 VSUBS 0.007509f
C322 B.n282 VSUBS 0.007509f
C323 B.n283 VSUBS 0.007509f
C324 B.n284 VSUBS 0.007509f
C325 B.n285 VSUBS 0.007509f
C326 B.n286 VSUBS 0.007509f
C327 B.n287 VSUBS 0.007509f
C328 B.n288 VSUBS 0.007509f
C329 B.n289 VSUBS 0.007509f
C330 B.n290 VSUBS 0.007509f
C331 B.n291 VSUBS 0.007509f
C332 B.n292 VSUBS 0.007509f
C333 B.n293 VSUBS 0.007509f
C334 B.n294 VSUBS 0.007509f
C335 B.n295 VSUBS 0.007509f
C336 B.n296 VSUBS 0.007509f
C337 B.n297 VSUBS 0.007509f
C338 B.n298 VSUBS 0.007509f
C339 B.n299 VSUBS 0.007509f
C340 B.n300 VSUBS 0.007509f
C341 B.n301 VSUBS 0.007509f
C342 B.n302 VSUBS 0.007509f
C343 B.n303 VSUBS 0.007509f
C344 B.n304 VSUBS 0.007509f
C345 B.n305 VSUBS 0.007509f
C346 B.n306 VSUBS 0.007509f
C347 B.n307 VSUBS 0.007509f
C348 B.n308 VSUBS 0.007509f
C349 B.n309 VSUBS 0.007509f
C350 B.n310 VSUBS 0.007509f
C351 B.n311 VSUBS 0.007509f
C352 B.n312 VSUBS 0.007509f
C353 B.n313 VSUBS 0.007509f
C354 B.n314 VSUBS 0.007509f
C355 B.n315 VSUBS 0.016654f
C356 B.n316 VSUBS 0.016654f
C357 B.n317 VSUBS 0.017577f
C358 B.n318 VSUBS 0.007509f
C359 B.n319 VSUBS 0.007509f
C360 B.n320 VSUBS 0.007509f
C361 B.n321 VSUBS 0.007509f
C362 B.n322 VSUBS 0.007509f
C363 B.n323 VSUBS 0.007509f
C364 B.n324 VSUBS 0.007509f
C365 B.n325 VSUBS 0.007509f
C366 B.n326 VSUBS 0.007509f
C367 B.n327 VSUBS 0.007509f
C368 B.n328 VSUBS 0.007509f
C369 B.n329 VSUBS 0.007509f
C370 B.n330 VSUBS 0.007509f
C371 B.n331 VSUBS 0.007509f
C372 B.n332 VSUBS 0.007509f
C373 B.n333 VSUBS 0.007509f
C374 B.n334 VSUBS 0.007509f
C375 B.n335 VSUBS 0.007509f
C376 B.n336 VSUBS 0.007509f
C377 B.n337 VSUBS 0.007509f
C378 B.n338 VSUBS 0.007509f
C379 B.n339 VSUBS 0.007509f
C380 B.n340 VSUBS 0.007509f
C381 B.n341 VSUBS 0.007509f
C382 B.n342 VSUBS 0.007509f
C383 B.n343 VSUBS 0.007509f
C384 B.n344 VSUBS 0.007509f
C385 B.n345 VSUBS 0.007509f
C386 B.n346 VSUBS 0.007509f
C387 B.n347 VSUBS 0.007509f
C388 B.n348 VSUBS 0.007509f
C389 B.n349 VSUBS 0.007509f
C390 B.n350 VSUBS 0.007509f
C391 B.n351 VSUBS 0.007509f
C392 B.n352 VSUBS 0.007509f
C393 B.n353 VSUBS 0.007509f
C394 B.n354 VSUBS 0.007509f
C395 B.n355 VSUBS 0.007509f
C396 B.n356 VSUBS 0.007509f
C397 B.n357 VSUBS 0.007509f
C398 B.n358 VSUBS 0.007509f
C399 B.n359 VSUBS 0.007509f
C400 B.n360 VSUBS 0.007509f
C401 B.n361 VSUBS 0.007509f
C402 B.n362 VSUBS 0.007509f
C403 B.n363 VSUBS 0.007509f
C404 B.n364 VSUBS 0.007509f
C405 B.n365 VSUBS 0.007509f
C406 B.n366 VSUBS 0.007509f
C407 B.n367 VSUBS 0.007509f
C408 B.n368 VSUBS 0.007509f
C409 B.n369 VSUBS 0.007509f
C410 B.n370 VSUBS 0.007509f
C411 B.n371 VSUBS 0.007509f
C412 B.n372 VSUBS 0.007509f
C413 B.n373 VSUBS 0.007509f
C414 B.n374 VSUBS 0.00519f
C415 B.n375 VSUBS 0.017397f
C416 B.n376 VSUBS 0.006073f
C417 B.n377 VSUBS 0.007509f
C418 B.n378 VSUBS 0.007509f
C419 B.n379 VSUBS 0.007509f
C420 B.n380 VSUBS 0.007509f
C421 B.n381 VSUBS 0.007509f
C422 B.n382 VSUBS 0.007509f
C423 B.n383 VSUBS 0.007509f
C424 B.n384 VSUBS 0.007509f
C425 B.n385 VSUBS 0.007509f
C426 B.n386 VSUBS 0.007509f
C427 B.n387 VSUBS 0.007509f
C428 B.n388 VSUBS 0.006073f
C429 B.n389 VSUBS 0.007509f
C430 B.n390 VSUBS 0.007509f
C431 B.n391 VSUBS 0.00519f
C432 B.n392 VSUBS 0.007509f
C433 B.n393 VSUBS 0.007509f
C434 B.n394 VSUBS 0.007509f
C435 B.n395 VSUBS 0.007509f
C436 B.n396 VSUBS 0.007509f
C437 B.n397 VSUBS 0.007509f
C438 B.n398 VSUBS 0.007509f
C439 B.n399 VSUBS 0.007509f
C440 B.n400 VSUBS 0.007509f
C441 B.n401 VSUBS 0.007509f
C442 B.n402 VSUBS 0.007509f
C443 B.n403 VSUBS 0.007509f
C444 B.n404 VSUBS 0.007509f
C445 B.n405 VSUBS 0.007509f
C446 B.n406 VSUBS 0.007509f
C447 B.n407 VSUBS 0.007509f
C448 B.n408 VSUBS 0.007509f
C449 B.n409 VSUBS 0.007509f
C450 B.n410 VSUBS 0.007509f
C451 B.n411 VSUBS 0.007509f
C452 B.n412 VSUBS 0.007509f
C453 B.n413 VSUBS 0.007509f
C454 B.n414 VSUBS 0.007509f
C455 B.n415 VSUBS 0.007509f
C456 B.n416 VSUBS 0.007509f
C457 B.n417 VSUBS 0.007509f
C458 B.n418 VSUBS 0.007509f
C459 B.n419 VSUBS 0.007509f
C460 B.n420 VSUBS 0.007509f
C461 B.n421 VSUBS 0.007509f
C462 B.n422 VSUBS 0.007509f
C463 B.n423 VSUBS 0.007509f
C464 B.n424 VSUBS 0.007509f
C465 B.n425 VSUBS 0.007509f
C466 B.n426 VSUBS 0.007509f
C467 B.n427 VSUBS 0.007509f
C468 B.n428 VSUBS 0.007509f
C469 B.n429 VSUBS 0.007509f
C470 B.n430 VSUBS 0.007509f
C471 B.n431 VSUBS 0.007509f
C472 B.n432 VSUBS 0.007509f
C473 B.n433 VSUBS 0.007509f
C474 B.n434 VSUBS 0.007509f
C475 B.n435 VSUBS 0.007509f
C476 B.n436 VSUBS 0.007509f
C477 B.n437 VSUBS 0.007509f
C478 B.n438 VSUBS 0.007509f
C479 B.n439 VSUBS 0.007509f
C480 B.n440 VSUBS 0.007509f
C481 B.n441 VSUBS 0.007509f
C482 B.n442 VSUBS 0.007509f
C483 B.n443 VSUBS 0.007509f
C484 B.n444 VSUBS 0.007509f
C485 B.n445 VSUBS 0.007509f
C486 B.n446 VSUBS 0.007509f
C487 B.n447 VSUBS 0.017577f
C488 B.n448 VSUBS 0.017577f
C489 B.n449 VSUBS 0.016654f
C490 B.n450 VSUBS 0.007509f
C491 B.n451 VSUBS 0.007509f
C492 B.n452 VSUBS 0.007509f
C493 B.n453 VSUBS 0.007509f
C494 B.n454 VSUBS 0.007509f
C495 B.n455 VSUBS 0.007509f
C496 B.n456 VSUBS 0.007509f
C497 B.n457 VSUBS 0.007509f
C498 B.n458 VSUBS 0.007509f
C499 B.n459 VSUBS 0.007509f
C500 B.n460 VSUBS 0.007509f
C501 B.n461 VSUBS 0.007509f
C502 B.n462 VSUBS 0.007509f
C503 B.n463 VSUBS 0.007509f
C504 B.n464 VSUBS 0.007509f
C505 B.n465 VSUBS 0.007509f
C506 B.n466 VSUBS 0.007509f
C507 B.n467 VSUBS 0.007509f
C508 B.n468 VSUBS 0.007509f
C509 B.n469 VSUBS 0.007509f
C510 B.n470 VSUBS 0.007509f
C511 B.n471 VSUBS 0.007509f
C512 B.n472 VSUBS 0.007509f
C513 B.n473 VSUBS 0.007509f
C514 B.n474 VSUBS 0.007509f
C515 B.n475 VSUBS 0.007509f
C516 B.n476 VSUBS 0.007509f
C517 B.n477 VSUBS 0.007509f
C518 B.n478 VSUBS 0.007509f
C519 B.n479 VSUBS 0.007509f
C520 B.n480 VSUBS 0.007509f
C521 B.n481 VSUBS 0.007509f
C522 B.n482 VSUBS 0.007509f
C523 B.n483 VSUBS 0.007509f
C524 B.n484 VSUBS 0.007509f
C525 B.n485 VSUBS 0.007509f
C526 B.n486 VSUBS 0.007509f
C527 B.n487 VSUBS 0.007509f
C528 B.n488 VSUBS 0.007509f
C529 B.n489 VSUBS 0.007509f
C530 B.n490 VSUBS 0.007509f
C531 B.n491 VSUBS 0.007509f
C532 B.n492 VSUBS 0.007509f
C533 B.n493 VSUBS 0.007509f
C534 B.n494 VSUBS 0.007509f
C535 B.n495 VSUBS 0.007509f
C536 B.n496 VSUBS 0.007509f
C537 B.n497 VSUBS 0.007509f
C538 B.n498 VSUBS 0.007509f
C539 B.n499 VSUBS 0.007509f
C540 B.n500 VSUBS 0.007509f
C541 B.n501 VSUBS 0.007509f
C542 B.n502 VSUBS 0.007509f
C543 B.n503 VSUBS 0.007509f
C544 B.n504 VSUBS 0.007509f
C545 B.n505 VSUBS 0.007509f
C546 B.n506 VSUBS 0.007509f
C547 B.n507 VSUBS 0.007509f
C548 B.n508 VSUBS 0.007509f
C549 B.n509 VSUBS 0.007509f
C550 B.n510 VSUBS 0.007509f
C551 B.n511 VSUBS 0.007509f
C552 B.n512 VSUBS 0.007509f
C553 B.n513 VSUBS 0.007509f
C554 B.n514 VSUBS 0.007509f
C555 B.n515 VSUBS 0.007509f
C556 B.n516 VSUBS 0.007509f
C557 B.n517 VSUBS 0.007509f
C558 B.n518 VSUBS 0.007509f
C559 B.n519 VSUBS 0.007509f
C560 B.n520 VSUBS 0.007509f
C561 B.n521 VSUBS 0.007509f
C562 B.n522 VSUBS 0.007509f
C563 B.n523 VSUBS 0.007509f
C564 B.n524 VSUBS 0.007509f
C565 B.n525 VSUBS 0.007509f
C566 B.n526 VSUBS 0.007509f
C567 B.n527 VSUBS 0.007509f
C568 B.n528 VSUBS 0.007509f
C569 B.n529 VSUBS 0.007509f
C570 B.n530 VSUBS 0.007509f
C571 B.n531 VSUBS 0.007509f
C572 B.n532 VSUBS 0.007509f
C573 B.n533 VSUBS 0.007509f
C574 B.n534 VSUBS 0.007509f
C575 B.n535 VSUBS 0.007509f
C576 B.n536 VSUBS 0.007509f
C577 B.n537 VSUBS 0.007509f
C578 B.n538 VSUBS 0.007509f
C579 B.n539 VSUBS 0.007509f
C580 B.n540 VSUBS 0.007509f
C581 B.n541 VSUBS 0.007509f
C582 B.n542 VSUBS 0.007509f
C583 B.n543 VSUBS 0.007509f
C584 B.n544 VSUBS 0.007509f
C585 B.n545 VSUBS 0.007509f
C586 B.n546 VSUBS 0.007509f
C587 B.n547 VSUBS 0.007509f
C588 B.n548 VSUBS 0.007509f
C589 B.n549 VSUBS 0.007509f
C590 B.n550 VSUBS 0.007509f
C591 B.n551 VSUBS 0.007509f
C592 B.n552 VSUBS 0.007509f
C593 B.n553 VSUBS 0.007509f
C594 B.n554 VSUBS 0.007509f
C595 B.n555 VSUBS 0.007509f
C596 B.n556 VSUBS 0.007509f
C597 B.n557 VSUBS 0.007509f
C598 B.n558 VSUBS 0.007509f
C599 B.n559 VSUBS 0.007509f
C600 B.n560 VSUBS 0.007509f
C601 B.n561 VSUBS 0.007509f
C602 B.n562 VSUBS 0.007509f
C603 B.n563 VSUBS 0.007509f
C604 B.n564 VSUBS 0.007509f
C605 B.n565 VSUBS 0.007509f
C606 B.n566 VSUBS 0.007509f
C607 B.n567 VSUBS 0.007509f
C608 B.n568 VSUBS 0.007509f
C609 B.n569 VSUBS 0.007509f
C610 B.n570 VSUBS 0.007509f
C611 B.n571 VSUBS 0.007509f
C612 B.n572 VSUBS 0.007509f
C613 B.n573 VSUBS 0.007509f
C614 B.n574 VSUBS 0.007509f
C615 B.n575 VSUBS 0.007509f
C616 B.n576 VSUBS 0.007509f
C617 B.n577 VSUBS 0.007509f
C618 B.n578 VSUBS 0.007509f
C619 B.n579 VSUBS 0.007509f
C620 B.n580 VSUBS 0.007509f
C621 B.n581 VSUBS 0.007509f
C622 B.n582 VSUBS 0.007509f
C623 B.n583 VSUBS 0.007509f
C624 B.n584 VSUBS 0.007509f
C625 B.n585 VSUBS 0.007509f
C626 B.n586 VSUBS 0.007509f
C627 B.n587 VSUBS 0.007509f
C628 B.n588 VSUBS 0.007509f
C629 B.n589 VSUBS 0.007509f
C630 B.n590 VSUBS 0.007509f
C631 B.n591 VSUBS 0.007509f
C632 B.n592 VSUBS 0.007509f
C633 B.n593 VSUBS 0.007509f
C634 B.n594 VSUBS 0.007509f
C635 B.n595 VSUBS 0.007509f
C636 B.n596 VSUBS 0.007509f
C637 B.n597 VSUBS 0.007509f
C638 B.n598 VSUBS 0.007509f
C639 B.n599 VSUBS 0.007509f
C640 B.n600 VSUBS 0.007509f
C641 B.n601 VSUBS 0.007509f
C642 B.n602 VSUBS 0.007509f
C643 B.n603 VSUBS 0.007509f
C644 B.n604 VSUBS 0.007509f
C645 B.n605 VSUBS 0.007509f
C646 B.n606 VSUBS 0.007509f
C647 B.n607 VSUBS 0.007509f
C648 B.n608 VSUBS 0.007509f
C649 B.n609 VSUBS 0.007509f
C650 B.n610 VSUBS 0.007509f
C651 B.n611 VSUBS 0.007509f
C652 B.n612 VSUBS 0.007509f
C653 B.n613 VSUBS 0.007509f
C654 B.n614 VSUBS 0.007509f
C655 B.n615 VSUBS 0.007509f
C656 B.n616 VSUBS 0.007509f
C657 B.n617 VSUBS 0.007509f
C658 B.n618 VSUBS 0.007509f
C659 B.n619 VSUBS 0.007509f
C660 B.n620 VSUBS 0.007509f
C661 B.n621 VSUBS 0.007509f
C662 B.n622 VSUBS 0.007509f
C663 B.n623 VSUBS 0.007509f
C664 B.n624 VSUBS 0.007509f
C665 B.n625 VSUBS 0.007509f
C666 B.n626 VSUBS 0.007509f
C667 B.n627 VSUBS 0.007509f
C668 B.n628 VSUBS 0.007509f
C669 B.n629 VSUBS 0.007509f
C670 B.n630 VSUBS 0.007509f
C671 B.n631 VSUBS 0.007509f
C672 B.n632 VSUBS 0.007509f
C673 B.n633 VSUBS 0.007509f
C674 B.n634 VSUBS 0.007509f
C675 B.n635 VSUBS 0.007509f
C676 B.n636 VSUBS 0.007509f
C677 B.n637 VSUBS 0.007509f
C678 B.n638 VSUBS 0.017577f
C679 B.n639 VSUBS 0.016654f
C680 B.n640 VSUBS 0.017577f
C681 B.n641 VSUBS 0.007509f
C682 B.n642 VSUBS 0.007509f
C683 B.n643 VSUBS 0.007509f
C684 B.n644 VSUBS 0.007509f
C685 B.n645 VSUBS 0.007509f
C686 B.n646 VSUBS 0.007509f
C687 B.n647 VSUBS 0.007509f
C688 B.n648 VSUBS 0.007509f
C689 B.n649 VSUBS 0.007509f
C690 B.n650 VSUBS 0.007509f
C691 B.n651 VSUBS 0.007509f
C692 B.n652 VSUBS 0.007509f
C693 B.n653 VSUBS 0.007509f
C694 B.n654 VSUBS 0.007509f
C695 B.n655 VSUBS 0.007509f
C696 B.n656 VSUBS 0.007509f
C697 B.n657 VSUBS 0.007509f
C698 B.n658 VSUBS 0.007509f
C699 B.n659 VSUBS 0.007509f
C700 B.n660 VSUBS 0.007509f
C701 B.n661 VSUBS 0.007509f
C702 B.n662 VSUBS 0.007509f
C703 B.n663 VSUBS 0.007509f
C704 B.n664 VSUBS 0.007509f
C705 B.n665 VSUBS 0.007509f
C706 B.n666 VSUBS 0.007509f
C707 B.n667 VSUBS 0.007509f
C708 B.n668 VSUBS 0.007509f
C709 B.n669 VSUBS 0.007509f
C710 B.n670 VSUBS 0.007509f
C711 B.n671 VSUBS 0.007509f
C712 B.n672 VSUBS 0.007509f
C713 B.n673 VSUBS 0.007509f
C714 B.n674 VSUBS 0.007509f
C715 B.n675 VSUBS 0.007509f
C716 B.n676 VSUBS 0.007509f
C717 B.n677 VSUBS 0.007509f
C718 B.n678 VSUBS 0.007509f
C719 B.n679 VSUBS 0.007509f
C720 B.n680 VSUBS 0.007509f
C721 B.n681 VSUBS 0.007509f
C722 B.n682 VSUBS 0.007509f
C723 B.n683 VSUBS 0.007509f
C724 B.n684 VSUBS 0.007509f
C725 B.n685 VSUBS 0.007509f
C726 B.n686 VSUBS 0.007509f
C727 B.n687 VSUBS 0.007509f
C728 B.n688 VSUBS 0.007509f
C729 B.n689 VSUBS 0.007509f
C730 B.n690 VSUBS 0.007509f
C731 B.n691 VSUBS 0.007509f
C732 B.n692 VSUBS 0.007509f
C733 B.n693 VSUBS 0.007509f
C734 B.n694 VSUBS 0.007509f
C735 B.n695 VSUBS 0.007509f
C736 B.n696 VSUBS 0.007509f
C737 B.n697 VSUBS 0.00519f
C738 B.n698 VSUBS 0.017397f
C739 B.n699 VSUBS 0.006073f
C740 B.n700 VSUBS 0.007509f
C741 B.n701 VSUBS 0.007509f
C742 B.n702 VSUBS 0.007509f
C743 B.n703 VSUBS 0.007509f
C744 B.n704 VSUBS 0.007509f
C745 B.n705 VSUBS 0.007509f
C746 B.n706 VSUBS 0.007509f
C747 B.n707 VSUBS 0.007509f
C748 B.n708 VSUBS 0.007509f
C749 B.n709 VSUBS 0.007509f
C750 B.n710 VSUBS 0.007509f
C751 B.n711 VSUBS 0.006073f
C752 B.n712 VSUBS 0.017397f
C753 B.n713 VSUBS 0.00519f
C754 B.n714 VSUBS 0.007509f
C755 B.n715 VSUBS 0.007509f
C756 B.n716 VSUBS 0.007509f
C757 B.n717 VSUBS 0.007509f
C758 B.n718 VSUBS 0.007509f
C759 B.n719 VSUBS 0.007509f
C760 B.n720 VSUBS 0.007509f
C761 B.n721 VSUBS 0.007509f
C762 B.n722 VSUBS 0.007509f
C763 B.n723 VSUBS 0.007509f
C764 B.n724 VSUBS 0.007509f
C765 B.n725 VSUBS 0.007509f
C766 B.n726 VSUBS 0.007509f
C767 B.n727 VSUBS 0.007509f
C768 B.n728 VSUBS 0.007509f
C769 B.n729 VSUBS 0.007509f
C770 B.n730 VSUBS 0.007509f
C771 B.n731 VSUBS 0.007509f
C772 B.n732 VSUBS 0.007509f
C773 B.n733 VSUBS 0.007509f
C774 B.n734 VSUBS 0.007509f
C775 B.n735 VSUBS 0.007509f
C776 B.n736 VSUBS 0.007509f
C777 B.n737 VSUBS 0.007509f
C778 B.n738 VSUBS 0.007509f
C779 B.n739 VSUBS 0.007509f
C780 B.n740 VSUBS 0.007509f
C781 B.n741 VSUBS 0.007509f
C782 B.n742 VSUBS 0.007509f
C783 B.n743 VSUBS 0.007509f
C784 B.n744 VSUBS 0.007509f
C785 B.n745 VSUBS 0.007509f
C786 B.n746 VSUBS 0.007509f
C787 B.n747 VSUBS 0.007509f
C788 B.n748 VSUBS 0.007509f
C789 B.n749 VSUBS 0.007509f
C790 B.n750 VSUBS 0.007509f
C791 B.n751 VSUBS 0.007509f
C792 B.n752 VSUBS 0.007509f
C793 B.n753 VSUBS 0.007509f
C794 B.n754 VSUBS 0.007509f
C795 B.n755 VSUBS 0.007509f
C796 B.n756 VSUBS 0.007509f
C797 B.n757 VSUBS 0.007509f
C798 B.n758 VSUBS 0.007509f
C799 B.n759 VSUBS 0.007509f
C800 B.n760 VSUBS 0.007509f
C801 B.n761 VSUBS 0.007509f
C802 B.n762 VSUBS 0.007509f
C803 B.n763 VSUBS 0.007509f
C804 B.n764 VSUBS 0.007509f
C805 B.n765 VSUBS 0.007509f
C806 B.n766 VSUBS 0.007509f
C807 B.n767 VSUBS 0.007509f
C808 B.n768 VSUBS 0.007509f
C809 B.n769 VSUBS 0.007509f
C810 B.n770 VSUBS 0.017577f
C811 B.n771 VSUBS 0.017577f
C812 B.n772 VSUBS 0.016654f
C813 B.n773 VSUBS 0.007509f
C814 B.n774 VSUBS 0.007509f
C815 B.n775 VSUBS 0.007509f
C816 B.n776 VSUBS 0.007509f
C817 B.n777 VSUBS 0.007509f
C818 B.n778 VSUBS 0.007509f
C819 B.n779 VSUBS 0.007509f
C820 B.n780 VSUBS 0.007509f
C821 B.n781 VSUBS 0.007509f
C822 B.n782 VSUBS 0.007509f
C823 B.n783 VSUBS 0.007509f
C824 B.n784 VSUBS 0.007509f
C825 B.n785 VSUBS 0.007509f
C826 B.n786 VSUBS 0.007509f
C827 B.n787 VSUBS 0.007509f
C828 B.n788 VSUBS 0.007509f
C829 B.n789 VSUBS 0.007509f
C830 B.n790 VSUBS 0.007509f
C831 B.n791 VSUBS 0.007509f
C832 B.n792 VSUBS 0.007509f
C833 B.n793 VSUBS 0.007509f
C834 B.n794 VSUBS 0.007509f
C835 B.n795 VSUBS 0.007509f
C836 B.n796 VSUBS 0.007509f
C837 B.n797 VSUBS 0.007509f
C838 B.n798 VSUBS 0.007509f
C839 B.n799 VSUBS 0.007509f
C840 B.n800 VSUBS 0.007509f
C841 B.n801 VSUBS 0.007509f
C842 B.n802 VSUBS 0.007509f
C843 B.n803 VSUBS 0.007509f
C844 B.n804 VSUBS 0.007509f
C845 B.n805 VSUBS 0.007509f
C846 B.n806 VSUBS 0.007509f
C847 B.n807 VSUBS 0.007509f
C848 B.n808 VSUBS 0.007509f
C849 B.n809 VSUBS 0.007509f
C850 B.n810 VSUBS 0.007509f
C851 B.n811 VSUBS 0.007509f
C852 B.n812 VSUBS 0.007509f
C853 B.n813 VSUBS 0.007509f
C854 B.n814 VSUBS 0.007509f
C855 B.n815 VSUBS 0.007509f
C856 B.n816 VSUBS 0.007509f
C857 B.n817 VSUBS 0.007509f
C858 B.n818 VSUBS 0.007509f
C859 B.n819 VSUBS 0.007509f
C860 B.n820 VSUBS 0.007509f
C861 B.n821 VSUBS 0.007509f
C862 B.n822 VSUBS 0.007509f
C863 B.n823 VSUBS 0.007509f
C864 B.n824 VSUBS 0.007509f
C865 B.n825 VSUBS 0.007509f
C866 B.n826 VSUBS 0.007509f
C867 B.n827 VSUBS 0.007509f
C868 B.n828 VSUBS 0.007509f
C869 B.n829 VSUBS 0.007509f
C870 B.n830 VSUBS 0.007509f
C871 B.n831 VSUBS 0.007509f
C872 B.n832 VSUBS 0.007509f
C873 B.n833 VSUBS 0.007509f
C874 B.n834 VSUBS 0.007509f
C875 B.n835 VSUBS 0.007509f
C876 B.n836 VSUBS 0.007509f
C877 B.n837 VSUBS 0.007509f
C878 B.n838 VSUBS 0.007509f
C879 B.n839 VSUBS 0.007509f
C880 B.n840 VSUBS 0.007509f
C881 B.n841 VSUBS 0.007509f
C882 B.n842 VSUBS 0.007509f
C883 B.n843 VSUBS 0.007509f
C884 B.n844 VSUBS 0.007509f
C885 B.n845 VSUBS 0.007509f
C886 B.n846 VSUBS 0.007509f
C887 B.n847 VSUBS 0.007509f
C888 B.n848 VSUBS 0.007509f
C889 B.n849 VSUBS 0.007509f
C890 B.n850 VSUBS 0.007509f
C891 B.n851 VSUBS 0.007509f
C892 B.n852 VSUBS 0.007509f
C893 B.n853 VSUBS 0.007509f
C894 B.n854 VSUBS 0.007509f
C895 B.n855 VSUBS 0.007509f
C896 B.n856 VSUBS 0.007509f
C897 B.n857 VSUBS 0.007509f
C898 B.n858 VSUBS 0.007509f
C899 B.n859 VSUBS 0.007509f
C900 B.n860 VSUBS 0.007509f
C901 B.n861 VSUBS 0.007509f
C902 B.n862 VSUBS 0.007509f
C903 B.n863 VSUBS 0.007509f
C904 B.n864 VSUBS 0.007509f
C905 B.n865 VSUBS 0.007509f
C906 B.n866 VSUBS 0.007509f
C907 B.n867 VSUBS 0.017002f
C908 VDD2.t1 VSUBS 0.265891f
C909 VDD2.t6 VSUBS 0.265891f
C910 VDD2.n0 VSUBS 2.06032f
C911 VDD2.t0 VSUBS 0.265891f
C912 VDD2.t4 VSUBS 0.265891f
C913 VDD2.n1 VSUBS 2.06032f
C914 VDD2.n2 VSUBS 5.12994f
C915 VDD2.t7 VSUBS 0.265891f
C916 VDD2.t2 VSUBS 0.265891f
C917 VDD2.n3 VSUBS 2.0388f
C918 VDD2.n4 VSUBS 4.17598f
C919 VDD2.t5 VSUBS 0.265891f
C920 VDD2.t3 VSUBS 0.265891f
C921 VDD2.n5 VSUBS 2.06026f
C922 VN.t3 VSUBS 2.64802f
C923 VN.n0 VSUBS 1.04358f
C924 VN.n1 VSUBS 0.026078f
C925 VN.n2 VSUBS 0.021216f
C926 VN.n3 VSUBS 0.026078f
C927 VN.t7 VSUBS 2.64802f
C928 VN.n4 VSUBS 0.934275f
C929 VN.n5 VSUBS 0.026078f
C930 VN.n6 VSUBS 0.03807f
C931 VN.n7 VSUBS 0.026078f
C932 VN.n8 VSUBS 0.030126f
C933 VN.t1 VSUBS 2.64802f
C934 VN.n9 VSUBS 1.01685f
C935 VN.t6 VSUBS 2.98381f
C936 VN.n10 VSUBS 0.967502f
C937 VN.n11 VSUBS 0.308509f
C938 VN.n12 VSUBS 0.026078f
C939 VN.n13 VSUBS 0.048603f
C940 VN.n14 VSUBS 0.048603f
C941 VN.n15 VSUBS 0.03807f
C942 VN.n16 VSUBS 0.026078f
C943 VN.n17 VSUBS 0.026078f
C944 VN.n18 VSUBS 0.026078f
C945 VN.n19 VSUBS 0.048603f
C946 VN.n20 VSUBS 0.048603f
C947 VN.n21 VSUBS 0.030126f
C948 VN.n22 VSUBS 0.026078f
C949 VN.n23 VSUBS 0.026078f
C950 VN.n24 VSUBS 0.043083f
C951 VN.n25 VSUBS 0.048603f
C952 VN.n26 VSUBS 0.051243f
C953 VN.n27 VSUBS 0.026078f
C954 VN.n28 VSUBS 0.026078f
C955 VN.n29 VSUBS 0.026078f
C956 VN.n30 VSUBS 0.052283f
C957 VN.n31 VSUBS 0.048603f
C958 VN.n32 VSUBS 0.041164f
C959 VN.n33 VSUBS 0.04209f
C960 VN.n34 VSUBS 0.061667f
C961 VN.t0 VSUBS 2.64802f
C962 VN.n35 VSUBS 1.04358f
C963 VN.n36 VSUBS 0.026078f
C964 VN.n37 VSUBS 0.021216f
C965 VN.n38 VSUBS 0.026078f
C966 VN.t5 VSUBS 2.64802f
C967 VN.n39 VSUBS 0.934275f
C968 VN.n40 VSUBS 0.026078f
C969 VN.n41 VSUBS 0.03807f
C970 VN.n42 VSUBS 0.026078f
C971 VN.n43 VSUBS 0.030126f
C972 VN.t4 VSUBS 2.98381f
C973 VN.t2 VSUBS 2.64802f
C974 VN.n44 VSUBS 1.01685f
C975 VN.n45 VSUBS 0.967502f
C976 VN.n46 VSUBS 0.308509f
C977 VN.n47 VSUBS 0.026078f
C978 VN.n48 VSUBS 0.048603f
C979 VN.n49 VSUBS 0.048603f
C980 VN.n50 VSUBS 0.03807f
C981 VN.n51 VSUBS 0.026078f
C982 VN.n52 VSUBS 0.026078f
C983 VN.n53 VSUBS 0.026078f
C984 VN.n54 VSUBS 0.048603f
C985 VN.n55 VSUBS 0.048603f
C986 VN.n56 VSUBS 0.030126f
C987 VN.n57 VSUBS 0.026078f
C988 VN.n58 VSUBS 0.026078f
C989 VN.n59 VSUBS 0.043083f
C990 VN.n60 VSUBS 0.048603f
C991 VN.n61 VSUBS 0.051243f
C992 VN.n62 VSUBS 0.026078f
C993 VN.n63 VSUBS 0.026078f
C994 VN.n64 VSUBS 0.026078f
C995 VN.n65 VSUBS 0.052283f
C996 VN.n66 VSUBS 0.048603f
C997 VN.n67 VSUBS 0.041164f
C998 VN.n68 VSUBS 0.04209f
C999 VN.n69 VSUBS 1.66669f
C1000 VTAIL.t3 VSUBS 0.228331f
C1001 VTAIL.t4 VSUBS 0.228331f
C1002 VTAIL.n0 VSUBS 1.61086f
C1003 VTAIL.n1 VSUBS 0.870244f
C1004 VTAIL.t2 VSUBS 2.13573f
C1005 VTAIL.n2 VSUBS 1.00297f
C1006 VTAIL.t11 VSUBS 2.13573f
C1007 VTAIL.n3 VSUBS 1.00297f
C1008 VTAIL.t10 VSUBS 0.228331f
C1009 VTAIL.t15 VSUBS 0.228331f
C1010 VTAIL.n4 VSUBS 1.61086f
C1011 VTAIL.n5 VSUBS 1.13772f
C1012 VTAIL.t8 VSUBS 2.13573f
C1013 VTAIL.n6 VSUBS 2.39533f
C1014 VTAIL.t0 VSUBS 2.13574f
C1015 VTAIL.n7 VSUBS 2.39531f
C1016 VTAIL.t6 VSUBS 0.228331f
C1017 VTAIL.t1 VSUBS 0.228331f
C1018 VTAIL.n8 VSUBS 1.61087f
C1019 VTAIL.n9 VSUBS 1.13772f
C1020 VTAIL.t7 VSUBS 2.13574f
C1021 VTAIL.n10 VSUBS 1.00295f
C1022 VTAIL.t9 VSUBS 2.13574f
C1023 VTAIL.n11 VSUBS 1.00295f
C1024 VTAIL.t12 VSUBS 0.228331f
C1025 VTAIL.t13 VSUBS 0.228331f
C1026 VTAIL.n12 VSUBS 1.61087f
C1027 VTAIL.n13 VSUBS 1.13772f
C1028 VTAIL.t14 VSUBS 2.13573f
C1029 VTAIL.n14 VSUBS 2.39533f
C1030 VTAIL.t5 VSUBS 2.13573f
C1031 VTAIL.n15 VSUBS 2.3904f
C1032 VDD1.t2 VSUBS 0.268245f
C1033 VDD1.t5 VSUBS 0.268245f
C1034 VDD1.n0 VSUBS 2.08035f
C1035 VDD1.t3 VSUBS 0.268245f
C1036 VDD1.t7 VSUBS 0.268245f
C1037 VDD1.n1 VSUBS 2.07856f
C1038 VDD1.t4 VSUBS 0.268245f
C1039 VDD1.t0 VSUBS 0.268245f
C1040 VDD1.n2 VSUBS 2.07856f
C1041 VDD1.n3 VSUBS 5.23921f
C1042 VDD1.t1 VSUBS 0.268245f
C1043 VDD1.t6 VSUBS 0.268245f
C1044 VDD1.n4 VSUBS 2.05684f
C1045 VDD1.n5 VSUBS 4.2516f
C1046 VP.t4 VSUBS 2.90248f
C1047 VP.n0 VSUBS 1.14386f
C1048 VP.n1 VSUBS 0.028584f
C1049 VP.n2 VSUBS 0.023255f
C1050 VP.n3 VSUBS 0.028584f
C1051 VP.t0 VSUBS 2.90248f
C1052 VP.n4 VSUBS 1.02405f
C1053 VP.n5 VSUBS 0.028584f
C1054 VP.n6 VSUBS 0.041728f
C1055 VP.n7 VSUBS 0.028584f
C1056 VP.n8 VSUBS 0.03302f
C1057 VP.n9 VSUBS 0.028584f
C1058 VP.n10 VSUBS 0.023255f
C1059 VP.n11 VSUBS 0.028584f
C1060 VP.t7 VSUBS 2.90248f
C1061 VP.n12 VSUBS 1.14386f
C1062 VP.t1 VSUBS 2.90248f
C1063 VP.n13 VSUBS 1.14386f
C1064 VP.n14 VSUBS 0.028584f
C1065 VP.n15 VSUBS 0.023255f
C1066 VP.n16 VSUBS 0.028584f
C1067 VP.t2 VSUBS 2.90248f
C1068 VP.n17 VSUBS 1.02405f
C1069 VP.n18 VSUBS 0.028584f
C1070 VP.n19 VSUBS 0.041728f
C1071 VP.n20 VSUBS 0.028584f
C1072 VP.n21 VSUBS 0.03302f
C1073 VP.t6 VSUBS 3.27054f
C1074 VP.t3 VSUBS 2.90248f
C1075 VP.n22 VSUBS 1.11456f
C1076 VP.n23 VSUBS 1.06047f
C1077 VP.n24 VSUBS 0.338156f
C1078 VP.n25 VSUBS 0.028584f
C1079 VP.n26 VSUBS 0.053274f
C1080 VP.n27 VSUBS 0.053274f
C1081 VP.n28 VSUBS 0.041728f
C1082 VP.n29 VSUBS 0.028584f
C1083 VP.n30 VSUBS 0.028584f
C1084 VP.n31 VSUBS 0.028584f
C1085 VP.n32 VSUBS 0.053274f
C1086 VP.n33 VSUBS 0.053274f
C1087 VP.n34 VSUBS 0.03302f
C1088 VP.n35 VSUBS 0.028584f
C1089 VP.n36 VSUBS 0.028584f
C1090 VP.n37 VSUBS 0.047223f
C1091 VP.n38 VSUBS 0.053274f
C1092 VP.n39 VSUBS 0.056167f
C1093 VP.n40 VSUBS 0.028584f
C1094 VP.n41 VSUBS 0.028584f
C1095 VP.n42 VSUBS 0.028584f
C1096 VP.n43 VSUBS 0.057307f
C1097 VP.n44 VSUBS 0.053274f
C1098 VP.n45 VSUBS 0.045119f
C1099 VP.n46 VSUBS 0.046134f
C1100 VP.n47 VSUBS 1.81547f
C1101 VP.n48 VSUBS 1.83448f
C1102 VP.n49 VSUBS 0.046134f
C1103 VP.n50 VSUBS 0.045119f
C1104 VP.n51 VSUBS 0.053274f
C1105 VP.n52 VSUBS 0.057307f
C1106 VP.n53 VSUBS 0.028584f
C1107 VP.n54 VSUBS 0.028584f
C1108 VP.n55 VSUBS 0.028584f
C1109 VP.n56 VSUBS 0.056167f
C1110 VP.n57 VSUBS 0.053274f
C1111 VP.t5 VSUBS 2.90248f
C1112 VP.n58 VSUBS 1.02405f
C1113 VP.n59 VSUBS 0.047223f
C1114 VP.n60 VSUBS 0.028584f
C1115 VP.n61 VSUBS 0.028584f
C1116 VP.n62 VSUBS 0.028584f
C1117 VP.n63 VSUBS 0.053274f
C1118 VP.n64 VSUBS 0.053274f
C1119 VP.n65 VSUBS 0.041728f
C1120 VP.n66 VSUBS 0.028584f
C1121 VP.n67 VSUBS 0.028584f
C1122 VP.n68 VSUBS 0.028584f
C1123 VP.n69 VSUBS 0.053274f
C1124 VP.n70 VSUBS 0.053274f
C1125 VP.n71 VSUBS 0.03302f
C1126 VP.n72 VSUBS 0.028584f
C1127 VP.n73 VSUBS 0.028584f
C1128 VP.n74 VSUBS 0.047223f
C1129 VP.n75 VSUBS 0.053274f
C1130 VP.n76 VSUBS 0.056167f
C1131 VP.n77 VSUBS 0.028584f
C1132 VP.n78 VSUBS 0.028584f
C1133 VP.n79 VSUBS 0.028584f
C1134 VP.n80 VSUBS 0.057307f
C1135 VP.n81 VSUBS 0.053274f
C1136 VP.n82 VSUBS 0.045119f
C1137 VP.n83 VSUBS 0.046134f
C1138 VP.n84 VSUBS 0.067592f
.ends

