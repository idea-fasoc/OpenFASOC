* NGSPICE file created from diff_pair_sample_0429.ext - technology: sky130A

.subckt diff_pair_sample_0429 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=2.08395 pd=12.96 as=4.9257 ps=26.04 w=12.63 l=1.09
X1 VTAIL.t8 VP.t1 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.08395 pd=12.96 as=2.08395 ps=12.96 w=12.63 l=1.09
X2 VDD1.t3 VP.t2 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=4.9257 pd=26.04 as=2.08395 ps=12.96 w=12.63 l=1.09
X3 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=4.9257 pd=26.04 as=0 ps=0 w=12.63 l=1.09
X4 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=4.9257 pd=26.04 as=0 ps=0 w=12.63 l=1.09
X5 VDD2.t5 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.9257 pd=26.04 as=2.08395 ps=12.96 w=12.63 l=1.09
X6 VTAIL.t0 VN.t1 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.08395 pd=12.96 as=2.08395 ps=12.96 w=12.63 l=1.09
X7 VDD2.t3 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.08395 pd=12.96 as=4.9257 ps=26.04 w=12.63 l=1.09
X8 VTAIL.t10 VP.t3 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.08395 pd=12.96 as=2.08395 ps=12.96 w=12.63 l=1.09
X9 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.9257 pd=26.04 as=0 ps=0 w=12.63 l=1.09
X10 VDD2.t2 VN.t3 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=4.9257 pd=26.04 as=2.08395 ps=12.96 w=12.63 l=1.09
X11 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.9257 pd=26.04 as=0 ps=0 w=12.63 l=1.09
X12 VDD2.t1 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.08395 pd=12.96 as=4.9257 ps=26.04 w=12.63 l=1.09
X13 VDD1.t1 VP.t4 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=2.08395 pd=12.96 as=4.9257 ps=26.04 w=12.63 l=1.09
X14 VDD1.t0 VP.t5 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=4.9257 pd=26.04 as=2.08395 ps=12.96 w=12.63 l=1.09
X15 VTAIL.t3 VN.t5 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=2.08395 pd=12.96 as=2.08395 ps=12.96 w=12.63 l=1.09
R0 VP.n3 VP.t2 338.505
R1 VP.n8 VP.t5 315.512
R2 VP.n14 VP.t0 315.512
R3 VP.n6 VP.t4 315.512
R4 VP.n12 VP.t1 279.25
R5 VP.n4 VP.t3 279.25
R6 VP.n5 VP.n2 161.3
R7 VP.n13 VP.n0 161.3
R8 VP.n12 VP.n11 161.3
R9 VP.n10 VP.n1 161.3
R10 VP.n7 VP.n6 80.6037
R11 VP.n15 VP.n14 80.6037
R12 VP.n9 VP.n8 80.6037
R13 VP.n8 VP.n1 50.4025
R14 VP.n14 VP.n13 50.4025
R15 VP.n6 VP.n5 50.4025
R16 VP.n9 VP.n7 43.4105
R17 VP.n4 VP.n3 32.6271
R18 VP.n3 VP.n2 28.1515
R19 VP.n12 VP.n1 24.4675
R20 VP.n13 VP.n12 24.4675
R21 VP.n5 VP.n4 24.4675
R22 VP.n7 VP.n2 0.285035
R23 VP.n10 VP.n9 0.285035
R24 VP.n15 VP.n0 0.285035
R25 VP.n11 VP.n10 0.189894
R26 VP.n11 VP.n0 0.189894
R27 VP VP.n15 0.146778
R28 VTAIL.n286 VTAIL.n285 289.615
R29 VTAIL.n70 VTAIL.n69 289.615
R30 VTAIL.n216 VTAIL.n215 289.615
R31 VTAIL.n144 VTAIL.n143 289.615
R32 VTAIL.n240 VTAIL.n239 185
R33 VTAIL.n245 VTAIL.n244 185
R34 VTAIL.n247 VTAIL.n246 185
R35 VTAIL.n236 VTAIL.n235 185
R36 VTAIL.n253 VTAIL.n252 185
R37 VTAIL.n255 VTAIL.n254 185
R38 VTAIL.n232 VTAIL.n231 185
R39 VTAIL.n261 VTAIL.n260 185
R40 VTAIL.n263 VTAIL.n262 185
R41 VTAIL.n228 VTAIL.n227 185
R42 VTAIL.n269 VTAIL.n268 185
R43 VTAIL.n271 VTAIL.n270 185
R44 VTAIL.n224 VTAIL.n223 185
R45 VTAIL.n277 VTAIL.n276 185
R46 VTAIL.n279 VTAIL.n278 185
R47 VTAIL.n220 VTAIL.n219 185
R48 VTAIL.n285 VTAIL.n284 185
R49 VTAIL.n24 VTAIL.n23 185
R50 VTAIL.n29 VTAIL.n28 185
R51 VTAIL.n31 VTAIL.n30 185
R52 VTAIL.n20 VTAIL.n19 185
R53 VTAIL.n37 VTAIL.n36 185
R54 VTAIL.n39 VTAIL.n38 185
R55 VTAIL.n16 VTAIL.n15 185
R56 VTAIL.n45 VTAIL.n44 185
R57 VTAIL.n47 VTAIL.n46 185
R58 VTAIL.n12 VTAIL.n11 185
R59 VTAIL.n53 VTAIL.n52 185
R60 VTAIL.n55 VTAIL.n54 185
R61 VTAIL.n8 VTAIL.n7 185
R62 VTAIL.n61 VTAIL.n60 185
R63 VTAIL.n63 VTAIL.n62 185
R64 VTAIL.n4 VTAIL.n3 185
R65 VTAIL.n69 VTAIL.n68 185
R66 VTAIL.n215 VTAIL.n214 185
R67 VTAIL.n150 VTAIL.n149 185
R68 VTAIL.n209 VTAIL.n208 185
R69 VTAIL.n207 VTAIL.n206 185
R70 VTAIL.n154 VTAIL.n153 185
R71 VTAIL.n201 VTAIL.n200 185
R72 VTAIL.n199 VTAIL.n198 185
R73 VTAIL.n158 VTAIL.n157 185
R74 VTAIL.n193 VTAIL.n192 185
R75 VTAIL.n191 VTAIL.n190 185
R76 VTAIL.n162 VTAIL.n161 185
R77 VTAIL.n185 VTAIL.n184 185
R78 VTAIL.n183 VTAIL.n182 185
R79 VTAIL.n166 VTAIL.n165 185
R80 VTAIL.n177 VTAIL.n176 185
R81 VTAIL.n175 VTAIL.n174 185
R82 VTAIL.n170 VTAIL.n169 185
R83 VTAIL.n143 VTAIL.n142 185
R84 VTAIL.n78 VTAIL.n77 185
R85 VTAIL.n137 VTAIL.n136 185
R86 VTAIL.n135 VTAIL.n134 185
R87 VTAIL.n82 VTAIL.n81 185
R88 VTAIL.n129 VTAIL.n128 185
R89 VTAIL.n127 VTAIL.n126 185
R90 VTAIL.n86 VTAIL.n85 185
R91 VTAIL.n121 VTAIL.n120 185
R92 VTAIL.n119 VTAIL.n118 185
R93 VTAIL.n90 VTAIL.n89 185
R94 VTAIL.n113 VTAIL.n112 185
R95 VTAIL.n111 VTAIL.n110 185
R96 VTAIL.n94 VTAIL.n93 185
R97 VTAIL.n105 VTAIL.n104 185
R98 VTAIL.n103 VTAIL.n102 185
R99 VTAIL.n98 VTAIL.n97 185
R100 VTAIL.n241 VTAIL.t2 147.659
R101 VTAIL.n25 VTAIL.t9 147.659
R102 VTAIL.n171 VTAIL.t7 147.659
R103 VTAIL.n99 VTAIL.t4 147.659
R104 VTAIL.n245 VTAIL.n239 104.615
R105 VTAIL.n246 VTAIL.n245 104.615
R106 VTAIL.n246 VTAIL.n235 104.615
R107 VTAIL.n253 VTAIL.n235 104.615
R108 VTAIL.n254 VTAIL.n253 104.615
R109 VTAIL.n254 VTAIL.n231 104.615
R110 VTAIL.n261 VTAIL.n231 104.615
R111 VTAIL.n262 VTAIL.n261 104.615
R112 VTAIL.n262 VTAIL.n227 104.615
R113 VTAIL.n269 VTAIL.n227 104.615
R114 VTAIL.n270 VTAIL.n269 104.615
R115 VTAIL.n270 VTAIL.n223 104.615
R116 VTAIL.n277 VTAIL.n223 104.615
R117 VTAIL.n278 VTAIL.n277 104.615
R118 VTAIL.n278 VTAIL.n219 104.615
R119 VTAIL.n285 VTAIL.n219 104.615
R120 VTAIL.n29 VTAIL.n23 104.615
R121 VTAIL.n30 VTAIL.n29 104.615
R122 VTAIL.n30 VTAIL.n19 104.615
R123 VTAIL.n37 VTAIL.n19 104.615
R124 VTAIL.n38 VTAIL.n37 104.615
R125 VTAIL.n38 VTAIL.n15 104.615
R126 VTAIL.n45 VTAIL.n15 104.615
R127 VTAIL.n46 VTAIL.n45 104.615
R128 VTAIL.n46 VTAIL.n11 104.615
R129 VTAIL.n53 VTAIL.n11 104.615
R130 VTAIL.n54 VTAIL.n53 104.615
R131 VTAIL.n54 VTAIL.n7 104.615
R132 VTAIL.n61 VTAIL.n7 104.615
R133 VTAIL.n62 VTAIL.n61 104.615
R134 VTAIL.n62 VTAIL.n3 104.615
R135 VTAIL.n69 VTAIL.n3 104.615
R136 VTAIL.n215 VTAIL.n149 104.615
R137 VTAIL.n208 VTAIL.n149 104.615
R138 VTAIL.n208 VTAIL.n207 104.615
R139 VTAIL.n207 VTAIL.n153 104.615
R140 VTAIL.n200 VTAIL.n153 104.615
R141 VTAIL.n200 VTAIL.n199 104.615
R142 VTAIL.n199 VTAIL.n157 104.615
R143 VTAIL.n192 VTAIL.n157 104.615
R144 VTAIL.n192 VTAIL.n191 104.615
R145 VTAIL.n191 VTAIL.n161 104.615
R146 VTAIL.n184 VTAIL.n161 104.615
R147 VTAIL.n184 VTAIL.n183 104.615
R148 VTAIL.n183 VTAIL.n165 104.615
R149 VTAIL.n176 VTAIL.n165 104.615
R150 VTAIL.n176 VTAIL.n175 104.615
R151 VTAIL.n175 VTAIL.n169 104.615
R152 VTAIL.n143 VTAIL.n77 104.615
R153 VTAIL.n136 VTAIL.n77 104.615
R154 VTAIL.n136 VTAIL.n135 104.615
R155 VTAIL.n135 VTAIL.n81 104.615
R156 VTAIL.n128 VTAIL.n81 104.615
R157 VTAIL.n128 VTAIL.n127 104.615
R158 VTAIL.n127 VTAIL.n85 104.615
R159 VTAIL.n120 VTAIL.n85 104.615
R160 VTAIL.n120 VTAIL.n119 104.615
R161 VTAIL.n119 VTAIL.n89 104.615
R162 VTAIL.n112 VTAIL.n89 104.615
R163 VTAIL.n112 VTAIL.n111 104.615
R164 VTAIL.n111 VTAIL.n93 104.615
R165 VTAIL.n104 VTAIL.n93 104.615
R166 VTAIL.n104 VTAIL.n103 104.615
R167 VTAIL.n103 VTAIL.n97 104.615
R168 VTAIL.t2 VTAIL.n239 52.3082
R169 VTAIL.t9 VTAIL.n23 52.3082
R170 VTAIL.t7 VTAIL.n169 52.3082
R171 VTAIL.t4 VTAIL.n97 52.3082
R172 VTAIL.n147 VTAIL.n146 47.4387
R173 VTAIL.n75 VTAIL.n74 47.4387
R174 VTAIL.n1 VTAIL.n0 47.4377
R175 VTAIL.n73 VTAIL.n72 47.4377
R176 VTAIL.n287 VTAIL.n286 34.7066
R177 VTAIL.n71 VTAIL.n70 34.7066
R178 VTAIL.n217 VTAIL.n216 34.7066
R179 VTAIL.n145 VTAIL.n144 34.7066
R180 VTAIL.n75 VTAIL.n73 25.7031
R181 VTAIL.n287 VTAIL.n217 24.4789
R182 VTAIL.n241 VTAIL.n240 15.6677
R183 VTAIL.n25 VTAIL.n24 15.6677
R184 VTAIL.n171 VTAIL.n170 15.6677
R185 VTAIL.n99 VTAIL.n98 15.6677
R186 VTAIL.n244 VTAIL.n243 12.8005
R187 VTAIL.n284 VTAIL.n218 12.8005
R188 VTAIL.n28 VTAIL.n27 12.8005
R189 VTAIL.n68 VTAIL.n2 12.8005
R190 VTAIL.n214 VTAIL.n148 12.8005
R191 VTAIL.n174 VTAIL.n173 12.8005
R192 VTAIL.n142 VTAIL.n76 12.8005
R193 VTAIL.n102 VTAIL.n101 12.8005
R194 VTAIL.n247 VTAIL.n238 12.0247
R195 VTAIL.n283 VTAIL.n220 12.0247
R196 VTAIL.n31 VTAIL.n22 12.0247
R197 VTAIL.n67 VTAIL.n4 12.0247
R198 VTAIL.n213 VTAIL.n150 12.0247
R199 VTAIL.n177 VTAIL.n168 12.0247
R200 VTAIL.n141 VTAIL.n78 12.0247
R201 VTAIL.n105 VTAIL.n96 12.0247
R202 VTAIL.n248 VTAIL.n236 11.249
R203 VTAIL.n280 VTAIL.n279 11.249
R204 VTAIL.n32 VTAIL.n20 11.249
R205 VTAIL.n64 VTAIL.n63 11.249
R206 VTAIL.n210 VTAIL.n209 11.249
R207 VTAIL.n178 VTAIL.n166 11.249
R208 VTAIL.n138 VTAIL.n137 11.249
R209 VTAIL.n106 VTAIL.n94 11.249
R210 VTAIL.n252 VTAIL.n251 10.4732
R211 VTAIL.n276 VTAIL.n222 10.4732
R212 VTAIL.n36 VTAIL.n35 10.4732
R213 VTAIL.n60 VTAIL.n6 10.4732
R214 VTAIL.n206 VTAIL.n152 10.4732
R215 VTAIL.n182 VTAIL.n181 10.4732
R216 VTAIL.n134 VTAIL.n80 10.4732
R217 VTAIL.n110 VTAIL.n109 10.4732
R218 VTAIL.n255 VTAIL.n234 9.69747
R219 VTAIL.n275 VTAIL.n224 9.69747
R220 VTAIL.n39 VTAIL.n18 9.69747
R221 VTAIL.n59 VTAIL.n8 9.69747
R222 VTAIL.n205 VTAIL.n154 9.69747
R223 VTAIL.n185 VTAIL.n164 9.69747
R224 VTAIL.n133 VTAIL.n82 9.69747
R225 VTAIL.n113 VTAIL.n92 9.69747
R226 VTAIL.n282 VTAIL.n218 9.45567
R227 VTAIL.n66 VTAIL.n2 9.45567
R228 VTAIL.n212 VTAIL.n148 9.45567
R229 VTAIL.n140 VTAIL.n76 9.45567
R230 VTAIL.n265 VTAIL.n264 9.3005
R231 VTAIL.n267 VTAIL.n266 9.3005
R232 VTAIL.n226 VTAIL.n225 9.3005
R233 VTAIL.n273 VTAIL.n272 9.3005
R234 VTAIL.n275 VTAIL.n274 9.3005
R235 VTAIL.n222 VTAIL.n221 9.3005
R236 VTAIL.n281 VTAIL.n280 9.3005
R237 VTAIL.n283 VTAIL.n282 9.3005
R238 VTAIL.n259 VTAIL.n258 9.3005
R239 VTAIL.n257 VTAIL.n256 9.3005
R240 VTAIL.n234 VTAIL.n233 9.3005
R241 VTAIL.n251 VTAIL.n250 9.3005
R242 VTAIL.n249 VTAIL.n248 9.3005
R243 VTAIL.n238 VTAIL.n237 9.3005
R244 VTAIL.n243 VTAIL.n242 9.3005
R245 VTAIL.n230 VTAIL.n229 9.3005
R246 VTAIL.n49 VTAIL.n48 9.3005
R247 VTAIL.n51 VTAIL.n50 9.3005
R248 VTAIL.n10 VTAIL.n9 9.3005
R249 VTAIL.n57 VTAIL.n56 9.3005
R250 VTAIL.n59 VTAIL.n58 9.3005
R251 VTAIL.n6 VTAIL.n5 9.3005
R252 VTAIL.n65 VTAIL.n64 9.3005
R253 VTAIL.n67 VTAIL.n66 9.3005
R254 VTAIL.n43 VTAIL.n42 9.3005
R255 VTAIL.n41 VTAIL.n40 9.3005
R256 VTAIL.n18 VTAIL.n17 9.3005
R257 VTAIL.n35 VTAIL.n34 9.3005
R258 VTAIL.n33 VTAIL.n32 9.3005
R259 VTAIL.n22 VTAIL.n21 9.3005
R260 VTAIL.n27 VTAIL.n26 9.3005
R261 VTAIL.n14 VTAIL.n13 9.3005
R262 VTAIL.n213 VTAIL.n212 9.3005
R263 VTAIL.n211 VTAIL.n210 9.3005
R264 VTAIL.n152 VTAIL.n151 9.3005
R265 VTAIL.n205 VTAIL.n204 9.3005
R266 VTAIL.n203 VTAIL.n202 9.3005
R267 VTAIL.n156 VTAIL.n155 9.3005
R268 VTAIL.n197 VTAIL.n196 9.3005
R269 VTAIL.n195 VTAIL.n194 9.3005
R270 VTAIL.n160 VTAIL.n159 9.3005
R271 VTAIL.n189 VTAIL.n188 9.3005
R272 VTAIL.n187 VTAIL.n186 9.3005
R273 VTAIL.n164 VTAIL.n163 9.3005
R274 VTAIL.n181 VTAIL.n180 9.3005
R275 VTAIL.n179 VTAIL.n178 9.3005
R276 VTAIL.n168 VTAIL.n167 9.3005
R277 VTAIL.n173 VTAIL.n172 9.3005
R278 VTAIL.n125 VTAIL.n124 9.3005
R279 VTAIL.n84 VTAIL.n83 9.3005
R280 VTAIL.n131 VTAIL.n130 9.3005
R281 VTAIL.n133 VTAIL.n132 9.3005
R282 VTAIL.n80 VTAIL.n79 9.3005
R283 VTAIL.n139 VTAIL.n138 9.3005
R284 VTAIL.n141 VTAIL.n140 9.3005
R285 VTAIL.n123 VTAIL.n122 9.3005
R286 VTAIL.n88 VTAIL.n87 9.3005
R287 VTAIL.n117 VTAIL.n116 9.3005
R288 VTAIL.n115 VTAIL.n114 9.3005
R289 VTAIL.n92 VTAIL.n91 9.3005
R290 VTAIL.n109 VTAIL.n108 9.3005
R291 VTAIL.n107 VTAIL.n106 9.3005
R292 VTAIL.n96 VTAIL.n95 9.3005
R293 VTAIL.n101 VTAIL.n100 9.3005
R294 VTAIL.n256 VTAIL.n232 8.92171
R295 VTAIL.n272 VTAIL.n271 8.92171
R296 VTAIL.n40 VTAIL.n16 8.92171
R297 VTAIL.n56 VTAIL.n55 8.92171
R298 VTAIL.n202 VTAIL.n201 8.92171
R299 VTAIL.n186 VTAIL.n162 8.92171
R300 VTAIL.n130 VTAIL.n129 8.92171
R301 VTAIL.n114 VTAIL.n90 8.92171
R302 VTAIL.n260 VTAIL.n259 8.14595
R303 VTAIL.n268 VTAIL.n226 8.14595
R304 VTAIL.n44 VTAIL.n43 8.14595
R305 VTAIL.n52 VTAIL.n10 8.14595
R306 VTAIL.n198 VTAIL.n156 8.14595
R307 VTAIL.n190 VTAIL.n189 8.14595
R308 VTAIL.n126 VTAIL.n84 8.14595
R309 VTAIL.n118 VTAIL.n117 8.14595
R310 VTAIL.n263 VTAIL.n230 7.3702
R311 VTAIL.n267 VTAIL.n228 7.3702
R312 VTAIL.n47 VTAIL.n14 7.3702
R313 VTAIL.n51 VTAIL.n12 7.3702
R314 VTAIL.n197 VTAIL.n158 7.3702
R315 VTAIL.n193 VTAIL.n160 7.3702
R316 VTAIL.n125 VTAIL.n86 7.3702
R317 VTAIL.n121 VTAIL.n88 7.3702
R318 VTAIL.n264 VTAIL.n263 6.59444
R319 VTAIL.n264 VTAIL.n228 6.59444
R320 VTAIL.n48 VTAIL.n47 6.59444
R321 VTAIL.n48 VTAIL.n12 6.59444
R322 VTAIL.n194 VTAIL.n158 6.59444
R323 VTAIL.n194 VTAIL.n193 6.59444
R324 VTAIL.n122 VTAIL.n86 6.59444
R325 VTAIL.n122 VTAIL.n121 6.59444
R326 VTAIL.n260 VTAIL.n230 5.81868
R327 VTAIL.n268 VTAIL.n267 5.81868
R328 VTAIL.n44 VTAIL.n14 5.81868
R329 VTAIL.n52 VTAIL.n51 5.81868
R330 VTAIL.n198 VTAIL.n197 5.81868
R331 VTAIL.n190 VTAIL.n160 5.81868
R332 VTAIL.n126 VTAIL.n125 5.81868
R333 VTAIL.n118 VTAIL.n88 5.81868
R334 VTAIL.n259 VTAIL.n232 5.04292
R335 VTAIL.n271 VTAIL.n226 5.04292
R336 VTAIL.n43 VTAIL.n16 5.04292
R337 VTAIL.n55 VTAIL.n10 5.04292
R338 VTAIL.n201 VTAIL.n156 5.04292
R339 VTAIL.n189 VTAIL.n162 5.04292
R340 VTAIL.n129 VTAIL.n84 5.04292
R341 VTAIL.n117 VTAIL.n90 5.04292
R342 VTAIL.n242 VTAIL.n241 4.38563
R343 VTAIL.n26 VTAIL.n25 4.38563
R344 VTAIL.n172 VTAIL.n171 4.38563
R345 VTAIL.n100 VTAIL.n99 4.38563
R346 VTAIL.n256 VTAIL.n255 4.26717
R347 VTAIL.n272 VTAIL.n224 4.26717
R348 VTAIL.n40 VTAIL.n39 4.26717
R349 VTAIL.n56 VTAIL.n8 4.26717
R350 VTAIL.n202 VTAIL.n154 4.26717
R351 VTAIL.n186 VTAIL.n185 4.26717
R352 VTAIL.n130 VTAIL.n82 4.26717
R353 VTAIL.n114 VTAIL.n113 4.26717
R354 VTAIL.n252 VTAIL.n234 3.49141
R355 VTAIL.n276 VTAIL.n275 3.49141
R356 VTAIL.n36 VTAIL.n18 3.49141
R357 VTAIL.n60 VTAIL.n59 3.49141
R358 VTAIL.n206 VTAIL.n205 3.49141
R359 VTAIL.n182 VTAIL.n164 3.49141
R360 VTAIL.n134 VTAIL.n133 3.49141
R361 VTAIL.n110 VTAIL.n92 3.49141
R362 VTAIL.n251 VTAIL.n236 2.71565
R363 VTAIL.n279 VTAIL.n222 2.71565
R364 VTAIL.n35 VTAIL.n20 2.71565
R365 VTAIL.n63 VTAIL.n6 2.71565
R366 VTAIL.n209 VTAIL.n152 2.71565
R367 VTAIL.n181 VTAIL.n166 2.71565
R368 VTAIL.n137 VTAIL.n80 2.71565
R369 VTAIL.n109 VTAIL.n94 2.71565
R370 VTAIL.n248 VTAIL.n247 1.93989
R371 VTAIL.n280 VTAIL.n220 1.93989
R372 VTAIL.n32 VTAIL.n31 1.93989
R373 VTAIL.n64 VTAIL.n4 1.93989
R374 VTAIL.n210 VTAIL.n150 1.93989
R375 VTAIL.n178 VTAIL.n177 1.93989
R376 VTAIL.n138 VTAIL.n78 1.93989
R377 VTAIL.n106 VTAIL.n105 1.93989
R378 VTAIL.n0 VTAIL.t11 1.5682
R379 VTAIL.n0 VTAIL.t0 1.5682
R380 VTAIL.n72 VTAIL.t5 1.5682
R381 VTAIL.n72 VTAIL.t8 1.5682
R382 VTAIL.n146 VTAIL.t6 1.5682
R383 VTAIL.n146 VTAIL.t10 1.5682
R384 VTAIL.n74 VTAIL.t1 1.5682
R385 VTAIL.n74 VTAIL.t3 1.5682
R386 VTAIL.n145 VTAIL.n75 1.22464
R387 VTAIL.n217 VTAIL.n147 1.22464
R388 VTAIL.n73 VTAIL.n71 1.22464
R389 VTAIL.n244 VTAIL.n238 1.16414
R390 VTAIL.n284 VTAIL.n283 1.16414
R391 VTAIL.n28 VTAIL.n22 1.16414
R392 VTAIL.n68 VTAIL.n67 1.16414
R393 VTAIL.n214 VTAIL.n213 1.16414
R394 VTAIL.n174 VTAIL.n168 1.16414
R395 VTAIL.n142 VTAIL.n141 1.16414
R396 VTAIL.n102 VTAIL.n96 1.16414
R397 VTAIL.n147 VTAIL.n145 1.0824
R398 VTAIL.n71 VTAIL.n1 1.0824
R399 VTAIL VTAIL.n287 0.860414
R400 VTAIL.n243 VTAIL.n240 0.388379
R401 VTAIL.n286 VTAIL.n218 0.388379
R402 VTAIL.n27 VTAIL.n24 0.388379
R403 VTAIL.n70 VTAIL.n2 0.388379
R404 VTAIL.n216 VTAIL.n148 0.388379
R405 VTAIL.n173 VTAIL.n170 0.388379
R406 VTAIL.n144 VTAIL.n76 0.388379
R407 VTAIL.n101 VTAIL.n98 0.388379
R408 VTAIL VTAIL.n1 0.364724
R409 VTAIL.n242 VTAIL.n237 0.155672
R410 VTAIL.n249 VTAIL.n237 0.155672
R411 VTAIL.n250 VTAIL.n249 0.155672
R412 VTAIL.n250 VTAIL.n233 0.155672
R413 VTAIL.n257 VTAIL.n233 0.155672
R414 VTAIL.n258 VTAIL.n257 0.155672
R415 VTAIL.n258 VTAIL.n229 0.155672
R416 VTAIL.n265 VTAIL.n229 0.155672
R417 VTAIL.n266 VTAIL.n265 0.155672
R418 VTAIL.n266 VTAIL.n225 0.155672
R419 VTAIL.n273 VTAIL.n225 0.155672
R420 VTAIL.n274 VTAIL.n273 0.155672
R421 VTAIL.n274 VTAIL.n221 0.155672
R422 VTAIL.n281 VTAIL.n221 0.155672
R423 VTAIL.n282 VTAIL.n281 0.155672
R424 VTAIL.n26 VTAIL.n21 0.155672
R425 VTAIL.n33 VTAIL.n21 0.155672
R426 VTAIL.n34 VTAIL.n33 0.155672
R427 VTAIL.n34 VTAIL.n17 0.155672
R428 VTAIL.n41 VTAIL.n17 0.155672
R429 VTAIL.n42 VTAIL.n41 0.155672
R430 VTAIL.n42 VTAIL.n13 0.155672
R431 VTAIL.n49 VTAIL.n13 0.155672
R432 VTAIL.n50 VTAIL.n49 0.155672
R433 VTAIL.n50 VTAIL.n9 0.155672
R434 VTAIL.n57 VTAIL.n9 0.155672
R435 VTAIL.n58 VTAIL.n57 0.155672
R436 VTAIL.n58 VTAIL.n5 0.155672
R437 VTAIL.n65 VTAIL.n5 0.155672
R438 VTAIL.n66 VTAIL.n65 0.155672
R439 VTAIL.n212 VTAIL.n211 0.155672
R440 VTAIL.n211 VTAIL.n151 0.155672
R441 VTAIL.n204 VTAIL.n151 0.155672
R442 VTAIL.n204 VTAIL.n203 0.155672
R443 VTAIL.n203 VTAIL.n155 0.155672
R444 VTAIL.n196 VTAIL.n155 0.155672
R445 VTAIL.n196 VTAIL.n195 0.155672
R446 VTAIL.n195 VTAIL.n159 0.155672
R447 VTAIL.n188 VTAIL.n159 0.155672
R448 VTAIL.n188 VTAIL.n187 0.155672
R449 VTAIL.n187 VTAIL.n163 0.155672
R450 VTAIL.n180 VTAIL.n163 0.155672
R451 VTAIL.n180 VTAIL.n179 0.155672
R452 VTAIL.n179 VTAIL.n167 0.155672
R453 VTAIL.n172 VTAIL.n167 0.155672
R454 VTAIL.n140 VTAIL.n139 0.155672
R455 VTAIL.n139 VTAIL.n79 0.155672
R456 VTAIL.n132 VTAIL.n79 0.155672
R457 VTAIL.n132 VTAIL.n131 0.155672
R458 VTAIL.n131 VTAIL.n83 0.155672
R459 VTAIL.n124 VTAIL.n83 0.155672
R460 VTAIL.n124 VTAIL.n123 0.155672
R461 VTAIL.n123 VTAIL.n87 0.155672
R462 VTAIL.n116 VTAIL.n87 0.155672
R463 VTAIL.n116 VTAIL.n115 0.155672
R464 VTAIL.n115 VTAIL.n91 0.155672
R465 VTAIL.n108 VTAIL.n91 0.155672
R466 VTAIL.n108 VTAIL.n107 0.155672
R467 VTAIL.n107 VTAIL.n95 0.155672
R468 VTAIL.n100 VTAIL.n95 0.155672
R469 VDD1.n68 VDD1.n67 289.615
R470 VDD1.n137 VDD1.n136 289.615
R471 VDD1.n67 VDD1.n66 185
R472 VDD1.n2 VDD1.n1 185
R473 VDD1.n61 VDD1.n60 185
R474 VDD1.n59 VDD1.n58 185
R475 VDD1.n6 VDD1.n5 185
R476 VDD1.n53 VDD1.n52 185
R477 VDD1.n51 VDD1.n50 185
R478 VDD1.n10 VDD1.n9 185
R479 VDD1.n45 VDD1.n44 185
R480 VDD1.n43 VDD1.n42 185
R481 VDD1.n14 VDD1.n13 185
R482 VDD1.n37 VDD1.n36 185
R483 VDD1.n35 VDD1.n34 185
R484 VDD1.n18 VDD1.n17 185
R485 VDD1.n29 VDD1.n28 185
R486 VDD1.n27 VDD1.n26 185
R487 VDD1.n22 VDD1.n21 185
R488 VDD1.n91 VDD1.n90 185
R489 VDD1.n96 VDD1.n95 185
R490 VDD1.n98 VDD1.n97 185
R491 VDD1.n87 VDD1.n86 185
R492 VDD1.n104 VDD1.n103 185
R493 VDD1.n106 VDD1.n105 185
R494 VDD1.n83 VDD1.n82 185
R495 VDD1.n112 VDD1.n111 185
R496 VDD1.n114 VDD1.n113 185
R497 VDD1.n79 VDD1.n78 185
R498 VDD1.n120 VDD1.n119 185
R499 VDD1.n122 VDD1.n121 185
R500 VDD1.n75 VDD1.n74 185
R501 VDD1.n128 VDD1.n127 185
R502 VDD1.n130 VDD1.n129 185
R503 VDD1.n71 VDD1.n70 185
R504 VDD1.n136 VDD1.n135 185
R505 VDD1.n92 VDD1.t0 147.659
R506 VDD1.n23 VDD1.t3 147.659
R507 VDD1.n67 VDD1.n1 104.615
R508 VDD1.n60 VDD1.n1 104.615
R509 VDD1.n60 VDD1.n59 104.615
R510 VDD1.n59 VDD1.n5 104.615
R511 VDD1.n52 VDD1.n5 104.615
R512 VDD1.n52 VDD1.n51 104.615
R513 VDD1.n51 VDD1.n9 104.615
R514 VDD1.n44 VDD1.n9 104.615
R515 VDD1.n44 VDD1.n43 104.615
R516 VDD1.n43 VDD1.n13 104.615
R517 VDD1.n36 VDD1.n13 104.615
R518 VDD1.n36 VDD1.n35 104.615
R519 VDD1.n35 VDD1.n17 104.615
R520 VDD1.n28 VDD1.n17 104.615
R521 VDD1.n28 VDD1.n27 104.615
R522 VDD1.n27 VDD1.n21 104.615
R523 VDD1.n96 VDD1.n90 104.615
R524 VDD1.n97 VDD1.n96 104.615
R525 VDD1.n97 VDD1.n86 104.615
R526 VDD1.n104 VDD1.n86 104.615
R527 VDD1.n105 VDD1.n104 104.615
R528 VDD1.n105 VDD1.n82 104.615
R529 VDD1.n112 VDD1.n82 104.615
R530 VDD1.n113 VDD1.n112 104.615
R531 VDD1.n113 VDD1.n78 104.615
R532 VDD1.n120 VDD1.n78 104.615
R533 VDD1.n121 VDD1.n120 104.615
R534 VDD1.n121 VDD1.n74 104.615
R535 VDD1.n128 VDD1.n74 104.615
R536 VDD1.n129 VDD1.n128 104.615
R537 VDD1.n129 VDD1.n70 104.615
R538 VDD1.n136 VDD1.n70 104.615
R539 VDD1.n139 VDD1.n138 64.3672
R540 VDD1.n141 VDD1.n140 64.1165
R541 VDD1 VDD1.n68 52.3616
R542 VDD1.t3 VDD1.n21 52.3082
R543 VDD1.t0 VDD1.n90 52.3082
R544 VDD1.n139 VDD1.n137 52.2481
R545 VDD1.n141 VDD1.n139 39.7768
R546 VDD1.n23 VDD1.n22 15.6677
R547 VDD1.n92 VDD1.n91 15.6677
R548 VDD1.n66 VDD1.n0 12.8005
R549 VDD1.n26 VDD1.n25 12.8005
R550 VDD1.n95 VDD1.n94 12.8005
R551 VDD1.n135 VDD1.n69 12.8005
R552 VDD1.n65 VDD1.n2 12.0247
R553 VDD1.n29 VDD1.n20 12.0247
R554 VDD1.n98 VDD1.n89 12.0247
R555 VDD1.n134 VDD1.n71 12.0247
R556 VDD1.n62 VDD1.n61 11.249
R557 VDD1.n30 VDD1.n18 11.249
R558 VDD1.n99 VDD1.n87 11.249
R559 VDD1.n131 VDD1.n130 11.249
R560 VDD1.n58 VDD1.n4 10.4732
R561 VDD1.n34 VDD1.n33 10.4732
R562 VDD1.n103 VDD1.n102 10.4732
R563 VDD1.n127 VDD1.n73 10.4732
R564 VDD1.n57 VDD1.n6 9.69747
R565 VDD1.n37 VDD1.n16 9.69747
R566 VDD1.n106 VDD1.n85 9.69747
R567 VDD1.n126 VDD1.n75 9.69747
R568 VDD1.n64 VDD1.n0 9.45567
R569 VDD1.n133 VDD1.n69 9.45567
R570 VDD1.n49 VDD1.n48 9.3005
R571 VDD1.n8 VDD1.n7 9.3005
R572 VDD1.n55 VDD1.n54 9.3005
R573 VDD1.n57 VDD1.n56 9.3005
R574 VDD1.n4 VDD1.n3 9.3005
R575 VDD1.n63 VDD1.n62 9.3005
R576 VDD1.n65 VDD1.n64 9.3005
R577 VDD1.n47 VDD1.n46 9.3005
R578 VDD1.n12 VDD1.n11 9.3005
R579 VDD1.n41 VDD1.n40 9.3005
R580 VDD1.n39 VDD1.n38 9.3005
R581 VDD1.n16 VDD1.n15 9.3005
R582 VDD1.n33 VDD1.n32 9.3005
R583 VDD1.n31 VDD1.n30 9.3005
R584 VDD1.n20 VDD1.n19 9.3005
R585 VDD1.n25 VDD1.n24 9.3005
R586 VDD1.n116 VDD1.n115 9.3005
R587 VDD1.n118 VDD1.n117 9.3005
R588 VDD1.n77 VDD1.n76 9.3005
R589 VDD1.n124 VDD1.n123 9.3005
R590 VDD1.n126 VDD1.n125 9.3005
R591 VDD1.n73 VDD1.n72 9.3005
R592 VDD1.n132 VDD1.n131 9.3005
R593 VDD1.n134 VDD1.n133 9.3005
R594 VDD1.n110 VDD1.n109 9.3005
R595 VDD1.n108 VDD1.n107 9.3005
R596 VDD1.n85 VDD1.n84 9.3005
R597 VDD1.n102 VDD1.n101 9.3005
R598 VDD1.n100 VDD1.n99 9.3005
R599 VDD1.n89 VDD1.n88 9.3005
R600 VDD1.n94 VDD1.n93 9.3005
R601 VDD1.n81 VDD1.n80 9.3005
R602 VDD1.n54 VDD1.n53 8.92171
R603 VDD1.n38 VDD1.n14 8.92171
R604 VDD1.n107 VDD1.n83 8.92171
R605 VDD1.n123 VDD1.n122 8.92171
R606 VDD1.n50 VDD1.n8 8.14595
R607 VDD1.n42 VDD1.n41 8.14595
R608 VDD1.n111 VDD1.n110 8.14595
R609 VDD1.n119 VDD1.n77 8.14595
R610 VDD1.n49 VDD1.n10 7.3702
R611 VDD1.n45 VDD1.n12 7.3702
R612 VDD1.n114 VDD1.n81 7.3702
R613 VDD1.n118 VDD1.n79 7.3702
R614 VDD1.n46 VDD1.n10 6.59444
R615 VDD1.n46 VDD1.n45 6.59444
R616 VDD1.n115 VDD1.n114 6.59444
R617 VDD1.n115 VDD1.n79 6.59444
R618 VDD1.n50 VDD1.n49 5.81868
R619 VDD1.n42 VDD1.n12 5.81868
R620 VDD1.n111 VDD1.n81 5.81868
R621 VDD1.n119 VDD1.n118 5.81868
R622 VDD1.n53 VDD1.n8 5.04292
R623 VDD1.n41 VDD1.n14 5.04292
R624 VDD1.n110 VDD1.n83 5.04292
R625 VDD1.n122 VDD1.n77 5.04292
R626 VDD1.n93 VDD1.n92 4.38563
R627 VDD1.n24 VDD1.n23 4.38563
R628 VDD1.n54 VDD1.n6 4.26717
R629 VDD1.n38 VDD1.n37 4.26717
R630 VDD1.n107 VDD1.n106 4.26717
R631 VDD1.n123 VDD1.n75 4.26717
R632 VDD1.n58 VDD1.n57 3.49141
R633 VDD1.n34 VDD1.n16 3.49141
R634 VDD1.n103 VDD1.n85 3.49141
R635 VDD1.n127 VDD1.n126 3.49141
R636 VDD1.n61 VDD1.n4 2.71565
R637 VDD1.n33 VDD1.n18 2.71565
R638 VDD1.n102 VDD1.n87 2.71565
R639 VDD1.n130 VDD1.n73 2.71565
R640 VDD1.n62 VDD1.n2 1.93989
R641 VDD1.n30 VDD1.n29 1.93989
R642 VDD1.n99 VDD1.n98 1.93989
R643 VDD1.n131 VDD1.n71 1.93989
R644 VDD1.n140 VDD1.t2 1.5682
R645 VDD1.n140 VDD1.t1 1.5682
R646 VDD1.n138 VDD1.t4 1.5682
R647 VDD1.n138 VDD1.t5 1.5682
R648 VDD1.n66 VDD1.n65 1.16414
R649 VDD1.n26 VDD1.n20 1.16414
R650 VDD1.n95 VDD1.n89 1.16414
R651 VDD1.n135 VDD1.n134 1.16414
R652 VDD1.n68 VDD1.n0 0.388379
R653 VDD1.n25 VDD1.n22 0.388379
R654 VDD1.n94 VDD1.n91 0.388379
R655 VDD1.n137 VDD1.n69 0.388379
R656 VDD1 VDD1.n141 0.248345
R657 VDD1.n64 VDD1.n63 0.155672
R658 VDD1.n63 VDD1.n3 0.155672
R659 VDD1.n56 VDD1.n3 0.155672
R660 VDD1.n56 VDD1.n55 0.155672
R661 VDD1.n55 VDD1.n7 0.155672
R662 VDD1.n48 VDD1.n7 0.155672
R663 VDD1.n48 VDD1.n47 0.155672
R664 VDD1.n47 VDD1.n11 0.155672
R665 VDD1.n40 VDD1.n11 0.155672
R666 VDD1.n40 VDD1.n39 0.155672
R667 VDD1.n39 VDD1.n15 0.155672
R668 VDD1.n32 VDD1.n15 0.155672
R669 VDD1.n32 VDD1.n31 0.155672
R670 VDD1.n31 VDD1.n19 0.155672
R671 VDD1.n24 VDD1.n19 0.155672
R672 VDD1.n93 VDD1.n88 0.155672
R673 VDD1.n100 VDD1.n88 0.155672
R674 VDD1.n101 VDD1.n100 0.155672
R675 VDD1.n101 VDD1.n84 0.155672
R676 VDD1.n108 VDD1.n84 0.155672
R677 VDD1.n109 VDD1.n108 0.155672
R678 VDD1.n109 VDD1.n80 0.155672
R679 VDD1.n116 VDD1.n80 0.155672
R680 VDD1.n117 VDD1.n116 0.155672
R681 VDD1.n117 VDD1.n76 0.155672
R682 VDD1.n124 VDD1.n76 0.155672
R683 VDD1.n125 VDD1.n124 0.155672
R684 VDD1.n125 VDD1.n72 0.155672
R685 VDD1.n132 VDD1.n72 0.155672
R686 VDD1.n133 VDD1.n132 0.155672
R687 B.n699 B.n698 585
R688 B.n700 B.n699 585
R689 B.n294 B.n97 585
R690 B.n293 B.n292 585
R691 B.n291 B.n290 585
R692 B.n289 B.n288 585
R693 B.n287 B.n286 585
R694 B.n285 B.n284 585
R695 B.n283 B.n282 585
R696 B.n281 B.n280 585
R697 B.n279 B.n278 585
R698 B.n277 B.n276 585
R699 B.n275 B.n274 585
R700 B.n273 B.n272 585
R701 B.n271 B.n270 585
R702 B.n269 B.n268 585
R703 B.n267 B.n266 585
R704 B.n265 B.n264 585
R705 B.n263 B.n262 585
R706 B.n261 B.n260 585
R707 B.n259 B.n258 585
R708 B.n257 B.n256 585
R709 B.n255 B.n254 585
R710 B.n253 B.n252 585
R711 B.n251 B.n250 585
R712 B.n249 B.n248 585
R713 B.n247 B.n246 585
R714 B.n245 B.n244 585
R715 B.n243 B.n242 585
R716 B.n241 B.n240 585
R717 B.n239 B.n238 585
R718 B.n237 B.n236 585
R719 B.n235 B.n234 585
R720 B.n233 B.n232 585
R721 B.n231 B.n230 585
R722 B.n229 B.n228 585
R723 B.n227 B.n226 585
R724 B.n225 B.n224 585
R725 B.n223 B.n222 585
R726 B.n221 B.n220 585
R727 B.n219 B.n218 585
R728 B.n217 B.n216 585
R729 B.n215 B.n214 585
R730 B.n213 B.n212 585
R731 B.n211 B.n210 585
R732 B.n208 B.n207 585
R733 B.n206 B.n205 585
R734 B.n204 B.n203 585
R735 B.n202 B.n201 585
R736 B.n200 B.n199 585
R737 B.n198 B.n197 585
R738 B.n196 B.n195 585
R739 B.n194 B.n193 585
R740 B.n192 B.n191 585
R741 B.n190 B.n189 585
R742 B.n188 B.n187 585
R743 B.n186 B.n185 585
R744 B.n184 B.n183 585
R745 B.n182 B.n181 585
R746 B.n180 B.n179 585
R747 B.n178 B.n177 585
R748 B.n176 B.n175 585
R749 B.n174 B.n173 585
R750 B.n172 B.n171 585
R751 B.n170 B.n169 585
R752 B.n168 B.n167 585
R753 B.n166 B.n165 585
R754 B.n164 B.n163 585
R755 B.n162 B.n161 585
R756 B.n160 B.n159 585
R757 B.n158 B.n157 585
R758 B.n156 B.n155 585
R759 B.n154 B.n153 585
R760 B.n152 B.n151 585
R761 B.n150 B.n149 585
R762 B.n148 B.n147 585
R763 B.n146 B.n145 585
R764 B.n144 B.n143 585
R765 B.n142 B.n141 585
R766 B.n140 B.n139 585
R767 B.n138 B.n137 585
R768 B.n136 B.n135 585
R769 B.n134 B.n133 585
R770 B.n132 B.n131 585
R771 B.n130 B.n129 585
R772 B.n128 B.n127 585
R773 B.n126 B.n125 585
R774 B.n124 B.n123 585
R775 B.n122 B.n121 585
R776 B.n120 B.n119 585
R777 B.n118 B.n117 585
R778 B.n116 B.n115 585
R779 B.n114 B.n113 585
R780 B.n112 B.n111 585
R781 B.n110 B.n109 585
R782 B.n108 B.n107 585
R783 B.n106 B.n105 585
R784 B.n104 B.n103 585
R785 B.n697 B.n48 585
R786 B.n701 B.n48 585
R787 B.n696 B.n47 585
R788 B.n702 B.n47 585
R789 B.n695 B.n694 585
R790 B.n694 B.n43 585
R791 B.n693 B.n42 585
R792 B.n708 B.n42 585
R793 B.n692 B.n41 585
R794 B.n709 B.n41 585
R795 B.n691 B.n40 585
R796 B.n710 B.n40 585
R797 B.n690 B.n689 585
R798 B.n689 B.n36 585
R799 B.n688 B.n35 585
R800 B.n716 B.n35 585
R801 B.n687 B.n34 585
R802 B.n717 B.n34 585
R803 B.n686 B.n33 585
R804 B.n718 B.n33 585
R805 B.n685 B.n684 585
R806 B.n684 B.n29 585
R807 B.n683 B.n28 585
R808 B.n724 B.n28 585
R809 B.n682 B.n27 585
R810 B.n725 B.n27 585
R811 B.n681 B.n26 585
R812 B.n726 B.n26 585
R813 B.n680 B.n679 585
R814 B.n679 B.n22 585
R815 B.n678 B.n21 585
R816 B.n732 B.n21 585
R817 B.n677 B.n20 585
R818 B.n733 B.n20 585
R819 B.n676 B.n19 585
R820 B.n734 B.n19 585
R821 B.n675 B.n674 585
R822 B.n674 B.n15 585
R823 B.n673 B.n14 585
R824 B.n740 B.n14 585
R825 B.n672 B.n13 585
R826 B.n741 B.n13 585
R827 B.n671 B.n12 585
R828 B.n742 B.n12 585
R829 B.n670 B.n669 585
R830 B.n669 B.n8 585
R831 B.n668 B.n7 585
R832 B.n748 B.n7 585
R833 B.n667 B.n6 585
R834 B.n749 B.n6 585
R835 B.n666 B.n5 585
R836 B.n750 B.n5 585
R837 B.n665 B.n664 585
R838 B.n664 B.n4 585
R839 B.n663 B.n295 585
R840 B.n663 B.n662 585
R841 B.n653 B.n296 585
R842 B.n297 B.n296 585
R843 B.n655 B.n654 585
R844 B.n656 B.n655 585
R845 B.n652 B.n302 585
R846 B.n302 B.n301 585
R847 B.n651 B.n650 585
R848 B.n650 B.n649 585
R849 B.n304 B.n303 585
R850 B.n305 B.n304 585
R851 B.n642 B.n641 585
R852 B.n643 B.n642 585
R853 B.n640 B.n310 585
R854 B.n310 B.n309 585
R855 B.n639 B.n638 585
R856 B.n638 B.n637 585
R857 B.n312 B.n311 585
R858 B.n313 B.n312 585
R859 B.n630 B.n629 585
R860 B.n631 B.n630 585
R861 B.n628 B.n317 585
R862 B.n321 B.n317 585
R863 B.n627 B.n626 585
R864 B.n626 B.n625 585
R865 B.n319 B.n318 585
R866 B.n320 B.n319 585
R867 B.n618 B.n617 585
R868 B.n619 B.n618 585
R869 B.n616 B.n326 585
R870 B.n326 B.n325 585
R871 B.n615 B.n614 585
R872 B.n614 B.n613 585
R873 B.n328 B.n327 585
R874 B.n329 B.n328 585
R875 B.n606 B.n605 585
R876 B.n607 B.n606 585
R877 B.n604 B.n334 585
R878 B.n334 B.n333 585
R879 B.n603 B.n602 585
R880 B.n602 B.n601 585
R881 B.n336 B.n335 585
R882 B.n337 B.n336 585
R883 B.n594 B.n593 585
R884 B.n595 B.n594 585
R885 B.n592 B.n342 585
R886 B.n342 B.n341 585
R887 B.n586 B.n585 585
R888 B.n584 B.n392 585
R889 B.n583 B.n391 585
R890 B.n588 B.n391 585
R891 B.n582 B.n581 585
R892 B.n580 B.n579 585
R893 B.n578 B.n577 585
R894 B.n576 B.n575 585
R895 B.n574 B.n573 585
R896 B.n572 B.n571 585
R897 B.n570 B.n569 585
R898 B.n568 B.n567 585
R899 B.n566 B.n565 585
R900 B.n564 B.n563 585
R901 B.n562 B.n561 585
R902 B.n560 B.n559 585
R903 B.n558 B.n557 585
R904 B.n556 B.n555 585
R905 B.n554 B.n553 585
R906 B.n552 B.n551 585
R907 B.n550 B.n549 585
R908 B.n548 B.n547 585
R909 B.n546 B.n545 585
R910 B.n544 B.n543 585
R911 B.n542 B.n541 585
R912 B.n540 B.n539 585
R913 B.n538 B.n537 585
R914 B.n536 B.n535 585
R915 B.n534 B.n533 585
R916 B.n532 B.n531 585
R917 B.n530 B.n529 585
R918 B.n528 B.n527 585
R919 B.n526 B.n525 585
R920 B.n524 B.n523 585
R921 B.n522 B.n521 585
R922 B.n520 B.n519 585
R923 B.n518 B.n517 585
R924 B.n516 B.n515 585
R925 B.n514 B.n513 585
R926 B.n512 B.n511 585
R927 B.n510 B.n509 585
R928 B.n508 B.n507 585
R929 B.n506 B.n505 585
R930 B.n504 B.n503 585
R931 B.n502 B.n501 585
R932 B.n499 B.n498 585
R933 B.n497 B.n496 585
R934 B.n495 B.n494 585
R935 B.n493 B.n492 585
R936 B.n491 B.n490 585
R937 B.n489 B.n488 585
R938 B.n487 B.n486 585
R939 B.n485 B.n484 585
R940 B.n483 B.n482 585
R941 B.n481 B.n480 585
R942 B.n479 B.n478 585
R943 B.n477 B.n476 585
R944 B.n475 B.n474 585
R945 B.n473 B.n472 585
R946 B.n471 B.n470 585
R947 B.n469 B.n468 585
R948 B.n467 B.n466 585
R949 B.n465 B.n464 585
R950 B.n463 B.n462 585
R951 B.n461 B.n460 585
R952 B.n459 B.n458 585
R953 B.n457 B.n456 585
R954 B.n455 B.n454 585
R955 B.n453 B.n452 585
R956 B.n451 B.n450 585
R957 B.n449 B.n448 585
R958 B.n447 B.n446 585
R959 B.n445 B.n444 585
R960 B.n443 B.n442 585
R961 B.n441 B.n440 585
R962 B.n439 B.n438 585
R963 B.n437 B.n436 585
R964 B.n435 B.n434 585
R965 B.n433 B.n432 585
R966 B.n431 B.n430 585
R967 B.n429 B.n428 585
R968 B.n427 B.n426 585
R969 B.n425 B.n424 585
R970 B.n423 B.n422 585
R971 B.n421 B.n420 585
R972 B.n419 B.n418 585
R973 B.n417 B.n416 585
R974 B.n415 B.n414 585
R975 B.n413 B.n412 585
R976 B.n411 B.n410 585
R977 B.n409 B.n408 585
R978 B.n407 B.n406 585
R979 B.n405 B.n404 585
R980 B.n403 B.n402 585
R981 B.n401 B.n400 585
R982 B.n399 B.n398 585
R983 B.n344 B.n343 585
R984 B.n591 B.n590 585
R985 B.n340 B.n339 585
R986 B.n341 B.n340 585
R987 B.n597 B.n596 585
R988 B.n596 B.n595 585
R989 B.n598 B.n338 585
R990 B.n338 B.n337 585
R991 B.n600 B.n599 585
R992 B.n601 B.n600 585
R993 B.n332 B.n331 585
R994 B.n333 B.n332 585
R995 B.n609 B.n608 585
R996 B.n608 B.n607 585
R997 B.n610 B.n330 585
R998 B.n330 B.n329 585
R999 B.n612 B.n611 585
R1000 B.n613 B.n612 585
R1001 B.n324 B.n323 585
R1002 B.n325 B.n324 585
R1003 B.n621 B.n620 585
R1004 B.n620 B.n619 585
R1005 B.n622 B.n322 585
R1006 B.n322 B.n320 585
R1007 B.n624 B.n623 585
R1008 B.n625 B.n624 585
R1009 B.n316 B.n315 585
R1010 B.n321 B.n316 585
R1011 B.n633 B.n632 585
R1012 B.n632 B.n631 585
R1013 B.n634 B.n314 585
R1014 B.n314 B.n313 585
R1015 B.n636 B.n635 585
R1016 B.n637 B.n636 585
R1017 B.n308 B.n307 585
R1018 B.n309 B.n308 585
R1019 B.n645 B.n644 585
R1020 B.n644 B.n643 585
R1021 B.n646 B.n306 585
R1022 B.n306 B.n305 585
R1023 B.n648 B.n647 585
R1024 B.n649 B.n648 585
R1025 B.n300 B.n299 585
R1026 B.n301 B.n300 585
R1027 B.n658 B.n657 585
R1028 B.n657 B.n656 585
R1029 B.n659 B.n298 585
R1030 B.n298 B.n297 585
R1031 B.n661 B.n660 585
R1032 B.n662 B.n661 585
R1033 B.n2 B.n0 585
R1034 B.n4 B.n2 585
R1035 B.n3 B.n1 585
R1036 B.n749 B.n3 585
R1037 B.n747 B.n746 585
R1038 B.n748 B.n747 585
R1039 B.n745 B.n9 585
R1040 B.n9 B.n8 585
R1041 B.n744 B.n743 585
R1042 B.n743 B.n742 585
R1043 B.n11 B.n10 585
R1044 B.n741 B.n11 585
R1045 B.n739 B.n738 585
R1046 B.n740 B.n739 585
R1047 B.n737 B.n16 585
R1048 B.n16 B.n15 585
R1049 B.n736 B.n735 585
R1050 B.n735 B.n734 585
R1051 B.n18 B.n17 585
R1052 B.n733 B.n18 585
R1053 B.n731 B.n730 585
R1054 B.n732 B.n731 585
R1055 B.n729 B.n23 585
R1056 B.n23 B.n22 585
R1057 B.n728 B.n727 585
R1058 B.n727 B.n726 585
R1059 B.n25 B.n24 585
R1060 B.n725 B.n25 585
R1061 B.n723 B.n722 585
R1062 B.n724 B.n723 585
R1063 B.n721 B.n30 585
R1064 B.n30 B.n29 585
R1065 B.n720 B.n719 585
R1066 B.n719 B.n718 585
R1067 B.n32 B.n31 585
R1068 B.n717 B.n32 585
R1069 B.n715 B.n714 585
R1070 B.n716 B.n715 585
R1071 B.n713 B.n37 585
R1072 B.n37 B.n36 585
R1073 B.n712 B.n711 585
R1074 B.n711 B.n710 585
R1075 B.n39 B.n38 585
R1076 B.n709 B.n39 585
R1077 B.n707 B.n706 585
R1078 B.n708 B.n707 585
R1079 B.n705 B.n44 585
R1080 B.n44 B.n43 585
R1081 B.n704 B.n703 585
R1082 B.n703 B.n702 585
R1083 B.n46 B.n45 585
R1084 B.n701 B.n46 585
R1085 B.n752 B.n751 585
R1086 B.n751 B.n750 585
R1087 B.n395 B.t6 482.752
R1088 B.n393 B.t17 482.752
R1089 B.n100 B.t10 482.752
R1090 B.n98 B.t14 482.752
R1091 B.n586 B.n340 430.038
R1092 B.n103 B.n46 430.038
R1093 B.n590 B.n342 430.038
R1094 B.n699 B.n48 430.038
R1095 B.n395 B.t9 320.291
R1096 B.n98 B.t15 320.291
R1097 B.n393 B.t19 320.291
R1098 B.n100 B.t12 320.291
R1099 B.n396 B.t8 292.75
R1100 B.n99 B.t16 292.75
R1101 B.n394 B.t18 292.75
R1102 B.n101 B.t13 292.75
R1103 B.n700 B.n96 256.663
R1104 B.n700 B.n95 256.663
R1105 B.n700 B.n94 256.663
R1106 B.n700 B.n93 256.663
R1107 B.n700 B.n92 256.663
R1108 B.n700 B.n91 256.663
R1109 B.n700 B.n90 256.663
R1110 B.n700 B.n89 256.663
R1111 B.n700 B.n88 256.663
R1112 B.n700 B.n87 256.663
R1113 B.n700 B.n86 256.663
R1114 B.n700 B.n85 256.663
R1115 B.n700 B.n84 256.663
R1116 B.n700 B.n83 256.663
R1117 B.n700 B.n82 256.663
R1118 B.n700 B.n81 256.663
R1119 B.n700 B.n80 256.663
R1120 B.n700 B.n79 256.663
R1121 B.n700 B.n78 256.663
R1122 B.n700 B.n77 256.663
R1123 B.n700 B.n76 256.663
R1124 B.n700 B.n75 256.663
R1125 B.n700 B.n74 256.663
R1126 B.n700 B.n73 256.663
R1127 B.n700 B.n72 256.663
R1128 B.n700 B.n71 256.663
R1129 B.n700 B.n70 256.663
R1130 B.n700 B.n69 256.663
R1131 B.n700 B.n68 256.663
R1132 B.n700 B.n67 256.663
R1133 B.n700 B.n66 256.663
R1134 B.n700 B.n65 256.663
R1135 B.n700 B.n64 256.663
R1136 B.n700 B.n63 256.663
R1137 B.n700 B.n62 256.663
R1138 B.n700 B.n61 256.663
R1139 B.n700 B.n60 256.663
R1140 B.n700 B.n59 256.663
R1141 B.n700 B.n58 256.663
R1142 B.n700 B.n57 256.663
R1143 B.n700 B.n56 256.663
R1144 B.n700 B.n55 256.663
R1145 B.n700 B.n54 256.663
R1146 B.n700 B.n53 256.663
R1147 B.n700 B.n52 256.663
R1148 B.n700 B.n51 256.663
R1149 B.n700 B.n50 256.663
R1150 B.n700 B.n49 256.663
R1151 B.n588 B.n587 256.663
R1152 B.n588 B.n345 256.663
R1153 B.n588 B.n346 256.663
R1154 B.n588 B.n347 256.663
R1155 B.n588 B.n348 256.663
R1156 B.n588 B.n349 256.663
R1157 B.n588 B.n350 256.663
R1158 B.n588 B.n351 256.663
R1159 B.n588 B.n352 256.663
R1160 B.n588 B.n353 256.663
R1161 B.n588 B.n354 256.663
R1162 B.n588 B.n355 256.663
R1163 B.n588 B.n356 256.663
R1164 B.n588 B.n357 256.663
R1165 B.n588 B.n358 256.663
R1166 B.n588 B.n359 256.663
R1167 B.n588 B.n360 256.663
R1168 B.n588 B.n361 256.663
R1169 B.n588 B.n362 256.663
R1170 B.n588 B.n363 256.663
R1171 B.n588 B.n364 256.663
R1172 B.n588 B.n365 256.663
R1173 B.n588 B.n366 256.663
R1174 B.n588 B.n367 256.663
R1175 B.n588 B.n368 256.663
R1176 B.n588 B.n369 256.663
R1177 B.n588 B.n370 256.663
R1178 B.n588 B.n371 256.663
R1179 B.n588 B.n372 256.663
R1180 B.n588 B.n373 256.663
R1181 B.n588 B.n374 256.663
R1182 B.n588 B.n375 256.663
R1183 B.n588 B.n376 256.663
R1184 B.n588 B.n377 256.663
R1185 B.n588 B.n378 256.663
R1186 B.n588 B.n379 256.663
R1187 B.n588 B.n380 256.663
R1188 B.n588 B.n381 256.663
R1189 B.n588 B.n382 256.663
R1190 B.n588 B.n383 256.663
R1191 B.n588 B.n384 256.663
R1192 B.n588 B.n385 256.663
R1193 B.n588 B.n386 256.663
R1194 B.n588 B.n387 256.663
R1195 B.n588 B.n388 256.663
R1196 B.n588 B.n389 256.663
R1197 B.n588 B.n390 256.663
R1198 B.n589 B.n588 256.663
R1199 B.n596 B.n340 163.367
R1200 B.n596 B.n338 163.367
R1201 B.n600 B.n338 163.367
R1202 B.n600 B.n332 163.367
R1203 B.n608 B.n332 163.367
R1204 B.n608 B.n330 163.367
R1205 B.n612 B.n330 163.367
R1206 B.n612 B.n324 163.367
R1207 B.n620 B.n324 163.367
R1208 B.n620 B.n322 163.367
R1209 B.n624 B.n322 163.367
R1210 B.n624 B.n316 163.367
R1211 B.n632 B.n316 163.367
R1212 B.n632 B.n314 163.367
R1213 B.n636 B.n314 163.367
R1214 B.n636 B.n308 163.367
R1215 B.n644 B.n308 163.367
R1216 B.n644 B.n306 163.367
R1217 B.n648 B.n306 163.367
R1218 B.n648 B.n300 163.367
R1219 B.n657 B.n300 163.367
R1220 B.n657 B.n298 163.367
R1221 B.n661 B.n298 163.367
R1222 B.n661 B.n2 163.367
R1223 B.n751 B.n2 163.367
R1224 B.n751 B.n3 163.367
R1225 B.n747 B.n3 163.367
R1226 B.n747 B.n9 163.367
R1227 B.n743 B.n9 163.367
R1228 B.n743 B.n11 163.367
R1229 B.n739 B.n11 163.367
R1230 B.n739 B.n16 163.367
R1231 B.n735 B.n16 163.367
R1232 B.n735 B.n18 163.367
R1233 B.n731 B.n18 163.367
R1234 B.n731 B.n23 163.367
R1235 B.n727 B.n23 163.367
R1236 B.n727 B.n25 163.367
R1237 B.n723 B.n25 163.367
R1238 B.n723 B.n30 163.367
R1239 B.n719 B.n30 163.367
R1240 B.n719 B.n32 163.367
R1241 B.n715 B.n32 163.367
R1242 B.n715 B.n37 163.367
R1243 B.n711 B.n37 163.367
R1244 B.n711 B.n39 163.367
R1245 B.n707 B.n39 163.367
R1246 B.n707 B.n44 163.367
R1247 B.n703 B.n44 163.367
R1248 B.n703 B.n46 163.367
R1249 B.n392 B.n391 163.367
R1250 B.n581 B.n391 163.367
R1251 B.n579 B.n578 163.367
R1252 B.n575 B.n574 163.367
R1253 B.n571 B.n570 163.367
R1254 B.n567 B.n566 163.367
R1255 B.n563 B.n562 163.367
R1256 B.n559 B.n558 163.367
R1257 B.n555 B.n554 163.367
R1258 B.n551 B.n550 163.367
R1259 B.n547 B.n546 163.367
R1260 B.n543 B.n542 163.367
R1261 B.n539 B.n538 163.367
R1262 B.n535 B.n534 163.367
R1263 B.n531 B.n530 163.367
R1264 B.n527 B.n526 163.367
R1265 B.n523 B.n522 163.367
R1266 B.n519 B.n518 163.367
R1267 B.n515 B.n514 163.367
R1268 B.n511 B.n510 163.367
R1269 B.n507 B.n506 163.367
R1270 B.n503 B.n502 163.367
R1271 B.n498 B.n497 163.367
R1272 B.n494 B.n493 163.367
R1273 B.n490 B.n489 163.367
R1274 B.n486 B.n485 163.367
R1275 B.n482 B.n481 163.367
R1276 B.n478 B.n477 163.367
R1277 B.n474 B.n473 163.367
R1278 B.n470 B.n469 163.367
R1279 B.n466 B.n465 163.367
R1280 B.n462 B.n461 163.367
R1281 B.n458 B.n457 163.367
R1282 B.n454 B.n453 163.367
R1283 B.n450 B.n449 163.367
R1284 B.n446 B.n445 163.367
R1285 B.n442 B.n441 163.367
R1286 B.n438 B.n437 163.367
R1287 B.n434 B.n433 163.367
R1288 B.n430 B.n429 163.367
R1289 B.n426 B.n425 163.367
R1290 B.n422 B.n421 163.367
R1291 B.n418 B.n417 163.367
R1292 B.n414 B.n413 163.367
R1293 B.n410 B.n409 163.367
R1294 B.n406 B.n405 163.367
R1295 B.n402 B.n401 163.367
R1296 B.n398 B.n344 163.367
R1297 B.n594 B.n342 163.367
R1298 B.n594 B.n336 163.367
R1299 B.n602 B.n336 163.367
R1300 B.n602 B.n334 163.367
R1301 B.n606 B.n334 163.367
R1302 B.n606 B.n328 163.367
R1303 B.n614 B.n328 163.367
R1304 B.n614 B.n326 163.367
R1305 B.n618 B.n326 163.367
R1306 B.n618 B.n319 163.367
R1307 B.n626 B.n319 163.367
R1308 B.n626 B.n317 163.367
R1309 B.n630 B.n317 163.367
R1310 B.n630 B.n312 163.367
R1311 B.n638 B.n312 163.367
R1312 B.n638 B.n310 163.367
R1313 B.n642 B.n310 163.367
R1314 B.n642 B.n304 163.367
R1315 B.n650 B.n304 163.367
R1316 B.n650 B.n302 163.367
R1317 B.n655 B.n302 163.367
R1318 B.n655 B.n296 163.367
R1319 B.n663 B.n296 163.367
R1320 B.n664 B.n663 163.367
R1321 B.n664 B.n5 163.367
R1322 B.n6 B.n5 163.367
R1323 B.n7 B.n6 163.367
R1324 B.n669 B.n7 163.367
R1325 B.n669 B.n12 163.367
R1326 B.n13 B.n12 163.367
R1327 B.n14 B.n13 163.367
R1328 B.n674 B.n14 163.367
R1329 B.n674 B.n19 163.367
R1330 B.n20 B.n19 163.367
R1331 B.n21 B.n20 163.367
R1332 B.n679 B.n21 163.367
R1333 B.n679 B.n26 163.367
R1334 B.n27 B.n26 163.367
R1335 B.n28 B.n27 163.367
R1336 B.n684 B.n28 163.367
R1337 B.n684 B.n33 163.367
R1338 B.n34 B.n33 163.367
R1339 B.n35 B.n34 163.367
R1340 B.n689 B.n35 163.367
R1341 B.n689 B.n40 163.367
R1342 B.n41 B.n40 163.367
R1343 B.n42 B.n41 163.367
R1344 B.n694 B.n42 163.367
R1345 B.n694 B.n47 163.367
R1346 B.n48 B.n47 163.367
R1347 B.n107 B.n106 163.367
R1348 B.n111 B.n110 163.367
R1349 B.n115 B.n114 163.367
R1350 B.n119 B.n118 163.367
R1351 B.n123 B.n122 163.367
R1352 B.n127 B.n126 163.367
R1353 B.n131 B.n130 163.367
R1354 B.n135 B.n134 163.367
R1355 B.n139 B.n138 163.367
R1356 B.n143 B.n142 163.367
R1357 B.n147 B.n146 163.367
R1358 B.n151 B.n150 163.367
R1359 B.n155 B.n154 163.367
R1360 B.n159 B.n158 163.367
R1361 B.n163 B.n162 163.367
R1362 B.n167 B.n166 163.367
R1363 B.n171 B.n170 163.367
R1364 B.n175 B.n174 163.367
R1365 B.n179 B.n178 163.367
R1366 B.n183 B.n182 163.367
R1367 B.n187 B.n186 163.367
R1368 B.n191 B.n190 163.367
R1369 B.n195 B.n194 163.367
R1370 B.n199 B.n198 163.367
R1371 B.n203 B.n202 163.367
R1372 B.n207 B.n206 163.367
R1373 B.n212 B.n211 163.367
R1374 B.n216 B.n215 163.367
R1375 B.n220 B.n219 163.367
R1376 B.n224 B.n223 163.367
R1377 B.n228 B.n227 163.367
R1378 B.n232 B.n231 163.367
R1379 B.n236 B.n235 163.367
R1380 B.n240 B.n239 163.367
R1381 B.n244 B.n243 163.367
R1382 B.n248 B.n247 163.367
R1383 B.n252 B.n251 163.367
R1384 B.n256 B.n255 163.367
R1385 B.n260 B.n259 163.367
R1386 B.n264 B.n263 163.367
R1387 B.n268 B.n267 163.367
R1388 B.n272 B.n271 163.367
R1389 B.n276 B.n275 163.367
R1390 B.n280 B.n279 163.367
R1391 B.n284 B.n283 163.367
R1392 B.n288 B.n287 163.367
R1393 B.n292 B.n291 163.367
R1394 B.n699 B.n97 163.367
R1395 B.n587 B.n586 71.676
R1396 B.n581 B.n345 71.676
R1397 B.n578 B.n346 71.676
R1398 B.n574 B.n347 71.676
R1399 B.n570 B.n348 71.676
R1400 B.n566 B.n349 71.676
R1401 B.n562 B.n350 71.676
R1402 B.n558 B.n351 71.676
R1403 B.n554 B.n352 71.676
R1404 B.n550 B.n353 71.676
R1405 B.n546 B.n354 71.676
R1406 B.n542 B.n355 71.676
R1407 B.n538 B.n356 71.676
R1408 B.n534 B.n357 71.676
R1409 B.n530 B.n358 71.676
R1410 B.n526 B.n359 71.676
R1411 B.n522 B.n360 71.676
R1412 B.n518 B.n361 71.676
R1413 B.n514 B.n362 71.676
R1414 B.n510 B.n363 71.676
R1415 B.n506 B.n364 71.676
R1416 B.n502 B.n365 71.676
R1417 B.n497 B.n366 71.676
R1418 B.n493 B.n367 71.676
R1419 B.n489 B.n368 71.676
R1420 B.n485 B.n369 71.676
R1421 B.n481 B.n370 71.676
R1422 B.n477 B.n371 71.676
R1423 B.n473 B.n372 71.676
R1424 B.n469 B.n373 71.676
R1425 B.n465 B.n374 71.676
R1426 B.n461 B.n375 71.676
R1427 B.n457 B.n376 71.676
R1428 B.n453 B.n377 71.676
R1429 B.n449 B.n378 71.676
R1430 B.n445 B.n379 71.676
R1431 B.n441 B.n380 71.676
R1432 B.n437 B.n381 71.676
R1433 B.n433 B.n382 71.676
R1434 B.n429 B.n383 71.676
R1435 B.n425 B.n384 71.676
R1436 B.n421 B.n385 71.676
R1437 B.n417 B.n386 71.676
R1438 B.n413 B.n387 71.676
R1439 B.n409 B.n388 71.676
R1440 B.n405 B.n389 71.676
R1441 B.n401 B.n390 71.676
R1442 B.n589 B.n344 71.676
R1443 B.n103 B.n49 71.676
R1444 B.n107 B.n50 71.676
R1445 B.n111 B.n51 71.676
R1446 B.n115 B.n52 71.676
R1447 B.n119 B.n53 71.676
R1448 B.n123 B.n54 71.676
R1449 B.n127 B.n55 71.676
R1450 B.n131 B.n56 71.676
R1451 B.n135 B.n57 71.676
R1452 B.n139 B.n58 71.676
R1453 B.n143 B.n59 71.676
R1454 B.n147 B.n60 71.676
R1455 B.n151 B.n61 71.676
R1456 B.n155 B.n62 71.676
R1457 B.n159 B.n63 71.676
R1458 B.n163 B.n64 71.676
R1459 B.n167 B.n65 71.676
R1460 B.n171 B.n66 71.676
R1461 B.n175 B.n67 71.676
R1462 B.n179 B.n68 71.676
R1463 B.n183 B.n69 71.676
R1464 B.n187 B.n70 71.676
R1465 B.n191 B.n71 71.676
R1466 B.n195 B.n72 71.676
R1467 B.n199 B.n73 71.676
R1468 B.n203 B.n74 71.676
R1469 B.n207 B.n75 71.676
R1470 B.n212 B.n76 71.676
R1471 B.n216 B.n77 71.676
R1472 B.n220 B.n78 71.676
R1473 B.n224 B.n79 71.676
R1474 B.n228 B.n80 71.676
R1475 B.n232 B.n81 71.676
R1476 B.n236 B.n82 71.676
R1477 B.n240 B.n83 71.676
R1478 B.n244 B.n84 71.676
R1479 B.n248 B.n85 71.676
R1480 B.n252 B.n86 71.676
R1481 B.n256 B.n87 71.676
R1482 B.n260 B.n88 71.676
R1483 B.n264 B.n89 71.676
R1484 B.n268 B.n90 71.676
R1485 B.n272 B.n91 71.676
R1486 B.n276 B.n92 71.676
R1487 B.n280 B.n93 71.676
R1488 B.n284 B.n94 71.676
R1489 B.n288 B.n95 71.676
R1490 B.n292 B.n96 71.676
R1491 B.n97 B.n96 71.676
R1492 B.n291 B.n95 71.676
R1493 B.n287 B.n94 71.676
R1494 B.n283 B.n93 71.676
R1495 B.n279 B.n92 71.676
R1496 B.n275 B.n91 71.676
R1497 B.n271 B.n90 71.676
R1498 B.n267 B.n89 71.676
R1499 B.n263 B.n88 71.676
R1500 B.n259 B.n87 71.676
R1501 B.n255 B.n86 71.676
R1502 B.n251 B.n85 71.676
R1503 B.n247 B.n84 71.676
R1504 B.n243 B.n83 71.676
R1505 B.n239 B.n82 71.676
R1506 B.n235 B.n81 71.676
R1507 B.n231 B.n80 71.676
R1508 B.n227 B.n79 71.676
R1509 B.n223 B.n78 71.676
R1510 B.n219 B.n77 71.676
R1511 B.n215 B.n76 71.676
R1512 B.n211 B.n75 71.676
R1513 B.n206 B.n74 71.676
R1514 B.n202 B.n73 71.676
R1515 B.n198 B.n72 71.676
R1516 B.n194 B.n71 71.676
R1517 B.n190 B.n70 71.676
R1518 B.n186 B.n69 71.676
R1519 B.n182 B.n68 71.676
R1520 B.n178 B.n67 71.676
R1521 B.n174 B.n66 71.676
R1522 B.n170 B.n65 71.676
R1523 B.n166 B.n64 71.676
R1524 B.n162 B.n63 71.676
R1525 B.n158 B.n62 71.676
R1526 B.n154 B.n61 71.676
R1527 B.n150 B.n60 71.676
R1528 B.n146 B.n59 71.676
R1529 B.n142 B.n58 71.676
R1530 B.n138 B.n57 71.676
R1531 B.n134 B.n56 71.676
R1532 B.n130 B.n55 71.676
R1533 B.n126 B.n54 71.676
R1534 B.n122 B.n53 71.676
R1535 B.n118 B.n52 71.676
R1536 B.n114 B.n51 71.676
R1537 B.n110 B.n50 71.676
R1538 B.n106 B.n49 71.676
R1539 B.n587 B.n392 71.676
R1540 B.n579 B.n345 71.676
R1541 B.n575 B.n346 71.676
R1542 B.n571 B.n347 71.676
R1543 B.n567 B.n348 71.676
R1544 B.n563 B.n349 71.676
R1545 B.n559 B.n350 71.676
R1546 B.n555 B.n351 71.676
R1547 B.n551 B.n352 71.676
R1548 B.n547 B.n353 71.676
R1549 B.n543 B.n354 71.676
R1550 B.n539 B.n355 71.676
R1551 B.n535 B.n356 71.676
R1552 B.n531 B.n357 71.676
R1553 B.n527 B.n358 71.676
R1554 B.n523 B.n359 71.676
R1555 B.n519 B.n360 71.676
R1556 B.n515 B.n361 71.676
R1557 B.n511 B.n362 71.676
R1558 B.n507 B.n363 71.676
R1559 B.n503 B.n364 71.676
R1560 B.n498 B.n365 71.676
R1561 B.n494 B.n366 71.676
R1562 B.n490 B.n367 71.676
R1563 B.n486 B.n368 71.676
R1564 B.n482 B.n369 71.676
R1565 B.n478 B.n370 71.676
R1566 B.n474 B.n371 71.676
R1567 B.n470 B.n372 71.676
R1568 B.n466 B.n373 71.676
R1569 B.n462 B.n374 71.676
R1570 B.n458 B.n375 71.676
R1571 B.n454 B.n376 71.676
R1572 B.n450 B.n377 71.676
R1573 B.n446 B.n378 71.676
R1574 B.n442 B.n379 71.676
R1575 B.n438 B.n380 71.676
R1576 B.n434 B.n381 71.676
R1577 B.n430 B.n382 71.676
R1578 B.n426 B.n383 71.676
R1579 B.n422 B.n384 71.676
R1580 B.n418 B.n385 71.676
R1581 B.n414 B.n386 71.676
R1582 B.n410 B.n387 71.676
R1583 B.n406 B.n388 71.676
R1584 B.n402 B.n389 71.676
R1585 B.n398 B.n390 71.676
R1586 B.n590 B.n589 71.676
R1587 B.n588 B.n341 68.1937
R1588 B.n701 B.n700 68.1937
R1589 B.n397 B.n396 59.5399
R1590 B.n500 B.n394 59.5399
R1591 B.n102 B.n101 59.5399
R1592 B.n209 B.n99 59.5399
R1593 B.n595 B.n341 41.7765
R1594 B.n595 B.n337 41.7765
R1595 B.n601 B.n337 41.7765
R1596 B.n601 B.n333 41.7765
R1597 B.n607 B.n333 41.7765
R1598 B.n613 B.n329 41.7765
R1599 B.n613 B.n325 41.7765
R1600 B.n619 B.n325 41.7765
R1601 B.n619 B.n320 41.7765
R1602 B.n625 B.n320 41.7765
R1603 B.n625 B.n321 41.7765
R1604 B.n631 B.n313 41.7765
R1605 B.n637 B.n313 41.7765
R1606 B.n637 B.n309 41.7765
R1607 B.n643 B.n309 41.7765
R1608 B.n649 B.n305 41.7765
R1609 B.n649 B.n301 41.7765
R1610 B.n656 B.n301 41.7765
R1611 B.n662 B.n297 41.7765
R1612 B.n662 B.n4 41.7765
R1613 B.n750 B.n4 41.7765
R1614 B.n750 B.n749 41.7765
R1615 B.n749 B.n748 41.7765
R1616 B.n748 B.n8 41.7765
R1617 B.n742 B.n741 41.7765
R1618 B.n741 B.n740 41.7765
R1619 B.n740 B.n15 41.7765
R1620 B.n734 B.n733 41.7765
R1621 B.n733 B.n732 41.7765
R1622 B.n732 B.n22 41.7765
R1623 B.n726 B.n22 41.7765
R1624 B.n725 B.n724 41.7765
R1625 B.n724 B.n29 41.7765
R1626 B.n718 B.n29 41.7765
R1627 B.n718 B.n717 41.7765
R1628 B.n717 B.n716 41.7765
R1629 B.n716 B.n36 41.7765
R1630 B.n710 B.n709 41.7765
R1631 B.n709 B.n708 41.7765
R1632 B.n708 B.n43 41.7765
R1633 B.n702 B.n43 41.7765
R1634 B.n702 B.n701 41.7765
R1635 B.n321 B.t1 39.9335
R1636 B.t2 B.n725 39.9335
R1637 B.t3 B.n305 36.2474
R1638 B.t0 B.n15 36.2474
R1639 B.t4 B.n297 28.8751
R1640 B.t5 B.n8 28.8751
R1641 B.n104 B.n45 27.942
R1642 B.n698 B.n697 27.942
R1643 B.n592 B.n591 27.942
R1644 B.n585 B.n339 27.942
R1645 B.n396 B.n395 27.5399
R1646 B.n394 B.n393 27.5399
R1647 B.n101 B.n100 27.5399
R1648 B.n99 B.n98 27.5399
R1649 B.n607 B.t7 23.9603
R1650 B.n710 B.t11 23.9603
R1651 B B.n752 18.0485
R1652 B.t7 B.n329 17.8168
R1653 B.t11 B.n36 17.8168
R1654 B.n656 B.t4 12.9019
R1655 B.n742 B.t5 12.9019
R1656 B.n105 B.n104 10.6151
R1657 B.n108 B.n105 10.6151
R1658 B.n109 B.n108 10.6151
R1659 B.n112 B.n109 10.6151
R1660 B.n113 B.n112 10.6151
R1661 B.n116 B.n113 10.6151
R1662 B.n117 B.n116 10.6151
R1663 B.n120 B.n117 10.6151
R1664 B.n121 B.n120 10.6151
R1665 B.n124 B.n121 10.6151
R1666 B.n125 B.n124 10.6151
R1667 B.n128 B.n125 10.6151
R1668 B.n129 B.n128 10.6151
R1669 B.n132 B.n129 10.6151
R1670 B.n133 B.n132 10.6151
R1671 B.n136 B.n133 10.6151
R1672 B.n137 B.n136 10.6151
R1673 B.n140 B.n137 10.6151
R1674 B.n141 B.n140 10.6151
R1675 B.n144 B.n141 10.6151
R1676 B.n145 B.n144 10.6151
R1677 B.n148 B.n145 10.6151
R1678 B.n149 B.n148 10.6151
R1679 B.n152 B.n149 10.6151
R1680 B.n153 B.n152 10.6151
R1681 B.n156 B.n153 10.6151
R1682 B.n157 B.n156 10.6151
R1683 B.n160 B.n157 10.6151
R1684 B.n161 B.n160 10.6151
R1685 B.n164 B.n161 10.6151
R1686 B.n165 B.n164 10.6151
R1687 B.n168 B.n165 10.6151
R1688 B.n169 B.n168 10.6151
R1689 B.n172 B.n169 10.6151
R1690 B.n173 B.n172 10.6151
R1691 B.n176 B.n173 10.6151
R1692 B.n177 B.n176 10.6151
R1693 B.n180 B.n177 10.6151
R1694 B.n181 B.n180 10.6151
R1695 B.n184 B.n181 10.6151
R1696 B.n185 B.n184 10.6151
R1697 B.n188 B.n185 10.6151
R1698 B.n189 B.n188 10.6151
R1699 B.n193 B.n192 10.6151
R1700 B.n196 B.n193 10.6151
R1701 B.n197 B.n196 10.6151
R1702 B.n200 B.n197 10.6151
R1703 B.n201 B.n200 10.6151
R1704 B.n204 B.n201 10.6151
R1705 B.n205 B.n204 10.6151
R1706 B.n208 B.n205 10.6151
R1707 B.n213 B.n210 10.6151
R1708 B.n214 B.n213 10.6151
R1709 B.n217 B.n214 10.6151
R1710 B.n218 B.n217 10.6151
R1711 B.n221 B.n218 10.6151
R1712 B.n222 B.n221 10.6151
R1713 B.n225 B.n222 10.6151
R1714 B.n226 B.n225 10.6151
R1715 B.n229 B.n226 10.6151
R1716 B.n230 B.n229 10.6151
R1717 B.n233 B.n230 10.6151
R1718 B.n234 B.n233 10.6151
R1719 B.n237 B.n234 10.6151
R1720 B.n238 B.n237 10.6151
R1721 B.n241 B.n238 10.6151
R1722 B.n242 B.n241 10.6151
R1723 B.n245 B.n242 10.6151
R1724 B.n246 B.n245 10.6151
R1725 B.n249 B.n246 10.6151
R1726 B.n250 B.n249 10.6151
R1727 B.n253 B.n250 10.6151
R1728 B.n254 B.n253 10.6151
R1729 B.n257 B.n254 10.6151
R1730 B.n258 B.n257 10.6151
R1731 B.n261 B.n258 10.6151
R1732 B.n262 B.n261 10.6151
R1733 B.n265 B.n262 10.6151
R1734 B.n266 B.n265 10.6151
R1735 B.n269 B.n266 10.6151
R1736 B.n270 B.n269 10.6151
R1737 B.n273 B.n270 10.6151
R1738 B.n274 B.n273 10.6151
R1739 B.n277 B.n274 10.6151
R1740 B.n278 B.n277 10.6151
R1741 B.n281 B.n278 10.6151
R1742 B.n282 B.n281 10.6151
R1743 B.n285 B.n282 10.6151
R1744 B.n286 B.n285 10.6151
R1745 B.n289 B.n286 10.6151
R1746 B.n290 B.n289 10.6151
R1747 B.n293 B.n290 10.6151
R1748 B.n294 B.n293 10.6151
R1749 B.n698 B.n294 10.6151
R1750 B.n593 B.n592 10.6151
R1751 B.n593 B.n335 10.6151
R1752 B.n603 B.n335 10.6151
R1753 B.n604 B.n603 10.6151
R1754 B.n605 B.n604 10.6151
R1755 B.n605 B.n327 10.6151
R1756 B.n615 B.n327 10.6151
R1757 B.n616 B.n615 10.6151
R1758 B.n617 B.n616 10.6151
R1759 B.n617 B.n318 10.6151
R1760 B.n627 B.n318 10.6151
R1761 B.n628 B.n627 10.6151
R1762 B.n629 B.n628 10.6151
R1763 B.n629 B.n311 10.6151
R1764 B.n639 B.n311 10.6151
R1765 B.n640 B.n639 10.6151
R1766 B.n641 B.n640 10.6151
R1767 B.n641 B.n303 10.6151
R1768 B.n651 B.n303 10.6151
R1769 B.n652 B.n651 10.6151
R1770 B.n654 B.n652 10.6151
R1771 B.n654 B.n653 10.6151
R1772 B.n653 B.n295 10.6151
R1773 B.n665 B.n295 10.6151
R1774 B.n666 B.n665 10.6151
R1775 B.n667 B.n666 10.6151
R1776 B.n668 B.n667 10.6151
R1777 B.n670 B.n668 10.6151
R1778 B.n671 B.n670 10.6151
R1779 B.n672 B.n671 10.6151
R1780 B.n673 B.n672 10.6151
R1781 B.n675 B.n673 10.6151
R1782 B.n676 B.n675 10.6151
R1783 B.n677 B.n676 10.6151
R1784 B.n678 B.n677 10.6151
R1785 B.n680 B.n678 10.6151
R1786 B.n681 B.n680 10.6151
R1787 B.n682 B.n681 10.6151
R1788 B.n683 B.n682 10.6151
R1789 B.n685 B.n683 10.6151
R1790 B.n686 B.n685 10.6151
R1791 B.n687 B.n686 10.6151
R1792 B.n688 B.n687 10.6151
R1793 B.n690 B.n688 10.6151
R1794 B.n691 B.n690 10.6151
R1795 B.n692 B.n691 10.6151
R1796 B.n693 B.n692 10.6151
R1797 B.n695 B.n693 10.6151
R1798 B.n696 B.n695 10.6151
R1799 B.n697 B.n696 10.6151
R1800 B.n585 B.n584 10.6151
R1801 B.n584 B.n583 10.6151
R1802 B.n583 B.n582 10.6151
R1803 B.n582 B.n580 10.6151
R1804 B.n580 B.n577 10.6151
R1805 B.n577 B.n576 10.6151
R1806 B.n576 B.n573 10.6151
R1807 B.n573 B.n572 10.6151
R1808 B.n572 B.n569 10.6151
R1809 B.n569 B.n568 10.6151
R1810 B.n568 B.n565 10.6151
R1811 B.n565 B.n564 10.6151
R1812 B.n564 B.n561 10.6151
R1813 B.n561 B.n560 10.6151
R1814 B.n560 B.n557 10.6151
R1815 B.n557 B.n556 10.6151
R1816 B.n556 B.n553 10.6151
R1817 B.n553 B.n552 10.6151
R1818 B.n552 B.n549 10.6151
R1819 B.n549 B.n548 10.6151
R1820 B.n548 B.n545 10.6151
R1821 B.n545 B.n544 10.6151
R1822 B.n544 B.n541 10.6151
R1823 B.n541 B.n540 10.6151
R1824 B.n540 B.n537 10.6151
R1825 B.n537 B.n536 10.6151
R1826 B.n536 B.n533 10.6151
R1827 B.n533 B.n532 10.6151
R1828 B.n532 B.n529 10.6151
R1829 B.n529 B.n528 10.6151
R1830 B.n528 B.n525 10.6151
R1831 B.n525 B.n524 10.6151
R1832 B.n524 B.n521 10.6151
R1833 B.n521 B.n520 10.6151
R1834 B.n520 B.n517 10.6151
R1835 B.n517 B.n516 10.6151
R1836 B.n516 B.n513 10.6151
R1837 B.n513 B.n512 10.6151
R1838 B.n512 B.n509 10.6151
R1839 B.n509 B.n508 10.6151
R1840 B.n508 B.n505 10.6151
R1841 B.n505 B.n504 10.6151
R1842 B.n504 B.n501 10.6151
R1843 B.n499 B.n496 10.6151
R1844 B.n496 B.n495 10.6151
R1845 B.n495 B.n492 10.6151
R1846 B.n492 B.n491 10.6151
R1847 B.n491 B.n488 10.6151
R1848 B.n488 B.n487 10.6151
R1849 B.n487 B.n484 10.6151
R1850 B.n484 B.n483 10.6151
R1851 B.n480 B.n479 10.6151
R1852 B.n479 B.n476 10.6151
R1853 B.n476 B.n475 10.6151
R1854 B.n475 B.n472 10.6151
R1855 B.n472 B.n471 10.6151
R1856 B.n471 B.n468 10.6151
R1857 B.n468 B.n467 10.6151
R1858 B.n467 B.n464 10.6151
R1859 B.n464 B.n463 10.6151
R1860 B.n463 B.n460 10.6151
R1861 B.n460 B.n459 10.6151
R1862 B.n459 B.n456 10.6151
R1863 B.n456 B.n455 10.6151
R1864 B.n455 B.n452 10.6151
R1865 B.n452 B.n451 10.6151
R1866 B.n451 B.n448 10.6151
R1867 B.n448 B.n447 10.6151
R1868 B.n447 B.n444 10.6151
R1869 B.n444 B.n443 10.6151
R1870 B.n443 B.n440 10.6151
R1871 B.n440 B.n439 10.6151
R1872 B.n439 B.n436 10.6151
R1873 B.n436 B.n435 10.6151
R1874 B.n435 B.n432 10.6151
R1875 B.n432 B.n431 10.6151
R1876 B.n431 B.n428 10.6151
R1877 B.n428 B.n427 10.6151
R1878 B.n427 B.n424 10.6151
R1879 B.n424 B.n423 10.6151
R1880 B.n423 B.n420 10.6151
R1881 B.n420 B.n419 10.6151
R1882 B.n419 B.n416 10.6151
R1883 B.n416 B.n415 10.6151
R1884 B.n415 B.n412 10.6151
R1885 B.n412 B.n411 10.6151
R1886 B.n411 B.n408 10.6151
R1887 B.n408 B.n407 10.6151
R1888 B.n407 B.n404 10.6151
R1889 B.n404 B.n403 10.6151
R1890 B.n403 B.n400 10.6151
R1891 B.n400 B.n399 10.6151
R1892 B.n399 B.n343 10.6151
R1893 B.n591 B.n343 10.6151
R1894 B.n597 B.n339 10.6151
R1895 B.n598 B.n597 10.6151
R1896 B.n599 B.n598 10.6151
R1897 B.n599 B.n331 10.6151
R1898 B.n609 B.n331 10.6151
R1899 B.n610 B.n609 10.6151
R1900 B.n611 B.n610 10.6151
R1901 B.n611 B.n323 10.6151
R1902 B.n621 B.n323 10.6151
R1903 B.n622 B.n621 10.6151
R1904 B.n623 B.n622 10.6151
R1905 B.n623 B.n315 10.6151
R1906 B.n633 B.n315 10.6151
R1907 B.n634 B.n633 10.6151
R1908 B.n635 B.n634 10.6151
R1909 B.n635 B.n307 10.6151
R1910 B.n645 B.n307 10.6151
R1911 B.n646 B.n645 10.6151
R1912 B.n647 B.n646 10.6151
R1913 B.n647 B.n299 10.6151
R1914 B.n658 B.n299 10.6151
R1915 B.n659 B.n658 10.6151
R1916 B.n660 B.n659 10.6151
R1917 B.n660 B.n0 10.6151
R1918 B.n746 B.n1 10.6151
R1919 B.n746 B.n745 10.6151
R1920 B.n745 B.n744 10.6151
R1921 B.n744 B.n10 10.6151
R1922 B.n738 B.n10 10.6151
R1923 B.n738 B.n737 10.6151
R1924 B.n737 B.n736 10.6151
R1925 B.n736 B.n17 10.6151
R1926 B.n730 B.n17 10.6151
R1927 B.n730 B.n729 10.6151
R1928 B.n729 B.n728 10.6151
R1929 B.n728 B.n24 10.6151
R1930 B.n722 B.n24 10.6151
R1931 B.n722 B.n721 10.6151
R1932 B.n721 B.n720 10.6151
R1933 B.n720 B.n31 10.6151
R1934 B.n714 B.n31 10.6151
R1935 B.n714 B.n713 10.6151
R1936 B.n713 B.n712 10.6151
R1937 B.n712 B.n38 10.6151
R1938 B.n706 B.n38 10.6151
R1939 B.n706 B.n705 10.6151
R1940 B.n705 B.n704 10.6151
R1941 B.n704 B.n45 10.6151
R1942 B.n192 B.n102 6.5566
R1943 B.n209 B.n208 6.5566
R1944 B.n500 B.n499 6.5566
R1945 B.n483 B.n397 6.5566
R1946 B.n643 B.t3 5.52968
R1947 B.n734 B.t0 5.52968
R1948 B.n189 B.n102 4.05904
R1949 B.n210 B.n209 4.05904
R1950 B.n501 B.n500 4.05904
R1951 B.n480 B.n397 4.05904
R1952 B.n752 B.n0 2.81026
R1953 B.n752 B.n1 2.81026
R1954 B.n631 B.t1 1.84356
R1955 B.n726 B.t2 1.84356
R1956 VN.n1 VN.t3 338.505
R1957 VN.n7 VN.t4 338.505
R1958 VN.n4 VN.t2 315.512
R1959 VN.n10 VN.t0 315.512
R1960 VN.n2 VN.t1 279.25
R1961 VN.n8 VN.t5 279.25
R1962 VN.n9 VN.n6 161.3
R1963 VN.n3 VN.n0 161.3
R1964 VN.n11 VN.n10 80.6037
R1965 VN.n5 VN.n4 80.6037
R1966 VN.n4 VN.n3 50.4025
R1967 VN.n10 VN.n9 50.4025
R1968 VN VN.n11 43.696
R1969 VN.n2 VN.n1 32.6271
R1970 VN.n8 VN.n7 32.6271
R1971 VN.n7 VN.n6 28.1515
R1972 VN.n1 VN.n0 28.1515
R1973 VN.n3 VN.n2 24.4675
R1974 VN.n9 VN.n8 24.4675
R1975 VN.n11 VN.n6 0.285035
R1976 VN.n5 VN.n0 0.285035
R1977 VN VN.n5 0.146778
R1978 VDD2.n139 VDD2.n138 289.615
R1979 VDD2.n68 VDD2.n67 289.615
R1980 VDD2.n138 VDD2.n137 185
R1981 VDD2.n73 VDD2.n72 185
R1982 VDD2.n132 VDD2.n131 185
R1983 VDD2.n130 VDD2.n129 185
R1984 VDD2.n77 VDD2.n76 185
R1985 VDD2.n124 VDD2.n123 185
R1986 VDD2.n122 VDD2.n121 185
R1987 VDD2.n81 VDD2.n80 185
R1988 VDD2.n116 VDD2.n115 185
R1989 VDD2.n114 VDD2.n113 185
R1990 VDD2.n85 VDD2.n84 185
R1991 VDD2.n108 VDD2.n107 185
R1992 VDD2.n106 VDD2.n105 185
R1993 VDD2.n89 VDD2.n88 185
R1994 VDD2.n100 VDD2.n99 185
R1995 VDD2.n98 VDD2.n97 185
R1996 VDD2.n93 VDD2.n92 185
R1997 VDD2.n22 VDD2.n21 185
R1998 VDD2.n27 VDD2.n26 185
R1999 VDD2.n29 VDD2.n28 185
R2000 VDD2.n18 VDD2.n17 185
R2001 VDD2.n35 VDD2.n34 185
R2002 VDD2.n37 VDD2.n36 185
R2003 VDD2.n14 VDD2.n13 185
R2004 VDD2.n43 VDD2.n42 185
R2005 VDD2.n45 VDD2.n44 185
R2006 VDD2.n10 VDD2.n9 185
R2007 VDD2.n51 VDD2.n50 185
R2008 VDD2.n53 VDD2.n52 185
R2009 VDD2.n6 VDD2.n5 185
R2010 VDD2.n59 VDD2.n58 185
R2011 VDD2.n61 VDD2.n60 185
R2012 VDD2.n2 VDD2.n1 185
R2013 VDD2.n67 VDD2.n66 185
R2014 VDD2.n23 VDD2.t2 147.659
R2015 VDD2.n94 VDD2.t5 147.659
R2016 VDD2.n138 VDD2.n72 104.615
R2017 VDD2.n131 VDD2.n72 104.615
R2018 VDD2.n131 VDD2.n130 104.615
R2019 VDD2.n130 VDD2.n76 104.615
R2020 VDD2.n123 VDD2.n76 104.615
R2021 VDD2.n123 VDD2.n122 104.615
R2022 VDD2.n122 VDD2.n80 104.615
R2023 VDD2.n115 VDD2.n80 104.615
R2024 VDD2.n115 VDD2.n114 104.615
R2025 VDD2.n114 VDD2.n84 104.615
R2026 VDD2.n107 VDD2.n84 104.615
R2027 VDD2.n107 VDD2.n106 104.615
R2028 VDD2.n106 VDD2.n88 104.615
R2029 VDD2.n99 VDD2.n88 104.615
R2030 VDD2.n99 VDD2.n98 104.615
R2031 VDD2.n98 VDD2.n92 104.615
R2032 VDD2.n27 VDD2.n21 104.615
R2033 VDD2.n28 VDD2.n27 104.615
R2034 VDD2.n28 VDD2.n17 104.615
R2035 VDD2.n35 VDD2.n17 104.615
R2036 VDD2.n36 VDD2.n35 104.615
R2037 VDD2.n36 VDD2.n13 104.615
R2038 VDD2.n43 VDD2.n13 104.615
R2039 VDD2.n44 VDD2.n43 104.615
R2040 VDD2.n44 VDD2.n9 104.615
R2041 VDD2.n51 VDD2.n9 104.615
R2042 VDD2.n52 VDD2.n51 104.615
R2043 VDD2.n52 VDD2.n5 104.615
R2044 VDD2.n59 VDD2.n5 104.615
R2045 VDD2.n60 VDD2.n59 104.615
R2046 VDD2.n60 VDD2.n1 104.615
R2047 VDD2.n67 VDD2.n1 104.615
R2048 VDD2.n70 VDD2.n69 64.3672
R2049 VDD2 VDD2.n141 64.3643
R2050 VDD2.t5 VDD2.n92 52.3082
R2051 VDD2.t2 VDD2.n21 52.3082
R2052 VDD2.n70 VDD2.n68 52.2481
R2053 VDD2.n140 VDD2.n139 51.3853
R2054 VDD2.n140 VDD2.n70 38.5817
R2055 VDD2.n94 VDD2.n93 15.6677
R2056 VDD2.n23 VDD2.n22 15.6677
R2057 VDD2.n137 VDD2.n71 12.8005
R2058 VDD2.n97 VDD2.n96 12.8005
R2059 VDD2.n26 VDD2.n25 12.8005
R2060 VDD2.n66 VDD2.n0 12.8005
R2061 VDD2.n136 VDD2.n73 12.0247
R2062 VDD2.n100 VDD2.n91 12.0247
R2063 VDD2.n29 VDD2.n20 12.0247
R2064 VDD2.n65 VDD2.n2 12.0247
R2065 VDD2.n133 VDD2.n132 11.249
R2066 VDD2.n101 VDD2.n89 11.249
R2067 VDD2.n30 VDD2.n18 11.249
R2068 VDD2.n62 VDD2.n61 11.249
R2069 VDD2.n129 VDD2.n75 10.4732
R2070 VDD2.n105 VDD2.n104 10.4732
R2071 VDD2.n34 VDD2.n33 10.4732
R2072 VDD2.n58 VDD2.n4 10.4732
R2073 VDD2.n128 VDD2.n77 9.69747
R2074 VDD2.n108 VDD2.n87 9.69747
R2075 VDD2.n37 VDD2.n16 9.69747
R2076 VDD2.n57 VDD2.n6 9.69747
R2077 VDD2.n135 VDD2.n71 9.45567
R2078 VDD2.n64 VDD2.n0 9.45567
R2079 VDD2.n120 VDD2.n119 9.3005
R2080 VDD2.n79 VDD2.n78 9.3005
R2081 VDD2.n126 VDD2.n125 9.3005
R2082 VDD2.n128 VDD2.n127 9.3005
R2083 VDD2.n75 VDD2.n74 9.3005
R2084 VDD2.n134 VDD2.n133 9.3005
R2085 VDD2.n136 VDD2.n135 9.3005
R2086 VDD2.n118 VDD2.n117 9.3005
R2087 VDD2.n83 VDD2.n82 9.3005
R2088 VDD2.n112 VDD2.n111 9.3005
R2089 VDD2.n110 VDD2.n109 9.3005
R2090 VDD2.n87 VDD2.n86 9.3005
R2091 VDD2.n104 VDD2.n103 9.3005
R2092 VDD2.n102 VDD2.n101 9.3005
R2093 VDD2.n91 VDD2.n90 9.3005
R2094 VDD2.n96 VDD2.n95 9.3005
R2095 VDD2.n47 VDD2.n46 9.3005
R2096 VDD2.n49 VDD2.n48 9.3005
R2097 VDD2.n8 VDD2.n7 9.3005
R2098 VDD2.n55 VDD2.n54 9.3005
R2099 VDD2.n57 VDD2.n56 9.3005
R2100 VDD2.n4 VDD2.n3 9.3005
R2101 VDD2.n63 VDD2.n62 9.3005
R2102 VDD2.n65 VDD2.n64 9.3005
R2103 VDD2.n41 VDD2.n40 9.3005
R2104 VDD2.n39 VDD2.n38 9.3005
R2105 VDD2.n16 VDD2.n15 9.3005
R2106 VDD2.n33 VDD2.n32 9.3005
R2107 VDD2.n31 VDD2.n30 9.3005
R2108 VDD2.n20 VDD2.n19 9.3005
R2109 VDD2.n25 VDD2.n24 9.3005
R2110 VDD2.n12 VDD2.n11 9.3005
R2111 VDD2.n125 VDD2.n124 8.92171
R2112 VDD2.n109 VDD2.n85 8.92171
R2113 VDD2.n38 VDD2.n14 8.92171
R2114 VDD2.n54 VDD2.n53 8.92171
R2115 VDD2.n121 VDD2.n79 8.14595
R2116 VDD2.n113 VDD2.n112 8.14595
R2117 VDD2.n42 VDD2.n41 8.14595
R2118 VDD2.n50 VDD2.n8 8.14595
R2119 VDD2.n120 VDD2.n81 7.3702
R2120 VDD2.n116 VDD2.n83 7.3702
R2121 VDD2.n45 VDD2.n12 7.3702
R2122 VDD2.n49 VDD2.n10 7.3702
R2123 VDD2.n117 VDD2.n81 6.59444
R2124 VDD2.n117 VDD2.n116 6.59444
R2125 VDD2.n46 VDD2.n45 6.59444
R2126 VDD2.n46 VDD2.n10 6.59444
R2127 VDD2.n121 VDD2.n120 5.81868
R2128 VDD2.n113 VDD2.n83 5.81868
R2129 VDD2.n42 VDD2.n12 5.81868
R2130 VDD2.n50 VDD2.n49 5.81868
R2131 VDD2.n124 VDD2.n79 5.04292
R2132 VDD2.n112 VDD2.n85 5.04292
R2133 VDD2.n41 VDD2.n14 5.04292
R2134 VDD2.n53 VDD2.n8 5.04292
R2135 VDD2.n24 VDD2.n23 4.38563
R2136 VDD2.n95 VDD2.n94 4.38563
R2137 VDD2.n125 VDD2.n77 4.26717
R2138 VDD2.n109 VDD2.n108 4.26717
R2139 VDD2.n38 VDD2.n37 4.26717
R2140 VDD2.n54 VDD2.n6 4.26717
R2141 VDD2.n129 VDD2.n128 3.49141
R2142 VDD2.n105 VDD2.n87 3.49141
R2143 VDD2.n34 VDD2.n16 3.49141
R2144 VDD2.n58 VDD2.n57 3.49141
R2145 VDD2.n132 VDD2.n75 2.71565
R2146 VDD2.n104 VDD2.n89 2.71565
R2147 VDD2.n33 VDD2.n18 2.71565
R2148 VDD2.n61 VDD2.n4 2.71565
R2149 VDD2.n133 VDD2.n73 1.93989
R2150 VDD2.n101 VDD2.n100 1.93989
R2151 VDD2.n30 VDD2.n29 1.93989
R2152 VDD2.n62 VDD2.n2 1.93989
R2153 VDD2.n141 VDD2.t0 1.5682
R2154 VDD2.n141 VDD2.t1 1.5682
R2155 VDD2.n69 VDD2.t4 1.5682
R2156 VDD2.n69 VDD2.t3 1.5682
R2157 VDD2.n137 VDD2.n136 1.16414
R2158 VDD2.n97 VDD2.n91 1.16414
R2159 VDD2.n26 VDD2.n20 1.16414
R2160 VDD2.n66 VDD2.n65 1.16414
R2161 VDD2 VDD2.n140 0.976793
R2162 VDD2.n139 VDD2.n71 0.388379
R2163 VDD2.n96 VDD2.n93 0.388379
R2164 VDD2.n25 VDD2.n22 0.388379
R2165 VDD2.n68 VDD2.n0 0.388379
R2166 VDD2.n135 VDD2.n134 0.155672
R2167 VDD2.n134 VDD2.n74 0.155672
R2168 VDD2.n127 VDD2.n74 0.155672
R2169 VDD2.n127 VDD2.n126 0.155672
R2170 VDD2.n126 VDD2.n78 0.155672
R2171 VDD2.n119 VDD2.n78 0.155672
R2172 VDD2.n119 VDD2.n118 0.155672
R2173 VDD2.n118 VDD2.n82 0.155672
R2174 VDD2.n111 VDD2.n82 0.155672
R2175 VDD2.n111 VDD2.n110 0.155672
R2176 VDD2.n110 VDD2.n86 0.155672
R2177 VDD2.n103 VDD2.n86 0.155672
R2178 VDD2.n103 VDD2.n102 0.155672
R2179 VDD2.n102 VDD2.n90 0.155672
R2180 VDD2.n95 VDD2.n90 0.155672
R2181 VDD2.n24 VDD2.n19 0.155672
R2182 VDD2.n31 VDD2.n19 0.155672
R2183 VDD2.n32 VDD2.n31 0.155672
R2184 VDD2.n32 VDD2.n15 0.155672
R2185 VDD2.n39 VDD2.n15 0.155672
R2186 VDD2.n40 VDD2.n39 0.155672
R2187 VDD2.n40 VDD2.n11 0.155672
R2188 VDD2.n47 VDD2.n11 0.155672
R2189 VDD2.n48 VDD2.n47 0.155672
R2190 VDD2.n48 VDD2.n7 0.155672
R2191 VDD2.n55 VDD2.n7 0.155672
R2192 VDD2.n56 VDD2.n55 0.155672
R2193 VDD2.n56 VDD2.n3 0.155672
R2194 VDD2.n63 VDD2.n3 0.155672
R2195 VDD2.n64 VDD2.n63 0.155672
C0 VN VDD1 0.148736f
C1 VDD2 VDD1 0.8543f
C2 VDD2 VN 5.52177f
C3 VTAIL VDD1 8.92772f
C4 VP VDD1 5.699471f
C5 VTAIL VN 5.29491f
C6 VDD2 VTAIL 8.965441f
C7 VN VP 5.57512f
C8 VDD2 VP 0.330679f
C9 VTAIL VP 5.309431f
C10 VDD2 B 4.903556f
C11 VDD1 B 4.956996f
C12 VTAIL B 6.963591f
C13 VN B 8.78387f
C14 VP B 6.997777f
C15 VDD2.n0 B 0.012498f
C16 VDD2.n1 B 0.028214f
C17 VDD2.n2 B 0.012639f
C18 VDD2.n3 B 0.022213f
C19 VDD2.n4 B 0.011936f
C20 VDD2.n5 B 0.028214f
C21 VDD2.n6 B 0.012639f
C22 VDD2.n7 B 0.022213f
C23 VDD2.n8 B 0.011936f
C24 VDD2.n9 B 0.028214f
C25 VDD2.n10 B 0.012639f
C26 VDD2.n11 B 0.022213f
C27 VDD2.n12 B 0.011936f
C28 VDD2.n13 B 0.028214f
C29 VDD2.n14 B 0.012639f
C30 VDD2.n15 B 0.022213f
C31 VDD2.n16 B 0.011936f
C32 VDD2.n17 B 0.028214f
C33 VDD2.n18 B 0.012639f
C34 VDD2.n19 B 0.022213f
C35 VDD2.n20 B 0.011936f
C36 VDD2.n21 B 0.02116f
C37 VDD2.n22 B 0.016667f
C38 VDD2.t2 B 0.04634f
C39 VDD2.n23 B 0.131681f
C40 VDD2.n24 B 1.20396f
C41 VDD2.n25 B 0.011936f
C42 VDD2.n26 B 0.012639f
C43 VDD2.n27 B 0.028214f
C44 VDD2.n28 B 0.028214f
C45 VDD2.n29 B 0.012639f
C46 VDD2.n30 B 0.011936f
C47 VDD2.n31 B 0.022213f
C48 VDD2.n32 B 0.022213f
C49 VDD2.n33 B 0.011936f
C50 VDD2.n34 B 0.012639f
C51 VDD2.n35 B 0.028214f
C52 VDD2.n36 B 0.028214f
C53 VDD2.n37 B 0.012639f
C54 VDD2.n38 B 0.011936f
C55 VDD2.n39 B 0.022213f
C56 VDD2.n40 B 0.022213f
C57 VDD2.n41 B 0.011936f
C58 VDD2.n42 B 0.012639f
C59 VDD2.n43 B 0.028214f
C60 VDD2.n44 B 0.028214f
C61 VDD2.n45 B 0.012639f
C62 VDD2.n46 B 0.011936f
C63 VDD2.n47 B 0.022213f
C64 VDD2.n48 B 0.022213f
C65 VDD2.n49 B 0.011936f
C66 VDD2.n50 B 0.012639f
C67 VDD2.n51 B 0.028214f
C68 VDD2.n52 B 0.028214f
C69 VDD2.n53 B 0.012639f
C70 VDD2.n54 B 0.011936f
C71 VDD2.n55 B 0.022213f
C72 VDD2.n56 B 0.022213f
C73 VDD2.n57 B 0.011936f
C74 VDD2.n58 B 0.012639f
C75 VDD2.n59 B 0.028214f
C76 VDD2.n60 B 0.028214f
C77 VDD2.n61 B 0.012639f
C78 VDD2.n62 B 0.011936f
C79 VDD2.n63 B 0.022213f
C80 VDD2.n64 B 0.055897f
C81 VDD2.n65 B 0.011936f
C82 VDD2.n66 B 0.012639f
C83 VDD2.n67 B 0.056572f
C84 VDD2.n68 B 0.064226f
C85 VDD2.t4 B 0.221703f
C86 VDD2.t3 B 0.221703f
C87 VDD2.n69 B 1.99077f
C88 VDD2.n70 B 1.82727f
C89 VDD2.n71 B 0.012498f
C90 VDD2.n72 B 0.028214f
C91 VDD2.n73 B 0.012639f
C92 VDD2.n74 B 0.022213f
C93 VDD2.n75 B 0.011936f
C94 VDD2.n76 B 0.028214f
C95 VDD2.n77 B 0.012639f
C96 VDD2.n78 B 0.022213f
C97 VDD2.n79 B 0.011936f
C98 VDD2.n80 B 0.028214f
C99 VDD2.n81 B 0.012639f
C100 VDD2.n82 B 0.022213f
C101 VDD2.n83 B 0.011936f
C102 VDD2.n84 B 0.028214f
C103 VDD2.n85 B 0.012639f
C104 VDD2.n86 B 0.022213f
C105 VDD2.n87 B 0.011936f
C106 VDD2.n88 B 0.028214f
C107 VDD2.n89 B 0.012639f
C108 VDD2.n90 B 0.022213f
C109 VDD2.n91 B 0.011936f
C110 VDD2.n92 B 0.02116f
C111 VDD2.n93 B 0.016667f
C112 VDD2.t5 B 0.04634f
C113 VDD2.n94 B 0.131681f
C114 VDD2.n95 B 1.20396f
C115 VDD2.n96 B 0.011936f
C116 VDD2.n97 B 0.012639f
C117 VDD2.n98 B 0.028214f
C118 VDD2.n99 B 0.028214f
C119 VDD2.n100 B 0.012639f
C120 VDD2.n101 B 0.011936f
C121 VDD2.n102 B 0.022213f
C122 VDD2.n103 B 0.022213f
C123 VDD2.n104 B 0.011936f
C124 VDD2.n105 B 0.012639f
C125 VDD2.n106 B 0.028214f
C126 VDD2.n107 B 0.028214f
C127 VDD2.n108 B 0.012639f
C128 VDD2.n109 B 0.011936f
C129 VDD2.n110 B 0.022213f
C130 VDD2.n111 B 0.022213f
C131 VDD2.n112 B 0.011936f
C132 VDD2.n113 B 0.012639f
C133 VDD2.n114 B 0.028214f
C134 VDD2.n115 B 0.028214f
C135 VDD2.n116 B 0.012639f
C136 VDD2.n117 B 0.011936f
C137 VDD2.n118 B 0.022213f
C138 VDD2.n119 B 0.022213f
C139 VDD2.n120 B 0.011936f
C140 VDD2.n121 B 0.012639f
C141 VDD2.n122 B 0.028214f
C142 VDD2.n123 B 0.028214f
C143 VDD2.n124 B 0.012639f
C144 VDD2.n125 B 0.011936f
C145 VDD2.n126 B 0.022213f
C146 VDD2.n127 B 0.022213f
C147 VDD2.n128 B 0.011936f
C148 VDD2.n129 B 0.012639f
C149 VDD2.n130 B 0.028214f
C150 VDD2.n131 B 0.028214f
C151 VDD2.n132 B 0.012639f
C152 VDD2.n133 B 0.011936f
C153 VDD2.n134 B 0.022213f
C154 VDD2.n135 B 0.055897f
C155 VDD2.n136 B 0.011936f
C156 VDD2.n137 B 0.012639f
C157 VDD2.n138 B 0.056572f
C158 VDD2.n139 B 0.062453f
C159 VDD2.n140 B 1.95615f
C160 VDD2.t0 B 0.221703f
C161 VDD2.t1 B 0.221703f
C162 VDD2.n141 B 1.99074f
C163 VN.n0 B 0.211747f
C164 VN.t1 B 1.43301f
C165 VN.t3 B 1.53745f
C166 VN.n1 B 0.574363f
C167 VN.n2 B 0.588096f
C168 VN.n3 B 0.049599f
C169 VN.t2 B 1.49672f
C170 VN.n4 B 0.589994f
C171 VN.n5 B 0.035729f
C172 VN.n6 B 0.211747f
C173 VN.t5 B 1.43301f
C174 VN.t4 B 1.53745f
C175 VN.n7 B 0.574363f
C176 VN.n8 B 0.588096f
C177 VN.n9 B 0.049599f
C178 VN.t0 B 1.49672f
C179 VN.n10 B 0.589994f
C180 VN.n11 B 1.69769f
C181 VDD1.n0 B 0.012514f
C182 VDD1.n1 B 0.028248f
C183 VDD1.n2 B 0.012654f
C184 VDD1.n3 B 0.022241f
C185 VDD1.n4 B 0.011951f
C186 VDD1.n5 B 0.028248f
C187 VDD1.n6 B 0.012654f
C188 VDD1.n7 B 0.022241f
C189 VDD1.n8 B 0.011951f
C190 VDD1.n9 B 0.028248f
C191 VDD1.n10 B 0.012654f
C192 VDD1.n11 B 0.022241f
C193 VDD1.n12 B 0.011951f
C194 VDD1.n13 B 0.028248f
C195 VDD1.n14 B 0.012654f
C196 VDD1.n15 B 0.022241f
C197 VDD1.n16 B 0.011951f
C198 VDD1.n17 B 0.028248f
C199 VDD1.n18 B 0.012654f
C200 VDD1.n19 B 0.022241f
C201 VDD1.n20 B 0.011951f
C202 VDD1.n21 B 0.021186f
C203 VDD1.n22 B 0.016687f
C204 VDD1.t3 B 0.046397f
C205 VDD1.n23 B 0.131843f
C206 VDD1.n24 B 1.20544f
C207 VDD1.n25 B 0.011951f
C208 VDD1.n26 B 0.012654f
C209 VDD1.n27 B 0.028248f
C210 VDD1.n28 B 0.028248f
C211 VDD1.n29 B 0.012654f
C212 VDD1.n30 B 0.011951f
C213 VDD1.n31 B 0.022241f
C214 VDD1.n32 B 0.022241f
C215 VDD1.n33 B 0.011951f
C216 VDD1.n34 B 0.012654f
C217 VDD1.n35 B 0.028248f
C218 VDD1.n36 B 0.028248f
C219 VDD1.n37 B 0.012654f
C220 VDD1.n38 B 0.011951f
C221 VDD1.n39 B 0.022241f
C222 VDD1.n40 B 0.022241f
C223 VDD1.n41 B 0.011951f
C224 VDD1.n42 B 0.012654f
C225 VDD1.n43 B 0.028248f
C226 VDD1.n44 B 0.028248f
C227 VDD1.n45 B 0.012654f
C228 VDD1.n46 B 0.011951f
C229 VDD1.n47 B 0.022241f
C230 VDD1.n48 B 0.022241f
C231 VDD1.n49 B 0.011951f
C232 VDD1.n50 B 0.012654f
C233 VDD1.n51 B 0.028248f
C234 VDD1.n52 B 0.028248f
C235 VDD1.n53 B 0.012654f
C236 VDD1.n54 B 0.011951f
C237 VDD1.n55 B 0.022241f
C238 VDD1.n56 B 0.022241f
C239 VDD1.n57 B 0.011951f
C240 VDD1.n58 B 0.012654f
C241 VDD1.n59 B 0.028248f
C242 VDD1.n60 B 0.028248f
C243 VDD1.n61 B 0.012654f
C244 VDD1.n62 B 0.011951f
C245 VDD1.n63 B 0.022241f
C246 VDD1.n64 B 0.055966f
C247 VDD1.n65 B 0.011951f
C248 VDD1.n66 B 0.012654f
C249 VDD1.n67 B 0.056642f
C250 VDD1.n68 B 0.064675f
C251 VDD1.n69 B 0.012514f
C252 VDD1.n70 B 0.028248f
C253 VDD1.n71 B 0.012654f
C254 VDD1.n72 B 0.022241f
C255 VDD1.n73 B 0.011951f
C256 VDD1.n74 B 0.028248f
C257 VDD1.n75 B 0.012654f
C258 VDD1.n76 B 0.022241f
C259 VDD1.n77 B 0.011951f
C260 VDD1.n78 B 0.028248f
C261 VDD1.n79 B 0.012654f
C262 VDD1.n80 B 0.022241f
C263 VDD1.n81 B 0.011951f
C264 VDD1.n82 B 0.028248f
C265 VDD1.n83 B 0.012654f
C266 VDD1.n84 B 0.022241f
C267 VDD1.n85 B 0.011951f
C268 VDD1.n86 B 0.028248f
C269 VDD1.n87 B 0.012654f
C270 VDD1.n88 B 0.022241f
C271 VDD1.n89 B 0.011951f
C272 VDD1.n90 B 0.021186f
C273 VDD1.n91 B 0.016687f
C274 VDD1.t0 B 0.046397f
C275 VDD1.n92 B 0.131843f
C276 VDD1.n93 B 1.20544f
C277 VDD1.n94 B 0.011951f
C278 VDD1.n95 B 0.012654f
C279 VDD1.n96 B 0.028248f
C280 VDD1.n97 B 0.028248f
C281 VDD1.n98 B 0.012654f
C282 VDD1.n99 B 0.011951f
C283 VDD1.n100 B 0.022241f
C284 VDD1.n101 B 0.022241f
C285 VDD1.n102 B 0.011951f
C286 VDD1.n103 B 0.012654f
C287 VDD1.n104 B 0.028248f
C288 VDD1.n105 B 0.028248f
C289 VDD1.n106 B 0.012654f
C290 VDD1.n107 B 0.011951f
C291 VDD1.n108 B 0.022241f
C292 VDD1.n109 B 0.022241f
C293 VDD1.n110 B 0.011951f
C294 VDD1.n111 B 0.012654f
C295 VDD1.n112 B 0.028248f
C296 VDD1.n113 B 0.028248f
C297 VDD1.n114 B 0.012654f
C298 VDD1.n115 B 0.011951f
C299 VDD1.n116 B 0.022241f
C300 VDD1.n117 B 0.022241f
C301 VDD1.n118 B 0.011951f
C302 VDD1.n119 B 0.012654f
C303 VDD1.n120 B 0.028248f
C304 VDD1.n121 B 0.028248f
C305 VDD1.n122 B 0.012654f
C306 VDD1.n123 B 0.011951f
C307 VDD1.n124 B 0.022241f
C308 VDD1.n125 B 0.022241f
C309 VDD1.n126 B 0.011951f
C310 VDD1.n127 B 0.012654f
C311 VDD1.n128 B 0.028248f
C312 VDD1.n129 B 0.028248f
C313 VDD1.n130 B 0.012654f
C314 VDD1.n131 B 0.011951f
C315 VDD1.n132 B 0.022241f
C316 VDD1.n133 B 0.055966f
C317 VDD1.n134 B 0.011951f
C318 VDD1.n135 B 0.012654f
C319 VDD1.n136 B 0.056642f
C320 VDD1.n137 B 0.064305f
C321 VDD1.t4 B 0.221976f
C322 VDD1.t5 B 0.221976f
C323 VDD1.n138 B 1.99322f
C324 VDD1.n139 B 1.90655f
C325 VDD1.t2 B 0.221976f
C326 VDD1.t1 B 0.221976f
C327 VDD1.n140 B 1.99207f
C328 VDD1.n141 B 2.13973f
C329 VTAIL.t11 B 0.232814f
C330 VTAIL.t0 B 0.232814f
C331 VTAIL.n0 B 2.02576f
C332 VTAIL.n1 B 0.325846f
C333 VTAIL.n2 B 0.013125f
C334 VTAIL.n3 B 0.029628f
C335 VTAIL.n4 B 0.013272f
C336 VTAIL.n5 B 0.023327f
C337 VTAIL.n6 B 0.012535f
C338 VTAIL.n7 B 0.029628f
C339 VTAIL.n8 B 0.013272f
C340 VTAIL.n9 B 0.023327f
C341 VTAIL.n10 B 0.012535f
C342 VTAIL.n11 B 0.029628f
C343 VTAIL.n12 B 0.013272f
C344 VTAIL.n13 B 0.023327f
C345 VTAIL.n14 B 0.012535f
C346 VTAIL.n15 B 0.029628f
C347 VTAIL.n16 B 0.013272f
C348 VTAIL.n17 B 0.023327f
C349 VTAIL.n18 B 0.012535f
C350 VTAIL.n19 B 0.029628f
C351 VTAIL.n20 B 0.013272f
C352 VTAIL.n21 B 0.023327f
C353 VTAIL.n22 B 0.012535f
C354 VTAIL.n23 B 0.022221f
C355 VTAIL.n24 B 0.017502f
C356 VTAIL.t9 B 0.048663f
C357 VTAIL.n25 B 0.138281f
C358 VTAIL.n26 B 1.2643f
C359 VTAIL.n27 B 0.012535f
C360 VTAIL.n28 B 0.013272f
C361 VTAIL.n29 B 0.029628f
C362 VTAIL.n30 B 0.029628f
C363 VTAIL.n31 B 0.013272f
C364 VTAIL.n32 B 0.012535f
C365 VTAIL.n33 B 0.023327f
C366 VTAIL.n34 B 0.023327f
C367 VTAIL.n35 B 0.012535f
C368 VTAIL.n36 B 0.013272f
C369 VTAIL.n37 B 0.029628f
C370 VTAIL.n38 B 0.029628f
C371 VTAIL.n39 B 0.013272f
C372 VTAIL.n40 B 0.012535f
C373 VTAIL.n41 B 0.023327f
C374 VTAIL.n42 B 0.023327f
C375 VTAIL.n43 B 0.012535f
C376 VTAIL.n44 B 0.013272f
C377 VTAIL.n45 B 0.029628f
C378 VTAIL.n46 B 0.029628f
C379 VTAIL.n47 B 0.013272f
C380 VTAIL.n48 B 0.012535f
C381 VTAIL.n49 B 0.023327f
C382 VTAIL.n50 B 0.023327f
C383 VTAIL.n51 B 0.012535f
C384 VTAIL.n52 B 0.013272f
C385 VTAIL.n53 B 0.029628f
C386 VTAIL.n54 B 0.029628f
C387 VTAIL.n55 B 0.013272f
C388 VTAIL.n56 B 0.012535f
C389 VTAIL.n57 B 0.023327f
C390 VTAIL.n58 B 0.023327f
C391 VTAIL.n59 B 0.012535f
C392 VTAIL.n60 B 0.013272f
C393 VTAIL.n61 B 0.029628f
C394 VTAIL.n62 B 0.029628f
C395 VTAIL.n63 B 0.013272f
C396 VTAIL.n64 B 0.012535f
C397 VTAIL.n65 B 0.023327f
C398 VTAIL.n66 B 0.058698f
C399 VTAIL.n67 B 0.012535f
C400 VTAIL.n68 B 0.013272f
C401 VTAIL.n69 B 0.059407f
C402 VTAIL.n70 B 0.049507f
C403 VTAIL.n71 B 0.195595f
C404 VTAIL.t5 B 0.232814f
C405 VTAIL.t8 B 0.232814f
C406 VTAIL.n72 B 2.02576f
C407 VTAIL.n73 B 1.62842f
C408 VTAIL.t1 B 0.232814f
C409 VTAIL.t3 B 0.232814f
C410 VTAIL.n74 B 2.02576f
C411 VTAIL.n75 B 1.62843f
C412 VTAIL.n76 B 0.013125f
C413 VTAIL.n77 B 0.029628f
C414 VTAIL.n78 B 0.013272f
C415 VTAIL.n79 B 0.023327f
C416 VTAIL.n80 B 0.012535f
C417 VTAIL.n81 B 0.029628f
C418 VTAIL.n82 B 0.013272f
C419 VTAIL.n83 B 0.023327f
C420 VTAIL.n84 B 0.012535f
C421 VTAIL.n85 B 0.029628f
C422 VTAIL.n86 B 0.013272f
C423 VTAIL.n87 B 0.023327f
C424 VTAIL.n88 B 0.012535f
C425 VTAIL.n89 B 0.029628f
C426 VTAIL.n90 B 0.013272f
C427 VTAIL.n91 B 0.023327f
C428 VTAIL.n92 B 0.012535f
C429 VTAIL.n93 B 0.029628f
C430 VTAIL.n94 B 0.013272f
C431 VTAIL.n95 B 0.023327f
C432 VTAIL.n96 B 0.012535f
C433 VTAIL.n97 B 0.022221f
C434 VTAIL.n98 B 0.017502f
C435 VTAIL.t4 B 0.048663f
C436 VTAIL.n99 B 0.138281f
C437 VTAIL.n100 B 1.2643f
C438 VTAIL.n101 B 0.012535f
C439 VTAIL.n102 B 0.013272f
C440 VTAIL.n103 B 0.029628f
C441 VTAIL.n104 B 0.029628f
C442 VTAIL.n105 B 0.013272f
C443 VTAIL.n106 B 0.012535f
C444 VTAIL.n107 B 0.023327f
C445 VTAIL.n108 B 0.023327f
C446 VTAIL.n109 B 0.012535f
C447 VTAIL.n110 B 0.013272f
C448 VTAIL.n111 B 0.029628f
C449 VTAIL.n112 B 0.029628f
C450 VTAIL.n113 B 0.013272f
C451 VTAIL.n114 B 0.012535f
C452 VTAIL.n115 B 0.023327f
C453 VTAIL.n116 B 0.023327f
C454 VTAIL.n117 B 0.012535f
C455 VTAIL.n118 B 0.013272f
C456 VTAIL.n119 B 0.029628f
C457 VTAIL.n120 B 0.029628f
C458 VTAIL.n121 B 0.013272f
C459 VTAIL.n122 B 0.012535f
C460 VTAIL.n123 B 0.023327f
C461 VTAIL.n124 B 0.023327f
C462 VTAIL.n125 B 0.012535f
C463 VTAIL.n126 B 0.013272f
C464 VTAIL.n127 B 0.029628f
C465 VTAIL.n128 B 0.029628f
C466 VTAIL.n129 B 0.013272f
C467 VTAIL.n130 B 0.012535f
C468 VTAIL.n131 B 0.023327f
C469 VTAIL.n132 B 0.023327f
C470 VTAIL.n133 B 0.012535f
C471 VTAIL.n134 B 0.013272f
C472 VTAIL.n135 B 0.029628f
C473 VTAIL.n136 B 0.029628f
C474 VTAIL.n137 B 0.013272f
C475 VTAIL.n138 B 0.012535f
C476 VTAIL.n139 B 0.023327f
C477 VTAIL.n140 B 0.058698f
C478 VTAIL.n141 B 0.012535f
C479 VTAIL.n142 B 0.013272f
C480 VTAIL.n143 B 0.059407f
C481 VTAIL.n144 B 0.049507f
C482 VTAIL.n145 B 0.195595f
C483 VTAIL.t6 B 0.232814f
C484 VTAIL.t10 B 0.232814f
C485 VTAIL.n146 B 2.02576f
C486 VTAIL.n147 B 0.390486f
C487 VTAIL.n148 B 0.013125f
C488 VTAIL.n149 B 0.029628f
C489 VTAIL.n150 B 0.013272f
C490 VTAIL.n151 B 0.023327f
C491 VTAIL.n152 B 0.012535f
C492 VTAIL.n153 B 0.029628f
C493 VTAIL.n154 B 0.013272f
C494 VTAIL.n155 B 0.023327f
C495 VTAIL.n156 B 0.012535f
C496 VTAIL.n157 B 0.029628f
C497 VTAIL.n158 B 0.013272f
C498 VTAIL.n159 B 0.023327f
C499 VTAIL.n160 B 0.012535f
C500 VTAIL.n161 B 0.029628f
C501 VTAIL.n162 B 0.013272f
C502 VTAIL.n163 B 0.023327f
C503 VTAIL.n164 B 0.012535f
C504 VTAIL.n165 B 0.029628f
C505 VTAIL.n166 B 0.013272f
C506 VTAIL.n167 B 0.023327f
C507 VTAIL.n168 B 0.012535f
C508 VTAIL.n169 B 0.022221f
C509 VTAIL.n170 B 0.017502f
C510 VTAIL.t7 B 0.048663f
C511 VTAIL.n171 B 0.138281f
C512 VTAIL.n172 B 1.2643f
C513 VTAIL.n173 B 0.012535f
C514 VTAIL.n174 B 0.013272f
C515 VTAIL.n175 B 0.029628f
C516 VTAIL.n176 B 0.029628f
C517 VTAIL.n177 B 0.013272f
C518 VTAIL.n178 B 0.012535f
C519 VTAIL.n179 B 0.023327f
C520 VTAIL.n180 B 0.023327f
C521 VTAIL.n181 B 0.012535f
C522 VTAIL.n182 B 0.013272f
C523 VTAIL.n183 B 0.029628f
C524 VTAIL.n184 B 0.029628f
C525 VTAIL.n185 B 0.013272f
C526 VTAIL.n186 B 0.012535f
C527 VTAIL.n187 B 0.023327f
C528 VTAIL.n188 B 0.023327f
C529 VTAIL.n189 B 0.012535f
C530 VTAIL.n190 B 0.013272f
C531 VTAIL.n191 B 0.029628f
C532 VTAIL.n192 B 0.029628f
C533 VTAIL.n193 B 0.013272f
C534 VTAIL.n194 B 0.012535f
C535 VTAIL.n195 B 0.023327f
C536 VTAIL.n196 B 0.023327f
C537 VTAIL.n197 B 0.012535f
C538 VTAIL.n198 B 0.013272f
C539 VTAIL.n199 B 0.029628f
C540 VTAIL.n200 B 0.029628f
C541 VTAIL.n201 B 0.013272f
C542 VTAIL.n202 B 0.012535f
C543 VTAIL.n203 B 0.023327f
C544 VTAIL.n204 B 0.023327f
C545 VTAIL.n205 B 0.012535f
C546 VTAIL.n206 B 0.013272f
C547 VTAIL.n207 B 0.029628f
C548 VTAIL.n208 B 0.029628f
C549 VTAIL.n209 B 0.013272f
C550 VTAIL.n210 B 0.012535f
C551 VTAIL.n211 B 0.023327f
C552 VTAIL.n212 B 0.058698f
C553 VTAIL.n213 B 0.012535f
C554 VTAIL.n214 B 0.013272f
C555 VTAIL.n215 B 0.059407f
C556 VTAIL.n216 B 0.049507f
C557 VTAIL.n217 B 1.34153f
C558 VTAIL.n218 B 0.013125f
C559 VTAIL.n219 B 0.029628f
C560 VTAIL.n220 B 0.013272f
C561 VTAIL.n221 B 0.023327f
C562 VTAIL.n222 B 0.012535f
C563 VTAIL.n223 B 0.029628f
C564 VTAIL.n224 B 0.013272f
C565 VTAIL.n225 B 0.023327f
C566 VTAIL.n226 B 0.012535f
C567 VTAIL.n227 B 0.029628f
C568 VTAIL.n228 B 0.013272f
C569 VTAIL.n229 B 0.023327f
C570 VTAIL.n230 B 0.012535f
C571 VTAIL.n231 B 0.029628f
C572 VTAIL.n232 B 0.013272f
C573 VTAIL.n233 B 0.023327f
C574 VTAIL.n234 B 0.012535f
C575 VTAIL.n235 B 0.029628f
C576 VTAIL.n236 B 0.013272f
C577 VTAIL.n237 B 0.023327f
C578 VTAIL.n238 B 0.012535f
C579 VTAIL.n239 B 0.022221f
C580 VTAIL.n240 B 0.017502f
C581 VTAIL.t2 B 0.048663f
C582 VTAIL.n241 B 0.138281f
C583 VTAIL.n242 B 1.2643f
C584 VTAIL.n243 B 0.012535f
C585 VTAIL.n244 B 0.013272f
C586 VTAIL.n245 B 0.029628f
C587 VTAIL.n246 B 0.029628f
C588 VTAIL.n247 B 0.013272f
C589 VTAIL.n248 B 0.012535f
C590 VTAIL.n249 B 0.023327f
C591 VTAIL.n250 B 0.023327f
C592 VTAIL.n251 B 0.012535f
C593 VTAIL.n252 B 0.013272f
C594 VTAIL.n253 B 0.029628f
C595 VTAIL.n254 B 0.029628f
C596 VTAIL.n255 B 0.013272f
C597 VTAIL.n256 B 0.012535f
C598 VTAIL.n257 B 0.023327f
C599 VTAIL.n258 B 0.023327f
C600 VTAIL.n259 B 0.012535f
C601 VTAIL.n260 B 0.013272f
C602 VTAIL.n261 B 0.029628f
C603 VTAIL.n262 B 0.029628f
C604 VTAIL.n263 B 0.013272f
C605 VTAIL.n264 B 0.012535f
C606 VTAIL.n265 B 0.023327f
C607 VTAIL.n266 B 0.023327f
C608 VTAIL.n267 B 0.012535f
C609 VTAIL.n268 B 0.013272f
C610 VTAIL.n269 B 0.029628f
C611 VTAIL.n270 B 0.029628f
C612 VTAIL.n271 B 0.013272f
C613 VTAIL.n272 B 0.012535f
C614 VTAIL.n273 B 0.023327f
C615 VTAIL.n274 B 0.023327f
C616 VTAIL.n275 B 0.012535f
C617 VTAIL.n276 B 0.013272f
C618 VTAIL.n277 B 0.029628f
C619 VTAIL.n278 B 0.029628f
C620 VTAIL.n279 B 0.013272f
C621 VTAIL.n280 B 0.012535f
C622 VTAIL.n281 B 0.023327f
C623 VTAIL.n282 B 0.058698f
C624 VTAIL.n283 B 0.012535f
C625 VTAIL.n284 B 0.013272f
C626 VTAIL.n285 B 0.059407f
C627 VTAIL.n286 B 0.049507f
C628 VTAIL.n287 B 1.31415f
C629 VP.n0 B 0.051696f
C630 VP.t1 B 1.45525f
C631 VP.n1 B 0.050368f
C632 VP.n2 B 0.215032f
C633 VP.t4 B 1.51994f
C634 VP.t3 B 1.45525f
C635 VP.t2 B 1.5613f
C636 VP.n3 B 0.583275f
C637 VP.n4 B 0.597221f
C638 VP.n5 B 0.050368f
C639 VP.n6 B 0.599148f
C640 VP.n7 B 1.70242f
C641 VP.t5 B 1.51994f
C642 VP.n8 B 0.599148f
C643 VP.n9 B 1.7345f
C644 VP.n10 B 0.051696f
C645 VP.n11 B 0.038742f
C646 VP.n12 B 0.570437f
C647 VP.n13 B 0.050368f
C648 VP.t0 B 1.51994f
C649 VP.n14 B 0.599148f
C650 VP.n15 B 0.036283f
.ends

