* NGSPICE file created from diff_pair_sample_1201.ext - technology: sky130A

.subckt diff_pair_sample_1201 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=2.8353 pd=15.32 as=0 ps=0 w=7.27 l=2.97
X1 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=2.8353 pd=15.32 as=0 ps=0 w=7.27 l=2.97
X2 VTAIL.t10 VP.t0 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.19955 pd=7.6 as=1.19955 ps=7.6 w=7.27 l=2.97
X3 VTAIL.t9 VP.t1 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.19955 pd=7.6 as=1.19955 ps=7.6 w=7.27 l=2.97
X4 VDD2.t5 VN.t0 VTAIL.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=2.8353 pd=15.32 as=1.19955 ps=7.6 w=7.27 l=2.97
X5 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.8353 pd=15.32 as=0 ps=0 w=7.27 l=2.97
X6 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.8353 pd=15.32 as=0 ps=0 w=7.27 l=2.97
X7 VTAIL.t3 VN.t1 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=1.19955 pd=7.6 as=1.19955 ps=7.6 w=7.27 l=2.97
X8 VTAIL.t1 VN.t2 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.19955 pd=7.6 as=1.19955 ps=7.6 w=7.27 l=2.97
X9 VDD2.t2 VN.t3 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=2.8353 pd=15.32 as=1.19955 ps=7.6 w=7.27 l=2.97
X10 VDD2.t1 VN.t4 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.19955 pd=7.6 as=2.8353 ps=15.32 w=7.27 l=2.97
X11 VDD1.t5 VP.t2 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=2.8353 pd=15.32 as=1.19955 ps=7.6 w=7.27 l=2.97
X12 VDD2.t0 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.19955 pd=7.6 as=2.8353 ps=15.32 w=7.27 l=2.97
X13 VDD1.t0 VP.t3 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.19955 pd=7.6 as=2.8353 ps=15.32 w=7.27 l=2.97
X14 VDD1.t4 VP.t4 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.8353 pd=15.32 as=1.19955 ps=7.6 w=7.27 l=2.97
X15 VDD1.t2 VP.t5 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.19955 pd=7.6 as=2.8353 ps=15.32 w=7.27 l=2.97
R0 B.n712 B.n711 585
R1 B.n713 B.n712 585
R2 B.n250 B.n120 585
R3 B.n249 B.n248 585
R4 B.n247 B.n246 585
R5 B.n245 B.n244 585
R6 B.n243 B.n242 585
R7 B.n241 B.n240 585
R8 B.n239 B.n238 585
R9 B.n237 B.n236 585
R10 B.n235 B.n234 585
R11 B.n233 B.n232 585
R12 B.n231 B.n230 585
R13 B.n229 B.n228 585
R14 B.n227 B.n226 585
R15 B.n225 B.n224 585
R16 B.n223 B.n222 585
R17 B.n221 B.n220 585
R18 B.n219 B.n218 585
R19 B.n217 B.n216 585
R20 B.n215 B.n214 585
R21 B.n213 B.n212 585
R22 B.n211 B.n210 585
R23 B.n209 B.n208 585
R24 B.n207 B.n206 585
R25 B.n205 B.n204 585
R26 B.n203 B.n202 585
R27 B.n201 B.n200 585
R28 B.n199 B.n198 585
R29 B.n196 B.n195 585
R30 B.n194 B.n193 585
R31 B.n192 B.n191 585
R32 B.n190 B.n189 585
R33 B.n188 B.n187 585
R34 B.n186 B.n185 585
R35 B.n184 B.n183 585
R36 B.n182 B.n181 585
R37 B.n180 B.n179 585
R38 B.n178 B.n177 585
R39 B.n176 B.n175 585
R40 B.n174 B.n173 585
R41 B.n172 B.n171 585
R42 B.n170 B.n169 585
R43 B.n168 B.n167 585
R44 B.n166 B.n165 585
R45 B.n164 B.n163 585
R46 B.n162 B.n161 585
R47 B.n160 B.n159 585
R48 B.n158 B.n157 585
R49 B.n156 B.n155 585
R50 B.n154 B.n153 585
R51 B.n152 B.n151 585
R52 B.n150 B.n149 585
R53 B.n148 B.n147 585
R54 B.n146 B.n145 585
R55 B.n144 B.n143 585
R56 B.n142 B.n141 585
R57 B.n140 B.n139 585
R58 B.n138 B.n137 585
R59 B.n136 B.n135 585
R60 B.n134 B.n133 585
R61 B.n132 B.n131 585
R62 B.n130 B.n129 585
R63 B.n128 B.n127 585
R64 B.n88 B.n87 585
R65 B.n716 B.n715 585
R66 B.n710 B.n121 585
R67 B.n121 B.n85 585
R68 B.n709 B.n84 585
R69 B.n720 B.n84 585
R70 B.n708 B.n83 585
R71 B.n721 B.n83 585
R72 B.n707 B.n82 585
R73 B.n722 B.n82 585
R74 B.n706 B.n705 585
R75 B.n705 B.n78 585
R76 B.n704 B.n77 585
R77 B.n728 B.n77 585
R78 B.n703 B.n76 585
R79 B.n729 B.n76 585
R80 B.n702 B.n75 585
R81 B.n730 B.n75 585
R82 B.n701 B.n700 585
R83 B.n700 B.n74 585
R84 B.n699 B.n70 585
R85 B.n736 B.n70 585
R86 B.n698 B.n69 585
R87 B.n737 B.n69 585
R88 B.n697 B.n68 585
R89 B.n738 B.n68 585
R90 B.n696 B.n695 585
R91 B.n695 B.n64 585
R92 B.n694 B.n63 585
R93 B.n744 B.n63 585
R94 B.n693 B.n62 585
R95 B.n745 B.n62 585
R96 B.n692 B.n61 585
R97 B.n746 B.n61 585
R98 B.n691 B.n690 585
R99 B.n690 B.n57 585
R100 B.n689 B.n56 585
R101 B.n752 B.n56 585
R102 B.n688 B.n55 585
R103 B.n753 B.n55 585
R104 B.n687 B.n54 585
R105 B.n754 B.n54 585
R106 B.n686 B.n685 585
R107 B.n685 B.n50 585
R108 B.n684 B.n49 585
R109 B.n760 B.n49 585
R110 B.n683 B.n48 585
R111 B.n761 B.n48 585
R112 B.n682 B.n47 585
R113 B.n762 B.n47 585
R114 B.n681 B.n680 585
R115 B.n680 B.n43 585
R116 B.n679 B.n42 585
R117 B.n768 B.n42 585
R118 B.n678 B.n41 585
R119 B.n769 B.n41 585
R120 B.n677 B.n40 585
R121 B.n770 B.n40 585
R122 B.n676 B.n675 585
R123 B.n675 B.n36 585
R124 B.n674 B.n35 585
R125 B.n776 B.n35 585
R126 B.n673 B.n34 585
R127 B.n777 B.n34 585
R128 B.n672 B.n33 585
R129 B.n778 B.n33 585
R130 B.n671 B.n670 585
R131 B.n670 B.n29 585
R132 B.n669 B.n28 585
R133 B.n784 B.n28 585
R134 B.n668 B.n27 585
R135 B.n785 B.n27 585
R136 B.n667 B.n26 585
R137 B.n786 B.n26 585
R138 B.n666 B.n665 585
R139 B.n665 B.n22 585
R140 B.n664 B.n21 585
R141 B.n792 B.n21 585
R142 B.n663 B.n20 585
R143 B.n793 B.n20 585
R144 B.n662 B.n19 585
R145 B.n794 B.n19 585
R146 B.n661 B.n660 585
R147 B.n660 B.n18 585
R148 B.n659 B.n14 585
R149 B.n800 B.n14 585
R150 B.n658 B.n13 585
R151 B.n801 B.n13 585
R152 B.n657 B.n12 585
R153 B.n802 B.n12 585
R154 B.n656 B.n655 585
R155 B.n655 B.n8 585
R156 B.n654 B.n7 585
R157 B.n808 B.n7 585
R158 B.n653 B.n6 585
R159 B.n809 B.n6 585
R160 B.n652 B.n5 585
R161 B.n810 B.n5 585
R162 B.n651 B.n650 585
R163 B.n650 B.n4 585
R164 B.n649 B.n251 585
R165 B.n649 B.n648 585
R166 B.n639 B.n252 585
R167 B.n253 B.n252 585
R168 B.n641 B.n640 585
R169 B.n642 B.n641 585
R170 B.n638 B.n258 585
R171 B.n258 B.n257 585
R172 B.n637 B.n636 585
R173 B.n636 B.n635 585
R174 B.n260 B.n259 585
R175 B.n628 B.n260 585
R176 B.n627 B.n626 585
R177 B.n629 B.n627 585
R178 B.n625 B.n265 585
R179 B.n265 B.n264 585
R180 B.n624 B.n623 585
R181 B.n623 B.n622 585
R182 B.n267 B.n266 585
R183 B.n268 B.n267 585
R184 B.n615 B.n614 585
R185 B.n616 B.n615 585
R186 B.n613 B.n273 585
R187 B.n273 B.n272 585
R188 B.n612 B.n611 585
R189 B.n611 B.n610 585
R190 B.n275 B.n274 585
R191 B.n276 B.n275 585
R192 B.n603 B.n602 585
R193 B.n604 B.n603 585
R194 B.n601 B.n280 585
R195 B.n284 B.n280 585
R196 B.n600 B.n599 585
R197 B.n599 B.n598 585
R198 B.n282 B.n281 585
R199 B.n283 B.n282 585
R200 B.n591 B.n590 585
R201 B.n592 B.n591 585
R202 B.n589 B.n289 585
R203 B.n289 B.n288 585
R204 B.n588 B.n587 585
R205 B.n587 B.n586 585
R206 B.n291 B.n290 585
R207 B.n292 B.n291 585
R208 B.n579 B.n578 585
R209 B.n580 B.n579 585
R210 B.n577 B.n297 585
R211 B.n297 B.n296 585
R212 B.n576 B.n575 585
R213 B.n575 B.n574 585
R214 B.n299 B.n298 585
R215 B.n300 B.n299 585
R216 B.n567 B.n566 585
R217 B.n568 B.n567 585
R218 B.n565 B.n305 585
R219 B.n305 B.n304 585
R220 B.n564 B.n563 585
R221 B.n563 B.n562 585
R222 B.n307 B.n306 585
R223 B.n308 B.n307 585
R224 B.n555 B.n554 585
R225 B.n556 B.n555 585
R226 B.n553 B.n313 585
R227 B.n313 B.n312 585
R228 B.n552 B.n551 585
R229 B.n551 B.n550 585
R230 B.n315 B.n314 585
R231 B.n316 B.n315 585
R232 B.n543 B.n542 585
R233 B.n544 B.n543 585
R234 B.n541 B.n321 585
R235 B.n321 B.n320 585
R236 B.n540 B.n539 585
R237 B.n539 B.n538 585
R238 B.n323 B.n322 585
R239 B.n531 B.n323 585
R240 B.n530 B.n529 585
R241 B.n532 B.n530 585
R242 B.n528 B.n328 585
R243 B.n328 B.n327 585
R244 B.n527 B.n526 585
R245 B.n526 B.n525 585
R246 B.n330 B.n329 585
R247 B.n331 B.n330 585
R248 B.n518 B.n517 585
R249 B.n519 B.n518 585
R250 B.n516 B.n336 585
R251 B.n336 B.n335 585
R252 B.n515 B.n514 585
R253 B.n514 B.n513 585
R254 B.n338 B.n337 585
R255 B.n339 B.n338 585
R256 B.n509 B.n508 585
R257 B.n342 B.n341 585
R258 B.n505 B.n504 585
R259 B.n506 B.n505 585
R260 B.n503 B.n374 585
R261 B.n502 B.n501 585
R262 B.n500 B.n499 585
R263 B.n498 B.n497 585
R264 B.n496 B.n495 585
R265 B.n494 B.n493 585
R266 B.n492 B.n491 585
R267 B.n490 B.n489 585
R268 B.n488 B.n487 585
R269 B.n486 B.n485 585
R270 B.n484 B.n483 585
R271 B.n482 B.n481 585
R272 B.n480 B.n479 585
R273 B.n478 B.n477 585
R274 B.n476 B.n475 585
R275 B.n474 B.n473 585
R276 B.n472 B.n471 585
R277 B.n470 B.n469 585
R278 B.n468 B.n467 585
R279 B.n466 B.n465 585
R280 B.n464 B.n463 585
R281 B.n462 B.n461 585
R282 B.n460 B.n459 585
R283 B.n458 B.n457 585
R284 B.n456 B.n455 585
R285 B.n453 B.n452 585
R286 B.n451 B.n450 585
R287 B.n449 B.n448 585
R288 B.n447 B.n446 585
R289 B.n445 B.n444 585
R290 B.n443 B.n442 585
R291 B.n441 B.n440 585
R292 B.n439 B.n438 585
R293 B.n437 B.n436 585
R294 B.n435 B.n434 585
R295 B.n433 B.n432 585
R296 B.n431 B.n430 585
R297 B.n429 B.n428 585
R298 B.n427 B.n426 585
R299 B.n425 B.n424 585
R300 B.n423 B.n422 585
R301 B.n421 B.n420 585
R302 B.n419 B.n418 585
R303 B.n417 B.n416 585
R304 B.n415 B.n414 585
R305 B.n413 B.n412 585
R306 B.n411 B.n410 585
R307 B.n409 B.n408 585
R308 B.n407 B.n406 585
R309 B.n405 B.n404 585
R310 B.n403 B.n402 585
R311 B.n401 B.n400 585
R312 B.n399 B.n398 585
R313 B.n397 B.n396 585
R314 B.n395 B.n394 585
R315 B.n393 B.n392 585
R316 B.n391 B.n390 585
R317 B.n389 B.n388 585
R318 B.n387 B.n386 585
R319 B.n385 B.n384 585
R320 B.n383 B.n382 585
R321 B.n381 B.n380 585
R322 B.n510 B.n340 585
R323 B.n340 B.n339 585
R324 B.n512 B.n511 585
R325 B.n513 B.n512 585
R326 B.n334 B.n333 585
R327 B.n335 B.n334 585
R328 B.n521 B.n520 585
R329 B.n520 B.n519 585
R330 B.n522 B.n332 585
R331 B.n332 B.n331 585
R332 B.n524 B.n523 585
R333 B.n525 B.n524 585
R334 B.n326 B.n325 585
R335 B.n327 B.n326 585
R336 B.n534 B.n533 585
R337 B.n533 B.n532 585
R338 B.n535 B.n324 585
R339 B.n531 B.n324 585
R340 B.n537 B.n536 585
R341 B.n538 B.n537 585
R342 B.n319 B.n318 585
R343 B.n320 B.n319 585
R344 B.n546 B.n545 585
R345 B.n545 B.n544 585
R346 B.n547 B.n317 585
R347 B.n317 B.n316 585
R348 B.n549 B.n548 585
R349 B.n550 B.n549 585
R350 B.n311 B.n310 585
R351 B.n312 B.n311 585
R352 B.n558 B.n557 585
R353 B.n557 B.n556 585
R354 B.n559 B.n309 585
R355 B.n309 B.n308 585
R356 B.n561 B.n560 585
R357 B.n562 B.n561 585
R358 B.n303 B.n302 585
R359 B.n304 B.n303 585
R360 B.n570 B.n569 585
R361 B.n569 B.n568 585
R362 B.n571 B.n301 585
R363 B.n301 B.n300 585
R364 B.n573 B.n572 585
R365 B.n574 B.n573 585
R366 B.n295 B.n294 585
R367 B.n296 B.n295 585
R368 B.n582 B.n581 585
R369 B.n581 B.n580 585
R370 B.n583 B.n293 585
R371 B.n293 B.n292 585
R372 B.n585 B.n584 585
R373 B.n586 B.n585 585
R374 B.n287 B.n286 585
R375 B.n288 B.n287 585
R376 B.n594 B.n593 585
R377 B.n593 B.n592 585
R378 B.n595 B.n285 585
R379 B.n285 B.n283 585
R380 B.n597 B.n596 585
R381 B.n598 B.n597 585
R382 B.n279 B.n278 585
R383 B.n284 B.n279 585
R384 B.n606 B.n605 585
R385 B.n605 B.n604 585
R386 B.n607 B.n277 585
R387 B.n277 B.n276 585
R388 B.n609 B.n608 585
R389 B.n610 B.n609 585
R390 B.n271 B.n270 585
R391 B.n272 B.n271 585
R392 B.n618 B.n617 585
R393 B.n617 B.n616 585
R394 B.n619 B.n269 585
R395 B.n269 B.n268 585
R396 B.n621 B.n620 585
R397 B.n622 B.n621 585
R398 B.n263 B.n262 585
R399 B.n264 B.n263 585
R400 B.n631 B.n630 585
R401 B.n630 B.n629 585
R402 B.n632 B.n261 585
R403 B.n628 B.n261 585
R404 B.n634 B.n633 585
R405 B.n635 B.n634 585
R406 B.n256 B.n255 585
R407 B.n257 B.n256 585
R408 B.n644 B.n643 585
R409 B.n643 B.n642 585
R410 B.n645 B.n254 585
R411 B.n254 B.n253 585
R412 B.n647 B.n646 585
R413 B.n648 B.n647 585
R414 B.n2 B.n0 585
R415 B.n4 B.n2 585
R416 B.n3 B.n1 585
R417 B.n809 B.n3 585
R418 B.n807 B.n806 585
R419 B.n808 B.n807 585
R420 B.n805 B.n9 585
R421 B.n9 B.n8 585
R422 B.n804 B.n803 585
R423 B.n803 B.n802 585
R424 B.n11 B.n10 585
R425 B.n801 B.n11 585
R426 B.n799 B.n798 585
R427 B.n800 B.n799 585
R428 B.n797 B.n15 585
R429 B.n18 B.n15 585
R430 B.n796 B.n795 585
R431 B.n795 B.n794 585
R432 B.n17 B.n16 585
R433 B.n793 B.n17 585
R434 B.n791 B.n790 585
R435 B.n792 B.n791 585
R436 B.n789 B.n23 585
R437 B.n23 B.n22 585
R438 B.n788 B.n787 585
R439 B.n787 B.n786 585
R440 B.n25 B.n24 585
R441 B.n785 B.n25 585
R442 B.n783 B.n782 585
R443 B.n784 B.n783 585
R444 B.n781 B.n30 585
R445 B.n30 B.n29 585
R446 B.n780 B.n779 585
R447 B.n779 B.n778 585
R448 B.n32 B.n31 585
R449 B.n777 B.n32 585
R450 B.n775 B.n774 585
R451 B.n776 B.n775 585
R452 B.n773 B.n37 585
R453 B.n37 B.n36 585
R454 B.n772 B.n771 585
R455 B.n771 B.n770 585
R456 B.n39 B.n38 585
R457 B.n769 B.n39 585
R458 B.n767 B.n766 585
R459 B.n768 B.n767 585
R460 B.n765 B.n44 585
R461 B.n44 B.n43 585
R462 B.n764 B.n763 585
R463 B.n763 B.n762 585
R464 B.n46 B.n45 585
R465 B.n761 B.n46 585
R466 B.n759 B.n758 585
R467 B.n760 B.n759 585
R468 B.n757 B.n51 585
R469 B.n51 B.n50 585
R470 B.n756 B.n755 585
R471 B.n755 B.n754 585
R472 B.n53 B.n52 585
R473 B.n753 B.n53 585
R474 B.n751 B.n750 585
R475 B.n752 B.n751 585
R476 B.n749 B.n58 585
R477 B.n58 B.n57 585
R478 B.n748 B.n747 585
R479 B.n747 B.n746 585
R480 B.n60 B.n59 585
R481 B.n745 B.n60 585
R482 B.n743 B.n742 585
R483 B.n744 B.n743 585
R484 B.n741 B.n65 585
R485 B.n65 B.n64 585
R486 B.n740 B.n739 585
R487 B.n739 B.n738 585
R488 B.n67 B.n66 585
R489 B.n737 B.n67 585
R490 B.n735 B.n734 585
R491 B.n736 B.n735 585
R492 B.n733 B.n71 585
R493 B.n74 B.n71 585
R494 B.n732 B.n731 585
R495 B.n731 B.n730 585
R496 B.n73 B.n72 585
R497 B.n729 B.n73 585
R498 B.n727 B.n726 585
R499 B.n728 B.n727 585
R500 B.n725 B.n79 585
R501 B.n79 B.n78 585
R502 B.n724 B.n723 585
R503 B.n723 B.n722 585
R504 B.n81 B.n80 585
R505 B.n721 B.n81 585
R506 B.n719 B.n718 585
R507 B.n720 B.n719 585
R508 B.n717 B.n86 585
R509 B.n86 B.n85 585
R510 B.n812 B.n811 585
R511 B.n811 B.n810 585
R512 B.n508 B.n340 487.695
R513 B.n715 B.n86 487.695
R514 B.n380 B.n338 487.695
R515 B.n712 B.n121 487.695
R516 B.n377 B.t14 267.536
R517 B.n375 B.t6 267.536
R518 B.n124 B.t10 267.536
R519 B.n122 B.t17 267.536
R520 B.n377 B.t16 264.616
R521 B.n122 B.t18 264.616
R522 B.n375 B.t9 264.616
R523 B.n124 B.t12 264.616
R524 B.n713 B.n119 256.663
R525 B.n713 B.n118 256.663
R526 B.n713 B.n117 256.663
R527 B.n713 B.n116 256.663
R528 B.n713 B.n115 256.663
R529 B.n713 B.n114 256.663
R530 B.n713 B.n113 256.663
R531 B.n713 B.n112 256.663
R532 B.n713 B.n111 256.663
R533 B.n713 B.n110 256.663
R534 B.n713 B.n109 256.663
R535 B.n713 B.n108 256.663
R536 B.n713 B.n107 256.663
R537 B.n713 B.n106 256.663
R538 B.n713 B.n105 256.663
R539 B.n713 B.n104 256.663
R540 B.n713 B.n103 256.663
R541 B.n713 B.n102 256.663
R542 B.n713 B.n101 256.663
R543 B.n713 B.n100 256.663
R544 B.n713 B.n99 256.663
R545 B.n713 B.n98 256.663
R546 B.n713 B.n97 256.663
R547 B.n713 B.n96 256.663
R548 B.n713 B.n95 256.663
R549 B.n713 B.n94 256.663
R550 B.n713 B.n93 256.663
R551 B.n713 B.n92 256.663
R552 B.n713 B.n91 256.663
R553 B.n713 B.n90 256.663
R554 B.n713 B.n89 256.663
R555 B.n714 B.n713 256.663
R556 B.n507 B.n506 256.663
R557 B.n506 B.n343 256.663
R558 B.n506 B.n344 256.663
R559 B.n506 B.n345 256.663
R560 B.n506 B.n346 256.663
R561 B.n506 B.n347 256.663
R562 B.n506 B.n348 256.663
R563 B.n506 B.n349 256.663
R564 B.n506 B.n350 256.663
R565 B.n506 B.n351 256.663
R566 B.n506 B.n352 256.663
R567 B.n506 B.n353 256.663
R568 B.n506 B.n354 256.663
R569 B.n506 B.n355 256.663
R570 B.n506 B.n356 256.663
R571 B.n506 B.n357 256.663
R572 B.n506 B.n358 256.663
R573 B.n506 B.n359 256.663
R574 B.n506 B.n360 256.663
R575 B.n506 B.n361 256.663
R576 B.n506 B.n362 256.663
R577 B.n506 B.n363 256.663
R578 B.n506 B.n364 256.663
R579 B.n506 B.n365 256.663
R580 B.n506 B.n366 256.663
R581 B.n506 B.n367 256.663
R582 B.n506 B.n368 256.663
R583 B.n506 B.n369 256.663
R584 B.n506 B.n370 256.663
R585 B.n506 B.n371 256.663
R586 B.n506 B.n372 256.663
R587 B.n506 B.n373 256.663
R588 B.n378 B.t15 200.617
R589 B.n123 B.t19 200.617
R590 B.n376 B.t8 200.617
R591 B.n125 B.t13 200.617
R592 B.n512 B.n340 163.367
R593 B.n512 B.n334 163.367
R594 B.n520 B.n334 163.367
R595 B.n520 B.n332 163.367
R596 B.n524 B.n332 163.367
R597 B.n524 B.n326 163.367
R598 B.n533 B.n326 163.367
R599 B.n533 B.n324 163.367
R600 B.n537 B.n324 163.367
R601 B.n537 B.n319 163.367
R602 B.n545 B.n319 163.367
R603 B.n545 B.n317 163.367
R604 B.n549 B.n317 163.367
R605 B.n549 B.n311 163.367
R606 B.n557 B.n311 163.367
R607 B.n557 B.n309 163.367
R608 B.n561 B.n309 163.367
R609 B.n561 B.n303 163.367
R610 B.n569 B.n303 163.367
R611 B.n569 B.n301 163.367
R612 B.n573 B.n301 163.367
R613 B.n573 B.n295 163.367
R614 B.n581 B.n295 163.367
R615 B.n581 B.n293 163.367
R616 B.n585 B.n293 163.367
R617 B.n585 B.n287 163.367
R618 B.n593 B.n287 163.367
R619 B.n593 B.n285 163.367
R620 B.n597 B.n285 163.367
R621 B.n597 B.n279 163.367
R622 B.n605 B.n279 163.367
R623 B.n605 B.n277 163.367
R624 B.n609 B.n277 163.367
R625 B.n609 B.n271 163.367
R626 B.n617 B.n271 163.367
R627 B.n617 B.n269 163.367
R628 B.n621 B.n269 163.367
R629 B.n621 B.n263 163.367
R630 B.n630 B.n263 163.367
R631 B.n630 B.n261 163.367
R632 B.n634 B.n261 163.367
R633 B.n634 B.n256 163.367
R634 B.n643 B.n256 163.367
R635 B.n643 B.n254 163.367
R636 B.n647 B.n254 163.367
R637 B.n647 B.n2 163.367
R638 B.n811 B.n2 163.367
R639 B.n811 B.n3 163.367
R640 B.n807 B.n3 163.367
R641 B.n807 B.n9 163.367
R642 B.n803 B.n9 163.367
R643 B.n803 B.n11 163.367
R644 B.n799 B.n11 163.367
R645 B.n799 B.n15 163.367
R646 B.n795 B.n15 163.367
R647 B.n795 B.n17 163.367
R648 B.n791 B.n17 163.367
R649 B.n791 B.n23 163.367
R650 B.n787 B.n23 163.367
R651 B.n787 B.n25 163.367
R652 B.n783 B.n25 163.367
R653 B.n783 B.n30 163.367
R654 B.n779 B.n30 163.367
R655 B.n779 B.n32 163.367
R656 B.n775 B.n32 163.367
R657 B.n775 B.n37 163.367
R658 B.n771 B.n37 163.367
R659 B.n771 B.n39 163.367
R660 B.n767 B.n39 163.367
R661 B.n767 B.n44 163.367
R662 B.n763 B.n44 163.367
R663 B.n763 B.n46 163.367
R664 B.n759 B.n46 163.367
R665 B.n759 B.n51 163.367
R666 B.n755 B.n51 163.367
R667 B.n755 B.n53 163.367
R668 B.n751 B.n53 163.367
R669 B.n751 B.n58 163.367
R670 B.n747 B.n58 163.367
R671 B.n747 B.n60 163.367
R672 B.n743 B.n60 163.367
R673 B.n743 B.n65 163.367
R674 B.n739 B.n65 163.367
R675 B.n739 B.n67 163.367
R676 B.n735 B.n67 163.367
R677 B.n735 B.n71 163.367
R678 B.n731 B.n71 163.367
R679 B.n731 B.n73 163.367
R680 B.n727 B.n73 163.367
R681 B.n727 B.n79 163.367
R682 B.n723 B.n79 163.367
R683 B.n723 B.n81 163.367
R684 B.n719 B.n81 163.367
R685 B.n719 B.n86 163.367
R686 B.n505 B.n342 163.367
R687 B.n505 B.n374 163.367
R688 B.n501 B.n500 163.367
R689 B.n497 B.n496 163.367
R690 B.n493 B.n492 163.367
R691 B.n489 B.n488 163.367
R692 B.n485 B.n484 163.367
R693 B.n481 B.n480 163.367
R694 B.n477 B.n476 163.367
R695 B.n473 B.n472 163.367
R696 B.n469 B.n468 163.367
R697 B.n465 B.n464 163.367
R698 B.n461 B.n460 163.367
R699 B.n457 B.n456 163.367
R700 B.n452 B.n451 163.367
R701 B.n448 B.n447 163.367
R702 B.n444 B.n443 163.367
R703 B.n440 B.n439 163.367
R704 B.n436 B.n435 163.367
R705 B.n432 B.n431 163.367
R706 B.n428 B.n427 163.367
R707 B.n424 B.n423 163.367
R708 B.n420 B.n419 163.367
R709 B.n416 B.n415 163.367
R710 B.n412 B.n411 163.367
R711 B.n408 B.n407 163.367
R712 B.n404 B.n403 163.367
R713 B.n400 B.n399 163.367
R714 B.n396 B.n395 163.367
R715 B.n392 B.n391 163.367
R716 B.n388 B.n387 163.367
R717 B.n384 B.n383 163.367
R718 B.n514 B.n338 163.367
R719 B.n514 B.n336 163.367
R720 B.n518 B.n336 163.367
R721 B.n518 B.n330 163.367
R722 B.n526 B.n330 163.367
R723 B.n526 B.n328 163.367
R724 B.n530 B.n328 163.367
R725 B.n530 B.n323 163.367
R726 B.n539 B.n323 163.367
R727 B.n539 B.n321 163.367
R728 B.n543 B.n321 163.367
R729 B.n543 B.n315 163.367
R730 B.n551 B.n315 163.367
R731 B.n551 B.n313 163.367
R732 B.n555 B.n313 163.367
R733 B.n555 B.n307 163.367
R734 B.n563 B.n307 163.367
R735 B.n563 B.n305 163.367
R736 B.n567 B.n305 163.367
R737 B.n567 B.n299 163.367
R738 B.n575 B.n299 163.367
R739 B.n575 B.n297 163.367
R740 B.n579 B.n297 163.367
R741 B.n579 B.n291 163.367
R742 B.n587 B.n291 163.367
R743 B.n587 B.n289 163.367
R744 B.n591 B.n289 163.367
R745 B.n591 B.n282 163.367
R746 B.n599 B.n282 163.367
R747 B.n599 B.n280 163.367
R748 B.n603 B.n280 163.367
R749 B.n603 B.n275 163.367
R750 B.n611 B.n275 163.367
R751 B.n611 B.n273 163.367
R752 B.n615 B.n273 163.367
R753 B.n615 B.n267 163.367
R754 B.n623 B.n267 163.367
R755 B.n623 B.n265 163.367
R756 B.n627 B.n265 163.367
R757 B.n627 B.n260 163.367
R758 B.n636 B.n260 163.367
R759 B.n636 B.n258 163.367
R760 B.n641 B.n258 163.367
R761 B.n641 B.n252 163.367
R762 B.n649 B.n252 163.367
R763 B.n650 B.n649 163.367
R764 B.n650 B.n5 163.367
R765 B.n6 B.n5 163.367
R766 B.n7 B.n6 163.367
R767 B.n655 B.n7 163.367
R768 B.n655 B.n12 163.367
R769 B.n13 B.n12 163.367
R770 B.n14 B.n13 163.367
R771 B.n660 B.n14 163.367
R772 B.n660 B.n19 163.367
R773 B.n20 B.n19 163.367
R774 B.n21 B.n20 163.367
R775 B.n665 B.n21 163.367
R776 B.n665 B.n26 163.367
R777 B.n27 B.n26 163.367
R778 B.n28 B.n27 163.367
R779 B.n670 B.n28 163.367
R780 B.n670 B.n33 163.367
R781 B.n34 B.n33 163.367
R782 B.n35 B.n34 163.367
R783 B.n675 B.n35 163.367
R784 B.n675 B.n40 163.367
R785 B.n41 B.n40 163.367
R786 B.n42 B.n41 163.367
R787 B.n680 B.n42 163.367
R788 B.n680 B.n47 163.367
R789 B.n48 B.n47 163.367
R790 B.n49 B.n48 163.367
R791 B.n685 B.n49 163.367
R792 B.n685 B.n54 163.367
R793 B.n55 B.n54 163.367
R794 B.n56 B.n55 163.367
R795 B.n690 B.n56 163.367
R796 B.n690 B.n61 163.367
R797 B.n62 B.n61 163.367
R798 B.n63 B.n62 163.367
R799 B.n695 B.n63 163.367
R800 B.n695 B.n68 163.367
R801 B.n69 B.n68 163.367
R802 B.n70 B.n69 163.367
R803 B.n700 B.n70 163.367
R804 B.n700 B.n75 163.367
R805 B.n76 B.n75 163.367
R806 B.n77 B.n76 163.367
R807 B.n705 B.n77 163.367
R808 B.n705 B.n82 163.367
R809 B.n83 B.n82 163.367
R810 B.n84 B.n83 163.367
R811 B.n121 B.n84 163.367
R812 B.n127 B.n88 163.367
R813 B.n131 B.n130 163.367
R814 B.n135 B.n134 163.367
R815 B.n139 B.n138 163.367
R816 B.n143 B.n142 163.367
R817 B.n147 B.n146 163.367
R818 B.n151 B.n150 163.367
R819 B.n155 B.n154 163.367
R820 B.n159 B.n158 163.367
R821 B.n163 B.n162 163.367
R822 B.n167 B.n166 163.367
R823 B.n171 B.n170 163.367
R824 B.n175 B.n174 163.367
R825 B.n179 B.n178 163.367
R826 B.n183 B.n182 163.367
R827 B.n187 B.n186 163.367
R828 B.n191 B.n190 163.367
R829 B.n195 B.n194 163.367
R830 B.n200 B.n199 163.367
R831 B.n204 B.n203 163.367
R832 B.n208 B.n207 163.367
R833 B.n212 B.n211 163.367
R834 B.n216 B.n215 163.367
R835 B.n220 B.n219 163.367
R836 B.n224 B.n223 163.367
R837 B.n228 B.n227 163.367
R838 B.n232 B.n231 163.367
R839 B.n236 B.n235 163.367
R840 B.n240 B.n239 163.367
R841 B.n244 B.n243 163.367
R842 B.n248 B.n247 163.367
R843 B.n712 B.n120 163.367
R844 B.n506 B.n339 104.344
R845 B.n713 B.n85 104.344
R846 B.n508 B.n507 71.676
R847 B.n374 B.n343 71.676
R848 B.n500 B.n344 71.676
R849 B.n496 B.n345 71.676
R850 B.n492 B.n346 71.676
R851 B.n488 B.n347 71.676
R852 B.n484 B.n348 71.676
R853 B.n480 B.n349 71.676
R854 B.n476 B.n350 71.676
R855 B.n472 B.n351 71.676
R856 B.n468 B.n352 71.676
R857 B.n464 B.n353 71.676
R858 B.n460 B.n354 71.676
R859 B.n456 B.n355 71.676
R860 B.n451 B.n356 71.676
R861 B.n447 B.n357 71.676
R862 B.n443 B.n358 71.676
R863 B.n439 B.n359 71.676
R864 B.n435 B.n360 71.676
R865 B.n431 B.n361 71.676
R866 B.n427 B.n362 71.676
R867 B.n423 B.n363 71.676
R868 B.n419 B.n364 71.676
R869 B.n415 B.n365 71.676
R870 B.n411 B.n366 71.676
R871 B.n407 B.n367 71.676
R872 B.n403 B.n368 71.676
R873 B.n399 B.n369 71.676
R874 B.n395 B.n370 71.676
R875 B.n391 B.n371 71.676
R876 B.n387 B.n372 71.676
R877 B.n383 B.n373 71.676
R878 B.n715 B.n714 71.676
R879 B.n127 B.n89 71.676
R880 B.n131 B.n90 71.676
R881 B.n135 B.n91 71.676
R882 B.n139 B.n92 71.676
R883 B.n143 B.n93 71.676
R884 B.n147 B.n94 71.676
R885 B.n151 B.n95 71.676
R886 B.n155 B.n96 71.676
R887 B.n159 B.n97 71.676
R888 B.n163 B.n98 71.676
R889 B.n167 B.n99 71.676
R890 B.n171 B.n100 71.676
R891 B.n175 B.n101 71.676
R892 B.n179 B.n102 71.676
R893 B.n183 B.n103 71.676
R894 B.n187 B.n104 71.676
R895 B.n191 B.n105 71.676
R896 B.n195 B.n106 71.676
R897 B.n200 B.n107 71.676
R898 B.n204 B.n108 71.676
R899 B.n208 B.n109 71.676
R900 B.n212 B.n110 71.676
R901 B.n216 B.n111 71.676
R902 B.n220 B.n112 71.676
R903 B.n224 B.n113 71.676
R904 B.n228 B.n114 71.676
R905 B.n232 B.n115 71.676
R906 B.n236 B.n116 71.676
R907 B.n240 B.n117 71.676
R908 B.n244 B.n118 71.676
R909 B.n248 B.n119 71.676
R910 B.n120 B.n119 71.676
R911 B.n247 B.n118 71.676
R912 B.n243 B.n117 71.676
R913 B.n239 B.n116 71.676
R914 B.n235 B.n115 71.676
R915 B.n231 B.n114 71.676
R916 B.n227 B.n113 71.676
R917 B.n223 B.n112 71.676
R918 B.n219 B.n111 71.676
R919 B.n215 B.n110 71.676
R920 B.n211 B.n109 71.676
R921 B.n207 B.n108 71.676
R922 B.n203 B.n107 71.676
R923 B.n199 B.n106 71.676
R924 B.n194 B.n105 71.676
R925 B.n190 B.n104 71.676
R926 B.n186 B.n103 71.676
R927 B.n182 B.n102 71.676
R928 B.n178 B.n101 71.676
R929 B.n174 B.n100 71.676
R930 B.n170 B.n99 71.676
R931 B.n166 B.n98 71.676
R932 B.n162 B.n97 71.676
R933 B.n158 B.n96 71.676
R934 B.n154 B.n95 71.676
R935 B.n150 B.n94 71.676
R936 B.n146 B.n93 71.676
R937 B.n142 B.n92 71.676
R938 B.n138 B.n91 71.676
R939 B.n134 B.n90 71.676
R940 B.n130 B.n89 71.676
R941 B.n714 B.n88 71.676
R942 B.n507 B.n342 71.676
R943 B.n501 B.n343 71.676
R944 B.n497 B.n344 71.676
R945 B.n493 B.n345 71.676
R946 B.n489 B.n346 71.676
R947 B.n485 B.n347 71.676
R948 B.n481 B.n348 71.676
R949 B.n477 B.n349 71.676
R950 B.n473 B.n350 71.676
R951 B.n469 B.n351 71.676
R952 B.n465 B.n352 71.676
R953 B.n461 B.n353 71.676
R954 B.n457 B.n354 71.676
R955 B.n452 B.n355 71.676
R956 B.n448 B.n356 71.676
R957 B.n444 B.n357 71.676
R958 B.n440 B.n358 71.676
R959 B.n436 B.n359 71.676
R960 B.n432 B.n360 71.676
R961 B.n428 B.n361 71.676
R962 B.n424 B.n362 71.676
R963 B.n420 B.n363 71.676
R964 B.n416 B.n364 71.676
R965 B.n412 B.n365 71.676
R966 B.n408 B.n366 71.676
R967 B.n404 B.n367 71.676
R968 B.n400 B.n368 71.676
R969 B.n396 B.n369 71.676
R970 B.n392 B.n370 71.676
R971 B.n388 B.n371 71.676
R972 B.n384 B.n372 71.676
R973 B.n380 B.n373 71.676
R974 B.n378 B.n377 64.0005
R975 B.n376 B.n375 64.0005
R976 B.n125 B.n124 64.0005
R977 B.n123 B.n122 64.0005
R978 B.n513 B.n339 59.6258
R979 B.n513 B.n335 59.6258
R980 B.n519 B.n335 59.6258
R981 B.n519 B.n331 59.6258
R982 B.n525 B.n331 59.6258
R983 B.n525 B.n327 59.6258
R984 B.n532 B.n327 59.6258
R985 B.n532 B.n531 59.6258
R986 B.n538 B.n320 59.6258
R987 B.n544 B.n320 59.6258
R988 B.n544 B.n316 59.6258
R989 B.n550 B.n316 59.6258
R990 B.n550 B.n312 59.6258
R991 B.n556 B.n312 59.6258
R992 B.n556 B.n308 59.6258
R993 B.n562 B.n308 59.6258
R994 B.n562 B.n304 59.6258
R995 B.n568 B.n304 59.6258
R996 B.n568 B.n300 59.6258
R997 B.n574 B.n300 59.6258
R998 B.n580 B.n296 59.6258
R999 B.n580 B.n292 59.6258
R1000 B.n586 B.n292 59.6258
R1001 B.n586 B.n288 59.6258
R1002 B.n592 B.n288 59.6258
R1003 B.n592 B.n283 59.6258
R1004 B.n598 B.n283 59.6258
R1005 B.n598 B.n284 59.6258
R1006 B.n604 B.n276 59.6258
R1007 B.n610 B.n276 59.6258
R1008 B.n610 B.n272 59.6258
R1009 B.n616 B.n272 59.6258
R1010 B.n616 B.n268 59.6258
R1011 B.n622 B.n268 59.6258
R1012 B.n622 B.n264 59.6258
R1013 B.n629 B.n264 59.6258
R1014 B.n629 B.n628 59.6258
R1015 B.n635 B.n257 59.6258
R1016 B.n642 B.n257 59.6258
R1017 B.n642 B.n253 59.6258
R1018 B.n648 B.n253 59.6258
R1019 B.n648 B.n4 59.6258
R1020 B.n810 B.n4 59.6258
R1021 B.n810 B.n809 59.6258
R1022 B.n809 B.n808 59.6258
R1023 B.n808 B.n8 59.6258
R1024 B.n802 B.n8 59.6258
R1025 B.n802 B.n801 59.6258
R1026 B.n801 B.n800 59.6258
R1027 B.n794 B.n18 59.6258
R1028 B.n794 B.n793 59.6258
R1029 B.n793 B.n792 59.6258
R1030 B.n792 B.n22 59.6258
R1031 B.n786 B.n22 59.6258
R1032 B.n786 B.n785 59.6258
R1033 B.n785 B.n784 59.6258
R1034 B.n784 B.n29 59.6258
R1035 B.n778 B.n29 59.6258
R1036 B.n777 B.n776 59.6258
R1037 B.n776 B.n36 59.6258
R1038 B.n770 B.n36 59.6258
R1039 B.n770 B.n769 59.6258
R1040 B.n769 B.n768 59.6258
R1041 B.n768 B.n43 59.6258
R1042 B.n762 B.n43 59.6258
R1043 B.n762 B.n761 59.6258
R1044 B.n760 B.n50 59.6258
R1045 B.n754 B.n50 59.6258
R1046 B.n754 B.n753 59.6258
R1047 B.n753 B.n752 59.6258
R1048 B.n752 B.n57 59.6258
R1049 B.n746 B.n57 59.6258
R1050 B.n746 B.n745 59.6258
R1051 B.n745 B.n744 59.6258
R1052 B.n744 B.n64 59.6258
R1053 B.n738 B.n64 59.6258
R1054 B.n738 B.n737 59.6258
R1055 B.n737 B.n736 59.6258
R1056 B.n730 B.n74 59.6258
R1057 B.n730 B.n729 59.6258
R1058 B.n729 B.n728 59.6258
R1059 B.n728 B.n78 59.6258
R1060 B.n722 B.n78 59.6258
R1061 B.n722 B.n721 59.6258
R1062 B.n721 B.n720 59.6258
R1063 B.n720 B.n85 59.6258
R1064 B.n379 B.n378 59.5399
R1065 B.n454 B.n376 59.5399
R1066 B.n126 B.n125 59.5399
R1067 B.n197 B.n123 59.5399
R1068 B.t5 B.n296 51.7343
R1069 B.n761 B.t0 51.7343
R1070 B.n284 B.t2 49.9806
R1071 B.t1 B.n777 49.9806
R1072 B.n538 B.t7 46.4732
R1073 B.n736 B.t11 46.4732
R1074 B.n628 B.t3 32.4437
R1075 B.n18 B.t4 32.4437
R1076 B.n717 B.n716 31.6883
R1077 B.n711 B.n710 31.6883
R1078 B.n381 B.n337 31.6883
R1079 B.n510 B.n509 31.6883
R1080 B.n635 B.t3 27.1826
R1081 B.n800 B.t4 27.1826
R1082 B B.n812 18.0485
R1083 B.n531 B.t7 13.1532
R1084 B.n74 B.t11 13.1532
R1085 B.n716 B.n87 10.6151
R1086 B.n128 B.n87 10.6151
R1087 B.n129 B.n128 10.6151
R1088 B.n132 B.n129 10.6151
R1089 B.n133 B.n132 10.6151
R1090 B.n136 B.n133 10.6151
R1091 B.n137 B.n136 10.6151
R1092 B.n140 B.n137 10.6151
R1093 B.n141 B.n140 10.6151
R1094 B.n144 B.n141 10.6151
R1095 B.n145 B.n144 10.6151
R1096 B.n148 B.n145 10.6151
R1097 B.n149 B.n148 10.6151
R1098 B.n152 B.n149 10.6151
R1099 B.n153 B.n152 10.6151
R1100 B.n156 B.n153 10.6151
R1101 B.n157 B.n156 10.6151
R1102 B.n160 B.n157 10.6151
R1103 B.n161 B.n160 10.6151
R1104 B.n164 B.n161 10.6151
R1105 B.n165 B.n164 10.6151
R1106 B.n168 B.n165 10.6151
R1107 B.n169 B.n168 10.6151
R1108 B.n172 B.n169 10.6151
R1109 B.n173 B.n172 10.6151
R1110 B.n176 B.n173 10.6151
R1111 B.n177 B.n176 10.6151
R1112 B.n181 B.n180 10.6151
R1113 B.n184 B.n181 10.6151
R1114 B.n185 B.n184 10.6151
R1115 B.n188 B.n185 10.6151
R1116 B.n189 B.n188 10.6151
R1117 B.n192 B.n189 10.6151
R1118 B.n193 B.n192 10.6151
R1119 B.n196 B.n193 10.6151
R1120 B.n201 B.n198 10.6151
R1121 B.n202 B.n201 10.6151
R1122 B.n205 B.n202 10.6151
R1123 B.n206 B.n205 10.6151
R1124 B.n209 B.n206 10.6151
R1125 B.n210 B.n209 10.6151
R1126 B.n213 B.n210 10.6151
R1127 B.n214 B.n213 10.6151
R1128 B.n217 B.n214 10.6151
R1129 B.n218 B.n217 10.6151
R1130 B.n221 B.n218 10.6151
R1131 B.n222 B.n221 10.6151
R1132 B.n225 B.n222 10.6151
R1133 B.n226 B.n225 10.6151
R1134 B.n229 B.n226 10.6151
R1135 B.n230 B.n229 10.6151
R1136 B.n233 B.n230 10.6151
R1137 B.n234 B.n233 10.6151
R1138 B.n237 B.n234 10.6151
R1139 B.n238 B.n237 10.6151
R1140 B.n241 B.n238 10.6151
R1141 B.n242 B.n241 10.6151
R1142 B.n245 B.n242 10.6151
R1143 B.n246 B.n245 10.6151
R1144 B.n249 B.n246 10.6151
R1145 B.n250 B.n249 10.6151
R1146 B.n711 B.n250 10.6151
R1147 B.n515 B.n337 10.6151
R1148 B.n516 B.n515 10.6151
R1149 B.n517 B.n516 10.6151
R1150 B.n517 B.n329 10.6151
R1151 B.n527 B.n329 10.6151
R1152 B.n528 B.n527 10.6151
R1153 B.n529 B.n528 10.6151
R1154 B.n529 B.n322 10.6151
R1155 B.n540 B.n322 10.6151
R1156 B.n541 B.n540 10.6151
R1157 B.n542 B.n541 10.6151
R1158 B.n542 B.n314 10.6151
R1159 B.n552 B.n314 10.6151
R1160 B.n553 B.n552 10.6151
R1161 B.n554 B.n553 10.6151
R1162 B.n554 B.n306 10.6151
R1163 B.n564 B.n306 10.6151
R1164 B.n565 B.n564 10.6151
R1165 B.n566 B.n565 10.6151
R1166 B.n566 B.n298 10.6151
R1167 B.n576 B.n298 10.6151
R1168 B.n577 B.n576 10.6151
R1169 B.n578 B.n577 10.6151
R1170 B.n578 B.n290 10.6151
R1171 B.n588 B.n290 10.6151
R1172 B.n589 B.n588 10.6151
R1173 B.n590 B.n589 10.6151
R1174 B.n590 B.n281 10.6151
R1175 B.n600 B.n281 10.6151
R1176 B.n601 B.n600 10.6151
R1177 B.n602 B.n601 10.6151
R1178 B.n602 B.n274 10.6151
R1179 B.n612 B.n274 10.6151
R1180 B.n613 B.n612 10.6151
R1181 B.n614 B.n613 10.6151
R1182 B.n614 B.n266 10.6151
R1183 B.n624 B.n266 10.6151
R1184 B.n625 B.n624 10.6151
R1185 B.n626 B.n625 10.6151
R1186 B.n626 B.n259 10.6151
R1187 B.n637 B.n259 10.6151
R1188 B.n638 B.n637 10.6151
R1189 B.n640 B.n638 10.6151
R1190 B.n640 B.n639 10.6151
R1191 B.n639 B.n251 10.6151
R1192 B.n651 B.n251 10.6151
R1193 B.n652 B.n651 10.6151
R1194 B.n653 B.n652 10.6151
R1195 B.n654 B.n653 10.6151
R1196 B.n656 B.n654 10.6151
R1197 B.n657 B.n656 10.6151
R1198 B.n658 B.n657 10.6151
R1199 B.n659 B.n658 10.6151
R1200 B.n661 B.n659 10.6151
R1201 B.n662 B.n661 10.6151
R1202 B.n663 B.n662 10.6151
R1203 B.n664 B.n663 10.6151
R1204 B.n666 B.n664 10.6151
R1205 B.n667 B.n666 10.6151
R1206 B.n668 B.n667 10.6151
R1207 B.n669 B.n668 10.6151
R1208 B.n671 B.n669 10.6151
R1209 B.n672 B.n671 10.6151
R1210 B.n673 B.n672 10.6151
R1211 B.n674 B.n673 10.6151
R1212 B.n676 B.n674 10.6151
R1213 B.n677 B.n676 10.6151
R1214 B.n678 B.n677 10.6151
R1215 B.n679 B.n678 10.6151
R1216 B.n681 B.n679 10.6151
R1217 B.n682 B.n681 10.6151
R1218 B.n683 B.n682 10.6151
R1219 B.n684 B.n683 10.6151
R1220 B.n686 B.n684 10.6151
R1221 B.n687 B.n686 10.6151
R1222 B.n688 B.n687 10.6151
R1223 B.n689 B.n688 10.6151
R1224 B.n691 B.n689 10.6151
R1225 B.n692 B.n691 10.6151
R1226 B.n693 B.n692 10.6151
R1227 B.n694 B.n693 10.6151
R1228 B.n696 B.n694 10.6151
R1229 B.n697 B.n696 10.6151
R1230 B.n698 B.n697 10.6151
R1231 B.n699 B.n698 10.6151
R1232 B.n701 B.n699 10.6151
R1233 B.n702 B.n701 10.6151
R1234 B.n703 B.n702 10.6151
R1235 B.n704 B.n703 10.6151
R1236 B.n706 B.n704 10.6151
R1237 B.n707 B.n706 10.6151
R1238 B.n708 B.n707 10.6151
R1239 B.n709 B.n708 10.6151
R1240 B.n710 B.n709 10.6151
R1241 B.n509 B.n341 10.6151
R1242 B.n504 B.n341 10.6151
R1243 B.n504 B.n503 10.6151
R1244 B.n503 B.n502 10.6151
R1245 B.n502 B.n499 10.6151
R1246 B.n499 B.n498 10.6151
R1247 B.n498 B.n495 10.6151
R1248 B.n495 B.n494 10.6151
R1249 B.n494 B.n491 10.6151
R1250 B.n491 B.n490 10.6151
R1251 B.n490 B.n487 10.6151
R1252 B.n487 B.n486 10.6151
R1253 B.n486 B.n483 10.6151
R1254 B.n483 B.n482 10.6151
R1255 B.n482 B.n479 10.6151
R1256 B.n479 B.n478 10.6151
R1257 B.n478 B.n475 10.6151
R1258 B.n475 B.n474 10.6151
R1259 B.n474 B.n471 10.6151
R1260 B.n471 B.n470 10.6151
R1261 B.n470 B.n467 10.6151
R1262 B.n467 B.n466 10.6151
R1263 B.n466 B.n463 10.6151
R1264 B.n463 B.n462 10.6151
R1265 B.n462 B.n459 10.6151
R1266 B.n459 B.n458 10.6151
R1267 B.n458 B.n455 10.6151
R1268 B.n453 B.n450 10.6151
R1269 B.n450 B.n449 10.6151
R1270 B.n449 B.n446 10.6151
R1271 B.n446 B.n445 10.6151
R1272 B.n445 B.n442 10.6151
R1273 B.n442 B.n441 10.6151
R1274 B.n441 B.n438 10.6151
R1275 B.n438 B.n437 10.6151
R1276 B.n434 B.n433 10.6151
R1277 B.n433 B.n430 10.6151
R1278 B.n430 B.n429 10.6151
R1279 B.n429 B.n426 10.6151
R1280 B.n426 B.n425 10.6151
R1281 B.n425 B.n422 10.6151
R1282 B.n422 B.n421 10.6151
R1283 B.n421 B.n418 10.6151
R1284 B.n418 B.n417 10.6151
R1285 B.n417 B.n414 10.6151
R1286 B.n414 B.n413 10.6151
R1287 B.n413 B.n410 10.6151
R1288 B.n410 B.n409 10.6151
R1289 B.n409 B.n406 10.6151
R1290 B.n406 B.n405 10.6151
R1291 B.n405 B.n402 10.6151
R1292 B.n402 B.n401 10.6151
R1293 B.n401 B.n398 10.6151
R1294 B.n398 B.n397 10.6151
R1295 B.n397 B.n394 10.6151
R1296 B.n394 B.n393 10.6151
R1297 B.n393 B.n390 10.6151
R1298 B.n390 B.n389 10.6151
R1299 B.n389 B.n386 10.6151
R1300 B.n386 B.n385 10.6151
R1301 B.n385 B.n382 10.6151
R1302 B.n382 B.n381 10.6151
R1303 B.n511 B.n510 10.6151
R1304 B.n511 B.n333 10.6151
R1305 B.n521 B.n333 10.6151
R1306 B.n522 B.n521 10.6151
R1307 B.n523 B.n522 10.6151
R1308 B.n523 B.n325 10.6151
R1309 B.n534 B.n325 10.6151
R1310 B.n535 B.n534 10.6151
R1311 B.n536 B.n535 10.6151
R1312 B.n536 B.n318 10.6151
R1313 B.n546 B.n318 10.6151
R1314 B.n547 B.n546 10.6151
R1315 B.n548 B.n547 10.6151
R1316 B.n548 B.n310 10.6151
R1317 B.n558 B.n310 10.6151
R1318 B.n559 B.n558 10.6151
R1319 B.n560 B.n559 10.6151
R1320 B.n560 B.n302 10.6151
R1321 B.n570 B.n302 10.6151
R1322 B.n571 B.n570 10.6151
R1323 B.n572 B.n571 10.6151
R1324 B.n572 B.n294 10.6151
R1325 B.n582 B.n294 10.6151
R1326 B.n583 B.n582 10.6151
R1327 B.n584 B.n583 10.6151
R1328 B.n584 B.n286 10.6151
R1329 B.n594 B.n286 10.6151
R1330 B.n595 B.n594 10.6151
R1331 B.n596 B.n595 10.6151
R1332 B.n596 B.n278 10.6151
R1333 B.n606 B.n278 10.6151
R1334 B.n607 B.n606 10.6151
R1335 B.n608 B.n607 10.6151
R1336 B.n608 B.n270 10.6151
R1337 B.n618 B.n270 10.6151
R1338 B.n619 B.n618 10.6151
R1339 B.n620 B.n619 10.6151
R1340 B.n620 B.n262 10.6151
R1341 B.n631 B.n262 10.6151
R1342 B.n632 B.n631 10.6151
R1343 B.n633 B.n632 10.6151
R1344 B.n633 B.n255 10.6151
R1345 B.n644 B.n255 10.6151
R1346 B.n645 B.n644 10.6151
R1347 B.n646 B.n645 10.6151
R1348 B.n646 B.n0 10.6151
R1349 B.n806 B.n1 10.6151
R1350 B.n806 B.n805 10.6151
R1351 B.n805 B.n804 10.6151
R1352 B.n804 B.n10 10.6151
R1353 B.n798 B.n10 10.6151
R1354 B.n798 B.n797 10.6151
R1355 B.n797 B.n796 10.6151
R1356 B.n796 B.n16 10.6151
R1357 B.n790 B.n16 10.6151
R1358 B.n790 B.n789 10.6151
R1359 B.n789 B.n788 10.6151
R1360 B.n788 B.n24 10.6151
R1361 B.n782 B.n24 10.6151
R1362 B.n782 B.n781 10.6151
R1363 B.n781 B.n780 10.6151
R1364 B.n780 B.n31 10.6151
R1365 B.n774 B.n31 10.6151
R1366 B.n774 B.n773 10.6151
R1367 B.n773 B.n772 10.6151
R1368 B.n772 B.n38 10.6151
R1369 B.n766 B.n38 10.6151
R1370 B.n766 B.n765 10.6151
R1371 B.n765 B.n764 10.6151
R1372 B.n764 B.n45 10.6151
R1373 B.n758 B.n45 10.6151
R1374 B.n758 B.n757 10.6151
R1375 B.n757 B.n756 10.6151
R1376 B.n756 B.n52 10.6151
R1377 B.n750 B.n52 10.6151
R1378 B.n750 B.n749 10.6151
R1379 B.n749 B.n748 10.6151
R1380 B.n748 B.n59 10.6151
R1381 B.n742 B.n59 10.6151
R1382 B.n742 B.n741 10.6151
R1383 B.n741 B.n740 10.6151
R1384 B.n740 B.n66 10.6151
R1385 B.n734 B.n66 10.6151
R1386 B.n734 B.n733 10.6151
R1387 B.n733 B.n732 10.6151
R1388 B.n732 B.n72 10.6151
R1389 B.n726 B.n72 10.6151
R1390 B.n726 B.n725 10.6151
R1391 B.n725 B.n724 10.6151
R1392 B.n724 B.n80 10.6151
R1393 B.n718 B.n80 10.6151
R1394 B.n718 B.n717 10.6151
R1395 B.n604 B.t2 9.64578
R1396 B.n778 B.t1 9.64578
R1397 B.n574 B.t5 7.89209
R1398 B.t0 B.n760 7.89209
R1399 B.n180 B.n126 6.5566
R1400 B.n197 B.n196 6.5566
R1401 B.n454 B.n453 6.5566
R1402 B.n437 B.n379 6.5566
R1403 B.n177 B.n126 4.05904
R1404 B.n198 B.n197 4.05904
R1405 B.n455 B.n454 4.05904
R1406 B.n434 B.n379 4.05904
R1407 B.n812 B.n0 2.81026
R1408 B.n812 B.n1 2.81026
R1409 VP.n14 VP.n11 161.3
R1410 VP.n16 VP.n15 161.3
R1411 VP.n17 VP.n10 161.3
R1412 VP.n19 VP.n18 161.3
R1413 VP.n20 VP.n9 161.3
R1414 VP.n22 VP.n21 161.3
R1415 VP.n23 VP.n8 161.3
R1416 VP.n48 VP.n0 161.3
R1417 VP.n47 VP.n46 161.3
R1418 VP.n45 VP.n1 161.3
R1419 VP.n44 VP.n43 161.3
R1420 VP.n42 VP.n2 161.3
R1421 VP.n41 VP.n40 161.3
R1422 VP.n39 VP.n3 161.3
R1423 VP.n38 VP.n37 161.3
R1424 VP.n35 VP.n4 161.3
R1425 VP.n34 VP.n33 161.3
R1426 VP.n32 VP.n5 161.3
R1427 VP.n31 VP.n30 161.3
R1428 VP.n29 VP.n6 161.3
R1429 VP.n28 VP.n27 161.3
R1430 VP.n26 VP.n7 108.309
R1431 VP.n50 VP.n49 108.309
R1432 VP.n25 VP.n24 108.309
R1433 VP.n13 VP.t2 91.8434
R1434 VP.n13 VP.n12 61.6401
R1435 VP.n7 VP.t4 58.9928
R1436 VP.n36 VP.t0 58.9928
R1437 VP.n49 VP.t3 58.9928
R1438 VP.n24 VP.t5 58.9928
R1439 VP.n12 VP.t1 58.9928
R1440 VP.n34 VP.n5 50.2061
R1441 VP.n43 VP.n42 50.2061
R1442 VP.n18 VP.n17 50.2061
R1443 VP.n26 VP.n25 46.5375
R1444 VP.n30 VP.n5 30.7807
R1445 VP.n43 VP.n1 30.7807
R1446 VP.n18 VP.n9 30.7807
R1447 VP.n29 VP.n28 24.4675
R1448 VP.n30 VP.n29 24.4675
R1449 VP.n35 VP.n34 24.4675
R1450 VP.n37 VP.n35 24.4675
R1451 VP.n41 VP.n3 24.4675
R1452 VP.n42 VP.n41 24.4675
R1453 VP.n47 VP.n1 24.4675
R1454 VP.n48 VP.n47 24.4675
R1455 VP.n22 VP.n9 24.4675
R1456 VP.n23 VP.n22 24.4675
R1457 VP.n16 VP.n11 24.4675
R1458 VP.n17 VP.n16 24.4675
R1459 VP.n37 VP.n36 12.234
R1460 VP.n36 VP.n3 12.234
R1461 VP.n12 VP.n11 12.234
R1462 VP.n14 VP.n13 5.10511
R1463 VP.n28 VP.n7 2.4472
R1464 VP.n49 VP.n48 2.4472
R1465 VP.n24 VP.n23 2.4472
R1466 VP.n25 VP.n8 0.278367
R1467 VP.n27 VP.n26 0.278367
R1468 VP.n50 VP.n0 0.278367
R1469 VP.n15 VP.n14 0.189894
R1470 VP.n15 VP.n10 0.189894
R1471 VP.n19 VP.n10 0.189894
R1472 VP.n20 VP.n19 0.189894
R1473 VP.n21 VP.n20 0.189894
R1474 VP.n21 VP.n8 0.189894
R1475 VP.n27 VP.n6 0.189894
R1476 VP.n31 VP.n6 0.189894
R1477 VP.n32 VP.n31 0.189894
R1478 VP.n33 VP.n32 0.189894
R1479 VP.n33 VP.n4 0.189894
R1480 VP.n38 VP.n4 0.189894
R1481 VP.n39 VP.n38 0.189894
R1482 VP.n40 VP.n39 0.189894
R1483 VP.n40 VP.n2 0.189894
R1484 VP.n44 VP.n2 0.189894
R1485 VP.n45 VP.n44 0.189894
R1486 VP.n46 VP.n45 0.189894
R1487 VP.n46 VP.n0 0.189894
R1488 VP VP.n50 0.153454
R1489 VDD1.n30 VDD1.n0 214.453
R1490 VDD1.n65 VDD1.n35 214.453
R1491 VDD1.n31 VDD1.n30 185
R1492 VDD1.n29 VDD1.n28 185
R1493 VDD1.n4 VDD1.n3 185
R1494 VDD1.n23 VDD1.n22 185
R1495 VDD1.n21 VDD1.n20 185
R1496 VDD1.n8 VDD1.n7 185
R1497 VDD1.n15 VDD1.n14 185
R1498 VDD1.n13 VDD1.n12 185
R1499 VDD1.n48 VDD1.n47 185
R1500 VDD1.n50 VDD1.n49 185
R1501 VDD1.n43 VDD1.n42 185
R1502 VDD1.n56 VDD1.n55 185
R1503 VDD1.n58 VDD1.n57 185
R1504 VDD1.n39 VDD1.n38 185
R1505 VDD1.n64 VDD1.n63 185
R1506 VDD1.n66 VDD1.n65 185
R1507 VDD1.n46 VDD1.t4 149.524
R1508 VDD1.n11 VDD1.t5 149.524
R1509 VDD1.n30 VDD1.n29 104.615
R1510 VDD1.n29 VDD1.n3 104.615
R1511 VDD1.n22 VDD1.n3 104.615
R1512 VDD1.n22 VDD1.n21 104.615
R1513 VDD1.n21 VDD1.n7 104.615
R1514 VDD1.n14 VDD1.n7 104.615
R1515 VDD1.n14 VDD1.n13 104.615
R1516 VDD1.n49 VDD1.n48 104.615
R1517 VDD1.n49 VDD1.n42 104.615
R1518 VDD1.n56 VDD1.n42 104.615
R1519 VDD1.n57 VDD1.n56 104.615
R1520 VDD1.n57 VDD1.n38 104.615
R1521 VDD1.n64 VDD1.n38 104.615
R1522 VDD1.n65 VDD1.n64 104.615
R1523 VDD1.n71 VDD1.n70 68.9755
R1524 VDD1.n73 VDD1.n72 68.3196
R1525 VDD1 VDD1.n34 54.7408
R1526 VDD1.n71 VDD1.n69 54.6273
R1527 VDD1.n13 VDD1.t5 52.3082
R1528 VDD1.n48 VDD1.t4 52.3082
R1529 VDD1.n73 VDD1.n71 41.2336
R1530 VDD1.n32 VDD1.n31 12.8005
R1531 VDD1.n67 VDD1.n66 12.8005
R1532 VDD1.n28 VDD1.n2 12.0247
R1533 VDD1.n63 VDD1.n37 12.0247
R1534 VDD1.n27 VDD1.n4 11.249
R1535 VDD1.n62 VDD1.n39 11.249
R1536 VDD1.n24 VDD1.n23 10.4732
R1537 VDD1.n59 VDD1.n58 10.4732
R1538 VDD1.n12 VDD1.n11 10.2747
R1539 VDD1.n47 VDD1.n46 10.2747
R1540 VDD1.n20 VDD1.n6 9.69747
R1541 VDD1.n55 VDD1.n41 9.69747
R1542 VDD1.n34 VDD1.n33 9.45567
R1543 VDD1.n69 VDD1.n68 9.45567
R1544 VDD1.n10 VDD1.n9 9.3005
R1545 VDD1.n17 VDD1.n16 9.3005
R1546 VDD1.n19 VDD1.n18 9.3005
R1547 VDD1.n6 VDD1.n5 9.3005
R1548 VDD1.n25 VDD1.n24 9.3005
R1549 VDD1.n27 VDD1.n26 9.3005
R1550 VDD1.n2 VDD1.n1 9.3005
R1551 VDD1.n33 VDD1.n32 9.3005
R1552 VDD1.n45 VDD1.n44 9.3005
R1553 VDD1.n52 VDD1.n51 9.3005
R1554 VDD1.n54 VDD1.n53 9.3005
R1555 VDD1.n41 VDD1.n40 9.3005
R1556 VDD1.n60 VDD1.n59 9.3005
R1557 VDD1.n62 VDD1.n61 9.3005
R1558 VDD1.n37 VDD1.n36 9.3005
R1559 VDD1.n68 VDD1.n67 9.3005
R1560 VDD1.n19 VDD1.n8 8.92171
R1561 VDD1.n54 VDD1.n43 8.92171
R1562 VDD1.n34 VDD1.n0 8.2187
R1563 VDD1.n69 VDD1.n35 8.2187
R1564 VDD1.n16 VDD1.n15 8.14595
R1565 VDD1.n51 VDD1.n50 8.14595
R1566 VDD1.n12 VDD1.n10 7.3702
R1567 VDD1.n47 VDD1.n45 7.3702
R1568 VDD1.n15 VDD1.n10 5.81868
R1569 VDD1.n50 VDD1.n45 5.81868
R1570 VDD1.n32 VDD1.n0 5.3904
R1571 VDD1.n67 VDD1.n35 5.3904
R1572 VDD1.n16 VDD1.n8 5.04292
R1573 VDD1.n51 VDD1.n43 5.04292
R1574 VDD1.n20 VDD1.n19 4.26717
R1575 VDD1.n55 VDD1.n54 4.26717
R1576 VDD1.n23 VDD1.n6 3.49141
R1577 VDD1.n58 VDD1.n41 3.49141
R1578 VDD1.n11 VDD1.n9 2.84305
R1579 VDD1.n46 VDD1.n44 2.84305
R1580 VDD1.n72 VDD1.t3 2.72402
R1581 VDD1.n72 VDD1.t2 2.72402
R1582 VDD1.n70 VDD1.t1 2.72402
R1583 VDD1.n70 VDD1.t0 2.72402
R1584 VDD1.n24 VDD1.n4 2.71565
R1585 VDD1.n59 VDD1.n39 2.71565
R1586 VDD1.n28 VDD1.n27 1.93989
R1587 VDD1.n63 VDD1.n62 1.93989
R1588 VDD1.n31 VDD1.n2 1.16414
R1589 VDD1.n66 VDD1.n37 1.16414
R1590 VDD1 VDD1.n73 0.653517
R1591 VDD1.n33 VDD1.n1 0.155672
R1592 VDD1.n26 VDD1.n1 0.155672
R1593 VDD1.n26 VDD1.n25 0.155672
R1594 VDD1.n25 VDD1.n5 0.155672
R1595 VDD1.n18 VDD1.n5 0.155672
R1596 VDD1.n18 VDD1.n17 0.155672
R1597 VDD1.n17 VDD1.n9 0.155672
R1598 VDD1.n52 VDD1.n44 0.155672
R1599 VDD1.n53 VDD1.n52 0.155672
R1600 VDD1.n53 VDD1.n40 0.155672
R1601 VDD1.n60 VDD1.n40 0.155672
R1602 VDD1.n61 VDD1.n60 0.155672
R1603 VDD1.n61 VDD1.n36 0.155672
R1604 VDD1.n68 VDD1.n36 0.155672
R1605 VTAIL.n146 VTAIL.n116 214.453
R1606 VTAIL.n32 VTAIL.n2 214.453
R1607 VTAIL.n110 VTAIL.n80 214.453
R1608 VTAIL.n72 VTAIL.n42 214.453
R1609 VTAIL.n129 VTAIL.n128 185
R1610 VTAIL.n131 VTAIL.n130 185
R1611 VTAIL.n124 VTAIL.n123 185
R1612 VTAIL.n137 VTAIL.n136 185
R1613 VTAIL.n139 VTAIL.n138 185
R1614 VTAIL.n120 VTAIL.n119 185
R1615 VTAIL.n145 VTAIL.n144 185
R1616 VTAIL.n147 VTAIL.n146 185
R1617 VTAIL.n15 VTAIL.n14 185
R1618 VTAIL.n17 VTAIL.n16 185
R1619 VTAIL.n10 VTAIL.n9 185
R1620 VTAIL.n23 VTAIL.n22 185
R1621 VTAIL.n25 VTAIL.n24 185
R1622 VTAIL.n6 VTAIL.n5 185
R1623 VTAIL.n31 VTAIL.n30 185
R1624 VTAIL.n33 VTAIL.n32 185
R1625 VTAIL.n111 VTAIL.n110 185
R1626 VTAIL.n109 VTAIL.n108 185
R1627 VTAIL.n84 VTAIL.n83 185
R1628 VTAIL.n103 VTAIL.n102 185
R1629 VTAIL.n101 VTAIL.n100 185
R1630 VTAIL.n88 VTAIL.n87 185
R1631 VTAIL.n95 VTAIL.n94 185
R1632 VTAIL.n93 VTAIL.n92 185
R1633 VTAIL.n73 VTAIL.n72 185
R1634 VTAIL.n71 VTAIL.n70 185
R1635 VTAIL.n46 VTAIL.n45 185
R1636 VTAIL.n65 VTAIL.n64 185
R1637 VTAIL.n63 VTAIL.n62 185
R1638 VTAIL.n50 VTAIL.n49 185
R1639 VTAIL.n57 VTAIL.n56 185
R1640 VTAIL.n55 VTAIL.n54 185
R1641 VTAIL.n127 VTAIL.t0 149.524
R1642 VTAIL.n13 VTAIL.t7 149.524
R1643 VTAIL.n91 VTAIL.t5 149.524
R1644 VTAIL.n53 VTAIL.t2 149.524
R1645 VTAIL.n130 VTAIL.n129 104.615
R1646 VTAIL.n130 VTAIL.n123 104.615
R1647 VTAIL.n137 VTAIL.n123 104.615
R1648 VTAIL.n138 VTAIL.n137 104.615
R1649 VTAIL.n138 VTAIL.n119 104.615
R1650 VTAIL.n145 VTAIL.n119 104.615
R1651 VTAIL.n146 VTAIL.n145 104.615
R1652 VTAIL.n16 VTAIL.n15 104.615
R1653 VTAIL.n16 VTAIL.n9 104.615
R1654 VTAIL.n23 VTAIL.n9 104.615
R1655 VTAIL.n24 VTAIL.n23 104.615
R1656 VTAIL.n24 VTAIL.n5 104.615
R1657 VTAIL.n31 VTAIL.n5 104.615
R1658 VTAIL.n32 VTAIL.n31 104.615
R1659 VTAIL.n110 VTAIL.n109 104.615
R1660 VTAIL.n109 VTAIL.n83 104.615
R1661 VTAIL.n102 VTAIL.n83 104.615
R1662 VTAIL.n102 VTAIL.n101 104.615
R1663 VTAIL.n101 VTAIL.n87 104.615
R1664 VTAIL.n94 VTAIL.n87 104.615
R1665 VTAIL.n94 VTAIL.n93 104.615
R1666 VTAIL.n72 VTAIL.n71 104.615
R1667 VTAIL.n71 VTAIL.n45 104.615
R1668 VTAIL.n64 VTAIL.n45 104.615
R1669 VTAIL.n64 VTAIL.n63 104.615
R1670 VTAIL.n63 VTAIL.n49 104.615
R1671 VTAIL.n56 VTAIL.n49 104.615
R1672 VTAIL.n56 VTAIL.n55 104.615
R1673 VTAIL.n129 VTAIL.t0 52.3082
R1674 VTAIL.n15 VTAIL.t7 52.3082
R1675 VTAIL.n93 VTAIL.t5 52.3082
R1676 VTAIL.n55 VTAIL.t2 52.3082
R1677 VTAIL.n79 VTAIL.n78 51.641
R1678 VTAIL.n41 VTAIL.n40 51.641
R1679 VTAIL.n1 VTAIL.n0 51.6408
R1680 VTAIL.n39 VTAIL.n38 51.6408
R1681 VTAIL.n151 VTAIL.n150 35.8702
R1682 VTAIL.n37 VTAIL.n36 35.8702
R1683 VTAIL.n115 VTAIL.n114 35.8702
R1684 VTAIL.n77 VTAIL.n76 35.8702
R1685 VTAIL.n41 VTAIL.n39 24.3238
R1686 VTAIL.n151 VTAIL.n115 21.4789
R1687 VTAIL.n148 VTAIL.n147 12.8005
R1688 VTAIL.n34 VTAIL.n33 12.8005
R1689 VTAIL.n112 VTAIL.n111 12.8005
R1690 VTAIL.n74 VTAIL.n73 12.8005
R1691 VTAIL.n144 VTAIL.n118 12.0247
R1692 VTAIL.n30 VTAIL.n4 12.0247
R1693 VTAIL.n108 VTAIL.n82 12.0247
R1694 VTAIL.n70 VTAIL.n44 12.0247
R1695 VTAIL.n143 VTAIL.n120 11.249
R1696 VTAIL.n29 VTAIL.n6 11.249
R1697 VTAIL.n107 VTAIL.n84 11.249
R1698 VTAIL.n69 VTAIL.n46 11.249
R1699 VTAIL.n140 VTAIL.n139 10.4732
R1700 VTAIL.n26 VTAIL.n25 10.4732
R1701 VTAIL.n104 VTAIL.n103 10.4732
R1702 VTAIL.n66 VTAIL.n65 10.4732
R1703 VTAIL.n128 VTAIL.n127 10.2747
R1704 VTAIL.n14 VTAIL.n13 10.2747
R1705 VTAIL.n92 VTAIL.n91 10.2747
R1706 VTAIL.n54 VTAIL.n53 10.2747
R1707 VTAIL.n136 VTAIL.n122 9.69747
R1708 VTAIL.n22 VTAIL.n8 9.69747
R1709 VTAIL.n100 VTAIL.n86 9.69747
R1710 VTAIL.n62 VTAIL.n48 9.69747
R1711 VTAIL.n150 VTAIL.n149 9.45567
R1712 VTAIL.n36 VTAIL.n35 9.45567
R1713 VTAIL.n114 VTAIL.n113 9.45567
R1714 VTAIL.n76 VTAIL.n75 9.45567
R1715 VTAIL.n126 VTAIL.n125 9.3005
R1716 VTAIL.n133 VTAIL.n132 9.3005
R1717 VTAIL.n135 VTAIL.n134 9.3005
R1718 VTAIL.n122 VTAIL.n121 9.3005
R1719 VTAIL.n141 VTAIL.n140 9.3005
R1720 VTAIL.n143 VTAIL.n142 9.3005
R1721 VTAIL.n118 VTAIL.n117 9.3005
R1722 VTAIL.n149 VTAIL.n148 9.3005
R1723 VTAIL.n12 VTAIL.n11 9.3005
R1724 VTAIL.n19 VTAIL.n18 9.3005
R1725 VTAIL.n21 VTAIL.n20 9.3005
R1726 VTAIL.n8 VTAIL.n7 9.3005
R1727 VTAIL.n27 VTAIL.n26 9.3005
R1728 VTAIL.n29 VTAIL.n28 9.3005
R1729 VTAIL.n4 VTAIL.n3 9.3005
R1730 VTAIL.n35 VTAIL.n34 9.3005
R1731 VTAIL.n90 VTAIL.n89 9.3005
R1732 VTAIL.n97 VTAIL.n96 9.3005
R1733 VTAIL.n99 VTAIL.n98 9.3005
R1734 VTAIL.n86 VTAIL.n85 9.3005
R1735 VTAIL.n105 VTAIL.n104 9.3005
R1736 VTAIL.n107 VTAIL.n106 9.3005
R1737 VTAIL.n82 VTAIL.n81 9.3005
R1738 VTAIL.n113 VTAIL.n112 9.3005
R1739 VTAIL.n52 VTAIL.n51 9.3005
R1740 VTAIL.n59 VTAIL.n58 9.3005
R1741 VTAIL.n61 VTAIL.n60 9.3005
R1742 VTAIL.n48 VTAIL.n47 9.3005
R1743 VTAIL.n67 VTAIL.n66 9.3005
R1744 VTAIL.n69 VTAIL.n68 9.3005
R1745 VTAIL.n44 VTAIL.n43 9.3005
R1746 VTAIL.n75 VTAIL.n74 9.3005
R1747 VTAIL.n135 VTAIL.n124 8.92171
R1748 VTAIL.n21 VTAIL.n10 8.92171
R1749 VTAIL.n99 VTAIL.n88 8.92171
R1750 VTAIL.n61 VTAIL.n50 8.92171
R1751 VTAIL.n150 VTAIL.n116 8.2187
R1752 VTAIL.n36 VTAIL.n2 8.2187
R1753 VTAIL.n114 VTAIL.n80 8.2187
R1754 VTAIL.n76 VTAIL.n42 8.2187
R1755 VTAIL.n132 VTAIL.n131 8.14595
R1756 VTAIL.n18 VTAIL.n17 8.14595
R1757 VTAIL.n96 VTAIL.n95 8.14595
R1758 VTAIL.n58 VTAIL.n57 8.14595
R1759 VTAIL.n128 VTAIL.n126 7.3702
R1760 VTAIL.n14 VTAIL.n12 7.3702
R1761 VTAIL.n92 VTAIL.n90 7.3702
R1762 VTAIL.n54 VTAIL.n52 7.3702
R1763 VTAIL.n131 VTAIL.n126 5.81868
R1764 VTAIL.n17 VTAIL.n12 5.81868
R1765 VTAIL.n95 VTAIL.n90 5.81868
R1766 VTAIL.n57 VTAIL.n52 5.81868
R1767 VTAIL.n148 VTAIL.n116 5.3904
R1768 VTAIL.n34 VTAIL.n2 5.3904
R1769 VTAIL.n112 VTAIL.n80 5.3904
R1770 VTAIL.n74 VTAIL.n42 5.3904
R1771 VTAIL.n132 VTAIL.n124 5.04292
R1772 VTAIL.n18 VTAIL.n10 5.04292
R1773 VTAIL.n96 VTAIL.n88 5.04292
R1774 VTAIL.n58 VTAIL.n50 5.04292
R1775 VTAIL.n136 VTAIL.n135 4.26717
R1776 VTAIL.n22 VTAIL.n21 4.26717
R1777 VTAIL.n100 VTAIL.n99 4.26717
R1778 VTAIL.n62 VTAIL.n61 4.26717
R1779 VTAIL.n139 VTAIL.n122 3.49141
R1780 VTAIL.n25 VTAIL.n8 3.49141
R1781 VTAIL.n103 VTAIL.n86 3.49141
R1782 VTAIL.n65 VTAIL.n48 3.49141
R1783 VTAIL.n77 VTAIL.n41 2.84533
R1784 VTAIL.n115 VTAIL.n79 2.84533
R1785 VTAIL.n39 VTAIL.n37 2.84533
R1786 VTAIL.n127 VTAIL.n125 2.84305
R1787 VTAIL.n13 VTAIL.n11 2.84305
R1788 VTAIL.n91 VTAIL.n89 2.84305
R1789 VTAIL.n53 VTAIL.n51 2.84305
R1790 VTAIL.n0 VTAIL.t11 2.72402
R1791 VTAIL.n0 VTAIL.t1 2.72402
R1792 VTAIL.n38 VTAIL.t6 2.72402
R1793 VTAIL.n38 VTAIL.t10 2.72402
R1794 VTAIL.n78 VTAIL.t8 2.72402
R1795 VTAIL.n78 VTAIL.t9 2.72402
R1796 VTAIL.n40 VTAIL.t4 2.72402
R1797 VTAIL.n40 VTAIL.t3 2.72402
R1798 VTAIL.n140 VTAIL.n120 2.71565
R1799 VTAIL.n26 VTAIL.n6 2.71565
R1800 VTAIL.n104 VTAIL.n84 2.71565
R1801 VTAIL.n66 VTAIL.n46 2.71565
R1802 VTAIL VTAIL.n151 2.07593
R1803 VTAIL.n144 VTAIL.n143 1.93989
R1804 VTAIL.n30 VTAIL.n29 1.93989
R1805 VTAIL.n108 VTAIL.n107 1.93989
R1806 VTAIL.n70 VTAIL.n69 1.93989
R1807 VTAIL.n79 VTAIL.n77 1.89274
R1808 VTAIL.n37 VTAIL.n1 1.89274
R1809 VTAIL.n147 VTAIL.n118 1.16414
R1810 VTAIL.n33 VTAIL.n4 1.16414
R1811 VTAIL.n111 VTAIL.n82 1.16414
R1812 VTAIL.n73 VTAIL.n44 1.16414
R1813 VTAIL VTAIL.n1 0.769897
R1814 VTAIL.n133 VTAIL.n125 0.155672
R1815 VTAIL.n134 VTAIL.n133 0.155672
R1816 VTAIL.n134 VTAIL.n121 0.155672
R1817 VTAIL.n141 VTAIL.n121 0.155672
R1818 VTAIL.n142 VTAIL.n141 0.155672
R1819 VTAIL.n142 VTAIL.n117 0.155672
R1820 VTAIL.n149 VTAIL.n117 0.155672
R1821 VTAIL.n19 VTAIL.n11 0.155672
R1822 VTAIL.n20 VTAIL.n19 0.155672
R1823 VTAIL.n20 VTAIL.n7 0.155672
R1824 VTAIL.n27 VTAIL.n7 0.155672
R1825 VTAIL.n28 VTAIL.n27 0.155672
R1826 VTAIL.n28 VTAIL.n3 0.155672
R1827 VTAIL.n35 VTAIL.n3 0.155672
R1828 VTAIL.n113 VTAIL.n81 0.155672
R1829 VTAIL.n106 VTAIL.n81 0.155672
R1830 VTAIL.n106 VTAIL.n105 0.155672
R1831 VTAIL.n105 VTAIL.n85 0.155672
R1832 VTAIL.n98 VTAIL.n85 0.155672
R1833 VTAIL.n98 VTAIL.n97 0.155672
R1834 VTAIL.n97 VTAIL.n89 0.155672
R1835 VTAIL.n75 VTAIL.n43 0.155672
R1836 VTAIL.n68 VTAIL.n43 0.155672
R1837 VTAIL.n68 VTAIL.n67 0.155672
R1838 VTAIL.n67 VTAIL.n47 0.155672
R1839 VTAIL.n60 VTAIL.n47 0.155672
R1840 VTAIL.n60 VTAIL.n59 0.155672
R1841 VTAIL.n59 VTAIL.n51 0.155672
R1842 VN.n33 VN.n18 161.3
R1843 VN.n32 VN.n31 161.3
R1844 VN.n30 VN.n19 161.3
R1845 VN.n29 VN.n28 161.3
R1846 VN.n27 VN.n20 161.3
R1847 VN.n26 VN.n25 161.3
R1848 VN.n24 VN.n21 161.3
R1849 VN.n15 VN.n0 161.3
R1850 VN.n14 VN.n13 161.3
R1851 VN.n12 VN.n1 161.3
R1852 VN.n11 VN.n10 161.3
R1853 VN.n9 VN.n2 161.3
R1854 VN.n8 VN.n7 161.3
R1855 VN.n6 VN.n3 161.3
R1856 VN.n17 VN.n16 108.309
R1857 VN.n35 VN.n34 108.309
R1858 VN.n5 VN.t3 91.8434
R1859 VN.n23 VN.t4 91.8434
R1860 VN.n5 VN.n4 61.6401
R1861 VN.n23 VN.n22 61.6401
R1862 VN.n4 VN.t2 58.9928
R1863 VN.n16 VN.t5 58.9928
R1864 VN.n22 VN.t1 58.9928
R1865 VN.n34 VN.t0 58.9928
R1866 VN.n10 VN.n9 50.2061
R1867 VN.n28 VN.n27 50.2061
R1868 VN VN.n35 46.8163
R1869 VN.n10 VN.n1 30.7807
R1870 VN.n28 VN.n19 30.7807
R1871 VN.n8 VN.n3 24.4675
R1872 VN.n9 VN.n8 24.4675
R1873 VN.n14 VN.n1 24.4675
R1874 VN.n15 VN.n14 24.4675
R1875 VN.n27 VN.n26 24.4675
R1876 VN.n26 VN.n21 24.4675
R1877 VN.n33 VN.n32 24.4675
R1878 VN.n32 VN.n19 24.4675
R1879 VN.n4 VN.n3 12.234
R1880 VN.n22 VN.n21 12.234
R1881 VN.n24 VN.n23 5.10511
R1882 VN.n6 VN.n5 5.10511
R1883 VN.n16 VN.n15 2.4472
R1884 VN.n34 VN.n33 2.4472
R1885 VN.n35 VN.n18 0.278367
R1886 VN.n17 VN.n0 0.278367
R1887 VN.n31 VN.n18 0.189894
R1888 VN.n31 VN.n30 0.189894
R1889 VN.n30 VN.n29 0.189894
R1890 VN.n29 VN.n20 0.189894
R1891 VN.n25 VN.n20 0.189894
R1892 VN.n25 VN.n24 0.189894
R1893 VN.n7 VN.n6 0.189894
R1894 VN.n7 VN.n2 0.189894
R1895 VN.n11 VN.n2 0.189894
R1896 VN.n12 VN.n11 0.189894
R1897 VN.n13 VN.n12 0.189894
R1898 VN.n13 VN.n0 0.189894
R1899 VN VN.n17 0.153454
R1900 VDD2.n67 VDD2.n37 214.453
R1901 VDD2.n30 VDD2.n0 214.453
R1902 VDD2.n68 VDD2.n67 185
R1903 VDD2.n66 VDD2.n65 185
R1904 VDD2.n41 VDD2.n40 185
R1905 VDD2.n60 VDD2.n59 185
R1906 VDD2.n58 VDD2.n57 185
R1907 VDD2.n45 VDD2.n44 185
R1908 VDD2.n52 VDD2.n51 185
R1909 VDD2.n50 VDD2.n49 185
R1910 VDD2.n13 VDD2.n12 185
R1911 VDD2.n15 VDD2.n14 185
R1912 VDD2.n8 VDD2.n7 185
R1913 VDD2.n21 VDD2.n20 185
R1914 VDD2.n23 VDD2.n22 185
R1915 VDD2.n4 VDD2.n3 185
R1916 VDD2.n29 VDD2.n28 185
R1917 VDD2.n31 VDD2.n30 185
R1918 VDD2.n11 VDD2.t2 149.524
R1919 VDD2.n48 VDD2.t5 149.524
R1920 VDD2.n67 VDD2.n66 104.615
R1921 VDD2.n66 VDD2.n40 104.615
R1922 VDD2.n59 VDD2.n40 104.615
R1923 VDD2.n59 VDD2.n58 104.615
R1924 VDD2.n58 VDD2.n44 104.615
R1925 VDD2.n51 VDD2.n44 104.615
R1926 VDD2.n51 VDD2.n50 104.615
R1927 VDD2.n14 VDD2.n13 104.615
R1928 VDD2.n14 VDD2.n7 104.615
R1929 VDD2.n21 VDD2.n7 104.615
R1930 VDD2.n22 VDD2.n21 104.615
R1931 VDD2.n22 VDD2.n3 104.615
R1932 VDD2.n29 VDD2.n3 104.615
R1933 VDD2.n30 VDD2.n29 104.615
R1934 VDD2.n36 VDD2.n35 68.9755
R1935 VDD2 VDD2.n73 68.9727
R1936 VDD2.n36 VDD2.n34 54.6273
R1937 VDD2.n72 VDD2.n71 52.549
R1938 VDD2.n50 VDD2.t5 52.3082
R1939 VDD2.n13 VDD2.t2 52.3082
R1940 VDD2.n72 VDD2.n36 39.2282
R1941 VDD2.n69 VDD2.n68 12.8005
R1942 VDD2.n32 VDD2.n31 12.8005
R1943 VDD2.n65 VDD2.n39 12.0247
R1944 VDD2.n28 VDD2.n2 12.0247
R1945 VDD2.n64 VDD2.n41 11.249
R1946 VDD2.n27 VDD2.n4 11.249
R1947 VDD2.n61 VDD2.n60 10.4732
R1948 VDD2.n24 VDD2.n23 10.4732
R1949 VDD2.n49 VDD2.n48 10.2747
R1950 VDD2.n12 VDD2.n11 10.2747
R1951 VDD2.n57 VDD2.n43 9.69747
R1952 VDD2.n20 VDD2.n6 9.69747
R1953 VDD2.n71 VDD2.n70 9.45567
R1954 VDD2.n34 VDD2.n33 9.45567
R1955 VDD2.n47 VDD2.n46 9.3005
R1956 VDD2.n54 VDD2.n53 9.3005
R1957 VDD2.n56 VDD2.n55 9.3005
R1958 VDD2.n43 VDD2.n42 9.3005
R1959 VDD2.n62 VDD2.n61 9.3005
R1960 VDD2.n64 VDD2.n63 9.3005
R1961 VDD2.n39 VDD2.n38 9.3005
R1962 VDD2.n70 VDD2.n69 9.3005
R1963 VDD2.n10 VDD2.n9 9.3005
R1964 VDD2.n17 VDD2.n16 9.3005
R1965 VDD2.n19 VDD2.n18 9.3005
R1966 VDD2.n6 VDD2.n5 9.3005
R1967 VDD2.n25 VDD2.n24 9.3005
R1968 VDD2.n27 VDD2.n26 9.3005
R1969 VDD2.n2 VDD2.n1 9.3005
R1970 VDD2.n33 VDD2.n32 9.3005
R1971 VDD2.n56 VDD2.n45 8.92171
R1972 VDD2.n19 VDD2.n8 8.92171
R1973 VDD2.n71 VDD2.n37 8.2187
R1974 VDD2.n34 VDD2.n0 8.2187
R1975 VDD2.n53 VDD2.n52 8.14595
R1976 VDD2.n16 VDD2.n15 8.14595
R1977 VDD2.n49 VDD2.n47 7.3702
R1978 VDD2.n12 VDD2.n10 7.3702
R1979 VDD2.n52 VDD2.n47 5.81868
R1980 VDD2.n15 VDD2.n10 5.81868
R1981 VDD2.n69 VDD2.n37 5.3904
R1982 VDD2.n32 VDD2.n0 5.3904
R1983 VDD2.n53 VDD2.n45 5.04292
R1984 VDD2.n16 VDD2.n8 5.04292
R1985 VDD2.n57 VDD2.n56 4.26717
R1986 VDD2.n20 VDD2.n19 4.26717
R1987 VDD2.n60 VDD2.n43 3.49141
R1988 VDD2.n23 VDD2.n6 3.49141
R1989 VDD2.n48 VDD2.n46 2.84305
R1990 VDD2.n11 VDD2.n9 2.84305
R1991 VDD2.n73 VDD2.t4 2.72402
R1992 VDD2.n73 VDD2.t1 2.72402
R1993 VDD2.n35 VDD2.t3 2.72402
R1994 VDD2.n35 VDD2.t0 2.72402
R1995 VDD2.n61 VDD2.n41 2.71565
R1996 VDD2.n24 VDD2.n4 2.71565
R1997 VDD2 VDD2.n72 2.19231
R1998 VDD2.n65 VDD2.n64 1.93989
R1999 VDD2.n28 VDD2.n27 1.93989
R2000 VDD2.n68 VDD2.n39 1.16414
R2001 VDD2.n31 VDD2.n2 1.16414
R2002 VDD2.n70 VDD2.n38 0.155672
R2003 VDD2.n63 VDD2.n38 0.155672
R2004 VDD2.n63 VDD2.n62 0.155672
R2005 VDD2.n62 VDD2.n42 0.155672
R2006 VDD2.n55 VDD2.n42 0.155672
R2007 VDD2.n55 VDD2.n54 0.155672
R2008 VDD2.n54 VDD2.n46 0.155672
R2009 VDD2.n17 VDD2.n9 0.155672
R2010 VDD2.n18 VDD2.n17 0.155672
R2011 VDD2.n18 VDD2.n5 0.155672
R2012 VDD2.n25 VDD2.n5 0.155672
R2013 VDD2.n26 VDD2.n25 0.155672
R2014 VDD2.n26 VDD2.n1 0.155672
R2015 VDD2.n33 VDD2.n1 0.155672
C0 VTAIL VP 4.80815f
C1 VN VTAIL 4.79395f
C2 VDD1 VDD2 1.55052f
C3 VDD2 VP 0.489311f
C4 VDD1 VP 4.66069f
C5 VN VDD2 4.32496f
C6 VN VDD1 0.151208f
C7 VN VP 6.40835f
C8 VTAIL VDD2 6.24044f
C9 VTAIL VDD1 6.1858f
C10 VDD2 B 5.421488f
C11 VDD1 B 5.582413f
C12 VTAIL B 6.14801f
C13 VN B 13.591811f
C14 VP B 12.297994f
C15 VDD2.n0 B 0.030001f
C16 VDD2.n1 B 0.02156f
C17 VDD2.n2 B 0.011586f
C18 VDD2.n3 B 0.027384f
C19 VDD2.n4 B 0.012267f
C20 VDD2.n5 B 0.02156f
C21 VDD2.n6 B 0.011586f
C22 VDD2.n7 B 0.027384f
C23 VDD2.n8 B 0.012267f
C24 VDD2.n9 B 0.634002f
C25 VDD2.n10 B 0.011586f
C26 VDD2.t2 B 0.045733f
C27 VDD2.n11 B 0.116352f
C28 VDD2.n12 B 0.019358f
C29 VDD2.n13 B 0.020538f
C30 VDD2.n14 B 0.027384f
C31 VDD2.n15 B 0.012267f
C32 VDD2.n16 B 0.011586f
C33 VDD2.n17 B 0.02156f
C34 VDD2.n18 B 0.02156f
C35 VDD2.n19 B 0.011586f
C36 VDD2.n20 B 0.012267f
C37 VDD2.n21 B 0.027384f
C38 VDD2.n22 B 0.027384f
C39 VDD2.n23 B 0.012267f
C40 VDD2.n24 B 0.011586f
C41 VDD2.n25 B 0.02156f
C42 VDD2.n26 B 0.02156f
C43 VDD2.n27 B 0.011586f
C44 VDD2.n28 B 0.012267f
C45 VDD2.n29 B 0.027384f
C46 VDD2.n30 B 0.056561f
C47 VDD2.n31 B 0.012267f
C48 VDD2.n32 B 0.022654f
C49 VDD2.n33 B 0.055432f
C50 VDD2.n34 B 0.081156f
C51 VDD2.t3 B 0.123864f
C52 VDD2.t0 B 0.123864f
C53 VDD2.n35 B 1.06846f
C54 VDD2.n36 B 2.19403f
C55 VDD2.n37 B 0.030001f
C56 VDD2.n38 B 0.02156f
C57 VDD2.n39 B 0.011586f
C58 VDD2.n40 B 0.027384f
C59 VDD2.n41 B 0.012267f
C60 VDD2.n42 B 0.02156f
C61 VDD2.n43 B 0.011586f
C62 VDD2.n44 B 0.027384f
C63 VDD2.n45 B 0.012267f
C64 VDD2.n46 B 0.634002f
C65 VDD2.n47 B 0.011586f
C66 VDD2.t5 B 0.045733f
C67 VDD2.n48 B 0.116352f
C68 VDD2.n49 B 0.019358f
C69 VDD2.n50 B 0.020538f
C70 VDD2.n51 B 0.027384f
C71 VDD2.n52 B 0.012267f
C72 VDD2.n53 B 0.011586f
C73 VDD2.n54 B 0.02156f
C74 VDD2.n55 B 0.02156f
C75 VDD2.n56 B 0.011586f
C76 VDD2.n57 B 0.012267f
C77 VDD2.n58 B 0.027384f
C78 VDD2.n59 B 0.027384f
C79 VDD2.n60 B 0.012267f
C80 VDD2.n61 B 0.011586f
C81 VDD2.n62 B 0.02156f
C82 VDD2.n63 B 0.02156f
C83 VDD2.n64 B 0.011586f
C84 VDD2.n65 B 0.012267f
C85 VDD2.n66 B 0.027384f
C86 VDD2.n67 B 0.056561f
C87 VDD2.n68 B 0.012267f
C88 VDD2.n69 B 0.022654f
C89 VDD2.n70 B 0.055432f
C90 VDD2.n71 B 0.073952f
C91 VDD2.n72 B 1.98163f
C92 VDD2.t4 B 0.123864f
C93 VDD2.t1 B 0.123864f
C94 VDD2.n73 B 1.06844f
C95 VN.n0 B 0.03054f
C96 VN.t5 B 1.33744f
C97 VN.n1 B 0.046407f
C98 VN.n2 B 0.023165f
C99 VN.n3 B 0.032516f
C100 VN.t3 B 1.56942f
C101 VN.t2 B 1.33744f
C102 VN.n4 B 0.561763f
C103 VN.n5 B 0.537782f
C104 VN.n6 B 0.247525f
C105 VN.n7 B 0.023165f
C106 VN.n8 B 0.043173f
C107 VN.n9 B 0.042515f
C108 VN.n10 B 0.021883f
C109 VN.n11 B 0.023165f
C110 VN.n12 B 0.023165f
C111 VN.n13 B 0.023165f
C112 VN.n14 B 0.043173f
C113 VN.n15 B 0.02399f
C114 VN.n16 B 0.567922f
C115 VN.n17 B 0.045017f
C116 VN.n18 B 0.03054f
C117 VN.t0 B 1.33744f
C118 VN.n19 B 0.046407f
C119 VN.n20 B 0.023165f
C120 VN.n21 B 0.032516f
C121 VN.t4 B 1.56942f
C122 VN.t1 B 1.33744f
C123 VN.n22 B 0.561763f
C124 VN.n23 B 0.537782f
C125 VN.n24 B 0.247525f
C126 VN.n25 B 0.023165f
C127 VN.n26 B 0.043173f
C128 VN.n27 B 0.042515f
C129 VN.n28 B 0.021883f
C130 VN.n29 B 0.023165f
C131 VN.n30 B 0.023165f
C132 VN.n31 B 0.023165f
C133 VN.n32 B 0.043173f
C134 VN.n33 B 0.02399f
C135 VN.n34 B 0.567922f
C136 VN.n35 B 1.17806f
C137 VTAIL.t11 B 0.149881f
C138 VTAIL.t1 B 0.149881f
C139 VTAIL.n0 B 1.22359f
C140 VTAIL.n1 B 0.457224f
C141 VTAIL.n2 B 0.036302f
C142 VTAIL.n3 B 0.026089f
C143 VTAIL.n4 B 0.014019f
C144 VTAIL.n5 B 0.033136f
C145 VTAIL.n6 B 0.014844f
C146 VTAIL.n7 B 0.026089f
C147 VTAIL.n8 B 0.014019f
C148 VTAIL.n9 B 0.033136f
C149 VTAIL.n10 B 0.014844f
C150 VTAIL.n11 B 0.76717f
C151 VTAIL.n12 B 0.014019f
C152 VTAIL.t7 B 0.055339f
C153 VTAIL.n13 B 0.140791f
C154 VTAIL.n14 B 0.023425f
C155 VTAIL.n15 B 0.024852f
C156 VTAIL.n16 B 0.033136f
C157 VTAIL.n17 B 0.014844f
C158 VTAIL.n18 B 0.014019f
C159 VTAIL.n19 B 0.026089f
C160 VTAIL.n20 B 0.026089f
C161 VTAIL.n21 B 0.014019f
C162 VTAIL.n22 B 0.014844f
C163 VTAIL.n23 B 0.033136f
C164 VTAIL.n24 B 0.033136f
C165 VTAIL.n25 B 0.014844f
C166 VTAIL.n26 B 0.014019f
C167 VTAIL.n27 B 0.026089f
C168 VTAIL.n28 B 0.026089f
C169 VTAIL.n29 B 0.014019f
C170 VTAIL.n30 B 0.014844f
C171 VTAIL.n31 B 0.033136f
C172 VTAIL.n32 B 0.068442f
C173 VTAIL.n33 B 0.014844f
C174 VTAIL.n34 B 0.027412f
C175 VTAIL.n35 B 0.067075f
C176 VTAIL.n36 B 0.071518f
C177 VTAIL.n37 B 0.424335f
C178 VTAIL.t6 B 0.149881f
C179 VTAIL.t10 B 0.149881f
C180 VTAIL.n38 B 1.22359f
C181 VTAIL.n39 B 1.83217f
C182 VTAIL.t4 B 0.149881f
C183 VTAIL.t3 B 0.149881f
C184 VTAIL.n40 B 1.2236f
C185 VTAIL.n41 B 1.83216f
C186 VTAIL.n42 B 0.036302f
C187 VTAIL.n43 B 0.026089f
C188 VTAIL.n44 B 0.014019f
C189 VTAIL.n45 B 0.033136f
C190 VTAIL.n46 B 0.014844f
C191 VTAIL.n47 B 0.026089f
C192 VTAIL.n48 B 0.014019f
C193 VTAIL.n49 B 0.033136f
C194 VTAIL.n50 B 0.014844f
C195 VTAIL.n51 B 0.76717f
C196 VTAIL.n52 B 0.014019f
C197 VTAIL.t2 B 0.055339f
C198 VTAIL.n53 B 0.140791f
C199 VTAIL.n54 B 0.023425f
C200 VTAIL.n55 B 0.024852f
C201 VTAIL.n56 B 0.033136f
C202 VTAIL.n57 B 0.014844f
C203 VTAIL.n58 B 0.014019f
C204 VTAIL.n59 B 0.026089f
C205 VTAIL.n60 B 0.026089f
C206 VTAIL.n61 B 0.014019f
C207 VTAIL.n62 B 0.014844f
C208 VTAIL.n63 B 0.033136f
C209 VTAIL.n64 B 0.033136f
C210 VTAIL.n65 B 0.014844f
C211 VTAIL.n66 B 0.014019f
C212 VTAIL.n67 B 0.026089f
C213 VTAIL.n68 B 0.026089f
C214 VTAIL.n69 B 0.014019f
C215 VTAIL.n70 B 0.014844f
C216 VTAIL.n71 B 0.033136f
C217 VTAIL.n72 B 0.068442f
C218 VTAIL.n73 B 0.014844f
C219 VTAIL.n74 B 0.027412f
C220 VTAIL.n75 B 0.067075f
C221 VTAIL.n76 B 0.071518f
C222 VTAIL.n77 B 0.424335f
C223 VTAIL.t8 B 0.149881f
C224 VTAIL.t9 B 0.149881f
C225 VTAIL.n78 B 1.2236f
C226 VTAIL.n79 B 0.631687f
C227 VTAIL.n80 B 0.036302f
C228 VTAIL.n81 B 0.026089f
C229 VTAIL.n82 B 0.014019f
C230 VTAIL.n83 B 0.033136f
C231 VTAIL.n84 B 0.014844f
C232 VTAIL.n85 B 0.026089f
C233 VTAIL.n86 B 0.014019f
C234 VTAIL.n87 B 0.033136f
C235 VTAIL.n88 B 0.014844f
C236 VTAIL.n89 B 0.76717f
C237 VTAIL.n90 B 0.014019f
C238 VTAIL.t5 B 0.055339f
C239 VTAIL.n91 B 0.140791f
C240 VTAIL.n92 B 0.023425f
C241 VTAIL.n93 B 0.024852f
C242 VTAIL.n94 B 0.033136f
C243 VTAIL.n95 B 0.014844f
C244 VTAIL.n96 B 0.014019f
C245 VTAIL.n97 B 0.026089f
C246 VTAIL.n98 B 0.026089f
C247 VTAIL.n99 B 0.014019f
C248 VTAIL.n100 B 0.014844f
C249 VTAIL.n101 B 0.033136f
C250 VTAIL.n102 B 0.033136f
C251 VTAIL.n103 B 0.014844f
C252 VTAIL.n104 B 0.014019f
C253 VTAIL.n105 B 0.026089f
C254 VTAIL.n106 B 0.026089f
C255 VTAIL.n107 B 0.014019f
C256 VTAIL.n108 B 0.014844f
C257 VTAIL.n109 B 0.033136f
C258 VTAIL.n110 B 0.068442f
C259 VTAIL.n111 B 0.014844f
C260 VTAIL.n112 B 0.027412f
C261 VTAIL.n113 B 0.067075f
C262 VTAIL.n114 B 0.071518f
C263 VTAIL.n115 B 1.38566f
C264 VTAIL.n116 B 0.036302f
C265 VTAIL.n117 B 0.026089f
C266 VTAIL.n118 B 0.014019f
C267 VTAIL.n119 B 0.033136f
C268 VTAIL.n120 B 0.014844f
C269 VTAIL.n121 B 0.026089f
C270 VTAIL.n122 B 0.014019f
C271 VTAIL.n123 B 0.033136f
C272 VTAIL.n124 B 0.014844f
C273 VTAIL.n125 B 0.76717f
C274 VTAIL.n126 B 0.014019f
C275 VTAIL.t0 B 0.055339f
C276 VTAIL.n127 B 0.140791f
C277 VTAIL.n128 B 0.023425f
C278 VTAIL.n129 B 0.024852f
C279 VTAIL.n130 B 0.033136f
C280 VTAIL.n131 B 0.014844f
C281 VTAIL.n132 B 0.014019f
C282 VTAIL.n133 B 0.026089f
C283 VTAIL.n134 B 0.026089f
C284 VTAIL.n135 B 0.014019f
C285 VTAIL.n136 B 0.014844f
C286 VTAIL.n137 B 0.033136f
C287 VTAIL.n138 B 0.033136f
C288 VTAIL.n139 B 0.014844f
C289 VTAIL.n140 B 0.014019f
C290 VTAIL.n141 B 0.026089f
C291 VTAIL.n142 B 0.026089f
C292 VTAIL.n143 B 0.014019f
C293 VTAIL.n144 B 0.014844f
C294 VTAIL.n145 B 0.033136f
C295 VTAIL.n146 B 0.068442f
C296 VTAIL.n147 B 0.014844f
C297 VTAIL.n148 B 0.027412f
C298 VTAIL.n149 B 0.067075f
C299 VTAIL.n150 B 0.071518f
C300 VTAIL.n151 B 1.32098f
C301 VDD1.n0 B 0.030909f
C302 VDD1.n1 B 0.022213f
C303 VDD1.n2 B 0.011936f
C304 VDD1.n3 B 0.028213f
C305 VDD1.n4 B 0.012639f
C306 VDD1.n5 B 0.022213f
C307 VDD1.n6 B 0.011936f
C308 VDD1.n7 B 0.028213f
C309 VDD1.n8 B 0.012639f
C310 VDD1.n9 B 0.6532f
C311 VDD1.n10 B 0.011936f
C312 VDD1.t5 B 0.047118f
C313 VDD1.n11 B 0.119876f
C314 VDD1.n12 B 0.019945f
C315 VDD1.n13 B 0.02116f
C316 VDD1.n14 B 0.028213f
C317 VDD1.n15 B 0.012639f
C318 VDD1.n16 B 0.011936f
C319 VDD1.n17 B 0.022213f
C320 VDD1.n18 B 0.022213f
C321 VDD1.n19 B 0.011936f
C322 VDD1.n20 B 0.012639f
C323 VDD1.n21 B 0.028213f
C324 VDD1.n22 B 0.028213f
C325 VDD1.n23 B 0.012639f
C326 VDD1.n24 B 0.011936f
C327 VDD1.n25 B 0.022213f
C328 VDD1.n26 B 0.022213f
C329 VDD1.n27 B 0.011936f
C330 VDD1.n28 B 0.012639f
C331 VDD1.n29 B 0.028213f
C332 VDD1.n30 B 0.058274f
C333 VDD1.n31 B 0.012639f
C334 VDD1.n32 B 0.02334f
C335 VDD1.n33 B 0.057111f
C336 VDD1.n34 B 0.084318f
C337 VDD1.n35 B 0.030909f
C338 VDD1.n36 B 0.022213f
C339 VDD1.n37 B 0.011936f
C340 VDD1.n38 B 0.028213f
C341 VDD1.n39 B 0.012639f
C342 VDD1.n40 B 0.022213f
C343 VDD1.n41 B 0.011936f
C344 VDD1.n42 B 0.028213f
C345 VDD1.n43 B 0.012639f
C346 VDD1.n44 B 0.6532f
C347 VDD1.n45 B 0.011936f
C348 VDD1.t4 B 0.047118f
C349 VDD1.n46 B 0.119876f
C350 VDD1.n47 B 0.019945f
C351 VDD1.n48 B 0.02116f
C352 VDD1.n49 B 0.028213f
C353 VDD1.n50 B 0.012639f
C354 VDD1.n51 B 0.011936f
C355 VDD1.n52 B 0.022213f
C356 VDD1.n53 B 0.022213f
C357 VDD1.n54 B 0.011936f
C358 VDD1.n55 B 0.012639f
C359 VDD1.n56 B 0.028213f
C360 VDD1.n57 B 0.028213f
C361 VDD1.n58 B 0.012639f
C362 VDD1.n59 B 0.011936f
C363 VDD1.n60 B 0.022213f
C364 VDD1.n61 B 0.022213f
C365 VDD1.n62 B 0.011936f
C366 VDD1.n63 B 0.012639f
C367 VDD1.n64 B 0.028213f
C368 VDD1.n65 B 0.058274f
C369 VDD1.n66 B 0.012639f
C370 VDD1.n67 B 0.02334f
C371 VDD1.n68 B 0.057111f
C372 VDD1.n69 B 0.083613f
C373 VDD1.t1 B 0.127615f
C374 VDD1.t0 B 0.127615f
C375 VDD1.n70 B 1.10082f
C376 VDD1.n71 B 2.37537f
C377 VDD1.t3 B 0.127615f
C378 VDD1.t2 B 0.127615f
C379 VDD1.n72 B 1.09669f
C380 VDD1.n73 B 2.23925f
C381 VP.n0 B 0.031394f
C382 VP.t3 B 1.37484f
C383 VP.n1 B 0.047705f
C384 VP.n2 B 0.023812f
C385 VP.n3 B 0.033425f
C386 VP.n4 B 0.023812f
C387 VP.n5 B 0.022495f
C388 VP.n6 B 0.023812f
C389 VP.t4 B 1.37484f
C390 VP.n7 B 0.583804f
C391 VP.n8 B 0.031394f
C392 VP.t5 B 1.37484f
C393 VP.n9 B 0.047705f
C394 VP.n10 B 0.023812f
C395 VP.n11 B 0.033425f
C396 VP.t2 B 1.61331f
C397 VP.t1 B 1.37484f
C398 VP.n12 B 0.577473f
C399 VP.n13 B 0.552821f
C400 VP.n14 B 0.254448f
C401 VP.n15 B 0.023812f
C402 VP.n16 B 0.04438f
C403 VP.n17 B 0.043704f
C404 VP.n18 B 0.022495f
C405 VP.n19 B 0.023812f
C406 VP.n20 B 0.023812f
C407 VP.n21 B 0.023812f
C408 VP.n22 B 0.04438f
C409 VP.n23 B 0.024661f
C410 VP.n24 B 0.583804f
C411 VP.n25 B 1.19806f
C412 VP.n26 B 1.21645f
C413 VP.n27 B 0.031394f
C414 VP.n28 B 0.024661f
C415 VP.n29 B 0.04438f
C416 VP.n30 B 0.047705f
C417 VP.n31 B 0.023812f
C418 VP.n32 B 0.023812f
C419 VP.n33 B 0.023812f
C420 VP.n34 B 0.043704f
C421 VP.n35 B 0.04438f
C422 VP.t0 B 1.37484f
C423 VP.n36 B 0.502213f
C424 VP.n37 B 0.033425f
C425 VP.n38 B 0.023812f
C426 VP.n39 B 0.023812f
C427 VP.n40 B 0.023812f
C428 VP.n41 B 0.04438f
C429 VP.n42 B 0.043704f
C430 VP.n43 B 0.022495f
C431 VP.n44 B 0.023812f
C432 VP.n45 B 0.023812f
C433 VP.n46 B 0.023812f
C434 VP.n47 B 0.04438f
C435 VP.n48 B 0.024661f
C436 VP.n49 B 0.583804f
C437 VP.n50 B 0.046276f
.ends

