* NGSPICE file created from diff_pair_sample_1088.ext - technology: sky130A

.subckt diff_pair_sample_1088 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.58885 pd=16.02 as=2.58885 ps=16.02 w=15.69 l=3.15
X1 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=6.1191 pd=32.16 as=0 ps=0 w=15.69 l=3.15
X2 VTAIL.t5 VN.t0 VDD2.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=6.1191 pd=32.16 as=2.58885 ps=16.02 w=15.69 l=3.15
X3 VDD1.t0 VP.t1 VTAIL.t14 B.t2 sky130_fd_pr__nfet_01v8 ad=2.58885 pd=16.02 as=2.58885 ps=16.02 w=15.69 l=3.15
X4 VDD2.t6 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.58885 pd=16.02 as=2.58885 ps=16.02 w=15.69 l=3.15
X5 VTAIL.t13 VP.t2 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=6.1191 pd=32.16 as=2.58885 ps=16.02 w=15.69 l=3.15
X6 VDD1.t4 VP.t3 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=2.58885 pd=16.02 as=6.1191 ps=32.16 w=15.69 l=3.15
X7 VDD2.t5 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.58885 pd=16.02 as=2.58885 ps=16.02 w=15.69 l=3.15
X8 VTAIL.t11 VP.t4 VDD1.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=2.58885 pd=16.02 as=2.58885 ps=16.02 w=15.69 l=3.15
X9 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=6.1191 pd=32.16 as=0 ps=0 w=15.69 l=3.15
X10 VDD1.t6 VP.t5 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=2.58885 pd=16.02 as=6.1191 ps=32.16 w=15.69 l=3.15
X11 VDD2.t4 VN.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.58885 pd=16.02 as=6.1191 ps=32.16 w=15.69 l=3.15
X12 VTAIL.t1 VN.t4 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=6.1191 pd=32.16 as=2.58885 ps=16.02 w=15.69 l=3.15
X13 VDD2.t2 VN.t5 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.58885 pd=16.02 as=6.1191 ps=32.16 w=15.69 l=3.15
X14 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=6.1191 pd=32.16 as=0 ps=0 w=15.69 l=3.15
X15 VDD1.t3 VP.t6 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=2.58885 pd=16.02 as=2.58885 ps=16.02 w=15.69 l=3.15
X16 VTAIL.t0 VN.t6 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.58885 pd=16.02 as=2.58885 ps=16.02 w=15.69 l=3.15
X17 VTAIL.t4 VN.t7 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=2.58885 pd=16.02 as=2.58885 ps=16.02 w=15.69 l=3.15
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.1191 pd=32.16 as=0 ps=0 w=15.69 l=3.15
X19 VTAIL.t8 VP.t7 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=6.1191 pd=32.16 as=2.58885 ps=16.02 w=15.69 l=3.15
R0 VP.n21 VP.n18 161.3
R1 VP.n23 VP.n22 161.3
R2 VP.n24 VP.n17 161.3
R3 VP.n26 VP.n25 161.3
R4 VP.n27 VP.n16 161.3
R5 VP.n29 VP.n28 161.3
R6 VP.n31 VP.n30 161.3
R7 VP.n32 VP.n14 161.3
R8 VP.n34 VP.n33 161.3
R9 VP.n35 VP.n13 161.3
R10 VP.n37 VP.n36 161.3
R11 VP.n38 VP.n12 161.3
R12 VP.n40 VP.n39 161.3
R13 VP.n75 VP.n74 161.3
R14 VP.n73 VP.n1 161.3
R15 VP.n72 VP.n71 161.3
R16 VP.n70 VP.n2 161.3
R17 VP.n69 VP.n68 161.3
R18 VP.n67 VP.n3 161.3
R19 VP.n66 VP.n65 161.3
R20 VP.n64 VP.n63 161.3
R21 VP.n62 VP.n5 161.3
R22 VP.n61 VP.n60 161.3
R23 VP.n59 VP.n6 161.3
R24 VP.n58 VP.n57 161.3
R25 VP.n56 VP.n7 161.3
R26 VP.n54 VP.n53 161.3
R27 VP.n52 VP.n8 161.3
R28 VP.n51 VP.n50 161.3
R29 VP.n49 VP.n9 161.3
R30 VP.n48 VP.n47 161.3
R31 VP.n46 VP.n10 161.3
R32 VP.n45 VP.n44 161.3
R33 VP.n19 VP.t7 153.446
R34 VP.n43 VP.t2 120.041
R35 VP.n55 VP.t6 120.041
R36 VP.n4 VP.t4 120.041
R37 VP.n0 VP.t5 120.041
R38 VP.n11 VP.t3 120.041
R39 VP.n15 VP.t0 120.041
R40 VP.n20 VP.t1 120.041
R41 VP.n43 VP.n42 67.0684
R42 VP.n76 VP.n0 67.0684
R43 VP.n41 VP.n11 67.0684
R44 VP.n49 VP.n48 56.5193
R45 VP.n61 VP.n6 56.5193
R46 VP.n72 VP.n2 56.5193
R47 VP.n37 VP.n13 56.5193
R48 VP.n26 VP.n17 56.5193
R49 VP.n42 VP.n41 56.469
R50 VP.n20 VP.n19 50.0328
R51 VP.n44 VP.n10 24.4675
R52 VP.n48 VP.n10 24.4675
R53 VP.n50 VP.n49 24.4675
R54 VP.n50 VP.n8 24.4675
R55 VP.n54 VP.n8 24.4675
R56 VP.n57 VP.n56 24.4675
R57 VP.n57 VP.n6 24.4675
R58 VP.n62 VP.n61 24.4675
R59 VP.n63 VP.n62 24.4675
R60 VP.n67 VP.n66 24.4675
R61 VP.n68 VP.n67 24.4675
R62 VP.n68 VP.n2 24.4675
R63 VP.n73 VP.n72 24.4675
R64 VP.n74 VP.n73 24.4675
R65 VP.n38 VP.n37 24.4675
R66 VP.n39 VP.n38 24.4675
R67 VP.n27 VP.n26 24.4675
R68 VP.n28 VP.n27 24.4675
R69 VP.n32 VP.n31 24.4675
R70 VP.n33 VP.n32 24.4675
R71 VP.n33 VP.n13 24.4675
R72 VP.n22 VP.n21 24.4675
R73 VP.n22 VP.n17 24.4675
R74 VP.n56 VP.n55 23.9782
R75 VP.n63 VP.n4 23.9782
R76 VP.n28 VP.n15 23.9782
R77 VP.n21 VP.n20 23.9782
R78 VP.n44 VP.n43 22.9995
R79 VP.n74 VP.n0 22.9995
R80 VP.n39 VP.n11 22.9995
R81 VP.n19 VP.n18 3.77028
R82 VP.n55 VP.n54 0.48984
R83 VP.n66 VP.n4 0.48984
R84 VP.n31 VP.n15 0.48984
R85 VP.n41 VP.n40 0.354971
R86 VP.n45 VP.n42 0.354971
R87 VP.n76 VP.n75 0.354971
R88 VP VP.n76 0.26696
R89 VP.n23 VP.n18 0.189894
R90 VP.n24 VP.n23 0.189894
R91 VP.n25 VP.n24 0.189894
R92 VP.n25 VP.n16 0.189894
R93 VP.n29 VP.n16 0.189894
R94 VP.n30 VP.n29 0.189894
R95 VP.n30 VP.n14 0.189894
R96 VP.n34 VP.n14 0.189894
R97 VP.n35 VP.n34 0.189894
R98 VP.n36 VP.n35 0.189894
R99 VP.n36 VP.n12 0.189894
R100 VP.n40 VP.n12 0.189894
R101 VP.n46 VP.n45 0.189894
R102 VP.n47 VP.n46 0.189894
R103 VP.n47 VP.n9 0.189894
R104 VP.n51 VP.n9 0.189894
R105 VP.n52 VP.n51 0.189894
R106 VP.n53 VP.n52 0.189894
R107 VP.n53 VP.n7 0.189894
R108 VP.n58 VP.n7 0.189894
R109 VP.n59 VP.n58 0.189894
R110 VP.n60 VP.n59 0.189894
R111 VP.n60 VP.n5 0.189894
R112 VP.n64 VP.n5 0.189894
R113 VP.n65 VP.n64 0.189894
R114 VP.n65 VP.n3 0.189894
R115 VP.n69 VP.n3 0.189894
R116 VP.n70 VP.n69 0.189894
R117 VP.n71 VP.n70 0.189894
R118 VP.n71 VP.n1 0.189894
R119 VP.n75 VP.n1 0.189894
R120 VDD1 VDD1.n0 61.7847
R121 VDD1.n3 VDD1.n2 61.6709
R122 VDD1.n3 VDD1.n1 61.6709
R123 VDD1.n5 VDD1.n4 60.2263
R124 VDD1.n5 VDD1.n3 51.3242
R125 VDD1 VDD1.n5 1.44231
R126 VDD1.n4 VDD1.t1 1.26245
R127 VDD1.n4 VDD1.t4 1.26245
R128 VDD1.n0 VDD1.t2 1.26245
R129 VDD1.n0 VDD1.t0 1.26245
R130 VDD1.n2 VDD1.t7 1.26245
R131 VDD1.n2 VDD1.t6 1.26245
R132 VDD1.n1 VDD1.t5 1.26245
R133 VDD1.n1 VDD1.t3 1.26245
R134 VTAIL.n11 VTAIL.t8 44.8096
R135 VTAIL.n10 VTAIL.t6 44.8096
R136 VTAIL.n7 VTAIL.t5 44.8096
R137 VTAIL.n15 VTAIL.t7 44.8095
R138 VTAIL.n2 VTAIL.t1 44.8095
R139 VTAIL.n3 VTAIL.t10 44.8095
R140 VTAIL.n6 VTAIL.t13 44.8095
R141 VTAIL.n14 VTAIL.t12 44.8095
R142 VTAIL.n13 VTAIL.n12 43.5477
R143 VTAIL.n9 VTAIL.n8 43.5477
R144 VTAIL.n1 VTAIL.n0 43.5474
R145 VTAIL.n5 VTAIL.n4 43.5474
R146 VTAIL.n15 VTAIL.n14 28.8927
R147 VTAIL.n7 VTAIL.n6 28.8927
R148 VTAIL.n9 VTAIL.n7 3.0005
R149 VTAIL.n10 VTAIL.n9 3.0005
R150 VTAIL.n13 VTAIL.n11 3.0005
R151 VTAIL.n14 VTAIL.n13 3.0005
R152 VTAIL.n6 VTAIL.n5 3.0005
R153 VTAIL.n5 VTAIL.n3 3.0005
R154 VTAIL.n2 VTAIL.n1 3.0005
R155 VTAIL VTAIL.n15 2.94231
R156 VTAIL.n0 VTAIL.t2 1.26245
R157 VTAIL.n0 VTAIL.t4 1.26245
R158 VTAIL.n4 VTAIL.t9 1.26245
R159 VTAIL.n4 VTAIL.t11 1.26245
R160 VTAIL.n12 VTAIL.t14 1.26245
R161 VTAIL.n12 VTAIL.t15 1.26245
R162 VTAIL.n8 VTAIL.t3 1.26245
R163 VTAIL.n8 VTAIL.t0 1.26245
R164 VTAIL.n11 VTAIL.n10 0.470328
R165 VTAIL.n3 VTAIL.n2 0.470328
R166 VTAIL VTAIL.n1 0.0586897
R167 B.n1055 B.n1054 585
R168 B.n394 B.n166 585
R169 B.n393 B.n392 585
R170 B.n391 B.n390 585
R171 B.n389 B.n388 585
R172 B.n387 B.n386 585
R173 B.n385 B.n384 585
R174 B.n383 B.n382 585
R175 B.n381 B.n380 585
R176 B.n379 B.n378 585
R177 B.n377 B.n376 585
R178 B.n375 B.n374 585
R179 B.n373 B.n372 585
R180 B.n371 B.n370 585
R181 B.n369 B.n368 585
R182 B.n367 B.n366 585
R183 B.n365 B.n364 585
R184 B.n363 B.n362 585
R185 B.n361 B.n360 585
R186 B.n359 B.n358 585
R187 B.n357 B.n356 585
R188 B.n355 B.n354 585
R189 B.n353 B.n352 585
R190 B.n351 B.n350 585
R191 B.n349 B.n348 585
R192 B.n347 B.n346 585
R193 B.n345 B.n344 585
R194 B.n343 B.n342 585
R195 B.n341 B.n340 585
R196 B.n339 B.n338 585
R197 B.n337 B.n336 585
R198 B.n335 B.n334 585
R199 B.n333 B.n332 585
R200 B.n331 B.n330 585
R201 B.n329 B.n328 585
R202 B.n327 B.n326 585
R203 B.n325 B.n324 585
R204 B.n323 B.n322 585
R205 B.n321 B.n320 585
R206 B.n319 B.n318 585
R207 B.n317 B.n316 585
R208 B.n315 B.n314 585
R209 B.n313 B.n312 585
R210 B.n311 B.n310 585
R211 B.n309 B.n308 585
R212 B.n307 B.n306 585
R213 B.n305 B.n304 585
R214 B.n303 B.n302 585
R215 B.n301 B.n300 585
R216 B.n299 B.n298 585
R217 B.n297 B.n296 585
R218 B.n295 B.n294 585
R219 B.n293 B.n292 585
R220 B.n291 B.n290 585
R221 B.n289 B.n288 585
R222 B.n287 B.n286 585
R223 B.n285 B.n284 585
R224 B.n283 B.n282 585
R225 B.n281 B.n280 585
R226 B.n279 B.n278 585
R227 B.n277 B.n276 585
R228 B.n275 B.n274 585
R229 B.n273 B.n272 585
R230 B.n271 B.n270 585
R231 B.n269 B.n268 585
R232 B.n267 B.n266 585
R233 B.n265 B.n264 585
R234 B.n263 B.n262 585
R235 B.n261 B.n260 585
R236 B.n259 B.n258 585
R237 B.n257 B.n256 585
R238 B.n255 B.n254 585
R239 B.n253 B.n252 585
R240 B.n251 B.n250 585
R241 B.n249 B.n248 585
R242 B.n247 B.n246 585
R243 B.n245 B.n244 585
R244 B.n243 B.n242 585
R245 B.n241 B.n240 585
R246 B.n239 B.n238 585
R247 B.n237 B.n236 585
R248 B.n235 B.n234 585
R249 B.n233 B.n232 585
R250 B.n231 B.n230 585
R251 B.n229 B.n228 585
R252 B.n227 B.n226 585
R253 B.n225 B.n224 585
R254 B.n223 B.n222 585
R255 B.n221 B.n220 585
R256 B.n219 B.n218 585
R257 B.n217 B.n216 585
R258 B.n215 B.n214 585
R259 B.n213 B.n212 585
R260 B.n211 B.n210 585
R261 B.n209 B.n208 585
R262 B.n207 B.n206 585
R263 B.n205 B.n204 585
R264 B.n203 B.n202 585
R265 B.n201 B.n200 585
R266 B.n199 B.n198 585
R267 B.n197 B.n196 585
R268 B.n195 B.n194 585
R269 B.n193 B.n192 585
R270 B.n191 B.n190 585
R271 B.n189 B.n188 585
R272 B.n187 B.n186 585
R273 B.n185 B.n184 585
R274 B.n183 B.n182 585
R275 B.n181 B.n180 585
R276 B.n179 B.n178 585
R277 B.n177 B.n176 585
R278 B.n175 B.n174 585
R279 B.n110 B.n109 585
R280 B.n1060 B.n1059 585
R281 B.n1053 B.n167 585
R282 B.n167 B.n107 585
R283 B.n1052 B.n106 585
R284 B.n1064 B.n106 585
R285 B.n1051 B.n105 585
R286 B.n1065 B.n105 585
R287 B.n1050 B.n104 585
R288 B.n1066 B.n104 585
R289 B.n1049 B.n1048 585
R290 B.n1048 B.n100 585
R291 B.n1047 B.n99 585
R292 B.n1072 B.n99 585
R293 B.n1046 B.n98 585
R294 B.n1073 B.n98 585
R295 B.n1045 B.n97 585
R296 B.n1074 B.n97 585
R297 B.n1044 B.n1043 585
R298 B.n1043 B.n96 585
R299 B.n1042 B.n92 585
R300 B.n1080 B.n92 585
R301 B.n1041 B.n91 585
R302 B.n1081 B.n91 585
R303 B.n1040 B.n90 585
R304 B.n1082 B.n90 585
R305 B.n1039 B.n1038 585
R306 B.n1038 B.n86 585
R307 B.n1037 B.n85 585
R308 B.n1088 B.n85 585
R309 B.n1036 B.n84 585
R310 B.n1089 B.n84 585
R311 B.n1035 B.n83 585
R312 B.n1090 B.n83 585
R313 B.n1034 B.n1033 585
R314 B.n1033 B.n79 585
R315 B.n1032 B.n78 585
R316 B.n1096 B.n78 585
R317 B.n1031 B.n77 585
R318 B.n1097 B.n77 585
R319 B.n1030 B.n76 585
R320 B.n1098 B.n76 585
R321 B.n1029 B.n1028 585
R322 B.n1028 B.n72 585
R323 B.n1027 B.n71 585
R324 B.n1104 B.n71 585
R325 B.n1026 B.n70 585
R326 B.n1105 B.n70 585
R327 B.n1025 B.n69 585
R328 B.n1106 B.n69 585
R329 B.n1024 B.n1023 585
R330 B.n1023 B.n65 585
R331 B.n1022 B.n64 585
R332 B.n1112 B.n64 585
R333 B.n1021 B.n63 585
R334 B.n1113 B.n63 585
R335 B.n1020 B.n62 585
R336 B.n1114 B.n62 585
R337 B.n1019 B.n1018 585
R338 B.n1018 B.n58 585
R339 B.n1017 B.n57 585
R340 B.n1120 B.n57 585
R341 B.n1016 B.n56 585
R342 B.n1121 B.n56 585
R343 B.n1015 B.n55 585
R344 B.n1122 B.n55 585
R345 B.n1014 B.n1013 585
R346 B.n1013 B.n54 585
R347 B.n1012 B.n50 585
R348 B.n1128 B.n50 585
R349 B.n1011 B.n49 585
R350 B.n1129 B.n49 585
R351 B.n1010 B.n48 585
R352 B.n1130 B.n48 585
R353 B.n1009 B.n1008 585
R354 B.n1008 B.n44 585
R355 B.n1007 B.n43 585
R356 B.n1136 B.n43 585
R357 B.n1006 B.n42 585
R358 B.n1137 B.n42 585
R359 B.n1005 B.n41 585
R360 B.n1138 B.n41 585
R361 B.n1004 B.n1003 585
R362 B.n1003 B.n37 585
R363 B.n1002 B.n36 585
R364 B.n1144 B.n36 585
R365 B.n1001 B.n35 585
R366 B.n1145 B.n35 585
R367 B.n1000 B.n34 585
R368 B.n1146 B.n34 585
R369 B.n999 B.n998 585
R370 B.n998 B.n30 585
R371 B.n997 B.n29 585
R372 B.n1152 B.n29 585
R373 B.n996 B.n28 585
R374 B.n1153 B.n28 585
R375 B.n995 B.n27 585
R376 B.n1154 B.n27 585
R377 B.n994 B.n993 585
R378 B.n993 B.n23 585
R379 B.n992 B.n22 585
R380 B.n1160 B.n22 585
R381 B.n991 B.n21 585
R382 B.n1161 B.n21 585
R383 B.n990 B.n20 585
R384 B.n1162 B.n20 585
R385 B.n989 B.n988 585
R386 B.n988 B.n19 585
R387 B.n987 B.n15 585
R388 B.n1168 B.n15 585
R389 B.n986 B.n14 585
R390 B.n1169 B.n14 585
R391 B.n985 B.n13 585
R392 B.n1170 B.n13 585
R393 B.n984 B.n983 585
R394 B.n983 B.n12 585
R395 B.n982 B.n981 585
R396 B.n982 B.n8 585
R397 B.n980 B.n7 585
R398 B.n1177 B.n7 585
R399 B.n979 B.n6 585
R400 B.n1178 B.n6 585
R401 B.n978 B.n5 585
R402 B.n1179 B.n5 585
R403 B.n977 B.n976 585
R404 B.n976 B.n4 585
R405 B.n975 B.n395 585
R406 B.n975 B.n974 585
R407 B.n965 B.n396 585
R408 B.n397 B.n396 585
R409 B.n967 B.n966 585
R410 B.n968 B.n967 585
R411 B.n964 B.n402 585
R412 B.n402 B.n401 585
R413 B.n963 B.n962 585
R414 B.n962 B.n961 585
R415 B.n404 B.n403 585
R416 B.n954 B.n404 585
R417 B.n953 B.n952 585
R418 B.n955 B.n953 585
R419 B.n951 B.n409 585
R420 B.n409 B.n408 585
R421 B.n950 B.n949 585
R422 B.n949 B.n948 585
R423 B.n411 B.n410 585
R424 B.n412 B.n411 585
R425 B.n941 B.n940 585
R426 B.n942 B.n941 585
R427 B.n939 B.n417 585
R428 B.n417 B.n416 585
R429 B.n938 B.n937 585
R430 B.n937 B.n936 585
R431 B.n419 B.n418 585
R432 B.n420 B.n419 585
R433 B.n929 B.n928 585
R434 B.n930 B.n929 585
R435 B.n927 B.n424 585
R436 B.n428 B.n424 585
R437 B.n926 B.n925 585
R438 B.n925 B.n924 585
R439 B.n426 B.n425 585
R440 B.n427 B.n426 585
R441 B.n917 B.n916 585
R442 B.n918 B.n917 585
R443 B.n915 B.n433 585
R444 B.n433 B.n432 585
R445 B.n914 B.n913 585
R446 B.n913 B.n912 585
R447 B.n435 B.n434 585
R448 B.n436 B.n435 585
R449 B.n905 B.n904 585
R450 B.n906 B.n905 585
R451 B.n903 B.n441 585
R452 B.n441 B.n440 585
R453 B.n902 B.n901 585
R454 B.n901 B.n900 585
R455 B.n443 B.n442 585
R456 B.n893 B.n443 585
R457 B.n892 B.n891 585
R458 B.n894 B.n892 585
R459 B.n890 B.n448 585
R460 B.n448 B.n447 585
R461 B.n889 B.n888 585
R462 B.n888 B.n887 585
R463 B.n450 B.n449 585
R464 B.n451 B.n450 585
R465 B.n880 B.n879 585
R466 B.n881 B.n880 585
R467 B.n878 B.n456 585
R468 B.n456 B.n455 585
R469 B.n877 B.n876 585
R470 B.n876 B.n875 585
R471 B.n458 B.n457 585
R472 B.n459 B.n458 585
R473 B.n868 B.n867 585
R474 B.n869 B.n868 585
R475 B.n866 B.n463 585
R476 B.n467 B.n463 585
R477 B.n865 B.n864 585
R478 B.n864 B.n863 585
R479 B.n465 B.n464 585
R480 B.n466 B.n465 585
R481 B.n856 B.n855 585
R482 B.n857 B.n856 585
R483 B.n854 B.n472 585
R484 B.n472 B.n471 585
R485 B.n853 B.n852 585
R486 B.n852 B.n851 585
R487 B.n474 B.n473 585
R488 B.n475 B.n474 585
R489 B.n844 B.n843 585
R490 B.n845 B.n844 585
R491 B.n842 B.n480 585
R492 B.n480 B.n479 585
R493 B.n841 B.n840 585
R494 B.n840 B.n839 585
R495 B.n482 B.n481 585
R496 B.n483 B.n482 585
R497 B.n832 B.n831 585
R498 B.n833 B.n832 585
R499 B.n830 B.n488 585
R500 B.n488 B.n487 585
R501 B.n829 B.n828 585
R502 B.n828 B.n827 585
R503 B.n490 B.n489 585
R504 B.n820 B.n490 585
R505 B.n819 B.n818 585
R506 B.n821 B.n819 585
R507 B.n817 B.n495 585
R508 B.n495 B.n494 585
R509 B.n816 B.n815 585
R510 B.n815 B.n814 585
R511 B.n497 B.n496 585
R512 B.n498 B.n497 585
R513 B.n807 B.n806 585
R514 B.n808 B.n807 585
R515 B.n805 B.n503 585
R516 B.n503 B.n502 585
R517 B.n804 B.n803 585
R518 B.n803 B.n802 585
R519 B.n505 B.n504 585
R520 B.n506 B.n505 585
R521 B.n798 B.n797 585
R522 B.n509 B.n508 585
R523 B.n794 B.n793 585
R524 B.n795 B.n794 585
R525 B.n792 B.n566 585
R526 B.n791 B.n790 585
R527 B.n789 B.n788 585
R528 B.n787 B.n786 585
R529 B.n785 B.n784 585
R530 B.n783 B.n782 585
R531 B.n781 B.n780 585
R532 B.n779 B.n778 585
R533 B.n777 B.n776 585
R534 B.n775 B.n774 585
R535 B.n773 B.n772 585
R536 B.n771 B.n770 585
R537 B.n769 B.n768 585
R538 B.n767 B.n766 585
R539 B.n765 B.n764 585
R540 B.n763 B.n762 585
R541 B.n761 B.n760 585
R542 B.n759 B.n758 585
R543 B.n757 B.n756 585
R544 B.n755 B.n754 585
R545 B.n753 B.n752 585
R546 B.n751 B.n750 585
R547 B.n749 B.n748 585
R548 B.n747 B.n746 585
R549 B.n745 B.n744 585
R550 B.n743 B.n742 585
R551 B.n741 B.n740 585
R552 B.n739 B.n738 585
R553 B.n737 B.n736 585
R554 B.n735 B.n734 585
R555 B.n733 B.n732 585
R556 B.n731 B.n730 585
R557 B.n729 B.n728 585
R558 B.n727 B.n726 585
R559 B.n725 B.n724 585
R560 B.n723 B.n722 585
R561 B.n721 B.n720 585
R562 B.n719 B.n718 585
R563 B.n717 B.n716 585
R564 B.n715 B.n714 585
R565 B.n713 B.n712 585
R566 B.n711 B.n710 585
R567 B.n709 B.n708 585
R568 B.n707 B.n706 585
R569 B.n705 B.n704 585
R570 B.n703 B.n702 585
R571 B.n701 B.n700 585
R572 B.n699 B.n698 585
R573 B.n697 B.n696 585
R574 B.n694 B.n693 585
R575 B.n692 B.n691 585
R576 B.n690 B.n689 585
R577 B.n688 B.n687 585
R578 B.n686 B.n685 585
R579 B.n684 B.n683 585
R580 B.n682 B.n681 585
R581 B.n680 B.n679 585
R582 B.n678 B.n677 585
R583 B.n676 B.n675 585
R584 B.n673 B.n672 585
R585 B.n671 B.n670 585
R586 B.n669 B.n668 585
R587 B.n667 B.n666 585
R588 B.n665 B.n664 585
R589 B.n663 B.n662 585
R590 B.n661 B.n660 585
R591 B.n659 B.n658 585
R592 B.n657 B.n656 585
R593 B.n655 B.n654 585
R594 B.n653 B.n652 585
R595 B.n651 B.n650 585
R596 B.n649 B.n648 585
R597 B.n647 B.n646 585
R598 B.n645 B.n644 585
R599 B.n643 B.n642 585
R600 B.n641 B.n640 585
R601 B.n639 B.n638 585
R602 B.n637 B.n636 585
R603 B.n635 B.n634 585
R604 B.n633 B.n632 585
R605 B.n631 B.n630 585
R606 B.n629 B.n628 585
R607 B.n627 B.n626 585
R608 B.n625 B.n624 585
R609 B.n623 B.n622 585
R610 B.n621 B.n620 585
R611 B.n619 B.n618 585
R612 B.n617 B.n616 585
R613 B.n615 B.n614 585
R614 B.n613 B.n612 585
R615 B.n611 B.n610 585
R616 B.n609 B.n608 585
R617 B.n607 B.n606 585
R618 B.n605 B.n604 585
R619 B.n603 B.n602 585
R620 B.n601 B.n600 585
R621 B.n599 B.n598 585
R622 B.n597 B.n596 585
R623 B.n595 B.n594 585
R624 B.n593 B.n592 585
R625 B.n591 B.n590 585
R626 B.n589 B.n588 585
R627 B.n587 B.n586 585
R628 B.n585 B.n584 585
R629 B.n583 B.n582 585
R630 B.n581 B.n580 585
R631 B.n579 B.n578 585
R632 B.n577 B.n576 585
R633 B.n575 B.n574 585
R634 B.n573 B.n572 585
R635 B.n571 B.n565 585
R636 B.n795 B.n565 585
R637 B.n799 B.n507 585
R638 B.n507 B.n506 585
R639 B.n801 B.n800 585
R640 B.n802 B.n801 585
R641 B.n501 B.n500 585
R642 B.n502 B.n501 585
R643 B.n810 B.n809 585
R644 B.n809 B.n808 585
R645 B.n811 B.n499 585
R646 B.n499 B.n498 585
R647 B.n813 B.n812 585
R648 B.n814 B.n813 585
R649 B.n493 B.n492 585
R650 B.n494 B.n493 585
R651 B.n823 B.n822 585
R652 B.n822 B.n821 585
R653 B.n824 B.n491 585
R654 B.n820 B.n491 585
R655 B.n826 B.n825 585
R656 B.n827 B.n826 585
R657 B.n486 B.n485 585
R658 B.n487 B.n486 585
R659 B.n835 B.n834 585
R660 B.n834 B.n833 585
R661 B.n836 B.n484 585
R662 B.n484 B.n483 585
R663 B.n838 B.n837 585
R664 B.n839 B.n838 585
R665 B.n478 B.n477 585
R666 B.n479 B.n478 585
R667 B.n847 B.n846 585
R668 B.n846 B.n845 585
R669 B.n848 B.n476 585
R670 B.n476 B.n475 585
R671 B.n850 B.n849 585
R672 B.n851 B.n850 585
R673 B.n470 B.n469 585
R674 B.n471 B.n470 585
R675 B.n859 B.n858 585
R676 B.n858 B.n857 585
R677 B.n860 B.n468 585
R678 B.n468 B.n466 585
R679 B.n862 B.n861 585
R680 B.n863 B.n862 585
R681 B.n462 B.n461 585
R682 B.n467 B.n462 585
R683 B.n871 B.n870 585
R684 B.n870 B.n869 585
R685 B.n872 B.n460 585
R686 B.n460 B.n459 585
R687 B.n874 B.n873 585
R688 B.n875 B.n874 585
R689 B.n454 B.n453 585
R690 B.n455 B.n454 585
R691 B.n883 B.n882 585
R692 B.n882 B.n881 585
R693 B.n884 B.n452 585
R694 B.n452 B.n451 585
R695 B.n886 B.n885 585
R696 B.n887 B.n886 585
R697 B.n446 B.n445 585
R698 B.n447 B.n446 585
R699 B.n896 B.n895 585
R700 B.n895 B.n894 585
R701 B.n897 B.n444 585
R702 B.n893 B.n444 585
R703 B.n899 B.n898 585
R704 B.n900 B.n899 585
R705 B.n439 B.n438 585
R706 B.n440 B.n439 585
R707 B.n908 B.n907 585
R708 B.n907 B.n906 585
R709 B.n909 B.n437 585
R710 B.n437 B.n436 585
R711 B.n911 B.n910 585
R712 B.n912 B.n911 585
R713 B.n431 B.n430 585
R714 B.n432 B.n431 585
R715 B.n920 B.n919 585
R716 B.n919 B.n918 585
R717 B.n921 B.n429 585
R718 B.n429 B.n427 585
R719 B.n923 B.n922 585
R720 B.n924 B.n923 585
R721 B.n423 B.n422 585
R722 B.n428 B.n423 585
R723 B.n932 B.n931 585
R724 B.n931 B.n930 585
R725 B.n933 B.n421 585
R726 B.n421 B.n420 585
R727 B.n935 B.n934 585
R728 B.n936 B.n935 585
R729 B.n415 B.n414 585
R730 B.n416 B.n415 585
R731 B.n944 B.n943 585
R732 B.n943 B.n942 585
R733 B.n945 B.n413 585
R734 B.n413 B.n412 585
R735 B.n947 B.n946 585
R736 B.n948 B.n947 585
R737 B.n407 B.n406 585
R738 B.n408 B.n407 585
R739 B.n957 B.n956 585
R740 B.n956 B.n955 585
R741 B.n958 B.n405 585
R742 B.n954 B.n405 585
R743 B.n960 B.n959 585
R744 B.n961 B.n960 585
R745 B.n400 B.n399 585
R746 B.n401 B.n400 585
R747 B.n970 B.n969 585
R748 B.n969 B.n968 585
R749 B.n971 B.n398 585
R750 B.n398 B.n397 585
R751 B.n973 B.n972 585
R752 B.n974 B.n973 585
R753 B.n3 B.n0 585
R754 B.n4 B.n3 585
R755 B.n1176 B.n1 585
R756 B.n1177 B.n1176 585
R757 B.n1175 B.n1174 585
R758 B.n1175 B.n8 585
R759 B.n1173 B.n9 585
R760 B.n12 B.n9 585
R761 B.n1172 B.n1171 585
R762 B.n1171 B.n1170 585
R763 B.n11 B.n10 585
R764 B.n1169 B.n11 585
R765 B.n1167 B.n1166 585
R766 B.n1168 B.n1167 585
R767 B.n1165 B.n16 585
R768 B.n19 B.n16 585
R769 B.n1164 B.n1163 585
R770 B.n1163 B.n1162 585
R771 B.n18 B.n17 585
R772 B.n1161 B.n18 585
R773 B.n1159 B.n1158 585
R774 B.n1160 B.n1159 585
R775 B.n1157 B.n24 585
R776 B.n24 B.n23 585
R777 B.n1156 B.n1155 585
R778 B.n1155 B.n1154 585
R779 B.n26 B.n25 585
R780 B.n1153 B.n26 585
R781 B.n1151 B.n1150 585
R782 B.n1152 B.n1151 585
R783 B.n1149 B.n31 585
R784 B.n31 B.n30 585
R785 B.n1148 B.n1147 585
R786 B.n1147 B.n1146 585
R787 B.n33 B.n32 585
R788 B.n1145 B.n33 585
R789 B.n1143 B.n1142 585
R790 B.n1144 B.n1143 585
R791 B.n1141 B.n38 585
R792 B.n38 B.n37 585
R793 B.n1140 B.n1139 585
R794 B.n1139 B.n1138 585
R795 B.n40 B.n39 585
R796 B.n1137 B.n40 585
R797 B.n1135 B.n1134 585
R798 B.n1136 B.n1135 585
R799 B.n1133 B.n45 585
R800 B.n45 B.n44 585
R801 B.n1132 B.n1131 585
R802 B.n1131 B.n1130 585
R803 B.n47 B.n46 585
R804 B.n1129 B.n47 585
R805 B.n1127 B.n1126 585
R806 B.n1128 B.n1127 585
R807 B.n1125 B.n51 585
R808 B.n54 B.n51 585
R809 B.n1124 B.n1123 585
R810 B.n1123 B.n1122 585
R811 B.n53 B.n52 585
R812 B.n1121 B.n53 585
R813 B.n1119 B.n1118 585
R814 B.n1120 B.n1119 585
R815 B.n1117 B.n59 585
R816 B.n59 B.n58 585
R817 B.n1116 B.n1115 585
R818 B.n1115 B.n1114 585
R819 B.n61 B.n60 585
R820 B.n1113 B.n61 585
R821 B.n1111 B.n1110 585
R822 B.n1112 B.n1111 585
R823 B.n1109 B.n66 585
R824 B.n66 B.n65 585
R825 B.n1108 B.n1107 585
R826 B.n1107 B.n1106 585
R827 B.n68 B.n67 585
R828 B.n1105 B.n68 585
R829 B.n1103 B.n1102 585
R830 B.n1104 B.n1103 585
R831 B.n1101 B.n73 585
R832 B.n73 B.n72 585
R833 B.n1100 B.n1099 585
R834 B.n1099 B.n1098 585
R835 B.n75 B.n74 585
R836 B.n1097 B.n75 585
R837 B.n1095 B.n1094 585
R838 B.n1096 B.n1095 585
R839 B.n1093 B.n80 585
R840 B.n80 B.n79 585
R841 B.n1092 B.n1091 585
R842 B.n1091 B.n1090 585
R843 B.n82 B.n81 585
R844 B.n1089 B.n82 585
R845 B.n1087 B.n1086 585
R846 B.n1088 B.n1087 585
R847 B.n1085 B.n87 585
R848 B.n87 B.n86 585
R849 B.n1084 B.n1083 585
R850 B.n1083 B.n1082 585
R851 B.n89 B.n88 585
R852 B.n1081 B.n89 585
R853 B.n1079 B.n1078 585
R854 B.n1080 B.n1079 585
R855 B.n1077 B.n93 585
R856 B.n96 B.n93 585
R857 B.n1076 B.n1075 585
R858 B.n1075 B.n1074 585
R859 B.n95 B.n94 585
R860 B.n1073 B.n95 585
R861 B.n1071 B.n1070 585
R862 B.n1072 B.n1071 585
R863 B.n1069 B.n101 585
R864 B.n101 B.n100 585
R865 B.n1068 B.n1067 585
R866 B.n1067 B.n1066 585
R867 B.n103 B.n102 585
R868 B.n1065 B.n103 585
R869 B.n1063 B.n1062 585
R870 B.n1064 B.n1063 585
R871 B.n1061 B.n108 585
R872 B.n108 B.n107 585
R873 B.n1180 B.n1179 585
R874 B.n1178 B.n2 585
R875 B.n1059 B.n108 506.916
R876 B.n1055 B.n167 506.916
R877 B.n565 B.n505 506.916
R878 B.n797 B.n507 506.916
R879 B.n171 B.t12 328.791
R880 B.n168 B.t19 328.791
R881 B.n569 B.t8 328.791
R882 B.n567 B.t16 328.791
R883 B.n1057 B.n1056 256.663
R884 B.n1057 B.n165 256.663
R885 B.n1057 B.n164 256.663
R886 B.n1057 B.n163 256.663
R887 B.n1057 B.n162 256.663
R888 B.n1057 B.n161 256.663
R889 B.n1057 B.n160 256.663
R890 B.n1057 B.n159 256.663
R891 B.n1057 B.n158 256.663
R892 B.n1057 B.n157 256.663
R893 B.n1057 B.n156 256.663
R894 B.n1057 B.n155 256.663
R895 B.n1057 B.n154 256.663
R896 B.n1057 B.n153 256.663
R897 B.n1057 B.n152 256.663
R898 B.n1057 B.n151 256.663
R899 B.n1057 B.n150 256.663
R900 B.n1057 B.n149 256.663
R901 B.n1057 B.n148 256.663
R902 B.n1057 B.n147 256.663
R903 B.n1057 B.n146 256.663
R904 B.n1057 B.n145 256.663
R905 B.n1057 B.n144 256.663
R906 B.n1057 B.n143 256.663
R907 B.n1057 B.n142 256.663
R908 B.n1057 B.n141 256.663
R909 B.n1057 B.n140 256.663
R910 B.n1057 B.n139 256.663
R911 B.n1057 B.n138 256.663
R912 B.n1057 B.n137 256.663
R913 B.n1057 B.n136 256.663
R914 B.n1057 B.n135 256.663
R915 B.n1057 B.n134 256.663
R916 B.n1057 B.n133 256.663
R917 B.n1057 B.n132 256.663
R918 B.n1057 B.n131 256.663
R919 B.n1057 B.n130 256.663
R920 B.n1057 B.n129 256.663
R921 B.n1057 B.n128 256.663
R922 B.n1057 B.n127 256.663
R923 B.n1057 B.n126 256.663
R924 B.n1057 B.n125 256.663
R925 B.n1057 B.n124 256.663
R926 B.n1057 B.n123 256.663
R927 B.n1057 B.n122 256.663
R928 B.n1057 B.n121 256.663
R929 B.n1057 B.n120 256.663
R930 B.n1057 B.n119 256.663
R931 B.n1057 B.n118 256.663
R932 B.n1057 B.n117 256.663
R933 B.n1057 B.n116 256.663
R934 B.n1057 B.n115 256.663
R935 B.n1057 B.n114 256.663
R936 B.n1057 B.n113 256.663
R937 B.n1057 B.n112 256.663
R938 B.n1057 B.n111 256.663
R939 B.n1058 B.n1057 256.663
R940 B.n796 B.n795 256.663
R941 B.n795 B.n510 256.663
R942 B.n795 B.n511 256.663
R943 B.n795 B.n512 256.663
R944 B.n795 B.n513 256.663
R945 B.n795 B.n514 256.663
R946 B.n795 B.n515 256.663
R947 B.n795 B.n516 256.663
R948 B.n795 B.n517 256.663
R949 B.n795 B.n518 256.663
R950 B.n795 B.n519 256.663
R951 B.n795 B.n520 256.663
R952 B.n795 B.n521 256.663
R953 B.n795 B.n522 256.663
R954 B.n795 B.n523 256.663
R955 B.n795 B.n524 256.663
R956 B.n795 B.n525 256.663
R957 B.n795 B.n526 256.663
R958 B.n795 B.n527 256.663
R959 B.n795 B.n528 256.663
R960 B.n795 B.n529 256.663
R961 B.n795 B.n530 256.663
R962 B.n795 B.n531 256.663
R963 B.n795 B.n532 256.663
R964 B.n795 B.n533 256.663
R965 B.n795 B.n534 256.663
R966 B.n795 B.n535 256.663
R967 B.n795 B.n536 256.663
R968 B.n795 B.n537 256.663
R969 B.n795 B.n538 256.663
R970 B.n795 B.n539 256.663
R971 B.n795 B.n540 256.663
R972 B.n795 B.n541 256.663
R973 B.n795 B.n542 256.663
R974 B.n795 B.n543 256.663
R975 B.n795 B.n544 256.663
R976 B.n795 B.n545 256.663
R977 B.n795 B.n546 256.663
R978 B.n795 B.n547 256.663
R979 B.n795 B.n548 256.663
R980 B.n795 B.n549 256.663
R981 B.n795 B.n550 256.663
R982 B.n795 B.n551 256.663
R983 B.n795 B.n552 256.663
R984 B.n795 B.n553 256.663
R985 B.n795 B.n554 256.663
R986 B.n795 B.n555 256.663
R987 B.n795 B.n556 256.663
R988 B.n795 B.n557 256.663
R989 B.n795 B.n558 256.663
R990 B.n795 B.n559 256.663
R991 B.n795 B.n560 256.663
R992 B.n795 B.n561 256.663
R993 B.n795 B.n562 256.663
R994 B.n795 B.n563 256.663
R995 B.n795 B.n564 256.663
R996 B.n1182 B.n1181 256.663
R997 B.n174 B.n110 163.367
R998 B.n178 B.n177 163.367
R999 B.n182 B.n181 163.367
R1000 B.n186 B.n185 163.367
R1001 B.n190 B.n189 163.367
R1002 B.n194 B.n193 163.367
R1003 B.n198 B.n197 163.367
R1004 B.n202 B.n201 163.367
R1005 B.n206 B.n205 163.367
R1006 B.n210 B.n209 163.367
R1007 B.n214 B.n213 163.367
R1008 B.n218 B.n217 163.367
R1009 B.n222 B.n221 163.367
R1010 B.n226 B.n225 163.367
R1011 B.n230 B.n229 163.367
R1012 B.n234 B.n233 163.367
R1013 B.n238 B.n237 163.367
R1014 B.n242 B.n241 163.367
R1015 B.n246 B.n245 163.367
R1016 B.n250 B.n249 163.367
R1017 B.n254 B.n253 163.367
R1018 B.n258 B.n257 163.367
R1019 B.n262 B.n261 163.367
R1020 B.n266 B.n265 163.367
R1021 B.n270 B.n269 163.367
R1022 B.n274 B.n273 163.367
R1023 B.n278 B.n277 163.367
R1024 B.n282 B.n281 163.367
R1025 B.n286 B.n285 163.367
R1026 B.n290 B.n289 163.367
R1027 B.n294 B.n293 163.367
R1028 B.n298 B.n297 163.367
R1029 B.n302 B.n301 163.367
R1030 B.n306 B.n305 163.367
R1031 B.n310 B.n309 163.367
R1032 B.n314 B.n313 163.367
R1033 B.n318 B.n317 163.367
R1034 B.n322 B.n321 163.367
R1035 B.n326 B.n325 163.367
R1036 B.n330 B.n329 163.367
R1037 B.n334 B.n333 163.367
R1038 B.n338 B.n337 163.367
R1039 B.n342 B.n341 163.367
R1040 B.n346 B.n345 163.367
R1041 B.n350 B.n349 163.367
R1042 B.n354 B.n353 163.367
R1043 B.n358 B.n357 163.367
R1044 B.n362 B.n361 163.367
R1045 B.n366 B.n365 163.367
R1046 B.n370 B.n369 163.367
R1047 B.n374 B.n373 163.367
R1048 B.n378 B.n377 163.367
R1049 B.n382 B.n381 163.367
R1050 B.n386 B.n385 163.367
R1051 B.n390 B.n389 163.367
R1052 B.n392 B.n166 163.367
R1053 B.n803 B.n505 163.367
R1054 B.n803 B.n503 163.367
R1055 B.n807 B.n503 163.367
R1056 B.n807 B.n497 163.367
R1057 B.n815 B.n497 163.367
R1058 B.n815 B.n495 163.367
R1059 B.n819 B.n495 163.367
R1060 B.n819 B.n490 163.367
R1061 B.n828 B.n490 163.367
R1062 B.n828 B.n488 163.367
R1063 B.n832 B.n488 163.367
R1064 B.n832 B.n482 163.367
R1065 B.n840 B.n482 163.367
R1066 B.n840 B.n480 163.367
R1067 B.n844 B.n480 163.367
R1068 B.n844 B.n474 163.367
R1069 B.n852 B.n474 163.367
R1070 B.n852 B.n472 163.367
R1071 B.n856 B.n472 163.367
R1072 B.n856 B.n465 163.367
R1073 B.n864 B.n465 163.367
R1074 B.n864 B.n463 163.367
R1075 B.n868 B.n463 163.367
R1076 B.n868 B.n458 163.367
R1077 B.n876 B.n458 163.367
R1078 B.n876 B.n456 163.367
R1079 B.n880 B.n456 163.367
R1080 B.n880 B.n450 163.367
R1081 B.n888 B.n450 163.367
R1082 B.n888 B.n448 163.367
R1083 B.n892 B.n448 163.367
R1084 B.n892 B.n443 163.367
R1085 B.n901 B.n443 163.367
R1086 B.n901 B.n441 163.367
R1087 B.n905 B.n441 163.367
R1088 B.n905 B.n435 163.367
R1089 B.n913 B.n435 163.367
R1090 B.n913 B.n433 163.367
R1091 B.n917 B.n433 163.367
R1092 B.n917 B.n426 163.367
R1093 B.n925 B.n426 163.367
R1094 B.n925 B.n424 163.367
R1095 B.n929 B.n424 163.367
R1096 B.n929 B.n419 163.367
R1097 B.n937 B.n419 163.367
R1098 B.n937 B.n417 163.367
R1099 B.n941 B.n417 163.367
R1100 B.n941 B.n411 163.367
R1101 B.n949 B.n411 163.367
R1102 B.n949 B.n409 163.367
R1103 B.n953 B.n409 163.367
R1104 B.n953 B.n404 163.367
R1105 B.n962 B.n404 163.367
R1106 B.n962 B.n402 163.367
R1107 B.n967 B.n402 163.367
R1108 B.n967 B.n396 163.367
R1109 B.n975 B.n396 163.367
R1110 B.n976 B.n975 163.367
R1111 B.n976 B.n5 163.367
R1112 B.n6 B.n5 163.367
R1113 B.n7 B.n6 163.367
R1114 B.n982 B.n7 163.367
R1115 B.n983 B.n982 163.367
R1116 B.n983 B.n13 163.367
R1117 B.n14 B.n13 163.367
R1118 B.n15 B.n14 163.367
R1119 B.n988 B.n15 163.367
R1120 B.n988 B.n20 163.367
R1121 B.n21 B.n20 163.367
R1122 B.n22 B.n21 163.367
R1123 B.n993 B.n22 163.367
R1124 B.n993 B.n27 163.367
R1125 B.n28 B.n27 163.367
R1126 B.n29 B.n28 163.367
R1127 B.n998 B.n29 163.367
R1128 B.n998 B.n34 163.367
R1129 B.n35 B.n34 163.367
R1130 B.n36 B.n35 163.367
R1131 B.n1003 B.n36 163.367
R1132 B.n1003 B.n41 163.367
R1133 B.n42 B.n41 163.367
R1134 B.n43 B.n42 163.367
R1135 B.n1008 B.n43 163.367
R1136 B.n1008 B.n48 163.367
R1137 B.n49 B.n48 163.367
R1138 B.n50 B.n49 163.367
R1139 B.n1013 B.n50 163.367
R1140 B.n1013 B.n55 163.367
R1141 B.n56 B.n55 163.367
R1142 B.n57 B.n56 163.367
R1143 B.n1018 B.n57 163.367
R1144 B.n1018 B.n62 163.367
R1145 B.n63 B.n62 163.367
R1146 B.n64 B.n63 163.367
R1147 B.n1023 B.n64 163.367
R1148 B.n1023 B.n69 163.367
R1149 B.n70 B.n69 163.367
R1150 B.n71 B.n70 163.367
R1151 B.n1028 B.n71 163.367
R1152 B.n1028 B.n76 163.367
R1153 B.n77 B.n76 163.367
R1154 B.n78 B.n77 163.367
R1155 B.n1033 B.n78 163.367
R1156 B.n1033 B.n83 163.367
R1157 B.n84 B.n83 163.367
R1158 B.n85 B.n84 163.367
R1159 B.n1038 B.n85 163.367
R1160 B.n1038 B.n90 163.367
R1161 B.n91 B.n90 163.367
R1162 B.n92 B.n91 163.367
R1163 B.n1043 B.n92 163.367
R1164 B.n1043 B.n97 163.367
R1165 B.n98 B.n97 163.367
R1166 B.n99 B.n98 163.367
R1167 B.n1048 B.n99 163.367
R1168 B.n1048 B.n104 163.367
R1169 B.n105 B.n104 163.367
R1170 B.n106 B.n105 163.367
R1171 B.n167 B.n106 163.367
R1172 B.n794 B.n509 163.367
R1173 B.n794 B.n566 163.367
R1174 B.n790 B.n789 163.367
R1175 B.n786 B.n785 163.367
R1176 B.n782 B.n781 163.367
R1177 B.n778 B.n777 163.367
R1178 B.n774 B.n773 163.367
R1179 B.n770 B.n769 163.367
R1180 B.n766 B.n765 163.367
R1181 B.n762 B.n761 163.367
R1182 B.n758 B.n757 163.367
R1183 B.n754 B.n753 163.367
R1184 B.n750 B.n749 163.367
R1185 B.n746 B.n745 163.367
R1186 B.n742 B.n741 163.367
R1187 B.n738 B.n737 163.367
R1188 B.n734 B.n733 163.367
R1189 B.n730 B.n729 163.367
R1190 B.n726 B.n725 163.367
R1191 B.n722 B.n721 163.367
R1192 B.n718 B.n717 163.367
R1193 B.n714 B.n713 163.367
R1194 B.n710 B.n709 163.367
R1195 B.n706 B.n705 163.367
R1196 B.n702 B.n701 163.367
R1197 B.n698 B.n697 163.367
R1198 B.n693 B.n692 163.367
R1199 B.n689 B.n688 163.367
R1200 B.n685 B.n684 163.367
R1201 B.n681 B.n680 163.367
R1202 B.n677 B.n676 163.367
R1203 B.n672 B.n671 163.367
R1204 B.n668 B.n667 163.367
R1205 B.n664 B.n663 163.367
R1206 B.n660 B.n659 163.367
R1207 B.n656 B.n655 163.367
R1208 B.n652 B.n651 163.367
R1209 B.n648 B.n647 163.367
R1210 B.n644 B.n643 163.367
R1211 B.n640 B.n639 163.367
R1212 B.n636 B.n635 163.367
R1213 B.n632 B.n631 163.367
R1214 B.n628 B.n627 163.367
R1215 B.n624 B.n623 163.367
R1216 B.n620 B.n619 163.367
R1217 B.n616 B.n615 163.367
R1218 B.n612 B.n611 163.367
R1219 B.n608 B.n607 163.367
R1220 B.n604 B.n603 163.367
R1221 B.n600 B.n599 163.367
R1222 B.n596 B.n595 163.367
R1223 B.n592 B.n591 163.367
R1224 B.n588 B.n587 163.367
R1225 B.n584 B.n583 163.367
R1226 B.n580 B.n579 163.367
R1227 B.n576 B.n575 163.367
R1228 B.n572 B.n565 163.367
R1229 B.n801 B.n507 163.367
R1230 B.n801 B.n501 163.367
R1231 B.n809 B.n501 163.367
R1232 B.n809 B.n499 163.367
R1233 B.n813 B.n499 163.367
R1234 B.n813 B.n493 163.367
R1235 B.n822 B.n493 163.367
R1236 B.n822 B.n491 163.367
R1237 B.n826 B.n491 163.367
R1238 B.n826 B.n486 163.367
R1239 B.n834 B.n486 163.367
R1240 B.n834 B.n484 163.367
R1241 B.n838 B.n484 163.367
R1242 B.n838 B.n478 163.367
R1243 B.n846 B.n478 163.367
R1244 B.n846 B.n476 163.367
R1245 B.n850 B.n476 163.367
R1246 B.n850 B.n470 163.367
R1247 B.n858 B.n470 163.367
R1248 B.n858 B.n468 163.367
R1249 B.n862 B.n468 163.367
R1250 B.n862 B.n462 163.367
R1251 B.n870 B.n462 163.367
R1252 B.n870 B.n460 163.367
R1253 B.n874 B.n460 163.367
R1254 B.n874 B.n454 163.367
R1255 B.n882 B.n454 163.367
R1256 B.n882 B.n452 163.367
R1257 B.n886 B.n452 163.367
R1258 B.n886 B.n446 163.367
R1259 B.n895 B.n446 163.367
R1260 B.n895 B.n444 163.367
R1261 B.n899 B.n444 163.367
R1262 B.n899 B.n439 163.367
R1263 B.n907 B.n439 163.367
R1264 B.n907 B.n437 163.367
R1265 B.n911 B.n437 163.367
R1266 B.n911 B.n431 163.367
R1267 B.n919 B.n431 163.367
R1268 B.n919 B.n429 163.367
R1269 B.n923 B.n429 163.367
R1270 B.n923 B.n423 163.367
R1271 B.n931 B.n423 163.367
R1272 B.n931 B.n421 163.367
R1273 B.n935 B.n421 163.367
R1274 B.n935 B.n415 163.367
R1275 B.n943 B.n415 163.367
R1276 B.n943 B.n413 163.367
R1277 B.n947 B.n413 163.367
R1278 B.n947 B.n407 163.367
R1279 B.n956 B.n407 163.367
R1280 B.n956 B.n405 163.367
R1281 B.n960 B.n405 163.367
R1282 B.n960 B.n400 163.367
R1283 B.n969 B.n400 163.367
R1284 B.n969 B.n398 163.367
R1285 B.n973 B.n398 163.367
R1286 B.n973 B.n3 163.367
R1287 B.n1180 B.n3 163.367
R1288 B.n1176 B.n2 163.367
R1289 B.n1176 B.n1175 163.367
R1290 B.n1175 B.n9 163.367
R1291 B.n1171 B.n9 163.367
R1292 B.n1171 B.n11 163.367
R1293 B.n1167 B.n11 163.367
R1294 B.n1167 B.n16 163.367
R1295 B.n1163 B.n16 163.367
R1296 B.n1163 B.n18 163.367
R1297 B.n1159 B.n18 163.367
R1298 B.n1159 B.n24 163.367
R1299 B.n1155 B.n24 163.367
R1300 B.n1155 B.n26 163.367
R1301 B.n1151 B.n26 163.367
R1302 B.n1151 B.n31 163.367
R1303 B.n1147 B.n31 163.367
R1304 B.n1147 B.n33 163.367
R1305 B.n1143 B.n33 163.367
R1306 B.n1143 B.n38 163.367
R1307 B.n1139 B.n38 163.367
R1308 B.n1139 B.n40 163.367
R1309 B.n1135 B.n40 163.367
R1310 B.n1135 B.n45 163.367
R1311 B.n1131 B.n45 163.367
R1312 B.n1131 B.n47 163.367
R1313 B.n1127 B.n47 163.367
R1314 B.n1127 B.n51 163.367
R1315 B.n1123 B.n51 163.367
R1316 B.n1123 B.n53 163.367
R1317 B.n1119 B.n53 163.367
R1318 B.n1119 B.n59 163.367
R1319 B.n1115 B.n59 163.367
R1320 B.n1115 B.n61 163.367
R1321 B.n1111 B.n61 163.367
R1322 B.n1111 B.n66 163.367
R1323 B.n1107 B.n66 163.367
R1324 B.n1107 B.n68 163.367
R1325 B.n1103 B.n68 163.367
R1326 B.n1103 B.n73 163.367
R1327 B.n1099 B.n73 163.367
R1328 B.n1099 B.n75 163.367
R1329 B.n1095 B.n75 163.367
R1330 B.n1095 B.n80 163.367
R1331 B.n1091 B.n80 163.367
R1332 B.n1091 B.n82 163.367
R1333 B.n1087 B.n82 163.367
R1334 B.n1087 B.n87 163.367
R1335 B.n1083 B.n87 163.367
R1336 B.n1083 B.n89 163.367
R1337 B.n1079 B.n89 163.367
R1338 B.n1079 B.n93 163.367
R1339 B.n1075 B.n93 163.367
R1340 B.n1075 B.n95 163.367
R1341 B.n1071 B.n95 163.367
R1342 B.n1071 B.n101 163.367
R1343 B.n1067 B.n101 163.367
R1344 B.n1067 B.n103 163.367
R1345 B.n1063 B.n103 163.367
R1346 B.n1063 B.n108 163.367
R1347 B.n168 B.t20 135.869
R1348 B.n569 B.t11 135.869
R1349 B.n171 B.t14 135.847
R1350 B.n567 B.t18 135.847
R1351 B.n1059 B.n1058 71.676
R1352 B.n174 B.n111 71.676
R1353 B.n178 B.n112 71.676
R1354 B.n182 B.n113 71.676
R1355 B.n186 B.n114 71.676
R1356 B.n190 B.n115 71.676
R1357 B.n194 B.n116 71.676
R1358 B.n198 B.n117 71.676
R1359 B.n202 B.n118 71.676
R1360 B.n206 B.n119 71.676
R1361 B.n210 B.n120 71.676
R1362 B.n214 B.n121 71.676
R1363 B.n218 B.n122 71.676
R1364 B.n222 B.n123 71.676
R1365 B.n226 B.n124 71.676
R1366 B.n230 B.n125 71.676
R1367 B.n234 B.n126 71.676
R1368 B.n238 B.n127 71.676
R1369 B.n242 B.n128 71.676
R1370 B.n246 B.n129 71.676
R1371 B.n250 B.n130 71.676
R1372 B.n254 B.n131 71.676
R1373 B.n258 B.n132 71.676
R1374 B.n262 B.n133 71.676
R1375 B.n266 B.n134 71.676
R1376 B.n270 B.n135 71.676
R1377 B.n274 B.n136 71.676
R1378 B.n278 B.n137 71.676
R1379 B.n282 B.n138 71.676
R1380 B.n286 B.n139 71.676
R1381 B.n290 B.n140 71.676
R1382 B.n294 B.n141 71.676
R1383 B.n298 B.n142 71.676
R1384 B.n302 B.n143 71.676
R1385 B.n306 B.n144 71.676
R1386 B.n310 B.n145 71.676
R1387 B.n314 B.n146 71.676
R1388 B.n318 B.n147 71.676
R1389 B.n322 B.n148 71.676
R1390 B.n326 B.n149 71.676
R1391 B.n330 B.n150 71.676
R1392 B.n334 B.n151 71.676
R1393 B.n338 B.n152 71.676
R1394 B.n342 B.n153 71.676
R1395 B.n346 B.n154 71.676
R1396 B.n350 B.n155 71.676
R1397 B.n354 B.n156 71.676
R1398 B.n358 B.n157 71.676
R1399 B.n362 B.n158 71.676
R1400 B.n366 B.n159 71.676
R1401 B.n370 B.n160 71.676
R1402 B.n374 B.n161 71.676
R1403 B.n378 B.n162 71.676
R1404 B.n382 B.n163 71.676
R1405 B.n386 B.n164 71.676
R1406 B.n390 B.n165 71.676
R1407 B.n1056 B.n166 71.676
R1408 B.n1056 B.n1055 71.676
R1409 B.n392 B.n165 71.676
R1410 B.n389 B.n164 71.676
R1411 B.n385 B.n163 71.676
R1412 B.n381 B.n162 71.676
R1413 B.n377 B.n161 71.676
R1414 B.n373 B.n160 71.676
R1415 B.n369 B.n159 71.676
R1416 B.n365 B.n158 71.676
R1417 B.n361 B.n157 71.676
R1418 B.n357 B.n156 71.676
R1419 B.n353 B.n155 71.676
R1420 B.n349 B.n154 71.676
R1421 B.n345 B.n153 71.676
R1422 B.n341 B.n152 71.676
R1423 B.n337 B.n151 71.676
R1424 B.n333 B.n150 71.676
R1425 B.n329 B.n149 71.676
R1426 B.n325 B.n148 71.676
R1427 B.n321 B.n147 71.676
R1428 B.n317 B.n146 71.676
R1429 B.n313 B.n145 71.676
R1430 B.n309 B.n144 71.676
R1431 B.n305 B.n143 71.676
R1432 B.n301 B.n142 71.676
R1433 B.n297 B.n141 71.676
R1434 B.n293 B.n140 71.676
R1435 B.n289 B.n139 71.676
R1436 B.n285 B.n138 71.676
R1437 B.n281 B.n137 71.676
R1438 B.n277 B.n136 71.676
R1439 B.n273 B.n135 71.676
R1440 B.n269 B.n134 71.676
R1441 B.n265 B.n133 71.676
R1442 B.n261 B.n132 71.676
R1443 B.n257 B.n131 71.676
R1444 B.n253 B.n130 71.676
R1445 B.n249 B.n129 71.676
R1446 B.n245 B.n128 71.676
R1447 B.n241 B.n127 71.676
R1448 B.n237 B.n126 71.676
R1449 B.n233 B.n125 71.676
R1450 B.n229 B.n124 71.676
R1451 B.n225 B.n123 71.676
R1452 B.n221 B.n122 71.676
R1453 B.n217 B.n121 71.676
R1454 B.n213 B.n120 71.676
R1455 B.n209 B.n119 71.676
R1456 B.n205 B.n118 71.676
R1457 B.n201 B.n117 71.676
R1458 B.n197 B.n116 71.676
R1459 B.n193 B.n115 71.676
R1460 B.n189 B.n114 71.676
R1461 B.n185 B.n113 71.676
R1462 B.n181 B.n112 71.676
R1463 B.n177 B.n111 71.676
R1464 B.n1058 B.n110 71.676
R1465 B.n797 B.n796 71.676
R1466 B.n566 B.n510 71.676
R1467 B.n789 B.n511 71.676
R1468 B.n785 B.n512 71.676
R1469 B.n781 B.n513 71.676
R1470 B.n777 B.n514 71.676
R1471 B.n773 B.n515 71.676
R1472 B.n769 B.n516 71.676
R1473 B.n765 B.n517 71.676
R1474 B.n761 B.n518 71.676
R1475 B.n757 B.n519 71.676
R1476 B.n753 B.n520 71.676
R1477 B.n749 B.n521 71.676
R1478 B.n745 B.n522 71.676
R1479 B.n741 B.n523 71.676
R1480 B.n737 B.n524 71.676
R1481 B.n733 B.n525 71.676
R1482 B.n729 B.n526 71.676
R1483 B.n725 B.n527 71.676
R1484 B.n721 B.n528 71.676
R1485 B.n717 B.n529 71.676
R1486 B.n713 B.n530 71.676
R1487 B.n709 B.n531 71.676
R1488 B.n705 B.n532 71.676
R1489 B.n701 B.n533 71.676
R1490 B.n697 B.n534 71.676
R1491 B.n692 B.n535 71.676
R1492 B.n688 B.n536 71.676
R1493 B.n684 B.n537 71.676
R1494 B.n680 B.n538 71.676
R1495 B.n676 B.n539 71.676
R1496 B.n671 B.n540 71.676
R1497 B.n667 B.n541 71.676
R1498 B.n663 B.n542 71.676
R1499 B.n659 B.n543 71.676
R1500 B.n655 B.n544 71.676
R1501 B.n651 B.n545 71.676
R1502 B.n647 B.n546 71.676
R1503 B.n643 B.n547 71.676
R1504 B.n639 B.n548 71.676
R1505 B.n635 B.n549 71.676
R1506 B.n631 B.n550 71.676
R1507 B.n627 B.n551 71.676
R1508 B.n623 B.n552 71.676
R1509 B.n619 B.n553 71.676
R1510 B.n615 B.n554 71.676
R1511 B.n611 B.n555 71.676
R1512 B.n607 B.n556 71.676
R1513 B.n603 B.n557 71.676
R1514 B.n599 B.n558 71.676
R1515 B.n595 B.n559 71.676
R1516 B.n591 B.n560 71.676
R1517 B.n587 B.n561 71.676
R1518 B.n583 B.n562 71.676
R1519 B.n579 B.n563 71.676
R1520 B.n575 B.n564 71.676
R1521 B.n796 B.n509 71.676
R1522 B.n790 B.n510 71.676
R1523 B.n786 B.n511 71.676
R1524 B.n782 B.n512 71.676
R1525 B.n778 B.n513 71.676
R1526 B.n774 B.n514 71.676
R1527 B.n770 B.n515 71.676
R1528 B.n766 B.n516 71.676
R1529 B.n762 B.n517 71.676
R1530 B.n758 B.n518 71.676
R1531 B.n754 B.n519 71.676
R1532 B.n750 B.n520 71.676
R1533 B.n746 B.n521 71.676
R1534 B.n742 B.n522 71.676
R1535 B.n738 B.n523 71.676
R1536 B.n734 B.n524 71.676
R1537 B.n730 B.n525 71.676
R1538 B.n726 B.n526 71.676
R1539 B.n722 B.n527 71.676
R1540 B.n718 B.n528 71.676
R1541 B.n714 B.n529 71.676
R1542 B.n710 B.n530 71.676
R1543 B.n706 B.n531 71.676
R1544 B.n702 B.n532 71.676
R1545 B.n698 B.n533 71.676
R1546 B.n693 B.n534 71.676
R1547 B.n689 B.n535 71.676
R1548 B.n685 B.n536 71.676
R1549 B.n681 B.n537 71.676
R1550 B.n677 B.n538 71.676
R1551 B.n672 B.n539 71.676
R1552 B.n668 B.n540 71.676
R1553 B.n664 B.n541 71.676
R1554 B.n660 B.n542 71.676
R1555 B.n656 B.n543 71.676
R1556 B.n652 B.n544 71.676
R1557 B.n648 B.n545 71.676
R1558 B.n644 B.n546 71.676
R1559 B.n640 B.n547 71.676
R1560 B.n636 B.n548 71.676
R1561 B.n632 B.n549 71.676
R1562 B.n628 B.n550 71.676
R1563 B.n624 B.n551 71.676
R1564 B.n620 B.n552 71.676
R1565 B.n616 B.n553 71.676
R1566 B.n612 B.n554 71.676
R1567 B.n608 B.n555 71.676
R1568 B.n604 B.n556 71.676
R1569 B.n600 B.n557 71.676
R1570 B.n596 B.n558 71.676
R1571 B.n592 B.n559 71.676
R1572 B.n588 B.n560 71.676
R1573 B.n584 B.n561 71.676
R1574 B.n580 B.n562 71.676
R1575 B.n576 B.n563 71.676
R1576 B.n572 B.n564 71.676
R1577 B.n1181 B.n1180 71.676
R1578 B.n1181 B.n2 71.676
R1579 B.n169 B.t21 68.377
R1580 B.n570 B.t10 68.377
R1581 B.n172 B.t15 68.3563
R1582 B.n568 B.t17 68.3563
R1583 B.n172 B.n171 67.4914
R1584 B.n169 B.n168 67.4914
R1585 B.n570 B.n569 67.4914
R1586 B.n568 B.n567 67.4914
R1587 B.n173 B.n172 59.5399
R1588 B.n170 B.n169 59.5399
R1589 B.n674 B.n570 59.5399
R1590 B.n695 B.n568 59.5399
R1591 B.n795 B.n506 57.1911
R1592 B.n1057 B.n107 57.1911
R1593 B.n802 B.n506 35.679
R1594 B.n802 B.n502 35.679
R1595 B.n808 B.n502 35.679
R1596 B.n808 B.n498 35.679
R1597 B.n814 B.n498 35.679
R1598 B.n814 B.n494 35.679
R1599 B.n821 B.n494 35.679
R1600 B.n821 B.n820 35.679
R1601 B.n827 B.n487 35.679
R1602 B.n833 B.n487 35.679
R1603 B.n833 B.n483 35.679
R1604 B.n839 B.n483 35.679
R1605 B.n839 B.n479 35.679
R1606 B.n845 B.n479 35.679
R1607 B.n845 B.n475 35.679
R1608 B.n851 B.n475 35.679
R1609 B.n851 B.n471 35.679
R1610 B.n857 B.n471 35.679
R1611 B.n857 B.n466 35.679
R1612 B.n863 B.n466 35.679
R1613 B.n863 B.n467 35.679
R1614 B.n869 B.n459 35.679
R1615 B.n875 B.n459 35.679
R1616 B.n875 B.n455 35.679
R1617 B.n881 B.n455 35.679
R1618 B.n881 B.n451 35.679
R1619 B.n887 B.n451 35.679
R1620 B.n887 B.n447 35.679
R1621 B.n894 B.n447 35.679
R1622 B.n894 B.n893 35.679
R1623 B.n900 B.n440 35.679
R1624 B.n906 B.n440 35.679
R1625 B.n906 B.n436 35.679
R1626 B.n912 B.n436 35.679
R1627 B.n912 B.n432 35.679
R1628 B.n918 B.n432 35.679
R1629 B.n918 B.n427 35.679
R1630 B.n924 B.n427 35.679
R1631 B.n924 B.n428 35.679
R1632 B.n930 B.n420 35.679
R1633 B.n936 B.n420 35.679
R1634 B.n936 B.n416 35.679
R1635 B.n942 B.n416 35.679
R1636 B.n942 B.n412 35.679
R1637 B.n948 B.n412 35.679
R1638 B.n948 B.n408 35.679
R1639 B.n955 B.n408 35.679
R1640 B.n955 B.n954 35.679
R1641 B.n961 B.n401 35.679
R1642 B.n968 B.n401 35.679
R1643 B.n968 B.n397 35.679
R1644 B.n974 B.n397 35.679
R1645 B.n974 B.n4 35.679
R1646 B.n1179 B.n4 35.679
R1647 B.n1179 B.n1178 35.679
R1648 B.n1178 B.n1177 35.679
R1649 B.n1177 B.n8 35.679
R1650 B.n12 B.n8 35.679
R1651 B.n1170 B.n12 35.679
R1652 B.n1170 B.n1169 35.679
R1653 B.n1169 B.n1168 35.679
R1654 B.n1162 B.n19 35.679
R1655 B.n1162 B.n1161 35.679
R1656 B.n1161 B.n1160 35.679
R1657 B.n1160 B.n23 35.679
R1658 B.n1154 B.n23 35.679
R1659 B.n1154 B.n1153 35.679
R1660 B.n1153 B.n1152 35.679
R1661 B.n1152 B.n30 35.679
R1662 B.n1146 B.n30 35.679
R1663 B.n1145 B.n1144 35.679
R1664 B.n1144 B.n37 35.679
R1665 B.n1138 B.n37 35.679
R1666 B.n1138 B.n1137 35.679
R1667 B.n1137 B.n1136 35.679
R1668 B.n1136 B.n44 35.679
R1669 B.n1130 B.n44 35.679
R1670 B.n1130 B.n1129 35.679
R1671 B.n1129 B.n1128 35.679
R1672 B.n1122 B.n54 35.679
R1673 B.n1122 B.n1121 35.679
R1674 B.n1121 B.n1120 35.679
R1675 B.n1120 B.n58 35.679
R1676 B.n1114 B.n58 35.679
R1677 B.n1114 B.n1113 35.679
R1678 B.n1113 B.n1112 35.679
R1679 B.n1112 B.n65 35.679
R1680 B.n1106 B.n65 35.679
R1681 B.n1105 B.n1104 35.679
R1682 B.n1104 B.n72 35.679
R1683 B.n1098 B.n72 35.679
R1684 B.n1098 B.n1097 35.679
R1685 B.n1097 B.n1096 35.679
R1686 B.n1096 B.n79 35.679
R1687 B.n1090 B.n79 35.679
R1688 B.n1090 B.n1089 35.679
R1689 B.n1089 B.n1088 35.679
R1690 B.n1088 B.n86 35.679
R1691 B.n1082 B.n86 35.679
R1692 B.n1082 B.n1081 35.679
R1693 B.n1081 B.n1080 35.679
R1694 B.n1074 B.n96 35.679
R1695 B.n1074 B.n1073 35.679
R1696 B.n1073 B.n1072 35.679
R1697 B.n1072 B.n100 35.679
R1698 B.n1066 B.n100 35.679
R1699 B.n1066 B.n1065 35.679
R1700 B.n1065 B.n1064 35.679
R1701 B.n1064 B.n107 35.679
R1702 B.n869 B.t5 33.0556
R1703 B.n1106 B.t7 33.0556
R1704 B.n799 B.n798 32.9371
R1705 B.n571 B.n504 32.9371
R1706 B.n1054 B.n1053 32.9371
R1707 B.n1061 B.n1060 32.9371
R1708 B.n954 B.t6 27.8088
R1709 B.n19 B.t1 27.8088
R1710 B.n900 B.t3 24.6606
R1711 B.n1128 B.t4 24.6606
R1712 B.n820 B.t9 22.5619
R1713 B.n96 B.t13 22.5619
R1714 B.n428 B.t0 19.4138
R1715 B.t2 B.n1145 19.4138
R1716 B B.n1182 18.0485
R1717 B.n930 B.t0 16.2657
R1718 B.n1146 B.t2 16.2657
R1719 B.n827 B.t9 13.1176
R1720 B.n1080 B.t13 13.1176
R1721 B.n893 B.t3 11.0189
R1722 B.n54 B.t4 11.0189
R1723 B.n800 B.n799 10.6151
R1724 B.n800 B.n500 10.6151
R1725 B.n810 B.n500 10.6151
R1726 B.n811 B.n810 10.6151
R1727 B.n812 B.n811 10.6151
R1728 B.n812 B.n492 10.6151
R1729 B.n823 B.n492 10.6151
R1730 B.n824 B.n823 10.6151
R1731 B.n825 B.n824 10.6151
R1732 B.n825 B.n485 10.6151
R1733 B.n835 B.n485 10.6151
R1734 B.n836 B.n835 10.6151
R1735 B.n837 B.n836 10.6151
R1736 B.n837 B.n477 10.6151
R1737 B.n847 B.n477 10.6151
R1738 B.n848 B.n847 10.6151
R1739 B.n849 B.n848 10.6151
R1740 B.n849 B.n469 10.6151
R1741 B.n859 B.n469 10.6151
R1742 B.n860 B.n859 10.6151
R1743 B.n861 B.n860 10.6151
R1744 B.n861 B.n461 10.6151
R1745 B.n871 B.n461 10.6151
R1746 B.n872 B.n871 10.6151
R1747 B.n873 B.n872 10.6151
R1748 B.n873 B.n453 10.6151
R1749 B.n883 B.n453 10.6151
R1750 B.n884 B.n883 10.6151
R1751 B.n885 B.n884 10.6151
R1752 B.n885 B.n445 10.6151
R1753 B.n896 B.n445 10.6151
R1754 B.n897 B.n896 10.6151
R1755 B.n898 B.n897 10.6151
R1756 B.n898 B.n438 10.6151
R1757 B.n908 B.n438 10.6151
R1758 B.n909 B.n908 10.6151
R1759 B.n910 B.n909 10.6151
R1760 B.n910 B.n430 10.6151
R1761 B.n920 B.n430 10.6151
R1762 B.n921 B.n920 10.6151
R1763 B.n922 B.n921 10.6151
R1764 B.n922 B.n422 10.6151
R1765 B.n932 B.n422 10.6151
R1766 B.n933 B.n932 10.6151
R1767 B.n934 B.n933 10.6151
R1768 B.n934 B.n414 10.6151
R1769 B.n944 B.n414 10.6151
R1770 B.n945 B.n944 10.6151
R1771 B.n946 B.n945 10.6151
R1772 B.n946 B.n406 10.6151
R1773 B.n957 B.n406 10.6151
R1774 B.n958 B.n957 10.6151
R1775 B.n959 B.n958 10.6151
R1776 B.n959 B.n399 10.6151
R1777 B.n970 B.n399 10.6151
R1778 B.n971 B.n970 10.6151
R1779 B.n972 B.n971 10.6151
R1780 B.n972 B.n0 10.6151
R1781 B.n798 B.n508 10.6151
R1782 B.n793 B.n508 10.6151
R1783 B.n793 B.n792 10.6151
R1784 B.n792 B.n791 10.6151
R1785 B.n791 B.n788 10.6151
R1786 B.n788 B.n787 10.6151
R1787 B.n787 B.n784 10.6151
R1788 B.n784 B.n783 10.6151
R1789 B.n783 B.n780 10.6151
R1790 B.n780 B.n779 10.6151
R1791 B.n779 B.n776 10.6151
R1792 B.n776 B.n775 10.6151
R1793 B.n775 B.n772 10.6151
R1794 B.n772 B.n771 10.6151
R1795 B.n771 B.n768 10.6151
R1796 B.n768 B.n767 10.6151
R1797 B.n767 B.n764 10.6151
R1798 B.n764 B.n763 10.6151
R1799 B.n763 B.n760 10.6151
R1800 B.n760 B.n759 10.6151
R1801 B.n759 B.n756 10.6151
R1802 B.n756 B.n755 10.6151
R1803 B.n755 B.n752 10.6151
R1804 B.n752 B.n751 10.6151
R1805 B.n751 B.n748 10.6151
R1806 B.n748 B.n747 10.6151
R1807 B.n747 B.n744 10.6151
R1808 B.n744 B.n743 10.6151
R1809 B.n743 B.n740 10.6151
R1810 B.n740 B.n739 10.6151
R1811 B.n739 B.n736 10.6151
R1812 B.n736 B.n735 10.6151
R1813 B.n735 B.n732 10.6151
R1814 B.n732 B.n731 10.6151
R1815 B.n731 B.n728 10.6151
R1816 B.n728 B.n727 10.6151
R1817 B.n727 B.n724 10.6151
R1818 B.n724 B.n723 10.6151
R1819 B.n723 B.n720 10.6151
R1820 B.n720 B.n719 10.6151
R1821 B.n719 B.n716 10.6151
R1822 B.n716 B.n715 10.6151
R1823 B.n715 B.n712 10.6151
R1824 B.n712 B.n711 10.6151
R1825 B.n711 B.n708 10.6151
R1826 B.n708 B.n707 10.6151
R1827 B.n707 B.n704 10.6151
R1828 B.n704 B.n703 10.6151
R1829 B.n703 B.n700 10.6151
R1830 B.n700 B.n699 10.6151
R1831 B.n699 B.n696 10.6151
R1832 B.n694 B.n691 10.6151
R1833 B.n691 B.n690 10.6151
R1834 B.n690 B.n687 10.6151
R1835 B.n687 B.n686 10.6151
R1836 B.n686 B.n683 10.6151
R1837 B.n683 B.n682 10.6151
R1838 B.n682 B.n679 10.6151
R1839 B.n679 B.n678 10.6151
R1840 B.n678 B.n675 10.6151
R1841 B.n673 B.n670 10.6151
R1842 B.n670 B.n669 10.6151
R1843 B.n669 B.n666 10.6151
R1844 B.n666 B.n665 10.6151
R1845 B.n665 B.n662 10.6151
R1846 B.n662 B.n661 10.6151
R1847 B.n661 B.n658 10.6151
R1848 B.n658 B.n657 10.6151
R1849 B.n657 B.n654 10.6151
R1850 B.n654 B.n653 10.6151
R1851 B.n653 B.n650 10.6151
R1852 B.n650 B.n649 10.6151
R1853 B.n649 B.n646 10.6151
R1854 B.n646 B.n645 10.6151
R1855 B.n645 B.n642 10.6151
R1856 B.n642 B.n641 10.6151
R1857 B.n641 B.n638 10.6151
R1858 B.n638 B.n637 10.6151
R1859 B.n637 B.n634 10.6151
R1860 B.n634 B.n633 10.6151
R1861 B.n633 B.n630 10.6151
R1862 B.n630 B.n629 10.6151
R1863 B.n629 B.n626 10.6151
R1864 B.n626 B.n625 10.6151
R1865 B.n625 B.n622 10.6151
R1866 B.n622 B.n621 10.6151
R1867 B.n621 B.n618 10.6151
R1868 B.n618 B.n617 10.6151
R1869 B.n617 B.n614 10.6151
R1870 B.n614 B.n613 10.6151
R1871 B.n613 B.n610 10.6151
R1872 B.n610 B.n609 10.6151
R1873 B.n609 B.n606 10.6151
R1874 B.n606 B.n605 10.6151
R1875 B.n605 B.n602 10.6151
R1876 B.n602 B.n601 10.6151
R1877 B.n601 B.n598 10.6151
R1878 B.n598 B.n597 10.6151
R1879 B.n597 B.n594 10.6151
R1880 B.n594 B.n593 10.6151
R1881 B.n593 B.n590 10.6151
R1882 B.n590 B.n589 10.6151
R1883 B.n589 B.n586 10.6151
R1884 B.n586 B.n585 10.6151
R1885 B.n585 B.n582 10.6151
R1886 B.n582 B.n581 10.6151
R1887 B.n581 B.n578 10.6151
R1888 B.n578 B.n577 10.6151
R1889 B.n577 B.n574 10.6151
R1890 B.n574 B.n573 10.6151
R1891 B.n573 B.n571 10.6151
R1892 B.n804 B.n504 10.6151
R1893 B.n805 B.n804 10.6151
R1894 B.n806 B.n805 10.6151
R1895 B.n806 B.n496 10.6151
R1896 B.n816 B.n496 10.6151
R1897 B.n817 B.n816 10.6151
R1898 B.n818 B.n817 10.6151
R1899 B.n818 B.n489 10.6151
R1900 B.n829 B.n489 10.6151
R1901 B.n830 B.n829 10.6151
R1902 B.n831 B.n830 10.6151
R1903 B.n831 B.n481 10.6151
R1904 B.n841 B.n481 10.6151
R1905 B.n842 B.n841 10.6151
R1906 B.n843 B.n842 10.6151
R1907 B.n843 B.n473 10.6151
R1908 B.n853 B.n473 10.6151
R1909 B.n854 B.n853 10.6151
R1910 B.n855 B.n854 10.6151
R1911 B.n855 B.n464 10.6151
R1912 B.n865 B.n464 10.6151
R1913 B.n866 B.n865 10.6151
R1914 B.n867 B.n866 10.6151
R1915 B.n867 B.n457 10.6151
R1916 B.n877 B.n457 10.6151
R1917 B.n878 B.n877 10.6151
R1918 B.n879 B.n878 10.6151
R1919 B.n879 B.n449 10.6151
R1920 B.n889 B.n449 10.6151
R1921 B.n890 B.n889 10.6151
R1922 B.n891 B.n890 10.6151
R1923 B.n891 B.n442 10.6151
R1924 B.n902 B.n442 10.6151
R1925 B.n903 B.n902 10.6151
R1926 B.n904 B.n903 10.6151
R1927 B.n904 B.n434 10.6151
R1928 B.n914 B.n434 10.6151
R1929 B.n915 B.n914 10.6151
R1930 B.n916 B.n915 10.6151
R1931 B.n916 B.n425 10.6151
R1932 B.n926 B.n425 10.6151
R1933 B.n927 B.n926 10.6151
R1934 B.n928 B.n927 10.6151
R1935 B.n928 B.n418 10.6151
R1936 B.n938 B.n418 10.6151
R1937 B.n939 B.n938 10.6151
R1938 B.n940 B.n939 10.6151
R1939 B.n940 B.n410 10.6151
R1940 B.n950 B.n410 10.6151
R1941 B.n951 B.n950 10.6151
R1942 B.n952 B.n951 10.6151
R1943 B.n952 B.n403 10.6151
R1944 B.n963 B.n403 10.6151
R1945 B.n964 B.n963 10.6151
R1946 B.n966 B.n964 10.6151
R1947 B.n966 B.n965 10.6151
R1948 B.n965 B.n395 10.6151
R1949 B.n977 B.n395 10.6151
R1950 B.n978 B.n977 10.6151
R1951 B.n979 B.n978 10.6151
R1952 B.n980 B.n979 10.6151
R1953 B.n981 B.n980 10.6151
R1954 B.n984 B.n981 10.6151
R1955 B.n985 B.n984 10.6151
R1956 B.n986 B.n985 10.6151
R1957 B.n987 B.n986 10.6151
R1958 B.n989 B.n987 10.6151
R1959 B.n990 B.n989 10.6151
R1960 B.n991 B.n990 10.6151
R1961 B.n992 B.n991 10.6151
R1962 B.n994 B.n992 10.6151
R1963 B.n995 B.n994 10.6151
R1964 B.n996 B.n995 10.6151
R1965 B.n997 B.n996 10.6151
R1966 B.n999 B.n997 10.6151
R1967 B.n1000 B.n999 10.6151
R1968 B.n1001 B.n1000 10.6151
R1969 B.n1002 B.n1001 10.6151
R1970 B.n1004 B.n1002 10.6151
R1971 B.n1005 B.n1004 10.6151
R1972 B.n1006 B.n1005 10.6151
R1973 B.n1007 B.n1006 10.6151
R1974 B.n1009 B.n1007 10.6151
R1975 B.n1010 B.n1009 10.6151
R1976 B.n1011 B.n1010 10.6151
R1977 B.n1012 B.n1011 10.6151
R1978 B.n1014 B.n1012 10.6151
R1979 B.n1015 B.n1014 10.6151
R1980 B.n1016 B.n1015 10.6151
R1981 B.n1017 B.n1016 10.6151
R1982 B.n1019 B.n1017 10.6151
R1983 B.n1020 B.n1019 10.6151
R1984 B.n1021 B.n1020 10.6151
R1985 B.n1022 B.n1021 10.6151
R1986 B.n1024 B.n1022 10.6151
R1987 B.n1025 B.n1024 10.6151
R1988 B.n1026 B.n1025 10.6151
R1989 B.n1027 B.n1026 10.6151
R1990 B.n1029 B.n1027 10.6151
R1991 B.n1030 B.n1029 10.6151
R1992 B.n1031 B.n1030 10.6151
R1993 B.n1032 B.n1031 10.6151
R1994 B.n1034 B.n1032 10.6151
R1995 B.n1035 B.n1034 10.6151
R1996 B.n1036 B.n1035 10.6151
R1997 B.n1037 B.n1036 10.6151
R1998 B.n1039 B.n1037 10.6151
R1999 B.n1040 B.n1039 10.6151
R2000 B.n1041 B.n1040 10.6151
R2001 B.n1042 B.n1041 10.6151
R2002 B.n1044 B.n1042 10.6151
R2003 B.n1045 B.n1044 10.6151
R2004 B.n1046 B.n1045 10.6151
R2005 B.n1047 B.n1046 10.6151
R2006 B.n1049 B.n1047 10.6151
R2007 B.n1050 B.n1049 10.6151
R2008 B.n1051 B.n1050 10.6151
R2009 B.n1052 B.n1051 10.6151
R2010 B.n1053 B.n1052 10.6151
R2011 B.n1174 B.n1 10.6151
R2012 B.n1174 B.n1173 10.6151
R2013 B.n1173 B.n1172 10.6151
R2014 B.n1172 B.n10 10.6151
R2015 B.n1166 B.n10 10.6151
R2016 B.n1166 B.n1165 10.6151
R2017 B.n1165 B.n1164 10.6151
R2018 B.n1164 B.n17 10.6151
R2019 B.n1158 B.n17 10.6151
R2020 B.n1158 B.n1157 10.6151
R2021 B.n1157 B.n1156 10.6151
R2022 B.n1156 B.n25 10.6151
R2023 B.n1150 B.n25 10.6151
R2024 B.n1150 B.n1149 10.6151
R2025 B.n1149 B.n1148 10.6151
R2026 B.n1148 B.n32 10.6151
R2027 B.n1142 B.n32 10.6151
R2028 B.n1142 B.n1141 10.6151
R2029 B.n1141 B.n1140 10.6151
R2030 B.n1140 B.n39 10.6151
R2031 B.n1134 B.n39 10.6151
R2032 B.n1134 B.n1133 10.6151
R2033 B.n1133 B.n1132 10.6151
R2034 B.n1132 B.n46 10.6151
R2035 B.n1126 B.n46 10.6151
R2036 B.n1126 B.n1125 10.6151
R2037 B.n1125 B.n1124 10.6151
R2038 B.n1124 B.n52 10.6151
R2039 B.n1118 B.n52 10.6151
R2040 B.n1118 B.n1117 10.6151
R2041 B.n1117 B.n1116 10.6151
R2042 B.n1116 B.n60 10.6151
R2043 B.n1110 B.n60 10.6151
R2044 B.n1110 B.n1109 10.6151
R2045 B.n1109 B.n1108 10.6151
R2046 B.n1108 B.n67 10.6151
R2047 B.n1102 B.n67 10.6151
R2048 B.n1102 B.n1101 10.6151
R2049 B.n1101 B.n1100 10.6151
R2050 B.n1100 B.n74 10.6151
R2051 B.n1094 B.n74 10.6151
R2052 B.n1094 B.n1093 10.6151
R2053 B.n1093 B.n1092 10.6151
R2054 B.n1092 B.n81 10.6151
R2055 B.n1086 B.n81 10.6151
R2056 B.n1086 B.n1085 10.6151
R2057 B.n1085 B.n1084 10.6151
R2058 B.n1084 B.n88 10.6151
R2059 B.n1078 B.n88 10.6151
R2060 B.n1078 B.n1077 10.6151
R2061 B.n1077 B.n1076 10.6151
R2062 B.n1076 B.n94 10.6151
R2063 B.n1070 B.n94 10.6151
R2064 B.n1070 B.n1069 10.6151
R2065 B.n1069 B.n1068 10.6151
R2066 B.n1068 B.n102 10.6151
R2067 B.n1062 B.n102 10.6151
R2068 B.n1062 B.n1061 10.6151
R2069 B.n1060 B.n109 10.6151
R2070 B.n175 B.n109 10.6151
R2071 B.n176 B.n175 10.6151
R2072 B.n179 B.n176 10.6151
R2073 B.n180 B.n179 10.6151
R2074 B.n183 B.n180 10.6151
R2075 B.n184 B.n183 10.6151
R2076 B.n187 B.n184 10.6151
R2077 B.n188 B.n187 10.6151
R2078 B.n191 B.n188 10.6151
R2079 B.n192 B.n191 10.6151
R2080 B.n195 B.n192 10.6151
R2081 B.n196 B.n195 10.6151
R2082 B.n199 B.n196 10.6151
R2083 B.n200 B.n199 10.6151
R2084 B.n203 B.n200 10.6151
R2085 B.n204 B.n203 10.6151
R2086 B.n207 B.n204 10.6151
R2087 B.n208 B.n207 10.6151
R2088 B.n211 B.n208 10.6151
R2089 B.n212 B.n211 10.6151
R2090 B.n215 B.n212 10.6151
R2091 B.n216 B.n215 10.6151
R2092 B.n219 B.n216 10.6151
R2093 B.n220 B.n219 10.6151
R2094 B.n223 B.n220 10.6151
R2095 B.n224 B.n223 10.6151
R2096 B.n227 B.n224 10.6151
R2097 B.n228 B.n227 10.6151
R2098 B.n231 B.n228 10.6151
R2099 B.n232 B.n231 10.6151
R2100 B.n235 B.n232 10.6151
R2101 B.n236 B.n235 10.6151
R2102 B.n239 B.n236 10.6151
R2103 B.n240 B.n239 10.6151
R2104 B.n243 B.n240 10.6151
R2105 B.n244 B.n243 10.6151
R2106 B.n247 B.n244 10.6151
R2107 B.n248 B.n247 10.6151
R2108 B.n251 B.n248 10.6151
R2109 B.n252 B.n251 10.6151
R2110 B.n255 B.n252 10.6151
R2111 B.n256 B.n255 10.6151
R2112 B.n259 B.n256 10.6151
R2113 B.n260 B.n259 10.6151
R2114 B.n263 B.n260 10.6151
R2115 B.n264 B.n263 10.6151
R2116 B.n267 B.n264 10.6151
R2117 B.n268 B.n267 10.6151
R2118 B.n271 B.n268 10.6151
R2119 B.n272 B.n271 10.6151
R2120 B.n276 B.n275 10.6151
R2121 B.n279 B.n276 10.6151
R2122 B.n280 B.n279 10.6151
R2123 B.n283 B.n280 10.6151
R2124 B.n284 B.n283 10.6151
R2125 B.n287 B.n284 10.6151
R2126 B.n288 B.n287 10.6151
R2127 B.n291 B.n288 10.6151
R2128 B.n292 B.n291 10.6151
R2129 B.n296 B.n295 10.6151
R2130 B.n299 B.n296 10.6151
R2131 B.n300 B.n299 10.6151
R2132 B.n303 B.n300 10.6151
R2133 B.n304 B.n303 10.6151
R2134 B.n307 B.n304 10.6151
R2135 B.n308 B.n307 10.6151
R2136 B.n311 B.n308 10.6151
R2137 B.n312 B.n311 10.6151
R2138 B.n315 B.n312 10.6151
R2139 B.n316 B.n315 10.6151
R2140 B.n319 B.n316 10.6151
R2141 B.n320 B.n319 10.6151
R2142 B.n323 B.n320 10.6151
R2143 B.n324 B.n323 10.6151
R2144 B.n327 B.n324 10.6151
R2145 B.n328 B.n327 10.6151
R2146 B.n331 B.n328 10.6151
R2147 B.n332 B.n331 10.6151
R2148 B.n335 B.n332 10.6151
R2149 B.n336 B.n335 10.6151
R2150 B.n339 B.n336 10.6151
R2151 B.n340 B.n339 10.6151
R2152 B.n343 B.n340 10.6151
R2153 B.n344 B.n343 10.6151
R2154 B.n347 B.n344 10.6151
R2155 B.n348 B.n347 10.6151
R2156 B.n351 B.n348 10.6151
R2157 B.n352 B.n351 10.6151
R2158 B.n355 B.n352 10.6151
R2159 B.n356 B.n355 10.6151
R2160 B.n359 B.n356 10.6151
R2161 B.n360 B.n359 10.6151
R2162 B.n363 B.n360 10.6151
R2163 B.n364 B.n363 10.6151
R2164 B.n367 B.n364 10.6151
R2165 B.n368 B.n367 10.6151
R2166 B.n371 B.n368 10.6151
R2167 B.n372 B.n371 10.6151
R2168 B.n375 B.n372 10.6151
R2169 B.n376 B.n375 10.6151
R2170 B.n379 B.n376 10.6151
R2171 B.n380 B.n379 10.6151
R2172 B.n383 B.n380 10.6151
R2173 B.n384 B.n383 10.6151
R2174 B.n387 B.n384 10.6151
R2175 B.n388 B.n387 10.6151
R2176 B.n391 B.n388 10.6151
R2177 B.n393 B.n391 10.6151
R2178 B.n394 B.n393 10.6151
R2179 B.n1054 B.n394 10.6151
R2180 B.n696 B.n695 9.36635
R2181 B.n674 B.n673 9.36635
R2182 B.n272 B.n173 9.36635
R2183 B.n295 B.n170 9.36635
R2184 B.n1182 B.n0 8.11757
R2185 B.n1182 B.n1 8.11757
R2186 B.n961 B.t6 7.87076
R2187 B.n1168 B.t1 7.87076
R2188 B.n467 B.t5 2.62392
R2189 B.t7 B.n1105 2.62392
R2190 B.n695 B.n694 1.24928
R2191 B.n675 B.n674 1.24928
R2192 B.n275 B.n173 1.24928
R2193 B.n292 B.n170 1.24928
R2194 VN.n60 VN.n59 161.3
R2195 VN.n58 VN.n32 161.3
R2196 VN.n57 VN.n56 161.3
R2197 VN.n55 VN.n33 161.3
R2198 VN.n54 VN.n53 161.3
R2199 VN.n52 VN.n34 161.3
R2200 VN.n51 VN.n50 161.3
R2201 VN.n49 VN.n48 161.3
R2202 VN.n47 VN.n36 161.3
R2203 VN.n46 VN.n45 161.3
R2204 VN.n44 VN.n37 161.3
R2205 VN.n43 VN.n42 161.3
R2206 VN.n41 VN.n38 161.3
R2207 VN.n29 VN.n28 161.3
R2208 VN.n27 VN.n1 161.3
R2209 VN.n26 VN.n25 161.3
R2210 VN.n24 VN.n2 161.3
R2211 VN.n23 VN.n22 161.3
R2212 VN.n21 VN.n3 161.3
R2213 VN.n20 VN.n19 161.3
R2214 VN.n18 VN.n17 161.3
R2215 VN.n16 VN.n5 161.3
R2216 VN.n15 VN.n14 161.3
R2217 VN.n13 VN.n6 161.3
R2218 VN.n12 VN.n11 161.3
R2219 VN.n10 VN.n7 161.3
R2220 VN.n39 VN.t3 153.446
R2221 VN.n8 VN.t4 153.446
R2222 VN.n9 VN.t2 120.041
R2223 VN.n4 VN.t7 120.041
R2224 VN.n0 VN.t5 120.041
R2225 VN.n40 VN.t6 120.041
R2226 VN.n35 VN.t1 120.041
R2227 VN.n31 VN.t0 120.041
R2228 VN.n30 VN.n0 67.0684
R2229 VN.n61 VN.n31 67.0684
R2230 VN VN.n61 56.6344
R2231 VN.n15 VN.n6 56.5193
R2232 VN.n26 VN.n2 56.5193
R2233 VN.n46 VN.n37 56.5193
R2234 VN.n57 VN.n33 56.5193
R2235 VN.n40 VN.n39 50.0328
R2236 VN.n9 VN.n8 50.0328
R2237 VN.n11 VN.n10 24.4675
R2238 VN.n11 VN.n6 24.4675
R2239 VN.n16 VN.n15 24.4675
R2240 VN.n17 VN.n16 24.4675
R2241 VN.n21 VN.n20 24.4675
R2242 VN.n22 VN.n21 24.4675
R2243 VN.n22 VN.n2 24.4675
R2244 VN.n27 VN.n26 24.4675
R2245 VN.n28 VN.n27 24.4675
R2246 VN.n42 VN.n37 24.4675
R2247 VN.n42 VN.n41 24.4675
R2248 VN.n53 VN.n33 24.4675
R2249 VN.n53 VN.n52 24.4675
R2250 VN.n52 VN.n51 24.4675
R2251 VN.n48 VN.n47 24.4675
R2252 VN.n47 VN.n46 24.4675
R2253 VN.n59 VN.n58 24.4675
R2254 VN.n58 VN.n57 24.4675
R2255 VN.n10 VN.n9 23.9782
R2256 VN.n17 VN.n4 23.9782
R2257 VN.n41 VN.n40 23.9782
R2258 VN.n48 VN.n35 23.9782
R2259 VN.n28 VN.n0 22.9995
R2260 VN.n59 VN.n31 22.9995
R2261 VN.n39 VN.n38 3.77031
R2262 VN.n8 VN.n7 3.77031
R2263 VN.n20 VN.n4 0.48984
R2264 VN.n51 VN.n35 0.48984
R2265 VN.n61 VN.n60 0.354971
R2266 VN.n30 VN.n29 0.354971
R2267 VN VN.n30 0.26696
R2268 VN.n60 VN.n32 0.189894
R2269 VN.n56 VN.n32 0.189894
R2270 VN.n56 VN.n55 0.189894
R2271 VN.n55 VN.n54 0.189894
R2272 VN.n54 VN.n34 0.189894
R2273 VN.n50 VN.n34 0.189894
R2274 VN.n50 VN.n49 0.189894
R2275 VN.n49 VN.n36 0.189894
R2276 VN.n45 VN.n36 0.189894
R2277 VN.n45 VN.n44 0.189894
R2278 VN.n44 VN.n43 0.189894
R2279 VN.n43 VN.n38 0.189894
R2280 VN.n12 VN.n7 0.189894
R2281 VN.n13 VN.n12 0.189894
R2282 VN.n14 VN.n13 0.189894
R2283 VN.n14 VN.n5 0.189894
R2284 VN.n18 VN.n5 0.189894
R2285 VN.n19 VN.n18 0.189894
R2286 VN.n19 VN.n3 0.189894
R2287 VN.n23 VN.n3 0.189894
R2288 VN.n24 VN.n23 0.189894
R2289 VN.n25 VN.n24 0.189894
R2290 VN.n25 VN.n1 0.189894
R2291 VN.n29 VN.n1 0.189894
R2292 VDD2.n2 VDD2.n1 61.6709
R2293 VDD2.n2 VDD2.n0 61.6709
R2294 VDD2 VDD2.n5 61.6681
R2295 VDD2.n4 VDD2.n3 60.2265
R2296 VDD2.n4 VDD2.n2 50.7412
R2297 VDD2 VDD2.n4 1.55869
R2298 VDD2.n5 VDD2.t1 1.26245
R2299 VDD2.n5 VDD2.t4 1.26245
R2300 VDD2.n3 VDD2.t7 1.26245
R2301 VDD2.n3 VDD2.t6 1.26245
R2302 VDD2.n1 VDD2.t0 1.26245
R2303 VDD2.n1 VDD2.t2 1.26245
R2304 VDD2.n0 VDD2.t3 1.26245
R2305 VDD2.n0 VDD2.t5 1.26245
C0 VDD1 VN 0.152847f
C1 VTAIL VP 12.0482f
C2 VDD1 VP 12.044f
C3 VN VP 9.01639f
C4 VTAIL VDD2 9.43462f
C5 VDD1 VDD2 2.0648f
C6 VN VDD2 11.6202f
C7 VDD2 VP 0.578322f
C8 VTAIL VDD1 9.376519f
C9 VTAIL VN 12.0341f
C10 VDD2 B 6.230631f
C11 VDD1 B 6.727162f
C12 VTAIL B 13.088223f
C13 VN B 17.90807f
C14 VP B 16.499443f
C15 VDD2.t3 B 0.328458f
C16 VDD2.t5 B 0.328458f
C17 VDD2.n0 B 2.98842f
C18 VDD2.t0 B 0.328458f
C19 VDD2.t2 B 0.328458f
C20 VDD2.n1 B 2.98842f
C21 VDD2.n2 B 4.058f
C22 VDD2.t7 B 0.328458f
C23 VDD2.t6 B 0.328458f
C24 VDD2.n3 B 2.97415f
C25 VDD2.n4 B 3.62469f
C26 VDD2.t1 B 0.328458f
C27 VDD2.t4 B 0.328458f
C28 VDD2.n5 B 2.98837f
C29 VN.t5 B 2.55232f
C30 VN.n0 B 0.968442f
C31 VN.n1 B 0.018827f
C32 VN.n2 B 0.026435f
C33 VN.n3 B 0.018827f
C34 VN.t7 B 2.55232f
C35 VN.n4 B 0.886566f
C36 VN.n5 B 0.018827f
C37 VN.n6 B 0.027484f
C38 VN.n7 B 0.214174f
C39 VN.t2 B 2.55232f
C40 VN.t4 B 2.7754f
C41 VN.n8 B 0.914128f
C42 VN.n9 B 0.957531f
C43 VN.n10 B 0.034743f
C44 VN.n11 B 0.035089f
C45 VN.n12 B 0.018827f
C46 VN.n13 B 0.018827f
C47 VN.n14 B 0.018827f
C48 VN.n15 B 0.027484f
C49 VN.n16 B 0.035089f
C50 VN.n17 B 0.034743f
C51 VN.n18 B 0.018827f
C52 VN.n19 B 0.018827f
C53 VN.n20 B 0.018112f
C54 VN.n21 B 0.035089f
C55 VN.n22 B 0.035089f
C56 VN.n23 B 0.018827f
C57 VN.n24 B 0.018827f
C58 VN.n25 B 0.018827f
C59 VN.n26 B 0.028534f
C60 VN.n27 B 0.035089f
C61 VN.n28 B 0.03405f
C62 VN.n29 B 0.030387f
C63 VN.n30 B 0.037228f
C64 VN.t0 B 2.55232f
C65 VN.n31 B 0.968442f
C66 VN.n32 B 0.018827f
C67 VN.n33 B 0.026435f
C68 VN.n34 B 0.018827f
C69 VN.t1 B 2.55232f
C70 VN.n35 B 0.886566f
C71 VN.n36 B 0.018827f
C72 VN.n37 B 0.027484f
C73 VN.n38 B 0.214174f
C74 VN.t6 B 2.55232f
C75 VN.t3 B 2.7754f
C76 VN.n39 B 0.914128f
C77 VN.n40 B 0.957531f
C78 VN.n41 B 0.034743f
C79 VN.n42 B 0.035089f
C80 VN.n43 B 0.018827f
C81 VN.n44 B 0.018827f
C82 VN.n45 B 0.018827f
C83 VN.n46 B 0.027484f
C84 VN.n47 B 0.035089f
C85 VN.n48 B 0.034743f
C86 VN.n49 B 0.018827f
C87 VN.n50 B 0.018827f
C88 VN.n51 B 0.018112f
C89 VN.n52 B 0.035089f
C90 VN.n53 B 0.035089f
C91 VN.n54 B 0.018827f
C92 VN.n55 B 0.018827f
C93 VN.n56 B 0.018827f
C94 VN.n57 B 0.028534f
C95 VN.n58 B 0.035089f
C96 VN.n59 B 0.03405f
C97 VN.n60 B 0.030387f
C98 VN.n61 B 1.27044f
C99 VTAIL.t2 B 0.238212f
C100 VTAIL.t4 B 0.238212f
C101 VTAIL.n0 B 2.09767f
C102 VTAIL.n1 B 0.381057f
C103 VTAIL.t1 B 2.67667f
C104 VTAIL.n2 B 0.477213f
C105 VTAIL.t10 B 2.67667f
C106 VTAIL.n3 B 0.477213f
C107 VTAIL.t9 B 0.238212f
C108 VTAIL.t11 B 0.238212f
C109 VTAIL.n4 B 2.09767f
C110 VTAIL.n5 B 0.563178f
C111 VTAIL.t13 B 2.67667f
C112 VTAIL.n6 B 1.73218f
C113 VTAIL.t5 B 2.67669f
C114 VTAIL.n7 B 1.73217f
C115 VTAIL.t3 B 0.238212f
C116 VTAIL.t0 B 0.238212f
C117 VTAIL.n8 B 2.09767f
C118 VTAIL.n9 B 0.563175f
C119 VTAIL.t6 B 2.67669f
C120 VTAIL.n10 B 0.477195f
C121 VTAIL.t8 B 2.67669f
C122 VTAIL.n11 B 0.477195f
C123 VTAIL.t14 B 0.238212f
C124 VTAIL.t15 B 0.238212f
C125 VTAIL.n12 B 2.09767f
C126 VTAIL.n13 B 0.563175f
C127 VTAIL.t12 B 2.67667f
C128 VTAIL.n14 B 1.73218f
C129 VTAIL.t7 B 2.67667f
C130 VTAIL.n15 B 1.72858f
C131 VDD1.t2 B 0.332737f
C132 VDD1.t0 B 0.332737f
C133 VDD1.n0 B 3.02869f
C134 VDD1.t5 B 0.332737f
C135 VDD1.t3 B 0.332737f
C136 VDD1.n1 B 3.02735f
C137 VDD1.t7 B 0.332737f
C138 VDD1.t6 B 0.332737f
C139 VDD1.n2 B 3.02735f
C140 VDD1.n3 B 4.16629f
C141 VDD1.t1 B 0.332737f
C142 VDD1.t4 B 0.332737f
C143 VDD1.n4 B 3.01288f
C144 VDD1.n5 B 3.70553f
C145 VP.t5 B 2.58574f
C146 VP.n0 B 0.981121f
C147 VP.n1 B 0.019074f
C148 VP.n2 B 0.026781f
C149 VP.n3 B 0.019074f
C150 VP.t4 B 2.58574f
C151 VP.n4 B 0.898173f
C152 VP.n5 B 0.019074f
C153 VP.n6 B 0.027844f
C154 VP.n7 B 0.019074f
C155 VP.t6 B 2.58574f
C156 VP.n8 B 0.035549f
C157 VP.n9 B 0.019074f
C158 VP.n10 B 0.035549f
C159 VP.t3 B 2.58574f
C160 VP.n11 B 0.981121f
C161 VP.n12 B 0.019074f
C162 VP.n13 B 0.026781f
C163 VP.n14 B 0.019074f
C164 VP.t0 B 2.58574f
C165 VP.n15 B 0.898173f
C166 VP.n16 B 0.019074f
C167 VP.n17 B 0.027844f
C168 VP.n18 B 0.216978f
C169 VP.t1 B 2.58574f
C170 VP.t7 B 2.81173f
C171 VP.n19 B 0.926097f
C172 VP.n20 B 0.970068f
C173 VP.n21 B 0.035198f
C174 VP.n22 B 0.035549f
C175 VP.n23 B 0.019074f
C176 VP.n24 B 0.019074f
C177 VP.n25 B 0.019074f
C178 VP.n26 B 0.027844f
C179 VP.n27 B 0.035549f
C180 VP.n28 B 0.035198f
C181 VP.n29 B 0.019074f
C182 VP.n30 B 0.019074f
C183 VP.n31 B 0.018349f
C184 VP.n32 B 0.035549f
C185 VP.n33 B 0.035549f
C186 VP.n34 B 0.019074f
C187 VP.n35 B 0.019074f
C188 VP.n36 B 0.019074f
C189 VP.n37 B 0.028907f
C190 VP.n38 B 0.035549f
C191 VP.n39 B 0.034496f
C192 VP.n40 B 0.030785f
C193 VP.n41 B 1.27958f
C194 VP.n42 B 1.29172f
C195 VP.t2 B 2.58574f
C196 VP.n43 B 0.981121f
C197 VP.n44 B 0.034496f
C198 VP.n45 B 0.030785f
C199 VP.n46 B 0.019074f
C200 VP.n47 B 0.019074f
C201 VP.n48 B 0.028907f
C202 VP.n49 B 0.026781f
C203 VP.n50 B 0.035549f
C204 VP.n51 B 0.019074f
C205 VP.n52 B 0.019074f
C206 VP.n53 B 0.019074f
C207 VP.n54 B 0.018349f
C208 VP.n55 B 0.898173f
C209 VP.n56 B 0.035198f
C210 VP.n57 B 0.035549f
C211 VP.n58 B 0.019074f
C212 VP.n59 B 0.019074f
C213 VP.n60 B 0.019074f
C214 VP.n61 B 0.027844f
C215 VP.n62 B 0.035549f
C216 VP.n63 B 0.035198f
C217 VP.n64 B 0.019074f
C218 VP.n65 B 0.019074f
C219 VP.n66 B 0.018349f
C220 VP.n67 B 0.035549f
C221 VP.n68 B 0.035549f
C222 VP.n69 B 0.019074f
C223 VP.n70 B 0.019074f
C224 VP.n71 B 0.019074f
C225 VP.n72 B 0.028907f
C226 VP.n73 B 0.035549f
C227 VP.n74 B 0.034496f
C228 VP.n75 B 0.030785f
C229 VP.n76 B 0.037716f
.ends

