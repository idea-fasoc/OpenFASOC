* NGSPICE file created from diff_pair_sample_0280.ext - technology: sky130A

.subckt diff_pair_sample_0280 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.7524 pd=4.89 as=1.7784 ps=9.9 w=4.56 l=2.54
X1 VTAIL.t3 VN.t0 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.7784 pd=9.9 as=0.7524 ps=4.89 w=4.56 l=2.54
X2 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=1.7784 pd=9.9 as=0 ps=0 w=4.56 l=2.54
X3 VTAIL.t0 VN.t1 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.7784 pd=9.9 as=0.7524 ps=4.89 w=4.56 l=2.54
X4 VTAIL.t5 VP.t1 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.7784 pd=9.9 as=0.7524 ps=4.89 w=4.56 l=2.54
X5 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=1.7784 pd=9.9 as=0 ps=0 w=4.56 l=2.54
X6 VDD1.t1 VP.t2 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7524 pd=4.89 as=1.7784 ps=9.9 w=4.56 l=2.54
X7 VTAIL.t4 VP.t3 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.7784 pd=9.9 as=0.7524 ps=4.89 w=4.56 l=2.54
X8 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.7784 pd=9.9 as=0 ps=0 w=4.56 l=2.54
X9 VDD2.t1 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7524 pd=4.89 as=1.7784 ps=9.9 w=4.56 l=2.54
X10 VDD2.t0 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.7524 pd=4.89 as=1.7784 ps=9.9 w=4.56 l=2.54
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.7784 pd=9.9 as=0 ps=0 w=4.56 l=2.54
R0 VP.n14 VP.n0 161.3
R1 VP.n13 VP.n12 161.3
R2 VP.n11 VP.n1 161.3
R3 VP.n10 VP.n9 161.3
R4 VP.n8 VP.n2 161.3
R5 VP.n7 VP.n6 161.3
R6 VP.n5 VP.n3 101.809
R7 VP.n16 VP.n15 101.809
R8 VP.n4 VP.t1 79.0883
R9 VP.n4 VP.t0 78.3227
R10 VP.n9 VP.n1 56.5617
R11 VP.n5 VP.n4 44.9031
R12 VP.n3 VP.t3 43.2666
R13 VP.n15 VP.t2 43.2666
R14 VP.n8 VP.n7 24.5923
R15 VP.n9 VP.n8 24.5923
R16 VP.n13 VP.n1 24.5923
R17 VP.n14 VP.n13 24.5923
R18 VP.n7 VP.n3 9.09948
R19 VP.n15 VP.n14 9.09948
R20 VP.n6 VP.n5 0.278335
R21 VP.n16 VP.n0 0.278335
R22 VP.n6 VP.n2 0.189894
R23 VP.n10 VP.n2 0.189894
R24 VP.n11 VP.n10 0.189894
R25 VP.n12 VP.n11 0.189894
R26 VP.n12 VP.n0 0.189894
R27 VP VP.n16 0.153485
R28 VTAIL.n186 VTAIL.n168 289.615
R29 VTAIL.n18 VTAIL.n0 289.615
R30 VTAIL.n42 VTAIL.n24 289.615
R31 VTAIL.n66 VTAIL.n48 289.615
R32 VTAIL.n162 VTAIL.n144 289.615
R33 VTAIL.n138 VTAIL.n120 289.615
R34 VTAIL.n114 VTAIL.n96 289.615
R35 VTAIL.n90 VTAIL.n72 289.615
R36 VTAIL.n177 VTAIL.n176 185
R37 VTAIL.n179 VTAIL.n178 185
R38 VTAIL.n172 VTAIL.n171 185
R39 VTAIL.n185 VTAIL.n184 185
R40 VTAIL.n187 VTAIL.n186 185
R41 VTAIL.n9 VTAIL.n8 185
R42 VTAIL.n11 VTAIL.n10 185
R43 VTAIL.n4 VTAIL.n3 185
R44 VTAIL.n17 VTAIL.n16 185
R45 VTAIL.n19 VTAIL.n18 185
R46 VTAIL.n33 VTAIL.n32 185
R47 VTAIL.n35 VTAIL.n34 185
R48 VTAIL.n28 VTAIL.n27 185
R49 VTAIL.n41 VTAIL.n40 185
R50 VTAIL.n43 VTAIL.n42 185
R51 VTAIL.n57 VTAIL.n56 185
R52 VTAIL.n59 VTAIL.n58 185
R53 VTAIL.n52 VTAIL.n51 185
R54 VTAIL.n65 VTAIL.n64 185
R55 VTAIL.n67 VTAIL.n66 185
R56 VTAIL.n163 VTAIL.n162 185
R57 VTAIL.n161 VTAIL.n160 185
R58 VTAIL.n148 VTAIL.n147 185
R59 VTAIL.n155 VTAIL.n154 185
R60 VTAIL.n153 VTAIL.n152 185
R61 VTAIL.n139 VTAIL.n138 185
R62 VTAIL.n137 VTAIL.n136 185
R63 VTAIL.n124 VTAIL.n123 185
R64 VTAIL.n131 VTAIL.n130 185
R65 VTAIL.n129 VTAIL.n128 185
R66 VTAIL.n115 VTAIL.n114 185
R67 VTAIL.n113 VTAIL.n112 185
R68 VTAIL.n100 VTAIL.n99 185
R69 VTAIL.n107 VTAIL.n106 185
R70 VTAIL.n105 VTAIL.n104 185
R71 VTAIL.n91 VTAIL.n90 185
R72 VTAIL.n89 VTAIL.n88 185
R73 VTAIL.n76 VTAIL.n75 185
R74 VTAIL.n83 VTAIL.n82 185
R75 VTAIL.n81 VTAIL.n80 185
R76 VTAIL.n175 VTAIL.t2 147.714
R77 VTAIL.n7 VTAIL.t3 147.714
R78 VTAIL.n31 VTAIL.t7 147.714
R79 VTAIL.n55 VTAIL.t4 147.714
R80 VTAIL.n151 VTAIL.t6 147.714
R81 VTAIL.n127 VTAIL.t5 147.714
R82 VTAIL.n103 VTAIL.t1 147.714
R83 VTAIL.n79 VTAIL.t0 147.714
R84 VTAIL.n178 VTAIL.n177 104.615
R85 VTAIL.n178 VTAIL.n171 104.615
R86 VTAIL.n185 VTAIL.n171 104.615
R87 VTAIL.n186 VTAIL.n185 104.615
R88 VTAIL.n10 VTAIL.n9 104.615
R89 VTAIL.n10 VTAIL.n3 104.615
R90 VTAIL.n17 VTAIL.n3 104.615
R91 VTAIL.n18 VTAIL.n17 104.615
R92 VTAIL.n34 VTAIL.n33 104.615
R93 VTAIL.n34 VTAIL.n27 104.615
R94 VTAIL.n41 VTAIL.n27 104.615
R95 VTAIL.n42 VTAIL.n41 104.615
R96 VTAIL.n58 VTAIL.n57 104.615
R97 VTAIL.n58 VTAIL.n51 104.615
R98 VTAIL.n65 VTAIL.n51 104.615
R99 VTAIL.n66 VTAIL.n65 104.615
R100 VTAIL.n162 VTAIL.n161 104.615
R101 VTAIL.n161 VTAIL.n147 104.615
R102 VTAIL.n154 VTAIL.n147 104.615
R103 VTAIL.n154 VTAIL.n153 104.615
R104 VTAIL.n138 VTAIL.n137 104.615
R105 VTAIL.n137 VTAIL.n123 104.615
R106 VTAIL.n130 VTAIL.n123 104.615
R107 VTAIL.n130 VTAIL.n129 104.615
R108 VTAIL.n114 VTAIL.n113 104.615
R109 VTAIL.n113 VTAIL.n99 104.615
R110 VTAIL.n106 VTAIL.n99 104.615
R111 VTAIL.n106 VTAIL.n105 104.615
R112 VTAIL.n90 VTAIL.n89 104.615
R113 VTAIL.n89 VTAIL.n75 104.615
R114 VTAIL.n82 VTAIL.n75 104.615
R115 VTAIL.n82 VTAIL.n81 104.615
R116 VTAIL.n177 VTAIL.t2 52.3082
R117 VTAIL.n9 VTAIL.t3 52.3082
R118 VTAIL.n33 VTAIL.t7 52.3082
R119 VTAIL.n57 VTAIL.t4 52.3082
R120 VTAIL.n153 VTAIL.t6 52.3082
R121 VTAIL.n129 VTAIL.t5 52.3082
R122 VTAIL.n105 VTAIL.t1 52.3082
R123 VTAIL.n81 VTAIL.t0 52.3082
R124 VTAIL.n191 VTAIL.n190 32.1853
R125 VTAIL.n23 VTAIL.n22 32.1853
R126 VTAIL.n47 VTAIL.n46 32.1853
R127 VTAIL.n71 VTAIL.n70 32.1853
R128 VTAIL.n167 VTAIL.n166 32.1853
R129 VTAIL.n143 VTAIL.n142 32.1853
R130 VTAIL.n119 VTAIL.n118 32.1853
R131 VTAIL.n95 VTAIL.n94 32.1853
R132 VTAIL.n191 VTAIL.n167 18.7721
R133 VTAIL.n95 VTAIL.n71 18.7721
R134 VTAIL.n176 VTAIL.n175 15.6631
R135 VTAIL.n8 VTAIL.n7 15.6631
R136 VTAIL.n32 VTAIL.n31 15.6631
R137 VTAIL.n56 VTAIL.n55 15.6631
R138 VTAIL.n152 VTAIL.n151 15.6631
R139 VTAIL.n128 VTAIL.n127 15.6631
R140 VTAIL.n104 VTAIL.n103 15.6631
R141 VTAIL.n80 VTAIL.n79 15.6631
R142 VTAIL.n179 VTAIL.n174 12.8005
R143 VTAIL.n11 VTAIL.n6 12.8005
R144 VTAIL.n35 VTAIL.n30 12.8005
R145 VTAIL.n59 VTAIL.n54 12.8005
R146 VTAIL.n155 VTAIL.n150 12.8005
R147 VTAIL.n131 VTAIL.n126 12.8005
R148 VTAIL.n107 VTAIL.n102 12.8005
R149 VTAIL.n83 VTAIL.n78 12.8005
R150 VTAIL.n180 VTAIL.n172 12.0247
R151 VTAIL.n12 VTAIL.n4 12.0247
R152 VTAIL.n36 VTAIL.n28 12.0247
R153 VTAIL.n60 VTAIL.n52 12.0247
R154 VTAIL.n156 VTAIL.n148 12.0247
R155 VTAIL.n132 VTAIL.n124 12.0247
R156 VTAIL.n108 VTAIL.n100 12.0247
R157 VTAIL.n84 VTAIL.n76 12.0247
R158 VTAIL.n184 VTAIL.n183 11.249
R159 VTAIL.n16 VTAIL.n15 11.249
R160 VTAIL.n40 VTAIL.n39 11.249
R161 VTAIL.n64 VTAIL.n63 11.249
R162 VTAIL.n160 VTAIL.n159 11.249
R163 VTAIL.n136 VTAIL.n135 11.249
R164 VTAIL.n112 VTAIL.n111 11.249
R165 VTAIL.n88 VTAIL.n87 11.249
R166 VTAIL.n187 VTAIL.n170 10.4732
R167 VTAIL.n19 VTAIL.n2 10.4732
R168 VTAIL.n43 VTAIL.n26 10.4732
R169 VTAIL.n67 VTAIL.n50 10.4732
R170 VTAIL.n163 VTAIL.n146 10.4732
R171 VTAIL.n139 VTAIL.n122 10.4732
R172 VTAIL.n115 VTAIL.n98 10.4732
R173 VTAIL.n91 VTAIL.n74 10.4732
R174 VTAIL.n188 VTAIL.n168 9.69747
R175 VTAIL.n20 VTAIL.n0 9.69747
R176 VTAIL.n44 VTAIL.n24 9.69747
R177 VTAIL.n68 VTAIL.n48 9.69747
R178 VTAIL.n164 VTAIL.n144 9.69747
R179 VTAIL.n140 VTAIL.n120 9.69747
R180 VTAIL.n116 VTAIL.n96 9.69747
R181 VTAIL.n92 VTAIL.n72 9.69747
R182 VTAIL.n190 VTAIL.n189 9.45567
R183 VTAIL.n22 VTAIL.n21 9.45567
R184 VTAIL.n46 VTAIL.n45 9.45567
R185 VTAIL.n70 VTAIL.n69 9.45567
R186 VTAIL.n166 VTAIL.n165 9.45567
R187 VTAIL.n142 VTAIL.n141 9.45567
R188 VTAIL.n118 VTAIL.n117 9.45567
R189 VTAIL.n94 VTAIL.n93 9.45567
R190 VTAIL.n189 VTAIL.n188 9.3005
R191 VTAIL.n170 VTAIL.n169 9.3005
R192 VTAIL.n183 VTAIL.n182 9.3005
R193 VTAIL.n181 VTAIL.n180 9.3005
R194 VTAIL.n174 VTAIL.n173 9.3005
R195 VTAIL.n21 VTAIL.n20 9.3005
R196 VTAIL.n2 VTAIL.n1 9.3005
R197 VTAIL.n15 VTAIL.n14 9.3005
R198 VTAIL.n13 VTAIL.n12 9.3005
R199 VTAIL.n6 VTAIL.n5 9.3005
R200 VTAIL.n45 VTAIL.n44 9.3005
R201 VTAIL.n26 VTAIL.n25 9.3005
R202 VTAIL.n39 VTAIL.n38 9.3005
R203 VTAIL.n37 VTAIL.n36 9.3005
R204 VTAIL.n30 VTAIL.n29 9.3005
R205 VTAIL.n69 VTAIL.n68 9.3005
R206 VTAIL.n50 VTAIL.n49 9.3005
R207 VTAIL.n63 VTAIL.n62 9.3005
R208 VTAIL.n61 VTAIL.n60 9.3005
R209 VTAIL.n54 VTAIL.n53 9.3005
R210 VTAIL.n165 VTAIL.n164 9.3005
R211 VTAIL.n146 VTAIL.n145 9.3005
R212 VTAIL.n159 VTAIL.n158 9.3005
R213 VTAIL.n157 VTAIL.n156 9.3005
R214 VTAIL.n150 VTAIL.n149 9.3005
R215 VTAIL.n141 VTAIL.n140 9.3005
R216 VTAIL.n122 VTAIL.n121 9.3005
R217 VTAIL.n135 VTAIL.n134 9.3005
R218 VTAIL.n133 VTAIL.n132 9.3005
R219 VTAIL.n126 VTAIL.n125 9.3005
R220 VTAIL.n117 VTAIL.n116 9.3005
R221 VTAIL.n98 VTAIL.n97 9.3005
R222 VTAIL.n111 VTAIL.n110 9.3005
R223 VTAIL.n109 VTAIL.n108 9.3005
R224 VTAIL.n102 VTAIL.n101 9.3005
R225 VTAIL.n93 VTAIL.n92 9.3005
R226 VTAIL.n74 VTAIL.n73 9.3005
R227 VTAIL.n87 VTAIL.n86 9.3005
R228 VTAIL.n85 VTAIL.n84 9.3005
R229 VTAIL.n78 VTAIL.n77 9.3005
R230 VTAIL.n175 VTAIL.n173 4.39059
R231 VTAIL.n7 VTAIL.n5 4.39059
R232 VTAIL.n31 VTAIL.n29 4.39059
R233 VTAIL.n55 VTAIL.n53 4.39059
R234 VTAIL.n151 VTAIL.n149 4.39059
R235 VTAIL.n127 VTAIL.n125 4.39059
R236 VTAIL.n103 VTAIL.n101 4.39059
R237 VTAIL.n79 VTAIL.n77 4.39059
R238 VTAIL.n190 VTAIL.n168 4.26717
R239 VTAIL.n22 VTAIL.n0 4.26717
R240 VTAIL.n46 VTAIL.n24 4.26717
R241 VTAIL.n70 VTAIL.n48 4.26717
R242 VTAIL.n166 VTAIL.n144 4.26717
R243 VTAIL.n142 VTAIL.n120 4.26717
R244 VTAIL.n118 VTAIL.n96 4.26717
R245 VTAIL.n94 VTAIL.n72 4.26717
R246 VTAIL.n188 VTAIL.n187 3.49141
R247 VTAIL.n20 VTAIL.n19 3.49141
R248 VTAIL.n44 VTAIL.n43 3.49141
R249 VTAIL.n68 VTAIL.n67 3.49141
R250 VTAIL.n164 VTAIL.n163 3.49141
R251 VTAIL.n140 VTAIL.n139 3.49141
R252 VTAIL.n116 VTAIL.n115 3.49141
R253 VTAIL.n92 VTAIL.n91 3.49141
R254 VTAIL.n184 VTAIL.n170 2.71565
R255 VTAIL.n16 VTAIL.n2 2.71565
R256 VTAIL.n40 VTAIL.n26 2.71565
R257 VTAIL.n64 VTAIL.n50 2.71565
R258 VTAIL.n160 VTAIL.n146 2.71565
R259 VTAIL.n136 VTAIL.n122 2.71565
R260 VTAIL.n112 VTAIL.n98 2.71565
R261 VTAIL.n88 VTAIL.n74 2.71565
R262 VTAIL.n119 VTAIL.n95 2.47464
R263 VTAIL.n167 VTAIL.n143 2.47464
R264 VTAIL.n71 VTAIL.n47 2.47464
R265 VTAIL.n183 VTAIL.n172 1.93989
R266 VTAIL.n15 VTAIL.n4 1.93989
R267 VTAIL.n39 VTAIL.n28 1.93989
R268 VTAIL.n63 VTAIL.n52 1.93989
R269 VTAIL.n159 VTAIL.n148 1.93989
R270 VTAIL.n135 VTAIL.n124 1.93989
R271 VTAIL.n111 VTAIL.n100 1.93989
R272 VTAIL.n87 VTAIL.n76 1.93989
R273 VTAIL VTAIL.n23 1.29576
R274 VTAIL VTAIL.n191 1.17938
R275 VTAIL.n180 VTAIL.n179 1.16414
R276 VTAIL.n12 VTAIL.n11 1.16414
R277 VTAIL.n36 VTAIL.n35 1.16414
R278 VTAIL.n60 VTAIL.n59 1.16414
R279 VTAIL.n156 VTAIL.n155 1.16414
R280 VTAIL.n132 VTAIL.n131 1.16414
R281 VTAIL.n108 VTAIL.n107 1.16414
R282 VTAIL.n84 VTAIL.n83 1.16414
R283 VTAIL.n143 VTAIL.n119 0.470328
R284 VTAIL.n47 VTAIL.n23 0.470328
R285 VTAIL.n176 VTAIL.n174 0.388379
R286 VTAIL.n8 VTAIL.n6 0.388379
R287 VTAIL.n32 VTAIL.n30 0.388379
R288 VTAIL.n56 VTAIL.n54 0.388379
R289 VTAIL.n152 VTAIL.n150 0.388379
R290 VTAIL.n128 VTAIL.n126 0.388379
R291 VTAIL.n104 VTAIL.n102 0.388379
R292 VTAIL.n80 VTAIL.n78 0.388379
R293 VTAIL.n181 VTAIL.n173 0.155672
R294 VTAIL.n182 VTAIL.n181 0.155672
R295 VTAIL.n182 VTAIL.n169 0.155672
R296 VTAIL.n189 VTAIL.n169 0.155672
R297 VTAIL.n13 VTAIL.n5 0.155672
R298 VTAIL.n14 VTAIL.n13 0.155672
R299 VTAIL.n14 VTAIL.n1 0.155672
R300 VTAIL.n21 VTAIL.n1 0.155672
R301 VTAIL.n37 VTAIL.n29 0.155672
R302 VTAIL.n38 VTAIL.n37 0.155672
R303 VTAIL.n38 VTAIL.n25 0.155672
R304 VTAIL.n45 VTAIL.n25 0.155672
R305 VTAIL.n61 VTAIL.n53 0.155672
R306 VTAIL.n62 VTAIL.n61 0.155672
R307 VTAIL.n62 VTAIL.n49 0.155672
R308 VTAIL.n69 VTAIL.n49 0.155672
R309 VTAIL.n165 VTAIL.n145 0.155672
R310 VTAIL.n158 VTAIL.n145 0.155672
R311 VTAIL.n158 VTAIL.n157 0.155672
R312 VTAIL.n157 VTAIL.n149 0.155672
R313 VTAIL.n141 VTAIL.n121 0.155672
R314 VTAIL.n134 VTAIL.n121 0.155672
R315 VTAIL.n134 VTAIL.n133 0.155672
R316 VTAIL.n133 VTAIL.n125 0.155672
R317 VTAIL.n117 VTAIL.n97 0.155672
R318 VTAIL.n110 VTAIL.n97 0.155672
R319 VTAIL.n110 VTAIL.n109 0.155672
R320 VTAIL.n109 VTAIL.n101 0.155672
R321 VTAIL.n93 VTAIL.n73 0.155672
R322 VTAIL.n86 VTAIL.n73 0.155672
R323 VTAIL.n86 VTAIL.n85 0.155672
R324 VTAIL.n85 VTAIL.n77 0.155672
R325 VDD1 VDD1.n1 106.234
R326 VDD1 VDD1.n0 70.6998
R327 VDD1.n0 VDD1.t2 4.34261
R328 VDD1.n0 VDD1.t3 4.34261
R329 VDD1.n1 VDD1.t0 4.34261
R330 VDD1.n1 VDD1.t1 4.34261
R331 B.n526 B.n525 585
R332 B.n527 B.n526 585
R333 B.n189 B.n88 585
R334 B.n188 B.n187 585
R335 B.n186 B.n185 585
R336 B.n184 B.n183 585
R337 B.n182 B.n181 585
R338 B.n180 B.n179 585
R339 B.n178 B.n177 585
R340 B.n176 B.n175 585
R341 B.n174 B.n173 585
R342 B.n172 B.n171 585
R343 B.n170 B.n169 585
R344 B.n168 B.n167 585
R345 B.n166 B.n165 585
R346 B.n164 B.n163 585
R347 B.n162 B.n161 585
R348 B.n160 B.n159 585
R349 B.n158 B.n157 585
R350 B.n156 B.n155 585
R351 B.n154 B.n153 585
R352 B.n151 B.n150 585
R353 B.n149 B.n148 585
R354 B.n147 B.n146 585
R355 B.n145 B.n144 585
R356 B.n143 B.n142 585
R357 B.n141 B.n140 585
R358 B.n139 B.n138 585
R359 B.n137 B.n136 585
R360 B.n135 B.n134 585
R361 B.n133 B.n132 585
R362 B.n131 B.n130 585
R363 B.n129 B.n128 585
R364 B.n127 B.n126 585
R365 B.n125 B.n124 585
R366 B.n123 B.n122 585
R367 B.n121 B.n120 585
R368 B.n119 B.n118 585
R369 B.n117 B.n116 585
R370 B.n115 B.n114 585
R371 B.n113 B.n112 585
R372 B.n111 B.n110 585
R373 B.n109 B.n108 585
R374 B.n107 B.n106 585
R375 B.n105 B.n104 585
R376 B.n103 B.n102 585
R377 B.n101 B.n100 585
R378 B.n99 B.n98 585
R379 B.n97 B.n96 585
R380 B.n95 B.n94 585
R381 B.n524 B.n63 585
R382 B.n528 B.n63 585
R383 B.n523 B.n62 585
R384 B.n529 B.n62 585
R385 B.n522 B.n521 585
R386 B.n521 B.n58 585
R387 B.n520 B.n57 585
R388 B.n535 B.n57 585
R389 B.n519 B.n56 585
R390 B.n536 B.n56 585
R391 B.n518 B.n55 585
R392 B.n537 B.n55 585
R393 B.n517 B.n516 585
R394 B.n516 B.n51 585
R395 B.n515 B.n50 585
R396 B.n543 B.n50 585
R397 B.n514 B.n49 585
R398 B.n544 B.n49 585
R399 B.n513 B.n48 585
R400 B.n545 B.n48 585
R401 B.n512 B.n511 585
R402 B.n511 B.n44 585
R403 B.n510 B.n43 585
R404 B.n551 B.n43 585
R405 B.n509 B.n42 585
R406 B.n552 B.n42 585
R407 B.n508 B.n41 585
R408 B.n553 B.n41 585
R409 B.n507 B.n506 585
R410 B.n506 B.n37 585
R411 B.n505 B.n36 585
R412 B.n559 B.n36 585
R413 B.n504 B.n35 585
R414 B.n560 B.n35 585
R415 B.n503 B.n34 585
R416 B.n561 B.n34 585
R417 B.n502 B.n501 585
R418 B.n501 B.n30 585
R419 B.n500 B.n29 585
R420 B.n567 B.n29 585
R421 B.n499 B.n28 585
R422 B.n568 B.n28 585
R423 B.n498 B.n27 585
R424 B.n569 B.n27 585
R425 B.n497 B.n496 585
R426 B.n496 B.n23 585
R427 B.n495 B.n22 585
R428 B.n575 B.n22 585
R429 B.n494 B.n21 585
R430 B.n576 B.n21 585
R431 B.n493 B.n20 585
R432 B.n577 B.n20 585
R433 B.n492 B.n491 585
R434 B.n491 B.n16 585
R435 B.n490 B.n15 585
R436 B.n583 B.n15 585
R437 B.n489 B.n14 585
R438 B.n584 B.n14 585
R439 B.n488 B.n13 585
R440 B.n585 B.n13 585
R441 B.n487 B.n486 585
R442 B.n486 B.n12 585
R443 B.n485 B.n484 585
R444 B.n485 B.n8 585
R445 B.n483 B.n7 585
R446 B.n592 B.n7 585
R447 B.n482 B.n6 585
R448 B.n593 B.n6 585
R449 B.n481 B.n5 585
R450 B.n594 B.n5 585
R451 B.n480 B.n479 585
R452 B.n479 B.n4 585
R453 B.n478 B.n190 585
R454 B.n478 B.n477 585
R455 B.n468 B.n191 585
R456 B.n192 B.n191 585
R457 B.n470 B.n469 585
R458 B.n471 B.n470 585
R459 B.n467 B.n197 585
R460 B.n197 B.n196 585
R461 B.n466 B.n465 585
R462 B.n465 B.n464 585
R463 B.n199 B.n198 585
R464 B.n200 B.n199 585
R465 B.n457 B.n456 585
R466 B.n458 B.n457 585
R467 B.n455 B.n205 585
R468 B.n205 B.n204 585
R469 B.n454 B.n453 585
R470 B.n453 B.n452 585
R471 B.n207 B.n206 585
R472 B.n208 B.n207 585
R473 B.n445 B.n444 585
R474 B.n446 B.n445 585
R475 B.n443 B.n213 585
R476 B.n213 B.n212 585
R477 B.n442 B.n441 585
R478 B.n441 B.n440 585
R479 B.n215 B.n214 585
R480 B.n216 B.n215 585
R481 B.n433 B.n432 585
R482 B.n434 B.n433 585
R483 B.n431 B.n221 585
R484 B.n221 B.n220 585
R485 B.n430 B.n429 585
R486 B.n429 B.n428 585
R487 B.n223 B.n222 585
R488 B.n224 B.n223 585
R489 B.n421 B.n420 585
R490 B.n422 B.n421 585
R491 B.n419 B.n229 585
R492 B.n229 B.n228 585
R493 B.n418 B.n417 585
R494 B.n417 B.n416 585
R495 B.n231 B.n230 585
R496 B.n232 B.n231 585
R497 B.n409 B.n408 585
R498 B.n410 B.n409 585
R499 B.n407 B.n237 585
R500 B.n237 B.n236 585
R501 B.n406 B.n405 585
R502 B.n405 B.n404 585
R503 B.n239 B.n238 585
R504 B.n240 B.n239 585
R505 B.n397 B.n396 585
R506 B.n398 B.n397 585
R507 B.n395 B.n245 585
R508 B.n245 B.n244 585
R509 B.n394 B.n393 585
R510 B.n393 B.n392 585
R511 B.n247 B.n246 585
R512 B.n248 B.n247 585
R513 B.n385 B.n384 585
R514 B.n386 B.n385 585
R515 B.n383 B.n253 585
R516 B.n253 B.n252 585
R517 B.n377 B.n376 585
R518 B.n375 B.n279 585
R519 B.n374 B.n278 585
R520 B.n379 B.n278 585
R521 B.n373 B.n372 585
R522 B.n371 B.n370 585
R523 B.n369 B.n368 585
R524 B.n367 B.n366 585
R525 B.n365 B.n364 585
R526 B.n363 B.n362 585
R527 B.n361 B.n360 585
R528 B.n359 B.n358 585
R529 B.n357 B.n356 585
R530 B.n355 B.n354 585
R531 B.n353 B.n352 585
R532 B.n351 B.n350 585
R533 B.n349 B.n348 585
R534 B.n347 B.n346 585
R535 B.n345 B.n344 585
R536 B.n343 B.n342 585
R537 B.n341 B.n340 585
R538 B.n338 B.n337 585
R539 B.n336 B.n335 585
R540 B.n334 B.n333 585
R541 B.n332 B.n331 585
R542 B.n330 B.n329 585
R543 B.n328 B.n327 585
R544 B.n326 B.n325 585
R545 B.n324 B.n323 585
R546 B.n322 B.n321 585
R547 B.n320 B.n319 585
R548 B.n318 B.n317 585
R549 B.n316 B.n315 585
R550 B.n314 B.n313 585
R551 B.n312 B.n311 585
R552 B.n310 B.n309 585
R553 B.n308 B.n307 585
R554 B.n306 B.n305 585
R555 B.n304 B.n303 585
R556 B.n302 B.n301 585
R557 B.n300 B.n299 585
R558 B.n298 B.n297 585
R559 B.n296 B.n295 585
R560 B.n294 B.n293 585
R561 B.n292 B.n291 585
R562 B.n290 B.n289 585
R563 B.n288 B.n287 585
R564 B.n286 B.n285 585
R565 B.n255 B.n254 585
R566 B.n382 B.n381 585
R567 B.n251 B.n250 585
R568 B.n252 B.n251 585
R569 B.n388 B.n387 585
R570 B.n387 B.n386 585
R571 B.n389 B.n249 585
R572 B.n249 B.n248 585
R573 B.n391 B.n390 585
R574 B.n392 B.n391 585
R575 B.n243 B.n242 585
R576 B.n244 B.n243 585
R577 B.n400 B.n399 585
R578 B.n399 B.n398 585
R579 B.n401 B.n241 585
R580 B.n241 B.n240 585
R581 B.n403 B.n402 585
R582 B.n404 B.n403 585
R583 B.n235 B.n234 585
R584 B.n236 B.n235 585
R585 B.n412 B.n411 585
R586 B.n411 B.n410 585
R587 B.n413 B.n233 585
R588 B.n233 B.n232 585
R589 B.n415 B.n414 585
R590 B.n416 B.n415 585
R591 B.n227 B.n226 585
R592 B.n228 B.n227 585
R593 B.n424 B.n423 585
R594 B.n423 B.n422 585
R595 B.n425 B.n225 585
R596 B.n225 B.n224 585
R597 B.n427 B.n426 585
R598 B.n428 B.n427 585
R599 B.n219 B.n218 585
R600 B.n220 B.n219 585
R601 B.n436 B.n435 585
R602 B.n435 B.n434 585
R603 B.n437 B.n217 585
R604 B.n217 B.n216 585
R605 B.n439 B.n438 585
R606 B.n440 B.n439 585
R607 B.n211 B.n210 585
R608 B.n212 B.n211 585
R609 B.n448 B.n447 585
R610 B.n447 B.n446 585
R611 B.n449 B.n209 585
R612 B.n209 B.n208 585
R613 B.n451 B.n450 585
R614 B.n452 B.n451 585
R615 B.n203 B.n202 585
R616 B.n204 B.n203 585
R617 B.n460 B.n459 585
R618 B.n459 B.n458 585
R619 B.n461 B.n201 585
R620 B.n201 B.n200 585
R621 B.n463 B.n462 585
R622 B.n464 B.n463 585
R623 B.n195 B.n194 585
R624 B.n196 B.n195 585
R625 B.n473 B.n472 585
R626 B.n472 B.n471 585
R627 B.n474 B.n193 585
R628 B.n193 B.n192 585
R629 B.n476 B.n475 585
R630 B.n477 B.n476 585
R631 B.n3 B.n0 585
R632 B.n4 B.n3 585
R633 B.n591 B.n1 585
R634 B.n592 B.n591 585
R635 B.n590 B.n589 585
R636 B.n590 B.n8 585
R637 B.n588 B.n9 585
R638 B.n12 B.n9 585
R639 B.n587 B.n586 585
R640 B.n586 B.n585 585
R641 B.n11 B.n10 585
R642 B.n584 B.n11 585
R643 B.n582 B.n581 585
R644 B.n583 B.n582 585
R645 B.n580 B.n17 585
R646 B.n17 B.n16 585
R647 B.n579 B.n578 585
R648 B.n578 B.n577 585
R649 B.n19 B.n18 585
R650 B.n576 B.n19 585
R651 B.n574 B.n573 585
R652 B.n575 B.n574 585
R653 B.n572 B.n24 585
R654 B.n24 B.n23 585
R655 B.n571 B.n570 585
R656 B.n570 B.n569 585
R657 B.n26 B.n25 585
R658 B.n568 B.n26 585
R659 B.n566 B.n565 585
R660 B.n567 B.n566 585
R661 B.n564 B.n31 585
R662 B.n31 B.n30 585
R663 B.n563 B.n562 585
R664 B.n562 B.n561 585
R665 B.n33 B.n32 585
R666 B.n560 B.n33 585
R667 B.n558 B.n557 585
R668 B.n559 B.n558 585
R669 B.n556 B.n38 585
R670 B.n38 B.n37 585
R671 B.n555 B.n554 585
R672 B.n554 B.n553 585
R673 B.n40 B.n39 585
R674 B.n552 B.n40 585
R675 B.n550 B.n549 585
R676 B.n551 B.n550 585
R677 B.n548 B.n45 585
R678 B.n45 B.n44 585
R679 B.n547 B.n546 585
R680 B.n546 B.n545 585
R681 B.n47 B.n46 585
R682 B.n544 B.n47 585
R683 B.n542 B.n541 585
R684 B.n543 B.n542 585
R685 B.n540 B.n52 585
R686 B.n52 B.n51 585
R687 B.n539 B.n538 585
R688 B.n538 B.n537 585
R689 B.n54 B.n53 585
R690 B.n536 B.n54 585
R691 B.n534 B.n533 585
R692 B.n535 B.n534 585
R693 B.n532 B.n59 585
R694 B.n59 B.n58 585
R695 B.n531 B.n530 585
R696 B.n530 B.n529 585
R697 B.n61 B.n60 585
R698 B.n528 B.n61 585
R699 B.n595 B.n594 585
R700 B.n593 B.n2 585
R701 B.n94 B.n61 492.5
R702 B.n526 B.n63 492.5
R703 B.n381 B.n253 492.5
R704 B.n377 B.n251 492.5
R705 B.n527 B.n87 256.663
R706 B.n527 B.n86 256.663
R707 B.n527 B.n85 256.663
R708 B.n527 B.n84 256.663
R709 B.n527 B.n83 256.663
R710 B.n527 B.n82 256.663
R711 B.n527 B.n81 256.663
R712 B.n527 B.n80 256.663
R713 B.n527 B.n79 256.663
R714 B.n527 B.n78 256.663
R715 B.n527 B.n77 256.663
R716 B.n527 B.n76 256.663
R717 B.n527 B.n75 256.663
R718 B.n527 B.n74 256.663
R719 B.n527 B.n73 256.663
R720 B.n527 B.n72 256.663
R721 B.n527 B.n71 256.663
R722 B.n527 B.n70 256.663
R723 B.n527 B.n69 256.663
R724 B.n527 B.n68 256.663
R725 B.n527 B.n67 256.663
R726 B.n527 B.n66 256.663
R727 B.n527 B.n65 256.663
R728 B.n527 B.n64 256.663
R729 B.n379 B.n378 256.663
R730 B.n379 B.n256 256.663
R731 B.n379 B.n257 256.663
R732 B.n379 B.n258 256.663
R733 B.n379 B.n259 256.663
R734 B.n379 B.n260 256.663
R735 B.n379 B.n261 256.663
R736 B.n379 B.n262 256.663
R737 B.n379 B.n263 256.663
R738 B.n379 B.n264 256.663
R739 B.n379 B.n265 256.663
R740 B.n379 B.n266 256.663
R741 B.n379 B.n267 256.663
R742 B.n379 B.n268 256.663
R743 B.n379 B.n269 256.663
R744 B.n379 B.n270 256.663
R745 B.n379 B.n271 256.663
R746 B.n379 B.n272 256.663
R747 B.n379 B.n273 256.663
R748 B.n379 B.n274 256.663
R749 B.n379 B.n275 256.663
R750 B.n379 B.n276 256.663
R751 B.n379 B.n277 256.663
R752 B.n380 B.n379 256.663
R753 B.n597 B.n596 256.663
R754 B.n91 B.t4 251.22
R755 B.n89 B.t12 251.22
R756 B.n282 B.t15 251.22
R757 B.n280 B.t8 251.22
R758 B.n89 B.t13 209.916
R759 B.n282 B.t17 209.916
R760 B.n91 B.t6 209.916
R761 B.n280 B.t11 209.916
R762 B.n98 B.n97 163.367
R763 B.n102 B.n101 163.367
R764 B.n106 B.n105 163.367
R765 B.n110 B.n109 163.367
R766 B.n114 B.n113 163.367
R767 B.n118 B.n117 163.367
R768 B.n122 B.n121 163.367
R769 B.n126 B.n125 163.367
R770 B.n130 B.n129 163.367
R771 B.n134 B.n133 163.367
R772 B.n138 B.n137 163.367
R773 B.n142 B.n141 163.367
R774 B.n146 B.n145 163.367
R775 B.n150 B.n149 163.367
R776 B.n155 B.n154 163.367
R777 B.n159 B.n158 163.367
R778 B.n163 B.n162 163.367
R779 B.n167 B.n166 163.367
R780 B.n171 B.n170 163.367
R781 B.n175 B.n174 163.367
R782 B.n179 B.n178 163.367
R783 B.n183 B.n182 163.367
R784 B.n187 B.n186 163.367
R785 B.n526 B.n88 163.367
R786 B.n385 B.n253 163.367
R787 B.n385 B.n247 163.367
R788 B.n393 B.n247 163.367
R789 B.n393 B.n245 163.367
R790 B.n397 B.n245 163.367
R791 B.n397 B.n239 163.367
R792 B.n405 B.n239 163.367
R793 B.n405 B.n237 163.367
R794 B.n409 B.n237 163.367
R795 B.n409 B.n231 163.367
R796 B.n417 B.n231 163.367
R797 B.n417 B.n229 163.367
R798 B.n421 B.n229 163.367
R799 B.n421 B.n223 163.367
R800 B.n429 B.n223 163.367
R801 B.n429 B.n221 163.367
R802 B.n433 B.n221 163.367
R803 B.n433 B.n215 163.367
R804 B.n441 B.n215 163.367
R805 B.n441 B.n213 163.367
R806 B.n445 B.n213 163.367
R807 B.n445 B.n207 163.367
R808 B.n453 B.n207 163.367
R809 B.n453 B.n205 163.367
R810 B.n457 B.n205 163.367
R811 B.n457 B.n199 163.367
R812 B.n465 B.n199 163.367
R813 B.n465 B.n197 163.367
R814 B.n470 B.n197 163.367
R815 B.n470 B.n191 163.367
R816 B.n478 B.n191 163.367
R817 B.n479 B.n478 163.367
R818 B.n479 B.n5 163.367
R819 B.n6 B.n5 163.367
R820 B.n7 B.n6 163.367
R821 B.n485 B.n7 163.367
R822 B.n486 B.n485 163.367
R823 B.n486 B.n13 163.367
R824 B.n14 B.n13 163.367
R825 B.n15 B.n14 163.367
R826 B.n491 B.n15 163.367
R827 B.n491 B.n20 163.367
R828 B.n21 B.n20 163.367
R829 B.n22 B.n21 163.367
R830 B.n496 B.n22 163.367
R831 B.n496 B.n27 163.367
R832 B.n28 B.n27 163.367
R833 B.n29 B.n28 163.367
R834 B.n501 B.n29 163.367
R835 B.n501 B.n34 163.367
R836 B.n35 B.n34 163.367
R837 B.n36 B.n35 163.367
R838 B.n506 B.n36 163.367
R839 B.n506 B.n41 163.367
R840 B.n42 B.n41 163.367
R841 B.n43 B.n42 163.367
R842 B.n511 B.n43 163.367
R843 B.n511 B.n48 163.367
R844 B.n49 B.n48 163.367
R845 B.n50 B.n49 163.367
R846 B.n516 B.n50 163.367
R847 B.n516 B.n55 163.367
R848 B.n56 B.n55 163.367
R849 B.n57 B.n56 163.367
R850 B.n521 B.n57 163.367
R851 B.n521 B.n62 163.367
R852 B.n63 B.n62 163.367
R853 B.n279 B.n278 163.367
R854 B.n372 B.n278 163.367
R855 B.n370 B.n369 163.367
R856 B.n366 B.n365 163.367
R857 B.n362 B.n361 163.367
R858 B.n358 B.n357 163.367
R859 B.n354 B.n353 163.367
R860 B.n350 B.n349 163.367
R861 B.n346 B.n345 163.367
R862 B.n342 B.n341 163.367
R863 B.n337 B.n336 163.367
R864 B.n333 B.n332 163.367
R865 B.n329 B.n328 163.367
R866 B.n325 B.n324 163.367
R867 B.n321 B.n320 163.367
R868 B.n317 B.n316 163.367
R869 B.n313 B.n312 163.367
R870 B.n309 B.n308 163.367
R871 B.n305 B.n304 163.367
R872 B.n301 B.n300 163.367
R873 B.n297 B.n296 163.367
R874 B.n293 B.n292 163.367
R875 B.n289 B.n288 163.367
R876 B.n285 B.n255 163.367
R877 B.n387 B.n251 163.367
R878 B.n387 B.n249 163.367
R879 B.n391 B.n249 163.367
R880 B.n391 B.n243 163.367
R881 B.n399 B.n243 163.367
R882 B.n399 B.n241 163.367
R883 B.n403 B.n241 163.367
R884 B.n403 B.n235 163.367
R885 B.n411 B.n235 163.367
R886 B.n411 B.n233 163.367
R887 B.n415 B.n233 163.367
R888 B.n415 B.n227 163.367
R889 B.n423 B.n227 163.367
R890 B.n423 B.n225 163.367
R891 B.n427 B.n225 163.367
R892 B.n427 B.n219 163.367
R893 B.n435 B.n219 163.367
R894 B.n435 B.n217 163.367
R895 B.n439 B.n217 163.367
R896 B.n439 B.n211 163.367
R897 B.n447 B.n211 163.367
R898 B.n447 B.n209 163.367
R899 B.n451 B.n209 163.367
R900 B.n451 B.n203 163.367
R901 B.n459 B.n203 163.367
R902 B.n459 B.n201 163.367
R903 B.n463 B.n201 163.367
R904 B.n463 B.n195 163.367
R905 B.n472 B.n195 163.367
R906 B.n472 B.n193 163.367
R907 B.n476 B.n193 163.367
R908 B.n476 B.n3 163.367
R909 B.n595 B.n3 163.367
R910 B.n591 B.n2 163.367
R911 B.n591 B.n590 163.367
R912 B.n590 B.n9 163.367
R913 B.n586 B.n9 163.367
R914 B.n586 B.n11 163.367
R915 B.n582 B.n11 163.367
R916 B.n582 B.n17 163.367
R917 B.n578 B.n17 163.367
R918 B.n578 B.n19 163.367
R919 B.n574 B.n19 163.367
R920 B.n574 B.n24 163.367
R921 B.n570 B.n24 163.367
R922 B.n570 B.n26 163.367
R923 B.n566 B.n26 163.367
R924 B.n566 B.n31 163.367
R925 B.n562 B.n31 163.367
R926 B.n562 B.n33 163.367
R927 B.n558 B.n33 163.367
R928 B.n558 B.n38 163.367
R929 B.n554 B.n38 163.367
R930 B.n554 B.n40 163.367
R931 B.n550 B.n40 163.367
R932 B.n550 B.n45 163.367
R933 B.n546 B.n45 163.367
R934 B.n546 B.n47 163.367
R935 B.n542 B.n47 163.367
R936 B.n542 B.n52 163.367
R937 B.n538 B.n52 163.367
R938 B.n538 B.n54 163.367
R939 B.n534 B.n54 163.367
R940 B.n534 B.n59 163.367
R941 B.n530 B.n59 163.367
R942 B.n530 B.n61 163.367
R943 B.n90 B.t14 154.255
R944 B.n283 B.t16 154.255
R945 B.n92 B.t7 154.255
R946 B.n281 B.t10 154.255
R947 B.n379 B.n252 133.096
R948 B.n528 B.n527 133.096
R949 B.n386 B.n252 76.0554
R950 B.n386 B.n248 76.0554
R951 B.n392 B.n248 76.0554
R952 B.n392 B.n244 76.0554
R953 B.n398 B.n244 76.0554
R954 B.n398 B.n240 76.0554
R955 B.n404 B.n240 76.0554
R956 B.n410 B.n236 76.0554
R957 B.n410 B.n232 76.0554
R958 B.n416 B.n232 76.0554
R959 B.n416 B.n228 76.0554
R960 B.n422 B.n228 76.0554
R961 B.n422 B.n224 76.0554
R962 B.n428 B.n224 76.0554
R963 B.n428 B.n220 76.0554
R964 B.n434 B.n220 76.0554
R965 B.n434 B.n216 76.0554
R966 B.n440 B.n216 76.0554
R967 B.n446 B.n212 76.0554
R968 B.n446 B.n208 76.0554
R969 B.n452 B.n208 76.0554
R970 B.n452 B.n204 76.0554
R971 B.n458 B.n204 76.0554
R972 B.n458 B.n200 76.0554
R973 B.n464 B.n200 76.0554
R974 B.n471 B.n196 76.0554
R975 B.n471 B.n192 76.0554
R976 B.n477 B.n192 76.0554
R977 B.n477 B.n4 76.0554
R978 B.n594 B.n4 76.0554
R979 B.n594 B.n593 76.0554
R980 B.n593 B.n592 76.0554
R981 B.n592 B.n8 76.0554
R982 B.n12 B.n8 76.0554
R983 B.n585 B.n12 76.0554
R984 B.n585 B.n584 76.0554
R985 B.n583 B.n16 76.0554
R986 B.n577 B.n16 76.0554
R987 B.n577 B.n576 76.0554
R988 B.n576 B.n575 76.0554
R989 B.n575 B.n23 76.0554
R990 B.n569 B.n23 76.0554
R991 B.n569 B.n568 76.0554
R992 B.n567 B.n30 76.0554
R993 B.n561 B.n30 76.0554
R994 B.n561 B.n560 76.0554
R995 B.n560 B.n559 76.0554
R996 B.n559 B.n37 76.0554
R997 B.n553 B.n37 76.0554
R998 B.n553 B.n552 76.0554
R999 B.n552 B.n551 76.0554
R1000 B.n551 B.n44 76.0554
R1001 B.n545 B.n44 76.0554
R1002 B.n545 B.n544 76.0554
R1003 B.n543 B.n51 76.0554
R1004 B.n537 B.n51 76.0554
R1005 B.n537 B.n536 76.0554
R1006 B.n536 B.n535 76.0554
R1007 B.n535 B.n58 76.0554
R1008 B.n529 B.n58 76.0554
R1009 B.n529 B.n528 76.0554
R1010 B.n94 B.n64 71.676
R1011 B.n98 B.n65 71.676
R1012 B.n102 B.n66 71.676
R1013 B.n106 B.n67 71.676
R1014 B.n110 B.n68 71.676
R1015 B.n114 B.n69 71.676
R1016 B.n118 B.n70 71.676
R1017 B.n122 B.n71 71.676
R1018 B.n126 B.n72 71.676
R1019 B.n130 B.n73 71.676
R1020 B.n134 B.n74 71.676
R1021 B.n138 B.n75 71.676
R1022 B.n142 B.n76 71.676
R1023 B.n146 B.n77 71.676
R1024 B.n150 B.n78 71.676
R1025 B.n155 B.n79 71.676
R1026 B.n159 B.n80 71.676
R1027 B.n163 B.n81 71.676
R1028 B.n167 B.n82 71.676
R1029 B.n171 B.n83 71.676
R1030 B.n175 B.n84 71.676
R1031 B.n179 B.n85 71.676
R1032 B.n183 B.n86 71.676
R1033 B.n187 B.n87 71.676
R1034 B.n88 B.n87 71.676
R1035 B.n186 B.n86 71.676
R1036 B.n182 B.n85 71.676
R1037 B.n178 B.n84 71.676
R1038 B.n174 B.n83 71.676
R1039 B.n170 B.n82 71.676
R1040 B.n166 B.n81 71.676
R1041 B.n162 B.n80 71.676
R1042 B.n158 B.n79 71.676
R1043 B.n154 B.n78 71.676
R1044 B.n149 B.n77 71.676
R1045 B.n145 B.n76 71.676
R1046 B.n141 B.n75 71.676
R1047 B.n137 B.n74 71.676
R1048 B.n133 B.n73 71.676
R1049 B.n129 B.n72 71.676
R1050 B.n125 B.n71 71.676
R1051 B.n121 B.n70 71.676
R1052 B.n117 B.n69 71.676
R1053 B.n113 B.n68 71.676
R1054 B.n109 B.n67 71.676
R1055 B.n105 B.n66 71.676
R1056 B.n101 B.n65 71.676
R1057 B.n97 B.n64 71.676
R1058 B.n378 B.n377 71.676
R1059 B.n372 B.n256 71.676
R1060 B.n369 B.n257 71.676
R1061 B.n365 B.n258 71.676
R1062 B.n361 B.n259 71.676
R1063 B.n357 B.n260 71.676
R1064 B.n353 B.n261 71.676
R1065 B.n349 B.n262 71.676
R1066 B.n345 B.n263 71.676
R1067 B.n341 B.n264 71.676
R1068 B.n336 B.n265 71.676
R1069 B.n332 B.n266 71.676
R1070 B.n328 B.n267 71.676
R1071 B.n324 B.n268 71.676
R1072 B.n320 B.n269 71.676
R1073 B.n316 B.n270 71.676
R1074 B.n312 B.n271 71.676
R1075 B.n308 B.n272 71.676
R1076 B.n304 B.n273 71.676
R1077 B.n300 B.n274 71.676
R1078 B.n296 B.n275 71.676
R1079 B.n292 B.n276 71.676
R1080 B.n288 B.n277 71.676
R1081 B.n380 B.n255 71.676
R1082 B.n378 B.n279 71.676
R1083 B.n370 B.n256 71.676
R1084 B.n366 B.n257 71.676
R1085 B.n362 B.n258 71.676
R1086 B.n358 B.n259 71.676
R1087 B.n354 B.n260 71.676
R1088 B.n350 B.n261 71.676
R1089 B.n346 B.n262 71.676
R1090 B.n342 B.n263 71.676
R1091 B.n337 B.n264 71.676
R1092 B.n333 B.n265 71.676
R1093 B.n329 B.n266 71.676
R1094 B.n325 B.n267 71.676
R1095 B.n321 B.n268 71.676
R1096 B.n317 B.n269 71.676
R1097 B.n313 B.n270 71.676
R1098 B.n309 B.n271 71.676
R1099 B.n305 B.n272 71.676
R1100 B.n301 B.n273 71.676
R1101 B.n297 B.n274 71.676
R1102 B.n293 B.n275 71.676
R1103 B.n289 B.n276 71.676
R1104 B.n285 B.n277 71.676
R1105 B.n381 B.n380 71.676
R1106 B.n596 B.n595 71.676
R1107 B.n596 B.n2 71.676
R1108 B.n93 B.n92 59.5399
R1109 B.n152 B.n90 59.5399
R1110 B.n284 B.n283 59.5399
R1111 B.n339 B.n281 59.5399
R1112 B.t0 B.n212 58.1601
R1113 B.n568 B.t2 58.1601
R1114 B.n92 B.n91 55.6611
R1115 B.n90 B.n89 55.6611
R1116 B.n283 B.n282 55.6611
R1117 B.n281 B.n280 55.6611
R1118 B.n464 B.t1 51.4494
R1119 B.t3 B.n583 51.4494
R1120 B.n404 B.t9 44.7387
R1121 B.t5 B.n543 44.7387
R1122 B.n376 B.n250 32.0005
R1123 B.n383 B.n382 32.0005
R1124 B.n525 B.n524 32.0005
R1125 B.n95 B.n60 32.0005
R1126 B.t9 B.n236 31.3172
R1127 B.n544 B.t5 31.3172
R1128 B.t1 B.n196 24.6065
R1129 B.n584 B.t3 24.6065
R1130 B B.n597 18.0485
R1131 B.n440 B.t0 17.8958
R1132 B.t2 B.n567 17.8958
R1133 B.n388 B.n250 10.6151
R1134 B.n389 B.n388 10.6151
R1135 B.n390 B.n389 10.6151
R1136 B.n390 B.n242 10.6151
R1137 B.n400 B.n242 10.6151
R1138 B.n401 B.n400 10.6151
R1139 B.n402 B.n401 10.6151
R1140 B.n402 B.n234 10.6151
R1141 B.n412 B.n234 10.6151
R1142 B.n413 B.n412 10.6151
R1143 B.n414 B.n413 10.6151
R1144 B.n414 B.n226 10.6151
R1145 B.n424 B.n226 10.6151
R1146 B.n425 B.n424 10.6151
R1147 B.n426 B.n425 10.6151
R1148 B.n426 B.n218 10.6151
R1149 B.n436 B.n218 10.6151
R1150 B.n437 B.n436 10.6151
R1151 B.n438 B.n437 10.6151
R1152 B.n438 B.n210 10.6151
R1153 B.n448 B.n210 10.6151
R1154 B.n449 B.n448 10.6151
R1155 B.n450 B.n449 10.6151
R1156 B.n450 B.n202 10.6151
R1157 B.n460 B.n202 10.6151
R1158 B.n461 B.n460 10.6151
R1159 B.n462 B.n461 10.6151
R1160 B.n462 B.n194 10.6151
R1161 B.n473 B.n194 10.6151
R1162 B.n474 B.n473 10.6151
R1163 B.n475 B.n474 10.6151
R1164 B.n475 B.n0 10.6151
R1165 B.n376 B.n375 10.6151
R1166 B.n375 B.n374 10.6151
R1167 B.n374 B.n373 10.6151
R1168 B.n373 B.n371 10.6151
R1169 B.n371 B.n368 10.6151
R1170 B.n368 B.n367 10.6151
R1171 B.n367 B.n364 10.6151
R1172 B.n364 B.n363 10.6151
R1173 B.n363 B.n360 10.6151
R1174 B.n360 B.n359 10.6151
R1175 B.n359 B.n356 10.6151
R1176 B.n356 B.n355 10.6151
R1177 B.n355 B.n352 10.6151
R1178 B.n352 B.n351 10.6151
R1179 B.n351 B.n348 10.6151
R1180 B.n348 B.n347 10.6151
R1181 B.n347 B.n344 10.6151
R1182 B.n344 B.n343 10.6151
R1183 B.n343 B.n340 10.6151
R1184 B.n338 B.n335 10.6151
R1185 B.n335 B.n334 10.6151
R1186 B.n334 B.n331 10.6151
R1187 B.n331 B.n330 10.6151
R1188 B.n330 B.n327 10.6151
R1189 B.n327 B.n326 10.6151
R1190 B.n326 B.n323 10.6151
R1191 B.n323 B.n322 10.6151
R1192 B.n319 B.n318 10.6151
R1193 B.n318 B.n315 10.6151
R1194 B.n315 B.n314 10.6151
R1195 B.n314 B.n311 10.6151
R1196 B.n311 B.n310 10.6151
R1197 B.n310 B.n307 10.6151
R1198 B.n307 B.n306 10.6151
R1199 B.n306 B.n303 10.6151
R1200 B.n303 B.n302 10.6151
R1201 B.n302 B.n299 10.6151
R1202 B.n299 B.n298 10.6151
R1203 B.n298 B.n295 10.6151
R1204 B.n295 B.n294 10.6151
R1205 B.n294 B.n291 10.6151
R1206 B.n291 B.n290 10.6151
R1207 B.n290 B.n287 10.6151
R1208 B.n287 B.n286 10.6151
R1209 B.n286 B.n254 10.6151
R1210 B.n382 B.n254 10.6151
R1211 B.n384 B.n383 10.6151
R1212 B.n384 B.n246 10.6151
R1213 B.n394 B.n246 10.6151
R1214 B.n395 B.n394 10.6151
R1215 B.n396 B.n395 10.6151
R1216 B.n396 B.n238 10.6151
R1217 B.n406 B.n238 10.6151
R1218 B.n407 B.n406 10.6151
R1219 B.n408 B.n407 10.6151
R1220 B.n408 B.n230 10.6151
R1221 B.n418 B.n230 10.6151
R1222 B.n419 B.n418 10.6151
R1223 B.n420 B.n419 10.6151
R1224 B.n420 B.n222 10.6151
R1225 B.n430 B.n222 10.6151
R1226 B.n431 B.n430 10.6151
R1227 B.n432 B.n431 10.6151
R1228 B.n432 B.n214 10.6151
R1229 B.n442 B.n214 10.6151
R1230 B.n443 B.n442 10.6151
R1231 B.n444 B.n443 10.6151
R1232 B.n444 B.n206 10.6151
R1233 B.n454 B.n206 10.6151
R1234 B.n455 B.n454 10.6151
R1235 B.n456 B.n455 10.6151
R1236 B.n456 B.n198 10.6151
R1237 B.n466 B.n198 10.6151
R1238 B.n467 B.n466 10.6151
R1239 B.n469 B.n467 10.6151
R1240 B.n469 B.n468 10.6151
R1241 B.n468 B.n190 10.6151
R1242 B.n480 B.n190 10.6151
R1243 B.n481 B.n480 10.6151
R1244 B.n482 B.n481 10.6151
R1245 B.n483 B.n482 10.6151
R1246 B.n484 B.n483 10.6151
R1247 B.n487 B.n484 10.6151
R1248 B.n488 B.n487 10.6151
R1249 B.n489 B.n488 10.6151
R1250 B.n490 B.n489 10.6151
R1251 B.n492 B.n490 10.6151
R1252 B.n493 B.n492 10.6151
R1253 B.n494 B.n493 10.6151
R1254 B.n495 B.n494 10.6151
R1255 B.n497 B.n495 10.6151
R1256 B.n498 B.n497 10.6151
R1257 B.n499 B.n498 10.6151
R1258 B.n500 B.n499 10.6151
R1259 B.n502 B.n500 10.6151
R1260 B.n503 B.n502 10.6151
R1261 B.n504 B.n503 10.6151
R1262 B.n505 B.n504 10.6151
R1263 B.n507 B.n505 10.6151
R1264 B.n508 B.n507 10.6151
R1265 B.n509 B.n508 10.6151
R1266 B.n510 B.n509 10.6151
R1267 B.n512 B.n510 10.6151
R1268 B.n513 B.n512 10.6151
R1269 B.n514 B.n513 10.6151
R1270 B.n515 B.n514 10.6151
R1271 B.n517 B.n515 10.6151
R1272 B.n518 B.n517 10.6151
R1273 B.n519 B.n518 10.6151
R1274 B.n520 B.n519 10.6151
R1275 B.n522 B.n520 10.6151
R1276 B.n523 B.n522 10.6151
R1277 B.n524 B.n523 10.6151
R1278 B.n589 B.n1 10.6151
R1279 B.n589 B.n588 10.6151
R1280 B.n588 B.n587 10.6151
R1281 B.n587 B.n10 10.6151
R1282 B.n581 B.n10 10.6151
R1283 B.n581 B.n580 10.6151
R1284 B.n580 B.n579 10.6151
R1285 B.n579 B.n18 10.6151
R1286 B.n573 B.n18 10.6151
R1287 B.n573 B.n572 10.6151
R1288 B.n572 B.n571 10.6151
R1289 B.n571 B.n25 10.6151
R1290 B.n565 B.n25 10.6151
R1291 B.n565 B.n564 10.6151
R1292 B.n564 B.n563 10.6151
R1293 B.n563 B.n32 10.6151
R1294 B.n557 B.n32 10.6151
R1295 B.n557 B.n556 10.6151
R1296 B.n556 B.n555 10.6151
R1297 B.n555 B.n39 10.6151
R1298 B.n549 B.n39 10.6151
R1299 B.n549 B.n548 10.6151
R1300 B.n548 B.n547 10.6151
R1301 B.n547 B.n46 10.6151
R1302 B.n541 B.n46 10.6151
R1303 B.n541 B.n540 10.6151
R1304 B.n540 B.n539 10.6151
R1305 B.n539 B.n53 10.6151
R1306 B.n533 B.n53 10.6151
R1307 B.n533 B.n532 10.6151
R1308 B.n532 B.n531 10.6151
R1309 B.n531 B.n60 10.6151
R1310 B.n96 B.n95 10.6151
R1311 B.n99 B.n96 10.6151
R1312 B.n100 B.n99 10.6151
R1313 B.n103 B.n100 10.6151
R1314 B.n104 B.n103 10.6151
R1315 B.n107 B.n104 10.6151
R1316 B.n108 B.n107 10.6151
R1317 B.n111 B.n108 10.6151
R1318 B.n112 B.n111 10.6151
R1319 B.n115 B.n112 10.6151
R1320 B.n116 B.n115 10.6151
R1321 B.n119 B.n116 10.6151
R1322 B.n120 B.n119 10.6151
R1323 B.n123 B.n120 10.6151
R1324 B.n124 B.n123 10.6151
R1325 B.n127 B.n124 10.6151
R1326 B.n128 B.n127 10.6151
R1327 B.n131 B.n128 10.6151
R1328 B.n132 B.n131 10.6151
R1329 B.n136 B.n135 10.6151
R1330 B.n139 B.n136 10.6151
R1331 B.n140 B.n139 10.6151
R1332 B.n143 B.n140 10.6151
R1333 B.n144 B.n143 10.6151
R1334 B.n147 B.n144 10.6151
R1335 B.n148 B.n147 10.6151
R1336 B.n151 B.n148 10.6151
R1337 B.n156 B.n153 10.6151
R1338 B.n157 B.n156 10.6151
R1339 B.n160 B.n157 10.6151
R1340 B.n161 B.n160 10.6151
R1341 B.n164 B.n161 10.6151
R1342 B.n165 B.n164 10.6151
R1343 B.n168 B.n165 10.6151
R1344 B.n169 B.n168 10.6151
R1345 B.n172 B.n169 10.6151
R1346 B.n173 B.n172 10.6151
R1347 B.n176 B.n173 10.6151
R1348 B.n177 B.n176 10.6151
R1349 B.n180 B.n177 10.6151
R1350 B.n181 B.n180 10.6151
R1351 B.n184 B.n181 10.6151
R1352 B.n185 B.n184 10.6151
R1353 B.n188 B.n185 10.6151
R1354 B.n189 B.n188 10.6151
R1355 B.n525 B.n189 10.6151
R1356 B.n597 B.n0 8.11757
R1357 B.n597 B.n1 8.11757
R1358 B.n339 B.n338 6.5566
R1359 B.n322 B.n284 6.5566
R1360 B.n135 B.n93 6.5566
R1361 B.n152 B.n151 6.5566
R1362 B.n340 B.n339 4.05904
R1363 B.n319 B.n284 4.05904
R1364 B.n132 B.n93 4.05904
R1365 B.n153 B.n152 4.05904
R1366 VN.n0 VN.t0 79.0883
R1367 VN.n1 VN.t2 79.0883
R1368 VN.n0 VN.t3 78.3227
R1369 VN.n1 VN.t1 78.3227
R1370 VN VN.n1 45.182
R1371 VN VN.n0 4.43574
R1372 VDD2.n2 VDD2.n0 105.71
R1373 VDD2.n2 VDD2.n1 70.6417
R1374 VDD2.n1 VDD2.t2 4.34261
R1375 VDD2.n1 VDD2.t1 4.34261
R1376 VDD2.n0 VDD2.t3 4.34261
R1377 VDD2.n0 VDD2.t0 4.34261
R1378 VDD2 VDD2.n2 0.0586897
C0 VTAIL VP 2.37079f
C1 VDD2 VN 1.99358f
C2 VTAIL VDD1 3.61275f
C3 VTAIL VDD2 3.66655f
C4 VTAIL VN 2.35669f
C5 VDD1 VP 2.23434f
C6 VDD2 VP 0.395311f
C7 VP VN 4.771471f
C8 VDD2 VDD1 1.01961f
C9 VDD1 VN 0.153384f
C10 VDD2 B 3.067492f
C11 VDD1 B 6.53016f
C12 VTAIL B 5.318185f
C13 VN B 9.5734f
C14 VP B 8.13698f
C15 VDD2.t3 B 0.065702f
C16 VDD2.t0 B 0.065702f
C17 VDD2.n0 B 0.79187f
C18 VDD2.t2 B 0.065702f
C19 VDD2.t1 B 0.065702f
C20 VDD2.n1 B 0.527799f
C21 VDD2.n2 B 1.96824f
C22 VN.t0 B 0.917455f
C23 VN.t3 B 0.913359f
C24 VN.n0 B 0.573381f
C25 VN.t2 B 0.917455f
C26 VN.t1 B 0.913359f
C27 VN.n1 B 1.64223f
C28 VDD1.t2 B 0.101151f
C29 VDD1.t3 B 0.101151f
C30 VDD1.n0 B 0.812951f
C31 VDD1.t0 B 0.101151f
C32 VDD1.t1 B 0.101151f
C33 VDD1.n1 B 1.24216f
C34 VTAIL.n0 B 0.028736f
C35 VTAIL.n1 B 0.021261f
C36 VTAIL.n2 B 0.011425f
C37 VTAIL.n3 B 0.027004f
C38 VTAIL.n4 B 0.012097f
C39 VTAIL.n5 B 0.364608f
C40 VTAIL.n6 B 0.011425f
C41 VTAIL.t3 B 0.044253f
C42 VTAIL.n7 B 0.083932f
C43 VTAIL.n8 B 0.015936f
C44 VTAIL.n9 B 0.020253f
C45 VTAIL.n10 B 0.027004f
C46 VTAIL.n11 B 0.012097f
C47 VTAIL.n12 B 0.011425f
C48 VTAIL.n13 B 0.021261f
C49 VTAIL.n14 B 0.021261f
C50 VTAIL.n15 B 0.011425f
C51 VTAIL.n16 B 0.012097f
C52 VTAIL.n17 B 0.027004f
C53 VTAIL.n18 B 0.056429f
C54 VTAIL.n19 B 0.012097f
C55 VTAIL.n20 B 0.011425f
C56 VTAIL.n21 B 0.049143f
C57 VTAIL.n22 B 0.031366f
C58 VTAIL.n23 B 0.139078f
C59 VTAIL.n24 B 0.028736f
C60 VTAIL.n25 B 0.021261f
C61 VTAIL.n26 B 0.011425f
C62 VTAIL.n27 B 0.027004f
C63 VTAIL.n28 B 0.012097f
C64 VTAIL.n29 B 0.364608f
C65 VTAIL.n30 B 0.011425f
C66 VTAIL.t7 B 0.044253f
C67 VTAIL.n31 B 0.083932f
C68 VTAIL.n32 B 0.015936f
C69 VTAIL.n33 B 0.020253f
C70 VTAIL.n34 B 0.027004f
C71 VTAIL.n35 B 0.012097f
C72 VTAIL.n36 B 0.011425f
C73 VTAIL.n37 B 0.021261f
C74 VTAIL.n38 B 0.021261f
C75 VTAIL.n39 B 0.011425f
C76 VTAIL.n40 B 0.012097f
C77 VTAIL.n41 B 0.027004f
C78 VTAIL.n42 B 0.056429f
C79 VTAIL.n43 B 0.012097f
C80 VTAIL.n44 B 0.011425f
C81 VTAIL.n45 B 0.049143f
C82 VTAIL.n46 B 0.031366f
C83 VTAIL.n47 B 0.219839f
C84 VTAIL.n48 B 0.028736f
C85 VTAIL.n49 B 0.021261f
C86 VTAIL.n50 B 0.011425f
C87 VTAIL.n51 B 0.027004f
C88 VTAIL.n52 B 0.012097f
C89 VTAIL.n53 B 0.364608f
C90 VTAIL.n54 B 0.011425f
C91 VTAIL.t4 B 0.044253f
C92 VTAIL.n55 B 0.083932f
C93 VTAIL.n56 B 0.015936f
C94 VTAIL.n57 B 0.020253f
C95 VTAIL.n58 B 0.027004f
C96 VTAIL.n59 B 0.012097f
C97 VTAIL.n60 B 0.011425f
C98 VTAIL.n61 B 0.021261f
C99 VTAIL.n62 B 0.021261f
C100 VTAIL.n63 B 0.011425f
C101 VTAIL.n64 B 0.012097f
C102 VTAIL.n65 B 0.027004f
C103 VTAIL.n66 B 0.056429f
C104 VTAIL.n67 B 0.012097f
C105 VTAIL.n68 B 0.011425f
C106 VTAIL.n69 B 0.049143f
C107 VTAIL.n70 B 0.031366f
C108 VTAIL.n71 B 0.91525f
C109 VTAIL.n72 B 0.028736f
C110 VTAIL.n73 B 0.021261f
C111 VTAIL.n74 B 0.011425f
C112 VTAIL.n75 B 0.027004f
C113 VTAIL.n76 B 0.012097f
C114 VTAIL.n77 B 0.364608f
C115 VTAIL.n78 B 0.011425f
C116 VTAIL.t0 B 0.044253f
C117 VTAIL.n79 B 0.083932f
C118 VTAIL.n80 B 0.015936f
C119 VTAIL.n81 B 0.020253f
C120 VTAIL.n82 B 0.027004f
C121 VTAIL.n83 B 0.012097f
C122 VTAIL.n84 B 0.011425f
C123 VTAIL.n85 B 0.021261f
C124 VTAIL.n86 B 0.021261f
C125 VTAIL.n87 B 0.011425f
C126 VTAIL.n88 B 0.012097f
C127 VTAIL.n89 B 0.027004f
C128 VTAIL.n90 B 0.056429f
C129 VTAIL.n91 B 0.012097f
C130 VTAIL.n92 B 0.011425f
C131 VTAIL.n93 B 0.049143f
C132 VTAIL.n94 B 0.031366f
C133 VTAIL.n95 B 0.91525f
C134 VTAIL.n96 B 0.028736f
C135 VTAIL.n97 B 0.021261f
C136 VTAIL.n98 B 0.011425f
C137 VTAIL.n99 B 0.027004f
C138 VTAIL.n100 B 0.012097f
C139 VTAIL.n101 B 0.364608f
C140 VTAIL.n102 B 0.011425f
C141 VTAIL.t1 B 0.044253f
C142 VTAIL.n103 B 0.083932f
C143 VTAIL.n104 B 0.015936f
C144 VTAIL.n105 B 0.020253f
C145 VTAIL.n106 B 0.027004f
C146 VTAIL.n107 B 0.012097f
C147 VTAIL.n108 B 0.011425f
C148 VTAIL.n109 B 0.021261f
C149 VTAIL.n110 B 0.021261f
C150 VTAIL.n111 B 0.011425f
C151 VTAIL.n112 B 0.012097f
C152 VTAIL.n113 B 0.027004f
C153 VTAIL.n114 B 0.056429f
C154 VTAIL.n115 B 0.012097f
C155 VTAIL.n116 B 0.011425f
C156 VTAIL.n117 B 0.049143f
C157 VTAIL.n118 B 0.031366f
C158 VTAIL.n119 B 0.219839f
C159 VTAIL.n120 B 0.028736f
C160 VTAIL.n121 B 0.021261f
C161 VTAIL.n122 B 0.011425f
C162 VTAIL.n123 B 0.027004f
C163 VTAIL.n124 B 0.012097f
C164 VTAIL.n125 B 0.364608f
C165 VTAIL.n126 B 0.011425f
C166 VTAIL.t5 B 0.044253f
C167 VTAIL.n127 B 0.083932f
C168 VTAIL.n128 B 0.015936f
C169 VTAIL.n129 B 0.020253f
C170 VTAIL.n130 B 0.027004f
C171 VTAIL.n131 B 0.012097f
C172 VTAIL.n132 B 0.011425f
C173 VTAIL.n133 B 0.021261f
C174 VTAIL.n134 B 0.021261f
C175 VTAIL.n135 B 0.011425f
C176 VTAIL.n136 B 0.012097f
C177 VTAIL.n137 B 0.027004f
C178 VTAIL.n138 B 0.056429f
C179 VTAIL.n139 B 0.012097f
C180 VTAIL.n140 B 0.011425f
C181 VTAIL.n141 B 0.049143f
C182 VTAIL.n142 B 0.031366f
C183 VTAIL.n143 B 0.219839f
C184 VTAIL.n144 B 0.028736f
C185 VTAIL.n145 B 0.021261f
C186 VTAIL.n146 B 0.011425f
C187 VTAIL.n147 B 0.027004f
C188 VTAIL.n148 B 0.012097f
C189 VTAIL.n149 B 0.364608f
C190 VTAIL.n150 B 0.011425f
C191 VTAIL.t6 B 0.044253f
C192 VTAIL.n151 B 0.083932f
C193 VTAIL.n152 B 0.015936f
C194 VTAIL.n153 B 0.020253f
C195 VTAIL.n154 B 0.027004f
C196 VTAIL.n155 B 0.012097f
C197 VTAIL.n156 B 0.011425f
C198 VTAIL.n157 B 0.021261f
C199 VTAIL.n158 B 0.021261f
C200 VTAIL.n159 B 0.011425f
C201 VTAIL.n160 B 0.012097f
C202 VTAIL.n161 B 0.027004f
C203 VTAIL.n162 B 0.056429f
C204 VTAIL.n163 B 0.012097f
C205 VTAIL.n164 B 0.011425f
C206 VTAIL.n165 B 0.049143f
C207 VTAIL.n166 B 0.031366f
C208 VTAIL.n167 B 0.91525f
C209 VTAIL.n168 B 0.028736f
C210 VTAIL.n169 B 0.021261f
C211 VTAIL.n170 B 0.011425f
C212 VTAIL.n171 B 0.027004f
C213 VTAIL.n172 B 0.012097f
C214 VTAIL.n173 B 0.364608f
C215 VTAIL.n174 B 0.011425f
C216 VTAIL.t2 B 0.044253f
C217 VTAIL.n175 B 0.083932f
C218 VTAIL.n176 B 0.015936f
C219 VTAIL.n177 B 0.020253f
C220 VTAIL.n178 B 0.027004f
C221 VTAIL.n179 B 0.012097f
C222 VTAIL.n180 B 0.011425f
C223 VTAIL.n181 B 0.021261f
C224 VTAIL.n182 B 0.021261f
C225 VTAIL.n183 B 0.011425f
C226 VTAIL.n184 B 0.012097f
C227 VTAIL.n185 B 0.027004f
C228 VTAIL.n186 B 0.056429f
C229 VTAIL.n187 B 0.012097f
C230 VTAIL.n188 B 0.011425f
C231 VTAIL.n189 B 0.049143f
C232 VTAIL.n190 B 0.031366f
C233 VTAIL.n191 B 0.826516f
C234 VP.n0 B 0.041463f
C235 VP.t2 B 0.946258f
C236 VP.n1 B 0.045719f
C237 VP.n2 B 0.031451f
C238 VP.t3 B 0.946258f
C239 VP.n3 B 0.469779f
C240 VP.t0 B 1.19805f
C241 VP.t1 B 1.20342f
C242 VP.n4 B 2.13735f
C243 VP.n5 B 1.44217f
C244 VP.n6 B 0.041463f
C245 VP.n7 B 0.040184f
C246 VP.n8 B 0.058323f
C247 VP.n9 B 0.045719f
C248 VP.n10 B 0.031451f
C249 VP.n11 B 0.031451f
C250 VP.n12 B 0.031451f
C251 VP.n13 B 0.058323f
C252 VP.n14 B 0.040184f
C253 VP.n15 B 0.469779f
C254 VP.n16 B 0.051283f
.ends

