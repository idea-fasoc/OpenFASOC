* NGSPICE file created from diff_pair_sample_1648.ext - technology: sky130A

.subckt diff_pair_sample_1648 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t5 VP.t0 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=5.5185 pd=29.08 as=2.33475 ps=14.48 w=14.15 l=2.01
X1 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=5.5185 pd=29.08 as=0 ps=0 w=14.15 l=2.01
X2 VDD1.t1 VP.t1 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.33475 pd=14.48 as=5.5185 ps=29.08 w=14.15 l=2.01
X3 VDD1.t0 VP.t2 VTAIL.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=2.33475 pd=14.48 as=5.5185 ps=29.08 w=14.15 l=2.01
X4 VTAIL.t1 VN.t0 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=5.5185 pd=29.08 as=2.33475 ps=14.48 w=14.15 l=2.01
X5 VDD2.t2 VN.t1 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=2.33475 pd=14.48 as=5.5185 ps=29.08 w=14.15 l=2.01
X6 VTAIL.t2 VP.t3 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=5.5185 pd=29.08 as=2.33475 ps=14.48 w=14.15 l=2.01
X7 VDD2.t1 VN.t2 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.33475 pd=14.48 as=5.5185 ps=29.08 w=14.15 l=2.01
X8 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=5.5185 pd=29.08 as=0 ps=0 w=14.15 l=2.01
X9 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=5.5185 pd=29.08 as=0 ps=0 w=14.15 l=2.01
X10 VTAIL.t0 VN.t3 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.5185 pd=29.08 as=2.33475 ps=14.48 w=14.15 l=2.01
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.5185 pd=29.08 as=0 ps=0 w=14.15 l=2.01
R0 VP.n2 VP.t3 205.304
R1 VP.n2 VP.t1 204.77
R2 VP.n4 VP.t0 169.66
R3 VP.n11 VP.t2 169.66
R4 VP.n10 VP.n0 161.3
R5 VP.n9 VP.n8 161.3
R6 VP.n7 VP.n1 161.3
R7 VP.n6 VP.n5 161.3
R8 VP.n4 VP.n3 90.2042
R9 VP.n12 VP.n11 90.2042
R10 VP.n9 VP.n1 56.5193
R11 VP.n3 VP.n2 53.3438
R12 VP.n5 VP.n1 24.4675
R13 VP.n10 VP.n9 24.4675
R14 VP.n5 VP.n4 20.5528
R15 VP.n11 VP.n10 20.5528
R16 VP.n6 VP.n3 0.278367
R17 VP.n12 VP.n0 0.278367
R18 VP.n7 VP.n6 0.189894
R19 VP.n8 VP.n7 0.189894
R20 VP.n8 VP.n0 0.189894
R21 VP VP.n12 0.153454
R22 VDD1 VDD1.n1 107.965
R23 VDD1 VDD1.n0 65.533
R24 VDD1.n0 VDD1.t3 1.39979
R25 VDD1.n0 VDD1.t1 1.39979
R26 VDD1.n1 VDD1.t2 1.39979
R27 VDD1.n1 VDD1.t0 1.39979
R28 VTAIL.n618 VTAIL.n546 289.615
R29 VTAIL.n72 VTAIL.n0 289.615
R30 VTAIL.n150 VTAIL.n78 289.615
R31 VTAIL.n228 VTAIL.n156 289.615
R32 VTAIL.n540 VTAIL.n468 289.615
R33 VTAIL.n462 VTAIL.n390 289.615
R34 VTAIL.n384 VTAIL.n312 289.615
R35 VTAIL.n306 VTAIL.n234 289.615
R36 VTAIL.n570 VTAIL.n569 185
R37 VTAIL.n575 VTAIL.n574 185
R38 VTAIL.n577 VTAIL.n576 185
R39 VTAIL.n566 VTAIL.n565 185
R40 VTAIL.n583 VTAIL.n582 185
R41 VTAIL.n585 VTAIL.n584 185
R42 VTAIL.n562 VTAIL.n561 185
R43 VTAIL.n591 VTAIL.n590 185
R44 VTAIL.n593 VTAIL.n592 185
R45 VTAIL.n558 VTAIL.n557 185
R46 VTAIL.n599 VTAIL.n598 185
R47 VTAIL.n601 VTAIL.n600 185
R48 VTAIL.n554 VTAIL.n553 185
R49 VTAIL.n607 VTAIL.n606 185
R50 VTAIL.n609 VTAIL.n608 185
R51 VTAIL.n550 VTAIL.n549 185
R52 VTAIL.n616 VTAIL.n615 185
R53 VTAIL.n617 VTAIL.n548 185
R54 VTAIL.n619 VTAIL.n618 185
R55 VTAIL.n24 VTAIL.n23 185
R56 VTAIL.n29 VTAIL.n28 185
R57 VTAIL.n31 VTAIL.n30 185
R58 VTAIL.n20 VTAIL.n19 185
R59 VTAIL.n37 VTAIL.n36 185
R60 VTAIL.n39 VTAIL.n38 185
R61 VTAIL.n16 VTAIL.n15 185
R62 VTAIL.n45 VTAIL.n44 185
R63 VTAIL.n47 VTAIL.n46 185
R64 VTAIL.n12 VTAIL.n11 185
R65 VTAIL.n53 VTAIL.n52 185
R66 VTAIL.n55 VTAIL.n54 185
R67 VTAIL.n8 VTAIL.n7 185
R68 VTAIL.n61 VTAIL.n60 185
R69 VTAIL.n63 VTAIL.n62 185
R70 VTAIL.n4 VTAIL.n3 185
R71 VTAIL.n70 VTAIL.n69 185
R72 VTAIL.n71 VTAIL.n2 185
R73 VTAIL.n73 VTAIL.n72 185
R74 VTAIL.n102 VTAIL.n101 185
R75 VTAIL.n107 VTAIL.n106 185
R76 VTAIL.n109 VTAIL.n108 185
R77 VTAIL.n98 VTAIL.n97 185
R78 VTAIL.n115 VTAIL.n114 185
R79 VTAIL.n117 VTAIL.n116 185
R80 VTAIL.n94 VTAIL.n93 185
R81 VTAIL.n123 VTAIL.n122 185
R82 VTAIL.n125 VTAIL.n124 185
R83 VTAIL.n90 VTAIL.n89 185
R84 VTAIL.n131 VTAIL.n130 185
R85 VTAIL.n133 VTAIL.n132 185
R86 VTAIL.n86 VTAIL.n85 185
R87 VTAIL.n139 VTAIL.n138 185
R88 VTAIL.n141 VTAIL.n140 185
R89 VTAIL.n82 VTAIL.n81 185
R90 VTAIL.n148 VTAIL.n147 185
R91 VTAIL.n149 VTAIL.n80 185
R92 VTAIL.n151 VTAIL.n150 185
R93 VTAIL.n180 VTAIL.n179 185
R94 VTAIL.n185 VTAIL.n184 185
R95 VTAIL.n187 VTAIL.n186 185
R96 VTAIL.n176 VTAIL.n175 185
R97 VTAIL.n193 VTAIL.n192 185
R98 VTAIL.n195 VTAIL.n194 185
R99 VTAIL.n172 VTAIL.n171 185
R100 VTAIL.n201 VTAIL.n200 185
R101 VTAIL.n203 VTAIL.n202 185
R102 VTAIL.n168 VTAIL.n167 185
R103 VTAIL.n209 VTAIL.n208 185
R104 VTAIL.n211 VTAIL.n210 185
R105 VTAIL.n164 VTAIL.n163 185
R106 VTAIL.n217 VTAIL.n216 185
R107 VTAIL.n219 VTAIL.n218 185
R108 VTAIL.n160 VTAIL.n159 185
R109 VTAIL.n226 VTAIL.n225 185
R110 VTAIL.n227 VTAIL.n158 185
R111 VTAIL.n229 VTAIL.n228 185
R112 VTAIL.n541 VTAIL.n540 185
R113 VTAIL.n539 VTAIL.n470 185
R114 VTAIL.n538 VTAIL.n537 185
R115 VTAIL.n473 VTAIL.n471 185
R116 VTAIL.n532 VTAIL.n531 185
R117 VTAIL.n530 VTAIL.n529 185
R118 VTAIL.n477 VTAIL.n476 185
R119 VTAIL.n524 VTAIL.n523 185
R120 VTAIL.n522 VTAIL.n521 185
R121 VTAIL.n481 VTAIL.n480 185
R122 VTAIL.n516 VTAIL.n515 185
R123 VTAIL.n514 VTAIL.n513 185
R124 VTAIL.n485 VTAIL.n484 185
R125 VTAIL.n508 VTAIL.n507 185
R126 VTAIL.n506 VTAIL.n505 185
R127 VTAIL.n489 VTAIL.n488 185
R128 VTAIL.n500 VTAIL.n499 185
R129 VTAIL.n498 VTAIL.n497 185
R130 VTAIL.n493 VTAIL.n492 185
R131 VTAIL.n463 VTAIL.n462 185
R132 VTAIL.n461 VTAIL.n392 185
R133 VTAIL.n460 VTAIL.n459 185
R134 VTAIL.n395 VTAIL.n393 185
R135 VTAIL.n454 VTAIL.n453 185
R136 VTAIL.n452 VTAIL.n451 185
R137 VTAIL.n399 VTAIL.n398 185
R138 VTAIL.n446 VTAIL.n445 185
R139 VTAIL.n444 VTAIL.n443 185
R140 VTAIL.n403 VTAIL.n402 185
R141 VTAIL.n438 VTAIL.n437 185
R142 VTAIL.n436 VTAIL.n435 185
R143 VTAIL.n407 VTAIL.n406 185
R144 VTAIL.n430 VTAIL.n429 185
R145 VTAIL.n428 VTAIL.n427 185
R146 VTAIL.n411 VTAIL.n410 185
R147 VTAIL.n422 VTAIL.n421 185
R148 VTAIL.n420 VTAIL.n419 185
R149 VTAIL.n415 VTAIL.n414 185
R150 VTAIL.n385 VTAIL.n384 185
R151 VTAIL.n383 VTAIL.n314 185
R152 VTAIL.n382 VTAIL.n381 185
R153 VTAIL.n317 VTAIL.n315 185
R154 VTAIL.n376 VTAIL.n375 185
R155 VTAIL.n374 VTAIL.n373 185
R156 VTAIL.n321 VTAIL.n320 185
R157 VTAIL.n368 VTAIL.n367 185
R158 VTAIL.n366 VTAIL.n365 185
R159 VTAIL.n325 VTAIL.n324 185
R160 VTAIL.n360 VTAIL.n359 185
R161 VTAIL.n358 VTAIL.n357 185
R162 VTAIL.n329 VTAIL.n328 185
R163 VTAIL.n352 VTAIL.n351 185
R164 VTAIL.n350 VTAIL.n349 185
R165 VTAIL.n333 VTAIL.n332 185
R166 VTAIL.n344 VTAIL.n343 185
R167 VTAIL.n342 VTAIL.n341 185
R168 VTAIL.n337 VTAIL.n336 185
R169 VTAIL.n307 VTAIL.n306 185
R170 VTAIL.n305 VTAIL.n236 185
R171 VTAIL.n304 VTAIL.n303 185
R172 VTAIL.n239 VTAIL.n237 185
R173 VTAIL.n298 VTAIL.n297 185
R174 VTAIL.n296 VTAIL.n295 185
R175 VTAIL.n243 VTAIL.n242 185
R176 VTAIL.n290 VTAIL.n289 185
R177 VTAIL.n288 VTAIL.n287 185
R178 VTAIL.n247 VTAIL.n246 185
R179 VTAIL.n282 VTAIL.n281 185
R180 VTAIL.n280 VTAIL.n279 185
R181 VTAIL.n251 VTAIL.n250 185
R182 VTAIL.n274 VTAIL.n273 185
R183 VTAIL.n272 VTAIL.n271 185
R184 VTAIL.n255 VTAIL.n254 185
R185 VTAIL.n266 VTAIL.n265 185
R186 VTAIL.n264 VTAIL.n263 185
R187 VTAIL.n259 VTAIL.n258 185
R188 VTAIL.n571 VTAIL.t6 147.659
R189 VTAIL.n25 VTAIL.t0 147.659
R190 VTAIL.n103 VTAIL.t3 147.659
R191 VTAIL.n181 VTAIL.t5 147.659
R192 VTAIL.n494 VTAIL.t4 147.659
R193 VTAIL.n416 VTAIL.t2 147.659
R194 VTAIL.n338 VTAIL.t7 147.659
R195 VTAIL.n260 VTAIL.t1 147.659
R196 VTAIL.n575 VTAIL.n569 104.615
R197 VTAIL.n576 VTAIL.n575 104.615
R198 VTAIL.n576 VTAIL.n565 104.615
R199 VTAIL.n583 VTAIL.n565 104.615
R200 VTAIL.n584 VTAIL.n583 104.615
R201 VTAIL.n584 VTAIL.n561 104.615
R202 VTAIL.n591 VTAIL.n561 104.615
R203 VTAIL.n592 VTAIL.n591 104.615
R204 VTAIL.n592 VTAIL.n557 104.615
R205 VTAIL.n599 VTAIL.n557 104.615
R206 VTAIL.n600 VTAIL.n599 104.615
R207 VTAIL.n600 VTAIL.n553 104.615
R208 VTAIL.n607 VTAIL.n553 104.615
R209 VTAIL.n608 VTAIL.n607 104.615
R210 VTAIL.n608 VTAIL.n549 104.615
R211 VTAIL.n616 VTAIL.n549 104.615
R212 VTAIL.n617 VTAIL.n616 104.615
R213 VTAIL.n618 VTAIL.n617 104.615
R214 VTAIL.n29 VTAIL.n23 104.615
R215 VTAIL.n30 VTAIL.n29 104.615
R216 VTAIL.n30 VTAIL.n19 104.615
R217 VTAIL.n37 VTAIL.n19 104.615
R218 VTAIL.n38 VTAIL.n37 104.615
R219 VTAIL.n38 VTAIL.n15 104.615
R220 VTAIL.n45 VTAIL.n15 104.615
R221 VTAIL.n46 VTAIL.n45 104.615
R222 VTAIL.n46 VTAIL.n11 104.615
R223 VTAIL.n53 VTAIL.n11 104.615
R224 VTAIL.n54 VTAIL.n53 104.615
R225 VTAIL.n54 VTAIL.n7 104.615
R226 VTAIL.n61 VTAIL.n7 104.615
R227 VTAIL.n62 VTAIL.n61 104.615
R228 VTAIL.n62 VTAIL.n3 104.615
R229 VTAIL.n70 VTAIL.n3 104.615
R230 VTAIL.n71 VTAIL.n70 104.615
R231 VTAIL.n72 VTAIL.n71 104.615
R232 VTAIL.n107 VTAIL.n101 104.615
R233 VTAIL.n108 VTAIL.n107 104.615
R234 VTAIL.n108 VTAIL.n97 104.615
R235 VTAIL.n115 VTAIL.n97 104.615
R236 VTAIL.n116 VTAIL.n115 104.615
R237 VTAIL.n116 VTAIL.n93 104.615
R238 VTAIL.n123 VTAIL.n93 104.615
R239 VTAIL.n124 VTAIL.n123 104.615
R240 VTAIL.n124 VTAIL.n89 104.615
R241 VTAIL.n131 VTAIL.n89 104.615
R242 VTAIL.n132 VTAIL.n131 104.615
R243 VTAIL.n132 VTAIL.n85 104.615
R244 VTAIL.n139 VTAIL.n85 104.615
R245 VTAIL.n140 VTAIL.n139 104.615
R246 VTAIL.n140 VTAIL.n81 104.615
R247 VTAIL.n148 VTAIL.n81 104.615
R248 VTAIL.n149 VTAIL.n148 104.615
R249 VTAIL.n150 VTAIL.n149 104.615
R250 VTAIL.n185 VTAIL.n179 104.615
R251 VTAIL.n186 VTAIL.n185 104.615
R252 VTAIL.n186 VTAIL.n175 104.615
R253 VTAIL.n193 VTAIL.n175 104.615
R254 VTAIL.n194 VTAIL.n193 104.615
R255 VTAIL.n194 VTAIL.n171 104.615
R256 VTAIL.n201 VTAIL.n171 104.615
R257 VTAIL.n202 VTAIL.n201 104.615
R258 VTAIL.n202 VTAIL.n167 104.615
R259 VTAIL.n209 VTAIL.n167 104.615
R260 VTAIL.n210 VTAIL.n209 104.615
R261 VTAIL.n210 VTAIL.n163 104.615
R262 VTAIL.n217 VTAIL.n163 104.615
R263 VTAIL.n218 VTAIL.n217 104.615
R264 VTAIL.n218 VTAIL.n159 104.615
R265 VTAIL.n226 VTAIL.n159 104.615
R266 VTAIL.n227 VTAIL.n226 104.615
R267 VTAIL.n228 VTAIL.n227 104.615
R268 VTAIL.n540 VTAIL.n539 104.615
R269 VTAIL.n539 VTAIL.n538 104.615
R270 VTAIL.n538 VTAIL.n471 104.615
R271 VTAIL.n531 VTAIL.n471 104.615
R272 VTAIL.n531 VTAIL.n530 104.615
R273 VTAIL.n530 VTAIL.n476 104.615
R274 VTAIL.n523 VTAIL.n476 104.615
R275 VTAIL.n523 VTAIL.n522 104.615
R276 VTAIL.n522 VTAIL.n480 104.615
R277 VTAIL.n515 VTAIL.n480 104.615
R278 VTAIL.n515 VTAIL.n514 104.615
R279 VTAIL.n514 VTAIL.n484 104.615
R280 VTAIL.n507 VTAIL.n484 104.615
R281 VTAIL.n507 VTAIL.n506 104.615
R282 VTAIL.n506 VTAIL.n488 104.615
R283 VTAIL.n499 VTAIL.n488 104.615
R284 VTAIL.n499 VTAIL.n498 104.615
R285 VTAIL.n498 VTAIL.n492 104.615
R286 VTAIL.n462 VTAIL.n461 104.615
R287 VTAIL.n461 VTAIL.n460 104.615
R288 VTAIL.n460 VTAIL.n393 104.615
R289 VTAIL.n453 VTAIL.n393 104.615
R290 VTAIL.n453 VTAIL.n452 104.615
R291 VTAIL.n452 VTAIL.n398 104.615
R292 VTAIL.n445 VTAIL.n398 104.615
R293 VTAIL.n445 VTAIL.n444 104.615
R294 VTAIL.n444 VTAIL.n402 104.615
R295 VTAIL.n437 VTAIL.n402 104.615
R296 VTAIL.n437 VTAIL.n436 104.615
R297 VTAIL.n436 VTAIL.n406 104.615
R298 VTAIL.n429 VTAIL.n406 104.615
R299 VTAIL.n429 VTAIL.n428 104.615
R300 VTAIL.n428 VTAIL.n410 104.615
R301 VTAIL.n421 VTAIL.n410 104.615
R302 VTAIL.n421 VTAIL.n420 104.615
R303 VTAIL.n420 VTAIL.n414 104.615
R304 VTAIL.n384 VTAIL.n383 104.615
R305 VTAIL.n383 VTAIL.n382 104.615
R306 VTAIL.n382 VTAIL.n315 104.615
R307 VTAIL.n375 VTAIL.n315 104.615
R308 VTAIL.n375 VTAIL.n374 104.615
R309 VTAIL.n374 VTAIL.n320 104.615
R310 VTAIL.n367 VTAIL.n320 104.615
R311 VTAIL.n367 VTAIL.n366 104.615
R312 VTAIL.n366 VTAIL.n324 104.615
R313 VTAIL.n359 VTAIL.n324 104.615
R314 VTAIL.n359 VTAIL.n358 104.615
R315 VTAIL.n358 VTAIL.n328 104.615
R316 VTAIL.n351 VTAIL.n328 104.615
R317 VTAIL.n351 VTAIL.n350 104.615
R318 VTAIL.n350 VTAIL.n332 104.615
R319 VTAIL.n343 VTAIL.n332 104.615
R320 VTAIL.n343 VTAIL.n342 104.615
R321 VTAIL.n342 VTAIL.n336 104.615
R322 VTAIL.n306 VTAIL.n305 104.615
R323 VTAIL.n305 VTAIL.n304 104.615
R324 VTAIL.n304 VTAIL.n237 104.615
R325 VTAIL.n297 VTAIL.n237 104.615
R326 VTAIL.n297 VTAIL.n296 104.615
R327 VTAIL.n296 VTAIL.n242 104.615
R328 VTAIL.n289 VTAIL.n242 104.615
R329 VTAIL.n289 VTAIL.n288 104.615
R330 VTAIL.n288 VTAIL.n246 104.615
R331 VTAIL.n281 VTAIL.n246 104.615
R332 VTAIL.n281 VTAIL.n280 104.615
R333 VTAIL.n280 VTAIL.n250 104.615
R334 VTAIL.n273 VTAIL.n250 104.615
R335 VTAIL.n273 VTAIL.n272 104.615
R336 VTAIL.n272 VTAIL.n254 104.615
R337 VTAIL.n265 VTAIL.n254 104.615
R338 VTAIL.n265 VTAIL.n264 104.615
R339 VTAIL.n264 VTAIL.n258 104.615
R340 VTAIL.t6 VTAIL.n569 52.3082
R341 VTAIL.t0 VTAIL.n23 52.3082
R342 VTAIL.t3 VTAIL.n101 52.3082
R343 VTAIL.t5 VTAIL.n179 52.3082
R344 VTAIL.t4 VTAIL.n492 52.3082
R345 VTAIL.t2 VTAIL.n414 52.3082
R346 VTAIL.t7 VTAIL.n336 52.3082
R347 VTAIL.t1 VTAIL.n258 52.3082
R348 VTAIL.n623 VTAIL.n622 36.646
R349 VTAIL.n77 VTAIL.n76 36.646
R350 VTAIL.n155 VTAIL.n154 36.646
R351 VTAIL.n233 VTAIL.n232 36.646
R352 VTAIL.n545 VTAIL.n544 36.646
R353 VTAIL.n467 VTAIL.n466 36.646
R354 VTAIL.n389 VTAIL.n388 36.646
R355 VTAIL.n311 VTAIL.n310 36.646
R356 VTAIL.n623 VTAIL.n545 26.5824
R357 VTAIL.n311 VTAIL.n233 26.5824
R358 VTAIL.n571 VTAIL.n570 15.6677
R359 VTAIL.n25 VTAIL.n24 15.6677
R360 VTAIL.n103 VTAIL.n102 15.6677
R361 VTAIL.n181 VTAIL.n180 15.6677
R362 VTAIL.n494 VTAIL.n493 15.6677
R363 VTAIL.n416 VTAIL.n415 15.6677
R364 VTAIL.n338 VTAIL.n337 15.6677
R365 VTAIL.n260 VTAIL.n259 15.6677
R366 VTAIL.n619 VTAIL.n548 13.1884
R367 VTAIL.n73 VTAIL.n2 13.1884
R368 VTAIL.n151 VTAIL.n80 13.1884
R369 VTAIL.n229 VTAIL.n158 13.1884
R370 VTAIL.n541 VTAIL.n470 13.1884
R371 VTAIL.n463 VTAIL.n392 13.1884
R372 VTAIL.n385 VTAIL.n314 13.1884
R373 VTAIL.n307 VTAIL.n236 13.1884
R374 VTAIL.n574 VTAIL.n573 12.8005
R375 VTAIL.n615 VTAIL.n614 12.8005
R376 VTAIL.n620 VTAIL.n546 12.8005
R377 VTAIL.n28 VTAIL.n27 12.8005
R378 VTAIL.n69 VTAIL.n68 12.8005
R379 VTAIL.n74 VTAIL.n0 12.8005
R380 VTAIL.n106 VTAIL.n105 12.8005
R381 VTAIL.n147 VTAIL.n146 12.8005
R382 VTAIL.n152 VTAIL.n78 12.8005
R383 VTAIL.n184 VTAIL.n183 12.8005
R384 VTAIL.n225 VTAIL.n224 12.8005
R385 VTAIL.n230 VTAIL.n156 12.8005
R386 VTAIL.n542 VTAIL.n468 12.8005
R387 VTAIL.n537 VTAIL.n472 12.8005
R388 VTAIL.n497 VTAIL.n496 12.8005
R389 VTAIL.n464 VTAIL.n390 12.8005
R390 VTAIL.n459 VTAIL.n394 12.8005
R391 VTAIL.n419 VTAIL.n418 12.8005
R392 VTAIL.n386 VTAIL.n312 12.8005
R393 VTAIL.n381 VTAIL.n316 12.8005
R394 VTAIL.n341 VTAIL.n340 12.8005
R395 VTAIL.n308 VTAIL.n234 12.8005
R396 VTAIL.n303 VTAIL.n238 12.8005
R397 VTAIL.n263 VTAIL.n262 12.8005
R398 VTAIL.n577 VTAIL.n568 12.0247
R399 VTAIL.n613 VTAIL.n550 12.0247
R400 VTAIL.n31 VTAIL.n22 12.0247
R401 VTAIL.n67 VTAIL.n4 12.0247
R402 VTAIL.n109 VTAIL.n100 12.0247
R403 VTAIL.n145 VTAIL.n82 12.0247
R404 VTAIL.n187 VTAIL.n178 12.0247
R405 VTAIL.n223 VTAIL.n160 12.0247
R406 VTAIL.n536 VTAIL.n473 12.0247
R407 VTAIL.n500 VTAIL.n491 12.0247
R408 VTAIL.n458 VTAIL.n395 12.0247
R409 VTAIL.n422 VTAIL.n413 12.0247
R410 VTAIL.n380 VTAIL.n317 12.0247
R411 VTAIL.n344 VTAIL.n335 12.0247
R412 VTAIL.n302 VTAIL.n239 12.0247
R413 VTAIL.n266 VTAIL.n257 12.0247
R414 VTAIL.n578 VTAIL.n566 11.249
R415 VTAIL.n610 VTAIL.n609 11.249
R416 VTAIL.n32 VTAIL.n20 11.249
R417 VTAIL.n64 VTAIL.n63 11.249
R418 VTAIL.n110 VTAIL.n98 11.249
R419 VTAIL.n142 VTAIL.n141 11.249
R420 VTAIL.n188 VTAIL.n176 11.249
R421 VTAIL.n220 VTAIL.n219 11.249
R422 VTAIL.n533 VTAIL.n532 11.249
R423 VTAIL.n501 VTAIL.n489 11.249
R424 VTAIL.n455 VTAIL.n454 11.249
R425 VTAIL.n423 VTAIL.n411 11.249
R426 VTAIL.n377 VTAIL.n376 11.249
R427 VTAIL.n345 VTAIL.n333 11.249
R428 VTAIL.n299 VTAIL.n298 11.249
R429 VTAIL.n267 VTAIL.n255 11.249
R430 VTAIL.n582 VTAIL.n581 10.4732
R431 VTAIL.n606 VTAIL.n552 10.4732
R432 VTAIL.n36 VTAIL.n35 10.4732
R433 VTAIL.n60 VTAIL.n6 10.4732
R434 VTAIL.n114 VTAIL.n113 10.4732
R435 VTAIL.n138 VTAIL.n84 10.4732
R436 VTAIL.n192 VTAIL.n191 10.4732
R437 VTAIL.n216 VTAIL.n162 10.4732
R438 VTAIL.n529 VTAIL.n475 10.4732
R439 VTAIL.n505 VTAIL.n504 10.4732
R440 VTAIL.n451 VTAIL.n397 10.4732
R441 VTAIL.n427 VTAIL.n426 10.4732
R442 VTAIL.n373 VTAIL.n319 10.4732
R443 VTAIL.n349 VTAIL.n348 10.4732
R444 VTAIL.n295 VTAIL.n241 10.4732
R445 VTAIL.n271 VTAIL.n270 10.4732
R446 VTAIL.n585 VTAIL.n564 9.69747
R447 VTAIL.n605 VTAIL.n554 9.69747
R448 VTAIL.n39 VTAIL.n18 9.69747
R449 VTAIL.n59 VTAIL.n8 9.69747
R450 VTAIL.n117 VTAIL.n96 9.69747
R451 VTAIL.n137 VTAIL.n86 9.69747
R452 VTAIL.n195 VTAIL.n174 9.69747
R453 VTAIL.n215 VTAIL.n164 9.69747
R454 VTAIL.n528 VTAIL.n477 9.69747
R455 VTAIL.n508 VTAIL.n487 9.69747
R456 VTAIL.n450 VTAIL.n399 9.69747
R457 VTAIL.n430 VTAIL.n409 9.69747
R458 VTAIL.n372 VTAIL.n321 9.69747
R459 VTAIL.n352 VTAIL.n331 9.69747
R460 VTAIL.n294 VTAIL.n243 9.69747
R461 VTAIL.n274 VTAIL.n253 9.69747
R462 VTAIL.n622 VTAIL.n621 9.45567
R463 VTAIL.n76 VTAIL.n75 9.45567
R464 VTAIL.n154 VTAIL.n153 9.45567
R465 VTAIL.n232 VTAIL.n231 9.45567
R466 VTAIL.n544 VTAIL.n543 9.45567
R467 VTAIL.n466 VTAIL.n465 9.45567
R468 VTAIL.n388 VTAIL.n387 9.45567
R469 VTAIL.n310 VTAIL.n309 9.45567
R470 VTAIL.n621 VTAIL.n620 9.3005
R471 VTAIL.n560 VTAIL.n559 9.3005
R472 VTAIL.n589 VTAIL.n588 9.3005
R473 VTAIL.n587 VTAIL.n586 9.3005
R474 VTAIL.n564 VTAIL.n563 9.3005
R475 VTAIL.n581 VTAIL.n580 9.3005
R476 VTAIL.n579 VTAIL.n578 9.3005
R477 VTAIL.n568 VTAIL.n567 9.3005
R478 VTAIL.n573 VTAIL.n572 9.3005
R479 VTAIL.n595 VTAIL.n594 9.3005
R480 VTAIL.n597 VTAIL.n596 9.3005
R481 VTAIL.n556 VTAIL.n555 9.3005
R482 VTAIL.n603 VTAIL.n602 9.3005
R483 VTAIL.n605 VTAIL.n604 9.3005
R484 VTAIL.n552 VTAIL.n551 9.3005
R485 VTAIL.n611 VTAIL.n610 9.3005
R486 VTAIL.n613 VTAIL.n612 9.3005
R487 VTAIL.n614 VTAIL.n547 9.3005
R488 VTAIL.n75 VTAIL.n74 9.3005
R489 VTAIL.n14 VTAIL.n13 9.3005
R490 VTAIL.n43 VTAIL.n42 9.3005
R491 VTAIL.n41 VTAIL.n40 9.3005
R492 VTAIL.n18 VTAIL.n17 9.3005
R493 VTAIL.n35 VTAIL.n34 9.3005
R494 VTAIL.n33 VTAIL.n32 9.3005
R495 VTAIL.n22 VTAIL.n21 9.3005
R496 VTAIL.n27 VTAIL.n26 9.3005
R497 VTAIL.n49 VTAIL.n48 9.3005
R498 VTAIL.n51 VTAIL.n50 9.3005
R499 VTAIL.n10 VTAIL.n9 9.3005
R500 VTAIL.n57 VTAIL.n56 9.3005
R501 VTAIL.n59 VTAIL.n58 9.3005
R502 VTAIL.n6 VTAIL.n5 9.3005
R503 VTAIL.n65 VTAIL.n64 9.3005
R504 VTAIL.n67 VTAIL.n66 9.3005
R505 VTAIL.n68 VTAIL.n1 9.3005
R506 VTAIL.n153 VTAIL.n152 9.3005
R507 VTAIL.n92 VTAIL.n91 9.3005
R508 VTAIL.n121 VTAIL.n120 9.3005
R509 VTAIL.n119 VTAIL.n118 9.3005
R510 VTAIL.n96 VTAIL.n95 9.3005
R511 VTAIL.n113 VTAIL.n112 9.3005
R512 VTAIL.n111 VTAIL.n110 9.3005
R513 VTAIL.n100 VTAIL.n99 9.3005
R514 VTAIL.n105 VTAIL.n104 9.3005
R515 VTAIL.n127 VTAIL.n126 9.3005
R516 VTAIL.n129 VTAIL.n128 9.3005
R517 VTAIL.n88 VTAIL.n87 9.3005
R518 VTAIL.n135 VTAIL.n134 9.3005
R519 VTAIL.n137 VTAIL.n136 9.3005
R520 VTAIL.n84 VTAIL.n83 9.3005
R521 VTAIL.n143 VTAIL.n142 9.3005
R522 VTAIL.n145 VTAIL.n144 9.3005
R523 VTAIL.n146 VTAIL.n79 9.3005
R524 VTAIL.n231 VTAIL.n230 9.3005
R525 VTAIL.n170 VTAIL.n169 9.3005
R526 VTAIL.n199 VTAIL.n198 9.3005
R527 VTAIL.n197 VTAIL.n196 9.3005
R528 VTAIL.n174 VTAIL.n173 9.3005
R529 VTAIL.n191 VTAIL.n190 9.3005
R530 VTAIL.n189 VTAIL.n188 9.3005
R531 VTAIL.n178 VTAIL.n177 9.3005
R532 VTAIL.n183 VTAIL.n182 9.3005
R533 VTAIL.n205 VTAIL.n204 9.3005
R534 VTAIL.n207 VTAIL.n206 9.3005
R535 VTAIL.n166 VTAIL.n165 9.3005
R536 VTAIL.n213 VTAIL.n212 9.3005
R537 VTAIL.n215 VTAIL.n214 9.3005
R538 VTAIL.n162 VTAIL.n161 9.3005
R539 VTAIL.n221 VTAIL.n220 9.3005
R540 VTAIL.n223 VTAIL.n222 9.3005
R541 VTAIL.n224 VTAIL.n157 9.3005
R542 VTAIL.n520 VTAIL.n519 9.3005
R543 VTAIL.n479 VTAIL.n478 9.3005
R544 VTAIL.n526 VTAIL.n525 9.3005
R545 VTAIL.n528 VTAIL.n527 9.3005
R546 VTAIL.n475 VTAIL.n474 9.3005
R547 VTAIL.n534 VTAIL.n533 9.3005
R548 VTAIL.n536 VTAIL.n535 9.3005
R549 VTAIL.n472 VTAIL.n469 9.3005
R550 VTAIL.n543 VTAIL.n542 9.3005
R551 VTAIL.n518 VTAIL.n517 9.3005
R552 VTAIL.n483 VTAIL.n482 9.3005
R553 VTAIL.n512 VTAIL.n511 9.3005
R554 VTAIL.n510 VTAIL.n509 9.3005
R555 VTAIL.n487 VTAIL.n486 9.3005
R556 VTAIL.n504 VTAIL.n503 9.3005
R557 VTAIL.n502 VTAIL.n501 9.3005
R558 VTAIL.n491 VTAIL.n490 9.3005
R559 VTAIL.n496 VTAIL.n495 9.3005
R560 VTAIL.n442 VTAIL.n441 9.3005
R561 VTAIL.n401 VTAIL.n400 9.3005
R562 VTAIL.n448 VTAIL.n447 9.3005
R563 VTAIL.n450 VTAIL.n449 9.3005
R564 VTAIL.n397 VTAIL.n396 9.3005
R565 VTAIL.n456 VTAIL.n455 9.3005
R566 VTAIL.n458 VTAIL.n457 9.3005
R567 VTAIL.n394 VTAIL.n391 9.3005
R568 VTAIL.n465 VTAIL.n464 9.3005
R569 VTAIL.n440 VTAIL.n439 9.3005
R570 VTAIL.n405 VTAIL.n404 9.3005
R571 VTAIL.n434 VTAIL.n433 9.3005
R572 VTAIL.n432 VTAIL.n431 9.3005
R573 VTAIL.n409 VTAIL.n408 9.3005
R574 VTAIL.n426 VTAIL.n425 9.3005
R575 VTAIL.n424 VTAIL.n423 9.3005
R576 VTAIL.n413 VTAIL.n412 9.3005
R577 VTAIL.n418 VTAIL.n417 9.3005
R578 VTAIL.n364 VTAIL.n363 9.3005
R579 VTAIL.n323 VTAIL.n322 9.3005
R580 VTAIL.n370 VTAIL.n369 9.3005
R581 VTAIL.n372 VTAIL.n371 9.3005
R582 VTAIL.n319 VTAIL.n318 9.3005
R583 VTAIL.n378 VTAIL.n377 9.3005
R584 VTAIL.n380 VTAIL.n379 9.3005
R585 VTAIL.n316 VTAIL.n313 9.3005
R586 VTAIL.n387 VTAIL.n386 9.3005
R587 VTAIL.n362 VTAIL.n361 9.3005
R588 VTAIL.n327 VTAIL.n326 9.3005
R589 VTAIL.n356 VTAIL.n355 9.3005
R590 VTAIL.n354 VTAIL.n353 9.3005
R591 VTAIL.n331 VTAIL.n330 9.3005
R592 VTAIL.n348 VTAIL.n347 9.3005
R593 VTAIL.n346 VTAIL.n345 9.3005
R594 VTAIL.n335 VTAIL.n334 9.3005
R595 VTAIL.n340 VTAIL.n339 9.3005
R596 VTAIL.n286 VTAIL.n285 9.3005
R597 VTAIL.n245 VTAIL.n244 9.3005
R598 VTAIL.n292 VTAIL.n291 9.3005
R599 VTAIL.n294 VTAIL.n293 9.3005
R600 VTAIL.n241 VTAIL.n240 9.3005
R601 VTAIL.n300 VTAIL.n299 9.3005
R602 VTAIL.n302 VTAIL.n301 9.3005
R603 VTAIL.n238 VTAIL.n235 9.3005
R604 VTAIL.n309 VTAIL.n308 9.3005
R605 VTAIL.n284 VTAIL.n283 9.3005
R606 VTAIL.n249 VTAIL.n248 9.3005
R607 VTAIL.n278 VTAIL.n277 9.3005
R608 VTAIL.n276 VTAIL.n275 9.3005
R609 VTAIL.n253 VTAIL.n252 9.3005
R610 VTAIL.n270 VTAIL.n269 9.3005
R611 VTAIL.n268 VTAIL.n267 9.3005
R612 VTAIL.n257 VTAIL.n256 9.3005
R613 VTAIL.n262 VTAIL.n261 9.3005
R614 VTAIL.n586 VTAIL.n562 8.92171
R615 VTAIL.n602 VTAIL.n601 8.92171
R616 VTAIL.n40 VTAIL.n16 8.92171
R617 VTAIL.n56 VTAIL.n55 8.92171
R618 VTAIL.n118 VTAIL.n94 8.92171
R619 VTAIL.n134 VTAIL.n133 8.92171
R620 VTAIL.n196 VTAIL.n172 8.92171
R621 VTAIL.n212 VTAIL.n211 8.92171
R622 VTAIL.n525 VTAIL.n524 8.92171
R623 VTAIL.n509 VTAIL.n485 8.92171
R624 VTAIL.n447 VTAIL.n446 8.92171
R625 VTAIL.n431 VTAIL.n407 8.92171
R626 VTAIL.n369 VTAIL.n368 8.92171
R627 VTAIL.n353 VTAIL.n329 8.92171
R628 VTAIL.n291 VTAIL.n290 8.92171
R629 VTAIL.n275 VTAIL.n251 8.92171
R630 VTAIL.n590 VTAIL.n589 8.14595
R631 VTAIL.n598 VTAIL.n556 8.14595
R632 VTAIL.n44 VTAIL.n43 8.14595
R633 VTAIL.n52 VTAIL.n10 8.14595
R634 VTAIL.n122 VTAIL.n121 8.14595
R635 VTAIL.n130 VTAIL.n88 8.14595
R636 VTAIL.n200 VTAIL.n199 8.14595
R637 VTAIL.n208 VTAIL.n166 8.14595
R638 VTAIL.n521 VTAIL.n479 8.14595
R639 VTAIL.n513 VTAIL.n512 8.14595
R640 VTAIL.n443 VTAIL.n401 8.14595
R641 VTAIL.n435 VTAIL.n434 8.14595
R642 VTAIL.n365 VTAIL.n323 8.14595
R643 VTAIL.n357 VTAIL.n356 8.14595
R644 VTAIL.n287 VTAIL.n245 8.14595
R645 VTAIL.n279 VTAIL.n278 8.14595
R646 VTAIL.n593 VTAIL.n560 7.3702
R647 VTAIL.n597 VTAIL.n558 7.3702
R648 VTAIL.n47 VTAIL.n14 7.3702
R649 VTAIL.n51 VTAIL.n12 7.3702
R650 VTAIL.n125 VTAIL.n92 7.3702
R651 VTAIL.n129 VTAIL.n90 7.3702
R652 VTAIL.n203 VTAIL.n170 7.3702
R653 VTAIL.n207 VTAIL.n168 7.3702
R654 VTAIL.n520 VTAIL.n481 7.3702
R655 VTAIL.n516 VTAIL.n483 7.3702
R656 VTAIL.n442 VTAIL.n403 7.3702
R657 VTAIL.n438 VTAIL.n405 7.3702
R658 VTAIL.n364 VTAIL.n325 7.3702
R659 VTAIL.n360 VTAIL.n327 7.3702
R660 VTAIL.n286 VTAIL.n247 7.3702
R661 VTAIL.n282 VTAIL.n249 7.3702
R662 VTAIL.n594 VTAIL.n593 6.59444
R663 VTAIL.n594 VTAIL.n558 6.59444
R664 VTAIL.n48 VTAIL.n47 6.59444
R665 VTAIL.n48 VTAIL.n12 6.59444
R666 VTAIL.n126 VTAIL.n125 6.59444
R667 VTAIL.n126 VTAIL.n90 6.59444
R668 VTAIL.n204 VTAIL.n203 6.59444
R669 VTAIL.n204 VTAIL.n168 6.59444
R670 VTAIL.n517 VTAIL.n481 6.59444
R671 VTAIL.n517 VTAIL.n516 6.59444
R672 VTAIL.n439 VTAIL.n403 6.59444
R673 VTAIL.n439 VTAIL.n438 6.59444
R674 VTAIL.n361 VTAIL.n325 6.59444
R675 VTAIL.n361 VTAIL.n360 6.59444
R676 VTAIL.n283 VTAIL.n247 6.59444
R677 VTAIL.n283 VTAIL.n282 6.59444
R678 VTAIL.n590 VTAIL.n560 5.81868
R679 VTAIL.n598 VTAIL.n597 5.81868
R680 VTAIL.n44 VTAIL.n14 5.81868
R681 VTAIL.n52 VTAIL.n51 5.81868
R682 VTAIL.n122 VTAIL.n92 5.81868
R683 VTAIL.n130 VTAIL.n129 5.81868
R684 VTAIL.n200 VTAIL.n170 5.81868
R685 VTAIL.n208 VTAIL.n207 5.81868
R686 VTAIL.n521 VTAIL.n520 5.81868
R687 VTAIL.n513 VTAIL.n483 5.81868
R688 VTAIL.n443 VTAIL.n442 5.81868
R689 VTAIL.n435 VTAIL.n405 5.81868
R690 VTAIL.n365 VTAIL.n364 5.81868
R691 VTAIL.n357 VTAIL.n327 5.81868
R692 VTAIL.n287 VTAIL.n286 5.81868
R693 VTAIL.n279 VTAIL.n249 5.81868
R694 VTAIL.n589 VTAIL.n562 5.04292
R695 VTAIL.n601 VTAIL.n556 5.04292
R696 VTAIL.n43 VTAIL.n16 5.04292
R697 VTAIL.n55 VTAIL.n10 5.04292
R698 VTAIL.n121 VTAIL.n94 5.04292
R699 VTAIL.n133 VTAIL.n88 5.04292
R700 VTAIL.n199 VTAIL.n172 5.04292
R701 VTAIL.n211 VTAIL.n166 5.04292
R702 VTAIL.n524 VTAIL.n479 5.04292
R703 VTAIL.n512 VTAIL.n485 5.04292
R704 VTAIL.n446 VTAIL.n401 5.04292
R705 VTAIL.n434 VTAIL.n407 5.04292
R706 VTAIL.n368 VTAIL.n323 5.04292
R707 VTAIL.n356 VTAIL.n329 5.04292
R708 VTAIL.n290 VTAIL.n245 5.04292
R709 VTAIL.n278 VTAIL.n251 5.04292
R710 VTAIL.n572 VTAIL.n571 4.38563
R711 VTAIL.n26 VTAIL.n25 4.38563
R712 VTAIL.n104 VTAIL.n103 4.38563
R713 VTAIL.n182 VTAIL.n181 4.38563
R714 VTAIL.n495 VTAIL.n494 4.38563
R715 VTAIL.n417 VTAIL.n416 4.38563
R716 VTAIL.n339 VTAIL.n338 4.38563
R717 VTAIL.n261 VTAIL.n260 4.38563
R718 VTAIL.n586 VTAIL.n585 4.26717
R719 VTAIL.n602 VTAIL.n554 4.26717
R720 VTAIL.n40 VTAIL.n39 4.26717
R721 VTAIL.n56 VTAIL.n8 4.26717
R722 VTAIL.n118 VTAIL.n117 4.26717
R723 VTAIL.n134 VTAIL.n86 4.26717
R724 VTAIL.n196 VTAIL.n195 4.26717
R725 VTAIL.n212 VTAIL.n164 4.26717
R726 VTAIL.n525 VTAIL.n477 4.26717
R727 VTAIL.n509 VTAIL.n508 4.26717
R728 VTAIL.n447 VTAIL.n399 4.26717
R729 VTAIL.n431 VTAIL.n430 4.26717
R730 VTAIL.n369 VTAIL.n321 4.26717
R731 VTAIL.n353 VTAIL.n352 4.26717
R732 VTAIL.n291 VTAIL.n243 4.26717
R733 VTAIL.n275 VTAIL.n274 4.26717
R734 VTAIL.n582 VTAIL.n564 3.49141
R735 VTAIL.n606 VTAIL.n605 3.49141
R736 VTAIL.n36 VTAIL.n18 3.49141
R737 VTAIL.n60 VTAIL.n59 3.49141
R738 VTAIL.n114 VTAIL.n96 3.49141
R739 VTAIL.n138 VTAIL.n137 3.49141
R740 VTAIL.n192 VTAIL.n174 3.49141
R741 VTAIL.n216 VTAIL.n215 3.49141
R742 VTAIL.n529 VTAIL.n528 3.49141
R743 VTAIL.n505 VTAIL.n487 3.49141
R744 VTAIL.n451 VTAIL.n450 3.49141
R745 VTAIL.n427 VTAIL.n409 3.49141
R746 VTAIL.n373 VTAIL.n372 3.49141
R747 VTAIL.n349 VTAIL.n331 3.49141
R748 VTAIL.n295 VTAIL.n294 3.49141
R749 VTAIL.n271 VTAIL.n253 3.49141
R750 VTAIL.n581 VTAIL.n566 2.71565
R751 VTAIL.n609 VTAIL.n552 2.71565
R752 VTAIL.n35 VTAIL.n20 2.71565
R753 VTAIL.n63 VTAIL.n6 2.71565
R754 VTAIL.n113 VTAIL.n98 2.71565
R755 VTAIL.n141 VTAIL.n84 2.71565
R756 VTAIL.n191 VTAIL.n176 2.71565
R757 VTAIL.n219 VTAIL.n162 2.71565
R758 VTAIL.n532 VTAIL.n475 2.71565
R759 VTAIL.n504 VTAIL.n489 2.71565
R760 VTAIL.n454 VTAIL.n397 2.71565
R761 VTAIL.n426 VTAIL.n411 2.71565
R762 VTAIL.n376 VTAIL.n319 2.71565
R763 VTAIL.n348 VTAIL.n333 2.71565
R764 VTAIL.n298 VTAIL.n241 2.71565
R765 VTAIL.n270 VTAIL.n255 2.71565
R766 VTAIL.n389 VTAIL.n311 2.01774
R767 VTAIL.n545 VTAIL.n467 2.01774
R768 VTAIL.n233 VTAIL.n155 2.01774
R769 VTAIL.n578 VTAIL.n577 1.93989
R770 VTAIL.n610 VTAIL.n550 1.93989
R771 VTAIL.n32 VTAIL.n31 1.93989
R772 VTAIL.n64 VTAIL.n4 1.93989
R773 VTAIL.n110 VTAIL.n109 1.93989
R774 VTAIL.n142 VTAIL.n82 1.93989
R775 VTAIL.n188 VTAIL.n187 1.93989
R776 VTAIL.n220 VTAIL.n160 1.93989
R777 VTAIL.n533 VTAIL.n473 1.93989
R778 VTAIL.n501 VTAIL.n500 1.93989
R779 VTAIL.n455 VTAIL.n395 1.93989
R780 VTAIL.n423 VTAIL.n422 1.93989
R781 VTAIL.n377 VTAIL.n317 1.93989
R782 VTAIL.n345 VTAIL.n344 1.93989
R783 VTAIL.n299 VTAIL.n239 1.93989
R784 VTAIL.n267 VTAIL.n266 1.93989
R785 VTAIL.n574 VTAIL.n568 1.16414
R786 VTAIL.n615 VTAIL.n613 1.16414
R787 VTAIL.n622 VTAIL.n546 1.16414
R788 VTAIL.n28 VTAIL.n22 1.16414
R789 VTAIL.n69 VTAIL.n67 1.16414
R790 VTAIL.n76 VTAIL.n0 1.16414
R791 VTAIL.n106 VTAIL.n100 1.16414
R792 VTAIL.n147 VTAIL.n145 1.16414
R793 VTAIL.n154 VTAIL.n78 1.16414
R794 VTAIL.n184 VTAIL.n178 1.16414
R795 VTAIL.n225 VTAIL.n223 1.16414
R796 VTAIL.n232 VTAIL.n156 1.16414
R797 VTAIL.n544 VTAIL.n468 1.16414
R798 VTAIL.n537 VTAIL.n536 1.16414
R799 VTAIL.n497 VTAIL.n491 1.16414
R800 VTAIL.n466 VTAIL.n390 1.16414
R801 VTAIL.n459 VTAIL.n458 1.16414
R802 VTAIL.n419 VTAIL.n413 1.16414
R803 VTAIL.n388 VTAIL.n312 1.16414
R804 VTAIL.n381 VTAIL.n380 1.16414
R805 VTAIL.n341 VTAIL.n335 1.16414
R806 VTAIL.n310 VTAIL.n234 1.16414
R807 VTAIL.n303 VTAIL.n302 1.16414
R808 VTAIL.n263 VTAIL.n257 1.16414
R809 VTAIL VTAIL.n77 1.06731
R810 VTAIL VTAIL.n623 0.950931
R811 VTAIL.n467 VTAIL.n389 0.470328
R812 VTAIL.n155 VTAIL.n77 0.470328
R813 VTAIL.n573 VTAIL.n570 0.388379
R814 VTAIL.n614 VTAIL.n548 0.388379
R815 VTAIL.n620 VTAIL.n619 0.388379
R816 VTAIL.n27 VTAIL.n24 0.388379
R817 VTAIL.n68 VTAIL.n2 0.388379
R818 VTAIL.n74 VTAIL.n73 0.388379
R819 VTAIL.n105 VTAIL.n102 0.388379
R820 VTAIL.n146 VTAIL.n80 0.388379
R821 VTAIL.n152 VTAIL.n151 0.388379
R822 VTAIL.n183 VTAIL.n180 0.388379
R823 VTAIL.n224 VTAIL.n158 0.388379
R824 VTAIL.n230 VTAIL.n229 0.388379
R825 VTAIL.n542 VTAIL.n541 0.388379
R826 VTAIL.n472 VTAIL.n470 0.388379
R827 VTAIL.n496 VTAIL.n493 0.388379
R828 VTAIL.n464 VTAIL.n463 0.388379
R829 VTAIL.n394 VTAIL.n392 0.388379
R830 VTAIL.n418 VTAIL.n415 0.388379
R831 VTAIL.n386 VTAIL.n385 0.388379
R832 VTAIL.n316 VTAIL.n314 0.388379
R833 VTAIL.n340 VTAIL.n337 0.388379
R834 VTAIL.n308 VTAIL.n307 0.388379
R835 VTAIL.n238 VTAIL.n236 0.388379
R836 VTAIL.n262 VTAIL.n259 0.388379
R837 VTAIL.n572 VTAIL.n567 0.155672
R838 VTAIL.n579 VTAIL.n567 0.155672
R839 VTAIL.n580 VTAIL.n579 0.155672
R840 VTAIL.n580 VTAIL.n563 0.155672
R841 VTAIL.n587 VTAIL.n563 0.155672
R842 VTAIL.n588 VTAIL.n587 0.155672
R843 VTAIL.n588 VTAIL.n559 0.155672
R844 VTAIL.n595 VTAIL.n559 0.155672
R845 VTAIL.n596 VTAIL.n595 0.155672
R846 VTAIL.n596 VTAIL.n555 0.155672
R847 VTAIL.n603 VTAIL.n555 0.155672
R848 VTAIL.n604 VTAIL.n603 0.155672
R849 VTAIL.n604 VTAIL.n551 0.155672
R850 VTAIL.n611 VTAIL.n551 0.155672
R851 VTAIL.n612 VTAIL.n611 0.155672
R852 VTAIL.n612 VTAIL.n547 0.155672
R853 VTAIL.n621 VTAIL.n547 0.155672
R854 VTAIL.n26 VTAIL.n21 0.155672
R855 VTAIL.n33 VTAIL.n21 0.155672
R856 VTAIL.n34 VTAIL.n33 0.155672
R857 VTAIL.n34 VTAIL.n17 0.155672
R858 VTAIL.n41 VTAIL.n17 0.155672
R859 VTAIL.n42 VTAIL.n41 0.155672
R860 VTAIL.n42 VTAIL.n13 0.155672
R861 VTAIL.n49 VTAIL.n13 0.155672
R862 VTAIL.n50 VTAIL.n49 0.155672
R863 VTAIL.n50 VTAIL.n9 0.155672
R864 VTAIL.n57 VTAIL.n9 0.155672
R865 VTAIL.n58 VTAIL.n57 0.155672
R866 VTAIL.n58 VTAIL.n5 0.155672
R867 VTAIL.n65 VTAIL.n5 0.155672
R868 VTAIL.n66 VTAIL.n65 0.155672
R869 VTAIL.n66 VTAIL.n1 0.155672
R870 VTAIL.n75 VTAIL.n1 0.155672
R871 VTAIL.n104 VTAIL.n99 0.155672
R872 VTAIL.n111 VTAIL.n99 0.155672
R873 VTAIL.n112 VTAIL.n111 0.155672
R874 VTAIL.n112 VTAIL.n95 0.155672
R875 VTAIL.n119 VTAIL.n95 0.155672
R876 VTAIL.n120 VTAIL.n119 0.155672
R877 VTAIL.n120 VTAIL.n91 0.155672
R878 VTAIL.n127 VTAIL.n91 0.155672
R879 VTAIL.n128 VTAIL.n127 0.155672
R880 VTAIL.n128 VTAIL.n87 0.155672
R881 VTAIL.n135 VTAIL.n87 0.155672
R882 VTAIL.n136 VTAIL.n135 0.155672
R883 VTAIL.n136 VTAIL.n83 0.155672
R884 VTAIL.n143 VTAIL.n83 0.155672
R885 VTAIL.n144 VTAIL.n143 0.155672
R886 VTAIL.n144 VTAIL.n79 0.155672
R887 VTAIL.n153 VTAIL.n79 0.155672
R888 VTAIL.n182 VTAIL.n177 0.155672
R889 VTAIL.n189 VTAIL.n177 0.155672
R890 VTAIL.n190 VTAIL.n189 0.155672
R891 VTAIL.n190 VTAIL.n173 0.155672
R892 VTAIL.n197 VTAIL.n173 0.155672
R893 VTAIL.n198 VTAIL.n197 0.155672
R894 VTAIL.n198 VTAIL.n169 0.155672
R895 VTAIL.n205 VTAIL.n169 0.155672
R896 VTAIL.n206 VTAIL.n205 0.155672
R897 VTAIL.n206 VTAIL.n165 0.155672
R898 VTAIL.n213 VTAIL.n165 0.155672
R899 VTAIL.n214 VTAIL.n213 0.155672
R900 VTAIL.n214 VTAIL.n161 0.155672
R901 VTAIL.n221 VTAIL.n161 0.155672
R902 VTAIL.n222 VTAIL.n221 0.155672
R903 VTAIL.n222 VTAIL.n157 0.155672
R904 VTAIL.n231 VTAIL.n157 0.155672
R905 VTAIL.n543 VTAIL.n469 0.155672
R906 VTAIL.n535 VTAIL.n469 0.155672
R907 VTAIL.n535 VTAIL.n534 0.155672
R908 VTAIL.n534 VTAIL.n474 0.155672
R909 VTAIL.n527 VTAIL.n474 0.155672
R910 VTAIL.n527 VTAIL.n526 0.155672
R911 VTAIL.n526 VTAIL.n478 0.155672
R912 VTAIL.n519 VTAIL.n478 0.155672
R913 VTAIL.n519 VTAIL.n518 0.155672
R914 VTAIL.n518 VTAIL.n482 0.155672
R915 VTAIL.n511 VTAIL.n482 0.155672
R916 VTAIL.n511 VTAIL.n510 0.155672
R917 VTAIL.n510 VTAIL.n486 0.155672
R918 VTAIL.n503 VTAIL.n486 0.155672
R919 VTAIL.n503 VTAIL.n502 0.155672
R920 VTAIL.n502 VTAIL.n490 0.155672
R921 VTAIL.n495 VTAIL.n490 0.155672
R922 VTAIL.n465 VTAIL.n391 0.155672
R923 VTAIL.n457 VTAIL.n391 0.155672
R924 VTAIL.n457 VTAIL.n456 0.155672
R925 VTAIL.n456 VTAIL.n396 0.155672
R926 VTAIL.n449 VTAIL.n396 0.155672
R927 VTAIL.n449 VTAIL.n448 0.155672
R928 VTAIL.n448 VTAIL.n400 0.155672
R929 VTAIL.n441 VTAIL.n400 0.155672
R930 VTAIL.n441 VTAIL.n440 0.155672
R931 VTAIL.n440 VTAIL.n404 0.155672
R932 VTAIL.n433 VTAIL.n404 0.155672
R933 VTAIL.n433 VTAIL.n432 0.155672
R934 VTAIL.n432 VTAIL.n408 0.155672
R935 VTAIL.n425 VTAIL.n408 0.155672
R936 VTAIL.n425 VTAIL.n424 0.155672
R937 VTAIL.n424 VTAIL.n412 0.155672
R938 VTAIL.n417 VTAIL.n412 0.155672
R939 VTAIL.n387 VTAIL.n313 0.155672
R940 VTAIL.n379 VTAIL.n313 0.155672
R941 VTAIL.n379 VTAIL.n378 0.155672
R942 VTAIL.n378 VTAIL.n318 0.155672
R943 VTAIL.n371 VTAIL.n318 0.155672
R944 VTAIL.n371 VTAIL.n370 0.155672
R945 VTAIL.n370 VTAIL.n322 0.155672
R946 VTAIL.n363 VTAIL.n322 0.155672
R947 VTAIL.n363 VTAIL.n362 0.155672
R948 VTAIL.n362 VTAIL.n326 0.155672
R949 VTAIL.n355 VTAIL.n326 0.155672
R950 VTAIL.n355 VTAIL.n354 0.155672
R951 VTAIL.n354 VTAIL.n330 0.155672
R952 VTAIL.n347 VTAIL.n330 0.155672
R953 VTAIL.n347 VTAIL.n346 0.155672
R954 VTAIL.n346 VTAIL.n334 0.155672
R955 VTAIL.n339 VTAIL.n334 0.155672
R956 VTAIL.n309 VTAIL.n235 0.155672
R957 VTAIL.n301 VTAIL.n235 0.155672
R958 VTAIL.n301 VTAIL.n300 0.155672
R959 VTAIL.n300 VTAIL.n240 0.155672
R960 VTAIL.n293 VTAIL.n240 0.155672
R961 VTAIL.n293 VTAIL.n292 0.155672
R962 VTAIL.n292 VTAIL.n244 0.155672
R963 VTAIL.n285 VTAIL.n244 0.155672
R964 VTAIL.n285 VTAIL.n284 0.155672
R965 VTAIL.n284 VTAIL.n248 0.155672
R966 VTAIL.n277 VTAIL.n248 0.155672
R967 VTAIL.n277 VTAIL.n276 0.155672
R968 VTAIL.n276 VTAIL.n252 0.155672
R969 VTAIL.n269 VTAIL.n252 0.155672
R970 VTAIL.n269 VTAIL.n268 0.155672
R971 VTAIL.n268 VTAIL.n256 0.155672
R972 VTAIL.n261 VTAIL.n256 0.155672
R973 B.n765 B.n764 585
R974 B.n766 B.n765 585
R975 B.n319 B.n108 585
R976 B.n318 B.n317 585
R977 B.n316 B.n315 585
R978 B.n314 B.n313 585
R979 B.n312 B.n311 585
R980 B.n310 B.n309 585
R981 B.n308 B.n307 585
R982 B.n306 B.n305 585
R983 B.n304 B.n303 585
R984 B.n302 B.n301 585
R985 B.n300 B.n299 585
R986 B.n298 B.n297 585
R987 B.n296 B.n295 585
R988 B.n294 B.n293 585
R989 B.n292 B.n291 585
R990 B.n290 B.n289 585
R991 B.n288 B.n287 585
R992 B.n286 B.n285 585
R993 B.n284 B.n283 585
R994 B.n282 B.n281 585
R995 B.n280 B.n279 585
R996 B.n278 B.n277 585
R997 B.n276 B.n275 585
R998 B.n274 B.n273 585
R999 B.n272 B.n271 585
R1000 B.n270 B.n269 585
R1001 B.n268 B.n267 585
R1002 B.n266 B.n265 585
R1003 B.n264 B.n263 585
R1004 B.n262 B.n261 585
R1005 B.n260 B.n259 585
R1006 B.n258 B.n257 585
R1007 B.n256 B.n255 585
R1008 B.n254 B.n253 585
R1009 B.n252 B.n251 585
R1010 B.n250 B.n249 585
R1011 B.n248 B.n247 585
R1012 B.n246 B.n245 585
R1013 B.n244 B.n243 585
R1014 B.n242 B.n241 585
R1015 B.n240 B.n239 585
R1016 B.n238 B.n237 585
R1017 B.n236 B.n235 585
R1018 B.n234 B.n233 585
R1019 B.n232 B.n231 585
R1020 B.n230 B.n229 585
R1021 B.n228 B.n227 585
R1022 B.n225 B.n224 585
R1023 B.n223 B.n222 585
R1024 B.n221 B.n220 585
R1025 B.n219 B.n218 585
R1026 B.n217 B.n216 585
R1027 B.n215 B.n214 585
R1028 B.n213 B.n212 585
R1029 B.n211 B.n210 585
R1030 B.n209 B.n208 585
R1031 B.n207 B.n206 585
R1032 B.n205 B.n204 585
R1033 B.n203 B.n202 585
R1034 B.n201 B.n200 585
R1035 B.n199 B.n198 585
R1036 B.n197 B.n196 585
R1037 B.n195 B.n194 585
R1038 B.n193 B.n192 585
R1039 B.n191 B.n190 585
R1040 B.n189 B.n188 585
R1041 B.n187 B.n186 585
R1042 B.n185 B.n184 585
R1043 B.n183 B.n182 585
R1044 B.n181 B.n180 585
R1045 B.n179 B.n178 585
R1046 B.n177 B.n176 585
R1047 B.n175 B.n174 585
R1048 B.n173 B.n172 585
R1049 B.n171 B.n170 585
R1050 B.n169 B.n168 585
R1051 B.n167 B.n166 585
R1052 B.n165 B.n164 585
R1053 B.n163 B.n162 585
R1054 B.n161 B.n160 585
R1055 B.n159 B.n158 585
R1056 B.n157 B.n156 585
R1057 B.n155 B.n154 585
R1058 B.n153 B.n152 585
R1059 B.n151 B.n150 585
R1060 B.n149 B.n148 585
R1061 B.n147 B.n146 585
R1062 B.n145 B.n144 585
R1063 B.n143 B.n142 585
R1064 B.n141 B.n140 585
R1065 B.n139 B.n138 585
R1066 B.n137 B.n136 585
R1067 B.n135 B.n134 585
R1068 B.n133 B.n132 585
R1069 B.n131 B.n130 585
R1070 B.n129 B.n128 585
R1071 B.n127 B.n126 585
R1072 B.n125 B.n124 585
R1073 B.n123 B.n122 585
R1074 B.n121 B.n120 585
R1075 B.n119 B.n118 585
R1076 B.n117 B.n116 585
R1077 B.n115 B.n114 585
R1078 B.n54 B.n53 585
R1079 B.n763 B.n55 585
R1080 B.n767 B.n55 585
R1081 B.n762 B.n761 585
R1082 B.n761 B.n51 585
R1083 B.n760 B.n50 585
R1084 B.n773 B.n50 585
R1085 B.n759 B.n49 585
R1086 B.n774 B.n49 585
R1087 B.n758 B.n48 585
R1088 B.n775 B.n48 585
R1089 B.n757 B.n756 585
R1090 B.n756 B.n44 585
R1091 B.n755 B.n43 585
R1092 B.n781 B.n43 585
R1093 B.n754 B.n42 585
R1094 B.n782 B.n42 585
R1095 B.n753 B.n41 585
R1096 B.n783 B.n41 585
R1097 B.n752 B.n751 585
R1098 B.n751 B.n37 585
R1099 B.n750 B.n36 585
R1100 B.n789 B.n36 585
R1101 B.n749 B.n35 585
R1102 B.n790 B.n35 585
R1103 B.n748 B.n34 585
R1104 B.n791 B.n34 585
R1105 B.n747 B.n746 585
R1106 B.n746 B.n30 585
R1107 B.n745 B.n29 585
R1108 B.n797 B.n29 585
R1109 B.n744 B.n28 585
R1110 B.n798 B.n28 585
R1111 B.n743 B.n27 585
R1112 B.n799 B.n27 585
R1113 B.n742 B.n741 585
R1114 B.n741 B.n23 585
R1115 B.n740 B.n22 585
R1116 B.n805 B.n22 585
R1117 B.n739 B.n21 585
R1118 B.n806 B.n21 585
R1119 B.n738 B.n20 585
R1120 B.n807 B.n20 585
R1121 B.n737 B.n736 585
R1122 B.n736 B.n16 585
R1123 B.n735 B.n15 585
R1124 B.n813 B.n15 585
R1125 B.n734 B.n14 585
R1126 B.n814 B.n14 585
R1127 B.n733 B.n13 585
R1128 B.n815 B.n13 585
R1129 B.n732 B.n731 585
R1130 B.n731 B.n12 585
R1131 B.n730 B.n729 585
R1132 B.n730 B.n8 585
R1133 B.n728 B.n7 585
R1134 B.n822 B.n7 585
R1135 B.n727 B.n6 585
R1136 B.n823 B.n6 585
R1137 B.n726 B.n5 585
R1138 B.n824 B.n5 585
R1139 B.n725 B.n724 585
R1140 B.n724 B.n4 585
R1141 B.n723 B.n320 585
R1142 B.n723 B.n722 585
R1143 B.n713 B.n321 585
R1144 B.n322 B.n321 585
R1145 B.n715 B.n714 585
R1146 B.n716 B.n715 585
R1147 B.n712 B.n326 585
R1148 B.n330 B.n326 585
R1149 B.n711 B.n710 585
R1150 B.n710 B.n709 585
R1151 B.n328 B.n327 585
R1152 B.n329 B.n328 585
R1153 B.n702 B.n701 585
R1154 B.n703 B.n702 585
R1155 B.n700 B.n335 585
R1156 B.n335 B.n334 585
R1157 B.n699 B.n698 585
R1158 B.n698 B.n697 585
R1159 B.n337 B.n336 585
R1160 B.n338 B.n337 585
R1161 B.n690 B.n689 585
R1162 B.n691 B.n690 585
R1163 B.n688 B.n343 585
R1164 B.n343 B.n342 585
R1165 B.n687 B.n686 585
R1166 B.n686 B.n685 585
R1167 B.n345 B.n344 585
R1168 B.n346 B.n345 585
R1169 B.n678 B.n677 585
R1170 B.n679 B.n678 585
R1171 B.n676 B.n351 585
R1172 B.n351 B.n350 585
R1173 B.n675 B.n674 585
R1174 B.n674 B.n673 585
R1175 B.n353 B.n352 585
R1176 B.n354 B.n353 585
R1177 B.n666 B.n665 585
R1178 B.n667 B.n666 585
R1179 B.n664 B.n359 585
R1180 B.n359 B.n358 585
R1181 B.n663 B.n662 585
R1182 B.n662 B.n661 585
R1183 B.n361 B.n360 585
R1184 B.n362 B.n361 585
R1185 B.n654 B.n653 585
R1186 B.n655 B.n654 585
R1187 B.n652 B.n367 585
R1188 B.n367 B.n366 585
R1189 B.n651 B.n650 585
R1190 B.n650 B.n649 585
R1191 B.n369 B.n368 585
R1192 B.n370 B.n369 585
R1193 B.n642 B.n641 585
R1194 B.n643 B.n642 585
R1195 B.n373 B.n372 585
R1196 B.n433 B.n431 585
R1197 B.n434 B.n430 585
R1198 B.n434 B.n374 585
R1199 B.n437 B.n436 585
R1200 B.n438 B.n429 585
R1201 B.n440 B.n439 585
R1202 B.n442 B.n428 585
R1203 B.n445 B.n444 585
R1204 B.n446 B.n427 585
R1205 B.n448 B.n447 585
R1206 B.n450 B.n426 585
R1207 B.n453 B.n452 585
R1208 B.n454 B.n425 585
R1209 B.n456 B.n455 585
R1210 B.n458 B.n424 585
R1211 B.n461 B.n460 585
R1212 B.n462 B.n423 585
R1213 B.n464 B.n463 585
R1214 B.n466 B.n422 585
R1215 B.n469 B.n468 585
R1216 B.n470 B.n421 585
R1217 B.n472 B.n471 585
R1218 B.n474 B.n420 585
R1219 B.n477 B.n476 585
R1220 B.n478 B.n419 585
R1221 B.n480 B.n479 585
R1222 B.n482 B.n418 585
R1223 B.n485 B.n484 585
R1224 B.n486 B.n417 585
R1225 B.n488 B.n487 585
R1226 B.n490 B.n416 585
R1227 B.n493 B.n492 585
R1228 B.n494 B.n415 585
R1229 B.n496 B.n495 585
R1230 B.n498 B.n414 585
R1231 B.n501 B.n500 585
R1232 B.n502 B.n413 585
R1233 B.n504 B.n503 585
R1234 B.n506 B.n412 585
R1235 B.n509 B.n508 585
R1236 B.n510 B.n411 585
R1237 B.n512 B.n511 585
R1238 B.n514 B.n410 585
R1239 B.n517 B.n516 585
R1240 B.n518 B.n409 585
R1241 B.n520 B.n519 585
R1242 B.n522 B.n408 585
R1243 B.n525 B.n524 585
R1244 B.n527 B.n405 585
R1245 B.n529 B.n528 585
R1246 B.n531 B.n404 585
R1247 B.n534 B.n533 585
R1248 B.n535 B.n403 585
R1249 B.n537 B.n536 585
R1250 B.n539 B.n402 585
R1251 B.n542 B.n541 585
R1252 B.n543 B.n399 585
R1253 B.n546 B.n545 585
R1254 B.n548 B.n398 585
R1255 B.n551 B.n550 585
R1256 B.n552 B.n397 585
R1257 B.n554 B.n553 585
R1258 B.n556 B.n396 585
R1259 B.n559 B.n558 585
R1260 B.n560 B.n395 585
R1261 B.n562 B.n561 585
R1262 B.n564 B.n394 585
R1263 B.n567 B.n566 585
R1264 B.n568 B.n393 585
R1265 B.n570 B.n569 585
R1266 B.n572 B.n392 585
R1267 B.n575 B.n574 585
R1268 B.n576 B.n391 585
R1269 B.n578 B.n577 585
R1270 B.n580 B.n390 585
R1271 B.n583 B.n582 585
R1272 B.n584 B.n389 585
R1273 B.n586 B.n585 585
R1274 B.n588 B.n388 585
R1275 B.n591 B.n590 585
R1276 B.n592 B.n387 585
R1277 B.n594 B.n593 585
R1278 B.n596 B.n386 585
R1279 B.n599 B.n598 585
R1280 B.n600 B.n385 585
R1281 B.n602 B.n601 585
R1282 B.n604 B.n384 585
R1283 B.n607 B.n606 585
R1284 B.n608 B.n383 585
R1285 B.n610 B.n609 585
R1286 B.n612 B.n382 585
R1287 B.n615 B.n614 585
R1288 B.n616 B.n381 585
R1289 B.n618 B.n617 585
R1290 B.n620 B.n380 585
R1291 B.n623 B.n622 585
R1292 B.n624 B.n379 585
R1293 B.n626 B.n625 585
R1294 B.n628 B.n378 585
R1295 B.n631 B.n630 585
R1296 B.n632 B.n377 585
R1297 B.n634 B.n633 585
R1298 B.n636 B.n376 585
R1299 B.n639 B.n638 585
R1300 B.n640 B.n375 585
R1301 B.n645 B.n644 585
R1302 B.n644 B.n643 585
R1303 B.n646 B.n371 585
R1304 B.n371 B.n370 585
R1305 B.n648 B.n647 585
R1306 B.n649 B.n648 585
R1307 B.n365 B.n364 585
R1308 B.n366 B.n365 585
R1309 B.n657 B.n656 585
R1310 B.n656 B.n655 585
R1311 B.n658 B.n363 585
R1312 B.n363 B.n362 585
R1313 B.n660 B.n659 585
R1314 B.n661 B.n660 585
R1315 B.n357 B.n356 585
R1316 B.n358 B.n357 585
R1317 B.n669 B.n668 585
R1318 B.n668 B.n667 585
R1319 B.n670 B.n355 585
R1320 B.n355 B.n354 585
R1321 B.n672 B.n671 585
R1322 B.n673 B.n672 585
R1323 B.n349 B.n348 585
R1324 B.n350 B.n349 585
R1325 B.n681 B.n680 585
R1326 B.n680 B.n679 585
R1327 B.n682 B.n347 585
R1328 B.n347 B.n346 585
R1329 B.n684 B.n683 585
R1330 B.n685 B.n684 585
R1331 B.n341 B.n340 585
R1332 B.n342 B.n341 585
R1333 B.n693 B.n692 585
R1334 B.n692 B.n691 585
R1335 B.n694 B.n339 585
R1336 B.n339 B.n338 585
R1337 B.n696 B.n695 585
R1338 B.n697 B.n696 585
R1339 B.n333 B.n332 585
R1340 B.n334 B.n333 585
R1341 B.n705 B.n704 585
R1342 B.n704 B.n703 585
R1343 B.n706 B.n331 585
R1344 B.n331 B.n329 585
R1345 B.n708 B.n707 585
R1346 B.n709 B.n708 585
R1347 B.n325 B.n324 585
R1348 B.n330 B.n325 585
R1349 B.n718 B.n717 585
R1350 B.n717 B.n716 585
R1351 B.n719 B.n323 585
R1352 B.n323 B.n322 585
R1353 B.n721 B.n720 585
R1354 B.n722 B.n721 585
R1355 B.n3 B.n0 585
R1356 B.n4 B.n3 585
R1357 B.n821 B.n1 585
R1358 B.n822 B.n821 585
R1359 B.n820 B.n819 585
R1360 B.n820 B.n8 585
R1361 B.n818 B.n9 585
R1362 B.n12 B.n9 585
R1363 B.n817 B.n816 585
R1364 B.n816 B.n815 585
R1365 B.n11 B.n10 585
R1366 B.n814 B.n11 585
R1367 B.n812 B.n811 585
R1368 B.n813 B.n812 585
R1369 B.n810 B.n17 585
R1370 B.n17 B.n16 585
R1371 B.n809 B.n808 585
R1372 B.n808 B.n807 585
R1373 B.n19 B.n18 585
R1374 B.n806 B.n19 585
R1375 B.n804 B.n803 585
R1376 B.n805 B.n804 585
R1377 B.n802 B.n24 585
R1378 B.n24 B.n23 585
R1379 B.n801 B.n800 585
R1380 B.n800 B.n799 585
R1381 B.n26 B.n25 585
R1382 B.n798 B.n26 585
R1383 B.n796 B.n795 585
R1384 B.n797 B.n796 585
R1385 B.n794 B.n31 585
R1386 B.n31 B.n30 585
R1387 B.n793 B.n792 585
R1388 B.n792 B.n791 585
R1389 B.n33 B.n32 585
R1390 B.n790 B.n33 585
R1391 B.n788 B.n787 585
R1392 B.n789 B.n788 585
R1393 B.n786 B.n38 585
R1394 B.n38 B.n37 585
R1395 B.n785 B.n784 585
R1396 B.n784 B.n783 585
R1397 B.n40 B.n39 585
R1398 B.n782 B.n40 585
R1399 B.n780 B.n779 585
R1400 B.n781 B.n780 585
R1401 B.n778 B.n45 585
R1402 B.n45 B.n44 585
R1403 B.n777 B.n776 585
R1404 B.n776 B.n775 585
R1405 B.n47 B.n46 585
R1406 B.n774 B.n47 585
R1407 B.n772 B.n771 585
R1408 B.n773 B.n772 585
R1409 B.n770 B.n52 585
R1410 B.n52 B.n51 585
R1411 B.n769 B.n768 585
R1412 B.n768 B.n767 585
R1413 B.n825 B.n824 585
R1414 B.n823 B.n2 585
R1415 B.n768 B.n54 578.989
R1416 B.n765 B.n55 578.989
R1417 B.n642 B.n375 578.989
R1418 B.n644 B.n373 578.989
R1419 B.n111 B.t11 376.601
R1420 B.n109 B.t15 376.601
R1421 B.n400 B.t4 376.601
R1422 B.n406 B.t8 376.601
R1423 B.n109 B.t16 364.661
R1424 B.n400 B.t7 364.661
R1425 B.n111 B.t13 364.661
R1426 B.n406 B.t10 364.661
R1427 B.n110 B.t17 319.279
R1428 B.n401 B.t6 319.279
R1429 B.n112 B.t14 319.279
R1430 B.n407 B.t9 319.279
R1431 B.n766 B.n107 256.663
R1432 B.n766 B.n106 256.663
R1433 B.n766 B.n105 256.663
R1434 B.n766 B.n104 256.663
R1435 B.n766 B.n103 256.663
R1436 B.n766 B.n102 256.663
R1437 B.n766 B.n101 256.663
R1438 B.n766 B.n100 256.663
R1439 B.n766 B.n99 256.663
R1440 B.n766 B.n98 256.663
R1441 B.n766 B.n97 256.663
R1442 B.n766 B.n96 256.663
R1443 B.n766 B.n95 256.663
R1444 B.n766 B.n94 256.663
R1445 B.n766 B.n93 256.663
R1446 B.n766 B.n92 256.663
R1447 B.n766 B.n91 256.663
R1448 B.n766 B.n90 256.663
R1449 B.n766 B.n89 256.663
R1450 B.n766 B.n88 256.663
R1451 B.n766 B.n87 256.663
R1452 B.n766 B.n86 256.663
R1453 B.n766 B.n85 256.663
R1454 B.n766 B.n84 256.663
R1455 B.n766 B.n83 256.663
R1456 B.n766 B.n82 256.663
R1457 B.n766 B.n81 256.663
R1458 B.n766 B.n80 256.663
R1459 B.n766 B.n79 256.663
R1460 B.n766 B.n78 256.663
R1461 B.n766 B.n77 256.663
R1462 B.n766 B.n76 256.663
R1463 B.n766 B.n75 256.663
R1464 B.n766 B.n74 256.663
R1465 B.n766 B.n73 256.663
R1466 B.n766 B.n72 256.663
R1467 B.n766 B.n71 256.663
R1468 B.n766 B.n70 256.663
R1469 B.n766 B.n69 256.663
R1470 B.n766 B.n68 256.663
R1471 B.n766 B.n67 256.663
R1472 B.n766 B.n66 256.663
R1473 B.n766 B.n65 256.663
R1474 B.n766 B.n64 256.663
R1475 B.n766 B.n63 256.663
R1476 B.n766 B.n62 256.663
R1477 B.n766 B.n61 256.663
R1478 B.n766 B.n60 256.663
R1479 B.n766 B.n59 256.663
R1480 B.n766 B.n58 256.663
R1481 B.n766 B.n57 256.663
R1482 B.n766 B.n56 256.663
R1483 B.n432 B.n374 256.663
R1484 B.n435 B.n374 256.663
R1485 B.n441 B.n374 256.663
R1486 B.n443 B.n374 256.663
R1487 B.n449 B.n374 256.663
R1488 B.n451 B.n374 256.663
R1489 B.n457 B.n374 256.663
R1490 B.n459 B.n374 256.663
R1491 B.n465 B.n374 256.663
R1492 B.n467 B.n374 256.663
R1493 B.n473 B.n374 256.663
R1494 B.n475 B.n374 256.663
R1495 B.n481 B.n374 256.663
R1496 B.n483 B.n374 256.663
R1497 B.n489 B.n374 256.663
R1498 B.n491 B.n374 256.663
R1499 B.n497 B.n374 256.663
R1500 B.n499 B.n374 256.663
R1501 B.n505 B.n374 256.663
R1502 B.n507 B.n374 256.663
R1503 B.n513 B.n374 256.663
R1504 B.n515 B.n374 256.663
R1505 B.n521 B.n374 256.663
R1506 B.n523 B.n374 256.663
R1507 B.n530 B.n374 256.663
R1508 B.n532 B.n374 256.663
R1509 B.n538 B.n374 256.663
R1510 B.n540 B.n374 256.663
R1511 B.n547 B.n374 256.663
R1512 B.n549 B.n374 256.663
R1513 B.n555 B.n374 256.663
R1514 B.n557 B.n374 256.663
R1515 B.n563 B.n374 256.663
R1516 B.n565 B.n374 256.663
R1517 B.n571 B.n374 256.663
R1518 B.n573 B.n374 256.663
R1519 B.n579 B.n374 256.663
R1520 B.n581 B.n374 256.663
R1521 B.n587 B.n374 256.663
R1522 B.n589 B.n374 256.663
R1523 B.n595 B.n374 256.663
R1524 B.n597 B.n374 256.663
R1525 B.n603 B.n374 256.663
R1526 B.n605 B.n374 256.663
R1527 B.n611 B.n374 256.663
R1528 B.n613 B.n374 256.663
R1529 B.n619 B.n374 256.663
R1530 B.n621 B.n374 256.663
R1531 B.n627 B.n374 256.663
R1532 B.n629 B.n374 256.663
R1533 B.n635 B.n374 256.663
R1534 B.n637 B.n374 256.663
R1535 B.n827 B.n826 256.663
R1536 B.n116 B.n115 163.367
R1537 B.n120 B.n119 163.367
R1538 B.n124 B.n123 163.367
R1539 B.n128 B.n127 163.367
R1540 B.n132 B.n131 163.367
R1541 B.n136 B.n135 163.367
R1542 B.n140 B.n139 163.367
R1543 B.n144 B.n143 163.367
R1544 B.n148 B.n147 163.367
R1545 B.n152 B.n151 163.367
R1546 B.n156 B.n155 163.367
R1547 B.n160 B.n159 163.367
R1548 B.n164 B.n163 163.367
R1549 B.n168 B.n167 163.367
R1550 B.n172 B.n171 163.367
R1551 B.n176 B.n175 163.367
R1552 B.n180 B.n179 163.367
R1553 B.n184 B.n183 163.367
R1554 B.n188 B.n187 163.367
R1555 B.n192 B.n191 163.367
R1556 B.n196 B.n195 163.367
R1557 B.n200 B.n199 163.367
R1558 B.n204 B.n203 163.367
R1559 B.n208 B.n207 163.367
R1560 B.n212 B.n211 163.367
R1561 B.n216 B.n215 163.367
R1562 B.n220 B.n219 163.367
R1563 B.n224 B.n223 163.367
R1564 B.n229 B.n228 163.367
R1565 B.n233 B.n232 163.367
R1566 B.n237 B.n236 163.367
R1567 B.n241 B.n240 163.367
R1568 B.n245 B.n244 163.367
R1569 B.n249 B.n248 163.367
R1570 B.n253 B.n252 163.367
R1571 B.n257 B.n256 163.367
R1572 B.n261 B.n260 163.367
R1573 B.n265 B.n264 163.367
R1574 B.n269 B.n268 163.367
R1575 B.n273 B.n272 163.367
R1576 B.n277 B.n276 163.367
R1577 B.n281 B.n280 163.367
R1578 B.n285 B.n284 163.367
R1579 B.n289 B.n288 163.367
R1580 B.n293 B.n292 163.367
R1581 B.n297 B.n296 163.367
R1582 B.n301 B.n300 163.367
R1583 B.n305 B.n304 163.367
R1584 B.n309 B.n308 163.367
R1585 B.n313 B.n312 163.367
R1586 B.n317 B.n316 163.367
R1587 B.n765 B.n108 163.367
R1588 B.n642 B.n369 163.367
R1589 B.n650 B.n369 163.367
R1590 B.n650 B.n367 163.367
R1591 B.n654 B.n367 163.367
R1592 B.n654 B.n361 163.367
R1593 B.n662 B.n361 163.367
R1594 B.n662 B.n359 163.367
R1595 B.n666 B.n359 163.367
R1596 B.n666 B.n353 163.367
R1597 B.n674 B.n353 163.367
R1598 B.n674 B.n351 163.367
R1599 B.n678 B.n351 163.367
R1600 B.n678 B.n345 163.367
R1601 B.n686 B.n345 163.367
R1602 B.n686 B.n343 163.367
R1603 B.n690 B.n343 163.367
R1604 B.n690 B.n337 163.367
R1605 B.n698 B.n337 163.367
R1606 B.n698 B.n335 163.367
R1607 B.n702 B.n335 163.367
R1608 B.n702 B.n328 163.367
R1609 B.n710 B.n328 163.367
R1610 B.n710 B.n326 163.367
R1611 B.n715 B.n326 163.367
R1612 B.n715 B.n321 163.367
R1613 B.n723 B.n321 163.367
R1614 B.n724 B.n723 163.367
R1615 B.n724 B.n5 163.367
R1616 B.n6 B.n5 163.367
R1617 B.n7 B.n6 163.367
R1618 B.n730 B.n7 163.367
R1619 B.n731 B.n730 163.367
R1620 B.n731 B.n13 163.367
R1621 B.n14 B.n13 163.367
R1622 B.n15 B.n14 163.367
R1623 B.n736 B.n15 163.367
R1624 B.n736 B.n20 163.367
R1625 B.n21 B.n20 163.367
R1626 B.n22 B.n21 163.367
R1627 B.n741 B.n22 163.367
R1628 B.n741 B.n27 163.367
R1629 B.n28 B.n27 163.367
R1630 B.n29 B.n28 163.367
R1631 B.n746 B.n29 163.367
R1632 B.n746 B.n34 163.367
R1633 B.n35 B.n34 163.367
R1634 B.n36 B.n35 163.367
R1635 B.n751 B.n36 163.367
R1636 B.n751 B.n41 163.367
R1637 B.n42 B.n41 163.367
R1638 B.n43 B.n42 163.367
R1639 B.n756 B.n43 163.367
R1640 B.n756 B.n48 163.367
R1641 B.n49 B.n48 163.367
R1642 B.n50 B.n49 163.367
R1643 B.n761 B.n50 163.367
R1644 B.n761 B.n55 163.367
R1645 B.n434 B.n433 163.367
R1646 B.n436 B.n434 163.367
R1647 B.n440 B.n429 163.367
R1648 B.n444 B.n442 163.367
R1649 B.n448 B.n427 163.367
R1650 B.n452 B.n450 163.367
R1651 B.n456 B.n425 163.367
R1652 B.n460 B.n458 163.367
R1653 B.n464 B.n423 163.367
R1654 B.n468 B.n466 163.367
R1655 B.n472 B.n421 163.367
R1656 B.n476 B.n474 163.367
R1657 B.n480 B.n419 163.367
R1658 B.n484 B.n482 163.367
R1659 B.n488 B.n417 163.367
R1660 B.n492 B.n490 163.367
R1661 B.n496 B.n415 163.367
R1662 B.n500 B.n498 163.367
R1663 B.n504 B.n413 163.367
R1664 B.n508 B.n506 163.367
R1665 B.n512 B.n411 163.367
R1666 B.n516 B.n514 163.367
R1667 B.n520 B.n409 163.367
R1668 B.n524 B.n522 163.367
R1669 B.n529 B.n405 163.367
R1670 B.n533 B.n531 163.367
R1671 B.n537 B.n403 163.367
R1672 B.n541 B.n539 163.367
R1673 B.n546 B.n399 163.367
R1674 B.n550 B.n548 163.367
R1675 B.n554 B.n397 163.367
R1676 B.n558 B.n556 163.367
R1677 B.n562 B.n395 163.367
R1678 B.n566 B.n564 163.367
R1679 B.n570 B.n393 163.367
R1680 B.n574 B.n572 163.367
R1681 B.n578 B.n391 163.367
R1682 B.n582 B.n580 163.367
R1683 B.n586 B.n389 163.367
R1684 B.n590 B.n588 163.367
R1685 B.n594 B.n387 163.367
R1686 B.n598 B.n596 163.367
R1687 B.n602 B.n385 163.367
R1688 B.n606 B.n604 163.367
R1689 B.n610 B.n383 163.367
R1690 B.n614 B.n612 163.367
R1691 B.n618 B.n381 163.367
R1692 B.n622 B.n620 163.367
R1693 B.n626 B.n379 163.367
R1694 B.n630 B.n628 163.367
R1695 B.n634 B.n377 163.367
R1696 B.n638 B.n636 163.367
R1697 B.n644 B.n371 163.367
R1698 B.n648 B.n371 163.367
R1699 B.n648 B.n365 163.367
R1700 B.n656 B.n365 163.367
R1701 B.n656 B.n363 163.367
R1702 B.n660 B.n363 163.367
R1703 B.n660 B.n357 163.367
R1704 B.n668 B.n357 163.367
R1705 B.n668 B.n355 163.367
R1706 B.n672 B.n355 163.367
R1707 B.n672 B.n349 163.367
R1708 B.n680 B.n349 163.367
R1709 B.n680 B.n347 163.367
R1710 B.n684 B.n347 163.367
R1711 B.n684 B.n341 163.367
R1712 B.n692 B.n341 163.367
R1713 B.n692 B.n339 163.367
R1714 B.n696 B.n339 163.367
R1715 B.n696 B.n333 163.367
R1716 B.n704 B.n333 163.367
R1717 B.n704 B.n331 163.367
R1718 B.n708 B.n331 163.367
R1719 B.n708 B.n325 163.367
R1720 B.n717 B.n325 163.367
R1721 B.n717 B.n323 163.367
R1722 B.n721 B.n323 163.367
R1723 B.n721 B.n3 163.367
R1724 B.n825 B.n3 163.367
R1725 B.n821 B.n2 163.367
R1726 B.n821 B.n820 163.367
R1727 B.n820 B.n9 163.367
R1728 B.n816 B.n9 163.367
R1729 B.n816 B.n11 163.367
R1730 B.n812 B.n11 163.367
R1731 B.n812 B.n17 163.367
R1732 B.n808 B.n17 163.367
R1733 B.n808 B.n19 163.367
R1734 B.n804 B.n19 163.367
R1735 B.n804 B.n24 163.367
R1736 B.n800 B.n24 163.367
R1737 B.n800 B.n26 163.367
R1738 B.n796 B.n26 163.367
R1739 B.n796 B.n31 163.367
R1740 B.n792 B.n31 163.367
R1741 B.n792 B.n33 163.367
R1742 B.n788 B.n33 163.367
R1743 B.n788 B.n38 163.367
R1744 B.n784 B.n38 163.367
R1745 B.n784 B.n40 163.367
R1746 B.n780 B.n40 163.367
R1747 B.n780 B.n45 163.367
R1748 B.n776 B.n45 163.367
R1749 B.n776 B.n47 163.367
R1750 B.n772 B.n47 163.367
R1751 B.n772 B.n52 163.367
R1752 B.n768 B.n52 163.367
R1753 B.n643 B.n374 79.8461
R1754 B.n767 B.n766 79.8461
R1755 B.n56 B.n54 71.676
R1756 B.n116 B.n57 71.676
R1757 B.n120 B.n58 71.676
R1758 B.n124 B.n59 71.676
R1759 B.n128 B.n60 71.676
R1760 B.n132 B.n61 71.676
R1761 B.n136 B.n62 71.676
R1762 B.n140 B.n63 71.676
R1763 B.n144 B.n64 71.676
R1764 B.n148 B.n65 71.676
R1765 B.n152 B.n66 71.676
R1766 B.n156 B.n67 71.676
R1767 B.n160 B.n68 71.676
R1768 B.n164 B.n69 71.676
R1769 B.n168 B.n70 71.676
R1770 B.n172 B.n71 71.676
R1771 B.n176 B.n72 71.676
R1772 B.n180 B.n73 71.676
R1773 B.n184 B.n74 71.676
R1774 B.n188 B.n75 71.676
R1775 B.n192 B.n76 71.676
R1776 B.n196 B.n77 71.676
R1777 B.n200 B.n78 71.676
R1778 B.n204 B.n79 71.676
R1779 B.n208 B.n80 71.676
R1780 B.n212 B.n81 71.676
R1781 B.n216 B.n82 71.676
R1782 B.n220 B.n83 71.676
R1783 B.n224 B.n84 71.676
R1784 B.n229 B.n85 71.676
R1785 B.n233 B.n86 71.676
R1786 B.n237 B.n87 71.676
R1787 B.n241 B.n88 71.676
R1788 B.n245 B.n89 71.676
R1789 B.n249 B.n90 71.676
R1790 B.n253 B.n91 71.676
R1791 B.n257 B.n92 71.676
R1792 B.n261 B.n93 71.676
R1793 B.n265 B.n94 71.676
R1794 B.n269 B.n95 71.676
R1795 B.n273 B.n96 71.676
R1796 B.n277 B.n97 71.676
R1797 B.n281 B.n98 71.676
R1798 B.n285 B.n99 71.676
R1799 B.n289 B.n100 71.676
R1800 B.n293 B.n101 71.676
R1801 B.n297 B.n102 71.676
R1802 B.n301 B.n103 71.676
R1803 B.n305 B.n104 71.676
R1804 B.n309 B.n105 71.676
R1805 B.n313 B.n106 71.676
R1806 B.n317 B.n107 71.676
R1807 B.n108 B.n107 71.676
R1808 B.n316 B.n106 71.676
R1809 B.n312 B.n105 71.676
R1810 B.n308 B.n104 71.676
R1811 B.n304 B.n103 71.676
R1812 B.n300 B.n102 71.676
R1813 B.n296 B.n101 71.676
R1814 B.n292 B.n100 71.676
R1815 B.n288 B.n99 71.676
R1816 B.n284 B.n98 71.676
R1817 B.n280 B.n97 71.676
R1818 B.n276 B.n96 71.676
R1819 B.n272 B.n95 71.676
R1820 B.n268 B.n94 71.676
R1821 B.n264 B.n93 71.676
R1822 B.n260 B.n92 71.676
R1823 B.n256 B.n91 71.676
R1824 B.n252 B.n90 71.676
R1825 B.n248 B.n89 71.676
R1826 B.n244 B.n88 71.676
R1827 B.n240 B.n87 71.676
R1828 B.n236 B.n86 71.676
R1829 B.n232 B.n85 71.676
R1830 B.n228 B.n84 71.676
R1831 B.n223 B.n83 71.676
R1832 B.n219 B.n82 71.676
R1833 B.n215 B.n81 71.676
R1834 B.n211 B.n80 71.676
R1835 B.n207 B.n79 71.676
R1836 B.n203 B.n78 71.676
R1837 B.n199 B.n77 71.676
R1838 B.n195 B.n76 71.676
R1839 B.n191 B.n75 71.676
R1840 B.n187 B.n74 71.676
R1841 B.n183 B.n73 71.676
R1842 B.n179 B.n72 71.676
R1843 B.n175 B.n71 71.676
R1844 B.n171 B.n70 71.676
R1845 B.n167 B.n69 71.676
R1846 B.n163 B.n68 71.676
R1847 B.n159 B.n67 71.676
R1848 B.n155 B.n66 71.676
R1849 B.n151 B.n65 71.676
R1850 B.n147 B.n64 71.676
R1851 B.n143 B.n63 71.676
R1852 B.n139 B.n62 71.676
R1853 B.n135 B.n61 71.676
R1854 B.n131 B.n60 71.676
R1855 B.n127 B.n59 71.676
R1856 B.n123 B.n58 71.676
R1857 B.n119 B.n57 71.676
R1858 B.n115 B.n56 71.676
R1859 B.n432 B.n373 71.676
R1860 B.n436 B.n435 71.676
R1861 B.n441 B.n440 71.676
R1862 B.n444 B.n443 71.676
R1863 B.n449 B.n448 71.676
R1864 B.n452 B.n451 71.676
R1865 B.n457 B.n456 71.676
R1866 B.n460 B.n459 71.676
R1867 B.n465 B.n464 71.676
R1868 B.n468 B.n467 71.676
R1869 B.n473 B.n472 71.676
R1870 B.n476 B.n475 71.676
R1871 B.n481 B.n480 71.676
R1872 B.n484 B.n483 71.676
R1873 B.n489 B.n488 71.676
R1874 B.n492 B.n491 71.676
R1875 B.n497 B.n496 71.676
R1876 B.n500 B.n499 71.676
R1877 B.n505 B.n504 71.676
R1878 B.n508 B.n507 71.676
R1879 B.n513 B.n512 71.676
R1880 B.n516 B.n515 71.676
R1881 B.n521 B.n520 71.676
R1882 B.n524 B.n523 71.676
R1883 B.n530 B.n529 71.676
R1884 B.n533 B.n532 71.676
R1885 B.n538 B.n537 71.676
R1886 B.n541 B.n540 71.676
R1887 B.n547 B.n546 71.676
R1888 B.n550 B.n549 71.676
R1889 B.n555 B.n554 71.676
R1890 B.n558 B.n557 71.676
R1891 B.n563 B.n562 71.676
R1892 B.n566 B.n565 71.676
R1893 B.n571 B.n570 71.676
R1894 B.n574 B.n573 71.676
R1895 B.n579 B.n578 71.676
R1896 B.n582 B.n581 71.676
R1897 B.n587 B.n586 71.676
R1898 B.n590 B.n589 71.676
R1899 B.n595 B.n594 71.676
R1900 B.n598 B.n597 71.676
R1901 B.n603 B.n602 71.676
R1902 B.n606 B.n605 71.676
R1903 B.n611 B.n610 71.676
R1904 B.n614 B.n613 71.676
R1905 B.n619 B.n618 71.676
R1906 B.n622 B.n621 71.676
R1907 B.n627 B.n626 71.676
R1908 B.n630 B.n629 71.676
R1909 B.n635 B.n634 71.676
R1910 B.n638 B.n637 71.676
R1911 B.n433 B.n432 71.676
R1912 B.n435 B.n429 71.676
R1913 B.n442 B.n441 71.676
R1914 B.n443 B.n427 71.676
R1915 B.n450 B.n449 71.676
R1916 B.n451 B.n425 71.676
R1917 B.n458 B.n457 71.676
R1918 B.n459 B.n423 71.676
R1919 B.n466 B.n465 71.676
R1920 B.n467 B.n421 71.676
R1921 B.n474 B.n473 71.676
R1922 B.n475 B.n419 71.676
R1923 B.n482 B.n481 71.676
R1924 B.n483 B.n417 71.676
R1925 B.n490 B.n489 71.676
R1926 B.n491 B.n415 71.676
R1927 B.n498 B.n497 71.676
R1928 B.n499 B.n413 71.676
R1929 B.n506 B.n505 71.676
R1930 B.n507 B.n411 71.676
R1931 B.n514 B.n513 71.676
R1932 B.n515 B.n409 71.676
R1933 B.n522 B.n521 71.676
R1934 B.n523 B.n405 71.676
R1935 B.n531 B.n530 71.676
R1936 B.n532 B.n403 71.676
R1937 B.n539 B.n538 71.676
R1938 B.n540 B.n399 71.676
R1939 B.n548 B.n547 71.676
R1940 B.n549 B.n397 71.676
R1941 B.n556 B.n555 71.676
R1942 B.n557 B.n395 71.676
R1943 B.n564 B.n563 71.676
R1944 B.n565 B.n393 71.676
R1945 B.n572 B.n571 71.676
R1946 B.n573 B.n391 71.676
R1947 B.n580 B.n579 71.676
R1948 B.n581 B.n389 71.676
R1949 B.n588 B.n587 71.676
R1950 B.n589 B.n387 71.676
R1951 B.n596 B.n595 71.676
R1952 B.n597 B.n385 71.676
R1953 B.n604 B.n603 71.676
R1954 B.n605 B.n383 71.676
R1955 B.n612 B.n611 71.676
R1956 B.n613 B.n381 71.676
R1957 B.n620 B.n619 71.676
R1958 B.n621 B.n379 71.676
R1959 B.n628 B.n627 71.676
R1960 B.n629 B.n377 71.676
R1961 B.n636 B.n635 71.676
R1962 B.n637 B.n375 71.676
R1963 B.n826 B.n825 71.676
R1964 B.n826 B.n2 71.676
R1965 B.n113 B.n112 59.5399
R1966 B.n226 B.n110 59.5399
R1967 B.n544 B.n401 59.5399
R1968 B.n526 B.n407 59.5399
R1969 B.n112 B.n111 45.3823
R1970 B.n110 B.n109 45.3823
R1971 B.n401 B.n400 45.3823
R1972 B.n407 B.n406 45.3823
R1973 B.n643 B.n370 38.5076
R1974 B.n649 B.n370 38.5076
R1975 B.n649 B.n366 38.5076
R1976 B.n655 B.n366 38.5076
R1977 B.n655 B.n362 38.5076
R1978 B.n661 B.n362 38.5076
R1979 B.n667 B.n358 38.5076
R1980 B.n667 B.n354 38.5076
R1981 B.n673 B.n354 38.5076
R1982 B.n673 B.n350 38.5076
R1983 B.n679 B.n350 38.5076
R1984 B.n679 B.n346 38.5076
R1985 B.n685 B.n346 38.5076
R1986 B.n685 B.n342 38.5076
R1987 B.n691 B.n342 38.5076
R1988 B.n697 B.n338 38.5076
R1989 B.n697 B.n334 38.5076
R1990 B.n703 B.n334 38.5076
R1991 B.n703 B.n329 38.5076
R1992 B.n709 B.n329 38.5076
R1993 B.n709 B.n330 38.5076
R1994 B.n716 B.n322 38.5076
R1995 B.n722 B.n322 38.5076
R1996 B.n722 B.n4 38.5076
R1997 B.n824 B.n4 38.5076
R1998 B.n824 B.n823 38.5076
R1999 B.n823 B.n822 38.5076
R2000 B.n822 B.n8 38.5076
R2001 B.n12 B.n8 38.5076
R2002 B.n815 B.n12 38.5076
R2003 B.n814 B.n813 38.5076
R2004 B.n813 B.n16 38.5076
R2005 B.n807 B.n16 38.5076
R2006 B.n807 B.n806 38.5076
R2007 B.n806 B.n805 38.5076
R2008 B.n805 B.n23 38.5076
R2009 B.n799 B.n798 38.5076
R2010 B.n798 B.n797 38.5076
R2011 B.n797 B.n30 38.5076
R2012 B.n791 B.n30 38.5076
R2013 B.n791 B.n790 38.5076
R2014 B.n790 B.n789 38.5076
R2015 B.n789 B.n37 38.5076
R2016 B.n783 B.n37 38.5076
R2017 B.n783 B.n782 38.5076
R2018 B.n781 B.n44 38.5076
R2019 B.n775 B.n44 38.5076
R2020 B.n775 B.n774 38.5076
R2021 B.n774 B.n773 38.5076
R2022 B.n773 B.n51 38.5076
R2023 B.n767 B.n51 38.5076
R2024 B.n645 B.n372 37.62
R2025 B.n641 B.n640 37.62
R2026 B.n764 B.n763 37.62
R2027 B.n769 B.n53 37.62
R2028 B.n691 B.t1 22.0854
R2029 B.n799 B.t3 22.0854
R2030 B.n716 B.t2 20.9529
R2031 B.n815 B.t0 20.9529
R2032 B.t5 B.n358 19.8203
R2033 B.n782 B.t12 19.8203
R2034 B.n661 B.t5 18.6878
R2035 B.t12 B.n781 18.6878
R2036 B B.n827 18.0485
R2037 B.n330 B.t2 17.5552
R2038 B.t0 B.n814 17.5552
R2039 B.t1 B.n338 16.4226
R2040 B.t3 B.n23 16.4226
R2041 B.n646 B.n645 10.6151
R2042 B.n647 B.n646 10.6151
R2043 B.n647 B.n364 10.6151
R2044 B.n657 B.n364 10.6151
R2045 B.n658 B.n657 10.6151
R2046 B.n659 B.n658 10.6151
R2047 B.n659 B.n356 10.6151
R2048 B.n669 B.n356 10.6151
R2049 B.n670 B.n669 10.6151
R2050 B.n671 B.n670 10.6151
R2051 B.n671 B.n348 10.6151
R2052 B.n681 B.n348 10.6151
R2053 B.n682 B.n681 10.6151
R2054 B.n683 B.n682 10.6151
R2055 B.n683 B.n340 10.6151
R2056 B.n693 B.n340 10.6151
R2057 B.n694 B.n693 10.6151
R2058 B.n695 B.n694 10.6151
R2059 B.n695 B.n332 10.6151
R2060 B.n705 B.n332 10.6151
R2061 B.n706 B.n705 10.6151
R2062 B.n707 B.n706 10.6151
R2063 B.n707 B.n324 10.6151
R2064 B.n718 B.n324 10.6151
R2065 B.n719 B.n718 10.6151
R2066 B.n720 B.n719 10.6151
R2067 B.n720 B.n0 10.6151
R2068 B.n431 B.n372 10.6151
R2069 B.n431 B.n430 10.6151
R2070 B.n437 B.n430 10.6151
R2071 B.n438 B.n437 10.6151
R2072 B.n439 B.n438 10.6151
R2073 B.n439 B.n428 10.6151
R2074 B.n445 B.n428 10.6151
R2075 B.n446 B.n445 10.6151
R2076 B.n447 B.n446 10.6151
R2077 B.n447 B.n426 10.6151
R2078 B.n453 B.n426 10.6151
R2079 B.n454 B.n453 10.6151
R2080 B.n455 B.n454 10.6151
R2081 B.n455 B.n424 10.6151
R2082 B.n461 B.n424 10.6151
R2083 B.n462 B.n461 10.6151
R2084 B.n463 B.n462 10.6151
R2085 B.n463 B.n422 10.6151
R2086 B.n469 B.n422 10.6151
R2087 B.n470 B.n469 10.6151
R2088 B.n471 B.n470 10.6151
R2089 B.n471 B.n420 10.6151
R2090 B.n477 B.n420 10.6151
R2091 B.n478 B.n477 10.6151
R2092 B.n479 B.n478 10.6151
R2093 B.n479 B.n418 10.6151
R2094 B.n485 B.n418 10.6151
R2095 B.n486 B.n485 10.6151
R2096 B.n487 B.n486 10.6151
R2097 B.n487 B.n416 10.6151
R2098 B.n493 B.n416 10.6151
R2099 B.n494 B.n493 10.6151
R2100 B.n495 B.n494 10.6151
R2101 B.n495 B.n414 10.6151
R2102 B.n501 B.n414 10.6151
R2103 B.n502 B.n501 10.6151
R2104 B.n503 B.n502 10.6151
R2105 B.n503 B.n412 10.6151
R2106 B.n509 B.n412 10.6151
R2107 B.n510 B.n509 10.6151
R2108 B.n511 B.n510 10.6151
R2109 B.n511 B.n410 10.6151
R2110 B.n517 B.n410 10.6151
R2111 B.n518 B.n517 10.6151
R2112 B.n519 B.n518 10.6151
R2113 B.n519 B.n408 10.6151
R2114 B.n525 B.n408 10.6151
R2115 B.n528 B.n527 10.6151
R2116 B.n528 B.n404 10.6151
R2117 B.n534 B.n404 10.6151
R2118 B.n535 B.n534 10.6151
R2119 B.n536 B.n535 10.6151
R2120 B.n536 B.n402 10.6151
R2121 B.n542 B.n402 10.6151
R2122 B.n543 B.n542 10.6151
R2123 B.n545 B.n398 10.6151
R2124 B.n551 B.n398 10.6151
R2125 B.n552 B.n551 10.6151
R2126 B.n553 B.n552 10.6151
R2127 B.n553 B.n396 10.6151
R2128 B.n559 B.n396 10.6151
R2129 B.n560 B.n559 10.6151
R2130 B.n561 B.n560 10.6151
R2131 B.n561 B.n394 10.6151
R2132 B.n567 B.n394 10.6151
R2133 B.n568 B.n567 10.6151
R2134 B.n569 B.n568 10.6151
R2135 B.n569 B.n392 10.6151
R2136 B.n575 B.n392 10.6151
R2137 B.n576 B.n575 10.6151
R2138 B.n577 B.n576 10.6151
R2139 B.n577 B.n390 10.6151
R2140 B.n583 B.n390 10.6151
R2141 B.n584 B.n583 10.6151
R2142 B.n585 B.n584 10.6151
R2143 B.n585 B.n388 10.6151
R2144 B.n591 B.n388 10.6151
R2145 B.n592 B.n591 10.6151
R2146 B.n593 B.n592 10.6151
R2147 B.n593 B.n386 10.6151
R2148 B.n599 B.n386 10.6151
R2149 B.n600 B.n599 10.6151
R2150 B.n601 B.n600 10.6151
R2151 B.n601 B.n384 10.6151
R2152 B.n607 B.n384 10.6151
R2153 B.n608 B.n607 10.6151
R2154 B.n609 B.n608 10.6151
R2155 B.n609 B.n382 10.6151
R2156 B.n615 B.n382 10.6151
R2157 B.n616 B.n615 10.6151
R2158 B.n617 B.n616 10.6151
R2159 B.n617 B.n380 10.6151
R2160 B.n623 B.n380 10.6151
R2161 B.n624 B.n623 10.6151
R2162 B.n625 B.n624 10.6151
R2163 B.n625 B.n378 10.6151
R2164 B.n631 B.n378 10.6151
R2165 B.n632 B.n631 10.6151
R2166 B.n633 B.n632 10.6151
R2167 B.n633 B.n376 10.6151
R2168 B.n639 B.n376 10.6151
R2169 B.n640 B.n639 10.6151
R2170 B.n641 B.n368 10.6151
R2171 B.n651 B.n368 10.6151
R2172 B.n652 B.n651 10.6151
R2173 B.n653 B.n652 10.6151
R2174 B.n653 B.n360 10.6151
R2175 B.n663 B.n360 10.6151
R2176 B.n664 B.n663 10.6151
R2177 B.n665 B.n664 10.6151
R2178 B.n665 B.n352 10.6151
R2179 B.n675 B.n352 10.6151
R2180 B.n676 B.n675 10.6151
R2181 B.n677 B.n676 10.6151
R2182 B.n677 B.n344 10.6151
R2183 B.n687 B.n344 10.6151
R2184 B.n688 B.n687 10.6151
R2185 B.n689 B.n688 10.6151
R2186 B.n689 B.n336 10.6151
R2187 B.n699 B.n336 10.6151
R2188 B.n700 B.n699 10.6151
R2189 B.n701 B.n700 10.6151
R2190 B.n701 B.n327 10.6151
R2191 B.n711 B.n327 10.6151
R2192 B.n712 B.n711 10.6151
R2193 B.n714 B.n712 10.6151
R2194 B.n714 B.n713 10.6151
R2195 B.n713 B.n320 10.6151
R2196 B.n725 B.n320 10.6151
R2197 B.n726 B.n725 10.6151
R2198 B.n727 B.n726 10.6151
R2199 B.n728 B.n727 10.6151
R2200 B.n729 B.n728 10.6151
R2201 B.n732 B.n729 10.6151
R2202 B.n733 B.n732 10.6151
R2203 B.n734 B.n733 10.6151
R2204 B.n735 B.n734 10.6151
R2205 B.n737 B.n735 10.6151
R2206 B.n738 B.n737 10.6151
R2207 B.n739 B.n738 10.6151
R2208 B.n740 B.n739 10.6151
R2209 B.n742 B.n740 10.6151
R2210 B.n743 B.n742 10.6151
R2211 B.n744 B.n743 10.6151
R2212 B.n745 B.n744 10.6151
R2213 B.n747 B.n745 10.6151
R2214 B.n748 B.n747 10.6151
R2215 B.n749 B.n748 10.6151
R2216 B.n750 B.n749 10.6151
R2217 B.n752 B.n750 10.6151
R2218 B.n753 B.n752 10.6151
R2219 B.n754 B.n753 10.6151
R2220 B.n755 B.n754 10.6151
R2221 B.n757 B.n755 10.6151
R2222 B.n758 B.n757 10.6151
R2223 B.n759 B.n758 10.6151
R2224 B.n760 B.n759 10.6151
R2225 B.n762 B.n760 10.6151
R2226 B.n763 B.n762 10.6151
R2227 B.n819 B.n1 10.6151
R2228 B.n819 B.n818 10.6151
R2229 B.n818 B.n817 10.6151
R2230 B.n817 B.n10 10.6151
R2231 B.n811 B.n10 10.6151
R2232 B.n811 B.n810 10.6151
R2233 B.n810 B.n809 10.6151
R2234 B.n809 B.n18 10.6151
R2235 B.n803 B.n18 10.6151
R2236 B.n803 B.n802 10.6151
R2237 B.n802 B.n801 10.6151
R2238 B.n801 B.n25 10.6151
R2239 B.n795 B.n25 10.6151
R2240 B.n795 B.n794 10.6151
R2241 B.n794 B.n793 10.6151
R2242 B.n793 B.n32 10.6151
R2243 B.n787 B.n32 10.6151
R2244 B.n787 B.n786 10.6151
R2245 B.n786 B.n785 10.6151
R2246 B.n785 B.n39 10.6151
R2247 B.n779 B.n39 10.6151
R2248 B.n779 B.n778 10.6151
R2249 B.n778 B.n777 10.6151
R2250 B.n777 B.n46 10.6151
R2251 B.n771 B.n46 10.6151
R2252 B.n771 B.n770 10.6151
R2253 B.n770 B.n769 10.6151
R2254 B.n114 B.n53 10.6151
R2255 B.n117 B.n114 10.6151
R2256 B.n118 B.n117 10.6151
R2257 B.n121 B.n118 10.6151
R2258 B.n122 B.n121 10.6151
R2259 B.n125 B.n122 10.6151
R2260 B.n126 B.n125 10.6151
R2261 B.n129 B.n126 10.6151
R2262 B.n130 B.n129 10.6151
R2263 B.n133 B.n130 10.6151
R2264 B.n134 B.n133 10.6151
R2265 B.n137 B.n134 10.6151
R2266 B.n138 B.n137 10.6151
R2267 B.n141 B.n138 10.6151
R2268 B.n142 B.n141 10.6151
R2269 B.n145 B.n142 10.6151
R2270 B.n146 B.n145 10.6151
R2271 B.n149 B.n146 10.6151
R2272 B.n150 B.n149 10.6151
R2273 B.n153 B.n150 10.6151
R2274 B.n154 B.n153 10.6151
R2275 B.n157 B.n154 10.6151
R2276 B.n158 B.n157 10.6151
R2277 B.n161 B.n158 10.6151
R2278 B.n162 B.n161 10.6151
R2279 B.n165 B.n162 10.6151
R2280 B.n166 B.n165 10.6151
R2281 B.n169 B.n166 10.6151
R2282 B.n170 B.n169 10.6151
R2283 B.n173 B.n170 10.6151
R2284 B.n174 B.n173 10.6151
R2285 B.n177 B.n174 10.6151
R2286 B.n178 B.n177 10.6151
R2287 B.n181 B.n178 10.6151
R2288 B.n182 B.n181 10.6151
R2289 B.n185 B.n182 10.6151
R2290 B.n186 B.n185 10.6151
R2291 B.n189 B.n186 10.6151
R2292 B.n190 B.n189 10.6151
R2293 B.n193 B.n190 10.6151
R2294 B.n194 B.n193 10.6151
R2295 B.n197 B.n194 10.6151
R2296 B.n198 B.n197 10.6151
R2297 B.n201 B.n198 10.6151
R2298 B.n202 B.n201 10.6151
R2299 B.n205 B.n202 10.6151
R2300 B.n206 B.n205 10.6151
R2301 B.n210 B.n209 10.6151
R2302 B.n213 B.n210 10.6151
R2303 B.n214 B.n213 10.6151
R2304 B.n217 B.n214 10.6151
R2305 B.n218 B.n217 10.6151
R2306 B.n221 B.n218 10.6151
R2307 B.n222 B.n221 10.6151
R2308 B.n225 B.n222 10.6151
R2309 B.n230 B.n227 10.6151
R2310 B.n231 B.n230 10.6151
R2311 B.n234 B.n231 10.6151
R2312 B.n235 B.n234 10.6151
R2313 B.n238 B.n235 10.6151
R2314 B.n239 B.n238 10.6151
R2315 B.n242 B.n239 10.6151
R2316 B.n243 B.n242 10.6151
R2317 B.n246 B.n243 10.6151
R2318 B.n247 B.n246 10.6151
R2319 B.n250 B.n247 10.6151
R2320 B.n251 B.n250 10.6151
R2321 B.n254 B.n251 10.6151
R2322 B.n255 B.n254 10.6151
R2323 B.n258 B.n255 10.6151
R2324 B.n259 B.n258 10.6151
R2325 B.n262 B.n259 10.6151
R2326 B.n263 B.n262 10.6151
R2327 B.n266 B.n263 10.6151
R2328 B.n267 B.n266 10.6151
R2329 B.n270 B.n267 10.6151
R2330 B.n271 B.n270 10.6151
R2331 B.n274 B.n271 10.6151
R2332 B.n275 B.n274 10.6151
R2333 B.n278 B.n275 10.6151
R2334 B.n279 B.n278 10.6151
R2335 B.n282 B.n279 10.6151
R2336 B.n283 B.n282 10.6151
R2337 B.n286 B.n283 10.6151
R2338 B.n287 B.n286 10.6151
R2339 B.n290 B.n287 10.6151
R2340 B.n291 B.n290 10.6151
R2341 B.n294 B.n291 10.6151
R2342 B.n295 B.n294 10.6151
R2343 B.n298 B.n295 10.6151
R2344 B.n299 B.n298 10.6151
R2345 B.n302 B.n299 10.6151
R2346 B.n303 B.n302 10.6151
R2347 B.n306 B.n303 10.6151
R2348 B.n307 B.n306 10.6151
R2349 B.n310 B.n307 10.6151
R2350 B.n311 B.n310 10.6151
R2351 B.n314 B.n311 10.6151
R2352 B.n315 B.n314 10.6151
R2353 B.n318 B.n315 10.6151
R2354 B.n319 B.n318 10.6151
R2355 B.n764 B.n319 10.6151
R2356 B.n827 B.n0 8.11757
R2357 B.n827 B.n1 8.11757
R2358 B.n527 B.n526 6.5566
R2359 B.n544 B.n543 6.5566
R2360 B.n209 B.n113 6.5566
R2361 B.n226 B.n225 6.5566
R2362 B.n526 B.n525 4.05904
R2363 B.n545 B.n544 4.05904
R2364 B.n206 B.n113 4.05904
R2365 B.n227 B.n226 4.05904
R2366 VN.n0 VN.t3 205.304
R2367 VN.n1 VN.t1 205.304
R2368 VN.n0 VN.t2 204.77
R2369 VN.n1 VN.t0 204.77
R2370 VN VN.n1 53.6227
R2371 VN VN.n0 7.24008
R2372 VDD2.n2 VDD2.n0 107.439
R2373 VDD2.n2 VDD2.n1 65.4748
R2374 VDD2.n1 VDD2.t3 1.39979
R2375 VDD2.n1 VDD2.t2 1.39979
R2376 VDD2.n0 VDD2.t0 1.39979
R2377 VDD2.n0 VDD2.t1 1.39979
R2378 VDD2 VDD2.n2 0.0586897
C0 VDD1 VP 5.46734f
C1 VDD2 VP 0.356888f
C2 VTAIL VP 5.01681f
C3 VN VDD1 0.148593f
C4 VN VDD2 5.25963f
C5 VN VTAIL 5.00271f
C6 VDD1 VDD2 0.886292f
C7 VTAIL VDD1 5.94815f
C8 VTAIL VDD2 5.99841f
C9 VN VP 6.1649f
C10 VDD2 B 3.601592f
C11 VDD1 B 7.76679f
C12 VTAIL B 11.007162f
C13 VN B 9.831599f
C14 VP B 7.833314f
C15 VDD2.t0 B 0.298443f
C16 VDD2.t1 B 0.298443f
C17 VDD2.n0 B 3.38284f
C18 VDD2.t3 B 0.298443f
C19 VDD2.t2 B 0.298443f
C20 VDD2.n1 B 2.69489f
C21 VDD2.n2 B 3.84926f
C22 VN.t3 B 2.45745f
C23 VN.t2 B 2.45494f
C24 VN.n0 B 1.66779f
C25 VN.t1 B 2.45745f
C26 VN.t0 B 2.45494f
C27 VN.n1 B 3.10231f
C28 VTAIL.n0 B 0.021878f
C29 VTAIL.n1 B 0.01564f
C30 VTAIL.n2 B 0.008652f
C31 VTAIL.n3 B 0.019865f
C32 VTAIL.n4 B 0.008899f
C33 VTAIL.n5 B 0.01564f
C34 VTAIL.n6 B 0.008404f
C35 VTAIL.n7 B 0.019865f
C36 VTAIL.n8 B 0.008899f
C37 VTAIL.n9 B 0.01564f
C38 VTAIL.n10 B 0.008404f
C39 VTAIL.n11 B 0.019865f
C40 VTAIL.n12 B 0.008899f
C41 VTAIL.n13 B 0.01564f
C42 VTAIL.n14 B 0.008404f
C43 VTAIL.n15 B 0.019865f
C44 VTAIL.n16 B 0.008899f
C45 VTAIL.n17 B 0.01564f
C46 VTAIL.n18 B 0.008404f
C47 VTAIL.n19 B 0.019865f
C48 VTAIL.n20 B 0.008899f
C49 VTAIL.n21 B 0.01564f
C50 VTAIL.n22 B 0.008404f
C51 VTAIL.n23 B 0.014899f
C52 VTAIL.n24 B 0.011735f
C53 VTAIL.t0 B 0.032709f
C54 VTAIL.n25 B 0.098676f
C55 VTAIL.n26 B 0.956651f
C56 VTAIL.n27 B 0.008404f
C57 VTAIL.n28 B 0.008899f
C58 VTAIL.n29 B 0.019865f
C59 VTAIL.n30 B 0.019865f
C60 VTAIL.n31 B 0.008899f
C61 VTAIL.n32 B 0.008404f
C62 VTAIL.n33 B 0.01564f
C63 VTAIL.n34 B 0.01564f
C64 VTAIL.n35 B 0.008404f
C65 VTAIL.n36 B 0.008899f
C66 VTAIL.n37 B 0.019865f
C67 VTAIL.n38 B 0.019865f
C68 VTAIL.n39 B 0.008899f
C69 VTAIL.n40 B 0.008404f
C70 VTAIL.n41 B 0.01564f
C71 VTAIL.n42 B 0.01564f
C72 VTAIL.n43 B 0.008404f
C73 VTAIL.n44 B 0.008899f
C74 VTAIL.n45 B 0.019865f
C75 VTAIL.n46 B 0.019865f
C76 VTAIL.n47 B 0.008899f
C77 VTAIL.n48 B 0.008404f
C78 VTAIL.n49 B 0.01564f
C79 VTAIL.n50 B 0.01564f
C80 VTAIL.n51 B 0.008404f
C81 VTAIL.n52 B 0.008899f
C82 VTAIL.n53 B 0.019865f
C83 VTAIL.n54 B 0.019865f
C84 VTAIL.n55 B 0.008899f
C85 VTAIL.n56 B 0.008404f
C86 VTAIL.n57 B 0.01564f
C87 VTAIL.n58 B 0.01564f
C88 VTAIL.n59 B 0.008404f
C89 VTAIL.n60 B 0.008899f
C90 VTAIL.n61 B 0.019865f
C91 VTAIL.n62 B 0.019865f
C92 VTAIL.n63 B 0.008899f
C93 VTAIL.n64 B 0.008404f
C94 VTAIL.n65 B 0.01564f
C95 VTAIL.n66 B 0.01564f
C96 VTAIL.n67 B 0.008404f
C97 VTAIL.n68 B 0.008404f
C98 VTAIL.n69 B 0.008899f
C99 VTAIL.n70 B 0.019865f
C100 VTAIL.n71 B 0.019865f
C101 VTAIL.n72 B 0.042818f
C102 VTAIL.n73 B 0.008652f
C103 VTAIL.n74 B 0.008404f
C104 VTAIL.n75 B 0.041066f
C105 VTAIL.n76 B 0.024082f
C106 VTAIL.n77 B 0.093581f
C107 VTAIL.n78 B 0.021878f
C108 VTAIL.n79 B 0.01564f
C109 VTAIL.n80 B 0.008652f
C110 VTAIL.n81 B 0.019865f
C111 VTAIL.n82 B 0.008899f
C112 VTAIL.n83 B 0.01564f
C113 VTAIL.n84 B 0.008404f
C114 VTAIL.n85 B 0.019865f
C115 VTAIL.n86 B 0.008899f
C116 VTAIL.n87 B 0.01564f
C117 VTAIL.n88 B 0.008404f
C118 VTAIL.n89 B 0.019865f
C119 VTAIL.n90 B 0.008899f
C120 VTAIL.n91 B 0.01564f
C121 VTAIL.n92 B 0.008404f
C122 VTAIL.n93 B 0.019865f
C123 VTAIL.n94 B 0.008899f
C124 VTAIL.n95 B 0.01564f
C125 VTAIL.n96 B 0.008404f
C126 VTAIL.n97 B 0.019865f
C127 VTAIL.n98 B 0.008899f
C128 VTAIL.n99 B 0.01564f
C129 VTAIL.n100 B 0.008404f
C130 VTAIL.n101 B 0.014899f
C131 VTAIL.n102 B 0.011735f
C132 VTAIL.t3 B 0.032709f
C133 VTAIL.n103 B 0.098676f
C134 VTAIL.n104 B 0.956651f
C135 VTAIL.n105 B 0.008404f
C136 VTAIL.n106 B 0.008899f
C137 VTAIL.n107 B 0.019865f
C138 VTAIL.n108 B 0.019865f
C139 VTAIL.n109 B 0.008899f
C140 VTAIL.n110 B 0.008404f
C141 VTAIL.n111 B 0.01564f
C142 VTAIL.n112 B 0.01564f
C143 VTAIL.n113 B 0.008404f
C144 VTAIL.n114 B 0.008899f
C145 VTAIL.n115 B 0.019865f
C146 VTAIL.n116 B 0.019865f
C147 VTAIL.n117 B 0.008899f
C148 VTAIL.n118 B 0.008404f
C149 VTAIL.n119 B 0.01564f
C150 VTAIL.n120 B 0.01564f
C151 VTAIL.n121 B 0.008404f
C152 VTAIL.n122 B 0.008899f
C153 VTAIL.n123 B 0.019865f
C154 VTAIL.n124 B 0.019865f
C155 VTAIL.n125 B 0.008899f
C156 VTAIL.n126 B 0.008404f
C157 VTAIL.n127 B 0.01564f
C158 VTAIL.n128 B 0.01564f
C159 VTAIL.n129 B 0.008404f
C160 VTAIL.n130 B 0.008899f
C161 VTAIL.n131 B 0.019865f
C162 VTAIL.n132 B 0.019865f
C163 VTAIL.n133 B 0.008899f
C164 VTAIL.n134 B 0.008404f
C165 VTAIL.n135 B 0.01564f
C166 VTAIL.n136 B 0.01564f
C167 VTAIL.n137 B 0.008404f
C168 VTAIL.n138 B 0.008899f
C169 VTAIL.n139 B 0.019865f
C170 VTAIL.n140 B 0.019865f
C171 VTAIL.n141 B 0.008899f
C172 VTAIL.n142 B 0.008404f
C173 VTAIL.n143 B 0.01564f
C174 VTAIL.n144 B 0.01564f
C175 VTAIL.n145 B 0.008404f
C176 VTAIL.n146 B 0.008404f
C177 VTAIL.n147 B 0.008899f
C178 VTAIL.n148 B 0.019865f
C179 VTAIL.n149 B 0.019865f
C180 VTAIL.n150 B 0.042818f
C181 VTAIL.n151 B 0.008652f
C182 VTAIL.n152 B 0.008404f
C183 VTAIL.n153 B 0.041066f
C184 VTAIL.n154 B 0.024082f
C185 VTAIL.n155 B 0.141479f
C186 VTAIL.n156 B 0.021878f
C187 VTAIL.n157 B 0.01564f
C188 VTAIL.n158 B 0.008652f
C189 VTAIL.n159 B 0.019865f
C190 VTAIL.n160 B 0.008899f
C191 VTAIL.n161 B 0.01564f
C192 VTAIL.n162 B 0.008404f
C193 VTAIL.n163 B 0.019865f
C194 VTAIL.n164 B 0.008899f
C195 VTAIL.n165 B 0.01564f
C196 VTAIL.n166 B 0.008404f
C197 VTAIL.n167 B 0.019865f
C198 VTAIL.n168 B 0.008899f
C199 VTAIL.n169 B 0.01564f
C200 VTAIL.n170 B 0.008404f
C201 VTAIL.n171 B 0.019865f
C202 VTAIL.n172 B 0.008899f
C203 VTAIL.n173 B 0.01564f
C204 VTAIL.n174 B 0.008404f
C205 VTAIL.n175 B 0.019865f
C206 VTAIL.n176 B 0.008899f
C207 VTAIL.n177 B 0.01564f
C208 VTAIL.n178 B 0.008404f
C209 VTAIL.n179 B 0.014899f
C210 VTAIL.n180 B 0.011735f
C211 VTAIL.t5 B 0.032709f
C212 VTAIL.n181 B 0.098676f
C213 VTAIL.n182 B 0.956651f
C214 VTAIL.n183 B 0.008404f
C215 VTAIL.n184 B 0.008899f
C216 VTAIL.n185 B 0.019865f
C217 VTAIL.n186 B 0.019865f
C218 VTAIL.n187 B 0.008899f
C219 VTAIL.n188 B 0.008404f
C220 VTAIL.n189 B 0.01564f
C221 VTAIL.n190 B 0.01564f
C222 VTAIL.n191 B 0.008404f
C223 VTAIL.n192 B 0.008899f
C224 VTAIL.n193 B 0.019865f
C225 VTAIL.n194 B 0.019865f
C226 VTAIL.n195 B 0.008899f
C227 VTAIL.n196 B 0.008404f
C228 VTAIL.n197 B 0.01564f
C229 VTAIL.n198 B 0.01564f
C230 VTAIL.n199 B 0.008404f
C231 VTAIL.n200 B 0.008899f
C232 VTAIL.n201 B 0.019865f
C233 VTAIL.n202 B 0.019865f
C234 VTAIL.n203 B 0.008899f
C235 VTAIL.n204 B 0.008404f
C236 VTAIL.n205 B 0.01564f
C237 VTAIL.n206 B 0.01564f
C238 VTAIL.n207 B 0.008404f
C239 VTAIL.n208 B 0.008899f
C240 VTAIL.n209 B 0.019865f
C241 VTAIL.n210 B 0.019865f
C242 VTAIL.n211 B 0.008899f
C243 VTAIL.n212 B 0.008404f
C244 VTAIL.n213 B 0.01564f
C245 VTAIL.n214 B 0.01564f
C246 VTAIL.n215 B 0.008404f
C247 VTAIL.n216 B 0.008899f
C248 VTAIL.n217 B 0.019865f
C249 VTAIL.n218 B 0.019865f
C250 VTAIL.n219 B 0.008899f
C251 VTAIL.n220 B 0.008404f
C252 VTAIL.n221 B 0.01564f
C253 VTAIL.n222 B 0.01564f
C254 VTAIL.n223 B 0.008404f
C255 VTAIL.n224 B 0.008404f
C256 VTAIL.n225 B 0.008899f
C257 VTAIL.n226 B 0.019865f
C258 VTAIL.n227 B 0.019865f
C259 VTAIL.n228 B 0.042818f
C260 VTAIL.n229 B 0.008652f
C261 VTAIL.n230 B 0.008404f
C262 VTAIL.n231 B 0.041066f
C263 VTAIL.n232 B 0.024082f
C264 VTAIL.n233 B 1.04667f
C265 VTAIL.n234 B 0.021878f
C266 VTAIL.n235 B 0.01564f
C267 VTAIL.n236 B 0.008652f
C268 VTAIL.n237 B 0.019865f
C269 VTAIL.n238 B 0.008404f
C270 VTAIL.n239 B 0.008899f
C271 VTAIL.n240 B 0.01564f
C272 VTAIL.n241 B 0.008404f
C273 VTAIL.n242 B 0.019865f
C274 VTAIL.n243 B 0.008899f
C275 VTAIL.n244 B 0.01564f
C276 VTAIL.n245 B 0.008404f
C277 VTAIL.n246 B 0.019865f
C278 VTAIL.n247 B 0.008899f
C279 VTAIL.n248 B 0.01564f
C280 VTAIL.n249 B 0.008404f
C281 VTAIL.n250 B 0.019865f
C282 VTAIL.n251 B 0.008899f
C283 VTAIL.n252 B 0.01564f
C284 VTAIL.n253 B 0.008404f
C285 VTAIL.n254 B 0.019865f
C286 VTAIL.n255 B 0.008899f
C287 VTAIL.n256 B 0.01564f
C288 VTAIL.n257 B 0.008404f
C289 VTAIL.n258 B 0.014899f
C290 VTAIL.n259 B 0.011735f
C291 VTAIL.t1 B 0.032709f
C292 VTAIL.n260 B 0.098676f
C293 VTAIL.n261 B 0.956651f
C294 VTAIL.n262 B 0.008404f
C295 VTAIL.n263 B 0.008899f
C296 VTAIL.n264 B 0.019865f
C297 VTAIL.n265 B 0.019865f
C298 VTAIL.n266 B 0.008899f
C299 VTAIL.n267 B 0.008404f
C300 VTAIL.n268 B 0.01564f
C301 VTAIL.n269 B 0.01564f
C302 VTAIL.n270 B 0.008404f
C303 VTAIL.n271 B 0.008899f
C304 VTAIL.n272 B 0.019865f
C305 VTAIL.n273 B 0.019865f
C306 VTAIL.n274 B 0.008899f
C307 VTAIL.n275 B 0.008404f
C308 VTAIL.n276 B 0.01564f
C309 VTAIL.n277 B 0.01564f
C310 VTAIL.n278 B 0.008404f
C311 VTAIL.n279 B 0.008899f
C312 VTAIL.n280 B 0.019865f
C313 VTAIL.n281 B 0.019865f
C314 VTAIL.n282 B 0.008899f
C315 VTAIL.n283 B 0.008404f
C316 VTAIL.n284 B 0.01564f
C317 VTAIL.n285 B 0.01564f
C318 VTAIL.n286 B 0.008404f
C319 VTAIL.n287 B 0.008899f
C320 VTAIL.n288 B 0.019865f
C321 VTAIL.n289 B 0.019865f
C322 VTAIL.n290 B 0.008899f
C323 VTAIL.n291 B 0.008404f
C324 VTAIL.n292 B 0.01564f
C325 VTAIL.n293 B 0.01564f
C326 VTAIL.n294 B 0.008404f
C327 VTAIL.n295 B 0.008899f
C328 VTAIL.n296 B 0.019865f
C329 VTAIL.n297 B 0.019865f
C330 VTAIL.n298 B 0.008899f
C331 VTAIL.n299 B 0.008404f
C332 VTAIL.n300 B 0.01564f
C333 VTAIL.n301 B 0.01564f
C334 VTAIL.n302 B 0.008404f
C335 VTAIL.n303 B 0.008899f
C336 VTAIL.n304 B 0.019865f
C337 VTAIL.n305 B 0.019865f
C338 VTAIL.n306 B 0.042818f
C339 VTAIL.n307 B 0.008652f
C340 VTAIL.n308 B 0.008404f
C341 VTAIL.n309 B 0.041066f
C342 VTAIL.n310 B 0.024082f
C343 VTAIL.n311 B 1.04667f
C344 VTAIL.n312 B 0.021878f
C345 VTAIL.n313 B 0.01564f
C346 VTAIL.n314 B 0.008652f
C347 VTAIL.n315 B 0.019865f
C348 VTAIL.n316 B 0.008404f
C349 VTAIL.n317 B 0.008899f
C350 VTAIL.n318 B 0.01564f
C351 VTAIL.n319 B 0.008404f
C352 VTAIL.n320 B 0.019865f
C353 VTAIL.n321 B 0.008899f
C354 VTAIL.n322 B 0.01564f
C355 VTAIL.n323 B 0.008404f
C356 VTAIL.n324 B 0.019865f
C357 VTAIL.n325 B 0.008899f
C358 VTAIL.n326 B 0.01564f
C359 VTAIL.n327 B 0.008404f
C360 VTAIL.n328 B 0.019865f
C361 VTAIL.n329 B 0.008899f
C362 VTAIL.n330 B 0.01564f
C363 VTAIL.n331 B 0.008404f
C364 VTAIL.n332 B 0.019865f
C365 VTAIL.n333 B 0.008899f
C366 VTAIL.n334 B 0.01564f
C367 VTAIL.n335 B 0.008404f
C368 VTAIL.n336 B 0.014899f
C369 VTAIL.n337 B 0.011735f
C370 VTAIL.t7 B 0.032709f
C371 VTAIL.n338 B 0.098676f
C372 VTAIL.n339 B 0.956651f
C373 VTAIL.n340 B 0.008404f
C374 VTAIL.n341 B 0.008899f
C375 VTAIL.n342 B 0.019865f
C376 VTAIL.n343 B 0.019865f
C377 VTAIL.n344 B 0.008899f
C378 VTAIL.n345 B 0.008404f
C379 VTAIL.n346 B 0.01564f
C380 VTAIL.n347 B 0.01564f
C381 VTAIL.n348 B 0.008404f
C382 VTAIL.n349 B 0.008899f
C383 VTAIL.n350 B 0.019865f
C384 VTAIL.n351 B 0.019865f
C385 VTAIL.n352 B 0.008899f
C386 VTAIL.n353 B 0.008404f
C387 VTAIL.n354 B 0.01564f
C388 VTAIL.n355 B 0.01564f
C389 VTAIL.n356 B 0.008404f
C390 VTAIL.n357 B 0.008899f
C391 VTAIL.n358 B 0.019865f
C392 VTAIL.n359 B 0.019865f
C393 VTAIL.n360 B 0.008899f
C394 VTAIL.n361 B 0.008404f
C395 VTAIL.n362 B 0.01564f
C396 VTAIL.n363 B 0.01564f
C397 VTAIL.n364 B 0.008404f
C398 VTAIL.n365 B 0.008899f
C399 VTAIL.n366 B 0.019865f
C400 VTAIL.n367 B 0.019865f
C401 VTAIL.n368 B 0.008899f
C402 VTAIL.n369 B 0.008404f
C403 VTAIL.n370 B 0.01564f
C404 VTAIL.n371 B 0.01564f
C405 VTAIL.n372 B 0.008404f
C406 VTAIL.n373 B 0.008899f
C407 VTAIL.n374 B 0.019865f
C408 VTAIL.n375 B 0.019865f
C409 VTAIL.n376 B 0.008899f
C410 VTAIL.n377 B 0.008404f
C411 VTAIL.n378 B 0.01564f
C412 VTAIL.n379 B 0.01564f
C413 VTAIL.n380 B 0.008404f
C414 VTAIL.n381 B 0.008899f
C415 VTAIL.n382 B 0.019865f
C416 VTAIL.n383 B 0.019865f
C417 VTAIL.n384 B 0.042818f
C418 VTAIL.n385 B 0.008652f
C419 VTAIL.n386 B 0.008404f
C420 VTAIL.n387 B 0.041066f
C421 VTAIL.n388 B 0.024082f
C422 VTAIL.n389 B 0.141479f
C423 VTAIL.n390 B 0.021878f
C424 VTAIL.n391 B 0.01564f
C425 VTAIL.n392 B 0.008652f
C426 VTAIL.n393 B 0.019865f
C427 VTAIL.n394 B 0.008404f
C428 VTAIL.n395 B 0.008899f
C429 VTAIL.n396 B 0.01564f
C430 VTAIL.n397 B 0.008404f
C431 VTAIL.n398 B 0.019865f
C432 VTAIL.n399 B 0.008899f
C433 VTAIL.n400 B 0.01564f
C434 VTAIL.n401 B 0.008404f
C435 VTAIL.n402 B 0.019865f
C436 VTAIL.n403 B 0.008899f
C437 VTAIL.n404 B 0.01564f
C438 VTAIL.n405 B 0.008404f
C439 VTAIL.n406 B 0.019865f
C440 VTAIL.n407 B 0.008899f
C441 VTAIL.n408 B 0.01564f
C442 VTAIL.n409 B 0.008404f
C443 VTAIL.n410 B 0.019865f
C444 VTAIL.n411 B 0.008899f
C445 VTAIL.n412 B 0.01564f
C446 VTAIL.n413 B 0.008404f
C447 VTAIL.n414 B 0.014899f
C448 VTAIL.n415 B 0.011735f
C449 VTAIL.t2 B 0.032709f
C450 VTAIL.n416 B 0.098676f
C451 VTAIL.n417 B 0.956651f
C452 VTAIL.n418 B 0.008404f
C453 VTAIL.n419 B 0.008899f
C454 VTAIL.n420 B 0.019865f
C455 VTAIL.n421 B 0.019865f
C456 VTAIL.n422 B 0.008899f
C457 VTAIL.n423 B 0.008404f
C458 VTAIL.n424 B 0.01564f
C459 VTAIL.n425 B 0.01564f
C460 VTAIL.n426 B 0.008404f
C461 VTAIL.n427 B 0.008899f
C462 VTAIL.n428 B 0.019865f
C463 VTAIL.n429 B 0.019865f
C464 VTAIL.n430 B 0.008899f
C465 VTAIL.n431 B 0.008404f
C466 VTAIL.n432 B 0.01564f
C467 VTAIL.n433 B 0.01564f
C468 VTAIL.n434 B 0.008404f
C469 VTAIL.n435 B 0.008899f
C470 VTAIL.n436 B 0.019865f
C471 VTAIL.n437 B 0.019865f
C472 VTAIL.n438 B 0.008899f
C473 VTAIL.n439 B 0.008404f
C474 VTAIL.n440 B 0.01564f
C475 VTAIL.n441 B 0.01564f
C476 VTAIL.n442 B 0.008404f
C477 VTAIL.n443 B 0.008899f
C478 VTAIL.n444 B 0.019865f
C479 VTAIL.n445 B 0.019865f
C480 VTAIL.n446 B 0.008899f
C481 VTAIL.n447 B 0.008404f
C482 VTAIL.n448 B 0.01564f
C483 VTAIL.n449 B 0.01564f
C484 VTAIL.n450 B 0.008404f
C485 VTAIL.n451 B 0.008899f
C486 VTAIL.n452 B 0.019865f
C487 VTAIL.n453 B 0.019865f
C488 VTAIL.n454 B 0.008899f
C489 VTAIL.n455 B 0.008404f
C490 VTAIL.n456 B 0.01564f
C491 VTAIL.n457 B 0.01564f
C492 VTAIL.n458 B 0.008404f
C493 VTAIL.n459 B 0.008899f
C494 VTAIL.n460 B 0.019865f
C495 VTAIL.n461 B 0.019865f
C496 VTAIL.n462 B 0.042818f
C497 VTAIL.n463 B 0.008652f
C498 VTAIL.n464 B 0.008404f
C499 VTAIL.n465 B 0.041066f
C500 VTAIL.n466 B 0.024082f
C501 VTAIL.n467 B 0.141479f
C502 VTAIL.n468 B 0.021878f
C503 VTAIL.n469 B 0.01564f
C504 VTAIL.n470 B 0.008652f
C505 VTAIL.n471 B 0.019865f
C506 VTAIL.n472 B 0.008404f
C507 VTAIL.n473 B 0.008899f
C508 VTAIL.n474 B 0.01564f
C509 VTAIL.n475 B 0.008404f
C510 VTAIL.n476 B 0.019865f
C511 VTAIL.n477 B 0.008899f
C512 VTAIL.n478 B 0.01564f
C513 VTAIL.n479 B 0.008404f
C514 VTAIL.n480 B 0.019865f
C515 VTAIL.n481 B 0.008899f
C516 VTAIL.n482 B 0.01564f
C517 VTAIL.n483 B 0.008404f
C518 VTAIL.n484 B 0.019865f
C519 VTAIL.n485 B 0.008899f
C520 VTAIL.n486 B 0.01564f
C521 VTAIL.n487 B 0.008404f
C522 VTAIL.n488 B 0.019865f
C523 VTAIL.n489 B 0.008899f
C524 VTAIL.n490 B 0.01564f
C525 VTAIL.n491 B 0.008404f
C526 VTAIL.n492 B 0.014899f
C527 VTAIL.n493 B 0.011735f
C528 VTAIL.t4 B 0.032709f
C529 VTAIL.n494 B 0.098676f
C530 VTAIL.n495 B 0.956651f
C531 VTAIL.n496 B 0.008404f
C532 VTAIL.n497 B 0.008899f
C533 VTAIL.n498 B 0.019865f
C534 VTAIL.n499 B 0.019865f
C535 VTAIL.n500 B 0.008899f
C536 VTAIL.n501 B 0.008404f
C537 VTAIL.n502 B 0.01564f
C538 VTAIL.n503 B 0.01564f
C539 VTAIL.n504 B 0.008404f
C540 VTAIL.n505 B 0.008899f
C541 VTAIL.n506 B 0.019865f
C542 VTAIL.n507 B 0.019865f
C543 VTAIL.n508 B 0.008899f
C544 VTAIL.n509 B 0.008404f
C545 VTAIL.n510 B 0.01564f
C546 VTAIL.n511 B 0.01564f
C547 VTAIL.n512 B 0.008404f
C548 VTAIL.n513 B 0.008899f
C549 VTAIL.n514 B 0.019865f
C550 VTAIL.n515 B 0.019865f
C551 VTAIL.n516 B 0.008899f
C552 VTAIL.n517 B 0.008404f
C553 VTAIL.n518 B 0.01564f
C554 VTAIL.n519 B 0.01564f
C555 VTAIL.n520 B 0.008404f
C556 VTAIL.n521 B 0.008899f
C557 VTAIL.n522 B 0.019865f
C558 VTAIL.n523 B 0.019865f
C559 VTAIL.n524 B 0.008899f
C560 VTAIL.n525 B 0.008404f
C561 VTAIL.n526 B 0.01564f
C562 VTAIL.n527 B 0.01564f
C563 VTAIL.n528 B 0.008404f
C564 VTAIL.n529 B 0.008899f
C565 VTAIL.n530 B 0.019865f
C566 VTAIL.n531 B 0.019865f
C567 VTAIL.n532 B 0.008899f
C568 VTAIL.n533 B 0.008404f
C569 VTAIL.n534 B 0.01564f
C570 VTAIL.n535 B 0.01564f
C571 VTAIL.n536 B 0.008404f
C572 VTAIL.n537 B 0.008899f
C573 VTAIL.n538 B 0.019865f
C574 VTAIL.n539 B 0.019865f
C575 VTAIL.n540 B 0.042818f
C576 VTAIL.n541 B 0.008652f
C577 VTAIL.n542 B 0.008404f
C578 VTAIL.n543 B 0.041066f
C579 VTAIL.n544 B 0.024082f
C580 VTAIL.n545 B 1.04667f
C581 VTAIL.n546 B 0.021878f
C582 VTAIL.n547 B 0.01564f
C583 VTAIL.n548 B 0.008652f
C584 VTAIL.n549 B 0.019865f
C585 VTAIL.n550 B 0.008899f
C586 VTAIL.n551 B 0.01564f
C587 VTAIL.n552 B 0.008404f
C588 VTAIL.n553 B 0.019865f
C589 VTAIL.n554 B 0.008899f
C590 VTAIL.n555 B 0.01564f
C591 VTAIL.n556 B 0.008404f
C592 VTAIL.n557 B 0.019865f
C593 VTAIL.n558 B 0.008899f
C594 VTAIL.n559 B 0.01564f
C595 VTAIL.n560 B 0.008404f
C596 VTAIL.n561 B 0.019865f
C597 VTAIL.n562 B 0.008899f
C598 VTAIL.n563 B 0.01564f
C599 VTAIL.n564 B 0.008404f
C600 VTAIL.n565 B 0.019865f
C601 VTAIL.n566 B 0.008899f
C602 VTAIL.n567 B 0.01564f
C603 VTAIL.n568 B 0.008404f
C604 VTAIL.n569 B 0.014899f
C605 VTAIL.n570 B 0.011735f
C606 VTAIL.t6 B 0.032709f
C607 VTAIL.n571 B 0.098676f
C608 VTAIL.n572 B 0.956651f
C609 VTAIL.n573 B 0.008404f
C610 VTAIL.n574 B 0.008899f
C611 VTAIL.n575 B 0.019865f
C612 VTAIL.n576 B 0.019865f
C613 VTAIL.n577 B 0.008899f
C614 VTAIL.n578 B 0.008404f
C615 VTAIL.n579 B 0.01564f
C616 VTAIL.n580 B 0.01564f
C617 VTAIL.n581 B 0.008404f
C618 VTAIL.n582 B 0.008899f
C619 VTAIL.n583 B 0.019865f
C620 VTAIL.n584 B 0.019865f
C621 VTAIL.n585 B 0.008899f
C622 VTAIL.n586 B 0.008404f
C623 VTAIL.n587 B 0.01564f
C624 VTAIL.n588 B 0.01564f
C625 VTAIL.n589 B 0.008404f
C626 VTAIL.n590 B 0.008899f
C627 VTAIL.n591 B 0.019865f
C628 VTAIL.n592 B 0.019865f
C629 VTAIL.n593 B 0.008899f
C630 VTAIL.n594 B 0.008404f
C631 VTAIL.n595 B 0.01564f
C632 VTAIL.n596 B 0.01564f
C633 VTAIL.n597 B 0.008404f
C634 VTAIL.n598 B 0.008899f
C635 VTAIL.n599 B 0.019865f
C636 VTAIL.n600 B 0.019865f
C637 VTAIL.n601 B 0.008899f
C638 VTAIL.n602 B 0.008404f
C639 VTAIL.n603 B 0.01564f
C640 VTAIL.n604 B 0.01564f
C641 VTAIL.n605 B 0.008404f
C642 VTAIL.n606 B 0.008899f
C643 VTAIL.n607 B 0.019865f
C644 VTAIL.n608 B 0.019865f
C645 VTAIL.n609 B 0.008899f
C646 VTAIL.n610 B 0.008404f
C647 VTAIL.n611 B 0.01564f
C648 VTAIL.n612 B 0.01564f
C649 VTAIL.n613 B 0.008404f
C650 VTAIL.n614 B 0.008404f
C651 VTAIL.n615 B 0.008899f
C652 VTAIL.n616 B 0.019865f
C653 VTAIL.n617 B 0.019865f
C654 VTAIL.n618 B 0.042818f
C655 VTAIL.n619 B 0.008652f
C656 VTAIL.n620 B 0.008404f
C657 VTAIL.n621 B 0.041066f
C658 VTAIL.n622 B 0.024082f
C659 VTAIL.n623 B 0.992905f
C660 VDD1.t3 B 0.29848f
C661 VDD1.t1 B 0.29848f
C662 VDD1.n0 B 2.69558f
C663 VDD1.t2 B 0.29848f
C664 VDD1.t0 B 0.29848f
C665 VDD1.n1 B 3.40941f
C666 VP.n0 B 0.039358f
C667 VP.t2 B 2.32342f
C668 VP.n1 B 0.04358f
C669 VP.t1 B 2.49094f
C670 VP.t3 B 2.49348f
C671 VP.n2 B 3.13255f
C672 VP.n3 B 1.70945f
C673 VP.t0 B 2.32342f
C674 VP.n4 B 0.913964f
C675 VP.n5 B 0.051243f
C676 VP.n6 B 0.039358f
C677 VP.n7 B 0.029853f
C678 VP.n8 B 0.029853f
C679 VP.n9 B 0.04358f
C680 VP.n10 B 0.051243f
C681 VP.n11 B 0.913964f
C682 VP.n12 B 0.035613f
.ends

