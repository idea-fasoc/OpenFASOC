* NGSPICE file created from diff_pair_sample_0733.ext - technology: sky130A

.subckt diff_pair_sample_0733 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=5.6238 pd=29.62 as=5.6238 ps=29.62 w=14.42 l=0.75
X1 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.6238 pd=29.62 as=5.6238 ps=29.62 w=14.42 l=0.75
X2 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=5.6238 pd=29.62 as=0 ps=0 w=14.42 l=0.75
X3 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=5.6238 pd=29.62 as=0 ps=0 w=14.42 l=0.75
X4 VDD1.t0 VP.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=5.6238 pd=29.62 as=5.6238 ps=29.62 w=14.42 l=0.75
X5 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=5.6238 pd=29.62 as=0 ps=0 w=14.42 l=0.75
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=5.6238 pd=29.62 as=0 ps=0 w=14.42 l=0.75
X7 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.6238 pd=29.62 as=5.6238 ps=29.62 w=14.42 l=0.75
R0 VP.n0 VP.t1 718.639
R1 VP.n0 VP.t0 677.04
R2 VP VP.n0 0.0516364
R3 VTAIL.n1 VTAIL.t1 48.3753
R4 VTAIL.n3 VTAIL.t0 48.3752
R5 VTAIL.n0 VTAIL.t3 48.3752
R6 VTAIL.n2 VTAIL.t2 48.3752
R7 VTAIL.n1 VTAIL.n0 26.6772
R8 VTAIL.n3 VTAIL.n2 25.7462
R9 VTAIL.n2 VTAIL.n1 0.935845
R10 VTAIL VTAIL.n0 0.761276
R11 VTAIL VTAIL.n3 0.175069
R12 VDD1 VDD1.t1 103.781
R13 VDD1 VDD1.t0 65.3449
R14 B.n56 B.t9 665.755
R15 B.n62 B.t13 665.755
R16 B.n149 B.t6 665.755
R17 B.n141 B.t2 665.755
R18 B.n451 B.n89 585
R19 B.n89 B.n30 585
R20 B.n453 B.n452 585
R21 B.n455 B.n88 585
R22 B.n458 B.n457 585
R23 B.n459 B.n87 585
R24 B.n461 B.n460 585
R25 B.n463 B.n86 585
R26 B.n466 B.n465 585
R27 B.n467 B.n85 585
R28 B.n469 B.n468 585
R29 B.n471 B.n84 585
R30 B.n474 B.n473 585
R31 B.n475 B.n83 585
R32 B.n477 B.n476 585
R33 B.n479 B.n82 585
R34 B.n482 B.n481 585
R35 B.n483 B.n81 585
R36 B.n485 B.n484 585
R37 B.n487 B.n80 585
R38 B.n490 B.n489 585
R39 B.n491 B.n79 585
R40 B.n493 B.n492 585
R41 B.n495 B.n78 585
R42 B.n498 B.n497 585
R43 B.n499 B.n77 585
R44 B.n501 B.n500 585
R45 B.n503 B.n76 585
R46 B.n506 B.n505 585
R47 B.n507 B.n75 585
R48 B.n509 B.n508 585
R49 B.n511 B.n74 585
R50 B.n514 B.n513 585
R51 B.n515 B.n73 585
R52 B.n517 B.n516 585
R53 B.n519 B.n72 585
R54 B.n522 B.n521 585
R55 B.n523 B.n71 585
R56 B.n525 B.n524 585
R57 B.n527 B.n70 585
R58 B.n530 B.n529 585
R59 B.n531 B.n69 585
R60 B.n533 B.n532 585
R61 B.n535 B.n68 585
R62 B.n538 B.n537 585
R63 B.n539 B.n67 585
R64 B.n541 B.n540 585
R65 B.n543 B.n66 585
R66 B.n545 B.n544 585
R67 B.n547 B.n546 585
R68 B.n550 B.n549 585
R69 B.n551 B.n61 585
R70 B.n553 B.n552 585
R71 B.n555 B.n60 585
R72 B.n558 B.n557 585
R73 B.n559 B.n59 585
R74 B.n561 B.n560 585
R75 B.n563 B.n58 585
R76 B.n566 B.n565 585
R77 B.n568 B.n55 585
R78 B.n570 B.n569 585
R79 B.n572 B.n54 585
R80 B.n575 B.n574 585
R81 B.n576 B.n53 585
R82 B.n578 B.n577 585
R83 B.n580 B.n52 585
R84 B.n583 B.n582 585
R85 B.n584 B.n51 585
R86 B.n586 B.n585 585
R87 B.n588 B.n50 585
R88 B.n591 B.n590 585
R89 B.n592 B.n49 585
R90 B.n594 B.n593 585
R91 B.n596 B.n48 585
R92 B.n599 B.n598 585
R93 B.n600 B.n47 585
R94 B.n602 B.n601 585
R95 B.n604 B.n46 585
R96 B.n607 B.n606 585
R97 B.n608 B.n45 585
R98 B.n610 B.n609 585
R99 B.n612 B.n44 585
R100 B.n615 B.n614 585
R101 B.n616 B.n43 585
R102 B.n618 B.n617 585
R103 B.n620 B.n42 585
R104 B.n623 B.n622 585
R105 B.n624 B.n41 585
R106 B.n626 B.n625 585
R107 B.n628 B.n40 585
R108 B.n631 B.n630 585
R109 B.n632 B.n39 585
R110 B.n634 B.n633 585
R111 B.n636 B.n38 585
R112 B.n639 B.n638 585
R113 B.n640 B.n37 585
R114 B.n642 B.n641 585
R115 B.n644 B.n36 585
R116 B.n647 B.n646 585
R117 B.n648 B.n35 585
R118 B.n650 B.n649 585
R119 B.n652 B.n34 585
R120 B.n655 B.n654 585
R121 B.n656 B.n33 585
R122 B.n658 B.n657 585
R123 B.n660 B.n32 585
R124 B.n663 B.n662 585
R125 B.n664 B.n31 585
R126 B.n450 B.n29 585
R127 B.n667 B.n29 585
R128 B.n449 B.n28 585
R129 B.n668 B.n28 585
R130 B.n448 B.n27 585
R131 B.n669 B.n27 585
R132 B.n447 B.n446 585
R133 B.n446 B.n23 585
R134 B.n445 B.n22 585
R135 B.n675 B.n22 585
R136 B.n444 B.n21 585
R137 B.n676 B.n21 585
R138 B.n443 B.n20 585
R139 B.n677 B.n20 585
R140 B.n442 B.n441 585
R141 B.n441 B.n16 585
R142 B.n440 B.n15 585
R143 B.n683 B.n15 585
R144 B.n439 B.n14 585
R145 B.n684 B.n14 585
R146 B.n438 B.n13 585
R147 B.n685 B.n13 585
R148 B.n437 B.n436 585
R149 B.n436 B.n12 585
R150 B.n435 B.n434 585
R151 B.n435 B.n8 585
R152 B.n433 B.n7 585
R153 B.n692 B.n7 585
R154 B.n432 B.n6 585
R155 B.n693 B.n6 585
R156 B.n431 B.n5 585
R157 B.n694 B.n5 585
R158 B.n430 B.n429 585
R159 B.n429 B.n4 585
R160 B.n428 B.n90 585
R161 B.n428 B.n427 585
R162 B.n417 B.n91 585
R163 B.n420 B.n91 585
R164 B.n419 B.n418 585
R165 B.n421 B.n419 585
R166 B.n416 B.n96 585
R167 B.n96 B.n95 585
R168 B.n415 B.n414 585
R169 B.n414 B.n413 585
R170 B.n98 B.n97 585
R171 B.n99 B.n98 585
R172 B.n406 B.n405 585
R173 B.n407 B.n406 585
R174 B.n404 B.n104 585
R175 B.n104 B.n103 585
R176 B.n403 B.n402 585
R177 B.n402 B.n401 585
R178 B.n106 B.n105 585
R179 B.n107 B.n106 585
R180 B.n394 B.n393 585
R181 B.n395 B.n394 585
R182 B.n392 B.n112 585
R183 B.n112 B.n111 585
R184 B.n391 B.n390 585
R185 B.n390 B.n389 585
R186 B.n386 B.n116 585
R187 B.n385 B.n384 585
R188 B.n382 B.n117 585
R189 B.n382 B.n115 585
R190 B.n381 B.n380 585
R191 B.n379 B.n378 585
R192 B.n377 B.n119 585
R193 B.n375 B.n374 585
R194 B.n373 B.n120 585
R195 B.n372 B.n371 585
R196 B.n369 B.n121 585
R197 B.n367 B.n366 585
R198 B.n365 B.n122 585
R199 B.n364 B.n363 585
R200 B.n361 B.n123 585
R201 B.n359 B.n358 585
R202 B.n357 B.n124 585
R203 B.n356 B.n355 585
R204 B.n353 B.n125 585
R205 B.n351 B.n350 585
R206 B.n349 B.n126 585
R207 B.n348 B.n347 585
R208 B.n345 B.n127 585
R209 B.n343 B.n342 585
R210 B.n341 B.n128 585
R211 B.n340 B.n339 585
R212 B.n337 B.n129 585
R213 B.n335 B.n334 585
R214 B.n333 B.n130 585
R215 B.n332 B.n331 585
R216 B.n329 B.n131 585
R217 B.n327 B.n326 585
R218 B.n325 B.n132 585
R219 B.n324 B.n323 585
R220 B.n321 B.n133 585
R221 B.n319 B.n318 585
R222 B.n317 B.n134 585
R223 B.n316 B.n315 585
R224 B.n313 B.n135 585
R225 B.n311 B.n310 585
R226 B.n309 B.n136 585
R227 B.n308 B.n307 585
R228 B.n305 B.n137 585
R229 B.n303 B.n302 585
R230 B.n301 B.n138 585
R231 B.n300 B.n299 585
R232 B.n297 B.n139 585
R233 B.n295 B.n294 585
R234 B.n293 B.n140 585
R235 B.n292 B.n291 585
R236 B.n289 B.n288 585
R237 B.n287 B.n286 585
R238 B.n285 B.n145 585
R239 B.n283 B.n282 585
R240 B.n281 B.n146 585
R241 B.n280 B.n279 585
R242 B.n277 B.n147 585
R243 B.n275 B.n274 585
R244 B.n273 B.n148 585
R245 B.n271 B.n270 585
R246 B.n268 B.n151 585
R247 B.n266 B.n265 585
R248 B.n264 B.n152 585
R249 B.n263 B.n262 585
R250 B.n260 B.n153 585
R251 B.n258 B.n257 585
R252 B.n256 B.n154 585
R253 B.n255 B.n254 585
R254 B.n252 B.n155 585
R255 B.n250 B.n249 585
R256 B.n248 B.n156 585
R257 B.n247 B.n246 585
R258 B.n244 B.n157 585
R259 B.n242 B.n241 585
R260 B.n240 B.n158 585
R261 B.n239 B.n238 585
R262 B.n236 B.n159 585
R263 B.n234 B.n233 585
R264 B.n232 B.n160 585
R265 B.n231 B.n230 585
R266 B.n228 B.n161 585
R267 B.n226 B.n225 585
R268 B.n224 B.n162 585
R269 B.n223 B.n222 585
R270 B.n220 B.n163 585
R271 B.n218 B.n217 585
R272 B.n216 B.n164 585
R273 B.n215 B.n214 585
R274 B.n212 B.n165 585
R275 B.n210 B.n209 585
R276 B.n208 B.n166 585
R277 B.n207 B.n206 585
R278 B.n204 B.n167 585
R279 B.n202 B.n201 585
R280 B.n200 B.n168 585
R281 B.n199 B.n198 585
R282 B.n196 B.n169 585
R283 B.n194 B.n193 585
R284 B.n192 B.n170 585
R285 B.n191 B.n190 585
R286 B.n188 B.n171 585
R287 B.n186 B.n185 585
R288 B.n184 B.n172 585
R289 B.n183 B.n182 585
R290 B.n180 B.n173 585
R291 B.n178 B.n177 585
R292 B.n176 B.n175 585
R293 B.n114 B.n113 585
R294 B.n388 B.n387 585
R295 B.n389 B.n388 585
R296 B.n110 B.n109 585
R297 B.n111 B.n110 585
R298 B.n397 B.n396 585
R299 B.n396 B.n395 585
R300 B.n398 B.n108 585
R301 B.n108 B.n107 585
R302 B.n400 B.n399 585
R303 B.n401 B.n400 585
R304 B.n102 B.n101 585
R305 B.n103 B.n102 585
R306 B.n409 B.n408 585
R307 B.n408 B.n407 585
R308 B.n410 B.n100 585
R309 B.n100 B.n99 585
R310 B.n412 B.n411 585
R311 B.n413 B.n412 585
R312 B.n94 B.n93 585
R313 B.n95 B.n94 585
R314 B.n423 B.n422 585
R315 B.n422 B.n421 585
R316 B.n424 B.n92 585
R317 B.n420 B.n92 585
R318 B.n426 B.n425 585
R319 B.n427 B.n426 585
R320 B.n3 B.n0 585
R321 B.n4 B.n3 585
R322 B.n691 B.n1 585
R323 B.n692 B.n691 585
R324 B.n690 B.n689 585
R325 B.n690 B.n8 585
R326 B.n688 B.n9 585
R327 B.n12 B.n9 585
R328 B.n687 B.n686 585
R329 B.n686 B.n685 585
R330 B.n11 B.n10 585
R331 B.n684 B.n11 585
R332 B.n682 B.n681 585
R333 B.n683 B.n682 585
R334 B.n680 B.n17 585
R335 B.n17 B.n16 585
R336 B.n679 B.n678 585
R337 B.n678 B.n677 585
R338 B.n19 B.n18 585
R339 B.n676 B.n19 585
R340 B.n674 B.n673 585
R341 B.n675 B.n674 585
R342 B.n672 B.n24 585
R343 B.n24 B.n23 585
R344 B.n671 B.n670 585
R345 B.n670 B.n669 585
R346 B.n26 B.n25 585
R347 B.n668 B.n26 585
R348 B.n666 B.n665 585
R349 B.n667 B.n666 585
R350 B.n695 B.n694 585
R351 B.n693 B.n2 585
R352 B.n666 B.n31 506.916
R353 B.n89 B.n29 506.916
R354 B.n390 B.n114 506.916
R355 B.n388 B.n116 506.916
R356 B.n454 B.n30 256.663
R357 B.n456 B.n30 256.663
R358 B.n462 B.n30 256.663
R359 B.n464 B.n30 256.663
R360 B.n470 B.n30 256.663
R361 B.n472 B.n30 256.663
R362 B.n478 B.n30 256.663
R363 B.n480 B.n30 256.663
R364 B.n486 B.n30 256.663
R365 B.n488 B.n30 256.663
R366 B.n494 B.n30 256.663
R367 B.n496 B.n30 256.663
R368 B.n502 B.n30 256.663
R369 B.n504 B.n30 256.663
R370 B.n510 B.n30 256.663
R371 B.n512 B.n30 256.663
R372 B.n518 B.n30 256.663
R373 B.n520 B.n30 256.663
R374 B.n526 B.n30 256.663
R375 B.n528 B.n30 256.663
R376 B.n534 B.n30 256.663
R377 B.n536 B.n30 256.663
R378 B.n542 B.n30 256.663
R379 B.n65 B.n30 256.663
R380 B.n548 B.n30 256.663
R381 B.n554 B.n30 256.663
R382 B.n556 B.n30 256.663
R383 B.n562 B.n30 256.663
R384 B.n564 B.n30 256.663
R385 B.n571 B.n30 256.663
R386 B.n573 B.n30 256.663
R387 B.n579 B.n30 256.663
R388 B.n581 B.n30 256.663
R389 B.n587 B.n30 256.663
R390 B.n589 B.n30 256.663
R391 B.n595 B.n30 256.663
R392 B.n597 B.n30 256.663
R393 B.n603 B.n30 256.663
R394 B.n605 B.n30 256.663
R395 B.n611 B.n30 256.663
R396 B.n613 B.n30 256.663
R397 B.n619 B.n30 256.663
R398 B.n621 B.n30 256.663
R399 B.n627 B.n30 256.663
R400 B.n629 B.n30 256.663
R401 B.n635 B.n30 256.663
R402 B.n637 B.n30 256.663
R403 B.n643 B.n30 256.663
R404 B.n645 B.n30 256.663
R405 B.n651 B.n30 256.663
R406 B.n653 B.n30 256.663
R407 B.n659 B.n30 256.663
R408 B.n661 B.n30 256.663
R409 B.n383 B.n115 256.663
R410 B.n118 B.n115 256.663
R411 B.n376 B.n115 256.663
R412 B.n370 B.n115 256.663
R413 B.n368 B.n115 256.663
R414 B.n362 B.n115 256.663
R415 B.n360 B.n115 256.663
R416 B.n354 B.n115 256.663
R417 B.n352 B.n115 256.663
R418 B.n346 B.n115 256.663
R419 B.n344 B.n115 256.663
R420 B.n338 B.n115 256.663
R421 B.n336 B.n115 256.663
R422 B.n330 B.n115 256.663
R423 B.n328 B.n115 256.663
R424 B.n322 B.n115 256.663
R425 B.n320 B.n115 256.663
R426 B.n314 B.n115 256.663
R427 B.n312 B.n115 256.663
R428 B.n306 B.n115 256.663
R429 B.n304 B.n115 256.663
R430 B.n298 B.n115 256.663
R431 B.n296 B.n115 256.663
R432 B.n290 B.n115 256.663
R433 B.n144 B.n115 256.663
R434 B.n284 B.n115 256.663
R435 B.n278 B.n115 256.663
R436 B.n276 B.n115 256.663
R437 B.n269 B.n115 256.663
R438 B.n267 B.n115 256.663
R439 B.n261 B.n115 256.663
R440 B.n259 B.n115 256.663
R441 B.n253 B.n115 256.663
R442 B.n251 B.n115 256.663
R443 B.n245 B.n115 256.663
R444 B.n243 B.n115 256.663
R445 B.n237 B.n115 256.663
R446 B.n235 B.n115 256.663
R447 B.n229 B.n115 256.663
R448 B.n227 B.n115 256.663
R449 B.n221 B.n115 256.663
R450 B.n219 B.n115 256.663
R451 B.n213 B.n115 256.663
R452 B.n211 B.n115 256.663
R453 B.n205 B.n115 256.663
R454 B.n203 B.n115 256.663
R455 B.n197 B.n115 256.663
R456 B.n195 B.n115 256.663
R457 B.n189 B.n115 256.663
R458 B.n187 B.n115 256.663
R459 B.n181 B.n115 256.663
R460 B.n179 B.n115 256.663
R461 B.n174 B.n115 256.663
R462 B.n697 B.n696 256.663
R463 B.n662 B.n660 163.367
R464 B.n658 B.n33 163.367
R465 B.n654 B.n652 163.367
R466 B.n650 B.n35 163.367
R467 B.n646 B.n644 163.367
R468 B.n642 B.n37 163.367
R469 B.n638 B.n636 163.367
R470 B.n634 B.n39 163.367
R471 B.n630 B.n628 163.367
R472 B.n626 B.n41 163.367
R473 B.n622 B.n620 163.367
R474 B.n618 B.n43 163.367
R475 B.n614 B.n612 163.367
R476 B.n610 B.n45 163.367
R477 B.n606 B.n604 163.367
R478 B.n602 B.n47 163.367
R479 B.n598 B.n596 163.367
R480 B.n594 B.n49 163.367
R481 B.n590 B.n588 163.367
R482 B.n586 B.n51 163.367
R483 B.n582 B.n580 163.367
R484 B.n578 B.n53 163.367
R485 B.n574 B.n572 163.367
R486 B.n570 B.n55 163.367
R487 B.n565 B.n563 163.367
R488 B.n561 B.n59 163.367
R489 B.n557 B.n555 163.367
R490 B.n553 B.n61 163.367
R491 B.n549 B.n547 163.367
R492 B.n544 B.n543 163.367
R493 B.n541 B.n67 163.367
R494 B.n537 B.n535 163.367
R495 B.n533 B.n69 163.367
R496 B.n529 B.n527 163.367
R497 B.n525 B.n71 163.367
R498 B.n521 B.n519 163.367
R499 B.n517 B.n73 163.367
R500 B.n513 B.n511 163.367
R501 B.n509 B.n75 163.367
R502 B.n505 B.n503 163.367
R503 B.n501 B.n77 163.367
R504 B.n497 B.n495 163.367
R505 B.n493 B.n79 163.367
R506 B.n489 B.n487 163.367
R507 B.n485 B.n81 163.367
R508 B.n481 B.n479 163.367
R509 B.n477 B.n83 163.367
R510 B.n473 B.n471 163.367
R511 B.n469 B.n85 163.367
R512 B.n465 B.n463 163.367
R513 B.n461 B.n87 163.367
R514 B.n457 B.n455 163.367
R515 B.n453 B.n89 163.367
R516 B.n390 B.n112 163.367
R517 B.n394 B.n112 163.367
R518 B.n394 B.n106 163.367
R519 B.n402 B.n106 163.367
R520 B.n402 B.n104 163.367
R521 B.n406 B.n104 163.367
R522 B.n406 B.n98 163.367
R523 B.n414 B.n98 163.367
R524 B.n414 B.n96 163.367
R525 B.n419 B.n96 163.367
R526 B.n419 B.n91 163.367
R527 B.n428 B.n91 163.367
R528 B.n429 B.n428 163.367
R529 B.n429 B.n5 163.367
R530 B.n6 B.n5 163.367
R531 B.n7 B.n6 163.367
R532 B.n435 B.n7 163.367
R533 B.n436 B.n435 163.367
R534 B.n436 B.n13 163.367
R535 B.n14 B.n13 163.367
R536 B.n15 B.n14 163.367
R537 B.n441 B.n15 163.367
R538 B.n441 B.n20 163.367
R539 B.n21 B.n20 163.367
R540 B.n22 B.n21 163.367
R541 B.n446 B.n22 163.367
R542 B.n446 B.n27 163.367
R543 B.n28 B.n27 163.367
R544 B.n29 B.n28 163.367
R545 B.n384 B.n382 163.367
R546 B.n382 B.n381 163.367
R547 B.n378 B.n377 163.367
R548 B.n375 B.n120 163.367
R549 B.n371 B.n369 163.367
R550 B.n367 B.n122 163.367
R551 B.n363 B.n361 163.367
R552 B.n359 B.n124 163.367
R553 B.n355 B.n353 163.367
R554 B.n351 B.n126 163.367
R555 B.n347 B.n345 163.367
R556 B.n343 B.n128 163.367
R557 B.n339 B.n337 163.367
R558 B.n335 B.n130 163.367
R559 B.n331 B.n329 163.367
R560 B.n327 B.n132 163.367
R561 B.n323 B.n321 163.367
R562 B.n319 B.n134 163.367
R563 B.n315 B.n313 163.367
R564 B.n311 B.n136 163.367
R565 B.n307 B.n305 163.367
R566 B.n303 B.n138 163.367
R567 B.n299 B.n297 163.367
R568 B.n295 B.n140 163.367
R569 B.n291 B.n289 163.367
R570 B.n286 B.n285 163.367
R571 B.n283 B.n146 163.367
R572 B.n279 B.n277 163.367
R573 B.n275 B.n148 163.367
R574 B.n270 B.n268 163.367
R575 B.n266 B.n152 163.367
R576 B.n262 B.n260 163.367
R577 B.n258 B.n154 163.367
R578 B.n254 B.n252 163.367
R579 B.n250 B.n156 163.367
R580 B.n246 B.n244 163.367
R581 B.n242 B.n158 163.367
R582 B.n238 B.n236 163.367
R583 B.n234 B.n160 163.367
R584 B.n230 B.n228 163.367
R585 B.n226 B.n162 163.367
R586 B.n222 B.n220 163.367
R587 B.n218 B.n164 163.367
R588 B.n214 B.n212 163.367
R589 B.n210 B.n166 163.367
R590 B.n206 B.n204 163.367
R591 B.n202 B.n168 163.367
R592 B.n198 B.n196 163.367
R593 B.n194 B.n170 163.367
R594 B.n190 B.n188 163.367
R595 B.n186 B.n172 163.367
R596 B.n182 B.n180 163.367
R597 B.n178 B.n175 163.367
R598 B.n388 B.n110 163.367
R599 B.n396 B.n110 163.367
R600 B.n396 B.n108 163.367
R601 B.n400 B.n108 163.367
R602 B.n400 B.n102 163.367
R603 B.n408 B.n102 163.367
R604 B.n408 B.n100 163.367
R605 B.n412 B.n100 163.367
R606 B.n412 B.n94 163.367
R607 B.n422 B.n94 163.367
R608 B.n422 B.n92 163.367
R609 B.n426 B.n92 163.367
R610 B.n426 B.n3 163.367
R611 B.n695 B.n3 163.367
R612 B.n691 B.n2 163.367
R613 B.n691 B.n690 163.367
R614 B.n690 B.n9 163.367
R615 B.n686 B.n9 163.367
R616 B.n686 B.n11 163.367
R617 B.n682 B.n11 163.367
R618 B.n682 B.n17 163.367
R619 B.n678 B.n17 163.367
R620 B.n678 B.n19 163.367
R621 B.n674 B.n19 163.367
R622 B.n674 B.n24 163.367
R623 B.n670 B.n24 163.367
R624 B.n670 B.n26 163.367
R625 B.n666 B.n26 163.367
R626 B.n62 B.t14 91.1771
R627 B.n149 B.t8 91.1771
R628 B.n56 B.t11 91.1584
R629 B.n141 B.t5 91.1584
R630 B.n661 B.n31 71.676
R631 B.n660 B.n659 71.676
R632 B.n653 B.n33 71.676
R633 B.n652 B.n651 71.676
R634 B.n645 B.n35 71.676
R635 B.n644 B.n643 71.676
R636 B.n637 B.n37 71.676
R637 B.n636 B.n635 71.676
R638 B.n629 B.n39 71.676
R639 B.n628 B.n627 71.676
R640 B.n621 B.n41 71.676
R641 B.n620 B.n619 71.676
R642 B.n613 B.n43 71.676
R643 B.n612 B.n611 71.676
R644 B.n605 B.n45 71.676
R645 B.n604 B.n603 71.676
R646 B.n597 B.n47 71.676
R647 B.n596 B.n595 71.676
R648 B.n589 B.n49 71.676
R649 B.n588 B.n587 71.676
R650 B.n581 B.n51 71.676
R651 B.n580 B.n579 71.676
R652 B.n573 B.n53 71.676
R653 B.n572 B.n571 71.676
R654 B.n564 B.n55 71.676
R655 B.n563 B.n562 71.676
R656 B.n556 B.n59 71.676
R657 B.n555 B.n554 71.676
R658 B.n548 B.n61 71.676
R659 B.n547 B.n65 71.676
R660 B.n543 B.n542 71.676
R661 B.n536 B.n67 71.676
R662 B.n535 B.n534 71.676
R663 B.n528 B.n69 71.676
R664 B.n527 B.n526 71.676
R665 B.n520 B.n71 71.676
R666 B.n519 B.n518 71.676
R667 B.n512 B.n73 71.676
R668 B.n511 B.n510 71.676
R669 B.n504 B.n75 71.676
R670 B.n503 B.n502 71.676
R671 B.n496 B.n77 71.676
R672 B.n495 B.n494 71.676
R673 B.n488 B.n79 71.676
R674 B.n487 B.n486 71.676
R675 B.n480 B.n81 71.676
R676 B.n479 B.n478 71.676
R677 B.n472 B.n83 71.676
R678 B.n471 B.n470 71.676
R679 B.n464 B.n85 71.676
R680 B.n463 B.n462 71.676
R681 B.n456 B.n87 71.676
R682 B.n455 B.n454 71.676
R683 B.n454 B.n453 71.676
R684 B.n457 B.n456 71.676
R685 B.n462 B.n461 71.676
R686 B.n465 B.n464 71.676
R687 B.n470 B.n469 71.676
R688 B.n473 B.n472 71.676
R689 B.n478 B.n477 71.676
R690 B.n481 B.n480 71.676
R691 B.n486 B.n485 71.676
R692 B.n489 B.n488 71.676
R693 B.n494 B.n493 71.676
R694 B.n497 B.n496 71.676
R695 B.n502 B.n501 71.676
R696 B.n505 B.n504 71.676
R697 B.n510 B.n509 71.676
R698 B.n513 B.n512 71.676
R699 B.n518 B.n517 71.676
R700 B.n521 B.n520 71.676
R701 B.n526 B.n525 71.676
R702 B.n529 B.n528 71.676
R703 B.n534 B.n533 71.676
R704 B.n537 B.n536 71.676
R705 B.n542 B.n541 71.676
R706 B.n544 B.n65 71.676
R707 B.n549 B.n548 71.676
R708 B.n554 B.n553 71.676
R709 B.n557 B.n556 71.676
R710 B.n562 B.n561 71.676
R711 B.n565 B.n564 71.676
R712 B.n571 B.n570 71.676
R713 B.n574 B.n573 71.676
R714 B.n579 B.n578 71.676
R715 B.n582 B.n581 71.676
R716 B.n587 B.n586 71.676
R717 B.n590 B.n589 71.676
R718 B.n595 B.n594 71.676
R719 B.n598 B.n597 71.676
R720 B.n603 B.n602 71.676
R721 B.n606 B.n605 71.676
R722 B.n611 B.n610 71.676
R723 B.n614 B.n613 71.676
R724 B.n619 B.n618 71.676
R725 B.n622 B.n621 71.676
R726 B.n627 B.n626 71.676
R727 B.n630 B.n629 71.676
R728 B.n635 B.n634 71.676
R729 B.n638 B.n637 71.676
R730 B.n643 B.n642 71.676
R731 B.n646 B.n645 71.676
R732 B.n651 B.n650 71.676
R733 B.n654 B.n653 71.676
R734 B.n659 B.n658 71.676
R735 B.n662 B.n661 71.676
R736 B.n383 B.n116 71.676
R737 B.n381 B.n118 71.676
R738 B.n377 B.n376 71.676
R739 B.n370 B.n120 71.676
R740 B.n369 B.n368 71.676
R741 B.n362 B.n122 71.676
R742 B.n361 B.n360 71.676
R743 B.n354 B.n124 71.676
R744 B.n353 B.n352 71.676
R745 B.n346 B.n126 71.676
R746 B.n345 B.n344 71.676
R747 B.n338 B.n128 71.676
R748 B.n337 B.n336 71.676
R749 B.n330 B.n130 71.676
R750 B.n329 B.n328 71.676
R751 B.n322 B.n132 71.676
R752 B.n321 B.n320 71.676
R753 B.n314 B.n134 71.676
R754 B.n313 B.n312 71.676
R755 B.n306 B.n136 71.676
R756 B.n305 B.n304 71.676
R757 B.n298 B.n138 71.676
R758 B.n297 B.n296 71.676
R759 B.n290 B.n140 71.676
R760 B.n289 B.n144 71.676
R761 B.n285 B.n284 71.676
R762 B.n278 B.n146 71.676
R763 B.n277 B.n276 71.676
R764 B.n269 B.n148 71.676
R765 B.n268 B.n267 71.676
R766 B.n261 B.n152 71.676
R767 B.n260 B.n259 71.676
R768 B.n253 B.n154 71.676
R769 B.n252 B.n251 71.676
R770 B.n245 B.n156 71.676
R771 B.n244 B.n243 71.676
R772 B.n237 B.n158 71.676
R773 B.n236 B.n235 71.676
R774 B.n229 B.n160 71.676
R775 B.n228 B.n227 71.676
R776 B.n221 B.n162 71.676
R777 B.n220 B.n219 71.676
R778 B.n213 B.n164 71.676
R779 B.n212 B.n211 71.676
R780 B.n205 B.n166 71.676
R781 B.n204 B.n203 71.676
R782 B.n197 B.n168 71.676
R783 B.n196 B.n195 71.676
R784 B.n189 B.n170 71.676
R785 B.n188 B.n187 71.676
R786 B.n181 B.n172 71.676
R787 B.n180 B.n179 71.676
R788 B.n175 B.n174 71.676
R789 B.n384 B.n383 71.676
R790 B.n378 B.n118 71.676
R791 B.n376 B.n375 71.676
R792 B.n371 B.n370 71.676
R793 B.n368 B.n367 71.676
R794 B.n363 B.n362 71.676
R795 B.n360 B.n359 71.676
R796 B.n355 B.n354 71.676
R797 B.n352 B.n351 71.676
R798 B.n347 B.n346 71.676
R799 B.n344 B.n343 71.676
R800 B.n339 B.n338 71.676
R801 B.n336 B.n335 71.676
R802 B.n331 B.n330 71.676
R803 B.n328 B.n327 71.676
R804 B.n323 B.n322 71.676
R805 B.n320 B.n319 71.676
R806 B.n315 B.n314 71.676
R807 B.n312 B.n311 71.676
R808 B.n307 B.n306 71.676
R809 B.n304 B.n303 71.676
R810 B.n299 B.n298 71.676
R811 B.n296 B.n295 71.676
R812 B.n291 B.n290 71.676
R813 B.n286 B.n144 71.676
R814 B.n284 B.n283 71.676
R815 B.n279 B.n278 71.676
R816 B.n276 B.n275 71.676
R817 B.n270 B.n269 71.676
R818 B.n267 B.n266 71.676
R819 B.n262 B.n261 71.676
R820 B.n259 B.n258 71.676
R821 B.n254 B.n253 71.676
R822 B.n251 B.n250 71.676
R823 B.n246 B.n245 71.676
R824 B.n243 B.n242 71.676
R825 B.n238 B.n237 71.676
R826 B.n235 B.n234 71.676
R827 B.n230 B.n229 71.676
R828 B.n227 B.n226 71.676
R829 B.n222 B.n221 71.676
R830 B.n219 B.n218 71.676
R831 B.n214 B.n213 71.676
R832 B.n211 B.n210 71.676
R833 B.n206 B.n205 71.676
R834 B.n203 B.n202 71.676
R835 B.n198 B.n197 71.676
R836 B.n195 B.n194 71.676
R837 B.n190 B.n189 71.676
R838 B.n187 B.n186 71.676
R839 B.n182 B.n181 71.676
R840 B.n179 B.n178 71.676
R841 B.n174 B.n114 71.676
R842 B.n696 B.n695 71.676
R843 B.n696 B.n2 71.676
R844 B.n63 B.t15 70.2316
R845 B.n150 B.t7 70.2316
R846 B.n57 B.t12 70.2129
R847 B.n142 B.t4 70.2129
R848 B.n389 B.n115 67.5125
R849 B.n667 B.n30 67.5125
R850 B.n567 B.n57 59.5399
R851 B.n64 B.n63 59.5399
R852 B.n272 B.n150 59.5399
R853 B.n143 B.n142 59.5399
R854 B.n389 B.n111 37.9412
R855 B.n395 B.n111 37.9412
R856 B.n395 B.n107 37.9412
R857 B.n401 B.n107 37.9412
R858 B.n407 B.n103 37.9412
R859 B.n407 B.n99 37.9412
R860 B.n413 B.n99 37.9412
R861 B.n413 B.n95 37.9412
R862 B.n421 B.n95 37.9412
R863 B.n421 B.n420 37.9412
R864 B.n427 B.n4 37.9412
R865 B.n694 B.n4 37.9412
R866 B.n694 B.n693 37.9412
R867 B.n693 B.n692 37.9412
R868 B.n692 B.n8 37.9412
R869 B.n685 B.n12 37.9412
R870 B.n685 B.n684 37.9412
R871 B.n684 B.n683 37.9412
R872 B.n683 B.n16 37.9412
R873 B.n677 B.n16 37.9412
R874 B.n677 B.n676 37.9412
R875 B.n675 B.n23 37.9412
R876 B.n669 B.n23 37.9412
R877 B.n669 B.n668 37.9412
R878 B.n668 B.n667 37.9412
R879 B.n401 B.t3 35.1514
R880 B.t10 B.n675 35.1514
R881 B.n387 B.n386 32.9371
R882 B.n391 B.n113 32.9371
R883 B.n451 B.n450 32.9371
R884 B.n665 B.n664 32.9371
R885 B.n427 B.t1 26.2242
R886 B.t0 B.n8 26.2242
R887 B.n57 B.n56 20.946
R888 B.n63 B.n62 20.946
R889 B.n150 B.n149 20.946
R890 B.n142 B.n141 20.946
R891 B B.n697 18.0485
R892 B.n420 B.t1 11.7175
R893 B.n12 B.t0 11.7175
R894 B.n387 B.n109 10.6151
R895 B.n397 B.n109 10.6151
R896 B.n398 B.n397 10.6151
R897 B.n399 B.n398 10.6151
R898 B.n399 B.n101 10.6151
R899 B.n409 B.n101 10.6151
R900 B.n410 B.n409 10.6151
R901 B.n411 B.n410 10.6151
R902 B.n411 B.n93 10.6151
R903 B.n423 B.n93 10.6151
R904 B.n424 B.n423 10.6151
R905 B.n425 B.n424 10.6151
R906 B.n425 B.n0 10.6151
R907 B.n386 B.n385 10.6151
R908 B.n385 B.n117 10.6151
R909 B.n380 B.n117 10.6151
R910 B.n380 B.n379 10.6151
R911 B.n379 B.n119 10.6151
R912 B.n374 B.n119 10.6151
R913 B.n374 B.n373 10.6151
R914 B.n373 B.n372 10.6151
R915 B.n372 B.n121 10.6151
R916 B.n366 B.n121 10.6151
R917 B.n366 B.n365 10.6151
R918 B.n365 B.n364 10.6151
R919 B.n364 B.n123 10.6151
R920 B.n358 B.n123 10.6151
R921 B.n358 B.n357 10.6151
R922 B.n357 B.n356 10.6151
R923 B.n356 B.n125 10.6151
R924 B.n350 B.n125 10.6151
R925 B.n350 B.n349 10.6151
R926 B.n349 B.n348 10.6151
R927 B.n348 B.n127 10.6151
R928 B.n342 B.n127 10.6151
R929 B.n342 B.n341 10.6151
R930 B.n341 B.n340 10.6151
R931 B.n340 B.n129 10.6151
R932 B.n334 B.n129 10.6151
R933 B.n334 B.n333 10.6151
R934 B.n333 B.n332 10.6151
R935 B.n332 B.n131 10.6151
R936 B.n326 B.n131 10.6151
R937 B.n326 B.n325 10.6151
R938 B.n325 B.n324 10.6151
R939 B.n324 B.n133 10.6151
R940 B.n318 B.n133 10.6151
R941 B.n318 B.n317 10.6151
R942 B.n317 B.n316 10.6151
R943 B.n316 B.n135 10.6151
R944 B.n310 B.n135 10.6151
R945 B.n310 B.n309 10.6151
R946 B.n309 B.n308 10.6151
R947 B.n308 B.n137 10.6151
R948 B.n302 B.n137 10.6151
R949 B.n302 B.n301 10.6151
R950 B.n301 B.n300 10.6151
R951 B.n300 B.n139 10.6151
R952 B.n294 B.n139 10.6151
R953 B.n294 B.n293 10.6151
R954 B.n293 B.n292 10.6151
R955 B.n288 B.n287 10.6151
R956 B.n287 B.n145 10.6151
R957 B.n282 B.n145 10.6151
R958 B.n282 B.n281 10.6151
R959 B.n281 B.n280 10.6151
R960 B.n280 B.n147 10.6151
R961 B.n274 B.n147 10.6151
R962 B.n274 B.n273 10.6151
R963 B.n271 B.n151 10.6151
R964 B.n265 B.n151 10.6151
R965 B.n265 B.n264 10.6151
R966 B.n264 B.n263 10.6151
R967 B.n263 B.n153 10.6151
R968 B.n257 B.n153 10.6151
R969 B.n257 B.n256 10.6151
R970 B.n256 B.n255 10.6151
R971 B.n255 B.n155 10.6151
R972 B.n249 B.n155 10.6151
R973 B.n249 B.n248 10.6151
R974 B.n248 B.n247 10.6151
R975 B.n247 B.n157 10.6151
R976 B.n241 B.n157 10.6151
R977 B.n241 B.n240 10.6151
R978 B.n240 B.n239 10.6151
R979 B.n239 B.n159 10.6151
R980 B.n233 B.n159 10.6151
R981 B.n233 B.n232 10.6151
R982 B.n232 B.n231 10.6151
R983 B.n231 B.n161 10.6151
R984 B.n225 B.n161 10.6151
R985 B.n225 B.n224 10.6151
R986 B.n224 B.n223 10.6151
R987 B.n223 B.n163 10.6151
R988 B.n217 B.n163 10.6151
R989 B.n217 B.n216 10.6151
R990 B.n216 B.n215 10.6151
R991 B.n215 B.n165 10.6151
R992 B.n209 B.n165 10.6151
R993 B.n209 B.n208 10.6151
R994 B.n208 B.n207 10.6151
R995 B.n207 B.n167 10.6151
R996 B.n201 B.n167 10.6151
R997 B.n201 B.n200 10.6151
R998 B.n200 B.n199 10.6151
R999 B.n199 B.n169 10.6151
R1000 B.n193 B.n169 10.6151
R1001 B.n193 B.n192 10.6151
R1002 B.n192 B.n191 10.6151
R1003 B.n191 B.n171 10.6151
R1004 B.n185 B.n171 10.6151
R1005 B.n185 B.n184 10.6151
R1006 B.n184 B.n183 10.6151
R1007 B.n183 B.n173 10.6151
R1008 B.n177 B.n173 10.6151
R1009 B.n177 B.n176 10.6151
R1010 B.n176 B.n113 10.6151
R1011 B.n392 B.n391 10.6151
R1012 B.n393 B.n392 10.6151
R1013 B.n393 B.n105 10.6151
R1014 B.n403 B.n105 10.6151
R1015 B.n404 B.n403 10.6151
R1016 B.n405 B.n404 10.6151
R1017 B.n405 B.n97 10.6151
R1018 B.n415 B.n97 10.6151
R1019 B.n416 B.n415 10.6151
R1020 B.n418 B.n416 10.6151
R1021 B.n418 B.n417 10.6151
R1022 B.n417 B.n90 10.6151
R1023 B.n430 B.n90 10.6151
R1024 B.n431 B.n430 10.6151
R1025 B.n432 B.n431 10.6151
R1026 B.n433 B.n432 10.6151
R1027 B.n434 B.n433 10.6151
R1028 B.n437 B.n434 10.6151
R1029 B.n438 B.n437 10.6151
R1030 B.n439 B.n438 10.6151
R1031 B.n440 B.n439 10.6151
R1032 B.n442 B.n440 10.6151
R1033 B.n443 B.n442 10.6151
R1034 B.n444 B.n443 10.6151
R1035 B.n445 B.n444 10.6151
R1036 B.n447 B.n445 10.6151
R1037 B.n448 B.n447 10.6151
R1038 B.n449 B.n448 10.6151
R1039 B.n450 B.n449 10.6151
R1040 B.n689 B.n1 10.6151
R1041 B.n689 B.n688 10.6151
R1042 B.n688 B.n687 10.6151
R1043 B.n687 B.n10 10.6151
R1044 B.n681 B.n10 10.6151
R1045 B.n681 B.n680 10.6151
R1046 B.n680 B.n679 10.6151
R1047 B.n679 B.n18 10.6151
R1048 B.n673 B.n18 10.6151
R1049 B.n673 B.n672 10.6151
R1050 B.n672 B.n671 10.6151
R1051 B.n671 B.n25 10.6151
R1052 B.n665 B.n25 10.6151
R1053 B.n664 B.n663 10.6151
R1054 B.n663 B.n32 10.6151
R1055 B.n657 B.n32 10.6151
R1056 B.n657 B.n656 10.6151
R1057 B.n656 B.n655 10.6151
R1058 B.n655 B.n34 10.6151
R1059 B.n649 B.n34 10.6151
R1060 B.n649 B.n648 10.6151
R1061 B.n648 B.n647 10.6151
R1062 B.n647 B.n36 10.6151
R1063 B.n641 B.n36 10.6151
R1064 B.n641 B.n640 10.6151
R1065 B.n640 B.n639 10.6151
R1066 B.n639 B.n38 10.6151
R1067 B.n633 B.n38 10.6151
R1068 B.n633 B.n632 10.6151
R1069 B.n632 B.n631 10.6151
R1070 B.n631 B.n40 10.6151
R1071 B.n625 B.n40 10.6151
R1072 B.n625 B.n624 10.6151
R1073 B.n624 B.n623 10.6151
R1074 B.n623 B.n42 10.6151
R1075 B.n617 B.n42 10.6151
R1076 B.n617 B.n616 10.6151
R1077 B.n616 B.n615 10.6151
R1078 B.n615 B.n44 10.6151
R1079 B.n609 B.n44 10.6151
R1080 B.n609 B.n608 10.6151
R1081 B.n608 B.n607 10.6151
R1082 B.n607 B.n46 10.6151
R1083 B.n601 B.n46 10.6151
R1084 B.n601 B.n600 10.6151
R1085 B.n600 B.n599 10.6151
R1086 B.n599 B.n48 10.6151
R1087 B.n593 B.n48 10.6151
R1088 B.n593 B.n592 10.6151
R1089 B.n592 B.n591 10.6151
R1090 B.n591 B.n50 10.6151
R1091 B.n585 B.n50 10.6151
R1092 B.n585 B.n584 10.6151
R1093 B.n584 B.n583 10.6151
R1094 B.n583 B.n52 10.6151
R1095 B.n577 B.n52 10.6151
R1096 B.n577 B.n576 10.6151
R1097 B.n576 B.n575 10.6151
R1098 B.n575 B.n54 10.6151
R1099 B.n569 B.n54 10.6151
R1100 B.n569 B.n568 10.6151
R1101 B.n566 B.n58 10.6151
R1102 B.n560 B.n58 10.6151
R1103 B.n560 B.n559 10.6151
R1104 B.n559 B.n558 10.6151
R1105 B.n558 B.n60 10.6151
R1106 B.n552 B.n60 10.6151
R1107 B.n552 B.n551 10.6151
R1108 B.n551 B.n550 10.6151
R1109 B.n546 B.n545 10.6151
R1110 B.n545 B.n66 10.6151
R1111 B.n540 B.n66 10.6151
R1112 B.n540 B.n539 10.6151
R1113 B.n539 B.n538 10.6151
R1114 B.n538 B.n68 10.6151
R1115 B.n532 B.n68 10.6151
R1116 B.n532 B.n531 10.6151
R1117 B.n531 B.n530 10.6151
R1118 B.n530 B.n70 10.6151
R1119 B.n524 B.n70 10.6151
R1120 B.n524 B.n523 10.6151
R1121 B.n523 B.n522 10.6151
R1122 B.n522 B.n72 10.6151
R1123 B.n516 B.n72 10.6151
R1124 B.n516 B.n515 10.6151
R1125 B.n515 B.n514 10.6151
R1126 B.n514 B.n74 10.6151
R1127 B.n508 B.n74 10.6151
R1128 B.n508 B.n507 10.6151
R1129 B.n507 B.n506 10.6151
R1130 B.n506 B.n76 10.6151
R1131 B.n500 B.n76 10.6151
R1132 B.n500 B.n499 10.6151
R1133 B.n499 B.n498 10.6151
R1134 B.n498 B.n78 10.6151
R1135 B.n492 B.n78 10.6151
R1136 B.n492 B.n491 10.6151
R1137 B.n491 B.n490 10.6151
R1138 B.n490 B.n80 10.6151
R1139 B.n484 B.n80 10.6151
R1140 B.n484 B.n483 10.6151
R1141 B.n483 B.n482 10.6151
R1142 B.n482 B.n82 10.6151
R1143 B.n476 B.n82 10.6151
R1144 B.n476 B.n475 10.6151
R1145 B.n475 B.n474 10.6151
R1146 B.n474 B.n84 10.6151
R1147 B.n468 B.n84 10.6151
R1148 B.n468 B.n467 10.6151
R1149 B.n467 B.n466 10.6151
R1150 B.n466 B.n86 10.6151
R1151 B.n460 B.n86 10.6151
R1152 B.n460 B.n459 10.6151
R1153 B.n459 B.n458 10.6151
R1154 B.n458 B.n88 10.6151
R1155 B.n452 B.n88 10.6151
R1156 B.n452 B.n451 10.6151
R1157 B.n697 B.n0 8.11757
R1158 B.n697 B.n1 8.11757
R1159 B.n288 B.n143 7.18099
R1160 B.n273 B.n272 7.18099
R1161 B.n567 B.n566 7.18099
R1162 B.n550 B.n64 7.18099
R1163 B.n292 B.n143 3.43465
R1164 B.n272 B.n271 3.43465
R1165 B.n568 B.n567 3.43465
R1166 B.n546 B.n64 3.43465
R1167 B.t3 B.n103 2.79025
R1168 B.n676 B.t10 2.79025
R1169 VN VN.t0 719.019
R1170 VN VN.t1 677.091
R1171 VDD2.n0 VDD2.t0 103.023
R1172 VDD2.n0 VDD2.t1 65.054
R1173 VDD2 VDD2.n0 0.291448
C0 VDD1 VP 2.50091f
C1 VTAIL VDD1 6.44976f
C2 VN VP 5.03041f
C3 VN VTAIL 1.79136f
C4 VDD2 VDD1 0.467613f
C5 VTAIL VP 1.80605f
C6 VN VDD2 2.39717f
C7 VDD2 VP 0.257769f
C8 VDD2 VTAIL 6.48282f
C9 VN VDD1 0.148945f
C10 VDD2 B 4.210034f
C11 VDD1 B 7.21595f
C12 VTAIL B 7.331822f
C13 VN B 8.66524f
C14 VP B 4.255111f
C15 VDD2.t0 B 3.26144f
C16 VDD2.t1 B 2.73851f
C17 VDD2.n0 B 2.84869f
C18 VN.t1 B 1.47078f
C19 VN.t0 B 1.59966f
C20 VDD1.t0 B 2.71613f
C21 VDD1.t1 B 3.25942f
C22 VTAIL.t3 B 2.0416f
C23 VTAIL.n0 B 1.19837f
C24 VTAIL.t1 B 2.04161f
C25 VTAIL.n1 B 1.20735f
C26 VTAIL.t2 B 2.0416f
C27 VTAIL.n2 B 1.15944f
C28 VTAIL.t0 B 2.0416f
C29 VTAIL.n3 B 1.12028f
C30 VP.t1 B 1.63206f
C31 VP.t0 B 1.50314f
C32 VP.n0 B 4.34781f
.ends

