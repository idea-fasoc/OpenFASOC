* NGSPICE file created from diff_pair_sample_0550.ext - technology: sky130A

.subckt diff_pair_sample_0550 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=0.58905 pd=3.9 as=1.3923 ps=7.92 w=3.57 l=3.28
X1 VDD2.t5 VN.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.3923 pd=7.92 as=0.58905 ps=3.9 w=3.57 l=3.28
X2 VTAIL.t3 VN.t1 VDD2.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.58905 pd=3.9 as=0.58905 ps=3.9 w=3.57 l=3.28
X3 VDD2.t3 VN.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.58905 pd=3.9 as=1.3923 ps=7.92 w=3.57 l=3.28
X4 VTAIL.t10 VP.t1 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.58905 pd=3.9 as=0.58905 ps=3.9 w=3.57 l=3.28
X5 VTAIL.t6 VP.t2 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.58905 pd=3.9 as=0.58905 ps=3.9 w=3.57 l=3.28
X6 VDD1.t2 VP.t3 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=1.3923 pd=7.92 as=0.58905 ps=3.9 w=3.57 l=3.28
X7 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=1.3923 pd=7.92 as=0 ps=0 w=3.57 l=3.28
X8 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=1.3923 pd=7.92 as=0 ps=0 w=3.57 l=3.28
X9 VTAIL.t2 VN.t3 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.58905 pd=3.9 as=0.58905 ps=3.9 w=3.57 l=3.28
X10 VDD1.t1 VP.t4 VTAIL.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=1.3923 pd=7.92 as=0.58905 ps=3.9 w=3.57 l=3.28
X11 VDD2.t1 VN.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.58905 pd=3.9 as=1.3923 ps=7.92 w=3.57 l=3.28
X12 VDD2.t0 VN.t5 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=1.3923 pd=7.92 as=0.58905 ps=3.9 w=3.57 l=3.28
X13 VDD1.t0 VP.t5 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=0.58905 pd=3.9 as=1.3923 ps=7.92 w=3.57 l=3.28
X14 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.3923 pd=7.92 as=0 ps=0 w=3.57 l=3.28
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.3923 pd=7.92 as=0 ps=0 w=3.57 l=3.28
R0 VP.n16 VP.n15 161.3
R1 VP.n17 VP.n12 161.3
R2 VP.n19 VP.n18 161.3
R3 VP.n20 VP.n11 161.3
R4 VP.n22 VP.n21 161.3
R5 VP.n23 VP.n10 161.3
R6 VP.n25 VP.n24 161.3
R7 VP.n49 VP.n48 161.3
R8 VP.n47 VP.n1 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n44 VP.n2 161.3
R11 VP.n43 VP.n42 161.3
R12 VP.n41 VP.n3 161.3
R13 VP.n40 VP.n39 161.3
R14 VP.n38 VP.n37 161.3
R15 VP.n36 VP.n5 161.3
R16 VP.n35 VP.n34 161.3
R17 VP.n33 VP.n6 161.3
R18 VP.n32 VP.n31 161.3
R19 VP.n30 VP.n7 161.3
R20 VP.n29 VP.n28 161.3
R21 VP.n27 VP.n8 72.4512
R22 VP.n50 VP.n0 72.4512
R23 VP.n26 VP.n9 72.4512
R24 VP.n14 VP.n13 62.0548
R25 VP.n14 VP.t3 59.4458
R26 VP.n31 VP.n6 45.8354
R27 VP.n46 VP.n2 45.8354
R28 VP.n22 VP.n11 45.8354
R29 VP.n27 VP.n26 45.1092
R30 VP.n35 VP.n6 35.1514
R31 VP.n42 VP.n2 35.1514
R32 VP.n18 VP.n11 35.1514
R33 VP.n8 VP.t4 26.2313
R34 VP.n4 VP.t2 26.2313
R35 VP.n0 VP.t0 26.2313
R36 VP.n9 VP.t5 26.2313
R37 VP.n13 VP.t1 26.2313
R38 VP.n30 VP.n29 24.4675
R39 VP.n31 VP.n30 24.4675
R40 VP.n36 VP.n35 24.4675
R41 VP.n37 VP.n36 24.4675
R42 VP.n41 VP.n40 24.4675
R43 VP.n42 VP.n41 24.4675
R44 VP.n47 VP.n46 24.4675
R45 VP.n48 VP.n47 24.4675
R46 VP.n23 VP.n22 24.4675
R47 VP.n24 VP.n23 24.4675
R48 VP.n17 VP.n16 24.4675
R49 VP.n18 VP.n17 24.4675
R50 VP.n29 VP.n8 17.6167
R51 VP.n48 VP.n0 17.6167
R52 VP.n24 VP.n9 17.6167
R53 VP.n37 VP.n4 12.234
R54 VP.n40 VP.n4 12.234
R55 VP.n16 VP.n13 12.234
R56 VP.n15 VP.n14 4.01735
R57 VP.n26 VP.n25 0.354971
R58 VP.n28 VP.n27 0.354971
R59 VP.n50 VP.n49 0.354971
R60 VP VP.n50 0.26696
R61 VP.n15 VP.n12 0.189894
R62 VP.n19 VP.n12 0.189894
R63 VP.n20 VP.n19 0.189894
R64 VP.n21 VP.n20 0.189894
R65 VP.n21 VP.n10 0.189894
R66 VP.n25 VP.n10 0.189894
R67 VP.n28 VP.n7 0.189894
R68 VP.n32 VP.n7 0.189894
R69 VP.n33 VP.n32 0.189894
R70 VP.n34 VP.n33 0.189894
R71 VP.n34 VP.n5 0.189894
R72 VP.n38 VP.n5 0.189894
R73 VP.n39 VP.n38 0.189894
R74 VP.n39 VP.n3 0.189894
R75 VP.n43 VP.n3 0.189894
R76 VP.n44 VP.n43 0.189894
R77 VP.n45 VP.n44 0.189894
R78 VP.n45 VP.n1 0.189894
R79 VP.n49 VP.n1 0.189894
R80 VTAIL.n7 VTAIL.t1 65.9734
R81 VTAIL.n11 VTAIL.t0 65.9734
R82 VTAIL.n2 VTAIL.t9 65.9734
R83 VTAIL.n10 VTAIL.t8 65.9734
R84 VTAIL.n9 VTAIL.n8 60.4273
R85 VTAIL.n6 VTAIL.n5 60.4273
R86 VTAIL.n1 VTAIL.n0 60.4271
R87 VTAIL.n4 VTAIL.n3 60.4271
R88 VTAIL.n6 VTAIL.n4 21.6686
R89 VTAIL.n11 VTAIL.n10 18.5565
R90 VTAIL.n0 VTAIL.t11 5.54672
R91 VTAIL.n0 VTAIL.t2 5.54672
R92 VTAIL.n3 VTAIL.t5 5.54672
R93 VTAIL.n3 VTAIL.t6 5.54672
R94 VTAIL.n8 VTAIL.t7 5.54672
R95 VTAIL.n8 VTAIL.t10 5.54672
R96 VTAIL.n5 VTAIL.t4 5.54672
R97 VTAIL.n5 VTAIL.t3 5.54672
R98 VTAIL.n7 VTAIL.n6 3.11257
R99 VTAIL.n10 VTAIL.n9 3.11257
R100 VTAIL.n4 VTAIL.n2 3.11257
R101 VTAIL VTAIL.n11 2.27636
R102 VTAIL.n9 VTAIL.n7 2.02636
R103 VTAIL.n2 VTAIL.n1 2.02636
R104 VTAIL VTAIL.n1 0.836707
R105 VDD1 VDD1.t2 85.0445
R106 VDD1.n1 VDD1.t1 84.9309
R107 VDD1.n1 VDD1.n0 77.8285
R108 VDD1.n3 VDD1.n2 77.106
R109 VDD1.n3 VDD1.n1 39.0462
R110 VDD1.n2 VDD1.t4 5.54672
R111 VDD1.n2 VDD1.t0 5.54672
R112 VDD1.n0 VDD1.t3 5.54672
R113 VDD1.n0 VDD1.t5 5.54672
R114 VDD1 VDD1.n3 0.720328
R115 B.n547 B.n120 585
R116 B.n120 B.n93 585
R117 B.n549 B.n548 585
R118 B.n551 B.n119 585
R119 B.n554 B.n553 585
R120 B.n555 B.n118 585
R121 B.n557 B.n556 585
R122 B.n559 B.n117 585
R123 B.n562 B.n561 585
R124 B.n563 B.n116 585
R125 B.n565 B.n564 585
R126 B.n567 B.n115 585
R127 B.n570 B.n569 585
R128 B.n571 B.n114 585
R129 B.n573 B.n572 585
R130 B.n575 B.n113 585
R131 B.n577 B.n576 585
R132 B.n579 B.n578 585
R133 B.n582 B.n581 585
R134 B.n583 B.n108 585
R135 B.n585 B.n584 585
R136 B.n587 B.n107 585
R137 B.n590 B.n589 585
R138 B.n591 B.n106 585
R139 B.n593 B.n592 585
R140 B.n595 B.n105 585
R141 B.n598 B.n597 585
R142 B.n600 B.n102 585
R143 B.n602 B.n601 585
R144 B.n604 B.n101 585
R145 B.n607 B.n606 585
R146 B.n608 B.n100 585
R147 B.n610 B.n609 585
R148 B.n612 B.n99 585
R149 B.n615 B.n614 585
R150 B.n616 B.n98 585
R151 B.n618 B.n617 585
R152 B.n620 B.n97 585
R153 B.n623 B.n622 585
R154 B.n624 B.n96 585
R155 B.n626 B.n625 585
R156 B.n628 B.n95 585
R157 B.n631 B.n630 585
R158 B.n632 B.n94 585
R159 B.n546 B.n92 585
R160 B.n635 B.n92 585
R161 B.n545 B.n91 585
R162 B.n636 B.n91 585
R163 B.n544 B.n90 585
R164 B.n637 B.n90 585
R165 B.n543 B.n542 585
R166 B.n542 B.n86 585
R167 B.n541 B.n85 585
R168 B.n643 B.n85 585
R169 B.n540 B.n84 585
R170 B.n644 B.n84 585
R171 B.n539 B.n83 585
R172 B.n645 B.n83 585
R173 B.n538 B.n537 585
R174 B.n537 B.n79 585
R175 B.n536 B.n78 585
R176 B.n651 B.n78 585
R177 B.n535 B.n77 585
R178 B.n652 B.n77 585
R179 B.n534 B.n76 585
R180 B.n653 B.n76 585
R181 B.n533 B.n532 585
R182 B.n532 B.n72 585
R183 B.n531 B.n71 585
R184 B.n659 B.n71 585
R185 B.n530 B.n70 585
R186 B.n660 B.n70 585
R187 B.n529 B.n69 585
R188 B.n661 B.n69 585
R189 B.n528 B.n527 585
R190 B.n527 B.n65 585
R191 B.n526 B.n64 585
R192 B.n667 B.n64 585
R193 B.n525 B.n63 585
R194 B.n668 B.n63 585
R195 B.n524 B.n62 585
R196 B.n669 B.n62 585
R197 B.n523 B.n522 585
R198 B.n522 B.n58 585
R199 B.n521 B.n57 585
R200 B.n675 B.n57 585
R201 B.n520 B.n56 585
R202 B.n676 B.n56 585
R203 B.n519 B.n55 585
R204 B.n677 B.n55 585
R205 B.n518 B.n517 585
R206 B.n517 B.n51 585
R207 B.n516 B.n50 585
R208 B.n683 B.n50 585
R209 B.n515 B.n49 585
R210 B.n684 B.n49 585
R211 B.n514 B.n48 585
R212 B.n685 B.n48 585
R213 B.n513 B.n512 585
R214 B.n512 B.n44 585
R215 B.n511 B.n43 585
R216 B.n691 B.n43 585
R217 B.n510 B.n42 585
R218 B.n692 B.n42 585
R219 B.n509 B.n41 585
R220 B.n693 B.n41 585
R221 B.n508 B.n507 585
R222 B.n507 B.n37 585
R223 B.n506 B.n36 585
R224 B.n699 B.n36 585
R225 B.n505 B.n35 585
R226 B.n700 B.n35 585
R227 B.n504 B.n34 585
R228 B.n701 B.n34 585
R229 B.n503 B.n502 585
R230 B.n502 B.n30 585
R231 B.n501 B.n29 585
R232 B.n707 B.n29 585
R233 B.n500 B.n28 585
R234 B.n708 B.n28 585
R235 B.n499 B.n27 585
R236 B.n709 B.n27 585
R237 B.n498 B.n497 585
R238 B.n497 B.n23 585
R239 B.n496 B.n22 585
R240 B.n715 B.n22 585
R241 B.n495 B.n21 585
R242 B.n716 B.n21 585
R243 B.n494 B.n20 585
R244 B.n717 B.n20 585
R245 B.n493 B.n492 585
R246 B.n492 B.n19 585
R247 B.n491 B.n15 585
R248 B.n723 B.n15 585
R249 B.n490 B.n14 585
R250 B.n724 B.n14 585
R251 B.n489 B.n13 585
R252 B.n725 B.n13 585
R253 B.n488 B.n487 585
R254 B.n487 B.n12 585
R255 B.n486 B.n485 585
R256 B.n486 B.n8 585
R257 B.n484 B.n7 585
R258 B.n732 B.n7 585
R259 B.n483 B.n6 585
R260 B.n733 B.n6 585
R261 B.n482 B.n5 585
R262 B.n734 B.n5 585
R263 B.n481 B.n480 585
R264 B.n480 B.n4 585
R265 B.n479 B.n121 585
R266 B.n479 B.n478 585
R267 B.n469 B.n122 585
R268 B.n123 B.n122 585
R269 B.n471 B.n470 585
R270 B.n472 B.n471 585
R271 B.n468 B.n128 585
R272 B.n128 B.n127 585
R273 B.n467 B.n466 585
R274 B.n466 B.n465 585
R275 B.n130 B.n129 585
R276 B.n458 B.n130 585
R277 B.n457 B.n456 585
R278 B.n459 B.n457 585
R279 B.n455 B.n135 585
R280 B.n135 B.n134 585
R281 B.n454 B.n453 585
R282 B.n453 B.n452 585
R283 B.n137 B.n136 585
R284 B.n138 B.n137 585
R285 B.n445 B.n444 585
R286 B.n446 B.n445 585
R287 B.n443 B.n143 585
R288 B.n143 B.n142 585
R289 B.n442 B.n441 585
R290 B.n441 B.n440 585
R291 B.n145 B.n144 585
R292 B.n146 B.n145 585
R293 B.n433 B.n432 585
R294 B.n434 B.n433 585
R295 B.n431 B.n151 585
R296 B.n151 B.n150 585
R297 B.n430 B.n429 585
R298 B.n429 B.n428 585
R299 B.n153 B.n152 585
R300 B.n154 B.n153 585
R301 B.n421 B.n420 585
R302 B.n422 B.n421 585
R303 B.n419 B.n159 585
R304 B.n159 B.n158 585
R305 B.n418 B.n417 585
R306 B.n417 B.n416 585
R307 B.n161 B.n160 585
R308 B.n162 B.n161 585
R309 B.n409 B.n408 585
R310 B.n410 B.n409 585
R311 B.n407 B.n167 585
R312 B.n167 B.n166 585
R313 B.n406 B.n405 585
R314 B.n405 B.n404 585
R315 B.n169 B.n168 585
R316 B.n170 B.n169 585
R317 B.n397 B.n396 585
R318 B.n398 B.n397 585
R319 B.n395 B.n175 585
R320 B.n175 B.n174 585
R321 B.n394 B.n393 585
R322 B.n393 B.n392 585
R323 B.n177 B.n176 585
R324 B.n178 B.n177 585
R325 B.n385 B.n384 585
R326 B.n386 B.n385 585
R327 B.n383 B.n183 585
R328 B.n183 B.n182 585
R329 B.n382 B.n381 585
R330 B.n381 B.n380 585
R331 B.n185 B.n184 585
R332 B.n186 B.n185 585
R333 B.n373 B.n372 585
R334 B.n374 B.n373 585
R335 B.n371 B.n191 585
R336 B.n191 B.n190 585
R337 B.n370 B.n369 585
R338 B.n369 B.n368 585
R339 B.n193 B.n192 585
R340 B.n194 B.n193 585
R341 B.n361 B.n360 585
R342 B.n362 B.n361 585
R343 B.n359 B.n199 585
R344 B.n199 B.n198 585
R345 B.n358 B.n357 585
R346 B.n357 B.n356 585
R347 B.n201 B.n200 585
R348 B.n202 B.n201 585
R349 B.n349 B.n348 585
R350 B.n350 B.n349 585
R351 B.n347 B.n207 585
R352 B.n207 B.n206 585
R353 B.n346 B.n345 585
R354 B.n345 B.n344 585
R355 B.n209 B.n208 585
R356 B.n210 B.n209 585
R357 B.n337 B.n336 585
R358 B.n338 B.n337 585
R359 B.n335 B.n215 585
R360 B.n215 B.n214 585
R361 B.n334 B.n333 585
R362 B.n333 B.n332 585
R363 B.n329 B.n219 585
R364 B.n328 B.n327 585
R365 B.n325 B.n220 585
R366 B.n325 B.n218 585
R367 B.n324 B.n323 585
R368 B.n322 B.n321 585
R369 B.n320 B.n222 585
R370 B.n318 B.n317 585
R371 B.n316 B.n223 585
R372 B.n315 B.n314 585
R373 B.n312 B.n224 585
R374 B.n310 B.n309 585
R375 B.n308 B.n225 585
R376 B.n307 B.n306 585
R377 B.n304 B.n226 585
R378 B.n302 B.n301 585
R379 B.n300 B.n227 585
R380 B.n299 B.n298 585
R381 B.n296 B.n295 585
R382 B.n294 B.n293 585
R383 B.n292 B.n232 585
R384 B.n290 B.n289 585
R385 B.n288 B.n233 585
R386 B.n287 B.n286 585
R387 B.n284 B.n234 585
R388 B.n282 B.n281 585
R389 B.n280 B.n235 585
R390 B.n278 B.n277 585
R391 B.n275 B.n238 585
R392 B.n273 B.n272 585
R393 B.n271 B.n239 585
R394 B.n270 B.n269 585
R395 B.n267 B.n240 585
R396 B.n265 B.n264 585
R397 B.n263 B.n241 585
R398 B.n262 B.n261 585
R399 B.n259 B.n242 585
R400 B.n257 B.n256 585
R401 B.n255 B.n243 585
R402 B.n254 B.n253 585
R403 B.n251 B.n244 585
R404 B.n249 B.n248 585
R405 B.n247 B.n246 585
R406 B.n217 B.n216 585
R407 B.n331 B.n330 585
R408 B.n332 B.n331 585
R409 B.n213 B.n212 585
R410 B.n214 B.n213 585
R411 B.n340 B.n339 585
R412 B.n339 B.n338 585
R413 B.n341 B.n211 585
R414 B.n211 B.n210 585
R415 B.n343 B.n342 585
R416 B.n344 B.n343 585
R417 B.n205 B.n204 585
R418 B.n206 B.n205 585
R419 B.n352 B.n351 585
R420 B.n351 B.n350 585
R421 B.n353 B.n203 585
R422 B.n203 B.n202 585
R423 B.n355 B.n354 585
R424 B.n356 B.n355 585
R425 B.n197 B.n196 585
R426 B.n198 B.n197 585
R427 B.n364 B.n363 585
R428 B.n363 B.n362 585
R429 B.n365 B.n195 585
R430 B.n195 B.n194 585
R431 B.n367 B.n366 585
R432 B.n368 B.n367 585
R433 B.n189 B.n188 585
R434 B.n190 B.n189 585
R435 B.n376 B.n375 585
R436 B.n375 B.n374 585
R437 B.n377 B.n187 585
R438 B.n187 B.n186 585
R439 B.n379 B.n378 585
R440 B.n380 B.n379 585
R441 B.n181 B.n180 585
R442 B.n182 B.n181 585
R443 B.n388 B.n387 585
R444 B.n387 B.n386 585
R445 B.n389 B.n179 585
R446 B.n179 B.n178 585
R447 B.n391 B.n390 585
R448 B.n392 B.n391 585
R449 B.n173 B.n172 585
R450 B.n174 B.n173 585
R451 B.n400 B.n399 585
R452 B.n399 B.n398 585
R453 B.n401 B.n171 585
R454 B.n171 B.n170 585
R455 B.n403 B.n402 585
R456 B.n404 B.n403 585
R457 B.n165 B.n164 585
R458 B.n166 B.n165 585
R459 B.n412 B.n411 585
R460 B.n411 B.n410 585
R461 B.n413 B.n163 585
R462 B.n163 B.n162 585
R463 B.n415 B.n414 585
R464 B.n416 B.n415 585
R465 B.n157 B.n156 585
R466 B.n158 B.n157 585
R467 B.n424 B.n423 585
R468 B.n423 B.n422 585
R469 B.n425 B.n155 585
R470 B.n155 B.n154 585
R471 B.n427 B.n426 585
R472 B.n428 B.n427 585
R473 B.n149 B.n148 585
R474 B.n150 B.n149 585
R475 B.n436 B.n435 585
R476 B.n435 B.n434 585
R477 B.n437 B.n147 585
R478 B.n147 B.n146 585
R479 B.n439 B.n438 585
R480 B.n440 B.n439 585
R481 B.n141 B.n140 585
R482 B.n142 B.n141 585
R483 B.n448 B.n447 585
R484 B.n447 B.n446 585
R485 B.n449 B.n139 585
R486 B.n139 B.n138 585
R487 B.n451 B.n450 585
R488 B.n452 B.n451 585
R489 B.n133 B.n132 585
R490 B.n134 B.n133 585
R491 B.n461 B.n460 585
R492 B.n460 B.n459 585
R493 B.n462 B.n131 585
R494 B.n458 B.n131 585
R495 B.n464 B.n463 585
R496 B.n465 B.n464 585
R497 B.n126 B.n125 585
R498 B.n127 B.n126 585
R499 B.n474 B.n473 585
R500 B.n473 B.n472 585
R501 B.n475 B.n124 585
R502 B.n124 B.n123 585
R503 B.n477 B.n476 585
R504 B.n478 B.n477 585
R505 B.n3 B.n0 585
R506 B.n4 B.n3 585
R507 B.n731 B.n1 585
R508 B.n732 B.n731 585
R509 B.n730 B.n729 585
R510 B.n730 B.n8 585
R511 B.n728 B.n9 585
R512 B.n12 B.n9 585
R513 B.n727 B.n726 585
R514 B.n726 B.n725 585
R515 B.n11 B.n10 585
R516 B.n724 B.n11 585
R517 B.n722 B.n721 585
R518 B.n723 B.n722 585
R519 B.n720 B.n16 585
R520 B.n19 B.n16 585
R521 B.n719 B.n718 585
R522 B.n718 B.n717 585
R523 B.n18 B.n17 585
R524 B.n716 B.n18 585
R525 B.n714 B.n713 585
R526 B.n715 B.n714 585
R527 B.n712 B.n24 585
R528 B.n24 B.n23 585
R529 B.n711 B.n710 585
R530 B.n710 B.n709 585
R531 B.n26 B.n25 585
R532 B.n708 B.n26 585
R533 B.n706 B.n705 585
R534 B.n707 B.n706 585
R535 B.n704 B.n31 585
R536 B.n31 B.n30 585
R537 B.n703 B.n702 585
R538 B.n702 B.n701 585
R539 B.n33 B.n32 585
R540 B.n700 B.n33 585
R541 B.n698 B.n697 585
R542 B.n699 B.n698 585
R543 B.n696 B.n38 585
R544 B.n38 B.n37 585
R545 B.n695 B.n694 585
R546 B.n694 B.n693 585
R547 B.n40 B.n39 585
R548 B.n692 B.n40 585
R549 B.n690 B.n689 585
R550 B.n691 B.n690 585
R551 B.n688 B.n45 585
R552 B.n45 B.n44 585
R553 B.n687 B.n686 585
R554 B.n686 B.n685 585
R555 B.n47 B.n46 585
R556 B.n684 B.n47 585
R557 B.n682 B.n681 585
R558 B.n683 B.n682 585
R559 B.n680 B.n52 585
R560 B.n52 B.n51 585
R561 B.n679 B.n678 585
R562 B.n678 B.n677 585
R563 B.n54 B.n53 585
R564 B.n676 B.n54 585
R565 B.n674 B.n673 585
R566 B.n675 B.n674 585
R567 B.n672 B.n59 585
R568 B.n59 B.n58 585
R569 B.n671 B.n670 585
R570 B.n670 B.n669 585
R571 B.n61 B.n60 585
R572 B.n668 B.n61 585
R573 B.n666 B.n665 585
R574 B.n667 B.n666 585
R575 B.n664 B.n66 585
R576 B.n66 B.n65 585
R577 B.n663 B.n662 585
R578 B.n662 B.n661 585
R579 B.n68 B.n67 585
R580 B.n660 B.n68 585
R581 B.n658 B.n657 585
R582 B.n659 B.n658 585
R583 B.n656 B.n73 585
R584 B.n73 B.n72 585
R585 B.n655 B.n654 585
R586 B.n654 B.n653 585
R587 B.n75 B.n74 585
R588 B.n652 B.n75 585
R589 B.n650 B.n649 585
R590 B.n651 B.n650 585
R591 B.n648 B.n80 585
R592 B.n80 B.n79 585
R593 B.n647 B.n646 585
R594 B.n646 B.n645 585
R595 B.n82 B.n81 585
R596 B.n644 B.n82 585
R597 B.n642 B.n641 585
R598 B.n643 B.n642 585
R599 B.n640 B.n87 585
R600 B.n87 B.n86 585
R601 B.n639 B.n638 585
R602 B.n638 B.n637 585
R603 B.n89 B.n88 585
R604 B.n636 B.n89 585
R605 B.n634 B.n633 585
R606 B.n635 B.n634 585
R607 B.n735 B.n734 585
R608 B.n733 B.n2 585
R609 B.n634 B.n94 530.939
R610 B.n120 B.n92 530.939
R611 B.n333 B.n217 530.939
R612 B.n331 B.n219 530.939
R613 B.n550 B.n93 256.663
R614 B.n552 B.n93 256.663
R615 B.n558 B.n93 256.663
R616 B.n560 B.n93 256.663
R617 B.n566 B.n93 256.663
R618 B.n568 B.n93 256.663
R619 B.n574 B.n93 256.663
R620 B.n112 B.n93 256.663
R621 B.n580 B.n93 256.663
R622 B.n586 B.n93 256.663
R623 B.n588 B.n93 256.663
R624 B.n594 B.n93 256.663
R625 B.n596 B.n93 256.663
R626 B.n603 B.n93 256.663
R627 B.n605 B.n93 256.663
R628 B.n611 B.n93 256.663
R629 B.n613 B.n93 256.663
R630 B.n619 B.n93 256.663
R631 B.n621 B.n93 256.663
R632 B.n627 B.n93 256.663
R633 B.n629 B.n93 256.663
R634 B.n326 B.n218 256.663
R635 B.n221 B.n218 256.663
R636 B.n319 B.n218 256.663
R637 B.n313 B.n218 256.663
R638 B.n311 B.n218 256.663
R639 B.n305 B.n218 256.663
R640 B.n303 B.n218 256.663
R641 B.n297 B.n218 256.663
R642 B.n231 B.n218 256.663
R643 B.n291 B.n218 256.663
R644 B.n285 B.n218 256.663
R645 B.n283 B.n218 256.663
R646 B.n276 B.n218 256.663
R647 B.n274 B.n218 256.663
R648 B.n268 B.n218 256.663
R649 B.n266 B.n218 256.663
R650 B.n260 B.n218 256.663
R651 B.n258 B.n218 256.663
R652 B.n252 B.n218 256.663
R653 B.n250 B.n218 256.663
R654 B.n245 B.n218 256.663
R655 B.n737 B.n736 256.663
R656 B.n103 B.t10 235.115
R657 B.n109 B.t14 235.115
R658 B.n236 B.t6 235.115
R659 B.n228 B.t17 235.115
R660 B.n630 B.n628 163.367
R661 B.n626 B.n96 163.367
R662 B.n622 B.n620 163.367
R663 B.n618 B.n98 163.367
R664 B.n614 B.n612 163.367
R665 B.n610 B.n100 163.367
R666 B.n606 B.n604 163.367
R667 B.n602 B.n102 163.367
R668 B.n597 B.n595 163.367
R669 B.n593 B.n106 163.367
R670 B.n589 B.n587 163.367
R671 B.n585 B.n108 163.367
R672 B.n581 B.n579 163.367
R673 B.n576 B.n575 163.367
R674 B.n573 B.n114 163.367
R675 B.n569 B.n567 163.367
R676 B.n565 B.n116 163.367
R677 B.n561 B.n559 163.367
R678 B.n557 B.n118 163.367
R679 B.n553 B.n551 163.367
R680 B.n549 B.n120 163.367
R681 B.n333 B.n215 163.367
R682 B.n337 B.n215 163.367
R683 B.n337 B.n209 163.367
R684 B.n345 B.n209 163.367
R685 B.n345 B.n207 163.367
R686 B.n349 B.n207 163.367
R687 B.n349 B.n201 163.367
R688 B.n357 B.n201 163.367
R689 B.n357 B.n199 163.367
R690 B.n361 B.n199 163.367
R691 B.n361 B.n193 163.367
R692 B.n369 B.n193 163.367
R693 B.n369 B.n191 163.367
R694 B.n373 B.n191 163.367
R695 B.n373 B.n185 163.367
R696 B.n381 B.n185 163.367
R697 B.n381 B.n183 163.367
R698 B.n385 B.n183 163.367
R699 B.n385 B.n177 163.367
R700 B.n393 B.n177 163.367
R701 B.n393 B.n175 163.367
R702 B.n397 B.n175 163.367
R703 B.n397 B.n169 163.367
R704 B.n405 B.n169 163.367
R705 B.n405 B.n167 163.367
R706 B.n409 B.n167 163.367
R707 B.n409 B.n161 163.367
R708 B.n417 B.n161 163.367
R709 B.n417 B.n159 163.367
R710 B.n421 B.n159 163.367
R711 B.n421 B.n153 163.367
R712 B.n429 B.n153 163.367
R713 B.n429 B.n151 163.367
R714 B.n433 B.n151 163.367
R715 B.n433 B.n145 163.367
R716 B.n441 B.n145 163.367
R717 B.n441 B.n143 163.367
R718 B.n445 B.n143 163.367
R719 B.n445 B.n137 163.367
R720 B.n453 B.n137 163.367
R721 B.n453 B.n135 163.367
R722 B.n457 B.n135 163.367
R723 B.n457 B.n130 163.367
R724 B.n466 B.n130 163.367
R725 B.n466 B.n128 163.367
R726 B.n471 B.n128 163.367
R727 B.n471 B.n122 163.367
R728 B.n479 B.n122 163.367
R729 B.n480 B.n479 163.367
R730 B.n480 B.n5 163.367
R731 B.n6 B.n5 163.367
R732 B.n7 B.n6 163.367
R733 B.n486 B.n7 163.367
R734 B.n487 B.n486 163.367
R735 B.n487 B.n13 163.367
R736 B.n14 B.n13 163.367
R737 B.n15 B.n14 163.367
R738 B.n492 B.n15 163.367
R739 B.n492 B.n20 163.367
R740 B.n21 B.n20 163.367
R741 B.n22 B.n21 163.367
R742 B.n497 B.n22 163.367
R743 B.n497 B.n27 163.367
R744 B.n28 B.n27 163.367
R745 B.n29 B.n28 163.367
R746 B.n502 B.n29 163.367
R747 B.n502 B.n34 163.367
R748 B.n35 B.n34 163.367
R749 B.n36 B.n35 163.367
R750 B.n507 B.n36 163.367
R751 B.n507 B.n41 163.367
R752 B.n42 B.n41 163.367
R753 B.n43 B.n42 163.367
R754 B.n512 B.n43 163.367
R755 B.n512 B.n48 163.367
R756 B.n49 B.n48 163.367
R757 B.n50 B.n49 163.367
R758 B.n517 B.n50 163.367
R759 B.n517 B.n55 163.367
R760 B.n56 B.n55 163.367
R761 B.n57 B.n56 163.367
R762 B.n522 B.n57 163.367
R763 B.n522 B.n62 163.367
R764 B.n63 B.n62 163.367
R765 B.n64 B.n63 163.367
R766 B.n527 B.n64 163.367
R767 B.n527 B.n69 163.367
R768 B.n70 B.n69 163.367
R769 B.n71 B.n70 163.367
R770 B.n532 B.n71 163.367
R771 B.n532 B.n76 163.367
R772 B.n77 B.n76 163.367
R773 B.n78 B.n77 163.367
R774 B.n537 B.n78 163.367
R775 B.n537 B.n83 163.367
R776 B.n84 B.n83 163.367
R777 B.n85 B.n84 163.367
R778 B.n542 B.n85 163.367
R779 B.n542 B.n90 163.367
R780 B.n91 B.n90 163.367
R781 B.n92 B.n91 163.367
R782 B.n327 B.n325 163.367
R783 B.n325 B.n324 163.367
R784 B.n321 B.n320 163.367
R785 B.n318 B.n223 163.367
R786 B.n314 B.n312 163.367
R787 B.n310 B.n225 163.367
R788 B.n306 B.n304 163.367
R789 B.n302 B.n227 163.367
R790 B.n298 B.n296 163.367
R791 B.n293 B.n292 163.367
R792 B.n290 B.n233 163.367
R793 B.n286 B.n284 163.367
R794 B.n282 B.n235 163.367
R795 B.n277 B.n275 163.367
R796 B.n273 B.n239 163.367
R797 B.n269 B.n267 163.367
R798 B.n265 B.n241 163.367
R799 B.n261 B.n259 163.367
R800 B.n257 B.n243 163.367
R801 B.n253 B.n251 163.367
R802 B.n249 B.n246 163.367
R803 B.n331 B.n213 163.367
R804 B.n339 B.n213 163.367
R805 B.n339 B.n211 163.367
R806 B.n343 B.n211 163.367
R807 B.n343 B.n205 163.367
R808 B.n351 B.n205 163.367
R809 B.n351 B.n203 163.367
R810 B.n355 B.n203 163.367
R811 B.n355 B.n197 163.367
R812 B.n363 B.n197 163.367
R813 B.n363 B.n195 163.367
R814 B.n367 B.n195 163.367
R815 B.n367 B.n189 163.367
R816 B.n375 B.n189 163.367
R817 B.n375 B.n187 163.367
R818 B.n379 B.n187 163.367
R819 B.n379 B.n181 163.367
R820 B.n387 B.n181 163.367
R821 B.n387 B.n179 163.367
R822 B.n391 B.n179 163.367
R823 B.n391 B.n173 163.367
R824 B.n399 B.n173 163.367
R825 B.n399 B.n171 163.367
R826 B.n403 B.n171 163.367
R827 B.n403 B.n165 163.367
R828 B.n411 B.n165 163.367
R829 B.n411 B.n163 163.367
R830 B.n415 B.n163 163.367
R831 B.n415 B.n157 163.367
R832 B.n423 B.n157 163.367
R833 B.n423 B.n155 163.367
R834 B.n427 B.n155 163.367
R835 B.n427 B.n149 163.367
R836 B.n435 B.n149 163.367
R837 B.n435 B.n147 163.367
R838 B.n439 B.n147 163.367
R839 B.n439 B.n141 163.367
R840 B.n447 B.n141 163.367
R841 B.n447 B.n139 163.367
R842 B.n451 B.n139 163.367
R843 B.n451 B.n133 163.367
R844 B.n460 B.n133 163.367
R845 B.n460 B.n131 163.367
R846 B.n464 B.n131 163.367
R847 B.n464 B.n126 163.367
R848 B.n473 B.n126 163.367
R849 B.n473 B.n124 163.367
R850 B.n477 B.n124 163.367
R851 B.n477 B.n3 163.367
R852 B.n735 B.n3 163.367
R853 B.n731 B.n2 163.367
R854 B.n731 B.n730 163.367
R855 B.n730 B.n9 163.367
R856 B.n726 B.n9 163.367
R857 B.n726 B.n11 163.367
R858 B.n722 B.n11 163.367
R859 B.n722 B.n16 163.367
R860 B.n718 B.n16 163.367
R861 B.n718 B.n18 163.367
R862 B.n714 B.n18 163.367
R863 B.n714 B.n24 163.367
R864 B.n710 B.n24 163.367
R865 B.n710 B.n26 163.367
R866 B.n706 B.n26 163.367
R867 B.n706 B.n31 163.367
R868 B.n702 B.n31 163.367
R869 B.n702 B.n33 163.367
R870 B.n698 B.n33 163.367
R871 B.n698 B.n38 163.367
R872 B.n694 B.n38 163.367
R873 B.n694 B.n40 163.367
R874 B.n690 B.n40 163.367
R875 B.n690 B.n45 163.367
R876 B.n686 B.n45 163.367
R877 B.n686 B.n47 163.367
R878 B.n682 B.n47 163.367
R879 B.n682 B.n52 163.367
R880 B.n678 B.n52 163.367
R881 B.n678 B.n54 163.367
R882 B.n674 B.n54 163.367
R883 B.n674 B.n59 163.367
R884 B.n670 B.n59 163.367
R885 B.n670 B.n61 163.367
R886 B.n666 B.n61 163.367
R887 B.n666 B.n66 163.367
R888 B.n662 B.n66 163.367
R889 B.n662 B.n68 163.367
R890 B.n658 B.n68 163.367
R891 B.n658 B.n73 163.367
R892 B.n654 B.n73 163.367
R893 B.n654 B.n75 163.367
R894 B.n650 B.n75 163.367
R895 B.n650 B.n80 163.367
R896 B.n646 B.n80 163.367
R897 B.n646 B.n82 163.367
R898 B.n642 B.n82 163.367
R899 B.n642 B.n87 163.367
R900 B.n638 B.n87 163.367
R901 B.n638 B.n89 163.367
R902 B.n634 B.n89 163.367
R903 B.n332 B.n218 160.43
R904 B.n635 B.n93 160.43
R905 B.n109 B.t15 145.816
R906 B.n236 B.t9 145.816
R907 B.n103 B.t12 145.814
R908 B.n228 B.t19 145.814
R909 B.n332 B.n214 84.5681
R910 B.n338 B.n214 84.5681
R911 B.n338 B.n210 84.5681
R912 B.n344 B.n210 84.5681
R913 B.n344 B.n206 84.5681
R914 B.n350 B.n206 84.5681
R915 B.n350 B.n202 84.5681
R916 B.n356 B.n202 84.5681
R917 B.n362 B.n198 84.5681
R918 B.n362 B.n194 84.5681
R919 B.n368 B.n194 84.5681
R920 B.n368 B.n190 84.5681
R921 B.n374 B.n190 84.5681
R922 B.n374 B.n186 84.5681
R923 B.n380 B.n186 84.5681
R924 B.n380 B.n182 84.5681
R925 B.n386 B.n182 84.5681
R926 B.n386 B.n178 84.5681
R927 B.n392 B.n178 84.5681
R928 B.n392 B.n174 84.5681
R929 B.n398 B.n174 84.5681
R930 B.n404 B.n170 84.5681
R931 B.n404 B.n166 84.5681
R932 B.n410 B.n166 84.5681
R933 B.n410 B.n162 84.5681
R934 B.n416 B.n162 84.5681
R935 B.n416 B.n158 84.5681
R936 B.n422 B.n158 84.5681
R937 B.n422 B.n154 84.5681
R938 B.n428 B.n154 84.5681
R939 B.n434 B.n150 84.5681
R940 B.n434 B.n146 84.5681
R941 B.n440 B.n146 84.5681
R942 B.n440 B.n142 84.5681
R943 B.n446 B.n142 84.5681
R944 B.n446 B.n138 84.5681
R945 B.n452 B.n138 84.5681
R946 B.n452 B.n134 84.5681
R947 B.n459 B.n134 84.5681
R948 B.n459 B.n458 84.5681
R949 B.n465 B.n127 84.5681
R950 B.n472 B.n127 84.5681
R951 B.n472 B.n123 84.5681
R952 B.n478 B.n123 84.5681
R953 B.n478 B.n4 84.5681
R954 B.n734 B.n4 84.5681
R955 B.n734 B.n733 84.5681
R956 B.n733 B.n732 84.5681
R957 B.n732 B.n8 84.5681
R958 B.n12 B.n8 84.5681
R959 B.n725 B.n12 84.5681
R960 B.n725 B.n724 84.5681
R961 B.n724 B.n723 84.5681
R962 B.n717 B.n19 84.5681
R963 B.n717 B.n716 84.5681
R964 B.n716 B.n715 84.5681
R965 B.n715 B.n23 84.5681
R966 B.n709 B.n23 84.5681
R967 B.n709 B.n708 84.5681
R968 B.n708 B.n707 84.5681
R969 B.n707 B.n30 84.5681
R970 B.n701 B.n30 84.5681
R971 B.n701 B.n700 84.5681
R972 B.n699 B.n37 84.5681
R973 B.n693 B.n37 84.5681
R974 B.n693 B.n692 84.5681
R975 B.n692 B.n691 84.5681
R976 B.n691 B.n44 84.5681
R977 B.n685 B.n44 84.5681
R978 B.n685 B.n684 84.5681
R979 B.n684 B.n683 84.5681
R980 B.n683 B.n51 84.5681
R981 B.n677 B.n676 84.5681
R982 B.n676 B.n675 84.5681
R983 B.n675 B.n58 84.5681
R984 B.n669 B.n58 84.5681
R985 B.n669 B.n668 84.5681
R986 B.n668 B.n667 84.5681
R987 B.n667 B.n65 84.5681
R988 B.n661 B.n65 84.5681
R989 B.n661 B.n660 84.5681
R990 B.n660 B.n659 84.5681
R991 B.n659 B.n72 84.5681
R992 B.n653 B.n72 84.5681
R993 B.n653 B.n652 84.5681
R994 B.n651 B.n79 84.5681
R995 B.n645 B.n79 84.5681
R996 B.n645 B.n644 84.5681
R997 B.n644 B.n643 84.5681
R998 B.n643 B.n86 84.5681
R999 B.n637 B.n86 84.5681
R1000 B.n637 B.n636 84.5681
R1001 B.n636 B.n635 84.5681
R1002 B.n428 B.t3 82.0808
R1003 B.t2 B.n699 82.0808
R1004 B.n110 B.t16 75.8048
R1005 B.n237 B.t8 75.8048
R1006 B.n104 B.t13 75.8018
R1007 B.n229 B.t18 75.8018
R1008 B.n629 B.n94 71.676
R1009 B.n628 B.n627 71.676
R1010 B.n621 B.n96 71.676
R1011 B.n620 B.n619 71.676
R1012 B.n613 B.n98 71.676
R1013 B.n612 B.n611 71.676
R1014 B.n605 B.n100 71.676
R1015 B.n604 B.n603 71.676
R1016 B.n596 B.n102 71.676
R1017 B.n595 B.n594 71.676
R1018 B.n588 B.n106 71.676
R1019 B.n587 B.n586 71.676
R1020 B.n580 B.n108 71.676
R1021 B.n579 B.n112 71.676
R1022 B.n575 B.n574 71.676
R1023 B.n568 B.n114 71.676
R1024 B.n567 B.n566 71.676
R1025 B.n560 B.n116 71.676
R1026 B.n559 B.n558 71.676
R1027 B.n552 B.n118 71.676
R1028 B.n551 B.n550 71.676
R1029 B.n550 B.n549 71.676
R1030 B.n553 B.n552 71.676
R1031 B.n558 B.n557 71.676
R1032 B.n561 B.n560 71.676
R1033 B.n566 B.n565 71.676
R1034 B.n569 B.n568 71.676
R1035 B.n574 B.n573 71.676
R1036 B.n576 B.n112 71.676
R1037 B.n581 B.n580 71.676
R1038 B.n586 B.n585 71.676
R1039 B.n589 B.n588 71.676
R1040 B.n594 B.n593 71.676
R1041 B.n597 B.n596 71.676
R1042 B.n603 B.n602 71.676
R1043 B.n606 B.n605 71.676
R1044 B.n611 B.n610 71.676
R1045 B.n614 B.n613 71.676
R1046 B.n619 B.n618 71.676
R1047 B.n622 B.n621 71.676
R1048 B.n627 B.n626 71.676
R1049 B.n630 B.n629 71.676
R1050 B.n326 B.n219 71.676
R1051 B.n324 B.n221 71.676
R1052 B.n320 B.n319 71.676
R1053 B.n313 B.n223 71.676
R1054 B.n312 B.n311 71.676
R1055 B.n305 B.n225 71.676
R1056 B.n304 B.n303 71.676
R1057 B.n297 B.n227 71.676
R1058 B.n296 B.n231 71.676
R1059 B.n292 B.n291 71.676
R1060 B.n285 B.n233 71.676
R1061 B.n284 B.n283 71.676
R1062 B.n276 B.n235 71.676
R1063 B.n275 B.n274 71.676
R1064 B.n268 B.n239 71.676
R1065 B.n267 B.n266 71.676
R1066 B.n260 B.n241 71.676
R1067 B.n259 B.n258 71.676
R1068 B.n252 B.n243 71.676
R1069 B.n251 B.n250 71.676
R1070 B.n246 B.n245 71.676
R1071 B.n327 B.n326 71.676
R1072 B.n321 B.n221 71.676
R1073 B.n319 B.n318 71.676
R1074 B.n314 B.n313 71.676
R1075 B.n311 B.n310 71.676
R1076 B.n306 B.n305 71.676
R1077 B.n303 B.n302 71.676
R1078 B.n298 B.n297 71.676
R1079 B.n293 B.n231 71.676
R1080 B.n291 B.n290 71.676
R1081 B.n286 B.n285 71.676
R1082 B.n283 B.n282 71.676
R1083 B.n277 B.n276 71.676
R1084 B.n274 B.n273 71.676
R1085 B.n269 B.n268 71.676
R1086 B.n266 B.n265 71.676
R1087 B.n261 B.n260 71.676
R1088 B.n258 B.n257 71.676
R1089 B.n253 B.n252 71.676
R1090 B.n250 B.n249 71.676
R1091 B.n245 B.n217 71.676
R1092 B.n736 B.n735 71.676
R1093 B.n736 B.n2 71.676
R1094 B.n104 B.n103 70.0126
R1095 B.n110 B.n109 70.0126
R1096 B.n237 B.n236 70.0126
R1097 B.n229 B.n228 70.0126
R1098 B.n599 B.n104 59.5399
R1099 B.n111 B.n110 59.5399
R1100 B.n279 B.n237 59.5399
R1101 B.n230 B.n229 59.5399
R1102 B.t4 B.n170 54.7207
R1103 B.t0 B.n51 54.7207
R1104 B.n458 B.t1 49.7461
R1105 B.n19 B.t5 49.7461
R1106 B.n356 B.t7 44.7716
R1107 B.t11 B.n651 44.7716
R1108 B.t7 B.n198 39.797
R1109 B.n652 B.t11 39.797
R1110 B.n465 B.t1 34.8224
R1111 B.n723 B.t5 34.8224
R1112 B.n330 B.n329 34.4981
R1113 B.n334 B.n216 34.4981
R1114 B.n547 B.n546 34.4981
R1115 B.n633 B.n632 34.4981
R1116 B.n398 B.t4 29.8479
R1117 B.n677 B.t0 29.8479
R1118 B B.n737 18.0485
R1119 B.n330 B.n212 10.6151
R1120 B.n340 B.n212 10.6151
R1121 B.n341 B.n340 10.6151
R1122 B.n342 B.n341 10.6151
R1123 B.n342 B.n204 10.6151
R1124 B.n352 B.n204 10.6151
R1125 B.n353 B.n352 10.6151
R1126 B.n354 B.n353 10.6151
R1127 B.n354 B.n196 10.6151
R1128 B.n364 B.n196 10.6151
R1129 B.n365 B.n364 10.6151
R1130 B.n366 B.n365 10.6151
R1131 B.n366 B.n188 10.6151
R1132 B.n376 B.n188 10.6151
R1133 B.n377 B.n376 10.6151
R1134 B.n378 B.n377 10.6151
R1135 B.n378 B.n180 10.6151
R1136 B.n388 B.n180 10.6151
R1137 B.n389 B.n388 10.6151
R1138 B.n390 B.n389 10.6151
R1139 B.n390 B.n172 10.6151
R1140 B.n400 B.n172 10.6151
R1141 B.n401 B.n400 10.6151
R1142 B.n402 B.n401 10.6151
R1143 B.n402 B.n164 10.6151
R1144 B.n412 B.n164 10.6151
R1145 B.n413 B.n412 10.6151
R1146 B.n414 B.n413 10.6151
R1147 B.n414 B.n156 10.6151
R1148 B.n424 B.n156 10.6151
R1149 B.n425 B.n424 10.6151
R1150 B.n426 B.n425 10.6151
R1151 B.n426 B.n148 10.6151
R1152 B.n436 B.n148 10.6151
R1153 B.n437 B.n436 10.6151
R1154 B.n438 B.n437 10.6151
R1155 B.n438 B.n140 10.6151
R1156 B.n448 B.n140 10.6151
R1157 B.n449 B.n448 10.6151
R1158 B.n450 B.n449 10.6151
R1159 B.n450 B.n132 10.6151
R1160 B.n461 B.n132 10.6151
R1161 B.n462 B.n461 10.6151
R1162 B.n463 B.n462 10.6151
R1163 B.n463 B.n125 10.6151
R1164 B.n474 B.n125 10.6151
R1165 B.n475 B.n474 10.6151
R1166 B.n476 B.n475 10.6151
R1167 B.n476 B.n0 10.6151
R1168 B.n329 B.n328 10.6151
R1169 B.n328 B.n220 10.6151
R1170 B.n323 B.n220 10.6151
R1171 B.n323 B.n322 10.6151
R1172 B.n322 B.n222 10.6151
R1173 B.n317 B.n222 10.6151
R1174 B.n317 B.n316 10.6151
R1175 B.n316 B.n315 10.6151
R1176 B.n315 B.n224 10.6151
R1177 B.n309 B.n224 10.6151
R1178 B.n309 B.n308 10.6151
R1179 B.n308 B.n307 10.6151
R1180 B.n307 B.n226 10.6151
R1181 B.n301 B.n226 10.6151
R1182 B.n301 B.n300 10.6151
R1183 B.n300 B.n299 10.6151
R1184 B.n295 B.n294 10.6151
R1185 B.n294 B.n232 10.6151
R1186 B.n289 B.n232 10.6151
R1187 B.n289 B.n288 10.6151
R1188 B.n288 B.n287 10.6151
R1189 B.n287 B.n234 10.6151
R1190 B.n281 B.n234 10.6151
R1191 B.n281 B.n280 10.6151
R1192 B.n278 B.n238 10.6151
R1193 B.n272 B.n238 10.6151
R1194 B.n272 B.n271 10.6151
R1195 B.n271 B.n270 10.6151
R1196 B.n270 B.n240 10.6151
R1197 B.n264 B.n240 10.6151
R1198 B.n264 B.n263 10.6151
R1199 B.n263 B.n262 10.6151
R1200 B.n262 B.n242 10.6151
R1201 B.n256 B.n242 10.6151
R1202 B.n256 B.n255 10.6151
R1203 B.n255 B.n254 10.6151
R1204 B.n254 B.n244 10.6151
R1205 B.n248 B.n244 10.6151
R1206 B.n248 B.n247 10.6151
R1207 B.n247 B.n216 10.6151
R1208 B.n335 B.n334 10.6151
R1209 B.n336 B.n335 10.6151
R1210 B.n336 B.n208 10.6151
R1211 B.n346 B.n208 10.6151
R1212 B.n347 B.n346 10.6151
R1213 B.n348 B.n347 10.6151
R1214 B.n348 B.n200 10.6151
R1215 B.n358 B.n200 10.6151
R1216 B.n359 B.n358 10.6151
R1217 B.n360 B.n359 10.6151
R1218 B.n360 B.n192 10.6151
R1219 B.n370 B.n192 10.6151
R1220 B.n371 B.n370 10.6151
R1221 B.n372 B.n371 10.6151
R1222 B.n372 B.n184 10.6151
R1223 B.n382 B.n184 10.6151
R1224 B.n383 B.n382 10.6151
R1225 B.n384 B.n383 10.6151
R1226 B.n384 B.n176 10.6151
R1227 B.n394 B.n176 10.6151
R1228 B.n395 B.n394 10.6151
R1229 B.n396 B.n395 10.6151
R1230 B.n396 B.n168 10.6151
R1231 B.n406 B.n168 10.6151
R1232 B.n407 B.n406 10.6151
R1233 B.n408 B.n407 10.6151
R1234 B.n408 B.n160 10.6151
R1235 B.n418 B.n160 10.6151
R1236 B.n419 B.n418 10.6151
R1237 B.n420 B.n419 10.6151
R1238 B.n420 B.n152 10.6151
R1239 B.n430 B.n152 10.6151
R1240 B.n431 B.n430 10.6151
R1241 B.n432 B.n431 10.6151
R1242 B.n432 B.n144 10.6151
R1243 B.n442 B.n144 10.6151
R1244 B.n443 B.n442 10.6151
R1245 B.n444 B.n443 10.6151
R1246 B.n444 B.n136 10.6151
R1247 B.n454 B.n136 10.6151
R1248 B.n455 B.n454 10.6151
R1249 B.n456 B.n455 10.6151
R1250 B.n456 B.n129 10.6151
R1251 B.n467 B.n129 10.6151
R1252 B.n468 B.n467 10.6151
R1253 B.n470 B.n468 10.6151
R1254 B.n470 B.n469 10.6151
R1255 B.n469 B.n121 10.6151
R1256 B.n481 B.n121 10.6151
R1257 B.n482 B.n481 10.6151
R1258 B.n483 B.n482 10.6151
R1259 B.n484 B.n483 10.6151
R1260 B.n485 B.n484 10.6151
R1261 B.n488 B.n485 10.6151
R1262 B.n489 B.n488 10.6151
R1263 B.n490 B.n489 10.6151
R1264 B.n491 B.n490 10.6151
R1265 B.n493 B.n491 10.6151
R1266 B.n494 B.n493 10.6151
R1267 B.n495 B.n494 10.6151
R1268 B.n496 B.n495 10.6151
R1269 B.n498 B.n496 10.6151
R1270 B.n499 B.n498 10.6151
R1271 B.n500 B.n499 10.6151
R1272 B.n501 B.n500 10.6151
R1273 B.n503 B.n501 10.6151
R1274 B.n504 B.n503 10.6151
R1275 B.n505 B.n504 10.6151
R1276 B.n506 B.n505 10.6151
R1277 B.n508 B.n506 10.6151
R1278 B.n509 B.n508 10.6151
R1279 B.n510 B.n509 10.6151
R1280 B.n511 B.n510 10.6151
R1281 B.n513 B.n511 10.6151
R1282 B.n514 B.n513 10.6151
R1283 B.n515 B.n514 10.6151
R1284 B.n516 B.n515 10.6151
R1285 B.n518 B.n516 10.6151
R1286 B.n519 B.n518 10.6151
R1287 B.n520 B.n519 10.6151
R1288 B.n521 B.n520 10.6151
R1289 B.n523 B.n521 10.6151
R1290 B.n524 B.n523 10.6151
R1291 B.n525 B.n524 10.6151
R1292 B.n526 B.n525 10.6151
R1293 B.n528 B.n526 10.6151
R1294 B.n529 B.n528 10.6151
R1295 B.n530 B.n529 10.6151
R1296 B.n531 B.n530 10.6151
R1297 B.n533 B.n531 10.6151
R1298 B.n534 B.n533 10.6151
R1299 B.n535 B.n534 10.6151
R1300 B.n536 B.n535 10.6151
R1301 B.n538 B.n536 10.6151
R1302 B.n539 B.n538 10.6151
R1303 B.n540 B.n539 10.6151
R1304 B.n541 B.n540 10.6151
R1305 B.n543 B.n541 10.6151
R1306 B.n544 B.n543 10.6151
R1307 B.n545 B.n544 10.6151
R1308 B.n546 B.n545 10.6151
R1309 B.n729 B.n1 10.6151
R1310 B.n729 B.n728 10.6151
R1311 B.n728 B.n727 10.6151
R1312 B.n727 B.n10 10.6151
R1313 B.n721 B.n10 10.6151
R1314 B.n721 B.n720 10.6151
R1315 B.n720 B.n719 10.6151
R1316 B.n719 B.n17 10.6151
R1317 B.n713 B.n17 10.6151
R1318 B.n713 B.n712 10.6151
R1319 B.n712 B.n711 10.6151
R1320 B.n711 B.n25 10.6151
R1321 B.n705 B.n25 10.6151
R1322 B.n705 B.n704 10.6151
R1323 B.n704 B.n703 10.6151
R1324 B.n703 B.n32 10.6151
R1325 B.n697 B.n32 10.6151
R1326 B.n697 B.n696 10.6151
R1327 B.n696 B.n695 10.6151
R1328 B.n695 B.n39 10.6151
R1329 B.n689 B.n39 10.6151
R1330 B.n689 B.n688 10.6151
R1331 B.n688 B.n687 10.6151
R1332 B.n687 B.n46 10.6151
R1333 B.n681 B.n46 10.6151
R1334 B.n681 B.n680 10.6151
R1335 B.n680 B.n679 10.6151
R1336 B.n679 B.n53 10.6151
R1337 B.n673 B.n53 10.6151
R1338 B.n673 B.n672 10.6151
R1339 B.n672 B.n671 10.6151
R1340 B.n671 B.n60 10.6151
R1341 B.n665 B.n60 10.6151
R1342 B.n665 B.n664 10.6151
R1343 B.n664 B.n663 10.6151
R1344 B.n663 B.n67 10.6151
R1345 B.n657 B.n67 10.6151
R1346 B.n657 B.n656 10.6151
R1347 B.n656 B.n655 10.6151
R1348 B.n655 B.n74 10.6151
R1349 B.n649 B.n74 10.6151
R1350 B.n649 B.n648 10.6151
R1351 B.n648 B.n647 10.6151
R1352 B.n647 B.n81 10.6151
R1353 B.n641 B.n81 10.6151
R1354 B.n641 B.n640 10.6151
R1355 B.n640 B.n639 10.6151
R1356 B.n639 B.n88 10.6151
R1357 B.n633 B.n88 10.6151
R1358 B.n632 B.n631 10.6151
R1359 B.n631 B.n95 10.6151
R1360 B.n625 B.n95 10.6151
R1361 B.n625 B.n624 10.6151
R1362 B.n624 B.n623 10.6151
R1363 B.n623 B.n97 10.6151
R1364 B.n617 B.n97 10.6151
R1365 B.n617 B.n616 10.6151
R1366 B.n616 B.n615 10.6151
R1367 B.n615 B.n99 10.6151
R1368 B.n609 B.n99 10.6151
R1369 B.n609 B.n608 10.6151
R1370 B.n608 B.n607 10.6151
R1371 B.n607 B.n101 10.6151
R1372 B.n601 B.n101 10.6151
R1373 B.n601 B.n600 10.6151
R1374 B.n598 B.n105 10.6151
R1375 B.n592 B.n105 10.6151
R1376 B.n592 B.n591 10.6151
R1377 B.n591 B.n590 10.6151
R1378 B.n590 B.n107 10.6151
R1379 B.n584 B.n107 10.6151
R1380 B.n584 B.n583 10.6151
R1381 B.n583 B.n582 10.6151
R1382 B.n578 B.n577 10.6151
R1383 B.n577 B.n113 10.6151
R1384 B.n572 B.n113 10.6151
R1385 B.n572 B.n571 10.6151
R1386 B.n571 B.n570 10.6151
R1387 B.n570 B.n115 10.6151
R1388 B.n564 B.n115 10.6151
R1389 B.n564 B.n563 10.6151
R1390 B.n563 B.n562 10.6151
R1391 B.n562 B.n117 10.6151
R1392 B.n556 B.n117 10.6151
R1393 B.n556 B.n555 10.6151
R1394 B.n555 B.n554 10.6151
R1395 B.n554 B.n119 10.6151
R1396 B.n548 B.n119 10.6151
R1397 B.n548 B.n547 10.6151
R1398 B.n737 B.n0 8.11757
R1399 B.n737 B.n1 8.11757
R1400 B.n295 B.n230 6.5566
R1401 B.n280 B.n279 6.5566
R1402 B.n599 B.n598 6.5566
R1403 B.n582 B.n111 6.5566
R1404 B.n299 B.n230 4.05904
R1405 B.n279 B.n278 4.05904
R1406 B.n600 B.n599 4.05904
R1407 B.n578 B.n111 4.05904
R1408 B.t3 B.n150 2.48778
R1409 B.n700 B.t2 2.48778
R1410 VN.n34 VN.n33 161.3
R1411 VN.n32 VN.n19 161.3
R1412 VN.n31 VN.n30 161.3
R1413 VN.n29 VN.n20 161.3
R1414 VN.n28 VN.n27 161.3
R1415 VN.n26 VN.n21 161.3
R1416 VN.n25 VN.n24 161.3
R1417 VN.n16 VN.n15 161.3
R1418 VN.n14 VN.n1 161.3
R1419 VN.n13 VN.n12 161.3
R1420 VN.n11 VN.n2 161.3
R1421 VN.n10 VN.n9 161.3
R1422 VN.n8 VN.n3 161.3
R1423 VN.n7 VN.n6 161.3
R1424 VN.n17 VN.n0 72.4512
R1425 VN.n35 VN.n18 72.4512
R1426 VN.n5 VN.n4 62.0548
R1427 VN.n23 VN.n22 62.0548
R1428 VN.n23 VN.t4 59.446
R1429 VN.n5 VN.t5 59.446
R1430 VN.n13 VN.n2 45.8354
R1431 VN.n31 VN.n20 45.8354
R1432 VN VN.n35 45.2745
R1433 VN.n9 VN.n2 35.1514
R1434 VN.n27 VN.n20 35.1514
R1435 VN.n4 VN.t3 26.2313
R1436 VN.n0 VN.t2 26.2313
R1437 VN.n22 VN.t1 26.2313
R1438 VN.n18 VN.t0 26.2313
R1439 VN.n8 VN.n7 24.4675
R1440 VN.n9 VN.n8 24.4675
R1441 VN.n14 VN.n13 24.4675
R1442 VN.n15 VN.n14 24.4675
R1443 VN.n27 VN.n26 24.4675
R1444 VN.n26 VN.n25 24.4675
R1445 VN.n33 VN.n32 24.4675
R1446 VN.n32 VN.n31 24.4675
R1447 VN.n15 VN.n0 17.6167
R1448 VN.n33 VN.n18 17.6167
R1449 VN.n7 VN.n4 12.234
R1450 VN.n25 VN.n22 12.234
R1451 VN.n6 VN.n5 4.01738
R1452 VN.n24 VN.n23 4.01738
R1453 VN.n35 VN.n34 0.354971
R1454 VN.n17 VN.n16 0.354971
R1455 VN VN.n17 0.26696
R1456 VN.n34 VN.n19 0.189894
R1457 VN.n30 VN.n19 0.189894
R1458 VN.n30 VN.n29 0.189894
R1459 VN.n29 VN.n28 0.189894
R1460 VN.n28 VN.n21 0.189894
R1461 VN.n24 VN.n21 0.189894
R1462 VN.n6 VN.n3 0.189894
R1463 VN.n10 VN.n3 0.189894
R1464 VN.n11 VN.n10 0.189894
R1465 VN.n12 VN.n11 0.189894
R1466 VN.n12 VN.n1 0.189894
R1467 VN.n16 VN.n1 0.189894
R1468 VDD2.n1 VDD2.t0 84.9309
R1469 VDD2.n2 VDD2.t5 82.6522
R1470 VDD2.n1 VDD2.n0 77.8285
R1471 VDD2 VDD2.n3 77.8258
R1472 VDD2.n2 VDD2.n1 36.9071
R1473 VDD2.n3 VDD2.t4 5.54672
R1474 VDD2.n3 VDD2.t1 5.54672
R1475 VDD2.n0 VDD2.t2 5.54672
R1476 VDD2.n0 VDD2.t3 5.54672
R1477 VDD2 VDD2.n2 2.39274
C0 VP VDD2 0.520557f
C1 VTAIL VP 3.31807f
C2 VN VDD1 0.156155f
C3 VDD1 VDD2 1.67067f
C4 VTAIL VDD1 5.11546f
C5 VN VDD2 2.36565f
C6 VTAIL VN 3.30393f
C7 VP VDD1 2.72739f
C8 VTAIL VDD2 5.17301f
C9 VP VN 6.03175f
C10 VDD2 B 5.008764f
C11 VDD1 B 5.34826f
C12 VTAIL B 4.422054f
C13 VN B 14.15192f
C14 VP B 12.768322f
C15 VDD2.t0 B 0.630864f
C16 VDD2.t2 B 0.06338f
C17 VDD2.t3 B 0.06338f
C18 VDD2.n0 B 0.491974f
C19 VDD2.n1 B 2.37833f
C20 VDD2.t5 B 0.620488f
C21 VDD2.n2 B 2.05285f
C22 VDD2.t4 B 0.06338f
C23 VDD2.t1 B 0.06338f
C24 VDD2.n3 B 0.491948f
C25 VN.t2 B 0.771328f
C26 VN.n0 B 0.413934f
C27 VN.n1 B 0.025926f
C28 VN.n2 B 0.021984f
C29 VN.n3 B 0.025926f
C30 VN.t3 B 0.771328f
C31 VN.n4 B 0.393684f
C32 VN.t5 B 1.04816f
C33 VN.n5 B 0.385365f
C34 VN.n6 B 0.3025f
C35 VN.n7 B 0.036391f
C36 VN.n8 B 0.048319f
C37 VN.n9 B 0.052379f
C38 VN.n10 B 0.025926f
C39 VN.n11 B 0.025926f
C40 VN.n12 B 0.025926f
C41 VN.n13 B 0.049653f
C42 VN.n14 B 0.048319f
C43 VN.n15 B 0.041639f
C44 VN.n16 B 0.041843f
C45 VN.n17 B 0.059281f
C46 VN.t0 B 0.771328f
C47 VN.n18 B 0.413934f
C48 VN.n19 B 0.025926f
C49 VN.n20 B 0.021984f
C50 VN.n21 B 0.025926f
C51 VN.t1 B 0.771328f
C52 VN.n22 B 0.393684f
C53 VN.t4 B 1.04816f
C54 VN.n23 B 0.385365f
C55 VN.n24 B 0.3025f
C56 VN.n25 B 0.036391f
C57 VN.n26 B 0.048319f
C58 VN.n27 B 0.052379f
C59 VN.n28 B 0.025926f
C60 VN.n29 B 0.025926f
C61 VN.n30 B 0.025926f
C62 VN.n31 B 0.049653f
C63 VN.n32 B 0.048319f
C64 VN.n33 B 0.041639f
C65 VN.n34 B 0.041843f
C66 VN.n35 B 1.27599f
C67 VDD1.t2 B 0.641214f
C68 VDD1.t1 B 0.640473f
C69 VDD1.t3 B 0.064346f
C70 VDD1.t5 B 0.064346f
C71 VDD1.n0 B 0.499467f
C72 VDD1.n1 B 2.53555f
C73 VDD1.t4 B 0.064346f
C74 VDD1.t0 B 0.064346f
C75 VDD1.n2 B 0.495131f
C76 VDD1.n3 B 2.11249f
C77 VTAIL.t11 B 0.088606f
C78 VTAIL.t2 B 0.088606f
C79 VTAIL.n0 B 0.616888f
C80 VTAIL.n1 B 0.553096f
C81 VTAIL.t9 B 0.793813f
C82 VTAIL.n2 B 0.848151f
C83 VTAIL.t5 B 0.088606f
C84 VTAIL.t6 B 0.088606f
C85 VTAIL.n3 B 0.616888f
C86 VTAIL.n4 B 1.94641f
C87 VTAIL.t4 B 0.088606f
C88 VTAIL.t3 B 0.088606f
C89 VTAIL.n5 B 0.616891f
C90 VTAIL.n6 B 1.94641f
C91 VTAIL.t1 B 0.793818f
C92 VTAIL.n7 B 0.848146f
C93 VTAIL.t7 B 0.088606f
C94 VTAIL.t10 B 0.088606f
C95 VTAIL.n8 B 0.616891f
C96 VTAIL.n9 B 0.78342f
C97 VTAIL.t8 B 0.793813f
C98 VTAIL.n10 B 1.69619f
C99 VTAIL.t0 B 0.793813f
C100 VTAIL.n11 B 1.61156f
C101 VP.t0 B 0.793578f
C102 VP.n0 B 0.425874f
C103 VP.n1 B 0.026673f
C104 VP.n2 B 0.022619f
C105 VP.n3 B 0.026673f
C106 VP.t2 B 0.793578f
C107 VP.n4 B 0.316312f
C108 VP.n5 B 0.026673f
C109 VP.n6 B 0.022619f
C110 VP.n7 B 0.026673f
C111 VP.t4 B 0.793578f
C112 VP.n8 B 0.425874f
C113 VP.t5 B 0.793578f
C114 VP.n9 B 0.425874f
C115 VP.n10 B 0.026673f
C116 VP.n11 B 0.022619f
C117 VP.n12 B 0.026673f
C118 VP.t1 B 0.793578f
C119 VP.n13 B 0.40504f
C120 VP.t3 B 1.07839f
C121 VP.n14 B 0.396482f
C122 VP.n15 B 0.311226f
C123 VP.n16 B 0.037441f
C124 VP.n17 B 0.049712f
C125 VP.n18 B 0.05389f
C126 VP.n19 B 0.026673f
C127 VP.n20 B 0.026673f
C128 VP.n21 B 0.026673f
C129 VP.n22 B 0.051085f
C130 VP.n23 B 0.049712f
C131 VP.n24 B 0.04284f
C132 VP.n25 B 0.04305f
C133 VP.n26 B 1.30149f
C134 VP.n27 B 1.32274f
C135 VP.n28 B 0.04305f
C136 VP.n29 B 0.04284f
C137 VP.n30 B 0.049712f
C138 VP.n31 B 0.051085f
C139 VP.n32 B 0.026673f
C140 VP.n33 B 0.026673f
C141 VP.n34 B 0.026673f
C142 VP.n35 B 0.05389f
C143 VP.n36 B 0.049712f
C144 VP.n37 B 0.037441f
C145 VP.n38 B 0.026673f
C146 VP.n39 B 0.026673f
C147 VP.n40 B 0.037441f
C148 VP.n41 B 0.049712f
C149 VP.n42 B 0.05389f
C150 VP.n43 B 0.026673f
C151 VP.n44 B 0.026673f
C152 VP.n45 B 0.026673f
C153 VP.n46 B 0.051085f
C154 VP.n47 B 0.049712f
C155 VP.n48 B 0.04284f
C156 VP.n49 B 0.04305f
C157 VP.n50 B 0.060991f
.ends

