* NGSPICE file created from diff_pair_sample_1768.ext - technology: sky130A

.subckt diff_pair_sample_1768 VTAIL VN VP B VDD2 VDD1
X0 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=7.5231 pd=39.36 as=0 ps=0 w=19.29 l=2.3
X1 VDD1.t5 VP.t0 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=3.18285 pd=19.62 as=7.5231 ps=39.36 w=19.29 l=2.3
X2 VTAIL.t10 VP.t1 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=3.18285 pd=19.62 as=3.18285 ps=19.62 w=19.29 l=2.3
X3 VDD1.t3 VP.t2 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=7.5231 pd=39.36 as=3.18285 ps=19.62 w=19.29 l=2.3
X4 VTAIL.t5 VP.t3 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.18285 pd=19.62 as=3.18285 ps=19.62 w=19.29 l=2.3
X5 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=7.5231 pd=39.36 as=0 ps=0 w=19.29 l=2.3
X6 B.t11 B.t9 B.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=7.5231 pd=39.36 as=0 ps=0 w=19.29 l=2.3
X7 VDD2.t5 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.18285 pd=19.62 as=7.5231 ps=39.36 w=19.29 l=2.3
X8 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=7.5231 pd=39.36 as=0 ps=0 w=19.29 l=2.3
X9 VTAIL.t2 VN.t1 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=3.18285 pd=19.62 as=3.18285 ps=19.62 w=19.29 l=2.3
X10 VDD2.t3 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.5231 pd=39.36 as=3.18285 ps=19.62 w=19.29 l=2.3
X11 VDD2.t2 VN.t3 VTAIL.t11 B.t19 sky130_fd_pr__nfet_01v8 ad=7.5231 pd=39.36 as=3.18285 ps=19.62 w=19.29 l=2.3
X12 VDD1.t1 VP.t4 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=3.18285 pd=19.62 as=7.5231 ps=39.36 w=19.29 l=2.3
X13 VTAIL.t0 VN.t4 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=3.18285 pd=19.62 as=3.18285 ps=19.62 w=19.29 l=2.3
X14 VDD2.t0 VN.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.18285 pd=19.62 as=7.5231 ps=39.36 w=19.29 l=2.3
X15 VDD1.t0 VP.t5 VTAIL.t9 B.t19 sky130_fd_pr__nfet_01v8 ad=7.5231 pd=39.36 as=3.18285 ps=19.62 w=19.29 l=2.3
R0 B.n1002 B.n1001 585
R1 B.n413 B.n141 585
R2 B.n412 B.n411 585
R3 B.n410 B.n409 585
R4 B.n408 B.n407 585
R5 B.n406 B.n405 585
R6 B.n404 B.n403 585
R7 B.n402 B.n401 585
R8 B.n400 B.n399 585
R9 B.n398 B.n397 585
R10 B.n396 B.n395 585
R11 B.n394 B.n393 585
R12 B.n392 B.n391 585
R13 B.n390 B.n389 585
R14 B.n388 B.n387 585
R15 B.n386 B.n385 585
R16 B.n384 B.n383 585
R17 B.n382 B.n381 585
R18 B.n380 B.n379 585
R19 B.n378 B.n377 585
R20 B.n376 B.n375 585
R21 B.n374 B.n373 585
R22 B.n372 B.n371 585
R23 B.n370 B.n369 585
R24 B.n368 B.n367 585
R25 B.n366 B.n365 585
R26 B.n364 B.n363 585
R27 B.n362 B.n361 585
R28 B.n360 B.n359 585
R29 B.n358 B.n357 585
R30 B.n356 B.n355 585
R31 B.n354 B.n353 585
R32 B.n352 B.n351 585
R33 B.n350 B.n349 585
R34 B.n348 B.n347 585
R35 B.n346 B.n345 585
R36 B.n344 B.n343 585
R37 B.n342 B.n341 585
R38 B.n340 B.n339 585
R39 B.n338 B.n337 585
R40 B.n336 B.n335 585
R41 B.n334 B.n333 585
R42 B.n332 B.n331 585
R43 B.n330 B.n329 585
R44 B.n328 B.n327 585
R45 B.n326 B.n325 585
R46 B.n324 B.n323 585
R47 B.n322 B.n321 585
R48 B.n320 B.n319 585
R49 B.n318 B.n317 585
R50 B.n316 B.n315 585
R51 B.n314 B.n313 585
R52 B.n312 B.n311 585
R53 B.n310 B.n309 585
R54 B.n308 B.n307 585
R55 B.n306 B.n305 585
R56 B.n304 B.n303 585
R57 B.n302 B.n301 585
R58 B.n300 B.n299 585
R59 B.n298 B.n297 585
R60 B.n296 B.n295 585
R61 B.n294 B.n293 585
R62 B.n292 B.n291 585
R63 B.n289 B.n288 585
R64 B.n287 B.n286 585
R65 B.n285 B.n284 585
R66 B.n283 B.n282 585
R67 B.n281 B.n280 585
R68 B.n279 B.n278 585
R69 B.n277 B.n276 585
R70 B.n275 B.n274 585
R71 B.n273 B.n272 585
R72 B.n271 B.n270 585
R73 B.n268 B.n267 585
R74 B.n266 B.n265 585
R75 B.n264 B.n263 585
R76 B.n262 B.n261 585
R77 B.n260 B.n259 585
R78 B.n258 B.n257 585
R79 B.n256 B.n255 585
R80 B.n254 B.n253 585
R81 B.n252 B.n251 585
R82 B.n250 B.n249 585
R83 B.n248 B.n247 585
R84 B.n246 B.n245 585
R85 B.n244 B.n243 585
R86 B.n242 B.n241 585
R87 B.n240 B.n239 585
R88 B.n238 B.n237 585
R89 B.n236 B.n235 585
R90 B.n234 B.n233 585
R91 B.n232 B.n231 585
R92 B.n230 B.n229 585
R93 B.n228 B.n227 585
R94 B.n226 B.n225 585
R95 B.n224 B.n223 585
R96 B.n222 B.n221 585
R97 B.n220 B.n219 585
R98 B.n218 B.n217 585
R99 B.n216 B.n215 585
R100 B.n214 B.n213 585
R101 B.n212 B.n211 585
R102 B.n210 B.n209 585
R103 B.n208 B.n207 585
R104 B.n206 B.n205 585
R105 B.n204 B.n203 585
R106 B.n202 B.n201 585
R107 B.n200 B.n199 585
R108 B.n198 B.n197 585
R109 B.n196 B.n195 585
R110 B.n194 B.n193 585
R111 B.n192 B.n191 585
R112 B.n190 B.n189 585
R113 B.n188 B.n187 585
R114 B.n186 B.n185 585
R115 B.n184 B.n183 585
R116 B.n182 B.n181 585
R117 B.n180 B.n179 585
R118 B.n178 B.n177 585
R119 B.n176 B.n175 585
R120 B.n174 B.n173 585
R121 B.n172 B.n171 585
R122 B.n170 B.n169 585
R123 B.n168 B.n167 585
R124 B.n166 B.n165 585
R125 B.n164 B.n163 585
R126 B.n162 B.n161 585
R127 B.n160 B.n159 585
R128 B.n158 B.n157 585
R129 B.n156 B.n155 585
R130 B.n154 B.n153 585
R131 B.n152 B.n151 585
R132 B.n150 B.n149 585
R133 B.n148 B.n147 585
R134 B.n74 B.n73 585
R135 B.n1007 B.n1006 585
R136 B.n1000 B.n142 585
R137 B.n142 B.n71 585
R138 B.n999 B.n70 585
R139 B.n1011 B.n70 585
R140 B.n998 B.n69 585
R141 B.n1012 B.n69 585
R142 B.n997 B.n68 585
R143 B.n1013 B.n68 585
R144 B.n996 B.n995 585
R145 B.n995 B.n64 585
R146 B.n994 B.n63 585
R147 B.n1019 B.n63 585
R148 B.n993 B.n62 585
R149 B.n1020 B.n62 585
R150 B.n992 B.n61 585
R151 B.n1021 B.n61 585
R152 B.n991 B.n990 585
R153 B.n990 B.n57 585
R154 B.n989 B.n56 585
R155 B.n1027 B.n56 585
R156 B.n988 B.n55 585
R157 B.n1028 B.n55 585
R158 B.n987 B.n54 585
R159 B.n1029 B.n54 585
R160 B.n986 B.n985 585
R161 B.n985 B.n50 585
R162 B.n984 B.n49 585
R163 B.n1035 B.n49 585
R164 B.n983 B.n48 585
R165 B.n1036 B.n48 585
R166 B.n982 B.n47 585
R167 B.n1037 B.n47 585
R168 B.n981 B.n980 585
R169 B.n980 B.n43 585
R170 B.n979 B.n42 585
R171 B.n1043 B.n42 585
R172 B.n978 B.n41 585
R173 B.n1044 B.n41 585
R174 B.n977 B.n40 585
R175 B.n1045 B.n40 585
R176 B.n976 B.n975 585
R177 B.n975 B.n36 585
R178 B.n974 B.n35 585
R179 B.n1051 B.n35 585
R180 B.n973 B.n34 585
R181 B.n1052 B.n34 585
R182 B.n972 B.n33 585
R183 B.n1053 B.n33 585
R184 B.n971 B.n970 585
R185 B.n970 B.n29 585
R186 B.n969 B.n28 585
R187 B.n1059 B.n28 585
R188 B.n968 B.n27 585
R189 B.n1060 B.n27 585
R190 B.n967 B.n26 585
R191 B.n1061 B.n26 585
R192 B.n966 B.n965 585
R193 B.n965 B.n22 585
R194 B.n964 B.n21 585
R195 B.n1067 B.n21 585
R196 B.n963 B.n20 585
R197 B.n1068 B.n20 585
R198 B.n962 B.n19 585
R199 B.n1069 B.n19 585
R200 B.n961 B.n960 585
R201 B.n960 B.n15 585
R202 B.n959 B.n14 585
R203 B.n1075 B.n14 585
R204 B.n958 B.n13 585
R205 B.n1076 B.n13 585
R206 B.n957 B.n12 585
R207 B.n1077 B.n12 585
R208 B.n956 B.n955 585
R209 B.n955 B.n8 585
R210 B.n954 B.n7 585
R211 B.n1083 B.n7 585
R212 B.n953 B.n6 585
R213 B.n1084 B.n6 585
R214 B.n952 B.n5 585
R215 B.n1085 B.n5 585
R216 B.n951 B.n950 585
R217 B.n950 B.n4 585
R218 B.n949 B.n414 585
R219 B.n949 B.n948 585
R220 B.n939 B.n415 585
R221 B.n416 B.n415 585
R222 B.n941 B.n940 585
R223 B.n942 B.n941 585
R224 B.n938 B.n421 585
R225 B.n421 B.n420 585
R226 B.n937 B.n936 585
R227 B.n936 B.n935 585
R228 B.n423 B.n422 585
R229 B.n424 B.n423 585
R230 B.n928 B.n927 585
R231 B.n929 B.n928 585
R232 B.n926 B.n429 585
R233 B.n429 B.n428 585
R234 B.n925 B.n924 585
R235 B.n924 B.n923 585
R236 B.n431 B.n430 585
R237 B.n432 B.n431 585
R238 B.n916 B.n915 585
R239 B.n917 B.n916 585
R240 B.n914 B.n437 585
R241 B.n437 B.n436 585
R242 B.n913 B.n912 585
R243 B.n912 B.n911 585
R244 B.n439 B.n438 585
R245 B.n440 B.n439 585
R246 B.n904 B.n903 585
R247 B.n905 B.n904 585
R248 B.n902 B.n445 585
R249 B.n445 B.n444 585
R250 B.n901 B.n900 585
R251 B.n900 B.n899 585
R252 B.n447 B.n446 585
R253 B.n448 B.n447 585
R254 B.n892 B.n891 585
R255 B.n893 B.n892 585
R256 B.n890 B.n452 585
R257 B.n456 B.n452 585
R258 B.n889 B.n888 585
R259 B.n888 B.n887 585
R260 B.n454 B.n453 585
R261 B.n455 B.n454 585
R262 B.n880 B.n879 585
R263 B.n881 B.n880 585
R264 B.n878 B.n461 585
R265 B.n461 B.n460 585
R266 B.n877 B.n876 585
R267 B.n876 B.n875 585
R268 B.n463 B.n462 585
R269 B.n464 B.n463 585
R270 B.n868 B.n867 585
R271 B.n869 B.n868 585
R272 B.n866 B.n469 585
R273 B.n469 B.n468 585
R274 B.n865 B.n864 585
R275 B.n864 B.n863 585
R276 B.n471 B.n470 585
R277 B.n472 B.n471 585
R278 B.n856 B.n855 585
R279 B.n857 B.n856 585
R280 B.n854 B.n477 585
R281 B.n477 B.n476 585
R282 B.n853 B.n852 585
R283 B.n852 B.n851 585
R284 B.n479 B.n478 585
R285 B.n480 B.n479 585
R286 B.n844 B.n843 585
R287 B.n845 B.n844 585
R288 B.n842 B.n485 585
R289 B.n485 B.n484 585
R290 B.n841 B.n840 585
R291 B.n840 B.n839 585
R292 B.n487 B.n486 585
R293 B.n488 B.n487 585
R294 B.n835 B.n834 585
R295 B.n491 B.n490 585
R296 B.n831 B.n830 585
R297 B.n832 B.n831 585
R298 B.n829 B.n559 585
R299 B.n828 B.n827 585
R300 B.n826 B.n825 585
R301 B.n824 B.n823 585
R302 B.n822 B.n821 585
R303 B.n820 B.n819 585
R304 B.n818 B.n817 585
R305 B.n816 B.n815 585
R306 B.n814 B.n813 585
R307 B.n812 B.n811 585
R308 B.n810 B.n809 585
R309 B.n808 B.n807 585
R310 B.n806 B.n805 585
R311 B.n804 B.n803 585
R312 B.n802 B.n801 585
R313 B.n800 B.n799 585
R314 B.n798 B.n797 585
R315 B.n796 B.n795 585
R316 B.n794 B.n793 585
R317 B.n792 B.n791 585
R318 B.n790 B.n789 585
R319 B.n788 B.n787 585
R320 B.n786 B.n785 585
R321 B.n784 B.n783 585
R322 B.n782 B.n781 585
R323 B.n780 B.n779 585
R324 B.n778 B.n777 585
R325 B.n776 B.n775 585
R326 B.n774 B.n773 585
R327 B.n772 B.n771 585
R328 B.n770 B.n769 585
R329 B.n768 B.n767 585
R330 B.n766 B.n765 585
R331 B.n764 B.n763 585
R332 B.n762 B.n761 585
R333 B.n760 B.n759 585
R334 B.n758 B.n757 585
R335 B.n756 B.n755 585
R336 B.n754 B.n753 585
R337 B.n752 B.n751 585
R338 B.n750 B.n749 585
R339 B.n748 B.n747 585
R340 B.n746 B.n745 585
R341 B.n744 B.n743 585
R342 B.n742 B.n741 585
R343 B.n740 B.n739 585
R344 B.n738 B.n737 585
R345 B.n736 B.n735 585
R346 B.n734 B.n733 585
R347 B.n732 B.n731 585
R348 B.n730 B.n729 585
R349 B.n728 B.n727 585
R350 B.n726 B.n725 585
R351 B.n724 B.n723 585
R352 B.n722 B.n721 585
R353 B.n720 B.n719 585
R354 B.n718 B.n717 585
R355 B.n716 B.n715 585
R356 B.n714 B.n713 585
R357 B.n712 B.n711 585
R358 B.n710 B.n709 585
R359 B.n708 B.n707 585
R360 B.n706 B.n705 585
R361 B.n704 B.n703 585
R362 B.n702 B.n701 585
R363 B.n700 B.n699 585
R364 B.n698 B.n697 585
R365 B.n696 B.n695 585
R366 B.n694 B.n693 585
R367 B.n692 B.n691 585
R368 B.n690 B.n689 585
R369 B.n688 B.n687 585
R370 B.n686 B.n685 585
R371 B.n684 B.n683 585
R372 B.n682 B.n681 585
R373 B.n680 B.n679 585
R374 B.n678 B.n677 585
R375 B.n676 B.n675 585
R376 B.n674 B.n673 585
R377 B.n672 B.n671 585
R378 B.n670 B.n669 585
R379 B.n668 B.n667 585
R380 B.n666 B.n665 585
R381 B.n664 B.n663 585
R382 B.n662 B.n661 585
R383 B.n660 B.n659 585
R384 B.n658 B.n657 585
R385 B.n656 B.n655 585
R386 B.n654 B.n653 585
R387 B.n652 B.n651 585
R388 B.n650 B.n649 585
R389 B.n648 B.n647 585
R390 B.n646 B.n645 585
R391 B.n644 B.n643 585
R392 B.n642 B.n641 585
R393 B.n640 B.n639 585
R394 B.n638 B.n637 585
R395 B.n636 B.n635 585
R396 B.n634 B.n633 585
R397 B.n632 B.n631 585
R398 B.n630 B.n629 585
R399 B.n628 B.n627 585
R400 B.n626 B.n625 585
R401 B.n624 B.n623 585
R402 B.n622 B.n621 585
R403 B.n620 B.n619 585
R404 B.n618 B.n617 585
R405 B.n616 B.n615 585
R406 B.n614 B.n613 585
R407 B.n612 B.n611 585
R408 B.n610 B.n609 585
R409 B.n608 B.n607 585
R410 B.n606 B.n605 585
R411 B.n604 B.n603 585
R412 B.n602 B.n601 585
R413 B.n600 B.n599 585
R414 B.n598 B.n597 585
R415 B.n596 B.n595 585
R416 B.n594 B.n593 585
R417 B.n592 B.n591 585
R418 B.n590 B.n589 585
R419 B.n588 B.n587 585
R420 B.n586 B.n585 585
R421 B.n584 B.n583 585
R422 B.n582 B.n581 585
R423 B.n580 B.n579 585
R424 B.n578 B.n577 585
R425 B.n576 B.n575 585
R426 B.n574 B.n573 585
R427 B.n572 B.n571 585
R428 B.n570 B.n569 585
R429 B.n568 B.n567 585
R430 B.n566 B.n558 585
R431 B.n832 B.n558 585
R432 B.n836 B.n489 585
R433 B.n489 B.n488 585
R434 B.n838 B.n837 585
R435 B.n839 B.n838 585
R436 B.n483 B.n482 585
R437 B.n484 B.n483 585
R438 B.n847 B.n846 585
R439 B.n846 B.n845 585
R440 B.n848 B.n481 585
R441 B.n481 B.n480 585
R442 B.n850 B.n849 585
R443 B.n851 B.n850 585
R444 B.n475 B.n474 585
R445 B.n476 B.n475 585
R446 B.n859 B.n858 585
R447 B.n858 B.n857 585
R448 B.n860 B.n473 585
R449 B.n473 B.n472 585
R450 B.n862 B.n861 585
R451 B.n863 B.n862 585
R452 B.n467 B.n466 585
R453 B.n468 B.n467 585
R454 B.n871 B.n870 585
R455 B.n870 B.n869 585
R456 B.n872 B.n465 585
R457 B.n465 B.n464 585
R458 B.n874 B.n873 585
R459 B.n875 B.n874 585
R460 B.n459 B.n458 585
R461 B.n460 B.n459 585
R462 B.n883 B.n882 585
R463 B.n882 B.n881 585
R464 B.n884 B.n457 585
R465 B.n457 B.n455 585
R466 B.n886 B.n885 585
R467 B.n887 B.n886 585
R468 B.n451 B.n450 585
R469 B.n456 B.n451 585
R470 B.n895 B.n894 585
R471 B.n894 B.n893 585
R472 B.n896 B.n449 585
R473 B.n449 B.n448 585
R474 B.n898 B.n897 585
R475 B.n899 B.n898 585
R476 B.n443 B.n442 585
R477 B.n444 B.n443 585
R478 B.n907 B.n906 585
R479 B.n906 B.n905 585
R480 B.n908 B.n441 585
R481 B.n441 B.n440 585
R482 B.n910 B.n909 585
R483 B.n911 B.n910 585
R484 B.n435 B.n434 585
R485 B.n436 B.n435 585
R486 B.n919 B.n918 585
R487 B.n918 B.n917 585
R488 B.n920 B.n433 585
R489 B.n433 B.n432 585
R490 B.n922 B.n921 585
R491 B.n923 B.n922 585
R492 B.n427 B.n426 585
R493 B.n428 B.n427 585
R494 B.n931 B.n930 585
R495 B.n930 B.n929 585
R496 B.n932 B.n425 585
R497 B.n425 B.n424 585
R498 B.n934 B.n933 585
R499 B.n935 B.n934 585
R500 B.n419 B.n418 585
R501 B.n420 B.n419 585
R502 B.n944 B.n943 585
R503 B.n943 B.n942 585
R504 B.n945 B.n417 585
R505 B.n417 B.n416 585
R506 B.n947 B.n946 585
R507 B.n948 B.n947 585
R508 B.n2 B.n0 585
R509 B.n4 B.n2 585
R510 B.n3 B.n1 585
R511 B.n1084 B.n3 585
R512 B.n1082 B.n1081 585
R513 B.n1083 B.n1082 585
R514 B.n1080 B.n9 585
R515 B.n9 B.n8 585
R516 B.n1079 B.n1078 585
R517 B.n1078 B.n1077 585
R518 B.n11 B.n10 585
R519 B.n1076 B.n11 585
R520 B.n1074 B.n1073 585
R521 B.n1075 B.n1074 585
R522 B.n1072 B.n16 585
R523 B.n16 B.n15 585
R524 B.n1071 B.n1070 585
R525 B.n1070 B.n1069 585
R526 B.n18 B.n17 585
R527 B.n1068 B.n18 585
R528 B.n1066 B.n1065 585
R529 B.n1067 B.n1066 585
R530 B.n1064 B.n23 585
R531 B.n23 B.n22 585
R532 B.n1063 B.n1062 585
R533 B.n1062 B.n1061 585
R534 B.n25 B.n24 585
R535 B.n1060 B.n25 585
R536 B.n1058 B.n1057 585
R537 B.n1059 B.n1058 585
R538 B.n1056 B.n30 585
R539 B.n30 B.n29 585
R540 B.n1055 B.n1054 585
R541 B.n1054 B.n1053 585
R542 B.n32 B.n31 585
R543 B.n1052 B.n32 585
R544 B.n1050 B.n1049 585
R545 B.n1051 B.n1050 585
R546 B.n1048 B.n37 585
R547 B.n37 B.n36 585
R548 B.n1047 B.n1046 585
R549 B.n1046 B.n1045 585
R550 B.n39 B.n38 585
R551 B.n1044 B.n39 585
R552 B.n1042 B.n1041 585
R553 B.n1043 B.n1042 585
R554 B.n1040 B.n44 585
R555 B.n44 B.n43 585
R556 B.n1039 B.n1038 585
R557 B.n1038 B.n1037 585
R558 B.n46 B.n45 585
R559 B.n1036 B.n46 585
R560 B.n1034 B.n1033 585
R561 B.n1035 B.n1034 585
R562 B.n1032 B.n51 585
R563 B.n51 B.n50 585
R564 B.n1031 B.n1030 585
R565 B.n1030 B.n1029 585
R566 B.n53 B.n52 585
R567 B.n1028 B.n53 585
R568 B.n1026 B.n1025 585
R569 B.n1027 B.n1026 585
R570 B.n1024 B.n58 585
R571 B.n58 B.n57 585
R572 B.n1023 B.n1022 585
R573 B.n1022 B.n1021 585
R574 B.n60 B.n59 585
R575 B.n1020 B.n60 585
R576 B.n1018 B.n1017 585
R577 B.n1019 B.n1018 585
R578 B.n1016 B.n65 585
R579 B.n65 B.n64 585
R580 B.n1015 B.n1014 585
R581 B.n1014 B.n1013 585
R582 B.n67 B.n66 585
R583 B.n1012 B.n67 585
R584 B.n1010 B.n1009 585
R585 B.n1011 B.n1010 585
R586 B.n1008 B.n72 585
R587 B.n72 B.n71 585
R588 B.n1087 B.n1086 585
R589 B.n1086 B.n1085 585
R590 B.n834 B.n489 482.89
R591 B.n1006 B.n72 482.89
R592 B.n558 B.n487 482.89
R593 B.n1002 B.n142 482.89
R594 B.n563 B.t9 409.671
R595 B.n560 B.t5 409.671
R596 B.n145 B.t12 409.671
R597 B.n143 B.t16 409.671
R598 B.n1004 B.n1003 256.663
R599 B.n1004 B.n140 256.663
R600 B.n1004 B.n139 256.663
R601 B.n1004 B.n138 256.663
R602 B.n1004 B.n137 256.663
R603 B.n1004 B.n136 256.663
R604 B.n1004 B.n135 256.663
R605 B.n1004 B.n134 256.663
R606 B.n1004 B.n133 256.663
R607 B.n1004 B.n132 256.663
R608 B.n1004 B.n131 256.663
R609 B.n1004 B.n130 256.663
R610 B.n1004 B.n129 256.663
R611 B.n1004 B.n128 256.663
R612 B.n1004 B.n127 256.663
R613 B.n1004 B.n126 256.663
R614 B.n1004 B.n125 256.663
R615 B.n1004 B.n124 256.663
R616 B.n1004 B.n123 256.663
R617 B.n1004 B.n122 256.663
R618 B.n1004 B.n121 256.663
R619 B.n1004 B.n120 256.663
R620 B.n1004 B.n119 256.663
R621 B.n1004 B.n118 256.663
R622 B.n1004 B.n117 256.663
R623 B.n1004 B.n116 256.663
R624 B.n1004 B.n115 256.663
R625 B.n1004 B.n114 256.663
R626 B.n1004 B.n113 256.663
R627 B.n1004 B.n112 256.663
R628 B.n1004 B.n111 256.663
R629 B.n1004 B.n110 256.663
R630 B.n1004 B.n109 256.663
R631 B.n1004 B.n108 256.663
R632 B.n1004 B.n107 256.663
R633 B.n1004 B.n106 256.663
R634 B.n1004 B.n105 256.663
R635 B.n1004 B.n104 256.663
R636 B.n1004 B.n103 256.663
R637 B.n1004 B.n102 256.663
R638 B.n1004 B.n101 256.663
R639 B.n1004 B.n100 256.663
R640 B.n1004 B.n99 256.663
R641 B.n1004 B.n98 256.663
R642 B.n1004 B.n97 256.663
R643 B.n1004 B.n96 256.663
R644 B.n1004 B.n95 256.663
R645 B.n1004 B.n94 256.663
R646 B.n1004 B.n93 256.663
R647 B.n1004 B.n92 256.663
R648 B.n1004 B.n91 256.663
R649 B.n1004 B.n90 256.663
R650 B.n1004 B.n89 256.663
R651 B.n1004 B.n88 256.663
R652 B.n1004 B.n87 256.663
R653 B.n1004 B.n86 256.663
R654 B.n1004 B.n85 256.663
R655 B.n1004 B.n84 256.663
R656 B.n1004 B.n83 256.663
R657 B.n1004 B.n82 256.663
R658 B.n1004 B.n81 256.663
R659 B.n1004 B.n80 256.663
R660 B.n1004 B.n79 256.663
R661 B.n1004 B.n78 256.663
R662 B.n1004 B.n77 256.663
R663 B.n1004 B.n76 256.663
R664 B.n1004 B.n75 256.663
R665 B.n1005 B.n1004 256.663
R666 B.n833 B.n832 256.663
R667 B.n832 B.n492 256.663
R668 B.n832 B.n493 256.663
R669 B.n832 B.n494 256.663
R670 B.n832 B.n495 256.663
R671 B.n832 B.n496 256.663
R672 B.n832 B.n497 256.663
R673 B.n832 B.n498 256.663
R674 B.n832 B.n499 256.663
R675 B.n832 B.n500 256.663
R676 B.n832 B.n501 256.663
R677 B.n832 B.n502 256.663
R678 B.n832 B.n503 256.663
R679 B.n832 B.n504 256.663
R680 B.n832 B.n505 256.663
R681 B.n832 B.n506 256.663
R682 B.n832 B.n507 256.663
R683 B.n832 B.n508 256.663
R684 B.n832 B.n509 256.663
R685 B.n832 B.n510 256.663
R686 B.n832 B.n511 256.663
R687 B.n832 B.n512 256.663
R688 B.n832 B.n513 256.663
R689 B.n832 B.n514 256.663
R690 B.n832 B.n515 256.663
R691 B.n832 B.n516 256.663
R692 B.n832 B.n517 256.663
R693 B.n832 B.n518 256.663
R694 B.n832 B.n519 256.663
R695 B.n832 B.n520 256.663
R696 B.n832 B.n521 256.663
R697 B.n832 B.n522 256.663
R698 B.n832 B.n523 256.663
R699 B.n832 B.n524 256.663
R700 B.n832 B.n525 256.663
R701 B.n832 B.n526 256.663
R702 B.n832 B.n527 256.663
R703 B.n832 B.n528 256.663
R704 B.n832 B.n529 256.663
R705 B.n832 B.n530 256.663
R706 B.n832 B.n531 256.663
R707 B.n832 B.n532 256.663
R708 B.n832 B.n533 256.663
R709 B.n832 B.n534 256.663
R710 B.n832 B.n535 256.663
R711 B.n832 B.n536 256.663
R712 B.n832 B.n537 256.663
R713 B.n832 B.n538 256.663
R714 B.n832 B.n539 256.663
R715 B.n832 B.n540 256.663
R716 B.n832 B.n541 256.663
R717 B.n832 B.n542 256.663
R718 B.n832 B.n543 256.663
R719 B.n832 B.n544 256.663
R720 B.n832 B.n545 256.663
R721 B.n832 B.n546 256.663
R722 B.n832 B.n547 256.663
R723 B.n832 B.n548 256.663
R724 B.n832 B.n549 256.663
R725 B.n832 B.n550 256.663
R726 B.n832 B.n551 256.663
R727 B.n832 B.n552 256.663
R728 B.n832 B.n553 256.663
R729 B.n832 B.n554 256.663
R730 B.n832 B.n555 256.663
R731 B.n832 B.n556 256.663
R732 B.n832 B.n557 256.663
R733 B.n838 B.n489 163.367
R734 B.n838 B.n483 163.367
R735 B.n846 B.n483 163.367
R736 B.n846 B.n481 163.367
R737 B.n850 B.n481 163.367
R738 B.n850 B.n475 163.367
R739 B.n858 B.n475 163.367
R740 B.n858 B.n473 163.367
R741 B.n862 B.n473 163.367
R742 B.n862 B.n467 163.367
R743 B.n870 B.n467 163.367
R744 B.n870 B.n465 163.367
R745 B.n874 B.n465 163.367
R746 B.n874 B.n459 163.367
R747 B.n882 B.n459 163.367
R748 B.n882 B.n457 163.367
R749 B.n886 B.n457 163.367
R750 B.n886 B.n451 163.367
R751 B.n894 B.n451 163.367
R752 B.n894 B.n449 163.367
R753 B.n898 B.n449 163.367
R754 B.n898 B.n443 163.367
R755 B.n906 B.n443 163.367
R756 B.n906 B.n441 163.367
R757 B.n910 B.n441 163.367
R758 B.n910 B.n435 163.367
R759 B.n918 B.n435 163.367
R760 B.n918 B.n433 163.367
R761 B.n922 B.n433 163.367
R762 B.n922 B.n427 163.367
R763 B.n930 B.n427 163.367
R764 B.n930 B.n425 163.367
R765 B.n934 B.n425 163.367
R766 B.n934 B.n419 163.367
R767 B.n943 B.n419 163.367
R768 B.n943 B.n417 163.367
R769 B.n947 B.n417 163.367
R770 B.n947 B.n2 163.367
R771 B.n1086 B.n2 163.367
R772 B.n1086 B.n3 163.367
R773 B.n1082 B.n3 163.367
R774 B.n1082 B.n9 163.367
R775 B.n1078 B.n9 163.367
R776 B.n1078 B.n11 163.367
R777 B.n1074 B.n11 163.367
R778 B.n1074 B.n16 163.367
R779 B.n1070 B.n16 163.367
R780 B.n1070 B.n18 163.367
R781 B.n1066 B.n18 163.367
R782 B.n1066 B.n23 163.367
R783 B.n1062 B.n23 163.367
R784 B.n1062 B.n25 163.367
R785 B.n1058 B.n25 163.367
R786 B.n1058 B.n30 163.367
R787 B.n1054 B.n30 163.367
R788 B.n1054 B.n32 163.367
R789 B.n1050 B.n32 163.367
R790 B.n1050 B.n37 163.367
R791 B.n1046 B.n37 163.367
R792 B.n1046 B.n39 163.367
R793 B.n1042 B.n39 163.367
R794 B.n1042 B.n44 163.367
R795 B.n1038 B.n44 163.367
R796 B.n1038 B.n46 163.367
R797 B.n1034 B.n46 163.367
R798 B.n1034 B.n51 163.367
R799 B.n1030 B.n51 163.367
R800 B.n1030 B.n53 163.367
R801 B.n1026 B.n53 163.367
R802 B.n1026 B.n58 163.367
R803 B.n1022 B.n58 163.367
R804 B.n1022 B.n60 163.367
R805 B.n1018 B.n60 163.367
R806 B.n1018 B.n65 163.367
R807 B.n1014 B.n65 163.367
R808 B.n1014 B.n67 163.367
R809 B.n1010 B.n67 163.367
R810 B.n1010 B.n72 163.367
R811 B.n831 B.n491 163.367
R812 B.n831 B.n559 163.367
R813 B.n827 B.n826 163.367
R814 B.n823 B.n822 163.367
R815 B.n819 B.n818 163.367
R816 B.n815 B.n814 163.367
R817 B.n811 B.n810 163.367
R818 B.n807 B.n806 163.367
R819 B.n803 B.n802 163.367
R820 B.n799 B.n798 163.367
R821 B.n795 B.n794 163.367
R822 B.n791 B.n790 163.367
R823 B.n787 B.n786 163.367
R824 B.n783 B.n782 163.367
R825 B.n779 B.n778 163.367
R826 B.n775 B.n774 163.367
R827 B.n771 B.n770 163.367
R828 B.n767 B.n766 163.367
R829 B.n763 B.n762 163.367
R830 B.n759 B.n758 163.367
R831 B.n755 B.n754 163.367
R832 B.n751 B.n750 163.367
R833 B.n747 B.n746 163.367
R834 B.n743 B.n742 163.367
R835 B.n739 B.n738 163.367
R836 B.n735 B.n734 163.367
R837 B.n731 B.n730 163.367
R838 B.n727 B.n726 163.367
R839 B.n723 B.n722 163.367
R840 B.n719 B.n718 163.367
R841 B.n715 B.n714 163.367
R842 B.n711 B.n710 163.367
R843 B.n707 B.n706 163.367
R844 B.n703 B.n702 163.367
R845 B.n699 B.n698 163.367
R846 B.n695 B.n694 163.367
R847 B.n691 B.n690 163.367
R848 B.n687 B.n686 163.367
R849 B.n683 B.n682 163.367
R850 B.n679 B.n678 163.367
R851 B.n675 B.n674 163.367
R852 B.n671 B.n670 163.367
R853 B.n667 B.n666 163.367
R854 B.n663 B.n662 163.367
R855 B.n659 B.n658 163.367
R856 B.n655 B.n654 163.367
R857 B.n651 B.n650 163.367
R858 B.n647 B.n646 163.367
R859 B.n643 B.n642 163.367
R860 B.n639 B.n638 163.367
R861 B.n635 B.n634 163.367
R862 B.n631 B.n630 163.367
R863 B.n627 B.n626 163.367
R864 B.n623 B.n622 163.367
R865 B.n619 B.n618 163.367
R866 B.n615 B.n614 163.367
R867 B.n611 B.n610 163.367
R868 B.n607 B.n606 163.367
R869 B.n603 B.n602 163.367
R870 B.n599 B.n598 163.367
R871 B.n595 B.n594 163.367
R872 B.n591 B.n590 163.367
R873 B.n587 B.n586 163.367
R874 B.n583 B.n582 163.367
R875 B.n579 B.n578 163.367
R876 B.n575 B.n574 163.367
R877 B.n571 B.n570 163.367
R878 B.n567 B.n558 163.367
R879 B.n840 B.n487 163.367
R880 B.n840 B.n485 163.367
R881 B.n844 B.n485 163.367
R882 B.n844 B.n479 163.367
R883 B.n852 B.n479 163.367
R884 B.n852 B.n477 163.367
R885 B.n856 B.n477 163.367
R886 B.n856 B.n471 163.367
R887 B.n864 B.n471 163.367
R888 B.n864 B.n469 163.367
R889 B.n868 B.n469 163.367
R890 B.n868 B.n463 163.367
R891 B.n876 B.n463 163.367
R892 B.n876 B.n461 163.367
R893 B.n880 B.n461 163.367
R894 B.n880 B.n454 163.367
R895 B.n888 B.n454 163.367
R896 B.n888 B.n452 163.367
R897 B.n892 B.n452 163.367
R898 B.n892 B.n447 163.367
R899 B.n900 B.n447 163.367
R900 B.n900 B.n445 163.367
R901 B.n904 B.n445 163.367
R902 B.n904 B.n439 163.367
R903 B.n912 B.n439 163.367
R904 B.n912 B.n437 163.367
R905 B.n916 B.n437 163.367
R906 B.n916 B.n431 163.367
R907 B.n924 B.n431 163.367
R908 B.n924 B.n429 163.367
R909 B.n928 B.n429 163.367
R910 B.n928 B.n423 163.367
R911 B.n936 B.n423 163.367
R912 B.n936 B.n421 163.367
R913 B.n941 B.n421 163.367
R914 B.n941 B.n415 163.367
R915 B.n949 B.n415 163.367
R916 B.n950 B.n949 163.367
R917 B.n950 B.n5 163.367
R918 B.n6 B.n5 163.367
R919 B.n7 B.n6 163.367
R920 B.n955 B.n7 163.367
R921 B.n955 B.n12 163.367
R922 B.n13 B.n12 163.367
R923 B.n14 B.n13 163.367
R924 B.n960 B.n14 163.367
R925 B.n960 B.n19 163.367
R926 B.n20 B.n19 163.367
R927 B.n21 B.n20 163.367
R928 B.n965 B.n21 163.367
R929 B.n965 B.n26 163.367
R930 B.n27 B.n26 163.367
R931 B.n28 B.n27 163.367
R932 B.n970 B.n28 163.367
R933 B.n970 B.n33 163.367
R934 B.n34 B.n33 163.367
R935 B.n35 B.n34 163.367
R936 B.n975 B.n35 163.367
R937 B.n975 B.n40 163.367
R938 B.n41 B.n40 163.367
R939 B.n42 B.n41 163.367
R940 B.n980 B.n42 163.367
R941 B.n980 B.n47 163.367
R942 B.n48 B.n47 163.367
R943 B.n49 B.n48 163.367
R944 B.n985 B.n49 163.367
R945 B.n985 B.n54 163.367
R946 B.n55 B.n54 163.367
R947 B.n56 B.n55 163.367
R948 B.n990 B.n56 163.367
R949 B.n990 B.n61 163.367
R950 B.n62 B.n61 163.367
R951 B.n63 B.n62 163.367
R952 B.n995 B.n63 163.367
R953 B.n995 B.n68 163.367
R954 B.n69 B.n68 163.367
R955 B.n70 B.n69 163.367
R956 B.n142 B.n70 163.367
R957 B.n147 B.n74 163.367
R958 B.n151 B.n150 163.367
R959 B.n155 B.n154 163.367
R960 B.n159 B.n158 163.367
R961 B.n163 B.n162 163.367
R962 B.n167 B.n166 163.367
R963 B.n171 B.n170 163.367
R964 B.n175 B.n174 163.367
R965 B.n179 B.n178 163.367
R966 B.n183 B.n182 163.367
R967 B.n187 B.n186 163.367
R968 B.n191 B.n190 163.367
R969 B.n195 B.n194 163.367
R970 B.n199 B.n198 163.367
R971 B.n203 B.n202 163.367
R972 B.n207 B.n206 163.367
R973 B.n211 B.n210 163.367
R974 B.n215 B.n214 163.367
R975 B.n219 B.n218 163.367
R976 B.n223 B.n222 163.367
R977 B.n227 B.n226 163.367
R978 B.n231 B.n230 163.367
R979 B.n235 B.n234 163.367
R980 B.n239 B.n238 163.367
R981 B.n243 B.n242 163.367
R982 B.n247 B.n246 163.367
R983 B.n251 B.n250 163.367
R984 B.n255 B.n254 163.367
R985 B.n259 B.n258 163.367
R986 B.n263 B.n262 163.367
R987 B.n267 B.n266 163.367
R988 B.n272 B.n271 163.367
R989 B.n276 B.n275 163.367
R990 B.n280 B.n279 163.367
R991 B.n284 B.n283 163.367
R992 B.n288 B.n287 163.367
R993 B.n293 B.n292 163.367
R994 B.n297 B.n296 163.367
R995 B.n301 B.n300 163.367
R996 B.n305 B.n304 163.367
R997 B.n309 B.n308 163.367
R998 B.n313 B.n312 163.367
R999 B.n317 B.n316 163.367
R1000 B.n321 B.n320 163.367
R1001 B.n325 B.n324 163.367
R1002 B.n329 B.n328 163.367
R1003 B.n333 B.n332 163.367
R1004 B.n337 B.n336 163.367
R1005 B.n341 B.n340 163.367
R1006 B.n345 B.n344 163.367
R1007 B.n349 B.n348 163.367
R1008 B.n353 B.n352 163.367
R1009 B.n357 B.n356 163.367
R1010 B.n361 B.n360 163.367
R1011 B.n365 B.n364 163.367
R1012 B.n369 B.n368 163.367
R1013 B.n373 B.n372 163.367
R1014 B.n377 B.n376 163.367
R1015 B.n381 B.n380 163.367
R1016 B.n385 B.n384 163.367
R1017 B.n389 B.n388 163.367
R1018 B.n393 B.n392 163.367
R1019 B.n397 B.n396 163.367
R1020 B.n401 B.n400 163.367
R1021 B.n405 B.n404 163.367
R1022 B.n409 B.n408 163.367
R1023 B.n411 B.n141 163.367
R1024 B.n563 B.t11 123.031
R1025 B.n143 B.t17 123.031
R1026 B.n560 B.t8 123.005
R1027 B.n145 B.t14 123.005
R1028 B.n564 B.t10 72.0253
R1029 B.n144 B.t18 72.0253
R1030 B.n561 B.t7 71.9996
R1031 B.n146 B.t15 71.9996
R1032 B.n834 B.n833 71.676
R1033 B.n559 B.n492 71.676
R1034 B.n826 B.n493 71.676
R1035 B.n822 B.n494 71.676
R1036 B.n818 B.n495 71.676
R1037 B.n814 B.n496 71.676
R1038 B.n810 B.n497 71.676
R1039 B.n806 B.n498 71.676
R1040 B.n802 B.n499 71.676
R1041 B.n798 B.n500 71.676
R1042 B.n794 B.n501 71.676
R1043 B.n790 B.n502 71.676
R1044 B.n786 B.n503 71.676
R1045 B.n782 B.n504 71.676
R1046 B.n778 B.n505 71.676
R1047 B.n774 B.n506 71.676
R1048 B.n770 B.n507 71.676
R1049 B.n766 B.n508 71.676
R1050 B.n762 B.n509 71.676
R1051 B.n758 B.n510 71.676
R1052 B.n754 B.n511 71.676
R1053 B.n750 B.n512 71.676
R1054 B.n746 B.n513 71.676
R1055 B.n742 B.n514 71.676
R1056 B.n738 B.n515 71.676
R1057 B.n734 B.n516 71.676
R1058 B.n730 B.n517 71.676
R1059 B.n726 B.n518 71.676
R1060 B.n722 B.n519 71.676
R1061 B.n718 B.n520 71.676
R1062 B.n714 B.n521 71.676
R1063 B.n710 B.n522 71.676
R1064 B.n706 B.n523 71.676
R1065 B.n702 B.n524 71.676
R1066 B.n698 B.n525 71.676
R1067 B.n694 B.n526 71.676
R1068 B.n690 B.n527 71.676
R1069 B.n686 B.n528 71.676
R1070 B.n682 B.n529 71.676
R1071 B.n678 B.n530 71.676
R1072 B.n674 B.n531 71.676
R1073 B.n670 B.n532 71.676
R1074 B.n666 B.n533 71.676
R1075 B.n662 B.n534 71.676
R1076 B.n658 B.n535 71.676
R1077 B.n654 B.n536 71.676
R1078 B.n650 B.n537 71.676
R1079 B.n646 B.n538 71.676
R1080 B.n642 B.n539 71.676
R1081 B.n638 B.n540 71.676
R1082 B.n634 B.n541 71.676
R1083 B.n630 B.n542 71.676
R1084 B.n626 B.n543 71.676
R1085 B.n622 B.n544 71.676
R1086 B.n618 B.n545 71.676
R1087 B.n614 B.n546 71.676
R1088 B.n610 B.n547 71.676
R1089 B.n606 B.n548 71.676
R1090 B.n602 B.n549 71.676
R1091 B.n598 B.n550 71.676
R1092 B.n594 B.n551 71.676
R1093 B.n590 B.n552 71.676
R1094 B.n586 B.n553 71.676
R1095 B.n582 B.n554 71.676
R1096 B.n578 B.n555 71.676
R1097 B.n574 B.n556 71.676
R1098 B.n570 B.n557 71.676
R1099 B.n1006 B.n1005 71.676
R1100 B.n147 B.n75 71.676
R1101 B.n151 B.n76 71.676
R1102 B.n155 B.n77 71.676
R1103 B.n159 B.n78 71.676
R1104 B.n163 B.n79 71.676
R1105 B.n167 B.n80 71.676
R1106 B.n171 B.n81 71.676
R1107 B.n175 B.n82 71.676
R1108 B.n179 B.n83 71.676
R1109 B.n183 B.n84 71.676
R1110 B.n187 B.n85 71.676
R1111 B.n191 B.n86 71.676
R1112 B.n195 B.n87 71.676
R1113 B.n199 B.n88 71.676
R1114 B.n203 B.n89 71.676
R1115 B.n207 B.n90 71.676
R1116 B.n211 B.n91 71.676
R1117 B.n215 B.n92 71.676
R1118 B.n219 B.n93 71.676
R1119 B.n223 B.n94 71.676
R1120 B.n227 B.n95 71.676
R1121 B.n231 B.n96 71.676
R1122 B.n235 B.n97 71.676
R1123 B.n239 B.n98 71.676
R1124 B.n243 B.n99 71.676
R1125 B.n247 B.n100 71.676
R1126 B.n251 B.n101 71.676
R1127 B.n255 B.n102 71.676
R1128 B.n259 B.n103 71.676
R1129 B.n263 B.n104 71.676
R1130 B.n267 B.n105 71.676
R1131 B.n272 B.n106 71.676
R1132 B.n276 B.n107 71.676
R1133 B.n280 B.n108 71.676
R1134 B.n284 B.n109 71.676
R1135 B.n288 B.n110 71.676
R1136 B.n293 B.n111 71.676
R1137 B.n297 B.n112 71.676
R1138 B.n301 B.n113 71.676
R1139 B.n305 B.n114 71.676
R1140 B.n309 B.n115 71.676
R1141 B.n313 B.n116 71.676
R1142 B.n317 B.n117 71.676
R1143 B.n321 B.n118 71.676
R1144 B.n325 B.n119 71.676
R1145 B.n329 B.n120 71.676
R1146 B.n333 B.n121 71.676
R1147 B.n337 B.n122 71.676
R1148 B.n341 B.n123 71.676
R1149 B.n345 B.n124 71.676
R1150 B.n349 B.n125 71.676
R1151 B.n353 B.n126 71.676
R1152 B.n357 B.n127 71.676
R1153 B.n361 B.n128 71.676
R1154 B.n365 B.n129 71.676
R1155 B.n369 B.n130 71.676
R1156 B.n373 B.n131 71.676
R1157 B.n377 B.n132 71.676
R1158 B.n381 B.n133 71.676
R1159 B.n385 B.n134 71.676
R1160 B.n389 B.n135 71.676
R1161 B.n393 B.n136 71.676
R1162 B.n397 B.n137 71.676
R1163 B.n401 B.n138 71.676
R1164 B.n405 B.n139 71.676
R1165 B.n409 B.n140 71.676
R1166 B.n1003 B.n141 71.676
R1167 B.n1003 B.n1002 71.676
R1168 B.n411 B.n140 71.676
R1169 B.n408 B.n139 71.676
R1170 B.n404 B.n138 71.676
R1171 B.n400 B.n137 71.676
R1172 B.n396 B.n136 71.676
R1173 B.n392 B.n135 71.676
R1174 B.n388 B.n134 71.676
R1175 B.n384 B.n133 71.676
R1176 B.n380 B.n132 71.676
R1177 B.n376 B.n131 71.676
R1178 B.n372 B.n130 71.676
R1179 B.n368 B.n129 71.676
R1180 B.n364 B.n128 71.676
R1181 B.n360 B.n127 71.676
R1182 B.n356 B.n126 71.676
R1183 B.n352 B.n125 71.676
R1184 B.n348 B.n124 71.676
R1185 B.n344 B.n123 71.676
R1186 B.n340 B.n122 71.676
R1187 B.n336 B.n121 71.676
R1188 B.n332 B.n120 71.676
R1189 B.n328 B.n119 71.676
R1190 B.n324 B.n118 71.676
R1191 B.n320 B.n117 71.676
R1192 B.n316 B.n116 71.676
R1193 B.n312 B.n115 71.676
R1194 B.n308 B.n114 71.676
R1195 B.n304 B.n113 71.676
R1196 B.n300 B.n112 71.676
R1197 B.n296 B.n111 71.676
R1198 B.n292 B.n110 71.676
R1199 B.n287 B.n109 71.676
R1200 B.n283 B.n108 71.676
R1201 B.n279 B.n107 71.676
R1202 B.n275 B.n106 71.676
R1203 B.n271 B.n105 71.676
R1204 B.n266 B.n104 71.676
R1205 B.n262 B.n103 71.676
R1206 B.n258 B.n102 71.676
R1207 B.n254 B.n101 71.676
R1208 B.n250 B.n100 71.676
R1209 B.n246 B.n99 71.676
R1210 B.n242 B.n98 71.676
R1211 B.n238 B.n97 71.676
R1212 B.n234 B.n96 71.676
R1213 B.n230 B.n95 71.676
R1214 B.n226 B.n94 71.676
R1215 B.n222 B.n93 71.676
R1216 B.n218 B.n92 71.676
R1217 B.n214 B.n91 71.676
R1218 B.n210 B.n90 71.676
R1219 B.n206 B.n89 71.676
R1220 B.n202 B.n88 71.676
R1221 B.n198 B.n87 71.676
R1222 B.n194 B.n86 71.676
R1223 B.n190 B.n85 71.676
R1224 B.n186 B.n84 71.676
R1225 B.n182 B.n83 71.676
R1226 B.n178 B.n82 71.676
R1227 B.n174 B.n81 71.676
R1228 B.n170 B.n80 71.676
R1229 B.n166 B.n79 71.676
R1230 B.n162 B.n78 71.676
R1231 B.n158 B.n77 71.676
R1232 B.n154 B.n76 71.676
R1233 B.n150 B.n75 71.676
R1234 B.n1005 B.n74 71.676
R1235 B.n833 B.n491 71.676
R1236 B.n827 B.n492 71.676
R1237 B.n823 B.n493 71.676
R1238 B.n819 B.n494 71.676
R1239 B.n815 B.n495 71.676
R1240 B.n811 B.n496 71.676
R1241 B.n807 B.n497 71.676
R1242 B.n803 B.n498 71.676
R1243 B.n799 B.n499 71.676
R1244 B.n795 B.n500 71.676
R1245 B.n791 B.n501 71.676
R1246 B.n787 B.n502 71.676
R1247 B.n783 B.n503 71.676
R1248 B.n779 B.n504 71.676
R1249 B.n775 B.n505 71.676
R1250 B.n771 B.n506 71.676
R1251 B.n767 B.n507 71.676
R1252 B.n763 B.n508 71.676
R1253 B.n759 B.n509 71.676
R1254 B.n755 B.n510 71.676
R1255 B.n751 B.n511 71.676
R1256 B.n747 B.n512 71.676
R1257 B.n743 B.n513 71.676
R1258 B.n739 B.n514 71.676
R1259 B.n735 B.n515 71.676
R1260 B.n731 B.n516 71.676
R1261 B.n727 B.n517 71.676
R1262 B.n723 B.n518 71.676
R1263 B.n719 B.n519 71.676
R1264 B.n715 B.n520 71.676
R1265 B.n711 B.n521 71.676
R1266 B.n707 B.n522 71.676
R1267 B.n703 B.n523 71.676
R1268 B.n699 B.n524 71.676
R1269 B.n695 B.n525 71.676
R1270 B.n691 B.n526 71.676
R1271 B.n687 B.n527 71.676
R1272 B.n683 B.n528 71.676
R1273 B.n679 B.n529 71.676
R1274 B.n675 B.n530 71.676
R1275 B.n671 B.n531 71.676
R1276 B.n667 B.n532 71.676
R1277 B.n663 B.n533 71.676
R1278 B.n659 B.n534 71.676
R1279 B.n655 B.n535 71.676
R1280 B.n651 B.n536 71.676
R1281 B.n647 B.n537 71.676
R1282 B.n643 B.n538 71.676
R1283 B.n639 B.n539 71.676
R1284 B.n635 B.n540 71.676
R1285 B.n631 B.n541 71.676
R1286 B.n627 B.n542 71.676
R1287 B.n623 B.n543 71.676
R1288 B.n619 B.n544 71.676
R1289 B.n615 B.n545 71.676
R1290 B.n611 B.n546 71.676
R1291 B.n607 B.n547 71.676
R1292 B.n603 B.n548 71.676
R1293 B.n599 B.n549 71.676
R1294 B.n595 B.n550 71.676
R1295 B.n591 B.n551 71.676
R1296 B.n587 B.n552 71.676
R1297 B.n583 B.n553 71.676
R1298 B.n579 B.n554 71.676
R1299 B.n575 B.n555 71.676
R1300 B.n571 B.n556 71.676
R1301 B.n567 B.n557 71.676
R1302 B.n565 B.n564 59.5399
R1303 B.n562 B.n561 59.5399
R1304 B.n269 B.n146 59.5399
R1305 B.n290 B.n144 59.5399
R1306 B.n832 B.n488 56.87
R1307 B.n1004 B.n71 56.87
R1308 B.n564 B.n563 51.0066
R1309 B.n561 B.n560 51.0066
R1310 B.n146 B.n145 51.0066
R1311 B.n144 B.n143 51.0066
R1312 B.n1008 B.n1007 31.3761
R1313 B.n1001 B.n1000 31.3761
R1314 B.n566 B.n486 31.3761
R1315 B.n836 B.n835 31.3761
R1316 B.n839 B.n488 30.4503
R1317 B.n839 B.n484 30.4503
R1318 B.n845 B.n484 30.4503
R1319 B.n845 B.n480 30.4503
R1320 B.n851 B.n480 30.4503
R1321 B.n851 B.n476 30.4503
R1322 B.n857 B.n476 30.4503
R1323 B.n863 B.n472 30.4503
R1324 B.n863 B.n468 30.4503
R1325 B.n869 B.n468 30.4503
R1326 B.n869 B.n464 30.4503
R1327 B.n875 B.n464 30.4503
R1328 B.n875 B.n460 30.4503
R1329 B.n881 B.n460 30.4503
R1330 B.n881 B.n455 30.4503
R1331 B.n887 B.n455 30.4503
R1332 B.n887 B.n456 30.4503
R1333 B.n893 B.n448 30.4503
R1334 B.n899 B.n448 30.4503
R1335 B.n899 B.n444 30.4503
R1336 B.n905 B.n444 30.4503
R1337 B.n905 B.n440 30.4503
R1338 B.n911 B.n440 30.4503
R1339 B.n917 B.n436 30.4503
R1340 B.n917 B.n432 30.4503
R1341 B.n923 B.n432 30.4503
R1342 B.n923 B.n428 30.4503
R1343 B.n929 B.n428 30.4503
R1344 B.n929 B.n424 30.4503
R1345 B.n935 B.n424 30.4503
R1346 B.n942 B.n420 30.4503
R1347 B.n942 B.n416 30.4503
R1348 B.n948 B.n416 30.4503
R1349 B.n948 B.n4 30.4503
R1350 B.n1085 B.n4 30.4503
R1351 B.n1085 B.n1084 30.4503
R1352 B.n1084 B.n1083 30.4503
R1353 B.n1083 B.n8 30.4503
R1354 B.n1077 B.n8 30.4503
R1355 B.n1077 B.n1076 30.4503
R1356 B.n1075 B.n15 30.4503
R1357 B.n1069 B.n15 30.4503
R1358 B.n1069 B.n1068 30.4503
R1359 B.n1068 B.n1067 30.4503
R1360 B.n1067 B.n22 30.4503
R1361 B.n1061 B.n22 30.4503
R1362 B.n1061 B.n1060 30.4503
R1363 B.n1059 B.n29 30.4503
R1364 B.n1053 B.n29 30.4503
R1365 B.n1053 B.n1052 30.4503
R1366 B.n1052 B.n1051 30.4503
R1367 B.n1051 B.n36 30.4503
R1368 B.n1045 B.n36 30.4503
R1369 B.n1044 B.n1043 30.4503
R1370 B.n1043 B.n43 30.4503
R1371 B.n1037 B.n43 30.4503
R1372 B.n1037 B.n1036 30.4503
R1373 B.n1036 B.n1035 30.4503
R1374 B.n1035 B.n50 30.4503
R1375 B.n1029 B.n50 30.4503
R1376 B.n1029 B.n1028 30.4503
R1377 B.n1028 B.n1027 30.4503
R1378 B.n1027 B.n57 30.4503
R1379 B.n1021 B.n1020 30.4503
R1380 B.n1020 B.n1019 30.4503
R1381 B.n1019 B.n64 30.4503
R1382 B.n1013 B.n64 30.4503
R1383 B.n1013 B.n1012 30.4503
R1384 B.n1012 B.n1011 30.4503
R1385 B.n1011 B.n71 30.4503
R1386 B.n893 B.t19 28.6592
R1387 B.n1045 B.t4 28.6592
R1388 B.t6 B.n472 26.868
R1389 B.t13 B.n57 26.868
R1390 B.n911 B.t2 24.1812
R1391 B.t0 B.n1059 24.1812
R1392 B B.n1087 18.0485
R1393 B.n935 B.t3 16.121
R1394 B.t1 B.n1075 16.121
R1395 B.t3 B.n420 14.3298
R1396 B.n1076 B.t1 14.3298
R1397 B.n1007 B.n73 10.6151
R1398 B.n148 B.n73 10.6151
R1399 B.n149 B.n148 10.6151
R1400 B.n152 B.n149 10.6151
R1401 B.n153 B.n152 10.6151
R1402 B.n156 B.n153 10.6151
R1403 B.n157 B.n156 10.6151
R1404 B.n160 B.n157 10.6151
R1405 B.n161 B.n160 10.6151
R1406 B.n164 B.n161 10.6151
R1407 B.n165 B.n164 10.6151
R1408 B.n168 B.n165 10.6151
R1409 B.n169 B.n168 10.6151
R1410 B.n172 B.n169 10.6151
R1411 B.n173 B.n172 10.6151
R1412 B.n176 B.n173 10.6151
R1413 B.n177 B.n176 10.6151
R1414 B.n180 B.n177 10.6151
R1415 B.n181 B.n180 10.6151
R1416 B.n184 B.n181 10.6151
R1417 B.n185 B.n184 10.6151
R1418 B.n188 B.n185 10.6151
R1419 B.n189 B.n188 10.6151
R1420 B.n192 B.n189 10.6151
R1421 B.n193 B.n192 10.6151
R1422 B.n196 B.n193 10.6151
R1423 B.n197 B.n196 10.6151
R1424 B.n200 B.n197 10.6151
R1425 B.n201 B.n200 10.6151
R1426 B.n204 B.n201 10.6151
R1427 B.n205 B.n204 10.6151
R1428 B.n208 B.n205 10.6151
R1429 B.n209 B.n208 10.6151
R1430 B.n212 B.n209 10.6151
R1431 B.n213 B.n212 10.6151
R1432 B.n216 B.n213 10.6151
R1433 B.n217 B.n216 10.6151
R1434 B.n220 B.n217 10.6151
R1435 B.n221 B.n220 10.6151
R1436 B.n224 B.n221 10.6151
R1437 B.n225 B.n224 10.6151
R1438 B.n228 B.n225 10.6151
R1439 B.n229 B.n228 10.6151
R1440 B.n232 B.n229 10.6151
R1441 B.n233 B.n232 10.6151
R1442 B.n236 B.n233 10.6151
R1443 B.n237 B.n236 10.6151
R1444 B.n240 B.n237 10.6151
R1445 B.n241 B.n240 10.6151
R1446 B.n244 B.n241 10.6151
R1447 B.n245 B.n244 10.6151
R1448 B.n248 B.n245 10.6151
R1449 B.n249 B.n248 10.6151
R1450 B.n252 B.n249 10.6151
R1451 B.n253 B.n252 10.6151
R1452 B.n256 B.n253 10.6151
R1453 B.n257 B.n256 10.6151
R1454 B.n260 B.n257 10.6151
R1455 B.n261 B.n260 10.6151
R1456 B.n264 B.n261 10.6151
R1457 B.n265 B.n264 10.6151
R1458 B.n268 B.n265 10.6151
R1459 B.n273 B.n270 10.6151
R1460 B.n274 B.n273 10.6151
R1461 B.n277 B.n274 10.6151
R1462 B.n278 B.n277 10.6151
R1463 B.n281 B.n278 10.6151
R1464 B.n282 B.n281 10.6151
R1465 B.n285 B.n282 10.6151
R1466 B.n286 B.n285 10.6151
R1467 B.n289 B.n286 10.6151
R1468 B.n294 B.n291 10.6151
R1469 B.n295 B.n294 10.6151
R1470 B.n298 B.n295 10.6151
R1471 B.n299 B.n298 10.6151
R1472 B.n302 B.n299 10.6151
R1473 B.n303 B.n302 10.6151
R1474 B.n306 B.n303 10.6151
R1475 B.n307 B.n306 10.6151
R1476 B.n310 B.n307 10.6151
R1477 B.n311 B.n310 10.6151
R1478 B.n314 B.n311 10.6151
R1479 B.n315 B.n314 10.6151
R1480 B.n318 B.n315 10.6151
R1481 B.n319 B.n318 10.6151
R1482 B.n322 B.n319 10.6151
R1483 B.n323 B.n322 10.6151
R1484 B.n326 B.n323 10.6151
R1485 B.n327 B.n326 10.6151
R1486 B.n330 B.n327 10.6151
R1487 B.n331 B.n330 10.6151
R1488 B.n334 B.n331 10.6151
R1489 B.n335 B.n334 10.6151
R1490 B.n338 B.n335 10.6151
R1491 B.n339 B.n338 10.6151
R1492 B.n342 B.n339 10.6151
R1493 B.n343 B.n342 10.6151
R1494 B.n346 B.n343 10.6151
R1495 B.n347 B.n346 10.6151
R1496 B.n350 B.n347 10.6151
R1497 B.n351 B.n350 10.6151
R1498 B.n354 B.n351 10.6151
R1499 B.n355 B.n354 10.6151
R1500 B.n358 B.n355 10.6151
R1501 B.n359 B.n358 10.6151
R1502 B.n362 B.n359 10.6151
R1503 B.n363 B.n362 10.6151
R1504 B.n366 B.n363 10.6151
R1505 B.n367 B.n366 10.6151
R1506 B.n370 B.n367 10.6151
R1507 B.n371 B.n370 10.6151
R1508 B.n374 B.n371 10.6151
R1509 B.n375 B.n374 10.6151
R1510 B.n378 B.n375 10.6151
R1511 B.n379 B.n378 10.6151
R1512 B.n382 B.n379 10.6151
R1513 B.n383 B.n382 10.6151
R1514 B.n386 B.n383 10.6151
R1515 B.n387 B.n386 10.6151
R1516 B.n390 B.n387 10.6151
R1517 B.n391 B.n390 10.6151
R1518 B.n394 B.n391 10.6151
R1519 B.n395 B.n394 10.6151
R1520 B.n398 B.n395 10.6151
R1521 B.n399 B.n398 10.6151
R1522 B.n402 B.n399 10.6151
R1523 B.n403 B.n402 10.6151
R1524 B.n406 B.n403 10.6151
R1525 B.n407 B.n406 10.6151
R1526 B.n410 B.n407 10.6151
R1527 B.n412 B.n410 10.6151
R1528 B.n413 B.n412 10.6151
R1529 B.n1001 B.n413 10.6151
R1530 B.n841 B.n486 10.6151
R1531 B.n842 B.n841 10.6151
R1532 B.n843 B.n842 10.6151
R1533 B.n843 B.n478 10.6151
R1534 B.n853 B.n478 10.6151
R1535 B.n854 B.n853 10.6151
R1536 B.n855 B.n854 10.6151
R1537 B.n855 B.n470 10.6151
R1538 B.n865 B.n470 10.6151
R1539 B.n866 B.n865 10.6151
R1540 B.n867 B.n866 10.6151
R1541 B.n867 B.n462 10.6151
R1542 B.n877 B.n462 10.6151
R1543 B.n878 B.n877 10.6151
R1544 B.n879 B.n878 10.6151
R1545 B.n879 B.n453 10.6151
R1546 B.n889 B.n453 10.6151
R1547 B.n890 B.n889 10.6151
R1548 B.n891 B.n890 10.6151
R1549 B.n891 B.n446 10.6151
R1550 B.n901 B.n446 10.6151
R1551 B.n902 B.n901 10.6151
R1552 B.n903 B.n902 10.6151
R1553 B.n903 B.n438 10.6151
R1554 B.n913 B.n438 10.6151
R1555 B.n914 B.n913 10.6151
R1556 B.n915 B.n914 10.6151
R1557 B.n915 B.n430 10.6151
R1558 B.n925 B.n430 10.6151
R1559 B.n926 B.n925 10.6151
R1560 B.n927 B.n926 10.6151
R1561 B.n927 B.n422 10.6151
R1562 B.n937 B.n422 10.6151
R1563 B.n938 B.n937 10.6151
R1564 B.n940 B.n938 10.6151
R1565 B.n940 B.n939 10.6151
R1566 B.n939 B.n414 10.6151
R1567 B.n951 B.n414 10.6151
R1568 B.n952 B.n951 10.6151
R1569 B.n953 B.n952 10.6151
R1570 B.n954 B.n953 10.6151
R1571 B.n956 B.n954 10.6151
R1572 B.n957 B.n956 10.6151
R1573 B.n958 B.n957 10.6151
R1574 B.n959 B.n958 10.6151
R1575 B.n961 B.n959 10.6151
R1576 B.n962 B.n961 10.6151
R1577 B.n963 B.n962 10.6151
R1578 B.n964 B.n963 10.6151
R1579 B.n966 B.n964 10.6151
R1580 B.n967 B.n966 10.6151
R1581 B.n968 B.n967 10.6151
R1582 B.n969 B.n968 10.6151
R1583 B.n971 B.n969 10.6151
R1584 B.n972 B.n971 10.6151
R1585 B.n973 B.n972 10.6151
R1586 B.n974 B.n973 10.6151
R1587 B.n976 B.n974 10.6151
R1588 B.n977 B.n976 10.6151
R1589 B.n978 B.n977 10.6151
R1590 B.n979 B.n978 10.6151
R1591 B.n981 B.n979 10.6151
R1592 B.n982 B.n981 10.6151
R1593 B.n983 B.n982 10.6151
R1594 B.n984 B.n983 10.6151
R1595 B.n986 B.n984 10.6151
R1596 B.n987 B.n986 10.6151
R1597 B.n988 B.n987 10.6151
R1598 B.n989 B.n988 10.6151
R1599 B.n991 B.n989 10.6151
R1600 B.n992 B.n991 10.6151
R1601 B.n993 B.n992 10.6151
R1602 B.n994 B.n993 10.6151
R1603 B.n996 B.n994 10.6151
R1604 B.n997 B.n996 10.6151
R1605 B.n998 B.n997 10.6151
R1606 B.n999 B.n998 10.6151
R1607 B.n1000 B.n999 10.6151
R1608 B.n835 B.n490 10.6151
R1609 B.n830 B.n490 10.6151
R1610 B.n830 B.n829 10.6151
R1611 B.n829 B.n828 10.6151
R1612 B.n828 B.n825 10.6151
R1613 B.n825 B.n824 10.6151
R1614 B.n824 B.n821 10.6151
R1615 B.n821 B.n820 10.6151
R1616 B.n820 B.n817 10.6151
R1617 B.n817 B.n816 10.6151
R1618 B.n816 B.n813 10.6151
R1619 B.n813 B.n812 10.6151
R1620 B.n812 B.n809 10.6151
R1621 B.n809 B.n808 10.6151
R1622 B.n808 B.n805 10.6151
R1623 B.n805 B.n804 10.6151
R1624 B.n804 B.n801 10.6151
R1625 B.n801 B.n800 10.6151
R1626 B.n800 B.n797 10.6151
R1627 B.n797 B.n796 10.6151
R1628 B.n796 B.n793 10.6151
R1629 B.n793 B.n792 10.6151
R1630 B.n792 B.n789 10.6151
R1631 B.n789 B.n788 10.6151
R1632 B.n788 B.n785 10.6151
R1633 B.n785 B.n784 10.6151
R1634 B.n784 B.n781 10.6151
R1635 B.n781 B.n780 10.6151
R1636 B.n780 B.n777 10.6151
R1637 B.n777 B.n776 10.6151
R1638 B.n776 B.n773 10.6151
R1639 B.n773 B.n772 10.6151
R1640 B.n772 B.n769 10.6151
R1641 B.n769 B.n768 10.6151
R1642 B.n768 B.n765 10.6151
R1643 B.n765 B.n764 10.6151
R1644 B.n764 B.n761 10.6151
R1645 B.n761 B.n760 10.6151
R1646 B.n760 B.n757 10.6151
R1647 B.n757 B.n756 10.6151
R1648 B.n756 B.n753 10.6151
R1649 B.n753 B.n752 10.6151
R1650 B.n752 B.n749 10.6151
R1651 B.n749 B.n748 10.6151
R1652 B.n748 B.n745 10.6151
R1653 B.n745 B.n744 10.6151
R1654 B.n744 B.n741 10.6151
R1655 B.n741 B.n740 10.6151
R1656 B.n740 B.n737 10.6151
R1657 B.n737 B.n736 10.6151
R1658 B.n736 B.n733 10.6151
R1659 B.n733 B.n732 10.6151
R1660 B.n732 B.n729 10.6151
R1661 B.n729 B.n728 10.6151
R1662 B.n728 B.n725 10.6151
R1663 B.n725 B.n724 10.6151
R1664 B.n724 B.n721 10.6151
R1665 B.n721 B.n720 10.6151
R1666 B.n720 B.n717 10.6151
R1667 B.n717 B.n716 10.6151
R1668 B.n716 B.n713 10.6151
R1669 B.n713 B.n712 10.6151
R1670 B.n709 B.n708 10.6151
R1671 B.n708 B.n705 10.6151
R1672 B.n705 B.n704 10.6151
R1673 B.n704 B.n701 10.6151
R1674 B.n701 B.n700 10.6151
R1675 B.n700 B.n697 10.6151
R1676 B.n697 B.n696 10.6151
R1677 B.n696 B.n693 10.6151
R1678 B.n693 B.n692 10.6151
R1679 B.n689 B.n688 10.6151
R1680 B.n688 B.n685 10.6151
R1681 B.n685 B.n684 10.6151
R1682 B.n684 B.n681 10.6151
R1683 B.n681 B.n680 10.6151
R1684 B.n680 B.n677 10.6151
R1685 B.n677 B.n676 10.6151
R1686 B.n676 B.n673 10.6151
R1687 B.n673 B.n672 10.6151
R1688 B.n672 B.n669 10.6151
R1689 B.n669 B.n668 10.6151
R1690 B.n668 B.n665 10.6151
R1691 B.n665 B.n664 10.6151
R1692 B.n664 B.n661 10.6151
R1693 B.n661 B.n660 10.6151
R1694 B.n660 B.n657 10.6151
R1695 B.n657 B.n656 10.6151
R1696 B.n656 B.n653 10.6151
R1697 B.n653 B.n652 10.6151
R1698 B.n652 B.n649 10.6151
R1699 B.n649 B.n648 10.6151
R1700 B.n648 B.n645 10.6151
R1701 B.n645 B.n644 10.6151
R1702 B.n644 B.n641 10.6151
R1703 B.n641 B.n640 10.6151
R1704 B.n640 B.n637 10.6151
R1705 B.n637 B.n636 10.6151
R1706 B.n636 B.n633 10.6151
R1707 B.n633 B.n632 10.6151
R1708 B.n632 B.n629 10.6151
R1709 B.n629 B.n628 10.6151
R1710 B.n628 B.n625 10.6151
R1711 B.n625 B.n624 10.6151
R1712 B.n624 B.n621 10.6151
R1713 B.n621 B.n620 10.6151
R1714 B.n620 B.n617 10.6151
R1715 B.n617 B.n616 10.6151
R1716 B.n616 B.n613 10.6151
R1717 B.n613 B.n612 10.6151
R1718 B.n612 B.n609 10.6151
R1719 B.n609 B.n608 10.6151
R1720 B.n608 B.n605 10.6151
R1721 B.n605 B.n604 10.6151
R1722 B.n604 B.n601 10.6151
R1723 B.n601 B.n600 10.6151
R1724 B.n600 B.n597 10.6151
R1725 B.n597 B.n596 10.6151
R1726 B.n596 B.n593 10.6151
R1727 B.n593 B.n592 10.6151
R1728 B.n592 B.n589 10.6151
R1729 B.n589 B.n588 10.6151
R1730 B.n588 B.n585 10.6151
R1731 B.n585 B.n584 10.6151
R1732 B.n584 B.n581 10.6151
R1733 B.n581 B.n580 10.6151
R1734 B.n580 B.n577 10.6151
R1735 B.n577 B.n576 10.6151
R1736 B.n576 B.n573 10.6151
R1737 B.n573 B.n572 10.6151
R1738 B.n572 B.n569 10.6151
R1739 B.n569 B.n568 10.6151
R1740 B.n568 B.n566 10.6151
R1741 B.n837 B.n836 10.6151
R1742 B.n837 B.n482 10.6151
R1743 B.n847 B.n482 10.6151
R1744 B.n848 B.n847 10.6151
R1745 B.n849 B.n848 10.6151
R1746 B.n849 B.n474 10.6151
R1747 B.n859 B.n474 10.6151
R1748 B.n860 B.n859 10.6151
R1749 B.n861 B.n860 10.6151
R1750 B.n861 B.n466 10.6151
R1751 B.n871 B.n466 10.6151
R1752 B.n872 B.n871 10.6151
R1753 B.n873 B.n872 10.6151
R1754 B.n873 B.n458 10.6151
R1755 B.n883 B.n458 10.6151
R1756 B.n884 B.n883 10.6151
R1757 B.n885 B.n884 10.6151
R1758 B.n885 B.n450 10.6151
R1759 B.n895 B.n450 10.6151
R1760 B.n896 B.n895 10.6151
R1761 B.n897 B.n896 10.6151
R1762 B.n897 B.n442 10.6151
R1763 B.n907 B.n442 10.6151
R1764 B.n908 B.n907 10.6151
R1765 B.n909 B.n908 10.6151
R1766 B.n909 B.n434 10.6151
R1767 B.n919 B.n434 10.6151
R1768 B.n920 B.n919 10.6151
R1769 B.n921 B.n920 10.6151
R1770 B.n921 B.n426 10.6151
R1771 B.n931 B.n426 10.6151
R1772 B.n932 B.n931 10.6151
R1773 B.n933 B.n932 10.6151
R1774 B.n933 B.n418 10.6151
R1775 B.n944 B.n418 10.6151
R1776 B.n945 B.n944 10.6151
R1777 B.n946 B.n945 10.6151
R1778 B.n946 B.n0 10.6151
R1779 B.n1081 B.n1 10.6151
R1780 B.n1081 B.n1080 10.6151
R1781 B.n1080 B.n1079 10.6151
R1782 B.n1079 B.n10 10.6151
R1783 B.n1073 B.n10 10.6151
R1784 B.n1073 B.n1072 10.6151
R1785 B.n1072 B.n1071 10.6151
R1786 B.n1071 B.n17 10.6151
R1787 B.n1065 B.n17 10.6151
R1788 B.n1065 B.n1064 10.6151
R1789 B.n1064 B.n1063 10.6151
R1790 B.n1063 B.n24 10.6151
R1791 B.n1057 B.n24 10.6151
R1792 B.n1057 B.n1056 10.6151
R1793 B.n1056 B.n1055 10.6151
R1794 B.n1055 B.n31 10.6151
R1795 B.n1049 B.n31 10.6151
R1796 B.n1049 B.n1048 10.6151
R1797 B.n1048 B.n1047 10.6151
R1798 B.n1047 B.n38 10.6151
R1799 B.n1041 B.n38 10.6151
R1800 B.n1041 B.n1040 10.6151
R1801 B.n1040 B.n1039 10.6151
R1802 B.n1039 B.n45 10.6151
R1803 B.n1033 B.n45 10.6151
R1804 B.n1033 B.n1032 10.6151
R1805 B.n1032 B.n1031 10.6151
R1806 B.n1031 B.n52 10.6151
R1807 B.n1025 B.n52 10.6151
R1808 B.n1025 B.n1024 10.6151
R1809 B.n1024 B.n1023 10.6151
R1810 B.n1023 B.n59 10.6151
R1811 B.n1017 B.n59 10.6151
R1812 B.n1017 B.n1016 10.6151
R1813 B.n1016 B.n1015 10.6151
R1814 B.n1015 B.n66 10.6151
R1815 B.n1009 B.n66 10.6151
R1816 B.n1009 B.n1008 10.6151
R1817 B.n269 B.n268 9.36635
R1818 B.n291 B.n290 9.36635
R1819 B.n712 B.n562 9.36635
R1820 B.n689 B.n565 9.36635
R1821 B.t2 B.n436 6.26958
R1822 B.n1060 B.t0 6.26958
R1823 B.n857 B.t6 3.58283
R1824 B.n1021 B.t13 3.58283
R1825 B.n1087 B.n0 2.81026
R1826 B.n1087 B.n1 2.81026
R1827 B.n456 B.t19 1.79167
R1828 B.t4 B.n1044 1.79167
R1829 B.n270 B.n269 1.24928
R1830 B.n290 B.n289 1.24928
R1831 B.n709 B.n562 1.24928
R1832 B.n692 B.n565 1.24928
R1833 VP.n9 VP.t2 235.775
R1834 VP.n5 VP.t5 202.126
R1835 VP.n29 VP.t3 202.126
R1836 VP.n37 VP.t4 202.126
R1837 VP.n18 VP.t0 202.126
R1838 VP.n10 VP.t1 202.126
R1839 VP.n11 VP.n8 161.3
R1840 VP.n13 VP.n12 161.3
R1841 VP.n14 VP.n7 161.3
R1842 VP.n16 VP.n15 161.3
R1843 VP.n17 VP.n6 161.3
R1844 VP.n36 VP.n0 161.3
R1845 VP.n35 VP.n34 161.3
R1846 VP.n33 VP.n1 161.3
R1847 VP.n32 VP.n31 161.3
R1848 VP.n30 VP.n2 161.3
R1849 VP.n28 VP.n27 161.3
R1850 VP.n26 VP.n3 161.3
R1851 VP.n25 VP.n24 161.3
R1852 VP.n23 VP.n4 161.3
R1853 VP.n22 VP.n21 161.3
R1854 VP.n20 VP.n5 92.1615
R1855 VP.n38 VP.n37 92.1615
R1856 VP.n19 VP.n18 92.1615
R1857 VP.n10 VP.n9 59.2386
R1858 VP.n20 VP.n19 53.1019
R1859 VP.n24 VP.n23 46.8066
R1860 VP.n35 VP.n1 46.8066
R1861 VP.n16 VP.n7 46.8066
R1862 VP.n24 VP.n3 34.1802
R1863 VP.n31 VP.n1 34.1802
R1864 VP.n12 VP.n7 34.1802
R1865 VP.n23 VP.n22 24.4675
R1866 VP.n28 VP.n3 24.4675
R1867 VP.n31 VP.n30 24.4675
R1868 VP.n36 VP.n35 24.4675
R1869 VP.n17 VP.n16 24.4675
R1870 VP.n12 VP.n11 24.4675
R1871 VP.n22 VP.n5 18.5954
R1872 VP.n37 VP.n36 18.5954
R1873 VP.n18 VP.n17 18.5954
R1874 VP.n29 VP.n28 12.234
R1875 VP.n30 VP.n29 12.234
R1876 VP.n11 VP.n10 12.234
R1877 VP.n9 VP.n8 9.10819
R1878 VP.n19 VP.n6 0.278367
R1879 VP.n21 VP.n20 0.278367
R1880 VP.n38 VP.n0 0.278367
R1881 VP.n13 VP.n8 0.189894
R1882 VP.n14 VP.n13 0.189894
R1883 VP.n15 VP.n14 0.189894
R1884 VP.n15 VP.n6 0.189894
R1885 VP.n21 VP.n4 0.189894
R1886 VP.n25 VP.n4 0.189894
R1887 VP.n26 VP.n25 0.189894
R1888 VP.n27 VP.n26 0.189894
R1889 VP.n27 VP.n2 0.189894
R1890 VP.n32 VP.n2 0.189894
R1891 VP.n33 VP.n32 0.189894
R1892 VP.n34 VP.n33 0.189894
R1893 VP.n34 VP.n0 0.189894
R1894 VP VP.n38 0.153454
R1895 VTAIL.n7 VTAIL.t3 44.377
R1896 VTAIL.n11 VTAIL.t4 44.3767
R1897 VTAIL.n2 VTAIL.t7 44.3767
R1898 VTAIL.n10 VTAIL.t6 44.3767
R1899 VTAIL.n9 VTAIL.n8 43.3505
R1900 VTAIL.n6 VTAIL.n5 43.3505
R1901 VTAIL.n1 VTAIL.n0 43.3505
R1902 VTAIL.n4 VTAIL.n3 43.3505
R1903 VTAIL.n6 VTAIL.n4 33.5307
R1904 VTAIL.n11 VTAIL.n10 31.2634
R1905 VTAIL.n7 VTAIL.n6 2.26774
R1906 VTAIL.n10 VTAIL.n9 2.26774
R1907 VTAIL.n4 VTAIL.n2 2.26774
R1908 VTAIL VTAIL.n11 1.64274
R1909 VTAIL.n9 VTAIL.n7 1.60395
R1910 VTAIL.n2 VTAIL.n1 1.60395
R1911 VTAIL.n0 VTAIL.t1 1.02694
R1912 VTAIL.n0 VTAIL.t0 1.02694
R1913 VTAIL.n3 VTAIL.t9 1.02694
R1914 VTAIL.n3 VTAIL.t5 1.02694
R1915 VTAIL.n8 VTAIL.t8 1.02694
R1916 VTAIL.n8 VTAIL.t10 1.02694
R1917 VTAIL.n5 VTAIL.t11 1.02694
R1918 VTAIL.n5 VTAIL.t2 1.02694
R1919 VTAIL VTAIL.n1 0.6255
R1920 VDD1 VDD1.t3 62.8144
R1921 VDD1.n1 VDD1.t0 62.7006
R1922 VDD1.n1 VDD1.n0 60.5407
R1923 VDD1.n3 VDD1.n2 60.0291
R1924 VDD1.n3 VDD1.n1 49.4298
R1925 VDD1.n2 VDD1.t4 1.02694
R1926 VDD1.n2 VDD1.t5 1.02694
R1927 VDD1.n0 VDD1.t2 1.02694
R1928 VDD1.n0 VDD1.t1 1.02694
R1929 VDD1 VDD1.n3 0.509121
R1930 VN.n3 VN.t2 235.775
R1931 VN.n17 VN.t0 235.775
R1932 VN.n4 VN.t4 202.126
R1933 VN.n12 VN.t5 202.126
R1934 VN.n18 VN.t1 202.126
R1935 VN.n26 VN.t3 202.126
R1936 VN.n25 VN.n14 161.3
R1937 VN.n24 VN.n23 161.3
R1938 VN.n22 VN.n15 161.3
R1939 VN.n21 VN.n20 161.3
R1940 VN.n19 VN.n16 161.3
R1941 VN.n11 VN.n0 161.3
R1942 VN.n10 VN.n9 161.3
R1943 VN.n8 VN.n1 161.3
R1944 VN.n7 VN.n6 161.3
R1945 VN.n5 VN.n2 161.3
R1946 VN.n13 VN.n12 92.1615
R1947 VN.n27 VN.n26 92.1615
R1948 VN.n4 VN.n3 59.2386
R1949 VN.n18 VN.n17 59.2386
R1950 VN VN.n27 53.3807
R1951 VN.n10 VN.n1 46.8066
R1952 VN.n24 VN.n15 46.8066
R1953 VN.n6 VN.n1 34.1802
R1954 VN.n20 VN.n15 34.1802
R1955 VN.n6 VN.n5 24.4675
R1956 VN.n11 VN.n10 24.4675
R1957 VN.n20 VN.n19 24.4675
R1958 VN.n25 VN.n24 24.4675
R1959 VN.n12 VN.n11 18.5954
R1960 VN.n26 VN.n25 18.5954
R1961 VN.n5 VN.n4 12.234
R1962 VN.n19 VN.n18 12.234
R1963 VN.n17 VN.n16 9.10819
R1964 VN.n3 VN.n2 9.10819
R1965 VN.n27 VN.n14 0.278367
R1966 VN.n13 VN.n0 0.278367
R1967 VN.n23 VN.n14 0.189894
R1968 VN.n23 VN.n22 0.189894
R1969 VN.n22 VN.n21 0.189894
R1970 VN.n21 VN.n16 0.189894
R1971 VN.n7 VN.n2 0.189894
R1972 VN.n8 VN.n7 0.189894
R1973 VN.n9 VN.n8 0.189894
R1974 VN.n9 VN.n0 0.189894
R1975 VN VN.n13 0.153454
R1976 VDD2.n1 VDD2.t3 62.7006
R1977 VDD2.n2 VDD2.t2 61.0558
R1978 VDD2.n1 VDD2.n0 60.5407
R1979 VDD2 VDD2.n3 60.5378
R1980 VDD2.n2 VDD2.n1 47.7131
R1981 VDD2 VDD2.n2 1.75912
R1982 VDD2.n3 VDD2.t4 1.02694
R1983 VDD2.n3 VDD2.t5 1.02694
R1984 VDD2.n0 VDD2.t1 1.02694
R1985 VDD2.n0 VDD2.t0 1.02694
C0 VDD2 VDD1 1.29036f
C1 VN VP 7.98291f
C2 VP VTAIL 10.1045f
C3 VN VTAIL 10.089999f
C4 VP VDD2 0.433428f
C5 VN VDD2 10.319799f
C6 VTAIL VDD2 10.5207f
C7 VP VDD1 10.598401f
C8 VN VDD1 0.15022f
C9 VTAIL VDD1 10.474099f
C10 VDD2 B 7.058592f
C11 VDD1 B 7.370756f
C12 VTAIL B 10.506323f
C13 VN B 12.67171f
C14 VP B 11.096176f
C15 VDD2.t3 B 3.77981f
C16 VDD2.t1 B 0.322929f
C17 VDD2.t0 B 0.322929f
C18 VDD2.n0 B 2.95184f
C19 VDD2.n1 B 2.74953f
C20 VDD2.t2 B 3.77041f
C21 VDD2.n2 B 2.77729f
C22 VDD2.t4 B 0.322929f
C23 VDD2.t5 B 0.322929f
C24 VDD2.n3 B 2.9518f
C25 VN.n0 B 0.031681f
C26 VN.t5 B 2.93617f
C27 VN.n1 B 0.020763f
C28 VN.n2 B 0.206761f
C29 VN.t4 B 2.93617f
C30 VN.t2 B 3.10106f
C31 VN.n3 B 1.06895f
C32 VN.n4 B 1.08171f
C33 VN.n5 B 0.03373f
C34 VN.n6 B 0.048555f
C35 VN.n7 B 0.02403f
C36 VN.n8 B 0.02403f
C37 VN.n9 B 0.02403f
C38 VN.n10 B 0.04563f
C39 VN.n11 B 0.039479f
C40 VN.n12 B 1.10078f
C41 VN.n13 B 0.031298f
C42 VN.n14 B 0.031681f
C43 VN.t3 B 2.93617f
C44 VN.n15 B 0.020763f
C45 VN.n16 B 0.206761f
C46 VN.t1 B 2.93617f
C47 VN.t0 B 3.10106f
C48 VN.n17 B 1.06895f
C49 VN.n18 B 1.08171f
C50 VN.n19 B 0.03373f
C51 VN.n20 B 0.048555f
C52 VN.n21 B 0.02403f
C53 VN.n22 B 0.02403f
C54 VN.n23 B 0.02403f
C55 VN.n24 B 0.04563f
C56 VN.n25 B 0.039479f
C57 VN.n26 B 1.10078f
C58 VN.n27 B 1.46425f
C59 VDD1.t3 B 3.8208f
C60 VDD1.t0 B 3.81995f
C61 VDD1.t2 B 0.326359f
C62 VDD1.t1 B 0.326359f
C63 VDD1.n0 B 2.98319f
C64 VDD1.n1 B 2.88209f
C65 VDD1.t4 B 0.326359f
C66 VDD1.t5 B 0.326359f
C67 VDD1.n2 B 2.97996f
C68 VDD1.n3 B 2.79312f
C69 VTAIL.t1 B 0.339534f
C70 VTAIL.t0 B 0.339534f
C71 VTAIL.n0 B 3.0299f
C72 VTAIL.n1 B 0.387154f
C73 VTAIL.t7 B 3.87225f
C74 VTAIL.n2 B 0.588679f
C75 VTAIL.t9 B 0.339534f
C76 VTAIL.t5 B 0.339534f
C77 VTAIL.n3 B 3.0299f
C78 VTAIL.n4 B 2.21146f
C79 VTAIL.t11 B 0.339534f
C80 VTAIL.t2 B 0.339534f
C81 VTAIL.n5 B 3.0299f
C82 VTAIL.n6 B 2.21147f
C83 VTAIL.t3 B 3.87225f
C84 VTAIL.n7 B 0.588675f
C85 VTAIL.t8 B 0.339534f
C86 VTAIL.t10 B 0.339534f
C87 VTAIL.n8 B 3.0299f
C88 VTAIL.n9 B 0.505027f
C89 VTAIL.t6 B 3.87225f
C90 VTAIL.n10 B 2.1324f
C91 VTAIL.t4 B 3.87225f
C92 VTAIL.n11 B 2.08754f
C93 VP.n0 B 0.032054f
C94 VP.t4 B 2.97072f
C95 VP.n1 B 0.021008f
C96 VP.n2 B 0.024313f
C97 VP.t3 B 2.97072f
C98 VP.n3 B 0.049127f
C99 VP.n4 B 0.024313f
C100 VP.t5 B 2.97072f
C101 VP.n5 B 1.11374f
C102 VP.n6 B 0.032054f
C103 VP.t0 B 2.97072f
C104 VP.n7 B 0.021008f
C105 VP.n8 B 0.209194f
C106 VP.t1 B 2.97072f
C107 VP.t2 B 3.13755f
C108 VP.n9 B 1.08153f
C109 VP.n10 B 1.09444f
C110 VP.n11 B 0.034127f
C111 VP.n12 B 0.049127f
C112 VP.n13 B 0.024313f
C113 VP.n14 B 0.024313f
C114 VP.n15 B 0.024313f
C115 VP.n16 B 0.046167f
C116 VP.n17 B 0.039944f
C117 VP.n18 B 1.11374f
C118 VP.n19 B 1.46853f
C119 VP.n20 B 1.48499f
C120 VP.n21 B 0.032054f
C121 VP.n22 B 0.039944f
C122 VP.n23 B 0.046167f
C123 VP.n24 B 0.021008f
C124 VP.n25 B 0.024313f
C125 VP.n26 B 0.024313f
C126 VP.n27 B 0.024313f
C127 VP.n28 B 0.034127f
C128 VP.n29 B 1.03002f
C129 VP.n30 B 0.034127f
C130 VP.n31 B 0.049127f
C131 VP.n32 B 0.024313f
C132 VP.n33 B 0.024313f
C133 VP.n34 B 0.024313f
C134 VP.n35 B 0.046167f
C135 VP.n36 B 0.039944f
C136 VP.n37 B 1.11374f
C137 VP.n38 B 0.031666f
.ends

