* NGSPICE file created from diff_pair_sample_0321.ext - technology: sky130A

.subckt diff_pair_sample_0321 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.4191 pd=2.87 as=0.9906 ps=5.86 w=2.54 l=0.19
X1 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9906 pd=5.86 as=0 ps=0 w=2.54 l=0.19
X2 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=0.9906 pd=5.86 as=0 ps=0 w=2.54 l=0.19
X3 VTAIL.t5 VN.t1 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9906 pd=5.86 as=0.4191 ps=2.87 w=2.54 l=0.19
X4 VTAIL.t2 VP.t0 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9906 pd=5.86 as=0.4191 ps=2.87 w=2.54 l=0.19
X5 VTAIL.t0 VP.t1 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9906 pd=5.86 as=0.4191 ps=2.87 w=2.54 l=0.19
X6 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.9906 pd=5.86 as=0 ps=0 w=2.54 l=0.19
X7 VDD1.t1 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.4191 pd=2.87 as=0.9906 ps=5.86 w=2.54 l=0.19
X8 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9906 pd=5.86 as=0 ps=0 w=2.54 l=0.19
X9 VDD1.t0 VP.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4191 pd=2.87 as=0.9906 ps=5.86 w=2.54 l=0.19
X10 VDD2.t1 VN.t2 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4191 pd=2.87 as=0.9906 ps=5.86 w=2.54 l=0.19
X11 VTAIL.t4 VN.t3 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9906 pd=5.86 as=0.4191 ps=2.87 w=2.54 l=0.19
R0 VN.n0 VN.t2 525.049
R1 VN.n0 VN.t3 525.049
R2 VN.n1 VN.t1 525.049
R3 VN.n1 VN.t0 525.049
R4 VN VN.n1 193.386
R5 VN VN.n0 161.351
R6 VTAIL.n90 VTAIL.n84 289.615
R7 VTAIL.n6 VTAIL.n0 289.615
R8 VTAIL.n18 VTAIL.n12 289.615
R9 VTAIL.n30 VTAIL.n24 289.615
R10 VTAIL.n78 VTAIL.n72 289.615
R11 VTAIL.n66 VTAIL.n60 289.615
R12 VTAIL.n54 VTAIL.n48 289.615
R13 VTAIL.n42 VTAIL.n36 289.615
R14 VTAIL.n89 VTAIL.n88 185
R15 VTAIL.n91 VTAIL.n90 185
R16 VTAIL.n5 VTAIL.n4 185
R17 VTAIL.n7 VTAIL.n6 185
R18 VTAIL.n17 VTAIL.n16 185
R19 VTAIL.n19 VTAIL.n18 185
R20 VTAIL.n29 VTAIL.n28 185
R21 VTAIL.n31 VTAIL.n30 185
R22 VTAIL.n79 VTAIL.n78 185
R23 VTAIL.n77 VTAIL.n76 185
R24 VTAIL.n67 VTAIL.n66 185
R25 VTAIL.n65 VTAIL.n64 185
R26 VTAIL.n55 VTAIL.n54 185
R27 VTAIL.n53 VTAIL.n52 185
R28 VTAIL.n43 VTAIL.n42 185
R29 VTAIL.n41 VTAIL.n40 185
R30 VTAIL.n87 VTAIL.t6 151.613
R31 VTAIL.n3 VTAIL.t4 151.613
R32 VTAIL.n15 VTAIL.t3 151.613
R33 VTAIL.n27 VTAIL.t2 151.613
R34 VTAIL.n75 VTAIL.t1 151.613
R35 VTAIL.n63 VTAIL.t0 151.613
R36 VTAIL.n51 VTAIL.t7 151.613
R37 VTAIL.n39 VTAIL.t5 151.613
R38 VTAIL.n90 VTAIL.n89 104.615
R39 VTAIL.n6 VTAIL.n5 104.615
R40 VTAIL.n18 VTAIL.n17 104.615
R41 VTAIL.n30 VTAIL.n29 104.615
R42 VTAIL.n78 VTAIL.n77 104.615
R43 VTAIL.n66 VTAIL.n65 104.615
R44 VTAIL.n54 VTAIL.n53 104.615
R45 VTAIL.n42 VTAIL.n41 104.615
R46 VTAIL.n89 VTAIL.t6 52.3082
R47 VTAIL.n5 VTAIL.t4 52.3082
R48 VTAIL.n17 VTAIL.t3 52.3082
R49 VTAIL.n29 VTAIL.t2 52.3082
R50 VTAIL.n77 VTAIL.t1 52.3082
R51 VTAIL.n65 VTAIL.t0 52.3082
R52 VTAIL.n53 VTAIL.t7 52.3082
R53 VTAIL.n41 VTAIL.t5 52.3082
R54 VTAIL.n95 VTAIL.n94 34.9005
R55 VTAIL.n11 VTAIL.n10 34.9005
R56 VTAIL.n23 VTAIL.n22 34.9005
R57 VTAIL.n35 VTAIL.n34 34.9005
R58 VTAIL.n83 VTAIL.n82 34.9005
R59 VTAIL.n71 VTAIL.n70 34.9005
R60 VTAIL.n59 VTAIL.n58 34.9005
R61 VTAIL.n47 VTAIL.n46 34.9005
R62 VTAIL.n88 VTAIL.n87 15.3979
R63 VTAIL.n4 VTAIL.n3 15.3979
R64 VTAIL.n16 VTAIL.n15 15.3979
R65 VTAIL.n28 VTAIL.n27 15.3979
R66 VTAIL.n76 VTAIL.n75 15.3979
R67 VTAIL.n64 VTAIL.n63 15.3979
R68 VTAIL.n52 VTAIL.n51 15.3979
R69 VTAIL.n40 VTAIL.n39 15.3979
R70 VTAIL.n95 VTAIL.n83 15.0221
R71 VTAIL.n47 VTAIL.n35 15.0221
R72 VTAIL.n91 VTAIL.n86 12.8005
R73 VTAIL.n7 VTAIL.n2 12.8005
R74 VTAIL.n19 VTAIL.n14 12.8005
R75 VTAIL.n31 VTAIL.n26 12.8005
R76 VTAIL.n79 VTAIL.n74 12.8005
R77 VTAIL.n67 VTAIL.n62 12.8005
R78 VTAIL.n55 VTAIL.n50 12.8005
R79 VTAIL.n43 VTAIL.n38 12.8005
R80 VTAIL.n92 VTAIL.n84 12.0247
R81 VTAIL.n8 VTAIL.n0 12.0247
R82 VTAIL.n20 VTAIL.n12 12.0247
R83 VTAIL.n32 VTAIL.n24 12.0247
R84 VTAIL.n80 VTAIL.n72 12.0247
R85 VTAIL.n68 VTAIL.n60 12.0247
R86 VTAIL.n56 VTAIL.n48 12.0247
R87 VTAIL.n44 VTAIL.n36 12.0247
R88 VTAIL.n94 VTAIL.n93 9.45567
R89 VTAIL.n10 VTAIL.n9 9.45567
R90 VTAIL.n22 VTAIL.n21 9.45567
R91 VTAIL.n34 VTAIL.n33 9.45567
R92 VTAIL.n82 VTAIL.n81 9.45567
R93 VTAIL.n70 VTAIL.n69 9.45567
R94 VTAIL.n58 VTAIL.n57 9.45567
R95 VTAIL.n46 VTAIL.n45 9.45567
R96 VTAIL.n93 VTAIL.n92 9.3005
R97 VTAIL.n86 VTAIL.n85 9.3005
R98 VTAIL.n9 VTAIL.n8 9.3005
R99 VTAIL.n2 VTAIL.n1 9.3005
R100 VTAIL.n21 VTAIL.n20 9.3005
R101 VTAIL.n14 VTAIL.n13 9.3005
R102 VTAIL.n33 VTAIL.n32 9.3005
R103 VTAIL.n26 VTAIL.n25 9.3005
R104 VTAIL.n81 VTAIL.n80 9.3005
R105 VTAIL.n74 VTAIL.n73 9.3005
R106 VTAIL.n69 VTAIL.n68 9.3005
R107 VTAIL.n62 VTAIL.n61 9.3005
R108 VTAIL.n57 VTAIL.n56 9.3005
R109 VTAIL.n50 VTAIL.n49 9.3005
R110 VTAIL.n45 VTAIL.n44 9.3005
R111 VTAIL.n38 VTAIL.n37 9.3005
R112 VTAIL.n87 VTAIL.n85 4.69785
R113 VTAIL.n3 VTAIL.n1 4.69785
R114 VTAIL.n15 VTAIL.n13 4.69785
R115 VTAIL.n27 VTAIL.n25 4.69785
R116 VTAIL.n75 VTAIL.n73 4.69785
R117 VTAIL.n63 VTAIL.n61 4.69785
R118 VTAIL.n51 VTAIL.n49 4.69785
R119 VTAIL.n39 VTAIL.n37 4.69785
R120 VTAIL.n94 VTAIL.n84 1.93989
R121 VTAIL.n10 VTAIL.n0 1.93989
R122 VTAIL.n22 VTAIL.n12 1.93989
R123 VTAIL.n34 VTAIL.n24 1.93989
R124 VTAIL.n82 VTAIL.n72 1.93989
R125 VTAIL.n70 VTAIL.n60 1.93989
R126 VTAIL.n58 VTAIL.n48 1.93989
R127 VTAIL.n46 VTAIL.n36 1.93989
R128 VTAIL.n92 VTAIL.n91 1.16414
R129 VTAIL.n8 VTAIL.n7 1.16414
R130 VTAIL.n20 VTAIL.n19 1.16414
R131 VTAIL.n32 VTAIL.n31 1.16414
R132 VTAIL.n80 VTAIL.n79 1.16414
R133 VTAIL.n68 VTAIL.n67 1.16414
R134 VTAIL.n56 VTAIL.n55 1.16414
R135 VTAIL.n44 VTAIL.n43 1.16414
R136 VTAIL.n71 VTAIL.n59 0.470328
R137 VTAIL.n23 VTAIL.n11 0.470328
R138 VTAIL.n59 VTAIL.n47 0.448776
R139 VTAIL.n83 VTAIL.n71 0.448776
R140 VTAIL.n35 VTAIL.n23 0.448776
R141 VTAIL.n88 VTAIL.n86 0.388379
R142 VTAIL.n4 VTAIL.n2 0.388379
R143 VTAIL.n16 VTAIL.n14 0.388379
R144 VTAIL.n28 VTAIL.n26 0.388379
R145 VTAIL.n76 VTAIL.n74 0.388379
R146 VTAIL.n64 VTAIL.n62 0.388379
R147 VTAIL.n52 VTAIL.n50 0.388379
R148 VTAIL.n40 VTAIL.n38 0.388379
R149 VTAIL VTAIL.n11 0.282828
R150 VTAIL VTAIL.n95 0.166448
R151 VTAIL.n93 VTAIL.n85 0.155672
R152 VTAIL.n9 VTAIL.n1 0.155672
R153 VTAIL.n21 VTAIL.n13 0.155672
R154 VTAIL.n33 VTAIL.n25 0.155672
R155 VTAIL.n81 VTAIL.n73 0.155672
R156 VTAIL.n69 VTAIL.n61 0.155672
R157 VTAIL.n57 VTAIL.n49 0.155672
R158 VTAIL.n45 VTAIL.n37 0.155672
R159 VDD2.n2 VDD2.n0 114.941
R160 VDD2.n2 VDD2.n1 87.6743
R161 VDD2.n1 VDD2.t2 7.79578
R162 VDD2.n1 VDD2.t3 7.79578
R163 VDD2.n0 VDD2.t0 7.79578
R164 VDD2.n0 VDD2.t1 7.79578
R165 VDD2 VDD2.n2 0.0586897
R166 B.n225 B.n224 585
R167 B.n225 B.n28 585
R168 B.n228 B.n227 585
R169 B.n229 B.n51 585
R170 B.n231 B.n230 585
R171 B.n233 B.n50 585
R172 B.n236 B.n235 585
R173 B.n237 B.n49 585
R174 B.n239 B.n238 585
R175 B.n241 B.n48 585
R176 B.n244 B.n243 585
R177 B.n245 B.n47 585
R178 B.n247 B.n246 585
R179 B.n249 B.n46 585
R180 B.n252 B.n251 585
R181 B.n254 B.n43 585
R182 B.n256 B.n255 585
R183 B.n258 B.n42 585
R184 B.n261 B.n260 585
R185 B.n262 B.n41 585
R186 B.n264 B.n263 585
R187 B.n266 B.n40 585
R188 B.n268 B.n267 585
R189 B.n270 B.n269 585
R190 B.n273 B.n272 585
R191 B.n274 B.n35 585
R192 B.n276 B.n275 585
R193 B.n278 B.n34 585
R194 B.n281 B.n280 585
R195 B.n282 B.n33 585
R196 B.n284 B.n283 585
R197 B.n286 B.n32 585
R198 B.n289 B.n288 585
R199 B.n290 B.n31 585
R200 B.n292 B.n291 585
R201 B.n294 B.n30 585
R202 B.n297 B.n296 585
R203 B.n298 B.n29 585
R204 B.n223 B.n27 585
R205 B.n301 B.n27 585
R206 B.n222 B.n26 585
R207 B.n302 B.n26 585
R208 B.n221 B.n25 585
R209 B.n303 B.n25 585
R210 B.n220 B.n219 585
R211 B.n219 B.n24 585
R212 B.n218 B.n20 585
R213 B.n309 B.n20 585
R214 B.n217 B.n19 585
R215 B.n310 B.n19 585
R216 B.n216 B.n18 585
R217 B.n311 B.n18 585
R218 B.n215 B.n214 585
R219 B.n214 B.n13 585
R220 B.n213 B.n12 585
R221 B.n317 B.n12 585
R222 B.n212 B.n11 585
R223 B.n318 B.n11 585
R224 B.n211 B.n10 585
R225 B.n319 B.n10 585
R226 B.n210 B.n7 585
R227 B.n322 B.n7 585
R228 B.n209 B.n6 585
R229 B.n323 B.n6 585
R230 B.n208 B.n5 585
R231 B.n324 B.n5 585
R232 B.n207 B.n206 585
R233 B.n206 B.n4 585
R234 B.n205 B.n52 585
R235 B.n205 B.n204 585
R236 B.n195 B.n53 585
R237 B.n54 B.n53 585
R238 B.n197 B.n196 585
R239 B.n198 B.n197 585
R240 B.n194 B.n59 585
R241 B.n59 B.n58 585
R242 B.n193 B.n192 585
R243 B.n192 B.n191 585
R244 B.n61 B.n60 585
R245 B.n62 B.n61 585
R246 B.n184 B.n183 585
R247 B.n185 B.n184 585
R248 B.n182 B.n66 585
R249 B.n70 B.n66 585
R250 B.n181 B.n180 585
R251 B.n180 B.n179 585
R252 B.n68 B.n67 585
R253 B.n69 B.n68 585
R254 B.n172 B.n171 585
R255 B.n173 B.n172 585
R256 B.n73 B.n72 585
R257 B.n98 B.n96 585
R258 B.n99 B.n95 585
R259 B.n99 B.n74 585
R260 B.n102 B.n101 585
R261 B.n103 B.n94 585
R262 B.n105 B.n104 585
R263 B.n107 B.n93 585
R264 B.n110 B.n109 585
R265 B.n111 B.n92 585
R266 B.n113 B.n112 585
R267 B.n115 B.n91 585
R268 B.n118 B.n117 585
R269 B.n119 B.n90 585
R270 B.n124 B.n123 585
R271 B.n126 B.n89 585
R272 B.n129 B.n128 585
R273 B.n130 B.n88 585
R274 B.n132 B.n131 585
R275 B.n134 B.n87 585
R276 B.n137 B.n136 585
R277 B.n138 B.n86 585
R278 B.n140 B.n139 585
R279 B.n142 B.n85 585
R280 B.n145 B.n144 585
R281 B.n146 B.n81 585
R282 B.n148 B.n147 585
R283 B.n150 B.n80 585
R284 B.n153 B.n152 585
R285 B.n154 B.n79 585
R286 B.n156 B.n155 585
R287 B.n158 B.n78 585
R288 B.n161 B.n160 585
R289 B.n162 B.n77 585
R290 B.n164 B.n163 585
R291 B.n166 B.n76 585
R292 B.n169 B.n168 585
R293 B.n170 B.n75 585
R294 B.n175 B.n174 585
R295 B.n174 B.n173 585
R296 B.n176 B.n71 585
R297 B.n71 B.n69 585
R298 B.n178 B.n177 585
R299 B.n179 B.n178 585
R300 B.n65 B.n64 585
R301 B.n70 B.n65 585
R302 B.n187 B.n186 585
R303 B.n186 B.n185 585
R304 B.n188 B.n63 585
R305 B.n63 B.n62 585
R306 B.n190 B.n189 585
R307 B.n191 B.n190 585
R308 B.n57 B.n56 585
R309 B.n58 B.n57 585
R310 B.n200 B.n199 585
R311 B.n199 B.n198 585
R312 B.n201 B.n55 585
R313 B.n55 B.n54 585
R314 B.n203 B.n202 585
R315 B.n204 B.n203 585
R316 B.n3 B.n0 585
R317 B.n4 B.n3 585
R318 B.n321 B.n1 585
R319 B.n322 B.n321 585
R320 B.n320 B.n9 585
R321 B.n320 B.n319 585
R322 B.n15 B.n8 585
R323 B.n318 B.n8 585
R324 B.n316 B.n315 585
R325 B.n317 B.n316 585
R326 B.n314 B.n14 585
R327 B.n14 B.n13 585
R328 B.n313 B.n312 585
R329 B.n312 B.n311 585
R330 B.n17 B.n16 585
R331 B.n310 B.n17 585
R332 B.n308 B.n307 585
R333 B.n309 B.n308 585
R334 B.n306 B.n21 585
R335 B.n24 B.n21 585
R336 B.n305 B.n304 585
R337 B.n304 B.n303 585
R338 B.n23 B.n22 585
R339 B.n302 B.n23 585
R340 B.n300 B.n299 585
R341 B.n301 B.n300 585
R342 B.n325 B.n324 585
R343 B.n323 B.n2 585
R344 B.n36 B.t15 561.701
R345 B.n44 B.t4 561.701
R346 B.n82 B.t8 561.701
R347 B.n120 B.t12 561.701
R348 B.n300 B.n29 554.963
R349 B.n225 B.n27 554.963
R350 B.n172 B.n75 554.963
R351 B.n174 B.n73 554.963
R352 B.n226 B.n28 256.663
R353 B.n232 B.n28 256.663
R354 B.n234 B.n28 256.663
R355 B.n240 B.n28 256.663
R356 B.n242 B.n28 256.663
R357 B.n248 B.n28 256.663
R358 B.n250 B.n28 256.663
R359 B.n257 B.n28 256.663
R360 B.n259 B.n28 256.663
R361 B.n265 B.n28 256.663
R362 B.n39 B.n28 256.663
R363 B.n271 B.n28 256.663
R364 B.n277 B.n28 256.663
R365 B.n279 B.n28 256.663
R366 B.n285 B.n28 256.663
R367 B.n287 B.n28 256.663
R368 B.n293 B.n28 256.663
R369 B.n295 B.n28 256.663
R370 B.n97 B.n74 256.663
R371 B.n100 B.n74 256.663
R372 B.n106 B.n74 256.663
R373 B.n108 B.n74 256.663
R374 B.n114 B.n74 256.663
R375 B.n116 B.n74 256.663
R376 B.n125 B.n74 256.663
R377 B.n127 B.n74 256.663
R378 B.n133 B.n74 256.663
R379 B.n135 B.n74 256.663
R380 B.n141 B.n74 256.663
R381 B.n143 B.n74 256.663
R382 B.n149 B.n74 256.663
R383 B.n151 B.n74 256.663
R384 B.n157 B.n74 256.663
R385 B.n159 B.n74 256.663
R386 B.n165 B.n74 256.663
R387 B.n167 B.n74 256.663
R388 B.n327 B.n326 256.663
R389 B.n173 B.n74 192.343
R390 B.n301 B.n28 192.343
R391 B.n296 B.n294 163.367
R392 B.n292 B.n31 163.367
R393 B.n288 B.n286 163.367
R394 B.n284 B.n33 163.367
R395 B.n280 B.n278 163.367
R396 B.n276 B.n35 163.367
R397 B.n272 B.n270 163.367
R398 B.n267 B.n266 163.367
R399 B.n264 B.n41 163.367
R400 B.n260 B.n258 163.367
R401 B.n256 B.n43 163.367
R402 B.n251 B.n249 163.367
R403 B.n247 B.n47 163.367
R404 B.n243 B.n241 163.367
R405 B.n239 B.n49 163.367
R406 B.n235 B.n233 163.367
R407 B.n231 B.n51 163.367
R408 B.n227 B.n225 163.367
R409 B.n172 B.n68 163.367
R410 B.n180 B.n68 163.367
R411 B.n180 B.n66 163.367
R412 B.n184 B.n66 163.367
R413 B.n184 B.n61 163.367
R414 B.n192 B.n61 163.367
R415 B.n192 B.n59 163.367
R416 B.n197 B.n59 163.367
R417 B.n197 B.n53 163.367
R418 B.n205 B.n53 163.367
R419 B.n206 B.n205 163.367
R420 B.n206 B.n5 163.367
R421 B.n6 B.n5 163.367
R422 B.n7 B.n6 163.367
R423 B.n10 B.n7 163.367
R424 B.n11 B.n10 163.367
R425 B.n12 B.n11 163.367
R426 B.n214 B.n12 163.367
R427 B.n214 B.n18 163.367
R428 B.n19 B.n18 163.367
R429 B.n20 B.n19 163.367
R430 B.n219 B.n20 163.367
R431 B.n219 B.n25 163.367
R432 B.n26 B.n25 163.367
R433 B.n27 B.n26 163.367
R434 B.n99 B.n98 163.367
R435 B.n101 B.n99 163.367
R436 B.n105 B.n94 163.367
R437 B.n109 B.n107 163.367
R438 B.n113 B.n92 163.367
R439 B.n117 B.n115 163.367
R440 B.n124 B.n90 163.367
R441 B.n128 B.n126 163.367
R442 B.n132 B.n88 163.367
R443 B.n136 B.n134 163.367
R444 B.n140 B.n86 163.367
R445 B.n144 B.n142 163.367
R446 B.n148 B.n81 163.367
R447 B.n152 B.n150 163.367
R448 B.n156 B.n79 163.367
R449 B.n160 B.n158 163.367
R450 B.n164 B.n77 163.367
R451 B.n168 B.n166 163.367
R452 B.n174 B.n71 163.367
R453 B.n178 B.n71 163.367
R454 B.n178 B.n65 163.367
R455 B.n186 B.n65 163.367
R456 B.n186 B.n63 163.367
R457 B.n190 B.n63 163.367
R458 B.n190 B.n57 163.367
R459 B.n199 B.n57 163.367
R460 B.n199 B.n55 163.367
R461 B.n203 B.n55 163.367
R462 B.n203 B.n3 163.367
R463 B.n325 B.n3 163.367
R464 B.n321 B.n2 163.367
R465 B.n321 B.n320 163.367
R466 B.n320 B.n8 163.367
R467 B.n316 B.n8 163.367
R468 B.n316 B.n14 163.367
R469 B.n312 B.n14 163.367
R470 B.n312 B.n17 163.367
R471 B.n308 B.n17 163.367
R472 B.n308 B.n21 163.367
R473 B.n304 B.n21 163.367
R474 B.n304 B.n23 163.367
R475 B.n300 B.n23 163.367
R476 B.n44 B.t6 133.56
R477 B.n82 B.t11 133.56
R478 B.n36 B.t16 133.56
R479 B.n120 B.t14 133.56
R480 B.n45 B.t7 123.475
R481 B.n83 B.t10 123.475
R482 B.n37 B.t17 123.475
R483 B.n121 B.t13 123.475
R484 B.n173 B.n69 95.4695
R485 B.n179 B.n69 95.4695
R486 B.n179 B.n70 95.4695
R487 B.n185 B.n62 95.4695
R488 B.n191 B.n62 95.4695
R489 B.n191 B.n58 95.4695
R490 B.n198 B.n58 95.4695
R491 B.n204 B.n54 95.4695
R492 B.n324 B.n4 95.4695
R493 B.n324 B.n323 95.4695
R494 B.n323 B.n322 95.4695
R495 B.n319 B.n318 95.4695
R496 B.n317 B.n13 95.4695
R497 B.n311 B.n13 95.4695
R498 B.n311 B.n310 95.4695
R499 B.n310 B.n309 95.4695
R500 B.n303 B.n24 95.4695
R501 B.n303 B.n302 95.4695
R502 B.n302 B.n301 95.4695
R503 B.n70 B.t9 82.8339
R504 B.t3 B.n4 82.8339
R505 B.n322 B.t0 82.8339
R506 B.n24 B.t5 82.8339
R507 B.n295 B.n29 71.676
R508 B.n294 B.n293 71.676
R509 B.n287 B.n31 71.676
R510 B.n286 B.n285 71.676
R511 B.n279 B.n33 71.676
R512 B.n278 B.n277 71.676
R513 B.n271 B.n35 71.676
R514 B.n270 B.n39 71.676
R515 B.n266 B.n265 71.676
R516 B.n259 B.n41 71.676
R517 B.n258 B.n257 71.676
R518 B.n250 B.n43 71.676
R519 B.n249 B.n248 71.676
R520 B.n242 B.n47 71.676
R521 B.n241 B.n240 71.676
R522 B.n234 B.n49 71.676
R523 B.n233 B.n232 71.676
R524 B.n226 B.n51 71.676
R525 B.n227 B.n226 71.676
R526 B.n232 B.n231 71.676
R527 B.n235 B.n234 71.676
R528 B.n240 B.n239 71.676
R529 B.n243 B.n242 71.676
R530 B.n248 B.n247 71.676
R531 B.n251 B.n250 71.676
R532 B.n257 B.n256 71.676
R533 B.n260 B.n259 71.676
R534 B.n265 B.n264 71.676
R535 B.n267 B.n39 71.676
R536 B.n272 B.n271 71.676
R537 B.n277 B.n276 71.676
R538 B.n280 B.n279 71.676
R539 B.n285 B.n284 71.676
R540 B.n288 B.n287 71.676
R541 B.n293 B.n292 71.676
R542 B.n296 B.n295 71.676
R543 B.n97 B.n73 71.676
R544 B.n101 B.n100 71.676
R545 B.n106 B.n105 71.676
R546 B.n109 B.n108 71.676
R547 B.n114 B.n113 71.676
R548 B.n117 B.n116 71.676
R549 B.n125 B.n124 71.676
R550 B.n128 B.n127 71.676
R551 B.n133 B.n132 71.676
R552 B.n136 B.n135 71.676
R553 B.n141 B.n140 71.676
R554 B.n144 B.n143 71.676
R555 B.n149 B.n148 71.676
R556 B.n152 B.n151 71.676
R557 B.n157 B.n156 71.676
R558 B.n160 B.n159 71.676
R559 B.n165 B.n164 71.676
R560 B.n168 B.n167 71.676
R561 B.n98 B.n97 71.676
R562 B.n100 B.n94 71.676
R563 B.n107 B.n106 71.676
R564 B.n108 B.n92 71.676
R565 B.n115 B.n114 71.676
R566 B.n116 B.n90 71.676
R567 B.n126 B.n125 71.676
R568 B.n127 B.n88 71.676
R569 B.n134 B.n133 71.676
R570 B.n135 B.n86 71.676
R571 B.n142 B.n141 71.676
R572 B.n143 B.n81 71.676
R573 B.n150 B.n149 71.676
R574 B.n151 B.n79 71.676
R575 B.n158 B.n157 71.676
R576 B.n159 B.n77 71.676
R577 B.n166 B.n165 71.676
R578 B.n167 B.n75 71.676
R579 B.n326 B.n325 71.676
R580 B.n326 B.n2 71.676
R581 B.n38 B.n37 59.5399
R582 B.n253 B.n45 59.5399
R583 B.n84 B.n83 59.5399
R584 B.n122 B.n121 59.5399
R585 B.n198 B.t2 57.5627
R586 B.t1 B.n317 57.5627
R587 B.t2 B.n54 37.9073
R588 B.n318 B.t1 37.9073
R589 B.n175 B.n72 36.059
R590 B.n171 B.n170 36.059
R591 B.n224 B.n223 36.059
R592 B.n299 B.n298 36.059
R593 B B.n327 18.0485
R594 B.n185 B.t9 12.6361
R595 B.n204 B.t3 12.6361
R596 B.n319 B.t0 12.6361
R597 B.n309 B.t5 12.6361
R598 B.n176 B.n175 10.6151
R599 B.n177 B.n176 10.6151
R600 B.n177 B.n64 10.6151
R601 B.n187 B.n64 10.6151
R602 B.n188 B.n187 10.6151
R603 B.n189 B.n188 10.6151
R604 B.n189 B.n56 10.6151
R605 B.n200 B.n56 10.6151
R606 B.n201 B.n200 10.6151
R607 B.n202 B.n201 10.6151
R608 B.n202 B.n0 10.6151
R609 B.n96 B.n72 10.6151
R610 B.n96 B.n95 10.6151
R611 B.n102 B.n95 10.6151
R612 B.n103 B.n102 10.6151
R613 B.n104 B.n103 10.6151
R614 B.n104 B.n93 10.6151
R615 B.n110 B.n93 10.6151
R616 B.n111 B.n110 10.6151
R617 B.n112 B.n111 10.6151
R618 B.n112 B.n91 10.6151
R619 B.n118 B.n91 10.6151
R620 B.n119 B.n118 10.6151
R621 B.n123 B.n119 10.6151
R622 B.n129 B.n89 10.6151
R623 B.n130 B.n129 10.6151
R624 B.n131 B.n130 10.6151
R625 B.n131 B.n87 10.6151
R626 B.n137 B.n87 10.6151
R627 B.n138 B.n137 10.6151
R628 B.n139 B.n138 10.6151
R629 B.n139 B.n85 10.6151
R630 B.n146 B.n145 10.6151
R631 B.n147 B.n146 10.6151
R632 B.n147 B.n80 10.6151
R633 B.n153 B.n80 10.6151
R634 B.n154 B.n153 10.6151
R635 B.n155 B.n154 10.6151
R636 B.n155 B.n78 10.6151
R637 B.n161 B.n78 10.6151
R638 B.n162 B.n161 10.6151
R639 B.n163 B.n162 10.6151
R640 B.n163 B.n76 10.6151
R641 B.n169 B.n76 10.6151
R642 B.n170 B.n169 10.6151
R643 B.n171 B.n67 10.6151
R644 B.n181 B.n67 10.6151
R645 B.n182 B.n181 10.6151
R646 B.n183 B.n182 10.6151
R647 B.n183 B.n60 10.6151
R648 B.n193 B.n60 10.6151
R649 B.n194 B.n193 10.6151
R650 B.n196 B.n194 10.6151
R651 B.n196 B.n195 10.6151
R652 B.n195 B.n52 10.6151
R653 B.n207 B.n52 10.6151
R654 B.n208 B.n207 10.6151
R655 B.n209 B.n208 10.6151
R656 B.n210 B.n209 10.6151
R657 B.n211 B.n210 10.6151
R658 B.n212 B.n211 10.6151
R659 B.n213 B.n212 10.6151
R660 B.n215 B.n213 10.6151
R661 B.n216 B.n215 10.6151
R662 B.n217 B.n216 10.6151
R663 B.n218 B.n217 10.6151
R664 B.n220 B.n218 10.6151
R665 B.n221 B.n220 10.6151
R666 B.n222 B.n221 10.6151
R667 B.n223 B.n222 10.6151
R668 B.n9 B.n1 10.6151
R669 B.n15 B.n9 10.6151
R670 B.n315 B.n15 10.6151
R671 B.n315 B.n314 10.6151
R672 B.n314 B.n313 10.6151
R673 B.n313 B.n16 10.6151
R674 B.n307 B.n16 10.6151
R675 B.n307 B.n306 10.6151
R676 B.n306 B.n305 10.6151
R677 B.n305 B.n22 10.6151
R678 B.n299 B.n22 10.6151
R679 B.n298 B.n297 10.6151
R680 B.n297 B.n30 10.6151
R681 B.n291 B.n30 10.6151
R682 B.n291 B.n290 10.6151
R683 B.n290 B.n289 10.6151
R684 B.n289 B.n32 10.6151
R685 B.n283 B.n32 10.6151
R686 B.n283 B.n282 10.6151
R687 B.n282 B.n281 10.6151
R688 B.n281 B.n34 10.6151
R689 B.n275 B.n34 10.6151
R690 B.n275 B.n274 10.6151
R691 B.n274 B.n273 10.6151
R692 B.n269 B.n268 10.6151
R693 B.n268 B.n40 10.6151
R694 B.n263 B.n40 10.6151
R695 B.n263 B.n262 10.6151
R696 B.n262 B.n261 10.6151
R697 B.n261 B.n42 10.6151
R698 B.n255 B.n42 10.6151
R699 B.n255 B.n254 10.6151
R700 B.n252 B.n46 10.6151
R701 B.n246 B.n46 10.6151
R702 B.n246 B.n245 10.6151
R703 B.n245 B.n244 10.6151
R704 B.n244 B.n48 10.6151
R705 B.n238 B.n48 10.6151
R706 B.n238 B.n237 10.6151
R707 B.n237 B.n236 10.6151
R708 B.n236 B.n50 10.6151
R709 B.n230 B.n50 10.6151
R710 B.n230 B.n229 10.6151
R711 B.n229 B.n228 10.6151
R712 B.n228 B.n224 10.6151
R713 B.n37 B.n36 10.0853
R714 B.n45 B.n44 10.0853
R715 B.n83 B.n82 10.0853
R716 B.n121 B.n120 10.0853
R717 B.n327 B.n0 8.11757
R718 B.n327 B.n1 8.11757
R719 B.n122 B.n89 7.18099
R720 B.n85 B.n84 7.18099
R721 B.n269 B.n38 7.18099
R722 B.n254 B.n253 7.18099
R723 B.n123 B.n122 3.43465
R724 B.n145 B.n84 3.43465
R725 B.n273 B.n38 3.43465
R726 B.n253 B.n252 3.43465
R727 VP.n1 VP.t2 525.049
R728 VP.n1 VP.t0 525.049
R729 VP.n0 VP.t1 525.049
R730 VP.n0 VP.t3 525.049
R731 VP.n2 VP.n0 193.006
R732 VP.n2 VP.n1 161.3
R733 VP VP.n2 0.0516364
R734 VDD1 VDD1.n1 115.466
R735 VDD1 VDD1.n0 87.7325
R736 VDD1.n0 VDD1.t2 7.79578
R737 VDD1.n0 VDD1.t0 7.79578
R738 VDD1.n1 VDD1.t3 7.79578
R739 VDD1.n1 VDD1.t1 7.79578
C0 VTAIL VDD1 3.3354f
C1 VP VDD2 0.248194f
C2 VDD2 VTAIL 3.37345f
C3 VP VN 2.70562f
C4 VTAIL VN 0.490589f
C5 VP VTAIL 0.504696f
C6 VDD2 VDD1 0.456355f
C7 VN VDD1 0.153553f
C8 VP VDD1 0.659275f
C9 VDD2 VN 0.565264f
C10 VDD2 B 1.652657f
C11 VDD1 B 3.85313f
C12 VTAIL B 2.885775f
C13 VN B 5.23989f
C14 VP B 3.073043f
C15 VDD1.t2 B 0.052523f
C16 VDD1.t0 B 0.052523f
C17 VDD1.n0 B 0.373331f
C18 VDD1.t3 B 0.052523f
C19 VDD1.t1 B 0.052523f
C20 VDD1.n1 B 0.598571f
C21 VP.t1 B 0.066046f
C22 VP.t3 B 0.066046f
C23 VP.n0 B 0.275289f
C24 VP.t0 B 0.066046f
C25 VP.t2 B 0.066046f
C26 VP.n1 B 0.095072f
C27 VP.n2 B 2.04958f
C28 VDD2.t0 B 0.055748f
C29 VDD2.t1 B 0.055748f
C30 VDD2.n0 B 0.618168f
C31 VDD2.t2 B 0.055748f
C32 VDD2.t3 B 0.055748f
C33 VDD2.n1 B 0.396076f
C34 VDD2.n2 B 2.11667f
C35 VTAIL.n0 B 0.029293f
C36 VTAIL.n1 B 0.164253f
C37 VTAIL.n2 B 0.011531f
C38 VTAIL.t4 B 0.047457f
C39 VTAIL.n3 B 0.076648f
C40 VTAIL.n4 B 0.015428f
C41 VTAIL.n5 B 0.020441f
C42 VTAIL.n6 B 0.057465f
C43 VTAIL.n7 B 0.012209f
C44 VTAIL.n8 B 0.011531f
C45 VTAIL.n9 B 0.053704f
C46 VTAIL.n10 B 0.032118f
C47 VTAIL.n11 B 0.072654f
C48 VTAIL.n12 B 0.029293f
C49 VTAIL.n13 B 0.164253f
C50 VTAIL.n14 B 0.011531f
C51 VTAIL.t3 B 0.047457f
C52 VTAIL.n15 B 0.076648f
C53 VTAIL.n16 B 0.015428f
C54 VTAIL.n17 B 0.020441f
C55 VTAIL.n18 B 0.057465f
C56 VTAIL.n19 B 0.012209f
C57 VTAIL.n20 B 0.011531f
C58 VTAIL.n21 B 0.053704f
C59 VTAIL.n22 B 0.032118f
C60 VTAIL.n23 B 0.084128f
C61 VTAIL.n24 B 0.029293f
C62 VTAIL.n25 B 0.164253f
C63 VTAIL.n26 B 0.011531f
C64 VTAIL.t2 B 0.047457f
C65 VTAIL.n27 B 0.076648f
C66 VTAIL.n28 B 0.015428f
C67 VTAIL.n29 B 0.020441f
C68 VTAIL.n30 B 0.057465f
C69 VTAIL.n31 B 0.012209f
C70 VTAIL.n32 B 0.011531f
C71 VTAIL.n33 B 0.053704f
C72 VTAIL.n34 B 0.032118f
C73 VTAIL.n35 B 0.526716f
C74 VTAIL.n36 B 0.029293f
C75 VTAIL.n37 B 0.164253f
C76 VTAIL.n38 B 0.011531f
C77 VTAIL.t5 B 0.047457f
C78 VTAIL.n39 B 0.076648f
C79 VTAIL.n40 B 0.015428f
C80 VTAIL.n41 B 0.020441f
C81 VTAIL.n42 B 0.057465f
C82 VTAIL.n43 B 0.012209f
C83 VTAIL.n44 B 0.011531f
C84 VTAIL.n45 B 0.053704f
C85 VTAIL.n46 B 0.032118f
C86 VTAIL.n47 B 0.526716f
C87 VTAIL.n48 B 0.029293f
C88 VTAIL.n49 B 0.164253f
C89 VTAIL.n50 B 0.011531f
C90 VTAIL.t7 B 0.047457f
C91 VTAIL.n51 B 0.076648f
C92 VTAIL.n52 B 0.015428f
C93 VTAIL.n53 B 0.020441f
C94 VTAIL.n54 B 0.057465f
C95 VTAIL.n55 B 0.012209f
C96 VTAIL.n56 B 0.011531f
C97 VTAIL.n57 B 0.053704f
C98 VTAIL.n58 B 0.032118f
C99 VTAIL.n59 B 0.084128f
C100 VTAIL.n60 B 0.029293f
C101 VTAIL.n61 B 0.164253f
C102 VTAIL.n62 B 0.011531f
C103 VTAIL.t0 B 0.047457f
C104 VTAIL.n63 B 0.076648f
C105 VTAIL.n64 B 0.015428f
C106 VTAIL.n65 B 0.020441f
C107 VTAIL.n66 B 0.057465f
C108 VTAIL.n67 B 0.012209f
C109 VTAIL.n68 B 0.011531f
C110 VTAIL.n69 B 0.053704f
C111 VTAIL.n70 B 0.032118f
C112 VTAIL.n71 B 0.084128f
C113 VTAIL.n72 B 0.029293f
C114 VTAIL.n73 B 0.164253f
C115 VTAIL.n74 B 0.011531f
C116 VTAIL.t1 B 0.047457f
C117 VTAIL.n75 B 0.076648f
C118 VTAIL.n76 B 0.015428f
C119 VTAIL.n77 B 0.020441f
C120 VTAIL.n78 B 0.057465f
C121 VTAIL.n79 B 0.012209f
C122 VTAIL.n80 B 0.011531f
C123 VTAIL.n81 B 0.053704f
C124 VTAIL.n82 B 0.032118f
C125 VTAIL.n83 B 0.526716f
C126 VTAIL.n84 B 0.029293f
C127 VTAIL.n85 B 0.164253f
C128 VTAIL.n86 B 0.011531f
C129 VTAIL.t6 B 0.047457f
C130 VTAIL.n87 B 0.076648f
C131 VTAIL.n88 B 0.015428f
C132 VTAIL.n89 B 0.020441f
C133 VTAIL.n90 B 0.057465f
C134 VTAIL.n91 B 0.012209f
C135 VTAIL.n92 B 0.011531f
C136 VTAIL.n93 B 0.053704f
C137 VTAIL.n94 B 0.032118f
C138 VTAIL.n95 B 0.507195f
C139 VN.t3 B 0.064542f
C140 VN.t2 B 0.064542f
C141 VN.n0 B 0.092919f
C142 VN.t1 B 0.064542f
C143 VN.t0 B 0.064542f
C144 VN.n1 B 0.275646f
.ends

