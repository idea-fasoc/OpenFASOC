* NGSPICE file created from diff_pair_sample_0578.ext - technology: sky130A

.subckt diff_pair_sample_0578 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=1.2837 pd=8.11 as=1.2837 ps=8.11 w=7.78 l=3.07
X1 VTAIL.t7 VP.t0 VDD1.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2837 pd=8.11 as=1.2837 ps=8.11 w=7.78 l=3.07
X2 VTAIL.t14 VN.t1 VDD2.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2837 pd=8.11 as=1.2837 ps=8.11 w=7.78 l=3.07
X3 VTAIL.t1 VP.t1 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=3.0342 pd=16.34 as=1.2837 ps=8.11 w=7.78 l=3.07
X4 VDD1.t5 VP.t2 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.2837 pd=8.11 as=3.0342 ps=16.34 w=7.78 l=3.07
X5 VTAIL.t5 VP.t3 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=3.0342 pd=16.34 as=1.2837 ps=8.11 w=7.78 l=3.07
X6 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=3.0342 pd=16.34 as=0 ps=0 w=7.78 l=3.07
X7 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=3.0342 pd=16.34 as=0 ps=0 w=7.78 l=3.07
X8 VDD2.t3 VN.t2 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2837 pd=8.11 as=1.2837 ps=8.11 w=7.78 l=3.07
X9 VTAIL.t12 VN.t3 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=3.0342 pd=16.34 as=1.2837 ps=8.11 w=7.78 l=3.07
X10 VTAIL.t11 VN.t4 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=3.0342 pd=16.34 as=1.2837 ps=8.11 w=7.78 l=3.07
X11 VDD1.t3 VP.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2837 pd=8.11 as=1.2837 ps=8.11 w=7.78 l=3.07
X12 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=3.0342 pd=16.34 as=0 ps=0 w=7.78 l=3.07
X13 VDD2.t6 VN.t5 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=1.2837 pd=8.11 as=1.2837 ps=8.11 w=7.78 l=3.07
X14 VDD2.t5 VN.t6 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2837 pd=8.11 as=3.0342 ps=16.34 w=7.78 l=3.07
X15 VDD2.t7 VN.t7 VTAIL.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=1.2837 pd=8.11 as=3.0342 ps=16.34 w=7.78 l=3.07
X16 VDD1.t2 VP.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.2837 pd=8.11 as=1.2837 ps=8.11 w=7.78 l=3.07
X17 VTAIL.t2 VP.t6 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.2837 pd=8.11 as=1.2837 ps=8.11 w=7.78 l=3.07
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.0342 pd=16.34 as=0 ps=0 w=7.78 l=3.07
X19 VDD1.t0 VP.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2837 pd=8.11 as=3.0342 ps=16.34 w=7.78 l=3.07
R0 VN.n60 VN.n59 161.3
R1 VN.n58 VN.n32 161.3
R2 VN.n57 VN.n56 161.3
R3 VN.n55 VN.n33 161.3
R4 VN.n54 VN.n53 161.3
R5 VN.n52 VN.n34 161.3
R6 VN.n51 VN.n50 161.3
R7 VN.n49 VN.n48 161.3
R8 VN.n47 VN.n36 161.3
R9 VN.n46 VN.n45 161.3
R10 VN.n44 VN.n37 161.3
R11 VN.n43 VN.n42 161.3
R12 VN.n41 VN.n38 161.3
R13 VN.n29 VN.n28 161.3
R14 VN.n27 VN.n1 161.3
R15 VN.n26 VN.n25 161.3
R16 VN.n24 VN.n2 161.3
R17 VN.n23 VN.n22 161.3
R18 VN.n21 VN.n3 161.3
R19 VN.n20 VN.n19 161.3
R20 VN.n18 VN.n17 161.3
R21 VN.n16 VN.n5 161.3
R22 VN.n15 VN.n14 161.3
R23 VN.n13 VN.n6 161.3
R24 VN.n12 VN.n11 161.3
R25 VN.n10 VN.n7 161.3
R26 VN.n8 VN.t4 94.2636
R27 VN.n39 VN.t7 94.2636
R28 VN.n30 VN.n0 72.8506
R29 VN.n61 VN.n31 72.8506
R30 VN.n9 VN.t2 61.0748
R31 VN.n4 VN.t0 61.0748
R32 VN.n0 VN.t6 61.0748
R33 VN.n40 VN.t1 61.0748
R34 VN.n35 VN.t5 61.0748
R35 VN.n31 VN.t3 61.0748
R36 VN.n15 VN.n6 56.4773
R37 VN.n46 VN.n37 56.4773
R38 VN.n26 VN.n2 55.0167
R39 VN.n57 VN.n33 55.0167
R40 VN.n9 VN.n8 51.6654
R41 VN.n40 VN.n39 51.6654
R42 VN VN.n61 50.157
R43 VN.n22 VN.n2 25.8045
R44 VN.n53 VN.n33 25.8045
R45 VN.n11 VN.n10 24.3439
R46 VN.n11 VN.n6 24.3439
R47 VN.n16 VN.n15 24.3439
R48 VN.n17 VN.n16 24.3439
R49 VN.n21 VN.n20 24.3439
R50 VN.n22 VN.n21 24.3439
R51 VN.n27 VN.n26 24.3439
R52 VN.n28 VN.n27 24.3439
R53 VN.n42 VN.n37 24.3439
R54 VN.n42 VN.n41 24.3439
R55 VN.n53 VN.n52 24.3439
R56 VN.n52 VN.n51 24.3439
R57 VN.n48 VN.n47 24.3439
R58 VN.n47 VN.n46 24.3439
R59 VN.n59 VN.n58 24.3439
R60 VN.n58 VN.n57 24.3439
R61 VN.n10 VN.n9 21.9096
R62 VN.n17 VN.n4 21.9096
R63 VN.n41 VN.n40 21.9096
R64 VN.n48 VN.n35 21.9096
R65 VN.n28 VN.n0 17.0409
R66 VN.n59 VN.n31 17.0409
R67 VN.n39 VN.n38 4.06494
R68 VN.n8 VN.n7 4.06494
R69 VN.n20 VN.n4 2.43484
R70 VN.n51 VN.n35 2.43484
R71 VN.n61 VN.n60 0.355081
R72 VN.n30 VN.n29 0.355081
R73 VN VN.n30 0.26685
R74 VN.n60 VN.n32 0.189894
R75 VN.n56 VN.n32 0.189894
R76 VN.n56 VN.n55 0.189894
R77 VN.n55 VN.n54 0.189894
R78 VN.n54 VN.n34 0.189894
R79 VN.n50 VN.n34 0.189894
R80 VN.n50 VN.n49 0.189894
R81 VN.n49 VN.n36 0.189894
R82 VN.n45 VN.n36 0.189894
R83 VN.n45 VN.n44 0.189894
R84 VN.n44 VN.n43 0.189894
R85 VN.n43 VN.n38 0.189894
R86 VN.n12 VN.n7 0.189894
R87 VN.n13 VN.n12 0.189894
R88 VN.n14 VN.n13 0.189894
R89 VN.n14 VN.n5 0.189894
R90 VN.n18 VN.n5 0.189894
R91 VN.n19 VN.n18 0.189894
R92 VN.n19 VN.n3 0.189894
R93 VN.n23 VN.n3 0.189894
R94 VN.n24 VN.n23 0.189894
R95 VN.n25 VN.n24 0.189894
R96 VN.n25 VN.n1 0.189894
R97 VN.n29 VN.n1 0.189894
R98 VDD2.n2 VDD2.n1 65.8549
R99 VDD2.n2 VDD2.n0 65.8549
R100 VDD2 VDD2.n5 65.8521
R101 VDD2.n4 VDD2.n3 64.4447
R102 VDD2.n4 VDD2.n2 43.6118
R103 VDD2.n5 VDD2.t0 2.54549
R104 VDD2.n5 VDD2.t7 2.54549
R105 VDD2.n3 VDD2.t2 2.54549
R106 VDD2.n3 VDD2.t6 2.54549
R107 VDD2.n1 VDD2.t4 2.54549
R108 VDD2.n1 VDD2.t5 2.54549
R109 VDD2.n0 VDD2.t1 2.54549
R110 VDD2.n0 VDD2.t3 2.54549
R111 VDD2 VDD2.n4 1.52421
R112 VTAIL.n14 VTAIL.t0 50.3109
R113 VTAIL.n11 VTAIL.t5 50.3109
R114 VTAIL.n10 VTAIL.t8 50.3109
R115 VTAIL.n7 VTAIL.t12 50.3109
R116 VTAIL.n15 VTAIL.t9 50.3108
R117 VTAIL.n2 VTAIL.t11 50.3108
R118 VTAIL.n3 VTAIL.t6 50.3108
R119 VTAIL.n6 VTAIL.t1 50.3108
R120 VTAIL.n13 VTAIL.n12 47.766
R121 VTAIL.n9 VTAIL.n8 47.766
R122 VTAIL.n1 VTAIL.n0 47.7659
R123 VTAIL.n5 VTAIL.n4 47.7659
R124 VTAIL.n15 VTAIL.n14 22.0048
R125 VTAIL.n7 VTAIL.n6 22.0048
R126 VTAIL.n9 VTAIL.n7 2.93153
R127 VTAIL.n10 VTAIL.n9 2.93153
R128 VTAIL.n13 VTAIL.n11 2.93153
R129 VTAIL.n14 VTAIL.n13 2.93153
R130 VTAIL.n6 VTAIL.n5 2.93153
R131 VTAIL.n5 VTAIL.n3 2.93153
R132 VTAIL.n2 VTAIL.n1 2.93153
R133 VTAIL VTAIL.n15 2.87334
R134 VTAIL.n0 VTAIL.t13 2.54549
R135 VTAIL.n0 VTAIL.t15 2.54549
R136 VTAIL.n4 VTAIL.t4 2.54549
R137 VTAIL.n4 VTAIL.t7 2.54549
R138 VTAIL.n12 VTAIL.t3 2.54549
R139 VTAIL.n12 VTAIL.t2 2.54549
R140 VTAIL.n8 VTAIL.t10 2.54549
R141 VTAIL.n8 VTAIL.t14 2.54549
R142 VTAIL.n11 VTAIL.n10 0.470328
R143 VTAIL.n3 VTAIL.n2 0.470328
R144 VTAIL VTAIL.n1 0.0586897
R145 B.n683 B.n682 585
R146 B.n685 B.n145 585
R147 B.n688 B.n687 585
R148 B.n689 B.n144 585
R149 B.n691 B.n690 585
R150 B.n693 B.n143 585
R151 B.n696 B.n695 585
R152 B.n697 B.n142 585
R153 B.n699 B.n698 585
R154 B.n701 B.n141 585
R155 B.n704 B.n703 585
R156 B.n705 B.n140 585
R157 B.n707 B.n706 585
R158 B.n709 B.n139 585
R159 B.n712 B.n711 585
R160 B.n713 B.n138 585
R161 B.n715 B.n714 585
R162 B.n717 B.n137 585
R163 B.n720 B.n719 585
R164 B.n721 B.n136 585
R165 B.n723 B.n722 585
R166 B.n725 B.n135 585
R167 B.n728 B.n727 585
R168 B.n729 B.n134 585
R169 B.n731 B.n730 585
R170 B.n733 B.n133 585
R171 B.n736 B.n735 585
R172 B.n737 B.n129 585
R173 B.n739 B.n738 585
R174 B.n741 B.n128 585
R175 B.n744 B.n743 585
R176 B.n745 B.n127 585
R177 B.n747 B.n746 585
R178 B.n749 B.n126 585
R179 B.n752 B.n751 585
R180 B.n753 B.n125 585
R181 B.n755 B.n754 585
R182 B.n757 B.n124 585
R183 B.n760 B.n759 585
R184 B.n762 B.n121 585
R185 B.n764 B.n763 585
R186 B.n766 B.n120 585
R187 B.n769 B.n768 585
R188 B.n770 B.n119 585
R189 B.n772 B.n771 585
R190 B.n774 B.n118 585
R191 B.n777 B.n776 585
R192 B.n778 B.n117 585
R193 B.n780 B.n779 585
R194 B.n782 B.n116 585
R195 B.n785 B.n784 585
R196 B.n786 B.n115 585
R197 B.n788 B.n787 585
R198 B.n790 B.n114 585
R199 B.n793 B.n792 585
R200 B.n794 B.n113 585
R201 B.n796 B.n795 585
R202 B.n798 B.n112 585
R203 B.n801 B.n800 585
R204 B.n802 B.n111 585
R205 B.n804 B.n803 585
R206 B.n806 B.n110 585
R207 B.n809 B.n808 585
R208 B.n810 B.n109 585
R209 B.n812 B.n811 585
R210 B.n814 B.n108 585
R211 B.n817 B.n816 585
R212 B.n818 B.n107 585
R213 B.n681 B.n105 585
R214 B.n821 B.n105 585
R215 B.n680 B.n104 585
R216 B.n822 B.n104 585
R217 B.n679 B.n103 585
R218 B.n823 B.n103 585
R219 B.n678 B.n677 585
R220 B.n677 B.n99 585
R221 B.n676 B.n98 585
R222 B.n829 B.n98 585
R223 B.n675 B.n97 585
R224 B.n830 B.n97 585
R225 B.n674 B.n96 585
R226 B.n831 B.n96 585
R227 B.n673 B.n672 585
R228 B.n672 B.n92 585
R229 B.n671 B.n91 585
R230 B.n837 B.n91 585
R231 B.n670 B.n90 585
R232 B.n838 B.n90 585
R233 B.n669 B.n89 585
R234 B.n839 B.n89 585
R235 B.n668 B.n667 585
R236 B.n667 B.n85 585
R237 B.n666 B.n84 585
R238 B.n845 B.n84 585
R239 B.n665 B.n83 585
R240 B.n846 B.n83 585
R241 B.n664 B.n82 585
R242 B.n847 B.n82 585
R243 B.n663 B.n662 585
R244 B.n662 B.n78 585
R245 B.n661 B.n77 585
R246 B.n853 B.n77 585
R247 B.n660 B.n76 585
R248 B.n854 B.n76 585
R249 B.n659 B.n75 585
R250 B.n855 B.n75 585
R251 B.n658 B.n657 585
R252 B.n657 B.n71 585
R253 B.n656 B.n70 585
R254 B.n861 B.n70 585
R255 B.n655 B.n69 585
R256 B.n862 B.n69 585
R257 B.n654 B.n68 585
R258 B.n863 B.n68 585
R259 B.n653 B.n652 585
R260 B.n652 B.n64 585
R261 B.n651 B.n63 585
R262 B.n869 B.n63 585
R263 B.n650 B.n62 585
R264 B.n870 B.n62 585
R265 B.n649 B.n61 585
R266 B.n871 B.n61 585
R267 B.n648 B.n647 585
R268 B.n647 B.n57 585
R269 B.n646 B.n56 585
R270 B.n877 B.n56 585
R271 B.n645 B.n55 585
R272 B.n878 B.n55 585
R273 B.n644 B.n54 585
R274 B.n879 B.n54 585
R275 B.n643 B.n642 585
R276 B.n642 B.n53 585
R277 B.n641 B.n49 585
R278 B.n885 B.n49 585
R279 B.n640 B.n48 585
R280 B.n886 B.n48 585
R281 B.n639 B.n47 585
R282 B.n887 B.n47 585
R283 B.n638 B.n637 585
R284 B.n637 B.n43 585
R285 B.n636 B.n42 585
R286 B.n893 B.n42 585
R287 B.n635 B.n41 585
R288 B.n894 B.n41 585
R289 B.n634 B.n40 585
R290 B.n895 B.n40 585
R291 B.n633 B.n632 585
R292 B.n632 B.n36 585
R293 B.n631 B.n35 585
R294 B.n901 B.n35 585
R295 B.n630 B.n34 585
R296 B.n902 B.n34 585
R297 B.n629 B.n33 585
R298 B.n903 B.n33 585
R299 B.n628 B.n627 585
R300 B.n627 B.n29 585
R301 B.n626 B.n28 585
R302 B.n909 B.n28 585
R303 B.n625 B.n27 585
R304 B.n910 B.n27 585
R305 B.n624 B.n26 585
R306 B.n911 B.n26 585
R307 B.n623 B.n622 585
R308 B.n622 B.n22 585
R309 B.n621 B.n21 585
R310 B.n917 B.n21 585
R311 B.n620 B.n20 585
R312 B.n918 B.n20 585
R313 B.n619 B.n19 585
R314 B.n919 B.n19 585
R315 B.n618 B.n617 585
R316 B.n617 B.n18 585
R317 B.n616 B.n14 585
R318 B.n925 B.n14 585
R319 B.n615 B.n13 585
R320 B.n926 B.n13 585
R321 B.n614 B.n12 585
R322 B.n927 B.n12 585
R323 B.n613 B.n612 585
R324 B.n612 B.n8 585
R325 B.n611 B.n7 585
R326 B.n933 B.n7 585
R327 B.n610 B.n6 585
R328 B.n934 B.n6 585
R329 B.n609 B.n5 585
R330 B.n935 B.n5 585
R331 B.n608 B.n607 585
R332 B.n607 B.n4 585
R333 B.n606 B.n146 585
R334 B.n606 B.n605 585
R335 B.n596 B.n147 585
R336 B.n148 B.n147 585
R337 B.n598 B.n597 585
R338 B.n599 B.n598 585
R339 B.n595 B.n153 585
R340 B.n153 B.n152 585
R341 B.n594 B.n593 585
R342 B.n593 B.n592 585
R343 B.n155 B.n154 585
R344 B.n585 B.n155 585
R345 B.n584 B.n583 585
R346 B.n586 B.n584 585
R347 B.n582 B.n160 585
R348 B.n160 B.n159 585
R349 B.n581 B.n580 585
R350 B.n580 B.n579 585
R351 B.n162 B.n161 585
R352 B.n163 B.n162 585
R353 B.n572 B.n571 585
R354 B.n573 B.n572 585
R355 B.n570 B.n168 585
R356 B.n168 B.n167 585
R357 B.n569 B.n568 585
R358 B.n568 B.n567 585
R359 B.n170 B.n169 585
R360 B.n171 B.n170 585
R361 B.n560 B.n559 585
R362 B.n561 B.n560 585
R363 B.n558 B.n175 585
R364 B.n179 B.n175 585
R365 B.n557 B.n556 585
R366 B.n556 B.n555 585
R367 B.n177 B.n176 585
R368 B.n178 B.n177 585
R369 B.n548 B.n547 585
R370 B.n549 B.n548 585
R371 B.n546 B.n184 585
R372 B.n184 B.n183 585
R373 B.n545 B.n544 585
R374 B.n544 B.n543 585
R375 B.n186 B.n185 585
R376 B.n187 B.n186 585
R377 B.n536 B.n535 585
R378 B.n537 B.n536 585
R379 B.n534 B.n192 585
R380 B.n192 B.n191 585
R381 B.n533 B.n532 585
R382 B.n532 B.n531 585
R383 B.n194 B.n193 585
R384 B.n524 B.n194 585
R385 B.n523 B.n522 585
R386 B.n525 B.n523 585
R387 B.n521 B.n199 585
R388 B.n199 B.n198 585
R389 B.n520 B.n519 585
R390 B.n519 B.n518 585
R391 B.n201 B.n200 585
R392 B.n202 B.n201 585
R393 B.n511 B.n510 585
R394 B.n512 B.n511 585
R395 B.n509 B.n207 585
R396 B.n207 B.n206 585
R397 B.n508 B.n507 585
R398 B.n507 B.n506 585
R399 B.n209 B.n208 585
R400 B.n210 B.n209 585
R401 B.n499 B.n498 585
R402 B.n500 B.n499 585
R403 B.n497 B.n214 585
R404 B.n218 B.n214 585
R405 B.n496 B.n495 585
R406 B.n495 B.n494 585
R407 B.n216 B.n215 585
R408 B.n217 B.n216 585
R409 B.n487 B.n486 585
R410 B.n488 B.n487 585
R411 B.n485 B.n223 585
R412 B.n223 B.n222 585
R413 B.n484 B.n483 585
R414 B.n483 B.n482 585
R415 B.n225 B.n224 585
R416 B.n226 B.n225 585
R417 B.n475 B.n474 585
R418 B.n476 B.n475 585
R419 B.n473 B.n231 585
R420 B.n231 B.n230 585
R421 B.n472 B.n471 585
R422 B.n471 B.n470 585
R423 B.n233 B.n232 585
R424 B.n234 B.n233 585
R425 B.n463 B.n462 585
R426 B.n464 B.n463 585
R427 B.n461 B.n239 585
R428 B.n239 B.n238 585
R429 B.n460 B.n459 585
R430 B.n459 B.n458 585
R431 B.n241 B.n240 585
R432 B.n242 B.n241 585
R433 B.n451 B.n450 585
R434 B.n452 B.n451 585
R435 B.n449 B.n247 585
R436 B.n247 B.n246 585
R437 B.n448 B.n447 585
R438 B.n447 B.n446 585
R439 B.n249 B.n248 585
R440 B.n250 B.n249 585
R441 B.n439 B.n438 585
R442 B.n440 B.n439 585
R443 B.n437 B.n255 585
R444 B.n255 B.n254 585
R445 B.n436 B.n435 585
R446 B.n435 B.n434 585
R447 B.n431 B.n259 585
R448 B.n430 B.n429 585
R449 B.n427 B.n260 585
R450 B.n427 B.n258 585
R451 B.n426 B.n425 585
R452 B.n424 B.n423 585
R453 B.n422 B.n262 585
R454 B.n420 B.n419 585
R455 B.n418 B.n263 585
R456 B.n417 B.n416 585
R457 B.n414 B.n264 585
R458 B.n412 B.n411 585
R459 B.n410 B.n265 585
R460 B.n409 B.n408 585
R461 B.n406 B.n266 585
R462 B.n404 B.n403 585
R463 B.n402 B.n267 585
R464 B.n401 B.n400 585
R465 B.n398 B.n268 585
R466 B.n396 B.n395 585
R467 B.n394 B.n269 585
R468 B.n393 B.n392 585
R469 B.n390 B.n270 585
R470 B.n388 B.n387 585
R471 B.n386 B.n271 585
R472 B.n385 B.n384 585
R473 B.n382 B.n272 585
R474 B.n380 B.n379 585
R475 B.n378 B.n273 585
R476 B.n377 B.n376 585
R477 B.n374 B.n373 585
R478 B.n372 B.n371 585
R479 B.n370 B.n278 585
R480 B.n368 B.n367 585
R481 B.n366 B.n279 585
R482 B.n365 B.n364 585
R483 B.n362 B.n280 585
R484 B.n360 B.n359 585
R485 B.n358 B.n281 585
R486 B.n357 B.n356 585
R487 B.n354 B.n353 585
R488 B.n352 B.n351 585
R489 B.n350 B.n286 585
R490 B.n348 B.n347 585
R491 B.n346 B.n287 585
R492 B.n345 B.n344 585
R493 B.n342 B.n288 585
R494 B.n340 B.n339 585
R495 B.n338 B.n289 585
R496 B.n337 B.n336 585
R497 B.n334 B.n290 585
R498 B.n332 B.n331 585
R499 B.n330 B.n291 585
R500 B.n329 B.n328 585
R501 B.n326 B.n292 585
R502 B.n324 B.n323 585
R503 B.n322 B.n293 585
R504 B.n321 B.n320 585
R505 B.n318 B.n294 585
R506 B.n316 B.n315 585
R507 B.n314 B.n295 585
R508 B.n313 B.n312 585
R509 B.n310 B.n296 585
R510 B.n308 B.n307 585
R511 B.n306 B.n297 585
R512 B.n305 B.n304 585
R513 B.n302 B.n298 585
R514 B.n300 B.n299 585
R515 B.n257 B.n256 585
R516 B.n258 B.n257 585
R517 B.n433 B.n432 585
R518 B.n434 B.n433 585
R519 B.n253 B.n252 585
R520 B.n254 B.n253 585
R521 B.n442 B.n441 585
R522 B.n441 B.n440 585
R523 B.n443 B.n251 585
R524 B.n251 B.n250 585
R525 B.n445 B.n444 585
R526 B.n446 B.n445 585
R527 B.n245 B.n244 585
R528 B.n246 B.n245 585
R529 B.n454 B.n453 585
R530 B.n453 B.n452 585
R531 B.n455 B.n243 585
R532 B.n243 B.n242 585
R533 B.n457 B.n456 585
R534 B.n458 B.n457 585
R535 B.n237 B.n236 585
R536 B.n238 B.n237 585
R537 B.n466 B.n465 585
R538 B.n465 B.n464 585
R539 B.n467 B.n235 585
R540 B.n235 B.n234 585
R541 B.n469 B.n468 585
R542 B.n470 B.n469 585
R543 B.n229 B.n228 585
R544 B.n230 B.n229 585
R545 B.n478 B.n477 585
R546 B.n477 B.n476 585
R547 B.n479 B.n227 585
R548 B.n227 B.n226 585
R549 B.n481 B.n480 585
R550 B.n482 B.n481 585
R551 B.n221 B.n220 585
R552 B.n222 B.n221 585
R553 B.n490 B.n489 585
R554 B.n489 B.n488 585
R555 B.n491 B.n219 585
R556 B.n219 B.n217 585
R557 B.n493 B.n492 585
R558 B.n494 B.n493 585
R559 B.n213 B.n212 585
R560 B.n218 B.n213 585
R561 B.n502 B.n501 585
R562 B.n501 B.n500 585
R563 B.n503 B.n211 585
R564 B.n211 B.n210 585
R565 B.n505 B.n504 585
R566 B.n506 B.n505 585
R567 B.n205 B.n204 585
R568 B.n206 B.n205 585
R569 B.n514 B.n513 585
R570 B.n513 B.n512 585
R571 B.n515 B.n203 585
R572 B.n203 B.n202 585
R573 B.n517 B.n516 585
R574 B.n518 B.n517 585
R575 B.n197 B.n196 585
R576 B.n198 B.n197 585
R577 B.n527 B.n526 585
R578 B.n526 B.n525 585
R579 B.n528 B.n195 585
R580 B.n524 B.n195 585
R581 B.n530 B.n529 585
R582 B.n531 B.n530 585
R583 B.n190 B.n189 585
R584 B.n191 B.n190 585
R585 B.n539 B.n538 585
R586 B.n538 B.n537 585
R587 B.n540 B.n188 585
R588 B.n188 B.n187 585
R589 B.n542 B.n541 585
R590 B.n543 B.n542 585
R591 B.n182 B.n181 585
R592 B.n183 B.n182 585
R593 B.n551 B.n550 585
R594 B.n550 B.n549 585
R595 B.n552 B.n180 585
R596 B.n180 B.n178 585
R597 B.n554 B.n553 585
R598 B.n555 B.n554 585
R599 B.n174 B.n173 585
R600 B.n179 B.n174 585
R601 B.n563 B.n562 585
R602 B.n562 B.n561 585
R603 B.n564 B.n172 585
R604 B.n172 B.n171 585
R605 B.n566 B.n565 585
R606 B.n567 B.n566 585
R607 B.n166 B.n165 585
R608 B.n167 B.n166 585
R609 B.n575 B.n574 585
R610 B.n574 B.n573 585
R611 B.n576 B.n164 585
R612 B.n164 B.n163 585
R613 B.n578 B.n577 585
R614 B.n579 B.n578 585
R615 B.n158 B.n157 585
R616 B.n159 B.n158 585
R617 B.n588 B.n587 585
R618 B.n587 B.n586 585
R619 B.n589 B.n156 585
R620 B.n585 B.n156 585
R621 B.n591 B.n590 585
R622 B.n592 B.n591 585
R623 B.n151 B.n150 585
R624 B.n152 B.n151 585
R625 B.n601 B.n600 585
R626 B.n600 B.n599 585
R627 B.n602 B.n149 585
R628 B.n149 B.n148 585
R629 B.n604 B.n603 585
R630 B.n605 B.n604 585
R631 B.n2 B.n0 585
R632 B.n4 B.n2 585
R633 B.n3 B.n1 585
R634 B.n934 B.n3 585
R635 B.n932 B.n931 585
R636 B.n933 B.n932 585
R637 B.n930 B.n9 585
R638 B.n9 B.n8 585
R639 B.n929 B.n928 585
R640 B.n928 B.n927 585
R641 B.n11 B.n10 585
R642 B.n926 B.n11 585
R643 B.n924 B.n923 585
R644 B.n925 B.n924 585
R645 B.n922 B.n15 585
R646 B.n18 B.n15 585
R647 B.n921 B.n920 585
R648 B.n920 B.n919 585
R649 B.n17 B.n16 585
R650 B.n918 B.n17 585
R651 B.n916 B.n915 585
R652 B.n917 B.n916 585
R653 B.n914 B.n23 585
R654 B.n23 B.n22 585
R655 B.n913 B.n912 585
R656 B.n912 B.n911 585
R657 B.n25 B.n24 585
R658 B.n910 B.n25 585
R659 B.n908 B.n907 585
R660 B.n909 B.n908 585
R661 B.n906 B.n30 585
R662 B.n30 B.n29 585
R663 B.n905 B.n904 585
R664 B.n904 B.n903 585
R665 B.n32 B.n31 585
R666 B.n902 B.n32 585
R667 B.n900 B.n899 585
R668 B.n901 B.n900 585
R669 B.n898 B.n37 585
R670 B.n37 B.n36 585
R671 B.n897 B.n896 585
R672 B.n896 B.n895 585
R673 B.n39 B.n38 585
R674 B.n894 B.n39 585
R675 B.n892 B.n891 585
R676 B.n893 B.n892 585
R677 B.n890 B.n44 585
R678 B.n44 B.n43 585
R679 B.n889 B.n888 585
R680 B.n888 B.n887 585
R681 B.n46 B.n45 585
R682 B.n886 B.n46 585
R683 B.n884 B.n883 585
R684 B.n885 B.n884 585
R685 B.n882 B.n50 585
R686 B.n53 B.n50 585
R687 B.n881 B.n880 585
R688 B.n880 B.n879 585
R689 B.n52 B.n51 585
R690 B.n878 B.n52 585
R691 B.n876 B.n875 585
R692 B.n877 B.n876 585
R693 B.n874 B.n58 585
R694 B.n58 B.n57 585
R695 B.n873 B.n872 585
R696 B.n872 B.n871 585
R697 B.n60 B.n59 585
R698 B.n870 B.n60 585
R699 B.n868 B.n867 585
R700 B.n869 B.n868 585
R701 B.n866 B.n65 585
R702 B.n65 B.n64 585
R703 B.n865 B.n864 585
R704 B.n864 B.n863 585
R705 B.n67 B.n66 585
R706 B.n862 B.n67 585
R707 B.n860 B.n859 585
R708 B.n861 B.n860 585
R709 B.n858 B.n72 585
R710 B.n72 B.n71 585
R711 B.n857 B.n856 585
R712 B.n856 B.n855 585
R713 B.n74 B.n73 585
R714 B.n854 B.n74 585
R715 B.n852 B.n851 585
R716 B.n853 B.n852 585
R717 B.n850 B.n79 585
R718 B.n79 B.n78 585
R719 B.n849 B.n848 585
R720 B.n848 B.n847 585
R721 B.n81 B.n80 585
R722 B.n846 B.n81 585
R723 B.n844 B.n843 585
R724 B.n845 B.n844 585
R725 B.n842 B.n86 585
R726 B.n86 B.n85 585
R727 B.n841 B.n840 585
R728 B.n840 B.n839 585
R729 B.n88 B.n87 585
R730 B.n838 B.n88 585
R731 B.n836 B.n835 585
R732 B.n837 B.n836 585
R733 B.n834 B.n93 585
R734 B.n93 B.n92 585
R735 B.n833 B.n832 585
R736 B.n832 B.n831 585
R737 B.n95 B.n94 585
R738 B.n830 B.n95 585
R739 B.n828 B.n827 585
R740 B.n829 B.n828 585
R741 B.n826 B.n100 585
R742 B.n100 B.n99 585
R743 B.n825 B.n824 585
R744 B.n824 B.n823 585
R745 B.n102 B.n101 585
R746 B.n822 B.n102 585
R747 B.n820 B.n819 585
R748 B.n821 B.n820 585
R749 B.n937 B.n936 585
R750 B.n936 B.n935 585
R751 B.n433 B.n259 516.524
R752 B.n820 B.n107 516.524
R753 B.n435 B.n257 516.524
R754 B.n683 B.n105 516.524
R755 B.n282 B.t8 270.404
R756 B.n130 B.t16 270.404
R757 B.n274 B.t19 270.115
R758 B.n122 B.t12 270.115
R759 B.n684 B.n106 256.663
R760 B.n686 B.n106 256.663
R761 B.n692 B.n106 256.663
R762 B.n694 B.n106 256.663
R763 B.n700 B.n106 256.663
R764 B.n702 B.n106 256.663
R765 B.n708 B.n106 256.663
R766 B.n710 B.n106 256.663
R767 B.n716 B.n106 256.663
R768 B.n718 B.n106 256.663
R769 B.n724 B.n106 256.663
R770 B.n726 B.n106 256.663
R771 B.n732 B.n106 256.663
R772 B.n734 B.n106 256.663
R773 B.n740 B.n106 256.663
R774 B.n742 B.n106 256.663
R775 B.n748 B.n106 256.663
R776 B.n750 B.n106 256.663
R777 B.n756 B.n106 256.663
R778 B.n758 B.n106 256.663
R779 B.n765 B.n106 256.663
R780 B.n767 B.n106 256.663
R781 B.n773 B.n106 256.663
R782 B.n775 B.n106 256.663
R783 B.n781 B.n106 256.663
R784 B.n783 B.n106 256.663
R785 B.n789 B.n106 256.663
R786 B.n791 B.n106 256.663
R787 B.n797 B.n106 256.663
R788 B.n799 B.n106 256.663
R789 B.n805 B.n106 256.663
R790 B.n807 B.n106 256.663
R791 B.n813 B.n106 256.663
R792 B.n815 B.n106 256.663
R793 B.n428 B.n258 256.663
R794 B.n261 B.n258 256.663
R795 B.n421 B.n258 256.663
R796 B.n415 B.n258 256.663
R797 B.n413 B.n258 256.663
R798 B.n407 B.n258 256.663
R799 B.n405 B.n258 256.663
R800 B.n399 B.n258 256.663
R801 B.n397 B.n258 256.663
R802 B.n391 B.n258 256.663
R803 B.n389 B.n258 256.663
R804 B.n383 B.n258 256.663
R805 B.n381 B.n258 256.663
R806 B.n375 B.n258 256.663
R807 B.n277 B.n258 256.663
R808 B.n369 B.n258 256.663
R809 B.n363 B.n258 256.663
R810 B.n361 B.n258 256.663
R811 B.n355 B.n258 256.663
R812 B.n285 B.n258 256.663
R813 B.n349 B.n258 256.663
R814 B.n343 B.n258 256.663
R815 B.n341 B.n258 256.663
R816 B.n335 B.n258 256.663
R817 B.n333 B.n258 256.663
R818 B.n327 B.n258 256.663
R819 B.n325 B.n258 256.663
R820 B.n319 B.n258 256.663
R821 B.n317 B.n258 256.663
R822 B.n311 B.n258 256.663
R823 B.n309 B.n258 256.663
R824 B.n303 B.n258 256.663
R825 B.n301 B.n258 256.663
R826 B.n433 B.n253 163.367
R827 B.n441 B.n253 163.367
R828 B.n441 B.n251 163.367
R829 B.n445 B.n251 163.367
R830 B.n445 B.n245 163.367
R831 B.n453 B.n245 163.367
R832 B.n453 B.n243 163.367
R833 B.n457 B.n243 163.367
R834 B.n457 B.n237 163.367
R835 B.n465 B.n237 163.367
R836 B.n465 B.n235 163.367
R837 B.n469 B.n235 163.367
R838 B.n469 B.n229 163.367
R839 B.n477 B.n229 163.367
R840 B.n477 B.n227 163.367
R841 B.n481 B.n227 163.367
R842 B.n481 B.n221 163.367
R843 B.n489 B.n221 163.367
R844 B.n489 B.n219 163.367
R845 B.n493 B.n219 163.367
R846 B.n493 B.n213 163.367
R847 B.n501 B.n213 163.367
R848 B.n501 B.n211 163.367
R849 B.n505 B.n211 163.367
R850 B.n505 B.n205 163.367
R851 B.n513 B.n205 163.367
R852 B.n513 B.n203 163.367
R853 B.n517 B.n203 163.367
R854 B.n517 B.n197 163.367
R855 B.n526 B.n197 163.367
R856 B.n526 B.n195 163.367
R857 B.n530 B.n195 163.367
R858 B.n530 B.n190 163.367
R859 B.n538 B.n190 163.367
R860 B.n538 B.n188 163.367
R861 B.n542 B.n188 163.367
R862 B.n542 B.n182 163.367
R863 B.n550 B.n182 163.367
R864 B.n550 B.n180 163.367
R865 B.n554 B.n180 163.367
R866 B.n554 B.n174 163.367
R867 B.n562 B.n174 163.367
R868 B.n562 B.n172 163.367
R869 B.n566 B.n172 163.367
R870 B.n566 B.n166 163.367
R871 B.n574 B.n166 163.367
R872 B.n574 B.n164 163.367
R873 B.n578 B.n164 163.367
R874 B.n578 B.n158 163.367
R875 B.n587 B.n158 163.367
R876 B.n587 B.n156 163.367
R877 B.n591 B.n156 163.367
R878 B.n591 B.n151 163.367
R879 B.n600 B.n151 163.367
R880 B.n600 B.n149 163.367
R881 B.n604 B.n149 163.367
R882 B.n604 B.n2 163.367
R883 B.n936 B.n2 163.367
R884 B.n936 B.n3 163.367
R885 B.n932 B.n3 163.367
R886 B.n932 B.n9 163.367
R887 B.n928 B.n9 163.367
R888 B.n928 B.n11 163.367
R889 B.n924 B.n11 163.367
R890 B.n924 B.n15 163.367
R891 B.n920 B.n15 163.367
R892 B.n920 B.n17 163.367
R893 B.n916 B.n17 163.367
R894 B.n916 B.n23 163.367
R895 B.n912 B.n23 163.367
R896 B.n912 B.n25 163.367
R897 B.n908 B.n25 163.367
R898 B.n908 B.n30 163.367
R899 B.n904 B.n30 163.367
R900 B.n904 B.n32 163.367
R901 B.n900 B.n32 163.367
R902 B.n900 B.n37 163.367
R903 B.n896 B.n37 163.367
R904 B.n896 B.n39 163.367
R905 B.n892 B.n39 163.367
R906 B.n892 B.n44 163.367
R907 B.n888 B.n44 163.367
R908 B.n888 B.n46 163.367
R909 B.n884 B.n46 163.367
R910 B.n884 B.n50 163.367
R911 B.n880 B.n50 163.367
R912 B.n880 B.n52 163.367
R913 B.n876 B.n52 163.367
R914 B.n876 B.n58 163.367
R915 B.n872 B.n58 163.367
R916 B.n872 B.n60 163.367
R917 B.n868 B.n60 163.367
R918 B.n868 B.n65 163.367
R919 B.n864 B.n65 163.367
R920 B.n864 B.n67 163.367
R921 B.n860 B.n67 163.367
R922 B.n860 B.n72 163.367
R923 B.n856 B.n72 163.367
R924 B.n856 B.n74 163.367
R925 B.n852 B.n74 163.367
R926 B.n852 B.n79 163.367
R927 B.n848 B.n79 163.367
R928 B.n848 B.n81 163.367
R929 B.n844 B.n81 163.367
R930 B.n844 B.n86 163.367
R931 B.n840 B.n86 163.367
R932 B.n840 B.n88 163.367
R933 B.n836 B.n88 163.367
R934 B.n836 B.n93 163.367
R935 B.n832 B.n93 163.367
R936 B.n832 B.n95 163.367
R937 B.n828 B.n95 163.367
R938 B.n828 B.n100 163.367
R939 B.n824 B.n100 163.367
R940 B.n824 B.n102 163.367
R941 B.n820 B.n102 163.367
R942 B.n429 B.n427 163.367
R943 B.n427 B.n426 163.367
R944 B.n423 B.n422 163.367
R945 B.n420 B.n263 163.367
R946 B.n416 B.n414 163.367
R947 B.n412 B.n265 163.367
R948 B.n408 B.n406 163.367
R949 B.n404 B.n267 163.367
R950 B.n400 B.n398 163.367
R951 B.n396 B.n269 163.367
R952 B.n392 B.n390 163.367
R953 B.n388 B.n271 163.367
R954 B.n384 B.n382 163.367
R955 B.n380 B.n273 163.367
R956 B.n376 B.n374 163.367
R957 B.n371 B.n370 163.367
R958 B.n368 B.n279 163.367
R959 B.n364 B.n362 163.367
R960 B.n360 B.n281 163.367
R961 B.n356 B.n354 163.367
R962 B.n351 B.n350 163.367
R963 B.n348 B.n287 163.367
R964 B.n344 B.n342 163.367
R965 B.n340 B.n289 163.367
R966 B.n336 B.n334 163.367
R967 B.n332 B.n291 163.367
R968 B.n328 B.n326 163.367
R969 B.n324 B.n293 163.367
R970 B.n320 B.n318 163.367
R971 B.n316 B.n295 163.367
R972 B.n312 B.n310 163.367
R973 B.n308 B.n297 163.367
R974 B.n304 B.n302 163.367
R975 B.n300 B.n257 163.367
R976 B.n435 B.n255 163.367
R977 B.n439 B.n255 163.367
R978 B.n439 B.n249 163.367
R979 B.n447 B.n249 163.367
R980 B.n447 B.n247 163.367
R981 B.n451 B.n247 163.367
R982 B.n451 B.n241 163.367
R983 B.n459 B.n241 163.367
R984 B.n459 B.n239 163.367
R985 B.n463 B.n239 163.367
R986 B.n463 B.n233 163.367
R987 B.n471 B.n233 163.367
R988 B.n471 B.n231 163.367
R989 B.n475 B.n231 163.367
R990 B.n475 B.n225 163.367
R991 B.n483 B.n225 163.367
R992 B.n483 B.n223 163.367
R993 B.n487 B.n223 163.367
R994 B.n487 B.n216 163.367
R995 B.n495 B.n216 163.367
R996 B.n495 B.n214 163.367
R997 B.n499 B.n214 163.367
R998 B.n499 B.n209 163.367
R999 B.n507 B.n209 163.367
R1000 B.n507 B.n207 163.367
R1001 B.n511 B.n207 163.367
R1002 B.n511 B.n201 163.367
R1003 B.n519 B.n201 163.367
R1004 B.n519 B.n199 163.367
R1005 B.n523 B.n199 163.367
R1006 B.n523 B.n194 163.367
R1007 B.n532 B.n194 163.367
R1008 B.n532 B.n192 163.367
R1009 B.n536 B.n192 163.367
R1010 B.n536 B.n186 163.367
R1011 B.n544 B.n186 163.367
R1012 B.n544 B.n184 163.367
R1013 B.n548 B.n184 163.367
R1014 B.n548 B.n177 163.367
R1015 B.n556 B.n177 163.367
R1016 B.n556 B.n175 163.367
R1017 B.n560 B.n175 163.367
R1018 B.n560 B.n170 163.367
R1019 B.n568 B.n170 163.367
R1020 B.n568 B.n168 163.367
R1021 B.n572 B.n168 163.367
R1022 B.n572 B.n162 163.367
R1023 B.n580 B.n162 163.367
R1024 B.n580 B.n160 163.367
R1025 B.n584 B.n160 163.367
R1026 B.n584 B.n155 163.367
R1027 B.n593 B.n155 163.367
R1028 B.n593 B.n153 163.367
R1029 B.n598 B.n153 163.367
R1030 B.n598 B.n147 163.367
R1031 B.n606 B.n147 163.367
R1032 B.n607 B.n606 163.367
R1033 B.n607 B.n5 163.367
R1034 B.n6 B.n5 163.367
R1035 B.n7 B.n6 163.367
R1036 B.n612 B.n7 163.367
R1037 B.n612 B.n12 163.367
R1038 B.n13 B.n12 163.367
R1039 B.n14 B.n13 163.367
R1040 B.n617 B.n14 163.367
R1041 B.n617 B.n19 163.367
R1042 B.n20 B.n19 163.367
R1043 B.n21 B.n20 163.367
R1044 B.n622 B.n21 163.367
R1045 B.n622 B.n26 163.367
R1046 B.n27 B.n26 163.367
R1047 B.n28 B.n27 163.367
R1048 B.n627 B.n28 163.367
R1049 B.n627 B.n33 163.367
R1050 B.n34 B.n33 163.367
R1051 B.n35 B.n34 163.367
R1052 B.n632 B.n35 163.367
R1053 B.n632 B.n40 163.367
R1054 B.n41 B.n40 163.367
R1055 B.n42 B.n41 163.367
R1056 B.n637 B.n42 163.367
R1057 B.n637 B.n47 163.367
R1058 B.n48 B.n47 163.367
R1059 B.n49 B.n48 163.367
R1060 B.n642 B.n49 163.367
R1061 B.n642 B.n54 163.367
R1062 B.n55 B.n54 163.367
R1063 B.n56 B.n55 163.367
R1064 B.n647 B.n56 163.367
R1065 B.n647 B.n61 163.367
R1066 B.n62 B.n61 163.367
R1067 B.n63 B.n62 163.367
R1068 B.n652 B.n63 163.367
R1069 B.n652 B.n68 163.367
R1070 B.n69 B.n68 163.367
R1071 B.n70 B.n69 163.367
R1072 B.n657 B.n70 163.367
R1073 B.n657 B.n75 163.367
R1074 B.n76 B.n75 163.367
R1075 B.n77 B.n76 163.367
R1076 B.n662 B.n77 163.367
R1077 B.n662 B.n82 163.367
R1078 B.n83 B.n82 163.367
R1079 B.n84 B.n83 163.367
R1080 B.n667 B.n84 163.367
R1081 B.n667 B.n89 163.367
R1082 B.n90 B.n89 163.367
R1083 B.n91 B.n90 163.367
R1084 B.n672 B.n91 163.367
R1085 B.n672 B.n96 163.367
R1086 B.n97 B.n96 163.367
R1087 B.n98 B.n97 163.367
R1088 B.n677 B.n98 163.367
R1089 B.n677 B.n103 163.367
R1090 B.n104 B.n103 163.367
R1091 B.n105 B.n104 163.367
R1092 B.n816 B.n814 163.367
R1093 B.n812 B.n109 163.367
R1094 B.n808 B.n806 163.367
R1095 B.n804 B.n111 163.367
R1096 B.n800 B.n798 163.367
R1097 B.n796 B.n113 163.367
R1098 B.n792 B.n790 163.367
R1099 B.n788 B.n115 163.367
R1100 B.n784 B.n782 163.367
R1101 B.n780 B.n117 163.367
R1102 B.n776 B.n774 163.367
R1103 B.n772 B.n119 163.367
R1104 B.n768 B.n766 163.367
R1105 B.n764 B.n121 163.367
R1106 B.n759 B.n757 163.367
R1107 B.n755 B.n125 163.367
R1108 B.n751 B.n749 163.367
R1109 B.n747 B.n127 163.367
R1110 B.n743 B.n741 163.367
R1111 B.n739 B.n129 163.367
R1112 B.n735 B.n733 163.367
R1113 B.n731 B.n134 163.367
R1114 B.n727 B.n725 163.367
R1115 B.n723 B.n136 163.367
R1116 B.n719 B.n717 163.367
R1117 B.n715 B.n138 163.367
R1118 B.n711 B.n709 163.367
R1119 B.n707 B.n140 163.367
R1120 B.n703 B.n701 163.367
R1121 B.n699 B.n142 163.367
R1122 B.n695 B.n693 163.367
R1123 B.n691 B.n144 163.367
R1124 B.n687 B.n685 163.367
R1125 B.n282 B.t11 140.631
R1126 B.n130 B.t17 140.631
R1127 B.n274 B.t21 140.623
R1128 B.n122 B.t14 140.623
R1129 B.n434 B.n258 110.379
R1130 B.n821 B.n106 110.379
R1131 B.n283 B.t10 74.6919
R1132 B.n131 B.t18 74.6919
R1133 B.n275 B.t20 74.6832
R1134 B.n123 B.t15 74.6832
R1135 B.n428 B.n259 71.676
R1136 B.n426 B.n261 71.676
R1137 B.n422 B.n421 71.676
R1138 B.n415 B.n263 71.676
R1139 B.n414 B.n413 71.676
R1140 B.n407 B.n265 71.676
R1141 B.n406 B.n405 71.676
R1142 B.n399 B.n267 71.676
R1143 B.n398 B.n397 71.676
R1144 B.n391 B.n269 71.676
R1145 B.n390 B.n389 71.676
R1146 B.n383 B.n271 71.676
R1147 B.n382 B.n381 71.676
R1148 B.n375 B.n273 71.676
R1149 B.n374 B.n277 71.676
R1150 B.n370 B.n369 71.676
R1151 B.n363 B.n279 71.676
R1152 B.n362 B.n361 71.676
R1153 B.n355 B.n281 71.676
R1154 B.n354 B.n285 71.676
R1155 B.n350 B.n349 71.676
R1156 B.n343 B.n287 71.676
R1157 B.n342 B.n341 71.676
R1158 B.n335 B.n289 71.676
R1159 B.n334 B.n333 71.676
R1160 B.n327 B.n291 71.676
R1161 B.n326 B.n325 71.676
R1162 B.n319 B.n293 71.676
R1163 B.n318 B.n317 71.676
R1164 B.n311 B.n295 71.676
R1165 B.n310 B.n309 71.676
R1166 B.n303 B.n297 71.676
R1167 B.n302 B.n301 71.676
R1168 B.n815 B.n107 71.676
R1169 B.n814 B.n813 71.676
R1170 B.n807 B.n109 71.676
R1171 B.n806 B.n805 71.676
R1172 B.n799 B.n111 71.676
R1173 B.n798 B.n797 71.676
R1174 B.n791 B.n113 71.676
R1175 B.n790 B.n789 71.676
R1176 B.n783 B.n115 71.676
R1177 B.n782 B.n781 71.676
R1178 B.n775 B.n117 71.676
R1179 B.n774 B.n773 71.676
R1180 B.n767 B.n119 71.676
R1181 B.n766 B.n765 71.676
R1182 B.n758 B.n121 71.676
R1183 B.n757 B.n756 71.676
R1184 B.n750 B.n125 71.676
R1185 B.n749 B.n748 71.676
R1186 B.n742 B.n127 71.676
R1187 B.n741 B.n740 71.676
R1188 B.n734 B.n129 71.676
R1189 B.n733 B.n732 71.676
R1190 B.n726 B.n134 71.676
R1191 B.n725 B.n724 71.676
R1192 B.n718 B.n136 71.676
R1193 B.n717 B.n716 71.676
R1194 B.n710 B.n138 71.676
R1195 B.n709 B.n708 71.676
R1196 B.n702 B.n140 71.676
R1197 B.n701 B.n700 71.676
R1198 B.n694 B.n142 71.676
R1199 B.n693 B.n692 71.676
R1200 B.n686 B.n144 71.676
R1201 B.n685 B.n684 71.676
R1202 B.n684 B.n683 71.676
R1203 B.n687 B.n686 71.676
R1204 B.n692 B.n691 71.676
R1205 B.n695 B.n694 71.676
R1206 B.n700 B.n699 71.676
R1207 B.n703 B.n702 71.676
R1208 B.n708 B.n707 71.676
R1209 B.n711 B.n710 71.676
R1210 B.n716 B.n715 71.676
R1211 B.n719 B.n718 71.676
R1212 B.n724 B.n723 71.676
R1213 B.n727 B.n726 71.676
R1214 B.n732 B.n731 71.676
R1215 B.n735 B.n734 71.676
R1216 B.n740 B.n739 71.676
R1217 B.n743 B.n742 71.676
R1218 B.n748 B.n747 71.676
R1219 B.n751 B.n750 71.676
R1220 B.n756 B.n755 71.676
R1221 B.n759 B.n758 71.676
R1222 B.n765 B.n764 71.676
R1223 B.n768 B.n767 71.676
R1224 B.n773 B.n772 71.676
R1225 B.n776 B.n775 71.676
R1226 B.n781 B.n780 71.676
R1227 B.n784 B.n783 71.676
R1228 B.n789 B.n788 71.676
R1229 B.n792 B.n791 71.676
R1230 B.n797 B.n796 71.676
R1231 B.n800 B.n799 71.676
R1232 B.n805 B.n804 71.676
R1233 B.n808 B.n807 71.676
R1234 B.n813 B.n812 71.676
R1235 B.n816 B.n815 71.676
R1236 B.n429 B.n428 71.676
R1237 B.n423 B.n261 71.676
R1238 B.n421 B.n420 71.676
R1239 B.n416 B.n415 71.676
R1240 B.n413 B.n412 71.676
R1241 B.n408 B.n407 71.676
R1242 B.n405 B.n404 71.676
R1243 B.n400 B.n399 71.676
R1244 B.n397 B.n396 71.676
R1245 B.n392 B.n391 71.676
R1246 B.n389 B.n388 71.676
R1247 B.n384 B.n383 71.676
R1248 B.n381 B.n380 71.676
R1249 B.n376 B.n375 71.676
R1250 B.n371 B.n277 71.676
R1251 B.n369 B.n368 71.676
R1252 B.n364 B.n363 71.676
R1253 B.n361 B.n360 71.676
R1254 B.n356 B.n355 71.676
R1255 B.n351 B.n285 71.676
R1256 B.n349 B.n348 71.676
R1257 B.n344 B.n343 71.676
R1258 B.n341 B.n340 71.676
R1259 B.n336 B.n335 71.676
R1260 B.n333 B.n332 71.676
R1261 B.n328 B.n327 71.676
R1262 B.n325 B.n324 71.676
R1263 B.n320 B.n319 71.676
R1264 B.n317 B.n316 71.676
R1265 B.n312 B.n311 71.676
R1266 B.n309 B.n308 71.676
R1267 B.n304 B.n303 71.676
R1268 B.n301 B.n300 71.676
R1269 B.n283 B.n282 65.9399
R1270 B.n275 B.n274 65.9399
R1271 B.n123 B.n122 65.9399
R1272 B.n131 B.n130 65.9399
R1273 B.n284 B.n283 59.5399
R1274 B.n276 B.n275 59.5399
R1275 B.n761 B.n123 59.5399
R1276 B.n132 B.n131 59.5399
R1277 B.n434 B.n254 57.2966
R1278 B.n440 B.n254 57.2966
R1279 B.n440 B.n250 57.2966
R1280 B.n446 B.n250 57.2966
R1281 B.n446 B.n246 57.2966
R1282 B.n452 B.n246 57.2966
R1283 B.n452 B.n242 57.2966
R1284 B.n458 B.n242 57.2966
R1285 B.n464 B.n238 57.2966
R1286 B.n464 B.n234 57.2966
R1287 B.n470 B.n234 57.2966
R1288 B.n470 B.n230 57.2966
R1289 B.n476 B.n230 57.2966
R1290 B.n476 B.n226 57.2966
R1291 B.n482 B.n226 57.2966
R1292 B.n482 B.n222 57.2966
R1293 B.n488 B.n222 57.2966
R1294 B.n488 B.n217 57.2966
R1295 B.n494 B.n217 57.2966
R1296 B.n494 B.n218 57.2966
R1297 B.n500 B.n210 57.2966
R1298 B.n506 B.n210 57.2966
R1299 B.n506 B.n206 57.2966
R1300 B.n512 B.n206 57.2966
R1301 B.n512 B.n202 57.2966
R1302 B.n518 B.n202 57.2966
R1303 B.n518 B.n198 57.2966
R1304 B.n525 B.n198 57.2966
R1305 B.n525 B.n524 57.2966
R1306 B.n531 B.n191 57.2966
R1307 B.n537 B.n191 57.2966
R1308 B.n537 B.n187 57.2966
R1309 B.n543 B.n187 57.2966
R1310 B.n543 B.n183 57.2966
R1311 B.n549 B.n183 57.2966
R1312 B.n549 B.n178 57.2966
R1313 B.n555 B.n178 57.2966
R1314 B.n555 B.n179 57.2966
R1315 B.n561 B.n171 57.2966
R1316 B.n567 B.n171 57.2966
R1317 B.n567 B.n167 57.2966
R1318 B.n573 B.n167 57.2966
R1319 B.n573 B.n163 57.2966
R1320 B.n579 B.n163 57.2966
R1321 B.n579 B.n159 57.2966
R1322 B.n586 B.n159 57.2966
R1323 B.n586 B.n585 57.2966
R1324 B.n592 B.n152 57.2966
R1325 B.n599 B.n152 57.2966
R1326 B.n599 B.n148 57.2966
R1327 B.n605 B.n148 57.2966
R1328 B.n605 B.n4 57.2966
R1329 B.n935 B.n4 57.2966
R1330 B.n935 B.n934 57.2966
R1331 B.n934 B.n933 57.2966
R1332 B.n933 B.n8 57.2966
R1333 B.n927 B.n8 57.2966
R1334 B.n927 B.n926 57.2966
R1335 B.n926 B.n925 57.2966
R1336 B.n919 B.n18 57.2966
R1337 B.n919 B.n918 57.2966
R1338 B.n918 B.n917 57.2966
R1339 B.n917 B.n22 57.2966
R1340 B.n911 B.n22 57.2966
R1341 B.n911 B.n910 57.2966
R1342 B.n910 B.n909 57.2966
R1343 B.n909 B.n29 57.2966
R1344 B.n903 B.n29 57.2966
R1345 B.n902 B.n901 57.2966
R1346 B.n901 B.n36 57.2966
R1347 B.n895 B.n36 57.2966
R1348 B.n895 B.n894 57.2966
R1349 B.n894 B.n893 57.2966
R1350 B.n893 B.n43 57.2966
R1351 B.n887 B.n43 57.2966
R1352 B.n887 B.n886 57.2966
R1353 B.n886 B.n885 57.2966
R1354 B.n879 B.n53 57.2966
R1355 B.n879 B.n878 57.2966
R1356 B.n878 B.n877 57.2966
R1357 B.n877 B.n57 57.2966
R1358 B.n871 B.n57 57.2966
R1359 B.n871 B.n870 57.2966
R1360 B.n870 B.n869 57.2966
R1361 B.n869 B.n64 57.2966
R1362 B.n863 B.n64 57.2966
R1363 B.n862 B.n861 57.2966
R1364 B.n861 B.n71 57.2966
R1365 B.n855 B.n71 57.2966
R1366 B.n855 B.n854 57.2966
R1367 B.n854 B.n853 57.2966
R1368 B.n853 B.n78 57.2966
R1369 B.n847 B.n78 57.2966
R1370 B.n847 B.n846 57.2966
R1371 B.n846 B.n845 57.2966
R1372 B.n845 B.n85 57.2966
R1373 B.n839 B.n85 57.2966
R1374 B.n839 B.n838 57.2966
R1375 B.n837 B.n92 57.2966
R1376 B.n831 B.n92 57.2966
R1377 B.n831 B.n830 57.2966
R1378 B.n830 B.n829 57.2966
R1379 B.n829 B.n99 57.2966
R1380 B.n823 B.n99 57.2966
R1381 B.n823 B.n822 57.2966
R1382 B.n822 B.n821 57.2966
R1383 B.t9 B.n238 46.3429
R1384 B.n838 B.t13 46.3429
R1385 B.n500 B.t1 34.5467
R1386 B.n531 B.t4 34.5467
R1387 B.n561 B.t7 34.5467
R1388 B.n592 B.t6 34.5467
R1389 B.n925 B.t5 34.5467
R1390 B.n903 B.t3 34.5467
R1391 B.n885 B.t2 34.5467
R1392 B.n863 B.t0 34.5467
R1393 B.n819 B.n818 33.5615
R1394 B.n682 B.n681 33.5615
R1395 B.n436 B.n256 33.5615
R1396 B.n432 B.n431 33.5615
R1397 B.n218 B.t1 22.7504
R1398 B.n524 B.t4 22.7504
R1399 B.n179 B.t7 22.7504
R1400 B.n585 B.t6 22.7504
R1401 B.n18 B.t5 22.7504
R1402 B.t3 B.n902 22.7504
R1403 B.n53 B.t2 22.7504
R1404 B.t0 B.n862 22.7504
R1405 B B.n937 18.0485
R1406 B.n458 B.t9 10.9542
R1407 B.t13 B.n837 10.9542
R1408 B.n818 B.n817 10.6151
R1409 B.n817 B.n108 10.6151
R1410 B.n811 B.n108 10.6151
R1411 B.n811 B.n810 10.6151
R1412 B.n810 B.n809 10.6151
R1413 B.n809 B.n110 10.6151
R1414 B.n803 B.n110 10.6151
R1415 B.n803 B.n802 10.6151
R1416 B.n802 B.n801 10.6151
R1417 B.n801 B.n112 10.6151
R1418 B.n795 B.n112 10.6151
R1419 B.n795 B.n794 10.6151
R1420 B.n794 B.n793 10.6151
R1421 B.n793 B.n114 10.6151
R1422 B.n787 B.n114 10.6151
R1423 B.n787 B.n786 10.6151
R1424 B.n786 B.n785 10.6151
R1425 B.n785 B.n116 10.6151
R1426 B.n779 B.n116 10.6151
R1427 B.n779 B.n778 10.6151
R1428 B.n778 B.n777 10.6151
R1429 B.n777 B.n118 10.6151
R1430 B.n771 B.n118 10.6151
R1431 B.n771 B.n770 10.6151
R1432 B.n770 B.n769 10.6151
R1433 B.n769 B.n120 10.6151
R1434 B.n763 B.n120 10.6151
R1435 B.n763 B.n762 10.6151
R1436 B.n760 B.n124 10.6151
R1437 B.n754 B.n124 10.6151
R1438 B.n754 B.n753 10.6151
R1439 B.n753 B.n752 10.6151
R1440 B.n752 B.n126 10.6151
R1441 B.n746 B.n126 10.6151
R1442 B.n746 B.n745 10.6151
R1443 B.n745 B.n744 10.6151
R1444 B.n744 B.n128 10.6151
R1445 B.n738 B.n737 10.6151
R1446 B.n737 B.n736 10.6151
R1447 B.n736 B.n133 10.6151
R1448 B.n730 B.n133 10.6151
R1449 B.n730 B.n729 10.6151
R1450 B.n729 B.n728 10.6151
R1451 B.n728 B.n135 10.6151
R1452 B.n722 B.n135 10.6151
R1453 B.n722 B.n721 10.6151
R1454 B.n721 B.n720 10.6151
R1455 B.n720 B.n137 10.6151
R1456 B.n714 B.n137 10.6151
R1457 B.n714 B.n713 10.6151
R1458 B.n713 B.n712 10.6151
R1459 B.n712 B.n139 10.6151
R1460 B.n706 B.n139 10.6151
R1461 B.n706 B.n705 10.6151
R1462 B.n705 B.n704 10.6151
R1463 B.n704 B.n141 10.6151
R1464 B.n698 B.n141 10.6151
R1465 B.n698 B.n697 10.6151
R1466 B.n697 B.n696 10.6151
R1467 B.n696 B.n143 10.6151
R1468 B.n690 B.n143 10.6151
R1469 B.n690 B.n689 10.6151
R1470 B.n689 B.n688 10.6151
R1471 B.n688 B.n145 10.6151
R1472 B.n682 B.n145 10.6151
R1473 B.n437 B.n436 10.6151
R1474 B.n438 B.n437 10.6151
R1475 B.n438 B.n248 10.6151
R1476 B.n448 B.n248 10.6151
R1477 B.n449 B.n448 10.6151
R1478 B.n450 B.n449 10.6151
R1479 B.n450 B.n240 10.6151
R1480 B.n460 B.n240 10.6151
R1481 B.n461 B.n460 10.6151
R1482 B.n462 B.n461 10.6151
R1483 B.n462 B.n232 10.6151
R1484 B.n472 B.n232 10.6151
R1485 B.n473 B.n472 10.6151
R1486 B.n474 B.n473 10.6151
R1487 B.n474 B.n224 10.6151
R1488 B.n484 B.n224 10.6151
R1489 B.n485 B.n484 10.6151
R1490 B.n486 B.n485 10.6151
R1491 B.n486 B.n215 10.6151
R1492 B.n496 B.n215 10.6151
R1493 B.n497 B.n496 10.6151
R1494 B.n498 B.n497 10.6151
R1495 B.n498 B.n208 10.6151
R1496 B.n508 B.n208 10.6151
R1497 B.n509 B.n508 10.6151
R1498 B.n510 B.n509 10.6151
R1499 B.n510 B.n200 10.6151
R1500 B.n520 B.n200 10.6151
R1501 B.n521 B.n520 10.6151
R1502 B.n522 B.n521 10.6151
R1503 B.n522 B.n193 10.6151
R1504 B.n533 B.n193 10.6151
R1505 B.n534 B.n533 10.6151
R1506 B.n535 B.n534 10.6151
R1507 B.n535 B.n185 10.6151
R1508 B.n545 B.n185 10.6151
R1509 B.n546 B.n545 10.6151
R1510 B.n547 B.n546 10.6151
R1511 B.n547 B.n176 10.6151
R1512 B.n557 B.n176 10.6151
R1513 B.n558 B.n557 10.6151
R1514 B.n559 B.n558 10.6151
R1515 B.n559 B.n169 10.6151
R1516 B.n569 B.n169 10.6151
R1517 B.n570 B.n569 10.6151
R1518 B.n571 B.n570 10.6151
R1519 B.n571 B.n161 10.6151
R1520 B.n581 B.n161 10.6151
R1521 B.n582 B.n581 10.6151
R1522 B.n583 B.n582 10.6151
R1523 B.n583 B.n154 10.6151
R1524 B.n594 B.n154 10.6151
R1525 B.n595 B.n594 10.6151
R1526 B.n597 B.n595 10.6151
R1527 B.n597 B.n596 10.6151
R1528 B.n596 B.n146 10.6151
R1529 B.n608 B.n146 10.6151
R1530 B.n609 B.n608 10.6151
R1531 B.n610 B.n609 10.6151
R1532 B.n611 B.n610 10.6151
R1533 B.n613 B.n611 10.6151
R1534 B.n614 B.n613 10.6151
R1535 B.n615 B.n614 10.6151
R1536 B.n616 B.n615 10.6151
R1537 B.n618 B.n616 10.6151
R1538 B.n619 B.n618 10.6151
R1539 B.n620 B.n619 10.6151
R1540 B.n621 B.n620 10.6151
R1541 B.n623 B.n621 10.6151
R1542 B.n624 B.n623 10.6151
R1543 B.n625 B.n624 10.6151
R1544 B.n626 B.n625 10.6151
R1545 B.n628 B.n626 10.6151
R1546 B.n629 B.n628 10.6151
R1547 B.n630 B.n629 10.6151
R1548 B.n631 B.n630 10.6151
R1549 B.n633 B.n631 10.6151
R1550 B.n634 B.n633 10.6151
R1551 B.n635 B.n634 10.6151
R1552 B.n636 B.n635 10.6151
R1553 B.n638 B.n636 10.6151
R1554 B.n639 B.n638 10.6151
R1555 B.n640 B.n639 10.6151
R1556 B.n641 B.n640 10.6151
R1557 B.n643 B.n641 10.6151
R1558 B.n644 B.n643 10.6151
R1559 B.n645 B.n644 10.6151
R1560 B.n646 B.n645 10.6151
R1561 B.n648 B.n646 10.6151
R1562 B.n649 B.n648 10.6151
R1563 B.n650 B.n649 10.6151
R1564 B.n651 B.n650 10.6151
R1565 B.n653 B.n651 10.6151
R1566 B.n654 B.n653 10.6151
R1567 B.n655 B.n654 10.6151
R1568 B.n656 B.n655 10.6151
R1569 B.n658 B.n656 10.6151
R1570 B.n659 B.n658 10.6151
R1571 B.n660 B.n659 10.6151
R1572 B.n661 B.n660 10.6151
R1573 B.n663 B.n661 10.6151
R1574 B.n664 B.n663 10.6151
R1575 B.n665 B.n664 10.6151
R1576 B.n666 B.n665 10.6151
R1577 B.n668 B.n666 10.6151
R1578 B.n669 B.n668 10.6151
R1579 B.n670 B.n669 10.6151
R1580 B.n671 B.n670 10.6151
R1581 B.n673 B.n671 10.6151
R1582 B.n674 B.n673 10.6151
R1583 B.n675 B.n674 10.6151
R1584 B.n676 B.n675 10.6151
R1585 B.n678 B.n676 10.6151
R1586 B.n679 B.n678 10.6151
R1587 B.n680 B.n679 10.6151
R1588 B.n681 B.n680 10.6151
R1589 B.n431 B.n430 10.6151
R1590 B.n430 B.n260 10.6151
R1591 B.n425 B.n260 10.6151
R1592 B.n425 B.n424 10.6151
R1593 B.n424 B.n262 10.6151
R1594 B.n419 B.n262 10.6151
R1595 B.n419 B.n418 10.6151
R1596 B.n418 B.n417 10.6151
R1597 B.n417 B.n264 10.6151
R1598 B.n411 B.n264 10.6151
R1599 B.n411 B.n410 10.6151
R1600 B.n410 B.n409 10.6151
R1601 B.n409 B.n266 10.6151
R1602 B.n403 B.n266 10.6151
R1603 B.n403 B.n402 10.6151
R1604 B.n402 B.n401 10.6151
R1605 B.n401 B.n268 10.6151
R1606 B.n395 B.n268 10.6151
R1607 B.n395 B.n394 10.6151
R1608 B.n394 B.n393 10.6151
R1609 B.n393 B.n270 10.6151
R1610 B.n387 B.n270 10.6151
R1611 B.n387 B.n386 10.6151
R1612 B.n386 B.n385 10.6151
R1613 B.n385 B.n272 10.6151
R1614 B.n379 B.n272 10.6151
R1615 B.n379 B.n378 10.6151
R1616 B.n378 B.n377 10.6151
R1617 B.n373 B.n372 10.6151
R1618 B.n372 B.n278 10.6151
R1619 B.n367 B.n278 10.6151
R1620 B.n367 B.n366 10.6151
R1621 B.n366 B.n365 10.6151
R1622 B.n365 B.n280 10.6151
R1623 B.n359 B.n280 10.6151
R1624 B.n359 B.n358 10.6151
R1625 B.n358 B.n357 10.6151
R1626 B.n353 B.n352 10.6151
R1627 B.n352 B.n286 10.6151
R1628 B.n347 B.n286 10.6151
R1629 B.n347 B.n346 10.6151
R1630 B.n346 B.n345 10.6151
R1631 B.n345 B.n288 10.6151
R1632 B.n339 B.n288 10.6151
R1633 B.n339 B.n338 10.6151
R1634 B.n338 B.n337 10.6151
R1635 B.n337 B.n290 10.6151
R1636 B.n331 B.n290 10.6151
R1637 B.n331 B.n330 10.6151
R1638 B.n330 B.n329 10.6151
R1639 B.n329 B.n292 10.6151
R1640 B.n323 B.n292 10.6151
R1641 B.n323 B.n322 10.6151
R1642 B.n322 B.n321 10.6151
R1643 B.n321 B.n294 10.6151
R1644 B.n315 B.n294 10.6151
R1645 B.n315 B.n314 10.6151
R1646 B.n314 B.n313 10.6151
R1647 B.n313 B.n296 10.6151
R1648 B.n307 B.n296 10.6151
R1649 B.n307 B.n306 10.6151
R1650 B.n306 B.n305 10.6151
R1651 B.n305 B.n298 10.6151
R1652 B.n299 B.n298 10.6151
R1653 B.n299 B.n256 10.6151
R1654 B.n432 B.n252 10.6151
R1655 B.n442 B.n252 10.6151
R1656 B.n443 B.n442 10.6151
R1657 B.n444 B.n443 10.6151
R1658 B.n444 B.n244 10.6151
R1659 B.n454 B.n244 10.6151
R1660 B.n455 B.n454 10.6151
R1661 B.n456 B.n455 10.6151
R1662 B.n456 B.n236 10.6151
R1663 B.n466 B.n236 10.6151
R1664 B.n467 B.n466 10.6151
R1665 B.n468 B.n467 10.6151
R1666 B.n468 B.n228 10.6151
R1667 B.n478 B.n228 10.6151
R1668 B.n479 B.n478 10.6151
R1669 B.n480 B.n479 10.6151
R1670 B.n480 B.n220 10.6151
R1671 B.n490 B.n220 10.6151
R1672 B.n491 B.n490 10.6151
R1673 B.n492 B.n491 10.6151
R1674 B.n492 B.n212 10.6151
R1675 B.n502 B.n212 10.6151
R1676 B.n503 B.n502 10.6151
R1677 B.n504 B.n503 10.6151
R1678 B.n504 B.n204 10.6151
R1679 B.n514 B.n204 10.6151
R1680 B.n515 B.n514 10.6151
R1681 B.n516 B.n515 10.6151
R1682 B.n516 B.n196 10.6151
R1683 B.n527 B.n196 10.6151
R1684 B.n528 B.n527 10.6151
R1685 B.n529 B.n528 10.6151
R1686 B.n529 B.n189 10.6151
R1687 B.n539 B.n189 10.6151
R1688 B.n540 B.n539 10.6151
R1689 B.n541 B.n540 10.6151
R1690 B.n541 B.n181 10.6151
R1691 B.n551 B.n181 10.6151
R1692 B.n552 B.n551 10.6151
R1693 B.n553 B.n552 10.6151
R1694 B.n553 B.n173 10.6151
R1695 B.n563 B.n173 10.6151
R1696 B.n564 B.n563 10.6151
R1697 B.n565 B.n564 10.6151
R1698 B.n565 B.n165 10.6151
R1699 B.n575 B.n165 10.6151
R1700 B.n576 B.n575 10.6151
R1701 B.n577 B.n576 10.6151
R1702 B.n577 B.n157 10.6151
R1703 B.n588 B.n157 10.6151
R1704 B.n589 B.n588 10.6151
R1705 B.n590 B.n589 10.6151
R1706 B.n590 B.n150 10.6151
R1707 B.n601 B.n150 10.6151
R1708 B.n602 B.n601 10.6151
R1709 B.n603 B.n602 10.6151
R1710 B.n603 B.n0 10.6151
R1711 B.n931 B.n1 10.6151
R1712 B.n931 B.n930 10.6151
R1713 B.n930 B.n929 10.6151
R1714 B.n929 B.n10 10.6151
R1715 B.n923 B.n10 10.6151
R1716 B.n923 B.n922 10.6151
R1717 B.n922 B.n921 10.6151
R1718 B.n921 B.n16 10.6151
R1719 B.n915 B.n16 10.6151
R1720 B.n915 B.n914 10.6151
R1721 B.n914 B.n913 10.6151
R1722 B.n913 B.n24 10.6151
R1723 B.n907 B.n24 10.6151
R1724 B.n907 B.n906 10.6151
R1725 B.n906 B.n905 10.6151
R1726 B.n905 B.n31 10.6151
R1727 B.n899 B.n31 10.6151
R1728 B.n899 B.n898 10.6151
R1729 B.n898 B.n897 10.6151
R1730 B.n897 B.n38 10.6151
R1731 B.n891 B.n38 10.6151
R1732 B.n891 B.n890 10.6151
R1733 B.n890 B.n889 10.6151
R1734 B.n889 B.n45 10.6151
R1735 B.n883 B.n45 10.6151
R1736 B.n883 B.n882 10.6151
R1737 B.n882 B.n881 10.6151
R1738 B.n881 B.n51 10.6151
R1739 B.n875 B.n51 10.6151
R1740 B.n875 B.n874 10.6151
R1741 B.n874 B.n873 10.6151
R1742 B.n873 B.n59 10.6151
R1743 B.n867 B.n59 10.6151
R1744 B.n867 B.n866 10.6151
R1745 B.n866 B.n865 10.6151
R1746 B.n865 B.n66 10.6151
R1747 B.n859 B.n66 10.6151
R1748 B.n859 B.n858 10.6151
R1749 B.n858 B.n857 10.6151
R1750 B.n857 B.n73 10.6151
R1751 B.n851 B.n73 10.6151
R1752 B.n851 B.n850 10.6151
R1753 B.n850 B.n849 10.6151
R1754 B.n849 B.n80 10.6151
R1755 B.n843 B.n80 10.6151
R1756 B.n843 B.n842 10.6151
R1757 B.n842 B.n841 10.6151
R1758 B.n841 B.n87 10.6151
R1759 B.n835 B.n87 10.6151
R1760 B.n835 B.n834 10.6151
R1761 B.n834 B.n833 10.6151
R1762 B.n833 B.n94 10.6151
R1763 B.n827 B.n94 10.6151
R1764 B.n827 B.n826 10.6151
R1765 B.n826 B.n825 10.6151
R1766 B.n825 B.n101 10.6151
R1767 B.n819 B.n101 10.6151
R1768 B.n762 B.n761 9.52245
R1769 B.n738 B.n132 9.52245
R1770 B.n377 B.n276 9.52245
R1771 B.n353 B.n284 9.52245
R1772 B.n937 B.n0 2.81026
R1773 B.n937 B.n1 2.81026
R1774 B.n761 B.n760 1.09318
R1775 B.n132 B.n128 1.09318
R1776 B.n373 B.n276 1.09318
R1777 B.n357 B.n284 1.09318
R1778 VP.n21 VP.n18 161.3
R1779 VP.n23 VP.n22 161.3
R1780 VP.n24 VP.n17 161.3
R1781 VP.n26 VP.n25 161.3
R1782 VP.n27 VP.n16 161.3
R1783 VP.n29 VP.n28 161.3
R1784 VP.n31 VP.n30 161.3
R1785 VP.n32 VP.n14 161.3
R1786 VP.n34 VP.n33 161.3
R1787 VP.n35 VP.n13 161.3
R1788 VP.n37 VP.n36 161.3
R1789 VP.n38 VP.n12 161.3
R1790 VP.n40 VP.n39 161.3
R1791 VP.n75 VP.n74 161.3
R1792 VP.n73 VP.n1 161.3
R1793 VP.n72 VP.n71 161.3
R1794 VP.n70 VP.n2 161.3
R1795 VP.n69 VP.n68 161.3
R1796 VP.n67 VP.n3 161.3
R1797 VP.n66 VP.n65 161.3
R1798 VP.n64 VP.n63 161.3
R1799 VP.n62 VP.n5 161.3
R1800 VP.n61 VP.n60 161.3
R1801 VP.n59 VP.n6 161.3
R1802 VP.n58 VP.n57 161.3
R1803 VP.n56 VP.n7 161.3
R1804 VP.n54 VP.n53 161.3
R1805 VP.n52 VP.n8 161.3
R1806 VP.n51 VP.n50 161.3
R1807 VP.n49 VP.n9 161.3
R1808 VP.n48 VP.n47 161.3
R1809 VP.n46 VP.n10 161.3
R1810 VP.n45 VP.n44 161.3
R1811 VP.n19 VP.t3 94.2633
R1812 VP.n43 VP.n42 72.8506
R1813 VP.n76 VP.n0 72.8506
R1814 VP.n41 VP.n11 72.8506
R1815 VP.n43 VP.t1 61.0748
R1816 VP.n55 VP.t5 61.0748
R1817 VP.n4 VP.t0 61.0748
R1818 VP.n0 VP.t2 61.0748
R1819 VP.n11 VP.t7 61.0748
R1820 VP.n15 VP.t6 61.0748
R1821 VP.n20 VP.t4 61.0748
R1822 VP.n61 VP.n6 56.4773
R1823 VP.n26 VP.n17 56.4773
R1824 VP.n49 VP.n48 55.0167
R1825 VP.n72 VP.n2 55.0167
R1826 VP.n37 VP.n13 55.0167
R1827 VP.n20 VP.n19 51.6654
R1828 VP.n42 VP.n41 49.9915
R1829 VP.n50 VP.n49 25.8045
R1830 VP.n68 VP.n2 25.8045
R1831 VP.n33 VP.n13 25.8045
R1832 VP.n44 VP.n10 24.3439
R1833 VP.n48 VP.n10 24.3439
R1834 VP.n50 VP.n8 24.3439
R1835 VP.n54 VP.n8 24.3439
R1836 VP.n57 VP.n56 24.3439
R1837 VP.n57 VP.n6 24.3439
R1838 VP.n62 VP.n61 24.3439
R1839 VP.n63 VP.n62 24.3439
R1840 VP.n67 VP.n66 24.3439
R1841 VP.n68 VP.n67 24.3439
R1842 VP.n73 VP.n72 24.3439
R1843 VP.n74 VP.n73 24.3439
R1844 VP.n38 VP.n37 24.3439
R1845 VP.n39 VP.n38 24.3439
R1846 VP.n27 VP.n26 24.3439
R1847 VP.n28 VP.n27 24.3439
R1848 VP.n32 VP.n31 24.3439
R1849 VP.n33 VP.n32 24.3439
R1850 VP.n22 VP.n21 24.3439
R1851 VP.n22 VP.n17 24.3439
R1852 VP.n56 VP.n55 21.9096
R1853 VP.n63 VP.n4 21.9096
R1854 VP.n28 VP.n15 21.9096
R1855 VP.n21 VP.n20 21.9096
R1856 VP.n44 VP.n43 17.0409
R1857 VP.n74 VP.n0 17.0409
R1858 VP.n39 VP.n11 17.0409
R1859 VP.n19 VP.n18 4.06491
R1860 VP.n55 VP.n54 2.43484
R1861 VP.n66 VP.n4 2.43484
R1862 VP.n31 VP.n15 2.43484
R1863 VP.n41 VP.n40 0.355081
R1864 VP.n45 VP.n42 0.355081
R1865 VP.n76 VP.n75 0.355081
R1866 VP VP.n76 0.26685
R1867 VP.n23 VP.n18 0.189894
R1868 VP.n24 VP.n23 0.189894
R1869 VP.n25 VP.n24 0.189894
R1870 VP.n25 VP.n16 0.189894
R1871 VP.n29 VP.n16 0.189894
R1872 VP.n30 VP.n29 0.189894
R1873 VP.n30 VP.n14 0.189894
R1874 VP.n34 VP.n14 0.189894
R1875 VP.n35 VP.n34 0.189894
R1876 VP.n36 VP.n35 0.189894
R1877 VP.n36 VP.n12 0.189894
R1878 VP.n40 VP.n12 0.189894
R1879 VP.n46 VP.n45 0.189894
R1880 VP.n47 VP.n46 0.189894
R1881 VP.n47 VP.n9 0.189894
R1882 VP.n51 VP.n9 0.189894
R1883 VP.n52 VP.n51 0.189894
R1884 VP.n53 VP.n52 0.189894
R1885 VP.n53 VP.n7 0.189894
R1886 VP.n58 VP.n7 0.189894
R1887 VP.n59 VP.n58 0.189894
R1888 VP.n60 VP.n59 0.189894
R1889 VP.n60 VP.n5 0.189894
R1890 VP.n64 VP.n5 0.189894
R1891 VP.n65 VP.n64 0.189894
R1892 VP.n65 VP.n3 0.189894
R1893 VP.n69 VP.n3 0.189894
R1894 VP.n70 VP.n69 0.189894
R1895 VP.n71 VP.n70 0.189894
R1896 VP.n71 VP.n1 0.189894
R1897 VP.n75 VP.n1 0.189894
R1898 VDD1 VDD1.n0 65.9684
R1899 VDD1.n3 VDD1.n2 65.8549
R1900 VDD1.n3 VDD1.n1 65.8549
R1901 VDD1.n5 VDD1.n4 64.4447
R1902 VDD1.n5 VDD1.n3 44.1949
R1903 VDD1.n4 VDD1.t1 2.54549
R1904 VDD1.n4 VDD1.t0 2.54549
R1905 VDD1.n0 VDD1.t4 2.54549
R1906 VDD1.n0 VDD1.t3 2.54549
R1907 VDD1.n2 VDD1.t7 2.54549
R1908 VDD1.n2 VDD1.t5 2.54549
R1909 VDD1.n1 VDD1.t6 2.54549
R1910 VDD1.n1 VDD1.t2 2.54549
R1911 VDD1 VDD1.n5 1.40783
C0 VDD2 VDD1 2.02259f
C1 VN VP 7.46581f
C2 VTAIL VP 6.73457f
C3 VDD1 VP 6.38414f
C4 VTAIL VN 6.72046f
C5 VDD1 VN 0.152316f
C6 VDD2 VP 0.56943f
C7 VDD1 VTAIL 6.9213f
C8 VDD2 VN 5.96867f
C9 VDD2 VTAIL 6.97887f
C10 VDD2 B 5.590075f
C11 VDD1 B 6.079427f
C12 VTAIL B 8.271098f
C13 VN B 17.041859f
C14 VP B 15.692099f
C15 VDD1.t4 B 0.174108f
C16 VDD1.t3 B 0.174108f
C17 VDD1.n0 B 1.50835f
C18 VDD1.t6 B 0.174108f
C19 VDD1.t2 B 0.174108f
C20 VDD1.n1 B 1.50703f
C21 VDD1.t7 B 0.174108f
C22 VDD1.t5 B 0.174108f
C23 VDD1.n2 B 1.50703f
C24 VDD1.n3 B 3.78808f
C25 VDD1.t1 B 0.174108f
C26 VDD1.t0 B 0.174108f
C27 VDD1.n4 B 1.49325f
C28 VDD1.n5 B 3.19765f
C29 VP.t2 B 1.39765f
C30 VP.n0 B 0.591732f
C31 VP.n1 B 0.021835f
C32 VP.n2 B 0.024981f
C33 VP.n3 B 0.021835f
C34 VP.t0 B 1.39765f
C35 VP.n4 B 0.507368f
C36 VP.n5 B 0.021835f
C37 VP.n6 B 0.032013f
C38 VP.n7 B 0.021835f
C39 VP.t5 B 1.39765f
C40 VP.n8 B 0.040898f
C41 VP.n9 B 0.021835f
C42 VP.n10 B 0.040898f
C43 VP.t7 B 1.39765f
C44 VP.n11 B 0.591732f
C45 VP.n12 B 0.021835f
C46 VP.n13 B 0.024981f
C47 VP.n14 B 0.021835f
C48 VP.t6 B 1.39765f
C49 VP.n15 B 0.507368f
C50 VP.n16 B 0.021835f
C51 VP.n17 B 0.032013f
C52 VP.n18 B 0.249681f
C53 VP.t4 B 1.39765f
C54 VP.t3 B 1.63007f
C55 VP.n19 B 0.553382f
C56 VP.n20 B 0.586826f
C57 VP.n21 B 0.038879f
C58 VP.n22 B 0.040898f
C59 VP.n23 B 0.021835f
C60 VP.n24 B 0.021835f
C61 VP.n25 B 0.021835f
C62 VP.n26 B 0.032013f
C63 VP.n27 B 0.040898f
C64 VP.n28 B 0.038879f
C65 VP.n29 B 0.021835f
C66 VP.n30 B 0.021835f
C67 VP.n31 B 0.022725f
C68 VP.n32 B 0.040898f
C69 VP.n33 B 0.041973f
C70 VP.n34 B 0.021835f
C71 VP.n35 B 0.021835f
C72 VP.n36 B 0.021835f
C73 VP.n37 B 0.037971f
C74 VP.n38 B 0.040898f
C75 VP.n39 B 0.034841f
C76 VP.n40 B 0.035246f
C77 VP.n41 B 1.23686f
C78 VP.n42 B 1.25252f
C79 VP.t1 B 1.39765f
C80 VP.n43 B 0.591732f
C81 VP.n44 B 0.034841f
C82 VP.n45 B 0.035246f
C83 VP.n46 B 0.021835f
C84 VP.n47 B 0.021835f
C85 VP.n48 B 0.037971f
C86 VP.n49 B 0.024981f
C87 VP.n50 B 0.041973f
C88 VP.n51 B 0.021835f
C89 VP.n52 B 0.021835f
C90 VP.n53 B 0.021835f
C91 VP.n54 B 0.022725f
C92 VP.n55 B 0.507368f
C93 VP.n56 B 0.038879f
C94 VP.n57 B 0.040898f
C95 VP.n58 B 0.021835f
C96 VP.n59 B 0.021835f
C97 VP.n60 B 0.021835f
C98 VP.n61 B 0.032013f
C99 VP.n62 B 0.040898f
C100 VP.n63 B 0.038879f
C101 VP.n64 B 0.021835f
C102 VP.n65 B 0.021835f
C103 VP.n66 B 0.022725f
C104 VP.n67 B 0.040898f
C105 VP.n68 B 0.041973f
C106 VP.n69 B 0.021835f
C107 VP.n70 B 0.021835f
C108 VP.n71 B 0.021835f
C109 VP.n72 B 0.037971f
C110 VP.n73 B 0.040898f
C111 VP.n74 B 0.034841f
C112 VP.n75 B 0.035246f
C113 VP.n76 B 0.048729f
C114 VTAIL.t13 B 0.135874f
C115 VTAIL.t15 B 0.135874f
C116 VTAIL.n0 B 1.10264f
C117 VTAIL.n1 B 0.429291f
C118 VTAIL.t11 B 1.40556f
C119 VTAIL.n2 B 0.52626f
C120 VTAIL.t6 B 1.40556f
C121 VTAIL.n3 B 0.52626f
C122 VTAIL.t4 B 0.135874f
C123 VTAIL.t7 B 0.135874f
C124 VTAIL.n4 B 1.10264f
C125 VTAIL.n5 B 0.633876f
C126 VTAIL.t1 B 1.40556f
C127 VTAIL.n6 B 1.47936f
C128 VTAIL.t12 B 1.40556f
C129 VTAIL.n7 B 1.47935f
C130 VTAIL.t10 B 0.135874f
C131 VTAIL.t14 B 0.135874f
C132 VTAIL.n8 B 1.10265f
C133 VTAIL.n9 B 0.633873f
C134 VTAIL.t8 B 1.40556f
C135 VTAIL.n10 B 0.526252f
C136 VTAIL.t5 B 1.40556f
C137 VTAIL.n11 B 0.526252f
C138 VTAIL.t3 B 0.135874f
C139 VTAIL.t2 B 0.135874f
C140 VTAIL.n12 B 1.10265f
C141 VTAIL.n13 B 0.633873f
C142 VTAIL.t0 B 1.40556f
C143 VTAIL.n14 B 1.47935f
C144 VTAIL.t9 B 1.40556f
C145 VTAIL.n15 B 1.47522f
C146 VDD2.t1 B 0.171869f
C147 VDD2.t3 B 0.171869f
C148 VDD2.n0 B 1.48765f
C149 VDD2.t4 B 0.171869f
C150 VDD2.t5 B 0.171869f
C151 VDD2.n1 B 1.48765f
C152 VDD2.n2 B 3.68128f
C153 VDD2.t2 B 0.171869f
C154 VDD2.t6 B 0.171869f
C155 VDD2.n3 B 1.47405f
C156 VDD2.n4 B 3.12185f
C157 VDD2.t0 B 0.171869f
C158 VDD2.t7 B 0.171869f
C159 VDD2.n5 B 1.48761f
C160 VN.t6 B 1.36847f
C161 VN.n0 B 0.579379f
C162 VN.n1 B 0.021379f
C163 VN.n2 B 0.02446f
C164 VN.n3 B 0.021379f
C165 VN.t0 B 1.36847f
C166 VN.n4 B 0.496776f
C167 VN.n5 B 0.021379f
C168 VN.n6 B 0.031345f
C169 VN.n7 B 0.244468f
C170 VN.t2 B 1.36847f
C171 VN.t4 B 1.59604f
C172 VN.n8 B 0.541828f
C173 VN.n9 B 0.574576f
C174 VN.n10 B 0.038067f
C175 VN.n11 B 0.040045f
C176 VN.n12 B 0.021379f
C177 VN.n13 B 0.021379f
C178 VN.n14 B 0.021379f
C179 VN.n15 B 0.031345f
C180 VN.n16 B 0.040045f
C181 VN.n17 B 0.038067f
C182 VN.n18 B 0.021379f
C183 VN.n19 B 0.021379f
C184 VN.n20 B 0.02225f
C185 VN.n21 B 0.040045f
C186 VN.n22 B 0.041097f
C187 VN.n23 B 0.021379f
C188 VN.n24 B 0.021379f
C189 VN.n25 B 0.021379f
C190 VN.n26 B 0.037179f
C191 VN.n27 B 0.040045f
C192 VN.n28 B 0.034113f
C193 VN.n29 B 0.034511f
C194 VN.n30 B 0.047711f
C195 VN.t3 B 1.36847f
C196 VN.n31 B 0.579379f
C197 VN.n32 B 0.021379f
C198 VN.n33 B 0.02446f
C199 VN.n34 B 0.021379f
C200 VN.t5 B 1.36847f
C201 VN.n35 B 0.496776f
C202 VN.n36 B 0.021379f
C203 VN.n37 B 0.031345f
C204 VN.n38 B 0.244468f
C205 VN.t1 B 1.36847f
C206 VN.t7 B 1.59604f
C207 VN.n39 B 0.541828f
C208 VN.n40 B 0.574576f
C209 VN.n41 B 0.038067f
C210 VN.n42 B 0.040045f
C211 VN.n43 B 0.021379f
C212 VN.n44 B 0.021379f
C213 VN.n45 B 0.021379f
C214 VN.n46 B 0.031345f
C215 VN.n47 B 0.040045f
C216 VN.n48 B 0.038067f
C217 VN.n49 B 0.021379f
C218 VN.n50 B 0.021379f
C219 VN.n51 B 0.02225f
C220 VN.n52 B 0.040045f
C221 VN.n53 B 0.041097f
C222 VN.n54 B 0.021379f
C223 VN.n55 B 0.021379f
C224 VN.n56 B 0.021379f
C225 VN.n57 B 0.037179f
C226 VN.n58 B 0.040045f
C227 VN.n59 B 0.034113f
C228 VN.n60 B 0.034511f
C229 VN.n61 B 1.2198f
.ends

