* NGSPICE file created from diff_pair_sample_0081.ext - technology: sky130A

.subckt diff_pair_sample_0081 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=2.5623 pd=13.92 as=0 ps=0 w=6.57 l=3.91
X1 VDD1.t5 VP.t0 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=2.5623 pd=13.92 as=1.08405 ps=6.9 w=6.57 l=3.91
X2 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=2.5623 pd=13.92 as=0 ps=0 w=6.57 l=3.91
X3 VDD1.t4 VP.t1 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=1.08405 pd=6.9 as=2.5623 ps=13.92 w=6.57 l=3.91
X4 VTAIL.t2 VN.t0 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.08405 pd=6.9 as=1.08405 ps=6.9 w=6.57 l=3.91
X5 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=2.5623 pd=13.92 as=0 ps=0 w=6.57 l=3.91
X6 VDD2.t4 VN.t1 VTAIL.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.08405 pd=6.9 as=2.5623 ps=13.92 w=6.57 l=3.91
X7 VTAIL.t5 VN.t2 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.08405 pd=6.9 as=1.08405 ps=6.9 w=6.57 l=3.91
X8 VDD2.t2 VN.t3 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.08405 pd=6.9 as=2.5623 ps=13.92 w=6.57 l=3.91
X9 VDD2.t1 VN.t4 VTAIL.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5623 pd=13.92 as=1.08405 ps=6.9 w=6.57 l=3.91
X10 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.5623 pd=13.92 as=0 ps=0 w=6.57 l=3.91
X11 VTAIL.t9 VP.t2 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.08405 pd=6.9 as=1.08405 ps=6.9 w=6.57 l=3.91
X12 VDD1.t2 VP.t3 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=1.08405 pd=6.9 as=2.5623 ps=13.92 w=6.57 l=3.91
X13 VDD2.t0 VN.t5 VTAIL.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.5623 pd=13.92 as=1.08405 ps=6.9 w=6.57 l=3.91
X14 VDD1.t1 VP.t4 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5623 pd=13.92 as=1.08405 ps=6.9 w=6.57 l=3.91
X15 VTAIL.t10 VP.t5 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.08405 pd=6.9 as=1.08405 ps=6.9 w=6.57 l=3.91
R0 B.n662 B.n661 585
R1 B.n662 B.n106 585
R2 B.n665 B.n664 585
R3 B.n666 B.n141 585
R4 B.n668 B.n667 585
R5 B.n670 B.n140 585
R6 B.n673 B.n672 585
R7 B.n674 B.n139 585
R8 B.n676 B.n675 585
R9 B.n678 B.n138 585
R10 B.n681 B.n680 585
R11 B.n682 B.n137 585
R12 B.n684 B.n683 585
R13 B.n686 B.n136 585
R14 B.n689 B.n688 585
R15 B.n690 B.n135 585
R16 B.n692 B.n691 585
R17 B.n694 B.n134 585
R18 B.n697 B.n696 585
R19 B.n698 B.n133 585
R20 B.n700 B.n699 585
R21 B.n702 B.n132 585
R22 B.n705 B.n704 585
R23 B.n706 B.n131 585
R24 B.n708 B.n707 585
R25 B.n710 B.n130 585
R26 B.n713 B.n712 585
R27 B.n715 B.n127 585
R28 B.n717 B.n716 585
R29 B.n719 B.n126 585
R30 B.n722 B.n721 585
R31 B.n723 B.n125 585
R32 B.n725 B.n724 585
R33 B.n727 B.n124 585
R34 B.n729 B.n728 585
R35 B.n731 B.n730 585
R36 B.n734 B.n733 585
R37 B.n735 B.n119 585
R38 B.n737 B.n736 585
R39 B.n739 B.n118 585
R40 B.n742 B.n741 585
R41 B.n743 B.n117 585
R42 B.n745 B.n744 585
R43 B.n747 B.n116 585
R44 B.n750 B.n749 585
R45 B.n751 B.n115 585
R46 B.n753 B.n752 585
R47 B.n755 B.n114 585
R48 B.n758 B.n757 585
R49 B.n759 B.n113 585
R50 B.n761 B.n760 585
R51 B.n763 B.n112 585
R52 B.n766 B.n765 585
R53 B.n767 B.n111 585
R54 B.n769 B.n768 585
R55 B.n771 B.n110 585
R56 B.n774 B.n773 585
R57 B.n775 B.n109 585
R58 B.n777 B.n776 585
R59 B.n779 B.n108 585
R60 B.n782 B.n781 585
R61 B.n783 B.n107 585
R62 B.n660 B.n105 585
R63 B.n786 B.n105 585
R64 B.n659 B.n104 585
R65 B.n787 B.n104 585
R66 B.n658 B.n103 585
R67 B.n788 B.n103 585
R68 B.n657 B.n656 585
R69 B.n656 B.n99 585
R70 B.n655 B.n98 585
R71 B.n794 B.n98 585
R72 B.n654 B.n97 585
R73 B.n795 B.n97 585
R74 B.n653 B.n96 585
R75 B.n796 B.n96 585
R76 B.n652 B.n651 585
R77 B.n651 B.n92 585
R78 B.n650 B.n91 585
R79 B.n802 B.n91 585
R80 B.n649 B.n90 585
R81 B.n803 B.n90 585
R82 B.n648 B.n89 585
R83 B.n804 B.n89 585
R84 B.n647 B.n646 585
R85 B.n646 B.n85 585
R86 B.n645 B.n84 585
R87 B.n810 B.n84 585
R88 B.n644 B.n83 585
R89 B.n811 B.n83 585
R90 B.n643 B.n82 585
R91 B.n812 B.n82 585
R92 B.n642 B.n641 585
R93 B.n641 B.n78 585
R94 B.n640 B.n77 585
R95 B.n818 B.n77 585
R96 B.n639 B.n76 585
R97 B.n819 B.n76 585
R98 B.n638 B.n75 585
R99 B.n820 B.n75 585
R100 B.n637 B.n636 585
R101 B.n636 B.n71 585
R102 B.n635 B.n70 585
R103 B.n826 B.n70 585
R104 B.n634 B.n69 585
R105 B.n827 B.n69 585
R106 B.n633 B.n68 585
R107 B.n828 B.n68 585
R108 B.n632 B.n631 585
R109 B.n631 B.n64 585
R110 B.n630 B.n63 585
R111 B.n834 B.n63 585
R112 B.n629 B.n62 585
R113 B.n835 B.n62 585
R114 B.n628 B.n61 585
R115 B.n836 B.n61 585
R116 B.n627 B.n626 585
R117 B.n626 B.n57 585
R118 B.n625 B.n56 585
R119 B.n842 B.n56 585
R120 B.n624 B.n55 585
R121 B.n843 B.n55 585
R122 B.n623 B.n54 585
R123 B.n844 B.n54 585
R124 B.n622 B.n621 585
R125 B.n621 B.n50 585
R126 B.n620 B.n49 585
R127 B.n850 B.n49 585
R128 B.n619 B.n48 585
R129 B.n851 B.n48 585
R130 B.n618 B.n47 585
R131 B.n852 B.n47 585
R132 B.n617 B.n616 585
R133 B.n616 B.n43 585
R134 B.n615 B.n42 585
R135 B.n858 B.n42 585
R136 B.n614 B.n41 585
R137 B.n859 B.n41 585
R138 B.n613 B.n40 585
R139 B.n860 B.n40 585
R140 B.n612 B.n611 585
R141 B.n611 B.n36 585
R142 B.n610 B.n35 585
R143 B.n866 B.n35 585
R144 B.n609 B.n34 585
R145 B.n867 B.n34 585
R146 B.n608 B.n33 585
R147 B.n868 B.n33 585
R148 B.n607 B.n606 585
R149 B.n606 B.n29 585
R150 B.n605 B.n28 585
R151 B.n874 B.n28 585
R152 B.n604 B.n27 585
R153 B.n875 B.n27 585
R154 B.n603 B.n26 585
R155 B.n876 B.n26 585
R156 B.n602 B.n601 585
R157 B.n601 B.n22 585
R158 B.n600 B.n21 585
R159 B.n882 B.n21 585
R160 B.n599 B.n20 585
R161 B.n883 B.n20 585
R162 B.n598 B.n19 585
R163 B.n884 B.n19 585
R164 B.n597 B.n596 585
R165 B.n596 B.n15 585
R166 B.n595 B.n14 585
R167 B.n890 B.n14 585
R168 B.n594 B.n13 585
R169 B.n891 B.n13 585
R170 B.n593 B.n12 585
R171 B.n892 B.n12 585
R172 B.n592 B.n591 585
R173 B.n591 B.n8 585
R174 B.n590 B.n7 585
R175 B.n898 B.n7 585
R176 B.n589 B.n6 585
R177 B.n899 B.n6 585
R178 B.n588 B.n5 585
R179 B.n900 B.n5 585
R180 B.n587 B.n586 585
R181 B.n586 B.n4 585
R182 B.n585 B.n142 585
R183 B.n585 B.n584 585
R184 B.n575 B.n143 585
R185 B.n144 B.n143 585
R186 B.n577 B.n576 585
R187 B.n578 B.n577 585
R188 B.n574 B.n149 585
R189 B.n149 B.n148 585
R190 B.n573 B.n572 585
R191 B.n572 B.n571 585
R192 B.n151 B.n150 585
R193 B.n152 B.n151 585
R194 B.n564 B.n563 585
R195 B.n565 B.n564 585
R196 B.n562 B.n157 585
R197 B.n157 B.n156 585
R198 B.n561 B.n560 585
R199 B.n560 B.n559 585
R200 B.n159 B.n158 585
R201 B.n160 B.n159 585
R202 B.n552 B.n551 585
R203 B.n553 B.n552 585
R204 B.n550 B.n165 585
R205 B.n165 B.n164 585
R206 B.n549 B.n548 585
R207 B.n548 B.n547 585
R208 B.n167 B.n166 585
R209 B.n168 B.n167 585
R210 B.n540 B.n539 585
R211 B.n541 B.n540 585
R212 B.n538 B.n173 585
R213 B.n173 B.n172 585
R214 B.n537 B.n536 585
R215 B.n536 B.n535 585
R216 B.n175 B.n174 585
R217 B.n176 B.n175 585
R218 B.n528 B.n527 585
R219 B.n529 B.n528 585
R220 B.n526 B.n180 585
R221 B.n184 B.n180 585
R222 B.n525 B.n524 585
R223 B.n524 B.n523 585
R224 B.n182 B.n181 585
R225 B.n183 B.n182 585
R226 B.n516 B.n515 585
R227 B.n517 B.n516 585
R228 B.n514 B.n189 585
R229 B.n189 B.n188 585
R230 B.n513 B.n512 585
R231 B.n512 B.n511 585
R232 B.n191 B.n190 585
R233 B.n192 B.n191 585
R234 B.n504 B.n503 585
R235 B.n505 B.n504 585
R236 B.n502 B.n197 585
R237 B.n197 B.n196 585
R238 B.n501 B.n500 585
R239 B.n500 B.n499 585
R240 B.n199 B.n198 585
R241 B.n200 B.n199 585
R242 B.n492 B.n491 585
R243 B.n493 B.n492 585
R244 B.n490 B.n204 585
R245 B.n208 B.n204 585
R246 B.n489 B.n488 585
R247 B.n488 B.n487 585
R248 B.n206 B.n205 585
R249 B.n207 B.n206 585
R250 B.n480 B.n479 585
R251 B.n481 B.n480 585
R252 B.n478 B.n213 585
R253 B.n213 B.n212 585
R254 B.n477 B.n476 585
R255 B.n476 B.n475 585
R256 B.n215 B.n214 585
R257 B.n216 B.n215 585
R258 B.n468 B.n467 585
R259 B.n469 B.n468 585
R260 B.n466 B.n221 585
R261 B.n221 B.n220 585
R262 B.n465 B.n464 585
R263 B.n464 B.n463 585
R264 B.n223 B.n222 585
R265 B.n224 B.n223 585
R266 B.n456 B.n455 585
R267 B.n457 B.n456 585
R268 B.n454 B.n229 585
R269 B.n229 B.n228 585
R270 B.n453 B.n452 585
R271 B.n452 B.n451 585
R272 B.n231 B.n230 585
R273 B.n232 B.n231 585
R274 B.n444 B.n443 585
R275 B.n445 B.n444 585
R276 B.n442 B.n236 585
R277 B.n240 B.n236 585
R278 B.n441 B.n440 585
R279 B.n440 B.n439 585
R280 B.n238 B.n237 585
R281 B.n239 B.n238 585
R282 B.n432 B.n431 585
R283 B.n433 B.n432 585
R284 B.n430 B.n245 585
R285 B.n245 B.n244 585
R286 B.n429 B.n428 585
R287 B.n428 B.n427 585
R288 B.n247 B.n246 585
R289 B.n248 B.n247 585
R290 B.n420 B.n419 585
R291 B.n421 B.n420 585
R292 B.n418 B.n253 585
R293 B.n253 B.n252 585
R294 B.n417 B.n416 585
R295 B.n416 B.n415 585
R296 B.n412 B.n257 585
R297 B.n411 B.n410 585
R298 B.n408 B.n258 585
R299 B.n408 B.n256 585
R300 B.n407 B.n406 585
R301 B.n405 B.n404 585
R302 B.n403 B.n260 585
R303 B.n401 B.n400 585
R304 B.n399 B.n261 585
R305 B.n398 B.n397 585
R306 B.n395 B.n262 585
R307 B.n393 B.n392 585
R308 B.n391 B.n263 585
R309 B.n390 B.n389 585
R310 B.n387 B.n264 585
R311 B.n385 B.n384 585
R312 B.n383 B.n265 585
R313 B.n382 B.n381 585
R314 B.n379 B.n266 585
R315 B.n377 B.n376 585
R316 B.n375 B.n267 585
R317 B.n374 B.n373 585
R318 B.n371 B.n268 585
R319 B.n369 B.n368 585
R320 B.n367 B.n269 585
R321 B.n366 B.n365 585
R322 B.n363 B.n270 585
R323 B.n361 B.n360 585
R324 B.n359 B.n271 585
R325 B.n358 B.n357 585
R326 B.n355 B.n275 585
R327 B.n353 B.n352 585
R328 B.n351 B.n276 585
R329 B.n350 B.n349 585
R330 B.n347 B.n277 585
R331 B.n345 B.n344 585
R332 B.n342 B.n278 585
R333 B.n341 B.n340 585
R334 B.n338 B.n281 585
R335 B.n336 B.n335 585
R336 B.n334 B.n282 585
R337 B.n333 B.n332 585
R338 B.n330 B.n283 585
R339 B.n328 B.n327 585
R340 B.n326 B.n284 585
R341 B.n325 B.n324 585
R342 B.n322 B.n285 585
R343 B.n320 B.n319 585
R344 B.n318 B.n286 585
R345 B.n317 B.n316 585
R346 B.n314 B.n287 585
R347 B.n312 B.n311 585
R348 B.n310 B.n288 585
R349 B.n309 B.n308 585
R350 B.n306 B.n289 585
R351 B.n304 B.n303 585
R352 B.n302 B.n290 585
R353 B.n301 B.n300 585
R354 B.n298 B.n291 585
R355 B.n296 B.n295 585
R356 B.n294 B.n293 585
R357 B.n255 B.n254 585
R358 B.n414 B.n413 585
R359 B.n415 B.n414 585
R360 B.n251 B.n250 585
R361 B.n252 B.n251 585
R362 B.n423 B.n422 585
R363 B.n422 B.n421 585
R364 B.n424 B.n249 585
R365 B.n249 B.n248 585
R366 B.n426 B.n425 585
R367 B.n427 B.n426 585
R368 B.n243 B.n242 585
R369 B.n244 B.n243 585
R370 B.n435 B.n434 585
R371 B.n434 B.n433 585
R372 B.n436 B.n241 585
R373 B.n241 B.n239 585
R374 B.n438 B.n437 585
R375 B.n439 B.n438 585
R376 B.n235 B.n234 585
R377 B.n240 B.n235 585
R378 B.n447 B.n446 585
R379 B.n446 B.n445 585
R380 B.n448 B.n233 585
R381 B.n233 B.n232 585
R382 B.n450 B.n449 585
R383 B.n451 B.n450 585
R384 B.n227 B.n226 585
R385 B.n228 B.n227 585
R386 B.n459 B.n458 585
R387 B.n458 B.n457 585
R388 B.n460 B.n225 585
R389 B.n225 B.n224 585
R390 B.n462 B.n461 585
R391 B.n463 B.n462 585
R392 B.n219 B.n218 585
R393 B.n220 B.n219 585
R394 B.n471 B.n470 585
R395 B.n470 B.n469 585
R396 B.n472 B.n217 585
R397 B.n217 B.n216 585
R398 B.n474 B.n473 585
R399 B.n475 B.n474 585
R400 B.n211 B.n210 585
R401 B.n212 B.n211 585
R402 B.n483 B.n482 585
R403 B.n482 B.n481 585
R404 B.n484 B.n209 585
R405 B.n209 B.n207 585
R406 B.n486 B.n485 585
R407 B.n487 B.n486 585
R408 B.n203 B.n202 585
R409 B.n208 B.n203 585
R410 B.n495 B.n494 585
R411 B.n494 B.n493 585
R412 B.n496 B.n201 585
R413 B.n201 B.n200 585
R414 B.n498 B.n497 585
R415 B.n499 B.n498 585
R416 B.n195 B.n194 585
R417 B.n196 B.n195 585
R418 B.n507 B.n506 585
R419 B.n506 B.n505 585
R420 B.n508 B.n193 585
R421 B.n193 B.n192 585
R422 B.n510 B.n509 585
R423 B.n511 B.n510 585
R424 B.n187 B.n186 585
R425 B.n188 B.n187 585
R426 B.n519 B.n518 585
R427 B.n518 B.n517 585
R428 B.n520 B.n185 585
R429 B.n185 B.n183 585
R430 B.n522 B.n521 585
R431 B.n523 B.n522 585
R432 B.n179 B.n178 585
R433 B.n184 B.n179 585
R434 B.n531 B.n530 585
R435 B.n530 B.n529 585
R436 B.n532 B.n177 585
R437 B.n177 B.n176 585
R438 B.n534 B.n533 585
R439 B.n535 B.n534 585
R440 B.n171 B.n170 585
R441 B.n172 B.n171 585
R442 B.n543 B.n542 585
R443 B.n542 B.n541 585
R444 B.n544 B.n169 585
R445 B.n169 B.n168 585
R446 B.n546 B.n545 585
R447 B.n547 B.n546 585
R448 B.n163 B.n162 585
R449 B.n164 B.n163 585
R450 B.n555 B.n554 585
R451 B.n554 B.n553 585
R452 B.n556 B.n161 585
R453 B.n161 B.n160 585
R454 B.n558 B.n557 585
R455 B.n559 B.n558 585
R456 B.n155 B.n154 585
R457 B.n156 B.n155 585
R458 B.n567 B.n566 585
R459 B.n566 B.n565 585
R460 B.n568 B.n153 585
R461 B.n153 B.n152 585
R462 B.n570 B.n569 585
R463 B.n571 B.n570 585
R464 B.n147 B.n146 585
R465 B.n148 B.n147 585
R466 B.n580 B.n579 585
R467 B.n579 B.n578 585
R468 B.n581 B.n145 585
R469 B.n145 B.n144 585
R470 B.n583 B.n582 585
R471 B.n584 B.n583 585
R472 B.n2 B.n0 585
R473 B.n4 B.n2 585
R474 B.n3 B.n1 585
R475 B.n899 B.n3 585
R476 B.n897 B.n896 585
R477 B.n898 B.n897 585
R478 B.n895 B.n9 585
R479 B.n9 B.n8 585
R480 B.n894 B.n893 585
R481 B.n893 B.n892 585
R482 B.n11 B.n10 585
R483 B.n891 B.n11 585
R484 B.n889 B.n888 585
R485 B.n890 B.n889 585
R486 B.n887 B.n16 585
R487 B.n16 B.n15 585
R488 B.n886 B.n885 585
R489 B.n885 B.n884 585
R490 B.n18 B.n17 585
R491 B.n883 B.n18 585
R492 B.n881 B.n880 585
R493 B.n882 B.n881 585
R494 B.n879 B.n23 585
R495 B.n23 B.n22 585
R496 B.n878 B.n877 585
R497 B.n877 B.n876 585
R498 B.n25 B.n24 585
R499 B.n875 B.n25 585
R500 B.n873 B.n872 585
R501 B.n874 B.n873 585
R502 B.n871 B.n30 585
R503 B.n30 B.n29 585
R504 B.n870 B.n869 585
R505 B.n869 B.n868 585
R506 B.n32 B.n31 585
R507 B.n867 B.n32 585
R508 B.n865 B.n864 585
R509 B.n866 B.n865 585
R510 B.n863 B.n37 585
R511 B.n37 B.n36 585
R512 B.n862 B.n861 585
R513 B.n861 B.n860 585
R514 B.n39 B.n38 585
R515 B.n859 B.n39 585
R516 B.n857 B.n856 585
R517 B.n858 B.n857 585
R518 B.n855 B.n44 585
R519 B.n44 B.n43 585
R520 B.n854 B.n853 585
R521 B.n853 B.n852 585
R522 B.n46 B.n45 585
R523 B.n851 B.n46 585
R524 B.n849 B.n848 585
R525 B.n850 B.n849 585
R526 B.n847 B.n51 585
R527 B.n51 B.n50 585
R528 B.n846 B.n845 585
R529 B.n845 B.n844 585
R530 B.n53 B.n52 585
R531 B.n843 B.n53 585
R532 B.n841 B.n840 585
R533 B.n842 B.n841 585
R534 B.n839 B.n58 585
R535 B.n58 B.n57 585
R536 B.n838 B.n837 585
R537 B.n837 B.n836 585
R538 B.n60 B.n59 585
R539 B.n835 B.n60 585
R540 B.n833 B.n832 585
R541 B.n834 B.n833 585
R542 B.n831 B.n65 585
R543 B.n65 B.n64 585
R544 B.n830 B.n829 585
R545 B.n829 B.n828 585
R546 B.n67 B.n66 585
R547 B.n827 B.n67 585
R548 B.n825 B.n824 585
R549 B.n826 B.n825 585
R550 B.n823 B.n72 585
R551 B.n72 B.n71 585
R552 B.n822 B.n821 585
R553 B.n821 B.n820 585
R554 B.n74 B.n73 585
R555 B.n819 B.n74 585
R556 B.n817 B.n816 585
R557 B.n818 B.n817 585
R558 B.n815 B.n79 585
R559 B.n79 B.n78 585
R560 B.n814 B.n813 585
R561 B.n813 B.n812 585
R562 B.n81 B.n80 585
R563 B.n811 B.n81 585
R564 B.n809 B.n808 585
R565 B.n810 B.n809 585
R566 B.n807 B.n86 585
R567 B.n86 B.n85 585
R568 B.n806 B.n805 585
R569 B.n805 B.n804 585
R570 B.n88 B.n87 585
R571 B.n803 B.n88 585
R572 B.n801 B.n800 585
R573 B.n802 B.n801 585
R574 B.n799 B.n93 585
R575 B.n93 B.n92 585
R576 B.n798 B.n797 585
R577 B.n797 B.n796 585
R578 B.n95 B.n94 585
R579 B.n795 B.n95 585
R580 B.n793 B.n792 585
R581 B.n794 B.n793 585
R582 B.n791 B.n100 585
R583 B.n100 B.n99 585
R584 B.n790 B.n789 585
R585 B.n789 B.n788 585
R586 B.n102 B.n101 585
R587 B.n787 B.n102 585
R588 B.n785 B.n784 585
R589 B.n786 B.n785 585
R590 B.n902 B.n901 585
R591 B.n901 B.n900 585
R592 B.n414 B.n257 487.695
R593 B.n785 B.n107 487.695
R594 B.n416 B.n255 487.695
R595 B.n662 B.n105 487.695
R596 B.n279 B.t9 270.762
R597 B.n128 B.t18 270.762
R598 B.n272 B.t12 270.762
R599 B.n120 B.t15 270.762
R600 B.n663 B.n106 256.663
R601 B.n669 B.n106 256.663
R602 B.n671 B.n106 256.663
R603 B.n677 B.n106 256.663
R604 B.n679 B.n106 256.663
R605 B.n685 B.n106 256.663
R606 B.n687 B.n106 256.663
R607 B.n693 B.n106 256.663
R608 B.n695 B.n106 256.663
R609 B.n701 B.n106 256.663
R610 B.n703 B.n106 256.663
R611 B.n709 B.n106 256.663
R612 B.n711 B.n106 256.663
R613 B.n718 B.n106 256.663
R614 B.n720 B.n106 256.663
R615 B.n726 B.n106 256.663
R616 B.n123 B.n106 256.663
R617 B.n732 B.n106 256.663
R618 B.n738 B.n106 256.663
R619 B.n740 B.n106 256.663
R620 B.n746 B.n106 256.663
R621 B.n748 B.n106 256.663
R622 B.n754 B.n106 256.663
R623 B.n756 B.n106 256.663
R624 B.n762 B.n106 256.663
R625 B.n764 B.n106 256.663
R626 B.n770 B.n106 256.663
R627 B.n772 B.n106 256.663
R628 B.n778 B.n106 256.663
R629 B.n780 B.n106 256.663
R630 B.n409 B.n256 256.663
R631 B.n259 B.n256 256.663
R632 B.n402 B.n256 256.663
R633 B.n396 B.n256 256.663
R634 B.n394 B.n256 256.663
R635 B.n388 B.n256 256.663
R636 B.n386 B.n256 256.663
R637 B.n380 B.n256 256.663
R638 B.n378 B.n256 256.663
R639 B.n372 B.n256 256.663
R640 B.n370 B.n256 256.663
R641 B.n364 B.n256 256.663
R642 B.n362 B.n256 256.663
R643 B.n356 B.n256 256.663
R644 B.n354 B.n256 256.663
R645 B.n348 B.n256 256.663
R646 B.n346 B.n256 256.663
R647 B.n339 B.n256 256.663
R648 B.n337 B.n256 256.663
R649 B.n331 B.n256 256.663
R650 B.n329 B.n256 256.663
R651 B.n323 B.n256 256.663
R652 B.n321 B.n256 256.663
R653 B.n315 B.n256 256.663
R654 B.n313 B.n256 256.663
R655 B.n307 B.n256 256.663
R656 B.n305 B.n256 256.663
R657 B.n299 B.n256 256.663
R658 B.n297 B.n256 256.663
R659 B.n292 B.n256 256.663
R660 B.n279 B.t6 249.923
R661 B.n272 B.t10 249.923
R662 B.n120 B.t13 249.923
R663 B.n128 B.t17 249.923
R664 B.n280 B.t8 188.531
R665 B.n129 B.t19 188.531
R666 B.n273 B.t11 188.531
R667 B.n121 B.t16 188.531
R668 B.n414 B.n251 163.367
R669 B.n422 B.n251 163.367
R670 B.n422 B.n249 163.367
R671 B.n426 B.n249 163.367
R672 B.n426 B.n243 163.367
R673 B.n434 B.n243 163.367
R674 B.n434 B.n241 163.367
R675 B.n438 B.n241 163.367
R676 B.n438 B.n235 163.367
R677 B.n446 B.n235 163.367
R678 B.n446 B.n233 163.367
R679 B.n450 B.n233 163.367
R680 B.n450 B.n227 163.367
R681 B.n458 B.n227 163.367
R682 B.n458 B.n225 163.367
R683 B.n462 B.n225 163.367
R684 B.n462 B.n219 163.367
R685 B.n470 B.n219 163.367
R686 B.n470 B.n217 163.367
R687 B.n474 B.n217 163.367
R688 B.n474 B.n211 163.367
R689 B.n482 B.n211 163.367
R690 B.n482 B.n209 163.367
R691 B.n486 B.n209 163.367
R692 B.n486 B.n203 163.367
R693 B.n494 B.n203 163.367
R694 B.n494 B.n201 163.367
R695 B.n498 B.n201 163.367
R696 B.n498 B.n195 163.367
R697 B.n506 B.n195 163.367
R698 B.n506 B.n193 163.367
R699 B.n510 B.n193 163.367
R700 B.n510 B.n187 163.367
R701 B.n518 B.n187 163.367
R702 B.n518 B.n185 163.367
R703 B.n522 B.n185 163.367
R704 B.n522 B.n179 163.367
R705 B.n530 B.n179 163.367
R706 B.n530 B.n177 163.367
R707 B.n534 B.n177 163.367
R708 B.n534 B.n171 163.367
R709 B.n542 B.n171 163.367
R710 B.n542 B.n169 163.367
R711 B.n546 B.n169 163.367
R712 B.n546 B.n163 163.367
R713 B.n554 B.n163 163.367
R714 B.n554 B.n161 163.367
R715 B.n558 B.n161 163.367
R716 B.n558 B.n155 163.367
R717 B.n566 B.n155 163.367
R718 B.n566 B.n153 163.367
R719 B.n570 B.n153 163.367
R720 B.n570 B.n147 163.367
R721 B.n579 B.n147 163.367
R722 B.n579 B.n145 163.367
R723 B.n583 B.n145 163.367
R724 B.n583 B.n2 163.367
R725 B.n901 B.n2 163.367
R726 B.n901 B.n3 163.367
R727 B.n897 B.n3 163.367
R728 B.n897 B.n9 163.367
R729 B.n893 B.n9 163.367
R730 B.n893 B.n11 163.367
R731 B.n889 B.n11 163.367
R732 B.n889 B.n16 163.367
R733 B.n885 B.n16 163.367
R734 B.n885 B.n18 163.367
R735 B.n881 B.n18 163.367
R736 B.n881 B.n23 163.367
R737 B.n877 B.n23 163.367
R738 B.n877 B.n25 163.367
R739 B.n873 B.n25 163.367
R740 B.n873 B.n30 163.367
R741 B.n869 B.n30 163.367
R742 B.n869 B.n32 163.367
R743 B.n865 B.n32 163.367
R744 B.n865 B.n37 163.367
R745 B.n861 B.n37 163.367
R746 B.n861 B.n39 163.367
R747 B.n857 B.n39 163.367
R748 B.n857 B.n44 163.367
R749 B.n853 B.n44 163.367
R750 B.n853 B.n46 163.367
R751 B.n849 B.n46 163.367
R752 B.n849 B.n51 163.367
R753 B.n845 B.n51 163.367
R754 B.n845 B.n53 163.367
R755 B.n841 B.n53 163.367
R756 B.n841 B.n58 163.367
R757 B.n837 B.n58 163.367
R758 B.n837 B.n60 163.367
R759 B.n833 B.n60 163.367
R760 B.n833 B.n65 163.367
R761 B.n829 B.n65 163.367
R762 B.n829 B.n67 163.367
R763 B.n825 B.n67 163.367
R764 B.n825 B.n72 163.367
R765 B.n821 B.n72 163.367
R766 B.n821 B.n74 163.367
R767 B.n817 B.n74 163.367
R768 B.n817 B.n79 163.367
R769 B.n813 B.n79 163.367
R770 B.n813 B.n81 163.367
R771 B.n809 B.n81 163.367
R772 B.n809 B.n86 163.367
R773 B.n805 B.n86 163.367
R774 B.n805 B.n88 163.367
R775 B.n801 B.n88 163.367
R776 B.n801 B.n93 163.367
R777 B.n797 B.n93 163.367
R778 B.n797 B.n95 163.367
R779 B.n793 B.n95 163.367
R780 B.n793 B.n100 163.367
R781 B.n789 B.n100 163.367
R782 B.n789 B.n102 163.367
R783 B.n785 B.n102 163.367
R784 B.n410 B.n408 163.367
R785 B.n408 B.n407 163.367
R786 B.n404 B.n403 163.367
R787 B.n401 B.n261 163.367
R788 B.n397 B.n395 163.367
R789 B.n393 B.n263 163.367
R790 B.n389 B.n387 163.367
R791 B.n385 B.n265 163.367
R792 B.n381 B.n379 163.367
R793 B.n377 B.n267 163.367
R794 B.n373 B.n371 163.367
R795 B.n369 B.n269 163.367
R796 B.n365 B.n363 163.367
R797 B.n361 B.n271 163.367
R798 B.n357 B.n355 163.367
R799 B.n353 B.n276 163.367
R800 B.n349 B.n347 163.367
R801 B.n345 B.n278 163.367
R802 B.n340 B.n338 163.367
R803 B.n336 B.n282 163.367
R804 B.n332 B.n330 163.367
R805 B.n328 B.n284 163.367
R806 B.n324 B.n322 163.367
R807 B.n320 B.n286 163.367
R808 B.n316 B.n314 163.367
R809 B.n312 B.n288 163.367
R810 B.n308 B.n306 163.367
R811 B.n304 B.n290 163.367
R812 B.n300 B.n298 163.367
R813 B.n296 B.n293 163.367
R814 B.n416 B.n253 163.367
R815 B.n420 B.n253 163.367
R816 B.n420 B.n247 163.367
R817 B.n428 B.n247 163.367
R818 B.n428 B.n245 163.367
R819 B.n432 B.n245 163.367
R820 B.n432 B.n238 163.367
R821 B.n440 B.n238 163.367
R822 B.n440 B.n236 163.367
R823 B.n444 B.n236 163.367
R824 B.n444 B.n231 163.367
R825 B.n452 B.n231 163.367
R826 B.n452 B.n229 163.367
R827 B.n456 B.n229 163.367
R828 B.n456 B.n223 163.367
R829 B.n464 B.n223 163.367
R830 B.n464 B.n221 163.367
R831 B.n468 B.n221 163.367
R832 B.n468 B.n215 163.367
R833 B.n476 B.n215 163.367
R834 B.n476 B.n213 163.367
R835 B.n480 B.n213 163.367
R836 B.n480 B.n206 163.367
R837 B.n488 B.n206 163.367
R838 B.n488 B.n204 163.367
R839 B.n492 B.n204 163.367
R840 B.n492 B.n199 163.367
R841 B.n500 B.n199 163.367
R842 B.n500 B.n197 163.367
R843 B.n504 B.n197 163.367
R844 B.n504 B.n191 163.367
R845 B.n512 B.n191 163.367
R846 B.n512 B.n189 163.367
R847 B.n516 B.n189 163.367
R848 B.n516 B.n182 163.367
R849 B.n524 B.n182 163.367
R850 B.n524 B.n180 163.367
R851 B.n528 B.n180 163.367
R852 B.n528 B.n175 163.367
R853 B.n536 B.n175 163.367
R854 B.n536 B.n173 163.367
R855 B.n540 B.n173 163.367
R856 B.n540 B.n167 163.367
R857 B.n548 B.n167 163.367
R858 B.n548 B.n165 163.367
R859 B.n552 B.n165 163.367
R860 B.n552 B.n159 163.367
R861 B.n560 B.n159 163.367
R862 B.n560 B.n157 163.367
R863 B.n564 B.n157 163.367
R864 B.n564 B.n151 163.367
R865 B.n572 B.n151 163.367
R866 B.n572 B.n149 163.367
R867 B.n577 B.n149 163.367
R868 B.n577 B.n143 163.367
R869 B.n585 B.n143 163.367
R870 B.n586 B.n585 163.367
R871 B.n586 B.n5 163.367
R872 B.n6 B.n5 163.367
R873 B.n7 B.n6 163.367
R874 B.n591 B.n7 163.367
R875 B.n591 B.n12 163.367
R876 B.n13 B.n12 163.367
R877 B.n14 B.n13 163.367
R878 B.n596 B.n14 163.367
R879 B.n596 B.n19 163.367
R880 B.n20 B.n19 163.367
R881 B.n21 B.n20 163.367
R882 B.n601 B.n21 163.367
R883 B.n601 B.n26 163.367
R884 B.n27 B.n26 163.367
R885 B.n28 B.n27 163.367
R886 B.n606 B.n28 163.367
R887 B.n606 B.n33 163.367
R888 B.n34 B.n33 163.367
R889 B.n35 B.n34 163.367
R890 B.n611 B.n35 163.367
R891 B.n611 B.n40 163.367
R892 B.n41 B.n40 163.367
R893 B.n42 B.n41 163.367
R894 B.n616 B.n42 163.367
R895 B.n616 B.n47 163.367
R896 B.n48 B.n47 163.367
R897 B.n49 B.n48 163.367
R898 B.n621 B.n49 163.367
R899 B.n621 B.n54 163.367
R900 B.n55 B.n54 163.367
R901 B.n56 B.n55 163.367
R902 B.n626 B.n56 163.367
R903 B.n626 B.n61 163.367
R904 B.n62 B.n61 163.367
R905 B.n63 B.n62 163.367
R906 B.n631 B.n63 163.367
R907 B.n631 B.n68 163.367
R908 B.n69 B.n68 163.367
R909 B.n70 B.n69 163.367
R910 B.n636 B.n70 163.367
R911 B.n636 B.n75 163.367
R912 B.n76 B.n75 163.367
R913 B.n77 B.n76 163.367
R914 B.n641 B.n77 163.367
R915 B.n641 B.n82 163.367
R916 B.n83 B.n82 163.367
R917 B.n84 B.n83 163.367
R918 B.n646 B.n84 163.367
R919 B.n646 B.n89 163.367
R920 B.n90 B.n89 163.367
R921 B.n91 B.n90 163.367
R922 B.n651 B.n91 163.367
R923 B.n651 B.n96 163.367
R924 B.n97 B.n96 163.367
R925 B.n98 B.n97 163.367
R926 B.n656 B.n98 163.367
R927 B.n656 B.n103 163.367
R928 B.n104 B.n103 163.367
R929 B.n105 B.n104 163.367
R930 B.n781 B.n779 163.367
R931 B.n777 B.n109 163.367
R932 B.n773 B.n771 163.367
R933 B.n769 B.n111 163.367
R934 B.n765 B.n763 163.367
R935 B.n761 B.n113 163.367
R936 B.n757 B.n755 163.367
R937 B.n753 B.n115 163.367
R938 B.n749 B.n747 163.367
R939 B.n745 B.n117 163.367
R940 B.n741 B.n739 163.367
R941 B.n737 B.n119 163.367
R942 B.n733 B.n731 163.367
R943 B.n728 B.n727 163.367
R944 B.n725 B.n125 163.367
R945 B.n721 B.n719 163.367
R946 B.n717 B.n127 163.367
R947 B.n712 B.n710 163.367
R948 B.n708 B.n131 163.367
R949 B.n704 B.n702 163.367
R950 B.n700 B.n133 163.367
R951 B.n696 B.n694 163.367
R952 B.n692 B.n135 163.367
R953 B.n688 B.n686 163.367
R954 B.n684 B.n137 163.367
R955 B.n680 B.n678 163.367
R956 B.n676 B.n139 163.367
R957 B.n672 B.n670 163.367
R958 B.n668 B.n141 163.367
R959 B.n664 B.n662 163.367
R960 B.n415 B.n256 114.225
R961 B.n786 B.n106 114.225
R962 B.n280 B.n279 82.2308
R963 B.n273 B.n272 82.2308
R964 B.n121 B.n120 82.2308
R965 B.n129 B.n128 82.2308
R966 B.n409 B.n257 71.676
R967 B.n407 B.n259 71.676
R968 B.n403 B.n402 71.676
R969 B.n396 B.n261 71.676
R970 B.n395 B.n394 71.676
R971 B.n388 B.n263 71.676
R972 B.n387 B.n386 71.676
R973 B.n380 B.n265 71.676
R974 B.n379 B.n378 71.676
R975 B.n372 B.n267 71.676
R976 B.n371 B.n370 71.676
R977 B.n364 B.n269 71.676
R978 B.n363 B.n362 71.676
R979 B.n356 B.n271 71.676
R980 B.n355 B.n354 71.676
R981 B.n348 B.n276 71.676
R982 B.n347 B.n346 71.676
R983 B.n339 B.n278 71.676
R984 B.n338 B.n337 71.676
R985 B.n331 B.n282 71.676
R986 B.n330 B.n329 71.676
R987 B.n323 B.n284 71.676
R988 B.n322 B.n321 71.676
R989 B.n315 B.n286 71.676
R990 B.n314 B.n313 71.676
R991 B.n307 B.n288 71.676
R992 B.n306 B.n305 71.676
R993 B.n299 B.n290 71.676
R994 B.n298 B.n297 71.676
R995 B.n293 B.n292 71.676
R996 B.n780 B.n107 71.676
R997 B.n779 B.n778 71.676
R998 B.n772 B.n109 71.676
R999 B.n771 B.n770 71.676
R1000 B.n764 B.n111 71.676
R1001 B.n763 B.n762 71.676
R1002 B.n756 B.n113 71.676
R1003 B.n755 B.n754 71.676
R1004 B.n748 B.n115 71.676
R1005 B.n747 B.n746 71.676
R1006 B.n740 B.n117 71.676
R1007 B.n739 B.n738 71.676
R1008 B.n732 B.n119 71.676
R1009 B.n731 B.n123 71.676
R1010 B.n727 B.n726 71.676
R1011 B.n720 B.n125 71.676
R1012 B.n719 B.n718 71.676
R1013 B.n711 B.n127 71.676
R1014 B.n710 B.n709 71.676
R1015 B.n703 B.n131 71.676
R1016 B.n702 B.n701 71.676
R1017 B.n695 B.n133 71.676
R1018 B.n694 B.n693 71.676
R1019 B.n687 B.n135 71.676
R1020 B.n686 B.n685 71.676
R1021 B.n679 B.n137 71.676
R1022 B.n678 B.n677 71.676
R1023 B.n671 B.n139 71.676
R1024 B.n670 B.n669 71.676
R1025 B.n663 B.n141 71.676
R1026 B.n664 B.n663 71.676
R1027 B.n669 B.n668 71.676
R1028 B.n672 B.n671 71.676
R1029 B.n677 B.n676 71.676
R1030 B.n680 B.n679 71.676
R1031 B.n685 B.n684 71.676
R1032 B.n688 B.n687 71.676
R1033 B.n693 B.n692 71.676
R1034 B.n696 B.n695 71.676
R1035 B.n701 B.n700 71.676
R1036 B.n704 B.n703 71.676
R1037 B.n709 B.n708 71.676
R1038 B.n712 B.n711 71.676
R1039 B.n718 B.n717 71.676
R1040 B.n721 B.n720 71.676
R1041 B.n726 B.n725 71.676
R1042 B.n728 B.n123 71.676
R1043 B.n733 B.n732 71.676
R1044 B.n738 B.n737 71.676
R1045 B.n741 B.n740 71.676
R1046 B.n746 B.n745 71.676
R1047 B.n749 B.n748 71.676
R1048 B.n754 B.n753 71.676
R1049 B.n757 B.n756 71.676
R1050 B.n762 B.n761 71.676
R1051 B.n765 B.n764 71.676
R1052 B.n770 B.n769 71.676
R1053 B.n773 B.n772 71.676
R1054 B.n778 B.n777 71.676
R1055 B.n781 B.n780 71.676
R1056 B.n410 B.n409 71.676
R1057 B.n404 B.n259 71.676
R1058 B.n402 B.n401 71.676
R1059 B.n397 B.n396 71.676
R1060 B.n394 B.n393 71.676
R1061 B.n389 B.n388 71.676
R1062 B.n386 B.n385 71.676
R1063 B.n381 B.n380 71.676
R1064 B.n378 B.n377 71.676
R1065 B.n373 B.n372 71.676
R1066 B.n370 B.n369 71.676
R1067 B.n365 B.n364 71.676
R1068 B.n362 B.n361 71.676
R1069 B.n357 B.n356 71.676
R1070 B.n354 B.n353 71.676
R1071 B.n349 B.n348 71.676
R1072 B.n346 B.n345 71.676
R1073 B.n340 B.n339 71.676
R1074 B.n337 B.n336 71.676
R1075 B.n332 B.n331 71.676
R1076 B.n329 B.n328 71.676
R1077 B.n324 B.n323 71.676
R1078 B.n321 B.n320 71.676
R1079 B.n316 B.n315 71.676
R1080 B.n313 B.n312 71.676
R1081 B.n308 B.n307 71.676
R1082 B.n305 B.n304 71.676
R1083 B.n300 B.n299 71.676
R1084 B.n297 B.n296 71.676
R1085 B.n292 B.n255 71.676
R1086 B.n415 B.n252 63.1495
R1087 B.n421 B.n252 63.1495
R1088 B.n421 B.n248 63.1495
R1089 B.n427 B.n248 63.1495
R1090 B.n427 B.n244 63.1495
R1091 B.n433 B.n244 63.1495
R1092 B.n433 B.n239 63.1495
R1093 B.n439 B.n239 63.1495
R1094 B.n439 B.n240 63.1495
R1095 B.n445 B.n232 63.1495
R1096 B.n451 B.n232 63.1495
R1097 B.n451 B.n228 63.1495
R1098 B.n457 B.n228 63.1495
R1099 B.n457 B.n224 63.1495
R1100 B.n463 B.n224 63.1495
R1101 B.n463 B.n220 63.1495
R1102 B.n469 B.n220 63.1495
R1103 B.n469 B.n216 63.1495
R1104 B.n475 B.n216 63.1495
R1105 B.n475 B.n212 63.1495
R1106 B.n481 B.n212 63.1495
R1107 B.n481 B.n207 63.1495
R1108 B.n487 B.n207 63.1495
R1109 B.n487 B.n208 63.1495
R1110 B.n493 B.n200 63.1495
R1111 B.n499 B.n200 63.1495
R1112 B.n499 B.n196 63.1495
R1113 B.n505 B.n196 63.1495
R1114 B.n505 B.n192 63.1495
R1115 B.n511 B.n192 63.1495
R1116 B.n511 B.n188 63.1495
R1117 B.n517 B.n188 63.1495
R1118 B.n517 B.n183 63.1495
R1119 B.n523 B.n183 63.1495
R1120 B.n523 B.n184 63.1495
R1121 B.n529 B.n176 63.1495
R1122 B.n535 B.n176 63.1495
R1123 B.n535 B.n172 63.1495
R1124 B.n541 B.n172 63.1495
R1125 B.n541 B.n168 63.1495
R1126 B.n547 B.n168 63.1495
R1127 B.n547 B.n164 63.1495
R1128 B.n553 B.n164 63.1495
R1129 B.n553 B.n160 63.1495
R1130 B.n559 B.n160 63.1495
R1131 B.n559 B.n156 63.1495
R1132 B.n565 B.n156 63.1495
R1133 B.n571 B.n152 63.1495
R1134 B.n571 B.n148 63.1495
R1135 B.n578 B.n148 63.1495
R1136 B.n578 B.n144 63.1495
R1137 B.n584 B.n144 63.1495
R1138 B.n584 B.n4 63.1495
R1139 B.n900 B.n4 63.1495
R1140 B.n900 B.n899 63.1495
R1141 B.n899 B.n898 63.1495
R1142 B.n898 B.n8 63.1495
R1143 B.n892 B.n8 63.1495
R1144 B.n892 B.n891 63.1495
R1145 B.n891 B.n890 63.1495
R1146 B.n890 B.n15 63.1495
R1147 B.n884 B.n883 63.1495
R1148 B.n883 B.n882 63.1495
R1149 B.n882 B.n22 63.1495
R1150 B.n876 B.n22 63.1495
R1151 B.n876 B.n875 63.1495
R1152 B.n875 B.n874 63.1495
R1153 B.n874 B.n29 63.1495
R1154 B.n868 B.n29 63.1495
R1155 B.n868 B.n867 63.1495
R1156 B.n867 B.n866 63.1495
R1157 B.n866 B.n36 63.1495
R1158 B.n860 B.n36 63.1495
R1159 B.n859 B.n858 63.1495
R1160 B.n858 B.n43 63.1495
R1161 B.n852 B.n43 63.1495
R1162 B.n852 B.n851 63.1495
R1163 B.n851 B.n850 63.1495
R1164 B.n850 B.n50 63.1495
R1165 B.n844 B.n50 63.1495
R1166 B.n844 B.n843 63.1495
R1167 B.n843 B.n842 63.1495
R1168 B.n842 B.n57 63.1495
R1169 B.n836 B.n57 63.1495
R1170 B.n835 B.n834 63.1495
R1171 B.n834 B.n64 63.1495
R1172 B.n828 B.n64 63.1495
R1173 B.n828 B.n827 63.1495
R1174 B.n827 B.n826 63.1495
R1175 B.n826 B.n71 63.1495
R1176 B.n820 B.n71 63.1495
R1177 B.n820 B.n819 63.1495
R1178 B.n819 B.n818 63.1495
R1179 B.n818 B.n78 63.1495
R1180 B.n812 B.n78 63.1495
R1181 B.n812 B.n811 63.1495
R1182 B.n811 B.n810 63.1495
R1183 B.n810 B.n85 63.1495
R1184 B.n804 B.n85 63.1495
R1185 B.n803 B.n802 63.1495
R1186 B.n802 B.n92 63.1495
R1187 B.n796 B.n92 63.1495
R1188 B.n796 B.n795 63.1495
R1189 B.n795 B.n794 63.1495
R1190 B.n794 B.n99 63.1495
R1191 B.n788 B.n99 63.1495
R1192 B.n788 B.n787 63.1495
R1193 B.n787 B.n786 63.1495
R1194 B.n343 B.n280 59.5399
R1195 B.n274 B.n273 59.5399
R1196 B.n122 B.n121 59.5399
R1197 B.n714 B.n129 59.5399
R1198 B.t1 B.n152 52.9342
R1199 B.t5 B.n15 52.9342
R1200 B.n493 B.t2 49.2196
R1201 B.n836 B.t4 49.2196
R1202 B.n184 B.t3 43.6476
R1203 B.t0 B.n859 43.6476
R1204 B.n240 B.t7 34.361
R1205 B.t14 B.n803 34.361
R1206 B.n784 B.n783 31.6883
R1207 B.n661 B.n660 31.6883
R1208 B.n417 B.n254 31.6883
R1209 B.n413 B.n412 31.6883
R1210 B.n445 B.t7 28.789
R1211 B.n804 B.t14 28.789
R1212 B.n529 B.t3 19.5024
R1213 B.n860 B.t0 19.5024
R1214 B B.n902 18.0485
R1215 B.n208 B.t2 13.9304
R1216 B.t4 B.n835 13.9304
R1217 B.n783 B.n782 10.6151
R1218 B.n782 B.n108 10.6151
R1219 B.n776 B.n108 10.6151
R1220 B.n776 B.n775 10.6151
R1221 B.n775 B.n774 10.6151
R1222 B.n774 B.n110 10.6151
R1223 B.n768 B.n110 10.6151
R1224 B.n768 B.n767 10.6151
R1225 B.n767 B.n766 10.6151
R1226 B.n766 B.n112 10.6151
R1227 B.n760 B.n112 10.6151
R1228 B.n760 B.n759 10.6151
R1229 B.n759 B.n758 10.6151
R1230 B.n758 B.n114 10.6151
R1231 B.n752 B.n114 10.6151
R1232 B.n752 B.n751 10.6151
R1233 B.n751 B.n750 10.6151
R1234 B.n750 B.n116 10.6151
R1235 B.n744 B.n116 10.6151
R1236 B.n744 B.n743 10.6151
R1237 B.n743 B.n742 10.6151
R1238 B.n742 B.n118 10.6151
R1239 B.n736 B.n118 10.6151
R1240 B.n736 B.n735 10.6151
R1241 B.n735 B.n734 10.6151
R1242 B.n730 B.n729 10.6151
R1243 B.n729 B.n124 10.6151
R1244 B.n724 B.n124 10.6151
R1245 B.n724 B.n723 10.6151
R1246 B.n723 B.n722 10.6151
R1247 B.n722 B.n126 10.6151
R1248 B.n716 B.n126 10.6151
R1249 B.n716 B.n715 10.6151
R1250 B.n713 B.n130 10.6151
R1251 B.n707 B.n130 10.6151
R1252 B.n707 B.n706 10.6151
R1253 B.n706 B.n705 10.6151
R1254 B.n705 B.n132 10.6151
R1255 B.n699 B.n132 10.6151
R1256 B.n699 B.n698 10.6151
R1257 B.n698 B.n697 10.6151
R1258 B.n697 B.n134 10.6151
R1259 B.n691 B.n134 10.6151
R1260 B.n691 B.n690 10.6151
R1261 B.n690 B.n689 10.6151
R1262 B.n689 B.n136 10.6151
R1263 B.n683 B.n136 10.6151
R1264 B.n683 B.n682 10.6151
R1265 B.n682 B.n681 10.6151
R1266 B.n681 B.n138 10.6151
R1267 B.n675 B.n138 10.6151
R1268 B.n675 B.n674 10.6151
R1269 B.n674 B.n673 10.6151
R1270 B.n673 B.n140 10.6151
R1271 B.n667 B.n140 10.6151
R1272 B.n667 B.n666 10.6151
R1273 B.n666 B.n665 10.6151
R1274 B.n665 B.n661 10.6151
R1275 B.n418 B.n417 10.6151
R1276 B.n419 B.n418 10.6151
R1277 B.n419 B.n246 10.6151
R1278 B.n429 B.n246 10.6151
R1279 B.n430 B.n429 10.6151
R1280 B.n431 B.n430 10.6151
R1281 B.n431 B.n237 10.6151
R1282 B.n441 B.n237 10.6151
R1283 B.n442 B.n441 10.6151
R1284 B.n443 B.n442 10.6151
R1285 B.n443 B.n230 10.6151
R1286 B.n453 B.n230 10.6151
R1287 B.n454 B.n453 10.6151
R1288 B.n455 B.n454 10.6151
R1289 B.n455 B.n222 10.6151
R1290 B.n465 B.n222 10.6151
R1291 B.n466 B.n465 10.6151
R1292 B.n467 B.n466 10.6151
R1293 B.n467 B.n214 10.6151
R1294 B.n477 B.n214 10.6151
R1295 B.n478 B.n477 10.6151
R1296 B.n479 B.n478 10.6151
R1297 B.n479 B.n205 10.6151
R1298 B.n489 B.n205 10.6151
R1299 B.n490 B.n489 10.6151
R1300 B.n491 B.n490 10.6151
R1301 B.n491 B.n198 10.6151
R1302 B.n501 B.n198 10.6151
R1303 B.n502 B.n501 10.6151
R1304 B.n503 B.n502 10.6151
R1305 B.n503 B.n190 10.6151
R1306 B.n513 B.n190 10.6151
R1307 B.n514 B.n513 10.6151
R1308 B.n515 B.n514 10.6151
R1309 B.n515 B.n181 10.6151
R1310 B.n525 B.n181 10.6151
R1311 B.n526 B.n525 10.6151
R1312 B.n527 B.n526 10.6151
R1313 B.n527 B.n174 10.6151
R1314 B.n537 B.n174 10.6151
R1315 B.n538 B.n537 10.6151
R1316 B.n539 B.n538 10.6151
R1317 B.n539 B.n166 10.6151
R1318 B.n549 B.n166 10.6151
R1319 B.n550 B.n549 10.6151
R1320 B.n551 B.n550 10.6151
R1321 B.n551 B.n158 10.6151
R1322 B.n561 B.n158 10.6151
R1323 B.n562 B.n561 10.6151
R1324 B.n563 B.n562 10.6151
R1325 B.n563 B.n150 10.6151
R1326 B.n573 B.n150 10.6151
R1327 B.n574 B.n573 10.6151
R1328 B.n576 B.n574 10.6151
R1329 B.n576 B.n575 10.6151
R1330 B.n575 B.n142 10.6151
R1331 B.n587 B.n142 10.6151
R1332 B.n588 B.n587 10.6151
R1333 B.n589 B.n588 10.6151
R1334 B.n590 B.n589 10.6151
R1335 B.n592 B.n590 10.6151
R1336 B.n593 B.n592 10.6151
R1337 B.n594 B.n593 10.6151
R1338 B.n595 B.n594 10.6151
R1339 B.n597 B.n595 10.6151
R1340 B.n598 B.n597 10.6151
R1341 B.n599 B.n598 10.6151
R1342 B.n600 B.n599 10.6151
R1343 B.n602 B.n600 10.6151
R1344 B.n603 B.n602 10.6151
R1345 B.n604 B.n603 10.6151
R1346 B.n605 B.n604 10.6151
R1347 B.n607 B.n605 10.6151
R1348 B.n608 B.n607 10.6151
R1349 B.n609 B.n608 10.6151
R1350 B.n610 B.n609 10.6151
R1351 B.n612 B.n610 10.6151
R1352 B.n613 B.n612 10.6151
R1353 B.n614 B.n613 10.6151
R1354 B.n615 B.n614 10.6151
R1355 B.n617 B.n615 10.6151
R1356 B.n618 B.n617 10.6151
R1357 B.n619 B.n618 10.6151
R1358 B.n620 B.n619 10.6151
R1359 B.n622 B.n620 10.6151
R1360 B.n623 B.n622 10.6151
R1361 B.n624 B.n623 10.6151
R1362 B.n625 B.n624 10.6151
R1363 B.n627 B.n625 10.6151
R1364 B.n628 B.n627 10.6151
R1365 B.n629 B.n628 10.6151
R1366 B.n630 B.n629 10.6151
R1367 B.n632 B.n630 10.6151
R1368 B.n633 B.n632 10.6151
R1369 B.n634 B.n633 10.6151
R1370 B.n635 B.n634 10.6151
R1371 B.n637 B.n635 10.6151
R1372 B.n638 B.n637 10.6151
R1373 B.n639 B.n638 10.6151
R1374 B.n640 B.n639 10.6151
R1375 B.n642 B.n640 10.6151
R1376 B.n643 B.n642 10.6151
R1377 B.n644 B.n643 10.6151
R1378 B.n645 B.n644 10.6151
R1379 B.n647 B.n645 10.6151
R1380 B.n648 B.n647 10.6151
R1381 B.n649 B.n648 10.6151
R1382 B.n650 B.n649 10.6151
R1383 B.n652 B.n650 10.6151
R1384 B.n653 B.n652 10.6151
R1385 B.n654 B.n653 10.6151
R1386 B.n655 B.n654 10.6151
R1387 B.n657 B.n655 10.6151
R1388 B.n658 B.n657 10.6151
R1389 B.n659 B.n658 10.6151
R1390 B.n660 B.n659 10.6151
R1391 B.n412 B.n411 10.6151
R1392 B.n411 B.n258 10.6151
R1393 B.n406 B.n258 10.6151
R1394 B.n406 B.n405 10.6151
R1395 B.n405 B.n260 10.6151
R1396 B.n400 B.n260 10.6151
R1397 B.n400 B.n399 10.6151
R1398 B.n399 B.n398 10.6151
R1399 B.n398 B.n262 10.6151
R1400 B.n392 B.n262 10.6151
R1401 B.n392 B.n391 10.6151
R1402 B.n391 B.n390 10.6151
R1403 B.n390 B.n264 10.6151
R1404 B.n384 B.n264 10.6151
R1405 B.n384 B.n383 10.6151
R1406 B.n383 B.n382 10.6151
R1407 B.n382 B.n266 10.6151
R1408 B.n376 B.n266 10.6151
R1409 B.n376 B.n375 10.6151
R1410 B.n375 B.n374 10.6151
R1411 B.n374 B.n268 10.6151
R1412 B.n368 B.n268 10.6151
R1413 B.n368 B.n367 10.6151
R1414 B.n367 B.n366 10.6151
R1415 B.n366 B.n270 10.6151
R1416 B.n360 B.n359 10.6151
R1417 B.n359 B.n358 10.6151
R1418 B.n358 B.n275 10.6151
R1419 B.n352 B.n275 10.6151
R1420 B.n352 B.n351 10.6151
R1421 B.n351 B.n350 10.6151
R1422 B.n350 B.n277 10.6151
R1423 B.n344 B.n277 10.6151
R1424 B.n342 B.n341 10.6151
R1425 B.n341 B.n281 10.6151
R1426 B.n335 B.n281 10.6151
R1427 B.n335 B.n334 10.6151
R1428 B.n334 B.n333 10.6151
R1429 B.n333 B.n283 10.6151
R1430 B.n327 B.n283 10.6151
R1431 B.n327 B.n326 10.6151
R1432 B.n326 B.n325 10.6151
R1433 B.n325 B.n285 10.6151
R1434 B.n319 B.n285 10.6151
R1435 B.n319 B.n318 10.6151
R1436 B.n318 B.n317 10.6151
R1437 B.n317 B.n287 10.6151
R1438 B.n311 B.n287 10.6151
R1439 B.n311 B.n310 10.6151
R1440 B.n310 B.n309 10.6151
R1441 B.n309 B.n289 10.6151
R1442 B.n303 B.n289 10.6151
R1443 B.n303 B.n302 10.6151
R1444 B.n302 B.n301 10.6151
R1445 B.n301 B.n291 10.6151
R1446 B.n295 B.n291 10.6151
R1447 B.n295 B.n294 10.6151
R1448 B.n294 B.n254 10.6151
R1449 B.n413 B.n250 10.6151
R1450 B.n423 B.n250 10.6151
R1451 B.n424 B.n423 10.6151
R1452 B.n425 B.n424 10.6151
R1453 B.n425 B.n242 10.6151
R1454 B.n435 B.n242 10.6151
R1455 B.n436 B.n435 10.6151
R1456 B.n437 B.n436 10.6151
R1457 B.n437 B.n234 10.6151
R1458 B.n447 B.n234 10.6151
R1459 B.n448 B.n447 10.6151
R1460 B.n449 B.n448 10.6151
R1461 B.n449 B.n226 10.6151
R1462 B.n459 B.n226 10.6151
R1463 B.n460 B.n459 10.6151
R1464 B.n461 B.n460 10.6151
R1465 B.n461 B.n218 10.6151
R1466 B.n471 B.n218 10.6151
R1467 B.n472 B.n471 10.6151
R1468 B.n473 B.n472 10.6151
R1469 B.n473 B.n210 10.6151
R1470 B.n483 B.n210 10.6151
R1471 B.n484 B.n483 10.6151
R1472 B.n485 B.n484 10.6151
R1473 B.n485 B.n202 10.6151
R1474 B.n495 B.n202 10.6151
R1475 B.n496 B.n495 10.6151
R1476 B.n497 B.n496 10.6151
R1477 B.n497 B.n194 10.6151
R1478 B.n507 B.n194 10.6151
R1479 B.n508 B.n507 10.6151
R1480 B.n509 B.n508 10.6151
R1481 B.n509 B.n186 10.6151
R1482 B.n519 B.n186 10.6151
R1483 B.n520 B.n519 10.6151
R1484 B.n521 B.n520 10.6151
R1485 B.n521 B.n178 10.6151
R1486 B.n531 B.n178 10.6151
R1487 B.n532 B.n531 10.6151
R1488 B.n533 B.n532 10.6151
R1489 B.n533 B.n170 10.6151
R1490 B.n543 B.n170 10.6151
R1491 B.n544 B.n543 10.6151
R1492 B.n545 B.n544 10.6151
R1493 B.n545 B.n162 10.6151
R1494 B.n555 B.n162 10.6151
R1495 B.n556 B.n555 10.6151
R1496 B.n557 B.n556 10.6151
R1497 B.n557 B.n154 10.6151
R1498 B.n567 B.n154 10.6151
R1499 B.n568 B.n567 10.6151
R1500 B.n569 B.n568 10.6151
R1501 B.n569 B.n146 10.6151
R1502 B.n580 B.n146 10.6151
R1503 B.n581 B.n580 10.6151
R1504 B.n582 B.n581 10.6151
R1505 B.n582 B.n0 10.6151
R1506 B.n896 B.n1 10.6151
R1507 B.n896 B.n895 10.6151
R1508 B.n895 B.n894 10.6151
R1509 B.n894 B.n10 10.6151
R1510 B.n888 B.n10 10.6151
R1511 B.n888 B.n887 10.6151
R1512 B.n887 B.n886 10.6151
R1513 B.n886 B.n17 10.6151
R1514 B.n880 B.n17 10.6151
R1515 B.n880 B.n879 10.6151
R1516 B.n879 B.n878 10.6151
R1517 B.n878 B.n24 10.6151
R1518 B.n872 B.n24 10.6151
R1519 B.n872 B.n871 10.6151
R1520 B.n871 B.n870 10.6151
R1521 B.n870 B.n31 10.6151
R1522 B.n864 B.n31 10.6151
R1523 B.n864 B.n863 10.6151
R1524 B.n863 B.n862 10.6151
R1525 B.n862 B.n38 10.6151
R1526 B.n856 B.n38 10.6151
R1527 B.n856 B.n855 10.6151
R1528 B.n855 B.n854 10.6151
R1529 B.n854 B.n45 10.6151
R1530 B.n848 B.n45 10.6151
R1531 B.n848 B.n847 10.6151
R1532 B.n847 B.n846 10.6151
R1533 B.n846 B.n52 10.6151
R1534 B.n840 B.n52 10.6151
R1535 B.n840 B.n839 10.6151
R1536 B.n839 B.n838 10.6151
R1537 B.n838 B.n59 10.6151
R1538 B.n832 B.n59 10.6151
R1539 B.n832 B.n831 10.6151
R1540 B.n831 B.n830 10.6151
R1541 B.n830 B.n66 10.6151
R1542 B.n824 B.n66 10.6151
R1543 B.n824 B.n823 10.6151
R1544 B.n823 B.n822 10.6151
R1545 B.n822 B.n73 10.6151
R1546 B.n816 B.n73 10.6151
R1547 B.n816 B.n815 10.6151
R1548 B.n815 B.n814 10.6151
R1549 B.n814 B.n80 10.6151
R1550 B.n808 B.n80 10.6151
R1551 B.n808 B.n807 10.6151
R1552 B.n807 B.n806 10.6151
R1553 B.n806 B.n87 10.6151
R1554 B.n800 B.n87 10.6151
R1555 B.n800 B.n799 10.6151
R1556 B.n799 B.n798 10.6151
R1557 B.n798 B.n94 10.6151
R1558 B.n792 B.n94 10.6151
R1559 B.n792 B.n791 10.6151
R1560 B.n791 B.n790 10.6151
R1561 B.n790 B.n101 10.6151
R1562 B.n784 B.n101 10.6151
R1563 B.n565 B.t1 10.2158
R1564 B.n884 B.t5 10.2158
R1565 B.n730 B.n122 6.5566
R1566 B.n715 B.n714 6.5566
R1567 B.n360 B.n274 6.5566
R1568 B.n344 B.n343 6.5566
R1569 B.n734 B.n122 4.05904
R1570 B.n714 B.n713 4.05904
R1571 B.n274 B.n270 4.05904
R1572 B.n343 B.n342 4.05904
R1573 B.n902 B.n0 2.81026
R1574 B.n902 B.n1 2.81026
R1575 VP.n15 VP.n14 161.3
R1576 VP.n16 VP.n11 161.3
R1577 VP.n18 VP.n17 161.3
R1578 VP.n19 VP.n10 161.3
R1579 VP.n21 VP.n20 161.3
R1580 VP.n22 VP.n9 161.3
R1581 VP.n24 VP.n23 161.3
R1582 VP.n25 VP.n8 161.3
R1583 VP.n54 VP.n0 161.3
R1584 VP.n53 VP.n52 161.3
R1585 VP.n51 VP.n1 161.3
R1586 VP.n50 VP.n49 161.3
R1587 VP.n48 VP.n2 161.3
R1588 VP.n47 VP.n46 161.3
R1589 VP.n45 VP.n3 161.3
R1590 VP.n44 VP.n43 161.3
R1591 VP.n41 VP.n4 161.3
R1592 VP.n40 VP.n39 161.3
R1593 VP.n38 VP.n5 161.3
R1594 VP.n37 VP.n36 161.3
R1595 VP.n35 VP.n6 161.3
R1596 VP.n34 VP.n33 161.3
R1597 VP.n32 VP.n7 161.3
R1598 VP.n31 VP.n30 161.3
R1599 VP.n12 VP.t4 72.5349
R1600 VP.n13 VP.n12 62.9129
R1601 VP.n29 VP.n28 58.2041
R1602 VP.n56 VP.n55 58.2041
R1603 VP.n27 VP.n26 58.2041
R1604 VP.n36 VP.n35 53.1199
R1605 VP.n49 VP.n48 53.1199
R1606 VP.n20 VP.n19 53.1199
R1607 VP.n28 VP.n27 49.9813
R1608 VP.n29 VP.t0 40.4959
R1609 VP.n42 VP.t5 40.4959
R1610 VP.n55 VP.t1 40.4959
R1611 VP.n26 VP.t3 40.4959
R1612 VP.n13 VP.t2 40.4959
R1613 VP.n35 VP.n34 27.8669
R1614 VP.n49 VP.n1 27.8669
R1615 VP.n20 VP.n9 27.8669
R1616 VP.n30 VP.n7 24.4675
R1617 VP.n34 VP.n7 24.4675
R1618 VP.n36 VP.n5 24.4675
R1619 VP.n40 VP.n5 24.4675
R1620 VP.n41 VP.n40 24.4675
R1621 VP.n43 VP.n3 24.4675
R1622 VP.n47 VP.n3 24.4675
R1623 VP.n48 VP.n47 24.4675
R1624 VP.n53 VP.n1 24.4675
R1625 VP.n54 VP.n53 24.4675
R1626 VP.n24 VP.n9 24.4675
R1627 VP.n25 VP.n24 24.4675
R1628 VP.n14 VP.n11 24.4675
R1629 VP.n18 VP.n11 24.4675
R1630 VP.n19 VP.n18 24.4675
R1631 VP.n30 VP.n29 23.9782
R1632 VP.n55 VP.n54 23.9782
R1633 VP.n26 VP.n25 23.9782
R1634 VP.n42 VP.n41 12.234
R1635 VP.n43 VP.n42 12.234
R1636 VP.n14 VP.n13 12.234
R1637 VP.n15 VP.n12 2.55161
R1638 VP.n27 VP.n8 0.417535
R1639 VP.n31 VP.n28 0.417535
R1640 VP.n56 VP.n0 0.417535
R1641 VP VP.n56 0.394291
R1642 VP.n16 VP.n15 0.189894
R1643 VP.n17 VP.n16 0.189894
R1644 VP.n17 VP.n10 0.189894
R1645 VP.n21 VP.n10 0.189894
R1646 VP.n22 VP.n21 0.189894
R1647 VP.n23 VP.n22 0.189894
R1648 VP.n23 VP.n8 0.189894
R1649 VP.n32 VP.n31 0.189894
R1650 VP.n33 VP.n32 0.189894
R1651 VP.n33 VP.n6 0.189894
R1652 VP.n37 VP.n6 0.189894
R1653 VP.n38 VP.n37 0.189894
R1654 VP.n39 VP.n38 0.189894
R1655 VP.n39 VP.n4 0.189894
R1656 VP.n44 VP.n4 0.189894
R1657 VP.n45 VP.n44 0.189894
R1658 VP.n46 VP.n45 0.189894
R1659 VP.n46 VP.n2 0.189894
R1660 VP.n50 VP.n2 0.189894
R1661 VP.n51 VP.n50 0.189894
R1662 VP.n52 VP.n51 0.189894
R1663 VP.n52 VP.n0 0.189894
R1664 VTAIL.n142 VTAIL.n141 289.615
R1665 VTAIL.n34 VTAIL.n33 289.615
R1666 VTAIL.n108 VTAIL.n107 289.615
R1667 VTAIL.n72 VTAIL.n71 289.615
R1668 VTAIL.n120 VTAIL.n119 185
R1669 VTAIL.n125 VTAIL.n124 185
R1670 VTAIL.n127 VTAIL.n126 185
R1671 VTAIL.n116 VTAIL.n115 185
R1672 VTAIL.n133 VTAIL.n132 185
R1673 VTAIL.n135 VTAIL.n134 185
R1674 VTAIL.n112 VTAIL.n111 185
R1675 VTAIL.n141 VTAIL.n140 185
R1676 VTAIL.n12 VTAIL.n11 185
R1677 VTAIL.n17 VTAIL.n16 185
R1678 VTAIL.n19 VTAIL.n18 185
R1679 VTAIL.n8 VTAIL.n7 185
R1680 VTAIL.n25 VTAIL.n24 185
R1681 VTAIL.n27 VTAIL.n26 185
R1682 VTAIL.n4 VTAIL.n3 185
R1683 VTAIL.n33 VTAIL.n32 185
R1684 VTAIL.n107 VTAIL.n106 185
R1685 VTAIL.n78 VTAIL.n77 185
R1686 VTAIL.n101 VTAIL.n100 185
R1687 VTAIL.n99 VTAIL.n98 185
R1688 VTAIL.n82 VTAIL.n81 185
R1689 VTAIL.n93 VTAIL.n92 185
R1690 VTAIL.n91 VTAIL.n90 185
R1691 VTAIL.n86 VTAIL.n85 185
R1692 VTAIL.n71 VTAIL.n70 185
R1693 VTAIL.n42 VTAIL.n41 185
R1694 VTAIL.n65 VTAIL.n64 185
R1695 VTAIL.n63 VTAIL.n62 185
R1696 VTAIL.n46 VTAIL.n45 185
R1697 VTAIL.n57 VTAIL.n56 185
R1698 VTAIL.n55 VTAIL.n54 185
R1699 VTAIL.n50 VTAIL.n49 185
R1700 VTAIL.n51 VTAIL.t0 149.525
R1701 VTAIL.n121 VTAIL.t3 149.525
R1702 VTAIL.n13 VTAIL.t11 149.525
R1703 VTAIL.n87 VTAIL.t6 149.525
R1704 VTAIL.n125 VTAIL.n119 104.615
R1705 VTAIL.n126 VTAIL.n125 104.615
R1706 VTAIL.n126 VTAIL.n115 104.615
R1707 VTAIL.n133 VTAIL.n115 104.615
R1708 VTAIL.n134 VTAIL.n133 104.615
R1709 VTAIL.n134 VTAIL.n111 104.615
R1710 VTAIL.n141 VTAIL.n111 104.615
R1711 VTAIL.n17 VTAIL.n11 104.615
R1712 VTAIL.n18 VTAIL.n17 104.615
R1713 VTAIL.n18 VTAIL.n7 104.615
R1714 VTAIL.n25 VTAIL.n7 104.615
R1715 VTAIL.n26 VTAIL.n25 104.615
R1716 VTAIL.n26 VTAIL.n3 104.615
R1717 VTAIL.n33 VTAIL.n3 104.615
R1718 VTAIL.n107 VTAIL.n77 104.615
R1719 VTAIL.n100 VTAIL.n77 104.615
R1720 VTAIL.n100 VTAIL.n99 104.615
R1721 VTAIL.n99 VTAIL.n81 104.615
R1722 VTAIL.n92 VTAIL.n81 104.615
R1723 VTAIL.n92 VTAIL.n91 104.615
R1724 VTAIL.n91 VTAIL.n85 104.615
R1725 VTAIL.n71 VTAIL.n41 104.615
R1726 VTAIL.n64 VTAIL.n41 104.615
R1727 VTAIL.n64 VTAIL.n63 104.615
R1728 VTAIL.n63 VTAIL.n45 104.615
R1729 VTAIL.n56 VTAIL.n45 104.615
R1730 VTAIL.n56 VTAIL.n55 104.615
R1731 VTAIL.n55 VTAIL.n49 104.615
R1732 VTAIL.n75 VTAIL.n74 52.808
R1733 VTAIL.n39 VTAIL.n38 52.808
R1734 VTAIL.n1 VTAIL.n0 52.807
R1735 VTAIL.n37 VTAIL.n36 52.807
R1736 VTAIL.t3 VTAIL.n119 52.3082
R1737 VTAIL.t11 VTAIL.n11 52.3082
R1738 VTAIL.t6 VTAIL.n85 52.3082
R1739 VTAIL.t0 VTAIL.n49 52.3082
R1740 VTAIL.n143 VTAIL.n142 35.8702
R1741 VTAIL.n35 VTAIL.n34 35.8702
R1742 VTAIL.n109 VTAIL.n108 35.8702
R1743 VTAIL.n73 VTAIL.n72 35.8702
R1744 VTAIL.n39 VTAIL.n37 25.341
R1745 VTAIL.n143 VTAIL.n109 21.6858
R1746 VTAIL.n140 VTAIL.n110 12.8005
R1747 VTAIL.n32 VTAIL.n2 12.8005
R1748 VTAIL.n106 VTAIL.n76 12.8005
R1749 VTAIL.n70 VTAIL.n40 12.8005
R1750 VTAIL.n139 VTAIL.n112 12.0247
R1751 VTAIL.n31 VTAIL.n4 12.0247
R1752 VTAIL.n105 VTAIL.n78 12.0247
R1753 VTAIL.n69 VTAIL.n42 12.0247
R1754 VTAIL.n136 VTAIL.n135 11.249
R1755 VTAIL.n28 VTAIL.n27 11.249
R1756 VTAIL.n102 VTAIL.n101 11.249
R1757 VTAIL.n66 VTAIL.n65 11.249
R1758 VTAIL.n132 VTAIL.n114 10.4732
R1759 VTAIL.n24 VTAIL.n6 10.4732
R1760 VTAIL.n98 VTAIL.n80 10.4732
R1761 VTAIL.n62 VTAIL.n44 10.4732
R1762 VTAIL.n121 VTAIL.n120 10.2746
R1763 VTAIL.n13 VTAIL.n12 10.2746
R1764 VTAIL.n87 VTAIL.n86 10.2746
R1765 VTAIL.n51 VTAIL.n50 10.2746
R1766 VTAIL.n131 VTAIL.n116 9.69747
R1767 VTAIL.n23 VTAIL.n8 9.69747
R1768 VTAIL.n97 VTAIL.n82 9.69747
R1769 VTAIL.n61 VTAIL.n46 9.69747
R1770 VTAIL.n138 VTAIL.n110 9.45567
R1771 VTAIL.n30 VTAIL.n2 9.45567
R1772 VTAIL.n104 VTAIL.n76 9.45567
R1773 VTAIL.n68 VTAIL.n40 9.45567
R1774 VTAIL.n123 VTAIL.n122 9.3005
R1775 VTAIL.n118 VTAIL.n117 9.3005
R1776 VTAIL.n129 VTAIL.n128 9.3005
R1777 VTAIL.n131 VTAIL.n130 9.3005
R1778 VTAIL.n114 VTAIL.n113 9.3005
R1779 VTAIL.n137 VTAIL.n136 9.3005
R1780 VTAIL.n139 VTAIL.n138 9.3005
R1781 VTAIL.n15 VTAIL.n14 9.3005
R1782 VTAIL.n10 VTAIL.n9 9.3005
R1783 VTAIL.n21 VTAIL.n20 9.3005
R1784 VTAIL.n23 VTAIL.n22 9.3005
R1785 VTAIL.n6 VTAIL.n5 9.3005
R1786 VTAIL.n29 VTAIL.n28 9.3005
R1787 VTAIL.n31 VTAIL.n30 9.3005
R1788 VTAIL.n105 VTAIL.n104 9.3005
R1789 VTAIL.n103 VTAIL.n102 9.3005
R1790 VTAIL.n80 VTAIL.n79 9.3005
R1791 VTAIL.n97 VTAIL.n96 9.3005
R1792 VTAIL.n95 VTAIL.n94 9.3005
R1793 VTAIL.n84 VTAIL.n83 9.3005
R1794 VTAIL.n89 VTAIL.n88 9.3005
R1795 VTAIL.n48 VTAIL.n47 9.3005
R1796 VTAIL.n59 VTAIL.n58 9.3005
R1797 VTAIL.n61 VTAIL.n60 9.3005
R1798 VTAIL.n44 VTAIL.n43 9.3005
R1799 VTAIL.n67 VTAIL.n66 9.3005
R1800 VTAIL.n69 VTAIL.n68 9.3005
R1801 VTAIL.n53 VTAIL.n52 9.3005
R1802 VTAIL.n128 VTAIL.n127 8.92171
R1803 VTAIL.n20 VTAIL.n19 8.92171
R1804 VTAIL.n94 VTAIL.n93 8.92171
R1805 VTAIL.n58 VTAIL.n57 8.92171
R1806 VTAIL.n124 VTAIL.n118 8.14595
R1807 VTAIL.n16 VTAIL.n10 8.14595
R1808 VTAIL.n90 VTAIL.n84 8.14595
R1809 VTAIL.n54 VTAIL.n48 8.14595
R1810 VTAIL.n123 VTAIL.n120 7.3702
R1811 VTAIL.n15 VTAIL.n12 7.3702
R1812 VTAIL.n89 VTAIL.n86 7.3702
R1813 VTAIL.n53 VTAIL.n50 7.3702
R1814 VTAIL.n124 VTAIL.n123 5.81868
R1815 VTAIL.n16 VTAIL.n15 5.81868
R1816 VTAIL.n90 VTAIL.n89 5.81868
R1817 VTAIL.n54 VTAIL.n53 5.81868
R1818 VTAIL.n127 VTAIL.n118 5.04292
R1819 VTAIL.n19 VTAIL.n10 5.04292
R1820 VTAIL.n93 VTAIL.n84 5.04292
R1821 VTAIL.n57 VTAIL.n48 5.04292
R1822 VTAIL.n128 VTAIL.n116 4.26717
R1823 VTAIL.n20 VTAIL.n8 4.26717
R1824 VTAIL.n94 VTAIL.n82 4.26717
R1825 VTAIL.n58 VTAIL.n46 4.26717
R1826 VTAIL.n73 VTAIL.n39 3.65567
R1827 VTAIL.n109 VTAIL.n75 3.65567
R1828 VTAIL.n37 VTAIL.n35 3.65567
R1829 VTAIL.n132 VTAIL.n131 3.49141
R1830 VTAIL.n24 VTAIL.n23 3.49141
R1831 VTAIL.n98 VTAIL.n97 3.49141
R1832 VTAIL.n62 VTAIL.n61 3.49141
R1833 VTAIL.n0 VTAIL.t4 3.0142
R1834 VTAIL.n0 VTAIL.t2 3.0142
R1835 VTAIL.n36 VTAIL.t7 3.0142
R1836 VTAIL.n36 VTAIL.t10 3.0142
R1837 VTAIL.n74 VTAIL.t8 3.0142
R1838 VTAIL.n74 VTAIL.t9 3.0142
R1839 VTAIL.n38 VTAIL.t1 3.0142
R1840 VTAIL.n38 VTAIL.t5 3.0142
R1841 VTAIL.n52 VTAIL.n51 2.84308
R1842 VTAIL.n122 VTAIL.n121 2.84308
R1843 VTAIL.n14 VTAIL.n13 2.84308
R1844 VTAIL.n88 VTAIL.n87 2.84308
R1845 VTAIL.n135 VTAIL.n114 2.71565
R1846 VTAIL.n27 VTAIL.n6 2.71565
R1847 VTAIL.n101 VTAIL.n80 2.71565
R1848 VTAIL.n65 VTAIL.n44 2.71565
R1849 VTAIL VTAIL.n143 2.68369
R1850 VTAIL.n75 VTAIL.n73 2.29791
R1851 VTAIL.n35 VTAIL.n1 2.29791
R1852 VTAIL.n136 VTAIL.n112 1.93989
R1853 VTAIL.n28 VTAIL.n4 1.93989
R1854 VTAIL.n102 VTAIL.n78 1.93989
R1855 VTAIL.n66 VTAIL.n42 1.93989
R1856 VTAIL.n140 VTAIL.n139 1.16414
R1857 VTAIL.n32 VTAIL.n31 1.16414
R1858 VTAIL.n106 VTAIL.n105 1.16414
R1859 VTAIL.n70 VTAIL.n69 1.16414
R1860 VTAIL VTAIL.n1 0.972483
R1861 VTAIL.n142 VTAIL.n110 0.388379
R1862 VTAIL.n34 VTAIL.n2 0.388379
R1863 VTAIL.n108 VTAIL.n76 0.388379
R1864 VTAIL.n72 VTAIL.n40 0.388379
R1865 VTAIL.n122 VTAIL.n117 0.155672
R1866 VTAIL.n129 VTAIL.n117 0.155672
R1867 VTAIL.n130 VTAIL.n129 0.155672
R1868 VTAIL.n130 VTAIL.n113 0.155672
R1869 VTAIL.n137 VTAIL.n113 0.155672
R1870 VTAIL.n138 VTAIL.n137 0.155672
R1871 VTAIL.n14 VTAIL.n9 0.155672
R1872 VTAIL.n21 VTAIL.n9 0.155672
R1873 VTAIL.n22 VTAIL.n21 0.155672
R1874 VTAIL.n22 VTAIL.n5 0.155672
R1875 VTAIL.n29 VTAIL.n5 0.155672
R1876 VTAIL.n30 VTAIL.n29 0.155672
R1877 VTAIL.n104 VTAIL.n103 0.155672
R1878 VTAIL.n103 VTAIL.n79 0.155672
R1879 VTAIL.n96 VTAIL.n79 0.155672
R1880 VTAIL.n96 VTAIL.n95 0.155672
R1881 VTAIL.n95 VTAIL.n83 0.155672
R1882 VTAIL.n88 VTAIL.n83 0.155672
R1883 VTAIL.n68 VTAIL.n67 0.155672
R1884 VTAIL.n67 VTAIL.n43 0.155672
R1885 VTAIL.n60 VTAIL.n43 0.155672
R1886 VTAIL.n60 VTAIL.n59 0.155672
R1887 VTAIL.n59 VTAIL.n47 0.155672
R1888 VTAIL.n52 VTAIL.n47 0.155672
R1889 VDD1.n32 VDD1.n31 289.615
R1890 VDD1.n65 VDD1.n64 289.615
R1891 VDD1.n31 VDD1.n30 185
R1892 VDD1.n2 VDD1.n1 185
R1893 VDD1.n25 VDD1.n24 185
R1894 VDD1.n23 VDD1.n22 185
R1895 VDD1.n6 VDD1.n5 185
R1896 VDD1.n17 VDD1.n16 185
R1897 VDD1.n15 VDD1.n14 185
R1898 VDD1.n10 VDD1.n9 185
R1899 VDD1.n43 VDD1.n42 185
R1900 VDD1.n48 VDD1.n47 185
R1901 VDD1.n50 VDD1.n49 185
R1902 VDD1.n39 VDD1.n38 185
R1903 VDD1.n56 VDD1.n55 185
R1904 VDD1.n58 VDD1.n57 185
R1905 VDD1.n35 VDD1.n34 185
R1906 VDD1.n64 VDD1.n63 185
R1907 VDD1.n11 VDD1.t1 149.525
R1908 VDD1.n44 VDD1.t5 149.525
R1909 VDD1.n31 VDD1.n1 104.615
R1910 VDD1.n24 VDD1.n1 104.615
R1911 VDD1.n24 VDD1.n23 104.615
R1912 VDD1.n23 VDD1.n5 104.615
R1913 VDD1.n16 VDD1.n5 104.615
R1914 VDD1.n16 VDD1.n15 104.615
R1915 VDD1.n15 VDD1.n9 104.615
R1916 VDD1.n48 VDD1.n42 104.615
R1917 VDD1.n49 VDD1.n48 104.615
R1918 VDD1.n49 VDD1.n38 104.615
R1919 VDD1.n56 VDD1.n38 104.615
R1920 VDD1.n57 VDD1.n56 104.615
R1921 VDD1.n57 VDD1.n34 104.615
R1922 VDD1.n64 VDD1.n34 104.615
R1923 VDD1.n67 VDD1.n66 70.3442
R1924 VDD1.n69 VDD1.n68 69.4856
R1925 VDD1 VDD1.n32 55.3486
R1926 VDD1.n67 VDD1.n65 55.235
R1927 VDD1.t1 VDD1.n9 52.3082
R1928 VDD1.t5 VDD1.n42 52.3082
R1929 VDD1.n69 VDD1.n67 43.669
R1930 VDD1.n30 VDD1.n0 12.8005
R1931 VDD1.n63 VDD1.n33 12.8005
R1932 VDD1.n29 VDD1.n2 12.0247
R1933 VDD1.n62 VDD1.n35 12.0247
R1934 VDD1.n26 VDD1.n25 11.249
R1935 VDD1.n59 VDD1.n58 11.249
R1936 VDD1.n22 VDD1.n4 10.4732
R1937 VDD1.n55 VDD1.n37 10.4732
R1938 VDD1.n11 VDD1.n10 10.2746
R1939 VDD1.n44 VDD1.n43 10.2746
R1940 VDD1.n21 VDD1.n6 9.69747
R1941 VDD1.n54 VDD1.n39 9.69747
R1942 VDD1.n28 VDD1.n0 9.45567
R1943 VDD1.n61 VDD1.n33 9.45567
R1944 VDD1.n8 VDD1.n7 9.3005
R1945 VDD1.n19 VDD1.n18 9.3005
R1946 VDD1.n21 VDD1.n20 9.3005
R1947 VDD1.n4 VDD1.n3 9.3005
R1948 VDD1.n27 VDD1.n26 9.3005
R1949 VDD1.n29 VDD1.n28 9.3005
R1950 VDD1.n13 VDD1.n12 9.3005
R1951 VDD1.n46 VDD1.n45 9.3005
R1952 VDD1.n41 VDD1.n40 9.3005
R1953 VDD1.n52 VDD1.n51 9.3005
R1954 VDD1.n54 VDD1.n53 9.3005
R1955 VDD1.n37 VDD1.n36 9.3005
R1956 VDD1.n60 VDD1.n59 9.3005
R1957 VDD1.n62 VDD1.n61 9.3005
R1958 VDD1.n18 VDD1.n17 8.92171
R1959 VDD1.n51 VDD1.n50 8.92171
R1960 VDD1.n14 VDD1.n8 8.14595
R1961 VDD1.n47 VDD1.n41 8.14595
R1962 VDD1.n13 VDD1.n10 7.3702
R1963 VDD1.n46 VDD1.n43 7.3702
R1964 VDD1.n14 VDD1.n13 5.81868
R1965 VDD1.n47 VDD1.n46 5.81868
R1966 VDD1.n17 VDD1.n8 5.04292
R1967 VDD1.n50 VDD1.n41 5.04292
R1968 VDD1.n18 VDD1.n6 4.26717
R1969 VDD1.n51 VDD1.n39 4.26717
R1970 VDD1.n22 VDD1.n21 3.49141
R1971 VDD1.n55 VDD1.n54 3.49141
R1972 VDD1.n68 VDD1.t3 3.0142
R1973 VDD1.n68 VDD1.t2 3.0142
R1974 VDD1.n66 VDD1.t0 3.0142
R1975 VDD1.n66 VDD1.t4 3.0142
R1976 VDD1.n12 VDD1.n11 2.84308
R1977 VDD1.n45 VDD1.n44 2.84308
R1978 VDD1.n25 VDD1.n4 2.71565
R1979 VDD1.n58 VDD1.n37 2.71565
R1980 VDD1.n26 VDD1.n2 1.93989
R1981 VDD1.n59 VDD1.n35 1.93989
R1982 VDD1.n30 VDD1.n29 1.16414
R1983 VDD1.n63 VDD1.n62 1.16414
R1984 VDD1 VDD1.n69 0.856103
R1985 VDD1.n32 VDD1.n0 0.388379
R1986 VDD1.n65 VDD1.n33 0.388379
R1987 VDD1.n28 VDD1.n27 0.155672
R1988 VDD1.n27 VDD1.n3 0.155672
R1989 VDD1.n20 VDD1.n3 0.155672
R1990 VDD1.n20 VDD1.n19 0.155672
R1991 VDD1.n19 VDD1.n7 0.155672
R1992 VDD1.n12 VDD1.n7 0.155672
R1993 VDD1.n45 VDD1.n40 0.155672
R1994 VDD1.n52 VDD1.n40 0.155672
R1995 VDD1.n53 VDD1.n52 0.155672
R1996 VDD1.n53 VDD1.n36 0.155672
R1997 VDD1.n60 VDD1.n36 0.155672
R1998 VDD1.n61 VDD1.n60 0.155672
R1999 VN.n37 VN.n20 161.3
R2000 VN.n36 VN.n35 161.3
R2001 VN.n34 VN.n21 161.3
R2002 VN.n33 VN.n32 161.3
R2003 VN.n31 VN.n22 161.3
R2004 VN.n30 VN.n29 161.3
R2005 VN.n28 VN.n23 161.3
R2006 VN.n27 VN.n26 161.3
R2007 VN.n17 VN.n0 161.3
R2008 VN.n16 VN.n15 161.3
R2009 VN.n14 VN.n1 161.3
R2010 VN.n13 VN.n12 161.3
R2011 VN.n11 VN.n2 161.3
R2012 VN.n10 VN.n9 161.3
R2013 VN.n8 VN.n3 161.3
R2014 VN.n7 VN.n6 161.3
R2015 VN.n4 VN.t4 72.5353
R2016 VN.n24 VN.t3 72.5353
R2017 VN.n5 VN.n4 62.9128
R2018 VN.n25 VN.n24 62.9128
R2019 VN.n19 VN.n18 58.2041
R2020 VN.n39 VN.n38 58.2041
R2021 VN.n12 VN.n11 53.1199
R2022 VN.n32 VN.n31 53.1199
R2023 VN VN.n39 50.0193
R2024 VN.n5 VN.t0 40.4959
R2025 VN.n18 VN.t1 40.4959
R2026 VN.n25 VN.t2 40.4959
R2027 VN.n38 VN.t5 40.4959
R2028 VN.n12 VN.n1 27.8669
R2029 VN.n32 VN.n21 27.8669
R2030 VN.n6 VN.n3 24.4675
R2031 VN.n10 VN.n3 24.4675
R2032 VN.n11 VN.n10 24.4675
R2033 VN.n16 VN.n1 24.4675
R2034 VN.n17 VN.n16 24.4675
R2035 VN.n31 VN.n30 24.4675
R2036 VN.n30 VN.n23 24.4675
R2037 VN.n26 VN.n23 24.4675
R2038 VN.n37 VN.n36 24.4675
R2039 VN.n36 VN.n21 24.4675
R2040 VN.n18 VN.n17 23.9782
R2041 VN.n38 VN.n37 23.9782
R2042 VN.n6 VN.n5 12.234
R2043 VN.n26 VN.n25 12.234
R2044 VN.n27 VN.n24 2.55164
R2045 VN.n7 VN.n4 2.55164
R2046 VN.n39 VN.n20 0.417535
R2047 VN.n19 VN.n0 0.417535
R2048 VN VN.n19 0.394291
R2049 VN.n35 VN.n20 0.189894
R2050 VN.n35 VN.n34 0.189894
R2051 VN.n34 VN.n33 0.189894
R2052 VN.n33 VN.n22 0.189894
R2053 VN.n29 VN.n22 0.189894
R2054 VN.n29 VN.n28 0.189894
R2055 VN.n28 VN.n27 0.189894
R2056 VN.n8 VN.n7 0.189894
R2057 VN.n9 VN.n8 0.189894
R2058 VN.n9 VN.n2 0.189894
R2059 VN.n13 VN.n2 0.189894
R2060 VN.n14 VN.n13 0.189894
R2061 VN.n15 VN.n14 0.189894
R2062 VN.n15 VN.n0 0.189894
R2063 VDD2.n67 VDD2.n66 289.615
R2064 VDD2.n32 VDD2.n31 289.615
R2065 VDD2.n66 VDD2.n65 185
R2066 VDD2.n37 VDD2.n36 185
R2067 VDD2.n60 VDD2.n59 185
R2068 VDD2.n58 VDD2.n57 185
R2069 VDD2.n41 VDD2.n40 185
R2070 VDD2.n52 VDD2.n51 185
R2071 VDD2.n50 VDD2.n49 185
R2072 VDD2.n45 VDD2.n44 185
R2073 VDD2.n10 VDD2.n9 185
R2074 VDD2.n15 VDD2.n14 185
R2075 VDD2.n17 VDD2.n16 185
R2076 VDD2.n6 VDD2.n5 185
R2077 VDD2.n23 VDD2.n22 185
R2078 VDD2.n25 VDD2.n24 185
R2079 VDD2.n2 VDD2.n1 185
R2080 VDD2.n31 VDD2.n30 185
R2081 VDD2.n46 VDD2.t0 149.525
R2082 VDD2.n11 VDD2.t1 149.525
R2083 VDD2.n66 VDD2.n36 104.615
R2084 VDD2.n59 VDD2.n36 104.615
R2085 VDD2.n59 VDD2.n58 104.615
R2086 VDD2.n58 VDD2.n40 104.615
R2087 VDD2.n51 VDD2.n40 104.615
R2088 VDD2.n51 VDD2.n50 104.615
R2089 VDD2.n50 VDD2.n44 104.615
R2090 VDD2.n15 VDD2.n9 104.615
R2091 VDD2.n16 VDD2.n15 104.615
R2092 VDD2.n16 VDD2.n5 104.615
R2093 VDD2.n23 VDD2.n5 104.615
R2094 VDD2.n24 VDD2.n23 104.615
R2095 VDD2.n24 VDD2.n1 104.615
R2096 VDD2.n31 VDD2.n1 104.615
R2097 VDD2.n34 VDD2.n33 70.3442
R2098 VDD2 VDD2.n69 70.3412
R2099 VDD2.n34 VDD2.n32 55.235
R2100 VDD2.n68 VDD2.n67 52.549
R2101 VDD2.t0 VDD2.n44 52.3082
R2102 VDD2.t1 VDD2.n9 52.3082
R2103 VDD2.n68 VDD2.n34 41.2584
R2104 VDD2.n65 VDD2.n35 12.8005
R2105 VDD2.n30 VDD2.n0 12.8005
R2106 VDD2.n64 VDD2.n37 12.0247
R2107 VDD2.n29 VDD2.n2 12.0247
R2108 VDD2.n61 VDD2.n60 11.249
R2109 VDD2.n26 VDD2.n25 11.249
R2110 VDD2.n57 VDD2.n39 10.4732
R2111 VDD2.n22 VDD2.n4 10.4732
R2112 VDD2.n46 VDD2.n45 10.2746
R2113 VDD2.n11 VDD2.n10 10.2746
R2114 VDD2.n56 VDD2.n41 9.69747
R2115 VDD2.n21 VDD2.n6 9.69747
R2116 VDD2.n63 VDD2.n35 9.45567
R2117 VDD2.n28 VDD2.n0 9.45567
R2118 VDD2.n43 VDD2.n42 9.3005
R2119 VDD2.n54 VDD2.n53 9.3005
R2120 VDD2.n56 VDD2.n55 9.3005
R2121 VDD2.n39 VDD2.n38 9.3005
R2122 VDD2.n62 VDD2.n61 9.3005
R2123 VDD2.n64 VDD2.n63 9.3005
R2124 VDD2.n48 VDD2.n47 9.3005
R2125 VDD2.n13 VDD2.n12 9.3005
R2126 VDD2.n8 VDD2.n7 9.3005
R2127 VDD2.n19 VDD2.n18 9.3005
R2128 VDD2.n21 VDD2.n20 9.3005
R2129 VDD2.n4 VDD2.n3 9.3005
R2130 VDD2.n27 VDD2.n26 9.3005
R2131 VDD2.n29 VDD2.n28 9.3005
R2132 VDD2.n53 VDD2.n52 8.92171
R2133 VDD2.n18 VDD2.n17 8.92171
R2134 VDD2.n49 VDD2.n43 8.14595
R2135 VDD2.n14 VDD2.n8 8.14595
R2136 VDD2.n48 VDD2.n45 7.3702
R2137 VDD2.n13 VDD2.n10 7.3702
R2138 VDD2.n49 VDD2.n48 5.81868
R2139 VDD2.n14 VDD2.n13 5.81868
R2140 VDD2.n52 VDD2.n43 5.04292
R2141 VDD2.n17 VDD2.n8 5.04292
R2142 VDD2.n53 VDD2.n41 4.26717
R2143 VDD2.n18 VDD2.n6 4.26717
R2144 VDD2.n57 VDD2.n56 3.49141
R2145 VDD2.n22 VDD2.n21 3.49141
R2146 VDD2.n69 VDD2.t3 3.0142
R2147 VDD2.n69 VDD2.t2 3.0142
R2148 VDD2.n33 VDD2.t5 3.0142
R2149 VDD2.n33 VDD2.t4 3.0142
R2150 VDD2.n47 VDD2.n46 2.84308
R2151 VDD2.n12 VDD2.n11 2.84308
R2152 VDD2 VDD2.n68 2.80007
R2153 VDD2.n60 VDD2.n39 2.71565
R2154 VDD2.n25 VDD2.n4 2.71565
R2155 VDD2.n61 VDD2.n37 1.93989
R2156 VDD2.n26 VDD2.n2 1.93989
R2157 VDD2.n65 VDD2.n64 1.16414
R2158 VDD2.n30 VDD2.n29 1.16414
R2159 VDD2.n67 VDD2.n35 0.388379
R2160 VDD2.n32 VDD2.n0 0.388379
R2161 VDD2.n63 VDD2.n62 0.155672
R2162 VDD2.n62 VDD2.n38 0.155672
R2163 VDD2.n55 VDD2.n38 0.155672
R2164 VDD2.n55 VDD2.n54 0.155672
R2165 VDD2.n54 VDD2.n42 0.155672
R2166 VDD2.n47 VDD2.n42 0.155672
R2167 VDD2.n12 VDD2.n7 0.155672
R2168 VDD2.n19 VDD2.n7 0.155672
R2169 VDD2.n20 VDD2.n19 0.155672
R2170 VDD2.n20 VDD2.n3 0.155672
R2171 VDD2.n27 VDD2.n3 0.155672
R2172 VDD2.n28 VDD2.n27 0.155672
C0 VP VN 7.19576f
C1 VTAIL VDD2 6.56666f
C2 VDD2 VN 4.11375f
C3 VTAIL VDD1 6.50521f
C4 VN VDD1 0.15256f
C5 VP VDD2 0.568786f
C6 VTAIL VN 5.04707f
C7 VP VDD1 4.52795f
C8 VDD2 VDD1 1.91805f
C9 VP VTAIL 5.0616f
C10 VDD2 B 6.024855f
C11 VDD1 B 6.225192f
C12 VTAIL B 5.988827f
C13 VN B 16.198881f
C14 VP B 14.909935f
C15 VDD2.n0 B 0.01233f
C16 VDD2.n1 B 0.027765f
C17 VDD2.n2 B 0.012438f
C18 VDD2.n3 B 0.02186f
C19 VDD2.n4 B 0.011747f
C20 VDD2.n5 B 0.027765f
C21 VDD2.n6 B 0.012438f
C22 VDD2.n7 B 0.02186f
C23 VDD2.n8 B 0.011747f
C24 VDD2.n9 B 0.020824f
C25 VDD2.n10 B 0.019628f
C26 VDD2.t1 B 0.046319f
C27 VDD2.n11 B 0.112154f
C28 VDD2.n12 B 0.57467f
C29 VDD2.n13 B 0.011747f
C30 VDD2.n14 B 0.012438f
C31 VDD2.n15 B 0.027765f
C32 VDD2.n16 B 0.027765f
C33 VDD2.n17 B 0.012438f
C34 VDD2.n18 B 0.011747f
C35 VDD2.n19 B 0.02186f
C36 VDD2.n20 B 0.02186f
C37 VDD2.n21 B 0.011747f
C38 VDD2.n22 B 0.012438f
C39 VDD2.n23 B 0.027765f
C40 VDD2.n24 B 0.027765f
C41 VDD2.n25 B 0.012438f
C42 VDD2.n26 B 0.011747f
C43 VDD2.n27 B 0.02186f
C44 VDD2.n28 B 0.056801f
C45 VDD2.n29 B 0.011747f
C46 VDD2.n30 B 0.012438f
C47 VDD2.n31 B 0.057238f
C48 VDD2.n32 B 0.074807f
C49 VDD2.t5 B 0.113495f
C50 VDD2.t4 B 0.113495f
C51 VDD2.n33 B 0.972022f
C52 VDD2.n34 B 2.53806f
C53 VDD2.n35 B 0.01233f
C54 VDD2.n36 B 0.027765f
C55 VDD2.n37 B 0.012438f
C56 VDD2.n38 B 0.02186f
C57 VDD2.n39 B 0.011747f
C58 VDD2.n40 B 0.027765f
C59 VDD2.n41 B 0.012438f
C60 VDD2.n42 B 0.02186f
C61 VDD2.n43 B 0.011747f
C62 VDD2.n44 B 0.020824f
C63 VDD2.n45 B 0.019628f
C64 VDD2.t0 B 0.046319f
C65 VDD2.n46 B 0.112154f
C66 VDD2.n47 B 0.57467f
C67 VDD2.n48 B 0.011747f
C68 VDD2.n49 B 0.012438f
C69 VDD2.n50 B 0.027765f
C70 VDD2.n51 B 0.027765f
C71 VDD2.n52 B 0.012438f
C72 VDD2.n53 B 0.011747f
C73 VDD2.n54 B 0.02186f
C74 VDD2.n55 B 0.02186f
C75 VDD2.n56 B 0.011747f
C76 VDD2.n57 B 0.012438f
C77 VDD2.n58 B 0.027765f
C78 VDD2.n59 B 0.027765f
C79 VDD2.n60 B 0.012438f
C80 VDD2.n61 B 0.011747f
C81 VDD2.n62 B 0.02186f
C82 VDD2.n63 B 0.056801f
C83 VDD2.n64 B 0.011747f
C84 VDD2.n65 B 0.012438f
C85 VDD2.n66 B 0.057238f
C86 VDD2.n67 B 0.063392f
C87 VDD2.n68 B 2.18789f
C88 VDD2.t3 B 0.113495f
C89 VDD2.t2 B 0.113495f
C90 VDD2.n69 B 0.971989f
C91 VN.n0 B 0.038414f
C92 VN.t1 B 1.39561f
C93 VN.n1 B 0.040031f
C94 VN.n2 B 0.020422f
C95 VN.n3 B 0.038061f
C96 VN.t4 B 1.69284f
C97 VN.n4 B 0.567423f
C98 VN.t0 B 1.39561f
C99 VN.n5 B 0.582988f
C100 VN.n6 B 0.028666f
C101 VN.n7 B 0.267176f
C102 VN.n8 B 0.020422f
C103 VN.n9 B 0.020422f
C104 VN.n10 B 0.038061f
C105 VN.n11 B 0.036235f
C106 VN.n12 B 0.021419f
C107 VN.n13 B 0.020422f
C108 VN.n14 B 0.020422f
C109 VN.n15 B 0.020422f
C110 VN.n16 B 0.038061f
C111 VN.n17 B 0.037685f
C112 VN.n18 B 0.603001f
C113 VN.n19 B 0.06006f
C114 VN.n20 B 0.038414f
C115 VN.t5 B 1.39561f
C116 VN.n21 B 0.040031f
C117 VN.n22 B 0.020422f
C118 VN.n23 B 0.038061f
C119 VN.t3 B 1.69284f
C120 VN.n24 B 0.567423f
C121 VN.t2 B 1.39561f
C122 VN.n25 B 0.582988f
C123 VN.n26 B 0.028666f
C124 VN.n27 B 0.267176f
C125 VN.n28 B 0.020422f
C126 VN.n29 B 0.020422f
C127 VN.n30 B 0.038061f
C128 VN.n31 B 0.036235f
C129 VN.n32 B 0.021419f
C130 VN.n33 B 0.020422f
C131 VN.n34 B 0.020422f
C132 VN.n35 B 0.020422f
C133 VN.n36 B 0.038061f
C134 VN.n37 B 0.037685f
C135 VN.n38 B 0.603001f
C136 VN.n39 B 1.18982f
C137 VDD1.n0 B 0.012581f
C138 VDD1.n1 B 0.02833f
C139 VDD1.n2 B 0.012691f
C140 VDD1.n3 B 0.022305f
C141 VDD1.n4 B 0.011986f
C142 VDD1.n5 B 0.02833f
C143 VDD1.n6 B 0.012691f
C144 VDD1.n7 B 0.022305f
C145 VDD1.n8 B 0.011986f
C146 VDD1.n9 B 0.021247f
C147 VDD1.n10 B 0.020027f
C148 VDD1.t1 B 0.047261f
C149 VDD1.n11 B 0.114435f
C150 VDD1.n12 B 0.586358f
C151 VDD1.n13 B 0.011986f
C152 VDD1.n14 B 0.012691f
C153 VDD1.n15 B 0.02833f
C154 VDD1.n16 B 0.02833f
C155 VDD1.n17 B 0.012691f
C156 VDD1.n18 B 0.011986f
C157 VDD1.n19 B 0.022305f
C158 VDD1.n20 B 0.022305f
C159 VDD1.n21 B 0.011986f
C160 VDD1.n22 B 0.012691f
C161 VDD1.n23 B 0.02833f
C162 VDD1.n24 B 0.02833f
C163 VDD1.n25 B 0.012691f
C164 VDD1.n26 B 0.011986f
C165 VDD1.n27 B 0.022305f
C166 VDD1.n28 B 0.057956f
C167 VDD1.n29 B 0.011986f
C168 VDD1.n30 B 0.012691f
C169 VDD1.n31 B 0.058402f
C170 VDD1.n32 B 0.077199f
C171 VDD1.n33 B 0.012581f
C172 VDD1.n34 B 0.02833f
C173 VDD1.n35 B 0.012691f
C174 VDD1.n36 B 0.022305f
C175 VDD1.n37 B 0.011986f
C176 VDD1.n38 B 0.02833f
C177 VDD1.n39 B 0.012691f
C178 VDD1.n40 B 0.022305f
C179 VDD1.n41 B 0.011986f
C180 VDD1.n42 B 0.021247f
C181 VDD1.n43 B 0.020027f
C182 VDD1.t5 B 0.047261f
C183 VDD1.n44 B 0.114435f
C184 VDD1.n45 B 0.586358f
C185 VDD1.n46 B 0.011986f
C186 VDD1.n47 B 0.012691f
C187 VDD1.n48 B 0.02833f
C188 VDD1.n49 B 0.02833f
C189 VDD1.n50 B 0.012691f
C190 VDD1.n51 B 0.011986f
C191 VDD1.n52 B 0.022305f
C192 VDD1.n53 B 0.022305f
C193 VDD1.n54 B 0.011986f
C194 VDD1.n55 B 0.012691f
C195 VDD1.n56 B 0.02833f
C196 VDD1.n57 B 0.02833f
C197 VDD1.n58 B 0.012691f
C198 VDD1.n59 B 0.011986f
C199 VDD1.n60 B 0.022305f
C200 VDD1.n61 B 0.057956f
C201 VDD1.n62 B 0.011986f
C202 VDD1.n63 B 0.012691f
C203 VDD1.n64 B 0.058402f
C204 VDD1.n65 B 0.076328f
C205 VDD1.t0 B 0.115803f
C206 VDD1.t4 B 0.115803f
C207 VDD1.n66 B 0.991791f
C208 VDD1.n67 B 2.72635f
C209 VDD1.t3 B 0.115803f
C210 VDD1.t2 B 0.115803f
C211 VDD1.n68 B 0.9856f
C212 VDD1.n69 B 2.43684f
C213 VTAIL.t4 B 0.146054f
C214 VTAIL.t2 B 0.146054f
C215 VTAIL.n0 B 1.17583f
C216 VTAIL.n1 B 0.5436f
C217 VTAIL.n2 B 0.015867f
C218 VTAIL.n3 B 0.03573f
C219 VTAIL.n4 B 0.016006f
C220 VTAIL.n5 B 0.028131f
C221 VTAIL.n6 B 0.015117f
C222 VTAIL.n7 B 0.03573f
C223 VTAIL.n8 B 0.016006f
C224 VTAIL.n9 B 0.028131f
C225 VTAIL.n10 B 0.015117f
C226 VTAIL.n11 B 0.026798f
C227 VTAIL.n12 B 0.025258f
C228 VTAIL.t11 B 0.059607f
C229 VTAIL.n13 B 0.144327f
C230 VTAIL.n14 B 0.739527f
C231 VTAIL.n15 B 0.015117f
C232 VTAIL.n16 B 0.016006f
C233 VTAIL.n17 B 0.03573f
C234 VTAIL.n18 B 0.03573f
C235 VTAIL.n19 B 0.016006f
C236 VTAIL.n20 B 0.015117f
C237 VTAIL.n21 B 0.028131f
C238 VTAIL.n22 B 0.028131f
C239 VTAIL.n23 B 0.015117f
C240 VTAIL.n24 B 0.016006f
C241 VTAIL.n25 B 0.03573f
C242 VTAIL.n26 B 0.03573f
C243 VTAIL.n27 B 0.016006f
C244 VTAIL.n28 B 0.015117f
C245 VTAIL.n29 B 0.028131f
C246 VTAIL.n30 B 0.073095f
C247 VTAIL.n31 B 0.015117f
C248 VTAIL.n32 B 0.016006f
C249 VTAIL.n33 B 0.073658f
C250 VTAIL.n34 B 0.062204f
C251 VTAIL.n35 B 0.567736f
C252 VTAIL.t7 B 0.146054f
C253 VTAIL.t10 B 0.146054f
C254 VTAIL.n36 B 1.17583f
C255 VTAIL.n37 B 2.13676f
C256 VTAIL.t1 B 0.146054f
C257 VTAIL.t5 B 0.146054f
C258 VTAIL.n38 B 1.17582f
C259 VTAIL.n39 B 2.13676f
C260 VTAIL.n40 B 0.015867f
C261 VTAIL.n41 B 0.03573f
C262 VTAIL.n42 B 0.016006f
C263 VTAIL.n43 B 0.028131f
C264 VTAIL.n44 B 0.015117f
C265 VTAIL.n45 B 0.03573f
C266 VTAIL.n46 B 0.016006f
C267 VTAIL.n47 B 0.028131f
C268 VTAIL.n48 B 0.015117f
C269 VTAIL.n49 B 0.026798f
C270 VTAIL.n50 B 0.025258f
C271 VTAIL.t0 B 0.059607f
C272 VTAIL.n51 B 0.144327f
C273 VTAIL.n52 B 0.739527f
C274 VTAIL.n53 B 0.015117f
C275 VTAIL.n54 B 0.016006f
C276 VTAIL.n55 B 0.03573f
C277 VTAIL.n56 B 0.03573f
C278 VTAIL.n57 B 0.016006f
C279 VTAIL.n58 B 0.015117f
C280 VTAIL.n59 B 0.028131f
C281 VTAIL.n60 B 0.028131f
C282 VTAIL.n61 B 0.015117f
C283 VTAIL.n62 B 0.016006f
C284 VTAIL.n63 B 0.03573f
C285 VTAIL.n64 B 0.03573f
C286 VTAIL.n65 B 0.016006f
C287 VTAIL.n66 B 0.015117f
C288 VTAIL.n67 B 0.028131f
C289 VTAIL.n68 B 0.073095f
C290 VTAIL.n69 B 0.015117f
C291 VTAIL.n70 B 0.016006f
C292 VTAIL.n71 B 0.073658f
C293 VTAIL.n72 B 0.062204f
C294 VTAIL.n73 B 0.567736f
C295 VTAIL.t8 B 0.146054f
C296 VTAIL.t9 B 0.146054f
C297 VTAIL.n74 B 1.17582f
C298 VTAIL.n75 B 0.786822f
C299 VTAIL.n76 B 0.015867f
C300 VTAIL.n77 B 0.03573f
C301 VTAIL.n78 B 0.016006f
C302 VTAIL.n79 B 0.028131f
C303 VTAIL.n80 B 0.015117f
C304 VTAIL.n81 B 0.03573f
C305 VTAIL.n82 B 0.016006f
C306 VTAIL.n83 B 0.028131f
C307 VTAIL.n84 B 0.015117f
C308 VTAIL.n85 B 0.026798f
C309 VTAIL.n86 B 0.025258f
C310 VTAIL.t6 B 0.059607f
C311 VTAIL.n87 B 0.144327f
C312 VTAIL.n88 B 0.739527f
C313 VTAIL.n89 B 0.015117f
C314 VTAIL.n90 B 0.016006f
C315 VTAIL.n91 B 0.03573f
C316 VTAIL.n92 B 0.03573f
C317 VTAIL.n93 B 0.016006f
C318 VTAIL.n94 B 0.015117f
C319 VTAIL.n95 B 0.028131f
C320 VTAIL.n96 B 0.028131f
C321 VTAIL.n97 B 0.015117f
C322 VTAIL.n98 B 0.016006f
C323 VTAIL.n99 B 0.03573f
C324 VTAIL.n100 B 0.03573f
C325 VTAIL.n101 B 0.016006f
C326 VTAIL.n102 B 0.015117f
C327 VTAIL.n103 B 0.028131f
C328 VTAIL.n104 B 0.073095f
C329 VTAIL.n105 B 0.015117f
C330 VTAIL.n106 B 0.016006f
C331 VTAIL.n107 B 0.073658f
C332 VTAIL.n108 B 0.062204f
C333 VTAIL.n109 B 1.58635f
C334 VTAIL.n110 B 0.015867f
C335 VTAIL.n111 B 0.03573f
C336 VTAIL.n112 B 0.016006f
C337 VTAIL.n113 B 0.028131f
C338 VTAIL.n114 B 0.015117f
C339 VTAIL.n115 B 0.03573f
C340 VTAIL.n116 B 0.016006f
C341 VTAIL.n117 B 0.028131f
C342 VTAIL.n118 B 0.015117f
C343 VTAIL.n119 B 0.026798f
C344 VTAIL.n120 B 0.025258f
C345 VTAIL.t3 B 0.059607f
C346 VTAIL.n121 B 0.144327f
C347 VTAIL.n122 B 0.739527f
C348 VTAIL.n123 B 0.015117f
C349 VTAIL.n124 B 0.016006f
C350 VTAIL.n125 B 0.03573f
C351 VTAIL.n126 B 0.03573f
C352 VTAIL.n127 B 0.016006f
C353 VTAIL.n128 B 0.015117f
C354 VTAIL.n129 B 0.028131f
C355 VTAIL.n130 B 0.028131f
C356 VTAIL.n131 B 0.015117f
C357 VTAIL.n132 B 0.016006f
C358 VTAIL.n133 B 0.03573f
C359 VTAIL.n134 B 0.03573f
C360 VTAIL.n135 B 0.016006f
C361 VTAIL.n136 B 0.015117f
C362 VTAIL.n137 B 0.028131f
C363 VTAIL.n138 B 0.073095f
C364 VTAIL.n139 B 0.015117f
C365 VTAIL.n140 B 0.016006f
C366 VTAIL.n141 B 0.073658f
C367 VTAIL.n142 B 0.062204f
C368 VTAIL.n143 B 1.49824f
C369 VP.n0 B 0.039662f
C370 VP.t1 B 1.44096f
C371 VP.n1 B 0.041332f
C372 VP.n2 B 0.021085f
C373 VP.n3 B 0.039298f
C374 VP.n4 B 0.021085f
C375 VP.t5 B 1.44096f
C376 VP.n5 B 0.039298f
C377 VP.n6 B 0.021085f
C378 VP.n7 B 0.039298f
C379 VP.n8 B 0.039662f
C380 VP.t3 B 1.44096f
C381 VP.n9 B 0.041332f
C382 VP.n10 B 0.021085f
C383 VP.n11 B 0.039298f
C384 VP.t4 B 1.74785f
C385 VP.n12 B 0.585862f
C386 VP.t2 B 1.44096f
C387 VP.n13 B 0.601932f
C388 VP.n14 B 0.029597f
C389 VP.n15 B 0.275858f
C390 VP.n16 B 0.021085f
C391 VP.n17 B 0.021085f
C392 VP.n18 B 0.039298f
C393 VP.n19 B 0.037412f
C394 VP.n20 B 0.022115f
C395 VP.n21 B 0.021085f
C396 VP.n22 B 0.021085f
C397 VP.n23 B 0.021085f
C398 VP.n24 B 0.039298f
C399 VP.n25 B 0.03891f
C400 VP.n26 B 0.622594f
C401 VP.n27 B 1.22297f
C402 VP.n28 B 1.23813f
C403 VP.t0 B 1.44096f
C404 VP.n29 B 0.622594f
C405 VP.n30 B 0.03891f
C406 VP.n31 B 0.039662f
C407 VP.n32 B 0.021085f
C408 VP.n33 B 0.021085f
C409 VP.n34 B 0.041332f
C410 VP.n35 B 0.022115f
C411 VP.n36 B 0.037412f
C412 VP.n37 B 0.021085f
C413 VP.n38 B 0.021085f
C414 VP.n39 B 0.021085f
C415 VP.n40 B 0.039298f
C416 VP.n41 B 0.029597f
C417 VP.n42 B 0.525393f
C418 VP.n43 B 0.029597f
C419 VP.n44 B 0.021085f
C420 VP.n45 B 0.021085f
C421 VP.n46 B 0.021085f
C422 VP.n47 B 0.039298f
C423 VP.n48 B 0.037412f
C424 VP.n49 B 0.022115f
C425 VP.n50 B 0.021085f
C426 VP.n51 B 0.021085f
C427 VP.n52 B 0.021085f
C428 VP.n53 B 0.039298f
C429 VP.n54 B 0.03891f
C430 VP.n55 B 0.622594f
C431 VP.n56 B 0.062012f
.ends

