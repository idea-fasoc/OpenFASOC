* NGSPICE file created from diff_pair_sample_1039.ext - technology: sky130A

.subckt diff_pair_sample_1039 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t3 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=2.74725 pd=16.98 as=2.74725 ps=16.98 w=16.65 l=1.35
X1 VDD2.t9 VN.t0 VTAIL.t9 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=2.74725 pd=16.98 as=6.4935 ps=34.08 w=16.65 l=1.35
X2 VDD1.t2 VP.t1 VTAIL.t18 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=6.4935 pd=34.08 as=2.74725 ps=16.98 w=16.65 l=1.35
X3 VTAIL.t8 VN.t1 VDD2.t8 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=2.74725 pd=16.98 as=2.74725 ps=16.98 w=16.65 l=1.35
X4 B.t11 B.t9 B.t10 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=6.4935 pd=34.08 as=0 ps=0 w=16.65 l=1.35
X5 VDD1.t5 VP.t2 VTAIL.t17 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=6.4935 pd=34.08 as=2.74725 ps=16.98 w=16.65 l=1.35
X6 VDD1.t4 VP.t3 VTAIL.t16 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=2.74725 pd=16.98 as=2.74725 ps=16.98 w=16.65 l=1.35
X7 VDD2.t7 VN.t2 VTAIL.t2 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=6.4935 pd=34.08 as=2.74725 ps=16.98 w=16.65 l=1.35
X8 B.t8 B.t6 B.t7 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=6.4935 pd=34.08 as=0 ps=0 w=16.65 l=1.35
X9 VDD2.t6 VN.t3 VTAIL.t7 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=2.74725 pd=16.98 as=6.4935 ps=34.08 w=16.65 l=1.35
X10 VDD2.t5 VN.t4 VTAIL.t1 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=2.74725 pd=16.98 as=2.74725 ps=16.98 w=16.65 l=1.35
X11 B.t5 B.t3 B.t4 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=6.4935 pd=34.08 as=0 ps=0 w=16.65 l=1.35
X12 VDD2.t4 VN.t5 VTAIL.t5 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=6.4935 pd=34.08 as=2.74725 ps=16.98 w=16.65 l=1.35
X13 VTAIL.t15 VP.t4 VDD1.t7 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=2.74725 pd=16.98 as=2.74725 ps=16.98 w=16.65 l=1.35
X14 VTAIL.t14 VP.t5 VDD1.t6 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=2.74725 pd=16.98 as=2.74725 ps=16.98 w=16.65 l=1.35
X15 VDD2.t3 VN.t6 VTAIL.t4 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=2.74725 pd=16.98 as=2.74725 ps=16.98 w=16.65 l=1.35
X16 VTAIL.t0 VN.t7 VDD2.t2 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=2.74725 pd=16.98 as=2.74725 ps=16.98 w=16.65 l=1.35
X17 VDD1.t9 VP.t6 VTAIL.t13 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=2.74725 pd=16.98 as=6.4935 ps=34.08 w=16.65 l=1.35
X18 VTAIL.t3 VN.t8 VDD2.t1 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=2.74725 pd=16.98 as=2.74725 ps=16.98 w=16.65 l=1.35
X19 B.t2 B.t0 B.t1 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=6.4935 pd=34.08 as=0 ps=0 w=16.65 l=1.35
X20 VDD1.t8 VP.t7 VTAIL.t12 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=2.74725 pd=16.98 as=2.74725 ps=16.98 w=16.65 l=1.35
X21 VDD1.t1 VP.t8 VTAIL.t11 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=2.74725 pd=16.98 as=6.4935 ps=34.08 w=16.65 l=1.35
X22 VTAIL.t6 VN.t9 VDD2.t0 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=2.74725 pd=16.98 as=2.74725 ps=16.98 w=16.65 l=1.35
X23 VTAIL.t10 VP.t9 VDD1.t0 w_n2986_n4298# sky130_fd_pr__pfet_01v8 ad=2.74725 pd=16.98 as=2.74725 ps=16.98 w=16.65 l=1.35
R0 VP.n13 VP.t1 344.692
R1 VP.n31 VP.t2 326.51
R2 VP.n49 VP.t6 326.51
R3 VP.n28 VP.t8 326.51
R4 VP.n3 VP.t3 297.233
R5 VP.n5 VP.t0 297.233
R6 VP.n1 VP.t9 297.233
R7 VP.n10 VP.t7 297.233
R8 VP.n8 VP.t4 297.233
R9 VP.n12 VP.t5 297.233
R10 VP.n15 VP.n14 161.3
R11 VP.n16 VP.n11 161.3
R12 VP.n18 VP.n17 161.3
R13 VP.n19 VP.n10 161.3
R14 VP.n21 VP.n20 161.3
R15 VP.n22 VP.n9 161.3
R16 VP.n24 VP.n23 161.3
R17 VP.n26 VP.n25 161.3
R18 VP.n27 VP.n7 161.3
R19 VP.n48 VP.n0 161.3
R20 VP.n47 VP.n46 161.3
R21 VP.n45 VP.n44 161.3
R22 VP.n43 VP.n2 161.3
R23 VP.n42 VP.n41 161.3
R24 VP.n40 VP.n3 161.3
R25 VP.n39 VP.n38 161.3
R26 VP.n37 VP.n4 161.3
R27 VP.n36 VP.n35 161.3
R28 VP.n34 VP.n33 161.3
R29 VP.n32 VP.n6 161.3
R30 VP.n29 VP.n28 80.6037
R31 VP.n50 VP.n49 80.6037
R32 VP.n31 VP.n30 80.6037
R33 VP.n38 VP.n37 56.0336
R34 VP.n43 VP.n42 56.0336
R35 VP.n22 VP.n21 56.0336
R36 VP.n17 VP.n16 56.0336
R37 VP.n30 VP.n29 50.0393
R38 VP.n13 VP.n12 49.0179
R39 VP.n33 VP.n32 38.5509
R40 VP.n48 VP.n47 38.5509
R41 VP.n27 VP.n26 38.5509
R42 VP.n14 VP.n13 29.8396
R43 VP.n32 VP.n31 27.0217
R44 VP.n49 VP.n48 27.0217
R45 VP.n28 VP.n27 27.0217
R46 VP.n37 VP.n36 24.9531
R47 VP.n44 VP.n43 24.9531
R48 VP.n23 VP.n22 24.9531
R49 VP.n16 VP.n15 24.9531
R50 VP.n38 VP.n3 24.4675
R51 VP.n42 VP.n3 24.4675
R52 VP.n17 VP.n10 24.4675
R53 VP.n21 VP.n10 24.4675
R54 VP.n33 VP.n5 15.6594
R55 VP.n47 VP.n1 15.6594
R56 VP.n26 VP.n8 15.6594
R57 VP.n36 VP.n5 8.80862
R58 VP.n44 VP.n1 8.80862
R59 VP.n23 VP.n8 8.80862
R60 VP.n15 VP.n12 8.80862
R61 VP.n29 VP.n7 0.285035
R62 VP.n30 VP.n6 0.285035
R63 VP.n50 VP.n0 0.285035
R64 VP.n14 VP.n11 0.189894
R65 VP.n18 VP.n11 0.189894
R66 VP.n19 VP.n18 0.189894
R67 VP.n20 VP.n19 0.189894
R68 VP.n20 VP.n9 0.189894
R69 VP.n24 VP.n9 0.189894
R70 VP.n25 VP.n24 0.189894
R71 VP.n25 VP.n7 0.189894
R72 VP.n34 VP.n6 0.189894
R73 VP.n35 VP.n34 0.189894
R74 VP.n35 VP.n4 0.189894
R75 VP.n39 VP.n4 0.189894
R76 VP.n40 VP.n39 0.189894
R77 VP.n41 VP.n40 0.189894
R78 VP.n41 VP.n2 0.189894
R79 VP.n45 VP.n2 0.189894
R80 VP.n46 VP.n45 0.189894
R81 VP.n46 VP.n0 0.189894
R82 VP VP.n50 0.146778
R83 VDD1.n1 VDD1.t2 77.0647
R84 VDD1.n3 VDD1.t5 77.0645
R85 VDD1.n5 VDD1.n4 74.6948
R86 VDD1.n1 VDD1.n0 73.6642
R87 VDD1.n7 VDD1.n6 73.664
R88 VDD1.n3 VDD1.n2 73.6639
R89 VDD1.n7 VDD1.n5 46.2552
R90 VDD1.n6 VDD1.t7 1.95275
R91 VDD1.n6 VDD1.t1 1.95275
R92 VDD1.n0 VDD1.t6 1.95275
R93 VDD1.n0 VDD1.t8 1.95275
R94 VDD1.n4 VDD1.t0 1.95275
R95 VDD1.n4 VDD1.t9 1.95275
R96 VDD1.n2 VDD1.t3 1.95275
R97 VDD1.n2 VDD1.t4 1.95275
R98 VDD1 VDD1.n7 1.02852
R99 VDD1 VDD1.n1 0.420759
R100 VDD1.n5 VDD1.n3 0.307223
R101 VTAIL.n11 VTAIL.t7 58.9377
R102 VTAIL.n17 VTAIL.t9 58.9374
R103 VTAIL.n2 VTAIL.t13 58.9374
R104 VTAIL.n16 VTAIL.t11 58.9374
R105 VTAIL.n15 VTAIL.n14 56.9854
R106 VTAIL.n13 VTAIL.n12 56.9854
R107 VTAIL.n10 VTAIL.n9 56.9854
R108 VTAIL.n8 VTAIL.n7 56.9854
R109 VTAIL.n19 VTAIL.n18 56.9852
R110 VTAIL.n1 VTAIL.n0 56.9852
R111 VTAIL.n4 VTAIL.n3 56.9852
R112 VTAIL.n6 VTAIL.n5 56.9852
R113 VTAIL.n8 VTAIL.n6 29.6169
R114 VTAIL.n17 VTAIL.n16 28.1686
R115 VTAIL.n18 VTAIL.t4 1.95275
R116 VTAIL.n18 VTAIL.t8 1.95275
R117 VTAIL.n0 VTAIL.t5 1.95275
R118 VTAIL.n0 VTAIL.t0 1.95275
R119 VTAIL.n3 VTAIL.t16 1.95275
R120 VTAIL.n3 VTAIL.t10 1.95275
R121 VTAIL.n5 VTAIL.t17 1.95275
R122 VTAIL.n5 VTAIL.t19 1.95275
R123 VTAIL.n14 VTAIL.t12 1.95275
R124 VTAIL.n14 VTAIL.t15 1.95275
R125 VTAIL.n12 VTAIL.t18 1.95275
R126 VTAIL.n12 VTAIL.t14 1.95275
R127 VTAIL.n9 VTAIL.t1 1.95275
R128 VTAIL.n9 VTAIL.t3 1.95275
R129 VTAIL.n7 VTAIL.t2 1.95275
R130 VTAIL.n7 VTAIL.t6 1.95275
R131 VTAIL.n10 VTAIL.n8 1.44878
R132 VTAIL.n11 VTAIL.n10 1.44878
R133 VTAIL.n15 VTAIL.n13 1.44878
R134 VTAIL.n16 VTAIL.n15 1.44878
R135 VTAIL.n6 VTAIL.n4 1.44878
R136 VTAIL.n4 VTAIL.n2 1.44878
R137 VTAIL.n19 VTAIL.n17 1.44878
R138 VTAIL.n13 VTAIL.n11 1.19447
R139 VTAIL.n2 VTAIL.n1 1.19447
R140 VTAIL VTAIL.n1 1.1449
R141 VTAIL VTAIL.n19 0.304379
R142 VN.n6 VN.t5 344.692
R143 VN.n29 VN.t3 344.692
R144 VN.n21 VN.t0 326.51
R145 VN.n44 VN.t2 326.51
R146 VN.n3 VN.t6 297.233
R147 VN.n5 VN.t7 297.233
R148 VN.n1 VN.t1 297.233
R149 VN.n26 VN.t4 297.233
R150 VN.n28 VN.t8 297.233
R151 VN.n24 VN.t9 297.233
R152 VN.n43 VN.n23 161.3
R153 VN.n42 VN.n41 161.3
R154 VN.n40 VN.n39 161.3
R155 VN.n38 VN.n25 161.3
R156 VN.n37 VN.n36 161.3
R157 VN.n35 VN.n26 161.3
R158 VN.n34 VN.n33 161.3
R159 VN.n32 VN.n27 161.3
R160 VN.n31 VN.n30 161.3
R161 VN.n20 VN.n0 161.3
R162 VN.n19 VN.n18 161.3
R163 VN.n17 VN.n16 161.3
R164 VN.n15 VN.n2 161.3
R165 VN.n14 VN.n13 161.3
R166 VN.n12 VN.n3 161.3
R167 VN.n11 VN.n10 161.3
R168 VN.n9 VN.n4 161.3
R169 VN.n8 VN.n7 161.3
R170 VN.n45 VN.n44 80.6037
R171 VN.n22 VN.n21 80.6037
R172 VN.n10 VN.n9 56.0336
R173 VN.n15 VN.n14 56.0336
R174 VN.n33 VN.n32 56.0336
R175 VN.n38 VN.n37 56.0336
R176 VN VN.n45 50.3248
R177 VN.n6 VN.n5 49.0179
R178 VN.n29 VN.n28 49.0179
R179 VN.n20 VN.n19 38.5509
R180 VN.n43 VN.n42 38.5509
R181 VN.n30 VN.n29 29.8396
R182 VN.n7 VN.n6 29.8396
R183 VN.n21 VN.n20 27.0217
R184 VN.n44 VN.n43 27.0217
R185 VN.n9 VN.n8 24.9531
R186 VN.n16 VN.n15 24.9531
R187 VN.n32 VN.n31 24.9531
R188 VN.n39 VN.n38 24.9531
R189 VN.n10 VN.n3 24.4675
R190 VN.n14 VN.n3 24.4675
R191 VN.n37 VN.n26 24.4675
R192 VN.n33 VN.n26 24.4675
R193 VN.n19 VN.n1 15.6594
R194 VN.n42 VN.n24 15.6594
R195 VN.n8 VN.n5 8.80862
R196 VN.n16 VN.n1 8.80862
R197 VN.n31 VN.n28 8.80862
R198 VN.n39 VN.n24 8.80862
R199 VN.n45 VN.n23 0.285035
R200 VN.n22 VN.n0 0.285035
R201 VN.n41 VN.n23 0.189894
R202 VN.n41 VN.n40 0.189894
R203 VN.n40 VN.n25 0.189894
R204 VN.n36 VN.n25 0.189894
R205 VN.n36 VN.n35 0.189894
R206 VN.n35 VN.n34 0.189894
R207 VN.n34 VN.n27 0.189894
R208 VN.n30 VN.n27 0.189894
R209 VN.n7 VN.n4 0.189894
R210 VN.n11 VN.n4 0.189894
R211 VN.n12 VN.n11 0.189894
R212 VN.n13 VN.n12 0.189894
R213 VN.n13 VN.n2 0.189894
R214 VN.n17 VN.n2 0.189894
R215 VN.n18 VN.n17 0.189894
R216 VN.n18 VN.n0 0.189894
R217 VN VN.n22 0.146778
R218 VDD2.n1 VDD2.t4 77.0645
R219 VDD2.n4 VDD2.t7 75.6165
R220 VDD2.n3 VDD2.n2 74.6948
R221 VDD2 VDD2.n7 74.692
R222 VDD2.n6 VDD2.n5 73.6642
R223 VDD2.n1 VDD2.n0 73.6639
R224 VDD2.n4 VDD2.n3 44.948
R225 VDD2.n7 VDD2.t1 1.95275
R226 VDD2.n7 VDD2.t6 1.95275
R227 VDD2.n5 VDD2.t0 1.95275
R228 VDD2.n5 VDD2.t5 1.95275
R229 VDD2.n2 VDD2.t8 1.95275
R230 VDD2.n2 VDD2.t9 1.95275
R231 VDD2.n0 VDD2.t2 1.95275
R232 VDD2.n0 VDD2.t3 1.95275
R233 VDD2.n6 VDD2.n4 1.44878
R234 VDD2 VDD2.n6 0.420759
R235 VDD2.n3 VDD2.n1 0.307223
R236 B.n440 B.n123 585
R237 B.n439 B.n438 585
R238 B.n437 B.n124 585
R239 B.n436 B.n435 585
R240 B.n434 B.n125 585
R241 B.n433 B.n432 585
R242 B.n431 B.n126 585
R243 B.n430 B.n429 585
R244 B.n428 B.n127 585
R245 B.n427 B.n426 585
R246 B.n425 B.n128 585
R247 B.n424 B.n423 585
R248 B.n422 B.n129 585
R249 B.n421 B.n420 585
R250 B.n419 B.n130 585
R251 B.n418 B.n417 585
R252 B.n416 B.n131 585
R253 B.n415 B.n414 585
R254 B.n413 B.n132 585
R255 B.n412 B.n411 585
R256 B.n410 B.n133 585
R257 B.n409 B.n408 585
R258 B.n407 B.n134 585
R259 B.n406 B.n405 585
R260 B.n404 B.n135 585
R261 B.n403 B.n402 585
R262 B.n401 B.n136 585
R263 B.n400 B.n399 585
R264 B.n398 B.n137 585
R265 B.n397 B.n396 585
R266 B.n395 B.n138 585
R267 B.n394 B.n393 585
R268 B.n392 B.n139 585
R269 B.n391 B.n390 585
R270 B.n389 B.n140 585
R271 B.n388 B.n387 585
R272 B.n386 B.n141 585
R273 B.n385 B.n384 585
R274 B.n383 B.n142 585
R275 B.n382 B.n381 585
R276 B.n380 B.n143 585
R277 B.n379 B.n378 585
R278 B.n377 B.n144 585
R279 B.n376 B.n375 585
R280 B.n374 B.n145 585
R281 B.n373 B.n372 585
R282 B.n371 B.n146 585
R283 B.n370 B.n369 585
R284 B.n368 B.n147 585
R285 B.n367 B.n366 585
R286 B.n365 B.n148 585
R287 B.n364 B.n363 585
R288 B.n362 B.n149 585
R289 B.n361 B.n360 585
R290 B.n359 B.n150 585
R291 B.n358 B.n357 585
R292 B.n353 B.n151 585
R293 B.n352 B.n351 585
R294 B.n350 B.n152 585
R295 B.n349 B.n348 585
R296 B.n347 B.n153 585
R297 B.n346 B.n345 585
R298 B.n344 B.n154 585
R299 B.n343 B.n342 585
R300 B.n341 B.n155 585
R301 B.n339 B.n338 585
R302 B.n337 B.n158 585
R303 B.n336 B.n335 585
R304 B.n334 B.n159 585
R305 B.n333 B.n332 585
R306 B.n331 B.n160 585
R307 B.n330 B.n329 585
R308 B.n328 B.n161 585
R309 B.n327 B.n326 585
R310 B.n325 B.n162 585
R311 B.n324 B.n323 585
R312 B.n322 B.n163 585
R313 B.n321 B.n320 585
R314 B.n319 B.n164 585
R315 B.n318 B.n317 585
R316 B.n316 B.n165 585
R317 B.n315 B.n314 585
R318 B.n313 B.n166 585
R319 B.n312 B.n311 585
R320 B.n310 B.n167 585
R321 B.n309 B.n308 585
R322 B.n307 B.n168 585
R323 B.n306 B.n305 585
R324 B.n304 B.n169 585
R325 B.n303 B.n302 585
R326 B.n301 B.n170 585
R327 B.n300 B.n299 585
R328 B.n298 B.n171 585
R329 B.n297 B.n296 585
R330 B.n295 B.n172 585
R331 B.n294 B.n293 585
R332 B.n292 B.n173 585
R333 B.n291 B.n290 585
R334 B.n289 B.n174 585
R335 B.n288 B.n287 585
R336 B.n286 B.n175 585
R337 B.n285 B.n284 585
R338 B.n283 B.n176 585
R339 B.n282 B.n281 585
R340 B.n280 B.n177 585
R341 B.n279 B.n278 585
R342 B.n277 B.n178 585
R343 B.n276 B.n275 585
R344 B.n274 B.n179 585
R345 B.n273 B.n272 585
R346 B.n271 B.n180 585
R347 B.n270 B.n269 585
R348 B.n268 B.n181 585
R349 B.n267 B.n266 585
R350 B.n265 B.n182 585
R351 B.n264 B.n263 585
R352 B.n262 B.n183 585
R353 B.n261 B.n260 585
R354 B.n259 B.n184 585
R355 B.n258 B.n257 585
R356 B.n442 B.n441 585
R357 B.n443 B.n122 585
R358 B.n445 B.n444 585
R359 B.n446 B.n121 585
R360 B.n448 B.n447 585
R361 B.n449 B.n120 585
R362 B.n451 B.n450 585
R363 B.n452 B.n119 585
R364 B.n454 B.n453 585
R365 B.n455 B.n118 585
R366 B.n457 B.n456 585
R367 B.n458 B.n117 585
R368 B.n460 B.n459 585
R369 B.n461 B.n116 585
R370 B.n463 B.n462 585
R371 B.n464 B.n115 585
R372 B.n466 B.n465 585
R373 B.n467 B.n114 585
R374 B.n469 B.n468 585
R375 B.n470 B.n113 585
R376 B.n472 B.n471 585
R377 B.n473 B.n112 585
R378 B.n475 B.n474 585
R379 B.n476 B.n111 585
R380 B.n478 B.n477 585
R381 B.n479 B.n110 585
R382 B.n481 B.n480 585
R383 B.n482 B.n109 585
R384 B.n484 B.n483 585
R385 B.n485 B.n108 585
R386 B.n487 B.n486 585
R387 B.n488 B.n107 585
R388 B.n490 B.n489 585
R389 B.n491 B.n106 585
R390 B.n493 B.n492 585
R391 B.n494 B.n105 585
R392 B.n496 B.n495 585
R393 B.n497 B.n104 585
R394 B.n499 B.n498 585
R395 B.n500 B.n103 585
R396 B.n502 B.n501 585
R397 B.n503 B.n102 585
R398 B.n505 B.n504 585
R399 B.n506 B.n101 585
R400 B.n508 B.n507 585
R401 B.n509 B.n100 585
R402 B.n511 B.n510 585
R403 B.n512 B.n99 585
R404 B.n514 B.n513 585
R405 B.n515 B.n98 585
R406 B.n517 B.n516 585
R407 B.n518 B.n97 585
R408 B.n520 B.n519 585
R409 B.n521 B.n96 585
R410 B.n523 B.n522 585
R411 B.n524 B.n95 585
R412 B.n526 B.n525 585
R413 B.n527 B.n94 585
R414 B.n529 B.n528 585
R415 B.n530 B.n93 585
R416 B.n532 B.n531 585
R417 B.n533 B.n92 585
R418 B.n535 B.n534 585
R419 B.n536 B.n91 585
R420 B.n538 B.n537 585
R421 B.n539 B.n90 585
R422 B.n541 B.n540 585
R423 B.n542 B.n89 585
R424 B.n544 B.n543 585
R425 B.n545 B.n88 585
R426 B.n547 B.n546 585
R427 B.n548 B.n87 585
R428 B.n550 B.n549 585
R429 B.n551 B.n86 585
R430 B.n553 B.n552 585
R431 B.n554 B.n85 585
R432 B.n736 B.n735 585
R433 B.n734 B.n21 585
R434 B.n733 B.n732 585
R435 B.n731 B.n22 585
R436 B.n730 B.n729 585
R437 B.n728 B.n23 585
R438 B.n727 B.n726 585
R439 B.n725 B.n24 585
R440 B.n724 B.n723 585
R441 B.n722 B.n25 585
R442 B.n721 B.n720 585
R443 B.n719 B.n26 585
R444 B.n718 B.n717 585
R445 B.n716 B.n27 585
R446 B.n715 B.n714 585
R447 B.n713 B.n28 585
R448 B.n712 B.n711 585
R449 B.n710 B.n29 585
R450 B.n709 B.n708 585
R451 B.n707 B.n30 585
R452 B.n706 B.n705 585
R453 B.n704 B.n31 585
R454 B.n703 B.n702 585
R455 B.n701 B.n32 585
R456 B.n700 B.n699 585
R457 B.n698 B.n33 585
R458 B.n697 B.n696 585
R459 B.n695 B.n34 585
R460 B.n694 B.n693 585
R461 B.n692 B.n35 585
R462 B.n691 B.n690 585
R463 B.n689 B.n36 585
R464 B.n688 B.n687 585
R465 B.n686 B.n37 585
R466 B.n685 B.n684 585
R467 B.n683 B.n38 585
R468 B.n682 B.n681 585
R469 B.n680 B.n39 585
R470 B.n679 B.n678 585
R471 B.n677 B.n40 585
R472 B.n676 B.n675 585
R473 B.n674 B.n41 585
R474 B.n673 B.n672 585
R475 B.n671 B.n42 585
R476 B.n670 B.n669 585
R477 B.n668 B.n43 585
R478 B.n667 B.n666 585
R479 B.n665 B.n44 585
R480 B.n664 B.n663 585
R481 B.n662 B.n45 585
R482 B.n661 B.n660 585
R483 B.n659 B.n46 585
R484 B.n658 B.n657 585
R485 B.n656 B.n47 585
R486 B.n655 B.n654 585
R487 B.n653 B.n652 585
R488 B.n651 B.n51 585
R489 B.n650 B.n649 585
R490 B.n648 B.n52 585
R491 B.n647 B.n646 585
R492 B.n645 B.n53 585
R493 B.n644 B.n643 585
R494 B.n642 B.n54 585
R495 B.n641 B.n640 585
R496 B.n639 B.n55 585
R497 B.n637 B.n636 585
R498 B.n635 B.n58 585
R499 B.n634 B.n633 585
R500 B.n632 B.n59 585
R501 B.n631 B.n630 585
R502 B.n629 B.n60 585
R503 B.n628 B.n627 585
R504 B.n626 B.n61 585
R505 B.n625 B.n624 585
R506 B.n623 B.n62 585
R507 B.n622 B.n621 585
R508 B.n620 B.n63 585
R509 B.n619 B.n618 585
R510 B.n617 B.n64 585
R511 B.n616 B.n615 585
R512 B.n614 B.n65 585
R513 B.n613 B.n612 585
R514 B.n611 B.n66 585
R515 B.n610 B.n609 585
R516 B.n608 B.n67 585
R517 B.n607 B.n606 585
R518 B.n605 B.n68 585
R519 B.n604 B.n603 585
R520 B.n602 B.n69 585
R521 B.n601 B.n600 585
R522 B.n599 B.n70 585
R523 B.n598 B.n597 585
R524 B.n596 B.n71 585
R525 B.n595 B.n594 585
R526 B.n593 B.n72 585
R527 B.n592 B.n591 585
R528 B.n590 B.n73 585
R529 B.n589 B.n588 585
R530 B.n587 B.n74 585
R531 B.n586 B.n585 585
R532 B.n584 B.n75 585
R533 B.n583 B.n582 585
R534 B.n581 B.n76 585
R535 B.n580 B.n579 585
R536 B.n578 B.n77 585
R537 B.n577 B.n576 585
R538 B.n575 B.n78 585
R539 B.n574 B.n573 585
R540 B.n572 B.n79 585
R541 B.n571 B.n570 585
R542 B.n569 B.n80 585
R543 B.n568 B.n567 585
R544 B.n566 B.n81 585
R545 B.n565 B.n564 585
R546 B.n563 B.n82 585
R547 B.n562 B.n561 585
R548 B.n560 B.n83 585
R549 B.n559 B.n558 585
R550 B.n557 B.n84 585
R551 B.n556 B.n555 585
R552 B.n737 B.n20 585
R553 B.n739 B.n738 585
R554 B.n740 B.n19 585
R555 B.n742 B.n741 585
R556 B.n743 B.n18 585
R557 B.n745 B.n744 585
R558 B.n746 B.n17 585
R559 B.n748 B.n747 585
R560 B.n749 B.n16 585
R561 B.n751 B.n750 585
R562 B.n752 B.n15 585
R563 B.n754 B.n753 585
R564 B.n755 B.n14 585
R565 B.n757 B.n756 585
R566 B.n758 B.n13 585
R567 B.n760 B.n759 585
R568 B.n761 B.n12 585
R569 B.n763 B.n762 585
R570 B.n764 B.n11 585
R571 B.n766 B.n765 585
R572 B.n767 B.n10 585
R573 B.n769 B.n768 585
R574 B.n770 B.n9 585
R575 B.n772 B.n771 585
R576 B.n773 B.n8 585
R577 B.n775 B.n774 585
R578 B.n776 B.n7 585
R579 B.n778 B.n777 585
R580 B.n779 B.n6 585
R581 B.n781 B.n780 585
R582 B.n782 B.n5 585
R583 B.n784 B.n783 585
R584 B.n785 B.n4 585
R585 B.n787 B.n786 585
R586 B.n788 B.n3 585
R587 B.n790 B.n789 585
R588 B.n791 B.n0 585
R589 B.n2 B.n1 585
R590 B.n204 B.n203 585
R591 B.n205 B.n202 585
R592 B.n207 B.n206 585
R593 B.n208 B.n201 585
R594 B.n210 B.n209 585
R595 B.n211 B.n200 585
R596 B.n213 B.n212 585
R597 B.n214 B.n199 585
R598 B.n216 B.n215 585
R599 B.n217 B.n198 585
R600 B.n219 B.n218 585
R601 B.n220 B.n197 585
R602 B.n222 B.n221 585
R603 B.n223 B.n196 585
R604 B.n225 B.n224 585
R605 B.n226 B.n195 585
R606 B.n228 B.n227 585
R607 B.n229 B.n194 585
R608 B.n231 B.n230 585
R609 B.n232 B.n193 585
R610 B.n234 B.n233 585
R611 B.n235 B.n192 585
R612 B.n237 B.n236 585
R613 B.n238 B.n191 585
R614 B.n240 B.n239 585
R615 B.n241 B.n190 585
R616 B.n243 B.n242 585
R617 B.n244 B.n189 585
R618 B.n246 B.n245 585
R619 B.n247 B.n188 585
R620 B.n249 B.n248 585
R621 B.n250 B.n187 585
R622 B.n252 B.n251 585
R623 B.n253 B.n186 585
R624 B.n255 B.n254 585
R625 B.n256 B.n185 585
R626 B.n258 B.n185 554.963
R627 B.n442 B.n123 554.963
R628 B.n556 B.n85 554.963
R629 B.n737 B.n736 554.963
R630 B.n156 B.t0 502.067
R631 B.n354 B.t3 502.067
R632 B.n56 B.t6 502.067
R633 B.n48 B.t9 502.067
R634 B.n793 B.n792 256.663
R635 B.n792 B.n791 235.042
R636 B.n792 B.n2 235.042
R637 B.n259 B.n258 163.367
R638 B.n260 B.n259 163.367
R639 B.n260 B.n183 163.367
R640 B.n264 B.n183 163.367
R641 B.n265 B.n264 163.367
R642 B.n266 B.n265 163.367
R643 B.n266 B.n181 163.367
R644 B.n270 B.n181 163.367
R645 B.n271 B.n270 163.367
R646 B.n272 B.n271 163.367
R647 B.n272 B.n179 163.367
R648 B.n276 B.n179 163.367
R649 B.n277 B.n276 163.367
R650 B.n278 B.n277 163.367
R651 B.n278 B.n177 163.367
R652 B.n282 B.n177 163.367
R653 B.n283 B.n282 163.367
R654 B.n284 B.n283 163.367
R655 B.n284 B.n175 163.367
R656 B.n288 B.n175 163.367
R657 B.n289 B.n288 163.367
R658 B.n290 B.n289 163.367
R659 B.n290 B.n173 163.367
R660 B.n294 B.n173 163.367
R661 B.n295 B.n294 163.367
R662 B.n296 B.n295 163.367
R663 B.n296 B.n171 163.367
R664 B.n300 B.n171 163.367
R665 B.n301 B.n300 163.367
R666 B.n302 B.n301 163.367
R667 B.n302 B.n169 163.367
R668 B.n306 B.n169 163.367
R669 B.n307 B.n306 163.367
R670 B.n308 B.n307 163.367
R671 B.n308 B.n167 163.367
R672 B.n312 B.n167 163.367
R673 B.n313 B.n312 163.367
R674 B.n314 B.n313 163.367
R675 B.n314 B.n165 163.367
R676 B.n318 B.n165 163.367
R677 B.n319 B.n318 163.367
R678 B.n320 B.n319 163.367
R679 B.n320 B.n163 163.367
R680 B.n324 B.n163 163.367
R681 B.n325 B.n324 163.367
R682 B.n326 B.n325 163.367
R683 B.n326 B.n161 163.367
R684 B.n330 B.n161 163.367
R685 B.n331 B.n330 163.367
R686 B.n332 B.n331 163.367
R687 B.n332 B.n159 163.367
R688 B.n336 B.n159 163.367
R689 B.n337 B.n336 163.367
R690 B.n338 B.n337 163.367
R691 B.n338 B.n155 163.367
R692 B.n343 B.n155 163.367
R693 B.n344 B.n343 163.367
R694 B.n345 B.n344 163.367
R695 B.n345 B.n153 163.367
R696 B.n349 B.n153 163.367
R697 B.n350 B.n349 163.367
R698 B.n351 B.n350 163.367
R699 B.n351 B.n151 163.367
R700 B.n358 B.n151 163.367
R701 B.n359 B.n358 163.367
R702 B.n360 B.n359 163.367
R703 B.n360 B.n149 163.367
R704 B.n364 B.n149 163.367
R705 B.n365 B.n364 163.367
R706 B.n366 B.n365 163.367
R707 B.n366 B.n147 163.367
R708 B.n370 B.n147 163.367
R709 B.n371 B.n370 163.367
R710 B.n372 B.n371 163.367
R711 B.n372 B.n145 163.367
R712 B.n376 B.n145 163.367
R713 B.n377 B.n376 163.367
R714 B.n378 B.n377 163.367
R715 B.n378 B.n143 163.367
R716 B.n382 B.n143 163.367
R717 B.n383 B.n382 163.367
R718 B.n384 B.n383 163.367
R719 B.n384 B.n141 163.367
R720 B.n388 B.n141 163.367
R721 B.n389 B.n388 163.367
R722 B.n390 B.n389 163.367
R723 B.n390 B.n139 163.367
R724 B.n394 B.n139 163.367
R725 B.n395 B.n394 163.367
R726 B.n396 B.n395 163.367
R727 B.n396 B.n137 163.367
R728 B.n400 B.n137 163.367
R729 B.n401 B.n400 163.367
R730 B.n402 B.n401 163.367
R731 B.n402 B.n135 163.367
R732 B.n406 B.n135 163.367
R733 B.n407 B.n406 163.367
R734 B.n408 B.n407 163.367
R735 B.n408 B.n133 163.367
R736 B.n412 B.n133 163.367
R737 B.n413 B.n412 163.367
R738 B.n414 B.n413 163.367
R739 B.n414 B.n131 163.367
R740 B.n418 B.n131 163.367
R741 B.n419 B.n418 163.367
R742 B.n420 B.n419 163.367
R743 B.n420 B.n129 163.367
R744 B.n424 B.n129 163.367
R745 B.n425 B.n424 163.367
R746 B.n426 B.n425 163.367
R747 B.n426 B.n127 163.367
R748 B.n430 B.n127 163.367
R749 B.n431 B.n430 163.367
R750 B.n432 B.n431 163.367
R751 B.n432 B.n125 163.367
R752 B.n436 B.n125 163.367
R753 B.n437 B.n436 163.367
R754 B.n438 B.n437 163.367
R755 B.n438 B.n123 163.367
R756 B.n552 B.n85 163.367
R757 B.n552 B.n551 163.367
R758 B.n551 B.n550 163.367
R759 B.n550 B.n87 163.367
R760 B.n546 B.n87 163.367
R761 B.n546 B.n545 163.367
R762 B.n545 B.n544 163.367
R763 B.n544 B.n89 163.367
R764 B.n540 B.n89 163.367
R765 B.n540 B.n539 163.367
R766 B.n539 B.n538 163.367
R767 B.n538 B.n91 163.367
R768 B.n534 B.n91 163.367
R769 B.n534 B.n533 163.367
R770 B.n533 B.n532 163.367
R771 B.n532 B.n93 163.367
R772 B.n528 B.n93 163.367
R773 B.n528 B.n527 163.367
R774 B.n527 B.n526 163.367
R775 B.n526 B.n95 163.367
R776 B.n522 B.n95 163.367
R777 B.n522 B.n521 163.367
R778 B.n521 B.n520 163.367
R779 B.n520 B.n97 163.367
R780 B.n516 B.n97 163.367
R781 B.n516 B.n515 163.367
R782 B.n515 B.n514 163.367
R783 B.n514 B.n99 163.367
R784 B.n510 B.n99 163.367
R785 B.n510 B.n509 163.367
R786 B.n509 B.n508 163.367
R787 B.n508 B.n101 163.367
R788 B.n504 B.n101 163.367
R789 B.n504 B.n503 163.367
R790 B.n503 B.n502 163.367
R791 B.n502 B.n103 163.367
R792 B.n498 B.n103 163.367
R793 B.n498 B.n497 163.367
R794 B.n497 B.n496 163.367
R795 B.n496 B.n105 163.367
R796 B.n492 B.n105 163.367
R797 B.n492 B.n491 163.367
R798 B.n491 B.n490 163.367
R799 B.n490 B.n107 163.367
R800 B.n486 B.n107 163.367
R801 B.n486 B.n485 163.367
R802 B.n485 B.n484 163.367
R803 B.n484 B.n109 163.367
R804 B.n480 B.n109 163.367
R805 B.n480 B.n479 163.367
R806 B.n479 B.n478 163.367
R807 B.n478 B.n111 163.367
R808 B.n474 B.n111 163.367
R809 B.n474 B.n473 163.367
R810 B.n473 B.n472 163.367
R811 B.n472 B.n113 163.367
R812 B.n468 B.n113 163.367
R813 B.n468 B.n467 163.367
R814 B.n467 B.n466 163.367
R815 B.n466 B.n115 163.367
R816 B.n462 B.n115 163.367
R817 B.n462 B.n461 163.367
R818 B.n461 B.n460 163.367
R819 B.n460 B.n117 163.367
R820 B.n456 B.n117 163.367
R821 B.n456 B.n455 163.367
R822 B.n455 B.n454 163.367
R823 B.n454 B.n119 163.367
R824 B.n450 B.n119 163.367
R825 B.n450 B.n449 163.367
R826 B.n449 B.n448 163.367
R827 B.n448 B.n121 163.367
R828 B.n444 B.n121 163.367
R829 B.n444 B.n443 163.367
R830 B.n443 B.n442 163.367
R831 B.n736 B.n21 163.367
R832 B.n732 B.n21 163.367
R833 B.n732 B.n731 163.367
R834 B.n731 B.n730 163.367
R835 B.n730 B.n23 163.367
R836 B.n726 B.n23 163.367
R837 B.n726 B.n725 163.367
R838 B.n725 B.n724 163.367
R839 B.n724 B.n25 163.367
R840 B.n720 B.n25 163.367
R841 B.n720 B.n719 163.367
R842 B.n719 B.n718 163.367
R843 B.n718 B.n27 163.367
R844 B.n714 B.n27 163.367
R845 B.n714 B.n713 163.367
R846 B.n713 B.n712 163.367
R847 B.n712 B.n29 163.367
R848 B.n708 B.n29 163.367
R849 B.n708 B.n707 163.367
R850 B.n707 B.n706 163.367
R851 B.n706 B.n31 163.367
R852 B.n702 B.n31 163.367
R853 B.n702 B.n701 163.367
R854 B.n701 B.n700 163.367
R855 B.n700 B.n33 163.367
R856 B.n696 B.n33 163.367
R857 B.n696 B.n695 163.367
R858 B.n695 B.n694 163.367
R859 B.n694 B.n35 163.367
R860 B.n690 B.n35 163.367
R861 B.n690 B.n689 163.367
R862 B.n689 B.n688 163.367
R863 B.n688 B.n37 163.367
R864 B.n684 B.n37 163.367
R865 B.n684 B.n683 163.367
R866 B.n683 B.n682 163.367
R867 B.n682 B.n39 163.367
R868 B.n678 B.n39 163.367
R869 B.n678 B.n677 163.367
R870 B.n677 B.n676 163.367
R871 B.n676 B.n41 163.367
R872 B.n672 B.n41 163.367
R873 B.n672 B.n671 163.367
R874 B.n671 B.n670 163.367
R875 B.n670 B.n43 163.367
R876 B.n666 B.n43 163.367
R877 B.n666 B.n665 163.367
R878 B.n665 B.n664 163.367
R879 B.n664 B.n45 163.367
R880 B.n660 B.n45 163.367
R881 B.n660 B.n659 163.367
R882 B.n659 B.n658 163.367
R883 B.n658 B.n47 163.367
R884 B.n654 B.n47 163.367
R885 B.n654 B.n653 163.367
R886 B.n653 B.n51 163.367
R887 B.n649 B.n51 163.367
R888 B.n649 B.n648 163.367
R889 B.n648 B.n647 163.367
R890 B.n647 B.n53 163.367
R891 B.n643 B.n53 163.367
R892 B.n643 B.n642 163.367
R893 B.n642 B.n641 163.367
R894 B.n641 B.n55 163.367
R895 B.n636 B.n55 163.367
R896 B.n636 B.n635 163.367
R897 B.n635 B.n634 163.367
R898 B.n634 B.n59 163.367
R899 B.n630 B.n59 163.367
R900 B.n630 B.n629 163.367
R901 B.n629 B.n628 163.367
R902 B.n628 B.n61 163.367
R903 B.n624 B.n61 163.367
R904 B.n624 B.n623 163.367
R905 B.n623 B.n622 163.367
R906 B.n622 B.n63 163.367
R907 B.n618 B.n63 163.367
R908 B.n618 B.n617 163.367
R909 B.n617 B.n616 163.367
R910 B.n616 B.n65 163.367
R911 B.n612 B.n65 163.367
R912 B.n612 B.n611 163.367
R913 B.n611 B.n610 163.367
R914 B.n610 B.n67 163.367
R915 B.n606 B.n67 163.367
R916 B.n606 B.n605 163.367
R917 B.n605 B.n604 163.367
R918 B.n604 B.n69 163.367
R919 B.n600 B.n69 163.367
R920 B.n600 B.n599 163.367
R921 B.n599 B.n598 163.367
R922 B.n598 B.n71 163.367
R923 B.n594 B.n71 163.367
R924 B.n594 B.n593 163.367
R925 B.n593 B.n592 163.367
R926 B.n592 B.n73 163.367
R927 B.n588 B.n73 163.367
R928 B.n588 B.n587 163.367
R929 B.n587 B.n586 163.367
R930 B.n586 B.n75 163.367
R931 B.n582 B.n75 163.367
R932 B.n582 B.n581 163.367
R933 B.n581 B.n580 163.367
R934 B.n580 B.n77 163.367
R935 B.n576 B.n77 163.367
R936 B.n576 B.n575 163.367
R937 B.n575 B.n574 163.367
R938 B.n574 B.n79 163.367
R939 B.n570 B.n79 163.367
R940 B.n570 B.n569 163.367
R941 B.n569 B.n568 163.367
R942 B.n568 B.n81 163.367
R943 B.n564 B.n81 163.367
R944 B.n564 B.n563 163.367
R945 B.n563 B.n562 163.367
R946 B.n562 B.n83 163.367
R947 B.n558 B.n83 163.367
R948 B.n558 B.n557 163.367
R949 B.n557 B.n556 163.367
R950 B.n738 B.n737 163.367
R951 B.n738 B.n19 163.367
R952 B.n742 B.n19 163.367
R953 B.n743 B.n742 163.367
R954 B.n744 B.n743 163.367
R955 B.n744 B.n17 163.367
R956 B.n748 B.n17 163.367
R957 B.n749 B.n748 163.367
R958 B.n750 B.n749 163.367
R959 B.n750 B.n15 163.367
R960 B.n754 B.n15 163.367
R961 B.n755 B.n754 163.367
R962 B.n756 B.n755 163.367
R963 B.n756 B.n13 163.367
R964 B.n760 B.n13 163.367
R965 B.n761 B.n760 163.367
R966 B.n762 B.n761 163.367
R967 B.n762 B.n11 163.367
R968 B.n766 B.n11 163.367
R969 B.n767 B.n766 163.367
R970 B.n768 B.n767 163.367
R971 B.n768 B.n9 163.367
R972 B.n772 B.n9 163.367
R973 B.n773 B.n772 163.367
R974 B.n774 B.n773 163.367
R975 B.n774 B.n7 163.367
R976 B.n778 B.n7 163.367
R977 B.n779 B.n778 163.367
R978 B.n780 B.n779 163.367
R979 B.n780 B.n5 163.367
R980 B.n784 B.n5 163.367
R981 B.n785 B.n784 163.367
R982 B.n786 B.n785 163.367
R983 B.n786 B.n3 163.367
R984 B.n790 B.n3 163.367
R985 B.n791 B.n790 163.367
R986 B.n204 B.n2 163.367
R987 B.n205 B.n204 163.367
R988 B.n206 B.n205 163.367
R989 B.n206 B.n201 163.367
R990 B.n210 B.n201 163.367
R991 B.n211 B.n210 163.367
R992 B.n212 B.n211 163.367
R993 B.n212 B.n199 163.367
R994 B.n216 B.n199 163.367
R995 B.n217 B.n216 163.367
R996 B.n218 B.n217 163.367
R997 B.n218 B.n197 163.367
R998 B.n222 B.n197 163.367
R999 B.n223 B.n222 163.367
R1000 B.n224 B.n223 163.367
R1001 B.n224 B.n195 163.367
R1002 B.n228 B.n195 163.367
R1003 B.n229 B.n228 163.367
R1004 B.n230 B.n229 163.367
R1005 B.n230 B.n193 163.367
R1006 B.n234 B.n193 163.367
R1007 B.n235 B.n234 163.367
R1008 B.n236 B.n235 163.367
R1009 B.n236 B.n191 163.367
R1010 B.n240 B.n191 163.367
R1011 B.n241 B.n240 163.367
R1012 B.n242 B.n241 163.367
R1013 B.n242 B.n189 163.367
R1014 B.n246 B.n189 163.367
R1015 B.n247 B.n246 163.367
R1016 B.n248 B.n247 163.367
R1017 B.n248 B.n187 163.367
R1018 B.n252 B.n187 163.367
R1019 B.n253 B.n252 163.367
R1020 B.n254 B.n253 163.367
R1021 B.n254 B.n185 163.367
R1022 B.n354 B.t4 145.331
R1023 B.n56 B.t8 145.331
R1024 B.n156 B.t1 145.31
R1025 B.n48 B.t11 145.31
R1026 B.n355 B.t5 112.749
R1027 B.n57 B.t7 112.749
R1028 B.n157 B.t2 112.728
R1029 B.n49 B.t10 112.728
R1030 B.n340 B.n157 59.5399
R1031 B.n356 B.n355 59.5399
R1032 B.n638 B.n57 59.5399
R1033 B.n50 B.n49 59.5399
R1034 B.n441 B.n440 36.059
R1035 B.n735 B.n20 36.059
R1036 B.n555 B.n554 36.059
R1037 B.n257 B.n256 36.059
R1038 B.n157 B.n156 32.5823
R1039 B.n355 B.n354 32.5823
R1040 B.n57 B.n56 32.5823
R1041 B.n49 B.n48 32.5823
R1042 B B.n793 18.0485
R1043 B.n739 B.n20 10.6151
R1044 B.n740 B.n739 10.6151
R1045 B.n741 B.n740 10.6151
R1046 B.n741 B.n18 10.6151
R1047 B.n745 B.n18 10.6151
R1048 B.n746 B.n745 10.6151
R1049 B.n747 B.n746 10.6151
R1050 B.n747 B.n16 10.6151
R1051 B.n751 B.n16 10.6151
R1052 B.n752 B.n751 10.6151
R1053 B.n753 B.n752 10.6151
R1054 B.n753 B.n14 10.6151
R1055 B.n757 B.n14 10.6151
R1056 B.n758 B.n757 10.6151
R1057 B.n759 B.n758 10.6151
R1058 B.n759 B.n12 10.6151
R1059 B.n763 B.n12 10.6151
R1060 B.n764 B.n763 10.6151
R1061 B.n765 B.n764 10.6151
R1062 B.n765 B.n10 10.6151
R1063 B.n769 B.n10 10.6151
R1064 B.n770 B.n769 10.6151
R1065 B.n771 B.n770 10.6151
R1066 B.n771 B.n8 10.6151
R1067 B.n775 B.n8 10.6151
R1068 B.n776 B.n775 10.6151
R1069 B.n777 B.n776 10.6151
R1070 B.n777 B.n6 10.6151
R1071 B.n781 B.n6 10.6151
R1072 B.n782 B.n781 10.6151
R1073 B.n783 B.n782 10.6151
R1074 B.n783 B.n4 10.6151
R1075 B.n787 B.n4 10.6151
R1076 B.n788 B.n787 10.6151
R1077 B.n789 B.n788 10.6151
R1078 B.n789 B.n0 10.6151
R1079 B.n735 B.n734 10.6151
R1080 B.n734 B.n733 10.6151
R1081 B.n733 B.n22 10.6151
R1082 B.n729 B.n22 10.6151
R1083 B.n729 B.n728 10.6151
R1084 B.n728 B.n727 10.6151
R1085 B.n727 B.n24 10.6151
R1086 B.n723 B.n24 10.6151
R1087 B.n723 B.n722 10.6151
R1088 B.n722 B.n721 10.6151
R1089 B.n721 B.n26 10.6151
R1090 B.n717 B.n26 10.6151
R1091 B.n717 B.n716 10.6151
R1092 B.n716 B.n715 10.6151
R1093 B.n715 B.n28 10.6151
R1094 B.n711 B.n28 10.6151
R1095 B.n711 B.n710 10.6151
R1096 B.n710 B.n709 10.6151
R1097 B.n709 B.n30 10.6151
R1098 B.n705 B.n30 10.6151
R1099 B.n705 B.n704 10.6151
R1100 B.n704 B.n703 10.6151
R1101 B.n703 B.n32 10.6151
R1102 B.n699 B.n32 10.6151
R1103 B.n699 B.n698 10.6151
R1104 B.n698 B.n697 10.6151
R1105 B.n697 B.n34 10.6151
R1106 B.n693 B.n34 10.6151
R1107 B.n693 B.n692 10.6151
R1108 B.n692 B.n691 10.6151
R1109 B.n691 B.n36 10.6151
R1110 B.n687 B.n36 10.6151
R1111 B.n687 B.n686 10.6151
R1112 B.n686 B.n685 10.6151
R1113 B.n685 B.n38 10.6151
R1114 B.n681 B.n38 10.6151
R1115 B.n681 B.n680 10.6151
R1116 B.n680 B.n679 10.6151
R1117 B.n679 B.n40 10.6151
R1118 B.n675 B.n40 10.6151
R1119 B.n675 B.n674 10.6151
R1120 B.n674 B.n673 10.6151
R1121 B.n673 B.n42 10.6151
R1122 B.n669 B.n42 10.6151
R1123 B.n669 B.n668 10.6151
R1124 B.n668 B.n667 10.6151
R1125 B.n667 B.n44 10.6151
R1126 B.n663 B.n44 10.6151
R1127 B.n663 B.n662 10.6151
R1128 B.n662 B.n661 10.6151
R1129 B.n661 B.n46 10.6151
R1130 B.n657 B.n46 10.6151
R1131 B.n657 B.n656 10.6151
R1132 B.n656 B.n655 10.6151
R1133 B.n652 B.n651 10.6151
R1134 B.n651 B.n650 10.6151
R1135 B.n650 B.n52 10.6151
R1136 B.n646 B.n52 10.6151
R1137 B.n646 B.n645 10.6151
R1138 B.n645 B.n644 10.6151
R1139 B.n644 B.n54 10.6151
R1140 B.n640 B.n54 10.6151
R1141 B.n640 B.n639 10.6151
R1142 B.n637 B.n58 10.6151
R1143 B.n633 B.n58 10.6151
R1144 B.n633 B.n632 10.6151
R1145 B.n632 B.n631 10.6151
R1146 B.n631 B.n60 10.6151
R1147 B.n627 B.n60 10.6151
R1148 B.n627 B.n626 10.6151
R1149 B.n626 B.n625 10.6151
R1150 B.n625 B.n62 10.6151
R1151 B.n621 B.n62 10.6151
R1152 B.n621 B.n620 10.6151
R1153 B.n620 B.n619 10.6151
R1154 B.n619 B.n64 10.6151
R1155 B.n615 B.n64 10.6151
R1156 B.n615 B.n614 10.6151
R1157 B.n614 B.n613 10.6151
R1158 B.n613 B.n66 10.6151
R1159 B.n609 B.n66 10.6151
R1160 B.n609 B.n608 10.6151
R1161 B.n608 B.n607 10.6151
R1162 B.n607 B.n68 10.6151
R1163 B.n603 B.n68 10.6151
R1164 B.n603 B.n602 10.6151
R1165 B.n602 B.n601 10.6151
R1166 B.n601 B.n70 10.6151
R1167 B.n597 B.n70 10.6151
R1168 B.n597 B.n596 10.6151
R1169 B.n596 B.n595 10.6151
R1170 B.n595 B.n72 10.6151
R1171 B.n591 B.n72 10.6151
R1172 B.n591 B.n590 10.6151
R1173 B.n590 B.n589 10.6151
R1174 B.n589 B.n74 10.6151
R1175 B.n585 B.n74 10.6151
R1176 B.n585 B.n584 10.6151
R1177 B.n584 B.n583 10.6151
R1178 B.n583 B.n76 10.6151
R1179 B.n579 B.n76 10.6151
R1180 B.n579 B.n578 10.6151
R1181 B.n578 B.n577 10.6151
R1182 B.n577 B.n78 10.6151
R1183 B.n573 B.n78 10.6151
R1184 B.n573 B.n572 10.6151
R1185 B.n572 B.n571 10.6151
R1186 B.n571 B.n80 10.6151
R1187 B.n567 B.n80 10.6151
R1188 B.n567 B.n566 10.6151
R1189 B.n566 B.n565 10.6151
R1190 B.n565 B.n82 10.6151
R1191 B.n561 B.n82 10.6151
R1192 B.n561 B.n560 10.6151
R1193 B.n560 B.n559 10.6151
R1194 B.n559 B.n84 10.6151
R1195 B.n555 B.n84 10.6151
R1196 B.n554 B.n553 10.6151
R1197 B.n553 B.n86 10.6151
R1198 B.n549 B.n86 10.6151
R1199 B.n549 B.n548 10.6151
R1200 B.n548 B.n547 10.6151
R1201 B.n547 B.n88 10.6151
R1202 B.n543 B.n88 10.6151
R1203 B.n543 B.n542 10.6151
R1204 B.n542 B.n541 10.6151
R1205 B.n541 B.n90 10.6151
R1206 B.n537 B.n90 10.6151
R1207 B.n537 B.n536 10.6151
R1208 B.n536 B.n535 10.6151
R1209 B.n535 B.n92 10.6151
R1210 B.n531 B.n92 10.6151
R1211 B.n531 B.n530 10.6151
R1212 B.n530 B.n529 10.6151
R1213 B.n529 B.n94 10.6151
R1214 B.n525 B.n94 10.6151
R1215 B.n525 B.n524 10.6151
R1216 B.n524 B.n523 10.6151
R1217 B.n523 B.n96 10.6151
R1218 B.n519 B.n96 10.6151
R1219 B.n519 B.n518 10.6151
R1220 B.n518 B.n517 10.6151
R1221 B.n517 B.n98 10.6151
R1222 B.n513 B.n98 10.6151
R1223 B.n513 B.n512 10.6151
R1224 B.n512 B.n511 10.6151
R1225 B.n511 B.n100 10.6151
R1226 B.n507 B.n100 10.6151
R1227 B.n507 B.n506 10.6151
R1228 B.n506 B.n505 10.6151
R1229 B.n505 B.n102 10.6151
R1230 B.n501 B.n102 10.6151
R1231 B.n501 B.n500 10.6151
R1232 B.n500 B.n499 10.6151
R1233 B.n499 B.n104 10.6151
R1234 B.n495 B.n104 10.6151
R1235 B.n495 B.n494 10.6151
R1236 B.n494 B.n493 10.6151
R1237 B.n493 B.n106 10.6151
R1238 B.n489 B.n106 10.6151
R1239 B.n489 B.n488 10.6151
R1240 B.n488 B.n487 10.6151
R1241 B.n487 B.n108 10.6151
R1242 B.n483 B.n108 10.6151
R1243 B.n483 B.n482 10.6151
R1244 B.n482 B.n481 10.6151
R1245 B.n481 B.n110 10.6151
R1246 B.n477 B.n110 10.6151
R1247 B.n477 B.n476 10.6151
R1248 B.n476 B.n475 10.6151
R1249 B.n475 B.n112 10.6151
R1250 B.n471 B.n112 10.6151
R1251 B.n471 B.n470 10.6151
R1252 B.n470 B.n469 10.6151
R1253 B.n469 B.n114 10.6151
R1254 B.n465 B.n114 10.6151
R1255 B.n465 B.n464 10.6151
R1256 B.n464 B.n463 10.6151
R1257 B.n463 B.n116 10.6151
R1258 B.n459 B.n116 10.6151
R1259 B.n459 B.n458 10.6151
R1260 B.n458 B.n457 10.6151
R1261 B.n457 B.n118 10.6151
R1262 B.n453 B.n118 10.6151
R1263 B.n453 B.n452 10.6151
R1264 B.n452 B.n451 10.6151
R1265 B.n451 B.n120 10.6151
R1266 B.n447 B.n120 10.6151
R1267 B.n447 B.n446 10.6151
R1268 B.n446 B.n445 10.6151
R1269 B.n445 B.n122 10.6151
R1270 B.n441 B.n122 10.6151
R1271 B.n203 B.n1 10.6151
R1272 B.n203 B.n202 10.6151
R1273 B.n207 B.n202 10.6151
R1274 B.n208 B.n207 10.6151
R1275 B.n209 B.n208 10.6151
R1276 B.n209 B.n200 10.6151
R1277 B.n213 B.n200 10.6151
R1278 B.n214 B.n213 10.6151
R1279 B.n215 B.n214 10.6151
R1280 B.n215 B.n198 10.6151
R1281 B.n219 B.n198 10.6151
R1282 B.n220 B.n219 10.6151
R1283 B.n221 B.n220 10.6151
R1284 B.n221 B.n196 10.6151
R1285 B.n225 B.n196 10.6151
R1286 B.n226 B.n225 10.6151
R1287 B.n227 B.n226 10.6151
R1288 B.n227 B.n194 10.6151
R1289 B.n231 B.n194 10.6151
R1290 B.n232 B.n231 10.6151
R1291 B.n233 B.n232 10.6151
R1292 B.n233 B.n192 10.6151
R1293 B.n237 B.n192 10.6151
R1294 B.n238 B.n237 10.6151
R1295 B.n239 B.n238 10.6151
R1296 B.n239 B.n190 10.6151
R1297 B.n243 B.n190 10.6151
R1298 B.n244 B.n243 10.6151
R1299 B.n245 B.n244 10.6151
R1300 B.n245 B.n188 10.6151
R1301 B.n249 B.n188 10.6151
R1302 B.n250 B.n249 10.6151
R1303 B.n251 B.n250 10.6151
R1304 B.n251 B.n186 10.6151
R1305 B.n255 B.n186 10.6151
R1306 B.n256 B.n255 10.6151
R1307 B.n257 B.n184 10.6151
R1308 B.n261 B.n184 10.6151
R1309 B.n262 B.n261 10.6151
R1310 B.n263 B.n262 10.6151
R1311 B.n263 B.n182 10.6151
R1312 B.n267 B.n182 10.6151
R1313 B.n268 B.n267 10.6151
R1314 B.n269 B.n268 10.6151
R1315 B.n269 B.n180 10.6151
R1316 B.n273 B.n180 10.6151
R1317 B.n274 B.n273 10.6151
R1318 B.n275 B.n274 10.6151
R1319 B.n275 B.n178 10.6151
R1320 B.n279 B.n178 10.6151
R1321 B.n280 B.n279 10.6151
R1322 B.n281 B.n280 10.6151
R1323 B.n281 B.n176 10.6151
R1324 B.n285 B.n176 10.6151
R1325 B.n286 B.n285 10.6151
R1326 B.n287 B.n286 10.6151
R1327 B.n287 B.n174 10.6151
R1328 B.n291 B.n174 10.6151
R1329 B.n292 B.n291 10.6151
R1330 B.n293 B.n292 10.6151
R1331 B.n293 B.n172 10.6151
R1332 B.n297 B.n172 10.6151
R1333 B.n298 B.n297 10.6151
R1334 B.n299 B.n298 10.6151
R1335 B.n299 B.n170 10.6151
R1336 B.n303 B.n170 10.6151
R1337 B.n304 B.n303 10.6151
R1338 B.n305 B.n304 10.6151
R1339 B.n305 B.n168 10.6151
R1340 B.n309 B.n168 10.6151
R1341 B.n310 B.n309 10.6151
R1342 B.n311 B.n310 10.6151
R1343 B.n311 B.n166 10.6151
R1344 B.n315 B.n166 10.6151
R1345 B.n316 B.n315 10.6151
R1346 B.n317 B.n316 10.6151
R1347 B.n317 B.n164 10.6151
R1348 B.n321 B.n164 10.6151
R1349 B.n322 B.n321 10.6151
R1350 B.n323 B.n322 10.6151
R1351 B.n323 B.n162 10.6151
R1352 B.n327 B.n162 10.6151
R1353 B.n328 B.n327 10.6151
R1354 B.n329 B.n328 10.6151
R1355 B.n329 B.n160 10.6151
R1356 B.n333 B.n160 10.6151
R1357 B.n334 B.n333 10.6151
R1358 B.n335 B.n334 10.6151
R1359 B.n335 B.n158 10.6151
R1360 B.n339 B.n158 10.6151
R1361 B.n342 B.n341 10.6151
R1362 B.n342 B.n154 10.6151
R1363 B.n346 B.n154 10.6151
R1364 B.n347 B.n346 10.6151
R1365 B.n348 B.n347 10.6151
R1366 B.n348 B.n152 10.6151
R1367 B.n352 B.n152 10.6151
R1368 B.n353 B.n352 10.6151
R1369 B.n357 B.n353 10.6151
R1370 B.n361 B.n150 10.6151
R1371 B.n362 B.n361 10.6151
R1372 B.n363 B.n362 10.6151
R1373 B.n363 B.n148 10.6151
R1374 B.n367 B.n148 10.6151
R1375 B.n368 B.n367 10.6151
R1376 B.n369 B.n368 10.6151
R1377 B.n369 B.n146 10.6151
R1378 B.n373 B.n146 10.6151
R1379 B.n374 B.n373 10.6151
R1380 B.n375 B.n374 10.6151
R1381 B.n375 B.n144 10.6151
R1382 B.n379 B.n144 10.6151
R1383 B.n380 B.n379 10.6151
R1384 B.n381 B.n380 10.6151
R1385 B.n381 B.n142 10.6151
R1386 B.n385 B.n142 10.6151
R1387 B.n386 B.n385 10.6151
R1388 B.n387 B.n386 10.6151
R1389 B.n387 B.n140 10.6151
R1390 B.n391 B.n140 10.6151
R1391 B.n392 B.n391 10.6151
R1392 B.n393 B.n392 10.6151
R1393 B.n393 B.n138 10.6151
R1394 B.n397 B.n138 10.6151
R1395 B.n398 B.n397 10.6151
R1396 B.n399 B.n398 10.6151
R1397 B.n399 B.n136 10.6151
R1398 B.n403 B.n136 10.6151
R1399 B.n404 B.n403 10.6151
R1400 B.n405 B.n404 10.6151
R1401 B.n405 B.n134 10.6151
R1402 B.n409 B.n134 10.6151
R1403 B.n410 B.n409 10.6151
R1404 B.n411 B.n410 10.6151
R1405 B.n411 B.n132 10.6151
R1406 B.n415 B.n132 10.6151
R1407 B.n416 B.n415 10.6151
R1408 B.n417 B.n416 10.6151
R1409 B.n417 B.n130 10.6151
R1410 B.n421 B.n130 10.6151
R1411 B.n422 B.n421 10.6151
R1412 B.n423 B.n422 10.6151
R1413 B.n423 B.n128 10.6151
R1414 B.n427 B.n128 10.6151
R1415 B.n428 B.n427 10.6151
R1416 B.n429 B.n428 10.6151
R1417 B.n429 B.n126 10.6151
R1418 B.n433 B.n126 10.6151
R1419 B.n434 B.n433 10.6151
R1420 B.n435 B.n434 10.6151
R1421 B.n435 B.n124 10.6151
R1422 B.n439 B.n124 10.6151
R1423 B.n440 B.n439 10.6151
R1424 B.n655 B.n50 9.36635
R1425 B.n638 B.n637 9.36635
R1426 B.n340 B.n339 9.36635
R1427 B.n356 B.n150 9.36635
R1428 B.n793 B.n0 8.11757
R1429 B.n793 B.n1 8.11757
R1430 B.n652 B.n50 1.24928
R1431 B.n639 B.n638 1.24928
R1432 B.n341 B.n340 1.24928
R1433 B.n357 B.n356 1.24928
C0 VTAIL VDD1 14.2665f
C1 w_n2986_n4298# VN 6.08777f
C2 B w_n2986_n4298# 9.74832f
C3 VP VDD2 0.424677f
C4 VN VDD1 0.150358f
C5 B VDD1 2.33144f
C6 VN VTAIL 12.155701f
C7 B VTAIL 4.05464f
C8 VP w_n2986_n4298# 6.47268f
C9 w_n2986_n4298# VDD2 2.72012f
C10 VP VDD1 12.4863f
C11 B VN 1.01975f
C12 VDD2 VDD1 1.36184f
C13 VP VTAIL 12.1703f
C14 VDD2 VTAIL 14.305201f
C15 VP VN 7.41371f
C16 VP B 1.66009f
C17 w_n2986_n4298# VDD1 2.64153f
C18 VDD2 VN 12.217401f
C19 B VDD2 2.40068f
C20 w_n2986_n4298# VTAIL 3.74644f
C21 VDD2 VSUBS 1.826911f
C22 VDD1 VSUBS 1.586637f
C23 VTAIL VSUBS 1.146989f
C24 VN VSUBS 6.022861f
C25 VP VSUBS 2.830906f
C26 B VSUBS 4.209857f
C27 w_n2986_n4298# VSUBS 0.157123p
C28 B.n0 VSUBS 0.007479f
C29 B.n1 VSUBS 0.007479f
C30 B.n2 VSUBS 0.011061f
C31 B.n3 VSUBS 0.008476f
C32 B.n4 VSUBS 0.008476f
C33 B.n5 VSUBS 0.008476f
C34 B.n6 VSUBS 0.008476f
C35 B.n7 VSUBS 0.008476f
C36 B.n8 VSUBS 0.008476f
C37 B.n9 VSUBS 0.008476f
C38 B.n10 VSUBS 0.008476f
C39 B.n11 VSUBS 0.008476f
C40 B.n12 VSUBS 0.008476f
C41 B.n13 VSUBS 0.008476f
C42 B.n14 VSUBS 0.008476f
C43 B.n15 VSUBS 0.008476f
C44 B.n16 VSUBS 0.008476f
C45 B.n17 VSUBS 0.008476f
C46 B.n18 VSUBS 0.008476f
C47 B.n19 VSUBS 0.008476f
C48 B.n20 VSUBS 0.020626f
C49 B.n21 VSUBS 0.008476f
C50 B.n22 VSUBS 0.008476f
C51 B.n23 VSUBS 0.008476f
C52 B.n24 VSUBS 0.008476f
C53 B.n25 VSUBS 0.008476f
C54 B.n26 VSUBS 0.008476f
C55 B.n27 VSUBS 0.008476f
C56 B.n28 VSUBS 0.008476f
C57 B.n29 VSUBS 0.008476f
C58 B.n30 VSUBS 0.008476f
C59 B.n31 VSUBS 0.008476f
C60 B.n32 VSUBS 0.008476f
C61 B.n33 VSUBS 0.008476f
C62 B.n34 VSUBS 0.008476f
C63 B.n35 VSUBS 0.008476f
C64 B.n36 VSUBS 0.008476f
C65 B.n37 VSUBS 0.008476f
C66 B.n38 VSUBS 0.008476f
C67 B.n39 VSUBS 0.008476f
C68 B.n40 VSUBS 0.008476f
C69 B.n41 VSUBS 0.008476f
C70 B.n42 VSUBS 0.008476f
C71 B.n43 VSUBS 0.008476f
C72 B.n44 VSUBS 0.008476f
C73 B.n45 VSUBS 0.008476f
C74 B.n46 VSUBS 0.008476f
C75 B.n47 VSUBS 0.008476f
C76 B.t10 VSUBS 0.676804f
C77 B.t11 VSUBS 0.692246f
C78 B.t9 VSUBS 1.15417f
C79 B.n48 VSUBS 0.289454f
C80 B.n49 VSUBS 0.080958f
C81 B.n50 VSUBS 0.019638f
C82 B.n51 VSUBS 0.008476f
C83 B.n52 VSUBS 0.008476f
C84 B.n53 VSUBS 0.008476f
C85 B.n54 VSUBS 0.008476f
C86 B.n55 VSUBS 0.008476f
C87 B.t7 VSUBS 0.676782f
C88 B.t8 VSUBS 0.692227f
C89 B.t6 VSUBS 1.15417f
C90 B.n56 VSUBS 0.289473f
C91 B.n57 VSUBS 0.08098f
C92 B.n58 VSUBS 0.008476f
C93 B.n59 VSUBS 0.008476f
C94 B.n60 VSUBS 0.008476f
C95 B.n61 VSUBS 0.008476f
C96 B.n62 VSUBS 0.008476f
C97 B.n63 VSUBS 0.008476f
C98 B.n64 VSUBS 0.008476f
C99 B.n65 VSUBS 0.008476f
C100 B.n66 VSUBS 0.008476f
C101 B.n67 VSUBS 0.008476f
C102 B.n68 VSUBS 0.008476f
C103 B.n69 VSUBS 0.008476f
C104 B.n70 VSUBS 0.008476f
C105 B.n71 VSUBS 0.008476f
C106 B.n72 VSUBS 0.008476f
C107 B.n73 VSUBS 0.008476f
C108 B.n74 VSUBS 0.008476f
C109 B.n75 VSUBS 0.008476f
C110 B.n76 VSUBS 0.008476f
C111 B.n77 VSUBS 0.008476f
C112 B.n78 VSUBS 0.008476f
C113 B.n79 VSUBS 0.008476f
C114 B.n80 VSUBS 0.008476f
C115 B.n81 VSUBS 0.008476f
C116 B.n82 VSUBS 0.008476f
C117 B.n83 VSUBS 0.008476f
C118 B.n84 VSUBS 0.008476f
C119 B.n85 VSUBS 0.020626f
C120 B.n86 VSUBS 0.008476f
C121 B.n87 VSUBS 0.008476f
C122 B.n88 VSUBS 0.008476f
C123 B.n89 VSUBS 0.008476f
C124 B.n90 VSUBS 0.008476f
C125 B.n91 VSUBS 0.008476f
C126 B.n92 VSUBS 0.008476f
C127 B.n93 VSUBS 0.008476f
C128 B.n94 VSUBS 0.008476f
C129 B.n95 VSUBS 0.008476f
C130 B.n96 VSUBS 0.008476f
C131 B.n97 VSUBS 0.008476f
C132 B.n98 VSUBS 0.008476f
C133 B.n99 VSUBS 0.008476f
C134 B.n100 VSUBS 0.008476f
C135 B.n101 VSUBS 0.008476f
C136 B.n102 VSUBS 0.008476f
C137 B.n103 VSUBS 0.008476f
C138 B.n104 VSUBS 0.008476f
C139 B.n105 VSUBS 0.008476f
C140 B.n106 VSUBS 0.008476f
C141 B.n107 VSUBS 0.008476f
C142 B.n108 VSUBS 0.008476f
C143 B.n109 VSUBS 0.008476f
C144 B.n110 VSUBS 0.008476f
C145 B.n111 VSUBS 0.008476f
C146 B.n112 VSUBS 0.008476f
C147 B.n113 VSUBS 0.008476f
C148 B.n114 VSUBS 0.008476f
C149 B.n115 VSUBS 0.008476f
C150 B.n116 VSUBS 0.008476f
C151 B.n117 VSUBS 0.008476f
C152 B.n118 VSUBS 0.008476f
C153 B.n119 VSUBS 0.008476f
C154 B.n120 VSUBS 0.008476f
C155 B.n121 VSUBS 0.008476f
C156 B.n122 VSUBS 0.008476f
C157 B.n123 VSUBS 0.021754f
C158 B.n124 VSUBS 0.008476f
C159 B.n125 VSUBS 0.008476f
C160 B.n126 VSUBS 0.008476f
C161 B.n127 VSUBS 0.008476f
C162 B.n128 VSUBS 0.008476f
C163 B.n129 VSUBS 0.008476f
C164 B.n130 VSUBS 0.008476f
C165 B.n131 VSUBS 0.008476f
C166 B.n132 VSUBS 0.008476f
C167 B.n133 VSUBS 0.008476f
C168 B.n134 VSUBS 0.008476f
C169 B.n135 VSUBS 0.008476f
C170 B.n136 VSUBS 0.008476f
C171 B.n137 VSUBS 0.008476f
C172 B.n138 VSUBS 0.008476f
C173 B.n139 VSUBS 0.008476f
C174 B.n140 VSUBS 0.008476f
C175 B.n141 VSUBS 0.008476f
C176 B.n142 VSUBS 0.008476f
C177 B.n143 VSUBS 0.008476f
C178 B.n144 VSUBS 0.008476f
C179 B.n145 VSUBS 0.008476f
C180 B.n146 VSUBS 0.008476f
C181 B.n147 VSUBS 0.008476f
C182 B.n148 VSUBS 0.008476f
C183 B.n149 VSUBS 0.008476f
C184 B.n150 VSUBS 0.007977f
C185 B.n151 VSUBS 0.008476f
C186 B.n152 VSUBS 0.008476f
C187 B.n153 VSUBS 0.008476f
C188 B.n154 VSUBS 0.008476f
C189 B.n155 VSUBS 0.008476f
C190 B.t2 VSUBS 0.676804f
C191 B.t1 VSUBS 0.692246f
C192 B.t0 VSUBS 1.15417f
C193 B.n156 VSUBS 0.289454f
C194 B.n157 VSUBS 0.080958f
C195 B.n158 VSUBS 0.008476f
C196 B.n159 VSUBS 0.008476f
C197 B.n160 VSUBS 0.008476f
C198 B.n161 VSUBS 0.008476f
C199 B.n162 VSUBS 0.008476f
C200 B.n163 VSUBS 0.008476f
C201 B.n164 VSUBS 0.008476f
C202 B.n165 VSUBS 0.008476f
C203 B.n166 VSUBS 0.008476f
C204 B.n167 VSUBS 0.008476f
C205 B.n168 VSUBS 0.008476f
C206 B.n169 VSUBS 0.008476f
C207 B.n170 VSUBS 0.008476f
C208 B.n171 VSUBS 0.008476f
C209 B.n172 VSUBS 0.008476f
C210 B.n173 VSUBS 0.008476f
C211 B.n174 VSUBS 0.008476f
C212 B.n175 VSUBS 0.008476f
C213 B.n176 VSUBS 0.008476f
C214 B.n177 VSUBS 0.008476f
C215 B.n178 VSUBS 0.008476f
C216 B.n179 VSUBS 0.008476f
C217 B.n180 VSUBS 0.008476f
C218 B.n181 VSUBS 0.008476f
C219 B.n182 VSUBS 0.008476f
C220 B.n183 VSUBS 0.008476f
C221 B.n184 VSUBS 0.008476f
C222 B.n185 VSUBS 0.020626f
C223 B.n186 VSUBS 0.008476f
C224 B.n187 VSUBS 0.008476f
C225 B.n188 VSUBS 0.008476f
C226 B.n189 VSUBS 0.008476f
C227 B.n190 VSUBS 0.008476f
C228 B.n191 VSUBS 0.008476f
C229 B.n192 VSUBS 0.008476f
C230 B.n193 VSUBS 0.008476f
C231 B.n194 VSUBS 0.008476f
C232 B.n195 VSUBS 0.008476f
C233 B.n196 VSUBS 0.008476f
C234 B.n197 VSUBS 0.008476f
C235 B.n198 VSUBS 0.008476f
C236 B.n199 VSUBS 0.008476f
C237 B.n200 VSUBS 0.008476f
C238 B.n201 VSUBS 0.008476f
C239 B.n202 VSUBS 0.008476f
C240 B.n203 VSUBS 0.008476f
C241 B.n204 VSUBS 0.008476f
C242 B.n205 VSUBS 0.008476f
C243 B.n206 VSUBS 0.008476f
C244 B.n207 VSUBS 0.008476f
C245 B.n208 VSUBS 0.008476f
C246 B.n209 VSUBS 0.008476f
C247 B.n210 VSUBS 0.008476f
C248 B.n211 VSUBS 0.008476f
C249 B.n212 VSUBS 0.008476f
C250 B.n213 VSUBS 0.008476f
C251 B.n214 VSUBS 0.008476f
C252 B.n215 VSUBS 0.008476f
C253 B.n216 VSUBS 0.008476f
C254 B.n217 VSUBS 0.008476f
C255 B.n218 VSUBS 0.008476f
C256 B.n219 VSUBS 0.008476f
C257 B.n220 VSUBS 0.008476f
C258 B.n221 VSUBS 0.008476f
C259 B.n222 VSUBS 0.008476f
C260 B.n223 VSUBS 0.008476f
C261 B.n224 VSUBS 0.008476f
C262 B.n225 VSUBS 0.008476f
C263 B.n226 VSUBS 0.008476f
C264 B.n227 VSUBS 0.008476f
C265 B.n228 VSUBS 0.008476f
C266 B.n229 VSUBS 0.008476f
C267 B.n230 VSUBS 0.008476f
C268 B.n231 VSUBS 0.008476f
C269 B.n232 VSUBS 0.008476f
C270 B.n233 VSUBS 0.008476f
C271 B.n234 VSUBS 0.008476f
C272 B.n235 VSUBS 0.008476f
C273 B.n236 VSUBS 0.008476f
C274 B.n237 VSUBS 0.008476f
C275 B.n238 VSUBS 0.008476f
C276 B.n239 VSUBS 0.008476f
C277 B.n240 VSUBS 0.008476f
C278 B.n241 VSUBS 0.008476f
C279 B.n242 VSUBS 0.008476f
C280 B.n243 VSUBS 0.008476f
C281 B.n244 VSUBS 0.008476f
C282 B.n245 VSUBS 0.008476f
C283 B.n246 VSUBS 0.008476f
C284 B.n247 VSUBS 0.008476f
C285 B.n248 VSUBS 0.008476f
C286 B.n249 VSUBS 0.008476f
C287 B.n250 VSUBS 0.008476f
C288 B.n251 VSUBS 0.008476f
C289 B.n252 VSUBS 0.008476f
C290 B.n253 VSUBS 0.008476f
C291 B.n254 VSUBS 0.008476f
C292 B.n255 VSUBS 0.008476f
C293 B.n256 VSUBS 0.020626f
C294 B.n257 VSUBS 0.021754f
C295 B.n258 VSUBS 0.021754f
C296 B.n259 VSUBS 0.008476f
C297 B.n260 VSUBS 0.008476f
C298 B.n261 VSUBS 0.008476f
C299 B.n262 VSUBS 0.008476f
C300 B.n263 VSUBS 0.008476f
C301 B.n264 VSUBS 0.008476f
C302 B.n265 VSUBS 0.008476f
C303 B.n266 VSUBS 0.008476f
C304 B.n267 VSUBS 0.008476f
C305 B.n268 VSUBS 0.008476f
C306 B.n269 VSUBS 0.008476f
C307 B.n270 VSUBS 0.008476f
C308 B.n271 VSUBS 0.008476f
C309 B.n272 VSUBS 0.008476f
C310 B.n273 VSUBS 0.008476f
C311 B.n274 VSUBS 0.008476f
C312 B.n275 VSUBS 0.008476f
C313 B.n276 VSUBS 0.008476f
C314 B.n277 VSUBS 0.008476f
C315 B.n278 VSUBS 0.008476f
C316 B.n279 VSUBS 0.008476f
C317 B.n280 VSUBS 0.008476f
C318 B.n281 VSUBS 0.008476f
C319 B.n282 VSUBS 0.008476f
C320 B.n283 VSUBS 0.008476f
C321 B.n284 VSUBS 0.008476f
C322 B.n285 VSUBS 0.008476f
C323 B.n286 VSUBS 0.008476f
C324 B.n287 VSUBS 0.008476f
C325 B.n288 VSUBS 0.008476f
C326 B.n289 VSUBS 0.008476f
C327 B.n290 VSUBS 0.008476f
C328 B.n291 VSUBS 0.008476f
C329 B.n292 VSUBS 0.008476f
C330 B.n293 VSUBS 0.008476f
C331 B.n294 VSUBS 0.008476f
C332 B.n295 VSUBS 0.008476f
C333 B.n296 VSUBS 0.008476f
C334 B.n297 VSUBS 0.008476f
C335 B.n298 VSUBS 0.008476f
C336 B.n299 VSUBS 0.008476f
C337 B.n300 VSUBS 0.008476f
C338 B.n301 VSUBS 0.008476f
C339 B.n302 VSUBS 0.008476f
C340 B.n303 VSUBS 0.008476f
C341 B.n304 VSUBS 0.008476f
C342 B.n305 VSUBS 0.008476f
C343 B.n306 VSUBS 0.008476f
C344 B.n307 VSUBS 0.008476f
C345 B.n308 VSUBS 0.008476f
C346 B.n309 VSUBS 0.008476f
C347 B.n310 VSUBS 0.008476f
C348 B.n311 VSUBS 0.008476f
C349 B.n312 VSUBS 0.008476f
C350 B.n313 VSUBS 0.008476f
C351 B.n314 VSUBS 0.008476f
C352 B.n315 VSUBS 0.008476f
C353 B.n316 VSUBS 0.008476f
C354 B.n317 VSUBS 0.008476f
C355 B.n318 VSUBS 0.008476f
C356 B.n319 VSUBS 0.008476f
C357 B.n320 VSUBS 0.008476f
C358 B.n321 VSUBS 0.008476f
C359 B.n322 VSUBS 0.008476f
C360 B.n323 VSUBS 0.008476f
C361 B.n324 VSUBS 0.008476f
C362 B.n325 VSUBS 0.008476f
C363 B.n326 VSUBS 0.008476f
C364 B.n327 VSUBS 0.008476f
C365 B.n328 VSUBS 0.008476f
C366 B.n329 VSUBS 0.008476f
C367 B.n330 VSUBS 0.008476f
C368 B.n331 VSUBS 0.008476f
C369 B.n332 VSUBS 0.008476f
C370 B.n333 VSUBS 0.008476f
C371 B.n334 VSUBS 0.008476f
C372 B.n335 VSUBS 0.008476f
C373 B.n336 VSUBS 0.008476f
C374 B.n337 VSUBS 0.008476f
C375 B.n338 VSUBS 0.008476f
C376 B.n339 VSUBS 0.007977f
C377 B.n340 VSUBS 0.019638f
C378 B.n341 VSUBS 0.004737f
C379 B.n342 VSUBS 0.008476f
C380 B.n343 VSUBS 0.008476f
C381 B.n344 VSUBS 0.008476f
C382 B.n345 VSUBS 0.008476f
C383 B.n346 VSUBS 0.008476f
C384 B.n347 VSUBS 0.008476f
C385 B.n348 VSUBS 0.008476f
C386 B.n349 VSUBS 0.008476f
C387 B.n350 VSUBS 0.008476f
C388 B.n351 VSUBS 0.008476f
C389 B.n352 VSUBS 0.008476f
C390 B.n353 VSUBS 0.008476f
C391 B.t5 VSUBS 0.676782f
C392 B.t4 VSUBS 0.692227f
C393 B.t3 VSUBS 1.15417f
C394 B.n354 VSUBS 0.289473f
C395 B.n355 VSUBS 0.08098f
C396 B.n356 VSUBS 0.019638f
C397 B.n357 VSUBS 0.004737f
C398 B.n358 VSUBS 0.008476f
C399 B.n359 VSUBS 0.008476f
C400 B.n360 VSUBS 0.008476f
C401 B.n361 VSUBS 0.008476f
C402 B.n362 VSUBS 0.008476f
C403 B.n363 VSUBS 0.008476f
C404 B.n364 VSUBS 0.008476f
C405 B.n365 VSUBS 0.008476f
C406 B.n366 VSUBS 0.008476f
C407 B.n367 VSUBS 0.008476f
C408 B.n368 VSUBS 0.008476f
C409 B.n369 VSUBS 0.008476f
C410 B.n370 VSUBS 0.008476f
C411 B.n371 VSUBS 0.008476f
C412 B.n372 VSUBS 0.008476f
C413 B.n373 VSUBS 0.008476f
C414 B.n374 VSUBS 0.008476f
C415 B.n375 VSUBS 0.008476f
C416 B.n376 VSUBS 0.008476f
C417 B.n377 VSUBS 0.008476f
C418 B.n378 VSUBS 0.008476f
C419 B.n379 VSUBS 0.008476f
C420 B.n380 VSUBS 0.008476f
C421 B.n381 VSUBS 0.008476f
C422 B.n382 VSUBS 0.008476f
C423 B.n383 VSUBS 0.008476f
C424 B.n384 VSUBS 0.008476f
C425 B.n385 VSUBS 0.008476f
C426 B.n386 VSUBS 0.008476f
C427 B.n387 VSUBS 0.008476f
C428 B.n388 VSUBS 0.008476f
C429 B.n389 VSUBS 0.008476f
C430 B.n390 VSUBS 0.008476f
C431 B.n391 VSUBS 0.008476f
C432 B.n392 VSUBS 0.008476f
C433 B.n393 VSUBS 0.008476f
C434 B.n394 VSUBS 0.008476f
C435 B.n395 VSUBS 0.008476f
C436 B.n396 VSUBS 0.008476f
C437 B.n397 VSUBS 0.008476f
C438 B.n398 VSUBS 0.008476f
C439 B.n399 VSUBS 0.008476f
C440 B.n400 VSUBS 0.008476f
C441 B.n401 VSUBS 0.008476f
C442 B.n402 VSUBS 0.008476f
C443 B.n403 VSUBS 0.008476f
C444 B.n404 VSUBS 0.008476f
C445 B.n405 VSUBS 0.008476f
C446 B.n406 VSUBS 0.008476f
C447 B.n407 VSUBS 0.008476f
C448 B.n408 VSUBS 0.008476f
C449 B.n409 VSUBS 0.008476f
C450 B.n410 VSUBS 0.008476f
C451 B.n411 VSUBS 0.008476f
C452 B.n412 VSUBS 0.008476f
C453 B.n413 VSUBS 0.008476f
C454 B.n414 VSUBS 0.008476f
C455 B.n415 VSUBS 0.008476f
C456 B.n416 VSUBS 0.008476f
C457 B.n417 VSUBS 0.008476f
C458 B.n418 VSUBS 0.008476f
C459 B.n419 VSUBS 0.008476f
C460 B.n420 VSUBS 0.008476f
C461 B.n421 VSUBS 0.008476f
C462 B.n422 VSUBS 0.008476f
C463 B.n423 VSUBS 0.008476f
C464 B.n424 VSUBS 0.008476f
C465 B.n425 VSUBS 0.008476f
C466 B.n426 VSUBS 0.008476f
C467 B.n427 VSUBS 0.008476f
C468 B.n428 VSUBS 0.008476f
C469 B.n429 VSUBS 0.008476f
C470 B.n430 VSUBS 0.008476f
C471 B.n431 VSUBS 0.008476f
C472 B.n432 VSUBS 0.008476f
C473 B.n433 VSUBS 0.008476f
C474 B.n434 VSUBS 0.008476f
C475 B.n435 VSUBS 0.008476f
C476 B.n436 VSUBS 0.008476f
C477 B.n437 VSUBS 0.008476f
C478 B.n438 VSUBS 0.008476f
C479 B.n439 VSUBS 0.008476f
C480 B.n440 VSUBS 0.020847f
C481 B.n441 VSUBS 0.021533f
C482 B.n442 VSUBS 0.020626f
C483 B.n443 VSUBS 0.008476f
C484 B.n444 VSUBS 0.008476f
C485 B.n445 VSUBS 0.008476f
C486 B.n446 VSUBS 0.008476f
C487 B.n447 VSUBS 0.008476f
C488 B.n448 VSUBS 0.008476f
C489 B.n449 VSUBS 0.008476f
C490 B.n450 VSUBS 0.008476f
C491 B.n451 VSUBS 0.008476f
C492 B.n452 VSUBS 0.008476f
C493 B.n453 VSUBS 0.008476f
C494 B.n454 VSUBS 0.008476f
C495 B.n455 VSUBS 0.008476f
C496 B.n456 VSUBS 0.008476f
C497 B.n457 VSUBS 0.008476f
C498 B.n458 VSUBS 0.008476f
C499 B.n459 VSUBS 0.008476f
C500 B.n460 VSUBS 0.008476f
C501 B.n461 VSUBS 0.008476f
C502 B.n462 VSUBS 0.008476f
C503 B.n463 VSUBS 0.008476f
C504 B.n464 VSUBS 0.008476f
C505 B.n465 VSUBS 0.008476f
C506 B.n466 VSUBS 0.008476f
C507 B.n467 VSUBS 0.008476f
C508 B.n468 VSUBS 0.008476f
C509 B.n469 VSUBS 0.008476f
C510 B.n470 VSUBS 0.008476f
C511 B.n471 VSUBS 0.008476f
C512 B.n472 VSUBS 0.008476f
C513 B.n473 VSUBS 0.008476f
C514 B.n474 VSUBS 0.008476f
C515 B.n475 VSUBS 0.008476f
C516 B.n476 VSUBS 0.008476f
C517 B.n477 VSUBS 0.008476f
C518 B.n478 VSUBS 0.008476f
C519 B.n479 VSUBS 0.008476f
C520 B.n480 VSUBS 0.008476f
C521 B.n481 VSUBS 0.008476f
C522 B.n482 VSUBS 0.008476f
C523 B.n483 VSUBS 0.008476f
C524 B.n484 VSUBS 0.008476f
C525 B.n485 VSUBS 0.008476f
C526 B.n486 VSUBS 0.008476f
C527 B.n487 VSUBS 0.008476f
C528 B.n488 VSUBS 0.008476f
C529 B.n489 VSUBS 0.008476f
C530 B.n490 VSUBS 0.008476f
C531 B.n491 VSUBS 0.008476f
C532 B.n492 VSUBS 0.008476f
C533 B.n493 VSUBS 0.008476f
C534 B.n494 VSUBS 0.008476f
C535 B.n495 VSUBS 0.008476f
C536 B.n496 VSUBS 0.008476f
C537 B.n497 VSUBS 0.008476f
C538 B.n498 VSUBS 0.008476f
C539 B.n499 VSUBS 0.008476f
C540 B.n500 VSUBS 0.008476f
C541 B.n501 VSUBS 0.008476f
C542 B.n502 VSUBS 0.008476f
C543 B.n503 VSUBS 0.008476f
C544 B.n504 VSUBS 0.008476f
C545 B.n505 VSUBS 0.008476f
C546 B.n506 VSUBS 0.008476f
C547 B.n507 VSUBS 0.008476f
C548 B.n508 VSUBS 0.008476f
C549 B.n509 VSUBS 0.008476f
C550 B.n510 VSUBS 0.008476f
C551 B.n511 VSUBS 0.008476f
C552 B.n512 VSUBS 0.008476f
C553 B.n513 VSUBS 0.008476f
C554 B.n514 VSUBS 0.008476f
C555 B.n515 VSUBS 0.008476f
C556 B.n516 VSUBS 0.008476f
C557 B.n517 VSUBS 0.008476f
C558 B.n518 VSUBS 0.008476f
C559 B.n519 VSUBS 0.008476f
C560 B.n520 VSUBS 0.008476f
C561 B.n521 VSUBS 0.008476f
C562 B.n522 VSUBS 0.008476f
C563 B.n523 VSUBS 0.008476f
C564 B.n524 VSUBS 0.008476f
C565 B.n525 VSUBS 0.008476f
C566 B.n526 VSUBS 0.008476f
C567 B.n527 VSUBS 0.008476f
C568 B.n528 VSUBS 0.008476f
C569 B.n529 VSUBS 0.008476f
C570 B.n530 VSUBS 0.008476f
C571 B.n531 VSUBS 0.008476f
C572 B.n532 VSUBS 0.008476f
C573 B.n533 VSUBS 0.008476f
C574 B.n534 VSUBS 0.008476f
C575 B.n535 VSUBS 0.008476f
C576 B.n536 VSUBS 0.008476f
C577 B.n537 VSUBS 0.008476f
C578 B.n538 VSUBS 0.008476f
C579 B.n539 VSUBS 0.008476f
C580 B.n540 VSUBS 0.008476f
C581 B.n541 VSUBS 0.008476f
C582 B.n542 VSUBS 0.008476f
C583 B.n543 VSUBS 0.008476f
C584 B.n544 VSUBS 0.008476f
C585 B.n545 VSUBS 0.008476f
C586 B.n546 VSUBS 0.008476f
C587 B.n547 VSUBS 0.008476f
C588 B.n548 VSUBS 0.008476f
C589 B.n549 VSUBS 0.008476f
C590 B.n550 VSUBS 0.008476f
C591 B.n551 VSUBS 0.008476f
C592 B.n552 VSUBS 0.008476f
C593 B.n553 VSUBS 0.008476f
C594 B.n554 VSUBS 0.020626f
C595 B.n555 VSUBS 0.021754f
C596 B.n556 VSUBS 0.021754f
C597 B.n557 VSUBS 0.008476f
C598 B.n558 VSUBS 0.008476f
C599 B.n559 VSUBS 0.008476f
C600 B.n560 VSUBS 0.008476f
C601 B.n561 VSUBS 0.008476f
C602 B.n562 VSUBS 0.008476f
C603 B.n563 VSUBS 0.008476f
C604 B.n564 VSUBS 0.008476f
C605 B.n565 VSUBS 0.008476f
C606 B.n566 VSUBS 0.008476f
C607 B.n567 VSUBS 0.008476f
C608 B.n568 VSUBS 0.008476f
C609 B.n569 VSUBS 0.008476f
C610 B.n570 VSUBS 0.008476f
C611 B.n571 VSUBS 0.008476f
C612 B.n572 VSUBS 0.008476f
C613 B.n573 VSUBS 0.008476f
C614 B.n574 VSUBS 0.008476f
C615 B.n575 VSUBS 0.008476f
C616 B.n576 VSUBS 0.008476f
C617 B.n577 VSUBS 0.008476f
C618 B.n578 VSUBS 0.008476f
C619 B.n579 VSUBS 0.008476f
C620 B.n580 VSUBS 0.008476f
C621 B.n581 VSUBS 0.008476f
C622 B.n582 VSUBS 0.008476f
C623 B.n583 VSUBS 0.008476f
C624 B.n584 VSUBS 0.008476f
C625 B.n585 VSUBS 0.008476f
C626 B.n586 VSUBS 0.008476f
C627 B.n587 VSUBS 0.008476f
C628 B.n588 VSUBS 0.008476f
C629 B.n589 VSUBS 0.008476f
C630 B.n590 VSUBS 0.008476f
C631 B.n591 VSUBS 0.008476f
C632 B.n592 VSUBS 0.008476f
C633 B.n593 VSUBS 0.008476f
C634 B.n594 VSUBS 0.008476f
C635 B.n595 VSUBS 0.008476f
C636 B.n596 VSUBS 0.008476f
C637 B.n597 VSUBS 0.008476f
C638 B.n598 VSUBS 0.008476f
C639 B.n599 VSUBS 0.008476f
C640 B.n600 VSUBS 0.008476f
C641 B.n601 VSUBS 0.008476f
C642 B.n602 VSUBS 0.008476f
C643 B.n603 VSUBS 0.008476f
C644 B.n604 VSUBS 0.008476f
C645 B.n605 VSUBS 0.008476f
C646 B.n606 VSUBS 0.008476f
C647 B.n607 VSUBS 0.008476f
C648 B.n608 VSUBS 0.008476f
C649 B.n609 VSUBS 0.008476f
C650 B.n610 VSUBS 0.008476f
C651 B.n611 VSUBS 0.008476f
C652 B.n612 VSUBS 0.008476f
C653 B.n613 VSUBS 0.008476f
C654 B.n614 VSUBS 0.008476f
C655 B.n615 VSUBS 0.008476f
C656 B.n616 VSUBS 0.008476f
C657 B.n617 VSUBS 0.008476f
C658 B.n618 VSUBS 0.008476f
C659 B.n619 VSUBS 0.008476f
C660 B.n620 VSUBS 0.008476f
C661 B.n621 VSUBS 0.008476f
C662 B.n622 VSUBS 0.008476f
C663 B.n623 VSUBS 0.008476f
C664 B.n624 VSUBS 0.008476f
C665 B.n625 VSUBS 0.008476f
C666 B.n626 VSUBS 0.008476f
C667 B.n627 VSUBS 0.008476f
C668 B.n628 VSUBS 0.008476f
C669 B.n629 VSUBS 0.008476f
C670 B.n630 VSUBS 0.008476f
C671 B.n631 VSUBS 0.008476f
C672 B.n632 VSUBS 0.008476f
C673 B.n633 VSUBS 0.008476f
C674 B.n634 VSUBS 0.008476f
C675 B.n635 VSUBS 0.008476f
C676 B.n636 VSUBS 0.008476f
C677 B.n637 VSUBS 0.007977f
C678 B.n638 VSUBS 0.019638f
C679 B.n639 VSUBS 0.004737f
C680 B.n640 VSUBS 0.008476f
C681 B.n641 VSUBS 0.008476f
C682 B.n642 VSUBS 0.008476f
C683 B.n643 VSUBS 0.008476f
C684 B.n644 VSUBS 0.008476f
C685 B.n645 VSUBS 0.008476f
C686 B.n646 VSUBS 0.008476f
C687 B.n647 VSUBS 0.008476f
C688 B.n648 VSUBS 0.008476f
C689 B.n649 VSUBS 0.008476f
C690 B.n650 VSUBS 0.008476f
C691 B.n651 VSUBS 0.008476f
C692 B.n652 VSUBS 0.004737f
C693 B.n653 VSUBS 0.008476f
C694 B.n654 VSUBS 0.008476f
C695 B.n655 VSUBS 0.007977f
C696 B.n656 VSUBS 0.008476f
C697 B.n657 VSUBS 0.008476f
C698 B.n658 VSUBS 0.008476f
C699 B.n659 VSUBS 0.008476f
C700 B.n660 VSUBS 0.008476f
C701 B.n661 VSUBS 0.008476f
C702 B.n662 VSUBS 0.008476f
C703 B.n663 VSUBS 0.008476f
C704 B.n664 VSUBS 0.008476f
C705 B.n665 VSUBS 0.008476f
C706 B.n666 VSUBS 0.008476f
C707 B.n667 VSUBS 0.008476f
C708 B.n668 VSUBS 0.008476f
C709 B.n669 VSUBS 0.008476f
C710 B.n670 VSUBS 0.008476f
C711 B.n671 VSUBS 0.008476f
C712 B.n672 VSUBS 0.008476f
C713 B.n673 VSUBS 0.008476f
C714 B.n674 VSUBS 0.008476f
C715 B.n675 VSUBS 0.008476f
C716 B.n676 VSUBS 0.008476f
C717 B.n677 VSUBS 0.008476f
C718 B.n678 VSUBS 0.008476f
C719 B.n679 VSUBS 0.008476f
C720 B.n680 VSUBS 0.008476f
C721 B.n681 VSUBS 0.008476f
C722 B.n682 VSUBS 0.008476f
C723 B.n683 VSUBS 0.008476f
C724 B.n684 VSUBS 0.008476f
C725 B.n685 VSUBS 0.008476f
C726 B.n686 VSUBS 0.008476f
C727 B.n687 VSUBS 0.008476f
C728 B.n688 VSUBS 0.008476f
C729 B.n689 VSUBS 0.008476f
C730 B.n690 VSUBS 0.008476f
C731 B.n691 VSUBS 0.008476f
C732 B.n692 VSUBS 0.008476f
C733 B.n693 VSUBS 0.008476f
C734 B.n694 VSUBS 0.008476f
C735 B.n695 VSUBS 0.008476f
C736 B.n696 VSUBS 0.008476f
C737 B.n697 VSUBS 0.008476f
C738 B.n698 VSUBS 0.008476f
C739 B.n699 VSUBS 0.008476f
C740 B.n700 VSUBS 0.008476f
C741 B.n701 VSUBS 0.008476f
C742 B.n702 VSUBS 0.008476f
C743 B.n703 VSUBS 0.008476f
C744 B.n704 VSUBS 0.008476f
C745 B.n705 VSUBS 0.008476f
C746 B.n706 VSUBS 0.008476f
C747 B.n707 VSUBS 0.008476f
C748 B.n708 VSUBS 0.008476f
C749 B.n709 VSUBS 0.008476f
C750 B.n710 VSUBS 0.008476f
C751 B.n711 VSUBS 0.008476f
C752 B.n712 VSUBS 0.008476f
C753 B.n713 VSUBS 0.008476f
C754 B.n714 VSUBS 0.008476f
C755 B.n715 VSUBS 0.008476f
C756 B.n716 VSUBS 0.008476f
C757 B.n717 VSUBS 0.008476f
C758 B.n718 VSUBS 0.008476f
C759 B.n719 VSUBS 0.008476f
C760 B.n720 VSUBS 0.008476f
C761 B.n721 VSUBS 0.008476f
C762 B.n722 VSUBS 0.008476f
C763 B.n723 VSUBS 0.008476f
C764 B.n724 VSUBS 0.008476f
C765 B.n725 VSUBS 0.008476f
C766 B.n726 VSUBS 0.008476f
C767 B.n727 VSUBS 0.008476f
C768 B.n728 VSUBS 0.008476f
C769 B.n729 VSUBS 0.008476f
C770 B.n730 VSUBS 0.008476f
C771 B.n731 VSUBS 0.008476f
C772 B.n732 VSUBS 0.008476f
C773 B.n733 VSUBS 0.008476f
C774 B.n734 VSUBS 0.008476f
C775 B.n735 VSUBS 0.021754f
C776 B.n736 VSUBS 0.021754f
C777 B.n737 VSUBS 0.020626f
C778 B.n738 VSUBS 0.008476f
C779 B.n739 VSUBS 0.008476f
C780 B.n740 VSUBS 0.008476f
C781 B.n741 VSUBS 0.008476f
C782 B.n742 VSUBS 0.008476f
C783 B.n743 VSUBS 0.008476f
C784 B.n744 VSUBS 0.008476f
C785 B.n745 VSUBS 0.008476f
C786 B.n746 VSUBS 0.008476f
C787 B.n747 VSUBS 0.008476f
C788 B.n748 VSUBS 0.008476f
C789 B.n749 VSUBS 0.008476f
C790 B.n750 VSUBS 0.008476f
C791 B.n751 VSUBS 0.008476f
C792 B.n752 VSUBS 0.008476f
C793 B.n753 VSUBS 0.008476f
C794 B.n754 VSUBS 0.008476f
C795 B.n755 VSUBS 0.008476f
C796 B.n756 VSUBS 0.008476f
C797 B.n757 VSUBS 0.008476f
C798 B.n758 VSUBS 0.008476f
C799 B.n759 VSUBS 0.008476f
C800 B.n760 VSUBS 0.008476f
C801 B.n761 VSUBS 0.008476f
C802 B.n762 VSUBS 0.008476f
C803 B.n763 VSUBS 0.008476f
C804 B.n764 VSUBS 0.008476f
C805 B.n765 VSUBS 0.008476f
C806 B.n766 VSUBS 0.008476f
C807 B.n767 VSUBS 0.008476f
C808 B.n768 VSUBS 0.008476f
C809 B.n769 VSUBS 0.008476f
C810 B.n770 VSUBS 0.008476f
C811 B.n771 VSUBS 0.008476f
C812 B.n772 VSUBS 0.008476f
C813 B.n773 VSUBS 0.008476f
C814 B.n774 VSUBS 0.008476f
C815 B.n775 VSUBS 0.008476f
C816 B.n776 VSUBS 0.008476f
C817 B.n777 VSUBS 0.008476f
C818 B.n778 VSUBS 0.008476f
C819 B.n779 VSUBS 0.008476f
C820 B.n780 VSUBS 0.008476f
C821 B.n781 VSUBS 0.008476f
C822 B.n782 VSUBS 0.008476f
C823 B.n783 VSUBS 0.008476f
C824 B.n784 VSUBS 0.008476f
C825 B.n785 VSUBS 0.008476f
C826 B.n786 VSUBS 0.008476f
C827 B.n787 VSUBS 0.008476f
C828 B.n788 VSUBS 0.008476f
C829 B.n789 VSUBS 0.008476f
C830 B.n790 VSUBS 0.008476f
C831 B.n791 VSUBS 0.011061f
C832 B.n792 VSUBS 0.011783f
C833 B.n793 VSUBS 0.023431f
C834 VDD2.t4 VSUBS 3.81309f
C835 VDD2.t2 VSUBS 0.353596f
C836 VDD2.t3 VSUBS 0.353596f
C837 VDD2.n0 VSUBS 2.92626f
C838 VDD2.n1 VSUBS 1.38106f
C839 VDD2.t8 VSUBS 0.353596f
C840 VDD2.t9 VSUBS 0.353596f
C841 VDD2.n2 VSUBS 2.93638f
C842 VDD2.n3 VSUBS 3.00959f
C843 VDD2.t7 VSUBS 3.7993f
C844 VDD2.n4 VSUBS 3.52725f
C845 VDD2.t0 VSUBS 0.353596f
C846 VDD2.t5 VSUBS 0.353596f
C847 VDD2.n5 VSUBS 2.92627f
C848 VDD2.n6 VSUBS 0.668448f
C849 VDD2.t1 VSUBS 0.353596f
C850 VDD2.t6 VSUBS 0.353596f
C851 VDD2.n7 VSUBS 2.93633f
C852 VN.n0 VSUBS 0.049581f
C853 VN.t1 VSUBS 2.29374f
C854 VN.n1 VSUBS 0.814388f
C855 VN.n2 VSUBS 0.037157f
C856 VN.t6 VSUBS 2.29374f
C857 VN.n3 VSUBS 0.849449f
C858 VN.n4 VSUBS 0.037157f
C859 VN.t7 VSUBS 2.29374f
C860 VN.n5 VSUBS 0.860908f
C861 VN.t5 VSUBS 2.4182f
C862 VN.n6 VSUBS 0.884644f
C863 VN.n7 VSUBS 0.197073f
C864 VN.n8 VSUBS 0.04802f
C865 VN.n9 VSUBS 0.044364f
C866 VN.n10 VSUBS 0.063469f
C867 VN.n11 VSUBS 0.037157f
C868 VN.n12 VSUBS 0.037157f
C869 VN.n13 VSUBS 0.037157f
C870 VN.n14 VSUBS 0.063469f
C871 VN.n15 VSUBS 0.044364f
C872 VN.n16 VSUBS 0.04802f
C873 VN.n17 VSUBS 0.037157f
C874 VN.n18 VSUBS 0.037157f
C875 VN.n19 VSUBS 0.062186f
C876 VN.n20 VSUBS 0.020866f
C877 VN.t0 VSUBS 2.37058f
C878 VN.n21 VSUBS 0.893955f
C879 VN.n22 VSUBS 0.034799f
C880 VN.n23 VSUBS 0.049581f
C881 VN.t9 VSUBS 2.29374f
C882 VN.n24 VSUBS 0.814388f
C883 VN.n25 VSUBS 0.037157f
C884 VN.t4 VSUBS 2.29374f
C885 VN.n26 VSUBS 0.849449f
C886 VN.n27 VSUBS 0.037157f
C887 VN.t8 VSUBS 2.29374f
C888 VN.n28 VSUBS 0.860908f
C889 VN.t3 VSUBS 2.4182f
C890 VN.n29 VSUBS 0.884644f
C891 VN.n30 VSUBS 0.197073f
C892 VN.n31 VSUBS 0.04802f
C893 VN.n32 VSUBS 0.044364f
C894 VN.n33 VSUBS 0.063469f
C895 VN.n34 VSUBS 0.037157f
C896 VN.n35 VSUBS 0.037157f
C897 VN.n36 VSUBS 0.037157f
C898 VN.n37 VSUBS 0.063469f
C899 VN.n38 VSUBS 0.044364f
C900 VN.n39 VSUBS 0.04802f
C901 VN.n40 VSUBS 0.037157f
C902 VN.n41 VSUBS 0.037157f
C903 VN.n42 VSUBS 0.062186f
C904 VN.n43 VSUBS 0.020866f
C905 VN.t2 VSUBS 2.37058f
C906 VN.n44 VSUBS 0.893955f
C907 VN.n45 VSUBS 2.05596f
C908 VTAIL.t5 VSUBS 0.359052f
C909 VTAIL.t0 VSUBS 0.359052f
C910 VTAIL.n0 VSUBS 2.82235f
C911 VTAIL.n1 VSUBS 0.832043f
C912 VTAIL.t13 VSUBS 3.68755f
C913 VTAIL.n2 VSUBS 0.972796f
C914 VTAIL.t16 VSUBS 0.359052f
C915 VTAIL.t10 VSUBS 0.359052f
C916 VTAIL.n3 VSUBS 2.82235f
C917 VTAIL.n4 VSUBS 0.881126f
C918 VTAIL.t17 VSUBS 0.359052f
C919 VTAIL.t19 VSUBS 0.359052f
C920 VTAIL.n5 VSUBS 2.82235f
C921 VTAIL.n6 VSUBS 2.64129f
C922 VTAIL.t2 VSUBS 0.359052f
C923 VTAIL.t6 VSUBS 0.359052f
C924 VTAIL.n7 VSUBS 2.82236f
C925 VTAIL.n8 VSUBS 2.64128f
C926 VTAIL.t1 VSUBS 0.359052f
C927 VTAIL.t3 VSUBS 0.359052f
C928 VTAIL.n9 VSUBS 2.82236f
C929 VTAIL.n10 VSUBS 0.88112f
C930 VTAIL.t7 VSUBS 3.68756f
C931 VTAIL.n11 VSUBS 0.97279f
C932 VTAIL.t18 VSUBS 0.359052f
C933 VTAIL.t14 VSUBS 0.359052f
C934 VTAIL.n12 VSUBS 2.82236f
C935 VTAIL.n13 VSUBS 0.858758f
C936 VTAIL.t12 VSUBS 0.359052f
C937 VTAIL.t15 VSUBS 0.359052f
C938 VTAIL.n14 VSUBS 2.82236f
C939 VTAIL.n15 VSUBS 0.88112f
C940 VTAIL.t11 VSUBS 3.68755f
C941 VTAIL.n16 VSUBS 2.62797f
C942 VTAIL.t9 VSUBS 3.68755f
C943 VTAIL.n17 VSUBS 2.62797f
C944 VTAIL.t4 VSUBS 0.359052f
C945 VTAIL.t8 VSUBS 0.359052f
C946 VTAIL.n18 VSUBS 2.82235f
C947 VTAIL.n19 VSUBS 0.780497f
C948 VDD1.t2 VSUBS 3.81319f
C949 VDD1.t6 VSUBS 0.353605f
C950 VDD1.t8 VSUBS 0.353605f
C951 VDD1.n0 VSUBS 2.92633f
C952 VDD1.n1 VSUBS 1.38888f
C953 VDD1.t5 VSUBS 3.81318f
C954 VDD1.t3 VSUBS 0.353605f
C955 VDD1.t4 VSUBS 0.353605f
C956 VDD1.n2 VSUBS 2.92633f
C957 VDD1.n3 VSUBS 1.38109f
C958 VDD1.t0 VSUBS 0.353605f
C959 VDD1.t9 VSUBS 0.353605f
C960 VDD1.n4 VSUBS 2.93644f
C961 VDD1.n5 VSUBS 3.11139f
C962 VDD1.t7 VSUBS 0.353605f
C963 VDD1.t1 VSUBS 0.353605f
C964 VDD1.n6 VSUBS 2.92632f
C965 VDD1.n7 VSUBS 3.52258f
C966 VP.n0 VSUBS 0.050566f
C967 VP.t9 VSUBS 2.33932f
C968 VP.n1 VSUBS 0.830574f
C969 VP.n2 VSUBS 0.037895f
C970 VP.t3 VSUBS 2.33932f
C971 VP.n3 VSUBS 0.866332f
C972 VP.n4 VSUBS 0.037895f
C973 VP.t0 VSUBS 2.33932f
C974 VP.n5 VSUBS 0.830574f
C975 VP.n6 VSUBS 0.050566f
C976 VP.n7 VSUBS 0.050566f
C977 VP.t8 VSUBS 2.4177f
C978 VP.t4 VSUBS 2.33932f
C979 VP.n8 VSUBS 0.830574f
C980 VP.n9 VSUBS 0.037895f
C981 VP.t7 VSUBS 2.33932f
C982 VP.n10 VSUBS 0.866332f
C983 VP.n11 VSUBS 0.037895f
C984 VP.t5 VSUBS 2.33932f
C985 VP.n12 VSUBS 0.878018f
C986 VP.t1 VSUBS 2.46626f
C987 VP.n13 VSUBS 0.902226f
C988 VP.n14 VSUBS 0.20099f
C989 VP.n15 VSUBS 0.048974f
C990 VP.n16 VSUBS 0.045246f
C991 VP.n17 VSUBS 0.064731f
C992 VP.n18 VSUBS 0.037895f
C993 VP.n19 VSUBS 0.037895f
C994 VP.n20 VSUBS 0.037895f
C995 VP.n21 VSUBS 0.064731f
C996 VP.n22 VSUBS 0.045246f
C997 VP.n23 VSUBS 0.048974f
C998 VP.n24 VSUBS 0.037895f
C999 VP.n25 VSUBS 0.037895f
C1000 VP.n26 VSUBS 0.063422f
C1001 VP.n27 VSUBS 0.021281f
C1002 VP.n28 VSUBS 0.911722f
C1003 VP.n29 VSUBS 2.07616f
C1004 VP.n30 VSUBS 2.10338f
C1005 VP.t2 VSUBS 2.4177f
C1006 VP.n31 VSUBS 0.911722f
C1007 VP.n32 VSUBS 0.021281f
C1008 VP.n33 VSUBS 0.063422f
C1009 VP.n34 VSUBS 0.037895f
C1010 VP.n35 VSUBS 0.037895f
C1011 VP.n36 VSUBS 0.048974f
C1012 VP.n37 VSUBS 0.045246f
C1013 VP.n38 VSUBS 0.064731f
C1014 VP.n39 VSUBS 0.037895f
C1015 VP.n40 VSUBS 0.037895f
C1016 VP.n41 VSUBS 0.037895f
C1017 VP.n42 VSUBS 0.064731f
C1018 VP.n43 VSUBS 0.045246f
C1019 VP.n44 VSUBS 0.048974f
C1020 VP.n45 VSUBS 0.037895f
C1021 VP.n46 VSUBS 0.037895f
C1022 VP.n47 VSUBS 0.063422f
C1023 VP.n48 VSUBS 0.021281f
C1024 VP.t6 VSUBS 2.4177f
C1025 VP.n49 VSUBS 0.911722f
C1026 VP.n50 VSUBS 0.03549f
.ends

