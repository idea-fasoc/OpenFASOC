* NGSPICE file created from diff_pair_sample_1525.ext - technology: sky130A

.subckt diff_pair_sample_1525 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t13 w_n1820_n3870# sky130_fd_pr__pfet_01v8 ad=2.39415 pd=14.84 as=5.6589 ps=29.8 w=14.51 l=0.52
X1 VTAIL.t1 VP.t0 VDD1.t7 w_n1820_n3870# sky130_fd_pr__pfet_01v8 ad=5.6589 pd=29.8 as=2.39415 ps=14.84 w=14.51 l=0.52
X2 VTAIL.t0 VP.t1 VDD1.t6 w_n1820_n3870# sky130_fd_pr__pfet_01v8 ad=2.39415 pd=14.84 as=2.39415 ps=14.84 w=14.51 l=0.52
X3 VDD2.t6 VN.t1 VTAIL.t11 w_n1820_n3870# sky130_fd_pr__pfet_01v8 ad=2.39415 pd=14.84 as=5.6589 ps=29.8 w=14.51 l=0.52
X4 VDD2.t5 VN.t2 VTAIL.t9 w_n1820_n3870# sky130_fd_pr__pfet_01v8 ad=2.39415 pd=14.84 as=2.39415 ps=14.84 w=14.51 l=0.52
X5 B.t11 B.t9 B.t10 w_n1820_n3870# sky130_fd_pr__pfet_01v8 ad=5.6589 pd=29.8 as=0 ps=0 w=14.51 l=0.52
X6 B.t8 B.t6 B.t7 w_n1820_n3870# sky130_fd_pr__pfet_01v8 ad=5.6589 pd=29.8 as=0 ps=0 w=14.51 l=0.52
X7 VDD2.t4 VN.t3 VTAIL.t14 w_n1820_n3870# sky130_fd_pr__pfet_01v8 ad=2.39415 pd=14.84 as=2.39415 ps=14.84 w=14.51 l=0.52
X8 B.t5 B.t3 B.t4 w_n1820_n3870# sky130_fd_pr__pfet_01v8 ad=5.6589 pd=29.8 as=0 ps=0 w=14.51 l=0.52
X9 VTAIL.t8 VN.t4 VDD2.t3 w_n1820_n3870# sky130_fd_pr__pfet_01v8 ad=2.39415 pd=14.84 as=2.39415 ps=14.84 w=14.51 l=0.52
X10 B.t2 B.t0 B.t1 w_n1820_n3870# sky130_fd_pr__pfet_01v8 ad=5.6589 pd=29.8 as=0 ps=0 w=14.51 l=0.52
X11 VTAIL.t15 VN.t5 VDD2.t2 w_n1820_n3870# sky130_fd_pr__pfet_01v8 ad=2.39415 pd=14.84 as=2.39415 ps=14.84 w=14.51 l=0.52
X12 VDD1.t5 VP.t2 VTAIL.t2 w_n1820_n3870# sky130_fd_pr__pfet_01v8 ad=2.39415 pd=14.84 as=2.39415 ps=14.84 w=14.51 l=0.52
X13 VTAIL.t12 VN.t6 VDD2.t1 w_n1820_n3870# sky130_fd_pr__pfet_01v8 ad=5.6589 pd=29.8 as=2.39415 ps=14.84 w=14.51 l=0.52
X14 VTAIL.t3 VP.t3 VDD1.t4 w_n1820_n3870# sky130_fd_pr__pfet_01v8 ad=5.6589 pd=29.8 as=2.39415 ps=14.84 w=14.51 l=0.52
X15 VTAIL.t5 VP.t4 VDD1.t3 w_n1820_n3870# sky130_fd_pr__pfet_01v8 ad=2.39415 pd=14.84 as=2.39415 ps=14.84 w=14.51 l=0.52
X16 VTAIL.t10 VN.t7 VDD2.t0 w_n1820_n3870# sky130_fd_pr__pfet_01v8 ad=5.6589 pd=29.8 as=2.39415 ps=14.84 w=14.51 l=0.52
X17 VDD1.t2 VP.t5 VTAIL.t7 w_n1820_n3870# sky130_fd_pr__pfet_01v8 ad=2.39415 pd=14.84 as=5.6589 ps=29.8 w=14.51 l=0.52
X18 VDD1.t1 VP.t6 VTAIL.t4 w_n1820_n3870# sky130_fd_pr__pfet_01v8 ad=2.39415 pd=14.84 as=2.39415 ps=14.84 w=14.51 l=0.52
X19 VDD1.t0 VP.t7 VTAIL.t6 w_n1820_n3870# sky130_fd_pr__pfet_01v8 ad=2.39415 pd=14.84 as=5.6589 ps=29.8 w=14.51 l=0.52
R0 VN.n2 VN.t7 770.828
R1 VN.n10 VN.t1 770.828
R2 VN.n6 VN.t0 750.682
R3 VN.n14 VN.t6 750.682
R4 VN.n1 VN.t2 748.49
R5 VN.n5 VN.t5 748.49
R6 VN.n9 VN.t4 748.49
R7 VN.n13 VN.t3 748.49
R8 VN.n7 VN.n6 161.3
R9 VN.n15 VN.n14 161.3
R10 VN.n13 VN.n8 161.3
R11 VN.n12 VN.n11 161.3
R12 VN.n5 VN.n0 161.3
R13 VN.n4 VN.n3 161.3
R14 VN.n11 VN.n10 70.8204
R15 VN.n3 VN.n2 70.8204
R16 VN.n6 VN.n5 46.0096
R17 VN.n14 VN.n13 46.0096
R18 VN VN.n15 43.563
R19 VN.n4 VN.n1 24.1005
R20 VN.n5 VN.n4 24.1005
R21 VN.n13 VN.n12 24.1005
R22 VN.n12 VN.n9 24.1005
R23 VN.n10 VN.n9 20.1238
R24 VN.n2 VN.n1 20.1238
R25 VN.n15 VN.n8 0.189894
R26 VN.n11 VN.n8 0.189894
R27 VN.n3 VN.n0 0.189894
R28 VN.n7 VN.n0 0.189894
R29 VN VN.n7 0.0516364
R30 VTAIL.n11 VTAIL.t3 61.0645
R31 VTAIL.n10 VTAIL.t11 61.0645
R32 VTAIL.n7 VTAIL.t12 61.0645
R33 VTAIL.n15 VTAIL.t13 61.0644
R34 VTAIL.n2 VTAIL.t10 61.0644
R35 VTAIL.n3 VTAIL.t7 61.0644
R36 VTAIL.n6 VTAIL.t1 61.0644
R37 VTAIL.n14 VTAIL.t6 61.0644
R38 VTAIL.n13 VTAIL.n12 58.8244
R39 VTAIL.n9 VTAIL.n8 58.8244
R40 VTAIL.n1 VTAIL.n0 58.8241
R41 VTAIL.n5 VTAIL.n4 58.8241
R42 VTAIL.n15 VTAIL.n14 25.6083
R43 VTAIL.n7 VTAIL.n6 25.6083
R44 VTAIL.n0 VTAIL.t9 2.24068
R45 VTAIL.n0 VTAIL.t15 2.24068
R46 VTAIL.n4 VTAIL.t2 2.24068
R47 VTAIL.n4 VTAIL.t0 2.24068
R48 VTAIL.n12 VTAIL.t4 2.24068
R49 VTAIL.n12 VTAIL.t5 2.24068
R50 VTAIL.n8 VTAIL.t14 2.24068
R51 VTAIL.n8 VTAIL.t8 2.24068
R52 VTAIL.n9 VTAIL.n7 0.733259
R53 VTAIL.n10 VTAIL.n9 0.733259
R54 VTAIL.n13 VTAIL.n11 0.733259
R55 VTAIL.n14 VTAIL.n13 0.733259
R56 VTAIL.n6 VTAIL.n5 0.733259
R57 VTAIL.n5 VTAIL.n3 0.733259
R58 VTAIL.n2 VTAIL.n1 0.733259
R59 VTAIL VTAIL.n15 0.675069
R60 VTAIL.n11 VTAIL.n10 0.470328
R61 VTAIL.n3 VTAIL.n2 0.470328
R62 VTAIL VTAIL.n1 0.0586897
R63 VDD2.n2 VDD2.n1 75.814
R64 VDD2.n2 VDD2.n0 75.814
R65 VDD2 VDD2.n5 75.8112
R66 VDD2.n4 VDD2.n3 75.5032
R67 VDD2.n4 VDD2.n2 39.5213
R68 VDD2.n5 VDD2.t3 2.24068
R69 VDD2.n5 VDD2.t6 2.24068
R70 VDD2.n3 VDD2.t1 2.24068
R71 VDD2.n3 VDD2.t4 2.24068
R72 VDD2.n1 VDD2.t2 2.24068
R73 VDD2.n1 VDD2.t7 2.24068
R74 VDD2.n0 VDD2.t0 2.24068
R75 VDD2.n0 VDD2.t5 2.24068
R76 VDD2 VDD2.n4 0.425069
R77 VP.n4 VP.t3 770.828
R78 VP.n16 VP.t5 750.682
R79 VP.n10 VP.t0 750.682
R80 VP.n8 VP.t7 750.682
R81 VP.n1 VP.t2 748.49
R82 VP.n15 VP.t1 748.49
R83 VP.n7 VP.t4 748.49
R84 VP.n3 VP.t6 748.49
R85 VP.n17 VP.n16 161.3
R86 VP.n6 VP.n5 161.3
R87 VP.n7 VP.n2 161.3
R88 VP.n9 VP.n8 161.3
R89 VP.n15 VP.n0 161.3
R90 VP.n14 VP.n13 161.3
R91 VP.n12 VP.n1 161.3
R92 VP.n11 VP.n10 161.3
R93 VP.n5 VP.n4 70.8204
R94 VP.n10 VP.n1 46.0096
R95 VP.n16 VP.n15 46.0096
R96 VP.n8 VP.n7 46.0096
R97 VP.n11 VP.n9 43.1823
R98 VP.n14 VP.n1 24.1005
R99 VP.n15 VP.n14 24.1005
R100 VP.n6 VP.n3 24.1005
R101 VP.n7 VP.n6 24.1005
R102 VP.n4 VP.n3 20.1238
R103 VP.n5 VP.n2 0.189894
R104 VP.n9 VP.n2 0.189894
R105 VP.n12 VP.n11 0.189894
R106 VP.n13 VP.n12 0.189894
R107 VP.n13 VP.n0 0.189894
R108 VP.n17 VP.n0 0.189894
R109 VP VP.n17 0.0516364
R110 VDD1 VDD1.n0 75.9278
R111 VDD1.n3 VDD1.n2 75.814
R112 VDD1.n3 VDD1.n1 75.814
R113 VDD1.n5 VDD1.n4 75.503
R114 VDD1.n5 VDD1.n3 40.1043
R115 VDD1.n4 VDD1.t3 2.24068
R116 VDD1.n4 VDD1.t0 2.24068
R117 VDD1.n0 VDD1.t4 2.24068
R118 VDD1.n0 VDD1.t1 2.24068
R119 VDD1.n2 VDD1.t6 2.24068
R120 VDD1.n2 VDD1.t2 2.24068
R121 VDD1.n1 VDD1.t7 2.24068
R122 VDD1.n1 VDD1.t5 2.24068
R123 VDD1 VDD1.n5 0.30869
R124 B.n258 B.t3 878.428
R125 B.n117 B.t0 878.428
R126 B.n45 B.t9 878.428
R127 B.n38 B.t6 878.428
R128 B.n351 B.n92 585
R129 B.n350 B.n349 585
R130 B.n348 B.n93 585
R131 B.n347 B.n346 585
R132 B.n345 B.n94 585
R133 B.n344 B.n343 585
R134 B.n342 B.n95 585
R135 B.n341 B.n340 585
R136 B.n339 B.n96 585
R137 B.n338 B.n337 585
R138 B.n336 B.n97 585
R139 B.n335 B.n334 585
R140 B.n333 B.n98 585
R141 B.n332 B.n331 585
R142 B.n330 B.n99 585
R143 B.n329 B.n328 585
R144 B.n327 B.n100 585
R145 B.n326 B.n325 585
R146 B.n324 B.n101 585
R147 B.n323 B.n322 585
R148 B.n321 B.n102 585
R149 B.n320 B.n319 585
R150 B.n318 B.n103 585
R151 B.n317 B.n316 585
R152 B.n315 B.n104 585
R153 B.n314 B.n313 585
R154 B.n312 B.n105 585
R155 B.n311 B.n310 585
R156 B.n309 B.n106 585
R157 B.n308 B.n307 585
R158 B.n306 B.n107 585
R159 B.n305 B.n304 585
R160 B.n303 B.n108 585
R161 B.n302 B.n301 585
R162 B.n300 B.n109 585
R163 B.n299 B.n298 585
R164 B.n297 B.n110 585
R165 B.n296 B.n295 585
R166 B.n294 B.n111 585
R167 B.n293 B.n292 585
R168 B.n291 B.n112 585
R169 B.n290 B.n289 585
R170 B.n288 B.n113 585
R171 B.n287 B.n286 585
R172 B.n285 B.n114 585
R173 B.n284 B.n283 585
R174 B.n282 B.n115 585
R175 B.n281 B.n280 585
R176 B.n279 B.n116 585
R177 B.n277 B.n276 585
R178 B.n275 B.n119 585
R179 B.n274 B.n273 585
R180 B.n272 B.n120 585
R181 B.n271 B.n270 585
R182 B.n269 B.n121 585
R183 B.n268 B.n267 585
R184 B.n266 B.n122 585
R185 B.n265 B.n264 585
R186 B.n263 B.n123 585
R187 B.n262 B.n261 585
R188 B.n257 B.n124 585
R189 B.n256 B.n255 585
R190 B.n254 B.n125 585
R191 B.n253 B.n252 585
R192 B.n251 B.n126 585
R193 B.n250 B.n249 585
R194 B.n248 B.n127 585
R195 B.n247 B.n246 585
R196 B.n245 B.n128 585
R197 B.n244 B.n243 585
R198 B.n242 B.n129 585
R199 B.n241 B.n240 585
R200 B.n239 B.n130 585
R201 B.n238 B.n237 585
R202 B.n236 B.n131 585
R203 B.n235 B.n234 585
R204 B.n233 B.n132 585
R205 B.n232 B.n231 585
R206 B.n230 B.n133 585
R207 B.n229 B.n228 585
R208 B.n227 B.n134 585
R209 B.n226 B.n225 585
R210 B.n224 B.n135 585
R211 B.n223 B.n222 585
R212 B.n221 B.n136 585
R213 B.n220 B.n219 585
R214 B.n218 B.n137 585
R215 B.n217 B.n216 585
R216 B.n215 B.n138 585
R217 B.n214 B.n213 585
R218 B.n212 B.n139 585
R219 B.n211 B.n210 585
R220 B.n209 B.n140 585
R221 B.n208 B.n207 585
R222 B.n206 B.n141 585
R223 B.n205 B.n204 585
R224 B.n203 B.n142 585
R225 B.n202 B.n201 585
R226 B.n200 B.n143 585
R227 B.n199 B.n198 585
R228 B.n197 B.n144 585
R229 B.n196 B.n195 585
R230 B.n194 B.n145 585
R231 B.n193 B.n192 585
R232 B.n191 B.n146 585
R233 B.n190 B.n189 585
R234 B.n188 B.n147 585
R235 B.n187 B.n186 585
R236 B.n353 B.n352 585
R237 B.n354 B.n91 585
R238 B.n356 B.n355 585
R239 B.n357 B.n90 585
R240 B.n359 B.n358 585
R241 B.n360 B.n89 585
R242 B.n362 B.n361 585
R243 B.n363 B.n88 585
R244 B.n365 B.n364 585
R245 B.n366 B.n87 585
R246 B.n368 B.n367 585
R247 B.n369 B.n86 585
R248 B.n371 B.n370 585
R249 B.n372 B.n85 585
R250 B.n374 B.n373 585
R251 B.n375 B.n84 585
R252 B.n377 B.n376 585
R253 B.n378 B.n83 585
R254 B.n380 B.n379 585
R255 B.n381 B.n82 585
R256 B.n383 B.n382 585
R257 B.n384 B.n81 585
R258 B.n386 B.n385 585
R259 B.n387 B.n80 585
R260 B.n389 B.n388 585
R261 B.n390 B.n79 585
R262 B.n392 B.n391 585
R263 B.n393 B.n78 585
R264 B.n395 B.n394 585
R265 B.n396 B.n77 585
R266 B.n398 B.n397 585
R267 B.n399 B.n76 585
R268 B.n401 B.n400 585
R269 B.n402 B.n75 585
R270 B.n404 B.n403 585
R271 B.n405 B.n74 585
R272 B.n407 B.n406 585
R273 B.n408 B.n73 585
R274 B.n410 B.n409 585
R275 B.n411 B.n72 585
R276 B.n413 B.n412 585
R277 B.n414 B.n71 585
R278 B.n577 B.n12 585
R279 B.n576 B.n575 585
R280 B.n574 B.n13 585
R281 B.n573 B.n572 585
R282 B.n571 B.n14 585
R283 B.n570 B.n569 585
R284 B.n568 B.n15 585
R285 B.n567 B.n566 585
R286 B.n565 B.n16 585
R287 B.n564 B.n563 585
R288 B.n562 B.n17 585
R289 B.n561 B.n560 585
R290 B.n559 B.n18 585
R291 B.n558 B.n557 585
R292 B.n556 B.n19 585
R293 B.n555 B.n554 585
R294 B.n553 B.n20 585
R295 B.n552 B.n551 585
R296 B.n550 B.n21 585
R297 B.n549 B.n548 585
R298 B.n547 B.n22 585
R299 B.n546 B.n545 585
R300 B.n544 B.n23 585
R301 B.n543 B.n542 585
R302 B.n541 B.n24 585
R303 B.n540 B.n539 585
R304 B.n538 B.n25 585
R305 B.n537 B.n536 585
R306 B.n535 B.n26 585
R307 B.n534 B.n533 585
R308 B.n532 B.n27 585
R309 B.n531 B.n530 585
R310 B.n529 B.n28 585
R311 B.n528 B.n527 585
R312 B.n526 B.n29 585
R313 B.n525 B.n524 585
R314 B.n523 B.n30 585
R315 B.n522 B.n521 585
R316 B.n520 B.n31 585
R317 B.n519 B.n518 585
R318 B.n517 B.n32 585
R319 B.n516 B.n515 585
R320 B.n514 B.n33 585
R321 B.n513 B.n512 585
R322 B.n511 B.n34 585
R323 B.n510 B.n509 585
R324 B.n508 B.n35 585
R325 B.n507 B.n506 585
R326 B.n505 B.n36 585
R327 B.n504 B.n503 585
R328 B.n502 B.n37 585
R329 B.n501 B.n500 585
R330 B.n499 B.n41 585
R331 B.n498 B.n497 585
R332 B.n496 B.n42 585
R333 B.n495 B.n494 585
R334 B.n493 B.n43 585
R335 B.n492 B.n491 585
R336 B.n490 B.n44 585
R337 B.n488 B.n487 585
R338 B.n486 B.n47 585
R339 B.n485 B.n484 585
R340 B.n483 B.n48 585
R341 B.n482 B.n481 585
R342 B.n480 B.n49 585
R343 B.n479 B.n478 585
R344 B.n477 B.n50 585
R345 B.n476 B.n475 585
R346 B.n474 B.n51 585
R347 B.n473 B.n472 585
R348 B.n471 B.n52 585
R349 B.n470 B.n469 585
R350 B.n468 B.n53 585
R351 B.n467 B.n466 585
R352 B.n465 B.n54 585
R353 B.n464 B.n463 585
R354 B.n462 B.n55 585
R355 B.n461 B.n460 585
R356 B.n459 B.n56 585
R357 B.n458 B.n457 585
R358 B.n456 B.n57 585
R359 B.n455 B.n454 585
R360 B.n453 B.n58 585
R361 B.n452 B.n451 585
R362 B.n450 B.n59 585
R363 B.n449 B.n448 585
R364 B.n447 B.n60 585
R365 B.n446 B.n445 585
R366 B.n444 B.n61 585
R367 B.n443 B.n442 585
R368 B.n441 B.n62 585
R369 B.n440 B.n439 585
R370 B.n438 B.n63 585
R371 B.n437 B.n436 585
R372 B.n435 B.n64 585
R373 B.n434 B.n433 585
R374 B.n432 B.n65 585
R375 B.n431 B.n430 585
R376 B.n429 B.n66 585
R377 B.n428 B.n427 585
R378 B.n426 B.n67 585
R379 B.n425 B.n424 585
R380 B.n423 B.n68 585
R381 B.n422 B.n421 585
R382 B.n420 B.n69 585
R383 B.n419 B.n418 585
R384 B.n417 B.n70 585
R385 B.n416 B.n415 585
R386 B.n579 B.n578 585
R387 B.n580 B.n11 585
R388 B.n582 B.n581 585
R389 B.n583 B.n10 585
R390 B.n585 B.n584 585
R391 B.n586 B.n9 585
R392 B.n588 B.n587 585
R393 B.n589 B.n8 585
R394 B.n591 B.n590 585
R395 B.n592 B.n7 585
R396 B.n594 B.n593 585
R397 B.n595 B.n6 585
R398 B.n597 B.n596 585
R399 B.n598 B.n5 585
R400 B.n600 B.n599 585
R401 B.n601 B.n4 585
R402 B.n603 B.n602 585
R403 B.n604 B.n3 585
R404 B.n606 B.n605 585
R405 B.n607 B.n0 585
R406 B.n2 B.n1 585
R407 B.n158 B.n157 585
R408 B.n160 B.n159 585
R409 B.n161 B.n156 585
R410 B.n163 B.n162 585
R411 B.n164 B.n155 585
R412 B.n166 B.n165 585
R413 B.n167 B.n154 585
R414 B.n169 B.n168 585
R415 B.n170 B.n153 585
R416 B.n172 B.n171 585
R417 B.n173 B.n152 585
R418 B.n175 B.n174 585
R419 B.n176 B.n151 585
R420 B.n178 B.n177 585
R421 B.n179 B.n150 585
R422 B.n181 B.n180 585
R423 B.n182 B.n149 585
R424 B.n184 B.n183 585
R425 B.n185 B.n148 585
R426 B.n187 B.n148 482.89
R427 B.n353 B.n92 482.89
R428 B.n415 B.n414 482.89
R429 B.n578 B.n577 482.89
R430 B.n609 B.n608 256.663
R431 B.n608 B.n607 235.042
R432 B.n608 B.n2 235.042
R433 B.n188 B.n187 163.367
R434 B.n189 B.n188 163.367
R435 B.n189 B.n146 163.367
R436 B.n193 B.n146 163.367
R437 B.n194 B.n193 163.367
R438 B.n195 B.n194 163.367
R439 B.n195 B.n144 163.367
R440 B.n199 B.n144 163.367
R441 B.n200 B.n199 163.367
R442 B.n201 B.n200 163.367
R443 B.n201 B.n142 163.367
R444 B.n205 B.n142 163.367
R445 B.n206 B.n205 163.367
R446 B.n207 B.n206 163.367
R447 B.n207 B.n140 163.367
R448 B.n211 B.n140 163.367
R449 B.n212 B.n211 163.367
R450 B.n213 B.n212 163.367
R451 B.n213 B.n138 163.367
R452 B.n217 B.n138 163.367
R453 B.n218 B.n217 163.367
R454 B.n219 B.n218 163.367
R455 B.n219 B.n136 163.367
R456 B.n223 B.n136 163.367
R457 B.n224 B.n223 163.367
R458 B.n225 B.n224 163.367
R459 B.n225 B.n134 163.367
R460 B.n229 B.n134 163.367
R461 B.n230 B.n229 163.367
R462 B.n231 B.n230 163.367
R463 B.n231 B.n132 163.367
R464 B.n235 B.n132 163.367
R465 B.n236 B.n235 163.367
R466 B.n237 B.n236 163.367
R467 B.n237 B.n130 163.367
R468 B.n241 B.n130 163.367
R469 B.n242 B.n241 163.367
R470 B.n243 B.n242 163.367
R471 B.n243 B.n128 163.367
R472 B.n247 B.n128 163.367
R473 B.n248 B.n247 163.367
R474 B.n249 B.n248 163.367
R475 B.n249 B.n126 163.367
R476 B.n253 B.n126 163.367
R477 B.n254 B.n253 163.367
R478 B.n255 B.n254 163.367
R479 B.n255 B.n124 163.367
R480 B.n262 B.n124 163.367
R481 B.n263 B.n262 163.367
R482 B.n264 B.n263 163.367
R483 B.n264 B.n122 163.367
R484 B.n268 B.n122 163.367
R485 B.n269 B.n268 163.367
R486 B.n270 B.n269 163.367
R487 B.n270 B.n120 163.367
R488 B.n274 B.n120 163.367
R489 B.n275 B.n274 163.367
R490 B.n276 B.n275 163.367
R491 B.n276 B.n116 163.367
R492 B.n281 B.n116 163.367
R493 B.n282 B.n281 163.367
R494 B.n283 B.n282 163.367
R495 B.n283 B.n114 163.367
R496 B.n287 B.n114 163.367
R497 B.n288 B.n287 163.367
R498 B.n289 B.n288 163.367
R499 B.n289 B.n112 163.367
R500 B.n293 B.n112 163.367
R501 B.n294 B.n293 163.367
R502 B.n295 B.n294 163.367
R503 B.n295 B.n110 163.367
R504 B.n299 B.n110 163.367
R505 B.n300 B.n299 163.367
R506 B.n301 B.n300 163.367
R507 B.n301 B.n108 163.367
R508 B.n305 B.n108 163.367
R509 B.n306 B.n305 163.367
R510 B.n307 B.n306 163.367
R511 B.n307 B.n106 163.367
R512 B.n311 B.n106 163.367
R513 B.n312 B.n311 163.367
R514 B.n313 B.n312 163.367
R515 B.n313 B.n104 163.367
R516 B.n317 B.n104 163.367
R517 B.n318 B.n317 163.367
R518 B.n319 B.n318 163.367
R519 B.n319 B.n102 163.367
R520 B.n323 B.n102 163.367
R521 B.n324 B.n323 163.367
R522 B.n325 B.n324 163.367
R523 B.n325 B.n100 163.367
R524 B.n329 B.n100 163.367
R525 B.n330 B.n329 163.367
R526 B.n331 B.n330 163.367
R527 B.n331 B.n98 163.367
R528 B.n335 B.n98 163.367
R529 B.n336 B.n335 163.367
R530 B.n337 B.n336 163.367
R531 B.n337 B.n96 163.367
R532 B.n341 B.n96 163.367
R533 B.n342 B.n341 163.367
R534 B.n343 B.n342 163.367
R535 B.n343 B.n94 163.367
R536 B.n347 B.n94 163.367
R537 B.n348 B.n347 163.367
R538 B.n349 B.n348 163.367
R539 B.n349 B.n92 163.367
R540 B.n414 B.n413 163.367
R541 B.n413 B.n72 163.367
R542 B.n409 B.n72 163.367
R543 B.n409 B.n408 163.367
R544 B.n408 B.n407 163.367
R545 B.n407 B.n74 163.367
R546 B.n403 B.n74 163.367
R547 B.n403 B.n402 163.367
R548 B.n402 B.n401 163.367
R549 B.n401 B.n76 163.367
R550 B.n397 B.n76 163.367
R551 B.n397 B.n396 163.367
R552 B.n396 B.n395 163.367
R553 B.n395 B.n78 163.367
R554 B.n391 B.n78 163.367
R555 B.n391 B.n390 163.367
R556 B.n390 B.n389 163.367
R557 B.n389 B.n80 163.367
R558 B.n385 B.n80 163.367
R559 B.n385 B.n384 163.367
R560 B.n384 B.n383 163.367
R561 B.n383 B.n82 163.367
R562 B.n379 B.n82 163.367
R563 B.n379 B.n378 163.367
R564 B.n378 B.n377 163.367
R565 B.n377 B.n84 163.367
R566 B.n373 B.n84 163.367
R567 B.n373 B.n372 163.367
R568 B.n372 B.n371 163.367
R569 B.n371 B.n86 163.367
R570 B.n367 B.n86 163.367
R571 B.n367 B.n366 163.367
R572 B.n366 B.n365 163.367
R573 B.n365 B.n88 163.367
R574 B.n361 B.n88 163.367
R575 B.n361 B.n360 163.367
R576 B.n360 B.n359 163.367
R577 B.n359 B.n90 163.367
R578 B.n355 B.n90 163.367
R579 B.n355 B.n354 163.367
R580 B.n354 B.n353 163.367
R581 B.n577 B.n576 163.367
R582 B.n576 B.n13 163.367
R583 B.n572 B.n13 163.367
R584 B.n572 B.n571 163.367
R585 B.n571 B.n570 163.367
R586 B.n570 B.n15 163.367
R587 B.n566 B.n15 163.367
R588 B.n566 B.n565 163.367
R589 B.n565 B.n564 163.367
R590 B.n564 B.n17 163.367
R591 B.n560 B.n17 163.367
R592 B.n560 B.n559 163.367
R593 B.n559 B.n558 163.367
R594 B.n558 B.n19 163.367
R595 B.n554 B.n19 163.367
R596 B.n554 B.n553 163.367
R597 B.n553 B.n552 163.367
R598 B.n552 B.n21 163.367
R599 B.n548 B.n21 163.367
R600 B.n548 B.n547 163.367
R601 B.n547 B.n546 163.367
R602 B.n546 B.n23 163.367
R603 B.n542 B.n23 163.367
R604 B.n542 B.n541 163.367
R605 B.n541 B.n540 163.367
R606 B.n540 B.n25 163.367
R607 B.n536 B.n25 163.367
R608 B.n536 B.n535 163.367
R609 B.n535 B.n534 163.367
R610 B.n534 B.n27 163.367
R611 B.n530 B.n27 163.367
R612 B.n530 B.n529 163.367
R613 B.n529 B.n528 163.367
R614 B.n528 B.n29 163.367
R615 B.n524 B.n29 163.367
R616 B.n524 B.n523 163.367
R617 B.n523 B.n522 163.367
R618 B.n522 B.n31 163.367
R619 B.n518 B.n31 163.367
R620 B.n518 B.n517 163.367
R621 B.n517 B.n516 163.367
R622 B.n516 B.n33 163.367
R623 B.n512 B.n33 163.367
R624 B.n512 B.n511 163.367
R625 B.n511 B.n510 163.367
R626 B.n510 B.n35 163.367
R627 B.n506 B.n35 163.367
R628 B.n506 B.n505 163.367
R629 B.n505 B.n504 163.367
R630 B.n504 B.n37 163.367
R631 B.n500 B.n37 163.367
R632 B.n500 B.n499 163.367
R633 B.n499 B.n498 163.367
R634 B.n498 B.n42 163.367
R635 B.n494 B.n42 163.367
R636 B.n494 B.n493 163.367
R637 B.n493 B.n492 163.367
R638 B.n492 B.n44 163.367
R639 B.n487 B.n44 163.367
R640 B.n487 B.n486 163.367
R641 B.n486 B.n485 163.367
R642 B.n485 B.n48 163.367
R643 B.n481 B.n48 163.367
R644 B.n481 B.n480 163.367
R645 B.n480 B.n479 163.367
R646 B.n479 B.n50 163.367
R647 B.n475 B.n50 163.367
R648 B.n475 B.n474 163.367
R649 B.n474 B.n473 163.367
R650 B.n473 B.n52 163.367
R651 B.n469 B.n52 163.367
R652 B.n469 B.n468 163.367
R653 B.n468 B.n467 163.367
R654 B.n467 B.n54 163.367
R655 B.n463 B.n54 163.367
R656 B.n463 B.n462 163.367
R657 B.n462 B.n461 163.367
R658 B.n461 B.n56 163.367
R659 B.n457 B.n56 163.367
R660 B.n457 B.n456 163.367
R661 B.n456 B.n455 163.367
R662 B.n455 B.n58 163.367
R663 B.n451 B.n58 163.367
R664 B.n451 B.n450 163.367
R665 B.n450 B.n449 163.367
R666 B.n449 B.n60 163.367
R667 B.n445 B.n60 163.367
R668 B.n445 B.n444 163.367
R669 B.n444 B.n443 163.367
R670 B.n443 B.n62 163.367
R671 B.n439 B.n62 163.367
R672 B.n439 B.n438 163.367
R673 B.n438 B.n437 163.367
R674 B.n437 B.n64 163.367
R675 B.n433 B.n64 163.367
R676 B.n433 B.n432 163.367
R677 B.n432 B.n431 163.367
R678 B.n431 B.n66 163.367
R679 B.n427 B.n66 163.367
R680 B.n427 B.n426 163.367
R681 B.n426 B.n425 163.367
R682 B.n425 B.n68 163.367
R683 B.n421 B.n68 163.367
R684 B.n421 B.n420 163.367
R685 B.n420 B.n419 163.367
R686 B.n419 B.n70 163.367
R687 B.n415 B.n70 163.367
R688 B.n578 B.n11 163.367
R689 B.n582 B.n11 163.367
R690 B.n583 B.n582 163.367
R691 B.n584 B.n583 163.367
R692 B.n584 B.n9 163.367
R693 B.n588 B.n9 163.367
R694 B.n589 B.n588 163.367
R695 B.n590 B.n589 163.367
R696 B.n590 B.n7 163.367
R697 B.n594 B.n7 163.367
R698 B.n595 B.n594 163.367
R699 B.n596 B.n595 163.367
R700 B.n596 B.n5 163.367
R701 B.n600 B.n5 163.367
R702 B.n601 B.n600 163.367
R703 B.n602 B.n601 163.367
R704 B.n602 B.n3 163.367
R705 B.n606 B.n3 163.367
R706 B.n607 B.n606 163.367
R707 B.n158 B.n2 163.367
R708 B.n159 B.n158 163.367
R709 B.n159 B.n156 163.367
R710 B.n163 B.n156 163.367
R711 B.n164 B.n163 163.367
R712 B.n165 B.n164 163.367
R713 B.n165 B.n154 163.367
R714 B.n169 B.n154 163.367
R715 B.n170 B.n169 163.367
R716 B.n171 B.n170 163.367
R717 B.n171 B.n152 163.367
R718 B.n175 B.n152 163.367
R719 B.n176 B.n175 163.367
R720 B.n177 B.n176 163.367
R721 B.n177 B.n150 163.367
R722 B.n181 B.n150 163.367
R723 B.n182 B.n181 163.367
R724 B.n183 B.n182 163.367
R725 B.n183 B.n148 163.367
R726 B.n117 B.t1 127.579
R727 B.n45 B.t11 127.579
R728 B.n258 B.t4 127.561
R729 B.n38 B.t8 127.561
R730 B.n118 B.t2 111.094
R731 B.n46 B.t10 111.094
R732 B.n259 B.t5 111.076
R733 B.n39 B.t7 111.076
R734 B.n260 B.n259 59.5399
R735 B.n278 B.n118 59.5399
R736 B.n489 B.n46 59.5399
R737 B.n40 B.n39 59.5399
R738 B.n579 B.n12 31.3761
R739 B.n416 B.n71 31.3761
R740 B.n352 B.n351 31.3761
R741 B.n186 B.n185 31.3761
R742 B B.n609 18.0485
R743 B.n259 B.n258 16.4853
R744 B.n118 B.n117 16.4853
R745 B.n46 B.n45 16.4853
R746 B.n39 B.n38 16.4853
R747 B.n580 B.n579 10.6151
R748 B.n581 B.n580 10.6151
R749 B.n581 B.n10 10.6151
R750 B.n585 B.n10 10.6151
R751 B.n586 B.n585 10.6151
R752 B.n587 B.n586 10.6151
R753 B.n587 B.n8 10.6151
R754 B.n591 B.n8 10.6151
R755 B.n592 B.n591 10.6151
R756 B.n593 B.n592 10.6151
R757 B.n593 B.n6 10.6151
R758 B.n597 B.n6 10.6151
R759 B.n598 B.n597 10.6151
R760 B.n599 B.n598 10.6151
R761 B.n599 B.n4 10.6151
R762 B.n603 B.n4 10.6151
R763 B.n604 B.n603 10.6151
R764 B.n605 B.n604 10.6151
R765 B.n605 B.n0 10.6151
R766 B.n575 B.n12 10.6151
R767 B.n575 B.n574 10.6151
R768 B.n574 B.n573 10.6151
R769 B.n573 B.n14 10.6151
R770 B.n569 B.n14 10.6151
R771 B.n569 B.n568 10.6151
R772 B.n568 B.n567 10.6151
R773 B.n567 B.n16 10.6151
R774 B.n563 B.n16 10.6151
R775 B.n563 B.n562 10.6151
R776 B.n562 B.n561 10.6151
R777 B.n561 B.n18 10.6151
R778 B.n557 B.n18 10.6151
R779 B.n557 B.n556 10.6151
R780 B.n556 B.n555 10.6151
R781 B.n555 B.n20 10.6151
R782 B.n551 B.n20 10.6151
R783 B.n551 B.n550 10.6151
R784 B.n550 B.n549 10.6151
R785 B.n549 B.n22 10.6151
R786 B.n545 B.n22 10.6151
R787 B.n545 B.n544 10.6151
R788 B.n544 B.n543 10.6151
R789 B.n543 B.n24 10.6151
R790 B.n539 B.n24 10.6151
R791 B.n539 B.n538 10.6151
R792 B.n538 B.n537 10.6151
R793 B.n537 B.n26 10.6151
R794 B.n533 B.n26 10.6151
R795 B.n533 B.n532 10.6151
R796 B.n532 B.n531 10.6151
R797 B.n531 B.n28 10.6151
R798 B.n527 B.n28 10.6151
R799 B.n527 B.n526 10.6151
R800 B.n526 B.n525 10.6151
R801 B.n525 B.n30 10.6151
R802 B.n521 B.n30 10.6151
R803 B.n521 B.n520 10.6151
R804 B.n520 B.n519 10.6151
R805 B.n519 B.n32 10.6151
R806 B.n515 B.n32 10.6151
R807 B.n515 B.n514 10.6151
R808 B.n514 B.n513 10.6151
R809 B.n513 B.n34 10.6151
R810 B.n509 B.n34 10.6151
R811 B.n509 B.n508 10.6151
R812 B.n508 B.n507 10.6151
R813 B.n507 B.n36 10.6151
R814 B.n503 B.n502 10.6151
R815 B.n502 B.n501 10.6151
R816 B.n501 B.n41 10.6151
R817 B.n497 B.n41 10.6151
R818 B.n497 B.n496 10.6151
R819 B.n496 B.n495 10.6151
R820 B.n495 B.n43 10.6151
R821 B.n491 B.n43 10.6151
R822 B.n491 B.n490 10.6151
R823 B.n488 B.n47 10.6151
R824 B.n484 B.n47 10.6151
R825 B.n484 B.n483 10.6151
R826 B.n483 B.n482 10.6151
R827 B.n482 B.n49 10.6151
R828 B.n478 B.n49 10.6151
R829 B.n478 B.n477 10.6151
R830 B.n477 B.n476 10.6151
R831 B.n476 B.n51 10.6151
R832 B.n472 B.n51 10.6151
R833 B.n472 B.n471 10.6151
R834 B.n471 B.n470 10.6151
R835 B.n470 B.n53 10.6151
R836 B.n466 B.n53 10.6151
R837 B.n466 B.n465 10.6151
R838 B.n465 B.n464 10.6151
R839 B.n464 B.n55 10.6151
R840 B.n460 B.n55 10.6151
R841 B.n460 B.n459 10.6151
R842 B.n459 B.n458 10.6151
R843 B.n458 B.n57 10.6151
R844 B.n454 B.n57 10.6151
R845 B.n454 B.n453 10.6151
R846 B.n453 B.n452 10.6151
R847 B.n452 B.n59 10.6151
R848 B.n448 B.n59 10.6151
R849 B.n448 B.n447 10.6151
R850 B.n447 B.n446 10.6151
R851 B.n446 B.n61 10.6151
R852 B.n442 B.n61 10.6151
R853 B.n442 B.n441 10.6151
R854 B.n441 B.n440 10.6151
R855 B.n440 B.n63 10.6151
R856 B.n436 B.n63 10.6151
R857 B.n436 B.n435 10.6151
R858 B.n435 B.n434 10.6151
R859 B.n434 B.n65 10.6151
R860 B.n430 B.n65 10.6151
R861 B.n430 B.n429 10.6151
R862 B.n429 B.n428 10.6151
R863 B.n428 B.n67 10.6151
R864 B.n424 B.n67 10.6151
R865 B.n424 B.n423 10.6151
R866 B.n423 B.n422 10.6151
R867 B.n422 B.n69 10.6151
R868 B.n418 B.n69 10.6151
R869 B.n418 B.n417 10.6151
R870 B.n417 B.n416 10.6151
R871 B.n412 B.n71 10.6151
R872 B.n412 B.n411 10.6151
R873 B.n411 B.n410 10.6151
R874 B.n410 B.n73 10.6151
R875 B.n406 B.n73 10.6151
R876 B.n406 B.n405 10.6151
R877 B.n405 B.n404 10.6151
R878 B.n404 B.n75 10.6151
R879 B.n400 B.n75 10.6151
R880 B.n400 B.n399 10.6151
R881 B.n399 B.n398 10.6151
R882 B.n398 B.n77 10.6151
R883 B.n394 B.n77 10.6151
R884 B.n394 B.n393 10.6151
R885 B.n393 B.n392 10.6151
R886 B.n392 B.n79 10.6151
R887 B.n388 B.n79 10.6151
R888 B.n388 B.n387 10.6151
R889 B.n387 B.n386 10.6151
R890 B.n386 B.n81 10.6151
R891 B.n382 B.n81 10.6151
R892 B.n382 B.n381 10.6151
R893 B.n381 B.n380 10.6151
R894 B.n380 B.n83 10.6151
R895 B.n376 B.n83 10.6151
R896 B.n376 B.n375 10.6151
R897 B.n375 B.n374 10.6151
R898 B.n374 B.n85 10.6151
R899 B.n370 B.n85 10.6151
R900 B.n370 B.n369 10.6151
R901 B.n369 B.n368 10.6151
R902 B.n368 B.n87 10.6151
R903 B.n364 B.n87 10.6151
R904 B.n364 B.n363 10.6151
R905 B.n363 B.n362 10.6151
R906 B.n362 B.n89 10.6151
R907 B.n358 B.n89 10.6151
R908 B.n358 B.n357 10.6151
R909 B.n357 B.n356 10.6151
R910 B.n356 B.n91 10.6151
R911 B.n352 B.n91 10.6151
R912 B.n157 B.n1 10.6151
R913 B.n160 B.n157 10.6151
R914 B.n161 B.n160 10.6151
R915 B.n162 B.n161 10.6151
R916 B.n162 B.n155 10.6151
R917 B.n166 B.n155 10.6151
R918 B.n167 B.n166 10.6151
R919 B.n168 B.n167 10.6151
R920 B.n168 B.n153 10.6151
R921 B.n172 B.n153 10.6151
R922 B.n173 B.n172 10.6151
R923 B.n174 B.n173 10.6151
R924 B.n174 B.n151 10.6151
R925 B.n178 B.n151 10.6151
R926 B.n179 B.n178 10.6151
R927 B.n180 B.n179 10.6151
R928 B.n180 B.n149 10.6151
R929 B.n184 B.n149 10.6151
R930 B.n185 B.n184 10.6151
R931 B.n186 B.n147 10.6151
R932 B.n190 B.n147 10.6151
R933 B.n191 B.n190 10.6151
R934 B.n192 B.n191 10.6151
R935 B.n192 B.n145 10.6151
R936 B.n196 B.n145 10.6151
R937 B.n197 B.n196 10.6151
R938 B.n198 B.n197 10.6151
R939 B.n198 B.n143 10.6151
R940 B.n202 B.n143 10.6151
R941 B.n203 B.n202 10.6151
R942 B.n204 B.n203 10.6151
R943 B.n204 B.n141 10.6151
R944 B.n208 B.n141 10.6151
R945 B.n209 B.n208 10.6151
R946 B.n210 B.n209 10.6151
R947 B.n210 B.n139 10.6151
R948 B.n214 B.n139 10.6151
R949 B.n215 B.n214 10.6151
R950 B.n216 B.n215 10.6151
R951 B.n216 B.n137 10.6151
R952 B.n220 B.n137 10.6151
R953 B.n221 B.n220 10.6151
R954 B.n222 B.n221 10.6151
R955 B.n222 B.n135 10.6151
R956 B.n226 B.n135 10.6151
R957 B.n227 B.n226 10.6151
R958 B.n228 B.n227 10.6151
R959 B.n228 B.n133 10.6151
R960 B.n232 B.n133 10.6151
R961 B.n233 B.n232 10.6151
R962 B.n234 B.n233 10.6151
R963 B.n234 B.n131 10.6151
R964 B.n238 B.n131 10.6151
R965 B.n239 B.n238 10.6151
R966 B.n240 B.n239 10.6151
R967 B.n240 B.n129 10.6151
R968 B.n244 B.n129 10.6151
R969 B.n245 B.n244 10.6151
R970 B.n246 B.n245 10.6151
R971 B.n246 B.n127 10.6151
R972 B.n250 B.n127 10.6151
R973 B.n251 B.n250 10.6151
R974 B.n252 B.n251 10.6151
R975 B.n252 B.n125 10.6151
R976 B.n256 B.n125 10.6151
R977 B.n257 B.n256 10.6151
R978 B.n261 B.n257 10.6151
R979 B.n265 B.n123 10.6151
R980 B.n266 B.n265 10.6151
R981 B.n267 B.n266 10.6151
R982 B.n267 B.n121 10.6151
R983 B.n271 B.n121 10.6151
R984 B.n272 B.n271 10.6151
R985 B.n273 B.n272 10.6151
R986 B.n273 B.n119 10.6151
R987 B.n277 B.n119 10.6151
R988 B.n280 B.n279 10.6151
R989 B.n280 B.n115 10.6151
R990 B.n284 B.n115 10.6151
R991 B.n285 B.n284 10.6151
R992 B.n286 B.n285 10.6151
R993 B.n286 B.n113 10.6151
R994 B.n290 B.n113 10.6151
R995 B.n291 B.n290 10.6151
R996 B.n292 B.n291 10.6151
R997 B.n292 B.n111 10.6151
R998 B.n296 B.n111 10.6151
R999 B.n297 B.n296 10.6151
R1000 B.n298 B.n297 10.6151
R1001 B.n298 B.n109 10.6151
R1002 B.n302 B.n109 10.6151
R1003 B.n303 B.n302 10.6151
R1004 B.n304 B.n303 10.6151
R1005 B.n304 B.n107 10.6151
R1006 B.n308 B.n107 10.6151
R1007 B.n309 B.n308 10.6151
R1008 B.n310 B.n309 10.6151
R1009 B.n310 B.n105 10.6151
R1010 B.n314 B.n105 10.6151
R1011 B.n315 B.n314 10.6151
R1012 B.n316 B.n315 10.6151
R1013 B.n316 B.n103 10.6151
R1014 B.n320 B.n103 10.6151
R1015 B.n321 B.n320 10.6151
R1016 B.n322 B.n321 10.6151
R1017 B.n322 B.n101 10.6151
R1018 B.n326 B.n101 10.6151
R1019 B.n327 B.n326 10.6151
R1020 B.n328 B.n327 10.6151
R1021 B.n328 B.n99 10.6151
R1022 B.n332 B.n99 10.6151
R1023 B.n333 B.n332 10.6151
R1024 B.n334 B.n333 10.6151
R1025 B.n334 B.n97 10.6151
R1026 B.n338 B.n97 10.6151
R1027 B.n339 B.n338 10.6151
R1028 B.n340 B.n339 10.6151
R1029 B.n340 B.n95 10.6151
R1030 B.n344 B.n95 10.6151
R1031 B.n345 B.n344 10.6151
R1032 B.n346 B.n345 10.6151
R1033 B.n346 B.n93 10.6151
R1034 B.n350 B.n93 10.6151
R1035 B.n351 B.n350 10.6151
R1036 B.n40 B.n36 9.36635
R1037 B.n489 B.n488 9.36635
R1038 B.n261 B.n260 9.36635
R1039 B.n279 B.n278 9.36635
R1040 B.n609 B.n0 8.11757
R1041 B.n609 B.n1 8.11757
R1042 B.n503 B.n40 1.24928
R1043 B.n490 B.n489 1.24928
R1044 B.n260 B.n123 1.24928
R1045 B.n278 B.n277 1.24928
C0 VDD2 B 1.11377f
C1 w_n1820_n3870# VTAIL 4.86945f
C2 VDD1 VTAIL 14.9494f
C3 VN VTAIL 5.16843f
C4 w_n1820_n3870# VDD1 1.29618f
C5 VDD2 VTAIL 14.989799f
C6 w_n1820_n3870# VN 3.16132f
C7 VDD1 VN 0.147934f
C8 VP B 1.14276f
C9 VDD2 w_n1820_n3870# 1.32356f
C10 VDD2 VDD1 0.737654f
C11 VDD2 VN 5.58047f
C12 VP VTAIL 5.18254f
C13 w_n1820_n3870# VP 3.39146f
C14 VTAIL B 4.34492f
C15 VDD1 VP 5.7305f
C16 VP VN 5.57994f
C17 w_n1820_n3870# B 7.63741f
C18 VDD1 B 1.08266f
C19 VDD2 VP 0.298303f
C20 VN B 0.768051f
C21 VDD2 VSUBS 1.383375f
C22 VDD1 VSUBS 1.653954f
C23 VTAIL VSUBS 0.927693f
C24 VN VSUBS 4.8066f
C25 VP VSUBS 1.564842f
C26 B VSUBS 2.890743f
C27 w_n1820_n3870# VSUBS 86.4209f
C28 B.n0 VSUBS 0.007141f
C29 B.n1 VSUBS 0.007141f
C30 B.n2 VSUBS 0.010561f
C31 B.n3 VSUBS 0.008093f
C32 B.n4 VSUBS 0.008093f
C33 B.n5 VSUBS 0.008093f
C34 B.n6 VSUBS 0.008093f
C35 B.n7 VSUBS 0.008093f
C36 B.n8 VSUBS 0.008093f
C37 B.n9 VSUBS 0.008093f
C38 B.n10 VSUBS 0.008093f
C39 B.n11 VSUBS 0.008093f
C40 B.n12 VSUBS 0.019189f
C41 B.n13 VSUBS 0.008093f
C42 B.n14 VSUBS 0.008093f
C43 B.n15 VSUBS 0.008093f
C44 B.n16 VSUBS 0.008093f
C45 B.n17 VSUBS 0.008093f
C46 B.n18 VSUBS 0.008093f
C47 B.n19 VSUBS 0.008093f
C48 B.n20 VSUBS 0.008093f
C49 B.n21 VSUBS 0.008093f
C50 B.n22 VSUBS 0.008093f
C51 B.n23 VSUBS 0.008093f
C52 B.n24 VSUBS 0.008093f
C53 B.n25 VSUBS 0.008093f
C54 B.n26 VSUBS 0.008093f
C55 B.n27 VSUBS 0.008093f
C56 B.n28 VSUBS 0.008093f
C57 B.n29 VSUBS 0.008093f
C58 B.n30 VSUBS 0.008093f
C59 B.n31 VSUBS 0.008093f
C60 B.n32 VSUBS 0.008093f
C61 B.n33 VSUBS 0.008093f
C62 B.n34 VSUBS 0.008093f
C63 B.n35 VSUBS 0.008093f
C64 B.n36 VSUBS 0.007617f
C65 B.n37 VSUBS 0.008093f
C66 B.t7 VSUBS 0.556908f
C67 B.t8 VSUBS 0.564878f
C68 B.t6 VSUBS 0.349486f
C69 B.n38 VSUBS 0.156745f
C70 B.n39 VSUBS 0.073214f
C71 B.n40 VSUBS 0.018752f
C72 B.n41 VSUBS 0.008093f
C73 B.n42 VSUBS 0.008093f
C74 B.n43 VSUBS 0.008093f
C75 B.n44 VSUBS 0.008093f
C76 B.t10 VSUBS 0.556893f
C77 B.t11 VSUBS 0.564864f
C78 B.t9 VSUBS 0.349486f
C79 B.n45 VSUBS 0.156759f
C80 B.n46 VSUBS 0.073228f
C81 B.n47 VSUBS 0.008093f
C82 B.n48 VSUBS 0.008093f
C83 B.n49 VSUBS 0.008093f
C84 B.n50 VSUBS 0.008093f
C85 B.n51 VSUBS 0.008093f
C86 B.n52 VSUBS 0.008093f
C87 B.n53 VSUBS 0.008093f
C88 B.n54 VSUBS 0.008093f
C89 B.n55 VSUBS 0.008093f
C90 B.n56 VSUBS 0.008093f
C91 B.n57 VSUBS 0.008093f
C92 B.n58 VSUBS 0.008093f
C93 B.n59 VSUBS 0.008093f
C94 B.n60 VSUBS 0.008093f
C95 B.n61 VSUBS 0.008093f
C96 B.n62 VSUBS 0.008093f
C97 B.n63 VSUBS 0.008093f
C98 B.n64 VSUBS 0.008093f
C99 B.n65 VSUBS 0.008093f
C100 B.n66 VSUBS 0.008093f
C101 B.n67 VSUBS 0.008093f
C102 B.n68 VSUBS 0.008093f
C103 B.n69 VSUBS 0.008093f
C104 B.n70 VSUBS 0.008093f
C105 B.n71 VSUBS 0.017708f
C106 B.n72 VSUBS 0.008093f
C107 B.n73 VSUBS 0.008093f
C108 B.n74 VSUBS 0.008093f
C109 B.n75 VSUBS 0.008093f
C110 B.n76 VSUBS 0.008093f
C111 B.n77 VSUBS 0.008093f
C112 B.n78 VSUBS 0.008093f
C113 B.n79 VSUBS 0.008093f
C114 B.n80 VSUBS 0.008093f
C115 B.n81 VSUBS 0.008093f
C116 B.n82 VSUBS 0.008093f
C117 B.n83 VSUBS 0.008093f
C118 B.n84 VSUBS 0.008093f
C119 B.n85 VSUBS 0.008093f
C120 B.n86 VSUBS 0.008093f
C121 B.n87 VSUBS 0.008093f
C122 B.n88 VSUBS 0.008093f
C123 B.n89 VSUBS 0.008093f
C124 B.n90 VSUBS 0.008093f
C125 B.n91 VSUBS 0.008093f
C126 B.n92 VSUBS 0.019189f
C127 B.n93 VSUBS 0.008093f
C128 B.n94 VSUBS 0.008093f
C129 B.n95 VSUBS 0.008093f
C130 B.n96 VSUBS 0.008093f
C131 B.n97 VSUBS 0.008093f
C132 B.n98 VSUBS 0.008093f
C133 B.n99 VSUBS 0.008093f
C134 B.n100 VSUBS 0.008093f
C135 B.n101 VSUBS 0.008093f
C136 B.n102 VSUBS 0.008093f
C137 B.n103 VSUBS 0.008093f
C138 B.n104 VSUBS 0.008093f
C139 B.n105 VSUBS 0.008093f
C140 B.n106 VSUBS 0.008093f
C141 B.n107 VSUBS 0.008093f
C142 B.n108 VSUBS 0.008093f
C143 B.n109 VSUBS 0.008093f
C144 B.n110 VSUBS 0.008093f
C145 B.n111 VSUBS 0.008093f
C146 B.n112 VSUBS 0.008093f
C147 B.n113 VSUBS 0.008093f
C148 B.n114 VSUBS 0.008093f
C149 B.n115 VSUBS 0.008093f
C150 B.n116 VSUBS 0.008093f
C151 B.t2 VSUBS 0.556893f
C152 B.t1 VSUBS 0.564864f
C153 B.t0 VSUBS 0.349486f
C154 B.n117 VSUBS 0.156759f
C155 B.n118 VSUBS 0.073228f
C156 B.n119 VSUBS 0.008093f
C157 B.n120 VSUBS 0.008093f
C158 B.n121 VSUBS 0.008093f
C159 B.n122 VSUBS 0.008093f
C160 B.n123 VSUBS 0.004523f
C161 B.n124 VSUBS 0.008093f
C162 B.n125 VSUBS 0.008093f
C163 B.n126 VSUBS 0.008093f
C164 B.n127 VSUBS 0.008093f
C165 B.n128 VSUBS 0.008093f
C166 B.n129 VSUBS 0.008093f
C167 B.n130 VSUBS 0.008093f
C168 B.n131 VSUBS 0.008093f
C169 B.n132 VSUBS 0.008093f
C170 B.n133 VSUBS 0.008093f
C171 B.n134 VSUBS 0.008093f
C172 B.n135 VSUBS 0.008093f
C173 B.n136 VSUBS 0.008093f
C174 B.n137 VSUBS 0.008093f
C175 B.n138 VSUBS 0.008093f
C176 B.n139 VSUBS 0.008093f
C177 B.n140 VSUBS 0.008093f
C178 B.n141 VSUBS 0.008093f
C179 B.n142 VSUBS 0.008093f
C180 B.n143 VSUBS 0.008093f
C181 B.n144 VSUBS 0.008093f
C182 B.n145 VSUBS 0.008093f
C183 B.n146 VSUBS 0.008093f
C184 B.n147 VSUBS 0.008093f
C185 B.n148 VSUBS 0.017708f
C186 B.n149 VSUBS 0.008093f
C187 B.n150 VSUBS 0.008093f
C188 B.n151 VSUBS 0.008093f
C189 B.n152 VSUBS 0.008093f
C190 B.n153 VSUBS 0.008093f
C191 B.n154 VSUBS 0.008093f
C192 B.n155 VSUBS 0.008093f
C193 B.n156 VSUBS 0.008093f
C194 B.n157 VSUBS 0.008093f
C195 B.n158 VSUBS 0.008093f
C196 B.n159 VSUBS 0.008093f
C197 B.n160 VSUBS 0.008093f
C198 B.n161 VSUBS 0.008093f
C199 B.n162 VSUBS 0.008093f
C200 B.n163 VSUBS 0.008093f
C201 B.n164 VSUBS 0.008093f
C202 B.n165 VSUBS 0.008093f
C203 B.n166 VSUBS 0.008093f
C204 B.n167 VSUBS 0.008093f
C205 B.n168 VSUBS 0.008093f
C206 B.n169 VSUBS 0.008093f
C207 B.n170 VSUBS 0.008093f
C208 B.n171 VSUBS 0.008093f
C209 B.n172 VSUBS 0.008093f
C210 B.n173 VSUBS 0.008093f
C211 B.n174 VSUBS 0.008093f
C212 B.n175 VSUBS 0.008093f
C213 B.n176 VSUBS 0.008093f
C214 B.n177 VSUBS 0.008093f
C215 B.n178 VSUBS 0.008093f
C216 B.n179 VSUBS 0.008093f
C217 B.n180 VSUBS 0.008093f
C218 B.n181 VSUBS 0.008093f
C219 B.n182 VSUBS 0.008093f
C220 B.n183 VSUBS 0.008093f
C221 B.n184 VSUBS 0.008093f
C222 B.n185 VSUBS 0.017708f
C223 B.n186 VSUBS 0.019189f
C224 B.n187 VSUBS 0.019189f
C225 B.n188 VSUBS 0.008093f
C226 B.n189 VSUBS 0.008093f
C227 B.n190 VSUBS 0.008093f
C228 B.n191 VSUBS 0.008093f
C229 B.n192 VSUBS 0.008093f
C230 B.n193 VSUBS 0.008093f
C231 B.n194 VSUBS 0.008093f
C232 B.n195 VSUBS 0.008093f
C233 B.n196 VSUBS 0.008093f
C234 B.n197 VSUBS 0.008093f
C235 B.n198 VSUBS 0.008093f
C236 B.n199 VSUBS 0.008093f
C237 B.n200 VSUBS 0.008093f
C238 B.n201 VSUBS 0.008093f
C239 B.n202 VSUBS 0.008093f
C240 B.n203 VSUBS 0.008093f
C241 B.n204 VSUBS 0.008093f
C242 B.n205 VSUBS 0.008093f
C243 B.n206 VSUBS 0.008093f
C244 B.n207 VSUBS 0.008093f
C245 B.n208 VSUBS 0.008093f
C246 B.n209 VSUBS 0.008093f
C247 B.n210 VSUBS 0.008093f
C248 B.n211 VSUBS 0.008093f
C249 B.n212 VSUBS 0.008093f
C250 B.n213 VSUBS 0.008093f
C251 B.n214 VSUBS 0.008093f
C252 B.n215 VSUBS 0.008093f
C253 B.n216 VSUBS 0.008093f
C254 B.n217 VSUBS 0.008093f
C255 B.n218 VSUBS 0.008093f
C256 B.n219 VSUBS 0.008093f
C257 B.n220 VSUBS 0.008093f
C258 B.n221 VSUBS 0.008093f
C259 B.n222 VSUBS 0.008093f
C260 B.n223 VSUBS 0.008093f
C261 B.n224 VSUBS 0.008093f
C262 B.n225 VSUBS 0.008093f
C263 B.n226 VSUBS 0.008093f
C264 B.n227 VSUBS 0.008093f
C265 B.n228 VSUBS 0.008093f
C266 B.n229 VSUBS 0.008093f
C267 B.n230 VSUBS 0.008093f
C268 B.n231 VSUBS 0.008093f
C269 B.n232 VSUBS 0.008093f
C270 B.n233 VSUBS 0.008093f
C271 B.n234 VSUBS 0.008093f
C272 B.n235 VSUBS 0.008093f
C273 B.n236 VSUBS 0.008093f
C274 B.n237 VSUBS 0.008093f
C275 B.n238 VSUBS 0.008093f
C276 B.n239 VSUBS 0.008093f
C277 B.n240 VSUBS 0.008093f
C278 B.n241 VSUBS 0.008093f
C279 B.n242 VSUBS 0.008093f
C280 B.n243 VSUBS 0.008093f
C281 B.n244 VSUBS 0.008093f
C282 B.n245 VSUBS 0.008093f
C283 B.n246 VSUBS 0.008093f
C284 B.n247 VSUBS 0.008093f
C285 B.n248 VSUBS 0.008093f
C286 B.n249 VSUBS 0.008093f
C287 B.n250 VSUBS 0.008093f
C288 B.n251 VSUBS 0.008093f
C289 B.n252 VSUBS 0.008093f
C290 B.n253 VSUBS 0.008093f
C291 B.n254 VSUBS 0.008093f
C292 B.n255 VSUBS 0.008093f
C293 B.n256 VSUBS 0.008093f
C294 B.n257 VSUBS 0.008093f
C295 B.t5 VSUBS 0.556908f
C296 B.t4 VSUBS 0.564878f
C297 B.t3 VSUBS 0.349486f
C298 B.n258 VSUBS 0.156745f
C299 B.n259 VSUBS 0.073214f
C300 B.n260 VSUBS 0.018752f
C301 B.n261 VSUBS 0.007617f
C302 B.n262 VSUBS 0.008093f
C303 B.n263 VSUBS 0.008093f
C304 B.n264 VSUBS 0.008093f
C305 B.n265 VSUBS 0.008093f
C306 B.n266 VSUBS 0.008093f
C307 B.n267 VSUBS 0.008093f
C308 B.n268 VSUBS 0.008093f
C309 B.n269 VSUBS 0.008093f
C310 B.n270 VSUBS 0.008093f
C311 B.n271 VSUBS 0.008093f
C312 B.n272 VSUBS 0.008093f
C313 B.n273 VSUBS 0.008093f
C314 B.n274 VSUBS 0.008093f
C315 B.n275 VSUBS 0.008093f
C316 B.n276 VSUBS 0.008093f
C317 B.n277 VSUBS 0.004523f
C318 B.n278 VSUBS 0.018752f
C319 B.n279 VSUBS 0.007617f
C320 B.n280 VSUBS 0.008093f
C321 B.n281 VSUBS 0.008093f
C322 B.n282 VSUBS 0.008093f
C323 B.n283 VSUBS 0.008093f
C324 B.n284 VSUBS 0.008093f
C325 B.n285 VSUBS 0.008093f
C326 B.n286 VSUBS 0.008093f
C327 B.n287 VSUBS 0.008093f
C328 B.n288 VSUBS 0.008093f
C329 B.n289 VSUBS 0.008093f
C330 B.n290 VSUBS 0.008093f
C331 B.n291 VSUBS 0.008093f
C332 B.n292 VSUBS 0.008093f
C333 B.n293 VSUBS 0.008093f
C334 B.n294 VSUBS 0.008093f
C335 B.n295 VSUBS 0.008093f
C336 B.n296 VSUBS 0.008093f
C337 B.n297 VSUBS 0.008093f
C338 B.n298 VSUBS 0.008093f
C339 B.n299 VSUBS 0.008093f
C340 B.n300 VSUBS 0.008093f
C341 B.n301 VSUBS 0.008093f
C342 B.n302 VSUBS 0.008093f
C343 B.n303 VSUBS 0.008093f
C344 B.n304 VSUBS 0.008093f
C345 B.n305 VSUBS 0.008093f
C346 B.n306 VSUBS 0.008093f
C347 B.n307 VSUBS 0.008093f
C348 B.n308 VSUBS 0.008093f
C349 B.n309 VSUBS 0.008093f
C350 B.n310 VSUBS 0.008093f
C351 B.n311 VSUBS 0.008093f
C352 B.n312 VSUBS 0.008093f
C353 B.n313 VSUBS 0.008093f
C354 B.n314 VSUBS 0.008093f
C355 B.n315 VSUBS 0.008093f
C356 B.n316 VSUBS 0.008093f
C357 B.n317 VSUBS 0.008093f
C358 B.n318 VSUBS 0.008093f
C359 B.n319 VSUBS 0.008093f
C360 B.n320 VSUBS 0.008093f
C361 B.n321 VSUBS 0.008093f
C362 B.n322 VSUBS 0.008093f
C363 B.n323 VSUBS 0.008093f
C364 B.n324 VSUBS 0.008093f
C365 B.n325 VSUBS 0.008093f
C366 B.n326 VSUBS 0.008093f
C367 B.n327 VSUBS 0.008093f
C368 B.n328 VSUBS 0.008093f
C369 B.n329 VSUBS 0.008093f
C370 B.n330 VSUBS 0.008093f
C371 B.n331 VSUBS 0.008093f
C372 B.n332 VSUBS 0.008093f
C373 B.n333 VSUBS 0.008093f
C374 B.n334 VSUBS 0.008093f
C375 B.n335 VSUBS 0.008093f
C376 B.n336 VSUBS 0.008093f
C377 B.n337 VSUBS 0.008093f
C378 B.n338 VSUBS 0.008093f
C379 B.n339 VSUBS 0.008093f
C380 B.n340 VSUBS 0.008093f
C381 B.n341 VSUBS 0.008093f
C382 B.n342 VSUBS 0.008093f
C383 B.n343 VSUBS 0.008093f
C384 B.n344 VSUBS 0.008093f
C385 B.n345 VSUBS 0.008093f
C386 B.n346 VSUBS 0.008093f
C387 B.n347 VSUBS 0.008093f
C388 B.n348 VSUBS 0.008093f
C389 B.n349 VSUBS 0.008093f
C390 B.n350 VSUBS 0.008093f
C391 B.n351 VSUBS 0.018193f
C392 B.n352 VSUBS 0.018703f
C393 B.n353 VSUBS 0.017708f
C394 B.n354 VSUBS 0.008093f
C395 B.n355 VSUBS 0.008093f
C396 B.n356 VSUBS 0.008093f
C397 B.n357 VSUBS 0.008093f
C398 B.n358 VSUBS 0.008093f
C399 B.n359 VSUBS 0.008093f
C400 B.n360 VSUBS 0.008093f
C401 B.n361 VSUBS 0.008093f
C402 B.n362 VSUBS 0.008093f
C403 B.n363 VSUBS 0.008093f
C404 B.n364 VSUBS 0.008093f
C405 B.n365 VSUBS 0.008093f
C406 B.n366 VSUBS 0.008093f
C407 B.n367 VSUBS 0.008093f
C408 B.n368 VSUBS 0.008093f
C409 B.n369 VSUBS 0.008093f
C410 B.n370 VSUBS 0.008093f
C411 B.n371 VSUBS 0.008093f
C412 B.n372 VSUBS 0.008093f
C413 B.n373 VSUBS 0.008093f
C414 B.n374 VSUBS 0.008093f
C415 B.n375 VSUBS 0.008093f
C416 B.n376 VSUBS 0.008093f
C417 B.n377 VSUBS 0.008093f
C418 B.n378 VSUBS 0.008093f
C419 B.n379 VSUBS 0.008093f
C420 B.n380 VSUBS 0.008093f
C421 B.n381 VSUBS 0.008093f
C422 B.n382 VSUBS 0.008093f
C423 B.n383 VSUBS 0.008093f
C424 B.n384 VSUBS 0.008093f
C425 B.n385 VSUBS 0.008093f
C426 B.n386 VSUBS 0.008093f
C427 B.n387 VSUBS 0.008093f
C428 B.n388 VSUBS 0.008093f
C429 B.n389 VSUBS 0.008093f
C430 B.n390 VSUBS 0.008093f
C431 B.n391 VSUBS 0.008093f
C432 B.n392 VSUBS 0.008093f
C433 B.n393 VSUBS 0.008093f
C434 B.n394 VSUBS 0.008093f
C435 B.n395 VSUBS 0.008093f
C436 B.n396 VSUBS 0.008093f
C437 B.n397 VSUBS 0.008093f
C438 B.n398 VSUBS 0.008093f
C439 B.n399 VSUBS 0.008093f
C440 B.n400 VSUBS 0.008093f
C441 B.n401 VSUBS 0.008093f
C442 B.n402 VSUBS 0.008093f
C443 B.n403 VSUBS 0.008093f
C444 B.n404 VSUBS 0.008093f
C445 B.n405 VSUBS 0.008093f
C446 B.n406 VSUBS 0.008093f
C447 B.n407 VSUBS 0.008093f
C448 B.n408 VSUBS 0.008093f
C449 B.n409 VSUBS 0.008093f
C450 B.n410 VSUBS 0.008093f
C451 B.n411 VSUBS 0.008093f
C452 B.n412 VSUBS 0.008093f
C453 B.n413 VSUBS 0.008093f
C454 B.n414 VSUBS 0.017708f
C455 B.n415 VSUBS 0.019189f
C456 B.n416 VSUBS 0.019189f
C457 B.n417 VSUBS 0.008093f
C458 B.n418 VSUBS 0.008093f
C459 B.n419 VSUBS 0.008093f
C460 B.n420 VSUBS 0.008093f
C461 B.n421 VSUBS 0.008093f
C462 B.n422 VSUBS 0.008093f
C463 B.n423 VSUBS 0.008093f
C464 B.n424 VSUBS 0.008093f
C465 B.n425 VSUBS 0.008093f
C466 B.n426 VSUBS 0.008093f
C467 B.n427 VSUBS 0.008093f
C468 B.n428 VSUBS 0.008093f
C469 B.n429 VSUBS 0.008093f
C470 B.n430 VSUBS 0.008093f
C471 B.n431 VSUBS 0.008093f
C472 B.n432 VSUBS 0.008093f
C473 B.n433 VSUBS 0.008093f
C474 B.n434 VSUBS 0.008093f
C475 B.n435 VSUBS 0.008093f
C476 B.n436 VSUBS 0.008093f
C477 B.n437 VSUBS 0.008093f
C478 B.n438 VSUBS 0.008093f
C479 B.n439 VSUBS 0.008093f
C480 B.n440 VSUBS 0.008093f
C481 B.n441 VSUBS 0.008093f
C482 B.n442 VSUBS 0.008093f
C483 B.n443 VSUBS 0.008093f
C484 B.n444 VSUBS 0.008093f
C485 B.n445 VSUBS 0.008093f
C486 B.n446 VSUBS 0.008093f
C487 B.n447 VSUBS 0.008093f
C488 B.n448 VSUBS 0.008093f
C489 B.n449 VSUBS 0.008093f
C490 B.n450 VSUBS 0.008093f
C491 B.n451 VSUBS 0.008093f
C492 B.n452 VSUBS 0.008093f
C493 B.n453 VSUBS 0.008093f
C494 B.n454 VSUBS 0.008093f
C495 B.n455 VSUBS 0.008093f
C496 B.n456 VSUBS 0.008093f
C497 B.n457 VSUBS 0.008093f
C498 B.n458 VSUBS 0.008093f
C499 B.n459 VSUBS 0.008093f
C500 B.n460 VSUBS 0.008093f
C501 B.n461 VSUBS 0.008093f
C502 B.n462 VSUBS 0.008093f
C503 B.n463 VSUBS 0.008093f
C504 B.n464 VSUBS 0.008093f
C505 B.n465 VSUBS 0.008093f
C506 B.n466 VSUBS 0.008093f
C507 B.n467 VSUBS 0.008093f
C508 B.n468 VSUBS 0.008093f
C509 B.n469 VSUBS 0.008093f
C510 B.n470 VSUBS 0.008093f
C511 B.n471 VSUBS 0.008093f
C512 B.n472 VSUBS 0.008093f
C513 B.n473 VSUBS 0.008093f
C514 B.n474 VSUBS 0.008093f
C515 B.n475 VSUBS 0.008093f
C516 B.n476 VSUBS 0.008093f
C517 B.n477 VSUBS 0.008093f
C518 B.n478 VSUBS 0.008093f
C519 B.n479 VSUBS 0.008093f
C520 B.n480 VSUBS 0.008093f
C521 B.n481 VSUBS 0.008093f
C522 B.n482 VSUBS 0.008093f
C523 B.n483 VSUBS 0.008093f
C524 B.n484 VSUBS 0.008093f
C525 B.n485 VSUBS 0.008093f
C526 B.n486 VSUBS 0.008093f
C527 B.n487 VSUBS 0.008093f
C528 B.n488 VSUBS 0.007617f
C529 B.n489 VSUBS 0.018752f
C530 B.n490 VSUBS 0.004523f
C531 B.n491 VSUBS 0.008093f
C532 B.n492 VSUBS 0.008093f
C533 B.n493 VSUBS 0.008093f
C534 B.n494 VSUBS 0.008093f
C535 B.n495 VSUBS 0.008093f
C536 B.n496 VSUBS 0.008093f
C537 B.n497 VSUBS 0.008093f
C538 B.n498 VSUBS 0.008093f
C539 B.n499 VSUBS 0.008093f
C540 B.n500 VSUBS 0.008093f
C541 B.n501 VSUBS 0.008093f
C542 B.n502 VSUBS 0.008093f
C543 B.n503 VSUBS 0.004523f
C544 B.n504 VSUBS 0.008093f
C545 B.n505 VSUBS 0.008093f
C546 B.n506 VSUBS 0.008093f
C547 B.n507 VSUBS 0.008093f
C548 B.n508 VSUBS 0.008093f
C549 B.n509 VSUBS 0.008093f
C550 B.n510 VSUBS 0.008093f
C551 B.n511 VSUBS 0.008093f
C552 B.n512 VSUBS 0.008093f
C553 B.n513 VSUBS 0.008093f
C554 B.n514 VSUBS 0.008093f
C555 B.n515 VSUBS 0.008093f
C556 B.n516 VSUBS 0.008093f
C557 B.n517 VSUBS 0.008093f
C558 B.n518 VSUBS 0.008093f
C559 B.n519 VSUBS 0.008093f
C560 B.n520 VSUBS 0.008093f
C561 B.n521 VSUBS 0.008093f
C562 B.n522 VSUBS 0.008093f
C563 B.n523 VSUBS 0.008093f
C564 B.n524 VSUBS 0.008093f
C565 B.n525 VSUBS 0.008093f
C566 B.n526 VSUBS 0.008093f
C567 B.n527 VSUBS 0.008093f
C568 B.n528 VSUBS 0.008093f
C569 B.n529 VSUBS 0.008093f
C570 B.n530 VSUBS 0.008093f
C571 B.n531 VSUBS 0.008093f
C572 B.n532 VSUBS 0.008093f
C573 B.n533 VSUBS 0.008093f
C574 B.n534 VSUBS 0.008093f
C575 B.n535 VSUBS 0.008093f
C576 B.n536 VSUBS 0.008093f
C577 B.n537 VSUBS 0.008093f
C578 B.n538 VSUBS 0.008093f
C579 B.n539 VSUBS 0.008093f
C580 B.n540 VSUBS 0.008093f
C581 B.n541 VSUBS 0.008093f
C582 B.n542 VSUBS 0.008093f
C583 B.n543 VSUBS 0.008093f
C584 B.n544 VSUBS 0.008093f
C585 B.n545 VSUBS 0.008093f
C586 B.n546 VSUBS 0.008093f
C587 B.n547 VSUBS 0.008093f
C588 B.n548 VSUBS 0.008093f
C589 B.n549 VSUBS 0.008093f
C590 B.n550 VSUBS 0.008093f
C591 B.n551 VSUBS 0.008093f
C592 B.n552 VSUBS 0.008093f
C593 B.n553 VSUBS 0.008093f
C594 B.n554 VSUBS 0.008093f
C595 B.n555 VSUBS 0.008093f
C596 B.n556 VSUBS 0.008093f
C597 B.n557 VSUBS 0.008093f
C598 B.n558 VSUBS 0.008093f
C599 B.n559 VSUBS 0.008093f
C600 B.n560 VSUBS 0.008093f
C601 B.n561 VSUBS 0.008093f
C602 B.n562 VSUBS 0.008093f
C603 B.n563 VSUBS 0.008093f
C604 B.n564 VSUBS 0.008093f
C605 B.n565 VSUBS 0.008093f
C606 B.n566 VSUBS 0.008093f
C607 B.n567 VSUBS 0.008093f
C608 B.n568 VSUBS 0.008093f
C609 B.n569 VSUBS 0.008093f
C610 B.n570 VSUBS 0.008093f
C611 B.n571 VSUBS 0.008093f
C612 B.n572 VSUBS 0.008093f
C613 B.n573 VSUBS 0.008093f
C614 B.n574 VSUBS 0.008093f
C615 B.n575 VSUBS 0.008093f
C616 B.n576 VSUBS 0.008093f
C617 B.n577 VSUBS 0.019189f
C618 B.n578 VSUBS 0.017708f
C619 B.n579 VSUBS 0.017708f
C620 B.n580 VSUBS 0.008093f
C621 B.n581 VSUBS 0.008093f
C622 B.n582 VSUBS 0.008093f
C623 B.n583 VSUBS 0.008093f
C624 B.n584 VSUBS 0.008093f
C625 B.n585 VSUBS 0.008093f
C626 B.n586 VSUBS 0.008093f
C627 B.n587 VSUBS 0.008093f
C628 B.n588 VSUBS 0.008093f
C629 B.n589 VSUBS 0.008093f
C630 B.n590 VSUBS 0.008093f
C631 B.n591 VSUBS 0.008093f
C632 B.n592 VSUBS 0.008093f
C633 B.n593 VSUBS 0.008093f
C634 B.n594 VSUBS 0.008093f
C635 B.n595 VSUBS 0.008093f
C636 B.n596 VSUBS 0.008093f
C637 B.n597 VSUBS 0.008093f
C638 B.n598 VSUBS 0.008093f
C639 B.n599 VSUBS 0.008093f
C640 B.n600 VSUBS 0.008093f
C641 B.n601 VSUBS 0.008093f
C642 B.n602 VSUBS 0.008093f
C643 B.n603 VSUBS 0.008093f
C644 B.n604 VSUBS 0.008093f
C645 B.n605 VSUBS 0.008093f
C646 B.n606 VSUBS 0.008093f
C647 B.n607 VSUBS 0.010561f
C648 B.n608 VSUBS 0.011251f
C649 B.n609 VSUBS 0.022373f
C650 VDD1.t4 VSUBS 0.333019f
C651 VDD1.t1 VSUBS 0.333019f
C652 VDD1.n0 VSUBS 2.71182f
C653 VDD1.t7 VSUBS 0.333019f
C654 VDD1.t5 VSUBS 0.333019f
C655 VDD1.n1 VSUBS 2.71081f
C656 VDD1.t6 VSUBS 0.333019f
C657 VDD1.t2 VSUBS 0.333019f
C658 VDD1.n2 VSUBS 2.71081f
C659 VDD1.n3 VSUBS 3.23124f
C660 VDD1.t3 VSUBS 0.333019f
C661 VDD1.t0 VSUBS 0.333019f
C662 VDD1.n4 VSUBS 2.70815f
C663 VDD1.n5 VSUBS 3.14362f
C664 VP.n0 VSUBS 0.059295f
C665 VP.t2 VSUBS 1.27223f
C666 VP.n1 VSUBS 0.503119f
C667 VP.n2 VSUBS 0.059295f
C668 VP.t4 VSUBS 1.27223f
C669 VP.t6 VSUBS 1.27223f
C670 VP.n3 VSUBS 0.503119f
C671 VP.t3 VSUBS 1.28663f
C672 VP.n4 VSUBS 0.484249f
C673 VP.n5 VSUBS 0.198256f
C674 VP.n6 VSUBS 0.013455f
C675 VP.n7 VSUBS 0.503119f
C676 VP.t7 VSUBS 1.27365f
C677 VP.n8 VSUBS 0.496769f
C678 VP.n9 VSUBS 2.56231f
C679 VP.t0 VSUBS 1.27365f
C680 VP.n10 VSUBS 0.496769f
C681 VP.n11 VSUBS 2.61167f
C682 VP.n12 VSUBS 0.059295f
C683 VP.n13 VSUBS 0.059295f
C684 VP.n14 VSUBS 0.013455f
C685 VP.t1 VSUBS 1.27223f
C686 VP.n15 VSUBS 0.503119f
C687 VP.t5 VSUBS 1.27365f
C688 VP.n16 VSUBS 0.496769f
C689 VP.n17 VSUBS 0.045951f
C690 VDD2.t0 VSUBS 0.334763f
C691 VDD2.t5 VSUBS 0.334763f
C692 VDD2.n0 VSUBS 2.725f
C693 VDD2.t2 VSUBS 0.334763f
C694 VDD2.t7 VSUBS 0.334763f
C695 VDD2.n1 VSUBS 2.725f
C696 VDD2.n2 VSUBS 3.18585f
C697 VDD2.t1 VSUBS 0.334763f
C698 VDD2.t4 VSUBS 0.334763f
C699 VDD2.n3 VSUBS 2.72234f
C700 VDD2.n4 VSUBS 3.12548f
C701 VDD2.t3 VSUBS 0.334763f
C702 VDD2.t6 VSUBS 0.334763f
C703 VDD2.n5 VSUBS 2.72496f
C704 VTAIL.t9 VSUBS 0.293444f
C705 VTAIL.t15 VSUBS 0.293444f
C706 VTAIL.n0 VSUBS 2.25418f
C707 VTAIL.n1 VSUBS 0.633547f
C708 VTAIL.t10 VSUBS 2.95318f
C709 VTAIL.n2 VSUBS 0.768792f
C710 VTAIL.t7 VSUBS 2.95318f
C711 VTAIL.n3 VSUBS 0.768792f
C712 VTAIL.t2 VSUBS 0.293444f
C713 VTAIL.t0 VSUBS 0.293444f
C714 VTAIL.n4 VSUBS 2.25418f
C715 VTAIL.n5 VSUBS 0.689174f
C716 VTAIL.t1 VSUBS 2.95318f
C717 VTAIL.n6 VSUBS 2.16961f
C718 VTAIL.t12 VSUBS 2.9532f
C719 VTAIL.n7 VSUBS 2.16959f
C720 VTAIL.t14 VSUBS 0.293444f
C721 VTAIL.t8 VSUBS 0.293444f
C722 VTAIL.n8 VSUBS 2.25418f
C723 VTAIL.n9 VSUBS 0.68917f
C724 VTAIL.t11 VSUBS 2.9532f
C725 VTAIL.n10 VSUBS 0.768769f
C726 VTAIL.t3 VSUBS 2.9532f
C727 VTAIL.n11 VSUBS 0.768769f
C728 VTAIL.t4 VSUBS 0.293444f
C729 VTAIL.t5 VSUBS 0.293444f
C730 VTAIL.n12 VSUBS 2.25418f
C731 VTAIL.n13 VSUBS 0.68917f
C732 VTAIL.t6 VSUBS 2.95318f
C733 VTAIL.n14 VSUBS 2.16961f
C734 VTAIL.t13 VSUBS 2.95318f
C735 VTAIL.n15 VSUBS 2.16481f
C736 VN.n0 VSUBS 0.058157f
C737 VN.t2 VSUBS 1.24783f
C738 VN.n1 VSUBS 0.493467f
C739 VN.t7 VSUBS 1.26195f
C740 VN.n2 VSUBS 0.47496f
C741 VN.n3 VSUBS 0.194452f
C742 VN.n4 VSUBS 0.013197f
C743 VN.t5 VSUBS 1.24783f
C744 VN.n5 VSUBS 0.493467f
C745 VN.t0 VSUBS 1.24921f
C746 VN.n6 VSUBS 0.487239f
C747 VN.n7 VSUBS 0.04507f
C748 VN.n8 VSUBS 0.058157f
C749 VN.t6 VSUBS 1.24921f
C750 VN.t4 VSUBS 1.24783f
C751 VN.n9 VSUBS 0.493467f
C752 VN.t1 VSUBS 1.26195f
C753 VN.n10 VSUBS 0.47496f
C754 VN.n11 VSUBS 0.194452f
C755 VN.n12 VSUBS 0.013197f
C756 VN.t3 VSUBS 1.24783f
C757 VN.n13 VSUBS 0.493467f
C758 VN.n14 VSUBS 0.487239f
C759 VN.n15 VSUBS 2.55127f
.ends

