* NGSPICE file created from diff_pair_sample_0529.ext - technology: sky130A

.subckt diff_pair_sample_0529 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t16 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.3366 pd=2.37 as=0.3366 ps=2.37 w=2.04 l=1.05
X1 B.t11 B.t9 B.t10 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.7956 pd=4.86 as=0 ps=0 w=2.04 l=1.05
X2 VTAIL.t6 VP.t0 VDD1.t9 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.3366 pd=2.37 as=0.3366 ps=2.37 w=2.04 l=1.05
X3 VTAIL.t1 VP.t1 VDD1.t8 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.3366 pd=2.37 as=0.3366 ps=2.37 w=2.04 l=1.05
X4 VDD2.t8 VN.t1 VTAIL.t14 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.3366 pd=2.37 as=0.7956 ps=4.86 w=2.04 l=1.05
X5 VDD1.t7 VP.t2 VTAIL.t8 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.3366 pd=2.37 as=0.3366 ps=2.37 w=2.04 l=1.05
X6 B.t8 B.t6 B.t7 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.7956 pd=4.86 as=0 ps=0 w=2.04 l=1.05
X7 VDD1.t6 VP.t3 VTAIL.t7 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.3366 pd=2.37 as=0.3366 ps=2.37 w=2.04 l=1.05
X8 B.t5 B.t3 B.t4 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.7956 pd=4.86 as=0 ps=0 w=2.04 l=1.05
X9 VTAIL.t19 VN.t2 VDD2.t7 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.3366 pd=2.37 as=0.3366 ps=2.37 w=2.04 l=1.05
X10 VTAIL.t10 VN.t3 VDD2.t6 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.3366 pd=2.37 as=0.3366 ps=2.37 w=2.04 l=1.05
X11 B.t2 B.t0 B.t1 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.7956 pd=4.86 as=0 ps=0 w=2.04 l=1.05
X12 VDD2.t5 VN.t4 VTAIL.t11 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.3366 pd=2.37 as=0.3366 ps=2.37 w=2.04 l=1.05
X13 VTAIL.t0 VP.t4 VDD1.t5 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.3366 pd=2.37 as=0.3366 ps=2.37 w=2.04 l=1.05
X14 VDD2.t4 VN.t5 VTAIL.t17 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.3366 pd=2.37 as=0.7956 ps=4.86 w=2.04 l=1.05
X15 VDD1.t4 VP.t5 VTAIL.t3 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.7956 pd=4.86 as=0.3366 ps=2.37 w=2.04 l=1.05
X16 VTAIL.t15 VN.t6 VDD2.t3 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.3366 pd=2.37 as=0.3366 ps=2.37 w=2.04 l=1.05
X17 VDD1.t3 VP.t6 VTAIL.t5 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.3366 pd=2.37 as=0.7956 ps=4.86 w=2.04 l=1.05
X18 VDD1.t2 VP.t7 VTAIL.t9 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.7956 pd=4.86 as=0.3366 ps=2.37 w=2.04 l=1.05
X19 VDD1.t1 VP.t8 VTAIL.t2 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.3366 pd=2.37 as=0.7956 ps=4.86 w=2.04 l=1.05
X20 VDD2.t2 VN.t7 VTAIL.t13 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.7956 pd=4.86 as=0.3366 ps=2.37 w=2.04 l=1.05
X21 VTAIL.t4 VP.t9 VDD1.t0 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.3366 pd=2.37 as=0.3366 ps=2.37 w=2.04 l=1.05
X22 VTAIL.t18 VN.t8 VDD2.t1 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.3366 pd=2.37 as=0.3366 ps=2.37 w=2.04 l=1.05
X23 VDD2.t0 VN.t9 VTAIL.t12 w_n2626_n1376# sky130_fd_pr__pfet_01v8 ad=0.7956 pd=4.86 as=0.3366 ps=2.37 w=2.04 l=1.05
R0 VN.n37 VN.n20 161.3
R1 VN.n35 VN.n34 161.3
R2 VN.n33 VN.n21 161.3
R3 VN.n32 VN.n31 161.3
R4 VN.n29 VN.n22 161.3
R5 VN.n28 VN.n27 161.3
R6 VN.n26 VN.n23 161.3
R7 VN.n17 VN.n0 161.3
R8 VN.n15 VN.n14 161.3
R9 VN.n13 VN.n1 161.3
R10 VN.n12 VN.n11 161.3
R11 VN.n9 VN.n2 161.3
R12 VN.n8 VN.n7 161.3
R13 VN.n6 VN.n3 161.3
R14 VN.n5 VN.t7 99.3881
R15 VN.n25 VN.t5 99.3881
R16 VN.n18 VN.t1 84.2357
R17 VN.n38 VN.t9 84.2357
R18 VN.n39 VN.n38 80.6037
R19 VN.n19 VN.n18 80.6037
R20 VN.n18 VN.n17 55.824
R21 VN.n38 VN.n37 55.824
R22 VN.n5 VN.n4 48.4137
R23 VN.n25 VN.n24 48.4137
R24 VN.n4 VN.t6 46.8234
R25 VN.n10 VN.t4 46.8234
R26 VN.n16 VN.t2 46.8234
R27 VN.n24 VN.t3 46.8234
R28 VN.n30 VN.t0 46.8234
R29 VN.n36 VN.t8 46.8234
R30 VN.n9 VN.n8 46.3896
R31 VN.n11 VN.n1 46.3896
R32 VN.n29 VN.n28 46.3896
R33 VN.n31 VN.n21 46.3896
R34 VN.n26 VN.n25 43.9713
R35 VN.n6 VN.n5 43.9713
R36 VN VN.n39 37.6657
R37 VN.n8 VN.n3 34.7644
R38 VN.n15 VN.n1 34.7644
R39 VN.n28 VN.n23 34.7644
R40 VN.n35 VN.n21 34.7644
R41 VN.n17 VN.n16 18.1985
R42 VN.n37 VN.n36 18.1985
R43 VN.n10 VN.n9 12.2964
R44 VN.n11 VN.n10 12.2964
R45 VN.n31 VN.n30 12.2964
R46 VN.n30 VN.n29 12.2964
R47 VN.n4 VN.n3 6.39438
R48 VN.n16 VN.n15 6.39438
R49 VN.n24 VN.n23 6.39438
R50 VN.n36 VN.n35 6.39438
R51 VN.n39 VN.n20 0.285035
R52 VN.n19 VN.n0 0.285035
R53 VN.n34 VN.n20 0.189894
R54 VN.n34 VN.n33 0.189894
R55 VN.n33 VN.n32 0.189894
R56 VN.n32 VN.n22 0.189894
R57 VN.n27 VN.n22 0.189894
R58 VN.n27 VN.n26 0.189894
R59 VN.n7 VN.n6 0.189894
R60 VN.n7 VN.n2 0.189894
R61 VN.n12 VN.n2 0.189894
R62 VN.n13 VN.n12 0.189894
R63 VN.n14 VN.n13 0.189894
R64 VN.n14 VN.n0 0.189894
R65 VN VN.n19 0.146778
R66 VTAIL.n17 VTAIL.t14 170.095
R67 VTAIL.n2 VTAIL.t5 170.095
R68 VTAIL.n16 VTAIL.t2 170.095
R69 VTAIL.n11 VTAIL.t17 170.095
R70 VTAIL.n15 VTAIL.n14 154.161
R71 VTAIL.n13 VTAIL.n12 154.161
R72 VTAIL.n10 VTAIL.n9 154.161
R73 VTAIL.n8 VTAIL.n7 154.161
R74 VTAIL.n19 VTAIL.n18 154.161
R75 VTAIL.n1 VTAIL.n0 154.161
R76 VTAIL.n4 VTAIL.n3 154.161
R77 VTAIL.n6 VTAIL.n5 154.161
R78 VTAIL.n8 VTAIL.n6 16.5048
R79 VTAIL.n18 VTAIL.t11 15.9343
R80 VTAIL.n18 VTAIL.t19 15.9343
R81 VTAIL.n0 VTAIL.t13 15.9343
R82 VTAIL.n0 VTAIL.t15 15.9343
R83 VTAIL.n3 VTAIL.t8 15.9343
R84 VTAIL.n3 VTAIL.t6 15.9343
R85 VTAIL.n5 VTAIL.t9 15.9343
R86 VTAIL.n5 VTAIL.t1 15.9343
R87 VTAIL.n14 VTAIL.t7 15.9343
R88 VTAIL.n14 VTAIL.t4 15.9343
R89 VTAIL.n12 VTAIL.t3 15.9343
R90 VTAIL.n12 VTAIL.t0 15.9343
R91 VTAIL.n9 VTAIL.t16 15.9343
R92 VTAIL.n9 VTAIL.t10 15.9343
R93 VTAIL.n7 VTAIL.t12 15.9343
R94 VTAIL.n7 VTAIL.t18 15.9343
R95 VTAIL.n17 VTAIL.n16 15.3152
R96 VTAIL.n10 VTAIL.n8 1.19016
R97 VTAIL.n11 VTAIL.n10 1.19016
R98 VTAIL.n15 VTAIL.n13 1.19016
R99 VTAIL.n16 VTAIL.n15 1.19016
R100 VTAIL.n6 VTAIL.n4 1.19016
R101 VTAIL.n4 VTAIL.n2 1.19016
R102 VTAIL.n19 VTAIL.n17 1.19016
R103 VTAIL.n13 VTAIL.n11 1.06516
R104 VTAIL.n2 VTAIL.n1 1.06516
R105 VTAIL VTAIL.n1 0.950931
R106 VTAIL VTAIL.n19 0.239724
R107 VDD2.n1 VDD2.t2 187.963
R108 VDD2.n4 VDD2.t0 186.774
R109 VDD2.n3 VDD2.n2 171.677
R110 VDD2 VDD2.n7 171.673
R111 VDD2.n6 VDD2.n5 170.839
R112 VDD2.n1 VDD2.n0 170.839
R113 VDD2.n4 VDD2.n3 31.1248
R114 VDD2.n7 VDD2.t6 15.9343
R115 VDD2.n7 VDD2.t4 15.9343
R116 VDD2.n5 VDD2.t1 15.9343
R117 VDD2.n5 VDD2.t9 15.9343
R118 VDD2.n2 VDD2.t7 15.9343
R119 VDD2.n2 VDD2.t8 15.9343
R120 VDD2.n0 VDD2.t3 15.9343
R121 VDD2.n0 VDD2.t5 15.9343
R122 VDD2.n6 VDD2.n4 1.19016
R123 VDD2 VDD2.n6 0.356103
R124 VDD2.n3 VDD2.n1 0.242568
R125 B.n208 B.n207 585
R126 B.n206 B.n73 585
R127 B.n205 B.n204 585
R128 B.n203 B.n74 585
R129 B.n202 B.n201 585
R130 B.n200 B.n75 585
R131 B.n199 B.n198 585
R132 B.n197 B.n76 585
R133 B.n196 B.n195 585
R134 B.n194 B.n77 585
R135 B.n193 B.n192 585
R136 B.n191 B.n78 585
R137 B.n190 B.n189 585
R138 B.n185 B.n79 585
R139 B.n184 B.n183 585
R140 B.n182 B.n80 585
R141 B.n181 B.n180 585
R142 B.n179 B.n81 585
R143 B.n178 B.n177 585
R144 B.n176 B.n82 585
R145 B.n175 B.n174 585
R146 B.n173 B.n83 585
R147 B.n171 B.n170 585
R148 B.n169 B.n86 585
R149 B.n168 B.n167 585
R150 B.n166 B.n87 585
R151 B.n165 B.n164 585
R152 B.n163 B.n88 585
R153 B.n162 B.n161 585
R154 B.n160 B.n89 585
R155 B.n159 B.n158 585
R156 B.n157 B.n90 585
R157 B.n156 B.n155 585
R158 B.n154 B.n91 585
R159 B.n209 B.n72 585
R160 B.n211 B.n210 585
R161 B.n212 B.n71 585
R162 B.n214 B.n213 585
R163 B.n215 B.n70 585
R164 B.n217 B.n216 585
R165 B.n218 B.n69 585
R166 B.n220 B.n219 585
R167 B.n221 B.n68 585
R168 B.n223 B.n222 585
R169 B.n224 B.n67 585
R170 B.n226 B.n225 585
R171 B.n227 B.n66 585
R172 B.n229 B.n228 585
R173 B.n230 B.n65 585
R174 B.n232 B.n231 585
R175 B.n233 B.n64 585
R176 B.n235 B.n234 585
R177 B.n236 B.n63 585
R178 B.n238 B.n237 585
R179 B.n239 B.n62 585
R180 B.n241 B.n240 585
R181 B.n242 B.n61 585
R182 B.n244 B.n243 585
R183 B.n245 B.n60 585
R184 B.n247 B.n246 585
R185 B.n248 B.n59 585
R186 B.n250 B.n249 585
R187 B.n251 B.n58 585
R188 B.n253 B.n252 585
R189 B.n254 B.n57 585
R190 B.n256 B.n255 585
R191 B.n257 B.n56 585
R192 B.n259 B.n258 585
R193 B.n260 B.n55 585
R194 B.n262 B.n261 585
R195 B.n263 B.n54 585
R196 B.n265 B.n264 585
R197 B.n266 B.n53 585
R198 B.n268 B.n267 585
R199 B.n269 B.n52 585
R200 B.n271 B.n270 585
R201 B.n272 B.n51 585
R202 B.n274 B.n273 585
R203 B.n275 B.n50 585
R204 B.n277 B.n276 585
R205 B.n278 B.n49 585
R206 B.n280 B.n279 585
R207 B.n281 B.n48 585
R208 B.n283 B.n282 585
R209 B.n284 B.n47 585
R210 B.n286 B.n285 585
R211 B.n287 B.n46 585
R212 B.n289 B.n288 585
R213 B.n290 B.n45 585
R214 B.n292 B.n291 585
R215 B.n293 B.n44 585
R216 B.n295 B.n294 585
R217 B.n296 B.n43 585
R218 B.n298 B.n297 585
R219 B.n299 B.n42 585
R220 B.n301 B.n300 585
R221 B.n302 B.n41 585
R222 B.n304 B.n303 585
R223 B.n305 B.n40 585
R224 B.n307 B.n306 585
R225 B.n359 B.n18 585
R226 B.n358 B.n357 585
R227 B.n356 B.n19 585
R228 B.n355 B.n354 585
R229 B.n353 B.n20 585
R230 B.n352 B.n351 585
R231 B.n350 B.n21 585
R232 B.n349 B.n348 585
R233 B.n347 B.n22 585
R234 B.n346 B.n345 585
R235 B.n344 B.n23 585
R236 B.n343 B.n342 585
R237 B.n341 B.n340 585
R238 B.n339 B.n27 585
R239 B.n338 B.n337 585
R240 B.n336 B.n28 585
R241 B.n335 B.n334 585
R242 B.n333 B.n29 585
R243 B.n332 B.n331 585
R244 B.n330 B.n30 585
R245 B.n329 B.n328 585
R246 B.n327 B.n31 585
R247 B.n325 B.n324 585
R248 B.n323 B.n34 585
R249 B.n322 B.n321 585
R250 B.n320 B.n35 585
R251 B.n319 B.n318 585
R252 B.n317 B.n36 585
R253 B.n316 B.n315 585
R254 B.n314 B.n37 585
R255 B.n313 B.n312 585
R256 B.n311 B.n38 585
R257 B.n310 B.n309 585
R258 B.n308 B.n39 585
R259 B.n361 B.n360 585
R260 B.n362 B.n17 585
R261 B.n364 B.n363 585
R262 B.n365 B.n16 585
R263 B.n367 B.n366 585
R264 B.n368 B.n15 585
R265 B.n370 B.n369 585
R266 B.n371 B.n14 585
R267 B.n373 B.n372 585
R268 B.n374 B.n13 585
R269 B.n376 B.n375 585
R270 B.n377 B.n12 585
R271 B.n379 B.n378 585
R272 B.n380 B.n11 585
R273 B.n382 B.n381 585
R274 B.n383 B.n10 585
R275 B.n385 B.n384 585
R276 B.n386 B.n9 585
R277 B.n388 B.n387 585
R278 B.n389 B.n8 585
R279 B.n391 B.n390 585
R280 B.n392 B.n7 585
R281 B.n394 B.n393 585
R282 B.n395 B.n6 585
R283 B.n397 B.n396 585
R284 B.n398 B.n5 585
R285 B.n400 B.n399 585
R286 B.n401 B.n4 585
R287 B.n403 B.n402 585
R288 B.n404 B.n3 585
R289 B.n406 B.n405 585
R290 B.n407 B.n0 585
R291 B.n2 B.n1 585
R292 B.n108 B.n107 585
R293 B.n109 B.n106 585
R294 B.n111 B.n110 585
R295 B.n112 B.n105 585
R296 B.n114 B.n113 585
R297 B.n115 B.n104 585
R298 B.n117 B.n116 585
R299 B.n118 B.n103 585
R300 B.n120 B.n119 585
R301 B.n121 B.n102 585
R302 B.n123 B.n122 585
R303 B.n124 B.n101 585
R304 B.n126 B.n125 585
R305 B.n127 B.n100 585
R306 B.n129 B.n128 585
R307 B.n130 B.n99 585
R308 B.n132 B.n131 585
R309 B.n133 B.n98 585
R310 B.n135 B.n134 585
R311 B.n136 B.n97 585
R312 B.n138 B.n137 585
R313 B.n139 B.n96 585
R314 B.n141 B.n140 585
R315 B.n142 B.n95 585
R316 B.n144 B.n143 585
R317 B.n145 B.n94 585
R318 B.n147 B.n146 585
R319 B.n148 B.n93 585
R320 B.n150 B.n149 585
R321 B.n151 B.n92 585
R322 B.n153 B.n152 585
R323 B.n152 B.n91 511.721
R324 B.n209 B.n208 511.721
R325 B.n306 B.n39 511.721
R326 B.n360 B.n359 511.721
R327 B.n409 B.n408 256.663
R328 B.n84 B.t6 250.077
R329 B.n186 B.t3 250.077
R330 B.n32 B.t9 250.077
R331 B.n24 B.t0 250.077
R332 B.n408 B.n407 235.042
R333 B.n408 B.n2 235.042
R334 B.n186 B.t4 197.667
R335 B.n32 B.t11 197.667
R336 B.n84 B.t7 197.667
R337 B.n24 B.t2 197.667
R338 B.n187 B.t5 170.904
R339 B.n33 B.t10 170.904
R340 B.n85 B.t8 170.904
R341 B.n25 B.t1 170.904
R342 B.n156 B.n91 163.367
R343 B.n157 B.n156 163.367
R344 B.n158 B.n157 163.367
R345 B.n158 B.n89 163.367
R346 B.n162 B.n89 163.367
R347 B.n163 B.n162 163.367
R348 B.n164 B.n163 163.367
R349 B.n164 B.n87 163.367
R350 B.n168 B.n87 163.367
R351 B.n169 B.n168 163.367
R352 B.n170 B.n169 163.367
R353 B.n170 B.n83 163.367
R354 B.n175 B.n83 163.367
R355 B.n176 B.n175 163.367
R356 B.n177 B.n176 163.367
R357 B.n177 B.n81 163.367
R358 B.n181 B.n81 163.367
R359 B.n182 B.n181 163.367
R360 B.n183 B.n182 163.367
R361 B.n183 B.n79 163.367
R362 B.n190 B.n79 163.367
R363 B.n191 B.n190 163.367
R364 B.n192 B.n191 163.367
R365 B.n192 B.n77 163.367
R366 B.n196 B.n77 163.367
R367 B.n197 B.n196 163.367
R368 B.n198 B.n197 163.367
R369 B.n198 B.n75 163.367
R370 B.n202 B.n75 163.367
R371 B.n203 B.n202 163.367
R372 B.n204 B.n203 163.367
R373 B.n204 B.n73 163.367
R374 B.n208 B.n73 163.367
R375 B.n306 B.n305 163.367
R376 B.n305 B.n304 163.367
R377 B.n304 B.n41 163.367
R378 B.n300 B.n41 163.367
R379 B.n300 B.n299 163.367
R380 B.n299 B.n298 163.367
R381 B.n298 B.n43 163.367
R382 B.n294 B.n43 163.367
R383 B.n294 B.n293 163.367
R384 B.n293 B.n292 163.367
R385 B.n292 B.n45 163.367
R386 B.n288 B.n45 163.367
R387 B.n288 B.n287 163.367
R388 B.n287 B.n286 163.367
R389 B.n286 B.n47 163.367
R390 B.n282 B.n47 163.367
R391 B.n282 B.n281 163.367
R392 B.n281 B.n280 163.367
R393 B.n280 B.n49 163.367
R394 B.n276 B.n49 163.367
R395 B.n276 B.n275 163.367
R396 B.n275 B.n274 163.367
R397 B.n274 B.n51 163.367
R398 B.n270 B.n51 163.367
R399 B.n270 B.n269 163.367
R400 B.n269 B.n268 163.367
R401 B.n268 B.n53 163.367
R402 B.n264 B.n53 163.367
R403 B.n264 B.n263 163.367
R404 B.n263 B.n262 163.367
R405 B.n262 B.n55 163.367
R406 B.n258 B.n55 163.367
R407 B.n258 B.n257 163.367
R408 B.n257 B.n256 163.367
R409 B.n256 B.n57 163.367
R410 B.n252 B.n57 163.367
R411 B.n252 B.n251 163.367
R412 B.n251 B.n250 163.367
R413 B.n250 B.n59 163.367
R414 B.n246 B.n59 163.367
R415 B.n246 B.n245 163.367
R416 B.n245 B.n244 163.367
R417 B.n244 B.n61 163.367
R418 B.n240 B.n61 163.367
R419 B.n240 B.n239 163.367
R420 B.n239 B.n238 163.367
R421 B.n238 B.n63 163.367
R422 B.n234 B.n63 163.367
R423 B.n234 B.n233 163.367
R424 B.n233 B.n232 163.367
R425 B.n232 B.n65 163.367
R426 B.n228 B.n65 163.367
R427 B.n228 B.n227 163.367
R428 B.n227 B.n226 163.367
R429 B.n226 B.n67 163.367
R430 B.n222 B.n67 163.367
R431 B.n222 B.n221 163.367
R432 B.n221 B.n220 163.367
R433 B.n220 B.n69 163.367
R434 B.n216 B.n69 163.367
R435 B.n216 B.n215 163.367
R436 B.n215 B.n214 163.367
R437 B.n214 B.n71 163.367
R438 B.n210 B.n71 163.367
R439 B.n210 B.n209 163.367
R440 B.n359 B.n358 163.367
R441 B.n358 B.n19 163.367
R442 B.n354 B.n19 163.367
R443 B.n354 B.n353 163.367
R444 B.n353 B.n352 163.367
R445 B.n352 B.n21 163.367
R446 B.n348 B.n21 163.367
R447 B.n348 B.n347 163.367
R448 B.n347 B.n346 163.367
R449 B.n346 B.n23 163.367
R450 B.n342 B.n23 163.367
R451 B.n342 B.n341 163.367
R452 B.n341 B.n27 163.367
R453 B.n337 B.n27 163.367
R454 B.n337 B.n336 163.367
R455 B.n336 B.n335 163.367
R456 B.n335 B.n29 163.367
R457 B.n331 B.n29 163.367
R458 B.n331 B.n330 163.367
R459 B.n330 B.n329 163.367
R460 B.n329 B.n31 163.367
R461 B.n324 B.n31 163.367
R462 B.n324 B.n323 163.367
R463 B.n323 B.n322 163.367
R464 B.n322 B.n35 163.367
R465 B.n318 B.n35 163.367
R466 B.n318 B.n317 163.367
R467 B.n317 B.n316 163.367
R468 B.n316 B.n37 163.367
R469 B.n312 B.n37 163.367
R470 B.n312 B.n311 163.367
R471 B.n311 B.n310 163.367
R472 B.n310 B.n39 163.367
R473 B.n360 B.n17 163.367
R474 B.n364 B.n17 163.367
R475 B.n365 B.n364 163.367
R476 B.n366 B.n365 163.367
R477 B.n366 B.n15 163.367
R478 B.n370 B.n15 163.367
R479 B.n371 B.n370 163.367
R480 B.n372 B.n371 163.367
R481 B.n372 B.n13 163.367
R482 B.n376 B.n13 163.367
R483 B.n377 B.n376 163.367
R484 B.n378 B.n377 163.367
R485 B.n378 B.n11 163.367
R486 B.n382 B.n11 163.367
R487 B.n383 B.n382 163.367
R488 B.n384 B.n383 163.367
R489 B.n384 B.n9 163.367
R490 B.n388 B.n9 163.367
R491 B.n389 B.n388 163.367
R492 B.n390 B.n389 163.367
R493 B.n390 B.n7 163.367
R494 B.n394 B.n7 163.367
R495 B.n395 B.n394 163.367
R496 B.n396 B.n395 163.367
R497 B.n396 B.n5 163.367
R498 B.n400 B.n5 163.367
R499 B.n401 B.n400 163.367
R500 B.n402 B.n401 163.367
R501 B.n402 B.n3 163.367
R502 B.n406 B.n3 163.367
R503 B.n407 B.n406 163.367
R504 B.n108 B.n2 163.367
R505 B.n109 B.n108 163.367
R506 B.n110 B.n109 163.367
R507 B.n110 B.n105 163.367
R508 B.n114 B.n105 163.367
R509 B.n115 B.n114 163.367
R510 B.n116 B.n115 163.367
R511 B.n116 B.n103 163.367
R512 B.n120 B.n103 163.367
R513 B.n121 B.n120 163.367
R514 B.n122 B.n121 163.367
R515 B.n122 B.n101 163.367
R516 B.n126 B.n101 163.367
R517 B.n127 B.n126 163.367
R518 B.n128 B.n127 163.367
R519 B.n128 B.n99 163.367
R520 B.n132 B.n99 163.367
R521 B.n133 B.n132 163.367
R522 B.n134 B.n133 163.367
R523 B.n134 B.n97 163.367
R524 B.n138 B.n97 163.367
R525 B.n139 B.n138 163.367
R526 B.n140 B.n139 163.367
R527 B.n140 B.n95 163.367
R528 B.n144 B.n95 163.367
R529 B.n145 B.n144 163.367
R530 B.n146 B.n145 163.367
R531 B.n146 B.n93 163.367
R532 B.n150 B.n93 163.367
R533 B.n151 B.n150 163.367
R534 B.n152 B.n151 163.367
R535 B.n172 B.n85 59.5399
R536 B.n188 B.n187 59.5399
R537 B.n326 B.n33 59.5399
R538 B.n26 B.n25 59.5399
R539 B.n361 B.n18 33.2493
R540 B.n308 B.n307 33.2493
R541 B.n207 B.n72 33.2493
R542 B.n154 B.n153 33.2493
R543 B.n85 B.n84 26.7641
R544 B.n187 B.n186 26.7641
R545 B.n33 B.n32 26.7641
R546 B.n25 B.n24 26.7641
R547 B B.n409 18.0485
R548 B.n362 B.n361 10.6151
R549 B.n363 B.n362 10.6151
R550 B.n363 B.n16 10.6151
R551 B.n367 B.n16 10.6151
R552 B.n368 B.n367 10.6151
R553 B.n369 B.n368 10.6151
R554 B.n369 B.n14 10.6151
R555 B.n373 B.n14 10.6151
R556 B.n374 B.n373 10.6151
R557 B.n375 B.n374 10.6151
R558 B.n375 B.n12 10.6151
R559 B.n379 B.n12 10.6151
R560 B.n380 B.n379 10.6151
R561 B.n381 B.n380 10.6151
R562 B.n381 B.n10 10.6151
R563 B.n385 B.n10 10.6151
R564 B.n386 B.n385 10.6151
R565 B.n387 B.n386 10.6151
R566 B.n387 B.n8 10.6151
R567 B.n391 B.n8 10.6151
R568 B.n392 B.n391 10.6151
R569 B.n393 B.n392 10.6151
R570 B.n393 B.n6 10.6151
R571 B.n397 B.n6 10.6151
R572 B.n398 B.n397 10.6151
R573 B.n399 B.n398 10.6151
R574 B.n399 B.n4 10.6151
R575 B.n403 B.n4 10.6151
R576 B.n404 B.n403 10.6151
R577 B.n405 B.n404 10.6151
R578 B.n405 B.n0 10.6151
R579 B.n357 B.n18 10.6151
R580 B.n357 B.n356 10.6151
R581 B.n356 B.n355 10.6151
R582 B.n355 B.n20 10.6151
R583 B.n351 B.n20 10.6151
R584 B.n351 B.n350 10.6151
R585 B.n350 B.n349 10.6151
R586 B.n349 B.n22 10.6151
R587 B.n345 B.n22 10.6151
R588 B.n345 B.n344 10.6151
R589 B.n344 B.n343 10.6151
R590 B.n340 B.n339 10.6151
R591 B.n339 B.n338 10.6151
R592 B.n338 B.n28 10.6151
R593 B.n334 B.n28 10.6151
R594 B.n334 B.n333 10.6151
R595 B.n333 B.n332 10.6151
R596 B.n332 B.n30 10.6151
R597 B.n328 B.n30 10.6151
R598 B.n328 B.n327 10.6151
R599 B.n325 B.n34 10.6151
R600 B.n321 B.n34 10.6151
R601 B.n321 B.n320 10.6151
R602 B.n320 B.n319 10.6151
R603 B.n319 B.n36 10.6151
R604 B.n315 B.n36 10.6151
R605 B.n315 B.n314 10.6151
R606 B.n314 B.n313 10.6151
R607 B.n313 B.n38 10.6151
R608 B.n309 B.n38 10.6151
R609 B.n309 B.n308 10.6151
R610 B.n307 B.n40 10.6151
R611 B.n303 B.n40 10.6151
R612 B.n303 B.n302 10.6151
R613 B.n302 B.n301 10.6151
R614 B.n301 B.n42 10.6151
R615 B.n297 B.n42 10.6151
R616 B.n297 B.n296 10.6151
R617 B.n296 B.n295 10.6151
R618 B.n295 B.n44 10.6151
R619 B.n291 B.n44 10.6151
R620 B.n291 B.n290 10.6151
R621 B.n290 B.n289 10.6151
R622 B.n289 B.n46 10.6151
R623 B.n285 B.n46 10.6151
R624 B.n285 B.n284 10.6151
R625 B.n284 B.n283 10.6151
R626 B.n283 B.n48 10.6151
R627 B.n279 B.n48 10.6151
R628 B.n279 B.n278 10.6151
R629 B.n278 B.n277 10.6151
R630 B.n277 B.n50 10.6151
R631 B.n273 B.n50 10.6151
R632 B.n273 B.n272 10.6151
R633 B.n272 B.n271 10.6151
R634 B.n271 B.n52 10.6151
R635 B.n267 B.n52 10.6151
R636 B.n267 B.n266 10.6151
R637 B.n266 B.n265 10.6151
R638 B.n265 B.n54 10.6151
R639 B.n261 B.n54 10.6151
R640 B.n261 B.n260 10.6151
R641 B.n260 B.n259 10.6151
R642 B.n259 B.n56 10.6151
R643 B.n255 B.n56 10.6151
R644 B.n255 B.n254 10.6151
R645 B.n254 B.n253 10.6151
R646 B.n253 B.n58 10.6151
R647 B.n249 B.n58 10.6151
R648 B.n249 B.n248 10.6151
R649 B.n248 B.n247 10.6151
R650 B.n247 B.n60 10.6151
R651 B.n243 B.n60 10.6151
R652 B.n243 B.n242 10.6151
R653 B.n242 B.n241 10.6151
R654 B.n241 B.n62 10.6151
R655 B.n237 B.n62 10.6151
R656 B.n237 B.n236 10.6151
R657 B.n236 B.n235 10.6151
R658 B.n235 B.n64 10.6151
R659 B.n231 B.n64 10.6151
R660 B.n231 B.n230 10.6151
R661 B.n230 B.n229 10.6151
R662 B.n229 B.n66 10.6151
R663 B.n225 B.n66 10.6151
R664 B.n225 B.n224 10.6151
R665 B.n224 B.n223 10.6151
R666 B.n223 B.n68 10.6151
R667 B.n219 B.n68 10.6151
R668 B.n219 B.n218 10.6151
R669 B.n218 B.n217 10.6151
R670 B.n217 B.n70 10.6151
R671 B.n213 B.n70 10.6151
R672 B.n213 B.n212 10.6151
R673 B.n212 B.n211 10.6151
R674 B.n211 B.n72 10.6151
R675 B.n107 B.n1 10.6151
R676 B.n107 B.n106 10.6151
R677 B.n111 B.n106 10.6151
R678 B.n112 B.n111 10.6151
R679 B.n113 B.n112 10.6151
R680 B.n113 B.n104 10.6151
R681 B.n117 B.n104 10.6151
R682 B.n118 B.n117 10.6151
R683 B.n119 B.n118 10.6151
R684 B.n119 B.n102 10.6151
R685 B.n123 B.n102 10.6151
R686 B.n124 B.n123 10.6151
R687 B.n125 B.n124 10.6151
R688 B.n125 B.n100 10.6151
R689 B.n129 B.n100 10.6151
R690 B.n130 B.n129 10.6151
R691 B.n131 B.n130 10.6151
R692 B.n131 B.n98 10.6151
R693 B.n135 B.n98 10.6151
R694 B.n136 B.n135 10.6151
R695 B.n137 B.n136 10.6151
R696 B.n137 B.n96 10.6151
R697 B.n141 B.n96 10.6151
R698 B.n142 B.n141 10.6151
R699 B.n143 B.n142 10.6151
R700 B.n143 B.n94 10.6151
R701 B.n147 B.n94 10.6151
R702 B.n148 B.n147 10.6151
R703 B.n149 B.n148 10.6151
R704 B.n149 B.n92 10.6151
R705 B.n153 B.n92 10.6151
R706 B.n155 B.n154 10.6151
R707 B.n155 B.n90 10.6151
R708 B.n159 B.n90 10.6151
R709 B.n160 B.n159 10.6151
R710 B.n161 B.n160 10.6151
R711 B.n161 B.n88 10.6151
R712 B.n165 B.n88 10.6151
R713 B.n166 B.n165 10.6151
R714 B.n167 B.n166 10.6151
R715 B.n167 B.n86 10.6151
R716 B.n171 B.n86 10.6151
R717 B.n174 B.n173 10.6151
R718 B.n174 B.n82 10.6151
R719 B.n178 B.n82 10.6151
R720 B.n179 B.n178 10.6151
R721 B.n180 B.n179 10.6151
R722 B.n180 B.n80 10.6151
R723 B.n184 B.n80 10.6151
R724 B.n185 B.n184 10.6151
R725 B.n189 B.n185 10.6151
R726 B.n193 B.n78 10.6151
R727 B.n194 B.n193 10.6151
R728 B.n195 B.n194 10.6151
R729 B.n195 B.n76 10.6151
R730 B.n199 B.n76 10.6151
R731 B.n200 B.n199 10.6151
R732 B.n201 B.n200 10.6151
R733 B.n201 B.n74 10.6151
R734 B.n205 B.n74 10.6151
R735 B.n206 B.n205 10.6151
R736 B.n207 B.n206 10.6151
R737 B.n343 B.n26 9.36635
R738 B.n326 B.n325 9.36635
R739 B.n172 B.n171 9.36635
R740 B.n188 B.n78 9.36635
R741 B.n409 B.n0 8.11757
R742 B.n409 B.n1 8.11757
R743 B.n340 B.n26 1.24928
R744 B.n327 B.n326 1.24928
R745 B.n173 B.n172 1.24928
R746 B.n189 B.n188 1.24928
R747 VP.n10 VP.n7 161.3
R748 VP.n12 VP.n11 161.3
R749 VP.n13 VP.n6 161.3
R750 VP.n16 VP.n15 161.3
R751 VP.n17 VP.n5 161.3
R752 VP.n19 VP.n18 161.3
R753 VP.n21 VP.n4 161.3
R754 VP.n40 VP.n0 161.3
R755 VP.n38 VP.n37 161.3
R756 VP.n36 VP.n1 161.3
R757 VP.n35 VP.n34 161.3
R758 VP.n32 VP.n2 161.3
R759 VP.n31 VP.n30 161.3
R760 VP.n29 VP.n3 161.3
R761 VP.n28 VP.n27 161.3
R762 VP.n9 VP.t5 99.3881
R763 VP.n25 VP.t7 84.2357
R764 VP.n41 VP.t6 84.2357
R765 VP.n22 VP.t8 84.2357
R766 VP.n23 VP.n22 80.6037
R767 VP.n42 VP.n41 80.6037
R768 VP.n25 VP.n24 80.6037
R769 VP.n27 VP.n25 55.824
R770 VP.n41 VP.n40 55.824
R771 VP.n22 VP.n21 55.824
R772 VP.n9 VP.n8 48.4137
R773 VP.n26 VP.t1 46.8234
R774 VP.n33 VP.t2 46.8234
R775 VP.n39 VP.t0 46.8234
R776 VP.n20 VP.t9 46.8234
R777 VP.n14 VP.t3 46.8234
R778 VP.n8 VP.t4 46.8234
R779 VP.n32 VP.n31 46.3896
R780 VP.n34 VP.n1 46.3896
R781 VP.n15 VP.n5 46.3896
R782 VP.n13 VP.n12 46.3896
R783 VP.n10 VP.n9 43.9713
R784 VP.n24 VP.n23 37.3802
R785 VP.n31 VP.n3 34.7644
R786 VP.n38 VP.n1 34.7644
R787 VP.n19 VP.n5 34.7644
R788 VP.n12 VP.n7 34.7644
R789 VP.n27 VP.n26 18.1985
R790 VP.n40 VP.n39 18.1985
R791 VP.n21 VP.n20 18.1985
R792 VP.n33 VP.n32 12.2964
R793 VP.n34 VP.n33 12.2964
R794 VP.n14 VP.n13 12.2964
R795 VP.n15 VP.n14 12.2964
R796 VP.n26 VP.n3 6.39438
R797 VP.n39 VP.n38 6.39438
R798 VP.n20 VP.n19 6.39438
R799 VP.n8 VP.n7 6.39438
R800 VP.n23 VP.n4 0.285035
R801 VP.n28 VP.n24 0.285035
R802 VP.n42 VP.n0 0.285035
R803 VP.n11 VP.n10 0.189894
R804 VP.n11 VP.n6 0.189894
R805 VP.n16 VP.n6 0.189894
R806 VP.n17 VP.n16 0.189894
R807 VP.n18 VP.n17 0.189894
R808 VP.n18 VP.n4 0.189894
R809 VP.n29 VP.n28 0.189894
R810 VP.n30 VP.n29 0.189894
R811 VP.n30 VP.n2 0.189894
R812 VP.n35 VP.n2 0.189894
R813 VP.n36 VP.n35 0.189894
R814 VP.n37 VP.n36 0.189894
R815 VP.n37 VP.n0 0.189894
R816 VP VP.n42 0.146778
R817 VDD1.n3 VDD1.t2 187.963
R818 VDD1.n1 VDD1.t4 187.963
R819 VDD1.n5 VDD1.n4 171.677
R820 VDD1.n1 VDD1.n0 170.839
R821 VDD1.n7 VDD1.n6 170.839
R822 VDD1.n3 VDD1.n2 170.839
R823 VDD1.n7 VDD1.n5 32.3026
R824 VDD1.n6 VDD1.t0 15.9343
R825 VDD1.n6 VDD1.t1 15.9343
R826 VDD1.n0 VDD1.t5 15.9343
R827 VDD1.n0 VDD1.t6 15.9343
R828 VDD1.n4 VDD1.t9 15.9343
R829 VDD1.n4 VDD1.t3 15.9343
R830 VDD1.n2 VDD1.t8 15.9343
R831 VDD1.n2 VDD1.t7 15.9343
R832 VDD1 VDD1.n7 0.834552
R833 VDD1 VDD1.n1 0.356103
R834 VDD1.n5 VDD1.n3 0.242568
C0 w_n2626_n1376# VDD2 1.52144f
C1 w_n2626_n1376# B 5.15214f
C2 w_n2626_n1376# VTAIL 1.485f
C3 VDD2 B 1.16811f
C4 VTAIL VDD2 4.536f
C5 VTAIL B 1.01623f
C6 VDD1 w_n2626_n1376# 1.45916f
C7 VDD1 VDD2 1.19029f
C8 w_n2626_n1376# VP 5.26071f
C9 w_n2626_n1376# VN 4.92805f
C10 VDD1 B 1.11019f
C11 VDD1 VTAIL 4.49368f
C12 VDD2 VP 0.392289f
C13 VDD2 VN 1.75988f
C14 B VP 1.32882f
C15 VN B 0.771237f
C16 VTAIL VP 2.32259f
C17 VTAIL VN 2.30842f
C18 VDD1 VP 1.9933f
C19 VDD1 VN 0.156472f
C20 VN VP 4.26923f
C21 VDD2 VSUBS 0.82398f
C22 VDD1 VSUBS 0.942118f
C23 VTAIL VSUBS 0.380931f
C24 VN VSUBS 4.72081f
C25 VP VSUBS 1.766486f
C26 B VSUBS 2.464391f
C27 w_n2626_n1376# VSUBS 46.102104f
C28 VDD1.t4 VSUBS 0.184017f
C29 VDD1.t5 VSUBS 0.027104f
C30 VDD1.t6 VSUBS 0.027104f
C31 VDD1.n0 VSUBS 0.122909f
C32 VDD1.n1 VSUBS 0.523292f
C33 VDD1.t2 VSUBS 0.184017f
C34 VDD1.t8 VSUBS 0.027104f
C35 VDD1.t7 VSUBS 0.027104f
C36 VDD1.n2 VSUBS 0.122909f
C37 VDD1.n3 VSUBS 0.518752f
C38 VDD1.t9 VSUBS 0.027104f
C39 VDD1.t3 VSUBS 0.027104f
C40 VDD1.n4 VSUBS 0.124346f
C41 VDD1.n5 VSUBS 1.10669f
C42 VDD1.t0 VSUBS 0.027104f
C43 VDD1.t1 VSUBS 0.027104f
C44 VDD1.n6 VSUBS 0.122908f
C45 VDD1.n7 VSUBS 1.20888f
C46 VP.n0 VSUBS 0.07824f
C47 VP.t0 VSUBS 0.294464f
C48 VP.n1 VSUBS 0.050104f
C49 VP.n2 VSUBS 0.058635f
C50 VP.t2 VSUBS 0.294464f
C51 VP.n3 VSUBS 0.07812f
C52 VP.n4 VSUBS 0.07824f
C53 VP.t8 VSUBS 0.388209f
C54 VP.t9 VSUBS 0.294464f
C55 VP.n5 VSUBS 0.050104f
C56 VP.n6 VSUBS 0.058635f
C57 VP.t3 VSUBS 0.294464f
C58 VP.n7 VSUBS 0.07812f
C59 VP.t4 VSUBS 0.294464f
C60 VP.n8 VSUBS 0.222434f
C61 VP.t5 VSUBS 0.429072f
C62 VP.n9 VSUBS 0.258985f
C63 VP.n10 VSUBS 0.253884f
C64 VP.n11 VSUBS 0.058635f
C65 VP.n12 VSUBS 0.050104f
C66 VP.n13 VSUBS 0.084415f
C67 VP.n14 VSUBS 0.171004f
C68 VP.n15 VSUBS 0.084415f
C69 VP.n16 VSUBS 0.058635f
C70 VP.n17 VSUBS 0.058635f
C71 VP.n18 VSUBS 0.058635f
C72 VP.n19 VSUBS 0.07812f
C73 VP.n20 VSUBS 0.171004f
C74 VP.n21 VSUBS 0.082406f
C75 VP.n22 VSUBS 0.267612f
C76 VP.n23 VSUBS 1.99703f
C77 VP.n24 VSUBS 2.05358f
C78 VP.t7 VSUBS 0.388209f
C79 VP.n25 VSUBS 0.267612f
C80 VP.t1 VSUBS 0.294464f
C81 VP.n26 VSUBS 0.171004f
C82 VP.n27 VSUBS 0.082406f
C83 VP.n28 VSUBS 0.07824f
C84 VP.n29 VSUBS 0.058635f
C85 VP.n30 VSUBS 0.058635f
C86 VP.n31 VSUBS 0.050104f
C87 VP.n32 VSUBS 0.084415f
C88 VP.n33 VSUBS 0.171004f
C89 VP.n34 VSUBS 0.084415f
C90 VP.n35 VSUBS 0.058635f
C91 VP.n36 VSUBS 0.058635f
C92 VP.n37 VSUBS 0.058635f
C93 VP.n38 VSUBS 0.07812f
C94 VP.n39 VSUBS 0.171004f
C95 VP.n40 VSUBS 0.082406f
C96 VP.t6 VSUBS 0.388209f
C97 VP.n41 VSUBS 0.267612f
C98 VP.n42 VSUBS 0.054914f
C99 B.n0 VSUBS 0.007566f
C100 B.n1 VSUBS 0.007566f
C101 B.n2 VSUBS 0.011189f
C102 B.n3 VSUBS 0.008574f
C103 B.n4 VSUBS 0.008574f
C104 B.n5 VSUBS 0.008574f
C105 B.n6 VSUBS 0.008574f
C106 B.n7 VSUBS 0.008574f
C107 B.n8 VSUBS 0.008574f
C108 B.n9 VSUBS 0.008574f
C109 B.n10 VSUBS 0.008574f
C110 B.n11 VSUBS 0.008574f
C111 B.n12 VSUBS 0.008574f
C112 B.n13 VSUBS 0.008574f
C113 B.n14 VSUBS 0.008574f
C114 B.n15 VSUBS 0.008574f
C115 B.n16 VSUBS 0.008574f
C116 B.n17 VSUBS 0.008574f
C117 B.n18 VSUBS 0.020653f
C118 B.n19 VSUBS 0.008574f
C119 B.n20 VSUBS 0.008574f
C120 B.n21 VSUBS 0.008574f
C121 B.n22 VSUBS 0.008574f
C122 B.n23 VSUBS 0.008574f
C123 B.t1 VSUBS 0.054312f
C124 B.t2 VSUBS 0.061279f
C125 B.t0 VSUBS 0.126469f
C126 B.n24 VSUBS 0.07048f
C127 B.n25 VSUBS 0.063689f
C128 B.n26 VSUBS 0.019866f
C129 B.n27 VSUBS 0.008574f
C130 B.n28 VSUBS 0.008574f
C131 B.n29 VSUBS 0.008574f
C132 B.n30 VSUBS 0.008574f
C133 B.n31 VSUBS 0.008574f
C134 B.t10 VSUBS 0.054312f
C135 B.t11 VSUBS 0.061279f
C136 B.t9 VSUBS 0.126469f
C137 B.n32 VSUBS 0.07048f
C138 B.n33 VSUBS 0.06369f
C139 B.n34 VSUBS 0.008574f
C140 B.n35 VSUBS 0.008574f
C141 B.n36 VSUBS 0.008574f
C142 B.n37 VSUBS 0.008574f
C143 B.n38 VSUBS 0.008574f
C144 B.n39 VSUBS 0.020653f
C145 B.n40 VSUBS 0.008574f
C146 B.n41 VSUBS 0.008574f
C147 B.n42 VSUBS 0.008574f
C148 B.n43 VSUBS 0.008574f
C149 B.n44 VSUBS 0.008574f
C150 B.n45 VSUBS 0.008574f
C151 B.n46 VSUBS 0.008574f
C152 B.n47 VSUBS 0.008574f
C153 B.n48 VSUBS 0.008574f
C154 B.n49 VSUBS 0.008574f
C155 B.n50 VSUBS 0.008574f
C156 B.n51 VSUBS 0.008574f
C157 B.n52 VSUBS 0.008574f
C158 B.n53 VSUBS 0.008574f
C159 B.n54 VSUBS 0.008574f
C160 B.n55 VSUBS 0.008574f
C161 B.n56 VSUBS 0.008574f
C162 B.n57 VSUBS 0.008574f
C163 B.n58 VSUBS 0.008574f
C164 B.n59 VSUBS 0.008574f
C165 B.n60 VSUBS 0.008574f
C166 B.n61 VSUBS 0.008574f
C167 B.n62 VSUBS 0.008574f
C168 B.n63 VSUBS 0.008574f
C169 B.n64 VSUBS 0.008574f
C170 B.n65 VSUBS 0.008574f
C171 B.n66 VSUBS 0.008574f
C172 B.n67 VSUBS 0.008574f
C173 B.n68 VSUBS 0.008574f
C174 B.n69 VSUBS 0.008574f
C175 B.n70 VSUBS 0.008574f
C176 B.n71 VSUBS 0.008574f
C177 B.n72 VSUBS 0.020944f
C178 B.n73 VSUBS 0.008574f
C179 B.n74 VSUBS 0.008574f
C180 B.n75 VSUBS 0.008574f
C181 B.n76 VSUBS 0.008574f
C182 B.n77 VSUBS 0.008574f
C183 B.n78 VSUBS 0.00807f
C184 B.n79 VSUBS 0.008574f
C185 B.n80 VSUBS 0.008574f
C186 B.n81 VSUBS 0.008574f
C187 B.n82 VSUBS 0.008574f
C188 B.n83 VSUBS 0.008574f
C189 B.t8 VSUBS 0.054312f
C190 B.t7 VSUBS 0.061279f
C191 B.t6 VSUBS 0.126469f
C192 B.n84 VSUBS 0.07048f
C193 B.n85 VSUBS 0.063689f
C194 B.n86 VSUBS 0.008574f
C195 B.n87 VSUBS 0.008574f
C196 B.n88 VSUBS 0.008574f
C197 B.n89 VSUBS 0.008574f
C198 B.n90 VSUBS 0.008574f
C199 B.n91 VSUBS 0.020653f
C200 B.n92 VSUBS 0.008574f
C201 B.n93 VSUBS 0.008574f
C202 B.n94 VSUBS 0.008574f
C203 B.n95 VSUBS 0.008574f
C204 B.n96 VSUBS 0.008574f
C205 B.n97 VSUBS 0.008574f
C206 B.n98 VSUBS 0.008574f
C207 B.n99 VSUBS 0.008574f
C208 B.n100 VSUBS 0.008574f
C209 B.n101 VSUBS 0.008574f
C210 B.n102 VSUBS 0.008574f
C211 B.n103 VSUBS 0.008574f
C212 B.n104 VSUBS 0.008574f
C213 B.n105 VSUBS 0.008574f
C214 B.n106 VSUBS 0.008574f
C215 B.n107 VSUBS 0.008574f
C216 B.n108 VSUBS 0.008574f
C217 B.n109 VSUBS 0.008574f
C218 B.n110 VSUBS 0.008574f
C219 B.n111 VSUBS 0.008574f
C220 B.n112 VSUBS 0.008574f
C221 B.n113 VSUBS 0.008574f
C222 B.n114 VSUBS 0.008574f
C223 B.n115 VSUBS 0.008574f
C224 B.n116 VSUBS 0.008574f
C225 B.n117 VSUBS 0.008574f
C226 B.n118 VSUBS 0.008574f
C227 B.n119 VSUBS 0.008574f
C228 B.n120 VSUBS 0.008574f
C229 B.n121 VSUBS 0.008574f
C230 B.n122 VSUBS 0.008574f
C231 B.n123 VSUBS 0.008574f
C232 B.n124 VSUBS 0.008574f
C233 B.n125 VSUBS 0.008574f
C234 B.n126 VSUBS 0.008574f
C235 B.n127 VSUBS 0.008574f
C236 B.n128 VSUBS 0.008574f
C237 B.n129 VSUBS 0.008574f
C238 B.n130 VSUBS 0.008574f
C239 B.n131 VSUBS 0.008574f
C240 B.n132 VSUBS 0.008574f
C241 B.n133 VSUBS 0.008574f
C242 B.n134 VSUBS 0.008574f
C243 B.n135 VSUBS 0.008574f
C244 B.n136 VSUBS 0.008574f
C245 B.n137 VSUBS 0.008574f
C246 B.n138 VSUBS 0.008574f
C247 B.n139 VSUBS 0.008574f
C248 B.n140 VSUBS 0.008574f
C249 B.n141 VSUBS 0.008574f
C250 B.n142 VSUBS 0.008574f
C251 B.n143 VSUBS 0.008574f
C252 B.n144 VSUBS 0.008574f
C253 B.n145 VSUBS 0.008574f
C254 B.n146 VSUBS 0.008574f
C255 B.n147 VSUBS 0.008574f
C256 B.n148 VSUBS 0.008574f
C257 B.n149 VSUBS 0.008574f
C258 B.n150 VSUBS 0.008574f
C259 B.n151 VSUBS 0.008574f
C260 B.n152 VSUBS 0.019949f
C261 B.n153 VSUBS 0.019949f
C262 B.n154 VSUBS 0.020653f
C263 B.n155 VSUBS 0.008574f
C264 B.n156 VSUBS 0.008574f
C265 B.n157 VSUBS 0.008574f
C266 B.n158 VSUBS 0.008574f
C267 B.n159 VSUBS 0.008574f
C268 B.n160 VSUBS 0.008574f
C269 B.n161 VSUBS 0.008574f
C270 B.n162 VSUBS 0.008574f
C271 B.n163 VSUBS 0.008574f
C272 B.n164 VSUBS 0.008574f
C273 B.n165 VSUBS 0.008574f
C274 B.n166 VSUBS 0.008574f
C275 B.n167 VSUBS 0.008574f
C276 B.n168 VSUBS 0.008574f
C277 B.n169 VSUBS 0.008574f
C278 B.n170 VSUBS 0.008574f
C279 B.n171 VSUBS 0.00807f
C280 B.n172 VSUBS 0.019866f
C281 B.n173 VSUBS 0.004792f
C282 B.n174 VSUBS 0.008574f
C283 B.n175 VSUBS 0.008574f
C284 B.n176 VSUBS 0.008574f
C285 B.n177 VSUBS 0.008574f
C286 B.n178 VSUBS 0.008574f
C287 B.n179 VSUBS 0.008574f
C288 B.n180 VSUBS 0.008574f
C289 B.n181 VSUBS 0.008574f
C290 B.n182 VSUBS 0.008574f
C291 B.n183 VSUBS 0.008574f
C292 B.n184 VSUBS 0.008574f
C293 B.n185 VSUBS 0.008574f
C294 B.t5 VSUBS 0.054312f
C295 B.t4 VSUBS 0.061279f
C296 B.t3 VSUBS 0.126469f
C297 B.n186 VSUBS 0.07048f
C298 B.n187 VSUBS 0.06369f
C299 B.n188 VSUBS 0.019866f
C300 B.n189 VSUBS 0.004792f
C301 B.n190 VSUBS 0.008574f
C302 B.n191 VSUBS 0.008574f
C303 B.n192 VSUBS 0.008574f
C304 B.n193 VSUBS 0.008574f
C305 B.n194 VSUBS 0.008574f
C306 B.n195 VSUBS 0.008574f
C307 B.n196 VSUBS 0.008574f
C308 B.n197 VSUBS 0.008574f
C309 B.n198 VSUBS 0.008574f
C310 B.n199 VSUBS 0.008574f
C311 B.n200 VSUBS 0.008574f
C312 B.n201 VSUBS 0.008574f
C313 B.n202 VSUBS 0.008574f
C314 B.n203 VSUBS 0.008574f
C315 B.n204 VSUBS 0.008574f
C316 B.n205 VSUBS 0.008574f
C317 B.n206 VSUBS 0.008574f
C318 B.n207 VSUBS 0.019658f
C319 B.n208 VSUBS 0.020653f
C320 B.n209 VSUBS 0.019949f
C321 B.n210 VSUBS 0.008574f
C322 B.n211 VSUBS 0.008574f
C323 B.n212 VSUBS 0.008574f
C324 B.n213 VSUBS 0.008574f
C325 B.n214 VSUBS 0.008574f
C326 B.n215 VSUBS 0.008574f
C327 B.n216 VSUBS 0.008574f
C328 B.n217 VSUBS 0.008574f
C329 B.n218 VSUBS 0.008574f
C330 B.n219 VSUBS 0.008574f
C331 B.n220 VSUBS 0.008574f
C332 B.n221 VSUBS 0.008574f
C333 B.n222 VSUBS 0.008574f
C334 B.n223 VSUBS 0.008574f
C335 B.n224 VSUBS 0.008574f
C336 B.n225 VSUBS 0.008574f
C337 B.n226 VSUBS 0.008574f
C338 B.n227 VSUBS 0.008574f
C339 B.n228 VSUBS 0.008574f
C340 B.n229 VSUBS 0.008574f
C341 B.n230 VSUBS 0.008574f
C342 B.n231 VSUBS 0.008574f
C343 B.n232 VSUBS 0.008574f
C344 B.n233 VSUBS 0.008574f
C345 B.n234 VSUBS 0.008574f
C346 B.n235 VSUBS 0.008574f
C347 B.n236 VSUBS 0.008574f
C348 B.n237 VSUBS 0.008574f
C349 B.n238 VSUBS 0.008574f
C350 B.n239 VSUBS 0.008574f
C351 B.n240 VSUBS 0.008574f
C352 B.n241 VSUBS 0.008574f
C353 B.n242 VSUBS 0.008574f
C354 B.n243 VSUBS 0.008574f
C355 B.n244 VSUBS 0.008574f
C356 B.n245 VSUBS 0.008574f
C357 B.n246 VSUBS 0.008574f
C358 B.n247 VSUBS 0.008574f
C359 B.n248 VSUBS 0.008574f
C360 B.n249 VSUBS 0.008574f
C361 B.n250 VSUBS 0.008574f
C362 B.n251 VSUBS 0.008574f
C363 B.n252 VSUBS 0.008574f
C364 B.n253 VSUBS 0.008574f
C365 B.n254 VSUBS 0.008574f
C366 B.n255 VSUBS 0.008574f
C367 B.n256 VSUBS 0.008574f
C368 B.n257 VSUBS 0.008574f
C369 B.n258 VSUBS 0.008574f
C370 B.n259 VSUBS 0.008574f
C371 B.n260 VSUBS 0.008574f
C372 B.n261 VSUBS 0.008574f
C373 B.n262 VSUBS 0.008574f
C374 B.n263 VSUBS 0.008574f
C375 B.n264 VSUBS 0.008574f
C376 B.n265 VSUBS 0.008574f
C377 B.n266 VSUBS 0.008574f
C378 B.n267 VSUBS 0.008574f
C379 B.n268 VSUBS 0.008574f
C380 B.n269 VSUBS 0.008574f
C381 B.n270 VSUBS 0.008574f
C382 B.n271 VSUBS 0.008574f
C383 B.n272 VSUBS 0.008574f
C384 B.n273 VSUBS 0.008574f
C385 B.n274 VSUBS 0.008574f
C386 B.n275 VSUBS 0.008574f
C387 B.n276 VSUBS 0.008574f
C388 B.n277 VSUBS 0.008574f
C389 B.n278 VSUBS 0.008574f
C390 B.n279 VSUBS 0.008574f
C391 B.n280 VSUBS 0.008574f
C392 B.n281 VSUBS 0.008574f
C393 B.n282 VSUBS 0.008574f
C394 B.n283 VSUBS 0.008574f
C395 B.n284 VSUBS 0.008574f
C396 B.n285 VSUBS 0.008574f
C397 B.n286 VSUBS 0.008574f
C398 B.n287 VSUBS 0.008574f
C399 B.n288 VSUBS 0.008574f
C400 B.n289 VSUBS 0.008574f
C401 B.n290 VSUBS 0.008574f
C402 B.n291 VSUBS 0.008574f
C403 B.n292 VSUBS 0.008574f
C404 B.n293 VSUBS 0.008574f
C405 B.n294 VSUBS 0.008574f
C406 B.n295 VSUBS 0.008574f
C407 B.n296 VSUBS 0.008574f
C408 B.n297 VSUBS 0.008574f
C409 B.n298 VSUBS 0.008574f
C410 B.n299 VSUBS 0.008574f
C411 B.n300 VSUBS 0.008574f
C412 B.n301 VSUBS 0.008574f
C413 B.n302 VSUBS 0.008574f
C414 B.n303 VSUBS 0.008574f
C415 B.n304 VSUBS 0.008574f
C416 B.n305 VSUBS 0.008574f
C417 B.n306 VSUBS 0.019949f
C418 B.n307 VSUBS 0.019949f
C419 B.n308 VSUBS 0.020653f
C420 B.n309 VSUBS 0.008574f
C421 B.n310 VSUBS 0.008574f
C422 B.n311 VSUBS 0.008574f
C423 B.n312 VSUBS 0.008574f
C424 B.n313 VSUBS 0.008574f
C425 B.n314 VSUBS 0.008574f
C426 B.n315 VSUBS 0.008574f
C427 B.n316 VSUBS 0.008574f
C428 B.n317 VSUBS 0.008574f
C429 B.n318 VSUBS 0.008574f
C430 B.n319 VSUBS 0.008574f
C431 B.n320 VSUBS 0.008574f
C432 B.n321 VSUBS 0.008574f
C433 B.n322 VSUBS 0.008574f
C434 B.n323 VSUBS 0.008574f
C435 B.n324 VSUBS 0.008574f
C436 B.n325 VSUBS 0.00807f
C437 B.n326 VSUBS 0.019866f
C438 B.n327 VSUBS 0.004792f
C439 B.n328 VSUBS 0.008574f
C440 B.n329 VSUBS 0.008574f
C441 B.n330 VSUBS 0.008574f
C442 B.n331 VSUBS 0.008574f
C443 B.n332 VSUBS 0.008574f
C444 B.n333 VSUBS 0.008574f
C445 B.n334 VSUBS 0.008574f
C446 B.n335 VSUBS 0.008574f
C447 B.n336 VSUBS 0.008574f
C448 B.n337 VSUBS 0.008574f
C449 B.n338 VSUBS 0.008574f
C450 B.n339 VSUBS 0.008574f
C451 B.n340 VSUBS 0.004792f
C452 B.n341 VSUBS 0.008574f
C453 B.n342 VSUBS 0.008574f
C454 B.n343 VSUBS 0.00807f
C455 B.n344 VSUBS 0.008574f
C456 B.n345 VSUBS 0.008574f
C457 B.n346 VSUBS 0.008574f
C458 B.n347 VSUBS 0.008574f
C459 B.n348 VSUBS 0.008574f
C460 B.n349 VSUBS 0.008574f
C461 B.n350 VSUBS 0.008574f
C462 B.n351 VSUBS 0.008574f
C463 B.n352 VSUBS 0.008574f
C464 B.n353 VSUBS 0.008574f
C465 B.n354 VSUBS 0.008574f
C466 B.n355 VSUBS 0.008574f
C467 B.n356 VSUBS 0.008574f
C468 B.n357 VSUBS 0.008574f
C469 B.n358 VSUBS 0.008574f
C470 B.n359 VSUBS 0.020653f
C471 B.n360 VSUBS 0.019949f
C472 B.n361 VSUBS 0.019949f
C473 B.n362 VSUBS 0.008574f
C474 B.n363 VSUBS 0.008574f
C475 B.n364 VSUBS 0.008574f
C476 B.n365 VSUBS 0.008574f
C477 B.n366 VSUBS 0.008574f
C478 B.n367 VSUBS 0.008574f
C479 B.n368 VSUBS 0.008574f
C480 B.n369 VSUBS 0.008574f
C481 B.n370 VSUBS 0.008574f
C482 B.n371 VSUBS 0.008574f
C483 B.n372 VSUBS 0.008574f
C484 B.n373 VSUBS 0.008574f
C485 B.n374 VSUBS 0.008574f
C486 B.n375 VSUBS 0.008574f
C487 B.n376 VSUBS 0.008574f
C488 B.n377 VSUBS 0.008574f
C489 B.n378 VSUBS 0.008574f
C490 B.n379 VSUBS 0.008574f
C491 B.n380 VSUBS 0.008574f
C492 B.n381 VSUBS 0.008574f
C493 B.n382 VSUBS 0.008574f
C494 B.n383 VSUBS 0.008574f
C495 B.n384 VSUBS 0.008574f
C496 B.n385 VSUBS 0.008574f
C497 B.n386 VSUBS 0.008574f
C498 B.n387 VSUBS 0.008574f
C499 B.n388 VSUBS 0.008574f
C500 B.n389 VSUBS 0.008574f
C501 B.n390 VSUBS 0.008574f
C502 B.n391 VSUBS 0.008574f
C503 B.n392 VSUBS 0.008574f
C504 B.n393 VSUBS 0.008574f
C505 B.n394 VSUBS 0.008574f
C506 B.n395 VSUBS 0.008574f
C507 B.n396 VSUBS 0.008574f
C508 B.n397 VSUBS 0.008574f
C509 B.n398 VSUBS 0.008574f
C510 B.n399 VSUBS 0.008574f
C511 B.n400 VSUBS 0.008574f
C512 B.n401 VSUBS 0.008574f
C513 B.n402 VSUBS 0.008574f
C514 B.n403 VSUBS 0.008574f
C515 B.n404 VSUBS 0.008574f
C516 B.n405 VSUBS 0.008574f
C517 B.n406 VSUBS 0.008574f
C518 B.n407 VSUBS 0.011189f
C519 B.n408 VSUBS 0.011919f
C520 B.n409 VSUBS 0.023703f
C521 VDD2.t2 VSUBS 0.186592f
C522 VDD2.t3 VSUBS 0.027483f
C523 VDD2.t5 VSUBS 0.027483f
C524 VDD2.n0 VSUBS 0.124628f
C525 VDD2.n1 VSUBS 0.526011f
C526 VDD2.t7 VSUBS 0.027483f
C527 VDD2.t8 VSUBS 0.027483f
C528 VDD2.n2 VSUBS 0.126086f
C529 VDD2.n3 VSUBS 1.06807f
C530 VDD2.t0 VSUBS 0.184901f
C531 VDD2.n4 VSUBS 1.18579f
C532 VDD2.t1 VSUBS 0.027483f
C533 VDD2.t9 VSUBS 0.027483f
C534 VDD2.n5 VSUBS 0.124629f
C535 VDD2.n6 VSUBS 0.265146f
C536 VDD2.t6 VSUBS 0.027483f
C537 VDD2.t4 VSUBS 0.027483f
C538 VDD2.n7 VSUBS 0.126078f
C539 VTAIL.t13 VSUBS 0.05261f
C540 VTAIL.t15 VSUBS 0.05261f
C541 VTAIL.n0 VSUBS 0.20191f
C542 VTAIL.n1 VSUBS 0.549266f
C543 VTAIL.t5 VSUBS 0.317965f
C544 VTAIL.n2 VSUBS 0.60185f
C545 VTAIL.t8 VSUBS 0.05261f
C546 VTAIL.t6 VSUBS 0.05261f
C547 VTAIL.n3 VSUBS 0.20191f
C548 VTAIL.n4 VSUBS 0.587567f
C549 VTAIL.t9 VSUBS 0.05261f
C550 VTAIL.t1 VSUBS 0.05261f
C551 VTAIL.n5 VSUBS 0.20191f
C552 VTAIL.n6 VSUBS 1.34091f
C553 VTAIL.t12 VSUBS 0.05261f
C554 VTAIL.t18 VSUBS 0.05261f
C555 VTAIL.n7 VSUBS 0.201911f
C556 VTAIL.n8 VSUBS 1.34091f
C557 VTAIL.t16 VSUBS 0.05261f
C558 VTAIL.t10 VSUBS 0.05261f
C559 VTAIL.n9 VSUBS 0.201911f
C560 VTAIL.n10 VSUBS 0.587566f
C561 VTAIL.t17 VSUBS 0.317966f
C562 VTAIL.n11 VSUBS 0.601848f
C563 VTAIL.t3 VSUBS 0.05261f
C564 VTAIL.t0 VSUBS 0.05261f
C565 VTAIL.n12 VSUBS 0.201911f
C566 VTAIL.n13 VSUBS 0.574422f
C567 VTAIL.t7 VSUBS 0.05261f
C568 VTAIL.t4 VSUBS 0.05261f
C569 VTAIL.n14 VSUBS 0.201911f
C570 VTAIL.n15 VSUBS 0.587566f
C571 VTAIL.t2 VSUBS 0.317965f
C572 VTAIL.n16 VSUBS 1.24323f
C573 VTAIL.t14 VSUBS 0.317965f
C574 VTAIL.n17 VSUBS 1.24323f
C575 VTAIL.t11 VSUBS 0.05261f
C576 VTAIL.t19 VSUBS 0.05261f
C577 VTAIL.n18 VSUBS 0.20191f
C578 VTAIL.n19 VSUBS 0.487622f
C579 VN.n0 VSUBS 0.07509f
C580 VN.t2 VSUBS 0.282609f
C581 VN.n1 VSUBS 0.048087f
C582 VN.n2 VSUBS 0.056274f
C583 VN.t4 VSUBS 0.282609f
C584 VN.n3 VSUBS 0.074975f
C585 VN.t7 VSUBS 0.411797f
C586 VN.t6 VSUBS 0.282609f
C587 VN.n4 VSUBS 0.213479f
C588 VN.n5 VSUBS 0.248558f
C589 VN.n6 VSUBS 0.243662f
C590 VN.n7 VSUBS 0.056274f
C591 VN.n8 VSUBS 0.048087f
C592 VN.n9 VSUBS 0.081017f
C593 VN.n10 VSUBS 0.164119f
C594 VN.n11 VSUBS 0.081017f
C595 VN.n12 VSUBS 0.056274f
C596 VN.n13 VSUBS 0.056274f
C597 VN.n14 VSUBS 0.056274f
C598 VN.n15 VSUBS 0.074975f
C599 VN.n16 VSUBS 0.164119f
C600 VN.n17 VSUBS 0.079089f
C601 VN.t1 VSUBS 0.37258f
C602 VN.n18 VSUBS 0.256837f
C603 VN.n19 VSUBS 0.052703f
C604 VN.n20 VSUBS 0.07509f
C605 VN.t8 VSUBS 0.282609f
C606 VN.n21 VSUBS 0.048087f
C607 VN.n22 VSUBS 0.056274f
C608 VN.t0 VSUBS 0.282609f
C609 VN.n23 VSUBS 0.074975f
C610 VN.t5 VSUBS 0.411797f
C611 VN.t3 VSUBS 0.282609f
C612 VN.n24 VSUBS 0.213479f
C613 VN.n25 VSUBS 0.248558f
C614 VN.n26 VSUBS 0.243662f
C615 VN.n27 VSUBS 0.056274f
C616 VN.n28 VSUBS 0.048087f
C617 VN.n29 VSUBS 0.081017f
C618 VN.n30 VSUBS 0.164119f
C619 VN.n31 VSUBS 0.081017f
C620 VN.n32 VSUBS 0.056274f
C621 VN.n33 VSUBS 0.056274f
C622 VN.n34 VSUBS 0.056274f
C623 VN.n35 VSUBS 0.074975f
C624 VN.n36 VSUBS 0.164119f
C625 VN.n37 VSUBS 0.079089f
C626 VN.t9 VSUBS 0.37258f
C627 VN.n38 VSUBS 0.256837f
C628 VN.n39 VSUBS 1.94889f
.ends

