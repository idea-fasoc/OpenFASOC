* NGSPICE file created from diff_pair_sample_0848.ext - technology: sky130A

.subckt diff_pair_sample_0848 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1170_n2790# sky130_fd_pr__pfet_01v8 ad=3.5451 pd=18.96 as=0 ps=0 w=9.09 l=0.17
X1 B.t8 B.t6 B.t7 w_n1170_n2790# sky130_fd_pr__pfet_01v8 ad=3.5451 pd=18.96 as=0 ps=0 w=9.09 l=0.17
X2 VDD1.t1 VP.t0 VTAIL.t2 w_n1170_n2790# sky130_fd_pr__pfet_01v8 ad=3.5451 pd=18.96 as=3.5451 ps=18.96 w=9.09 l=0.17
X3 B.t5 B.t3 B.t4 w_n1170_n2790# sky130_fd_pr__pfet_01v8 ad=3.5451 pd=18.96 as=0 ps=0 w=9.09 l=0.17
X4 VDD1.t0 VP.t1 VTAIL.t3 w_n1170_n2790# sky130_fd_pr__pfet_01v8 ad=3.5451 pd=18.96 as=3.5451 ps=18.96 w=9.09 l=0.17
X5 VDD2.t1 VN.t0 VTAIL.t1 w_n1170_n2790# sky130_fd_pr__pfet_01v8 ad=3.5451 pd=18.96 as=3.5451 ps=18.96 w=9.09 l=0.17
X6 VDD2.t0 VN.t1 VTAIL.t0 w_n1170_n2790# sky130_fd_pr__pfet_01v8 ad=3.5451 pd=18.96 as=3.5451 ps=18.96 w=9.09 l=0.17
X7 B.t2 B.t0 B.t1 w_n1170_n2790# sky130_fd_pr__pfet_01v8 ad=3.5451 pd=18.96 as=0 ps=0 w=9.09 l=0.17
R0 B.n78 B.t6 1535.62
R1 B.n86 B.t9 1535.62
R2 B.n24 B.t0 1535.62
R3 B.n32 B.t3 1535.62
R4 B.n275 B.n274 585
R5 B.n276 B.n49 585
R6 B.n278 B.n277 585
R7 B.n279 B.n48 585
R8 B.n281 B.n280 585
R9 B.n282 B.n47 585
R10 B.n284 B.n283 585
R11 B.n285 B.n46 585
R12 B.n287 B.n286 585
R13 B.n288 B.n45 585
R14 B.n290 B.n289 585
R15 B.n291 B.n44 585
R16 B.n293 B.n292 585
R17 B.n294 B.n43 585
R18 B.n296 B.n295 585
R19 B.n297 B.n42 585
R20 B.n299 B.n298 585
R21 B.n300 B.n41 585
R22 B.n302 B.n301 585
R23 B.n303 B.n40 585
R24 B.n305 B.n304 585
R25 B.n306 B.n39 585
R26 B.n308 B.n307 585
R27 B.n309 B.n38 585
R28 B.n311 B.n310 585
R29 B.n312 B.n37 585
R30 B.n314 B.n313 585
R31 B.n315 B.n36 585
R32 B.n317 B.n316 585
R33 B.n318 B.n35 585
R34 B.n320 B.n319 585
R35 B.n321 B.n34 585
R36 B.n323 B.n322 585
R37 B.n325 B.n31 585
R38 B.n327 B.n326 585
R39 B.n328 B.n30 585
R40 B.n330 B.n329 585
R41 B.n331 B.n29 585
R42 B.n333 B.n332 585
R43 B.n334 B.n28 585
R44 B.n336 B.n335 585
R45 B.n337 B.n27 585
R46 B.n339 B.n338 585
R47 B.n341 B.n340 585
R48 B.n342 B.n23 585
R49 B.n344 B.n343 585
R50 B.n345 B.n22 585
R51 B.n347 B.n346 585
R52 B.n348 B.n21 585
R53 B.n350 B.n349 585
R54 B.n351 B.n20 585
R55 B.n353 B.n352 585
R56 B.n354 B.n19 585
R57 B.n356 B.n355 585
R58 B.n357 B.n18 585
R59 B.n359 B.n358 585
R60 B.n360 B.n17 585
R61 B.n362 B.n361 585
R62 B.n363 B.n16 585
R63 B.n365 B.n364 585
R64 B.n366 B.n15 585
R65 B.n368 B.n367 585
R66 B.n369 B.n14 585
R67 B.n371 B.n370 585
R68 B.n372 B.n13 585
R69 B.n374 B.n373 585
R70 B.n375 B.n12 585
R71 B.n377 B.n376 585
R72 B.n378 B.n11 585
R73 B.n380 B.n379 585
R74 B.n381 B.n10 585
R75 B.n383 B.n382 585
R76 B.n384 B.n9 585
R77 B.n386 B.n385 585
R78 B.n387 B.n8 585
R79 B.n389 B.n388 585
R80 B.n273 B.n50 585
R81 B.n272 B.n271 585
R82 B.n270 B.n51 585
R83 B.n269 B.n268 585
R84 B.n267 B.n52 585
R85 B.n266 B.n265 585
R86 B.n264 B.n53 585
R87 B.n263 B.n262 585
R88 B.n261 B.n54 585
R89 B.n260 B.n259 585
R90 B.n258 B.n55 585
R91 B.n257 B.n256 585
R92 B.n255 B.n56 585
R93 B.n254 B.n253 585
R94 B.n252 B.n57 585
R95 B.n251 B.n250 585
R96 B.n249 B.n58 585
R97 B.n248 B.n247 585
R98 B.n246 B.n59 585
R99 B.n245 B.n244 585
R100 B.n243 B.n60 585
R101 B.n242 B.n241 585
R102 B.n240 B.n61 585
R103 B.n125 B.n124 585
R104 B.n126 B.n103 585
R105 B.n128 B.n127 585
R106 B.n129 B.n102 585
R107 B.n131 B.n130 585
R108 B.n132 B.n101 585
R109 B.n134 B.n133 585
R110 B.n135 B.n100 585
R111 B.n137 B.n136 585
R112 B.n138 B.n99 585
R113 B.n140 B.n139 585
R114 B.n141 B.n98 585
R115 B.n143 B.n142 585
R116 B.n144 B.n97 585
R117 B.n146 B.n145 585
R118 B.n147 B.n96 585
R119 B.n149 B.n148 585
R120 B.n150 B.n95 585
R121 B.n152 B.n151 585
R122 B.n153 B.n94 585
R123 B.n155 B.n154 585
R124 B.n156 B.n93 585
R125 B.n158 B.n157 585
R126 B.n159 B.n92 585
R127 B.n161 B.n160 585
R128 B.n162 B.n91 585
R129 B.n164 B.n163 585
R130 B.n165 B.n90 585
R131 B.n167 B.n166 585
R132 B.n168 B.n89 585
R133 B.n170 B.n169 585
R134 B.n171 B.n88 585
R135 B.n173 B.n172 585
R136 B.n175 B.n85 585
R137 B.n177 B.n176 585
R138 B.n178 B.n84 585
R139 B.n180 B.n179 585
R140 B.n181 B.n83 585
R141 B.n183 B.n182 585
R142 B.n184 B.n82 585
R143 B.n186 B.n185 585
R144 B.n187 B.n81 585
R145 B.n189 B.n188 585
R146 B.n191 B.n190 585
R147 B.n192 B.n77 585
R148 B.n194 B.n193 585
R149 B.n195 B.n76 585
R150 B.n197 B.n196 585
R151 B.n198 B.n75 585
R152 B.n200 B.n199 585
R153 B.n201 B.n74 585
R154 B.n203 B.n202 585
R155 B.n204 B.n73 585
R156 B.n206 B.n205 585
R157 B.n207 B.n72 585
R158 B.n209 B.n208 585
R159 B.n210 B.n71 585
R160 B.n212 B.n211 585
R161 B.n213 B.n70 585
R162 B.n215 B.n214 585
R163 B.n216 B.n69 585
R164 B.n218 B.n217 585
R165 B.n219 B.n68 585
R166 B.n221 B.n220 585
R167 B.n222 B.n67 585
R168 B.n224 B.n223 585
R169 B.n225 B.n66 585
R170 B.n227 B.n226 585
R171 B.n228 B.n65 585
R172 B.n230 B.n229 585
R173 B.n231 B.n64 585
R174 B.n233 B.n232 585
R175 B.n234 B.n63 585
R176 B.n236 B.n235 585
R177 B.n237 B.n62 585
R178 B.n239 B.n238 585
R179 B.n123 B.n104 585
R180 B.n122 B.n121 585
R181 B.n120 B.n105 585
R182 B.n119 B.n118 585
R183 B.n117 B.n106 585
R184 B.n116 B.n115 585
R185 B.n114 B.n107 585
R186 B.n113 B.n112 585
R187 B.n111 B.n108 585
R188 B.n110 B.n109 585
R189 B.n2 B.n0 585
R190 B.n405 B.n1 585
R191 B.n404 B.n403 585
R192 B.n402 B.n3 585
R193 B.n401 B.n400 585
R194 B.n399 B.n4 585
R195 B.n398 B.n397 585
R196 B.n396 B.n5 585
R197 B.n395 B.n394 585
R198 B.n393 B.n6 585
R199 B.n392 B.n391 585
R200 B.n390 B.n7 585
R201 B.n407 B.n406 585
R202 B.n124 B.n123 492.5
R203 B.n388 B.n7 492.5
R204 B.n238 B.n61 492.5
R205 B.n274 B.n273 492.5
R206 B.n123 B.n122 163.367
R207 B.n122 B.n105 163.367
R208 B.n118 B.n105 163.367
R209 B.n118 B.n117 163.367
R210 B.n117 B.n116 163.367
R211 B.n116 B.n107 163.367
R212 B.n112 B.n107 163.367
R213 B.n112 B.n111 163.367
R214 B.n111 B.n110 163.367
R215 B.n110 B.n2 163.367
R216 B.n406 B.n2 163.367
R217 B.n406 B.n405 163.367
R218 B.n405 B.n404 163.367
R219 B.n404 B.n3 163.367
R220 B.n400 B.n3 163.367
R221 B.n400 B.n399 163.367
R222 B.n399 B.n398 163.367
R223 B.n398 B.n5 163.367
R224 B.n394 B.n5 163.367
R225 B.n394 B.n393 163.367
R226 B.n393 B.n392 163.367
R227 B.n392 B.n7 163.367
R228 B.n124 B.n103 163.367
R229 B.n128 B.n103 163.367
R230 B.n129 B.n128 163.367
R231 B.n130 B.n129 163.367
R232 B.n130 B.n101 163.367
R233 B.n134 B.n101 163.367
R234 B.n135 B.n134 163.367
R235 B.n136 B.n135 163.367
R236 B.n136 B.n99 163.367
R237 B.n140 B.n99 163.367
R238 B.n141 B.n140 163.367
R239 B.n142 B.n141 163.367
R240 B.n142 B.n97 163.367
R241 B.n146 B.n97 163.367
R242 B.n147 B.n146 163.367
R243 B.n148 B.n147 163.367
R244 B.n148 B.n95 163.367
R245 B.n152 B.n95 163.367
R246 B.n153 B.n152 163.367
R247 B.n154 B.n153 163.367
R248 B.n154 B.n93 163.367
R249 B.n158 B.n93 163.367
R250 B.n159 B.n158 163.367
R251 B.n160 B.n159 163.367
R252 B.n160 B.n91 163.367
R253 B.n164 B.n91 163.367
R254 B.n165 B.n164 163.367
R255 B.n166 B.n165 163.367
R256 B.n166 B.n89 163.367
R257 B.n170 B.n89 163.367
R258 B.n171 B.n170 163.367
R259 B.n172 B.n171 163.367
R260 B.n172 B.n85 163.367
R261 B.n177 B.n85 163.367
R262 B.n178 B.n177 163.367
R263 B.n179 B.n178 163.367
R264 B.n179 B.n83 163.367
R265 B.n183 B.n83 163.367
R266 B.n184 B.n183 163.367
R267 B.n185 B.n184 163.367
R268 B.n185 B.n81 163.367
R269 B.n189 B.n81 163.367
R270 B.n190 B.n189 163.367
R271 B.n190 B.n77 163.367
R272 B.n194 B.n77 163.367
R273 B.n195 B.n194 163.367
R274 B.n196 B.n195 163.367
R275 B.n196 B.n75 163.367
R276 B.n200 B.n75 163.367
R277 B.n201 B.n200 163.367
R278 B.n202 B.n201 163.367
R279 B.n202 B.n73 163.367
R280 B.n206 B.n73 163.367
R281 B.n207 B.n206 163.367
R282 B.n208 B.n207 163.367
R283 B.n208 B.n71 163.367
R284 B.n212 B.n71 163.367
R285 B.n213 B.n212 163.367
R286 B.n214 B.n213 163.367
R287 B.n214 B.n69 163.367
R288 B.n218 B.n69 163.367
R289 B.n219 B.n218 163.367
R290 B.n220 B.n219 163.367
R291 B.n220 B.n67 163.367
R292 B.n224 B.n67 163.367
R293 B.n225 B.n224 163.367
R294 B.n226 B.n225 163.367
R295 B.n226 B.n65 163.367
R296 B.n230 B.n65 163.367
R297 B.n231 B.n230 163.367
R298 B.n232 B.n231 163.367
R299 B.n232 B.n63 163.367
R300 B.n236 B.n63 163.367
R301 B.n237 B.n236 163.367
R302 B.n238 B.n237 163.367
R303 B.n242 B.n61 163.367
R304 B.n243 B.n242 163.367
R305 B.n244 B.n243 163.367
R306 B.n244 B.n59 163.367
R307 B.n248 B.n59 163.367
R308 B.n249 B.n248 163.367
R309 B.n250 B.n249 163.367
R310 B.n250 B.n57 163.367
R311 B.n254 B.n57 163.367
R312 B.n255 B.n254 163.367
R313 B.n256 B.n255 163.367
R314 B.n256 B.n55 163.367
R315 B.n260 B.n55 163.367
R316 B.n261 B.n260 163.367
R317 B.n262 B.n261 163.367
R318 B.n262 B.n53 163.367
R319 B.n266 B.n53 163.367
R320 B.n267 B.n266 163.367
R321 B.n268 B.n267 163.367
R322 B.n268 B.n51 163.367
R323 B.n272 B.n51 163.367
R324 B.n273 B.n272 163.367
R325 B.n388 B.n387 163.367
R326 B.n387 B.n386 163.367
R327 B.n386 B.n9 163.367
R328 B.n382 B.n9 163.367
R329 B.n382 B.n381 163.367
R330 B.n381 B.n380 163.367
R331 B.n380 B.n11 163.367
R332 B.n376 B.n11 163.367
R333 B.n376 B.n375 163.367
R334 B.n375 B.n374 163.367
R335 B.n374 B.n13 163.367
R336 B.n370 B.n13 163.367
R337 B.n370 B.n369 163.367
R338 B.n369 B.n368 163.367
R339 B.n368 B.n15 163.367
R340 B.n364 B.n15 163.367
R341 B.n364 B.n363 163.367
R342 B.n363 B.n362 163.367
R343 B.n362 B.n17 163.367
R344 B.n358 B.n17 163.367
R345 B.n358 B.n357 163.367
R346 B.n357 B.n356 163.367
R347 B.n356 B.n19 163.367
R348 B.n352 B.n19 163.367
R349 B.n352 B.n351 163.367
R350 B.n351 B.n350 163.367
R351 B.n350 B.n21 163.367
R352 B.n346 B.n21 163.367
R353 B.n346 B.n345 163.367
R354 B.n345 B.n344 163.367
R355 B.n344 B.n23 163.367
R356 B.n340 B.n23 163.367
R357 B.n340 B.n339 163.367
R358 B.n339 B.n27 163.367
R359 B.n335 B.n27 163.367
R360 B.n335 B.n334 163.367
R361 B.n334 B.n333 163.367
R362 B.n333 B.n29 163.367
R363 B.n329 B.n29 163.367
R364 B.n329 B.n328 163.367
R365 B.n328 B.n327 163.367
R366 B.n327 B.n31 163.367
R367 B.n322 B.n31 163.367
R368 B.n322 B.n321 163.367
R369 B.n321 B.n320 163.367
R370 B.n320 B.n35 163.367
R371 B.n316 B.n35 163.367
R372 B.n316 B.n315 163.367
R373 B.n315 B.n314 163.367
R374 B.n314 B.n37 163.367
R375 B.n310 B.n37 163.367
R376 B.n310 B.n309 163.367
R377 B.n309 B.n308 163.367
R378 B.n308 B.n39 163.367
R379 B.n304 B.n39 163.367
R380 B.n304 B.n303 163.367
R381 B.n303 B.n302 163.367
R382 B.n302 B.n41 163.367
R383 B.n298 B.n41 163.367
R384 B.n298 B.n297 163.367
R385 B.n297 B.n296 163.367
R386 B.n296 B.n43 163.367
R387 B.n292 B.n43 163.367
R388 B.n292 B.n291 163.367
R389 B.n291 B.n290 163.367
R390 B.n290 B.n45 163.367
R391 B.n286 B.n45 163.367
R392 B.n286 B.n285 163.367
R393 B.n285 B.n284 163.367
R394 B.n284 B.n47 163.367
R395 B.n280 B.n47 163.367
R396 B.n280 B.n279 163.367
R397 B.n279 B.n278 163.367
R398 B.n278 B.n49 163.367
R399 B.n274 B.n49 163.367
R400 B.n78 B.t8 122.603
R401 B.n32 B.t4 122.603
R402 B.n86 B.t11 122.594
R403 B.n24 B.t1 122.594
R404 B.n79 B.t7 112.906
R405 B.n33 B.t5 112.906
R406 B.n87 B.t10 112.897
R407 B.n25 B.t2 112.897
R408 B.n80 B.n79 59.5399
R409 B.n174 B.n87 59.5399
R410 B.n26 B.n25 59.5399
R411 B.n324 B.n33 59.5399
R412 B.n390 B.n389 32.0005
R413 B.n275 B.n50 32.0005
R414 B.n240 B.n239 32.0005
R415 B.n125 B.n104 32.0005
R416 B B.n407 18.0485
R417 B.n389 B.n8 10.6151
R418 B.n385 B.n8 10.6151
R419 B.n385 B.n384 10.6151
R420 B.n384 B.n383 10.6151
R421 B.n383 B.n10 10.6151
R422 B.n379 B.n10 10.6151
R423 B.n379 B.n378 10.6151
R424 B.n378 B.n377 10.6151
R425 B.n377 B.n12 10.6151
R426 B.n373 B.n12 10.6151
R427 B.n373 B.n372 10.6151
R428 B.n372 B.n371 10.6151
R429 B.n371 B.n14 10.6151
R430 B.n367 B.n14 10.6151
R431 B.n367 B.n366 10.6151
R432 B.n366 B.n365 10.6151
R433 B.n365 B.n16 10.6151
R434 B.n361 B.n16 10.6151
R435 B.n361 B.n360 10.6151
R436 B.n360 B.n359 10.6151
R437 B.n359 B.n18 10.6151
R438 B.n355 B.n18 10.6151
R439 B.n355 B.n354 10.6151
R440 B.n354 B.n353 10.6151
R441 B.n353 B.n20 10.6151
R442 B.n349 B.n20 10.6151
R443 B.n349 B.n348 10.6151
R444 B.n348 B.n347 10.6151
R445 B.n347 B.n22 10.6151
R446 B.n343 B.n22 10.6151
R447 B.n343 B.n342 10.6151
R448 B.n342 B.n341 10.6151
R449 B.n338 B.n337 10.6151
R450 B.n337 B.n336 10.6151
R451 B.n336 B.n28 10.6151
R452 B.n332 B.n28 10.6151
R453 B.n332 B.n331 10.6151
R454 B.n331 B.n330 10.6151
R455 B.n330 B.n30 10.6151
R456 B.n326 B.n30 10.6151
R457 B.n326 B.n325 10.6151
R458 B.n323 B.n34 10.6151
R459 B.n319 B.n34 10.6151
R460 B.n319 B.n318 10.6151
R461 B.n318 B.n317 10.6151
R462 B.n317 B.n36 10.6151
R463 B.n313 B.n36 10.6151
R464 B.n313 B.n312 10.6151
R465 B.n312 B.n311 10.6151
R466 B.n311 B.n38 10.6151
R467 B.n307 B.n38 10.6151
R468 B.n307 B.n306 10.6151
R469 B.n306 B.n305 10.6151
R470 B.n305 B.n40 10.6151
R471 B.n301 B.n40 10.6151
R472 B.n301 B.n300 10.6151
R473 B.n300 B.n299 10.6151
R474 B.n299 B.n42 10.6151
R475 B.n295 B.n42 10.6151
R476 B.n295 B.n294 10.6151
R477 B.n294 B.n293 10.6151
R478 B.n293 B.n44 10.6151
R479 B.n289 B.n44 10.6151
R480 B.n289 B.n288 10.6151
R481 B.n288 B.n287 10.6151
R482 B.n287 B.n46 10.6151
R483 B.n283 B.n46 10.6151
R484 B.n283 B.n282 10.6151
R485 B.n282 B.n281 10.6151
R486 B.n281 B.n48 10.6151
R487 B.n277 B.n48 10.6151
R488 B.n277 B.n276 10.6151
R489 B.n276 B.n275 10.6151
R490 B.n241 B.n240 10.6151
R491 B.n241 B.n60 10.6151
R492 B.n245 B.n60 10.6151
R493 B.n246 B.n245 10.6151
R494 B.n247 B.n246 10.6151
R495 B.n247 B.n58 10.6151
R496 B.n251 B.n58 10.6151
R497 B.n252 B.n251 10.6151
R498 B.n253 B.n252 10.6151
R499 B.n253 B.n56 10.6151
R500 B.n257 B.n56 10.6151
R501 B.n258 B.n257 10.6151
R502 B.n259 B.n258 10.6151
R503 B.n259 B.n54 10.6151
R504 B.n263 B.n54 10.6151
R505 B.n264 B.n263 10.6151
R506 B.n265 B.n264 10.6151
R507 B.n265 B.n52 10.6151
R508 B.n269 B.n52 10.6151
R509 B.n270 B.n269 10.6151
R510 B.n271 B.n270 10.6151
R511 B.n271 B.n50 10.6151
R512 B.n126 B.n125 10.6151
R513 B.n127 B.n126 10.6151
R514 B.n127 B.n102 10.6151
R515 B.n131 B.n102 10.6151
R516 B.n132 B.n131 10.6151
R517 B.n133 B.n132 10.6151
R518 B.n133 B.n100 10.6151
R519 B.n137 B.n100 10.6151
R520 B.n138 B.n137 10.6151
R521 B.n139 B.n138 10.6151
R522 B.n139 B.n98 10.6151
R523 B.n143 B.n98 10.6151
R524 B.n144 B.n143 10.6151
R525 B.n145 B.n144 10.6151
R526 B.n145 B.n96 10.6151
R527 B.n149 B.n96 10.6151
R528 B.n150 B.n149 10.6151
R529 B.n151 B.n150 10.6151
R530 B.n151 B.n94 10.6151
R531 B.n155 B.n94 10.6151
R532 B.n156 B.n155 10.6151
R533 B.n157 B.n156 10.6151
R534 B.n157 B.n92 10.6151
R535 B.n161 B.n92 10.6151
R536 B.n162 B.n161 10.6151
R537 B.n163 B.n162 10.6151
R538 B.n163 B.n90 10.6151
R539 B.n167 B.n90 10.6151
R540 B.n168 B.n167 10.6151
R541 B.n169 B.n168 10.6151
R542 B.n169 B.n88 10.6151
R543 B.n173 B.n88 10.6151
R544 B.n176 B.n175 10.6151
R545 B.n176 B.n84 10.6151
R546 B.n180 B.n84 10.6151
R547 B.n181 B.n180 10.6151
R548 B.n182 B.n181 10.6151
R549 B.n182 B.n82 10.6151
R550 B.n186 B.n82 10.6151
R551 B.n187 B.n186 10.6151
R552 B.n188 B.n187 10.6151
R553 B.n192 B.n191 10.6151
R554 B.n193 B.n192 10.6151
R555 B.n193 B.n76 10.6151
R556 B.n197 B.n76 10.6151
R557 B.n198 B.n197 10.6151
R558 B.n199 B.n198 10.6151
R559 B.n199 B.n74 10.6151
R560 B.n203 B.n74 10.6151
R561 B.n204 B.n203 10.6151
R562 B.n205 B.n204 10.6151
R563 B.n205 B.n72 10.6151
R564 B.n209 B.n72 10.6151
R565 B.n210 B.n209 10.6151
R566 B.n211 B.n210 10.6151
R567 B.n211 B.n70 10.6151
R568 B.n215 B.n70 10.6151
R569 B.n216 B.n215 10.6151
R570 B.n217 B.n216 10.6151
R571 B.n217 B.n68 10.6151
R572 B.n221 B.n68 10.6151
R573 B.n222 B.n221 10.6151
R574 B.n223 B.n222 10.6151
R575 B.n223 B.n66 10.6151
R576 B.n227 B.n66 10.6151
R577 B.n228 B.n227 10.6151
R578 B.n229 B.n228 10.6151
R579 B.n229 B.n64 10.6151
R580 B.n233 B.n64 10.6151
R581 B.n234 B.n233 10.6151
R582 B.n235 B.n234 10.6151
R583 B.n235 B.n62 10.6151
R584 B.n239 B.n62 10.6151
R585 B.n121 B.n104 10.6151
R586 B.n121 B.n120 10.6151
R587 B.n120 B.n119 10.6151
R588 B.n119 B.n106 10.6151
R589 B.n115 B.n106 10.6151
R590 B.n115 B.n114 10.6151
R591 B.n114 B.n113 10.6151
R592 B.n113 B.n108 10.6151
R593 B.n109 B.n108 10.6151
R594 B.n109 B.n0 10.6151
R595 B.n403 B.n1 10.6151
R596 B.n403 B.n402 10.6151
R597 B.n402 B.n401 10.6151
R598 B.n401 B.n4 10.6151
R599 B.n397 B.n4 10.6151
R600 B.n397 B.n396 10.6151
R601 B.n396 B.n395 10.6151
R602 B.n395 B.n6 10.6151
R603 B.n391 B.n6 10.6151
R604 B.n391 B.n390 10.6151
R605 B.n79 B.n78 9.69747
R606 B.n87 B.n86 9.69747
R607 B.n25 B.n24 9.69747
R608 B.n33 B.n32 9.69747
R609 B.n341 B.n26 8.74196
R610 B.n324 B.n323 8.74196
R611 B.n174 B.n173 8.74196
R612 B.n191 B.n80 8.74196
R613 B.n407 B.n0 2.81026
R614 B.n407 B.n1 2.81026
R615 B.n338 B.n26 1.87367
R616 B.n325 B.n324 1.87367
R617 B.n175 B.n174 1.87367
R618 B.n188 B.n80 1.87367
R619 VP.n0 VP.t1 1695.78
R620 VP.n0 VP.t0 1659.75
R621 VP VP.n0 0.0516364
R622 VTAIL.n1 VTAIL.t0 70.3754
R623 VTAIL.n2 VTAIL.t3 70.3751
R624 VTAIL.n3 VTAIL.t1 70.3751
R625 VTAIL.n0 VTAIL.t2 70.3751
R626 VTAIL.n1 VTAIL.n0 21.0824
R627 VTAIL.n3 VTAIL.n2 20.6514
R628 VTAIL.n2 VTAIL.n1 0.685845
R629 VTAIL VTAIL.n0 0.636276
R630 VTAIL VTAIL.n3 0.050069
R631 VDD1 VDD1.t1 120.061
R632 VDD1 VDD1.t0 87.2199
R633 VN VN.t1 1696.16
R634 VN VN.t0 1659.8
R635 VDD2.n0 VDD2.t1 119.428
R636 VDD2.n0 VDD2.t0 87.0539
R637 VDD2 VDD2.n0 0.166448
C0 VDD1 VP 1.04631f
C1 B VN 0.601431f
C2 VTAIL VN 0.497159f
C3 w_n1170_n2790# B 5.43685f
C4 VP VN 3.79255f
C5 w_n1170_n2790# VTAIL 2.51204f
C6 w_n1170_n2790# VP 1.56143f
C7 VDD2 B 1.12201f
C8 VDD2 VTAIL 6.38367f
C9 VDD2 VP 0.232488f
C10 VDD1 VN 0.148323f
C11 w_n1170_n2790# VDD1 1.29112f
C12 VTAIL B 1.89438f
C13 VP B 0.82809f
C14 w_n1170_n2790# VN 1.41763f
C15 VTAIL VP 0.511808f
C16 VDD2 VDD1 0.421713f
C17 VDD2 VN 0.966173f
C18 w_n1170_n2790# VDD2 1.29059f
C19 VDD1 B 1.11084f
C20 VDD1 VTAIL 6.35377f
C21 VDD2 VSUBS 0.602395f
C22 VDD1 VSUBS 3.605638f
C23 VTAIL VSUBS 0.204332f
C24 VN VSUBS 4.62415f
C25 VP VSUBS 0.853304f
C26 B VSUBS 1.861911f
C27 w_n1170_n2790# VSUBS 40.3931f
C28 VDD2.t1 VSUBS 1.94637f
C29 VDD2.t0 VSUBS 1.57163f
C30 VDD2.n0 VSUBS 2.85398f
C31 VN.t0 VSUBS 0.22427f
C32 VN.t1 VSUBS 0.259663f
C33 VDD1.t0 VSUBS 1.55255f
C34 VDD1.t1 VSUBS 1.94059f
C35 VTAIL.t2 VSUBS 1.90262f
C36 VTAIL.n0 VSUBS 1.93784f
C37 VTAIL.t0 VSUBS 1.90263f
C38 VTAIL.n1 VSUBS 1.94245f
C39 VTAIL.t3 VSUBS 1.90262f
C40 VTAIL.n2 VSUBS 1.9023f
C41 VTAIL.t1 VSUBS 1.90262f
C42 VTAIL.n3 VSUBS 1.84308f
C43 VP.t1 VSUBS 0.263357f
C44 VP.t0 VSUBS 0.228379f
C45 VP.n0 VSUBS 3.30231f
C46 B.n0 VSUBS 0.003937f
C47 B.n1 VSUBS 0.003937f
C48 B.n2 VSUBS 0.006226f
C49 B.n3 VSUBS 0.006226f
C50 B.n4 VSUBS 0.006226f
C51 B.n5 VSUBS 0.006226f
C52 B.n6 VSUBS 0.006226f
C53 B.n7 VSUBS 0.013925f
C54 B.n8 VSUBS 0.006226f
C55 B.n9 VSUBS 0.006226f
C56 B.n10 VSUBS 0.006226f
C57 B.n11 VSUBS 0.006226f
C58 B.n12 VSUBS 0.006226f
C59 B.n13 VSUBS 0.006226f
C60 B.n14 VSUBS 0.006226f
C61 B.n15 VSUBS 0.006226f
C62 B.n16 VSUBS 0.006226f
C63 B.n17 VSUBS 0.006226f
C64 B.n18 VSUBS 0.006226f
C65 B.n19 VSUBS 0.006226f
C66 B.n20 VSUBS 0.006226f
C67 B.n21 VSUBS 0.006226f
C68 B.n22 VSUBS 0.006226f
C69 B.n23 VSUBS 0.006226f
C70 B.t2 VSUBS 0.254444f
C71 B.t1 VSUBS 0.258067f
C72 B.t0 VSUBS 0.0534f
C73 B.n24 VSUBS 0.066352f
C74 B.n25 VSUBS 0.054692f
C75 B.n26 VSUBS 0.014424f
C76 B.n27 VSUBS 0.006226f
C77 B.n28 VSUBS 0.006226f
C78 B.n29 VSUBS 0.006226f
C79 B.n30 VSUBS 0.006226f
C80 B.n31 VSUBS 0.006226f
C81 B.t5 VSUBS 0.254441f
C82 B.t4 VSUBS 0.258064f
C83 B.t3 VSUBS 0.0534f
C84 B.n32 VSUBS 0.066355f
C85 B.n33 VSUBS 0.054695f
C86 B.n34 VSUBS 0.006226f
C87 B.n35 VSUBS 0.006226f
C88 B.n36 VSUBS 0.006226f
C89 B.n37 VSUBS 0.006226f
C90 B.n38 VSUBS 0.006226f
C91 B.n39 VSUBS 0.006226f
C92 B.n40 VSUBS 0.006226f
C93 B.n41 VSUBS 0.006226f
C94 B.n42 VSUBS 0.006226f
C95 B.n43 VSUBS 0.006226f
C96 B.n44 VSUBS 0.006226f
C97 B.n45 VSUBS 0.006226f
C98 B.n46 VSUBS 0.006226f
C99 B.n47 VSUBS 0.006226f
C100 B.n48 VSUBS 0.006226f
C101 B.n49 VSUBS 0.006226f
C102 B.n50 VSUBS 0.014676f
C103 B.n51 VSUBS 0.006226f
C104 B.n52 VSUBS 0.006226f
C105 B.n53 VSUBS 0.006226f
C106 B.n54 VSUBS 0.006226f
C107 B.n55 VSUBS 0.006226f
C108 B.n56 VSUBS 0.006226f
C109 B.n57 VSUBS 0.006226f
C110 B.n58 VSUBS 0.006226f
C111 B.n59 VSUBS 0.006226f
C112 B.n60 VSUBS 0.006226f
C113 B.n61 VSUBS 0.013925f
C114 B.n62 VSUBS 0.006226f
C115 B.n63 VSUBS 0.006226f
C116 B.n64 VSUBS 0.006226f
C117 B.n65 VSUBS 0.006226f
C118 B.n66 VSUBS 0.006226f
C119 B.n67 VSUBS 0.006226f
C120 B.n68 VSUBS 0.006226f
C121 B.n69 VSUBS 0.006226f
C122 B.n70 VSUBS 0.006226f
C123 B.n71 VSUBS 0.006226f
C124 B.n72 VSUBS 0.006226f
C125 B.n73 VSUBS 0.006226f
C126 B.n74 VSUBS 0.006226f
C127 B.n75 VSUBS 0.006226f
C128 B.n76 VSUBS 0.006226f
C129 B.n77 VSUBS 0.006226f
C130 B.t7 VSUBS 0.254441f
C131 B.t8 VSUBS 0.258064f
C132 B.t6 VSUBS 0.0534f
C133 B.n78 VSUBS 0.066355f
C134 B.n79 VSUBS 0.054695f
C135 B.n80 VSUBS 0.014424f
C136 B.n81 VSUBS 0.006226f
C137 B.n82 VSUBS 0.006226f
C138 B.n83 VSUBS 0.006226f
C139 B.n84 VSUBS 0.006226f
C140 B.n85 VSUBS 0.006226f
C141 B.t10 VSUBS 0.254444f
C142 B.t11 VSUBS 0.258067f
C143 B.t9 VSUBS 0.0534f
C144 B.n86 VSUBS 0.066352f
C145 B.n87 VSUBS 0.054692f
C146 B.n88 VSUBS 0.006226f
C147 B.n89 VSUBS 0.006226f
C148 B.n90 VSUBS 0.006226f
C149 B.n91 VSUBS 0.006226f
C150 B.n92 VSUBS 0.006226f
C151 B.n93 VSUBS 0.006226f
C152 B.n94 VSUBS 0.006226f
C153 B.n95 VSUBS 0.006226f
C154 B.n96 VSUBS 0.006226f
C155 B.n97 VSUBS 0.006226f
C156 B.n98 VSUBS 0.006226f
C157 B.n99 VSUBS 0.006226f
C158 B.n100 VSUBS 0.006226f
C159 B.n101 VSUBS 0.006226f
C160 B.n102 VSUBS 0.006226f
C161 B.n103 VSUBS 0.006226f
C162 B.n104 VSUBS 0.013925f
C163 B.n105 VSUBS 0.006226f
C164 B.n106 VSUBS 0.006226f
C165 B.n107 VSUBS 0.006226f
C166 B.n108 VSUBS 0.006226f
C167 B.n109 VSUBS 0.006226f
C168 B.n110 VSUBS 0.006226f
C169 B.n111 VSUBS 0.006226f
C170 B.n112 VSUBS 0.006226f
C171 B.n113 VSUBS 0.006226f
C172 B.n114 VSUBS 0.006226f
C173 B.n115 VSUBS 0.006226f
C174 B.n116 VSUBS 0.006226f
C175 B.n117 VSUBS 0.006226f
C176 B.n118 VSUBS 0.006226f
C177 B.n119 VSUBS 0.006226f
C178 B.n120 VSUBS 0.006226f
C179 B.n121 VSUBS 0.006226f
C180 B.n122 VSUBS 0.006226f
C181 B.n123 VSUBS 0.013925f
C182 B.n124 VSUBS 0.014823f
C183 B.n125 VSUBS 0.014823f
C184 B.n126 VSUBS 0.006226f
C185 B.n127 VSUBS 0.006226f
C186 B.n128 VSUBS 0.006226f
C187 B.n129 VSUBS 0.006226f
C188 B.n130 VSUBS 0.006226f
C189 B.n131 VSUBS 0.006226f
C190 B.n132 VSUBS 0.006226f
C191 B.n133 VSUBS 0.006226f
C192 B.n134 VSUBS 0.006226f
C193 B.n135 VSUBS 0.006226f
C194 B.n136 VSUBS 0.006226f
C195 B.n137 VSUBS 0.006226f
C196 B.n138 VSUBS 0.006226f
C197 B.n139 VSUBS 0.006226f
C198 B.n140 VSUBS 0.006226f
C199 B.n141 VSUBS 0.006226f
C200 B.n142 VSUBS 0.006226f
C201 B.n143 VSUBS 0.006226f
C202 B.n144 VSUBS 0.006226f
C203 B.n145 VSUBS 0.006226f
C204 B.n146 VSUBS 0.006226f
C205 B.n147 VSUBS 0.006226f
C206 B.n148 VSUBS 0.006226f
C207 B.n149 VSUBS 0.006226f
C208 B.n150 VSUBS 0.006226f
C209 B.n151 VSUBS 0.006226f
C210 B.n152 VSUBS 0.006226f
C211 B.n153 VSUBS 0.006226f
C212 B.n154 VSUBS 0.006226f
C213 B.n155 VSUBS 0.006226f
C214 B.n156 VSUBS 0.006226f
C215 B.n157 VSUBS 0.006226f
C216 B.n158 VSUBS 0.006226f
C217 B.n159 VSUBS 0.006226f
C218 B.n160 VSUBS 0.006226f
C219 B.n161 VSUBS 0.006226f
C220 B.n162 VSUBS 0.006226f
C221 B.n163 VSUBS 0.006226f
C222 B.n164 VSUBS 0.006226f
C223 B.n165 VSUBS 0.006226f
C224 B.n166 VSUBS 0.006226f
C225 B.n167 VSUBS 0.006226f
C226 B.n168 VSUBS 0.006226f
C227 B.n169 VSUBS 0.006226f
C228 B.n170 VSUBS 0.006226f
C229 B.n171 VSUBS 0.006226f
C230 B.n172 VSUBS 0.006226f
C231 B.n173 VSUBS 0.005676f
C232 B.n174 VSUBS 0.014424f
C233 B.n175 VSUBS 0.003662f
C234 B.n176 VSUBS 0.006226f
C235 B.n177 VSUBS 0.006226f
C236 B.n178 VSUBS 0.006226f
C237 B.n179 VSUBS 0.006226f
C238 B.n180 VSUBS 0.006226f
C239 B.n181 VSUBS 0.006226f
C240 B.n182 VSUBS 0.006226f
C241 B.n183 VSUBS 0.006226f
C242 B.n184 VSUBS 0.006226f
C243 B.n185 VSUBS 0.006226f
C244 B.n186 VSUBS 0.006226f
C245 B.n187 VSUBS 0.006226f
C246 B.n188 VSUBS 0.003662f
C247 B.n189 VSUBS 0.006226f
C248 B.n190 VSUBS 0.006226f
C249 B.n191 VSUBS 0.005676f
C250 B.n192 VSUBS 0.006226f
C251 B.n193 VSUBS 0.006226f
C252 B.n194 VSUBS 0.006226f
C253 B.n195 VSUBS 0.006226f
C254 B.n196 VSUBS 0.006226f
C255 B.n197 VSUBS 0.006226f
C256 B.n198 VSUBS 0.006226f
C257 B.n199 VSUBS 0.006226f
C258 B.n200 VSUBS 0.006226f
C259 B.n201 VSUBS 0.006226f
C260 B.n202 VSUBS 0.006226f
C261 B.n203 VSUBS 0.006226f
C262 B.n204 VSUBS 0.006226f
C263 B.n205 VSUBS 0.006226f
C264 B.n206 VSUBS 0.006226f
C265 B.n207 VSUBS 0.006226f
C266 B.n208 VSUBS 0.006226f
C267 B.n209 VSUBS 0.006226f
C268 B.n210 VSUBS 0.006226f
C269 B.n211 VSUBS 0.006226f
C270 B.n212 VSUBS 0.006226f
C271 B.n213 VSUBS 0.006226f
C272 B.n214 VSUBS 0.006226f
C273 B.n215 VSUBS 0.006226f
C274 B.n216 VSUBS 0.006226f
C275 B.n217 VSUBS 0.006226f
C276 B.n218 VSUBS 0.006226f
C277 B.n219 VSUBS 0.006226f
C278 B.n220 VSUBS 0.006226f
C279 B.n221 VSUBS 0.006226f
C280 B.n222 VSUBS 0.006226f
C281 B.n223 VSUBS 0.006226f
C282 B.n224 VSUBS 0.006226f
C283 B.n225 VSUBS 0.006226f
C284 B.n226 VSUBS 0.006226f
C285 B.n227 VSUBS 0.006226f
C286 B.n228 VSUBS 0.006226f
C287 B.n229 VSUBS 0.006226f
C288 B.n230 VSUBS 0.006226f
C289 B.n231 VSUBS 0.006226f
C290 B.n232 VSUBS 0.006226f
C291 B.n233 VSUBS 0.006226f
C292 B.n234 VSUBS 0.006226f
C293 B.n235 VSUBS 0.006226f
C294 B.n236 VSUBS 0.006226f
C295 B.n237 VSUBS 0.006226f
C296 B.n238 VSUBS 0.014823f
C297 B.n239 VSUBS 0.014823f
C298 B.n240 VSUBS 0.013925f
C299 B.n241 VSUBS 0.006226f
C300 B.n242 VSUBS 0.006226f
C301 B.n243 VSUBS 0.006226f
C302 B.n244 VSUBS 0.006226f
C303 B.n245 VSUBS 0.006226f
C304 B.n246 VSUBS 0.006226f
C305 B.n247 VSUBS 0.006226f
C306 B.n248 VSUBS 0.006226f
C307 B.n249 VSUBS 0.006226f
C308 B.n250 VSUBS 0.006226f
C309 B.n251 VSUBS 0.006226f
C310 B.n252 VSUBS 0.006226f
C311 B.n253 VSUBS 0.006226f
C312 B.n254 VSUBS 0.006226f
C313 B.n255 VSUBS 0.006226f
C314 B.n256 VSUBS 0.006226f
C315 B.n257 VSUBS 0.006226f
C316 B.n258 VSUBS 0.006226f
C317 B.n259 VSUBS 0.006226f
C318 B.n260 VSUBS 0.006226f
C319 B.n261 VSUBS 0.006226f
C320 B.n262 VSUBS 0.006226f
C321 B.n263 VSUBS 0.006226f
C322 B.n264 VSUBS 0.006226f
C323 B.n265 VSUBS 0.006226f
C324 B.n266 VSUBS 0.006226f
C325 B.n267 VSUBS 0.006226f
C326 B.n268 VSUBS 0.006226f
C327 B.n269 VSUBS 0.006226f
C328 B.n270 VSUBS 0.006226f
C329 B.n271 VSUBS 0.006226f
C330 B.n272 VSUBS 0.006226f
C331 B.n273 VSUBS 0.013925f
C332 B.n274 VSUBS 0.014823f
C333 B.n275 VSUBS 0.014072f
C334 B.n276 VSUBS 0.006226f
C335 B.n277 VSUBS 0.006226f
C336 B.n278 VSUBS 0.006226f
C337 B.n279 VSUBS 0.006226f
C338 B.n280 VSUBS 0.006226f
C339 B.n281 VSUBS 0.006226f
C340 B.n282 VSUBS 0.006226f
C341 B.n283 VSUBS 0.006226f
C342 B.n284 VSUBS 0.006226f
C343 B.n285 VSUBS 0.006226f
C344 B.n286 VSUBS 0.006226f
C345 B.n287 VSUBS 0.006226f
C346 B.n288 VSUBS 0.006226f
C347 B.n289 VSUBS 0.006226f
C348 B.n290 VSUBS 0.006226f
C349 B.n291 VSUBS 0.006226f
C350 B.n292 VSUBS 0.006226f
C351 B.n293 VSUBS 0.006226f
C352 B.n294 VSUBS 0.006226f
C353 B.n295 VSUBS 0.006226f
C354 B.n296 VSUBS 0.006226f
C355 B.n297 VSUBS 0.006226f
C356 B.n298 VSUBS 0.006226f
C357 B.n299 VSUBS 0.006226f
C358 B.n300 VSUBS 0.006226f
C359 B.n301 VSUBS 0.006226f
C360 B.n302 VSUBS 0.006226f
C361 B.n303 VSUBS 0.006226f
C362 B.n304 VSUBS 0.006226f
C363 B.n305 VSUBS 0.006226f
C364 B.n306 VSUBS 0.006226f
C365 B.n307 VSUBS 0.006226f
C366 B.n308 VSUBS 0.006226f
C367 B.n309 VSUBS 0.006226f
C368 B.n310 VSUBS 0.006226f
C369 B.n311 VSUBS 0.006226f
C370 B.n312 VSUBS 0.006226f
C371 B.n313 VSUBS 0.006226f
C372 B.n314 VSUBS 0.006226f
C373 B.n315 VSUBS 0.006226f
C374 B.n316 VSUBS 0.006226f
C375 B.n317 VSUBS 0.006226f
C376 B.n318 VSUBS 0.006226f
C377 B.n319 VSUBS 0.006226f
C378 B.n320 VSUBS 0.006226f
C379 B.n321 VSUBS 0.006226f
C380 B.n322 VSUBS 0.006226f
C381 B.n323 VSUBS 0.005676f
C382 B.n324 VSUBS 0.014424f
C383 B.n325 VSUBS 0.003662f
C384 B.n326 VSUBS 0.006226f
C385 B.n327 VSUBS 0.006226f
C386 B.n328 VSUBS 0.006226f
C387 B.n329 VSUBS 0.006226f
C388 B.n330 VSUBS 0.006226f
C389 B.n331 VSUBS 0.006226f
C390 B.n332 VSUBS 0.006226f
C391 B.n333 VSUBS 0.006226f
C392 B.n334 VSUBS 0.006226f
C393 B.n335 VSUBS 0.006226f
C394 B.n336 VSUBS 0.006226f
C395 B.n337 VSUBS 0.006226f
C396 B.n338 VSUBS 0.003662f
C397 B.n339 VSUBS 0.006226f
C398 B.n340 VSUBS 0.006226f
C399 B.n341 VSUBS 0.005676f
C400 B.n342 VSUBS 0.006226f
C401 B.n343 VSUBS 0.006226f
C402 B.n344 VSUBS 0.006226f
C403 B.n345 VSUBS 0.006226f
C404 B.n346 VSUBS 0.006226f
C405 B.n347 VSUBS 0.006226f
C406 B.n348 VSUBS 0.006226f
C407 B.n349 VSUBS 0.006226f
C408 B.n350 VSUBS 0.006226f
C409 B.n351 VSUBS 0.006226f
C410 B.n352 VSUBS 0.006226f
C411 B.n353 VSUBS 0.006226f
C412 B.n354 VSUBS 0.006226f
C413 B.n355 VSUBS 0.006226f
C414 B.n356 VSUBS 0.006226f
C415 B.n357 VSUBS 0.006226f
C416 B.n358 VSUBS 0.006226f
C417 B.n359 VSUBS 0.006226f
C418 B.n360 VSUBS 0.006226f
C419 B.n361 VSUBS 0.006226f
C420 B.n362 VSUBS 0.006226f
C421 B.n363 VSUBS 0.006226f
C422 B.n364 VSUBS 0.006226f
C423 B.n365 VSUBS 0.006226f
C424 B.n366 VSUBS 0.006226f
C425 B.n367 VSUBS 0.006226f
C426 B.n368 VSUBS 0.006226f
C427 B.n369 VSUBS 0.006226f
C428 B.n370 VSUBS 0.006226f
C429 B.n371 VSUBS 0.006226f
C430 B.n372 VSUBS 0.006226f
C431 B.n373 VSUBS 0.006226f
C432 B.n374 VSUBS 0.006226f
C433 B.n375 VSUBS 0.006226f
C434 B.n376 VSUBS 0.006226f
C435 B.n377 VSUBS 0.006226f
C436 B.n378 VSUBS 0.006226f
C437 B.n379 VSUBS 0.006226f
C438 B.n380 VSUBS 0.006226f
C439 B.n381 VSUBS 0.006226f
C440 B.n382 VSUBS 0.006226f
C441 B.n383 VSUBS 0.006226f
C442 B.n384 VSUBS 0.006226f
C443 B.n385 VSUBS 0.006226f
C444 B.n386 VSUBS 0.006226f
C445 B.n387 VSUBS 0.006226f
C446 B.n388 VSUBS 0.014823f
C447 B.n389 VSUBS 0.014823f
C448 B.n390 VSUBS 0.013925f
C449 B.n391 VSUBS 0.006226f
C450 B.n392 VSUBS 0.006226f
C451 B.n393 VSUBS 0.006226f
C452 B.n394 VSUBS 0.006226f
C453 B.n395 VSUBS 0.006226f
C454 B.n396 VSUBS 0.006226f
C455 B.n397 VSUBS 0.006226f
C456 B.n398 VSUBS 0.006226f
C457 B.n399 VSUBS 0.006226f
C458 B.n400 VSUBS 0.006226f
C459 B.n401 VSUBS 0.006226f
C460 B.n402 VSUBS 0.006226f
C461 B.n403 VSUBS 0.006226f
C462 B.n404 VSUBS 0.006226f
C463 B.n405 VSUBS 0.006226f
C464 B.n406 VSUBS 0.006226f
C465 B.n407 VSUBS 0.014097f
.ends

