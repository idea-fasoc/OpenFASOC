* NGSPICE file created from diff_pair_sample_1469.ext - technology: sky130A

.subckt diff_pair_sample_1469 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=2.9913 pd=16.12 as=1.26555 ps=8 w=7.67 l=3.45
X1 VDD1.t7 VP.t1 VTAIL.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=1.26555 pd=8 as=2.9913 ps=16.12 w=7.67 l=3.45
X2 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=2.9913 pd=16.12 as=0 ps=0 w=7.67 l=3.45
X3 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=2.9913 pd=16.12 as=0 ps=0 w=7.67 l=3.45
X4 VDD1.t6 VP.t2 VTAIL.t13 B.t1 sky130_fd_pr__nfet_01v8 ad=1.26555 pd=8 as=1.26555 ps=8 w=7.67 l=3.45
X5 VTAIL.t3 VN.t0 VDD2.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.26555 pd=8 as=1.26555 ps=8 w=7.67 l=3.45
X6 VDD2.t6 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.26555 pd=8 as=1.26555 ps=8 w=7.67 l=3.45
X7 VDD2.t5 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.26555 pd=8 as=1.26555 ps=8 w=7.67 l=3.45
X8 VDD1.t2 VP.t3 VTAIL.t12 B.t0 sky130_fd_pr__nfet_01v8 ad=1.26555 pd=8 as=2.9913 ps=16.12 w=7.67 l=3.45
X9 VTAIL.t11 VP.t4 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.26555 pd=8 as=1.26555 ps=8 w=7.67 l=3.45
X10 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=2.9913 pd=16.12 as=0 ps=0 w=7.67 l=3.45
X11 VDD2.t4 VN.t3 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.26555 pd=8 as=2.9913 ps=16.12 w=7.67 l=3.45
X12 VTAIL.t6 VN.t4 VDD2.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=1.26555 pd=8 as=1.26555 ps=8 w=7.67 l=3.45
X13 VTAIL.t10 VP.t5 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.9913 pd=16.12 as=1.26555 ps=8 w=7.67 l=3.45
X14 VDD1.t1 VP.t6 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=1.26555 pd=8 as=1.26555 ps=8 w=7.67 l=3.45
X15 VDD2.t2 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.26555 pd=8 as=2.9913 ps=16.12 w=7.67 l=3.45
X16 VTAIL.t8 VP.t7 VDD1.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=1.26555 pd=8 as=1.26555 ps=8 w=7.67 l=3.45
X17 VTAIL.t5 VN.t6 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=2.9913 pd=16.12 as=1.26555 ps=8 w=7.67 l=3.45
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.9913 pd=16.12 as=0 ps=0 w=7.67 l=3.45
X19 VTAIL.t4 VN.t7 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=2.9913 pd=16.12 as=1.26555 ps=8 w=7.67 l=3.45
R0 VP.n24 VP.n23 161.3
R1 VP.n25 VP.n20 161.3
R2 VP.n27 VP.n26 161.3
R3 VP.n28 VP.n19 161.3
R4 VP.n30 VP.n29 161.3
R5 VP.n31 VP.n18 161.3
R6 VP.n34 VP.n33 161.3
R7 VP.n35 VP.n17 161.3
R8 VP.n37 VP.n36 161.3
R9 VP.n38 VP.n16 161.3
R10 VP.n40 VP.n39 161.3
R11 VP.n41 VP.n15 161.3
R12 VP.n43 VP.n42 161.3
R13 VP.n44 VP.n14 161.3
R14 VP.n46 VP.n45 161.3
R15 VP.n85 VP.n84 161.3
R16 VP.n83 VP.n1 161.3
R17 VP.n82 VP.n81 161.3
R18 VP.n80 VP.n2 161.3
R19 VP.n79 VP.n78 161.3
R20 VP.n77 VP.n3 161.3
R21 VP.n76 VP.n75 161.3
R22 VP.n74 VP.n4 161.3
R23 VP.n73 VP.n72 161.3
R24 VP.n70 VP.n5 161.3
R25 VP.n69 VP.n68 161.3
R26 VP.n67 VP.n6 161.3
R27 VP.n66 VP.n65 161.3
R28 VP.n64 VP.n7 161.3
R29 VP.n63 VP.n62 161.3
R30 VP.n61 VP.n60 161.3
R31 VP.n59 VP.n9 161.3
R32 VP.n58 VP.n57 161.3
R33 VP.n56 VP.n10 161.3
R34 VP.n55 VP.n54 161.3
R35 VP.n53 VP.n11 161.3
R36 VP.n52 VP.n51 161.3
R37 VP.n50 VP.n12 161.3
R38 VP.n22 VP.t5 86.6911
R39 VP.n49 VP.n48 81.7486
R40 VP.n86 VP.n0 81.7486
R41 VP.n47 VP.n13 81.7486
R42 VP.n54 VP.n10 56.5193
R43 VP.n78 VP.n2 56.5193
R44 VP.n39 VP.n15 56.5193
R45 VP.n22 VP.n21 55.4655
R46 VP.n48 VP.t0 53.5793
R47 VP.n8 VP.t6 53.5793
R48 VP.n71 VP.t4 53.5793
R49 VP.n0 VP.t1 53.5793
R50 VP.n13 VP.t3 53.5793
R51 VP.n32 VP.t7 53.5793
R52 VP.n21 VP.t2 53.5793
R53 VP.n49 VP.n47 51.6433
R54 VP.n65 VP.n6 40.4934
R55 VP.n69 VP.n6 40.4934
R56 VP.n30 VP.n19 40.4934
R57 VP.n26 VP.n19 40.4934
R58 VP.n52 VP.n12 24.4675
R59 VP.n53 VP.n52 24.4675
R60 VP.n54 VP.n53 24.4675
R61 VP.n58 VP.n10 24.4675
R62 VP.n59 VP.n58 24.4675
R63 VP.n60 VP.n59 24.4675
R64 VP.n64 VP.n63 24.4675
R65 VP.n65 VP.n64 24.4675
R66 VP.n70 VP.n69 24.4675
R67 VP.n72 VP.n70 24.4675
R68 VP.n76 VP.n4 24.4675
R69 VP.n77 VP.n76 24.4675
R70 VP.n78 VP.n77 24.4675
R71 VP.n82 VP.n2 24.4675
R72 VP.n83 VP.n82 24.4675
R73 VP.n84 VP.n83 24.4675
R74 VP.n43 VP.n15 24.4675
R75 VP.n44 VP.n43 24.4675
R76 VP.n45 VP.n44 24.4675
R77 VP.n31 VP.n30 24.4675
R78 VP.n33 VP.n31 24.4675
R79 VP.n37 VP.n17 24.4675
R80 VP.n38 VP.n37 24.4675
R81 VP.n39 VP.n38 24.4675
R82 VP.n25 VP.n24 24.4675
R83 VP.n26 VP.n25 24.4675
R84 VP.n63 VP.n8 19.0848
R85 VP.n72 VP.n71 19.0848
R86 VP.n33 VP.n32 19.0848
R87 VP.n24 VP.n21 19.0848
R88 VP.n48 VP.n12 8.31928
R89 VP.n84 VP.n0 8.31928
R90 VP.n45 VP.n13 8.31928
R91 VP.n60 VP.n8 5.38324
R92 VP.n71 VP.n4 5.38324
R93 VP.n32 VP.n17 5.38324
R94 VP.n23 VP.n22 3.21182
R95 VP.n47 VP.n46 0.354971
R96 VP.n50 VP.n49 0.354971
R97 VP.n86 VP.n85 0.354971
R98 VP VP.n86 0.26696
R99 VP.n23 VP.n20 0.189894
R100 VP.n27 VP.n20 0.189894
R101 VP.n28 VP.n27 0.189894
R102 VP.n29 VP.n28 0.189894
R103 VP.n29 VP.n18 0.189894
R104 VP.n34 VP.n18 0.189894
R105 VP.n35 VP.n34 0.189894
R106 VP.n36 VP.n35 0.189894
R107 VP.n36 VP.n16 0.189894
R108 VP.n40 VP.n16 0.189894
R109 VP.n41 VP.n40 0.189894
R110 VP.n42 VP.n41 0.189894
R111 VP.n42 VP.n14 0.189894
R112 VP.n46 VP.n14 0.189894
R113 VP.n51 VP.n50 0.189894
R114 VP.n51 VP.n11 0.189894
R115 VP.n55 VP.n11 0.189894
R116 VP.n56 VP.n55 0.189894
R117 VP.n57 VP.n56 0.189894
R118 VP.n57 VP.n9 0.189894
R119 VP.n61 VP.n9 0.189894
R120 VP.n62 VP.n61 0.189894
R121 VP.n62 VP.n7 0.189894
R122 VP.n66 VP.n7 0.189894
R123 VP.n67 VP.n66 0.189894
R124 VP.n68 VP.n67 0.189894
R125 VP.n68 VP.n5 0.189894
R126 VP.n73 VP.n5 0.189894
R127 VP.n74 VP.n73 0.189894
R128 VP.n75 VP.n74 0.189894
R129 VP.n75 VP.n3 0.189894
R130 VP.n79 VP.n3 0.189894
R131 VP.n80 VP.n79 0.189894
R132 VP.n81 VP.n80 0.189894
R133 VP.n81 VP.n1 0.189894
R134 VP.n85 VP.n1 0.189894
R135 VDD1 VDD1.n0 70.4394
R136 VDD1.n3 VDD1.n2 70.3257
R137 VDD1.n3 VDD1.n1 70.3257
R138 VDD1.n5 VDD1.n4 68.7517
R139 VDD1.n5 VDD1.n3 45.5742
R140 VDD1.n4 VDD1.t4 2.58199
R141 VDD1.n4 VDD1.t2 2.58199
R142 VDD1.n0 VDD1.t5 2.58199
R143 VDD1.n0 VDD1.t6 2.58199
R144 VDD1.n2 VDD1.t3 2.58199
R145 VDD1.n2 VDD1.t7 2.58199
R146 VDD1.n1 VDD1.t0 2.58199
R147 VDD1.n1 VDD1.t1 2.58199
R148 VDD1 VDD1.n5 1.57162
R149 VTAIL.n11 VTAIL.t10 54.6546
R150 VTAIL.n10 VTAIL.t7 54.6546
R151 VTAIL.n7 VTAIL.t5 54.6546
R152 VTAIL.n15 VTAIL.t0 54.6544
R153 VTAIL.n2 VTAIL.t4 54.6544
R154 VTAIL.n3 VTAIL.t14 54.6544
R155 VTAIL.n6 VTAIL.t15 54.6544
R156 VTAIL.n14 VTAIL.t12 54.6544
R157 VTAIL.n13 VTAIL.n12 52.0731
R158 VTAIL.n9 VTAIL.n8 52.0731
R159 VTAIL.n1 VTAIL.n0 52.0729
R160 VTAIL.n5 VTAIL.n4 52.0729
R161 VTAIL.n15 VTAIL.n14 22.2376
R162 VTAIL.n7 VTAIL.n6 22.2376
R163 VTAIL.n9 VTAIL.n7 3.25912
R164 VTAIL.n10 VTAIL.n9 3.25912
R165 VTAIL.n13 VTAIL.n11 3.25912
R166 VTAIL.n14 VTAIL.n13 3.25912
R167 VTAIL.n6 VTAIL.n5 3.25912
R168 VTAIL.n5 VTAIL.n3 3.25912
R169 VTAIL.n2 VTAIL.n1 3.25912
R170 VTAIL VTAIL.n15 3.20093
R171 VTAIL.n0 VTAIL.t1 2.58199
R172 VTAIL.n0 VTAIL.t6 2.58199
R173 VTAIL.n4 VTAIL.t9 2.58199
R174 VTAIL.n4 VTAIL.t11 2.58199
R175 VTAIL.n12 VTAIL.t13 2.58199
R176 VTAIL.n12 VTAIL.t8 2.58199
R177 VTAIL.n8 VTAIL.t2 2.58199
R178 VTAIL.n8 VTAIL.t3 2.58199
R179 VTAIL.n11 VTAIL.n10 0.470328
R180 VTAIL.n3 VTAIL.n2 0.470328
R181 VTAIL VTAIL.n1 0.0586897
R182 B.n853 B.n852 585
R183 B.n854 B.n853 585
R184 B.n284 B.n150 585
R185 B.n283 B.n282 585
R186 B.n281 B.n280 585
R187 B.n279 B.n278 585
R188 B.n277 B.n276 585
R189 B.n275 B.n274 585
R190 B.n273 B.n272 585
R191 B.n271 B.n270 585
R192 B.n269 B.n268 585
R193 B.n267 B.n266 585
R194 B.n265 B.n264 585
R195 B.n263 B.n262 585
R196 B.n261 B.n260 585
R197 B.n259 B.n258 585
R198 B.n257 B.n256 585
R199 B.n255 B.n254 585
R200 B.n253 B.n252 585
R201 B.n251 B.n250 585
R202 B.n249 B.n248 585
R203 B.n247 B.n246 585
R204 B.n245 B.n244 585
R205 B.n243 B.n242 585
R206 B.n241 B.n240 585
R207 B.n239 B.n238 585
R208 B.n237 B.n236 585
R209 B.n235 B.n234 585
R210 B.n233 B.n232 585
R211 B.n231 B.n230 585
R212 B.n229 B.n228 585
R213 B.n227 B.n226 585
R214 B.n225 B.n224 585
R215 B.n223 B.n222 585
R216 B.n221 B.n220 585
R217 B.n219 B.n218 585
R218 B.n217 B.n216 585
R219 B.n215 B.n214 585
R220 B.n213 B.n212 585
R221 B.n210 B.n209 585
R222 B.n208 B.n207 585
R223 B.n206 B.n205 585
R224 B.n204 B.n203 585
R225 B.n202 B.n201 585
R226 B.n200 B.n199 585
R227 B.n198 B.n197 585
R228 B.n196 B.n195 585
R229 B.n194 B.n193 585
R230 B.n192 B.n191 585
R231 B.n190 B.n189 585
R232 B.n188 B.n187 585
R233 B.n186 B.n185 585
R234 B.n184 B.n183 585
R235 B.n182 B.n181 585
R236 B.n180 B.n179 585
R237 B.n178 B.n177 585
R238 B.n176 B.n175 585
R239 B.n174 B.n173 585
R240 B.n172 B.n171 585
R241 B.n170 B.n169 585
R242 B.n168 B.n167 585
R243 B.n166 B.n165 585
R244 B.n164 B.n163 585
R245 B.n162 B.n161 585
R246 B.n160 B.n159 585
R247 B.n158 B.n157 585
R248 B.n117 B.n116 585
R249 B.n857 B.n856 585
R250 B.n851 B.n151 585
R251 B.n151 B.n114 585
R252 B.n850 B.n113 585
R253 B.n861 B.n113 585
R254 B.n849 B.n112 585
R255 B.n862 B.n112 585
R256 B.n848 B.n111 585
R257 B.n863 B.n111 585
R258 B.n847 B.n846 585
R259 B.n846 B.n107 585
R260 B.n845 B.n106 585
R261 B.n869 B.n106 585
R262 B.n844 B.n105 585
R263 B.n870 B.n105 585
R264 B.n843 B.n104 585
R265 B.n871 B.n104 585
R266 B.n842 B.n841 585
R267 B.n841 B.n103 585
R268 B.n840 B.n99 585
R269 B.n877 B.n99 585
R270 B.n839 B.n98 585
R271 B.n878 B.n98 585
R272 B.n838 B.n97 585
R273 B.n879 B.n97 585
R274 B.n837 B.n836 585
R275 B.n836 B.n93 585
R276 B.n835 B.n92 585
R277 B.n885 B.n92 585
R278 B.n834 B.n91 585
R279 B.n886 B.n91 585
R280 B.n833 B.n90 585
R281 B.n887 B.n90 585
R282 B.n832 B.n831 585
R283 B.n831 B.n86 585
R284 B.n830 B.n85 585
R285 B.n893 B.n85 585
R286 B.n829 B.n84 585
R287 B.n894 B.n84 585
R288 B.n828 B.n83 585
R289 B.n895 B.n83 585
R290 B.n827 B.n826 585
R291 B.n826 B.n79 585
R292 B.n825 B.n78 585
R293 B.n901 B.n78 585
R294 B.n824 B.n77 585
R295 B.n902 B.n77 585
R296 B.n823 B.n76 585
R297 B.n903 B.n76 585
R298 B.n822 B.n821 585
R299 B.n821 B.n72 585
R300 B.n820 B.n71 585
R301 B.n909 B.n71 585
R302 B.n819 B.n70 585
R303 B.n910 B.n70 585
R304 B.n818 B.n69 585
R305 B.n911 B.n69 585
R306 B.n817 B.n816 585
R307 B.n816 B.n65 585
R308 B.n815 B.n64 585
R309 B.n917 B.n64 585
R310 B.n814 B.n63 585
R311 B.n918 B.n63 585
R312 B.n813 B.n62 585
R313 B.n919 B.n62 585
R314 B.n812 B.n811 585
R315 B.n811 B.n58 585
R316 B.n810 B.n57 585
R317 B.n925 B.n57 585
R318 B.n809 B.n56 585
R319 B.n926 B.n56 585
R320 B.n808 B.n55 585
R321 B.n927 B.n55 585
R322 B.n807 B.n806 585
R323 B.n806 B.n51 585
R324 B.n805 B.n50 585
R325 B.n933 B.n50 585
R326 B.n804 B.n49 585
R327 B.n934 B.n49 585
R328 B.n803 B.n48 585
R329 B.n935 B.n48 585
R330 B.n802 B.n801 585
R331 B.n801 B.n44 585
R332 B.n800 B.n43 585
R333 B.n941 B.n43 585
R334 B.n799 B.n42 585
R335 B.n942 B.n42 585
R336 B.n798 B.n41 585
R337 B.n943 B.n41 585
R338 B.n797 B.n796 585
R339 B.n796 B.n37 585
R340 B.n795 B.n36 585
R341 B.n949 B.n36 585
R342 B.n794 B.n35 585
R343 B.n950 B.n35 585
R344 B.n793 B.n34 585
R345 B.n951 B.n34 585
R346 B.n792 B.n791 585
R347 B.n791 B.n30 585
R348 B.n790 B.n29 585
R349 B.n957 B.n29 585
R350 B.n789 B.n28 585
R351 B.n958 B.n28 585
R352 B.n788 B.n27 585
R353 B.n959 B.n27 585
R354 B.n787 B.n786 585
R355 B.n786 B.n23 585
R356 B.n785 B.n22 585
R357 B.n965 B.n22 585
R358 B.n784 B.n21 585
R359 B.n966 B.n21 585
R360 B.n783 B.n20 585
R361 B.n967 B.n20 585
R362 B.n782 B.n781 585
R363 B.n781 B.n19 585
R364 B.n780 B.n15 585
R365 B.n973 B.n15 585
R366 B.n779 B.n14 585
R367 B.n974 B.n14 585
R368 B.n778 B.n13 585
R369 B.n975 B.n13 585
R370 B.n777 B.n776 585
R371 B.n776 B.n12 585
R372 B.n775 B.n774 585
R373 B.n775 B.n8 585
R374 B.n773 B.n7 585
R375 B.n982 B.n7 585
R376 B.n772 B.n6 585
R377 B.n983 B.n6 585
R378 B.n771 B.n5 585
R379 B.n984 B.n5 585
R380 B.n770 B.n769 585
R381 B.n769 B.n4 585
R382 B.n768 B.n285 585
R383 B.n768 B.n767 585
R384 B.n758 B.n286 585
R385 B.n287 B.n286 585
R386 B.n760 B.n759 585
R387 B.n761 B.n760 585
R388 B.n757 B.n292 585
R389 B.n292 B.n291 585
R390 B.n756 B.n755 585
R391 B.n755 B.n754 585
R392 B.n294 B.n293 585
R393 B.n747 B.n294 585
R394 B.n746 B.n745 585
R395 B.n748 B.n746 585
R396 B.n744 B.n299 585
R397 B.n299 B.n298 585
R398 B.n743 B.n742 585
R399 B.n742 B.n741 585
R400 B.n301 B.n300 585
R401 B.n302 B.n301 585
R402 B.n734 B.n733 585
R403 B.n735 B.n734 585
R404 B.n732 B.n307 585
R405 B.n307 B.n306 585
R406 B.n731 B.n730 585
R407 B.n730 B.n729 585
R408 B.n309 B.n308 585
R409 B.n310 B.n309 585
R410 B.n722 B.n721 585
R411 B.n723 B.n722 585
R412 B.n720 B.n315 585
R413 B.n315 B.n314 585
R414 B.n719 B.n718 585
R415 B.n718 B.n717 585
R416 B.n317 B.n316 585
R417 B.n318 B.n317 585
R418 B.n710 B.n709 585
R419 B.n711 B.n710 585
R420 B.n708 B.n323 585
R421 B.n323 B.n322 585
R422 B.n707 B.n706 585
R423 B.n706 B.n705 585
R424 B.n325 B.n324 585
R425 B.n326 B.n325 585
R426 B.n698 B.n697 585
R427 B.n699 B.n698 585
R428 B.n696 B.n331 585
R429 B.n331 B.n330 585
R430 B.n695 B.n694 585
R431 B.n694 B.n693 585
R432 B.n333 B.n332 585
R433 B.n334 B.n333 585
R434 B.n686 B.n685 585
R435 B.n687 B.n686 585
R436 B.n684 B.n338 585
R437 B.n342 B.n338 585
R438 B.n683 B.n682 585
R439 B.n682 B.n681 585
R440 B.n340 B.n339 585
R441 B.n341 B.n340 585
R442 B.n674 B.n673 585
R443 B.n675 B.n674 585
R444 B.n672 B.n347 585
R445 B.n347 B.n346 585
R446 B.n671 B.n670 585
R447 B.n670 B.n669 585
R448 B.n349 B.n348 585
R449 B.n350 B.n349 585
R450 B.n662 B.n661 585
R451 B.n663 B.n662 585
R452 B.n660 B.n355 585
R453 B.n355 B.n354 585
R454 B.n659 B.n658 585
R455 B.n658 B.n657 585
R456 B.n357 B.n356 585
R457 B.n358 B.n357 585
R458 B.n650 B.n649 585
R459 B.n651 B.n650 585
R460 B.n648 B.n362 585
R461 B.n366 B.n362 585
R462 B.n647 B.n646 585
R463 B.n646 B.n645 585
R464 B.n364 B.n363 585
R465 B.n365 B.n364 585
R466 B.n638 B.n637 585
R467 B.n639 B.n638 585
R468 B.n636 B.n371 585
R469 B.n371 B.n370 585
R470 B.n635 B.n634 585
R471 B.n634 B.n633 585
R472 B.n373 B.n372 585
R473 B.n374 B.n373 585
R474 B.n626 B.n625 585
R475 B.n627 B.n626 585
R476 B.n624 B.n379 585
R477 B.n379 B.n378 585
R478 B.n623 B.n622 585
R479 B.n622 B.n621 585
R480 B.n381 B.n380 585
R481 B.n382 B.n381 585
R482 B.n614 B.n613 585
R483 B.n615 B.n614 585
R484 B.n612 B.n387 585
R485 B.n387 B.n386 585
R486 B.n611 B.n610 585
R487 B.n610 B.n609 585
R488 B.n389 B.n388 585
R489 B.n602 B.n389 585
R490 B.n601 B.n600 585
R491 B.n603 B.n601 585
R492 B.n599 B.n394 585
R493 B.n394 B.n393 585
R494 B.n598 B.n597 585
R495 B.n597 B.n596 585
R496 B.n396 B.n395 585
R497 B.n397 B.n396 585
R498 B.n589 B.n588 585
R499 B.n590 B.n589 585
R500 B.n587 B.n402 585
R501 B.n402 B.n401 585
R502 B.n586 B.n585 585
R503 B.n585 B.n584 585
R504 B.n404 B.n403 585
R505 B.n405 B.n404 585
R506 B.n580 B.n579 585
R507 B.n408 B.n407 585
R508 B.n576 B.n575 585
R509 B.n577 B.n576 585
R510 B.n574 B.n441 585
R511 B.n573 B.n572 585
R512 B.n571 B.n570 585
R513 B.n569 B.n568 585
R514 B.n567 B.n566 585
R515 B.n565 B.n564 585
R516 B.n563 B.n562 585
R517 B.n561 B.n560 585
R518 B.n559 B.n558 585
R519 B.n557 B.n556 585
R520 B.n555 B.n554 585
R521 B.n553 B.n552 585
R522 B.n551 B.n550 585
R523 B.n549 B.n548 585
R524 B.n547 B.n546 585
R525 B.n545 B.n544 585
R526 B.n543 B.n542 585
R527 B.n541 B.n540 585
R528 B.n539 B.n538 585
R529 B.n537 B.n536 585
R530 B.n535 B.n534 585
R531 B.n533 B.n532 585
R532 B.n531 B.n530 585
R533 B.n529 B.n528 585
R534 B.n527 B.n526 585
R535 B.n525 B.n524 585
R536 B.n523 B.n522 585
R537 B.n521 B.n520 585
R538 B.n519 B.n518 585
R539 B.n517 B.n516 585
R540 B.n515 B.n514 585
R541 B.n513 B.n512 585
R542 B.n511 B.n510 585
R543 B.n509 B.n508 585
R544 B.n507 B.n506 585
R545 B.n504 B.n503 585
R546 B.n502 B.n501 585
R547 B.n500 B.n499 585
R548 B.n498 B.n497 585
R549 B.n496 B.n495 585
R550 B.n494 B.n493 585
R551 B.n492 B.n491 585
R552 B.n490 B.n489 585
R553 B.n488 B.n487 585
R554 B.n486 B.n485 585
R555 B.n484 B.n483 585
R556 B.n482 B.n481 585
R557 B.n480 B.n479 585
R558 B.n478 B.n477 585
R559 B.n476 B.n475 585
R560 B.n474 B.n473 585
R561 B.n472 B.n471 585
R562 B.n470 B.n469 585
R563 B.n468 B.n467 585
R564 B.n466 B.n465 585
R565 B.n464 B.n463 585
R566 B.n462 B.n461 585
R567 B.n460 B.n459 585
R568 B.n458 B.n457 585
R569 B.n456 B.n455 585
R570 B.n454 B.n453 585
R571 B.n452 B.n451 585
R572 B.n450 B.n449 585
R573 B.n448 B.n447 585
R574 B.n581 B.n406 585
R575 B.n406 B.n405 585
R576 B.n583 B.n582 585
R577 B.n584 B.n583 585
R578 B.n400 B.n399 585
R579 B.n401 B.n400 585
R580 B.n592 B.n591 585
R581 B.n591 B.n590 585
R582 B.n593 B.n398 585
R583 B.n398 B.n397 585
R584 B.n595 B.n594 585
R585 B.n596 B.n595 585
R586 B.n392 B.n391 585
R587 B.n393 B.n392 585
R588 B.n605 B.n604 585
R589 B.n604 B.n603 585
R590 B.n606 B.n390 585
R591 B.n602 B.n390 585
R592 B.n608 B.n607 585
R593 B.n609 B.n608 585
R594 B.n385 B.n384 585
R595 B.n386 B.n385 585
R596 B.n617 B.n616 585
R597 B.n616 B.n615 585
R598 B.n618 B.n383 585
R599 B.n383 B.n382 585
R600 B.n620 B.n619 585
R601 B.n621 B.n620 585
R602 B.n377 B.n376 585
R603 B.n378 B.n377 585
R604 B.n629 B.n628 585
R605 B.n628 B.n627 585
R606 B.n630 B.n375 585
R607 B.n375 B.n374 585
R608 B.n632 B.n631 585
R609 B.n633 B.n632 585
R610 B.n369 B.n368 585
R611 B.n370 B.n369 585
R612 B.n641 B.n640 585
R613 B.n640 B.n639 585
R614 B.n642 B.n367 585
R615 B.n367 B.n365 585
R616 B.n644 B.n643 585
R617 B.n645 B.n644 585
R618 B.n361 B.n360 585
R619 B.n366 B.n361 585
R620 B.n653 B.n652 585
R621 B.n652 B.n651 585
R622 B.n654 B.n359 585
R623 B.n359 B.n358 585
R624 B.n656 B.n655 585
R625 B.n657 B.n656 585
R626 B.n353 B.n352 585
R627 B.n354 B.n353 585
R628 B.n665 B.n664 585
R629 B.n664 B.n663 585
R630 B.n666 B.n351 585
R631 B.n351 B.n350 585
R632 B.n668 B.n667 585
R633 B.n669 B.n668 585
R634 B.n345 B.n344 585
R635 B.n346 B.n345 585
R636 B.n677 B.n676 585
R637 B.n676 B.n675 585
R638 B.n678 B.n343 585
R639 B.n343 B.n341 585
R640 B.n680 B.n679 585
R641 B.n681 B.n680 585
R642 B.n337 B.n336 585
R643 B.n342 B.n337 585
R644 B.n689 B.n688 585
R645 B.n688 B.n687 585
R646 B.n690 B.n335 585
R647 B.n335 B.n334 585
R648 B.n692 B.n691 585
R649 B.n693 B.n692 585
R650 B.n329 B.n328 585
R651 B.n330 B.n329 585
R652 B.n701 B.n700 585
R653 B.n700 B.n699 585
R654 B.n702 B.n327 585
R655 B.n327 B.n326 585
R656 B.n704 B.n703 585
R657 B.n705 B.n704 585
R658 B.n321 B.n320 585
R659 B.n322 B.n321 585
R660 B.n713 B.n712 585
R661 B.n712 B.n711 585
R662 B.n714 B.n319 585
R663 B.n319 B.n318 585
R664 B.n716 B.n715 585
R665 B.n717 B.n716 585
R666 B.n313 B.n312 585
R667 B.n314 B.n313 585
R668 B.n725 B.n724 585
R669 B.n724 B.n723 585
R670 B.n726 B.n311 585
R671 B.n311 B.n310 585
R672 B.n728 B.n727 585
R673 B.n729 B.n728 585
R674 B.n305 B.n304 585
R675 B.n306 B.n305 585
R676 B.n737 B.n736 585
R677 B.n736 B.n735 585
R678 B.n738 B.n303 585
R679 B.n303 B.n302 585
R680 B.n740 B.n739 585
R681 B.n741 B.n740 585
R682 B.n297 B.n296 585
R683 B.n298 B.n297 585
R684 B.n750 B.n749 585
R685 B.n749 B.n748 585
R686 B.n751 B.n295 585
R687 B.n747 B.n295 585
R688 B.n753 B.n752 585
R689 B.n754 B.n753 585
R690 B.n290 B.n289 585
R691 B.n291 B.n290 585
R692 B.n763 B.n762 585
R693 B.n762 B.n761 585
R694 B.n764 B.n288 585
R695 B.n288 B.n287 585
R696 B.n766 B.n765 585
R697 B.n767 B.n766 585
R698 B.n3 B.n0 585
R699 B.n4 B.n3 585
R700 B.n981 B.n1 585
R701 B.n982 B.n981 585
R702 B.n980 B.n979 585
R703 B.n980 B.n8 585
R704 B.n978 B.n9 585
R705 B.n12 B.n9 585
R706 B.n977 B.n976 585
R707 B.n976 B.n975 585
R708 B.n11 B.n10 585
R709 B.n974 B.n11 585
R710 B.n972 B.n971 585
R711 B.n973 B.n972 585
R712 B.n970 B.n16 585
R713 B.n19 B.n16 585
R714 B.n969 B.n968 585
R715 B.n968 B.n967 585
R716 B.n18 B.n17 585
R717 B.n966 B.n18 585
R718 B.n964 B.n963 585
R719 B.n965 B.n964 585
R720 B.n962 B.n24 585
R721 B.n24 B.n23 585
R722 B.n961 B.n960 585
R723 B.n960 B.n959 585
R724 B.n26 B.n25 585
R725 B.n958 B.n26 585
R726 B.n956 B.n955 585
R727 B.n957 B.n956 585
R728 B.n954 B.n31 585
R729 B.n31 B.n30 585
R730 B.n953 B.n952 585
R731 B.n952 B.n951 585
R732 B.n33 B.n32 585
R733 B.n950 B.n33 585
R734 B.n948 B.n947 585
R735 B.n949 B.n948 585
R736 B.n946 B.n38 585
R737 B.n38 B.n37 585
R738 B.n945 B.n944 585
R739 B.n944 B.n943 585
R740 B.n40 B.n39 585
R741 B.n942 B.n40 585
R742 B.n940 B.n939 585
R743 B.n941 B.n940 585
R744 B.n938 B.n45 585
R745 B.n45 B.n44 585
R746 B.n937 B.n936 585
R747 B.n936 B.n935 585
R748 B.n47 B.n46 585
R749 B.n934 B.n47 585
R750 B.n932 B.n931 585
R751 B.n933 B.n932 585
R752 B.n930 B.n52 585
R753 B.n52 B.n51 585
R754 B.n929 B.n928 585
R755 B.n928 B.n927 585
R756 B.n54 B.n53 585
R757 B.n926 B.n54 585
R758 B.n924 B.n923 585
R759 B.n925 B.n924 585
R760 B.n922 B.n59 585
R761 B.n59 B.n58 585
R762 B.n921 B.n920 585
R763 B.n920 B.n919 585
R764 B.n61 B.n60 585
R765 B.n918 B.n61 585
R766 B.n916 B.n915 585
R767 B.n917 B.n916 585
R768 B.n914 B.n66 585
R769 B.n66 B.n65 585
R770 B.n913 B.n912 585
R771 B.n912 B.n911 585
R772 B.n68 B.n67 585
R773 B.n910 B.n68 585
R774 B.n908 B.n907 585
R775 B.n909 B.n908 585
R776 B.n906 B.n73 585
R777 B.n73 B.n72 585
R778 B.n905 B.n904 585
R779 B.n904 B.n903 585
R780 B.n75 B.n74 585
R781 B.n902 B.n75 585
R782 B.n900 B.n899 585
R783 B.n901 B.n900 585
R784 B.n898 B.n80 585
R785 B.n80 B.n79 585
R786 B.n897 B.n896 585
R787 B.n896 B.n895 585
R788 B.n82 B.n81 585
R789 B.n894 B.n82 585
R790 B.n892 B.n891 585
R791 B.n893 B.n892 585
R792 B.n890 B.n87 585
R793 B.n87 B.n86 585
R794 B.n889 B.n888 585
R795 B.n888 B.n887 585
R796 B.n89 B.n88 585
R797 B.n886 B.n89 585
R798 B.n884 B.n883 585
R799 B.n885 B.n884 585
R800 B.n882 B.n94 585
R801 B.n94 B.n93 585
R802 B.n881 B.n880 585
R803 B.n880 B.n879 585
R804 B.n96 B.n95 585
R805 B.n878 B.n96 585
R806 B.n876 B.n875 585
R807 B.n877 B.n876 585
R808 B.n874 B.n100 585
R809 B.n103 B.n100 585
R810 B.n873 B.n872 585
R811 B.n872 B.n871 585
R812 B.n102 B.n101 585
R813 B.n870 B.n102 585
R814 B.n868 B.n867 585
R815 B.n869 B.n868 585
R816 B.n866 B.n108 585
R817 B.n108 B.n107 585
R818 B.n865 B.n864 585
R819 B.n864 B.n863 585
R820 B.n110 B.n109 585
R821 B.n862 B.n110 585
R822 B.n860 B.n859 585
R823 B.n861 B.n860 585
R824 B.n858 B.n115 585
R825 B.n115 B.n114 585
R826 B.n985 B.n984 585
R827 B.n983 B.n2 585
R828 B.n856 B.n115 559.769
R829 B.n853 B.n151 559.769
R830 B.n447 B.n404 559.769
R831 B.n579 B.n406 559.769
R832 B.n155 B.t12 262.627
R833 B.n152 B.t19 262.627
R834 B.n445 B.t16 262.627
R835 B.n442 B.t8 262.627
R836 B.n854 B.n149 256.663
R837 B.n854 B.n148 256.663
R838 B.n854 B.n147 256.663
R839 B.n854 B.n146 256.663
R840 B.n854 B.n145 256.663
R841 B.n854 B.n144 256.663
R842 B.n854 B.n143 256.663
R843 B.n854 B.n142 256.663
R844 B.n854 B.n141 256.663
R845 B.n854 B.n140 256.663
R846 B.n854 B.n139 256.663
R847 B.n854 B.n138 256.663
R848 B.n854 B.n137 256.663
R849 B.n854 B.n136 256.663
R850 B.n854 B.n135 256.663
R851 B.n854 B.n134 256.663
R852 B.n854 B.n133 256.663
R853 B.n854 B.n132 256.663
R854 B.n854 B.n131 256.663
R855 B.n854 B.n130 256.663
R856 B.n854 B.n129 256.663
R857 B.n854 B.n128 256.663
R858 B.n854 B.n127 256.663
R859 B.n854 B.n126 256.663
R860 B.n854 B.n125 256.663
R861 B.n854 B.n124 256.663
R862 B.n854 B.n123 256.663
R863 B.n854 B.n122 256.663
R864 B.n854 B.n121 256.663
R865 B.n854 B.n120 256.663
R866 B.n854 B.n119 256.663
R867 B.n854 B.n118 256.663
R868 B.n855 B.n854 256.663
R869 B.n578 B.n577 256.663
R870 B.n577 B.n409 256.663
R871 B.n577 B.n410 256.663
R872 B.n577 B.n411 256.663
R873 B.n577 B.n412 256.663
R874 B.n577 B.n413 256.663
R875 B.n577 B.n414 256.663
R876 B.n577 B.n415 256.663
R877 B.n577 B.n416 256.663
R878 B.n577 B.n417 256.663
R879 B.n577 B.n418 256.663
R880 B.n577 B.n419 256.663
R881 B.n577 B.n420 256.663
R882 B.n577 B.n421 256.663
R883 B.n577 B.n422 256.663
R884 B.n577 B.n423 256.663
R885 B.n577 B.n424 256.663
R886 B.n577 B.n425 256.663
R887 B.n577 B.n426 256.663
R888 B.n577 B.n427 256.663
R889 B.n577 B.n428 256.663
R890 B.n577 B.n429 256.663
R891 B.n577 B.n430 256.663
R892 B.n577 B.n431 256.663
R893 B.n577 B.n432 256.663
R894 B.n577 B.n433 256.663
R895 B.n577 B.n434 256.663
R896 B.n577 B.n435 256.663
R897 B.n577 B.n436 256.663
R898 B.n577 B.n437 256.663
R899 B.n577 B.n438 256.663
R900 B.n577 B.n439 256.663
R901 B.n577 B.n440 256.663
R902 B.n987 B.n986 256.663
R903 B.n157 B.n117 163.367
R904 B.n161 B.n160 163.367
R905 B.n165 B.n164 163.367
R906 B.n169 B.n168 163.367
R907 B.n173 B.n172 163.367
R908 B.n177 B.n176 163.367
R909 B.n181 B.n180 163.367
R910 B.n185 B.n184 163.367
R911 B.n189 B.n188 163.367
R912 B.n193 B.n192 163.367
R913 B.n197 B.n196 163.367
R914 B.n201 B.n200 163.367
R915 B.n205 B.n204 163.367
R916 B.n209 B.n208 163.367
R917 B.n214 B.n213 163.367
R918 B.n218 B.n217 163.367
R919 B.n222 B.n221 163.367
R920 B.n226 B.n225 163.367
R921 B.n230 B.n229 163.367
R922 B.n234 B.n233 163.367
R923 B.n238 B.n237 163.367
R924 B.n242 B.n241 163.367
R925 B.n246 B.n245 163.367
R926 B.n250 B.n249 163.367
R927 B.n254 B.n253 163.367
R928 B.n258 B.n257 163.367
R929 B.n262 B.n261 163.367
R930 B.n266 B.n265 163.367
R931 B.n270 B.n269 163.367
R932 B.n274 B.n273 163.367
R933 B.n278 B.n277 163.367
R934 B.n282 B.n281 163.367
R935 B.n853 B.n150 163.367
R936 B.n585 B.n404 163.367
R937 B.n585 B.n402 163.367
R938 B.n589 B.n402 163.367
R939 B.n589 B.n396 163.367
R940 B.n597 B.n396 163.367
R941 B.n597 B.n394 163.367
R942 B.n601 B.n394 163.367
R943 B.n601 B.n389 163.367
R944 B.n610 B.n389 163.367
R945 B.n610 B.n387 163.367
R946 B.n614 B.n387 163.367
R947 B.n614 B.n381 163.367
R948 B.n622 B.n381 163.367
R949 B.n622 B.n379 163.367
R950 B.n626 B.n379 163.367
R951 B.n626 B.n373 163.367
R952 B.n634 B.n373 163.367
R953 B.n634 B.n371 163.367
R954 B.n638 B.n371 163.367
R955 B.n638 B.n364 163.367
R956 B.n646 B.n364 163.367
R957 B.n646 B.n362 163.367
R958 B.n650 B.n362 163.367
R959 B.n650 B.n357 163.367
R960 B.n658 B.n357 163.367
R961 B.n658 B.n355 163.367
R962 B.n662 B.n355 163.367
R963 B.n662 B.n349 163.367
R964 B.n670 B.n349 163.367
R965 B.n670 B.n347 163.367
R966 B.n674 B.n347 163.367
R967 B.n674 B.n340 163.367
R968 B.n682 B.n340 163.367
R969 B.n682 B.n338 163.367
R970 B.n686 B.n338 163.367
R971 B.n686 B.n333 163.367
R972 B.n694 B.n333 163.367
R973 B.n694 B.n331 163.367
R974 B.n698 B.n331 163.367
R975 B.n698 B.n325 163.367
R976 B.n706 B.n325 163.367
R977 B.n706 B.n323 163.367
R978 B.n710 B.n323 163.367
R979 B.n710 B.n317 163.367
R980 B.n718 B.n317 163.367
R981 B.n718 B.n315 163.367
R982 B.n722 B.n315 163.367
R983 B.n722 B.n309 163.367
R984 B.n730 B.n309 163.367
R985 B.n730 B.n307 163.367
R986 B.n734 B.n307 163.367
R987 B.n734 B.n301 163.367
R988 B.n742 B.n301 163.367
R989 B.n742 B.n299 163.367
R990 B.n746 B.n299 163.367
R991 B.n746 B.n294 163.367
R992 B.n755 B.n294 163.367
R993 B.n755 B.n292 163.367
R994 B.n760 B.n292 163.367
R995 B.n760 B.n286 163.367
R996 B.n768 B.n286 163.367
R997 B.n769 B.n768 163.367
R998 B.n769 B.n5 163.367
R999 B.n6 B.n5 163.367
R1000 B.n7 B.n6 163.367
R1001 B.n775 B.n7 163.367
R1002 B.n776 B.n775 163.367
R1003 B.n776 B.n13 163.367
R1004 B.n14 B.n13 163.367
R1005 B.n15 B.n14 163.367
R1006 B.n781 B.n15 163.367
R1007 B.n781 B.n20 163.367
R1008 B.n21 B.n20 163.367
R1009 B.n22 B.n21 163.367
R1010 B.n786 B.n22 163.367
R1011 B.n786 B.n27 163.367
R1012 B.n28 B.n27 163.367
R1013 B.n29 B.n28 163.367
R1014 B.n791 B.n29 163.367
R1015 B.n791 B.n34 163.367
R1016 B.n35 B.n34 163.367
R1017 B.n36 B.n35 163.367
R1018 B.n796 B.n36 163.367
R1019 B.n796 B.n41 163.367
R1020 B.n42 B.n41 163.367
R1021 B.n43 B.n42 163.367
R1022 B.n801 B.n43 163.367
R1023 B.n801 B.n48 163.367
R1024 B.n49 B.n48 163.367
R1025 B.n50 B.n49 163.367
R1026 B.n806 B.n50 163.367
R1027 B.n806 B.n55 163.367
R1028 B.n56 B.n55 163.367
R1029 B.n57 B.n56 163.367
R1030 B.n811 B.n57 163.367
R1031 B.n811 B.n62 163.367
R1032 B.n63 B.n62 163.367
R1033 B.n64 B.n63 163.367
R1034 B.n816 B.n64 163.367
R1035 B.n816 B.n69 163.367
R1036 B.n70 B.n69 163.367
R1037 B.n71 B.n70 163.367
R1038 B.n821 B.n71 163.367
R1039 B.n821 B.n76 163.367
R1040 B.n77 B.n76 163.367
R1041 B.n78 B.n77 163.367
R1042 B.n826 B.n78 163.367
R1043 B.n826 B.n83 163.367
R1044 B.n84 B.n83 163.367
R1045 B.n85 B.n84 163.367
R1046 B.n831 B.n85 163.367
R1047 B.n831 B.n90 163.367
R1048 B.n91 B.n90 163.367
R1049 B.n92 B.n91 163.367
R1050 B.n836 B.n92 163.367
R1051 B.n836 B.n97 163.367
R1052 B.n98 B.n97 163.367
R1053 B.n99 B.n98 163.367
R1054 B.n841 B.n99 163.367
R1055 B.n841 B.n104 163.367
R1056 B.n105 B.n104 163.367
R1057 B.n106 B.n105 163.367
R1058 B.n846 B.n106 163.367
R1059 B.n846 B.n111 163.367
R1060 B.n112 B.n111 163.367
R1061 B.n113 B.n112 163.367
R1062 B.n151 B.n113 163.367
R1063 B.n576 B.n408 163.367
R1064 B.n576 B.n441 163.367
R1065 B.n572 B.n571 163.367
R1066 B.n568 B.n567 163.367
R1067 B.n564 B.n563 163.367
R1068 B.n560 B.n559 163.367
R1069 B.n556 B.n555 163.367
R1070 B.n552 B.n551 163.367
R1071 B.n548 B.n547 163.367
R1072 B.n544 B.n543 163.367
R1073 B.n540 B.n539 163.367
R1074 B.n536 B.n535 163.367
R1075 B.n532 B.n531 163.367
R1076 B.n528 B.n527 163.367
R1077 B.n524 B.n523 163.367
R1078 B.n520 B.n519 163.367
R1079 B.n516 B.n515 163.367
R1080 B.n512 B.n511 163.367
R1081 B.n508 B.n507 163.367
R1082 B.n503 B.n502 163.367
R1083 B.n499 B.n498 163.367
R1084 B.n495 B.n494 163.367
R1085 B.n491 B.n490 163.367
R1086 B.n487 B.n486 163.367
R1087 B.n483 B.n482 163.367
R1088 B.n479 B.n478 163.367
R1089 B.n475 B.n474 163.367
R1090 B.n471 B.n470 163.367
R1091 B.n467 B.n466 163.367
R1092 B.n463 B.n462 163.367
R1093 B.n459 B.n458 163.367
R1094 B.n455 B.n454 163.367
R1095 B.n451 B.n450 163.367
R1096 B.n583 B.n406 163.367
R1097 B.n583 B.n400 163.367
R1098 B.n591 B.n400 163.367
R1099 B.n591 B.n398 163.367
R1100 B.n595 B.n398 163.367
R1101 B.n595 B.n392 163.367
R1102 B.n604 B.n392 163.367
R1103 B.n604 B.n390 163.367
R1104 B.n608 B.n390 163.367
R1105 B.n608 B.n385 163.367
R1106 B.n616 B.n385 163.367
R1107 B.n616 B.n383 163.367
R1108 B.n620 B.n383 163.367
R1109 B.n620 B.n377 163.367
R1110 B.n628 B.n377 163.367
R1111 B.n628 B.n375 163.367
R1112 B.n632 B.n375 163.367
R1113 B.n632 B.n369 163.367
R1114 B.n640 B.n369 163.367
R1115 B.n640 B.n367 163.367
R1116 B.n644 B.n367 163.367
R1117 B.n644 B.n361 163.367
R1118 B.n652 B.n361 163.367
R1119 B.n652 B.n359 163.367
R1120 B.n656 B.n359 163.367
R1121 B.n656 B.n353 163.367
R1122 B.n664 B.n353 163.367
R1123 B.n664 B.n351 163.367
R1124 B.n668 B.n351 163.367
R1125 B.n668 B.n345 163.367
R1126 B.n676 B.n345 163.367
R1127 B.n676 B.n343 163.367
R1128 B.n680 B.n343 163.367
R1129 B.n680 B.n337 163.367
R1130 B.n688 B.n337 163.367
R1131 B.n688 B.n335 163.367
R1132 B.n692 B.n335 163.367
R1133 B.n692 B.n329 163.367
R1134 B.n700 B.n329 163.367
R1135 B.n700 B.n327 163.367
R1136 B.n704 B.n327 163.367
R1137 B.n704 B.n321 163.367
R1138 B.n712 B.n321 163.367
R1139 B.n712 B.n319 163.367
R1140 B.n716 B.n319 163.367
R1141 B.n716 B.n313 163.367
R1142 B.n724 B.n313 163.367
R1143 B.n724 B.n311 163.367
R1144 B.n728 B.n311 163.367
R1145 B.n728 B.n305 163.367
R1146 B.n736 B.n305 163.367
R1147 B.n736 B.n303 163.367
R1148 B.n740 B.n303 163.367
R1149 B.n740 B.n297 163.367
R1150 B.n749 B.n297 163.367
R1151 B.n749 B.n295 163.367
R1152 B.n753 B.n295 163.367
R1153 B.n753 B.n290 163.367
R1154 B.n762 B.n290 163.367
R1155 B.n762 B.n288 163.367
R1156 B.n766 B.n288 163.367
R1157 B.n766 B.n3 163.367
R1158 B.n985 B.n3 163.367
R1159 B.n981 B.n2 163.367
R1160 B.n981 B.n980 163.367
R1161 B.n980 B.n9 163.367
R1162 B.n976 B.n9 163.367
R1163 B.n976 B.n11 163.367
R1164 B.n972 B.n11 163.367
R1165 B.n972 B.n16 163.367
R1166 B.n968 B.n16 163.367
R1167 B.n968 B.n18 163.367
R1168 B.n964 B.n18 163.367
R1169 B.n964 B.n24 163.367
R1170 B.n960 B.n24 163.367
R1171 B.n960 B.n26 163.367
R1172 B.n956 B.n26 163.367
R1173 B.n956 B.n31 163.367
R1174 B.n952 B.n31 163.367
R1175 B.n952 B.n33 163.367
R1176 B.n948 B.n33 163.367
R1177 B.n948 B.n38 163.367
R1178 B.n944 B.n38 163.367
R1179 B.n944 B.n40 163.367
R1180 B.n940 B.n40 163.367
R1181 B.n940 B.n45 163.367
R1182 B.n936 B.n45 163.367
R1183 B.n936 B.n47 163.367
R1184 B.n932 B.n47 163.367
R1185 B.n932 B.n52 163.367
R1186 B.n928 B.n52 163.367
R1187 B.n928 B.n54 163.367
R1188 B.n924 B.n54 163.367
R1189 B.n924 B.n59 163.367
R1190 B.n920 B.n59 163.367
R1191 B.n920 B.n61 163.367
R1192 B.n916 B.n61 163.367
R1193 B.n916 B.n66 163.367
R1194 B.n912 B.n66 163.367
R1195 B.n912 B.n68 163.367
R1196 B.n908 B.n68 163.367
R1197 B.n908 B.n73 163.367
R1198 B.n904 B.n73 163.367
R1199 B.n904 B.n75 163.367
R1200 B.n900 B.n75 163.367
R1201 B.n900 B.n80 163.367
R1202 B.n896 B.n80 163.367
R1203 B.n896 B.n82 163.367
R1204 B.n892 B.n82 163.367
R1205 B.n892 B.n87 163.367
R1206 B.n888 B.n87 163.367
R1207 B.n888 B.n89 163.367
R1208 B.n884 B.n89 163.367
R1209 B.n884 B.n94 163.367
R1210 B.n880 B.n94 163.367
R1211 B.n880 B.n96 163.367
R1212 B.n876 B.n96 163.367
R1213 B.n876 B.n100 163.367
R1214 B.n872 B.n100 163.367
R1215 B.n872 B.n102 163.367
R1216 B.n868 B.n102 163.367
R1217 B.n868 B.n108 163.367
R1218 B.n864 B.n108 163.367
R1219 B.n864 B.n110 163.367
R1220 B.n860 B.n110 163.367
R1221 B.n860 B.n115 163.367
R1222 B.n152 B.t20 145.71
R1223 B.n445 B.t18 145.71
R1224 B.n155 B.t14 145.702
R1225 B.n442 B.t11 145.702
R1226 B.n577 B.n405 116.416
R1227 B.n854 B.n114 116.416
R1228 B.n156 B.n155 73.3096
R1229 B.n153 B.n152 73.3096
R1230 B.n446 B.n445 73.3096
R1231 B.n443 B.n442 73.3096
R1232 B.n153 B.t21 72.4011
R1233 B.n446 B.t17 72.4011
R1234 B.n156 B.t15 72.3924
R1235 B.n443 B.t10 72.3924
R1236 B.n856 B.n855 71.676
R1237 B.n157 B.n118 71.676
R1238 B.n161 B.n119 71.676
R1239 B.n165 B.n120 71.676
R1240 B.n169 B.n121 71.676
R1241 B.n173 B.n122 71.676
R1242 B.n177 B.n123 71.676
R1243 B.n181 B.n124 71.676
R1244 B.n185 B.n125 71.676
R1245 B.n189 B.n126 71.676
R1246 B.n193 B.n127 71.676
R1247 B.n197 B.n128 71.676
R1248 B.n201 B.n129 71.676
R1249 B.n205 B.n130 71.676
R1250 B.n209 B.n131 71.676
R1251 B.n214 B.n132 71.676
R1252 B.n218 B.n133 71.676
R1253 B.n222 B.n134 71.676
R1254 B.n226 B.n135 71.676
R1255 B.n230 B.n136 71.676
R1256 B.n234 B.n137 71.676
R1257 B.n238 B.n138 71.676
R1258 B.n242 B.n139 71.676
R1259 B.n246 B.n140 71.676
R1260 B.n250 B.n141 71.676
R1261 B.n254 B.n142 71.676
R1262 B.n258 B.n143 71.676
R1263 B.n262 B.n144 71.676
R1264 B.n266 B.n145 71.676
R1265 B.n270 B.n146 71.676
R1266 B.n274 B.n147 71.676
R1267 B.n278 B.n148 71.676
R1268 B.n282 B.n149 71.676
R1269 B.n150 B.n149 71.676
R1270 B.n281 B.n148 71.676
R1271 B.n277 B.n147 71.676
R1272 B.n273 B.n146 71.676
R1273 B.n269 B.n145 71.676
R1274 B.n265 B.n144 71.676
R1275 B.n261 B.n143 71.676
R1276 B.n257 B.n142 71.676
R1277 B.n253 B.n141 71.676
R1278 B.n249 B.n140 71.676
R1279 B.n245 B.n139 71.676
R1280 B.n241 B.n138 71.676
R1281 B.n237 B.n137 71.676
R1282 B.n233 B.n136 71.676
R1283 B.n229 B.n135 71.676
R1284 B.n225 B.n134 71.676
R1285 B.n221 B.n133 71.676
R1286 B.n217 B.n132 71.676
R1287 B.n213 B.n131 71.676
R1288 B.n208 B.n130 71.676
R1289 B.n204 B.n129 71.676
R1290 B.n200 B.n128 71.676
R1291 B.n196 B.n127 71.676
R1292 B.n192 B.n126 71.676
R1293 B.n188 B.n125 71.676
R1294 B.n184 B.n124 71.676
R1295 B.n180 B.n123 71.676
R1296 B.n176 B.n122 71.676
R1297 B.n172 B.n121 71.676
R1298 B.n168 B.n120 71.676
R1299 B.n164 B.n119 71.676
R1300 B.n160 B.n118 71.676
R1301 B.n855 B.n117 71.676
R1302 B.n579 B.n578 71.676
R1303 B.n441 B.n409 71.676
R1304 B.n571 B.n410 71.676
R1305 B.n567 B.n411 71.676
R1306 B.n563 B.n412 71.676
R1307 B.n559 B.n413 71.676
R1308 B.n555 B.n414 71.676
R1309 B.n551 B.n415 71.676
R1310 B.n547 B.n416 71.676
R1311 B.n543 B.n417 71.676
R1312 B.n539 B.n418 71.676
R1313 B.n535 B.n419 71.676
R1314 B.n531 B.n420 71.676
R1315 B.n527 B.n421 71.676
R1316 B.n523 B.n422 71.676
R1317 B.n519 B.n423 71.676
R1318 B.n515 B.n424 71.676
R1319 B.n511 B.n425 71.676
R1320 B.n507 B.n426 71.676
R1321 B.n502 B.n427 71.676
R1322 B.n498 B.n428 71.676
R1323 B.n494 B.n429 71.676
R1324 B.n490 B.n430 71.676
R1325 B.n486 B.n431 71.676
R1326 B.n482 B.n432 71.676
R1327 B.n478 B.n433 71.676
R1328 B.n474 B.n434 71.676
R1329 B.n470 B.n435 71.676
R1330 B.n466 B.n436 71.676
R1331 B.n462 B.n437 71.676
R1332 B.n458 B.n438 71.676
R1333 B.n454 B.n439 71.676
R1334 B.n450 B.n440 71.676
R1335 B.n578 B.n408 71.676
R1336 B.n572 B.n409 71.676
R1337 B.n568 B.n410 71.676
R1338 B.n564 B.n411 71.676
R1339 B.n560 B.n412 71.676
R1340 B.n556 B.n413 71.676
R1341 B.n552 B.n414 71.676
R1342 B.n548 B.n415 71.676
R1343 B.n544 B.n416 71.676
R1344 B.n540 B.n417 71.676
R1345 B.n536 B.n418 71.676
R1346 B.n532 B.n419 71.676
R1347 B.n528 B.n420 71.676
R1348 B.n524 B.n421 71.676
R1349 B.n520 B.n422 71.676
R1350 B.n516 B.n423 71.676
R1351 B.n512 B.n424 71.676
R1352 B.n508 B.n425 71.676
R1353 B.n503 B.n426 71.676
R1354 B.n499 B.n427 71.676
R1355 B.n495 B.n428 71.676
R1356 B.n491 B.n429 71.676
R1357 B.n487 B.n430 71.676
R1358 B.n483 B.n431 71.676
R1359 B.n479 B.n432 71.676
R1360 B.n475 B.n433 71.676
R1361 B.n471 B.n434 71.676
R1362 B.n467 B.n435 71.676
R1363 B.n463 B.n436 71.676
R1364 B.n459 B.n437 71.676
R1365 B.n455 B.n438 71.676
R1366 B.n451 B.n439 71.676
R1367 B.n447 B.n440 71.676
R1368 B.n986 B.n985 71.676
R1369 B.n986 B.n2 71.676
R1370 B.n211 B.n156 59.5399
R1371 B.n154 B.n153 59.5399
R1372 B.n505 B.n446 59.5399
R1373 B.n444 B.n443 59.5399
R1374 B.n584 B.n405 57.7834
R1375 B.n584 B.n401 57.7834
R1376 B.n590 B.n401 57.7834
R1377 B.n590 B.n397 57.7834
R1378 B.n596 B.n397 57.7834
R1379 B.n596 B.n393 57.7834
R1380 B.n603 B.n393 57.7834
R1381 B.n603 B.n602 57.7834
R1382 B.n609 B.n386 57.7834
R1383 B.n615 B.n386 57.7834
R1384 B.n615 B.n382 57.7834
R1385 B.n621 B.n382 57.7834
R1386 B.n621 B.n378 57.7834
R1387 B.n627 B.n378 57.7834
R1388 B.n627 B.n374 57.7834
R1389 B.n633 B.n374 57.7834
R1390 B.n633 B.n370 57.7834
R1391 B.n639 B.n370 57.7834
R1392 B.n639 B.n365 57.7834
R1393 B.n645 B.n365 57.7834
R1394 B.n645 B.n366 57.7834
R1395 B.n651 B.n358 57.7834
R1396 B.n657 B.n358 57.7834
R1397 B.n657 B.n354 57.7834
R1398 B.n663 B.n354 57.7834
R1399 B.n663 B.n350 57.7834
R1400 B.n669 B.n350 57.7834
R1401 B.n669 B.n346 57.7834
R1402 B.n675 B.n346 57.7834
R1403 B.n675 B.n341 57.7834
R1404 B.n681 B.n341 57.7834
R1405 B.n681 B.n342 57.7834
R1406 B.n687 B.n334 57.7834
R1407 B.n693 B.n334 57.7834
R1408 B.n693 B.n330 57.7834
R1409 B.n699 B.n330 57.7834
R1410 B.n699 B.n326 57.7834
R1411 B.n705 B.n326 57.7834
R1412 B.n705 B.n322 57.7834
R1413 B.n711 B.n322 57.7834
R1414 B.n711 B.n318 57.7834
R1415 B.n717 B.n318 57.7834
R1416 B.n723 B.n314 57.7834
R1417 B.n723 B.n310 57.7834
R1418 B.n729 B.n310 57.7834
R1419 B.n729 B.n306 57.7834
R1420 B.n735 B.n306 57.7834
R1421 B.n735 B.n302 57.7834
R1422 B.n741 B.n302 57.7834
R1423 B.n741 B.n298 57.7834
R1424 B.n748 B.n298 57.7834
R1425 B.n748 B.n747 57.7834
R1426 B.n754 B.n291 57.7834
R1427 B.n761 B.n291 57.7834
R1428 B.n761 B.n287 57.7834
R1429 B.n767 B.n287 57.7834
R1430 B.n767 B.n4 57.7834
R1431 B.n984 B.n4 57.7834
R1432 B.n984 B.n983 57.7834
R1433 B.n983 B.n982 57.7834
R1434 B.n982 B.n8 57.7834
R1435 B.n12 B.n8 57.7834
R1436 B.n975 B.n12 57.7834
R1437 B.n975 B.n974 57.7834
R1438 B.n974 B.n973 57.7834
R1439 B.n967 B.n19 57.7834
R1440 B.n967 B.n966 57.7834
R1441 B.n966 B.n965 57.7834
R1442 B.n965 B.n23 57.7834
R1443 B.n959 B.n23 57.7834
R1444 B.n959 B.n958 57.7834
R1445 B.n958 B.n957 57.7834
R1446 B.n957 B.n30 57.7834
R1447 B.n951 B.n30 57.7834
R1448 B.n951 B.n950 57.7834
R1449 B.n949 B.n37 57.7834
R1450 B.n943 B.n37 57.7834
R1451 B.n943 B.n942 57.7834
R1452 B.n942 B.n941 57.7834
R1453 B.n941 B.n44 57.7834
R1454 B.n935 B.n44 57.7834
R1455 B.n935 B.n934 57.7834
R1456 B.n934 B.n933 57.7834
R1457 B.n933 B.n51 57.7834
R1458 B.n927 B.n51 57.7834
R1459 B.n926 B.n925 57.7834
R1460 B.n925 B.n58 57.7834
R1461 B.n919 B.n58 57.7834
R1462 B.n919 B.n918 57.7834
R1463 B.n918 B.n917 57.7834
R1464 B.n917 B.n65 57.7834
R1465 B.n911 B.n65 57.7834
R1466 B.n911 B.n910 57.7834
R1467 B.n910 B.n909 57.7834
R1468 B.n909 B.n72 57.7834
R1469 B.n903 B.n72 57.7834
R1470 B.n902 B.n901 57.7834
R1471 B.n901 B.n79 57.7834
R1472 B.n895 B.n79 57.7834
R1473 B.n895 B.n894 57.7834
R1474 B.n894 B.n893 57.7834
R1475 B.n893 B.n86 57.7834
R1476 B.n887 B.n86 57.7834
R1477 B.n887 B.n886 57.7834
R1478 B.n886 B.n885 57.7834
R1479 B.n885 B.n93 57.7834
R1480 B.n879 B.n93 57.7834
R1481 B.n879 B.n878 57.7834
R1482 B.n878 B.n877 57.7834
R1483 B.n871 B.n103 57.7834
R1484 B.n871 B.n870 57.7834
R1485 B.n870 B.n869 57.7834
R1486 B.n869 B.n107 57.7834
R1487 B.n863 B.n107 57.7834
R1488 B.n863 B.n862 57.7834
R1489 B.n862 B.n861 57.7834
R1490 B.n861 B.n114 57.7834
R1491 B.n366 B.t5 56.9337
R1492 B.t0 B.n902 56.9337
R1493 B.n687 B.t2 51.8352
R1494 B.n927 B.t6 51.8352
R1495 B.t3 B.n314 45.0372
R1496 B.n950 B.t1 45.0372
R1497 B.n602 B.t9 38.2392
R1498 B.n754 B.t7 38.2392
R1499 B.n973 B.t4 38.2392
R1500 B.n103 B.t13 38.2392
R1501 B.n581 B.n580 36.3712
R1502 B.n448 B.n403 36.3712
R1503 B.n852 B.n851 36.3712
R1504 B.n858 B.n857 36.3712
R1505 B.n609 B.t9 19.5447
R1506 B.n747 B.t7 19.5447
R1507 B.n19 B.t4 19.5447
R1508 B.n877 B.t13 19.5447
R1509 B B.n987 18.0485
R1510 B.n717 B.t3 12.7467
R1511 B.t1 B.n949 12.7467
R1512 B.n582 B.n581 10.6151
R1513 B.n582 B.n399 10.6151
R1514 B.n592 B.n399 10.6151
R1515 B.n593 B.n592 10.6151
R1516 B.n594 B.n593 10.6151
R1517 B.n594 B.n391 10.6151
R1518 B.n605 B.n391 10.6151
R1519 B.n606 B.n605 10.6151
R1520 B.n607 B.n606 10.6151
R1521 B.n607 B.n384 10.6151
R1522 B.n617 B.n384 10.6151
R1523 B.n618 B.n617 10.6151
R1524 B.n619 B.n618 10.6151
R1525 B.n619 B.n376 10.6151
R1526 B.n629 B.n376 10.6151
R1527 B.n630 B.n629 10.6151
R1528 B.n631 B.n630 10.6151
R1529 B.n631 B.n368 10.6151
R1530 B.n641 B.n368 10.6151
R1531 B.n642 B.n641 10.6151
R1532 B.n643 B.n642 10.6151
R1533 B.n643 B.n360 10.6151
R1534 B.n653 B.n360 10.6151
R1535 B.n654 B.n653 10.6151
R1536 B.n655 B.n654 10.6151
R1537 B.n655 B.n352 10.6151
R1538 B.n665 B.n352 10.6151
R1539 B.n666 B.n665 10.6151
R1540 B.n667 B.n666 10.6151
R1541 B.n667 B.n344 10.6151
R1542 B.n677 B.n344 10.6151
R1543 B.n678 B.n677 10.6151
R1544 B.n679 B.n678 10.6151
R1545 B.n679 B.n336 10.6151
R1546 B.n689 B.n336 10.6151
R1547 B.n690 B.n689 10.6151
R1548 B.n691 B.n690 10.6151
R1549 B.n691 B.n328 10.6151
R1550 B.n701 B.n328 10.6151
R1551 B.n702 B.n701 10.6151
R1552 B.n703 B.n702 10.6151
R1553 B.n703 B.n320 10.6151
R1554 B.n713 B.n320 10.6151
R1555 B.n714 B.n713 10.6151
R1556 B.n715 B.n714 10.6151
R1557 B.n715 B.n312 10.6151
R1558 B.n725 B.n312 10.6151
R1559 B.n726 B.n725 10.6151
R1560 B.n727 B.n726 10.6151
R1561 B.n727 B.n304 10.6151
R1562 B.n737 B.n304 10.6151
R1563 B.n738 B.n737 10.6151
R1564 B.n739 B.n738 10.6151
R1565 B.n739 B.n296 10.6151
R1566 B.n750 B.n296 10.6151
R1567 B.n751 B.n750 10.6151
R1568 B.n752 B.n751 10.6151
R1569 B.n752 B.n289 10.6151
R1570 B.n763 B.n289 10.6151
R1571 B.n764 B.n763 10.6151
R1572 B.n765 B.n764 10.6151
R1573 B.n765 B.n0 10.6151
R1574 B.n580 B.n407 10.6151
R1575 B.n575 B.n407 10.6151
R1576 B.n575 B.n574 10.6151
R1577 B.n574 B.n573 10.6151
R1578 B.n573 B.n570 10.6151
R1579 B.n570 B.n569 10.6151
R1580 B.n569 B.n566 10.6151
R1581 B.n566 B.n565 10.6151
R1582 B.n565 B.n562 10.6151
R1583 B.n562 B.n561 10.6151
R1584 B.n561 B.n558 10.6151
R1585 B.n558 B.n557 10.6151
R1586 B.n557 B.n554 10.6151
R1587 B.n554 B.n553 10.6151
R1588 B.n553 B.n550 10.6151
R1589 B.n550 B.n549 10.6151
R1590 B.n549 B.n546 10.6151
R1591 B.n546 B.n545 10.6151
R1592 B.n545 B.n542 10.6151
R1593 B.n542 B.n541 10.6151
R1594 B.n541 B.n538 10.6151
R1595 B.n538 B.n537 10.6151
R1596 B.n537 B.n534 10.6151
R1597 B.n534 B.n533 10.6151
R1598 B.n533 B.n530 10.6151
R1599 B.n530 B.n529 10.6151
R1600 B.n529 B.n526 10.6151
R1601 B.n526 B.n525 10.6151
R1602 B.n522 B.n521 10.6151
R1603 B.n521 B.n518 10.6151
R1604 B.n518 B.n517 10.6151
R1605 B.n517 B.n514 10.6151
R1606 B.n514 B.n513 10.6151
R1607 B.n513 B.n510 10.6151
R1608 B.n510 B.n509 10.6151
R1609 B.n509 B.n506 10.6151
R1610 B.n504 B.n501 10.6151
R1611 B.n501 B.n500 10.6151
R1612 B.n500 B.n497 10.6151
R1613 B.n497 B.n496 10.6151
R1614 B.n496 B.n493 10.6151
R1615 B.n493 B.n492 10.6151
R1616 B.n492 B.n489 10.6151
R1617 B.n489 B.n488 10.6151
R1618 B.n488 B.n485 10.6151
R1619 B.n485 B.n484 10.6151
R1620 B.n484 B.n481 10.6151
R1621 B.n481 B.n480 10.6151
R1622 B.n480 B.n477 10.6151
R1623 B.n477 B.n476 10.6151
R1624 B.n476 B.n473 10.6151
R1625 B.n473 B.n472 10.6151
R1626 B.n472 B.n469 10.6151
R1627 B.n469 B.n468 10.6151
R1628 B.n468 B.n465 10.6151
R1629 B.n465 B.n464 10.6151
R1630 B.n464 B.n461 10.6151
R1631 B.n461 B.n460 10.6151
R1632 B.n460 B.n457 10.6151
R1633 B.n457 B.n456 10.6151
R1634 B.n456 B.n453 10.6151
R1635 B.n453 B.n452 10.6151
R1636 B.n452 B.n449 10.6151
R1637 B.n449 B.n448 10.6151
R1638 B.n586 B.n403 10.6151
R1639 B.n587 B.n586 10.6151
R1640 B.n588 B.n587 10.6151
R1641 B.n588 B.n395 10.6151
R1642 B.n598 B.n395 10.6151
R1643 B.n599 B.n598 10.6151
R1644 B.n600 B.n599 10.6151
R1645 B.n600 B.n388 10.6151
R1646 B.n611 B.n388 10.6151
R1647 B.n612 B.n611 10.6151
R1648 B.n613 B.n612 10.6151
R1649 B.n613 B.n380 10.6151
R1650 B.n623 B.n380 10.6151
R1651 B.n624 B.n623 10.6151
R1652 B.n625 B.n624 10.6151
R1653 B.n625 B.n372 10.6151
R1654 B.n635 B.n372 10.6151
R1655 B.n636 B.n635 10.6151
R1656 B.n637 B.n636 10.6151
R1657 B.n637 B.n363 10.6151
R1658 B.n647 B.n363 10.6151
R1659 B.n648 B.n647 10.6151
R1660 B.n649 B.n648 10.6151
R1661 B.n649 B.n356 10.6151
R1662 B.n659 B.n356 10.6151
R1663 B.n660 B.n659 10.6151
R1664 B.n661 B.n660 10.6151
R1665 B.n661 B.n348 10.6151
R1666 B.n671 B.n348 10.6151
R1667 B.n672 B.n671 10.6151
R1668 B.n673 B.n672 10.6151
R1669 B.n673 B.n339 10.6151
R1670 B.n683 B.n339 10.6151
R1671 B.n684 B.n683 10.6151
R1672 B.n685 B.n684 10.6151
R1673 B.n685 B.n332 10.6151
R1674 B.n695 B.n332 10.6151
R1675 B.n696 B.n695 10.6151
R1676 B.n697 B.n696 10.6151
R1677 B.n697 B.n324 10.6151
R1678 B.n707 B.n324 10.6151
R1679 B.n708 B.n707 10.6151
R1680 B.n709 B.n708 10.6151
R1681 B.n709 B.n316 10.6151
R1682 B.n719 B.n316 10.6151
R1683 B.n720 B.n719 10.6151
R1684 B.n721 B.n720 10.6151
R1685 B.n721 B.n308 10.6151
R1686 B.n731 B.n308 10.6151
R1687 B.n732 B.n731 10.6151
R1688 B.n733 B.n732 10.6151
R1689 B.n733 B.n300 10.6151
R1690 B.n743 B.n300 10.6151
R1691 B.n744 B.n743 10.6151
R1692 B.n745 B.n744 10.6151
R1693 B.n745 B.n293 10.6151
R1694 B.n756 B.n293 10.6151
R1695 B.n757 B.n756 10.6151
R1696 B.n759 B.n757 10.6151
R1697 B.n759 B.n758 10.6151
R1698 B.n758 B.n285 10.6151
R1699 B.n770 B.n285 10.6151
R1700 B.n771 B.n770 10.6151
R1701 B.n772 B.n771 10.6151
R1702 B.n773 B.n772 10.6151
R1703 B.n774 B.n773 10.6151
R1704 B.n777 B.n774 10.6151
R1705 B.n778 B.n777 10.6151
R1706 B.n779 B.n778 10.6151
R1707 B.n780 B.n779 10.6151
R1708 B.n782 B.n780 10.6151
R1709 B.n783 B.n782 10.6151
R1710 B.n784 B.n783 10.6151
R1711 B.n785 B.n784 10.6151
R1712 B.n787 B.n785 10.6151
R1713 B.n788 B.n787 10.6151
R1714 B.n789 B.n788 10.6151
R1715 B.n790 B.n789 10.6151
R1716 B.n792 B.n790 10.6151
R1717 B.n793 B.n792 10.6151
R1718 B.n794 B.n793 10.6151
R1719 B.n795 B.n794 10.6151
R1720 B.n797 B.n795 10.6151
R1721 B.n798 B.n797 10.6151
R1722 B.n799 B.n798 10.6151
R1723 B.n800 B.n799 10.6151
R1724 B.n802 B.n800 10.6151
R1725 B.n803 B.n802 10.6151
R1726 B.n804 B.n803 10.6151
R1727 B.n805 B.n804 10.6151
R1728 B.n807 B.n805 10.6151
R1729 B.n808 B.n807 10.6151
R1730 B.n809 B.n808 10.6151
R1731 B.n810 B.n809 10.6151
R1732 B.n812 B.n810 10.6151
R1733 B.n813 B.n812 10.6151
R1734 B.n814 B.n813 10.6151
R1735 B.n815 B.n814 10.6151
R1736 B.n817 B.n815 10.6151
R1737 B.n818 B.n817 10.6151
R1738 B.n819 B.n818 10.6151
R1739 B.n820 B.n819 10.6151
R1740 B.n822 B.n820 10.6151
R1741 B.n823 B.n822 10.6151
R1742 B.n824 B.n823 10.6151
R1743 B.n825 B.n824 10.6151
R1744 B.n827 B.n825 10.6151
R1745 B.n828 B.n827 10.6151
R1746 B.n829 B.n828 10.6151
R1747 B.n830 B.n829 10.6151
R1748 B.n832 B.n830 10.6151
R1749 B.n833 B.n832 10.6151
R1750 B.n834 B.n833 10.6151
R1751 B.n835 B.n834 10.6151
R1752 B.n837 B.n835 10.6151
R1753 B.n838 B.n837 10.6151
R1754 B.n839 B.n838 10.6151
R1755 B.n840 B.n839 10.6151
R1756 B.n842 B.n840 10.6151
R1757 B.n843 B.n842 10.6151
R1758 B.n844 B.n843 10.6151
R1759 B.n845 B.n844 10.6151
R1760 B.n847 B.n845 10.6151
R1761 B.n848 B.n847 10.6151
R1762 B.n849 B.n848 10.6151
R1763 B.n850 B.n849 10.6151
R1764 B.n851 B.n850 10.6151
R1765 B.n979 B.n1 10.6151
R1766 B.n979 B.n978 10.6151
R1767 B.n978 B.n977 10.6151
R1768 B.n977 B.n10 10.6151
R1769 B.n971 B.n10 10.6151
R1770 B.n971 B.n970 10.6151
R1771 B.n970 B.n969 10.6151
R1772 B.n969 B.n17 10.6151
R1773 B.n963 B.n17 10.6151
R1774 B.n963 B.n962 10.6151
R1775 B.n962 B.n961 10.6151
R1776 B.n961 B.n25 10.6151
R1777 B.n955 B.n25 10.6151
R1778 B.n955 B.n954 10.6151
R1779 B.n954 B.n953 10.6151
R1780 B.n953 B.n32 10.6151
R1781 B.n947 B.n32 10.6151
R1782 B.n947 B.n946 10.6151
R1783 B.n946 B.n945 10.6151
R1784 B.n945 B.n39 10.6151
R1785 B.n939 B.n39 10.6151
R1786 B.n939 B.n938 10.6151
R1787 B.n938 B.n937 10.6151
R1788 B.n937 B.n46 10.6151
R1789 B.n931 B.n46 10.6151
R1790 B.n931 B.n930 10.6151
R1791 B.n930 B.n929 10.6151
R1792 B.n929 B.n53 10.6151
R1793 B.n923 B.n53 10.6151
R1794 B.n923 B.n922 10.6151
R1795 B.n922 B.n921 10.6151
R1796 B.n921 B.n60 10.6151
R1797 B.n915 B.n60 10.6151
R1798 B.n915 B.n914 10.6151
R1799 B.n914 B.n913 10.6151
R1800 B.n913 B.n67 10.6151
R1801 B.n907 B.n67 10.6151
R1802 B.n907 B.n906 10.6151
R1803 B.n906 B.n905 10.6151
R1804 B.n905 B.n74 10.6151
R1805 B.n899 B.n74 10.6151
R1806 B.n899 B.n898 10.6151
R1807 B.n898 B.n897 10.6151
R1808 B.n897 B.n81 10.6151
R1809 B.n891 B.n81 10.6151
R1810 B.n891 B.n890 10.6151
R1811 B.n890 B.n889 10.6151
R1812 B.n889 B.n88 10.6151
R1813 B.n883 B.n88 10.6151
R1814 B.n883 B.n882 10.6151
R1815 B.n882 B.n881 10.6151
R1816 B.n881 B.n95 10.6151
R1817 B.n875 B.n95 10.6151
R1818 B.n875 B.n874 10.6151
R1819 B.n874 B.n873 10.6151
R1820 B.n873 B.n101 10.6151
R1821 B.n867 B.n101 10.6151
R1822 B.n867 B.n866 10.6151
R1823 B.n866 B.n865 10.6151
R1824 B.n865 B.n109 10.6151
R1825 B.n859 B.n109 10.6151
R1826 B.n859 B.n858 10.6151
R1827 B.n857 B.n116 10.6151
R1828 B.n158 B.n116 10.6151
R1829 B.n159 B.n158 10.6151
R1830 B.n162 B.n159 10.6151
R1831 B.n163 B.n162 10.6151
R1832 B.n166 B.n163 10.6151
R1833 B.n167 B.n166 10.6151
R1834 B.n170 B.n167 10.6151
R1835 B.n171 B.n170 10.6151
R1836 B.n174 B.n171 10.6151
R1837 B.n175 B.n174 10.6151
R1838 B.n178 B.n175 10.6151
R1839 B.n179 B.n178 10.6151
R1840 B.n182 B.n179 10.6151
R1841 B.n183 B.n182 10.6151
R1842 B.n186 B.n183 10.6151
R1843 B.n187 B.n186 10.6151
R1844 B.n190 B.n187 10.6151
R1845 B.n191 B.n190 10.6151
R1846 B.n194 B.n191 10.6151
R1847 B.n195 B.n194 10.6151
R1848 B.n198 B.n195 10.6151
R1849 B.n199 B.n198 10.6151
R1850 B.n202 B.n199 10.6151
R1851 B.n203 B.n202 10.6151
R1852 B.n206 B.n203 10.6151
R1853 B.n207 B.n206 10.6151
R1854 B.n210 B.n207 10.6151
R1855 B.n215 B.n212 10.6151
R1856 B.n216 B.n215 10.6151
R1857 B.n219 B.n216 10.6151
R1858 B.n220 B.n219 10.6151
R1859 B.n223 B.n220 10.6151
R1860 B.n224 B.n223 10.6151
R1861 B.n227 B.n224 10.6151
R1862 B.n228 B.n227 10.6151
R1863 B.n232 B.n231 10.6151
R1864 B.n235 B.n232 10.6151
R1865 B.n236 B.n235 10.6151
R1866 B.n239 B.n236 10.6151
R1867 B.n240 B.n239 10.6151
R1868 B.n243 B.n240 10.6151
R1869 B.n244 B.n243 10.6151
R1870 B.n247 B.n244 10.6151
R1871 B.n248 B.n247 10.6151
R1872 B.n251 B.n248 10.6151
R1873 B.n252 B.n251 10.6151
R1874 B.n255 B.n252 10.6151
R1875 B.n256 B.n255 10.6151
R1876 B.n259 B.n256 10.6151
R1877 B.n260 B.n259 10.6151
R1878 B.n263 B.n260 10.6151
R1879 B.n264 B.n263 10.6151
R1880 B.n267 B.n264 10.6151
R1881 B.n268 B.n267 10.6151
R1882 B.n271 B.n268 10.6151
R1883 B.n272 B.n271 10.6151
R1884 B.n275 B.n272 10.6151
R1885 B.n276 B.n275 10.6151
R1886 B.n279 B.n276 10.6151
R1887 B.n280 B.n279 10.6151
R1888 B.n283 B.n280 10.6151
R1889 B.n284 B.n283 10.6151
R1890 B.n852 B.n284 10.6151
R1891 B.n987 B.n0 8.11757
R1892 B.n987 B.n1 8.11757
R1893 B.n522 B.n444 6.5566
R1894 B.n506 B.n505 6.5566
R1895 B.n212 B.n211 6.5566
R1896 B.n228 B.n154 6.5566
R1897 B.n342 B.t2 5.94874
R1898 B.t6 B.n926 5.94874
R1899 B.n525 B.n444 4.05904
R1900 B.n505 B.n504 4.05904
R1901 B.n211 B.n210 4.05904
R1902 B.n231 B.n154 4.05904
R1903 B.n651 B.t5 0.850249
R1904 B.n903 B.t0 0.850249
R1905 VN.n68 VN.n67 161.3
R1906 VN.n66 VN.n36 161.3
R1907 VN.n65 VN.n64 161.3
R1908 VN.n63 VN.n37 161.3
R1909 VN.n62 VN.n61 161.3
R1910 VN.n60 VN.n38 161.3
R1911 VN.n59 VN.n58 161.3
R1912 VN.n57 VN.n39 161.3
R1913 VN.n56 VN.n55 161.3
R1914 VN.n54 VN.n40 161.3
R1915 VN.n53 VN.n52 161.3
R1916 VN.n51 VN.n42 161.3
R1917 VN.n50 VN.n49 161.3
R1918 VN.n48 VN.n43 161.3
R1919 VN.n47 VN.n46 161.3
R1920 VN.n33 VN.n32 161.3
R1921 VN.n31 VN.n1 161.3
R1922 VN.n30 VN.n29 161.3
R1923 VN.n28 VN.n2 161.3
R1924 VN.n27 VN.n26 161.3
R1925 VN.n25 VN.n3 161.3
R1926 VN.n24 VN.n23 161.3
R1927 VN.n22 VN.n4 161.3
R1928 VN.n21 VN.n20 161.3
R1929 VN.n18 VN.n5 161.3
R1930 VN.n17 VN.n16 161.3
R1931 VN.n15 VN.n6 161.3
R1932 VN.n14 VN.n13 161.3
R1933 VN.n12 VN.n7 161.3
R1934 VN.n11 VN.n10 161.3
R1935 VN.n45 VN.t3 86.6913
R1936 VN.n9 VN.t7 86.6913
R1937 VN.n34 VN.n0 81.7486
R1938 VN.n69 VN.n35 81.7486
R1939 VN.n26 VN.n2 56.5193
R1940 VN.n61 VN.n37 56.5193
R1941 VN.n45 VN.n44 55.4655
R1942 VN.n9 VN.n8 55.4655
R1943 VN.n8 VN.t2 53.5793
R1944 VN.n19 VN.t4 53.5793
R1945 VN.n0 VN.t5 53.5793
R1946 VN.n44 VN.t0 53.5793
R1947 VN.n41 VN.t1 53.5793
R1948 VN.n35 VN.t6 53.5793
R1949 VN VN.n69 51.8086
R1950 VN.n13 VN.n6 40.4934
R1951 VN.n17 VN.n6 40.4934
R1952 VN.n49 VN.n42 40.4934
R1953 VN.n53 VN.n42 40.4934
R1954 VN.n12 VN.n11 24.4675
R1955 VN.n13 VN.n12 24.4675
R1956 VN.n18 VN.n17 24.4675
R1957 VN.n20 VN.n18 24.4675
R1958 VN.n24 VN.n4 24.4675
R1959 VN.n25 VN.n24 24.4675
R1960 VN.n26 VN.n25 24.4675
R1961 VN.n30 VN.n2 24.4675
R1962 VN.n31 VN.n30 24.4675
R1963 VN.n32 VN.n31 24.4675
R1964 VN.n49 VN.n48 24.4675
R1965 VN.n48 VN.n47 24.4675
R1966 VN.n61 VN.n60 24.4675
R1967 VN.n60 VN.n59 24.4675
R1968 VN.n59 VN.n39 24.4675
R1969 VN.n55 VN.n54 24.4675
R1970 VN.n54 VN.n53 24.4675
R1971 VN.n67 VN.n66 24.4675
R1972 VN.n66 VN.n65 24.4675
R1973 VN.n65 VN.n37 24.4675
R1974 VN.n11 VN.n8 19.0848
R1975 VN.n20 VN.n19 19.0848
R1976 VN.n47 VN.n44 19.0848
R1977 VN.n55 VN.n41 19.0848
R1978 VN.n32 VN.n0 8.31928
R1979 VN.n67 VN.n35 8.31928
R1980 VN.n19 VN.n4 5.38324
R1981 VN.n41 VN.n39 5.38324
R1982 VN.n10 VN.n9 3.21184
R1983 VN.n46 VN.n45 3.21184
R1984 VN.n69 VN.n68 0.354971
R1985 VN.n34 VN.n33 0.354971
R1986 VN VN.n34 0.26696
R1987 VN.n68 VN.n36 0.189894
R1988 VN.n64 VN.n36 0.189894
R1989 VN.n64 VN.n63 0.189894
R1990 VN.n63 VN.n62 0.189894
R1991 VN.n62 VN.n38 0.189894
R1992 VN.n58 VN.n38 0.189894
R1993 VN.n58 VN.n57 0.189894
R1994 VN.n57 VN.n56 0.189894
R1995 VN.n56 VN.n40 0.189894
R1996 VN.n52 VN.n40 0.189894
R1997 VN.n52 VN.n51 0.189894
R1998 VN.n51 VN.n50 0.189894
R1999 VN.n50 VN.n43 0.189894
R2000 VN.n46 VN.n43 0.189894
R2001 VN.n10 VN.n7 0.189894
R2002 VN.n14 VN.n7 0.189894
R2003 VN.n15 VN.n14 0.189894
R2004 VN.n16 VN.n15 0.189894
R2005 VN.n16 VN.n5 0.189894
R2006 VN.n21 VN.n5 0.189894
R2007 VN.n22 VN.n21 0.189894
R2008 VN.n23 VN.n22 0.189894
R2009 VN.n23 VN.n3 0.189894
R2010 VN.n27 VN.n3 0.189894
R2011 VN.n28 VN.n27 0.189894
R2012 VN.n29 VN.n28 0.189894
R2013 VN.n29 VN.n1 0.189894
R2014 VN.n33 VN.n1 0.189894
R2015 VDD2.n2 VDD2.n1 70.3257
R2016 VDD2.n2 VDD2.n0 70.3257
R2017 VDD2 VDD2.n5 70.3228
R2018 VDD2.n4 VDD2.n3 68.7519
R2019 VDD2.n4 VDD2.n2 44.9912
R2020 VDD2.n5 VDD2.t7 2.58199
R2021 VDD2.n5 VDD2.t4 2.58199
R2022 VDD2.n3 VDD2.t1 2.58199
R2023 VDD2.n3 VDD2.t6 2.58199
R2024 VDD2.n1 VDD2.t3 2.58199
R2025 VDD2.n1 VDD2.t2 2.58199
R2026 VDD2.n0 VDD2.t0 2.58199
R2027 VDD2.n0 VDD2.t5 2.58199
R2028 VDD2 VDD2.n4 1.688
C0 VDD2 VDD1 2.21862f
C1 VTAIL VDD1 7.14461f
C2 VP VDD1 6.4529f
C3 VN VDD1 0.1534f
C4 VDD2 VTAIL 7.20473f
C5 VP VDD2 0.610255f
C6 VDD2 VN 5.99787f
C7 VP VTAIL 6.90475f
C8 VTAIL VN 6.89065f
C9 VP VN 7.90326f
C10 VDD2 B 5.952732f
C11 VDD1 B 6.487932f
C12 VTAIL B 8.447101f
C13 VN B 18.48483f
C14 VP B 17.14646f
C15 VDD2.t0 B 0.170067f
C16 VDD2.t5 B 0.170067f
C17 VDD2.n0 B 1.48399f
C18 VDD2.t3 B 0.170067f
C19 VDD2.t2 B 0.170067f
C20 VDD2.n1 B 1.48399f
C21 VDD2.n2 B 3.90986f
C22 VDD2.t1 B 0.170067f
C23 VDD2.t6 B 0.170067f
C24 VDD2.n3 B 1.46901f
C25 VDD2.n4 B 3.26042f
C26 VDD2.t7 B 0.170067f
C27 VDD2.t4 B 0.170067f
C28 VDD2.n5 B 1.48395f
C29 VN.t5 B 1.41627f
C30 VN.n0 B 0.586008f
C31 VN.n1 B 0.019966f
C32 VN.n2 B 0.027477f
C33 VN.n3 B 0.019966f
C34 VN.n4 B 0.022882f
C35 VN.n5 B 0.019966f
C36 VN.n6 B 0.01614f
C37 VN.n7 B 0.019966f
C38 VN.t2 B 1.41627f
C39 VN.n8 B 0.585747f
C40 VN.t7 B 1.66817f
C41 VN.n9 B 0.554418f
C42 VN.n10 B 0.246062f
C43 VN.n11 B 0.03317f
C44 VN.n12 B 0.037211f
C45 VN.n13 B 0.039682f
C46 VN.n14 B 0.019966f
C47 VN.n15 B 0.019966f
C48 VN.n16 B 0.019966f
C49 VN.n17 B 0.039682f
C50 VN.n18 B 0.037211f
C51 VN.t4 B 1.41627f
C52 VN.n19 B 0.511911f
C53 VN.n20 B 0.03317f
C54 VN.n21 B 0.019966f
C55 VN.n22 B 0.019966f
C56 VN.n23 B 0.019966f
C57 VN.n24 B 0.037211f
C58 VN.n25 B 0.037211f
C59 VN.n26 B 0.030816f
C60 VN.n27 B 0.019966f
C61 VN.n28 B 0.019966f
C62 VN.n29 B 0.019966f
C63 VN.n30 B 0.037211f
C64 VN.n31 B 0.037211f
C65 VN.n32 B 0.025086f
C66 VN.n33 B 0.032224f
C67 VN.n34 B 0.054284f
C68 VN.t6 B 1.41627f
C69 VN.n35 B 0.586008f
C70 VN.n36 B 0.019966f
C71 VN.n37 B 0.027477f
C72 VN.n38 B 0.019966f
C73 VN.n39 B 0.022882f
C74 VN.n40 B 0.019966f
C75 VN.t1 B 1.41627f
C76 VN.n41 B 0.511911f
C77 VN.n42 B 0.01614f
C78 VN.n43 B 0.019966f
C79 VN.t0 B 1.41627f
C80 VN.n44 B 0.585747f
C81 VN.t3 B 1.66817f
C82 VN.n45 B 0.554418f
C83 VN.n46 B 0.246062f
C84 VN.n47 B 0.03317f
C85 VN.n48 B 0.037211f
C86 VN.n49 B 0.039682f
C87 VN.n50 B 0.019966f
C88 VN.n51 B 0.019966f
C89 VN.n52 B 0.019966f
C90 VN.n53 B 0.039682f
C91 VN.n54 B 0.037211f
C92 VN.n55 B 0.03317f
C93 VN.n56 B 0.019966f
C94 VN.n57 B 0.019966f
C95 VN.n58 B 0.019966f
C96 VN.n59 B 0.037211f
C97 VN.n60 B 0.037211f
C98 VN.n61 B 0.030816f
C99 VN.n62 B 0.019966f
C100 VN.n63 B 0.019966f
C101 VN.n64 B 0.019966f
C102 VN.n65 B 0.037211f
C103 VN.n66 B 0.037211f
C104 VN.n67 B 0.025086f
C105 VN.n68 B 0.032224f
C106 VN.n69 B 1.20282f
C107 VTAIL.t1 B 0.137061f
C108 VTAIL.t6 B 0.137061f
C109 VTAIL.n0 B 1.12834f
C110 VTAIL.n1 B 0.444298f
C111 VTAIL.t4 B 1.43766f
C112 VTAIL.n2 B 0.53877f
C113 VTAIL.t14 B 1.43766f
C114 VTAIL.n3 B 0.53877f
C115 VTAIL.t9 B 0.137061f
C116 VTAIL.t11 B 0.137061f
C117 VTAIL.n4 B 1.12834f
C118 VTAIL.n5 B 0.677498f
C119 VTAIL.t15 B 1.43766f
C120 VTAIL.n6 B 1.53094f
C121 VTAIL.t5 B 1.43767f
C122 VTAIL.n7 B 1.53094f
C123 VTAIL.t2 B 0.137061f
C124 VTAIL.t3 B 0.137061f
C125 VTAIL.n8 B 1.12834f
C126 VTAIL.n9 B 0.677495f
C127 VTAIL.t7 B 1.43767f
C128 VTAIL.n10 B 0.538767f
C129 VTAIL.t10 B 1.43767f
C130 VTAIL.n11 B 0.538767f
C131 VTAIL.t13 B 0.137061f
C132 VTAIL.t8 B 0.137061f
C133 VTAIL.n12 B 1.12834f
C134 VTAIL.n13 B 0.677495f
C135 VTAIL.t12 B 1.43766f
C136 VTAIL.n14 B 1.53094f
C137 VTAIL.t0 B 1.43766f
C138 VTAIL.n15 B 1.5267f
C139 VDD1.t5 B 0.173318f
C140 VDD1.t6 B 0.173318f
C141 VDD1.n0 B 1.51367f
C142 VDD1.t0 B 0.173318f
C143 VDD1.t1 B 0.173318f
C144 VDD1.n1 B 1.51235f
C145 VDD1.t3 B 0.173318f
C146 VDD1.t7 B 0.173318f
C147 VDD1.n2 B 1.51235f
C148 VDD1.n3 B 4.04379f
C149 VDD1.t4 B 0.173318f
C150 VDD1.t2 B 0.173318f
C151 VDD1.n4 B 1.49709f
C152 VDD1.n5 B 3.35845f
C153 VP.t1 B 1.45228f
C154 VP.n0 B 0.600905f
C155 VP.n1 B 0.020473f
C156 VP.n2 B 0.028176f
C157 VP.n3 B 0.020473f
C158 VP.n4 B 0.023463f
C159 VP.n5 B 0.020473f
C160 VP.n6 B 0.016551f
C161 VP.n7 B 0.020473f
C162 VP.t6 B 1.45228f
C163 VP.n8 B 0.524924f
C164 VP.n9 B 0.020473f
C165 VP.n10 B 0.031599f
C166 VP.n11 B 0.020473f
C167 VP.n12 B 0.025724f
C168 VP.t3 B 1.45228f
C169 VP.n13 B 0.600905f
C170 VP.n14 B 0.020473f
C171 VP.n15 B 0.028176f
C172 VP.n16 B 0.020473f
C173 VP.n17 B 0.023463f
C174 VP.n18 B 0.020473f
C175 VP.n19 B 0.016551f
C176 VP.n20 B 0.020473f
C177 VP.t2 B 1.45228f
C178 VP.n21 B 0.600638f
C179 VP.t5 B 1.71058f
C180 VP.n22 B 0.568513f
C181 VP.n23 B 0.252318f
C182 VP.n24 B 0.034013f
C183 VP.n25 B 0.038157f
C184 VP.n26 B 0.040691f
C185 VP.n27 B 0.020473f
C186 VP.n28 B 0.020473f
C187 VP.n29 B 0.020473f
C188 VP.n30 B 0.040691f
C189 VP.n31 B 0.038157f
C190 VP.t7 B 1.45228f
C191 VP.n32 B 0.524924f
C192 VP.n33 B 0.034013f
C193 VP.n34 B 0.020473f
C194 VP.n35 B 0.020473f
C195 VP.n36 B 0.020473f
C196 VP.n37 B 0.038157f
C197 VP.n38 B 0.038157f
C198 VP.n39 B 0.031599f
C199 VP.n40 B 0.020473f
C200 VP.n41 B 0.020473f
C201 VP.n42 B 0.020473f
C202 VP.n43 B 0.038157f
C203 VP.n44 B 0.038157f
C204 VP.n45 B 0.025724f
C205 VP.n46 B 0.033044f
C206 VP.n47 B 1.22511f
C207 VP.t0 B 1.45228f
C208 VP.n48 B 0.600905f
C209 VP.n49 B 1.23936f
C210 VP.n50 B 0.033044f
C211 VP.n51 B 0.020473f
C212 VP.n52 B 0.038157f
C213 VP.n53 B 0.038157f
C214 VP.n54 B 0.028176f
C215 VP.n55 B 0.020473f
C216 VP.n56 B 0.020473f
C217 VP.n57 B 0.020473f
C218 VP.n58 B 0.038157f
C219 VP.n59 B 0.038157f
C220 VP.n60 B 0.023463f
C221 VP.n61 B 0.020473f
C222 VP.n62 B 0.020473f
C223 VP.n63 B 0.034013f
C224 VP.n64 B 0.038157f
C225 VP.n65 B 0.040691f
C226 VP.n66 B 0.020473f
C227 VP.n67 B 0.020473f
C228 VP.n68 B 0.020473f
C229 VP.n69 B 0.040691f
C230 VP.n70 B 0.038157f
C231 VP.t4 B 1.45228f
C232 VP.n71 B 0.524924f
C233 VP.n72 B 0.034013f
C234 VP.n73 B 0.020473f
C235 VP.n74 B 0.020473f
C236 VP.n75 B 0.020473f
C237 VP.n76 B 0.038157f
C238 VP.n77 B 0.038157f
C239 VP.n78 B 0.031599f
C240 VP.n79 B 0.020473f
C241 VP.n80 B 0.020473f
C242 VP.n81 B 0.020473f
C243 VP.n82 B 0.038157f
C244 VP.n83 B 0.038157f
C245 VP.n84 B 0.025724f
C246 VP.n85 B 0.033044f
C247 VP.n86 B 0.055664f
.ends

