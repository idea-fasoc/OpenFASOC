* NGSPICE file created from diff_pair_sample_0896.ext - technology: sky130A

.subckt diff_pair_sample_0896 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 w_n1974_n3928# sky130_fd_pr__pfet_01v8 ad=5.772 pd=30.38 as=5.772 ps=30.38 w=14.8 l=2.18
X1 B.t11 B.t9 B.t10 w_n1974_n3928# sky130_fd_pr__pfet_01v8 ad=5.772 pd=30.38 as=0 ps=0 w=14.8 l=2.18
X2 VDD1.t0 VP.t1 VTAIL.t3 w_n1974_n3928# sky130_fd_pr__pfet_01v8 ad=5.772 pd=30.38 as=5.772 ps=30.38 w=14.8 l=2.18
X3 VDD2.t1 VN.t0 VTAIL.t1 w_n1974_n3928# sky130_fd_pr__pfet_01v8 ad=5.772 pd=30.38 as=5.772 ps=30.38 w=14.8 l=2.18
X4 VDD2.t0 VN.t1 VTAIL.t0 w_n1974_n3928# sky130_fd_pr__pfet_01v8 ad=5.772 pd=30.38 as=5.772 ps=30.38 w=14.8 l=2.18
X5 B.t8 B.t6 B.t7 w_n1974_n3928# sky130_fd_pr__pfet_01v8 ad=5.772 pd=30.38 as=0 ps=0 w=14.8 l=2.18
X6 B.t5 B.t3 B.t4 w_n1974_n3928# sky130_fd_pr__pfet_01v8 ad=5.772 pd=30.38 as=0 ps=0 w=14.8 l=2.18
X7 B.t2 B.t0 B.t1 w_n1974_n3928# sky130_fd_pr__pfet_01v8 ad=5.772 pd=30.38 as=0 ps=0 w=14.8 l=2.18
R0 VP.n0 VP.t1 258.495
R1 VP.n0 VP.t0 212.831
R2 VP VP.n0 0.336784
R3 VTAIL.n322 VTAIL.n246 756.745
R4 VTAIL.n76 VTAIL.n0 756.745
R5 VTAIL.n240 VTAIL.n164 756.745
R6 VTAIL.n158 VTAIL.n82 756.745
R7 VTAIL.n273 VTAIL.n272 585
R8 VTAIL.n270 VTAIL.n269 585
R9 VTAIL.n279 VTAIL.n278 585
R10 VTAIL.n281 VTAIL.n280 585
R11 VTAIL.n266 VTAIL.n265 585
R12 VTAIL.n287 VTAIL.n286 585
R13 VTAIL.n289 VTAIL.n288 585
R14 VTAIL.n262 VTAIL.n261 585
R15 VTAIL.n295 VTAIL.n294 585
R16 VTAIL.n297 VTAIL.n296 585
R17 VTAIL.n258 VTAIL.n257 585
R18 VTAIL.n303 VTAIL.n302 585
R19 VTAIL.n305 VTAIL.n304 585
R20 VTAIL.n254 VTAIL.n253 585
R21 VTAIL.n311 VTAIL.n310 585
R22 VTAIL.n314 VTAIL.n313 585
R23 VTAIL.n312 VTAIL.n250 585
R24 VTAIL.n319 VTAIL.n249 585
R25 VTAIL.n321 VTAIL.n320 585
R26 VTAIL.n323 VTAIL.n322 585
R27 VTAIL.n27 VTAIL.n26 585
R28 VTAIL.n24 VTAIL.n23 585
R29 VTAIL.n33 VTAIL.n32 585
R30 VTAIL.n35 VTAIL.n34 585
R31 VTAIL.n20 VTAIL.n19 585
R32 VTAIL.n41 VTAIL.n40 585
R33 VTAIL.n43 VTAIL.n42 585
R34 VTAIL.n16 VTAIL.n15 585
R35 VTAIL.n49 VTAIL.n48 585
R36 VTAIL.n51 VTAIL.n50 585
R37 VTAIL.n12 VTAIL.n11 585
R38 VTAIL.n57 VTAIL.n56 585
R39 VTAIL.n59 VTAIL.n58 585
R40 VTAIL.n8 VTAIL.n7 585
R41 VTAIL.n65 VTAIL.n64 585
R42 VTAIL.n68 VTAIL.n67 585
R43 VTAIL.n66 VTAIL.n4 585
R44 VTAIL.n73 VTAIL.n3 585
R45 VTAIL.n75 VTAIL.n74 585
R46 VTAIL.n77 VTAIL.n76 585
R47 VTAIL.n241 VTAIL.n240 585
R48 VTAIL.n239 VTAIL.n238 585
R49 VTAIL.n237 VTAIL.n167 585
R50 VTAIL.n171 VTAIL.n168 585
R51 VTAIL.n232 VTAIL.n231 585
R52 VTAIL.n230 VTAIL.n229 585
R53 VTAIL.n173 VTAIL.n172 585
R54 VTAIL.n224 VTAIL.n223 585
R55 VTAIL.n222 VTAIL.n221 585
R56 VTAIL.n177 VTAIL.n176 585
R57 VTAIL.n216 VTAIL.n215 585
R58 VTAIL.n214 VTAIL.n213 585
R59 VTAIL.n181 VTAIL.n180 585
R60 VTAIL.n208 VTAIL.n207 585
R61 VTAIL.n206 VTAIL.n205 585
R62 VTAIL.n185 VTAIL.n184 585
R63 VTAIL.n200 VTAIL.n199 585
R64 VTAIL.n198 VTAIL.n197 585
R65 VTAIL.n189 VTAIL.n188 585
R66 VTAIL.n192 VTAIL.n191 585
R67 VTAIL.n159 VTAIL.n158 585
R68 VTAIL.n157 VTAIL.n156 585
R69 VTAIL.n155 VTAIL.n85 585
R70 VTAIL.n89 VTAIL.n86 585
R71 VTAIL.n150 VTAIL.n149 585
R72 VTAIL.n148 VTAIL.n147 585
R73 VTAIL.n91 VTAIL.n90 585
R74 VTAIL.n142 VTAIL.n141 585
R75 VTAIL.n140 VTAIL.n139 585
R76 VTAIL.n95 VTAIL.n94 585
R77 VTAIL.n134 VTAIL.n133 585
R78 VTAIL.n132 VTAIL.n131 585
R79 VTAIL.n99 VTAIL.n98 585
R80 VTAIL.n126 VTAIL.n125 585
R81 VTAIL.n124 VTAIL.n123 585
R82 VTAIL.n103 VTAIL.n102 585
R83 VTAIL.n118 VTAIL.n117 585
R84 VTAIL.n116 VTAIL.n115 585
R85 VTAIL.n107 VTAIL.n106 585
R86 VTAIL.n110 VTAIL.n109 585
R87 VTAIL.t3 VTAIL.n190 327.466
R88 VTAIL.t1 VTAIL.n108 327.466
R89 VTAIL.t0 VTAIL.n271 327.466
R90 VTAIL.t2 VTAIL.n25 327.466
R91 VTAIL.n272 VTAIL.n269 171.744
R92 VTAIL.n279 VTAIL.n269 171.744
R93 VTAIL.n280 VTAIL.n279 171.744
R94 VTAIL.n280 VTAIL.n265 171.744
R95 VTAIL.n287 VTAIL.n265 171.744
R96 VTAIL.n288 VTAIL.n287 171.744
R97 VTAIL.n288 VTAIL.n261 171.744
R98 VTAIL.n295 VTAIL.n261 171.744
R99 VTAIL.n296 VTAIL.n295 171.744
R100 VTAIL.n296 VTAIL.n257 171.744
R101 VTAIL.n303 VTAIL.n257 171.744
R102 VTAIL.n304 VTAIL.n303 171.744
R103 VTAIL.n304 VTAIL.n253 171.744
R104 VTAIL.n311 VTAIL.n253 171.744
R105 VTAIL.n313 VTAIL.n311 171.744
R106 VTAIL.n313 VTAIL.n312 171.744
R107 VTAIL.n312 VTAIL.n249 171.744
R108 VTAIL.n321 VTAIL.n249 171.744
R109 VTAIL.n322 VTAIL.n321 171.744
R110 VTAIL.n26 VTAIL.n23 171.744
R111 VTAIL.n33 VTAIL.n23 171.744
R112 VTAIL.n34 VTAIL.n33 171.744
R113 VTAIL.n34 VTAIL.n19 171.744
R114 VTAIL.n41 VTAIL.n19 171.744
R115 VTAIL.n42 VTAIL.n41 171.744
R116 VTAIL.n42 VTAIL.n15 171.744
R117 VTAIL.n49 VTAIL.n15 171.744
R118 VTAIL.n50 VTAIL.n49 171.744
R119 VTAIL.n50 VTAIL.n11 171.744
R120 VTAIL.n57 VTAIL.n11 171.744
R121 VTAIL.n58 VTAIL.n57 171.744
R122 VTAIL.n58 VTAIL.n7 171.744
R123 VTAIL.n65 VTAIL.n7 171.744
R124 VTAIL.n67 VTAIL.n65 171.744
R125 VTAIL.n67 VTAIL.n66 171.744
R126 VTAIL.n66 VTAIL.n3 171.744
R127 VTAIL.n75 VTAIL.n3 171.744
R128 VTAIL.n76 VTAIL.n75 171.744
R129 VTAIL.n240 VTAIL.n239 171.744
R130 VTAIL.n239 VTAIL.n167 171.744
R131 VTAIL.n171 VTAIL.n167 171.744
R132 VTAIL.n231 VTAIL.n171 171.744
R133 VTAIL.n231 VTAIL.n230 171.744
R134 VTAIL.n230 VTAIL.n172 171.744
R135 VTAIL.n223 VTAIL.n172 171.744
R136 VTAIL.n223 VTAIL.n222 171.744
R137 VTAIL.n222 VTAIL.n176 171.744
R138 VTAIL.n215 VTAIL.n176 171.744
R139 VTAIL.n215 VTAIL.n214 171.744
R140 VTAIL.n214 VTAIL.n180 171.744
R141 VTAIL.n207 VTAIL.n180 171.744
R142 VTAIL.n207 VTAIL.n206 171.744
R143 VTAIL.n206 VTAIL.n184 171.744
R144 VTAIL.n199 VTAIL.n184 171.744
R145 VTAIL.n199 VTAIL.n198 171.744
R146 VTAIL.n198 VTAIL.n188 171.744
R147 VTAIL.n191 VTAIL.n188 171.744
R148 VTAIL.n158 VTAIL.n157 171.744
R149 VTAIL.n157 VTAIL.n85 171.744
R150 VTAIL.n89 VTAIL.n85 171.744
R151 VTAIL.n149 VTAIL.n89 171.744
R152 VTAIL.n149 VTAIL.n148 171.744
R153 VTAIL.n148 VTAIL.n90 171.744
R154 VTAIL.n141 VTAIL.n90 171.744
R155 VTAIL.n141 VTAIL.n140 171.744
R156 VTAIL.n140 VTAIL.n94 171.744
R157 VTAIL.n133 VTAIL.n94 171.744
R158 VTAIL.n133 VTAIL.n132 171.744
R159 VTAIL.n132 VTAIL.n98 171.744
R160 VTAIL.n125 VTAIL.n98 171.744
R161 VTAIL.n125 VTAIL.n124 171.744
R162 VTAIL.n124 VTAIL.n102 171.744
R163 VTAIL.n117 VTAIL.n102 171.744
R164 VTAIL.n117 VTAIL.n116 171.744
R165 VTAIL.n116 VTAIL.n106 171.744
R166 VTAIL.n109 VTAIL.n106 171.744
R167 VTAIL.n272 VTAIL.t0 85.8723
R168 VTAIL.n26 VTAIL.t2 85.8723
R169 VTAIL.n191 VTAIL.t3 85.8723
R170 VTAIL.n109 VTAIL.t1 85.8723
R171 VTAIL.n327 VTAIL.n326 35.2884
R172 VTAIL.n81 VTAIL.n80 35.2884
R173 VTAIL.n245 VTAIL.n244 35.2884
R174 VTAIL.n163 VTAIL.n162 35.2884
R175 VTAIL.n163 VTAIL.n81 29.4531
R176 VTAIL.n327 VTAIL.n245 27.2893
R177 VTAIL.n273 VTAIL.n271 16.3895
R178 VTAIL.n27 VTAIL.n25 16.3895
R179 VTAIL.n192 VTAIL.n190 16.3895
R180 VTAIL.n110 VTAIL.n108 16.3895
R181 VTAIL.n320 VTAIL.n319 13.1884
R182 VTAIL.n74 VTAIL.n73 13.1884
R183 VTAIL.n238 VTAIL.n237 13.1884
R184 VTAIL.n156 VTAIL.n155 13.1884
R185 VTAIL.n274 VTAIL.n270 12.8005
R186 VTAIL.n318 VTAIL.n250 12.8005
R187 VTAIL.n323 VTAIL.n248 12.8005
R188 VTAIL.n28 VTAIL.n24 12.8005
R189 VTAIL.n72 VTAIL.n4 12.8005
R190 VTAIL.n77 VTAIL.n2 12.8005
R191 VTAIL.n241 VTAIL.n166 12.8005
R192 VTAIL.n236 VTAIL.n168 12.8005
R193 VTAIL.n193 VTAIL.n189 12.8005
R194 VTAIL.n159 VTAIL.n84 12.8005
R195 VTAIL.n154 VTAIL.n86 12.8005
R196 VTAIL.n111 VTAIL.n107 12.8005
R197 VTAIL.n278 VTAIL.n277 12.0247
R198 VTAIL.n315 VTAIL.n314 12.0247
R199 VTAIL.n324 VTAIL.n246 12.0247
R200 VTAIL.n32 VTAIL.n31 12.0247
R201 VTAIL.n69 VTAIL.n68 12.0247
R202 VTAIL.n78 VTAIL.n0 12.0247
R203 VTAIL.n242 VTAIL.n164 12.0247
R204 VTAIL.n233 VTAIL.n232 12.0247
R205 VTAIL.n197 VTAIL.n196 12.0247
R206 VTAIL.n160 VTAIL.n82 12.0247
R207 VTAIL.n151 VTAIL.n150 12.0247
R208 VTAIL.n115 VTAIL.n114 12.0247
R209 VTAIL.n281 VTAIL.n268 11.249
R210 VTAIL.n310 VTAIL.n252 11.249
R211 VTAIL.n35 VTAIL.n22 11.249
R212 VTAIL.n64 VTAIL.n6 11.249
R213 VTAIL.n229 VTAIL.n170 11.249
R214 VTAIL.n200 VTAIL.n187 11.249
R215 VTAIL.n147 VTAIL.n88 11.249
R216 VTAIL.n118 VTAIL.n105 11.249
R217 VTAIL.n282 VTAIL.n266 10.4732
R218 VTAIL.n309 VTAIL.n254 10.4732
R219 VTAIL.n36 VTAIL.n20 10.4732
R220 VTAIL.n63 VTAIL.n8 10.4732
R221 VTAIL.n228 VTAIL.n173 10.4732
R222 VTAIL.n201 VTAIL.n185 10.4732
R223 VTAIL.n146 VTAIL.n91 10.4732
R224 VTAIL.n119 VTAIL.n103 10.4732
R225 VTAIL.n286 VTAIL.n285 9.69747
R226 VTAIL.n306 VTAIL.n305 9.69747
R227 VTAIL.n40 VTAIL.n39 9.69747
R228 VTAIL.n60 VTAIL.n59 9.69747
R229 VTAIL.n225 VTAIL.n224 9.69747
R230 VTAIL.n205 VTAIL.n204 9.69747
R231 VTAIL.n143 VTAIL.n142 9.69747
R232 VTAIL.n123 VTAIL.n122 9.69747
R233 VTAIL.n326 VTAIL.n325 9.45567
R234 VTAIL.n80 VTAIL.n79 9.45567
R235 VTAIL.n244 VTAIL.n243 9.45567
R236 VTAIL.n162 VTAIL.n161 9.45567
R237 VTAIL.n325 VTAIL.n324 9.3005
R238 VTAIL.n248 VTAIL.n247 9.3005
R239 VTAIL.n293 VTAIL.n292 9.3005
R240 VTAIL.n291 VTAIL.n290 9.3005
R241 VTAIL.n264 VTAIL.n263 9.3005
R242 VTAIL.n285 VTAIL.n284 9.3005
R243 VTAIL.n283 VTAIL.n282 9.3005
R244 VTAIL.n268 VTAIL.n267 9.3005
R245 VTAIL.n277 VTAIL.n276 9.3005
R246 VTAIL.n275 VTAIL.n274 9.3005
R247 VTAIL.n260 VTAIL.n259 9.3005
R248 VTAIL.n299 VTAIL.n298 9.3005
R249 VTAIL.n301 VTAIL.n300 9.3005
R250 VTAIL.n256 VTAIL.n255 9.3005
R251 VTAIL.n307 VTAIL.n306 9.3005
R252 VTAIL.n309 VTAIL.n308 9.3005
R253 VTAIL.n252 VTAIL.n251 9.3005
R254 VTAIL.n316 VTAIL.n315 9.3005
R255 VTAIL.n318 VTAIL.n317 9.3005
R256 VTAIL.n79 VTAIL.n78 9.3005
R257 VTAIL.n2 VTAIL.n1 9.3005
R258 VTAIL.n47 VTAIL.n46 9.3005
R259 VTAIL.n45 VTAIL.n44 9.3005
R260 VTAIL.n18 VTAIL.n17 9.3005
R261 VTAIL.n39 VTAIL.n38 9.3005
R262 VTAIL.n37 VTAIL.n36 9.3005
R263 VTAIL.n22 VTAIL.n21 9.3005
R264 VTAIL.n31 VTAIL.n30 9.3005
R265 VTAIL.n29 VTAIL.n28 9.3005
R266 VTAIL.n14 VTAIL.n13 9.3005
R267 VTAIL.n53 VTAIL.n52 9.3005
R268 VTAIL.n55 VTAIL.n54 9.3005
R269 VTAIL.n10 VTAIL.n9 9.3005
R270 VTAIL.n61 VTAIL.n60 9.3005
R271 VTAIL.n63 VTAIL.n62 9.3005
R272 VTAIL.n6 VTAIL.n5 9.3005
R273 VTAIL.n70 VTAIL.n69 9.3005
R274 VTAIL.n72 VTAIL.n71 9.3005
R275 VTAIL.n218 VTAIL.n217 9.3005
R276 VTAIL.n220 VTAIL.n219 9.3005
R277 VTAIL.n175 VTAIL.n174 9.3005
R278 VTAIL.n226 VTAIL.n225 9.3005
R279 VTAIL.n228 VTAIL.n227 9.3005
R280 VTAIL.n170 VTAIL.n169 9.3005
R281 VTAIL.n234 VTAIL.n233 9.3005
R282 VTAIL.n236 VTAIL.n235 9.3005
R283 VTAIL.n243 VTAIL.n242 9.3005
R284 VTAIL.n166 VTAIL.n165 9.3005
R285 VTAIL.n179 VTAIL.n178 9.3005
R286 VTAIL.n212 VTAIL.n211 9.3005
R287 VTAIL.n210 VTAIL.n209 9.3005
R288 VTAIL.n183 VTAIL.n182 9.3005
R289 VTAIL.n204 VTAIL.n203 9.3005
R290 VTAIL.n202 VTAIL.n201 9.3005
R291 VTAIL.n187 VTAIL.n186 9.3005
R292 VTAIL.n196 VTAIL.n195 9.3005
R293 VTAIL.n194 VTAIL.n193 9.3005
R294 VTAIL.n136 VTAIL.n135 9.3005
R295 VTAIL.n138 VTAIL.n137 9.3005
R296 VTAIL.n93 VTAIL.n92 9.3005
R297 VTAIL.n144 VTAIL.n143 9.3005
R298 VTAIL.n146 VTAIL.n145 9.3005
R299 VTAIL.n88 VTAIL.n87 9.3005
R300 VTAIL.n152 VTAIL.n151 9.3005
R301 VTAIL.n154 VTAIL.n153 9.3005
R302 VTAIL.n161 VTAIL.n160 9.3005
R303 VTAIL.n84 VTAIL.n83 9.3005
R304 VTAIL.n97 VTAIL.n96 9.3005
R305 VTAIL.n130 VTAIL.n129 9.3005
R306 VTAIL.n128 VTAIL.n127 9.3005
R307 VTAIL.n101 VTAIL.n100 9.3005
R308 VTAIL.n122 VTAIL.n121 9.3005
R309 VTAIL.n120 VTAIL.n119 9.3005
R310 VTAIL.n105 VTAIL.n104 9.3005
R311 VTAIL.n114 VTAIL.n113 9.3005
R312 VTAIL.n112 VTAIL.n111 9.3005
R313 VTAIL.n289 VTAIL.n264 8.92171
R314 VTAIL.n302 VTAIL.n256 8.92171
R315 VTAIL.n43 VTAIL.n18 8.92171
R316 VTAIL.n56 VTAIL.n10 8.92171
R317 VTAIL.n221 VTAIL.n175 8.92171
R318 VTAIL.n208 VTAIL.n183 8.92171
R319 VTAIL.n139 VTAIL.n93 8.92171
R320 VTAIL.n126 VTAIL.n101 8.92171
R321 VTAIL.n290 VTAIL.n262 8.14595
R322 VTAIL.n301 VTAIL.n258 8.14595
R323 VTAIL.n44 VTAIL.n16 8.14595
R324 VTAIL.n55 VTAIL.n12 8.14595
R325 VTAIL.n220 VTAIL.n177 8.14595
R326 VTAIL.n209 VTAIL.n181 8.14595
R327 VTAIL.n138 VTAIL.n95 8.14595
R328 VTAIL.n127 VTAIL.n99 8.14595
R329 VTAIL.n294 VTAIL.n293 7.3702
R330 VTAIL.n298 VTAIL.n297 7.3702
R331 VTAIL.n48 VTAIL.n47 7.3702
R332 VTAIL.n52 VTAIL.n51 7.3702
R333 VTAIL.n217 VTAIL.n216 7.3702
R334 VTAIL.n213 VTAIL.n212 7.3702
R335 VTAIL.n135 VTAIL.n134 7.3702
R336 VTAIL.n131 VTAIL.n130 7.3702
R337 VTAIL.n294 VTAIL.n260 6.59444
R338 VTAIL.n297 VTAIL.n260 6.59444
R339 VTAIL.n48 VTAIL.n14 6.59444
R340 VTAIL.n51 VTAIL.n14 6.59444
R341 VTAIL.n216 VTAIL.n179 6.59444
R342 VTAIL.n213 VTAIL.n179 6.59444
R343 VTAIL.n134 VTAIL.n97 6.59444
R344 VTAIL.n131 VTAIL.n97 6.59444
R345 VTAIL.n293 VTAIL.n262 5.81868
R346 VTAIL.n298 VTAIL.n258 5.81868
R347 VTAIL.n47 VTAIL.n16 5.81868
R348 VTAIL.n52 VTAIL.n12 5.81868
R349 VTAIL.n217 VTAIL.n177 5.81868
R350 VTAIL.n212 VTAIL.n181 5.81868
R351 VTAIL.n135 VTAIL.n95 5.81868
R352 VTAIL.n130 VTAIL.n99 5.81868
R353 VTAIL.n290 VTAIL.n289 5.04292
R354 VTAIL.n302 VTAIL.n301 5.04292
R355 VTAIL.n44 VTAIL.n43 5.04292
R356 VTAIL.n56 VTAIL.n55 5.04292
R357 VTAIL.n221 VTAIL.n220 5.04292
R358 VTAIL.n209 VTAIL.n208 5.04292
R359 VTAIL.n139 VTAIL.n138 5.04292
R360 VTAIL.n127 VTAIL.n126 5.04292
R361 VTAIL.n286 VTAIL.n264 4.26717
R362 VTAIL.n305 VTAIL.n256 4.26717
R363 VTAIL.n40 VTAIL.n18 4.26717
R364 VTAIL.n59 VTAIL.n10 4.26717
R365 VTAIL.n224 VTAIL.n175 4.26717
R366 VTAIL.n205 VTAIL.n183 4.26717
R367 VTAIL.n142 VTAIL.n93 4.26717
R368 VTAIL.n123 VTAIL.n101 4.26717
R369 VTAIL.n275 VTAIL.n271 3.70982
R370 VTAIL.n29 VTAIL.n25 3.70982
R371 VTAIL.n194 VTAIL.n190 3.70982
R372 VTAIL.n112 VTAIL.n108 3.70982
R373 VTAIL.n285 VTAIL.n266 3.49141
R374 VTAIL.n306 VTAIL.n254 3.49141
R375 VTAIL.n39 VTAIL.n20 3.49141
R376 VTAIL.n60 VTAIL.n8 3.49141
R377 VTAIL.n225 VTAIL.n173 3.49141
R378 VTAIL.n204 VTAIL.n185 3.49141
R379 VTAIL.n143 VTAIL.n91 3.49141
R380 VTAIL.n122 VTAIL.n103 3.49141
R381 VTAIL.n282 VTAIL.n281 2.71565
R382 VTAIL.n310 VTAIL.n309 2.71565
R383 VTAIL.n36 VTAIL.n35 2.71565
R384 VTAIL.n64 VTAIL.n63 2.71565
R385 VTAIL.n229 VTAIL.n228 2.71565
R386 VTAIL.n201 VTAIL.n200 2.71565
R387 VTAIL.n147 VTAIL.n146 2.71565
R388 VTAIL.n119 VTAIL.n118 2.71565
R389 VTAIL.n278 VTAIL.n268 1.93989
R390 VTAIL.n314 VTAIL.n252 1.93989
R391 VTAIL.n326 VTAIL.n246 1.93989
R392 VTAIL.n32 VTAIL.n22 1.93989
R393 VTAIL.n68 VTAIL.n6 1.93989
R394 VTAIL.n80 VTAIL.n0 1.93989
R395 VTAIL.n244 VTAIL.n164 1.93989
R396 VTAIL.n232 VTAIL.n170 1.93989
R397 VTAIL.n197 VTAIL.n187 1.93989
R398 VTAIL.n162 VTAIL.n82 1.93989
R399 VTAIL.n150 VTAIL.n88 1.93989
R400 VTAIL.n115 VTAIL.n105 1.93989
R401 VTAIL.n245 VTAIL.n163 1.55222
R402 VTAIL.n277 VTAIL.n270 1.16414
R403 VTAIL.n315 VTAIL.n250 1.16414
R404 VTAIL.n324 VTAIL.n323 1.16414
R405 VTAIL.n31 VTAIL.n24 1.16414
R406 VTAIL.n69 VTAIL.n4 1.16414
R407 VTAIL.n78 VTAIL.n77 1.16414
R408 VTAIL.n242 VTAIL.n241 1.16414
R409 VTAIL.n233 VTAIL.n168 1.16414
R410 VTAIL.n196 VTAIL.n189 1.16414
R411 VTAIL.n160 VTAIL.n159 1.16414
R412 VTAIL.n151 VTAIL.n86 1.16414
R413 VTAIL.n114 VTAIL.n107 1.16414
R414 VTAIL VTAIL.n81 1.06947
R415 VTAIL VTAIL.n327 0.483259
R416 VTAIL.n274 VTAIL.n273 0.388379
R417 VTAIL.n319 VTAIL.n318 0.388379
R418 VTAIL.n320 VTAIL.n248 0.388379
R419 VTAIL.n28 VTAIL.n27 0.388379
R420 VTAIL.n73 VTAIL.n72 0.388379
R421 VTAIL.n74 VTAIL.n2 0.388379
R422 VTAIL.n238 VTAIL.n166 0.388379
R423 VTAIL.n237 VTAIL.n236 0.388379
R424 VTAIL.n193 VTAIL.n192 0.388379
R425 VTAIL.n156 VTAIL.n84 0.388379
R426 VTAIL.n155 VTAIL.n154 0.388379
R427 VTAIL.n111 VTAIL.n110 0.388379
R428 VTAIL.n276 VTAIL.n275 0.155672
R429 VTAIL.n276 VTAIL.n267 0.155672
R430 VTAIL.n283 VTAIL.n267 0.155672
R431 VTAIL.n284 VTAIL.n283 0.155672
R432 VTAIL.n284 VTAIL.n263 0.155672
R433 VTAIL.n291 VTAIL.n263 0.155672
R434 VTAIL.n292 VTAIL.n291 0.155672
R435 VTAIL.n292 VTAIL.n259 0.155672
R436 VTAIL.n299 VTAIL.n259 0.155672
R437 VTAIL.n300 VTAIL.n299 0.155672
R438 VTAIL.n300 VTAIL.n255 0.155672
R439 VTAIL.n307 VTAIL.n255 0.155672
R440 VTAIL.n308 VTAIL.n307 0.155672
R441 VTAIL.n308 VTAIL.n251 0.155672
R442 VTAIL.n316 VTAIL.n251 0.155672
R443 VTAIL.n317 VTAIL.n316 0.155672
R444 VTAIL.n317 VTAIL.n247 0.155672
R445 VTAIL.n325 VTAIL.n247 0.155672
R446 VTAIL.n30 VTAIL.n29 0.155672
R447 VTAIL.n30 VTAIL.n21 0.155672
R448 VTAIL.n37 VTAIL.n21 0.155672
R449 VTAIL.n38 VTAIL.n37 0.155672
R450 VTAIL.n38 VTAIL.n17 0.155672
R451 VTAIL.n45 VTAIL.n17 0.155672
R452 VTAIL.n46 VTAIL.n45 0.155672
R453 VTAIL.n46 VTAIL.n13 0.155672
R454 VTAIL.n53 VTAIL.n13 0.155672
R455 VTAIL.n54 VTAIL.n53 0.155672
R456 VTAIL.n54 VTAIL.n9 0.155672
R457 VTAIL.n61 VTAIL.n9 0.155672
R458 VTAIL.n62 VTAIL.n61 0.155672
R459 VTAIL.n62 VTAIL.n5 0.155672
R460 VTAIL.n70 VTAIL.n5 0.155672
R461 VTAIL.n71 VTAIL.n70 0.155672
R462 VTAIL.n71 VTAIL.n1 0.155672
R463 VTAIL.n79 VTAIL.n1 0.155672
R464 VTAIL.n243 VTAIL.n165 0.155672
R465 VTAIL.n235 VTAIL.n165 0.155672
R466 VTAIL.n235 VTAIL.n234 0.155672
R467 VTAIL.n234 VTAIL.n169 0.155672
R468 VTAIL.n227 VTAIL.n169 0.155672
R469 VTAIL.n227 VTAIL.n226 0.155672
R470 VTAIL.n226 VTAIL.n174 0.155672
R471 VTAIL.n219 VTAIL.n174 0.155672
R472 VTAIL.n219 VTAIL.n218 0.155672
R473 VTAIL.n218 VTAIL.n178 0.155672
R474 VTAIL.n211 VTAIL.n178 0.155672
R475 VTAIL.n211 VTAIL.n210 0.155672
R476 VTAIL.n210 VTAIL.n182 0.155672
R477 VTAIL.n203 VTAIL.n182 0.155672
R478 VTAIL.n203 VTAIL.n202 0.155672
R479 VTAIL.n202 VTAIL.n186 0.155672
R480 VTAIL.n195 VTAIL.n186 0.155672
R481 VTAIL.n195 VTAIL.n194 0.155672
R482 VTAIL.n161 VTAIL.n83 0.155672
R483 VTAIL.n153 VTAIL.n83 0.155672
R484 VTAIL.n153 VTAIL.n152 0.155672
R485 VTAIL.n152 VTAIL.n87 0.155672
R486 VTAIL.n145 VTAIL.n87 0.155672
R487 VTAIL.n145 VTAIL.n144 0.155672
R488 VTAIL.n144 VTAIL.n92 0.155672
R489 VTAIL.n137 VTAIL.n92 0.155672
R490 VTAIL.n137 VTAIL.n136 0.155672
R491 VTAIL.n136 VTAIL.n96 0.155672
R492 VTAIL.n129 VTAIL.n96 0.155672
R493 VTAIL.n129 VTAIL.n128 0.155672
R494 VTAIL.n128 VTAIL.n100 0.155672
R495 VTAIL.n121 VTAIL.n100 0.155672
R496 VTAIL.n121 VTAIL.n120 0.155672
R497 VTAIL.n120 VTAIL.n104 0.155672
R498 VTAIL.n113 VTAIL.n104 0.155672
R499 VTAIL.n113 VTAIL.n112 0.155672
R500 VDD1.n76 VDD1.n0 756.745
R501 VDD1.n157 VDD1.n81 756.745
R502 VDD1.n77 VDD1.n76 585
R503 VDD1.n75 VDD1.n74 585
R504 VDD1.n73 VDD1.n3 585
R505 VDD1.n7 VDD1.n4 585
R506 VDD1.n68 VDD1.n67 585
R507 VDD1.n66 VDD1.n65 585
R508 VDD1.n9 VDD1.n8 585
R509 VDD1.n60 VDD1.n59 585
R510 VDD1.n58 VDD1.n57 585
R511 VDD1.n13 VDD1.n12 585
R512 VDD1.n52 VDD1.n51 585
R513 VDD1.n50 VDD1.n49 585
R514 VDD1.n17 VDD1.n16 585
R515 VDD1.n44 VDD1.n43 585
R516 VDD1.n42 VDD1.n41 585
R517 VDD1.n21 VDD1.n20 585
R518 VDD1.n36 VDD1.n35 585
R519 VDD1.n34 VDD1.n33 585
R520 VDD1.n25 VDD1.n24 585
R521 VDD1.n28 VDD1.n27 585
R522 VDD1.n108 VDD1.n107 585
R523 VDD1.n105 VDD1.n104 585
R524 VDD1.n114 VDD1.n113 585
R525 VDD1.n116 VDD1.n115 585
R526 VDD1.n101 VDD1.n100 585
R527 VDD1.n122 VDD1.n121 585
R528 VDD1.n124 VDD1.n123 585
R529 VDD1.n97 VDD1.n96 585
R530 VDD1.n130 VDD1.n129 585
R531 VDD1.n132 VDD1.n131 585
R532 VDD1.n93 VDD1.n92 585
R533 VDD1.n138 VDD1.n137 585
R534 VDD1.n140 VDD1.n139 585
R535 VDD1.n89 VDD1.n88 585
R536 VDD1.n146 VDD1.n145 585
R537 VDD1.n149 VDD1.n148 585
R538 VDD1.n147 VDD1.n85 585
R539 VDD1.n154 VDD1.n84 585
R540 VDD1.n156 VDD1.n155 585
R541 VDD1.n158 VDD1.n157 585
R542 VDD1.t0 VDD1.n26 327.466
R543 VDD1.t1 VDD1.n106 327.466
R544 VDD1.n76 VDD1.n75 171.744
R545 VDD1.n75 VDD1.n3 171.744
R546 VDD1.n7 VDD1.n3 171.744
R547 VDD1.n67 VDD1.n7 171.744
R548 VDD1.n67 VDD1.n66 171.744
R549 VDD1.n66 VDD1.n8 171.744
R550 VDD1.n59 VDD1.n8 171.744
R551 VDD1.n59 VDD1.n58 171.744
R552 VDD1.n58 VDD1.n12 171.744
R553 VDD1.n51 VDD1.n12 171.744
R554 VDD1.n51 VDD1.n50 171.744
R555 VDD1.n50 VDD1.n16 171.744
R556 VDD1.n43 VDD1.n16 171.744
R557 VDD1.n43 VDD1.n42 171.744
R558 VDD1.n42 VDD1.n20 171.744
R559 VDD1.n35 VDD1.n20 171.744
R560 VDD1.n35 VDD1.n34 171.744
R561 VDD1.n34 VDD1.n24 171.744
R562 VDD1.n27 VDD1.n24 171.744
R563 VDD1.n107 VDD1.n104 171.744
R564 VDD1.n114 VDD1.n104 171.744
R565 VDD1.n115 VDD1.n114 171.744
R566 VDD1.n115 VDD1.n100 171.744
R567 VDD1.n122 VDD1.n100 171.744
R568 VDD1.n123 VDD1.n122 171.744
R569 VDD1.n123 VDD1.n96 171.744
R570 VDD1.n130 VDD1.n96 171.744
R571 VDD1.n131 VDD1.n130 171.744
R572 VDD1.n131 VDD1.n92 171.744
R573 VDD1.n138 VDD1.n92 171.744
R574 VDD1.n139 VDD1.n138 171.744
R575 VDD1.n139 VDD1.n88 171.744
R576 VDD1.n146 VDD1.n88 171.744
R577 VDD1.n148 VDD1.n146 171.744
R578 VDD1.n148 VDD1.n147 171.744
R579 VDD1.n147 VDD1.n84 171.744
R580 VDD1.n156 VDD1.n84 171.744
R581 VDD1.n157 VDD1.n156 171.744
R582 VDD1 VDD1.n161 93.7786
R583 VDD1.n27 VDD1.t0 85.8723
R584 VDD1.n107 VDD1.t1 85.8723
R585 VDD1 VDD1.n80 52.5663
R586 VDD1.n28 VDD1.n26 16.3895
R587 VDD1.n108 VDD1.n106 16.3895
R588 VDD1.n74 VDD1.n73 13.1884
R589 VDD1.n155 VDD1.n154 13.1884
R590 VDD1.n77 VDD1.n2 12.8005
R591 VDD1.n72 VDD1.n4 12.8005
R592 VDD1.n29 VDD1.n25 12.8005
R593 VDD1.n109 VDD1.n105 12.8005
R594 VDD1.n153 VDD1.n85 12.8005
R595 VDD1.n158 VDD1.n83 12.8005
R596 VDD1.n78 VDD1.n0 12.0247
R597 VDD1.n69 VDD1.n68 12.0247
R598 VDD1.n33 VDD1.n32 12.0247
R599 VDD1.n113 VDD1.n112 12.0247
R600 VDD1.n150 VDD1.n149 12.0247
R601 VDD1.n159 VDD1.n81 12.0247
R602 VDD1.n65 VDD1.n6 11.249
R603 VDD1.n36 VDD1.n23 11.249
R604 VDD1.n116 VDD1.n103 11.249
R605 VDD1.n145 VDD1.n87 11.249
R606 VDD1.n64 VDD1.n9 10.4732
R607 VDD1.n37 VDD1.n21 10.4732
R608 VDD1.n117 VDD1.n101 10.4732
R609 VDD1.n144 VDD1.n89 10.4732
R610 VDD1.n61 VDD1.n60 9.69747
R611 VDD1.n41 VDD1.n40 9.69747
R612 VDD1.n121 VDD1.n120 9.69747
R613 VDD1.n141 VDD1.n140 9.69747
R614 VDD1.n80 VDD1.n79 9.45567
R615 VDD1.n161 VDD1.n160 9.45567
R616 VDD1.n54 VDD1.n53 9.3005
R617 VDD1.n56 VDD1.n55 9.3005
R618 VDD1.n11 VDD1.n10 9.3005
R619 VDD1.n62 VDD1.n61 9.3005
R620 VDD1.n64 VDD1.n63 9.3005
R621 VDD1.n6 VDD1.n5 9.3005
R622 VDD1.n70 VDD1.n69 9.3005
R623 VDD1.n72 VDD1.n71 9.3005
R624 VDD1.n79 VDD1.n78 9.3005
R625 VDD1.n2 VDD1.n1 9.3005
R626 VDD1.n15 VDD1.n14 9.3005
R627 VDD1.n48 VDD1.n47 9.3005
R628 VDD1.n46 VDD1.n45 9.3005
R629 VDD1.n19 VDD1.n18 9.3005
R630 VDD1.n40 VDD1.n39 9.3005
R631 VDD1.n38 VDD1.n37 9.3005
R632 VDD1.n23 VDD1.n22 9.3005
R633 VDD1.n32 VDD1.n31 9.3005
R634 VDD1.n30 VDD1.n29 9.3005
R635 VDD1.n160 VDD1.n159 9.3005
R636 VDD1.n83 VDD1.n82 9.3005
R637 VDD1.n128 VDD1.n127 9.3005
R638 VDD1.n126 VDD1.n125 9.3005
R639 VDD1.n99 VDD1.n98 9.3005
R640 VDD1.n120 VDD1.n119 9.3005
R641 VDD1.n118 VDD1.n117 9.3005
R642 VDD1.n103 VDD1.n102 9.3005
R643 VDD1.n112 VDD1.n111 9.3005
R644 VDD1.n110 VDD1.n109 9.3005
R645 VDD1.n95 VDD1.n94 9.3005
R646 VDD1.n134 VDD1.n133 9.3005
R647 VDD1.n136 VDD1.n135 9.3005
R648 VDD1.n91 VDD1.n90 9.3005
R649 VDD1.n142 VDD1.n141 9.3005
R650 VDD1.n144 VDD1.n143 9.3005
R651 VDD1.n87 VDD1.n86 9.3005
R652 VDD1.n151 VDD1.n150 9.3005
R653 VDD1.n153 VDD1.n152 9.3005
R654 VDD1.n57 VDD1.n11 8.92171
R655 VDD1.n44 VDD1.n19 8.92171
R656 VDD1.n124 VDD1.n99 8.92171
R657 VDD1.n137 VDD1.n91 8.92171
R658 VDD1.n56 VDD1.n13 8.14595
R659 VDD1.n45 VDD1.n17 8.14595
R660 VDD1.n125 VDD1.n97 8.14595
R661 VDD1.n136 VDD1.n93 8.14595
R662 VDD1.n53 VDD1.n52 7.3702
R663 VDD1.n49 VDD1.n48 7.3702
R664 VDD1.n129 VDD1.n128 7.3702
R665 VDD1.n133 VDD1.n132 7.3702
R666 VDD1.n52 VDD1.n15 6.59444
R667 VDD1.n49 VDD1.n15 6.59444
R668 VDD1.n129 VDD1.n95 6.59444
R669 VDD1.n132 VDD1.n95 6.59444
R670 VDD1.n53 VDD1.n13 5.81868
R671 VDD1.n48 VDD1.n17 5.81868
R672 VDD1.n128 VDD1.n97 5.81868
R673 VDD1.n133 VDD1.n93 5.81868
R674 VDD1.n57 VDD1.n56 5.04292
R675 VDD1.n45 VDD1.n44 5.04292
R676 VDD1.n125 VDD1.n124 5.04292
R677 VDD1.n137 VDD1.n136 5.04292
R678 VDD1.n60 VDD1.n11 4.26717
R679 VDD1.n41 VDD1.n19 4.26717
R680 VDD1.n121 VDD1.n99 4.26717
R681 VDD1.n140 VDD1.n91 4.26717
R682 VDD1.n30 VDD1.n26 3.70982
R683 VDD1.n110 VDD1.n106 3.70982
R684 VDD1.n61 VDD1.n9 3.49141
R685 VDD1.n40 VDD1.n21 3.49141
R686 VDD1.n120 VDD1.n101 3.49141
R687 VDD1.n141 VDD1.n89 3.49141
R688 VDD1.n65 VDD1.n64 2.71565
R689 VDD1.n37 VDD1.n36 2.71565
R690 VDD1.n117 VDD1.n116 2.71565
R691 VDD1.n145 VDD1.n144 2.71565
R692 VDD1.n80 VDD1.n0 1.93989
R693 VDD1.n68 VDD1.n6 1.93989
R694 VDD1.n33 VDD1.n23 1.93989
R695 VDD1.n113 VDD1.n103 1.93989
R696 VDD1.n149 VDD1.n87 1.93989
R697 VDD1.n161 VDD1.n81 1.93989
R698 VDD1.n78 VDD1.n77 1.16414
R699 VDD1.n69 VDD1.n4 1.16414
R700 VDD1.n32 VDD1.n25 1.16414
R701 VDD1.n112 VDD1.n105 1.16414
R702 VDD1.n150 VDD1.n85 1.16414
R703 VDD1.n159 VDD1.n158 1.16414
R704 VDD1.n74 VDD1.n2 0.388379
R705 VDD1.n73 VDD1.n72 0.388379
R706 VDD1.n29 VDD1.n28 0.388379
R707 VDD1.n109 VDD1.n108 0.388379
R708 VDD1.n154 VDD1.n153 0.388379
R709 VDD1.n155 VDD1.n83 0.388379
R710 VDD1.n79 VDD1.n1 0.155672
R711 VDD1.n71 VDD1.n1 0.155672
R712 VDD1.n71 VDD1.n70 0.155672
R713 VDD1.n70 VDD1.n5 0.155672
R714 VDD1.n63 VDD1.n5 0.155672
R715 VDD1.n63 VDD1.n62 0.155672
R716 VDD1.n62 VDD1.n10 0.155672
R717 VDD1.n55 VDD1.n10 0.155672
R718 VDD1.n55 VDD1.n54 0.155672
R719 VDD1.n54 VDD1.n14 0.155672
R720 VDD1.n47 VDD1.n14 0.155672
R721 VDD1.n47 VDD1.n46 0.155672
R722 VDD1.n46 VDD1.n18 0.155672
R723 VDD1.n39 VDD1.n18 0.155672
R724 VDD1.n39 VDD1.n38 0.155672
R725 VDD1.n38 VDD1.n22 0.155672
R726 VDD1.n31 VDD1.n22 0.155672
R727 VDD1.n31 VDD1.n30 0.155672
R728 VDD1.n111 VDD1.n110 0.155672
R729 VDD1.n111 VDD1.n102 0.155672
R730 VDD1.n118 VDD1.n102 0.155672
R731 VDD1.n119 VDD1.n118 0.155672
R732 VDD1.n119 VDD1.n98 0.155672
R733 VDD1.n126 VDD1.n98 0.155672
R734 VDD1.n127 VDD1.n126 0.155672
R735 VDD1.n127 VDD1.n94 0.155672
R736 VDD1.n134 VDD1.n94 0.155672
R737 VDD1.n135 VDD1.n134 0.155672
R738 VDD1.n135 VDD1.n90 0.155672
R739 VDD1.n142 VDD1.n90 0.155672
R740 VDD1.n143 VDD1.n142 0.155672
R741 VDD1.n143 VDD1.n86 0.155672
R742 VDD1.n151 VDD1.n86 0.155672
R743 VDD1.n152 VDD1.n151 0.155672
R744 VDD1.n152 VDD1.n82 0.155672
R745 VDD1.n160 VDD1.n82 0.155672
R746 B.n436 B.n435 585
R747 B.n437 B.n72 585
R748 B.n439 B.n438 585
R749 B.n440 B.n71 585
R750 B.n442 B.n441 585
R751 B.n443 B.n70 585
R752 B.n445 B.n444 585
R753 B.n446 B.n69 585
R754 B.n448 B.n447 585
R755 B.n449 B.n68 585
R756 B.n451 B.n450 585
R757 B.n452 B.n67 585
R758 B.n454 B.n453 585
R759 B.n455 B.n66 585
R760 B.n457 B.n456 585
R761 B.n458 B.n65 585
R762 B.n460 B.n459 585
R763 B.n461 B.n64 585
R764 B.n463 B.n462 585
R765 B.n464 B.n63 585
R766 B.n466 B.n465 585
R767 B.n467 B.n62 585
R768 B.n469 B.n468 585
R769 B.n470 B.n61 585
R770 B.n472 B.n471 585
R771 B.n473 B.n60 585
R772 B.n475 B.n474 585
R773 B.n476 B.n59 585
R774 B.n478 B.n477 585
R775 B.n479 B.n58 585
R776 B.n481 B.n480 585
R777 B.n482 B.n57 585
R778 B.n484 B.n483 585
R779 B.n485 B.n56 585
R780 B.n487 B.n486 585
R781 B.n488 B.n55 585
R782 B.n490 B.n489 585
R783 B.n491 B.n54 585
R784 B.n493 B.n492 585
R785 B.n494 B.n53 585
R786 B.n496 B.n495 585
R787 B.n497 B.n52 585
R788 B.n499 B.n498 585
R789 B.n500 B.n51 585
R790 B.n502 B.n501 585
R791 B.n503 B.n50 585
R792 B.n505 B.n504 585
R793 B.n506 B.n49 585
R794 B.n508 B.n507 585
R795 B.n509 B.n46 585
R796 B.n512 B.n511 585
R797 B.n513 B.n45 585
R798 B.n515 B.n514 585
R799 B.n516 B.n44 585
R800 B.n518 B.n517 585
R801 B.n519 B.n43 585
R802 B.n521 B.n520 585
R803 B.n522 B.n39 585
R804 B.n524 B.n523 585
R805 B.n525 B.n38 585
R806 B.n527 B.n526 585
R807 B.n528 B.n37 585
R808 B.n530 B.n529 585
R809 B.n531 B.n36 585
R810 B.n533 B.n532 585
R811 B.n534 B.n35 585
R812 B.n536 B.n535 585
R813 B.n537 B.n34 585
R814 B.n539 B.n538 585
R815 B.n540 B.n33 585
R816 B.n542 B.n541 585
R817 B.n543 B.n32 585
R818 B.n545 B.n544 585
R819 B.n546 B.n31 585
R820 B.n548 B.n547 585
R821 B.n549 B.n30 585
R822 B.n551 B.n550 585
R823 B.n552 B.n29 585
R824 B.n554 B.n553 585
R825 B.n555 B.n28 585
R826 B.n557 B.n556 585
R827 B.n558 B.n27 585
R828 B.n560 B.n559 585
R829 B.n561 B.n26 585
R830 B.n563 B.n562 585
R831 B.n564 B.n25 585
R832 B.n566 B.n565 585
R833 B.n567 B.n24 585
R834 B.n569 B.n568 585
R835 B.n570 B.n23 585
R836 B.n572 B.n571 585
R837 B.n573 B.n22 585
R838 B.n575 B.n574 585
R839 B.n576 B.n21 585
R840 B.n578 B.n577 585
R841 B.n579 B.n20 585
R842 B.n581 B.n580 585
R843 B.n582 B.n19 585
R844 B.n584 B.n583 585
R845 B.n585 B.n18 585
R846 B.n587 B.n586 585
R847 B.n588 B.n17 585
R848 B.n590 B.n589 585
R849 B.n591 B.n16 585
R850 B.n593 B.n592 585
R851 B.n594 B.n15 585
R852 B.n596 B.n595 585
R853 B.n597 B.n14 585
R854 B.n599 B.n598 585
R855 B.n434 B.n73 585
R856 B.n433 B.n432 585
R857 B.n431 B.n74 585
R858 B.n430 B.n429 585
R859 B.n428 B.n75 585
R860 B.n427 B.n426 585
R861 B.n425 B.n76 585
R862 B.n424 B.n423 585
R863 B.n422 B.n77 585
R864 B.n421 B.n420 585
R865 B.n419 B.n78 585
R866 B.n418 B.n417 585
R867 B.n416 B.n79 585
R868 B.n415 B.n414 585
R869 B.n413 B.n80 585
R870 B.n412 B.n411 585
R871 B.n410 B.n81 585
R872 B.n409 B.n408 585
R873 B.n407 B.n82 585
R874 B.n406 B.n405 585
R875 B.n404 B.n83 585
R876 B.n403 B.n402 585
R877 B.n401 B.n84 585
R878 B.n400 B.n399 585
R879 B.n398 B.n85 585
R880 B.n397 B.n396 585
R881 B.n395 B.n86 585
R882 B.n394 B.n393 585
R883 B.n392 B.n87 585
R884 B.n391 B.n390 585
R885 B.n389 B.n88 585
R886 B.n388 B.n387 585
R887 B.n386 B.n89 585
R888 B.n385 B.n384 585
R889 B.n383 B.n90 585
R890 B.n382 B.n381 585
R891 B.n380 B.n91 585
R892 B.n379 B.n378 585
R893 B.n377 B.n92 585
R894 B.n376 B.n375 585
R895 B.n374 B.n93 585
R896 B.n373 B.n372 585
R897 B.n371 B.n94 585
R898 B.n370 B.n369 585
R899 B.n368 B.n95 585
R900 B.n367 B.n366 585
R901 B.n365 B.n96 585
R902 B.n198 B.n197 585
R903 B.n199 B.n152 585
R904 B.n201 B.n200 585
R905 B.n202 B.n151 585
R906 B.n204 B.n203 585
R907 B.n205 B.n150 585
R908 B.n207 B.n206 585
R909 B.n208 B.n149 585
R910 B.n210 B.n209 585
R911 B.n211 B.n148 585
R912 B.n213 B.n212 585
R913 B.n214 B.n147 585
R914 B.n216 B.n215 585
R915 B.n217 B.n146 585
R916 B.n219 B.n218 585
R917 B.n220 B.n145 585
R918 B.n222 B.n221 585
R919 B.n223 B.n144 585
R920 B.n225 B.n224 585
R921 B.n226 B.n143 585
R922 B.n228 B.n227 585
R923 B.n229 B.n142 585
R924 B.n231 B.n230 585
R925 B.n232 B.n141 585
R926 B.n234 B.n233 585
R927 B.n235 B.n140 585
R928 B.n237 B.n236 585
R929 B.n238 B.n139 585
R930 B.n240 B.n239 585
R931 B.n241 B.n138 585
R932 B.n243 B.n242 585
R933 B.n244 B.n137 585
R934 B.n246 B.n245 585
R935 B.n247 B.n136 585
R936 B.n249 B.n248 585
R937 B.n250 B.n135 585
R938 B.n252 B.n251 585
R939 B.n253 B.n134 585
R940 B.n255 B.n254 585
R941 B.n256 B.n133 585
R942 B.n258 B.n257 585
R943 B.n259 B.n132 585
R944 B.n261 B.n260 585
R945 B.n262 B.n131 585
R946 B.n264 B.n263 585
R947 B.n265 B.n130 585
R948 B.n267 B.n266 585
R949 B.n268 B.n129 585
R950 B.n270 B.n269 585
R951 B.n271 B.n126 585
R952 B.n274 B.n273 585
R953 B.n275 B.n125 585
R954 B.n277 B.n276 585
R955 B.n278 B.n124 585
R956 B.n280 B.n279 585
R957 B.n281 B.n123 585
R958 B.n283 B.n282 585
R959 B.n284 B.n122 585
R960 B.n289 B.n288 585
R961 B.n290 B.n121 585
R962 B.n292 B.n291 585
R963 B.n293 B.n120 585
R964 B.n295 B.n294 585
R965 B.n296 B.n119 585
R966 B.n298 B.n297 585
R967 B.n299 B.n118 585
R968 B.n301 B.n300 585
R969 B.n302 B.n117 585
R970 B.n304 B.n303 585
R971 B.n305 B.n116 585
R972 B.n307 B.n306 585
R973 B.n308 B.n115 585
R974 B.n310 B.n309 585
R975 B.n311 B.n114 585
R976 B.n313 B.n312 585
R977 B.n314 B.n113 585
R978 B.n316 B.n315 585
R979 B.n317 B.n112 585
R980 B.n319 B.n318 585
R981 B.n320 B.n111 585
R982 B.n322 B.n321 585
R983 B.n323 B.n110 585
R984 B.n325 B.n324 585
R985 B.n326 B.n109 585
R986 B.n328 B.n327 585
R987 B.n329 B.n108 585
R988 B.n331 B.n330 585
R989 B.n332 B.n107 585
R990 B.n334 B.n333 585
R991 B.n335 B.n106 585
R992 B.n337 B.n336 585
R993 B.n338 B.n105 585
R994 B.n340 B.n339 585
R995 B.n341 B.n104 585
R996 B.n343 B.n342 585
R997 B.n344 B.n103 585
R998 B.n346 B.n345 585
R999 B.n347 B.n102 585
R1000 B.n349 B.n348 585
R1001 B.n350 B.n101 585
R1002 B.n352 B.n351 585
R1003 B.n353 B.n100 585
R1004 B.n355 B.n354 585
R1005 B.n356 B.n99 585
R1006 B.n358 B.n357 585
R1007 B.n359 B.n98 585
R1008 B.n361 B.n360 585
R1009 B.n362 B.n97 585
R1010 B.n364 B.n363 585
R1011 B.n196 B.n153 585
R1012 B.n195 B.n194 585
R1013 B.n193 B.n154 585
R1014 B.n192 B.n191 585
R1015 B.n190 B.n155 585
R1016 B.n189 B.n188 585
R1017 B.n187 B.n156 585
R1018 B.n186 B.n185 585
R1019 B.n184 B.n157 585
R1020 B.n183 B.n182 585
R1021 B.n181 B.n158 585
R1022 B.n180 B.n179 585
R1023 B.n178 B.n159 585
R1024 B.n177 B.n176 585
R1025 B.n175 B.n160 585
R1026 B.n174 B.n173 585
R1027 B.n172 B.n161 585
R1028 B.n171 B.n170 585
R1029 B.n169 B.n162 585
R1030 B.n168 B.n167 585
R1031 B.n166 B.n163 585
R1032 B.n165 B.n164 585
R1033 B.n2 B.n0 585
R1034 B.n633 B.n1 585
R1035 B.n632 B.n631 585
R1036 B.n630 B.n3 585
R1037 B.n629 B.n628 585
R1038 B.n627 B.n4 585
R1039 B.n626 B.n625 585
R1040 B.n624 B.n5 585
R1041 B.n623 B.n622 585
R1042 B.n621 B.n6 585
R1043 B.n620 B.n619 585
R1044 B.n618 B.n7 585
R1045 B.n617 B.n616 585
R1046 B.n615 B.n8 585
R1047 B.n614 B.n613 585
R1048 B.n612 B.n9 585
R1049 B.n611 B.n610 585
R1050 B.n609 B.n10 585
R1051 B.n608 B.n607 585
R1052 B.n606 B.n11 585
R1053 B.n605 B.n604 585
R1054 B.n603 B.n12 585
R1055 B.n602 B.n601 585
R1056 B.n600 B.n13 585
R1057 B.n635 B.n634 585
R1058 B.n197 B.n196 502.111
R1059 B.n598 B.n13 502.111
R1060 B.n363 B.n96 502.111
R1061 B.n435 B.n434 502.111
R1062 B.n285 B.t2 474.75
R1063 B.n47 B.t10 474.75
R1064 B.n127 B.t5 474.75
R1065 B.n40 B.t7 474.75
R1066 B.n286 B.t1 426.072
R1067 B.n48 B.t11 426.072
R1068 B.n128 B.t4 426.072
R1069 B.n41 B.t8 426.072
R1070 B.n285 B.t0 370.925
R1071 B.n127 B.t3 370.925
R1072 B.n40 B.t6 370.925
R1073 B.n47 B.t9 370.925
R1074 B.n196 B.n195 163.367
R1075 B.n195 B.n154 163.367
R1076 B.n191 B.n154 163.367
R1077 B.n191 B.n190 163.367
R1078 B.n190 B.n189 163.367
R1079 B.n189 B.n156 163.367
R1080 B.n185 B.n156 163.367
R1081 B.n185 B.n184 163.367
R1082 B.n184 B.n183 163.367
R1083 B.n183 B.n158 163.367
R1084 B.n179 B.n158 163.367
R1085 B.n179 B.n178 163.367
R1086 B.n178 B.n177 163.367
R1087 B.n177 B.n160 163.367
R1088 B.n173 B.n160 163.367
R1089 B.n173 B.n172 163.367
R1090 B.n172 B.n171 163.367
R1091 B.n171 B.n162 163.367
R1092 B.n167 B.n162 163.367
R1093 B.n167 B.n166 163.367
R1094 B.n166 B.n165 163.367
R1095 B.n165 B.n2 163.367
R1096 B.n634 B.n2 163.367
R1097 B.n634 B.n633 163.367
R1098 B.n633 B.n632 163.367
R1099 B.n632 B.n3 163.367
R1100 B.n628 B.n3 163.367
R1101 B.n628 B.n627 163.367
R1102 B.n627 B.n626 163.367
R1103 B.n626 B.n5 163.367
R1104 B.n622 B.n5 163.367
R1105 B.n622 B.n621 163.367
R1106 B.n621 B.n620 163.367
R1107 B.n620 B.n7 163.367
R1108 B.n616 B.n7 163.367
R1109 B.n616 B.n615 163.367
R1110 B.n615 B.n614 163.367
R1111 B.n614 B.n9 163.367
R1112 B.n610 B.n9 163.367
R1113 B.n610 B.n609 163.367
R1114 B.n609 B.n608 163.367
R1115 B.n608 B.n11 163.367
R1116 B.n604 B.n11 163.367
R1117 B.n604 B.n603 163.367
R1118 B.n603 B.n602 163.367
R1119 B.n602 B.n13 163.367
R1120 B.n197 B.n152 163.367
R1121 B.n201 B.n152 163.367
R1122 B.n202 B.n201 163.367
R1123 B.n203 B.n202 163.367
R1124 B.n203 B.n150 163.367
R1125 B.n207 B.n150 163.367
R1126 B.n208 B.n207 163.367
R1127 B.n209 B.n208 163.367
R1128 B.n209 B.n148 163.367
R1129 B.n213 B.n148 163.367
R1130 B.n214 B.n213 163.367
R1131 B.n215 B.n214 163.367
R1132 B.n215 B.n146 163.367
R1133 B.n219 B.n146 163.367
R1134 B.n220 B.n219 163.367
R1135 B.n221 B.n220 163.367
R1136 B.n221 B.n144 163.367
R1137 B.n225 B.n144 163.367
R1138 B.n226 B.n225 163.367
R1139 B.n227 B.n226 163.367
R1140 B.n227 B.n142 163.367
R1141 B.n231 B.n142 163.367
R1142 B.n232 B.n231 163.367
R1143 B.n233 B.n232 163.367
R1144 B.n233 B.n140 163.367
R1145 B.n237 B.n140 163.367
R1146 B.n238 B.n237 163.367
R1147 B.n239 B.n238 163.367
R1148 B.n239 B.n138 163.367
R1149 B.n243 B.n138 163.367
R1150 B.n244 B.n243 163.367
R1151 B.n245 B.n244 163.367
R1152 B.n245 B.n136 163.367
R1153 B.n249 B.n136 163.367
R1154 B.n250 B.n249 163.367
R1155 B.n251 B.n250 163.367
R1156 B.n251 B.n134 163.367
R1157 B.n255 B.n134 163.367
R1158 B.n256 B.n255 163.367
R1159 B.n257 B.n256 163.367
R1160 B.n257 B.n132 163.367
R1161 B.n261 B.n132 163.367
R1162 B.n262 B.n261 163.367
R1163 B.n263 B.n262 163.367
R1164 B.n263 B.n130 163.367
R1165 B.n267 B.n130 163.367
R1166 B.n268 B.n267 163.367
R1167 B.n269 B.n268 163.367
R1168 B.n269 B.n126 163.367
R1169 B.n274 B.n126 163.367
R1170 B.n275 B.n274 163.367
R1171 B.n276 B.n275 163.367
R1172 B.n276 B.n124 163.367
R1173 B.n280 B.n124 163.367
R1174 B.n281 B.n280 163.367
R1175 B.n282 B.n281 163.367
R1176 B.n282 B.n122 163.367
R1177 B.n289 B.n122 163.367
R1178 B.n290 B.n289 163.367
R1179 B.n291 B.n290 163.367
R1180 B.n291 B.n120 163.367
R1181 B.n295 B.n120 163.367
R1182 B.n296 B.n295 163.367
R1183 B.n297 B.n296 163.367
R1184 B.n297 B.n118 163.367
R1185 B.n301 B.n118 163.367
R1186 B.n302 B.n301 163.367
R1187 B.n303 B.n302 163.367
R1188 B.n303 B.n116 163.367
R1189 B.n307 B.n116 163.367
R1190 B.n308 B.n307 163.367
R1191 B.n309 B.n308 163.367
R1192 B.n309 B.n114 163.367
R1193 B.n313 B.n114 163.367
R1194 B.n314 B.n313 163.367
R1195 B.n315 B.n314 163.367
R1196 B.n315 B.n112 163.367
R1197 B.n319 B.n112 163.367
R1198 B.n320 B.n319 163.367
R1199 B.n321 B.n320 163.367
R1200 B.n321 B.n110 163.367
R1201 B.n325 B.n110 163.367
R1202 B.n326 B.n325 163.367
R1203 B.n327 B.n326 163.367
R1204 B.n327 B.n108 163.367
R1205 B.n331 B.n108 163.367
R1206 B.n332 B.n331 163.367
R1207 B.n333 B.n332 163.367
R1208 B.n333 B.n106 163.367
R1209 B.n337 B.n106 163.367
R1210 B.n338 B.n337 163.367
R1211 B.n339 B.n338 163.367
R1212 B.n339 B.n104 163.367
R1213 B.n343 B.n104 163.367
R1214 B.n344 B.n343 163.367
R1215 B.n345 B.n344 163.367
R1216 B.n345 B.n102 163.367
R1217 B.n349 B.n102 163.367
R1218 B.n350 B.n349 163.367
R1219 B.n351 B.n350 163.367
R1220 B.n351 B.n100 163.367
R1221 B.n355 B.n100 163.367
R1222 B.n356 B.n355 163.367
R1223 B.n357 B.n356 163.367
R1224 B.n357 B.n98 163.367
R1225 B.n361 B.n98 163.367
R1226 B.n362 B.n361 163.367
R1227 B.n363 B.n362 163.367
R1228 B.n367 B.n96 163.367
R1229 B.n368 B.n367 163.367
R1230 B.n369 B.n368 163.367
R1231 B.n369 B.n94 163.367
R1232 B.n373 B.n94 163.367
R1233 B.n374 B.n373 163.367
R1234 B.n375 B.n374 163.367
R1235 B.n375 B.n92 163.367
R1236 B.n379 B.n92 163.367
R1237 B.n380 B.n379 163.367
R1238 B.n381 B.n380 163.367
R1239 B.n381 B.n90 163.367
R1240 B.n385 B.n90 163.367
R1241 B.n386 B.n385 163.367
R1242 B.n387 B.n386 163.367
R1243 B.n387 B.n88 163.367
R1244 B.n391 B.n88 163.367
R1245 B.n392 B.n391 163.367
R1246 B.n393 B.n392 163.367
R1247 B.n393 B.n86 163.367
R1248 B.n397 B.n86 163.367
R1249 B.n398 B.n397 163.367
R1250 B.n399 B.n398 163.367
R1251 B.n399 B.n84 163.367
R1252 B.n403 B.n84 163.367
R1253 B.n404 B.n403 163.367
R1254 B.n405 B.n404 163.367
R1255 B.n405 B.n82 163.367
R1256 B.n409 B.n82 163.367
R1257 B.n410 B.n409 163.367
R1258 B.n411 B.n410 163.367
R1259 B.n411 B.n80 163.367
R1260 B.n415 B.n80 163.367
R1261 B.n416 B.n415 163.367
R1262 B.n417 B.n416 163.367
R1263 B.n417 B.n78 163.367
R1264 B.n421 B.n78 163.367
R1265 B.n422 B.n421 163.367
R1266 B.n423 B.n422 163.367
R1267 B.n423 B.n76 163.367
R1268 B.n427 B.n76 163.367
R1269 B.n428 B.n427 163.367
R1270 B.n429 B.n428 163.367
R1271 B.n429 B.n74 163.367
R1272 B.n433 B.n74 163.367
R1273 B.n434 B.n433 163.367
R1274 B.n598 B.n597 163.367
R1275 B.n597 B.n596 163.367
R1276 B.n596 B.n15 163.367
R1277 B.n592 B.n15 163.367
R1278 B.n592 B.n591 163.367
R1279 B.n591 B.n590 163.367
R1280 B.n590 B.n17 163.367
R1281 B.n586 B.n17 163.367
R1282 B.n586 B.n585 163.367
R1283 B.n585 B.n584 163.367
R1284 B.n584 B.n19 163.367
R1285 B.n580 B.n19 163.367
R1286 B.n580 B.n579 163.367
R1287 B.n579 B.n578 163.367
R1288 B.n578 B.n21 163.367
R1289 B.n574 B.n21 163.367
R1290 B.n574 B.n573 163.367
R1291 B.n573 B.n572 163.367
R1292 B.n572 B.n23 163.367
R1293 B.n568 B.n23 163.367
R1294 B.n568 B.n567 163.367
R1295 B.n567 B.n566 163.367
R1296 B.n566 B.n25 163.367
R1297 B.n562 B.n25 163.367
R1298 B.n562 B.n561 163.367
R1299 B.n561 B.n560 163.367
R1300 B.n560 B.n27 163.367
R1301 B.n556 B.n27 163.367
R1302 B.n556 B.n555 163.367
R1303 B.n555 B.n554 163.367
R1304 B.n554 B.n29 163.367
R1305 B.n550 B.n29 163.367
R1306 B.n550 B.n549 163.367
R1307 B.n549 B.n548 163.367
R1308 B.n548 B.n31 163.367
R1309 B.n544 B.n31 163.367
R1310 B.n544 B.n543 163.367
R1311 B.n543 B.n542 163.367
R1312 B.n542 B.n33 163.367
R1313 B.n538 B.n33 163.367
R1314 B.n538 B.n537 163.367
R1315 B.n537 B.n536 163.367
R1316 B.n536 B.n35 163.367
R1317 B.n532 B.n35 163.367
R1318 B.n532 B.n531 163.367
R1319 B.n531 B.n530 163.367
R1320 B.n530 B.n37 163.367
R1321 B.n526 B.n37 163.367
R1322 B.n526 B.n525 163.367
R1323 B.n525 B.n524 163.367
R1324 B.n524 B.n39 163.367
R1325 B.n520 B.n39 163.367
R1326 B.n520 B.n519 163.367
R1327 B.n519 B.n518 163.367
R1328 B.n518 B.n44 163.367
R1329 B.n514 B.n44 163.367
R1330 B.n514 B.n513 163.367
R1331 B.n513 B.n512 163.367
R1332 B.n512 B.n46 163.367
R1333 B.n507 B.n46 163.367
R1334 B.n507 B.n506 163.367
R1335 B.n506 B.n505 163.367
R1336 B.n505 B.n50 163.367
R1337 B.n501 B.n50 163.367
R1338 B.n501 B.n500 163.367
R1339 B.n500 B.n499 163.367
R1340 B.n499 B.n52 163.367
R1341 B.n495 B.n52 163.367
R1342 B.n495 B.n494 163.367
R1343 B.n494 B.n493 163.367
R1344 B.n493 B.n54 163.367
R1345 B.n489 B.n54 163.367
R1346 B.n489 B.n488 163.367
R1347 B.n488 B.n487 163.367
R1348 B.n487 B.n56 163.367
R1349 B.n483 B.n56 163.367
R1350 B.n483 B.n482 163.367
R1351 B.n482 B.n481 163.367
R1352 B.n481 B.n58 163.367
R1353 B.n477 B.n58 163.367
R1354 B.n477 B.n476 163.367
R1355 B.n476 B.n475 163.367
R1356 B.n475 B.n60 163.367
R1357 B.n471 B.n60 163.367
R1358 B.n471 B.n470 163.367
R1359 B.n470 B.n469 163.367
R1360 B.n469 B.n62 163.367
R1361 B.n465 B.n62 163.367
R1362 B.n465 B.n464 163.367
R1363 B.n464 B.n463 163.367
R1364 B.n463 B.n64 163.367
R1365 B.n459 B.n64 163.367
R1366 B.n459 B.n458 163.367
R1367 B.n458 B.n457 163.367
R1368 B.n457 B.n66 163.367
R1369 B.n453 B.n66 163.367
R1370 B.n453 B.n452 163.367
R1371 B.n452 B.n451 163.367
R1372 B.n451 B.n68 163.367
R1373 B.n447 B.n68 163.367
R1374 B.n447 B.n446 163.367
R1375 B.n446 B.n445 163.367
R1376 B.n445 B.n70 163.367
R1377 B.n441 B.n70 163.367
R1378 B.n441 B.n440 163.367
R1379 B.n440 B.n439 163.367
R1380 B.n439 B.n72 163.367
R1381 B.n435 B.n72 163.367
R1382 B.n287 B.n286 59.5399
R1383 B.n272 B.n128 59.5399
R1384 B.n42 B.n41 59.5399
R1385 B.n510 B.n48 59.5399
R1386 B.n286 B.n285 48.6793
R1387 B.n128 B.n127 48.6793
R1388 B.n41 B.n40 48.6793
R1389 B.n48 B.n47 48.6793
R1390 B.n600 B.n599 32.6249
R1391 B.n436 B.n73 32.6249
R1392 B.n365 B.n364 32.6249
R1393 B.n198 B.n153 32.6249
R1394 B B.n635 18.0485
R1395 B.n599 B.n14 10.6151
R1396 B.n595 B.n14 10.6151
R1397 B.n595 B.n594 10.6151
R1398 B.n594 B.n593 10.6151
R1399 B.n593 B.n16 10.6151
R1400 B.n589 B.n16 10.6151
R1401 B.n589 B.n588 10.6151
R1402 B.n588 B.n587 10.6151
R1403 B.n587 B.n18 10.6151
R1404 B.n583 B.n18 10.6151
R1405 B.n583 B.n582 10.6151
R1406 B.n582 B.n581 10.6151
R1407 B.n581 B.n20 10.6151
R1408 B.n577 B.n20 10.6151
R1409 B.n577 B.n576 10.6151
R1410 B.n576 B.n575 10.6151
R1411 B.n575 B.n22 10.6151
R1412 B.n571 B.n22 10.6151
R1413 B.n571 B.n570 10.6151
R1414 B.n570 B.n569 10.6151
R1415 B.n569 B.n24 10.6151
R1416 B.n565 B.n24 10.6151
R1417 B.n565 B.n564 10.6151
R1418 B.n564 B.n563 10.6151
R1419 B.n563 B.n26 10.6151
R1420 B.n559 B.n26 10.6151
R1421 B.n559 B.n558 10.6151
R1422 B.n558 B.n557 10.6151
R1423 B.n557 B.n28 10.6151
R1424 B.n553 B.n28 10.6151
R1425 B.n553 B.n552 10.6151
R1426 B.n552 B.n551 10.6151
R1427 B.n551 B.n30 10.6151
R1428 B.n547 B.n30 10.6151
R1429 B.n547 B.n546 10.6151
R1430 B.n546 B.n545 10.6151
R1431 B.n545 B.n32 10.6151
R1432 B.n541 B.n32 10.6151
R1433 B.n541 B.n540 10.6151
R1434 B.n540 B.n539 10.6151
R1435 B.n539 B.n34 10.6151
R1436 B.n535 B.n34 10.6151
R1437 B.n535 B.n534 10.6151
R1438 B.n534 B.n533 10.6151
R1439 B.n533 B.n36 10.6151
R1440 B.n529 B.n36 10.6151
R1441 B.n529 B.n528 10.6151
R1442 B.n528 B.n527 10.6151
R1443 B.n527 B.n38 10.6151
R1444 B.n523 B.n522 10.6151
R1445 B.n522 B.n521 10.6151
R1446 B.n521 B.n43 10.6151
R1447 B.n517 B.n43 10.6151
R1448 B.n517 B.n516 10.6151
R1449 B.n516 B.n515 10.6151
R1450 B.n515 B.n45 10.6151
R1451 B.n511 B.n45 10.6151
R1452 B.n509 B.n508 10.6151
R1453 B.n508 B.n49 10.6151
R1454 B.n504 B.n49 10.6151
R1455 B.n504 B.n503 10.6151
R1456 B.n503 B.n502 10.6151
R1457 B.n502 B.n51 10.6151
R1458 B.n498 B.n51 10.6151
R1459 B.n498 B.n497 10.6151
R1460 B.n497 B.n496 10.6151
R1461 B.n496 B.n53 10.6151
R1462 B.n492 B.n53 10.6151
R1463 B.n492 B.n491 10.6151
R1464 B.n491 B.n490 10.6151
R1465 B.n490 B.n55 10.6151
R1466 B.n486 B.n55 10.6151
R1467 B.n486 B.n485 10.6151
R1468 B.n485 B.n484 10.6151
R1469 B.n484 B.n57 10.6151
R1470 B.n480 B.n57 10.6151
R1471 B.n480 B.n479 10.6151
R1472 B.n479 B.n478 10.6151
R1473 B.n478 B.n59 10.6151
R1474 B.n474 B.n59 10.6151
R1475 B.n474 B.n473 10.6151
R1476 B.n473 B.n472 10.6151
R1477 B.n472 B.n61 10.6151
R1478 B.n468 B.n61 10.6151
R1479 B.n468 B.n467 10.6151
R1480 B.n467 B.n466 10.6151
R1481 B.n466 B.n63 10.6151
R1482 B.n462 B.n63 10.6151
R1483 B.n462 B.n461 10.6151
R1484 B.n461 B.n460 10.6151
R1485 B.n460 B.n65 10.6151
R1486 B.n456 B.n65 10.6151
R1487 B.n456 B.n455 10.6151
R1488 B.n455 B.n454 10.6151
R1489 B.n454 B.n67 10.6151
R1490 B.n450 B.n67 10.6151
R1491 B.n450 B.n449 10.6151
R1492 B.n449 B.n448 10.6151
R1493 B.n448 B.n69 10.6151
R1494 B.n444 B.n69 10.6151
R1495 B.n444 B.n443 10.6151
R1496 B.n443 B.n442 10.6151
R1497 B.n442 B.n71 10.6151
R1498 B.n438 B.n71 10.6151
R1499 B.n438 B.n437 10.6151
R1500 B.n437 B.n436 10.6151
R1501 B.n366 B.n365 10.6151
R1502 B.n366 B.n95 10.6151
R1503 B.n370 B.n95 10.6151
R1504 B.n371 B.n370 10.6151
R1505 B.n372 B.n371 10.6151
R1506 B.n372 B.n93 10.6151
R1507 B.n376 B.n93 10.6151
R1508 B.n377 B.n376 10.6151
R1509 B.n378 B.n377 10.6151
R1510 B.n378 B.n91 10.6151
R1511 B.n382 B.n91 10.6151
R1512 B.n383 B.n382 10.6151
R1513 B.n384 B.n383 10.6151
R1514 B.n384 B.n89 10.6151
R1515 B.n388 B.n89 10.6151
R1516 B.n389 B.n388 10.6151
R1517 B.n390 B.n389 10.6151
R1518 B.n390 B.n87 10.6151
R1519 B.n394 B.n87 10.6151
R1520 B.n395 B.n394 10.6151
R1521 B.n396 B.n395 10.6151
R1522 B.n396 B.n85 10.6151
R1523 B.n400 B.n85 10.6151
R1524 B.n401 B.n400 10.6151
R1525 B.n402 B.n401 10.6151
R1526 B.n402 B.n83 10.6151
R1527 B.n406 B.n83 10.6151
R1528 B.n407 B.n406 10.6151
R1529 B.n408 B.n407 10.6151
R1530 B.n408 B.n81 10.6151
R1531 B.n412 B.n81 10.6151
R1532 B.n413 B.n412 10.6151
R1533 B.n414 B.n413 10.6151
R1534 B.n414 B.n79 10.6151
R1535 B.n418 B.n79 10.6151
R1536 B.n419 B.n418 10.6151
R1537 B.n420 B.n419 10.6151
R1538 B.n420 B.n77 10.6151
R1539 B.n424 B.n77 10.6151
R1540 B.n425 B.n424 10.6151
R1541 B.n426 B.n425 10.6151
R1542 B.n426 B.n75 10.6151
R1543 B.n430 B.n75 10.6151
R1544 B.n431 B.n430 10.6151
R1545 B.n432 B.n431 10.6151
R1546 B.n432 B.n73 10.6151
R1547 B.n199 B.n198 10.6151
R1548 B.n200 B.n199 10.6151
R1549 B.n200 B.n151 10.6151
R1550 B.n204 B.n151 10.6151
R1551 B.n205 B.n204 10.6151
R1552 B.n206 B.n205 10.6151
R1553 B.n206 B.n149 10.6151
R1554 B.n210 B.n149 10.6151
R1555 B.n211 B.n210 10.6151
R1556 B.n212 B.n211 10.6151
R1557 B.n212 B.n147 10.6151
R1558 B.n216 B.n147 10.6151
R1559 B.n217 B.n216 10.6151
R1560 B.n218 B.n217 10.6151
R1561 B.n218 B.n145 10.6151
R1562 B.n222 B.n145 10.6151
R1563 B.n223 B.n222 10.6151
R1564 B.n224 B.n223 10.6151
R1565 B.n224 B.n143 10.6151
R1566 B.n228 B.n143 10.6151
R1567 B.n229 B.n228 10.6151
R1568 B.n230 B.n229 10.6151
R1569 B.n230 B.n141 10.6151
R1570 B.n234 B.n141 10.6151
R1571 B.n235 B.n234 10.6151
R1572 B.n236 B.n235 10.6151
R1573 B.n236 B.n139 10.6151
R1574 B.n240 B.n139 10.6151
R1575 B.n241 B.n240 10.6151
R1576 B.n242 B.n241 10.6151
R1577 B.n242 B.n137 10.6151
R1578 B.n246 B.n137 10.6151
R1579 B.n247 B.n246 10.6151
R1580 B.n248 B.n247 10.6151
R1581 B.n248 B.n135 10.6151
R1582 B.n252 B.n135 10.6151
R1583 B.n253 B.n252 10.6151
R1584 B.n254 B.n253 10.6151
R1585 B.n254 B.n133 10.6151
R1586 B.n258 B.n133 10.6151
R1587 B.n259 B.n258 10.6151
R1588 B.n260 B.n259 10.6151
R1589 B.n260 B.n131 10.6151
R1590 B.n264 B.n131 10.6151
R1591 B.n265 B.n264 10.6151
R1592 B.n266 B.n265 10.6151
R1593 B.n266 B.n129 10.6151
R1594 B.n270 B.n129 10.6151
R1595 B.n271 B.n270 10.6151
R1596 B.n273 B.n125 10.6151
R1597 B.n277 B.n125 10.6151
R1598 B.n278 B.n277 10.6151
R1599 B.n279 B.n278 10.6151
R1600 B.n279 B.n123 10.6151
R1601 B.n283 B.n123 10.6151
R1602 B.n284 B.n283 10.6151
R1603 B.n288 B.n284 10.6151
R1604 B.n292 B.n121 10.6151
R1605 B.n293 B.n292 10.6151
R1606 B.n294 B.n293 10.6151
R1607 B.n294 B.n119 10.6151
R1608 B.n298 B.n119 10.6151
R1609 B.n299 B.n298 10.6151
R1610 B.n300 B.n299 10.6151
R1611 B.n300 B.n117 10.6151
R1612 B.n304 B.n117 10.6151
R1613 B.n305 B.n304 10.6151
R1614 B.n306 B.n305 10.6151
R1615 B.n306 B.n115 10.6151
R1616 B.n310 B.n115 10.6151
R1617 B.n311 B.n310 10.6151
R1618 B.n312 B.n311 10.6151
R1619 B.n312 B.n113 10.6151
R1620 B.n316 B.n113 10.6151
R1621 B.n317 B.n316 10.6151
R1622 B.n318 B.n317 10.6151
R1623 B.n318 B.n111 10.6151
R1624 B.n322 B.n111 10.6151
R1625 B.n323 B.n322 10.6151
R1626 B.n324 B.n323 10.6151
R1627 B.n324 B.n109 10.6151
R1628 B.n328 B.n109 10.6151
R1629 B.n329 B.n328 10.6151
R1630 B.n330 B.n329 10.6151
R1631 B.n330 B.n107 10.6151
R1632 B.n334 B.n107 10.6151
R1633 B.n335 B.n334 10.6151
R1634 B.n336 B.n335 10.6151
R1635 B.n336 B.n105 10.6151
R1636 B.n340 B.n105 10.6151
R1637 B.n341 B.n340 10.6151
R1638 B.n342 B.n341 10.6151
R1639 B.n342 B.n103 10.6151
R1640 B.n346 B.n103 10.6151
R1641 B.n347 B.n346 10.6151
R1642 B.n348 B.n347 10.6151
R1643 B.n348 B.n101 10.6151
R1644 B.n352 B.n101 10.6151
R1645 B.n353 B.n352 10.6151
R1646 B.n354 B.n353 10.6151
R1647 B.n354 B.n99 10.6151
R1648 B.n358 B.n99 10.6151
R1649 B.n359 B.n358 10.6151
R1650 B.n360 B.n359 10.6151
R1651 B.n360 B.n97 10.6151
R1652 B.n364 B.n97 10.6151
R1653 B.n194 B.n153 10.6151
R1654 B.n194 B.n193 10.6151
R1655 B.n193 B.n192 10.6151
R1656 B.n192 B.n155 10.6151
R1657 B.n188 B.n155 10.6151
R1658 B.n188 B.n187 10.6151
R1659 B.n187 B.n186 10.6151
R1660 B.n186 B.n157 10.6151
R1661 B.n182 B.n157 10.6151
R1662 B.n182 B.n181 10.6151
R1663 B.n181 B.n180 10.6151
R1664 B.n180 B.n159 10.6151
R1665 B.n176 B.n159 10.6151
R1666 B.n176 B.n175 10.6151
R1667 B.n175 B.n174 10.6151
R1668 B.n174 B.n161 10.6151
R1669 B.n170 B.n161 10.6151
R1670 B.n170 B.n169 10.6151
R1671 B.n169 B.n168 10.6151
R1672 B.n168 B.n163 10.6151
R1673 B.n164 B.n163 10.6151
R1674 B.n164 B.n0 10.6151
R1675 B.n631 B.n1 10.6151
R1676 B.n631 B.n630 10.6151
R1677 B.n630 B.n629 10.6151
R1678 B.n629 B.n4 10.6151
R1679 B.n625 B.n4 10.6151
R1680 B.n625 B.n624 10.6151
R1681 B.n624 B.n623 10.6151
R1682 B.n623 B.n6 10.6151
R1683 B.n619 B.n6 10.6151
R1684 B.n619 B.n618 10.6151
R1685 B.n618 B.n617 10.6151
R1686 B.n617 B.n8 10.6151
R1687 B.n613 B.n8 10.6151
R1688 B.n613 B.n612 10.6151
R1689 B.n612 B.n611 10.6151
R1690 B.n611 B.n10 10.6151
R1691 B.n607 B.n10 10.6151
R1692 B.n607 B.n606 10.6151
R1693 B.n606 B.n605 10.6151
R1694 B.n605 B.n12 10.6151
R1695 B.n601 B.n12 10.6151
R1696 B.n601 B.n600 10.6151
R1697 B.n523 B.n42 6.5566
R1698 B.n511 B.n510 6.5566
R1699 B.n273 B.n272 6.5566
R1700 B.n288 B.n287 6.5566
R1701 B.n42 B.n38 4.05904
R1702 B.n510 B.n509 4.05904
R1703 B.n272 B.n271 4.05904
R1704 B.n287 B.n121 4.05904
R1705 B.n635 B.n0 2.81026
R1706 B.n635 B.n1 2.81026
R1707 VN VN.t0 258.591
R1708 VN VN.t1 213.167
R1709 VDD2.n157 VDD2.n81 756.745
R1710 VDD2.n76 VDD2.n0 756.745
R1711 VDD2.n158 VDD2.n157 585
R1712 VDD2.n156 VDD2.n155 585
R1713 VDD2.n154 VDD2.n84 585
R1714 VDD2.n88 VDD2.n85 585
R1715 VDD2.n149 VDD2.n148 585
R1716 VDD2.n147 VDD2.n146 585
R1717 VDD2.n90 VDD2.n89 585
R1718 VDD2.n141 VDD2.n140 585
R1719 VDD2.n139 VDD2.n138 585
R1720 VDD2.n94 VDD2.n93 585
R1721 VDD2.n133 VDD2.n132 585
R1722 VDD2.n131 VDD2.n130 585
R1723 VDD2.n98 VDD2.n97 585
R1724 VDD2.n125 VDD2.n124 585
R1725 VDD2.n123 VDD2.n122 585
R1726 VDD2.n102 VDD2.n101 585
R1727 VDD2.n117 VDD2.n116 585
R1728 VDD2.n115 VDD2.n114 585
R1729 VDD2.n106 VDD2.n105 585
R1730 VDD2.n109 VDD2.n108 585
R1731 VDD2.n27 VDD2.n26 585
R1732 VDD2.n24 VDD2.n23 585
R1733 VDD2.n33 VDD2.n32 585
R1734 VDD2.n35 VDD2.n34 585
R1735 VDD2.n20 VDD2.n19 585
R1736 VDD2.n41 VDD2.n40 585
R1737 VDD2.n43 VDD2.n42 585
R1738 VDD2.n16 VDD2.n15 585
R1739 VDD2.n49 VDD2.n48 585
R1740 VDD2.n51 VDD2.n50 585
R1741 VDD2.n12 VDD2.n11 585
R1742 VDD2.n57 VDD2.n56 585
R1743 VDD2.n59 VDD2.n58 585
R1744 VDD2.n8 VDD2.n7 585
R1745 VDD2.n65 VDD2.n64 585
R1746 VDD2.n68 VDD2.n67 585
R1747 VDD2.n66 VDD2.n4 585
R1748 VDD2.n73 VDD2.n3 585
R1749 VDD2.n75 VDD2.n74 585
R1750 VDD2.n77 VDD2.n76 585
R1751 VDD2.t1 VDD2.n107 327.466
R1752 VDD2.t0 VDD2.n25 327.466
R1753 VDD2.n157 VDD2.n156 171.744
R1754 VDD2.n156 VDD2.n84 171.744
R1755 VDD2.n88 VDD2.n84 171.744
R1756 VDD2.n148 VDD2.n88 171.744
R1757 VDD2.n148 VDD2.n147 171.744
R1758 VDD2.n147 VDD2.n89 171.744
R1759 VDD2.n140 VDD2.n89 171.744
R1760 VDD2.n140 VDD2.n139 171.744
R1761 VDD2.n139 VDD2.n93 171.744
R1762 VDD2.n132 VDD2.n93 171.744
R1763 VDD2.n132 VDD2.n131 171.744
R1764 VDD2.n131 VDD2.n97 171.744
R1765 VDD2.n124 VDD2.n97 171.744
R1766 VDD2.n124 VDD2.n123 171.744
R1767 VDD2.n123 VDD2.n101 171.744
R1768 VDD2.n116 VDD2.n101 171.744
R1769 VDD2.n116 VDD2.n115 171.744
R1770 VDD2.n115 VDD2.n105 171.744
R1771 VDD2.n108 VDD2.n105 171.744
R1772 VDD2.n26 VDD2.n23 171.744
R1773 VDD2.n33 VDD2.n23 171.744
R1774 VDD2.n34 VDD2.n33 171.744
R1775 VDD2.n34 VDD2.n19 171.744
R1776 VDD2.n41 VDD2.n19 171.744
R1777 VDD2.n42 VDD2.n41 171.744
R1778 VDD2.n42 VDD2.n15 171.744
R1779 VDD2.n49 VDD2.n15 171.744
R1780 VDD2.n50 VDD2.n49 171.744
R1781 VDD2.n50 VDD2.n11 171.744
R1782 VDD2.n57 VDD2.n11 171.744
R1783 VDD2.n58 VDD2.n57 171.744
R1784 VDD2.n58 VDD2.n7 171.744
R1785 VDD2.n65 VDD2.n7 171.744
R1786 VDD2.n67 VDD2.n65 171.744
R1787 VDD2.n67 VDD2.n66 171.744
R1788 VDD2.n66 VDD2.n3 171.744
R1789 VDD2.n75 VDD2.n3 171.744
R1790 VDD2.n76 VDD2.n75 171.744
R1791 VDD2.n162 VDD2.n80 92.7128
R1792 VDD2.n108 VDD2.t1 85.8723
R1793 VDD2.n26 VDD2.t0 85.8723
R1794 VDD2.n162 VDD2.n161 51.9672
R1795 VDD2.n109 VDD2.n107 16.3895
R1796 VDD2.n27 VDD2.n25 16.3895
R1797 VDD2.n155 VDD2.n154 13.1884
R1798 VDD2.n74 VDD2.n73 13.1884
R1799 VDD2.n158 VDD2.n83 12.8005
R1800 VDD2.n153 VDD2.n85 12.8005
R1801 VDD2.n110 VDD2.n106 12.8005
R1802 VDD2.n28 VDD2.n24 12.8005
R1803 VDD2.n72 VDD2.n4 12.8005
R1804 VDD2.n77 VDD2.n2 12.8005
R1805 VDD2.n159 VDD2.n81 12.0247
R1806 VDD2.n150 VDD2.n149 12.0247
R1807 VDD2.n114 VDD2.n113 12.0247
R1808 VDD2.n32 VDD2.n31 12.0247
R1809 VDD2.n69 VDD2.n68 12.0247
R1810 VDD2.n78 VDD2.n0 12.0247
R1811 VDD2.n146 VDD2.n87 11.249
R1812 VDD2.n117 VDD2.n104 11.249
R1813 VDD2.n35 VDD2.n22 11.249
R1814 VDD2.n64 VDD2.n6 11.249
R1815 VDD2.n145 VDD2.n90 10.4732
R1816 VDD2.n118 VDD2.n102 10.4732
R1817 VDD2.n36 VDD2.n20 10.4732
R1818 VDD2.n63 VDD2.n8 10.4732
R1819 VDD2.n142 VDD2.n141 9.69747
R1820 VDD2.n122 VDD2.n121 9.69747
R1821 VDD2.n40 VDD2.n39 9.69747
R1822 VDD2.n60 VDD2.n59 9.69747
R1823 VDD2.n161 VDD2.n160 9.45567
R1824 VDD2.n80 VDD2.n79 9.45567
R1825 VDD2.n135 VDD2.n134 9.3005
R1826 VDD2.n137 VDD2.n136 9.3005
R1827 VDD2.n92 VDD2.n91 9.3005
R1828 VDD2.n143 VDD2.n142 9.3005
R1829 VDD2.n145 VDD2.n144 9.3005
R1830 VDD2.n87 VDD2.n86 9.3005
R1831 VDD2.n151 VDD2.n150 9.3005
R1832 VDD2.n153 VDD2.n152 9.3005
R1833 VDD2.n160 VDD2.n159 9.3005
R1834 VDD2.n83 VDD2.n82 9.3005
R1835 VDD2.n96 VDD2.n95 9.3005
R1836 VDD2.n129 VDD2.n128 9.3005
R1837 VDD2.n127 VDD2.n126 9.3005
R1838 VDD2.n100 VDD2.n99 9.3005
R1839 VDD2.n121 VDD2.n120 9.3005
R1840 VDD2.n119 VDD2.n118 9.3005
R1841 VDD2.n104 VDD2.n103 9.3005
R1842 VDD2.n113 VDD2.n112 9.3005
R1843 VDD2.n111 VDD2.n110 9.3005
R1844 VDD2.n79 VDD2.n78 9.3005
R1845 VDD2.n2 VDD2.n1 9.3005
R1846 VDD2.n47 VDD2.n46 9.3005
R1847 VDD2.n45 VDD2.n44 9.3005
R1848 VDD2.n18 VDD2.n17 9.3005
R1849 VDD2.n39 VDD2.n38 9.3005
R1850 VDD2.n37 VDD2.n36 9.3005
R1851 VDD2.n22 VDD2.n21 9.3005
R1852 VDD2.n31 VDD2.n30 9.3005
R1853 VDD2.n29 VDD2.n28 9.3005
R1854 VDD2.n14 VDD2.n13 9.3005
R1855 VDD2.n53 VDD2.n52 9.3005
R1856 VDD2.n55 VDD2.n54 9.3005
R1857 VDD2.n10 VDD2.n9 9.3005
R1858 VDD2.n61 VDD2.n60 9.3005
R1859 VDD2.n63 VDD2.n62 9.3005
R1860 VDD2.n6 VDD2.n5 9.3005
R1861 VDD2.n70 VDD2.n69 9.3005
R1862 VDD2.n72 VDD2.n71 9.3005
R1863 VDD2.n138 VDD2.n92 8.92171
R1864 VDD2.n125 VDD2.n100 8.92171
R1865 VDD2.n43 VDD2.n18 8.92171
R1866 VDD2.n56 VDD2.n10 8.92171
R1867 VDD2.n137 VDD2.n94 8.14595
R1868 VDD2.n126 VDD2.n98 8.14595
R1869 VDD2.n44 VDD2.n16 8.14595
R1870 VDD2.n55 VDD2.n12 8.14595
R1871 VDD2.n134 VDD2.n133 7.3702
R1872 VDD2.n130 VDD2.n129 7.3702
R1873 VDD2.n48 VDD2.n47 7.3702
R1874 VDD2.n52 VDD2.n51 7.3702
R1875 VDD2.n133 VDD2.n96 6.59444
R1876 VDD2.n130 VDD2.n96 6.59444
R1877 VDD2.n48 VDD2.n14 6.59444
R1878 VDD2.n51 VDD2.n14 6.59444
R1879 VDD2.n134 VDD2.n94 5.81868
R1880 VDD2.n129 VDD2.n98 5.81868
R1881 VDD2.n47 VDD2.n16 5.81868
R1882 VDD2.n52 VDD2.n12 5.81868
R1883 VDD2.n138 VDD2.n137 5.04292
R1884 VDD2.n126 VDD2.n125 5.04292
R1885 VDD2.n44 VDD2.n43 5.04292
R1886 VDD2.n56 VDD2.n55 5.04292
R1887 VDD2.n141 VDD2.n92 4.26717
R1888 VDD2.n122 VDD2.n100 4.26717
R1889 VDD2.n40 VDD2.n18 4.26717
R1890 VDD2.n59 VDD2.n10 4.26717
R1891 VDD2.n111 VDD2.n107 3.70982
R1892 VDD2.n29 VDD2.n25 3.70982
R1893 VDD2.n142 VDD2.n90 3.49141
R1894 VDD2.n121 VDD2.n102 3.49141
R1895 VDD2.n39 VDD2.n20 3.49141
R1896 VDD2.n60 VDD2.n8 3.49141
R1897 VDD2.n146 VDD2.n145 2.71565
R1898 VDD2.n118 VDD2.n117 2.71565
R1899 VDD2.n36 VDD2.n35 2.71565
R1900 VDD2.n64 VDD2.n63 2.71565
R1901 VDD2.n161 VDD2.n81 1.93989
R1902 VDD2.n149 VDD2.n87 1.93989
R1903 VDD2.n114 VDD2.n104 1.93989
R1904 VDD2.n32 VDD2.n22 1.93989
R1905 VDD2.n68 VDD2.n6 1.93989
R1906 VDD2.n80 VDD2.n0 1.93989
R1907 VDD2.n159 VDD2.n158 1.16414
R1908 VDD2.n150 VDD2.n85 1.16414
R1909 VDD2.n113 VDD2.n106 1.16414
R1910 VDD2.n31 VDD2.n24 1.16414
R1911 VDD2.n69 VDD2.n4 1.16414
R1912 VDD2.n78 VDD2.n77 1.16414
R1913 VDD2 VDD2.n162 0.599638
R1914 VDD2.n155 VDD2.n83 0.388379
R1915 VDD2.n154 VDD2.n153 0.388379
R1916 VDD2.n110 VDD2.n109 0.388379
R1917 VDD2.n28 VDD2.n27 0.388379
R1918 VDD2.n73 VDD2.n72 0.388379
R1919 VDD2.n74 VDD2.n2 0.388379
R1920 VDD2.n160 VDD2.n82 0.155672
R1921 VDD2.n152 VDD2.n82 0.155672
R1922 VDD2.n152 VDD2.n151 0.155672
R1923 VDD2.n151 VDD2.n86 0.155672
R1924 VDD2.n144 VDD2.n86 0.155672
R1925 VDD2.n144 VDD2.n143 0.155672
R1926 VDD2.n143 VDD2.n91 0.155672
R1927 VDD2.n136 VDD2.n91 0.155672
R1928 VDD2.n136 VDD2.n135 0.155672
R1929 VDD2.n135 VDD2.n95 0.155672
R1930 VDD2.n128 VDD2.n95 0.155672
R1931 VDD2.n128 VDD2.n127 0.155672
R1932 VDD2.n127 VDD2.n99 0.155672
R1933 VDD2.n120 VDD2.n99 0.155672
R1934 VDD2.n120 VDD2.n119 0.155672
R1935 VDD2.n119 VDD2.n103 0.155672
R1936 VDD2.n112 VDD2.n103 0.155672
R1937 VDD2.n112 VDD2.n111 0.155672
R1938 VDD2.n30 VDD2.n29 0.155672
R1939 VDD2.n30 VDD2.n21 0.155672
R1940 VDD2.n37 VDD2.n21 0.155672
R1941 VDD2.n38 VDD2.n37 0.155672
R1942 VDD2.n38 VDD2.n17 0.155672
R1943 VDD2.n45 VDD2.n17 0.155672
R1944 VDD2.n46 VDD2.n45 0.155672
R1945 VDD2.n46 VDD2.n13 0.155672
R1946 VDD2.n53 VDD2.n13 0.155672
R1947 VDD2.n54 VDD2.n53 0.155672
R1948 VDD2.n54 VDD2.n9 0.155672
R1949 VDD2.n61 VDD2.n9 0.155672
R1950 VDD2.n62 VDD2.n61 0.155672
R1951 VDD2.n62 VDD2.n5 0.155672
R1952 VDD2.n70 VDD2.n5 0.155672
R1953 VDD2.n71 VDD2.n70 0.155672
R1954 VDD2.n71 VDD2.n1 0.155672
R1955 VDD2.n79 VDD2.n1 0.155672
C0 VDD2 VDD1 0.624898f
C1 VDD1 VP 3.43712f
C2 B VN 1.01528f
C3 VDD2 VN 3.27268f
C4 VP VN 5.77743f
C5 B VTAIL 4.08865f
C6 B w_n1974_n3928# 9.141129f
C7 VDD2 VTAIL 5.83657f
C8 VDD2 w_n1974_n3928# 1.95122f
C9 VP VTAIL 2.78948f
C10 VP w_n1974_n3928# 3.00125f
C11 VDD1 VN 0.148263f
C12 VDD2 B 1.89365f
C13 VDD1 VTAIL 5.79005f
C14 VDD1 w_n1974_n3928# 1.9304f
C15 B VP 1.4255f
C16 VDD2 VP 0.316037f
C17 VN VTAIL 2.7751f
C18 VN w_n1974_n3928# 2.7507f
C19 w_n1974_n3928# VTAIL 3.17782f
C20 VDD1 B 1.86729f
C21 VDD2 VSUBS 0.941421f
C22 VDD1 VSUBS 3.85889f
C23 VTAIL VSUBS 1.05693f
C24 VN VSUBS 8.43357f
C25 VP VSUBS 1.668743f
C26 B VSUBS 3.815037f
C27 w_n1974_n3928# VSUBS 95.1073f
C28 VDD2.n0 VSUBS 0.021586f
C29 VDD2.n1 VSUBS 0.02003f
C30 VDD2.n2 VSUBS 0.010763f
C31 VDD2.n3 VSUBS 0.025441f
C32 VDD2.n4 VSUBS 0.011397f
C33 VDD2.n5 VSUBS 0.02003f
C34 VDD2.n6 VSUBS 0.010763f
C35 VDD2.n7 VSUBS 0.025441f
C36 VDD2.n8 VSUBS 0.011397f
C37 VDD2.n9 VSUBS 0.02003f
C38 VDD2.n10 VSUBS 0.010763f
C39 VDD2.n11 VSUBS 0.025441f
C40 VDD2.n12 VSUBS 0.011397f
C41 VDD2.n13 VSUBS 0.02003f
C42 VDD2.n14 VSUBS 0.010763f
C43 VDD2.n15 VSUBS 0.025441f
C44 VDD2.n16 VSUBS 0.011397f
C45 VDD2.n17 VSUBS 0.02003f
C46 VDD2.n18 VSUBS 0.010763f
C47 VDD2.n19 VSUBS 0.025441f
C48 VDD2.n20 VSUBS 0.011397f
C49 VDD2.n21 VSUBS 0.02003f
C50 VDD2.n22 VSUBS 0.010763f
C51 VDD2.n23 VSUBS 0.025441f
C52 VDD2.n24 VSUBS 0.011397f
C53 VDD2.n25 VSUBS 0.140014f
C54 VDD2.t0 VSUBS 0.054453f
C55 VDD2.n26 VSUBS 0.01908f
C56 VDD2.n27 VSUBS 0.016184f
C57 VDD2.n28 VSUBS 0.010763f
C58 VDD2.n29 VSUBS 1.26078f
C59 VDD2.n30 VSUBS 0.02003f
C60 VDD2.n31 VSUBS 0.010763f
C61 VDD2.n32 VSUBS 0.011397f
C62 VDD2.n33 VSUBS 0.025441f
C63 VDD2.n34 VSUBS 0.025441f
C64 VDD2.n35 VSUBS 0.011397f
C65 VDD2.n36 VSUBS 0.010763f
C66 VDD2.n37 VSUBS 0.02003f
C67 VDD2.n38 VSUBS 0.02003f
C68 VDD2.n39 VSUBS 0.010763f
C69 VDD2.n40 VSUBS 0.011397f
C70 VDD2.n41 VSUBS 0.025441f
C71 VDD2.n42 VSUBS 0.025441f
C72 VDD2.n43 VSUBS 0.011397f
C73 VDD2.n44 VSUBS 0.010763f
C74 VDD2.n45 VSUBS 0.02003f
C75 VDD2.n46 VSUBS 0.02003f
C76 VDD2.n47 VSUBS 0.010763f
C77 VDD2.n48 VSUBS 0.011397f
C78 VDD2.n49 VSUBS 0.025441f
C79 VDD2.n50 VSUBS 0.025441f
C80 VDD2.n51 VSUBS 0.011397f
C81 VDD2.n52 VSUBS 0.010763f
C82 VDD2.n53 VSUBS 0.02003f
C83 VDD2.n54 VSUBS 0.02003f
C84 VDD2.n55 VSUBS 0.010763f
C85 VDD2.n56 VSUBS 0.011397f
C86 VDD2.n57 VSUBS 0.025441f
C87 VDD2.n58 VSUBS 0.025441f
C88 VDD2.n59 VSUBS 0.011397f
C89 VDD2.n60 VSUBS 0.010763f
C90 VDD2.n61 VSUBS 0.02003f
C91 VDD2.n62 VSUBS 0.02003f
C92 VDD2.n63 VSUBS 0.010763f
C93 VDD2.n64 VSUBS 0.011397f
C94 VDD2.n65 VSUBS 0.025441f
C95 VDD2.n66 VSUBS 0.025441f
C96 VDD2.n67 VSUBS 0.025441f
C97 VDD2.n68 VSUBS 0.011397f
C98 VDD2.n69 VSUBS 0.010763f
C99 VDD2.n70 VSUBS 0.02003f
C100 VDD2.n71 VSUBS 0.02003f
C101 VDD2.n72 VSUBS 0.010763f
C102 VDD2.n73 VSUBS 0.01108f
C103 VDD2.n74 VSUBS 0.01108f
C104 VDD2.n75 VSUBS 0.025441f
C105 VDD2.n76 VSUBS 0.060147f
C106 VDD2.n77 VSUBS 0.011397f
C107 VDD2.n78 VSUBS 0.010763f
C108 VDD2.n79 VSUBS 0.050677f
C109 VDD2.n80 VSUBS 0.627992f
C110 VDD2.n81 VSUBS 0.021586f
C111 VDD2.n82 VSUBS 0.02003f
C112 VDD2.n83 VSUBS 0.010763f
C113 VDD2.n84 VSUBS 0.025441f
C114 VDD2.n85 VSUBS 0.011397f
C115 VDD2.n86 VSUBS 0.02003f
C116 VDD2.n87 VSUBS 0.010763f
C117 VDD2.n88 VSUBS 0.025441f
C118 VDD2.n89 VSUBS 0.025441f
C119 VDD2.n90 VSUBS 0.011397f
C120 VDD2.n91 VSUBS 0.02003f
C121 VDD2.n92 VSUBS 0.010763f
C122 VDD2.n93 VSUBS 0.025441f
C123 VDD2.n94 VSUBS 0.011397f
C124 VDD2.n95 VSUBS 0.02003f
C125 VDD2.n96 VSUBS 0.010763f
C126 VDD2.n97 VSUBS 0.025441f
C127 VDD2.n98 VSUBS 0.011397f
C128 VDD2.n99 VSUBS 0.02003f
C129 VDD2.n100 VSUBS 0.010763f
C130 VDD2.n101 VSUBS 0.025441f
C131 VDD2.n102 VSUBS 0.011397f
C132 VDD2.n103 VSUBS 0.02003f
C133 VDD2.n104 VSUBS 0.010763f
C134 VDD2.n105 VSUBS 0.025441f
C135 VDD2.n106 VSUBS 0.011397f
C136 VDD2.n107 VSUBS 0.140014f
C137 VDD2.t1 VSUBS 0.054453f
C138 VDD2.n108 VSUBS 0.01908f
C139 VDD2.n109 VSUBS 0.016184f
C140 VDD2.n110 VSUBS 0.010763f
C141 VDD2.n111 VSUBS 1.26078f
C142 VDD2.n112 VSUBS 0.02003f
C143 VDD2.n113 VSUBS 0.010763f
C144 VDD2.n114 VSUBS 0.011397f
C145 VDD2.n115 VSUBS 0.025441f
C146 VDD2.n116 VSUBS 0.025441f
C147 VDD2.n117 VSUBS 0.011397f
C148 VDD2.n118 VSUBS 0.010763f
C149 VDD2.n119 VSUBS 0.02003f
C150 VDD2.n120 VSUBS 0.02003f
C151 VDD2.n121 VSUBS 0.010763f
C152 VDD2.n122 VSUBS 0.011397f
C153 VDD2.n123 VSUBS 0.025441f
C154 VDD2.n124 VSUBS 0.025441f
C155 VDD2.n125 VSUBS 0.011397f
C156 VDD2.n126 VSUBS 0.010763f
C157 VDD2.n127 VSUBS 0.02003f
C158 VDD2.n128 VSUBS 0.02003f
C159 VDD2.n129 VSUBS 0.010763f
C160 VDD2.n130 VSUBS 0.011397f
C161 VDD2.n131 VSUBS 0.025441f
C162 VDD2.n132 VSUBS 0.025441f
C163 VDD2.n133 VSUBS 0.011397f
C164 VDD2.n134 VSUBS 0.010763f
C165 VDD2.n135 VSUBS 0.02003f
C166 VDD2.n136 VSUBS 0.02003f
C167 VDD2.n137 VSUBS 0.010763f
C168 VDD2.n138 VSUBS 0.011397f
C169 VDD2.n139 VSUBS 0.025441f
C170 VDD2.n140 VSUBS 0.025441f
C171 VDD2.n141 VSUBS 0.011397f
C172 VDD2.n142 VSUBS 0.010763f
C173 VDD2.n143 VSUBS 0.02003f
C174 VDD2.n144 VSUBS 0.02003f
C175 VDD2.n145 VSUBS 0.010763f
C176 VDD2.n146 VSUBS 0.011397f
C177 VDD2.n147 VSUBS 0.025441f
C178 VDD2.n148 VSUBS 0.025441f
C179 VDD2.n149 VSUBS 0.011397f
C180 VDD2.n150 VSUBS 0.010763f
C181 VDD2.n151 VSUBS 0.02003f
C182 VDD2.n152 VSUBS 0.02003f
C183 VDD2.n153 VSUBS 0.010763f
C184 VDD2.n154 VSUBS 0.01108f
C185 VDD2.n155 VSUBS 0.01108f
C186 VDD2.n156 VSUBS 0.025441f
C187 VDD2.n157 VSUBS 0.060147f
C188 VDD2.n158 VSUBS 0.011397f
C189 VDD2.n159 VSUBS 0.010763f
C190 VDD2.n160 VSUBS 0.050677f
C191 VDD2.n161 VSUBS 0.044112f
C192 VDD2.n162 VSUBS 2.63531f
C193 VN.t1 VSUBS 4.02221f
C194 VN.t0 VSUBS 4.60388f
C195 B.n0 VSUBS 0.003739f
C196 B.n1 VSUBS 0.003739f
C197 B.n2 VSUBS 0.005913f
C198 B.n3 VSUBS 0.005913f
C199 B.n4 VSUBS 0.005913f
C200 B.n5 VSUBS 0.005913f
C201 B.n6 VSUBS 0.005913f
C202 B.n7 VSUBS 0.005913f
C203 B.n8 VSUBS 0.005913f
C204 B.n9 VSUBS 0.005913f
C205 B.n10 VSUBS 0.005913f
C206 B.n11 VSUBS 0.005913f
C207 B.n12 VSUBS 0.005913f
C208 B.n13 VSUBS 0.013647f
C209 B.n14 VSUBS 0.005913f
C210 B.n15 VSUBS 0.005913f
C211 B.n16 VSUBS 0.005913f
C212 B.n17 VSUBS 0.005913f
C213 B.n18 VSUBS 0.005913f
C214 B.n19 VSUBS 0.005913f
C215 B.n20 VSUBS 0.005913f
C216 B.n21 VSUBS 0.005913f
C217 B.n22 VSUBS 0.005913f
C218 B.n23 VSUBS 0.005913f
C219 B.n24 VSUBS 0.005913f
C220 B.n25 VSUBS 0.005913f
C221 B.n26 VSUBS 0.005913f
C222 B.n27 VSUBS 0.005913f
C223 B.n28 VSUBS 0.005913f
C224 B.n29 VSUBS 0.005913f
C225 B.n30 VSUBS 0.005913f
C226 B.n31 VSUBS 0.005913f
C227 B.n32 VSUBS 0.005913f
C228 B.n33 VSUBS 0.005913f
C229 B.n34 VSUBS 0.005913f
C230 B.n35 VSUBS 0.005913f
C231 B.n36 VSUBS 0.005913f
C232 B.n37 VSUBS 0.005913f
C233 B.n38 VSUBS 0.004087f
C234 B.n39 VSUBS 0.005913f
C235 B.t8 VSUBS 0.232274f
C236 B.t7 VSUBS 0.256302f
C237 B.t6 VSUBS 1.20916f
C238 B.n40 VSUBS 0.391962f
C239 B.n41 VSUBS 0.242777f
C240 B.n42 VSUBS 0.013701f
C241 B.n43 VSUBS 0.005913f
C242 B.n44 VSUBS 0.005913f
C243 B.n45 VSUBS 0.005913f
C244 B.n46 VSUBS 0.005913f
C245 B.t11 VSUBS 0.232277f
C246 B.t10 VSUBS 0.256305f
C247 B.t9 VSUBS 1.20916f
C248 B.n47 VSUBS 0.391959f
C249 B.n48 VSUBS 0.242774f
C250 B.n49 VSUBS 0.005913f
C251 B.n50 VSUBS 0.005913f
C252 B.n51 VSUBS 0.005913f
C253 B.n52 VSUBS 0.005913f
C254 B.n53 VSUBS 0.005913f
C255 B.n54 VSUBS 0.005913f
C256 B.n55 VSUBS 0.005913f
C257 B.n56 VSUBS 0.005913f
C258 B.n57 VSUBS 0.005913f
C259 B.n58 VSUBS 0.005913f
C260 B.n59 VSUBS 0.005913f
C261 B.n60 VSUBS 0.005913f
C262 B.n61 VSUBS 0.005913f
C263 B.n62 VSUBS 0.005913f
C264 B.n63 VSUBS 0.005913f
C265 B.n64 VSUBS 0.005913f
C266 B.n65 VSUBS 0.005913f
C267 B.n66 VSUBS 0.005913f
C268 B.n67 VSUBS 0.005913f
C269 B.n68 VSUBS 0.005913f
C270 B.n69 VSUBS 0.005913f
C271 B.n70 VSUBS 0.005913f
C272 B.n71 VSUBS 0.005913f
C273 B.n72 VSUBS 0.005913f
C274 B.n73 VSUBS 0.014347f
C275 B.n74 VSUBS 0.005913f
C276 B.n75 VSUBS 0.005913f
C277 B.n76 VSUBS 0.005913f
C278 B.n77 VSUBS 0.005913f
C279 B.n78 VSUBS 0.005913f
C280 B.n79 VSUBS 0.005913f
C281 B.n80 VSUBS 0.005913f
C282 B.n81 VSUBS 0.005913f
C283 B.n82 VSUBS 0.005913f
C284 B.n83 VSUBS 0.005913f
C285 B.n84 VSUBS 0.005913f
C286 B.n85 VSUBS 0.005913f
C287 B.n86 VSUBS 0.005913f
C288 B.n87 VSUBS 0.005913f
C289 B.n88 VSUBS 0.005913f
C290 B.n89 VSUBS 0.005913f
C291 B.n90 VSUBS 0.005913f
C292 B.n91 VSUBS 0.005913f
C293 B.n92 VSUBS 0.005913f
C294 B.n93 VSUBS 0.005913f
C295 B.n94 VSUBS 0.005913f
C296 B.n95 VSUBS 0.005913f
C297 B.n96 VSUBS 0.013647f
C298 B.n97 VSUBS 0.005913f
C299 B.n98 VSUBS 0.005913f
C300 B.n99 VSUBS 0.005913f
C301 B.n100 VSUBS 0.005913f
C302 B.n101 VSUBS 0.005913f
C303 B.n102 VSUBS 0.005913f
C304 B.n103 VSUBS 0.005913f
C305 B.n104 VSUBS 0.005913f
C306 B.n105 VSUBS 0.005913f
C307 B.n106 VSUBS 0.005913f
C308 B.n107 VSUBS 0.005913f
C309 B.n108 VSUBS 0.005913f
C310 B.n109 VSUBS 0.005913f
C311 B.n110 VSUBS 0.005913f
C312 B.n111 VSUBS 0.005913f
C313 B.n112 VSUBS 0.005913f
C314 B.n113 VSUBS 0.005913f
C315 B.n114 VSUBS 0.005913f
C316 B.n115 VSUBS 0.005913f
C317 B.n116 VSUBS 0.005913f
C318 B.n117 VSUBS 0.005913f
C319 B.n118 VSUBS 0.005913f
C320 B.n119 VSUBS 0.005913f
C321 B.n120 VSUBS 0.005913f
C322 B.n121 VSUBS 0.004087f
C323 B.n122 VSUBS 0.005913f
C324 B.n123 VSUBS 0.005913f
C325 B.n124 VSUBS 0.005913f
C326 B.n125 VSUBS 0.005913f
C327 B.n126 VSUBS 0.005913f
C328 B.t4 VSUBS 0.232274f
C329 B.t5 VSUBS 0.256302f
C330 B.t3 VSUBS 1.20916f
C331 B.n127 VSUBS 0.391962f
C332 B.n128 VSUBS 0.242777f
C333 B.n129 VSUBS 0.005913f
C334 B.n130 VSUBS 0.005913f
C335 B.n131 VSUBS 0.005913f
C336 B.n132 VSUBS 0.005913f
C337 B.n133 VSUBS 0.005913f
C338 B.n134 VSUBS 0.005913f
C339 B.n135 VSUBS 0.005913f
C340 B.n136 VSUBS 0.005913f
C341 B.n137 VSUBS 0.005913f
C342 B.n138 VSUBS 0.005913f
C343 B.n139 VSUBS 0.005913f
C344 B.n140 VSUBS 0.005913f
C345 B.n141 VSUBS 0.005913f
C346 B.n142 VSUBS 0.005913f
C347 B.n143 VSUBS 0.005913f
C348 B.n144 VSUBS 0.005913f
C349 B.n145 VSUBS 0.005913f
C350 B.n146 VSUBS 0.005913f
C351 B.n147 VSUBS 0.005913f
C352 B.n148 VSUBS 0.005913f
C353 B.n149 VSUBS 0.005913f
C354 B.n150 VSUBS 0.005913f
C355 B.n151 VSUBS 0.005913f
C356 B.n152 VSUBS 0.005913f
C357 B.n153 VSUBS 0.013647f
C358 B.n154 VSUBS 0.005913f
C359 B.n155 VSUBS 0.005913f
C360 B.n156 VSUBS 0.005913f
C361 B.n157 VSUBS 0.005913f
C362 B.n158 VSUBS 0.005913f
C363 B.n159 VSUBS 0.005913f
C364 B.n160 VSUBS 0.005913f
C365 B.n161 VSUBS 0.005913f
C366 B.n162 VSUBS 0.005913f
C367 B.n163 VSUBS 0.005913f
C368 B.n164 VSUBS 0.005913f
C369 B.n165 VSUBS 0.005913f
C370 B.n166 VSUBS 0.005913f
C371 B.n167 VSUBS 0.005913f
C372 B.n168 VSUBS 0.005913f
C373 B.n169 VSUBS 0.005913f
C374 B.n170 VSUBS 0.005913f
C375 B.n171 VSUBS 0.005913f
C376 B.n172 VSUBS 0.005913f
C377 B.n173 VSUBS 0.005913f
C378 B.n174 VSUBS 0.005913f
C379 B.n175 VSUBS 0.005913f
C380 B.n176 VSUBS 0.005913f
C381 B.n177 VSUBS 0.005913f
C382 B.n178 VSUBS 0.005913f
C383 B.n179 VSUBS 0.005913f
C384 B.n180 VSUBS 0.005913f
C385 B.n181 VSUBS 0.005913f
C386 B.n182 VSUBS 0.005913f
C387 B.n183 VSUBS 0.005913f
C388 B.n184 VSUBS 0.005913f
C389 B.n185 VSUBS 0.005913f
C390 B.n186 VSUBS 0.005913f
C391 B.n187 VSUBS 0.005913f
C392 B.n188 VSUBS 0.005913f
C393 B.n189 VSUBS 0.005913f
C394 B.n190 VSUBS 0.005913f
C395 B.n191 VSUBS 0.005913f
C396 B.n192 VSUBS 0.005913f
C397 B.n193 VSUBS 0.005913f
C398 B.n194 VSUBS 0.005913f
C399 B.n195 VSUBS 0.005913f
C400 B.n196 VSUBS 0.013647f
C401 B.n197 VSUBS 0.014006f
C402 B.n198 VSUBS 0.014006f
C403 B.n199 VSUBS 0.005913f
C404 B.n200 VSUBS 0.005913f
C405 B.n201 VSUBS 0.005913f
C406 B.n202 VSUBS 0.005913f
C407 B.n203 VSUBS 0.005913f
C408 B.n204 VSUBS 0.005913f
C409 B.n205 VSUBS 0.005913f
C410 B.n206 VSUBS 0.005913f
C411 B.n207 VSUBS 0.005913f
C412 B.n208 VSUBS 0.005913f
C413 B.n209 VSUBS 0.005913f
C414 B.n210 VSUBS 0.005913f
C415 B.n211 VSUBS 0.005913f
C416 B.n212 VSUBS 0.005913f
C417 B.n213 VSUBS 0.005913f
C418 B.n214 VSUBS 0.005913f
C419 B.n215 VSUBS 0.005913f
C420 B.n216 VSUBS 0.005913f
C421 B.n217 VSUBS 0.005913f
C422 B.n218 VSUBS 0.005913f
C423 B.n219 VSUBS 0.005913f
C424 B.n220 VSUBS 0.005913f
C425 B.n221 VSUBS 0.005913f
C426 B.n222 VSUBS 0.005913f
C427 B.n223 VSUBS 0.005913f
C428 B.n224 VSUBS 0.005913f
C429 B.n225 VSUBS 0.005913f
C430 B.n226 VSUBS 0.005913f
C431 B.n227 VSUBS 0.005913f
C432 B.n228 VSUBS 0.005913f
C433 B.n229 VSUBS 0.005913f
C434 B.n230 VSUBS 0.005913f
C435 B.n231 VSUBS 0.005913f
C436 B.n232 VSUBS 0.005913f
C437 B.n233 VSUBS 0.005913f
C438 B.n234 VSUBS 0.005913f
C439 B.n235 VSUBS 0.005913f
C440 B.n236 VSUBS 0.005913f
C441 B.n237 VSUBS 0.005913f
C442 B.n238 VSUBS 0.005913f
C443 B.n239 VSUBS 0.005913f
C444 B.n240 VSUBS 0.005913f
C445 B.n241 VSUBS 0.005913f
C446 B.n242 VSUBS 0.005913f
C447 B.n243 VSUBS 0.005913f
C448 B.n244 VSUBS 0.005913f
C449 B.n245 VSUBS 0.005913f
C450 B.n246 VSUBS 0.005913f
C451 B.n247 VSUBS 0.005913f
C452 B.n248 VSUBS 0.005913f
C453 B.n249 VSUBS 0.005913f
C454 B.n250 VSUBS 0.005913f
C455 B.n251 VSUBS 0.005913f
C456 B.n252 VSUBS 0.005913f
C457 B.n253 VSUBS 0.005913f
C458 B.n254 VSUBS 0.005913f
C459 B.n255 VSUBS 0.005913f
C460 B.n256 VSUBS 0.005913f
C461 B.n257 VSUBS 0.005913f
C462 B.n258 VSUBS 0.005913f
C463 B.n259 VSUBS 0.005913f
C464 B.n260 VSUBS 0.005913f
C465 B.n261 VSUBS 0.005913f
C466 B.n262 VSUBS 0.005913f
C467 B.n263 VSUBS 0.005913f
C468 B.n264 VSUBS 0.005913f
C469 B.n265 VSUBS 0.005913f
C470 B.n266 VSUBS 0.005913f
C471 B.n267 VSUBS 0.005913f
C472 B.n268 VSUBS 0.005913f
C473 B.n269 VSUBS 0.005913f
C474 B.n270 VSUBS 0.005913f
C475 B.n271 VSUBS 0.004087f
C476 B.n272 VSUBS 0.013701f
C477 B.n273 VSUBS 0.004783f
C478 B.n274 VSUBS 0.005913f
C479 B.n275 VSUBS 0.005913f
C480 B.n276 VSUBS 0.005913f
C481 B.n277 VSUBS 0.005913f
C482 B.n278 VSUBS 0.005913f
C483 B.n279 VSUBS 0.005913f
C484 B.n280 VSUBS 0.005913f
C485 B.n281 VSUBS 0.005913f
C486 B.n282 VSUBS 0.005913f
C487 B.n283 VSUBS 0.005913f
C488 B.n284 VSUBS 0.005913f
C489 B.t1 VSUBS 0.232277f
C490 B.t2 VSUBS 0.256305f
C491 B.t0 VSUBS 1.20916f
C492 B.n285 VSUBS 0.391959f
C493 B.n286 VSUBS 0.242774f
C494 B.n287 VSUBS 0.013701f
C495 B.n288 VSUBS 0.004783f
C496 B.n289 VSUBS 0.005913f
C497 B.n290 VSUBS 0.005913f
C498 B.n291 VSUBS 0.005913f
C499 B.n292 VSUBS 0.005913f
C500 B.n293 VSUBS 0.005913f
C501 B.n294 VSUBS 0.005913f
C502 B.n295 VSUBS 0.005913f
C503 B.n296 VSUBS 0.005913f
C504 B.n297 VSUBS 0.005913f
C505 B.n298 VSUBS 0.005913f
C506 B.n299 VSUBS 0.005913f
C507 B.n300 VSUBS 0.005913f
C508 B.n301 VSUBS 0.005913f
C509 B.n302 VSUBS 0.005913f
C510 B.n303 VSUBS 0.005913f
C511 B.n304 VSUBS 0.005913f
C512 B.n305 VSUBS 0.005913f
C513 B.n306 VSUBS 0.005913f
C514 B.n307 VSUBS 0.005913f
C515 B.n308 VSUBS 0.005913f
C516 B.n309 VSUBS 0.005913f
C517 B.n310 VSUBS 0.005913f
C518 B.n311 VSUBS 0.005913f
C519 B.n312 VSUBS 0.005913f
C520 B.n313 VSUBS 0.005913f
C521 B.n314 VSUBS 0.005913f
C522 B.n315 VSUBS 0.005913f
C523 B.n316 VSUBS 0.005913f
C524 B.n317 VSUBS 0.005913f
C525 B.n318 VSUBS 0.005913f
C526 B.n319 VSUBS 0.005913f
C527 B.n320 VSUBS 0.005913f
C528 B.n321 VSUBS 0.005913f
C529 B.n322 VSUBS 0.005913f
C530 B.n323 VSUBS 0.005913f
C531 B.n324 VSUBS 0.005913f
C532 B.n325 VSUBS 0.005913f
C533 B.n326 VSUBS 0.005913f
C534 B.n327 VSUBS 0.005913f
C535 B.n328 VSUBS 0.005913f
C536 B.n329 VSUBS 0.005913f
C537 B.n330 VSUBS 0.005913f
C538 B.n331 VSUBS 0.005913f
C539 B.n332 VSUBS 0.005913f
C540 B.n333 VSUBS 0.005913f
C541 B.n334 VSUBS 0.005913f
C542 B.n335 VSUBS 0.005913f
C543 B.n336 VSUBS 0.005913f
C544 B.n337 VSUBS 0.005913f
C545 B.n338 VSUBS 0.005913f
C546 B.n339 VSUBS 0.005913f
C547 B.n340 VSUBS 0.005913f
C548 B.n341 VSUBS 0.005913f
C549 B.n342 VSUBS 0.005913f
C550 B.n343 VSUBS 0.005913f
C551 B.n344 VSUBS 0.005913f
C552 B.n345 VSUBS 0.005913f
C553 B.n346 VSUBS 0.005913f
C554 B.n347 VSUBS 0.005913f
C555 B.n348 VSUBS 0.005913f
C556 B.n349 VSUBS 0.005913f
C557 B.n350 VSUBS 0.005913f
C558 B.n351 VSUBS 0.005913f
C559 B.n352 VSUBS 0.005913f
C560 B.n353 VSUBS 0.005913f
C561 B.n354 VSUBS 0.005913f
C562 B.n355 VSUBS 0.005913f
C563 B.n356 VSUBS 0.005913f
C564 B.n357 VSUBS 0.005913f
C565 B.n358 VSUBS 0.005913f
C566 B.n359 VSUBS 0.005913f
C567 B.n360 VSUBS 0.005913f
C568 B.n361 VSUBS 0.005913f
C569 B.n362 VSUBS 0.005913f
C570 B.n363 VSUBS 0.014006f
C571 B.n364 VSUBS 0.014006f
C572 B.n365 VSUBS 0.013647f
C573 B.n366 VSUBS 0.005913f
C574 B.n367 VSUBS 0.005913f
C575 B.n368 VSUBS 0.005913f
C576 B.n369 VSUBS 0.005913f
C577 B.n370 VSUBS 0.005913f
C578 B.n371 VSUBS 0.005913f
C579 B.n372 VSUBS 0.005913f
C580 B.n373 VSUBS 0.005913f
C581 B.n374 VSUBS 0.005913f
C582 B.n375 VSUBS 0.005913f
C583 B.n376 VSUBS 0.005913f
C584 B.n377 VSUBS 0.005913f
C585 B.n378 VSUBS 0.005913f
C586 B.n379 VSUBS 0.005913f
C587 B.n380 VSUBS 0.005913f
C588 B.n381 VSUBS 0.005913f
C589 B.n382 VSUBS 0.005913f
C590 B.n383 VSUBS 0.005913f
C591 B.n384 VSUBS 0.005913f
C592 B.n385 VSUBS 0.005913f
C593 B.n386 VSUBS 0.005913f
C594 B.n387 VSUBS 0.005913f
C595 B.n388 VSUBS 0.005913f
C596 B.n389 VSUBS 0.005913f
C597 B.n390 VSUBS 0.005913f
C598 B.n391 VSUBS 0.005913f
C599 B.n392 VSUBS 0.005913f
C600 B.n393 VSUBS 0.005913f
C601 B.n394 VSUBS 0.005913f
C602 B.n395 VSUBS 0.005913f
C603 B.n396 VSUBS 0.005913f
C604 B.n397 VSUBS 0.005913f
C605 B.n398 VSUBS 0.005913f
C606 B.n399 VSUBS 0.005913f
C607 B.n400 VSUBS 0.005913f
C608 B.n401 VSUBS 0.005913f
C609 B.n402 VSUBS 0.005913f
C610 B.n403 VSUBS 0.005913f
C611 B.n404 VSUBS 0.005913f
C612 B.n405 VSUBS 0.005913f
C613 B.n406 VSUBS 0.005913f
C614 B.n407 VSUBS 0.005913f
C615 B.n408 VSUBS 0.005913f
C616 B.n409 VSUBS 0.005913f
C617 B.n410 VSUBS 0.005913f
C618 B.n411 VSUBS 0.005913f
C619 B.n412 VSUBS 0.005913f
C620 B.n413 VSUBS 0.005913f
C621 B.n414 VSUBS 0.005913f
C622 B.n415 VSUBS 0.005913f
C623 B.n416 VSUBS 0.005913f
C624 B.n417 VSUBS 0.005913f
C625 B.n418 VSUBS 0.005913f
C626 B.n419 VSUBS 0.005913f
C627 B.n420 VSUBS 0.005913f
C628 B.n421 VSUBS 0.005913f
C629 B.n422 VSUBS 0.005913f
C630 B.n423 VSUBS 0.005913f
C631 B.n424 VSUBS 0.005913f
C632 B.n425 VSUBS 0.005913f
C633 B.n426 VSUBS 0.005913f
C634 B.n427 VSUBS 0.005913f
C635 B.n428 VSUBS 0.005913f
C636 B.n429 VSUBS 0.005913f
C637 B.n430 VSUBS 0.005913f
C638 B.n431 VSUBS 0.005913f
C639 B.n432 VSUBS 0.005913f
C640 B.n433 VSUBS 0.005913f
C641 B.n434 VSUBS 0.013647f
C642 B.n435 VSUBS 0.014006f
C643 B.n436 VSUBS 0.013306f
C644 B.n437 VSUBS 0.005913f
C645 B.n438 VSUBS 0.005913f
C646 B.n439 VSUBS 0.005913f
C647 B.n440 VSUBS 0.005913f
C648 B.n441 VSUBS 0.005913f
C649 B.n442 VSUBS 0.005913f
C650 B.n443 VSUBS 0.005913f
C651 B.n444 VSUBS 0.005913f
C652 B.n445 VSUBS 0.005913f
C653 B.n446 VSUBS 0.005913f
C654 B.n447 VSUBS 0.005913f
C655 B.n448 VSUBS 0.005913f
C656 B.n449 VSUBS 0.005913f
C657 B.n450 VSUBS 0.005913f
C658 B.n451 VSUBS 0.005913f
C659 B.n452 VSUBS 0.005913f
C660 B.n453 VSUBS 0.005913f
C661 B.n454 VSUBS 0.005913f
C662 B.n455 VSUBS 0.005913f
C663 B.n456 VSUBS 0.005913f
C664 B.n457 VSUBS 0.005913f
C665 B.n458 VSUBS 0.005913f
C666 B.n459 VSUBS 0.005913f
C667 B.n460 VSUBS 0.005913f
C668 B.n461 VSUBS 0.005913f
C669 B.n462 VSUBS 0.005913f
C670 B.n463 VSUBS 0.005913f
C671 B.n464 VSUBS 0.005913f
C672 B.n465 VSUBS 0.005913f
C673 B.n466 VSUBS 0.005913f
C674 B.n467 VSUBS 0.005913f
C675 B.n468 VSUBS 0.005913f
C676 B.n469 VSUBS 0.005913f
C677 B.n470 VSUBS 0.005913f
C678 B.n471 VSUBS 0.005913f
C679 B.n472 VSUBS 0.005913f
C680 B.n473 VSUBS 0.005913f
C681 B.n474 VSUBS 0.005913f
C682 B.n475 VSUBS 0.005913f
C683 B.n476 VSUBS 0.005913f
C684 B.n477 VSUBS 0.005913f
C685 B.n478 VSUBS 0.005913f
C686 B.n479 VSUBS 0.005913f
C687 B.n480 VSUBS 0.005913f
C688 B.n481 VSUBS 0.005913f
C689 B.n482 VSUBS 0.005913f
C690 B.n483 VSUBS 0.005913f
C691 B.n484 VSUBS 0.005913f
C692 B.n485 VSUBS 0.005913f
C693 B.n486 VSUBS 0.005913f
C694 B.n487 VSUBS 0.005913f
C695 B.n488 VSUBS 0.005913f
C696 B.n489 VSUBS 0.005913f
C697 B.n490 VSUBS 0.005913f
C698 B.n491 VSUBS 0.005913f
C699 B.n492 VSUBS 0.005913f
C700 B.n493 VSUBS 0.005913f
C701 B.n494 VSUBS 0.005913f
C702 B.n495 VSUBS 0.005913f
C703 B.n496 VSUBS 0.005913f
C704 B.n497 VSUBS 0.005913f
C705 B.n498 VSUBS 0.005913f
C706 B.n499 VSUBS 0.005913f
C707 B.n500 VSUBS 0.005913f
C708 B.n501 VSUBS 0.005913f
C709 B.n502 VSUBS 0.005913f
C710 B.n503 VSUBS 0.005913f
C711 B.n504 VSUBS 0.005913f
C712 B.n505 VSUBS 0.005913f
C713 B.n506 VSUBS 0.005913f
C714 B.n507 VSUBS 0.005913f
C715 B.n508 VSUBS 0.005913f
C716 B.n509 VSUBS 0.004087f
C717 B.n510 VSUBS 0.013701f
C718 B.n511 VSUBS 0.004783f
C719 B.n512 VSUBS 0.005913f
C720 B.n513 VSUBS 0.005913f
C721 B.n514 VSUBS 0.005913f
C722 B.n515 VSUBS 0.005913f
C723 B.n516 VSUBS 0.005913f
C724 B.n517 VSUBS 0.005913f
C725 B.n518 VSUBS 0.005913f
C726 B.n519 VSUBS 0.005913f
C727 B.n520 VSUBS 0.005913f
C728 B.n521 VSUBS 0.005913f
C729 B.n522 VSUBS 0.005913f
C730 B.n523 VSUBS 0.004783f
C731 B.n524 VSUBS 0.005913f
C732 B.n525 VSUBS 0.005913f
C733 B.n526 VSUBS 0.005913f
C734 B.n527 VSUBS 0.005913f
C735 B.n528 VSUBS 0.005913f
C736 B.n529 VSUBS 0.005913f
C737 B.n530 VSUBS 0.005913f
C738 B.n531 VSUBS 0.005913f
C739 B.n532 VSUBS 0.005913f
C740 B.n533 VSUBS 0.005913f
C741 B.n534 VSUBS 0.005913f
C742 B.n535 VSUBS 0.005913f
C743 B.n536 VSUBS 0.005913f
C744 B.n537 VSUBS 0.005913f
C745 B.n538 VSUBS 0.005913f
C746 B.n539 VSUBS 0.005913f
C747 B.n540 VSUBS 0.005913f
C748 B.n541 VSUBS 0.005913f
C749 B.n542 VSUBS 0.005913f
C750 B.n543 VSUBS 0.005913f
C751 B.n544 VSUBS 0.005913f
C752 B.n545 VSUBS 0.005913f
C753 B.n546 VSUBS 0.005913f
C754 B.n547 VSUBS 0.005913f
C755 B.n548 VSUBS 0.005913f
C756 B.n549 VSUBS 0.005913f
C757 B.n550 VSUBS 0.005913f
C758 B.n551 VSUBS 0.005913f
C759 B.n552 VSUBS 0.005913f
C760 B.n553 VSUBS 0.005913f
C761 B.n554 VSUBS 0.005913f
C762 B.n555 VSUBS 0.005913f
C763 B.n556 VSUBS 0.005913f
C764 B.n557 VSUBS 0.005913f
C765 B.n558 VSUBS 0.005913f
C766 B.n559 VSUBS 0.005913f
C767 B.n560 VSUBS 0.005913f
C768 B.n561 VSUBS 0.005913f
C769 B.n562 VSUBS 0.005913f
C770 B.n563 VSUBS 0.005913f
C771 B.n564 VSUBS 0.005913f
C772 B.n565 VSUBS 0.005913f
C773 B.n566 VSUBS 0.005913f
C774 B.n567 VSUBS 0.005913f
C775 B.n568 VSUBS 0.005913f
C776 B.n569 VSUBS 0.005913f
C777 B.n570 VSUBS 0.005913f
C778 B.n571 VSUBS 0.005913f
C779 B.n572 VSUBS 0.005913f
C780 B.n573 VSUBS 0.005913f
C781 B.n574 VSUBS 0.005913f
C782 B.n575 VSUBS 0.005913f
C783 B.n576 VSUBS 0.005913f
C784 B.n577 VSUBS 0.005913f
C785 B.n578 VSUBS 0.005913f
C786 B.n579 VSUBS 0.005913f
C787 B.n580 VSUBS 0.005913f
C788 B.n581 VSUBS 0.005913f
C789 B.n582 VSUBS 0.005913f
C790 B.n583 VSUBS 0.005913f
C791 B.n584 VSUBS 0.005913f
C792 B.n585 VSUBS 0.005913f
C793 B.n586 VSUBS 0.005913f
C794 B.n587 VSUBS 0.005913f
C795 B.n588 VSUBS 0.005913f
C796 B.n589 VSUBS 0.005913f
C797 B.n590 VSUBS 0.005913f
C798 B.n591 VSUBS 0.005913f
C799 B.n592 VSUBS 0.005913f
C800 B.n593 VSUBS 0.005913f
C801 B.n594 VSUBS 0.005913f
C802 B.n595 VSUBS 0.005913f
C803 B.n596 VSUBS 0.005913f
C804 B.n597 VSUBS 0.005913f
C805 B.n598 VSUBS 0.014006f
C806 B.n599 VSUBS 0.014006f
C807 B.n600 VSUBS 0.013647f
C808 B.n601 VSUBS 0.005913f
C809 B.n602 VSUBS 0.005913f
C810 B.n603 VSUBS 0.005913f
C811 B.n604 VSUBS 0.005913f
C812 B.n605 VSUBS 0.005913f
C813 B.n606 VSUBS 0.005913f
C814 B.n607 VSUBS 0.005913f
C815 B.n608 VSUBS 0.005913f
C816 B.n609 VSUBS 0.005913f
C817 B.n610 VSUBS 0.005913f
C818 B.n611 VSUBS 0.005913f
C819 B.n612 VSUBS 0.005913f
C820 B.n613 VSUBS 0.005913f
C821 B.n614 VSUBS 0.005913f
C822 B.n615 VSUBS 0.005913f
C823 B.n616 VSUBS 0.005913f
C824 B.n617 VSUBS 0.005913f
C825 B.n618 VSUBS 0.005913f
C826 B.n619 VSUBS 0.005913f
C827 B.n620 VSUBS 0.005913f
C828 B.n621 VSUBS 0.005913f
C829 B.n622 VSUBS 0.005913f
C830 B.n623 VSUBS 0.005913f
C831 B.n624 VSUBS 0.005913f
C832 B.n625 VSUBS 0.005913f
C833 B.n626 VSUBS 0.005913f
C834 B.n627 VSUBS 0.005913f
C835 B.n628 VSUBS 0.005913f
C836 B.n629 VSUBS 0.005913f
C837 B.n630 VSUBS 0.005913f
C838 B.n631 VSUBS 0.005913f
C839 B.n632 VSUBS 0.005913f
C840 B.n633 VSUBS 0.005913f
C841 B.n634 VSUBS 0.005913f
C842 B.n635 VSUBS 0.01339f
C843 VDD1.n0 VSUBS 0.021647f
C844 VDD1.n1 VSUBS 0.020087f
C845 VDD1.n2 VSUBS 0.010794f
C846 VDD1.n3 VSUBS 0.025513f
C847 VDD1.n4 VSUBS 0.011429f
C848 VDD1.n5 VSUBS 0.020087f
C849 VDD1.n6 VSUBS 0.010794f
C850 VDD1.n7 VSUBS 0.025513f
C851 VDD1.n8 VSUBS 0.025513f
C852 VDD1.n9 VSUBS 0.011429f
C853 VDD1.n10 VSUBS 0.020087f
C854 VDD1.n11 VSUBS 0.010794f
C855 VDD1.n12 VSUBS 0.025513f
C856 VDD1.n13 VSUBS 0.011429f
C857 VDD1.n14 VSUBS 0.020087f
C858 VDD1.n15 VSUBS 0.010794f
C859 VDD1.n16 VSUBS 0.025513f
C860 VDD1.n17 VSUBS 0.011429f
C861 VDD1.n18 VSUBS 0.020087f
C862 VDD1.n19 VSUBS 0.010794f
C863 VDD1.n20 VSUBS 0.025513f
C864 VDD1.n21 VSUBS 0.011429f
C865 VDD1.n22 VSUBS 0.020087f
C866 VDD1.n23 VSUBS 0.010794f
C867 VDD1.n24 VSUBS 0.025513f
C868 VDD1.n25 VSUBS 0.011429f
C869 VDD1.n26 VSUBS 0.140411f
C870 VDD1.t0 VSUBS 0.054608f
C871 VDD1.n27 VSUBS 0.019135f
C872 VDD1.n28 VSUBS 0.01623f
C873 VDD1.n29 VSUBS 0.010794f
C874 VDD1.n30 VSUBS 1.26436f
C875 VDD1.n31 VSUBS 0.020087f
C876 VDD1.n32 VSUBS 0.010794f
C877 VDD1.n33 VSUBS 0.011429f
C878 VDD1.n34 VSUBS 0.025513f
C879 VDD1.n35 VSUBS 0.025513f
C880 VDD1.n36 VSUBS 0.011429f
C881 VDD1.n37 VSUBS 0.010794f
C882 VDD1.n38 VSUBS 0.020087f
C883 VDD1.n39 VSUBS 0.020087f
C884 VDD1.n40 VSUBS 0.010794f
C885 VDD1.n41 VSUBS 0.011429f
C886 VDD1.n42 VSUBS 0.025513f
C887 VDD1.n43 VSUBS 0.025513f
C888 VDD1.n44 VSUBS 0.011429f
C889 VDD1.n45 VSUBS 0.010794f
C890 VDD1.n46 VSUBS 0.020087f
C891 VDD1.n47 VSUBS 0.020087f
C892 VDD1.n48 VSUBS 0.010794f
C893 VDD1.n49 VSUBS 0.011429f
C894 VDD1.n50 VSUBS 0.025513f
C895 VDD1.n51 VSUBS 0.025513f
C896 VDD1.n52 VSUBS 0.011429f
C897 VDD1.n53 VSUBS 0.010794f
C898 VDD1.n54 VSUBS 0.020087f
C899 VDD1.n55 VSUBS 0.020087f
C900 VDD1.n56 VSUBS 0.010794f
C901 VDD1.n57 VSUBS 0.011429f
C902 VDD1.n58 VSUBS 0.025513f
C903 VDD1.n59 VSUBS 0.025513f
C904 VDD1.n60 VSUBS 0.011429f
C905 VDD1.n61 VSUBS 0.010794f
C906 VDD1.n62 VSUBS 0.020087f
C907 VDD1.n63 VSUBS 0.020087f
C908 VDD1.n64 VSUBS 0.010794f
C909 VDD1.n65 VSUBS 0.011429f
C910 VDD1.n66 VSUBS 0.025513f
C911 VDD1.n67 VSUBS 0.025513f
C912 VDD1.n68 VSUBS 0.011429f
C913 VDD1.n69 VSUBS 0.010794f
C914 VDD1.n70 VSUBS 0.020087f
C915 VDD1.n71 VSUBS 0.020087f
C916 VDD1.n72 VSUBS 0.010794f
C917 VDD1.n73 VSUBS 0.011111f
C918 VDD1.n74 VSUBS 0.011111f
C919 VDD1.n75 VSUBS 0.025513f
C920 VDD1.n76 VSUBS 0.060317f
C921 VDD1.n77 VSUBS 0.011429f
C922 VDD1.n78 VSUBS 0.010794f
C923 VDD1.n79 VSUBS 0.050821f
C924 VDD1.n80 VSUBS 0.045148f
C925 VDD1.n81 VSUBS 0.021647f
C926 VDD1.n82 VSUBS 0.020087f
C927 VDD1.n83 VSUBS 0.010794f
C928 VDD1.n84 VSUBS 0.025513f
C929 VDD1.n85 VSUBS 0.011429f
C930 VDD1.n86 VSUBS 0.020087f
C931 VDD1.n87 VSUBS 0.010794f
C932 VDD1.n88 VSUBS 0.025513f
C933 VDD1.n89 VSUBS 0.011429f
C934 VDD1.n90 VSUBS 0.020087f
C935 VDD1.n91 VSUBS 0.010794f
C936 VDD1.n92 VSUBS 0.025513f
C937 VDD1.n93 VSUBS 0.011429f
C938 VDD1.n94 VSUBS 0.020087f
C939 VDD1.n95 VSUBS 0.010794f
C940 VDD1.n96 VSUBS 0.025513f
C941 VDD1.n97 VSUBS 0.011429f
C942 VDD1.n98 VSUBS 0.020087f
C943 VDD1.n99 VSUBS 0.010794f
C944 VDD1.n100 VSUBS 0.025513f
C945 VDD1.n101 VSUBS 0.011429f
C946 VDD1.n102 VSUBS 0.020087f
C947 VDD1.n103 VSUBS 0.010794f
C948 VDD1.n104 VSUBS 0.025513f
C949 VDD1.n105 VSUBS 0.011429f
C950 VDD1.n106 VSUBS 0.140411f
C951 VDD1.t1 VSUBS 0.054608f
C952 VDD1.n107 VSUBS 0.019135f
C953 VDD1.n108 VSUBS 0.01623f
C954 VDD1.n109 VSUBS 0.010794f
C955 VDD1.n110 VSUBS 1.26436f
C956 VDD1.n111 VSUBS 0.020087f
C957 VDD1.n112 VSUBS 0.010794f
C958 VDD1.n113 VSUBS 0.011429f
C959 VDD1.n114 VSUBS 0.025513f
C960 VDD1.n115 VSUBS 0.025513f
C961 VDD1.n116 VSUBS 0.011429f
C962 VDD1.n117 VSUBS 0.010794f
C963 VDD1.n118 VSUBS 0.020087f
C964 VDD1.n119 VSUBS 0.020087f
C965 VDD1.n120 VSUBS 0.010794f
C966 VDD1.n121 VSUBS 0.011429f
C967 VDD1.n122 VSUBS 0.025513f
C968 VDD1.n123 VSUBS 0.025513f
C969 VDD1.n124 VSUBS 0.011429f
C970 VDD1.n125 VSUBS 0.010794f
C971 VDD1.n126 VSUBS 0.020087f
C972 VDD1.n127 VSUBS 0.020087f
C973 VDD1.n128 VSUBS 0.010794f
C974 VDD1.n129 VSUBS 0.011429f
C975 VDD1.n130 VSUBS 0.025513f
C976 VDD1.n131 VSUBS 0.025513f
C977 VDD1.n132 VSUBS 0.011429f
C978 VDD1.n133 VSUBS 0.010794f
C979 VDD1.n134 VSUBS 0.020087f
C980 VDD1.n135 VSUBS 0.020087f
C981 VDD1.n136 VSUBS 0.010794f
C982 VDD1.n137 VSUBS 0.011429f
C983 VDD1.n138 VSUBS 0.025513f
C984 VDD1.n139 VSUBS 0.025513f
C985 VDD1.n140 VSUBS 0.011429f
C986 VDD1.n141 VSUBS 0.010794f
C987 VDD1.n142 VSUBS 0.020087f
C988 VDD1.n143 VSUBS 0.020087f
C989 VDD1.n144 VSUBS 0.010794f
C990 VDD1.n145 VSUBS 0.011429f
C991 VDD1.n146 VSUBS 0.025513f
C992 VDD1.n147 VSUBS 0.025513f
C993 VDD1.n148 VSUBS 0.025513f
C994 VDD1.n149 VSUBS 0.011429f
C995 VDD1.n150 VSUBS 0.010794f
C996 VDD1.n151 VSUBS 0.020087f
C997 VDD1.n152 VSUBS 0.020087f
C998 VDD1.n153 VSUBS 0.010794f
C999 VDD1.n154 VSUBS 0.011111f
C1000 VDD1.n155 VSUBS 0.011111f
C1001 VDD1.n156 VSUBS 0.025513f
C1002 VDD1.n157 VSUBS 0.060317f
C1003 VDD1.n158 VSUBS 0.011429f
C1004 VDD1.n159 VSUBS 0.010794f
C1005 VDD1.n160 VSUBS 0.050821f
C1006 VDD1.n161 VSUBS 0.666954f
C1007 VTAIL.n0 VSUBS 0.030769f
C1008 VTAIL.n1 VSUBS 0.028552f
C1009 VTAIL.n2 VSUBS 0.015343f
C1010 VTAIL.n3 VSUBS 0.036265f
C1011 VTAIL.n4 VSUBS 0.016245f
C1012 VTAIL.n5 VSUBS 0.028552f
C1013 VTAIL.n6 VSUBS 0.015343f
C1014 VTAIL.n7 VSUBS 0.036265f
C1015 VTAIL.n8 VSUBS 0.016245f
C1016 VTAIL.n9 VSUBS 0.028552f
C1017 VTAIL.n10 VSUBS 0.015343f
C1018 VTAIL.n11 VSUBS 0.036265f
C1019 VTAIL.n12 VSUBS 0.016245f
C1020 VTAIL.n13 VSUBS 0.028552f
C1021 VTAIL.n14 VSUBS 0.015343f
C1022 VTAIL.n15 VSUBS 0.036265f
C1023 VTAIL.n16 VSUBS 0.016245f
C1024 VTAIL.n17 VSUBS 0.028552f
C1025 VTAIL.n18 VSUBS 0.015343f
C1026 VTAIL.n19 VSUBS 0.036265f
C1027 VTAIL.n20 VSUBS 0.016245f
C1028 VTAIL.n21 VSUBS 0.028552f
C1029 VTAIL.n22 VSUBS 0.015343f
C1030 VTAIL.n23 VSUBS 0.036265f
C1031 VTAIL.n24 VSUBS 0.016245f
C1032 VTAIL.n25 VSUBS 0.199585f
C1033 VTAIL.t2 VSUBS 0.077621f
C1034 VTAIL.n26 VSUBS 0.027198f
C1035 VTAIL.n27 VSUBS 0.02307f
C1036 VTAIL.n28 VSUBS 0.015343f
C1037 VTAIL.n29 VSUBS 1.7972f
C1038 VTAIL.n30 VSUBS 0.028552f
C1039 VTAIL.n31 VSUBS 0.015343f
C1040 VTAIL.n32 VSUBS 0.016245f
C1041 VTAIL.n33 VSUBS 0.036265f
C1042 VTAIL.n34 VSUBS 0.036265f
C1043 VTAIL.n35 VSUBS 0.016245f
C1044 VTAIL.n36 VSUBS 0.015343f
C1045 VTAIL.n37 VSUBS 0.028552f
C1046 VTAIL.n38 VSUBS 0.028552f
C1047 VTAIL.n39 VSUBS 0.015343f
C1048 VTAIL.n40 VSUBS 0.016245f
C1049 VTAIL.n41 VSUBS 0.036265f
C1050 VTAIL.n42 VSUBS 0.036265f
C1051 VTAIL.n43 VSUBS 0.016245f
C1052 VTAIL.n44 VSUBS 0.015343f
C1053 VTAIL.n45 VSUBS 0.028552f
C1054 VTAIL.n46 VSUBS 0.028552f
C1055 VTAIL.n47 VSUBS 0.015343f
C1056 VTAIL.n48 VSUBS 0.016245f
C1057 VTAIL.n49 VSUBS 0.036265f
C1058 VTAIL.n50 VSUBS 0.036265f
C1059 VTAIL.n51 VSUBS 0.016245f
C1060 VTAIL.n52 VSUBS 0.015343f
C1061 VTAIL.n53 VSUBS 0.028552f
C1062 VTAIL.n54 VSUBS 0.028552f
C1063 VTAIL.n55 VSUBS 0.015343f
C1064 VTAIL.n56 VSUBS 0.016245f
C1065 VTAIL.n57 VSUBS 0.036265f
C1066 VTAIL.n58 VSUBS 0.036265f
C1067 VTAIL.n59 VSUBS 0.016245f
C1068 VTAIL.n60 VSUBS 0.015343f
C1069 VTAIL.n61 VSUBS 0.028552f
C1070 VTAIL.n62 VSUBS 0.028552f
C1071 VTAIL.n63 VSUBS 0.015343f
C1072 VTAIL.n64 VSUBS 0.016245f
C1073 VTAIL.n65 VSUBS 0.036265f
C1074 VTAIL.n66 VSUBS 0.036265f
C1075 VTAIL.n67 VSUBS 0.036265f
C1076 VTAIL.n68 VSUBS 0.016245f
C1077 VTAIL.n69 VSUBS 0.015343f
C1078 VTAIL.n70 VSUBS 0.028552f
C1079 VTAIL.n71 VSUBS 0.028552f
C1080 VTAIL.n72 VSUBS 0.015343f
C1081 VTAIL.n73 VSUBS 0.015794f
C1082 VTAIL.n74 VSUBS 0.015794f
C1083 VTAIL.n75 VSUBS 0.036265f
C1084 VTAIL.n76 VSUBS 0.085737f
C1085 VTAIL.n77 VSUBS 0.016245f
C1086 VTAIL.n78 VSUBS 0.015343f
C1087 VTAIL.n79 VSUBS 0.072238f
C1088 VTAIL.n80 VSUBS 0.043209f
C1089 VTAIL.n81 VSUBS 2.08607f
C1090 VTAIL.n82 VSUBS 0.030769f
C1091 VTAIL.n83 VSUBS 0.028552f
C1092 VTAIL.n84 VSUBS 0.015343f
C1093 VTAIL.n85 VSUBS 0.036265f
C1094 VTAIL.n86 VSUBS 0.016245f
C1095 VTAIL.n87 VSUBS 0.028552f
C1096 VTAIL.n88 VSUBS 0.015343f
C1097 VTAIL.n89 VSUBS 0.036265f
C1098 VTAIL.n90 VSUBS 0.036265f
C1099 VTAIL.n91 VSUBS 0.016245f
C1100 VTAIL.n92 VSUBS 0.028552f
C1101 VTAIL.n93 VSUBS 0.015343f
C1102 VTAIL.n94 VSUBS 0.036265f
C1103 VTAIL.n95 VSUBS 0.016245f
C1104 VTAIL.n96 VSUBS 0.028552f
C1105 VTAIL.n97 VSUBS 0.015343f
C1106 VTAIL.n98 VSUBS 0.036265f
C1107 VTAIL.n99 VSUBS 0.016245f
C1108 VTAIL.n100 VSUBS 0.028552f
C1109 VTAIL.n101 VSUBS 0.015343f
C1110 VTAIL.n102 VSUBS 0.036265f
C1111 VTAIL.n103 VSUBS 0.016245f
C1112 VTAIL.n104 VSUBS 0.028552f
C1113 VTAIL.n105 VSUBS 0.015343f
C1114 VTAIL.n106 VSUBS 0.036265f
C1115 VTAIL.n107 VSUBS 0.016245f
C1116 VTAIL.n108 VSUBS 0.199585f
C1117 VTAIL.t1 VSUBS 0.077621f
C1118 VTAIL.n109 VSUBS 0.027198f
C1119 VTAIL.n110 VSUBS 0.02307f
C1120 VTAIL.n111 VSUBS 0.015343f
C1121 VTAIL.n112 VSUBS 1.7972f
C1122 VTAIL.n113 VSUBS 0.028552f
C1123 VTAIL.n114 VSUBS 0.015343f
C1124 VTAIL.n115 VSUBS 0.016245f
C1125 VTAIL.n116 VSUBS 0.036265f
C1126 VTAIL.n117 VSUBS 0.036265f
C1127 VTAIL.n118 VSUBS 0.016245f
C1128 VTAIL.n119 VSUBS 0.015343f
C1129 VTAIL.n120 VSUBS 0.028552f
C1130 VTAIL.n121 VSUBS 0.028552f
C1131 VTAIL.n122 VSUBS 0.015343f
C1132 VTAIL.n123 VSUBS 0.016245f
C1133 VTAIL.n124 VSUBS 0.036265f
C1134 VTAIL.n125 VSUBS 0.036265f
C1135 VTAIL.n126 VSUBS 0.016245f
C1136 VTAIL.n127 VSUBS 0.015343f
C1137 VTAIL.n128 VSUBS 0.028552f
C1138 VTAIL.n129 VSUBS 0.028552f
C1139 VTAIL.n130 VSUBS 0.015343f
C1140 VTAIL.n131 VSUBS 0.016245f
C1141 VTAIL.n132 VSUBS 0.036265f
C1142 VTAIL.n133 VSUBS 0.036265f
C1143 VTAIL.n134 VSUBS 0.016245f
C1144 VTAIL.n135 VSUBS 0.015343f
C1145 VTAIL.n136 VSUBS 0.028552f
C1146 VTAIL.n137 VSUBS 0.028552f
C1147 VTAIL.n138 VSUBS 0.015343f
C1148 VTAIL.n139 VSUBS 0.016245f
C1149 VTAIL.n140 VSUBS 0.036265f
C1150 VTAIL.n141 VSUBS 0.036265f
C1151 VTAIL.n142 VSUBS 0.016245f
C1152 VTAIL.n143 VSUBS 0.015343f
C1153 VTAIL.n144 VSUBS 0.028552f
C1154 VTAIL.n145 VSUBS 0.028552f
C1155 VTAIL.n146 VSUBS 0.015343f
C1156 VTAIL.n147 VSUBS 0.016245f
C1157 VTAIL.n148 VSUBS 0.036265f
C1158 VTAIL.n149 VSUBS 0.036265f
C1159 VTAIL.n150 VSUBS 0.016245f
C1160 VTAIL.n151 VSUBS 0.015343f
C1161 VTAIL.n152 VSUBS 0.028552f
C1162 VTAIL.n153 VSUBS 0.028552f
C1163 VTAIL.n154 VSUBS 0.015343f
C1164 VTAIL.n155 VSUBS 0.015794f
C1165 VTAIL.n156 VSUBS 0.015794f
C1166 VTAIL.n157 VSUBS 0.036265f
C1167 VTAIL.n158 VSUBS 0.085737f
C1168 VTAIL.n159 VSUBS 0.016245f
C1169 VTAIL.n160 VSUBS 0.015343f
C1170 VTAIL.n161 VSUBS 0.072238f
C1171 VTAIL.n162 VSUBS 0.043209f
C1172 VTAIL.n163 VSUBS 2.13049f
C1173 VTAIL.n164 VSUBS 0.030769f
C1174 VTAIL.n165 VSUBS 0.028552f
C1175 VTAIL.n166 VSUBS 0.015343f
C1176 VTAIL.n167 VSUBS 0.036265f
C1177 VTAIL.n168 VSUBS 0.016245f
C1178 VTAIL.n169 VSUBS 0.028552f
C1179 VTAIL.n170 VSUBS 0.015343f
C1180 VTAIL.n171 VSUBS 0.036265f
C1181 VTAIL.n172 VSUBS 0.036265f
C1182 VTAIL.n173 VSUBS 0.016245f
C1183 VTAIL.n174 VSUBS 0.028552f
C1184 VTAIL.n175 VSUBS 0.015343f
C1185 VTAIL.n176 VSUBS 0.036265f
C1186 VTAIL.n177 VSUBS 0.016245f
C1187 VTAIL.n178 VSUBS 0.028552f
C1188 VTAIL.n179 VSUBS 0.015343f
C1189 VTAIL.n180 VSUBS 0.036265f
C1190 VTAIL.n181 VSUBS 0.016245f
C1191 VTAIL.n182 VSUBS 0.028552f
C1192 VTAIL.n183 VSUBS 0.015343f
C1193 VTAIL.n184 VSUBS 0.036265f
C1194 VTAIL.n185 VSUBS 0.016245f
C1195 VTAIL.n186 VSUBS 0.028552f
C1196 VTAIL.n187 VSUBS 0.015343f
C1197 VTAIL.n188 VSUBS 0.036265f
C1198 VTAIL.n189 VSUBS 0.016245f
C1199 VTAIL.n190 VSUBS 0.199585f
C1200 VTAIL.t3 VSUBS 0.077621f
C1201 VTAIL.n191 VSUBS 0.027198f
C1202 VTAIL.n192 VSUBS 0.02307f
C1203 VTAIL.n193 VSUBS 0.015343f
C1204 VTAIL.n194 VSUBS 1.7972f
C1205 VTAIL.n195 VSUBS 0.028552f
C1206 VTAIL.n196 VSUBS 0.015343f
C1207 VTAIL.n197 VSUBS 0.016245f
C1208 VTAIL.n198 VSUBS 0.036265f
C1209 VTAIL.n199 VSUBS 0.036265f
C1210 VTAIL.n200 VSUBS 0.016245f
C1211 VTAIL.n201 VSUBS 0.015343f
C1212 VTAIL.n202 VSUBS 0.028552f
C1213 VTAIL.n203 VSUBS 0.028552f
C1214 VTAIL.n204 VSUBS 0.015343f
C1215 VTAIL.n205 VSUBS 0.016245f
C1216 VTAIL.n206 VSUBS 0.036265f
C1217 VTAIL.n207 VSUBS 0.036265f
C1218 VTAIL.n208 VSUBS 0.016245f
C1219 VTAIL.n209 VSUBS 0.015343f
C1220 VTAIL.n210 VSUBS 0.028552f
C1221 VTAIL.n211 VSUBS 0.028552f
C1222 VTAIL.n212 VSUBS 0.015343f
C1223 VTAIL.n213 VSUBS 0.016245f
C1224 VTAIL.n214 VSUBS 0.036265f
C1225 VTAIL.n215 VSUBS 0.036265f
C1226 VTAIL.n216 VSUBS 0.016245f
C1227 VTAIL.n217 VSUBS 0.015343f
C1228 VTAIL.n218 VSUBS 0.028552f
C1229 VTAIL.n219 VSUBS 0.028552f
C1230 VTAIL.n220 VSUBS 0.015343f
C1231 VTAIL.n221 VSUBS 0.016245f
C1232 VTAIL.n222 VSUBS 0.036265f
C1233 VTAIL.n223 VSUBS 0.036265f
C1234 VTAIL.n224 VSUBS 0.016245f
C1235 VTAIL.n225 VSUBS 0.015343f
C1236 VTAIL.n226 VSUBS 0.028552f
C1237 VTAIL.n227 VSUBS 0.028552f
C1238 VTAIL.n228 VSUBS 0.015343f
C1239 VTAIL.n229 VSUBS 0.016245f
C1240 VTAIL.n230 VSUBS 0.036265f
C1241 VTAIL.n231 VSUBS 0.036265f
C1242 VTAIL.n232 VSUBS 0.016245f
C1243 VTAIL.n233 VSUBS 0.015343f
C1244 VTAIL.n234 VSUBS 0.028552f
C1245 VTAIL.n235 VSUBS 0.028552f
C1246 VTAIL.n236 VSUBS 0.015343f
C1247 VTAIL.n237 VSUBS 0.015794f
C1248 VTAIL.n238 VSUBS 0.015794f
C1249 VTAIL.n239 VSUBS 0.036265f
C1250 VTAIL.n240 VSUBS 0.085737f
C1251 VTAIL.n241 VSUBS 0.016245f
C1252 VTAIL.n242 VSUBS 0.015343f
C1253 VTAIL.n243 VSUBS 0.072238f
C1254 VTAIL.n244 VSUBS 0.043209f
C1255 VTAIL.n245 VSUBS 1.93142f
C1256 VTAIL.n246 VSUBS 0.030769f
C1257 VTAIL.n247 VSUBS 0.028552f
C1258 VTAIL.n248 VSUBS 0.015343f
C1259 VTAIL.n249 VSUBS 0.036265f
C1260 VTAIL.n250 VSUBS 0.016245f
C1261 VTAIL.n251 VSUBS 0.028552f
C1262 VTAIL.n252 VSUBS 0.015343f
C1263 VTAIL.n253 VSUBS 0.036265f
C1264 VTAIL.n254 VSUBS 0.016245f
C1265 VTAIL.n255 VSUBS 0.028552f
C1266 VTAIL.n256 VSUBS 0.015343f
C1267 VTAIL.n257 VSUBS 0.036265f
C1268 VTAIL.n258 VSUBS 0.016245f
C1269 VTAIL.n259 VSUBS 0.028552f
C1270 VTAIL.n260 VSUBS 0.015343f
C1271 VTAIL.n261 VSUBS 0.036265f
C1272 VTAIL.n262 VSUBS 0.016245f
C1273 VTAIL.n263 VSUBS 0.028552f
C1274 VTAIL.n264 VSUBS 0.015343f
C1275 VTAIL.n265 VSUBS 0.036265f
C1276 VTAIL.n266 VSUBS 0.016245f
C1277 VTAIL.n267 VSUBS 0.028552f
C1278 VTAIL.n268 VSUBS 0.015343f
C1279 VTAIL.n269 VSUBS 0.036265f
C1280 VTAIL.n270 VSUBS 0.016245f
C1281 VTAIL.n271 VSUBS 0.199585f
C1282 VTAIL.t0 VSUBS 0.077621f
C1283 VTAIL.n272 VSUBS 0.027198f
C1284 VTAIL.n273 VSUBS 0.02307f
C1285 VTAIL.n274 VSUBS 0.015343f
C1286 VTAIL.n275 VSUBS 1.7972f
C1287 VTAIL.n276 VSUBS 0.028552f
C1288 VTAIL.n277 VSUBS 0.015343f
C1289 VTAIL.n278 VSUBS 0.016245f
C1290 VTAIL.n279 VSUBS 0.036265f
C1291 VTAIL.n280 VSUBS 0.036265f
C1292 VTAIL.n281 VSUBS 0.016245f
C1293 VTAIL.n282 VSUBS 0.015343f
C1294 VTAIL.n283 VSUBS 0.028552f
C1295 VTAIL.n284 VSUBS 0.028552f
C1296 VTAIL.n285 VSUBS 0.015343f
C1297 VTAIL.n286 VSUBS 0.016245f
C1298 VTAIL.n287 VSUBS 0.036265f
C1299 VTAIL.n288 VSUBS 0.036265f
C1300 VTAIL.n289 VSUBS 0.016245f
C1301 VTAIL.n290 VSUBS 0.015343f
C1302 VTAIL.n291 VSUBS 0.028552f
C1303 VTAIL.n292 VSUBS 0.028552f
C1304 VTAIL.n293 VSUBS 0.015343f
C1305 VTAIL.n294 VSUBS 0.016245f
C1306 VTAIL.n295 VSUBS 0.036265f
C1307 VTAIL.n296 VSUBS 0.036265f
C1308 VTAIL.n297 VSUBS 0.016245f
C1309 VTAIL.n298 VSUBS 0.015343f
C1310 VTAIL.n299 VSUBS 0.028552f
C1311 VTAIL.n300 VSUBS 0.028552f
C1312 VTAIL.n301 VSUBS 0.015343f
C1313 VTAIL.n302 VSUBS 0.016245f
C1314 VTAIL.n303 VSUBS 0.036265f
C1315 VTAIL.n304 VSUBS 0.036265f
C1316 VTAIL.n305 VSUBS 0.016245f
C1317 VTAIL.n306 VSUBS 0.015343f
C1318 VTAIL.n307 VSUBS 0.028552f
C1319 VTAIL.n308 VSUBS 0.028552f
C1320 VTAIL.n309 VSUBS 0.015343f
C1321 VTAIL.n310 VSUBS 0.016245f
C1322 VTAIL.n311 VSUBS 0.036265f
C1323 VTAIL.n312 VSUBS 0.036265f
C1324 VTAIL.n313 VSUBS 0.036265f
C1325 VTAIL.n314 VSUBS 0.016245f
C1326 VTAIL.n315 VSUBS 0.015343f
C1327 VTAIL.n316 VSUBS 0.028552f
C1328 VTAIL.n317 VSUBS 0.028552f
C1329 VTAIL.n318 VSUBS 0.015343f
C1330 VTAIL.n319 VSUBS 0.015794f
C1331 VTAIL.n320 VSUBS 0.015794f
C1332 VTAIL.n321 VSUBS 0.036265f
C1333 VTAIL.n322 VSUBS 0.085737f
C1334 VTAIL.n323 VSUBS 0.016245f
C1335 VTAIL.n324 VSUBS 0.015343f
C1336 VTAIL.n325 VSUBS 0.072238f
C1337 VTAIL.n326 VSUBS 0.043209f
C1338 VTAIL.n327 VSUBS 1.83307f
C1339 VP.t1 VSUBS 4.71291f
C1340 VP.t0 VSUBS 4.11851f
C1341 VP.n0 VSUBS 6.08329f
.ends

