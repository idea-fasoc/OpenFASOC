.subcircuit ind_top
XL1 outp outn VDD sky130_fd_pr__ind_05_220
.ends 
