* NGSPICE file created from diff_pair_sample_1428.ext - technology: sky130A

.subckt diff_pair_sample_1428 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=2.1801 pd=11.96 as=0 ps=0 w=5.59 l=2.94
X1 VTAIL.t7 VN.t0 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1801 pd=11.96 as=0.92235 ps=5.92 w=5.59 l=2.94
X2 VDD1.t3 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.92235 pd=5.92 as=2.1801 ps=11.96 w=5.59 l=2.94
X3 VTAIL.t6 VN.t1 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1801 pd=11.96 as=0.92235 ps=5.92 w=5.59 l=2.94
X4 VDD1.t2 VP.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.92235 pd=5.92 as=2.1801 ps=11.96 w=5.59 l=2.94
X5 VTAIL.t0 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1801 pd=11.96 as=0.92235 ps=5.92 w=5.59 l=2.94
X6 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=2.1801 pd=11.96 as=0 ps=0 w=5.59 l=2.94
X7 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.1801 pd=11.96 as=0 ps=0 w=5.59 l=2.94
X8 VDD2.t1 VN.t2 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=0.92235 pd=5.92 as=2.1801 ps=11.96 w=5.59 l=2.94
X9 VTAIL.t2 VP.t3 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1801 pd=11.96 as=0.92235 ps=5.92 w=5.59 l=2.94
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.1801 pd=11.96 as=0 ps=0 w=5.59 l=2.94
X11 VDD2.t0 VN.t3 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.92235 pd=5.92 as=2.1801 ps=11.96 w=5.59 l=2.94
R0 B.n585 B.n584 585
R1 B.n586 B.n585 585
R2 B.n210 B.n97 585
R3 B.n209 B.n208 585
R4 B.n207 B.n206 585
R5 B.n205 B.n204 585
R6 B.n203 B.n202 585
R7 B.n201 B.n200 585
R8 B.n199 B.n198 585
R9 B.n197 B.n196 585
R10 B.n195 B.n194 585
R11 B.n193 B.n192 585
R12 B.n191 B.n190 585
R13 B.n189 B.n188 585
R14 B.n187 B.n186 585
R15 B.n185 B.n184 585
R16 B.n183 B.n182 585
R17 B.n181 B.n180 585
R18 B.n179 B.n178 585
R19 B.n177 B.n176 585
R20 B.n175 B.n174 585
R21 B.n173 B.n172 585
R22 B.n171 B.n170 585
R23 B.n169 B.n168 585
R24 B.n167 B.n166 585
R25 B.n165 B.n164 585
R26 B.n163 B.n162 585
R27 B.n161 B.n160 585
R28 B.n159 B.n158 585
R29 B.n157 B.n156 585
R30 B.n155 B.n154 585
R31 B.n153 B.n152 585
R32 B.n151 B.n150 585
R33 B.n148 B.n147 585
R34 B.n146 B.n145 585
R35 B.n144 B.n143 585
R36 B.n142 B.n141 585
R37 B.n140 B.n139 585
R38 B.n138 B.n137 585
R39 B.n136 B.n135 585
R40 B.n134 B.n133 585
R41 B.n132 B.n131 585
R42 B.n130 B.n129 585
R43 B.n128 B.n127 585
R44 B.n126 B.n125 585
R45 B.n124 B.n123 585
R46 B.n122 B.n121 585
R47 B.n120 B.n119 585
R48 B.n118 B.n117 585
R49 B.n116 B.n115 585
R50 B.n114 B.n113 585
R51 B.n112 B.n111 585
R52 B.n110 B.n109 585
R53 B.n108 B.n107 585
R54 B.n106 B.n105 585
R55 B.n104 B.n103 585
R56 B.n583 B.n69 585
R57 B.n587 B.n69 585
R58 B.n582 B.n68 585
R59 B.n588 B.n68 585
R60 B.n581 B.n580 585
R61 B.n580 B.n64 585
R62 B.n579 B.n63 585
R63 B.n594 B.n63 585
R64 B.n578 B.n62 585
R65 B.n595 B.n62 585
R66 B.n577 B.n61 585
R67 B.n596 B.n61 585
R68 B.n576 B.n575 585
R69 B.n575 B.n57 585
R70 B.n574 B.n56 585
R71 B.n602 B.n56 585
R72 B.n573 B.n55 585
R73 B.n603 B.n55 585
R74 B.n572 B.n54 585
R75 B.n604 B.n54 585
R76 B.n571 B.n570 585
R77 B.n570 B.n50 585
R78 B.n569 B.n49 585
R79 B.n610 B.n49 585
R80 B.n568 B.n48 585
R81 B.n611 B.n48 585
R82 B.n567 B.n47 585
R83 B.n612 B.n47 585
R84 B.n566 B.n565 585
R85 B.n565 B.n43 585
R86 B.n564 B.n42 585
R87 B.n618 B.n42 585
R88 B.n563 B.n41 585
R89 B.n619 B.n41 585
R90 B.n562 B.n40 585
R91 B.n620 B.n40 585
R92 B.n561 B.n560 585
R93 B.n560 B.n36 585
R94 B.n559 B.n35 585
R95 B.n626 B.n35 585
R96 B.n558 B.n34 585
R97 B.n627 B.n34 585
R98 B.n557 B.n33 585
R99 B.n628 B.n33 585
R100 B.n556 B.n555 585
R101 B.n555 B.n29 585
R102 B.n554 B.n28 585
R103 B.n634 B.n28 585
R104 B.n553 B.n27 585
R105 B.n635 B.n27 585
R106 B.n552 B.n26 585
R107 B.n636 B.n26 585
R108 B.n551 B.n550 585
R109 B.n550 B.n22 585
R110 B.n549 B.n21 585
R111 B.n642 B.n21 585
R112 B.n548 B.n20 585
R113 B.n643 B.n20 585
R114 B.n547 B.n19 585
R115 B.n644 B.n19 585
R116 B.n546 B.n545 585
R117 B.n545 B.n18 585
R118 B.n544 B.n14 585
R119 B.n650 B.n14 585
R120 B.n543 B.n13 585
R121 B.n651 B.n13 585
R122 B.n542 B.n12 585
R123 B.n652 B.n12 585
R124 B.n541 B.n540 585
R125 B.n540 B.n8 585
R126 B.n539 B.n7 585
R127 B.n658 B.n7 585
R128 B.n538 B.n6 585
R129 B.n659 B.n6 585
R130 B.n537 B.n5 585
R131 B.n660 B.n5 585
R132 B.n536 B.n535 585
R133 B.n535 B.n4 585
R134 B.n534 B.n211 585
R135 B.n534 B.n533 585
R136 B.n524 B.n212 585
R137 B.n213 B.n212 585
R138 B.n526 B.n525 585
R139 B.n527 B.n526 585
R140 B.n523 B.n218 585
R141 B.n218 B.n217 585
R142 B.n522 B.n521 585
R143 B.n521 B.n520 585
R144 B.n220 B.n219 585
R145 B.n513 B.n220 585
R146 B.n512 B.n511 585
R147 B.n514 B.n512 585
R148 B.n510 B.n225 585
R149 B.n225 B.n224 585
R150 B.n509 B.n508 585
R151 B.n508 B.n507 585
R152 B.n227 B.n226 585
R153 B.n228 B.n227 585
R154 B.n500 B.n499 585
R155 B.n501 B.n500 585
R156 B.n498 B.n233 585
R157 B.n233 B.n232 585
R158 B.n497 B.n496 585
R159 B.n496 B.n495 585
R160 B.n235 B.n234 585
R161 B.n236 B.n235 585
R162 B.n488 B.n487 585
R163 B.n489 B.n488 585
R164 B.n486 B.n240 585
R165 B.n244 B.n240 585
R166 B.n485 B.n484 585
R167 B.n484 B.n483 585
R168 B.n242 B.n241 585
R169 B.n243 B.n242 585
R170 B.n476 B.n475 585
R171 B.n477 B.n476 585
R172 B.n474 B.n249 585
R173 B.n249 B.n248 585
R174 B.n473 B.n472 585
R175 B.n472 B.n471 585
R176 B.n251 B.n250 585
R177 B.n252 B.n251 585
R178 B.n464 B.n463 585
R179 B.n465 B.n464 585
R180 B.n462 B.n257 585
R181 B.n257 B.n256 585
R182 B.n461 B.n460 585
R183 B.n460 B.n459 585
R184 B.n259 B.n258 585
R185 B.n260 B.n259 585
R186 B.n452 B.n451 585
R187 B.n453 B.n452 585
R188 B.n450 B.n264 585
R189 B.n268 B.n264 585
R190 B.n449 B.n448 585
R191 B.n448 B.n447 585
R192 B.n266 B.n265 585
R193 B.n267 B.n266 585
R194 B.n440 B.n439 585
R195 B.n441 B.n440 585
R196 B.n438 B.n273 585
R197 B.n273 B.n272 585
R198 B.n437 B.n436 585
R199 B.n436 B.n435 585
R200 B.n275 B.n274 585
R201 B.n276 B.n275 585
R202 B.n428 B.n427 585
R203 B.n429 B.n428 585
R204 B.n426 B.n281 585
R205 B.n281 B.n280 585
R206 B.n420 B.n419 585
R207 B.n418 B.n310 585
R208 B.n417 B.n309 585
R209 B.n422 B.n309 585
R210 B.n416 B.n415 585
R211 B.n414 B.n413 585
R212 B.n412 B.n411 585
R213 B.n410 B.n409 585
R214 B.n408 B.n407 585
R215 B.n406 B.n405 585
R216 B.n404 B.n403 585
R217 B.n402 B.n401 585
R218 B.n400 B.n399 585
R219 B.n398 B.n397 585
R220 B.n396 B.n395 585
R221 B.n394 B.n393 585
R222 B.n392 B.n391 585
R223 B.n390 B.n389 585
R224 B.n388 B.n387 585
R225 B.n386 B.n385 585
R226 B.n384 B.n383 585
R227 B.n382 B.n381 585
R228 B.n380 B.n379 585
R229 B.n378 B.n377 585
R230 B.n376 B.n375 585
R231 B.n374 B.n373 585
R232 B.n372 B.n371 585
R233 B.n370 B.n369 585
R234 B.n368 B.n367 585
R235 B.n366 B.n365 585
R236 B.n364 B.n363 585
R237 B.n362 B.n361 585
R238 B.n360 B.n359 585
R239 B.n357 B.n356 585
R240 B.n355 B.n354 585
R241 B.n353 B.n352 585
R242 B.n351 B.n350 585
R243 B.n349 B.n348 585
R244 B.n347 B.n346 585
R245 B.n345 B.n344 585
R246 B.n343 B.n342 585
R247 B.n341 B.n340 585
R248 B.n339 B.n338 585
R249 B.n337 B.n336 585
R250 B.n335 B.n334 585
R251 B.n333 B.n332 585
R252 B.n331 B.n330 585
R253 B.n329 B.n328 585
R254 B.n327 B.n326 585
R255 B.n325 B.n324 585
R256 B.n323 B.n322 585
R257 B.n321 B.n320 585
R258 B.n319 B.n318 585
R259 B.n317 B.n316 585
R260 B.n283 B.n282 585
R261 B.n425 B.n424 585
R262 B.n279 B.n278 585
R263 B.n280 B.n279 585
R264 B.n431 B.n430 585
R265 B.n430 B.n429 585
R266 B.n432 B.n277 585
R267 B.n277 B.n276 585
R268 B.n434 B.n433 585
R269 B.n435 B.n434 585
R270 B.n271 B.n270 585
R271 B.n272 B.n271 585
R272 B.n443 B.n442 585
R273 B.n442 B.n441 585
R274 B.n444 B.n269 585
R275 B.n269 B.n267 585
R276 B.n446 B.n445 585
R277 B.n447 B.n446 585
R278 B.n263 B.n262 585
R279 B.n268 B.n263 585
R280 B.n455 B.n454 585
R281 B.n454 B.n453 585
R282 B.n456 B.n261 585
R283 B.n261 B.n260 585
R284 B.n458 B.n457 585
R285 B.n459 B.n458 585
R286 B.n255 B.n254 585
R287 B.n256 B.n255 585
R288 B.n467 B.n466 585
R289 B.n466 B.n465 585
R290 B.n468 B.n253 585
R291 B.n253 B.n252 585
R292 B.n470 B.n469 585
R293 B.n471 B.n470 585
R294 B.n247 B.n246 585
R295 B.n248 B.n247 585
R296 B.n479 B.n478 585
R297 B.n478 B.n477 585
R298 B.n480 B.n245 585
R299 B.n245 B.n243 585
R300 B.n482 B.n481 585
R301 B.n483 B.n482 585
R302 B.n239 B.n238 585
R303 B.n244 B.n239 585
R304 B.n491 B.n490 585
R305 B.n490 B.n489 585
R306 B.n492 B.n237 585
R307 B.n237 B.n236 585
R308 B.n494 B.n493 585
R309 B.n495 B.n494 585
R310 B.n231 B.n230 585
R311 B.n232 B.n231 585
R312 B.n503 B.n502 585
R313 B.n502 B.n501 585
R314 B.n504 B.n229 585
R315 B.n229 B.n228 585
R316 B.n506 B.n505 585
R317 B.n507 B.n506 585
R318 B.n223 B.n222 585
R319 B.n224 B.n223 585
R320 B.n516 B.n515 585
R321 B.n515 B.n514 585
R322 B.n517 B.n221 585
R323 B.n513 B.n221 585
R324 B.n519 B.n518 585
R325 B.n520 B.n519 585
R326 B.n216 B.n215 585
R327 B.n217 B.n216 585
R328 B.n529 B.n528 585
R329 B.n528 B.n527 585
R330 B.n530 B.n214 585
R331 B.n214 B.n213 585
R332 B.n532 B.n531 585
R333 B.n533 B.n532 585
R334 B.n2 B.n0 585
R335 B.n4 B.n2 585
R336 B.n3 B.n1 585
R337 B.n659 B.n3 585
R338 B.n657 B.n656 585
R339 B.n658 B.n657 585
R340 B.n655 B.n9 585
R341 B.n9 B.n8 585
R342 B.n654 B.n653 585
R343 B.n653 B.n652 585
R344 B.n11 B.n10 585
R345 B.n651 B.n11 585
R346 B.n649 B.n648 585
R347 B.n650 B.n649 585
R348 B.n647 B.n15 585
R349 B.n18 B.n15 585
R350 B.n646 B.n645 585
R351 B.n645 B.n644 585
R352 B.n17 B.n16 585
R353 B.n643 B.n17 585
R354 B.n641 B.n640 585
R355 B.n642 B.n641 585
R356 B.n639 B.n23 585
R357 B.n23 B.n22 585
R358 B.n638 B.n637 585
R359 B.n637 B.n636 585
R360 B.n25 B.n24 585
R361 B.n635 B.n25 585
R362 B.n633 B.n632 585
R363 B.n634 B.n633 585
R364 B.n631 B.n30 585
R365 B.n30 B.n29 585
R366 B.n630 B.n629 585
R367 B.n629 B.n628 585
R368 B.n32 B.n31 585
R369 B.n627 B.n32 585
R370 B.n625 B.n624 585
R371 B.n626 B.n625 585
R372 B.n623 B.n37 585
R373 B.n37 B.n36 585
R374 B.n622 B.n621 585
R375 B.n621 B.n620 585
R376 B.n39 B.n38 585
R377 B.n619 B.n39 585
R378 B.n617 B.n616 585
R379 B.n618 B.n617 585
R380 B.n615 B.n44 585
R381 B.n44 B.n43 585
R382 B.n614 B.n613 585
R383 B.n613 B.n612 585
R384 B.n46 B.n45 585
R385 B.n611 B.n46 585
R386 B.n609 B.n608 585
R387 B.n610 B.n609 585
R388 B.n607 B.n51 585
R389 B.n51 B.n50 585
R390 B.n606 B.n605 585
R391 B.n605 B.n604 585
R392 B.n53 B.n52 585
R393 B.n603 B.n53 585
R394 B.n601 B.n600 585
R395 B.n602 B.n601 585
R396 B.n599 B.n58 585
R397 B.n58 B.n57 585
R398 B.n598 B.n597 585
R399 B.n597 B.n596 585
R400 B.n60 B.n59 585
R401 B.n595 B.n60 585
R402 B.n593 B.n592 585
R403 B.n594 B.n593 585
R404 B.n591 B.n65 585
R405 B.n65 B.n64 585
R406 B.n590 B.n589 585
R407 B.n589 B.n588 585
R408 B.n67 B.n66 585
R409 B.n587 B.n67 585
R410 B.n662 B.n661 585
R411 B.n661 B.n660 585
R412 B.n420 B.n279 502.111
R413 B.n103 B.n67 502.111
R414 B.n424 B.n281 502.111
R415 B.n585 B.n69 502.111
R416 B.n586 B.n96 256.663
R417 B.n586 B.n95 256.663
R418 B.n586 B.n94 256.663
R419 B.n586 B.n93 256.663
R420 B.n586 B.n92 256.663
R421 B.n586 B.n91 256.663
R422 B.n586 B.n90 256.663
R423 B.n586 B.n89 256.663
R424 B.n586 B.n88 256.663
R425 B.n586 B.n87 256.663
R426 B.n586 B.n86 256.663
R427 B.n586 B.n85 256.663
R428 B.n586 B.n84 256.663
R429 B.n586 B.n83 256.663
R430 B.n586 B.n82 256.663
R431 B.n586 B.n81 256.663
R432 B.n586 B.n80 256.663
R433 B.n586 B.n79 256.663
R434 B.n586 B.n78 256.663
R435 B.n586 B.n77 256.663
R436 B.n586 B.n76 256.663
R437 B.n586 B.n75 256.663
R438 B.n586 B.n74 256.663
R439 B.n586 B.n73 256.663
R440 B.n586 B.n72 256.663
R441 B.n586 B.n71 256.663
R442 B.n586 B.n70 256.663
R443 B.n422 B.n421 256.663
R444 B.n422 B.n284 256.663
R445 B.n422 B.n285 256.663
R446 B.n422 B.n286 256.663
R447 B.n422 B.n287 256.663
R448 B.n422 B.n288 256.663
R449 B.n422 B.n289 256.663
R450 B.n422 B.n290 256.663
R451 B.n422 B.n291 256.663
R452 B.n422 B.n292 256.663
R453 B.n422 B.n293 256.663
R454 B.n422 B.n294 256.663
R455 B.n422 B.n295 256.663
R456 B.n422 B.n296 256.663
R457 B.n422 B.n297 256.663
R458 B.n422 B.n298 256.663
R459 B.n422 B.n299 256.663
R460 B.n422 B.n300 256.663
R461 B.n422 B.n301 256.663
R462 B.n422 B.n302 256.663
R463 B.n422 B.n303 256.663
R464 B.n422 B.n304 256.663
R465 B.n422 B.n305 256.663
R466 B.n422 B.n306 256.663
R467 B.n422 B.n307 256.663
R468 B.n422 B.n308 256.663
R469 B.n423 B.n422 256.663
R470 B.n314 B.t8 254.332
R471 B.n311 B.t4 254.332
R472 B.n101 B.t11 254.332
R473 B.n98 B.t15 254.332
R474 B.n430 B.n279 163.367
R475 B.n430 B.n277 163.367
R476 B.n434 B.n277 163.367
R477 B.n434 B.n271 163.367
R478 B.n442 B.n271 163.367
R479 B.n442 B.n269 163.367
R480 B.n446 B.n269 163.367
R481 B.n446 B.n263 163.367
R482 B.n454 B.n263 163.367
R483 B.n454 B.n261 163.367
R484 B.n458 B.n261 163.367
R485 B.n458 B.n255 163.367
R486 B.n466 B.n255 163.367
R487 B.n466 B.n253 163.367
R488 B.n470 B.n253 163.367
R489 B.n470 B.n247 163.367
R490 B.n478 B.n247 163.367
R491 B.n478 B.n245 163.367
R492 B.n482 B.n245 163.367
R493 B.n482 B.n239 163.367
R494 B.n490 B.n239 163.367
R495 B.n490 B.n237 163.367
R496 B.n494 B.n237 163.367
R497 B.n494 B.n231 163.367
R498 B.n502 B.n231 163.367
R499 B.n502 B.n229 163.367
R500 B.n506 B.n229 163.367
R501 B.n506 B.n223 163.367
R502 B.n515 B.n223 163.367
R503 B.n515 B.n221 163.367
R504 B.n519 B.n221 163.367
R505 B.n519 B.n216 163.367
R506 B.n528 B.n216 163.367
R507 B.n528 B.n214 163.367
R508 B.n532 B.n214 163.367
R509 B.n532 B.n2 163.367
R510 B.n661 B.n2 163.367
R511 B.n661 B.n3 163.367
R512 B.n657 B.n3 163.367
R513 B.n657 B.n9 163.367
R514 B.n653 B.n9 163.367
R515 B.n653 B.n11 163.367
R516 B.n649 B.n11 163.367
R517 B.n649 B.n15 163.367
R518 B.n645 B.n15 163.367
R519 B.n645 B.n17 163.367
R520 B.n641 B.n17 163.367
R521 B.n641 B.n23 163.367
R522 B.n637 B.n23 163.367
R523 B.n637 B.n25 163.367
R524 B.n633 B.n25 163.367
R525 B.n633 B.n30 163.367
R526 B.n629 B.n30 163.367
R527 B.n629 B.n32 163.367
R528 B.n625 B.n32 163.367
R529 B.n625 B.n37 163.367
R530 B.n621 B.n37 163.367
R531 B.n621 B.n39 163.367
R532 B.n617 B.n39 163.367
R533 B.n617 B.n44 163.367
R534 B.n613 B.n44 163.367
R535 B.n613 B.n46 163.367
R536 B.n609 B.n46 163.367
R537 B.n609 B.n51 163.367
R538 B.n605 B.n51 163.367
R539 B.n605 B.n53 163.367
R540 B.n601 B.n53 163.367
R541 B.n601 B.n58 163.367
R542 B.n597 B.n58 163.367
R543 B.n597 B.n60 163.367
R544 B.n593 B.n60 163.367
R545 B.n593 B.n65 163.367
R546 B.n589 B.n65 163.367
R547 B.n589 B.n67 163.367
R548 B.n310 B.n309 163.367
R549 B.n415 B.n309 163.367
R550 B.n413 B.n412 163.367
R551 B.n409 B.n408 163.367
R552 B.n405 B.n404 163.367
R553 B.n401 B.n400 163.367
R554 B.n397 B.n396 163.367
R555 B.n393 B.n392 163.367
R556 B.n389 B.n388 163.367
R557 B.n385 B.n384 163.367
R558 B.n381 B.n380 163.367
R559 B.n377 B.n376 163.367
R560 B.n373 B.n372 163.367
R561 B.n369 B.n368 163.367
R562 B.n365 B.n364 163.367
R563 B.n361 B.n360 163.367
R564 B.n356 B.n355 163.367
R565 B.n352 B.n351 163.367
R566 B.n348 B.n347 163.367
R567 B.n344 B.n343 163.367
R568 B.n340 B.n339 163.367
R569 B.n336 B.n335 163.367
R570 B.n332 B.n331 163.367
R571 B.n328 B.n327 163.367
R572 B.n324 B.n323 163.367
R573 B.n320 B.n319 163.367
R574 B.n316 B.n283 163.367
R575 B.n428 B.n281 163.367
R576 B.n428 B.n275 163.367
R577 B.n436 B.n275 163.367
R578 B.n436 B.n273 163.367
R579 B.n440 B.n273 163.367
R580 B.n440 B.n266 163.367
R581 B.n448 B.n266 163.367
R582 B.n448 B.n264 163.367
R583 B.n452 B.n264 163.367
R584 B.n452 B.n259 163.367
R585 B.n460 B.n259 163.367
R586 B.n460 B.n257 163.367
R587 B.n464 B.n257 163.367
R588 B.n464 B.n251 163.367
R589 B.n472 B.n251 163.367
R590 B.n472 B.n249 163.367
R591 B.n476 B.n249 163.367
R592 B.n476 B.n242 163.367
R593 B.n484 B.n242 163.367
R594 B.n484 B.n240 163.367
R595 B.n488 B.n240 163.367
R596 B.n488 B.n235 163.367
R597 B.n496 B.n235 163.367
R598 B.n496 B.n233 163.367
R599 B.n500 B.n233 163.367
R600 B.n500 B.n227 163.367
R601 B.n508 B.n227 163.367
R602 B.n508 B.n225 163.367
R603 B.n512 B.n225 163.367
R604 B.n512 B.n220 163.367
R605 B.n521 B.n220 163.367
R606 B.n521 B.n218 163.367
R607 B.n526 B.n218 163.367
R608 B.n526 B.n212 163.367
R609 B.n534 B.n212 163.367
R610 B.n535 B.n534 163.367
R611 B.n535 B.n5 163.367
R612 B.n6 B.n5 163.367
R613 B.n7 B.n6 163.367
R614 B.n540 B.n7 163.367
R615 B.n540 B.n12 163.367
R616 B.n13 B.n12 163.367
R617 B.n14 B.n13 163.367
R618 B.n545 B.n14 163.367
R619 B.n545 B.n19 163.367
R620 B.n20 B.n19 163.367
R621 B.n21 B.n20 163.367
R622 B.n550 B.n21 163.367
R623 B.n550 B.n26 163.367
R624 B.n27 B.n26 163.367
R625 B.n28 B.n27 163.367
R626 B.n555 B.n28 163.367
R627 B.n555 B.n33 163.367
R628 B.n34 B.n33 163.367
R629 B.n35 B.n34 163.367
R630 B.n560 B.n35 163.367
R631 B.n560 B.n40 163.367
R632 B.n41 B.n40 163.367
R633 B.n42 B.n41 163.367
R634 B.n565 B.n42 163.367
R635 B.n565 B.n47 163.367
R636 B.n48 B.n47 163.367
R637 B.n49 B.n48 163.367
R638 B.n570 B.n49 163.367
R639 B.n570 B.n54 163.367
R640 B.n55 B.n54 163.367
R641 B.n56 B.n55 163.367
R642 B.n575 B.n56 163.367
R643 B.n575 B.n61 163.367
R644 B.n62 B.n61 163.367
R645 B.n63 B.n62 163.367
R646 B.n580 B.n63 163.367
R647 B.n580 B.n68 163.367
R648 B.n69 B.n68 163.367
R649 B.n107 B.n106 163.367
R650 B.n111 B.n110 163.367
R651 B.n115 B.n114 163.367
R652 B.n119 B.n118 163.367
R653 B.n123 B.n122 163.367
R654 B.n127 B.n126 163.367
R655 B.n131 B.n130 163.367
R656 B.n135 B.n134 163.367
R657 B.n139 B.n138 163.367
R658 B.n143 B.n142 163.367
R659 B.n147 B.n146 163.367
R660 B.n152 B.n151 163.367
R661 B.n156 B.n155 163.367
R662 B.n160 B.n159 163.367
R663 B.n164 B.n163 163.367
R664 B.n168 B.n167 163.367
R665 B.n172 B.n171 163.367
R666 B.n176 B.n175 163.367
R667 B.n180 B.n179 163.367
R668 B.n184 B.n183 163.367
R669 B.n188 B.n187 163.367
R670 B.n192 B.n191 163.367
R671 B.n196 B.n195 163.367
R672 B.n200 B.n199 163.367
R673 B.n204 B.n203 163.367
R674 B.n208 B.n207 163.367
R675 B.n585 B.n97 163.367
R676 B.n314 B.t10 136.034
R677 B.n98 B.t16 136.034
R678 B.n311 B.t7 136.028
R679 B.n101 B.t13 136.028
R680 B.n422 B.n280 122.504
R681 B.n587 B.n586 122.504
R682 B.n315 B.t9 72.6155
R683 B.n99 B.t17 72.6155
R684 B.n312 B.t6 72.6097
R685 B.n102 B.t14 72.6097
R686 B.n421 B.n420 71.676
R687 B.n415 B.n284 71.676
R688 B.n412 B.n285 71.676
R689 B.n408 B.n286 71.676
R690 B.n404 B.n287 71.676
R691 B.n400 B.n288 71.676
R692 B.n396 B.n289 71.676
R693 B.n392 B.n290 71.676
R694 B.n388 B.n291 71.676
R695 B.n384 B.n292 71.676
R696 B.n380 B.n293 71.676
R697 B.n376 B.n294 71.676
R698 B.n372 B.n295 71.676
R699 B.n368 B.n296 71.676
R700 B.n364 B.n297 71.676
R701 B.n360 B.n298 71.676
R702 B.n355 B.n299 71.676
R703 B.n351 B.n300 71.676
R704 B.n347 B.n301 71.676
R705 B.n343 B.n302 71.676
R706 B.n339 B.n303 71.676
R707 B.n335 B.n304 71.676
R708 B.n331 B.n305 71.676
R709 B.n327 B.n306 71.676
R710 B.n323 B.n307 71.676
R711 B.n319 B.n308 71.676
R712 B.n423 B.n283 71.676
R713 B.n103 B.n70 71.676
R714 B.n107 B.n71 71.676
R715 B.n111 B.n72 71.676
R716 B.n115 B.n73 71.676
R717 B.n119 B.n74 71.676
R718 B.n123 B.n75 71.676
R719 B.n127 B.n76 71.676
R720 B.n131 B.n77 71.676
R721 B.n135 B.n78 71.676
R722 B.n139 B.n79 71.676
R723 B.n143 B.n80 71.676
R724 B.n147 B.n81 71.676
R725 B.n152 B.n82 71.676
R726 B.n156 B.n83 71.676
R727 B.n160 B.n84 71.676
R728 B.n164 B.n85 71.676
R729 B.n168 B.n86 71.676
R730 B.n172 B.n87 71.676
R731 B.n176 B.n88 71.676
R732 B.n180 B.n89 71.676
R733 B.n184 B.n90 71.676
R734 B.n188 B.n91 71.676
R735 B.n192 B.n92 71.676
R736 B.n196 B.n93 71.676
R737 B.n200 B.n94 71.676
R738 B.n204 B.n95 71.676
R739 B.n208 B.n96 71.676
R740 B.n97 B.n96 71.676
R741 B.n207 B.n95 71.676
R742 B.n203 B.n94 71.676
R743 B.n199 B.n93 71.676
R744 B.n195 B.n92 71.676
R745 B.n191 B.n91 71.676
R746 B.n187 B.n90 71.676
R747 B.n183 B.n89 71.676
R748 B.n179 B.n88 71.676
R749 B.n175 B.n87 71.676
R750 B.n171 B.n86 71.676
R751 B.n167 B.n85 71.676
R752 B.n163 B.n84 71.676
R753 B.n159 B.n83 71.676
R754 B.n155 B.n82 71.676
R755 B.n151 B.n81 71.676
R756 B.n146 B.n80 71.676
R757 B.n142 B.n79 71.676
R758 B.n138 B.n78 71.676
R759 B.n134 B.n77 71.676
R760 B.n130 B.n76 71.676
R761 B.n126 B.n75 71.676
R762 B.n122 B.n74 71.676
R763 B.n118 B.n73 71.676
R764 B.n114 B.n72 71.676
R765 B.n110 B.n71 71.676
R766 B.n106 B.n70 71.676
R767 B.n421 B.n310 71.676
R768 B.n413 B.n284 71.676
R769 B.n409 B.n285 71.676
R770 B.n405 B.n286 71.676
R771 B.n401 B.n287 71.676
R772 B.n397 B.n288 71.676
R773 B.n393 B.n289 71.676
R774 B.n389 B.n290 71.676
R775 B.n385 B.n291 71.676
R776 B.n381 B.n292 71.676
R777 B.n377 B.n293 71.676
R778 B.n373 B.n294 71.676
R779 B.n369 B.n295 71.676
R780 B.n365 B.n296 71.676
R781 B.n361 B.n297 71.676
R782 B.n356 B.n298 71.676
R783 B.n352 B.n299 71.676
R784 B.n348 B.n300 71.676
R785 B.n344 B.n301 71.676
R786 B.n340 B.n302 71.676
R787 B.n336 B.n303 71.676
R788 B.n332 B.n304 71.676
R789 B.n328 B.n305 71.676
R790 B.n324 B.n306 71.676
R791 B.n320 B.n307 71.676
R792 B.n316 B.n308 71.676
R793 B.n424 B.n423 71.676
R794 B.n429 B.n280 68.8454
R795 B.n429 B.n276 68.8454
R796 B.n435 B.n276 68.8454
R797 B.n435 B.n272 68.8454
R798 B.n441 B.n272 68.8454
R799 B.n441 B.n267 68.8454
R800 B.n447 B.n267 68.8454
R801 B.n447 B.n268 68.8454
R802 B.n453 B.n260 68.8454
R803 B.n459 B.n260 68.8454
R804 B.n459 B.n256 68.8454
R805 B.n465 B.n256 68.8454
R806 B.n465 B.n252 68.8454
R807 B.n471 B.n252 68.8454
R808 B.n471 B.n248 68.8454
R809 B.n477 B.n248 68.8454
R810 B.n477 B.n243 68.8454
R811 B.n483 B.n243 68.8454
R812 B.n483 B.n244 68.8454
R813 B.n489 B.n236 68.8454
R814 B.n495 B.n236 68.8454
R815 B.n495 B.n232 68.8454
R816 B.n501 B.n232 68.8454
R817 B.n501 B.n228 68.8454
R818 B.n507 B.n228 68.8454
R819 B.n507 B.n224 68.8454
R820 B.n514 B.n224 68.8454
R821 B.n514 B.n513 68.8454
R822 B.n520 B.n217 68.8454
R823 B.n527 B.n217 68.8454
R824 B.n527 B.n213 68.8454
R825 B.n533 B.n213 68.8454
R826 B.n533 B.n4 68.8454
R827 B.n660 B.n4 68.8454
R828 B.n660 B.n659 68.8454
R829 B.n659 B.n658 68.8454
R830 B.n658 B.n8 68.8454
R831 B.n652 B.n8 68.8454
R832 B.n652 B.n651 68.8454
R833 B.n651 B.n650 68.8454
R834 B.n644 B.n18 68.8454
R835 B.n644 B.n643 68.8454
R836 B.n643 B.n642 68.8454
R837 B.n642 B.n22 68.8454
R838 B.n636 B.n22 68.8454
R839 B.n636 B.n635 68.8454
R840 B.n635 B.n634 68.8454
R841 B.n634 B.n29 68.8454
R842 B.n628 B.n29 68.8454
R843 B.n627 B.n626 68.8454
R844 B.n626 B.n36 68.8454
R845 B.n620 B.n36 68.8454
R846 B.n620 B.n619 68.8454
R847 B.n619 B.n618 68.8454
R848 B.n618 B.n43 68.8454
R849 B.n612 B.n43 68.8454
R850 B.n612 B.n611 68.8454
R851 B.n611 B.n610 68.8454
R852 B.n610 B.n50 68.8454
R853 B.n604 B.n50 68.8454
R854 B.n603 B.n602 68.8454
R855 B.n602 B.n57 68.8454
R856 B.n596 B.n57 68.8454
R857 B.n596 B.n595 68.8454
R858 B.n595 B.n594 68.8454
R859 B.n594 B.n64 68.8454
R860 B.n588 B.n64 68.8454
R861 B.n588 B.n587 68.8454
R862 B.n244 B.t0 66.8206
R863 B.t1 B.n627 66.8206
R864 B.n315 B.n314 63.4187
R865 B.n312 B.n311 63.4187
R866 B.n102 B.n101 63.4187
R867 B.n99 B.n98 63.4187
R868 B.n358 B.n315 59.5399
R869 B.n313 B.n312 59.5399
R870 B.n149 B.n102 59.5399
R871 B.n100 B.n99 59.5399
R872 B.n453 B.t5 58.7212
R873 B.n604 B.t12 58.7212
R874 B.n513 B.t3 40.4975
R875 B.n18 B.t2 40.4975
R876 B.n104 B.n66 32.6249
R877 B.n584 B.n583 32.6249
R878 B.n426 B.n425 32.6249
R879 B.n419 B.n278 32.6249
R880 B.n520 B.t3 28.3484
R881 B.n650 B.t2 28.3484
R882 B B.n662 18.0485
R883 B.n105 B.n104 10.6151
R884 B.n108 B.n105 10.6151
R885 B.n109 B.n108 10.6151
R886 B.n112 B.n109 10.6151
R887 B.n113 B.n112 10.6151
R888 B.n116 B.n113 10.6151
R889 B.n117 B.n116 10.6151
R890 B.n120 B.n117 10.6151
R891 B.n121 B.n120 10.6151
R892 B.n124 B.n121 10.6151
R893 B.n125 B.n124 10.6151
R894 B.n128 B.n125 10.6151
R895 B.n129 B.n128 10.6151
R896 B.n132 B.n129 10.6151
R897 B.n133 B.n132 10.6151
R898 B.n136 B.n133 10.6151
R899 B.n137 B.n136 10.6151
R900 B.n140 B.n137 10.6151
R901 B.n141 B.n140 10.6151
R902 B.n144 B.n141 10.6151
R903 B.n145 B.n144 10.6151
R904 B.n148 B.n145 10.6151
R905 B.n153 B.n150 10.6151
R906 B.n154 B.n153 10.6151
R907 B.n157 B.n154 10.6151
R908 B.n158 B.n157 10.6151
R909 B.n161 B.n158 10.6151
R910 B.n162 B.n161 10.6151
R911 B.n165 B.n162 10.6151
R912 B.n166 B.n165 10.6151
R913 B.n170 B.n169 10.6151
R914 B.n173 B.n170 10.6151
R915 B.n174 B.n173 10.6151
R916 B.n177 B.n174 10.6151
R917 B.n178 B.n177 10.6151
R918 B.n181 B.n178 10.6151
R919 B.n182 B.n181 10.6151
R920 B.n185 B.n182 10.6151
R921 B.n186 B.n185 10.6151
R922 B.n189 B.n186 10.6151
R923 B.n190 B.n189 10.6151
R924 B.n193 B.n190 10.6151
R925 B.n194 B.n193 10.6151
R926 B.n197 B.n194 10.6151
R927 B.n198 B.n197 10.6151
R928 B.n201 B.n198 10.6151
R929 B.n202 B.n201 10.6151
R930 B.n205 B.n202 10.6151
R931 B.n206 B.n205 10.6151
R932 B.n209 B.n206 10.6151
R933 B.n210 B.n209 10.6151
R934 B.n584 B.n210 10.6151
R935 B.n427 B.n426 10.6151
R936 B.n427 B.n274 10.6151
R937 B.n437 B.n274 10.6151
R938 B.n438 B.n437 10.6151
R939 B.n439 B.n438 10.6151
R940 B.n439 B.n265 10.6151
R941 B.n449 B.n265 10.6151
R942 B.n450 B.n449 10.6151
R943 B.n451 B.n450 10.6151
R944 B.n451 B.n258 10.6151
R945 B.n461 B.n258 10.6151
R946 B.n462 B.n461 10.6151
R947 B.n463 B.n462 10.6151
R948 B.n463 B.n250 10.6151
R949 B.n473 B.n250 10.6151
R950 B.n474 B.n473 10.6151
R951 B.n475 B.n474 10.6151
R952 B.n475 B.n241 10.6151
R953 B.n485 B.n241 10.6151
R954 B.n486 B.n485 10.6151
R955 B.n487 B.n486 10.6151
R956 B.n487 B.n234 10.6151
R957 B.n497 B.n234 10.6151
R958 B.n498 B.n497 10.6151
R959 B.n499 B.n498 10.6151
R960 B.n499 B.n226 10.6151
R961 B.n509 B.n226 10.6151
R962 B.n510 B.n509 10.6151
R963 B.n511 B.n510 10.6151
R964 B.n511 B.n219 10.6151
R965 B.n522 B.n219 10.6151
R966 B.n523 B.n522 10.6151
R967 B.n525 B.n523 10.6151
R968 B.n525 B.n524 10.6151
R969 B.n524 B.n211 10.6151
R970 B.n536 B.n211 10.6151
R971 B.n537 B.n536 10.6151
R972 B.n538 B.n537 10.6151
R973 B.n539 B.n538 10.6151
R974 B.n541 B.n539 10.6151
R975 B.n542 B.n541 10.6151
R976 B.n543 B.n542 10.6151
R977 B.n544 B.n543 10.6151
R978 B.n546 B.n544 10.6151
R979 B.n547 B.n546 10.6151
R980 B.n548 B.n547 10.6151
R981 B.n549 B.n548 10.6151
R982 B.n551 B.n549 10.6151
R983 B.n552 B.n551 10.6151
R984 B.n553 B.n552 10.6151
R985 B.n554 B.n553 10.6151
R986 B.n556 B.n554 10.6151
R987 B.n557 B.n556 10.6151
R988 B.n558 B.n557 10.6151
R989 B.n559 B.n558 10.6151
R990 B.n561 B.n559 10.6151
R991 B.n562 B.n561 10.6151
R992 B.n563 B.n562 10.6151
R993 B.n564 B.n563 10.6151
R994 B.n566 B.n564 10.6151
R995 B.n567 B.n566 10.6151
R996 B.n568 B.n567 10.6151
R997 B.n569 B.n568 10.6151
R998 B.n571 B.n569 10.6151
R999 B.n572 B.n571 10.6151
R1000 B.n573 B.n572 10.6151
R1001 B.n574 B.n573 10.6151
R1002 B.n576 B.n574 10.6151
R1003 B.n577 B.n576 10.6151
R1004 B.n578 B.n577 10.6151
R1005 B.n579 B.n578 10.6151
R1006 B.n581 B.n579 10.6151
R1007 B.n582 B.n581 10.6151
R1008 B.n583 B.n582 10.6151
R1009 B.n419 B.n418 10.6151
R1010 B.n418 B.n417 10.6151
R1011 B.n417 B.n416 10.6151
R1012 B.n416 B.n414 10.6151
R1013 B.n414 B.n411 10.6151
R1014 B.n411 B.n410 10.6151
R1015 B.n410 B.n407 10.6151
R1016 B.n407 B.n406 10.6151
R1017 B.n406 B.n403 10.6151
R1018 B.n403 B.n402 10.6151
R1019 B.n402 B.n399 10.6151
R1020 B.n399 B.n398 10.6151
R1021 B.n398 B.n395 10.6151
R1022 B.n395 B.n394 10.6151
R1023 B.n394 B.n391 10.6151
R1024 B.n391 B.n390 10.6151
R1025 B.n390 B.n387 10.6151
R1026 B.n387 B.n386 10.6151
R1027 B.n386 B.n383 10.6151
R1028 B.n383 B.n382 10.6151
R1029 B.n382 B.n379 10.6151
R1030 B.n379 B.n378 10.6151
R1031 B.n375 B.n374 10.6151
R1032 B.n374 B.n371 10.6151
R1033 B.n371 B.n370 10.6151
R1034 B.n370 B.n367 10.6151
R1035 B.n367 B.n366 10.6151
R1036 B.n366 B.n363 10.6151
R1037 B.n363 B.n362 10.6151
R1038 B.n362 B.n359 10.6151
R1039 B.n357 B.n354 10.6151
R1040 B.n354 B.n353 10.6151
R1041 B.n353 B.n350 10.6151
R1042 B.n350 B.n349 10.6151
R1043 B.n349 B.n346 10.6151
R1044 B.n346 B.n345 10.6151
R1045 B.n345 B.n342 10.6151
R1046 B.n342 B.n341 10.6151
R1047 B.n341 B.n338 10.6151
R1048 B.n338 B.n337 10.6151
R1049 B.n337 B.n334 10.6151
R1050 B.n334 B.n333 10.6151
R1051 B.n333 B.n330 10.6151
R1052 B.n330 B.n329 10.6151
R1053 B.n329 B.n326 10.6151
R1054 B.n326 B.n325 10.6151
R1055 B.n325 B.n322 10.6151
R1056 B.n322 B.n321 10.6151
R1057 B.n321 B.n318 10.6151
R1058 B.n318 B.n317 10.6151
R1059 B.n317 B.n282 10.6151
R1060 B.n425 B.n282 10.6151
R1061 B.n431 B.n278 10.6151
R1062 B.n432 B.n431 10.6151
R1063 B.n433 B.n432 10.6151
R1064 B.n433 B.n270 10.6151
R1065 B.n443 B.n270 10.6151
R1066 B.n444 B.n443 10.6151
R1067 B.n445 B.n444 10.6151
R1068 B.n445 B.n262 10.6151
R1069 B.n455 B.n262 10.6151
R1070 B.n456 B.n455 10.6151
R1071 B.n457 B.n456 10.6151
R1072 B.n457 B.n254 10.6151
R1073 B.n467 B.n254 10.6151
R1074 B.n468 B.n467 10.6151
R1075 B.n469 B.n468 10.6151
R1076 B.n469 B.n246 10.6151
R1077 B.n479 B.n246 10.6151
R1078 B.n480 B.n479 10.6151
R1079 B.n481 B.n480 10.6151
R1080 B.n481 B.n238 10.6151
R1081 B.n491 B.n238 10.6151
R1082 B.n492 B.n491 10.6151
R1083 B.n493 B.n492 10.6151
R1084 B.n493 B.n230 10.6151
R1085 B.n503 B.n230 10.6151
R1086 B.n504 B.n503 10.6151
R1087 B.n505 B.n504 10.6151
R1088 B.n505 B.n222 10.6151
R1089 B.n516 B.n222 10.6151
R1090 B.n517 B.n516 10.6151
R1091 B.n518 B.n517 10.6151
R1092 B.n518 B.n215 10.6151
R1093 B.n529 B.n215 10.6151
R1094 B.n530 B.n529 10.6151
R1095 B.n531 B.n530 10.6151
R1096 B.n531 B.n0 10.6151
R1097 B.n656 B.n1 10.6151
R1098 B.n656 B.n655 10.6151
R1099 B.n655 B.n654 10.6151
R1100 B.n654 B.n10 10.6151
R1101 B.n648 B.n10 10.6151
R1102 B.n648 B.n647 10.6151
R1103 B.n647 B.n646 10.6151
R1104 B.n646 B.n16 10.6151
R1105 B.n640 B.n16 10.6151
R1106 B.n640 B.n639 10.6151
R1107 B.n639 B.n638 10.6151
R1108 B.n638 B.n24 10.6151
R1109 B.n632 B.n24 10.6151
R1110 B.n632 B.n631 10.6151
R1111 B.n631 B.n630 10.6151
R1112 B.n630 B.n31 10.6151
R1113 B.n624 B.n31 10.6151
R1114 B.n624 B.n623 10.6151
R1115 B.n623 B.n622 10.6151
R1116 B.n622 B.n38 10.6151
R1117 B.n616 B.n38 10.6151
R1118 B.n616 B.n615 10.6151
R1119 B.n615 B.n614 10.6151
R1120 B.n614 B.n45 10.6151
R1121 B.n608 B.n45 10.6151
R1122 B.n608 B.n607 10.6151
R1123 B.n607 B.n606 10.6151
R1124 B.n606 B.n52 10.6151
R1125 B.n600 B.n52 10.6151
R1126 B.n600 B.n599 10.6151
R1127 B.n599 B.n598 10.6151
R1128 B.n598 B.n59 10.6151
R1129 B.n592 B.n59 10.6151
R1130 B.n592 B.n591 10.6151
R1131 B.n591 B.n590 10.6151
R1132 B.n590 B.n66 10.6151
R1133 B.n268 B.t5 10.1248
R1134 B.t12 B.n603 10.1248
R1135 B.n150 B.n149 6.5566
R1136 B.n166 B.n100 6.5566
R1137 B.n375 B.n313 6.5566
R1138 B.n359 B.n358 6.5566
R1139 B.n149 B.n148 4.05904
R1140 B.n169 B.n100 4.05904
R1141 B.n378 B.n313 4.05904
R1142 B.n358 B.n357 4.05904
R1143 B.n662 B.n0 2.81026
R1144 B.n662 B.n1 2.81026
R1145 B.n489 B.t0 2.02535
R1146 B.n628 B.t1 2.02535
R1147 VN.n1 VN.t2 80.1836
R1148 VN.n0 VN.t0 80.1836
R1149 VN.n0 VN.t3 79.2059
R1150 VN.n1 VN.t1 79.2059
R1151 VN VN.n1 45.7807
R1152 VN VN.n0 3.11784
R1153 VDD2.n2 VDD2.n0 103.891
R1154 VDD2.n2 VDD2.n1 66.9002
R1155 VDD2.n1 VDD2.t3 3.54254
R1156 VDD2.n1 VDD2.t1 3.54254
R1157 VDD2.n0 VDD2.t2 3.54254
R1158 VDD2.n0 VDD2.t0 3.54254
R1159 VDD2 VDD2.n2 0.0586897
R1160 VTAIL.n5 VTAIL.t2 53.7636
R1161 VTAIL.n4 VTAIL.t5 53.7636
R1162 VTAIL.n3 VTAIL.t6 53.7636
R1163 VTAIL.n7 VTAIL.t4 53.7634
R1164 VTAIL.n0 VTAIL.t7 53.7634
R1165 VTAIL.n1 VTAIL.t3 53.7634
R1166 VTAIL.n2 VTAIL.t0 53.7634
R1167 VTAIL.n6 VTAIL.t1 53.7634
R1168 VTAIL.n7 VTAIL.n6 20.0048
R1169 VTAIL.n3 VTAIL.n2 20.0048
R1170 VTAIL.n4 VTAIL.n3 2.81947
R1171 VTAIL.n6 VTAIL.n5 2.81947
R1172 VTAIL.n2 VTAIL.n1 2.81947
R1173 VTAIL VTAIL.n0 1.46817
R1174 VTAIL VTAIL.n7 1.35179
R1175 VTAIL.n5 VTAIL.n4 0.470328
R1176 VTAIL.n1 VTAIL.n0 0.470328
R1177 VP.n15 VP.n14 161.3
R1178 VP.n13 VP.n1 161.3
R1179 VP.n12 VP.n11 161.3
R1180 VP.n10 VP.n2 161.3
R1181 VP.n9 VP.n8 161.3
R1182 VP.n7 VP.n3 161.3
R1183 VP.n4 VP.t3 80.1833
R1184 VP.n4 VP.t0 79.206
R1185 VP.n6 VP.n5 71.2278
R1186 VP.n16 VP.n0 71.2278
R1187 VP.n12 VP.n2 56.5193
R1188 VP.n6 VP.t2 45.8233
R1189 VP.n0 VP.t1 45.8233
R1190 VP.n5 VP.n4 45.6153
R1191 VP.n8 VP.n7 24.4675
R1192 VP.n8 VP.n2 24.4675
R1193 VP.n13 VP.n12 24.4675
R1194 VP.n14 VP.n13 24.4675
R1195 VP.n7 VP.n6 18.8401
R1196 VP.n14 VP.n0 18.8401
R1197 VP.n5 VP.n3 0.354971
R1198 VP.n16 VP.n15 0.354971
R1199 VP VP.n16 0.26696
R1200 VP.n9 VP.n3 0.189894
R1201 VP.n10 VP.n9 0.189894
R1202 VP.n11 VP.n10 0.189894
R1203 VP.n11 VP.n1 0.189894
R1204 VP.n15 VP.n1 0.189894
R1205 VDD1 VDD1.n1 104.415
R1206 VDD1 VDD1.n0 66.9584
R1207 VDD1.n0 VDD1.t0 3.54254
R1208 VDD1.n0 VDD1.t3 3.54254
R1209 VDD1.n1 VDD1.t1 3.54254
R1210 VDD1.n1 VDD1.t2 3.54254
C0 VP VTAIL 2.83145f
C1 VDD2 VN 2.4307f
C2 VTAIL VDD1 4.01938f
C3 VP VN 5.25271f
C4 VDD1 VN 0.149448f
C5 VP VDD2 0.416081f
C6 VDD1 VDD2 1.10789f
C7 VP VDD1 2.69651f
C8 VTAIL VN 2.81734f
C9 VTAIL VDD2 4.075861f
C10 VDD2 B 3.470067f
C11 VDD1 B 7.13461f
C12 VTAIL B 6.122786f
C13 VN B 10.79484f
C14 VP B 9.103848f
C15 VDD1.t0 B 0.125067f
C16 VDD1.t3 B 0.125067f
C17 VDD1.n0 B 1.034f
C18 VDD1.t1 B 0.125067f
C19 VDD1.t2 B 0.125067f
C20 VDD1.n1 B 1.53441f
C21 VP.t1 B 1.2116f
C22 VP.n0 B 0.561604f
C23 VP.n1 B 0.027974f
C24 VP.n2 B 0.040837f
C25 VP.n3 B 0.04515f
C26 VP.t2 B 1.2116f
C27 VP.t3 B 1.49034f
C28 VP.t0 B 1.48252f
C29 VP.n4 B 2.31968f
C30 VP.n5 B 1.36911f
C31 VP.n6 B 0.561604f
C32 VP.n7 B 0.046216f
C33 VP.n8 B 0.052137f
C34 VP.n9 B 0.027974f
C35 VP.n10 B 0.027974f
C36 VP.n11 B 0.027974f
C37 VP.n12 B 0.040837f
C38 VP.n13 B 0.052137f
C39 VP.n14 B 0.046216f
C40 VP.n15 B 0.04515f
C41 VP.n16 B 0.059071f
C42 VTAIL.t7 B 0.878611f
C43 VTAIL.n0 B 0.372328f
C44 VTAIL.t3 B 0.878611f
C45 VTAIL.n1 B 0.460882f
C46 VTAIL.t0 B 0.878611f
C47 VTAIL.n2 B 1.2069f
C48 VTAIL.t6 B 0.878615f
C49 VTAIL.n3 B 1.20689f
C50 VTAIL.t5 B 0.878615f
C51 VTAIL.n4 B 0.460879f
C52 VTAIL.t2 B 0.878615f
C53 VTAIL.n5 B 0.460879f
C54 VTAIL.t1 B 0.878611f
C55 VTAIL.n6 B 1.2069f
C56 VTAIL.t4 B 0.878611f
C57 VTAIL.n7 B 1.11071f
C58 VDD2.t2 B 0.123257f
C59 VDD2.t0 B 0.123257f
C60 VDD2.n0 B 1.48782f
C61 VDD2.t3 B 0.123257f
C62 VDD2.t1 B 0.123257f
C63 VDD2.n1 B 1.01861f
C64 VDD2.n2 B 3.24108f
C65 VN.t3 B 1.43611f
C66 VN.t0 B 1.44368f
C67 VN.n0 B 0.884571f
C68 VN.t2 B 1.44368f
C69 VN.t1 B 1.43611f
C70 VN.n1 B 2.25841f
.ends

