* NGSPICE file created from diff_pair_sample_0755.ext - technology: sky130A

.subckt diff_pair_sample_0755 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.6747 pd=4.24 as=0.6747 ps=4.24 w=1.73 l=2.19
X1 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=0.6747 pd=4.24 as=0 ps=0 w=1.73 l=2.19
X2 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.6747 pd=4.24 as=0.6747 ps=4.24 w=1.73 l=2.19
X3 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=0.6747 pd=4.24 as=0 ps=0 w=1.73 l=2.19
X4 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.6747 pd=4.24 as=0 ps=0 w=1.73 l=2.19
X5 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.6747 pd=4.24 as=0.6747 ps=4.24 w=1.73 l=2.19
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.6747 pd=4.24 as=0 ps=0 w=1.73 l=2.19
X7 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.6747 pd=4.24 as=0.6747 ps=4.24 w=1.73 l=2.19
R0 VP.n0 VP.t1 103.998
R1 VP.n0 VP.t0 68.2087
R2 VP VP.n0 0.336784
R3 VTAIL.n26 VTAIL.n24 289.615
R4 VTAIL.n2 VTAIL.n0 289.615
R5 VTAIL.n18 VTAIL.n16 289.615
R6 VTAIL.n10 VTAIL.n8 289.615
R7 VTAIL.n27 VTAIL.n26 185
R8 VTAIL.n3 VTAIL.n2 185
R9 VTAIL.n19 VTAIL.n18 185
R10 VTAIL.n11 VTAIL.n10 185
R11 VTAIL.t3 VTAIL.n25 164.876
R12 VTAIL.t2 VTAIL.n1 164.876
R13 VTAIL.t1 VTAIL.n17 164.876
R14 VTAIL.t0 VTAIL.n9 164.876
R15 VTAIL.n26 VTAIL.t3 52.3082
R16 VTAIL.n2 VTAIL.t2 52.3082
R17 VTAIL.n18 VTAIL.t1 52.3082
R18 VTAIL.n10 VTAIL.t0 52.3082
R19 VTAIL.n31 VTAIL.n30 33.155
R20 VTAIL.n7 VTAIL.n6 33.155
R21 VTAIL.n23 VTAIL.n22 33.155
R22 VTAIL.n15 VTAIL.n14 33.155
R23 VTAIL.n15 VTAIL.n7 18.2031
R24 VTAIL.n31 VTAIL.n23 16.0307
R25 VTAIL.n27 VTAIL.n25 14.7318
R26 VTAIL.n3 VTAIL.n1 14.7318
R27 VTAIL.n19 VTAIL.n17 14.7318
R28 VTAIL.n11 VTAIL.n9 14.7318
R29 VTAIL.n28 VTAIL.n24 12.8005
R30 VTAIL.n4 VTAIL.n0 12.8005
R31 VTAIL.n20 VTAIL.n16 12.8005
R32 VTAIL.n12 VTAIL.n8 12.8005
R33 VTAIL.n30 VTAIL.n29 9.45567
R34 VTAIL.n6 VTAIL.n5 9.45567
R35 VTAIL.n22 VTAIL.n21 9.45567
R36 VTAIL.n14 VTAIL.n13 9.45567
R37 VTAIL.n29 VTAIL.n28 9.3005
R38 VTAIL.n5 VTAIL.n4 9.3005
R39 VTAIL.n21 VTAIL.n20 9.3005
R40 VTAIL.n13 VTAIL.n12 9.3005
R41 VTAIL.n29 VTAIL.n25 5.62509
R42 VTAIL.n5 VTAIL.n1 5.62509
R43 VTAIL.n21 VTAIL.n17 5.62509
R44 VTAIL.n13 VTAIL.n9 5.62509
R45 VTAIL.n23 VTAIL.n15 1.55653
R46 VTAIL.n30 VTAIL.n24 1.16414
R47 VTAIL.n6 VTAIL.n0 1.16414
R48 VTAIL.n22 VTAIL.n16 1.16414
R49 VTAIL.n14 VTAIL.n8 1.16414
R50 VTAIL VTAIL.n7 1.07162
R51 VTAIL VTAIL.n31 0.485414
R52 VTAIL.n28 VTAIL.n27 0.388379
R53 VTAIL.n4 VTAIL.n3 0.388379
R54 VTAIL.n20 VTAIL.n19 0.388379
R55 VTAIL.n12 VTAIL.n11 0.388379
R56 VDD1.n2 VDD1.n0 289.615
R57 VDD1.n9 VDD1.n7 289.615
R58 VDD1.n3 VDD1.n2 185
R59 VDD1.n10 VDD1.n9 185
R60 VDD1.t0 VDD1.n1 164.876
R61 VDD1.t1 VDD1.n8 164.876
R62 VDD1 VDD1.n13 80.3974
R63 VDD1.n2 VDD1.t0 52.3082
R64 VDD1.n9 VDD1.t1 52.3082
R65 VDD1 VDD1.n6 50.4351
R66 VDD1.n3 VDD1.n1 14.7318
R67 VDD1.n10 VDD1.n8 14.7318
R68 VDD1.n4 VDD1.n0 12.8005
R69 VDD1.n11 VDD1.n7 12.8005
R70 VDD1.n6 VDD1.n5 9.45567
R71 VDD1.n13 VDD1.n12 9.45567
R72 VDD1.n5 VDD1.n4 9.3005
R73 VDD1.n12 VDD1.n11 9.3005
R74 VDD1.n5 VDD1.n1 5.62509
R75 VDD1.n12 VDD1.n8 5.62509
R76 VDD1.n6 VDD1.n0 1.16414
R77 VDD1.n13 VDD1.n7 1.16414
R78 VDD1.n4 VDD1.n3 0.388379
R79 VDD1.n11 VDD1.n10 0.388379
R80 B.n354 B.n353 585
R81 B.n125 B.n61 585
R82 B.n124 B.n123 585
R83 B.n122 B.n121 585
R84 B.n120 B.n119 585
R85 B.n118 B.n117 585
R86 B.n116 B.n115 585
R87 B.n114 B.n113 585
R88 B.n112 B.n111 585
R89 B.n110 B.n109 585
R90 B.n108 B.n107 585
R91 B.n105 B.n104 585
R92 B.n103 B.n102 585
R93 B.n101 B.n100 585
R94 B.n99 B.n98 585
R95 B.n97 B.n96 585
R96 B.n95 B.n94 585
R97 B.n93 B.n92 585
R98 B.n91 B.n90 585
R99 B.n89 B.n88 585
R100 B.n87 B.n86 585
R101 B.n84 B.n83 585
R102 B.n82 B.n81 585
R103 B.n80 B.n79 585
R104 B.n78 B.n77 585
R105 B.n76 B.n75 585
R106 B.n74 B.n73 585
R107 B.n72 B.n71 585
R108 B.n70 B.n69 585
R109 B.n68 B.n67 585
R110 B.n46 B.n45 585
R111 B.n359 B.n358 585
R112 B.n352 B.n62 585
R113 B.n62 B.n43 585
R114 B.n351 B.n42 585
R115 B.n363 B.n42 585
R116 B.n350 B.n41 585
R117 B.n364 B.n41 585
R118 B.n349 B.n40 585
R119 B.n365 B.n40 585
R120 B.n348 B.n347 585
R121 B.n347 B.n36 585
R122 B.n346 B.n35 585
R123 B.n371 B.n35 585
R124 B.n345 B.n34 585
R125 B.n372 B.n34 585
R126 B.n344 B.n33 585
R127 B.n373 B.n33 585
R128 B.n343 B.n342 585
R129 B.n342 B.n29 585
R130 B.n341 B.n28 585
R131 B.n379 B.n28 585
R132 B.n340 B.n27 585
R133 B.n380 B.n27 585
R134 B.n339 B.n26 585
R135 B.n381 B.n26 585
R136 B.n338 B.n337 585
R137 B.n337 B.n22 585
R138 B.n336 B.n21 585
R139 B.n387 B.n21 585
R140 B.n335 B.n20 585
R141 B.n388 B.n20 585
R142 B.n334 B.n19 585
R143 B.n389 B.n19 585
R144 B.n333 B.n332 585
R145 B.n332 B.n15 585
R146 B.n331 B.n14 585
R147 B.n395 B.n14 585
R148 B.n330 B.n13 585
R149 B.n396 B.n13 585
R150 B.n329 B.n12 585
R151 B.n397 B.n12 585
R152 B.n328 B.n327 585
R153 B.n327 B.n8 585
R154 B.n326 B.n7 585
R155 B.n403 B.n7 585
R156 B.n325 B.n6 585
R157 B.n404 B.n6 585
R158 B.n324 B.n5 585
R159 B.n405 B.n5 585
R160 B.n323 B.n322 585
R161 B.n322 B.n4 585
R162 B.n321 B.n126 585
R163 B.n321 B.n320 585
R164 B.n311 B.n127 585
R165 B.n128 B.n127 585
R166 B.n313 B.n312 585
R167 B.n314 B.n313 585
R168 B.n310 B.n133 585
R169 B.n133 B.n132 585
R170 B.n309 B.n308 585
R171 B.n308 B.n307 585
R172 B.n135 B.n134 585
R173 B.n136 B.n135 585
R174 B.n300 B.n299 585
R175 B.n301 B.n300 585
R176 B.n298 B.n141 585
R177 B.n141 B.n140 585
R178 B.n297 B.n296 585
R179 B.n296 B.n295 585
R180 B.n143 B.n142 585
R181 B.n144 B.n143 585
R182 B.n288 B.n287 585
R183 B.n289 B.n288 585
R184 B.n286 B.n149 585
R185 B.n149 B.n148 585
R186 B.n285 B.n284 585
R187 B.n284 B.n283 585
R188 B.n151 B.n150 585
R189 B.n152 B.n151 585
R190 B.n276 B.n275 585
R191 B.n277 B.n276 585
R192 B.n274 B.n157 585
R193 B.n157 B.n156 585
R194 B.n273 B.n272 585
R195 B.n272 B.n271 585
R196 B.n159 B.n158 585
R197 B.n160 B.n159 585
R198 B.n264 B.n263 585
R199 B.n265 B.n264 585
R200 B.n262 B.n165 585
R201 B.n165 B.n164 585
R202 B.n261 B.n260 585
R203 B.n260 B.n259 585
R204 B.n167 B.n166 585
R205 B.n168 B.n167 585
R206 B.n255 B.n254 585
R207 B.n171 B.n170 585
R208 B.n251 B.n250 585
R209 B.n252 B.n251 585
R210 B.n249 B.n187 585
R211 B.n248 B.n247 585
R212 B.n246 B.n245 585
R213 B.n244 B.n243 585
R214 B.n242 B.n241 585
R215 B.n240 B.n239 585
R216 B.n238 B.n237 585
R217 B.n236 B.n235 585
R218 B.n234 B.n233 585
R219 B.n232 B.n231 585
R220 B.n230 B.n229 585
R221 B.n228 B.n227 585
R222 B.n226 B.n225 585
R223 B.n224 B.n223 585
R224 B.n222 B.n221 585
R225 B.n220 B.n219 585
R226 B.n218 B.n217 585
R227 B.n216 B.n215 585
R228 B.n214 B.n213 585
R229 B.n212 B.n211 585
R230 B.n210 B.n209 585
R231 B.n208 B.n207 585
R232 B.n206 B.n205 585
R233 B.n204 B.n203 585
R234 B.n202 B.n201 585
R235 B.n200 B.n199 585
R236 B.n198 B.n197 585
R237 B.n196 B.n195 585
R238 B.n194 B.n186 585
R239 B.n252 B.n186 585
R240 B.n256 B.n169 585
R241 B.n169 B.n168 585
R242 B.n258 B.n257 585
R243 B.n259 B.n258 585
R244 B.n163 B.n162 585
R245 B.n164 B.n163 585
R246 B.n267 B.n266 585
R247 B.n266 B.n265 585
R248 B.n268 B.n161 585
R249 B.n161 B.n160 585
R250 B.n270 B.n269 585
R251 B.n271 B.n270 585
R252 B.n155 B.n154 585
R253 B.n156 B.n155 585
R254 B.n279 B.n278 585
R255 B.n278 B.n277 585
R256 B.n280 B.n153 585
R257 B.n153 B.n152 585
R258 B.n282 B.n281 585
R259 B.n283 B.n282 585
R260 B.n147 B.n146 585
R261 B.n148 B.n147 585
R262 B.n291 B.n290 585
R263 B.n290 B.n289 585
R264 B.n292 B.n145 585
R265 B.n145 B.n144 585
R266 B.n294 B.n293 585
R267 B.n295 B.n294 585
R268 B.n139 B.n138 585
R269 B.n140 B.n139 585
R270 B.n303 B.n302 585
R271 B.n302 B.n301 585
R272 B.n304 B.n137 585
R273 B.n137 B.n136 585
R274 B.n306 B.n305 585
R275 B.n307 B.n306 585
R276 B.n131 B.n130 585
R277 B.n132 B.n131 585
R278 B.n316 B.n315 585
R279 B.n315 B.n314 585
R280 B.n317 B.n129 585
R281 B.n129 B.n128 585
R282 B.n319 B.n318 585
R283 B.n320 B.n319 585
R284 B.n2 B.n0 585
R285 B.n4 B.n2 585
R286 B.n3 B.n1 585
R287 B.n404 B.n3 585
R288 B.n402 B.n401 585
R289 B.n403 B.n402 585
R290 B.n400 B.n9 585
R291 B.n9 B.n8 585
R292 B.n399 B.n398 585
R293 B.n398 B.n397 585
R294 B.n11 B.n10 585
R295 B.n396 B.n11 585
R296 B.n394 B.n393 585
R297 B.n395 B.n394 585
R298 B.n392 B.n16 585
R299 B.n16 B.n15 585
R300 B.n391 B.n390 585
R301 B.n390 B.n389 585
R302 B.n18 B.n17 585
R303 B.n388 B.n18 585
R304 B.n386 B.n385 585
R305 B.n387 B.n386 585
R306 B.n384 B.n23 585
R307 B.n23 B.n22 585
R308 B.n383 B.n382 585
R309 B.n382 B.n381 585
R310 B.n25 B.n24 585
R311 B.n380 B.n25 585
R312 B.n378 B.n377 585
R313 B.n379 B.n378 585
R314 B.n376 B.n30 585
R315 B.n30 B.n29 585
R316 B.n375 B.n374 585
R317 B.n374 B.n373 585
R318 B.n32 B.n31 585
R319 B.n372 B.n32 585
R320 B.n370 B.n369 585
R321 B.n371 B.n370 585
R322 B.n368 B.n37 585
R323 B.n37 B.n36 585
R324 B.n367 B.n366 585
R325 B.n366 B.n365 585
R326 B.n39 B.n38 585
R327 B.n364 B.n39 585
R328 B.n362 B.n361 585
R329 B.n363 B.n362 585
R330 B.n360 B.n44 585
R331 B.n44 B.n43 585
R332 B.n407 B.n406 585
R333 B.n406 B.n405 585
R334 B.n254 B.n169 521.33
R335 B.n358 B.n44 521.33
R336 B.n186 B.n167 521.33
R337 B.n354 B.n62 521.33
R338 B.n356 B.n355 256.663
R339 B.n356 B.n60 256.663
R340 B.n356 B.n59 256.663
R341 B.n356 B.n58 256.663
R342 B.n356 B.n57 256.663
R343 B.n356 B.n56 256.663
R344 B.n356 B.n55 256.663
R345 B.n356 B.n54 256.663
R346 B.n356 B.n53 256.663
R347 B.n356 B.n52 256.663
R348 B.n356 B.n51 256.663
R349 B.n356 B.n50 256.663
R350 B.n356 B.n49 256.663
R351 B.n356 B.n48 256.663
R352 B.n356 B.n47 256.663
R353 B.n357 B.n356 256.663
R354 B.n253 B.n252 256.663
R355 B.n252 B.n172 256.663
R356 B.n252 B.n173 256.663
R357 B.n252 B.n174 256.663
R358 B.n252 B.n175 256.663
R359 B.n252 B.n176 256.663
R360 B.n252 B.n177 256.663
R361 B.n252 B.n178 256.663
R362 B.n252 B.n179 256.663
R363 B.n252 B.n180 256.663
R364 B.n252 B.n181 256.663
R365 B.n252 B.n182 256.663
R366 B.n252 B.n183 256.663
R367 B.n252 B.n184 256.663
R368 B.n252 B.n185 256.663
R369 B.n191 B.t13 226.369
R370 B.n188 B.t9 226.369
R371 B.n65 B.t2 226.369
R372 B.n63 B.t6 226.369
R373 B.n252 B.n168 186.868
R374 B.n356 B.n43 186.868
R375 B.n191 B.t15 166.655
R376 B.n63 B.t7 166.655
R377 B.n188 B.t12 166.655
R378 B.n65 B.t4 166.655
R379 B.n258 B.n169 163.367
R380 B.n258 B.n163 163.367
R381 B.n266 B.n163 163.367
R382 B.n266 B.n161 163.367
R383 B.n270 B.n161 163.367
R384 B.n270 B.n155 163.367
R385 B.n278 B.n155 163.367
R386 B.n278 B.n153 163.367
R387 B.n282 B.n153 163.367
R388 B.n282 B.n147 163.367
R389 B.n290 B.n147 163.367
R390 B.n290 B.n145 163.367
R391 B.n294 B.n145 163.367
R392 B.n294 B.n139 163.367
R393 B.n302 B.n139 163.367
R394 B.n302 B.n137 163.367
R395 B.n306 B.n137 163.367
R396 B.n306 B.n131 163.367
R397 B.n315 B.n131 163.367
R398 B.n315 B.n129 163.367
R399 B.n319 B.n129 163.367
R400 B.n319 B.n2 163.367
R401 B.n406 B.n2 163.367
R402 B.n406 B.n3 163.367
R403 B.n402 B.n3 163.367
R404 B.n402 B.n9 163.367
R405 B.n398 B.n9 163.367
R406 B.n398 B.n11 163.367
R407 B.n394 B.n11 163.367
R408 B.n394 B.n16 163.367
R409 B.n390 B.n16 163.367
R410 B.n390 B.n18 163.367
R411 B.n386 B.n18 163.367
R412 B.n386 B.n23 163.367
R413 B.n382 B.n23 163.367
R414 B.n382 B.n25 163.367
R415 B.n378 B.n25 163.367
R416 B.n378 B.n30 163.367
R417 B.n374 B.n30 163.367
R418 B.n374 B.n32 163.367
R419 B.n370 B.n32 163.367
R420 B.n370 B.n37 163.367
R421 B.n366 B.n37 163.367
R422 B.n366 B.n39 163.367
R423 B.n362 B.n39 163.367
R424 B.n362 B.n44 163.367
R425 B.n251 B.n171 163.367
R426 B.n251 B.n187 163.367
R427 B.n247 B.n246 163.367
R428 B.n243 B.n242 163.367
R429 B.n239 B.n238 163.367
R430 B.n235 B.n234 163.367
R431 B.n231 B.n230 163.367
R432 B.n227 B.n226 163.367
R433 B.n223 B.n222 163.367
R434 B.n219 B.n218 163.367
R435 B.n215 B.n214 163.367
R436 B.n211 B.n210 163.367
R437 B.n207 B.n206 163.367
R438 B.n203 B.n202 163.367
R439 B.n199 B.n198 163.367
R440 B.n195 B.n186 163.367
R441 B.n260 B.n167 163.367
R442 B.n260 B.n165 163.367
R443 B.n264 B.n165 163.367
R444 B.n264 B.n159 163.367
R445 B.n272 B.n159 163.367
R446 B.n272 B.n157 163.367
R447 B.n276 B.n157 163.367
R448 B.n276 B.n151 163.367
R449 B.n284 B.n151 163.367
R450 B.n284 B.n149 163.367
R451 B.n288 B.n149 163.367
R452 B.n288 B.n143 163.367
R453 B.n296 B.n143 163.367
R454 B.n296 B.n141 163.367
R455 B.n300 B.n141 163.367
R456 B.n300 B.n135 163.367
R457 B.n308 B.n135 163.367
R458 B.n308 B.n133 163.367
R459 B.n313 B.n133 163.367
R460 B.n313 B.n127 163.367
R461 B.n321 B.n127 163.367
R462 B.n322 B.n321 163.367
R463 B.n322 B.n5 163.367
R464 B.n6 B.n5 163.367
R465 B.n7 B.n6 163.367
R466 B.n327 B.n7 163.367
R467 B.n327 B.n12 163.367
R468 B.n13 B.n12 163.367
R469 B.n14 B.n13 163.367
R470 B.n332 B.n14 163.367
R471 B.n332 B.n19 163.367
R472 B.n20 B.n19 163.367
R473 B.n21 B.n20 163.367
R474 B.n337 B.n21 163.367
R475 B.n337 B.n26 163.367
R476 B.n27 B.n26 163.367
R477 B.n28 B.n27 163.367
R478 B.n342 B.n28 163.367
R479 B.n342 B.n33 163.367
R480 B.n34 B.n33 163.367
R481 B.n35 B.n34 163.367
R482 B.n347 B.n35 163.367
R483 B.n347 B.n40 163.367
R484 B.n41 B.n40 163.367
R485 B.n42 B.n41 163.367
R486 B.n62 B.n42 163.367
R487 B.n67 B.n46 163.367
R488 B.n71 B.n70 163.367
R489 B.n75 B.n74 163.367
R490 B.n79 B.n78 163.367
R491 B.n83 B.n82 163.367
R492 B.n88 B.n87 163.367
R493 B.n92 B.n91 163.367
R494 B.n96 B.n95 163.367
R495 B.n100 B.n99 163.367
R496 B.n104 B.n103 163.367
R497 B.n109 B.n108 163.367
R498 B.n113 B.n112 163.367
R499 B.n117 B.n116 163.367
R500 B.n121 B.n120 163.367
R501 B.n123 B.n61 163.367
R502 B.n192 B.t14 117.782
R503 B.n64 B.t8 117.782
R504 B.n189 B.t11 117.781
R505 B.n66 B.t5 117.781
R506 B.n259 B.n168 106.781
R507 B.n259 B.n164 106.781
R508 B.n265 B.n164 106.781
R509 B.n265 B.n160 106.781
R510 B.n271 B.n160 106.781
R511 B.n271 B.n156 106.781
R512 B.n277 B.n156 106.781
R513 B.n283 B.n152 106.781
R514 B.n283 B.n148 106.781
R515 B.n289 B.n148 106.781
R516 B.n289 B.n144 106.781
R517 B.n295 B.n144 106.781
R518 B.n295 B.n140 106.781
R519 B.n301 B.n140 106.781
R520 B.n301 B.n136 106.781
R521 B.n307 B.n136 106.781
R522 B.n314 B.n132 106.781
R523 B.n314 B.n128 106.781
R524 B.n320 B.n128 106.781
R525 B.n320 B.n4 106.781
R526 B.n405 B.n4 106.781
R527 B.n405 B.n404 106.781
R528 B.n404 B.n403 106.781
R529 B.n403 B.n8 106.781
R530 B.n397 B.n8 106.781
R531 B.n397 B.n396 106.781
R532 B.n395 B.n15 106.781
R533 B.n389 B.n15 106.781
R534 B.n389 B.n388 106.781
R535 B.n388 B.n387 106.781
R536 B.n387 B.n22 106.781
R537 B.n381 B.n22 106.781
R538 B.n381 B.n380 106.781
R539 B.n380 B.n379 106.781
R540 B.n379 B.n29 106.781
R541 B.n373 B.n372 106.781
R542 B.n372 B.n371 106.781
R543 B.n371 B.n36 106.781
R544 B.n365 B.n36 106.781
R545 B.n365 B.n364 106.781
R546 B.n364 B.n363 106.781
R547 B.n363 B.n43 106.781
R548 B.t10 B.n152 98.9298
R549 B.t3 B.n29 98.9298
R550 B.n307 B.t0 73.8049
R551 B.t1 B.n395 73.8049
R552 B.n254 B.n253 71.676
R553 B.n187 B.n172 71.676
R554 B.n246 B.n173 71.676
R555 B.n242 B.n174 71.676
R556 B.n238 B.n175 71.676
R557 B.n234 B.n176 71.676
R558 B.n230 B.n177 71.676
R559 B.n226 B.n178 71.676
R560 B.n222 B.n179 71.676
R561 B.n218 B.n180 71.676
R562 B.n214 B.n181 71.676
R563 B.n210 B.n182 71.676
R564 B.n206 B.n183 71.676
R565 B.n202 B.n184 71.676
R566 B.n198 B.n185 71.676
R567 B.n358 B.n357 71.676
R568 B.n67 B.n47 71.676
R569 B.n71 B.n48 71.676
R570 B.n75 B.n49 71.676
R571 B.n79 B.n50 71.676
R572 B.n83 B.n51 71.676
R573 B.n88 B.n52 71.676
R574 B.n92 B.n53 71.676
R575 B.n96 B.n54 71.676
R576 B.n100 B.n55 71.676
R577 B.n104 B.n56 71.676
R578 B.n109 B.n57 71.676
R579 B.n113 B.n58 71.676
R580 B.n117 B.n59 71.676
R581 B.n121 B.n60 71.676
R582 B.n355 B.n61 71.676
R583 B.n355 B.n354 71.676
R584 B.n123 B.n60 71.676
R585 B.n120 B.n59 71.676
R586 B.n116 B.n58 71.676
R587 B.n112 B.n57 71.676
R588 B.n108 B.n56 71.676
R589 B.n103 B.n55 71.676
R590 B.n99 B.n54 71.676
R591 B.n95 B.n53 71.676
R592 B.n91 B.n52 71.676
R593 B.n87 B.n51 71.676
R594 B.n82 B.n50 71.676
R595 B.n78 B.n49 71.676
R596 B.n74 B.n48 71.676
R597 B.n70 B.n47 71.676
R598 B.n357 B.n46 71.676
R599 B.n253 B.n171 71.676
R600 B.n247 B.n172 71.676
R601 B.n243 B.n173 71.676
R602 B.n239 B.n174 71.676
R603 B.n235 B.n175 71.676
R604 B.n231 B.n176 71.676
R605 B.n227 B.n177 71.676
R606 B.n223 B.n178 71.676
R607 B.n219 B.n179 71.676
R608 B.n215 B.n180 71.676
R609 B.n211 B.n181 71.676
R610 B.n207 B.n182 71.676
R611 B.n203 B.n183 71.676
R612 B.n199 B.n184 71.676
R613 B.n195 B.n185 71.676
R614 B.n193 B.n192 59.5399
R615 B.n190 B.n189 59.5399
R616 B.n85 B.n66 59.5399
R617 B.n106 B.n64 59.5399
R618 B.n192 B.n191 48.8732
R619 B.n189 B.n188 48.8732
R620 B.n66 B.n65 48.8732
R621 B.n64 B.n63 48.8732
R622 B.n360 B.n359 33.8737
R623 B.n353 B.n352 33.8737
R624 B.n194 B.n166 33.8737
R625 B.n256 B.n255 33.8737
R626 B.t0 B.n132 32.9769
R627 B.n396 B.t1 32.9769
R628 B B.n407 18.0485
R629 B.n359 B.n45 10.6151
R630 B.n68 B.n45 10.6151
R631 B.n69 B.n68 10.6151
R632 B.n72 B.n69 10.6151
R633 B.n73 B.n72 10.6151
R634 B.n76 B.n73 10.6151
R635 B.n77 B.n76 10.6151
R636 B.n80 B.n77 10.6151
R637 B.n81 B.n80 10.6151
R638 B.n84 B.n81 10.6151
R639 B.n89 B.n86 10.6151
R640 B.n90 B.n89 10.6151
R641 B.n93 B.n90 10.6151
R642 B.n94 B.n93 10.6151
R643 B.n97 B.n94 10.6151
R644 B.n98 B.n97 10.6151
R645 B.n101 B.n98 10.6151
R646 B.n102 B.n101 10.6151
R647 B.n105 B.n102 10.6151
R648 B.n110 B.n107 10.6151
R649 B.n111 B.n110 10.6151
R650 B.n114 B.n111 10.6151
R651 B.n115 B.n114 10.6151
R652 B.n118 B.n115 10.6151
R653 B.n119 B.n118 10.6151
R654 B.n122 B.n119 10.6151
R655 B.n124 B.n122 10.6151
R656 B.n125 B.n124 10.6151
R657 B.n353 B.n125 10.6151
R658 B.n261 B.n166 10.6151
R659 B.n262 B.n261 10.6151
R660 B.n263 B.n262 10.6151
R661 B.n263 B.n158 10.6151
R662 B.n273 B.n158 10.6151
R663 B.n274 B.n273 10.6151
R664 B.n275 B.n274 10.6151
R665 B.n275 B.n150 10.6151
R666 B.n285 B.n150 10.6151
R667 B.n286 B.n285 10.6151
R668 B.n287 B.n286 10.6151
R669 B.n287 B.n142 10.6151
R670 B.n297 B.n142 10.6151
R671 B.n298 B.n297 10.6151
R672 B.n299 B.n298 10.6151
R673 B.n299 B.n134 10.6151
R674 B.n309 B.n134 10.6151
R675 B.n310 B.n309 10.6151
R676 B.n312 B.n310 10.6151
R677 B.n312 B.n311 10.6151
R678 B.n311 B.n126 10.6151
R679 B.n323 B.n126 10.6151
R680 B.n324 B.n323 10.6151
R681 B.n325 B.n324 10.6151
R682 B.n326 B.n325 10.6151
R683 B.n328 B.n326 10.6151
R684 B.n329 B.n328 10.6151
R685 B.n330 B.n329 10.6151
R686 B.n331 B.n330 10.6151
R687 B.n333 B.n331 10.6151
R688 B.n334 B.n333 10.6151
R689 B.n335 B.n334 10.6151
R690 B.n336 B.n335 10.6151
R691 B.n338 B.n336 10.6151
R692 B.n339 B.n338 10.6151
R693 B.n340 B.n339 10.6151
R694 B.n341 B.n340 10.6151
R695 B.n343 B.n341 10.6151
R696 B.n344 B.n343 10.6151
R697 B.n345 B.n344 10.6151
R698 B.n346 B.n345 10.6151
R699 B.n348 B.n346 10.6151
R700 B.n349 B.n348 10.6151
R701 B.n350 B.n349 10.6151
R702 B.n351 B.n350 10.6151
R703 B.n352 B.n351 10.6151
R704 B.n255 B.n170 10.6151
R705 B.n250 B.n170 10.6151
R706 B.n250 B.n249 10.6151
R707 B.n249 B.n248 10.6151
R708 B.n248 B.n245 10.6151
R709 B.n245 B.n244 10.6151
R710 B.n244 B.n241 10.6151
R711 B.n241 B.n240 10.6151
R712 B.n240 B.n237 10.6151
R713 B.n237 B.n236 10.6151
R714 B.n233 B.n232 10.6151
R715 B.n232 B.n229 10.6151
R716 B.n229 B.n228 10.6151
R717 B.n228 B.n225 10.6151
R718 B.n225 B.n224 10.6151
R719 B.n224 B.n221 10.6151
R720 B.n221 B.n220 10.6151
R721 B.n220 B.n217 10.6151
R722 B.n217 B.n216 10.6151
R723 B.n213 B.n212 10.6151
R724 B.n212 B.n209 10.6151
R725 B.n209 B.n208 10.6151
R726 B.n208 B.n205 10.6151
R727 B.n205 B.n204 10.6151
R728 B.n204 B.n201 10.6151
R729 B.n201 B.n200 10.6151
R730 B.n200 B.n197 10.6151
R731 B.n197 B.n196 10.6151
R732 B.n196 B.n194 10.6151
R733 B.n257 B.n256 10.6151
R734 B.n257 B.n162 10.6151
R735 B.n267 B.n162 10.6151
R736 B.n268 B.n267 10.6151
R737 B.n269 B.n268 10.6151
R738 B.n269 B.n154 10.6151
R739 B.n279 B.n154 10.6151
R740 B.n280 B.n279 10.6151
R741 B.n281 B.n280 10.6151
R742 B.n281 B.n146 10.6151
R743 B.n291 B.n146 10.6151
R744 B.n292 B.n291 10.6151
R745 B.n293 B.n292 10.6151
R746 B.n293 B.n138 10.6151
R747 B.n303 B.n138 10.6151
R748 B.n304 B.n303 10.6151
R749 B.n305 B.n304 10.6151
R750 B.n305 B.n130 10.6151
R751 B.n316 B.n130 10.6151
R752 B.n317 B.n316 10.6151
R753 B.n318 B.n317 10.6151
R754 B.n318 B.n0 10.6151
R755 B.n401 B.n1 10.6151
R756 B.n401 B.n400 10.6151
R757 B.n400 B.n399 10.6151
R758 B.n399 B.n10 10.6151
R759 B.n393 B.n10 10.6151
R760 B.n393 B.n392 10.6151
R761 B.n392 B.n391 10.6151
R762 B.n391 B.n17 10.6151
R763 B.n385 B.n17 10.6151
R764 B.n385 B.n384 10.6151
R765 B.n384 B.n383 10.6151
R766 B.n383 B.n24 10.6151
R767 B.n377 B.n24 10.6151
R768 B.n377 B.n376 10.6151
R769 B.n376 B.n375 10.6151
R770 B.n375 B.n31 10.6151
R771 B.n369 B.n31 10.6151
R772 B.n369 B.n368 10.6151
R773 B.n368 B.n367 10.6151
R774 B.n367 B.n38 10.6151
R775 B.n361 B.n38 10.6151
R776 B.n361 B.n360 10.6151
R777 B.n85 B.n84 9.36635
R778 B.n107 B.n106 9.36635
R779 B.n236 B.n190 9.36635
R780 B.n213 B.n193 9.36635
R781 B.n277 B.t10 7.85203
R782 B.n373 B.t3 7.85203
R783 B.n407 B.n0 2.81026
R784 B.n407 B.n1 2.81026
R785 B.n86 B.n85 1.24928
R786 B.n106 B.n105 1.24928
R787 B.n233 B.n190 1.24928
R788 B.n216 B.n193 1.24928
R789 VN VN.t1 104.094
R790 VN VN.t0 68.545
R791 VDD2.n9 VDD2.n7 289.615
R792 VDD2.n2 VDD2.n0 289.615
R793 VDD2.n10 VDD2.n9 185
R794 VDD2.n3 VDD2.n2 185
R795 VDD2.t0 VDD2.n8 164.876
R796 VDD2.t1 VDD2.n1 164.876
R797 VDD2.n14 VDD2.n6 79.3295
R798 VDD2.n9 VDD2.t0 52.3082
R799 VDD2.n2 VDD2.t1 52.3082
R800 VDD2.n14 VDD2.n13 49.8338
R801 VDD2.n10 VDD2.n8 14.7318
R802 VDD2.n3 VDD2.n1 14.7318
R803 VDD2.n11 VDD2.n7 12.8005
R804 VDD2.n4 VDD2.n0 12.8005
R805 VDD2.n13 VDD2.n12 9.45567
R806 VDD2.n6 VDD2.n5 9.45567
R807 VDD2.n12 VDD2.n11 9.3005
R808 VDD2.n5 VDD2.n4 9.3005
R809 VDD2.n12 VDD2.n8 5.62509
R810 VDD2.n5 VDD2.n1 5.62509
R811 VDD2.n13 VDD2.n7 1.16414
R812 VDD2.n6 VDD2.n0 1.16414
R813 VDD2 VDD2.n14 0.601793
R814 VDD2.n11 VDD2.n10 0.388379
R815 VDD2.n4 VDD2.n3 0.388379
C0 VDD1 VN 0.154633f
C1 VDD2 VP 0.322469f
C2 VDD2 VTAIL 2.27101f
C3 VDD2 VN 0.606378f
C4 VDD1 VDD2 0.624297f
C5 VP VTAIL 0.877975f
C6 VP VN 3.37217f
C7 VDD1 VP 0.772582f
C8 VTAIL VN 0.863837f
C9 VDD1 VTAIL 2.22084f
C10 VDD2 B 2.409207f
C11 VDD1 B 3.87301f
C12 VTAIL B 2.722439f
C13 VN B 7.07783f
C14 VP B 4.9987f
C15 VDD2.n0 B 0.022786f
C16 VDD2.n1 B 0.053375f
C17 VDD2.t1 B 0.038574f
C18 VDD2.n2 B 0.039338f
C19 VDD2.n3 B 0.011808f
C20 VDD2.n4 B 0.009585f
C21 VDD2.n5 B 0.103492f
C22 VDD2.n6 B 0.271973f
C23 VDD2.n7 B 0.022786f
C24 VDD2.n8 B 0.053375f
C25 VDD2.t0 B 0.038574f
C26 VDD2.n9 B 0.039338f
C27 VDD2.n10 B 0.011808f
C28 VDD2.n11 B 0.009585f
C29 VDD2.n12 B 0.103492f
C30 VDD2.n13 B 0.037109f
C31 VDD2.n14 B 1.33551f
C32 VN.t0 B 0.497312f
C33 VN.t1 B 0.902683f
C34 VDD1.n0 B 0.021188f
C35 VDD1.n1 B 0.049633f
C36 VDD1.t0 B 0.03587f
C37 VDD1.n2 B 0.03658f
C38 VDD1.n3 B 0.01098f
C39 VDD1.n4 B 0.008913f
C40 VDD1.n5 B 0.096236f
C41 VDD1.n6 B 0.035279f
C42 VDD1.n7 B 0.021188f
C43 VDD1.n8 B 0.049633f
C44 VDD1.t1 B 0.03587f
C45 VDD1.n9 B 0.03658f
C46 VDD1.n10 B 0.01098f
C47 VDD1.n11 B 0.008913f
C48 VDD1.n12 B 0.096236f
C49 VDD1.n13 B 0.27645f
C50 VTAIL.n0 B 0.027729f
C51 VTAIL.n1 B 0.064955f
C52 VTAIL.t2 B 0.046943f
C53 VTAIL.n2 B 0.047873f
C54 VTAIL.n3 B 0.01437f
C55 VTAIL.n4 B 0.011665f
C56 VTAIL.n5 B 0.125946f
C57 VTAIL.n6 B 0.030183f
C58 VTAIL.n7 B 0.797394f
C59 VTAIL.n8 B 0.027729f
C60 VTAIL.n9 B 0.064955f
C61 VTAIL.t0 B 0.046943f
C62 VTAIL.n10 B 0.047873f
C63 VTAIL.n11 B 0.01437f
C64 VTAIL.n12 B 0.011665f
C65 VTAIL.n13 B 0.125946f
C66 VTAIL.n14 B 0.030183f
C67 VTAIL.n15 B 0.831312f
C68 VTAIL.n16 B 0.027729f
C69 VTAIL.n17 B 0.064955f
C70 VTAIL.t1 B 0.046943f
C71 VTAIL.n18 B 0.047873f
C72 VTAIL.n19 B 0.01437f
C73 VTAIL.n20 B 0.011665f
C74 VTAIL.n21 B 0.125946f
C75 VTAIL.n22 B 0.030183f
C76 VTAIL.n23 B 0.679359f
C77 VTAIL.n24 B 0.027729f
C78 VTAIL.n25 B 0.064955f
C79 VTAIL.t3 B 0.046943f
C80 VTAIL.n26 B 0.047873f
C81 VTAIL.n27 B 0.01437f
C82 VTAIL.n28 B 0.011665f
C83 VTAIL.n29 B 0.125946f
C84 VTAIL.n30 B 0.030183f
C85 VTAIL.n31 B 0.604437f
C86 VP.t1 B 0.909356f
C87 VP.t0 B 0.502776f
C88 VP.n0 B 1.92444f
.ends

