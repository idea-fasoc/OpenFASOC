* NGSPICE file created from diff_pair_sample_1082.ext - technology: sky130A

.subckt diff_pair_sample_1082 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8976 pd=5.77 as=0.8976 ps=5.77 w=5.44 l=3.27
X1 VDD1.t7 VP.t0 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.8976 pd=5.77 as=0.8976 ps=5.77 w=5.44 l=3.27
X2 VTAIL.t7 VP.t1 VDD1.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=2.1216 pd=11.66 as=0.8976 ps=5.77 w=5.44 l=3.27
X3 VTAIL.t2 VP.t2 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1216 pd=11.66 as=0.8976 ps=5.77 w=5.44 l=3.27
X4 VDD1.t4 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.8976 pd=5.77 as=2.1216 ps=11.66 w=5.44 l=3.27
X5 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=2.1216 pd=11.66 as=0 ps=0 w=5.44 l=3.27
X6 VTAIL.t1 VP.t4 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8976 pd=5.77 as=0.8976 ps=5.77 w=5.44 l=3.27
X7 VDD1.t2 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.8976 pd=5.77 as=2.1216 ps=11.66 w=5.44 l=3.27
X8 VDD2.t6 VN.t1 VTAIL.t14 B.t5 sky130_fd_pr__nfet_01v8 ad=0.8976 pd=5.77 as=0.8976 ps=5.77 w=5.44 l=3.27
X9 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=2.1216 pd=11.66 as=0 ps=0 w=5.44 l=3.27
X10 VDD2.t0 VN.t2 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=0.8976 pd=5.77 as=2.1216 ps=11.66 w=5.44 l=3.27
X11 VDD2.t7 VN.t3 VTAIL.t12 B.t3 sky130_fd_pr__nfet_01v8 ad=0.8976 pd=5.77 as=2.1216 ps=11.66 w=5.44 l=3.27
X12 VDD1.t1 VP.t6 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.8976 pd=5.77 as=0.8976 ps=5.77 w=5.44 l=3.27
X13 VTAIL.t11 VN.t4 VDD2.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=0.8976 pd=5.77 as=0.8976 ps=5.77 w=5.44 l=3.27
X14 VTAIL.t10 VN.t5 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1216 pd=11.66 as=0.8976 ps=5.77 w=5.44 l=3.27
X15 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=2.1216 pd=11.66 as=0 ps=0 w=5.44 l=3.27
X16 VTAIL.t6 VP.t7 VDD1.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=0.8976 pd=5.77 as=0.8976 ps=5.77 w=5.44 l=3.27
X17 VTAIL.t9 VN.t6 VDD2.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=2.1216 pd=11.66 as=0.8976 ps=5.77 w=5.44 l=3.27
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.1216 pd=11.66 as=0 ps=0 w=5.44 l=3.27
X19 VDD2.t5 VN.t7 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=0.8976 pd=5.77 as=0.8976 ps=5.77 w=5.44 l=3.27
R0 VN.n64 VN.n63 161.3
R1 VN.n62 VN.n34 161.3
R2 VN.n61 VN.n60 161.3
R3 VN.n59 VN.n35 161.3
R4 VN.n58 VN.n57 161.3
R5 VN.n56 VN.n36 161.3
R6 VN.n55 VN.n54 161.3
R7 VN.n53 VN.n52 161.3
R8 VN.n51 VN.n38 161.3
R9 VN.n50 VN.n49 161.3
R10 VN.n48 VN.n39 161.3
R11 VN.n47 VN.n46 161.3
R12 VN.n45 VN.n40 161.3
R13 VN.n44 VN.n43 161.3
R14 VN.n31 VN.n30 161.3
R15 VN.n29 VN.n1 161.3
R16 VN.n28 VN.n27 161.3
R17 VN.n26 VN.n2 161.3
R18 VN.n25 VN.n24 161.3
R19 VN.n23 VN.n3 161.3
R20 VN.n22 VN.n21 161.3
R21 VN.n20 VN.n19 161.3
R22 VN.n18 VN.n5 161.3
R23 VN.n17 VN.n16 161.3
R24 VN.n15 VN.n6 161.3
R25 VN.n14 VN.n13 161.3
R26 VN.n12 VN.n7 161.3
R27 VN.n11 VN.n10 161.3
R28 VN.n42 VN.t3 73.5144
R29 VN.n9 VN.t5 73.5144
R30 VN.n32 VN.n0 70.5721
R31 VN.n65 VN.n33 70.5721
R32 VN.n42 VN.n41 59.6504
R33 VN.n9 VN.n8 59.6504
R34 VN.n28 VN.n2 50.2647
R35 VN.n61 VN.n35 50.2647
R36 VN VN.n65 49.4072
R37 VN.n13 VN.n6 40.577
R38 VN.n17 VN.n6 40.577
R39 VN.n46 VN.n39 40.577
R40 VN.n50 VN.n39 40.577
R41 VN.n8 VN.t7 40.0935
R42 VN.n4 VN.t4 40.0935
R43 VN.n0 VN.t2 40.0935
R44 VN.n41 VN.t0 40.0935
R45 VN.n37 VN.t1 40.0935
R46 VN.n33 VN.t6 40.0935
R47 VN.n24 VN.n2 30.8893
R48 VN.n57 VN.n35 30.8893
R49 VN.n12 VN.n11 24.5923
R50 VN.n13 VN.n12 24.5923
R51 VN.n18 VN.n17 24.5923
R52 VN.n19 VN.n18 24.5923
R53 VN.n23 VN.n22 24.5923
R54 VN.n24 VN.n23 24.5923
R55 VN.n29 VN.n28 24.5923
R56 VN.n30 VN.n29 24.5923
R57 VN.n46 VN.n45 24.5923
R58 VN.n45 VN.n44 24.5923
R59 VN.n57 VN.n56 24.5923
R60 VN.n56 VN.n55 24.5923
R61 VN.n52 VN.n51 24.5923
R62 VN.n51 VN.n50 24.5923
R63 VN.n63 VN.n62 24.5923
R64 VN.n62 VN.n61 24.5923
R65 VN.n30 VN.n0 19.674
R66 VN.n63 VN.n33 19.674
R67 VN.n11 VN.n8 14.7556
R68 VN.n19 VN.n4 14.7556
R69 VN.n44 VN.n41 14.7556
R70 VN.n52 VN.n37 14.7556
R71 VN.n22 VN.n4 9.83723
R72 VN.n55 VN.n37 9.83723
R73 VN.n43 VN.n42 3.91115
R74 VN.n10 VN.n9 3.91115
R75 VN.n65 VN.n64 0.354861
R76 VN.n32 VN.n31 0.354861
R77 VN VN.n32 0.267071
R78 VN.n64 VN.n34 0.189894
R79 VN.n60 VN.n34 0.189894
R80 VN.n60 VN.n59 0.189894
R81 VN.n59 VN.n58 0.189894
R82 VN.n58 VN.n36 0.189894
R83 VN.n54 VN.n36 0.189894
R84 VN.n54 VN.n53 0.189894
R85 VN.n53 VN.n38 0.189894
R86 VN.n49 VN.n38 0.189894
R87 VN.n49 VN.n48 0.189894
R88 VN.n48 VN.n47 0.189894
R89 VN.n47 VN.n40 0.189894
R90 VN.n43 VN.n40 0.189894
R91 VN.n10 VN.n7 0.189894
R92 VN.n14 VN.n7 0.189894
R93 VN.n15 VN.n14 0.189894
R94 VN.n16 VN.n15 0.189894
R95 VN.n16 VN.n5 0.189894
R96 VN.n20 VN.n5 0.189894
R97 VN.n21 VN.n20 0.189894
R98 VN.n21 VN.n3 0.189894
R99 VN.n25 VN.n3 0.189894
R100 VN.n26 VN.n25 0.189894
R101 VN.n27 VN.n26 0.189894
R102 VN.n27 VN.n1 0.189894
R103 VN.n31 VN.n1 0.189894
R104 VDD2.n2 VDD2.n1 71.566
R105 VDD2.n2 VDD2.n0 71.566
R106 VDD2 VDD2.n5 71.5624
R107 VDD2.n4 VDD2.n3 70.0698
R108 VDD2.n4 VDD2.n2 42.3705
R109 VDD2.n5 VDD2.t1 3.64021
R110 VDD2.n5 VDD2.t7 3.64021
R111 VDD2.n3 VDD2.t2 3.64021
R112 VDD2.n3 VDD2.t6 3.64021
R113 VDD2.n1 VDD2.t3 3.64021
R114 VDD2.n1 VDD2.t0 3.64021
R115 VDD2.n0 VDD2.t4 3.64021
R116 VDD2.n0 VDD2.t5 3.64021
R117 VDD2 VDD2.n4 1.61041
R118 VTAIL.n11 VTAIL.t2 57.0307
R119 VTAIL.n10 VTAIL.t12 57.0307
R120 VTAIL.n7 VTAIL.t9 57.0307
R121 VTAIL.n14 VTAIL.t0 57.0298
R122 VTAIL.n15 VTAIL.t13 57.0297
R123 VTAIL.n2 VTAIL.t10 57.0297
R124 VTAIL.n3 VTAIL.t3 57.0297
R125 VTAIL.n6 VTAIL.t7 57.0297
R126 VTAIL.n13 VTAIL.n12 53.391
R127 VTAIL.n9 VTAIL.n8 53.391
R128 VTAIL.n1 VTAIL.n0 53.3909
R129 VTAIL.n5 VTAIL.n4 53.3909
R130 VTAIL.n15 VTAIL.n14 20.16
R131 VTAIL.n7 VTAIL.n6 20.16
R132 VTAIL.n0 VTAIL.t8 3.64021
R133 VTAIL.n0 VTAIL.t11 3.64021
R134 VTAIL.n4 VTAIL.t5 3.64021
R135 VTAIL.n4 VTAIL.t1 3.64021
R136 VTAIL.n12 VTAIL.t4 3.64021
R137 VTAIL.n12 VTAIL.t6 3.64021
R138 VTAIL.n8 VTAIL.t14 3.64021
R139 VTAIL.n8 VTAIL.t15 3.64021
R140 VTAIL.n9 VTAIL.n7 3.10395
R141 VTAIL.n10 VTAIL.n9 3.10395
R142 VTAIL.n13 VTAIL.n11 3.10395
R143 VTAIL.n14 VTAIL.n13 3.10395
R144 VTAIL.n6 VTAIL.n5 3.10395
R145 VTAIL.n5 VTAIL.n3 3.10395
R146 VTAIL.n2 VTAIL.n1 3.10395
R147 VTAIL VTAIL.n15 3.04576
R148 VTAIL.n11 VTAIL.n10 0.470328
R149 VTAIL.n3 VTAIL.n2 0.470328
R150 VTAIL VTAIL.n1 0.0586897
R151 B.n771 B.n770 585
R152 B.n249 B.n138 585
R153 B.n248 B.n247 585
R154 B.n246 B.n245 585
R155 B.n244 B.n243 585
R156 B.n242 B.n241 585
R157 B.n240 B.n239 585
R158 B.n238 B.n237 585
R159 B.n236 B.n235 585
R160 B.n234 B.n233 585
R161 B.n232 B.n231 585
R162 B.n230 B.n229 585
R163 B.n228 B.n227 585
R164 B.n226 B.n225 585
R165 B.n224 B.n223 585
R166 B.n222 B.n221 585
R167 B.n220 B.n219 585
R168 B.n218 B.n217 585
R169 B.n216 B.n215 585
R170 B.n214 B.n213 585
R171 B.n212 B.n211 585
R172 B.n210 B.n209 585
R173 B.n208 B.n207 585
R174 B.n206 B.n205 585
R175 B.n204 B.n203 585
R176 B.n202 B.n201 585
R177 B.n200 B.n199 585
R178 B.n198 B.n197 585
R179 B.n196 B.n195 585
R180 B.n194 B.n193 585
R181 B.n192 B.n191 585
R182 B.n190 B.n189 585
R183 B.n188 B.n187 585
R184 B.n186 B.n185 585
R185 B.n184 B.n183 585
R186 B.n182 B.n181 585
R187 B.n180 B.n179 585
R188 B.n178 B.n177 585
R189 B.n176 B.n175 585
R190 B.n174 B.n173 585
R191 B.n172 B.n171 585
R192 B.n170 B.n169 585
R193 B.n168 B.n167 585
R194 B.n166 B.n165 585
R195 B.n164 B.n163 585
R196 B.n162 B.n161 585
R197 B.n160 B.n159 585
R198 B.n158 B.n157 585
R199 B.n156 B.n155 585
R200 B.n154 B.n153 585
R201 B.n152 B.n151 585
R202 B.n150 B.n149 585
R203 B.n148 B.n147 585
R204 B.n146 B.n145 585
R205 B.n769 B.n111 585
R206 B.n774 B.n111 585
R207 B.n768 B.n110 585
R208 B.n775 B.n110 585
R209 B.n767 B.n766 585
R210 B.n766 B.n106 585
R211 B.n765 B.n105 585
R212 B.n781 B.n105 585
R213 B.n764 B.n104 585
R214 B.n782 B.n104 585
R215 B.n763 B.n103 585
R216 B.n783 B.n103 585
R217 B.n762 B.n761 585
R218 B.n761 B.n99 585
R219 B.n760 B.n98 585
R220 B.n789 B.n98 585
R221 B.n759 B.n97 585
R222 B.n790 B.n97 585
R223 B.n758 B.n96 585
R224 B.n791 B.n96 585
R225 B.n757 B.n756 585
R226 B.n756 B.n92 585
R227 B.n755 B.n91 585
R228 B.n797 B.n91 585
R229 B.n754 B.n90 585
R230 B.n798 B.n90 585
R231 B.n753 B.n89 585
R232 B.n799 B.n89 585
R233 B.n752 B.n751 585
R234 B.n751 B.n85 585
R235 B.n750 B.n84 585
R236 B.n805 B.n84 585
R237 B.n749 B.n83 585
R238 B.n806 B.n83 585
R239 B.n748 B.n82 585
R240 B.n807 B.n82 585
R241 B.n747 B.n746 585
R242 B.n746 B.n78 585
R243 B.n745 B.n77 585
R244 B.n813 B.n77 585
R245 B.n744 B.n76 585
R246 B.n814 B.n76 585
R247 B.n743 B.n75 585
R248 B.n815 B.n75 585
R249 B.n742 B.n741 585
R250 B.n741 B.n74 585
R251 B.n740 B.n70 585
R252 B.n821 B.n70 585
R253 B.n739 B.n69 585
R254 B.n822 B.n69 585
R255 B.n738 B.n68 585
R256 B.n823 B.n68 585
R257 B.n737 B.n736 585
R258 B.n736 B.n64 585
R259 B.n735 B.n63 585
R260 B.n829 B.n63 585
R261 B.n734 B.n62 585
R262 B.n830 B.n62 585
R263 B.n733 B.n61 585
R264 B.n831 B.n61 585
R265 B.n732 B.n731 585
R266 B.n731 B.n57 585
R267 B.n730 B.n56 585
R268 B.n837 B.n56 585
R269 B.n729 B.n55 585
R270 B.n838 B.n55 585
R271 B.n728 B.n54 585
R272 B.n839 B.n54 585
R273 B.n727 B.n726 585
R274 B.n726 B.n50 585
R275 B.n725 B.n49 585
R276 B.n845 B.n49 585
R277 B.n724 B.n48 585
R278 B.n846 B.n48 585
R279 B.n723 B.n47 585
R280 B.n847 B.n47 585
R281 B.n722 B.n721 585
R282 B.n721 B.n43 585
R283 B.n720 B.n42 585
R284 B.n853 B.n42 585
R285 B.n719 B.n41 585
R286 B.n854 B.n41 585
R287 B.n718 B.n40 585
R288 B.n855 B.n40 585
R289 B.n717 B.n716 585
R290 B.n716 B.n36 585
R291 B.n715 B.n35 585
R292 B.n861 B.n35 585
R293 B.n714 B.n34 585
R294 B.n862 B.n34 585
R295 B.n713 B.n33 585
R296 B.n863 B.n33 585
R297 B.n712 B.n711 585
R298 B.n711 B.n29 585
R299 B.n710 B.n28 585
R300 B.n869 B.n28 585
R301 B.n709 B.n27 585
R302 B.n870 B.n27 585
R303 B.n708 B.n26 585
R304 B.n871 B.n26 585
R305 B.n707 B.n706 585
R306 B.n706 B.n22 585
R307 B.n705 B.n21 585
R308 B.n877 B.n21 585
R309 B.n704 B.n20 585
R310 B.n878 B.n20 585
R311 B.n703 B.n19 585
R312 B.n879 B.n19 585
R313 B.n702 B.n701 585
R314 B.n701 B.n18 585
R315 B.n700 B.n14 585
R316 B.n885 B.n14 585
R317 B.n699 B.n13 585
R318 B.n886 B.n13 585
R319 B.n698 B.n12 585
R320 B.n887 B.n12 585
R321 B.n697 B.n696 585
R322 B.n696 B.n8 585
R323 B.n695 B.n7 585
R324 B.n893 B.n7 585
R325 B.n694 B.n6 585
R326 B.n894 B.n6 585
R327 B.n693 B.n5 585
R328 B.n895 B.n5 585
R329 B.n692 B.n691 585
R330 B.n691 B.n4 585
R331 B.n690 B.n250 585
R332 B.n690 B.n689 585
R333 B.n680 B.n251 585
R334 B.n252 B.n251 585
R335 B.n682 B.n681 585
R336 B.n683 B.n682 585
R337 B.n679 B.n257 585
R338 B.n257 B.n256 585
R339 B.n678 B.n677 585
R340 B.n677 B.n676 585
R341 B.n259 B.n258 585
R342 B.n669 B.n259 585
R343 B.n668 B.n667 585
R344 B.n670 B.n668 585
R345 B.n666 B.n264 585
R346 B.n264 B.n263 585
R347 B.n665 B.n664 585
R348 B.n664 B.n663 585
R349 B.n266 B.n265 585
R350 B.n267 B.n266 585
R351 B.n656 B.n655 585
R352 B.n657 B.n656 585
R353 B.n654 B.n272 585
R354 B.n272 B.n271 585
R355 B.n653 B.n652 585
R356 B.n652 B.n651 585
R357 B.n274 B.n273 585
R358 B.n275 B.n274 585
R359 B.n644 B.n643 585
R360 B.n645 B.n644 585
R361 B.n642 B.n280 585
R362 B.n280 B.n279 585
R363 B.n641 B.n640 585
R364 B.n640 B.n639 585
R365 B.n282 B.n281 585
R366 B.n283 B.n282 585
R367 B.n632 B.n631 585
R368 B.n633 B.n632 585
R369 B.n630 B.n288 585
R370 B.n288 B.n287 585
R371 B.n629 B.n628 585
R372 B.n628 B.n627 585
R373 B.n290 B.n289 585
R374 B.n291 B.n290 585
R375 B.n620 B.n619 585
R376 B.n621 B.n620 585
R377 B.n618 B.n296 585
R378 B.n296 B.n295 585
R379 B.n617 B.n616 585
R380 B.n616 B.n615 585
R381 B.n298 B.n297 585
R382 B.n299 B.n298 585
R383 B.n608 B.n607 585
R384 B.n609 B.n608 585
R385 B.n606 B.n303 585
R386 B.n307 B.n303 585
R387 B.n605 B.n604 585
R388 B.n604 B.n603 585
R389 B.n305 B.n304 585
R390 B.n306 B.n305 585
R391 B.n596 B.n595 585
R392 B.n597 B.n596 585
R393 B.n594 B.n312 585
R394 B.n312 B.n311 585
R395 B.n593 B.n592 585
R396 B.n592 B.n591 585
R397 B.n314 B.n313 585
R398 B.n315 B.n314 585
R399 B.n584 B.n583 585
R400 B.n585 B.n584 585
R401 B.n582 B.n320 585
R402 B.n320 B.n319 585
R403 B.n581 B.n580 585
R404 B.n580 B.n579 585
R405 B.n322 B.n321 585
R406 B.n572 B.n322 585
R407 B.n571 B.n570 585
R408 B.n573 B.n571 585
R409 B.n569 B.n327 585
R410 B.n327 B.n326 585
R411 B.n568 B.n567 585
R412 B.n567 B.n566 585
R413 B.n329 B.n328 585
R414 B.n330 B.n329 585
R415 B.n559 B.n558 585
R416 B.n560 B.n559 585
R417 B.n557 B.n335 585
R418 B.n335 B.n334 585
R419 B.n556 B.n555 585
R420 B.n555 B.n554 585
R421 B.n337 B.n336 585
R422 B.n338 B.n337 585
R423 B.n547 B.n546 585
R424 B.n548 B.n547 585
R425 B.n545 B.n343 585
R426 B.n343 B.n342 585
R427 B.n544 B.n543 585
R428 B.n543 B.n542 585
R429 B.n345 B.n344 585
R430 B.n346 B.n345 585
R431 B.n535 B.n534 585
R432 B.n536 B.n535 585
R433 B.n533 B.n350 585
R434 B.n354 B.n350 585
R435 B.n532 B.n531 585
R436 B.n531 B.n530 585
R437 B.n352 B.n351 585
R438 B.n353 B.n352 585
R439 B.n523 B.n522 585
R440 B.n524 B.n523 585
R441 B.n521 B.n359 585
R442 B.n359 B.n358 585
R443 B.n520 B.n519 585
R444 B.n519 B.n518 585
R445 B.n361 B.n360 585
R446 B.n362 B.n361 585
R447 B.n511 B.n510 585
R448 B.n512 B.n511 585
R449 B.n509 B.n367 585
R450 B.n367 B.n366 585
R451 B.n504 B.n503 585
R452 B.n502 B.n396 585
R453 B.n501 B.n395 585
R454 B.n506 B.n395 585
R455 B.n500 B.n499 585
R456 B.n498 B.n497 585
R457 B.n496 B.n495 585
R458 B.n494 B.n493 585
R459 B.n492 B.n491 585
R460 B.n490 B.n489 585
R461 B.n488 B.n487 585
R462 B.n486 B.n485 585
R463 B.n484 B.n483 585
R464 B.n482 B.n481 585
R465 B.n480 B.n479 585
R466 B.n478 B.n477 585
R467 B.n476 B.n475 585
R468 B.n474 B.n473 585
R469 B.n472 B.n471 585
R470 B.n470 B.n469 585
R471 B.n468 B.n467 585
R472 B.n466 B.n465 585
R473 B.n464 B.n463 585
R474 B.n461 B.n460 585
R475 B.n459 B.n458 585
R476 B.n457 B.n456 585
R477 B.n455 B.n454 585
R478 B.n453 B.n452 585
R479 B.n451 B.n450 585
R480 B.n449 B.n448 585
R481 B.n447 B.n446 585
R482 B.n445 B.n444 585
R483 B.n443 B.n442 585
R484 B.n440 B.n439 585
R485 B.n438 B.n437 585
R486 B.n436 B.n435 585
R487 B.n434 B.n433 585
R488 B.n432 B.n431 585
R489 B.n430 B.n429 585
R490 B.n428 B.n427 585
R491 B.n426 B.n425 585
R492 B.n424 B.n423 585
R493 B.n422 B.n421 585
R494 B.n420 B.n419 585
R495 B.n418 B.n417 585
R496 B.n416 B.n415 585
R497 B.n414 B.n413 585
R498 B.n412 B.n411 585
R499 B.n410 B.n409 585
R500 B.n408 B.n407 585
R501 B.n406 B.n405 585
R502 B.n404 B.n403 585
R503 B.n402 B.n401 585
R504 B.n369 B.n368 585
R505 B.n508 B.n507 585
R506 B.n507 B.n506 585
R507 B.n365 B.n364 585
R508 B.n366 B.n365 585
R509 B.n514 B.n513 585
R510 B.n513 B.n512 585
R511 B.n515 B.n363 585
R512 B.n363 B.n362 585
R513 B.n517 B.n516 585
R514 B.n518 B.n517 585
R515 B.n357 B.n356 585
R516 B.n358 B.n357 585
R517 B.n526 B.n525 585
R518 B.n525 B.n524 585
R519 B.n527 B.n355 585
R520 B.n355 B.n353 585
R521 B.n529 B.n528 585
R522 B.n530 B.n529 585
R523 B.n349 B.n348 585
R524 B.n354 B.n349 585
R525 B.n538 B.n537 585
R526 B.n537 B.n536 585
R527 B.n539 B.n347 585
R528 B.n347 B.n346 585
R529 B.n541 B.n540 585
R530 B.n542 B.n541 585
R531 B.n341 B.n340 585
R532 B.n342 B.n341 585
R533 B.n550 B.n549 585
R534 B.n549 B.n548 585
R535 B.n551 B.n339 585
R536 B.n339 B.n338 585
R537 B.n553 B.n552 585
R538 B.n554 B.n553 585
R539 B.n333 B.n332 585
R540 B.n334 B.n333 585
R541 B.n562 B.n561 585
R542 B.n561 B.n560 585
R543 B.n563 B.n331 585
R544 B.n331 B.n330 585
R545 B.n565 B.n564 585
R546 B.n566 B.n565 585
R547 B.n325 B.n324 585
R548 B.n326 B.n325 585
R549 B.n575 B.n574 585
R550 B.n574 B.n573 585
R551 B.n576 B.n323 585
R552 B.n572 B.n323 585
R553 B.n578 B.n577 585
R554 B.n579 B.n578 585
R555 B.n318 B.n317 585
R556 B.n319 B.n318 585
R557 B.n587 B.n586 585
R558 B.n586 B.n585 585
R559 B.n588 B.n316 585
R560 B.n316 B.n315 585
R561 B.n590 B.n589 585
R562 B.n591 B.n590 585
R563 B.n310 B.n309 585
R564 B.n311 B.n310 585
R565 B.n599 B.n598 585
R566 B.n598 B.n597 585
R567 B.n600 B.n308 585
R568 B.n308 B.n306 585
R569 B.n602 B.n601 585
R570 B.n603 B.n602 585
R571 B.n302 B.n301 585
R572 B.n307 B.n302 585
R573 B.n611 B.n610 585
R574 B.n610 B.n609 585
R575 B.n612 B.n300 585
R576 B.n300 B.n299 585
R577 B.n614 B.n613 585
R578 B.n615 B.n614 585
R579 B.n294 B.n293 585
R580 B.n295 B.n294 585
R581 B.n623 B.n622 585
R582 B.n622 B.n621 585
R583 B.n624 B.n292 585
R584 B.n292 B.n291 585
R585 B.n626 B.n625 585
R586 B.n627 B.n626 585
R587 B.n286 B.n285 585
R588 B.n287 B.n286 585
R589 B.n635 B.n634 585
R590 B.n634 B.n633 585
R591 B.n636 B.n284 585
R592 B.n284 B.n283 585
R593 B.n638 B.n637 585
R594 B.n639 B.n638 585
R595 B.n278 B.n277 585
R596 B.n279 B.n278 585
R597 B.n647 B.n646 585
R598 B.n646 B.n645 585
R599 B.n648 B.n276 585
R600 B.n276 B.n275 585
R601 B.n650 B.n649 585
R602 B.n651 B.n650 585
R603 B.n270 B.n269 585
R604 B.n271 B.n270 585
R605 B.n659 B.n658 585
R606 B.n658 B.n657 585
R607 B.n660 B.n268 585
R608 B.n268 B.n267 585
R609 B.n662 B.n661 585
R610 B.n663 B.n662 585
R611 B.n262 B.n261 585
R612 B.n263 B.n262 585
R613 B.n672 B.n671 585
R614 B.n671 B.n670 585
R615 B.n673 B.n260 585
R616 B.n669 B.n260 585
R617 B.n675 B.n674 585
R618 B.n676 B.n675 585
R619 B.n255 B.n254 585
R620 B.n256 B.n255 585
R621 B.n685 B.n684 585
R622 B.n684 B.n683 585
R623 B.n686 B.n253 585
R624 B.n253 B.n252 585
R625 B.n688 B.n687 585
R626 B.n689 B.n688 585
R627 B.n2 B.n0 585
R628 B.n4 B.n2 585
R629 B.n3 B.n1 585
R630 B.n894 B.n3 585
R631 B.n892 B.n891 585
R632 B.n893 B.n892 585
R633 B.n890 B.n9 585
R634 B.n9 B.n8 585
R635 B.n889 B.n888 585
R636 B.n888 B.n887 585
R637 B.n11 B.n10 585
R638 B.n886 B.n11 585
R639 B.n884 B.n883 585
R640 B.n885 B.n884 585
R641 B.n882 B.n15 585
R642 B.n18 B.n15 585
R643 B.n881 B.n880 585
R644 B.n880 B.n879 585
R645 B.n17 B.n16 585
R646 B.n878 B.n17 585
R647 B.n876 B.n875 585
R648 B.n877 B.n876 585
R649 B.n874 B.n23 585
R650 B.n23 B.n22 585
R651 B.n873 B.n872 585
R652 B.n872 B.n871 585
R653 B.n25 B.n24 585
R654 B.n870 B.n25 585
R655 B.n868 B.n867 585
R656 B.n869 B.n868 585
R657 B.n866 B.n30 585
R658 B.n30 B.n29 585
R659 B.n865 B.n864 585
R660 B.n864 B.n863 585
R661 B.n32 B.n31 585
R662 B.n862 B.n32 585
R663 B.n860 B.n859 585
R664 B.n861 B.n860 585
R665 B.n858 B.n37 585
R666 B.n37 B.n36 585
R667 B.n857 B.n856 585
R668 B.n856 B.n855 585
R669 B.n39 B.n38 585
R670 B.n854 B.n39 585
R671 B.n852 B.n851 585
R672 B.n853 B.n852 585
R673 B.n850 B.n44 585
R674 B.n44 B.n43 585
R675 B.n849 B.n848 585
R676 B.n848 B.n847 585
R677 B.n46 B.n45 585
R678 B.n846 B.n46 585
R679 B.n844 B.n843 585
R680 B.n845 B.n844 585
R681 B.n842 B.n51 585
R682 B.n51 B.n50 585
R683 B.n841 B.n840 585
R684 B.n840 B.n839 585
R685 B.n53 B.n52 585
R686 B.n838 B.n53 585
R687 B.n836 B.n835 585
R688 B.n837 B.n836 585
R689 B.n834 B.n58 585
R690 B.n58 B.n57 585
R691 B.n833 B.n832 585
R692 B.n832 B.n831 585
R693 B.n60 B.n59 585
R694 B.n830 B.n60 585
R695 B.n828 B.n827 585
R696 B.n829 B.n828 585
R697 B.n826 B.n65 585
R698 B.n65 B.n64 585
R699 B.n825 B.n824 585
R700 B.n824 B.n823 585
R701 B.n67 B.n66 585
R702 B.n822 B.n67 585
R703 B.n820 B.n819 585
R704 B.n821 B.n820 585
R705 B.n818 B.n71 585
R706 B.n74 B.n71 585
R707 B.n817 B.n816 585
R708 B.n816 B.n815 585
R709 B.n73 B.n72 585
R710 B.n814 B.n73 585
R711 B.n812 B.n811 585
R712 B.n813 B.n812 585
R713 B.n810 B.n79 585
R714 B.n79 B.n78 585
R715 B.n809 B.n808 585
R716 B.n808 B.n807 585
R717 B.n81 B.n80 585
R718 B.n806 B.n81 585
R719 B.n804 B.n803 585
R720 B.n805 B.n804 585
R721 B.n802 B.n86 585
R722 B.n86 B.n85 585
R723 B.n801 B.n800 585
R724 B.n800 B.n799 585
R725 B.n88 B.n87 585
R726 B.n798 B.n88 585
R727 B.n796 B.n795 585
R728 B.n797 B.n796 585
R729 B.n794 B.n93 585
R730 B.n93 B.n92 585
R731 B.n793 B.n792 585
R732 B.n792 B.n791 585
R733 B.n95 B.n94 585
R734 B.n790 B.n95 585
R735 B.n788 B.n787 585
R736 B.n789 B.n788 585
R737 B.n786 B.n100 585
R738 B.n100 B.n99 585
R739 B.n785 B.n784 585
R740 B.n784 B.n783 585
R741 B.n102 B.n101 585
R742 B.n782 B.n102 585
R743 B.n780 B.n779 585
R744 B.n781 B.n780 585
R745 B.n778 B.n107 585
R746 B.n107 B.n106 585
R747 B.n777 B.n776 585
R748 B.n776 B.n775 585
R749 B.n109 B.n108 585
R750 B.n774 B.n109 585
R751 B.n897 B.n896 585
R752 B.n896 B.n895 585
R753 B.n504 B.n365 526.135
R754 B.n145 B.n109 526.135
R755 B.n507 B.n367 526.135
R756 B.n771 B.n111 526.135
R757 B.n773 B.n772 256.663
R758 B.n773 B.n137 256.663
R759 B.n773 B.n136 256.663
R760 B.n773 B.n135 256.663
R761 B.n773 B.n134 256.663
R762 B.n773 B.n133 256.663
R763 B.n773 B.n132 256.663
R764 B.n773 B.n131 256.663
R765 B.n773 B.n130 256.663
R766 B.n773 B.n129 256.663
R767 B.n773 B.n128 256.663
R768 B.n773 B.n127 256.663
R769 B.n773 B.n126 256.663
R770 B.n773 B.n125 256.663
R771 B.n773 B.n124 256.663
R772 B.n773 B.n123 256.663
R773 B.n773 B.n122 256.663
R774 B.n773 B.n121 256.663
R775 B.n773 B.n120 256.663
R776 B.n773 B.n119 256.663
R777 B.n773 B.n118 256.663
R778 B.n773 B.n117 256.663
R779 B.n773 B.n116 256.663
R780 B.n773 B.n115 256.663
R781 B.n773 B.n114 256.663
R782 B.n773 B.n113 256.663
R783 B.n773 B.n112 256.663
R784 B.n506 B.n505 256.663
R785 B.n506 B.n370 256.663
R786 B.n506 B.n371 256.663
R787 B.n506 B.n372 256.663
R788 B.n506 B.n373 256.663
R789 B.n506 B.n374 256.663
R790 B.n506 B.n375 256.663
R791 B.n506 B.n376 256.663
R792 B.n506 B.n377 256.663
R793 B.n506 B.n378 256.663
R794 B.n506 B.n379 256.663
R795 B.n506 B.n380 256.663
R796 B.n506 B.n381 256.663
R797 B.n506 B.n382 256.663
R798 B.n506 B.n383 256.663
R799 B.n506 B.n384 256.663
R800 B.n506 B.n385 256.663
R801 B.n506 B.n386 256.663
R802 B.n506 B.n387 256.663
R803 B.n506 B.n388 256.663
R804 B.n506 B.n389 256.663
R805 B.n506 B.n390 256.663
R806 B.n506 B.n391 256.663
R807 B.n506 B.n392 256.663
R808 B.n506 B.n393 256.663
R809 B.n506 B.n394 256.663
R810 B.n399 B.t12 248.968
R811 B.n397 B.t16 248.968
R812 B.n142 B.t8 248.968
R813 B.n139 B.t19 248.968
R814 B.n513 B.n365 163.367
R815 B.n513 B.n363 163.367
R816 B.n517 B.n363 163.367
R817 B.n517 B.n357 163.367
R818 B.n525 B.n357 163.367
R819 B.n525 B.n355 163.367
R820 B.n529 B.n355 163.367
R821 B.n529 B.n349 163.367
R822 B.n537 B.n349 163.367
R823 B.n537 B.n347 163.367
R824 B.n541 B.n347 163.367
R825 B.n541 B.n341 163.367
R826 B.n549 B.n341 163.367
R827 B.n549 B.n339 163.367
R828 B.n553 B.n339 163.367
R829 B.n553 B.n333 163.367
R830 B.n561 B.n333 163.367
R831 B.n561 B.n331 163.367
R832 B.n565 B.n331 163.367
R833 B.n565 B.n325 163.367
R834 B.n574 B.n325 163.367
R835 B.n574 B.n323 163.367
R836 B.n578 B.n323 163.367
R837 B.n578 B.n318 163.367
R838 B.n586 B.n318 163.367
R839 B.n586 B.n316 163.367
R840 B.n590 B.n316 163.367
R841 B.n590 B.n310 163.367
R842 B.n598 B.n310 163.367
R843 B.n598 B.n308 163.367
R844 B.n602 B.n308 163.367
R845 B.n602 B.n302 163.367
R846 B.n610 B.n302 163.367
R847 B.n610 B.n300 163.367
R848 B.n614 B.n300 163.367
R849 B.n614 B.n294 163.367
R850 B.n622 B.n294 163.367
R851 B.n622 B.n292 163.367
R852 B.n626 B.n292 163.367
R853 B.n626 B.n286 163.367
R854 B.n634 B.n286 163.367
R855 B.n634 B.n284 163.367
R856 B.n638 B.n284 163.367
R857 B.n638 B.n278 163.367
R858 B.n646 B.n278 163.367
R859 B.n646 B.n276 163.367
R860 B.n650 B.n276 163.367
R861 B.n650 B.n270 163.367
R862 B.n658 B.n270 163.367
R863 B.n658 B.n268 163.367
R864 B.n662 B.n268 163.367
R865 B.n662 B.n262 163.367
R866 B.n671 B.n262 163.367
R867 B.n671 B.n260 163.367
R868 B.n675 B.n260 163.367
R869 B.n675 B.n255 163.367
R870 B.n684 B.n255 163.367
R871 B.n684 B.n253 163.367
R872 B.n688 B.n253 163.367
R873 B.n688 B.n2 163.367
R874 B.n896 B.n2 163.367
R875 B.n896 B.n3 163.367
R876 B.n892 B.n3 163.367
R877 B.n892 B.n9 163.367
R878 B.n888 B.n9 163.367
R879 B.n888 B.n11 163.367
R880 B.n884 B.n11 163.367
R881 B.n884 B.n15 163.367
R882 B.n880 B.n15 163.367
R883 B.n880 B.n17 163.367
R884 B.n876 B.n17 163.367
R885 B.n876 B.n23 163.367
R886 B.n872 B.n23 163.367
R887 B.n872 B.n25 163.367
R888 B.n868 B.n25 163.367
R889 B.n868 B.n30 163.367
R890 B.n864 B.n30 163.367
R891 B.n864 B.n32 163.367
R892 B.n860 B.n32 163.367
R893 B.n860 B.n37 163.367
R894 B.n856 B.n37 163.367
R895 B.n856 B.n39 163.367
R896 B.n852 B.n39 163.367
R897 B.n852 B.n44 163.367
R898 B.n848 B.n44 163.367
R899 B.n848 B.n46 163.367
R900 B.n844 B.n46 163.367
R901 B.n844 B.n51 163.367
R902 B.n840 B.n51 163.367
R903 B.n840 B.n53 163.367
R904 B.n836 B.n53 163.367
R905 B.n836 B.n58 163.367
R906 B.n832 B.n58 163.367
R907 B.n832 B.n60 163.367
R908 B.n828 B.n60 163.367
R909 B.n828 B.n65 163.367
R910 B.n824 B.n65 163.367
R911 B.n824 B.n67 163.367
R912 B.n820 B.n67 163.367
R913 B.n820 B.n71 163.367
R914 B.n816 B.n71 163.367
R915 B.n816 B.n73 163.367
R916 B.n812 B.n73 163.367
R917 B.n812 B.n79 163.367
R918 B.n808 B.n79 163.367
R919 B.n808 B.n81 163.367
R920 B.n804 B.n81 163.367
R921 B.n804 B.n86 163.367
R922 B.n800 B.n86 163.367
R923 B.n800 B.n88 163.367
R924 B.n796 B.n88 163.367
R925 B.n796 B.n93 163.367
R926 B.n792 B.n93 163.367
R927 B.n792 B.n95 163.367
R928 B.n788 B.n95 163.367
R929 B.n788 B.n100 163.367
R930 B.n784 B.n100 163.367
R931 B.n784 B.n102 163.367
R932 B.n780 B.n102 163.367
R933 B.n780 B.n107 163.367
R934 B.n776 B.n107 163.367
R935 B.n776 B.n109 163.367
R936 B.n396 B.n395 163.367
R937 B.n499 B.n395 163.367
R938 B.n497 B.n496 163.367
R939 B.n493 B.n492 163.367
R940 B.n489 B.n488 163.367
R941 B.n485 B.n484 163.367
R942 B.n481 B.n480 163.367
R943 B.n477 B.n476 163.367
R944 B.n473 B.n472 163.367
R945 B.n469 B.n468 163.367
R946 B.n465 B.n464 163.367
R947 B.n460 B.n459 163.367
R948 B.n456 B.n455 163.367
R949 B.n452 B.n451 163.367
R950 B.n448 B.n447 163.367
R951 B.n444 B.n443 163.367
R952 B.n439 B.n438 163.367
R953 B.n435 B.n434 163.367
R954 B.n431 B.n430 163.367
R955 B.n427 B.n426 163.367
R956 B.n423 B.n422 163.367
R957 B.n419 B.n418 163.367
R958 B.n415 B.n414 163.367
R959 B.n411 B.n410 163.367
R960 B.n407 B.n406 163.367
R961 B.n403 B.n402 163.367
R962 B.n507 B.n369 163.367
R963 B.n511 B.n367 163.367
R964 B.n511 B.n361 163.367
R965 B.n519 B.n361 163.367
R966 B.n519 B.n359 163.367
R967 B.n523 B.n359 163.367
R968 B.n523 B.n352 163.367
R969 B.n531 B.n352 163.367
R970 B.n531 B.n350 163.367
R971 B.n535 B.n350 163.367
R972 B.n535 B.n345 163.367
R973 B.n543 B.n345 163.367
R974 B.n543 B.n343 163.367
R975 B.n547 B.n343 163.367
R976 B.n547 B.n337 163.367
R977 B.n555 B.n337 163.367
R978 B.n555 B.n335 163.367
R979 B.n559 B.n335 163.367
R980 B.n559 B.n329 163.367
R981 B.n567 B.n329 163.367
R982 B.n567 B.n327 163.367
R983 B.n571 B.n327 163.367
R984 B.n571 B.n322 163.367
R985 B.n580 B.n322 163.367
R986 B.n580 B.n320 163.367
R987 B.n584 B.n320 163.367
R988 B.n584 B.n314 163.367
R989 B.n592 B.n314 163.367
R990 B.n592 B.n312 163.367
R991 B.n596 B.n312 163.367
R992 B.n596 B.n305 163.367
R993 B.n604 B.n305 163.367
R994 B.n604 B.n303 163.367
R995 B.n608 B.n303 163.367
R996 B.n608 B.n298 163.367
R997 B.n616 B.n298 163.367
R998 B.n616 B.n296 163.367
R999 B.n620 B.n296 163.367
R1000 B.n620 B.n290 163.367
R1001 B.n628 B.n290 163.367
R1002 B.n628 B.n288 163.367
R1003 B.n632 B.n288 163.367
R1004 B.n632 B.n282 163.367
R1005 B.n640 B.n282 163.367
R1006 B.n640 B.n280 163.367
R1007 B.n644 B.n280 163.367
R1008 B.n644 B.n274 163.367
R1009 B.n652 B.n274 163.367
R1010 B.n652 B.n272 163.367
R1011 B.n656 B.n272 163.367
R1012 B.n656 B.n266 163.367
R1013 B.n664 B.n266 163.367
R1014 B.n664 B.n264 163.367
R1015 B.n668 B.n264 163.367
R1016 B.n668 B.n259 163.367
R1017 B.n677 B.n259 163.367
R1018 B.n677 B.n257 163.367
R1019 B.n682 B.n257 163.367
R1020 B.n682 B.n251 163.367
R1021 B.n690 B.n251 163.367
R1022 B.n691 B.n690 163.367
R1023 B.n691 B.n5 163.367
R1024 B.n6 B.n5 163.367
R1025 B.n7 B.n6 163.367
R1026 B.n696 B.n7 163.367
R1027 B.n696 B.n12 163.367
R1028 B.n13 B.n12 163.367
R1029 B.n14 B.n13 163.367
R1030 B.n701 B.n14 163.367
R1031 B.n701 B.n19 163.367
R1032 B.n20 B.n19 163.367
R1033 B.n21 B.n20 163.367
R1034 B.n706 B.n21 163.367
R1035 B.n706 B.n26 163.367
R1036 B.n27 B.n26 163.367
R1037 B.n28 B.n27 163.367
R1038 B.n711 B.n28 163.367
R1039 B.n711 B.n33 163.367
R1040 B.n34 B.n33 163.367
R1041 B.n35 B.n34 163.367
R1042 B.n716 B.n35 163.367
R1043 B.n716 B.n40 163.367
R1044 B.n41 B.n40 163.367
R1045 B.n42 B.n41 163.367
R1046 B.n721 B.n42 163.367
R1047 B.n721 B.n47 163.367
R1048 B.n48 B.n47 163.367
R1049 B.n49 B.n48 163.367
R1050 B.n726 B.n49 163.367
R1051 B.n726 B.n54 163.367
R1052 B.n55 B.n54 163.367
R1053 B.n56 B.n55 163.367
R1054 B.n731 B.n56 163.367
R1055 B.n731 B.n61 163.367
R1056 B.n62 B.n61 163.367
R1057 B.n63 B.n62 163.367
R1058 B.n736 B.n63 163.367
R1059 B.n736 B.n68 163.367
R1060 B.n69 B.n68 163.367
R1061 B.n70 B.n69 163.367
R1062 B.n741 B.n70 163.367
R1063 B.n741 B.n75 163.367
R1064 B.n76 B.n75 163.367
R1065 B.n77 B.n76 163.367
R1066 B.n746 B.n77 163.367
R1067 B.n746 B.n82 163.367
R1068 B.n83 B.n82 163.367
R1069 B.n84 B.n83 163.367
R1070 B.n751 B.n84 163.367
R1071 B.n751 B.n89 163.367
R1072 B.n90 B.n89 163.367
R1073 B.n91 B.n90 163.367
R1074 B.n756 B.n91 163.367
R1075 B.n756 B.n96 163.367
R1076 B.n97 B.n96 163.367
R1077 B.n98 B.n97 163.367
R1078 B.n761 B.n98 163.367
R1079 B.n761 B.n103 163.367
R1080 B.n104 B.n103 163.367
R1081 B.n105 B.n104 163.367
R1082 B.n766 B.n105 163.367
R1083 B.n766 B.n110 163.367
R1084 B.n111 B.n110 163.367
R1085 B.n149 B.n148 163.367
R1086 B.n153 B.n152 163.367
R1087 B.n157 B.n156 163.367
R1088 B.n161 B.n160 163.367
R1089 B.n165 B.n164 163.367
R1090 B.n169 B.n168 163.367
R1091 B.n173 B.n172 163.367
R1092 B.n177 B.n176 163.367
R1093 B.n181 B.n180 163.367
R1094 B.n185 B.n184 163.367
R1095 B.n189 B.n188 163.367
R1096 B.n193 B.n192 163.367
R1097 B.n197 B.n196 163.367
R1098 B.n201 B.n200 163.367
R1099 B.n205 B.n204 163.367
R1100 B.n209 B.n208 163.367
R1101 B.n213 B.n212 163.367
R1102 B.n217 B.n216 163.367
R1103 B.n221 B.n220 163.367
R1104 B.n225 B.n224 163.367
R1105 B.n229 B.n228 163.367
R1106 B.n233 B.n232 163.367
R1107 B.n237 B.n236 163.367
R1108 B.n241 B.n240 163.367
R1109 B.n245 B.n244 163.367
R1110 B.n247 B.n138 163.367
R1111 B.n399 B.t15 139.623
R1112 B.n139 B.t20 139.623
R1113 B.n397 B.t18 139.617
R1114 B.n142 B.t10 139.617
R1115 B.n506 B.n366 130.379
R1116 B.n774 B.n773 130.379
R1117 B.n505 B.n504 71.676
R1118 B.n499 B.n370 71.676
R1119 B.n496 B.n371 71.676
R1120 B.n492 B.n372 71.676
R1121 B.n488 B.n373 71.676
R1122 B.n484 B.n374 71.676
R1123 B.n480 B.n375 71.676
R1124 B.n476 B.n376 71.676
R1125 B.n472 B.n377 71.676
R1126 B.n468 B.n378 71.676
R1127 B.n464 B.n379 71.676
R1128 B.n459 B.n380 71.676
R1129 B.n455 B.n381 71.676
R1130 B.n451 B.n382 71.676
R1131 B.n447 B.n383 71.676
R1132 B.n443 B.n384 71.676
R1133 B.n438 B.n385 71.676
R1134 B.n434 B.n386 71.676
R1135 B.n430 B.n387 71.676
R1136 B.n426 B.n388 71.676
R1137 B.n422 B.n389 71.676
R1138 B.n418 B.n390 71.676
R1139 B.n414 B.n391 71.676
R1140 B.n410 B.n392 71.676
R1141 B.n406 B.n393 71.676
R1142 B.n402 B.n394 71.676
R1143 B.n145 B.n112 71.676
R1144 B.n149 B.n113 71.676
R1145 B.n153 B.n114 71.676
R1146 B.n157 B.n115 71.676
R1147 B.n161 B.n116 71.676
R1148 B.n165 B.n117 71.676
R1149 B.n169 B.n118 71.676
R1150 B.n173 B.n119 71.676
R1151 B.n177 B.n120 71.676
R1152 B.n181 B.n121 71.676
R1153 B.n185 B.n122 71.676
R1154 B.n189 B.n123 71.676
R1155 B.n193 B.n124 71.676
R1156 B.n197 B.n125 71.676
R1157 B.n201 B.n126 71.676
R1158 B.n205 B.n127 71.676
R1159 B.n209 B.n128 71.676
R1160 B.n213 B.n129 71.676
R1161 B.n217 B.n130 71.676
R1162 B.n221 B.n131 71.676
R1163 B.n225 B.n132 71.676
R1164 B.n229 B.n133 71.676
R1165 B.n233 B.n134 71.676
R1166 B.n237 B.n135 71.676
R1167 B.n241 B.n136 71.676
R1168 B.n245 B.n137 71.676
R1169 B.n772 B.n138 71.676
R1170 B.n772 B.n771 71.676
R1171 B.n247 B.n137 71.676
R1172 B.n244 B.n136 71.676
R1173 B.n240 B.n135 71.676
R1174 B.n236 B.n134 71.676
R1175 B.n232 B.n133 71.676
R1176 B.n228 B.n132 71.676
R1177 B.n224 B.n131 71.676
R1178 B.n220 B.n130 71.676
R1179 B.n216 B.n129 71.676
R1180 B.n212 B.n128 71.676
R1181 B.n208 B.n127 71.676
R1182 B.n204 B.n126 71.676
R1183 B.n200 B.n125 71.676
R1184 B.n196 B.n124 71.676
R1185 B.n192 B.n123 71.676
R1186 B.n188 B.n122 71.676
R1187 B.n184 B.n121 71.676
R1188 B.n180 B.n120 71.676
R1189 B.n176 B.n119 71.676
R1190 B.n172 B.n118 71.676
R1191 B.n168 B.n117 71.676
R1192 B.n164 B.n116 71.676
R1193 B.n160 B.n115 71.676
R1194 B.n156 B.n114 71.676
R1195 B.n152 B.n113 71.676
R1196 B.n148 B.n112 71.676
R1197 B.n505 B.n396 71.676
R1198 B.n497 B.n370 71.676
R1199 B.n493 B.n371 71.676
R1200 B.n489 B.n372 71.676
R1201 B.n485 B.n373 71.676
R1202 B.n481 B.n374 71.676
R1203 B.n477 B.n375 71.676
R1204 B.n473 B.n376 71.676
R1205 B.n469 B.n377 71.676
R1206 B.n465 B.n378 71.676
R1207 B.n460 B.n379 71.676
R1208 B.n456 B.n380 71.676
R1209 B.n452 B.n381 71.676
R1210 B.n448 B.n382 71.676
R1211 B.n444 B.n383 71.676
R1212 B.n439 B.n384 71.676
R1213 B.n435 B.n385 71.676
R1214 B.n431 B.n386 71.676
R1215 B.n427 B.n387 71.676
R1216 B.n423 B.n388 71.676
R1217 B.n419 B.n389 71.676
R1218 B.n415 B.n390 71.676
R1219 B.n411 B.n391 71.676
R1220 B.n407 B.n392 71.676
R1221 B.n403 B.n393 71.676
R1222 B.n394 B.n369 71.676
R1223 B.n400 B.n399 69.8187
R1224 B.n398 B.n397 69.8187
R1225 B.n143 B.n142 69.8187
R1226 B.n140 B.n139 69.8187
R1227 B.n512 B.n366 69.8092
R1228 B.n512 B.n362 69.8092
R1229 B.n518 B.n362 69.8092
R1230 B.n518 B.n358 69.8092
R1231 B.n524 B.n358 69.8092
R1232 B.n524 B.n353 69.8092
R1233 B.n530 B.n353 69.8092
R1234 B.n530 B.n354 69.8092
R1235 B.n536 B.n346 69.8092
R1236 B.n542 B.n346 69.8092
R1237 B.n542 B.n342 69.8092
R1238 B.n548 B.n342 69.8092
R1239 B.n548 B.n338 69.8092
R1240 B.n554 B.n338 69.8092
R1241 B.n554 B.n334 69.8092
R1242 B.n560 B.n334 69.8092
R1243 B.n560 B.n330 69.8092
R1244 B.n566 B.n330 69.8092
R1245 B.n566 B.n326 69.8092
R1246 B.n573 B.n326 69.8092
R1247 B.n573 B.n572 69.8092
R1248 B.n579 B.n319 69.8092
R1249 B.n585 B.n319 69.8092
R1250 B.n585 B.n315 69.8092
R1251 B.n591 B.n315 69.8092
R1252 B.n591 B.n311 69.8092
R1253 B.n597 B.n311 69.8092
R1254 B.n597 B.n306 69.8092
R1255 B.n603 B.n306 69.8092
R1256 B.n603 B.n307 69.8092
R1257 B.n609 B.n299 69.8092
R1258 B.n615 B.n299 69.8092
R1259 B.n615 B.n295 69.8092
R1260 B.n621 B.n295 69.8092
R1261 B.n621 B.n291 69.8092
R1262 B.n627 B.n291 69.8092
R1263 B.n627 B.n287 69.8092
R1264 B.n633 B.n287 69.8092
R1265 B.n633 B.n283 69.8092
R1266 B.n639 B.n283 69.8092
R1267 B.n645 B.n279 69.8092
R1268 B.n645 B.n275 69.8092
R1269 B.n651 B.n275 69.8092
R1270 B.n651 B.n271 69.8092
R1271 B.n657 B.n271 69.8092
R1272 B.n657 B.n267 69.8092
R1273 B.n663 B.n267 69.8092
R1274 B.n663 B.n263 69.8092
R1275 B.n670 B.n263 69.8092
R1276 B.n670 B.n669 69.8092
R1277 B.n676 B.n256 69.8092
R1278 B.n683 B.n256 69.8092
R1279 B.n683 B.n252 69.8092
R1280 B.n689 B.n252 69.8092
R1281 B.n689 B.n4 69.8092
R1282 B.n895 B.n4 69.8092
R1283 B.n895 B.n894 69.8092
R1284 B.n894 B.n893 69.8092
R1285 B.n893 B.n8 69.8092
R1286 B.n887 B.n8 69.8092
R1287 B.n887 B.n886 69.8092
R1288 B.n886 B.n885 69.8092
R1289 B.n879 B.n18 69.8092
R1290 B.n879 B.n878 69.8092
R1291 B.n878 B.n877 69.8092
R1292 B.n877 B.n22 69.8092
R1293 B.n871 B.n22 69.8092
R1294 B.n871 B.n870 69.8092
R1295 B.n870 B.n869 69.8092
R1296 B.n869 B.n29 69.8092
R1297 B.n863 B.n29 69.8092
R1298 B.n863 B.n862 69.8092
R1299 B.n861 B.n36 69.8092
R1300 B.n855 B.n36 69.8092
R1301 B.n855 B.n854 69.8092
R1302 B.n854 B.n853 69.8092
R1303 B.n853 B.n43 69.8092
R1304 B.n847 B.n43 69.8092
R1305 B.n847 B.n846 69.8092
R1306 B.n846 B.n845 69.8092
R1307 B.n845 B.n50 69.8092
R1308 B.n839 B.n50 69.8092
R1309 B.n838 B.n837 69.8092
R1310 B.n837 B.n57 69.8092
R1311 B.n831 B.n57 69.8092
R1312 B.n831 B.n830 69.8092
R1313 B.n830 B.n829 69.8092
R1314 B.n829 B.n64 69.8092
R1315 B.n823 B.n64 69.8092
R1316 B.n823 B.n822 69.8092
R1317 B.n822 B.n821 69.8092
R1318 B.n815 B.n74 69.8092
R1319 B.n815 B.n814 69.8092
R1320 B.n814 B.n813 69.8092
R1321 B.n813 B.n78 69.8092
R1322 B.n807 B.n78 69.8092
R1323 B.n807 B.n806 69.8092
R1324 B.n806 B.n805 69.8092
R1325 B.n805 B.n85 69.8092
R1326 B.n799 B.n85 69.8092
R1327 B.n799 B.n798 69.8092
R1328 B.n798 B.n797 69.8092
R1329 B.n797 B.n92 69.8092
R1330 B.n791 B.n92 69.8092
R1331 B.n790 B.n789 69.8092
R1332 B.n789 B.n99 69.8092
R1333 B.n783 B.n99 69.8092
R1334 B.n783 B.n782 69.8092
R1335 B.n782 B.n781 69.8092
R1336 B.n781 B.n106 69.8092
R1337 B.n775 B.n106 69.8092
R1338 B.n775 B.n774 69.8092
R1339 B.n400 B.t14 69.8041
R1340 B.n140 B.t21 69.8041
R1341 B.n398 B.t17 69.7983
R1342 B.n143 B.t11 69.7983
R1343 B.n307 B.t5 64.6762
R1344 B.t6 B.n838 64.6762
R1345 B.n676 B.t3 62.623
R1346 B.n885 B.t2 62.623
R1347 B.n441 B.n400 59.5399
R1348 B.n462 B.n398 59.5399
R1349 B.n144 B.n143 59.5399
R1350 B.n141 B.n140 59.5399
R1351 B.n579 B.t7 46.1974
R1352 B.n821 B.t0 46.1974
R1353 B.n354 B.t13 37.9846
R1354 B.t9 B.n790 37.9846
R1355 B.n639 B.t1 35.9314
R1356 B.t4 B.n861 35.9314
R1357 B.n146 B.n108 34.1859
R1358 B.n770 B.n769 34.1859
R1359 B.n509 B.n508 34.1859
R1360 B.n503 B.n364 34.1859
R1361 B.t1 B.n279 33.8782
R1362 B.n862 B.t4 33.8782
R1363 B.n536 B.t13 31.825
R1364 B.n791 B.t9 31.825
R1365 B.n572 B.t7 23.6123
R1366 B.n74 B.t0 23.6123
R1367 B B.n897 18.0485
R1368 B.n147 B.n146 10.6151
R1369 B.n150 B.n147 10.6151
R1370 B.n151 B.n150 10.6151
R1371 B.n154 B.n151 10.6151
R1372 B.n155 B.n154 10.6151
R1373 B.n158 B.n155 10.6151
R1374 B.n159 B.n158 10.6151
R1375 B.n162 B.n159 10.6151
R1376 B.n163 B.n162 10.6151
R1377 B.n166 B.n163 10.6151
R1378 B.n167 B.n166 10.6151
R1379 B.n170 B.n167 10.6151
R1380 B.n171 B.n170 10.6151
R1381 B.n174 B.n171 10.6151
R1382 B.n175 B.n174 10.6151
R1383 B.n178 B.n175 10.6151
R1384 B.n179 B.n178 10.6151
R1385 B.n182 B.n179 10.6151
R1386 B.n183 B.n182 10.6151
R1387 B.n186 B.n183 10.6151
R1388 B.n187 B.n186 10.6151
R1389 B.n191 B.n190 10.6151
R1390 B.n194 B.n191 10.6151
R1391 B.n195 B.n194 10.6151
R1392 B.n198 B.n195 10.6151
R1393 B.n199 B.n198 10.6151
R1394 B.n202 B.n199 10.6151
R1395 B.n203 B.n202 10.6151
R1396 B.n206 B.n203 10.6151
R1397 B.n207 B.n206 10.6151
R1398 B.n211 B.n210 10.6151
R1399 B.n214 B.n211 10.6151
R1400 B.n215 B.n214 10.6151
R1401 B.n218 B.n215 10.6151
R1402 B.n219 B.n218 10.6151
R1403 B.n222 B.n219 10.6151
R1404 B.n223 B.n222 10.6151
R1405 B.n226 B.n223 10.6151
R1406 B.n227 B.n226 10.6151
R1407 B.n230 B.n227 10.6151
R1408 B.n231 B.n230 10.6151
R1409 B.n234 B.n231 10.6151
R1410 B.n235 B.n234 10.6151
R1411 B.n238 B.n235 10.6151
R1412 B.n239 B.n238 10.6151
R1413 B.n242 B.n239 10.6151
R1414 B.n243 B.n242 10.6151
R1415 B.n246 B.n243 10.6151
R1416 B.n248 B.n246 10.6151
R1417 B.n249 B.n248 10.6151
R1418 B.n770 B.n249 10.6151
R1419 B.n510 B.n509 10.6151
R1420 B.n510 B.n360 10.6151
R1421 B.n520 B.n360 10.6151
R1422 B.n521 B.n520 10.6151
R1423 B.n522 B.n521 10.6151
R1424 B.n522 B.n351 10.6151
R1425 B.n532 B.n351 10.6151
R1426 B.n533 B.n532 10.6151
R1427 B.n534 B.n533 10.6151
R1428 B.n534 B.n344 10.6151
R1429 B.n544 B.n344 10.6151
R1430 B.n545 B.n544 10.6151
R1431 B.n546 B.n545 10.6151
R1432 B.n546 B.n336 10.6151
R1433 B.n556 B.n336 10.6151
R1434 B.n557 B.n556 10.6151
R1435 B.n558 B.n557 10.6151
R1436 B.n558 B.n328 10.6151
R1437 B.n568 B.n328 10.6151
R1438 B.n569 B.n568 10.6151
R1439 B.n570 B.n569 10.6151
R1440 B.n570 B.n321 10.6151
R1441 B.n581 B.n321 10.6151
R1442 B.n582 B.n581 10.6151
R1443 B.n583 B.n582 10.6151
R1444 B.n583 B.n313 10.6151
R1445 B.n593 B.n313 10.6151
R1446 B.n594 B.n593 10.6151
R1447 B.n595 B.n594 10.6151
R1448 B.n595 B.n304 10.6151
R1449 B.n605 B.n304 10.6151
R1450 B.n606 B.n605 10.6151
R1451 B.n607 B.n606 10.6151
R1452 B.n607 B.n297 10.6151
R1453 B.n617 B.n297 10.6151
R1454 B.n618 B.n617 10.6151
R1455 B.n619 B.n618 10.6151
R1456 B.n619 B.n289 10.6151
R1457 B.n629 B.n289 10.6151
R1458 B.n630 B.n629 10.6151
R1459 B.n631 B.n630 10.6151
R1460 B.n631 B.n281 10.6151
R1461 B.n641 B.n281 10.6151
R1462 B.n642 B.n641 10.6151
R1463 B.n643 B.n642 10.6151
R1464 B.n643 B.n273 10.6151
R1465 B.n653 B.n273 10.6151
R1466 B.n654 B.n653 10.6151
R1467 B.n655 B.n654 10.6151
R1468 B.n655 B.n265 10.6151
R1469 B.n665 B.n265 10.6151
R1470 B.n666 B.n665 10.6151
R1471 B.n667 B.n666 10.6151
R1472 B.n667 B.n258 10.6151
R1473 B.n678 B.n258 10.6151
R1474 B.n679 B.n678 10.6151
R1475 B.n681 B.n679 10.6151
R1476 B.n681 B.n680 10.6151
R1477 B.n680 B.n250 10.6151
R1478 B.n692 B.n250 10.6151
R1479 B.n693 B.n692 10.6151
R1480 B.n694 B.n693 10.6151
R1481 B.n695 B.n694 10.6151
R1482 B.n697 B.n695 10.6151
R1483 B.n698 B.n697 10.6151
R1484 B.n699 B.n698 10.6151
R1485 B.n700 B.n699 10.6151
R1486 B.n702 B.n700 10.6151
R1487 B.n703 B.n702 10.6151
R1488 B.n704 B.n703 10.6151
R1489 B.n705 B.n704 10.6151
R1490 B.n707 B.n705 10.6151
R1491 B.n708 B.n707 10.6151
R1492 B.n709 B.n708 10.6151
R1493 B.n710 B.n709 10.6151
R1494 B.n712 B.n710 10.6151
R1495 B.n713 B.n712 10.6151
R1496 B.n714 B.n713 10.6151
R1497 B.n715 B.n714 10.6151
R1498 B.n717 B.n715 10.6151
R1499 B.n718 B.n717 10.6151
R1500 B.n719 B.n718 10.6151
R1501 B.n720 B.n719 10.6151
R1502 B.n722 B.n720 10.6151
R1503 B.n723 B.n722 10.6151
R1504 B.n724 B.n723 10.6151
R1505 B.n725 B.n724 10.6151
R1506 B.n727 B.n725 10.6151
R1507 B.n728 B.n727 10.6151
R1508 B.n729 B.n728 10.6151
R1509 B.n730 B.n729 10.6151
R1510 B.n732 B.n730 10.6151
R1511 B.n733 B.n732 10.6151
R1512 B.n734 B.n733 10.6151
R1513 B.n735 B.n734 10.6151
R1514 B.n737 B.n735 10.6151
R1515 B.n738 B.n737 10.6151
R1516 B.n739 B.n738 10.6151
R1517 B.n740 B.n739 10.6151
R1518 B.n742 B.n740 10.6151
R1519 B.n743 B.n742 10.6151
R1520 B.n744 B.n743 10.6151
R1521 B.n745 B.n744 10.6151
R1522 B.n747 B.n745 10.6151
R1523 B.n748 B.n747 10.6151
R1524 B.n749 B.n748 10.6151
R1525 B.n750 B.n749 10.6151
R1526 B.n752 B.n750 10.6151
R1527 B.n753 B.n752 10.6151
R1528 B.n754 B.n753 10.6151
R1529 B.n755 B.n754 10.6151
R1530 B.n757 B.n755 10.6151
R1531 B.n758 B.n757 10.6151
R1532 B.n759 B.n758 10.6151
R1533 B.n760 B.n759 10.6151
R1534 B.n762 B.n760 10.6151
R1535 B.n763 B.n762 10.6151
R1536 B.n764 B.n763 10.6151
R1537 B.n765 B.n764 10.6151
R1538 B.n767 B.n765 10.6151
R1539 B.n768 B.n767 10.6151
R1540 B.n769 B.n768 10.6151
R1541 B.n503 B.n502 10.6151
R1542 B.n502 B.n501 10.6151
R1543 B.n501 B.n500 10.6151
R1544 B.n500 B.n498 10.6151
R1545 B.n498 B.n495 10.6151
R1546 B.n495 B.n494 10.6151
R1547 B.n494 B.n491 10.6151
R1548 B.n491 B.n490 10.6151
R1549 B.n490 B.n487 10.6151
R1550 B.n487 B.n486 10.6151
R1551 B.n486 B.n483 10.6151
R1552 B.n483 B.n482 10.6151
R1553 B.n482 B.n479 10.6151
R1554 B.n479 B.n478 10.6151
R1555 B.n478 B.n475 10.6151
R1556 B.n475 B.n474 10.6151
R1557 B.n474 B.n471 10.6151
R1558 B.n471 B.n470 10.6151
R1559 B.n470 B.n467 10.6151
R1560 B.n467 B.n466 10.6151
R1561 B.n466 B.n463 10.6151
R1562 B.n461 B.n458 10.6151
R1563 B.n458 B.n457 10.6151
R1564 B.n457 B.n454 10.6151
R1565 B.n454 B.n453 10.6151
R1566 B.n453 B.n450 10.6151
R1567 B.n450 B.n449 10.6151
R1568 B.n449 B.n446 10.6151
R1569 B.n446 B.n445 10.6151
R1570 B.n445 B.n442 10.6151
R1571 B.n440 B.n437 10.6151
R1572 B.n437 B.n436 10.6151
R1573 B.n436 B.n433 10.6151
R1574 B.n433 B.n432 10.6151
R1575 B.n432 B.n429 10.6151
R1576 B.n429 B.n428 10.6151
R1577 B.n428 B.n425 10.6151
R1578 B.n425 B.n424 10.6151
R1579 B.n424 B.n421 10.6151
R1580 B.n421 B.n420 10.6151
R1581 B.n420 B.n417 10.6151
R1582 B.n417 B.n416 10.6151
R1583 B.n416 B.n413 10.6151
R1584 B.n413 B.n412 10.6151
R1585 B.n412 B.n409 10.6151
R1586 B.n409 B.n408 10.6151
R1587 B.n408 B.n405 10.6151
R1588 B.n405 B.n404 10.6151
R1589 B.n404 B.n401 10.6151
R1590 B.n401 B.n368 10.6151
R1591 B.n508 B.n368 10.6151
R1592 B.n514 B.n364 10.6151
R1593 B.n515 B.n514 10.6151
R1594 B.n516 B.n515 10.6151
R1595 B.n516 B.n356 10.6151
R1596 B.n526 B.n356 10.6151
R1597 B.n527 B.n526 10.6151
R1598 B.n528 B.n527 10.6151
R1599 B.n528 B.n348 10.6151
R1600 B.n538 B.n348 10.6151
R1601 B.n539 B.n538 10.6151
R1602 B.n540 B.n539 10.6151
R1603 B.n540 B.n340 10.6151
R1604 B.n550 B.n340 10.6151
R1605 B.n551 B.n550 10.6151
R1606 B.n552 B.n551 10.6151
R1607 B.n552 B.n332 10.6151
R1608 B.n562 B.n332 10.6151
R1609 B.n563 B.n562 10.6151
R1610 B.n564 B.n563 10.6151
R1611 B.n564 B.n324 10.6151
R1612 B.n575 B.n324 10.6151
R1613 B.n576 B.n575 10.6151
R1614 B.n577 B.n576 10.6151
R1615 B.n577 B.n317 10.6151
R1616 B.n587 B.n317 10.6151
R1617 B.n588 B.n587 10.6151
R1618 B.n589 B.n588 10.6151
R1619 B.n589 B.n309 10.6151
R1620 B.n599 B.n309 10.6151
R1621 B.n600 B.n599 10.6151
R1622 B.n601 B.n600 10.6151
R1623 B.n601 B.n301 10.6151
R1624 B.n611 B.n301 10.6151
R1625 B.n612 B.n611 10.6151
R1626 B.n613 B.n612 10.6151
R1627 B.n613 B.n293 10.6151
R1628 B.n623 B.n293 10.6151
R1629 B.n624 B.n623 10.6151
R1630 B.n625 B.n624 10.6151
R1631 B.n625 B.n285 10.6151
R1632 B.n635 B.n285 10.6151
R1633 B.n636 B.n635 10.6151
R1634 B.n637 B.n636 10.6151
R1635 B.n637 B.n277 10.6151
R1636 B.n647 B.n277 10.6151
R1637 B.n648 B.n647 10.6151
R1638 B.n649 B.n648 10.6151
R1639 B.n649 B.n269 10.6151
R1640 B.n659 B.n269 10.6151
R1641 B.n660 B.n659 10.6151
R1642 B.n661 B.n660 10.6151
R1643 B.n661 B.n261 10.6151
R1644 B.n672 B.n261 10.6151
R1645 B.n673 B.n672 10.6151
R1646 B.n674 B.n673 10.6151
R1647 B.n674 B.n254 10.6151
R1648 B.n685 B.n254 10.6151
R1649 B.n686 B.n685 10.6151
R1650 B.n687 B.n686 10.6151
R1651 B.n687 B.n0 10.6151
R1652 B.n891 B.n1 10.6151
R1653 B.n891 B.n890 10.6151
R1654 B.n890 B.n889 10.6151
R1655 B.n889 B.n10 10.6151
R1656 B.n883 B.n10 10.6151
R1657 B.n883 B.n882 10.6151
R1658 B.n882 B.n881 10.6151
R1659 B.n881 B.n16 10.6151
R1660 B.n875 B.n16 10.6151
R1661 B.n875 B.n874 10.6151
R1662 B.n874 B.n873 10.6151
R1663 B.n873 B.n24 10.6151
R1664 B.n867 B.n24 10.6151
R1665 B.n867 B.n866 10.6151
R1666 B.n866 B.n865 10.6151
R1667 B.n865 B.n31 10.6151
R1668 B.n859 B.n31 10.6151
R1669 B.n859 B.n858 10.6151
R1670 B.n858 B.n857 10.6151
R1671 B.n857 B.n38 10.6151
R1672 B.n851 B.n38 10.6151
R1673 B.n851 B.n850 10.6151
R1674 B.n850 B.n849 10.6151
R1675 B.n849 B.n45 10.6151
R1676 B.n843 B.n45 10.6151
R1677 B.n843 B.n842 10.6151
R1678 B.n842 B.n841 10.6151
R1679 B.n841 B.n52 10.6151
R1680 B.n835 B.n52 10.6151
R1681 B.n835 B.n834 10.6151
R1682 B.n834 B.n833 10.6151
R1683 B.n833 B.n59 10.6151
R1684 B.n827 B.n59 10.6151
R1685 B.n827 B.n826 10.6151
R1686 B.n826 B.n825 10.6151
R1687 B.n825 B.n66 10.6151
R1688 B.n819 B.n66 10.6151
R1689 B.n819 B.n818 10.6151
R1690 B.n818 B.n817 10.6151
R1691 B.n817 B.n72 10.6151
R1692 B.n811 B.n72 10.6151
R1693 B.n811 B.n810 10.6151
R1694 B.n810 B.n809 10.6151
R1695 B.n809 B.n80 10.6151
R1696 B.n803 B.n80 10.6151
R1697 B.n803 B.n802 10.6151
R1698 B.n802 B.n801 10.6151
R1699 B.n801 B.n87 10.6151
R1700 B.n795 B.n87 10.6151
R1701 B.n795 B.n794 10.6151
R1702 B.n794 B.n793 10.6151
R1703 B.n793 B.n94 10.6151
R1704 B.n787 B.n94 10.6151
R1705 B.n787 B.n786 10.6151
R1706 B.n786 B.n785 10.6151
R1707 B.n785 B.n101 10.6151
R1708 B.n779 B.n101 10.6151
R1709 B.n779 B.n778 10.6151
R1710 B.n778 B.n777 10.6151
R1711 B.n777 B.n108 10.6151
R1712 B.n187 B.n144 9.36635
R1713 B.n210 B.n141 9.36635
R1714 B.n463 B.n462 9.36635
R1715 B.n441 B.n440 9.36635
R1716 B.n669 B.t3 7.18669
R1717 B.n18 B.t2 7.18669
R1718 B.n609 B.t5 5.13349
R1719 B.n839 B.t6 5.13349
R1720 B.n897 B.n0 2.81026
R1721 B.n897 B.n1 2.81026
R1722 B.n190 B.n144 1.24928
R1723 B.n207 B.n141 1.24928
R1724 B.n462 B.n461 1.24928
R1725 B.n442 B.n441 1.24928
R1726 VP.n24 VP.n23 161.3
R1727 VP.n25 VP.n20 161.3
R1728 VP.n27 VP.n26 161.3
R1729 VP.n28 VP.n19 161.3
R1730 VP.n30 VP.n29 161.3
R1731 VP.n31 VP.n18 161.3
R1732 VP.n33 VP.n32 161.3
R1733 VP.n35 VP.n34 161.3
R1734 VP.n36 VP.n16 161.3
R1735 VP.n38 VP.n37 161.3
R1736 VP.n39 VP.n15 161.3
R1737 VP.n41 VP.n40 161.3
R1738 VP.n42 VP.n14 161.3
R1739 VP.n44 VP.n43 161.3
R1740 VP.n79 VP.n78 161.3
R1741 VP.n77 VP.n1 161.3
R1742 VP.n76 VP.n75 161.3
R1743 VP.n74 VP.n2 161.3
R1744 VP.n73 VP.n72 161.3
R1745 VP.n71 VP.n3 161.3
R1746 VP.n70 VP.n69 161.3
R1747 VP.n68 VP.n67 161.3
R1748 VP.n66 VP.n5 161.3
R1749 VP.n65 VP.n64 161.3
R1750 VP.n63 VP.n6 161.3
R1751 VP.n62 VP.n61 161.3
R1752 VP.n60 VP.n7 161.3
R1753 VP.n59 VP.n58 161.3
R1754 VP.n57 VP.n56 161.3
R1755 VP.n55 VP.n9 161.3
R1756 VP.n54 VP.n53 161.3
R1757 VP.n52 VP.n10 161.3
R1758 VP.n51 VP.n50 161.3
R1759 VP.n49 VP.n11 161.3
R1760 VP.n48 VP.n47 161.3
R1761 VP.n22 VP.t2 73.5142
R1762 VP.n46 VP.n12 70.5721
R1763 VP.n80 VP.n0 70.5721
R1764 VP.n45 VP.n13 70.5721
R1765 VP.n22 VP.n21 59.6505
R1766 VP.n50 VP.n10 50.2647
R1767 VP.n76 VP.n2 50.2647
R1768 VP.n41 VP.n15 50.2647
R1769 VP.n46 VP.n45 49.242
R1770 VP.n61 VP.n6 40.577
R1771 VP.n65 VP.n6 40.577
R1772 VP.n30 VP.n19 40.577
R1773 VP.n26 VP.n19 40.577
R1774 VP.n12 VP.t1 40.0935
R1775 VP.n8 VP.t0 40.0935
R1776 VP.n4 VP.t4 40.0935
R1777 VP.n0 VP.t5 40.0935
R1778 VP.n13 VP.t3 40.0935
R1779 VP.n17 VP.t7 40.0935
R1780 VP.n21 VP.t6 40.0935
R1781 VP.n54 VP.n10 30.8893
R1782 VP.n72 VP.n2 30.8893
R1783 VP.n37 VP.n15 30.8893
R1784 VP.n49 VP.n48 24.5923
R1785 VP.n50 VP.n49 24.5923
R1786 VP.n55 VP.n54 24.5923
R1787 VP.n56 VP.n55 24.5923
R1788 VP.n60 VP.n59 24.5923
R1789 VP.n61 VP.n60 24.5923
R1790 VP.n66 VP.n65 24.5923
R1791 VP.n67 VP.n66 24.5923
R1792 VP.n71 VP.n70 24.5923
R1793 VP.n72 VP.n71 24.5923
R1794 VP.n77 VP.n76 24.5923
R1795 VP.n78 VP.n77 24.5923
R1796 VP.n42 VP.n41 24.5923
R1797 VP.n43 VP.n42 24.5923
R1798 VP.n31 VP.n30 24.5923
R1799 VP.n32 VP.n31 24.5923
R1800 VP.n36 VP.n35 24.5923
R1801 VP.n37 VP.n36 24.5923
R1802 VP.n25 VP.n24 24.5923
R1803 VP.n26 VP.n25 24.5923
R1804 VP.n48 VP.n12 19.674
R1805 VP.n78 VP.n0 19.674
R1806 VP.n43 VP.n13 19.674
R1807 VP.n59 VP.n8 14.7556
R1808 VP.n67 VP.n4 14.7556
R1809 VP.n32 VP.n17 14.7556
R1810 VP.n24 VP.n21 14.7556
R1811 VP.n56 VP.n8 9.83723
R1812 VP.n70 VP.n4 9.83723
R1813 VP.n35 VP.n17 9.83723
R1814 VP.n23 VP.n22 3.91112
R1815 VP.n45 VP.n44 0.354861
R1816 VP.n47 VP.n46 0.354861
R1817 VP.n80 VP.n79 0.354861
R1818 VP VP.n80 0.267071
R1819 VP.n23 VP.n20 0.189894
R1820 VP.n27 VP.n20 0.189894
R1821 VP.n28 VP.n27 0.189894
R1822 VP.n29 VP.n28 0.189894
R1823 VP.n29 VP.n18 0.189894
R1824 VP.n33 VP.n18 0.189894
R1825 VP.n34 VP.n33 0.189894
R1826 VP.n34 VP.n16 0.189894
R1827 VP.n38 VP.n16 0.189894
R1828 VP.n39 VP.n38 0.189894
R1829 VP.n40 VP.n39 0.189894
R1830 VP.n40 VP.n14 0.189894
R1831 VP.n44 VP.n14 0.189894
R1832 VP.n47 VP.n11 0.189894
R1833 VP.n51 VP.n11 0.189894
R1834 VP.n52 VP.n51 0.189894
R1835 VP.n53 VP.n52 0.189894
R1836 VP.n53 VP.n9 0.189894
R1837 VP.n57 VP.n9 0.189894
R1838 VP.n58 VP.n57 0.189894
R1839 VP.n58 VP.n7 0.189894
R1840 VP.n62 VP.n7 0.189894
R1841 VP.n63 VP.n62 0.189894
R1842 VP.n64 VP.n63 0.189894
R1843 VP.n64 VP.n5 0.189894
R1844 VP.n68 VP.n5 0.189894
R1845 VP.n69 VP.n68 0.189894
R1846 VP.n69 VP.n3 0.189894
R1847 VP.n73 VP.n3 0.189894
R1848 VP.n74 VP.n73 0.189894
R1849 VP.n75 VP.n74 0.189894
R1850 VP.n75 VP.n1 0.189894
R1851 VP.n79 VP.n1 0.189894
R1852 VDD1 VDD1.n0 71.6797
R1853 VDD1.n3 VDD1.n2 71.566
R1854 VDD1.n3 VDD1.n1 71.566
R1855 VDD1.n5 VDD1.n4 70.0689
R1856 VDD1.n5 VDD1.n3 42.9535
R1857 VDD1.n4 VDD1.t0 3.64021
R1858 VDD1.n4 VDD1.t4 3.64021
R1859 VDD1.n0 VDD1.t5 3.64021
R1860 VDD1.n0 VDD1.t1 3.64021
R1861 VDD1.n2 VDD1.t3 3.64021
R1862 VDD1.n2 VDD1.t2 3.64021
R1863 VDD1.n1 VDD1.t6 3.64021
R1864 VDD1.n1 VDD1.t7 3.64021
R1865 VDD1 VDD1.n5 1.49403
C0 VDD1 VDD2 2.12564f
C1 VP VTAIL 5.52441f
C2 VP VN 7.25852f
C3 VN VTAIL 5.5103f
C4 VDD1 VP 4.79945f
C5 VDD1 VTAIL 6.35366f
C6 VP VDD2 0.59507f
C7 VDD2 VTAIL 6.41256f
C8 VDD1 VN 0.153154f
C9 VDD2 VN 4.3632f
C10 VDD2 B 5.605489f
C11 VDD1 B 6.129807f
C12 VTAIL B 6.518911f
C13 VN B 17.43302f
C14 VP B 16.046871f
C15 VDD1.t5 B 0.126779f
C16 VDD1.t1 B 0.126779f
C17 VDD1.n0 B 1.07234f
C18 VDD1.t6 B 0.126779f
C19 VDD1.t7 B 0.126779f
C20 VDD1.n1 B 1.07106f
C21 VDD1.t3 B 0.126779f
C22 VDD1.t2 B 0.126779f
C23 VDD1.n2 B 1.07106f
C24 VDD1.n3 B 3.87274f
C25 VDD1.t0 B 0.126779f
C26 VDD1.t4 B 0.126779f
C27 VDD1.n4 B 1.05697f
C28 VDD1.n5 B 3.17789f
C29 VP.t5 B 1.0765f
C30 VP.n0 B 0.500092f
C31 VP.n1 B 0.023003f
C32 VP.n2 B 0.021689f
C33 VP.n3 B 0.023003f
C34 VP.t4 B 1.0765f
C35 VP.n4 B 0.403314f
C36 VP.n5 B 0.023003f
C37 VP.n6 B 0.018579f
C38 VP.n7 B 0.023003f
C39 VP.t0 B 1.0765f
C40 VP.n8 B 0.403314f
C41 VP.n9 B 0.023003f
C42 VP.n10 B 0.021689f
C43 VP.n11 B 0.023003f
C44 VP.t1 B 1.0765f
C45 VP.n12 B 0.500092f
C46 VP.t3 B 1.0765f
C47 VP.n13 B 0.500092f
C48 VP.n14 B 0.023003f
C49 VP.n15 B 0.021689f
C50 VP.n16 B 0.023003f
C51 VP.t7 B 1.0765f
C52 VP.n17 B 0.403314f
C53 VP.n18 B 0.023003f
C54 VP.n19 B 0.018579f
C55 VP.n20 B 0.023003f
C56 VP.t6 B 1.0765f
C57 VP.n21 B 0.481222f
C58 VP.t2 B 1.33606f
C59 VP.n22 B 0.458548f
C60 VP.n23 B 0.266867f
C61 VP.n24 B 0.034234f
C62 VP.n25 B 0.042657f
C63 VP.n26 B 0.045478f
C64 VP.n27 B 0.023003f
C65 VP.n28 B 0.023003f
C66 VP.n29 B 0.023003f
C67 VP.n30 B 0.045478f
C68 VP.n31 B 0.042657f
C69 VP.n32 B 0.034234f
C70 VP.n33 B 0.023003f
C71 VP.n34 B 0.023003f
C72 VP.n35 B 0.030022f
C73 VP.n36 B 0.042657f
C74 VP.n37 B 0.045834f
C75 VP.n38 B 0.023003f
C76 VP.n39 B 0.023003f
C77 VP.n40 B 0.023003f
C78 VP.n41 B 0.042012f
C79 VP.n42 B 0.042657f
C80 VP.n43 B 0.038445f
C81 VP.n44 B 0.037121f
C82 VP.n45 B 1.27619f
C83 VP.n46 B 1.29303f
C84 VP.n47 B 0.037121f
C85 VP.n48 B 0.038445f
C86 VP.n49 B 0.042657f
C87 VP.n50 B 0.042012f
C88 VP.n51 B 0.023003f
C89 VP.n52 B 0.023003f
C90 VP.n53 B 0.023003f
C91 VP.n54 B 0.045834f
C92 VP.n55 B 0.042657f
C93 VP.n56 B 0.030022f
C94 VP.n57 B 0.023003f
C95 VP.n58 B 0.023003f
C96 VP.n59 B 0.034234f
C97 VP.n60 B 0.042657f
C98 VP.n61 B 0.045478f
C99 VP.n62 B 0.023003f
C100 VP.n63 B 0.023003f
C101 VP.n64 B 0.023003f
C102 VP.n65 B 0.045478f
C103 VP.n66 B 0.042657f
C104 VP.n67 B 0.034234f
C105 VP.n68 B 0.023003f
C106 VP.n69 B 0.023003f
C107 VP.n70 B 0.030022f
C108 VP.n71 B 0.042657f
C109 VP.n72 B 0.045834f
C110 VP.n73 B 0.023003f
C111 VP.n74 B 0.023003f
C112 VP.n75 B 0.023003f
C113 VP.n76 B 0.042012f
C114 VP.n77 B 0.042657f
C115 VP.n78 B 0.038445f
C116 VP.n79 B 0.037121f
C117 VP.n80 B 0.050358f
C118 VTAIL.t8 B 0.107235f
C119 VTAIL.t11 B 0.107235f
C120 VTAIL.n0 B 0.83623f
C121 VTAIL.n1 B 0.467828f
C122 VTAIL.t10 B 1.0635f
C123 VTAIL.n2 B 0.566102f
C124 VTAIL.t3 B 1.0635f
C125 VTAIL.n3 B 0.566102f
C126 VTAIL.t5 B 0.107235f
C127 VTAIL.t1 B 0.107235f
C128 VTAIL.n4 B 0.83623f
C129 VTAIL.n5 B 0.712603f
C130 VTAIL.t7 B 1.0635f
C131 VTAIL.n6 B 1.49359f
C132 VTAIL.t9 B 1.0635f
C133 VTAIL.n7 B 1.49359f
C134 VTAIL.t14 B 0.107235f
C135 VTAIL.t15 B 0.107235f
C136 VTAIL.n8 B 0.836234f
C137 VTAIL.n9 B 0.712599f
C138 VTAIL.t12 B 1.0635f
C139 VTAIL.n10 B 0.566101f
C140 VTAIL.t2 B 1.0635f
C141 VTAIL.n11 B 0.566101f
C142 VTAIL.t4 B 0.107235f
C143 VTAIL.t6 B 0.107235f
C144 VTAIL.n12 B 0.836234f
C145 VTAIL.n13 B 0.712599f
C146 VTAIL.t0 B 1.0635f
C147 VTAIL.n14 B 1.49359f
C148 VTAIL.t13 B 1.0635f
C149 VTAIL.n15 B 1.48891f
C150 VDD2.t4 B 0.123981f
C151 VDD2.t5 B 0.123981f
C152 VDD2.n0 B 1.04743f
C153 VDD2.t3 B 0.123981f
C154 VDD2.t0 B 0.123981f
C155 VDD2.n1 B 1.04743f
C156 VDD2.n2 B 3.72742f
C157 VDD2.t2 B 0.123981f
C158 VDD2.t6 B 0.123981f
C159 VDD2.n3 B 1.03365f
C160 VDD2.n4 B 3.07191f
C161 VDD2.t1 B 0.123981f
C162 VDD2.t7 B 0.123981f
C163 VDD2.n5 B 1.04739f
C164 VN.t2 B 1.0501f
C165 VN.n0 B 0.48783f
C166 VN.n1 B 0.022439f
C167 VN.n2 B 0.021157f
C168 VN.n3 B 0.022439f
C169 VN.t4 B 1.0501f
C170 VN.n4 B 0.393425f
C171 VN.n5 B 0.022439f
C172 VN.n6 B 0.018123f
C173 VN.n7 B 0.022439f
C174 VN.t7 B 1.0501f
C175 VN.n8 B 0.469423f
C176 VN.t5 B 1.3033f
C177 VN.n9 B 0.447304f
C178 VN.n10 B 0.260323f
C179 VN.n11 B 0.033394f
C180 VN.n12 B 0.041611f
C181 VN.n13 B 0.044363f
C182 VN.n14 B 0.022439f
C183 VN.n15 B 0.022439f
C184 VN.n16 B 0.022439f
C185 VN.n17 B 0.044363f
C186 VN.n18 B 0.041611f
C187 VN.n19 B 0.033394f
C188 VN.n20 B 0.022439f
C189 VN.n21 B 0.022439f
C190 VN.n22 B 0.029286f
C191 VN.n23 B 0.041611f
C192 VN.n24 B 0.04471f
C193 VN.n25 B 0.022439f
C194 VN.n26 B 0.022439f
C195 VN.n27 B 0.022439f
C196 VN.n28 B 0.040982f
C197 VN.n29 B 0.041611f
C198 VN.n30 B 0.037503f
C199 VN.n31 B 0.036211f
C200 VN.n32 B 0.049123f
C201 VN.t6 B 1.0501f
C202 VN.n33 B 0.48783f
C203 VN.n34 B 0.022439f
C204 VN.n35 B 0.021157f
C205 VN.n36 B 0.022439f
C206 VN.t1 B 1.0501f
C207 VN.n37 B 0.393425f
C208 VN.n38 B 0.022439f
C209 VN.n39 B 0.018123f
C210 VN.n40 B 0.022439f
C211 VN.t0 B 1.0501f
C212 VN.n41 B 0.469423f
C213 VN.t3 B 1.3033f
C214 VN.n42 B 0.447304f
C215 VN.n43 B 0.260323f
C216 VN.n44 B 0.033394f
C217 VN.n45 B 0.041611f
C218 VN.n46 B 0.044363f
C219 VN.n47 B 0.022439f
C220 VN.n48 B 0.022439f
C221 VN.n49 B 0.022439f
C222 VN.n50 B 0.044363f
C223 VN.n51 B 0.041611f
C224 VN.n52 B 0.033394f
C225 VN.n53 B 0.022439f
C226 VN.n54 B 0.022439f
C227 VN.n55 B 0.029286f
C228 VN.n56 B 0.041611f
C229 VN.n57 B 0.04471f
C230 VN.n58 B 0.022439f
C231 VN.n59 B 0.022439f
C232 VN.n60 B 0.022439f
C233 VN.n61 B 0.040982f
C234 VN.n62 B 0.041611f
C235 VN.n63 B 0.037503f
C236 VN.n64 B 0.036211f
C237 VN.n65 B 1.25411f
.ends

