* NGSPICE file created from diff_pair_sample_0706.ext - technology: sky130A

.subckt diff_pair_sample_0706 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 w_n1382_n4218# sky130_fd_pr__pfet_01v8 ad=6.3297 pd=33.24 as=6.3297 ps=33.24 w=16.23 l=0.7
X1 B.t11 B.t9 B.t10 w_n1382_n4218# sky130_fd_pr__pfet_01v8 ad=6.3297 pd=33.24 as=0 ps=0 w=16.23 l=0.7
X2 VDD1.t0 VP.t1 VTAIL.t1 w_n1382_n4218# sky130_fd_pr__pfet_01v8 ad=6.3297 pd=33.24 as=6.3297 ps=33.24 w=16.23 l=0.7
X3 B.t8 B.t6 B.t7 w_n1382_n4218# sky130_fd_pr__pfet_01v8 ad=6.3297 pd=33.24 as=0 ps=0 w=16.23 l=0.7
X4 VDD2.t1 VN.t0 VTAIL.t0 w_n1382_n4218# sky130_fd_pr__pfet_01v8 ad=6.3297 pd=33.24 as=6.3297 ps=33.24 w=16.23 l=0.7
X5 VDD2.t0 VN.t1 VTAIL.t3 w_n1382_n4218# sky130_fd_pr__pfet_01v8 ad=6.3297 pd=33.24 as=6.3297 ps=33.24 w=16.23 l=0.7
X6 B.t5 B.t3 B.t4 w_n1382_n4218# sky130_fd_pr__pfet_01v8 ad=6.3297 pd=33.24 as=0 ps=0 w=16.23 l=0.7
X7 B.t2 B.t0 B.t1 w_n1382_n4218# sky130_fd_pr__pfet_01v8 ad=6.3297 pd=33.24 as=0 ps=0 w=16.23 l=0.7
R0 VP.n0 VP.t0 819.376
R1 VP.n0 VP.t1 776.539
R2 VP VP.n0 0.0516364
R3 VTAIL.n354 VTAIL.n270 756.745
R4 VTAIL.n84 VTAIL.n0 756.745
R5 VTAIL.n264 VTAIL.n180 756.745
R6 VTAIL.n174 VTAIL.n90 756.745
R7 VTAIL.n298 VTAIL.n297 585
R8 VTAIL.n303 VTAIL.n302 585
R9 VTAIL.n305 VTAIL.n304 585
R10 VTAIL.n294 VTAIL.n293 585
R11 VTAIL.n311 VTAIL.n310 585
R12 VTAIL.n313 VTAIL.n312 585
R13 VTAIL.n290 VTAIL.n289 585
R14 VTAIL.n319 VTAIL.n318 585
R15 VTAIL.n321 VTAIL.n320 585
R16 VTAIL.n286 VTAIL.n285 585
R17 VTAIL.n327 VTAIL.n326 585
R18 VTAIL.n329 VTAIL.n328 585
R19 VTAIL.n282 VTAIL.n281 585
R20 VTAIL.n335 VTAIL.n334 585
R21 VTAIL.n337 VTAIL.n336 585
R22 VTAIL.n278 VTAIL.n277 585
R23 VTAIL.n344 VTAIL.n343 585
R24 VTAIL.n345 VTAIL.n276 585
R25 VTAIL.n347 VTAIL.n346 585
R26 VTAIL.n274 VTAIL.n273 585
R27 VTAIL.n353 VTAIL.n352 585
R28 VTAIL.n355 VTAIL.n354 585
R29 VTAIL.n28 VTAIL.n27 585
R30 VTAIL.n33 VTAIL.n32 585
R31 VTAIL.n35 VTAIL.n34 585
R32 VTAIL.n24 VTAIL.n23 585
R33 VTAIL.n41 VTAIL.n40 585
R34 VTAIL.n43 VTAIL.n42 585
R35 VTAIL.n20 VTAIL.n19 585
R36 VTAIL.n49 VTAIL.n48 585
R37 VTAIL.n51 VTAIL.n50 585
R38 VTAIL.n16 VTAIL.n15 585
R39 VTAIL.n57 VTAIL.n56 585
R40 VTAIL.n59 VTAIL.n58 585
R41 VTAIL.n12 VTAIL.n11 585
R42 VTAIL.n65 VTAIL.n64 585
R43 VTAIL.n67 VTAIL.n66 585
R44 VTAIL.n8 VTAIL.n7 585
R45 VTAIL.n74 VTAIL.n73 585
R46 VTAIL.n75 VTAIL.n6 585
R47 VTAIL.n77 VTAIL.n76 585
R48 VTAIL.n4 VTAIL.n3 585
R49 VTAIL.n83 VTAIL.n82 585
R50 VTAIL.n85 VTAIL.n84 585
R51 VTAIL.n265 VTAIL.n264 585
R52 VTAIL.n263 VTAIL.n262 585
R53 VTAIL.n184 VTAIL.n183 585
R54 VTAIL.n257 VTAIL.n256 585
R55 VTAIL.n255 VTAIL.n186 585
R56 VTAIL.n254 VTAIL.n253 585
R57 VTAIL.n189 VTAIL.n187 585
R58 VTAIL.n248 VTAIL.n247 585
R59 VTAIL.n246 VTAIL.n245 585
R60 VTAIL.n193 VTAIL.n192 585
R61 VTAIL.n240 VTAIL.n239 585
R62 VTAIL.n238 VTAIL.n237 585
R63 VTAIL.n197 VTAIL.n196 585
R64 VTAIL.n232 VTAIL.n231 585
R65 VTAIL.n230 VTAIL.n229 585
R66 VTAIL.n201 VTAIL.n200 585
R67 VTAIL.n224 VTAIL.n223 585
R68 VTAIL.n222 VTAIL.n221 585
R69 VTAIL.n205 VTAIL.n204 585
R70 VTAIL.n216 VTAIL.n215 585
R71 VTAIL.n214 VTAIL.n213 585
R72 VTAIL.n209 VTAIL.n208 585
R73 VTAIL.n175 VTAIL.n174 585
R74 VTAIL.n173 VTAIL.n172 585
R75 VTAIL.n94 VTAIL.n93 585
R76 VTAIL.n167 VTAIL.n166 585
R77 VTAIL.n165 VTAIL.n96 585
R78 VTAIL.n164 VTAIL.n163 585
R79 VTAIL.n99 VTAIL.n97 585
R80 VTAIL.n158 VTAIL.n157 585
R81 VTAIL.n156 VTAIL.n155 585
R82 VTAIL.n103 VTAIL.n102 585
R83 VTAIL.n150 VTAIL.n149 585
R84 VTAIL.n148 VTAIL.n147 585
R85 VTAIL.n107 VTAIL.n106 585
R86 VTAIL.n142 VTAIL.n141 585
R87 VTAIL.n140 VTAIL.n139 585
R88 VTAIL.n111 VTAIL.n110 585
R89 VTAIL.n134 VTAIL.n133 585
R90 VTAIL.n132 VTAIL.n131 585
R91 VTAIL.n115 VTAIL.n114 585
R92 VTAIL.n126 VTAIL.n125 585
R93 VTAIL.n124 VTAIL.n123 585
R94 VTAIL.n119 VTAIL.n118 585
R95 VTAIL.n299 VTAIL.t0 327.466
R96 VTAIL.n29 VTAIL.t1 327.466
R97 VTAIL.n210 VTAIL.t2 327.466
R98 VTAIL.n120 VTAIL.t3 327.466
R99 VTAIL.n303 VTAIL.n297 171.744
R100 VTAIL.n304 VTAIL.n303 171.744
R101 VTAIL.n304 VTAIL.n293 171.744
R102 VTAIL.n311 VTAIL.n293 171.744
R103 VTAIL.n312 VTAIL.n311 171.744
R104 VTAIL.n312 VTAIL.n289 171.744
R105 VTAIL.n319 VTAIL.n289 171.744
R106 VTAIL.n320 VTAIL.n319 171.744
R107 VTAIL.n320 VTAIL.n285 171.744
R108 VTAIL.n327 VTAIL.n285 171.744
R109 VTAIL.n328 VTAIL.n327 171.744
R110 VTAIL.n328 VTAIL.n281 171.744
R111 VTAIL.n335 VTAIL.n281 171.744
R112 VTAIL.n336 VTAIL.n335 171.744
R113 VTAIL.n336 VTAIL.n277 171.744
R114 VTAIL.n344 VTAIL.n277 171.744
R115 VTAIL.n345 VTAIL.n344 171.744
R116 VTAIL.n346 VTAIL.n345 171.744
R117 VTAIL.n346 VTAIL.n273 171.744
R118 VTAIL.n353 VTAIL.n273 171.744
R119 VTAIL.n354 VTAIL.n353 171.744
R120 VTAIL.n33 VTAIL.n27 171.744
R121 VTAIL.n34 VTAIL.n33 171.744
R122 VTAIL.n34 VTAIL.n23 171.744
R123 VTAIL.n41 VTAIL.n23 171.744
R124 VTAIL.n42 VTAIL.n41 171.744
R125 VTAIL.n42 VTAIL.n19 171.744
R126 VTAIL.n49 VTAIL.n19 171.744
R127 VTAIL.n50 VTAIL.n49 171.744
R128 VTAIL.n50 VTAIL.n15 171.744
R129 VTAIL.n57 VTAIL.n15 171.744
R130 VTAIL.n58 VTAIL.n57 171.744
R131 VTAIL.n58 VTAIL.n11 171.744
R132 VTAIL.n65 VTAIL.n11 171.744
R133 VTAIL.n66 VTAIL.n65 171.744
R134 VTAIL.n66 VTAIL.n7 171.744
R135 VTAIL.n74 VTAIL.n7 171.744
R136 VTAIL.n75 VTAIL.n74 171.744
R137 VTAIL.n76 VTAIL.n75 171.744
R138 VTAIL.n76 VTAIL.n3 171.744
R139 VTAIL.n83 VTAIL.n3 171.744
R140 VTAIL.n84 VTAIL.n83 171.744
R141 VTAIL.n264 VTAIL.n263 171.744
R142 VTAIL.n263 VTAIL.n183 171.744
R143 VTAIL.n256 VTAIL.n183 171.744
R144 VTAIL.n256 VTAIL.n255 171.744
R145 VTAIL.n255 VTAIL.n254 171.744
R146 VTAIL.n254 VTAIL.n187 171.744
R147 VTAIL.n247 VTAIL.n187 171.744
R148 VTAIL.n247 VTAIL.n246 171.744
R149 VTAIL.n246 VTAIL.n192 171.744
R150 VTAIL.n239 VTAIL.n192 171.744
R151 VTAIL.n239 VTAIL.n238 171.744
R152 VTAIL.n238 VTAIL.n196 171.744
R153 VTAIL.n231 VTAIL.n196 171.744
R154 VTAIL.n231 VTAIL.n230 171.744
R155 VTAIL.n230 VTAIL.n200 171.744
R156 VTAIL.n223 VTAIL.n200 171.744
R157 VTAIL.n223 VTAIL.n222 171.744
R158 VTAIL.n222 VTAIL.n204 171.744
R159 VTAIL.n215 VTAIL.n204 171.744
R160 VTAIL.n215 VTAIL.n214 171.744
R161 VTAIL.n214 VTAIL.n208 171.744
R162 VTAIL.n174 VTAIL.n173 171.744
R163 VTAIL.n173 VTAIL.n93 171.744
R164 VTAIL.n166 VTAIL.n93 171.744
R165 VTAIL.n166 VTAIL.n165 171.744
R166 VTAIL.n165 VTAIL.n164 171.744
R167 VTAIL.n164 VTAIL.n97 171.744
R168 VTAIL.n157 VTAIL.n97 171.744
R169 VTAIL.n157 VTAIL.n156 171.744
R170 VTAIL.n156 VTAIL.n102 171.744
R171 VTAIL.n149 VTAIL.n102 171.744
R172 VTAIL.n149 VTAIL.n148 171.744
R173 VTAIL.n148 VTAIL.n106 171.744
R174 VTAIL.n141 VTAIL.n106 171.744
R175 VTAIL.n141 VTAIL.n140 171.744
R176 VTAIL.n140 VTAIL.n110 171.744
R177 VTAIL.n133 VTAIL.n110 171.744
R178 VTAIL.n133 VTAIL.n132 171.744
R179 VTAIL.n132 VTAIL.n114 171.744
R180 VTAIL.n125 VTAIL.n114 171.744
R181 VTAIL.n125 VTAIL.n124 171.744
R182 VTAIL.n124 VTAIL.n118 171.744
R183 VTAIL.t0 VTAIL.n297 85.8723
R184 VTAIL.t1 VTAIL.n27 85.8723
R185 VTAIL.t2 VTAIL.n208 85.8723
R186 VTAIL.t3 VTAIL.n118 85.8723
R187 VTAIL.n359 VTAIL.n358 35.0944
R188 VTAIL.n89 VTAIL.n88 35.0944
R189 VTAIL.n269 VTAIL.n268 35.0944
R190 VTAIL.n179 VTAIL.n178 35.0944
R191 VTAIL.n179 VTAIL.n89 28.1514
R192 VTAIL.n359 VTAIL.n269 27.2634
R193 VTAIL.n299 VTAIL.n298 16.3895
R194 VTAIL.n29 VTAIL.n28 16.3895
R195 VTAIL.n210 VTAIL.n209 16.3895
R196 VTAIL.n120 VTAIL.n119 16.3895
R197 VTAIL.n347 VTAIL.n276 13.1884
R198 VTAIL.n77 VTAIL.n6 13.1884
R199 VTAIL.n257 VTAIL.n186 13.1884
R200 VTAIL.n167 VTAIL.n96 13.1884
R201 VTAIL.n302 VTAIL.n301 12.8005
R202 VTAIL.n343 VTAIL.n342 12.8005
R203 VTAIL.n348 VTAIL.n274 12.8005
R204 VTAIL.n32 VTAIL.n31 12.8005
R205 VTAIL.n73 VTAIL.n72 12.8005
R206 VTAIL.n78 VTAIL.n4 12.8005
R207 VTAIL.n258 VTAIL.n184 12.8005
R208 VTAIL.n253 VTAIL.n188 12.8005
R209 VTAIL.n213 VTAIL.n212 12.8005
R210 VTAIL.n168 VTAIL.n94 12.8005
R211 VTAIL.n163 VTAIL.n98 12.8005
R212 VTAIL.n123 VTAIL.n122 12.8005
R213 VTAIL.n305 VTAIL.n296 12.0247
R214 VTAIL.n341 VTAIL.n278 12.0247
R215 VTAIL.n352 VTAIL.n351 12.0247
R216 VTAIL.n35 VTAIL.n26 12.0247
R217 VTAIL.n71 VTAIL.n8 12.0247
R218 VTAIL.n82 VTAIL.n81 12.0247
R219 VTAIL.n262 VTAIL.n261 12.0247
R220 VTAIL.n252 VTAIL.n189 12.0247
R221 VTAIL.n216 VTAIL.n207 12.0247
R222 VTAIL.n172 VTAIL.n171 12.0247
R223 VTAIL.n162 VTAIL.n99 12.0247
R224 VTAIL.n126 VTAIL.n117 12.0247
R225 VTAIL.n306 VTAIL.n294 11.249
R226 VTAIL.n338 VTAIL.n337 11.249
R227 VTAIL.n355 VTAIL.n272 11.249
R228 VTAIL.n36 VTAIL.n24 11.249
R229 VTAIL.n68 VTAIL.n67 11.249
R230 VTAIL.n85 VTAIL.n2 11.249
R231 VTAIL.n265 VTAIL.n182 11.249
R232 VTAIL.n249 VTAIL.n248 11.249
R233 VTAIL.n217 VTAIL.n205 11.249
R234 VTAIL.n175 VTAIL.n92 11.249
R235 VTAIL.n159 VTAIL.n158 11.249
R236 VTAIL.n127 VTAIL.n115 11.249
R237 VTAIL.n310 VTAIL.n309 10.4732
R238 VTAIL.n334 VTAIL.n280 10.4732
R239 VTAIL.n356 VTAIL.n270 10.4732
R240 VTAIL.n40 VTAIL.n39 10.4732
R241 VTAIL.n64 VTAIL.n10 10.4732
R242 VTAIL.n86 VTAIL.n0 10.4732
R243 VTAIL.n266 VTAIL.n180 10.4732
R244 VTAIL.n245 VTAIL.n191 10.4732
R245 VTAIL.n221 VTAIL.n220 10.4732
R246 VTAIL.n176 VTAIL.n90 10.4732
R247 VTAIL.n155 VTAIL.n101 10.4732
R248 VTAIL.n131 VTAIL.n130 10.4732
R249 VTAIL.n313 VTAIL.n292 9.69747
R250 VTAIL.n333 VTAIL.n282 9.69747
R251 VTAIL.n43 VTAIL.n22 9.69747
R252 VTAIL.n63 VTAIL.n12 9.69747
R253 VTAIL.n244 VTAIL.n193 9.69747
R254 VTAIL.n224 VTAIL.n203 9.69747
R255 VTAIL.n154 VTAIL.n103 9.69747
R256 VTAIL.n134 VTAIL.n113 9.69747
R257 VTAIL.n358 VTAIL.n357 9.45567
R258 VTAIL.n88 VTAIL.n87 9.45567
R259 VTAIL.n268 VTAIL.n267 9.45567
R260 VTAIL.n178 VTAIL.n177 9.45567
R261 VTAIL.n357 VTAIL.n356 9.3005
R262 VTAIL.n272 VTAIL.n271 9.3005
R263 VTAIL.n351 VTAIL.n350 9.3005
R264 VTAIL.n349 VTAIL.n348 9.3005
R265 VTAIL.n288 VTAIL.n287 9.3005
R266 VTAIL.n317 VTAIL.n316 9.3005
R267 VTAIL.n315 VTAIL.n314 9.3005
R268 VTAIL.n292 VTAIL.n291 9.3005
R269 VTAIL.n309 VTAIL.n308 9.3005
R270 VTAIL.n307 VTAIL.n306 9.3005
R271 VTAIL.n296 VTAIL.n295 9.3005
R272 VTAIL.n301 VTAIL.n300 9.3005
R273 VTAIL.n323 VTAIL.n322 9.3005
R274 VTAIL.n325 VTAIL.n324 9.3005
R275 VTAIL.n284 VTAIL.n283 9.3005
R276 VTAIL.n331 VTAIL.n330 9.3005
R277 VTAIL.n333 VTAIL.n332 9.3005
R278 VTAIL.n280 VTAIL.n279 9.3005
R279 VTAIL.n339 VTAIL.n338 9.3005
R280 VTAIL.n341 VTAIL.n340 9.3005
R281 VTAIL.n342 VTAIL.n275 9.3005
R282 VTAIL.n87 VTAIL.n86 9.3005
R283 VTAIL.n2 VTAIL.n1 9.3005
R284 VTAIL.n81 VTAIL.n80 9.3005
R285 VTAIL.n79 VTAIL.n78 9.3005
R286 VTAIL.n18 VTAIL.n17 9.3005
R287 VTAIL.n47 VTAIL.n46 9.3005
R288 VTAIL.n45 VTAIL.n44 9.3005
R289 VTAIL.n22 VTAIL.n21 9.3005
R290 VTAIL.n39 VTAIL.n38 9.3005
R291 VTAIL.n37 VTAIL.n36 9.3005
R292 VTAIL.n26 VTAIL.n25 9.3005
R293 VTAIL.n31 VTAIL.n30 9.3005
R294 VTAIL.n53 VTAIL.n52 9.3005
R295 VTAIL.n55 VTAIL.n54 9.3005
R296 VTAIL.n14 VTAIL.n13 9.3005
R297 VTAIL.n61 VTAIL.n60 9.3005
R298 VTAIL.n63 VTAIL.n62 9.3005
R299 VTAIL.n10 VTAIL.n9 9.3005
R300 VTAIL.n69 VTAIL.n68 9.3005
R301 VTAIL.n71 VTAIL.n70 9.3005
R302 VTAIL.n72 VTAIL.n5 9.3005
R303 VTAIL.n236 VTAIL.n235 9.3005
R304 VTAIL.n195 VTAIL.n194 9.3005
R305 VTAIL.n242 VTAIL.n241 9.3005
R306 VTAIL.n244 VTAIL.n243 9.3005
R307 VTAIL.n191 VTAIL.n190 9.3005
R308 VTAIL.n250 VTAIL.n249 9.3005
R309 VTAIL.n252 VTAIL.n251 9.3005
R310 VTAIL.n188 VTAIL.n185 9.3005
R311 VTAIL.n267 VTAIL.n266 9.3005
R312 VTAIL.n182 VTAIL.n181 9.3005
R313 VTAIL.n261 VTAIL.n260 9.3005
R314 VTAIL.n259 VTAIL.n258 9.3005
R315 VTAIL.n234 VTAIL.n233 9.3005
R316 VTAIL.n199 VTAIL.n198 9.3005
R317 VTAIL.n228 VTAIL.n227 9.3005
R318 VTAIL.n226 VTAIL.n225 9.3005
R319 VTAIL.n203 VTAIL.n202 9.3005
R320 VTAIL.n220 VTAIL.n219 9.3005
R321 VTAIL.n218 VTAIL.n217 9.3005
R322 VTAIL.n207 VTAIL.n206 9.3005
R323 VTAIL.n212 VTAIL.n211 9.3005
R324 VTAIL.n146 VTAIL.n145 9.3005
R325 VTAIL.n105 VTAIL.n104 9.3005
R326 VTAIL.n152 VTAIL.n151 9.3005
R327 VTAIL.n154 VTAIL.n153 9.3005
R328 VTAIL.n101 VTAIL.n100 9.3005
R329 VTAIL.n160 VTAIL.n159 9.3005
R330 VTAIL.n162 VTAIL.n161 9.3005
R331 VTAIL.n98 VTAIL.n95 9.3005
R332 VTAIL.n177 VTAIL.n176 9.3005
R333 VTAIL.n92 VTAIL.n91 9.3005
R334 VTAIL.n171 VTAIL.n170 9.3005
R335 VTAIL.n169 VTAIL.n168 9.3005
R336 VTAIL.n144 VTAIL.n143 9.3005
R337 VTAIL.n109 VTAIL.n108 9.3005
R338 VTAIL.n138 VTAIL.n137 9.3005
R339 VTAIL.n136 VTAIL.n135 9.3005
R340 VTAIL.n113 VTAIL.n112 9.3005
R341 VTAIL.n130 VTAIL.n129 9.3005
R342 VTAIL.n128 VTAIL.n127 9.3005
R343 VTAIL.n117 VTAIL.n116 9.3005
R344 VTAIL.n122 VTAIL.n121 9.3005
R345 VTAIL.n314 VTAIL.n290 8.92171
R346 VTAIL.n330 VTAIL.n329 8.92171
R347 VTAIL.n44 VTAIL.n20 8.92171
R348 VTAIL.n60 VTAIL.n59 8.92171
R349 VTAIL.n241 VTAIL.n240 8.92171
R350 VTAIL.n225 VTAIL.n201 8.92171
R351 VTAIL.n151 VTAIL.n150 8.92171
R352 VTAIL.n135 VTAIL.n111 8.92171
R353 VTAIL.n318 VTAIL.n317 8.14595
R354 VTAIL.n326 VTAIL.n284 8.14595
R355 VTAIL.n48 VTAIL.n47 8.14595
R356 VTAIL.n56 VTAIL.n14 8.14595
R357 VTAIL.n237 VTAIL.n195 8.14595
R358 VTAIL.n229 VTAIL.n228 8.14595
R359 VTAIL.n147 VTAIL.n105 8.14595
R360 VTAIL.n139 VTAIL.n138 8.14595
R361 VTAIL.n321 VTAIL.n288 7.3702
R362 VTAIL.n325 VTAIL.n286 7.3702
R363 VTAIL.n51 VTAIL.n18 7.3702
R364 VTAIL.n55 VTAIL.n16 7.3702
R365 VTAIL.n236 VTAIL.n197 7.3702
R366 VTAIL.n232 VTAIL.n199 7.3702
R367 VTAIL.n146 VTAIL.n107 7.3702
R368 VTAIL.n142 VTAIL.n109 7.3702
R369 VTAIL.n322 VTAIL.n321 6.59444
R370 VTAIL.n322 VTAIL.n286 6.59444
R371 VTAIL.n52 VTAIL.n51 6.59444
R372 VTAIL.n52 VTAIL.n16 6.59444
R373 VTAIL.n233 VTAIL.n197 6.59444
R374 VTAIL.n233 VTAIL.n232 6.59444
R375 VTAIL.n143 VTAIL.n107 6.59444
R376 VTAIL.n143 VTAIL.n142 6.59444
R377 VTAIL.n318 VTAIL.n288 5.81868
R378 VTAIL.n326 VTAIL.n325 5.81868
R379 VTAIL.n48 VTAIL.n18 5.81868
R380 VTAIL.n56 VTAIL.n55 5.81868
R381 VTAIL.n237 VTAIL.n236 5.81868
R382 VTAIL.n229 VTAIL.n199 5.81868
R383 VTAIL.n147 VTAIL.n146 5.81868
R384 VTAIL.n139 VTAIL.n109 5.81868
R385 VTAIL.n317 VTAIL.n290 5.04292
R386 VTAIL.n329 VTAIL.n284 5.04292
R387 VTAIL.n47 VTAIL.n20 5.04292
R388 VTAIL.n59 VTAIL.n14 5.04292
R389 VTAIL.n240 VTAIL.n195 5.04292
R390 VTAIL.n228 VTAIL.n201 5.04292
R391 VTAIL.n150 VTAIL.n105 5.04292
R392 VTAIL.n138 VTAIL.n111 5.04292
R393 VTAIL.n314 VTAIL.n313 4.26717
R394 VTAIL.n330 VTAIL.n282 4.26717
R395 VTAIL.n44 VTAIL.n43 4.26717
R396 VTAIL.n60 VTAIL.n12 4.26717
R397 VTAIL.n241 VTAIL.n193 4.26717
R398 VTAIL.n225 VTAIL.n224 4.26717
R399 VTAIL.n151 VTAIL.n103 4.26717
R400 VTAIL.n135 VTAIL.n134 4.26717
R401 VTAIL.n300 VTAIL.n299 3.70982
R402 VTAIL.n30 VTAIL.n29 3.70982
R403 VTAIL.n211 VTAIL.n210 3.70982
R404 VTAIL.n121 VTAIL.n120 3.70982
R405 VTAIL.n310 VTAIL.n292 3.49141
R406 VTAIL.n334 VTAIL.n333 3.49141
R407 VTAIL.n358 VTAIL.n270 3.49141
R408 VTAIL.n40 VTAIL.n22 3.49141
R409 VTAIL.n64 VTAIL.n63 3.49141
R410 VTAIL.n88 VTAIL.n0 3.49141
R411 VTAIL.n268 VTAIL.n180 3.49141
R412 VTAIL.n245 VTAIL.n244 3.49141
R413 VTAIL.n221 VTAIL.n203 3.49141
R414 VTAIL.n178 VTAIL.n90 3.49141
R415 VTAIL.n155 VTAIL.n154 3.49141
R416 VTAIL.n131 VTAIL.n113 3.49141
R417 VTAIL.n309 VTAIL.n294 2.71565
R418 VTAIL.n337 VTAIL.n280 2.71565
R419 VTAIL.n356 VTAIL.n355 2.71565
R420 VTAIL.n39 VTAIL.n24 2.71565
R421 VTAIL.n67 VTAIL.n10 2.71565
R422 VTAIL.n86 VTAIL.n85 2.71565
R423 VTAIL.n266 VTAIL.n265 2.71565
R424 VTAIL.n248 VTAIL.n191 2.71565
R425 VTAIL.n220 VTAIL.n205 2.71565
R426 VTAIL.n176 VTAIL.n175 2.71565
R427 VTAIL.n158 VTAIL.n101 2.71565
R428 VTAIL.n130 VTAIL.n115 2.71565
R429 VTAIL.n306 VTAIL.n305 1.93989
R430 VTAIL.n338 VTAIL.n278 1.93989
R431 VTAIL.n352 VTAIL.n272 1.93989
R432 VTAIL.n36 VTAIL.n35 1.93989
R433 VTAIL.n68 VTAIL.n8 1.93989
R434 VTAIL.n82 VTAIL.n2 1.93989
R435 VTAIL.n262 VTAIL.n182 1.93989
R436 VTAIL.n249 VTAIL.n189 1.93989
R437 VTAIL.n217 VTAIL.n216 1.93989
R438 VTAIL.n172 VTAIL.n92 1.93989
R439 VTAIL.n159 VTAIL.n99 1.93989
R440 VTAIL.n127 VTAIL.n126 1.93989
R441 VTAIL.n302 VTAIL.n296 1.16414
R442 VTAIL.n343 VTAIL.n341 1.16414
R443 VTAIL.n351 VTAIL.n274 1.16414
R444 VTAIL.n32 VTAIL.n26 1.16414
R445 VTAIL.n73 VTAIL.n71 1.16414
R446 VTAIL.n81 VTAIL.n4 1.16414
R447 VTAIL.n261 VTAIL.n184 1.16414
R448 VTAIL.n253 VTAIL.n252 1.16414
R449 VTAIL.n213 VTAIL.n207 1.16414
R450 VTAIL.n171 VTAIL.n94 1.16414
R451 VTAIL.n163 VTAIL.n162 1.16414
R452 VTAIL.n123 VTAIL.n117 1.16414
R453 VTAIL.n269 VTAIL.n179 0.914293
R454 VTAIL VTAIL.n89 0.7505
R455 VTAIL.n301 VTAIL.n298 0.388379
R456 VTAIL.n342 VTAIL.n276 0.388379
R457 VTAIL.n348 VTAIL.n347 0.388379
R458 VTAIL.n31 VTAIL.n28 0.388379
R459 VTAIL.n72 VTAIL.n6 0.388379
R460 VTAIL.n78 VTAIL.n77 0.388379
R461 VTAIL.n258 VTAIL.n257 0.388379
R462 VTAIL.n188 VTAIL.n186 0.388379
R463 VTAIL.n212 VTAIL.n209 0.388379
R464 VTAIL.n168 VTAIL.n167 0.388379
R465 VTAIL.n98 VTAIL.n96 0.388379
R466 VTAIL.n122 VTAIL.n119 0.388379
R467 VTAIL VTAIL.n359 0.164293
R468 VTAIL.n300 VTAIL.n295 0.155672
R469 VTAIL.n307 VTAIL.n295 0.155672
R470 VTAIL.n308 VTAIL.n307 0.155672
R471 VTAIL.n308 VTAIL.n291 0.155672
R472 VTAIL.n315 VTAIL.n291 0.155672
R473 VTAIL.n316 VTAIL.n315 0.155672
R474 VTAIL.n316 VTAIL.n287 0.155672
R475 VTAIL.n323 VTAIL.n287 0.155672
R476 VTAIL.n324 VTAIL.n323 0.155672
R477 VTAIL.n324 VTAIL.n283 0.155672
R478 VTAIL.n331 VTAIL.n283 0.155672
R479 VTAIL.n332 VTAIL.n331 0.155672
R480 VTAIL.n332 VTAIL.n279 0.155672
R481 VTAIL.n339 VTAIL.n279 0.155672
R482 VTAIL.n340 VTAIL.n339 0.155672
R483 VTAIL.n340 VTAIL.n275 0.155672
R484 VTAIL.n349 VTAIL.n275 0.155672
R485 VTAIL.n350 VTAIL.n349 0.155672
R486 VTAIL.n350 VTAIL.n271 0.155672
R487 VTAIL.n357 VTAIL.n271 0.155672
R488 VTAIL.n30 VTAIL.n25 0.155672
R489 VTAIL.n37 VTAIL.n25 0.155672
R490 VTAIL.n38 VTAIL.n37 0.155672
R491 VTAIL.n38 VTAIL.n21 0.155672
R492 VTAIL.n45 VTAIL.n21 0.155672
R493 VTAIL.n46 VTAIL.n45 0.155672
R494 VTAIL.n46 VTAIL.n17 0.155672
R495 VTAIL.n53 VTAIL.n17 0.155672
R496 VTAIL.n54 VTAIL.n53 0.155672
R497 VTAIL.n54 VTAIL.n13 0.155672
R498 VTAIL.n61 VTAIL.n13 0.155672
R499 VTAIL.n62 VTAIL.n61 0.155672
R500 VTAIL.n62 VTAIL.n9 0.155672
R501 VTAIL.n69 VTAIL.n9 0.155672
R502 VTAIL.n70 VTAIL.n69 0.155672
R503 VTAIL.n70 VTAIL.n5 0.155672
R504 VTAIL.n79 VTAIL.n5 0.155672
R505 VTAIL.n80 VTAIL.n79 0.155672
R506 VTAIL.n80 VTAIL.n1 0.155672
R507 VTAIL.n87 VTAIL.n1 0.155672
R508 VTAIL.n267 VTAIL.n181 0.155672
R509 VTAIL.n260 VTAIL.n181 0.155672
R510 VTAIL.n260 VTAIL.n259 0.155672
R511 VTAIL.n259 VTAIL.n185 0.155672
R512 VTAIL.n251 VTAIL.n185 0.155672
R513 VTAIL.n251 VTAIL.n250 0.155672
R514 VTAIL.n250 VTAIL.n190 0.155672
R515 VTAIL.n243 VTAIL.n190 0.155672
R516 VTAIL.n243 VTAIL.n242 0.155672
R517 VTAIL.n242 VTAIL.n194 0.155672
R518 VTAIL.n235 VTAIL.n194 0.155672
R519 VTAIL.n235 VTAIL.n234 0.155672
R520 VTAIL.n234 VTAIL.n198 0.155672
R521 VTAIL.n227 VTAIL.n198 0.155672
R522 VTAIL.n227 VTAIL.n226 0.155672
R523 VTAIL.n226 VTAIL.n202 0.155672
R524 VTAIL.n219 VTAIL.n202 0.155672
R525 VTAIL.n219 VTAIL.n218 0.155672
R526 VTAIL.n218 VTAIL.n206 0.155672
R527 VTAIL.n211 VTAIL.n206 0.155672
R528 VTAIL.n177 VTAIL.n91 0.155672
R529 VTAIL.n170 VTAIL.n91 0.155672
R530 VTAIL.n170 VTAIL.n169 0.155672
R531 VTAIL.n169 VTAIL.n95 0.155672
R532 VTAIL.n161 VTAIL.n95 0.155672
R533 VTAIL.n161 VTAIL.n160 0.155672
R534 VTAIL.n160 VTAIL.n100 0.155672
R535 VTAIL.n153 VTAIL.n100 0.155672
R536 VTAIL.n153 VTAIL.n152 0.155672
R537 VTAIL.n152 VTAIL.n104 0.155672
R538 VTAIL.n145 VTAIL.n104 0.155672
R539 VTAIL.n145 VTAIL.n144 0.155672
R540 VTAIL.n144 VTAIL.n108 0.155672
R541 VTAIL.n137 VTAIL.n108 0.155672
R542 VTAIL.n137 VTAIL.n136 0.155672
R543 VTAIL.n136 VTAIL.n112 0.155672
R544 VTAIL.n129 VTAIL.n112 0.155672
R545 VTAIL.n129 VTAIL.n128 0.155672
R546 VTAIL.n128 VTAIL.n116 0.155672
R547 VTAIL.n121 VTAIL.n116 0.155672
R548 VDD1.n84 VDD1.n0 756.745
R549 VDD1.n173 VDD1.n89 756.745
R550 VDD1.n85 VDD1.n84 585
R551 VDD1.n83 VDD1.n82 585
R552 VDD1.n4 VDD1.n3 585
R553 VDD1.n77 VDD1.n76 585
R554 VDD1.n75 VDD1.n6 585
R555 VDD1.n74 VDD1.n73 585
R556 VDD1.n9 VDD1.n7 585
R557 VDD1.n68 VDD1.n67 585
R558 VDD1.n66 VDD1.n65 585
R559 VDD1.n13 VDD1.n12 585
R560 VDD1.n60 VDD1.n59 585
R561 VDD1.n58 VDD1.n57 585
R562 VDD1.n17 VDD1.n16 585
R563 VDD1.n52 VDD1.n51 585
R564 VDD1.n50 VDD1.n49 585
R565 VDD1.n21 VDD1.n20 585
R566 VDD1.n44 VDD1.n43 585
R567 VDD1.n42 VDD1.n41 585
R568 VDD1.n25 VDD1.n24 585
R569 VDD1.n36 VDD1.n35 585
R570 VDD1.n34 VDD1.n33 585
R571 VDD1.n29 VDD1.n28 585
R572 VDD1.n117 VDD1.n116 585
R573 VDD1.n122 VDD1.n121 585
R574 VDD1.n124 VDD1.n123 585
R575 VDD1.n113 VDD1.n112 585
R576 VDD1.n130 VDD1.n129 585
R577 VDD1.n132 VDD1.n131 585
R578 VDD1.n109 VDD1.n108 585
R579 VDD1.n138 VDD1.n137 585
R580 VDD1.n140 VDD1.n139 585
R581 VDD1.n105 VDD1.n104 585
R582 VDD1.n146 VDD1.n145 585
R583 VDD1.n148 VDD1.n147 585
R584 VDD1.n101 VDD1.n100 585
R585 VDD1.n154 VDD1.n153 585
R586 VDD1.n156 VDD1.n155 585
R587 VDD1.n97 VDD1.n96 585
R588 VDD1.n163 VDD1.n162 585
R589 VDD1.n164 VDD1.n95 585
R590 VDD1.n166 VDD1.n165 585
R591 VDD1.n93 VDD1.n92 585
R592 VDD1.n172 VDD1.n171 585
R593 VDD1.n174 VDD1.n173 585
R594 VDD1.n30 VDD1.t1 327.466
R595 VDD1.n118 VDD1.t0 327.466
R596 VDD1.n84 VDD1.n83 171.744
R597 VDD1.n83 VDD1.n3 171.744
R598 VDD1.n76 VDD1.n3 171.744
R599 VDD1.n76 VDD1.n75 171.744
R600 VDD1.n75 VDD1.n74 171.744
R601 VDD1.n74 VDD1.n7 171.744
R602 VDD1.n67 VDD1.n7 171.744
R603 VDD1.n67 VDD1.n66 171.744
R604 VDD1.n66 VDD1.n12 171.744
R605 VDD1.n59 VDD1.n12 171.744
R606 VDD1.n59 VDD1.n58 171.744
R607 VDD1.n58 VDD1.n16 171.744
R608 VDD1.n51 VDD1.n16 171.744
R609 VDD1.n51 VDD1.n50 171.744
R610 VDD1.n50 VDD1.n20 171.744
R611 VDD1.n43 VDD1.n20 171.744
R612 VDD1.n43 VDD1.n42 171.744
R613 VDD1.n42 VDD1.n24 171.744
R614 VDD1.n35 VDD1.n24 171.744
R615 VDD1.n35 VDD1.n34 171.744
R616 VDD1.n34 VDD1.n28 171.744
R617 VDD1.n122 VDD1.n116 171.744
R618 VDD1.n123 VDD1.n122 171.744
R619 VDD1.n123 VDD1.n112 171.744
R620 VDD1.n130 VDD1.n112 171.744
R621 VDD1.n131 VDD1.n130 171.744
R622 VDD1.n131 VDD1.n108 171.744
R623 VDD1.n138 VDD1.n108 171.744
R624 VDD1.n139 VDD1.n138 171.744
R625 VDD1.n139 VDD1.n104 171.744
R626 VDD1.n146 VDD1.n104 171.744
R627 VDD1.n147 VDD1.n146 171.744
R628 VDD1.n147 VDD1.n100 171.744
R629 VDD1.n154 VDD1.n100 171.744
R630 VDD1.n155 VDD1.n154 171.744
R631 VDD1.n155 VDD1.n96 171.744
R632 VDD1.n163 VDD1.n96 171.744
R633 VDD1.n164 VDD1.n163 171.744
R634 VDD1.n165 VDD1.n164 171.744
R635 VDD1.n165 VDD1.n92 171.744
R636 VDD1.n172 VDD1.n92 171.744
R637 VDD1.n173 VDD1.n172 171.744
R638 VDD1 VDD1.n177 91.964
R639 VDD1.t1 VDD1.n28 85.8723
R640 VDD1.t0 VDD1.n116 85.8723
R641 VDD1 VDD1.n88 52.0534
R642 VDD1.n30 VDD1.n29 16.3895
R643 VDD1.n118 VDD1.n117 16.3895
R644 VDD1.n77 VDD1.n6 13.1884
R645 VDD1.n166 VDD1.n95 13.1884
R646 VDD1.n78 VDD1.n4 12.8005
R647 VDD1.n73 VDD1.n8 12.8005
R648 VDD1.n33 VDD1.n32 12.8005
R649 VDD1.n121 VDD1.n120 12.8005
R650 VDD1.n162 VDD1.n161 12.8005
R651 VDD1.n167 VDD1.n93 12.8005
R652 VDD1.n82 VDD1.n81 12.0247
R653 VDD1.n72 VDD1.n9 12.0247
R654 VDD1.n36 VDD1.n27 12.0247
R655 VDD1.n124 VDD1.n115 12.0247
R656 VDD1.n160 VDD1.n97 12.0247
R657 VDD1.n171 VDD1.n170 12.0247
R658 VDD1.n85 VDD1.n2 11.249
R659 VDD1.n69 VDD1.n68 11.249
R660 VDD1.n37 VDD1.n25 11.249
R661 VDD1.n125 VDD1.n113 11.249
R662 VDD1.n157 VDD1.n156 11.249
R663 VDD1.n174 VDD1.n91 11.249
R664 VDD1.n86 VDD1.n0 10.4732
R665 VDD1.n65 VDD1.n11 10.4732
R666 VDD1.n41 VDD1.n40 10.4732
R667 VDD1.n129 VDD1.n128 10.4732
R668 VDD1.n153 VDD1.n99 10.4732
R669 VDD1.n175 VDD1.n89 10.4732
R670 VDD1.n64 VDD1.n13 9.69747
R671 VDD1.n44 VDD1.n23 9.69747
R672 VDD1.n132 VDD1.n111 9.69747
R673 VDD1.n152 VDD1.n101 9.69747
R674 VDD1.n88 VDD1.n87 9.45567
R675 VDD1.n177 VDD1.n176 9.45567
R676 VDD1.n56 VDD1.n55 9.3005
R677 VDD1.n15 VDD1.n14 9.3005
R678 VDD1.n62 VDD1.n61 9.3005
R679 VDD1.n64 VDD1.n63 9.3005
R680 VDD1.n11 VDD1.n10 9.3005
R681 VDD1.n70 VDD1.n69 9.3005
R682 VDD1.n72 VDD1.n71 9.3005
R683 VDD1.n8 VDD1.n5 9.3005
R684 VDD1.n87 VDD1.n86 9.3005
R685 VDD1.n2 VDD1.n1 9.3005
R686 VDD1.n81 VDD1.n80 9.3005
R687 VDD1.n79 VDD1.n78 9.3005
R688 VDD1.n54 VDD1.n53 9.3005
R689 VDD1.n19 VDD1.n18 9.3005
R690 VDD1.n48 VDD1.n47 9.3005
R691 VDD1.n46 VDD1.n45 9.3005
R692 VDD1.n23 VDD1.n22 9.3005
R693 VDD1.n40 VDD1.n39 9.3005
R694 VDD1.n38 VDD1.n37 9.3005
R695 VDD1.n27 VDD1.n26 9.3005
R696 VDD1.n32 VDD1.n31 9.3005
R697 VDD1.n176 VDD1.n175 9.3005
R698 VDD1.n91 VDD1.n90 9.3005
R699 VDD1.n170 VDD1.n169 9.3005
R700 VDD1.n168 VDD1.n167 9.3005
R701 VDD1.n107 VDD1.n106 9.3005
R702 VDD1.n136 VDD1.n135 9.3005
R703 VDD1.n134 VDD1.n133 9.3005
R704 VDD1.n111 VDD1.n110 9.3005
R705 VDD1.n128 VDD1.n127 9.3005
R706 VDD1.n126 VDD1.n125 9.3005
R707 VDD1.n115 VDD1.n114 9.3005
R708 VDD1.n120 VDD1.n119 9.3005
R709 VDD1.n142 VDD1.n141 9.3005
R710 VDD1.n144 VDD1.n143 9.3005
R711 VDD1.n103 VDD1.n102 9.3005
R712 VDD1.n150 VDD1.n149 9.3005
R713 VDD1.n152 VDD1.n151 9.3005
R714 VDD1.n99 VDD1.n98 9.3005
R715 VDD1.n158 VDD1.n157 9.3005
R716 VDD1.n160 VDD1.n159 9.3005
R717 VDD1.n161 VDD1.n94 9.3005
R718 VDD1.n61 VDD1.n60 8.92171
R719 VDD1.n45 VDD1.n21 8.92171
R720 VDD1.n133 VDD1.n109 8.92171
R721 VDD1.n149 VDD1.n148 8.92171
R722 VDD1.n57 VDD1.n15 8.14595
R723 VDD1.n49 VDD1.n48 8.14595
R724 VDD1.n137 VDD1.n136 8.14595
R725 VDD1.n145 VDD1.n103 8.14595
R726 VDD1.n56 VDD1.n17 7.3702
R727 VDD1.n52 VDD1.n19 7.3702
R728 VDD1.n140 VDD1.n107 7.3702
R729 VDD1.n144 VDD1.n105 7.3702
R730 VDD1.n53 VDD1.n17 6.59444
R731 VDD1.n53 VDD1.n52 6.59444
R732 VDD1.n141 VDD1.n140 6.59444
R733 VDD1.n141 VDD1.n105 6.59444
R734 VDD1.n57 VDD1.n56 5.81868
R735 VDD1.n49 VDD1.n19 5.81868
R736 VDD1.n137 VDD1.n107 5.81868
R737 VDD1.n145 VDD1.n144 5.81868
R738 VDD1.n60 VDD1.n15 5.04292
R739 VDD1.n48 VDD1.n21 5.04292
R740 VDD1.n136 VDD1.n109 5.04292
R741 VDD1.n148 VDD1.n103 5.04292
R742 VDD1.n61 VDD1.n13 4.26717
R743 VDD1.n45 VDD1.n44 4.26717
R744 VDD1.n133 VDD1.n132 4.26717
R745 VDD1.n149 VDD1.n101 4.26717
R746 VDD1.n31 VDD1.n30 3.70982
R747 VDD1.n119 VDD1.n118 3.70982
R748 VDD1.n88 VDD1.n0 3.49141
R749 VDD1.n65 VDD1.n64 3.49141
R750 VDD1.n41 VDD1.n23 3.49141
R751 VDD1.n129 VDD1.n111 3.49141
R752 VDD1.n153 VDD1.n152 3.49141
R753 VDD1.n177 VDD1.n89 3.49141
R754 VDD1.n86 VDD1.n85 2.71565
R755 VDD1.n68 VDD1.n11 2.71565
R756 VDD1.n40 VDD1.n25 2.71565
R757 VDD1.n128 VDD1.n113 2.71565
R758 VDD1.n156 VDD1.n99 2.71565
R759 VDD1.n175 VDD1.n174 2.71565
R760 VDD1.n82 VDD1.n2 1.93989
R761 VDD1.n69 VDD1.n9 1.93989
R762 VDD1.n37 VDD1.n36 1.93989
R763 VDD1.n125 VDD1.n124 1.93989
R764 VDD1.n157 VDD1.n97 1.93989
R765 VDD1.n171 VDD1.n91 1.93989
R766 VDD1.n81 VDD1.n4 1.16414
R767 VDD1.n73 VDD1.n72 1.16414
R768 VDD1.n33 VDD1.n27 1.16414
R769 VDD1.n121 VDD1.n115 1.16414
R770 VDD1.n162 VDD1.n160 1.16414
R771 VDD1.n170 VDD1.n93 1.16414
R772 VDD1.n78 VDD1.n77 0.388379
R773 VDD1.n8 VDD1.n6 0.388379
R774 VDD1.n32 VDD1.n29 0.388379
R775 VDD1.n120 VDD1.n117 0.388379
R776 VDD1.n161 VDD1.n95 0.388379
R777 VDD1.n167 VDD1.n166 0.388379
R778 VDD1.n87 VDD1.n1 0.155672
R779 VDD1.n80 VDD1.n1 0.155672
R780 VDD1.n80 VDD1.n79 0.155672
R781 VDD1.n79 VDD1.n5 0.155672
R782 VDD1.n71 VDD1.n5 0.155672
R783 VDD1.n71 VDD1.n70 0.155672
R784 VDD1.n70 VDD1.n10 0.155672
R785 VDD1.n63 VDD1.n10 0.155672
R786 VDD1.n63 VDD1.n62 0.155672
R787 VDD1.n62 VDD1.n14 0.155672
R788 VDD1.n55 VDD1.n14 0.155672
R789 VDD1.n55 VDD1.n54 0.155672
R790 VDD1.n54 VDD1.n18 0.155672
R791 VDD1.n47 VDD1.n18 0.155672
R792 VDD1.n47 VDD1.n46 0.155672
R793 VDD1.n46 VDD1.n22 0.155672
R794 VDD1.n39 VDD1.n22 0.155672
R795 VDD1.n39 VDD1.n38 0.155672
R796 VDD1.n38 VDD1.n26 0.155672
R797 VDD1.n31 VDD1.n26 0.155672
R798 VDD1.n119 VDD1.n114 0.155672
R799 VDD1.n126 VDD1.n114 0.155672
R800 VDD1.n127 VDD1.n126 0.155672
R801 VDD1.n127 VDD1.n110 0.155672
R802 VDD1.n134 VDD1.n110 0.155672
R803 VDD1.n135 VDD1.n134 0.155672
R804 VDD1.n135 VDD1.n106 0.155672
R805 VDD1.n142 VDD1.n106 0.155672
R806 VDD1.n143 VDD1.n142 0.155672
R807 VDD1.n143 VDD1.n102 0.155672
R808 VDD1.n150 VDD1.n102 0.155672
R809 VDD1.n151 VDD1.n150 0.155672
R810 VDD1.n151 VDD1.n98 0.155672
R811 VDD1.n158 VDD1.n98 0.155672
R812 VDD1.n159 VDD1.n158 0.155672
R813 VDD1.n159 VDD1.n94 0.155672
R814 VDD1.n168 VDD1.n94 0.155672
R815 VDD1.n169 VDD1.n168 0.155672
R816 VDD1.n169 VDD1.n90 0.155672
R817 VDD1.n176 VDD1.n90 0.155672
R818 B.n114 B.t9 761.74
R819 B.n122 B.t3 761.74
R820 B.n36 B.t6 761.74
R821 B.n44 B.t0 761.74
R822 B.n399 B.n72 585
R823 B.n401 B.n400 585
R824 B.n402 B.n71 585
R825 B.n404 B.n403 585
R826 B.n405 B.n70 585
R827 B.n407 B.n406 585
R828 B.n408 B.n69 585
R829 B.n410 B.n409 585
R830 B.n411 B.n68 585
R831 B.n413 B.n412 585
R832 B.n414 B.n67 585
R833 B.n416 B.n415 585
R834 B.n417 B.n66 585
R835 B.n419 B.n418 585
R836 B.n420 B.n65 585
R837 B.n422 B.n421 585
R838 B.n423 B.n64 585
R839 B.n425 B.n424 585
R840 B.n426 B.n63 585
R841 B.n428 B.n427 585
R842 B.n429 B.n62 585
R843 B.n431 B.n430 585
R844 B.n432 B.n61 585
R845 B.n434 B.n433 585
R846 B.n435 B.n60 585
R847 B.n437 B.n436 585
R848 B.n438 B.n59 585
R849 B.n440 B.n439 585
R850 B.n441 B.n58 585
R851 B.n443 B.n442 585
R852 B.n444 B.n57 585
R853 B.n446 B.n445 585
R854 B.n447 B.n56 585
R855 B.n449 B.n448 585
R856 B.n450 B.n55 585
R857 B.n452 B.n451 585
R858 B.n453 B.n54 585
R859 B.n455 B.n454 585
R860 B.n456 B.n53 585
R861 B.n458 B.n457 585
R862 B.n459 B.n52 585
R863 B.n461 B.n460 585
R864 B.n462 B.n51 585
R865 B.n464 B.n463 585
R866 B.n465 B.n50 585
R867 B.n467 B.n466 585
R868 B.n468 B.n49 585
R869 B.n470 B.n469 585
R870 B.n471 B.n48 585
R871 B.n473 B.n472 585
R872 B.n474 B.n47 585
R873 B.n476 B.n475 585
R874 B.n477 B.n46 585
R875 B.n479 B.n478 585
R876 B.n481 B.n43 585
R877 B.n483 B.n482 585
R878 B.n484 B.n42 585
R879 B.n486 B.n485 585
R880 B.n487 B.n41 585
R881 B.n489 B.n488 585
R882 B.n490 B.n40 585
R883 B.n492 B.n491 585
R884 B.n493 B.n39 585
R885 B.n495 B.n494 585
R886 B.n497 B.n496 585
R887 B.n498 B.n35 585
R888 B.n500 B.n499 585
R889 B.n501 B.n34 585
R890 B.n503 B.n502 585
R891 B.n504 B.n33 585
R892 B.n506 B.n505 585
R893 B.n507 B.n32 585
R894 B.n509 B.n508 585
R895 B.n510 B.n31 585
R896 B.n512 B.n511 585
R897 B.n513 B.n30 585
R898 B.n515 B.n514 585
R899 B.n516 B.n29 585
R900 B.n518 B.n517 585
R901 B.n519 B.n28 585
R902 B.n521 B.n520 585
R903 B.n522 B.n27 585
R904 B.n524 B.n523 585
R905 B.n525 B.n26 585
R906 B.n527 B.n526 585
R907 B.n528 B.n25 585
R908 B.n530 B.n529 585
R909 B.n531 B.n24 585
R910 B.n533 B.n532 585
R911 B.n534 B.n23 585
R912 B.n536 B.n535 585
R913 B.n537 B.n22 585
R914 B.n539 B.n538 585
R915 B.n540 B.n21 585
R916 B.n542 B.n541 585
R917 B.n543 B.n20 585
R918 B.n545 B.n544 585
R919 B.n546 B.n19 585
R920 B.n548 B.n547 585
R921 B.n549 B.n18 585
R922 B.n551 B.n550 585
R923 B.n552 B.n17 585
R924 B.n554 B.n553 585
R925 B.n555 B.n16 585
R926 B.n557 B.n556 585
R927 B.n558 B.n15 585
R928 B.n560 B.n559 585
R929 B.n561 B.n14 585
R930 B.n563 B.n562 585
R931 B.n564 B.n13 585
R932 B.n566 B.n565 585
R933 B.n567 B.n12 585
R934 B.n569 B.n568 585
R935 B.n570 B.n11 585
R936 B.n572 B.n571 585
R937 B.n573 B.n10 585
R938 B.n575 B.n574 585
R939 B.n576 B.n9 585
R940 B.n398 B.n397 585
R941 B.n396 B.n73 585
R942 B.n395 B.n394 585
R943 B.n393 B.n74 585
R944 B.n392 B.n391 585
R945 B.n390 B.n75 585
R946 B.n389 B.n388 585
R947 B.n387 B.n76 585
R948 B.n386 B.n385 585
R949 B.n384 B.n77 585
R950 B.n383 B.n382 585
R951 B.n381 B.n78 585
R952 B.n380 B.n379 585
R953 B.n378 B.n79 585
R954 B.n377 B.n376 585
R955 B.n375 B.n80 585
R956 B.n374 B.n373 585
R957 B.n372 B.n81 585
R958 B.n371 B.n370 585
R959 B.n369 B.n82 585
R960 B.n368 B.n367 585
R961 B.n366 B.n83 585
R962 B.n365 B.n364 585
R963 B.n363 B.n84 585
R964 B.n362 B.n361 585
R965 B.n360 B.n85 585
R966 B.n359 B.n358 585
R967 B.n357 B.n86 585
R968 B.n356 B.n355 585
R969 B.n177 B.n150 585
R970 B.n179 B.n178 585
R971 B.n180 B.n149 585
R972 B.n182 B.n181 585
R973 B.n183 B.n148 585
R974 B.n185 B.n184 585
R975 B.n186 B.n147 585
R976 B.n188 B.n187 585
R977 B.n189 B.n146 585
R978 B.n191 B.n190 585
R979 B.n192 B.n145 585
R980 B.n194 B.n193 585
R981 B.n195 B.n144 585
R982 B.n197 B.n196 585
R983 B.n198 B.n143 585
R984 B.n200 B.n199 585
R985 B.n201 B.n142 585
R986 B.n203 B.n202 585
R987 B.n204 B.n141 585
R988 B.n206 B.n205 585
R989 B.n207 B.n140 585
R990 B.n209 B.n208 585
R991 B.n210 B.n139 585
R992 B.n212 B.n211 585
R993 B.n213 B.n138 585
R994 B.n215 B.n214 585
R995 B.n216 B.n137 585
R996 B.n218 B.n217 585
R997 B.n219 B.n136 585
R998 B.n221 B.n220 585
R999 B.n222 B.n135 585
R1000 B.n224 B.n223 585
R1001 B.n225 B.n134 585
R1002 B.n227 B.n226 585
R1003 B.n228 B.n133 585
R1004 B.n230 B.n229 585
R1005 B.n231 B.n132 585
R1006 B.n233 B.n232 585
R1007 B.n234 B.n131 585
R1008 B.n236 B.n235 585
R1009 B.n237 B.n130 585
R1010 B.n239 B.n238 585
R1011 B.n240 B.n129 585
R1012 B.n242 B.n241 585
R1013 B.n243 B.n128 585
R1014 B.n245 B.n244 585
R1015 B.n246 B.n127 585
R1016 B.n248 B.n247 585
R1017 B.n249 B.n126 585
R1018 B.n251 B.n250 585
R1019 B.n252 B.n125 585
R1020 B.n254 B.n253 585
R1021 B.n255 B.n124 585
R1022 B.n257 B.n256 585
R1023 B.n259 B.n121 585
R1024 B.n261 B.n260 585
R1025 B.n262 B.n120 585
R1026 B.n264 B.n263 585
R1027 B.n265 B.n119 585
R1028 B.n267 B.n266 585
R1029 B.n268 B.n118 585
R1030 B.n270 B.n269 585
R1031 B.n271 B.n117 585
R1032 B.n273 B.n272 585
R1033 B.n275 B.n274 585
R1034 B.n276 B.n113 585
R1035 B.n278 B.n277 585
R1036 B.n279 B.n112 585
R1037 B.n281 B.n280 585
R1038 B.n282 B.n111 585
R1039 B.n284 B.n283 585
R1040 B.n285 B.n110 585
R1041 B.n287 B.n286 585
R1042 B.n288 B.n109 585
R1043 B.n290 B.n289 585
R1044 B.n291 B.n108 585
R1045 B.n293 B.n292 585
R1046 B.n294 B.n107 585
R1047 B.n296 B.n295 585
R1048 B.n297 B.n106 585
R1049 B.n299 B.n298 585
R1050 B.n300 B.n105 585
R1051 B.n302 B.n301 585
R1052 B.n303 B.n104 585
R1053 B.n305 B.n304 585
R1054 B.n306 B.n103 585
R1055 B.n308 B.n307 585
R1056 B.n309 B.n102 585
R1057 B.n311 B.n310 585
R1058 B.n312 B.n101 585
R1059 B.n314 B.n313 585
R1060 B.n315 B.n100 585
R1061 B.n317 B.n316 585
R1062 B.n318 B.n99 585
R1063 B.n320 B.n319 585
R1064 B.n321 B.n98 585
R1065 B.n323 B.n322 585
R1066 B.n324 B.n97 585
R1067 B.n326 B.n325 585
R1068 B.n327 B.n96 585
R1069 B.n329 B.n328 585
R1070 B.n330 B.n95 585
R1071 B.n332 B.n331 585
R1072 B.n333 B.n94 585
R1073 B.n335 B.n334 585
R1074 B.n336 B.n93 585
R1075 B.n338 B.n337 585
R1076 B.n339 B.n92 585
R1077 B.n341 B.n340 585
R1078 B.n342 B.n91 585
R1079 B.n344 B.n343 585
R1080 B.n345 B.n90 585
R1081 B.n347 B.n346 585
R1082 B.n348 B.n89 585
R1083 B.n350 B.n349 585
R1084 B.n351 B.n88 585
R1085 B.n353 B.n352 585
R1086 B.n354 B.n87 585
R1087 B.n176 B.n175 585
R1088 B.n174 B.n151 585
R1089 B.n173 B.n172 585
R1090 B.n171 B.n152 585
R1091 B.n170 B.n169 585
R1092 B.n168 B.n153 585
R1093 B.n167 B.n166 585
R1094 B.n165 B.n154 585
R1095 B.n164 B.n163 585
R1096 B.n162 B.n155 585
R1097 B.n161 B.n160 585
R1098 B.n159 B.n156 585
R1099 B.n158 B.n157 585
R1100 B.n2 B.n0 585
R1101 B.n597 B.n1 585
R1102 B.n596 B.n595 585
R1103 B.n594 B.n3 585
R1104 B.n593 B.n592 585
R1105 B.n591 B.n4 585
R1106 B.n590 B.n589 585
R1107 B.n588 B.n5 585
R1108 B.n587 B.n586 585
R1109 B.n585 B.n6 585
R1110 B.n584 B.n583 585
R1111 B.n582 B.n7 585
R1112 B.n581 B.n580 585
R1113 B.n579 B.n8 585
R1114 B.n578 B.n577 585
R1115 B.n599 B.n598 585
R1116 B.n177 B.n176 511.721
R1117 B.n578 B.n9 511.721
R1118 B.n356 B.n87 511.721
R1119 B.n399 B.n398 511.721
R1120 B.n114 B.t11 471.901
R1121 B.n44 B.t1 471.901
R1122 B.n122 B.t5 471.901
R1123 B.n36 B.t7 471.901
R1124 B.n115 B.t10 451.925
R1125 B.n45 B.t2 451.925
R1126 B.n123 B.t4 451.925
R1127 B.n37 B.t8 451.925
R1128 B.n176 B.n151 163.367
R1129 B.n172 B.n151 163.367
R1130 B.n172 B.n171 163.367
R1131 B.n171 B.n170 163.367
R1132 B.n170 B.n153 163.367
R1133 B.n166 B.n153 163.367
R1134 B.n166 B.n165 163.367
R1135 B.n165 B.n164 163.367
R1136 B.n164 B.n155 163.367
R1137 B.n160 B.n155 163.367
R1138 B.n160 B.n159 163.367
R1139 B.n159 B.n158 163.367
R1140 B.n158 B.n2 163.367
R1141 B.n598 B.n2 163.367
R1142 B.n598 B.n597 163.367
R1143 B.n597 B.n596 163.367
R1144 B.n596 B.n3 163.367
R1145 B.n592 B.n3 163.367
R1146 B.n592 B.n591 163.367
R1147 B.n591 B.n590 163.367
R1148 B.n590 B.n5 163.367
R1149 B.n586 B.n5 163.367
R1150 B.n586 B.n585 163.367
R1151 B.n585 B.n584 163.367
R1152 B.n584 B.n7 163.367
R1153 B.n580 B.n7 163.367
R1154 B.n580 B.n579 163.367
R1155 B.n579 B.n578 163.367
R1156 B.n178 B.n177 163.367
R1157 B.n178 B.n149 163.367
R1158 B.n182 B.n149 163.367
R1159 B.n183 B.n182 163.367
R1160 B.n184 B.n183 163.367
R1161 B.n184 B.n147 163.367
R1162 B.n188 B.n147 163.367
R1163 B.n189 B.n188 163.367
R1164 B.n190 B.n189 163.367
R1165 B.n190 B.n145 163.367
R1166 B.n194 B.n145 163.367
R1167 B.n195 B.n194 163.367
R1168 B.n196 B.n195 163.367
R1169 B.n196 B.n143 163.367
R1170 B.n200 B.n143 163.367
R1171 B.n201 B.n200 163.367
R1172 B.n202 B.n201 163.367
R1173 B.n202 B.n141 163.367
R1174 B.n206 B.n141 163.367
R1175 B.n207 B.n206 163.367
R1176 B.n208 B.n207 163.367
R1177 B.n208 B.n139 163.367
R1178 B.n212 B.n139 163.367
R1179 B.n213 B.n212 163.367
R1180 B.n214 B.n213 163.367
R1181 B.n214 B.n137 163.367
R1182 B.n218 B.n137 163.367
R1183 B.n219 B.n218 163.367
R1184 B.n220 B.n219 163.367
R1185 B.n220 B.n135 163.367
R1186 B.n224 B.n135 163.367
R1187 B.n225 B.n224 163.367
R1188 B.n226 B.n225 163.367
R1189 B.n226 B.n133 163.367
R1190 B.n230 B.n133 163.367
R1191 B.n231 B.n230 163.367
R1192 B.n232 B.n231 163.367
R1193 B.n232 B.n131 163.367
R1194 B.n236 B.n131 163.367
R1195 B.n237 B.n236 163.367
R1196 B.n238 B.n237 163.367
R1197 B.n238 B.n129 163.367
R1198 B.n242 B.n129 163.367
R1199 B.n243 B.n242 163.367
R1200 B.n244 B.n243 163.367
R1201 B.n244 B.n127 163.367
R1202 B.n248 B.n127 163.367
R1203 B.n249 B.n248 163.367
R1204 B.n250 B.n249 163.367
R1205 B.n250 B.n125 163.367
R1206 B.n254 B.n125 163.367
R1207 B.n255 B.n254 163.367
R1208 B.n256 B.n255 163.367
R1209 B.n256 B.n121 163.367
R1210 B.n261 B.n121 163.367
R1211 B.n262 B.n261 163.367
R1212 B.n263 B.n262 163.367
R1213 B.n263 B.n119 163.367
R1214 B.n267 B.n119 163.367
R1215 B.n268 B.n267 163.367
R1216 B.n269 B.n268 163.367
R1217 B.n269 B.n117 163.367
R1218 B.n273 B.n117 163.367
R1219 B.n274 B.n273 163.367
R1220 B.n274 B.n113 163.367
R1221 B.n278 B.n113 163.367
R1222 B.n279 B.n278 163.367
R1223 B.n280 B.n279 163.367
R1224 B.n280 B.n111 163.367
R1225 B.n284 B.n111 163.367
R1226 B.n285 B.n284 163.367
R1227 B.n286 B.n285 163.367
R1228 B.n286 B.n109 163.367
R1229 B.n290 B.n109 163.367
R1230 B.n291 B.n290 163.367
R1231 B.n292 B.n291 163.367
R1232 B.n292 B.n107 163.367
R1233 B.n296 B.n107 163.367
R1234 B.n297 B.n296 163.367
R1235 B.n298 B.n297 163.367
R1236 B.n298 B.n105 163.367
R1237 B.n302 B.n105 163.367
R1238 B.n303 B.n302 163.367
R1239 B.n304 B.n303 163.367
R1240 B.n304 B.n103 163.367
R1241 B.n308 B.n103 163.367
R1242 B.n309 B.n308 163.367
R1243 B.n310 B.n309 163.367
R1244 B.n310 B.n101 163.367
R1245 B.n314 B.n101 163.367
R1246 B.n315 B.n314 163.367
R1247 B.n316 B.n315 163.367
R1248 B.n316 B.n99 163.367
R1249 B.n320 B.n99 163.367
R1250 B.n321 B.n320 163.367
R1251 B.n322 B.n321 163.367
R1252 B.n322 B.n97 163.367
R1253 B.n326 B.n97 163.367
R1254 B.n327 B.n326 163.367
R1255 B.n328 B.n327 163.367
R1256 B.n328 B.n95 163.367
R1257 B.n332 B.n95 163.367
R1258 B.n333 B.n332 163.367
R1259 B.n334 B.n333 163.367
R1260 B.n334 B.n93 163.367
R1261 B.n338 B.n93 163.367
R1262 B.n339 B.n338 163.367
R1263 B.n340 B.n339 163.367
R1264 B.n340 B.n91 163.367
R1265 B.n344 B.n91 163.367
R1266 B.n345 B.n344 163.367
R1267 B.n346 B.n345 163.367
R1268 B.n346 B.n89 163.367
R1269 B.n350 B.n89 163.367
R1270 B.n351 B.n350 163.367
R1271 B.n352 B.n351 163.367
R1272 B.n352 B.n87 163.367
R1273 B.n357 B.n356 163.367
R1274 B.n358 B.n357 163.367
R1275 B.n358 B.n85 163.367
R1276 B.n362 B.n85 163.367
R1277 B.n363 B.n362 163.367
R1278 B.n364 B.n363 163.367
R1279 B.n364 B.n83 163.367
R1280 B.n368 B.n83 163.367
R1281 B.n369 B.n368 163.367
R1282 B.n370 B.n369 163.367
R1283 B.n370 B.n81 163.367
R1284 B.n374 B.n81 163.367
R1285 B.n375 B.n374 163.367
R1286 B.n376 B.n375 163.367
R1287 B.n376 B.n79 163.367
R1288 B.n380 B.n79 163.367
R1289 B.n381 B.n380 163.367
R1290 B.n382 B.n381 163.367
R1291 B.n382 B.n77 163.367
R1292 B.n386 B.n77 163.367
R1293 B.n387 B.n386 163.367
R1294 B.n388 B.n387 163.367
R1295 B.n388 B.n75 163.367
R1296 B.n392 B.n75 163.367
R1297 B.n393 B.n392 163.367
R1298 B.n394 B.n393 163.367
R1299 B.n394 B.n73 163.367
R1300 B.n398 B.n73 163.367
R1301 B.n574 B.n9 163.367
R1302 B.n574 B.n573 163.367
R1303 B.n573 B.n572 163.367
R1304 B.n572 B.n11 163.367
R1305 B.n568 B.n11 163.367
R1306 B.n568 B.n567 163.367
R1307 B.n567 B.n566 163.367
R1308 B.n566 B.n13 163.367
R1309 B.n562 B.n13 163.367
R1310 B.n562 B.n561 163.367
R1311 B.n561 B.n560 163.367
R1312 B.n560 B.n15 163.367
R1313 B.n556 B.n15 163.367
R1314 B.n556 B.n555 163.367
R1315 B.n555 B.n554 163.367
R1316 B.n554 B.n17 163.367
R1317 B.n550 B.n17 163.367
R1318 B.n550 B.n549 163.367
R1319 B.n549 B.n548 163.367
R1320 B.n548 B.n19 163.367
R1321 B.n544 B.n19 163.367
R1322 B.n544 B.n543 163.367
R1323 B.n543 B.n542 163.367
R1324 B.n542 B.n21 163.367
R1325 B.n538 B.n21 163.367
R1326 B.n538 B.n537 163.367
R1327 B.n537 B.n536 163.367
R1328 B.n536 B.n23 163.367
R1329 B.n532 B.n23 163.367
R1330 B.n532 B.n531 163.367
R1331 B.n531 B.n530 163.367
R1332 B.n530 B.n25 163.367
R1333 B.n526 B.n25 163.367
R1334 B.n526 B.n525 163.367
R1335 B.n525 B.n524 163.367
R1336 B.n524 B.n27 163.367
R1337 B.n520 B.n27 163.367
R1338 B.n520 B.n519 163.367
R1339 B.n519 B.n518 163.367
R1340 B.n518 B.n29 163.367
R1341 B.n514 B.n29 163.367
R1342 B.n514 B.n513 163.367
R1343 B.n513 B.n512 163.367
R1344 B.n512 B.n31 163.367
R1345 B.n508 B.n31 163.367
R1346 B.n508 B.n507 163.367
R1347 B.n507 B.n506 163.367
R1348 B.n506 B.n33 163.367
R1349 B.n502 B.n33 163.367
R1350 B.n502 B.n501 163.367
R1351 B.n501 B.n500 163.367
R1352 B.n500 B.n35 163.367
R1353 B.n496 B.n35 163.367
R1354 B.n496 B.n495 163.367
R1355 B.n495 B.n39 163.367
R1356 B.n491 B.n39 163.367
R1357 B.n491 B.n490 163.367
R1358 B.n490 B.n489 163.367
R1359 B.n489 B.n41 163.367
R1360 B.n485 B.n41 163.367
R1361 B.n485 B.n484 163.367
R1362 B.n484 B.n483 163.367
R1363 B.n483 B.n43 163.367
R1364 B.n478 B.n43 163.367
R1365 B.n478 B.n477 163.367
R1366 B.n477 B.n476 163.367
R1367 B.n476 B.n47 163.367
R1368 B.n472 B.n47 163.367
R1369 B.n472 B.n471 163.367
R1370 B.n471 B.n470 163.367
R1371 B.n470 B.n49 163.367
R1372 B.n466 B.n49 163.367
R1373 B.n466 B.n465 163.367
R1374 B.n465 B.n464 163.367
R1375 B.n464 B.n51 163.367
R1376 B.n460 B.n51 163.367
R1377 B.n460 B.n459 163.367
R1378 B.n459 B.n458 163.367
R1379 B.n458 B.n53 163.367
R1380 B.n454 B.n53 163.367
R1381 B.n454 B.n453 163.367
R1382 B.n453 B.n452 163.367
R1383 B.n452 B.n55 163.367
R1384 B.n448 B.n55 163.367
R1385 B.n448 B.n447 163.367
R1386 B.n447 B.n446 163.367
R1387 B.n446 B.n57 163.367
R1388 B.n442 B.n57 163.367
R1389 B.n442 B.n441 163.367
R1390 B.n441 B.n440 163.367
R1391 B.n440 B.n59 163.367
R1392 B.n436 B.n59 163.367
R1393 B.n436 B.n435 163.367
R1394 B.n435 B.n434 163.367
R1395 B.n434 B.n61 163.367
R1396 B.n430 B.n61 163.367
R1397 B.n430 B.n429 163.367
R1398 B.n429 B.n428 163.367
R1399 B.n428 B.n63 163.367
R1400 B.n424 B.n63 163.367
R1401 B.n424 B.n423 163.367
R1402 B.n423 B.n422 163.367
R1403 B.n422 B.n65 163.367
R1404 B.n418 B.n65 163.367
R1405 B.n418 B.n417 163.367
R1406 B.n417 B.n416 163.367
R1407 B.n416 B.n67 163.367
R1408 B.n412 B.n67 163.367
R1409 B.n412 B.n411 163.367
R1410 B.n411 B.n410 163.367
R1411 B.n410 B.n69 163.367
R1412 B.n406 B.n69 163.367
R1413 B.n406 B.n405 163.367
R1414 B.n405 B.n404 163.367
R1415 B.n404 B.n71 163.367
R1416 B.n400 B.n71 163.367
R1417 B.n400 B.n399 163.367
R1418 B.n116 B.n115 59.5399
R1419 B.n258 B.n123 59.5399
R1420 B.n38 B.n37 59.5399
R1421 B.n480 B.n45 59.5399
R1422 B.n577 B.n576 33.2493
R1423 B.n397 B.n72 33.2493
R1424 B.n355 B.n354 33.2493
R1425 B.n175 B.n150 33.2493
R1426 B.n115 B.n114 19.9763
R1427 B.n123 B.n122 19.9763
R1428 B.n37 B.n36 19.9763
R1429 B.n45 B.n44 19.9763
R1430 B B.n599 18.0485
R1431 B.n576 B.n575 10.6151
R1432 B.n575 B.n10 10.6151
R1433 B.n571 B.n10 10.6151
R1434 B.n571 B.n570 10.6151
R1435 B.n570 B.n569 10.6151
R1436 B.n569 B.n12 10.6151
R1437 B.n565 B.n12 10.6151
R1438 B.n565 B.n564 10.6151
R1439 B.n564 B.n563 10.6151
R1440 B.n563 B.n14 10.6151
R1441 B.n559 B.n14 10.6151
R1442 B.n559 B.n558 10.6151
R1443 B.n558 B.n557 10.6151
R1444 B.n557 B.n16 10.6151
R1445 B.n553 B.n16 10.6151
R1446 B.n553 B.n552 10.6151
R1447 B.n552 B.n551 10.6151
R1448 B.n551 B.n18 10.6151
R1449 B.n547 B.n18 10.6151
R1450 B.n547 B.n546 10.6151
R1451 B.n546 B.n545 10.6151
R1452 B.n545 B.n20 10.6151
R1453 B.n541 B.n20 10.6151
R1454 B.n541 B.n540 10.6151
R1455 B.n540 B.n539 10.6151
R1456 B.n539 B.n22 10.6151
R1457 B.n535 B.n22 10.6151
R1458 B.n535 B.n534 10.6151
R1459 B.n534 B.n533 10.6151
R1460 B.n533 B.n24 10.6151
R1461 B.n529 B.n24 10.6151
R1462 B.n529 B.n528 10.6151
R1463 B.n528 B.n527 10.6151
R1464 B.n527 B.n26 10.6151
R1465 B.n523 B.n26 10.6151
R1466 B.n523 B.n522 10.6151
R1467 B.n522 B.n521 10.6151
R1468 B.n521 B.n28 10.6151
R1469 B.n517 B.n28 10.6151
R1470 B.n517 B.n516 10.6151
R1471 B.n516 B.n515 10.6151
R1472 B.n515 B.n30 10.6151
R1473 B.n511 B.n30 10.6151
R1474 B.n511 B.n510 10.6151
R1475 B.n510 B.n509 10.6151
R1476 B.n509 B.n32 10.6151
R1477 B.n505 B.n32 10.6151
R1478 B.n505 B.n504 10.6151
R1479 B.n504 B.n503 10.6151
R1480 B.n503 B.n34 10.6151
R1481 B.n499 B.n34 10.6151
R1482 B.n499 B.n498 10.6151
R1483 B.n498 B.n497 10.6151
R1484 B.n494 B.n493 10.6151
R1485 B.n493 B.n492 10.6151
R1486 B.n492 B.n40 10.6151
R1487 B.n488 B.n40 10.6151
R1488 B.n488 B.n487 10.6151
R1489 B.n487 B.n486 10.6151
R1490 B.n486 B.n42 10.6151
R1491 B.n482 B.n42 10.6151
R1492 B.n482 B.n481 10.6151
R1493 B.n479 B.n46 10.6151
R1494 B.n475 B.n46 10.6151
R1495 B.n475 B.n474 10.6151
R1496 B.n474 B.n473 10.6151
R1497 B.n473 B.n48 10.6151
R1498 B.n469 B.n48 10.6151
R1499 B.n469 B.n468 10.6151
R1500 B.n468 B.n467 10.6151
R1501 B.n467 B.n50 10.6151
R1502 B.n463 B.n50 10.6151
R1503 B.n463 B.n462 10.6151
R1504 B.n462 B.n461 10.6151
R1505 B.n461 B.n52 10.6151
R1506 B.n457 B.n52 10.6151
R1507 B.n457 B.n456 10.6151
R1508 B.n456 B.n455 10.6151
R1509 B.n455 B.n54 10.6151
R1510 B.n451 B.n54 10.6151
R1511 B.n451 B.n450 10.6151
R1512 B.n450 B.n449 10.6151
R1513 B.n449 B.n56 10.6151
R1514 B.n445 B.n56 10.6151
R1515 B.n445 B.n444 10.6151
R1516 B.n444 B.n443 10.6151
R1517 B.n443 B.n58 10.6151
R1518 B.n439 B.n58 10.6151
R1519 B.n439 B.n438 10.6151
R1520 B.n438 B.n437 10.6151
R1521 B.n437 B.n60 10.6151
R1522 B.n433 B.n60 10.6151
R1523 B.n433 B.n432 10.6151
R1524 B.n432 B.n431 10.6151
R1525 B.n431 B.n62 10.6151
R1526 B.n427 B.n62 10.6151
R1527 B.n427 B.n426 10.6151
R1528 B.n426 B.n425 10.6151
R1529 B.n425 B.n64 10.6151
R1530 B.n421 B.n64 10.6151
R1531 B.n421 B.n420 10.6151
R1532 B.n420 B.n419 10.6151
R1533 B.n419 B.n66 10.6151
R1534 B.n415 B.n66 10.6151
R1535 B.n415 B.n414 10.6151
R1536 B.n414 B.n413 10.6151
R1537 B.n413 B.n68 10.6151
R1538 B.n409 B.n68 10.6151
R1539 B.n409 B.n408 10.6151
R1540 B.n408 B.n407 10.6151
R1541 B.n407 B.n70 10.6151
R1542 B.n403 B.n70 10.6151
R1543 B.n403 B.n402 10.6151
R1544 B.n402 B.n401 10.6151
R1545 B.n401 B.n72 10.6151
R1546 B.n355 B.n86 10.6151
R1547 B.n359 B.n86 10.6151
R1548 B.n360 B.n359 10.6151
R1549 B.n361 B.n360 10.6151
R1550 B.n361 B.n84 10.6151
R1551 B.n365 B.n84 10.6151
R1552 B.n366 B.n365 10.6151
R1553 B.n367 B.n366 10.6151
R1554 B.n367 B.n82 10.6151
R1555 B.n371 B.n82 10.6151
R1556 B.n372 B.n371 10.6151
R1557 B.n373 B.n372 10.6151
R1558 B.n373 B.n80 10.6151
R1559 B.n377 B.n80 10.6151
R1560 B.n378 B.n377 10.6151
R1561 B.n379 B.n378 10.6151
R1562 B.n379 B.n78 10.6151
R1563 B.n383 B.n78 10.6151
R1564 B.n384 B.n383 10.6151
R1565 B.n385 B.n384 10.6151
R1566 B.n385 B.n76 10.6151
R1567 B.n389 B.n76 10.6151
R1568 B.n390 B.n389 10.6151
R1569 B.n391 B.n390 10.6151
R1570 B.n391 B.n74 10.6151
R1571 B.n395 B.n74 10.6151
R1572 B.n396 B.n395 10.6151
R1573 B.n397 B.n396 10.6151
R1574 B.n179 B.n150 10.6151
R1575 B.n180 B.n179 10.6151
R1576 B.n181 B.n180 10.6151
R1577 B.n181 B.n148 10.6151
R1578 B.n185 B.n148 10.6151
R1579 B.n186 B.n185 10.6151
R1580 B.n187 B.n186 10.6151
R1581 B.n187 B.n146 10.6151
R1582 B.n191 B.n146 10.6151
R1583 B.n192 B.n191 10.6151
R1584 B.n193 B.n192 10.6151
R1585 B.n193 B.n144 10.6151
R1586 B.n197 B.n144 10.6151
R1587 B.n198 B.n197 10.6151
R1588 B.n199 B.n198 10.6151
R1589 B.n199 B.n142 10.6151
R1590 B.n203 B.n142 10.6151
R1591 B.n204 B.n203 10.6151
R1592 B.n205 B.n204 10.6151
R1593 B.n205 B.n140 10.6151
R1594 B.n209 B.n140 10.6151
R1595 B.n210 B.n209 10.6151
R1596 B.n211 B.n210 10.6151
R1597 B.n211 B.n138 10.6151
R1598 B.n215 B.n138 10.6151
R1599 B.n216 B.n215 10.6151
R1600 B.n217 B.n216 10.6151
R1601 B.n217 B.n136 10.6151
R1602 B.n221 B.n136 10.6151
R1603 B.n222 B.n221 10.6151
R1604 B.n223 B.n222 10.6151
R1605 B.n223 B.n134 10.6151
R1606 B.n227 B.n134 10.6151
R1607 B.n228 B.n227 10.6151
R1608 B.n229 B.n228 10.6151
R1609 B.n229 B.n132 10.6151
R1610 B.n233 B.n132 10.6151
R1611 B.n234 B.n233 10.6151
R1612 B.n235 B.n234 10.6151
R1613 B.n235 B.n130 10.6151
R1614 B.n239 B.n130 10.6151
R1615 B.n240 B.n239 10.6151
R1616 B.n241 B.n240 10.6151
R1617 B.n241 B.n128 10.6151
R1618 B.n245 B.n128 10.6151
R1619 B.n246 B.n245 10.6151
R1620 B.n247 B.n246 10.6151
R1621 B.n247 B.n126 10.6151
R1622 B.n251 B.n126 10.6151
R1623 B.n252 B.n251 10.6151
R1624 B.n253 B.n252 10.6151
R1625 B.n253 B.n124 10.6151
R1626 B.n257 B.n124 10.6151
R1627 B.n260 B.n259 10.6151
R1628 B.n260 B.n120 10.6151
R1629 B.n264 B.n120 10.6151
R1630 B.n265 B.n264 10.6151
R1631 B.n266 B.n265 10.6151
R1632 B.n266 B.n118 10.6151
R1633 B.n270 B.n118 10.6151
R1634 B.n271 B.n270 10.6151
R1635 B.n272 B.n271 10.6151
R1636 B.n276 B.n275 10.6151
R1637 B.n277 B.n276 10.6151
R1638 B.n277 B.n112 10.6151
R1639 B.n281 B.n112 10.6151
R1640 B.n282 B.n281 10.6151
R1641 B.n283 B.n282 10.6151
R1642 B.n283 B.n110 10.6151
R1643 B.n287 B.n110 10.6151
R1644 B.n288 B.n287 10.6151
R1645 B.n289 B.n288 10.6151
R1646 B.n289 B.n108 10.6151
R1647 B.n293 B.n108 10.6151
R1648 B.n294 B.n293 10.6151
R1649 B.n295 B.n294 10.6151
R1650 B.n295 B.n106 10.6151
R1651 B.n299 B.n106 10.6151
R1652 B.n300 B.n299 10.6151
R1653 B.n301 B.n300 10.6151
R1654 B.n301 B.n104 10.6151
R1655 B.n305 B.n104 10.6151
R1656 B.n306 B.n305 10.6151
R1657 B.n307 B.n306 10.6151
R1658 B.n307 B.n102 10.6151
R1659 B.n311 B.n102 10.6151
R1660 B.n312 B.n311 10.6151
R1661 B.n313 B.n312 10.6151
R1662 B.n313 B.n100 10.6151
R1663 B.n317 B.n100 10.6151
R1664 B.n318 B.n317 10.6151
R1665 B.n319 B.n318 10.6151
R1666 B.n319 B.n98 10.6151
R1667 B.n323 B.n98 10.6151
R1668 B.n324 B.n323 10.6151
R1669 B.n325 B.n324 10.6151
R1670 B.n325 B.n96 10.6151
R1671 B.n329 B.n96 10.6151
R1672 B.n330 B.n329 10.6151
R1673 B.n331 B.n330 10.6151
R1674 B.n331 B.n94 10.6151
R1675 B.n335 B.n94 10.6151
R1676 B.n336 B.n335 10.6151
R1677 B.n337 B.n336 10.6151
R1678 B.n337 B.n92 10.6151
R1679 B.n341 B.n92 10.6151
R1680 B.n342 B.n341 10.6151
R1681 B.n343 B.n342 10.6151
R1682 B.n343 B.n90 10.6151
R1683 B.n347 B.n90 10.6151
R1684 B.n348 B.n347 10.6151
R1685 B.n349 B.n348 10.6151
R1686 B.n349 B.n88 10.6151
R1687 B.n353 B.n88 10.6151
R1688 B.n354 B.n353 10.6151
R1689 B.n175 B.n174 10.6151
R1690 B.n174 B.n173 10.6151
R1691 B.n173 B.n152 10.6151
R1692 B.n169 B.n152 10.6151
R1693 B.n169 B.n168 10.6151
R1694 B.n168 B.n167 10.6151
R1695 B.n167 B.n154 10.6151
R1696 B.n163 B.n154 10.6151
R1697 B.n163 B.n162 10.6151
R1698 B.n162 B.n161 10.6151
R1699 B.n161 B.n156 10.6151
R1700 B.n157 B.n156 10.6151
R1701 B.n157 B.n0 10.6151
R1702 B.n595 B.n1 10.6151
R1703 B.n595 B.n594 10.6151
R1704 B.n594 B.n593 10.6151
R1705 B.n593 B.n4 10.6151
R1706 B.n589 B.n4 10.6151
R1707 B.n589 B.n588 10.6151
R1708 B.n588 B.n587 10.6151
R1709 B.n587 B.n6 10.6151
R1710 B.n583 B.n6 10.6151
R1711 B.n583 B.n582 10.6151
R1712 B.n582 B.n581 10.6151
R1713 B.n581 B.n8 10.6151
R1714 B.n577 B.n8 10.6151
R1715 B.n497 B.n38 8.74196
R1716 B.n480 B.n479 8.74196
R1717 B.n258 B.n257 8.74196
R1718 B.n275 B.n116 8.74196
R1719 B.n599 B.n0 2.81026
R1720 B.n599 B.n1 2.81026
R1721 B.n494 B.n38 1.87367
R1722 B.n481 B.n480 1.87367
R1723 B.n259 B.n258 1.87367
R1724 B.n272 B.n116 1.87367
R1725 VN VN.t1 819.756
R1726 VN VN.t0 776.591
R1727 VDD2.n173 VDD2.n89 756.745
R1728 VDD2.n84 VDD2.n0 756.745
R1729 VDD2.n174 VDD2.n173 585
R1730 VDD2.n172 VDD2.n171 585
R1731 VDD2.n93 VDD2.n92 585
R1732 VDD2.n166 VDD2.n165 585
R1733 VDD2.n164 VDD2.n95 585
R1734 VDD2.n163 VDD2.n162 585
R1735 VDD2.n98 VDD2.n96 585
R1736 VDD2.n157 VDD2.n156 585
R1737 VDD2.n155 VDD2.n154 585
R1738 VDD2.n102 VDD2.n101 585
R1739 VDD2.n149 VDD2.n148 585
R1740 VDD2.n147 VDD2.n146 585
R1741 VDD2.n106 VDD2.n105 585
R1742 VDD2.n141 VDD2.n140 585
R1743 VDD2.n139 VDD2.n138 585
R1744 VDD2.n110 VDD2.n109 585
R1745 VDD2.n133 VDD2.n132 585
R1746 VDD2.n131 VDD2.n130 585
R1747 VDD2.n114 VDD2.n113 585
R1748 VDD2.n125 VDD2.n124 585
R1749 VDD2.n123 VDD2.n122 585
R1750 VDD2.n118 VDD2.n117 585
R1751 VDD2.n28 VDD2.n27 585
R1752 VDD2.n33 VDD2.n32 585
R1753 VDD2.n35 VDD2.n34 585
R1754 VDD2.n24 VDD2.n23 585
R1755 VDD2.n41 VDD2.n40 585
R1756 VDD2.n43 VDD2.n42 585
R1757 VDD2.n20 VDD2.n19 585
R1758 VDD2.n49 VDD2.n48 585
R1759 VDD2.n51 VDD2.n50 585
R1760 VDD2.n16 VDD2.n15 585
R1761 VDD2.n57 VDD2.n56 585
R1762 VDD2.n59 VDD2.n58 585
R1763 VDD2.n12 VDD2.n11 585
R1764 VDD2.n65 VDD2.n64 585
R1765 VDD2.n67 VDD2.n66 585
R1766 VDD2.n8 VDD2.n7 585
R1767 VDD2.n74 VDD2.n73 585
R1768 VDD2.n75 VDD2.n6 585
R1769 VDD2.n77 VDD2.n76 585
R1770 VDD2.n4 VDD2.n3 585
R1771 VDD2.n83 VDD2.n82 585
R1772 VDD2.n85 VDD2.n84 585
R1773 VDD2.n119 VDD2.t0 327.466
R1774 VDD2.n29 VDD2.t1 327.466
R1775 VDD2.n173 VDD2.n172 171.744
R1776 VDD2.n172 VDD2.n92 171.744
R1777 VDD2.n165 VDD2.n92 171.744
R1778 VDD2.n165 VDD2.n164 171.744
R1779 VDD2.n164 VDD2.n163 171.744
R1780 VDD2.n163 VDD2.n96 171.744
R1781 VDD2.n156 VDD2.n96 171.744
R1782 VDD2.n156 VDD2.n155 171.744
R1783 VDD2.n155 VDD2.n101 171.744
R1784 VDD2.n148 VDD2.n101 171.744
R1785 VDD2.n148 VDD2.n147 171.744
R1786 VDD2.n147 VDD2.n105 171.744
R1787 VDD2.n140 VDD2.n105 171.744
R1788 VDD2.n140 VDD2.n139 171.744
R1789 VDD2.n139 VDD2.n109 171.744
R1790 VDD2.n132 VDD2.n109 171.744
R1791 VDD2.n132 VDD2.n131 171.744
R1792 VDD2.n131 VDD2.n113 171.744
R1793 VDD2.n124 VDD2.n113 171.744
R1794 VDD2.n124 VDD2.n123 171.744
R1795 VDD2.n123 VDD2.n117 171.744
R1796 VDD2.n33 VDD2.n27 171.744
R1797 VDD2.n34 VDD2.n33 171.744
R1798 VDD2.n34 VDD2.n23 171.744
R1799 VDD2.n41 VDD2.n23 171.744
R1800 VDD2.n42 VDD2.n41 171.744
R1801 VDD2.n42 VDD2.n19 171.744
R1802 VDD2.n49 VDD2.n19 171.744
R1803 VDD2.n50 VDD2.n49 171.744
R1804 VDD2.n50 VDD2.n15 171.744
R1805 VDD2.n57 VDD2.n15 171.744
R1806 VDD2.n58 VDD2.n57 171.744
R1807 VDD2.n58 VDD2.n11 171.744
R1808 VDD2.n65 VDD2.n11 171.744
R1809 VDD2.n66 VDD2.n65 171.744
R1810 VDD2.n66 VDD2.n7 171.744
R1811 VDD2.n74 VDD2.n7 171.744
R1812 VDD2.n75 VDD2.n74 171.744
R1813 VDD2.n76 VDD2.n75 171.744
R1814 VDD2.n76 VDD2.n3 171.744
R1815 VDD2.n83 VDD2.n3 171.744
R1816 VDD2.n84 VDD2.n83 171.744
R1817 VDD2.n178 VDD2.n88 91.2172
R1818 VDD2.t0 VDD2.n117 85.8723
R1819 VDD2.t1 VDD2.n27 85.8723
R1820 VDD2.n178 VDD2.n177 51.7732
R1821 VDD2.n119 VDD2.n118 16.3895
R1822 VDD2.n29 VDD2.n28 16.3895
R1823 VDD2.n166 VDD2.n95 13.1884
R1824 VDD2.n77 VDD2.n6 13.1884
R1825 VDD2.n167 VDD2.n93 12.8005
R1826 VDD2.n162 VDD2.n97 12.8005
R1827 VDD2.n122 VDD2.n121 12.8005
R1828 VDD2.n32 VDD2.n31 12.8005
R1829 VDD2.n73 VDD2.n72 12.8005
R1830 VDD2.n78 VDD2.n4 12.8005
R1831 VDD2.n171 VDD2.n170 12.0247
R1832 VDD2.n161 VDD2.n98 12.0247
R1833 VDD2.n125 VDD2.n116 12.0247
R1834 VDD2.n35 VDD2.n26 12.0247
R1835 VDD2.n71 VDD2.n8 12.0247
R1836 VDD2.n82 VDD2.n81 12.0247
R1837 VDD2.n174 VDD2.n91 11.249
R1838 VDD2.n158 VDD2.n157 11.249
R1839 VDD2.n126 VDD2.n114 11.249
R1840 VDD2.n36 VDD2.n24 11.249
R1841 VDD2.n68 VDD2.n67 11.249
R1842 VDD2.n85 VDD2.n2 11.249
R1843 VDD2.n175 VDD2.n89 10.4732
R1844 VDD2.n154 VDD2.n100 10.4732
R1845 VDD2.n130 VDD2.n129 10.4732
R1846 VDD2.n40 VDD2.n39 10.4732
R1847 VDD2.n64 VDD2.n10 10.4732
R1848 VDD2.n86 VDD2.n0 10.4732
R1849 VDD2.n153 VDD2.n102 9.69747
R1850 VDD2.n133 VDD2.n112 9.69747
R1851 VDD2.n43 VDD2.n22 9.69747
R1852 VDD2.n63 VDD2.n12 9.69747
R1853 VDD2.n177 VDD2.n176 9.45567
R1854 VDD2.n88 VDD2.n87 9.45567
R1855 VDD2.n145 VDD2.n144 9.3005
R1856 VDD2.n104 VDD2.n103 9.3005
R1857 VDD2.n151 VDD2.n150 9.3005
R1858 VDD2.n153 VDD2.n152 9.3005
R1859 VDD2.n100 VDD2.n99 9.3005
R1860 VDD2.n159 VDD2.n158 9.3005
R1861 VDD2.n161 VDD2.n160 9.3005
R1862 VDD2.n97 VDD2.n94 9.3005
R1863 VDD2.n176 VDD2.n175 9.3005
R1864 VDD2.n91 VDD2.n90 9.3005
R1865 VDD2.n170 VDD2.n169 9.3005
R1866 VDD2.n168 VDD2.n167 9.3005
R1867 VDD2.n143 VDD2.n142 9.3005
R1868 VDD2.n108 VDD2.n107 9.3005
R1869 VDD2.n137 VDD2.n136 9.3005
R1870 VDD2.n135 VDD2.n134 9.3005
R1871 VDD2.n112 VDD2.n111 9.3005
R1872 VDD2.n129 VDD2.n128 9.3005
R1873 VDD2.n127 VDD2.n126 9.3005
R1874 VDD2.n116 VDD2.n115 9.3005
R1875 VDD2.n121 VDD2.n120 9.3005
R1876 VDD2.n87 VDD2.n86 9.3005
R1877 VDD2.n2 VDD2.n1 9.3005
R1878 VDD2.n81 VDD2.n80 9.3005
R1879 VDD2.n79 VDD2.n78 9.3005
R1880 VDD2.n18 VDD2.n17 9.3005
R1881 VDD2.n47 VDD2.n46 9.3005
R1882 VDD2.n45 VDD2.n44 9.3005
R1883 VDD2.n22 VDD2.n21 9.3005
R1884 VDD2.n39 VDD2.n38 9.3005
R1885 VDD2.n37 VDD2.n36 9.3005
R1886 VDD2.n26 VDD2.n25 9.3005
R1887 VDD2.n31 VDD2.n30 9.3005
R1888 VDD2.n53 VDD2.n52 9.3005
R1889 VDD2.n55 VDD2.n54 9.3005
R1890 VDD2.n14 VDD2.n13 9.3005
R1891 VDD2.n61 VDD2.n60 9.3005
R1892 VDD2.n63 VDD2.n62 9.3005
R1893 VDD2.n10 VDD2.n9 9.3005
R1894 VDD2.n69 VDD2.n68 9.3005
R1895 VDD2.n71 VDD2.n70 9.3005
R1896 VDD2.n72 VDD2.n5 9.3005
R1897 VDD2.n150 VDD2.n149 8.92171
R1898 VDD2.n134 VDD2.n110 8.92171
R1899 VDD2.n44 VDD2.n20 8.92171
R1900 VDD2.n60 VDD2.n59 8.92171
R1901 VDD2.n146 VDD2.n104 8.14595
R1902 VDD2.n138 VDD2.n137 8.14595
R1903 VDD2.n48 VDD2.n47 8.14595
R1904 VDD2.n56 VDD2.n14 8.14595
R1905 VDD2.n145 VDD2.n106 7.3702
R1906 VDD2.n141 VDD2.n108 7.3702
R1907 VDD2.n51 VDD2.n18 7.3702
R1908 VDD2.n55 VDD2.n16 7.3702
R1909 VDD2.n142 VDD2.n106 6.59444
R1910 VDD2.n142 VDD2.n141 6.59444
R1911 VDD2.n52 VDD2.n51 6.59444
R1912 VDD2.n52 VDD2.n16 6.59444
R1913 VDD2.n146 VDD2.n145 5.81868
R1914 VDD2.n138 VDD2.n108 5.81868
R1915 VDD2.n48 VDD2.n18 5.81868
R1916 VDD2.n56 VDD2.n55 5.81868
R1917 VDD2.n149 VDD2.n104 5.04292
R1918 VDD2.n137 VDD2.n110 5.04292
R1919 VDD2.n47 VDD2.n20 5.04292
R1920 VDD2.n59 VDD2.n14 5.04292
R1921 VDD2.n150 VDD2.n102 4.26717
R1922 VDD2.n134 VDD2.n133 4.26717
R1923 VDD2.n44 VDD2.n43 4.26717
R1924 VDD2.n60 VDD2.n12 4.26717
R1925 VDD2.n120 VDD2.n119 3.70982
R1926 VDD2.n30 VDD2.n29 3.70982
R1927 VDD2.n177 VDD2.n89 3.49141
R1928 VDD2.n154 VDD2.n153 3.49141
R1929 VDD2.n130 VDD2.n112 3.49141
R1930 VDD2.n40 VDD2.n22 3.49141
R1931 VDD2.n64 VDD2.n63 3.49141
R1932 VDD2.n88 VDD2.n0 3.49141
R1933 VDD2.n175 VDD2.n174 2.71565
R1934 VDD2.n157 VDD2.n100 2.71565
R1935 VDD2.n129 VDD2.n114 2.71565
R1936 VDD2.n39 VDD2.n24 2.71565
R1937 VDD2.n67 VDD2.n10 2.71565
R1938 VDD2.n86 VDD2.n85 2.71565
R1939 VDD2.n171 VDD2.n91 1.93989
R1940 VDD2.n158 VDD2.n98 1.93989
R1941 VDD2.n126 VDD2.n125 1.93989
R1942 VDD2.n36 VDD2.n35 1.93989
R1943 VDD2.n68 VDD2.n8 1.93989
R1944 VDD2.n82 VDD2.n2 1.93989
R1945 VDD2.n170 VDD2.n93 1.16414
R1946 VDD2.n162 VDD2.n161 1.16414
R1947 VDD2.n122 VDD2.n116 1.16414
R1948 VDD2.n32 VDD2.n26 1.16414
R1949 VDD2.n73 VDD2.n71 1.16414
R1950 VDD2.n81 VDD2.n4 1.16414
R1951 VDD2.n167 VDD2.n166 0.388379
R1952 VDD2.n97 VDD2.n95 0.388379
R1953 VDD2.n121 VDD2.n118 0.388379
R1954 VDD2.n31 VDD2.n28 0.388379
R1955 VDD2.n72 VDD2.n6 0.388379
R1956 VDD2.n78 VDD2.n77 0.388379
R1957 VDD2 VDD2.n178 0.280672
R1958 VDD2.n176 VDD2.n90 0.155672
R1959 VDD2.n169 VDD2.n90 0.155672
R1960 VDD2.n169 VDD2.n168 0.155672
R1961 VDD2.n168 VDD2.n94 0.155672
R1962 VDD2.n160 VDD2.n94 0.155672
R1963 VDD2.n160 VDD2.n159 0.155672
R1964 VDD2.n159 VDD2.n99 0.155672
R1965 VDD2.n152 VDD2.n99 0.155672
R1966 VDD2.n152 VDD2.n151 0.155672
R1967 VDD2.n151 VDD2.n103 0.155672
R1968 VDD2.n144 VDD2.n103 0.155672
R1969 VDD2.n144 VDD2.n143 0.155672
R1970 VDD2.n143 VDD2.n107 0.155672
R1971 VDD2.n136 VDD2.n107 0.155672
R1972 VDD2.n136 VDD2.n135 0.155672
R1973 VDD2.n135 VDD2.n111 0.155672
R1974 VDD2.n128 VDD2.n111 0.155672
R1975 VDD2.n128 VDD2.n127 0.155672
R1976 VDD2.n127 VDD2.n115 0.155672
R1977 VDD2.n120 VDD2.n115 0.155672
R1978 VDD2.n30 VDD2.n25 0.155672
R1979 VDD2.n37 VDD2.n25 0.155672
R1980 VDD2.n38 VDD2.n37 0.155672
R1981 VDD2.n38 VDD2.n21 0.155672
R1982 VDD2.n45 VDD2.n21 0.155672
R1983 VDD2.n46 VDD2.n45 0.155672
R1984 VDD2.n46 VDD2.n17 0.155672
R1985 VDD2.n53 VDD2.n17 0.155672
R1986 VDD2.n54 VDD2.n53 0.155672
R1987 VDD2.n54 VDD2.n13 0.155672
R1988 VDD2.n61 VDD2.n13 0.155672
R1989 VDD2.n62 VDD2.n61 0.155672
R1990 VDD2.n62 VDD2.n9 0.155672
R1991 VDD2.n69 VDD2.n9 0.155672
R1992 VDD2.n70 VDD2.n69 0.155672
R1993 VDD2.n70 VDD2.n5 0.155672
R1994 VDD2.n79 VDD2.n5 0.155672
R1995 VDD2.n80 VDD2.n79 0.155672
R1996 VDD2.n80 VDD2.n1 0.155672
R1997 VDD2.n87 VDD2.n1 0.155672
C0 B VDD1 1.72333f
C1 B w_n1382_n4218# 7.94573f
C2 VP VN 5.3451f
C3 VP VDD2 0.255642f
C4 VN VDD2 2.60324f
C5 VP VTAIL 1.92239f
C6 VN VTAIL 1.90761f
C7 VTAIL VDD2 7.24671f
C8 VP B 1.05217f
C9 VN B 0.777109f
C10 B VDD2 1.73783f
C11 B VTAIL 3.50998f
C12 VDD1 w_n1382_n4218# 1.88404f
C13 VP VDD1 2.70448f
C14 VP w_n1382_n4218# 1.99837f
C15 VN VDD1 0.148589f
C16 VN w_n1382_n4218# 1.82643f
C17 VDD2 VDD1 0.463311f
C18 VDD2 w_n1382_n4218# 1.88869f
C19 VTAIL VDD1 7.21522f
C20 VTAIL w_n1382_n4218# 3.60845f
C21 VDD2 VSUBS 0.890893f
C22 VDD1 VSUBS 3.712862f
C23 VTAIL VSUBS 0.9031f
C24 VN VSUBS 6.45709f
C25 VP VSUBS 1.266088f
C26 B VSUBS 2.854248f
C27 w_n1382_n4218# VSUBS 71.394104f
C28 VDD2.n0 VSUBS 0.023014f
C29 VDD2.n1 VSUBS 0.020783f
C30 VDD2.n2 VSUBS 0.011168f
C31 VDD2.n3 VSUBS 0.026397f
C32 VDD2.n4 VSUBS 0.011825f
C33 VDD2.n5 VSUBS 0.020783f
C34 VDD2.n6 VSUBS 0.011496f
C35 VDD2.n7 VSUBS 0.026397f
C36 VDD2.n8 VSUBS 0.011825f
C37 VDD2.n9 VSUBS 0.020783f
C38 VDD2.n10 VSUBS 0.011168f
C39 VDD2.n11 VSUBS 0.026397f
C40 VDD2.n12 VSUBS 0.011825f
C41 VDD2.n13 VSUBS 0.020783f
C42 VDD2.n14 VSUBS 0.011168f
C43 VDD2.n15 VSUBS 0.026397f
C44 VDD2.n16 VSUBS 0.011825f
C45 VDD2.n17 VSUBS 0.020783f
C46 VDD2.n18 VSUBS 0.011168f
C47 VDD2.n19 VSUBS 0.026397f
C48 VDD2.n20 VSUBS 0.011825f
C49 VDD2.n21 VSUBS 0.020783f
C50 VDD2.n22 VSUBS 0.011168f
C51 VDD2.n23 VSUBS 0.026397f
C52 VDD2.n24 VSUBS 0.011825f
C53 VDD2.n25 VSUBS 0.020783f
C54 VDD2.n26 VSUBS 0.011168f
C55 VDD2.n27 VSUBS 0.019798f
C56 VDD2.n28 VSUBS 0.016792f
C57 VDD2.t1 VSUBS 0.056574f
C58 VDD2.n29 VSUBS 0.154042f
C59 VDD2.n30 VSUBS 1.44309f
C60 VDD2.n31 VSUBS 0.011168f
C61 VDD2.n32 VSUBS 0.011825f
C62 VDD2.n33 VSUBS 0.026397f
C63 VDD2.n34 VSUBS 0.026397f
C64 VDD2.n35 VSUBS 0.011825f
C65 VDD2.n36 VSUBS 0.011168f
C66 VDD2.n37 VSUBS 0.020783f
C67 VDD2.n38 VSUBS 0.020783f
C68 VDD2.n39 VSUBS 0.011168f
C69 VDD2.n40 VSUBS 0.011825f
C70 VDD2.n41 VSUBS 0.026397f
C71 VDD2.n42 VSUBS 0.026397f
C72 VDD2.n43 VSUBS 0.011825f
C73 VDD2.n44 VSUBS 0.011168f
C74 VDD2.n45 VSUBS 0.020783f
C75 VDD2.n46 VSUBS 0.020783f
C76 VDD2.n47 VSUBS 0.011168f
C77 VDD2.n48 VSUBS 0.011825f
C78 VDD2.n49 VSUBS 0.026397f
C79 VDD2.n50 VSUBS 0.026397f
C80 VDD2.n51 VSUBS 0.011825f
C81 VDD2.n52 VSUBS 0.011168f
C82 VDD2.n53 VSUBS 0.020783f
C83 VDD2.n54 VSUBS 0.020783f
C84 VDD2.n55 VSUBS 0.011168f
C85 VDD2.n56 VSUBS 0.011825f
C86 VDD2.n57 VSUBS 0.026397f
C87 VDD2.n58 VSUBS 0.026397f
C88 VDD2.n59 VSUBS 0.011825f
C89 VDD2.n60 VSUBS 0.011168f
C90 VDD2.n61 VSUBS 0.020783f
C91 VDD2.n62 VSUBS 0.020783f
C92 VDD2.n63 VSUBS 0.011168f
C93 VDD2.n64 VSUBS 0.011825f
C94 VDD2.n65 VSUBS 0.026397f
C95 VDD2.n66 VSUBS 0.026397f
C96 VDD2.n67 VSUBS 0.011825f
C97 VDD2.n68 VSUBS 0.011168f
C98 VDD2.n69 VSUBS 0.020783f
C99 VDD2.n70 VSUBS 0.020783f
C100 VDD2.n71 VSUBS 0.011168f
C101 VDD2.n72 VSUBS 0.011168f
C102 VDD2.n73 VSUBS 0.011825f
C103 VDD2.n74 VSUBS 0.026397f
C104 VDD2.n75 VSUBS 0.026397f
C105 VDD2.n76 VSUBS 0.026397f
C106 VDD2.n77 VSUBS 0.011496f
C107 VDD2.n78 VSUBS 0.011168f
C108 VDD2.n79 VSUBS 0.020783f
C109 VDD2.n80 VSUBS 0.020783f
C110 VDD2.n81 VSUBS 0.011168f
C111 VDD2.n82 VSUBS 0.011825f
C112 VDD2.n83 VSUBS 0.026397f
C113 VDD2.n84 VSUBS 0.064508f
C114 VDD2.n85 VSUBS 0.011825f
C115 VDD2.n86 VSUBS 0.011168f
C116 VDD2.n87 VSUBS 0.052298f
C117 VDD2.n88 VSUBS 0.616217f
C118 VDD2.n89 VSUBS 0.023014f
C119 VDD2.n90 VSUBS 0.020783f
C120 VDD2.n91 VSUBS 0.011168f
C121 VDD2.n92 VSUBS 0.026397f
C122 VDD2.n93 VSUBS 0.011825f
C123 VDD2.n94 VSUBS 0.020783f
C124 VDD2.n95 VSUBS 0.011496f
C125 VDD2.n96 VSUBS 0.026397f
C126 VDD2.n97 VSUBS 0.011168f
C127 VDD2.n98 VSUBS 0.011825f
C128 VDD2.n99 VSUBS 0.020783f
C129 VDD2.n100 VSUBS 0.011168f
C130 VDD2.n101 VSUBS 0.026397f
C131 VDD2.n102 VSUBS 0.011825f
C132 VDD2.n103 VSUBS 0.020783f
C133 VDD2.n104 VSUBS 0.011168f
C134 VDD2.n105 VSUBS 0.026397f
C135 VDD2.n106 VSUBS 0.011825f
C136 VDD2.n107 VSUBS 0.020783f
C137 VDD2.n108 VSUBS 0.011168f
C138 VDD2.n109 VSUBS 0.026397f
C139 VDD2.n110 VSUBS 0.011825f
C140 VDD2.n111 VSUBS 0.020783f
C141 VDD2.n112 VSUBS 0.011168f
C142 VDD2.n113 VSUBS 0.026397f
C143 VDD2.n114 VSUBS 0.011825f
C144 VDD2.n115 VSUBS 0.020783f
C145 VDD2.n116 VSUBS 0.011168f
C146 VDD2.n117 VSUBS 0.019798f
C147 VDD2.n118 VSUBS 0.016792f
C148 VDD2.t0 VSUBS 0.056574f
C149 VDD2.n119 VSUBS 0.154042f
C150 VDD2.n120 VSUBS 1.44309f
C151 VDD2.n121 VSUBS 0.011168f
C152 VDD2.n122 VSUBS 0.011825f
C153 VDD2.n123 VSUBS 0.026397f
C154 VDD2.n124 VSUBS 0.026397f
C155 VDD2.n125 VSUBS 0.011825f
C156 VDD2.n126 VSUBS 0.011168f
C157 VDD2.n127 VSUBS 0.020783f
C158 VDD2.n128 VSUBS 0.020783f
C159 VDD2.n129 VSUBS 0.011168f
C160 VDD2.n130 VSUBS 0.011825f
C161 VDD2.n131 VSUBS 0.026397f
C162 VDD2.n132 VSUBS 0.026397f
C163 VDD2.n133 VSUBS 0.011825f
C164 VDD2.n134 VSUBS 0.011168f
C165 VDD2.n135 VSUBS 0.020783f
C166 VDD2.n136 VSUBS 0.020783f
C167 VDD2.n137 VSUBS 0.011168f
C168 VDD2.n138 VSUBS 0.011825f
C169 VDD2.n139 VSUBS 0.026397f
C170 VDD2.n140 VSUBS 0.026397f
C171 VDD2.n141 VSUBS 0.011825f
C172 VDD2.n142 VSUBS 0.011168f
C173 VDD2.n143 VSUBS 0.020783f
C174 VDD2.n144 VSUBS 0.020783f
C175 VDD2.n145 VSUBS 0.011168f
C176 VDD2.n146 VSUBS 0.011825f
C177 VDD2.n147 VSUBS 0.026397f
C178 VDD2.n148 VSUBS 0.026397f
C179 VDD2.n149 VSUBS 0.011825f
C180 VDD2.n150 VSUBS 0.011168f
C181 VDD2.n151 VSUBS 0.020783f
C182 VDD2.n152 VSUBS 0.020783f
C183 VDD2.n153 VSUBS 0.011168f
C184 VDD2.n154 VSUBS 0.011825f
C185 VDD2.n155 VSUBS 0.026397f
C186 VDD2.n156 VSUBS 0.026397f
C187 VDD2.n157 VSUBS 0.011825f
C188 VDD2.n158 VSUBS 0.011168f
C189 VDD2.n159 VSUBS 0.020783f
C190 VDD2.n160 VSUBS 0.020783f
C191 VDD2.n161 VSUBS 0.011168f
C192 VDD2.n162 VSUBS 0.011825f
C193 VDD2.n163 VSUBS 0.026397f
C194 VDD2.n164 VSUBS 0.026397f
C195 VDD2.n165 VSUBS 0.026397f
C196 VDD2.n166 VSUBS 0.011496f
C197 VDD2.n167 VSUBS 0.011168f
C198 VDD2.n168 VSUBS 0.020783f
C199 VDD2.n169 VSUBS 0.020783f
C200 VDD2.n170 VSUBS 0.011168f
C201 VDD2.n171 VSUBS 0.011825f
C202 VDD2.n172 VSUBS 0.026397f
C203 VDD2.n173 VSUBS 0.064508f
C204 VDD2.n174 VSUBS 0.011825f
C205 VDD2.n175 VSUBS 0.011168f
C206 VDD2.n176 VSUBS 0.052298f
C207 VDD2.n177 VSUBS 0.046913f
C208 VDD2.n178 VSUBS 2.61757f
C209 VN.t0 VSUBS 1.55597f
C210 VN.t1 VSUBS 1.68105f
C211 B.n0 VSUBS 0.00439f
C212 B.n1 VSUBS 0.00439f
C213 B.n2 VSUBS 0.006943f
C214 B.n3 VSUBS 0.006943f
C215 B.n4 VSUBS 0.006943f
C216 B.n5 VSUBS 0.006943f
C217 B.n6 VSUBS 0.006943f
C218 B.n7 VSUBS 0.006943f
C219 B.n8 VSUBS 0.006943f
C220 B.n9 VSUBS 0.016998f
C221 B.n10 VSUBS 0.006943f
C222 B.n11 VSUBS 0.006943f
C223 B.n12 VSUBS 0.006943f
C224 B.n13 VSUBS 0.006943f
C225 B.n14 VSUBS 0.006943f
C226 B.n15 VSUBS 0.006943f
C227 B.n16 VSUBS 0.006943f
C228 B.n17 VSUBS 0.006943f
C229 B.n18 VSUBS 0.006943f
C230 B.n19 VSUBS 0.006943f
C231 B.n20 VSUBS 0.006943f
C232 B.n21 VSUBS 0.006943f
C233 B.n22 VSUBS 0.006943f
C234 B.n23 VSUBS 0.006943f
C235 B.n24 VSUBS 0.006943f
C236 B.n25 VSUBS 0.006943f
C237 B.n26 VSUBS 0.006943f
C238 B.n27 VSUBS 0.006943f
C239 B.n28 VSUBS 0.006943f
C240 B.n29 VSUBS 0.006943f
C241 B.n30 VSUBS 0.006943f
C242 B.n31 VSUBS 0.006943f
C243 B.n32 VSUBS 0.006943f
C244 B.n33 VSUBS 0.006943f
C245 B.n34 VSUBS 0.006943f
C246 B.n35 VSUBS 0.006943f
C247 B.t8 VSUBS 0.306222f
C248 B.t7 VSUBS 0.318364f
C249 B.t6 VSUBS 0.456695f
C250 B.n36 VSUBS 0.397702f
C251 B.n37 VSUBS 0.296727f
C252 B.n38 VSUBS 0.016086f
C253 B.n39 VSUBS 0.006943f
C254 B.n40 VSUBS 0.006943f
C255 B.n41 VSUBS 0.006943f
C256 B.n42 VSUBS 0.006943f
C257 B.n43 VSUBS 0.006943f
C258 B.t2 VSUBS 0.306226f
C259 B.t1 VSUBS 0.318367f
C260 B.t0 VSUBS 0.456695f
C261 B.n44 VSUBS 0.397699f
C262 B.n45 VSUBS 0.296724f
C263 B.n46 VSUBS 0.006943f
C264 B.n47 VSUBS 0.006943f
C265 B.n48 VSUBS 0.006943f
C266 B.n49 VSUBS 0.006943f
C267 B.n50 VSUBS 0.006943f
C268 B.n51 VSUBS 0.006943f
C269 B.n52 VSUBS 0.006943f
C270 B.n53 VSUBS 0.006943f
C271 B.n54 VSUBS 0.006943f
C272 B.n55 VSUBS 0.006943f
C273 B.n56 VSUBS 0.006943f
C274 B.n57 VSUBS 0.006943f
C275 B.n58 VSUBS 0.006943f
C276 B.n59 VSUBS 0.006943f
C277 B.n60 VSUBS 0.006943f
C278 B.n61 VSUBS 0.006943f
C279 B.n62 VSUBS 0.006943f
C280 B.n63 VSUBS 0.006943f
C281 B.n64 VSUBS 0.006943f
C282 B.n65 VSUBS 0.006943f
C283 B.n66 VSUBS 0.006943f
C284 B.n67 VSUBS 0.006943f
C285 B.n68 VSUBS 0.006943f
C286 B.n69 VSUBS 0.006943f
C287 B.n70 VSUBS 0.006943f
C288 B.n71 VSUBS 0.006943f
C289 B.n72 VSUBS 0.016192f
C290 B.n73 VSUBS 0.006943f
C291 B.n74 VSUBS 0.006943f
C292 B.n75 VSUBS 0.006943f
C293 B.n76 VSUBS 0.006943f
C294 B.n77 VSUBS 0.006943f
C295 B.n78 VSUBS 0.006943f
C296 B.n79 VSUBS 0.006943f
C297 B.n80 VSUBS 0.006943f
C298 B.n81 VSUBS 0.006943f
C299 B.n82 VSUBS 0.006943f
C300 B.n83 VSUBS 0.006943f
C301 B.n84 VSUBS 0.006943f
C302 B.n85 VSUBS 0.006943f
C303 B.n86 VSUBS 0.006943f
C304 B.n87 VSUBS 0.016998f
C305 B.n88 VSUBS 0.006943f
C306 B.n89 VSUBS 0.006943f
C307 B.n90 VSUBS 0.006943f
C308 B.n91 VSUBS 0.006943f
C309 B.n92 VSUBS 0.006943f
C310 B.n93 VSUBS 0.006943f
C311 B.n94 VSUBS 0.006943f
C312 B.n95 VSUBS 0.006943f
C313 B.n96 VSUBS 0.006943f
C314 B.n97 VSUBS 0.006943f
C315 B.n98 VSUBS 0.006943f
C316 B.n99 VSUBS 0.006943f
C317 B.n100 VSUBS 0.006943f
C318 B.n101 VSUBS 0.006943f
C319 B.n102 VSUBS 0.006943f
C320 B.n103 VSUBS 0.006943f
C321 B.n104 VSUBS 0.006943f
C322 B.n105 VSUBS 0.006943f
C323 B.n106 VSUBS 0.006943f
C324 B.n107 VSUBS 0.006943f
C325 B.n108 VSUBS 0.006943f
C326 B.n109 VSUBS 0.006943f
C327 B.n110 VSUBS 0.006943f
C328 B.n111 VSUBS 0.006943f
C329 B.n112 VSUBS 0.006943f
C330 B.n113 VSUBS 0.006943f
C331 B.t10 VSUBS 0.306226f
C332 B.t11 VSUBS 0.318367f
C333 B.t9 VSUBS 0.456695f
C334 B.n114 VSUBS 0.397699f
C335 B.n115 VSUBS 0.296724f
C336 B.n116 VSUBS 0.016086f
C337 B.n117 VSUBS 0.006943f
C338 B.n118 VSUBS 0.006943f
C339 B.n119 VSUBS 0.006943f
C340 B.n120 VSUBS 0.006943f
C341 B.n121 VSUBS 0.006943f
C342 B.t4 VSUBS 0.306222f
C343 B.t5 VSUBS 0.318364f
C344 B.t3 VSUBS 0.456695f
C345 B.n122 VSUBS 0.397702f
C346 B.n123 VSUBS 0.296727f
C347 B.n124 VSUBS 0.006943f
C348 B.n125 VSUBS 0.006943f
C349 B.n126 VSUBS 0.006943f
C350 B.n127 VSUBS 0.006943f
C351 B.n128 VSUBS 0.006943f
C352 B.n129 VSUBS 0.006943f
C353 B.n130 VSUBS 0.006943f
C354 B.n131 VSUBS 0.006943f
C355 B.n132 VSUBS 0.006943f
C356 B.n133 VSUBS 0.006943f
C357 B.n134 VSUBS 0.006943f
C358 B.n135 VSUBS 0.006943f
C359 B.n136 VSUBS 0.006943f
C360 B.n137 VSUBS 0.006943f
C361 B.n138 VSUBS 0.006943f
C362 B.n139 VSUBS 0.006943f
C363 B.n140 VSUBS 0.006943f
C364 B.n141 VSUBS 0.006943f
C365 B.n142 VSUBS 0.006943f
C366 B.n143 VSUBS 0.006943f
C367 B.n144 VSUBS 0.006943f
C368 B.n145 VSUBS 0.006943f
C369 B.n146 VSUBS 0.006943f
C370 B.n147 VSUBS 0.006943f
C371 B.n148 VSUBS 0.006943f
C372 B.n149 VSUBS 0.006943f
C373 B.n150 VSUBS 0.016998f
C374 B.n151 VSUBS 0.006943f
C375 B.n152 VSUBS 0.006943f
C376 B.n153 VSUBS 0.006943f
C377 B.n154 VSUBS 0.006943f
C378 B.n155 VSUBS 0.006943f
C379 B.n156 VSUBS 0.006943f
C380 B.n157 VSUBS 0.006943f
C381 B.n158 VSUBS 0.006943f
C382 B.n159 VSUBS 0.006943f
C383 B.n160 VSUBS 0.006943f
C384 B.n161 VSUBS 0.006943f
C385 B.n162 VSUBS 0.006943f
C386 B.n163 VSUBS 0.006943f
C387 B.n164 VSUBS 0.006943f
C388 B.n165 VSUBS 0.006943f
C389 B.n166 VSUBS 0.006943f
C390 B.n167 VSUBS 0.006943f
C391 B.n168 VSUBS 0.006943f
C392 B.n169 VSUBS 0.006943f
C393 B.n170 VSUBS 0.006943f
C394 B.n171 VSUBS 0.006943f
C395 B.n172 VSUBS 0.006943f
C396 B.n173 VSUBS 0.006943f
C397 B.n174 VSUBS 0.006943f
C398 B.n175 VSUBS 0.015878f
C399 B.n176 VSUBS 0.015878f
C400 B.n177 VSUBS 0.016998f
C401 B.n178 VSUBS 0.006943f
C402 B.n179 VSUBS 0.006943f
C403 B.n180 VSUBS 0.006943f
C404 B.n181 VSUBS 0.006943f
C405 B.n182 VSUBS 0.006943f
C406 B.n183 VSUBS 0.006943f
C407 B.n184 VSUBS 0.006943f
C408 B.n185 VSUBS 0.006943f
C409 B.n186 VSUBS 0.006943f
C410 B.n187 VSUBS 0.006943f
C411 B.n188 VSUBS 0.006943f
C412 B.n189 VSUBS 0.006943f
C413 B.n190 VSUBS 0.006943f
C414 B.n191 VSUBS 0.006943f
C415 B.n192 VSUBS 0.006943f
C416 B.n193 VSUBS 0.006943f
C417 B.n194 VSUBS 0.006943f
C418 B.n195 VSUBS 0.006943f
C419 B.n196 VSUBS 0.006943f
C420 B.n197 VSUBS 0.006943f
C421 B.n198 VSUBS 0.006943f
C422 B.n199 VSUBS 0.006943f
C423 B.n200 VSUBS 0.006943f
C424 B.n201 VSUBS 0.006943f
C425 B.n202 VSUBS 0.006943f
C426 B.n203 VSUBS 0.006943f
C427 B.n204 VSUBS 0.006943f
C428 B.n205 VSUBS 0.006943f
C429 B.n206 VSUBS 0.006943f
C430 B.n207 VSUBS 0.006943f
C431 B.n208 VSUBS 0.006943f
C432 B.n209 VSUBS 0.006943f
C433 B.n210 VSUBS 0.006943f
C434 B.n211 VSUBS 0.006943f
C435 B.n212 VSUBS 0.006943f
C436 B.n213 VSUBS 0.006943f
C437 B.n214 VSUBS 0.006943f
C438 B.n215 VSUBS 0.006943f
C439 B.n216 VSUBS 0.006943f
C440 B.n217 VSUBS 0.006943f
C441 B.n218 VSUBS 0.006943f
C442 B.n219 VSUBS 0.006943f
C443 B.n220 VSUBS 0.006943f
C444 B.n221 VSUBS 0.006943f
C445 B.n222 VSUBS 0.006943f
C446 B.n223 VSUBS 0.006943f
C447 B.n224 VSUBS 0.006943f
C448 B.n225 VSUBS 0.006943f
C449 B.n226 VSUBS 0.006943f
C450 B.n227 VSUBS 0.006943f
C451 B.n228 VSUBS 0.006943f
C452 B.n229 VSUBS 0.006943f
C453 B.n230 VSUBS 0.006943f
C454 B.n231 VSUBS 0.006943f
C455 B.n232 VSUBS 0.006943f
C456 B.n233 VSUBS 0.006943f
C457 B.n234 VSUBS 0.006943f
C458 B.n235 VSUBS 0.006943f
C459 B.n236 VSUBS 0.006943f
C460 B.n237 VSUBS 0.006943f
C461 B.n238 VSUBS 0.006943f
C462 B.n239 VSUBS 0.006943f
C463 B.n240 VSUBS 0.006943f
C464 B.n241 VSUBS 0.006943f
C465 B.n242 VSUBS 0.006943f
C466 B.n243 VSUBS 0.006943f
C467 B.n244 VSUBS 0.006943f
C468 B.n245 VSUBS 0.006943f
C469 B.n246 VSUBS 0.006943f
C470 B.n247 VSUBS 0.006943f
C471 B.n248 VSUBS 0.006943f
C472 B.n249 VSUBS 0.006943f
C473 B.n250 VSUBS 0.006943f
C474 B.n251 VSUBS 0.006943f
C475 B.n252 VSUBS 0.006943f
C476 B.n253 VSUBS 0.006943f
C477 B.n254 VSUBS 0.006943f
C478 B.n255 VSUBS 0.006943f
C479 B.n256 VSUBS 0.006943f
C480 B.n257 VSUBS 0.00633f
C481 B.n258 VSUBS 0.016086f
C482 B.n259 VSUBS 0.004084f
C483 B.n260 VSUBS 0.006943f
C484 B.n261 VSUBS 0.006943f
C485 B.n262 VSUBS 0.006943f
C486 B.n263 VSUBS 0.006943f
C487 B.n264 VSUBS 0.006943f
C488 B.n265 VSUBS 0.006943f
C489 B.n266 VSUBS 0.006943f
C490 B.n267 VSUBS 0.006943f
C491 B.n268 VSUBS 0.006943f
C492 B.n269 VSUBS 0.006943f
C493 B.n270 VSUBS 0.006943f
C494 B.n271 VSUBS 0.006943f
C495 B.n272 VSUBS 0.004084f
C496 B.n273 VSUBS 0.006943f
C497 B.n274 VSUBS 0.006943f
C498 B.n275 VSUBS 0.00633f
C499 B.n276 VSUBS 0.006943f
C500 B.n277 VSUBS 0.006943f
C501 B.n278 VSUBS 0.006943f
C502 B.n279 VSUBS 0.006943f
C503 B.n280 VSUBS 0.006943f
C504 B.n281 VSUBS 0.006943f
C505 B.n282 VSUBS 0.006943f
C506 B.n283 VSUBS 0.006943f
C507 B.n284 VSUBS 0.006943f
C508 B.n285 VSUBS 0.006943f
C509 B.n286 VSUBS 0.006943f
C510 B.n287 VSUBS 0.006943f
C511 B.n288 VSUBS 0.006943f
C512 B.n289 VSUBS 0.006943f
C513 B.n290 VSUBS 0.006943f
C514 B.n291 VSUBS 0.006943f
C515 B.n292 VSUBS 0.006943f
C516 B.n293 VSUBS 0.006943f
C517 B.n294 VSUBS 0.006943f
C518 B.n295 VSUBS 0.006943f
C519 B.n296 VSUBS 0.006943f
C520 B.n297 VSUBS 0.006943f
C521 B.n298 VSUBS 0.006943f
C522 B.n299 VSUBS 0.006943f
C523 B.n300 VSUBS 0.006943f
C524 B.n301 VSUBS 0.006943f
C525 B.n302 VSUBS 0.006943f
C526 B.n303 VSUBS 0.006943f
C527 B.n304 VSUBS 0.006943f
C528 B.n305 VSUBS 0.006943f
C529 B.n306 VSUBS 0.006943f
C530 B.n307 VSUBS 0.006943f
C531 B.n308 VSUBS 0.006943f
C532 B.n309 VSUBS 0.006943f
C533 B.n310 VSUBS 0.006943f
C534 B.n311 VSUBS 0.006943f
C535 B.n312 VSUBS 0.006943f
C536 B.n313 VSUBS 0.006943f
C537 B.n314 VSUBS 0.006943f
C538 B.n315 VSUBS 0.006943f
C539 B.n316 VSUBS 0.006943f
C540 B.n317 VSUBS 0.006943f
C541 B.n318 VSUBS 0.006943f
C542 B.n319 VSUBS 0.006943f
C543 B.n320 VSUBS 0.006943f
C544 B.n321 VSUBS 0.006943f
C545 B.n322 VSUBS 0.006943f
C546 B.n323 VSUBS 0.006943f
C547 B.n324 VSUBS 0.006943f
C548 B.n325 VSUBS 0.006943f
C549 B.n326 VSUBS 0.006943f
C550 B.n327 VSUBS 0.006943f
C551 B.n328 VSUBS 0.006943f
C552 B.n329 VSUBS 0.006943f
C553 B.n330 VSUBS 0.006943f
C554 B.n331 VSUBS 0.006943f
C555 B.n332 VSUBS 0.006943f
C556 B.n333 VSUBS 0.006943f
C557 B.n334 VSUBS 0.006943f
C558 B.n335 VSUBS 0.006943f
C559 B.n336 VSUBS 0.006943f
C560 B.n337 VSUBS 0.006943f
C561 B.n338 VSUBS 0.006943f
C562 B.n339 VSUBS 0.006943f
C563 B.n340 VSUBS 0.006943f
C564 B.n341 VSUBS 0.006943f
C565 B.n342 VSUBS 0.006943f
C566 B.n343 VSUBS 0.006943f
C567 B.n344 VSUBS 0.006943f
C568 B.n345 VSUBS 0.006943f
C569 B.n346 VSUBS 0.006943f
C570 B.n347 VSUBS 0.006943f
C571 B.n348 VSUBS 0.006943f
C572 B.n349 VSUBS 0.006943f
C573 B.n350 VSUBS 0.006943f
C574 B.n351 VSUBS 0.006943f
C575 B.n352 VSUBS 0.006943f
C576 B.n353 VSUBS 0.006943f
C577 B.n354 VSUBS 0.016998f
C578 B.n355 VSUBS 0.015878f
C579 B.n356 VSUBS 0.015878f
C580 B.n357 VSUBS 0.006943f
C581 B.n358 VSUBS 0.006943f
C582 B.n359 VSUBS 0.006943f
C583 B.n360 VSUBS 0.006943f
C584 B.n361 VSUBS 0.006943f
C585 B.n362 VSUBS 0.006943f
C586 B.n363 VSUBS 0.006943f
C587 B.n364 VSUBS 0.006943f
C588 B.n365 VSUBS 0.006943f
C589 B.n366 VSUBS 0.006943f
C590 B.n367 VSUBS 0.006943f
C591 B.n368 VSUBS 0.006943f
C592 B.n369 VSUBS 0.006943f
C593 B.n370 VSUBS 0.006943f
C594 B.n371 VSUBS 0.006943f
C595 B.n372 VSUBS 0.006943f
C596 B.n373 VSUBS 0.006943f
C597 B.n374 VSUBS 0.006943f
C598 B.n375 VSUBS 0.006943f
C599 B.n376 VSUBS 0.006943f
C600 B.n377 VSUBS 0.006943f
C601 B.n378 VSUBS 0.006943f
C602 B.n379 VSUBS 0.006943f
C603 B.n380 VSUBS 0.006943f
C604 B.n381 VSUBS 0.006943f
C605 B.n382 VSUBS 0.006943f
C606 B.n383 VSUBS 0.006943f
C607 B.n384 VSUBS 0.006943f
C608 B.n385 VSUBS 0.006943f
C609 B.n386 VSUBS 0.006943f
C610 B.n387 VSUBS 0.006943f
C611 B.n388 VSUBS 0.006943f
C612 B.n389 VSUBS 0.006943f
C613 B.n390 VSUBS 0.006943f
C614 B.n391 VSUBS 0.006943f
C615 B.n392 VSUBS 0.006943f
C616 B.n393 VSUBS 0.006943f
C617 B.n394 VSUBS 0.006943f
C618 B.n395 VSUBS 0.006943f
C619 B.n396 VSUBS 0.006943f
C620 B.n397 VSUBS 0.016684f
C621 B.n398 VSUBS 0.015878f
C622 B.n399 VSUBS 0.016998f
C623 B.n400 VSUBS 0.006943f
C624 B.n401 VSUBS 0.006943f
C625 B.n402 VSUBS 0.006943f
C626 B.n403 VSUBS 0.006943f
C627 B.n404 VSUBS 0.006943f
C628 B.n405 VSUBS 0.006943f
C629 B.n406 VSUBS 0.006943f
C630 B.n407 VSUBS 0.006943f
C631 B.n408 VSUBS 0.006943f
C632 B.n409 VSUBS 0.006943f
C633 B.n410 VSUBS 0.006943f
C634 B.n411 VSUBS 0.006943f
C635 B.n412 VSUBS 0.006943f
C636 B.n413 VSUBS 0.006943f
C637 B.n414 VSUBS 0.006943f
C638 B.n415 VSUBS 0.006943f
C639 B.n416 VSUBS 0.006943f
C640 B.n417 VSUBS 0.006943f
C641 B.n418 VSUBS 0.006943f
C642 B.n419 VSUBS 0.006943f
C643 B.n420 VSUBS 0.006943f
C644 B.n421 VSUBS 0.006943f
C645 B.n422 VSUBS 0.006943f
C646 B.n423 VSUBS 0.006943f
C647 B.n424 VSUBS 0.006943f
C648 B.n425 VSUBS 0.006943f
C649 B.n426 VSUBS 0.006943f
C650 B.n427 VSUBS 0.006943f
C651 B.n428 VSUBS 0.006943f
C652 B.n429 VSUBS 0.006943f
C653 B.n430 VSUBS 0.006943f
C654 B.n431 VSUBS 0.006943f
C655 B.n432 VSUBS 0.006943f
C656 B.n433 VSUBS 0.006943f
C657 B.n434 VSUBS 0.006943f
C658 B.n435 VSUBS 0.006943f
C659 B.n436 VSUBS 0.006943f
C660 B.n437 VSUBS 0.006943f
C661 B.n438 VSUBS 0.006943f
C662 B.n439 VSUBS 0.006943f
C663 B.n440 VSUBS 0.006943f
C664 B.n441 VSUBS 0.006943f
C665 B.n442 VSUBS 0.006943f
C666 B.n443 VSUBS 0.006943f
C667 B.n444 VSUBS 0.006943f
C668 B.n445 VSUBS 0.006943f
C669 B.n446 VSUBS 0.006943f
C670 B.n447 VSUBS 0.006943f
C671 B.n448 VSUBS 0.006943f
C672 B.n449 VSUBS 0.006943f
C673 B.n450 VSUBS 0.006943f
C674 B.n451 VSUBS 0.006943f
C675 B.n452 VSUBS 0.006943f
C676 B.n453 VSUBS 0.006943f
C677 B.n454 VSUBS 0.006943f
C678 B.n455 VSUBS 0.006943f
C679 B.n456 VSUBS 0.006943f
C680 B.n457 VSUBS 0.006943f
C681 B.n458 VSUBS 0.006943f
C682 B.n459 VSUBS 0.006943f
C683 B.n460 VSUBS 0.006943f
C684 B.n461 VSUBS 0.006943f
C685 B.n462 VSUBS 0.006943f
C686 B.n463 VSUBS 0.006943f
C687 B.n464 VSUBS 0.006943f
C688 B.n465 VSUBS 0.006943f
C689 B.n466 VSUBS 0.006943f
C690 B.n467 VSUBS 0.006943f
C691 B.n468 VSUBS 0.006943f
C692 B.n469 VSUBS 0.006943f
C693 B.n470 VSUBS 0.006943f
C694 B.n471 VSUBS 0.006943f
C695 B.n472 VSUBS 0.006943f
C696 B.n473 VSUBS 0.006943f
C697 B.n474 VSUBS 0.006943f
C698 B.n475 VSUBS 0.006943f
C699 B.n476 VSUBS 0.006943f
C700 B.n477 VSUBS 0.006943f
C701 B.n478 VSUBS 0.006943f
C702 B.n479 VSUBS 0.00633f
C703 B.n480 VSUBS 0.016086f
C704 B.n481 VSUBS 0.004084f
C705 B.n482 VSUBS 0.006943f
C706 B.n483 VSUBS 0.006943f
C707 B.n484 VSUBS 0.006943f
C708 B.n485 VSUBS 0.006943f
C709 B.n486 VSUBS 0.006943f
C710 B.n487 VSUBS 0.006943f
C711 B.n488 VSUBS 0.006943f
C712 B.n489 VSUBS 0.006943f
C713 B.n490 VSUBS 0.006943f
C714 B.n491 VSUBS 0.006943f
C715 B.n492 VSUBS 0.006943f
C716 B.n493 VSUBS 0.006943f
C717 B.n494 VSUBS 0.004084f
C718 B.n495 VSUBS 0.006943f
C719 B.n496 VSUBS 0.006943f
C720 B.n497 VSUBS 0.00633f
C721 B.n498 VSUBS 0.006943f
C722 B.n499 VSUBS 0.006943f
C723 B.n500 VSUBS 0.006943f
C724 B.n501 VSUBS 0.006943f
C725 B.n502 VSUBS 0.006943f
C726 B.n503 VSUBS 0.006943f
C727 B.n504 VSUBS 0.006943f
C728 B.n505 VSUBS 0.006943f
C729 B.n506 VSUBS 0.006943f
C730 B.n507 VSUBS 0.006943f
C731 B.n508 VSUBS 0.006943f
C732 B.n509 VSUBS 0.006943f
C733 B.n510 VSUBS 0.006943f
C734 B.n511 VSUBS 0.006943f
C735 B.n512 VSUBS 0.006943f
C736 B.n513 VSUBS 0.006943f
C737 B.n514 VSUBS 0.006943f
C738 B.n515 VSUBS 0.006943f
C739 B.n516 VSUBS 0.006943f
C740 B.n517 VSUBS 0.006943f
C741 B.n518 VSUBS 0.006943f
C742 B.n519 VSUBS 0.006943f
C743 B.n520 VSUBS 0.006943f
C744 B.n521 VSUBS 0.006943f
C745 B.n522 VSUBS 0.006943f
C746 B.n523 VSUBS 0.006943f
C747 B.n524 VSUBS 0.006943f
C748 B.n525 VSUBS 0.006943f
C749 B.n526 VSUBS 0.006943f
C750 B.n527 VSUBS 0.006943f
C751 B.n528 VSUBS 0.006943f
C752 B.n529 VSUBS 0.006943f
C753 B.n530 VSUBS 0.006943f
C754 B.n531 VSUBS 0.006943f
C755 B.n532 VSUBS 0.006943f
C756 B.n533 VSUBS 0.006943f
C757 B.n534 VSUBS 0.006943f
C758 B.n535 VSUBS 0.006943f
C759 B.n536 VSUBS 0.006943f
C760 B.n537 VSUBS 0.006943f
C761 B.n538 VSUBS 0.006943f
C762 B.n539 VSUBS 0.006943f
C763 B.n540 VSUBS 0.006943f
C764 B.n541 VSUBS 0.006943f
C765 B.n542 VSUBS 0.006943f
C766 B.n543 VSUBS 0.006943f
C767 B.n544 VSUBS 0.006943f
C768 B.n545 VSUBS 0.006943f
C769 B.n546 VSUBS 0.006943f
C770 B.n547 VSUBS 0.006943f
C771 B.n548 VSUBS 0.006943f
C772 B.n549 VSUBS 0.006943f
C773 B.n550 VSUBS 0.006943f
C774 B.n551 VSUBS 0.006943f
C775 B.n552 VSUBS 0.006943f
C776 B.n553 VSUBS 0.006943f
C777 B.n554 VSUBS 0.006943f
C778 B.n555 VSUBS 0.006943f
C779 B.n556 VSUBS 0.006943f
C780 B.n557 VSUBS 0.006943f
C781 B.n558 VSUBS 0.006943f
C782 B.n559 VSUBS 0.006943f
C783 B.n560 VSUBS 0.006943f
C784 B.n561 VSUBS 0.006943f
C785 B.n562 VSUBS 0.006943f
C786 B.n563 VSUBS 0.006943f
C787 B.n564 VSUBS 0.006943f
C788 B.n565 VSUBS 0.006943f
C789 B.n566 VSUBS 0.006943f
C790 B.n567 VSUBS 0.006943f
C791 B.n568 VSUBS 0.006943f
C792 B.n569 VSUBS 0.006943f
C793 B.n570 VSUBS 0.006943f
C794 B.n571 VSUBS 0.006943f
C795 B.n572 VSUBS 0.006943f
C796 B.n573 VSUBS 0.006943f
C797 B.n574 VSUBS 0.006943f
C798 B.n575 VSUBS 0.006943f
C799 B.n576 VSUBS 0.016998f
C800 B.n577 VSUBS 0.015878f
C801 B.n578 VSUBS 0.015878f
C802 B.n579 VSUBS 0.006943f
C803 B.n580 VSUBS 0.006943f
C804 B.n581 VSUBS 0.006943f
C805 B.n582 VSUBS 0.006943f
C806 B.n583 VSUBS 0.006943f
C807 B.n584 VSUBS 0.006943f
C808 B.n585 VSUBS 0.006943f
C809 B.n586 VSUBS 0.006943f
C810 B.n587 VSUBS 0.006943f
C811 B.n588 VSUBS 0.006943f
C812 B.n589 VSUBS 0.006943f
C813 B.n590 VSUBS 0.006943f
C814 B.n591 VSUBS 0.006943f
C815 B.n592 VSUBS 0.006943f
C816 B.n593 VSUBS 0.006943f
C817 B.n594 VSUBS 0.006943f
C818 B.n595 VSUBS 0.006943f
C819 B.n596 VSUBS 0.006943f
C820 B.n597 VSUBS 0.006943f
C821 B.n598 VSUBS 0.006943f
C822 B.n599 VSUBS 0.015721f
C823 VDD1.n0 VSUBS 0.023068f
C824 VDD1.n1 VSUBS 0.020832f
C825 VDD1.n2 VSUBS 0.011194f
C826 VDD1.n3 VSUBS 0.026459f
C827 VDD1.n4 VSUBS 0.011853f
C828 VDD1.n5 VSUBS 0.020832f
C829 VDD1.n6 VSUBS 0.011523f
C830 VDD1.n7 VSUBS 0.026459f
C831 VDD1.n8 VSUBS 0.011194f
C832 VDD1.n9 VSUBS 0.011853f
C833 VDD1.n10 VSUBS 0.020832f
C834 VDD1.n11 VSUBS 0.011194f
C835 VDD1.n12 VSUBS 0.026459f
C836 VDD1.n13 VSUBS 0.011853f
C837 VDD1.n14 VSUBS 0.020832f
C838 VDD1.n15 VSUBS 0.011194f
C839 VDD1.n16 VSUBS 0.026459f
C840 VDD1.n17 VSUBS 0.011853f
C841 VDD1.n18 VSUBS 0.020832f
C842 VDD1.n19 VSUBS 0.011194f
C843 VDD1.n20 VSUBS 0.026459f
C844 VDD1.n21 VSUBS 0.011853f
C845 VDD1.n22 VSUBS 0.020832f
C846 VDD1.n23 VSUBS 0.011194f
C847 VDD1.n24 VSUBS 0.026459f
C848 VDD1.n25 VSUBS 0.011853f
C849 VDD1.n26 VSUBS 0.020832f
C850 VDD1.n27 VSUBS 0.011194f
C851 VDD1.n28 VSUBS 0.019844f
C852 VDD1.n29 VSUBS 0.016832f
C853 VDD1.t1 VSUBS 0.056707f
C854 VDD1.n30 VSUBS 0.154405f
C855 VDD1.n31 VSUBS 1.44648f
C856 VDD1.n32 VSUBS 0.011194f
C857 VDD1.n33 VSUBS 0.011853f
C858 VDD1.n34 VSUBS 0.026459f
C859 VDD1.n35 VSUBS 0.026459f
C860 VDD1.n36 VSUBS 0.011853f
C861 VDD1.n37 VSUBS 0.011194f
C862 VDD1.n38 VSUBS 0.020832f
C863 VDD1.n39 VSUBS 0.020832f
C864 VDD1.n40 VSUBS 0.011194f
C865 VDD1.n41 VSUBS 0.011853f
C866 VDD1.n42 VSUBS 0.026459f
C867 VDD1.n43 VSUBS 0.026459f
C868 VDD1.n44 VSUBS 0.011853f
C869 VDD1.n45 VSUBS 0.011194f
C870 VDD1.n46 VSUBS 0.020832f
C871 VDD1.n47 VSUBS 0.020832f
C872 VDD1.n48 VSUBS 0.011194f
C873 VDD1.n49 VSUBS 0.011853f
C874 VDD1.n50 VSUBS 0.026459f
C875 VDD1.n51 VSUBS 0.026459f
C876 VDD1.n52 VSUBS 0.011853f
C877 VDD1.n53 VSUBS 0.011194f
C878 VDD1.n54 VSUBS 0.020832f
C879 VDD1.n55 VSUBS 0.020832f
C880 VDD1.n56 VSUBS 0.011194f
C881 VDD1.n57 VSUBS 0.011853f
C882 VDD1.n58 VSUBS 0.026459f
C883 VDD1.n59 VSUBS 0.026459f
C884 VDD1.n60 VSUBS 0.011853f
C885 VDD1.n61 VSUBS 0.011194f
C886 VDD1.n62 VSUBS 0.020832f
C887 VDD1.n63 VSUBS 0.020832f
C888 VDD1.n64 VSUBS 0.011194f
C889 VDD1.n65 VSUBS 0.011853f
C890 VDD1.n66 VSUBS 0.026459f
C891 VDD1.n67 VSUBS 0.026459f
C892 VDD1.n68 VSUBS 0.011853f
C893 VDD1.n69 VSUBS 0.011194f
C894 VDD1.n70 VSUBS 0.020832f
C895 VDD1.n71 VSUBS 0.020832f
C896 VDD1.n72 VSUBS 0.011194f
C897 VDD1.n73 VSUBS 0.011853f
C898 VDD1.n74 VSUBS 0.026459f
C899 VDD1.n75 VSUBS 0.026459f
C900 VDD1.n76 VSUBS 0.026459f
C901 VDD1.n77 VSUBS 0.011523f
C902 VDD1.n78 VSUBS 0.011194f
C903 VDD1.n79 VSUBS 0.020832f
C904 VDD1.n80 VSUBS 0.020832f
C905 VDD1.n81 VSUBS 0.011194f
C906 VDD1.n82 VSUBS 0.011853f
C907 VDD1.n83 VSUBS 0.026459f
C908 VDD1.n84 VSUBS 0.06466f
C909 VDD1.n85 VSUBS 0.011853f
C910 VDD1.n86 VSUBS 0.011194f
C911 VDD1.n87 VSUBS 0.052421f
C912 VDD1.n88 VSUBS 0.047354f
C913 VDD1.n89 VSUBS 0.023068f
C914 VDD1.n90 VSUBS 0.020832f
C915 VDD1.n91 VSUBS 0.011194f
C916 VDD1.n92 VSUBS 0.026459f
C917 VDD1.n93 VSUBS 0.011853f
C918 VDD1.n94 VSUBS 0.020832f
C919 VDD1.n95 VSUBS 0.011523f
C920 VDD1.n96 VSUBS 0.026459f
C921 VDD1.n97 VSUBS 0.011853f
C922 VDD1.n98 VSUBS 0.020832f
C923 VDD1.n99 VSUBS 0.011194f
C924 VDD1.n100 VSUBS 0.026459f
C925 VDD1.n101 VSUBS 0.011853f
C926 VDD1.n102 VSUBS 0.020832f
C927 VDD1.n103 VSUBS 0.011194f
C928 VDD1.n104 VSUBS 0.026459f
C929 VDD1.n105 VSUBS 0.011853f
C930 VDD1.n106 VSUBS 0.020832f
C931 VDD1.n107 VSUBS 0.011194f
C932 VDD1.n108 VSUBS 0.026459f
C933 VDD1.n109 VSUBS 0.011853f
C934 VDD1.n110 VSUBS 0.020832f
C935 VDD1.n111 VSUBS 0.011194f
C936 VDD1.n112 VSUBS 0.026459f
C937 VDD1.n113 VSUBS 0.011853f
C938 VDD1.n114 VSUBS 0.020832f
C939 VDD1.n115 VSUBS 0.011194f
C940 VDD1.n116 VSUBS 0.019844f
C941 VDD1.n117 VSUBS 0.016832f
C942 VDD1.t0 VSUBS 0.056707f
C943 VDD1.n118 VSUBS 0.154405f
C944 VDD1.n119 VSUBS 1.44648f
C945 VDD1.n120 VSUBS 0.011194f
C946 VDD1.n121 VSUBS 0.011853f
C947 VDD1.n122 VSUBS 0.026459f
C948 VDD1.n123 VSUBS 0.026459f
C949 VDD1.n124 VSUBS 0.011853f
C950 VDD1.n125 VSUBS 0.011194f
C951 VDD1.n126 VSUBS 0.020832f
C952 VDD1.n127 VSUBS 0.020832f
C953 VDD1.n128 VSUBS 0.011194f
C954 VDD1.n129 VSUBS 0.011853f
C955 VDD1.n130 VSUBS 0.026459f
C956 VDD1.n131 VSUBS 0.026459f
C957 VDD1.n132 VSUBS 0.011853f
C958 VDD1.n133 VSUBS 0.011194f
C959 VDD1.n134 VSUBS 0.020832f
C960 VDD1.n135 VSUBS 0.020832f
C961 VDD1.n136 VSUBS 0.011194f
C962 VDD1.n137 VSUBS 0.011853f
C963 VDD1.n138 VSUBS 0.026459f
C964 VDD1.n139 VSUBS 0.026459f
C965 VDD1.n140 VSUBS 0.011853f
C966 VDD1.n141 VSUBS 0.011194f
C967 VDD1.n142 VSUBS 0.020832f
C968 VDD1.n143 VSUBS 0.020832f
C969 VDD1.n144 VSUBS 0.011194f
C970 VDD1.n145 VSUBS 0.011853f
C971 VDD1.n146 VSUBS 0.026459f
C972 VDD1.n147 VSUBS 0.026459f
C973 VDD1.n148 VSUBS 0.011853f
C974 VDD1.n149 VSUBS 0.011194f
C975 VDD1.n150 VSUBS 0.020832f
C976 VDD1.n151 VSUBS 0.020832f
C977 VDD1.n152 VSUBS 0.011194f
C978 VDD1.n153 VSUBS 0.011853f
C979 VDD1.n154 VSUBS 0.026459f
C980 VDD1.n155 VSUBS 0.026459f
C981 VDD1.n156 VSUBS 0.011853f
C982 VDD1.n157 VSUBS 0.011194f
C983 VDD1.n158 VSUBS 0.020832f
C984 VDD1.n159 VSUBS 0.020832f
C985 VDD1.n160 VSUBS 0.011194f
C986 VDD1.n161 VSUBS 0.011194f
C987 VDD1.n162 VSUBS 0.011853f
C988 VDD1.n163 VSUBS 0.026459f
C989 VDD1.n164 VSUBS 0.026459f
C990 VDD1.n165 VSUBS 0.026459f
C991 VDD1.n166 VSUBS 0.011523f
C992 VDD1.n167 VSUBS 0.011194f
C993 VDD1.n168 VSUBS 0.020832f
C994 VDD1.n169 VSUBS 0.020832f
C995 VDD1.n170 VSUBS 0.011194f
C996 VDD1.n171 VSUBS 0.011853f
C997 VDD1.n172 VSUBS 0.026459f
C998 VDD1.n173 VSUBS 0.06466f
C999 VDD1.n174 VSUBS 0.011853f
C1000 VDD1.n175 VSUBS 0.011194f
C1001 VDD1.n176 VSUBS 0.052421f
C1002 VDD1.n177 VSUBS 0.646561f
C1003 VTAIL.n0 VSUBS 0.026552f
C1004 VTAIL.n1 VSUBS 0.023979f
C1005 VTAIL.n2 VSUBS 0.012885f
C1006 VTAIL.n3 VSUBS 0.030455f
C1007 VTAIL.n4 VSUBS 0.013643f
C1008 VTAIL.n5 VSUBS 0.023979f
C1009 VTAIL.n6 VSUBS 0.013264f
C1010 VTAIL.n7 VSUBS 0.030455f
C1011 VTAIL.n8 VSUBS 0.013643f
C1012 VTAIL.n9 VSUBS 0.023979f
C1013 VTAIL.n10 VSUBS 0.012885f
C1014 VTAIL.n11 VSUBS 0.030455f
C1015 VTAIL.n12 VSUBS 0.013643f
C1016 VTAIL.n13 VSUBS 0.023979f
C1017 VTAIL.n14 VSUBS 0.012885f
C1018 VTAIL.n15 VSUBS 0.030455f
C1019 VTAIL.n16 VSUBS 0.013643f
C1020 VTAIL.n17 VSUBS 0.023979f
C1021 VTAIL.n18 VSUBS 0.012885f
C1022 VTAIL.n19 VSUBS 0.030455f
C1023 VTAIL.n20 VSUBS 0.013643f
C1024 VTAIL.n21 VSUBS 0.023979f
C1025 VTAIL.n22 VSUBS 0.012885f
C1026 VTAIL.n23 VSUBS 0.030455f
C1027 VTAIL.n24 VSUBS 0.013643f
C1028 VTAIL.n25 VSUBS 0.023979f
C1029 VTAIL.n26 VSUBS 0.012885f
C1030 VTAIL.n27 VSUBS 0.022842f
C1031 VTAIL.n28 VSUBS 0.019374f
C1032 VTAIL.t1 VSUBS 0.065272f
C1033 VTAIL.n29 VSUBS 0.177727f
C1034 VTAIL.n30 VSUBS 1.66497f
C1035 VTAIL.n31 VSUBS 0.012885f
C1036 VTAIL.n32 VSUBS 0.013643f
C1037 VTAIL.n33 VSUBS 0.030455f
C1038 VTAIL.n34 VSUBS 0.030455f
C1039 VTAIL.n35 VSUBS 0.013643f
C1040 VTAIL.n36 VSUBS 0.012885f
C1041 VTAIL.n37 VSUBS 0.023979f
C1042 VTAIL.n38 VSUBS 0.023979f
C1043 VTAIL.n39 VSUBS 0.012885f
C1044 VTAIL.n40 VSUBS 0.013643f
C1045 VTAIL.n41 VSUBS 0.030455f
C1046 VTAIL.n42 VSUBS 0.030455f
C1047 VTAIL.n43 VSUBS 0.013643f
C1048 VTAIL.n44 VSUBS 0.012885f
C1049 VTAIL.n45 VSUBS 0.023979f
C1050 VTAIL.n46 VSUBS 0.023979f
C1051 VTAIL.n47 VSUBS 0.012885f
C1052 VTAIL.n48 VSUBS 0.013643f
C1053 VTAIL.n49 VSUBS 0.030455f
C1054 VTAIL.n50 VSUBS 0.030455f
C1055 VTAIL.n51 VSUBS 0.013643f
C1056 VTAIL.n52 VSUBS 0.012885f
C1057 VTAIL.n53 VSUBS 0.023979f
C1058 VTAIL.n54 VSUBS 0.023979f
C1059 VTAIL.n55 VSUBS 0.012885f
C1060 VTAIL.n56 VSUBS 0.013643f
C1061 VTAIL.n57 VSUBS 0.030455f
C1062 VTAIL.n58 VSUBS 0.030455f
C1063 VTAIL.n59 VSUBS 0.013643f
C1064 VTAIL.n60 VSUBS 0.012885f
C1065 VTAIL.n61 VSUBS 0.023979f
C1066 VTAIL.n62 VSUBS 0.023979f
C1067 VTAIL.n63 VSUBS 0.012885f
C1068 VTAIL.n64 VSUBS 0.013643f
C1069 VTAIL.n65 VSUBS 0.030455f
C1070 VTAIL.n66 VSUBS 0.030455f
C1071 VTAIL.n67 VSUBS 0.013643f
C1072 VTAIL.n68 VSUBS 0.012885f
C1073 VTAIL.n69 VSUBS 0.023979f
C1074 VTAIL.n70 VSUBS 0.023979f
C1075 VTAIL.n71 VSUBS 0.012885f
C1076 VTAIL.n72 VSUBS 0.012885f
C1077 VTAIL.n73 VSUBS 0.013643f
C1078 VTAIL.n74 VSUBS 0.030455f
C1079 VTAIL.n75 VSUBS 0.030455f
C1080 VTAIL.n76 VSUBS 0.030455f
C1081 VTAIL.n77 VSUBS 0.013264f
C1082 VTAIL.n78 VSUBS 0.012885f
C1083 VTAIL.n79 VSUBS 0.023979f
C1084 VTAIL.n80 VSUBS 0.023979f
C1085 VTAIL.n81 VSUBS 0.012885f
C1086 VTAIL.n82 VSUBS 0.013643f
C1087 VTAIL.n83 VSUBS 0.030455f
C1088 VTAIL.n84 VSUBS 0.074427f
C1089 VTAIL.n85 VSUBS 0.013643f
C1090 VTAIL.n86 VSUBS 0.012885f
C1091 VTAIL.n87 VSUBS 0.060339f
C1092 VTAIL.n88 VSUBS 0.037605f
C1093 VTAIL.n89 VSUBS 1.6265f
C1094 VTAIL.n90 VSUBS 0.026552f
C1095 VTAIL.n91 VSUBS 0.023979f
C1096 VTAIL.n92 VSUBS 0.012885f
C1097 VTAIL.n93 VSUBS 0.030455f
C1098 VTAIL.n94 VSUBS 0.013643f
C1099 VTAIL.n95 VSUBS 0.023979f
C1100 VTAIL.n96 VSUBS 0.013264f
C1101 VTAIL.n97 VSUBS 0.030455f
C1102 VTAIL.n98 VSUBS 0.012885f
C1103 VTAIL.n99 VSUBS 0.013643f
C1104 VTAIL.n100 VSUBS 0.023979f
C1105 VTAIL.n101 VSUBS 0.012885f
C1106 VTAIL.n102 VSUBS 0.030455f
C1107 VTAIL.n103 VSUBS 0.013643f
C1108 VTAIL.n104 VSUBS 0.023979f
C1109 VTAIL.n105 VSUBS 0.012885f
C1110 VTAIL.n106 VSUBS 0.030455f
C1111 VTAIL.n107 VSUBS 0.013643f
C1112 VTAIL.n108 VSUBS 0.023979f
C1113 VTAIL.n109 VSUBS 0.012885f
C1114 VTAIL.n110 VSUBS 0.030455f
C1115 VTAIL.n111 VSUBS 0.013643f
C1116 VTAIL.n112 VSUBS 0.023979f
C1117 VTAIL.n113 VSUBS 0.012885f
C1118 VTAIL.n114 VSUBS 0.030455f
C1119 VTAIL.n115 VSUBS 0.013643f
C1120 VTAIL.n116 VSUBS 0.023979f
C1121 VTAIL.n117 VSUBS 0.012885f
C1122 VTAIL.n118 VSUBS 0.022842f
C1123 VTAIL.n119 VSUBS 0.019374f
C1124 VTAIL.t3 VSUBS 0.065272f
C1125 VTAIL.n120 VSUBS 0.177727f
C1126 VTAIL.n121 VSUBS 1.66497f
C1127 VTAIL.n122 VSUBS 0.012885f
C1128 VTAIL.n123 VSUBS 0.013643f
C1129 VTAIL.n124 VSUBS 0.030455f
C1130 VTAIL.n125 VSUBS 0.030455f
C1131 VTAIL.n126 VSUBS 0.013643f
C1132 VTAIL.n127 VSUBS 0.012885f
C1133 VTAIL.n128 VSUBS 0.023979f
C1134 VTAIL.n129 VSUBS 0.023979f
C1135 VTAIL.n130 VSUBS 0.012885f
C1136 VTAIL.n131 VSUBS 0.013643f
C1137 VTAIL.n132 VSUBS 0.030455f
C1138 VTAIL.n133 VSUBS 0.030455f
C1139 VTAIL.n134 VSUBS 0.013643f
C1140 VTAIL.n135 VSUBS 0.012885f
C1141 VTAIL.n136 VSUBS 0.023979f
C1142 VTAIL.n137 VSUBS 0.023979f
C1143 VTAIL.n138 VSUBS 0.012885f
C1144 VTAIL.n139 VSUBS 0.013643f
C1145 VTAIL.n140 VSUBS 0.030455f
C1146 VTAIL.n141 VSUBS 0.030455f
C1147 VTAIL.n142 VSUBS 0.013643f
C1148 VTAIL.n143 VSUBS 0.012885f
C1149 VTAIL.n144 VSUBS 0.023979f
C1150 VTAIL.n145 VSUBS 0.023979f
C1151 VTAIL.n146 VSUBS 0.012885f
C1152 VTAIL.n147 VSUBS 0.013643f
C1153 VTAIL.n148 VSUBS 0.030455f
C1154 VTAIL.n149 VSUBS 0.030455f
C1155 VTAIL.n150 VSUBS 0.013643f
C1156 VTAIL.n151 VSUBS 0.012885f
C1157 VTAIL.n152 VSUBS 0.023979f
C1158 VTAIL.n153 VSUBS 0.023979f
C1159 VTAIL.n154 VSUBS 0.012885f
C1160 VTAIL.n155 VSUBS 0.013643f
C1161 VTAIL.n156 VSUBS 0.030455f
C1162 VTAIL.n157 VSUBS 0.030455f
C1163 VTAIL.n158 VSUBS 0.013643f
C1164 VTAIL.n159 VSUBS 0.012885f
C1165 VTAIL.n160 VSUBS 0.023979f
C1166 VTAIL.n161 VSUBS 0.023979f
C1167 VTAIL.n162 VSUBS 0.012885f
C1168 VTAIL.n163 VSUBS 0.013643f
C1169 VTAIL.n164 VSUBS 0.030455f
C1170 VTAIL.n165 VSUBS 0.030455f
C1171 VTAIL.n166 VSUBS 0.030455f
C1172 VTAIL.n167 VSUBS 0.013264f
C1173 VTAIL.n168 VSUBS 0.012885f
C1174 VTAIL.n169 VSUBS 0.023979f
C1175 VTAIL.n170 VSUBS 0.023979f
C1176 VTAIL.n171 VSUBS 0.012885f
C1177 VTAIL.n172 VSUBS 0.013643f
C1178 VTAIL.n173 VSUBS 0.030455f
C1179 VTAIL.n174 VSUBS 0.074427f
C1180 VTAIL.n175 VSUBS 0.013643f
C1181 VTAIL.n176 VSUBS 0.012885f
C1182 VTAIL.n177 VSUBS 0.060339f
C1183 VTAIL.n178 VSUBS 0.037605f
C1184 VTAIL.n179 VSUBS 1.63916f
C1185 VTAIL.n180 VSUBS 0.026552f
C1186 VTAIL.n181 VSUBS 0.023979f
C1187 VTAIL.n182 VSUBS 0.012885f
C1188 VTAIL.n183 VSUBS 0.030455f
C1189 VTAIL.n184 VSUBS 0.013643f
C1190 VTAIL.n185 VSUBS 0.023979f
C1191 VTAIL.n186 VSUBS 0.013264f
C1192 VTAIL.n187 VSUBS 0.030455f
C1193 VTAIL.n188 VSUBS 0.012885f
C1194 VTAIL.n189 VSUBS 0.013643f
C1195 VTAIL.n190 VSUBS 0.023979f
C1196 VTAIL.n191 VSUBS 0.012885f
C1197 VTAIL.n192 VSUBS 0.030455f
C1198 VTAIL.n193 VSUBS 0.013643f
C1199 VTAIL.n194 VSUBS 0.023979f
C1200 VTAIL.n195 VSUBS 0.012885f
C1201 VTAIL.n196 VSUBS 0.030455f
C1202 VTAIL.n197 VSUBS 0.013643f
C1203 VTAIL.n198 VSUBS 0.023979f
C1204 VTAIL.n199 VSUBS 0.012885f
C1205 VTAIL.n200 VSUBS 0.030455f
C1206 VTAIL.n201 VSUBS 0.013643f
C1207 VTAIL.n202 VSUBS 0.023979f
C1208 VTAIL.n203 VSUBS 0.012885f
C1209 VTAIL.n204 VSUBS 0.030455f
C1210 VTAIL.n205 VSUBS 0.013643f
C1211 VTAIL.n206 VSUBS 0.023979f
C1212 VTAIL.n207 VSUBS 0.012885f
C1213 VTAIL.n208 VSUBS 0.022842f
C1214 VTAIL.n209 VSUBS 0.019374f
C1215 VTAIL.t2 VSUBS 0.065272f
C1216 VTAIL.n210 VSUBS 0.177727f
C1217 VTAIL.n211 VSUBS 1.66497f
C1218 VTAIL.n212 VSUBS 0.012885f
C1219 VTAIL.n213 VSUBS 0.013643f
C1220 VTAIL.n214 VSUBS 0.030455f
C1221 VTAIL.n215 VSUBS 0.030455f
C1222 VTAIL.n216 VSUBS 0.013643f
C1223 VTAIL.n217 VSUBS 0.012885f
C1224 VTAIL.n218 VSUBS 0.023979f
C1225 VTAIL.n219 VSUBS 0.023979f
C1226 VTAIL.n220 VSUBS 0.012885f
C1227 VTAIL.n221 VSUBS 0.013643f
C1228 VTAIL.n222 VSUBS 0.030455f
C1229 VTAIL.n223 VSUBS 0.030455f
C1230 VTAIL.n224 VSUBS 0.013643f
C1231 VTAIL.n225 VSUBS 0.012885f
C1232 VTAIL.n226 VSUBS 0.023979f
C1233 VTAIL.n227 VSUBS 0.023979f
C1234 VTAIL.n228 VSUBS 0.012885f
C1235 VTAIL.n229 VSUBS 0.013643f
C1236 VTAIL.n230 VSUBS 0.030455f
C1237 VTAIL.n231 VSUBS 0.030455f
C1238 VTAIL.n232 VSUBS 0.013643f
C1239 VTAIL.n233 VSUBS 0.012885f
C1240 VTAIL.n234 VSUBS 0.023979f
C1241 VTAIL.n235 VSUBS 0.023979f
C1242 VTAIL.n236 VSUBS 0.012885f
C1243 VTAIL.n237 VSUBS 0.013643f
C1244 VTAIL.n238 VSUBS 0.030455f
C1245 VTAIL.n239 VSUBS 0.030455f
C1246 VTAIL.n240 VSUBS 0.013643f
C1247 VTAIL.n241 VSUBS 0.012885f
C1248 VTAIL.n242 VSUBS 0.023979f
C1249 VTAIL.n243 VSUBS 0.023979f
C1250 VTAIL.n244 VSUBS 0.012885f
C1251 VTAIL.n245 VSUBS 0.013643f
C1252 VTAIL.n246 VSUBS 0.030455f
C1253 VTAIL.n247 VSUBS 0.030455f
C1254 VTAIL.n248 VSUBS 0.013643f
C1255 VTAIL.n249 VSUBS 0.012885f
C1256 VTAIL.n250 VSUBS 0.023979f
C1257 VTAIL.n251 VSUBS 0.023979f
C1258 VTAIL.n252 VSUBS 0.012885f
C1259 VTAIL.n253 VSUBS 0.013643f
C1260 VTAIL.n254 VSUBS 0.030455f
C1261 VTAIL.n255 VSUBS 0.030455f
C1262 VTAIL.n256 VSUBS 0.030455f
C1263 VTAIL.n257 VSUBS 0.013264f
C1264 VTAIL.n258 VSUBS 0.012885f
C1265 VTAIL.n259 VSUBS 0.023979f
C1266 VTAIL.n260 VSUBS 0.023979f
C1267 VTAIL.n261 VSUBS 0.012885f
C1268 VTAIL.n262 VSUBS 0.013643f
C1269 VTAIL.n263 VSUBS 0.030455f
C1270 VTAIL.n264 VSUBS 0.074427f
C1271 VTAIL.n265 VSUBS 0.013643f
C1272 VTAIL.n266 VSUBS 0.012885f
C1273 VTAIL.n267 VSUBS 0.060339f
C1274 VTAIL.n268 VSUBS 0.037605f
C1275 VTAIL.n269 VSUBS 1.57055f
C1276 VTAIL.n270 VSUBS 0.026552f
C1277 VTAIL.n271 VSUBS 0.023979f
C1278 VTAIL.n272 VSUBS 0.012885f
C1279 VTAIL.n273 VSUBS 0.030455f
C1280 VTAIL.n274 VSUBS 0.013643f
C1281 VTAIL.n275 VSUBS 0.023979f
C1282 VTAIL.n276 VSUBS 0.013264f
C1283 VTAIL.n277 VSUBS 0.030455f
C1284 VTAIL.n278 VSUBS 0.013643f
C1285 VTAIL.n279 VSUBS 0.023979f
C1286 VTAIL.n280 VSUBS 0.012885f
C1287 VTAIL.n281 VSUBS 0.030455f
C1288 VTAIL.n282 VSUBS 0.013643f
C1289 VTAIL.n283 VSUBS 0.023979f
C1290 VTAIL.n284 VSUBS 0.012885f
C1291 VTAIL.n285 VSUBS 0.030455f
C1292 VTAIL.n286 VSUBS 0.013643f
C1293 VTAIL.n287 VSUBS 0.023979f
C1294 VTAIL.n288 VSUBS 0.012885f
C1295 VTAIL.n289 VSUBS 0.030455f
C1296 VTAIL.n290 VSUBS 0.013643f
C1297 VTAIL.n291 VSUBS 0.023979f
C1298 VTAIL.n292 VSUBS 0.012885f
C1299 VTAIL.n293 VSUBS 0.030455f
C1300 VTAIL.n294 VSUBS 0.013643f
C1301 VTAIL.n295 VSUBS 0.023979f
C1302 VTAIL.n296 VSUBS 0.012885f
C1303 VTAIL.n297 VSUBS 0.022842f
C1304 VTAIL.n298 VSUBS 0.019374f
C1305 VTAIL.t0 VSUBS 0.065272f
C1306 VTAIL.n299 VSUBS 0.177727f
C1307 VTAIL.n300 VSUBS 1.66497f
C1308 VTAIL.n301 VSUBS 0.012885f
C1309 VTAIL.n302 VSUBS 0.013643f
C1310 VTAIL.n303 VSUBS 0.030455f
C1311 VTAIL.n304 VSUBS 0.030455f
C1312 VTAIL.n305 VSUBS 0.013643f
C1313 VTAIL.n306 VSUBS 0.012885f
C1314 VTAIL.n307 VSUBS 0.023979f
C1315 VTAIL.n308 VSUBS 0.023979f
C1316 VTAIL.n309 VSUBS 0.012885f
C1317 VTAIL.n310 VSUBS 0.013643f
C1318 VTAIL.n311 VSUBS 0.030455f
C1319 VTAIL.n312 VSUBS 0.030455f
C1320 VTAIL.n313 VSUBS 0.013643f
C1321 VTAIL.n314 VSUBS 0.012885f
C1322 VTAIL.n315 VSUBS 0.023979f
C1323 VTAIL.n316 VSUBS 0.023979f
C1324 VTAIL.n317 VSUBS 0.012885f
C1325 VTAIL.n318 VSUBS 0.013643f
C1326 VTAIL.n319 VSUBS 0.030455f
C1327 VTAIL.n320 VSUBS 0.030455f
C1328 VTAIL.n321 VSUBS 0.013643f
C1329 VTAIL.n322 VSUBS 0.012885f
C1330 VTAIL.n323 VSUBS 0.023979f
C1331 VTAIL.n324 VSUBS 0.023979f
C1332 VTAIL.n325 VSUBS 0.012885f
C1333 VTAIL.n326 VSUBS 0.013643f
C1334 VTAIL.n327 VSUBS 0.030455f
C1335 VTAIL.n328 VSUBS 0.030455f
C1336 VTAIL.n329 VSUBS 0.013643f
C1337 VTAIL.n330 VSUBS 0.012885f
C1338 VTAIL.n331 VSUBS 0.023979f
C1339 VTAIL.n332 VSUBS 0.023979f
C1340 VTAIL.n333 VSUBS 0.012885f
C1341 VTAIL.n334 VSUBS 0.013643f
C1342 VTAIL.n335 VSUBS 0.030455f
C1343 VTAIL.n336 VSUBS 0.030455f
C1344 VTAIL.n337 VSUBS 0.013643f
C1345 VTAIL.n338 VSUBS 0.012885f
C1346 VTAIL.n339 VSUBS 0.023979f
C1347 VTAIL.n340 VSUBS 0.023979f
C1348 VTAIL.n341 VSUBS 0.012885f
C1349 VTAIL.n342 VSUBS 0.012885f
C1350 VTAIL.n343 VSUBS 0.013643f
C1351 VTAIL.n344 VSUBS 0.030455f
C1352 VTAIL.n345 VSUBS 0.030455f
C1353 VTAIL.n346 VSUBS 0.030455f
C1354 VTAIL.n347 VSUBS 0.013264f
C1355 VTAIL.n348 VSUBS 0.012885f
C1356 VTAIL.n349 VSUBS 0.023979f
C1357 VTAIL.n350 VSUBS 0.023979f
C1358 VTAIL.n351 VSUBS 0.012885f
C1359 VTAIL.n352 VSUBS 0.013643f
C1360 VTAIL.n353 VSUBS 0.030455f
C1361 VTAIL.n354 VSUBS 0.074427f
C1362 VTAIL.n355 VSUBS 0.013643f
C1363 VTAIL.n356 VSUBS 0.012885f
C1364 VTAIL.n357 VSUBS 0.060339f
C1365 VTAIL.n358 VSUBS 0.037605f
C1366 VTAIL.n359 VSUBS 1.51261f
C1367 VP.t0 VSUBS 1.71335f
C1368 VP.t1 VSUBS 1.58828f
C1369 VP.n0 VSUBS 4.68246f
.ends

