* NGSPICE file created from diff_pair_sample_0368.ext - technology: sky130A

.subckt diff_pair_sample_0368 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1324_n3436# sky130_fd_pr__pfet_01v8 ad=4.8048 pd=25.42 as=0 ps=0 w=12.32 l=0.26
X1 VTAIL.t7 VN.t0 VDD2.t3 w_n1324_n3436# sky130_fd_pr__pfet_01v8 ad=4.8048 pd=25.42 as=2.0328 ps=12.65 w=12.32 l=0.26
X2 B.t8 B.t6 B.t7 w_n1324_n3436# sky130_fd_pr__pfet_01v8 ad=4.8048 pd=25.42 as=0 ps=0 w=12.32 l=0.26
X3 VDD2.t0 VN.t1 VTAIL.t6 w_n1324_n3436# sky130_fd_pr__pfet_01v8 ad=2.0328 pd=12.65 as=4.8048 ps=25.42 w=12.32 l=0.26
X4 VDD1.t3 VP.t0 VTAIL.t1 w_n1324_n3436# sky130_fd_pr__pfet_01v8 ad=2.0328 pd=12.65 as=4.8048 ps=25.42 w=12.32 l=0.26
X5 B.t5 B.t3 B.t4 w_n1324_n3436# sky130_fd_pr__pfet_01v8 ad=4.8048 pd=25.42 as=0 ps=0 w=12.32 l=0.26
X6 VTAIL.t2 VP.t1 VDD1.t2 w_n1324_n3436# sky130_fd_pr__pfet_01v8 ad=4.8048 pd=25.42 as=2.0328 ps=12.65 w=12.32 l=0.26
X7 VTAIL.t5 VN.t2 VDD2.t2 w_n1324_n3436# sky130_fd_pr__pfet_01v8 ad=4.8048 pd=25.42 as=2.0328 ps=12.65 w=12.32 l=0.26
X8 VTAIL.t3 VP.t2 VDD1.t1 w_n1324_n3436# sky130_fd_pr__pfet_01v8 ad=4.8048 pd=25.42 as=2.0328 ps=12.65 w=12.32 l=0.26
X9 B.t2 B.t0 B.t1 w_n1324_n3436# sky130_fd_pr__pfet_01v8 ad=4.8048 pd=25.42 as=0 ps=0 w=12.32 l=0.26
X10 VDD2.t1 VN.t3 VTAIL.t4 w_n1324_n3436# sky130_fd_pr__pfet_01v8 ad=2.0328 pd=12.65 as=4.8048 ps=25.42 w=12.32 l=0.26
X11 VDD1.t0 VP.t3 VTAIL.t0 w_n1324_n3436# sky130_fd_pr__pfet_01v8 ad=2.0328 pd=12.65 as=4.8048 ps=25.42 w=12.32 l=0.26
R0 B.n104 B.t6 1364.42
R1 B.n96 B.t3 1364.42
R2 B.n38 B.t0 1364.42
R3 B.n30 B.t9 1364.42
R4 B.n294 B.n293 585
R5 B.n292 B.n75 585
R6 B.n291 B.n290 585
R7 B.n289 B.n76 585
R8 B.n288 B.n287 585
R9 B.n286 B.n77 585
R10 B.n285 B.n284 585
R11 B.n283 B.n78 585
R12 B.n282 B.n281 585
R13 B.n280 B.n79 585
R14 B.n279 B.n278 585
R15 B.n277 B.n80 585
R16 B.n276 B.n275 585
R17 B.n274 B.n81 585
R18 B.n273 B.n272 585
R19 B.n271 B.n82 585
R20 B.n270 B.n269 585
R21 B.n268 B.n83 585
R22 B.n267 B.n266 585
R23 B.n265 B.n84 585
R24 B.n264 B.n263 585
R25 B.n262 B.n85 585
R26 B.n261 B.n260 585
R27 B.n259 B.n86 585
R28 B.n258 B.n257 585
R29 B.n256 B.n87 585
R30 B.n255 B.n254 585
R31 B.n253 B.n88 585
R32 B.n252 B.n251 585
R33 B.n250 B.n89 585
R34 B.n249 B.n248 585
R35 B.n247 B.n90 585
R36 B.n246 B.n245 585
R37 B.n244 B.n91 585
R38 B.n243 B.n242 585
R39 B.n241 B.n92 585
R40 B.n240 B.n239 585
R41 B.n238 B.n93 585
R42 B.n237 B.n236 585
R43 B.n235 B.n94 585
R44 B.n234 B.n233 585
R45 B.n232 B.n95 585
R46 B.n231 B.n230 585
R47 B.n229 B.n228 585
R48 B.n227 B.n99 585
R49 B.n226 B.n225 585
R50 B.n224 B.n100 585
R51 B.n223 B.n222 585
R52 B.n221 B.n101 585
R53 B.n220 B.n219 585
R54 B.n218 B.n102 585
R55 B.n217 B.n216 585
R56 B.n214 B.n103 585
R57 B.n213 B.n212 585
R58 B.n211 B.n106 585
R59 B.n210 B.n209 585
R60 B.n208 B.n107 585
R61 B.n207 B.n206 585
R62 B.n205 B.n108 585
R63 B.n204 B.n203 585
R64 B.n202 B.n109 585
R65 B.n201 B.n200 585
R66 B.n199 B.n110 585
R67 B.n198 B.n197 585
R68 B.n196 B.n111 585
R69 B.n195 B.n194 585
R70 B.n193 B.n112 585
R71 B.n192 B.n191 585
R72 B.n190 B.n113 585
R73 B.n189 B.n188 585
R74 B.n187 B.n114 585
R75 B.n186 B.n185 585
R76 B.n184 B.n115 585
R77 B.n183 B.n182 585
R78 B.n181 B.n116 585
R79 B.n180 B.n179 585
R80 B.n178 B.n117 585
R81 B.n177 B.n176 585
R82 B.n175 B.n118 585
R83 B.n174 B.n173 585
R84 B.n172 B.n119 585
R85 B.n171 B.n170 585
R86 B.n169 B.n120 585
R87 B.n168 B.n167 585
R88 B.n166 B.n121 585
R89 B.n165 B.n164 585
R90 B.n163 B.n122 585
R91 B.n162 B.n161 585
R92 B.n160 B.n123 585
R93 B.n159 B.n158 585
R94 B.n157 B.n124 585
R95 B.n156 B.n155 585
R96 B.n154 B.n125 585
R97 B.n153 B.n152 585
R98 B.n151 B.n126 585
R99 B.n295 B.n74 585
R100 B.n297 B.n296 585
R101 B.n298 B.n73 585
R102 B.n300 B.n299 585
R103 B.n301 B.n72 585
R104 B.n303 B.n302 585
R105 B.n304 B.n71 585
R106 B.n306 B.n305 585
R107 B.n307 B.n70 585
R108 B.n309 B.n308 585
R109 B.n310 B.n69 585
R110 B.n312 B.n311 585
R111 B.n313 B.n68 585
R112 B.n315 B.n314 585
R113 B.n316 B.n67 585
R114 B.n318 B.n317 585
R115 B.n319 B.n66 585
R116 B.n321 B.n320 585
R117 B.n322 B.n65 585
R118 B.n324 B.n323 585
R119 B.n325 B.n64 585
R120 B.n327 B.n326 585
R121 B.n328 B.n63 585
R122 B.n330 B.n329 585
R123 B.n331 B.n62 585
R124 B.n333 B.n332 585
R125 B.n334 B.n61 585
R126 B.n336 B.n335 585
R127 B.n480 B.n479 585
R128 B.n478 B.n9 585
R129 B.n477 B.n476 585
R130 B.n475 B.n10 585
R131 B.n474 B.n473 585
R132 B.n472 B.n11 585
R133 B.n471 B.n470 585
R134 B.n469 B.n12 585
R135 B.n468 B.n467 585
R136 B.n466 B.n13 585
R137 B.n465 B.n464 585
R138 B.n463 B.n14 585
R139 B.n462 B.n461 585
R140 B.n460 B.n15 585
R141 B.n459 B.n458 585
R142 B.n457 B.n16 585
R143 B.n456 B.n455 585
R144 B.n454 B.n17 585
R145 B.n453 B.n452 585
R146 B.n451 B.n18 585
R147 B.n450 B.n449 585
R148 B.n448 B.n19 585
R149 B.n447 B.n446 585
R150 B.n445 B.n20 585
R151 B.n444 B.n443 585
R152 B.n442 B.n21 585
R153 B.n441 B.n440 585
R154 B.n439 B.n22 585
R155 B.n438 B.n437 585
R156 B.n436 B.n23 585
R157 B.n435 B.n434 585
R158 B.n433 B.n24 585
R159 B.n432 B.n431 585
R160 B.n430 B.n25 585
R161 B.n429 B.n428 585
R162 B.n427 B.n26 585
R163 B.n426 B.n425 585
R164 B.n424 B.n27 585
R165 B.n423 B.n422 585
R166 B.n421 B.n28 585
R167 B.n420 B.n419 585
R168 B.n418 B.n29 585
R169 B.n417 B.n416 585
R170 B.n415 B.n414 585
R171 B.n413 B.n33 585
R172 B.n412 B.n411 585
R173 B.n410 B.n34 585
R174 B.n409 B.n408 585
R175 B.n407 B.n35 585
R176 B.n406 B.n405 585
R177 B.n404 B.n36 585
R178 B.n403 B.n402 585
R179 B.n400 B.n37 585
R180 B.n399 B.n398 585
R181 B.n397 B.n40 585
R182 B.n396 B.n395 585
R183 B.n394 B.n41 585
R184 B.n393 B.n392 585
R185 B.n391 B.n42 585
R186 B.n390 B.n389 585
R187 B.n388 B.n43 585
R188 B.n387 B.n386 585
R189 B.n385 B.n44 585
R190 B.n384 B.n383 585
R191 B.n382 B.n45 585
R192 B.n381 B.n380 585
R193 B.n379 B.n46 585
R194 B.n378 B.n377 585
R195 B.n376 B.n47 585
R196 B.n375 B.n374 585
R197 B.n373 B.n48 585
R198 B.n372 B.n371 585
R199 B.n370 B.n49 585
R200 B.n369 B.n368 585
R201 B.n367 B.n50 585
R202 B.n366 B.n365 585
R203 B.n364 B.n51 585
R204 B.n363 B.n362 585
R205 B.n361 B.n52 585
R206 B.n360 B.n359 585
R207 B.n358 B.n53 585
R208 B.n357 B.n356 585
R209 B.n355 B.n54 585
R210 B.n354 B.n353 585
R211 B.n352 B.n55 585
R212 B.n351 B.n350 585
R213 B.n349 B.n56 585
R214 B.n348 B.n347 585
R215 B.n346 B.n57 585
R216 B.n345 B.n344 585
R217 B.n343 B.n58 585
R218 B.n342 B.n341 585
R219 B.n340 B.n59 585
R220 B.n339 B.n338 585
R221 B.n337 B.n60 585
R222 B.n481 B.n8 585
R223 B.n483 B.n482 585
R224 B.n484 B.n7 585
R225 B.n486 B.n485 585
R226 B.n487 B.n6 585
R227 B.n489 B.n488 585
R228 B.n490 B.n5 585
R229 B.n492 B.n491 585
R230 B.n493 B.n4 585
R231 B.n495 B.n494 585
R232 B.n496 B.n3 585
R233 B.n498 B.n497 585
R234 B.n499 B.n0 585
R235 B.n2 B.n1 585
R236 B.n133 B.n132 585
R237 B.n135 B.n134 585
R238 B.n136 B.n131 585
R239 B.n138 B.n137 585
R240 B.n139 B.n130 585
R241 B.n141 B.n140 585
R242 B.n142 B.n129 585
R243 B.n144 B.n143 585
R244 B.n145 B.n128 585
R245 B.n147 B.n146 585
R246 B.n148 B.n127 585
R247 B.n150 B.n149 585
R248 B.n151 B.n150 454.062
R249 B.n295 B.n294 454.062
R250 B.n337 B.n336 454.062
R251 B.n481 B.n480 454.062
R252 B.n501 B.n500 256.663
R253 B.n500 B.n499 235.042
R254 B.n500 B.n2 235.042
R255 B.n152 B.n151 163.367
R256 B.n152 B.n125 163.367
R257 B.n156 B.n125 163.367
R258 B.n157 B.n156 163.367
R259 B.n158 B.n157 163.367
R260 B.n158 B.n123 163.367
R261 B.n162 B.n123 163.367
R262 B.n163 B.n162 163.367
R263 B.n164 B.n163 163.367
R264 B.n164 B.n121 163.367
R265 B.n168 B.n121 163.367
R266 B.n169 B.n168 163.367
R267 B.n170 B.n169 163.367
R268 B.n170 B.n119 163.367
R269 B.n174 B.n119 163.367
R270 B.n175 B.n174 163.367
R271 B.n176 B.n175 163.367
R272 B.n176 B.n117 163.367
R273 B.n180 B.n117 163.367
R274 B.n181 B.n180 163.367
R275 B.n182 B.n181 163.367
R276 B.n182 B.n115 163.367
R277 B.n186 B.n115 163.367
R278 B.n187 B.n186 163.367
R279 B.n188 B.n187 163.367
R280 B.n188 B.n113 163.367
R281 B.n192 B.n113 163.367
R282 B.n193 B.n192 163.367
R283 B.n194 B.n193 163.367
R284 B.n194 B.n111 163.367
R285 B.n198 B.n111 163.367
R286 B.n199 B.n198 163.367
R287 B.n200 B.n199 163.367
R288 B.n200 B.n109 163.367
R289 B.n204 B.n109 163.367
R290 B.n205 B.n204 163.367
R291 B.n206 B.n205 163.367
R292 B.n206 B.n107 163.367
R293 B.n210 B.n107 163.367
R294 B.n211 B.n210 163.367
R295 B.n212 B.n211 163.367
R296 B.n212 B.n103 163.367
R297 B.n217 B.n103 163.367
R298 B.n218 B.n217 163.367
R299 B.n219 B.n218 163.367
R300 B.n219 B.n101 163.367
R301 B.n223 B.n101 163.367
R302 B.n224 B.n223 163.367
R303 B.n225 B.n224 163.367
R304 B.n225 B.n99 163.367
R305 B.n229 B.n99 163.367
R306 B.n230 B.n229 163.367
R307 B.n230 B.n95 163.367
R308 B.n234 B.n95 163.367
R309 B.n235 B.n234 163.367
R310 B.n236 B.n235 163.367
R311 B.n236 B.n93 163.367
R312 B.n240 B.n93 163.367
R313 B.n241 B.n240 163.367
R314 B.n242 B.n241 163.367
R315 B.n242 B.n91 163.367
R316 B.n246 B.n91 163.367
R317 B.n247 B.n246 163.367
R318 B.n248 B.n247 163.367
R319 B.n248 B.n89 163.367
R320 B.n252 B.n89 163.367
R321 B.n253 B.n252 163.367
R322 B.n254 B.n253 163.367
R323 B.n254 B.n87 163.367
R324 B.n258 B.n87 163.367
R325 B.n259 B.n258 163.367
R326 B.n260 B.n259 163.367
R327 B.n260 B.n85 163.367
R328 B.n264 B.n85 163.367
R329 B.n265 B.n264 163.367
R330 B.n266 B.n265 163.367
R331 B.n266 B.n83 163.367
R332 B.n270 B.n83 163.367
R333 B.n271 B.n270 163.367
R334 B.n272 B.n271 163.367
R335 B.n272 B.n81 163.367
R336 B.n276 B.n81 163.367
R337 B.n277 B.n276 163.367
R338 B.n278 B.n277 163.367
R339 B.n278 B.n79 163.367
R340 B.n282 B.n79 163.367
R341 B.n283 B.n282 163.367
R342 B.n284 B.n283 163.367
R343 B.n284 B.n77 163.367
R344 B.n288 B.n77 163.367
R345 B.n289 B.n288 163.367
R346 B.n290 B.n289 163.367
R347 B.n290 B.n75 163.367
R348 B.n294 B.n75 163.367
R349 B.n336 B.n61 163.367
R350 B.n332 B.n61 163.367
R351 B.n332 B.n331 163.367
R352 B.n331 B.n330 163.367
R353 B.n330 B.n63 163.367
R354 B.n326 B.n63 163.367
R355 B.n326 B.n325 163.367
R356 B.n325 B.n324 163.367
R357 B.n324 B.n65 163.367
R358 B.n320 B.n65 163.367
R359 B.n320 B.n319 163.367
R360 B.n319 B.n318 163.367
R361 B.n318 B.n67 163.367
R362 B.n314 B.n67 163.367
R363 B.n314 B.n313 163.367
R364 B.n313 B.n312 163.367
R365 B.n312 B.n69 163.367
R366 B.n308 B.n69 163.367
R367 B.n308 B.n307 163.367
R368 B.n307 B.n306 163.367
R369 B.n306 B.n71 163.367
R370 B.n302 B.n71 163.367
R371 B.n302 B.n301 163.367
R372 B.n301 B.n300 163.367
R373 B.n300 B.n73 163.367
R374 B.n296 B.n73 163.367
R375 B.n296 B.n295 163.367
R376 B.n480 B.n9 163.367
R377 B.n476 B.n9 163.367
R378 B.n476 B.n475 163.367
R379 B.n475 B.n474 163.367
R380 B.n474 B.n11 163.367
R381 B.n470 B.n11 163.367
R382 B.n470 B.n469 163.367
R383 B.n469 B.n468 163.367
R384 B.n468 B.n13 163.367
R385 B.n464 B.n13 163.367
R386 B.n464 B.n463 163.367
R387 B.n463 B.n462 163.367
R388 B.n462 B.n15 163.367
R389 B.n458 B.n15 163.367
R390 B.n458 B.n457 163.367
R391 B.n457 B.n456 163.367
R392 B.n456 B.n17 163.367
R393 B.n452 B.n17 163.367
R394 B.n452 B.n451 163.367
R395 B.n451 B.n450 163.367
R396 B.n450 B.n19 163.367
R397 B.n446 B.n19 163.367
R398 B.n446 B.n445 163.367
R399 B.n445 B.n444 163.367
R400 B.n444 B.n21 163.367
R401 B.n440 B.n21 163.367
R402 B.n440 B.n439 163.367
R403 B.n439 B.n438 163.367
R404 B.n438 B.n23 163.367
R405 B.n434 B.n23 163.367
R406 B.n434 B.n433 163.367
R407 B.n433 B.n432 163.367
R408 B.n432 B.n25 163.367
R409 B.n428 B.n25 163.367
R410 B.n428 B.n427 163.367
R411 B.n427 B.n426 163.367
R412 B.n426 B.n27 163.367
R413 B.n422 B.n27 163.367
R414 B.n422 B.n421 163.367
R415 B.n421 B.n420 163.367
R416 B.n420 B.n29 163.367
R417 B.n416 B.n29 163.367
R418 B.n416 B.n415 163.367
R419 B.n415 B.n33 163.367
R420 B.n411 B.n33 163.367
R421 B.n411 B.n410 163.367
R422 B.n410 B.n409 163.367
R423 B.n409 B.n35 163.367
R424 B.n405 B.n35 163.367
R425 B.n405 B.n404 163.367
R426 B.n404 B.n403 163.367
R427 B.n403 B.n37 163.367
R428 B.n398 B.n37 163.367
R429 B.n398 B.n397 163.367
R430 B.n397 B.n396 163.367
R431 B.n396 B.n41 163.367
R432 B.n392 B.n41 163.367
R433 B.n392 B.n391 163.367
R434 B.n391 B.n390 163.367
R435 B.n390 B.n43 163.367
R436 B.n386 B.n43 163.367
R437 B.n386 B.n385 163.367
R438 B.n385 B.n384 163.367
R439 B.n384 B.n45 163.367
R440 B.n380 B.n45 163.367
R441 B.n380 B.n379 163.367
R442 B.n379 B.n378 163.367
R443 B.n378 B.n47 163.367
R444 B.n374 B.n47 163.367
R445 B.n374 B.n373 163.367
R446 B.n373 B.n372 163.367
R447 B.n372 B.n49 163.367
R448 B.n368 B.n49 163.367
R449 B.n368 B.n367 163.367
R450 B.n367 B.n366 163.367
R451 B.n366 B.n51 163.367
R452 B.n362 B.n51 163.367
R453 B.n362 B.n361 163.367
R454 B.n361 B.n360 163.367
R455 B.n360 B.n53 163.367
R456 B.n356 B.n53 163.367
R457 B.n356 B.n355 163.367
R458 B.n355 B.n354 163.367
R459 B.n354 B.n55 163.367
R460 B.n350 B.n55 163.367
R461 B.n350 B.n349 163.367
R462 B.n349 B.n348 163.367
R463 B.n348 B.n57 163.367
R464 B.n344 B.n57 163.367
R465 B.n344 B.n343 163.367
R466 B.n343 B.n342 163.367
R467 B.n342 B.n59 163.367
R468 B.n338 B.n59 163.367
R469 B.n338 B.n337 163.367
R470 B.n482 B.n481 163.367
R471 B.n482 B.n7 163.367
R472 B.n486 B.n7 163.367
R473 B.n487 B.n486 163.367
R474 B.n488 B.n487 163.367
R475 B.n488 B.n5 163.367
R476 B.n492 B.n5 163.367
R477 B.n493 B.n492 163.367
R478 B.n494 B.n493 163.367
R479 B.n494 B.n3 163.367
R480 B.n498 B.n3 163.367
R481 B.n499 B.n498 163.367
R482 B.n133 B.n2 163.367
R483 B.n134 B.n133 163.367
R484 B.n134 B.n131 163.367
R485 B.n138 B.n131 163.367
R486 B.n139 B.n138 163.367
R487 B.n140 B.n139 163.367
R488 B.n140 B.n129 163.367
R489 B.n144 B.n129 163.367
R490 B.n145 B.n144 163.367
R491 B.n146 B.n145 163.367
R492 B.n146 B.n127 163.367
R493 B.n150 B.n127 163.367
R494 B.n96 B.t4 120.028
R495 B.n38 B.t2 120.028
R496 B.n104 B.t7 120.013
R497 B.n30 B.t11 120.013
R498 B.n97 B.t5 108.585
R499 B.n39 B.t1 108.585
R500 B.n105 B.t8 108.57
R501 B.n31 B.t10 108.57
R502 B.n215 B.n105 59.5399
R503 B.n98 B.n97 59.5399
R504 B.n401 B.n39 59.5399
R505 B.n32 B.n31 59.5399
R506 B.n479 B.n8 29.5029
R507 B.n335 B.n60 29.5029
R508 B.n149 B.n126 29.5029
R509 B.n293 B.n74 29.5029
R510 B B.n501 18.0485
R511 B.n105 B.n104 11.4429
R512 B.n97 B.n96 11.4429
R513 B.n39 B.n38 11.4429
R514 B.n31 B.n30 11.4429
R515 B.n483 B.n8 10.6151
R516 B.n484 B.n483 10.6151
R517 B.n485 B.n484 10.6151
R518 B.n485 B.n6 10.6151
R519 B.n489 B.n6 10.6151
R520 B.n490 B.n489 10.6151
R521 B.n491 B.n490 10.6151
R522 B.n491 B.n4 10.6151
R523 B.n495 B.n4 10.6151
R524 B.n496 B.n495 10.6151
R525 B.n497 B.n496 10.6151
R526 B.n497 B.n0 10.6151
R527 B.n479 B.n478 10.6151
R528 B.n478 B.n477 10.6151
R529 B.n477 B.n10 10.6151
R530 B.n473 B.n10 10.6151
R531 B.n473 B.n472 10.6151
R532 B.n472 B.n471 10.6151
R533 B.n471 B.n12 10.6151
R534 B.n467 B.n12 10.6151
R535 B.n467 B.n466 10.6151
R536 B.n466 B.n465 10.6151
R537 B.n465 B.n14 10.6151
R538 B.n461 B.n14 10.6151
R539 B.n461 B.n460 10.6151
R540 B.n460 B.n459 10.6151
R541 B.n459 B.n16 10.6151
R542 B.n455 B.n16 10.6151
R543 B.n455 B.n454 10.6151
R544 B.n454 B.n453 10.6151
R545 B.n453 B.n18 10.6151
R546 B.n449 B.n18 10.6151
R547 B.n449 B.n448 10.6151
R548 B.n448 B.n447 10.6151
R549 B.n447 B.n20 10.6151
R550 B.n443 B.n20 10.6151
R551 B.n443 B.n442 10.6151
R552 B.n442 B.n441 10.6151
R553 B.n441 B.n22 10.6151
R554 B.n437 B.n22 10.6151
R555 B.n437 B.n436 10.6151
R556 B.n436 B.n435 10.6151
R557 B.n435 B.n24 10.6151
R558 B.n431 B.n24 10.6151
R559 B.n431 B.n430 10.6151
R560 B.n430 B.n429 10.6151
R561 B.n429 B.n26 10.6151
R562 B.n425 B.n26 10.6151
R563 B.n425 B.n424 10.6151
R564 B.n424 B.n423 10.6151
R565 B.n423 B.n28 10.6151
R566 B.n419 B.n28 10.6151
R567 B.n419 B.n418 10.6151
R568 B.n418 B.n417 10.6151
R569 B.n414 B.n413 10.6151
R570 B.n413 B.n412 10.6151
R571 B.n412 B.n34 10.6151
R572 B.n408 B.n34 10.6151
R573 B.n408 B.n407 10.6151
R574 B.n407 B.n406 10.6151
R575 B.n406 B.n36 10.6151
R576 B.n402 B.n36 10.6151
R577 B.n400 B.n399 10.6151
R578 B.n399 B.n40 10.6151
R579 B.n395 B.n40 10.6151
R580 B.n395 B.n394 10.6151
R581 B.n394 B.n393 10.6151
R582 B.n393 B.n42 10.6151
R583 B.n389 B.n42 10.6151
R584 B.n389 B.n388 10.6151
R585 B.n388 B.n387 10.6151
R586 B.n387 B.n44 10.6151
R587 B.n383 B.n44 10.6151
R588 B.n383 B.n382 10.6151
R589 B.n382 B.n381 10.6151
R590 B.n381 B.n46 10.6151
R591 B.n377 B.n46 10.6151
R592 B.n377 B.n376 10.6151
R593 B.n376 B.n375 10.6151
R594 B.n375 B.n48 10.6151
R595 B.n371 B.n48 10.6151
R596 B.n371 B.n370 10.6151
R597 B.n370 B.n369 10.6151
R598 B.n369 B.n50 10.6151
R599 B.n365 B.n50 10.6151
R600 B.n365 B.n364 10.6151
R601 B.n364 B.n363 10.6151
R602 B.n363 B.n52 10.6151
R603 B.n359 B.n52 10.6151
R604 B.n359 B.n358 10.6151
R605 B.n358 B.n357 10.6151
R606 B.n357 B.n54 10.6151
R607 B.n353 B.n54 10.6151
R608 B.n353 B.n352 10.6151
R609 B.n352 B.n351 10.6151
R610 B.n351 B.n56 10.6151
R611 B.n347 B.n56 10.6151
R612 B.n347 B.n346 10.6151
R613 B.n346 B.n345 10.6151
R614 B.n345 B.n58 10.6151
R615 B.n341 B.n58 10.6151
R616 B.n341 B.n340 10.6151
R617 B.n340 B.n339 10.6151
R618 B.n339 B.n60 10.6151
R619 B.n335 B.n334 10.6151
R620 B.n334 B.n333 10.6151
R621 B.n333 B.n62 10.6151
R622 B.n329 B.n62 10.6151
R623 B.n329 B.n328 10.6151
R624 B.n328 B.n327 10.6151
R625 B.n327 B.n64 10.6151
R626 B.n323 B.n64 10.6151
R627 B.n323 B.n322 10.6151
R628 B.n322 B.n321 10.6151
R629 B.n321 B.n66 10.6151
R630 B.n317 B.n66 10.6151
R631 B.n317 B.n316 10.6151
R632 B.n316 B.n315 10.6151
R633 B.n315 B.n68 10.6151
R634 B.n311 B.n68 10.6151
R635 B.n311 B.n310 10.6151
R636 B.n310 B.n309 10.6151
R637 B.n309 B.n70 10.6151
R638 B.n305 B.n70 10.6151
R639 B.n305 B.n304 10.6151
R640 B.n304 B.n303 10.6151
R641 B.n303 B.n72 10.6151
R642 B.n299 B.n72 10.6151
R643 B.n299 B.n298 10.6151
R644 B.n298 B.n297 10.6151
R645 B.n297 B.n74 10.6151
R646 B.n132 B.n1 10.6151
R647 B.n135 B.n132 10.6151
R648 B.n136 B.n135 10.6151
R649 B.n137 B.n136 10.6151
R650 B.n137 B.n130 10.6151
R651 B.n141 B.n130 10.6151
R652 B.n142 B.n141 10.6151
R653 B.n143 B.n142 10.6151
R654 B.n143 B.n128 10.6151
R655 B.n147 B.n128 10.6151
R656 B.n148 B.n147 10.6151
R657 B.n149 B.n148 10.6151
R658 B.n153 B.n126 10.6151
R659 B.n154 B.n153 10.6151
R660 B.n155 B.n154 10.6151
R661 B.n155 B.n124 10.6151
R662 B.n159 B.n124 10.6151
R663 B.n160 B.n159 10.6151
R664 B.n161 B.n160 10.6151
R665 B.n161 B.n122 10.6151
R666 B.n165 B.n122 10.6151
R667 B.n166 B.n165 10.6151
R668 B.n167 B.n166 10.6151
R669 B.n167 B.n120 10.6151
R670 B.n171 B.n120 10.6151
R671 B.n172 B.n171 10.6151
R672 B.n173 B.n172 10.6151
R673 B.n173 B.n118 10.6151
R674 B.n177 B.n118 10.6151
R675 B.n178 B.n177 10.6151
R676 B.n179 B.n178 10.6151
R677 B.n179 B.n116 10.6151
R678 B.n183 B.n116 10.6151
R679 B.n184 B.n183 10.6151
R680 B.n185 B.n184 10.6151
R681 B.n185 B.n114 10.6151
R682 B.n189 B.n114 10.6151
R683 B.n190 B.n189 10.6151
R684 B.n191 B.n190 10.6151
R685 B.n191 B.n112 10.6151
R686 B.n195 B.n112 10.6151
R687 B.n196 B.n195 10.6151
R688 B.n197 B.n196 10.6151
R689 B.n197 B.n110 10.6151
R690 B.n201 B.n110 10.6151
R691 B.n202 B.n201 10.6151
R692 B.n203 B.n202 10.6151
R693 B.n203 B.n108 10.6151
R694 B.n207 B.n108 10.6151
R695 B.n208 B.n207 10.6151
R696 B.n209 B.n208 10.6151
R697 B.n209 B.n106 10.6151
R698 B.n213 B.n106 10.6151
R699 B.n214 B.n213 10.6151
R700 B.n216 B.n102 10.6151
R701 B.n220 B.n102 10.6151
R702 B.n221 B.n220 10.6151
R703 B.n222 B.n221 10.6151
R704 B.n222 B.n100 10.6151
R705 B.n226 B.n100 10.6151
R706 B.n227 B.n226 10.6151
R707 B.n228 B.n227 10.6151
R708 B.n232 B.n231 10.6151
R709 B.n233 B.n232 10.6151
R710 B.n233 B.n94 10.6151
R711 B.n237 B.n94 10.6151
R712 B.n238 B.n237 10.6151
R713 B.n239 B.n238 10.6151
R714 B.n239 B.n92 10.6151
R715 B.n243 B.n92 10.6151
R716 B.n244 B.n243 10.6151
R717 B.n245 B.n244 10.6151
R718 B.n245 B.n90 10.6151
R719 B.n249 B.n90 10.6151
R720 B.n250 B.n249 10.6151
R721 B.n251 B.n250 10.6151
R722 B.n251 B.n88 10.6151
R723 B.n255 B.n88 10.6151
R724 B.n256 B.n255 10.6151
R725 B.n257 B.n256 10.6151
R726 B.n257 B.n86 10.6151
R727 B.n261 B.n86 10.6151
R728 B.n262 B.n261 10.6151
R729 B.n263 B.n262 10.6151
R730 B.n263 B.n84 10.6151
R731 B.n267 B.n84 10.6151
R732 B.n268 B.n267 10.6151
R733 B.n269 B.n268 10.6151
R734 B.n269 B.n82 10.6151
R735 B.n273 B.n82 10.6151
R736 B.n274 B.n273 10.6151
R737 B.n275 B.n274 10.6151
R738 B.n275 B.n80 10.6151
R739 B.n279 B.n80 10.6151
R740 B.n280 B.n279 10.6151
R741 B.n281 B.n280 10.6151
R742 B.n281 B.n78 10.6151
R743 B.n285 B.n78 10.6151
R744 B.n286 B.n285 10.6151
R745 B.n287 B.n286 10.6151
R746 B.n287 B.n76 10.6151
R747 B.n291 B.n76 10.6151
R748 B.n292 B.n291 10.6151
R749 B.n293 B.n292 10.6151
R750 B.n501 B.n0 8.11757
R751 B.n501 B.n1 8.11757
R752 B.n414 B.n32 7.18099
R753 B.n402 B.n401 7.18099
R754 B.n216 B.n215 7.18099
R755 B.n228 B.n98 7.18099
R756 B.n417 B.n32 3.43465
R757 B.n401 B.n400 3.43465
R758 B.n215 B.n214 3.43465
R759 B.n231 B.n98 3.43465
R760 VN.n0 VN.t1 1307.41
R761 VN.n0 VN.t0 1307.41
R762 VN.n1 VN.t2 1307.41
R763 VN.n1 VN.t3 1307.41
R764 VN VN.n1 201.06
R765 VN VN.n0 161.351
R766 VDD2.n2 VDD2.n0 112.781
R767 VDD2.n2 VDD2.n1 76.901
R768 VDD2.n1 VDD2.t2 2.63889
R769 VDD2.n1 VDD2.t1 2.63889
R770 VDD2.n0 VDD2.t3 2.63889
R771 VDD2.n0 VDD2.t0 2.63889
R772 VDD2 VDD2.n2 0.0586897
R773 VTAIL.n5 VTAIL.t3 62.8618
R774 VTAIL.n4 VTAIL.t4 62.8618
R775 VTAIL.n3 VTAIL.t5 62.8618
R776 VTAIL.n7 VTAIL.t6 62.8607
R777 VTAIL.n0 VTAIL.t7 62.8607
R778 VTAIL.n1 VTAIL.t1 62.8607
R779 VTAIL.n2 VTAIL.t2 62.8607
R780 VTAIL.n6 VTAIL.t0 62.8606
R781 VTAIL.n7 VTAIL.n6 23.5134
R782 VTAIL.n3 VTAIL.n2 23.5134
R783 VTAIL.n4 VTAIL.n3 0.509121
R784 VTAIL.n6 VTAIL.n5 0.509121
R785 VTAIL.n2 VTAIL.n1 0.509121
R786 VTAIL.n5 VTAIL.n4 0.470328
R787 VTAIL.n1 VTAIL.n0 0.470328
R788 VTAIL VTAIL.n0 0.313
R789 VTAIL VTAIL.n7 0.196621
R790 VP.n1 VP.t0 1307.41
R791 VP.n1 VP.t1 1307.41
R792 VP.n0 VP.t2 1307.41
R793 VP.n0 VP.t3 1307.41
R794 VP.n2 VP.n0 200.679
R795 VP.n2 VP.n1 161.3
R796 VP VP.n2 0.0516364
R797 VDD1 VDD1.n1 113.305
R798 VDD1 VDD1.n0 76.9592
R799 VDD1.n0 VDD1.t1 2.63889
R800 VDD1.n0 VDD1.t0 2.63889
R801 VDD1.n1 VDD1.t2 2.63889
R802 VDD1.n1 VDD1.t3 2.63889
C0 VN VTAIL 1.423f
C1 VP VN 4.56197f
C2 B VTAIL 3.55876f
C3 VDD2 VTAIL 10.238701f
C4 w_n1324_n3436# VN 1.8221f
C5 VP B 0.923744f
C6 VP VDD2 0.246213f
C7 w_n1324_n3436# B 6.49226f
C8 w_n1324_n3436# VDD2 0.973117f
C9 VDD1 VN 0.147691f
C10 VDD1 B 0.856572f
C11 VP VTAIL 1.43711f
C12 VDD1 VDD2 0.470294f
C13 w_n1324_n3436# VTAIL 4.37921f
C14 VP w_n1324_n3436# 1.98639f
C15 VN B 0.662007f
C16 VDD2 VN 1.98075f
C17 VDD1 VTAIL 10.2001f
C18 VDD2 B 0.872061f
C19 VDD1 VP 2.07913f
C20 VDD1 w_n1324_n3436# 0.967081f
C21 VDD2 VSUBS 0.624198f
C22 VDD1 VSUBS 5.643883f
C23 VTAIL VSUBS 0.722956f
C24 VN VSUBS 4.05657f
C25 VP VSUBS 1.07711f
C26 B VSUBS 2.272499f
C27 w_n1324_n3436# VSUBS 55.973396f
C28 VDD1.t1 VSUBS 0.333185f
C29 VDD1.t0 VSUBS 0.333185f
C30 VDD1.n0 VSUBS 2.64366f
C31 VDD1.t2 VSUBS 0.333185f
C32 VDD1.t3 VSUBS 0.333185f
C33 VDD1.n1 VSUBS 3.40442f
C34 VP.t2 VSUBS 0.484331f
C35 VP.t3 VSUBS 0.484331f
C36 VP.n0 VSUBS 0.778889f
C37 VP.t1 VSUBS 0.484331f
C38 VP.t0 VSUBS 0.484331f
C39 VP.n1 VSUBS 0.39361f
C40 VP.n2 VSUBS 3.5669f
C41 VTAIL.t7 VSUBS 2.28915f
C42 VTAIL.n0 VSUBS 0.668248f
C43 VTAIL.t1 VSUBS 2.28915f
C44 VTAIL.n1 VSUBS 0.683456f
C45 VTAIL.t2 VSUBS 2.28915f
C46 VTAIL.n2 VSUBS 1.83824f
C47 VTAIL.t5 VSUBS 2.28916f
C48 VTAIL.n3 VSUBS 1.83823f
C49 VTAIL.t4 VSUBS 2.28916f
C50 VTAIL.n4 VSUBS 0.683453f
C51 VTAIL.t3 VSUBS 2.28916f
C52 VTAIL.n5 VSUBS 0.683453f
C53 VTAIL.t0 VSUBS 2.28915f
C54 VTAIL.n6 VSUBS 1.83824f
C55 VTAIL.t6 VSUBS 2.28915f
C56 VTAIL.n7 VSUBS 1.81401f
C57 VDD2.t3 VSUBS 0.279169f
C58 VDD2.t0 VSUBS 0.279169f
C59 VDD2.n0 VSUBS 2.82764f
C60 VDD2.t2 VSUBS 0.279169f
C61 VDD2.t1 VSUBS 0.279169f
C62 VDD2.n1 VSUBS 2.21463f
C63 VDD2.n2 VSUBS 3.98788f
C64 VN.t0 VSUBS 0.328884f
C65 VN.t1 VSUBS 0.328884f
C66 VN.n0 VSUBS 0.267291f
C67 VN.t2 VSUBS 0.328884f
C68 VN.t3 VSUBS 0.328884f
C69 VN.n1 VSUBS 0.535604f
C70 B.n0 VSUBS 0.007794f
C71 B.n1 VSUBS 0.007794f
C72 B.n2 VSUBS 0.011527f
C73 B.n3 VSUBS 0.008834f
C74 B.n4 VSUBS 0.008834f
C75 B.n5 VSUBS 0.008834f
C76 B.n6 VSUBS 0.008834f
C77 B.n7 VSUBS 0.008834f
C78 B.n8 VSUBS 0.018891f
C79 B.n9 VSUBS 0.008834f
C80 B.n10 VSUBS 0.008834f
C81 B.n11 VSUBS 0.008834f
C82 B.n12 VSUBS 0.008834f
C83 B.n13 VSUBS 0.008834f
C84 B.n14 VSUBS 0.008834f
C85 B.n15 VSUBS 0.008834f
C86 B.n16 VSUBS 0.008834f
C87 B.n17 VSUBS 0.008834f
C88 B.n18 VSUBS 0.008834f
C89 B.n19 VSUBS 0.008834f
C90 B.n20 VSUBS 0.008834f
C91 B.n21 VSUBS 0.008834f
C92 B.n22 VSUBS 0.008834f
C93 B.n23 VSUBS 0.008834f
C94 B.n24 VSUBS 0.008834f
C95 B.n25 VSUBS 0.008834f
C96 B.n26 VSUBS 0.008834f
C97 B.n27 VSUBS 0.008834f
C98 B.n28 VSUBS 0.008834f
C99 B.n29 VSUBS 0.008834f
C100 B.t10 VSUBS 0.508057f
C101 B.t11 VSUBS 0.514331f
C102 B.t9 VSUBS 0.157791f
C103 B.n30 VSUBS 0.117793f
C104 B.n31 VSUBS 0.078406f
C105 B.n32 VSUBS 0.020466f
C106 B.n33 VSUBS 0.008834f
C107 B.n34 VSUBS 0.008834f
C108 B.n35 VSUBS 0.008834f
C109 B.n36 VSUBS 0.008834f
C110 B.n37 VSUBS 0.008834f
C111 B.t1 VSUBS 0.508046f
C112 B.t2 VSUBS 0.514321f
C113 B.t0 VSUBS 0.157791f
C114 B.n38 VSUBS 0.117803f
C115 B.n39 VSUBS 0.078417f
C116 B.n40 VSUBS 0.008834f
C117 B.n41 VSUBS 0.008834f
C118 B.n42 VSUBS 0.008834f
C119 B.n43 VSUBS 0.008834f
C120 B.n44 VSUBS 0.008834f
C121 B.n45 VSUBS 0.008834f
C122 B.n46 VSUBS 0.008834f
C123 B.n47 VSUBS 0.008834f
C124 B.n48 VSUBS 0.008834f
C125 B.n49 VSUBS 0.008834f
C126 B.n50 VSUBS 0.008834f
C127 B.n51 VSUBS 0.008834f
C128 B.n52 VSUBS 0.008834f
C129 B.n53 VSUBS 0.008834f
C130 B.n54 VSUBS 0.008834f
C131 B.n55 VSUBS 0.008834f
C132 B.n56 VSUBS 0.008834f
C133 B.n57 VSUBS 0.008834f
C134 B.n58 VSUBS 0.008834f
C135 B.n59 VSUBS 0.008834f
C136 B.n60 VSUBS 0.019821f
C137 B.n61 VSUBS 0.008834f
C138 B.n62 VSUBS 0.008834f
C139 B.n63 VSUBS 0.008834f
C140 B.n64 VSUBS 0.008834f
C141 B.n65 VSUBS 0.008834f
C142 B.n66 VSUBS 0.008834f
C143 B.n67 VSUBS 0.008834f
C144 B.n68 VSUBS 0.008834f
C145 B.n69 VSUBS 0.008834f
C146 B.n70 VSUBS 0.008834f
C147 B.n71 VSUBS 0.008834f
C148 B.n72 VSUBS 0.008834f
C149 B.n73 VSUBS 0.008834f
C150 B.n74 VSUBS 0.020046f
C151 B.n75 VSUBS 0.008834f
C152 B.n76 VSUBS 0.008834f
C153 B.n77 VSUBS 0.008834f
C154 B.n78 VSUBS 0.008834f
C155 B.n79 VSUBS 0.008834f
C156 B.n80 VSUBS 0.008834f
C157 B.n81 VSUBS 0.008834f
C158 B.n82 VSUBS 0.008834f
C159 B.n83 VSUBS 0.008834f
C160 B.n84 VSUBS 0.008834f
C161 B.n85 VSUBS 0.008834f
C162 B.n86 VSUBS 0.008834f
C163 B.n87 VSUBS 0.008834f
C164 B.n88 VSUBS 0.008834f
C165 B.n89 VSUBS 0.008834f
C166 B.n90 VSUBS 0.008834f
C167 B.n91 VSUBS 0.008834f
C168 B.n92 VSUBS 0.008834f
C169 B.n93 VSUBS 0.008834f
C170 B.n94 VSUBS 0.008834f
C171 B.n95 VSUBS 0.008834f
C172 B.t5 VSUBS 0.508046f
C173 B.t4 VSUBS 0.514321f
C174 B.t3 VSUBS 0.157791f
C175 B.n96 VSUBS 0.117803f
C176 B.n97 VSUBS 0.078417f
C177 B.n98 VSUBS 0.020466f
C178 B.n99 VSUBS 0.008834f
C179 B.n100 VSUBS 0.008834f
C180 B.n101 VSUBS 0.008834f
C181 B.n102 VSUBS 0.008834f
C182 B.n103 VSUBS 0.008834f
C183 B.t8 VSUBS 0.508057f
C184 B.t7 VSUBS 0.514331f
C185 B.t6 VSUBS 0.157791f
C186 B.n104 VSUBS 0.117793f
C187 B.n105 VSUBS 0.078406f
C188 B.n106 VSUBS 0.008834f
C189 B.n107 VSUBS 0.008834f
C190 B.n108 VSUBS 0.008834f
C191 B.n109 VSUBS 0.008834f
C192 B.n110 VSUBS 0.008834f
C193 B.n111 VSUBS 0.008834f
C194 B.n112 VSUBS 0.008834f
C195 B.n113 VSUBS 0.008834f
C196 B.n114 VSUBS 0.008834f
C197 B.n115 VSUBS 0.008834f
C198 B.n116 VSUBS 0.008834f
C199 B.n117 VSUBS 0.008834f
C200 B.n118 VSUBS 0.008834f
C201 B.n119 VSUBS 0.008834f
C202 B.n120 VSUBS 0.008834f
C203 B.n121 VSUBS 0.008834f
C204 B.n122 VSUBS 0.008834f
C205 B.n123 VSUBS 0.008834f
C206 B.n124 VSUBS 0.008834f
C207 B.n125 VSUBS 0.008834f
C208 B.n126 VSUBS 0.019821f
C209 B.n127 VSUBS 0.008834f
C210 B.n128 VSUBS 0.008834f
C211 B.n129 VSUBS 0.008834f
C212 B.n130 VSUBS 0.008834f
C213 B.n131 VSUBS 0.008834f
C214 B.n132 VSUBS 0.008834f
C215 B.n133 VSUBS 0.008834f
C216 B.n134 VSUBS 0.008834f
C217 B.n135 VSUBS 0.008834f
C218 B.n136 VSUBS 0.008834f
C219 B.n137 VSUBS 0.008834f
C220 B.n138 VSUBS 0.008834f
C221 B.n139 VSUBS 0.008834f
C222 B.n140 VSUBS 0.008834f
C223 B.n141 VSUBS 0.008834f
C224 B.n142 VSUBS 0.008834f
C225 B.n143 VSUBS 0.008834f
C226 B.n144 VSUBS 0.008834f
C227 B.n145 VSUBS 0.008834f
C228 B.n146 VSUBS 0.008834f
C229 B.n147 VSUBS 0.008834f
C230 B.n148 VSUBS 0.008834f
C231 B.n149 VSUBS 0.018891f
C232 B.n150 VSUBS 0.018891f
C233 B.n151 VSUBS 0.019821f
C234 B.n152 VSUBS 0.008834f
C235 B.n153 VSUBS 0.008834f
C236 B.n154 VSUBS 0.008834f
C237 B.n155 VSUBS 0.008834f
C238 B.n156 VSUBS 0.008834f
C239 B.n157 VSUBS 0.008834f
C240 B.n158 VSUBS 0.008834f
C241 B.n159 VSUBS 0.008834f
C242 B.n160 VSUBS 0.008834f
C243 B.n161 VSUBS 0.008834f
C244 B.n162 VSUBS 0.008834f
C245 B.n163 VSUBS 0.008834f
C246 B.n164 VSUBS 0.008834f
C247 B.n165 VSUBS 0.008834f
C248 B.n166 VSUBS 0.008834f
C249 B.n167 VSUBS 0.008834f
C250 B.n168 VSUBS 0.008834f
C251 B.n169 VSUBS 0.008834f
C252 B.n170 VSUBS 0.008834f
C253 B.n171 VSUBS 0.008834f
C254 B.n172 VSUBS 0.008834f
C255 B.n173 VSUBS 0.008834f
C256 B.n174 VSUBS 0.008834f
C257 B.n175 VSUBS 0.008834f
C258 B.n176 VSUBS 0.008834f
C259 B.n177 VSUBS 0.008834f
C260 B.n178 VSUBS 0.008834f
C261 B.n179 VSUBS 0.008834f
C262 B.n180 VSUBS 0.008834f
C263 B.n181 VSUBS 0.008834f
C264 B.n182 VSUBS 0.008834f
C265 B.n183 VSUBS 0.008834f
C266 B.n184 VSUBS 0.008834f
C267 B.n185 VSUBS 0.008834f
C268 B.n186 VSUBS 0.008834f
C269 B.n187 VSUBS 0.008834f
C270 B.n188 VSUBS 0.008834f
C271 B.n189 VSUBS 0.008834f
C272 B.n190 VSUBS 0.008834f
C273 B.n191 VSUBS 0.008834f
C274 B.n192 VSUBS 0.008834f
C275 B.n193 VSUBS 0.008834f
C276 B.n194 VSUBS 0.008834f
C277 B.n195 VSUBS 0.008834f
C278 B.n196 VSUBS 0.008834f
C279 B.n197 VSUBS 0.008834f
C280 B.n198 VSUBS 0.008834f
C281 B.n199 VSUBS 0.008834f
C282 B.n200 VSUBS 0.008834f
C283 B.n201 VSUBS 0.008834f
C284 B.n202 VSUBS 0.008834f
C285 B.n203 VSUBS 0.008834f
C286 B.n204 VSUBS 0.008834f
C287 B.n205 VSUBS 0.008834f
C288 B.n206 VSUBS 0.008834f
C289 B.n207 VSUBS 0.008834f
C290 B.n208 VSUBS 0.008834f
C291 B.n209 VSUBS 0.008834f
C292 B.n210 VSUBS 0.008834f
C293 B.n211 VSUBS 0.008834f
C294 B.n212 VSUBS 0.008834f
C295 B.n213 VSUBS 0.008834f
C296 B.n214 VSUBS 0.005846f
C297 B.n215 VSUBS 0.020466f
C298 B.n216 VSUBS 0.007405f
C299 B.n217 VSUBS 0.008834f
C300 B.n218 VSUBS 0.008834f
C301 B.n219 VSUBS 0.008834f
C302 B.n220 VSUBS 0.008834f
C303 B.n221 VSUBS 0.008834f
C304 B.n222 VSUBS 0.008834f
C305 B.n223 VSUBS 0.008834f
C306 B.n224 VSUBS 0.008834f
C307 B.n225 VSUBS 0.008834f
C308 B.n226 VSUBS 0.008834f
C309 B.n227 VSUBS 0.008834f
C310 B.n228 VSUBS 0.007405f
C311 B.n229 VSUBS 0.008834f
C312 B.n230 VSUBS 0.008834f
C313 B.n231 VSUBS 0.005846f
C314 B.n232 VSUBS 0.008834f
C315 B.n233 VSUBS 0.008834f
C316 B.n234 VSUBS 0.008834f
C317 B.n235 VSUBS 0.008834f
C318 B.n236 VSUBS 0.008834f
C319 B.n237 VSUBS 0.008834f
C320 B.n238 VSUBS 0.008834f
C321 B.n239 VSUBS 0.008834f
C322 B.n240 VSUBS 0.008834f
C323 B.n241 VSUBS 0.008834f
C324 B.n242 VSUBS 0.008834f
C325 B.n243 VSUBS 0.008834f
C326 B.n244 VSUBS 0.008834f
C327 B.n245 VSUBS 0.008834f
C328 B.n246 VSUBS 0.008834f
C329 B.n247 VSUBS 0.008834f
C330 B.n248 VSUBS 0.008834f
C331 B.n249 VSUBS 0.008834f
C332 B.n250 VSUBS 0.008834f
C333 B.n251 VSUBS 0.008834f
C334 B.n252 VSUBS 0.008834f
C335 B.n253 VSUBS 0.008834f
C336 B.n254 VSUBS 0.008834f
C337 B.n255 VSUBS 0.008834f
C338 B.n256 VSUBS 0.008834f
C339 B.n257 VSUBS 0.008834f
C340 B.n258 VSUBS 0.008834f
C341 B.n259 VSUBS 0.008834f
C342 B.n260 VSUBS 0.008834f
C343 B.n261 VSUBS 0.008834f
C344 B.n262 VSUBS 0.008834f
C345 B.n263 VSUBS 0.008834f
C346 B.n264 VSUBS 0.008834f
C347 B.n265 VSUBS 0.008834f
C348 B.n266 VSUBS 0.008834f
C349 B.n267 VSUBS 0.008834f
C350 B.n268 VSUBS 0.008834f
C351 B.n269 VSUBS 0.008834f
C352 B.n270 VSUBS 0.008834f
C353 B.n271 VSUBS 0.008834f
C354 B.n272 VSUBS 0.008834f
C355 B.n273 VSUBS 0.008834f
C356 B.n274 VSUBS 0.008834f
C357 B.n275 VSUBS 0.008834f
C358 B.n276 VSUBS 0.008834f
C359 B.n277 VSUBS 0.008834f
C360 B.n278 VSUBS 0.008834f
C361 B.n279 VSUBS 0.008834f
C362 B.n280 VSUBS 0.008834f
C363 B.n281 VSUBS 0.008834f
C364 B.n282 VSUBS 0.008834f
C365 B.n283 VSUBS 0.008834f
C366 B.n284 VSUBS 0.008834f
C367 B.n285 VSUBS 0.008834f
C368 B.n286 VSUBS 0.008834f
C369 B.n287 VSUBS 0.008834f
C370 B.n288 VSUBS 0.008834f
C371 B.n289 VSUBS 0.008834f
C372 B.n290 VSUBS 0.008834f
C373 B.n291 VSUBS 0.008834f
C374 B.n292 VSUBS 0.008834f
C375 B.n293 VSUBS 0.018665f
C376 B.n294 VSUBS 0.019821f
C377 B.n295 VSUBS 0.018891f
C378 B.n296 VSUBS 0.008834f
C379 B.n297 VSUBS 0.008834f
C380 B.n298 VSUBS 0.008834f
C381 B.n299 VSUBS 0.008834f
C382 B.n300 VSUBS 0.008834f
C383 B.n301 VSUBS 0.008834f
C384 B.n302 VSUBS 0.008834f
C385 B.n303 VSUBS 0.008834f
C386 B.n304 VSUBS 0.008834f
C387 B.n305 VSUBS 0.008834f
C388 B.n306 VSUBS 0.008834f
C389 B.n307 VSUBS 0.008834f
C390 B.n308 VSUBS 0.008834f
C391 B.n309 VSUBS 0.008834f
C392 B.n310 VSUBS 0.008834f
C393 B.n311 VSUBS 0.008834f
C394 B.n312 VSUBS 0.008834f
C395 B.n313 VSUBS 0.008834f
C396 B.n314 VSUBS 0.008834f
C397 B.n315 VSUBS 0.008834f
C398 B.n316 VSUBS 0.008834f
C399 B.n317 VSUBS 0.008834f
C400 B.n318 VSUBS 0.008834f
C401 B.n319 VSUBS 0.008834f
C402 B.n320 VSUBS 0.008834f
C403 B.n321 VSUBS 0.008834f
C404 B.n322 VSUBS 0.008834f
C405 B.n323 VSUBS 0.008834f
C406 B.n324 VSUBS 0.008834f
C407 B.n325 VSUBS 0.008834f
C408 B.n326 VSUBS 0.008834f
C409 B.n327 VSUBS 0.008834f
C410 B.n328 VSUBS 0.008834f
C411 B.n329 VSUBS 0.008834f
C412 B.n330 VSUBS 0.008834f
C413 B.n331 VSUBS 0.008834f
C414 B.n332 VSUBS 0.008834f
C415 B.n333 VSUBS 0.008834f
C416 B.n334 VSUBS 0.008834f
C417 B.n335 VSUBS 0.018891f
C418 B.n336 VSUBS 0.018891f
C419 B.n337 VSUBS 0.019821f
C420 B.n338 VSUBS 0.008834f
C421 B.n339 VSUBS 0.008834f
C422 B.n340 VSUBS 0.008834f
C423 B.n341 VSUBS 0.008834f
C424 B.n342 VSUBS 0.008834f
C425 B.n343 VSUBS 0.008834f
C426 B.n344 VSUBS 0.008834f
C427 B.n345 VSUBS 0.008834f
C428 B.n346 VSUBS 0.008834f
C429 B.n347 VSUBS 0.008834f
C430 B.n348 VSUBS 0.008834f
C431 B.n349 VSUBS 0.008834f
C432 B.n350 VSUBS 0.008834f
C433 B.n351 VSUBS 0.008834f
C434 B.n352 VSUBS 0.008834f
C435 B.n353 VSUBS 0.008834f
C436 B.n354 VSUBS 0.008834f
C437 B.n355 VSUBS 0.008834f
C438 B.n356 VSUBS 0.008834f
C439 B.n357 VSUBS 0.008834f
C440 B.n358 VSUBS 0.008834f
C441 B.n359 VSUBS 0.008834f
C442 B.n360 VSUBS 0.008834f
C443 B.n361 VSUBS 0.008834f
C444 B.n362 VSUBS 0.008834f
C445 B.n363 VSUBS 0.008834f
C446 B.n364 VSUBS 0.008834f
C447 B.n365 VSUBS 0.008834f
C448 B.n366 VSUBS 0.008834f
C449 B.n367 VSUBS 0.008834f
C450 B.n368 VSUBS 0.008834f
C451 B.n369 VSUBS 0.008834f
C452 B.n370 VSUBS 0.008834f
C453 B.n371 VSUBS 0.008834f
C454 B.n372 VSUBS 0.008834f
C455 B.n373 VSUBS 0.008834f
C456 B.n374 VSUBS 0.008834f
C457 B.n375 VSUBS 0.008834f
C458 B.n376 VSUBS 0.008834f
C459 B.n377 VSUBS 0.008834f
C460 B.n378 VSUBS 0.008834f
C461 B.n379 VSUBS 0.008834f
C462 B.n380 VSUBS 0.008834f
C463 B.n381 VSUBS 0.008834f
C464 B.n382 VSUBS 0.008834f
C465 B.n383 VSUBS 0.008834f
C466 B.n384 VSUBS 0.008834f
C467 B.n385 VSUBS 0.008834f
C468 B.n386 VSUBS 0.008834f
C469 B.n387 VSUBS 0.008834f
C470 B.n388 VSUBS 0.008834f
C471 B.n389 VSUBS 0.008834f
C472 B.n390 VSUBS 0.008834f
C473 B.n391 VSUBS 0.008834f
C474 B.n392 VSUBS 0.008834f
C475 B.n393 VSUBS 0.008834f
C476 B.n394 VSUBS 0.008834f
C477 B.n395 VSUBS 0.008834f
C478 B.n396 VSUBS 0.008834f
C479 B.n397 VSUBS 0.008834f
C480 B.n398 VSUBS 0.008834f
C481 B.n399 VSUBS 0.008834f
C482 B.n400 VSUBS 0.005846f
C483 B.n401 VSUBS 0.020466f
C484 B.n402 VSUBS 0.007405f
C485 B.n403 VSUBS 0.008834f
C486 B.n404 VSUBS 0.008834f
C487 B.n405 VSUBS 0.008834f
C488 B.n406 VSUBS 0.008834f
C489 B.n407 VSUBS 0.008834f
C490 B.n408 VSUBS 0.008834f
C491 B.n409 VSUBS 0.008834f
C492 B.n410 VSUBS 0.008834f
C493 B.n411 VSUBS 0.008834f
C494 B.n412 VSUBS 0.008834f
C495 B.n413 VSUBS 0.008834f
C496 B.n414 VSUBS 0.007405f
C497 B.n415 VSUBS 0.008834f
C498 B.n416 VSUBS 0.008834f
C499 B.n417 VSUBS 0.005846f
C500 B.n418 VSUBS 0.008834f
C501 B.n419 VSUBS 0.008834f
C502 B.n420 VSUBS 0.008834f
C503 B.n421 VSUBS 0.008834f
C504 B.n422 VSUBS 0.008834f
C505 B.n423 VSUBS 0.008834f
C506 B.n424 VSUBS 0.008834f
C507 B.n425 VSUBS 0.008834f
C508 B.n426 VSUBS 0.008834f
C509 B.n427 VSUBS 0.008834f
C510 B.n428 VSUBS 0.008834f
C511 B.n429 VSUBS 0.008834f
C512 B.n430 VSUBS 0.008834f
C513 B.n431 VSUBS 0.008834f
C514 B.n432 VSUBS 0.008834f
C515 B.n433 VSUBS 0.008834f
C516 B.n434 VSUBS 0.008834f
C517 B.n435 VSUBS 0.008834f
C518 B.n436 VSUBS 0.008834f
C519 B.n437 VSUBS 0.008834f
C520 B.n438 VSUBS 0.008834f
C521 B.n439 VSUBS 0.008834f
C522 B.n440 VSUBS 0.008834f
C523 B.n441 VSUBS 0.008834f
C524 B.n442 VSUBS 0.008834f
C525 B.n443 VSUBS 0.008834f
C526 B.n444 VSUBS 0.008834f
C527 B.n445 VSUBS 0.008834f
C528 B.n446 VSUBS 0.008834f
C529 B.n447 VSUBS 0.008834f
C530 B.n448 VSUBS 0.008834f
C531 B.n449 VSUBS 0.008834f
C532 B.n450 VSUBS 0.008834f
C533 B.n451 VSUBS 0.008834f
C534 B.n452 VSUBS 0.008834f
C535 B.n453 VSUBS 0.008834f
C536 B.n454 VSUBS 0.008834f
C537 B.n455 VSUBS 0.008834f
C538 B.n456 VSUBS 0.008834f
C539 B.n457 VSUBS 0.008834f
C540 B.n458 VSUBS 0.008834f
C541 B.n459 VSUBS 0.008834f
C542 B.n460 VSUBS 0.008834f
C543 B.n461 VSUBS 0.008834f
C544 B.n462 VSUBS 0.008834f
C545 B.n463 VSUBS 0.008834f
C546 B.n464 VSUBS 0.008834f
C547 B.n465 VSUBS 0.008834f
C548 B.n466 VSUBS 0.008834f
C549 B.n467 VSUBS 0.008834f
C550 B.n468 VSUBS 0.008834f
C551 B.n469 VSUBS 0.008834f
C552 B.n470 VSUBS 0.008834f
C553 B.n471 VSUBS 0.008834f
C554 B.n472 VSUBS 0.008834f
C555 B.n473 VSUBS 0.008834f
C556 B.n474 VSUBS 0.008834f
C557 B.n475 VSUBS 0.008834f
C558 B.n476 VSUBS 0.008834f
C559 B.n477 VSUBS 0.008834f
C560 B.n478 VSUBS 0.008834f
C561 B.n479 VSUBS 0.019821f
C562 B.n480 VSUBS 0.019821f
C563 B.n481 VSUBS 0.018891f
C564 B.n482 VSUBS 0.008834f
C565 B.n483 VSUBS 0.008834f
C566 B.n484 VSUBS 0.008834f
C567 B.n485 VSUBS 0.008834f
C568 B.n486 VSUBS 0.008834f
C569 B.n487 VSUBS 0.008834f
C570 B.n488 VSUBS 0.008834f
C571 B.n489 VSUBS 0.008834f
C572 B.n490 VSUBS 0.008834f
C573 B.n491 VSUBS 0.008834f
C574 B.n492 VSUBS 0.008834f
C575 B.n493 VSUBS 0.008834f
C576 B.n494 VSUBS 0.008834f
C577 B.n495 VSUBS 0.008834f
C578 B.n496 VSUBS 0.008834f
C579 B.n497 VSUBS 0.008834f
C580 B.n498 VSUBS 0.008834f
C581 B.n499 VSUBS 0.011527f
C582 B.n500 VSUBS 0.01228f
C583 B.n501 VSUBS 0.024419f
.ends

