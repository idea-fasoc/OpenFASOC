* NGSPICE file created from diff_pair_sample_0301.ext - technology: sky130A

.subckt diff_pair_sample_0301 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 w_n2670_n3862# sky130_fd_pr__pfet_01v8 ad=5.6433 pd=29.72 as=5.6433 ps=29.72 w=14.47 l=3.92
X1 VDD1.t0 VP.t1 VTAIL.t3 w_n2670_n3862# sky130_fd_pr__pfet_01v8 ad=5.6433 pd=29.72 as=5.6433 ps=29.72 w=14.47 l=3.92
X2 B.t11 B.t9 B.t10 w_n2670_n3862# sky130_fd_pr__pfet_01v8 ad=5.6433 pd=29.72 as=0 ps=0 w=14.47 l=3.92
X3 VDD2.t1 VN.t0 VTAIL.t1 w_n2670_n3862# sky130_fd_pr__pfet_01v8 ad=5.6433 pd=29.72 as=5.6433 ps=29.72 w=14.47 l=3.92
X4 B.t8 B.t6 B.t7 w_n2670_n3862# sky130_fd_pr__pfet_01v8 ad=5.6433 pd=29.72 as=0 ps=0 w=14.47 l=3.92
X5 B.t5 B.t3 B.t4 w_n2670_n3862# sky130_fd_pr__pfet_01v8 ad=5.6433 pd=29.72 as=0 ps=0 w=14.47 l=3.92
X6 B.t2 B.t0 B.t1 w_n2670_n3862# sky130_fd_pr__pfet_01v8 ad=5.6433 pd=29.72 as=0 ps=0 w=14.47 l=3.92
X7 VDD2.t0 VN.t1 VTAIL.t0 w_n2670_n3862# sky130_fd_pr__pfet_01v8 ad=5.6433 pd=29.72 as=5.6433 ps=29.72 w=14.47 l=3.92
R0 VP.n0 VP.t0 174.026
R1 VP.n0 VP.t1 123.999
R2 VP VP.n0 0.621237
R3 VTAIL.n1 VTAIL.t1 60.295
R4 VTAIL.n3 VTAIL.t0 60.2948
R5 VTAIL.n0 VTAIL.t3 60.2948
R6 VTAIL.n2 VTAIL.t2 60.2948
R7 VTAIL.n1 VTAIL.n0 32.1686
R8 VTAIL.n3 VTAIL.n2 28.5048
R9 VTAIL.n2 VTAIL.n1 2.30222
R10 VTAIL VTAIL.n0 1.44447
R11 VTAIL VTAIL.n3 0.858259
R12 VDD1 VDD1.t0 121.876
R13 VDD1 VDD1.t1 77.9478
R14 B.n495 B.n494 585
R15 B.n496 B.n75 585
R16 B.n498 B.n497 585
R17 B.n499 B.n74 585
R18 B.n501 B.n500 585
R19 B.n502 B.n73 585
R20 B.n504 B.n503 585
R21 B.n505 B.n72 585
R22 B.n507 B.n506 585
R23 B.n508 B.n71 585
R24 B.n510 B.n509 585
R25 B.n511 B.n70 585
R26 B.n513 B.n512 585
R27 B.n514 B.n69 585
R28 B.n516 B.n515 585
R29 B.n517 B.n68 585
R30 B.n519 B.n518 585
R31 B.n520 B.n67 585
R32 B.n522 B.n521 585
R33 B.n523 B.n66 585
R34 B.n525 B.n524 585
R35 B.n526 B.n65 585
R36 B.n528 B.n527 585
R37 B.n529 B.n64 585
R38 B.n531 B.n530 585
R39 B.n532 B.n63 585
R40 B.n534 B.n533 585
R41 B.n535 B.n62 585
R42 B.n537 B.n536 585
R43 B.n538 B.n61 585
R44 B.n540 B.n539 585
R45 B.n541 B.n60 585
R46 B.n543 B.n542 585
R47 B.n544 B.n59 585
R48 B.n546 B.n545 585
R49 B.n547 B.n58 585
R50 B.n549 B.n548 585
R51 B.n550 B.n57 585
R52 B.n552 B.n551 585
R53 B.n553 B.n56 585
R54 B.n555 B.n554 585
R55 B.n556 B.n55 585
R56 B.n558 B.n557 585
R57 B.n559 B.n54 585
R58 B.n561 B.n560 585
R59 B.n562 B.n53 585
R60 B.n564 B.n563 585
R61 B.n565 B.n52 585
R62 B.n567 B.n566 585
R63 B.n569 B.n49 585
R64 B.n571 B.n570 585
R65 B.n572 B.n48 585
R66 B.n574 B.n573 585
R67 B.n575 B.n47 585
R68 B.n577 B.n576 585
R69 B.n578 B.n46 585
R70 B.n580 B.n579 585
R71 B.n581 B.n43 585
R72 B.n584 B.n583 585
R73 B.n585 B.n42 585
R74 B.n587 B.n586 585
R75 B.n588 B.n41 585
R76 B.n590 B.n589 585
R77 B.n591 B.n40 585
R78 B.n593 B.n592 585
R79 B.n594 B.n39 585
R80 B.n596 B.n595 585
R81 B.n597 B.n38 585
R82 B.n599 B.n598 585
R83 B.n600 B.n37 585
R84 B.n602 B.n601 585
R85 B.n603 B.n36 585
R86 B.n605 B.n604 585
R87 B.n606 B.n35 585
R88 B.n608 B.n607 585
R89 B.n609 B.n34 585
R90 B.n611 B.n610 585
R91 B.n612 B.n33 585
R92 B.n614 B.n613 585
R93 B.n615 B.n32 585
R94 B.n617 B.n616 585
R95 B.n618 B.n31 585
R96 B.n620 B.n619 585
R97 B.n621 B.n30 585
R98 B.n623 B.n622 585
R99 B.n624 B.n29 585
R100 B.n626 B.n625 585
R101 B.n627 B.n28 585
R102 B.n629 B.n628 585
R103 B.n630 B.n27 585
R104 B.n632 B.n631 585
R105 B.n633 B.n26 585
R106 B.n635 B.n634 585
R107 B.n636 B.n25 585
R108 B.n638 B.n637 585
R109 B.n639 B.n24 585
R110 B.n641 B.n640 585
R111 B.n642 B.n23 585
R112 B.n644 B.n643 585
R113 B.n645 B.n22 585
R114 B.n647 B.n646 585
R115 B.n648 B.n21 585
R116 B.n650 B.n649 585
R117 B.n651 B.n20 585
R118 B.n653 B.n652 585
R119 B.n654 B.n19 585
R120 B.n656 B.n655 585
R121 B.n493 B.n76 585
R122 B.n492 B.n491 585
R123 B.n490 B.n77 585
R124 B.n489 B.n488 585
R125 B.n487 B.n78 585
R126 B.n486 B.n485 585
R127 B.n484 B.n79 585
R128 B.n483 B.n482 585
R129 B.n481 B.n80 585
R130 B.n480 B.n479 585
R131 B.n478 B.n81 585
R132 B.n477 B.n476 585
R133 B.n475 B.n82 585
R134 B.n474 B.n473 585
R135 B.n472 B.n83 585
R136 B.n471 B.n470 585
R137 B.n469 B.n84 585
R138 B.n468 B.n467 585
R139 B.n466 B.n85 585
R140 B.n465 B.n464 585
R141 B.n463 B.n86 585
R142 B.n462 B.n461 585
R143 B.n460 B.n87 585
R144 B.n459 B.n458 585
R145 B.n457 B.n88 585
R146 B.n456 B.n455 585
R147 B.n454 B.n89 585
R148 B.n453 B.n452 585
R149 B.n451 B.n90 585
R150 B.n450 B.n449 585
R151 B.n448 B.n91 585
R152 B.n447 B.n446 585
R153 B.n445 B.n92 585
R154 B.n444 B.n443 585
R155 B.n442 B.n93 585
R156 B.n441 B.n440 585
R157 B.n439 B.n94 585
R158 B.n438 B.n437 585
R159 B.n436 B.n95 585
R160 B.n435 B.n434 585
R161 B.n433 B.n96 585
R162 B.n432 B.n431 585
R163 B.n430 B.n97 585
R164 B.n429 B.n428 585
R165 B.n427 B.n98 585
R166 B.n426 B.n425 585
R167 B.n424 B.n99 585
R168 B.n423 B.n422 585
R169 B.n421 B.n100 585
R170 B.n420 B.n419 585
R171 B.n418 B.n101 585
R172 B.n417 B.n416 585
R173 B.n415 B.n102 585
R174 B.n414 B.n413 585
R175 B.n412 B.n103 585
R176 B.n411 B.n410 585
R177 B.n409 B.n104 585
R178 B.n408 B.n407 585
R179 B.n406 B.n105 585
R180 B.n405 B.n404 585
R181 B.n403 B.n106 585
R182 B.n402 B.n401 585
R183 B.n400 B.n107 585
R184 B.n399 B.n398 585
R185 B.n397 B.n108 585
R186 B.n396 B.n395 585
R187 B.n394 B.n109 585
R188 B.n232 B.n167 585
R189 B.n234 B.n233 585
R190 B.n235 B.n166 585
R191 B.n237 B.n236 585
R192 B.n238 B.n165 585
R193 B.n240 B.n239 585
R194 B.n241 B.n164 585
R195 B.n243 B.n242 585
R196 B.n244 B.n163 585
R197 B.n246 B.n245 585
R198 B.n247 B.n162 585
R199 B.n249 B.n248 585
R200 B.n250 B.n161 585
R201 B.n252 B.n251 585
R202 B.n253 B.n160 585
R203 B.n255 B.n254 585
R204 B.n256 B.n159 585
R205 B.n258 B.n257 585
R206 B.n259 B.n158 585
R207 B.n261 B.n260 585
R208 B.n262 B.n157 585
R209 B.n264 B.n263 585
R210 B.n265 B.n156 585
R211 B.n267 B.n266 585
R212 B.n268 B.n155 585
R213 B.n270 B.n269 585
R214 B.n271 B.n154 585
R215 B.n273 B.n272 585
R216 B.n274 B.n153 585
R217 B.n276 B.n275 585
R218 B.n277 B.n152 585
R219 B.n279 B.n278 585
R220 B.n280 B.n151 585
R221 B.n282 B.n281 585
R222 B.n283 B.n150 585
R223 B.n285 B.n284 585
R224 B.n286 B.n149 585
R225 B.n288 B.n287 585
R226 B.n289 B.n148 585
R227 B.n291 B.n290 585
R228 B.n292 B.n147 585
R229 B.n294 B.n293 585
R230 B.n295 B.n146 585
R231 B.n297 B.n296 585
R232 B.n298 B.n145 585
R233 B.n300 B.n299 585
R234 B.n301 B.n144 585
R235 B.n303 B.n302 585
R236 B.n304 B.n141 585
R237 B.n307 B.n306 585
R238 B.n308 B.n140 585
R239 B.n310 B.n309 585
R240 B.n311 B.n139 585
R241 B.n313 B.n312 585
R242 B.n314 B.n138 585
R243 B.n316 B.n315 585
R244 B.n317 B.n137 585
R245 B.n319 B.n318 585
R246 B.n321 B.n320 585
R247 B.n322 B.n133 585
R248 B.n324 B.n323 585
R249 B.n325 B.n132 585
R250 B.n327 B.n326 585
R251 B.n328 B.n131 585
R252 B.n330 B.n329 585
R253 B.n331 B.n130 585
R254 B.n333 B.n332 585
R255 B.n334 B.n129 585
R256 B.n336 B.n335 585
R257 B.n337 B.n128 585
R258 B.n339 B.n338 585
R259 B.n340 B.n127 585
R260 B.n342 B.n341 585
R261 B.n343 B.n126 585
R262 B.n345 B.n344 585
R263 B.n346 B.n125 585
R264 B.n348 B.n347 585
R265 B.n349 B.n124 585
R266 B.n351 B.n350 585
R267 B.n352 B.n123 585
R268 B.n354 B.n353 585
R269 B.n355 B.n122 585
R270 B.n357 B.n356 585
R271 B.n358 B.n121 585
R272 B.n360 B.n359 585
R273 B.n361 B.n120 585
R274 B.n363 B.n362 585
R275 B.n364 B.n119 585
R276 B.n366 B.n365 585
R277 B.n367 B.n118 585
R278 B.n369 B.n368 585
R279 B.n370 B.n117 585
R280 B.n372 B.n371 585
R281 B.n373 B.n116 585
R282 B.n375 B.n374 585
R283 B.n376 B.n115 585
R284 B.n378 B.n377 585
R285 B.n379 B.n114 585
R286 B.n381 B.n380 585
R287 B.n382 B.n113 585
R288 B.n384 B.n383 585
R289 B.n385 B.n112 585
R290 B.n387 B.n386 585
R291 B.n388 B.n111 585
R292 B.n390 B.n389 585
R293 B.n391 B.n110 585
R294 B.n393 B.n392 585
R295 B.n231 B.n230 585
R296 B.n229 B.n168 585
R297 B.n228 B.n227 585
R298 B.n226 B.n169 585
R299 B.n225 B.n224 585
R300 B.n223 B.n170 585
R301 B.n222 B.n221 585
R302 B.n220 B.n171 585
R303 B.n219 B.n218 585
R304 B.n217 B.n172 585
R305 B.n216 B.n215 585
R306 B.n214 B.n173 585
R307 B.n213 B.n212 585
R308 B.n211 B.n174 585
R309 B.n210 B.n209 585
R310 B.n208 B.n175 585
R311 B.n207 B.n206 585
R312 B.n205 B.n176 585
R313 B.n204 B.n203 585
R314 B.n202 B.n177 585
R315 B.n201 B.n200 585
R316 B.n199 B.n178 585
R317 B.n198 B.n197 585
R318 B.n196 B.n179 585
R319 B.n195 B.n194 585
R320 B.n193 B.n180 585
R321 B.n192 B.n191 585
R322 B.n190 B.n181 585
R323 B.n189 B.n188 585
R324 B.n187 B.n182 585
R325 B.n186 B.n185 585
R326 B.n184 B.n183 585
R327 B.n2 B.n0 585
R328 B.n705 B.n1 585
R329 B.n704 B.n703 585
R330 B.n702 B.n3 585
R331 B.n701 B.n700 585
R332 B.n699 B.n4 585
R333 B.n698 B.n697 585
R334 B.n696 B.n5 585
R335 B.n695 B.n694 585
R336 B.n693 B.n6 585
R337 B.n692 B.n691 585
R338 B.n690 B.n7 585
R339 B.n689 B.n688 585
R340 B.n687 B.n8 585
R341 B.n686 B.n685 585
R342 B.n684 B.n9 585
R343 B.n683 B.n682 585
R344 B.n681 B.n10 585
R345 B.n680 B.n679 585
R346 B.n678 B.n11 585
R347 B.n677 B.n676 585
R348 B.n675 B.n12 585
R349 B.n674 B.n673 585
R350 B.n672 B.n13 585
R351 B.n671 B.n670 585
R352 B.n669 B.n14 585
R353 B.n668 B.n667 585
R354 B.n666 B.n15 585
R355 B.n665 B.n664 585
R356 B.n663 B.n16 585
R357 B.n662 B.n661 585
R358 B.n660 B.n17 585
R359 B.n659 B.n658 585
R360 B.n657 B.n18 585
R361 B.n707 B.n706 585
R362 B.n230 B.n167 545.355
R363 B.n657 B.n656 545.355
R364 B.n392 B.n109 545.355
R365 B.n494 B.n493 545.355
R366 B.n134 B.t9 298.396
R367 B.n142 B.t6 298.396
R368 B.n44 B.t3 298.396
R369 B.n50 B.t0 298.396
R370 B.n134 B.t11 192.75
R371 B.n50 B.t1 192.75
R372 B.n142 B.t8 192.732
R373 B.n44 B.t4 192.732
R374 B.n230 B.n229 163.367
R375 B.n229 B.n228 163.367
R376 B.n228 B.n169 163.367
R377 B.n224 B.n169 163.367
R378 B.n224 B.n223 163.367
R379 B.n223 B.n222 163.367
R380 B.n222 B.n171 163.367
R381 B.n218 B.n171 163.367
R382 B.n218 B.n217 163.367
R383 B.n217 B.n216 163.367
R384 B.n216 B.n173 163.367
R385 B.n212 B.n173 163.367
R386 B.n212 B.n211 163.367
R387 B.n211 B.n210 163.367
R388 B.n210 B.n175 163.367
R389 B.n206 B.n175 163.367
R390 B.n206 B.n205 163.367
R391 B.n205 B.n204 163.367
R392 B.n204 B.n177 163.367
R393 B.n200 B.n177 163.367
R394 B.n200 B.n199 163.367
R395 B.n199 B.n198 163.367
R396 B.n198 B.n179 163.367
R397 B.n194 B.n179 163.367
R398 B.n194 B.n193 163.367
R399 B.n193 B.n192 163.367
R400 B.n192 B.n181 163.367
R401 B.n188 B.n181 163.367
R402 B.n188 B.n187 163.367
R403 B.n187 B.n186 163.367
R404 B.n186 B.n183 163.367
R405 B.n183 B.n2 163.367
R406 B.n706 B.n2 163.367
R407 B.n706 B.n705 163.367
R408 B.n705 B.n704 163.367
R409 B.n704 B.n3 163.367
R410 B.n700 B.n3 163.367
R411 B.n700 B.n699 163.367
R412 B.n699 B.n698 163.367
R413 B.n698 B.n5 163.367
R414 B.n694 B.n5 163.367
R415 B.n694 B.n693 163.367
R416 B.n693 B.n692 163.367
R417 B.n692 B.n7 163.367
R418 B.n688 B.n7 163.367
R419 B.n688 B.n687 163.367
R420 B.n687 B.n686 163.367
R421 B.n686 B.n9 163.367
R422 B.n682 B.n9 163.367
R423 B.n682 B.n681 163.367
R424 B.n681 B.n680 163.367
R425 B.n680 B.n11 163.367
R426 B.n676 B.n11 163.367
R427 B.n676 B.n675 163.367
R428 B.n675 B.n674 163.367
R429 B.n674 B.n13 163.367
R430 B.n670 B.n13 163.367
R431 B.n670 B.n669 163.367
R432 B.n669 B.n668 163.367
R433 B.n668 B.n15 163.367
R434 B.n664 B.n15 163.367
R435 B.n664 B.n663 163.367
R436 B.n663 B.n662 163.367
R437 B.n662 B.n17 163.367
R438 B.n658 B.n17 163.367
R439 B.n658 B.n657 163.367
R440 B.n234 B.n167 163.367
R441 B.n235 B.n234 163.367
R442 B.n236 B.n235 163.367
R443 B.n236 B.n165 163.367
R444 B.n240 B.n165 163.367
R445 B.n241 B.n240 163.367
R446 B.n242 B.n241 163.367
R447 B.n242 B.n163 163.367
R448 B.n246 B.n163 163.367
R449 B.n247 B.n246 163.367
R450 B.n248 B.n247 163.367
R451 B.n248 B.n161 163.367
R452 B.n252 B.n161 163.367
R453 B.n253 B.n252 163.367
R454 B.n254 B.n253 163.367
R455 B.n254 B.n159 163.367
R456 B.n258 B.n159 163.367
R457 B.n259 B.n258 163.367
R458 B.n260 B.n259 163.367
R459 B.n260 B.n157 163.367
R460 B.n264 B.n157 163.367
R461 B.n265 B.n264 163.367
R462 B.n266 B.n265 163.367
R463 B.n266 B.n155 163.367
R464 B.n270 B.n155 163.367
R465 B.n271 B.n270 163.367
R466 B.n272 B.n271 163.367
R467 B.n272 B.n153 163.367
R468 B.n276 B.n153 163.367
R469 B.n277 B.n276 163.367
R470 B.n278 B.n277 163.367
R471 B.n278 B.n151 163.367
R472 B.n282 B.n151 163.367
R473 B.n283 B.n282 163.367
R474 B.n284 B.n283 163.367
R475 B.n284 B.n149 163.367
R476 B.n288 B.n149 163.367
R477 B.n289 B.n288 163.367
R478 B.n290 B.n289 163.367
R479 B.n290 B.n147 163.367
R480 B.n294 B.n147 163.367
R481 B.n295 B.n294 163.367
R482 B.n296 B.n295 163.367
R483 B.n296 B.n145 163.367
R484 B.n300 B.n145 163.367
R485 B.n301 B.n300 163.367
R486 B.n302 B.n301 163.367
R487 B.n302 B.n141 163.367
R488 B.n307 B.n141 163.367
R489 B.n308 B.n307 163.367
R490 B.n309 B.n308 163.367
R491 B.n309 B.n139 163.367
R492 B.n313 B.n139 163.367
R493 B.n314 B.n313 163.367
R494 B.n315 B.n314 163.367
R495 B.n315 B.n137 163.367
R496 B.n319 B.n137 163.367
R497 B.n320 B.n319 163.367
R498 B.n320 B.n133 163.367
R499 B.n324 B.n133 163.367
R500 B.n325 B.n324 163.367
R501 B.n326 B.n325 163.367
R502 B.n326 B.n131 163.367
R503 B.n330 B.n131 163.367
R504 B.n331 B.n330 163.367
R505 B.n332 B.n331 163.367
R506 B.n332 B.n129 163.367
R507 B.n336 B.n129 163.367
R508 B.n337 B.n336 163.367
R509 B.n338 B.n337 163.367
R510 B.n338 B.n127 163.367
R511 B.n342 B.n127 163.367
R512 B.n343 B.n342 163.367
R513 B.n344 B.n343 163.367
R514 B.n344 B.n125 163.367
R515 B.n348 B.n125 163.367
R516 B.n349 B.n348 163.367
R517 B.n350 B.n349 163.367
R518 B.n350 B.n123 163.367
R519 B.n354 B.n123 163.367
R520 B.n355 B.n354 163.367
R521 B.n356 B.n355 163.367
R522 B.n356 B.n121 163.367
R523 B.n360 B.n121 163.367
R524 B.n361 B.n360 163.367
R525 B.n362 B.n361 163.367
R526 B.n362 B.n119 163.367
R527 B.n366 B.n119 163.367
R528 B.n367 B.n366 163.367
R529 B.n368 B.n367 163.367
R530 B.n368 B.n117 163.367
R531 B.n372 B.n117 163.367
R532 B.n373 B.n372 163.367
R533 B.n374 B.n373 163.367
R534 B.n374 B.n115 163.367
R535 B.n378 B.n115 163.367
R536 B.n379 B.n378 163.367
R537 B.n380 B.n379 163.367
R538 B.n380 B.n113 163.367
R539 B.n384 B.n113 163.367
R540 B.n385 B.n384 163.367
R541 B.n386 B.n385 163.367
R542 B.n386 B.n111 163.367
R543 B.n390 B.n111 163.367
R544 B.n391 B.n390 163.367
R545 B.n392 B.n391 163.367
R546 B.n396 B.n109 163.367
R547 B.n397 B.n396 163.367
R548 B.n398 B.n397 163.367
R549 B.n398 B.n107 163.367
R550 B.n402 B.n107 163.367
R551 B.n403 B.n402 163.367
R552 B.n404 B.n403 163.367
R553 B.n404 B.n105 163.367
R554 B.n408 B.n105 163.367
R555 B.n409 B.n408 163.367
R556 B.n410 B.n409 163.367
R557 B.n410 B.n103 163.367
R558 B.n414 B.n103 163.367
R559 B.n415 B.n414 163.367
R560 B.n416 B.n415 163.367
R561 B.n416 B.n101 163.367
R562 B.n420 B.n101 163.367
R563 B.n421 B.n420 163.367
R564 B.n422 B.n421 163.367
R565 B.n422 B.n99 163.367
R566 B.n426 B.n99 163.367
R567 B.n427 B.n426 163.367
R568 B.n428 B.n427 163.367
R569 B.n428 B.n97 163.367
R570 B.n432 B.n97 163.367
R571 B.n433 B.n432 163.367
R572 B.n434 B.n433 163.367
R573 B.n434 B.n95 163.367
R574 B.n438 B.n95 163.367
R575 B.n439 B.n438 163.367
R576 B.n440 B.n439 163.367
R577 B.n440 B.n93 163.367
R578 B.n444 B.n93 163.367
R579 B.n445 B.n444 163.367
R580 B.n446 B.n445 163.367
R581 B.n446 B.n91 163.367
R582 B.n450 B.n91 163.367
R583 B.n451 B.n450 163.367
R584 B.n452 B.n451 163.367
R585 B.n452 B.n89 163.367
R586 B.n456 B.n89 163.367
R587 B.n457 B.n456 163.367
R588 B.n458 B.n457 163.367
R589 B.n458 B.n87 163.367
R590 B.n462 B.n87 163.367
R591 B.n463 B.n462 163.367
R592 B.n464 B.n463 163.367
R593 B.n464 B.n85 163.367
R594 B.n468 B.n85 163.367
R595 B.n469 B.n468 163.367
R596 B.n470 B.n469 163.367
R597 B.n470 B.n83 163.367
R598 B.n474 B.n83 163.367
R599 B.n475 B.n474 163.367
R600 B.n476 B.n475 163.367
R601 B.n476 B.n81 163.367
R602 B.n480 B.n81 163.367
R603 B.n481 B.n480 163.367
R604 B.n482 B.n481 163.367
R605 B.n482 B.n79 163.367
R606 B.n486 B.n79 163.367
R607 B.n487 B.n486 163.367
R608 B.n488 B.n487 163.367
R609 B.n488 B.n77 163.367
R610 B.n492 B.n77 163.367
R611 B.n493 B.n492 163.367
R612 B.n656 B.n19 163.367
R613 B.n652 B.n19 163.367
R614 B.n652 B.n651 163.367
R615 B.n651 B.n650 163.367
R616 B.n650 B.n21 163.367
R617 B.n646 B.n21 163.367
R618 B.n646 B.n645 163.367
R619 B.n645 B.n644 163.367
R620 B.n644 B.n23 163.367
R621 B.n640 B.n23 163.367
R622 B.n640 B.n639 163.367
R623 B.n639 B.n638 163.367
R624 B.n638 B.n25 163.367
R625 B.n634 B.n25 163.367
R626 B.n634 B.n633 163.367
R627 B.n633 B.n632 163.367
R628 B.n632 B.n27 163.367
R629 B.n628 B.n27 163.367
R630 B.n628 B.n627 163.367
R631 B.n627 B.n626 163.367
R632 B.n626 B.n29 163.367
R633 B.n622 B.n29 163.367
R634 B.n622 B.n621 163.367
R635 B.n621 B.n620 163.367
R636 B.n620 B.n31 163.367
R637 B.n616 B.n31 163.367
R638 B.n616 B.n615 163.367
R639 B.n615 B.n614 163.367
R640 B.n614 B.n33 163.367
R641 B.n610 B.n33 163.367
R642 B.n610 B.n609 163.367
R643 B.n609 B.n608 163.367
R644 B.n608 B.n35 163.367
R645 B.n604 B.n35 163.367
R646 B.n604 B.n603 163.367
R647 B.n603 B.n602 163.367
R648 B.n602 B.n37 163.367
R649 B.n598 B.n37 163.367
R650 B.n598 B.n597 163.367
R651 B.n597 B.n596 163.367
R652 B.n596 B.n39 163.367
R653 B.n592 B.n39 163.367
R654 B.n592 B.n591 163.367
R655 B.n591 B.n590 163.367
R656 B.n590 B.n41 163.367
R657 B.n586 B.n41 163.367
R658 B.n586 B.n585 163.367
R659 B.n585 B.n584 163.367
R660 B.n584 B.n43 163.367
R661 B.n579 B.n43 163.367
R662 B.n579 B.n578 163.367
R663 B.n578 B.n577 163.367
R664 B.n577 B.n47 163.367
R665 B.n573 B.n47 163.367
R666 B.n573 B.n572 163.367
R667 B.n572 B.n571 163.367
R668 B.n571 B.n49 163.367
R669 B.n566 B.n49 163.367
R670 B.n566 B.n565 163.367
R671 B.n565 B.n564 163.367
R672 B.n564 B.n53 163.367
R673 B.n560 B.n53 163.367
R674 B.n560 B.n559 163.367
R675 B.n559 B.n558 163.367
R676 B.n558 B.n55 163.367
R677 B.n554 B.n55 163.367
R678 B.n554 B.n553 163.367
R679 B.n553 B.n552 163.367
R680 B.n552 B.n57 163.367
R681 B.n548 B.n57 163.367
R682 B.n548 B.n547 163.367
R683 B.n547 B.n546 163.367
R684 B.n546 B.n59 163.367
R685 B.n542 B.n59 163.367
R686 B.n542 B.n541 163.367
R687 B.n541 B.n540 163.367
R688 B.n540 B.n61 163.367
R689 B.n536 B.n61 163.367
R690 B.n536 B.n535 163.367
R691 B.n535 B.n534 163.367
R692 B.n534 B.n63 163.367
R693 B.n530 B.n63 163.367
R694 B.n530 B.n529 163.367
R695 B.n529 B.n528 163.367
R696 B.n528 B.n65 163.367
R697 B.n524 B.n65 163.367
R698 B.n524 B.n523 163.367
R699 B.n523 B.n522 163.367
R700 B.n522 B.n67 163.367
R701 B.n518 B.n67 163.367
R702 B.n518 B.n517 163.367
R703 B.n517 B.n516 163.367
R704 B.n516 B.n69 163.367
R705 B.n512 B.n69 163.367
R706 B.n512 B.n511 163.367
R707 B.n511 B.n510 163.367
R708 B.n510 B.n71 163.367
R709 B.n506 B.n71 163.367
R710 B.n506 B.n505 163.367
R711 B.n505 B.n504 163.367
R712 B.n504 B.n73 163.367
R713 B.n500 B.n73 163.367
R714 B.n500 B.n499 163.367
R715 B.n499 B.n498 163.367
R716 B.n498 B.n75 163.367
R717 B.n494 B.n75 163.367
R718 B.n135 B.t10 110.325
R719 B.n51 B.t2 110.325
R720 B.n143 B.t7 110.306
R721 B.n45 B.t5 110.306
R722 B.n135 B.n134 82.4247
R723 B.n143 B.n142 82.4247
R724 B.n45 B.n44 82.4247
R725 B.n51 B.n50 82.4247
R726 B.n136 B.n135 59.5399
R727 B.n305 B.n143 59.5399
R728 B.n582 B.n45 59.5399
R729 B.n568 B.n51 59.5399
R730 B.n655 B.n18 35.4346
R731 B.n394 B.n393 35.4346
R732 B.n232 B.n231 35.4346
R733 B.n495 B.n76 35.4346
R734 B B.n707 18.0485
R735 B.n655 B.n654 10.6151
R736 B.n654 B.n653 10.6151
R737 B.n653 B.n20 10.6151
R738 B.n649 B.n20 10.6151
R739 B.n649 B.n648 10.6151
R740 B.n648 B.n647 10.6151
R741 B.n647 B.n22 10.6151
R742 B.n643 B.n22 10.6151
R743 B.n643 B.n642 10.6151
R744 B.n642 B.n641 10.6151
R745 B.n641 B.n24 10.6151
R746 B.n637 B.n24 10.6151
R747 B.n637 B.n636 10.6151
R748 B.n636 B.n635 10.6151
R749 B.n635 B.n26 10.6151
R750 B.n631 B.n26 10.6151
R751 B.n631 B.n630 10.6151
R752 B.n630 B.n629 10.6151
R753 B.n629 B.n28 10.6151
R754 B.n625 B.n28 10.6151
R755 B.n625 B.n624 10.6151
R756 B.n624 B.n623 10.6151
R757 B.n623 B.n30 10.6151
R758 B.n619 B.n30 10.6151
R759 B.n619 B.n618 10.6151
R760 B.n618 B.n617 10.6151
R761 B.n617 B.n32 10.6151
R762 B.n613 B.n32 10.6151
R763 B.n613 B.n612 10.6151
R764 B.n612 B.n611 10.6151
R765 B.n611 B.n34 10.6151
R766 B.n607 B.n34 10.6151
R767 B.n607 B.n606 10.6151
R768 B.n606 B.n605 10.6151
R769 B.n605 B.n36 10.6151
R770 B.n601 B.n36 10.6151
R771 B.n601 B.n600 10.6151
R772 B.n600 B.n599 10.6151
R773 B.n599 B.n38 10.6151
R774 B.n595 B.n38 10.6151
R775 B.n595 B.n594 10.6151
R776 B.n594 B.n593 10.6151
R777 B.n593 B.n40 10.6151
R778 B.n589 B.n40 10.6151
R779 B.n589 B.n588 10.6151
R780 B.n588 B.n587 10.6151
R781 B.n587 B.n42 10.6151
R782 B.n583 B.n42 10.6151
R783 B.n581 B.n580 10.6151
R784 B.n580 B.n46 10.6151
R785 B.n576 B.n46 10.6151
R786 B.n576 B.n575 10.6151
R787 B.n575 B.n574 10.6151
R788 B.n574 B.n48 10.6151
R789 B.n570 B.n48 10.6151
R790 B.n570 B.n569 10.6151
R791 B.n567 B.n52 10.6151
R792 B.n563 B.n52 10.6151
R793 B.n563 B.n562 10.6151
R794 B.n562 B.n561 10.6151
R795 B.n561 B.n54 10.6151
R796 B.n557 B.n54 10.6151
R797 B.n557 B.n556 10.6151
R798 B.n556 B.n555 10.6151
R799 B.n555 B.n56 10.6151
R800 B.n551 B.n56 10.6151
R801 B.n551 B.n550 10.6151
R802 B.n550 B.n549 10.6151
R803 B.n549 B.n58 10.6151
R804 B.n545 B.n58 10.6151
R805 B.n545 B.n544 10.6151
R806 B.n544 B.n543 10.6151
R807 B.n543 B.n60 10.6151
R808 B.n539 B.n60 10.6151
R809 B.n539 B.n538 10.6151
R810 B.n538 B.n537 10.6151
R811 B.n537 B.n62 10.6151
R812 B.n533 B.n62 10.6151
R813 B.n533 B.n532 10.6151
R814 B.n532 B.n531 10.6151
R815 B.n531 B.n64 10.6151
R816 B.n527 B.n64 10.6151
R817 B.n527 B.n526 10.6151
R818 B.n526 B.n525 10.6151
R819 B.n525 B.n66 10.6151
R820 B.n521 B.n66 10.6151
R821 B.n521 B.n520 10.6151
R822 B.n520 B.n519 10.6151
R823 B.n519 B.n68 10.6151
R824 B.n515 B.n68 10.6151
R825 B.n515 B.n514 10.6151
R826 B.n514 B.n513 10.6151
R827 B.n513 B.n70 10.6151
R828 B.n509 B.n70 10.6151
R829 B.n509 B.n508 10.6151
R830 B.n508 B.n507 10.6151
R831 B.n507 B.n72 10.6151
R832 B.n503 B.n72 10.6151
R833 B.n503 B.n502 10.6151
R834 B.n502 B.n501 10.6151
R835 B.n501 B.n74 10.6151
R836 B.n497 B.n74 10.6151
R837 B.n497 B.n496 10.6151
R838 B.n496 B.n495 10.6151
R839 B.n395 B.n394 10.6151
R840 B.n395 B.n108 10.6151
R841 B.n399 B.n108 10.6151
R842 B.n400 B.n399 10.6151
R843 B.n401 B.n400 10.6151
R844 B.n401 B.n106 10.6151
R845 B.n405 B.n106 10.6151
R846 B.n406 B.n405 10.6151
R847 B.n407 B.n406 10.6151
R848 B.n407 B.n104 10.6151
R849 B.n411 B.n104 10.6151
R850 B.n412 B.n411 10.6151
R851 B.n413 B.n412 10.6151
R852 B.n413 B.n102 10.6151
R853 B.n417 B.n102 10.6151
R854 B.n418 B.n417 10.6151
R855 B.n419 B.n418 10.6151
R856 B.n419 B.n100 10.6151
R857 B.n423 B.n100 10.6151
R858 B.n424 B.n423 10.6151
R859 B.n425 B.n424 10.6151
R860 B.n425 B.n98 10.6151
R861 B.n429 B.n98 10.6151
R862 B.n430 B.n429 10.6151
R863 B.n431 B.n430 10.6151
R864 B.n431 B.n96 10.6151
R865 B.n435 B.n96 10.6151
R866 B.n436 B.n435 10.6151
R867 B.n437 B.n436 10.6151
R868 B.n437 B.n94 10.6151
R869 B.n441 B.n94 10.6151
R870 B.n442 B.n441 10.6151
R871 B.n443 B.n442 10.6151
R872 B.n443 B.n92 10.6151
R873 B.n447 B.n92 10.6151
R874 B.n448 B.n447 10.6151
R875 B.n449 B.n448 10.6151
R876 B.n449 B.n90 10.6151
R877 B.n453 B.n90 10.6151
R878 B.n454 B.n453 10.6151
R879 B.n455 B.n454 10.6151
R880 B.n455 B.n88 10.6151
R881 B.n459 B.n88 10.6151
R882 B.n460 B.n459 10.6151
R883 B.n461 B.n460 10.6151
R884 B.n461 B.n86 10.6151
R885 B.n465 B.n86 10.6151
R886 B.n466 B.n465 10.6151
R887 B.n467 B.n466 10.6151
R888 B.n467 B.n84 10.6151
R889 B.n471 B.n84 10.6151
R890 B.n472 B.n471 10.6151
R891 B.n473 B.n472 10.6151
R892 B.n473 B.n82 10.6151
R893 B.n477 B.n82 10.6151
R894 B.n478 B.n477 10.6151
R895 B.n479 B.n478 10.6151
R896 B.n479 B.n80 10.6151
R897 B.n483 B.n80 10.6151
R898 B.n484 B.n483 10.6151
R899 B.n485 B.n484 10.6151
R900 B.n485 B.n78 10.6151
R901 B.n489 B.n78 10.6151
R902 B.n490 B.n489 10.6151
R903 B.n491 B.n490 10.6151
R904 B.n491 B.n76 10.6151
R905 B.n233 B.n232 10.6151
R906 B.n233 B.n166 10.6151
R907 B.n237 B.n166 10.6151
R908 B.n238 B.n237 10.6151
R909 B.n239 B.n238 10.6151
R910 B.n239 B.n164 10.6151
R911 B.n243 B.n164 10.6151
R912 B.n244 B.n243 10.6151
R913 B.n245 B.n244 10.6151
R914 B.n245 B.n162 10.6151
R915 B.n249 B.n162 10.6151
R916 B.n250 B.n249 10.6151
R917 B.n251 B.n250 10.6151
R918 B.n251 B.n160 10.6151
R919 B.n255 B.n160 10.6151
R920 B.n256 B.n255 10.6151
R921 B.n257 B.n256 10.6151
R922 B.n257 B.n158 10.6151
R923 B.n261 B.n158 10.6151
R924 B.n262 B.n261 10.6151
R925 B.n263 B.n262 10.6151
R926 B.n263 B.n156 10.6151
R927 B.n267 B.n156 10.6151
R928 B.n268 B.n267 10.6151
R929 B.n269 B.n268 10.6151
R930 B.n269 B.n154 10.6151
R931 B.n273 B.n154 10.6151
R932 B.n274 B.n273 10.6151
R933 B.n275 B.n274 10.6151
R934 B.n275 B.n152 10.6151
R935 B.n279 B.n152 10.6151
R936 B.n280 B.n279 10.6151
R937 B.n281 B.n280 10.6151
R938 B.n281 B.n150 10.6151
R939 B.n285 B.n150 10.6151
R940 B.n286 B.n285 10.6151
R941 B.n287 B.n286 10.6151
R942 B.n287 B.n148 10.6151
R943 B.n291 B.n148 10.6151
R944 B.n292 B.n291 10.6151
R945 B.n293 B.n292 10.6151
R946 B.n293 B.n146 10.6151
R947 B.n297 B.n146 10.6151
R948 B.n298 B.n297 10.6151
R949 B.n299 B.n298 10.6151
R950 B.n299 B.n144 10.6151
R951 B.n303 B.n144 10.6151
R952 B.n304 B.n303 10.6151
R953 B.n306 B.n140 10.6151
R954 B.n310 B.n140 10.6151
R955 B.n311 B.n310 10.6151
R956 B.n312 B.n311 10.6151
R957 B.n312 B.n138 10.6151
R958 B.n316 B.n138 10.6151
R959 B.n317 B.n316 10.6151
R960 B.n318 B.n317 10.6151
R961 B.n322 B.n321 10.6151
R962 B.n323 B.n322 10.6151
R963 B.n323 B.n132 10.6151
R964 B.n327 B.n132 10.6151
R965 B.n328 B.n327 10.6151
R966 B.n329 B.n328 10.6151
R967 B.n329 B.n130 10.6151
R968 B.n333 B.n130 10.6151
R969 B.n334 B.n333 10.6151
R970 B.n335 B.n334 10.6151
R971 B.n335 B.n128 10.6151
R972 B.n339 B.n128 10.6151
R973 B.n340 B.n339 10.6151
R974 B.n341 B.n340 10.6151
R975 B.n341 B.n126 10.6151
R976 B.n345 B.n126 10.6151
R977 B.n346 B.n345 10.6151
R978 B.n347 B.n346 10.6151
R979 B.n347 B.n124 10.6151
R980 B.n351 B.n124 10.6151
R981 B.n352 B.n351 10.6151
R982 B.n353 B.n352 10.6151
R983 B.n353 B.n122 10.6151
R984 B.n357 B.n122 10.6151
R985 B.n358 B.n357 10.6151
R986 B.n359 B.n358 10.6151
R987 B.n359 B.n120 10.6151
R988 B.n363 B.n120 10.6151
R989 B.n364 B.n363 10.6151
R990 B.n365 B.n364 10.6151
R991 B.n365 B.n118 10.6151
R992 B.n369 B.n118 10.6151
R993 B.n370 B.n369 10.6151
R994 B.n371 B.n370 10.6151
R995 B.n371 B.n116 10.6151
R996 B.n375 B.n116 10.6151
R997 B.n376 B.n375 10.6151
R998 B.n377 B.n376 10.6151
R999 B.n377 B.n114 10.6151
R1000 B.n381 B.n114 10.6151
R1001 B.n382 B.n381 10.6151
R1002 B.n383 B.n382 10.6151
R1003 B.n383 B.n112 10.6151
R1004 B.n387 B.n112 10.6151
R1005 B.n388 B.n387 10.6151
R1006 B.n389 B.n388 10.6151
R1007 B.n389 B.n110 10.6151
R1008 B.n393 B.n110 10.6151
R1009 B.n231 B.n168 10.6151
R1010 B.n227 B.n168 10.6151
R1011 B.n227 B.n226 10.6151
R1012 B.n226 B.n225 10.6151
R1013 B.n225 B.n170 10.6151
R1014 B.n221 B.n170 10.6151
R1015 B.n221 B.n220 10.6151
R1016 B.n220 B.n219 10.6151
R1017 B.n219 B.n172 10.6151
R1018 B.n215 B.n172 10.6151
R1019 B.n215 B.n214 10.6151
R1020 B.n214 B.n213 10.6151
R1021 B.n213 B.n174 10.6151
R1022 B.n209 B.n174 10.6151
R1023 B.n209 B.n208 10.6151
R1024 B.n208 B.n207 10.6151
R1025 B.n207 B.n176 10.6151
R1026 B.n203 B.n176 10.6151
R1027 B.n203 B.n202 10.6151
R1028 B.n202 B.n201 10.6151
R1029 B.n201 B.n178 10.6151
R1030 B.n197 B.n178 10.6151
R1031 B.n197 B.n196 10.6151
R1032 B.n196 B.n195 10.6151
R1033 B.n195 B.n180 10.6151
R1034 B.n191 B.n180 10.6151
R1035 B.n191 B.n190 10.6151
R1036 B.n190 B.n189 10.6151
R1037 B.n189 B.n182 10.6151
R1038 B.n185 B.n182 10.6151
R1039 B.n185 B.n184 10.6151
R1040 B.n184 B.n0 10.6151
R1041 B.n703 B.n1 10.6151
R1042 B.n703 B.n702 10.6151
R1043 B.n702 B.n701 10.6151
R1044 B.n701 B.n4 10.6151
R1045 B.n697 B.n4 10.6151
R1046 B.n697 B.n696 10.6151
R1047 B.n696 B.n695 10.6151
R1048 B.n695 B.n6 10.6151
R1049 B.n691 B.n6 10.6151
R1050 B.n691 B.n690 10.6151
R1051 B.n690 B.n689 10.6151
R1052 B.n689 B.n8 10.6151
R1053 B.n685 B.n8 10.6151
R1054 B.n685 B.n684 10.6151
R1055 B.n684 B.n683 10.6151
R1056 B.n683 B.n10 10.6151
R1057 B.n679 B.n10 10.6151
R1058 B.n679 B.n678 10.6151
R1059 B.n678 B.n677 10.6151
R1060 B.n677 B.n12 10.6151
R1061 B.n673 B.n12 10.6151
R1062 B.n673 B.n672 10.6151
R1063 B.n672 B.n671 10.6151
R1064 B.n671 B.n14 10.6151
R1065 B.n667 B.n14 10.6151
R1066 B.n667 B.n666 10.6151
R1067 B.n666 B.n665 10.6151
R1068 B.n665 B.n16 10.6151
R1069 B.n661 B.n16 10.6151
R1070 B.n661 B.n660 10.6151
R1071 B.n660 B.n659 10.6151
R1072 B.n659 B.n18 10.6151
R1073 B.n582 B.n581 6.5566
R1074 B.n569 B.n568 6.5566
R1075 B.n306 B.n305 6.5566
R1076 B.n318 B.n136 6.5566
R1077 B.n583 B.n582 4.05904
R1078 B.n568 B.n567 4.05904
R1079 B.n305 B.n304 4.05904
R1080 B.n321 B.n136 4.05904
R1081 B.n707 B.n0 2.81026
R1082 B.n707 B.n1 2.81026
R1083 VN VN.t0 173.839
R1084 VN VN.t1 124.62
R1085 VDD2.n0 VDD2.t0 120.434
R1086 VDD2.n0 VDD2.t1 76.9736
R1087 VDD2 VDD2.n0 0.974638
C0 w_n2670_n3862# VDD1 2.09403f
C1 B VN 1.3007f
C2 VTAIL VN 3.10884f
C3 VDD2 VP 0.387878f
C4 B VDD2 2.12033f
C5 VP VDD1 3.71873f
C6 w_n2670_n3862# VP 4.20108f
C7 VTAIL VDD2 6.01674f
C8 B VDD1 2.07838f
C9 B w_n2670_n3862# 10.9275f
C10 VTAIL VDD1 5.95662f
C11 VTAIL w_n2670_n3862# 3.11065f
C12 VDD2 VN 3.48112f
C13 VDD1 VN 0.148729f
C14 w_n2670_n3862# VN 3.85813f
C15 B VP 1.86983f
C16 VTAIL VP 3.12388f
C17 VDD2 VDD1 0.823385f
C18 VTAIL B 4.72382f
C19 w_n2670_n3862# VDD2 2.13615f
C20 VP VN 6.53288f
C21 VDD2 VSUBS 1.174351f
C22 VDD1 VSUBS 6.94738f
C23 VTAIL VSUBS 1.232913f
C24 VN VSUBS 8.73482f
C25 VP VSUBS 2.162678f
C26 B VSUBS 5.086574f
C27 w_n2670_n3862# VSUBS 0.126526p
C28 VDD2.t0 VSUBS 4.522141f
C29 VDD2.t1 VSUBS 3.53576f
C30 VDD2.n0 VSUBS 5.37652f
C31 VN.t1 VSUBS 5.20537f
C32 VN.t0 VSUBS 6.13509f
C33 B.n0 VSUBS 0.004158f
C34 B.n1 VSUBS 0.004158f
C35 B.n2 VSUBS 0.006576f
C36 B.n3 VSUBS 0.006576f
C37 B.n4 VSUBS 0.006576f
C38 B.n5 VSUBS 0.006576f
C39 B.n6 VSUBS 0.006576f
C40 B.n7 VSUBS 0.006576f
C41 B.n8 VSUBS 0.006576f
C42 B.n9 VSUBS 0.006576f
C43 B.n10 VSUBS 0.006576f
C44 B.n11 VSUBS 0.006576f
C45 B.n12 VSUBS 0.006576f
C46 B.n13 VSUBS 0.006576f
C47 B.n14 VSUBS 0.006576f
C48 B.n15 VSUBS 0.006576f
C49 B.n16 VSUBS 0.006576f
C50 B.n17 VSUBS 0.006576f
C51 B.n18 VSUBS 0.01594f
C52 B.n19 VSUBS 0.006576f
C53 B.n20 VSUBS 0.006576f
C54 B.n21 VSUBS 0.006576f
C55 B.n22 VSUBS 0.006576f
C56 B.n23 VSUBS 0.006576f
C57 B.n24 VSUBS 0.006576f
C58 B.n25 VSUBS 0.006576f
C59 B.n26 VSUBS 0.006576f
C60 B.n27 VSUBS 0.006576f
C61 B.n28 VSUBS 0.006576f
C62 B.n29 VSUBS 0.006576f
C63 B.n30 VSUBS 0.006576f
C64 B.n31 VSUBS 0.006576f
C65 B.n32 VSUBS 0.006576f
C66 B.n33 VSUBS 0.006576f
C67 B.n34 VSUBS 0.006576f
C68 B.n35 VSUBS 0.006576f
C69 B.n36 VSUBS 0.006576f
C70 B.n37 VSUBS 0.006576f
C71 B.n38 VSUBS 0.006576f
C72 B.n39 VSUBS 0.006576f
C73 B.n40 VSUBS 0.006576f
C74 B.n41 VSUBS 0.006576f
C75 B.n42 VSUBS 0.006576f
C76 B.n43 VSUBS 0.006576f
C77 B.t5 VSUBS 0.451119f
C78 B.t4 VSUBS 0.478207f
C79 B.t3 VSUBS 2.46449f
C80 B.n44 VSUBS 0.285701f
C81 B.n45 VSUBS 0.072719f
C82 B.n46 VSUBS 0.006576f
C83 B.n47 VSUBS 0.006576f
C84 B.n48 VSUBS 0.006576f
C85 B.n49 VSUBS 0.006576f
C86 B.t2 VSUBS 0.451107f
C87 B.t1 VSUBS 0.478198f
C88 B.t0 VSUBS 2.46449f
C89 B.n50 VSUBS 0.28571f
C90 B.n51 VSUBS 0.07273f
C91 B.n52 VSUBS 0.006576f
C92 B.n53 VSUBS 0.006576f
C93 B.n54 VSUBS 0.006576f
C94 B.n55 VSUBS 0.006576f
C95 B.n56 VSUBS 0.006576f
C96 B.n57 VSUBS 0.006576f
C97 B.n58 VSUBS 0.006576f
C98 B.n59 VSUBS 0.006576f
C99 B.n60 VSUBS 0.006576f
C100 B.n61 VSUBS 0.006576f
C101 B.n62 VSUBS 0.006576f
C102 B.n63 VSUBS 0.006576f
C103 B.n64 VSUBS 0.006576f
C104 B.n65 VSUBS 0.006576f
C105 B.n66 VSUBS 0.006576f
C106 B.n67 VSUBS 0.006576f
C107 B.n68 VSUBS 0.006576f
C108 B.n69 VSUBS 0.006576f
C109 B.n70 VSUBS 0.006576f
C110 B.n71 VSUBS 0.006576f
C111 B.n72 VSUBS 0.006576f
C112 B.n73 VSUBS 0.006576f
C113 B.n74 VSUBS 0.006576f
C114 B.n75 VSUBS 0.006576f
C115 B.n76 VSUBS 0.016657f
C116 B.n77 VSUBS 0.006576f
C117 B.n78 VSUBS 0.006576f
C118 B.n79 VSUBS 0.006576f
C119 B.n80 VSUBS 0.006576f
C120 B.n81 VSUBS 0.006576f
C121 B.n82 VSUBS 0.006576f
C122 B.n83 VSUBS 0.006576f
C123 B.n84 VSUBS 0.006576f
C124 B.n85 VSUBS 0.006576f
C125 B.n86 VSUBS 0.006576f
C126 B.n87 VSUBS 0.006576f
C127 B.n88 VSUBS 0.006576f
C128 B.n89 VSUBS 0.006576f
C129 B.n90 VSUBS 0.006576f
C130 B.n91 VSUBS 0.006576f
C131 B.n92 VSUBS 0.006576f
C132 B.n93 VSUBS 0.006576f
C133 B.n94 VSUBS 0.006576f
C134 B.n95 VSUBS 0.006576f
C135 B.n96 VSUBS 0.006576f
C136 B.n97 VSUBS 0.006576f
C137 B.n98 VSUBS 0.006576f
C138 B.n99 VSUBS 0.006576f
C139 B.n100 VSUBS 0.006576f
C140 B.n101 VSUBS 0.006576f
C141 B.n102 VSUBS 0.006576f
C142 B.n103 VSUBS 0.006576f
C143 B.n104 VSUBS 0.006576f
C144 B.n105 VSUBS 0.006576f
C145 B.n106 VSUBS 0.006576f
C146 B.n107 VSUBS 0.006576f
C147 B.n108 VSUBS 0.006576f
C148 B.n109 VSUBS 0.01594f
C149 B.n110 VSUBS 0.006576f
C150 B.n111 VSUBS 0.006576f
C151 B.n112 VSUBS 0.006576f
C152 B.n113 VSUBS 0.006576f
C153 B.n114 VSUBS 0.006576f
C154 B.n115 VSUBS 0.006576f
C155 B.n116 VSUBS 0.006576f
C156 B.n117 VSUBS 0.006576f
C157 B.n118 VSUBS 0.006576f
C158 B.n119 VSUBS 0.006576f
C159 B.n120 VSUBS 0.006576f
C160 B.n121 VSUBS 0.006576f
C161 B.n122 VSUBS 0.006576f
C162 B.n123 VSUBS 0.006576f
C163 B.n124 VSUBS 0.006576f
C164 B.n125 VSUBS 0.006576f
C165 B.n126 VSUBS 0.006576f
C166 B.n127 VSUBS 0.006576f
C167 B.n128 VSUBS 0.006576f
C168 B.n129 VSUBS 0.006576f
C169 B.n130 VSUBS 0.006576f
C170 B.n131 VSUBS 0.006576f
C171 B.n132 VSUBS 0.006576f
C172 B.n133 VSUBS 0.006576f
C173 B.t10 VSUBS 0.451107f
C174 B.t11 VSUBS 0.478198f
C175 B.t9 VSUBS 2.46449f
C176 B.n134 VSUBS 0.28571f
C177 B.n135 VSUBS 0.07273f
C178 B.n136 VSUBS 0.015235f
C179 B.n137 VSUBS 0.006576f
C180 B.n138 VSUBS 0.006576f
C181 B.n139 VSUBS 0.006576f
C182 B.n140 VSUBS 0.006576f
C183 B.n141 VSUBS 0.006576f
C184 B.t7 VSUBS 0.451119f
C185 B.t8 VSUBS 0.478207f
C186 B.t6 VSUBS 2.46449f
C187 B.n142 VSUBS 0.285701f
C188 B.n143 VSUBS 0.072719f
C189 B.n144 VSUBS 0.006576f
C190 B.n145 VSUBS 0.006576f
C191 B.n146 VSUBS 0.006576f
C192 B.n147 VSUBS 0.006576f
C193 B.n148 VSUBS 0.006576f
C194 B.n149 VSUBS 0.006576f
C195 B.n150 VSUBS 0.006576f
C196 B.n151 VSUBS 0.006576f
C197 B.n152 VSUBS 0.006576f
C198 B.n153 VSUBS 0.006576f
C199 B.n154 VSUBS 0.006576f
C200 B.n155 VSUBS 0.006576f
C201 B.n156 VSUBS 0.006576f
C202 B.n157 VSUBS 0.006576f
C203 B.n158 VSUBS 0.006576f
C204 B.n159 VSUBS 0.006576f
C205 B.n160 VSUBS 0.006576f
C206 B.n161 VSUBS 0.006576f
C207 B.n162 VSUBS 0.006576f
C208 B.n163 VSUBS 0.006576f
C209 B.n164 VSUBS 0.006576f
C210 B.n165 VSUBS 0.006576f
C211 B.n166 VSUBS 0.006576f
C212 B.n167 VSUBS 0.016552f
C213 B.n168 VSUBS 0.006576f
C214 B.n169 VSUBS 0.006576f
C215 B.n170 VSUBS 0.006576f
C216 B.n171 VSUBS 0.006576f
C217 B.n172 VSUBS 0.006576f
C218 B.n173 VSUBS 0.006576f
C219 B.n174 VSUBS 0.006576f
C220 B.n175 VSUBS 0.006576f
C221 B.n176 VSUBS 0.006576f
C222 B.n177 VSUBS 0.006576f
C223 B.n178 VSUBS 0.006576f
C224 B.n179 VSUBS 0.006576f
C225 B.n180 VSUBS 0.006576f
C226 B.n181 VSUBS 0.006576f
C227 B.n182 VSUBS 0.006576f
C228 B.n183 VSUBS 0.006576f
C229 B.n184 VSUBS 0.006576f
C230 B.n185 VSUBS 0.006576f
C231 B.n186 VSUBS 0.006576f
C232 B.n187 VSUBS 0.006576f
C233 B.n188 VSUBS 0.006576f
C234 B.n189 VSUBS 0.006576f
C235 B.n190 VSUBS 0.006576f
C236 B.n191 VSUBS 0.006576f
C237 B.n192 VSUBS 0.006576f
C238 B.n193 VSUBS 0.006576f
C239 B.n194 VSUBS 0.006576f
C240 B.n195 VSUBS 0.006576f
C241 B.n196 VSUBS 0.006576f
C242 B.n197 VSUBS 0.006576f
C243 B.n198 VSUBS 0.006576f
C244 B.n199 VSUBS 0.006576f
C245 B.n200 VSUBS 0.006576f
C246 B.n201 VSUBS 0.006576f
C247 B.n202 VSUBS 0.006576f
C248 B.n203 VSUBS 0.006576f
C249 B.n204 VSUBS 0.006576f
C250 B.n205 VSUBS 0.006576f
C251 B.n206 VSUBS 0.006576f
C252 B.n207 VSUBS 0.006576f
C253 B.n208 VSUBS 0.006576f
C254 B.n209 VSUBS 0.006576f
C255 B.n210 VSUBS 0.006576f
C256 B.n211 VSUBS 0.006576f
C257 B.n212 VSUBS 0.006576f
C258 B.n213 VSUBS 0.006576f
C259 B.n214 VSUBS 0.006576f
C260 B.n215 VSUBS 0.006576f
C261 B.n216 VSUBS 0.006576f
C262 B.n217 VSUBS 0.006576f
C263 B.n218 VSUBS 0.006576f
C264 B.n219 VSUBS 0.006576f
C265 B.n220 VSUBS 0.006576f
C266 B.n221 VSUBS 0.006576f
C267 B.n222 VSUBS 0.006576f
C268 B.n223 VSUBS 0.006576f
C269 B.n224 VSUBS 0.006576f
C270 B.n225 VSUBS 0.006576f
C271 B.n226 VSUBS 0.006576f
C272 B.n227 VSUBS 0.006576f
C273 B.n228 VSUBS 0.006576f
C274 B.n229 VSUBS 0.006576f
C275 B.n230 VSUBS 0.01594f
C276 B.n231 VSUBS 0.01594f
C277 B.n232 VSUBS 0.016552f
C278 B.n233 VSUBS 0.006576f
C279 B.n234 VSUBS 0.006576f
C280 B.n235 VSUBS 0.006576f
C281 B.n236 VSUBS 0.006576f
C282 B.n237 VSUBS 0.006576f
C283 B.n238 VSUBS 0.006576f
C284 B.n239 VSUBS 0.006576f
C285 B.n240 VSUBS 0.006576f
C286 B.n241 VSUBS 0.006576f
C287 B.n242 VSUBS 0.006576f
C288 B.n243 VSUBS 0.006576f
C289 B.n244 VSUBS 0.006576f
C290 B.n245 VSUBS 0.006576f
C291 B.n246 VSUBS 0.006576f
C292 B.n247 VSUBS 0.006576f
C293 B.n248 VSUBS 0.006576f
C294 B.n249 VSUBS 0.006576f
C295 B.n250 VSUBS 0.006576f
C296 B.n251 VSUBS 0.006576f
C297 B.n252 VSUBS 0.006576f
C298 B.n253 VSUBS 0.006576f
C299 B.n254 VSUBS 0.006576f
C300 B.n255 VSUBS 0.006576f
C301 B.n256 VSUBS 0.006576f
C302 B.n257 VSUBS 0.006576f
C303 B.n258 VSUBS 0.006576f
C304 B.n259 VSUBS 0.006576f
C305 B.n260 VSUBS 0.006576f
C306 B.n261 VSUBS 0.006576f
C307 B.n262 VSUBS 0.006576f
C308 B.n263 VSUBS 0.006576f
C309 B.n264 VSUBS 0.006576f
C310 B.n265 VSUBS 0.006576f
C311 B.n266 VSUBS 0.006576f
C312 B.n267 VSUBS 0.006576f
C313 B.n268 VSUBS 0.006576f
C314 B.n269 VSUBS 0.006576f
C315 B.n270 VSUBS 0.006576f
C316 B.n271 VSUBS 0.006576f
C317 B.n272 VSUBS 0.006576f
C318 B.n273 VSUBS 0.006576f
C319 B.n274 VSUBS 0.006576f
C320 B.n275 VSUBS 0.006576f
C321 B.n276 VSUBS 0.006576f
C322 B.n277 VSUBS 0.006576f
C323 B.n278 VSUBS 0.006576f
C324 B.n279 VSUBS 0.006576f
C325 B.n280 VSUBS 0.006576f
C326 B.n281 VSUBS 0.006576f
C327 B.n282 VSUBS 0.006576f
C328 B.n283 VSUBS 0.006576f
C329 B.n284 VSUBS 0.006576f
C330 B.n285 VSUBS 0.006576f
C331 B.n286 VSUBS 0.006576f
C332 B.n287 VSUBS 0.006576f
C333 B.n288 VSUBS 0.006576f
C334 B.n289 VSUBS 0.006576f
C335 B.n290 VSUBS 0.006576f
C336 B.n291 VSUBS 0.006576f
C337 B.n292 VSUBS 0.006576f
C338 B.n293 VSUBS 0.006576f
C339 B.n294 VSUBS 0.006576f
C340 B.n295 VSUBS 0.006576f
C341 B.n296 VSUBS 0.006576f
C342 B.n297 VSUBS 0.006576f
C343 B.n298 VSUBS 0.006576f
C344 B.n299 VSUBS 0.006576f
C345 B.n300 VSUBS 0.006576f
C346 B.n301 VSUBS 0.006576f
C347 B.n302 VSUBS 0.006576f
C348 B.n303 VSUBS 0.006576f
C349 B.n304 VSUBS 0.004545f
C350 B.n305 VSUBS 0.015235f
C351 B.n306 VSUBS 0.005319f
C352 B.n307 VSUBS 0.006576f
C353 B.n308 VSUBS 0.006576f
C354 B.n309 VSUBS 0.006576f
C355 B.n310 VSUBS 0.006576f
C356 B.n311 VSUBS 0.006576f
C357 B.n312 VSUBS 0.006576f
C358 B.n313 VSUBS 0.006576f
C359 B.n314 VSUBS 0.006576f
C360 B.n315 VSUBS 0.006576f
C361 B.n316 VSUBS 0.006576f
C362 B.n317 VSUBS 0.006576f
C363 B.n318 VSUBS 0.005319f
C364 B.n319 VSUBS 0.006576f
C365 B.n320 VSUBS 0.006576f
C366 B.n321 VSUBS 0.004545f
C367 B.n322 VSUBS 0.006576f
C368 B.n323 VSUBS 0.006576f
C369 B.n324 VSUBS 0.006576f
C370 B.n325 VSUBS 0.006576f
C371 B.n326 VSUBS 0.006576f
C372 B.n327 VSUBS 0.006576f
C373 B.n328 VSUBS 0.006576f
C374 B.n329 VSUBS 0.006576f
C375 B.n330 VSUBS 0.006576f
C376 B.n331 VSUBS 0.006576f
C377 B.n332 VSUBS 0.006576f
C378 B.n333 VSUBS 0.006576f
C379 B.n334 VSUBS 0.006576f
C380 B.n335 VSUBS 0.006576f
C381 B.n336 VSUBS 0.006576f
C382 B.n337 VSUBS 0.006576f
C383 B.n338 VSUBS 0.006576f
C384 B.n339 VSUBS 0.006576f
C385 B.n340 VSUBS 0.006576f
C386 B.n341 VSUBS 0.006576f
C387 B.n342 VSUBS 0.006576f
C388 B.n343 VSUBS 0.006576f
C389 B.n344 VSUBS 0.006576f
C390 B.n345 VSUBS 0.006576f
C391 B.n346 VSUBS 0.006576f
C392 B.n347 VSUBS 0.006576f
C393 B.n348 VSUBS 0.006576f
C394 B.n349 VSUBS 0.006576f
C395 B.n350 VSUBS 0.006576f
C396 B.n351 VSUBS 0.006576f
C397 B.n352 VSUBS 0.006576f
C398 B.n353 VSUBS 0.006576f
C399 B.n354 VSUBS 0.006576f
C400 B.n355 VSUBS 0.006576f
C401 B.n356 VSUBS 0.006576f
C402 B.n357 VSUBS 0.006576f
C403 B.n358 VSUBS 0.006576f
C404 B.n359 VSUBS 0.006576f
C405 B.n360 VSUBS 0.006576f
C406 B.n361 VSUBS 0.006576f
C407 B.n362 VSUBS 0.006576f
C408 B.n363 VSUBS 0.006576f
C409 B.n364 VSUBS 0.006576f
C410 B.n365 VSUBS 0.006576f
C411 B.n366 VSUBS 0.006576f
C412 B.n367 VSUBS 0.006576f
C413 B.n368 VSUBS 0.006576f
C414 B.n369 VSUBS 0.006576f
C415 B.n370 VSUBS 0.006576f
C416 B.n371 VSUBS 0.006576f
C417 B.n372 VSUBS 0.006576f
C418 B.n373 VSUBS 0.006576f
C419 B.n374 VSUBS 0.006576f
C420 B.n375 VSUBS 0.006576f
C421 B.n376 VSUBS 0.006576f
C422 B.n377 VSUBS 0.006576f
C423 B.n378 VSUBS 0.006576f
C424 B.n379 VSUBS 0.006576f
C425 B.n380 VSUBS 0.006576f
C426 B.n381 VSUBS 0.006576f
C427 B.n382 VSUBS 0.006576f
C428 B.n383 VSUBS 0.006576f
C429 B.n384 VSUBS 0.006576f
C430 B.n385 VSUBS 0.006576f
C431 B.n386 VSUBS 0.006576f
C432 B.n387 VSUBS 0.006576f
C433 B.n388 VSUBS 0.006576f
C434 B.n389 VSUBS 0.006576f
C435 B.n390 VSUBS 0.006576f
C436 B.n391 VSUBS 0.006576f
C437 B.n392 VSUBS 0.016552f
C438 B.n393 VSUBS 0.016552f
C439 B.n394 VSUBS 0.01594f
C440 B.n395 VSUBS 0.006576f
C441 B.n396 VSUBS 0.006576f
C442 B.n397 VSUBS 0.006576f
C443 B.n398 VSUBS 0.006576f
C444 B.n399 VSUBS 0.006576f
C445 B.n400 VSUBS 0.006576f
C446 B.n401 VSUBS 0.006576f
C447 B.n402 VSUBS 0.006576f
C448 B.n403 VSUBS 0.006576f
C449 B.n404 VSUBS 0.006576f
C450 B.n405 VSUBS 0.006576f
C451 B.n406 VSUBS 0.006576f
C452 B.n407 VSUBS 0.006576f
C453 B.n408 VSUBS 0.006576f
C454 B.n409 VSUBS 0.006576f
C455 B.n410 VSUBS 0.006576f
C456 B.n411 VSUBS 0.006576f
C457 B.n412 VSUBS 0.006576f
C458 B.n413 VSUBS 0.006576f
C459 B.n414 VSUBS 0.006576f
C460 B.n415 VSUBS 0.006576f
C461 B.n416 VSUBS 0.006576f
C462 B.n417 VSUBS 0.006576f
C463 B.n418 VSUBS 0.006576f
C464 B.n419 VSUBS 0.006576f
C465 B.n420 VSUBS 0.006576f
C466 B.n421 VSUBS 0.006576f
C467 B.n422 VSUBS 0.006576f
C468 B.n423 VSUBS 0.006576f
C469 B.n424 VSUBS 0.006576f
C470 B.n425 VSUBS 0.006576f
C471 B.n426 VSUBS 0.006576f
C472 B.n427 VSUBS 0.006576f
C473 B.n428 VSUBS 0.006576f
C474 B.n429 VSUBS 0.006576f
C475 B.n430 VSUBS 0.006576f
C476 B.n431 VSUBS 0.006576f
C477 B.n432 VSUBS 0.006576f
C478 B.n433 VSUBS 0.006576f
C479 B.n434 VSUBS 0.006576f
C480 B.n435 VSUBS 0.006576f
C481 B.n436 VSUBS 0.006576f
C482 B.n437 VSUBS 0.006576f
C483 B.n438 VSUBS 0.006576f
C484 B.n439 VSUBS 0.006576f
C485 B.n440 VSUBS 0.006576f
C486 B.n441 VSUBS 0.006576f
C487 B.n442 VSUBS 0.006576f
C488 B.n443 VSUBS 0.006576f
C489 B.n444 VSUBS 0.006576f
C490 B.n445 VSUBS 0.006576f
C491 B.n446 VSUBS 0.006576f
C492 B.n447 VSUBS 0.006576f
C493 B.n448 VSUBS 0.006576f
C494 B.n449 VSUBS 0.006576f
C495 B.n450 VSUBS 0.006576f
C496 B.n451 VSUBS 0.006576f
C497 B.n452 VSUBS 0.006576f
C498 B.n453 VSUBS 0.006576f
C499 B.n454 VSUBS 0.006576f
C500 B.n455 VSUBS 0.006576f
C501 B.n456 VSUBS 0.006576f
C502 B.n457 VSUBS 0.006576f
C503 B.n458 VSUBS 0.006576f
C504 B.n459 VSUBS 0.006576f
C505 B.n460 VSUBS 0.006576f
C506 B.n461 VSUBS 0.006576f
C507 B.n462 VSUBS 0.006576f
C508 B.n463 VSUBS 0.006576f
C509 B.n464 VSUBS 0.006576f
C510 B.n465 VSUBS 0.006576f
C511 B.n466 VSUBS 0.006576f
C512 B.n467 VSUBS 0.006576f
C513 B.n468 VSUBS 0.006576f
C514 B.n469 VSUBS 0.006576f
C515 B.n470 VSUBS 0.006576f
C516 B.n471 VSUBS 0.006576f
C517 B.n472 VSUBS 0.006576f
C518 B.n473 VSUBS 0.006576f
C519 B.n474 VSUBS 0.006576f
C520 B.n475 VSUBS 0.006576f
C521 B.n476 VSUBS 0.006576f
C522 B.n477 VSUBS 0.006576f
C523 B.n478 VSUBS 0.006576f
C524 B.n479 VSUBS 0.006576f
C525 B.n480 VSUBS 0.006576f
C526 B.n481 VSUBS 0.006576f
C527 B.n482 VSUBS 0.006576f
C528 B.n483 VSUBS 0.006576f
C529 B.n484 VSUBS 0.006576f
C530 B.n485 VSUBS 0.006576f
C531 B.n486 VSUBS 0.006576f
C532 B.n487 VSUBS 0.006576f
C533 B.n488 VSUBS 0.006576f
C534 B.n489 VSUBS 0.006576f
C535 B.n490 VSUBS 0.006576f
C536 B.n491 VSUBS 0.006576f
C537 B.n492 VSUBS 0.006576f
C538 B.n493 VSUBS 0.01594f
C539 B.n494 VSUBS 0.016552f
C540 B.n495 VSUBS 0.015836f
C541 B.n496 VSUBS 0.006576f
C542 B.n497 VSUBS 0.006576f
C543 B.n498 VSUBS 0.006576f
C544 B.n499 VSUBS 0.006576f
C545 B.n500 VSUBS 0.006576f
C546 B.n501 VSUBS 0.006576f
C547 B.n502 VSUBS 0.006576f
C548 B.n503 VSUBS 0.006576f
C549 B.n504 VSUBS 0.006576f
C550 B.n505 VSUBS 0.006576f
C551 B.n506 VSUBS 0.006576f
C552 B.n507 VSUBS 0.006576f
C553 B.n508 VSUBS 0.006576f
C554 B.n509 VSUBS 0.006576f
C555 B.n510 VSUBS 0.006576f
C556 B.n511 VSUBS 0.006576f
C557 B.n512 VSUBS 0.006576f
C558 B.n513 VSUBS 0.006576f
C559 B.n514 VSUBS 0.006576f
C560 B.n515 VSUBS 0.006576f
C561 B.n516 VSUBS 0.006576f
C562 B.n517 VSUBS 0.006576f
C563 B.n518 VSUBS 0.006576f
C564 B.n519 VSUBS 0.006576f
C565 B.n520 VSUBS 0.006576f
C566 B.n521 VSUBS 0.006576f
C567 B.n522 VSUBS 0.006576f
C568 B.n523 VSUBS 0.006576f
C569 B.n524 VSUBS 0.006576f
C570 B.n525 VSUBS 0.006576f
C571 B.n526 VSUBS 0.006576f
C572 B.n527 VSUBS 0.006576f
C573 B.n528 VSUBS 0.006576f
C574 B.n529 VSUBS 0.006576f
C575 B.n530 VSUBS 0.006576f
C576 B.n531 VSUBS 0.006576f
C577 B.n532 VSUBS 0.006576f
C578 B.n533 VSUBS 0.006576f
C579 B.n534 VSUBS 0.006576f
C580 B.n535 VSUBS 0.006576f
C581 B.n536 VSUBS 0.006576f
C582 B.n537 VSUBS 0.006576f
C583 B.n538 VSUBS 0.006576f
C584 B.n539 VSUBS 0.006576f
C585 B.n540 VSUBS 0.006576f
C586 B.n541 VSUBS 0.006576f
C587 B.n542 VSUBS 0.006576f
C588 B.n543 VSUBS 0.006576f
C589 B.n544 VSUBS 0.006576f
C590 B.n545 VSUBS 0.006576f
C591 B.n546 VSUBS 0.006576f
C592 B.n547 VSUBS 0.006576f
C593 B.n548 VSUBS 0.006576f
C594 B.n549 VSUBS 0.006576f
C595 B.n550 VSUBS 0.006576f
C596 B.n551 VSUBS 0.006576f
C597 B.n552 VSUBS 0.006576f
C598 B.n553 VSUBS 0.006576f
C599 B.n554 VSUBS 0.006576f
C600 B.n555 VSUBS 0.006576f
C601 B.n556 VSUBS 0.006576f
C602 B.n557 VSUBS 0.006576f
C603 B.n558 VSUBS 0.006576f
C604 B.n559 VSUBS 0.006576f
C605 B.n560 VSUBS 0.006576f
C606 B.n561 VSUBS 0.006576f
C607 B.n562 VSUBS 0.006576f
C608 B.n563 VSUBS 0.006576f
C609 B.n564 VSUBS 0.006576f
C610 B.n565 VSUBS 0.006576f
C611 B.n566 VSUBS 0.006576f
C612 B.n567 VSUBS 0.004545f
C613 B.n568 VSUBS 0.015235f
C614 B.n569 VSUBS 0.005319f
C615 B.n570 VSUBS 0.006576f
C616 B.n571 VSUBS 0.006576f
C617 B.n572 VSUBS 0.006576f
C618 B.n573 VSUBS 0.006576f
C619 B.n574 VSUBS 0.006576f
C620 B.n575 VSUBS 0.006576f
C621 B.n576 VSUBS 0.006576f
C622 B.n577 VSUBS 0.006576f
C623 B.n578 VSUBS 0.006576f
C624 B.n579 VSUBS 0.006576f
C625 B.n580 VSUBS 0.006576f
C626 B.n581 VSUBS 0.005319f
C627 B.n582 VSUBS 0.015235f
C628 B.n583 VSUBS 0.004545f
C629 B.n584 VSUBS 0.006576f
C630 B.n585 VSUBS 0.006576f
C631 B.n586 VSUBS 0.006576f
C632 B.n587 VSUBS 0.006576f
C633 B.n588 VSUBS 0.006576f
C634 B.n589 VSUBS 0.006576f
C635 B.n590 VSUBS 0.006576f
C636 B.n591 VSUBS 0.006576f
C637 B.n592 VSUBS 0.006576f
C638 B.n593 VSUBS 0.006576f
C639 B.n594 VSUBS 0.006576f
C640 B.n595 VSUBS 0.006576f
C641 B.n596 VSUBS 0.006576f
C642 B.n597 VSUBS 0.006576f
C643 B.n598 VSUBS 0.006576f
C644 B.n599 VSUBS 0.006576f
C645 B.n600 VSUBS 0.006576f
C646 B.n601 VSUBS 0.006576f
C647 B.n602 VSUBS 0.006576f
C648 B.n603 VSUBS 0.006576f
C649 B.n604 VSUBS 0.006576f
C650 B.n605 VSUBS 0.006576f
C651 B.n606 VSUBS 0.006576f
C652 B.n607 VSUBS 0.006576f
C653 B.n608 VSUBS 0.006576f
C654 B.n609 VSUBS 0.006576f
C655 B.n610 VSUBS 0.006576f
C656 B.n611 VSUBS 0.006576f
C657 B.n612 VSUBS 0.006576f
C658 B.n613 VSUBS 0.006576f
C659 B.n614 VSUBS 0.006576f
C660 B.n615 VSUBS 0.006576f
C661 B.n616 VSUBS 0.006576f
C662 B.n617 VSUBS 0.006576f
C663 B.n618 VSUBS 0.006576f
C664 B.n619 VSUBS 0.006576f
C665 B.n620 VSUBS 0.006576f
C666 B.n621 VSUBS 0.006576f
C667 B.n622 VSUBS 0.006576f
C668 B.n623 VSUBS 0.006576f
C669 B.n624 VSUBS 0.006576f
C670 B.n625 VSUBS 0.006576f
C671 B.n626 VSUBS 0.006576f
C672 B.n627 VSUBS 0.006576f
C673 B.n628 VSUBS 0.006576f
C674 B.n629 VSUBS 0.006576f
C675 B.n630 VSUBS 0.006576f
C676 B.n631 VSUBS 0.006576f
C677 B.n632 VSUBS 0.006576f
C678 B.n633 VSUBS 0.006576f
C679 B.n634 VSUBS 0.006576f
C680 B.n635 VSUBS 0.006576f
C681 B.n636 VSUBS 0.006576f
C682 B.n637 VSUBS 0.006576f
C683 B.n638 VSUBS 0.006576f
C684 B.n639 VSUBS 0.006576f
C685 B.n640 VSUBS 0.006576f
C686 B.n641 VSUBS 0.006576f
C687 B.n642 VSUBS 0.006576f
C688 B.n643 VSUBS 0.006576f
C689 B.n644 VSUBS 0.006576f
C690 B.n645 VSUBS 0.006576f
C691 B.n646 VSUBS 0.006576f
C692 B.n647 VSUBS 0.006576f
C693 B.n648 VSUBS 0.006576f
C694 B.n649 VSUBS 0.006576f
C695 B.n650 VSUBS 0.006576f
C696 B.n651 VSUBS 0.006576f
C697 B.n652 VSUBS 0.006576f
C698 B.n653 VSUBS 0.006576f
C699 B.n654 VSUBS 0.006576f
C700 B.n655 VSUBS 0.016552f
C701 B.n656 VSUBS 0.016552f
C702 B.n657 VSUBS 0.01594f
C703 B.n658 VSUBS 0.006576f
C704 B.n659 VSUBS 0.006576f
C705 B.n660 VSUBS 0.006576f
C706 B.n661 VSUBS 0.006576f
C707 B.n662 VSUBS 0.006576f
C708 B.n663 VSUBS 0.006576f
C709 B.n664 VSUBS 0.006576f
C710 B.n665 VSUBS 0.006576f
C711 B.n666 VSUBS 0.006576f
C712 B.n667 VSUBS 0.006576f
C713 B.n668 VSUBS 0.006576f
C714 B.n669 VSUBS 0.006576f
C715 B.n670 VSUBS 0.006576f
C716 B.n671 VSUBS 0.006576f
C717 B.n672 VSUBS 0.006576f
C718 B.n673 VSUBS 0.006576f
C719 B.n674 VSUBS 0.006576f
C720 B.n675 VSUBS 0.006576f
C721 B.n676 VSUBS 0.006576f
C722 B.n677 VSUBS 0.006576f
C723 B.n678 VSUBS 0.006576f
C724 B.n679 VSUBS 0.006576f
C725 B.n680 VSUBS 0.006576f
C726 B.n681 VSUBS 0.006576f
C727 B.n682 VSUBS 0.006576f
C728 B.n683 VSUBS 0.006576f
C729 B.n684 VSUBS 0.006576f
C730 B.n685 VSUBS 0.006576f
C731 B.n686 VSUBS 0.006576f
C732 B.n687 VSUBS 0.006576f
C733 B.n688 VSUBS 0.006576f
C734 B.n689 VSUBS 0.006576f
C735 B.n690 VSUBS 0.006576f
C736 B.n691 VSUBS 0.006576f
C737 B.n692 VSUBS 0.006576f
C738 B.n693 VSUBS 0.006576f
C739 B.n694 VSUBS 0.006576f
C740 B.n695 VSUBS 0.006576f
C741 B.n696 VSUBS 0.006576f
C742 B.n697 VSUBS 0.006576f
C743 B.n698 VSUBS 0.006576f
C744 B.n699 VSUBS 0.006576f
C745 B.n700 VSUBS 0.006576f
C746 B.n701 VSUBS 0.006576f
C747 B.n702 VSUBS 0.006576f
C748 B.n703 VSUBS 0.006576f
C749 B.n704 VSUBS 0.006576f
C750 B.n705 VSUBS 0.006576f
C751 B.n706 VSUBS 0.006576f
C752 B.n707 VSUBS 0.01489f
C753 VDD1.t1 VSUBS 3.56861f
C754 VDD1.t0 VSUBS 4.6172f
C755 VTAIL.t3 VSUBS 3.38975f
C756 VTAIL.n0 VSUBS 3.20296f
C757 VTAIL.t1 VSUBS 3.38977f
C758 VTAIL.n1 VSUBS 3.28457f
C759 VTAIL.t2 VSUBS 3.38975f
C760 VTAIL.n2 VSUBS 2.93591f
C761 VTAIL.t0 VSUBS 3.38975f
C762 VTAIL.n3 VSUBS 2.79849f
C763 VP.t0 VSUBS 6.33392f
C764 VP.t1 VSUBS 5.36362f
C765 VP.n0 VSUBS 5.66573f
.ends

