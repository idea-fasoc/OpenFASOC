* NGSPICE file created from diff_pair_sample_1070.ext - technology: sky130A

.subckt diff_pair_sample_1070 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7144 pd=14.7 as=2.7144 ps=14.7 w=6.96 l=0.5
X1 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=2.7144 pd=14.7 as=0 ps=0 w=6.96 l=0.5
X2 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=2.7144 pd=14.7 as=0 ps=0 w=6.96 l=0.5
X3 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7144 pd=14.7 as=2.7144 ps=14.7 w=6.96 l=0.5
X4 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7144 pd=14.7 as=2.7144 ps=14.7 w=6.96 l=0.5
X5 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7144 pd=14.7 as=0 ps=0 w=6.96 l=0.5
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7144 pd=14.7 as=0 ps=0 w=6.96 l=0.5
X7 VDD2.t0 VN.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7144 pd=14.7 as=2.7144 ps=14.7 w=6.96 l=0.5
R0 VN VN.t0 611.004
R1 VN VN.t1 575.389
R2 VTAIL.n1 VTAIL.t3 49.45
R3 VTAIL.n3 VTAIL.t2 49.4498
R4 VTAIL.n0 VTAIL.t0 49.4498
R5 VTAIL.n2 VTAIL.t1 49.4498
R6 VTAIL.n1 VTAIL.n0 19.8152
R7 VTAIL.n3 VTAIL.n2 19.0996
R8 VTAIL.n2 VTAIL.n1 0.828086
R9 VTAIL VTAIL.n0 0.707397
R10 VTAIL VTAIL.n3 0.12119
R11 VDD2.n0 VDD2.t0 97.2363
R12 VDD2.n0 VDD2.t1 66.1286
R13 VDD2 VDD2.n0 0.237569
R14 B.n433 B.n432 585
R15 B.n434 B.n433 585
R16 B.n188 B.n59 585
R17 B.n187 B.n186 585
R18 B.n185 B.n184 585
R19 B.n183 B.n182 585
R20 B.n181 B.n180 585
R21 B.n179 B.n178 585
R22 B.n177 B.n176 585
R23 B.n175 B.n174 585
R24 B.n173 B.n172 585
R25 B.n171 B.n170 585
R26 B.n169 B.n168 585
R27 B.n167 B.n166 585
R28 B.n165 B.n164 585
R29 B.n163 B.n162 585
R30 B.n161 B.n160 585
R31 B.n159 B.n158 585
R32 B.n157 B.n156 585
R33 B.n155 B.n154 585
R34 B.n153 B.n152 585
R35 B.n151 B.n150 585
R36 B.n149 B.n148 585
R37 B.n147 B.n146 585
R38 B.n145 B.n144 585
R39 B.n143 B.n142 585
R40 B.n141 B.n140 585
R41 B.n139 B.n138 585
R42 B.n137 B.n136 585
R43 B.n135 B.n134 585
R44 B.n133 B.n132 585
R45 B.n131 B.n130 585
R46 B.n129 B.n128 585
R47 B.n127 B.n126 585
R48 B.n125 B.n124 585
R49 B.n123 B.n122 585
R50 B.n121 B.n120 585
R51 B.n118 B.n117 585
R52 B.n116 B.n115 585
R53 B.n114 B.n113 585
R54 B.n112 B.n111 585
R55 B.n110 B.n109 585
R56 B.n108 B.n107 585
R57 B.n106 B.n105 585
R58 B.n104 B.n103 585
R59 B.n102 B.n101 585
R60 B.n100 B.n99 585
R61 B.n98 B.n97 585
R62 B.n96 B.n95 585
R63 B.n94 B.n93 585
R64 B.n92 B.n91 585
R65 B.n90 B.n89 585
R66 B.n88 B.n87 585
R67 B.n86 B.n85 585
R68 B.n84 B.n83 585
R69 B.n82 B.n81 585
R70 B.n80 B.n79 585
R71 B.n78 B.n77 585
R72 B.n76 B.n75 585
R73 B.n74 B.n73 585
R74 B.n72 B.n71 585
R75 B.n70 B.n69 585
R76 B.n68 B.n67 585
R77 B.n66 B.n65 585
R78 B.n431 B.n27 585
R79 B.n435 B.n27 585
R80 B.n430 B.n26 585
R81 B.n436 B.n26 585
R82 B.n429 B.n428 585
R83 B.n428 B.n22 585
R84 B.n427 B.n21 585
R85 B.n442 B.n21 585
R86 B.n426 B.n20 585
R87 B.n443 B.n20 585
R88 B.n425 B.n19 585
R89 B.n444 B.n19 585
R90 B.n424 B.n423 585
R91 B.n423 B.n15 585
R92 B.n422 B.n14 585
R93 B.n450 B.n14 585
R94 B.n421 B.n13 585
R95 B.n451 B.n13 585
R96 B.n420 B.n12 585
R97 B.n452 B.n12 585
R98 B.n419 B.n418 585
R99 B.n418 B.n11 585
R100 B.n417 B.n7 585
R101 B.n458 B.n7 585
R102 B.n416 B.n6 585
R103 B.n459 B.n6 585
R104 B.n415 B.n5 585
R105 B.n460 B.n5 585
R106 B.n414 B.n413 585
R107 B.n413 B.n4 585
R108 B.n412 B.n189 585
R109 B.n412 B.n411 585
R110 B.n401 B.n190 585
R111 B.n404 B.n190 585
R112 B.n403 B.n402 585
R113 B.n405 B.n403 585
R114 B.n400 B.n195 585
R115 B.n195 B.n194 585
R116 B.n399 B.n398 585
R117 B.n398 B.n397 585
R118 B.n197 B.n196 585
R119 B.n198 B.n197 585
R120 B.n390 B.n389 585
R121 B.n391 B.n390 585
R122 B.n388 B.n202 585
R123 B.n206 B.n202 585
R124 B.n387 B.n386 585
R125 B.n386 B.n385 585
R126 B.n204 B.n203 585
R127 B.n205 B.n204 585
R128 B.n378 B.n377 585
R129 B.n379 B.n378 585
R130 B.n376 B.n211 585
R131 B.n211 B.n210 585
R132 B.n370 B.n369 585
R133 B.n368 B.n244 585
R134 B.n367 B.n243 585
R135 B.n372 B.n243 585
R136 B.n366 B.n365 585
R137 B.n364 B.n363 585
R138 B.n362 B.n361 585
R139 B.n360 B.n359 585
R140 B.n358 B.n357 585
R141 B.n356 B.n355 585
R142 B.n354 B.n353 585
R143 B.n352 B.n351 585
R144 B.n350 B.n349 585
R145 B.n348 B.n347 585
R146 B.n346 B.n345 585
R147 B.n344 B.n343 585
R148 B.n342 B.n341 585
R149 B.n340 B.n339 585
R150 B.n338 B.n337 585
R151 B.n336 B.n335 585
R152 B.n334 B.n333 585
R153 B.n332 B.n331 585
R154 B.n330 B.n329 585
R155 B.n328 B.n327 585
R156 B.n326 B.n325 585
R157 B.n324 B.n323 585
R158 B.n322 B.n321 585
R159 B.n320 B.n319 585
R160 B.n318 B.n317 585
R161 B.n316 B.n315 585
R162 B.n314 B.n313 585
R163 B.n312 B.n311 585
R164 B.n310 B.n309 585
R165 B.n308 B.n307 585
R166 B.n306 B.n305 585
R167 B.n304 B.n303 585
R168 B.n302 B.n301 585
R169 B.n299 B.n298 585
R170 B.n297 B.n296 585
R171 B.n295 B.n294 585
R172 B.n293 B.n292 585
R173 B.n291 B.n290 585
R174 B.n289 B.n288 585
R175 B.n287 B.n286 585
R176 B.n285 B.n284 585
R177 B.n283 B.n282 585
R178 B.n281 B.n280 585
R179 B.n279 B.n278 585
R180 B.n277 B.n276 585
R181 B.n275 B.n274 585
R182 B.n273 B.n272 585
R183 B.n271 B.n270 585
R184 B.n269 B.n268 585
R185 B.n267 B.n266 585
R186 B.n265 B.n264 585
R187 B.n263 B.n262 585
R188 B.n261 B.n260 585
R189 B.n259 B.n258 585
R190 B.n257 B.n256 585
R191 B.n255 B.n254 585
R192 B.n253 B.n252 585
R193 B.n251 B.n250 585
R194 B.n213 B.n212 585
R195 B.n375 B.n374 585
R196 B.n209 B.n208 585
R197 B.n210 B.n209 585
R198 B.n381 B.n380 585
R199 B.n380 B.n379 585
R200 B.n382 B.n207 585
R201 B.n207 B.n205 585
R202 B.n384 B.n383 585
R203 B.n385 B.n384 585
R204 B.n201 B.n200 585
R205 B.n206 B.n201 585
R206 B.n393 B.n392 585
R207 B.n392 B.n391 585
R208 B.n394 B.n199 585
R209 B.n199 B.n198 585
R210 B.n396 B.n395 585
R211 B.n397 B.n396 585
R212 B.n193 B.n192 585
R213 B.n194 B.n193 585
R214 B.n407 B.n406 585
R215 B.n406 B.n405 585
R216 B.n408 B.n191 585
R217 B.n404 B.n191 585
R218 B.n410 B.n409 585
R219 B.n411 B.n410 585
R220 B.n2 B.n0 585
R221 B.n4 B.n2 585
R222 B.n3 B.n1 585
R223 B.n459 B.n3 585
R224 B.n457 B.n456 585
R225 B.n458 B.n457 585
R226 B.n455 B.n8 585
R227 B.n11 B.n8 585
R228 B.n454 B.n453 585
R229 B.n453 B.n452 585
R230 B.n10 B.n9 585
R231 B.n451 B.n10 585
R232 B.n449 B.n448 585
R233 B.n450 B.n449 585
R234 B.n447 B.n16 585
R235 B.n16 B.n15 585
R236 B.n446 B.n445 585
R237 B.n445 B.n444 585
R238 B.n18 B.n17 585
R239 B.n443 B.n18 585
R240 B.n441 B.n440 585
R241 B.n442 B.n441 585
R242 B.n439 B.n23 585
R243 B.n23 B.n22 585
R244 B.n438 B.n437 585
R245 B.n437 B.n436 585
R246 B.n25 B.n24 585
R247 B.n435 B.n25 585
R248 B.n462 B.n461 585
R249 B.n461 B.n460 585
R250 B.n248 B.t9 541.88
R251 B.n245 B.t13 541.88
R252 B.n63 B.t6 541.88
R253 B.n60 B.t2 541.88
R254 B.n370 B.n209 521.33
R255 B.n65 B.n25 521.33
R256 B.n374 B.n211 521.33
R257 B.n433 B.n27 521.33
R258 B.n434 B.n58 256.663
R259 B.n434 B.n57 256.663
R260 B.n434 B.n56 256.663
R261 B.n434 B.n55 256.663
R262 B.n434 B.n54 256.663
R263 B.n434 B.n53 256.663
R264 B.n434 B.n52 256.663
R265 B.n434 B.n51 256.663
R266 B.n434 B.n50 256.663
R267 B.n434 B.n49 256.663
R268 B.n434 B.n48 256.663
R269 B.n434 B.n47 256.663
R270 B.n434 B.n46 256.663
R271 B.n434 B.n45 256.663
R272 B.n434 B.n44 256.663
R273 B.n434 B.n43 256.663
R274 B.n434 B.n42 256.663
R275 B.n434 B.n41 256.663
R276 B.n434 B.n40 256.663
R277 B.n434 B.n39 256.663
R278 B.n434 B.n38 256.663
R279 B.n434 B.n37 256.663
R280 B.n434 B.n36 256.663
R281 B.n434 B.n35 256.663
R282 B.n434 B.n34 256.663
R283 B.n434 B.n33 256.663
R284 B.n434 B.n32 256.663
R285 B.n434 B.n31 256.663
R286 B.n434 B.n30 256.663
R287 B.n434 B.n29 256.663
R288 B.n434 B.n28 256.663
R289 B.n372 B.n371 256.663
R290 B.n372 B.n214 256.663
R291 B.n372 B.n215 256.663
R292 B.n372 B.n216 256.663
R293 B.n372 B.n217 256.663
R294 B.n372 B.n218 256.663
R295 B.n372 B.n219 256.663
R296 B.n372 B.n220 256.663
R297 B.n372 B.n221 256.663
R298 B.n372 B.n222 256.663
R299 B.n372 B.n223 256.663
R300 B.n372 B.n224 256.663
R301 B.n372 B.n225 256.663
R302 B.n372 B.n226 256.663
R303 B.n372 B.n227 256.663
R304 B.n372 B.n228 256.663
R305 B.n372 B.n229 256.663
R306 B.n372 B.n230 256.663
R307 B.n372 B.n231 256.663
R308 B.n372 B.n232 256.663
R309 B.n372 B.n233 256.663
R310 B.n372 B.n234 256.663
R311 B.n372 B.n235 256.663
R312 B.n372 B.n236 256.663
R313 B.n372 B.n237 256.663
R314 B.n372 B.n238 256.663
R315 B.n372 B.n239 256.663
R316 B.n372 B.n240 256.663
R317 B.n372 B.n241 256.663
R318 B.n372 B.n242 256.663
R319 B.n373 B.n372 256.663
R320 B.n380 B.n209 163.367
R321 B.n380 B.n207 163.367
R322 B.n384 B.n207 163.367
R323 B.n384 B.n201 163.367
R324 B.n392 B.n201 163.367
R325 B.n392 B.n199 163.367
R326 B.n396 B.n199 163.367
R327 B.n396 B.n193 163.367
R328 B.n406 B.n193 163.367
R329 B.n406 B.n191 163.367
R330 B.n410 B.n191 163.367
R331 B.n410 B.n2 163.367
R332 B.n461 B.n2 163.367
R333 B.n461 B.n3 163.367
R334 B.n457 B.n3 163.367
R335 B.n457 B.n8 163.367
R336 B.n453 B.n8 163.367
R337 B.n453 B.n10 163.367
R338 B.n449 B.n10 163.367
R339 B.n449 B.n16 163.367
R340 B.n445 B.n16 163.367
R341 B.n445 B.n18 163.367
R342 B.n441 B.n18 163.367
R343 B.n441 B.n23 163.367
R344 B.n437 B.n23 163.367
R345 B.n437 B.n25 163.367
R346 B.n244 B.n243 163.367
R347 B.n365 B.n243 163.367
R348 B.n363 B.n362 163.367
R349 B.n359 B.n358 163.367
R350 B.n355 B.n354 163.367
R351 B.n351 B.n350 163.367
R352 B.n347 B.n346 163.367
R353 B.n343 B.n342 163.367
R354 B.n339 B.n338 163.367
R355 B.n335 B.n334 163.367
R356 B.n331 B.n330 163.367
R357 B.n327 B.n326 163.367
R358 B.n323 B.n322 163.367
R359 B.n319 B.n318 163.367
R360 B.n315 B.n314 163.367
R361 B.n311 B.n310 163.367
R362 B.n307 B.n306 163.367
R363 B.n303 B.n302 163.367
R364 B.n298 B.n297 163.367
R365 B.n294 B.n293 163.367
R366 B.n290 B.n289 163.367
R367 B.n286 B.n285 163.367
R368 B.n282 B.n281 163.367
R369 B.n278 B.n277 163.367
R370 B.n274 B.n273 163.367
R371 B.n270 B.n269 163.367
R372 B.n266 B.n265 163.367
R373 B.n262 B.n261 163.367
R374 B.n258 B.n257 163.367
R375 B.n254 B.n253 163.367
R376 B.n250 B.n213 163.367
R377 B.n378 B.n211 163.367
R378 B.n378 B.n204 163.367
R379 B.n386 B.n204 163.367
R380 B.n386 B.n202 163.367
R381 B.n390 B.n202 163.367
R382 B.n390 B.n197 163.367
R383 B.n398 B.n197 163.367
R384 B.n398 B.n195 163.367
R385 B.n403 B.n195 163.367
R386 B.n403 B.n190 163.367
R387 B.n412 B.n190 163.367
R388 B.n413 B.n412 163.367
R389 B.n413 B.n5 163.367
R390 B.n6 B.n5 163.367
R391 B.n7 B.n6 163.367
R392 B.n418 B.n7 163.367
R393 B.n418 B.n12 163.367
R394 B.n13 B.n12 163.367
R395 B.n14 B.n13 163.367
R396 B.n423 B.n14 163.367
R397 B.n423 B.n19 163.367
R398 B.n20 B.n19 163.367
R399 B.n21 B.n20 163.367
R400 B.n428 B.n21 163.367
R401 B.n428 B.n26 163.367
R402 B.n27 B.n26 163.367
R403 B.n69 B.n68 163.367
R404 B.n73 B.n72 163.367
R405 B.n77 B.n76 163.367
R406 B.n81 B.n80 163.367
R407 B.n85 B.n84 163.367
R408 B.n89 B.n88 163.367
R409 B.n93 B.n92 163.367
R410 B.n97 B.n96 163.367
R411 B.n101 B.n100 163.367
R412 B.n105 B.n104 163.367
R413 B.n109 B.n108 163.367
R414 B.n113 B.n112 163.367
R415 B.n117 B.n116 163.367
R416 B.n122 B.n121 163.367
R417 B.n126 B.n125 163.367
R418 B.n130 B.n129 163.367
R419 B.n134 B.n133 163.367
R420 B.n138 B.n137 163.367
R421 B.n142 B.n141 163.367
R422 B.n146 B.n145 163.367
R423 B.n150 B.n149 163.367
R424 B.n154 B.n153 163.367
R425 B.n158 B.n157 163.367
R426 B.n162 B.n161 163.367
R427 B.n166 B.n165 163.367
R428 B.n170 B.n169 163.367
R429 B.n174 B.n173 163.367
R430 B.n178 B.n177 163.367
R431 B.n182 B.n181 163.367
R432 B.n186 B.n185 163.367
R433 B.n433 B.n59 163.367
R434 B.n372 B.n210 110.404
R435 B.n435 B.n434 110.404
R436 B.n248 B.t12 88.1813
R437 B.n60 B.t4 88.1813
R438 B.n245 B.t15 88.1735
R439 B.n63 B.t7 88.1735
R440 B.n249 B.t11 72.0843
R441 B.n61 B.t5 72.0843
R442 B.n246 B.t14 72.0765
R443 B.n64 B.t8 72.0765
R444 B.n371 B.n370 71.676
R445 B.n365 B.n214 71.676
R446 B.n362 B.n215 71.676
R447 B.n358 B.n216 71.676
R448 B.n354 B.n217 71.676
R449 B.n350 B.n218 71.676
R450 B.n346 B.n219 71.676
R451 B.n342 B.n220 71.676
R452 B.n338 B.n221 71.676
R453 B.n334 B.n222 71.676
R454 B.n330 B.n223 71.676
R455 B.n326 B.n224 71.676
R456 B.n322 B.n225 71.676
R457 B.n318 B.n226 71.676
R458 B.n314 B.n227 71.676
R459 B.n310 B.n228 71.676
R460 B.n306 B.n229 71.676
R461 B.n302 B.n230 71.676
R462 B.n297 B.n231 71.676
R463 B.n293 B.n232 71.676
R464 B.n289 B.n233 71.676
R465 B.n285 B.n234 71.676
R466 B.n281 B.n235 71.676
R467 B.n277 B.n236 71.676
R468 B.n273 B.n237 71.676
R469 B.n269 B.n238 71.676
R470 B.n265 B.n239 71.676
R471 B.n261 B.n240 71.676
R472 B.n257 B.n241 71.676
R473 B.n253 B.n242 71.676
R474 B.n373 B.n213 71.676
R475 B.n65 B.n28 71.676
R476 B.n69 B.n29 71.676
R477 B.n73 B.n30 71.676
R478 B.n77 B.n31 71.676
R479 B.n81 B.n32 71.676
R480 B.n85 B.n33 71.676
R481 B.n89 B.n34 71.676
R482 B.n93 B.n35 71.676
R483 B.n97 B.n36 71.676
R484 B.n101 B.n37 71.676
R485 B.n105 B.n38 71.676
R486 B.n109 B.n39 71.676
R487 B.n113 B.n40 71.676
R488 B.n117 B.n41 71.676
R489 B.n122 B.n42 71.676
R490 B.n126 B.n43 71.676
R491 B.n130 B.n44 71.676
R492 B.n134 B.n45 71.676
R493 B.n138 B.n46 71.676
R494 B.n142 B.n47 71.676
R495 B.n146 B.n48 71.676
R496 B.n150 B.n49 71.676
R497 B.n154 B.n50 71.676
R498 B.n158 B.n51 71.676
R499 B.n162 B.n52 71.676
R500 B.n166 B.n53 71.676
R501 B.n170 B.n54 71.676
R502 B.n174 B.n55 71.676
R503 B.n178 B.n56 71.676
R504 B.n182 B.n57 71.676
R505 B.n186 B.n58 71.676
R506 B.n59 B.n58 71.676
R507 B.n185 B.n57 71.676
R508 B.n181 B.n56 71.676
R509 B.n177 B.n55 71.676
R510 B.n173 B.n54 71.676
R511 B.n169 B.n53 71.676
R512 B.n165 B.n52 71.676
R513 B.n161 B.n51 71.676
R514 B.n157 B.n50 71.676
R515 B.n153 B.n49 71.676
R516 B.n149 B.n48 71.676
R517 B.n145 B.n47 71.676
R518 B.n141 B.n46 71.676
R519 B.n137 B.n45 71.676
R520 B.n133 B.n44 71.676
R521 B.n129 B.n43 71.676
R522 B.n125 B.n42 71.676
R523 B.n121 B.n41 71.676
R524 B.n116 B.n40 71.676
R525 B.n112 B.n39 71.676
R526 B.n108 B.n38 71.676
R527 B.n104 B.n37 71.676
R528 B.n100 B.n36 71.676
R529 B.n96 B.n35 71.676
R530 B.n92 B.n34 71.676
R531 B.n88 B.n33 71.676
R532 B.n84 B.n32 71.676
R533 B.n80 B.n31 71.676
R534 B.n76 B.n30 71.676
R535 B.n72 B.n29 71.676
R536 B.n68 B.n28 71.676
R537 B.n371 B.n244 71.676
R538 B.n363 B.n214 71.676
R539 B.n359 B.n215 71.676
R540 B.n355 B.n216 71.676
R541 B.n351 B.n217 71.676
R542 B.n347 B.n218 71.676
R543 B.n343 B.n219 71.676
R544 B.n339 B.n220 71.676
R545 B.n335 B.n221 71.676
R546 B.n331 B.n222 71.676
R547 B.n327 B.n223 71.676
R548 B.n323 B.n224 71.676
R549 B.n319 B.n225 71.676
R550 B.n315 B.n226 71.676
R551 B.n311 B.n227 71.676
R552 B.n307 B.n228 71.676
R553 B.n303 B.n229 71.676
R554 B.n298 B.n230 71.676
R555 B.n294 B.n231 71.676
R556 B.n290 B.n232 71.676
R557 B.n286 B.n233 71.676
R558 B.n282 B.n234 71.676
R559 B.n278 B.n235 71.676
R560 B.n274 B.n236 71.676
R561 B.n270 B.n237 71.676
R562 B.n266 B.n238 71.676
R563 B.n262 B.n239 71.676
R564 B.n258 B.n240 71.676
R565 B.n254 B.n241 71.676
R566 B.n250 B.n242 71.676
R567 B.n374 B.n373 71.676
R568 B.n379 B.n210 61.0368
R569 B.n379 B.n205 61.0368
R570 B.n385 B.n205 61.0368
R571 B.n385 B.n206 61.0368
R572 B.n391 B.n198 61.0368
R573 B.n397 B.n198 61.0368
R574 B.n397 B.n194 61.0368
R575 B.n405 B.n194 61.0368
R576 B.n405 B.n404 61.0368
R577 B.n411 B.n4 61.0368
R578 B.n460 B.n4 61.0368
R579 B.n460 B.n459 61.0368
R580 B.n459 B.n458 61.0368
R581 B.n452 B.n11 61.0368
R582 B.n452 B.n451 61.0368
R583 B.n451 B.n450 61.0368
R584 B.n450 B.n15 61.0368
R585 B.n444 B.n15 61.0368
R586 B.n443 B.n442 61.0368
R587 B.n442 B.n22 61.0368
R588 B.n436 B.n22 61.0368
R589 B.n436 B.n435 61.0368
R590 B.n300 B.n249 59.5399
R591 B.n247 B.n246 59.5399
R592 B.n119 B.n64 59.5399
R593 B.n62 B.n61 59.5399
R594 B.n411 B.t0 50.2657
R595 B.n458 B.t1 50.2657
R596 B.n66 B.n24 33.8737
R597 B.n432 B.n431 33.8737
R598 B.n376 B.n375 33.8737
R599 B.n369 B.n208 33.8737
R600 B.n206 B.t10 32.3138
R601 B.t3 B.n443 32.3138
R602 B.n391 B.t10 28.7235
R603 B.n444 B.t3 28.7235
R604 B B.n462 18.0485
R605 B.n249 B.n248 16.0975
R606 B.n246 B.n245 16.0975
R607 B.n64 B.n63 16.0975
R608 B.n61 B.n60 16.0975
R609 B.n404 B.t0 10.7716
R610 B.n11 B.t1 10.7716
R611 B.n67 B.n66 10.6151
R612 B.n70 B.n67 10.6151
R613 B.n71 B.n70 10.6151
R614 B.n74 B.n71 10.6151
R615 B.n75 B.n74 10.6151
R616 B.n78 B.n75 10.6151
R617 B.n79 B.n78 10.6151
R618 B.n82 B.n79 10.6151
R619 B.n83 B.n82 10.6151
R620 B.n86 B.n83 10.6151
R621 B.n87 B.n86 10.6151
R622 B.n90 B.n87 10.6151
R623 B.n91 B.n90 10.6151
R624 B.n94 B.n91 10.6151
R625 B.n95 B.n94 10.6151
R626 B.n98 B.n95 10.6151
R627 B.n99 B.n98 10.6151
R628 B.n102 B.n99 10.6151
R629 B.n103 B.n102 10.6151
R630 B.n106 B.n103 10.6151
R631 B.n107 B.n106 10.6151
R632 B.n110 B.n107 10.6151
R633 B.n111 B.n110 10.6151
R634 B.n114 B.n111 10.6151
R635 B.n115 B.n114 10.6151
R636 B.n118 B.n115 10.6151
R637 B.n123 B.n120 10.6151
R638 B.n124 B.n123 10.6151
R639 B.n127 B.n124 10.6151
R640 B.n128 B.n127 10.6151
R641 B.n131 B.n128 10.6151
R642 B.n132 B.n131 10.6151
R643 B.n135 B.n132 10.6151
R644 B.n136 B.n135 10.6151
R645 B.n140 B.n139 10.6151
R646 B.n143 B.n140 10.6151
R647 B.n144 B.n143 10.6151
R648 B.n147 B.n144 10.6151
R649 B.n148 B.n147 10.6151
R650 B.n151 B.n148 10.6151
R651 B.n152 B.n151 10.6151
R652 B.n155 B.n152 10.6151
R653 B.n156 B.n155 10.6151
R654 B.n159 B.n156 10.6151
R655 B.n160 B.n159 10.6151
R656 B.n163 B.n160 10.6151
R657 B.n164 B.n163 10.6151
R658 B.n167 B.n164 10.6151
R659 B.n168 B.n167 10.6151
R660 B.n171 B.n168 10.6151
R661 B.n172 B.n171 10.6151
R662 B.n175 B.n172 10.6151
R663 B.n176 B.n175 10.6151
R664 B.n179 B.n176 10.6151
R665 B.n180 B.n179 10.6151
R666 B.n183 B.n180 10.6151
R667 B.n184 B.n183 10.6151
R668 B.n187 B.n184 10.6151
R669 B.n188 B.n187 10.6151
R670 B.n432 B.n188 10.6151
R671 B.n377 B.n376 10.6151
R672 B.n377 B.n203 10.6151
R673 B.n387 B.n203 10.6151
R674 B.n388 B.n387 10.6151
R675 B.n389 B.n388 10.6151
R676 B.n389 B.n196 10.6151
R677 B.n399 B.n196 10.6151
R678 B.n400 B.n399 10.6151
R679 B.n402 B.n400 10.6151
R680 B.n402 B.n401 10.6151
R681 B.n401 B.n189 10.6151
R682 B.n414 B.n189 10.6151
R683 B.n415 B.n414 10.6151
R684 B.n416 B.n415 10.6151
R685 B.n417 B.n416 10.6151
R686 B.n419 B.n417 10.6151
R687 B.n420 B.n419 10.6151
R688 B.n421 B.n420 10.6151
R689 B.n422 B.n421 10.6151
R690 B.n424 B.n422 10.6151
R691 B.n425 B.n424 10.6151
R692 B.n426 B.n425 10.6151
R693 B.n427 B.n426 10.6151
R694 B.n429 B.n427 10.6151
R695 B.n430 B.n429 10.6151
R696 B.n431 B.n430 10.6151
R697 B.n369 B.n368 10.6151
R698 B.n368 B.n367 10.6151
R699 B.n367 B.n366 10.6151
R700 B.n366 B.n364 10.6151
R701 B.n364 B.n361 10.6151
R702 B.n361 B.n360 10.6151
R703 B.n360 B.n357 10.6151
R704 B.n357 B.n356 10.6151
R705 B.n356 B.n353 10.6151
R706 B.n353 B.n352 10.6151
R707 B.n352 B.n349 10.6151
R708 B.n349 B.n348 10.6151
R709 B.n348 B.n345 10.6151
R710 B.n345 B.n344 10.6151
R711 B.n344 B.n341 10.6151
R712 B.n341 B.n340 10.6151
R713 B.n340 B.n337 10.6151
R714 B.n337 B.n336 10.6151
R715 B.n336 B.n333 10.6151
R716 B.n333 B.n332 10.6151
R717 B.n332 B.n329 10.6151
R718 B.n329 B.n328 10.6151
R719 B.n328 B.n325 10.6151
R720 B.n325 B.n324 10.6151
R721 B.n324 B.n321 10.6151
R722 B.n321 B.n320 10.6151
R723 B.n317 B.n316 10.6151
R724 B.n316 B.n313 10.6151
R725 B.n313 B.n312 10.6151
R726 B.n312 B.n309 10.6151
R727 B.n309 B.n308 10.6151
R728 B.n308 B.n305 10.6151
R729 B.n305 B.n304 10.6151
R730 B.n304 B.n301 10.6151
R731 B.n299 B.n296 10.6151
R732 B.n296 B.n295 10.6151
R733 B.n295 B.n292 10.6151
R734 B.n292 B.n291 10.6151
R735 B.n291 B.n288 10.6151
R736 B.n288 B.n287 10.6151
R737 B.n287 B.n284 10.6151
R738 B.n284 B.n283 10.6151
R739 B.n283 B.n280 10.6151
R740 B.n280 B.n279 10.6151
R741 B.n279 B.n276 10.6151
R742 B.n276 B.n275 10.6151
R743 B.n275 B.n272 10.6151
R744 B.n272 B.n271 10.6151
R745 B.n271 B.n268 10.6151
R746 B.n268 B.n267 10.6151
R747 B.n267 B.n264 10.6151
R748 B.n264 B.n263 10.6151
R749 B.n263 B.n260 10.6151
R750 B.n260 B.n259 10.6151
R751 B.n259 B.n256 10.6151
R752 B.n256 B.n255 10.6151
R753 B.n255 B.n252 10.6151
R754 B.n252 B.n251 10.6151
R755 B.n251 B.n212 10.6151
R756 B.n375 B.n212 10.6151
R757 B.n381 B.n208 10.6151
R758 B.n382 B.n381 10.6151
R759 B.n383 B.n382 10.6151
R760 B.n383 B.n200 10.6151
R761 B.n393 B.n200 10.6151
R762 B.n394 B.n393 10.6151
R763 B.n395 B.n394 10.6151
R764 B.n395 B.n192 10.6151
R765 B.n407 B.n192 10.6151
R766 B.n408 B.n407 10.6151
R767 B.n409 B.n408 10.6151
R768 B.n409 B.n0 10.6151
R769 B.n456 B.n1 10.6151
R770 B.n456 B.n455 10.6151
R771 B.n455 B.n454 10.6151
R772 B.n454 B.n9 10.6151
R773 B.n448 B.n9 10.6151
R774 B.n448 B.n447 10.6151
R775 B.n447 B.n446 10.6151
R776 B.n446 B.n17 10.6151
R777 B.n440 B.n17 10.6151
R778 B.n440 B.n439 10.6151
R779 B.n439 B.n438 10.6151
R780 B.n438 B.n24 10.6151
R781 B.n120 B.n119 7.18099
R782 B.n136 B.n62 7.18099
R783 B.n317 B.n247 7.18099
R784 B.n301 B.n300 7.18099
R785 B.n119 B.n118 3.43465
R786 B.n139 B.n62 3.43465
R787 B.n320 B.n247 3.43465
R788 B.n300 B.n299 3.43465
R789 B.n462 B.n0 2.81026
R790 B.n462 B.n1 2.81026
R791 VP.n0 VP.t1 610.622
R792 VP.n0 VP.t0 575.338
R793 VP VP.n0 0.0516364
R794 VDD1 VDD1.t1 97.94
R795 VDD1 VDD1.t0 66.3657
C0 VDD2 VN 1.11144f
C1 VDD1 VN 0.148831f
C2 VTAIL VDD2 4.06492f
C3 VTAIL VDD1 4.03012f
C4 VDD2 VDD1 0.442093f
C5 VP VN 3.53595f
C6 VTAIL VP 0.851526f
C7 VP VDD2 0.246206f
C8 VP VDD1 1.20602f
C9 VTAIL VN 0.837089f
C10 VDD2 B 2.765902f
C11 VDD1 B 4.62206f
C12 VTAIL B 3.974728f
C13 VN B 6.05593f
C14 VP B 3.405639f
C15 VDD1.t0 B 0.9794f
C16 VDD1.t1 B 1.25575f
C17 VP.t1 B 0.511214f
C18 VP.t0 B 0.43647f
C19 VP.n0 B 2.5436f
C20 VDD2.t0 B 1.28961f
C21 VDD2.t1 B 1.01872f
C22 VDD2.n0 B 1.75819f
C23 VTAIL.t0 B 1.04688f
C24 VTAIL.n0 B 0.992493f
C25 VTAIL.t3 B 1.04689f
C26 VTAIL.n1 B 0.999806f
C27 VTAIL.t1 B 1.04688f
C28 VTAIL.n2 B 0.956427f
C29 VTAIL.t2 B 1.04688f
C30 VTAIL.n3 B 0.913567f
C31 VN.t1 B 0.429795f
C32 VN.t0 B 0.505607f
.ends

