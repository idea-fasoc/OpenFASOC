* NGSPICE file created from diff_pair_sample_0547.ext - technology: sky130A

.subckt diff_pair_sample_0547 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1444_n3284# sky130_fd_pr__pfet_01v8 ad=4.5162 pd=23.94 as=0 ps=0 w=11.58 l=0.46
X1 VTAIL.t7 VP.t0 VDD1.t1 w_n1444_n3284# sky130_fd_pr__pfet_01v8 ad=4.5162 pd=23.94 as=1.9107 ps=11.91 w=11.58 l=0.46
X2 B.t8 B.t6 B.t7 w_n1444_n3284# sky130_fd_pr__pfet_01v8 ad=4.5162 pd=23.94 as=0 ps=0 w=11.58 l=0.46
X3 B.t5 B.t3 B.t4 w_n1444_n3284# sky130_fd_pr__pfet_01v8 ad=4.5162 pd=23.94 as=0 ps=0 w=11.58 l=0.46
X4 VDD2.t3 VN.t0 VTAIL.t0 w_n1444_n3284# sky130_fd_pr__pfet_01v8 ad=1.9107 pd=11.91 as=4.5162 ps=23.94 w=11.58 l=0.46
X5 VDD1.t0 VP.t1 VTAIL.t6 w_n1444_n3284# sky130_fd_pr__pfet_01v8 ad=1.9107 pd=11.91 as=4.5162 ps=23.94 w=11.58 l=0.46
X6 VTAIL.t2 VN.t1 VDD2.t2 w_n1444_n3284# sky130_fd_pr__pfet_01v8 ad=4.5162 pd=23.94 as=1.9107 ps=11.91 w=11.58 l=0.46
X7 VTAIL.t1 VN.t2 VDD2.t1 w_n1444_n3284# sky130_fd_pr__pfet_01v8 ad=4.5162 pd=23.94 as=1.9107 ps=11.91 w=11.58 l=0.46
X8 VTAIL.t5 VP.t2 VDD1.t3 w_n1444_n3284# sky130_fd_pr__pfet_01v8 ad=4.5162 pd=23.94 as=1.9107 ps=11.91 w=11.58 l=0.46
X9 VDD2.t0 VN.t3 VTAIL.t3 w_n1444_n3284# sky130_fd_pr__pfet_01v8 ad=1.9107 pd=11.91 as=4.5162 ps=23.94 w=11.58 l=0.46
X10 VDD1.t2 VP.t3 VTAIL.t4 w_n1444_n3284# sky130_fd_pr__pfet_01v8 ad=1.9107 pd=11.91 as=4.5162 ps=23.94 w=11.58 l=0.46
X11 B.t2 B.t0 B.t1 w_n1444_n3284# sky130_fd_pr__pfet_01v8 ad=4.5162 pd=23.94 as=0 ps=0 w=11.58 l=0.46
R0 B.n95 B.t3 814.148
R1 B.n103 B.t0 814.148
R2 B.n30 B.t9 814.148
R3 B.n38 B.t6 814.148
R4 B.n336 B.n59 585
R5 B.n338 B.n337 585
R6 B.n339 B.n58 585
R7 B.n341 B.n340 585
R8 B.n342 B.n57 585
R9 B.n344 B.n343 585
R10 B.n345 B.n56 585
R11 B.n347 B.n346 585
R12 B.n348 B.n55 585
R13 B.n350 B.n349 585
R14 B.n351 B.n54 585
R15 B.n353 B.n352 585
R16 B.n354 B.n53 585
R17 B.n356 B.n355 585
R18 B.n357 B.n52 585
R19 B.n359 B.n358 585
R20 B.n360 B.n51 585
R21 B.n362 B.n361 585
R22 B.n363 B.n50 585
R23 B.n365 B.n364 585
R24 B.n366 B.n49 585
R25 B.n368 B.n367 585
R26 B.n369 B.n48 585
R27 B.n371 B.n370 585
R28 B.n372 B.n47 585
R29 B.n374 B.n373 585
R30 B.n375 B.n46 585
R31 B.n377 B.n376 585
R32 B.n378 B.n45 585
R33 B.n380 B.n379 585
R34 B.n381 B.n44 585
R35 B.n383 B.n382 585
R36 B.n384 B.n43 585
R37 B.n386 B.n385 585
R38 B.n387 B.n42 585
R39 B.n389 B.n388 585
R40 B.n390 B.n41 585
R41 B.n392 B.n391 585
R42 B.n393 B.n37 585
R43 B.n395 B.n394 585
R44 B.n396 B.n36 585
R45 B.n398 B.n397 585
R46 B.n399 B.n35 585
R47 B.n401 B.n400 585
R48 B.n402 B.n34 585
R49 B.n404 B.n403 585
R50 B.n405 B.n33 585
R51 B.n407 B.n406 585
R52 B.n408 B.n32 585
R53 B.n410 B.n409 585
R54 B.n412 B.n29 585
R55 B.n414 B.n413 585
R56 B.n415 B.n28 585
R57 B.n417 B.n416 585
R58 B.n418 B.n27 585
R59 B.n420 B.n419 585
R60 B.n421 B.n26 585
R61 B.n423 B.n422 585
R62 B.n424 B.n25 585
R63 B.n426 B.n425 585
R64 B.n427 B.n24 585
R65 B.n429 B.n428 585
R66 B.n430 B.n23 585
R67 B.n432 B.n431 585
R68 B.n433 B.n22 585
R69 B.n435 B.n434 585
R70 B.n436 B.n21 585
R71 B.n438 B.n437 585
R72 B.n439 B.n20 585
R73 B.n441 B.n440 585
R74 B.n442 B.n19 585
R75 B.n444 B.n443 585
R76 B.n445 B.n18 585
R77 B.n447 B.n446 585
R78 B.n448 B.n17 585
R79 B.n450 B.n449 585
R80 B.n451 B.n16 585
R81 B.n453 B.n452 585
R82 B.n454 B.n15 585
R83 B.n456 B.n455 585
R84 B.n457 B.n14 585
R85 B.n459 B.n458 585
R86 B.n460 B.n13 585
R87 B.n462 B.n461 585
R88 B.n463 B.n12 585
R89 B.n465 B.n464 585
R90 B.n466 B.n11 585
R91 B.n468 B.n467 585
R92 B.n469 B.n10 585
R93 B.n471 B.n470 585
R94 B.n335 B.n334 585
R95 B.n333 B.n60 585
R96 B.n332 B.n331 585
R97 B.n330 B.n61 585
R98 B.n329 B.n328 585
R99 B.n327 B.n62 585
R100 B.n326 B.n325 585
R101 B.n324 B.n63 585
R102 B.n323 B.n322 585
R103 B.n321 B.n64 585
R104 B.n320 B.n319 585
R105 B.n318 B.n65 585
R106 B.n317 B.n316 585
R107 B.n315 B.n66 585
R108 B.n314 B.n313 585
R109 B.n312 B.n67 585
R110 B.n311 B.n310 585
R111 B.n309 B.n68 585
R112 B.n308 B.n307 585
R113 B.n306 B.n69 585
R114 B.n305 B.n304 585
R115 B.n303 B.n70 585
R116 B.n302 B.n301 585
R117 B.n300 B.n71 585
R118 B.n299 B.n298 585
R119 B.n297 B.n72 585
R120 B.n296 B.n295 585
R121 B.n294 B.n73 585
R122 B.n293 B.n292 585
R123 B.n291 B.n74 585
R124 B.n290 B.n289 585
R125 B.n153 B.n124 585
R126 B.n155 B.n154 585
R127 B.n156 B.n123 585
R128 B.n158 B.n157 585
R129 B.n159 B.n122 585
R130 B.n161 B.n160 585
R131 B.n162 B.n121 585
R132 B.n164 B.n163 585
R133 B.n165 B.n120 585
R134 B.n167 B.n166 585
R135 B.n168 B.n119 585
R136 B.n170 B.n169 585
R137 B.n171 B.n118 585
R138 B.n173 B.n172 585
R139 B.n174 B.n117 585
R140 B.n176 B.n175 585
R141 B.n177 B.n116 585
R142 B.n179 B.n178 585
R143 B.n180 B.n115 585
R144 B.n182 B.n181 585
R145 B.n183 B.n114 585
R146 B.n185 B.n184 585
R147 B.n186 B.n113 585
R148 B.n188 B.n187 585
R149 B.n189 B.n112 585
R150 B.n191 B.n190 585
R151 B.n192 B.n111 585
R152 B.n194 B.n193 585
R153 B.n195 B.n110 585
R154 B.n197 B.n196 585
R155 B.n198 B.n109 585
R156 B.n200 B.n199 585
R157 B.n201 B.n108 585
R158 B.n203 B.n202 585
R159 B.n204 B.n107 585
R160 B.n206 B.n205 585
R161 B.n207 B.n106 585
R162 B.n209 B.n208 585
R163 B.n210 B.n105 585
R164 B.n212 B.n211 585
R165 B.n214 B.n102 585
R166 B.n216 B.n215 585
R167 B.n217 B.n101 585
R168 B.n219 B.n218 585
R169 B.n220 B.n100 585
R170 B.n222 B.n221 585
R171 B.n223 B.n99 585
R172 B.n225 B.n224 585
R173 B.n226 B.n98 585
R174 B.n228 B.n227 585
R175 B.n230 B.n229 585
R176 B.n231 B.n94 585
R177 B.n233 B.n232 585
R178 B.n234 B.n93 585
R179 B.n236 B.n235 585
R180 B.n237 B.n92 585
R181 B.n239 B.n238 585
R182 B.n240 B.n91 585
R183 B.n242 B.n241 585
R184 B.n243 B.n90 585
R185 B.n245 B.n244 585
R186 B.n246 B.n89 585
R187 B.n248 B.n247 585
R188 B.n249 B.n88 585
R189 B.n251 B.n250 585
R190 B.n252 B.n87 585
R191 B.n254 B.n253 585
R192 B.n255 B.n86 585
R193 B.n257 B.n256 585
R194 B.n258 B.n85 585
R195 B.n260 B.n259 585
R196 B.n261 B.n84 585
R197 B.n263 B.n262 585
R198 B.n264 B.n83 585
R199 B.n266 B.n265 585
R200 B.n267 B.n82 585
R201 B.n269 B.n268 585
R202 B.n270 B.n81 585
R203 B.n272 B.n271 585
R204 B.n273 B.n80 585
R205 B.n275 B.n274 585
R206 B.n276 B.n79 585
R207 B.n278 B.n277 585
R208 B.n279 B.n78 585
R209 B.n281 B.n280 585
R210 B.n282 B.n77 585
R211 B.n284 B.n283 585
R212 B.n285 B.n76 585
R213 B.n287 B.n286 585
R214 B.n288 B.n75 585
R215 B.n152 B.n151 585
R216 B.n150 B.n125 585
R217 B.n149 B.n148 585
R218 B.n147 B.n126 585
R219 B.n146 B.n145 585
R220 B.n144 B.n127 585
R221 B.n143 B.n142 585
R222 B.n141 B.n128 585
R223 B.n140 B.n139 585
R224 B.n138 B.n129 585
R225 B.n137 B.n136 585
R226 B.n135 B.n130 585
R227 B.n134 B.n133 585
R228 B.n132 B.n131 585
R229 B.n2 B.n0 585
R230 B.n493 B.n1 585
R231 B.n492 B.n491 585
R232 B.n490 B.n3 585
R233 B.n489 B.n488 585
R234 B.n487 B.n4 585
R235 B.n486 B.n485 585
R236 B.n484 B.n5 585
R237 B.n483 B.n482 585
R238 B.n481 B.n6 585
R239 B.n480 B.n479 585
R240 B.n478 B.n7 585
R241 B.n477 B.n476 585
R242 B.n475 B.n8 585
R243 B.n474 B.n473 585
R244 B.n472 B.n9 585
R245 B.n495 B.n494 585
R246 B.n151 B.n124 540.549
R247 B.n470 B.n9 540.549
R248 B.n289 B.n288 540.549
R249 B.n336 B.n335 540.549
R250 B.n151 B.n150 163.367
R251 B.n150 B.n149 163.367
R252 B.n149 B.n126 163.367
R253 B.n145 B.n126 163.367
R254 B.n145 B.n144 163.367
R255 B.n144 B.n143 163.367
R256 B.n143 B.n128 163.367
R257 B.n139 B.n128 163.367
R258 B.n139 B.n138 163.367
R259 B.n138 B.n137 163.367
R260 B.n137 B.n130 163.367
R261 B.n133 B.n130 163.367
R262 B.n133 B.n132 163.367
R263 B.n132 B.n2 163.367
R264 B.n494 B.n2 163.367
R265 B.n494 B.n493 163.367
R266 B.n493 B.n492 163.367
R267 B.n492 B.n3 163.367
R268 B.n488 B.n3 163.367
R269 B.n488 B.n487 163.367
R270 B.n487 B.n486 163.367
R271 B.n486 B.n5 163.367
R272 B.n482 B.n5 163.367
R273 B.n482 B.n481 163.367
R274 B.n481 B.n480 163.367
R275 B.n480 B.n7 163.367
R276 B.n476 B.n7 163.367
R277 B.n476 B.n475 163.367
R278 B.n475 B.n474 163.367
R279 B.n474 B.n9 163.367
R280 B.n155 B.n124 163.367
R281 B.n156 B.n155 163.367
R282 B.n157 B.n156 163.367
R283 B.n157 B.n122 163.367
R284 B.n161 B.n122 163.367
R285 B.n162 B.n161 163.367
R286 B.n163 B.n162 163.367
R287 B.n163 B.n120 163.367
R288 B.n167 B.n120 163.367
R289 B.n168 B.n167 163.367
R290 B.n169 B.n168 163.367
R291 B.n169 B.n118 163.367
R292 B.n173 B.n118 163.367
R293 B.n174 B.n173 163.367
R294 B.n175 B.n174 163.367
R295 B.n175 B.n116 163.367
R296 B.n179 B.n116 163.367
R297 B.n180 B.n179 163.367
R298 B.n181 B.n180 163.367
R299 B.n181 B.n114 163.367
R300 B.n185 B.n114 163.367
R301 B.n186 B.n185 163.367
R302 B.n187 B.n186 163.367
R303 B.n187 B.n112 163.367
R304 B.n191 B.n112 163.367
R305 B.n192 B.n191 163.367
R306 B.n193 B.n192 163.367
R307 B.n193 B.n110 163.367
R308 B.n197 B.n110 163.367
R309 B.n198 B.n197 163.367
R310 B.n199 B.n198 163.367
R311 B.n199 B.n108 163.367
R312 B.n203 B.n108 163.367
R313 B.n204 B.n203 163.367
R314 B.n205 B.n204 163.367
R315 B.n205 B.n106 163.367
R316 B.n209 B.n106 163.367
R317 B.n210 B.n209 163.367
R318 B.n211 B.n210 163.367
R319 B.n211 B.n102 163.367
R320 B.n216 B.n102 163.367
R321 B.n217 B.n216 163.367
R322 B.n218 B.n217 163.367
R323 B.n218 B.n100 163.367
R324 B.n222 B.n100 163.367
R325 B.n223 B.n222 163.367
R326 B.n224 B.n223 163.367
R327 B.n224 B.n98 163.367
R328 B.n228 B.n98 163.367
R329 B.n229 B.n228 163.367
R330 B.n229 B.n94 163.367
R331 B.n233 B.n94 163.367
R332 B.n234 B.n233 163.367
R333 B.n235 B.n234 163.367
R334 B.n235 B.n92 163.367
R335 B.n239 B.n92 163.367
R336 B.n240 B.n239 163.367
R337 B.n241 B.n240 163.367
R338 B.n241 B.n90 163.367
R339 B.n245 B.n90 163.367
R340 B.n246 B.n245 163.367
R341 B.n247 B.n246 163.367
R342 B.n247 B.n88 163.367
R343 B.n251 B.n88 163.367
R344 B.n252 B.n251 163.367
R345 B.n253 B.n252 163.367
R346 B.n253 B.n86 163.367
R347 B.n257 B.n86 163.367
R348 B.n258 B.n257 163.367
R349 B.n259 B.n258 163.367
R350 B.n259 B.n84 163.367
R351 B.n263 B.n84 163.367
R352 B.n264 B.n263 163.367
R353 B.n265 B.n264 163.367
R354 B.n265 B.n82 163.367
R355 B.n269 B.n82 163.367
R356 B.n270 B.n269 163.367
R357 B.n271 B.n270 163.367
R358 B.n271 B.n80 163.367
R359 B.n275 B.n80 163.367
R360 B.n276 B.n275 163.367
R361 B.n277 B.n276 163.367
R362 B.n277 B.n78 163.367
R363 B.n281 B.n78 163.367
R364 B.n282 B.n281 163.367
R365 B.n283 B.n282 163.367
R366 B.n283 B.n76 163.367
R367 B.n287 B.n76 163.367
R368 B.n288 B.n287 163.367
R369 B.n289 B.n74 163.367
R370 B.n293 B.n74 163.367
R371 B.n294 B.n293 163.367
R372 B.n295 B.n294 163.367
R373 B.n295 B.n72 163.367
R374 B.n299 B.n72 163.367
R375 B.n300 B.n299 163.367
R376 B.n301 B.n300 163.367
R377 B.n301 B.n70 163.367
R378 B.n305 B.n70 163.367
R379 B.n306 B.n305 163.367
R380 B.n307 B.n306 163.367
R381 B.n307 B.n68 163.367
R382 B.n311 B.n68 163.367
R383 B.n312 B.n311 163.367
R384 B.n313 B.n312 163.367
R385 B.n313 B.n66 163.367
R386 B.n317 B.n66 163.367
R387 B.n318 B.n317 163.367
R388 B.n319 B.n318 163.367
R389 B.n319 B.n64 163.367
R390 B.n323 B.n64 163.367
R391 B.n324 B.n323 163.367
R392 B.n325 B.n324 163.367
R393 B.n325 B.n62 163.367
R394 B.n329 B.n62 163.367
R395 B.n330 B.n329 163.367
R396 B.n331 B.n330 163.367
R397 B.n331 B.n60 163.367
R398 B.n335 B.n60 163.367
R399 B.n470 B.n469 163.367
R400 B.n469 B.n468 163.367
R401 B.n468 B.n11 163.367
R402 B.n464 B.n11 163.367
R403 B.n464 B.n463 163.367
R404 B.n463 B.n462 163.367
R405 B.n462 B.n13 163.367
R406 B.n458 B.n13 163.367
R407 B.n458 B.n457 163.367
R408 B.n457 B.n456 163.367
R409 B.n456 B.n15 163.367
R410 B.n452 B.n15 163.367
R411 B.n452 B.n451 163.367
R412 B.n451 B.n450 163.367
R413 B.n450 B.n17 163.367
R414 B.n446 B.n17 163.367
R415 B.n446 B.n445 163.367
R416 B.n445 B.n444 163.367
R417 B.n444 B.n19 163.367
R418 B.n440 B.n19 163.367
R419 B.n440 B.n439 163.367
R420 B.n439 B.n438 163.367
R421 B.n438 B.n21 163.367
R422 B.n434 B.n21 163.367
R423 B.n434 B.n433 163.367
R424 B.n433 B.n432 163.367
R425 B.n432 B.n23 163.367
R426 B.n428 B.n23 163.367
R427 B.n428 B.n427 163.367
R428 B.n427 B.n426 163.367
R429 B.n426 B.n25 163.367
R430 B.n422 B.n25 163.367
R431 B.n422 B.n421 163.367
R432 B.n421 B.n420 163.367
R433 B.n420 B.n27 163.367
R434 B.n416 B.n27 163.367
R435 B.n416 B.n415 163.367
R436 B.n415 B.n414 163.367
R437 B.n414 B.n29 163.367
R438 B.n409 B.n29 163.367
R439 B.n409 B.n408 163.367
R440 B.n408 B.n407 163.367
R441 B.n407 B.n33 163.367
R442 B.n403 B.n33 163.367
R443 B.n403 B.n402 163.367
R444 B.n402 B.n401 163.367
R445 B.n401 B.n35 163.367
R446 B.n397 B.n35 163.367
R447 B.n397 B.n396 163.367
R448 B.n396 B.n395 163.367
R449 B.n395 B.n37 163.367
R450 B.n391 B.n37 163.367
R451 B.n391 B.n390 163.367
R452 B.n390 B.n389 163.367
R453 B.n389 B.n42 163.367
R454 B.n385 B.n42 163.367
R455 B.n385 B.n384 163.367
R456 B.n384 B.n383 163.367
R457 B.n383 B.n44 163.367
R458 B.n379 B.n44 163.367
R459 B.n379 B.n378 163.367
R460 B.n378 B.n377 163.367
R461 B.n377 B.n46 163.367
R462 B.n373 B.n46 163.367
R463 B.n373 B.n372 163.367
R464 B.n372 B.n371 163.367
R465 B.n371 B.n48 163.367
R466 B.n367 B.n48 163.367
R467 B.n367 B.n366 163.367
R468 B.n366 B.n365 163.367
R469 B.n365 B.n50 163.367
R470 B.n361 B.n50 163.367
R471 B.n361 B.n360 163.367
R472 B.n360 B.n359 163.367
R473 B.n359 B.n52 163.367
R474 B.n355 B.n52 163.367
R475 B.n355 B.n354 163.367
R476 B.n354 B.n353 163.367
R477 B.n353 B.n54 163.367
R478 B.n349 B.n54 163.367
R479 B.n349 B.n348 163.367
R480 B.n348 B.n347 163.367
R481 B.n347 B.n56 163.367
R482 B.n343 B.n56 163.367
R483 B.n343 B.n342 163.367
R484 B.n342 B.n341 163.367
R485 B.n341 B.n58 163.367
R486 B.n337 B.n58 163.367
R487 B.n337 B.n336 163.367
R488 B.n95 B.t5 122.913
R489 B.n38 B.t7 122.913
R490 B.n103 B.t2 122.9
R491 B.n30 B.t10 122.9
R492 B.n96 B.t4 107.593
R493 B.n39 B.t8 107.593
R494 B.n104 B.t1 107.579
R495 B.n31 B.t11 107.579
R496 B.n97 B.n96 59.5399
R497 B.n213 B.n104 59.5399
R498 B.n411 B.n31 59.5399
R499 B.n40 B.n39 59.5399
R500 B.n472 B.n471 35.1225
R501 B.n290 B.n75 35.1225
R502 B.n153 B.n152 35.1225
R503 B.n334 B.n59 35.1224
R504 B B.n495 18.0485
R505 B.n96 B.n95 15.3217
R506 B.n104 B.n103 15.3217
R507 B.n31 B.n30 15.3217
R508 B.n39 B.n38 15.3217
R509 B.n471 B.n10 10.6151
R510 B.n467 B.n10 10.6151
R511 B.n467 B.n466 10.6151
R512 B.n466 B.n465 10.6151
R513 B.n465 B.n12 10.6151
R514 B.n461 B.n12 10.6151
R515 B.n461 B.n460 10.6151
R516 B.n460 B.n459 10.6151
R517 B.n459 B.n14 10.6151
R518 B.n455 B.n14 10.6151
R519 B.n455 B.n454 10.6151
R520 B.n454 B.n453 10.6151
R521 B.n453 B.n16 10.6151
R522 B.n449 B.n16 10.6151
R523 B.n449 B.n448 10.6151
R524 B.n448 B.n447 10.6151
R525 B.n447 B.n18 10.6151
R526 B.n443 B.n18 10.6151
R527 B.n443 B.n442 10.6151
R528 B.n442 B.n441 10.6151
R529 B.n441 B.n20 10.6151
R530 B.n437 B.n20 10.6151
R531 B.n437 B.n436 10.6151
R532 B.n436 B.n435 10.6151
R533 B.n435 B.n22 10.6151
R534 B.n431 B.n22 10.6151
R535 B.n431 B.n430 10.6151
R536 B.n430 B.n429 10.6151
R537 B.n429 B.n24 10.6151
R538 B.n425 B.n24 10.6151
R539 B.n425 B.n424 10.6151
R540 B.n424 B.n423 10.6151
R541 B.n423 B.n26 10.6151
R542 B.n419 B.n26 10.6151
R543 B.n419 B.n418 10.6151
R544 B.n418 B.n417 10.6151
R545 B.n417 B.n28 10.6151
R546 B.n413 B.n28 10.6151
R547 B.n413 B.n412 10.6151
R548 B.n410 B.n32 10.6151
R549 B.n406 B.n32 10.6151
R550 B.n406 B.n405 10.6151
R551 B.n405 B.n404 10.6151
R552 B.n404 B.n34 10.6151
R553 B.n400 B.n34 10.6151
R554 B.n400 B.n399 10.6151
R555 B.n399 B.n398 10.6151
R556 B.n398 B.n36 10.6151
R557 B.n394 B.n393 10.6151
R558 B.n393 B.n392 10.6151
R559 B.n392 B.n41 10.6151
R560 B.n388 B.n41 10.6151
R561 B.n388 B.n387 10.6151
R562 B.n387 B.n386 10.6151
R563 B.n386 B.n43 10.6151
R564 B.n382 B.n43 10.6151
R565 B.n382 B.n381 10.6151
R566 B.n381 B.n380 10.6151
R567 B.n380 B.n45 10.6151
R568 B.n376 B.n45 10.6151
R569 B.n376 B.n375 10.6151
R570 B.n375 B.n374 10.6151
R571 B.n374 B.n47 10.6151
R572 B.n370 B.n47 10.6151
R573 B.n370 B.n369 10.6151
R574 B.n369 B.n368 10.6151
R575 B.n368 B.n49 10.6151
R576 B.n364 B.n49 10.6151
R577 B.n364 B.n363 10.6151
R578 B.n363 B.n362 10.6151
R579 B.n362 B.n51 10.6151
R580 B.n358 B.n51 10.6151
R581 B.n358 B.n357 10.6151
R582 B.n357 B.n356 10.6151
R583 B.n356 B.n53 10.6151
R584 B.n352 B.n53 10.6151
R585 B.n352 B.n351 10.6151
R586 B.n351 B.n350 10.6151
R587 B.n350 B.n55 10.6151
R588 B.n346 B.n55 10.6151
R589 B.n346 B.n345 10.6151
R590 B.n345 B.n344 10.6151
R591 B.n344 B.n57 10.6151
R592 B.n340 B.n57 10.6151
R593 B.n340 B.n339 10.6151
R594 B.n339 B.n338 10.6151
R595 B.n338 B.n59 10.6151
R596 B.n291 B.n290 10.6151
R597 B.n292 B.n291 10.6151
R598 B.n292 B.n73 10.6151
R599 B.n296 B.n73 10.6151
R600 B.n297 B.n296 10.6151
R601 B.n298 B.n297 10.6151
R602 B.n298 B.n71 10.6151
R603 B.n302 B.n71 10.6151
R604 B.n303 B.n302 10.6151
R605 B.n304 B.n303 10.6151
R606 B.n304 B.n69 10.6151
R607 B.n308 B.n69 10.6151
R608 B.n309 B.n308 10.6151
R609 B.n310 B.n309 10.6151
R610 B.n310 B.n67 10.6151
R611 B.n314 B.n67 10.6151
R612 B.n315 B.n314 10.6151
R613 B.n316 B.n315 10.6151
R614 B.n316 B.n65 10.6151
R615 B.n320 B.n65 10.6151
R616 B.n321 B.n320 10.6151
R617 B.n322 B.n321 10.6151
R618 B.n322 B.n63 10.6151
R619 B.n326 B.n63 10.6151
R620 B.n327 B.n326 10.6151
R621 B.n328 B.n327 10.6151
R622 B.n328 B.n61 10.6151
R623 B.n332 B.n61 10.6151
R624 B.n333 B.n332 10.6151
R625 B.n334 B.n333 10.6151
R626 B.n154 B.n153 10.6151
R627 B.n154 B.n123 10.6151
R628 B.n158 B.n123 10.6151
R629 B.n159 B.n158 10.6151
R630 B.n160 B.n159 10.6151
R631 B.n160 B.n121 10.6151
R632 B.n164 B.n121 10.6151
R633 B.n165 B.n164 10.6151
R634 B.n166 B.n165 10.6151
R635 B.n166 B.n119 10.6151
R636 B.n170 B.n119 10.6151
R637 B.n171 B.n170 10.6151
R638 B.n172 B.n171 10.6151
R639 B.n172 B.n117 10.6151
R640 B.n176 B.n117 10.6151
R641 B.n177 B.n176 10.6151
R642 B.n178 B.n177 10.6151
R643 B.n178 B.n115 10.6151
R644 B.n182 B.n115 10.6151
R645 B.n183 B.n182 10.6151
R646 B.n184 B.n183 10.6151
R647 B.n184 B.n113 10.6151
R648 B.n188 B.n113 10.6151
R649 B.n189 B.n188 10.6151
R650 B.n190 B.n189 10.6151
R651 B.n190 B.n111 10.6151
R652 B.n194 B.n111 10.6151
R653 B.n195 B.n194 10.6151
R654 B.n196 B.n195 10.6151
R655 B.n196 B.n109 10.6151
R656 B.n200 B.n109 10.6151
R657 B.n201 B.n200 10.6151
R658 B.n202 B.n201 10.6151
R659 B.n202 B.n107 10.6151
R660 B.n206 B.n107 10.6151
R661 B.n207 B.n206 10.6151
R662 B.n208 B.n207 10.6151
R663 B.n208 B.n105 10.6151
R664 B.n212 B.n105 10.6151
R665 B.n215 B.n214 10.6151
R666 B.n215 B.n101 10.6151
R667 B.n219 B.n101 10.6151
R668 B.n220 B.n219 10.6151
R669 B.n221 B.n220 10.6151
R670 B.n221 B.n99 10.6151
R671 B.n225 B.n99 10.6151
R672 B.n226 B.n225 10.6151
R673 B.n227 B.n226 10.6151
R674 B.n231 B.n230 10.6151
R675 B.n232 B.n231 10.6151
R676 B.n232 B.n93 10.6151
R677 B.n236 B.n93 10.6151
R678 B.n237 B.n236 10.6151
R679 B.n238 B.n237 10.6151
R680 B.n238 B.n91 10.6151
R681 B.n242 B.n91 10.6151
R682 B.n243 B.n242 10.6151
R683 B.n244 B.n243 10.6151
R684 B.n244 B.n89 10.6151
R685 B.n248 B.n89 10.6151
R686 B.n249 B.n248 10.6151
R687 B.n250 B.n249 10.6151
R688 B.n250 B.n87 10.6151
R689 B.n254 B.n87 10.6151
R690 B.n255 B.n254 10.6151
R691 B.n256 B.n255 10.6151
R692 B.n256 B.n85 10.6151
R693 B.n260 B.n85 10.6151
R694 B.n261 B.n260 10.6151
R695 B.n262 B.n261 10.6151
R696 B.n262 B.n83 10.6151
R697 B.n266 B.n83 10.6151
R698 B.n267 B.n266 10.6151
R699 B.n268 B.n267 10.6151
R700 B.n268 B.n81 10.6151
R701 B.n272 B.n81 10.6151
R702 B.n273 B.n272 10.6151
R703 B.n274 B.n273 10.6151
R704 B.n274 B.n79 10.6151
R705 B.n278 B.n79 10.6151
R706 B.n279 B.n278 10.6151
R707 B.n280 B.n279 10.6151
R708 B.n280 B.n77 10.6151
R709 B.n284 B.n77 10.6151
R710 B.n285 B.n284 10.6151
R711 B.n286 B.n285 10.6151
R712 B.n286 B.n75 10.6151
R713 B.n152 B.n125 10.6151
R714 B.n148 B.n125 10.6151
R715 B.n148 B.n147 10.6151
R716 B.n147 B.n146 10.6151
R717 B.n146 B.n127 10.6151
R718 B.n142 B.n127 10.6151
R719 B.n142 B.n141 10.6151
R720 B.n141 B.n140 10.6151
R721 B.n140 B.n129 10.6151
R722 B.n136 B.n129 10.6151
R723 B.n136 B.n135 10.6151
R724 B.n135 B.n134 10.6151
R725 B.n134 B.n131 10.6151
R726 B.n131 B.n0 10.6151
R727 B.n491 B.n1 10.6151
R728 B.n491 B.n490 10.6151
R729 B.n490 B.n489 10.6151
R730 B.n489 B.n4 10.6151
R731 B.n485 B.n4 10.6151
R732 B.n485 B.n484 10.6151
R733 B.n484 B.n483 10.6151
R734 B.n483 B.n6 10.6151
R735 B.n479 B.n6 10.6151
R736 B.n479 B.n478 10.6151
R737 B.n478 B.n477 10.6151
R738 B.n477 B.n8 10.6151
R739 B.n473 B.n8 10.6151
R740 B.n473 B.n472 10.6151
R741 B.n412 B.n411 9.36635
R742 B.n394 B.n40 9.36635
R743 B.n213 B.n212 9.36635
R744 B.n230 B.n97 9.36635
R745 B.n495 B.n0 2.81026
R746 B.n495 B.n1 2.81026
R747 B.n411 B.n410 1.24928
R748 B.n40 B.n36 1.24928
R749 B.n214 B.n213 1.24928
R750 B.n227 B.n97 1.24928
R751 VP.n0 VP.t2 713.072
R752 VP.n0 VP.t1 713.047
R753 VP.n2 VP.t0 692.09
R754 VP.n3 VP.t3 692.09
R755 VP.n4 VP.n3 161.3
R756 VP.n2 VP.n1 161.3
R757 VP.n1 VP.n0 109.585
R758 VP.n3 VP.n2 48.2005
R759 VP.n4 VP.n1 0.189894
R760 VP VP.n4 0.0516364
R761 VDD1 VDD1.n1 113.591
R762 VDD1 VDD1.n0 77.383
R763 VDD1.n0 VDD1.t3 2.80749
R764 VDD1.n0 VDD1.t0 2.80749
R765 VDD1.n1 VDD1.t1 2.80749
R766 VDD1.n1 VDD1.t2 2.80749
R767 VTAIL.n5 VTAIL.t5 63.4542
R768 VTAIL.n4 VTAIL.t0 63.4542
R769 VTAIL.n3 VTAIL.t2 63.4542
R770 VTAIL.n7 VTAIL.t3 63.4532
R771 VTAIL.n0 VTAIL.t1 63.4532
R772 VTAIL.n1 VTAIL.t4 63.4532
R773 VTAIL.n2 VTAIL.t7 63.4532
R774 VTAIL.n6 VTAIL.t6 63.453
R775 VTAIL.n7 VTAIL.n6 23.0307
R776 VTAIL.n3 VTAIL.n2 23.0307
R777 VTAIL.n4 VTAIL.n3 0.681535
R778 VTAIL.n6 VTAIL.n5 0.681535
R779 VTAIL.n2 VTAIL.n1 0.681535
R780 VTAIL.n5 VTAIL.n4 0.470328
R781 VTAIL.n1 VTAIL.n0 0.470328
R782 VTAIL VTAIL.n0 0.399207
R783 VTAIL VTAIL.n7 0.282828
R784 VN.n0 VN.t2 713.072
R785 VN.n1 VN.t0 713.072
R786 VN.n0 VN.t3 713.047
R787 VN.n1 VN.t1 713.047
R788 VN VN.n1 109.966
R789 VN VN.n0 70.265
R790 VDD2.n2 VDD2.n0 113.066
R791 VDD2.n2 VDD2.n1 77.3248
R792 VDD2.n1 VDD2.t2 2.80749
R793 VDD2.n1 VDD2.t3 2.80749
R794 VDD2.n0 VDD2.t1 2.80749
R795 VDD2.n0 VDD2.t0 2.80749
R796 VDD2 VDD2.n2 0.0586897
C0 VDD2 w_n1444_n3284# 1.00922f
C1 VDD2 VTAIL 7.77163f
C2 VDD1 w_n1444_n3284# 0.999348f
C3 w_n1444_n3284# B 6.49489f
C4 VTAIL VDD1 7.73177f
C5 VTAIL B 3.52005f
C6 VP VN 4.5706f
C7 VTAIL w_n1444_n3284# 4.09851f
C8 VDD2 VN 2.497f
C9 VN B 0.696339f
C10 VDD1 VN 0.147503f
C11 VN w_n1444_n3284# 2.0426f
C12 VTAIL VN 2.05397f
C13 VDD2 VP 0.25857f
C14 VP VDD1 2.60787f
C15 VP B 0.985445f
C16 VDD2 VDD1 0.51474f
C17 VDD2 B 0.890049f
C18 VP w_n1444_n3284# 2.22282f
C19 VTAIL VP 2.06807f
C20 VDD1 B 0.87188f
C21 VDD2 VSUBS 0.637434f
C22 VDD1 VSUBS 4.999456f
C23 VTAIL VSUBS 0.775441f
C24 VN VSUBS 6.10266f
C25 VP VSUBS 1.15628f
C26 B VSUBS 2.378699f
C27 w_n1444_n3284# VSUBS 58.4127f
C28 VDD2.t1 VSUBS 0.276568f
C29 VDD2.t0 VSUBS 0.276568f
C30 VDD2.n0 VSUBS 2.7985f
C31 VDD2.t2 VSUBS 0.276568f
C32 VDD2.t3 VSUBS 0.276568f
C33 VDD2.n1 VSUBS 2.17128f
C34 VDD2.n2 VSUBS 4.15111f
C35 VN.t2 VSUBS 1.0497f
C36 VN.t3 VSUBS 1.04968f
C37 VN.n0 VSUBS 0.819834f
C38 VN.t0 VSUBS 1.0497f
C39 VN.t1 VSUBS 1.04968f
C40 VN.n1 VSUBS 1.77649f
C41 VTAIL.t1 VSUBS 2.15019f
C42 VTAIL.n0 VSUBS 0.67484f
C43 VTAIL.t4 VSUBS 2.15019f
C44 VTAIL.n1 VSUBS 0.696992f
C45 VTAIL.t7 VSUBS 2.15019f
C46 VTAIL.n2 VSUBS 1.82763f
C47 VTAIL.t2 VSUBS 2.15019f
C48 VTAIL.n3 VSUBS 1.82763f
C49 VTAIL.t0 VSUBS 2.15019f
C50 VTAIL.n4 VSUBS 0.696986f
C51 VTAIL.t5 VSUBS 2.15019f
C52 VTAIL.n5 VSUBS 0.696986f
C53 VTAIL.t6 VSUBS 2.15018f
C54 VTAIL.n6 VSUBS 1.82764f
C55 VTAIL.t3 VSUBS 2.15019f
C56 VTAIL.n7 VSUBS 1.79635f
C57 VDD1.t3 VSUBS 0.273602f
C58 VDD1.t0 VSUBS 0.273602f
C59 VDD1.n0 VSUBS 2.14847f
C60 VDD1.t1 VSUBS 0.273602f
C61 VDD1.t2 VSUBS 0.273602f
C62 VDD1.n1 VSUBS 2.79413f
C63 VP.t1 VSUBS 1.08711f
C64 VP.t2 VSUBS 1.08712f
C65 VP.n0 VSUBS 1.81702f
C66 VP.n1 VSUBS 4.40407f
C67 VP.t0 VSUBS 1.07426f
C68 VP.n2 VSUBS 0.437297f
C69 VP.t3 VSUBS 1.07426f
C70 VP.n3 VSUBS 0.437297f
C71 VP.n4 VSUBS 0.054774f
C72 B.n0 VSUBS 0.005396f
C73 B.n1 VSUBS 0.005396f
C74 B.n2 VSUBS 0.008533f
C75 B.n3 VSUBS 0.008533f
C76 B.n4 VSUBS 0.008533f
C77 B.n5 VSUBS 0.008533f
C78 B.n6 VSUBS 0.008533f
C79 B.n7 VSUBS 0.008533f
C80 B.n8 VSUBS 0.008533f
C81 B.n9 VSUBS 0.02058f
C82 B.n10 VSUBS 0.008533f
C83 B.n11 VSUBS 0.008533f
C84 B.n12 VSUBS 0.008533f
C85 B.n13 VSUBS 0.008533f
C86 B.n14 VSUBS 0.008533f
C87 B.n15 VSUBS 0.008533f
C88 B.n16 VSUBS 0.008533f
C89 B.n17 VSUBS 0.008533f
C90 B.n18 VSUBS 0.008533f
C91 B.n19 VSUBS 0.008533f
C92 B.n20 VSUBS 0.008533f
C93 B.n21 VSUBS 0.008533f
C94 B.n22 VSUBS 0.008533f
C95 B.n23 VSUBS 0.008533f
C96 B.n24 VSUBS 0.008533f
C97 B.n25 VSUBS 0.008533f
C98 B.n26 VSUBS 0.008533f
C99 B.n27 VSUBS 0.008533f
C100 B.n28 VSUBS 0.008533f
C101 B.n29 VSUBS 0.008533f
C102 B.t11 VSUBS 0.458235f
C103 B.t10 VSUBS 0.466279f
C104 B.t9 VSUBS 0.261269f
C105 B.n30 VSUBS 0.135942f
C106 B.n31 VSUBS 0.076701f
C107 B.n32 VSUBS 0.008533f
C108 B.n33 VSUBS 0.008533f
C109 B.n34 VSUBS 0.008533f
C110 B.n35 VSUBS 0.008533f
C111 B.n36 VSUBS 0.004769f
C112 B.n37 VSUBS 0.008533f
C113 B.t8 VSUBS 0.458226f
C114 B.t7 VSUBS 0.466271f
C115 B.t6 VSUBS 0.261269f
C116 B.n38 VSUBS 0.135951f
C117 B.n39 VSUBS 0.07671f
C118 B.n40 VSUBS 0.019771f
C119 B.n41 VSUBS 0.008533f
C120 B.n42 VSUBS 0.008533f
C121 B.n43 VSUBS 0.008533f
C122 B.n44 VSUBS 0.008533f
C123 B.n45 VSUBS 0.008533f
C124 B.n46 VSUBS 0.008533f
C125 B.n47 VSUBS 0.008533f
C126 B.n48 VSUBS 0.008533f
C127 B.n49 VSUBS 0.008533f
C128 B.n50 VSUBS 0.008533f
C129 B.n51 VSUBS 0.008533f
C130 B.n52 VSUBS 0.008533f
C131 B.n53 VSUBS 0.008533f
C132 B.n54 VSUBS 0.008533f
C133 B.n55 VSUBS 0.008533f
C134 B.n56 VSUBS 0.008533f
C135 B.n57 VSUBS 0.008533f
C136 B.n58 VSUBS 0.008533f
C137 B.n59 VSUBS 0.020397f
C138 B.n60 VSUBS 0.008533f
C139 B.n61 VSUBS 0.008533f
C140 B.n62 VSUBS 0.008533f
C141 B.n63 VSUBS 0.008533f
C142 B.n64 VSUBS 0.008533f
C143 B.n65 VSUBS 0.008533f
C144 B.n66 VSUBS 0.008533f
C145 B.n67 VSUBS 0.008533f
C146 B.n68 VSUBS 0.008533f
C147 B.n69 VSUBS 0.008533f
C148 B.n70 VSUBS 0.008533f
C149 B.n71 VSUBS 0.008533f
C150 B.n72 VSUBS 0.008533f
C151 B.n73 VSUBS 0.008533f
C152 B.n74 VSUBS 0.008533f
C153 B.n75 VSUBS 0.021335f
C154 B.n76 VSUBS 0.008533f
C155 B.n77 VSUBS 0.008533f
C156 B.n78 VSUBS 0.008533f
C157 B.n79 VSUBS 0.008533f
C158 B.n80 VSUBS 0.008533f
C159 B.n81 VSUBS 0.008533f
C160 B.n82 VSUBS 0.008533f
C161 B.n83 VSUBS 0.008533f
C162 B.n84 VSUBS 0.008533f
C163 B.n85 VSUBS 0.008533f
C164 B.n86 VSUBS 0.008533f
C165 B.n87 VSUBS 0.008533f
C166 B.n88 VSUBS 0.008533f
C167 B.n89 VSUBS 0.008533f
C168 B.n90 VSUBS 0.008533f
C169 B.n91 VSUBS 0.008533f
C170 B.n92 VSUBS 0.008533f
C171 B.n93 VSUBS 0.008533f
C172 B.n94 VSUBS 0.008533f
C173 B.t4 VSUBS 0.458226f
C174 B.t5 VSUBS 0.466271f
C175 B.t3 VSUBS 0.261269f
C176 B.n95 VSUBS 0.135951f
C177 B.n96 VSUBS 0.07671f
C178 B.n97 VSUBS 0.019771f
C179 B.n98 VSUBS 0.008533f
C180 B.n99 VSUBS 0.008533f
C181 B.n100 VSUBS 0.008533f
C182 B.n101 VSUBS 0.008533f
C183 B.n102 VSUBS 0.008533f
C184 B.t1 VSUBS 0.458235f
C185 B.t2 VSUBS 0.466279f
C186 B.t0 VSUBS 0.261269f
C187 B.n103 VSUBS 0.135942f
C188 B.n104 VSUBS 0.076701f
C189 B.n105 VSUBS 0.008533f
C190 B.n106 VSUBS 0.008533f
C191 B.n107 VSUBS 0.008533f
C192 B.n108 VSUBS 0.008533f
C193 B.n109 VSUBS 0.008533f
C194 B.n110 VSUBS 0.008533f
C195 B.n111 VSUBS 0.008533f
C196 B.n112 VSUBS 0.008533f
C197 B.n113 VSUBS 0.008533f
C198 B.n114 VSUBS 0.008533f
C199 B.n115 VSUBS 0.008533f
C200 B.n116 VSUBS 0.008533f
C201 B.n117 VSUBS 0.008533f
C202 B.n118 VSUBS 0.008533f
C203 B.n119 VSUBS 0.008533f
C204 B.n120 VSUBS 0.008533f
C205 B.n121 VSUBS 0.008533f
C206 B.n122 VSUBS 0.008533f
C207 B.n123 VSUBS 0.008533f
C208 B.n124 VSUBS 0.021335f
C209 B.n125 VSUBS 0.008533f
C210 B.n126 VSUBS 0.008533f
C211 B.n127 VSUBS 0.008533f
C212 B.n128 VSUBS 0.008533f
C213 B.n129 VSUBS 0.008533f
C214 B.n130 VSUBS 0.008533f
C215 B.n131 VSUBS 0.008533f
C216 B.n132 VSUBS 0.008533f
C217 B.n133 VSUBS 0.008533f
C218 B.n134 VSUBS 0.008533f
C219 B.n135 VSUBS 0.008533f
C220 B.n136 VSUBS 0.008533f
C221 B.n137 VSUBS 0.008533f
C222 B.n138 VSUBS 0.008533f
C223 B.n139 VSUBS 0.008533f
C224 B.n140 VSUBS 0.008533f
C225 B.n141 VSUBS 0.008533f
C226 B.n142 VSUBS 0.008533f
C227 B.n143 VSUBS 0.008533f
C228 B.n144 VSUBS 0.008533f
C229 B.n145 VSUBS 0.008533f
C230 B.n146 VSUBS 0.008533f
C231 B.n147 VSUBS 0.008533f
C232 B.n148 VSUBS 0.008533f
C233 B.n149 VSUBS 0.008533f
C234 B.n150 VSUBS 0.008533f
C235 B.n151 VSUBS 0.02058f
C236 B.n152 VSUBS 0.02058f
C237 B.n153 VSUBS 0.021335f
C238 B.n154 VSUBS 0.008533f
C239 B.n155 VSUBS 0.008533f
C240 B.n156 VSUBS 0.008533f
C241 B.n157 VSUBS 0.008533f
C242 B.n158 VSUBS 0.008533f
C243 B.n159 VSUBS 0.008533f
C244 B.n160 VSUBS 0.008533f
C245 B.n161 VSUBS 0.008533f
C246 B.n162 VSUBS 0.008533f
C247 B.n163 VSUBS 0.008533f
C248 B.n164 VSUBS 0.008533f
C249 B.n165 VSUBS 0.008533f
C250 B.n166 VSUBS 0.008533f
C251 B.n167 VSUBS 0.008533f
C252 B.n168 VSUBS 0.008533f
C253 B.n169 VSUBS 0.008533f
C254 B.n170 VSUBS 0.008533f
C255 B.n171 VSUBS 0.008533f
C256 B.n172 VSUBS 0.008533f
C257 B.n173 VSUBS 0.008533f
C258 B.n174 VSUBS 0.008533f
C259 B.n175 VSUBS 0.008533f
C260 B.n176 VSUBS 0.008533f
C261 B.n177 VSUBS 0.008533f
C262 B.n178 VSUBS 0.008533f
C263 B.n179 VSUBS 0.008533f
C264 B.n180 VSUBS 0.008533f
C265 B.n181 VSUBS 0.008533f
C266 B.n182 VSUBS 0.008533f
C267 B.n183 VSUBS 0.008533f
C268 B.n184 VSUBS 0.008533f
C269 B.n185 VSUBS 0.008533f
C270 B.n186 VSUBS 0.008533f
C271 B.n187 VSUBS 0.008533f
C272 B.n188 VSUBS 0.008533f
C273 B.n189 VSUBS 0.008533f
C274 B.n190 VSUBS 0.008533f
C275 B.n191 VSUBS 0.008533f
C276 B.n192 VSUBS 0.008533f
C277 B.n193 VSUBS 0.008533f
C278 B.n194 VSUBS 0.008533f
C279 B.n195 VSUBS 0.008533f
C280 B.n196 VSUBS 0.008533f
C281 B.n197 VSUBS 0.008533f
C282 B.n198 VSUBS 0.008533f
C283 B.n199 VSUBS 0.008533f
C284 B.n200 VSUBS 0.008533f
C285 B.n201 VSUBS 0.008533f
C286 B.n202 VSUBS 0.008533f
C287 B.n203 VSUBS 0.008533f
C288 B.n204 VSUBS 0.008533f
C289 B.n205 VSUBS 0.008533f
C290 B.n206 VSUBS 0.008533f
C291 B.n207 VSUBS 0.008533f
C292 B.n208 VSUBS 0.008533f
C293 B.n209 VSUBS 0.008533f
C294 B.n210 VSUBS 0.008533f
C295 B.n211 VSUBS 0.008533f
C296 B.n212 VSUBS 0.008031f
C297 B.n213 VSUBS 0.019771f
C298 B.n214 VSUBS 0.004769f
C299 B.n215 VSUBS 0.008533f
C300 B.n216 VSUBS 0.008533f
C301 B.n217 VSUBS 0.008533f
C302 B.n218 VSUBS 0.008533f
C303 B.n219 VSUBS 0.008533f
C304 B.n220 VSUBS 0.008533f
C305 B.n221 VSUBS 0.008533f
C306 B.n222 VSUBS 0.008533f
C307 B.n223 VSUBS 0.008533f
C308 B.n224 VSUBS 0.008533f
C309 B.n225 VSUBS 0.008533f
C310 B.n226 VSUBS 0.008533f
C311 B.n227 VSUBS 0.004769f
C312 B.n228 VSUBS 0.008533f
C313 B.n229 VSUBS 0.008533f
C314 B.n230 VSUBS 0.008031f
C315 B.n231 VSUBS 0.008533f
C316 B.n232 VSUBS 0.008533f
C317 B.n233 VSUBS 0.008533f
C318 B.n234 VSUBS 0.008533f
C319 B.n235 VSUBS 0.008533f
C320 B.n236 VSUBS 0.008533f
C321 B.n237 VSUBS 0.008533f
C322 B.n238 VSUBS 0.008533f
C323 B.n239 VSUBS 0.008533f
C324 B.n240 VSUBS 0.008533f
C325 B.n241 VSUBS 0.008533f
C326 B.n242 VSUBS 0.008533f
C327 B.n243 VSUBS 0.008533f
C328 B.n244 VSUBS 0.008533f
C329 B.n245 VSUBS 0.008533f
C330 B.n246 VSUBS 0.008533f
C331 B.n247 VSUBS 0.008533f
C332 B.n248 VSUBS 0.008533f
C333 B.n249 VSUBS 0.008533f
C334 B.n250 VSUBS 0.008533f
C335 B.n251 VSUBS 0.008533f
C336 B.n252 VSUBS 0.008533f
C337 B.n253 VSUBS 0.008533f
C338 B.n254 VSUBS 0.008533f
C339 B.n255 VSUBS 0.008533f
C340 B.n256 VSUBS 0.008533f
C341 B.n257 VSUBS 0.008533f
C342 B.n258 VSUBS 0.008533f
C343 B.n259 VSUBS 0.008533f
C344 B.n260 VSUBS 0.008533f
C345 B.n261 VSUBS 0.008533f
C346 B.n262 VSUBS 0.008533f
C347 B.n263 VSUBS 0.008533f
C348 B.n264 VSUBS 0.008533f
C349 B.n265 VSUBS 0.008533f
C350 B.n266 VSUBS 0.008533f
C351 B.n267 VSUBS 0.008533f
C352 B.n268 VSUBS 0.008533f
C353 B.n269 VSUBS 0.008533f
C354 B.n270 VSUBS 0.008533f
C355 B.n271 VSUBS 0.008533f
C356 B.n272 VSUBS 0.008533f
C357 B.n273 VSUBS 0.008533f
C358 B.n274 VSUBS 0.008533f
C359 B.n275 VSUBS 0.008533f
C360 B.n276 VSUBS 0.008533f
C361 B.n277 VSUBS 0.008533f
C362 B.n278 VSUBS 0.008533f
C363 B.n279 VSUBS 0.008533f
C364 B.n280 VSUBS 0.008533f
C365 B.n281 VSUBS 0.008533f
C366 B.n282 VSUBS 0.008533f
C367 B.n283 VSUBS 0.008533f
C368 B.n284 VSUBS 0.008533f
C369 B.n285 VSUBS 0.008533f
C370 B.n286 VSUBS 0.008533f
C371 B.n287 VSUBS 0.008533f
C372 B.n288 VSUBS 0.021335f
C373 B.n289 VSUBS 0.02058f
C374 B.n290 VSUBS 0.02058f
C375 B.n291 VSUBS 0.008533f
C376 B.n292 VSUBS 0.008533f
C377 B.n293 VSUBS 0.008533f
C378 B.n294 VSUBS 0.008533f
C379 B.n295 VSUBS 0.008533f
C380 B.n296 VSUBS 0.008533f
C381 B.n297 VSUBS 0.008533f
C382 B.n298 VSUBS 0.008533f
C383 B.n299 VSUBS 0.008533f
C384 B.n300 VSUBS 0.008533f
C385 B.n301 VSUBS 0.008533f
C386 B.n302 VSUBS 0.008533f
C387 B.n303 VSUBS 0.008533f
C388 B.n304 VSUBS 0.008533f
C389 B.n305 VSUBS 0.008533f
C390 B.n306 VSUBS 0.008533f
C391 B.n307 VSUBS 0.008533f
C392 B.n308 VSUBS 0.008533f
C393 B.n309 VSUBS 0.008533f
C394 B.n310 VSUBS 0.008533f
C395 B.n311 VSUBS 0.008533f
C396 B.n312 VSUBS 0.008533f
C397 B.n313 VSUBS 0.008533f
C398 B.n314 VSUBS 0.008533f
C399 B.n315 VSUBS 0.008533f
C400 B.n316 VSUBS 0.008533f
C401 B.n317 VSUBS 0.008533f
C402 B.n318 VSUBS 0.008533f
C403 B.n319 VSUBS 0.008533f
C404 B.n320 VSUBS 0.008533f
C405 B.n321 VSUBS 0.008533f
C406 B.n322 VSUBS 0.008533f
C407 B.n323 VSUBS 0.008533f
C408 B.n324 VSUBS 0.008533f
C409 B.n325 VSUBS 0.008533f
C410 B.n326 VSUBS 0.008533f
C411 B.n327 VSUBS 0.008533f
C412 B.n328 VSUBS 0.008533f
C413 B.n329 VSUBS 0.008533f
C414 B.n330 VSUBS 0.008533f
C415 B.n331 VSUBS 0.008533f
C416 B.n332 VSUBS 0.008533f
C417 B.n333 VSUBS 0.008533f
C418 B.n334 VSUBS 0.021517f
C419 B.n335 VSUBS 0.02058f
C420 B.n336 VSUBS 0.021335f
C421 B.n337 VSUBS 0.008533f
C422 B.n338 VSUBS 0.008533f
C423 B.n339 VSUBS 0.008533f
C424 B.n340 VSUBS 0.008533f
C425 B.n341 VSUBS 0.008533f
C426 B.n342 VSUBS 0.008533f
C427 B.n343 VSUBS 0.008533f
C428 B.n344 VSUBS 0.008533f
C429 B.n345 VSUBS 0.008533f
C430 B.n346 VSUBS 0.008533f
C431 B.n347 VSUBS 0.008533f
C432 B.n348 VSUBS 0.008533f
C433 B.n349 VSUBS 0.008533f
C434 B.n350 VSUBS 0.008533f
C435 B.n351 VSUBS 0.008533f
C436 B.n352 VSUBS 0.008533f
C437 B.n353 VSUBS 0.008533f
C438 B.n354 VSUBS 0.008533f
C439 B.n355 VSUBS 0.008533f
C440 B.n356 VSUBS 0.008533f
C441 B.n357 VSUBS 0.008533f
C442 B.n358 VSUBS 0.008533f
C443 B.n359 VSUBS 0.008533f
C444 B.n360 VSUBS 0.008533f
C445 B.n361 VSUBS 0.008533f
C446 B.n362 VSUBS 0.008533f
C447 B.n363 VSUBS 0.008533f
C448 B.n364 VSUBS 0.008533f
C449 B.n365 VSUBS 0.008533f
C450 B.n366 VSUBS 0.008533f
C451 B.n367 VSUBS 0.008533f
C452 B.n368 VSUBS 0.008533f
C453 B.n369 VSUBS 0.008533f
C454 B.n370 VSUBS 0.008533f
C455 B.n371 VSUBS 0.008533f
C456 B.n372 VSUBS 0.008533f
C457 B.n373 VSUBS 0.008533f
C458 B.n374 VSUBS 0.008533f
C459 B.n375 VSUBS 0.008533f
C460 B.n376 VSUBS 0.008533f
C461 B.n377 VSUBS 0.008533f
C462 B.n378 VSUBS 0.008533f
C463 B.n379 VSUBS 0.008533f
C464 B.n380 VSUBS 0.008533f
C465 B.n381 VSUBS 0.008533f
C466 B.n382 VSUBS 0.008533f
C467 B.n383 VSUBS 0.008533f
C468 B.n384 VSUBS 0.008533f
C469 B.n385 VSUBS 0.008533f
C470 B.n386 VSUBS 0.008533f
C471 B.n387 VSUBS 0.008533f
C472 B.n388 VSUBS 0.008533f
C473 B.n389 VSUBS 0.008533f
C474 B.n390 VSUBS 0.008533f
C475 B.n391 VSUBS 0.008533f
C476 B.n392 VSUBS 0.008533f
C477 B.n393 VSUBS 0.008533f
C478 B.n394 VSUBS 0.008031f
C479 B.n395 VSUBS 0.008533f
C480 B.n396 VSUBS 0.008533f
C481 B.n397 VSUBS 0.008533f
C482 B.n398 VSUBS 0.008533f
C483 B.n399 VSUBS 0.008533f
C484 B.n400 VSUBS 0.008533f
C485 B.n401 VSUBS 0.008533f
C486 B.n402 VSUBS 0.008533f
C487 B.n403 VSUBS 0.008533f
C488 B.n404 VSUBS 0.008533f
C489 B.n405 VSUBS 0.008533f
C490 B.n406 VSUBS 0.008533f
C491 B.n407 VSUBS 0.008533f
C492 B.n408 VSUBS 0.008533f
C493 B.n409 VSUBS 0.008533f
C494 B.n410 VSUBS 0.004769f
C495 B.n411 VSUBS 0.019771f
C496 B.n412 VSUBS 0.008031f
C497 B.n413 VSUBS 0.008533f
C498 B.n414 VSUBS 0.008533f
C499 B.n415 VSUBS 0.008533f
C500 B.n416 VSUBS 0.008533f
C501 B.n417 VSUBS 0.008533f
C502 B.n418 VSUBS 0.008533f
C503 B.n419 VSUBS 0.008533f
C504 B.n420 VSUBS 0.008533f
C505 B.n421 VSUBS 0.008533f
C506 B.n422 VSUBS 0.008533f
C507 B.n423 VSUBS 0.008533f
C508 B.n424 VSUBS 0.008533f
C509 B.n425 VSUBS 0.008533f
C510 B.n426 VSUBS 0.008533f
C511 B.n427 VSUBS 0.008533f
C512 B.n428 VSUBS 0.008533f
C513 B.n429 VSUBS 0.008533f
C514 B.n430 VSUBS 0.008533f
C515 B.n431 VSUBS 0.008533f
C516 B.n432 VSUBS 0.008533f
C517 B.n433 VSUBS 0.008533f
C518 B.n434 VSUBS 0.008533f
C519 B.n435 VSUBS 0.008533f
C520 B.n436 VSUBS 0.008533f
C521 B.n437 VSUBS 0.008533f
C522 B.n438 VSUBS 0.008533f
C523 B.n439 VSUBS 0.008533f
C524 B.n440 VSUBS 0.008533f
C525 B.n441 VSUBS 0.008533f
C526 B.n442 VSUBS 0.008533f
C527 B.n443 VSUBS 0.008533f
C528 B.n444 VSUBS 0.008533f
C529 B.n445 VSUBS 0.008533f
C530 B.n446 VSUBS 0.008533f
C531 B.n447 VSUBS 0.008533f
C532 B.n448 VSUBS 0.008533f
C533 B.n449 VSUBS 0.008533f
C534 B.n450 VSUBS 0.008533f
C535 B.n451 VSUBS 0.008533f
C536 B.n452 VSUBS 0.008533f
C537 B.n453 VSUBS 0.008533f
C538 B.n454 VSUBS 0.008533f
C539 B.n455 VSUBS 0.008533f
C540 B.n456 VSUBS 0.008533f
C541 B.n457 VSUBS 0.008533f
C542 B.n458 VSUBS 0.008533f
C543 B.n459 VSUBS 0.008533f
C544 B.n460 VSUBS 0.008533f
C545 B.n461 VSUBS 0.008533f
C546 B.n462 VSUBS 0.008533f
C547 B.n463 VSUBS 0.008533f
C548 B.n464 VSUBS 0.008533f
C549 B.n465 VSUBS 0.008533f
C550 B.n466 VSUBS 0.008533f
C551 B.n467 VSUBS 0.008533f
C552 B.n468 VSUBS 0.008533f
C553 B.n469 VSUBS 0.008533f
C554 B.n470 VSUBS 0.021335f
C555 B.n471 VSUBS 0.021335f
C556 B.n472 VSUBS 0.02058f
C557 B.n473 VSUBS 0.008533f
C558 B.n474 VSUBS 0.008533f
C559 B.n475 VSUBS 0.008533f
C560 B.n476 VSUBS 0.008533f
C561 B.n477 VSUBS 0.008533f
C562 B.n478 VSUBS 0.008533f
C563 B.n479 VSUBS 0.008533f
C564 B.n480 VSUBS 0.008533f
C565 B.n481 VSUBS 0.008533f
C566 B.n482 VSUBS 0.008533f
C567 B.n483 VSUBS 0.008533f
C568 B.n484 VSUBS 0.008533f
C569 B.n485 VSUBS 0.008533f
C570 B.n486 VSUBS 0.008533f
C571 B.n487 VSUBS 0.008533f
C572 B.n488 VSUBS 0.008533f
C573 B.n489 VSUBS 0.008533f
C574 B.n490 VSUBS 0.008533f
C575 B.n491 VSUBS 0.008533f
C576 B.n492 VSUBS 0.008533f
C577 B.n493 VSUBS 0.008533f
C578 B.n494 VSUBS 0.008533f
C579 B.n495 VSUBS 0.019323f
.ends

