* NGSPICE file created from diff_pair_sample_0558.ext - technology: sky130A

.subckt diff_pair_sample_0558 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=6.1815 pd=32.48 as=0 ps=0 w=15.85 l=2.27
X1 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=6.1815 pd=32.48 as=0 ps=0 w=15.85 l=2.27
X2 VTAIL.t19 VN.t0 VDD2.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.61525 pd=16.18 as=2.61525 ps=16.18 w=15.85 l=2.27
X3 VTAIL.t18 VN.t1 VDD2.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=2.61525 pd=16.18 as=2.61525 ps=16.18 w=15.85 l=2.27
X4 VDD1.t9 VP.t0 VTAIL.t7 B.t8 sky130_fd_pr__nfet_01v8 ad=2.61525 pd=16.18 as=2.61525 ps=16.18 w=15.85 l=2.27
X5 VDD2.t1 VN.t2 VTAIL.t17 B.t2 sky130_fd_pr__nfet_01v8 ad=2.61525 pd=16.18 as=6.1815 ps=32.48 w=15.85 l=2.27
X6 VDD2.t2 VN.t3 VTAIL.t16 B.t3 sky130_fd_pr__nfet_01v8 ad=2.61525 pd=16.18 as=2.61525 ps=16.18 w=15.85 l=2.27
X7 VDD1.t8 VP.t1 VTAIL.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=2.61525 pd=16.18 as=6.1815 ps=32.48 w=15.85 l=2.27
X8 VTAIL.t5 VP.t2 VDD1.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.61525 pd=16.18 as=2.61525 ps=16.18 w=15.85 l=2.27
X9 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=6.1815 pd=32.48 as=0 ps=0 w=15.85 l=2.27
X10 VTAIL.t15 VN.t4 VDD2.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=2.61525 pd=16.18 as=2.61525 ps=16.18 w=15.85 l=2.27
X11 VDD2.t8 VN.t5 VTAIL.t14 B.t9 sky130_fd_pr__nfet_01v8 ad=2.61525 pd=16.18 as=6.1815 ps=32.48 w=15.85 l=2.27
X12 VDD1.t6 VP.t3 VTAIL.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=6.1815 pd=32.48 as=2.61525 ps=16.18 w=15.85 l=2.27
X13 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.1815 pd=32.48 as=0 ps=0 w=15.85 l=2.27
X14 VDD1.t5 VP.t4 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=2.61525 pd=16.18 as=6.1815 ps=32.48 w=15.85 l=2.27
X15 VTAIL.t1 VP.t5 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.61525 pd=16.18 as=2.61525 ps=16.18 w=15.85 l=2.27
X16 VDD2.t5 VN.t6 VTAIL.t13 B.t8 sky130_fd_pr__nfet_01v8 ad=2.61525 pd=16.18 as=2.61525 ps=16.18 w=15.85 l=2.27
X17 VDD2.t4 VN.t7 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=6.1815 pd=32.48 as=2.61525 ps=16.18 w=15.85 l=2.27
X18 VTAIL.t8 VP.t6 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=2.61525 pd=16.18 as=2.61525 ps=16.18 w=15.85 l=2.27
X19 VDD1.t2 VP.t7 VTAIL.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=6.1815 pd=32.48 as=2.61525 ps=16.18 w=15.85 l=2.27
X20 VDD2.t3 VN.t8 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=6.1815 pd=32.48 as=2.61525 ps=16.18 w=15.85 l=2.27
X21 VDD1.t1 VP.t8 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.61525 pd=16.18 as=2.61525 ps=16.18 w=15.85 l=2.27
X22 VTAIL.t0 VP.t9 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.61525 pd=16.18 as=2.61525 ps=16.18 w=15.85 l=2.27
X23 VTAIL.t10 VN.t9 VDD2.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.61525 pd=16.18 as=2.61525 ps=16.18 w=15.85 l=2.27
R0 B.n792 B.n162 585
R1 B.n162 B.n99 585
R2 B.n794 B.n793 585
R3 B.n796 B.n161 585
R4 B.n799 B.n798 585
R5 B.n800 B.n160 585
R6 B.n802 B.n801 585
R7 B.n804 B.n159 585
R8 B.n807 B.n806 585
R9 B.n808 B.n158 585
R10 B.n810 B.n809 585
R11 B.n812 B.n157 585
R12 B.n815 B.n814 585
R13 B.n816 B.n156 585
R14 B.n818 B.n817 585
R15 B.n820 B.n155 585
R16 B.n823 B.n822 585
R17 B.n824 B.n154 585
R18 B.n826 B.n825 585
R19 B.n828 B.n153 585
R20 B.n831 B.n830 585
R21 B.n832 B.n152 585
R22 B.n834 B.n833 585
R23 B.n836 B.n151 585
R24 B.n839 B.n838 585
R25 B.n840 B.n150 585
R26 B.n842 B.n841 585
R27 B.n844 B.n149 585
R28 B.n847 B.n846 585
R29 B.n848 B.n148 585
R30 B.n850 B.n849 585
R31 B.n852 B.n147 585
R32 B.n855 B.n854 585
R33 B.n856 B.n146 585
R34 B.n858 B.n857 585
R35 B.n860 B.n145 585
R36 B.n863 B.n862 585
R37 B.n864 B.n144 585
R38 B.n866 B.n865 585
R39 B.n868 B.n143 585
R40 B.n871 B.n870 585
R41 B.n872 B.n142 585
R42 B.n874 B.n873 585
R43 B.n876 B.n141 585
R44 B.n879 B.n878 585
R45 B.n880 B.n140 585
R46 B.n882 B.n881 585
R47 B.n884 B.n139 585
R48 B.n887 B.n886 585
R49 B.n888 B.n138 585
R50 B.n890 B.n889 585
R51 B.n892 B.n137 585
R52 B.n894 B.n893 585
R53 B.n896 B.n895 585
R54 B.n899 B.n898 585
R55 B.n900 B.n132 585
R56 B.n902 B.n901 585
R57 B.n904 B.n131 585
R58 B.n907 B.n906 585
R59 B.n908 B.n130 585
R60 B.n910 B.n909 585
R61 B.n912 B.n129 585
R62 B.n915 B.n914 585
R63 B.n917 B.n126 585
R64 B.n919 B.n918 585
R65 B.n921 B.n125 585
R66 B.n924 B.n923 585
R67 B.n925 B.n124 585
R68 B.n927 B.n926 585
R69 B.n929 B.n123 585
R70 B.n932 B.n931 585
R71 B.n933 B.n122 585
R72 B.n935 B.n934 585
R73 B.n937 B.n121 585
R74 B.n940 B.n939 585
R75 B.n941 B.n120 585
R76 B.n943 B.n942 585
R77 B.n945 B.n119 585
R78 B.n948 B.n947 585
R79 B.n949 B.n118 585
R80 B.n951 B.n950 585
R81 B.n953 B.n117 585
R82 B.n956 B.n955 585
R83 B.n957 B.n116 585
R84 B.n959 B.n958 585
R85 B.n961 B.n115 585
R86 B.n964 B.n963 585
R87 B.n965 B.n114 585
R88 B.n967 B.n966 585
R89 B.n969 B.n113 585
R90 B.n972 B.n971 585
R91 B.n973 B.n112 585
R92 B.n975 B.n974 585
R93 B.n977 B.n111 585
R94 B.n980 B.n979 585
R95 B.n981 B.n110 585
R96 B.n983 B.n982 585
R97 B.n985 B.n109 585
R98 B.n988 B.n987 585
R99 B.n989 B.n108 585
R100 B.n991 B.n990 585
R101 B.n993 B.n107 585
R102 B.n996 B.n995 585
R103 B.n997 B.n106 585
R104 B.n999 B.n998 585
R105 B.n1001 B.n105 585
R106 B.n1004 B.n1003 585
R107 B.n1005 B.n104 585
R108 B.n1007 B.n1006 585
R109 B.n1009 B.n103 585
R110 B.n1012 B.n1011 585
R111 B.n1013 B.n102 585
R112 B.n1015 B.n1014 585
R113 B.n1017 B.n101 585
R114 B.n1020 B.n1019 585
R115 B.n1021 B.n100 585
R116 B.n791 B.n98 585
R117 B.n1024 B.n98 585
R118 B.n790 B.n97 585
R119 B.n1025 B.n97 585
R120 B.n789 B.n96 585
R121 B.n1026 B.n96 585
R122 B.n788 B.n787 585
R123 B.n787 B.n92 585
R124 B.n786 B.n91 585
R125 B.n1032 B.n91 585
R126 B.n785 B.n90 585
R127 B.n1033 B.n90 585
R128 B.n784 B.n89 585
R129 B.n1034 B.n89 585
R130 B.n783 B.n782 585
R131 B.n782 B.n88 585
R132 B.n781 B.n84 585
R133 B.n1040 B.n84 585
R134 B.n780 B.n83 585
R135 B.n1041 B.n83 585
R136 B.n779 B.n82 585
R137 B.n1042 B.n82 585
R138 B.n778 B.n777 585
R139 B.n777 B.n78 585
R140 B.n776 B.n77 585
R141 B.n1048 B.n77 585
R142 B.n775 B.n76 585
R143 B.n1049 B.n76 585
R144 B.n774 B.n75 585
R145 B.n1050 B.n75 585
R146 B.n773 B.n772 585
R147 B.n772 B.n71 585
R148 B.n771 B.n70 585
R149 B.n1056 B.n70 585
R150 B.n770 B.n69 585
R151 B.n1057 B.n69 585
R152 B.n769 B.n68 585
R153 B.n1058 B.n68 585
R154 B.n768 B.n767 585
R155 B.n767 B.n64 585
R156 B.n766 B.n63 585
R157 B.n1064 B.n63 585
R158 B.n765 B.n62 585
R159 B.n1065 B.n62 585
R160 B.n764 B.n61 585
R161 B.n1066 B.n61 585
R162 B.n763 B.n762 585
R163 B.n762 B.n57 585
R164 B.n761 B.n56 585
R165 B.n1072 B.n56 585
R166 B.n760 B.n55 585
R167 B.n1073 B.n55 585
R168 B.n759 B.n54 585
R169 B.n1074 B.n54 585
R170 B.n758 B.n757 585
R171 B.n757 B.n50 585
R172 B.n756 B.n49 585
R173 B.n1080 B.n49 585
R174 B.n755 B.n48 585
R175 B.n1081 B.n48 585
R176 B.n754 B.n47 585
R177 B.n1082 B.n47 585
R178 B.n753 B.n752 585
R179 B.n752 B.n43 585
R180 B.n751 B.n42 585
R181 B.n1088 B.n42 585
R182 B.n750 B.n41 585
R183 B.n1089 B.n41 585
R184 B.n749 B.n40 585
R185 B.n1090 B.n40 585
R186 B.n748 B.n747 585
R187 B.n747 B.n36 585
R188 B.n746 B.n35 585
R189 B.n1096 B.n35 585
R190 B.n745 B.n34 585
R191 B.n1097 B.n34 585
R192 B.n744 B.n33 585
R193 B.n1098 B.n33 585
R194 B.n743 B.n742 585
R195 B.n742 B.n29 585
R196 B.n741 B.n28 585
R197 B.n1104 B.n28 585
R198 B.n740 B.n27 585
R199 B.n1105 B.n27 585
R200 B.n739 B.n26 585
R201 B.n1106 B.n26 585
R202 B.n738 B.n737 585
R203 B.n737 B.n22 585
R204 B.n736 B.n21 585
R205 B.n1112 B.n21 585
R206 B.n735 B.n20 585
R207 B.n1113 B.n20 585
R208 B.n734 B.n19 585
R209 B.n1114 B.n19 585
R210 B.n733 B.n732 585
R211 B.n732 B.n15 585
R212 B.n731 B.n14 585
R213 B.n1120 B.n14 585
R214 B.n730 B.n13 585
R215 B.n1121 B.n13 585
R216 B.n729 B.n12 585
R217 B.n1122 B.n12 585
R218 B.n728 B.n727 585
R219 B.n727 B.n8 585
R220 B.n726 B.n7 585
R221 B.n1128 B.n7 585
R222 B.n725 B.n6 585
R223 B.n1129 B.n6 585
R224 B.n724 B.n5 585
R225 B.n1130 B.n5 585
R226 B.n723 B.n722 585
R227 B.n722 B.n4 585
R228 B.n721 B.n163 585
R229 B.n721 B.n720 585
R230 B.n711 B.n164 585
R231 B.n165 B.n164 585
R232 B.n713 B.n712 585
R233 B.n714 B.n713 585
R234 B.n710 B.n170 585
R235 B.n170 B.n169 585
R236 B.n709 B.n708 585
R237 B.n708 B.n707 585
R238 B.n172 B.n171 585
R239 B.n173 B.n172 585
R240 B.n700 B.n699 585
R241 B.n701 B.n700 585
R242 B.n698 B.n178 585
R243 B.n178 B.n177 585
R244 B.n697 B.n696 585
R245 B.n696 B.n695 585
R246 B.n180 B.n179 585
R247 B.n181 B.n180 585
R248 B.n688 B.n687 585
R249 B.n689 B.n688 585
R250 B.n686 B.n186 585
R251 B.n186 B.n185 585
R252 B.n685 B.n684 585
R253 B.n684 B.n683 585
R254 B.n188 B.n187 585
R255 B.n189 B.n188 585
R256 B.n676 B.n675 585
R257 B.n677 B.n676 585
R258 B.n674 B.n194 585
R259 B.n194 B.n193 585
R260 B.n673 B.n672 585
R261 B.n672 B.n671 585
R262 B.n196 B.n195 585
R263 B.n197 B.n196 585
R264 B.n664 B.n663 585
R265 B.n665 B.n664 585
R266 B.n662 B.n201 585
R267 B.n205 B.n201 585
R268 B.n661 B.n660 585
R269 B.n660 B.n659 585
R270 B.n203 B.n202 585
R271 B.n204 B.n203 585
R272 B.n652 B.n651 585
R273 B.n653 B.n652 585
R274 B.n650 B.n210 585
R275 B.n210 B.n209 585
R276 B.n649 B.n648 585
R277 B.n648 B.n647 585
R278 B.n212 B.n211 585
R279 B.n213 B.n212 585
R280 B.n640 B.n639 585
R281 B.n641 B.n640 585
R282 B.n638 B.n217 585
R283 B.n221 B.n217 585
R284 B.n637 B.n636 585
R285 B.n636 B.n635 585
R286 B.n219 B.n218 585
R287 B.n220 B.n219 585
R288 B.n628 B.n627 585
R289 B.n629 B.n628 585
R290 B.n626 B.n226 585
R291 B.n226 B.n225 585
R292 B.n625 B.n624 585
R293 B.n624 B.n623 585
R294 B.n228 B.n227 585
R295 B.n229 B.n228 585
R296 B.n616 B.n615 585
R297 B.n617 B.n616 585
R298 B.n614 B.n233 585
R299 B.n237 B.n233 585
R300 B.n613 B.n612 585
R301 B.n612 B.n611 585
R302 B.n235 B.n234 585
R303 B.n236 B.n235 585
R304 B.n604 B.n603 585
R305 B.n605 B.n604 585
R306 B.n602 B.n242 585
R307 B.n242 B.n241 585
R308 B.n601 B.n600 585
R309 B.n600 B.n599 585
R310 B.n244 B.n243 585
R311 B.n245 B.n244 585
R312 B.n592 B.n591 585
R313 B.n593 B.n592 585
R314 B.n590 B.n250 585
R315 B.n250 B.n249 585
R316 B.n589 B.n588 585
R317 B.n588 B.n587 585
R318 B.n252 B.n251 585
R319 B.n580 B.n252 585
R320 B.n579 B.n578 585
R321 B.n581 B.n579 585
R322 B.n577 B.n257 585
R323 B.n257 B.n256 585
R324 B.n576 B.n575 585
R325 B.n575 B.n574 585
R326 B.n259 B.n258 585
R327 B.n260 B.n259 585
R328 B.n567 B.n566 585
R329 B.n568 B.n567 585
R330 B.n565 B.n265 585
R331 B.n265 B.n264 585
R332 B.n564 B.n563 585
R333 B.n563 B.n562 585
R334 B.n559 B.n269 585
R335 B.n558 B.n557 585
R336 B.n555 B.n270 585
R337 B.n555 B.n268 585
R338 B.n554 B.n553 585
R339 B.n552 B.n551 585
R340 B.n550 B.n272 585
R341 B.n548 B.n547 585
R342 B.n546 B.n273 585
R343 B.n545 B.n544 585
R344 B.n542 B.n274 585
R345 B.n540 B.n539 585
R346 B.n538 B.n275 585
R347 B.n537 B.n536 585
R348 B.n534 B.n276 585
R349 B.n532 B.n531 585
R350 B.n530 B.n277 585
R351 B.n529 B.n528 585
R352 B.n526 B.n278 585
R353 B.n524 B.n523 585
R354 B.n522 B.n279 585
R355 B.n521 B.n520 585
R356 B.n518 B.n280 585
R357 B.n516 B.n515 585
R358 B.n514 B.n281 585
R359 B.n513 B.n512 585
R360 B.n510 B.n282 585
R361 B.n508 B.n507 585
R362 B.n506 B.n283 585
R363 B.n505 B.n504 585
R364 B.n502 B.n284 585
R365 B.n500 B.n499 585
R366 B.n498 B.n285 585
R367 B.n497 B.n496 585
R368 B.n494 B.n286 585
R369 B.n492 B.n491 585
R370 B.n490 B.n287 585
R371 B.n489 B.n488 585
R372 B.n486 B.n288 585
R373 B.n484 B.n483 585
R374 B.n482 B.n289 585
R375 B.n481 B.n480 585
R376 B.n478 B.n290 585
R377 B.n476 B.n475 585
R378 B.n474 B.n291 585
R379 B.n473 B.n472 585
R380 B.n470 B.n292 585
R381 B.n468 B.n467 585
R382 B.n466 B.n293 585
R383 B.n465 B.n464 585
R384 B.n462 B.n294 585
R385 B.n460 B.n459 585
R386 B.n458 B.n295 585
R387 B.n457 B.n456 585
R388 B.n454 B.n453 585
R389 B.n452 B.n451 585
R390 B.n450 B.n300 585
R391 B.n448 B.n447 585
R392 B.n446 B.n301 585
R393 B.n445 B.n444 585
R394 B.n442 B.n302 585
R395 B.n440 B.n439 585
R396 B.n438 B.n303 585
R397 B.n436 B.n435 585
R398 B.n433 B.n306 585
R399 B.n431 B.n430 585
R400 B.n429 B.n307 585
R401 B.n428 B.n427 585
R402 B.n425 B.n308 585
R403 B.n423 B.n422 585
R404 B.n421 B.n309 585
R405 B.n420 B.n419 585
R406 B.n417 B.n310 585
R407 B.n415 B.n414 585
R408 B.n413 B.n311 585
R409 B.n412 B.n411 585
R410 B.n409 B.n312 585
R411 B.n407 B.n406 585
R412 B.n405 B.n313 585
R413 B.n404 B.n403 585
R414 B.n401 B.n314 585
R415 B.n399 B.n398 585
R416 B.n397 B.n315 585
R417 B.n396 B.n395 585
R418 B.n393 B.n316 585
R419 B.n391 B.n390 585
R420 B.n389 B.n317 585
R421 B.n388 B.n387 585
R422 B.n385 B.n318 585
R423 B.n383 B.n382 585
R424 B.n381 B.n319 585
R425 B.n380 B.n379 585
R426 B.n377 B.n320 585
R427 B.n375 B.n374 585
R428 B.n373 B.n321 585
R429 B.n372 B.n371 585
R430 B.n369 B.n322 585
R431 B.n367 B.n366 585
R432 B.n365 B.n323 585
R433 B.n364 B.n363 585
R434 B.n361 B.n324 585
R435 B.n359 B.n358 585
R436 B.n357 B.n325 585
R437 B.n356 B.n355 585
R438 B.n353 B.n326 585
R439 B.n351 B.n350 585
R440 B.n349 B.n327 585
R441 B.n348 B.n347 585
R442 B.n345 B.n328 585
R443 B.n343 B.n342 585
R444 B.n341 B.n329 585
R445 B.n340 B.n339 585
R446 B.n337 B.n330 585
R447 B.n335 B.n334 585
R448 B.n333 B.n332 585
R449 B.n267 B.n266 585
R450 B.n561 B.n560 585
R451 B.n562 B.n561 585
R452 B.n263 B.n262 585
R453 B.n264 B.n263 585
R454 B.n570 B.n569 585
R455 B.n569 B.n568 585
R456 B.n571 B.n261 585
R457 B.n261 B.n260 585
R458 B.n573 B.n572 585
R459 B.n574 B.n573 585
R460 B.n255 B.n254 585
R461 B.n256 B.n255 585
R462 B.n583 B.n582 585
R463 B.n582 B.n581 585
R464 B.n584 B.n253 585
R465 B.n580 B.n253 585
R466 B.n586 B.n585 585
R467 B.n587 B.n586 585
R468 B.n248 B.n247 585
R469 B.n249 B.n248 585
R470 B.n595 B.n594 585
R471 B.n594 B.n593 585
R472 B.n596 B.n246 585
R473 B.n246 B.n245 585
R474 B.n598 B.n597 585
R475 B.n599 B.n598 585
R476 B.n240 B.n239 585
R477 B.n241 B.n240 585
R478 B.n607 B.n606 585
R479 B.n606 B.n605 585
R480 B.n608 B.n238 585
R481 B.n238 B.n236 585
R482 B.n610 B.n609 585
R483 B.n611 B.n610 585
R484 B.n232 B.n231 585
R485 B.n237 B.n232 585
R486 B.n619 B.n618 585
R487 B.n618 B.n617 585
R488 B.n620 B.n230 585
R489 B.n230 B.n229 585
R490 B.n622 B.n621 585
R491 B.n623 B.n622 585
R492 B.n224 B.n223 585
R493 B.n225 B.n224 585
R494 B.n631 B.n630 585
R495 B.n630 B.n629 585
R496 B.n632 B.n222 585
R497 B.n222 B.n220 585
R498 B.n634 B.n633 585
R499 B.n635 B.n634 585
R500 B.n216 B.n215 585
R501 B.n221 B.n216 585
R502 B.n643 B.n642 585
R503 B.n642 B.n641 585
R504 B.n644 B.n214 585
R505 B.n214 B.n213 585
R506 B.n646 B.n645 585
R507 B.n647 B.n646 585
R508 B.n208 B.n207 585
R509 B.n209 B.n208 585
R510 B.n655 B.n654 585
R511 B.n654 B.n653 585
R512 B.n656 B.n206 585
R513 B.n206 B.n204 585
R514 B.n658 B.n657 585
R515 B.n659 B.n658 585
R516 B.n200 B.n199 585
R517 B.n205 B.n200 585
R518 B.n667 B.n666 585
R519 B.n666 B.n665 585
R520 B.n668 B.n198 585
R521 B.n198 B.n197 585
R522 B.n670 B.n669 585
R523 B.n671 B.n670 585
R524 B.n192 B.n191 585
R525 B.n193 B.n192 585
R526 B.n679 B.n678 585
R527 B.n678 B.n677 585
R528 B.n680 B.n190 585
R529 B.n190 B.n189 585
R530 B.n682 B.n681 585
R531 B.n683 B.n682 585
R532 B.n184 B.n183 585
R533 B.n185 B.n184 585
R534 B.n691 B.n690 585
R535 B.n690 B.n689 585
R536 B.n692 B.n182 585
R537 B.n182 B.n181 585
R538 B.n694 B.n693 585
R539 B.n695 B.n694 585
R540 B.n176 B.n175 585
R541 B.n177 B.n176 585
R542 B.n703 B.n702 585
R543 B.n702 B.n701 585
R544 B.n704 B.n174 585
R545 B.n174 B.n173 585
R546 B.n706 B.n705 585
R547 B.n707 B.n706 585
R548 B.n168 B.n167 585
R549 B.n169 B.n168 585
R550 B.n716 B.n715 585
R551 B.n715 B.n714 585
R552 B.n717 B.n166 585
R553 B.n166 B.n165 585
R554 B.n719 B.n718 585
R555 B.n720 B.n719 585
R556 B.n2 B.n0 585
R557 B.n4 B.n2 585
R558 B.n3 B.n1 585
R559 B.n1129 B.n3 585
R560 B.n1127 B.n1126 585
R561 B.n1128 B.n1127 585
R562 B.n1125 B.n9 585
R563 B.n9 B.n8 585
R564 B.n1124 B.n1123 585
R565 B.n1123 B.n1122 585
R566 B.n11 B.n10 585
R567 B.n1121 B.n11 585
R568 B.n1119 B.n1118 585
R569 B.n1120 B.n1119 585
R570 B.n1117 B.n16 585
R571 B.n16 B.n15 585
R572 B.n1116 B.n1115 585
R573 B.n1115 B.n1114 585
R574 B.n18 B.n17 585
R575 B.n1113 B.n18 585
R576 B.n1111 B.n1110 585
R577 B.n1112 B.n1111 585
R578 B.n1109 B.n23 585
R579 B.n23 B.n22 585
R580 B.n1108 B.n1107 585
R581 B.n1107 B.n1106 585
R582 B.n25 B.n24 585
R583 B.n1105 B.n25 585
R584 B.n1103 B.n1102 585
R585 B.n1104 B.n1103 585
R586 B.n1101 B.n30 585
R587 B.n30 B.n29 585
R588 B.n1100 B.n1099 585
R589 B.n1099 B.n1098 585
R590 B.n32 B.n31 585
R591 B.n1097 B.n32 585
R592 B.n1095 B.n1094 585
R593 B.n1096 B.n1095 585
R594 B.n1093 B.n37 585
R595 B.n37 B.n36 585
R596 B.n1092 B.n1091 585
R597 B.n1091 B.n1090 585
R598 B.n39 B.n38 585
R599 B.n1089 B.n39 585
R600 B.n1087 B.n1086 585
R601 B.n1088 B.n1087 585
R602 B.n1085 B.n44 585
R603 B.n44 B.n43 585
R604 B.n1084 B.n1083 585
R605 B.n1083 B.n1082 585
R606 B.n46 B.n45 585
R607 B.n1081 B.n46 585
R608 B.n1079 B.n1078 585
R609 B.n1080 B.n1079 585
R610 B.n1077 B.n51 585
R611 B.n51 B.n50 585
R612 B.n1076 B.n1075 585
R613 B.n1075 B.n1074 585
R614 B.n53 B.n52 585
R615 B.n1073 B.n53 585
R616 B.n1071 B.n1070 585
R617 B.n1072 B.n1071 585
R618 B.n1069 B.n58 585
R619 B.n58 B.n57 585
R620 B.n1068 B.n1067 585
R621 B.n1067 B.n1066 585
R622 B.n60 B.n59 585
R623 B.n1065 B.n60 585
R624 B.n1063 B.n1062 585
R625 B.n1064 B.n1063 585
R626 B.n1061 B.n65 585
R627 B.n65 B.n64 585
R628 B.n1060 B.n1059 585
R629 B.n1059 B.n1058 585
R630 B.n67 B.n66 585
R631 B.n1057 B.n67 585
R632 B.n1055 B.n1054 585
R633 B.n1056 B.n1055 585
R634 B.n1053 B.n72 585
R635 B.n72 B.n71 585
R636 B.n1052 B.n1051 585
R637 B.n1051 B.n1050 585
R638 B.n74 B.n73 585
R639 B.n1049 B.n74 585
R640 B.n1047 B.n1046 585
R641 B.n1048 B.n1047 585
R642 B.n1045 B.n79 585
R643 B.n79 B.n78 585
R644 B.n1044 B.n1043 585
R645 B.n1043 B.n1042 585
R646 B.n81 B.n80 585
R647 B.n1041 B.n81 585
R648 B.n1039 B.n1038 585
R649 B.n1040 B.n1039 585
R650 B.n1037 B.n85 585
R651 B.n88 B.n85 585
R652 B.n1036 B.n1035 585
R653 B.n1035 B.n1034 585
R654 B.n87 B.n86 585
R655 B.n1033 B.n87 585
R656 B.n1031 B.n1030 585
R657 B.n1032 B.n1031 585
R658 B.n1029 B.n93 585
R659 B.n93 B.n92 585
R660 B.n1028 B.n1027 585
R661 B.n1027 B.n1026 585
R662 B.n95 B.n94 585
R663 B.n1025 B.n95 585
R664 B.n1023 B.n1022 585
R665 B.n1024 B.n1023 585
R666 B.n1132 B.n1131 585
R667 B.n1131 B.n1130 585
R668 B.n561 B.n269 535.745
R669 B.n1023 B.n100 535.745
R670 B.n563 B.n267 535.745
R671 B.n162 B.n98 535.745
R672 B.n304 B.t10 375.764
R673 B.n296 B.t18 375.764
R674 B.n127 B.t21 375.764
R675 B.n133 B.t14 375.764
R676 B.n795 B.n99 256.663
R677 B.n797 B.n99 256.663
R678 B.n803 B.n99 256.663
R679 B.n805 B.n99 256.663
R680 B.n811 B.n99 256.663
R681 B.n813 B.n99 256.663
R682 B.n819 B.n99 256.663
R683 B.n821 B.n99 256.663
R684 B.n827 B.n99 256.663
R685 B.n829 B.n99 256.663
R686 B.n835 B.n99 256.663
R687 B.n837 B.n99 256.663
R688 B.n843 B.n99 256.663
R689 B.n845 B.n99 256.663
R690 B.n851 B.n99 256.663
R691 B.n853 B.n99 256.663
R692 B.n859 B.n99 256.663
R693 B.n861 B.n99 256.663
R694 B.n867 B.n99 256.663
R695 B.n869 B.n99 256.663
R696 B.n875 B.n99 256.663
R697 B.n877 B.n99 256.663
R698 B.n883 B.n99 256.663
R699 B.n885 B.n99 256.663
R700 B.n891 B.n99 256.663
R701 B.n136 B.n99 256.663
R702 B.n897 B.n99 256.663
R703 B.n903 B.n99 256.663
R704 B.n905 B.n99 256.663
R705 B.n911 B.n99 256.663
R706 B.n913 B.n99 256.663
R707 B.n920 B.n99 256.663
R708 B.n922 B.n99 256.663
R709 B.n928 B.n99 256.663
R710 B.n930 B.n99 256.663
R711 B.n936 B.n99 256.663
R712 B.n938 B.n99 256.663
R713 B.n944 B.n99 256.663
R714 B.n946 B.n99 256.663
R715 B.n952 B.n99 256.663
R716 B.n954 B.n99 256.663
R717 B.n960 B.n99 256.663
R718 B.n962 B.n99 256.663
R719 B.n968 B.n99 256.663
R720 B.n970 B.n99 256.663
R721 B.n976 B.n99 256.663
R722 B.n978 B.n99 256.663
R723 B.n984 B.n99 256.663
R724 B.n986 B.n99 256.663
R725 B.n992 B.n99 256.663
R726 B.n994 B.n99 256.663
R727 B.n1000 B.n99 256.663
R728 B.n1002 B.n99 256.663
R729 B.n1008 B.n99 256.663
R730 B.n1010 B.n99 256.663
R731 B.n1016 B.n99 256.663
R732 B.n1018 B.n99 256.663
R733 B.n556 B.n268 256.663
R734 B.n271 B.n268 256.663
R735 B.n549 B.n268 256.663
R736 B.n543 B.n268 256.663
R737 B.n541 B.n268 256.663
R738 B.n535 B.n268 256.663
R739 B.n533 B.n268 256.663
R740 B.n527 B.n268 256.663
R741 B.n525 B.n268 256.663
R742 B.n519 B.n268 256.663
R743 B.n517 B.n268 256.663
R744 B.n511 B.n268 256.663
R745 B.n509 B.n268 256.663
R746 B.n503 B.n268 256.663
R747 B.n501 B.n268 256.663
R748 B.n495 B.n268 256.663
R749 B.n493 B.n268 256.663
R750 B.n487 B.n268 256.663
R751 B.n485 B.n268 256.663
R752 B.n479 B.n268 256.663
R753 B.n477 B.n268 256.663
R754 B.n471 B.n268 256.663
R755 B.n469 B.n268 256.663
R756 B.n463 B.n268 256.663
R757 B.n461 B.n268 256.663
R758 B.n455 B.n268 256.663
R759 B.n299 B.n268 256.663
R760 B.n449 B.n268 256.663
R761 B.n443 B.n268 256.663
R762 B.n441 B.n268 256.663
R763 B.n434 B.n268 256.663
R764 B.n432 B.n268 256.663
R765 B.n426 B.n268 256.663
R766 B.n424 B.n268 256.663
R767 B.n418 B.n268 256.663
R768 B.n416 B.n268 256.663
R769 B.n410 B.n268 256.663
R770 B.n408 B.n268 256.663
R771 B.n402 B.n268 256.663
R772 B.n400 B.n268 256.663
R773 B.n394 B.n268 256.663
R774 B.n392 B.n268 256.663
R775 B.n386 B.n268 256.663
R776 B.n384 B.n268 256.663
R777 B.n378 B.n268 256.663
R778 B.n376 B.n268 256.663
R779 B.n370 B.n268 256.663
R780 B.n368 B.n268 256.663
R781 B.n362 B.n268 256.663
R782 B.n360 B.n268 256.663
R783 B.n354 B.n268 256.663
R784 B.n352 B.n268 256.663
R785 B.n346 B.n268 256.663
R786 B.n344 B.n268 256.663
R787 B.n338 B.n268 256.663
R788 B.n336 B.n268 256.663
R789 B.n331 B.n268 256.663
R790 B.n561 B.n263 163.367
R791 B.n569 B.n263 163.367
R792 B.n569 B.n261 163.367
R793 B.n573 B.n261 163.367
R794 B.n573 B.n255 163.367
R795 B.n582 B.n255 163.367
R796 B.n582 B.n253 163.367
R797 B.n586 B.n253 163.367
R798 B.n586 B.n248 163.367
R799 B.n594 B.n248 163.367
R800 B.n594 B.n246 163.367
R801 B.n598 B.n246 163.367
R802 B.n598 B.n240 163.367
R803 B.n606 B.n240 163.367
R804 B.n606 B.n238 163.367
R805 B.n610 B.n238 163.367
R806 B.n610 B.n232 163.367
R807 B.n618 B.n232 163.367
R808 B.n618 B.n230 163.367
R809 B.n622 B.n230 163.367
R810 B.n622 B.n224 163.367
R811 B.n630 B.n224 163.367
R812 B.n630 B.n222 163.367
R813 B.n634 B.n222 163.367
R814 B.n634 B.n216 163.367
R815 B.n642 B.n216 163.367
R816 B.n642 B.n214 163.367
R817 B.n646 B.n214 163.367
R818 B.n646 B.n208 163.367
R819 B.n654 B.n208 163.367
R820 B.n654 B.n206 163.367
R821 B.n658 B.n206 163.367
R822 B.n658 B.n200 163.367
R823 B.n666 B.n200 163.367
R824 B.n666 B.n198 163.367
R825 B.n670 B.n198 163.367
R826 B.n670 B.n192 163.367
R827 B.n678 B.n192 163.367
R828 B.n678 B.n190 163.367
R829 B.n682 B.n190 163.367
R830 B.n682 B.n184 163.367
R831 B.n690 B.n184 163.367
R832 B.n690 B.n182 163.367
R833 B.n694 B.n182 163.367
R834 B.n694 B.n176 163.367
R835 B.n702 B.n176 163.367
R836 B.n702 B.n174 163.367
R837 B.n706 B.n174 163.367
R838 B.n706 B.n168 163.367
R839 B.n715 B.n168 163.367
R840 B.n715 B.n166 163.367
R841 B.n719 B.n166 163.367
R842 B.n719 B.n2 163.367
R843 B.n1131 B.n2 163.367
R844 B.n1131 B.n3 163.367
R845 B.n1127 B.n3 163.367
R846 B.n1127 B.n9 163.367
R847 B.n1123 B.n9 163.367
R848 B.n1123 B.n11 163.367
R849 B.n1119 B.n11 163.367
R850 B.n1119 B.n16 163.367
R851 B.n1115 B.n16 163.367
R852 B.n1115 B.n18 163.367
R853 B.n1111 B.n18 163.367
R854 B.n1111 B.n23 163.367
R855 B.n1107 B.n23 163.367
R856 B.n1107 B.n25 163.367
R857 B.n1103 B.n25 163.367
R858 B.n1103 B.n30 163.367
R859 B.n1099 B.n30 163.367
R860 B.n1099 B.n32 163.367
R861 B.n1095 B.n32 163.367
R862 B.n1095 B.n37 163.367
R863 B.n1091 B.n37 163.367
R864 B.n1091 B.n39 163.367
R865 B.n1087 B.n39 163.367
R866 B.n1087 B.n44 163.367
R867 B.n1083 B.n44 163.367
R868 B.n1083 B.n46 163.367
R869 B.n1079 B.n46 163.367
R870 B.n1079 B.n51 163.367
R871 B.n1075 B.n51 163.367
R872 B.n1075 B.n53 163.367
R873 B.n1071 B.n53 163.367
R874 B.n1071 B.n58 163.367
R875 B.n1067 B.n58 163.367
R876 B.n1067 B.n60 163.367
R877 B.n1063 B.n60 163.367
R878 B.n1063 B.n65 163.367
R879 B.n1059 B.n65 163.367
R880 B.n1059 B.n67 163.367
R881 B.n1055 B.n67 163.367
R882 B.n1055 B.n72 163.367
R883 B.n1051 B.n72 163.367
R884 B.n1051 B.n74 163.367
R885 B.n1047 B.n74 163.367
R886 B.n1047 B.n79 163.367
R887 B.n1043 B.n79 163.367
R888 B.n1043 B.n81 163.367
R889 B.n1039 B.n81 163.367
R890 B.n1039 B.n85 163.367
R891 B.n1035 B.n85 163.367
R892 B.n1035 B.n87 163.367
R893 B.n1031 B.n87 163.367
R894 B.n1031 B.n93 163.367
R895 B.n1027 B.n93 163.367
R896 B.n1027 B.n95 163.367
R897 B.n1023 B.n95 163.367
R898 B.n557 B.n555 163.367
R899 B.n555 B.n554 163.367
R900 B.n551 B.n550 163.367
R901 B.n548 B.n273 163.367
R902 B.n544 B.n542 163.367
R903 B.n540 B.n275 163.367
R904 B.n536 B.n534 163.367
R905 B.n532 B.n277 163.367
R906 B.n528 B.n526 163.367
R907 B.n524 B.n279 163.367
R908 B.n520 B.n518 163.367
R909 B.n516 B.n281 163.367
R910 B.n512 B.n510 163.367
R911 B.n508 B.n283 163.367
R912 B.n504 B.n502 163.367
R913 B.n500 B.n285 163.367
R914 B.n496 B.n494 163.367
R915 B.n492 B.n287 163.367
R916 B.n488 B.n486 163.367
R917 B.n484 B.n289 163.367
R918 B.n480 B.n478 163.367
R919 B.n476 B.n291 163.367
R920 B.n472 B.n470 163.367
R921 B.n468 B.n293 163.367
R922 B.n464 B.n462 163.367
R923 B.n460 B.n295 163.367
R924 B.n456 B.n454 163.367
R925 B.n451 B.n450 163.367
R926 B.n448 B.n301 163.367
R927 B.n444 B.n442 163.367
R928 B.n440 B.n303 163.367
R929 B.n435 B.n433 163.367
R930 B.n431 B.n307 163.367
R931 B.n427 B.n425 163.367
R932 B.n423 B.n309 163.367
R933 B.n419 B.n417 163.367
R934 B.n415 B.n311 163.367
R935 B.n411 B.n409 163.367
R936 B.n407 B.n313 163.367
R937 B.n403 B.n401 163.367
R938 B.n399 B.n315 163.367
R939 B.n395 B.n393 163.367
R940 B.n391 B.n317 163.367
R941 B.n387 B.n385 163.367
R942 B.n383 B.n319 163.367
R943 B.n379 B.n377 163.367
R944 B.n375 B.n321 163.367
R945 B.n371 B.n369 163.367
R946 B.n367 B.n323 163.367
R947 B.n363 B.n361 163.367
R948 B.n359 B.n325 163.367
R949 B.n355 B.n353 163.367
R950 B.n351 B.n327 163.367
R951 B.n347 B.n345 163.367
R952 B.n343 B.n329 163.367
R953 B.n339 B.n337 163.367
R954 B.n335 B.n332 163.367
R955 B.n563 B.n265 163.367
R956 B.n567 B.n265 163.367
R957 B.n567 B.n259 163.367
R958 B.n575 B.n259 163.367
R959 B.n575 B.n257 163.367
R960 B.n579 B.n257 163.367
R961 B.n579 B.n252 163.367
R962 B.n588 B.n252 163.367
R963 B.n588 B.n250 163.367
R964 B.n592 B.n250 163.367
R965 B.n592 B.n244 163.367
R966 B.n600 B.n244 163.367
R967 B.n600 B.n242 163.367
R968 B.n604 B.n242 163.367
R969 B.n604 B.n235 163.367
R970 B.n612 B.n235 163.367
R971 B.n612 B.n233 163.367
R972 B.n616 B.n233 163.367
R973 B.n616 B.n228 163.367
R974 B.n624 B.n228 163.367
R975 B.n624 B.n226 163.367
R976 B.n628 B.n226 163.367
R977 B.n628 B.n219 163.367
R978 B.n636 B.n219 163.367
R979 B.n636 B.n217 163.367
R980 B.n640 B.n217 163.367
R981 B.n640 B.n212 163.367
R982 B.n648 B.n212 163.367
R983 B.n648 B.n210 163.367
R984 B.n652 B.n210 163.367
R985 B.n652 B.n203 163.367
R986 B.n660 B.n203 163.367
R987 B.n660 B.n201 163.367
R988 B.n664 B.n201 163.367
R989 B.n664 B.n196 163.367
R990 B.n672 B.n196 163.367
R991 B.n672 B.n194 163.367
R992 B.n676 B.n194 163.367
R993 B.n676 B.n188 163.367
R994 B.n684 B.n188 163.367
R995 B.n684 B.n186 163.367
R996 B.n688 B.n186 163.367
R997 B.n688 B.n180 163.367
R998 B.n696 B.n180 163.367
R999 B.n696 B.n178 163.367
R1000 B.n700 B.n178 163.367
R1001 B.n700 B.n172 163.367
R1002 B.n708 B.n172 163.367
R1003 B.n708 B.n170 163.367
R1004 B.n713 B.n170 163.367
R1005 B.n713 B.n164 163.367
R1006 B.n721 B.n164 163.367
R1007 B.n722 B.n721 163.367
R1008 B.n722 B.n5 163.367
R1009 B.n6 B.n5 163.367
R1010 B.n7 B.n6 163.367
R1011 B.n727 B.n7 163.367
R1012 B.n727 B.n12 163.367
R1013 B.n13 B.n12 163.367
R1014 B.n14 B.n13 163.367
R1015 B.n732 B.n14 163.367
R1016 B.n732 B.n19 163.367
R1017 B.n20 B.n19 163.367
R1018 B.n21 B.n20 163.367
R1019 B.n737 B.n21 163.367
R1020 B.n737 B.n26 163.367
R1021 B.n27 B.n26 163.367
R1022 B.n28 B.n27 163.367
R1023 B.n742 B.n28 163.367
R1024 B.n742 B.n33 163.367
R1025 B.n34 B.n33 163.367
R1026 B.n35 B.n34 163.367
R1027 B.n747 B.n35 163.367
R1028 B.n747 B.n40 163.367
R1029 B.n41 B.n40 163.367
R1030 B.n42 B.n41 163.367
R1031 B.n752 B.n42 163.367
R1032 B.n752 B.n47 163.367
R1033 B.n48 B.n47 163.367
R1034 B.n49 B.n48 163.367
R1035 B.n757 B.n49 163.367
R1036 B.n757 B.n54 163.367
R1037 B.n55 B.n54 163.367
R1038 B.n56 B.n55 163.367
R1039 B.n762 B.n56 163.367
R1040 B.n762 B.n61 163.367
R1041 B.n62 B.n61 163.367
R1042 B.n63 B.n62 163.367
R1043 B.n767 B.n63 163.367
R1044 B.n767 B.n68 163.367
R1045 B.n69 B.n68 163.367
R1046 B.n70 B.n69 163.367
R1047 B.n772 B.n70 163.367
R1048 B.n772 B.n75 163.367
R1049 B.n76 B.n75 163.367
R1050 B.n77 B.n76 163.367
R1051 B.n777 B.n77 163.367
R1052 B.n777 B.n82 163.367
R1053 B.n83 B.n82 163.367
R1054 B.n84 B.n83 163.367
R1055 B.n782 B.n84 163.367
R1056 B.n782 B.n89 163.367
R1057 B.n90 B.n89 163.367
R1058 B.n91 B.n90 163.367
R1059 B.n787 B.n91 163.367
R1060 B.n787 B.n96 163.367
R1061 B.n97 B.n96 163.367
R1062 B.n98 B.n97 163.367
R1063 B.n1019 B.n1017 163.367
R1064 B.n1015 B.n102 163.367
R1065 B.n1011 B.n1009 163.367
R1066 B.n1007 B.n104 163.367
R1067 B.n1003 B.n1001 163.367
R1068 B.n999 B.n106 163.367
R1069 B.n995 B.n993 163.367
R1070 B.n991 B.n108 163.367
R1071 B.n987 B.n985 163.367
R1072 B.n983 B.n110 163.367
R1073 B.n979 B.n977 163.367
R1074 B.n975 B.n112 163.367
R1075 B.n971 B.n969 163.367
R1076 B.n967 B.n114 163.367
R1077 B.n963 B.n961 163.367
R1078 B.n959 B.n116 163.367
R1079 B.n955 B.n953 163.367
R1080 B.n951 B.n118 163.367
R1081 B.n947 B.n945 163.367
R1082 B.n943 B.n120 163.367
R1083 B.n939 B.n937 163.367
R1084 B.n935 B.n122 163.367
R1085 B.n931 B.n929 163.367
R1086 B.n927 B.n124 163.367
R1087 B.n923 B.n921 163.367
R1088 B.n919 B.n126 163.367
R1089 B.n914 B.n912 163.367
R1090 B.n910 B.n130 163.367
R1091 B.n906 B.n904 163.367
R1092 B.n902 B.n132 163.367
R1093 B.n898 B.n896 163.367
R1094 B.n893 B.n892 163.367
R1095 B.n890 B.n138 163.367
R1096 B.n886 B.n884 163.367
R1097 B.n882 B.n140 163.367
R1098 B.n878 B.n876 163.367
R1099 B.n874 B.n142 163.367
R1100 B.n870 B.n868 163.367
R1101 B.n866 B.n144 163.367
R1102 B.n862 B.n860 163.367
R1103 B.n858 B.n146 163.367
R1104 B.n854 B.n852 163.367
R1105 B.n850 B.n148 163.367
R1106 B.n846 B.n844 163.367
R1107 B.n842 B.n150 163.367
R1108 B.n838 B.n836 163.367
R1109 B.n834 B.n152 163.367
R1110 B.n830 B.n828 163.367
R1111 B.n826 B.n154 163.367
R1112 B.n822 B.n820 163.367
R1113 B.n818 B.n156 163.367
R1114 B.n814 B.n812 163.367
R1115 B.n810 B.n158 163.367
R1116 B.n806 B.n804 163.367
R1117 B.n802 B.n160 163.367
R1118 B.n798 B.n796 163.367
R1119 B.n794 B.n162 163.367
R1120 B.n304 B.t13 121.891
R1121 B.n133 B.t16 121.891
R1122 B.n296 B.t20 121.871
R1123 B.n127 B.t22 121.871
R1124 B.n556 B.n269 71.676
R1125 B.n554 B.n271 71.676
R1126 B.n550 B.n549 71.676
R1127 B.n543 B.n273 71.676
R1128 B.n542 B.n541 71.676
R1129 B.n535 B.n275 71.676
R1130 B.n534 B.n533 71.676
R1131 B.n527 B.n277 71.676
R1132 B.n526 B.n525 71.676
R1133 B.n519 B.n279 71.676
R1134 B.n518 B.n517 71.676
R1135 B.n511 B.n281 71.676
R1136 B.n510 B.n509 71.676
R1137 B.n503 B.n283 71.676
R1138 B.n502 B.n501 71.676
R1139 B.n495 B.n285 71.676
R1140 B.n494 B.n493 71.676
R1141 B.n487 B.n287 71.676
R1142 B.n486 B.n485 71.676
R1143 B.n479 B.n289 71.676
R1144 B.n478 B.n477 71.676
R1145 B.n471 B.n291 71.676
R1146 B.n470 B.n469 71.676
R1147 B.n463 B.n293 71.676
R1148 B.n462 B.n461 71.676
R1149 B.n455 B.n295 71.676
R1150 B.n454 B.n299 71.676
R1151 B.n450 B.n449 71.676
R1152 B.n443 B.n301 71.676
R1153 B.n442 B.n441 71.676
R1154 B.n434 B.n303 71.676
R1155 B.n433 B.n432 71.676
R1156 B.n426 B.n307 71.676
R1157 B.n425 B.n424 71.676
R1158 B.n418 B.n309 71.676
R1159 B.n417 B.n416 71.676
R1160 B.n410 B.n311 71.676
R1161 B.n409 B.n408 71.676
R1162 B.n402 B.n313 71.676
R1163 B.n401 B.n400 71.676
R1164 B.n394 B.n315 71.676
R1165 B.n393 B.n392 71.676
R1166 B.n386 B.n317 71.676
R1167 B.n385 B.n384 71.676
R1168 B.n378 B.n319 71.676
R1169 B.n377 B.n376 71.676
R1170 B.n370 B.n321 71.676
R1171 B.n369 B.n368 71.676
R1172 B.n362 B.n323 71.676
R1173 B.n361 B.n360 71.676
R1174 B.n354 B.n325 71.676
R1175 B.n353 B.n352 71.676
R1176 B.n346 B.n327 71.676
R1177 B.n345 B.n344 71.676
R1178 B.n338 B.n329 71.676
R1179 B.n337 B.n336 71.676
R1180 B.n332 B.n331 71.676
R1181 B.n1018 B.n100 71.676
R1182 B.n1017 B.n1016 71.676
R1183 B.n1010 B.n102 71.676
R1184 B.n1009 B.n1008 71.676
R1185 B.n1002 B.n104 71.676
R1186 B.n1001 B.n1000 71.676
R1187 B.n994 B.n106 71.676
R1188 B.n993 B.n992 71.676
R1189 B.n986 B.n108 71.676
R1190 B.n985 B.n984 71.676
R1191 B.n978 B.n110 71.676
R1192 B.n977 B.n976 71.676
R1193 B.n970 B.n112 71.676
R1194 B.n969 B.n968 71.676
R1195 B.n962 B.n114 71.676
R1196 B.n961 B.n960 71.676
R1197 B.n954 B.n116 71.676
R1198 B.n953 B.n952 71.676
R1199 B.n946 B.n118 71.676
R1200 B.n945 B.n944 71.676
R1201 B.n938 B.n120 71.676
R1202 B.n937 B.n936 71.676
R1203 B.n930 B.n122 71.676
R1204 B.n929 B.n928 71.676
R1205 B.n922 B.n124 71.676
R1206 B.n921 B.n920 71.676
R1207 B.n913 B.n126 71.676
R1208 B.n912 B.n911 71.676
R1209 B.n905 B.n130 71.676
R1210 B.n904 B.n903 71.676
R1211 B.n897 B.n132 71.676
R1212 B.n896 B.n136 71.676
R1213 B.n892 B.n891 71.676
R1214 B.n885 B.n138 71.676
R1215 B.n884 B.n883 71.676
R1216 B.n877 B.n140 71.676
R1217 B.n876 B.n875 71.676
R1218 B.n869 B.n142 71.676
R1219 B.n868 B.n867 71.676
R1220 B.n861 B.n144 71.676
R1221 B.n860 B.n859 71.676
R1222 B.n853 B.n146 71.676
R1223 B.n852 B.n851 71.676
R1224 B.n845 B.n148 71.676
R1225 B.n844 B.n843 71.676
R1226 B.n837 B.n150 71.676
R1227 B.n836 B.n835 71.676
R1228 B.n829 B.n152 71.676
R1229 B.n828 B.n827 71.676
R1230 B.n821 B.n154 71.676
R1231 B.n820 B.n819 71.676
R1232 B.n813 B.n156 71.676
R1233 B.n812 B.n811 71.676
R1234 B.n805 B.n158 71.676
R1235 B.n804 B.n803 71.676
R1236 B.n797 B.n160 71.676
R1237 B.n796 B.n795 71.676
R1238 B.n795 B.n794 71.676
R1239 B.n798 B.n797 71.676
R1240 B.n803 B.n802 71.676
R1241 B.n806 B.n805 71.676
R1242 B.n811 B.n810 71.676
R1243 B.n814 B.n813 71.676
R1244 B.n819 B.n818 71.676
R1245 B.n822 B.n821 71.676
R1246 B.n827 B.n826 71.676
R1247 B.n830 B.n829 71.676
R1248 B.n835 B.n834 71.676
R1249 B.n838 B.n837 71.676
R1250 B.n843 B.n842 71.676
R1251 B.n846 B.n845 71.676
R1252 B.n851 B.n850 71.676
R1253 B.n854 B.n853 71.676
R1254 B.n859 B.n858 71.676
R1255 B.n862 B.n861 71.676
R1256 B.n867 B.n866 71.676
R1257 B.n870 B.n869 71.676
R1258 B.n875 B.n874 71.676
R1259 B.n878 B.n877 71.676
R1260 B.n883 B.n882 71.676
R1261 B.n886 B.n885 71.676
R1262 B.n891 B.n890 71.676
R1263 B.n893 B.n136 71.676
R1264 B.n898 B.n897 71.676
R1265 B.n903 B.n902 71.676
R1266 B.n906 B.n905 71.676
R1267 B.n911 B.n910 71.676
R1268 B.n914 B.n913 71.676
R1269 B.n920 B.n919 71.676
R1270 B.n923 B.n922 71.676
R1271 B.n928 B.n927 71.676
R1272 B.n931 B.n930 71.676
R1273 B.n936 B.n935 71.676
R1274 B.n939 B.n938 71.676
R1275 B.n944 B.n943 71.676
R1276 B.n947 B.n946 71.676
R1277 B.n952 B.n951 71.676
R1278 B.n955 B.n954 71.676
R1279 B.n960 B.n959 71.676
R1280 B.n963 B.n962 71.676
R1281 B.n968 B.n967 71.676
R1282 B.n971 B.n970 71.676
R1283 B.n976 B.n975 71.676
R1284 B.n979 B.n978 71.676
R1285 B.n984 B.n983 71.676
R1286 B.n987 B.n986 71.676
R1287 B.n992 B.n991 71.676
R1288 B.n995 B.n994 71.676
R1289 B.n1000 B.n999 71.676
R1290 B.n1003 B.n1002 71.676
R1291 B.n1008 B.n1007 71.676
R1292 B.n1011 B.n1010 71.676
R1293 B.n1016 B.n1015 71.676
R1294 B.n1019 B.n1018 71.676
R1295 B.n557 B.n556 71.676
R1296 B.n551 B.n271 71.676
R1297 B.n549 B.n548 71.676
R1298 B.n544 B.n543 71.676
R1299 B.n541 B.n540 71.676
R1300 B.n536 B.n535 71.676
R1301 B.n533 B.n532 71.676
R1302 B.n528 B.n527 71.676
R1303 B.n525 B.n524 71.676
R1304 B.n520 B.n519 71.676
R1305 B.n517 B.n516 71.676
R1306 B.n512 B.n511 71.676
R1307 B.n509 B.n508 71.676
R1308 B.n504 B.n503 71.676
R1309 B.n501 B.n500 71.676
R1310 B.n496 B.n495 71.676
R1311 B.n493 B.n492 71.676
R1312 B.n488 B.n487 71.676
R1313 B.n485 B.n484 71.676
R1314 B.n480 B.n479 71.676
R1315 B.n477 B.n476 71.676
R1316 B.n472 B.n471 71.676
R1317 B.n469 B.n468 71.676
R1318 B.n464 B.n463 71.676
R1319 B.n461 B.n460 71.676
R1320 B.n456 B.n455 71.676
R1321 B.n451 B.n299 71.676
R1322 B.n449 B.n448 71.676
R1323 B.n444 B.n443 71.676
R1324 B.n441 B.n440 71.676
R1325 B.n435 B.n434 71.676
R1326 B.n432 B.n431 71.676
R1327 B.n427 B.n426 71.676
R1328 B.n424 B.n423 71.676
R1329 B.n419 B.n418 71.676
R1330 B.n416 B.n415 71.676
R1331 B.n411 B.n410 71.676
R1332 B.n408 B.n407 71.676
R1333 B.n403 B.n402 71.676
R1334 B.n400 B.n399 71.676
R1335 B.n395 B.n394 71.676
R1336 B.n392 B.n391 71.676
R1337 B.n387 B.n386 71.676
R1338 B.n384 B.n383 71.676
R1339 B.n379 B.n378 71.676
R1340 B.n376 B.n375 71.676
R1341 B.n371 B.n370 71.676
R1342 B.n368 B.n367 71.676
R1343 B.n363 B.n362 71.676
R1344 B.n360 B.n359 71.676
R1345 B.n355 B.n354 71.676
R1346 B.n352 B.n351 71.676
R1347 B.n347 B.n346 71.676
R1348 B.n344 B.n343 71.676
R1349 B.n339 B.n338 71.676
R1350 B.n336 B.n335 71.676
R1351 B.n331 B.n267 71.676
R1352 B.n305 B.t12 71.4673
R1353 B.n134 B.t17 71.4673
R1354 B.n297 B.t19 71.4466
R1355 B.n128 B.t23 71.4466
R1356 B.n562 B.n268 64.0478
R1357 B.n1024 B.n99 64.0478
R1358 B.n437 B.n305 59.5399
R1359 B.n298 B.n297 59.5399
R1360 B.n916 B.n128 59.5399
R1361 B.n135 B.n134 59.5399
R1362 B.n305 B.n304 50.4247
R1363 B.n297 B.n296 50.4247
R1364 B.n128 B.n127 50.4247
R1365 B.n134 B.n133 50.4247
R1366 B.n562 B.n264 35.4088
R1367 B.n568 B.n264 35.4088
R1368 B.n568 B.n260 35.4088
R1369 B.n574 B.n260 35.4088
R1370 B.n574 B.n256 35.4088
R1371 B.n581 B.n256 35.4088
R1372 B.n581 B.n580 35.4088
R1373 B.n587 B.n249 35.4088
R1374 B.n593 B.n249 35.4088
R1375 B.n593 B.n245 35.4088
R1376 B.n599 B.n245 35.4088
R1377 B.n599 B.n241 35.4088
R1378 B.n605 B.n241 35.4088
R1379 B.n605 B.n236 35.4088
R1380 B.n611 B.n236 35.4088
R1381 B.n611 B.n237 35.4088
R1382 B.n617 B.n229 35.4088
R1383 B.n623 B.n229 35.4088
R1384 B.n623 B.n225 35.4088
R1385 B.n629 B.n225 35.4088
R1386 B.n629 B.n220 35.4088
R1387 B.n635 B.n220 35.4088
R1388 B.n635 B.n221 35.4088
R1389 B.n641 B.n213 35.4088
R1390 B.n647 B.n213 35.4088
R1391 B.n647 B.n209 35.4088
R1392 B.n653 B.n209 35.4088
R1393 B.n653 B.n204 35.4088
R1394 B.n659 B.n204 35.4088
R1395 B.n659 B.n205 35.4088
R1396 B.n665 B.n197 35.4088
R1397 B.n671 B.n197 35.4088
R1398 B.n671 B.n193 35.4088
R1399 B.n677 B.n193 35.4088
R1400 B.n677 B.n189 35.4088
R1401 B.n683 B.n189 35.4088
R1402 B.n689 B.n185 35.4088
R1403 B.n689 B.n181 35.4088
R1404 B.n695 B.n181 35.4088
R1405 B.n695 B.n177 35.4088
R1406 B.n701 B.n177 35.4088
R1407 B.n701 B.n173 35.4088
R1408 B.n707 B.n173 35.4088
R1409 B.n714 B.n169 35.4088
R1410 B.n714 B.n165 35.4088
R1411 B.n720 B.n165 35.4088
R1412 B.n720 B.n4 35.4088
R1413 B.n1130 B.n4 35.4088
R1414 B.n1130 B.n1129 35.4088
R1415 B.n1129 B.n1128 35.4088
R1416 B.n1128 B.n8 35.4088
R1417 B.n1122 B.n8 35.4088
R1418 B.n1122 B.n1121 35.4088
R1419 B.n1120 B.n15 35.4088
R1420 B.n1114 B.n15 35.4088
R1421 B.n1114 B.n1113 35.4088
R1422 B.n1113 B.n1112 35.4088
R1423 B.n1112 B.n22 35.4088
R1424 B.n1106 B.n22 35.4088
R1425 B.n1106 B.n1105 35.4088
R1426 B.n1104 B.n29 35.4088
R1427 B.n1098 B.n29 35.4088
R1428 B.n1098 B.n1097 35.4088
R1429 B.n1097 B.n1096 35.4088
R1430 B.n1096 B.n36 35.4088
R1431 B.n1090 B.n36 35.4088
R1432 B.n1089 B.n1088 35.4088
R1433 B.n1088 B.n43 35.4088
R1434 B.n1082 B.n43 35.4088
R1435 B.n1082 B.n1081 35.4088
R1436 B.n1081 B.n1080 35.4088
R1437 B.n1080 B.n50 35.4088
R1438 B.n1074 B.n50 35.4088
R1439 B.n1073 B.n1072 35.4088
R1440 B.n1072 B.n57 35.4088
R1441 B.n1066 B.n57 35.4088
R1442 B.n1066 B.n1065 35.4088
R1443 B.n1065 B.n1064 35.4088
R1444 B.n1064 B.n64 35.4088
R1445 B.n1058 B.n64 35.4088
R1446 B.n1057 B.n1056 35.4088
R1447 B.n1056 B.n71 35.4088
R1448 B.n1050 B.n71 35.4088
R1449 B.n1050 B.n1049 35.4088
R1450 B.n1049 B.n1048 35.4088
R1451 B.n1048 B.n78 35.4088
R1452 B.n1042 B.n78 35.4088
R1453 B.n1042 B.n1041 35.4088
R1454 B.n1041 B.n1040 35.4088
R1455 B.n1034 B.n88 35.4088
R1456 B.n1034 B.n1033 35.4088
R1457 B.n1033 B.n1032 35.4088
R1458 B.n1032 B.n92 35.4088
R1459 B.n1026 B.n92 35.4088
R1460 B.n1026 B.n1025 35.4088
R1461 B.n1025 B.n1024 35.4088
R1462 B.n237 B.t6 34.8881
R1463 B.t2 B.n1057 34.8881
R1464 B.n1022 B.n1021 34.8103
R1465 B.n792 B.n791 34.8103
R1466 B.n564 B.n266 34.8103
R1467 B.n560 B.n559 34.8103
R1468 B.n683 B.t7 32.8052
R1469 B.t0 B.n1104 32.8052
R1470 B.n587 B.t11 30.7224
R1471 B.n1040 B.t15 30.7224
R1472 B.n665 B.t8 25.5153
R1473 B.n1090 B.t3 25.5153
R1474 B.n221 B.t5 22.391
R1475 B.t1 B.n1073 22.391
R1476 B.n707 B.t9 20.3082
R1477 B.t4 B.n1120 20.3082
R1478 B B.n1132 18.0485
R1479 B.t9 B.n169 15.1011
R1480 B.n1121 B.t4 15.1011
R1481 B.n641 B.t5 13.0183
R1482 B.n1074 B.t1 13.0183
R1483 B.n1021 B.n1020 10.6151
R1484 B.n1020 B.n101 10.6151
R1485 B.n1014 B.n101 10.6151
R1486 B.n1014 B.n1013 10.6151
R1487 B.n1013 B.n1012 10.6151
R1488 B.n1012 B.n103 10.6151
R1489 B.n1006 B.n103 10.6151
R1490 B.n1006 B.n1005 10.6151
R1491 B.n1005 B.n1004 10.6151
R1492 B.n1004 B.n105 10.6151
R1493 B.n998 B.n105 10.6151
R1494 B.n998 B.n997 10.6151
R1495 B.n997 B.n996 10.6151
R1496 B.n996 B.n107 10.6151
R1497 B.n990 B.n107 10.6151
R1498 B.n990 B.n989 10.6151
R1499 B.n989 B.n988 10.6151
R1500 B.n988 B.n109 10.6151
R1501 B.n982 B.n109 10.6151
R1502 B.n982 B.n981 10.6151
R1503 B.n981 B.n980 10.6151
R1504 B.n980 B.n111 10.6151
R1505 B.n974 B.n111 10.6151
R1506 B.n974 B.n973 10.6151
R1507 B.n973 B.n972 10.6151
R1508 B.n972 B.n113 10.6151
R1509 B.n966 B.n113 10.6151
R1510 B.n966 B.n965 10.6151
R1511 B.n965 B.n964 10.6151
R1512 B.n964 B.n115 10.6151
R1513 B.n958 B.n115 10.6151
R1514 B.n958 B.n957 10.6151
R1515 B.n957 B.n956 10.6151
R1516 B.n956 B.n117 10.6151
R1517 B.n950 B.n117 10.6151
R1518 B.n950 B.n949 10.6151
R1519 B.n949 B.n948 10.6151
R1520 B.n948 B.n119 10.6151
R1521 B.n942 B.n119 10.6151
R1522 B.n942 B.n941 10.6151
R1523 B.n941 B.n940 10.6151
R1524 B.n940 B.n121 10.6151
R1525 B.n934 B.n121 10.6151
R1526 B.n934 B.n933 10.6151
R1527 B.n933 B.n932 10.6151
R1528 B.n932 B.n123 10.6151
R1529 B.n926 B.n123 10.6151
R1530 B.n926 B.n925 10.6151
R1531 B.n925 B.n924 10.6151
R1532 B.n924 B.n125 10.6151
R1533 B.n918 B.n125 10.6151
R1534 B.n918 B.n917 10.6151
R1535 B.n915 B.n129 10.6151
R1536 B.n909 B.n129 10.6151
R1537 B.n909 B.n908 10.6151
R1538 B.n908 B.n907 10.6151
R1539 B.n907 B.n131 10.6151
R1540 B.n901 B.n131 10.6151
R1541 B.n901 B.n900 10.6151
R1542 B.n900 B.n899 10.6151
R1543 B.n895 B.n894 10.6151
R1544 B.n894 B.n137 10.6151
R1545 B.n889 B.n137 10.6151
R1546 B.n889 B.n888 10.6151
R1547 B.n888 B.n887 10.6151
R1548 B.n887 B.n139 10.6151
R1549 B.n881 B.n139 10.6151
R1550 B.n881 B.n880 10.6151
R1551 B.n880 B.n879 10.6151
R1552 B.n879 B.n141 10.6151
R1553 B.n873 B.n141 10.6151
R1554 B.n873 B.n872 10.6151
R1555 B.n872 B.n871 10.6151
R1556 B.n871 B.n143 10.6151
R1557 B.n865 B.n143 10.6151
R1558 B.n865 B.n864 10.6151
R1559 B.n864 B.n863 10.6151
R1560 B.n863 B.n145 10.6151
R1561 B.n857 B.n145 10.6151
R1562 B.n857 B.n856 10.6151
R1563 B.n856 B.n855 10.6151
R1564 B.n855 B.n147 10.6151
R1565 B.n849 B.n147 10.6151
R1566 B.n849 B.n848 10.6151
R1567 B.n848 B.n847 10.6151
R1568 B.n847 B.n149 10.6151
R1569 B.n841 B.n149 10.6151
R1570 B.n841 B.n840 10.6151
R1571 B.n840 B.n839 10.6151
R1572 B.n839 B.n151 10.6151
R1573 B.n833 B.n151 10.6151
R1574 B.n833 B.n832 10.6151
R1575 B.n832 B.n831 10.6151
R1576 B.n831 B.n153 10.6151
R1577 B.n825 B.n153 10.6151
R1578 B.n825 B.n824 10.6151
R1579 B.n824 B.n823 10.6151
R1580 B.n823 B.n155 10.6151
R1581 B.n817 B.n155 10.6151
R1582 B.n817 B.n816 10.6151
R1583 B.n816 B.n815 10.6151
R1584 B.n815 B.n157 10.6151
R1585 B.n809 B.n157 10.6151
R1586 B.n809 B.n808 10.6151
R1587 B.n808 B.n807 10.6151
R1588 B.n807 B.n159 10.6151
R1589 B.n801 B.n159 10.6151
R1590 B.n801 B.n800 10.6151
R1591 B.n800 B.n799 10.6151
R1592 B.n799 B.n161 10.6151
R1593 B.n793 B.n161 10.6151
R1594 B.n793 B.n792 10.6151
R1595 B.n565 B.n564 10.6151
R1596 B.n566 B.n565 10.6151
R1597 B.n566 B.n258 10.6151
R1598 B.n576 B.n258 10.6151
R1599 B.n577 B.n576 10.6151
R1600 B.n578 B.n577 10.6151
R1601 B.n578 B.n251 10.6151
R1602 B.n589 B.n251 10.6151
R1603 B.n590 B.n589 10.6151
R1604 B.n591 B.n590 10.6151
R1605 B.n591 B.n243 10.6151
R1606 B.n601 B.n243 10.6151
R1607 B.n602 B.n601 10.6151
R1608 B.n603 B.n602 10.6151
R1609 B.n603 B.n234 10.6151
R1610 B.n613 B.n234 10.6151
R1611 B.n614 B.n613 10.6151
R1612 B.n615 B.n614 10.6151
R1613 B.n615 B.n227 10.6151
R1614 B.n625 B.n227 10.6151
R1615 B.n626 B.n625 10.6151
R1616 B.n627 B.n626 10.6151
R1617 B.n627 B.n218 10.6151
R1618 B.n637 B.n218 10.6151
R1619 B.n638 B.n637 10.6151
R1620 B.n639 B.n638 10.6151
R1621 B.n639 B.n211 10.6151
R1622 B.n649 B.n211 10.6151
R1623 B.n650 B.n649 10.6151
R1624 B.n651 B.n650 10.6151
R1625 B.n651 B.n202 10.6151
R1626 B.n661 B.n202 10.6151
R1627 B.n662 B.n661 10.6151
R1628 B.n663 B.n662 10.6151
R1629 B.n663 B.n195 10.6151
R1630 B.n673 B.n195 10.6151
R1631 B.n674 B.n673 10.6151
R1632 B.n675 B.n674 10.6151
R1633 B.n675 B.n187 10.6151
R1634 B.n685 B.n187 10.6151
R1635 B.n686 B.n685 10.6151
R1636 B.n687 B.n686 10.6151
R1637 B.n687 B.n179 10.6151
R1638 B.n697 B.n179 10.6151
R1639 B.n698 B.n697 10.6151
R1640 B.n699 B.n698 10.6151
R1641 B.n699 B.n171 10.6151
R1642 B.n709 B.n171 10.6151
R1643 B.n710 B.n709 10.6151
R1644 B.n712 B.n710 10.6151
R1645 B.n712 B.n711 10.6151
R1646 B.n711 B.n163 10.6151
R1647 B.n723 B.n163 10.6151
R1648 B.n724 B.n723 10.6151
R1649 B.n725 B.n724 10.6151
R1650 B.n726 B.n725 10.6151
R1651 B.n728 B.n726 10.6151
R1652 B.n729 B.n728 10.6151
R1653 B.n730 B.n729 10.6151
R1654 B.n731 B.n730 10.6151
R1655 B.n733 B.n731 10.6151
R1656 B.n734 B.n733 10.6151
R1657 B.n735 B.n734 10.6151
R1658 B.n736 B.n735 10.6151
R1659 B.n738 B.n736 10.6151
R1660 B.n739 B.n738 10.6151
R1661 B.n740 B.n739 10.6151
R1662 B.n741 B.n740 10.6151
R1663 B.n743 B.n741 10.6151
R1664 B.n744 B.n743 10.6151
R1665 B.n745 B.n744 10.6151
R1666 B.n746 B.n745 10.6151
R1667 B.n748 B.n746 10.6151
R1668 B.n749 B.n748 10.6151
R1669 B.n750 B.n749 10.6151
R1670 B.n751 B.n750 10.6151
R1671 B.n753 B.n751 10.6151
R1672 B.n754 B.n753 10.6151
R1673 B.n755 B.n754 10.6151
R1674 B.n756 B.n755 10.6151
R1675 B.n758 B.n756 10.6151
R1676 B.n759 B.n758 10.6151
R1677 B.n760 B.n759 10.6151
R1678 B.n761 B.n760 10.6151
R1679 B.n763 B.n761 10.6151
R1680 B.n764 B.n763 10.6151
R1681 B.n765 B.n764 10.6151
R1682 B.n766 B.n765 10.6151
R1683 B.n768 B.n766 10.6151
R1684 B.n769 B.n768 10.6151
R1685 B.n770 B.n769 10.6151
R1686 B.n771 B.n770 10.6151
R1687 B.n773 B.n771 10.6151
R1688 B.n774 B.n773 10.6151
R1689 B.n775 B.n774 10.6151
R1690 B.n776 B.n775 10.6151
R1691 B.n778 B.n776 10.6151
R1692 B.n779 B.n778 10.6151
R1693 B.n780 B.n779 10.6151
R1694 B.n781 B.n780 10.6151
R1695 B.n783 B.n781 10.6151
R1696 B.n784 B.n783 10.6151
R1697 B.n785 B.n784 10.6151
R1698 B.n786 B.n785 10.6151
R1699 B.n788 B.n786 10.6151
R1700 B.n789 B.n788 10.6151
R1701 B.n790 B.n789 10.6151
R1702 B.n791 B.n790 10.6151
R1703 B.n559 B.n558 10.6151
R1704 B.n558 B.n270 10.6151
R1705 B.n553 B.n270 10.6151
R1706 B.n553 B.n552 10.6151
R1707 B.n552 B.n272 10.6151
R1708 B.n547 B.n272 10.6151
R1709 B.n547 B.n546 10.6151
R1710 B.n546 B.n545 10.6151
R1711 B.n545 B.n274 10.6151
R1712 B.n539 B.n274 10.6151
R1713 B.n539 B.n538 10.6151
R1714 B.n538 B.n537 10.6151
R1715 B.n537 B.n276 10.6151
R1716 B.n531 B.n276 10.6151
R1717 B.n531 B.n530 10.6151
R1718 B.n530 B.n529 10.6151
R1719 B.n529 B.n278 10.6151
R1720 B.n523 B.n278 10.6151
R1721 B.n523 B.n522 10.6151
R1722 B.n522 B.n521 10.6151
R1723 B.n521 B.n280 10.6151
R1724 B.n515 B.n280 10.6151
R1725 B.n515 B.n514 10.6151
R1726 B.n514 B.n513 10.6151
R1727 B.n513 B.n282 10.6151
R1728 B.n507 B.n282 10.6151
R1729 B.n507 B.n506 10.6151
R1730 B.n506 B.n505 10.6151
R1731 B.n505 B.n284 10.6151
R1732 B.n499 B.n284 10.6151
R1733 B.n499 B.n498 10.6151
R1734 B.n498 B.n497 10.6151
R1735 B.n497 B.n286 10.6151
R1736 B.n491 B.n286 10.6151
R1737 B.n491 B.n490 10.6151
R1738 B.n490 B.n489 10.6151
R1739 B.n489 B.n288 10.6151
R1740 B.n483 B.n288 10.6151
R1741 B.n483 B.n482 10.6151
R1742 B.n482 B.n481 10.6151
R1743 B.n481 B.n290 10.6151
R1744 B.n475 B.n290 10.6151
R1745 B.n475 B.n474 10.6151
R1746 B.n474 B.n473 10.6151
R1747 B.n473 B.n292 10.6151
R1748 B.n467 B.n292 10.6151
R1749 B.n467 B.n466 10.6151
R1750 B.n466 B.n465 10.6151
R1751 B.n465 B.n294 10.6151
R1752 B.n459 B.n294 10.6151
R1753 B.n459 B.n458 10.6151
R1754 B.n458 B.n457 10.6151
R1755 B.n453 B.n452 10.6151
R1756 B.n452 B.n300 10.6151
R1757 B.n447 B.n300 10.6151
R1758 B.n447 B.n446 10.6151
R1759 B.n446 B.n445 10.6151
R1760 B.n445 B.n302 10.6151
R1761 B.n439 B.n302 10.6151
R1762 B.n439 B.n438 10.6151
R1763 B.n436 B.n306 10.6151
R1764 B.n430 B.n306 10.6151
R1765 B.n430 B.n429 10.6151
R1766 B.n429 B.n428 10.6151
R1767 B.n428 B.n308 10.6151
R1768 B.n422 B.n308 10.6151
R1769 B.n422 B.n421 10.6151
R1770 B.n421 B.n420 10.6151
R1771 B.n420 B.n310 10.6151
R1772 B.n414 B.n310 10.6151
R1773 B.n414 B.n413 10.6151
R1774 B.n413 B.n412 10.6151
R1775 B.n412 B.n312 10.6151
R1776 B.n406 B.n312 10.6151
R1777 B.n406 B.n405 10.6151
R1778 B.n405 B.n404 10.6151
R1779 B.n404 B.n314 10.6151
R1780 B.n398 B.n314 10.6151
R1781 B.n398 B.n397 10.6151
R1782 B.n397 B.n396 10.6151
R1783 B.n396 B.n316 10.6151
R1784 B.n390 B.n316 10.6151
R1785 B.n390 B.n389 10.6151
R1786 B.n389 B.n388 10.6151
R1787 B.n388 B.n318 10.6151
R1788 B.n382 B.n318 10.6151
R1789 B.n382 B.n381 10.6151
R1790 B.n381 B.n380 10.6151
R1791 B.n380 B.n320 10.6151
R1792 B.n374 B.n320 10.6151
R1793 B.n374 B.n373 10.6151
R1794 B.n373 B.n372 10.6151
R1795 B.n372 B.n322 10.6151
R1796 B.n366 B.n322 10.6151
R1797 B.n366 B.n365 10.6151
R1798 B.n365 B.n364 10.6151
R1799 B.n364 B.n324 10.6151
R1800 B.n358 B.n324 10.6151
R1801 B.n358 B.n357 10.6151
R1802 B.n357 B.n356 10.6151
R1803 B.n356 B.n326 10.6151
R1804 B.n350 B.n326 10.6151
R1805 B.n350 B.n349 10.6151
R1806 B.n349 B.n348 10.6151
R1807 B.n348 B.n328 10.6151
R1808 B.n342 B.n328 10.6151
R1809 B.n342 B.n341 10.6151
R1810 B.n341 B.n340 10.6151
R1811 B.n340 B.n330 10.6151
R1812 B.n334 B.n330 10.6151
R1813 B.n334 B.n333 10.6151
R1814 B.n333 B.n266 10.6151
R1815 B.n560 B.n262 10.6151
R1816 B.n570 B.n262 10.6151
R1817 B.n571 B.n570 10.6151
R1818 B.n572 B.n571 10.6151
R1819 B.n572 B.n254 10.6151
R1820 B.n583 B.n254 10.6151
R1821 B.n584 B.n583 10.6151
R1822 B.n585 B.n584 10.6151
R1823 B.n585 B.n247 10.6151
R1824 B.n595 B.n247 10.6151
R1825 B.n596 B.n595 10.6151
R1826 B.n597 B.n596 10.6151
R1827 B.n597 B.n239 10.6151
R1828 B.n607 B.n239 10.6151
R1829 B.n608 B.n607 10.6151
R1830 B.n609 B.n608 10.6151
R1831 B.n609 B.n231 10.6151
R1832 B.n619 B.n231 10.6151
R1833 B.n620 B.n619 10.6151
R1834 B.n621 B.n620 10.6151
R1835 B.n621 B.n223 10.6151
R1836 B.n631 B.n223 10.6151
R1837 B.n632 B.n631 10.6151
R1838 B.n633 B.n632 10.6151
R1839 B.n633 B.n215 10.6151
R1840 B.n643 B.n215 10.6151
R1841 B.n644 B.n643 10.6151
R1842 B.n645 B.n644 10.6151
R1843 B.n645 B.n207 10.6151
R1844 B.n655 B.n207 10.6151
R1845 B.n656 B.n655 10.6151
R1846 B.n657 B.n656 10.6151
R1847 B.n657 B.n199 10.6151
R1848 B.n667 B.n199 10.6151
R1849 B.n668 B.n667 10.6151
R1850 B.n669 B.n668 10.6151
R1851 B.n669 B.n191 10.6151
R1852 B.n679 B.n191 10.6151
R1853 B.n680 B.n679 10.6151
R1854 B.n681 B.n680 10.6151
R1855 B.n681 B.n183 10.6151
R1856 B.n691 B.n183 10.6151
R1857 B.n692 B.n691 10.6151
R1858 B.n693 B.n692 10.6151
R1859 B.n693 B.n175 10.6151
R1860 B.n703 B.n175 10.6151
R1861 B.n704 B.n703 10.6151
R1862 B.n705 B.n704 10.6151
R1863 B.n705 B.n167 10.6151
R1864 B.n716 B.n167 10.6151
R1865 B.n717 B.n716 10.6151
R1866 B.n718 B.n717 10.6151
R1867 B.n718 B.n0 10.6151
R1868 B.n1126 B.n1 10.6151
R1869 B.n1126 B.n1125 10.6151
R1870 B.n1125 B.n1124 10.6151
R1871 B.n1124 B.n10 10.6151
R1872 B.n1118 B.n10 10.6151
R1873 B.n1118 B.n1117 10.6151
R1874 B.n1117 B.n1116 10.6151
R1875 B.n1116 B.n17 10.6151
R1876 B.n1110 B.n17 10.6151
R1877 B.n1110 B.n1109 10.6151
R1878 B.n1109 B.n1108 10.6151
R1879 B.n1108 B.n24 10.6151
R1880 B.n1102 B.n24 10.6151
R1881 B.n1102 B.n1101 10.6151
R1882 B.n1101 B.n1100 10.6151
R1883 B.n1100 B.n31 10.6151
R1884 B.n1094 B.n31 10.6151
R1885 B.n1094 B.n1093 10.6151
R1886 B.n1093 B.n1092 10.6151
R1887 B.n1092 B.n38 10.6151
R1888 B.n1086 B.n38 10.6151
R1889 B.n1086 B.n1085 10.6151
R1890 B.n1085 B.n1084 10.6151
R1891 B.n1084 B.n45 10.6151
R1892 B.n1078 B.n45 10.6151
R1893 B.n1078 B.n1077 10.6151
R1894 B.n1077 B.n1076 10.6151
R1895 B.n1076 B.n52 10.6151
R1896 B.n1070 B.n52 10.6151
R1897 B.n1070 B.n1069 10.6151
R1898 B.n1069 B.n1068 10.6151
R1899 B.n1068 B.n59 10.6151
R1900 B.n1062 B.n59 10.6151
R1901 B.n1062 B.n1061 10.6151
R1902 B.n1061 B.n1060 10.6151
R1903 B.n1060 B.n66 10.6151
R1904 B.n1054 B.n66 10.6151
R1905 B.n1054 B.n1053 10.6151
R1906 B.n1053 B.n1052 10.6151
R1907 B.n1052 B.n73 10.6151
R1908 B.n1046 B.n73 10.6151
R1909 B.n1046 B.n1045 10.6151
R1910 B.n1045 B.n1044 10.6151
R1911 B.n1044 B.n80 10.6151
R1912 B.n1038 B.n80 10.6151
R1913 B.n1038 B.n1037 10.6151
R1914 B.n1037 B.n1036 10.6151
R1915 B.n1036 B.n86 10.6151
R1916 B.n1030 B.n86 10.6151
R1917 B.n1030 B.n1029 10.6151
R1918 B.n1029 B.n1028 10.6151
R1919 B.n1028 B.n94 10.6151
R1920 B.n1022 B.n94 10.6151
R1921 B.n205 B.t8 9.89399
R1922 B.t3 B.n1089 9.89399
R1923 B.n916 B.n915 6.5566
R1924 B.n899 B.n135 6.5566
R1925 B.n453 B.n298 6.5566
R1926 B.n438 B.n437 6.5566
R1927 B.n580 B.t11 4.68689
R1928 B.n88 B.t15 4.68689
R1929 B.n917 B.n916 4.05904
R1930 B.n895 B.n135 4.05904
R1931 B.n457 B.n298 4.05904
R1932 B.n437 B.n436 4.05904
R1933 B.n1132 B.n0 2.81026
R1934 B.n1132 B.n1 2.81026
R1935 B.t7 B.n185 2.60405
R1936 B.n1105 B.t0 2.60405
R1937 B.n617 B.t6 0.52121
R1938 B.n1058 B.t2 0.52121
R1939 VN.n8 VN.t8 199.149
R1940 VN.n45 VN.t5 199.149
R1941 VN.n5 VN.t3 168.275
R1942 VN.n9 VN.t1 168.275
R1943 VN.n27 VN.t0 168.275
R1944 VN.n35 VN.t2 168.275
R1945 VN.n42 VN.t6 168.275
R1946 VN.n46 VN.t4 168.275
R1947 VN.n64 VN.t9 168.275
R1948 VN.n72 VN.t7 168.275
R1949 VN.n71 VN.n37 161.3
R1950 VN.n70 VN.n69 161.3
R1951 VN.n68 VN.n38 161.3
R1952 VN.n67 VN.n66 161.3
R1953 VN.n65 VN.n39 161.3
R1954 VN.n63 VN.n62 161.3
R1955 VN.n61 VN.n40 161.3
R1956 VN.n60 VN.n59 161.3
R1957 VN.n58 VN.n41 161.3
R1958 VN.n57 VN.n56 161.3
R1959 VN.n55 VN.n42 161.3
R1960 VN.n54 VN.n53 161.3
R1961 VN.n52 VN.n43 161.3
R1962 VN.n51 VN.n50 161.3
R1963 VN.n49 VN.n44 161.3
R1964 VN.n48 VN.n47 161.3
R1965 VN.n34 VN.n0 161.3
R1966 VN.n33 VN.n32 161.3
R1967 VN.n31 VN.n1 161.3
R1968 VN.n30 VN.n29 161.3
R1969 VN.n28 VN.n2 161.3
R1970 VN.n26 VN.n25 161.3
R1971 VN.n24 VN.n3 161.3
R1972 VN.n23 VN.n22 161.3
R1973 VN.n21 VN.n4 161.3
R1974 VN.n20 VN.n19 161.3
R1975 VN.n18 VN.n5 161.3
R1976 VN.n17 VN.n16 161.3
R1977 VN.n15 VN.n6 161.3
R1978 VN.n14 VN.n13 161.3
R1979 VN.n12 VN.n7 161.3
R1980 VN.n11 VN.n10 161.3
R1981 VN.n36 VN.n35 100.969
R1982 VN.n73 VN.n72 100.969
R1983 VN.n9 VN.n8 67.1934
R1984 VN.n46 VN.n45 67.1934
R1985 VN.n15 VN.n14 56.5193
R1986 VN.n22 VN.n21 56.5193
R1987 VN.n52 VN.n51 56.5193
R1988 VN.n59 VN.n58 56.5193
R1989 VN VN.n73 54.4527
R1990 VN.n29 VN.n1 50.2061
R1991 VN.n66 VN.n38 50.2061
R1992 VN.n33 VN.n1 30.7807
R1993 VN.n70 VN.n38 30.7807
R1994 VN.n10 VN.n7 24.4675
R1995 VN.n14 VN.n7 24.4675
R1996 VN.n16 VN.n15 24.4675
R1997 VN.n16 VN.n5 24.4675
R1998 VN.n20 VN.n5 24.4675
R1999 VN.n21 VN.n20 24.4675
R2000 VN.n22 VN.n3 24.4675
R2001 VN.n26 VN.n3 24.4675
R2002 VN.n29 VN.n28 24.4675
R2003 VN.n34 VN.n33 24.4675
R2004 VN.n51 VN.n44 24.4675
R2005 VN.n47 VN.n44 24.4675
R2006 VN.n58 VN.n57 24.4675
R2007 VN.n57 VN.n42 24.4675
R2008 VN.n53 VN.n42 24.4675
R2009 VN.n53 VN.n52 24.4675
R2010 VN.n66 VN.n65 24.4675
R2011 VN.n63 VN.n40 24.4675
R2012 VN.n59 VN.n40 24.4675
R2013 VN.n71 VN.n70 24.4675
R2014 VN.n28 VN.n27 19.5741
R2015 VN.n65 VN.n64 19.5741
R2016 VN.n48 VN.n45 10.026
R2017 VN.n11 VN.n8 10.026
R2018 VN.n35 VN.n34 9.7873
R2019 VN.n72 VN.n71 9.7873
R2020 VN.n10 VN.n9 4.8939
R2021 VN.n27 VN.n26 4.8939
R2022 VN.n47 VN.n46 4.8939
R2023 VN.n64 VN.n63 4.8939
R2024 VN.n73 VN.n37 0.278367
R2025 VN.n36 VN.n0 0.278367
R2026 VN.n69 VN.n37 0.189894
R2027 VN.n69 VN.n68 0.189894
R2028 VN.n68 VN.n67 0.189894
R2029 VN.n67 VN.n39 0.189894
R2030 VN.n62 VN.n39 0.189894
R2031 VN.n62 VN.n61 0.189894
R2032 VN.n61 VN.n60 0.189894
R2033 VN.n60 VN.n41 0.189894
R2034 VN.n56 VN.n41 0.189894
R2035 VN.n56 VN.n55 0.189894
R2036 VN.n55 VN.n54 0.189894
R2037 VN.n54 VN.n43 0.189894
R2038 VN.n50 VN.n43 0.189894
R2039 VN.n50 VN.n49 0.189894
R2040 VN.n49 VN.n48 0.189894
R2041 VN.n12 VN.n11 0.189894
R2042 VN.n13 VN.n12 0.189894
R2043 VN.n13 VN.n6 0.189894
R2044 VN.n17 VN.n6 0.189894
R2045 VN.n18 VN.n17 0.189894
R2046 VN.n19 VN.n18 0.189894
R2047 VN.n19 VN.n4 0.189894
R2048 VN.n23 VN.n4 0.189894
R2049 VN.n24 VN.n23 0.189894
R2050 VN.n25 VN.n24 0.189894
R2051 VN.n25 VN.n2 0.189894
R2052 VN.n30 VN.n2 0.189894
R2053 VN.n31 VN.n30 0.189894
R2054 VN.n32 VN.n31 0.189894
R2055 VN.n32 VN.n0 0.189894
R2056 VN VN.n36 0.153454
R2057 VDD2.n1 VDD2.t3 66.8199
R2058 VDD2.n3 VDD2.n2 64.955
R2059 VDD2 VDD2.n7 64.9522
R2060 VDD2.n4 VDD2.t4 64.5787
R2061 VDD2.n6 VDD2.n5 63.3295
R2062 VDD2.n1 VDD2.n0 63.3293
R2063 VDD2.n4 VDD2.n3 48.0256
R2064 VDD2.n6 VDD2.n4 2.24188
R2065 VDD2.n7 VDD2.t0 1.24971
R2066 VDD2.n7 VDD2.t8 1.24971
R2067 VDD2.n5 VDD2.t9 1.24971
R2068 VDD2.n5 VDD2.t5 1.24971
R2069 VDD2.n2 VDD2.t6 1.24971
R2070 VDD2.n2 VDD2.t1 1.24971
R2071 VDD2.n0 VDD2.t7 1.24971
R2072 VDD2.n0 VDD2.t2 1.24971
R2073 VDD2 VDD2.n6 0.619035
R2074 VDD2.n3 VDD2.n1 0.505499
R2075 VTAIL.n11 VTAIL.t14 47.8999
R2076 VTAIL.n17 VTAIL.t17 47.8998
R2077 VTAIL.n2 VTAIL.t6 47.8998
R2078 VTAIL.n16 VTAIL.t9 47.8998
R2079 VTAIL.n15 VTAIL.n14 46.6507
R2080 VTAIL.n13 VTAIL.n12 46.6507
R2081 VTAIL.n10 VTAIL.n9 46.6507
R2082 VTAIL.n8 VTAIL.n7 46.6507
R2083 VTAIL.n19 VTAIL.n18 46.6505
R2084 VTAIL.n1 VTAIL.n0 46.6505
R2085 VTAIL.n4 VTAIL.n3 46.6505
R2086 VTAIL.n6 VTAIL.n5 46.6505
R2087 VTAIL.n8 VTAIL.n6 30.5134
R2088 VTAIL.n17 VTAIL.n16 28.2721
R2089 VTAIL.n10 VTAIL.n8 2.24188
R2090 VTAIL.n11 VTAIL.n10 2.24188
R2091 VTAIL.n15 VTAIL.n13 2.24188
R2092 VTAIL.n16 VTAIL.n15 2.24188
R2093 VTAIL.n6 VTAIL.n4 2.24188
R2094 VTAIL.n4 VTAIL.n2 2.24188
R2095 VTAIL.n19 VTAIL.n17 2.24188
R2096 VTAIL VTAIL.n1 1.73972
R2097 VTAIL.n13 VTAIL.n11 1.59102
R2098 VTAIL.n2 VTAIL.n1 1.59102
R2099 VTAIL.n18 VTAIL.t16 1.24971
R2100 VTAIL.n18 VTAIL.t19 1.24971
R2101 VTAIL.n0 VTAIL.t11 1.24971
R2102 VTAIL.n0 VTAIL.t18 1.24971
R2103 VTAIL.n3 VTAIL.t7 1.24971
R2104 VTAIL.n3 VTAIL.t5 1.24971
R2105 VTAIL.n5 VTAIL.t4 1.24971
R2106 VTAIL.n5 VTAIL.t8 1.24971
R2107 VTAIL.n14 VTAIL.t2 1.24971
R2108 VTAIL.n14 VTAIL.t1 1.24971
R2109 VTAIL.n12 VTAIL.t3 1.24971
R2110 VTAIL.n12 VTAIL.t0 1.24971
R2111 VTAIL.n9 VTAIL.t13 1.24971
R2112 VTAIL.n9 VTAIL.t15 1.24971
R2113 VTAIL.n7 VTAIL.t12 1.24971
R2114 VTAIL.n7 VTAIL.t10 1.24971
R2115 VTAIL VTAIL.n19 0.502655
R2116 VP.n19 VP.t7 199.149
R2117 VP.n5 VP.t0 168.275
R2118 VP.n49 VP.t3 168.275
R2119 VP.n57 VP.t6 168.275
R2120 VP.n75 VP.t2 168.275
R2121 VP.n83 VP.t1 168.275
R2122 VP.n16 VP.t8 168.275
R2123 VP.n46 VP.t4 168.275
R2124 VP.n38 VP.t5 168.275
R2125 VP.n20 VP.t9 168.275
R2126 VP.n22 VP.n21 161.3
R2127 VP.n23 VP.n18 161.3
R2128 VP.n25 VP.n24 161.3
R2129 VP.n26 VP.n17 161.3
R2130 VP.n28 VP.n27 161.3
R2131 VP.n29 VP.n16 161.3
R2132 VP.n31 VP.n30 161.3
R2133 VP.n32 VP.n15 161.3
R2134 VP.n34 VP.n33 161.3
R2135 VP.n35 VP.n14 161.3
R2136 VP.n37 VP.n36 161.3
R2137 VP.n39 VP.n13 161.3
R2138 VP.n41 VP.n40 161.3
R2139 VP.n42 VP.n12 161.3
R2140 VP.n44 VP.n43 161.3
R2141 VP.n45 VP.n11 161.3
R2142 VP.n82 VP.n0 161.3
R2143 VP.n81 VP.n80 161.3
R2144 VP.n79 VP.n1 161.3
R2145 VP.n78 VP.n77 161.3
R2146 VP.n76 VP.n2 161.3
R2147 VP.n74 VP.n73 161.3
R2148 VP.n72 VP.n3 161.3
R2149 VP.n71 VP.n70 161.3
R2150 VP.n69 VP.n4 161.3
R2151 VP.n68 VP.n67 161.3
R2152 VP.n66 VP.n5 161.3
R2153 VP.n65 VP.n64 161.3
R2154 VP.n63 VP.n6 161.3
R2155 VP.n62 VP.n61 161.3
R2156 VP.n60 VP.n7 161.3
R2157 VP.n59 VP.n58 161.3
R2158 VP.n56 VP.n8 161.3
R2159 VP.n55 VP.n54 161.3
R2160 VP.n53 VP.n9 161.3
R2161 VP.n52 VP.n51 161.3
R2162 VP.n50 VP.n10 161.3
R2163 VP.n49 VP.n48 100.969
R2164 VP.n84 VP.n83 100.969
R2165 VP.n47 VP.n46 100.969
R2166 VP.n20 VP.n19 67.1934
R2167 VP.n63 VP.n62 56.5193
R2168 VP.n70 VP.n69 56.5193
R2169 VP.n33 VP.n32 56.5193
R2170 VP.n26 VP.n25 56.5193
R2171 VP.n48 VP.n47 54.1738
R2172 VP.n55 VP.n9 50.2061
R2173 VP.n77 VP.n1 50.2061
R2174 VP.n40 VP.n12 50.2061
R2175 VP.n51 VP.n9 30.7807
R2176 VP.n81 VP.n1 30.7807
R2177 VP.n44 VP.n12 30.7807
R2178 VP.n51 VP.n50 24.4675
R2179 VP.n56 VP.n55 24.4675
R2180 VP.n58 VP.n7 24.4675
R2181 VP.n62 VP.n7 24.4675
R2182 VP.n64 VP.n63 24.4675
R2183 VP.n64 VP.n5 24.4675
R2184 VP.n68 VP.n5 24.4675
R2185 VP.n69 VP.n68 24.4675
R2186 VP.n70 VP.n3 24.4675
R2187 VP.n74 VP.n3 24.4675
R2188 VP.n77 VP.n76 24.4675
R2189 VP.n82 VP.n81 24.4675
R2190 VP.n45 VP.n44 24.4675
R2191 VP.n33 VP.n14 24.4675
R2192 VP.n37 VP.n14 24.4675
R2193 VP.n40 VP.n39 24.4675
R2194 VP.n27 VP.n26 24.4675
R2195 VP.n27 VP.n16 24.4675
R2196 VP.n31 VP.n16 24.4675
R2197 VP.n32 VP.n31 24.4675
R2198 VP.n21 VP.n18 24.4675
R2199 VP.n25 VP.n18 24.4675
R2200 VP.n57 VP.n56 19.5741
R2201 VP.n76 VP.n75 19.5741
R2202 VP.n39 VP.n38 19.5741
R2203 VP.n22 VP.n19 10.026
R2204 VP.n50 VP.n49 9.7873
R2205 VP.n83 VP.n82 9.7873
R2206 VP.n46 VP.n45 9.7873
R2207 VP.n58 VP.n57 4.8939
R2208 VP.n75 VP.n74 4.8939
R2209 VP.n38 VP.n37 4.8939
R2210 VP.n21 VP.n20 4.8939
R2211 VP.n47 VP.n11 0.278367
R2212 VP.n48 VP.n10 0.278367
R2213 VP.n84 VP.n0 0.278367
R2214 VP.n23 VP.n22 0.189894
R2215 VP.n24 VP.n23 0.189894
R2216 VP.n24 VP.n17 0.189894
R2217 VP.n28 VP.n17 0.189894
R2218 VP.n29 VP.n28 0.189894
R2219 VP.n30 VP.n29 0.189894
R2220 VP.n30 VP.n15 0.189894
R2221 VP.n34 VP.n15 0.189894
R2222 VP.n35 VP.n34 0.189894
R2223 VP.n36 VP.n35 0.189894
R2224 VP.n36 VP.n13 0.189894
R2225 VP.n41 VP.n13 0.189894
R2226 VP.n42 VP.n41 0.189894
R2227 VP.n43 VP.n42 0.189894
R2228 VP.n43 VP.n11 0.189894
R2229 VP.n52 VP.n10 0.189894
R2230 VP.n53 VP.n52 0.189894
R2231 VP.n54 VP.n53 0.189894
R2232 VP.n54 VP.n8 0.189894
R2233 VP.n59 VP.n8 0.189894
R2234 VP.n60 VP.n59 0.189894
R2235 VP.n61 VP.n60 0.189894
R2236 VP.n61 VP.n6 0.189894
R2237 VP.n65 VP.n6 0.189894
R2238 VP.n66 VP.n65 0.189894
R2239 VP.n67 VP.n66 0.189894
R2240 VP.n67 VP.n4 0.189894
R2241 VP.n71 VP.n4 0.189894
R2242 VP.n72 VP.n71 0.189894
R2243 VP.n73 VP.n72 0.189894
R2244 VP.n73 VP.n2 0.189894
R2245 VP.n78 VP.n2 0.189894
R2246 VP.n79 VP.n78 0.189894
R2247 VP.n80 VP.n79 0.189894
R2248 VP.n80 VP.n0 0.189894
R2249 VP VP.n84 0.153454
R2250 VDD1.n1 VDD1.t2 66.82
R2251 VDD1.n3 VDD1.t6 66.8199
R2252 VDD1.n5 VDD1.n4 64.955
R2253 VDD1.n1 VDD1.n0 63.3295
R2254 VDD1.n7 VDD1.n6 63.3293
R2255 VDD1.n3 VDD1.n2 63.3293
R2256 VDD1.n7 VDD1.n5 49.7293
R2257 VDD1 VDD1.n7 1.62334
R2258 VDD1.n6 VDD1.t4 1.24971
R2259 VDD1.n6 VDD1.t5 1.24971
R2260 VDD1.n0 VDD1.t0 1.24971
R2261 VDD1.n0 VDD1.t1 1.24971
R2262 VDD1.n4 VDD1.t7 1.24971
R2263 VDD1.n4 VDD1.t8 1.24971
R2264 VDD1.n2 VDD1.t3 1.24971
R2265 VDD1.n2 VDD1.t9 1.24971
R2266 VDD1 VDD1.n1 0.619035
R2267 VDD1.n5 VDD1.n3 0.505499
C0 VDD1 VTAIL 12.275499f
C1 VP VN 8.6291f
C2 VDD2 VN 13.5261f
C3 VP VDD2 0.541864f
C4 VN VTAIL 13.8628f
C5 VP VTAIL 13.8772f
C6 VDD2 VTAIL 12.3228f
C7 VDD1 VN 0.152635f
C8 VP VDD1 13.9108f
C9 VDD1 VDD2 1.96039f
C10 VDD2 B 7.464177f
C11 VDD1 B 7.468984f
C12 VTAIL B 9.469768f
C13 VN B 16.92205f
C14 VP B 15.345453f
C15 VDD1.t2 B 3.23565f
C16 VDD1.t0 B 0.278025f
C17 VDD1.t1 B 0.278025f
C18 VDD1.n0 B 2.5218f
C19 VDD1.n1 B 0.778476f
C20 VDD1.t6 B 3.23564f
C21 VDD1.t3 B 0.278025f
C22 VDD1.t9 B 0.278025f
C23 VDD1.n2 B 2.5218f
C24 VDD1.n3 B 0.77139f
C25 VDD1.t7 B 0.278025f
C26 VDD1.t8 B 0.278025f
C27 VDD1.n4 B 2.53346f
C28 VDD1.n5 B 2.74204f
C29 VDD1.t4 B 0.278025f
C30 VDD1.t5 B 0.278025f
C31 VDD1.n6 B 2.52179f
C32 VDD1.n7 B 2.95345f
C33 VP.n0 B 0.030339f
C34 VP.t1 B 2.27155f
C35 VP.n1 B 0.021739f
C36 VP.n2 B 0.023012f
C37 VP.t2 B 2.27155f
C38 VP.n3 B 0.042889f
C39 VP.n4 B 0.023012f
C40 VP.t0 B 2.27155f
C41 VP.n5 B 0.816336f
C42 VP.n6 B 0.023012f
C43 VP.n7 B 0.042889f
C44 VP.n8 B 0.023012f
C45 VP.t6 B 2.27155f
C46 VP.n9 B 0.021739f
C47 VP.n10 B 0.030339f
C48 VP.t3 B 2.27155f
C49 VP.n11 B 0.030339f
C50 VP.t4 B 2.27155f
C51 VP.n12 B 0.021739f
C52 VP.n13 B 0.023012f
C53 VP.t5 B 2.27155f
C54 VP.n14 B 0.042889f
C55 VP.n15 B 0.023012f
C56 VP.t8 B 2.27155f
C57 VP.n16 B 0.816336f
C58 VP.n17 B 0.023012f
C59 VP.n18 B 0.042889f
C60 VP.t7 B 2.41381f
C61 VP.n19 B 0.849954f
C62 VP.t9 B 2.27155f
C63 VP.n20 B 0.849813f
C64 VP.n21 B 0.025949f
C65 VP.n22 B 0.19714f
C66 VP.n23 B 0.023012f
C67 VP.n24 B 0.023012f
C68 VP.n25 B 0.030387f
C69 VP.n26 B 0.0368f
C70 VP.n27 B 0.042889f
C71 VP.n28 B 0.023012f
C72 VP.n29 B 0.023012f
C73 VP.n30 B 0.023012f
C74 VP.n31 B 0.042889f
C75 VP.n32 B 0.0368f
C76 VP.n33 B 0.030387f
C77 VP.n34 B 0.023012f
C78 VP.n35 B 0.023012f
C79 VP.n36 B 0.023012f
C80 VP.n37 B 0.025949f
C81 VP.n38 B 0.794622f
C82 VP.n39 B 0.038654f
C83 VP.n40 B 0.042236f
C84 VP.n41 B 0.023012f
C85 VP.n42 B 0.023012f
C86 VP.n43 B 0.023012f
C87 VP.n44 B 0.046101f
C88 VP.n45 B 0.030184f
C89 VP.n46 B 0.861205f
C90 VP.n47 B 1.43405f
C91 VP.n48 B 1.44932f
C92 VP.n49 B 0.861205f
C93 VP.n50 B 0.030184f
C94 VP.n51 B 0.046101f
C95 VP.n52 B 0.023012f
C96 VP.n53 B 0.023012f
C97 VP.n54 B 0.023012f
C98 VP.n55 B 0.042236f
C99 VP.n56 B 0.038654f
C100 VP.n57 B 0.794622f
C101 VP.n58 B 0.025949f
C102 VP.n59 B 0.023012f
C103 VP.n60 B 0.023012f
C104 VP.n61 B 0.023012f
C105 VP.n62 B 0.030387f
C106 VP.n63 B 0.0368f
C107 VP.n64 B 0.042889f
C108 VP.n65 B 0.023012f
C109 VP.n66 B 0.023012f
C110 VP.n67 B 0.023012f
C111 VP.n68 B 0.042889f
C112 VP.n69 B 0.0368f
C113 VP.n70 B 0.030387f
C114 VP.n71 B 0.023012f
C115 VP.n72 B 0.023012f
C116 VP.n73 B 0.023012f
C117 VP.n74 B 0.025949f
C118 VP.n75 B 0.794622f
C119 VP.n76 B 0.038654f
C120 VP.n77 B 0.042236f
C121 VP.n78 B 0.023012f
C122 VP.n79 B 0.023012f
C123 VP.n80 B 0.023012f
C124 VP.n81 B 0.046101f
C125 VP.n82 B 0.030184f
C126 VP.n83 B 0.861205f
C127 VP.n84 B 0.03518f
C128 VTAIL.t11 B 0.299518f
C129 VTAIL.t18 B 0.299518f
C130 VTAIL.n0 B 2.64899f
C131 VTAIL.n1 B 0.485885f
C132 VTAIL.t6 B 3.38327f
C133 VTAIL.n2 B 0.607165f
C134 VTAIL.t7 B 0.299518f
C135 VTAIL.t5 B 0.299518f
C136 VTAIL.n3 B 2.64899f
C137 VTAIL.n4 B 0.57473f
C138 VTAIL.t4 B 0.299518f
C139 VTAIL.t8 B 0.299518f
C140 VTAIL.n5 B 2.64899f
C141 VTAIL.n6 B 2.12512f
C142 VTAIL.t12 B 0.299518f
C143 VTAIL.t10 B 0.299518f
C144 VTAIL.n7 B 2.649f
C145 VTAIL.n8 B 2.12512f
C146 VTAIL.t13 B 0.299518f
C147 VTAIL.t15 B 0.299518f
C148 VTAIL.n9 B 2.649f
C149 VTAIL.n10 B 0.574726f
C150 VTAIL.t14 B 3.3833f
C151 VTAIL.n11 B 0.607144f
C152 VTAIL.t3 B 0.299518f
C153 VTAIL.t0 B 0.299518f
C154 VTAIL.n12 B 2.649f
C155 VTAIL.n13 B 0.524575f
C156 VTAIL.t2 B 0.299518f
C157 VTAIL.t1 B 0.299518f
C158 VTAIL.n14 B 2.649f
C159 VTAIL.n15 B 0.574726f
C160 VTAIL.t9 B 3.38327f
C161 VTAIL.n16 B 2.035f
C162 VTAIL.t17 B 3.38327f
C163 VTAIL.n17 B 2.035f
C164 VTAIL.t16 B 0.299518f
C165 VTAIL.t19 B 0.299518f
C166 VTAIL.n18 B 2.64899f
C167 VTAIL.n19 B 0.440715f
C168 VDD2.t3 B 3.19624f
C169 VDD2.t7 B 0.27464f
C170 VDD2.t2 B 0.27464f
C171 VDD2.n0 B 2.49109f
C172 VDD2.n1 B 0.761998f
C173 VDD2.t6 B 0.27464f
C174 VDD2.t1 B 0.27464f
C175 VDD2.n2 B 2.50261f
C176 VDD2.n3 B 2.6047f
C177 VDD2.t4 B 3.18275f
C178 VDD2.n4 B 2.88314f
C179 VDD2.t9 B 0.27464f
C180 VDD2.t5 B 0.27464f
C181 VDD2.n5 B 2.49109f
C182 VDD2.n6 B 0.380005f
C183 VDD2.t0 B 0.27464f
C184 VDD2.t8 B 0.27464f
C185 VDD2.n7 B 2.50257f
C186 VN.n0 B 0.029979f
C187 VN.t2 B 2.24459f
C188 VN.n1 B 0.021481f
C189 VN.n2 B 0.022739f
C190 VN.t0 B 2.24459f
C191 VN.n3 B 0.04238f
C192 VN.n4 B 0.022739f
C193 VN.t3 B 2.24459f
C194 VN.n5 B 0.806649f
C195 VN.n6 B 0.022739f
C196 VN.n7 B 0.04238f
C197 VN.t8 B 2.38517f
C198 VN.n8 B 0.839867f
C199 VN.t1 B 2.24459f
C200 VN.n9 B 0.839728f
C201 VN.n10 B 0.025641f
C202 VN.n11 B 0.1948f
C203 VN.n12 B 0.022739f
C204 VN.n13 B 0.022739f
C205 VN.n14 B 0.030027f
C206 VN.n15 B 0.036363f
C207 VN.n16 B 0.04238f
C208 VN.n17 B 0.022739f
C209 VN.n18 B 0.022739f
C210 VN.n19 B 0.022739f
C211 VN.n20 B 0.04238f
C212 VN.n21 B 0.036363f
C213 VN.n22 B 0.030027f
C214 VN.n23 B 0.022739f
C215 VN.n24 B 0.022739f
C216 VN.n25 B 0.022739f
C217 VN.n26 B 0.025641f
C218 VN.n27 B 0.785192f
C219 VN.n28 B 0.038195f
C220 VN.n29 B 0.041734f
C221 VN.n30 B 0.022739f
C222 VN.n31 B 0.022739f
C223 VN.n32 B 0.022739f
C224 VN.n33 B 0.045554f
C225 VN.n34 B 0.029826f
C226 VN.n35 B 0.850984f
C227 VN.n36 B 0.034763f
C228 VN.n37 B 0.029979f
C229 VN.t7 B 2.24459f
C230 VN.n38 B 0.021481f
C231 VN.n39 B 0.022739f
C232 VN.t9 B 2.24459f
C233 VN.n40 B 0.04238f
C234 VN.n41 B 0.022739f
C235 VN.t6 B 2.24459f
C236 VN.n42 B 0.806649f
C237 VN.n43 B 0.022739f
C238 VN.n44 B 0.04238f
C239 VN.t5 B 2.38517f
C240 VN.n45 B 0.839867f
C241 VN.t4 B 2.24459f
C242 VN.n46 B 0.839728f
C243 VN.n47 B 0.025641f
C244 VN.n48 B 0.1948f
C245 VN.n49 B 0.022739f
C246 VN.n50 B 0.022739f
C247 VN.n51 B 0.030027f
C248 VN.n52 B 0.036363f
C249 VN.n53 B 0.04238f
C250 VN.n54 B 0.022739f
C251 VN.n55 B 0.022739f
C252 VN.n56 B 0.022739f
C253 VN.n57 B 0.04238f
C254 VN.n58 B 0.036363f
C255 VN.n59 B 0.030027f
C256 VN.n60 B 0.022739f
C257 VN.n61 B 0.022739f
C258 VN.n62 B 0.022739f
C259 VN.n63 B 0.025641f
C260 VN.n64 B 0.785192f
C261 VN.n65 B 0.038195f
C262 VN.n66 B 0.041734f
C263 VN.n67 B 0.022739f
C264 VN.n68 B 0.022739f
C265 VN.n69 B 0.022739f
C266 VN.n70 B 0.045554f
C267 VN.n71 B 0.029826f
C268 VN.n72 B 0.850984f
C269 VN.n73 B 1.4291f
.ends

