* NGSPICE file created from diff_pair_sample_0481.ext - technology: sky130A

.subckt diff_pair_sample_0481 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t15 w_n2810_n4916# sky130_fd_pr__pfet_01v8 ad=3.2571 pd=20.07 as=3.2571 ps=20.07 w=19.74 l=1.51
X1 VTAIL.t14 VN.t1 VDD2.t6 w_n2810_n4916# sky130_fd_pr__pfet_01v8 ad=7.6986 pd=40.26 as=3.2571 ps=20.07 w=19.74 l=1.51
X2 VDD1.t7 VP.t0 VTAIL.t2 w_n2810_n4916# sky130_fd_pr__pfet_01v8 ad=3.2571 pd=20.07 as=7.6986 ps=40.26 w=19.74 l=1.51
X3 B.t11 B.t9 B.t10 w_n2810_n4916# sky130_fd_pr__pfet_01v8 ad=7.6986 pd=40.26 as=0 ps=0 w=19.74 l=1.51
X4 VTAIL.t6 VP.t1 VDD1.t6 w_n2810_n4916# sky130_fd_pr__pfet_01v8 ad=7.6986 pd=40.26 as=3.2571 ps=20.07 w=19.74 l=1.51
X5 VDD2.t5 VN.t2 VTAIL.t8 w_n2810_n4916# sky130_fd_pr__pfet_01v8 ad=3.2571 pd=20.07 as=7.6986 ps=40.26 w=19.74 l=1.51
X6 VDD1.t5 VP.t2 VTAIL.t7 w_n2810_n4916# sky130_fd_pr__pfet_01v8 ad=3.2571 pd=20.07 as=3.2571 ps=20.07 w=19.74 l=1.51
X7 B.t8 B.t6 B.t7 w_n2810_n4916# sky130_fd_pr__pfet_01v8 ad=7.6986 pd=40.26 as=0 ps=0 w=19.74 l=1.51
X8 VTAIL.t9 VN.t3 VDD2.t4 w_n2810_n4916# sky130_fd_pr__pfet_01v8 ad=3.2571 pd=20.07 as=3.2571 ps=20.07 w=19.74 l=1.51
X9 VDD2.t3 VN.t4 VTAIL.t12 w_n2810_n4916# sky130_fd_pr__pfet_01v8 ad=3.2571 pd=20.07 as=3.2571 ps=20.07 w=19.74 l=1.51
X10 VTAIL.t5 VP.t3 VDD1.t4 w_n2810_n4916# sky130_fd_pr__pfet_01v8 ad=3.2571 pd=20.07 as=3.2571 ps=20.07 w=19.74 l=1.51
X11 B.t5 B.t3 B.t4 w_n2810_n4916# sky130_fd_pr__pfet_01v8 ad=7.6986 pd=40.26 as=0 ps=0 w=19.74 l=1.51
X12 B.t2 B.t0 B.t1 w_n2810_n4916# sky130_fd_pr__pfet_01v8 ad=7.6986 pd=40.26 as=0 ps=0 w=19.74 l=1.51
X13 VDD1.t3 VP.t4 VTAIL.t0 w_n2810_n4916# sky130_fd_pr__pfet_01v8 ad=3.2571 pd=20.07 as=7.6986 ps=40.26 w=19.74 l=1.51
X14 VTAIL.t1 VP.t5 VDD1.t2 w_n2810_n4916# sky130_fd_pr__pfet_01v8 ad=7.6986 pd=40.26 as=3.2571 ps=20.07 w=19.74 l=1.51
X15 VDD2.t2 VN.t5 VTAIL.t10 w_n2810_n4916# sky130_fd_pr__pfet_01v8 ad=3.2571 pd=20.07 as=7.6986 ps=40.26 w=19.74 l=1.51
X16 VTAIL.t4 VP.t6 VDD1.t1 w_n2810_n4916# sky130_fd_pr__pfet_01v8 ad=3.2571 pd=20.07 as=3.2571 ps=20.07 w=19.74 l=1.51
X17 VTAIL.t13 VN.t6 VDD2.t1 w_n2810_n4916# sky130_fd_pr__pfet_01v8 ad=3.2571 pd=20.07 as=3.2571 ps=20.07 w=19.74 l=1.51
X18 VTAIL.t11 VN.t7 VDD2.t0 w_n2810_n4916# sky130_fd_pr__pfet_01v8 ad=7.6986 pd=40.26 as=3.2571 ps=20.07 w=19.74 l=1.51
X19 VDD1.t0 VP.t7 VTAIL.t3 w_n2810_n4916# sky130_fd_pr__pfet_01v8 ad=3.2571 pd=20.07 as=3.2571 ps=20.07 w=19.74 l=1.51
R0 VN.n5 VN.t1 350.332
R1 VN.n24 VN.t2 350.332
R2 VN.n4 VN.t0 315.057
R3 VN.n10 VN.t6 315.057
R4 VN.n17 VN.t5 315.057
R5 VN.n23 VN.t3 315.057
R6 VN.n29 VN.t4 315.057
R7 VN.n36 VN.t7 315.057
R8 VN.n18 VN.n17 173.105
R9 VN.n37 VN.n36 173.105
R10 VN.n35 VN.n19 161.3
R11 VN.n34 VN.n33 161.3
R12 VN.n32 VN.n20 161.3
R13 VN.n31 VN.n30 161.3
R14 VN.n28 VN.n21 161.3
R15 VN.n27 VN.n26 161.3
R16 VN.n25 VN.n22 161.3
R17 VN.n16 VN.n0 161.3
R18 VN.n15 VN.n14 161.3
R19 VN.n13 VN.n1 161.3
R20 VN.n12 VN.n11 161.3
R21 VN.n9 VN.n2 161.3
R22 VN.n8 VN.n7 161.3
R23 VN.n6 VN.n3 161.3
R24 VN.n15 VN.n1 56.0773
R25 VN.n34 VN.n20 56.0773
R26 VN VN.n37 52.01
R27 VN.n5 VN.n4 46.1603
R28 VN.n24 VN.n23 46.1603
R29 VN.n8 VN.n3 40.577
R30 VN.n9 VN.n8 40.577
R31 VN.n27 VN.n22 40.577
R32 VN.n28 VN.n27 40.577
R33 VN.n16 VN.n15 25.0767
R34 VN.n35 VN.n34 25.0767
R35 VN.n11 VN.n1 24.5923
R36 VN.n30 VN.n20 24.5923
R37 VN.n4 VN.n3 20.6576
R38 VN.n10 VN.n9 20.6576
R39 VN.n23 VN.n22 20.6576
R40 VN.n29 VN.n28 20.6576
R41 VN.n25 VN.n24 17.4856
R42 VN.n6 VN.n5 17.4856
R43 VN.n17 VN.n16 12.7883
R44 VN.n36 VN.n35 12.7883
R45 VN.n11 VN.n10 3.93519
R46 VN.n30 VN.n29 3.93519
R47 VN.n37 VN.n19 0.189894
R48 VN.n33 VN.n19 0.189894
R49 VN.n33 VN.n32 0.189894
R50 VN.n32 VN.n31 0.189894
R51 VN.n31 VN.n21 0.189894
R52 VN.n26 VN.n21 0.189894
R53 VN.n26 VN.n25 0.189894
R54 VN.n7 VN.n6 0.189894
R55 VN.n7 VN.n2 0.189894
R56 VN.n12 VN.n2 0.189894
R57 VN.n13 VN.n12 0.189894
R58 VN.n14 VN.n13 0.189894
R59 VN.n14 VN.n0 0.189894
R60 VN.n18 VN.n0 0.189894
R61 VN VN.n18 0.0516364
R62 VTAIL.n11 VTAIL.t1 53.8537
R63 VTAIL.n10 VTAIL.t8 53.8537
R64 VTAIL.n7 VTAIL.t11 53.8537
R65 VTAIL.n15 VTAIL.t10 53.8535
R66 VTAIL.n2 VTAIL.t14 53.8535
R67 VTAIL.n3 VTAIL.t0 53.8535
R68 VTAIL.n6 VTAIL.t6 53.8535
R69 VTAIL.n14 VTAIL.t2 53.8535
R70 VTAIL.n13 VTAIL.n12 52.207
R71 VTAIL.n9 VTAIL.n8 52.207
R72 VTAIL.n1 VTAIL.n0 52.2068
R73 VTAIL.n5 VTAIL.n4 52.2068
R74 VTAIL.n15 VTAIL.n14 30.9703
R75 VTAIL.n7 VTAIL.n6 30.9703
R76 VTAIL.n0 VTAIL.t15 1.64716
R77 VTAIL.n0 VTAIL.t13 1.64716
R78 VTAIL.n4 VTAIL.t7 1.64716
R79 VTAIL.n4 VTAIL.t5 1.64716
R80 VTAIL.n12 VTAIL.t3 1.64716
R81 VTAIL.n12 VTAIL.t4 1.64716
R82 VTAIL.n8 VTAIL.t12 1.64716
R83 VTAIL.n8 VTAIL.t9 1.64716
R84 VTAIL.n9 VTAIL.n7 1.58671
R85 VTAIL.n10 VTAIL.n9 1.58671
R86 VTAIL.n13 VTAIL.n11 1.58671
R87 VTAIL.n14 VTAIL.n13 1.58671
R88 VTAIL.n6 VTAIL.n5 1.58671
R89 VTAIL.n5 VTAIL.n3 1.58671
R90 VTAIL.n2 VTAIL.n1 1.58671
R91 VTAIL VTAIL.n15 1.52852
R92 VTAIL.n11 VTAIL.n10 0.470328
R93 VTAIL.n3 VTAIL.n2 0.470328
R94 VTAIL VTAIL.n1 0.0586897
R95 VDD2.n2 VDD2.n1 69.6234
R96 VDD2.n2 VDD2.n0 69.6234
R97 VDD2 VDD2.n5 69.6206
R98 VDD2.n4 VDD2.n3 68.8858
R99 VDD2.n4 VDD2.n2 47.8705
R100 VDD2.n5 VDD2.t4 1.64716
R101 VDD2.n5 VDD2.t5 1.64716
R102 VDD2.n3 VDD2.t0 1.64716
R103 VDD2.n3 VDD2.t3 1.64716
R104 VDD2.n1 VDD2.t1 1.64716
R105 VDD2.n1 VDD2.t2 1.64716
R106 VDD2.n0 VDD2.t6 1.64716
R107 VDD2.n0 VDD2.t7 1.64716
R108 VDD2 VDD2.n4 0.851793
R109 VP.n11 VP.t5 350.332
R110 VP.n25 VP.t1 315.057
R111 VP.n31 VP.t2 315.057
R112 VP.n38 VP.t3 315.057
R113 VP.n45 VP.t4 315.057
R114 VP.n23 VP.t0 315.057
R115 VP.n16 VP.t6 315.057
R116 VP.n10 VP.t7 315.057
R117 VP.n26 VP.n25 173.105
R118 VP.n46 VP.n45 173.105
R119 VP.n24 VP.n23 173.105
R120 VP.n12 VP.n9 161.3
R121 VP.n14 VP.n13 161.3
R122 VP.n15 VP.n8 161.3
R123 VP.n18 VP.n17 161.3
R124 VP.n19 VP.n7 161.3
R125 VP.n21 VP.n20 161.3
R126 VP.n22 VP.n6 161.3
R127 VP.n44 VP.n0 161.3
R128 VP.n43 VP.n42 161.3
R129 VP.n41 VP.n1 161.3
R130 VP.n40 VP.n39 161.3
R131 VP.n37 VP.n2 161.3
R132 VP.n36 VP.n35 161.3
R133 VP.n34 VP.n3 161.3
R134 VP.n33 VP.n32 161.3
R135 VP.n30 VP.n4 161.3
R136 VP.n29 VP.n28 161.3
R137 VP.n27 VP.n5 161.3
R138 VP.n30 VP.n29 56.0773
R139 VP.n43 VP.n1 56.0773
R140 VP.n21 VP.n7 56.0773
R141 VP.n26 VP.n24 51.6293
R142 VP.n11 VP.n10 46.1603
R143 VP.n36 VP.n3 40.577
R144 VP.n37 VP.n36 40.577
R145 VP.n15 VP.n14 40.577
R146 VP.n14 VP.n9 40.577
R147 VP.n29 VP.n5 25.0767
R148 VP.n44 VP.n43 25.0767
R149 VP.n22 VP.n21 25.0767
R150 VP.n32 VP.n30 24.5923
R151 VP.n39 VP.n1 24.5923
R152 VP.n17 VP.n7 24.5923
R153 VP.n31 VP.n3 20.6576
R154 VP.n38 VP.n37 20.6576
R155 VP.n16 VP.n15 20.6576
R156 VP.n10 VP.n9 20.6576
R157 VP.n12 VP.n11 17.4856
R158 VP.n25 VP.n5 12.7883
R159 VP.n45 VP.n44 12.7883
R160 VP.n23 VP.n22 12.7883
R161 VP.n32 VP.n31 3.93519
R162 VP.n39 VP.n38 3.93519
R163 VP.n17 VP.n16 3.93519
R164 VP.n13 VP.n12 0.189894
R165 VP.n13 VP.n8 0.189894
R166 VP.n18 VP.n8 0.189894
R167 VP.n19 VP.n18 0.189894
R168 VP.n20 VP.n19 0.189894
R169 VP.n20 VP.n6 0.189894
R170 VP.n24 VP.n6 0.189894
R171 VP.n27 VP.n26 0.189894
R172 VP.n28 VP.n27 0.189894
R173 VP.n28 VP.n4 0.189894
R174 VP.n33 VP.n4 0.189894
R175 VP.n34 VP.n33 0.189894
R176 VP.n35 VP.n34 0.189894
R177 VP.n35 VP.n2 0.189894
R178 VP.n40 VP.n2 0.189894
R179 VP.n41 VP.n40 0.189894
R180 VP.n42 VP.n41 0.189894
R181 VP.n42 VP.n0 0.189894
R182 VP.n46 VP.n0 0.189894
R183 VP VP.n46 0.0516364
R184 VDD1 VDD1.n0 69.7371
R185 VDD1.n3 VDD1.n2 69.6234
R186 VDD1.n3 VDD1.n1 69.6234
R187 VDD1.n5 VDD1.n4 68.8857
R188 VDD1.n5 VDD1.n3 48.4535
R189 VDD1.n4 VDD1.t1 1.64716
R190 VDD1.n4 VDD1.t7 1.64716
R191 VDD1.n0 VDD1.t2 1.64716
R192 VDD1.n0 VDD1.t0 1.64716
R193 VDD1.n2 VDD1.t4 1.64716
R194 VDD1.n2 VDD1.t3 1.64716
R195 VDD1.n1 VDD1.t6 1.64716
R196 VDD1.n1 VDD1.t5 1.64716
R197 VDD1 VDD1.n5 0.735414
R198 B.n586 B.n93 585
R199 B.n588 B.n587 585
R200 B.n589 B.n92 585
R201 B.n591 B.n590 585
R202 B.n592 B.n91 585
R203 B.n594 B.n593 585
R204 B.n595 B.n90 585
R205 B.n597 B.n596 585
R206 B.n598 B.n89 585
R207 B.n600 B.n599 585
R208 B.n601 B.n88 585
R209 B.n603 B.n602 585
R210 B.n604 B.n87 585
R211 B.n606 B.n605 585
R212 B.n607 B.n86 585
R213 B.n609 B.n608 585
R214 B.n610 B.n85 585
R215 B.n612 B.n611 585
R216 B.n613 B.n84 585
R217 B.n615 B.n614 585
R218 B.n616 B.n83 585
R219 B.n618 B.n617 585
R220 B.n619 B.n82 585
R221 B.n621 B.n620 585
R222 B.n622 B.n81 585
R223 B.n624 B.n623 585
R224 B.n625 B.n80 585
R225 B.n627 B.n626 585
R226 B.n628 B.n79 585
R227 B.n630 B.n629 585
R228 B.n631 B.n78 585
R229 B.n633 B.n632 585
R230 B.n634 B.n77 585
R231 B.n636 B.n635 585
R232 B.n637 B.n76 585
R233 B.n639 B.n638 585
R234 B.n640 B.n75 585
R235 B.n642 B.n641 585
R236 B.n643 B.n74 585
R237 B.n645 B.n644 585
R238 B.n646 B.n73 585
R239 B.n648 B.n647 585
R240 B.n649 B.n72 585
R241 B.n651 B.n650 585
R242 B.n652 B.n71 585
R243 B.n654 B.n653 585
R244 B.n655 B.n70 585
R245 B.n657 B.n656 585
R246 B.n658 B.n69 585
R247 B.n660 B.n659 585
R248 B.n661 B.n68 585
R249 B.n663 B.n662 585
R250 B.n664 B.n67 585
R251 B.n666 B.n665 585
R252 B.n667 B.n66 585
R253 B.n669 B.n668 585
R254 B.n670 B.n65 585
R255 B.n672 B.n671 585
R256 B.n673 B.n64 585
R257 B.n675 B.n674 585
R258 B.n676 B.n63 585
R259 B.n678 B.n677 585
R260 B.n679 B.n59 585
R261 B.n681 B.n680 585
R262 B.n682 B.n58 585
R263 B.n684 B.n683 585
R264 B.n685 B.n57 585
R265 B.n687 B.n686 585
R266 B.n688 B.n56 585
R267 B.n690 B.n689 585
R268 B.n691 B.n55 585
R269 B.n693 B.n692 585
R270 B.n694 B.n54 585
R271 B.n696 B.n695 585
R272 B.n698 B.n51 585
R273 B.n700 B.n699 585
R274 B.n701 B.n50 585
R275 B.n703 B.n702 585
R276 B.n704 B.n49 585
R277 B.n706 B.n705 585
R278 B.n707 B.n48 585
R279 B.n709 B.n708 585
R280 B.n710 B.n47 585
R281 B.n712 B.n711 585
R282 B.n713 B.n46 585
R283 B.n715 B.n714 585
R284 B.n716 B.n45 585
R285 B.n718 B.n717 585
R286 B.n719 B.n44 585
R287 B.n721 B.n720 585
R288 B.n722 B.n43 585
R289 B.n724 B.n723 585
R290 B.n725 B.n42 585
R291 B.n727 B.n726 585
R292 B.n728 B.n41 585
R293 B.n730 B.n729 585
R294 B.n731 B.n40 585
R295 B.n733 B.n732 585
R296 B.n734 B.n39 585
R297 B.n736 B.n735 585
R298 B.n737 B.n38 585
R299 B.n739 B.n738 585
R300 B.n740 B.n37 585
R301 B.n742 B.n741 585
R302 B.n743 B.n36 585
R303 B.n745 B.n744 585
R304 B.n746 B.n35 585
R305 B.n748 B.n747 585
R306 B.n749 B.n34 585
R307 B.n751 B.n750 585
R308 B.n752 B.n33 585
R309 B.n754 B.n753 585
R310 B.n755 B.n32 585
R311 B.n757 B.n756 585
R312 B.n758 B.n31 585
R313 B.n760 B.n759 585
R314 B.n761 B.n30 585
R315 B.n763 B.n762 585
R316 B.n764 B.n29 585
R317 B.n766 B.n765 585
R318 B.n767 B.n28 585
R319 B.n769 B.n768 585
R320 B.n770 B.n27 585
R321 B.n772 B.n771 585
R322 B.n773 B.n26 585
R323 B.n775 B.n774 585
R324 B.n776 B.n25 585
R325 B.n778 B.n777 585
R326 B.n779 B.n24 585
R327 B.n781 B.n780 585
R328 B.n782 B.n23 585
R329 B.n784 B.n783 585
R330 B.n785 B.n22 585
R331 B.n787 B.n786 585
R332 B.n788 B.n21 585
R333 B.n790 B.n789 585
R334 B.n791 B.n20 585
R335 B.n793 B.n792 585
R336 B.n585 B.n584 585
R337 B.n583 B.n94 585
R338 B.n582 B.n581 585
R339 B.n580 B.n95 585
R340 B.n579 B.n578 585
R341 B.n577 B.n96 585
R342 B.n576 B.n575 585
R343 B.n574 B.n97 585
R344 B.n573 B.n572 585
R345 B.n571 B.n98 585
R346 B.n570 B.n569 585
R347 B.n568 B.n99 585
R348 B.n567 B.n566 585
R349 B.n565 B.n100 585
R350 B.n564 B.n563 585
R351 B.n562 B.n101 585
R352 B.n561 B.n560 585
R353 B.n559 B.n102 585
R354 B.n558 B.n557 585
R355 B.n556 B.n103 585
R356 B.n555 B.n554 585
R357 B.n553 B.n104 585
R358 B.n552 B.n551 585
R359 B.n550 B.n105 585
R360 B.n549 B.n548 585
R361 B.n547 B.n106 585
R362 B.n546 B.n545 585
R363 B.n544 B.n107 585
R364 B.n543 B.n542 585
R365 B.n541 B.n108 585
R366 B.n540 B.n539 585
R367 B.n538 B.n109 585
R368 B.n537 B.n536 585
R369 B.n535 B.n110 585
R370 B.n534 B.n533 585
R371 B.n532 B.n111 585
R372 B.n531 B.n530 585
R373 B.n529 B.n112 585
R374 B.n528 B.n527 585
R375 B.n526 B.n113 585
R376 B.n525 B.n524 585
R377 B.n523 B.n114 585
R378 B.n522 B.n521 585
R379 B.n520 B.n115 585
R380 B.n519 B.n518 585
R381 B.n517 B.n116 585
R382 B.n516 B.n515 585
R383 B.n514 B.n117 585
R384 B.n513 B.n512 585
R385 B.n511 B.n118 585
R386 B.n510 B.n509 585
R387 B.n508 B.n119 585
R388 B.n507 B.n506 585
R389 B.n505 B.n120 585
R390 B.n504 B.n503 585
R391 B.n502 B.n121 585
R392 B.n501 B.n500 585
R393 B.n499 B.n122 585
R394 B.n498 B.n497 585
R395 B.n496 B.n123 585
R396 B.n495 B.n494 585
R397 B.n493 B.n124 585
R398 B.n492 B.n491 585
R399 B.n490 B.n125 585
R400 B.n489 B.n488 585
R401 B.n487 B.n126 585
R402 B.n486 B.n485 585
R403 B.n484 B.n127 585
R404 B.n483 B.n482 585
R405 B.n481 B.n128 585
R406 B.n480 B.n479 585
R407 B.n271 B.n202 585
R408 B.n273 B.n272 585
R409 B.n274 B.n201 585
R410 B.n276 B.n275 585
R411 B.n277 B.n200 585
R412 B.n279 B.n278 585
R413 B.n280 B.n199 585
R414 B.n282 B.n281 585
R415 B.n283 B.n198 585
R416 B.n285 B.n284 585
R417 B.n286 B.n197 585
R418 B.n288 B.n287 585
R419 B.n289 B.n196 585
R420 B.n291 B.n290 585
R421 B.n292 B.n195 585
R422 B.n294 B.n293 585
R423 B.n295 B.n194 585
R424 B.n297 B.n296 585
R425 B.n298 B.n193 585
R426 B.n300 B.n299 585
R427 B.n301 B.n192 585
R428 B.n303 B.n302 585
R429 B.n304 B.n191 585
R430 B.n306 B.n305 585
R431 B.n307 B.n190 585
R432 B.n309 B.n308 585
R433 B.n310 B.n189 585
R434 B.n312 B.n311 585
R435 B.n313 B.n188 585
R436 B.n315 B.n314 585
R437 B.n316 B.n187 585
R438 B.n318 B.n317 585
R439 B.n319 B.n186 585
R440 B.n321 B.n320 585
R441 B.n322 B.n185 585
R442 B.n324 B.n323 585
R443 B.n325 B.n184 585
R444 B.n327 B.n326 585
R445 B.n328 B.n183 585
R446 B.n330 B.n329 585
R447 B.n331 B.n182 585
R448 B.n333 B.n332 585
R449 B.n334 B.n181 585
R450 B.n336 B.n335 585
R451 B.n337 B.n180 585
R452 B.n339 B.n338 585
R453 B.n340 B.n179 585
R454 B.n342 B.n341 585
R455 B.n343 B.n178 585
R456 B.n345 B.n344 585
R457 B.n346 B.n177 585
R458 B.n348 B.n347 585
R459 B.n349 B.n176 585
R460 B.n351 B.n350 585
R461 B.n352 B.n175 585
R462 B.n354 B.n353 585
R463 B.n355 B.n174 585
R464 B.n357 B.n356 585
R465 B.n358 B.n173 585
R466 B.n360 B.n359 585
R467 B.n361 B.n172 585
R468 B.n363 B.n362 585
R469 B.n364 B.n171 585
R470 B.n366 B.n365 585
R471 B.n368 B.n168 585
R472 B.n370 B.n369 585
R473 B.n371 B.n167 585
R474 B.n373 B.n372 585
R475 B.n374 B.n166 585
R476 B.n376 B.n375 585
R477 B.n377 B.n165 585
R478 B.n379 B.n378 585
R479 B.n380 B.n164 585
R480 B.n382 B.n381 585
R481 B.n384 B.n383 585
R482 B.n385 B.n160 585
R483 B.n387 B.n386 585
R484 B.n388 B.n159 585
R485 B.n390 B.n389 585
R486 B.n391 B.n158 585
R487 B.n393 B.n392 585
R488 B.n394 B.n157 585
R489 B.n396 B.n395 585
R490 B.n397 B.n156 585
R491 B.n399 B.n398 585
R492 B.n400 B.n155 585
R493 B.n402 B.n401 585
R494 B.n403 B.n154 585
R495 B.n405 B.n404 585
R496 B.n406 B.n153 585
R497 B.n408 B.n407 585
R498 B.n409 B.n152 585
R499 B.n411 B.n410 585
R500 B.n412 B.n151 585
R501 B.n414 B.n413 585
R502 B.n415 B.n150 585
R503 B.n417 B.n416 585
R504 B.n418 B.n149 585
R505 B.n420 B.n419 585
R506 B.n421 B.n148 585
R507 B.n423 B.n422 585
R508 B.n424 B.n147 585
R509 B.n426 B.n425 585
R510 B.n427 B.n146 585
R511 B.n429 B.n428 585
R512 B.n430 B.n145 585
R513 B.n432 B.n431 585
R514 B.n433 B.n144 585
R515 B.n435 B.n434 585
R516 B.n436 B.n143 585
R517 B.n438 B.n437 585
R518 B.n439 B.n142 585
R519 B.n441 B.n440 585
R520 B.n442 B.n141 585
R521 B.n444 B.n443 585
R522 B.n445 B.n140 585
R523 B.n447 B.n446 585
R524 B.n448 B.n139 585
R525 B.n450 B.n449 585
R526 B.n451 B.n138 585
R527 B.n453 B.n452 585
R528 B.n454 B.n137 585
R529 B.n456 B.n455 585
R530 B.n457 B.n136 585
R531 B.n459 B.n458 585
R532 B.n460 B.n135 585
R533 B.n462 B.n461 585
R534 B.n463 B.n134 585
R535 B.n465 B.n464 585
R536 B.n466 B.n133 585
R537 B.n468 B.n467 585
R538 B.n469 B.n132 585
R539 B.n471 B.n470 585
R540 B.n472 B.n131 585
R541 B.n474 B.n473 585
R542 B.n475 B.n130 585
R543 B.n477 B.n476 585
R544 B.n478 B.n129 585
R545 B.n270 B.n269 585
R546 B.n268 B.n203 585
R547 B.n267 B.n266 585
R548 B.n265 B.n204 585
R549 B.n264 B.n263 585
R550 B.n262 B.n205 585
R551 B.n261 B.n260 585
R552 B.n259 B.n206 585
R553 B.n258 B.n257 585
R554 B.n256 B.n207 585
R555 B.n255 B.n254 585
R556 B.n253 B.n208 585
R557 B.n252 B.n251 585
R558 B.n250 B.n209 585
R559 B.n249 B.n248 585
R560 B.n247 B.n210 585
R561 B.n246 B.n245 585
R562 B.n244 B.n211 585
R563 B.n243 B.n242 585
R564 B.n241 B.n212 585
R565 B.n240 B.n239 585
R566 B.n238 B.n213 585
R567 B.n237 B.n236 585
R568 B.n235 B.n214 585
R569 B.n234 B.n233 585
R570 B.n232 B.n215 585
R571 B.n231 B.n230 585
R572 B.n229 B.n216 585
R573 B.n228 B.n227 585
R574 B.n226 B.n217 585
R575 B.n225 B.n224 585
R576 B.n223 B.n218 585
R577 B.n222 B.n221 585
R578 B.n220 B.n219 585
R579 B.n2 B.n0 585
R580 B.n845 B.n1 585
R581 B.n844 B.n843 585
R582 B.n842 B.n3 585
R583 B.n841 B.n840 585
R584 B.n839 B.n4 585
R585 B.n838 B.n837 585
R586 B.n836 B.n5 585
R587 B.n835 B.n834 585
R588 B.n833 B.n6 585
R589 B.n832 B.n831 585
R590 B.n830 B.n7 585
R591 B.n829 B.n828 585
R592 B.n827 B.n8 585
R593 B.n826 B.n825 585
R594 B.n824 B.n9 585
R595 B.n823 B.n822 585
R596 B.n821 B.n10 585
R597 B.n820 B.n819 585
R598 B.n818 B.n11 585
R599 B.n817 B.n816 585
R600 B.n815 B.n12 585
R601 B.n814 B.n813 585
R602 B.n812 B.n13 585
R603 B.n811 B.n810 585
R604 B.n809 B.n14 585
R605 B.n808 B.n807 585
R606 B.n806 B.n15 585
R607 B.n805 B.n804 585
R608 B.n803 B.n16 585
R609 B.n802 B.n801 585
R610 B.n800 B.n17 585
R611 B.n799 B.n798 585
R612 B.n797 B.n18 585
R613 B.n796 B.n795 585
R614 B.n794 B.n19 585
R615 B.n847 B.n846 585
R616 B.n269 B.n202 554.963
R617 B.n792 B.n19 554.963
R618 B.n479 B.n478 554.963
R619 B.n586 B.n585 554.963
R620 B.n161 B.t9 520.533
R621 B.n169 B.t0 520.533
R622 B.n52 B.t6 520.533
R623 B.n60 B.t3 520.533
R624 B.n269 B.n268 163.367
R625 B.n268 B.n267 163.367
R626 B.n267 B.n204 163.367
R627 B.n263 B.n204 163.367
R628 B.n263 B.n262 163.367
R629 B.n262 B.n261 163.367
R630 B.n261 B.n206 163.367
R631 B.n257 B.n206 163.367
R632 B.n257 B.n256 163.367
R633 B.n256 B.n255 163.367
R634 B.n255 B.n208 163.367
R635 B.n251 B.n208 163.367
R636 B.n251 B.n250 163.367
R637 B.n250 B.n249 163.367
R638 B.n249 B.n210 163.367
R639 B.n245 B.n210 163.367
R640 B.n245 B.n244 163.367
R641 B.n244 B.n243 163.367
R642 B.n243 B.n212 163.367
R643 B.n239 B.n212 163.367
R644 B.n239 B.n238 163.367
R645 B.n238 B.n237 163.367
R646 B.n237 B.n214 163.367
R647 B.n233 B.n214 163.367
R648 B.n233 B.n232 163.367
R649 B.n232 B.n231 163.367
R650 B.n231 B.n216 163.367
R651 B.n227 B.n216 163.367
R652 B.n227 B.n226 163.367
R653 B.n226 B.n225 163.367
R654 B.n225 B.n218 163.367
R655 B.n221 B.n218 163.367
R656 B.n221 B.n220 163.367
R657 B.n220 B.n2 163.367
R658 B.n846 B.n2 163.367
R659 B.n846 B.n845 163.367
R660 B.n845 B.n844 163.367
R661 B.n844 B.n3 163.367
R662 B.n840 B.n3 163.367
R663 B.n840 B.n839 163.367
R664 B.n839 B.n838 163.367
R665 B.n838 B.n5 163.367
R666 B.n834 B.n5 163.367
R667 B.n834 B.n833 163.367
R668 B.n833 B.n832 163.367
R669 B.n832 B.n7 163.367
R670 B.n828 B.n7 163.367
R671 B.n828 B.n827 163.367
R672 B.n827 B.n826 163.367
R673 B.n826 B.n9 163.367
R674 B.n822 B.n9 163.367
R675 B.n822 B.n821 163.367
R676 B.n821 B.n820 163.367
R677 B.n820 B.n11 163.367
R678 B.n816 B.n11 163.367
R679 B.n816 B.n815 163.367
R680 B.n815 B.n814 163.367
R681 B.n814 B.n13 163.367
R682 B.n810 B.n13 163.367
R683 B.n810 B.n809 163.367
R684 B.n809 B.n808 163.367
R685 B.n808 B.n15 163.367
R686 B.n804 B.n15 163.367
R687 B.n804 B.n803 163.367
R688 B.n803 B.n802 163.367
R689 B.n802 B.n17 163.367
R690 B.n798 B.n17 163.367
R691 B.n798 B.n797 163.367
R692 B.n797 B.n796 163.367
R693 B.n796 B.n19 163.367
R694 B.n273 B.n202 163.367
R695 B.n274 B.n273 163.367
R696 B.n275 B.n274 163.367
R697 B.n275 B.n200 163.367
R698 B.n279 B.n200 163.367
R699 B.n280 B.n279 163.367
R700 B.n281 B.n280 163.367
R701 B.n281 B.n198 163.367
R702 B.n285 B.n198 163.367
R703 B.n286 B.n285 163.367
R704 B.n287 B.n286 163.367
R705 B.n287 B.n196 163.367
R706 B.n291 B.n196 163.367
R707 B.n292 B.n291 163.367
R708 B.n293 B.n292 163.367
R709 B.n293 B.n194 163.367
R710 B.n297 B.n194 163.367
R711 B.n298 B.n297 163.367
R712 B.n299 B.n298 163.367
R713 B.n299 B.n192 163.367
R714 B.n303 B.n192 163.367
R715 B.n304 B.n303 163.367
R716 B.n305 B.n304 163.367
R717 B.n305 B.n190 163.367
R718 B.n309 B.n190 163.367
R719 B.n310 B.n309 163.367
R720 B.n311 B.n310 163.367
R721 B.n311 B.n188 163.367
R722 B.n315 B.n188 163.367
R723 B.n316 B.n315 163.367
R724 B.n317 B.n316 163.367
R725 B.n317 B.n186 163.367
R726 B.n321 B.n186 163.367
R727 B.n322 B.n321 163.367
R728 B.n323 B.n322 163.367
R729 B.n323 B.n184 163.367
R730 B.n327 B.n184 163.367
R731 B.n328 B.n327 163.367
R732 B.n329 B.n328 163.367
R733 B.n329 B.n182 163.367
R734 B.n333 B.n182 163.367
R735 B.n334 B.n333 163.367
R736 B.n335 B.n334 163.367
R737 B.n335 B.n180 163.367
R738 B.n339 B.n180 163.367
R739 B.n340 B.n339 163.367
R740 B.n341 B.n340 163.367
R741 B.n341 B.n178 163.367
R742 B.n345 B.n178 163.367
R743 B.n346 B.n345 163.367
R744 B.n347 B.n346 163.367
R745 B.n347 B.n176 163.367
R746 B.n351 B.n176 163.367
R747 B.n352 B.n351 163.367
R748 B.n353 B.n352 163.367
R749 B.n353 B.n174 163.367
R750 B.n357 B.n174 163.367
R751 B.n358 B.n357 163.367
R752 B.n359 B.n358 163.367
R753 B.n359 B.n172 163.367
R754 B.n363 B.n172 163.367
R755 B.n364 B.n363 163.367
R756 B.n365 B.n364 163.367
R757 B.n365 B.n168 163.367
R758 B.n370 B.n168 163.367
R759 B.n371 B.n370 163.367
R760 B.n372 B.n371 163.367
R761 B.n372 B.n166 163.367
R762 B.n376 B.n166 163.367
R763 B.n377 B.n376 163.367
R764 B.n378 B.n377 163.367
R765 B.n378 B.n164 163.367
R766 B.n382 B.n164 163.367
R767 B.n383 B.n382 163.367
R768 B.n383 B.n160 163.367
R769 B.n387 B.n160 163.367
R770 B.n388 B.n387 163.367
R771 B.n389 B.n388 163.367
R772 B.n389 B.n158 163.367
R773 B.n393 B.n158 163.367
R774 B.n394 B.n393 163.367
R775 B.n395 B.n394 163.367
R776 B.n395 B.n156 163.367
R777 B.n399 B.n156 163.367
R778 B.n400 B.n399 163.367
R779 B.n401 B.n400 163.367
R780 B.n401 B.n154 163.367
R781 B.n405 B.n154 163.367
R782 B.n406 B.n405 163.367
R783 B.n407 B.n406 163.367
R784 B.n407 B.n152 163.367
R785 B.n411 B.n152 163.367
R786 B.n412 B.n411 163.367
R787 B.n413 B.n412 163.367
R788 B.n413 B.n150 163.367
R789 B.n417 B.n150 163.367
R790 B.n418 B.n417 163.367
R791 B.n419 B.n418 163.367
R792 B.n419 B.n148 163.367
R793 B.n423 B.n148 163.367
R794 B.n424 B.n423 163.367
R795 B.n425 B.n424 163.367
R796 B.n425 B.n146 163.367
R797 B.n429 B.n146 163.367
R798 B.n430 B.n429 163.367
R799 B.n431 B.n430 163.367
R800 B.n431 B.n144 163.367
R801 B.n435 B.n144 163.367
R802 B.n436 B.n435 163.367
R803 B.n437 B.n436 163.367
R804 B.n437 B.n142 163.367
R805 B.n441 B.n142 163.367
R806 B.n442 B.n441 163.367
R807 B.n443 B.n442 163.367
R808 B.n443 B.n140 163.367
R809 B.n447 B.n140 163.367
R810 B.n448 B.n447 163.367
R811 B.n449 B.n448 163.367
R812 B.n449 B.n138 163.367
R813 B.n453 B.n138 163.367
R814 B.n454 B.n453 163.367
R815 B.n455 B.n454 163.367
R816 B.n455 B.n136 163.367
R817 B.n459 B.n136 163.367
R818 B.n460 B.n459 163.367
R819 B.n461 B.n460 163.367
R820 B.n461 B.n134 163.367
R821 B.n465 B.n134 163.367
R822 B.n466 B.n465 163.367
R823 B.n467 B.n466 163.367
R824 B.n467 B.n132 163.367
R825 B.n471 B.n132 163.367
R826 B.n472 B.n471 163.367
R827 B.n473 B.n472 163.367
R828 B.n473 B.n130 163.367
R829 B.n477 B.n130 163.367
R830 B.n478 B.n477 163.367
R831 B.n479 B.n128 163.367
R832 B.n483 B.n128 163.367
R833 B.n484 B.n483 163.367
R834 B.n485 B.n484 163.367
R835 B.n485 B.n126 163.367
R836 B.n489 B.n126 163.367
R837 B.n490 B.n489 163.367
R838 B.n491 B.n490 163.367
R839 B.n491 B.n124 163.367
R840 B.n495 B.n124 163.367
R841 B.n496 B.n495 163.367
R842 B.n497 B.n496 163.367
R843 B.n497 B.n122 163.367
R844 B.n501 B.n122 163.367
R845 B.n502 B.n501 163.367
R846 B.n503 B.n502 163.367
R847 B.n503 B.n120 163.367
R848 B.n507 B.n120 163.367
R849 B.n508 B.n507 163.367
R850 B.n509 B.n508 163.367
R851 B.n509 B.n118 163.367
R852 B.n513 B.n118 163.367
R853 B.n514 B.n513 163.367
R854 B.n515 B.n514 163.367
R855 B.n515 B.n116 163.367
R856 B.n519 B.n116 163.367
R857 B.n520 B.n519 163.367
R858 B.n521 B.n520 163.367
R859 B.n521 B.n114 163.367
R860 B.n525 B.n114 163.367
R861 B.n526 B.n525 163.367
R862 B.n527 B.n526 163.367
R863 B.n527 B.n112 163.367
R864 B.n531 B.n112 163.367
R865 B.n532 B.n531 163.367
R866 B.n533 B.n532 163.367
R867 B.n533 B.n110 163.367
R868 B.n537 B.n110 163.367
R869 B.n538 B.n537 163.367
R870 B.n539 B.n538 163.367
R871 B.n539 B.n108 163.367
R872 B.n543 B.n108 163.367
R873 B.n544 B.n543 163.367
R874 B.n545 B.n544 163.367
R875 B.n545 B.n106 163.367
R876 B.n549 B.n106 163.367
R877 B.n550 B.n549 163.367
R878 B.n551 B.n550 163.367
R879 B.n551 B.n104 163.367
R880 B.n555 B.n104 163.367
R881 B.n556 B.n555 163.367
R882 B.n557 B.n556 163.367
R883 B.n557 B.n102 163.367
R884 B.n561 B.n102 163.367
R885 B.n562 B.n561 163.367
R886 B.n563 B.n562 163.367
R887 B.n563 B.n100 163.367
R888 B.n567 B.n100 163.367
R889 B.n568 B.n567 163.367
R890 B.n569 B.n568 163.367
R891 B.n569 B.n98 163.367
R892 B.n573 B.n98 163.367
R893 B.n574 B.n573 163.367
R894 B.n575 B.n574 163.367
R895 B.n575 B.n96 163.367
R896 B.n579 B.n96 163.367
R897 B.n580 B.n579 163.367
R898 B.n581 B.n580 163.367
R899 B.n581 B.n94 163.367
R900 B.n585 B.n94 163.367
R901 B.n792 B.n791 163.367
R902 B.n791 B.n790 163.367
R903 B.n790 B.n21 163.367
R904 B.n786 B.n21 163.367
R905 B.n786 B.n785 163.367
R906 B.n785 B.n784 163.367
R907 B.n784 B.n23 163.367
R908 B.n780 B.n23 163.367
R909 B.n780 B.n779 163.367
R910 B.n779 B.n778 163.367
R911 B.n778 B.n25 163.367
R912 B.n774 B.n25 163.367
R913 B.n774 B.n773 163.367
R914 B.n773 B.n772 163.367
R915 B.n772 B.n27 163.367
R916 B.n768 B.n27 163.367
R917 B.n768 B.n767 163.367
R918 B.n767 B.n766 163.367
R919 B.n766 B.n29 163.367
R920 B.n762 B.n29 163.367
R921 B.n762 B.n761 163.367
R922 B.n761 B.n760 163.367
R923 B.n760 B.n31 163.367
R924 B.n756 B.n31 163.367
R925 B.n756 B.n755 163.367
R926 B.n755 B.n754 163.367
R927 B.n754 B.n33 163.367
R928 B.n750 B.n33 163.367
R929 B.n750 B.n749 163.367
R930 B.n749 B.n748 163.367
R931 B.n748 B.n35 163.367
R932 B.n744 B.n35 163.367
R933 B.n744 B.n743 163.367
R934 B.n743 B.n742 163.367
R935 B.n742 B.n37 163.367
R936 B.n738 B.n37 163.367
R937 B.n738 B.n737 163.367
R938 B.n737 B.n736 163.367
R939 B.n736 B.n39 163.367
R940 B.n732 B.n39 163.367
R941 B.n732 B.n731 163.367
R942 B.n731 B.n730 163.367
R943 B.n730 B.n41 163.367
R944 B.n726 B.n41 163.367
R945 B.n726 B.n725 163.367
R946 B.n725 B.n724 163.367
R947 B.n724 B.n43 163.367
R948 B.n720 B.n43 163.367
R949 B.n720 B.n719 163.367
R950 B.n719 B.n718 163.367
R951 B.n718 B.n45 163.367
R952 B.n714 B.n45 163.367
R953 B.n714 B.n713 163.367
R954 B.n713 B.n712 163.367
R955 B.n712 B.n47 163.367
R956 B.n708 B.n47 163.367
R957 B.n708 B.n707 163.367
R958 B.n707 B.n706 163.367
R959 B.n706 B.n49 163.367
R960 B.n702 B.n49 163.367
R961 B.n702 B.n701 163.367
R962 B.n701 B.n700 163.367
R963 B.n700 B.n51 163.367
R964 B.n695 B.n51 163.367
R965 B.n695 B.n694 163.367
R966 B.n694 B.n693 163.367
R967 B.n693 B.n55 163.367
R968 B.n689 B.n55 163.367
R969 B.n689 B.n688 163.367
R970 B.n688 B.n687 163.367
R971 B.n687 B.n57 163.367
R972 B.n683 B.n57 163.367
R973 B.n683 B.n682 163.367
R974 B.n682 B.n681 163.367
R975 B.n681 B.n59 163.367
R976 B.n677 B.n59 163.367
R977 B.n677 B.n676 163.367
R978 B.n676 B.n675 163.367
R979 B.n675 B.n64 163.367
R980 B.n671 B.n64 163.367
R981 B.n671 B.n670 163.367
R982 B.n670 B.n669 163.367
R983 B.n669 B.n66 163.367
R984 B.n665 B.n66 163.367
R985 B.n665 B.n664 163.367
R986 B.n664 B.n663 163.367
R987 B.n663 B.n68 163.367
R988 B.n659 B.n68 163.367
R989 B.n659 B.n658 163.367
R990 B.n658 B.n657 163.367
R991 B.n657 B.n70 163.367
R992 B.n653 B.n70 163.367
R993 B.n653 B.n652 163.367
R994 B.n652 B.n651 163.367
R995 B.n651 B.n72 163.367
R996 B.n647 B.n72 163.367
R997 B.n647 B.n646 163.367
R998 B.n646 B.n645 163.367
R999 B.n645 B.n74 163.367
R1000 B.n641 B.n74 163.367
R1001 B.n641 B.n640 163.367
R1002 B.n640 B.n639 163.367
R1003 B.n639 B.n76 163.367
R1004 B.n635 B.n76 163.367
R1005 B.n635 B.n634 163.367
R1006 B.n634 B.n633 163.367
R1007 B.n633 B.n78 163.367
R1008 B.n629 B.n78 163.367
R1009 B.n629 B.n628 163.367
R1010 B.n628 B.n627 163.367
R1011 B.n627 B.n80 163.367
R1012 B.n623 B.n80 163.367
R1013 B.n623 B.n622 163.367
R1014 B.n622 B.n621 163.367
R1015 B.n621 B.n82 163.367
R1016 B.n617 B.n82 163.367
R1017 B.n617 B.n616 163.367
R1018 B.n616 B.n615 163.367
R1019 B.n615 B.n84 163.367
R1020 B.n611 B.n84 163.367
R1021 B.n611 B.n610 163.367
R1022 B.n610 B.n609 163.367
R1023 B.n609 B.n86 163.367
R1024 B.n605 B.n86 163.367
R1025 B.n605 B.n604 163.367
R1026 B.n604 B.n603 163.367
R1027 B.n603 B.n88 163.367
R1028 B.n599 B.n88 163.367
R1029 B.n599 B.n598 163.367
R1030 B.n598 B.n597 163.367
R1031 B.n597 B.n90 163.367
R1032 B.n593 B.n90 163.367
R1033 B.n593 B.n592 163.367
R1034 B.n592 B.n591 163.367
R1035 B.n591 B.n92 163.367
R1036 B.n587 B.n92 163.367
R1037 B.n587 B.n586 163.367
R1038 B.n161 B.t11 142.12
R1039 B.n60 B.t4 142.12
R1040 B.n169 B.t2 142.095
R1041 B.n52 B.t7 142.095
R1042 B.n162 B.t10 106.436
R1043 B.n61 B.t5 106.436
R1044 B.n170 B.t1 106.409
R1045 B.n53 B.t8 106.409
R1046 B.n163 B.n162 59.5399
R1047 B.n367 B.n170 59.5399
R1048 B.n697 B.n53 59.5399
R1049 B.n62 B.n61 59.5399
R1050 B.n794 B.n793 36.059
R1051 B.n584 B.n93 36.059
R1052 B.n480 B.n129 36.059
R1053 B.n271 B.n270 36.059
R1054 B.n162 B.n161 35.6853
R1055 B.n170 B.n169 35.6853
R1056 B.n53 B.n52 35.6853
R1057 B.n61 B.n60 35.6853
R1058 B B.n847 18.0485
R1059 B.n793 B.n20 10.6151
R1060 B.n789 B.n20 10.6151
R1061 B.n789 B.n788 10.6151
R1062 B.n788 B.n787 10.6151
R1063 B.n787 B.n22 10.6151
R1064 B.n783 B.n22 10.6151
R1065 B.n783 B.n782 10.6151
R1066 B.n782 B.n781 10.6151
R1067 B.n781 B.n24 10.6151
R1068 B.n777 B.n24 10.6151
R1069 B.n777 B.n776 10.6151
R1070 B.n776 B.n775 10.6151
R1071 B.n775 B.n26 10.6151
R1072 B.n771 B.n26 10.6151
R1073 B.n771 B.n770 10.6151
R1074 B.n770 B.n769 10.6151
R1075 B.n769 B.n28 10.6151
R1076 B.n765 B.n28 10.6151
R1077 B.n765 B.n764 10.6151
R1078 B.n764 B.n763 10.6151
R1079 B.n763 B.n30 10.6151
R1080 B.n759 B.n30 10.6151
R1081 B.n759 B.n758 10.6151
R1082 B.n758 B.n757 10.6151
R1083 B.n757 B.n32 10.6151
R1084 B.n753 B.n32 10.6151
R1085 B.n753 B.n752 10.6151
R1086 B.n752 B.n751 10.6151
R1087 B.n751 B.n34 10.6151
R1088 B.n747 B.n34 10.6151
R1089 B.n747 B.n746 10.6151
R1090 B.n746 B.n745 10.6151
R1091 B.n745 B.n36 10.6151
R1092 B.n741 B.n36 10.6151
R1093 B.n741 B.n740 10.6151
R1094 B.n740 B.n739 10.6151
R1095 B.n739 B.n38 10.6151
R1096 B.n735 B.n38 10.6151
R1097 B.n735 B.n734 10.6151
R1098 B.n734 B.n733 10.6151
R1099 B.n733 B.n40 10.6151
R1100 B.n729 B.n40 10.6151
R1101 B.n729 B.n728 10.6151
R1102 B.n728 B.n727 10.6151
R1103 B.n727 B.n42 10.6151
R1104 B.n723 B.n42 10.6151
R1105 B.n723 B.n722 10.6151
R1106 B.n722 B.n721 10.6151
R1107 B.n721 B.n44 10.6151
R1108 B.n717 B.n44 10.6151
R1109 B.n717 B.n716 10.6151
R1110 B.n716 B.n715 10.6151
R1111 B.n715 B.n46 10.6151
R1112 B.n711 B.n46 10.6151
R1113 B.n711 B.n710 10.6151
R1114 B.n710 B.n709 10.6151
R1115 B.n709 B.n48 10.6151
R1116 B.n705 B.n48 10.6151
R1117 B.n705 B.n704 10.6151
R1118 B.n704 B.n703 10.6151
R1119 B.n703 B.n50 10.6151
R1120 B.n699 B.n50 10.6151
R1121 B.n699 B.n698 10.6151
R1122 B.n696 B.n54 10.6151
R1123 B.n692 B.n54 10.6151
R1124 B.n692 B.n691 10.6151
R1125 B.n691 B.n690 10.6151
R1126 B.n690 B.n56 10.6151
R1127 B.n686 B.n56 10.6151
R1128 B.n686 B.n685 10.6151
R1129 B.n685 B.n684 10.6151
R1130 B.n684 B.n58 10.6151
R1131 B.n680 B.n679 10.6151
R1132 B.n679 B.n678 10.6151
R1133 B.n678 B.n63 10.6151
R1134 B.n674 B.n63 10.6151
R1135 B.n674 B.n673 10.6151
R1136 B.n673 B.n672 10.6151
R1137 B.n672 B.n65 10.6151
R1138 B.n668 B.n65 10.6151
R1139 B.n668 B.n667 10.6151
R1140 B.n667 B.n666 10.6151
R1141 B.n666 B.n67 10.6151
R1142 B.n662 B.n67 10.6151
R1143 B.n662 B.n661 10.6151
R1144 B.n661 B.n660 10.6151
R1145 B.n660 B.n69 10.6151
R1146 B.n656 B.n69 10.6151
R1147 B.n656 B.n655 10.6151
R1148 B.n655 B.n654 10.6151
R1149 B.n654 B.n71 10.6151
R1150 B.n650 B.n71 10.6151
R1151 B.n650 B.n649 10.6151
R1152 B.n649 B.n648 10.6151
R1153 B.n648 B.n73 10.6151
R1154 B.n644 B.n73 10.6151
R1155 B.n644 B.n643 10.6151
R1156 B.n643 B.n642 10.6151
R1157 B.n642 B.n75 10.6151
R1158 B.n638 B.n75 10.6151
R1159 B.n638 B.n637 10.6151
R1160 B.n637 B.n636 10.6151
R1161 B.n636 B.n77 10.6151
R1162 B.n632 B.n77 10.6151
R1163 B.n632 B.n631 10.6151
R1164 B.n631 B.n630 10.6151
R1165 B.n630 B.n79 10.6151
R1166 B.n626 B.n79 10.6151
R1167 B.n626 B.n625 10.6151
R1168 B.n625 B.n624 10.6151
R1169 B.n624 B.n81 10.6151
R1170 B.n620 B.n81 10.6151
R1171 B.n620 B.n619 10.6151
R1172 B.n619 B.n618 10.6151
R1173 B.n618 B.n83 10.6151
R1174 B.n614 B.n83 10.6151
R1175 B.n614 B.n613 10.6151
R1176 B.n613 B.n612 10.6151
R1177 B.n612 B.n85 10.6151
R1178 B.n608 B.n85 10.6151
R1179 B.n608 B.n607 10.6151
R1180 B.n607 B.n606 10.6151
R1181 B.n606 B.n87 10.6151
R1182 B.n602 B.n87 10.6151
R1183 B.n602 B.n601 10.6151
R1184 B.n601 B.n600 10.6151
R1185 B.n600 B.n89 10.6151
R1186 B.n596 B.n89 10.6151
R1187 B.n596 B.n595 10.6151
R1188 B.n595 B.n594 10.6151
R1189 B.n594 B.n91 10.6151
R1190 B.n590 B.n91 10.6151
R1191 B.n590 B.n589 10.6151
R1192 B.n589 B.n588 10.6151
R1193 B.n588 B.n93 10.6151
R1194 B.n481 B.n480 10.6151
R1195 B.n482 B.n481 10.6151
R1196 B.n482 B.n127 10.6151
R1197 B.n486 B.n127 10.6151
R1198 B.n487 B.n486 10.6151
R1199 B.n488 B.n487 10.6151
R1200 B.n488 B.n125 10.6151
R1201 B.n492 B.n125 10.6151
R1202 B.n493 B.n492 10.6151
R1203 B.n494 B.n493 10.6151
R1204 B.n494 B.n123 10.6151
R1205 B.n498 B.n123 10.6151
R1206 B.n499 B.n498 10.6151
R1207 B.n500 B.n499 10.6151
R1208 B.n500 B.n121 10.6151
R1209 B.n504 B.n121 10.6151
R1210 B.n505 B.n504 10.6151
R1211 B.n506 B.n505 10.6151
R1212 B.n506 B.n119 10.6151
R1213 B.n510 B.n119 10.6151
R1214 B.n511 B.n510 10.6151
R1215 B.n512 B.n511 10.6151
R1216 B.n512 B.n117 10.6151
R1217 B.n516 B.n117 10.6151
R1218 B.n517 B.n516 10.6151
R1219 B.n518 B.n517 10.6151
R1220 B.n518 B.n115 10.6151
R1221 B.n522 B.n115 10.6151
R1222 B.n523 B.n522 10.6151
R1223 B.n524 B.n523 10.6151
R1224 B.n524 B.n113 10.6151
R1225 B.n528 B.n113 10.6151
R1226 B.n529 B.n528 10.6151
R1227 B.n530 B.n529 10.6151
R1228 B.n530 B.n111 10.6151
R1229 B.n534 B.n111 10.6151
R1230 B.n535 B.n534 10.6151
R1231 B.n536 B.n535 10.6151
R1232 B.n536 B.n109 10.6151
R1233 B.n540 B.n109 10.6151
R1234 B.n541 B.n540 10.6151
R1235 B.n542 B.n541 10.6151
R1236 B.n542 B.n107 10.6151
R1237 B.n546 B.n107 10.6151
R1238 B.n547 B.n546 10.6151
R1239 B.n548 B.n547 10.6151
R1240 B.n548 B.n105 10.6151
R1241 B.n552 B.n105 10.6151
R1242 B.n553 B.n552 10.6151
R1243 B.n554 B.n553 10.6151
R1244 B.n554 B.n103 10.6151
R1245 B.n558 B.n103 10.6151
R1246 B.n559 B.n558 10.6151
R1247 B.n560 B.n559 10.6151
R1248 B.n560 B.n101 10.6151
R1249 B.n564 B.n101 10.6151
R1250 B.n565 B.n564 10.6151
R1251 B.n566 B.n565 10.6151
R1252 B.n566 B.n99 10.6151
R1253 B.n570 B.n99 10.6151
R1254 B.n571 B.n570 10.6151
R1255 B.n572 B.n571 10.6151
R1256 B.n572 B.n97 10.6151
R1257 B.n576 B.n97 10.6151
R1258 B.n577 B.n576 10.6151
R1259 B.n578 B.n577 10.6151
R1260 B.n578 B.n95 10.6151
R1261 B.n582 B.n95 10.6151
R1262 B.n583 B.n582 10.6151
R1263 B.n584 B.n583 10.6151
R1264 B.n272 B.n271 10.6151
R1265 B.n272 B.n201 10.6151
R1266 B.n276 B.n201 10.6151
R1267 B.n277 B.n276 10.6151
R1268 B.n278 B.n277 10.6151
R1269 B.n278 B.n199 10.6151
R1270 B.n282 B.n199 10.6151
R1271 B.n283 B.n282 10.6151
R1272 B.n284 B.n283 10.6151
R1273 B.n284 B.n197 10.6151
R1274 B.n288 B.n197 10.6151
R1275 B.n289 B.n288 10.6151
R1276 B.n290 B.n289 10.6151
R1277 B.n290 B.n195 10.6151
R1278 B.n294 B.n195 10.6151
R1279 B.n295 B.n294 10.6151
R1280 B.n296 B.n295 10.6151
R1281 B.n296 B.n193 10.6151
R1282 B.n300 B.n193 10.6151
R1283 B.n301 B.n300 10.6151
R1284 B.n302 B.n301 10.6151
R1285 B.n302 B.n191 10.6151
R1286 B.n306 B.n191 10.6151
R1287 B.n307 B.n306 10.6151
R1288 B.n308 B.n307 10.6151
R1289 B.n308 B.n189 10.6151
R1290 B.n312 B.n189 10.6151
R1291 B.n313 B.n312 10.6151
R1292 B.n314 B.n313 10.6151
R1293 B.n314 B.n187 10.6151
R1294 B.n318 B.n187 10.6151
R1295 B.n319 B.n318 10.6151
R1296 B.n320 B.n319 10.6151
R1297 B.n320 B.n185 10.6151
R1298 B.n324 B.n185 10.6151
R1299 B.n325 B.n324 10.6151
R1300 B.n326 B.n325 10.6151
R1301 B.n326 B.n183 10.6151
R1302 B.n330 B.n183 10.6151
R1303 B.n331 B.n330 10.6151
R1304 B.n332 B.n331 10.6151
R1305 B.n332 B.n181 10.6151
R1306 B.n336 B.n181 10.6151
R1307 B.n337 B.n336 10.6151
R1308 B.n338 B.n337 10.6151
R1309 B.n338 B.n179 10.6151
R1310 B.n342 B.n179 10.6151
R1311 B.n343 B.n342 10.6151
R1312 B.n344 B.n343 10.6151
R1313 B.n344 B.n177 10.6151
R1314 B.n348 B.n177 10.6151
R1315 B.n349 B.n348 10.6151
R1316 B.n350 B.n349 10.6151
R1317 B.n350 B.n175 10.6151
R1318 B.n354 B.n175 10.6151
R1319 B.n355 B.n354 10.6151
R1320 B.n356 B.n355 10.6151
R1321 B.n356 B.n173 10.6151
R1322 B.n360 B.n173 10.6151
R1323 B.n361 B.n360 10.6151
R1324 B.n362 B.n361 10.6151
R1325 B.n362 B.n171 10.6151
R1326 B.n366 B.n171 10.6151
R1327 B.n369 B.n368 10.6151
R1328 B.n369 B.n167 10.6151
R1329 B.n373 B.n167 10.6151
R1330 B.n374 B.n373 10.6151
R1331 B.n375 B.n374 10.6151
R1332 B.n375 B.n165 10.6151
R1333 B.n379 B.n165 10.6151
R1334 B.n380 B.n379 10.6151
R1335 B.n381 B.n380 10.6151
R1336 B.n385 B.n384 10.6151
R1337 B.n386 B.n385 10.6151
R1338 B.n386 B.n159 10.6151
R1339 B.n390 B.n159 10.6151
R1340 B.n391 B.n390 10.6151
R1341 B.n392 B.n391 10.6151
R1342 B.n392 B.n157 10.6151
R1343 B.n396 B.n157 10.6151
R1344 B.n397 B.n396 10.6151
R1345 B.n398 B.n397 10.6151
R1346 B.n398 B.n155 10.6151
R1347 B.n402 B.n155 10.6151
R1348 B.n403 B.n402 10.6151
R1349 B.n404 B.n403 10.6151
R1350 B.n404 B.n153 10.6151
R1351 B.n408 B.n153 10.6151
R1352 B.n409 B.n408 10.6151
R1353 B.n410 B.n409 10.6151
R1354 B.n410 B.n151 10.6151
R1355 B.n414 B.n151 10.6151
R1356 B.n415 B.n414 10.6151
R1357 B.n416 B.n415 10.6151
R1358 B.n416 B.n149 10.6151
R1359 B.n420 B.n149 10.6151
R1360 B.n421 B.n420 10.6151
R1361 B.n422 B.n421 10.6151
R1362 B.n422 B.n147 10.6151
R1363 B.n426 B.n147 10.6151
R1364 B.n427 B.n426 10.6151
R1365 B.n428 B.n427 10.6151
R1366 B.n428 B.n145 10.6151
R1367 B.n432 B.n145 10.6151
R1368 B.n433 B.n432 10.6151
R1369 B.n434 B.n433 10.6151
R1370 B.n434 B.n143 10.6151
R1371 B.n438 B.n143 10.6151
R1372 B.n439 B.n438 10.6151
R1373 B.n440 B.n439 10.6151
R1374 B.n440 B.n141 10.6151
R1375 B.n444 B.n141 10.6151
R1376 B.n445 B.n444 10.6151
R1377 B.n446 B.n445 10.6151
R1378 B.n446 B.n139 10.6151
R1379 B.n450 B.n139 10.6151
R1380 B.n451 B.n450 10.6151
R1381 B.n452 B.n451 10.6151
R1382 B.n452 B.n137 10.6151
R1383 B.n456 B.n137 10.6151
R1384 B.n457 B.n456 10.6151
R1385 B.n458 B.n457 10.6151
R1386 B.n458 B.n135 10.6151
R1387 B.n462 B.n135 10.6151
R1388 B.n463 B.n462 10.6151
R1389 B.n464 B.n463 10.6151
R1390 B.n464 B.n133 10.6151
R1391 B.n468 B.n133 10.6151
R1392 B.n469 B.n468 10.6151
R1393 B.n470 B.n469 10.6151
R1394 B.n470 B.n131 10.6151
R1395 B.n474 B.n131 10.6151
R1396 B.n475 B.n474 10.6151
R1397 B.n476 B.n475 10.6151
R1398 B.n476 B.n129 10.6151
R1399 B.n270 B.n203 10.6151
R1400 B.n266 B.n203 10.6151
R1401 B.n266 B.n265 10.6151
R1402 B.n265 B.n264 10.6151
R1403 B.n264 B.n205 10.6151
R1404 B.n260 B.n205 10.6151
R1405 B.n260 B.n259 10.6151
R1406 B.n259 B.n258 10.6151
R1407 B.n258 B.n207 10.6151
R1408 B.n254 B.n207 10.6151
R1409 B.n254 B.n253 10.6151
R1410 B.n253 B.n252 10.6151
R1411 B.n252 B.n209 10.6151
R1412 B.n248 B.n209 10.6151
R1413 B.n248 B.n247 10.6151
R1414 B.n247 B.n246 10.6151
R1415 B.n246 B.n211 10.6151
R1416 B.n242 B.n211 10.6151
R1417 B.n242 B.n241 10.6151
R1418 B.n241 B.n240 10.6151
R1419 B.n240 B.n213 10.6151
R1420 B.n236 B.n213 10.6151
R1421 B.n236 B.n235 10.6151
R1422 B.n235 B.n234 10.6151
R1423 B.n234 B.n215 10.6151
R1424 B.n230 B.n215 10.6151
R1425 B.n230 B.n229 10.6151
R1426 B.n229 B.n228 10.6151
R1427 B.n228 B.n217 10.6151
R1428 B.n224 B.n217 10.6151
R1429 B.n224 B.n223 10.6151
R1430 B.n223 B.n222 10.6151
R1431 B.n222 B.n219 10.6151
R1432 B.n219 B.n0 10.6151
R1433 B.n843 B.n1 10.6151
R1434 B.n843 B.n842 10.6151
R1435 B.n842 B.n841 10.6151
R1436 B.n841 B.n4 10.6151
R1437 B.n837 B.n4 10.6151
R1438 B.n837 B.n836 10.6151
R1439 B.n836 B.n835 10.6151
R1440 B.n835 B.n6 10.6151
R1441 B.n831 B.n6 10.6151
R1442 B.n831 B.n830 10.6151
R1443 B.n830 B.n829 10.6151
R1444 B.n829 B.n8 10.6151
R1445 B.n825 B.n8 10.6151
R1446 B.n825 B.n824 10.6151
R1447 B.n824 B.n823 10.6151
R1448 B.n823 B.n10 10.6151
R1449 B.n819 B.n10 10.6151
R1450 B.n819 B.n818 10.6151
R1451 B.n818 B.n817 10.6151
R1452 B.n817 B.n12 10.6151
R1453 B.n813 B.n12 10.6151
R1454 B.n813 B.n812 10.6151
R1455 B.n812 B.n811 10.6151
R1456 B.n811 B.n14 10.6151
R1457 B.n807 B.n14 10.6151
R1458 B.n807 B.n806 10.6151
R1459 B.n806 B.n805 10.6151
R1460 B.n805 B.n16 10.6151
R1461 B.n801 B.n16 10.6151
R1462 B.n801 B.n800 10.6151
R1463 B.n800 B.n799 10.6151
R1464 B.n799 B.n18 10.6151
R1465 B.n795 B.n18 10.6151
R1466 B.n795 B.n794 10.6151
R1467 B.n698 B.n697 9.36635
R1468 B.n680 B.n62 9.36635
R1469 B.n367 B.n366 9.36635
R1470 B.n384 B.n163 9.36635
R1471 B.n847 B.n0 2.81026
R1472 B.n847 B.n1 2.81026
R1473 B.n697 B.n696 1.24928
R1474 B.n62 B.n58 1.24928
R1475 B.n368 B.n367 1.24928
R1476 B.n381 B.n163 1.24928
C0 VDD1 VN 0.150123f
C1 VP VN 7.756259f
C2 VDD1 VDD2 1.22582f
C3 VN w_n2810_n4916# 5.54681f
C4 VDD2 VP 0.404049f
C5 VDD2 w_n2810_n4916# 1.87306f
C6 VN B 1.06525f
C7 VDD2 B 1.58784f
C8 VDD1 VTAIL 12.026401f
C9 VTAIL VP 11.9533f
C10 VTAIL w_n2810_n4916# 5.97444f
C11 VDD2 VN 12.198099f
C12 VTAIL B 6.74074f
C13 VDD1 VP 12.4512f
C14 VDD1 w_n2810_n4916# 1.80406f
C15 VP w_n2810_n4916# 5.9084f
C16 VTAIL VN 11.9392f
C17 VDD1 B 1.52607f
C18 VP B 1.66558f
C19 VDD2 VTAIL 12.0735f
C20 w_n2810_n4916# B 10.6159f
C21 VDD2 VSUBS 1.701976f
C22 VDD1 VSUBS 2.152258f
C23 VTAIL VSUBS 1.470678f
C24 VN VSUBS 5.85426f
C25 VP VSUBS 2.748576f
C26 B VSUBS 4.440797f
C27 w_n2810_n4916# VSUBS 0.168701p
C28 B.n0 VSUBS 0.00425f
C29 B.n1 VSUBS 0.00425f
C30 B.n2 VSUBS 0.006721f
C31 B.n3 VSUBS 0.006721f
C32 B.n4 VSUBS 0.006721f
C33 B.n5 VSUBS 0.006721f
C34 B.n6 VSUBS 0.006721f
C35 B.n7 VSUBS 0.006721f
C36 B.n8 VSUBS 0.006721f
C37 B.n9 VSUBS 0.006721f
C38 B.n10 VSUBS 0.006721f
C39 B.n11 VSUBS 0.006721f
C40 B.n12 VSUBS 0.006721f
C41 B.n13 VSUBS 0.006721f
C42 B.n14 VSUBS 0.006721f
C43 B.n15 VSUBS 0.006721f
C44 B.n16 VSUBS 0.006721f
C45 B.n17 VSUBS 0.006721f
C46 B.n18 VSUBS 0.006721f
C47 B.n19 VSUBS 0.01646f
C48 B.n20 VSUBS 0.006721f
C49 B.n21 VSUBS 0.006721f
C50 B.n22 VSUBS 0.006721f
C51 B.n23 VSUBS 0.006721f
C52 B.n24 VSUBS 0.006721f
C53 B.n25 VSUBS 0.006721f
C54 B.n26 VSUBS 0.006721f
C55 B.n27 VSUBS 0.006721f
C56 B.n28 VSUBS 0.006721f
C57 B.n29 VSUBS 0.006721f
C58 B.n30 VSUBS 0.006721f
C59 B.n31 VSUBS 0.006721f
C60 B.n32 VSUBS 0.006721f
C61 B.n33 VSUBS 0.006721f
C62 B.n34 VSUBS 0.006721f
C63 B.n35 VSUBS 0.006721f
C64 B.n36 VSUBS 0.006721f
C65 B.n37 VSUBS 0.006721f
C66 B.n38 VSUBS 0.006721f
C67 B.n39 VSUBS 0.006721f
C68 B.n40 VSUBS 0.006721f
C69 B.n41 VSUBS 0.006721f
C70 B.n42 VSUBS 0.006721f
C71 B.n43 VSUBS 0.006721f
C72 B.n44 VSUBS 0.006721f
C73 B.n45 VSUBS 0.006721f
C74 B.n46 VSUBS 0.006721f
C75 B.n47 VSUBS 0.006721f
C76 B.n48 VSUBS 0.006721f
C77 B.n49 VSUBS 0.006721f
C78 B.n50 VSUBS 0.006721f
C79 B.n51 VSUBS 0.006721f
C80 B.t8 VSUBS 0.643727f
C81 B.t7 VSUBS 0.657644f
C82 B.t6 VSUBS 1.21002f
C83 B.n52 VSUBS 0.288431f
C84 B.n53 VSUBS 0.065002f
C85 B.n54 VSUBS 0.006721f
C86 B.n55 VSUBS 0.006721f
C87 B.n56 VSUBS 0.006721f
C88 B.n57 VSUBS 0.006721f
C89 B.n58 VSUBS 0.003756f
C90 B.n59 VSUBS 0.006721f
C91 B.t5 VSUBS 0.643699f
C92 B.t4 VSUBS 0.657621f
C93 B.t3 VSUBS 1.21002f
C94 B.n60 VSUBS 0.288455f
C95 B.n61 VSUBS 0.06503f
C96 B.n62 VSUBS 0.015571f
C97 B.n63 VSUBS 0.006721f
C98 B.n64 VSUBS 0.006721f
C99 B.n65 VSUBS 0.006721f
C100 B.n66 VSUBS 0.006721f
C101 B.n67 VSUBS 0.006721f
C102 B.n68 VSUBS 0.006721f
C103 B.n69 VSUBS 0.006721f
C104 B.n70 VSUBS 0.006721f
C105 B.n71 VSUBS 0.006721f
C106 B.n72 VSUBS 0.006721f
C107 B.n73 VSUBS 0.006721f
C108 B.n74 VSUBS 0.006721f
C109 B.n75 VSUBS 0.006721f
C110 B.n76 VSUBS 0.006721f
C111 B.n77 VSUBS 0.006721f
C112 B.n78 VSUBS 0.006721f
C113 B.n79 VSUBS 0.006721f
C114 B.n80 VSUBS 0.006721f
C115 B.n81 VSUBS 0.006721f
C116 B.n82 VSUBS 0.006721f
C117 B.n83 VSUBS 0.006721f
C118 B.n84 VSUBS 0.006721f
C119 B.n85 VSUBS 0.006721f
C120 B.n86 VSUBS 0.006721f
C121 B.n87 VSUBS 0.006721f
C122 B.n88 VSUBS 0.006721f
C123 B.n89 VSUBS 0.006721f
C124 B.n90 VSUBS 0.006721f
C125 B.n91 VSUBS 0.006721f
C126 B.n92 VSUBS 0.006721f
C127 B.n93 VSUBS 0.016425f
C128 B.n94 VSUBS 0.006721f
C129 B.n95 VSUBS 0.006721f
C130 B.n96 VSUBS 0.006721f
C131 B.n97 VSUBS 0.006721f
C132 B.n98 VSUBS 0.006721f
C133 B.n99 VSUBS 0.006721f
C134 B.n100 VSUBS 0.006721f
C135 B.n101 VSUBS 0.006721f
C136 B.n102 VSUBS 0.006721f
C137 B.n103 VSUBS 0.006721f
C138 B.n104 VSUBS 0.006721f
C139 B.n105 VSUBS 0.006721f
C140 B.n106 VSUBS 0.006721f
C141 B.n107 VSUBS 0.006721f
C142 B.n108 VSUBS 0.006721f
C143 B.n109 VSUBS 0.006721f
C144 B.n110 VSUBS 0.006721f
C145 B.n111 VSUBS 0.006721f
C146 B.n112 VSUBS 0.006721f
C147 B.n113 VSUBS 0.006721f
C148 B.n114 VSUBS 0.006721f
C149 B.n115 VSUBS 0.006721f
C150 B.n116 VSUBS 0.006721f
C151 B.n117 VSUBS 0.006721f
C152 B.n118 VSUBS 0.006721f
C153 B.n119 VSUBS 0.006721f
C154 B.n120 VSUBS 0.006721f
C155 B.n121 VSUBS 0.006721f
C156 B.n122 VSUBS 0.006721f
C157 B.n123 VSUBS 0.006721f
C158 B.n124 VSUBS 0.006721f
C159 B.n125 VSUBS 0.006721f
C160 B.n126 VSUBS 0.006721f
C161 B.n127 VSUBS 0.006721f
C162 B.n128 VSUBS 0.006721f
C163 B.n129 VSUBS 0.017144f
C164 B.n130 VSUBS 0.006721f
C165 B.n131 VSUBS 0.006721f
C166 B.n132 VSUBS 0.006721f
C167 B.n133 VSUBS 0.006721f
C168 B.n134 VSUBS 0.006721f
C169 B.n135 VSUBS 0.006721f
C170 B.n136 VSUBS 0.006721f
C171 B.n137 VSUBS 0.006721f
C172 B.n138 VSUBS 0.006721f
C173 B.n139 VSUBS 0.006721f
C174 B.n140 VSUBS 0.006721f
C175 B.n141 VSUBS 0.006721f
C176 B.n142 VSUBS 0.006721f
C177 B.n143 VSUBS 0.006721f
C178 B.n144 VSUBS 0.006721f
C179 B.n145 VSUBS 0.006721f
C180 B.n146 VSUBS 0.006721f
C181 B.n147 VSUBS 0.006721f
C182 B.n148 VSUBS 0.006721f
C183 B.n149 VSUBS 0.006721f
C184 B.n150 VSUBS 0.006721f
C185 B.n151 VSUBS 0.006721f
C186 B.n152 VSUBS 0.006721f
C187 B.n153 VSUBS 0.006721f
C188 B.n154 VSUBS 0.006721f
C189 B.n155 VSUBS 0.006721f
C190 B.n156 VSUBS 0.006721f
C191 B.n157 VSUBS 0.006721f
C192 B.n158 VSUBS 0.006721f
C193 B.n159 VSUBS 0.006721f
C194 B.n160 VSUBS 0.006721f
C195 B.t10 VSUBS 0.643699f
C196 B.t11 VSUBS 0.657621f
C197 B.t9 VSUBS 1.21002f
C198 B.n161 VSUBS 0.288455f
C199 B.n162 VSUBS 0.06503f
C200 B.n163 VSUBS 0.015571f
C201 B.n164 VSUBS 0.006721f
C202 B.n165 VSUBS 0.006721f
C203 B.n166 VSUBS 0.006721f
C204 B.n167 VSUBS 0.006721f
C205 B.n168 VSUBS 0.006721f
C206 B.t1 VSUBS 0.643727f
C207 B.t2 VSUBS 0.657644f
C208 B.t0 VSUBS 1.21002f
C209 B.n169 VSUBS 0.288431f
C210 B.n170 VSUBS 0.065002f
C211 B.n171 VSUBS 0.006721f
C212 B.n172 VSUBS 0.006721f
C213 B.n173 VSUBS 0.006721f
C214 B.n174 VSUBS 0.006721f
C215 B.n175 VSUBS 0.006721f
C216 B.n176 VSUBS 0.006721f
C217 B.n177 VSUBS 0.006721f
C218 B.n178 VSUBS 0.006721f
C219 B.n179 VSUBS 0.006721f
C220 B.n180 VSUBS 0.006721f
C221 B.n181 VSUBS 0.006721f
C222 B.n182 VSUBS 0.006721f
C223 B.n183 VSUBS 0.006721f
C224 B.n184 VSUBS 0.006721f
C225 B.n185 VSUBS 0.006721f
C226 B.n186 VSUBS 0.006721f
C227 B.n187 VSUBS 0.006721f
C228 B.n188 VSUBS 0.006721f
C229 B.n189 VSUBS 0.006721f
C230 B.n190 VSUBS 0.006721f
C231 B.n191 VSUBS 0.006721f
C232 B.n192 VSUBS 0.006721f
C233 B.n193 VSUBS 0.006721f
C234 B.n194 VSUBS 0.006721f
C235 B.n195 VSUBS 0.006721f
C236 B.n196 VSUBS 0.006721f
C237 B.n197 VSUBS 0.006721f
C238 B.n198 VSUBS 0.006721f
C239 B.n199 VSUBS 0.006721f
C240 B.n200 VSUBS 0.006721f
C241 B.n201 VSUBS 0.006721f
C242 B.n202 VSUBS 0.017144f
C243 B.n203 VSUBS 0.006721f
C244 B.n204 VSUBS 0.006721f
C245 B.n205 VSUBS 0.006721f
C246 B.n206 VSUBS 0.006721f
C247 B.n207 VSUBS 0.006721f
C248 B.n208 VSUBS 0.006721f
C249 B.n209 VSUBS 0.006721f
C250 B.n210 VSUBS 0.006721f
C251 B.n211 VSUBS 0.006721f
C252 B.n212 VSUBS 0.006721f
C253 B.n213 VSUBS 0.006721f
C254 B.n214 VSUBS 0.006721f
C255 B.n215 VSUBS 0.006721f
C256 B.n216 VSUBS 0.006721f
C257 B.n217 VSUBS 0.006721f
C258 B.n218 VSUBS 0.006721f
C259 B.n219 VSUBS 0.006721f
C260 B.n220 VSUBS 0.006721f
C261 B.n221 VSUBS 0.006721f
C262 B.n222 VSUBS 0.006721f
C263 B.n223 VSUBS 0.006721f
C264 B.n224 VSUBS 0.006721f
C265 B.n225 VSUBS 0.006721f
C266 B.n226 VSUBS 0.006721f
C267 B.n227 VSUBS 0.006721f
C268 B.n228 VSUBS 0.006721f
C269 B.n229 VSUBS 0.006721f
C270 B.n230 VSUBS 0.006721f
C271 B.n231 VSUBS 0.006721f
C272 B.n232 VSUBS 0.006721f
C273 B.n233 VSUBS 0.006721f
C274 B.n234 VSUBS 0.006721f
C275 B.n235 VSUBS 0.006721f
C276 B.n236 VSUBS 0.006721f
C277 B.n237 VSUBS 0.006721f
C278 B.n238 VSUBS 0.006721f
C279 B.n239 VSUBS 0.006721f
C280 B.n240 VSUBS 0.006721f
C281 B.n241 VSUBS 0.006721f
C282 B.n242 VSUBS 0.006721f
C283 B.n243 VSUBS 0.006721f
C284 B.n244 VSUBS 0.006721f
C285 B.n245 VSUBS 0.006721f
C286 B.n246 VSUBS 0.006721f
C287 B.n247 VSUBS 0.006721f
C288 B.n248 VSUBS 0.006721f
C289 B.n249 VSUBS 0.006721f
C290 B.n250 VSUBS 0.006721f
C291 B.n251 VSUBS 0.006721f
C292 B.n252 VSUBS 0.006721f
C293 B.n253 VSUBS 0.006721f
C294 B.n254 VSUBS 0.006721f
C295 B.n255 VSUBS 0.006721f
C296 B.n256 VSUBS 0.006721f
C297 B.n257 VSUBS 0.006721f
C298 B.n258 VSUBS 0.006721f
C299 B.n259 VSUBS 0.006721f
C300 B.n260 VSUBS 0.006721f
C301 B.n261 VSUBS 0.006721f
C302 B.n262 VSUBS 0.006721f
C303 B.n263 VSUBS 0.006721f
C304 B.n264 VSUBS 0.006721f
C305 B.n265 VSUBS 0.006721f
C306 B.n266 VSUBS 0.006721f
C307 B.n267 VSUBS 0.006721f
C308 B.n268 VSUBS 0.006721f
C309 B.n269 VSUBS 0.01646f
C310 B.n270 VSUBS 0.01646f
C311 B.n271 VSUBS 0.017144f
C312 B.n272 VSUBS 0.006721f
C313 B.n273 VSUBS 0.006721f
C314 B.n274 VSUBS 0.006721f
C315 B.n275 VSUBS 0.006721f
C316 B.n276 VSUBS 0.006721f
C317 B.n277 VSUBS 0.006721f
C318 B.n278 VSUBS 0.006721f
C319 B.n279 VSUBS 0.006721f
C320 B.n280 VSUBS 0.006721f
C321 B.n281 VSUBS 0.006721f
C322 B.n282 VSUBS 0.006721f
C323 B.n283 VSUBS 0.006721f
C324 B.n284 VSUBS 0.006721f
C325 B.n285 VSUBS 0.006721f
C326 B.n286 VSUBS 0.006721f
C327 B.n287 VSUBS 0.006721f
C328 B.n288 VSUBS 0.006721f
C329 B.n289 VSUBS 0.006721f
C330 B.n290 VSUBS 0.006721f
C331 B.n291 VSUBS 0.006721f
C332 B.n292 VSUBS 0.006721f
C333 B.n293 VSUBS 0.006721f
C334 B.n294 VSUBS 0.006721f
C335 B.n295 VSUBS 0.006721f
C336 B.n296 VSUBS 0.006721f
C337 B.n297 VSUBS 0.006721f
C338 B.n298 VSUBS 0.006721f
C339 B.n299 VSUBS 0.006721f
C340 B.n300 VSUBS 0.006721f
C341 B.n301 VSUBS 0.006721f
C342 B.n302 VSUBS 0.006721f
C343 B.n303 VSUBS 0.006721f
C344 B.n304 VSUBS 0.006721f
C345 B.n305 VSUBS 0.006721f
C346 B.n306 VSUBS 0.006721f
C347 B.n307 VSUBS 0.006721f
C348 B.n308 VSUBS 0.006721f
C349 B.n309 VSUBS 0.006721f
C350 B.n310 VSUBS 0.006721f
C351 B.n311 VSUBS 0.006721f
C352 B.n312 VSUBS 0.006721f
C353 B.n313 VSUBS 0.006721f
C354 B.n314 VSUBS 0.006721f
C355 B.n315 VSUBS 0.006721f
C356 B.n316 VSUBS 0.006721f
C357 B.n317 VSUBS 0.006721f
C358 B.n318 VSUBS 0.006721f
C359 B.n319 VSUBS 0.006721f
C360 B.n320 VSUBS 0.006721f
C361 B.n321 VSUBS 0.006721f
C362 B.n322 VSUBS 0.006721f
C363 B.n323 VSUBS 0.006721f
C364 B.n324 VSUBS 0.006721f
C365 B.n325 VSUBS 0.006721f
C366 B.n326 VSUBS 0.006721f
C367 B.n327 VSUBS 0.006721f
C368 B.n328 VSUBS 0.006721f
C369 B.n329 VSUBS 0.006721f
C370 B.n330 VSUBS 0.006721f
C371 B.n331 VSUBS 0.006721f
C372 B.n332 VSUBS 0.006721f
C373 B.n333 VSUBS 0.006721f
C374 B.n334 VSUBS 0.006721f
C375 B.n335 VSUBS 0.006721f
C376 B.n336 VSUBS 0.006721f
C377 B.n337 VSUBS 0.006721f
C378 B.n338 VSUBS 0.006721f
C379 B.n339 VSUBS 0.006721f
C380 B.n340 VSUBS 0.006721f
C381 B.n341 VSUBS 0.006721f
C382 B.n342 VSUBS 0.006721f
C383 B.n343 VSUBS 0.006721f
C384 B.n344 VSUBS 0.006721f
C385 B.n345 VSUBS 0.006721f
C386 B.n346 VSUBS 0.006721f
C387 B.n347 VSUBS 0.006721f
C388 B.n348 VSUBS 0.006721f
C389 B.n349 VSUBS 0.006721f
C390 B.n350 VSUBS 0.006721f
C391 B.n351 VSUBS 0.006721f
C392 B.n352 VSUBS 0.006721f
C393 B.n353 VSUBS 0.006721f
C394 B.n354 VSUBS 0.006721f
C395 B.n355 VSUBS 0.006721f
C396 B.n356 VSUBS 0.006721f
C397 B.n357 VSUBS 0.006721f
C398 B.n358 VSUBS 0.006721f
C399 B.n359 VSUBS 0.006721f
C400 B.n360 VSUBS 0.006721f
C401 B.n361 VSUBS 0.006721f
C402 B.n362 VSUBS 0.006721f
C403 B.n363 VSUBS 0.006721f
C404 B.n364 VSUBS 0.006721f
C405 B.n365 VSUBS 0.006721f
C406 B.n366 VSUBS 0.006325f
C407 B.n367 VSUBS 0.015571f
C408 B.n368 VSUBS 0.003756f
C409 B.n369 VSUBS 0.006721f
C410 B.n370 VSUBS 0.006721f
C411 B.n371 VSUBS 0.006721f
C412 B.n372 VSUBS 0.006721f
C413 B.n373 VSUBS 0.006721f
C414 B.n374 VSUBS 0.006721f
C415 B.n375 VSUBS 0.006721f
C416 B.n376 VSUBS 0.006721f
C417 B.n377 VSUBS 0.006721f
C418 B.n378 VSUBS 0.006721f
C419 B.n379 VSUBS 0.006721f
C420 B.n380 VSUBS 0.006721f
C421 B.n381 VSUBS 0.003756f
C422 B.n382 VSUBS 0.006721f
C423 B.n383 VSUBS 0.006721f
C424 B.n384 VSUBS 0.006325f
C425 B.n385 VSUBS 0.006721f
C426 B.n386 VSUBS 0.006721f
C427 B.n387 VSUBS 0.006721f
C428 B.n388 VSUBS 0.006721f
C429 B.n389 VSUBS 0.006721f
C430 B.n390 VSUBS 0.006721f
C431 B.n391 VSUBS 0.006721f
C432 B.n392 VSUBS 0.006721f
C433 B.n393 VSUBS 0.006721f
C434 B.n394 VSUBS 0.006721f
C435 B.n395 VSUBS 0.006721f
C436 B.n396 VSUBS 0.006721f
C437 B.n397 VSUBS 0.006721f
C438 B.n398 VSUBS 0.006721f
C439 B.n399 VSUBS 0.006721f
C440 B.n400 VSUBS 0.006721f
C441 B.n401 VSUBS 0.006721f
C442 B.n402 VSUBS 0.006721f
C443 B.n403 VSUBS 0.006721f
C444 B.n404 VSUBS 0.006721f
C445 B.n405 VSUBS 0.006721f
C446 B.n406 VSUBS 0.006721f
C447 B.n407 VSUBS 0.006721f
C448 B.n408 VSUBS 0.006721f
C449 B.n409 VSUBS 0.006721f
C450 B.n410 VSUBS 0.006721f
C451 B.n411 VSUBS 0.006721f
C452 B.n412 VSUBS 0.006721f
C453 B.n413 VSUBS 0.006721f
C454 B.n414 VSUBS 0.006721f
C455 B.n415 VSUBS 0.006721f
C456 B.n416 VSUBS 0.006721f
C457 B.n417 VSUBS 0.006721f
C458 B.n418 VSUBS 0.006721f
C459 B.n419 VSUBS 0.006721f
C460 B.n420 VSUBS 0.006721f
C461 B.n421 VSUBS 0.006721f
C462 B.n422 VSUBS 0.006721f
C463 B.n423 VSUBS 0.006721f
C464 B.n424 VSUBS 0.006721f
C465 B.n425 VSUBS 0.006721f
C466 B.n426 VSUBS 0.006721f
C467 B.n427 VSUBS 0.006721f
C468 B.n428 VSUBS 0.006721f
C469 B.n429 VSUBS 0.006721f
C470 B.n430 VSUBS 0.006721f
C471 B.n431 VSUBS 0.006721f
C472 B.n432 VSUBS 0.006721f
C473 B.n433 VSUBS 0.006721f
C474 B.n434 VSUBS 0.006721f
C475 B.n435 VSUBS 0.006721f
C476 B.n436 VSUBS 0.006721f
C477 B.n437 VSUBS 0.006721f
C478 B.n438 VSUBS 0.006721f
C479 B.n439 VSUBS 0.006721f
C480 B.n440 VSUBS 0.006721f
C481 B.n441 VSUBS 0.006721f
C482 B.n442 VSUBS 0.006721f
C483 B.n443 VSUBS 0.006721f
C484 B.n444 VSUBS 0.006721f
C485 B.n445 VSUBS 0.006721f
C486 B.n446 VSUBS 0.006721f
C487 B.n447 VSUBS 0.006721f
C488 B.n448 VSUBS 0.006721f
C489 B.n449 VSUBS 0.006721f
C490 B.n450 VSUBS 0.006721f
C491 B.n451 VSUBS 0.006721f
C492 B.n452 VSUBS 0.006721f
C493 B.n453 VSUBS 0.006721f
C494 B.n454 VSUBS 0.006721f
C495 B.n455 VSUBS 0.006721f
C496 B.n456 VSUBS 0.006721f
C497 B.n457 VSUBS 0.006721f
C498 B.n458 VSUBS 0.006721f
C499 B.n459 VSUBS 0.006721f
C500 B.n460 VSUBS 0.006721f
C501 B.n461 VSUBS 0.006721f
C502 B.n462 VSUBS 0.006721f
C503 B.n463 VSUBS 0.006721f
C504 B.n464 VSUBS 0.006721f
C505 B.n465 VSUBS 0.006721f
C506 B.n466 VSUBS 0.006721f
C507 B.n467 VSUBS 0.006721f
C508 B.n468 VSUBS 0.006721f
C509 B.n469 VSUBS 0.006721f
C510 B.n470 VSUBS 0.006721f
C511 B.n471 VSUBS 0.006721f
C512 B.n472 VSUBS 0.006721f
C513 B.n473 VSUBS 0.006721f
C514 B.n474 VSUBS 0.006721f
C515 B.n475 VSUBS 0.006721f
C516 B.n476 VSUBS 0.006721f
C517 B.n477 VSUBS 0.006721f
C518 B.n478 VSUBS 0.017144f
C519 B.n479 VSUBS 0.01646f
C520 B.n480 VSUBS 0.01646f
C521 B.n481 VSUBS 0.006721f
C522 B.n482 VSUBS 0.006721f
C523 B.n483 VSUBS 0.006721f
C524 B.n484 VSUBS 0.006721f
C525 B.n485 VSUBS 0.006721f
C526 B.n486 VSUBS 0.006721f
C527 B.n487 VSUBS 0.006721f
C528 B.n488 VSUBS 0.006721f
C529 B.n489 VSUBS 0.006721f
C530 B.n490 VSUBS 0.006721f
C531 B.n491 VSUBS 0.006721f
C532 B.n492 VSUBS 0.006721f
C533 B.n493 VSUBS 0.006721f
C534 B.n494 VSUBS 0.006721f
C535 B.n495 VSUBS 0.006721f
C536 B.n496 VSUBS 0.006721f
C537 B.n497 VSUBS 0.006721f
C538 B.n498 VSUBS 0.006721f
C539 B.n499 VSUBS 0.006721f
C540 B.n500 VSUBS 0.006721f
C541 B.n501 VSUBS 0.006721f
C542 B.n502 VSUBS 0.006721f
C543 B.n503 VSUBS 0.006721f
C544 B.n504 VSUBS 0.006721f
C545 B.n505 VSUBS 0.006721f
C546 B.n506 VSUBS 0.006721f
C547 B.n507 VSUBS 0.006721f
C548 B.n508 VSUBS 0.006721f
C549 B.n509 VSUBS 0.006721f
C550 B.n510 VSUBS 0.006721f
C551 B.n511 VSUBS 0.006721f
C552 B.n512 VSUBS 0.006721f
C553 B.n513 VSUBS 0.006721f
C554 B.n514 VSUBS 0.006721f
C555 B.n515 VSUBS 0.006721f
C556 B.n516 VSUBS 0.006721f
C557 B.n517 VSUBS 0.006721f
C558 B.n518 VSUBS 0.006721f
C559 B.n519 VSUBS 0.006721f
C560 B.n520 VSUBS 0.006721f
C561 B.n521 VSUBS 0.006721f
C562 B.n522 VSUBS 0.006721f
C563 B.n523 VSUBS 0.006721f
C564 B.n524 VSUBS 0.006721f
C565 B.n525 VSUBS 0.006721f
C566 B.n526 VSUBS 0.006721f
C567 B.n527 VSUBS 0.006721f
C568 B.n528 VSUBS 0.006721f
C569 B.n529 VSUBS 0.006721f
C570 B.n530 VSUBS 0.006721f
C571 B.n531 VSUBS 0.006721f
C572 B.n532 VSUBS 0.006721f
C573 B.n533 VSUBS 0.006721f
C574 B.n534 VSUBS 0.006721f
C575 B.n535 VSUBS 0.006721f
C576 B.n536 VSUBS 0.006721f
C577 B.n537 VSUBS 0.006721f
C578 B.n538 VSUBS 0.006721f
C579 B.n539 VSUBS 0.006721f
C580 B.n540 VSUBS 0.006721f
C581 B.n541 VSUBS 0.006721f
C582 B.n542 VSUBS 0.006721f
C583 B.n543 VSUBS 0.006721f
C584 B.n544 VSUBS 0.006721f
C585 B.n545 VSUBS 0.006721f
C586 B.n546 VSUBS 0.006721f
C587 B.n547 VSUBS 0.006721f
C588 B.n548 VSUBS 0.006721f
C589 B.n549 VSUBS 0.006721f
C590 B.n550 VSUBS 0.006721f
C591 B.n551 VSUBS 0.006721f
C592 B.n552 VSUBS 0.006721f
C593 B.n553 VSUBS 0.006721f
C594 B.n554 VSUBS 0.006721f
C595 B.n555 VSUBS 0.006721f
C596 B.n556 VSUBS 0.006721f
C597 B.n557 VSUBS 0.006721f
C598 B.n558 VSUBS 0.006721f
C599 B.n559 VSUBS 0.006721f
C600 B.n560 VSUBS 0.006721f
C601 B.n561 VSUBS 0.006721f
C602 B.n562 VSUBS 0.006721f
C603 B.n563 VSUBS 0.006721f
C604 B.n564 VSUBS 0.006721f
C605 B.n565 VSUBS 0.006721f
C606 B.n566 VSUBS 0.006721f
C607 B.n567 VSUBS 0.006721f
C608 B.n568 VSUBS 0.006721f
C609 B.n569 VSUBS 0.006721f
C610 B.n570 VSUBS 0.006721f
C611 B.n571 VSUBS 0.006721f
C612 B.n572 VSUBS 0.006721f
C613 B.n573 VSUBS 0.006721f
C614 B.n574 VSUBS 0.006721f
C615 B.n575 VSUBS 0.006721f
C616 B.n576 VSUBS 0.006721f
C617 B.n577 VSUBS 0.006721f
C618 B.n578 VSUBS 0.006721f
C619 B.n579 VSUBS 0.006721f
C620 B.n580 VSUBS 0.006721f
C621 B.n581 VSUBS 0.006721f
C622 B.n582 VSUBS 0.006721f
C623 B.n583 VSUBS 0.006721f
C624 B.n584 VSUBS 0.017179f
C625 B.n585 VSUBS 0.01646f
C626 B.n586 VSUBS 0.017144f
C627 B.n587 VSUBS 0.006721f
C628 B.n588 VSUBS 0.006721f
C629 B.n589 VSUBS 0.006721f
C630 B.n590 VSUBS 0.006721f
C631 B.n591 VSUBS 0.006721f
C632 B.n592 VSUBS 0.006721f
C633 B.n593 VSUBS 0.006721f
C634 B.n594 VSUBS 0.006721f
C635 B.n595 VSUBS 0.006721f
C636 B.n596 VSUBS 0.006721f
C637 B.n597 VSUBS 0.006721f
C638 B.n598 VSUBS 0.006721f
C639 B.n599 VSUBS 0.006721f
C640 B.n600 VSUBS 0.006721f
C641 B.n601 VSUBS 0.006721f
C642 B.n602 VSUBS 0.006721f
C643 B.n603 VSUBS 0.006721f
C644 B.n604 VSUBS 0.006721f
C645 B.n605 VSUBS 0.006721f
C646 B.n606 VSUBS 0.006721f
C647 B.n607 VSUBS 0.006721f
C648 B.n608 VSUBS 0.006721f
C649 B.n609 VSUBS 0.006721f
C650 B.n610 VSUBS 0.006721f
C651 B.n611 VSUBS 0.006721f
C652 B.n612 VSUBS 0.006721f
C653 B.n613 VSUBS 0.006721f
C654 B.n614 VSUBS 0.006721f
C655 B.n615 VSUBS 0.006721f
C656 B.n616 VSUBS 0.006721f
C657 B.n617 VSUBS 0.006721f
C658 B.n618 VSUBS 0.006721f
C659 B.n619 VSUBS 0.006721f
C660 B.n620 VSUBS 0.006721f
C661 B.n621 VSUBS 0.006721f
C662 B.n622 VSUBS 0.006721f
C663 B.n623 VSUBS 0.006721f
C664 B.n624 VSUBS 0.006721f
C665 B.n625 VSUBS 0.006721f
C666 B.n626 VSUBS 0.006721f
C667 B.n627 VSUBS 0.006721f
C668 B.n628 VSUBS 0.006721f
C669 B.n629 VSUBS 0.006721f
C670 B.n630 VSUBS 0.006721f
C671 B.n631 VSUBS 0.006721f
C672 B.n632 VSUBS 0.006721f
C673 B.n633 VSUBS 0.006721f
C674 B.n634 VSUBS 0.006721f
C675 B.n635 VSUBS 0.006721f
C676 B.n636 VSUBS 0.006721f
C677 B.n637 VSUBS 0.006721f
C678 B.n638 VSUBS 0.006721f
C679 B.n639 VSUBS 0.006721f
C680 B.n640 VSUBS 0.006721f
C681 B.n641 VSUBS 0.006721f
C682 B.n642 VSUBS 0.006721f
C683 B.n643 VSUBS 0.006721f
C684 B.n644 VSUBS 0.006721f
C685 B.n645 VSUBS 0.006721f
C686 B.n646 VSUBS 0.006721f
C687 B.n647 VSUBS 0.006721f
C688 B.n648 VSUBS 0.006721f
C689 B.n649 VSUBS 0.006721f
C690 B.n650 VSUBS 0.006721f
C691 B.n651 VSUBS 0.006721f
C692 B.n652 VSUBS 0.006721f
C693 B.n653 VSUBS 0.006721f
C694 B.n654 VSUBS 0.006721f
C695 B.n655 VSUBS 0.006721f
C696 B.n656 VSUBS 0.006721f
C697 B.n657 VSUBS 0.006721f
C698 B.n658 VSUBS 0.006721f
C699 B.n659 VSUBS 0.006721f
C700 B.n660 VSUBS 0.006721f
C701 B.n661 VSUBS 0.006721f
C702 B.n662 VSUBS 0.006721f
C703 B.n663 VSUBS 0.006721f
C704 B.n664 VSUBS 0.006721f
C705 B.n665 VSUBS 0.006721f
C706 B.n666 VSUBS 0.006721f
C707 B.n667 VSUBS 0.006721f
C708 B.n668 VSUBS 0.006721f
C709 B.n669 VSUBS 0.006721f
C710 B.n670 VSUBS 0.006721f
C711 B.n671 VSUBS 0.006721f
C712 B.n672 VSUBS 0.006721f
C713 B.n673 VSUBS 0.006721f
C714 B.n674 VSUBS 0.006721f
C715 B.n675 VSUBS 0.006721f
C716 B.n676 VSUBS 0.006721f
C717 B.n677 VSUBS 0.006721f
C718 B.n678 VSUBS 0.006721f
C719 B.n679 VSUBS 0.006721f
C720 B.n680 VSUBS 0.006325f
C721 B.n681 VSUBS 0.006721f
C722 B.n682 VSUBS 0.006721f
C723 B.n683 VSUBS 0.006721f
C724 B.n684 VSUBS 0.006721f
C725 B.n685 VSUBS 0.006721f
C726 B.n686 VSUBS 0.006721f
C727 B.n687 VSUBS 0.006721f
C728 B.n688 VSUBS 0.006721f
C729 B.n689 VSUBS 0.006721f
C730 B.n690 VSUBS 0.006721f
C731 B.n691 VSUBS 0.006721f
C732 B.n692 VSUBS 0.006721f
C733 B.n693 VSUBS 0.006721f
C734 B.n694 VSUBS 0.006721f
C735 B.n695 VSUBS 0.006721f
C736 B.n696 VSUBS 0.003756f
C737 B.n697 VSUBS 0.015571f
C738 B.n698 VSUBS 0.006325f
C739 B.n699 VSUBS 0.006721f
C740 B.n700 VSUBS 0.006721f
C741 B.n701 VSUBS 0.006721f
C742 B.n702 VSUBS 0.006721f
C743 B.n703 VSUBS 0.006721f
C744 B.n704 VSUBS 0.006721f
C745 B.n705 VSUBS 0.006721f
C746 B.n706 VSUBS 0.006721f
C747 B.n707 VSUBS 0.006721f
C748 B.n708 VSUBS 0.006721f
C749 B.n709 VSUBS 0.006721f
C750 B.n710 VSUBS 0.006721f
C751 B.n711 VSUBS 0.006721f
C752 B.n712 VSUBS 0.006721f
C753 B.n713 VSUBS 0.006721f
C754 B.n714 VSUBS 0.006721f
C755 B.n715 VSUBS 0.006721f
C756 B.n716 VSUBS 0.006721f
C757 B.n717 VSUBS 0.006721f
C758 B.n718 VSUBS 0.006721f
C759 B.n719 VSUBS 0.006721f
C760 B.n720 VSUBS 0.006721f
C761 B.n721 VSUBS 0.006721f
C762 B.n722 VSUBS 0.006721f
C763 B.n723 VSUBS 0.006721f
C764 B.n724 VSUBS 0.006721f
C765 B.n725 VSUBS 0.006721f
C766 B.n726 VSUBS 0.006721f
C767 B.n727 VSUBS 0.006721f
C768 B.n728 VSUBS 0.006721f
C769 B.n729 VSUBS 0.006721f
C770 B.n730 VSUBS 0.006721f
C771 B.n731 VSUBS 0.006721f
C772 B.n732 VSUBS 0.006721f
C773 B.n733 VSUBS 0.006721f
C774 B.n734 VSUBS 0.006721f
C775 B.n735 VSUBS 0.006721f
C776 B.n736 VSUBS 0.006721f
C777 B.n737 VSUBS 0.006721f
C778 B.n738 VSUBS 0.006721f
C779 B.n739 VSUBS 0.006721f
C780 B.n740 VSUBS 0.006721f
C781 B.n741 VSUBS 0.006721f
C782 B.n742 VSUBS 0.006721f
C783 B.n743 VSUBS 0.006721f
C784 B.n744 VSUBS 0.006721f
C785 B.n745 VSUBS 0.006721f
C786 B.n746 VSUBS 0.006721f
C787 B.n747 VSUBS 0.006721f
C788 B.n748 VSUBS 0.006721f
C789 B.n749 VSUBS 0.006721f
C790 B.n750 VSUBS 0.006721f
C791 B.n751 VSUBS 0.006721f
C792 B.n752 VSUBS 0.006721f
C793 B.n753 VSUBS 0.006721f
C794 B.n754 VSUBS 0.006721f
C795 B.n755 VSUBS 0.006721f
C796 B.n756 VSUBS 0.006721f
C797 B.n757 VSUBS 0.006721f
C798 B.n758 VSUBS 0.006721f
C799 B.n759 VSUBS 0.006721f
C800 B.n760 VSUBS 0.006721f
C801 B.n761 VSUBS 0.006721f
C802 B.n762 VSUBS 0.006721f
C803 B.n763 VSUBS 0.006721f
C804 B.n764 VSUBS 0.006721f
C805 B.n765 VSUBS 0.006721f
C806 B.n766 VSUBS 0.006721f
C807 B.n767 VSUBS 0.006721f
C808 B.n768 VSUBS 0.006721f
C809 B.n769 VSUBS 0.006721f
C810 B.n770 VSUBS 0.006721f
C811 B.n771 VSUBS 0.006721f
C812 B.n772 VSUBS 0.006721f
C813 B.n773 VSUBS 0.006721f
C814 B.n774 VSUBS 0.006721f
C815 B.n775 VSUBS 0.006721f
C816 B.n776 VSUBS 0.006721f
C817 B.n777 VSUBS 0.006721f
C818 B.n778 VSUBS 0.006721f
C819 B.n779 VSUBS 0.006721f
C820 B.n780 VSUBS 0.006721f
C821 B.n781 VSUBS 0.006721f
C822 B.n782 VSUBS 0.006721f
C823 B.n783 VSUBS 0.006721f
C824 B.n784 VSUBS 0.006721f
C825 B.n785 VSUBS 0.006721f
C826 B.n786 VSUBS 0.006721f
C827 B.n787 VSUBS 0.006721f
C828 B.n788 VSUBS 0.006721f
C829 B.n789 VSUBS 0.006721f
C830 B.n790 VSUBS 0.006721f
C831 B.n791 VSUBS 0.006721f
C832 B.n792 VSUBS 0.017144f
C833 B.n793 VSUBS 0.017144f
C834 B.n794 VSUBS 0.01646f
C835 B.n795 VSUBS 0.006721f
C836 B.n796 VSUBS 0.006721f
C837 B.n797 VSUBS 0.006721f
C838 B.n798 VSUBS 0.006721f
C839 B.n799 VSUBS 0.006721f
C840 B.n800 VSUBS 0.006721f
C841 B.n801 VSUBS 0.006721f
C842 B.n802 VSUBS 0.006721f
C843 B.n803 VSUBS 0.006721f
C844 B.n804 VSUBS 0.006721f
C845 B.n805 VSUBS 0.006721f
C846 B.n806 VSUBS 0.006721f
C847 B.n807 VSUBS 0.006721f
C848 B.n808 VSUBS 0.006721f
C849 B.n809 VSUBS 0.006721f
C850 B.n810 VSUBS 0.006721f
C851 B.n811 VSUBS 0.006721f
C852 B.n812 VSUBS 0.006721f
C853 B.n813 VSUBS 0.006721f
C854 B.n814 VSUBS 0.006721f
C855 B.n815 VSUBS 0.006721f
C856 B.n816 VSUBS 0.006721f
C857 B.n817 VSUBS 0.006721f
C858 B.n818 VSUBS 0.006721f
C859 B.n819 VSUBS 0.006721f
C860 B.n820 VSUBS 0.006721f
C861 B.n821 VSUBS 0.006721f
C862 B.n822 VSUBS 0.006721f
C863 B.n823 VSUBS 0.006721f
C864 B.n824 VSUBS 0.006721f
C865 B.n825 VSUBS 0.006721f
C866 B.n826 VSUBS 0.006721f
C867 B.n827 VSUBS 0.006721f
C868 B.n828 VSUBS 0.006721f
C869 B.n829 VSUBS 0.006721f
C870 B.n830 VSUBS 0.006721f
C871 B.n831 VSUBS 0.006721f
C872 B.n832 VSUBS 0.006721f
C873 B.n833 VSUBS 0.006721f
C874 B.n834 VSUBS 0.006721f
C875 B.n835 VSUBS 0.006721f
C876 B.n836 VSUBS 0.006721f
C877 B.n837 VSUBS 0.006721f
C878 B.n838 VSUBS 0.006721f
C879 B.n839 VSUBS 0.006721f
C880 B.n840 VSUBS 0.006721f
C881 B.n841 VSUBS 0.006721f
C882 B.n842 VSUBS 0.006721f
C883 B.n843 VSUBS 0.006721f
C884 B.n844 VSUBS 0.006721f
C885 B.n845 VSUBS 0.006721f
C886 B.n846 VSUBS 0.006721f
C887 B.n847 VSUBS 0.015218f
C888 VDD1.t2 VSUBS 0.392905f
C889 VDD1.t0 VSUBS 0.392905f
C890 VDD1.n0 VSUBS 3.32084f
C891 VDD1.t6 VSUBS 0.392905f
C892 VDD1.t5 VSUBS 0.392905f
C893 VDD1.n1 VSUBS 3.31963f
C894 VDD1.t4 VSUBS 0.392905f
C895 VDD1.t3 VSUBS 0.392905f
C896 VDD1.n2 VSUBS 3.31963f
C897 VDD1.n3 VSUBS 3.76839f
C898 VDD1.t1 VSUBS 0.392905f
C899 VDD1.t7 VSUBS 0.392905f
C900 VDD1.n4 VSUBS 3.31231f
C901 VDD1.n5 VSUBS 3.49747f
C902 VP.n0 VSUBS 0.03582f
C903 VP.t4 VSUBS 2.94167f
C904 VP.n1 VSUBS 0.060901f
C905 VP.n2 VSUBS 0.03582f
C906 VP.t3 VSUBS 2.94167f
C907 VP.n3 VSUBS 0.06557f
C908 VP.n4 VSUBS 0.03582f
C909 VP.n5 VSUBS 0.051305f
C910 VP.n6 VSUBS 0.03582f
C911 VP.t0 VSUBS 2.94167f
C912 VP.n7 VSUBS 0.060901f
C913 VP.n8 VSUBS 0.03582f
C914 VP.t6 VSUBS 2.94167f
C915 VP.n9 VSUBS 0.06557f
C916 VP.t5 VSUBS 3.05957f
C917 VP.t7 VSUBS 2.94167f
C918 VP.n10 VSUBS 1.10847f
C919 VP.n11 VSUBS 1.11008f
C920 VP.n12 VSUBS 0.228387f
C921 VP.n13 VSUBS 0.03582f
C922 VP.n14 VSUBS 0.028931f
C923 VP.n15 VSUBS 0.06557f
C924 VP.n16 VSUBS 1.03019f
C925 VP.n17 VSUBS 0.038879f
C926 VP.n18 VSUBS 0.03582f
C927 VP.n19 VSUBS 0.03582f
C928 VP.n20 VSUBS 0.03582f
C929 VP.n21 VSUBS 0.042618f
C930 VP.n22 VSUBS 0.051305f
C931 VP.n23 VSUBS 1.10859f
C932 VP.n24 VSUBS 2.04851f
C933 VP.t1 VSUBS 2.94167f
C934 VP.n25 VSUBS 1.10859f
C935 VP.n26 VSUBS 2.07353f
C936 VP.n27 VSUBS 0.03582f
C937 VP.n28 VSUBS 0.03582f
C938 VP.n29 VSUBS 0.042618f
C939 VP.n30 VSUBS 0.060901f
C940 VP.t2 VSUBS 2.94167f
C941 VP.n31 VSUBS 1.03019f
C942 VP.n32 VSUBS 0.038879f
C943 VP.n33 VSUBS 0.03582f
C944 VP.n34 VSUBS 0.03582f
C945 VP.n35 VSUBS 0.03582f
C946 VP.n36 VSUBS 0.028931f
C947 VP.n37 VSUBS 0.06557f
C948 VP.n38 VSUBS 1.03019f
C949 VP.n39 VSUBS 0.038879f
C950 VP.n40 VSUBS 0.03582f
C951 VP.n41 VSUBS 0.03582f
C952 VP.n42 VSUBS 0.03582f
C953 VP.n43 VSUBS 0.042618f
C954 VP.n44 VSUBS 0.051305f
C955 VP.n45 VSUBS 1.10859f
C956 VP.n46 VSUBS 0.033496f
C957 VDD2.t6 VSUBS 0.391183f
C958 VDD2.t7 VSUBS 0.391183f
C959 VDD2.n0 VSUBS 3.30508f
C960 VDD2.t1 VSUBS 0.391183f
C961 VDD2.t2 VSUBS 0.391183f
C962 VDD2.n1 VSUBS 3.30508f
C963 VDD2.n2 VSUBS 3.69936f
C964 VDD2.t0 VSUBS 0.391183f
C965 VDD2.t3 VSUBS 0.391183f
C966 VDD2.n3 VSUBS 3.2978f
C967 VDD2.n4 VSUBS 3.45142f
C968 VDD2.t4 VSUBS 0.391183f
C969 VDD2.t5 VSUBS 0.391183f
C970 VDD2.n5 VSUBS 3.30503f
C971 VTAIL.t15 VSUBS 0.35833f
C972 VTAIL.t13 VSUBS 0.35833f
C973 VTAIL.n0 VSUBS 2.87937f
C974 VTAIL.n1 VSUBS 0.679135f
C975 VTAIL.t14 VSUBS 3.74967f
C976 VTAIL.n2 VSUBS 0.81657f
C977 VTAIL.t0 VSUBS 3.74967f
C978 VTAIL.n3 VSUBS 0.81657f
C979 VTAIL.t7 VSUBS 0.35833f
C980 VTAIL.t5 VSUBS 0.35833f
C981 VTAIL.n4 VSUBS 2.87937f
C982 VTAIL.n5 VSUBS 0.792235f
C983 VTAIL.t6 VSUBS 3.74967f
C984 VTAIL.n6 VSUBS 2.47082f
C985 VTAIL.t11 VSUBS 3.74967f
C986 VTAIL.n7 VSUBS 2.47082f
C987 VTAIL.t12 VSUBS 0.35833f
C988 VTAIL.t9 VSUBS 0.35833f
C989 VTAIL.n8 VSUBS 2.87937f
C990 VTAIL.n9 VSUBS 0.792235f
C991 VTAIL.t8 VSUBS 3.74967f
C992 VTAIL.n10 VSUBS 0.816569f
C993 VTAIL.t1 VSUBS 3.74967f
C994 VTAIL.n11 VSUBS 0.816569f
C995 VTAIL.t3 VSUBS 0.35833f
C996 VTAIL.t4 VSUBS 0.35833f
C997 VTAIL.n12 VSUBS 2.87937f
C998 VTAIL.n13 VSUBS 0.792235f
C999 VTAIL.t2 VSUBS 3.74967f
C1000 VTAIL.n14 VSUBS 2.47082f
C1001 VTAIL.t10 VSUBS 3.74967f
C1002 VTAIL.n15 VSUBS 2.46652f
C1003 VN.n0 VSUBS 0.035024f
C1004 VN.t5 VSUBS 2.87627f
C1005 VN.n1 VSUBS 0.059547f
C1006 VN.n2 VSUBS 0.035024f
C1007 VN.t6 VSUBS 2.87627f
C1008 VN.n3 VSUBS 0.064113f
C1009 VN.t1 VSUBS 2.99155f
C1010 VN.t0 VSUBS 2.87627f
C1011 VN.n4 VSUBS 1.08382f
C1012 VN.n5 VSUBS 1.08541f
C1013 VN.n6 VSUBS 0.22331f
C1014 VN.n7 VSUBS 0.035024f
C1015 VN.n8 VSUBS 0.028287f
C1016 VN.n9 VSUBS 0.064113f
C1017 VN.n10 VSUBS 1.00729f
C1018 VN.n11 VSUBS 0.038015f
C1019 VN.n12 VSUBS 0.035024f
C1020 VN.n13 VSUBS 0.035024f
C1021 VN.n14 VSUBS 0.035024f
C1022 VN.n15 VSUBS 0.04167f
C1023 VN.n16 VSUBS 0.050165f
C1024 VN.n17 VSUBS 1.08394f
C1025 VN.n18 VSUBS 0.032751f
C1026 VN.n19 VSUBS 0.035024f
C1027 VN.t7 VSUBS 2.87627f
C1028 VN.n20 VSUBS 0.059547f
C1029 VN.n21 VSUBS 0.035024f
C1030 VN.t4 VSUBS 2.87627f
C1031 VN.n22 VSUBS 0.064113f
C1032 VN.t2 VSUBS 2.99155f
C1033 VN.t3 VSUBS 2.87627f
C1034 VN.n23 VSUBS 1.08382f
C1035 VN.n24 VSUBS 1.08541f
C1036 VN.n25 VSUBS 0.22331f
C1037 VN.n26 VSUBS 0.035024f
C1038 VN.n27 VSUBS 0.028287f
C1039 VN.n28 VSUBS 0.064113f
C1040 VN.n29 VSUBS 1.00729f
C1041 VN.n30 VSUBS 0.038015f
C1042 VN.n31 VSUBS 0.035024f
C1043 VN.n32 VSUBS 0.035024f
C1044 VN.n33 VSUBS 0.035024f
C1045 VN.n34 VSUBS 0.04167f
C1046 VN.n35 VSUBS 0.050165f
C1047 VN.n36 VSUBS 1.08394f
C1048 VN.n37 VSUBS 2.02571f
.ends

