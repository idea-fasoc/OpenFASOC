* NGSPICE file created from diff_pair_sample_0950.ext - technology: sky130A

.subckt diff_pair_sample_0950 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1762_n3218# sky130_fd_pr__pfet_01v8 ad=4.3875 pd=23.28 as=0 ps=0 w=11.25 l=1.65
X1 B.t8 B.t6 B.t7 w_n1762_n3218# sky130_fd_pr__pfet_01v8 ad=4.3875 pd=23.28 as=0 ps=0 w=11.25 l=1.65
X2 VDD2.t1 VN.t0 VTAIL.t3 w_n1762_n3218# sky130_fd_pr__pfet_01v8 ad=4.3875 pd=23.28 as=4.3875 ps=23.28 w=11.25 l=1.65
X3 VDD1.t1 VP.t0 VTAIL.t0 w_n1762_n3218# sky130_fd_pr__pfet_01v8 ad=4.3875 pd=23.28 as=4.3875 ps=23.28 w=11.25 l=1.65
X4 B.t5 B.t3 B.t4 w_n1762_n3218# sky130_fd_pr__pfet_01v8 ad=4.3875 pd=23.28 as=0 ps=0 w=11.25 l=1.65
X5 VDD1.t0 VP.t1 VTAIL.t1 w_n1762_n3218# sky130_fd_pr__pfet_01v8 ad=4.3875 pd=23.28 as=4.3875 ps=23.28 w=11.25 l=1.65
X6 B.t2 B.t0 B.t1 w_n1762_n3218# sky130_fd_pr__pfet_01v8 ad=4.3875 pd=23.28 as=0 ps=0 w=11.25 l=1.65
X7 VDD2.t0 VN.t1 VTAIL.t2 w_n1762_n3218# sky130_fd_pr__pfet_01v8 ad=4.3875 pd=23.28 as=4.3875 ps=23.28 w=11.25 l=1.65
R0 B.n297 B.n80 585
R1 B.n296 B.n295 585
R2 B.n294 B.n81 585
R3 B.n293 B.n292 585
R4 B.n291 B.n82 585
R5 B.n290 B.n289 585
R6 B.n288 B.n83 585
R7 B.n287 B.n286 585
R8 B.n285 B.n84 585
R9 B.n284 B.n283 585
R10 B.n282 B.n85 585
R11 B.n281 B.n280 585
R12 B.n279 B.n86 585
R13 B.n278 B.n277 585
R14 B.n276 B.n87 585
R15 B.n275 B.n274 585
R16 B.n273 B.n88 585
R17 B.n272 B.n271 585
R18 B.n270 B.n89 585
R19 B.n269 B.n268 585
R20 B.n267 B.n90 585
R21 B.n266 B.n265 585
R22 B.n264 B.n91 585
R23 B.n263 B.n262 585
R24 B.n261 B.n92 585
R25 B.n260 B.n259 585
R26 B.n258 B.n93 585
R27 B.n257 B.n256 585
R28 B.n255 B.n94 585
R29 B.n254 B.n253 585
R30 B.n252 B.n95 585
R31 B.n251 B.n250 585
R32 B.n249 B.n96 585
R33 B.n248 B.n247 585
R34 B.n246 B.n97 585
R35 B.n245 B.n244 585
R36 B.n243 B.n98 585
R37 B.n242 B.n241 585
R38 B.n240 B.n99 585
R39 B.n238 B.n237 585
R40 B.n236 B.n102 585
R41 B.n235 B.n234 585
R42 B.n233 B.n103 585
R43 B.n232 B.n231 585
R44 B.n230 B.n104 585
R45 B.n229 B.n228 585
R46 B.n227 B.n105 585
R47 B.n226 B.n225 585
R48 B.n224 B.n106 585
R49 B.n223 B.n222 585
R50 B.n218 B.n107 585
R51 B.n217 B.n216 585
R52 B.n215 B.n108 585
R53 B.n214 B.n213 585
R54 B.n212 B.n109 585
R55 B.n211 B.n210 585
R56 B.n209 B.n110 585
R57 B.n208 B.n207 585
R58 B.n206 B.n111 585
R59 B.n205 B.n204 585
R60 B.n203 B.n112 585
R61 B.n202 B.n201 585
R62 B.n200 B.n113 585
R63 B.n199 B.n198 585
R64 B.n197 B.n114 585
R65 B.n196 B.n195 585
R66 B.n194 B.n115 585
R67 B.n193 B.n192 585
R68 B.n191 B.n116 585
R69 B.n190 B.n189 585
R70 B.n188 B.n117 585
R71 B.n187 B.n186 585
R72 B.n185 B.n118 585
R73 B.n184 B.n183 585
R74 B.n182 B.n119 585
R75 B.n181 B.n180 585
R76 B.n179 B.n120 585
R77 B.n178 B.n177 585
R78 B.n176 B.n121 585
R79 B.n175 B.n174 585
R80 B.n173 B.n122 585
R81 B.n172 B.n171 585
R82 B.n170 B.n123 585
R83 B.n169 B.n168 585
R84 B.n167 B.n124 585
R85 B.n166 B.n165 585
R86 B.n164 B.n125 585
R87 B.n163 B.n162 585
R88 B.n299 B.n298 585
R89 B.n300 B.n79 585
R90 B.n302 B.n301 585
R91 B.n303 B.n78 585
R92 B.n305 B.n304 585
R93 B.n306 B.n77 585
R94 B.n308 B.n307 585
R95 B.n309 B.n76 585
R96 B.n311 B.n310 585
R97 B.n312 B.n75 585
R98 B.n314 B.n313 585
R99 B.n315 B.n74 585
R100 B.n317 B.n316 585
R101 B.n318 B.n73 585
R102 B.n320 B.n319 585
R103 B.n321 B.n72 585
R104 B.n323 B.n322 585
R105 B.n324 B.n71 585
R106 B.n326 B.n325 585
R107 B.n327 B.n70 585
R108 B.n329 B.n328 585
R109 B.n330 B.n69 585
R110 B.n332 B.n331 585
R111 B.n333 B.n68 585
R112 B.n335 B.n334 585
R113 B.n336 B.n67 585
R114 B.n338 B.n337 585
R115 B.n339 B.n66 585
R116 B.n341 B.n340 585
R117 B.n342 B.n65 585
R118 B.n344 B.n343 585
R119 B.n345 B.n64 585
R120 B.n347 B.n346 585
R121 B.n348 B.n63 585
R122 B.n350 B.n349 585
R123 B.n351 B.n62 585
R124 B.n353 B.n352 585
R125 B.n354 B.n61 585
R126 B.n356 B.n355 585
R127 B.n357 B.n60 585
R128 B.n491 B.n490 585
R129 B.n489 B.n12 585
R130 B.n488 B.n487 585
R131 B.n486 B.n13 585
R132 B.n485 B.n484 585
R133 B.n483 B.n14 585
R134 B.n482 B.n481 585
R135 B.n480 B.n15 585
R136 B.n479 B.n478 585
R137 B.n477 B.n16 585
R138 B.n476 B.n475 585
R139 B.n474 B.n17 585
R140 B.n473 B.n472 585
R141 B.n471 B.n18 585
R142 B.n470 B.n469 585
R143 B.n468 B.n19 585
R144 B.n467 B.n466 585
R145 B.n465 B.n20 585
R146 B.n464 B.n463 585
R147 B.n462 B.n21 585
R148 B.n461 B.n460 585
R149 B.n459 B.n22 585
R150 B.n458 B.n457 585
R151 B.n456 B.n23 585
R152 B.n455 B.n454 585
R153 B.n453 B.n24 585
R154 B.n452 B.n451 585
R155 B.n450 B.n25 585
R156 B.n449 B.n448 585
R157 B.n447 B.n26 585
R158 B.n446 B.n445 585
R159 B.n444 B.n27 585
R160 B.n443 B.n442 585
R161 B.n441 B.n28 585
R162 B.n440 B.n439 585
R163 B.n438 B.n29 585
R164 B.n437 B.n436 585
R165 B.n435 B.n30 585
R166 B.n434 B.n433 585
R167 B.n431 B.n31 585
R168 B.n430 B.n429 585
R169 B.n428 B.n34 585
R170 B.n427 B.n426 585
R171 B.n425 B.n35 585
R172 B.n424 B.n423 585
R173 B.n422 B.n36 585
R174 B.n421 B.n420 585
R175 B.n419 B.n37 585
R176 B.n418 B.n417 585
R177 B.n416 B.n415 585
R178 B.n414 B.n41 585
R179 B.n413 B.n412 585
R180 B.n411 B.n42 585
R181 B.n410 B.n409 585
R182 B.n408 B.n43 585
R183 B.n407 B.n406 585
R184 B.n405 B.n44 585
R185 B.n404 B.n403 585
R186 B.n402 B.n45 585
R187 B.n401 B.n400 585
R188 B.n399 B.n46 585
R189 B.n398 B.n397 585
R190 B.n396 B.n47 585
R191 B.n395 B.n394 585
R192 B.n393 B.n48 585
R193 B.n392 B.n391 585
R194 B.n390 B.n49 585
R195 B.n389 B.n388 585
R196 B.n387 B.n50 585
R197 B.n386 B.n385 585
R198 B.n384 B.n51 585
R199 B.n383 B.n382 585
R200 B.n381 B.n52 585
R201 B.n380 B.n379 585
R202 B.n378 B.n53 585
R203 B.n377 B.n376 585
R204 B.n375 B.n54 585
R205 B.n374 B.n373 585
R206 B.n372 B.n55 585
R207 B.n371 B.n370 585
R208 B.n369 B.n56 585
R209 B.n368 B.n367 585
R210 B.n366 B.n57 585
R211 B.n365 B.n364 585
R212 B.n363 B.n58 585
R213 B.n362 B.n361 585
R214 B.n360 B.n59 585
R215 B.n359 B.n358 585
R216 B.n492 B.n11 585
R217 B.n494 B.n493 585
R218 B.n495 B.n10 585
R219 B.n497 B.n496 585
R220 B.n498 B.n9 585
R221 B.n500 B.n499 585
R222 B.n501 B.n8 585
R223 B.n503 B.n502 585
R224 B.n504 B.n7 585
R225 B.n506 B.n505 585
R226 B.n507 B.n6 585
R227 B.n509 B.n508 585
R228 B.n510 B.n5 585
R229 B.n512 B.n511 585
R230 B.n513 B.n4 585
R231 B.n515 B.n514 585
R232 B.n516 B.n3 585
R233 B.n518 B.n517 585
R234 B.n519 B.n0 585
R235 B.n2 B.n1 585
R236 B.n136 B.n135 585
R237 B.n137 B.n134 585
R238 B.n139 B.n138 585
R239 B.n140 B.n133 585
R240 B.n142 B.n141 585
R241 B.n143 B.n132 585
R242 B.n145 B.n144 585
R243 B.n146 B.n131 585
R244 B.n148 B.n147 585
R245 B.n149 B.n130 585
R246 B.n151 B.n150 585
R247 B.n152 B.n129 585
R248 B.n154 B.n153 585
R249 B.n155 B.n128 585
R250 B.n157 B.n156 585
R251 B.n158 B.n127 585
R252 B.n160 B.n159 585
R253 B.n161 B.n126 585
R254 B.n162 B.n161 574.183
R255 B.n298 B.n297 574.183
R256 B.n358 B.n357 574.183
R257 B.n490 B.n11 574.183
R258 B.n100 B.t1 400.327
R259 B.n38 B.t5 400.327
R260 B.n219 B.t7 400.327
R261 B.n32 B.t11 400.327
R262 B.n219 B.t6 370.276
R263 B.n100 B.t0 370.276
R264 B.n38 B.t3 370.276
R265 B.n32 B.t9 370.276
R266 B.n101 B.t2 361.926
R267 B.n39 B.t4 361.926
R268 B.n220 B.t8 361.926
R269 B.n33 B.t10 361.926
R270 B.n521 B.n520 256.663
R271 B.n520 B.n519 235.042
R272 B.n520 B.n2 235.042
R273 B.n162 B.n125 163.367
R274 B.n166 B.n125 163.367
R275 B.n167 B.n166 163.367
R276 B.n168 B.n167 163.367
R277 B.n168 B.n123 163.367
R278 B.n172 B.n123 163.367
R279 B.n173 B.n172 163.367
R280 B.n174 B.n173 163.367
R281 B.n174 B.n121 163.367
R282 B.n178 B.n121 163.367
R283 B.n179 B.n178 163.367
R284 B.n180 B.n179 163.367
R285 B.n180 B.n119 163.367
R286 B.n184 B.n119 163.367
R287 B.n185 B.n184 163.367
R288 B.n186 B.n185 163.367
R289 B.n186 B.n117 163.367
R290 B.n190 B.n117 163.367
R291 B.n191 B.n190 163.367
R292 B.n192 B.n191 163.367
R293 B.n192 B.n115 163.367
R294 B.n196 B.n115 163.367
R295 B.n197 B.n196 163.367
R296 B.n198 B.n197 163.367
R297 B.n198 B.n113 163.367
R298 B.n202 B.n113 163.367
R299 B.n203 B.n202 163.367
R300 B.n204 B.n203 163.367
R301 B.n204 B.n111 163.367
R302 B.n208 B.n111 163.367
R303 B.n209 B.n208 163.367
R304 B.n210 B.n209 163.367
R305 B.n210 B.n109 163.367
R306 B.n214 B.n109 163.367
R307 B.n215 B.n214 163.367
R308 B.n216 B.n215 163.367
R309 B.n216 B.n107 163.367
R310 B.n223 B.n107 163.367
R311 B.n224 B.n223 163.367
R312 B.n225 B.n224 163.367
R313 B.n225 B.n105 163.367
R314 B.n229 B.n105 163.367
R315 B.n230 B.n229 163.367
R316 B.n231 B.n230 163.367
R317 B.n231 B.n103 163.367
R318 B.n235 B.n103 163.367
R319 B.n236 B.n235 163.367
R320 B.n237 B.n236 163.367
R321 B.n237 B.n99 163.367
R322 B.n242 B.n99 163.367
R323 B.n243 B.n242 163.367
R324 B.n244 B.n243 163.367
R325 B.n244 B.n97 163.367
R326 B.n248 B.n97 163.367
R327 B.n249 B.n248 163.367
R328 B.n250 B.n249 163.367
R329 B.n250 B.n95 163.367
R330 B.n254 B.n95 163.367
R331 B.n255 B.n254 163.367
R332 B.n256 B.n255 163.367
R333 B.n256 B.n93 163.367
R334 B.n260 B.n93 163.367
R335 B.n261 B.n260 163.367
R336 B.n262 B.n261 163.367
R337 B.n262 B.n91 163.367
R338 B.n266 B.n91 163.367
R339 B.n267 B.n266 163.367
R340 B.n268 B.n267 163.367
R341 B.n268 B.n89 163.367
R342 B.n272 B.n89 163.367
R343 B.n273 B.n272 163.367
R344 B.n274 B.n273 163.367
R345 B.n274 B.n87 163.367
R346 B.n278 B.n87 163.367
R347 B.n279 B.n278 163.367
R348 B.n280 B.n279 163.367
R349 B.n280 B.n85 163.367
R350 B.n284 B.n85 163.367
R351 B.n285 B.n284 163.367
R352 B.n286 B.n285 163.367
R353 B.n286 B.n83 163.367
R354 B.n290 B.n83 163.367
R355 B.n291 B.n290 163.367
R356 B.n292 B.n291 163.367
R357 B.n292 B.n81 163.367
R358 B.n296 B.n81 163.367
R359 B.n297 B.n296 163.367
R360 B.n357 B.n356 163.367
R361 B.n356 B.n61 163.367
R362 B.n352 B.n61 163.367
R363 B.n352 B.n351 163.367
R364 B.n351 B.n350 163.367
R365 B.n350 B.n63 163.367
R366 B.n346 B.n63 163.367
R367 B.n346 B.n345 163.367
R368 B.n345 B.n344 163.367
R369 B.n344 B.n65 163.367
R370 B.n340 B.n65 163.367
R371 B.n340 B.n339 163.367
R372 B.n339 B.n338 163.367
R373 B.n338 B.n67 163.367
R374 B.n334 B.n67 163.367
R375 B.n334 B.n333 163.367
R376 B.n333 B.n332 163.367
R377 B.n332 B.n69 163.367
R378 B.n328 B.n69 163.367
R379 B.n328 B.n327 163.367
R380 B.n327 B.n326 163.367
R381 B.n326 B.n71 163.367
R382 B.n322 B.n71 163.367
R383 B.n322 B.n321 163.367
R384 B.n321 B.n320 163.367
R385 B.n320 B.n73 163.367
R386 B.n316 B.n73 163.367
R387 B.n316 B.n315 163.367
R388 B.n315 B.n314 163.367
R389 B.n314 B.n75 163.367
R390 B.n310 B.n75 163.367
R391 B.n310 B.n309 163.367
R392 B.n309 B.n308 163.367
R393 B.n308 B.n77 163.367
R394 B.n304 B.n77 163.367
R395 B.n304 B.n303 163.367
R396 B.n303 B.n302 163.367
R397 B.n302 B.n79 163.367
R398 B.n298 B.n79 163.367
R399 B.n490 B.n489 163.367
R400 B.n489 B.n488 163.367
R401 B.n488 B.n13 163.367
R402 B.n484 B.n13 163.367
R403 B.n484 B.n483 163.367
R404 B.n483 B.n482 163.367
R405 B.n482 B.n15 163.367
R406 B.n478 B.n15 163.367
R407 B.n478 B.n477 163.367
R408 B.n477 B.n476 163.367
R409 B.n476 B.n17 163.367
R410 B.n472 B.n17 163.367
R411 B.n472 B.n471 163.367
R412 B.n471 B.n470 163.367
R413 B.n470 B.n19 163.367
R414 B.n466 B.n19 163.367
R415 B.n466 B.n465 163.367
R416 B.n465 B.n464 163.367
R417 B.n464 B.n21 163.367
R418 B.n460 B.n21 163.367
R419 B.n460 B.n459 163.367
R420 B.n459 B.n458 163.367
R421 B.n458 B.n23 163.367
R422 B.n454 B.n23 163.367
R423 B.n454 B.n453 163.367
R424 B.n453 B.n452 163.367
R425 B.n452 B.n25 163.367
R426 B.n448 B.n25 163.367
R427 B.n448 B.n447 163.367
R428 B.n447 B.n446 163.367
R429 B.n446 B.n27 163.367
R430 B.n442 B.n27 163.367
R431 B.n442 B.n441 163.367
R432 B.n441 B.n440 163.367
R433 B.n440 B.n29 163.367
R434 B.n436 B.n29 163.367
R435 B.n436 B.n435 163.367
R436 B.n435 B.n434 163.367
R437 B.n434 B.n31 163.367
R438 B.n429 B.n31 163.367
R439 B.n429 B.n428 163.367
R440 B.n428 B.n427 163.367
R441 B.n427 B.n35 163.367
R442 B.n423 B.n35 163.367
R443 B.n423 B.n422 163.367
R444 B.n422 B.n421 163.367
R445 B.n421 B.n37 163.367
R446 B.n417 B.n37 163.367
R447 B.n417 B.n416 163.367
R448 B.n416 B.n41 163.367
R449 B.n412 B.n41 163.367
R450 B.n412 B.n411 163.367
R451 B.n411 B.n410 163.367
R452 B.n410 B.n43 163.367
R453 B.n406 B.n43 163.367
R454 B.n406 B.n405 163.367
R455 B.n405 B.n404 163.367
R456 B.n404 B.n45 163.367
R457 B.n400 B.n45 163.367
R458 B.n400 B.n399 163.367
R459 B.n399 B.n398 163.367
R460 B.n398 B.n47 163.367
R461 B.n394 B.n47 163.367
R462 B.n394 B.n393 163.367
R463 B.n393 B.n392 163.367
R464 B.n392 B.n49 163.367
R465 B.n388 B.n49 163.367
R466 B.n388 B.n387 163.367
R467 B.n387 B.n386 163.367
R468 B.n386 B.n51 163.367
R469 B.n382 B.n51 163.367
R470 B.n382 B.n381 163.367
R471 B.n381 B.n380 163.367
R472 B.n380 B.n53 163.367
R473 B.n376 B.n53 163.367
R474 B.n376 B.n375 163.367
R475 B.n375 B.n374 163.367
R476 B.n374 B.n55 163.367
R477 B.n370 B.n55 163.367
R478 B.n370 B.n369 163.367
R479 B.n369 B.n368 163.367
R480 B.n368 B.n57 163.367
R481 B.n364 B.n57 163.367
R482 B.n364 B.n363 163.367
R483 B.n363 B.n362 163.367
R484 B.n362 B.n59 163.367
R485 B.n358 B.n59 163.367
R486 B.n494 B.n11 163.367
R487 B.n495 B.n494 163.367
R488 B.n496 B.n495 163.367
R489 B.n496 B.n9 163.367
R490 B.n500 B.n9 163.367
R491 B.n501 B.n500 163.367
R492 B.n502 B.n501 163.367
R493 B.n502 B.n7 163.367
R494 B.n506 B.n7 163.367
R495 B.n507 B.n506 163.367
R496 B.n508 B.n507 163.367
R497 B.n508 B.n5 163.367
R498 B.n512 B.n5 163.367
R499 B.n513 B.n512 163.367
R500 B.n514 B.n513 163.367
R501 B.n514 B.n3 163.367
R502 B.n518 B.n3 163.367
R503 B.n519 B.n518 163.367
R504 B.n136 B.n2 163.367
R505 B.n137 B.n136 163.367
R506 B.n138 B.n137 163.367
R507 B.n138 B.n133 163.367
R508 B.n142 B.n133 163.367
R509 B.n143 B.n142 163.367
R510 B.n144 B.n143 163.367
R511 B.n144 B.n131 163.367
R512 B.n148 B.n131 163.367
R513 B.n149 B.n148 163.367
R514 B.n150 B.n149 163.367
R515 B.n150 B.n129 163.367
R516 B.n154 B.n129 163.367
R517 B.n155 B.n154 163.367
R518 B.n156 B.n155 163.367
R519 B.n156 B.n127 163.367
R520 B.n160 B.n127 163.367
R521 B.n161 B.n160 163.367
R522 B.n221 B.n220 59.5399
R523 B.n239 B.n101 59.5399
R524 B.n40 B.n39 59.5399
R525 B.n432 B.n33 59.5399
R526 B.n220 B.n219 38.4005
R527 B.n101 B.n100 38.4005
R528 B.n39 B.n38 38.4005
R529 B.n33 B.n32 38.4005
R530 B.n492 B.n491 37.3078
R531 B.n359 B.n60 37.3078
R532 B.n299 B.n80 37.3078
R533 B.n163 B.n126 37.3078
R534 B B.n521 18.0485
R535 B.n493 B.n492 10.6151
R536 B.n493 B.n10 10.6151
R537 B.n497 B.n10 10.6151
R538 B.n498 B.n497 10.6151
R539 B.n499 B.n498 10.6151
R540 B.n499 B.n8 10.6151
R541 B.n503 B.n8 10.6151
R542 B.n504 B.n503 10.6151
R543 B.n505 B.n504 10.6151
R544 B.n505 B.n6 10.6151
R545 B.n509 B.n6 10.6151
R546 B.n510 B.n509 10.6151
R547 B.n511 B.n510 10.6151
R548 B.n511 B.n4 10.6151
R549 B.n515 B.n4 10.6151
R550 B.n516 B.n515 10.6151
R551 B.n517 B.n516 10.6151
R552 B.n517 B.n0 10.6151
R553 B.n491 B.n12 10.6151
R554 B.n487 B.n12 10.6151
R555 B.n487 B.n486 10.6151
R556 B.n486 B.n485 10.6151
R557 B.n485 B.n14 10.6151
R558 B.n481 B.n14 10.6151
R559 B.n481 B.n480 10.6151
R560 B.n480 B.n479 10.6151
R561 B.n479 B.n16 10.6151
R562 B.n475 B.n16 10.6151
R563 B.n475 B.n474 10.6151
R564 B.n474 B.n473 10.6151
R565 B.n473 B.n18 10.6151
R566 B.n469 B.n18 10.6151
R567 B.n469 B.n468 10.6151
R568 B.n468 B.n467 10.6151
R569 B.n467 B.n20 10.6151
R570 B.n463 B.n20 10.6151
R571 B.n463 B.n462 10.6151
R572 B.n462 B.n461 10.6151
R573 B.n461 B.n22 10.6151
R574 B.n457 B.n22 10.6151
R575 B.n457 B.n456 10.6151
R576 B.n456 B.n455 10.6151
R577 B.n455 B.n24 10.6151
R578 B.n451 B.n24 10.6151
R579 B.n451 B.n450 10.6151
R580 B.n450 B.n449 10.6151
R581 B.n449 B.n26 10.6151
R582 B.n445 B.n26 10.6151
R583 B.n445 B.n444 10.6151
R584 B.n444 B.n443 10.6151
R585 B.n443 B.n28 10.6151
R586 B.n439 B.n28 10.6151
R587 B.n439 B.n438 10.6151
R588 B.n438 B.n437 10.6151
R589 B.n437 B.n30 10.6151
R590 B.n433 B.n30 10.6151
R591 B.n431 B.n430 10.6151
R592 B.n430 B.n34 10.6151
R593 B.n426 B.n34 10.6151
R594 B.n426 B.n425 10.6151
R595 B.n425 B.n424 10.6151
R596 B.n424 B.n36 10.6151
R597 B.n420 B.n36 10.6151
R598 B.n420 B.n419 10.6151
R599 B.n419 B.n418 10.6151
R600 B.n415 B.n414 10.6151
R601 B.n414 B.n413 10.6151
R602 B.n413 B.n42 10.6151
R603 B.n409 B.n42 10.6151
R604 B.n409 B.n408 10.6151
R605 B.n408 B.n407 10.6151
R606 B.n407 B.n44 10.6151
R607 B.n403 B.n44 10.6151
R608 B.n403 B.n402 10.6151
R609 B.n402 B.n401 10.6151
R610 B.n401 B.n46 10.6151
R611 B.n397 B.n46 10.6151
R612 B.n397 B.n396 10.6151
R613 B.n396 B.n395 10.6151
R614 B.n395 B.n48 10.6151
R615 B.n391 B.n48 10.6151
R616 B.n391 B.n390 10.6151
R617 B.n390 B.n389 10.6151
R618 B.n389 B.n50 10.6151
R619 B.n385 B.n50 10.6151
R620 B.n385 B.n384 10.6151
R621 B.n384 B.n383 10.6151
R622 B.n383 B.n52 10.6151
R623 B.n379 B.n52 10.6151
R624 B.n379 B.n378 10.6151
R625 B.n378 B.n377 10.6151
R626 B.n377 B.n54 10.6151
R627 B.n373 B.n54 10.6151
R628 B.n373 B.n372 10.6151
R629 B.n372 B.n371 10.6151
R630 B.n371 B.n56 10.6151
R631 B.n367 B.n56 10.6151
R632 B.n367 B.n366 10.6151
R633 B.n366 B.n365 10.6151
R634 B.n365 B.n58 10.6151
R635 B.n361 B.n58 10.6151
R636 B.n361 B.n360 10.6151
R637 B.n360 B.n359 10.6151
R638 B.n355 B.n60 10.6151
R639 B.n355 B.n354 10.6151
R640 B.n354 B.n353 10.6151
R641 B.n353 B.n62 10.6151
R642 B.n349 B.n62 10.6151
R643 B.n349 B.n348 10.6151
R644 B.n348 B.n347 10.6151
R645 B.n347 B.n64 10.6151
R646 B.n343 B.n64 10.6151
R647 B.n343 B.n342 10.6151
R648 B.n342 B.n341 10.6151
R649 B.n341 B.n66 10.6151
R650 B.n337 B.n66 10.6151
R651 B.n337 B.n336 10.6151
R652 B.n336 B.n335 10.6151
R653 B.n335 B.n68 10.6151
R654 B.n331 B.n68 10.6151
R655 B.n331 B.n330 10.6151
R656 B.n330 B.n329 10.6151
R657 B.n329 B.n70 10.6151
R658 B.n325 B.n70 10.6151
R659 B.n325 B.n324 10.6151
R660 B.n324 B.n323 10.6151
R661 B.n323 B.n72 10.6151
R662 B.n319 B.n72 10.6151
R663 B.n319 B.n318 10.6151
R664 B.n318 B.n317 10.6151
R665 B.n317 B.n74 10.6151
R666 B.n313 B.n74 10.6151
R667 B.n313 B.n312 10.6151
R668 B.n312 B.n311 10.6151
R669 B.n311 B.n76 10.6151
R670 B.n307 B.n76 10.6151
R671 B.n307 B.n306 10.6151
R672 B.n306 B.n305 10.6151
R673 B.n305 B.n78 10.6151
R674 B.n301 B.n78 10.6151
R675 B.n301 B.n300 10.6151
R676 B.n300 B.n299 10.6151
R677 B.n135 B.n1 10.6151
R678 B.n135 B.n134 10.6151
R679 B.n139 B.n134 10.6151
R680 B.n140 B.n139 10.6151
R681 B.n141 B.n140 10.6151
R682 B.n141 B.n132 10.6151
R683 B.n145 B.n132 10.6151
R684 B.n146 B.n145 10.6151
R685 B.n147 B.n146 10.6151
R686 B.n147 B.n130 10.6151
R687 B.n151 B.n130 10.6151
R688 B.n152 B.n151 10.6151
R689 B.n153 B.n152 10.6151
R690 B.n153 B.n128 10.6151
R691 B.n157 B.n128 10.6151
R692 B.n158 B.n157 10.6151
R693 B.n159 B.n158 10.6151
R694 B.n159 B.n126 10.6151
R695 B.n164 B.n163 10.6151
R696 B.n165 B.n164 10.6151
R697 B.n165 B.n124 10.6151
R698 B.n169 B.n124 10.6151
R699 B.n170 B.n169 10.6151
R700 B.n171 B.n170 10.6151
R701 B.n171 B.n122 10.6151
R702 B.n175 B.n122 10.6151
R703 B.n176 B.n175 10.6151
R704 B.n177 B.n176 10.6151
R705 B.n177 B.n120 10.6151
R706 B.n181 B.n120 10.6151
R707 B.n182 B.n181 10.6151
R708 B.n183 B.n182 10.6151
R709 B.n183 B.n118 10.6151
R710 B.n187 B.n118 10.6151
R711 B.n188 B.n187 10.6151
R712 B.n189 B.n188 10.6151
R713 B.n189 B.n116 10.6151
R714 B.n193 B.n116 10.6151
R715 B.n194 B.n193 10.6151
R716 B.n195 B.n194 10.6151
R717 B.n195 B.n114 10.6151
R718 B.n199 B.n114 10.6151
R719 B.n200 B.n199 10.6151
R720 B.n201 B.n200 10.6151
R721 B.n201 B.n112 10.6151
R722 B.n205 B.n112 10.6151
R723 B.n206 B.n205 10.6151
R724 B.n207 B.n206 10.6151
R725 B.n207 B.n110 10.6151
R726 B.n211 B.n110 10.6151
R727 B.n212 B.n211 10.6151
R728 B.n213 B.n212 10.6151
R729 B.n213 B.n108 10.6151
R730 B.n217 B.n108 10.6151
R731 B.n218 B.n217 10.6151
R732 B.n222 B.n218 10.6151
R733 B.n226 B.n106 10.6151
R734 B.n227 B.n226 10.6151
R735 B.n228 B.n227 10.6151
R736 B.n228 B.n104 10.6151
R737 B.n232 B.n104 10.6151
R738 B.n233 B.n232 10.6151
R739 B.n234 B.n233 10.6151
R740 B.n234 B.n102 10.6151
R741 B.n238 B.n102 10.6151
R742 B.n241 B.n240 10.6151
R743 B.n241 B.n98 10.6151
R744 B.n245 B.n98 10.6151
R745 B.n246 B.n245 10.6151
R746 B.n247 B.n246 10.6151
R747 B.n247 B.n96 10.6151
R748 B.n251 B.n96 10.6151
R749 B.n252 B.n251 10.6151
R750 B.n253 B.n252 10.6151
R751 B.n253 B.n94 10.6151
R752 B.n257 B.n94 10.6151
R753 B.n258 B.n257 10.6151
R754 B.n259 B.n258 10.6151
R755 B.n259 B.n92 10.6151
R756 B.n263 B.n92 10.6151
R757 B.n264 B.n263 10.6151
R758 B.n265 B.n264 10.6151
R759 B.n265 B.n90 10.6151
R760 B.n269 B.n90 10.6151
R761 B.n270 B.n269 10.6151
R762 B.n271 B.n270 10.6151
R763 B.n271 B.n88 10.6151
R764 B.n275 B.n88 10.6151
R765 B.n276 B.n275 10.6151
R766 B.n277 B.n276 10.6151
R767 B.n277 B.n86 10.6151
R768 B.n281 B.n86 10.6151
R769 B.n282 B.n281 10.6151
R770 B.n283 B.n282 10.6151
R771 B.n283 B.n84 10.6151
R772 B.n287 B.n84 10.6151
R773 B.n288 B.n287 10.6151
R774 B.n289 B.n288 10.6151
R775 B.n289 B.n82 10.6151
R776 B.n293 B.n82 10.6151
R777 B.n294 B.n293 10.6151
R778 B.n295 B.n294 10.6151
R779 B.n295 B.n80 10.6151
R780 B.n433 B.n432 9.36635
R781 B.n415 B.n40 9.36635
R782 B.n222 B.n221 9.36635
R783 B.n240 B.n239 9.36635
R784 B.n521 B.n0 8.11757
R785 B.n521 B.n1 8.11757
R786 B.n432 B.n431 1.24928
R787 B.n418 B.n40 1.24928
R788 B.n221 B.n106 1.24928
R789 B.n239 B.n238 1.24928
R790 VN VN.t0 264.94
R791 VN VN.t1 223.421
R792 VTAIL.n246 VTAIL.n245 756.745
R793 VTAIL.n60 VTAIL.n59 756.745
R794 VTAIL.n184 VTAIL.n183 756.745
R795 VTAIL.n122 VTAIL.n121 756.745
R796 VTAIL.n207 VTAIL.n206 585
R797 VTAIL.n204 VTAIL.n203 585
R798 VTAIL.n213 VTAIL.n212 585
R799 VTAIL.n215 VTAIL.n214 585
R800 VTAIL.n200 VTAIL.n199 585
R801 VTAIL.n221 VTAIL.n220 585
R802 VTAIL.n223 VTAIL.n222 585
R803 VTAIL.n196 VTAIL.n195 585
R804 VTAIL.n229 VTAIL.n228 585
R805 VTAIL.n231 VTAIL.n230 585
R806 VTAIL.n192 VTAIL.n191 585
R807 VTAIL.n237 VTAIL.n236 585
R808 VTAIL.n239 VTAIL.n238 585
R809 VTAIL.n188 VTAIL.n187 585
R810 VTAIL.n245 VTAIL.n244 585
R811 VTAIL.n21 VTAIL.n20 585
R812 VTAIL.n18 VTAIL.n17 585
R813 VTAIL.n27 VTAIL.n26 585
R814 VTAIL.n29 VTAIL.n28 585
R815 VTAIL.n14 VTAIL.n13 585
R816 VTAIL.n35 VTAIL.n34 585
R817 VTAIL.n37 VTAIL.n36 585
R818 VTAIL.n10 VTAIL.n9 585
R819 VTAIL.n43 VTAIL.n42 585
R820 VTAIL.n45 VTAIL.n44 585
R821 VTAIL.n6 VTAIL.n5 585
R822 VTAIL.n51 VTAIL.n50 585
R823 VTAIL.n53 VTAIL.n52 585
R824 VTAIL.n2 VTAIL.n1 585
R825 VTAIL.n59 VTAIL.n58 585
R826 VTAIL.n183 VTAIL.n182 585
R827 VTAIL.n126 VTAIL.n125 585
R828 VTAIL.n177 VTAIL.n176 585
R829 VTAIL.n175 VTAIL.n174 585
R830 VTAIL.n130 VTAIL.n129 585
R831 VTAIL.n169 VTAIL.n168 585
R832 VTAIL.n167 VTAIL.n166 585
R833 VTAIL.n134 VTAIL.n133 585
R834 VTAIL.n161 VTAIL.n160 585
R835 VTAIL.n159 VTAIL.n158 585
R836 VTAIL.n138 VTAIL.n137 585
R837 VTAIL.n153 VTAIL.n152 585
R838 VTAIL.n151 VTAIL.n150 585
R839 VTAIL.n142 VTAIL.n141 585
R840 VTAIL.n145 VTAIL.n144 585
R841 VTAIL.n121 VTAIL.n120 585
R842 VTAIL.n64 VTAIL.n63 585
R843 VTAIL.n115 VTAIL.n114 585
R844 VTAIL.n113 VTAIL.n112 585
R845 VTAIL.n68 VTAIL.n67 585
R846 VTAIL.n107 VTAIL.n106 585
R847 VTAIL.n105 VTAIL.n104 585
R848 VTAIL.n72 VTAIL.n71 585
R849 VTAIL.n99 VTAIL.n98 585
R850 VTAIL.n97 VTAIL.n96 585
R851 VTAIL.n76 VTAIL.n75 585
R852 VTAIL.n91 VTAIL.n90 585
R853 VTAIL.n89 VTAIL.n88 585
R854 VTAIL.n80 VTAIL.n79 585
R855 VTAIL.n83 VTAIL.n82 585
R856 VTAIL.t2 VTAIL.n205 327.466
R857 VTAIL.t0 VTAIL.n19 327.466
R858 VTAIL.t1 VTAIL.n143 327.466
R859 VTAIL.t3 VTAIL.n81 327.466
R860 VTAIL.n206 VTAIL.n203 171.744
R861 VTAIL.n213 VTAIL.n203 171.744
R862 VTAIL.n214 VTAIL.n213 171.744
R863 VTAIL.n214 VTAIL.n199 171.744
R864 VTAIL.n221 VTAIL.n199 171.744
R865 VTAIL.n222 VTAIL.n221 171.744
R866 VTAIL.n222 VTAIL.n195 171.744
R867 VTAIL.n229 VTAIL.n195 171.744
R868 VTAIL.n230 VTAIL.n229 171.744
R869 VTAIL.n230 VTAIL.n191 171.744
R870 VTAIL.n237 VTAIL.n191 171.744
R871 VTAIL.n238 VTAIL.n237 171.744
R872 VTAIL.n238 VTAIL.n187 171.744
R873 VTAIL.n245 VTAIL.n187 171.744
R874 VTAIL.n20 VTAIL.n17 171.744
R875 VTAIL.n27 VTAIL.n17 171.744
R876 VTAIL.n28 VTAIL.n27 171.744
R877 VTAIL.n28 VTAIL.n13 171.744
R878 VTAIL.n35 VTAIL.n13 171.744
R879 VTAIL.n36 VTAIL.n35 171.744
R880 VTAIL.n36 VTAIL.n9 171.744
R881 VTAIL.n43 VTAIL.n9 171.744
R882 VTAIL.n44 VTAIL.n43 171.744
R883 VTAIL.n44 VTAIL.n5 171.744
R884 VTAIL.n51 VTAIL.n5 171.744
R885 VTAIL.n52 VTAIL.n51 171.744
R886 VTAIL.n52 VTAIL.n1 171.744
R887 VTAIL.n59 VTAIL.n1 171.744
R888 VTAIL.n183 VTAIL.n125 171.744
R889 VTAIL.n176 VTAIL.n125 171.744
R890 VTAIL.n176 VTAIL.n175 171.744
R891 VTAIL.n175 VTAIL.n129 171.744
R892 VTAIL.n168 VTAIL.n129 171.744
R893 VTAIL.n168 VTAIL.n167 171.744
R894 VTAIL.n167 VTAIL.n133 171.744
R895 VTAIL.n160 VTAIL.n133 171.744
R896 VTAIL.n160 VTAIL.n159 171.744
R897 VTAIL.n159 VTAIL.n137 171.744
R898 VTAIL.n152 VTAIL.n137 171.744
R899 VTAIL.n152 VTAIL.n151 171.744
R900 VTAIL.n151 VTAIL.n141 171.744
R901 VTAIL.n144 VTAIL.n141 171.744
R902 VTAIL.n121 VTAIL.n63 171.744
R903 VTAIL.n114 VTAIL.n63 171.744
R904 VTAIL.n114 VTAIL.n113 171.744
R905 VTAIL.n113 VTAIL.n67 171.744
R906 VTAIL.n106 VTAIL.n67 171.744
R907 VTAIL.n106 VTAIL.n105 171.744
R908 VTAIL.n105 VTAIL.n71 171.744
R909 VTAIL.n98 VTAIL.n71 171.744
R910 VTAIL.n98 VTAIL.n97 171.744
R911 VTAIL.n97 VTAIL.n75 171.744
R912 VTAIL.n90 VTAIL.n75 171.744
R913 VTAIL.n90 VTAIL.n89 171.744
R914 VTAIL.n89 VTAIL.n79 171.744
R915 VTAIL.n82 VTAIL.n79 171.744
R916 VTAIL.n206 VTAIL.t2 85.8723
R917 VTAIL.n20 VTAIL.t0 85.8723
R918 VTAIL.n144 VTAIL.t1 85.8723
R919 VTAIL.n82 VTAIL.t3 85.8723
R920 VTAIL.n247 VTAIL.n246 34.3187
R921 VTAIL.n61 VTAIL.n60 34.3187
R922 VTAIL.n185 VTAIL.n184 34.3187
R923 VTAIL.n123 VTAIL.n122 34.3187
R924 VTAIL.n123 VTAIL.n61 25.4789
R925 VTAIL.n247 VTAIL.n185 23.7721
R926 VTAIL.n207 VTAIL.n205 16.3895
R927 VTAIL.n21 VTAIL.n19 16.3895
R928 VTAIL.n145 VTAIL.n143 16.3895
R929 VTAIL.n83 VTAIL.n81 16.3895
R930 VTAIL.n208 VTAIL.n204 12.8005
R931 VTAIL.n22 VTAIL.n18 12.8005
R932 VTAIL.n146 VTAIL.n142 12.8005
R933 VTAIL.n84 VTAIL.n80 12.8005
R934 VTAIL.n212 VTAIL.n211 12.0247
R935 VTAIL.n26 VTAIL.n25 12.0247
R936 VTAIL.n150 VTAIL.n149 12.0247
R937 VTAIL.n88 VTAIL.n87 12.0247
R938 VTAIL.n215 VTAIL.n202 11.249
R939 VTAIL.n244 VTAIL.n186 11.249
R940 VTAIL.n29 VTAIL.n16 11.249
R941 VTAIL.n58 VTAIL.n0 11.249
R942 VTAIL.n182 VTAIL.n124 11.249
R943 VTAIL.n153 VTAIL.n140 11.249
R944 VTAIL.n120 VTAIL.n62 11.249
R945 VTAIL.n91 VTAIL.n78 11.249
R946 VTAIL.n216 VTAIL.n200 10.4732
R947 VTAIL.n243 VTAIL.n188 10.4732
R948 VTAIL.n30 VTAIL.n14 10.4732
R949 VTAIL.n57 VTAIL.n2 10.4732
R950 VTAIL.n181 VTAIL.n126 10.4732
R951 VTAIL.n154 VTAIL.n138 10.4732
R952 VTAIL.n119 VTAIL.n64 10.4732
R953 VTAIL.n92 VTAIL.n76 10.4732
R954 VTAIL.n220 VTAIL.n219 9.69747
R955 VTAIL.n240 VTAIL.n239 9.69747
R956 VTAIL.n34 VTAIL.n33 9.69747
R957 VTAIL.n54 VTAIL.n53 9.69747
R958 VTAIL.n178 VTAIL.n177 9.69747
R959 VTAIL.n158 VTAIL.n157 9.69747
R960 VTAIL.n116 VTAIL.n115 9.69747
R961 VTAIL.n96 VTAIL.n95 9.69747
R962 VTAIL.n242 VTAIL.n186 9.45567
R963 VTAIL.n56 VTAIL.n0 9.45567
R964 VTAIL.n180 VTAIL.n124 9.45567
R965 VTAIL.n118 VTAIL.n62 9.45567
R966 VTAIL.n194 VTAIL.n193 9.3005
R967 VTAIL.n233 VTAIL.n232 9.3005
R968 VTAIL.n235 VTAIL.n234 9.3005
R969 VTAIL.n190 VTAIL.n189 9.3005
R970 VTAIL.n241 VTAIL.n240 9.3005
R971 VTAIL.n243 VTAIL.n242 9.3005
R972 VTAIL.n225 VTAIL.n224 9.3005
R973 VTAIL.n198 VTAIL.n197 9.3005
R974 VTAIL.n219 VTAIL.n218 9.3005
R975 VTAIL.n217 VTAIL.n216 9.3005
R976 VTAIL.n202 VTAIL.n201 9.3005
R977 VTAIL.n211 VTAIL.n210 9.3005
R978 VTAIL.n209 VTAIL.n208 9.3005
R979 VTAIL.n227 VTAIL.n226 9.3005
R980 VTAIL.n8 VTAIL.n7 9.3005
R981 VTAIL.n47 VTAIL.n46 9.3005
R982 VTAIL.n49 VTAIL.n48 9.3005
R983 VTAIL.n4 VTAIL.n3 9.3005
R984 VTAIL.n55 VTAIL.n54 9.3005
R985 VTAIL.n57 VTAIL.n56 9.3005
R986 VTAIL.n39 VTAIL.n38 9.3005
R987 VTAIL.n12 VTAIL.n11 9.3005
R988 VTAIL.n33 VTAIL.n32 9.3005
R989 VTAIL.n31 VTAIL.n30 9.3005
R990 VTAIL.n16 VTAIL.n15 9.3005
R991 VTAIL.n25 VTAIL.n24 9.3005
R992 VTAIL.n23 VTAIL.n22 9.3005
R993 VTAIL.n41 VTAIL.n40 9.3005
R994 VTAIL.n181 VTAIL.n180 9.3005
R995 VTAIL.n179 VTAIL.n178 9.3005
R996 VTAIL.n128 VTAIL.n127 9.3005
R997 VTAIL.n173 VTAIL.n172 9.3005
R998 VTAIL.n171 VTAIL.n170 9.3005
R999 VTAIL.n132 VTAIL.n131 9.3005
R1000 VTAIL.n165 VTAIL.n164 9.3005
R1001 VTAIL.n163 VTAIL.n162 9.3005
R1002 VTAIL.n136 VTAIL.n135 9.3005
R1003 VTAIL.n157 VTAIL.n156 9.3005
R1004 VTAIL.n155 VTAIL.n154 9.3005
R1005 VTAIL.n140 VTAIL.n139 9.3005
R1006 VTAIL.n149 VTAIL.n148 9.3005
R1007 VTAIL.n147 VTAIL.n146 9.3005
R1008 VTAIL.n109 VTAIL.n108 9.3005
R1009 VTAIL.n111 VTAIL.n110 9.3005
R1010 VTAIL.n66 VTAIL.n65 9.3005
R1011 VTAIL.n117 VTAIL.n116 9.3005
R1012 VTAIL.n119 VTAIL.n118 9.3005
R1013 VTAIL.n70 VTAIL.n69 9.3005
R1014 VTAIL.n103 VTAIL.n102 9.3005
R1015 VTAIL.n101 VTAIL.n100 9.3005
R1016 VTAIL.n74 VTAIL.n73 9.3005
R1017 VTAIL.n95 VTAIL.n94 9.3005
R1018 VTAIL.n93 VTAIL.n92 9.3005
R1019 VTAIL.n78 VTAIL.n77 9.3005
R1020 VTAIL.n87 VTAIL.n86 9.3005
R1021 VTAIL.n85 VTAIL.n84 9.3005
R1022 VTAIL.n223 VTAIL.n198 8.92171
R1023 VTAIL.n236 VTAIL.n190 8.92171
R1024 VTAIL.n37 VTAIL.n12 8.92171
R1025 VTAIL.n50 VTAIL.n4 8.92171
R1026 VTAIL.n174 VTAIL.n128 8.92171
R1027 VTAIL.n161 VTAIL.n136 8.92171
R1028 VTAIL.n112 VTAIL.n66 8.92171
R1029 VTAIL.n99 VTAIL.n74 8.92171
R1030 VTAIL.n224 VTAIL.n196 8.14595
R1031 VTAIL.n235 VTAIL.n192 8.14595
R1032 VTAIL.n38 VTAIL.n10 8.14595
R1033 VTAIL.n49 VTAIL.n6 8.14595
R1034 VTAIL.n173 VTAIL.n130 8.14595
R1035 VTAIL.n162 VTAIL.n134 8.14595
R1036 VTAIL.n111 VTAIL.n68 8.14595
R1037 VTAIL.n100 VTAIL.n72 8.14595
R1038 VTAIL.n228 VTAIL.n227 7.3702
R1039 VTAIL.n232 VTAIL.n231 7.3702
R1040 VTAIL.n42 VTAIL.n41 7.3702
R1041 VTAIL.n46 VTAIL.n45 7.3702
R1042 VTAIL.n170 VTAIL.n169 7.3702
R1043 VTAIL.n166 VTAIL.n165 7.3702
R1044 VTAIL.n108 VTAIL.n107 7.3702
R1045 VTAIL.n104 VTAIL.n103 7.3702
R1046 VTAIL.n228 VTAIL.n194 6.59444
R1047 VTAIL.n231 VTAIL.n194 6.59444
R1048 VTAIL.n42 VTAIL.n8 6.59444
R1049 VTAIL.n45 VTAIL.n8 6.59444
R1050 VTAIL.n169 VTAIL.n132 6.59444
R1051 VTAIL.n166 VTAIL.n132 6.59444
R1052 VTAIL.n107 VTAIL.n70 6.59444
R1053 VTAIL.n104 VTAIL.n70 6.59444
R1054 VTAIL.n227 VTAIL.n196 5.81868
R1055 VTAIL.n232 VTAIL.n192 5.81868
R1056 VTAIL.n41 VTAIL.n10 5.81868
R1057 VTAIL.n46 VTAIL.n6 5.81868
R1058 VTAIL.n170 VTAIL.n130 5.81868
R1059 VTAIL.n165 VTAIL.n134 5.81868
R1060 VTAIL.n108 VTAIL.n68 5.81868
R1061 VTAIL.n103 VTAIL.n72 5.81868
R1062 VTAIL.n224 VTAIL.n223 5.04292
R1063 VTAIL.n236 VTAIL.n235 5.04292
R1064 VTAIL.n38 VTAIL.n37 5.04292
R1065 VTAIL.n50 VTAIL.n49 5.04292
R1066 VTAIL.n174 VTAIL.n173 5.04292
R1067 VTAIL.n162 VTAIL.n161 5.04292
R1068 VTAIL.n112 VTAIL.n111 5.04292
R1069 VTAIL.n100 VTAIL.n99 5.04292
R1070 VTAIL.n220 VTAIL.n198 4.26717
R1071 VTAIL.n239 VTAIL.n190 4.26717
R1072 VTAIL.n34 VTAIL.n12 4.26717
R1073 VTAIL.n53 VTAIL.n4 4.26717
R1074 VTAIL.n177 VTAIL.n128 4.26717
R1075 VTAIL.n158 VTAIL.n136 4.26717
R1076 VTAIL.n115 VTAIL.n66 4.26717
R1077 VTAIL.n96 VTAIL.n74 4.26717
R1078 VTAIL.n209 VTAIL.n205 3.70982
R1079 VTAIL.n23 VTAIL.n19 3.70982
R1080 VTAIL.n147 VTAIL.n143 3.70982
R1081 VTAIL.n85 VTAIL.n81 3.70982
R1082 VTAIL.n219 VTAIL.n200 3.49141
R1083 VTAIL.n240 VTAIL.n188 3.49141
R1084 VTAIL.n33 VTAIL.n14 3.49141
R1085 VTAIL.n54 VTAIL.n2 3.49141
R1086 VTAIL.n178 VTAIL.n126 3.49141
R1087 VTAIL.n157 VTAIL.n138 3.49141
R1088 VTAIL.n116 VTAIL.n64 3.49141
R1089 VTAIL.n95 VTAIL.n76 3.49141
R1090 VTAIL.n216 VTAIL.n215 2.71565
R1091 VTAIL.n244 VTAIL.n243 2.71565
R1092 VTAIL.n30 VTAIL.n29 2.71565
R1093 VTAIL.n58 VTAIL.n57 2.71565
R1094 VTAIL.n182 VTAIL.n181 2.71565
R1095 VTAIL.n154 VTAIL.n153 2.71565
R1096 VTAIL.n120 VTAIL.n119 2.71565
R1097 VTAIL.n92 VTAIL.n91 2.71565
R1098 VTAIL.n212 VTAIL.n202 1.93989
R1099 VTAIL.n246 VTAIL.n186 1.93989
R1100 VTAIL.n26 VTAIL.n16 1.93989
R1101 VTAIL.n60 VTAIL.n0 1.93989
R1102 VTAIL.n184 VTAIL.n124 1.93989
R1103 VTAIL.n150 VTAIL.n140 1.93989
R1104 VTAIL.n122 VTAIL.n62 1.93989
R1105 VTAIL.n88 VTAIL.n78 1.93989
R1106 VTAIL.n185 VTAIL.n123 1.32378
R1107 VTAIL.n211 VTAIL.n204 1.16414
R1108 VTAIL.n25 VTAIL.n18 1.16414
R1109 VTAIL.n149 VTAIL.n142 1.16414
R1110 VTAIL.n87 VTAIL.n80 1.16414
R1111 VTAIL VTAIL.n61 0.955241
R1112 VTAIL.n208 VTAIL.n207 0.388379
R1113 VTAIL.n22 VTAIL.n21 0.388379
R1114 VTAIL.n146 VTAIL.n145 0.388379
R1115 VTAIL.n84 VTAIL.n83 0.388379
R1116 VTAIL VTAIL.n247 0.369034
R1117 VTAIL.n210 VTAIL.n209 0.155672
R1118 VTAIL.n210 VTAIL.n201 0.155672
R1119 VTAIL.n217 VTAIL.n201 0.155672
R1120 VTAIL.n218 VTAIL.n217 0.155672
R1121 VTAIL.n218 VTAIL.n197 0.155672
R1122 VTAIL.n225 VTAIL.n197 0.155672
R1123 VTAIL.n226 VTAIL.n225 0.155672
R1124 VTAIL.n226 VTAIL.n193 0.155672
R1125 VTAIL.n233 VTAIL.n193 0.155672
R1126 VTAIL.n234 VTAIL.n233 0.155672
R1127 VTAIL.n234 VTAIL.n189 0.155672
R1128 VTAIL.n241 VTAIL.n189 0.155672
R1129 VTAIL.n242 VTAIL.n241 0.155672
R1130 VTAIL.n24 VTAIL.n23 0.155672
R1131 VTAIL.n24 VTAIL.n15 0.155672
R1132 VTAIL.n31 VTAIL.n15 0.155672
R1133 VTAIL.n32 VTAIL.n31 0.155672
R1134 VTAIL.n32 VTAIL.n11 0.155672
R1135 VTAIL.n39 VTAIL.n11 0.155672
R1136 VTAIL.n40 VTAIL.n39 0.155672
R1137 VTAIL.n40 VTAIL.n7 0.155672
R1138 VTAIL.n47 VTAIL.n7 0.155672
R1139 VTAIL.n48 VTAIL.n47 0.155672
R1140 VTAIL.n48 VTAIL.n3 0.155672
R1141 VTAIL.n55 VTAIL.n3 0.155672
R1142 VTAIL.n56 VTAIL.n55 0.155672
R1143 VTAIL.n180 VTAIL.n179 0.155672
R1144 VTAIL.n179 VTAIL.n127 0.155672
R1145 VTAIL.n172 VTAIL.n127 0.155672
R1146 VTAIL.n172 VTAIL.n171 0.155672
R1147 VTAIL.n171 VTAIL.n131 0.155672
R1148 VTAIL.n164 VTAIL.n131 0.155672
R1149 VTAIL.n164 VTAIL.n163 0.155672
R1150 VTAIL.n163 VTAIL.n135 0.155672
R1151 VTAIL.n156 VTAIL.n135 0.155672
R1152 VTAIL.n156 VTAIL.n155 0.155672
R1153 VTAIL.n155 VTAIL.n139 0.155672
R1154 VTAIL.n148 VTAIL.n139 0.155672
R1155 VTAIL.n148 VTAIL.n147 0.155672
R1156 VTAIL.n118 VTAIL.n117 0.155672
R1157 VTAIL.n117 VTAIL.n65 0.155672
R1158 VTAIL.n110 VTAIL.n65 0.155672
R1159 VTAIL.n110 VTAIL.n109 0.155672
R1160 VTAIL.n109 VTAIL.n69 0.155672
R1161 VTAIL.n102 VTAIL.n69 0.155672
R1162 VTAIL.n102 VTAIL.n101 0.155672
R1163 VTAIL.n101 VTAIL.n73 0.155672
R1164 VTAIL.n94 VTAIL.n73 0.155672
R1165 VTAIL.n94 VTAIL.n93 0.155672
R1166 VTAIL.n93 VTAIL.n77 0.155672
R1167 VTAIL.n86 VTAIL.n77 0.155672
R1168 VTAIL.n86 VTAIL.n85 0.155672
R1169 VDD2.n121 VDD2.n120 756.745
R1170 VDD2.n60 VDD2.n59 756.745
R1171 VDD2.n120 VDD2.n119 585
R1172 VDD2.n63 VDD2.n62 585
R1173 VDD2.n114 VDD2.n113 585
R1174 VDD2.n112 VDD2.n111 585
R1175 VDD2.n67 VDD2.n66 585
R1176 VDD2.n106 VDD2.n105 585
R1177 VDD2.n104 VDD2.n103 585
R1178 VDD2.n71 VDD2.n70 585
R1179 VDD2.n98 VDD2.n97 585
R1180 VDD2.n96 VDD2.n95 585
R1181 VDD2.n75 VDD2.n74 585
R1182 VDD2.n90 VDD2.n89 585
R1183 VDD2.n88 VDD2.n87 585
R1184 VDD2.n79 VDD2.n78 585
R1185 VDD2.n82 VDD2.n81 585
R1186 VDD2.n21 VDD2.n20 585
R1187 VDD2.n18 VDD2.n17 585
R1188 VDD2.n27 VDD2.n26 585
R1189 VDD2.n29 VDD2.n28 585
R1190 VDD2.n14 VDD2.n13 585
R1191 VDD2.n35 VDD2.n34 585
R1192 VDD2.n37 VDD2.n36 585
R1193 VDD2.n10 VDD2.n9 585
R1194 VDD2.n43 VDD2.n42 585
R1195 VDD2.n45 VDD2.n44 585
R1196 VDD2.n6 VDD2.n5 585
R1197 VDD2.n51 VDD2.n50 585
R1198 VDD2.n53 VDD2.n52 585
R1199 VDD2.n2 VDD2.n1 585
R1200 VDD2.n59 VDD2.n58 585
R1201 VDD2.t1 VDD2.n80 327.466
R1202 VDD2.t0 VDD2.n19 327.466
R1203 VDD2.n120 VDD2.n62 171.744
R1204 VDD2.n113 VDD2.n62 171.744
R1205 VDD2.n113 VDD2.n112 171.744
R1206 VDD2.n112 VDD2.n66 171.744
R1207 VDD2.n105 VDD2.n66 171.744
R1208 VDD2.n105 VDD2.n104 171.744
R1209 VDD2.n104 VDD2.n70 171.744
R1210 VDD2.n97 VDD2.n70 171.744
R1211 VDD2.n97 VDD2.n96 171.744
R1212 VDD2.n96 VDD2.n74 171.744
R1213 VDD2.n89 VDD2.n74 171.744
R1214 VDD2.n89 VDD2.n88 171.744
R1215 VDD2.n88 VDD2.n78 171.744
R1216 VDD2.n81 VDD2.n78 171.744
R1217 VDD2.n20 VDD2.n17 171.744
R1218 VDD2.n27 VDD2.n17 171.744
R1219 VDD2.n28 VDD2.n27 171.744
R1220 VDD2.n28 VDD2.n13 171.744
R1221 VDD2.n35 VDD2.n13 171.744
R1222 VDD2.n36 VDD2.n35 171.744
R1223 VDD2.n36 VDD2.n9 171.744
R1224 VDD2.n43 VDD2.n9 171.744
R1225 VDD2.n44 VDD2.n43 171.744
R1226 VDD2.n44 VDD2.n5 171.744
R1227 VDD2.n51 VDD2.n5 171.744
R1228 VDD2.n52 VDD2.n51 171.744
R1229 VDD2.n52 VDD2.n1 171.744
R1230 VDD2.n59 VDD2.n1 171.744
R1231 VDD2.n122 VDD2.n60 87.769
R1232 VDD2.n81 VDD2.t1 85.8723
R1233 VDD2.n20 VDD2.t0 85.8723
R1234 VDD2.n122 VDD2.n121 50.9975
R1235 VDD2.n82 VDD2.n80 16.3895
R1236 VDD2.n21 VDD2.n19 16.3895
R1237 VDD2.n83 VDD2.n79 12.8005
R1238 VDD2.n22 VDD2.n18 12.8005
R1239 VDD2.n87 VDD2.n86 12.0247
R1240 VDD2.n26 VDD2.n25 12.0247
R1241 VDD2.n119 VDD2.n61 11.249
R1242 VDD2.n90 VDD2.n77 11.249
R1243 VDD2.n29 VDD2.n16 11.249
R1244 VDD2.n58 VDD2.n0 11.249
R1245 VDD2.n118 VDD2.n63 10.4732
R1246 VDD2.n91 VDD2.n75 10.4732
R1247 VDD2.n30 VDD2.n14 10.4732
R1248 VDD2.n57 VDD2.n2 10.4732
R1249 VDD2.n115 VDD2.n114 9.69747
R1250 VDD2.n95 VDD2.n94 9.69747
R1251 VDD2.n34 VDD2.n33 9.69747
R1252 VDD2.n54 VDD2.n53 9.69747
R1253 VDD2.n117 VDD2.n61 9.45567
R1254 VDD2.n56 VDD2.n0 9.45567
R1255 VDD2.n118 VDD2.n117 9.3005
R1256 VDD2.n116 VDD2.n115 9.3005
R1257 VDD2.n65 VDD2.n64 9.3005
R1258 VDD2.n110 VDD2.n109 9.3005
R1259 VDD2.n108 VDD2.n107 9.3005
R1260 VDD2.n69 VDD2.n68 9.3005
R1261 VDD2.n102 VDD2.n101 9.3005
R1262 VDD2.n100 VDD2.n99 9.3005
R1263 VDD2.n73 VDD2.n72 9.3005
R1264 VDD2.n94 VDD2.n93 9.3005
R1265 VDD2.n92 VDD2.n91 9.3005
R1266 VDD2.n77 VDD2.n76 9.3005
R1267 VDD2.n86 VDD2.n85 9.3005
R1268 VDD2.n84 VDD2.n83 9.3005
R1269 VDD2.n8 VDD2.n7 9.3005
R1270 VDD2.n47 VDD2.n46 9.3005
R1271 VDD2.n49 VDD2.n48 9.3005
R1272 VDD2.n4 VDD2.n3 9.3005
R1273 VDD2.n55 VDD2.n54 9.3005
R1274 VDD2.n57 VDD2.n56 9.3005
R1275 VDD2.n39 VDD2.n38 9.3005
R1276 VDD2.n12 VDD2.n11 9.3005
R1277 VDD2.n33 VDD2.n32 9.3005
R1278 VDD2.n31 VDD2.n30 9.3005
R1279 VDD2.n16 VDD2.n15 9.3005
R1280 VDD2.n25 VDD2.n24 9.3005
R1281 VDD2.n23 VDD2.n22 9.3005
R1282 VDD2.n41 VDD2.n40 9.3005
R1283 VDD2.n111 VDD2.n65 8.92171
R1284 VDD2.n98 VDD2.n73 8.92171
R1285 VDD2.n37 VDD2.n12 8.92171
R1286 VDD2.n50 VDD2.n4 8.92171
R1287 VDD2.n110 VDD2.n67 8.14595
R1288 VDD2.n99 VDD2.n71 8.14595
R1289 VDD2.n38 VDD2.n10 8.14595
R1290 VDD2.n49 VDD2.n6 8.14595
R1291 VDD2.n107 VDD2.n106 7.3702
R1292 VDD2.n103 VDD2.n102 7.3702
R1293 VDD2.n42 VDD2.n41 7.3702
R1294 VDD2.n46 VDD2.n45 7.3702
R1295 VDD2.n106 VDD2.n69 6.59444
R1296 VDD2.n103 VDD2.n69 6.59444
R1297 VDD2.n42 VDD2.n8 6.59444
R1298 VDD2.n45 VDD2.n8 6.59444
R1299 VDD2.n107 VDD2.n67 5.81868
R1300 VDD2.n102 VDD2.n71 5.81868
R1301 VDD2.n41 VDD2.n10 5.81868
R1302 VDD2.n46 VDD2.n6 5.81868
R1303 VDD2.n111 VDD2.n110 5.04292
R1304 VDD2.n99 VDD2.n98 5.04292
R1305 VDD2.n38 VDD2.n37 5.04292
R1306 VDD2.n50 VDD2.n49 5.04292
R1307 VDD2.n114 VDD2.n65 4.26717
R1308 VDD2.n95 VDD2.n73 4.26717
R1309 VDD2.n34 VDD2.n12 4.26717
R1310 VDD2.n53 VDD2.n4 4.26717
R1311 VDD2.n84 VDD2.n80 3.70982
R1312 VDD2.n23 VDD2.n19 3.70982
R1313 VDD2.n115 VDD2.n63 3.49141
R1314 VDD2.n94 VDD2.n75 3.49141
R1315 VDD2.n33 VDD2.n14 3.49141
R1316 VDD2.n54 VDD2.n2 3.49141
R1317 VDD2.n119 VDD2.n118 2.71565
R1318 VDD2.n91 VDD2.n90 2.71565
R1319 VDD2.n30 VDD2.n29 2.71565
R1320 VDD2.n58 VDD2.n57 2.71565
R1321 VDD2.n121 VDD2.n61 1.93989
R1322 VDD2.n87 VDD2.n77 1.93989
R1323 VDD2.n26 VDD2.n16 1.93989
R1324 VDD2.n60 VDD2.n0 1.93989
R1325 VDD2.n86 VDD2.n79 1.16414
R1326 VDD2.n25 VDD2.n18 1.16414
R1327 VDD2 VDD2.n122 0.485414
R1328 VDD2.n83 VDD2.n82 0.388379
R1329 VDD2.n22 VDD2.n21 0.388379
R1330 VDD2.n117 VDD2.n116 0.155672
R1331 VDD2.n116 VDD2.n64 0.155672
R1332 VDD2.n109 VDD2.n64 0.155672
R1333 VDD2.n109 VDD2.n108 0.155672
R1334 VDD2.n108 VDD2.n68 0.155672
R1335 VDD2.n101 VDD2.n68 0.155672
R1336 VDD2.n101 VDD2.n100 0.155672
R1337 VDD2.n100 VDD2.n72 0.155672
R1338 VDD2.n93 VDD2.n72 0.155672
R1339 VDD2.n93 VDD2.n92 0.155672
R1340 VDD2.n92 VDD2.n76 0.155672
R1341 VDD2.n85 VDD2.n76 0.155672
R1342 VDD2.n85 VDD2.n84 0.155672
R1343 VDD2.n24 VDD2.n23 0.155672
R1344 VDD2.n24 VDD2.n15 0.155672
R1345 VDD2.n31 VDD2.n15 0.155672
R1346 VDD2.n32 VDD2.n31 0.155672
R1347 VDD2.n32 VDD2.n11 0.155672
R1348 VDD2.n39 VDD2.n11 0.155672
R1349 VDD2.n40 VDD2.n39 0.155672
R1350 VDD2.n40 VDD2.n7 0.155672
R1351 VDD2.n47 VDD2.n7 0.155672
R1352 VDD2.n48 VDD2.n47 0.155672
R1353 VDD2.n48 VDD2.n3 0.155672
R1354 VDD2.n55 VDD2.n3 0.155672
R1355 VDD2.n56 VDD2.n55 0.155672
R1356 VP.n0 VP.t1 264.748
R1357 VP.n0 VP.t0 223.179
R1358 VP VP.n0 0.241678
R1359 VDD1.n60 VDD1.n59 756.745
R1360 VDD1.n121 VDD1.n120 756.745
R1361 VDD1.n59 VDD1.n58 585
R1362 VDD1.n2 VDD1.n1 585
R1363 VDD1.n53 VDD1.n52 585
R1364 VDD1.n51 VDD1.n50 585
R1365 VDD1.n6 VDD1.n5 585
R1366 VDD1.n45 VDD1.n44 585
R1367 VDD1.n43 VDD1.n42 585
R1368 VDD1.n10 VDD1.n9 585
R1369 VDD1.n37 VDD1.n36 585
R1370 VDD1.n35 VDD1.n34 585
R1371 VDD1.n14 VDD1.n13 585
R1372 VDD1.n29 VDD1.n28 585
R1373 VDD1.n27 VDD1.n26 585
R1374 VDD1.n18 VDD1.n17 585
R1375 VDD1.n21 VDD1.n20 585
R1376 VDD1.n82 VDD1.n81 585
R1377 VDD1.n79 VDD1.n78 585
R1378 VDD1.n88 VDD1.n87 585
R1379 VDD1.n90 VDD1.n89 585
R1380 VDD1.n75 VDD1.n74 585
R1381 VDD1.n96 VDD1.n95 585
R1382 VDD1.n98 VDD1.n97 585
R1383 VDD1.n71 VDD1.n70 585
R1384 VDD1.n104 VDD1.n103 585
R1385 VDD1.n106 VDD1.n105 585
R1386 VDD1.n67 VDD1.n66 585
R1387 VDD1.n112 VDD1.n111 585
R1388 VDD1.n114 VDD1.n113 585
R1389 VDD1.n63 VDD1.n62 585
R1390 VDD1.n120 VDD1.n119 585
R1391 VDD1.t0 VDD1.n19 327.466
R1392 VDD1.t1 VDD1.n80 327.466
R1393 VDD1.n59 VDD1.n1 171.744
R1394 VDD1.n52 VDD1.n1 171.744
R1395 VDD1.n52 VDD1.n51 171.744
R1396 VDD1.n51 VDD1.n5 171.744
R1397 VDD1.n44 VDD1.n5 171.744
R1398 VDD1.n44 VDD1.n43 171.744
R1399 VDD1.n43 VDD1.n9 171.744
R1400 VDD1.n36 VDD1.n9 171.744
R1401 VDD1.n36 VDD1.n35 171.744
R1402 VDD1.n35 VDD1.n13 171.744
R1403 VDD1.n28 VDD1.n13 171.744
R1404 VDD1.n28 VDD1.n27 171.744
R1405 VDD1.n27 VDD1.n17 171.744
R1406 VDD1.n20 VDD1.n17 171.744
R1407 VDD1.n81 VDD1.n78 171.744
R1408 VDD1.n88 VDD1.n78 171.744
R1409 VDD1.n89 VDD1.n88 171.744
R1410 VDD1.n89 VDD1.n74 171.744
R1411 VDD1.n96 VDD1.n74 171.744
R1412 VDD1.n97 VDD1.n96 171.744
R1413 VDD1.n97 VDD1.n70 171.744
R1414 VDD1.n104 VDD1.n70 171.744
R1415 VDD1.n105 VDD1.n104 171.744
R1416 VDD1.n105 VDD1.n66 171.744
R1417 VDD1.n112 VDD1.n66 171.744
R1418 VDD1.n113 VDD1.n112 171.744
R1419 VDD1.n113 VDD1.n62 171.744
R1420 VDD1.n120 VDD1.n62 171.744
R1421 VDD1 VDD1.n121 88.7205
R1422 VDD1.n20 VDD1.t0 85.8723
R1423 VDD1.n81 VDD1.t1 85.8723
R1424 VDD1 VDD1.n60 51.4824
R1425 VDD1.n21 VDD1.n19 16.3895
R1426 VDD1.n82 VDD1.n80 16.3895
R1427 VDD1.n22 VDD1.n18 12.8005
R1428 VDD1.n83 VDD1.n79 12.8005
R1429 VDD1.n26 VDD1.n25 12.0247
R1430 VDD1.n87 VDD1.n86 12.0247
R1431 VDD1.n58 VDD1.n0 11.249
R1432 VDD1.n29 VDD1.n16 11.249
R1433 VDD1.n90 VDD1.n77 11.249
R1434 VDD1.n119 VDD1.n61 11.249
R1435 VDD1.n57 VDD1.n2 10.4732
R1436 VDD1.n30 VDD1.n14 10.4732
R1437 VDD1.n91 VDD1.n75 10.4732
R1438 VDD1.n118 VDD1.n63 10.4732
R1439 VDD1.n54 VDD1.n53 9.69747
R1440 VDD1.n34 VDD1.n33 9.69747
R1441 VDD1.n95 VDD1.n94 9.69747
R1442 VDD1.n115 VDD1.n114 9.69747
R1443 VDD1.n56 VDD1.n0 9.45567
R1444 VDD1.n117 VDD1.n61 9.45567
R1445 VDD1.n57 VDD1.n56 9.3005
R1446 VDD1.n55 VDD1.n54 9.3005
R1447 VDD1.n4 VDD1.n3 9.3005
R1448 VDD1.n49 VDD1.n48 9.3005
R1449 VDD1.n47 VDD1.n46 9.3005
R1450 VDD1.n8 VDD1.n7 9.3005
R1451 VDD1.n41 VDD1.n40 9.3005
R1452 VDD1.n39 VDD1.n38 9.3005
R1453 VDD1.n12 VDD1.n11 9.3005
R1454 VDD1.n33 VDD1.n32 9.3005
R1455 VDD1.n31 VDD1.n30 9.3005
R1456 VDD1.n16 VDD1.n15 9.3005
R1457 VDD1.n25 VDD1.n24 9.3005
R1458 VDD1.n23 VDD1.n22 9.3005
R1459 VDD1.n69 VDD1.n68 9.3005
R1460 VDD1.n108 VDD1.n107 9.3005
R1461 VDD1.n110 VDD1.n109 9.3005
R1462 VDD1.n65 VDD1.n64 9.3005
R1463 VDD1.n116 VDD1.n115 9.3005
R1464 VDD1.n118 VDD1.n117 9.3005
R1465 VDD1.n100 VDD1.n99 9.3005
R1466 VDD1.n73 VDD1.n72 9.3005
R1467 VDD1.n94 VDD1.n93 9.3005
R1468 VDD1.n92 VDD1.n91 9.3005
R1469 VDD1.n77 VDD1.n76 9.3005
R1470 VDD1.n86 VDD1.n85 9.3005
R1471 VDD1.n84 VDD1.n83 9.3005
R1472 VDD1.n102 VDD1.n101 9.3005
R1473 VDD1.n50 VDD1.n4 8.92171
R1474 VDD1.n37 VDD1.n12 8.92171
R1475 VDD1.n98 VDD1.n73 8.92171
R1476 VDD1.n111 VDD1.n65 8.92171
R1477 VDD1.n49 VDD1.n6 8.14595
R1478 VDD1.n38 VDD1.n10 8.14595
R1479 VDD1.n99 VDD1.n71 8.14595
R1480 VDD1.n110 VDD1.n67 8.14595
R1481 VDD1.n46 VDD1.n45 7.3702
R1482 VDD1.n42 VDD1.n41 7.3702
R1483 VDD1.n103 VDD1.n102 7.3702
R1484 VDD1.n107 VDD1.n106 7.3702
R1485 VDD1.n45 VDD1.n8 6.59444
R1486 VDD1.n42 VDD1.n8 6.59444
R1487 VDD1.n103 VDD1.n69 6.59444
R1488 VDD1.n106 VDD1.n69 6.59444
R1489 VDD1.n46 VDD1.n6 5.81868
R1490 VDD1.n41 VDD1.n10 5.81868
R1491 VDD1.n102 VDD1.n71 5.81868
R1492 VDD1.n107 VDD1.n67 5.81868
R1493 VDD1.n50 VDD1.n49 5.04292
R1494 VDD1.n38 VDD1.n37 5.04292
R1495 VDD1.n99 VDD1.n98 5.04292
R1496 VDD1.n111 VDD1.n110 5.04292
R1497 VDD1.n53 VDD1.n4 4.26717
R1498 VDD1.n34 VDD1.n12 4.26717
R1499 VDD1.n95 VDD1.n73 4.26717
R1500 VDD1.n114 VDD1.n65 4.26717
R1501 VDD1.n23 VDD1.n19 3.70982
R1502 VDD1.n84 VDD1.n80 3.70982
R1503 VDD1.n54 VDD1.n2 3.49141
R1504 VDD1.n33 VDD1.n14 3.49141
R1505 VDD1.n94 VDD1.n75 3.49141
R1506 VDD1.n115 VDD1.n63 3.49141
R1507 VDD1.n58 VDD1.n57 2.71565
R1508 VDD1.n30 VDD1.n29 2.71565
R1509 VDD1.n91 VDD1.n90 2.71565
R1510 VDD1.n119 VDD1.n118 2.71565
R1511 VDD1.n60 VDD1.n0 1.93989
R1512 VDD1.n26 VDD1.n16 1.93989
R1513 VDD1.n87 VDD1.n77 1.93989
R1514 VDD1.n121 VDD1.n61 1.93989
R1515 VDD1.n25 VDD1.n18 1.16414
R1516 VDD1.n86 VDD1.n79 1.16414
R1517 VDD1.n22 VDD1.n21 0.388379
R1518 VDD1.n83 VDD1.n82 0.388379
R1519 VDD1.n56 VDD1.n55 0.155672
R1520 VDD1.n55 VDD1.n3 0.155672
R1521 VDD1.n48 VDD1.n3 0.155672
R1522 VDD1.n48 VDD1.n47 0.155672
R1523 VDD1.n47 VDD1.n7 0.155672
R1524 VDD1.n40 VDD1.n7 0.155672
R1525 VDD1.n40 VDD1.n39 0.155672
R1526 VDD1.n39 VDD1.n11 0.155672
R1527 VDD1.n32 VDD1.n11 0.155672
R1528 VDD1.n32 VDD1.n31 0.155672
R1529 VDD1.n31 VDD1.n15 0.155672
R1530 VDD1.n24 VDD1.n15 0.155672
R1531 VDD1.n24 VDD1.n23 0.155672
R1532 VDD1.n85 VDD1.n84 0.155672
R1533 VDD1.n85 VDD1.n76 0.155672
R1534 VDD1.n92 VDD1.n76 0.155672
R1535 VDD1.n93 VDD1.n92 0.155672
R1536 VDD1.n93 VDD1.n72 0.155672
R1537 VDD1.n100 VDD1.n72 0.155672
R1538 VDD1.n101 VDD1.n100 0.155672
R1539 VDD1.n101 VDD1.n68 0.155672
R1540 VDD1.n108 VDD1.n68 0.155672
R1541 VDD1.n109 VDD1.n108 0.155672
R1542 VDD1.n109 VDD1.n64 0.155672
R1543 VDD1.n116 VDD1.n64 0.155672
R1544 VDD1.n117 VDD1.n116 0.155672
C0 w_n1762_n3218# VP 2.56825f
C1 w_n1762_n3218# VDD1 1.62189f
C2 VP VDD2 0.29318f
C3 B VTAIL 3.07819f
C4 VDD2 VDD1 0.56295f
C5 w_n1762_n3218# B 7.57192f
C6 VDD2 B 1.53543f
C7 VP VDD1 2.55169f
C8 VP B 1.24236f
C9 B VDD1 1.51375f
C10 VN VTAIL 2.04337f
C11 w_n1762_n3218# VN 2.34585f
C12 VDD2 VN 2.4092f
C13 w_n1762_n3218# VTAIL 2.67386f
C14 VDD2 VTAIL 4.86457f
C15 w_n1762_n3218# VDD2 1.63638f
C16 VP VN 4.8743f
C17 VN VDD1 0.147686f
C18 VP VTAIL 2.05775f
C19 VTAIL VDD1 4.82145f
C20 VN B 0.880537f
C21 VDD2 VSUBS 0.790625f
C22 VDD1 VSUBS 3.33414f
C23 VTAIL VSUBS 0.869419f
C24 VN VSUBS 7.53892f
C25 VP VSUBS 1.385371f
C26 B VSUBS 3.127038f
C27 w_n1762_n3218# VSUBS 69.8809f
C28 VDD1.n0 VSUBS 0.011499f
C29 VDD1.n1 VSUBS 0.025894f
C30 VDD1.n2 VSUBS 0.0116f
C31 VDD1.n3 VSUBS 0.020387f
C32 VDD1.n4 VSUBS 0.010955f
C33 VDD1.n5 VSUBS 0.025894f
C34 VDD1.n6 VSUBS 0.0116f
C35 VDD1.n7 VSUBS 0.020387f
C36 VDD1.n8 VSUBS 0.010955f
C37 VDD1.n9 VSUBS 0.025894f
C38 VDD1.n10 VSUBS 0.0116f
C39 VDD1.n11 VSUBS 0.020387f
C40 VDD1.n12 VSUBS 0.010955f
C41 VDD1.n13 VSUBS 0.025894f
C42 VDD1.n14 VSUBS 0.0116f
C43 VDD1.n15 VSUBS 0.020387f
C44 VDD1.n16 VSUBS 0.010955f
C45 VDD1.n17 VSUBS 0.025894f
C46 VDD1.n18 VSUBS 0.0116f
C47 VDD1.n19 VSUBS 0.121167f
C48 VDD1.t0 VSUBS 0.055249f
C49 VDD1.n20 VSUBS 0.019421f
C50 VDD1.n21 VSUBS 0.016473f
C51 VDD1.n22 VSUBS 0.010955f
C52 VDD1.n23 VSUBS 0.954681f
C53 VDD1.n24 VSUBS 0.020387f
C54 VDD1.n25 VSUBS 0.010955f
C55 VDD1.n26 VSUBS 0.0116f
C56 VDD1.n27 VSUBS 0.025894f
C57 VDD1.n28 VSUBS 0.025894f
C58 VDD1.n29 VSUBS 0.0116f
C59 VDD1.n30 VSUBS 0.010955f
C60 VDD1.n31 VSUBS 0.020387f
C61 VDD1.n32 VSUBS 0.020387f
C62 VDD1.n33 VSUBS 0.010955f
C63 VDD1.n34 VSUBS 0.0116f
C64 VDD1.n35 VSUBS 0.025894f
C65 VDD1.n36 VSUBS 0.025894f
C66 VDD1.n37 VSUBS 0.0116f
C67 VDD1.n38 VSUBS 0.010955f
C68 VDD1.n39 VSUBS 0.020387f
C69 VDD1.n40 VSUBS 0.020387f
C70 VDD1.n41 VSUBS 0.010955f
C71 VDD1.n42 VSUBS 0.0116f
C72 VDD1.n43 VSUBS 0.025894f
C73 VDD1.n44 VSUBS 0.025894f
C74 VDD1.n45 VSUBS 0.0116f
C75 VDD1.n46 VSUBS 0.010955f
C76 VDD1.n47 VSUBS 0.020387f
C77 VDD1.n48 VSUBS 0.020387f
C78 VDD1.n49 VSUBS 0.010955f
C79 VDD1.n50 VSUBS 0.0116f
C80 VDD1.n51 VSUBS 0.025894f
C81 VDD1.n52 VSUBS 0.025894f
C82 VDD1.n53 VSUBS 0.0116f
C83 VDD1.n54 VSUBS 0.010955f
C84 VDD1.n55 VSUBS 0.020387f
C85 VDD1.n56 VSUBS 0.052973f
C86 VDD1.n57 VSUBS 0.010955f
C87 VDD1.n58 VSUBS 0.0116f
C88 VDD1.n59 VSUBS 0.056803f
C89 VDD1.n60 VSUBS 0.053325f
C90 VDD1.n61 VSUBS 0.011499f
C91 VDD1.n62 VSUBS 0.025894f
C92 VDD1.n63 VSUBS 0.0116f
C93 VDD1.n64 VSUBS 0.020387f
C94 VDD1.n65 VSUBS 0.010955f
C95 VDD1.n66 VSUBS 0.025894f
C96 VDD1.n67 VSUBS 0.0116f
C97 VDD1.n68 VSUBS 0.020387f
C98 VDD1.n69 VSUBS 0.010955f
C99 VDD1.n70 VSUBS 0.025894f
C100 VDD1.n71 VSUBS 0.0116f
C101 VDD1.n72 VSUBS 0.020387f
C102 VDD1.n73 VSUBS 0.010955f
C103 VDD1.n74 VSUBS 0.025894f
C104 VDD1.n75 VSUBS 0.0116f
C105 VDD1.n76 VSUBS 0.020387f
C106 VDD1.n77 VSUBS 0.010955f
C107 VDD1.n78 VSUBS 0.025894f
C108 VDD1.n79 VSUBS 0.0116f
C109 VDD1.n80 VSUBS 0.121167f
C110 VDD1.t1 VSUBS 0.055249f
C111 VDD1.n81 VSUBS 0.019421f
C112 VDD1.n82 VSUBS 0.016473f
C113 VDD1.n83 VSUBS 0.010955f
C114 VDD1.n84 VSUBS 0.954681f
C115 VDD1.n85 VSUBS 0.020387f
C116 VDD1.n86 VSUBS 0.010955f
C117 VDD1.n87 VSUBS 0.0116f
C118 VDD1.n88 VSUBS 0.025894f
C119 VDD1.n89 VSUBS 0.025894f
C120 VDD1.n90 VSUBS 0.0116f
C121 VDD1.n91 VSUBS 0.010955f
C122 VDD1.n92 VSUBS 0.020387f
C123 VDD1.n93 VSUBS 0.020387f
C124 VDD1.n94 VSUBS 0.010955f
C125 VDD1.n95 VSUBS 0.0116f
C126 VDD1.n96 VSUBS 0.025894f
C127 VDD1.n97 VSUBS 0.025894f
C128 VDD1.n98 VSUBS 0.0116f
C129 VDD1.n99 VSUBS 0.010955f
C130 VDD1.n100 VSUBS 0.020387f
C131 VDD1.n101 VSUBS 0.020387f
C132 VDD1.n102 VSUBS 0.010955f
C133 VDD1.n103 VSUBS 0.0116f
C134 VDD1.n104 VSUBS 0.025894f
C135 VDD1.n105 VSUBS 0.025894f
C136 VDD1.n106 VSUBS 0.0116f
C137 VDD1.n107 VSUBS 0.010955f
C138 VDD1.n108 VSUBS 0.020387f
C139 VDD1.n109 VSUBS 0.020387f
C140 VDD1.n110 VSUBS 0.010955f
C141 VDD1.n111 VSUBS 0.0116f
C142 VDD1.n112 VSUBS 0.025894f
C143 VDD1.n113 VSUBS 0.025894f
C144 VDD1.n114 VSUBS 0.0116f
C145 VDD1.n115 VSUBS 0.010955f
C146 VDD1.n116 VSUBS 0.020387f
C147 VDD1.n117 VSUBS 0.052973f
C148 VDD1.n118 VSUBS 0.010955f
C149 VDD1.n119 VSUBS 0.0116f
C150 VDD1.n120 VSUBS 0.056803f
C151 VDD1.n121 VSUBS 0.556844f
C152 VP.t1 VSUBS 3.45042f
C153 VP.t0 VSUBS 2.96112f
C154 VP.n0 VSUBS 5.71506f
C155 VDD2.n0 VSUBS 0.01146f
C156 VDD2.n1 VSUBS 0.025807f
C157 VDD2.n2 VSUBS 0.01156f
C158 VDD2.n3 VSUBS 0.020318f
C159 VDD2.n4 VSUBS 0.010918f
C160 VDD2.n5 VSUBS 0.025807f
C161 VDD2.n6 VSUBS 0.01156f
C162 VDD2.n7 VSUBS 0.020318f
C163 VDD2.n8 VSUBS 0.010918f
C164 VDD2.n9 VSUBS 0.025807f
C165 VDD2.n10 VSUBS 0.01156f
C166 VDD2.n11 VSUBS 0.020318f
C167 VDD2.n12 VSUBS 0.010918f
C168 VDD2.n13 VSUBS 0.025807f
C169 VDD2.n14 VSUBS 0.01156f
C170 VDD2.n15 VSUBS 0.020318f
C171 VDD2.n16 VSUBS 0.010918f
C172 VDD2.n17 VSUBS 0.025807f
C173 VDD2.n18 VSUBS 0.01156f
C174 VDD2.n19 VSUBS 0.120759f
C175 VDD2.t0 VSUBS 0.055063f
C176 VDD2.n20 VSUBS 0.019355f
C177 VDD2.n21 VSUBS 0.016417f
C178 VDD2.n22 VSUBS 0.010918f
C179 VDD2.n23 VSUBS 0.951461f
C180 VDD2.n24 VSUBS 0.020318f
C181 VDD2.n25 VSUBS 0.010918f
C182 VDD2.n26 VSUBS 0.01156f
C183 VDD2.n27 VSUBS 0.025807f
C184 VDD2.n28 VSUBS 0.025807f
C185 VDD2.n29 VSUBS 0.01156f
C186 VDD2.n30 VSUBS 0.010918f
C187 VDD2.n31 VSUBS 0.020318f
C188 VDD2.n32 VSUBS 0.020318f
C189 VDD2.n33 VSUBS 0.010918f
C190 VDD2.n34 VSUBS 0.01156f
C191 VDD2.n35 VSUBS 0.025807f
C192 VDD2.n36 VSUBS 0.025807f
C193 VDD2.n37 VSUBS 0.01156f
C194 VDD2.n38 VSUBS 0.010918f
C195 VDD2.n39 VSUBS 0.020318f
C196 VDD2.n40 VSUBS 0.020318f
C197 VDD2.n41 VSUBS 0.010918f
C198 VDD2.n42 VSUBS 0.01156f
C199 VDD2.n43 VSUBS 0.025807f
C200 VDD2.n44 VSUBS 0.025807f
C201 VDD2.n45 VSUBS 0.01156f
C202 VDD2.n46 VSUBS 0.010918f
C203 VDD2.n47 VSUBS 0.020318f
C204 VDD2.n48 VSUBS 0.020318f
C205 VDD2.n49 VSUBS 0.010918f
C206 VDD2.n50 VSUBS 0.01156f
C207 VDD2.n51 VSUBS 0.025807f
C208 VDD2.n52 VSUBS 0.025807f
C209 VDD2.n53 VSUBS 0.01156f
C210 VDD2.n54 VSUBS 0.010918f
C211 VDD2.n55 VSUBS 0.020318f
C212 VDD2.n56 VSUBS 0.052794f
C213 VDD2.n57 VSUBS 0.010918f
C214 VDD2.n58 VSUBS 0.01156f
C215 VDD2.n59 VSUBS 0.056612f
C216 VDD2.n60 VSUBS 0.522793f
C217 VDD2.n61 VSUBS 0.01146f
C218 VDD2.n62 VSUBS 0.025807f
C219 VDD2.n63 VSUBS 0.01156f
C220 VDD2.n64 VSUBS 0.020318f
C221 VDD2.n65 VSUBS 0.010918f
C222 VDD2.n66 VSUBS 0.025807f
C223 VDD2.n67 VSUBS 0.01156f
C224 VDD2.n68 VSUBS 0.020318f
C225 VDD2.n69 VSUBS 0.010918f
C226 VDD2.n70 VSUBS 0.025807f
C227 VDD2.n71 VSUBS 0.01156f
C228 VDD2.n72 VSUBS 0.020318f
C229 VDD2.n73 VSUBS 0.010918f
C230 VDD2.n74 VSUBS 0.025807f
C231 VDD2.n75 VSUBS 0.01156f
C232 VDD2.n76 VSUBS 0.020318f
C233 VDD2.n77 VSUBS 0.010918f
C234 VDD2.n78 VSUBS 0.025807f
C235 VDD2.n79 VSUBS 0.01156f
C236 VDD2.n80 VSUBS 0.120759f
C237 VDD2.t1 VSUBS 0.055063f
C238 VDD2.n81 VSUBS 0.019355f
C239 VDD2.n82 VSUBS 0.016417f
C240 VDD2.n83 VSUBS 0.010918f
C241 VDD2.n84 VSUBS 0.951461f
C242 VDD2.n85 VSUBS 0.020318f
C243 VDD2.n86 VSUBS 0.010918f
C244 VDD2.n87 VSUBS 0.01156f
C245 VDD2.n88 VSUBS 0.025807f
C246 VDD2.n89 VSUBS 0.025807f
C247 VDD2.n90 VSUBS 0.01156f
C248 VDD2.n91 VSUBS 0.010918f
C249 VDD2.n92 VSUBS 0.020318f
C250 VDD2.n93 VSUBS 0.020318f
C251 VDD2.n94 VSUBS 0.010918f
C252 VDD2.n95 VSUBS 0.01156f
C253 VDD2.n96 VSUBS 0.025807f
C254 VDD2.n97 VSUBS 0.025807f
C255 VDD2.n98 VSUBS 0.01156f
C256 VDD2.n99 VSUBS 0.010918f
C257 VDD2.n100 VSUBS 0.020318f
C258 VDD2.n101 VSUBS 0.020318f
C259 VDD2.n102 VSUBS 0.010918f
C260 VDD2.n103 VSUBS 0.01156f
C261 VDD2.n104 VSUBS 0.025807f
C262 VDD2.n105 VSUBS 0.025807f
C263 VDD2.n106 VSUBS 0.01156f
C264 VDD2.n107 VSUBS 0.010918f
C265 VDD2.n108 VSUBS 0.020318f
C266 VDD2.n109 VSUBS 0.020318f
C267 VDD2.n110 VSUBS 0.010918f
C268 VDD2.n111 VSUBS 0.01156f
C269 VDD2.n112 VSUBS 0.025807f
C270 VDD2.n113 VSUBS 0.025807f
C271 VDD2.n114 VSUBS 0.01156f
C272 VDD2.n115 VSUBS 0.010918f
C273 VDD2.n116 VSUBS 0.020318f
C274 VDD2.n117 VSUBS 0.052794f
C275 VDD2.n118 VSUBS 0.010918f
C276 VDD2.n119 VSUBS 0.01156f
C277 VDD2.n120 VSUBS 0.056612f
C278 VDD2.n121 VSUBS 0.052461f
C279 VDD2.n122 VSUBS 2.28069f
C280 VTAIL.n0 VSUBS 0.016513f
C281 VTAIL.n1 VSUBS 0.037185f
C282 VTAIL.n2 VSUBS 0.016657f
C283 VTAIL.n3 VSUBS 0.029277f
C284 VTAIL.n4 VSUBS 0.015732f
C285 VTAIL.n5 VSUBS 0.037185f
C286 VTAIL.n6 VSUBS 0.016657f
C287 VTAIL.n7 VSUBS 0.029277f
C288 VTAIL.n8 VSUBS 0.015732f
C289 VTAIL.n9 VSUBS 0.037185f
C290 VTAIL.n10 VSUBS 0.016657f
C291 VTAIL.n11 VSUBS 0.029277f
C292 VTAIL.n12 VSUBS 0.015732f
C293 VTAIL.n13 VSUBS 0.037185f
C294 VTAIL.n14 VSUBS 0.016657f
C295 VTAIL.n15 VSUBS 0.029277f
C296 VTAIL.n16 VSUBS 0.015732f
C297 VTAIL.n17 VSUBS 0.037185f
C298 VTAIL.n18 VSUBS 0.016657f
C299 VTAIL.n19 VSUBS 0.174f
C300 VTAIL.t0 VSUBS 0.07934f
C301 VTAIL.n20 VSUBS 0.027889f
C302 VTAIL.n21 VSUBS 0.023655f
C303 VTAIL.n22 VSUBS 0.015732f
C304 VTAIL.n23 VSUBS 1.37095f
C305 VTAIL.n24 VSUBS 0.029277f
C306 VTAIL.n25 VSUBS 0.015732f
C307 VTAIL.n26 VSUBS 0.016657f
C308 VTAIL.n27 VSUBS 0.037185f
C309 VTAIL.n28 VSUBS 0.037185f
C310 VTAIL.n29 VSUBS 0.016657f
C311 VTAIL.n30 VSUBS 0.015732f
C312 VTAIL.n31 VSUBS 0.029277f
C313 VTAIL.n32 VSUBS 0.029277f
C314 VTAIL.n33 VSUBS 0.015732f
C315 VTAIL.n34 VSUBS 0.016657f
C316 VTAIL.n35 VSUBS 0.037185f
C317 VTAIL.n36 VSUBS 0.037185f
C318 VTAIL.n37 VSUBS 0.016657f
C319 VTAIL.n38 VSUBS 0.015732f
C320 VTAIL.n39 VSUBS 0.029277f
C321 VTAIL.n40 VSUBS 0.029277f
C322 VTAIL.n41 VSUBS 0.015732f
C323 VTAIL.n42 VSUBS 0.016657f
C324 VTAIL.n43 VSUBS 0.037185f
C325 VTAIL.n44 VSUBS 0.037185f
C326 VTAIL.n45 VSUBS 0.016657f
C327 VTAIL.n46 VSUBS 0.015732f
C328 VTAIL.n47 VSUBS 0.029277f
C329 VTAIL.n48 VSUBS 0.029277f
C330 VTAIL.n49 VSUBS 0.015732f
C331 VTAIL.n50 VSUBS 0.016657f
C332 VTAIL.n51 VSUBS 0.037185f
C333 VTAIL.n52 VSUBS 0.037185f
C334 VTAIL.n53 VSUBS 0.016657f
C335 VTAIL.n54 VSUBS 0.015732f
C336 VTAIL.n55 VSUBS 0.029277f
C337 VTAIL.n56 VSUBS 0.07607f
C338 VTAIL.n57 VSUBS 0.015732f
C339 VTAIL.n58 VSUBS 0.016657f
C340 VTAIL.n59 VSUBS 0.081571f
C341 VTAIL.n60 VSUBS 0.055408f
C342 VTAIL.n61 VSUBS 1.75218f
C343 VTAIL.n62 VSUBS 0.016513f
C344 VTAIL.n63 VSUBS 0.037185f
C345 VTAIL.n64 VSUBS 0.016657f
C346 VTAIL.n65 VSUBS 0.029277f
C347 VTAIL.n66 VSUBS 0.015732f
C348 VTAIL.n67 VSUBS 0.037185f
C349 VTAIL.n68 VSUBS 0.016657f
C350 VTAIL.n69 VSUBS 0.029277f
C351 VTAIL.n70 VSUBS 0.015732f
C352 VTAIL.n71 VSUBS 0.037185f
C353 VTAIL.n72 VSUBS 0.016657f
C354 VTAIL.n73 VSUBS 0.029277f
C355 VTAIL.n74 VSUBS 0.015732f
C356 VTAIL.n75 VSUBS 0.037185f
C357 VTAIL.n76 VSUBS 0.016657f
C358 VTAIL.n77 VSUBS 0.029277f
C359 VTAIL.n78 VSUBS 0.015732f
C360 VTAIL.n79 VSUBS 0.037185f
C361 VTAIL.n80 VSUBS 0.016657f
C362 VTAIL.n81 VSUBS 0.174f
C363 VTAIL.t3 VSUBS 0.07934f
C364 VTAIL.n82 VSUBS 0.027889f
C365 VTAIL.n83 VSUBS 0.023655f
C366 VTAIL.n84 VSUBS 0.015732f
C367 VTAIL.n85 VSUBS 1.37095f
C368 VTAIL.n86 VSUBS 0.029277f
C369 VTAIL.n87 VSUBS 0.015732f
C370 VTAIL.n88 VSUBS 0.016657f
C371 VTAIL.n89 VSUBS 0.037185f
C372 VTAIL.n90 VSUBS 0.037185f
C373 VTAIL.n91 VSUBS 0.016657f
C374 VTAIL.n92 VSUBS 0.015732f
C375 VTAIL.n93 VSUBS 0.029277f
C376 VTAIL.n94 VSUBS 0.029277f
C377 VTAIL.n95 VSUBS 0.015732f
C378 VTAIL.n96 VSUBS 0.016657f
C379 VTAIL.n97 VSUBS 0.037185f
C380 VTAIL.n98 VSUBS 0.037185f
C381 VTAIL.n99 VSUBS 0.016657f
C382 VTAIL.n100 VSUBS 0.015732f
C383 VTAIL.n101 VSUBS 0.029277f
C384 VTAIL.n102 VSUBS 0.029277f
C385 VTAIL.n103 VSUBS 0.015732f
C386 VTAIL.n104 VSUBS 0.016657f
C387 VTAIL.n105 VSUBS 0.037185f
C388 VTAIL.n106 VSUBS 0.037185f
C389 VTAIL.n107 VSUBS 0.016657f
C390 VTAIL.n108 VSUBS 0.015732f
C391 VTAIL.n109 VSUBS 0.029277f
C392 VTAIL.n110 VSUBS 0.029277f
C393 VTAIL.n111 VSUBS 0.015732f
C394 VTAIL.n112 VSUBS 0.016657f
C395 VTAIL.n113 VSUBS 0.037185f
C396 VTAIL.n114 VSUBS 0.037185f
C397 VTAIL.n115 VSUBS 0.016657f
C398 VTAIL.n116 VSUBS 0.015732f
C399 VTAIL.n117 VSUBS 0.029277f
C400 VTAIL.n118 VSUBS 0.07607f
C401 VTAIL.n119 VSUBS 0.015732f
C402 VTAIL.n120 VSUBS 0.016657f
C403 VTAIL.n121 VSUBS 0.081571f
C404 VTAIL.n122 VSUBS 0.055408f
C405 VTAIL.n123 VSUBS 1.78695f
C406 VTAIL.n124 VSUBS 0.016513f
C407 VTAIL.n125 VSUBS 0.037185f
C408 VTAIL.n126 VSUBS 0.016657f
C409 VTAIL.n127 VSUBS 0.029277f
C410 VTAIL.n128 VSUBS 0.015732f
C411 VTAIL.n129 VSUBS 0.037185f
C412 VTAIL.n130 VSUBS 0.016657f
C413 VTAIL.n131 VSUBS 0.029277f
C414 VTAIL.n132 VSUBS 0.015732f
C415 VTAIL.n133 VSUBS 0.037185f
C416 VTAIL.n134 VSUBS 0.016657f
C417 VTAIL.n135 VSUBS 0.029277f
C418 VTAIL.n136 VSUBS 0.015732f
C419 VTAIL.n137 VSUBS 0.037185f
C420 VTAIL.n138 VSUBS 0.016657f
C421 VTAIL.n139 VSUBS 0.029277f
C422 VTAIL.n140 VSUBS 0.015732f
C423 VTAIL.n141 VSUBS 0.037185f
C424 VTAIL.n142 VSUBS 0.016657f
C425 VTAIL.n143 VSUBS 0.174f
C426 VTAIL.t1 VSUBS 0.07934f
C427 VTAIL.n144 VSUBS 0.027889f
C428 VTAIL.n145 VSUBS 0.023655f
C429 VTAIL.n146 VSUBS 0.015732f
C430 VTAIL.n147 VSUBS 1.37095f
C431 VTAIL.n148 VSUBS 0.029277f
C432 VTAIL.n149 VSUBS 0.015732f
C433 VTAIL.n150 VSUBS 0.016657f
C434 VTAIL.n151 VSUBS 0.037185f
C435 VTAIL.n152 VSUBS 0.037185f
C436 VTAIL.n153 VSUBS 0.016657f
C437 VTAIL.n154 VSUBS 0.015732f
C438 VTAIL.n155 VSUBS 0.029277f
C439 VTAIL.n156 VSUBS 0.029277f
C440 VTAIL.n157 VSUBS 0.015732f
C441 VTAIL.n158 VSUBS 0.016657f
C442 VTAIL.n159 VSUBS 0.037185f
C443 VTAIL.n160 VSUBS 0.037185f
C444 VTAIL.n161 VSUBS 0.016657f
C445 VTAIL.n162 VSUBS 0.015732f
C446 VTAIL.n163 VSUBS 0.029277f
C447 VTAIL.n164 VSUBS 0.029277f
C448 VTAIL.n165 VSUBS 0.015732f
C449 VTAIL.n166 VSUBS 0.016657f
C450 VTAIL.n167 VSUBS 0.037185f
C451 VTAIL.n168 VSUBS 0.037185f
C452 VTAIL.n169 VSUBS 0.016657f
C453 VTAIL.n170 VSUBS 0.015732f
C454 VTAIL.n171 VSUBS 0.029277f
C455 VTAIL.n172 VSUBS 0.029277f
C456 VTAIL.n173 VSUBS 0.015732f
C457 VTAIL.n174 VSUBS 0.016657f
C458 VTAIL.n175 VSUBS 0.037185f
C459 VTAIL.n176 VSUBS 0.037185f
C460 VTAIL.n177 VSUBS 0.016657f
C461 VTAIL.n178 VSUBS 0.015732f
C462 VTAIL.n179 VSUBS 0.029277f
C463 VTAIL.n180 VSUBS 0.07607f
C464 VTAIL.n181 VSUBS 0.015732f
C465 VTAIL.n182 VSUBS 0.016657f
C466 VTAIL.n183 VSUBS 0.081571f
C467 VTAIL.n184 VSUBS 0.055408f
C468 VTAIL.n185 VSUBS 1.62593f
C469 VTAIL.n186 VSUBS 0.016513f
C470 VTAIL.n187 VSUBS 0.037185f
C471 VTAIL.n188 VSUBS 0.016657f
C472 VTAIL.n189 VSUBS 0.029277f
C473 VTAIL.n190 VSUBS 0.015732f
C474 VTAIL.n191 VSUBS 0.037185f
C475 VTAIL.n192 VSUBS 0.016657f
C476 VTAIL.n193 VSUBS 0.029277f
C477 VTAIL.n194 VSUBS 0.015732f
C478 VTAIL.n195 VSUBS 0.037185f
C479 VTAIL.n196 VSUBS 0.016657f
C480 VTAIL.n197 VSUBS 0.029277f
C481 VTAIL.n198 VSUBS 0.015732f
C482 VTAIL.n199 VSUBS 0.037185f
C483 VTAIL.n200 VSUBS 0.016657f
C484 VTAIL.n201 VSUBS 0.029277f
C485 VTAIL.n202 VSUBS 0.015732f
C486 VTAIL.n203 VSUBS 0.037185f
C487 VTAIL.n204 VSUBS 0.016657f
C488 VTAIL.n205 VSUBS 0.174f
C489 VTAIL.t2 VSUBS 0.07934f
C490 VTAIL.n206 VSUBS 0.027889f
C491 VTAIL.n207 VSUBS 0.023655f
C492 VTAIL.n208 VSUBS 0.015732f
C493 VTAIL.n209 VSUBS 1.37095f
C494 VTAIL.n210 VSUBS 0.029277f
C495 VTAIL.n211 VSUBS 0.015732f
C496 VTAIL.n212 VSUBS 0.016657f
C497 VTAIL.n213 VSUBS 0.037185f
C498 VTAIL.n214 VSUBS 0.037185f
C499 VTAIL.n215 VSUBS 0.016657f
C500 VTAIL.n216 VSUBS 0.015732f
C501 VTAIL.n217 VSUBS 0.029277f
C502 VTAIL.n218 VSUBS 0.029277f
C503 VTAIL.n219 VSUBS 0.015732f
C504 VTAIL.n220 VSUBS 0.016657f
C505 VTAIL.n221 VSUBS 0.037185f
C506 VTAIL.n222 VSUBS 0.037185f
C507 VTAIL.n223 VSUBS 0.016657f
C508 VTAIL.n224 VSUBS 0.015732f
C509 VTAIL.n225 VSUBS 0.029277f
C510 VTAIL.n226 VSUBS 0.029277f
C511 VTAIL.n227 VSUBS 0.015732f
C512 VTAIL.n228 VSUBS 0.016657f
C513 VTAIL.n229 VSUBS 0.037185f
C514 VTAIL.n230 VSUBS 0.037185f
C515 VTAIL.n231 VSUBS 0.016657f
C516 VTAIL.n232 VSUBS 0.015732f
C517 VTAIL.n233 VSUBS 0.029277f
C518 VTAIL.n234 VSUBS 0.029277f
C519 VTAIL.n235 VSUBS 0.015732f
C520 VTAIL.n236 VSUBS 0.016657f
C521 VTAIL.n237 VSUBS 0.037185f
C522 VTAIL.n238 VSUBS 0.037185f
C523 VTAIL.n239 VSUBS 0.016657f
C524 VTAIL.n240 VSUBS 0.015732f
C525 VTAIL.n241 VSUBS 0.029277f
C526 VTAIL.n242 VSUBS 0.07607f
C527 VTAIL.n243 VSUBS 0.015732f
C528 VTAIL.n244 VSUBS 0.016657f
C529 VTAIL.n245 VSUBS 0.081571f
C530 VTAIL.n246 VSUBS 0.055408f
C531 VTAIL.n247 VSUBS 1.53586f
C532 VN.t1 VSUBS 2.79963f
C533 VN.t0 VSUBS 3.26646f
C534 B.n0 VSUBS 0.005979f
C535 B.n1 VSUBS 0.005979f
C536 B.n2 VSUBS 0.008843f
C537 B.n3 VSUBS 0.006777f
C538 B.n4 VSUBS 0.006777f
C539 B.n5 VSUBS 0.006777f
C540 B.n6 VSUBS 0.006777f
C541 B.n7 VSUBS 0.006777f
C542 B.n8 VSUBS 0.006777f
C543 B.n9 VSUBS 0.006777f
C544 B.n10 VSUBS 0.006777f
C545 B.n11 VSUBS 0.016973f
C546 B.n12 VSUBS 0.006777f
C547 B.n13 VSUBS 0.006777f
C548 B.n14 VSUBS 0.006777f
C549 B.n15 VSUBS 0.006777f
C550 B.n16 VSUBS 0.006777f
C551 B.n17 VSUBS 0.006777f
C552 B.n18 VSUBS 0.006777f
C553 B.n19 VSUBS 0.006777f
C554 B.n20 VSUBS 0.006777f
C555 B.n21 VSUBS 0.006777f
C556 B.n22 VSUBS 0.006777f
C557 B.n23 VSUBS 0.006777f
C558 B.n24 VSUBS 0.006777f
C559 B.n25 VSUBS 0.006777f
C560 B.n26 VSUBS 0.006777f
C561 B.n27 VSUBS 0.006777f
C562 B.n28 VSUBS 0.006777f
C563 B.n29 VSUBS 0.006777f
C564 B.n30 VSUBS 0.006777f
C565 B.n31 VSUBS 0.006777f
C566 B.t10 VSUBS 0.188043f
C567 B.t11 VSUBS 0.209177f
C568 B.t9 VSUBS 0.795368f
C569 B.n32 VSUBS 0.327392f
C570 B.n33 VSUBS 0.229992f
C571 B.n34 VSUBS 0.006777f
C572 B.n35 VSUBS 0.006777f
C573 B.n36 VSUBS 0.006777f
C574 B.n37 VSUBS 0.006777f
C575 B.t4 VSUBS 0.188045f
C576 B.t5 VSUBS 0.209179f
C577 B.t3 VSUBS 0.795368f
C578 B.n38 VSUBS 0.327389f
C579 B.n39 VSUBS 0.229989f
C580 B.n40 VSUBS 0.015701f
C581 B.n41 VSUBS 0.006777f
C582 B.n42 VSUBS 0.006777f
C583 B.n43 VSUBS 0.006777f
C584 B.n44 VSUBS 0.006777f
C585 B.n45 VSUBS 0.006777f
C586 B.n46 VSUBS 0.006777f
C587 B.n47 VSUBS 0.006777f
C588 B.n48 VSUBS 0.006777f
C589 B.n49 VSUBS 0.006777f
C590 B.n50 VSUBS 0.006777f
C591 B.n51 VSUBS 0.006777f
C592 B.n52 VSUBS 0.006777f
C593 B.n53 VSUBS 0.006777f
C594 B.n54 VSUBS 0.006777f
C595 B.n55 VSUBS 0.006777f
C596 B.n56 VSUBS 0.006777f
C597 B.n57 VSUBS 0.006777f
C598 B.n58 VSUBS 0.006777f
C599 B.n59 VSUBS 0.006777f
C600 B.n60 VSUBS 0.016973f
C601 B.n61 VSUBS 0.006777f
C602 B.n62 VSUBS 0.006777f
C603 B.n63 VSUBS 0.006777f
C604 B.n64 VSUBS 0.006777f
C605 B.n65 VSUBS 0.006777f
C606 B.n66 VSUBS 0.006777f
C607 B.n67 VSUBS 0.006777f
C608 B.n68 VSUBS 0.006777f
C609 B.n69 VSUBS 0.006777f
C610 B.n70 VSUBS 0.006777f
C611 B.n71 VSUBS 0.006777f
C612 B.n72 VSUBS 0.006777f
C613 B.n73 VSUBS 0.006777f
C614 B.n74 VSUBS 0.006777f
C615 B.n75 VSUBS 0.006777f
C616 B.n76 VSUBS 0.006777f
C617 B.n77 VSUBS 0.006777f
C618 B.n78 VSUBS 0.006777f
C619 B.n79 VSUBS 0.006777f
C620 B.n80 VSUBS 0.017007f
C621 B.n81 VSUBS 0.006777f
C622 B.n82 VSUBS 0.006777f
C623 B.n83 VSUBS 0.006777f
C624 B.n84 VSUBS 0.006777f
C625 B.n85 VSUBS 0.006777f
C626 B.n86 VSUBS 0.006777f
C627 B.n87 VSUBS 0.006777f
C628 B.n88 VSUBS 0.006777f
C629 B.n89 VSUBS 0.006777f
C630 B.n90 VSUBS 0.006777f
C631 B.n91 VSUBS 0.006777f
C632 B.n92 VSUBS 0.006777f
C633 B.n93 VSUBS 0.006777f
C634 B.n94 VSUBS 0.006777f
C635 B.n95 VSUBS 0.006777f
C636 B.n96 VSUBS 0.006777f
C637 B.n97 VSUBS 0.006777f
C638 B.n98 VSUBS 0.006777f
C639 B.n99 VSUBS 0.006777f
C640 B.t2 VSUBS 0.188045f
C641 B.t1 VSUBS 0.209179f
C642 B.t0 VSUBS 0.795368f
C643 B.n100 VSUBS 0.327389f
C644 B.n101 VSUBS 0.229989f
C645 B.n102 VSUBS 0.006777f
C646 B.n103 VSUBS 0.006777f
C647 B.n104 VSUBS 0.006777f
C648 B.n105 VSUBS 0.006777f
C649 B.n106 VSUBS 0.003787f
C650 B.n107 VSUBS 0.006777f
C651 B.n108 VSUBS 0.006777f
C652 B.n109 VSUBS 0.006777f
C653 B.n110 VSUBS 0.006777f
C654 B.n111 VSUBS 0.006777f
C655 B.n112 VSUBS 0.006777f
C656 B.n113 VSUBS 0.006777f
C657 B.n114 VSUBS 0.006777f
C658 B.n115 VSUBS 0.006777f
C659 B.n116 VSUBS 0.006777f
C660 B.n117 VSUBS 0.006777f
C661 B.n118 VSUBS 0.006777f
C662 B.n119 VSUBS 0.006777f
C663 B.n120 VSUBS 0.006777f
C664 B.n121 VSUBS 0.006777f
C665 B.n122 VSUBS 0.006777f
C666 B.n123 VSUBS 0.006777f
C667 B.n124 VSUBS 0.006777f
C668 B.n125 VSUBS 0.006777f
C669 B.n126 VSUBS 0.016973f
C670 B.n127 VSUBS 0.006777f
C671 B.n128 VSUBS 0.006777f
C672 B.n129 VSUBS 0.006777f
C673 B.n130 VSUBS 0.006777f
C674 B.n131 VSUBS 0.006777f
C675 B.n132 VSUBS 0.006777f
C676 B.n133 VSUBS 0.006777f
C677 B.n134 VSUBS 0.006777f
C678 B.n135 VSUBS 0.006777f
C679 B.n136 VSUBS 0.006777f
C680 B.n137 VSUBS 0.006777f
C681 B.n138 VSUBS 0.006777f
C682 B.n139 VSUBS 0.006777f
C683 B.n140 VSUBS 0.006777f
C684 B.n141 VSUBS 0.006777f
C685 B.n142 VSUBS 0.006777f
C686 B.n143 VSUBS 0.006777f
C687 B.n144 VSUBS 0.006777f
C688 B.n145 VSUBS 0.006777f
C689 B.n146 VSUBS 0.006777f
C690 B.n147 VSUBS 0.006777f
C691 B.n148 VSUBS 0.006777f
C692 B.n149 VSUBS 0.006777f
C693 B.n150 VSUBS 0.006777f
C694 B.n151 VSUBS 0.006777f
C695 B.n152 VSUBS 0.006777f
C696 B.n153 VSUBS 0.006777f
C697 B.n154 VSUBS 0.006777f
C698 B.n155 VSUBS 0.006777f
C699 B.n156 VSUBS 0.006777f
C700 B.n157 VSUBS 0.006777f
C701 B.n158 VSUBS 0.006777f
C702 B.n159 VSUBS 0.006777f
C703 B.n160 VSUBS 0.006777f
C704 B.n161 VSUBS 0.016973f
C705 B.n162 VSUBS 0.017708f
C706 B.n163 VSUBS 0.017708f
C707 B.n164 VSUBS 0.006777f
C708 B.n165 VSUBS 0.006777f
C709 B.n166 VSUBS 0.006777f
C710 B.n167 VSUBS 0.006777f
C711 B.n168 VSUBS 0.006777f
C712 B.n169 VSUBS 0.006777f
C713 B.n170 VSUBS 0.006777f
C714 B.n171 VSUBS 0.006777f
C715 B.n172 VSUBS 0.006777f
C716 B.n173 VSUBS 0.006777f
C717 B.n174 VSUBS 0.006777f
C718 B.n175 VSUBS 0.006777f
C719 B.n176 VSUBS 0.006777f
C720 B.n177 VSUBS 0.006777f
C721 B.n178 VSUBS 0.006777f
C722 B.n179 VSUBS 0.006777f
C723 B.n180 VSUBS 0.006777f
C724 B.n181 VSUBS 0.006777f
C725 B.n182 VSUBS 0.006777f
C726 B.n183 VSUBS 0.006777f
C727 B.n184 VSUBS 0.006777f
C728 B.n185 VSUBS 0.006777f
C729 B.n186 VSUBS 0.006777f
C730 B.n187 VSUBS 0.006777f
C731 B.n188 VSUBS 0.006777f
C732 B.n189 VSUBS 0.006777f
C733 B.n190 VSUBS 0.006777f
C734 B.n191 VSUBS 0.006777f
C735 B.n192 VSUBS 0.006777f
C736 B.n193 VSUBS 0.006777f
C737 B.n194 VSUBS 0.006777f
C738 B.n195 VSUBS 0.006777f
C739 B.n196 VSUBS 0.006777f
C740 B.n197 VSUBS 0.006777f
C741 B.n198 VSUBS 0.006777f
C742 B.n199 VSUBS 0.006777f
C743 B.n200 VSUBS 0.006777f
C744 B.n201 VSUBS 0.006777f
C745 B.n202 VSUBS 0.006777f
C746 B.n203 VSUBS 0.006777f
C747 B.n204 VSUBS 0.006777f
C748 B.n205 VSUBS 0.006777f
C749 B.n206 VSUBS 0.006777f
C750 B.n207 VSUBS 0.006777f
C751 B.n208 VSUBS 0.006777f
C752 B.n209 VSUBS 0.006777f
C753 B.n210 VSUBS 0.006777f
C754 B.n211 VSUBS 0.006777f
C755 B.n212 VSUBS 0.006777f
C756 B.n213 VSUBS 0.006777f
C757 B.n214 VSUBS 0.006777f
C758 B.n215 VSUBS 0.006777f
C759 B.n216 VSUBS 0.006777f
C760 B.n217 VSUBS 0.006777f
C761 B.n218 VSUBS 0.006777f
C762 B.t8 VSUBS 0.188043f
C763 B.t7 VSUBS 0.209177f
C764 B.t6 VSUBS 0.795368f
C765 B.n219 VSUBS 0.327392f
C766 B.n220 VSUBS 0.229992f
C767 B.n221 VSUBS 0.015701f
C768 B.n222 VSUBS 0.006378f
C769 B.n223 VSUBS 0.006777f
C770 B.n224 VSUBS 0.006777f
C771 B.n225 VSUBS 0.006777f
C772 B.n226 VSUBS 0.006777f
C773 B.n227 VSUBS 0.006777f
C774 B.n228 VSUBS 0.006777f
C775 B.n229 VSUBS 0.006777f
C776 B.n230 VSUBS 0.006777f
C777 B.n231 VSUBS 0.006777f
C778 B.n232 VSUBS 0.006777f
C779 B.n233 VSUBS 0.006777f
C780 B.n234 VSUBS 0.006777f
C781 B.n235 VSUBS 0.006777f
C782 B.n236 VSUBS 0.006777f
C783 B.n237 VSUBS 0.006777f
C784 B.n238 VSUBS 0.003787f
C785 B.n239 VSUBS 0.015701f
C786 B.n240 VSUBS 0.006378f
C787 B.n241 VSUBS 0.006777f
C788 B.n242 VSUBS 0.006777f
C789 B.n243 VSUBS 0.006777f
C790 B.n244 VSUBS 0.006777f
C791 B.n245 VSUBS 0.006777f
C792 B.n246 VSUBS 0.006777f
C793 B.n247 VSUBS 0.006777f
C794 B.n248 VSUBS 0.006777f
C795 B.n249 VSUBS 0.006777f
C796 B.n250 VSUBS 0.006777f
C797 B.n251 VSUBS 0.006777f
C798 B.n252 VSUBS 0.006777f
C799 B.n253 VSUBS 0.006777f
C800 B.n254 VSUBS 0.006777f
C801 B.n255 VSUBS 0.006777f
C802 B.n256 VSUBS 0.006777f
C803 B.n257 VSUBS 0.006777f
C804 B.n258 VSUBS 0.006777f
C805 B.n259 VSUBS 0.006777f
C806 B.n260 VSUBS 0.006777f
C807 B.n261 VSUBS 0.006777f
C808 B.n262 VSUBS 0.006777f
C809 B.n263 VSUBS 0.006777f
C810 B.n264 VSUBS 0.006777f
C811 B.n265 VSUBS 0.006777f
C812 B.n266 VSUBS 0.006777f
C813 B.n267 VSUBS 0.006777f
C814 B.n268 VSUBS 0.006777f
C815 B.n269 VSUBS 0.006777f
C816 B.n270 VSUBS 0.006777f
C817 B.n271 VSUBS 0.006777f
C818 B.n272 VSUBS 0.006777f
C819 B.n273 VSUBS 0.006777f
C820 B.n274 VSUBS 0.006777f
C821 B.n275 VSUBS 0.006777f
C822 B.n276 VSUBS 0.006777f
C823 B.n277 VSUBS 0.006777f
C824 B.n278 VSUBS 0.006777f
C825 B.n279 VSUBS 0.006777f
C826 B.n280 VSUBS 0.006777f
C827 B.n281 VSUBS 0.006777f
C828 B.n282 VSUBS 0.006777f
C829 B.n283 VSUBS 0.006777f
C830 B.n284 VSUBS 0.006777f
C831 B.n285 VSUBS 0.006777f
C832 B.n286 VSUBS 0.006777f
C833 B.n287 VSUBS 0.006777f
C834 B.n288 VSUBS 0.006777f
C835 B.n289 VSUBS 0.006777f
C836 B.n290 VSUBS 0.006777f
C837 B.n291 VSUBS 0.006777f
C838 B.n292 VSUBS 0.006777f
C839 B.n293 VSUBS 0.006777f
C840 B.n294 VSUBS 0.006777f
C841 B.n295 VSUBS 0.006777f
C842 B.n296 VSUBS 0.006777f
C843 B.n297 VSUBS 0.017708f
C844 B.n298 VSUBS 0.016973f
C845 B.n299 VSUBS 0.017674f
C846 B.n300 VSUBS 0.006777f
C847 B.n301 VSUBS 0.006777f
C848 B.n302 VSUBS 0.006777f
C849 B.n303 VSUBS 0.006777f
C850 B.n304 VSUBS 0.006777f
C851 B.n305 VSUBS 0.006777f
C852 B.n306 VSUBS 0.006777f
C853 B.n307 VSUBS 0.006777f
C854 B.n308 VSUBS 0.006777f
C855 B.n309 VSUBS 0.006777f
C856 B.n310 VSUBS 0.006777f
C857 B.n311 VSUBS 0.006777f
C858 B.n312 VSUBS 0.006777f
C859 B.n313 VSUBS 0.006777f
C860 B.n314 VSUBS 0.006777f
C861 B.n315 VSUBS 0.006777f
C862 B.n316 VSUBS 0.006777f
C863 B.n317 VSUBS 0.006777f
C864 B.n318 VSUBS 0.006777f
C865 B.n319 VSUBS 0.006777f
C866 B.n320 VSUBS 0.006777f
C867 B.n321 VSUBS 0.006777f
C868 B.n322 VSUBS 0.006777f
C869 B.n323 VSUBS 0.006777f
C870 B.n324 VSUBS 0.006777f
C871 B.n325 VSUBS 0.006777f
C872 B.n326 VSUBS 0.006777f
C873 B.n327 VSUBS 0.006777f
C874 B.n328 VSUBS 0.006777f
C875 B.n329 VSUBS 0.006777f
C876 B.n330 VSUBS 0.006777f
C877 B.n331 VSUBS 0.006777f
C878 B.n332 VSUBS 0.006777f
C879 B.n333 VSUBS 0.006777f
C880 B.n334 VSUBS 0.006777f
C881 B.n335 VSUBS 0.006777f
C882 B.n336 VSUBS 0.006777f
C883 B.n337 VSUBS 0.006777f
C884 B.n338 VSUBS 0.006777f
C885 B.n339 VSUBS 0.006777f
C886 B.n340 VSUBS 0.006777f
C887 B.n341 VSUBS 0.006777f
C888 B.n342 VSUBS 0.006777f
C889 B.n343 VSUBS 0.006777f
C890 B.n344 VSUBS 0.006777f
C891 B.n345 VSUBS 0.006777f
C892 B.n346 VSUBS 0.006777f
C893 B.n347 VSUBS 0.006777f
C894 B.n348 VSUBS 0.006777f
C895 B.n349 VSUBS 0.006777f
C896 B.n350 VSUBS 0.006777f
C897 B.n351 VSUBS 0.006777f
C898 B.n352 VSUBS 0.006777f
C899 B.n353 VSUBS 0.006777f
C900 B.n354 VSUBS 0.006777f
C901 B.n355 VSUBS 0.006777f
C902 B.n356 VSUBS 0.006777f
C903 B.n357 VSUBS 0.016973f
C904 B.n358 VSUBS 0.017708f
C905 B.n359 VSUBS 0.017708f
C906 B.n360 VSUBS 0.006777f
C907 B.n361 VSUBS 0.006777f
C908 B.n362 VSUBS 0.006777f
C909 B.n363 VSUBS 0.006777f
C910 B.n364 VSUBS 0.006777f
C911 B.n365 VSUBS 0.006777f
C912 B.n366 VSUBS 0.006777f
C913 B.n367 VSUBS 0.006777f
C914 B.n368 VSUBS 0.006777f
C915 B.n369 VSUBS 0.006777f
C916 B.n370 VSUBS 0.006777f
C917 B.n371 VSUBS 0.006777f
C918 B.n372 VSUBS 0.006777f
C919 B.n373 VSUBS 0.006777f
C920 B.n374 VSUBS 0.006777f
C921 B.n375 VSUBS 0.006777f
C922 B.n376 VSUBS 0.006777f
C923 B.n377 VSUBS 0.006777f
C924 B.n378 VSUBS 0.006777f
C925 B.n379 VSUBS 0.006777f
C926 B.n380 VSUBS 0.006777f
C927 B.n381 VSUBS 0.006777f
C928 B.n382 VSUBS 0.006777f
C929 B.n383 VSUBS 0.006777f
C930 B.n384 VSUBS 0.006777f
C931 B.n385 VSUBS 0.006777f
C932 B.n386 VSUBS 0.006777f
C933 B.n387 VSUBS 0.006777f
C934 B.n388 VSUBS 0.006777f
C935 B.n389 VSUBS 0.006777f
C936 B.n390 VSUBS 0.006777f
C937 B.n391 VSUBS 0.006777f
C938 B.n392 VSUBS 0.006777f
C939 B.n393 VSUBS 0.006777f
C940 B.n394 VSUBS 0.006777f
C941 B.n395 VSUBS 0.006777f
C942 B.n396 VSUBS 0.006777f
C943 B.n397 VSUBS 0.006777f
C944 B.n398 VSUBS 0.006777f
C945 B.n399 VSUBS 0.006777f
C946 B.n400 VSUBS 0.006777f
C947 B.n401 VSUBS 0.006777f
C948 B.n402 VSUBS 0.006777f
C949 B.n403 VSUBS 0.006777f
C950 B.n404 VSUBS 0.006777f
C951 B.n405 VSUBS 0.006777f
C952 B.n406 VSUBS 0.006777f
C953 B.n407 VSUBS 0.006777f
C954 B.n408 VSUBS 0.006777f
C955 B.n409 VSUBS 0.006777f
C956 B.n410 VSUBS 0.006777f
C957 B.n411 VSUBS 0.006777f
C958 B.n412 VSUBS 0.006777f
C959 B.n413 VSUBS 0.006777f
C960 B.n414 VSUBS 0.006777f
C961 B.n415 VSUBS 0.006378f
C962 B.n416 VSUBS 0.006777f
C963 B.n417 VSUBS 0.006777f
C964 B.n418 VSUBS 0.003787f
C965 B.n419 VSUBS 0.006777f
C966 B.n420 VSUBS 0.006777f
C967 B.n421 VSUBS 0.006777f
C968 B.n422 VSUBS 0.006777f
C969 B.n423 VSUBS 0.006777f
C970 B.n424 VSUBS 0.006777f
C971 B.n425 VSUBS 0.006777f
C972 B.n426 VSUBS 0.006777f
C973 B.n427 VSUBS 0.006777f
C974 B.n428 VSUBS 0.006777f
C975 B.n429 VSUBS 0.006777f
C976 B.n430 VSUBS 0.006777f
C977 B.n431 VSUBS 0.003787f
C978 B.n432 VSUBS 0.015701f
C979 B.n433 VSUBS 0.006378f
C980 B.n434 VSUBS 0.006777f
C981 B.n435 VSUBS 0.006777f
C982 B.n436 VSUBS 0.006777f
C983 B.n437 VSUBS 0.006777f
C984 B.n438 VSUBS 0.006777f
C985 B.n439 VSUBS 0.006777f
C986 B.n440 VSUBS 0.006777f
C987 B.n441 VSUBS 0.006777f
C988 B.n442 VSUBS 0.006777f
C989 B.n443 VSUBS 0.006777f
C990 B.n444 VSUBS 0.006777f
C991 B.n445 VSUBS 0.006777f
C992 B.n446 VSUBS 0.006777f
C993 B.n447 VSUBS 0.006777f
C994 B.n448 VSUBS 0.006777f
C995 B.n449 VSUBS 0.006777f
C996 B.n450 VSUBS 0.006777f
C997 B.n451 VSUBS 0.006777f
C998 B.n452 VSUBS 0.006777f
C999 B.n453 VSUBS 0.006777f
C1000 B.n454 VSUBS 0.006777f
C1001 B.n455 VSUBS 0.006777f
C1002 B.n456 VSUBS 0.006777f
C1003 B.n457 VSUBS 0.006777f
C1004 B.n458 VSUBS 0.006777f
C1005 B.n459 VSUBS 0.006777f
C1006 B.n460 VSUBS 0.006777f
C1007 B.n461 VSUBS 0.006777f
C1008 B.n462 VSUBS 0.006777f
C1009 B.n463 VSUBS 0.006777f
C1010 B.n464 VSUBS 0.006777f
C1011 B.n465 VSUBS 0.006777f
C1012 B.n466 VSUBS 0.006777f
C1013 B.n467 VSUBS 0.006777f
C1014 B.n468 VSUBS 0.006777f
C1015 B.n469 VSUBS 0.006777f
C1016 B.n470 VSUBS 0.006777f
C1017 B.n471 VSUBS 0.006777f
C1018 B.n472 VSUBS 0.006777f
C1019 B.n473 VSUBS 0.006777f
C1020 B.n474 VSUBS 0.006777f
C1021 B.n475 VSUBS 0.006777f
C1022 B.n476 VSUBS 0.006777f
C1023 B.n477 VSUBS 0.006777f
C1024 B.n478 VSUBS 0.006777f
C1025 B.n479 VSUBS 0.006777f
C1026 B.n480 VSUBS 0.006777f
C1027 B.n481 VSUBS 0.006777f
C1028 B.n482 VSUBS 0.006777f
C1029 B.n483 VSUBS 0.006777f
C1030 B.n484 VSUBS 0.006777f
C1031 B.n485 VSUBS 0.006777f
C1032 B.n486 VSUBS 0.006777f
C1033 B.n487 VSUBS 0.006777f
C1034 B.n488 VSUBS 0.006777f
C1035 B.n489 VSUBS 0.006777f
C1036 B.n490 VSUBS 0.017708f
C1037 B.n491 VSUBS 0.017708f
C1038 B.n492 VSUBS 0.016973f
C1039 B.n493 VSUBS 0.006777f
C1040 B.n494 VSUBS 0.006777f
C1041 B.n495 VSUBS 0.006777f
C1042 B.n496 VSUBS 0.006777f
C1043 B.n497 VSUBS 0.006777f
C1044 B.n498 VSUBS 0.006777f
C1045 B.n499 VSUBS 0.006777f
C1046 B.n500 VSUBS 0.006777f
C1047 B.n501 VSUBS 0.006777f
C1048 B.n502 VSUBS 0.006777f
C1049 B.n503 VSUBS 0.006777f
C1050 B.n504 VSUBS 0.006777f
C1051 B.n505 VSUBS 0.006777f
C1052 B.n506 VSUBS 0.006777f
C1053 B.n507 VSUBS 0.006777f
C1054 B.n508 VSUBS 0.006777f
C1055 B.n509 VSUBS 0.006777f
C1056 B.n510 VSUBS 0.006777f
C1057 B.n511 VSUBS 0.006777f
C1058 B.n512 VSUBS 0.006777f
C1059 B.n513 VSUBS 0.006777f
C1060 B.n514 VSUBS 0.006777f
C1061 B.n515 VSUBS 0.006777f
C1062 B.n516 VSUBS 0.006777f
C1063 B.n517 VSUBS 0.006777f
C1064 B.n518 VSUBS 0.006777f
C1065 B.n519 VSUBS 0.008843f
C1066 B.n520 VSUBS 0.00942f
C1067 B.n521 VSUBS 0.018733f
.ends

