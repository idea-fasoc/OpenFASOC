* NGSPICE file created from diff_pair_sample_0348.ext - technology: sky130A

.subckt diff_pair_sample_0348 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t17 VP.t0 VDD1.t9 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=1.23255 pd=7.8 as=1.23255 ps=7.8 w=7.47 l=3.14
X1 VDD2.t9 VN.t0 VTAIL.t19 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=1.23255 pd=7.8 as=2.9133 ps=15.72 w=7.47 l=3.14
X2 VTAIL.t16 VP.t1 VDD1.t5 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=1.23255 pd=7.8 as=1.23255 ps=7.8 w=7.47 l=3.14
X3 VDD2.t8 VN.t1 VTAIL.t18 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=1.23255 pd=7.8 as=1.23255 ps=7.8 w=7.47 l=3.14
X4 VDD2.t7 VN.t2 VTAIL.t7 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=2.9133 pd=15.72 as=1.23255 ps=7.8 w=7.47 l=3.14
X5 VDD1.t0 VP.t2 VTAIL.t15 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=1.23255 pd=7.8 as=2.9133 ps=15.72 w=7.47 l=3.14
X6 VTAIL.t6 VN.t3 VDD2.t6 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=1.23255 pd=7.8 as=1.23255 ps=7.8 w=7.47 l=3.14
X7 B.t11 B.t9 B.t10 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=2.9133 pd=15.72 as=0 ps=0 w=7.47 l=3.14
X8 VTAIL.t5 VN.t4 VDD2.t5 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=1.23255 pd=7.8 as=1.23255 ps=7.8 w=7.47 l=3.14
X9 VDD1.t8 VP.t3 VTAIL.t14 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=1.23255 pd=7.8 as=2.9133 ps=15.72 w=7.47 l=3.14
X10 VDD2.t4 VN.t5 VTAIL.t0 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=1.23255 pd=7.8 as=2.9133 ps=15.72 w=7.47 l=3.14
X11 B.t8 B.t6 B.t7 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=2.9133 pd=15.72 as=0 ps=0 w=7.47 l=3.14
X12 B.t5 B.t3 B.t4 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=2.9133 pd=15.72 as=0 ps=0 w=7.47 l=3.14
X13 VDD1.t2 VP.t4 VTAIL.t13 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=2.9133 pd=15.72 as=1.23255 ps=7.8 w=7.47 l=3.14
X14 VDD1.t3 VP.t5 VTAIL.t12 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=2.9133 pd=15.72 as=1.23255 ps=7.8 w=7.47 l=3.14
X15 VTAIL.t11 VP.t6 VDD1.t4 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=1.23255 pd=7.8 as=1.23255 ps=7.8 w=7.47 l=3.14
X16 VDD2.t3 VN.t6 VTAIL.t3 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=1.23255 pd=7.8 as=1.23255 ps=7.8 w=7.47 l=3.14
X17 VDD2.t2 VN.t7 VTAIL.t4 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=2.9133 pd=15.72 as=1.23255 ps=7.8 w=7.47 l=3.14
X18 VDD1.t7 VP.t7 VTAIL.t10 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=1.23255 pd=7.8 as=1.23255 ps=7.8 w=7.47 l=3.14
X19 VTAIL.t9 VP.t8 VDD1.t6 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=1.23255 pd=7.8 as=1.23255 ps=7.8 w=7.47 l=3.14
X20 VDD1.t1 VP.t9 VTAIL.t8 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=1.23255 pd=7.8 as=1.23255 ps=7.8 w=7.47 l=3.14
X21 VTAIL.t2 VN.t8 VDD2.t1 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=1.23255 pd=7.8 as=1.23255 ps=7.8 w=7.47 l=3.14
X22 VTAIL.t1 VN.t9 VDD2.t0 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=1.23255 pd=7.8 as=1.23255 ps=7.8 w=7.47 l=3.14
X23 B.t2 B.t0 B.t1 w_n5134_n2462# sky130_fd_pr__pfet_01v8 ad=2.9133 pd=15.72 as=0 ps=0 w=7.47 l=3.14
R0 VP.n29 VP.n28 161.3
R1 VP.n30 VP.n25 161.3
R2 VP.n32 VP.n31 161.3
R3 VP.n33 VP.n24 161.3
R4 VP.n35 VP.n34 161.3
R5 VP.n36 VP.n23 161.3
R6 VP.n38 VP.n37 161.3
R7 VP.n39 VP.n22 161.3
R8 VP.n41 VP.n40 161.3
R9 VP.n42 VP.n21 161.3
R10 VP.n44 VP.n43 161.3
R11 VP.n45 VP.n20 161.3
R12 VP.n47 VP.n46 161.3
R13 VP.n49 VP.n48 161.3
R14 VP.n50 VP.n18 161.3
R15 VP.n52 VP.n51 161.3
R16 VP.n53 VP.n17 161.3
R17 VP.n55 VP.n54 161.3
R18 VP.n56 VP.n16 161.3
R19 VP.n58 VP.n57 161.3
R20 VP.n103 VP.n102 161.3
R21 VP.n101 VP.n1 161.3
R22 VP.n100 VP.n99 161.3
R23 VP.n98 VP.n2 161.3
R24 VP.n97 VP.n96 161.3
R25 VP.n95 VP.n3 161.3
R26 VP.n94 VP.n93 161.3
R27 VP.n92 VP.n91 161.3
R28 VP.n90 VP.n5 161.3
R29 VP.n89 VP.n88 161.3
R30 VP.n87 VP.n6 161.3
R31 VP.n86 VP.n85 161.3
R32 VP.n84 VP.n7 161.3
R33 VP.n83 VP.n82 161.3
R34 VP.n81 VP.n8 161.3
R35 VP.n80 VP.n79 161.3
R36 VP.n78 VP.n9 161.3
R37 VP.n77 VP.n76 161.3
R38 VP.n75 VP.n10 161.3
R39 VP.n74 VP.n73 161.3
R40 VP.n71 VP.n11 161.3
R41 VP.n70 VP.n69 161.3
R42 VP.n68 VP.n12 161.3
R43 VP.n67 VP.n66 161.3
R44 VP.n65 VP.n13 161.3
R45 VP.n64 VP.n63 161.3
R46 VP.n62 VP.n14 161.3
R47 VP.n26 VP.t4 90.7512
R48 VP.n61 VP.n60 68.5364
R49 VP.n104 VP.n0 68.5364
R50 VP.n59 VP.n15 68.5364
R51 VP.n83 VP.t7 57.3339
R52 VP.n60 VP.t5 57.3339
R53 VP.n72 VP.t0 57.3339
R54 VP.n4 VP.t8 57.3339
R55 VP.n0 VP.t3 57.3339
R56 VP.n38 VP.t9 57.3339
R57 VP.n15 VP.t2 57.3339
R58 VP.n19 VP.t6 57.3339
R59 VP.n27 VP.t1 57.3339
R60 VP.n66 VP.n65 56.5193
R61 VP.n78 VP.n77 56.5193
R62 VP.n89 VP.n6 56.5193
R63 VP.n100 VP.n2 56.5193
R64 VP.n55 VP.n17 56.5193
R65 VP.n44 VP.n21 56.5193
R66 VP.n33 VP.n32 56.5193
R67 VP.n61 VP.n59 52.7986
R68 VP.n27 VP.n26 50.9408
R69 VP.n64 VP.n14 24.4675
R70 VP.n65 VP.n64 24.4675
R71 VP.n66 VP.n12 24.4675
R72 VP.n70 VP.n12 24.4675
R73 VP.n71 VP.n70 24.4675
R74 VP.n73 VP.n10 24.4675
R75 VP.n77 VP.n10 24.4675
R76 VP.n79 VP.n78 24.4675
R77 VP.n79 VP.n8 24.4675
R78 VP.n83 VP.n8 24.4675
R79 VP.n84 VP.n83 24.4675
R80 VP.n85 VP.n84 24.4675
R81 VP.n85 VP.n6 24.4675
R82 VP.n90 VP.n89 24.4675
R83 VP.n91 VP.n90 24.4675
R84 VP.n95 VP.n94 24.4675
R85 VP.n96 VP.n95 24.4675
R86 VP.n96 VP.n2 24.4675
R87 VP.n101 VP.n100 24.4675
R88 VP.n102 VP.n101 24.4675
R89 VP.n56 VP.n55 24.4675
R90 VP.n57 VP.n56 24.4675
R91 VP.n45 VP.n44 24.4675
R92 VP.n46 VP.n45 24.4675
R93 VP.n50 VP.n49 24.4675
R94 VP.n51 VP.n50 24.4675
R95 VP.n51 VP.n17 24.4675
R96 VP.n34 VP.n33 24.4675
R97 VP.n34 VP.n23 24.4675
R98 VP.n38 VP.n23 24.4675
R99 VP.n39 VP.n38 24.4675
R100 VP.n40 VP.n39 24.4675
R101 VP.n40 VP.n21 24.4675
R102 VP.n28 VP.n25 24.4675
R103 VP.n32 VP.n25 24.4675
R104 VP.n73 VP.n72 22.9995
R105 VP.n91 VP.n4 22.9995
R106 VP.n46 VP.n19 22.9995
R107 VP.n28 VP.n27 22.9995
R108 VP.n60 VP.n14 21.5315
R109 VP.n102 VP.n0 21.5315
R110 VP.n57 VP.n15 21.5315
R111 VP.n29 VP.n26 3.84097
R112 VP.n72 VP.n71 1.46852
R113 VP.n94 VP.n4 1.46852
R114 VP.n49 VP.n19 1.46852
R115 VP.n59 VP.n58 0.354971
R116 VP.n62 VP.n61 0.354971
R117 VP.n104 VP.n103 0.354971
R118 VP VP.n104 0.26696
R119 VP.n30 VP.n29 0.189894
R120 VP.n31 VP.n30 0.189894
R121 VP.n31 VP.n24 0.189894
R122 VP.n35 VP.n24 0.189894
R123 VP.n36 VP.n35 0.189894
R124 VP.n37 VP.n36 0.189894
R125 VP.n37 VP.n22 0.189894
R126 VP.n41 VP.n22 0.189894
R127 VP.n42 VP.n41 0.189894
R128 VP.n43 VP.n42 0.189894
R129 VP.n43 VP.n20 0.189894
R130 VP.n47 VP.n20 0.189894
R131 VP.n48 VP.n47 0.189894
R132 VP.n48 VP.n18 0.189894
R133 VP.n52 VP.n18 0.189894
R134 VP.n53 VP.n52 0.189894
R135 VP.n54 VP.n53 0.189894
R136 VP.n54 VP.n16 0.189894
R137 VP.n58 VP.n16 0.189894
R138 VP.n63 VP.n62 0.189894
R139 VP.n63 VP.n13 0.189894
R140 VP.n67 VP.n13 0.189894
R141 VP.n68 VP.n67 0.189894
R142 VP.n69 VP.n68 0.189894
R143 VP.n69 VP.n11 0.189894
R144 VP.n74 VP.n11 0.189894
R145 VP.n75 VP.n74 0.189894
R146 VP.n76 VP.n75 0.189894
R147 VP.n76 VP.n9 0.189894
R148 VP.n80 VP.n9 0.189894
R149 VP.n81 VP.n80 0.189894
R150 VP.n82 VP.n81 0.189894
R151 VP.n82 VP.n7 0.189894
R152 VP.n86 VP.n7 0.189894
R153 VP.n87 VP.n86 0.189894
R154 VP.n88 VP.n87 0.189894
R155 VP.n88 VP.n5 0.189894
R156 VP.n92 VP.n5 0.189894
R157 VP.n93 VP.n92 0.189894
R158 VP.n93 VP.n3 0.189894
R159 VP.n97 VP.n3 0.189894
R160 VP.n98 VP.n97 0.189894
R161 VP.n99 VP.n98 0.189894
R162 VP.n99 VP.n1 0.189894
R163 VP.n103 VP.n1 0.189894
R164 VDD1.n34 VDD1.n0 756.745
R165 VDD1.n75 VDD1.n41 756.745
R166 VDD1.n35 VDD1.n34 585
R167 VDD1.n33 VDD1.n32 585
R168 VDD1.n4 VDD1.n3 585
R169 VDD1.n27 VDD1.n26 585
R170 VDD1.n25 VDD1.n24 585
R171 VDD1.n8 VDD1.n7 585
R172 VDD1.n19 VDD1.n18 585
R173 VDD1.n17 VDD1.n16 585
R174 VDD1.n12 VDD1.n11 585
R175 VDD1.n53 VDD1.n52 585
R176 VDD1.n58 VDD1.n57 585
R177 VDD1.n60 VDD1.n59 585
R178 VDD1.n49 VDD1.n48 585
R179 VDD1.n66 VDD1.n65 585
R180 VDD1.n68 VDD1.n67 585
R181 VDD1.n45 VDD1.n44 585
R182 VDD1.n74 VDD1.n73 585
R183 VDD1.n76 VDD1.n75 585
R184 VDD1.n13 VDD1.t2 327.483
R185 VDD1.n54 VDD1.t3 327.483
R186 VDD1.n34 VDD1.n33 171.744
R187 VDD1.n33 VDD1.n3 171.744
R188 VDD1.n26 VDD1.n3 171.744
R189 VDD1.n26 VDD1.n25 171.744
R190 VDD1.n25 VDD1.n7 171.744
R191 VDD1.n18 VDD1.n7 171.744
R192 VDD1.n18 VDD1.n17 171.744
R193 VDD1.n17 VDD1.n11 171.744
R194 VDD1.n58 VDD1.n52 171.744
R195 VDD1.n59 VDD1.n58 171.744
R196 VDD1.n59 VDD1.n48 171.744
R197 VDD1.n66 VDD1.n48 171.744
R198 VDD1.n67 VDD1.n66 171.744
R199 VDD1.n67 VDD1.n44 171.744
R200 VDD1.n74 VDD1.n44 171.744
R201 VDD1.n75 VDD1.n74 171.744
R202 VDD1.n83 VDD1.n82 88.0724
R203 VDD1.n40 VDD1.n39 85.8844
R204 VDD1.n85 VDD1.n84 85.8842
R205 VDD1.n81 VDD1.n80 85.8842
R206 VDD1.t2 VDD1.n11 85.8723
R207 VDD1.t3 VDD1.n52 85.8723
R208 VDD1.n40 VDD1.n38 52.4373
R209 VDD1.n81 VDD1.n79 52.4373
R210 VDD1.n85 VDD1.n83 46.4427
R211 VDD1.n13 VDD1.n12 16.3891
R212 VDD1.n54 VDD1.n53 16.3891
R213 VDD1.n16 VDD1.n15 12.8005
R214 VDD1.n57 VDD1.n56 12.8005
R215 VDD1.n19 VDD1.n10 12.0247
R216 VDD1.n60 VDD1.n51 12.0247
R217 VDD1.n20 VDD1.n8 11.249
R218 VDD1.n61 VDD1.n49 11.249
R219 VDD1.n24 VDD1.n23 10.4732
R220 VDD1.n65 VDD1.n64 10.4732
R221 VDD1.n27 VDD1.n6 9.69747
R222 VDD1.n68 VDD1.n47 9.69747
R223 VDD1.n38 VDD1.n37 9.45567
R224 VDD1.n79 VDD1.n78 9.45567
R225 VDD1.n37 VDD1.n36 9.3005
R226 VDD1.n2 VDD1.n1 9.3005
R227 VDD1.n31 VDD1.n30 9.3005
R228 VDD1.n29 VDD1.n28 9.3005
R229 VDD1.n6 VDD1.n5 9.3005
R230 VDD1.n23 VDD1.n22 9.3005
R231 VDD1.n21 VDD1.n20 9.3005
R232 VDD1.n10 VDD1.n9 9.3005
R233 VDD1.n15 VDD1.n14 9.3005
R234 VDD1.n78 VDD1.n77 9.3005
R235 VDD1.n72 VDD1.n71 9.3005
R236 VDD1.n70 VDD1.n69 9.3005
R237 VDD1.n47 VDD1.n46 9.3005
R238 VDD1.n64 VDD1.n63 9.3005
R239 VDD1.n62 VDD1.n61 9.3005
R240 VDD1.n51 VDD1.n50 9.3005
R241 VDD1.n56 VDD1.n55 9.3005
R242 VDD1.n43 VDD1.n42 9.3005
R243 VDD1.n28 VDD1.n4 8.92171
R244 VDD1.n69 VDD1.n45 8.92171
R245 VDD1.n32 VDD1.n31 8.14595
R246 VDD1.n73 VDD1.n72 8.14595
R247 VDD1.n38 VDD1.n0 7.3702
R248 VDD1.n35 VDD1.n2 7.3702
R249 VDD1.n76 VDD1.n43 7.3702
R250 VDD1.n79 VDD1.n41 7.3702
R251 VDD1.n36 VDD1.n0 6.59444
R252 VDD1.n36 VDD1.n35 6.59444
R253 VDD1.n77 VDD1.n76 6.59444
R254 VDD1.n77 VDD1.n41 6.59444
R255 VDD1.n32 VDD1.n2 5.81868
R256 VDD1.n73 VDD1.n43 5.81868
R257 VDD1.n31 VDD1.n4 5.04292
R258 VDD1.n72 VDD1.n45 5.04292
R259 VDD1.n84 VDD1.t4 4.35191
R260 VDD1.n84 VDD1.t0 4.35191
R261 VDD1.n39 VDD1.t5 4.35191
R262 VDD1.n39 VDD1.t1 4.35191
R263 VDD1.n82 VDD1.t6 4.35191
R264 VDD1.n82 VDD1.t8 4.35191
R265 VDD1.n80 VDD1.t9 4.35191
R266 VDD1.n80 VDD1.t7 4.35191
R267 VDD1.n28 VDD1.n27 4.26717
R268 VDD1.n69 VDD1.n68 4.26717
R269 VDD1.n14 VDD1.n13 3.71019
R270 VDD1.n55 VDD1.n54 3.71019
R271 VDD1.n24 VDD1.n6 3.49141
R272 VDD1.n65 VDD1.n47 3.49141
R273 VDD1.n23 VDD1.n8 2.71565
R274 VDD1.n64 VDD1.n49 2.71565
R275 VDD1 VDD1.n85 2.18584
R276 VDD1.n20 VDD1.n19 1.93989
R277 VDD1.n61 VDD1.n60 1.93989
R278 VDD1.n16 VDD1.n10 1.16414
R279 VDD1.n57 VDD1.n51 1.16414
R280 VDD1 VDD1.n40 0.806535
R281 VDD1.n83 VDD1.n81 0.692999
R282 VDD1.n15 VDD1.n12 0.388379
R283 VDD1.n56 VDD1.n53 0.388379
R284 VDD1.n37 VDD1.n1 0.155672
R285 VDD1.n30 VDD1.n1 0.155672
R286 VDD1.n30 VDD1.n29 0.155672
R287 VDD1.n29 VDD1.n5 0.155672
R288 VDD1.n22 VDD1.n5 0.155672
R289 VDD1.n22 VDD1.n21 0.155672
R290 VDD1.n21 VDD1.n9 0.155672
R291 VDD1.n14 VDD1.n9 0.155672
R292 VDD1.n55 VDD1.n50 0.155672
R293 VDD1.n62 VDD1.n50 0.155672
R294 VDD1.n63 VDD1.n62 0.155672
R295 VDD1.n63 VDD1.n46 0.155672
R296 VDD1.n70 VDD1.n46 0.155672
R297 VDD1.n71 VDD1.n70 0.155672
R298 VDD1.n71 VDD1.n42 0.155672
R299 VDD1.n78 VDD1.n42 0.155672
R300 VTAIL.n168 VTAIL.n134 756.745
R301 VTAIL.n36 VTAIL.n2 756.745
R302 VTAIL.n128 VTAIL.n94 756.745
R303 VTAIL.n84 VTAIL.n50 756.745
R304 VTAIL.n146 VTAIL.n145 585
R305 VTAIL.n151 VTAIL.n150 585
R306 VTAIL.n153 VTAIL.n152 585
R307 VTAIL.n142 VTAIL.n141 585
R308 VTAIL.n159 VTAIL.n158 585
R309 VTAIL.n161 VTAIL.n160 585
R310 VTAIL.n138 VTAIL.n137 585
R311 VTAIL.n167 VTAIL.n166 585
R312 VTAIL.n169 VTAIL.n168 585
R313 VTAIL.n14 VTAIL.n13 585
R314 VTAIL.n19 VTAIL.n18 585
R315 VTAIL.n21 VTAIL.n20 585
R316 VTAIL.n10 VTAIL.n9 585
R317 VTAIL.n27 VTAIL.n26 585
R318 VTAIL.n29 VTAIL.n28 585
R319 VTAIL.n6 VTAIL.n5 585
R320 VTAIL.n35 VTAIL.n34 585
R321 VTAIL.n37 VTAIL.n36 585
R322 VTAIL.n129 VTAIL.n128 585
R323 VTAIL.n127 VTAIL.n126 585
R324 VTAIL.n98 VTAIL.n97 585
R325 VTAIL.n121 VTAIL.n120 585
R326 VTAIL.n119 VTAIL.n118 585
R327 VTAIL.n102 VTAIL.n101 585
R328 VTAIL.n113 VTAIL.n112 585
R329 VTAIL.n111 VTAIL.n110 585
R330 VTAIL.n106 VTAIL.n105 585
R331 VTAIL.n85 VTAIL.n84 585
R332 VTAIL.n83 VTAIL.n82 585
R333 VTAIL.n54 VTAIL.n53 585
R334 VTAIL.n77 VTAIL.n76 585
R335 VTAIL.n75 VTAIL.n74 585
R336 VTAIL.n58 VTAIL.n57 585
R337 VTAIL.n69 VTAIL.n68 585
R338 VTAIL.n67 VTAIL.n66 585
R339 VTAIL.n62 VTAIL.n61 585
R340 VTAIL.n147 VTAIL.t19 327.483
R341 VTAIL.n15 VTAIL.t14 327.483
R342 VTAIL.n107 VTAIL.t15 327.483
R343 VTAIL.n63 VTAIL.t0 327.483
R344 VTAIL.n151 VTAIL.n145 171.744
R345 VTAIL.n152 VTAIL.n151 171.744
R346 VTAIL.n152 VTAIL.n141 171.744
R347 VTAIL.n159 VTAIL.n141 171.744
R348 VTAIL.n160 VTAIL.n159 171.744
R349 VTAIL.n160 VTAIL.n137 171.744
R350 VTAIL.n167 VTAIL.n137 171.744
R351 VTAIL.n168 VTAIL.n167 171.744
R352 VTAIL.n19 VTAIL.n13 171.744
R353 VTAIL.n20 VTAIL.n19 171.744
R354 VTAIL.n20 VTAIL.n9 171.744
R355 VTAIL.n27 VTAIL.n9 171.744
R356 VTAIL.n28 VTAIL.n27 171.744
R357 VTAIL.n28 VTAIL.n5 171.744
R358 VTAIL.n35 VTAIL.n5 171.744
R359 VTAIL.n36 VTAIL.n35 171.744
R360 VTAIL.n128 VTAIL.n127 171.744
R361 VTAIL.n127 VTAIL.n97 171.744
R362 VTAIL.n120 VTAIL.n97 171.744
R363 VTAIL.n120 VTAIL.n119 171.744
R364 VTAIL.n119 VTAIL.n101 171.744
R365 VTAIL.n112 VTAIL.n101 171.744
R366 VTAIL.n112 VTAIL.n111 171.744
R367 VTAIL.n111 VTAIL.n105 171.744
R368 VTAIL.n84 VTAIL.n83 171.744
R369 VTAIL.n83 VTAIL.n53 171.744
R370 VTAIL.n76 VTAIL.n53 171.744
R371 VTAIL.n76 VTAIL.n75 171.744
R372 VTAIL.n75 VTAIL.n57 171.744
R373 VTAIL.n68 VTAIL.n57 171.744
R374 VTAIL.n68 VTAIL.n67 171.744
R375 VTAIL.n67 VTAIL.n61 171.744
R376 VTAIL.t19 VTAIL.n145 85.8723
R377 VTAIL.t14 VTAIL.n13 85.8723
R378 VTAIL.t15 VTAIL.n105 85.8723
R379 VTAIL.t0 VTAIL.n61 85.8723
R380 VTAIL.n93 VTAIL.n92 69.2056
R381 VTAIL.n91 VTAIL.n90 69.2056
R382 VTAIL.n49 VTAIL.n48 69.2056
R383 VTAIL.n47 VTAIL.n46 69.2056
R384 VTAIL.n175 VTAIL.n174 69.2054
R385 VTAIL.n1 VTAIL.n0 69.2054
R386 VTAIL.n43 VTAIL.n42 69.2054
R387 VTAIL.n45 VTAIL.n44 69.2054
R388 VTAIL.n173 VTAIL.n172 32.7672
R389 VTAIL.n41 VTAIL.n40 32.7672
R390 VTAIL.n133 VTAIL.n132 32.7672
R391 VTAIL.n89 VTAIL.n88 32.7672
R392 VTAIL.n47 VTAIL.n45 24.7893
R393 VTAIL.n173 VTAIL.n133 21.7979
R394 VTAIL.n147 VTAIL.n146 16.3891
R395 VTAIL.n15 VTAIL.n14 16.3891
R396 VTAIL.n107 VTAIL.n106 16.3891
R397 VTAIL.n63 VTAIL.n62 16.3891
R398 VTAIL.n150 VTAIL.n149 12.8005
R399 VTAIL.n18 VTAIL.n17 12.8005
R400 VTAIL.n110 VTAIL.n109 12.8005
R401 VTAIL.n66 VTAIL.n65 12.8005
R402 VTAIL.n153 VTAIL.n144 12.0247
R403 VTAIL.n21 VTAIL.n12 12.0247
R404 VTAIL.n113 VTAIL.n104 12.0247
R405 VTAIL.n69 VTAIL.n60 12.0247
R406 VTAIL.n154 VTAIL.n142 11.249
R407 VTAIL.n22 VTAIL.n10 11.249
R408 VTAIL.n114 VTAIL.n102 11.249
R409 VTAIL.n70 VTAIL.n58 11.249
R410 VTAIL.n158 VTAIL.n157 10.4732
R411 VTAIL.n26 VTAIL.n25 10.4732
R412 VTAIL.n118 VTAIL.n117 10.4732
R413 VTAIL.n74 VTAIL.n73 10.4732
R414 VTAIL.n161 VTAIL.n140 9.69747
R415 VTAIL.n29 VTAIL.n8 9.69747
R416 VTAIL.n121 VTAIL.n100 9.69747
R417 VTAIL.n77 VTAIL.n56 9.69747
R418 VTAIL.n172 VTAIL.n171 9.45567
R419 VTAIL.n40 VTAIL.n39 9.45567
R420 VTAIL.n132 VTAIL.n131 9.45567
R421 VTAIL.n88 VTAIL.n87 9.45567
R422 VTAIL.n171 VTAIL.n170 9.3005
R423 VTAIL.n165 VTAIL.n164 9.3005
R424 VTAIL.n163 VTAIL.n162 9.3005
R425 VTAIL.n140 VTAIL.n139 9.3005
R426 VTAIL.n157 VTAIL.n156 9.3005
R427 VTAIL.n155 VTAIL.n154 9.3005
R428 VTAIL.n144 VTAIL.n143 9.3005
R429 VTAIL.n149 VTAIL.n148 9.3005
R430 VTAIL.n136 VTAIL.n135 9.3005
R431 VTAIL.n39 VTAIL.n38 9.3005
R432 VTAIL.n33 VTAIL.n32 9.3005
R433 VTAIL.n31 VTAIL.n30 9.3005
R434 VTAIL.n8 VTAIL.n7 9.3005
R435 VTAIL.n25 VTAIL.n24 9.3005
R436 VTAIL.n23 VTAIL.n22 9.3005
R437 VTAIL.n12 VTAIL.n11 9.3005
R438 VTAIL.n17 VTAIL.n16 9.3005
R439 VTAIL.n4 VTAIL.n3 9.3005
R440 VTAIL.n131 VTAIL.n130 9.3005
R441 VTAIL.n96 VTAIL.n95 9.3005
R442 VTAIL.n125 VTAIL.n124 9.3005
R443 VTAIL.n123 VTAIL.n122 9.3005
R444 VTAIL.n100 VTAIL.n99 9.3005
R445 VTAIL.n117 VTAIL.n116 9.3005
R446 VTAIL.n115 VTAIL.n114 9.3005
R447 VTAIL.n104 VTAIL.n103 9.3005
R448 VTAIL.n109 VTAIL.n108 9.3005
R449 VTAIL.n87 VTAIL.n86 9.3005
R450 VTAIL.n52 VTAIL.n51 9.3005
R451 VTAIL.n81 VTAIL.n80 9.3005
R452 VTAIL.n79 VTAIL.n78 9.3005
R453 VTAIL.n56 VTAIL.n55 9.3005
R454 VTAIL.n73 VTAIL.n72 9.3005
R455 VTAIL.n71 VTAIL.n70 9.3005
R456 VTAIL.n60 VTAIL.n59 9.3005
R457 VTAIL.n65 VTAIL.n64 9.3005
R458 VTAIL.n162 VTAIL.n138 8.92171
R459 VTAIL.n30 VTAIL.n6 8.92171
R460 VTAIL.n122 VTAIL.n98 8.92171
R461 VTAIL.n78 VTAIL.n54 8.92171
R462 VTAIL.n166 VTAIL.n165 8.14595
R463 VTAIL.n34 VTAIL.n33 8.14595
R464 VTAIL.n126 VTAIL.n125 8.14595
R465 VTAIL.n82 VTAIL.n81 8.14595
R466 VTAIL.n169 VTAIL.n136 7.3702
R467 VTAIL.n172 VTAIL.n134 7.3702
R468 VTAIL.n37 VTAIL.n4 7.3702
R469 VTAIL.n40 VTAIL.n2 7.3702
R470 VTAIL.n132 VTAIL.n94 7.3702
R471 VTAIL.n129 VTAIL.n96 7.3702
R472 VTAIL.n88 VTAIL.n50 7.3702
R473 VTAIL.n85 VTAIL.n52 7.3702
R474 VTAIL.n170 VTAIL.n169 6.59444
R475 VTAIL.n170 VTAIL.n134 6.59444
R476 VTAIL.n38 VTAIL.n37 6.59444
R477 VTAIL.n38 VTAIL.n2 6.59444
R478 VTAIL.n130 VTAIL.n94 6.59444
R479 VTAIL.n130 VTAIL.n129 6.59444
R480 VTAIL.n86 VTAIL.n50 6.59444
R481 VTAIL.n86 VTAIL.n85 6.59444
R482 VTAIL.n166 VTAIL.n136 5.81868
R483 VTAIL.n34 VTAIL.n4 5.81868
R484 VTAIL.n126 VTAIL.n96 5.81868
R485 VTAIL.n82 VTAIL.n52 5.81868
R486 VTAIL.n165 VTAIL.n138 5.04292
R487 VTAIL.n33 VTAIL.n6 5.04292
R488 VTAIL.n125 VTAIL.n98 5.04292
R489 VTAIL.n81 VTAIL.n54 5.04292
R490 VTAIL.n174 VTAIL.t3 4.35191
R491 VTAIL.n174 VTAIL.t2 4.35191
R492 VTAIL.n0 VTAIL.t7 4.35191
R493 VTAIL.n0 VTAIL.t5 4.35191
R494 VTAIL.n42 VTAIL.t10 4.35191
R495 VTAIL.n42 VTAIL.t9 4.35191
R496 VTAIL.n44 VTAIL.t12 4.35191
R497 VTAIL.n44 VTAIL.t17 4.35191
R498 VTAIL.n92 VTAIL.t8 4.35191
R499 VTAIL.n92 VTAIL.t11 4.35191
R500 VTAIL.n90 VTAIL.t13 4.35191
R501 VTAIL.n90 VTAIL.t16 4.35191
R502 VTAIL.n48 VTAIL.t18 4.35191
R503 VTAIL.n48 VTAIL.t6 4.35191
R504 VTAIL.n46 VTAIL.t4 4.35191
R505 VTAIL.n46 VTAIL.t1 4.35191
R506 VTAIL.n162 VTAIL.n161 4.26717
R507 VTAIL.n30 VTAIL.n29 4.26717
R508 VTAIL.n122 VTAIL.n121 4.26717
R509 VTAIL.n78 VTAIL.n77 4.26717
R510 VTAIL.n148 VTAIL.n147 3.71019
R511 VTAIL.n16 VTAIL.n15 3.71019
R512 VTAIL.n108 VTAIL.n107 3.71019
R513 VTAIL.n64 VTAIL.n63 3.71019
R514 VTAIL.n158 VTAIL.n140 3.49141
R515 VTAIL.n26 VTAIL.n8 3.49141
R516 VTAIL.n118 VTAIL.n100 3.49141
R517 VTAIL.n74 VTAIL.n56 3.49141
R518 VTAIL.n49 VTAIL.n47 2.99188
R519 VTAIL.n89 VTAIL.n49 2.99188
R520 VTAIL.n93 VTAIL.n91 2.99188
R521 VTAIL.n133 VTAIL.n93 2.99188
R522 VTAIL.n45 VTAIL.n43 2.99188
R523 VTAIL.n43 VTAIL.n41 2.99188
R524 VTAIL.n175 VTAIL.n173 2.99188
R525 VTAIL.n157 VTAIL.n142 2.71565
R526 VTAIL.n25 VTAIL.n10 2.71565
R527 VTAIL.n117 VTAIL.n102 2.71565
R528 VTAIL.n73 VTAIL.n58 2.71565
R529 VTAIL VTAIL.n1 2.30222
R530 VTAIL.n91 VTAIL.n89 1.96602
R531 VTAIL.n41 VTAIL.n1 1.96602
R532 VTAIL.n154 VTAIL.n153 1.93989
R533 VTAIL.n22 VTAIL.n21 1.93989
R534 VTAIL.n114 VTAIL.n113 1.93989
R535 VTAIL.n70 VTAIL.n69 1.93989
R536 VTAIL.n150 VTAIL.n144 1.16414
R537 VTAIL.n18 VTAIL.n12 1.16414
R538 VTAIL.n110 VTAIL.n104 1.16414
R539 VTAIL.n66 VTAIL.n60 1.16414
R540 VTAIL VTAIL.n175 0.690155
R541 VTAIL.n149 VTAIL.n146 0.388379
R542 VTAIL.n17 VTAIL.n14 0.388379
R543 VTAIL.n109 VTAIL.n106 0.388379
R544 VTAIL.n65 VTAIL.n62 0.388379
R545 VTAIL.n148 VTAIL.n143 0.155672
R546 VTAIL.n155 VTAIL.n143 0.155672
R547 VTAIL.n156 VTAIL.n155 0.155672
R548 VTAIL.n156 VTAIL.n139 0.155672
R549 VTAIL.n163 VTAIL.n139 0.155672
R550 VTAIL.n164 VTAIL.n163 0.155672
R551 VTAIL.n164 VTAIL.n135 0.155672
R552 VTAIL.n171 VTAIL.n135 0.155672
R553 VTAIL.n16 VTAIL.n11 0.155672
R554 VTAIL.n23 VTAIL.n11 0.155672
R555 VTAIL.n24 VTAIL.n23 0.155672
R556 VTAIL.n24 VTAIL.n7 0.155672
R557 VTAIL.n31 VTAIL.n7 0.155672
R558 VTAIL.n32 VTAIL.n31 0.155672
R559 VTAIL.n32 VTAIL.n3 0.155672
R560 VTAIL.n39 VTAIL.n3 0.155672
R561 VTAIL.n131 VTAIL.n95 0.155672
R562 VTAIL.n124 VTAIL.n95 0.155672
R563 VTAIL.n124 VTAIL.n123 0.155672
R564 VTAIL.n123 VTAIL.n99 0.155672
R565 VTAIL.n116 VTAIL.n99 0.155672
R566 VTAIL.n116 VTAIL.n115 0.155672
R567 VTAIL.n115 VTAIL.n103 0.155672
R568 VTAIL.n108 VTAIL.n103 0.155672
R569 VTAIL.n87 VTAIL.n51 0.155672
R570 VTAIL.n80 VTAIL.n51 0.155672
R571 VTAIL.n80 VTAIL.n79 0.155672
R572 VTAIL.n79 VTAIL.n55 0.155672
R573 VTAIL.n72 VTAIL.n55 0.155672
R574 VTAIL.n72 VTAIL.n71 0.155672
R575 VTAIL.n71 VTAIL.n59 0.155672
R576 VTAIL.n64 VTAIL.n59 0.155672
R577 VN.n88 VN.n87 161.3
R578 VN.n86 VN.n46 161.3
R579 VN.n85 VN.n84 161.3
R580 VN.n83 VN.n47 161.3
R581 VN.n82 VN.n81 161.3
R582 VN.n80 VN.n48 161.3
R583 VN.n79 VN.n78 161.3
R584 VN.n77 VN.n76 161.3
R585 VN.n75 VN.n50 161.3
R586 VN.n74 VN.n73 161.3
R587 VN.n72 VN.n51 161.3
R588 VN.n71 VN.n70 161.3
R589 VN.n69 VN.n52 161.3
R590 VN.n68 VN.n67 161.3
R591 VN.n66 VN.n53 161.3
R592 VN.n65 VN.n64 161.3
R593 VN.n63 VN.n54 161.3
R594 VN.n62 VN.n61 161.3
R595 VN.n60 VN.n55 161.3
R596 VN.n59 VN.n58 161.3
R597 VN.n43 VN.n42 161.3
R598 VN.n41 VN.n1 161.3
R599 VN.n40 VN.n39 161.3
R600 VN.n38 VN.n2 161.3
R601 VN.n37 VN.n36 161.3
R602 VN.n35 VN.n3 161.3
R603 VN.n34 VN.n33 161.3
R604 VN.n32 VN.n31 161.3
R605 VN.n30 VN.n5 161.3
R606 VN.n29 VN.n28 161.3
R607 VN.n27 VN.n6 161.3
R608 VN.n26 VN.n25 161.3
R609 VN.n24 VN.n7 161.3
R610 VN.n23 VN.n22 161.3
R611 VN.n21 VN.n8 161.3
R612 VN.n20 VN.n19 161.3
R613 VN.n18 VN.n9 161.3
R614 VN.n17 VN.n16 161.3
R615 VN.n15 VN.n10 161.3
R616 VN.n14 VN.n13 161.3
R617 VN.n56 VN.t5 90.7515
R618 VN.n11 VN.t2 90.7515
R619 VN.n44 VN.n0 68.5364
R620 VN.n89 VN.n45 68.5364
R621 VN.n23 VN.t6 57.3339
R622 VN.n12 VN.t4 57.3339
R623 VN.n4 VN.t8 57.3339
R624 VN.n0 VN.t0 57.3339
R625 VN.n68 VN.t1 57.3339
R626 VN.n57 VN.t3 57.3339
R627 VN.n49 VN.t9 57.3339
R628 VN.n45 VN.t7 57.3339
R629 VN.n18 VN.n17 56.5193
R630 VN.n29 VN.n6 56.5193
R631 VN.n40 VN.n2 56.5193
R632 VN.n63 VN.n62 56.5193
R633 VN.n74 VN.n51 56.5193
R634 VN.n85 VN.n47 56.5193
R635 VN VN.n89 52.9639
R636 VN.n12 VN.n11 50.9408
R637 VN.n57 VN.n56 50.9408
R638 VN.n13 VN.n10 24.4675
R639 VN.n17 VN.n10 24.4675
R640 VN.n19 VN.n18 24.4675
R641 VN.n19 VN.n8 24.4675
R642 VN.n23 VN.n8 24.4675
R643 VN.n24 VN.n23 24.4675
R644 VN.n25 VN.n24 24.4675
R645 VN.n25 VN.n6 24.4675
R646 VN.n30 VN.n29 24.4675
R647 VN.n31 VN.n30 24.4675
R648 VN.n35 VN.n34 24.4675
R649 VN.n36 VN.n35 24.4675
R650 VN.n36 VN.n2 24.4675
R651 VN.n41 VN.n40 24.4675
R652 VN.n42 VN.n41 24.4675
R653 VN.n62 VN.n55 24.4675
R654 VN.n58 VN.n55 24.4675
R655 VN.n70 VN.n51 24.4675
R656 VN.n70 VN.n69 24.4675
R657 VN.n69 VN.n68 24.4675
R658 VN.n68 VN.n53 24.4675
R659 VN.n64 VN.n53 24.4675
R660 VN.n64 VN.n63 24.4675
R661 VN.n81 VN.n47 24.4675
R662 VN.n81 VN.n80 24.4675
R663 VN.n80 VN.n79 24.4675
R664 VN.n76 VN.n75 24.4675
R665 VN.n75 VN.n74 24.4675
R666 VN.n87 VN.n86 24.4675
R667 VN.n86 VN.n85 24.4675
R668 VN.n13 VN.n12 22.9995
R669 VN.n31 VN.n4 22.9995
R670 VN.n58 VN.n57 22.9995
R671 VN.n76 VN.n49 22.9995
R672 VN.n42 VN.n0 21.5315
R673 VN.n87 VN.n45 21.5315
R674 VN.n59 VN.n56 3.84099
R675 VN.n14 VN.n11 3.84099
R676 VN.n34 VN.n4 1.46852
R677 VN.n79 VN.n49 1.46852
R678 VN.n89 VN.n88 0.354971
R679 VN.n44 VN.n43 0.354971
R680 VN VN.n44 0.26696
R681 VN.n88 VN.n46 0.189894
R682 VN.n84 VN.n46 0.189894
R683 VN.n84 VN.n83 0.189894
R684 VN.n83 VN.n82 0.189894
R685 VN.n82 VN.n48 0.189894
R686 VN.n78 VN.n48 0.189894
R687 VN.n78 VN.n77 0.189894
R688 VN.n77 VN.n50 0.189894
R689 VN.n73 VN.n50 0.189894
R690 VN.n73 VN.n72 0.189894
R691 VN.n72 VN.n71 0.189894
R692 VN.n71 VN.n52 0.189894
R693 VN.n67 VN.n52 0.189894
R694 VN.n67 VN.n66 0.189894
R695 VN.n66 VN.n65 0.189894
R696 VN.n65 VN.n54 0.189894
R697 VN.n61 VN.n54 0.189894
R698 VN.n61 VN.n60 0.189894
R699 VN.n60 VN.n59 0.189894
R700 VN.n15 VN.n14 0.189894
R701 VN.n16 VN.n15 0.189894
R702 VN.n16 VN.n9 0.189894
R703 VN.n20 VN.n9 0.189894
R704 VN.n21 VN.n20 0.189894
R705 VN.n22 VN.n21 0.189894
R706 VN.n22 VN.n7 0.189894
R707 VN.n26 VN.n7 0.189894
R708 VN.n27 VN.n26 0.189894
R709 VN.n28 VN.n27 0.189894
R710 VN.n28 VN.n5 0.189894
R711 VN.n32 VN.n5 0.189894
R712 VN.n33 VN.n32 0.189894
R713 VN.n33 VN.n3 0.189894
R714 VN.n37 VN.n3 0.189894
R715 VN.n38 VN.n37 0.189894
R716 VN.n39 VN.n38 0.189894
R717 VN.n39 VN.n1 0.189894
R718 VN.n43 VN.n1 0.189894
R719 VDD2.n77 VDD2.n43 756.745
R720 VDD2.n34 VDD2.n0 756.745
R721 VDD2.n78 VDD2.n77 585
R722 VDD2.n76 VDD2.n75 585
R723 VDD2.n47 VDD2.n46 585
R724 VDD2.n70 VDD2.n69 585
R725 VDD2.n68 VDD2.n67 585
R726 VDD2.n51 VDD2.n50 585
R727 VDD2.n62 VDD2.n61 585
R728 VDD2.n60 VDD2.n59 585
R729 VDD2.n55 VDD2.n54 585
R730 VDD2.n12 VDD2.n11 585
R731 VDD2.n17 VDD2.n16 585
R732 VDD2.n19 VDD2.n18 585
R733 VDD2.n8 VDD2.n7 585
R734 VDD2.n25 VDD2.n24 585
R735 VDD2.n27 VDD2.n26 585
R736 VDD2.n4 VDD2.n3 585
R737 VDD2.n33 VDD2.n32 585
R738 VDD2.n35 VDD2.n34 585
R739 VDD2.n56 VDD2.t2 327.483
R740 VDD2.n13 VDD2.t7 327.483
R741 VDD2.n77 VDD2.n76 171.744
R742 VDD2.n76 VDD2.n46 171.744
R743 VDD2.n69 VDD2.n46 171.744
R744 VDD2.n69 VDD2.n68 171.744
R745 VDD2.n68 VDD2.n50 171.744
R746 VDD2.n61 VDD2.n50 171.744
R747 VDD2.n61 VDD2.n60 171.744
R748 VDD2.n60 VDD2.n54 171.744
R749 VDD2.n17 VDD2.n11 171.744
R750 VDD2.n18 VDD2.n17 171.744
R751 VDD2.n18 VDD2.n7 171.744
R752 VDD2.n25 VDD2.n7 171.744
R753 VDD2.n26 VDD2.n25 171.744
R754 VDD2.n26 VDD2.n3 171.744
R755 VDD2.n33 VDD2.n3 171.744
R756 VDD2.n34 VDD2.n33 171.744
R757 VDD2.n42 VDD2.n41 88.0724
R758 VDD2 VDD2.n85 88.0695
R759 VDD2.n84 VDD2.n83 85.8844
R760 VDD2.n40 VDD2.n39 85.8842
R761 VDD2.t2 VDD2.n54 85.8723
R762 VDD2.t7 VDD2.n11 85.8723
R763 VDD2.n40 VDD2.n38 52.4373
R764 VDD2.n82 VDD2.n81 49.446
R765 VDD2.n82 VDD2.n42 44.364
R766 VDD2.n56 VDD2.n55 16.3891
R767 VDD2.n13 VDD2.n12 16.3891
R768 VDD2.n59 VDD2.n58 12.8005
R769 VDD2.n16 VDD2.n15 12.8005
R770 VDD2.n62 VDD2.n53 12.0247
R771 VDD2.n19 VDD2.n10 12.0247
R772 VDD2.n63 VDD2.n51 11.249
R773 VDD2.n20 VDD2.n8 11.249
R774 VDD2.n67 VDD2.n66 10.4732
R775 VDD2.n24 VDD2.n23 10.4732
R776 VDD2.n70 VDD2.n49 9.69747
R777 VDD2.n27 VDD2.n6 9.69747
R778 VDD2.n81 VDD2.n80 9.45567
R779 VDD2.n38 VDD2.n37 9.45567
R780 VDD2.n80 VDD2.n79 9.3005
R781 VDD2.n45 VDD2.n44 9.3005
R782 VDD2.n74 VDD2.n73 9.3005
R783 VDD2.n72 VDD2.n71 9.3005
R784 VDD2.n49 VDD2.n48 9.3005
R785 VDD2.n66 VDD2.n65 9.3005
R786 VDD2.n64 VDD2.n63 9.3005
R787 VDD2.n53 VDD2.n52 9.3005
R788 VDD2.n58 VDD2.n57 9.3005
R789 VDD2.n37 VDD2.n36 9.3005
R790 VDD2.n31 VDD2.n30 9.3005
R791 VDD2.n29 VDD2.n28 9.3005
R792 VDD2.n6 VDD2.n5 9.3005
R793 VDD2.n23 VDD2.n22 9.3005
R794 VDD2.n21 VDD2.n20 9.3005
R795 VDD2.n10 VDD2.n9 9.3005
R796 VDD2.n15 VDD2.n14 9.3005
R797 VDD2.n2 VDD2.n1 9.3005
R798 VDD2.n71 VDD2.n47 8.92171
R799 VDD2.n28 VDD2.n4 8.92171
R800 VDD2.n75 VDD2.n74 8.14595
R801 VDD2.n32 VDD2.n31 8.14595
R802 VDD2.n81 VDD2.n43 7.3702
R803 VDD2.n78 VDD2.n45 7.3702
R804 VDD2.n35 VDD2.n2 7.3702
R805 VDD2.n38 VDD2.n0 7.3702
R806 VDD2.n79 VDD2.n43 6.59444
R807 VDD2.n79 VDD2.n78 6.59444
R808 VDD2.n36 VDD2.n35 6.59444
R809 VDD2.n36 VDD2.n0 6.59444
R810 VDD2.n75 VDD2.n45 5.81868
R811 VDD2.n32 VDD2.n2 5.81868
R812 VDD2.n74 VDD2.n47 5.04292
R813 VDD2.n31 VDD2.n4 5.04292
R814 VDD2.n85 VDD2.t6 4.35191
R815 VDD2.n85 VDD2.t4 4.35191
R816 VDD2.n83 VDD2.t0 4.35191
R817 VDD2.n83 VDD2.t8 4.35191
R818 VDD2.n41 VDD2.t1 4.35191
R819 VDD2.n41 VDD2.t9 4.35191
R820 VDD2.n39 VDD2.t5 4.35191
R821 VDD2.n39 VDD2.t3 4.35191
R822 VDD2.n71 VDD2.n70 4.26717
R823 VDD2.n28 VDD2.n27 4.26717
R824 VDD2.n57 VDD2.n56 3.71019
R825 VDD2.n14 VDD2.n13 3.71019
R826 VDD2.n67 VDD2.n49 3.49141
R827 VDD2.n24 VDD2.n6 3.49141
R828 VDD2.n84 VDD2.n82 2.99188
R829 VDD2.n66 VDD2.n51 2.71565
R830 VDD2.n23 VDD2.n8 2.71565
R831 VDD2.n63 VDD2.n62 1.93989
R832 VDD2.n20 VDD2.n19 1.93989
R833 VDD2.n59 VDD2.n53 1.16414
R834 VDD2.n16 VDD2.n10 1.16414
R835 VDD2 VDD2.n84 0.806535
R836 VDD2.n42 VDD2.n40 0.692999
R837 VDD2.n58 VDD2.n55 0.388379
R838 VDD2.n15 VDD2.n12 0.388379
R839 VDD2.n80 VDD2.n44 0.155672
R840 VDD2.n73 VDD2.n44 0.155672
R841 VDD2.n73 VDD2.n72 0.155672
R842 VDD2.n72 VDD2.n48 0.155672
R843 VDD2.n65 VDD2.n48 0.155672
R844 VDD2.n65 VDD2.n64 0.155672
R845 VDD2.n64 VDD2.n52 0.155672
R846 VDD2.n57 VDD2.n52 0.155672
R847 VDD2.n14 VDD2.n9 0.155672
R848 VDD2.n21 VDD2.n9 0.155672
R849 VDD2.n22 VDD2.n21 0.155672
R850 VDD2.n22 VDD2.n5 0.155672
R851 VDD2.n29 VDD2.n5 0.155672
R852 VDD2.n30 VDD2.n29 0.155672
R853 VDD2.n30 VDD2.n1 0.155672
R854 VDD2.n37 VDD2.n1 0.155672
R855 B.n418 B.n417 585
R856 B.n416 B.n145 585
R857 B.n415 B.n414 585
R858 B.n413 B.n146 585
R859 B.n412 B.n411 585
R860 B.n410 B.n147 585
R861 B.n409 B.n408 585
R862 B.n407 B.n148 585
R863 B.n406 B.n405 585
R864 B.n404 B.n149 585
R865 B.n403 B.n402 585
R866 B.n401 B.n150 585
R867 B.n400 B.n399 585
R868 B.n398 B.n151 585
R869 B.n397 B.n396 585
R870 B.n395 B.n152 585
R871 B.n394 B.n393 585
R872 B.n392 B.n153 585
R873 B.n391 B.n390 585
R874 B.n389 B.n154 585
R875 B.n388 B.n387 585
R876 B.n386 B.n155 585
R877 B.n385 B.n384 585
R878 B.n383 B.n156 585
R879 B.n382 B.n381 585
R880 B.n380 B.n157 585
R881 B.n379 B.n378 585
R882 B.n377 B.n158 585
R883 B.n375 B.n374 585
R884 B.n373 B.n161 585
R885 B.n372 B.n371 585
R886 B.n370 B.n162 585
R887 B.n369 B.n368 585
R888 B.n367 B.n163 585
R889 B.n366 B.n365 585
R890 B.n364 B.n164 585
R891 B.n363 B.n362 585
R892 B.n361 B.n165 585
R893 B.n360 B.n359 585
R894 B.n355 B.n166 585
R895 B.n354 B.n353 585
R896 B.n352 B.n167 585
R897 B.n351 B.n350 585
R898 B.n349 B.n168 585
R899 B.n348 B.n347 585
R900 B.n346 B.n169 585
R901 B.n345 B.n344 585
R902 B.n343 B.n170 585
R903 B.n342 B.n341 585
R904 B.n340 B.n171 585
R905 B.n339 B.n338 585
R906 B.n337 B.n172 585
R907 B.n336 B.n335 585
R908 B.n334 B.n173 585
R909 B.n333 B.n332 585
R910 B.n331 B.n174 585
R911 B.n330 B.n329 585
R912 B.n328 B.n175 585
R913 B.n327 B.n326 585
R914 B.n325 B.n176 585
R915 B.n324 B.n323 585
R916 B.n322 B.n177 585
R917 B.n321 B.n320 585
R918 B.n319 B.n178 585
R919 B.n318 B.n317 585
R920 B.n316 B.n179 585
R921 B.n419 B.n144 585
R922 B.n421 B.n420 585
R923 B.n422 B.n143 585
R924 B.n424 B.n423 585
R925 B.n425 B.n142 585
R926 B.n427 B.n426 585
R927 B.n428 B.n141 585
R928 B.n430 B.n429 585
R929 B.n431 B.n140 585
R930 B.n433 B.n432 585
R931 B.n434 B.n139 585
R932 B.n436 B.n435 585
R933 B.n437 B.n138 585
R934 B.n439 B.n438 585
R935 B.n440 B.n137 585
R936 B.n442 B.n441 585
R937 B.n443 B.n136 585
R938 B.n445 B.n444 585
R939 B.n446 B.n135 585
R940 B.n448 B.n447 585
R941 B.n449 B.n134 585
R942 B.n451 B.n450 585
R943 B.n452 B.n133 585
R944 B.n454 B.n453 585
R945 B.n455 B.n132 585
R946 B.n457 B.n456 585
R947 B.n458 B.n131 585
R948 B.n460 B.n459 585
R949 B.n461 B.n130 585
R950 B.n463 B.n462 585
R951 B.n464 B.n129 585
R952 B.n466 B.n465 585
R953 B.n467 B.n128 585
R954 B.n469 B.n468 585
R955 B.n470 B.n127 585
R956 B.n472 B.n471 585
R957 B.n473 B.n126 585
R958 B.n475 B.n474 585
R959 B.n476 B.n125 585
R960 B.n478 B.n477 585
R961 B.n479 B.n124 585
R962 B.n481 B.n480 585
R963 B.n482 B.n123 585
R964 B.n484 B.n483 585
R965 B.n485 B.n122 585
R966 B.n487 B.n486 585
R967 B.n488 B.n121 585
R968 B.n490 B.n489 585
R969 B.n491 B.n120 585
R970 B.n493 B.n492 585
R971 B.n494 B.n119 585
R972 B.n496 B.n495 585
R973 B.n497 B.n118 585
R974 B.n499 B.n498 585
R975 B.n500 B.n117 585
R976 B.n502 B.n501 585
R977 B.n503 B.n116 585
R978 B.n505 B.n504 585
R979 B.n506 B.n115 585
R980 B.n508 B.n507 585
R981 B.n509 B.n114 585
R982 B.n511 B.n510 585
R983 B.n512 B.n113 585
R984 B.n514 B.n513 585
R985 B.n515 B.n112 585
R986 B.n517 B.n516 585
R987 B.n518 B.n111 585
R988 B.n520 B.n519 585
R989 B.n521 B.n110 585
R990 B.n523 B.n522 585
R991 B.n524 B.n109 585
R992 B.n526 B.n525 585
R993 B.n527 B.n108 585
R994 B.n529 B.n528 585
R995 B.n530 B.n107 585
R996 B.n532 B.n531 585
R997 B.n533 B.n106 585
R998 B.n535 B.n534 585
R999 B.n536 B.n105 585
R1000 B.n538 B.n537 585
R1001 B.n539 B.n104 585
R1002 B.n541 B.n540 585
R1003 B.n542 B.n103 585
R1004 B.n544 B.n543 585
R1005 B.n545 B.n102 585
R1006 B.n547 B.n546 585
R1007 B.n548 B.n101 585
R1008 B.n550 B.n549 585
R1009 B.n551 B.n100 585
R1010 B.n553 B.n552 585
R1011 B.n554 B.n99 585
R1012 B.n556 B.n555 585
R1013 B.n557 B.n98 585
R1014 B.n559 B.n558 585
R1015 B.n560 B.n97 585
R1016 B.n562 B.n561 585
R1017 B.n563 B.n96 585
R1018 B.n565 B.n564 585
R1019 B.n566 B.n95 585
R1020 B.n568 B.n567 585
R1021 B.n569 B.n94 585
R1022 B.n571 B.n570 585
R1023 B.n572 B.n93 585
R1024 B.n574 B.n573 585
R1025 B.n575 B.n92 585
R1026 B.n577 B.n576 585
R1027 B.n578 B.n91 585
R1028 B.n580 B.n579 585
R1029 B.n581 B.n90 585
R1030 B.n583 B.n582 585
R1031 B.n584 B.n89 585
R1032 B.n586 B.n585 585
R1033 B.n587 B.n88 585
R1034 B.n589 B.n588 585
R1035 B.n590 B.n87 585
R1036 B.n592 B.n591 585
R1037 B.n593 B.n86 585
R1038 B.n595 B.n594 585
R1039 B.n596 B.n85 585
R1040 B.n598 B.n597 585
R1041 B.n599 B.n84 585
R1042 B.n601 B.n600 585
R1043 B.n602 B.n83 585
R1044 B.n604 B.n603 585
R1045 B.n605 B.n82 585
R1046 B.n607 B.n606 585
R1047 B.n608 B.n81 585
R1048 B.n610 B.n609 585
R1049 B.n611 B.n80 585
R1050 B.n613 B.n612 585
R1051 B.n614 B.n79 585
R1052 B.n616 B.n615 585
R1053 B.n617 B.n78 585
R1054 B.n619 B.n618 585
R1055 B.n620 B.n77 585
R1056 B.n622 B.n621 585
R1057 B.n623 B.n76 585
R1058 B.n625 B.n624 585
R1059 B.n626 B.n75 585
R1060 B.n628 B.n627 585
R1061 B.n728 B.n727 585
R1062 B.n726 B.n37 585
R1063 B.n725 B.n724 585
R1064 B.n723 B.n38 585
R1065 B.n722 B.n721 585
R1066 B.n720 B.n39 585
R1067 B.n719 B.n718 585
R1068 B.n717 B.n40 585
R1069 B.n716 B.n715 585
R1070 B.n714 B.n41 585
R1071 B.n713 B.n712 585
R1072 B.n711 B.n42 585
R1073 B.n710 B.n709 585
R1074 B.n708 B.n43 585
R1075 B.n707 B.n706 585
R1076 B.n705 B.n44 585
R1077 B.n704 B.n703 585
R1078 B.n702 B.n45 585
R1079 B.n701 B.n700 585
R1080 B.n699 B.n46 585
R1081 B.n698 B.n697 585
R1082 B.n696 B.n47 585
R1083 B.n695 B.n694 585
R1084 B.n693 B.n48 585
R1085 B.n692 B.n691 585
R1086 B.n690 B.n49 585
R1087 B.n689 B.n688 585
R1088 B.n687 B.n50 585
R1089 B.n686 B.n685 585
R1090 B.n684 B.n51 585
R1091 B.n683 B.n682 585
R1092 B.n681 B.n55 585
R1093 B.n680 B.n679 585
R1094 B.n678 B.n56 585
R1095 B.n677 B.n676 585
R1096 B.n675 B.n57 585
R1097 B.n674 B.n673 585
R1098 B.n672 B.n58 585
R1099 B.n670 B.n669 585
R1100 B.n668 B.n61 585
R1101 B.n667 B.n666 585
R1102 B.n665 B.n62 585
R1103 B.n664 B.n663 585
R1104 B.n662 B.n63 585
R1105 B.n661 B.n660 585
R1106 B.n659 B.n64 585
R1107 B.n658 B.n657 585
R1108 B.n656 B.n65 585
R1109 B.n655 B.n654 585
R1110 B.n653 B.n66 585
R1111 B.n652 B.n651 585
R1112 B.n650 B.n67 585
R1113 B.n649 B.n648 585
R1114 B.n647 B.n68 585
R1115 B.n646 B.n645 585
R1116 B.n644 B.n69 585
R1117 B.n643 B.n642 585
R1118 B.n641 B.n70 585
R1119 B.n640 B.n639 585
R1120 B.n638 B.n71 585
R1121 B.n637 B.n636 585
R1122 B.n635 B.n72 585
R1123 B.n634 B.n633 585
R1124 B.n632 B.n73 585
R1125 B.n631 B.n630 585
R1126 B.n629 B.n74 585
R1127 B.n729 B.n36 585
R1128 B.n731 B.n730 585
R1129 B.n732 B.n35 585
R1130 B.n734 B.n733 585
R1131 B.n735 B.n34 585
R1132 B.n737 B.n736 585
R1133 B.n738 B.n33 585
R1134 B.n740 B.n739 585
R1135 B.n741 B.n32 585
R1136 B.n743 B.n742 585
R1137 B.n744 B.n31 585
R1138 B.n746 B.n745 585
R1139 B.n747 B.n30 585
R1140 B.n749 B.n748 585
R1141 B.n750 B.n29 585
R1142 B.n752 B.n751 585
R1143 B.n753 B.n28 585
R1144 B.n755 B.n754 585
R1145 B.n756 B.n27 585
R1146 B.n758 B.n757 585
R1147 B.n759 B.n26 585
R1148 B.n761 B.n760 585
R1149 B.n762 B.n25 585
R1150 B.n764 B.n763 585
R1151 B.n765 B.n24 585
R1152 B.n767 B.n766 585
R1153 B.n768 B.n23 585
R1154 B.n770 B.n769 585
R1155 B.n771 B.n22 585
R1156 B.n773 B.n772 585
R1157 B.n774 B.n21 585
R1158 B.n776 B.n775 585
R1159 B.n777 B.n20 585
R1160 B.n779 B.n778 585
R1161 B.n780 B.n19 585
R1162 B.n782 B.n781 585
R1163 B.n783 B.n18 585
R1164 B.n785 B.n784 585
R1165 B.n786 B.n17 585
R1166 B.n788 B.n787 585
R1167 B.n789 B.n16 585
R1168 B.n791 B.n790 585
R1169 B.n792 B.n15 585
R1170 B.n794 B.n793 585
R1171 B.n795 B.n14 585
R1172 B.n797 B.n796 585
R1173 B.n798 B.n13 585
R1174 B.n800 B.n799 585
R1175 B.n801 B.n12 585
R1176 B.n803 B.n802 585
R1177 B.n804 B.n11 585
R1178 B.n806 B.n805 585
R1179 B.n807 B.n10 585
R1180 B.n809 B.n808 585
R1181 B.n810 B.n9 585
R1182 B.n812 B.n811 585
R1183 B.n813 B.n8 585
R1184 B.n815 B.n814 585
R1185 B.n816 B.n7 585
R1186 B.n818 B.n817 585
R1187 B.n819 B.n6 585
R1188 B.n821 B.n820 585
R1189 B.n822 B.n5 585
R1190 B.n824 B.n823 585
R1191 B.n825 B.n4 585
R1192 B.n827 B.n826 585
R1193 B.n828 B.n3 585
R1194 B.n830 B.n829 585
R1195 B.n831 B.n0 585
R1196 B.n2 B.n1 585
R1197 B.n214 B.n213 585
R1198 B.n216 B.n215 585
R1199 B.n217 B.n212 585
R1200 B.n219 B.n218 585
R1201 B.n220 B.n211 585
R1202 B.n222 B.n221 585
R1203 B.n223 B.n210 585
R1204 B.n225 B.n224 585
R1205 B.n226 B.n209 585
R1206 B.n228 B.n227 585
R1207 B.n229 B.n208 585
R1208 B.n231 B.n230 585
R1209 B.n232 B.n207 585
R1210 B.n234 B.n233 585
R1211 B.n235 B.n206 585
R1212 B.n237 B.n236 585
R1213 B.n238 B.n205 585
R1214 B.n240 B.n239 585
R1215 B.n241 B.n204 585
R1216 B.n243 B.n242 585
R1217 B.n244 B.n203 585
R1218 B.n246 B.n245 585
R1219 B.n247 B.n202 585
R1220 B.n249 B.n248 585
R1221 B.n250 B.n201 585
R1222 B.n252 B.n251 585
R1223 B.n253 B.n200 585
R1224 B.n255 B.n254 585
R1225 B.n256 B.n199 585
R1226 B.n258 B.n257 585
R1227 B.n259 B.n198 585
R1228 B.n261 B.n260 585
R1229 B.n262 B.n197 585
R1230 B.n264 B.n263 585
R1231 B.n265 B.n196 585
R1232 B.n267 B.n266 585
R1233 B.n268 B.n195 585
R1234 B.n270 B.n269 585
R1235 B.n271 B.n194 585
R1236 B.n273 B.n272 585
R1237 B.n274 B.n193 585
R1238 B.n276 B.n275 585
R1239 B.n277 B.n192 585
R1240 B.n279 B.n278 585
R1241 B.n280 B.n191 585
R1242 B.n282 B.n281 585
R1243 B.n283 B.n190 585
R1244 B.n285 B.n284 585
R1245 B.n286 B.n189 585
R1246 B.n288 B.n287 585
R1247 B.n289 B.n188 585
R1248 B.n291 B.n290 585
R1249 B.n292 B.n187 585
R1250 B.n294 B.n293 585
R1251 B.n295 B.n186 585
R1252 B.n297 B.n296 585
R1253 B.n298 B.n185 585
R1254 B.n300 B.n299 585
R1255 B.n301 B.n184 585
R1256 B.n303 B.n302 585
R1257 B.n304 B.n183 585
R1258 B.n306 B.n305 585
R1259 B.n307 B.n182 585
R1260 B.n309 B.n308 585
R1261 B.n310 B.n181 585
R1262 B.n312 B.n311 585
R1263 B.n313 B.n180 585
R1264 B.n315 B.n314 585
R1265 B.n316 B.n315 487.695
R1266 B.n417 B.n144 487.695
R1267 B.n627 B.n74 487.695
R1268 B.n729 B.n728 487.695
R1269 B.n159 B.t10 361.726
R1270 B.n59 B.t8 361.726
R1271 B.n356 B.t4 361.726
R1272 B.n52 B.t2 361.726
R1273 B.n160 B.t11 294.428
R1274 B.n60 B.t7 294.428
R1275 B.n357 B.t5 294.428
R1276 B.n53 B.t1 294.428
R1277 B.n356 B.t3 266.072
R1278 B.n159 B.t9 266.072
R1279 B.n59 B.t6 266.072
R1280 B.n52 B.t0 266.072
R1281 B.n833 B.n832 256.663
R1282 B.n832 B.n831 235.042
R1283 B.n832 B.n2 235.042
R1284 B.n317 B.n316 163.367
R1285 B.n317 B.n178 163.367
R1286 B.n321 B.n178 163.367
R1287 B.n322 B.n321 163.367
R1288 B.n323 B.n322 163.367
R1289 B.n323 B.n176 163.367
R1290 B.n327 B.n176 163.367
R1291 B.n328 B.n327 163.367
R1292 B.n329 B.n328 163.367
R1293 B.n329 B.n174 163.367
R1294 B.n333 B.n174 163.367
R1295 B.n334 B.n333 163.367
R1296 B.n335 B.n334 163.367
R1297 B.n335 B.n172 163.367
R1298 B.n339 B.n172 163.367
R1299 B.n340 B.n339 163.367
R1300 B.n341 B.n340 163.367
R1301 B.n341 B.n170 163.367
R1302 B.n345 B.n170 163.367
R1303 B.n346 B.n345 163.367
R1304 B.n347 B.n346 163.367
R1305 B.n347 B.n168 163.367
R1306 B.n351 B.n168 163.367
R1307 B.n352 B.n351 163.367
R1308 B.n353 B.n352 163.367
R1309 B.n353 B.n166 163.367
R1310 B.n360 B.n166 163.367
R1311 B.n361 B.n360 163.367
R1312 B.n362 B.n361 163.367
R1313 B.n362 B.n164 163.367
R1314 B.n366 B.n164 163.367
R1315 B.n367 B.n366 163.367
R1316 B.n368 B.n367 163.367
R1317 B.n368 B.n162 163.367
R1318 B.n372 B.n162 163.367
R1319 B.n373 B.n372 163.367
R1320 B.n374 B.n373 163.367
R1321 B.n374 B.n158 163.367
R1322 B.n379 B.n158 163.367
R1323 B.n380 B.n379 163.367
R1324 B.n381 B.n380 163.367
R1325 B.n381 B.n156 163.367
R1326 B.n385 B.n156 163.367
R1327 B.n386 B.n385 163.367
R1328 B.n387 B.n386 163.367
R1329 B.n387 B.n154 163.367
R1330 B.n391 B.n154 163.367
R1331 B.n392 B.n391 163.367
R1332 B.n393 B.n392 163.367
R1333 B.n393 B.n152 163.367
R1334 B.n397 B.n152 163.367
R1335 B.n398 B.n397 163.367
R1336 B.n399 B.n398 163.367
R1337 B.n399 B.n150 163.367
R1338 B.n403 B.n150 163.367
R1339 B.n404 B.n403 163.367
R1340 B.n405 B.n404 163.367
R1341 B.n405 B.n148 163.367
R1342 B.n409 B.n148 163.367
R1343 B.n410 B.n409 163.367
R1344 B.n411 B.n410 163.367
R1345 B.n411 B.n146 163.367
R1346 B.n415 B.n146 163.367
R1347 B.n416 B.n415 163.367
R1348 B.n417 B.n416 163.367
R1349 B.n627 B.n626 163.367
R1350 B.n626 B.n625 163.367
R1351 B.n625 B.n76 163.367
R1352 B.n621 B.n76 163.367
R1353 B.n621 B.n620 163.367
R1354 B.n620 B.n619 163.367
R1355 B.n619 B.n78 163.367
R1356 B.n615 B.n78 163.367
R1357 B.n615 B.n614 163.367
R1358 B.n614 B.n613 163.367
R1359 B.n613 B.n80 163.367
R1360 B.n609 B.n80 163.367
R1361 B.n609 B.n608 163.367
R1362 B.n608 B.n607 163.367
R1363 B.n607 B.n82 163.367
R1364 B.n603 B.n82 163.367
R1365 B.n603 B.n602 163.367
R1366 B.n602 B.n601 163.367
R1367 B.n601 B.n84 163.367
R1368 B.n597 B.n84 163.367
R1369 B.n597 B.n596 163.367
R1370 B.n596 B.n595 163.367
R1371 B.n595 B.n86 163.367
R1372 B.n591 B.n86 163.367
R1373 B.n591 B.n590 163.367
R1374 B.n590 B.n589 163.367
R1375 B.n589 B.n88 163.367
R1376 B.n585 B.n88 163.367
R1377 B.n585 B.n584 163.367
R1378 B.n584 B.n583 163.367
R1379 B.n583 B.n90 163.367
R1380 B.n579 B.n90 163.367
R1381 B.n579 B.n578 163.367
R1382 B.n578 B.n577 163.367
R1383 B.n577 B.n92 163.367
R1384 B.n573 B.n92 163.367
R1385 B.n573 B.n572 163.367
R1386 B.n572 B.n571 163.367
R1387 B.n571 B.n94 163.367
R1388 B.n567 B.n94 163.367
R1389 B.n567 B.n566 163.367
R1390 B.n566 B.n565 163.367
R1391 B.n565 B.n96 163.367
R1392 B.n561 B.n96 163.367
R1393 B.n561 B.n560 163.367
R1394 B.n560 B.n559 163.367
R1395 B.n559 B.n98 163.367
R1396 B.n555 B.n98 163.367
R1397 B.n555 B.n554 163.367
R1398 B.n554 B.n553 163.367
R1399 B.n553 B.n100 163.367
R1400 B.n549 B.n100 163.367
R1401 B.n549 B.n548 163.367
R1402 B.n548 B.n547 163.367
R1403 B.n547 B.n102 163.367
R1404 B.n543 B.n102 163.367
R1405 B.n543 B.n542 163.367
R1406 B.n542 B.n541 163.367
R1407 B.n541 B.n104 163.367
R1408 B.n537 B.n104 163.367
R1409 B.n537 B.n536 163.367
R1410 B.n536 B.n535 163.367
R1411 B.n535 B.n106 163.367
R1412 B.n531 B.n106 163.367
R1413 B.n531 B.n530 163.367
R1414 B.n530 B.n529 163.367
R1415 B.n529 B.n108 163.367
R1416 B.n525 B.n108 163.367
R1417 B.n525 B.n524 163.367
R1418 B.n524 B.n523 163.367
R1419 B.n523 B.n110 163.367
R1420 B.n519 B.n110 163.367
R1421 B.n519 B.n518 163.367
R1422 B.n518 B.n517 163.367
R1423 B.n517 B.n112 163.367
R1424 B.n513 B.n112 163.367
R1425 B.n513 B.n512 163.367
R1426 B.n512 B.n511 163.367
R1427 B.n511 B.n114 163.367
R1428 B.n507 B.n114 163.367
R1429 B.n507 B.n506 163.367
R1430 B.n506 B.n505 163.367
R1431 B.n505 B.n116 163.367
R1432 B.n501 B.n116 163.367
R1433 B.n501 B.n500 163.367
R1434 B.n500 B.n499 163.367
R1435 B.n499 B.n118 163.367
R1436 B.n495 B.n118 163.367
R1437 B.n495 B.n494 163.367
R1438 B.n494 B.n493 163.367
R1439 B.n493 B.n120 163.367
R1440 B.n489 B.n120 163.367
R1441 B.n489 B.n488 163.367
R1442 B.n488 B.n487 163.367
R1443 B.n487 B.n122 163.367
R1444 B.n483 B.n122 163.367
R1445 B.n483 B.n482 163.367
R1446 B.n482 B.n481 163.367
R1447 B.n481 B.n124 163.367
R1448 B.n477 B.n124 163.367
R1449 B.n477 B.n476 163.367
R1450 B.n476 B.n475 163.367
R1451 B.n475 B.n126 163.367
R1452 B.n471 B.n126 163.367
R1453 B.n471 B.n470 163.367
R1454 B.n470 B.n469 163.367
R1455 B.n469 B.n128 163.367
R1456 B.n465 B.n128 163.367
R1457 B.n465 B.n464 163.367
R1458 B.n464 B.n463 163.367
R1459 B.n463 B.n130 163.367
R1460 B.n459 B.n130 163.367
R1461 B.n459 B.n458 163.367
R1462 B.n458 B.n457 163.367
R1463 B.n457 B.n132 163.367
R1464 B.n453 B.n132 163.367
R1465 B.n453 B.n452 163.367
R1466 B.n452 B.n451 163.367
R1467 B.n451 B.n134 163.367
R1468 B.n447 B.n134 163.367
R1469 B.n447 B.n446 163.367
R1470 B.n446 B.n445 163.367
R1471 B.n445 B.n136 163.367
R1472 B.n441 B.n136 163.367
R1473 B.n441 B.n440 163.367
R1474 B.n440 B.n439 163.367
R1475 B.n439 B.n138 163.367
R1476 B.n435 B.n138 163.367
R1477 B.n435 B.n434 163.367
R1478 B.n434 B.n433 163.367
R1479 B.n433 B.n140 163.367
R1480 B.n429 B.n140 163.367
R1481 B.n429 B.n428 163.367
R1482 B.n428 B.n427 163.367
R1483 B.n427 B.n142 163.367
R1484 B.n423 B.n142 163.367
R1485 B.n423 B.n422 163.367
R1486 B.n422 B.n421 163.367
R1487 B.n421 B.n144 163.367
R1488 B.n728 B.n37 163.367
R1489 B.n724 B.n37 163.367
R1490 B.n724 B.n723 163.367
R1491 B.n723 B.n722 163.367
R1492 B.n722 B.n39 163.367
R1493 B.n718 B.n39 163.367
R1494 B.n718 B.n717 163.367
R1495 B.n717 B.n716 163.367
R1496 B.n716 B.n41 163.367
R1497 B.n712 B.n41 163.367
R1498 B.n712 B.n711 163.367
R1499 B.n711 B.n710 163.367
R1500 B.n710 B.n43 163.367
R1501 B.n706 B.n43 163.367
R1502 B.n706 B.n705 163.367
R1503 B.n705 B.n704 163.367
R1504 B.n704 B.n45 163.367
R1505 B.n700 B.n45 163.367
R1506 B.n700 B.n699 163.367
R1507 B.n699 B.n698 163.367
R1508 B.n698 B.n47 163.367
R1509 B.n694 B.n47 163.367
R1510 B.n694 B.n693 163.367
R1511 B.n693 B.n692 163.367
R1512 B.n692 B.n49 163.367
R1513 B.n688 B.n49 163.367
R1514 B.n688 B.n687 163.367
R1515 B.n687 B.n686 163.367
R1516 B.n686 B.n51 163.367
R1517 B.n682 B.n51 163.367
R1518 B.n682 B.n681 163.367
R1519 B.n681 B.n680 163.367
R1520 B.n680 B.n56 163.367
R1521 B.n676 B.n56 163.367
R1522 B.n676 B.n675 163.367
R1523 B.n675 B.n674 163.367
R1524 B.n674 B.n58 163.367
R1525 B.n669 B.n58 163.367
R1526 B.n669 B.n668 163.367
R1527 B.n668 B.n667 163.367
R1528 B.n667 B.n62 163.367
R1529 B.n663 B.n62 163.367
R1530 B.n663 B.n662 163.367
R1531 B.n662 B.n661 163.367
R1532 B.n661 B.n64 163.367
R1533 B.n657 B.n64 163.367
R1534 B.n657 B.n656 163.367
R1535 B.n656 B.n655 163.367
R1536 B.n655 B.n66 163.367
R1537 B.n651 B.n66 163.367
R1538 B.n651 B.n650 163.367
R1539 B.n650 B.n649 163.367
R1540 B.n649 B.n68 163.367
R1541 B.n645 B.n68 163.367
R1542 B.n645 B.n644 163.367
R1543 B.n644 B.n643 163.367
R1544 B.n643 B.n70 163.367
R1545 B.n639 B.n70 163.367
R1546 B.n639 B.n638 163.367
R1547 B.n638 B.n637 163.367
R1548 B.n637 B.n72 163.367
R1549 B.n633 B.n72 163.367
R1550 B.n633 B.n632 163.367
R1551 B.n632 B.n631 163.367
R1552 B.n631 B.n74 163.367
R1553 B.n730 B.n729 163.367
R1554 B.n730 B.n35 163.367
R1555 B.n734 B.n35 163.367
R1556 B.n735 B.n734 163.367
R1557 B.n736 B.n735 163.367
R1558 B.n736 B.n33 163.367
R1559 B.n740 B.n33 163.367
R1560 B.n741 B.n740 163.367
R1561 B.n742 B.n741 163.367
R1562 B.n742 B.n31 163.367
R1563 B.n746 B.n31 163.367
R1564 B.n747 B.n746 163.367
R1565 B.n748 B.n747 163.367
R1566 B.n748 B.n29 163.367
R1567 B.n752 B.n29 163.367
R1568 B.n753 B.n752 163.367
R1569 B.n754 B.n753 163.367
R1570 B.n754 B.n27 163.367
R1571 B.n758 B.n27 163.367
R1572 B.n759 B.n758 163.367
R1573 B.n760 B.n759 163.367
R1574 B.n760 B.n25 163.367
R1575 B.n764 B.n25 163.367
R1576 B.n765 B.n764 163.367
R1577 B.n766 B.n765 163.367
R1578 B.n766 B.n23 163.367
R1579 B.n770 B.n23 163.367
R1580 B.n771 B.n770 163.367
R1581 B.n772 B.n771 163.367
R1582 B.n772 B.n21 163.367
R1583 B.n776 B.n21 163.367
R1584 B.n777 B.n776 163.367
R1585 B.n778 B.n777 163.367
R1586 B.n778 B.n19 163.367
R1587 B.n782 B.n19 163.367
R1588 B.n783 B.n782 163.367
R1589 B.n784 B.n783 163.367
R1590 B.n784 B.n17 163.367
R1591 B.n788 B.n17 163.367
R1592 B.n789 B.n788 163.367
R1593 B.n790 B.n789 163.367
R1594 B.n790 B.n15 163.367
R1595 B.n794 B.n15 163.367
R1596 B.n795 B.n794 163.367
R1597 B.n796 B.n795 163.367
R1598 B.n796 B.n13 163.367
R1599 B.n800 B.n13 163.367
R1600 B.n801 B.n800 163.367
R1601 B.n802 B.n801 163.367
R1602 B.n802 B.n11 163.367
R1603 B.n806 B.n11 163.367
R1604 B.n807 B.n806 163.367
R1605 B.n808 B.n807 163.367
R1606 B.n808 B.n9 163.367
R1607 B.n812 B.n9 163.367
R1608 B.n813 B.n812 163.367
R1609 B.n814 B.n813 163.367
R1610 B.n814 B.n7 163.367
R1611 B.n818 B.n7 163.367
R1612 B.n819 B.n818 163.367
R1613 B.n820 B.n819 163.367
R1614 B.n820 B.n5 163.367
R1615 B.n824 B.n5 163.367
R1616 B.n825 B.n824 163.367
R1617 B.n826 B.n825 163.367
R1618 B.n826 B.n3 163.367
R1619 B.n830 B.n3 163.367
R1620 B.n831 B.n830 163.367
R1621 B.n214 B.n2 163.367
R1622 B.n215 B.n214 163.367
R1623 B.n215 B.n212 163.367
R1624 B.n219 B.n212 163.367
R1625 B.n220 B.n219 163.367
R1626 B.n221 B.n220 163.367
R1627 B.n221 B.n210 163.367
R1628 B.n225 B.n210 163.367
R1629 B.n226 B.n225 163.367
R1630 B.n227 B.n226 163.367
R1631 B.n227 B.n208 163.367
R1632 B.n231 B.n208 163.367
R1633 B.n232 B.n231 163.367
R1634 B.n233 B.n232 163.367
R1635 B.n233 B.n206 163.367
R1636 B.n237 B.n206 163.367
R1637 B.n238 B.n237 163.367
R1638 B.n239 B.n238 163.367
R1639 B.n239 B.n204 163.367
R1640 B.n243 B.n204 163.367
R1641 B.n244 B.n243 163.367
R1642 B.n245 B.n244 163.367
R1643 B.n245 B.n202 163.367
R1644 B.n249 B.n202 163.367
R1645 B.n250 B.n249 163.367
R1646 B.n251 B.n250 163.367
R1647 B.n251 B.n200 163.367
R1648 B.n255 B.n200 163.367
R1649 B.n256 B.n255 163.367
R1650 B.n257 B.n256 163.367
R1651 B.n257 B.n198 163.367
R1652 B.n261 B.n198 163.367
R1653 B.n262 B.n261 163.367
R1654 B.n263 B.n262 163.367
R1655 B.n263 B.n196 163.367
R1656 B.n267 B.n196 163.367
R1657 B.n268 B.n267 163.367
R1658 B.n269 B.n268 163.367
R1659 B.n269 B.n194 163.367
R1660 B.n273 B.n194 163.367
R1661 B.n274 B.n273 163.367
R1662 B.n275 B.n274 163.367
R1663 B.n275 B.n192 163.367
R1664 B.n279 B.n192 163.367
R1665 B.n280 B.n279 163.367
R1666 B.n281 B.n280 163.367
R1667 B.n281 B.n190 163.367
R1668 B.n285 B.n190 163.367
R1669 B.n286 B.n285 163.367
R1670 B.n287 B.n286 163.367
R1671 B.n287 B.n188 163.367
R1672 B.n291 B.n188 163.367
R1673 B.n292 B.n291 163.367
R1674 B.n293 B.n292 163.367
R1675 B.n293 B.n186 163.367
R1676 B.n297 B.n186 163.367
R1677 B.n298 B.n297 163.367
R1678 B.n299 B.n298 163.367
R1679 B.n299 B.n184 163.367
R1680 B.n303 B.n184 163.367
R1681 B.n304 B.n303 163.367
R1682 B.n305 B.n304 163.367
R1683 B.n305 B.n182 163.367
R1684 B.n309 B.n182 163.367
R1685 B.n310 B.n309 163.367
R1686 B.n311 B.n310 163.367
R1687 B.n311 B.n180 163.367
R1688 B.n315 B.n180 163.367
R1689 B.n357 B.n356 67.2975
R1690 B.n160 B.n159 67.2975
R1691 B.n60 B.n59 67.2975
R1692 B.n53 B.n52 67.2975
R1693 B.n358 B.n357 59.5399
R1694 B.n376 B.n160 59.5399
R1695 B.n671 B.n60 59.5399
R1696 B.n54 B.n53 59.5399
R1697 B.n727 B.n36 31.6883
R1698 B.n629 B.n628 31.6883
R1699 B.n419 B.n418 31.6883
R1700 B.n314 B.n179 31.6883
R1701 B B.n833 18.0485
R1702 B.n731 B.n36 10.6151
R1703 B.n732 B.n731 10.6151
R1704 B.n733 B.n732 10.6151
R1705 B.n733 B.n34 10.6151
R1706 B.n737 B.n34 10.6151
R1707 B.n738 B.n737 10.6151
R1708 B.n739 B.n738 10.6151
R1709 B.n739 B.n32 10.6151
R1710 B.n743 B.n32 10.6151
R1711 B.n744 B.n743 10.6151
R1712 B.n745 B.n744 10.6151
R1713 B.n745 B.n30 10.6151
R1714 B.n749 B.n30 10.6151
R1715 B.n750 B.n749 10.6151
R1716 B.n751 B.n750 10.6151
R1717 B.n751 B.n28 10.6151
R1718 B.n755 B.n28 10.6151
R1719 B.n756 B.n755 10.6151
R1720 B.n757 B.n756 10.6151
R1721 B.n757 B.n26 10.6151
R1722 B.n761 B.n26 10.6151
R1723 B.n762 B.n761 10.6151
R1724 B.n763 B.n762 10.6151
R1725 B.n763 B.n24 10.6151
R1726 B.n767 B.n24 10.6151
R1727 B.n768 B.n767 10.6151
R1728 B.n769 B.n768 10.6151
R1729 B.n769 B.n22 10.6151
R1730 B.n773 B.n22 10.6151
R1731 B.n774 B.n773 10.6151
R1732 B.n775 B.n774 10.6151
R1733 B.n775 B.n20 10.6151
R1734 B.n779 B.n20 10.6151
R1735 B.n780 B.n779 10.6151
R1736 B.n781 B.n780 10.6151
R1737 B.n781 B.n18 10.6151
R1738 B.n785 B.n18 10.6151
R1739 B.n786 B.n785 10.6151
R1740 B.n787 B.n786 10.6151
R1741 B.n787 B.n16 10.6151
R1742 B.n791 B.n16 10.6151
R1743 B.n792 B.n791 10.6151
R1744 B.n793 B.n792 10.6151
R1745 B.n793 B.n14 10.6151
R1746 B.n797 B.n14 10.6151
R1747 B.n798 B.n797 10.6151
R1748 B.n799 B.n798 10.6151
R1749 B.n799 B.n12 10.6151
R1750 B.n803 B.n12 10.6151
R1751 B.n804 B.n803 10.6151
R1752 B.n805 B.n804 10.6151
R1753 B.n805 B.n10 10.6151
R1754 B.n809 B.n10 10.6151
R1755 B.n810 B.n809 10.6151
R1756 B.n811 B.n810 10.6151
R1757 B.n811 B.n8 10.6151
R1758 B.n815 B.n8 10.6151
R1759 B.n816 B.n815 10.6151
R1760 B.n817 B.n816 10.6151
R1761 B.n817 B.n6 10.6151
R1762 B.n821 B.n6 10.6151
R1763 B.n822 B.n821 10.6151
R1764 B.n823 B.n822 10.6151
R1765 B.n823 B.n4 10.6151
R1766 B.n827 B.n4 10.6151
R1767 B.n828 B.n827 10.6151
R1768 B.n829 B.n828 10.6151
R1769 B.n829 B.n0 10.6151
R1770 B.n727 B.n726 10.6151
R1771 B.n726 B.n725 10.6151
R1772 B.n725 B.n38 10.6151
R1773 B.n721 B.n38 10.6151
R1774 B.n721 B.n720 10.6151
R1775 B.n720 B.n719 10.6151
R1776 B.n719 B.n40 10.6151
R1777 B.n715 B.n40 10.6151
R1778 B.n715 B.n714 10.6151
R1779 B.n714 B.n713 10.6151
R1780 B.n713 B.n42 10.6151
R1781 B.n709 B.n42 10.6151
R1782 B.n709 B.n708 10.6151
R1783 B.n708 B.n707 10.6151
R1784 B.n707 B.n44 10.6151
R1785 B.n703 B.n44 10.6151
R1786 B.n703 B.n702 10.6151
R1787 B.n702 B.n701 10.6151
R1788 B.n701 B.n46 10.6151
R1789 B.n697 B.n46 10.6151
R1790 B.n697 B.n696 10.6151
R1791 B.n696 B.n695 10.6151
R1792 B.n695 B.n48 10.6151
R1793 B.n691 B.n48 10.6151
R1794 B.n691 B.n690 10.6151
R1795 B.n690 B.n689 10.6151
R1796 B.n689 B.n50 10.6151
R1797 B.n685 B.n684 10.6151
R1798 B.n684 B.n683 10.6151
R1799 B.n683 B.n55 10.6151
R1800 B.n679 B.n55 10.6151
R1801 B.n679 B.n678 10.6151
R1802 B.n678 B.n677 10.6151
R1803 B.n677 B.n57 10.6151
R1804 B.n673 B.n57 10.6151
R1805 B.n673 B.n672 10.6151
R1806 B.n670 B.n61 10.6151
R1807 B.n666 B.n61 10.6151
R1808 B.n666 B.n665 10.6151
R1809 B.n665 B.n664 10.6151
R1810 B.n664 B.n63 10.6151
R1811 B.n660 B.n63 10.6151
R1812 B.n660 B.n659 10.6151
R1813 B.n659 B.n658 10.6151
R1814 B.n658 B.n65 10.6151
R1815 B.n654 B.n65 10.6151
R1816 B.n654 B.n653 10.6151
R1817 B.n653 B.n652 10.6151
R1818 B.n652 B.n67 10.6151
R1819 B.n648 B.n67 10.6151
R1820 B.n648 B.n647 10.6151
R1821 B.n647 B.n646 10.6151
R1822 B.n646 B.n69 10.6151
R1823 B.n642 B.n69 10.6151
R1824 B.n642 B.n641 10.6151
R1825 B.n641 B.n640 10.6151
R1826 B.n640 B.n71 10.6151
R1827 B.n636 B.n71 10.6151
R1828 B.n636 B.n635 10.6151
R1829 B.n635 B.n634 10.6151
R1830 B.n634 B.n73 10.6151
R1831 B.n630 B.n73 10.6151
R1832 B.n630 B.n629 10.6151
R1833 B.n628 B.n75 10.6151
R1834 B.n624 B.n75 10.6151
R1835 B.n624 B.n623 10.6151
R1836 B.n623 B.n622 10.6151
R1837 B.n622 B.n77 10.6151
R1838 B.n618 B.n77 10.6151
R1839 B.n618 B.n617 10.6151
R1840 B.n617 B.n616 10.6151
R1841 B.n616 B.n79 10.6151
R1842 B.n612 B.n79 10.6151
R1843 B.n612 B.n611 10.6151
R1844 B.n611 B.n610 10.6151
R1845 B.n610 B.n81 10.6151
R1846 B.n606 B.n81 10.6151
R1847 B.n606 B.n605 10.6151
R1848 B.n605 B.n604 10.6151
R1849 B.n604 B.n83 10.6151
R1850 B.n600 B.n83 10.6151
R1851 B.n600 B.n599 10.6151
R1852 B.n599 B.n598 10.6151
R1853 B.n598 B.n85 10.6151
R1854 B.n594 B.n85 10.6151
R1855 B.n594 B.n593 10.6151
R1856 B.n593 B.n592 10.6151
R1857 B.n592 B.n87 10.6151
R1858 B.n588 B.n87 10.6151
R1859 B.n588 B.n587 10.6151
R1860 B.n587 B.n586 10.6151
R1861 B.n586 B.n89 10.6151
R1862 B.n582 B.n89 10.6151
R1863 B.n582 B.n581 10.6151
R1864 B.n581 B.n580 10.6151
R1865 B.n580 B.n91 10.6151
R1866 B.n576 B.n91 10.6151
R1867 B.n576 B.n575 10.6151
R1868 B.n575 B.n574 10.6151
R1869 B.n574 B.n93 10.6151
R1870 B.n570 B.n93 10.6151
R1871 B.n570 B.n569 10.6151
R1872 B.n569 B.n568 10.6151
R1873 B.n568 B.n95 10.6151
R1874 B.n564 B.n95 10.6151
R1875 B.n564 B.n563 10.6151
R1876 B.n563 B.n562 10.6151
R1877 B.n562 B.n97 10.6151
R1878 B.n558 B.n97 10.6151
R1879 B.n558 B.n557 10.6151
R1880 B.n557 B.n556 10.6151
R1881 B.n556 B.n99 10.6151
R1882 B.n552 B.n99 10.6151
R1883 B.n552 B.n551 10.6151
R1884 B.n551 B.n550 10.6151
R1885 B.n550 B.n101 10.6151
R1886 B.n546 B.n101 10.6151
R1887 B.n546 B.n545 10.6151
R1888 B.n545 B.n544 10.6151
R1889 B.n544 B.n103 10.6151
R1890 B.n540 B.n103 10.6151
R1891 B.n540 B.n539 10.6151
R1892 B.n539 B.n538 10.6151
R1893 B.n538 B.n105 10.6151
R1894 B.n534 B.n105 10.6151
R1895 B.n534 B.n533 10.6151
R1896 B.n533 B.n532 10.6151
R1897 B.n532 B.n107 10.6151
R1898 B.n528 B.n107 10.6151
R1899 B.n528 B.n527 10.6151
R1900 B.n527 B.n526 10.6151
R1901 B.n526 B.n109 10.6151
R1902 B.n522 B.n109 10.6151
R1903 B.n522 B.n521 10.6151
R1904 B.n521 B.n520 10.6151
R1905 B.n520 B.n111 10.6151
R1906 B.n516 B.n111 10.6151
R1907 B.n516 B.n515 10.6151
R1908 B.n515 B.n514 10.6151
R1909 B.n514 B.n113 10.6151
R1910 B.n510 B.n113 10.6151
R1911 B.n510 B.n509 10.6151
R1912 B.n509 B.n508 10.6151
R1913 B.n508 B.n115 10.6151
R1914 B.n504 B.n115 10.6151
R1915 B.n504 B.n503 10.6151
R1916 B.n503 B.n502 10.6151
R1917 B.n502 B.n117 10.6151
R1918 B.n498 B.n117 10.6151
R1919 B.n498 B.n497 10.6151
R1920 B.n497 B.n496 10.6151
R1921 B.n496 B.n119 10.6151
R1922 B.n492 B.n119 10.6151
R1923 B.n492 B.n491 10.6151
R1924 B.n491 B.n490 10.6151
R1925 B.n490 B.n121 10.6151
R1926 B.n486 B.n121 10.6151
R1927 B.n486 B.n485 10.6151
R1928 B.n485 B.n484 10.6151
R1929 B.n484 B.n123 10.6151
R1930 B.n480 B.n123 10.6151
R1931 B.n480 B.n479 10.6151
R1932 B.n479 B.n478 10.6151
R1933 B.n478 B.n125 10.6151
R1934 B.n474 B.n125 10.6151
R1935 B.n474 B.n473 10.6151
R1936 B.n473 B.n472 10.6151
R1937 B.n472 B.n127 10.6151
R1938 B.n468 B.n127 10.6151
R1939 B.n468 B.n467 10.6151
R1940 B.n467 B.n466 10.6151
R1941 B.n466 B.n129 10.6151
R1942 B.n462 B.n129 10.6151
R1943 B.n462 B.n461 10.6151
R1944 B.n461 B.n460 10.6151
R1945 B.n460 B.n131 10.6151
R1946 B.n456 B.n131 10.6151
R1947 B.n456 B.n455 10.6151
R1948 B.n455 B.n454 10.6151
R1949 B.n454 B.n133 10.6151
R1950 B.n450 B.n133 10.6151
R1951 B.n450 B.n449 10.6151
R1952 B.n449 B.n448 10.6151
R1953 B.n448 B.n135 10.6151
R1954 B.n444 B.n135 10.6151
R1955 B.n444 B.n443 10.6151
R1956 B.n443 B.n442 10.6151
R1957 B.n442 B.n137 10.6151
R1958 B.n438 B.n137 10.6151
R1959 B.n438 B.n437 10.6151
R1960 B.n437 B.n436 10.6151
R1961 B.n436 B.n139 10.6151
R1962 B.n432 B.n139 10.6151
R1963 B.n432 B.n431 10.6151
R1964 B.n431 B.n430 10.6151
R1965 B.n430 B.n141 10.6151
R1966 B.n426 B.n141 10.6151
R1967 B.n426 B.n425 10.6151
R1968 B.n425 B.n424 10.6151
R1969 B.n424 B.n143 10.6151
R1970 B.n420 B.n143 10.6151
R1971 B.n420 B.n419 10.6151
R1972 B.n213 B.n1 10.6151
R1973 B.n216 B.n213 10.6151
R1974 B.n217 B.n216 10.6151
R1975 B.n218 B.n217 10.6151
R1976 B.n218 B.n211 10.6151
R1977 B.n222 B.n211 10.6151
R1978 B.n223 B.n222 10.6151
R1979 B.n224 B.n223 10.6151
R1980 B.n224 B.n209 10.6151
R1981 B.n228 B.n209 10.6151
R1982 B.n229 B.n228 10.6151
R1983 B.n230 B.n229 10.6151
R1984 B.n230 B.n207 10.6151
R1985 B.n234 B.n207 10.6151
R1986 B.n235 B.n234 10.6151
R1987 B.n236 B.n235 10.6151
R1988 B.n236 B.n205 10.6151
R1989 B.n240 B.n205 10.6151
R1990 B.n241 B.n240 10.6151
R1991 B.n242 B.n241 10.6151
R1992 B.n242 B.n203 10.6151
R1993 B.n246 B.n203 10.6151
R1994 B.n247 B.n246 10.6151
R1995 B.n248 B.n247 10.6151
R1996 B.n248 B.n201 10.6151
R1997 B.n252 B.n201 10.6151
R1998 B.n253 B.n252 10.6151
R1999 B.n254 B.n253 10.6151
R2000 B.n254 B.n199 10.6151
R2001 B.n258 B.n199 10.6151
R2002 B.n259 B.n258 10.6151
R2003 B.n260 B.n259 10.6151
R2004 B.n260 B.n197 10.6151
R2005 B.n264 B.n197 10.6151
R2006 B.n265 B.n264 10.6151
R2007 B.n266 B.n265 10.6151
R2008 B.n266 B.n195 10.6151
R2009 B.n270 B.n195 10.6151
R2010 B.n271 B.n270 10.6151
R2011 B.n272 B.n271 10.6151
R2012 B.n272 B.n193 10.6151
R2013 B.n276 B.n193 10.6151
R2014 B.n277 B.n276 10.6151
R2015 B.n278 B.n277 10.6151
R2016 B.n278 B.n191 10.6151
R2017 B.n282 B.n191 10.6151
R2018 B.n283 B.n282 10.6151
R2019 B.n284 B.n283 10.6151
R2020 B.n284 B.n189 10.6151
R2021 B.n288 B.n189 10.6151
R2022 B.n289 B.n288 10.6151
R2023 B.n290 B.n289 10.6151
R2024 B.n290 B.n187 10.6151
R2025 B.n294 B.n187 10.6151
R2026 B.n295 B.n294 10.6151
R2027 B.n296 B.n295 10.6151
R2028 B.n296 B.n185 10.6151
R2029 B.n300 B.n185 10.6151
R2030 B.n301 B.n300 10.6151
R2031 B.n302 B.n301 10.6151
R2032 B.n302 B.n183 10.6151
R2033 B.n306 B.n183 10.6151
R2034 B.n307 B.n306 10.6151
R2035 B.n308 B.n307 10.6151
R2036 B.n308 B.n181 10.6151
R2037 B.n312 B.n181 10.6151
R2038 B.n313 B.n312 10.6151
R2039 B.n314 B.n313 10.6151
R2040 B.n318 B.n179 10.6151
R2041 B.n319 B.n318 10.6151
R2042 B.n320 B.n319 10.6151
R2043 B.n320 B.n177 10.6151
R2044 B.n324 B.n177 10.6151
R2045 B.n325 B.n324 10.6151
R2046 B.n326 B.n325 10.6151
R2047 B.n326 B.n175 10.6151
R2048 B.n330 B.n175 10.6151
R2049 B.n331 B.n330 10.6151
R2050 B.n332 B.n331 10.6151
R2051 B.n332 B.n173 10.6151
R2052 B.n336 B.n173 10.6151
R2053 B.n337 B.n336 10.6151
R2054 B.n338 B.n337 10.6151
R2055 B.n338 B.n171 10.6151
R2056 B.n342 B.n171 10.6151
R2057 B.n343 B.n342 10.6151
R2058 B.n344 B.n343 10.6151
R2059 B.n344 B.n169 10.6151
R2060 B.n348 B.n169 10.6151
R2061 B.n349 B.n348 10.6151
R2062 B.n350 B.n349 10.6151
R2063 B.n350 B.n167 10.6151
R2064 B.n354 B.n167 10.6151
R2065 B.n355 B.n354 10.6151
R2066 B.n359 B.n355 10.6151
R2067 B.n363 B.n165 10.6151
R2068 B.n364 B.n363 10.6151
R2069 B.n365 B.n364 10.6151
R2070 B.n365 B.n163 10.6151
R2071 B.n369 B.n163 10.6151
R2072 B.n370 B.n369 10.6151
R2073 B.n371 B.n370 10.6151
R2074 B.n371 B.n161 10.6151
R2075 B.n375 B.n161 10.6151
R2076 B.n378 B.n377 10.6151
R2077 B.n378 B.n157 10.6151
R2078 B.n382 B.n157 10.6151
R2079 B.n383 B.n382 10.6151
R2080 B.n384 B.n383 10.6151
R2081 B.n384 B.n155 10.6151
R2082 B.n388 B.n155 10.6151
R2083 B.n389 B.n388 10.6151
R2084 B.n390 B.n389 10.6151
R2085 B.n390 B.n153 10.6151
R2086 B.n394 B.n153 10.6151
R2087 B.n395 B.n394 10.6151
R2088 B.n396 B.n395 10.6151
R2089 B.n396 B.n151 10.6151
R2090 B.n400 B.n151 10.6151
R2091 B.n401 B.n400 10.6151
R2092 B.n402 B.n401 10.6151
R2093 B.n402 B.n149 10.6151
R2094 B.n406 B.n149 10.6151
R2095 B.n407 B.n406 10.6151
R2096 B.n408 B.n407 10.6151
R2097 B.n408 B.n147 10.6151
R2098 B.n412 B.n147 10.6151
R2099 B.n413 B.n412 10.6151
R2100 B.n414 B.n413 10.6151
R2101 B.n414 B.n145 10.6151
R2102 B.n418 B.n145 10.6151
R2103 B.n54 B.n50 9.36635
R2104 B.n671 B.n670 9.36635
R2105 B.n359 B.n358 9.36635
R2106 B.n377 B.n376 9.36635
R2107 B.n833 B.n0 8.11757
R2108 B.n833 B.n1 8.11757
R2109 B.n685 B.n54 1.24928
R2110 B.n672 B.n671 1.24928
R2111 B.n358 B.n165 1.24928
R2112 B.n376 B.n375 1.24928
C0 VDD2 VP 0.652329f
C1 B VTAIL 2.89551f
C2 VTAIL VDD1 8.683081f
C3 VN VTAIL 8.15266f
C4 B VDD1 2.32908f
C5 B VN 1.36748f
C6 VN VDD1 0.154763f
C7 w_n5134_n2462# VTAIL 2.67221f
C8 VTAIL VP 8.16686f
C9 w_n5134_n2462# B 10.1852f
C10 w_n5134_n2462# VDD1 2.68522f
C11 w_n5134_n2462# VN 11.051499f
C12 VDD2 VTAIL 8.739019f
C13 B VP 2.49725f
C14 VDD1 VP 7.56371f
C15 VN VP 8.35467f
C16 VDD2 B 2.46802f
C17 VDD2 VDD1 2.52685f
C18 VDD2 VN 7.06935f
C19 w_n5134_n2462# VP 11.7216f
C20 w_n5134_n2462# VDD2 2.85683f
C21 VDD2 VSUBS 2.324104f
C22 VDD1 VSUBS 2.079118f
C23 VTAIL VSUBS 1.294289f
C24 VN VSUBS 8.564559f
C25 VP VSUBS 4.782906f
C26 B VSUBS 5.655603f
C27 w_n5134_n2462# VSUBS 0.157039p
C28 B.n0 VSUBS 0.009549f
C29 B.n1 VSUBS 0.009549f
C30 B.n2 VSUBS 0.014122f
C31 B.n3 VSUBS 0.010822f
C32 B.n4 VSUBS 0.010822f
C33 B.n5 VSUBS 0.010822f
C34 B.n6 VSUBS 0.010822f
C35 B.n7 VSUBS 0.010822f
C36 B.n8 VSUBS 0.010822f
C37 B.n9 VSUBS 0.010822f
C38 B.n10 VSUBS 0.010822f
C39 B.n11 VSUBS 0.010822f
C40 B.n12 VSUBS 0.010822f
C41 B.n13 VSUBS 0.010822f
C42 B.n14 VSUBS 0.010822f
C43 B.n15 VSUBS 0.010822f
C44 B.n16 VSUBS 0.010822f
C45 B.n17 VSUBS 0.010822f
C46 B.n18 VSUBS 0.010822f
C47 B.n19 VSUBS 0.010822f
C48 B.n20 VSUBS 0.010822f
C49 B.n21 VSUBS 0.010822f
C50 B.n22 VSUBS 0.010822f
C51 B.n23 VSUBS 0.010822f
C52 B.n24 VSUBS 0.010822f
C53 B.n25 VSUBS 0.010822f
C54 B.n26 VSUBS 0.010822f
C55 B.n27 VSUBS 0.010822f
C56 B.n28 VSUBS 0.010822f
C57 B.n29 VSUBS 0.010822f
C58 B.n30 VSUBS 0.010822f
C59 B.n31 VSUBS 0.010822f
C60 B.n32 VSUBS 0.010822f
C61 B.n33 VSUBS 0.010822f
C62 B.n34 VSUBS 0.010822f
C63 B.n35 VSUBS 0.010822f
C64 B.n36 VSUBS 0.024458f
C65 B.n37 VSUBS 0.010822f
C66 B.n38 VSUBS 0.010822f
C67 B.n39 VSUBS 0.010822f
C68 B.n40 VSUBS 0.010822f
C69 B.n41 VSUBS 0.010822f
C70 B.n42 VSUBS 0.010822f
C71 B.n43 VSUBS 0.010822f
C72 B.n44 VSUBS 0.010822f
C73 B.n45 VSUBS 0.010822f
C74 B.n46 VSUBS 0.010822f
C75 B.n47 VSUBS 0.010822f
C76 B.n48 VSUBS 0.010822f
C77 B.n49 VSUBS 0.010822f
C78 B.n50 VSUBS 0.010185f
C79 B.n51 VSUBS 0.010822f
C80 B.t1 VSUBS 0.180326f
C81 B.t2 VSUBS 0.230572f
C82 B.t0 VSUBS 1.71365f
C83 B.n52 VSUBS 0.380046f
C84 B.n53 VSUBS 0.285511f
C85 B.n54 VSUBS 0.025074f
C86 B.n55 VSUBS 0.010822f
C87 B.n56 VSUBS 0.010822f
C88 B.n57 VSUBS 0.010822f
C89 B.n58 VSUBS 0.010822f
C90 B.t7 VSUBS 0.18033f
C91 B.t8 VSUBS 0.230575f
C92 B.t6 VSUBS 1.71365f
C93 B.n59 VSUBS 0.380043f
C94 B.n60 VSUBS 0.285508f
C95 B.n61 VSUBS 0.010822f
C96 B.n62 VSUBS 0.010822f
C97 B.n63 VSUBS 0.010822f
C98 B.n64 VSUBS 0.010822f
C99 B.n65 VSUBS 0.010822f
C100 B.n66 VSUBS 0.010822f
C101 B.n67 VSUBS 0.010822f
C102 B.n68 VSUBS 0.010822f
C103 B.n69 VSUBS 0.010822f
C104 B.n70 VSUBS 0.010822f
C105 B.n71 VSUBS 0.010822f
C106 B.n72 VSUBS 0.010822f
C107 B.n73 VSUBS 0.010822f
C108 B.n74 VSUBS 0.025197f
C109 B.n75 VSUBS 0.010822f
C110 B.n76 VSUBS 0.010822f
C111 B.n77 VSUBS 0.010822f
C112 B.n78 VSUBS 0.010822f
C113 B.n79 VSUBS 0.010822f
C114 B.n80 VSUBS 0.010822f
C115 B.n81 VSUBS 0.010822f
C116 B.n82 VSUBS 0.010822f
C117 B.n83 VSUBS 0.010822f
C118 B.n84 VSUBS 0.010822f
C119 B.n85 VSUBS 0.010822f
C120 B.n86 VSUBS 0.010822f
C121 B.n87 VSUBS 0.010822f
C122 B.n88 VSUBS 0.010822f
C123 B.n89 VSUBS 0.010822f
C124 B.n90 VSUBS 0.010822f
C125 B.n91 VSUBS 0.010822f
C126 B.n92 VSUBS 0.010822f
C127 B.n93 VSUBS 0.010822f
C128 B.n94 VSUBS 0.010822f
C129 B.n95 VSUBS 0.010822f
C130 B.n96 VSUBS 0.010822f
C131 B.n97 VSUBS 0.010822f
C132 B.n98 VSUBS 0.010822f
C133 B.n99 VSUBS 0.010822f
C134 B.n100 VSUBS 0.010822f
C135 B.n101 VSUBS 0.010822f
C136 B.n102 VSUBS 0.010822f
C137 B.n103 VSUBS 0.010822f
C138 B.n104 VSUBS 0.010822f
C139 B.n105 VSUBS 0.010822f
C140 B.n106 VSUBS 0.010822f
C141 B.n107 VSUBS 0.010822f
C142 B.n108 VSUBS 0.010822f
C143 B.n109 VSUBS 0.010822f
C144 B.n110 VSUBS 0.010822f
C145 B.n111 VSUBS 0.010822f
C146 B.n112 VSUBS 0.010822f
C147 B.n113 VSUBS 0.010822f
C148 B.n114 VSUBS 0.010822f
C149 B.n115 VSUBS 0.010822f
C150 B.n116 VSUBS 0.010822f
C151 B.n117 VSUBS 0.010822f
C152 B.n118 VSUBS 0.010822f
C153 B.n119 VSUBS 0.010822f
C154 B.n120 VSUBS 0.010822f
C155 B.n121 VSUBS 0.010822f
C156 B.n122 VSUBS 0.010822f
C157 B.n123 VSUBS 0.010822f
C158 B.n124 VSUBS 0.010822f
C159 B.n125 VSUBS 0.010822f
C160 B.n126 VSUBS 0.010822f
C161 B.n127 VSUBS 0.010822f
C162 B.n128 VSUBS 0.010822f
C163 B.n129 VSUBS 0.010822f
C164 B.n130 VSUBS 0.010822f
C165 B.n131 VSUBS 0.010822f
C166 B.n132 VSUBS 0.010822f
C167 B.n133 VSUBS 0.010822f
C168 B.n134 VSUBS 0.010822f
C169 B.n135 VSUBS 0.010822f
C170 B.n136 VSUBS 0.010822f
C171 B.n137 VSUBS 0.010822f
C172 B.n138 VSUBS 0.010822f
C173 B.n139 VSUBS 0.010822f
C174 B.n140 VSUBS 0.010822f
C175 B.n141 VSUBS 0.010822f
C176 B.n142 VSUBS 0.010822f
C177 B.n143 VSUBS 0.010822f
C178 B.n144 VSUBS 0.024458f
C179 B.n145 VSUBS 0.010822f
C180 B.n146 VSUBS 0.010822f
C181 B.n147 VSUBS 0.010822f
C182 B.n148 VSUBS 0.010822f
C183 B.n149 VSUBS 0.010822f
C184 B.n150 VSUBS 0.010822f
C185 B.n151 VSUBS 0.010822f
C186 B.n152 VSUBS 0.010822f
C187 B.n153 VSUBS 0.010822f
C188 B.n154 VSUBS 0.010822f
C189 B.n155 VSUBS 0.010822f
C190 B.n156 VSUBS 0.010822f
C191 B.n157 VSUBS 0.010822f
C192 B.n158 VSUBS 0.010822f
C193 B.t11 VSUBS 0.18033f
C194 B.t10 VSUBS 0.230575f
C195 B.t9 VSUBS 1.71365f
C196 B.n159 VSUBS 0.380043f
C197 B.n160 VSUBS 0.285508f
C198 B.n161 VSUBS 0.010822f
C199 B.n162 VSUBS 0.010822f
C200 B.n163 VSUBS 0.010822f
C201 B.n164 VSUBS 0.010822f
C202 B.n165 VSUBS 0.006048f
C203 B.n166 VSUBS 0.010822f
C204 B.n167 VSUBS 0.010822f
C205 B.n168 VSUBS 0.010822f
C206 B.n169 VSUBS 0.010822f
C207 B.n170 VSUBS 0.010822f
C208 B.n171 VSUBS 0.010822f
C209 B.n172 VSUBS 0.010822f
C210 B.n173 VSUBS 0.010822f
C211 B.n174 VSUBS 0.010822f
C212 B.n175 VSUBS 0.010822f
C213 B.n176 VSUBS 0.010822f
C214 B.n177 VSUBS 0.010822f
C215 B.n178 VSUBS 0.010822f
C216 B.n179 VSUBS 0.025197f
C217 B.n180 VSUBS 0.010822f
C218 B.n181 VSUBS 0.010822f
C219 B.n182 VSUBS 0.010822f
C220 B.n183 VSUBS 0.010822f
C221 B.n184 VSUBS 0.010822f
C222 B.n185 VSUBS 0.010822f
C223 B.n186 VSUBS 0.010822f
C224 B.n187 VSUBS 0.010822f
C225 B.n188 VSUBS 0.010822f
C226 B.n189 VSUBS 0.010822f
C227 B.n190 VSUBS 0.010822f
C228 B.n191 VSUBS 0.010822f
C229 B.n192 VSUBS 0.010822f
C230 B.n193 VSUBS 0.010822f
C231 B.n194 VSUBS 0.010822f
C232 B.n195 VSUBS 0.010822f
C233 B.n196 VSUBS 0.010822f
C234 B.n197 VSUBS 0.010822f
C235 B.n198 VSUBS 0.010822f
C236 B.n199 VSUBS 0.010822f
C237 B.n200 VSUBS 0.010822f
C238 B.n201 VSUBS 0.010822f
C239 B.n202 VSUBS 0.010822f
C240 B.n203 VSUBS 0.010822f
C241 B.n204 VSUBS 0.010822f
C242 B.n205 VSUBS 0.010822f
C243 B.n206 VSUBS 0.010822f
C244 B.n207 VSUBS 0.010822f
C245 B.n208 VSUBS 0.010822f
C246 B.n209 VSUBS 0.010822f
C247 B.n210 VSUBS 0.010822f
C248 B.n211 VSUBS 0.010822f
C249 B.n212 VSUBS 0.010822f
C250 B.n213 VSUBS 0.010822f
C251 B.n214 VSUBS 0.010822f
C252 B.n215 VSUBS 0.010822f
C253 B.n216 VSUBS 0.010822f
C254 B.n217 VSUBS 0.010822f
C255 B.n218 VSUBS 0.010822f
C256 B.n219 VSUBS 0.010822f
C257 B.n220 VSUBS 0.010822f
C258 B.n221 VSUBS 0.010822f
C259 B.n222 VSUBS 0.010822f
C260 B.n223 VSUBS 0.010822f
C261 B.n224 VSUBS 0.010822f
C262 B.n225 VSUBS 0.010822f
C263 B.n226 VSUBS 0.010822f
C264 B.n227 VSUBS 0.010822f
C265 B.n228 VSUBS 0.010822f
C266 B.n229 VSUBS 0.010822f
C267 B.n230 VSUBS 0.010822f
C268 B.n231 VSUBS 0.010822f
C269 B.n232 VSUBS 0.010822f
C270 B.n233 VSUBS 0.010822f
C271 B.n234 VSUBS 0.010822f
C272 B.n235 VSUBS 0.010822f
C273 B.n236 VSUBS 0.010822f
C274 B.n237 VSUBS 0.010822f
C275 B.n238 VSUBS 0.010822f
C276 B.n239 VSUBS 0.010822f
C277 B.n240 VSUBS 0.010822f
C278 B.n241 VSUBS 0.010822f
C279 B.n242 VSUBS 0.010822f
C280 B.n243 VSUBS 0.010822f
C281 B.n244 VSUBS 0.010822f
C282 B.n245 VSUBS 0.010822f
C283 B.n246 VSUBS 0.010822f
C284 B.n247 VSUBS 0.010822f
C285 B.n248 VSUBS 0.010822f
C286 B.n249 VSUBS 0.010822f
C287 B.n250 VSUBS 0.010822f
C288 B.n251 VSUBS 0.010822f
C289 B.n252 VSUBS 0.010822f
C290 B.n253 VSUBS 0.010822f
C291 B.n254 VSUBS 0.010822f
C292 B.n255 VSUBS 0.010822f
C293 B.n256 VSUBS 0.010822f
C294 B.n257 VSUBS 0.010822f
C295 B.n258 VSUBS 0.010822f
C296 B.n259 VSUBS 0.010822f
C297 B.n260 VSUBS 0.010822f
C298 B.n261 VSUBS 0.010822f
C299 B.n262 VSUBS 0.010822f
C300 B.n263 VSUBS 0.010822f
C301 B.n264 VSUBS 0.010822f
C302 B.n265 VSUBS 0.010822f
C303 B.n266 VSUBS 0.010822f
C304 B.n267 VSUBS 0.010822f
C305 B.n268 VSUBS 0.010822f
C306 B.n269 VSUBS 0.010822f
C307 B.n270 VSUBS 0.010822f
C308 B.n271 VSUBS 0.010822f
C309 B.n272 VSUBS 0.010822f
C310 B.n273 VSUBS 0.010822f
C311 B.n274 VSUBS 0.010822f
C312 B.n275 VSUBS 0.010822f
C313 B.n276 VSUBS 0.010822f
C314 B.n277 VSUBS 0.010822f
C315 B.n278 VSUBS 0.010822f
C316 B.n279 VSUBS 0.010822f
C317 B.n280 VSUBS 0.010822f
C318 B.n281 VSUBS 0.010822f
C319 B.n282 VSUBS 0.010822f
C320 B.n283 VSUBS 0.010822f
C321 B.n284 VSUBS 0.010822f
C322 B.n285 VSUBS 0.010822f
C323 B.n286 VSUBS 0.010822f
C324 B.n287 VSUBS 0.010822f
C325 B.n288 VSUBS 0.010822f
C326 B.n289 VSUBS 0.010822f
C327 B.n290 VSUBS 0.010822f
C328 B.n291 VSUBS 0.010822f
C329 B.n292 VSUBS 0.010822f
C330 B.n293 VSUBS 0.010822f
C331 B.n294 VSUBS 0.010822f
C332 B.n295 VSUBS 0.010822f
C333 B.n296 VSUBS 0.010822f
C334 B.n297 VSUBS 0.010822f
C335 B.n298 VSUBS 0.010822f
C336 B.n299 VSUBS 0.010822f
C337 B.n300 VSUBS 0.010822f
C338 B.n301 VSUBS 0.010822f
C339 B.n302 VSUBS 0.010822f
C340 B.n303 VSUBS 0.010822f
C341 B.n304 VSUBS 0.010822f
C342 B.n305 VSUBS 0.010822f
C343 B.n306 VSUBS 0.010822f
C344 B.n307 VSUBS 0.010822f
C345 B.n308 VSUBS 0.010822f
C346 B.n309 VSUBS 0.010822f
C347 B.n310 VSUBS 0.010822f
C348 B.n311 VSUBS 0.010822f
C349 B.n312 VSUBS 0.010822f
C350 B.n313 VSUBS 0.010822f
C351 B.n314 VSUBS 0.024458f
C352 B.n315 VSUBS 0.024458f
C353 B.n316 VSUBS 0.025197f
C354 B.n317 VSUBS 0.010822f
C355 B.n318 VSUBS 0.010822f
C356 B.n319 VSUBS 0.010822f
C357 B.n320 VSUBS 0.010822f
C358 B.n321 VSUBS 0.010822f
C359 B.n322 VSUBS 0.010822f
C360 B.n323 VSUBS 0.010822f
C361 B.n324 VSUBS 0.010822f
C362 B.n325 VSUBS 0.010822f
C363 B.n326 VSUBS 0.010822f
C364 B.n327 VSUBS 0.010822f
C365 B.n328 VSUBS 0.010822f
C366 B.n329 VSUBS 0.010822f
C367 B.n330 VSUBS 0.010822f
C368 B.n331 VSUBS 0.010822f
C369 B.n332 VSUBS 0.010822f
C370 B.n333 VSUBS 0.010822f
C371 B.n334 VSUBS 0.010822f
C372 B.n335 VSUBS 0.010822f
C373 B.n336 VSUBS 0.010822f
C374 B.n337 VSUBS 0.010822f
C375 B.n338 VSUBS 0.010822f
C376 B.n339 VSUBS 0.010822f
C377 B.n340 VSUBS 0.010822f
C378 B.n341 VSUBS 0.010822f
C379 B.n342 VSUBS 0.010822f
C380 B.n343 VSUBS 0.010822f
C381 B.n344 VSUBS 0.010822f
C382 B.n345 VSUBS 0.010822f
C383 B.n346 VSUBS 0.010822f
C384 B.n347 VSUBS 0.010822f
C385 B.n348 VSUBS 0.010822f
C386 B.n349 VSUBS 0.010822f
C387 B.n350 VSUBS 0.010822f
C388 B.n351 VSUBS 0.010822f
C389 B.n352 VSUBS 0.010822f
C390 B.n353 VSUBS 0.010822f
C391 B.n354 VSUBS 0.010822f
C392 B.n355 VSUBS 0.010822f
C393 B.t5 VSUBS 0.180326f
C394 B.t4 VSUBS 0.230572f
C395 B.t3 VSUBS 1.71365f
C396 B.n356 VSUBS 0.380046f
C397 B.n357 VSUBS 0.285511f
C398 B.n358 VSUBS 0.025074f
C399 B.n359 VSUBS 0.010185f
C400 B.n360 VSUBS 0.010822f
C401 B.n361 VSUBS 0.010822f
C402 B.n362 VSUBS 0.010822f
C403 B.n363 VSUBS 0.010822f
C404 B.n364 VSUBS 0.010822f
C405 B.n365 VSUBS 0.010822f
C406 B.n366 VSUBS 0.010822f
C407 B.n367 VSUBS 0.010822f
C408 B.n368 VSUBS 0.010822f
C409 B.n369 VSUBS 0.010822f
C410 B.n370 VSUBS 0.010822f
C411 B.n371 VSUBS 0.010822f
C412 B.n372 VSUBS 0.010822f
C413 B.n373 VSUBS 0.010822f
C414 B.n374 VSUBS 0.010822f
C415 B.n375 VSUBS 0.006048f
C416 B.n376 VSUBS 0.025074f
C417 B.n377 VSUBS 0.010185f
C418 B.n378 VSUBS 0.010822f
C419 B.n379 VSUBS 0.010822f
C420 B.n380 VSUBS 0.010822f
C421 B.n381 VSUBS 0.010822f
C422 B.n382 VSUBS 0.010822f
C423 B.n383 VSUBS 0.010822f
C424 B.n384 VSUBS 0.010822f
C425 B.n385 VSUBS 0.010822f
C426 B.n386 VSUBS 0.010822f
C427 B.n387 VSUBS 0.010822f
C428 B.n388 VSUBS 0.010822f
C429 B.n389 VSUBS 0.010822f
C430 B.n390 VSUBS 0.010822f
C431 B.n391 VSUBS 0.010822f
C432 B.n392 VSUBS 0.010822f
C433 B.n393 VSUBS 0.010822f
C434 B.n394 VSUBS 0.010822f
C435 B.n395 VSUBS 0.010822f
C436 B.n396 VSUBS 0.010822f
C437 B.n397 VSUBS 0.010822f
C438 B.n398 VSUBS 0.010822f
C439 B.n399 VSUBS 0.010822f
C440 B.n400 VSUBS 0.010822f
C441 B.n401 VSUBS 0.010822f
C442 B.n402 VSUBS 0.010822f
C443 B.n403 VSUBS 0.010822f
C444 B.n404 VSUBS 0.010822f
C445 B.n405 VSUBS 0.010822f
C446 B.n406 VSUBS 0.010822f
C447 B.n407 VSUBS 0.010822f
C448 B.n408 VSUBS 0.010822f
C449 B.n409 VSUBS 0.010822f
C450 B.n410 VSUBS 0.010822f
C451 B.n411 VSUBS 0.010822f
C452 B.n412 VSUBS 0.010822f
C453 B.n413 VSUBS 0.010822f
C454 B.n414 VSUBS 0.010822f
C455 B.n415 VSUBS 0.010822f
C456 B.n416 VSUBS 0.010822f
C457 B.n417 VSUBS 0.025197f
C458 B.n418 VSUBS 0.023879f
C459 B.n419 VSUBS 0.025775f
C460 B.n420 VSUBS 0.010822f
C461 B.n421 VSUBS 0.010822f
C462 B.n422 VSUBS 0.010822f
C463 B.n423 VSUBS 0.010822f
C464 B.n424 VSUBS 0.010822f
C465 B.n425 VSUBS 0.010822f
C466 B.n426 VSUBS 0.010822f
C467 B.n427 VSUBS 0.010822f
C468 B.n428 VSUBS 0.010822f
C469 B.n429 VSUBS 0.010822f
C470 B.n430 VSUBS 0.010822f
C471 B.n431 VSUBS 0.010822f
C472 B.n432 VSUBS 0.010822f
C473 B.n433 VSUBS 0.010822f
C474 B.n434 VSUBS 0.010822f
C475 B.n435 VSUBS 0.010822f
C476 B.n436 VSUBS 0.010822f
C477 B.n437 VSUBS 0.010822f
C478 B.n438 VSUBS 0.010822f
C479 B.n439 VSUBS 0.010822f
C480 B.n440 VSUBS 0.010822f
C481 B.n441 VSUBS 0.010822f
C482 B.n442 VSUBS 0.010822f
C483 B.n443 VSUBS 0.010822f
C484 B.n444 VSUBS 0.010822f
C485 B.n445 VSUBS 0.010822f
C486 B.n446 VSUBS 0.010822f
C487 B.n447 VSUBS 0.010822f
C488 B.n448 VSUBS 0.010822f
C489 B.n449 VSUBS 0.010822f
C490 B.n450 VSUBS 0.010822f
C491 B.n451 VSUBS 0.010822f
C492 B.n452 VSUBS 0.010822f
C493 B.n453 VSUBS 0.010822f
C494 B.n454 VSUBS 0.010822f
C495 B.n455 VSUBS 0.010822f
C496 B.n456 VSUBS 0.010822f
C497 B.n457 VSUBS 0.010822f
C498 B.n458 VSUBS 0.010822f
C499 B.n459 VSUBS 0.010822f
C500 B.n460 VSUBS 0.010822f
C501 B.n461 VSUBS 0.010822f
C502 B.n462 VSUBS 0.010822f
C503 B.n463 VSUBS 0.010822f
C504 B.n464 VSUBS 0.010822f
C505 B.n465 VSUBS 0.010822f
C506 B.n466 VSUBS 0.010822f
C507 B.n467 VSUBS 0.010822f
C508 B.n468 VSUBS 0.010822f
C509 B.n469 VSUBS 0.010822f
C510 B.n470 VSUBS 0.010822f
C511 B.n471 VSUBS 0.010822f
C512 B.n472 VSUBS 0.010822f
C513 B.n473 VSUBS 0.010822f
C514 B.n474 VSUBS 0.010822f
C515 B.n475 VSUBS 0.010822f
C516 B.n476 VSUBS 0.010822f
C517 B.n477 VSUBS 0.010822f
C518 B.n478 VSUBS 0.010822f
C519 B.n479 VSUBS 0.010822f
C520 B.n480 VSUBS 0.010822f
C521 B.n481 VSUBS 0.010822f
C522 B.n482 VSUBS 0.010822f
C523 B.n483 VSUBS 0.010822f
C524 B.n484 VSUBS 0.010822f
C525 B.n485 VSUBS 0.010822f
C526 B.n486 VSUBS 0.010822f
C527 B.n487 VSUBS 0.010822f
C528 B.n488 VSUBS 0.010822f
C529 B.n489 VSUBS 0.010822f
C530 B.n490 VSUBS 0.010822f
C531 B.n491 VSUBS 0.010822f
C532 B.n492 VSUBS 0.010822f
C533 B.n493 VSUBS 0.010822f
C534 B.n494 VSUBS 0.010822f
C535 B.n495 VSUBS 0.010822f
C536 B.n496 VSUBS 0.010822f
C537 B.n497 VSUBS 0.010822f
C538 B.n498 VSUBS 0.010822f
C539 B.n499 VSUBS 0.010822f
C540 B.n500 VSUBS 0.010822f
C541 B.n501 VSUBS 0.010822f
C542 B.n502 VSUBS 0.010822f
C543 B.n503 VSUBS 0.010822f
C544 B.n504 VSUBS 0.010822f
C545 B.n505 VSUBS 0.010822f
C546 B.n506 VSUBS 0.010822f
C547 B.n507 VSUBS 0.010822f
C548 B.n508 VSUBS 0.010822f
C549 B.n509 VSUBS 0.010822f
C550 B.n510 VSUBS 0.010822f
C551 B.n511 VSUBS 0.010822f
C552 B.n512 VSUBS 0.010822f
C553 B.n513 VSUBS 0.010822f
C554 B.n514 VSUBS 0.010822f
C555 B.n515 VSUBS 0.010822f
C556 B.n516 VSUBS 0.010822f
C557 B.n517 VSUBS 0.010822f
C558 B.n518 VSUBS 0.010822f
C559 B.n519 VSUBS 0.010822f
C560 B.n520 VSUBS 0.010822f
C561 B.n521 VSUBS 0.010822f
C562 B.n522 VSUBS 0.010822f
C563 B.n523 VSUBS 0.010822f
C564 B.n524 VSUBS 0.010822f
C565 B.n525 VSUBS 0.010822f
C566 B.n526 VSUBS 0.010822f
C567 B.n527 VSUBS 0.010822f
C568 B.n528 VSUBS 0.010822f
C569 B.n529 VSUBS 0.010822f
C570 B.n530 VSUBS 0.010822f
C571 B.n531 VSUBS 0.010822f
C572 B.n532 VSUBS 0.010822f
C573 B.n533 VSUBS 0.010822f
C574 B.n534 VSUBS 0.010822f
C575 B.n535 VSUBS 0.010822f
C576 B.n536 VSUBS 0.010822f
C577 B.n537 VSUBS 0.010822f
C578 B.n538 VSUBS 0.010822f
C579 B.n539 VSUBS 0.010822f
C580 B.n540 VSUBS 0.010822f
C581 B.n541 VSUBS 0.010822f
C582 B.n542 VSUBS 0.010822f
C583 B.n543 VSUBS 0.010822f
C584 B.n544 VSUBS 0.010822f
C585 B.n545 VSUBS 0.010822f
C586 B.n546 VSUBS 0.010822f
C587 B.n547 VSUBS 0.010822f
C588 B.n548 VSUBS 0.010822f
C589 B.n549 VSUBS 0.010822f
C590 B.n550 VSUBS 0.010822f
C591 B.n551 VSUBS 0.010822f
C592 B.n552 VSUBS 0.010822f
C593 B.n553 VSUBS 0.010822f
C594 B.n554 VSUBS 0.010822f
C595 B.n555 VSUBS 0.010822f
C596 B.n556 VSUBS 0.010822f
C597 B.n557 VSUBS 0.010822f
C598 B.n558 VSUBS 0.010822f
C599 B.n559 VSUBS 0.010822f
C600 B.n560 VSUBS 0.010822f
C601 B.n561 VSUBS 0.010822f
C602 B.n562 VSUBS 0.010822f
C603 B.n563 VSUBS 0.010822f
C604 B.n564 VSUBS 0.010822f
C605 B.n565 VSUBS 0.010822f
C606 B.n566 VSUBS 0.010822f
C607 B.n567 VSUBS 0.010822f
C608 B.n568 VSUBS 0.010822f
C609 B.n569 VSUBS 0.010822f
C610 B.n570 VSUBS 0.010822f
C611 B.n571 VSUBS 0.010822f
C612 B.n572 VSUBS 0.010822f
C613 B.n573 VSUBS 0.010822f
C614 B.n574 VSUBS 0.010822f
C615 B.n575 VSUBS 0.010822f
C616 B.n576 VSUBS 0.010822f
C617 B.n577 VSUBS 0.010822f
C618 B.n578 VSUBS 0.010822f
C619 B.n579 VSUBS 0.010822f
C620 B.n580 VSUBS 0.010822f
C621 B.n581 VSUBS 0.010822f
C622 B.n582 VSUBS 0.010822f
C623 B.n583 VSUBS 0.010822f
C624 B.n584 VSUBS 0.010822f
C625 B.n585 VSUBS 0.010822f
C626 B.n586 VSUBS 0.010822f
C627 B.n587 VSUBS 0.010822f
C628 B.n588 VSUBS 0.010822f
C629 B.n589 VSUBS 0.010822f
C630 B.n590 VSUBS 0.010822f
C631 B.n591 VSUBS 0.010822f
C632 B.n592 VSUBS 0.010822f
C633 B.n593 VSUBS 0.010822f
C634 B.n594 VSUBS 0.010822f
C635 B.n595 VSUBS 0.010822f
C636 B.n596 VSUBS 0.010822f
C637 B.n597 VSUBS 0.010822f
C638 B.n598 VSUBS 0.010822f
C639 B.n599 VSUBS 0.010822f
C640 B.n600 VSUBS 0.010822f
C641 B.n601 VSUBS 0.010822f
C642 B.n602 VSUBS 0.010822f
C643 B.n603 VSUBS 0.010822f
C644 B.n604 VSUBS 0.010822f
C645 B.n605 VSUBS 0.010822f
C646 B.n606 VSUBS 0.010822f
C647 B.n607 VSUBS 0.010822f
C648 B.n608 VSUBS 0.010822f
C649 B.n609 VSUBS 0.010822f
C650 B.n610 VSUBS 0.010822f
C651 B.n611 VSUBS 0.010822f
C652 B.n612 VSUBS 0.010822f
C653 B.n613 VSUBS 0.010822f
C654 B.n614 VSUBS 0.010822f
C655 B.n615 VSUBS 0.010822f
C656 B.n616 VSUBS 0.010822f
C657 B.n617 VSUBS 0.010822f
C658 B.n618 VSUBS 0.010822f
C659 B.n619 VSUBS 0.010822f
C660 B.n620 VSUBS 0.010822f
C661 B.n621 VSUBS 0.010822f
C662 B.n622 VSUBS 0.010822f
C663 B.n623 VSUBS 0.010822f
C664 B.n624 VSUBS 0.010822f
C665 B.n625 VSUBS 0.010822f
C666 B.n626 VSUBS 0.010822f
C667 B.n627 VSUBS 0.024458f
C668 B.n628 VSUBS 0.024458f
C669 B.n629 VSUBS 0.025197f
C670 B.n630 VSUBS 0.010822f
C671 B.n631 VSUBS 0.010822f
C672 B.n632 VSUBS 0.010822f
C673 B.n633 VSUBS 0.010822f
C674 B.n634 VSUBS 0.010822f
C675 B.n635 VSUBS 0.010822f
C676 B.n636 VSUBS 0.010822f
C677 B.n637 VSUBS 0.010822f
C678 B.n638 VSUBS 0.010822f
C679 B.n639 VSUBS 0.010822f
C680 B.n640 VSUBS 0.010822f
C681 B.n641 VSUBS 0.010822f
C682 B.n642 VSUBS 0.010822f
C683 B.n643 VSUBS 0.010822f
C684 B.n644 VSUBS 0.010822f
C685 B.n645 VSUBS 0.010822f
C686 B.n646 VSUBS 0.010822f
C687 B.n647 VSUBS 0.010822f
C688 B.n648 VSUBS 0.010822f
C689 B.n649 VSUBS 0.010822f
C690 B.n650 VSUBS 0.010822f
C691 B.n651 VSUBS 0.010822f
C692 B.n652 VSUBS 0.010822f
C693 B.n653 VSUBS 0.010822f
C694 B.n654 VSUBS 0.010822f
C695 B.n655 VSUBS 0.010822f
C696 B.n656 VSUBS 0.010822f
C697 B.n657 VSUBS 0.010822f
C698 B.n658 VSUBS 0.010822f
C699 B.n659 VSUBS 0.010822f
C700 B.n660 VSUBS 0.010822f
C701 B.n661 VSUBS 0.010822f
C702 B.n662 VSUBS 0.010822f
C703 B.n663 VSUBS 0.010822f
C704 B.n664 VSUBS 0.010822f
C705 B.n665 VSUBS 0.010822f
C706 B.n666 VSUBS 0.010822f
C707 B.n667 VSUBS 0.010822f
C708 B.n668 VSUBS 0.010822f
C709 B.n669 VSUBS 0.010822f
C710 B.n670 VSUBS 0.010185f
C711 B.n671 VSUBS 0.025074f
C712 B.n672 VSUBS 0.006048f
C713 B.n673 VSUBS 0.010822f
C714 B.n674 VSUBS 0.010822f
C715 B.n675 VSUBS 0.010822f
C716 B.n676 VSUBS 0.010822f
C717 B.n677 VSUBS 0.010822f
C718 B.n678 VSUBS 0.010822f
C719 B.n679 VSUBS 0.010822f
C720 B.n680 VSUBS 0.010822f
C721 B.n681 VSUBS 0.010822f
C722 B.n682 VSUBS 0.010822f
C723 B.n683 VSUBS 0.010822f
C724 B.n684 VSUBS 0.010822f
C725 B.n685 VSUBS 0.006048f
C726 B.n686 VSUBS 0.010822f
C727 B.n687 VSUBS 0.010822f
C728 B.n688 VSUBS 0.010822f
C729 B.n689 VSUBS 0.010822f
C730 B.n690 VSUBS 0.010822f
C731 B.n691 VSUBS 0.010822f
C732 B.n692 VSUBS 0.010822f
C733 B.n693 VSUBS 0.010822f
C734 B.n694 VSUBS 0.010822f
C735 B.n695 VSUBS 0.010822f
C736 B.n696 VSUBS 0.010822f
C737 B.n697 VSUBS 0.010822f
C738 B.n698 VSUBS 0.010822f
C739 B.n699 VSUBS 0.010822f
C740 B.n700 VSUBS 0.010822f
C741 B.n701 VSUBS 0.010822f
C742 B.n702 VSUBS 0.010822f
C743 B.n703 VSUBS 0.010822f
C744 B.n704 VSUBS 0.010822f
C745 B.n705 VSUBS 0.010822f
C746 B.n706 VSUBS 0.010822f
C747 B.n707 VSUBS 0.010822f
C748 B.n708 VSUBS 0.010822f
C749 B.n709 VSUBS 0.010822f
C750 B.n710 VSUBS 0.010822f
C751 B.n711 VSUBS 0.010822f
C752 B.n712 VSUBS 0.010822f
C753 B.n713 VSUBS 0.010822f
C754 B.n714 VSUBS 0.010822f
C755 B.n715 VSUBS 0.010822f
C756 B.n716 VSUBS 0.010822f
C757 B.n717 VSUBS 0.010822f
C758 B.n718 VSUBS 0.010822f
C759 B.n719 VSUBS 0.010822f
C760 B.n720 VSUBS 0.010822f
C761 B.n721 VSUBS 0.010822f
C762 B.n722 VSUBS 0.010822f
C763 B.n723 VSUBS 0.010822f
C764 B.n724 VSUBS 0.010822f
C765 B.n725 VSUBS 0.010822f
C766 B.n726 VSUBS 0.010822f
C767 B.n727 VSUBS 0.025197f
C768 B.n728 VSUBS 0.025197f
C769 B.n729 VSUBS 0.024458f
C770 B.n730 VSUBS 0.010822f
C771 B.n731 VSUBS 0.010822f
C772 B.n732 VSUBS 0.010822f
C773 B.n733 VSUBS 0.010822f
C774 B.n734 VSUBS 0.010822f
C775 B.n735 VSUBS 0.010822f
C776 B.n736 VSUBS 0.010822f
C777 B.n737 VSUBS 0.010822f
C778 B.n738 VSUBS 0.010822f
C779 B.n739 VSUBS 0.010822f
C780 B.n740 VSUBS 0.010822f
C781 B.n741 VSUBS 0.010822f
C782 B.n742 VSUBS 0.010822f
C783 B.n743 VSUBS 0.010822f
C784 B.n744 VSUBS 0.010822f
C785 B.n745 VSUBS 0.010822f
C786 B.n746 VSUBS 0.010822f
C787 B.n747 VSUBS 0.010822f
C788 B.n748 VSUBS 0.010822f
C789 B.n749 VSUBS 0.010822f
C790 B.n750 VSUBS 0.010822f
C791 B.n751 VSUBS 0.010822f
C792 B.n752 VSUBS 0.010822f
C793 B.n753 VSUBS 0.010822f
C794 B.n754 VSUBS 0.010822f
C795 B.n755 VSUBS 0.010822f
C796 B.n756 VSUBS 0.010822f
C797 B.n757 VSUBS 0.010822f
C798 B.n758 VSUBS 0.010822f
C799 B.n759 VSUBS 0.010822f
C800 B.n760 VSUBS 0.010822f
C801 B.n761 VSUBS 0.010822f
C802 B.n762 VSUBS 0.010822f
C803 B.n763 VSUBS 0.010822f
C804 B.n764 VSUBS 0.010822f
C805 B.n765 VSUBS 0.010822f
C806 B.n766 VSUBS 0.010822f
C807 B.n767 VSUBS 0.010822f
C808 B.n768 VSUBS 0.010822f
C809 B.n769 VSUBS 0.010822f
C810 B.n770 VSUBS 0.010822f
C811 B.n771 VSUBS 0.010822f
C812 B.n772 VSUBS 0.010822f
C813 B.n773 VSUBS 0.010822f
C814 B.n774 VSUBS 0.010822f
C815 B.n775 VSUBS 0.010822f
C816 B.n776 VSUBS 0.010822f
C817 B.n777 VSUBS 0.010822f
C818 B.n778 VSUBS 0.010822f
C819 B.n779 VSUBS 0.010822f
C820 B.n780 VSUBS 0.010822f
C821 B.n781 VSUBS 0.010822f
C822 B.n782 VSUBS 0.010822f
C823 B.n783 VSUBS 0.010822f
C824 B.n784 VSUBS 0.010822f
C825 B.n785 VSUBS 0.010822f
C826 B.n786 VSUBS 0.010822f
C827 B.n787 VSUBS 0.010822f
C828 B.n788 VSUBS 0.010822f
C829 B.n789 VSUBS 0.010822f
C830 B.n790 VSUBS 0.010822f
C831 B.n791 VSUBS 0.010822f
C832 B.n792 VSUBS 0.010822f
C833 B.n793 VSUBS 0.010822f
C834 B.n794 VSUBS 0.010822f
C835 B.n795 VSUBS 0.010822f
C836 B.n796 VSUBS 0.010822f
C837 B.n797 VSUBS 0.010822f
C838 B.n798 VSUBS 0.010822f
C839 B.n799 VSUBS 0.010822f
C840 B.n800 VSUBS 0.010822f
C841 B.n801 VSUBS 0.010822f
C842 B.n802 VSUBS 0.010822f
C843 B.n803 VSUBS 0.010822f
C844 B.n804 VSUBS 0.010822f
C845 B.n805 VSUBS 0.010822f
C846 B.n806 VSUBS 0.010822f
C847 B.n807 VSUBS 0.010822f
C848 B.n808 VSUBS 0.010822f
C849 B.n809 VSUBS 0.010822f
C850 B.n810 VSUBS 0.010822f
C851 B.n811 VSUBS 0.010822f
C852 B.n812 VSUBS 0.010822f
C853 B.n813 VSUBS 0.010822f
C854 B.n814 VSUBS 0.010822f
C855 B.n815 VSUBS 0.010822f
C856 B.n816 VSUBS 0.010822f
C857 B.n817 VSUBS 0.010822f
C858 B.n818 VSUBS 0.010822f
C859 B.n819 VSUBS 0.010822f
C860 B.n820 VSUBS 0.010822f
C861 B.n821 VSUBS 0.010822f
C862 B.n822 VSUBS 0.010822f
C863 B.n823 VSUBS 0.010822f
C864 B.n824 VSUBS 0.010822f
C865 B.n825 VSUBS 0.010822f
C866 B.n826 VSUBS 0.010822f
C867 B.n827 VSUBS 0.010822f
C868 B.n828 VSUBS 0.010822f
C869 B.n829 VSUBS 0.010822f
C870 B.n830 VSUBS 0.010822f
C871 B.n831 VSUBS 0.014122f
C872 B.n832 VSUBS 0.015044f
C873 B.n833 VSUBS 0.029916f
C874 VDD2.n0 VSUBS 0.038093f
C875 VDD2.n1 VSUBS 0.033379f
C876 VDD2.n2 VSUBS 0.017936f
C877 VDD2.n3 VSUBS 0.042395f
C878 VDD2.n4 VSUBS 0.018991f
C879 VDD2.n5 VSUBS 0.033379f
C880 VDD2.n6 VSUBS 0.017936f
C881 VDD2.n7 VSUBS 0.042395f
C882 VDD2.n8 VSUBS 0.018991f
C883 VDD2.n9 VSUBS 0.033379f
C884 VDD2.n10 VSUBS 0.017936f
C885 VDD2.n11 VSUBS 0.031796f
C886 VDD2.n12 VSUBS 0.026968f
C887 VDD2.t7 VSUBS 0.090541f
C888 VDD2.n13 VSUBS 0.161555f
C889 VDD2.n14 VSUBS 0.989467f
C890 VDD2.n15 VSUBS 0.017936f
C891 VDD2.n16 VSUBS 0.018991f
C892 VDD2.n17 VSUBS 0.042395f
C893 VDD2.n18 VSUBS 0.042395f
C894 VDD2.n19 VSUBS 0.018991f
C895 VDD2.n20 VSUBS 0.017936f
C896 VDD2.n21 VSUBS 0.033379f
C897 VDD2.n22 VSUBS 0.033379f
C898 VDD2.n23 VSUBS 0.017936f
C899 VDD2.n24 VSUBS 0.018991f
C900 VDD2.n25 VSUBS 0.042395f
C901 VDD2.n26 VSUBS 0.042395f
C902 VDD2.n27 VSUBS 0.018991f
C903 VDD2.n28 VSUBS 0.017936f
C904 VDD2.n29 VSUBS 0.033379f
C905 VDD2.n30 VSUBS 0.033379f
C906 VDD2.n31 VSUBS 0.017936f
C907 VDD2.n32 VSUBS 0.018991f
C908 VDD2.n33 VSUBS 0.042395f
C909 VDD2.n34 VSUBS 0.107459f
C910 VDD2.n35 VSUBS 0.018991f
C911 VDD2.n36 VSUBS 0.017936f
C912 VDD2.n37 VSUBS 0.078521f
C913 VDD2.n38 VSUBS 0.099398f
C914 VDD2.t5 VSUBS 0.197034f
C915 VDD2.t3 VSUBS 0.197034f
C916 VDD2.n39 VSUBS 1.38376f
C917 VDD2.n40 VSUBS 1.33804f
C918 VDD2.t1 VSUBS 0.197034f
C919 VDD2.t9 VSUBS 0.197034f
C920 VDD2.n41 VSUBS 1.41225f
C921 VDD2.n42 VSUBS 4.18435f
C922 VDD2.n43 VSUBS 0.038093f
C923 VDD2.n44 VSUBS 0.033379f
C924 VDD2.n45 VSUBS 0.017936f
C925 VDD2.n46 VSUBS 0.042395f
C926 VDD2.n47 VSUBS 0.018991f
C927 VDD2.n48 VSUBS 0.033379f
C928 VDD2.n49 VSUBS 0.017936f
C929 VDD2.n50 VSUBS 0.042395f
C930 VDD2.n51 VSUBS 0.018991f
C931 VDD2.n52 VSUBS 0.033379f
C932 VDD2.n53 VSUBS 0.017936f
C933 VDD2.n54 VSUBS 0.031796f
C934 VDD2.n55 VSUBS 0.026968f
C935 VDD2.t2 VSUBS 0.090541f
C936 VDD2.n56 VSUBS 0.161555f
C937 VDD2.n57 VSUBS 0.989467f
C938 VDD2.n58 VSUBS 0.017936f
C939 VDD2.n59 VSUBS 0.018991f
C940 VDD2.n60 VSUBS 0.042395f
C941 VDD2.n61 VSUBS 0.042395f
C942 VDD2.n62 VSUBS 0.018991f
C943 VDD2.n63 VSUBS 0.017936f
C944 VDD2.n64 VSUBS 0.033379f
C945 VDD2.n65 VSUBS 0.033379f
C946 VDD2.n66 VSUBS 0.017936f
C947 VDD2.n67 VSUBS 0.018991f
C948 VDD2.n68 VSUBS 0.042395f
C949 VDD2.n69 VSUBS 0.042395f
C950 VDD2.n70 VSUBS 0.018991f
C951 VDD2.n71 VSUBS 0.017936f
C952 VDD2.n72 VSUBS 0.033379f
C953 VDD2.n73 VSUBS 0.033379f
C954 VDD2.n74 VSUBS 0.017936f
C955 VDD2.n75 VSUBS 0.018991f
C956 VDD2.n76 VSUBS 0.042395f
C957 VDD2.n77 VSUBS 0.107459f
C958 VDD2.n78 VSUBS 0.018991f
C959 VDD2.n79 VSUBS 0.017936f
C960 VDD2.n80 VSUBS 0.078521f
C961 VDD2.n81 VSUBS 0.077332f
C962 VDD2.n82 VSUBS 3.67239f
C963 VDD2.t0 VSUBS 0.197034f
C964 VDD2.t8 VSUBS 0.197034f
C965 VDD2.n83 VSUBS 1.38377f
C966 VDD2.n84 VSUBS 0.984402f
C967 VDD2.t6 VSUBS 0.197034f
C968 VDD2.t4 VSUBS 0.197034f
C969 VDD2.n85 VSUBS 1.4122f
C970 VN.t0 VSUBS 1.89925f
C971 VN.n0 VSUBS 0.818255f
C972 VN.n1 VSUBS 0.030242f
C973 VN.n2 VSUBS 0.040359f
C974 VN.n3 VSUBS 0.030242f
C975 VN.t8 VSUBS 1.89925f
C976 VN.n4 VSUBS 0.690479f
C977 VN.n5 VSUBS 0.030242f
C978 VN.n6 VSUBS 0.042887f
C979 VN.n7 VSUBS 0.030242f
C980 VN.t6 VSUBS 1.89925f
C981 VN.n8 VSUBS 0.056364f
C982 VN.n9 VSUBS 0.030242f
C983 VN.n10 VSUBS 0.056364f
C984 VN.t2 VSUBS 2.2342f
C985 VN.n11 VSUBS 0.754901f
C986 VN.t4 VSUBS 1.89925f
C987 VN.n12 VSUBS 0.802617f
C988 VN.n13 VSUBS 0.054694f
C989 VN.n14 VSUBS 0.345017f
C990 VN.n15 VSUBS 0.030242f
C991 VN.n16 VSUBS 0.030242f
C992 VN.n17 VSUBS 0.045415f
C993 VN.n18 VSUBS 0.042887f
C994 VN.n19 VSUBS 0.056364f
C995 VN.n20 VSUBS 0.030242f
C996 VN.n21 VSUBS 0.030242f
C997 VN.n22 VSUBS 0.030242f
C998 VN.n23 VSUBS 0.719016f
C999 VN.n24 VSUBS 0.056364f
C1000 VN.n25 VSUBS 0.056364f
C1001 VN.n26 VSUBS 0.030242f
C1002 VN.n27 VSUBS 0.030242f
C1003 VN.n28 VSUBS 0.030242f
C1004 VN.n29 VSUBS 0.045415f
C1005 VN.n30 VSUBS 0.056364f
C1006 VN.n31 VSUBS 0.054694f
C1007 VN.n32 VSUBS 0.030242f
C1008 VN.n33 VSUBS 0.030242f
C1009 VN.n34 VSUBS 0.030206f
C1010 VN.n35 VSUBS 0.056364f
C1011 VN.n36 VSUBS 0.056364f
C1012 VN.n37 VSUBS 0.030242f
C1013 VN.n38 VSUBS 0.030242f
C1014 VN.n39 VSUBS 0.030242f
C1015 VN.n40 VSUBS 0.047943f
C1016 VN.n41 VSUBS 0.056364f
C1017 VN.n42 VSUBS 0.053025f
C1018 VN.n43 VSUBS 0.048811f
C1019 VN.n44 VSUBS 0.062048f
C1020 VN.t7 VSUBS 1.89925f
C1021 VN.n45 VSUBS 0.818255f
C1022 VN.n46 VSUBS 0.030242f
C1023 VN.n47 VSUBS 0.040359f
C1024 VN.n48 VSUBS 0.030242f
C1025 VN.t9 VSUBS 1.89925f
C1026 VN.n49 VSUBS 0.690479f
C1027 VN.n50 VSUBS 0.030242f
C1028 VN.n51 VSUBS 0.042887f
C1029 VN.n52 VSUBS 0.030242f
C1030 VN.t1 VSUBS 1.89925f
C1031 VN.n53 VSUBS 0.056364f
C1032 VN.n54 VSUBS 0.030242f
C1033 VN.n55 VSUBS 0.056364f
C1034 VN.t5 VSUBS 2.2342f
C1035 VN.n56 VSUBS 0.754901f
C1036 VN.t3 VSUBS 1.89925f
C1037 VN.n57 VSUBS 0.802617f
C1038 VN.n58 VSUBS 0.054694f
C1039 VN.n59 VSUBS 0.345017f
C1040 VN.n60 VSUBS 0.030242f
C1041 VN.n61 VSUBS 0.030242f
C1042 VN.n62 VSUBS 0.045415f
C1043 VN.n63 VSUBS 0.042887f
C1044 VN.n64 VSUBS 0.056364f
C1045 VN.n65 VSUBS 0.030242f
C1046 VN.n66 VSUBS 0.030242f
C1047 VN.n67 VSUBS 0.030242f
C1048 VN.n68 VSUBS 0.719016f
C1049 VN.n69 VSUBS 0.056364f
C1050 VN.n70 VSUBS 0.056364f
C1051 VN.n71 VSUBS 0.030242f
C1052 VN.n72 VSUBS 0.030242f
C1053 VN.n73 VSUBS 0.030242f
C1054 VN.n74 VSUBS 0.045415f
C1055 VN.n75 VSUBS 0.056364f
C1056 VN.n76 VSUBS 0.054694f
C1057 VN.n77 VSUBS 0.030242f
C1058 VN.n78 VSUBS 0.030242f
C1059 VN.n79 VSUBS 0.030206f
C1060 VN.n80 VSUBS 0.056364f
C1061 VN.n81 VSUBS 0.056364f
C1062 VN.n82 VSUBS 0.030242f
C1063 VN.n83 VSUBS 0.030242f
C1064 VN.n84 VSUBS 0.030242f
C1065 VN.n85 VSUBS 0.047943f
C1066 VN.n86 VSUBS 0.056364f
C1067 VN.n87 VSUBS 0.053025f
C1068 VN.n88 VSUBS 0.048811f
C1069 VN.n89 VSUBS 1.86114f
C1070 VTAIL.t7 VSUBS 0.190356f
C1071 VTAIL.t5 VSUBS 0.190356f
C1072 VTAIL.n0 VSUBS 1.20423f
C1073 VTAIL.n1 VSUBS 1.08866f
C1074 VTAIL.n2 VSUBS 0.036802f
C1075 VTAIL.n3 VSUBS 0.032247f
C1076 VTAIL.n4 VSUBS 0.017328f
C1077 VTAIL.n5 VSUBS 0.040958f
C1078 VTAIL.n6 VSUBS 0.018348f
C1079 VTAIL.n7 VSUBS 0.032247f
C1080 VTAIL.n8 VSUBS 0.017328f
C1081 VTAIL.n9 VSUBS 0.040958f
C1082 VTAIL.n10 VSUBS 0.018348f
C1083 VTAIL.n11 VSUBS 0.032247f
C1084 VTAIL.n12 VSUBS 0.017328f
C1085 VTAIL.n13 VSUBS 0.030718f
C1086 VTAIL.n14 VSUBS 0.026054f
C1087 VTAIL.t14 VSUBS 0.087472f
C1088 VTAIL.n15 VSUBS 0.156079f
C1089 VTAIL.n16 VSUBS 0.955929f
C1090 VTAIL.n17 VSUBS 0.017328f
C1091 VTAIL.n18 VSUBS 0.018348f
C1092 VTAIL.n19 VSUBS 0.040958f
C1093 VTAIL.n20 VSUBS 0.040958f
C1094 VTAIL.n21 VSUBS 0.018348f
C1095 VTAIL.n22 VSUBS 0.017328f
C1096 VTAIL.n23 VSUBS 0.032247f
C1097 VTAIL.n24 VSUBS 0.032247f
C1098 VTAIL.n25 VSUBS 0.017328f
C1099 VTAIL.n26 VSUBS 0.018348f
C1100 VTAIL.n27 VSUBS 0.040958f
C1101 VTAIL.n28 VSUBS 0.040958f
C1102 VTAIL.n29 VSUBS 0.018348f
C1103 VTAIL.n30 VSUBS 0.017328f
C1104 VTAIL.n31 VSUBS 0.032247f
C1105 VTAIL.n32 VSUBS 0.032247f
C1106 VTAIL.n33 VSUBS 0.017328f
C1107 VTAIL.n34 VSUBS 0.018348f
C1108 VTAIL.n35 VSUBS 0.040958f
C1109 VTAIL.n36 VSUBS 0.103817f
C1110 VTAIL.n37 VSUBS 0.018348f
C1111 VTAIL.n38 VSUBS 0.017328f
C1112 VTAIL.n39 VSUBS 0.075859f
C1113 VTAIL.n40 VSUBS 0.052456f
C1114 VTAIL.n41 VSUBS 0.543348f
C1115 VTAIL.t10 VSUBS 0.190356f
C1116 VTAIL.t9 VSUBS 0.190356f
C1117 VTAIL.n42 VSUBS 1.20423f
C1118 VTAIL.n43 VSUBS 1.26692f
C1119 VTAIL.t12 VSUBS 0.190356f
C1120 VTAIL.t17 VSUBS 0.190356f
C1121 VTAIL.n44 VSUBS 1.20423f
C1122 VTAIL.n45 VSUBS 2.68492f
C1123 VTAIL.t4 VSUBS 0.190356f
C1124 VTAIL.t1 VSUBS 0.190356f
C1125 VTAIL.n46 VSUBS 1.20424f
C1126 VTAIL.n47 VSUBS 2.68491f
C1127 VTAIL.t18 VSUBS 0.190356f
C1128 VTAIL.t6 VSUBS 0.190356f
C1129 VTAIL.n48 VSUBS 1.20424f
C1130 VTAIL.n49 VSUBS 1.26691f
C1131 VTAIL.n50 VSUBS 0.036802f
C1132 VTAIL.n51 VSUBS 0.032247f
C1133 VTAIL.n52 VSUBS 0.017328f
C1134 VTAIL.n53 VSUBS 0.040958f
C1135 VTAIL.n54 VSUBS 0.018348f
C1136 VTAIL.n55 VSUBS 0.032247f
C1137 VTAIL.n56 VSUBS 0.017328f
C1138 VTAIL.n57 VSUBS 0.040958f
C1139 VTAIL.n58 VSUBS 0.018348f
C1140 VTAIL.n59 VSUBS 0.032247f
C1141 VTAIL.n60 VSUBS 0.017328f
C1142 VTAIL.n61 VSUBS 0.030718f
C1143 VTAIL.n62 VSUBS 0.026054f
C1144 VTAIL.t0 VSUBS 0.087472f
C1145 VTAIL.n63 VSUBS 0.156079f
C1146 VTAIL.n64 VSUBS 0.955929f
C1147 VTAIL.n65 VSUBS 0.017328f
C1148 VTAIL.n66 VSUBS 0.018348f
C1149 VTAIL.n67 VSUBS 0.040958f
C1150 VTAIL.n68 VSUBS 0.040958f
C1151 VTAIL.n69 VSUBS 0.018348f
C1152 VTAIL.n70 VSUBS 0.017328f
C1153 VTAIL.n71 VSUBS 0.032247f
C1154 VTAIL.n72 VSUBS 0.032247f
C1155 VTAIL.n73 VSUBS 0.017328f
C1156 VTAIL.n74 VSUBS 0.018348f
C1157 VTAIL.n75 VSUBS 0.040958f
C1158 VTAIL.n76 VSUBS 0.040958f
C1159 VTAIL.n77 VSUBS 0.018348f
C1160 VTAIL.n78 VSUBS 0.017328f
C1161 VTAIL.n79 VSUBS 0.032247f
C1162 VTAIL.n80 VSUBS 0.032247f
C1163 VTAIL.n81 VSUBS 0.017328f
C1164 VTAIL.n82 VSUBS 0.018348f
C1165 VTAIL.n83 VSUBS 0.040958f
C1166 VTAIL.n84 VSUBS 0.103817f
C1167 VTAIL.n85 VSUBS 0.018348f
C1168 VTAIL.n86 VSUBS 0.017328f
C1169 VTAIL.n87 VSUBS 0.075859f
C1170 VTAIL.n88 VSUBS 0.052456f
C1171 VTAIL.n89 VSUBS 0.543348f
C1172 VTAIL.t13 VSUBS 0.190356f
C1173 VTAIL.t16 VSUBS 0.190356f
C1174 VTAIL.n90 VSUBS 1.20424f
C1175 VTAIL.n91 VSUBS 1.16031f
C1176 VTAIL.t8 VSUBS 0.190356f
C1177 VTAIL.t11 VSUBS 0.190356f
C1178 VTAIL.n92 VSUBS 1.20424f
C1179 VTAIL.n93 VSUBS 1.26691f
C1180 VTAIL.n94 VSUBS 0.036802f
C1181 VTAIL.n95 VSUBS 0.032247f
C1182 VTAIL.n96 VSUBS 0.017328f
C1183 VTAIL.n97 VSUBS 0.040958f
C1184 VTAIL.n98 VSUBS 0.018348f
C1185 VTAIL.n99 VSUBS 0.032247f
C1186 VTAIL.n100 VSUBS 0.017328f
C1187 VTAIL.n101 VSUBS 0.040958f
C1188 VTAIL.n102 VSUBS 0.018348f
C1189 VTAIL.n103 VSUBS 0.032247f
C1190 VTAIL.n104 VSUBS 0.017328f
C1191 VTAIL.n105 VSUBS 0.030718f
C1192 VTAIL.n106 VSUBS 0.026054f
C1193 VTAIL.t15 VSUBS 0.087472f
C1194 VTAIL.n107 VSUBS 0.156079f
C1195 VTAIL.n108 VSUBS 0.955929f
C1196 VTAIL.n109 VSUBS 0.017328f
C1197 VTAIL.n110 VSUBS 0.018348f
C1198 VTAIL.n111 VSUBS 0.040958f
C1199 VTAIL.n112 VSUBS 0.040958f
C1200 VTAIL.n113 VSUBS 0.018348f
C1201 VTAIL.n114 VSUBS 0.017328f
C1202 VTAIL.n115 VSUBS 0.032247f
C1203 VTAIL.n116 VSUBS 0.032247f
C1204 VTAIL.n117 VSUBS 0.017328f
C1205 VTAIL.n118 VSUBS 0.018348f
C1206 VTAIL.n119 VSUBS 0.040958f
C1207 VTAIL.n120 VSUBS 0.040958f
C1208 VTAIL.n121 VSUBS 0.018348f
C1209 VTAIL.n122 VSUBS 0.017328f
C1210 VTAIL.n123 VSUBS 0.032247f
C1211 VTAIL.n124 VSUBS 0.032247f
C1212 VTAIL.n125 VSUBS 0.017328f
C1213 VTAIL.n126 VSUBS 0.018348f
C1214 VTAIL.n127 VSUBS 0.040958f
C1215 VTAIL.n128 VSUBS 0.103817f
C1216 VTAIL.n129 VSUBS 0.018348f
C1217 VTAIL.n130 VSUBS 0.017328f
C1218 VTAIL.n131 VSUBS 0.075859f
C1219 VTAIL.n132 VSUBS 0.052456f
C1220 VTAIL.n133 VSUBS 1.75711f
C1221 VTAIL.n134 VSUBS 0.036802f
C1222 VTAIL.n135 VSUBS 0.032247f
C1223 VTAIL.n136 VSUBS 0.017328f
C1224 VTAIL.n137 VSUBS 0.040958f
C1225 VTAIL.n138 VSUBS 0.018348f
C1226 VTAIL.n139 VSUBS 0.032247f
C1227 VTAIL.n140 VSUBS 0.017328f
C1228 VTAIL.n141 VSUBS 0.040958f
C1229 VTAIL.n142 VSUBS 0.018348f
C1230 VTAIL.n143 VSUBS 0.032247f
C1231 VTAIL.n144 VSUBS 0.017328f
C1232 VTAIL.n145 VSUBS 0.030718f
C1233 VTAIL.n146 VSUBS 0.026054f
C1234 VTAIL.t19 VSUBS 0.087472f
C1235 VTAIL.n147 VSUBS 0.156079f
C1236 VTAIL.n148 VSUBS 0.955929f
C1237 VTAIL.n149 VSUBS 0.017328f
C1238 VTAIL.n150 VSUBS 0.018348f
C1239 VTAIL.n151 VSUBS 0.040958f
C1240 VTAIL.n152 VSUBS 0.040958f
C1241 VTAIL.n153 VSUBS 0.018348f
C1242 VTAIL.n154 VSUBS 0.017328f
C1243 VTAIL.n155 VSUBS 0.032247f
C1244 VTAIL.n156 VSUBS 0.032247f
C1245 VTAIL.n157 VSUBS 0.017328f
C1246 VTAIL.n158 VSUBS 0.018348f
C1247 VTAIL.n159 VSUBS 0.040958f
C1248 VTAIL.n160 VSUBS 0.040958f
C1249 VTAIL.n161 VSUBS 0.018348f
C1250 VTAIL.n162 VSUBS 0.017328f
C1251 VTAIL.n163 VSUBS 0.032247f
C1252 VTAIL.n164 VSUBS 0.032247f
C1253 VTAIL.n165 VSUBS 0.017328f
C1254 VTAIL.n166 VSUBS 0.018348f
C1255 VTAIL.n167 VSUBS 0.040958f
C1256 VTAIL.n168 VSUBS 0.103817f
C1257 VTAIL.n169 VSUBS 0.018348f
C1258 VTAIL.n170 VSUBS 0.017328f
C1259 VTAIL.n171 VSUBS 0.075859f
C1260 VTAIL.n172 VSUBS 0.052456f
C1261 VTAIL.n173 VSUBS 1.75711f
C1262 VTAIL.t3 VSUBS 0.190356f
C1263 VTAIL.t2 VSUBS 0.190356f
C1264 VTAIL.n174 VSUBS 1.20423f
C1265 VTAIL.n175 VSUBS 1.02775f
C1266 VDD1.n0 VSUBS 0.038055f
C1267 VDD1.n1 VSUBS 0.033346f
C1268 VDD1.n2 VSUBS 0.017919f
C1269 VDD1.n3 VSUBS 0.042353f
C1270 VDD1.n4 VSUBS 0.018973f
C1271 VDD1.n5 VSUBS 0.033346f
C1272 VDD1.n6 VSUBS 0.017919f
C1273 VDD1.n7 VSUBS 0.042353f
C1274 VDD1.n8 VSUBS 0.018973f
C1275 VDD1.n9 VSUBS 0.033346f
C1276 VDD1.n10 VSUBS 0.017919f
C1277 VDD1.n11 VSUBS 0.031765f
C1278 VDD1.n12 VSUBS 0.026941f
C1279 VDD1.t2 VSUBS 0.090452f
C1280 VDD1.n13 VSUBS 0.161397f
C1281 VDD1.n14 VSUBS 0.9885f
C1282 VDD1.n15 VSUBS 0.017919f
C1283 VDD1.n16 VSUBS 0.018973f
C1284 VDD1.n17 VSUBS 0.042353f
C1285 VDD1.n18 VSUBS 0.042353f
C1286 VDD1.n19 VSUBS 0.018973f
C1287 VDD1.n20 VSUBS 0.017919f
C1288 VDD1.n21 VSUBS 0.033346f
C1289 VDD1.n22 VSUBS 0.033346f
C1290 VDD1.n23 VSUBS 0.017919f
C1291 VDD1.n24 VSUBS 0.018973f
C1292 VDD1.n25 VSUBS 0.042353f
C1293 VDD1.n26 VSUBS 0.042353f
C1294 VDD1.n27 VSUBS 0.018973f
C1295 VDD1.n28 VSUBS 0.017919f
C1296 VDD1.n29 VSUBS 0.033346f
C1297 VDD1.n30 VSUBS 0.033346f
C1298 VDD1.n31 VSUBS 0.017919f
C1299 VDD1.n32 VSUBS 0.018973f
C1300 VDD1.n33 VSUBS 0.042353f
C1301 VDD1.n34 VSUBS 0.107354f
C1302 VDD1.n35 VSUBS 0.018973f
C1303 VDD1.n36 VSUBS 0.017919f
C1304 VDD1.n37 VSUBS 0.078444f
C1305 VDD1.n38 VSUBS 0.099301f
C1306 VDD1.t5 VSUBS 0.196842f
C1307 VDD1.t1 VSUBS 0.196842f
C1308 VDD1.n39 VSUBS 1.38241f
C1309 VDD1.n40 VSUBS 1.34781f
C1310 VDD1.n41 VSUBS 0.038055f
C1311 VDD1.n42 VSUBS 0.033346f
C1312 VDD1.n43 VSUBS 0.017919f
C1313 VDD1.n44 VSUBS 0.042353f
C1314 VDD1.n45 VSUBS 0.018973f
C1315 VDD1.n46 VSUBS 0.033346f
C1316 VDD1.n47 VSUBS 0.017919f
C1317 VDD1.n48 VSUBS 0.042353f
C1318 VDD1.n49 VSUBS 0.018973f
C1319 VDD1.n50 VSUBS 0.033346f
C1320 VDD1.n51 VSUBS 0.017919f
C1321 VDD1.n52 VSUBS 0.031765f
C1322 VDD1.n53 VSUBS 0.026941f
C1323 VDD1.t3 VSUBS 0.090452f
C1324 VDD1.n54 VSUBS 0.161397f
C1325 VDD1.n55 VSUBS 0.9885f
C1326 VDD1.n56 VSUBS 0.017919f
C1327 VDD1.n57 VSUBS 0.018973f
C1328 VDD1.n58 VSUBS 0.042353f
C1329 VDD1.n59 VSUBS 0.042353f
C1330 VDD1.n60 VSUBS 0.018973f
C1331 VDD1.n61 VSUBS 0.017919f
C1332 VDD1.n62 VSUBS 0.033346f
C1333 VDD1.n63 VSUBS 0.033346f
C1334 VDD1.n64 VSUBS 0.017919f
C1335 VDD1.n65 VSUBS 0.018973f
C1336 VDD1.n66 VSUBS 0.042353f
C1337 VDD1.n67 VSUBS 0.042353f
C1338 VDD1.n68 VSUBS 0.018973f
C1339 VDD1.n69 VSUBS 0.017919f
C1340 VDD1.n70 VSUBS 0.033346f
C1341 VDD1.n71 VSUBS 0.033346f
C1342 VDD1.n72 VSUBS 0.017919f
C1343 VDD1.n73 VSUBS 0.018973f
C1344 VDD1.n74 VSUBS 0.042353f
C1345 VDD1.n75 VSUBS 0.107354f
C1346 VDD1.n76 VSUBS 0.018973f
C1347 VDD1.n77 VSUBS 0.017919f
C1348 VDD1.n78 VSUBS 0.078444f
C1349 VDD1.n79 VSUBS 0.099301f
C1350 VDD1.t9 VSUBS 0.196842f
C1351 VDD1.t7 VSUBS 0.196842f
C1352 VDD1.n80 VSUBS 1.38241f
C1353 VDD1.n81 VSUBS 1.33673f
C1354 VDD1.t6 VSUBS 0.196842f
C1355 VDD1.t8 VSUBS 0.196842f
C1356 VDD1.n82 VSUBS 1.41087f
C1357 VDD1.n83 VSUBS 4.36161f
C1358 VDD1.t4 VSUBS 0.196842f
C1359 VDD1.t0 VSUBS 0.196842f
C1360 VDD1.n84 VSUBS 1.38241f
C1361 VDD1.n85 VSUBS 4.36929f
C1362 VP.t3 VSUBS 2.09828f
C1363 VP.n0 VSUBS 0.904007f
C1364 VP.n1 VSUBS 0.033412f
C1365 VP.n2 VSUBS 0.044589f
C1366 VP.n3 VSUBS 0.033412f
C1367 VP.t8 VSUBS 2.09828f
C1368 VP.n4 VSUBS 0.762839f
C1369 VP.n5 VSUBS 0.033412f
C1370 VP.n6 VSUBS 0.047382f
C1371 VP.n7 VSUBS 0.033412f
C1372 VP.t7 VSUBS 2.09828f
C1373 VP.n8 VSUBS 0.062271f
C1374 VP.n9 VSUBS 0.033412f
C1375 VP.n10 VSUBS 0.062271f
C1376 VP.n11 VSUBS 0.033412f
C1377 VP.t0 VSUBS 2.09828f
C1378 VP.n12 VSUBS 0.062271f
C1379 VP.n13 VSUBS 0.033412f
C1380 VP.n14 VSUBS 0.058582f
C1381 VP.t2 VSUBS 2.09828f
C1382 VP.n15 VSUBS 0.904007f
C1383 VP.n16 VSUBS 0.033412f
C1384 VP.n17 VSUBS 0.044589f
C1385 VP.n18 VSUBS 0.033412f
C1386 VP.t6 VSUBS 2.09828f
C1387 VP.n19 VSUBS 0.762839f
C1388 VP.n20 VSUBS 0.033412f
C1389 VP.n21 VSUBS 0.047382f
C1390 VP.n22 VSUBS 0.033412f
C1391 VP.t9 VSUBS 2.09828f
C1392 VP.n23 VSUBS 0.062271f
C1393 VP.n24 VSUBS 0.033412f
C1394 VP.n25 VSUBS 0.062271f
C1395 VP.t4 VSUBS 2.46834f
C1396 VP.n26 VSUBS 0.834015f
C1397 VP.t1 VSUBS 2.09828f
C1398 VP.n27 VSUBS 0.88673f
C1399 VP.n28 VSUBS 0.060426f
C1400 VP.n29 VSUBS 0.381174f
C1401 VP.n30 VSUBS 0.033412f
C1402 VP.n31 VSUBS 0.033412f
C1403 VP.n32 VSUBS 0.050175f
C1404 VP.n33 VSUBS 0.047382f
C1405 VP.n34 VSUBS 0.062271f
C1406 VP.n35 VSUBS 0.033412f
C1407 VP.n36 VSUBS 0.033412f
C1408 VP.n37 VSUBS 0.033412f
C1409 VP.n38 VSUBS 0.794367f
C1410 VP.n39 VSUBS 0.062271f
C1411 VP.n40 VSUBS 0.062271f
C1412 VP.n41 VSUBS 0.033412f
C1413 VP.n42 VSUBS 0.033412f
C1414 VP.n43 VSUBS 0.033412f
C1415 VP.n44 VSUBS 0.050175f
C1416 VP.n45 VSUBS 0.062271f
C1417 VP.n46 VSUBS 0.060426f
C1418 VP.n47 VSUBS 0.033412f
C1419 VP.n48 VSUBS 0.033412f
C1420 VP.n49 VSUBS 0.033372f
C1421 VP.n50 VSUBS 0.062271f
C1422 VP.n51 VSUBS 0.062271f
C1423 VP.n52 VSUBS 0.033412f
C1424 VP.n53 VSUBS 0.033412f
C1425 VP.n54 VSUBS 0.033412f
C1426 VP.n55 VSUBS 0.052968f
C1427 VP.n56 VSUBS 0.062271f
C1428 VP.n57 VSUBS 0.058582f
C1429 VP.n58 VSUBS 0.053926f
C1430 VP.n59 VSUBS 2.04277f
C1431 VP.t5 VSUBS 2.09828f
C1432 VP.n60 VSUBS 0.904007f
C1433 VP.n61 VSUBS 2.06552f
C1434 VP.n62 VSUBS 0.053926f
C1435 VP.n63 VSUBS 0.033412f
C1436 VP.n64 VSUBS 0.062271f
C1437 VP.n65 VSUBS 0.052968f
C1438 VP.n66 VSUBS 0.044589f
C1439 VP.n67 VSUBS 0.033412f
C1440 VP.n68 VSUBS 0.033412f
C1441 VP.n69 VSUBS 0.033412f
C1442 VP.n70 VSUBS 0.062271f
C1443 VP.n71 VSUBS 0.033372f
C1444 VP.n72 VSUBS 0.762839f
C1445 VP.n73 VSUBS 0.060426f
C1446 VP.n74 VSUBS 0.033412f
C1447 VP.n75 VSUBS 0.033412f
C1448 VP.n76 VSUBS 0.033412f
C1449 VP.n77 VSUBS 0.050175f
C1450 VP.n78 VSUBS 0.047382f
C1451 VP.n79 VSUBS 0.062271f
C1452 VP.n80 VSUBS 0.033412f
C1453 VP.n81 VSUBS 0.033412f
C1454 VP.n82 VSUBS 0.033412f
C1455 VP.n83 VSUBS 0.794367f
C1456 VP.n84 VSUBS 0.062271f
C1457 VP.n85 VSUBS 0.062271f
C1458 VP.n86 VSUBS 0.033412f
C1459 VP.n87 VSUBS 0.033412f
C1460 VP.n88 VSUBS 0.033412f
C1461 VP.n89 VSUBS 0.050175f
C1462 VP.n90 VSUBS 0.062271f
C1463 VP.n91 VSUBS 0.060426f
C1464 VP.n92 VSUBS 0.033412f
C1465 VP.n93 VSUBS 0.033412f
C1466 VP.n94 VSUBS 0.033372f
C1467 VP.n95 VSUBS 0.062271f
C1468 VP.n96 VSUBS 0.062271f
C1469 VP.n97 VSUBS 0.033412f
C1470 VP.n98 VSUBS 0.033412f
C1471 VP.n99 VSUBS 0.033412f
C1472 VP.n100 VSUBS 0.052968f
C1473 VP.n101 VSUBS 0.062271f
C1474 VP.n102 VSUBS 0.058582f
C1475 VP.n103 VSUBS 0.053926f
C1476 VP.n104 VSUBS 0.068551f
.ends

