* NGSPICE file created from diff_pair_sample_0329.ext - technology: sky130A

.subckt diff_pair_sample_0329 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=3.4047 pd=18.24 as=0 ps=0 w=8.73 l=2.78
X1 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=3.4047 pd=18.24 as=0 ps=0 w=8.73 l=2.78
X2 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=3.4047 pd=18.24 as=0 ps=0 w=8.73 l=2.78
X3 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.4047 pd=18.24 as=0 ps=0 w=8.73 l=2.78
X4 VDD2.t1 VN.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=3.4047 pd=18.24 as=3.4047 ps=18.24 w=8.73 l=2.78
X5 VDD2.t0 VN.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=3.4047 pd=18.24 as=3.4047 ps=18.24 w=8.73 l=2.78
X6 VDD1.t1 VP.t0 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=3.4047 pd=18.24 as=3.4047 ps=18.24 w=8.73 l=2.78
X7 VDD1.t0 VP.t1 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=3.4047 pd=18.24 as=3.4047 ps=18.24 w=8.73 l=2.78
R0 B.n448 B.n447 585
R1 B.n450 B.n93 585
R2 B.n453 B.n452 585
R3 B.n454 B.n92 585
R4 B.n456 B.n455 585
R5 B.n458 B.n91 585
R6 B.n461 B.n460 585
R7 B.n462 B.n90 585
R8 B.n464 B.n463 585
R9 B.n466 B.n89 585
R10 B.n469 B.n468 585
R11 B.n470 B.n88 585
R12 B.n472 B.n471 585
R13 B.n474 B.n87 585
R14 B.n477 B.n476 585
R15 B.n478 B.n86 585
R16 B.n480 B.n479 585
R17 B.n482 B.n85 585
R18 B.n485 B.n484 585
R19 B.n486 B.n84 585
R20 B.n488 B.n487 585
R21 B.n490 B.n83 585
R22 B.n493 B.n492 585
R23 B.n494 B.n82 585
R24 B.n496 B.n495 585
R25 B.n498 B.n81 585
R26 B.n501 B.n500 585
R27 B.n502 B.n80 585
R28 B.n504 B.n503 585
R29 B.n506 B.n79 585
R30 B.n508 B.n507 585
R31 B.n510 B.n509 585
R32 B.n513 B.n512 585
R33 B.n514 B.n74 585
R34 B.n516 B.n515 585
R35 B.n518 B.n73 585
R36 B.n521 B.n520 585
R37 B.n522 B.n72 585
R38 B.n524 B.n523 585
R39 B.n526 B.n71 585
R40 B.n529 B.n528 585
R41 B.n530 B.n68 585
R42 B.n533 B.n532 585
R43 B.n535 B.n67 585
R44 B.n538 B.n537 585
R45 B.n539 B.n66 585
R46 B.n541 B.n540 585
R47 B.n543 B.n65 585
R48 B.n546 B.n545 585
R49 B.n547 B.n64 585
R50 B.n549 B.n548 585
R51 B.n551 B.n63 585
R52 B.n554 B.n553 585
R53 B.n555 B.n62 585
R54 B.n557 B.n556 585
R55 B.n559 B.n61 585
R56 B.n562 B.n561 585
R57 B.n563 B.n60 585
R58 B.n565 B.n564 585
R59 B.n567 B.n59 585
R60 B.n570 B.n569 585
R61 B.n571 B.n58 585
R62 B.n573 B.n572 585
R63 B.n575 B.n57 585
R64 B.n578 B.n577 585
R65 B.n579 B.n56 585
R66 B.n581 B.n580 585
R67 B.n583 B.n55 585
R68 B.n586 B.n585 585
R69 B.n587 B.n54 585
R70 B.n589 B.n588 585
R71 B.n591 B.n53 585
R72 B.n594 B.n593 585
R73 B.n595 B.n52 585
R74 B.n446 B.n50 585
R75 B.n598 B.n50 585
R76 B.n445 B.n49 585
R77 B.n599 B.n49 585
R78 B.n444 B.n48 585
R79 B.n600 B.n48 585
R80 B.n443 B.n442 585
R81 B.n442 B.n44 585
R82 B.n441 B.n43 585
R83 B.n606 B.n43 585
R84 B.n440 B.n42 585
R85 B.n607 B.n42 585
R86 B.n439 B.n41 585
R87 B.n608 B.n41 585
R88 B.n438 B.n437 585
R89 B.n437 B.n40 585
R90 B.n436 B.n36 585
R91 B.n614 B.n36 585
R92 B.n435 B.n35 585
R93 B.n615 B.n35 585
R94 B.n434 B.n34 585
R95 B.n616 B.n34 585
R96 B.n433 B.n432 585
R97 B.n432 B.n30 585
R98 B.n431 B.n29 585
R99 B.n622 B.n29 585
R100 B.n430 B.n28 585
R101 B.n623 B.n28 585
R102 B.n429 B.n27 585
R103 B.n624 B.n27 585
R104 B.n428 B.n427 585
R105 B.n427 B.n23 585
R106 B.n426 B.n22 585
R107 B.n630 B.n22 585
R108 B.n425 B.n21 585
R109 B.n631 B.n21 585
R110 B.n424 B.n20 585
R111 B.n632 B.n20 585
R112 B.n423 B.n422 585
R113 B.n422 B.n16 585
R114 B.n421 B.n15 585
R115 B.n638 B.n15 585
R116 B.n420 B.n14 585
R117 B.n639 B.n14 585
R118 B.n419 B.n13 585
R119 B.n640 B.n13 585
R120 B.n418 B.n417 585
R121 B.n417 B.n12 585
R122 B.n416 B.n415 585
R123 B.n416 B.n8 585
R124 B.n414 B.n7 585
R125 B.n647 B.n7 585
R126 B.n413 B.n6 585
R127 B.n648 B.n6 585
R128 B.n412 B.n5 585
R129 B.n649 B.n5 585
R130 B.n411 B.n410 585
R131 B.n410 B.n4 585
R132 B.n409 B.n94 585
R133 B.n409 B.n408 585
R134 B.n399 B.n95 585
R135 B.n96 B.n95 585
R136 B.n401 B.n400 585
R137 B.n402 B.n401 585
R138 B.n398 B.n101 585
R139 B.n101 B.n100 585
R140 B.n397 B.n396 585
R141 B.n396 B.n395 585
R142 B.n103 B.n102 585
R143 B.n104 B.n103 585
R144 B.n388 B.n387 585
R145 B.n389 B.n388 585
R146 B.n386 B.n109 585
R147 B.n109 B.n108 585
R148 B.n385 B.n384 585
R149 B.n384 B.n383 585
R150 B.n111 B.n110 585
R151 B.n112 B.n111 585
R152 B.n376 B.n375 585
R153 B.n377 B.n376 585
R154 B.n374 B.n117 585
R155 B.n117 B.n116 585
R156 B.n373 B.n372 585
R157 B.n372 B.n371 585
R158 B.n119 B.n118 585
R159 B.n120 B.n119 585
R160 B.n364 B.n363 585
R161 B.n365 B.n364 585
R162 B.n362 B.n125 585
R163 B.n125 B.n124 585
R164 B.n361 B.n360 585
R165 B.n360 B.n359 585
R166 B.n127 B.n126 585
R167 B.n352 B.n127 585
R168 B.n351 B.n350 585
R169 B.n353 B.n351 585
R170 B.n349 B.n132 585
R171 B.n132 B.n131 585
R172 B.n348 B.n347 585
R173 B.n347 B.n346 585
R174 B.n134 B.n133 585
R175 B.n135 B.n134 585
R176 B.n339 B.n338 585
R177 B.n340 B.n339 585
R178 B.n337 B.n140 585
R179 B.n140 B.n139 585
R180 B.n336 B.n335 585
R181 B.n335 B.n334 585
R182 B.n331 B.n144 585
R183 B.n330 B.n329 585
R184 B.n327 B.n145 585
R185 B.n327 B.n143 585
R186 B.n326 B.n325 585
R187 B.n324 B.n323 585
R188 B.n322 B.n147 585
R189 B.n320 B.n319 585
R190 B.n318 B.n148 585
R191 B.n317 B.n316 585
R192 B.n314 B.n149 585
R193 B.n312 B.n311 585
R194 B.n310 B.n150 585
R195 B.n309 B.n308 585
R196 B.n306 B.n151 585
R197 B.n304 B.n303 585
R198 B.n302 B.n152 585
R199 B.n301 B.n300 585
R200 B.n298 B.n153 585
R201 B.n296 B.n295 585
R202 B.n294 B.n154 585
R203 B.n293 B.n292 585
R204 B.n290 B.n155 585
R205 B.n288 B.n287 585
R206 B.n286 B.n156 585
R207 B.n285 B.n284 585
R208 B.n282 B.n157 585
R209 B.n280 B.n279 585
R210 B.n278 B.n158 585
R211 B.n277 B.n276 585
R212 B.n274 B.n159 585
R213 B.n272 B.n271 585
R214 B.n270 B.n160 585
R215 B.n268 B.n267 585
R216 B.n265 B.n163 585
R217 B.n263 B.n262 585
R218 B.n261 B.n164 585
R219 B.n260 B.n259 585
R220 B.n257 B.n165 585
R221 B.n255 B.n254 585
R222 B.n253 B.n166 585
R223 B.n252 B.n251 585
R224 B.n249 B.n167 585
R225 B.n247 B.n246 585
R226 B.n245 B.n168 585
R227 B.n244 B.n243 585
R228 B.n241 B.n172 585
R229 B.n239 B.n238 585
R230 B.n237 B.n173 585
R231 B.n236 B.n235 585
R232 B.n233 B.n174 585
R233 B.n231 B.n230 585
R234 B.n229 B.n175 585
R235 B.n228 B.n227 585
R236 B.n225 B.n176 585
R237 B.n223 B.n222 585
R238 B.n221 B.n177 585
R239 B.n220 B.n219 585
R240 B.n217 B.n178 585
R241 B.n215 B.n214 585
R242 B.n213 B.n179 585
R243 B.n212 B.n211 585
R244 B.n209 B.n180 585
R245 B.n207 B.n206 585
R246 B.n205 B.n181 585
R247 B.n204 B.n203 585
R248 B.n201 B.n182 585
R249 B.n199 B.n198 585
R250 B.n197 B.n183 585
R251 B.n196 B.n195 585
R252 B.n193 B.n184 585
R253 B.n191 B.n190 585
R254 B.n189 B.n185 585
R255 B.n188 B.n187 585
R256 B.n142 B.n141 585
R257 B.n143 B.n142 585
R258 B.n333 B.n332 585
R259 B.n334 B.n333 585
R260 B.n138 B.n137 585
R261 B.n139 B.n138 585
R262 B.n342 B.n341 585
R263 B.n341 B.n340 585
R264 B.n343 B.n136 585
R265 B.n136 B.n135 585
R266 B.n345 B.n344 585
R267 B.n346 B.n345 585
R268 B.n130 B.n129 585
R269 B.n131 B.n130 585
R270 B.n355 B.n354 585
R271 B.n354 B.n353 585
R272 B.n356 B.n128 585
R273 B.n352 B.n128 585
R274 B.n358 B.n357 585
R275 B.n359 B.n358 585
R276 B.n123 B.n122 585
R277 B.n124 B.n123 585
R278 B.n367 B.n366 585
R279 B.n366 B.n365 585
R280 B.n368 B.n121 585
R281 B.n121 B.n120 585
R282 B.n370 B.n369 585
R283 B.n371 B.n370 585
R284 B.n115 B.n114 585
R285 B.n116 B.n115 585
R286 B.n379 B.n378 585
R287 B.n378 B.n377 585
R288 B.n380 B.n113 585
R289 B.n113 B.n112 585
R290 B.n382 B.n381 585
R291 B.n383 B.n382 585
R292 B.n107 B.n106 585
R293 B.n108 B.n107 585
R294 B.n391 B.n390 585
R295 B.n390 B.n389 585
R296 B.n392 B.n105 585
R297 B.n105 B.n104 585
R298 B.n394 B.n393 585
R299 B.n395 B.n394 585
R300 B.n99 B.n98 585
R301 B.n100 B.n99 585
R302 B.n404 B.n403 585
R303 B.n403 B.n402 585
R304 B.n405 B.n97 585
R305 B.n97 B.n96 585
R306 B.n407 B.n406 585
R307 B.n408 B.n407 585
R308 B.n3 B.n0 585
R309 B.n4 B.n3 585
R310 B.n646 B.n1 585
R311 B.n647 B.n646 585
R312 B.n645 B.n644 585
R313 B.n645 B.n8 585
R314 B.n643 B.n9 585
R315 B.n12 B.n9 585
R316 B.n642 B.n641 585
R317 B.n641 B.n640 585
R318 B.n11 B.n10 585
R319 B.n639 B.n11 585
R320 B.n637 B.n636 585
R321 B.n638 B.n637 585
R322 B.n635 B.n17 585
R323 B.n17 B.n16 585
R324 B.n634 B.n633 585
R325 B.n633 B.n632 585
R326 B.n19 B.n18 585
R327 B.n631 B.n19 585
R328 B.n629 B.n628 585
R329 B.n630 B.n629 585
R330 B.n627 B.n24 585
R331 B.n24 B.n23 585
R332 B.n626 B.n625 585
R333 B.n625 B.n624 585
R334 B.n26 B.n25 585
R335 B.n623 B.n26 585
R336 B.n621 B.n620 585
R337 B.n622 B.n621 585
R338 B.n619 B.n31 585
R339 B.n31 B.n30 585
R340 B.n618 B.n617 585
R341 B.n617 B.n616 585
R342 B.n33 B.n32 585
R343 B.n615 B.n33 585
R344 B.n613 B.n612 585
R345 B.n614 B.n613 585
R346 B.n611 B.n37 585
R347 B.n40 B.n37 585
R348 B.n610 B.n609 585
R349 B.n609 B.n608 585
R350 B.n39 B.n38 585
R351 B.n607 B.n39 585
R352 B.n605 B.n604 585
R353 B.n606 B.n605 585
R354 B.n603 B.n45 585
R355 B.n45 B.n44 585
R356 B.n602 B.n601 585
R357 B.n601 B.n600 585
R358 B.n47 B.n46 585
R359 B.n599 B.n47 585
R360 B.n597 B.n596 585
R361 B.n598 B.n597 585
R362 B.n650 B.n649 585
R363 B.n648 B.n2 585
R364 B.n597 B.n52 449.257
R365 B.n448 B.n50 449.257
R366 B.n335 B.n142 449.257
R367 B.n333 B.n144 449.257
R368 B.n75 B.t7 286.286
R369 B.n169 B.t12 286.286
R370 B.n69 B.t4 286.286
R371 B.n161 B.t15 286.286
R372 B.n69 B.t2 283.985
R373 B.n75 B.t6 283.985
R374 B.n169 B.t9 283.985
R375 B.n161 B.t13 283.985
R376 B.n449 B.n51 256.663
R377 B.n451 B.n51 256.663
R378 B.n457 B.n51 256.663
R379 B.n459 B.n51 256.663
R380 B.n465 B.n51 256.663
R381 B.n467 B.n51 256.663
R382 B.n473 B.n51 256.663
R383 B.n475 B.n51 256.663
R384 B.n481 B.n51 256.663
R385 B.n483 B.n51 256.663
R386 B.n489 B.n51 256.663
R387 B.n491 B.n51 256.663
R388 B.n497 B.n51 256.663
R389 B.n499 B.n51 256.663
R390 B.n505 B.n51 256.663
R391 B.n78 B.n51 256.663
R392 B.n511 B.n51 256.663
R393 B.n517 B.n51 256.663
R394 B.n519 B.n51 256.663
R395 B.n525 B.n51 256.663
R396 B.n527 B.n51 256.663
R397 B.n534 B.n51 256.663
R398 B.n536 B.n51 256.663
R399 B.n542 B.n51 256.663
R400 B.n544 B.n51 256.663
R401 B.n550 B.n51 256.663
R402 B.n552 B.n51 256.663
R403 B.n558 B.n51 256.663
R404 B.n560 B.n51 256.663
R405 B.n566 B.n51 256.663
R406 B.n568 B.n51 256.663
R407 B.n574 B.n51 256.663
R408 B.n576 B.n51 256.663
R409 B.n582 B.n51 256.663
R410 B.n584 B.n51 256.663
R411 B.n590 B.n51 256.663
R412 B.n592 B.n51 256.663
R413 B.n328 B.n143 256.663
R414 B.n146 B.n143 256.663
R415 B.n321 B.n143 256.663
R416 B.n315 B.n143 256.663
R417 B.n313 B.n143 256.663
R418 B.n307 B.n143 256.663
R419 B.n305 B.n143 256.663
R420 B.n299 B.n143 256.663
R421 B.n297 B.n143 256.663
R422 B.n291 B.n143 256.663
R423 B.n289 B.n143 256.663
R424 B.n283 B.n143 256.663
R425 B.n281 B.n143 256.663
R426 B.n275 B.n143 256.663
R427 B.n273 B.n143 256.663
R428 B.n266 B.n143 256.663
R429 B.n264 B.n143 256.663
R430 B.n258 B.n143 256.663
R431 B.n256 B.n143 256.663
R432 B.n250 B.n143 256.663
R433 B.n248 B.n143 256.663
R434 B.n242 B.n143 256.663
R435 B.n240 B.n143 256.663
R436 B.n234 B.n143 256.663
R437 B.n232 B.n143 256.663
R438 B.n226 B.n143 256.663
R439 B.n224 B.n143 256.663
R440 B.n218 B.n143 256.663
R441 B.n216 B.n143 256.663
R442 B.n210 B.n143 256.663
R443 B.n208 B.n143 256.663
R444 B.n202 B.n143 256.663
R445 B.n200 B.n143 256.663
R446 B.n194 B.n143 256.663
R447 B.n192 B.n143 256.663
R448 B.n186 B.n143 256.663
R449 B.n652 B.n651 256.663
R450 B.n76 B.t8 225.97
R451 B.n170 B.t11 225.97
R452 B.n70 B.t5 225.97
R453 B.n162 B.t14 225.97
R454 B.n593 B.n591 163.367
R455 B.n589 B.n54 163.367
R456 B.n585 B.n583 163.367
R457 B.n581 B.n56 163.367
R458 B.n577 B.n575 163.367
R459 B.n573 B.n58 163.367
R460 B.n569 B.n567 163.367
R461 B.n565 B.n60 163.367
R462 B.n561 B.n559 163.367
R463 B.n557 B.n62 163.367
R464 B.n553 B.n551 163.367
R465 B.n549 B.n64 163.367
R466 B.n545 B.n543 163.367
R467 B.n541 B.n66 163.367
R468 B.n537 B.n535 163.367
R469 B.n533 B.n68 163.367
R470 B.n528 B.n526 163.367
R471 B.n524 B.n72 163.367
R472 B.n520 B.n518 163.367
R473 B.n516 B.n74 163.367
R474 B.n512 B.n510 163.367
R475 B.n507 B.n506 163.367
R476 B.n504 B.n80 163.367
R477 B.n500 B.n498 163.367
R478 B.n496 B.n82 163.367
R479 B.n492 B.n490 163.367
R480 B.n488 B.n84 163.367
R481 B.n484 B.n482 163.367
R482 B.n480 B.n86 163.367
R483 B.n476 B.n474 163.367
R484 B.n472 B.n88 163.367
R485 B.n468 B.n466 163.367
R486 B.n464 B.n90 163.367
R487 B.n460 B.n458 163.367
R488 B.n456 B.n92 163.367
R489 B.n452 B.n450 163.367
R490 B.n335 B.n140 163.367
R491 B.n339 B.n140 163.367
R492 B.n339 B.n134 163.367
R493 B.n347 B.n134 163.367
R494 B.n347 B.n132 163.367
R495 B.n351 B.n132 163.367
R496 B.n351 B.n127 163.367
R497 B.n360 B.n127 163.367
R498 B.n360 B.n125 163.367
R499 B.n364 B.n125 163.367
R500 B.n364 B.n119 163.367
R501 B.n372 B.n119 163.367
R502 B.n372 B.n117 163.367
R503 B.n376 B.n117 163.367
R504 B.n376 B.n111 163.367
R505 B.n384 B.n111 163.367
R506 B.n384 B.n109 163.367
R507 B.n388 B.n109 163.367
R508 B.n388 B.n103 163.367
R509 B.n396 B.n103 163.367
R510 B.n396 B.n101 163.367
R511 B.n401 B.n101 163.367
R512 B.n401 B.n95 163.367
R513 B.n409 B.n95 163.367
R514 B.n410 B.n409 163.367
R515 B.n410 B.n5 163.367
R516 B.n6 B.n5 163.367
R517 B.n7 B.n6 163.367
R518 B.n416 B.n7 163.367
R519 B.n417 B.n416 163.367
R520 B.n417 B.n13 163.367
R521 B.n14 B.n13 163.367
R522 B.n15 B.n14 163.367
R523 B.n422 B.n15 163.367
R524 B.n422 B.n20 163.367
R525 B.n21 B.n20 163.367
R526 B.n22 B.n21 163.367
R527 B.n427 B.n22 163.367
R528 B.n427 B.n27 163.367
R529 B.n28 B.n27 163.367
R530 B.n29 B.n28 163.367
R531 B.n432 B.n29 163.367
R532 B.n432 B.n34 163.367
R533 B.n35 B.n34 163.367
R534 B.n36 B.n35 163.367
R535 B.n437 B.n36 163.367
R536 B.n437 B.n41 163.367
R537 B.n42 B.n41 163.367
R538 B.n43 B.n42 163.367
R539 B.n442 B.n43 163.367
R540 B.n442 B.n48 163.367
R541 B.n49 B.n48 163.367
R542 B.n50 B.n49 163.367
R543 B.n329 B.n327 163.367
R544 B.n327 B.n326 163.367
R545 B.n323 B.n322 163.367
R546 B.n320 B.n148 163.367
R547 B.n316 B.n314 163.367
R548 B.n312 B.n150 163.367
R549 B.n308 B.n306 163.367
R550 B.n304 B.n152 163.367
R551 B.n300 B.n298 163.367
R552 B.n296 B.n154 163.367
R553 B.n292 B.n290 163.367
R554 B.n288 B.n156 163.367
R555 B.n284 B.n282 163.367
R556 B.n280 B.n158 163.367
R557 B.n276 B.n274 163.367
R558 B.n272 B.n160 163.367
R559 B.n267 B.n265 163.367
R560 B.n263 B.n164 163.367
R561 B.n259 B.n257 163.367
R562 B.n255 B.n166 163.367
R563 B.n251 B.n249 163.367
R564 B.n247 B.n168 163.367
R565 B.n243 B.n241 163.367
R566 B.n239 B.n173 163.367
R567 B.n235 B.n233 163.367
R568 B.n231 B.n175 163.367
R569 B.n227 B.n225 163.367
R570 B.n223 B.n177 163.367
R571 B.n219 B.n217 163.367
R572 B.n215 B.n179 163.367
R573 B.n211 B.n209 163.367
R574 B.n207 B.n181 163.367
R575 B.n203 B.n201 163.367
R576 B.n199 B.n183 163.367
R577 B.n195 B.n193 163.367
R578 B.n191 B.n185 163.367
R579 B.n187 B.n142 163.367
R580 B.n333 B.n138 163.367
R581 B.n341 B.n138 163.367
R582 B.n341 B.n136 163.367
R583 B.n345 B.n136 163.367
R584 B.n345 B.n130 163.367
R585 B.n354 B.n130 163.367
R586 B.n354 B.n128 163.367
R587 B.n358 B.n128 163.367
R588 B.n358 B.n123 163.367
R589 B.n366 B.n123 163.367
R590 B.n366 B.n121 163.367
R591 B.n370 B.n121 163.367
R592 B.n370 B.n115 163.367
R593 B.n378 B.n115 163.367
R594 B.n378 B.n113 163.367
R595 B.n382 B.n113 163.367
R596 B.n382 B.n107 163.367
R597 B.n390 B.n107 163.367
R598 B.n390 B.n105 163.367
R599 B.n394 B.n105 163.367
R600 B.n394 B.n99 163.367
R601 B.n403 B.n99 163.367
R602 B.n403 B.n97 163.367
R603 B.n407 B.n97 163.367
R604 B.n407 B.n3 163.367
R605 B.n650 B.n3 163.367
R606 B.n646 B.n2 163.367
R607 B.n646 B.n645 163.367
R608 B.n645 B.n9 163.367
R609 B.n641 B.n9 163.367
R610 B.n641 B.n11 163.367
R611 B.n637 B.n11 163.367
R612 B.n637 B.n17 163.367
R613 B.n633 B.n17 163.367
R614 B.n633 B.n19 163.367
R615 B.n629 B.n19 163.367
R616 B.n629 B.n24 163.367
R617 B.n625 B.n24 163.367
R618 B.n625 B.n26 163.367
R619 B.n621 B.n26 163.367
R620 B.n621 B.n31 163.367
R621 B.n617 B.n31 163.367
R622 B.n617 B.n33 163.367
R623 B.n613 B.n33 163.367
R624 B.n613 B.n37 163.367
R625 B.n609 B.n37 163.367
R626 B.n609 B.n39 163.367
R627 B.n605 B.n39 163.367
R628 B.n605 B.n45 163.367
R629 B.n601 B.n45 163.367
R630 B.n601 B.n47 163.367
R631 B.n597 B.n47 163.367
R632 B.n334 B.n143 91.8963
R633 B.n598 B.n51 91.8963
R634 B.n592 B.n52 71.676
R635 B.n591 B.n590 71.676
R636 B.n584 B.n54 71.676
R637 B.n583 B.n582 71.676
R638 B.n576 B.n56 71.676
R639 B.n575 B.n574 71.676
R640 B.n568 B.n58 71.676
R641 B.n567 B.n566 71.676
R642 B.n560 B.n60 71.676
R643 B.n559 B.n558 71.676
R644 B.n552 B.n62 71.676
R645 B.n551 B.n550 71.676
R646 B.n544 B.n64 71.676
R647 B.n543 B.n542 71.676
R648 B.n536 B.n66 71.676
R649 B.n535 B.n534 71.676
R650 B.n527 B.n68 71.676
R651 B.n526 B.n525 71.676
R652 B.n519 B.n72 71.676
R653 B.n518 B.n517 71.676
R654 B.n511 B.n74 71.676
R655 B.n510 B.n78 71.676
R656 B.n506 B.n505 71.676
R657 B.n499 B.n80 71.676
R658 B.n498 B.n497 71.676
R659 B.n491 B.n82 71.676
R660 B.n490 B.n489 71.676
R661 B.n483 B.n84 71.676
R662 B.n482 B.n481 71.676
R663 B.n475 B.n86 71.676
R664 B.n474 B.n473 71.676
R665 B.n467 B.n88 71.676
R666 B.n466 B.n465 71.676
R667 B.n459 B.n90 71.676
R668 B.n458 B.n457 71.676
R669 B.n451 B.n92 71.676
R670 B.n450 B.n449 71.676
R671 B.n449 B.n448 71.676
R672 B.n452 B.n451 71.676
R673 B.n457 B.n456 71.676
R674 B.n460 B.n459 71.676
R675 B.n465 B.n464 71.676
R676 B.n468 B.n467 71.676
R677 B.n473 B.n472 71.676
R678 B.n476 B.n475 71.676
R679 B.n481 B.n480 71.676
R680 B.n484 B.n483 71.676
R681 B.n489 B.n488 71.676
R682 B.n492 B.n491 71.676
R683 B.n497 B.n496 71.676
R684 B.n500 B.n499 71.676
R685 B.n505 B.n504 71.676
R686 B.n507 B.n78 71.676
R687 B.n512 B.n511 71.676
R688 B.n517 B.n516 71.676
R689 B.n520 B.n519 71.676
R690 B.n525 B.n524 71.676
R691 B.n528 B.n527 71.676
R692 B.n534 B.n533 71.676
R693 B.n537 B.n536 71.676
R694 B.n542 B.n541 71.676
R695 B.n545 B.n544 71.676
R696 B.n550 B.n549 71.676
R697 B.n553 B.n552 71.676
R698 B.n558 B.n557 71.676
R699 B.n561 B.n560 71.676
R700 B.n566 B.n565 71.676
R701 B.n569 B.n568 71.676
R702 B.n574 B.n573 71.676
R703 B.n577 B.n576 71.676
R704 B.n582 B.n581 71.676
R705 B.n585 B.n584 71.676
R706 B.n590 B.n589 71.676
R707 B.n593 B.n592 71.676
R708 B.n328 B.n144 71.676
R709 B.n326 B.n146 71.676
R710 B.n322 B.n321 71.676
R711 B.n315 B.n148 71.676
R712 B.n314 B.n313 71.676
R713 B.n307 B.n150 71.676
R714 B.n306 B.n305 71.676
R715 B.n299 B.n152 71.676
R716 B.n298 B.n297 71.676
R717 B.n291 B.n154 71.676
R718 B.n290 B.n289 71.676
R719 B.n283 B.n156 71.676
R720 B.n282 B.n281 71.676
R721 B.n275 B.n158 71.676
R722 B.n274 B.n273 71.676
R723 B.n266 B.n160 71.676
R724 B.n265 B.n264 71.676
R725 B.n258 B.n164 71.676
R726 B.n257 B.n256 71.676
R727 B.n250 B.n166 71.676
R728 B.n249 B.n248 71.676
R729 B.n242 B.n168 71.676
R730 B.n241 B.n240 71.676
R731 B.n234 B.n173 71.676
R732 B.n233 B.n232 71.676
R733 B.n226 B.n175 71.676
R734 B.n225 B.n224 71.676
R735 B.n218 B.n177 71.676
R736 B.n217 B.n216 71.676
R737 B.n210 B.n179 71.676
R738 B.n209 B.n208 71.676
R739 B.n202 B.n181 71.676
R740 B.n201 B.n200 71.676
R741 B.n194 B.n183 71.676
R742 B.n193 B.n192 71.676
R743 B.n186 B.n185 71.676
R744 B.n329 B.n328 71.676
R745 B.n323 B.n146 71.676
R746 B.n321 B.n320 71.676
R747 B.n316 B.n315 71.676
R748 B.n313 B.n312 71.676
R749 B.n308 B.n307 71.676
R750 B.n305 B.n304 71.676
R751 B.n300 B.n299 71.676
R752 B.n297 B.n296 71.676
R753 B.n292 B.n291 71.676
R754 B.n289 B.n288 71.676
R755 B.n284 B.n283 71.676
R756 B.n281 B.n280 71.676
R757 B.n276 B.n275 71.676
R758 B.n273 B.n272 71.676
R759 B.n267 B.n266 71.676
R760 B.n264 B.n263 71.676
R761 B.n259 B.n258 71.676
R762 B.n256 B.n255 71.676
R763 B.n251 B.n250 71.676
R764 B.n248 B.n247 71.676
R765 B.n243 B.n242 71.676
R766 B.n240 B.n239 71.676
R767 B.n235 B.n234 71.676
R768 B.n232 B.n231 71.676
R769 B.n227 B.n226 71.676
R770 B.n224 B.n223 71.676
R771 B.n219 B.n218 71.676
R772 B.n216 B.n215 71.676
R773 B.n211 B.n210 71.676
R774 B.n208 B.n207 71.676
R775 B.n203 B.n202 71.676
R776 B.n200 B.n199 71.676
R777 B.n195 B.n194 71.676
R778 B.n192 B.n191 71.676
R779 B.n187 B.n186 71.676
R780 B.n651 B.n650 71.676
R781 B.n651 B.n2 71.676
R782 B.n70 B.n69 60.3157
R783 B.n76 B.n75 60.3157
R784 B.n170 B.n169 60.3157
R785 B.n162 B.n161 60.3157
R786 B.n531 B.n70 59.5399
R787 B.n77 B.n76 59.5399
R788 B.n171 B.n170 59.5399
R789 B.n269 B.n162 59.5399
R790 B.n334 B.n139 53.41
R791 B.n340 B.n139 53.41
R792 B.n340 B.n135 53.41
R793 B.n346 B.n135 53.41
R794 B.n346 B.n131 53.41
R795 B.n353 B.n131 53.41
R796 B.n353 B.n352 53.41
R797 B.n359 B.n124 53.41
R798 B.n365 B.n124 53.41
R799 B.n365 B.n120 53.41
R800 B.n371 B.n120 53.41
R801 B.n371 B.n116 53.41
R802 B.n377 B.n116 53.41
R803 B.n377 B.n112 53.41
R804 B.n383 B.n112 53.41
R805 B.n383 B.n108 53.41
R806 B.n389 B.n108 53.41
R807 B.n389 B.n104 53.41
R808 B.n395 B.n104 53.41
R809 B.n402 B.n100 53.41
R810 B.n402 B.n96 53.41
R811 B.n408 B.n96 53.41
R812 B.n408 B.n4 53.41
R813 B.n649 B.n4 53.41
R814 B.n649 B.n648 53.41
R815 B.n648 B.n647 53.41
R816 B.n647 B.n8 53.41
R817 B.n12 B.n8 53.41
R818 B.n640 B.n12 53.41
R819 B.n640 B.n639 53.41
R820 B.n638 B.n16 53.41
R821 B.n632 B.n16 53.41
R822 B.n632 B.n631 53.41
R823 B.n631 B.n630 53.41
R824 B.n630 B.n23 53.41
R825 B.n624 B.n23 53.41
R826 B.n624 B.n623 53.41
R827 B.n623 B.n622 53.41
R828 B.n622 B.n30 53.41
R829 B.n616 B.n30 53.41
R830 B.n616 B.n615 53.41
R831 B.n615 B.n614 53.41
R832 B.n608 B.n40 53.41
R833 B.n608 B.n607 53.41
R834 B.n607 B.n606 53.41
R835 B.n606 B.n44 53.41
R836 B.n600 B.n44 53.41
R837 B.n600 B.n599 53.41
R838 B.n599 B.n598 53.41
R839 B.n352 B.t10 51.8391
R840 B.n40 B.t3 51.8391
R841 B.t0 B.n100 36.1305
R842 B.n639 B.t1 36.1305
R843 B.n447 B.n446 29.1907
R844 B.n332 B.n331 29.1907
R845 B.n336 B.n141 29.1907
R846 B.n596 B.n595 29.1907
R847 B B.n652 18.0485
R848 B.n395 B.t0 17.28
R849 B.t1 B.n638 17.28
R850 B.n332 B.n137 10.6151
R851 B.n342 B.n137 10.6151
R852 B.n343 B.n342 10.6151
R853 B.n344 B.n343 10.6151
R854 B.n344 B.n129 10.6151
R855 B.n355 B.n129 10.6151
R856 B.n356 B.n355 10.6151
R857 B.n357 B.n356 10.6151
R858 B.n357 B.n122 10.6151
R859 B.n367 B.n122 10.6151
R860 B.n368 B.n367 10.6151
R861 B.n369 B.n368 10.6151
R862 B.n369 B.n114 10.6151
R863 B.n379 B.n114 10.6151
R864 B.n380 B.n379 10.6151
R865 B.n381 B.n380 10.6151
R866 B.n381 B.n106 10.6151
R867 B.n391 B.n106 10.6151
R868 B.n392 B.n391 10.6151
R869 B.n393 B.n392 10.6151
R870 B.n393 B.n98 10.6151
R871 B.n404 B.n98 10.6151
R872 B.n405 B.n404 10.6151
R873 B.n406 B.n405 10.6151
R874 B.n406 B.n0 10.6151
R875 B.n331 B.n330 10.6151
R876 B.n330 B.n145 10.6151
R877 B.n325 B.n145 10.6151
R878 B.n325 B.n324 10.6151
R879 B.n324 B.n147 10.6151
R880 B.n319 B.n147 10.6151
R881 B.n319 B.n318 10.6151
R882 B.n318 B.n317 10.6151
R883 B.n317 B.n149 10.6151
R884 B.n311 B.n149 10.6151
R885 B.n311 B.n310 10.6151
R886 B.n310 B.n309 10.6151
R887 B.n309 B.n151 10.6151
R888 B.n303 B.n151 10.6151
R889 B.n303 B.n302 10.6151
R890 B.n302 B.n301 10.6151
R891 B.n301 B.n153 10.6151
R892 B.n295 B.n153 10.6151
R893 B.n295 B.n294 10.6151
R894 B.n294 B.n293 10.6151
R895 B.n293 B.n155 10.6151
R896 B.n287 B.n155 10.6151
R897 B.n287 B.n286 10.6151
R898 B.n286 B.n285 10.6151
R899 B.n285 B.n157 10.6151
R900 B.n279 B.n157 10.6151
R901 B.n279 B.n278 10.6151
R902 B.n278 B.n277 10.6151
R903 B.n277 B.n159 10.6151
R904 B.n271 B.n159 10.6151
R905 B.n271 B.n270 10.6151
R906 B.n268 B.n163 10.6151
R907 B.n262 B.n163 10.6151
R908 B.n262 B.n261 10.6151
R909 B.n261 B.n260 10.6151
R910 B.n260 B.n165 10.6151
R911 B.n254 B.n165 10.6151
R912 B.n254 B.n253 10.6151
R913 B.n253 B.n252 10.6151
R914 B.n252 B.n167 10.6151
R915 B.n246 B.n245 10.6151
R916 B.n245 B.n244 10.6151
R917 B.n244 B.n172 10.6151
R918 B.n238 B.n172 10.6151
R919 B.n238 B.n237 10.6151
R920 B.n237 B.n236 10.6151
R921 B.n236 B.n174 10.6151
R922 B.n230 B.n174 10.6151
R923 B.n230 B.n229 10.6151
R924 B.n229 B.n228 10.6151
R925 B.n228 B.n176 10.6151
R926 B.n222 B.n176 10.6151
R927 B.n222 B.n221 10.6151
R928 B.n221 B.n220 10.6151
R929 B.n220 B.n178 10.6151
R930 B.n214 B.n178 10.6151
R931 B.n214 B.n213 10.6151
R932 B.n213 B.n212 10.6151
R933 B.n212 B.n180 10.6151
R934 B.n206 B.n180 10.6151
R935 B.n206 B.n205 10.6151
R936 B.n205 B.n204 10.6151
R937 B.n204 B.n182 10.6151
R938 B.n198 B.n182 10.6151
R939 B.n198 B.n197 10.6151
R940 B.n197 B.n196 10.6151
R941 B.n196 B.n184 10.6151
R942 B.n190 B.n184 10.6151
R943 B.n190 B.n189 10.6151
R944 B.n189 B.n188 10.6151
R945 B.n188 B.n141 10.6151
R946 B.n337 B.n336 10.6151
R947 B.n338 B.n337 10.6151
R948 B.n338 B.n133 10.6151
R949 B.n348 B.n133 10.6151
R950 B.n349 B.n348 10.6151
R951 B.n350 B.n349 10.6151
R952 B.n350 B.n126 10.6151
R953 B.n361 B.n126 10.6151
R954 B.n362 B.n361 10.6151
R955 B.n363 B.n362 10.6151
R956 B.n363 B.n118 10.6151
R957 B.n373 B.n118 10.6151
R958 B.n374 B.n373 10.6151
R959 B.n375 B.n374 10.6151
R960 B.n375 B.n110 10.6151
R961 B.n385 B.n110 10.6151
R962 B.n386 B.n385 10.6151
R963 B.n387 B.n386 10.6151
R964 B.n387 B.n102 10.6151
R965 B.n397 B.n102 10.6151
R966 B.n398 B.n397 10.6151
R967 B.n400 B.n398 10.6151
R968 B.n400 B.n399 10.6151
R969 B.n399 B.n94 10.6151
R970 B.n411 B.n94 10.6151
R971 B.n412 B.n411 10.6151
R972 B.n413 B.n412 10.6151
R973 B.n414 B.n413 10.6151
R974 B.n415 B.n414 10.6151
R975 B.n418 B.n415 10.6151
R976 B.n419 B.n418 10.6151
R977 B.n420 B.n419 10.6151
R978 B.n421 B.n420 10.6151
R979 B.n423 B.n421 10.6151
R980 B.n424 B.n423 10.6151
R981 B.n425 B.n424 10.6151
R982 B.n426 B.n425 10.6151
R983 B.n428 B.n426 10.6151
R984 B.n429 B.n428 10.6151
R985 B.n430 B.n429 10.6151
R986 B.n431 B.n430 10.6151
R987 B.n433 B.n431 10.6151
R988 B.n434 B.n433 10.6151
R989 B.n435 B.n434 10.6151
R990 B.n436 B.n435 10.6151
R991 B.n438 B.n436 10.6151
R992 B.n439 B.n438 10.6151
R993 B.n440 B.n439 10.6151
R994 B.n441 B.n440 10.6151
R995 B.n443 B.n441 10.6151
R996 B.n444 B.n443 10.6151
R997 B.n445 B.n444 10.6151
R998 B.n446 B.n445 10.6151
R999 B.n644 B.n1 10.6151
R1000 B.n644 B.n643 10.6151
R1001 B.n643 B.n642 10.6151
R1002 B.n642 B.n10 10.6151
R1003 B.n636 B.n10 10.6151
R1004 B.n636 B.n635 10.6151
R1005 B.n635 B.n634 10.6151
R1006 B.n634 B.n18 10.6151
R1007 B.n628 B.n18 10.6151
R1008 B.n628 B.n627 10.6151
R1009 B.n627 B.n626 10.6151
R1010 B.n626 B.n25 10.6151
R1011 B.n620 B.n25 10.6151
R1012 B.n620 B.n619 10.6151
R1013 B.n619 B.n618 10.6151
R1014 B.n618 B.n32 10.6151
R1015 B.n612 B.n32 10.6151
R1016 B.n612 B.n611 10.6151
R1017 B.n611 B.n610 10.6151
R1018 B.n610 B.n38 10.6151
R1019 B.n604 B.n38 10.6151
R1020 B.n604 B.n603 10.6151
R1021 B.n603 B.n602 10.6151
R1022 B.n602 B.n46 10.6151
R1023 B.n596 B.n46 10.6151
R1024 B.n595 B.n594 10.6151
R1025 B.n594 B.n53 10.6151
R1026 B.n588 B.n53 10.6151
R1027 B.n588 B.n587 10.6151
R1028 B.n587 B.n586 10.6151
R1029 B.n586 B.n55 10.6151
R1030 B.n580 B.n55 10.6151
R1031 B.n580 B.n579 10.6151
R1032 B.n579 B.n578 10.6151
R1033 B.n578 B.n57 10.6151
R1034 B.n572 B.n57 10.6151
R1035 B.n572 B.n571 10.6151
R1036 B.n571 B.n570 10.6151
R1037 B.n570 B.n59 10.6151
R1038 B.n564 B.n59 10.6151
R1039 B.n564 B.n563 10.6151
R1040 B.n563 B.n562 10.6151
R1041 B.n562 B.n61 10.6151
R1042 B.n556 B.n61 10.6151
R1043 B.n556 B.n555 10.6151
R1044 B.n555 B.n554 10.6151
R1045 B.n554 B.n63 10.6151
R1046 B.n548 B.n63 10.6151
R1047 B.n548 B.n547 10.6151
R1048 B.n547 B.n546 10.6151
R1049 B.n546 B.n65 10.6151
R1050 B.n540 B.n65 10.6151
R1051 B.n540 B.n539 10.6151
R1052 B.n539 B.n538 10.6151
R1053 B.n538 B.n67 10.6151
R1054 B.n532 B.n67 10.6151
R1055 B.n530 B.n529 10.6151
R1056 B.n529 B.n71 10.6151
R1057 B.n523 B.n71 10.6151
R1058 B.n523 B.n522 10.6151
R1059 B.n522 B.n521 10.6151
R1060 B.n521 B.n73 10.6151
R1061 B.n515 B.n73 10.6151
R1062 B.n515 B.n514 10.6151
R1063 B.n514 B.n513 10.6151
R1064 B.n509 B.n508 10.6151
R1065 B.n508 B.n79 10.6151
R1066 B.n503 B.n79 10.6151
R1067 B.n503 B.n502 10.6151
R1068 B.n502 B.n501 10.6151
R1069 B.n501 B.n81 10.6151
R1070 B.n495 B.n81 10.6151
R1071 B.n495 B.n494 10.6151
R1072 B.n494 B.n493 10.6151
R1073 B.n493 B.n83 10.6151
R1074 B.n487 B.n83 10.6151
R1075 B.n487 B.n486 10.6151
R1076 B.n486 B.n485 10.6151
R1077 B.n485 B.n85 10.6151
R1078 B.n479 B.n85 10.6151
R1079 B.n479 B.n478 10.6151
R1080 B.n478 B.n477 10.6151
R1081 B.n477 B.n87 10.6151
R1082 B.n471 B.n87 10.6151
R1083 B.n471 B.n470 10.6151
R1084 B.n470 B.n469 10.6151
R1085 B.n469 B.n89 10.6151
R1086 B.n463 B.n89 10.6151
R1087 B.n463 B.n462 10.6151
R1088 B.n462 B.n461 10.6151
R1089 B.n461 B.n91 10.6151
R1090 B.n455 B.n91 10.6151
R1091 B.n455 B.n454 10.6151
R1092 B.n454 B.n453 10.6151
R1093 B.n453 B.n93 10.6151
R1094 B.n447 B.n93 10.6151
R1095 B.n270 B.n269 9.36635
R1096 B.n246 B.n171 9.36635
R1097 B.n532 B.n531 9.36635
R1098 B.n509 B.n77 9.36635
R1099 B.n652 B.n0 8.11757
R1100 B.n652 B.n1 8.11757
R1101 B.n359 B.t10 1.57137
R1102 B.n614 B.t3 1.57137
R1103 B.n269 B.n268 1.24928
R1104 B.n171 B.n167 1.24928
R1105 B.n531 B.n530 1.24928
R1106 B.n513 B.n77 1.24928
R1107 VN VN.t0 159.435
R1108 VN VN.t1 117.209
R1109 VTAIL.n178 VTAIL.n138 289.615
R1110 VTAIL.n40 VTAIL.n0 289.615
R1111 VTAIL.n132 VTAIL.n92 289.615
R1112 VTAIL.n86 VTAIL.n46 289.615
R1113 VTAIL.n153 VTAIL.n152 185
R1114 VTAIL.n150 VTAIL.n149 185
R1115 VTAIL.n159 VTAIL.n158 185
R1116 VTAIL.n161 VTAIL.n160 185
R1117 VTAIL.n146 VTAIL.n145 185
R1118 VTAIL.n167 VTAIL.n166 185
R1119 VTAIL.n170 VTAIL.n169 185
R1120 VTAIL.n168 VTAIL.n142 185
R1121 VTAIL.n175 VTAIL.n141 185
R1122 VTAIL.n177 VTAIL.n176 185
R1123 VTAIL.n179 VTAIL.n178 185
R1124 VTAIL.n15 VTAIL.n14 185
R1125 VTAIL.n12 VTAIL.n11 185
R1126 VTAIL.n21 VTAIL.n20 185
R1127 VTAIL.n23 VTAIL.n22 185
R1128 VTAIL.n8 VTAIL.n7 185
R1129 VTAIL.n29 VTAIL.n28 185
R1130 VTAIL.n32 VTAIL.n31 185
R1131 VTAIL.n30 VTAIL.n4 185
R1132 VTAIL.n37 VTAIL.n3 185
R1133 VTAIL.n39 VTAIL.n38 185
R1134 VTAIL.n41 VTAIL.n40 185
R1135 VTAIL.n133 VTAIL.n132 185
R1136 VTAIL.n131 VTAIL.n130 185
R1137 VTAIL.n129 VTAIL.n95 185
R1138 VTAIL.n99 VTAIL.n96 185
R1139 VTAIL.n124 VTAIL.n123 185
R1140 VTAIL.n122 VTAIL.n121 185
R1141 VTAIL.n101 VTAIL.n100 185
R1142 VTAIL.n116 VTAIL.n115 185
R1143 VTAIL.n114 VTAIL.n113 185
R1144 VTAIL.n105 VTAIL.n104 185
R1145 VTAIL.n108 VTAIL.n107 185
R1146 VTAIL.n87 VTAIL.n86 185
R1147 VTAIL.n85 VTAIL.n84 185
R1148 VTAIL.n83 VTAIL.n49 185
R1149 VTAIL.n53 VTAIL.n50 185
R1150 VTAIL.n78 VTAIL.n77 185
R1151 VTAIL.n76 VTAIL.n75 185
R1152 VTAIL.n55 VTAIL.n54 185
R1153 VTAIL.n70 VTAIL.n69 185
R1154 VTAIL.n68 VTAIL.n67 185
R1155 VTAIL.n59 VTAIL.n58 185
R1156 VTAIL.n62 VTAIL.n61 185
R1157 VTAIL.t2 VTAIL.n151 149.524
R1158 VTAIL.t1 VTAIL.n13 149.524
R1159 VTAIL.t0 VTAIL.n106 149.524
R1160 VTAIL.t3 VTAIL.n60 149.524
R1161 VTAIL.n152 VTAIL.n149 104.615
R1162 VTAIL.n159 VTAIL.n149 104.615
R1163 VTAIL.n160 VTAIL.n159 104.615
R1164 VTAIL.n160 VTAIL.n145 104.615
R1165 VTAIL.n167 VTAIL.n145 104.615
R1166 VTAIL.n169 VTAIL.n167 104.615
R1167 VTAIL.n169 VTAIL.n168 104.615
R1168 VTAIL.n168 VTAIL.n141 104.615
R1169 VTAIL.n177 VTAIL.n141 104.615
R1170 VTAIL.n178 VTAIL.n177 104.615
R1171 VTAIL.n14 VTAIL.n11 104.615
R1172 VTAIL.n21 VTAIL.n11 104.615
R1173 VTAIL.n22 VTAIL.n21 104.615
R1174 VTAIL.n22 VTAIL.n7 104.615
R1175 VTAIL.n29 VTAIL.n7 104.615
R1176 VTAIL.n31 VTAIL.n29 104.615
R1177 VTAIL.n31 VTAIL.n30 104.615
R1178 VTAIL.n30 VTAIL.n3 104.615
R1179 VTAIL.n39 VTAIL.n3 104.615
R1180 VTAIL.n40 VTAIL.n39 104.615
R1181 VTAIL.n132 VTAIL.n131 104.615
R1182 VTAIL.n131 VTAIL.n95 104.615
R1183 VTAIL.n99 VTAIL.n95 104.615
R1184 VTAIL.n123 VTAIL.n99 104.615
R1185 VTAIL.n123 VTAIL.n122 104.615
R1186 VTAIL.n122 VTAIL.n100 104.615
R1187 VTAIL.n115 VTAIL.n100 104.615
R1188 VTAIL.n115 VTAIL.n114 104.615
R1189 VTAIL.n114 VTAIL.n104 104.615
R1190 VTAIL.n107 VTAIL.n104 104.615
R1191 VTAIL.n86 VTAIL.n85 104.615
R1192 VTAIL.n85 VTAIL.n49 104.615
R1193 VTAIL.n53 VTAIL.n49 104.615
R1194 VTAIL.n77 VTAIL.n53 104.615
R1195 VTAIL.n77 VTAIL.n76 104.615
R1196 VTAIL.n76 VTAIL.n54 104.615
R1197 VTAIL.n69 VTAIL.n54 104.615
R1198 VTAIL.n69 VTAIL.n68 104.615
R1199 VTAIL.n68 VTAIL.n58 104.615
R1200 VTAIL.n61 VTAIL.n58 104.615
R1201 VTAIL.n152 VTAIL.t2 52.3082
R1202 VTAIL.n14 VTAIL.t1 52.3082
R1203 VTAIL.n107 VTAIL.t0 52.3082
R1204 VTAIL.n61 VTAIL.t3 52.3082
R1205 VTAIL.n183 VTAIL.n182 36.2581
R1206 VTAIL.n45 VTAIL.n44 36.2581
R1207 VTAIL.n137 VTAIL.n136 36.2581
R1208 VTAIL.n91 VTAIL.n90 36.2581
R1209 VTAIL.n91 VTAIL.n45 25.2548
R1210 VTAIL.n183 VTAIL.n137 22.5738
R1211 VTAIL.n176 VTAIL.n175 13.1884
R1212 VTAIL.n38 VTAIL.n37 13.1884
R1213 VTAIL.n130 VTAIL.n129 13.1884
R1214 VTAIL.n84 VTAIL.n83 13.1884
R1215 VTAIL.n174 VTAIL.n142 12.8005
R1216 VTAIL.n179 VTAIL.n140 12.8005
R1217 VTAIL.n36 VTAIL.n4 12.8005
R1218 VTAIL.n41 VTAIL.n2 12.8005
R1219 VTAIL.n133 VTAIL.n94 12.8005
R1220 VTAIL.n128 VTAIL.n96 12.8005
R1221 VTAIL.n87 VTAIL.n48 12.8005
R1222 VTAIL.n82 VTAIL.n50 12.8005
R1223 VTAIL.n171 VTAIL.n170 12.0247
R1224 VTAIL.n180 VTAIL.n138 12.0247
R1225 VTAIL.n33 VTAIL.n32 12.0247
R1226 VTAIL.n42 VTAIL.n0 12.0247
R1227 VTAIL.n134 VTAIL.n92 12.0247
R1228 VTAIL.n125 VTAIL.n124 12.0247
R1229 VTAIL.n88 VTAIL.n46 12.0247
R1230 VTAIL.n79 VTAIL.n78 12.0247
R1231 VTAIL.n166 VTAIL.n144 11.249
R1232 VTAIL.n28 VTAIL.n6 11.249
R1233 VTAIL.n121 VTAIL.n98 11.249
R1234 VTAIL.n75 VTAIL.n52 11.249
R1235 VTAIL.n165 VTAIL.n146 10.4732
R1236 VTAIL.n27 VTAIL.n8 10.4732
R1237 VTAIL.n120 VTAIL.n101 10.4732
R1238 VTAIL.n74 VTAIL.n55 10.4732
R1239 VTAIL.n153 VTAIL.n151 10.2747
R1240 VTAIL.n15 VTAIL.n13 10.2747
R1241 VTAIL.n108 VTAIL.n106 10.2747
R1242 VTAIL.n62 VTAIL.n60 10.2747
R1243 VTAIL.n162 VTAIL.n161 9.69747
R1244 VTAIL.n24 VTAIL.n23 9.69747
R1245 VTAIL.n117 VTAIL.n116 9.69747
R1246 VTAIL.n71 VTAIL.n70 9.69747
R1247 VTAIL.n182 VTAIL.n181 9.45567
R1248 VTAIL.n44 VTAIL.n43 9.45567
R1249 VTAIL.n136 VTAIL.n135 9.45567
R1250 VTAIL.n90 VTAIL.n89 9.45567
R1251 VTAIL.n181 VTAIL.n180 9.3005
R1252 VTAIL.n140 VTAIL.n139 9.3005
R1253 VTAIL.n155 VTAIL.n154 9.3005
R1254 VTAIL.n157 VTAIL.n156 9.3005
R1255 VTAIL.n148 VTAIL.n147 9.3005
R1256 VTAIL.n163 VTAIL.n162 9.3005
R1257 VTAIL.n165 VTAIL.n164 9.3005
R1258 VTAIL.n144 VTAIL.n143 9.3005
R1259 VTAIL.n172 VTAIL.n171 9.3005
R1260 VTAIL.n174 VTAIL.n173 9.3005
R1261 VTAIL.n43 VTAIL.n42 9.3005
R1262 VTAIL.n2 VTAIL.n1 9.3005
R1263 VTAIL.n17 VTAIL.n16 9.3005
R1264 VTAIL.n19 VTAIL.n18 9.3005
R1265 VTAIL.n10 VTAIL.n9 9.3005
R1266 VTAIL.n25 VTAIL.n24 9.3005
R1267 VTAIL.n27 VTAIL.n26 9.3005
R1268 VTAIL.n6 VTAIL.n5 9.3005
R1269 VTAIL.n34 VTAIL.n33 9.3005
R1270 VTAIL.n36 VTAIL.n35 9.3005
R1271 VTAIL.n110 VTAIL.n109 9.3005
R1272 VTAIL.n112 VTAIL.n111 9.3005
R1273 VTAIL.n103 VTAIL.n102 9.3005
R1274 VTAIL.n118 VTAIL.n117 9.3005
R1275 VTAIL.n120 VTAIL.n119 9.3005
R1276 VTAIL.n98 VTAIL.n97 9.3005
R1277 VTAIL.n126 VTAIL.n125 9.3005
R1278 VTAIL.n128 VTAIL.n127 9.3005
R1279 VTAIL.n135 VTAIL.n134 9.3005
R1280 VTAIL.n94 VTAIL.n93 9.3005
R1281 VTAIL.n64 VTAIL.n63 9.3005
R1282 VTAIL.n66 VTAIL.n65 9.3005
R1283 VTAIL.n57 VTAIL.n56 9.3005
R1284 VTAIL.n72 VTAIL.n71 9.3005
R1285 VTAIL.n74 VTAIL.n73 9.3005
R1286 VTAIL.n52 VTAIL.n51 9.3005
R1287 VTAIL.n80 VTAIL.n79 9.3005
R1288 VTAIL.n82 VTAIL.n81 9.3005
R1289 VTAIL.n89 VTAIL.n88 9.3005
R1290 VTAIL.n48 VTAIL.n47 9.3005
R1291 VTAIL.n158 VTAIL.n148 8.92171
R1292 VTAIL.n20 VTAIL.n10 8.92171
R1293 VTAIL.n113 VTAIL.n103 8.92171
R1294 VTAIL.n67 VTAIL.n57 8.92171
R1295 VTAIL.n157 VTAIL.n150 8.14595
R1296 VTAIL.n19 VTAIL.n12 8.14595
R1297 VTAIL.n112 VTAIL.n105 8.14595
R1298 VTAIL.n66 VTAIL.n59 8.14595
R1299 VTAIL.n154 VTAIL.n153 7.3702
R1300 VTAIL.n16 VTAIL.n15 7.3702
R1301 VTAIL.n109 VTAIL.n108 7.3702
R1302 VTAIL.n63 VTAIL.n62 7.3702
R1303 VTAIL.n154 VTAIL.n150 5.81868
R1304 VTAIL.n16 VTAIL.n12 5.81868
R1305 VTAIL.n109 VTAIL.n105 5.81868
R1306 VTAIL.n63 VTAIL.n59 5.81868
R1307 VTAIL.n158 VTAIL.n157 5.04292
R1308 VTAIL.n20 VTAIL.n19 5.04292
R1309 VTAIL.n113 VTAIL.n112 5.04292
R1310 VTAIL.n67 VTAIL.n66 5.04292
R1311 VTAIL.n161 VTAIL.n148 4.26717
R1312 VTAIL.n23 VTAIL.n10 4.26717
R1313 VTAIL.n116 VTAIL.n103 4.26717
R1314 VTAIL.n70 VTAIL.n57 4.26717
R1315 VTAIL.n162 VTAIL.n146 3.49141
R1316 VTAIL.n24 VTAIL.n8 3.49141
R1317 VTAIL.n117 VTAIL.n101 3.49141
R1318 VTAIL.n71 VTAIL.n55 3.49141
R1319 VTAIL.n155 VTAIL.n151 2.84303
R1320 VTAIL.n17 VTAIL.n13 2.84303
R1321 VTAIL.n110 VTAIL.n106 2.84303
R1322 VTAIL.n64 VTAIL.n60 2.84303
R1323 VTAIL.n166 VTAIL.n165 2.71565
R1324 VTAIL.n28 VTAIL.n27 2.71565
R1325 VTAIL.n121 VTAIL.n120 2.71565
R1326 VTAIL.n75 VTAIL.n74 2.71565
R1327 VTAIL.n170 VTAIL.n144 1.93989
R1328 VTAIL.n182 VTAIL.n138 1.93989
R1329 VTAIL.n32 VTAIL.n6 1.93989
R1330 VTAIL.n44 VTAIL.n0 1.93989
R1331 VTAIL.n136 VTAIL.n92 1.93989
R1332 VTAIL.n124 VTAIL.n98 1.93989
R1333 VTAIL.n90 VTAIL.n46 1.93989
R1334 VTAIL.n78 VTAIL.n52 1.93989
R1335 VTAIL.n137 VTAIL.n91 1.81084
R1336 VTAIL VTAIL.n45 1.19878
R1337 VTAIL.n171 VTAIL.n142 1.16414
R1338 VTAIL.n180 VTAIL.n179 1.16414
R1339 VTAIL.n33 VTAIL.n4 1.16414
R1340 VTAIL.n42 VTAIL.n41 1.16414
R1341 VTAIL.n134 VTAIL.n133 1.16414
R1342 VTAIL.n125 VTAIL.n96 1.16414
R1343 VTAIL.n88 VTAIL.n87 1.16414
R1344 VTAIL.n79 VTAIL.n50 1.16414
R1345 VTAIL VTAIL.n183 0.612569
R1346 VTAIL.n175 VTAIL.n174 0.388379
R1347 VTAIL.n176 VTAIL.n140 0.388379
R1348 VTAIL.n37 VTAIL.n36 0.388379
R1349 VTAIL.n38 VTAIL.n2 0.388379
R1350 VTAIL.n130 VTAIL.n94 0.388379
R1351 VTAIL.n129 VTAIL.n128 0.388379
R1352 VTAIL.n84 VTAIL.n48 0.388379
R1353 VTAIL.n83 VTAIL.n82 0.388379
R1354 VTAIL.n156 VTAIL.n155 0.155672
R1355 VTAIL.n156 VTAIL.n147 0.155672
R1356 VTAIL.n163 VTAIL.n147 0.155672
R1357 VTAIL.n164 VTAIL.n163 0.155672
R1358 VTAIL.n164 VTAIL.n143 0.155672
R1359 VTAIL.n172 VTAIL.n143 0.155672
R1360 VTAIL.n173 VTAIL.n172 0.155672
R1361 VTAIL.n173 VTAIL.n139 0.155672
R1362 VTAIL.n181 VTAIL.n139 0.155672
R1363 VTAIL.n18 VTAIL.n17 0.155672
R1364 VTAIL.n18 VTAIL.n9 0.155672
R1365 VTAIL.n25 VTAIL.n9 0.155672
R1366 VTAIL.n26 VTAIL.n25 0.155672
R1367 VTAIL.n26 VTAIL.n5 0.155672
R1368 VTAIL.n34 VTAIL.n5 0.155672
R1369 VTAIL.n35 VTAIL.n34 0.155672
R1370 VTAIL.n35 VTAIL.n1 0.155672
R1371 VTAIL.n43 VTAIL.n1 0.155672
R1372 VTAIL.n135 VTAIL.n93 0.155672
R1373 VTAIL.n127 VTAIL.n93 0.155672
R1374 VTAIL.n127 VTAIL.n126 0.155672
R1375 VTAIL.n126 VTAIL.n97 0.155672
R1376 VTAIL.n119 VTAIL.n97 0.155672
R1377 VTAIL.n119 VTAIL.n118 0.155672
R1378 VTAIL.n118 VTAIL.n102 0.155672
R1379 VTAIL.n111 VTAIL.n102 0.155672
R1380 VTAIL.n111 VTAIL.n110 0.155672
R1381 VTAIL.n89 VTAIL.n47 0.155672
R1382 VTAIL.n81 VTAIL.n47 0.155672
R1383 VTAIL.n81 VTAIL.n80 0.155672
R1384 VTAIL.n80 VTAIL.n51 0.155672
R1385 VTAIL.n73 VTAIL.n51 0.155672
R1386 VTAIL.n73 VTAIL.n72 0.155672
R1387 VTAIL.n72 VTAIL.n56 0.155672
R1388 VTAIL.n65 VTAIL.n56 0.155672
R1389 VTAIL.n65 VTAIL.n64 0.155672
R1390 VDD2.n85 VDD2.n45 289.615
R1391 VDD2.n40 VDD2.n0 289.615
R1392 VDD2.n86 VDD2.n85 185
R1393 VDD2.n84 VDD2.n83 185
R1394 VDD2.n82 VDD2.n48 185
R1395 VDD2.n52 VDD2.n49 185
R1396 VDD2.n77 VDD2.n76 185
R1397 VDD2.n75 VDD2.n74 185
R1398 VDD2.n54 VDD2.n53 185
R1399 VDD2.n69 VDD2.n68 185
R1400 VDD2.n67 VDD2.n66 185
R1401 VDD2.n58 VDD2.n57 185
R1402 VDD2.n61 VDD2.n60 185
R1403 VDD2.n15 VDD2.n14 185
R1404 VDD2.n12 VDD2.n11 185
R1405 VDD2.n21 VDD2.n20 185
R1406 VDD2.n23 VDD2.n22 185
R1407 VDD2.n8 VDD2.n7 185
R1408 VDD2.n29 VDD2.n28 185
R1409 VDD2.n32 VDD2.n31 185
R1410 VDD2.n30 VDD2.n4 185
R1411 VDD2.n37 VDD2.n3 185
R1412 VDD2.n39 VDD2.n38 185
R1413 VDD2.n41 VDD2.n40 185
R1414 VDD2.t1 VDD2.n59 149.524
R1415 VDD2.t0 VDD2.n13 149.524
R1416 VDD2.n85 VDD2.n84 104.615
R1417 VDD2.n84 VDD2.n48 104.615
R1418 VDD2.n52 VDD2.n48 104.615
R1419 VDD2.n76 VDD2.n52 104.615
R1420 VDD2.n76 VDD2.n75 104.615
R1421 VDD2.n75 VDD2.n53 104.615
R1422 VDD2.n68 VDD2.n53 104.615
R1423 VDD2.n68 VDD2.n67 104.615
R1424 VDD2.n67 VDD2.n57 104.615
R1425 VDD2.n60 VDD2.n57 104.615
R1426 VDD2.n14 VDD2.n11 104.615
R1427 VDD2.n21 VDD2.n11 104.615
R1428 VDD2.n22 VDD2.n21 104.615
R1429 VDD2.n22 VDD2.n7 104.615
R1430 VDD2.n29 VDD2.n7 104.615
R1431 VDD2.n31 VDD2.n29 104.615
R1432 VDD2.n31 VDD2.n30 104.615
R1433 VDD2.n30 VDD2.n3 104.615
R1434 VDD2.n39 VDD2.n3 104.615
R1435 VDD2.n40 VDD2.n39 104.615
R1436 VDD2.n90 VDD2.n44 89.4842
R1437 VDD2.n90 VDD2.n89 52.9369
R1438 VDD2.n60 VDD2.t1 52.3082
R1439 VDD2.n14 VDD2.t0 52.3082
R1440 VDD2.n83 VDD2.n82 13.1884
R1441 VDD2.n38 VDD2.n37 13.1884
R1442 VDD2.n86 VDD2.n47 12.8005
R1443 VDD2.n81 VDD2.n49 12.8005
R1444 VDD2.n36 VDD2.n4 12.8005
R1445 VDD2.n41 VDD2.n2 12.8005
R1446 VDD2.n87 VDD2.n45 12.0247
R1447 VDD2.n78 VDD2.n77 12.0247
R1448 VDD2.n33 VDD2.n32 12.0247
R1449 VDD2.n42 VDD2.n0 12.0247
R1450 VDD2.n74 VDD2.n51 11.249
R1451 VDD2.n28 VDD2.n6 11.249
R1452 VDD2.n73 VDD2.n54 10.4732
R1453 VDD2.n27 VDD2.n8 10.4732
R1454 VDD2.n61 VDD2.n59 10.2747
R1455 VDD2.n15 VDD2.n13 10.2747
R1456 VDD2.n70 VDD2.n69 9.69747
R1457 VDD2.n24 VDD2.n23 9.69747
R1458 VDD2.n89 VDD2.n88 9.45567
R1459 VDD2.n44 VDD2.n43 9.45567
R1460 VDD2.n63 VDD2.n62 9.3005
R1461 VDD2.n65 VDD2.n64 9.3005
R1462 VDD2.n56 VDD2.n55 9.3005
R1463 VDD2.n71 VDD2.n70 9.3005
R1464 VDD2.n73 VDD2.n72 9.3005
R1465 VDD2.n51 VDD2.n50 9.3005
R1466 VDD2.n79 VDD2.n78 9.3005
R1467 VDD2.n81 VDD2.n80 9.3005
R1468 VDD2.n88 VDD2.n87 9.3005
R1469 VDD2.n47 VDD2.n46 9.3005
R1470 VDD2.n43 VDD2.n42 9.3005
R1471 VDD2.n2 VDD2.n1 9.3005
R1472 VDD2.n17 VDD2.n16 9.3005
R1473 VDD2.n19 VDD2.n18 9.3005
R1474 VDD2.n10 VDD2.n9 9.3005
R1475 VDD2.n25 VDD2.n24 9.3005
R1476 VDD2.n27 VDD2.n26 9.3005
R1477 VDD2.n6 VDD2.n5 9.3005
R1478 VDD2.n34 VDD2.n33 9.3005
R1479 VDD2.n36 VDD2.n35 9.3005
R1480 VDD2.n66 VDD2.n56 8.92171
R1481 VDD2.n20 VDD2.n10 8.92171
R1482 VDD2.n65 VDD2.n58 8.14595
R1483 VDD2.n19 VDD2.n12 8.14595
R1484 VDD2.n62 VDD2.n61 7.3702
R1485 VDD2.n16 VDD2.n15 7.3702
R1486 VDD2.n62 VDD2.n58 5.81868
R1487 VDD2.n16 VDD2.n12 5.81868
R1488 VDD2.n66 VDD2.n65 5.04292
R1489 VDD2.n20 VDD2.n19 5.04292
R1490 VDD2.n69 VDD2.n56 4.26717
R1491 VDD2.n23 VDD2.n10 4.26717
R1492 VDD2.n70 VDD2.n54 3.49141
R1493 VDD2.n24 VDD2.n8 3.49141
R1494 VDD2.n17 VDD2.n13 2.84303
R1495 VDD2.n63 VDD2.n59 2.84303
R1496 VDD2.n74 VDD2.n73 2.71565
R1497 VDD2.n28 VDD2.n27 2.71565
R1498 VDD2.n89 VDD2.n45 1.93989
R1499 VDD2.n77 VDD2.n51 1.93989
R1500 VDD2.n32 VDD2.n6 1.93989
R1501 VDD2.n44 VDD2.n0 1.93989
R1502 VDD2.n87 VDD2.n86 1.16414
R1503 VDD2.n78 VDD2.n49 1.16414
R1504 VDD2.n33 VDD2.n4 1.16414
R1505 VDD2.n42 VDD2.n41 1.16414
R1506 VDD2 VDD2.n90 0.728948
R1507 VDD2.n83 VDD2.n47 0.388379
R1508 VDD2.n82 VDD2.n81 0.388379
R1509 VDD2.n37 VDD2.n36 0.388379
R1510 VDD2.n38 VDD2.n2 0.388379
R1511 VDD2.n88 VDD2.n46 0.155672
R1512 VDD2.n80 VDD2.n46 0.155672
R1513 VDD2.n80 VDD2.n79 0.155672
R1514 VDD2.n79 VDD2.n50 0.155672
R1515 VDD2.n72 VDD2.n50 0.155672
R1516 VDD2.n72 VDD2.n71 0.155672
R1517 VDD2.n71 VDD2.n55 0.155672
R1518 VDD2.n64 VDD2.n55 0.155672
R1519 VDD2.n64 VDD2.n63 0.155672
R1520 VDD2.n18 VDD2.n17 0.155672
R1521 VDD2.n18 VDD2.n9 0.155672
R1522 VDD2.n25 VDD2.n9 0.155672
R1523 VDD2.n26 VDD2.n25 0.155672
R1524 VDD2.n26 VDD2.n5 0.155672
R1525 VDD2.n34 VDD2.n5 0.155672
R1526 VDD2.n35 VDD2.n34 0.155672
R1527 VDD2.n35 VDD2.n1 0.155672
R1528 VDD2.n43 VDD2.n1 0.155672
R1529 VP.n0 VP.t0 159.435
R1530 VP.n0 VP.t1 116.778
R1531 VP VP.n0 0.431811
R1532 VDD1.n40 VDD1.n0 289.615
R1533 VDD1.n85 VDD1.n45 289.615
R1534 VDD1.n41 VDD1.n40 185
R1535 VDD1.n39 VDD1.n38 185
R1536 VDD1.n37 VDD1.n3 185
R1537 VDD1.n7 VDD1.n4 185
R1538 VDD1.n32 VDD1.n31 185
R1539 VDD1.n30 VDD1.n29 185
R1540 VDD1.n9 VDD1.n8 185
R1541 VDD1.n24 VDD1.n23 185
R1542 VDD1.n22 VDD1.n21 185
R1543 VDD1.n13 VDD1.n12 185
R1544 VDD1.n16 VDD1.n15 185
R1545 VDD1.n60 VDD1.n59 185
R1546 VDD1.n57 VDD1.n56 185
R1547 VDD1.n66 VDD1.n65 185
R1548 VDD1.n68 VDD1.n67 185
R1549 VDD1.n53 VDD1.n52 185
R1550 VDD1.n74 VDD1.n73 185
R1551 VDD1.n77 VDD1.n76 185
R1552 VDD1.n75 VDD1.n49 185
R1553 VDD1.n82 VDD1.n48 185
R1554 VDD1.n84 VDD1.n83 185
R1555 VDD1.n86 VDD1.n85 185
R1556 VDD1.t1 VDD1.n14 149.524
R1557 VDD1.t0 VDD1.n58 149.524
R1558 VDD1.n40 VDD1.n39 104.615
R1559 VDD1.n39 VDD1.n3 104.615
R1560 VDD1.n7 VDD1.n3 104.615
R1561 VDD1.n31 VDD1.n7 104.615
R1562 VDD1.n31 VDD1.n30 104.615
R1563 VDD1.n30 VDD1.n8 104.615
R1564 VDD1.n23 VDD1.n8 104.615
R1565 VDD1.n23 VDD1.n22 104.615
R1566 VDD1.n22 VDD1.n12 104.615
R1567 VDD1.n15 VDD1.n12 104.615
R1568 VDD1.n59 VDD1.n56 104.615
R1569 VDD1.n66 VDD1.n56 104.615
R1570 VDD1.n67 VDD1.n66 104.615
R1571 VDD1.n67 VDD1.n52 104.615
R1572 VDD1.n74 VDD1.n52 104.615
R1573 VDD1.n76 VDD1.n74 104.615
R1574 VDD1.n76 VDD1.n75 104.615
R1575 VDD1.n75 VDD1.n48 104.615
R1576 VDD1.n84 VDD1.n48 104.615
R1577 VDD1.n85 VDD1.n84 104.615
R1578 VDD1 VDD1.n89 90.6793
R1579 VDD1 VDD1.n44 53.6653
R1580 VDD1.n15 VDD1.t1 52.3082
R1581 VDD1.n59 VDD1.t0 52.3082
R1582 VDD1.n38 VDD1.n37 13.1884
R1583 VDD1.n83 VDD1.n82 13.1884
R1584 VDD1.n41 VDD1.n2 12.8005
R1585 VDD1.n36 VDD1.n4 12.8005
R1586 VDD1.n81 VDD1.n49 12.8005
R1587 VDD1.n86 VDD1.n47 12.8005
R1588 VDD1.n42 VDD1.n0 12.0247
R1589 VDD1.n33 VDD1.n32 12.0247
R1590 VDD1.n78 VDD1.n77 12.0247
R1591 VDD1.n87 VDD1.n45 12.0247
R1592 VDD1.n29 VDD1.n6 11.249
R1593 VDD1.n73 VDD1.n51 11.249
R1594 VDD1.n28 VDD1.n9 10.4732
R1595 VDD1.n72 VDD1.n53 10.4732
R1596 VDD1.n16 VDD1.n14 10.2747
R1597 VDD1.n60 VDD1.n58 10.2747
R1598 VDD1.n25 VDD1.n24 9.69747
R1599 VDD1.n69 VDD1.n68 9.69747
R1600 VDD1.n44 VDD1.n43 9.45567
R1601 VDD1.n89 VDD1.n88 9.45567
R1602 VDD1.n18 VDD1.n17 9.3005
R1603 VDD1.n20 VDD1.n19 9.3005
R1604 VDD1.n11 VDD1.n10 9.3005
R1605 VDD1.n26 VDD1.n25 9.3005
R1606 VDD1.n28 VDD1.n27 9.3005
R1607 VDD1.n6 VDD1.n5 9.3005
R1608 VDD1.n34 VDD1.n33 9.3005
R1609 VDD1.n36 VDD1.n35 9.3005
R1610 VDD1.n43 VDD1.n42 9.3005
R1611 VDD1.n2 VDD1.n1 9.3005
R1612 VDD1.n88 VDD1.n87 9.3005
R1613 VDD1.n47 VDD1.n46 9.3005
R1614 VDD1.n62 VDD1.n61 9.3005
R1615 VDD1.n64 VDD1.n63 9.3005
R1616 VDD1.n55 VDD1.n54 9.3005
R1617 VDD1.n70 VDD1.n69 9.3005
R1618 VDD1.n72 VDD1.n71 9.3005
R1619 VDD1.n51 VDD1.n50 9.3005
R1620 VDD1.n79 VDD1.n78 9.3005
R1621 VDD1.n81 VDD1.n80 9.3005
R1622 VDD1.n21 VDD1.n11 8.92171
R1623 VDD1.n65 VDD1.n55 8.92171
R1624 VDD1.n20 VDD1.n13 8.14595
R1625 VDD1.n64 VDD1.n57 8.14595
R1626 VDD1.n17 VDD1.n16 7.3702
R1627 VDD1.n61 VDD1.n60 7.3702
R1628 VDD1.n17 VDD1.n13 5.81868
R1629 VDD1.n61 VDD1.n57 5.81868
R1630 VDD1.n21 VDD1.n20 5.04292
R1631 VDD1.n65 VDD1.n64 5.04292
R1632 VDD1.n24 VDD1.n11 4.26717
R1633 VDD1.n68 VDD1.n55 4.26717
R1634 VDD1.n25 VDD1.n9 3.49141
R1635 VDD1.n69 VDD1.n53 3.49141
R1636 VDD1.n62 VDD1.n58 2.84303
R1637 VDD1.n18 VDD1.n14 2.84303
R1638 VDD1.n29 VDD1.n28 2.71565
R1639 VDD1.n73 VDD1.n72 2.71565
R1640 VDD1.n44 VDD1.n0 1.93989
R1641 VDD1.n32 VDD1.n6 1.93989
R1642 VDD1.n77 VDD1.n51 1.93989
R1643 VDD1.n89 VDD1.n45 1.93989
R1644 VDD1.n42 VDD1.n41 1.16414
R1645 VDD1.n33 VDD1.n4 1.16414
R1646 VDD1.n78 VDD1.n49 1.16414
R1647 VDD1.n87 VDD1.n86 1.16414
R1648 VDD1.n38 VDD1.n2 0.388379
R1649 VDD1.n37 VDD1.n36 0.388379
R1650 VDD1.n82 VDD1.n81 0.388379
R1651 VDD1.n83 VDD1.n47 0.388379
R1652 VDD1.n43 VDD1.n1 0.155672
R1653 VDD1.n35 VDD1.n1 0.155672
R1654 VDD1.n35 VDD1.n34 0.155672
R1655 VDD1.n34 VDD1.n5 0.155672
R1656 VDD1.n27 VDD1.n5 0.155672
R1657 VDD1.n27 VDD1.n26 0.155672
R1658 VDD1.n26 VDD1.n10 0.155672
R1659 VDD1.n19 VDD1.n10 0.155672
R1660 VDD1.n19 VDD1.n18 0.155672
R1661 VDD1.n63 VDD1.n62 0.155672
R1662 VDD1.n63 VDD1.n54 0.155672
R1663 VDD1.n70 VDD1.n54 0.155672
R1664 VDD1.n71 VDD1.n70 0.155672
R1665 VDD1.n71 VDD1.n50 0.155672
R1666 VDD1.n79 VDD1.n50 0.155672
R1667 VDD1.n80 VDD1.n79 0.155672
R1668 VDD1.n80 VDD1.n46 0.155672
R1669 VDD1.n88 VDD1.n46 0.155672
C0 VP VDD2 0.340375f
C1 VDD1 VTAIL 4.24009f
C2 VP VN 4.93655f
C3 VDD1 VDD2 0.696006f
C4 VTAIL VDD2 4.29281f
C5 VDD1 VN 0.148205f
C6 VN VTAIL 1.93999f
C7 VN VDD2 2.1105f
C8 VDD1 VP 2.30076f
C9 VP VTAIL 1.95422f
C10 VDD2 B 3.90835f
C11 VDD1 B 6.45324f
C12 VTAIL B 6.08107f
C13 VN B 9.32488f
C14 VP B 6.393656f
C15 VDD1.n0 B 0.029205f
C16 VDD1.n1 B 0.020678f
C17 VDD1.n2 B 0.011112f
C18 VDD1.n3 B 0.026264f
C19 VDD1.n4 B 0.011765f
C20 VDD1.n5 B 0.020678f
C21 VDD1.n6 B 0.011112f
C22 VDD1.n7 B 0.026264f
C23 VDD1.n8 B 0.026264f
C24 VDD1.n9 B 0.011765f
C25 VDD1.n10 B 0.020678f
C26 VDD1.n11 B 0.011112f
C27 VDD1.n12 B 0.026264f
C28 VDD1.n13 B 0.011765f
C29 VDD1.n14 B 0.123143f
C30 VDD1.t1 B 0.044002f
C31 VDD1.n15 B 0.019698f
C32 VDD1.n16 B 0.018566f
C33 VDD1.n17 B 0.011112f
C34 VDD1.n18 B 0.742404f
C35 VDD1.n19 B 0.020678f
C36 VDD1.n20 B 0.011112f
C37 VDD1.n21 B 0.011765f
C38 VDD1.n22 B 0.026264f
C39 VDD1.n23 B 0.026264f
C40 VDD1.n24 B 0.011765f
C41 VDD1.n25 B 0.011112f
C42 VDD1.n26 B 0.020678f
C43 VDD1.n27 B 0.020678f
C44 VDD1.n28 B 0.011112f
C45 VDD1.n29 B 0.011765f
C46 VDD1.n30 B 0.026264f
C47 VDD1.n31 B 0.026264f
C48 VDD1.n32 B 0.011765f
C49 VDD1.n33 B 0.011112f
C50 VDD1.n34 B 0.020678f
C51 VDD1.n35 B 0.020678f
C52 VDD1.n36 B 0.011112f
C53 VDD1.n37 B 0.011438f
C54 VDD1.n38 B 0.011438f
C55 VDD1.n39 B 0.026264f
C56 VDD1.n40 B 0.057103f
C57 VDD1.n41 B 0.011765f
C58 VDD1.n42 B 0.011112f
C59 VDD1.n43 B 0.053729f
C60 VDD1.n44 B 0.047633f
C61 VDD1.n45 B 0.029205f
C62 VDD1.n46 B 0.020678f
C63 VDD1.n47 B 0.011112f
C64 VDD1.n48 B 0.026264f
C65 VDD1.n49 B 0.011765f
C66 VDD1.n50 B 0.020678f
C67 VDD1.n51 B 0.011112f
C68 VDD1.n52 B 0.026264f
C69 VDD1.n53 B 0.011765f
C70 VDD1.n54 B 0.020678f
C71 VDD1.n55 B 0.011112f
C72 VDD1.n56 B 0.026264f
C73 VDD1.n57 B 0.011765f
C74 VDD1.n58 B 0.123143f
C75 VDD1.t0 B 0.044002f
C76 VDD1.n59 B 0.019698f
C77 VDD1.n60 B 0.018566f
C78 VDD1.n61 B 0.011112f
C79 VDD1.n62 B 0.742404f
C80 VDD1.n63 B 0.020678f
C81 VDD1.n64 B 0.011112f
C82 VDD1.n65 B 0.011765f
C83 VDD1.n66 B 0.026264f
C84 VDD1.n67 B 0.026264f
C85 VDD1.n68 B 0.011765f
C86 VDD1.n69 B 0.011112f
C87 VDD1.n70 B 0.020678f
C88 VDD1.n71 B 0.020678f
C89 VDD1.n72 B 0.011112f
C90 VDD1.n73 B 0.011765f
C91 VDD1.n74 B 0.026264f
C92 VDD1.n75 B 0.026264f
C93 VDD1.n76 B 0.026264f
C94 VDD1.n77 B 0.011765f
C95 VDD1.n78 B 0.011112f
C96 VDD1.n79 B 0.020678f
C97 VDD1.n80 B 0.020678f
C98 VDD1.n81 B 0.011112f
C99 VDD1.n82 B 0.011438f
C100 VDD1.n83 B 0.011438f
C101 VDD1.n84 B 0.026264f
C102 VDD1.n85 B 0.057103f
C103 VDD1.n86 B 0.011765f
C104 VDD1.n87 B 0.011112f
C105 VDD1.n88 B 0.053729f
C106 VDD1.n89 B 0.542249f
C107 VP.t1 B 1.90318f
C108 VP.t0 B 2.35436f
C109 VP.n0 B 2.8738f
C110 VDD2.n0 B 0.029097f
C111 VDD2.n1 B 0.020602f
C112 VDD2.n2 B 0.011071f
C113 VDD2.n3 B 0.026167f
C114 VDD2.n4 B 0.011722f
C115 VDD2.n5 B 0.020602f
C116 VDD2.n6 B 0.011071f
C117 VDD2.n7 B 0.026167f
C118 VDD2.n8 B 0.011722f
C119 VDD2.n9 B 0.020602f
C120 VDD2.n10 B 0.011071f
C121 VDD2.n11 B 0.026167f
C122 VDD2.n12 B 0.011722f
C123 VDD2.n13 B 0.122691f
C124 VDD2.t0 B 0.043841f
C125 VDD2.n14 B 0.019625f
C126 VDD2.n15 B 0.018498f
C127 VDD2.n16 B 0.011071f
C128 VDD2.n17 B 0.739673f
C129 VDD2.n18 B 0.020602f
C130 VDD2.n19 B 0.011071f
C131 VDD2.n20 B 0.011722f
C132 VDD2.n21 B 0.026167f
C133 VDD2.n22 B 0.026167f
C134 VDD2.n23 B 0.011722f
C135 VDD2.n24 B 0.011071f
C136 VDD2.n25 B 0.020602f
C137 VDD2.n26 B 0.020602f
C138 VDD2.n27 B 0.011071f
C139 VDD2.n28 B 0.011722f
C140 VDD2.n29 B 0.026167f
C141 VDD2.n30 B 0.026167f
C142 VDD2.n31 B 0.026167f
C143 VDD2.n32 B 0.011722f
C144 VDD2.n33 B 0.011071f
C145 VDD2.n34 B 0.020602f
C146 VDD2.n35 B 0.020602f
C147 VDD2.n36 B 0.011071f
C148 VDD2.n37 B 0.011396f
C149 VDD2.n38 B 0.011396f
C150 VDD2.n39 B 0.026167f
C151 VDD2.n40 B 0.056893f
C152 VDD2.n41 B 0.011722f
C153 VDD2.n42 B 0.011071f
C154 VDD2.n43 B 0.053531f
C155 VDD2.n44 B 0.502441f
C156 VDD2.n45 B 0.029097f
C157 VDD2.n46 B 0.020602f
C158 VDD2.n47 B 0.011071f
C159 VDD2.n48 B 0.026167f
C160 VDD2.n49 B 0.011722f
C161 VDD2.n50 B 0.020602f
C162 VDD2.n51 B 0.011071f
C163 VDD2.n52 B 0.026167f
C164 VDD2.n53 B 0.026167f
C165 VDD2.n54 B 0.011722f
C166 VDD2.n55 B 0.020602f
C167 VDD2.n56 B 0.011071f
C168 VDD2.n57 B 0.026167f
C169 VDD2.n58 B 0.011722f
C170 VDD2.n59 B 0.122691f
C171 VDD2.t1 B 0.043841f
C172 VDD2.n60 B 0.019625f
C173 VDD2.n61 B 0.018498f
C174 VDD2.n62 B 0.011071f
C175 VDD2.n63 B 0.739673f
C176 VDD2.n64 B 0.020602f
C177 VDD2.n65 B 0.011071f
C178 VDD2.n66 B 0.011722f
C179 VDD2.n67 B 0.026167f
C180 VDD2.n68 B 0.026167f
C181 VDD2.n69 B 0.011722f
C182 VDD2.n70 B 0.011071f
C183 VDD2.n71 B 0.020602f
C184 VDD2.n72 B 0.020602f
C185 VDD2.n73 B 0.011071f
C186 VDD2.n74 B 0.011722f
C187 VDD2.n75 B 0.026167f
C188 VDD2.n76 B 0.026167f
C189 VDD2.n77 B 0.011722f
C190 VDD2.n78 B 0.011071f
C191 VDD2.n79 B 0.020602f
C192 VDD2.n80 B 0.020602f
C193 VDD2.n81 B 0.011071f
C194 VDD2.n82 B 0.011396f
C195 VDD2.n83 B 0.011396f
C196 VDD2.n84 B 0.026167f
C197 VDD2.n85 B 0.056893f
C198 VDD2.n86 B 0.011722f
C199 VDD2.n87 B 0.011071f
C200 VDD2.n88 B 0.053531f
C201 VDD2.n89 B 0.046216f
C202 VDD2.n90 B 2.29053f
C203 VTAIL.n0 B 0.021096f
C204 VTAIL.n1 B 0.014937f
C205 VTAIL.n2 B 0.008026f
C206 VTAIL.n3 B 0.018971f
C207 VTAIL.n4 B 0.008498f
C208 VTAIL.n5 B 0.014937f
C209 VTAIL.n6 B 0.008026f
C210 VTAIL.n7 B 0.018971f
C211 VTAIL.n8 B 0.008498f
C212 VTAIL.n9 B 0.014937f
C213 VTAIL.n10 B 0.008026f
C214 VTAIL.n11 B 0.018971f
C215 VTAIL.n12 B 0.008498f
C216 VTAIL.n13 B 0.088951f
C217 VTAIL.t1 B 0.031784f
C218 VTAIL.n14 B 0.014228f
C219 VTAIL.n15 B 0.013411f
C220 VTAIL.n16 B 0.008026f
C221 VTAIL.n17 B 0.536264f
C222 VTAIL.n18 B 0.014937f
C223 VTAIL.n19 B 0.008026f
C224 VTAIL.n20 B 0.008498f
C225 VTAIL.n21 B 0.018971f
C226 VTAIL.n22 B 0.018971f
C227 VTAIL.n23 B 0.008498f
C228 VTAIL.n24 B 0.008026f
C229 VTAIL.n25 B 0.014937f
C230 VTAIL.n26 B 0.014937f
C231 VTAIL.n27 B 0.008026f
C232 VTAIL.n28 B 0.008498f
C233 VTAIL.n29 B 0.018971f
C234 VTAIL.n30 B 0.018971f
C235 VTAIL.n31 B 0.018971f
C236 VTAIL.n32 B 0.008498f
C237 VTAIL.n33 B 0.008026f
C238 VTAIL.n34 B 0.014937f
C239 VTAIL.n35 B 0.014937f
C240 VTAIL.n36 B 0.008026f
C241 VTAIL.n37 B 0.008262f
C242 VTAIL.n38 B 0.008262f
C243 VTAIL.n39 B 0.018971f
C244 VTAIL.n40 B 0.041248f
C245 VTAIL.n41 B 0.008498f
C246 VTAIL.n42 B 0.008026f
C247 VTAIL.n43 B 0.03881f
C248 VTAIL.n44 B 0.023223f
C249 VTAIL.n45 B 0.896035f
C250 VTAIL.n46 B 0.021096f
C251 VTAIL.n47 B 0.014937f
C252 VTAIL.n48 B 0.008026f
C253 VTAIL.n49 B 0.018971f
C254 VTAIL.n50 B 0.008498f
C255 VTAIL.n51 B 0.014937f
C256 VTAIL.n52 B 0.008026f
C257 VTAIL.n53 B 0.018971f
C258 VTAIL.n54 B 0.018971f
C259 VTAIL.n55 B 0.008498f
C260 VTAIL.n56 B 0.014937f
C261 VTAIL.n57 B 0.008026f
C262 VTAIL.n58 B 0.018971f
C263 VTAIL.n59 B 0.008498f
C264 VTAIL.n60 B 0.088951f
C265 VTAIL.t3 B 0.031784f
C266 VTAIL.n61 B 0.014228f
C267 VTAIL.n62 B 0.013411f
C268 VTAIL.n63 B 0.008026f
C269 VTAIL.n64 B 0.536264f
C270 VTAIL.n65 B 0.014937f
C271 VTAIL.n66 B 0.008026f
C272 VTAIL.n67 B 0.008498f
C273 VTAIL.n68 B 0.018971f
C274 VTAIL.n69 B 0.018971f
C275 VTAIL.n70 B 0.008498f
C276 VTAIL.n71 B 0.008026f
C277 VTAIL.n72 B 0.014937f
C278 VTAIL.n73 B 0.014937f
C279 VTAIL.n74 B 0.008026f
C280 VTAIL.n75 B 0.008498f
C281 VTAIL.n76 B 0.018971f
C282 VTAIL.n77 B 0.018971f
C283 VTAIL.n78 B 0.008498f
C284 VTAIL.n79 B 0.008026f
C285 VTAIL.n80 B 0.014937f
C286 VTAIL.n81 B 0.014937f
C287 VTAIL.n82 B 0.008026f
C288 VTAIL.n83 B 0.008262f
C289 VTAIL.n84 B 0.008262f
C290 VTAIL.n85 B 0.018971f
C291 VTAIL.n86 B 0.041248f
C292 VTAIL.n87 B 0.008498f
C293 VTAIL.n88 B 0.008026f
C294 VTAIL.n89 B 0.03881f
C295 VTAIL.n90 B 0.023223f
C296 VTAIL.n91 B 0.925494f
C297 VTAIL.n92 B 0.021096f
C298 VTAIL.n93 B 0.014937f
C299 VTAIL.n94 B 0.008026f
C300 VTAIL.n95 B 0.018971f
C301 VTAIL.n96 B 0.008498f
C302 VTAIL.n97 B 0.014937f
C303 VTAIL.n98 B 0.008026f
C304 VTAIL.n99 B 0.018971f
C305 VTAIL.n100 B 0.018971f
C306 VTAIL.n101 B 0.008498f
C307 VTAIL.n102 B 0.014937f
C308 VTAIL.n103 B 0.008026f
C309 VTAIL.n104 B 0.018971f
C310 VTAIL.n105 B 0.008498f
C311 VTAIL.n106 B 0.088951f
C312 VTAIL.t0 B 0.031784f
C313 VTAIL.n107 B 0.014228f
C314 VTAIL.n108 B 0.013411f
C315 VTAIL.n109 B 0.008026f
C316 VTAIL.n110 B 0.536264f
C317 VTAIL.n111 B 0.014937f
C318 VTAIL.n112 B 0.008026f
C319 VTAIL.n113 B 0.008498f
C320 VTAIL.n114 B 0.018971f
C321 VTAIL.n115 B 0.018971f
C322 VTAIL.n116 B 0.008498f
C323 VTAIL.n117 B 0.008026f
C324 VTAIL.n118 B 0.014937f
C325 VTAIL.n119 B 0.014937f
C326 VTAIL.n120 B 0.008026f
C327 VTAIL.n121 B 0.008498f
C328 VTAIL.n122 B 0.018971f
C329 VTAIL.n123 B 0.018971f
C330 VTAIL.n124 B 0.008498f
C331 VTAIL.n125 B 0.008026f
C332 VTAIL.n126 B 0.014937f
C333 VTAIL.n127 B 0.014937f
C334 VTAIL.n128 B 0.008026f
C335 VTAIL.n129 B 0.008262f
C336 VTAIL.n130 B 0.008262f
C337 VTAIL.n131 B 0.018971f
C338 VTAIL.n132 B 0.041248f
C339 VTAIL.n133 B 0.008498f
C340 VTAIL.n134 B 0.008026f
C341 VTAIL.n135 B 0.03881f
C342 VTAIL.n136 B 0.023223f
C343 VTAIL.n137 B 0.796458f
C344 VTAIL.n138 B 0.021096f
C345 VTAIL.n139 B 0.014937f
C346 VTAIL.n140 B 0.008026f
C347 VTAIL.n141 B 0.018971f
C348 VTAIL.n142 B 0.008498f
C349 VTAIL.n143 B 0.014937f
C350 VTAIL.n144 B 0.008026f
C351 VTAIL.n145 B 0.018971f
C352 VTAIL.n146 B 0.008498f
C353 VTAIL.n147 B 0.014937f
C354 VTAIL.n148 B 0.008026f
C355 VTAIL.n149 B 0.018971f
C356 VTAIL.n150 B 0.008498f
C357 VTAIL.n151 B 0.088951f
C358 VTAIL.t2 B 0.031784f
C359 VTAIL.n152 B 0.014228f
C360 VTAIL.n153 B 0.013411f
C361 VTAIL.n154 B 0.008026f
C362 VTAIL.n155 B 0.536264f
C363 VTAIL.n156 B 0.014937f
C364 VTAIL.n157 B 0.008026f
C365 VTAIL.n158 B 0.008498f
C366 VTAIL.n159 B 0.018971f
C367 VTAIL.n160 B 0.018971f
C368 VTAIL.n161 B 0.008498f
C369 VTAIL.n162 B 0.008026f
C370 VTAIL.n163 B 0.014937f
C371 VTAIL.n164 B 0.014937f
C372 VTAIL.n165 B 0.008026f
C373 VTAIL.n166 B 0.008498f
C374 VTAIL.n167 B 0.018971f
C375 VTAIL.n168 B 0.018971f
C376 VTAIL.n169 B 0.018971f
C377 VTAIL.n170 B 0.008498f
C378 VTAIL.n171 B 0.008026f
C379 VTAIL.n172 B 0.014937f
C380 VTAIL.n173 B 0.014937f
C381 VTAIL.n174 B 0.008026f
C382 VTAIL.n175 B 0.008262f
C383 VTAIL.n176 B 0.008262f
C384 VTAIL.n177 B 0.018971f
C385 VTAIL.n178 B 0.041248f
C386 VTAIL.n179 B 0.008498f
C387 VTAIL.n180 B 0.008026f
C388 VTAIL.n181 B 0.03881f
C389 VTAIL.n182 B 0.023223f
C390 VTAIL.n183 B 0.738786f
C391 VN.t1 B 1.84354f
C392 VN.t0 B 2.27954f
.ends

