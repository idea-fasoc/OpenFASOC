* NGSPICE file created from diff_pair_sample_1232.ext - technology: sky130A

.subckt diff_pair_sample_1232 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 w_n1766_n2264# sky130_fd_pr__pfet_01v8 ad=2.5272 pd=13.74 as=2.5272 ps=13.74 w=6.48 l=1.66
X1 B.t11 B.t9 B.t10 w_n1766_n2264# sky130_fd_pr__pfet_01v8 ad=2.5272 pd=13.74 as=0 ps=0 w=6.48 l=1.66
X2 VDD2.t1 VN.t0 VTAIL.t0 w_n1766_n2264# sky130_fd_pr__pfet_01v8 ad=2.5272 pd=13.74 as=2.5272 ps=13.74 w=6.48 l=1.66
X3 VDD2.t0 VN.t1 VTAIL.t1 w_n1766_n2264# sky130_fd_pr__pfet_01v8 ad=2.5272 pd=13.74 as=2.5272 ps=13.74 w=6.48 l=1.66
X4 B.t8 B.t6 B.t7 w_n1766_n2264# sky130_fd_pr__pfet_01v8 ad=2.5272 pd=13.74 as=0 ps=0 w=6.48 l=1.66
X5 VDD1.t0 VP.t1 VTAIL.t3 w_n1766_n2264# sky130_fd_pr__pfet_01v8 ad=2.5272 pd=13.74 as=2.5272 ps=13.74 w=6.48 l=1.66
X6 B.t5 B.t3 B.t4 w_n1766_n2264# sky130_fd_pr__pfet_01v8 ad=2.5272 pd=13.74 as=0 ps=0 w=6.48 l=1.66
X7 B.t2 B.t0 B.t1 w_n1766_n2264# sky130_fd_pr__pfet_01v8 ad=2.5272 pd=13.74 as=0 ps=0 w=6.48 l=1.66
R0 VP.n0 VP.t0 190.946
R1 VP.n0 VP.t1 152.964
R2 VP VP.n0 0.241678
R3 VTAIL.n134 VTAIL.n133 756.745
R4 VTAIL.n32 VTAIL.n31 756.745
R5 VTAIL.n100 VTAIL.n99 756.745
R6 VTAIL.n66 VTAIL.n65 756.745
R7 VTAIL.n112 VTAIL.n111 585
R8 VTAIL.n117 VTAIL.n116 585
R9 VTAIL.n119 VTAIL.n118 585
R10 VTAIL.n108 VTAIL.n107 585
R11 VTAIL.n125 VTAIL.n124 585
R12 VTAIL.n127 VTAIL.n126 585
R13 VTAIL.n104 VTAIL.n103 585
R14 VTAIL.n133 VTAIL.n132 585
R15 VTAIL.n10 VTAIL.n9 585
R16 VTAIL.n15 VTAIL.n14 585
R17 VTAIL.n17 VTAIL.n16 585
R18 VTAIL.n6 VTAIL.n5 585
R19 VTAIL.n23 VTAIL.n22 585
R20 VTAIL.n25 VTAIL.n24 585
R21 VTAIL.n2 VTAIL.n1 585
R22 VTAIL.n31 VTAIL.n30 585
R23 VTAIL.n99 VTAIL.n98 585
R24 VTAIL.n70 VTAIL.n69 585
R25 VTAIL.n93 VTAIL.n92 585
R26 VTAIL.n91 VTAIL.n90 585
R27 VTAIL.n74 VTAIL.n73 585
R28 VTAIL.n85 VTAIL.n84 585
R29 VTAIL.n83 VTAIL.n82 585
R30 VTAIL.n78 VTAIL.n77 585
R31 VTAIL.n65 VTAIL.n64 585
R32 VTAIL.n36 VTAIL.n35 585
R33 VTAIL.n59 VTAIL.n58 585
R34 VTAIL.n57 VTAIL.n56 585
R35 VTAIL.n40 VTAIL.n39 585
R36 VTAIL.n51 VTAIL.n50 585
R37 VTAIL.n49 VTAIL.n48 585
R38 VTAIL.n44 VTAIL.n43 585
R39 VTAIL.n113 VTAIL.t0 329.084
R40 VTAIL.n11 VTAIL.t3 329.084
R41 VTAIL.n79 VTAIL.t2 329.084
R42 VTAIL.n45 VTAIL.t1 329.084
R43 VTAIL.n117 VTAIL.n111 171.744
R44 VTAIL.n118 VTAIL.n117 171.744
R45 VTAIL.n118 VTAIL.n107 171.744
R46 VTAIL.n125 VTAIL.n107 171.744
R47 VTAIL.n126 VTAIL.n125 171.744
R48 VTAIL.n126 VTAIL.n103 171.744
R49 VTAIL.n133 VTAIL.n103 171.744
R50 VTAIL.n15 VTAIL.n9 171.744
R51 VTAIL.n16 VTAIL.n15 171.744
R52 VTAIL.n16 VTAIL.n5 171.744
R53 VTAIL.n23 VTAIL.n5 171.744
R54 VTAIL.n24 VTAIL.n23 171.744
R55 VTAIL.n24 VTAIL.n1 171.744
R56 VTAIL.n31 VTAIL.n1 171.744
R57 VTAIL.n99 VTAIL.n69 171.744
R58 VTAIL.n92 VTAIL.n69 171.744
R59 VTAIL.n92 VTAIL.n91 171.744
R60 VTAIL.n91 VTAIL.n73 171.744
R61 VTAIL.n84 VTAIL.n73 171.744
R62 VTAIL.n84 VTAIL.n83 171.744
R63 VTAIL.n83 VTAIL.n77 171.744
R64 VTAIL.n65 VTAIL.n35 171.744
R65 VTAIL.n58 VTAIL.n35 171.744
R66 VTAIL.n58 VTAIL.n57 171.744
R67 VTAIL.n57 VTAIL.n39 171.744
R68 VTAIL.n50 VTAIL.n39 171.744
R69 VTAIL.n50 VTAIL.n49 171.744
R70 VTAIL.n49 VTAIL.n43 171.744
R71 VTAIL.t0 VTAIL.n111 85.8723
R72 VTAIL.t3 VTAIL.n9 85.8723
R73 VTAIL.t2 VTAIL.n77 85.8723
R74 VTAIL.t1 VTAIL.n43 85.8723
R75 VTAIL.n135 VTAIL.n134 34.1247
R76 VTAIL.n33 VTAIL.n32 34.1247
R77 VTAIL.n101 VTAIL.n100 34.1247
R78 VTAIL.n67 VTAIL.n66 34.1247
R79 VTAIL.n67 VTAIL.n33 21.3841
R80 VTAIL.n135 VTAIL.n101 19.6686
R81 VTAIL.n132 VTAIL.n102 12.8005
R82 VTAIL.n30 VTAIL.n0 12.8005
R83 VTAIL.n98 VTAIL.n68 12.8005
R84 VTAIL.n64 VTAIL.n34 12.8005
R85 VTAIL.n131 VTAIL.n104 12.0247
R86 VTAIL.n29 VTAIL.n2 12.0247
R87 VTAIL.n97 VTAIL.n70 12.0247
R88 VTAIL.n63 VTAIL.n36 12.0247
R89 VTAIL.n128 VTAIL.n127 11.249
R90 VTAIL.n26 VTAIL.n25 11.249
R91 VTAIL.n94 VTAIL.n93 11.249
R92 VTAIL.n60 VTAIL.n59 11.249
R93 VTAIL.n113 VTAIL.n112 10.7233
R94 VTAIL.n11 VTAIL.n10 10.7233
R95 VTAIL.n79 VTAIL.n78 10.7233
R96 VTAIL.n45 VTAIL.n44 10.7233
R97 VTAIL.n124 VTAIL.n106 10.4732
R98 VTAIL.n22 VTAIL.n4 10.4732
R99 VTAIL.n90 VTAIL.n72 10.4732
R100 VTAIL.n56 VTAIL.n38 10.4732
R101 VTAIL.n123 VTAIL.n108 9.69747
R102 VTAIL.n21 VTAIL.n6 9.69747
R103 VTAIL.n89 VTAIL.n74 9.69747
R104 VTAIL.n55 VTAIL.n40 9.69747
R105 VTAIL.n130 VTAIL.n102 9.45567
R106 VTAIL.n28 VTAIL.n0 9.45567
R107 VTAIL.n96 VTAIL.n68 9.45567
R108 VTAIL.n62 VTAIL.n34 9.45567
R109 VTAIL.n115 VTAIL.n114 9.3005
R110 VTAIL.n110 VTAIL.n109 9.3005
R111 VTAIL.n121 VTAIL.n120 9.3005
R112 VTAIL.n123 VTAIL.n122 9.3005
R113 VTAIL.n106 VTAIL.n105 9.3005
R114 VTAIL.n129 VTAIL.n128 9.3005
R115 VTAIL.n131 VTAIL.n130 9.3005
R116 VTAIL.n13 VTAIL.n12 9.3005
R117 VTAIL.n8 VTAIL.n7 9.3005
R118 VTAIL.n19 VTAIL.n18 9.3005
R119 VTAIL.n21 VTAIL.n20 9.3005
R120 VTAIL.n4 VTAIL.n3 9.3005
R121 VTAIL.n27 VTAIL.n26 9.3005
R122 VTAIL.n29 VTAIL.n28 9.3005
R123 VTAIL.n97 VTAIL.n96 9.3005
R124 VTAIL.n95 VTAIL.n94 9.3005
R125 VTAIL.n72 VTAIL.n71 9.3005
R126 VTAIL.n89 VTAIL.n88 9.3005
R127 VTAIL.n87 VTAIL.n86 9.3005
R128 VTAIL.n76 VTAIL.n75 9.3005
R129 VTAIL.n81 VTAIL.n80 9.3005
R130 VTAIL.n42 VTAIL.n41 9.3005
R131 VTAIL.n53 VTAIL.n52 9.3005
R132 VTAIL.n55 VTAIL.n54 9.3005
R133 VTAIL.n38 VTAIL.n37 9.3005
R134 VTAIL.n61 VTAIL.n60 9.3005
R135 VTAIL.n63 VTAIL.n62 9.3005
R136 VTAIL.n47 VTAIL.n46 9.3005
R137 VTAIL.n120 VTAIL.n119 8.92171
R138 VTAIL.n18 VTAIL.n17 8.92171
R139 VTAIL.n86 VTAIL.n85 8.92171
R140 VTAIL.n52 VTAIL.n51 8.92171
R141 VTAIL.n116 VTAIL.n110 8.14595
R142 VTAIL.n14 VTAIL.n8 8.14595
R143 VTAIL.n82 VTAIL.n76 8.14595
R144 VTAIL.n48 VTAIL.n42 8.14595
R145 VTAIL.n115 VTAIL.n112 7.3702
R146 VTAIL.n13 VTAIL.n10 7.3702
R147 VTAIL.n81 VTAIL.n78 7.3702
R148 VTAIL.n47 VTAIL.n44 7.3702
R149 VTAIL.n116 VTAIL.n115 5.81868
R150 VTAIL.n14 VTAIL.n13 5.81868
R151 VTAIL.n82 VTAIL.n81 5.81868
R152 VTAIL.n48 VTAIL.n47 5.81868
R153 VTAIL.n119 VTAIL.n110 5.04292
R154 VTAIL.n17 VTAIL.n8 5.04292
R155 VTAIL.n85 VTAIL.n76 5.04292
R156 VTAIL.n51 VTAIL.n42 5.04292
R157 VTAIL.n120 VTAIL.n108 4.26717
R158 VTAIL.n18 VTAIL.n6 4.26717
R159 VTAIL.n86 VTAIL.n74 4.26717
R160 VTAIL.n52 VTAIL.n40 4.26717
R161 VTAIL.n124 VTAIL.n123 3.49141
R162 VTAIL.n22 VTAIL.n21 3.49141
R163 VTAIL.n90 VTAIL.n89 3.49141
R164 VTAIL.n56 VTAIL.n55 3.49141
R165 VTAIL.n127 VTAIL.n106 2.71565
R166 VTAIL.n25 VTAIL.n4 2.71565
R167 VTAIL.n93 VTAIL.n72 2.71565
R168 VTAIL.n59 VTAIL.n38 2.71565
R169 VTAIL.n46 VTAIL.n45 2.41347
R170 VTAIL.n114 VTAIL.n113 2.41347
R171 VTAIL.n12 VTAIL.n11 2.41347
R172 VTAIL.n80 VTAIL.n79 2.41347
R173 VTAIL.n128 VTAIL.n104 1.93989
R174 VTAIL.n26 VTAIL.n2 1.93989
R175 VTAIL.n94 VTAIL.n70 1.93989
R176 VTAIL.n60 VTAIL.n36 1.93989
R177 VTAIL.n101 VTAIL.n67 1.32809
R178 VTAIL.n132 VTAIL.n131 1.16414
R179 VTAIL.n30 VTAIL.n29 1.16414
R180 VTAIL.n98 VTAIL.n97 1.16414
R181 VTAIL.n64 VTAIL.n63 1.16414
R182 VTAIL VTAIL.n33 0.957397
R183 VTAIL.n134 VTAIL.n102 0.388379
R184 VTAIL.n32 VTAIL.n0 0.388379
R185 VTAIL.n100 VTAIL.n68 0.388379
R186 VTAIL.n66 VTAIL.n34 0.388379
R187 VTAIL VTAIL.n135 0.37119
R188 VTAIL.n114 VTAIL.n109 0.155672
R189 VTAIL.n121 VTAIL.n109 0.155672
R190 VTAIL.n122 VTAIL.n121 0.155672
R191 VTAIL.n122 VTAIL.n105 0.155672
R192 VTAIL.n129 VTAIL.n105 0.155672
R193 VTAIL.n130 VTAIL.n129 0.155672
R194 VTAIL.n12 VTAIL.n7 0.155672
R195 VTAIL.n19 VTAIL.n7 0.155672
R196 VTAIL.n20 VTAIL.n19 0.155672
R197 VTAIL.n20 VTAIL.n3 0.155672
R198 VTAIL.n27 VTAIL.n3 0.155672
R199 VTAIL.n28 VTAIL.n27 0.155672
R200 VTAIL.n96 VTAIL.n95 0.155672
R201 VTAIL.n95 VTAIL.n71 0.155672
R202 VTAIL.n88 VTAIL.n71 0.155672
R203 VTAIL.n88 VTAIL.n87 0.155672
R204 VTAIL.n87 VTAIL.n75 0.155672
R205 VTAIL.n80 VTAIL.n75 0.155672
R206 VTAIL.n62 VTAIL.n61 0.155672
R207 VTAIL.n61 VTAIL.n37 0.155672
R208 VTAIL.n54 VTAIL.n37 0.155672
R209 VTAIL.n54 VTAIL.n53 0.155672
R210 VTAIL.n53 VTAIL.n41 0.155672
R211 VTAIL.n46 VTAIL.n41 0.155672
R212 VDD1.n32 VDD1.n31 756.745
R213 VDD1.n65 VDD1.n64 756.745
R214 VDD1.n31 VDD1.n30 585
R215 VDD1.n2 VDD1.n1 585
R216 VDD1.n25 VDD1.n24 585
R217 VDD1.n23 VDD1.n22 585
R218 VDD1.n6 VDD1.n5 585
R219 VDD1.n17 VDD1.n16 585
R220 VDD1.n15 VDD1.n14 585
R221 VDD1.n10 VDD1.n9 585
R222 VDD1.n43 VDD1.n42 585
R223 VDD1.n48 VDD1.n47 585
R224 VDD1.n50 VDD1.n49 585
R225 VDD1.n39 VDD1.n38 585
R226 VDD1.n56 VDD1.n55 585
R227 VDD1.n58 VDD1.n57 585
R228 VDD1.n35 VDD1.n34 585
R229 VDD1.n64 VDD1.n63 585
R230 VDD1.n11 VDD1.t1 329.084
R231 VDD1.n44 VDD1.t0 329.084
R232 VDD1.n31 VDD1.n1 171.744
R233 VDD1.n24 VDD1.n1 171.744
R234 VDD1.n24 VDD1.n23 171.744
R235 VDD1.n23 VDD1.n5 171.744
R236 VDD1.n16 VDD1.n5 171.744
R237 VDD1.n16 VDD1.n15 171.744
R238 VDD1.n15 VDD1.n9 171.744
R239 VDD1.n48 VDD1.n42 171.744
R240 VDD1.n49 VDD1.n48 171.744
R241 VDD1.n49 VDD1.n38 171.744
R242 VDD1.n56 VDD1.n38 171.744
R243 VDD1.n57 VDD1.n56 171.744
R244 VDD1.n57 VDD1.n34 171.744
R245 VDD1.n64 VDD1.n34 171.744
R246 VDD1.t1 VDD1.n9 85.8723
R247 VDD1.t0 VDD1.n42 85.8723
R248 VDD1 VDD1.n65 84.4339
R249 VDD1 VDD1.n32 51.2906
R250 VDD1.n30 VDD1.n0 12.8005
R251 VDD1.n63 VDD1.n33 12.8005
R252 VDD1.n29 VDD1.n2 12.0247
R253 VDD1.n62 VDD1.n35 12.0247
R254 VDD1.n26 VDD1.n25 11.249
R255 VDD1.n59 VDD1.n58 11.249
R256 VDD1.n11 VDD1.n10 10.7233
R257 VDD1.n44 VDD1.n43 10.7233
R258 VDD1.n22 VDD1.n4 10.4732
R259 VDD1.n55 VDD1.n37 10.4732
R260 VDD1.n21 VDD1.n6 9.69747
R261 VDD1.n54 VDD1.n39 9.69747
R262 VDD1.n28 VDD1.n0 9.45567
R263 VDD1.n61 VDD1.n33 9.45567
R264 VDD1.n29 VDD1.n28 9.3005
R265 VDD1.n27 VDD1.n26 9.3005
R266 VDD1.n4 VDD1.n3 9.3005
R267 VDD1.n21 VDD1.n20 9.3005
R268 VDD1.n19 VDD1.n18 9.3005
R269 VDD1.n8 VDD1.n7 9.3005
R270 VDD1.n13 VDD1.n12 9.3005
R271 VDD1.n46 VDD1.n45 9.3005
R272 VDD1.n41 VDD1.n40 9.3005
R273 VDD1.n52 VDD1.n51 9.3005
R274 VDD1.n54 VDD1.n53 9.3005
R275 VDD1.n37 VDD1.n36 9.3005
R276 VDD1.n60 VDD1.n59 9.3005
R277 VDD1.n62 VDD1.n61 9.3005
R278 VDD1.n18 VDD1.n17 8.92171
R279 VDD1.n51 VDD1.n50 8.92171
R280 VDD1.n14 VDD1.n8 8.14595
R281 VDD1.n47 VDD1.n41 8.14595
R282 VDD1.n13 VDD1.n10 7.3702
R283 VDD1.n46 VDD1.n43 7.3702
R284 VDD1.n14 VDD1.n13 5.81868
R285 VDD1.n47 VDD1.n46 5.81868
R286 VDD1.n17 VDD1.n8 5.04292
R287 VDD1.n50 VDD1.n41 5.04292
R288 VDD1.n18 VDD1.n6 4.26717
R289 VDD1.n51 VDD1.n39 4.26717
R290 VDD1.n22 VDD1.n21 3.49141
R291 VDD1.n55 VDD1.n54 3.49141
R292 VDD1.n25 VDD1.n4 2.71565
R293 VDD1.n58 VDD1.n37 2.71565
R294 VDD1.n12 VDD1.n11 2.41347
R295 VDD1.n45 VDD1.n44 2.41347
R296 VDD1.n26 VDD1.n2 1.93989
R297 VDD1.n59 VDD1.n35 1.93989
R298 VDD1.n30 VDD1.n29 1.16414
R299 VDD1.n63 VDD1.n62 1.16414
R300 VDD1.n32 VDD1.n0 0.388379
R301 VDD1.n65 VDD1.n33 0.388379
R302 VDD1.n28 VDD1.n27 0.155672
R303 VDD1.n27 VDD1.n3 0.155672
R304 VDD1.n20 VDD1.n3 0.155672
R305 VDD1.n20 VDD1.n19 0.155672
R306 VDD1.n19 VDD1.n7 0.155672
R307 VDD1.n12 VDD1.n7 0.155672
R308 VDD1.n45 VDD1.n40 0.155672
R309 VDD1.n52 VDD1.n40 0.155672
R310 VDD1.n53 VDD1.n52 0.155672
R311 VDD1.n53 VDD1.n36 0.155672
R312 VDD1.n60 VDD1.n36 0.155672
R313 VDD1.n61 VDD1.n60 0.155672
R314 B.n294 B.n293 585
R315 B.n295 B.n46 585
R316 B.n297 B.n296 585
R317 B.n298 B.n45 585
R318 B.n300 B.n299 585
R319 B.n301 B.n44 585
R320 B.n303 B.n302 585
R321 B.n304 B.n43 585
R322 B.n306 B.n305 585
R323 B.n307 B.n42 585
R324 B.n309 B.n308 585
R325 B.n310 B.n41 585
R326 B.n312 B.n311 585
R327 B.n313 B.n40 585
R328 B.n315 B.n314 585
R329 B.n316 B.n39 585
R330 B.n318 B.n317 585
R331 B.n319 B.n38 585
R332 B.n321 B.n320 585
R333 B.n322 B.n37 585
R334 B.n324 B.n323 585
R335 B.n325 B.n36 585
R336 B.n327 B.n326 585
R337 B.n328 B.n35 585
R338 B.n330 B.n329 585
R339 B.n332 B.n32 585
R340 B.n334 B.n333 585
R341 B.n335 B.n31 585
R342 B.n337 B.n336 585
R343 B.n338 B.n30 585
R344 B.n340 B.n339 585
R345 B.n341 B.n29 585
R346 B.n343 B.n342 585
R347 B.n344 B.n25 585
R348 B.n346 B.n345 585
R349 B.n347 B.n24 585
R350 B.n349 B.n348 585
R351 B.n350 B.n23 585
R352 B.n352 B.n351 585
R353 B.n353 B.n22 585
R354 B.n355 B.n354 585
R355 B.n356 B.n21 585
R356 B.n358 B.n357 585
R357 B.n359 B.n20 585
R358 B.n361 B.n360 585
R359 B.n362 B.n19 585
R360 B.n364 B.n363 585
R361 B.n365 B.n18 585
R362 B.n367 B.n366 585
R363 B.n368 B.n17 585
R364 B.n370 B.n369 585
R365 B.n371 B.n16 585
R366 B.n373 B.n372 585
R367 B.n374 B.n15 585
R368 B.n376 B.n375 585
R369 B.n377 B.n14 585
R370 B.n379 B.n378 585
R371 B.n380 B.n13 585
R372 B.n382 B.n381 585
R373 B.n383 B.n12 585
R374 B.n292 B.n47 585
R375 B.n291 B.n290 585
R376 B.n289 B.n48 585
R377 B.n288 B.n287 585
R378 B.n286 B.n49 585
R379 B.n285 B.n284 585
R380 B.n283 B.n50 585
R381 B.n282 B.n281 585
R382 B.n280 B.n51 585
R383 B.n279 B.n278 585
R384 B.n277 B.n52 585
R385 B.n276 B.n275 585
R386 B.n274 B.n53 585
R387 B.n273 B.n272 585
R388 B.n271 B.n54 585
R389 B.n270 B.n269 585
R390 B.n268 B.n55 585
R391 B.n267 B.n266 585
R392 B.n265 B.n56 585
R393 B.n264 B.n263 585
R394 B.n262 B.n57 585
R395 B.n261 B.n260 585
R396 B.n259 B.n58 585
R397 B.n258 B.n257 585
R398 B.n256 B.n59 585
R399 B.n255 B.n254 585
R400 B.n253 B.n60 585
R401 B.n252 B.n251 585
R402 B.n250 B.n61 585
R403 B.n249 B.n248 585
R404 B.n247 B.n62 585
R405 B.n246 B.n245 585
R406 B.n244 B.n63 585
R407 B.n243 B.n242 585
R408 B.n241 B.n64 585
R409 B.n240 B.n239 585
R410 B.n238 B.n65 585
R411 B.n237 B.n236 585
R412 B.n235 B.n66 585
R413 B.n234 B.n233 585
R414 B.n232 B.n67 585
R415 B.n141 B.n140 585
R416 B.n142 B.n101 585
R417 B.n144 B.n143 585
R418 B.n145 B.n100 585
R419 B.n147 B.n146 585
R420 B.n148 B.n99 585
R421 B.n150 B.n149 585
R422 B.n151 B.n98 585
R423 B.n153 B.n152 585
R424 B.n154 B.n97 585
R425 B.n156 B.n155 585
R426 B.n157 B.n96 585
R427 B.n159 B.n158 585
R428 B.n160 B.n95 585
R429 B.n162 B.n161 585
R430 B.n163 B.n94 585
R431 B.n165 B.n164 585
R432 B.n166 B.n93 585
R433 B.n168 B.n167 585
R434 B.n169 B.n92 585
R435 B.n171 B.n170 585
R436 B.n172 B.n91 585
R437 B.n174 B.n173 585
R438 B.n175 B.n90 585
R439 B.n177 B.n176 585
R440 B.n179 B.n178 585
R441 B.n180 B.n86 585
R442 B.n182 B.n181 585
R443 B.n183 B.n85 585
R444 B.n185 B.n184 585
R445 B.n186 B.n84 585
R446 B.n188 B.n187 585
R447 B.n189 B.n83 585
R448 B.n191 B.n190 585
R449 B.n192 B.n80 585
R450 B.n195 B.n194 585
R451 B.n196 B.n79 585
R452 B.n198 B.n197 585
R453 B.n199 B.n78 585
R454 B.n201 B.n200 585
R455 B.n202 B.n77 585
R456 B.n204 B.n203 585
R457 B.n205 B.n76 585
R458 B.n207 B.n206 585
R459 B.n208 B.n75 585
R460 B.n210 B.n209 585
R461 B.n211 B.n74 585
R462 B.n213 B.n212 585
R463 B.n214 B.n73 585
R464 B.n216 B.n215 585
R465 B.n217 B.n72 585
R466 B.n219 B.n218 585
R467 B.n220 B.n71 585
R468 B.n222 B.n221 585
R469 B.n223 B.n70 585
R470 B.n225 B.n224 585
R471 B.n226 B.n69 585
R472 B.n228 B.n227 585
R473 B.n229 B.n68 585
R474 B.n231 B.n230 585
R475 B.n139 B.n102 585
R476 B.n138 B.n137 585
R477 B.n136 B.n103 585
R478 B.n135 B.n134 585
R479 B.n133 B.n104 585
R480 B.n132 B.n131 585
R481 B.n130 B.n105 585
R482 B.n129 B.n128 585
R483 B.n127 B.n106 585
R484 B.n126 B.n125 585
R485 B.n124 B.n107 585
R486 B.n123 B.n122 585
R487 B.n121 B.n108 585
R488 B.n120 B.n119 585
R489 B.n118 B.n109 585
R490 B.n117 B.n116 585
R491 B.n115 B.n110 585
R492 B.n114 B.n113 585
R493 B.n112 B.n111 585
R494 B.n2 B.n0 585
R495 B.n413 B.n1 585
R496 B.n412 B.n411 585
R497 B.n410 B.n3 585
R498 B.n409 B.n408 585
R499 B.n407 B.n4 585
R500 B.n406 B.n405 585
R501 B.n404 B.n5 585
R502 B.n403 B.n402 585
R503 B.n401 B.n6 585
R504 B.n400 B.n399 585
R505 B.n398 B.n7 585
R506 B.n397 B.n396 585
R507 B.n395 B.n8 585
R508 B.n394 B.n393 585
R509 B.n392 B.n9 585
R510 B.n391 B.n390 585
R511 B.n389 B.n10 585
R512 B.n388 B.n387 585
R513 B.n386 B.n11 585
R514 B.n385 B.n384 585
R515 B.n415 B.n414 585
R516 B.n141 B.n102 497.305
R517 B.n384 B.n383 497.305
R518 B.n232 B.n231 497.305
R519 B.n293 B.n292 497.305
R520 B.n81 B.t11 314.901
R521 B.n33 B.t4 314.901
R522 B.n87 B.t8 314.901
R523 B.n26 B.t1 314.901
R524 B.n81 B.t9 300.067
R525 B.n87 B.t6 300.067
R526 B.n26 B.t0 300.067
R527 B.n33 B.t3 300.067
R528 B.n82 B.t10 276.308
R529 B.n34 B.t5 276.308
R530 B.n88 B.t7 276.308
R531 B.n27 B.t2 276.308
R532 B.n137 B.n102 163.367
R533 B.n137 B.n136 163.367
R534 B.n136 B.n135 163.367
R535 B.n135 B.n104 163.367
R536 B.n131 B.n104 163.367
R537 B.n131 B.n130 163.367
R538 B.n130 B.n129 163.367
R539 B.n129 B.n106 163.367
R540 B.n125 B.n106 163.367
R541 B.n125 B.n124 163.367
R542 B.n124 B.n123 163.367
R543 B.n123 B.n108 163.367
R544 B.n119 B.n108 163.367
R545 B.n119 B.n118 163.367
R546 B.n118 B.n117 163.367
R547 B.n117 B.n110 163.367
R548 B.n113 B.n110 163.367
R549 B.n113 B.n112 163.367
R550 B.n112 B.n2 163.367
R551 B.n414 B.n2 163.367
R552 B.n414 B.n413 163.367
R553 B.n413 B.n412 163.367
R554 B.n412 B.n3 163.367
R555 B.n408 B.n3 163.367
R556 B.n408 B.n407 163.367
R557 B.n407 B.n406 163.367
R558 B.n406 B.n5 163.367
R559 B.n402 B.n5 163.367
R560 B.n402 B.n401 163.367
R561 B.n401 B.n400 163.367
R562 B.n400 B.n7 163.367
R563 B.n396 B.n7 163.367
R564 B.n396 B.n395 163.367
R565 B.n395 B.n394 163.367
R566 B.n394 B.n9 163.367
R567 B.n390 B.n9 163.367
R568 B.n390 B.n389 163.367
R569 B.n389 B.n388 163.367
R570 B.n388 B.n11 163.367
R571 B.n384 B.n11 163.367
R572 B.n142 B.n141 163.367
R573 B.n143 B.n142 163.367
R574 B.n143 B.n100 163.367
R575 B.n147 B.n100 163.367
R576 B.n148 B.n147 163.367
R577 B.n149 B.n148 163.367
R578 B.n149 B.n98 163.367
R579 B.n153 B.n98 163.367
R580 B.n154 B.n153 163.367
R581 B.n155 B.n154 163.367
R582 B.n155 B.n96 163.367
R583 B.n159 B.n96 163.367
R584 B.n160 B.n159 163.367
R585 B.n161 B.n160 163.367
R586 B.n161 B.n94 163.367
R587 B.n165 B.n94 163.367
R588 B.n166 B.n165 163.367
R589 B.n167 B.n166 163.367
R590 B.n167 B.n92 163.367
R591 B.n171 B.n92 163.367
R592 B.n172 B.n171 163.367
R593 B.n173 B.n172 163.367
R594 B.n173 B.n90 163.367
R595 B.n177 B.n90 163.367
R596 B.n178 B.n177 163.367
R597 B.n178 B.n86 163.367
R598 B.n182 B.n86 163.367
R599 B.n183 B.n182 163.367
R600 B.n184 B.n183 163.367
R601 B.n184 B.n84 163.367
R602 B.n188 B.n84 163.367
R603 B.n189 B.n188 163.367
R604 B.n190 B.n189 163.367
R605 B.n190 B.n80 163.367
R606 B.n195 B.n80 163.367
R607 B.n196 B.n195 163.367
R608 B.n197 B.n196 163.367
R609 B.n197 B.n78 163.367
R610 B.n201 B.n78 163.367
R611 B.n202 B.n201 163.367
R612 B.n203 B.n202 163.367
R613 B.n203 B.n76 163.367
R614 B.n207 B.n76 163.367
R615 B.n208 B.n207 163.367
R616 B.n209 B.n208 163.367
R617 B.n209 B.n74 163.367
R618 B.n213 B.n74 163.367
R619 B.n214 B.n213 163.367
R620 B.n215 B.n214 163.367
R621 B.n215 B.n72 163.367
R622 B.n219 B.n72 163.367
R623 B.n220 B.n219 163.367
R624 B.n221 B.n220 163.367
R625 B.n221 B.n70 163.367
R626 B.n225 B.n70 163.367
R627 B.n226 B.n225 163.367
R628 B.n227 B.n226 163.367
R629 B.n227 B.n68 163.367
R630 B.n231 B.n68 163.367
R631 B.n233 B.n232 163.367
R632 B.n233 B.n66 163.367
R633 B.n237 B.n66 163.367
R634 B.n238 B.n237 163.367
R635 B.n239 B.n238 163.367
R636 B.n239 B.n64 163.367
R637 B.n243 B.n64 163.367
R638 B.n244 B.n243 163.367
R639 B.n245 B.n244 163.367
R640 B.n245 B.n62 163.367
R641 B.n249 B.n62 163.367
R642 B.n250 B.n249 163.367
R643 B.n251 B.n250 163.367
R644 B.n251 B.n60 163.367
R645 B.n255 B.n60 163.367
R646 B.n256 B.n255 163.367
R647 B.n257 B.n256 163.367
R648 B.n257 B.n58 163.367
R649 B.n261 B.n58 163.367
R650 B.n262 B.n261 163.367
R651 B.n263 B.n262 163.367
R652 B.n263 B.n56 163.367
R653 B.n267 B.n56 163.367
R654 B.n268 B.n267 163.367
R655 B.n269 B.n268 163.367
R656 B.n269 B.n54 163.367
R657 B.n273 B.n54 163.367
R658 B.n274 B.n273 163.367
R659 B.n275 B.n274 163.367
R660 B.n275 B.n52 163.367
R661 B.n279 B.n52 163.367
R662 B.n280 B.n279 163.367
R663 B.n281 B.n280 163.367
R664 B.n281 B.n50 163.367
R665 B.n285 B.n50 163.367
R666 B.n286 B.n285 163.367
R667 B.n287 B.n286 163.367
R668 B.n287 B.n48 163.367
R669 B.n291 B.n48 163.367
R670 B.n292 B.n291 163.367
R671 B.n383 B.n382 163.367
R672 B.n382 B.n13 163.367
R673 B.n378 B.n13 163.367
R674 B.n378 B.n377 163.367
R675 B.n377 B.n376 163.367
R676 B.n376 B.n15 163.367
R677 B.n372 B.n15 163.367
R678 B.n372 B.n371 163.367
R679 B.n371 B.n370 163.367
R680 B.n370 B.n17 163.367
R681 B.n366 B.n17 163.367
R682 B.n366 B.n365 163.367
R683 B.n365 B.n364 163.367
R684 B.n364 B.n19 163.367
R685 B.n360 B.n19 163.367
R686 B.n360 B.n359 163.367
R687 B.n359 B.n358 163.367
R688 B.n358 B.n21 163.367
R689 B.n354 B.n21 163.367
R690 B.n354 B.n353 163.367
R691 B.n353 B.n352 163.367
R692 B.n352 B.n23 163.367
R693 B.n348 B.n23 163.367
R694 B.n348 B.n347 163.367
R695 B.n347 B.n346 163.367
R696 B.n346 B.n25 163.367
R697 B.n342 B.n25 163.367
R698 B.n342 B.n341 163.367
R699 B.n341 B.n340 163.367
R700 B.n340 B.n30 163.367
R701 B.n336 B.n30 163.367
R702 B.n336 B.n335 163.367
R703 B.n335 B.n334 163.367
R704 B.n334 B.n32 163.367
R705 B.n329 B.n32 163.367
R706 B.n329 B.n328 163.367
R707 B.n328 B.n327 163.367
R708 B.n327 B.n36 163.367
R709 B.n323 B.n36 163.367
R710 B.n323 B.n322 163.367
R711 B.n322 B.n321 163.367
R712 B.n321 B.n38 163.367
R713 B.n317 B.n38 163.367
R714 B.n317 B.n316 163.367
R715 B.n316 B.n315 163.367
R716 B.n315 B.n40 163.367
R717 B.n311 B.n40 163.367
R718 B.n311 B.n310 163.367
R719 B.n310 B.n309 163.367
R720 B.n309 B.n42 163.367
R721 B.n305 B.n42 163.367
R722 B.n305 B.n304 163.367
R723 B.n304 B.n303 163.367
R724 B.n303 B.n44 163.367
R725 B.n299 B.n44 163.367
R726 B.n299 B.n298 163.367
R727 B.n298 B.n297 163.367
R728 B.n297 B.n46 163.367
R729 B.n293 B.n46 163.367
R730 B.n193 B.n82 59.5399
R731 B.n89 B.n88 59.5399
R732 B.n28 B.n27 59.5399
R733 B.n331 B.n34 59.5399
R734 B.n82 B.n81 38.5944
R735 B.n88 B.n87 38.5944
R736 B.n27 B.n26 38.5944
R737 B.n34 B.n33 38.5944
R738 B.n385 B.n12 32.3127
R739 B.n294 B.n47 32.3127
R740 B.n230 B.n67 32.3127
R741 B.n140 B.n139 32.3127
R742 B B.n415 18.0485
R743 B.n381 B.n12 10.6151
R744 B.n381 B.n380 10.6151
R745 B.n380 B.n379 10.6151
R746 B.n379 B.n14 10.6151
R747 B.n375 B.n14 10.6151
R748 B.n375 B.n374 10.6151
R749 B.n374 B.n373 10.6151
R750 B.n373 B.n16 10.6151
R751 B.n369 B.n16 10.6151
R752 B.n369 B.n368 10.6151
R753 B.n368 B.n367 10.6151
R754 B.n367 B.n18 10.6151
R755 B.n363 B.n18 10.6151
R756 B.n363 B.n362 10.6151
R757 B.n362 B.n361 10.6151
R758 B.n361 B.n20 10.6151
R759 B.n357 B.n20 10.6151
R760 B.n357 B.n356 10.6151
R761 B.n356 B.n355 10.6151
R762 B.n355 B.n22 10.6151
R763 B.n351 B.n22 10.6151
R764 B.n351 B.n350 10.6151
R765 B.n350 B.n349 10.6151
R766 B.n349 B.n24 10.6151
R767 B.n345 B.n344 10.6151
R768 B.n344 B.n343 10.6151
R769 B.n343 B.n29 10.6151
R770 B.n339 B.n29 10.6151
R771 B.n339 B.n338 10.6151
R772 B.n338 B.n337 10.6151
R773 B.n337 B.n31 10.6151
R774 B.n333 B.n31 10.6151
R775 B.n333 B.n332 10.6151
R776 B.n330 B.n35 10.6151
R777 B.n326 B.n35 10.6151
R778 B.n326 B.n325 10.6151
R779 B.n325 B.n324 10.6151
R780 B.n324 B.n37 10.6151
R781 B.n320 B.n37 10.6151
R782 B.n320 B.n319 10.6151
R783 B.n319 B.n318 10.6151
R784 B.n318 B.n39 10.6151
R785 B.n314 B.n39 10.6151
R786 B.n314 B.n313 10.6151
R787 B.n313 B.n312 10.6151
R788 B.n312 B.n41 10.6151
R789 B.n308 B.n41 10.6151
R790 B.n308 B.n307 10.6151
R791 B.n307 B.n306 10.6151
R792 B.n306 B.n43 10.6151
R793 B.n302 B.n43 10.6151
R794 B.n302 B.n301 10.6151
R795 B.n301 B.n300 10.6151
R796 B.n300 B.n45 10.6151
R797 B.n296 B.n45 10.6151
R798 B.n296 B.n295 10.6151
R799 B.n295 B.n294 10.6151
R800 B.n234 B.n67 10.6151
R801 B.n235 B.n234 10.6151
R802 B.n236 B.n235 10.6151
R803 B.n236 B.n65 10.6151
R804 B.n240 B.n65 10.6151
R805 B.n241 B.n240 10.6151
R806 B.n242 B.n241 10.6151
R807 B.n242 B.n63 10.6151
R808 B.n246 B.n63 10.6151
R809 B.n247 B.n246 10.6151
R810 B.n248 B.n247 10.6151
R811 B.n248 B.n61 10.6151
R812 B.n252 B.n61 10.6151
R813 B.n253 B.n252 10.6151
R814 B.n254 B.n253 10.6151
R815 B.n254 B.n59 10.6151
R816 B.n258 B.n59 10.6151
R817 B.n259 B.n258 10.6151
R818 B.n260 B.n259 10.6151
R819 B.n260 B.n57 10.6151
R820 B.n264 B.n57 10.6151
R821 B.n265 B.n264 10.6151
R822 B.n266 B.n265 10.6151
R823 B.n266 B.n55 10.6151
R824 B.n270 B.n55 10.6151
R825 B.n271 B.n270 10.6151
R826 B.n272 B.n271 10.6151
R827 B.n272 B.n53 10.6151
R828 B.n276 B.n53 10.6151
R829 B.n277 B.n276 10.6151
R830 B.n278 B.n277 10.6151
R831 B.n278 B.n51 10.6151
R832 B.n282 B.n51 10.6151
R833 B.n283 B.n282 10.6151
R834 B.n284 B.n283 10.6151
R835 B.n284 B.n49 10.6151
R836 B.n288 B.n49 10.6151
R837 B.n289 B.n288 10.6151
R838 B.n290 B.n289 10.6151
R839 B.n290 B.n47 10.6151
R840 B.n140 B.n101 10.6151
R841 B.n144 B.n101 10.6151
R842 B.n145 B.n144 10.6151
R843 B.n146 B.n145 10.6151
R844 B.n146 B.n99 10.6151
R845 B.n150 B.n99 10.6151
R846 B.n151 B.n150 10.6151
R847 B.n152 B.n151 10.6151
R848 B.n152 B.n97 10.6151
R849 B.n156 B.n97 10.6151
R850 B.n157 B.n156 10.6151
R851 B.n158 B.n157 10.6151
R852 B.n158 B.n95 10.6151
R853 B.n162 B.n95 10.6151
R854 B.n163 B.n162 10.6151
R855 B.n164 B.n163 10.6151
R856 B.n164 B.n93 10.6151
R857 B.n168 B.n93 10.6151
R858 B.n169 B.n168 10.6151
R859 B.n170 B.n169 10.6151
R860 B.n170 B.n91 10.6151
R861 B.n174 B.n91 10.6151
R862 B.n175 B.n174 10.6151
R863 B.n176 B.n175 10.6151
R864 B.n180 B.n179 10.6151
R865 B.n181 B.n180 10.6151
R866 B.n181 B.n85 10.6151
R867 B.n185 B.n85 10.6151
R868 B.n186 B.n185 10.6151
R869 B.n187 B.n186 10.6151
R870 B.n187 B.n83 10.6151
R871 B.n191 B.n83 10.6151
R872 B.n192 B.n191 10.6151
R873 B.n194 B.n79 10.6151
R874 B.n198 B.n79 10.6151
R875 B.n199 B.n198 10.6151
R876 B.n200 B.n199 10.6151
R877 B.n200 B.n77 10.6151
R878 B.n204 B.n77 10.6151
R879 B.n205 B.n204 10.6151
R880 B.n206 B.n205 10.6151
R881 B.n206 B.n75 10.6151
R882 B.n210 B.n75 10.6151
R883 B.n211 B.n210 10.6151
R884 B.n212 B.n211 10.6151
R885 B.n212 B.n73 10.6151
R886 B.n216 B.n73 10.6151
R887 B.n217 B.n216 10.6151
R888 B.n218 B.n217 10.6151
R889 B.n218 B.n71 10.6151
R890 B.n222 B.n71 10.6151
R891 B.n223 B.n222 10.6151
R892 B.n224 B.n223 10.6151
R893 B.n224 B.n69 10.6151
R894 B.n228 B.n69 10.6151
R895 B.n229 B.n228 10.6151
R896 B.n230 B.n229 10.6151
R897 B.n139 B.n138 10.6151
R898 B.n138 B.n103 10.6151
R899 B.n134 B.n103 10.6151
R900 B.n134 B.n133 10.6151
R901 B.n133 B.n132 10.6151
R902 B.n132 B.n105 10.6151
R903 B.n128 B.n105 10.6151
R904 B.n128 B.n127 10.6151
R905 B.n127 B.n126 10.6151
R906 B.n126 B.n107 10.6151
R907 B.n122 B.n107 10.6151
R908 B.n122 B.n121 10.6151
R909 B.n121 B.n120 10.6151
R910 B.n120 B.n109 10.6151
R911 B.n116 B.n109 10.6151
R912 B.n116 B.n115 10.6151
R913 B.n115 B.n114 10.6151
R914 B.n114 B.n111 10.6151
R915 B.n111 B.n0 10.6151
R916 B.n411 B.n1 10.6151
R917 B.n411 B.n410 10.6151
R918 B.n410 B.n409 10.6151
R919 B.n409 B.n4 10.6151
R920 B.n405 B.n4 10.6151
R921 B.n405 B.n404 10.6151
R922 B.n404 B.n403 10.6151
R923 B.n403 B.n6 10.6151
R924 B.n399 B.n6 10.6151
R925 B.n399 B.n398 10.6151
R926 B.n398 B.n397 10.6151
R927 B.n397 B.n8 10.6151
R928 B.n393 B.n8 10.6151
R929 B.n393 B.n392 10.6151
R930 B.n392 B.n391 10.6151
R931 B.n391 B.n10 10.6151
R932 B.n387 B.n10 10.6151
R933 B.n387 B.n386 10.6151
R934 B.n386 B.n385 10.6151
R935 B.n28 B.n24 9.36635
R936 B.n331 B.n330 9.36635
R937 B.n176 B.n89 9.36635
R938 B.n194 B.n193 9.36635
R939 B.n415 B.n0 2.81026
R940 B.n415 B.n1 2.81026
R941 B.n345 B.n28 1.24928
R942 B.n332 B.n331 1.24928
R943 B.n179 B.n89 1.24928
R944 B.n193 B.n192 1.24928
R945 VN VN.t1 191.137
R946 VN VN.t0 153.204
R947 VDD2.n65 VDD2.n64 756.745
R948 VDD2.n32 VDD2.n31 756.745
R949 VDD2.n64 VDD2.n63 585
R950 VDD2.n35 VDD2.n34 585
R951 VDD2.n58 VDD2.n57 585
R952 VDD2.n56 VDD2.n55 585
R953 VDD2.n39 VDD2.n38 585
R954 VDD2.n50 VDD2.n49 585
R955 VDD2.n48 VDD2.n47 585
R956 VDD2.n43 VDD2.n42 585
R957 VDD2.n10 VDD2.n9 585
R958 VDD2.n15 VDD2.n14 585
R959 VDD2.n17 VDD2.n16 585
R960 VDD2.n6 VDD2.n5 585
R961 VDD2.n23 VDD2.n22 585
R962 VDD2.n25 VDD2.n24 585
R963 VDD2.n2 VDD2.n1 585
R964 VDD2.n31 VDD2.n30 585
R965 VDD2.n44 VDD2.t0 329.084
R966 VDD2.n11 VDD2.t1 329.084
R967 VDD2.n64 VDD2.n34 171.744
R968 VDD2.n57 VDD2.n34 171.744
R969 VDD2.n57 VDD2.n56 171.744
R970 VDD2.n56 VDD2.n38 171.744
R971 VDD2.n49 VDD2.n38 171.744
R972 VDD2.n49 VDD2.n48 171.744
R973 VDD2.n48 VDD2.n42 171.744
R974 VDD2.n15 VDD2.n9 171.744
R975 VDD2.n16 VDD2.n15 171.744
R976 VDD2.n16 VDD2.n5 171.744
R977 VDD2.n23 VDD2.n5 171.744
R978 VDD2.n24 VDD2.n23 171.744
R979 VDD2.n24 VDD2.n1 171.744
R980 VDD2.n31 VDD2.n1 171.744
R981 VDD2.t0 VDD2.n42 85.8723
R982 VDD2.t1 VDD2.n9 85.8723
R983 VDD2.n66 VDD2.n32 83.4802
R984 VDD2.n66 VDD2.n65 50.8035
R985 VDD2.n63 VDD2.n33 12.8005
R986 VDD2.n30 VDD2.n0 12.8005
R987 VDD2.n62 VDD2.n35 12.0247
R988 VDD2.n29 VDD2.n2 12.0247
R989 VDD2.n59 VDD2.n58 11.249
R990 VDD2.n26 VDD2.n25 11.249
R991 VDD2.n44 VDD2.n43 10.7233
R992 VDD2.n11 VDD2.n10 10.7233
R993 VDD2.n55 VDD2.n37 10.4732
R994 VDD2.n22 VDD2.n4 10.4732
R995 VDD2.n54 VDD2.n39 9.69747
R996 VDD2.n21 VDD2.n6 9.69747
R997 VDD2.n61 VDD2.n33 9.45567
R998 VDD2.n28 VDD2.n0 9.45567
R999 VDD2.n62 VDD2.n61 9.3005
R1000 VDD2.n60 VDD2.n59 9.3005
R1001 VDD2.n37 VDD2.n36 9.3005
R1002 VDD2.n54 VDD2.n53 9.3005
R1003 VDD2.n52 VDD2.n51 9.3005
R1004 VDD2.n41 VDD2.n40 9.3005
R1005 VDD2.n46 VDD2.n45 9.3005
R1006 VDD2.n13 VDD2.n12 9.3005
R1007 VDD2.n8 VDD2.n7 9.3005
R1008 VDD2.n19 VDD2.n18 9.3005
R1009 VDD2.n21 VDD2.n20 9.3005
R1010 VDD2.n4 VDD2.n3 9.3005
R1011 VDD2.n27 VDD2.n26 9.3005
R1012 VDD2.n29 VDD2.n28 9.3005
R1013 VDD2.n51 VDD2.n50 8.92171
R1014 VDD2.n18 VDD2.n17 8.92171
R1015 VDD2.n47 VDD2.n41 8.14595
R1016 VDD2.n14 VDD2.n8 8.14595
R1017 VDD2.n46 VDD2.n43 7.3702
R1018 VDD2.n13 VDD2.n10 7.3702
R1019 VDD2.n47 VDD2.n46 5.81868
R1020 VDD2.n14 VDD2.n13 5.81868
R1021 VDD2.n50 VDD2.n41 5.04292
R1022 VDD2.n17 VDD2.n8 5.04292
R1023 VDD2.n51 VDD2.n39 4.26717
R1024 VDD2.n18 VDD2.n6 4.26717
R1025 VDD2.n55 VDD2.n54 3.49141
R1026 VDD2.n22 VDD2.n21 3.49141
R1027 VDD2.n58 VDD2.n37 2.71565
R1028 VDD2.n25 VDD2.n4 2.71565
R1029 VDD2.n45 VDD2.n44 2.41347
R1030 VDD2.n12 VDD2.n11 2.41347
R1031 VDD2.n59 VDD2.n35 1.93989
R1032 VDD2.n26 VDD2.n2 1.93989
R1033 VDD2.n63 VDD2.n62 1.16414
R1034 VDD2.n30 VDD2.n29 1.16414
R1035 VDD2 VDD2.n66 0.487569
R1036 VDD2.n65 VDD2.n33 0.388379
R1037 VDD2.n32 VDD2.n0 0.388379
R1038 VDD2.n61 VDD2.n60 0.155672
R1039 VDD2.n60 VDD2.n36 0.155672
R1040 VDD2.n53 VDD2.n36 0.155672
R1041 VDD2.n53 VDD2.n52 0.155672
R1042 VDD2.n52 VDD2.n40 0.155672
R1043 VDD2.n45 VDD2.n40 0.155672
R1044 VDD2.n12 VDD2.n7 0.155672
R1045 VDD2.n19 VDD2.n7 0.155672
R1046 VDD2.n20 VDD2.n19 0.155672
R1047 VDD2.n20 VDD2.n3 0.155672
R1048 VDD2.n27 VDD2.n3 0.155672
R1049 VDD2.n28 VDD2.n27 0.155672
C0 VP VN 3.9929f
C1 VN B 0.827371f
C2 VP B 1.1901f
C3 VDD1 VTAIL 3.43898f
C4 VTAIL VDD2 3.48382f
C5 VDD1 VDD2 0.563269f
C6 w_n1766_n2264# VTAIL 1.9595f
C7 VDD1 w_n1766_n2264# 1.28384f
C8 w_n1766_n2264# VDD2 1.29845f
C9 VN VTAIL 1.39686f
C10 VDD1 VN 0.148025f
C11 VP VTAIL 1.41112f
C12 VTAIL B 2.09563f
C13 VN VDD2 1.49577f
C14 VP VDD1 1.63931f
C15 VDD1 B 1.1493f
C16 VP VDD2 0.293422f
C17 VDD2 B 1.17107f
C18 w_n1766_n2264# VN 2.25988f
C19 VP w_n1766_n2264# 2.48281f
C20 w_n1766_n2264# B 6.24976f
C21 VDD2 VSUBS 0.60787f
C22 VDD1 VSUBS 2.126272f
C23 VTAIL VSUBS 0.511168f
C24 VN VSUBS 5.04424f
C25 VP VSUBS 1.11989f
C26 B VSUBS 2.732141f
C27 w_n1766_n2264# VSUBS 49.8224f
C28 VDD2.n0 VSUBS 0.008175f
C29 VDD2.n1 VSUBS 0.018475f
C30 VDD2.n2 VSUBS 0.008276f
C31 VDD2.n3 VSUBS 0.014546f
C32 VDD2.n4 VSUBS 0.007817f
C33 VDD2.n5 VSUBS 0.018475f
C34 VDD2.n6 VSUBS 0.008276f
C35 VDD2.n7 VSUBS 0.014546f
C36 VDD2.n8 VSUBS 0.007817f
C37 VDD2.n9 VSUBS 0.013857f
C38 VDD2.n10 VSUBS 0.013896f
C39 VDD2.t1 VSUBS 0.039698f
C40 VDD2.n11 VSUBS 0.07838f
C41 VDD2.n12 VSUBS 0.362599f
C42 VDD2.n13 VSUBS 0.007817f
C43 VDD2.n14 VSUBS 0.008276f
C44 VDD2.n15 VSUBS 0.018475f
C45 VDD2.n16 VSUBS 0.018475f
C46 VDD2.n17 VSUBS 0.008276f
C47 VDD2.n18 VSUBS 0.007817f
C48 VDD2.n19 VSUBS 0.014546f
C49 VDD2.n20 VSUBS 0.014546f
C50 VDD2.n21 VSUBS 0.007817f
C51 VDD2.n22 VSUBS 0.008276f
C52 VDD2.n23 VSUBS 0.018475f
C53 VDD2.n24 VSUBS 0.018475f
C54 VDD2.n25 VSUBS 0.008276f
C55 VDD2.n26 VSUBS 0.007817f
C56 VDD2.n27 VSUBS 0.014546f
C57 VDD2.n28 VSUBS 0.036008f
C58 VDD2.n29 VSUBS 0.007817f
C59 VDD2.n30 VSUBS 0.008276f
C60 VDD2.n31 VSUBS 0.040319f
C61 VDD2.n32 VSUBS 0.286745f
C62 VDD2.n33 VSUBS 0.008175f
C63 VDD2.n34 VSUBS 0.018475f
C64 VDD2.n35 VSUBS 0.008276f
C65 VDD2.n36 VSUBS 0.014546f
C66 VDD2.n37 VSUBS 0.007817f
C67 VDD2.n38 VSUBS 0.018475f
C68 VDD2.n39 VSUBS 0.008276f
C69 VDD2.n40 VSUBS 0.014546f
C70 VDD2.n41 VSUBS 0.007817f
C71 VDD2.n42 VSUBS 0.013857f
C72 VDD2.n43 VSUBS 0.013896f
C73 VDD2.t0 VSUBS 0.039698f
C74 VDD2.n44 VSUBS 0.07838f
C75 VDD2.n45 VSUBS 0.362599f
C76 VDD2.n46 VSUBS 0.007817f
C77 VDD2.n47 VSUBS 0.008276f
C78 VDD2.n48 VSUBS 0.018475f
C79 VDD2.n49 VSUBS 0.018475f
C80 VDD2.n50 VSUBS 0.008276f
C81 VDD2.n51 VSUBS 0.007817f
C82 VDD2.n52 VSUBS 0.014546f
C83 VDD2.n53 VSUBS 0.014546f
C84 VDD2.n54 VSUBS 0.007817f
C85 VDD2.n55 VSUBS 0.008276f
C86 VDD2.n56 VSUBS 0.018475f
C87 VDD2.n57 VSUBS 0.018475f
C88 VDD2.n58 VSUBS 0.008276f
C89 VDD2.n59 VSUBS 0.007817f
C90 VDD2.n60 VSUBS 0.014546f
C91 VDD2.n61 VSUBS 0.036008f
C92 VDD2.n62 VSUBS 0.007817f
C93 VDD2.n63 VSUBS 0.008276f
C94 VDD2.n64 VSUBS 0.040319f
C95 VDD2.n65 VSUBS 0.03646f
C96 VDD2.n66 VSUBS 1.33503f
C97 VN.t0 VSUBS 1.32803f
C98 VN.t1 VSUBS 1.68599f
C99 B.n0 VSUBS 0.005017f
C100 B.n1 VSUBS 0.005017f
C101 B.n2 VSUBS 0.007934f
C102 B.n3 VSUBS 0.007934f
C103 B.n4 VSUBS 0.007934f
C104 B.n5 VSUBS 0.007934f
C105 B.n6 VSUBS 0.007934f
C106 B.n7 VSUBS 0.007934f
C107 B.n8 VSUBS 0.007934f
C108 B.n9 VSUBS 0.007934f
C109 B.n10 VSUBS 0.007934f
C110 B.n11 VSUBS 0.007934f
C111 B.n12 VSUBS 0.018607f
C112 B.n13 VSUBS 0.007934f
C113 B.n14 VSUBS 0.007934f
C114 B.n15 VSUBS 0.007934f
C115 B.n16 VSUBS 0.007934f
C116 B.n17 VSUBS 0.007934f
C117 B.n18 VSUBS 0.007934f
C118 B.n19 VSUBS 0.007934f
C119 B.n20 VSUBS 0.007934f
C120 B.n21 VSUBS 0.007934f
C121 B.n22 VSUBS 0.007934f
C122 B.n23 VSUBS 0.007934f
C123 B.n24 VSUBS 0.007467f
C124 B.n25 VSUBS 0.007934f
C125 B.t2 VSUBS 0.110645f
C126 B.t1 VSUBS 0.131728f
C127 B.t0 VSUBS 0.55968f
C128 B.n26 VSUBS 0.228342f
C129 B.n27 VSUBS 0.183339f
C130 B.n28 VSUBS 0.018381f
C131 B.n29 VSUBS 0.007934f
C132 B.n30 VSUBS 0.007934f
C133 B.n31 VSUBS 0.007934f
C134 B.n32 VSUBS 0.007934f
C135 B.t5 VSUBS 0.110648f
C136 B.t4 VSUBS 0.13173f
C137 B.t3 VSUBS 0.55968f
C138 B.n33 VSUBS 0.22834f
C139 B.n34 VSUBS 0.183337f
C140 B.n35 VSUBS 0.007934f
C141 B.n36 VSUBS 0.007934f
C142 B.n37 VSUBS 0.007934f
C143 B.n38 VSUBS 0.007934f
C144 B.n39 VSUBS 0.007934f
C145 B.n40 VSUBS 0.007934f
C146 B.n41 VSUBS 0.007934f
C147 B.n42 VSUBS 0.007934f
C148 B.n43 VSUBS 0.007934f
C149 B.n44 VSUBS 0.007934f
C150 B.n45 VSUBS 0.007934f
C151 B.n46 VSUBS 0.007934f
C152 B.n47 VSUBS 0.019208f
C153 B.n48 VSUBS 0.007934f
C154 B.n49 VSUBS 0.007934f
C155 B.n50 VSUBS 0.007934f
C156 B.n51 VSUBS 0.007934f
C157 B.n52 VSUBS 0.007934f
C158 B.n53 VSUBS 0.007934f
C159 B.n54 VSUBS 0.007934f
C160 B.n55 VSUBS 0.007934f
C161 B.n56 VSUBS 0.007934f
C162 B.n57 VSUBS 0.007934f
C163 B.n58 VSUBS 0.007934f
C164 B.n59 VSUBS 0.007934f
C165 B.n60 VSUBS 0.007934f
C166 B.n61 VSUBS 0.007934f
C167 B.n62 VSUBS 0.007934f
C168 B.n63 VSUBS 0.007934f
C169 B.n64 VSUBS 0.007934f
C170 B.n65 VSUBS 0.007934f
C171 B.n66 VSUBS 0.007934f
C172 B.n67 VSUBS 0.018261f
C173 B.n68 VSUBS 0.007934f
C174 B.n69 VSUBS 0.007934f
C175 B.n70 VSUBS 0.007934f
C176 B.n71 VSUBS 0.007934f
C177 B.n72 VSUBS 0.007934f
C178 B.n73 VSUBS 0.007934f
C179 B.n74 VSUBS 0.007934f
C180 B.n75 VSUBS 0.007934f
C181 B.n76 VSUBS 0.007934f
C182 B.n77 VSUBS 0.007934f
C183 B.n78 VSUBS 0.007934f
C184 B.n79 VSUBS 0.007934f
C185 B.n80 VSUBS 0.007934f
C186 B.t10 VSUBS 0.110648f
C187 B.t11 VSUBS 0.13173f
C188 B.t9 VSUBS 0.55968f
C189 B.n81 VSUBS 0.22834f
C190 B.n82 VSUBS 0.183337f
C191 B.n83 VSUBS 0.007934f
C192 B.n84 VSUBS 0.007934f
C193 B.n85 VSUBS 0.007934f
C194 B.n86 VSUBS 0.007934f
C195 B.t7 VSUBS 0.110645f
C196 B.t8 VSUBS 0.131728f
C197 B.t6 VSUBS 0.55968f
C198 B.n87 VSUBS 0.228342f
C199 B.n88 VSUBS 0.183339f
C200 B.n89 VSUBS 0.018381f
C201 B.n90 VSUBS 0.007934f
C202 B.n91 VSUBS 0.007934f
C203 B.n92 VSUBS 0.007934f
C204 B.n93 VSUBS 0.007934f
C205 B.n94 VSUBS 0.007934f
C206 B.n95 VSUBS 0.007934f
C207 B.n96 VSUBS 0.007934f
C208 B.n97 VSUBS 0.007934f
C209 B.n98 VSUBS 0.007934f
C210 B.n99 VSUBS 0.007934f
C211 B.n100 VSUBS 0.007934f
C212 B.n101 VSUBS 0.007934f
C213 B.n102 VSUBS 0.018261f
C214 B.n103 VSUBS 0.007934f
C215 B.n104 VSUBS 0.007934f
C216 B.n105 VSUBS 0.007934f
C217 B.n106 VSUBS 0.007934f
C218 B.n107 VSUBS 0.007934f
C219 B.n108 VSUBS 0.007934f
C220 B.n109 VSUBS 0.007934f
C221 B.n110 VSUBS 0.007934f
C222 B.n111 VSUBS 0.007934f
C223 B.n112 VSUBS 0.007934f
C224 B.n113 VSUBS 0.007934f
C225 B.n114 VSUBS 0.007934f
C226 B.n115 VSUBS 0.007934f
C227 B.n116 VSUBS 0.007934f
C228 B.n117 VSUBS 0.007934f
C229 B.n118 VSUBS 0.007934f
C230 B.n119 VSUBS 0.007934f
C231 B.n120 VSUBS 0.007934f
C232 B.n121 VSUBS 0.007934f
C233 B.n122 VSUBS 0.007934f
C234 B.n123 VSUBS 0.007934f
C235 B.n124 VSUBS 0.007934f
C236 B.n125 VSUBS 0.007934f
C237 B.n126 VSUBS 0.007934f
C238 B.n127 VSUBS 0.007934f
C239 B.n128 VSUBS 0.007934f
C240 B.n129 VSUBS 0.007934f
C241 B.n130 VSUBS 0.007934f
C242 B.n131 VSUBS 0.007934f
C243 B.n132 VSUBS 0.007934f
C244 B.n133 VSUBS 0.007934f
C245 B.n134 VSUBS 0.007934f
C246 B.n135 VSUBS 0.007934f
C247 B.n136 VSUBS 0.007934f
C248 B.n137 VSUBS 0.007934f
C249 B.n138 VSUBS 0.007934f
C250 B.n139 VSUBS 0.018261f
C251 B.n140 VSUBS 0.018607f
C252 B.n141 VSUBS 0.018607f
C253 B.n142 VSUBS 0.007934f
C254 B.n143 VSUBS 0.007934f
C255 B.n144 VSUBS 0.007934f
C256 B.n145 VSUBS 0.007934f
C257 B.n146 VSUBS 0.007934f
C258 B.n147 VSUBS 0.007934f
C259 B.n148 VSUBS 0.007934f
C260 B.n149 VSUBS 0.007934f
C261 B.n150 VSUBS 0.007934f
C262 B.n151 VSUBS 0.007934f
C263 B.n152 VSUBS 0.007934f
C264 B.n153 VSUBS 0.007934f
C265 B.n154 VSUBS 0.007934f
C266 B.n155 VSUBS 0.007934f
C267 B.n156 VSUBS 0.007934f
C268 B.n157 VSUBS 0.007934f
C269 B.n158 VSUBS 0.007934f
C270 B.n159 VSUBS 0.007934f
C271 B.n160 VSUBS 0.007934f
C272 B.n161 VSUBS 0.007934f
C273 B.n162 VSUBS 0.007934f
C274 B.n163 VSUBS 0.007934f
C275 B.n164 VSUBS 0.007934f
C276 B.n165 VSUBS 0.007934f
C277 B.n166 VSUBS 0.007934f
C278 B.n167 VSUBS 0.007934f
C279 B.n168 VSUBS 0.007934f
C280 B.n169 VSUBS 0.007934f
C281 B.n170 VSUBS 0.007934f
C282 B.n171 VSUBS 0.007934f
C283 B.n172 VSUBS 0.007934f
C284 B.n173 VSUBS 0.007934f
C285 B.n174 VSUBS 0.007934f
C286 B.n175 VSUBS 0.007934f
C287 B.n176 VSUBS 0.007467f
C288 B.n177 VSUBS 0.007934f
C289 B.n178 VSUBS 0.007934f
C290 B.n179 VSUBS 0.004433f
C291 B.n180 VSUBS 0.007934f
C292 B.n181 VSUBS 0.007934f
C293 B.n182 VSUBS 0.007934f
C294 B.n183 VSUBS 0.007934f
C295 B.n184 VSUBS 0.007934f
C296 B.n185 VSUBS 0.007934f
C297 B.n186 VSUBS 0.007934f
C298 B.n187 VSUBS 0.007934f
C299 B.n188 VSUBS 0.007934f
C300 B.n189 VSUBS 0.007934f
C301 B.n190 VSUBS 0.007934f
C302 B.n191 VSUBS 0.007934f
C303 B.n192 VSUBS 0.004433f
C304 B.n193 VSUBS 0.018381f
C305 B.n194 VSUBS 0.007467f
C306 B.n195 VSUBS 0.007934f
C307 B.n196 VSUBS 0.007934f
C308 B.n197 VSUBS 0.007934f
C309 B.n198 VSUBS 0.007934f
C310 B.n199 VSUBS 0.007934f
C311 B.n200 VSUBS 0.007934f
C312 B.n201 VSUBS 0.007934f
C313 B.n202 VSUBS 0.007934f
C314 B.n203 VSUBS 0.007934f
C315 B.n204 VSUBS 0.007934f
C316 B.n205 VSUBS 0.007934f
C317 B.n206 VSUBS 0.007934f
C318 B.n207 VSUBS 0.007934f
C319 B.n208 VSUBS 0.007934f
C320 B.n209 VSUBS 0.007934f
C321 B.n210 VSUBS 0.007934f
C322 B.n211 VSUBS 0.007934f
C323 B.n212 VSUBS 0.007934f
C324 B.n213 VSUBS 0.007934f
C325 B.n214 VSUBS 0.007934f
C326 B.n215 VSUBS 0.007934f
C327 B.n216 VSUBS 0.007934f
C328 B.n217 VSUBS 0.007934f
C329 B.n218 VSUBS 0.007934f
C330 B.n219 VSUBS 0.007934f
C331 B.n220 VSUBS 0.007934f
C332 B.n221 VSUBS 0.007934f
C333 B.n222 VSUBS 0.007934f
C334 B.n223 VSUBS 0.007934f
C335 B.n224 VSUBS 0.007934f
C336 B.n225 VSUBS 0.007934f
C337 B.n226 VSUBS 0.007934f
C338 B.n227 VSUBS 0.007934f
C339 B.n228 VSUBS 0.007934f
C340 B.n229 VSUBS 0.007934f
C341 B.n230 VSUBS 0.018607f
C342 B.n231 VSUBS 0.018607f
C343 B.n232 VSUBS 0.018261f
C344 B.n233 VSUBS 0.007934f
C345 B.n234 VSUBS 0.007934f
C346 B.n235 VSUBS 0.007934f
C347 B.n236 VSUBS 0.007934f
C348 B.n237 VSUBS 0.007934f
C349 B.n238 VSUBS 0.007934f
C350 B.n239 VSUBS 0.007934f
C351 B.n240 VSUBS 0.007934f
C352 B.n241 VSUBS 0.007934f
C353 B.n242 VSUBS 0.007934f
C354 B.n243 VSUBS 0.007934f
C355 B.n244 VSUBS 0.007934f
C356 B.n245 VSUBS 0.007934f
C357 B.n246 VSUBS 0.007934f
C358 B.n247 VSUBS 0.007934f
C359 B.n248 VSUBS 0.007934f
C360 B.n249 VSUBS 0.007934f
C361 B.n250 VSUBS 0.007934f
C362 B.n251 VSUBS 0.007934f
C363 B.n252 VSUBS 0.007934f
C364 B.n253 VSUBS 0.007934f
C365 B.n254 VSUBS 0.007934f
C366 B.n255 VSUBS 0.007934f
C367 B.n256 VSUBS 0.007934f
C368 B.n257 VSUBS 0.007934f
C369 B.n258 VSUBS 0.007934f
C370 B.n259 VSUBS 0.007934f
C371 B.n260 VSUBS 0.007934f
C372 B.n261 VSUBS 0.007934f
C373 B.n262 VSUBS 0.007934f
C374 B.n263 VSUBS 0.007934f
C375 B.n264 VSUBS 0.007934f
C376 B.n265 VSUBS 0.007934f
C377 B.n266 VSUBS 0.007934f
C378 B.n267 VSUBS 0.007934f
C379 B.n268 VSUBS 0.007934f
C380 B.n269 VSUBS 0.007934f
C381 B.n270 VSUBS 0.007934f
C382 B.n271 VSUBS 0.007934f
C383 B.n272 VSUBS 0.007934f
C384 B.n273 VSUBS 0.007934f
C385 B.n274 VSUBS 0.007934f
C386 B.n275 VSUBS 0.007934f
C387 B.n276 VSUBS 0.007934f
C388 B.n277 VSUBS 0.007934f
C389 B.n278 VSUBS 0.007934f
C390 B.n279 VSUBS 0.007934f
C391 B.n280 VSUBS 0.007934f
C392 B.n281 VSUBS 0.007934f
C393 B.n282 VSUBS 0.007934f
C394 B.n283 VSUBS 0.007934f
C395 B.n284 VSUBS 0.007934f
C396 B.n285 VSUBS 0.007934f
C397 B.n286 VSUBS 0.007934f
C398 B.n287 VSUBS 0.007934f
C399 B.n288 VSUBS 0.007934f
C400 B.n289 VSUBS 0.007934f
C401 B.n290 VSUBS 0.007934f
C402 B.n291 VSUBS 0.007934f
C403 B.n292 VSUBS 0.018261f
C404 B.n293 VSUBS 0.018607f
C405 B.n294 VSUBS 0.01766f
C406 B.n295 VSUBS 0.007934f
C407 B.n296 VSUBS 0.007934f
C408 B.n297 VSUBS 0.007934f
C409 B.n298 VSUBS 0.007934f
C410 B.n299 VSUBS 0.007934f
C411 B.n300 VSUBS 0.007934f
C412 B.n301 VSUBS 0.007934f
C413 B.n302 VSUBS 0.007934f
C414 B.n303 VSUBS 0.007934f
C415 B.n304 VSUBS 0.007934f
C416 B.n305 VSUBS 0.007934f
C417 B.n306 VSUBS 0.007934f
C418 B.n307 VSUBS 0.007934f
C419 B.n308 VSUBS 0.007934f
C420 B.n309 VSUBS 0.007934f
C421 B.n310 VSUBS 0.007934f
C422 B.n311 VSUBS 0.007934f
C423 B.n312 VSUBS 0.007934f
C424 B.n313 VSUBS 0.007934f
C425 B.n314 VSUBS 0.007934f
C426 B.n315 VSUBS 0.007934f
C427 B.n316 VSUBS 0.007934f
C428 B.n317 VSUBS 0.007934f
C429 B.n318 VSUBS 0.007934f
C430 B.n319 VSUBS 0.007934f
C431 B.n320 VSUBS 0.007934f
C432 B.n321 VSUBS 0.007934f
C433 B.n322 VSUBS 0.007934f
C434 B.n323 VSUBS 0.007934f
C435 B.n324 VSUBS 0.007934f
C436 B.n325 VSUBS 0.007934f
C437 B.n326 VSUBS 0.007934f
C438 B.n327 VSUBS 0.007934f
C439 B.n328 VSUBS 0.007934f
C440 B.n329 VSUBS 0.007934f
C441 B.n330 VSUBS 0.007467f
C442 B.n331 VSUBS 0.018381f
C443 B.n332 VSUBS 0.004433f
C444 B.n333 VSUBS 0.007934f
C445 B.n334 VSUBS 0.007934f
C446 B.n335 VSUBS 0.007934f
C447 B.n336 VSUBS 0.007934f
C448 B.n337 VSUBS 0.007934f
C449 B.n338 VSUBS 0.007934f
C450 B.n339 VSUBS 0.007934f
C451 B.n340 VSUBS 0.007934f
C452 B.n341 VSUBS 0.007934f
C453 B.n342 VSUBS 0.007934f
C454 B.n343 VSUBS 0.007934f
C455 B.n344 VSUBS 0.007934f
C456 B.n345 VSUBS 0.004433f
C457 B.n346 VSUBS 0.007934f
C458 B.n347 VSUBS 0.007934f
C459 B.n348 VSUBS 0.007934f
C460 B.n349 VSUBS 0.007934f
C461 B.n350 VSUBS 0.007934f
C462 B.n351 VSUBS 0.007934f
C463 B.n352 VSUBS 0.007934f
C464 B.n353 VSUBS 0.007934f
C465 B.n354 VSUBS 0.007934f
C466 B.n355 VSUBS 0.007934f
C467 B.n356 VSUBS 0.007934f
C468 B.n357 VSUBS 0.007934f
C469 B.n358 VSUBS 0.007934f
C470 B.n359 VSUBS 0.007934f
C471 B.n360 VSUBS 0.007934f
C472 B.n361 VSUBS 0.007934f
C473 B.n362 VSUBS 0.007934f
C474 B.n363 VSUBS 0.007934f
C475 B.n364 VSUBS 0.007934f
C476 B.n365 VSUBS 0.007934f
C477 B.n366 VSUBS 0.007934f
C478 B.n367 VSUBS 0.007934f
C479 B.n368 VSUBS 0.007934f
C480 B.n369 VSUBS 0.007934f
C481 B.n370 VSUBS 0.007934f
C482 B.n371 VSUBS 0.007934f
C483 B.n372 VSUBS 0.007934f
C484 B.n373 VSUBS 0.007934f
C485 B.n374 VSUBS 0.007934f
C486 B.n375 VSUBS 0.007934f
C487 B.n376 VSUBS 0.007934f
C488 B.n377 VSUBS 0.007934f
C489 B.n378 VSUBS 0.007934f
C490 B.n379 VSUBS 0.007934f
C491 B.n380 VSUBS 0.007934f
C492 B.n381 VSUBS 0.007934f
C493 B.n382 VSUBS 0.007934f
C494 B.n383 VSUBS 0.018607f
C495 B.n384 VSUBS 0.018261f
C496 B.n385 VSUBS 0.018261f
C497 B.n386 VSUBS 0.007934f
C498 B.n387 VSUBS 0.007934f
C499 B.n388 VSUBS 0.007934f
C500 B.n389 VSUBS 0.007934f
C501 B.n390 VSUBS 0.007934f
C502 B.n391 VSUBS 0.007934f
C503 B.n392 VSUBS 0.007934f
C504 B.n393 VSUBS 0.007934f
C505 B.n394 VSUBS 0.007934f
C506 B.n395 VSUBS 0.007934f
C507 B.n396 VSUBS 0.007934f
C508 B.n397 VSUBS 0.007934f
C509 B.n398 VSUBS 0.007934f
C510 B.n399 VSUBS 0.007934f
C511 B.n400 VSUBS 0.007934f
C512 B.n401 VSUBS 0.007934f
C513 B.n402 VSUBS 0.007934f
C514 B.n403 VSUBS 0.007934f
C515 B.n404 VSUBS 0.007934f
C516 B.n405 VSUBS 0.007934f
C517 B.n406 VSUBS 0.007934f
C518 B.n407 VSUBS 0.007934f
C519 B.n408 VSUBS 0.007934f
C520 B.n409 VSUBS 0.007934f
C521 B.n410 VSUBS 0.007934f
C522 B.n411 VSUBS 0.007934f
C523 B.n412 VSUBS 0.007934f
C524 B.n413 VSUBS 0.007934f
C525 B.n414 VSUBS 0.007934f
C526 B.n415 VSUBS 0.017964f
C527 VDD1.n0 VSUBS 0.007821f
C528 VDD1.n1 VSUBS 0.017676f
C529 VDD1.n2 VSUBS 0.007918f
C530 VDD1.n3 VSUBS 0.013917f
C531 VDD1.n4 VSUBS 0.007478f
C532 VDD1.n5 VSUBS 0.017676f
C533 VDD1.n6 VSUBS 0.007918f
C534 VDD1.n7 VSUBS 0.013917f
C535 VDD1.n8 VSUBS 0.007478f
C536 VDD1.n9 VSUBS 0.013257f
C537 VDD1.n10 VSUBS 0.013295f
C538 VDD1.t1 VSUBS 0.037981f
C539 VDD1.n11 VSUBS 0.074989f
C540 VDD1.n12 VSUBS 0.346914f
C541 VDD1.n13 VSUBS 0.007478f
C542 VDD1.n14 VSUBS 0.007918f
C543 VDD1.n15 VSUBS 0.017676f
C544 VDD1.n16 VSUBS 0.017676f
C545 VDD1.n17 VSUBS 0.007918f
C546 VDD1.n18 VSUBS 0.007478f
C547 VDD1.n19 VSUBS 0.013917f
C548 VDD1.n20 VSUBS 0.013917f
C549 VDD1.n21 VSUBS 0.007478f
C550 VDD1.n22 VSUBS 0.007918f
C551 VDD1.n23 VSUBS 0.017676f
C552 VDD1.n24 VSUBS 0.017676f
C553 VDD1.n25 VSUBS 0.007918f
C554 VDD1.n26 VSUBS 0.007478f
C555 VDD1.n27 VSUBS 0.013917f
C556 VDD1.n28 VSUBS 0.03445f
C557 VDD1.n29 VSUBS 0.007478f
C558 VDD1.n30 VSUBS 0.007918f
C559 VDD1.n31 VSUBS 0.038575f
C560 VDD1.n32 VSUBS 0.035355f
C561 VDD1.n33 VSUBS 0.007821f
C562 VDD1.n34 VSUBS 0.017676f
C563 VDD1.n35 VSUBS 0.007918f
C564 VDD1.n36 VSUBS 0.013917f
C565 VDD1.n37 VSUBS 0.007478f
C566 VDD1.n38 VSUBS 0.017676f
C567 VDD1.n39 VSUBS 0.007918f
C568 VDD1.n40 VSUBS 0.013917f
C569 VDD1.n41 VSUBS 0.007478f
C570 VDD1.n42 VSUBS 0.013257f
C571 VDD1.n43 VSUBS 0.013295f
C572 VDD1.t0 VSUBS 0.037981f
C573 VDD1.n44 VSUBS 0.074989f
C574 VDD1.n45 VSUBS 0.346914f
C575 VDD1.n46 VSUBS 0.007478f
C576 VDD1.n47 VSUBS 0.007918f
C577 VDD1.n48 VSUBS 0.017676f
C578 VDD1.n49 VSUBS 0.017676f
C579 VDD1.n50 VSUBS 0.007918f
C580 VDD1.n51 VSUBS 0.007478f
C581 VDD1.n52 VSUBS 0.013917f
C582 VDD1.n53 VSUBS 0.013917f
C583 VDD1.n54 VSUBS 0.007478f
C584 VDD1.n55 VSUBS 0.007918f
C585 VDD1.n56 VSUBS 0.017676f
C586 VDD1.n57 VSUBS 0.017676f
C587 VDD1.n58 VSUBS 0.007918f
C588 VDD1.n59 VSUBS 0.007478f
C589 VDD1.n60 VSUBS 0.013917f
C590 VDD1.n61 VSUBS 0.03445f
C591 VDD1.n62 VSUBS 0.007478f
C592 VDD1.n63 VSUBS 0.007918f
C593 VDD1.n64 VSUBS 0.038575f
C594 VDD1.n65 VSUBS 0.294362f
C595 VTAIL.n0 VSUBS 0.011705f
C596 VTAIL.n1 VSUBS 0.026454f
C597 VTAIL.n2 VSUBS 0.01185f
C598 VTAIL.n3 VSUBS 0.020828f
C599 VTAIL.n4 VSUBS 0.011192f
C600 VTAIL.n5 VSUBS 0.026454f
C601 VTAIL.n6 VSUBS 0.01185f
C602 VTAIL.n7 VSUBS 0.020828f
C603 VTAIL.n8 VSUBS 0.011192f
C604 VTAIL.n9 VSUBS 0.01984f
C605 VTAIL.n10 VSUBS 0.019897f
C606 VTAIL.t3 VSUBS 0.056841f
C607 VTAIL.n11 VSUBS 0.112228f
C608 VTAIL.n12 VSUBS 0.519183f
C609 VTAIL.n13 VSUBS 0.011192f
C610 VTAIL.n14 VSUBS 0.01185f
C611 VTAIL.n15 VSUBS 0.026454f
C612 VTAIL.n16 VSUBS 0.026454f
C613 VTAIL.n17 VSUBS 0.01185f
C614 VTAIL.n18 VSUBS 0.011192f
C615 VTAIL.n19 VSUBS 0.020828f
C616 VTAIL.n20 VSUBS 0.020828f
C617 VTAIL.n21 VSUBS 0.011192f
C618 VTAIL.n22 VSUBS 0.01185f
C619 VTAIL.n23 VSUBS 0.026454f
C620 VTAIL.n24 VSUBS 0.026454f
C621 VTAIL.n25 VSUBS 0.01185f
C622 VTAIL.n26 VSUBS 0.011192f
C623 VTAIL.n27 VSUBS 0.020828f
C624 VTAIL.n28 VSUBS 0.051557f
C625 VTAIL.n29 VSUBS 0.011192f
C626 VTAIL.n30 VSUBS 0.01185f
C627 VTAIL.n31 VSUBS 0.05773f
C628 VTAIL.n32 VSUBS 0.037845f
C629 VTAIL.n33 VSUBS 0.971704f
C630 VTAIL.n34 VSUBS 0.011705f
C631 VTAIL.n35 VSUBS 0.026454f
C632 VTAIL.n36 VSUBS 0.01185f
C633 VTAIL.n37 VSUBS 0.020828f
C634 VTAIL.n38 VSUBS 0.011192f
C635 VTAIL.n39 VSUBS 0.026454f
C636 VTAIL.n40 VSUBS 0.01185f
C637 VTAIL.n41 VSUBS 0.020828f
C638 VTAIL.n42 VSUBS 0.011192f
C639 VTAIL.n43 VSUBS 0.01984f
C640 VTAIL.n44 VSUBS 0.019897f
C641 VTAIL.t1 VSUBS 0.056841f
C642 VTAIL.n45 VSUBS 0.112228f
C643 VTAIL.n46 VSUBS 0.519183f
C644 VTAIL.n47 VSUBS 0.011192f
C645 VTAIL.n48 VSUBS 0.01185f
C646 VTAIL.n49 VSUBS 0.026454f
C647 VTAIL.n50 VSUBS 0.026454f
C648 VTAIL.n51 VSUBS 0.01185f
C649 VTAIL.n52 VSUBS 0.011192f
C650 VTAIL.n53 VSUBS 0.020828f
C651 VTAIL.n54 VSUBS 0.020828f
C652 VTAIL.n55 VSUBS 0.011192f
C653 VTAIL.n56 VSUBS 0.01185f
C654 VTAIL.n57 VSUBS 0.026454f
C655 VTAIL.n58 VSUBS 0.026454f
C656 VTAIL.n59 VSUBS 0.01185f
C657 VTAIL.n60 VSUBS 0.011192f
C658 VTAIL.n61 VSUBS 0.020828f
C659 VTAIL.n62 VSUBS 0.051557f
C660 VTAIL.n63 VSUBS 0.011192f
C661 VTAIL.n64 VSUBS 0.01185f
C662 VTAIL.n65 VSUBS 0.05773f
C663 VTAIL.n66 VSUBS 0.037845f
C664 VTAIL.n67 VSUBS 0.996581f
C665 VTAIL.n68 VSUBS 0.011705f
C666 VTAIL.n69 VSUBS 0.026454f
C667 VTAIL.n70 VSUBS 0.01185f
C668 VTAIL.n71 VSUBS 0.020828f
C669 VTAIL.n72 VSUBS 0.011192f
C670 VTAIL.n73 VSUBS 0.026454f
C671 VTAIL.n74 VSUBS 0.01185f
C672 VTAIL.n75 VSUBS 0.020828f
C673 VTAIL.n76 VSUBS 0.011192f
C674 VTAIL.n77 VSUBS 0.01984f
C675 VTAIL.n78 VSUBS 0.019897f
C676 VTAIL.t2 VSUBS 0.056841f
C677 VTAIL.n79 VSUBS 0.112228f
C678 VTAIL.n80 VSUBS 0.519183f
C679 VTAIL.n81 VSUBS 0.011192f
C680 VTAIL.n82 VSUBS 0.01185f
C681 VTAIL.n83 VSUBS 0.026454f
C682 VTAIL.n84 VSUBS 0.026454f
C683 VTAIL.n85 VSUBS 0.01185f
C684 VTAIL.n86 VSUBS 0.011192f
C685 VTAIL.n87 VSUBS 0.020828f
C686 VTAIL.n88 VSUBS 0.020828f
C687 VTAIL.n89 VSUBS 0.011192f
C688 VTAIL.n90 VSUBS 0.01185f
C689 VTAIL.n91 VSUBS 0.026454f
C690 VTAIL.n92 VSUBS 0.026454f
C691 VTAIL.n93 VSUBS 0.01185f
C692 VTAIL.n94 VSUBS 0.011192f
C693 VTAIL.n95 VSUBS 0.020828f
C694 VTAIL.n96 VSUBS 0.051557f
C695 VTAIL.n97 VSUBS 0.011192f
C696 VTAIL.n98 VSUBS 0.01185f
C697 VTAIL.n99 VSUBS 0.05773f
C698 VTAIL.n100 VSUBS 0.037845f
C699 VTAIL.n101 VSUBS 0.88145f
C700 VTAIL.n102 VSUBS 0.011705f
C701 VTAIL.n103 VSUBS 0.026454f
C702 VTAIL.n104 VSUBS 0.01185f
C703 VTAIL.n105 VSUBS 0.020828f
C704 VTAIL.n106 VSUBS 0.011192f
C705 VTAIL.n107 VSUBS 0.026454f
C706 VTAIL.n108 VSUBS 0.01185f
C707 VTAIL.n109 VSUBS 0.020828f
C708 VTAIL.n110 VSUBS 0.011192f
C709 VTAIL.n111 VSUBS 0.01984f
C710 VTAIL.n112 VSUBS 0.019897f
C711 VTAIL.t0 VSUBS 0.056841f
C712 VTAIL.n113 VSUBS 0.112228f
C713 VTAIL.n114 VSUBS 0.519183f
C714 VTAIL.n115 VSUBS 0.011192f
C715 VTAIL.n116 VSUBS 0.01185f
C716 VTAIL.n117 VSUBS 0.026454f
C717 VTAIL.n118 VSUBS 0.026454f
C718 VTAIL.n119 VSUBS 0.01185f
C719 VTAIL.n120 VSUBS 0.011192f
C720 VTAIL.n121 VSUBS 0.020828f
C721 VTAIL.n122 VSUBS 0.020828f
C722 VTAIL.n123 VSUBS 0.011192f
C723 VTAIL.n124 VSUBS 0.01185f
C724 VTAIL.n125 VSUBS 0.026454f
C725 VTAIL.n126 VSUBS 0.026454f
C726 VTAIL.n127 VSUBS 0.01185f
C727 VTAIL.n128 VSUBS 0.011192f
C728 VTAIL.n129 VSUBS 0.020828f
C729 VTAIL.n130 VSUBS 0.051557f
C730 VTAIL.n131 VSUBS 0.011192f
C731 VTAIL.n132 VSUBS 0.01185f
C732 VTAIL.n133 VSUBS 0.05773f
C733 VTAIL.n134 VSUBS 0.037845f
C734 VTAIL.n135 VSUBS 0.81723f
C735 VP.t0 VSUBS 1.74922f
C736 VP.t1 VSUBS 1.38126f
C737 VP.n0 VSUBS 3.31329f
.ends

