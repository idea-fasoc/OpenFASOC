* NGSPICE file created from diff_pair_sample_1191.ext - technology: sky130A

.subckt diff_pair_sample_1191 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=2.53
X1 VDD1.t9 VP.t0 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=0.9555 pd=5.68 as=0.40425 ps=2.78 w=2.45 l=2.53
X2 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=2.53
X3 VDD2.t0 VN.t1 VTAIL.t18 B.t4 sky130_fd_pr__nfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=2.53
X4 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=2.53
X5 VTAIL.t17 VN.t2 VDD2.t1 B.t8 sky130_fd_pr__nfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=2.53
X6 VDD2.t2 VN.t3 VTAIL.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=0.9555 pd=5.68 as=0.40425 ps=2.78 w=2.45 l=2.53
X7 VTAIL.t8 VP.t1 VDD1.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=2.53
X8 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=2.53
X9 VDD1.t7 VP.t2 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=2.53
X10 VTAIL.t6 VP.t3 VDD1.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=2.53
X11 VTAIL.t15 VN.t4 VDD2.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=2.53
X12 VDD1.t5 VP.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9555 pd=5.68 as=0.40425 ps=2.78 w=2.45 l=2.53
X13 VDD2.t6 VN.t5 VTAIL.t14 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9555 pd=5.68 as=0.40425 ps=2.78 w=2.45 l=2.53
X14 VDD2.t9 VN.t6 VTAIL.t13 B.t1 sky130_fd_pr__nfet_01v8 ad=0.40425 pd=2.78 as=0.9555 ps=5.68 w=2.45 l=2.53
X15 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=2.53
X16 VDD2.t8 VN.t7 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=2.53
X17 VDD1.t4 VP.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.40425 pd=2.78 as=0.9555 ps=5.68 w=2.45 l=2.53
X18 VTAIL.t0 VP.t6 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=2.53
X19 VDD1.t2 VP.t7 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.40425 pd=2.78 as=0.9555 ps=5.68 w=2.45 l=2.53
X20 VTAIL.t3 VP.t8 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=2.53
X21 VTAIL.t11 VN.t8 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=2.53
X22 VDD2.t3 VN.t9 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=0.40425 pd=2.78 as=0.9555 ps=5.68 w=2.45 l=2.53
X23 VDD1.t0 VP.t9 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=2.53
R0 VN.n75 VN.n39 161.3
R1 VN.n74 VN.n73 161.3
R2 VN.n72 VN.n40 161.3
R3 VN.n71 VN.n70 161.3
R4 VN.n69 VN.n41 161.3
R5 VN.n68 VN.n67 161.3
R6 VN.n66 VN.n65 161.3
R7 VN.n64 VN.n43 161.3
R8 VN.n63 VN.n62 161.3
R9 VN.n61 VN.n44 161.3
R10 VN.n60 VN.n59 161.3
R11 VN.n58 VN.n45 161.3
R12 VN.n57 VN.n56 161.3
R13 VN.n55 VN.n46 161.3
R14 VN.n54 VN.n53 161.3
R15 VN.n52 VN.n47 161.3
R16 VN.n51 VN.n50 161.3
R17 VN.n36 VN.n0 161.3
R18 VN.n35 VN.n34 161.3
R19 VN.n33 VN.n1 161.3
R20 VN.n32 VN.n31 161.3
R21 VN.n30 VN.n2 161.3
R22 VN.n29 VN.n28 161.3
R23 VN.n27 VN.n26 161.3
R24 VN.n25 VN.n4 161.3
R25 VN.n24 VN.n23 161.3
R26 VN.n22 VN.n5 161.3
R27 VN.n21 VN.n20 161.3
R28 VN.n19 VN.n6 161.3
R29 VN.n18 VN.n17 161.3
R30 VN.n16 VN.n7 161.3
R31 VN.n15 VN.n14 161.3
R32 VN.n13 VN.n8 161.3
R33 VN.n12 VN.n11 161.3
R34 VN.n38 VN.n37 99.991
R35 VN.n77 VN.n76 99.991
R36 VN.n10 VN.t3 57.1567
R37 VN.n49 VN.t6 57.1567
R38 VN.n31 VN.n1 56.5193
R39 VN.n70 VN.n40 56.5193
R40 VN.n10 VN.n9 54.8849
R41 VN.n49 VN.n48 54.8849
R42 VN.n14 VN.n7 47.2923
R43 VN.n24 VN.n5 47.2923
R44 VN.n53 VN.n46 47.2923
R45 VN.n63 VN.n44 47.2923
R46 VN VN.n77 45.7936
R47 VN.n14 VN.n13 33.6945
R48 VN.n25 VN.n24 33.6945
R49 VN.n53 VN.n52 33.6945
R50 VN.n64 VN.n63 33.6945
R51 VN.n13 VN.n12 24.4675
R52 VN.n18 VN.n7 24.4675
R53 VN.n19 VN.n18 24.4675
R54 VN.n20 VN.n19 24.4675
R55 VN.n20 VN.n5 24.4675
R56 VN.n26 VN.n25 24.4675
R57 VN.n30 VN.n29 24.4675
R58 VN.n31 VN.n30 24.4675
R59 VN.n35 VN.n1 24.4675
R60 VN.n36 VN.n35 24.4675
R61 VN.n52 VN.n51 24.4675
R62 VN.n59 VN.n44 24.4675
R63 VN.n59 VN.n58 24.4675
R64 VN.n58 VN.n57 24.4675
R65 VN.n57 VN.n46 24.4675
R66 VN.n70 VN.n69 24.4675
R67 VN.n69 VN.n68 24.4675
R68 VN.n65 VN.n64 24.4675
R69 VN.n75 VN.n74 24.4675
R70 VN.n74 VN.n40 24.4675
R71 VN.n19 VN.t7 23.3384
R72 VN.n9 VN.t2 23.3384
R73 VN.n3 VN.t0 23.3384
R74 VN.n37 VN.t9 23.3384
R75 VN.n58 VN.t1 23.3384
R76 VN.n48 VN.t8 23.3384
R77 VN.n42 VN.t4 23.3384
R78 VN.n76 VN.t5 23.3384
R79 VN.n12 VN.n9 17.6167
R80 VN.n26 VN.n3 17.6167
R81 VN.n51 VN.n48 17.6167
R82 VN.n65 VN.n42 17.6167
R83 VN.n37 VN.n36 10.766
R84 VN.n76 VN.n75 10.766
R85 VN.n29 VN.n3 6.85126
R86 VN.n68 VN.n42 6.85126
R87 VN.n50 VN.n49 6.80183
R88 VN.n11 VN.n10 6.80183
R89 VN.n77 VN.n39 0.278367
R90 VN.n38 VN.n0 0.278367
R91 VN.n73 VN.n39 0.189894
R92 VN.n73 VN.n72 0.189894
R93 VN.n72 VN.n71 0.189894
R94 VN.n71 VN.n41 0.189894
R95 VN.n67 VN.n41 0.189894
R96 VN.n67 VN.n66 0.189894
R97 VN.n66 VN.n43 0.189894
R98 VN.n62 VN.n43 0.189894
R99 VN.n62 VN.n61 0.189894
R100 VN.n61 VN.n60 0.189894
R101 VN.n60 VN.n45 0.189894
R102 VN.n56 VN.n45 0.189894
R103 VN.n56 VN.n55 0.189894
R104 VN.n55 VN.n54 0.189894
R105 VN.n54 VN.n47 0.189894
R106 VN.n50 VN.n47 0.189894
R107 VN.n11 VN.n8 0.189894
R108 VN.n15 VN.n8 0.189894
R109 VN.n16 VN.n15 0.189894
R110 VN.n17 VN.n16 0.189894
R111 VN.n17 VN.n6 0.189894
R112 VN.n21 VN.n6 0.189894
R113 VN.n22 VN.n21 0.189894
R114 VN.n23 VN.n22 0.189894
R115 VN.n23 VN.n4 0.189894
R116 VN.n27 VN.n4 0.189894
R117 VN.n28 VN.n27 0.189894
R118 VN.n28 VN.n2 0.189894
R119 VN.n32 VN.n2 0.189894
R120 VN.n33 VN.n32 0.189894
R121 VN.n34 VN.n33 0.189894
R122 VN.n34 VN.n0 0.189894
R123 VN VN.n38 0.153454
R124 VDD2.n21 VDD2.n15 289.615
R125 VDD2.n6 VDD2.n0 289.615
R126 VDD2.n22 VDD2.n21 185
R127 VDD2.n20 VDD2.n19 185
R128 VDD2.n5 VDD2.n4 185
R129 VDD2.n7 VDD2.n6 185
R130 VDD2.n18 VDD2.t6 151.613
R131 VDD2.n3 VDD2.t2 151.613
R132 VDD2.n21 VDD2.n20 104.615
R133 VDD2.n6 VDD2.n5 104.615
R134 VDD2.n14 VDD2.n13 87.7227
R135 VDD2 VDD2.n29 87.7198
R136 VDD2.n28 VDD2.n27 85.929
R137 VDD2.n12 VDD2.n11 85.9289
R138 VDD2.n20 VDD2.t6 52.3082
R139 VDD2.n5 VDD2.t2 52.3082
R140 VDD2.n12 VDD2.n10 52.2994
R141 VDD2.n26 VDD2.n25 49.8338
R142 VDD2.n26 VDD2.n14 37.5386
R143 VDD2.n19 VDD2.n18 15.3979
R144 VDD2.n4 VDD2.n3 15.3979
R145 VDD2.n22 VDD2.n17 12.8005
R146 VDD2.n7 VDD2.n2 12.8005
R147 VDD2.n23 VDD2.n15 12.0247
R148 VDD2.n8 VDD2.n0 12.0247
R149 VDD2.n25 VDD2.n24 9.45567
R150 VDD2.n10 VDD2.n9 9.45567
R151 VDD2.n24 VDD2.n23 9.3005
R152 VDD2.n17 VDD2.n16 9.3005
R153 VDD2.n9 VDD2.n8 9.3005
R154 VDD2.n2 VDD2.n1 9.3005
R155 VDD2.n29 VDD2.t5 8.08213
R156 VDD2.n29 VDD2.t9 8.08213
R157 VDD2.n27 VDD2.t4 8.08213
R158 VDD2.n27 VDD2.t0 8.08213
R159 VDD2.n13 VDD2.t7 8.08213
R160 VDD2.n13 VDD2.t3 8.08213
R161 VDD2.n11 VDD2.t1 8.08213
R162 VDD2.n11 VDD2.t8 8.08213
R163 VDD2.n18 VDD2.n16 4.69785
R164 VDD2.n3 VDD2.n1 4.69785
R165 VDD2.n28 VDD2.n26 2.46602
R166 VDD2.n25 VDD2.n15 1.93989
R167 VDD2.n10 VDD2.n0 1.93989
R168 VDD2.n23 VDD2.n22 1.16414
R169 VDD2.n8 VDD2.n7 1.16414
R170 VDD2 VDD2.n28 0.675069
R171 VDD2.n14 VDD2.n12 0.561533
R172 VDD2.n19 VDD2.n17 0.388379
R173 VDD2.n4 VDD2.n2 0.388379
R174 VDD2.n24 VDD2.n16 0.155672
R175 VDD2.n9 VDD2.n1 0.155672
R176 VTAIL.n56 VTAIL.n50 289.615
R177 VTAIL.n8 VTAIL.n2 289.615
R178 VTAIL.n44 VTAIL.n38 289.615
R179 VTAIL.n28 VTAIL.n22 289.615
R180 VTAIL.n55 VTAIL.n54 185
R181 VTAIL.n57 VTAIL.n56 185
R182 VTAIL.n7 VTAIL.n6 185
R183 VTAIL.n9 VTAIL.n8 185
R184 VTAIL.n45 VTAIL.n44 185
R185 VTAIL.n43 VTAIL.n42 185
R186 VTAIL.n29 VTAIL.n28 185
R187 VTAIL.n27 VTAIL.n26 185
R188 VTAIL.n53 VTAIL.t10 151.613
R189 VTAIL.n5 VTAIL.t1 151.613
R190 VTAIL.n41 VTAIL.t5 151.613
R191 VTAIL.n25 VTAIL.t13 151.613
R192 VTAIL.n56 VTAIL.n55 104.615
R193 VTAIL.n8 VTAIL.n7 104.615
R194 VTAIL.n44 VTAIL.n43 104.615
R195 VTAIL.n28 VTAIL.n27 104.615
R196 VTAIL.n37 VTAIL.n36 69.2502
R197 VTAIL.n35 VTAIL.n34 69.2502
R198 VTAIL.n21 VTAIL.n20 69.2502
R199 VTAIL.n19 VTAIL.n18 69.2502
R200 VTAIL.n63 VTAIL.n62 69.2501
R201 VTAIL.n1 VTAIL.n0 69.2501
R202 VTAIL.n15 VTAIL.n14 69.2501
R203 VTAIL.n17 VTAIL.n16 69.2501
R204 VTAIL.n55 VTAIL.t10 52.3082
R205 VTAIL.n7 VTAIL.t1 52.3082
R206 VTAIL.n43 VTAIL.t5 52.3082
R207 VTAIL.n27 VTAIL.t13 52.3082
R208 VTAIL.n61 VTAIL.n60 33.155
R209 VTAIL.n13 VTAIL.n12 33.155
R210 VTAIL.n49 VTAIL.n48 33.155
R211 VTAIL.n33 VTAIL.n32 33.155
R212 VTAIL.n19 VTAIL.n17 19.41
R213 VTAIL.n61 VTAIL.n49 16.9445
R214 VTAIL.n54 VTAIL.n53 15.3979
R215 VTAIL.n6 VTAIL.n5 15.3979
R216 VTAIL.n42 VTAIL.n41 15.3979
R217 VTAIL.n26 VTAIL.n25 15.3979
R218 VTAIL.n57 VTAIL.n52 12.8005
R219 VTAIL.n9 VTAIL.n4 12.8005
R220 VTAIL.n45 VTAIL.n40 12.8005
R221 VTAIL.n29 VTAIL.n24 12.8005
R222 VTAIL.n58 VTAIL.n50 12.0247
R223 VTAIL.n10 VTAIL.n2 12.0247
R224 VTAIL.n46 VTAIL.n38 12.0247
R225 VTAIL.n30 VTAIL.n22 12.0247
R226 VTAIL.n60 VTAIL.n59 9.45567
R227 VTAIL.n12 VTAIL.n11 9.45567
R228 VTAIL.n48 VTAIL.n47 9.45567
R229 VTAIL.n32 VTAIL.n31 9.45567
R230 VTAIL.n59 VTAIL.n58 9.3005
R231 VTAIL.n52 VTAIL.n51 9.3005
R232 VTAIL.n11 VTAIL.n10 9.3005
R233 VTAIL.n4 VTAIL.n3 9.3005
R234 VTAIL.n47 VTAIL.n46 9.3005
R235 VTAIL.n40 VTAIL.n39 9.3005
R236 VTAIL.n31 VTAIL.n30 9.3005
R237 VTAIL.n24 VTAIL.n23 9.3005
R238 VTAIL.n62 VTAIL.t12 8.08213
R239 VTAIL.n62 VTAIL.t19 8.08213
R240 VTAIL.n0 VTAIL.t16 8.08213
R241 VTAIL.n0 VTAIL.t17 8.08213
R242 VTAIL.n14 VTAIL.t4 8.08213
R243 VTAIL.n14 VTAIL.t0 8.08213
R244 VTAIL.n16 VTAIL.t2 8.08213
R245 VTAIL.n16 VTAIL.t3 8.08213
R246 VTAIL.n36 VTAIL.t7 8.08213
R247 VTAIL.n36 VTAIL.t6 8.08213
R248 VTAIL.n34 VTAIL.t9 8.08213
R249 VTAIL.n34 VTAIL.t8 8.08213
R250 VTAIL.n20 VTAIL.t18 8.08213
R251 VTAIL.n20 VTAIL.t11 8.08213
R252 VTAIL.n18 VTAIL.t14 8.08213
R253 VTAIL.n18 VTAIL.t15 8.08213
R254 VTAIL.n53 VTAIL.n51 4.69785
R255 VTAIL.n5 VTAIL.n3 4.69785
R256 VTAIL.n41 VTAIL.n39 4.69785
R257 VTAIL.n25 VTAIL.n23 4.69785
R258 VTAIL.n21 VTAIL.n19 2.46602
R259 VTAIL.n33 VTAIL.n21 2.46602
R260 VTAIL.n37 VTAIL.n35 2.46602
R261 VTAIL.n49 VTAIL.n37 2.46602
R262 VTAIL.n17 VTAIL.n15 2.46602
R263 VTAIL.n15 VTAIL.n13 2.46602
R264 VTAIL.n63 VTAIL.n61 2.46602
R265 VTAIL.n60 VTAIL.n50 1.93989
R266 VTAIL.n12 VTAIL.n2 1.93989
R267 VTAIL.n48 VTAIL.n38 1.93989
R268 VTAIL.n32 VTAIL.n22 1.93989
R269 VTAIL VTAIL.n1 1.90783
R270 VTAIL.n35 VTAIL.n33 1.70309
R271 VTAIL.n13 VTAIL.n1 1.70309
R272 VTAIL.n58 VTAIL.n57 1.16414
R273 VTAIL.n10 VTAIL.n9 1.16414
R274 VTAIL.n46 VTAIL.n45 1.16414
R275 VTAIL.n30 VTAIL.n29 1.16414
R276 VTAIL VTAIL.n63 0.55869
R277 VTAIL.n54 VTAIL.n52 0.388379
R278 VTAIL.n6 VTAIL.n4 0.388379
R279 VTAIL.n42 VTAIL.n40 0.388379
R280 VTAIL.n26 VTAIL.n24 0.388379
R281 VTAIL.n59 VTAIL.n51 0.155672
R282 VTAIL.n11 VTAIL.n3 0.155672
R283 VTAIL.n47 VTAIL.n39 0.155672
R284 VTAIL.n31 VTAIL.n23 0.155672
R285 B.n593 B.n592 585
R286 B.n593 B.n107 585
R287 B.n596 B.n595 585
R288 B.n597 B.n130 585
R289 B.n599 B.n598 585
R290 B.n601 B.n129 585
R291 B.n604 B.n603 585
R292 B.n605 B.n128 585
R293 B.n607 B.n606 585
R294 B.n609 B.n127 585
R295 B.n612 B.n611 585
R296 B.n613 B.n126 585
R297 B.n615 B.n614 585
R298 B.n617 B.n125 585
R299 B.n620 B.n619 585
R300 B.n622 B.n122 585
R301 B.n624 B.n623 585
R302 B.n626 B.n121 585
R303 B.n629 B.n628 585
R304 B.n630 B.n120 585
R305 B.n632 B.n631 585
R306 B.n634 B.n119 585
R307 B.n636 B.n635 585
R308 B.n638 B.n637 585
R309 B.n641 B.n640 585
R310 B.n642 B.n114 585
R311 B.n644 B.n643 585
R312 B.n646 B.n113 585
R313 B.n649 B.n648 585
R314 B.n650 B.n112 585
R315 B.n652 B.n651 585
R316 B.n654 B.n111 585
R317 B.n657 B.n656 585
R318 B.n658 B.n110 585
R319 B.n660 B.n659 585
R320 B.n662 B.n109 585
R321 B.n665 B.n664 585
R322 B.n666 B.n108 585
R323 B.n591 B.n106 585
R324 B.n669 B.n106 585
R325 B.n590 B.n105 585
R326 B.n670 B.n105 585
R327 B.n589 B.n104 585
R328 B.n671 B.n104 585
R329 B.n588 B.n587 585
R330 B.n587 B.n100 585
R331 B.n586 B.n99 585
R332 B.n677 B.n99 585
R333 B.n585 B.n98 585
R334 B.n678 B.n98 585
R335 B.n584 B.n97 585
R336 B.n679 B.n97 585
R337 B.n583 B.n582 585
R338 B.n582 B.n96 585
R339 B.n581 B.n92 585
R340 B.n685 B.n92 585
R341 B.n580 B.n91 585
R342 B.n686 B.n91 585
R343 B.n579 B.n90 585
R344 B.n687 B.n90 585
R345 B.n578 B.n577 585
R346 B.n577 B.n86 585
R347 B.n576 B.n85 585
R348 B.n693 B.n85 585
R349 B.n575 B.n84 585
R350 B.n694 B.n84 585
R351 B.n574 B.n83 585
R352 B.n695 B.n83 585
R353 B.n573 B.n572 585
R354 B.n572 B.n79 585
R355 B.n571 B.n78 585
R356 B.n701 B.n78 585
R357 B.n570 B.n77 585
R358 B.n702 B.n77 585
R359 B.n569 B.n76 585
R360 B.n703 B.n76 585
R361 B.n568 B.n567 585
R362 B.n567 B.n75 585
R363 B.n566 B.n71 585
R364 B.n709 B.n71 585
R365 B.n565 B.n70 585
R366 B.n710 B.n70 585
R367 B.n564 B.n69 585
R368 B.n711 B.n69 585
R369 B.n563 B.n562 585
R370 B.n562 B.n65 585
R371 B.n561 B.n64 585
R372 B.n717 B.n64 585
R373 B.n560 B.n63 585
R374 B.n718 B.n63 585
R375 B.n559 B.n62 585
R376 B.n719 B.n62 585
R377 B.n558 B.n557 585
R378 B.n557 B.n61 585
R379 B.n556 B.n57 585
R380 B.n725 B.n57 585
R381 B.n555 B.n56 585
R382 B.n726 B.n56 585
R383 B.n554 B.n55 585
R384 B.n727 B.n55 585
R385 B.n553 B.n552 585
R386 B.n552 B.n51 585
R387 B.n551 B.n50 585
R388 B.n733 B.n50 585
R389 B.n550 B.n49 585
R390 B.n734 B.n49 585
R391 B.n549 B.n48 585
R392 B.n735 B.n48 585
R393 B.n548 B.n547 585
R394 B.n547 B.n47 585
R395 B.n546 B.n43 585
R396 B.n741 B.n43 585
R397 B.n545 B.n42 585
R398 B.n742 B.n42 585
R399 B.n544 B.n41 585
R400 B.n743 B.n41 585
R401 B.n543 B.n542 585
R402 B.n542 B.n37 585
R403 B.n541 B.n36 585
R404 B.n749 B.n36 585
R405 B.n540 B.n35 585
R406 B.n750 B.n35 585
R407 B.n539 B.n34 585
R408 B.n751 B.n34 585
R409 B.n538 B.n537 585
R410 B.n537 B.n30 585
R411 B.n536 B.n29 585
R412 B.n757 B.n29 585
R413 B.n535 B.n28 585
R414 B.n758 B.n28 585
R415 B.n534 B.n27 585
R416 B.n759 B.n27 585
R417 B.n533 B.n532 585
R418 B.n532 B.n23 585
R419 B.n531 B.n22 585
R420 B.n765 B.n22 585
R421 B.n530 B.n21 585
R422 B.n766 B.n21 585
R423 B.n529 B.n20 585
R424 B.n767 B.n20 585
R425 B.n528 B.n527 585
R426 B.n527 B.n16 585
R427 B.n526 B.n15 585
R428 B.n773 B.n15 585
R429 B.n525 B.n14 585
R430 B.n774 B.n14 585
R431 B.n524 B.n13 585
R432 B.n775 B.n13 585
R433 B.n523 B.n522 585
R434 B.n522 B.n12 585
R435 B.n521 B.n520 585
R436 B.n521 B.n8 585
R437 B.n519 B.n7 585
R438 B.n782 B.n7 585
R439 B.n518 B.n6 585
R440 B.n783 B.n6 585
R441 B.n517 B.n5 585
R442 B.n784 B.n5 585
R443 B.n516 B.n515 585
R444 B.n515 B.n4 585
R445 B.n514 B.n131 585
R446 B.n514 B.n513 585
R447 B.n504 B.n132 585
R448 B.n133 B.n132 585
R449 B.n506 B.n505 585
R450 B.n507 B.n506 585
R451 B.n503 B.n138 585
R452 B.n138 B.n137 585
R453 B.n502 B.n501 585
R454 B.n501 B.n500 585
R455 B.n140 B.n139 585
R456 B.n141 B.n140 585
R457 B.n493 B.n492 585
R458 B.n494 B.n493 585
R459 B.n491 B.n146 585
R460 B.n146 B.n145 585
R461 B.n490 B.n489 585
R462 B.n489 B.n488 585
R463 B.n148 B.n147 585
R464 B.n149 B.n148 585
R465 B.n481 B.n480 585
R466 B.n482 B.n481 585
R467 B.n479 B.n154 585
R468 B.n154 B.n153 585
R469 B.n478 B.n477 585
R470 B.n477 B.n476 585
R471 B.n156 B.n155 585
R472 B.n157 B.n156 585
R473 B.n469 B.n468 585
R474 B.n470 B.n469 585
R475 B.n467 B.n162 585
R476 B.n162 B.n161 585
R477 B.n466 B.n465 585
R478 B.n465 B.n464 585
R479 B.n164 B.n163 585
R480 B.n165 B.n164 585
R481 B.n457 B.n456 585
R482 B.n458 B.n457 585
R483 B.n455 B.n170 585
R484 B.n170 B.n169 585
R485 B.n454 B.n453 585
R486 B.n453 B.n452 585
R487 B.n172 B.n171 585
R488 B.n445 B.n172 585
R489 B.n444 B.n443 585
R490 B.n446 B.n444 585
R491 B.n442 B.n177 585
R492 B.n177 B.n176 585
R493 B.n441 B.n440 585
R494 B.n440 B.n439 585
R495 B.n179 B.n178 585
R496 B.n180 B.n179 585
R497 B.n432 B.n431 585
R498 B.n433 B.n432 585
R499 B.n430 B.n185 585
R500 B.n185 B.n184 585
R501 B.n429 B.n428 585
R502 B.n428 B.n427 585
R503 B.n187 B.n186 585
R504 B.n420 B.n187 585
R505 B.n419 B.n418 585
R506 B.n421 B.n419 585
R507 B.n417 B.n192 585
R508 B.n192 B.n191 585
R509 B.n416 B.n415 585
R510 B.n415 B.n414 585
R511 B.n194 B.n193 585
R512 B.n195 B.n194 585
R513 B.n407 B.n406 585
R514 B.n408 B.n407 585
R515 B.n405 B.n200 585
R516 B.n200 B.n199 585
R517 B.n404 B.n403 585
R518 B.n403 B.n402 585
R519 B.n202 B.n201 585
R520 B.n395 B.n202 585
R521 B.n394 B.n393 585
R522 B.n396 B.n394 585
R523 B.n392 B.n207 585
R524 B.n207 B.n206 585
R525 B.n391 B.n390 585
R526 B.n390 B.n389 585
R527 B.n209 B.n208 585
R528 B.n210 B.n209 585
R529 B.n382 B.n381 585
R530 B.n383 B.n382 585
R531 B.n380 B.n215 585
R532 B.n215 B.n214 585
R533 B.n379 B.n378 585
R534 B.n378 B.n377 585
R535 B.n217 B.n216 585
R536 B.n218 B.n217 585
R537 B.n370 B.n369 585
R538 B.n371 B.n370 585
R539 B.n368 B.n223 585
R540 B.n223 B.n222 585
R541 B.n367 B.n366 585
R542 B.n366 B.n365 585
R543 B.n225 B.n224 585
R544 B.n358 B.n225 585
R545 B.n357 B.n356 585
R546 B.n359 B.n357 585
R547 B.n355 B.n230 585
R548 B.n230 B.n229 585
R549 B.n354 B.n353 585
R550 B.n353 B.n352 585
R551 B.n232 B.n231 585
R552 B.n233 B.n232 585
R553 B.n345 B.n344 585
R554 B.n346 B.n345 585
R555 B.n343 B.n238 585
R556 B.n238 B.n237 585
R557 B.n342 B.n341 585
R558 B.n341 B.n340 585
R559 B.n337 B.n242 585
R560 B.n336 B.n335 585
R561 B.n333 B.n243 585
R562 B.n333 B.n241 585
R563 B.n332 B.n331 585
R564 B.n330 B.n329 585
R565 B.n328 B.n245 585
R566 B.n326 B.n325 585
R567 B.n324 B.n246 585
R568 B.n323 B.n322 585
R569 B.n320 B.n247 585
R570 B.n318 B.n317 585
R571 B.n316 B.n248 585
R572 B.n315 B.n314 585
R573 B.n312 B.n249 585
R574 B.n310 B.n309 585
R575 B.n308 B.n250 585
R576 B.n307 B.n306 585
R577 B.n304 B.n254 585
R578 B.n302 B.n301 585
R579 B.n300 B.n255 585
R580 B.n299 B.n298 585
R581 B.n296 B.n256 585
R582 B.n294 B.n293 585
R583 B.n291 B.n257 585
R584 B.n290 B.n289 585
R585 B.n287 B.n260 585
R586 B.n285 B.n284 585
R587 B.n283 B.n261 585
R588 B.n282 B.n281 585
R589 B.n279 B.n262 585
R590 B.n277 B.n276 585
R591 B.n275 B.n263 585
R592 B.n274 B.n273 585
R593 B.n271 B.n264 585
R594 B.n269 B.n268 585
R595 B.n267 B.n266 585
R596 B.n240 B.n239 585
R597 B.n339 B.n338 585
R598 B.n340 B.n339 585
R599 B.n236 B.n235 585
R600 B.n237 B.n236 585
R601 B.n348 B.n347 585
R602 B.n347 B.n346 585
R603 B.n349 B.n234 585
R604 B.n234 B.n233 585
R605 B.n351 B.n350 585
R606 B.n352 B.n351 585
R607 B.n228 B.n227 585
R608 B.n229 B.n228 585
R609 B.n361 B.n360 585
R610 B.n360 B.n359 585
R611 B.n362 B.n226 585
R612 B.n358 B.n226 585
R613 B.n364 B.n363 585
R614 B.n365 B.n364 585
R615 B.n221 B.n220 585
R616 B.n222 B.n221 585
R617 B.n373 B.n372 585
R618 B.n372 B.n371 585
R619 B.n374 B.n219 585
R620 B.n219 B.n218 585
R621 B.n376 B.n375 585
R622 B.n377 B.n376 585
R623 B.n213 B.n212 585
R624 B.n214 B.n213 585
R625 B.n385 B.n384 585
R626 B.n384 B.n383 585
R627 B.n386 B.n211 585
R628 B.n211 B.n210 585
R629 B.n388 B.n387 585
R630 B.n389 B.n388 585
R631 B.n205 B.n204 585
R632 B.n206 B.n205 585
R633 B.n398 B.n397 585
R634 B.n397 B.n396 585
R635 B.n399 B.n203 585
R636 B.n395 B.n203 585
R637 B.n401 B.n400 585
R638 B.n402 B.n401 585
R639 B.n198 B.n197 585
R640 B.n199 B.n198 585
R641 B.n410 B.n409 585
R642 B.n409 B.n408 585
R643 B.n411 B.n196 585
R644 B.n196 B.n195 585
R645 B.n413 B.n412 585
R646 B.n414 B.n413 585
R647 B.n190 B.n189 585
R648 B.n191 B.n190 585
R649 B.n423 B.n422 585
R650 B.n422 B.n421 585
R651 B.n424 B.n188 585
R652 B.n420 B.n188 585
R653 B.n426 B.n425 585
R654 B.n427 B.n426 585
R655 B.n183 B.n182 585
R656 B.n184 B.n183 585
R657 B.n435 B.n434 585
R658 B.n434 B.n433 585
R659 B.n436 B.n181 585
R660 B.n181 B.n180 585
R661 B.n438 B.n437 585
R662 B.n439 B.n438 585
R663 B.n175 B.n174 585
R664 B.n176 B.n175 585
R665 B.n448 B.n447 585
R666 B.n447 B.n446 585
R667 B.n449 B.n173 585
R668 B.n445 B.n173 585
R669 B.n451 B.n450 585
R670 B.n452 B.n451 585
R671 B.n168 B.n167 585
R672 B.n169 B.n168 585
R673 B.n460 B.n459 585
R674 B.n459 B.n458 585
R675 B.n461 B.n166 585
R676 B.n166 B.n165 585
R677 B.n463 B.n462 585
R678 B.n464 B.n463 585
R679 B.n160 B.n159 585
R680 B.n161 B.n160 585
R681 B.n472 B.n471 585
R682 B.n471 B.n470 585
R683 B.n473 B.n158 585
R684 B.n158 B.n157 585
R685 B.n475 B.n474 585
R686 B.n476 B.n475 585
R687 B.n152 B.n151 585
R688 B.n153 B.n152 585
R689 B.n484 B.n483 585
R690 B.n483 B.n482 585
R691 B.n485 B.n150 585
R692 B.n150 B.n149 585
R693 B.n487 B.n486 585
R694 B.n488 B.n487 585
R695 B.n144 B.n143 585
R696 B.n145 B.n144 585
R697 B.n496 B.n495 585
R698 B.n495 B.n494 585
R699 B.n497 B.n142 585
R700 B.n142 B.n141 585
R701 B.n499 B.n498 585
R702 B.n500 B.n499 585
R703 B.n136 B.n135 585
R704 B.n137 B.n136 585
R705 B.n509 B.n508 585
R706 B.n508 B.n507 585
R707 B.n510 B.n134 585
R708 B.n134 B.n133 585
R709 B.n512 B.n511 585
R710 B.n513 B.n512 585
R711 B.n3 B.n0 585
R712 B.n4 B.n3 585
R713 B.n781 B.n1 585
R714 B.n782 B.n781 585
R715 B.n780 B.n779 585
R716 B.n780 B.n8 585
R717 B.n778 B.n9 585
R718 B.n12 B.n9 585
R719 B.n777 B.n776 585
R720 B.n776 B.n775 585
R721 B.n11 B.n10 585
R722 B.n774 B.n11 585
R723 B.n772 B.n771 585
R724 B.n773 B.n772 585
R725 B.n770 B.n17 585
R726 B.n17 B.n16 585
R727 B.n769 B.n768 585
R728 B.n768 B.n767 585
R729 B.n19 B.n18 585
R730 B.n766 B.n19 585
R731 B.n764 B.n763 585
R732 B.n765 B.n764 585
R733 B.n762 B.n24 585
R734 B.n24 B.n23 585
R735 B.n761 B.n760 585
R736 B.n760 B.n759 585
R737 B.n26 B.n25 585
R738 B.n758 B.n26 585
R739 B.n756 B.n755 585
R740 B.n757 B.n756 585
R741 B.n754 B.n31 585
R742 B.n31 B.n30 585
R743 B.n753 B.n752 585
R744 B.n752 B.n751 585
R745 B.n33 B.n32 585
R746 B.n750 B.n33 585
R747 B.n748 B.n747 585
R748 B.n749 B.n748 585
R749 B.n746 B.n38 585
R750 B.n38 B.n37 585
R751 B.n745 B.n744 585
R752 B.n744 B.n743 585
R753 B.n40 B.n39 585
R754 B.n742 B.n40 585
R755 B.n740 B.n739 585
R756 B.n741 B.n740 585
R757 B.n738 B.n44 585
R758 B.n47 B.n44 585
R759 B.n737 B.n736 585
R760 B.n736 B.n735 585
R761 B.n46 B.n45 585
R762 B.n734 B.n46 585
R763 B.n732 B.n731 585
R764 B.n733 B.n732 585
R765 B.n730 B.n52 585
R766 B.n52 B.n51 585
R767 B.n729 B.n728 585
R768 B.n728 B.n727 585
R769 B.n54 B.n53 585
R770 B.n726 B.n54 585
R771 B.n724 B.n723 585
R772 B.n725 B.n724 585
R773 B.n722 B.n58 585
R774 B.n61 B.n58 585
R775 B.n721 B.n720 585
R776 B.n720 B.n719 585
R777 B.n60 B.n59 585
R778 B.n718 B.n60 585
R779 B.n716 B.n715 585
R780 B.n717 B.n716 585
R781 B.n714 B.n66 585
R782 B.n66 B.n65 585
R783 B.n713 B.n712 585
R784 B.n712 B.n711 585
R785 B.n68 B.n67 585
R786 B.n710 B.n68 585
R787 B.n708 B.n707 585
R788 B.n709 B.n708 585
R789 B.n706 B.n72 585
R790 B.n75 B.n72 585
R791 B.n705 B.n704 585
R792 B.n704 B.n703 585
R793 B.n74 B.n73 585
R794 B.n702 B.n74 585
R795 B.n700 B.n699 585
R796 B.n701 B.n700 585
R797 B.n698 B.n80 585
R798 B.n80 B.n79 585
R799 B.n697 B.n696 585
R800 B.n696 B.n695 585
R801 B.n82 B.n81 585
R802 B.n694 B.n82 585
R803 B.n692 B.n691 585
R804 B.n693 B.n692 585
R805 B.n690 B.n87 585
R806 B.n87 B.n86 585
R807 B.n689 B.n688 585
R808 B.n688 B.n687 585
R809 B.n89 B.n88 585
R810 B.n686 B.n89 585
R811 B.n684 B.n683 585
R812 B.n685 B.n684 585
R813 B.n682 B.n93 585
R814 B.n96 B.n93 585
R815 B.n681 B.n680 585
R816 B.n680 B.n679 585
R817 B.n95 B.n94 585
R818 B.n678 B.n95 585
R819 B.n676 B.n675 585
R820 B.n677 B.n676 585
R821 B.n674 B.n101 585
R822 B.n101 B.n100 585
R823 B.n673 B.n672 585
R824 B.n672 B.n671 585
R825 B.n103 B.n102 585
R826 B.n670 B.n103 585
R827 B.n668 B.n667 585
R828 B.n669 B.n668 585
R829 B.n785 B.n784 585
R830 B.n783 B.n2 585
R831 B.n668 B.n108 482.89
R832 B.n593 B.n106 482.89
R833 B.n341 B.n240 482.89
R834 B.n339 B.n242 482.89
R835 B.n594 B.n107 256.663
R836 B.n600 B.n107 256.663
R837 B.n602 B.n107 256.663
R838 B.n608 B.n107 256.663
R839 B.n610 B.n107 256.663
R840 B.n616 B.n107 256.663
R841 B.n618 B.n107 256.663
R842 B.n625 B.n107 256.663
R843 B.n627 B.n107 256.663
R844 B.n633 B.n107 256.663
R845 B.n118 B.n107 256.663
R846 B.n639 B.n107 256.663
R847 B.n645 B.n107 256.663
R848 B.n647 B.n107 256.663
R849 B.n653 B.n107 256.663
R850 B.n655 B.n107 256.663
R851 B.n661 B.n107 256.663
R852 B.n663 B.n107 256.663
R853 B.n334 B.n241 256.663
R854 B.n244 B.n241 256.663
R855 B.n327 B.n241 256.663
R856 B.n321 B.n241 256.663
R857 B.n319 B.n241 256.663
R858 B.n313 B.n241 256.663
R859 B.n311 B.n241 256.663
R860 B.n305 B.n241 256.663
R861 B.n303 B.n241 256.663
R862 B.n297 B.n241 256.663
R863 B.n295 B.n241 256.663
R864 B.n288 B.n241 256.663
R865 B.n286 B.n241 256.663
R866 B.n280 B.n241 256.663
R867 B.n278 B.n241 256.663
R868 B.n272 B.n241 256.663
R869 B.n270 B.n241 256.663
R870 B.n265 B.n241 256.663
R871 B.n787 B.n786 256.663
R872 B.n115 B.t14 231.276
R873 B.n123 B.t10 231.276
R874 B.n258 B.t17 231.276
R875 B.n251 B.t21 231.276
R876 B.n340 B.n241 183.69
R877 B.n669 B.n107 183.69
R878 B.n123 B.t12 177.196
R879 B.n258 B.t20 177.196
R880 B.n115 B.t15 177.196
R881 B.n251 B.t23 177.196
R882 B.n664 B.n662 163.367
R883 B.n660 B.n110 163.367
R884 B.n656 B.n654 163.367
R885 B.n652 B.n112 163.367
R886 B.n648 B.n646 163.367
R887 B.n644 B.n114 163.367
R888 B.n640 B.n638 163.367
R889 B.n635 B.n634 163.367
R890 B.n632 B.n120 163.367
R891 B.n628 B.n626 163.367
R892 B.n624 B.n122 163.367
R893 B.n619 B.n617 163.367
R894 B.n615 B.n126 163.367
R895 B.n611 B.n609 163.367
R896 B.n607 B.n128 163.367
R897 B.n603 B.n601 163.367
R898 B.n599 B.n130 163.367
R899 B.n595 B.n593 163.367
R900 B.n341 B.n238 163.367
R901 B.n345 B.n238 163.367
R902 B.n345 B.n232 163.367
R903 B.n353 B.n232 163.367
R904 B.n353 B.n230 163.367
R905 B.n357 B.n230 163.367
R906 B.n357 B.n225 163.367
R907 B.n366 B.n225 163.367
R908 B.n366 B.n223 163.367
R909 B.n370 B.n223 163.367
R910 B.n370 B.n217 163.367
R911 B.n378 B.n217 163.367
R912 B.n378 B.n215 163.367
R913 B.n382 B.n215 163.367
R914 B.n382 B.n209 163.367
R915 B.n390 B.n209 163.367
R916 B.n390 B.n207 163.367
R917 B.n394 B.n207 163.367
R918 B.n394 B.n202 163.367
R919 B.n403 B.n202 163.367
R920 B.n403 B.n200 163.367
R921 B.n407 B.n200 163.367
R922 B.n407 B.n194 163.367
R923 B.n415 B.n194 163.367
R924 B.n415 B.n192 163.367
R925 B.n419 B.n192 163.367
R926 B.n419 B.n187 163.367
R927 B.n428 B.n187 163.367
R928 B.n428 B.n185 163.367
R929 B.n432 B.n185 163.367
R930 B.n432 B.n179 163.367
R931 B.n440 B.n179 163.367
R932 B.n440 B.n177 163.367
R933 B.n444 B.n177 163.367
R934 B.n444 B.n172 163.367
R935 B.n453 B.n172 163.367
R936 B.n453 B.n170 163.367
R937 B.n457 B.n170 163.367
R938 B.n457 B.n164 163.367
R939 B.n465 B.n164 163.367
R940 B.n465 B.n162 163.367
R941 B.n469 B.n162 163.367
R942 B.n469 B.n156 163.367
R943 B.n477 B.n156 163.367
R944 B.n477 B.n154 163.367
R945 B.n481 B.n154 163.367
R946 B.n481 B.n148 163.367
R947 B.n489 B.n148 163.367
R948 B.n489 B.n146 163.367
R949 B.n493 B.n146 163.367
R950 B.n493 B.n140 163.367
R951 B.n501 B.n140 163.367
R952 B.n501 B.n138 163.367
R953 B.n506 B.n138 163.367
R954 B.n506 B.n132 163.367
R955 B.n514 B.n132 163.367
R956 B.n515 B.n514 163.367
R957 B.n515 B.n5 163.367
R958 B.n6 B.n5 163.367
R959 B.n7 B.n6 163.367
R960 B.n521 B.n7 163.367
R961 B.n522 B.n521 163.367
R962 B.n522 B.n13 163.367
R963 B.n14 B.n13 163.367
R964 B.n15 B.n14 163.367
R965 B.n527 B.n15 163.367
R966 B.n527 B.n20 163.367
R967 B.n21 B.n20 163.367
R968 B.n22 B.n21 163.367
R969 B.n532 B.n22 163.367
R970 B.n532 B.n27 163.367
R971 B.n28 B.n27 163.367
R972 B.n29 B.n28 163.367
R973 B.n537 B.n29 163.367
R974 B.n537 B.n34 163.367
R975 B.n35 B.n34 163.367
R976 B.n36 B.n35 163.367
R977 B.n542 B.n36 163.367
R978 B.n542 B.n41 163.367
R979 B.n42 B.n41 163.367
R980 B.n43 B.n42 163.367
R981 B.n547 B.n43 163.367
R982 B.n547 B.n48 163.367
R983 B.n49 B.n48 163.367
R984 B.n50 B.n49 163.367
R985 B.n552 B.n50 163.367
R986 B.n552 B.n55 163.367
R987 B.n56 B.n55 163.367
R988 B.n57 B.n56 163.367
R989 B.n557 B.n57 163.367
R990 B.n557 B.n62 163.367
R991 B.n63 B.n62 163.367
R992 B.n64 B.n63 163.367
R993 B.n562 B.n64 163.367
R994 B.n562 B.n69 163.367
R995 B.n70 B.n69 163.367
R996 B.n71 B.n70 163.367
R997 B.n567 B.n71 163.367
R998 B.n567 B.n76 163.367
R999 B.n77 B.n76 163.367
R1000 B.n78 B.n77 163.367
R1001 B.n572 B.n78 163.367
R1002 B.n572 B.n83 163.367
R1003 B.n84 B.n83 163.367
R1004 B.n85 B.n84 163.367
R1005 B.n577 B.n85 163.367
R1006 B.n577 B.n90 163.367
R1007 B.n91 B.n90 163.367
R1008 B.n92 B.n91 163.367
R1009 B.n582 B.n92 163.367
R1010 B.n582 B.n97 163.367
R1011 B.n98 B.n97 163.367
R1012 B.n99 B.n98 163.367
R1013 B.n587 B.n99 163.367
R1014 B.n587 B.n104 163.367
R1015 B.n105 B.n104 163.367
R1016 B.n106 B.n105 163.367
R1017 B.n335 B.n333 163.367
R1018 B.n333 B.n332 163.367
R1019 B.n329 B.n328 163.367
R1020 B.n326 B.n246 163.367
R1021 B.n322 B.n320 163.367
R1022 B.n318 B.n248 163.367
R1023 B.n314 B.n312 163.367
R1024 B.n310 B.n250 163.367
R1025 B.n306 B.n304 163.367
R1026 B.n302 B.n255 163.367
R1027 B.n298 B.n296 163.367
R1028 B.n294 B.n257 163.367
R1029 B.n289 B.n287 163.367
R1030 B.n285 B.n261 163.367
R1031 B.n281 B.n279 163.367
R1032 B.n277 B.n263 163.367
R1033 B.n273 B.n271 163.367
R1034 B.n269 B.n266 163.367
R1035 B.n339 B.n236 163.367
R1036 B.n347 B.n236 163.367
R1037 B.n347 B.n234 163.367
R1038 B.n351 B.n234 163.367
R1039 B.n351 B.n228 163.367
R1040 B.n360 B.n228 163.367
R1041 B.n360 B.n226 163.367
R1042 B.n364 B.n226 163.367
R1043 B.n364 B.n221 163.367
R1044 B.n372 B.n221 163.367
R1045 B.n372 B.n219 163.367
R1046 B.n376 B.n219 163.367
R1047 B.n376 B.n213 163.367
R1048 B.n384 B.n213 163.367
R1049 B.n384 B.n211 163.367
R1050 B.n388 B.n211 163.367
R1051 B.n388 B.n205 163.367
R1052 B.n397 B.n205 163.367
R1053 B.n397 B.n203 163.367
R1054 B.n401 B.n203 163.367
R1055 B.n401 B.n198 163.367
R1056 B.n409 B.n198 163.367
R1057 B.n409 B.n196 163.367
R1058 B.n413 B.n196 163.367
R1059 B.n413 B.n190 163.367
R1060 B.n422 B.n190 163.367
R1061 B.n422 B.n188 163.367
R1062 B.n426 B.n188 163.367
R1063 B.n426 B.n183 163.367
R1064 B.n434 B.n183 163.367
R1065 B.n434 B.n181 163.367
R1066 B.n438 B.n181 163.367
R1067 B.n438 B.n175 163.367
R1068 B.n447 B.n175 163.367
R1069 B.n447 B.n173 163.367
R1070 B.n451 B.n173 163.367
R1071 B.n451 B.n168 163.367
R1072 B.n459 B.n168 163.367
R1073 B.n459 B.n166 163.367
R1074 B.n463 B.n166 163.367
R1075 B.n463 B.n160 163.367
R1076 B.n471 B.n160 163.367
R1077 B.n471 B.n158 163.367
R1078 B.n475 B.n158 163.367
R1079 B.n475 B.n152 163.367
R1080 B.n483 B.n152 163.367
R1081 B.n483 B.n150 163.367
R1082 B.n487 B.n150 163.367
R1083 B.n487 B.n144 163.367
R1084 B.n495 B.n144 163.367
R1085 B.n495 B.n142 163.367
R1086 B.n499 B.n142 163.367
R1087 B.n499 B.n136 163.367
R1088 B.n508 B.n136 163.367
R1089 B.n508 B.n134 163.367
R1090 B.n512 B.n134 163.367
R1091 B.n512 B.n3 163.367
R1092 B.n785 B.n3 163.367
R1093 B.n781 B.n2 163.367
R1094 B.n781 B.n780 163.367
R1095 B.n780 B.n9 163.367
R1096 B.n776 B.n9 163.367
R1097 B.n776 B.n11 163.367
R1098 B.n772 B.n11 163.367
R1099 B.n772 B.n17 163.367
R1100 B.n768 B.n17 163.367
R1101 B.n768 B.n19 163.367
R1102 B.n764 B.n19 163.367
R1103 B.n764 B.n24 163.367
R1104 B.n760 B.n24 163.367
R1105 B.n760 B.n26 163.367
R1106 B.n756 B.n26 163.367
R1107 B.n756 B.n31 163.367
R1108 B.n752 B.n31 163.367
R1109 B.n752 B.n33 163.367
R1110 B.n748 B.n33 163.367
R1111 B.n748 B.n38 163.367
R1112 B.n744 B.n38 163.367
R1113 B.n744 B.n40 163.367
R1114 B.n740 B.n40 163.367
R1115 B.n740 B.n44 163.367
R1116 B.n736 B.n44 163.367
R1117 B.n736 B.n46 163.367
R1118 B.n732 B.n46 163.367
R1119 B.n732 B.n52 163.367
R1120 B.n728 B.n52 163.367
R1121 B.n728 B.n54 163.367
R1122 B.n724 B.n54 163.367
R1123 B.n724 B.n58 163.367
R1124 B.n720 B.n58 163.367
R1125 B.n720 B.n60 163.367
R1126 B.n716 B.n60 163.367
R1127 B.n716 B.n66 163.367
R1128 B.n712 B.n66 163.367
R1129 B.n712 B.n68 163.367
R1130 B.n708 B.n68 163.367
R1131 B.n708 B.n72 163.367
R1132 B.n704 B.n72 163.367
R1133 B.n704 B.n74 163.367
R1134 B.n700 B.n74 163.367
R1135 B.n700 B.n80 163.367
R1136 B.n696 B.n80 163.367
R1137 B.n696 B.n82 163.367
R1138 B.n692 B.n82 163.367
R1139 B.n692 B.n87 163.367
R1140 B.n688 B.n87 163.367
R1141 B.n688 B.n89 163.367
R1142 B.n684 B.n89 163.367
R1143 B.n684 B.n93 163.367
R1144 B.n680 B.n93 163.367
R1145 B.n680 B.n95 163.367
R1146 B.n676 B.n95 163.367
R1147 B.n676 B.n101 163.367
R1148 B.n672 B.n101 163.367
R1149 B.n672 B.n103 163.367
R1150 B.n668 B.n103 163.367
R1151 B.n124 B.t13 121.73
R1152 B.n259 B.t19 121.73
R1153 B.n116 B.t16 121.73
R1154 B.n252 B.t22 121.73
R1155 B.n340 B.n237 96.829
R1156 B.n346 B.n237 96.829
R1157 B.n346 B.n233 96.829
R1158 B.n352 B.n233 96.829
R1159 B.n352 B.n229 96.829
R1160 B.n359 B.n229 96.829
R1161 B.n359 B.n358 96.829
R1162 B.n365 B.n222 96.829
R1163 B.n371 B.n222 96.829
R1164 B.n371 B.n218 96.829
R1165 B.n377 B.n218 96.829
R1166 B.n377 B.n214 96.829
R1167 B.n383 B.n214 96.829
R1168 B.n383 B.n210 96.829
R1169 B.n389 B.n210 96.829
R1170 B.n389 B.n206 96.829
R1171 B.n396 B.n206 96.829
R1172 B.n396 B.n395 96.829
R1173 B.n402 B.n199 96.829
R1174 B.n408 B.n199 96.829
R1175 B.n408 B.n195 96.829
R1176 B.n414 B.n195 96.829
R1177 B.n414 B.n191 96.829
R1178 B.n421 B.n191 96.829
R1179 B.n421 B.n420 96.829
R1180 B.n427 B.n184 96.829
R1181 B.n433 B.n184 96.829
R1182 B.n433 B.n180 96.829
R1183 B.n439 B.n180 96.829
R1184 B.n439 B.n176 96.829
R1185 B.n446 B.n176 96.829
R1186 B.n446 B.n445 96.829
R1187 B.n452 B.n169 96.829
R1188 B.n458 B.n169 96.829
R1189 B.n458 B.n165 96.829
R1190 B.n464 B.n165 96.829
R1191 B.n464 B.n161 96.829
R1192 B.n470 B.n161 96.829
R1193 B.n470 B.n157 96.829
R1194 B.n476 B.n157 96.829
R1195 B.n482 B.n153 96.829
R1196 B.n482 B.n149 96.829
R1197 B.n488 B.n149 96.829
R1198 B.n488 B.n145 96.829
R1199 B.n494 B.n145 96.829
R1200 B.n494 B.n141 96.829
R1201 B.n500 B.n141 96.829
R1202 B.n507 B.n137 96.829
R1203 B.n507 B.n133 96.829
R1204 B.n513 B.n133 96.829
R1205 B.n513 B.n4 96.829
R1206 B.n784 B.n4 96.829
R1207 B.n784 B.n783 96.829
R1208 B.n783 B.n782 96.829
R1209 B.n782 B.n8 96.829
R1210 B.n12 B.n8 96.829
R1211 B.n775 B.n12 96.829
R1212 B.n775 B.n774 96.829
R1213 B.n773 B.n16 96.829
R1214 B.n767 B.n16 96.829
R1215 B.n767 B.n766 96.829
R1216 B.n766 B.n765 96.829
R1217 B.n765 B.n23 96.829
R1218 B.n759 B.n23 96.829
R1219 B.n759 B.n758 96.829
R1220 B.n757 B.n30 96.829
R1221 B.n751 B.n30 96.829
R1222 B.n751 B.n750 96.829
R1223 B.n750 B.n749 96.829
R1224 B.n749 B.n37 96.829
R1225 B.n743 B.n37 96.829
R1226 B.n743 B.n742 96.829
R1227 B.n742 B.n741 96.829
R1228 B.n735 B.n47 96.829
R1229 B.n735 B.n734 96.829
R1230 B.n734 B.n733 96.829
R1231 B.n733 B.n51 96.829
R1232 B.n727 B.n51 96.829
R1233 B.n727 B.n726 96.829
R1234 B.n726 B.n725 96.829
R1235 B.n719 B.n61 96.829
R1236 B.n719 B.n718 96.829
R1237 B.n718 B.n717 96.829
R1238 B.n717 B.n65 96.829
R1239 B.n711 B.n65 96.829
R1240 B.n711 B.n710 96.829
R1241 B.n710 B.n709 96.829
R1242 B.n703 B.n75 96.829
R1243 B.n703 B.n702 96.829
R1244 B.n702 B.n701 96.829
R1245 B.n701 B.n79 96.829
R1246 B.n695 B.n79 96.829
R1247 B.n695 B.n694 96.829
R1248 B.n694 B.n693 96.829
R1249 B.n693 B.n86 96.829
R1250 B.n687 B.n86 96.829
R1251 B.n687 B.n686 96.829
R1252 B.n686 B.n685 96.829
R1253 B.n679 B.n96 96.829
R1254 B.n679 B.n678 96.829
R1255 B.n678 B.n677 96.829
R1256 B.n677 B.n100 96.829
R1257 B.n671 B.n100 96.829
R1258 B.n671 B.n670 96.829
R1259 B.n670 B.n669 96.829
R1260 B.n402 B.t2 92.5571
R1261 B.n709 B.t5 92.5571
R1262 B.n445 B.t4 84.0134
R1263 B.n47 B.t7 84.0134
R1264 B.n663 B.n108 71.676
R1265 B.n662 B.n661 71.676
R1266 B.n655 B.n110 71.676
R1267 B.n654 B.n653 71.676
R1268 B.n647 B.n112 71.676
R1269 B.n646 B.n645 71.676
R1270 B.n639 B.n114 71.676
R1271 B.n638 B.n118 71.676
R1272 B.n634 B.n633 71.676
R1273 B.n627 B.n120 71.676
R1274 B.n626 B.n625 71.676
R1275 B.n618 B.n122 71.676
R1276 B.n617 B.n616 71.676
R1277 B.n610 B.n126 71.676
R1278 B.n609 B.n608 71.676
R1279 B.n602 B.n128 71.676
R1280 B.n601 B.n600 71.676
R1281 B.n594 B.n130 71.676
R1282 B.n595 B.n594 71.676
R1283 B.n600 B.n599 71.676
R1284 B.n603 B.n602 71.676
R1285 B.n608 B.n607 71.676
R1286 B.n611 B.n610 71.676
R1287 B.n616 B.n615 71.676
R1288 B.n619 B.n618 71.676
R1289 B.n625 B.n624 71.676
R1290 B.n628 B.n627 71.676
R1291 B.n633 B.n632 71.676
R1292 B.n635 B.n118 71.676
R1293 B.n640 B.n639 71.676
R1294 B.n645 B.n644 71.676
R1295 B.n648 B.n647 71.676
R1296 B.n653 B.n652 71.676
R1297 B.n656 B.n655 71.676
R1298 B.n661 B.n660 71.676
R1299 B.n664 B.n663 71.676
R1300 B.n334 B.n242 71.676
R1301 B.n332 B.n244 71.676
R1302 B.n328 B.n327 71.676
R1303 B.n321 B.n246 71.676
R1304 B.n320 B.n319 71.676
R1305 B.n313 B.n248 71.676
R1306 B.n312 B.n311 71.676
R1307 B.n305 B.n250 71.676
R1308 B.n304 B.n303 71.676
R1309 B.n297 B.n255 71.676
R1310 B.n296 B.n295 71.676
R1311 B.n288 B.n257 71.676
R1312 B.n287 B.n286 71.676
R1313 B.n280 B.n261 71.676
R1314 B.n279 B.n278 71.676
R1315 B.n272 B.n263 71.676
R1316 B.n271 B.n270 71.676
R1317 B.n266 B.n265 71.676
R1318 B.n335 B.n334 71.676
R1319 B.n329 B.n244 71.676
R1320 B.n327 B.n326 71.676
R1321 B.n322 B.n321 71.676
R1322 B.n319 B.n318 71.676
R1323 B.n314 B.n313 71.676
R1324 B.n311 B.n310 71.676
R1325 B.n306 B.n305 71.676
R1326 B.n303 B.n302 71.676
R1327 B.n298 B.n297 71.676
R1328 B.n295 B.n294 71.676
R1329 B.n289 B.n288 71.676
R1330 B.n286 B.n285 71.676
R1331 B.n281 B.n280 71.676
R1332 B.n278 B.n277 71.676
R1333 B.n273 B.n272 71.676
R1334 B.n270 B.n269 71.676
R1335 B.n265 B.n240 71.676
R1336 B.n786 B.n785 71.676
R1337 B.n786 B.n2 71.676
R1338 B.t0 B.n153 69.774
R1339 B.n758 B.t8 69.774
R1340 B.n500 B.t1 66.9261
R1341 B.t9 B.n773 66.9261
R1342 B.n117 B.n116 59.5399
R1343 B.n621 B.n124 59.5399
R1344 B.n292 B.n259 59.5399
R1345 B.n253 B.n252 59.5399
R1346 B.n365 B.t18 55.5345
R1347 B.n685 B.t11 55.5345
R1348 B.n116 B.n115 55.4672
R1349 B.n124 B.n123 55.4672
R1350 B.n259 B.n258 55.4672
R1351 B.n252 B.n251 55.4672
R1352 B.n427 B.t3 52.6866
R1353 B.n725 B.t6 52.6866
R1354 B.n420 B.t3 44.1429
R1355 B.n61 B.t6 44.1429
R1356 B.n358 B.t18 41.295
R1357 B.n96 B.t11 41.295
R1358 B.n338 B.n337 31.3761
R1359 B.n342 B.n239 31.3761
R1360 B.n592 B.n591 31.3761
R1361 B.n667 B.n666 31.3761
R1362 B.t1 B.n137 29.9034
R1363 B.n774 B.t9 29.9034
R1364 B.n476 B.t0 27.0555
R1365 B.t8 B.n757 27.0555
R1366 B B.n787 18.0485
R1367 B.n452 B.t4 12.816
R1368 B.n741 B.t7 12.816
R1369 B.n338 B.n235 10.6151
R1370 B.n348 B.n235 10.6151
R1371 B.n349 B.n348 10.6151
R1372 B.n350 B.n349 10.6151
R1373 B.n350 B.n227 10.6151
R1374 B.n361 B.n227 10.6151
R1375 B.n362 B.n361 10.6151
R1376 B.n363 B.n362 10.6151
R1377 B.n363 B.n220 10.6151
R1378 B.n373 B.n220 10.6151
R1379 B.n374 B.n373 10.6151
R1380 B.n375 B.n374 10.6151
R1381 B.n375 B.n212 10.6151
R1382 B.n385 B.n212 10.6151
R1383 B.n386 B.n385 10.6151
R1384 B.n387 B.n386 10.6151
R1385 B.n387 B.n204 10.6151
R1386 B.n398 B.n204 10.6151
R1387 B.n399 B.n398 10.6151
R1388 B.n400 B.n399 10.6151
R1389 B.n400 B.n197 10.6151
R1390 B.n410 B.n197 10.6151
R1391 B.n411 B.n410 10.6151
R1392 B.n412 B.n411 10.6151
R1393 B.n412 B.n189 10.6151
R1394 B.n423 B.n189 10.6151
R1395 B.n424 B.n423 10.6151
R1396 B.n425 B.n424 10.6151
R1397 B.n425 B.n182 10.6151
R1398 B.n435 B.n182 10.6151
R1399 B.n436 B.n435 10.6151
R1400 B.n437 B.n436 10.6151
R1401 B.n437 B.n174 10.6151
R1402 B.n448 B.n174 10.6151
R1403 B.n449 B.n448 10.6151
R1404 B.n450 B.n449 10.6151
R1405 B.n450 B.n167 10.6151
R1406 B.n460 B.n167 10.6151
R1407 B.n461 B.n460 10.6151
R1408 B.n462 B.n461 10.6151
R1409 B.n462 B.n159 10.6151
R1410 B.n472 B.n159 10.6151
R1411 B.n473 B.n472 10.6151
R1412 B.n474 B.n473 10.6151
R1413 B.n474 B.n151 10.6151
R1414 B.n484 B.n151 10.6151
R1415 B.n485 B.n484 10.6151
R1416 B.n486 B.n485 10.6151
R1417 B.n486 B.n143 10.6151
R1418 B.n496 B.n143 10.6151
R1419 B.n497 B.n496 10.6151
R1420 B.n498 B.n497 10.6151
R1421 B.n498 B.n135 10.6151
R1422 B.n509 B.n135 10.6151
R1423 B.n510 B.n509 10.6151
R1424 B.n511 B.n510 10.6151
R1425 B.n511 B.n0 10.6151
R1426 B.n337 B.n336 10.6151
R1427 B.n336 B.n243 10.6151
R1428 B.n331 B.n243 10.6151
R1429 B.n331 B.n330 10.6151
R1430 B.n330 B.n245 10.6151
R1431 B.n325 B.n245 10.6151
R1432 B.n325 B.n324 10.6151
R1433 B.n324 B.n323 10.6151
R1434 B.n323 B.n247 10.6151
R1435 B.n317 B.n247 10.6151
R1436 B.n317 B.n316 10.6151
R1437 B.n316 B.n315 10.6151
R1438 B.n315 B.n249 10.6151
R1439 B.n309 B.n308 10.6151
R1440 B.n308 B.n307 10.6151
R1441 B.n307 B.n254 10.6151
R1442 B.n301 B.n254 10.6151
R1443 B.n301 B.n300 10.6151
R1444 B.n300 B.n299 10.6151
R1445 B.n299 B.n256 10.6151
R1446 B.n293 B.n256 10.6151
R1447 B.n291 B.n290 10.6151
R1448 B.n290 B.n260 10.6151
R1449 B.n284 B.n260 10.6151
R1450 B.n284 B.n283 10.6151
R1451 B.n283 B.n282 10.6151
R1452 B.n282 B.n262 10.6151
R1453 B.n276 B.n262 10.6151
R1454 B.n276 B.n275 10.6151
R1455 B.n275 B.n274 10.6151
R1456 B.n274 B.n264 10.6151
R1457 B.n268 B.n264 10.6151
R1458 B.n268 B.n267 10.6151
R1459 B.n267 B.n239 10.6151
R1460 B.n343 B.n342 10.6151
R1461 B.n344 B.n343 10.6151
R1462 B.n344 B.n231 10.6151
R1463 B.n354 B.n231 10.6151
R1464 B.n355 B.n354 10.6151
R1465 B.n356 B.n355 10.6151
R1466 B.n356 B.n224 10.6151
R1467 B.n367 B.n224 10.6151
R1468 B.n368 B.n367 10.6151
R1469 B.n369 B.n368 10.6151
R1470 B.n369 B.n216 10.6151
R1471 B.n379 B.n216 10.6151
R1472 B.n380 B.n379 10.6151
R1473 B.n381 B.n380 10.6151
R1474 B.n381 B.n208 10.6151
R1475 B.n391 B.n208 10.6151
R1476 B.n392 B.n391 10.6151
R1477 B.n393 B.n392 10.6151
R1478 B.n393 B.n201 10.6151
R1479 B.n404 B.n201 10.6151
R1480 B.n405 B.n404 10.6151
R1481 B.n406 B.n405 10.6151
R1482 B.n406 B.n193 10.6151
R1483 B.n416 B.n193 10.6151
R1484 B.n417 B.n416 10.6151
R1485 B.n418 B.n417 10.6151
R1486 B.n418 B.n186 10.6151
R1487 B.n429 B.n186 10.6151
R1488 B.n430 B.n429 10.6151
R1489 B.n431 B.n430 10.6151
R1490 B.n431 B.n178 10.6151
R1491 B.n441 B.n178 10.6151
R1492 B.n442 B.n441 10.6151
R1493 B.n443 B.n442 10.6151
R1494 B.n443 B.n171 10.6151
R1495 B.n454 B.n171 10.6151
R1496 B.n455 B.n454 10.6151
R1497 B.n456 B.n455 10.6151
R1498 B.n456 B.n163 10.6151
R1499 B.n466 B.n163 10.6151
R1500 B.n467 B.n466 10.6151
R1501 B.n468 B.n467 10.6151
R1502 B.n468 B.n155 10.6151
R1503 B.n478 B.n155 10.6151
R1504 B.n479 B.n478 10.6151
R1505 B.n480 B.n479 10.6151
R1506 B.n480 B.n147 10.6151
R1507 B.n490 B.n147 10.6151
R1508 B.n491 B.n490 10.6151
R1509 B.n492 B.n491 10.6151
R1510 B.n492 B.n139 10.6151
R1511 B.n502 B.n139 10.6151
R1512 B.n503 B.n502 10.6151
R1513 B.n505 B.n503 10.6151
R1514 B.n505 B.n504 10.6151
R1515 B.n504 B.n131 10.6151
R1516 B.n516 B.n131 10.6151
R1517 B.n517 B.n516 10.6151
R1518 B.n518 B.n517 10.6151
R1519 B.n519 B.n518 10.6151
R1520 B.n520 B.n519 10.6151
R1521 B.n523 B.n520 10.6151
R1522 B.n524 B.n523 10.6151
R1523 B.n525 B.n524 10.6151
R1524 B.n526 B.n525 10.6151
R1525 B.n528 B.n526 10.6151
R1526 B.n529 B.n528 10.6151
R1527 B.n530 B.n529 10.6151
R1528 B.n531 B.n530 10.6151
R1529 B.n533 B.n531 10.6151
R1530 B.n534 B.n533 10.6151
R1531 B.n535 B.n534 10.6151
R1532 B.n536 B.n535 10.6151
R1533 B.n538 B.n536 10.6151
R1534 B.n539 B.n538 10.6151
R1535 B.n540 B.n539 10.6151
R1536 B.n541 B.n540 10.6151
R1537 B.n543 B.n541 10.6151
R1538 B.n544 B.n543 10.6151
R1539 B.n545 B.n544 10.6151
R1540 B.n546 B.n545 10.6151
R1541 B.n548 B.n546 10.6151
R1542 B.n549 B.n548 10.6151
R1543 B.n550 B.n549 10.6151
R1544 B.n551 B.n550 10.6151
R1545 B.n553 B.n551 10.6151
R1546 B.n554 B.n553 10.6151
R1547 B.n555 B.n554 10.6151
R1548 B.n556 B.n555 10.6151
R1549 B.n558 B.n556 10.6151
R1550 B.n559 B.n558 10.6151
R1551 B.n560 B.n559 10.6151
R1552 B.n561 B.n560 10.6151
R1553 B.n563 B.n561 10.6151
R1554 B.n564 B.n563 10.6151
R1555 B.n565 B.n564 10.6151
R1556 B.n566 B.n565 10.6151
R1557 B.n568 B.n566 10.6151
R1558 B.n569 B.n568 10.6151
R1559 B.n570 B.n569 10.6151
R1560 B.n571 B.n570 10.6151
R1561 B.n573 B.n571 10.6151
R1562 B.n574 B.n573 10.6151
R1563 B.n575 B.n574 10.6151
R1564 B.n576 B.n575 10.6151
R1565 B.n578 B.n576 10.6151
R1566 B.n579 B.n578 10.6151
R1567 B.n580 B.n579 10.6151
R1568 B.n581 B.n580 10.6151
R1569 B.n583 B.n581 10.6151
R1570 B.n584 B.n583 10.6151
R1571 B.n585 B.n584 10.6151
R1572 B.n586 B.n585 10.6151
R1573 B.n588 B.n586 10.6151
R1574 B.n589 B.n588 10.6151
R1575 B.n590 B.n589 10.6151
R1576 B.n591 B.n590 10.6151
R1577 B.n779 B.n1 10.6151
R1578 B.n779 B.n778 10.6151
R1579 B.n778 B.n777 10.6151
R1580 B.n777 B.n10 10.6151
R1581 B.n771 B.n10 10.6151
R1582 B.n771 B.n770 10.6151
R1583 B.n770 B.n769 10.6151
R1584 B.n769 B.n18 10.6151
R1585 B.n763 B.n18 10.6151
R1586 B.n763 B.n762 10.6151
R1587 B.n762 B.n761 10.6151
R1588 B.n761 B.n25 10.6151
R1589 B.n755 B.n25 10.6151
R1590 B.n755 B.n754 10.6151
R1591 B.n754 B.n753 10.6151
R1592 B.n753 B.n32 10.6151
R1593 B.n747 B.n32 10.6151
R1594 B.n747 B.n746 10.6151
R1595 B.n746 B.n745 10.6151
R1596 B.n745 B.n39 10.6151
R1597 B.n739 B.n39 10.6151
R1598 B.n739 B.n738 10.6151
R1599 B.n738 B.n737 10.6151
R1600 B.n737 B.n45 10.6151
R1601 B.n731 B.n45 10.6151
R1602 B.n731 B.n730 10.6151
R1603 B.n730 B.n729 10.6151
R1604 B.n729 B.n53 10.6151
R1605 B.n723 B.n53 10.6151
R1606 B.n723 B.n722 10.6151
R1607 B.n722 B.n721 10.6151
R1608 B.n721 B.n59 10.6151
R1609 B.n715 B.n59 10.6151
R1610 B.n715 B.n714 10.6151
R1611 B.n714 B.n713 10.6151
R1612 B.n713 B.n67 10.6151
R1613 B.n707 B.n67 10.6151
R1614 B.n707 B.n706 10.6151
R1615 B.n706 B.n705 10.6151
R1616 B.n705 B.n73 10.6151
R1617 B.n699 B.n73 10.6151
R1618 B.n699 B.n698 10.6151
R1619 B.n698 B.n697 10.6151
R1620 B.n697 B.n81 10.6151
R1621 B.n691 B.n81 10.6151
R1622 B.n691 B.n690 10.6151
R1623 B.n690 B.n689 10.6151
R1624 B.n689 B.n88 10.6151
R1625 B.n683 B.n88 10.6151
R1626 B.n683 B.n682 10.6151
R1627 B.n682 B.n681 10.6151
R1628 B.n681 B.n94 10.6151
R1629 B.n675 B.n94 10.6151
R1630 B.n675 B.n674 10.6151
R1631 B.n674 B.n673 10.6151
R1632 B.n673 B.n102 10.6151
R1633 B.n667 B.n102 10.6151
R1634 B.n666 B.n665 10.6151
R1635 B.n665 B.n109 10.6151
R1636 B.n659 B.n109 10.6151
R1637 B.n659 B.n658 10.6151
R1638 B.n658 B.n657 10.6151
R1639 B.n657 B.n111 10.6151
R1640 B.n651 B.n111 10.6151
R1641 B.n651 B.n650 10.6151
R1642 B.n650 B.n649 10.6151
R1643 B.n649 B.n113 10.6151
R1644 B.n643 B.n113 10.6151
R1645 B.n643 B.n642 10.6151
R1646 B.n642 B.n641 10.6151
R1647 B.n637 B.n636 10.6151
R1648 B.n636 B.n119 10.6151
R1649 B.n631 B.n119 10.6151
R1650 B.n631 B.n630 10.6151
R1651 B.n630 B.n629 10.6151
R1652 B.n629 B.n121 10.6151
R1653 B.n623 B.n121 10.6151
R1654 B.n623 B.n622 10.6151
R1655 B.n620 B.n125 10.6151
R1656 B.n614 B.n125 10.6151
R1657 B.n614 B.n613 10.6151
R1658 B.n613 B.n612 10.6151
R1659 B.n612 B.n127 10.6151
R1660 B.n606 B.n127 10.6151
R1661 B.n606 B.n605 10.6151
R1662 B.n605 B.n604 10.6151
R1663 B.n604 B.n129 10.6151
R1664 B.n598 B.n129 10.6151
R1665 B.n598 B.n597 10.6151
R1666 B.n597 B.n596 10.6151
R1667 B.n596 B.n592 10.6151
R1668 B.n787 B.n0 8.11757
R1669 B.n787 B.n1 8.11757
R1670 B.n309 B.n253 6.5566
R1671 B.n293 B.n292 6.5566
R1672 B.n637 B.n117 6.5566
R1673 B.n622 B.n621 6.5566
R1674 B.n395 B.t2 4.27234
R1675 B.n75 B.t5 4.27234
R1676 B.n253 B.n249 4.05904
R1677 B.n292 B.n291 4.05904
R1678 B.n641 B.n117 4.05904
R1679 B.n621 B.n620 4.05904
R1680 VP.n25 VP.n24 161.3
R1681 VP.n26 VP.n21 161.3
R1682 VP.n28 VP.n27 161.3
R1683 VP.n29 VP.n20 161.3
R1684 VP.n31 VP.n30 161.3
R1685 VP.n32 VP.n19 161.3
R1686 VP.n34 VP.n33 161.3
R1687 VP.n35 VP.n18 161.3
R1688 VP.n37 VP.n36 161.3
R1689 VP.n38 VP.n17 161.3
R1690 VP.n40 VP.n39 161.3
R1691 VP.n42 VP.n41 161.3
R1692 VP.n43 VP.n15 161.3
R1693 VP.n45 VP.n44 161.3
R1694 VP.n46 VP.n14 161.3
R1695 VP.n48 VP.n47 161.3
R1696 VP.n49 VP.n13 161.3
R1697 VP.n88 VP.n0 161.3
R1698 VP.n87 VP.n86 161.3
R1699 VP.n85 VP.n1 161.3
R1700 VP.n84 VP.n83 161.3
R1701 VP.n82 VP.n2 161.3
R1702 VP.n81 VP.n80 161.3
R1703 VP.n79 VP.n78 161.3
R1704 VP.n77 VP.n4 161.3
R1705 VP.n76 VP.n75 161.3
R1706 VP.n74 VP.n5 161.3
R1707 VP.n73 VP.n72 161.3
R1708 VP.n71 VP.n6 161.3
R1709 VP.n70 VP.n69 161.3
R1710 VP.n68 VP.n7 161.3
R1711 VP.n67 VP.n66 161.3
R1712 VP.n65 VP.n8 161.3
R1713 VP.n64 VP.n63 161.3
R1714 VP.n62 VP.n61 161.3
R1715 VP.n60 VP.n10 161.3
R1716 VP.n59 VP.n58 161.3
R1717 VP.n57 VP.n11 161.3
R1718 VP.n56 VP.n55 161.3
R1719 VP.n54 VP.n12 161.3
R1720 VP.n53 VP.n52 99.991
R1721 VP.n90 VP.n89 99.991
R1722 VP.n51 VP.n50 99.991
R1723 VP.n23 VP.t0 57.1567
R1724 VP.n59 VP.n11 56.5193
R1725 VP.n83 VP.n1 56.5193
R1726 VP.n44 VP.n14 56.5193
R1727 VP.n23 VP.n22 54.8849
R1728 VP.n66 VP.n7 47.2923
R1729 VP.n76 VP.n5 47.2923
R1730 VP.n37 VP.n18 47.2923
R1731 VP.n27 VP.n20 47.2923
R1732 VP.n52 VP.n51 45.5147
R1733 VP.n66 VP.n65 33.6945
R1734 VP.n77 VP.n76 33.6945
R1735 VP.n38 VP.n37 33.6945
R1736 VP.n27 VP.n26 33.6945
R1737 VP.n55 VP.n54 24.4675
R1738 VP.n55 VP.n11 24.4675
R1739 VP.n60 VP.n59 24.4675
R1740 VP.n61 VP.n60 24.4675
R1741 VP.n65 VP.n64 24.4675
R1742 VP.n70 VP.n7 24.4675
R1743 VP.n71 VP.n70 24.4675
R1744 VP.n72 VP.n71 24.4675
R1745 VP.n72 VP.n5 24.4675
R1746 VP.n78 VP.n77 24.4675
R1747 VP.n82 VP.n81 24.4675
R1748 VP.n83 VP.n82 24.4675
R1749 VP.n87 VP.n1 24.4675
R1750 VP.n88 VP.n87 24.4675
R1751 VP.n48 VP.n14 24.4675
R1752 VP.n49 VP.n48 24.4675
R1753 VP.n39 VP.n38 24.4675
R1754 VP.n43 VP.n42 24.4675
R1755 VP.n44 VP.n43 24.4675
R1756 VP.n31 VP.n20 24.4675
R1757 VP.n32 VP.n31 24.4675
R1758 VP.n33 VP.n32 24.4675
R1759 VP.n33 VP.n18 24.4675
R1760 VP.n26 VP.n25 24.4675
R1761 VP.n71 VP.t9 23.3384
R1762 VP.n53 VP.t4 23.3384
R1763 VP.n9 VP.t8 23.3384
R1764 VP.n3 VP.t6 23.3384
R1765 VP.n89 VP.t7 23.3384
R1766 VP.n32 VP.t2 23.3384
R1767 VP.n50 VP.t5 23.3384
R1768 VP.n16 VP.t3 23.3384
R1769 VP.n22 VP.t1 23.3384
R1770 VP.n64 VP.n9 17.6167
R1771 VP.n78 VP.n3 17.6167
R1772 VP.n39 VP.n16 17.6167
R1773 VP.n25 VP.n22 17.6167
R1774 VP.n54 VP.n53 10.766
R1775 VP.n89 VP.n88 10.766
R1776 VP.n50 VP.n49 10.766
R1777 VP.n61 VP.n9 6.85126
R1778 VP.n81 VP.n3 6.85126
R1779 VP.n42 VP.n16 6.85126
R1780 VP.n24 VP.n23 6.80183
R1781 VP.n51 VP.n13 0.278367
R1782 VP.n52 VP.n12 0.278367
R1783 VP.n90 VP.n0 0.278367
R1784 VP.n24 VP.n21 0.189894
R1785 VP.n28 VP.n21 0.189894
R1786 VP.n29 VP.n28 0.189894
R1787 VP.n30 VP.n29 0.189894
R1788 VP.n30 VP.n19 0.189894
R1789 VP.n34 VP.n19 0.189894
R1790 VP.n35 VP.n34 0.189894
R1791 VP.n36 VP.n35 0.189894
R1792 VP.n36 VP.n17 0.189894
R1793 VP.n40 VP.n17 0.189894
R1794 VP.n41 VP.n40 0.189894
R1795 VP.n41 VP.n15 0.189894
R1796 VP.n45 VP.n15 0.189894
R1797 VP.n46 VP.n45 0.189894
R1798 VP.n47 VP.n46 0.189894
R1799 VP.n47 VP.n13 0.189894
R1800 VP.n56 VP.n12 0.189894
R1801 VP.n57 VP.n56 0.189894
R1802 VP.n58 VP.n57 0.189894
R1803 VP.n58 VP.n10 0.189894
R1804 VP.n62 VP.n10 0.189894
R1805 VP.n63 VP.n62 0.189894
R1806 VP.n63 VP.n8 0.189894
R1807 VP.n67 VP.n8 0.189894
R1808 VP.n68 VP.n67 0.189894
R1809 VP.n69 VP.n68 0.189894
R1810 VP.n69 VP.n6 0.189894
R1811 VP.n73 VP.n6 0.189894
R1812 VP.n74 VP.n73 0.189894
R1813 VP.n75 VP.n74 0.189894
R1814 VP.n75 VP.n4 0.189894
R1815 VP.n79 VP.n4 0.189894
R1816 VP.n80 VP.n79 0.189894
R1817 VP.n80 VP.n2 0.189894
R1818 VP.n84 VP.n2 0.189894
R1819 VP.n85 VP.n84 0.189894
R1820 VP.n86 VP.n85 0.189894
R1821 VP.n86 VP.n0 0.189894
R1822 VP VP.n90 0.153454
R1823 VDD1.n6 VDD1.n0 289.615
R1824 VDD1.n19 VDD1.n13 289.615
R1825 VDD1.n7 VDD1.n6 185
R1826 VDD1.n5 VDD1.n4 185
R1827 VDD1.n18 VDD1.n17 185
R1828 VDD1.n20 VDD1.n19 185
R1829 VDD1.n3 VDD1.t9 151.613
R1830 VDD1.n16 VDD1.t5 151.613
R1831 VDD1.n6 VDD1.n5 104.615
R1832 VDD1.n19 VDD1.n18 104.615
R1833 VDD1.n27 VDD1.n26 87.7227
R1834 VDD1.n12 VDD1.n11 85.929
R1835 VDD1.n29 VDD1.n28 85.9289
R1836 VDD1.n25 VDD1.n24 85.9289
R1837 VDD1.n5 VDD1.t9 52.3082
R1838 VDD1.n18 VDD1.t5 52.3082
R1839 VDD1.n12 VDD1.n10 52.2994
R1840 VDD1.n25 VDD1.n23 52.2994
R1841 VDD1.n29 VDD1.n27 39.3543
R1842 VDD1.n4 VDD1.n3 15.3979
R1843 VDD1.n17 VDD1.n16 15.3979
R1844 VDD1.n7 VDD1.n2 12.8005
R1845 VDD1.n20 VDD1.n15 12.8005
R1846 VDD1.n8 VDD1.n0 12.0247
R1847 VDD1.n21 VDD1.n13 12.0247
R1848 VDD1.n10 VDD1.n9 9.45567
R1849 VDD1.n23 VDD1.n22 9.45567
R1850 VDD1.n9 VDD1.n8 9.3005
R1851 VDD1.n2 VDD1.n1 9.3005
R1852 VDD1.n22 VDD1.n21 9.3005
R1853 VDD1.n15 VDD1.n14 9.3005
R1854 VDD1.n28 VDD1.t6 8.08213
R1855 VDD1.n28 VDD1.t4 8.08213
R1856 VDD1.n11 VDD1.t8 8.08213
R1857 VDD1.n11 VDD1.t7 8.08213
R1858 VDD1.n26 VDD1.t3 8.08213
R1859 VDD1.n26 VDD1.t2 8.08213
R1860 VDD1.n24 VDD1.t1 8.08213
R1861 VDD1.n24 VDD1.t0 8.08213
R1862 VDD1.n3 VDD1.n1 4.69785
R1863 VDD1.n16 VDD1.n14 4.69785
R1864 VDD1.n10 VDD1.n0 1.93989
R1865 VDD1.n23 VDD1.n13 1.93989
R1866 VDD1 VDD1.n29 1.79145
R1867 VDD1.n8 VDD1.n7 1.16414
R1868 VDD1.n21 VDD1.n20 1.16414
R1869 VDD1 VDD1.n12 0.675069
R1870 VDD1.n27 VDD1.n25 0.561533
R1871 VDD1.n4 VDD1.n2 0.388379
R1872 VDD1.n17 VDD1.n15 0.388379
R1873 VDD1.n9 VDD1.n1 0.155672
R1874 VDD1.n22 VDD1.n14 0.155672
C0 VDD1 VTAIL 5.91498f
C1 VDD2 VTAIL 5.96766f
C2 VP VN 6.53328f
C3 VDD1 VP 2.99708f
C4 VDD1 VN 0.159009f
C5 VDD2 VP 0.580777f
C6 VDD2 VN 2.57883f
C7 VDD2 VDD1 2.12756f
C8 VP VTAIL 3.91967f
C9 VTAIL VN 3.90552f
C10 VDD2 B 5.549469f
C11 VDD1 B 5.431669f
C12 VTAIL B 3.877965f
C13 VN B 16.97071f
C14 VP B 15.414915f
C15 VDD1.n0 B 0.038472f
C16 VDD1.n1 B 0.216867f
C17 VDD1.n2 B 0.015849f
C18 VDD1.t9 B 0.06409f
C19 VDD1.n3 B 0.102556f
C20 VDD1.n4 B 0.021206f
C21 VDD1.n5 B 0.028096f
C22 VDD1.n6 B 0.07582f
C23 VDD1.n7 B 0.016781f
C24 VDD1.n8 B 0.015849f
C25 VDD1.n9 B 0.07019f
C26 VDD1.n10 B 0.076071f
C27 VDD1.t8 B 0.057104f
C28 VDD1.t7 B 0.057104f
C29 VDD1.n11 B 0.404301f
C30 VDD1.n12 B 0.791016f
C31 VDD1.n13 B 0.038472f
C32 VDD1.n14 B 0.216867f
C33 VDD1.n15 B 0.015849f
C34 VDD1.t5 B 0.06409f
C35 VDD1.n16 B 0.102556f
C36 VDD1.n17 B 0.021206f
C37 VDD1.n18 B 0.028096f
C38 VDD1.n19 B 0.07582f
C39 VDD1.n20 B 0.016781f
C40 VDD1.n21 B 0.015849f
C41 VDD1.n22 B 0.07019f
C42 VDD1.n23 B 0.076071f
C43 VDD1.t1 B 0.057104f
C44 VDD1.t0 B 0.057104f
C45 VDD1.n24 B 0.4043f
C46 VDD1.n25 B 0.781446f
C47 VDD1.t3 B 0.057104f
C48 VDD1.t2 B 0.057104f
C49 VDD1.n26 B 0.417206f
C50 VDD1.n27 B 2.81877f
C51 VDD1.t6 B 0.057104f
C52 VDD1.t4 B 0.057104f
C53 VDD1.n28 B 0.4043f
C54 VDD1.n29 B 2.80382f
C55 VP.n0 B 0.039052f
C56 VP.t7 B 0.444537f
C57 VP.n1 B 0.039939f
C58 VP.n2 B 0.029621f
C59 VP.t6 B 0.444537f
C60 VP.n3 B 0.198769f
C61 VP.n4 B 0.029621f
C62 VP.n5 B 0.055992f
C63 VP.n6 B 0.029621f
C64 VP.t9 B 0.444537f
C65 VP.n7 B 0.055992f
C66 VP.n8 B 0.029621f
C67 VP.t8 B 0.444537f
C68 VP.n9 B 0.198769f
C69 VP.n10 B 0.029621f
C70 VP.n11 B 0.039939f
C71 VP.n12 B 0.039052f
C72 VP.t4 B 0.444537f
C73 VP.n13 B 0.039052f
C74 VP.t5 B 0.444537f
C75 VP.n14 B 0.039939f
C76 VP.n15 B 0.029621f
C77 VP.t3 B 0.444537f
C78 VP.n16 B 0.198769f
C79 VP.n17 B 0.029621f
C80 VP.n18 B 0.055992f
C81 VP.n19 B 0.029621f
C82 VP.t2 B 0.444537f
C83 VP.n20 B 0.055992f
C84 VP.n21 B 0.029621f
C85 VP.t1 B 0.444537f
C86 VP.n22 B 0.289299f
C87 VP.t0 B 0.669107f
C88 VP.n23 B 0.271039f
C89 VP.n24 B 0.284254f
C90 VP.n25 B 0.047574f
C91 VP.n26 B 0.059831f
C92 VP.n27 B 0.025864f
C93 VP.n28 B 0.029621f
C94 VP.n29 B 0.029621f
C95 VP.n30 B 0.029621f
C96 VP.n31 B 0.055205f
C97 VP.n32 B 0.22672f
C98 VP.n33 B 0.055205f
C99 VP.n34 B 0.029621f
C100 VP.n35 B 0.029621f
C101 VP.n36 B 0.029621f
C102 VP.n37 B 0.025864f
C103 VP.n38 B 0.059831f
C104 VP.n39 B 0.047574f
C105 VP.n40 B 0.029621f
C106 VP.n41 B 0.029621f
C107 VP.n42 B 0.035582f
C108 VP.n43 B 0.055205f
C109 VP.n44 B 0.046542f
C110 VP.n45 B 0.029621f
C111 VP.n46 B 0.029621f
C112 VP.n47 B 0.029621f
C113 VP.n48 B 0.055205f
C114 VP.n49 B 0.039942f
C115 VP.n50 B 0.296624f
C116 VP.n51 B 1.42964f
C117 VP.n52 B 1.45303f
C118 VP.n53 B 0.296624f
C119 VP.n54 B 0.039942f
C120 VP.n55 B 0.055205f
C121 VP.n56 B 0.029621f
C122 VP.n57 B 0.029621f
C123 VP.n58 B 0.029621f
C124 VP.n59 B 0.046542f
C125 VP.n60 B 0.055205f
C126 VP.n61 B 0.035582f
C127 VP.n62 B 0.029621f
C128 VP.n63 B 0.029621f
C129 VP.n64 B 0.047574f
C130 VP.n65 B 0.059831f
C131 VP.n66 B 0.025864f
C132 VP.n67 B 0.029621f
C133 VP.n68 B 0.029621f
C134 VP.n69 B 0.029621f
C135 VP.n70 B 0.055205f
C136 VP.n71 B 0.22672f
C137 VP.n72 B 0.055205f
C138 VP.n73 B 0.029621f
C139 VP.n74 B 0.029621f
C140 VP.n75 B 0.029621f
C141 VP.n76 B 0.025864f
C142 VP.n77 B 0.059831f
C143 VP.n78 B 0.047574f
C144 VP.n79 B 0.029621f
C145 VP.n80 B 0.029621f
C146 VP.n81 B 0.035582f
C147 VP.n82 B 0.055205f
C148 VP.n83 B 0.046542f
C149 VP.n84 B 0.029621f
C150 VP.n85 B 0.029621f
C151 VP.n86 B 0.029621f
C152 VP.n87 B 0.055205f
C153 VP.n88 B 0.039942f
C154 VP.n89 B 0.296624f
C155 VP.n90 B 0.046961f
C156 VTAIL.t16 B 0.067426f
C157 VTAIL.t17 B 0.067426f
C158 VTAIL.n0 B 0.418092f
C159 VTAIL.n1 B 0.669854f
C160 VTAIL.n2 B 0.045427f
C161 VTAIL.n3 B 0.256069f
C162 VTAIL.n4 B 0.018714f
C163 VTAIL.t1 B 0.075675f
C164 VTAIL.n5 B 0.121094f
C165 VTAIL.n6 B 0.025039f
C166 VTAIL.n7 B 0.033175f
C167 VTAIL.n8 B 0.089525f
C168 VTAIL.n9 B 0.019815f
C169 VTAIL.n10 B 0.018714f
C170 VTAIL.n11 B 0.082878f
C171 VTAIL.n12 B 0.049524f
C172 VTAIL.n13 B 0.498824f
C173 VTAIL.t4 B 0.067426f
C174 VTAIL.t0 B 0.067426f
C175 VTAIL.n14 B 0.418092f
C176 VTAIL.n15 B 0.818108f
C177 VTAIL.t2 B 0.067426f
C178 VTAIL.t3 B 0.067426f
C179 VTAIL.n16 B 0.418092f
C180 VTAIL.n17 B 1.80487f
C181 VTAIL.t14 B 0.067426f
C182 VTAIL.t15 B 0.067426f
C183 VTAIL.n18 B 0.418095f
C184 VTAIL.n19 B 1.80487f
C185 VTAIL.t18 B 0.067426f
C186 VTAIL.t11 B 0.067426f
C187 VTAIL.n20 B 0.418095f
C188 VTAIL.n21 B 0.818105f
C189 VTAIL.n22 B 0.045427f
C190 VTAIL.n23 B 0.256069f
C191 VTAIL.n24 B 0.018714f
C192 VTAIL.t13 B 0.075675f
C193 VTAIL.n25 B 0.121094f
C194 VTAIL.n26 B 0.025039f
C195 VTAIL.n27 B 0.033175f
C196 VTAIL.n28 B 0.089525f
C197 VTAIL.n29 B 0.019815f
C198 VTAIL.n30 B 0.018714f
C199 VTAIL.n31 B 0.082878f
C200 VTAIL.n32 B 0.049524f
C201 VTAIL.n33 B 0.498824f
C202 VTAIL.t9 B 0.067426f
C203 VTAIL.t8 B 0.067426f
C204 VTAIL.n34 B 0.418095f
C205 VTAIL.n35 B 0.73249f
C206 VTAIL.t7 B 0.067426f
C207 VTAIL.t6 B 0.067426f
C208 VTAIL.n36 B 0.418095f
C209 VTAIL.n37 B 0.818105f
C210 VTAIL.n38 B 0.045427f
C211 VTAIL.n39 B 0.256069f
C212 VTAIL.n40 B 0.018714f
C213 VTAIL.t5 B 0.075675f
C214 VTAIL.n41 B 0.121094f
C215 VTAIL.n42 B 0.025039f
C216 VTAIL.n43 B 0.033175f
C217 VTAIL.n44 B 0.089525f
C218 VTAIL.n45 B 0.019815f
C219 VTAIL.n46 B 0.018714f
C220 VTAIL.n47 B 0.082878f
C221 VTAIL.n48 B 0.049524f
C222 VTAIL.n49 B 1.29452f
C223 VTAIL.n50 B 0.045427f
C224 VTAIL.n51 B 0.256069f
C225 VTAIL.n52 B 0.018714f
C226 VTAIL.t10 B 0.075675f
C227 VTAIL.n53 B 0.121094f
C228 VTAIL.n54 B 0.025039f
C229 VTAIL.n55 B 0.033175f
C230 VTAIL.n56 B 0.089525f
C231 VTAIL.n57 B 0.019815f
C232 VTAIL.n58 B 0.018714f
C233 VTAIL.n59 B 0.082878f
C234 VTAIL.n60 B 0.049524f
C235 VTAIL.n61 B 1.29452f
C236 VTAIL.t12 B 0.067426f
C237 VTAIL.t19 B 0.067426f
C238 VTAIL.n62 B 0.418092f
C239 VTAIL.n63 B 0.604071f
C240 VDD2.n0 B 0.037798f
C241 VDD2.n1 B 0.213063f
C242 VDD2.n2 B 0.015571f
C243 VDD2.t2 B 0.062965f
C244 VDD2.n3 B 0.100756f
C245 VDD2.n4 B 0.020834f
C246 VDD2.n5 B 0.027603f
C247 VDD2.n6 B 0.074489f
C248 VDD2.n7 B 0.016487f
C249 VDD2.n8 B 0.015571f
C250 VDD2.n9 B 0.068959f
C251 VDD2.n10 B 0.074736f
C252 VDD2.t1 B 0.056102f
C253 VDD2.t8 B 0.056102f
C254 VDD2.n11 B 0.397207f
C255 VDD2.n12 B 0.767737f
C256 VDD2.t7 B 0.056102f
C257 VDD2.t3 B 0.056102f
C258 VDD2.n13 B 0.409887f
C259 VDD2.n14 B 2.63648f
C260 VDD2.n15 B 0.037798f
C261 VDD2.n16 B 0.213063f
C262 VDD2.n17 B 0.015571f
C263 VDD2.t6 B 0.062965f
C264 VDD2.n18 B 0.100756f
C265 VDD2.n19 B 0.020834f
C266 VDD2.n20 B 0.027603f
C267 VDD2.n21 B 0.074489f
C268 VDD2.n22 B 0.016487f
C269 VDD2.n23 B 0.015571f
C270 VDD2.n24 B 0.068959f
C271 VDD2.n25 B 0.0612f
C272 VDD2.n26 B 2.44814f
C273 VDD2.t4 B 0.056102f
C274 VDD2.t0 B 0.056102f
C275 VDD2.n27 B 0.397209f
C276 VDD2.n28 B 0.503536f
C277 VDD2.t5 B 0.056102f
C278 VDD2.t9 B 0.056102f
C279 VDD2.n29 B 0.409854f
C280 VN.n0 B 0.037769f
C281 VN.t9 B 0.429931f
C282 VN.n1 B 0.038627f
C283 VN.n2 B 0.028647f
C284 VN.t0 B 0.429931f
C285 VN.n3 B 0.192239f
C286 VN.n4 B 0.028647f
C287 VN.n5 B 0.054153f
C288 VN.n6 B 0.028647f
C289 VN.t7 B 0.429931f
C290 VN.n7 B 0.054153f
C291 VN.n8 B 0.028647f
C292 VN.t2 B 0.429931f
C293 VN.n9 B 0.279794f
C294 VN.t3 B 0.647123f
C295 VN.n10 B 0.262134f
C296 VN.n11 B 0.274915f
C297 VN.n12 B 0.046011f
C298 VN.n13 B 0.057865f
C299 VN.n14 B 0.025014f
C300 VN.n15 B 0.028647f
C301 VN.n16 B 0.028647f
C302 VN.n17 B 0.028647f
C303 VN.n18 B 0.053392f
C304 VN.n19 B 0.21927f
C305 VN.n20 B 0.053392f
C306 VN.n21 B 0.028647f
C307 VN.n22 B 0.028647f
C308 VN.n23 B 0.028647f
C309 VN.n24 B 0.025014f
C310 VN.n25 B 0.057865f
C311 VN.n26 B 0.046011f
C312 VN.n27 B 0.028647f
C313 VN.n28 B 0.028647f
C314 VN.n29 B 0.034413f
C315 VN.n30 B 0.053392f
C316 VN.n31 B 0.045013f
C317 VN.n32 B 0.028647f
C318 VN.n33 B 0.028647f
C319 VN.n34 B 0.028647f
C320 VN.n35 B 0.053392f
C321 VN.n36 B 0.03863f
C322 VN.n37 B 0.286878f
C323 VN.n38 B 0.045418f
C324 VN.n39 B 0.037769f
C325 VN.t5 B 0.429931f
C326 VN.n40 B 0.038627f
C327 VN.n41 B 0.028647f
C328 VN.t4 B 0.429931f
C329 VN.n42 B 0.192239f
C330 VN.n43 B 0.028647f
C331 VN.n44 B 0.054153f
C332 VN.n45 B 0.028647f
C333 VN.t1 B 0.429931f
C334 VN.n46 B 0.054153f
C335 VN.n47 B 0.028647f
C336 VN.t8 B 0.429931f
C337 VN.n48 B 0.279794f
C338 VN.t6 B 0.647123f
C339 VN.n49 B 0.262134f
C340 VN.n50 B 0.274915f
C341 VN.n51 B 0.046011f
C342 VN.n52 B 0.057865f
C343 VN.n53 B 0.025014f
C344 VN.n54 B 0.028647f
C345 VN.n55 B 0.028647f
C346 VN.n56 B 0.028647f
C347 VN.n57 B 0.053392f
C348 VN.n58 B 0.21927f
C349 VN.n59 B 0.053392f
C350 VN.n60 B 0.028647f
C351 VN.n61 B 0.028647f
C352 VN.n62 B 0.028647f
C353 VN.n63 B 0.025014f
C354 VN.n64 B 0.057865f
C355 VN.n65 B 0.046011f
C356 VN.n66 B 0.028647f
C357 VN.n67 B 0.028647f
C358 VN.n68 B 0.034413f
C359 VN.n69 B 0.053392f
C360 VN.n70 B 0.045013f
C361 VN.n71 B 0.028647f
C362 VN.n72 B 0.028647f
C363 VN.n73 B 0.028647f
C364 VN.n74 B 0.053392f
C365 VN.n75 B 0.03863f
C366 VN.n76 B 0.286878f
C367 VN.n77 B 1.3983f
.ends

