* NGSPICE file created from diff_pair_sample_0741.ext - technology: sky130A

.subckt diff_pair_sample_0741 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1564_n4646# sky130_fd_pr__pfet_01v8 ad=7.1721 pd=37.56 as=0 ps=0 w=18.39 l=0.66
X1 VTAIL.t7 VP.t0 VDD1.t1 w_n1564_n4646# sky130_fd_pr__pfet_01v8 ad=7.1721 pd=37.56 as=3.03435 ps=18.72 w=18.39 l=0.66
X2 B.t8 B.t6 B.t7 w_n1564_n4646# sky130_fd_pr__pfet_01v8 ad=7.1721 pd=37.56 as=0 ps=0 w=18.39 l=0.66
X3 VDD2.t3 VN.t0 VTAIL.t1 w_n1564_n4646# sky130_fd_pr__pfet_01v8 ad=3.03435 pd=18.72 as=7.1721 ps=37.56 w=18.39 l=0.66
X4 VTAIL.t2 VN.t1 VDD2.t2 w_n1564_n4646# sky130_fd_pr__pfet_01v8 ad=7.1721 pd=37.56 as=3.03435 ps=18.72 w=18.39 l=0.66
X5 B.t5 B.t3 B.t4 w_n1564_n4646# sky130_fd_pr__pfet_01v8 ad=7.1721 pd=37.56 as=0 ps=0 w=18.39 l=0.66
X6 VTAIL.t3 VN.t2 VDD2.t1 w_n1564_n4646# sky130_fd_pr__pfet_01v8 ad=7.1721 pd=37.56 as=3.03435 ps=18.72 w=18.39 l=0.66
X7 VTAIL.t6 VP.t1 VDD1.t0 w_n1564_n4646# sky130_fd_pr__pfet_01v8 ad=7.1721 pd=37.56 as=3.03435 ps=18.72 w=18.39 l=0.66
X8 VDD1.t3 VP.t2 VTAIL.t5 w_n1564_n4646# sky130_fd_pr__pfet_01v8 ad=3.03435 pd=18.72 as=7.1721 ps=37.56 w=18.39 l=0.66
X9 VDD1.t2 VP.t3 VTAIL.t4 w_n1564_n4646# sky130_fd_pr__pfet_01v8 ad=3.03435 pd=18.72 as=7.1721 ps=37.56 w=18.39 l=0.66
X10 B.t2 B.t0 B.t1 w_n1564_n4646# sky130_fd_pr__pfet_01v8 ad=7.1721 pd=37.56 as=0 ps=0 w=18.39 l=0.66
X11 VDD2.t0 VN.t3 VTAIL.t0 w_n1564_n4646# sky130_fd_pr__pfet_01v8 ad=3.03435 pd=18.72 as=7.1721 ps=37.56 w=18.39 l=0.66
R0 B.n129 B.t0 875
R1 B.n135 B.t9 875
R2 B.n42 B.t6 875
R3 B.n49 B.t3 875
R4 B.n449 B.n80 585
R5 B.n451 B.n450 585
R6 B.n452 B.n79 585
R7 B.n454 B.n453 585
R8 B.n455 B.n78 585
R9 B.n457 B.n456 585
R10 B.n458 B.n77 585
R11 B.n460 B.n459 585
R12 B.n461 B.n76 585
R13 B.n463 B.n462 585
R14 B.n464 B.n75 585
R15 B.n466 B.n465 585
R16 B.n467 B.n74 585
R17 B.n469 B.n468 585
R18 B.n470 B.n73 585
R19 B.n472 B.n471 585
R20 B.n473 B.n72 585
R21 B.n475 B.n474 585
R22 B.n476 B.n71 585
R23 B.n478 B.n477 585
R24 B.n479 B.n70 585
R25 B.n481 B.n480 585
R26 B.n482 B.n69 585
R27 B.n484 B.n483 585
R28 B.n485 B.n68 585
R29 B.n487 B.n486 585
R30 B.n488 B.n67 585
R31 B.n490 B.n489 585
R32 B.n491 B.n66 585
R33 B.n493 B.n492 585
R34 B.n494 B.n65 585
R35 B.n496 B.n495 585
R36 B.n497 B.n64 585
R37 B.n499 B.n498 585
R38 B.n500 B.n63 585
R39 B.n502 B.n501 585
R40 B.n503 B.n62 585
R41 B.n505 B.n504 585
R42 B.n506 B.n61 585
R43 B.n508 B.n507 585
R44 B.n509 B.n60 585
R45 B.n511 B.n510 585
R46 B.n512 B.n59 585
R47 B.n514 B.n513 585
R48 B.n515 B.n58 585
R49 B.n517 B.n516 585
R50 B.n518 B.n57 585
R51 B.n520 B.n519 585
R52 B.n521 B.n56 585
R53 B.n523 B.n522 585
R54 B.n524 B.n55 585
R55 B.n526 B.n525 585
R56 B.n527 B.n54 585
R57 B.n529 B.n528 585
R58 B.n530 B.n53 585
R59 B.n532 B.n531 585
R60 B.n533 B.n52 585
R61 B.n535 B.n534 585
R62 B.n536 B.n51 585
R63 B.n538 B.n537 585
R64 B.n540 B.n48 585
R65 B.n542 B.n541 585
R66 B.n543 B.n47 585
R67 B.n545 B.n544 585
R68 B.n546 B.n46 585
R69 B.n548 B.n547 585
R70 B.n549 B.n45 585
R71 B.n551 B.n550 585
R72 B.n552 B.n41 585
R73 B.n554 B.n553 585
R74 B.n555 B.n40 585
R75 B.n557 B.n556 585
R76 B.n558 B.n39 585
R77 B.n560 B.n559 585
R78 B.n561 B.n38 585
R79 B.n563 B.n562 585
R80 B.n564 B.n37 585
R81 B.n566 B.n565 585
R82 B.n567 B.n36 585
R83 B.n569 B.n568 585
R84 B.n570 B.n35 585
R85 B.n572 B.n571 585
R86 B.n573 B.n34 585
R87 B.n575 B.n574 585
R88 B.n576 B.n33 585
R89 B.n578 B.n577 585
R90 B.n579 B.n32 585
R91 B.n581 B.n580 585
R92 B.n582 B.n31 585
R93 B.n584 B.n583 585
R94 B.n585 B.n30 585
R95 B.n587 B.n586 585
R96 B.n588 B.n29 585
R97 B.n590 B.n589 585
R98 B.n591 B.n28 585
R99 B.n593 B.n592 585
R100 B.n594 B.n27 585
R101 B.n596 B.n595 585
R102 B.n597 B.n26 585
R103 B.n599 B.n598 585
R104 B.n600 B.n25 585
R105 B.n602 B.n601 585
R106 B.n603 B.n24 585
R107 B.n605 B.n604 585
R108 B.n606 B.n23 585
R109 B.n608 B.n607 585
R110 B.n609 B.n22 585
R111 B.n611 B.n610 585
R112 B.n612 B.n21 585
R113 B.n614 B.n613 585
R114 B.n615 B.n20 585
R115 B.n617 B.n616 585
R116 B.n618 B.n19 585
R117 B.n620 B.n619 585
R118 B.n621 B.n18 585
R119 B.n623 B.n622 585
R120 B.n624 B.n17 585
R121 B.n626 B.n625 585
R122 B.n627 B.n16 585
R123 B.n629 B.n628 585
R124 B.n630 B.n15 585
R125 B.n632 B.n631 585
R126 B.n633 B.n14 585
R127 B.n635 B.n634 585
R128 B.n636 B.n13 585
R129 B.n638 B.n637 585
R130 B.n639 B.n12 585
R131 B.n641 B.n640 585
R132 B.n642 B.n11 585
R133 B.n644 B.n643 585
R134 B.n448 B.n447 585
R135 B.n446 B.n81 585
R136 B.n445 B.n444 585
R137 B.n443 B.n82 585
R138 B.n442 B.n441 585
R139 B.n440 B.n83 585
R140 B.n439 B.n438 585
R141 B.n437 B.n84 585
R142 B.n436 B.n435 585
R143 B.n434 B.n85 585
R144 B.n433 B.n432 585
R145 B.n431 B.n86 585
R146 B.n430 B.n429 585
R147 B.n428 B.n87 585
R148 B.n427 B.n426 585
R149 B.n425 B.n88 585
R150 B.n424 B.n423 585
R151 B.n422 B.n89 585
R152 B.n421 B.n420 585
R153 B.n419 B.n90 585
R154 B.n418 B.n417 585
R155 B.n416 B.n91 585
R156 B.n415 B.n414 585
R157 B.n413 B.n92 585
R158 B.n412 B.n411 585
R159 B.n410 B.n93 585
R160 B.n409 B.n408 585
R161 B.n407 B.n94 585
R162 B.n406 B.n405 585
R163 B.n404 B.n95 585
R164 B.n403 B.n402 585
R165 B.n401 B.n96 585
R166 B.n400 B.n399 585
R167 B.n398 B.n97 585
R168 B.n397 B.n396 585
R169 B.n200 B.n167 585
R170 B.n202 B.n201 585
R171 B.n203 B.n166 585
R172 B.n205 B.n204 585
R173 B.n206 B.n165 585
R174 B.n208 B.n207 585
R175 B.n209 B.n164 585
R176 B.n211 B.n210 585
R177 B.n212 B.n163 585
R178 B.n214 B.n213 585
R179 B.n215 B.n162 585
R180 B.n217 B.n216 585
R181 B.n218 B.n161 585
R182 B.n220 B.n219 585
R183 B.n221 B.n160 585
R184 B.n223 B.n222 585
R185 B.n224 B.n159 585
R186 B.n226 B.n225 585
R187 B.n227 B.n158 585
R188 B.n229 B.n228 585
R189 B.n230 B.n157 585
R190 B.n232 B.n231 585
R191 B.n233 B.n156 585
R192 B.n235 B.n234 585
R193 B.n236 B.n155 585
R194 B.n238 B.n237 585
R195 B.n239 B.n154 585
R196 B.n241 B.n240 585
R197 B.n242 B.n153 585
R198 B.n244 B.n243 585
R199 B.n245 B.n152 585
R200 B.n247 B.n246 585
R201 B.n248 B.n151 585
R202 B.n250 B.n249 585
R203 B.n251 B.n150 585
R204 B.n253 B.n252 585
R205 B.n254 B.n149 585
R206 B.n256 B.n255 585
R207 B.n257 B.n148 585
R208 B.n259 B.n258 585
R209 B.n260 B.n147 585
R210 B.n262 B.n261 585
R211 B.n263 B.n146 585
R212 B.n265 B.n264 585
R213 B.n266 B.n145 585
R214 B.n268 B.n267 585
R215 B.n269 B.n144 585
R216 B.n271 B.n270 585
R217 B.n272 B.n143 585
R218 B.n274 B.n273 585
R219 B.n275 B.n142 585
R220 B.n277 B.n276 585
R221 B.n278 B.n141 585
R222 B.n280 B.n279 585
R223 B.n281 B.n140 585
R224 B.n283 B.n282 585
R225 B.n284 B.n139 585
R226 B.n286 B.n285 585
R227 B.n287 B.n138 585
R228 B.n289 B.n288 585
R229 B.n291 B.n290 585
R230 B.n292 B.n134 585
R231 B.n294 B.n293 585
R232 B.n295 B.n133 585
R233 B.n297 B.n296 585
R234 B.n298 B.n132 585
R235 B.n300 B.n299 585
R236 B.n301 B.n131 585
R237 B.n303 B.n302 585
R238 B.n304 B.n128 585
R239 B.n307 B.n306 585
R240 B.n308 B.n127 585
R241 B.n310 B.n309 585
R242 B.n311 B.n126 585
R243 B.n313 B.n312 585
R244 B.n314 B.n125 585
R245 B.n316 B.n315 585
R246 B.n317 B.n124 585
R247 B.n319 B.n318 585
R248 B.n320 B.n123 585
R249 B.n322 B.n321 585
R250 B.n323 B.n122 585
R251 B.n325 B.n324 585
R252 B.n326 B.n121 585
R253 B.n328 B.n327 585
R254 B.n329 B.n120 585
R255 B.n331 B.n330 585
R256 B.n332 B.n119 585
R257 B.n334 B.n333 585
R258 B.n335 B.n118 585
R259 B.n337 B.n336 585
R260 B.n338 B.n117 585
R261 B.n340 B.n339 585
R262 B.n341 B.n116 585
R263 B.n343 B.n342 585
R264 B.n344 B.n115 585
R265 B.n346 B.n345 585
R266 B.n347 B.n114 585
R267 B.n349 B.n348 585
R268 B.n350 B.n113 585
R269 B.n352 B.n351 585
R270 B.n353 B.n112 585
R271 B.n355 B.n354 585
R272 B.n356 B.n111 585
R273 B.n358 B.n357 585
R274 B.n359 B.n110 585
R275 B.n361 B.n360 585
R276 B.n362 B.n109 585
R277 B.n364 B.n363 585
R278 B.n365 B.n108 585
R279 B.n367 B.n366 585
R280 B.n368 B.n107 585
R281 B.n370 B.n369 585
R282 B.n371 B.n106 585
R283 B.n373 B.n372 585
R284 B.n374 B.n105 585
R285 B.n376 B.n375 585
R286 B.n377 B.n104 585
R287 B.n379 B.n378 585
R288 B.n380 B.n103 585
R289 B.n382 B.n381 585
R290 B.n383 B.n102 585
R291 B.n385 B.n384 585
R292 B.n386 B.n101 585
R293 B.n388 B.n387 585
R294 B.n389 B.n100 585
R295 B.n391 B.n390 585
R296 B.n392 B.n99 585
R297 B.n394 B.n393 585
R298 B.n395 B.n98 585
R299 B.n199 B.n198 585
R300 B.n197 B.n168 585
R301 B.n196 B.n195 585
R302 B.n194 B.n169 585
R303 B.n193 B.n192 585
R304 B.n191 B.n170 585
R305 B.n190 B.n189 585
R306 B.n188 B.n171 585
R307 B.n187 B.n186 585
R308 B.n185 B.n172 585
R309 B.n184 B.n183 585
R310 B.n182 B.n173 585
R311 B.n181 B.n180 585
R312 B.n179 B.n174 585
R313 B.n178 B.n177 585
R314 B.n176 B.n175 585
R315 B.n2 B.n0 585
R316 B.n669 B.n1 585
R317 B.n668 B.n667 585
R318 B.n666 B.n3 585
R319 B.n665 B.n664 585
R320 B.n663 B.n4 585
R321 B.n662 B.n661 585
R322 B.n660 B.n5 585
R323 B.n659 B.n658 585
R324 B.n657 B.n6 585
R325 B.n656 B.n655 585
R326 B.n654 B.n7 585
R327 B.n653 B.n652 585
R328 B.n651 B.n8 585
R329 B.n650 B.n649 585
R330 B.n648 B.n9 585
R331 B.n647 B.n646 585
R332 B.n645 B.n10 585
R333 B.n671 B.n670 585
R334 B.n200 B.n199 506.916
R335 B.n645 B.n644 506.916
R336 B.n397 B.n98 506.916
R337 B.n447 B.n80 506.916
R338 B.n199 B.n168 163.367
R339 B.n195 B.n168 163.367
R340 B.n195 B.n194 163.367
R341 B.n194 B.n193 163.367
R342 B.n193 B.n170 163.367
R343 B.n189 B.n170 163.367
R344 B.n189 B.n188 163.367
R345 B.n188 B.n187 163.367
R346 B.n187 B.n172 163.367
R347 B.n183 B.n172 163.367
R348 B.n183 B.n182 163.367
R349 B.n182 B.n181 163.367
R350 B.n181 B.n174 163.367
R351 B.n177 B.n174 163.367
R352 B.n177 B.n176 163.367
R353 B.n176 B.n2 163.367
R354 B.n670 B.n2 163.367
R355 B.n670 B.n669 163.367
R356 B.n669 B.n668 163.367
R357 B.n668 B.n3 163.367
R358 B.n664 B.n3 163.367
R359 B.n664 B.n663 163.367
R360 B.n663 B.n662 163.367
R361 B.n662 B.n5 163.367
R362 B.n658 B.n5 163.367
R363 B.n658 B.n657 163.367
R364 B.n657 B.n656 163.367
R365 B.n656 B.n7 163.367
R366 B.n652 B.n7 163.367
R367 B.n652 B.n651 163.367
R368 B.n651 B.n650 163.367
R369 B.n650 B.n9 163.367
R370 B.n646 B.n9 163.367
R371 B.n646 B.n645 163.367
R372 B.n201 B.n200 163.367
R373 B.n201 B.n166 163.367
R374 B.n205 B.n166 163.367
R375 B.n206 B.n205 163.367
R376 B.n207 B.n206 163.367
R377 B.n207 B.n164 163.367
R378 B.n211 B.n164 163.367
R379 B.n212 B.n211 163.367
R380 B.n213 B.n212 163.367
R381 B.n213 B.n162 163.367
R382 B.n217 B.n162 163.367
R383 B.n218 B.n217 163.367
R384 B.n219 B.n218 163.367
R385 B.n219 B.n160 163.367
R386 B.n223 B.n160 163.367
R387 B.n224 B.n223 163.367
R388 B.n225 B.n224 163.367
R389 B.n225 B.n158 163.367
R390 B.n229 B.n158 163.367
R391 B.n230 B.n229 163.367
R392 B.n231 B.n230 163.367
R393 B.n231 B.n156 163.367
R394 B.n235 B.n156 163.367
R395 B.n236 B.n235 163.367
R396 B.n237 B.n236 163.367
R397 B.n237 B.n154 163.367
R398 B.n241 B.n154 163.367
R399 B.n242 B.n241 163.367
R400 B.n243 B.n242 163.367
R401 B.n243 B.n152 163.367
R402 B.n247 B.n152 163.367
R403 B.n248 B.n247 163.367
R404 B.n249 B.n248 163.367
R405 B.n249 B.n150 163.367
R406 B.n253 B.n150 163.367
R407 B.n254 B.n253 163.367
R408 B.n255 B.n254 163.367
R409 B.n255 B.n148 163.367
R410 B.n259 B.n148 163.367
R411 B.n260 B.n259 163.367
R412 B.n261 B.n260 163.367
R413 B.n261 B.n146 163.367
R414 B.n265 B.n146 163.367
R415 B.n266 B.n265 163.367
R416 B.n267 B.n266 163.367
R417 B.n267 B.n144 163.367
R418 B.n271 B.n144 163.367
R419 B.n272 B.n271 163.367
R420 B.n273 B.n272 163.367
R421 B.n273 B.n142 163.367
R422 B.n277 B.n142 163.367
R423 B.n278 B.n277 163.367
R424 B.n279 B.n278 163.367
R425 B.n279 B.n140 163.367
R426 B.n283 B.n140 163.367
R427 B.n284 B.n283 163.367
R428 B.n285 B.n284 163.367
R429 B.n285 B.n138 163.367
R430 B.n289 B.n138 163.367
R431 B.n290 B.n289 163.367
R432 B.n290 B.n134 163.367
R433 B.n294 B.n134 163.367
R434 B.n295 B.n294 163.367
R435 B.n296 B.n295 163.367
R436 B.n296 B.n132 163.367
R437 B.n300 B.n132 163.367
R438 B.n301 B.n300 163.367
R439 B.n302 B.n301 163.367
R440 B.n302 B.n128 163.367
R441 B.n307 B.n128 163.367
R442 B.n308 B.n307 163.367
R443 B.n309 B.n308 163.367
R444 B.n309 B.n126 163.367
R445 B.n313 B.n126 163.367
R446 B.n314 B.n313 163.367
R447 B.n315 B.n314 163.367
R448 B.n315 B.n124 163.367
R449 B.n319 B.n124 163.367
R450 B.n320 B.n319 163.367
R451 B.n321 B.n320 163.367
R452 B.n321 B.n122 163.367
R453 B.n325 B.n122 163.367
R454 B.n326 B.n325 163.367
R455 B.n327 B.n326 163.367
R456 B.n327 B.n120 163.367
R457 B.n331 B.n120 163.367
R458 B.n332 B.n331 163.367
R459 B.n333 B.n332 163.367
R460 B.n333 B.n118 163.367
R461 B.n337 B.n118 163.367
R462 B.n338 B.n337 163.367
R463 B.n339 B.n338 163.367
R464 B.n339 B.n116 163.367
R465 B.n343 B.n116 163.367
R466 B.n344 B.n343 163.367
R467 B.n345 B.n344 163.367
R468 B.n345 B.n114 163.367
R469 B.n349 B.n114 163.367
R470 B.n350 B.n349 163.367
R471 B.n351 B.n350 163.367
R472 B.n351 B.n112 163.367
R473 B.n355 B.n112 163.367
R474 B.n356 B.n355 163.367
R475 B.n357 B.n356 163.367
R476 B.n357 B.n110 163.367
R477 B.n361 B.n110 163.367
R478 B.n362 B.n361 163.367
R479 B.n363 B.n362 163.367
R480 B.n363 B.n108 163.367
R481 B.n367 B.n108 163.367
R482 B.n368 B.n367 163.367
R483 B.n369 B.n368 163.367
R484 B.n369 B.n106 163.367
R485 B.n373 B.n106 163.367
R486 B.n374 B.n373 163.367
R487 B.n375 B.n374 163.367
R488 B.n375 B.n104 163.367
R489 B.n379 B.n104 163.367
R490 B.n380 B.n379 163.367
R491 B.n381 B.n380 163.367
R492 B.n381 B.n102 163.367
R493 B.n385 B.n102 163.367
R494 B.n386 B.n385 163.367
R495 B.n387 B.n386 163.367
R496 B.n387 B.n100 163.367
R497 B.n391 B.n100 163.367
R498 B.n392 B.n391 163.367
R499 B.n393 B.n392 163.367
R500 B.n393 B.n98 163.367
R501 B.n398 B.n397 163.367
R502 B.n399 B.n398 163.367
R503 B.n399 B.n96 163.367
R504 B.n403 B.n96 163.367
R505 B.n404 B.n403 163.367
R506 B.n405 B.n404 163.367
R507 B.n405 B.n94 163.367
R508 B.n409 B.n94 163.367
R509 B.n410 B.n409 163.367
R510 B.n411 B.n410 163.367
R511 B.n411 B.n92 163.367
R512 B.n415 B.n92 163.367
R513 B.n416 B.n415 163.367
R514 B.n417 B.n416 163.367
R515 B.n417 B.n90 163.367
R516 B.n421 B.n90 163.367
R517 B.n422 B.n421 163.367
R518 B.n423 B.n422 163.367
R519 B.n423 B.n88 163.367
R520 B.n427 B.n88 163.367
R521 B.n428 B.n427 163.367
R522 B.n429 B.n428 163.367
R523 B.n429 B.n86 163.367
R524 B.n433 B.n86 163.367
R525 B.n434 B.n433 163.367
R526 B.n435 B.n434 163.367
R527 B.n435 B.n84 163.367
R528 B.n439 B.n84 163.367
R529 B.n440 B.n439 163.367
R530 B.n441 B.n440 163.367
R531 B.n441 B.n82 163.367
R532 B.n445 B.n82 163.367
R533 B.n446 B.n445 163.367
R534 B.n447 B.n446 163.367
R535 B.n644 B.n11 163.367
R536 B.n640 B.n11 163.367
R537 B.n640 B.n639 163.367
R538 B.n639 B.n638 163.367
R539 B.n638 B.n13 163.367
R540 B.n634 B.n13 163.367
R541 B.n634 B.n633 163.367
R542 B.n633 B.n632 163.367
R543 B.n632 B.n15 163.367
R544 B.n628 B.n15 163.367
R545 B.n628 B.n627 163.367
R546 B.n627 B.n626 163.367
R547 B.n626 B.n17 163.367
R548 B.n622 B.n17 163.367
R549 B.n622 B.n621 163.367
R550 B.n621 B.n620 163.367
R551 B.n620 B.n19 163.367
R552 B.n616 B.n19 163.367
R553 B.n616 B.n615 163.367
R554 B.n615 B.n614 163.367
R555 B.n614 B.n21 163.367
R556 B.n610 B.n21 163.367
R557 B.n610 B.n609 163.367
R558 B.n609 B.n608 163.367
R559 B.n608 B.n23 163.367
R560 B.n604 B.n23 163.367
R561 B.n604 B.n603 163.367
R562 B.n603 B.n602 163.367
R563 B.n602 B.n25 163.367
R564 B.n598 B.n25 163.367
R565 B.n598 B.n597 163.367
R566 B.n597 B.n596 163.367
R567 B.n596 B.n27 163.367
R568 B.n592 B.n27 163.367
R569 B.n592 B.n591 163.367
R570 B.n591 B.n590 163.367
R571 B.n590 B.n29 163.367
R572 B.n586 B.n29 163.367
R573 B.n586 B.n585 163.367
R574 B.n585 B.n584 163.367
R575 B.n584 B.n31 163.367
R576 B.n580 B.n31 163.367
R577 B.n580 B.n579 163.367
R578 B.n579 B.n578 163.367
R579 B.n578 B.n33 163.367
R580 B.n574 B.n33 163.367
R581 B.n574 B.n573 163.367
R582 B.n573 B.n572 163.367
R583 B.n572 B.n35 163.367
R584 B.n568 B.n35 163.367
R585 B.n568 B.n567 163.367
R586 B.n567 B.n566 163.367
R587 B.n566 B.n37 163.367
R588 B.n562 B.n37 163.367
R589 B.n562 B.n561 163.367
R590 B.n561 B.n560 163.367
R591 B.n560 B.n39 163.367
R592 B.n556 B.n39 163.367
R593 B.n556 B.n555 163.367
R594 B.n555 B.n554 163.367
R595 B.n554 B.n41 163.367
R596 B.n550 B.n41 163.367
R597 B.n550 B.n549 163.367
R598 B.n549 B.n548 163.367
R599 B.n548 B.n46 163.367
R600 B.n544 B.n46 163.367
R601 B.n544 B.n543 163.367
R602 B.n543 B.n542 163.367
R603 B.n542 B.n48 163.367
R604 B.n537 B.n48 163.367
R605 B.n537 B.n536 163.367
R606 B.n536 B.n535 163.367
R607 B.n535 B.n52 163.367
R608 B.n531 B.n52 163.367
R609 B.n531 B.n530 163.367
R610 B.n530 B.n529 163.367
R611 B.n529 B.n54 163.367
R612 B.n525 B.n54 163.367
R613 B.n525 B.n524 163.367
R614 B.n524 B.n523 163.367
R615 B.n523 B.n56 163.367
R616 B.n519 B.n56 163.367
R617 B.n519 B.n518 163.367
R618 B.n518 B.n517 163.367
R619 B.n517 B.n58 163.367
R620 B.n513 B.n58 163.367
R621 B.n513 B.n512 163.367
R622 B.n512 B.n511 163.367
R623 B.n511 B.n60 163.367
R624 B.n507 B.n60 163.367
R625 B.n507 B.n506 163.367
R626 B.n506 B.n505 163.367
R627 B.n505 B.n62 163.367
R628 B.n501 B.n62 163.367
R629 B.n501 B.n500 163.367
R630 B.n500 B.n499 163.367
R631 B.n499 B.n64 163.367
R632 B.n495 B.n64 163.367
R633 B.n495 B.n494 163.367
R634 B.n494 B.n493 163.367
R635 B.n493 B.n66 163.367
R636 B.n489 B.n66 163.367
R637 B.n489 B.n488 163.367
R638 B.n488 B.n487 163.367
R639 B.n487 B.n68 163.367
R640 B.n483 B.n68 163.367
R641 B.n483 B.n482 163.367
R642 B.n482 B.n481 163.367
R643 B.n481 B.n70 163.367
R644 B.n477 B.n70 163.367
R645 B.n477 B.n476 163.367
R646 B.n476 B.n475 163.367
R647 B.n475 B.n72 163.367
R648 B.n471 B.n72 163.367
R649 B.n471 B.n470 163.367
R650 B.n470 B.n469 163.367
R651 B.n469 B.n74 163.367
R652 B.n465 B.n74 163.367
R653 B.n465 B.n464 163.367
R654 B.n464 B.n463 163.367
R655 B.n463 B.n76 163.367
R656 B.n459 B.n76 163.367
R657 B.n459 B.n458 163.367
R658 B.n458 B.n457 163.367
R659 B.n457 B.n78 163.367
R660 B.n453 B.n78 163.367
R661 B.n453 B.n452 163.367
R662 B.n452 B.n451 163.367
R663 B.n451 B.n80 163.367
R664 B.n129 B.t2 125.948
R665 B.n49 B.t4 125.948
R666 B.n135 B.t11 125.924
R667 B.n42 B.t7 125.924
R668 B.n130 B.t1 106.749
R669 B.n50 B.t5 106.749
R670 B.n136 B.t10 106.725
R671 B.n43 B.t8 106.725
R672 B.n305 B.n130 59.5399
R673 B.n137 B.n136 59.5399
R674 B.n44 B.n43 59.5399
R675 B.n539 B.n50 59.5399
R676 B.n643 B.n10 32.9371
R677 B.n449 B.n448 32.9371
R678 B.n396 B.n395 32.9371
R679 B.n198 B.n167 32.9371
R680 B.n130 B.n129 19.2005
R681 B.n136 B.n135 19.2005
R682 B.n43 B.n42 19.2005
R683 B.n50 B.n49 19.2005
R684 B B.n671 18.0485
R685 B.n643 B.n642 10.6151
R686 B.n642 B.n641 10.6151
R687 B.n641 B.n12 10.6151
R688 B.n637 B.n12 10.6151
R689 B.n637 B.n636 10.6151
R690 B.n636 B.n635 10.6151
R691 B.n635 B.n14 10.6151
R692 B.n631 B.n14 10.6151
R693 B.n631 B.n630 10.6151
R694 B.n630 B.n629 10.6151
R695 B.n629 B.n16 10.6151
R696 B.n625 B.n16 10.6151
R697 B.n625 B.n624 10.6151
R698 B.n624 B.n623 10.6151
R699 B.n623 B.n18 10.6151
R700 B.n619 B.n18 10.6151
R701 B.n619 B.n618 10.6151
R702 B.n618 B.n617 10.6151
R703 B.n617 B.n20 10.6151
R704 B.n613 B.n20 10.6151
R705 B.n613 B.n612 10.6151
R706 B.n612 B.n611 10.6151
R707 B.n611 B.n22 10.6151
R708 B.n607 B.n22 10.6151
R709 B.n607 B.n606 10.6151
R710 B.n606 B.n605 10.6151
R711 B.n605 B.n24 10.6151
R712 B.n601 B.n24 10.6151
R713 B.n601 B.n600 10.6151
R714 B.n600 B.n599 10.6151
R715 B.n599 B.n26 10.6151
R716 B.n595 B.n26 10.6151
R717 B.n595 B.n594 10.6151
R718 B.n594 B.n593 10.6151
R719 B.n593 B.n28 10.6151
R720 B.n589 B.n28 10.6151
R721 B.n589 B.n588 10.6151
R722 B.n588 B.n587 10.6151
R723 B.n587 B.n30 10.6151
R724 B.n583 B.n30 10.6151
R725 B.n583 B.n582 10.6151
R726 B.n582 B.n581 10.6151
R727 B.n581 B.n32 10.6151
R728 B.n577 B.n32 10.6151
R729 B.n577 B.n576 10.6151
R730 B.n576 B.n575 10.6151
R731 B.n575 B.n34 10.6151
R732 B.n571 B.n34 10.6151
R733 B.n571 B.n570 10.6151
R734 B.n570 B.n569 10.6151
R735 B.n569 B.n36 10.6151
R736 B.n565 B.n36 10.6151
R737 B.n565 B.n564 10.6151
R738 B.n564 B.n563 10.6151
R739 B.n563 B.n38 10.6151
R740 B.n559 B.n38 10.6151
R741 B.n559 B.n558 10.6151
R742 B.n558 B.n557 10.6151
R743 B.n557 B.n40 10.6151
R744 B.n553 B.n552 10.6151
R745 B.n552 B.n551 10.6151
R746 B.n551 B.n45 10.6151
R747 B.n547 B.n45 10.6151
R748 B.n547 B.n546 10.6151
R749 B.n546 B.n545 10.6151
R750 B.n545 B.n47 10.6151
R751 B.n541 B.n47 10.6151
R752 B.n541 B.n540 10.6151
R753 B.n538 B.n51 10.6151
R754 B.n534 B.n51 10.6151
R755 B.n534 B.n533 10.6151
R756 B.n533 B.n532 10.6151
R757 B.n532 B.n53 10.6151
R758 B.n528 B.n53 10.6151
R759 B.n528 B.n527 10.6151
R760 B.n527 B.n526 10.6151
R761 B.n526 B.n55 10.6151
R762 B.n522 B.n55 10.6151
R763 B.n522 B.n521 10.6151
R764 B.n521 B.n520 10.6151
R765 B.n520 B.n57 10.6151
R766 B.n516 B.n57 10.6151
R767 B.n516 B.n515 10.6151
R768 B.n515 B.n514 10.6151
R769 B.n514 B.n59 10.6151
R770 B.n510 B.n59 10.6151
R771 B.n510 B.n509 10.6151
R772 B.n509 B.n508 10.6151
R773 B.n508 B.n61 10.6151
R774 B.n504 B.n61 10.6151
R775 B.n504 B.n503 10.6151
R776 B.n503 B.n502 10.6151
R777 B.n502 B.n63 10.6151
R778 B.n498 B.n63 10.6151
R779 B.n498 B.n497 10.6151
R780 B.n497 B.n496 10.6151
R781 B.n496 B.n65 10.6151
R782 B.n492 B.n65 10.6151
R783 B.n492 B.n491 10.6151
R784 B.n491 B.n490 10.6151
R785 B.n490 B.n67 10.6151
R786 B.n486 B.n67 10.6151
R787 B.n486 B.n485 10.6151
R788 B.n485 B.n484 10.6151
R789 B.n484 B.n69 10.6151
R790 B.n480 B.n69 10.6151
R791 B.n480 B.n479 10.6151
R792 B.n479 B.n478 10.6151
R793 B.n478 B.n71 10.6151
R794 B.n474 B.n71 10.6151
R795 B.n474 B.n473 10.6151
R796 B.n473 B.n472 10.6151
R797 B.n472 B.n73 10.6151
R798 B.n468 B.n73 10.6151
R799 B.n468 B.n467 10.6151
R800 B.n467 B.n466 10.6151
R801 B.n466 B.n75 10.6151
R802 B.n462 B.n75 10.6151
R803 B.n462 B.n461 10.6151
R804 B.n461 B.n460 10.6151
R805 B.n460 B.n77 10.6151
R806 B.n456 B.n77 10.6151
R807 B.n456 B.n455 10.6151
R808 B.n455 B.n454 10.6151
R809 B.n454 B.n79 10.6151
R810 B.n450 B.n79 10.6151
R811 B.n450 B.n449 10.6151
R812 B.n396 B.n97 10.6151
R813 B.n400 B.n97 10.6151
R814 B.n401 B.n400 10.6151
R815 B.n402 B.n401 10.6151
R816 B.n402 B.n95 10.6151
R817 B.n406 B.n95 10.6151
R818 B.n407 B.n406 10.6151
R819 B.n408 B.n407 10.6151
R820 B.n408 B.n93 10.6151
R821 B.n412 B.n93 10.6151
R822 B.n413 B.n412 10.6151
R823 B.n414 B.n413 10.6151
R824 B.n414 B.n91 10.6151
R825 B.n418 B.n91 10.6151
R826 B.n419 B.n418 10.6151
R827 B.n420 B.n419 10.6151
R828 B.n420 B.n89 10.6151
R829 B.n424 B.n89 10.6151
R830 B.n425 B.n424 10.6151
R831 B.n426 B.n425 10.6151
R832 B.n426 B.n87 10.6151
R833 B.n430 B.n87 10.6151
R834 B.n431 B.n430 10.6151
R835 B.n432 B.n431 10.6151
R836 B.n432 B.n85 10.6151
R837 B.n436 B.n85 10.6151
R838 B.n437 B.n436 10.6151
R839 B.n438 B.n437 10.6151
R840 B.n438 B.n83 10.6151
R841 B.n442 B.n83 10.6151
R842 B.n443 B.n442 10.6151
R843 B.n444 B.n443 10.6151
R844 B.n444 B.n81 10.6151
R845 B.n448 B.n81 10.6151
R846 B.n202 B.n167 10.6151
R847 B.n203 B.n202 10.6151
R848 B.n204 B.n203 10.6151
R849 B.n204 B.n165 10.6151
R850 B.n208 B.n165 10.6151
R851 B.n209 B.n208 10.6151
R852 B.n210 B.n209 10.6151
R853 B.n210 B.n163 10.6151
R854 B.n214 B.n163 10.6151
R855 B.n215 B.n214 10.6151
R856 B.n216 B.n215 10.6151
R857 B.n216 B.n161 10.6151
R858 B.n220 B.n161 10.6151
R859 B.n221 B.n220 10.6151
R860 B.n222 B.n221 10.6151
R861 B.n222 B.n159 10.6151
R862 B.n226 B.n159 10.6151
R863 B.n227 B.n226 10.6151
R864 B.n228 B.n227 10.6151
R865 B.n228 B.n157 10.6151
R866 B.n232 B.n157 10.6151
R867 B.n233 B.n232 10.6151
R868 B.n234 B.n233 10.6151
R869 B.n234 B.n155 10.6151
R870 B.n238 B.n155 10.6151
R871 B.n239 B.n238 10.6151
R872 B.n240 B.n239 10.6151
R873 B.n240 B.n153 10.6151
R874 B.n244 B.n153 10.6151
R875 B.n245 B.n244 10.6151
R876 B.n246 B.n245 10.6151
R877 B.n246 B.n151 10.6151
R878 B.n250 B.n151 10.6151
R879 B.n251 B.n250 10.6151
R880 B.n252 B.n251 10.6151
R881 B.n252 B.n149 10.6151
R882 B.n256 B.n149 10.6151
R883 B.n257 B.n256 10.6151
R884 B.n258 B.n257 10.6151
R885 B.n258 B.n147 10.6151
R886 B.n262 B.n147 10.6151
R887 B.n263 B.n262 10.6151
R888 B.n264 B.n263 10.6151
R889 B.n264 B.n145 10.6151
R890 B.n268 B.n145 10.6151
R891 B.n269 B.n268 10.6151
R892 B.n270 B.n269 10.6151
R893 B.n270 B.n143 10.6151
R894 B.n274 B.n143 10.6151
R895 B.n275 B.n274 10.6151
R896 B.n276 B.n275 10.6151
R897 B.n276 B.n141 10.6151
R898 B.n280 B.n141 10.6151
R899 B.n281 B.n280 10.6151
R900 B.n282 B.n281 10.6151
R901 B.n282 B.n139 10.6151
R902 B.n286 B.n139 10.6151
R903 B.n287 B.n286 10.6151
R904 B.n288 B.n287 10.6151
R905 B.n292 B.n291 10.6151
R906 B.n293 B.n292 10.6151
R907 B.n293 B.n133 10.6151
R908 B.n297 B.n133 10.6151
R909 B.n298 B.n297 10.6151
R910 B.n299 B.n298 10.6151
R911 B.n299 B.n131 10.6151
R912 B.n303 B.n131 10.6151
R913 B.n304 B.n303 10.6151
R914 B.n306 B.n127 10.6151
R915 B.n310 B.n127 10.6151
R916 B.n311 B.n310 10.6151
R917 B.n312 B.n311 10.6151
R918 B.n312 B.n125 10.6151
R919 B.n316 B.n125 10.6151
R920 B.n317 B.n316 10.6151
R921 B.n318 B.n317 10.6151
R922 B.n318 B.n123 10.6151
R923 B.n322 B.n123 10.6151
R924 B.n323 B.n322 10.6151
R925 B.n324 B.n323 10.6151
R926 B.n324 B.n121 10.6151
R927 B.n328 B.n121 10.6151
R928 B.n329 B.n328 10.6151
R929 B.n330 B.n329 10.6151
R930 B.n330 B.n119 10.6151
R931 B.n334 B.n119 10.6151
R932 B.n335 B.n334 10.6151
R933 B.n336 B.n335 10.6151
R934 B.n336 B.n117 10.6151
R935 B.n340 B.n117 10.6151
R936 B.n341 B.n340 10.6151
R937 B.n342 B.n341 10.6151
R938 B.n342 B.n115 10.6151
R939 B.n346 B.n115 10.6151
R940 B.n347 B.n346 10.6151
R941 B.n348 B.n347 10.6151
R942 B.n348 B.n113 10.6151
R943 B.n352 B.n113 10.6151
R944 B.n353 B.n352 10.6151
R945 B.n354 B.n353 10.6151
R946 B.n354 B.n111 10.6151
R947 B.n358 B.n111 10.6151
R948 B.n359 B.n358 10.6151
R949 B.n360 B.n359 10.6151
R950 B.n360 B.n109 10.6151
R951 B.n364 B.n109 10.6151
R952 B.n365 B.n364 10.6151
R953 B.n366 B.n365 10.6151
R954 B.n366 B.n107 10.6151
R955 B.n370 B.n107 10.6151
R956 B.n371 B.n370 10.6151
R957 B.n372 B.n371 10.6151
R958 B.n372 B.n105 10.6151
R959 B.n376 B.n105 10.6151
R960 B.n377 B.n376 10.6151
R961 B.n378 B.n377 10.6151
R962 B.n378 B.n103 10.6151
R963 B.n382 B.n103 10.6151
R964 B.n383 B.n382 10.6151
R965 B.n384 B.n383 10.6151
R966 B.n384 B.n101 10.6151
R967 B.n388 B.n101 10.6151
R968 B.n389 B.n388 10.6151
R969 B.n390 B.n389 10.6151
R970 B.n390 B.n99 10.6151
R971 B.n394 B.n99 10.6151
R972 B.n395 B.n394 10.6151
R973 B.n198 B.n197 10.6151
R974 B.n197 B.n196 10.6151
R975 B.n196 B.n169 10.6151
R976 B.n192 B.n169 10.6151
R977 B.n192 B.n191 10.6151
R978 B.n191 B.n190 10.6151
R979 B.n190 B.n171 10.6151
R980 B.n186 B.n171 10.6151
R981 B.n186 B.n185 10.6151
R982 B.n185 B.n184 10.6151
R983 B.n184 B.n173 10.6151
R984 B.n180 B.n173 10.6151
R985 B.n180 B.n179 10.6151
R986 B.n179 B.n178 10.6151
R987 B.n178 B.n175 10.6151
R988 B.n175 B.n0 10.6151
R989 B.n667 B.n1 10.6151
R990 B.n667 B.n666 10.6151
R991 B.n666 B.n665 10.6151
R992 B.n665 B.n4 10.6151
R993 B.n661 B.n4 10.6151
R994 B.n661 B.n660 10.6151
R995 B.n660 B.n659 10.6151
R996 B.n659 B.n6 10.6151
R997 B.n655 B.n6 10.6151
R998 B.n655 B.n654 10.6151
R999 B.n654 B.n653 10.6151
R1000 B.n653 B.n8 10.6151
R1001 B.n649 B.n8 10.6151
R1002 B.n649 B.n648 10.6151
R1003 B.n648 B.n647 10.6151
R1004 B.n647 B.n10 10.6151
R1005 B.n44 B.n40 9.36635
R1006 B.n539 B.n538 9.36635
R1007 B.n288 B.n137 9.36635
R1008 B.n306 B.n305 9.36635
R1009 B.n671 B.n0 2.81026
R1010 B.n671 B.n1 2.81026
R1011 B.n553 B.n44 1.24928
R1012 B.n540 B.n539 1.24928
R1013 B.n291 B.n137 1.24928
R1014 B.n305 B.n304 1.24928
R1015 VP.n1 VP.t1 752.395
R1016 VP.n1 VP.t2 752.346
R1017 VP.n3 VP.t0 731.399
R1018 VP.n5 VP.t3 731.399
R1019 VP.n6 VP.n5 161.3
R1020 VP.n4 VP.n0 161.3
R1021 VP.n3 VP.n2 161.3
R1022 VP.n2 VP.n1 89.7606
R1023 VP.n4 VP.n3 24.1005
R1024 VP.n5 VP.n4 24.1005
R1025 VP.n2 VP.n0 0.189894
R1026 VP.n6 VP.n0 0.189894
R1027 VP VP.n6 0.0516364
R1028 VDD1 VDD1.n1 113.772
R1029 VDD1 VDD1.n0 71.1759
R1030 VDD1.n0 VDD1.t0 1.76804
R1031 VDD1.n0 VDD1.t3 1.76804
R1032 VDD1.n1 VDD1.t1 1.76804
R1033 VDD1.n1 VDD1.t2 1.76804
R1034 VTAIL.n5 VTAIL.t6 56.2076
R1035 VTAIL.n4 VTAIL.t1 56.2076
R1036 VTAIL.n3 VTAIL.t2 56.2076
R1037 VTAIL.n7 VTAIL.t0 56.2066
R1038 VTAIL.n0 VTAIL.t3 56.2066
R1039 VTAIL.n1 VTAIL.t4 56.2066
R1040 VTAIL.n2 VTAIL.t7 56.2066
R1041 VTAIL.n6 VTAIL.t5 56.2065
R1042 VTAIL.n7 VTAIL.n6 29.0738
R1043 VTAIL.n3 VTAIL.n2 29.0738
R1044 VTAIL.n4 VTAIL.n3 0.853948
R1045 VTAIL.n6 VTAIL.n5 0.853948
R1046 VTAIL.n2 VTAIL.n1 0.853948
R1047 VTAIL VTAIL.n0 0.485414
R1048 VTAIL.n5 VTAIL.n4 0.470328
R1049 VTAIL.n1 VTAIL.n0 0.470328
R1050 VTAIL VTAIL.n7 0.369034
R1051 VN.n0 VN.t2 752.395
R1052 VN.n1 VN.t0 752.395
R1053 VN.n0 VN.t3 752.346
R1054 VN.n1 VN.t1 752.346
R1055 VN VN.n1 90.1413
R1056 VN VN.n0 44.7132
R1057 VDD2.n2 VDD2.n0 113.248
R1058 VDD2.n2 VDD2.n1 71.1177
R1059 VDD2.n1 VDD2.t2 1.76804
R1060 VDD2.n1 VDD2.t3 1.76804
R1061 VDD2.n0 VDD2.t1 1.76804
R1062 VDD2.n0 VDD2.t0 1.76804
R1063 VDD2 VDD2.n2 0.0586897
C0 VDD1 VN 0.147052f
C1 w_n1564_n4646# VN 2.42061f
C2 B VP 1.13006f
C3 VTAIL VDD1 9.85699f
C4 VTAIL w_n1564_n4646# 5.75635f
C5 VDD2 VP 0.270665f
C6 B VDD2 1.11207f
C7 VDD1 VP 4.69115f
C8 VTAIL VN 3.90116f
C9 B VDD1 1.0911f
C10 w_n1564_n4646# VP 2.61676f
C11 B w_n1564_n4646# 8.64988f
C12 VDD2 VDD1 0.557286f
C13 VN VP 5.97977f
C14 VDD2 w_n1564_n4646# 1.23695f
C15 B VN 0.813588f
C16 VTAIL VP 3.91527f
C17 w_n1564_n4646# VDD1 1.22322f
C18 VTAIL B 5.49632f
C19 VDD2 VN 4.56779f
C20 VTAIL VDD2 9.89819f
C21 VDD2 VSUBS 0.827728f
C22 VDD1 VSUBS 5.947123f
C23 VTAIL VSUBS 1.106628f
C24 VN VSUBS 6.45004f
C25 VP VSUBS 1.504129f
C26 B VSUBS 3.125859f
C27 w_n1564_n4646# VSUBS 88.8289f
C28 VDD2.t1 VSUBS 0.416979f
C29 VDD2.t0 VSUBS 0.416979f
C30 VDD2.n0 VSUBS 4.39576f
C31 VDD2.t2 VSUBS 0.416979f
C32 VDD2.t3 VSUBS 0.416979f
C33 VDD2.n1 VSUBS 3.4967f
C34 VDD2.n2 VSUBS 4.85454f
C35 VN.t2 VSUBS 2.03539f
C36 VN.t3 VSUBS 2.03533f
C37 VN.n0 VSUBS 1.47967f
C38 VN.t0 VSUBS 2.03539f
C39 VN.t1 VSUBS 2.03533f
C40 VN.n1 VSUBS 2.92931f
C41 VTAIL.t3 VSUBS 3.4013f
C42 VTAIL.n0 VSUBS 0.693778f
C43 VTAIL.t4 VSUBS 3.4013f
C44 VTAIL.n1 VSUBS 0.720472f
C45 VTAIL.t7 VSUBS 3.4013f
C46 VTAIL.n2 VSUBS 2.20192f
C47 VTAIL.t2 VSUBS 3.4013f
C48 VTAIL.n3 VSUBS 2.20192f
C49 VTAIL.t1 VSUBS 3.4013f
C50 VTAIL.n4 VSUBS 0.720474f
C51 VTAIL.t6 VSUBS 3.4013f
C52 VTAIL.n5 VSUBS 0.720474f
C53 VTAIL.t5 VSUBS 3.40129f
C54 VTAIL.n6 VSUBS 2.20193f
C55 VTAIL.t0 VSUBS 3.4013f
C56 VTAIL.n7 VSUBS 2.1668f
C57 VDD1.t0 VSUBS 0.416808f
C58 VDD1.t3 VSUBS 0.416808f
C59 VDD1.n0 VSUBS 3.4958f
C60 VDD1.t1 VSUBS 0.416808f
C61 VDD1.t2 VSUBS 0.416808f
C62 VDD1.n1 VSUBS 4.42246f
C63 VP.n0 VSUBS 0.059868f
C64 VP.t2 VSUBS 2.0816f
C65 VP.t1 VSUBS 2.08165f
C66 VP.n1 VSUBS 2.97006f
C67 VP.n2 VSUBS 4.26545f
C68 VP.t0 VSUBS 2.06001f
C69 VP.n3 VSUBS 0.771185f
C70 VP.n4 VSUBS 0.013585f
C71 VP.t3 VSUBS 2.06001f
C72 VP.n5 VSUBS 0.771185f
C73 VP.n6 VSUBS 0.046395f
C74 B.n0 VSUBS 0.004886f
C75 B.n1 VSUBS 0.004886f
C76 B.n2 VSUBS 0.007726f
C77 B.n3 VSUBS 0.007726f
C78 B.n4 VSUBS 0.007726f
C79 B.n5 VSUBS 0.007726f
C80 B.n6 VSUBS 0.007726f
C81 B.n7 VSUBS 0.007726f
C82 B.n8 VSUBS 0.007726f
C83 B.n9 VSUBS 0.007726f
C84 B.n10 VSUBS 0.018014f
C85 B.n11 VSUBS 0.007726f
C86 B.n12 VSUBS 0.007726f
C87 B.n13 VSUBS 0.007726f
C88 B.n14 VSUBS 0.007726f
C89 B.n15 VSUBS 0.007726f
C90 B.n16 VSUBS 0.007726f
C91 B.n17 VSUBS 0.007726f
C92 B.n18 VSUBS 0.007726f
C93 B.n19 VSUBS 0.007726f
C94 B.n20 VSUBS 0.007726f
C95 B.n21 VSUBS 0.007726f
C96 B.n22 VSUBS 0.007726f
C97 B.n23 VSUBS 0.007726f
C98 B.n24 VSUBS 0.007726f
C99 B.n25 VSUBS 0.007726f
C100 B.n26 VSUBS 0.007726f
C101 B.n27 VSUBS 0.007726f
C102 B.n28 VSUBS 0.007726f
C103 B.n29 VSUBS 0.007726f
C104 B.n30 VSUBS 0.007726f
C105 B.n31 VSUBS 0.007726f
C106 B.n32 VSUBS 0.007726f
C107 B.n33 VSUBS 0.007726f
C108 B.n34 VSUBS 0.007726f
C109 B.n35 VSUBS 0.007726f
C110 B.n36 VSUBS 0.007726f
C111 B.n37 VSUBS 0.007726f
C112 B.n38 VSUBS 0.007726f
C113 B.n39 VSUBS 0.007726f
C114 B.n40 VSUBS 0.007272f
C115 B.n41 VSUBS 0.007726f
C116 B.t8 VSUBS 0.686236f
C117 B.t7 VSUBS 0.695349f
C118 B.t6 VSUBS 0.537632f
C119 B.n42 VSUBS 0.200833f
C120 B.n43 VSUBS 0.070784f
C121 B.n44 VSUBS 0.017901f
C122 B.n45 VSUBS 0.007726f
C123 B.n46 VSUBS 0.007726f
C124 B.n47 VSUBS 0.007726f
C125 B.n48 VSUBS 0.007726f
C126 B.t5 VSUBS 0.68621f
C127 B.t4 VSUBS 0.695324f
C128 B.t3 VSUBS 0.537632f
C129 B.n49 VSUBS 0.200857f
C130 B.n50 VSUBS 0.070811f
C131 B.n51 VSUBS 0.007726f
C132 B.n52 VSUBS 0.007726f
C133 B.n53 VSUBS 0.007726f
C134 B.n54 VSUBS 0.007726f
C135 B.n55 VSUBS 0.007726f
C136 B.n56 VSUBS 0.007726f
C137 B.n57 VSUBS 0.007726f
C138 B.n58 VSUBS 0.007726f
C139 B.n59 VSUBS 0.007726f
C140 B.n60 VSUBS 0.007726f
C141 B.n61 VSUBS 0.007726f
C142 B.n62 VSUBS 0.007726f
C143 B.n63 VSUBS 0.007726f
C144 B.n64 VSUBS 0.007726f
C145 B.n65 VSUBS 0.007726f
C146 B.n66 VSUBS 0.007726f
C147 B.n67 VSUBS 0.007726f
C148 B.n68 VSUBS 0.007726f
C149 B.n69 VSUBS 0.007726f
C150 B.n70 VSUBS 0.007726f
C151 B.n71 VSUBS 0.007726f
C152 B.n72 VSUBS 0.007726f
C153 B.n73 VSUBS 0.007726f
C154 B.n74 VSUBS 0.007726f
C155 B.n75 VSUBS 0.007726f
C156 B.n76 VSUBS 0.007726f
C157 B.n77 VSUBS 0.007726f
C158 B.n78 VSUBS 0.007726f
C159 B.n79 VSUBS 0.007726f
C160 B.n80 VSUBS 0.018345f
C161 B.n81 VSUBS 0.007726f
C162 B.n82 VSUBS 0.007726f
C163 B.n83 VSUBS 0.007726f
C164 B.n84 VSUBS 0.007726f
C165 B.n85 VSUBS 0.007726f
C166 B.n86 VSUBS 0.007726f
C167 B.n87 VSUBS 0.007726f
C168 B.n88 VSUBS 0.007726f
C169 B.n89 VSUBS 0.007726f
C170 B.n90 VSUBS 0.007726f
C171 B.n91 VSUBS 0.007726f
C172 B.n92 VSUBS 0.007726f
C173 B.n93 VSUBS 0.007726f
C174 B.n94 VSUBS 0.007726f
C175 B.n95 VSUBS 0.007726f
C176 B.n96 VSUBS 0.007726f
C177 B.n97 VSUBS 0.007726f
C178 B.n98 VSUBS 0.018345f
C179 B.n99 VSUBS 0.007726f
C180 B.n100 VSUBS 0.007726f
C181 B.n101 VSUBS 0.007726f
C182 B.n102 VSUBS 0.007726f
C183 B.n103 VSUBS 0.007726f
C184 B.n104 VSUBS 0.007726f
C185 B.n105 VSUBS 0.007726f
C186 B.n106 VSUBS 0.007726f
C187 B.n107 VSUBS 0.007726f
C188 B.n108 VSUBS 0.007726f
C189 B.n109 VSUBS 0.007726f
C190 B.n110 VSUBS 0.007726f
C191 B.n111 VSUBS 0.007726f
C192 B.n112 VSUBS 0.007726f
C193 B.n113 VSUBS 0.007726f
C194 B.n114 VSUBS 0.007726f
C195 B.n115 VSUBS 0.007726f
C196 B.n116 VSUBS 0.007726f
C197 B.n117 VSUBS 0.007726f
C198 B.n118 VSUBS 0.007726f
C199 B.n119 VSUBS 0.007726f
C200 B.n120 VSUBS 0.007726f
C201 B.n121 VSUBS 0.007726f
C202 B.n122 VSUBS 0.007726f
C203 B.n123 VSUBS 0.007726f
C204 B.n124 VSUBS 0.007726f
C205 B.n125 VSUBS 0.007726f
C206 B.n126 VSUBS 0.007726f
C207 B.n127 VSUBS 0.007726f
C208 B.n128 VSUBS 0.007726f
C209 B.t1 VSUBS 0.68621f
C210 B.t2 VSUBS 0.695324f
C211 B.t0 VSUBS 0.537632f
C212 B.n129 VSUBS 0.200857f
C213 B.n130 VSUBS 0.070811f
C214 B.n131 VSUBS 0.007726f
C215 B.n132 VSUBS 0.007726f
C216 B.n133 VSUBS 0.007726f
C217 B.n134 VSUBS 0.007726f
C218 B.t10 VSUBS 0.686236f
C219 B.t11 VSUBS 0.695349f
C220 B.t9 VSUBS 0.537632f
C221 B.n135 VSUBS 0.200833f
C222 B.n136 VSUBS 0.070784f
C223 B.n137 VSUBS 0.017901f
C224 B.n138 VSUBS 0.007726f
C225 B.n139 VSUBS 0.007726f
C226 B.n140 VSUBS 0.007726f
C227 B.n141 VSUBS 0.007726f
C228 B.n142 VSUBS 0.007726f
C229 B.n143 VSUBS 0.007726f
C230 B.n144 VSUBS 0.007726f
C231 B.n145 VSUBS 0.007726f
C232 B.n146 VSUBS 0.007726f
C233 B.n147 VSUBS 0.007726f
C234 B.n148 VSUBS 0.007726f
C235 B.n149 VSUBS 0.007726f
C236 B.n150 VSUBS 0.007726f
C237 B.n151 VSUBS 0.007726f
C238 B.n152 VSUBS 0.007726f
C239 B.n153 VSUBS 0.007726f
C240 B.n154 VSUBS 0.007726f
C241 B.n155 VSUBS 0.007726f
C242 B.n156 VSUBS 0.007726f
C243 B.n157 VSUBS 0.007726f
C244 B.n158 VSUBS 0.007726f
C245 B.n159 VSUBS 0.007726f
C246 B.n160 VSUBS 0.007726f
C247 B.n161 VSUBS 0.007726f
C248 B.n162 VSUBS 0.007726f
C249 B.n163 VSUBS 0.007726f
C250 B.n164 VSUBS 0.007726f
C251 B.n165 VSUBS 0.007726f
C252 B.n166 VSUBS 0.007726f
C253 B.n167 VSUBS 0.018345f
C254 B.n168 VSUBS 0.007726f
C255 B.n169 VSUBS 0.007726f
C256 B.n170 VSUBS 0.007726f
C257 B.n171 VSUBS 0.007726f
C258 B.n172 VSUBS 0.007726f
C259 B.n173 VSUBS 0.007726f
C260 B.n174 VSUBS 0.007726f
C261 B.n175 VSUBS 0.007726f
C262 B.n176 VSUBS 0.007726f
C263 B.n177 VSUBS 0.007726f
C264 B.n178 VSUBS 0.007726f
C265 B.n179 VSUBS 0.007726f
C266 B.n180 VSUBS 0.007726f
C267 B.n181 VSUBS 0.007726f
C268 B.n182 VSUBS 0.007726f
C269 B.n183 VSUBS 0.007726f
C270 B.n184 VSUBS 0.007726f
C271 B.n185 VSUBS 0.007726f
C272 B.n186 VSUBS 0.007726f
C273 B.n187 VSUBS 0.007726f
C274 B.n188 VSUBS 0.007726f
C275 B.n189 VSUBS 0.007726f
C276 B.n190 VSUBS 0.007726f
C277 B.n191 VSUBS 0.007726f
C278 B.n192 VSUBS 0.007726f
C279 B.n193 VSUBS 0.007726f
C280 B.n194 VSUBS 0.007726f
C281 B.n195 VSUBS 0.007726f
C282 B.n196 VSUBS 0.007726f
C283 B.n197 VSUBS 0.007726f
C284 B.n198 VSUBS 0.018014f
C285 B.n199 VSUBS 0.018014f
C286 B.n200 VSUBS 0.018345f
C287 B.n201 VSUBS 0.007726f
C288 B.n202 VSUBS 0.007726f
C289 B.n203 VSUBS 0.007726f
C290 B.n204 VSUBS 0.007726f
C291 B.n205 VSUBS 0.007726f
C292 B.n206 VSUBS 0.007726f
C293 B.n207 VSUBS 0.007726f
C294 B.n208 VSUBS 0.007726f
C295 B.n209 VSUBS 0.007726f
C296 B.n210 VSUBS 0.007726f
C297 B.n211 VSUBS 0.007726f
C298 B.n212 VSUBS 0.007726f
C299 B.n213 VSUBS 0.007726f
C300 B.n214 VSUBS 0.007726f
C301 B.n215 VSUBS 0.007726f
C302 B.n216 VSUBS 0.007726f
C303 B.n217 VSUBS 0.007726f
C304 B.n218 VSUBS 0.007726f
C305 B.n219 VSUBS 0.007726f
C306 B.n220 VSUBS 0.007726f
C307 B.n221 VSUBS 0.007726f
C308 B.n222 VSUBS 0.007726f
C309 B.n223 VSUBS 0.007726f
C310 B.n224 VSUBS 0.007726f
C311 B.n225 VSUBS 0.007726f
C312 B.n226 VSUBS 0.007726f
C313 B.n227 VSUBS 0.007726f
C314 B.n228 VSUBS 0.007726f
C315 B.n229 VSUBS 0.007726f
C316 B.n230 VSUBS 0.007726f
C317 B.n231 VSUBS 0.007726f
C318 B.n232 VSUBS 0.007726f
C319 B.n233 VSUBS 0.007726f
C320 B.n234 VSUBS 0.007726f
C321 B.n235 VSUBS 0.007726f
C322 B.n236 VSUBS 0.007726f
C323 B.n237 VSUBS 0.007726f
C324 B.n238 VSUBS 0.007726f
C325 B.n239 VSUBS 0.007726f
C326 B.n240 VSUBS 0.007726f
C327 B.n241 VSUBS 0.007726f
C328 B.n242 VSUBS 0.007726f
C329 B.n243 VSUBS 0.007726f
C330 B.n244 VSUBS 0.007726f
C331 B.n245 VSUBS 0.007726f
C332 B.n246 VSUBS 0.007726f
C333 B.n247 VSUBS 0.007726f
C334 B.n248 VSUBS 0.007726f
C335 B.n249 VSUBS 0.007726f
C336 B.n250 VSUBS 0.007726f
C337 B.n251 VSUBS 0.007726f
C338 B.n252 VSUBS 0.007726f
C339 B.n253 VSUBS 0.007726f
C340 B.n254 VSUBS 0.007726f
C341 B.n255 VSUBS 0.007726f
C342 B.n256 VSUBS 0.007726f
C343 B.n257 VSUBS 0.007726f
C344 B.n258 VSUBS 0.007726f
C345 B.n259 VSUBS 0.007726f
C346 B.n260 VSUBS 0.007726f
C347 B.n261 VSUBS 0.007726f
C348 B.n262 VSUBS 0.007726f
C349 B.n263 VSUBS 0.007726f
C350 B.n264 VSUBS 0.007726f
C351 B.n265 VSUBS 0.007726f
C352 B.n266 VSUBS 0.007726f
C353 B.n267 VSUBS 0.007726f
C354 B.n268 VSUBS 0.007726f
C355 B.n269 VSUBS 0.007726f
C356 B.n270 VSUBS 0.007726f
C357 B.n271 VSUBS 0.007726f
C358 B.n272 VSUBS 0.007726f
C359 B.n273 VSUBS 0.007726f
C360 B.n274 VSUBS 0.007726f
C361 B.n275 VSUBS 0.007726f
C362 B.n276 VSUBS 0.007726f
C363 B.n277 VSUBS 0.007726f
C364 B.n278 VSUBS 0.007726f
C365 B.n279 VSUBS 0.007726f
C366 B.n280 VSUBS 0.007726f
C367 B.n281 VSUBS 0.007726f
C368 B.n282 VSUBS 0.007726f
C369 B.n283 VSUBS 0.007726f
C370 B.n284 VSUBS 0.007726f
C371 B.n285 VSUBS 0.007726f
C372 B.n286 VSUBS 0.007726f
C373 B.n287 VSUBS 0.007726f
C374 B.n288 VSUBS 0.007272f
C375 B.n289 VSUBS 0.007726f
C376 B.n290 VSUBS 0.007726f
C377 B.n291 VSUBS 0.004318f
C378 B.n292 VSUBS 0.007726f
C379 B.n293 VSUBS 0.007726f
C380 B.n294 VSUBS 0.007726f
C381 B.n295 VSUBS 0.007726f
C382 B.n296 VSUBS 0.007726f
C383 B.n297 VSUBS 0.007726f
C384 B.n298 VSUBS 0.007726f
C385 B.n299 VSUBS 0.007726f
C386 B.n300 VSUBS 0.007726f
C387 B.n301 VSUBS 0.007726f
C388 B.n302 VSUBS 0.007726f
C389 B.n303 VSUBS 0.007726f
C390 B.n304 VSUBS 0.004318f
C391 B.n305 VSUBS 0.017901f
C392 B.n306 VSUBS 0.007272f
C393 B.n307 VSUBS 0.007726f
C394 B.n308 VSUBS 0.007726f
C395 B.n309 VSUBS 0.007726f
C396 B.n310 VSUBS 0.007726f
C397 B.n311 VSUBS 0.007726f
C398 B.n312 VSUBS 0.007726f
C399 B.n313 VSUBS 0.007726f
C400 B.n314 VSUBS 0.007726f
C401 B.n315 VSUBS 0.007726f
C402 B.n316 VSUBS 0.007726f
C403 B.n317 VSUBS 0.007726f
C404 B.n318 VSUBS 0.007726f
C405 B.n319 VSUBS 0.007726f
C406 B.n320 VSUBS 0.007726f
C407 B.n321 VSUBS 0.007726f
C408 B.n322 VSUBS 0.007726f
C409 B.n323 VSUBS 0.007726f
C410 B.n324 VSUBS 0.007726f
C411 B.n325 VSUBS 0.007726f
C412 B.n326 VSUBS 0.007726f
C413 B.n327 VSUBS 0.007726f
C414 B.n328 VSUBS 0.007726f
C415 B.n329 VSUBS 0.007726f
C416 B.n330 VSUBS 0.007726f
C417 B.n331 VSUBS 0.007726f
C418 B.n332 VSUBS 0.007726f
C419 B.n333 VSUBS 0.007726f
C420 B.n334 VSUBS 0.007726f
C421 B.n335 VSUBS 0.007726f
C422 B.n336 VSUBS 0.007726f
C423 B.n337 VSUBS 0.007726f
C424 B.n338 VSUBS 0.007726f
C425 B.n339 VSUBS 0.007726f
C426 B.n340 VSUBS 0.007726f
C427 B.n341 VSUBS 0.007726f
C428 B.n342 VSUBS 0.007726f
C429 B.n343 VSUBS 0.007726f
C430 B.n344 VSUBS 0.007726f
C431 B.n345 VSUBS 0.007726f
C432 B.n346 VSUBS 0.007726f
C433 B.n347 VSUBS 0.007726f
C434 B.n348 VSUBS 0.007726f
C435 B.n349 VSUBS 0.007726f
C436 B.n350 VSUBS 0.007726f
C437 B.n351 VSUBS 0.007726f
C438 B.n352 VSUBS 0.007726f
C439 B.n353 VSUBS 0.007726f
C440 B.n354 VSUBS 0.007726f
C441 B.n355 VSUBS 0.007726f
C442 B.n356 VSUBS 0.007726f
C443 B.n357 VSUBS 0.007726f
C444 B.n358 VSUBS 0.007726f
C445 B.n359 VSUBS 0.007726f
C446 B.n360 VSUBS 0.007726f
C447 B.n361 VSUBS 0.007726f
C448 B.n362 VSUBS 0.007726f
C449 B.n363 VSUBS 0.007726f
C450 B.n364 VSUBS 0.007726f
C451 B.n365 VSUBS 0.007726f
C452 B.n366 VSUBS 0.007726f
C453 B.n367 VSUBS 0.007726f
C454 B.n368 VSUBS 0.007726f
C455 B.n369 VSUBS 0.007726f
C456 B.n370 VSUBS 0.007726f
C457 B.n371 VSUBS 0.007726f
C458 B.n372 VSUBS 0.007726f
C459 B.n373 VSUBS 0.007726f
C460 B.n374 VSUBS 0.007726f
C461 B.n375 VSUBS 0.007726f
C462 B.n376 VSUBS 0.007726f
C463 B.n377 VSUBS 0.007726f
C464 B.n378 VSUBS 0.007726f
C465 B.n379 VSUBS 0.007726f
C466 B.n380 VSUBS 0.007726f
C467 B.n381 VSUBS 0.007726f
C468 B.n382 VSUBS 0.007726f
C469 B.n383 VSUBS 0.007726f
C470 B.n384 VSUBS 0.007726f
C471 B.n385 VSUBS 0.007726f
C472 B.n386 VSUBS 0.007726f
C473 B.n387 VSUBS 0.007726f
C474 B.n388 VSUBS 0.007726f
C475 B.n389 VSUBS 0.007726f
C476 B.n390 VSUBS 0.007726f
C477 B.n391 VSUBS 0.007726f
C478 B.n392 VSUBS 0.007726f
C479 B.n393 VSUBS 0.007726f
C480 B.n394 VSUBS 0.007726f
C481 B.n395 VSUBS 0.018345f
C482 B.n396 VSUBS 0.018014f
C483 B.n397 VSUBS 0.018014f
C484 B.n398 VSUBS 0.007726f
C485 B.n399 VSUBS 0.007726f
C486 B.n400 VSUBS 0.007726f
C487 B.n401 VSUBS 0.007726f
C488 B.n402 VSUBS 0.007726f
C489 B.n403 VSUBS 0.007726f
C490 B.n404 VSUBS 0.007726f
C491 B.n405 VSUBS 0.007726f
C492 B.n406 VSUBS 0.007726f
C493 B.n407 VSUBS 0.007726f
C494 B.n408 VSUBS 0.007726f
C495 B.n409 VSUBS 0.007726f
C496 B.n410 VSUBS 0.007726f
C497 B.n411 VSUBS 0.007726f
C498 B.n412 VSUBS 0.007726f
C499 B.n413 VSUBS 0.007726f
C500 B.n414 VSUBS 0.007726f
C501 B.n415 VSUBS 0.007726f
C502 B.n416 VSUBS 0.007726f
C503 B.n417 VSUBS 0.007726f
C504 B.n418 VSUBS 0.007726f
C505 B.n419 VSUBS 0.007726f
C506 B.n420 VSUBS 0.007726f
C507 B.n421 VSUBS 0.007726f
C508 B.n422 VSUBS 0.007726f
C509 B.n423 VSUBS 0.007726f
C510 B.n424 VSUBS 0.007726f
C511 B.n425 VSUBS 0.007726f
C512 B.n426 VSUBS 0.007726f
C513 B.n427 VSUBS 0.007726f
C514 B.n428 VSUBS 0.007726f
C515 B.n429 VSUBS 0.007726f
C516 B.n430 VSUBS 0.007726f
C517 B.n431 VSUBS 0.007726f
C518 B.n432 VSUBS 0.007726f
C519 B.n433 VSUBS 0.007726f
C520 B.n434 VSUBS 0.007726f
C521 B.n435 VSUBS 0.007726f
C522 B.n436 VSUBS 0.007726f
C523 B.n437 VSUBS 0.007726f
C524 B.n438 VSUBS 0.007726f
C525 B.n439 VSUBS 0.007726f
C526 B.n440 VSUBS 0.007726f
C527 B.n441 VSUBS 0.007726f
C528 B.n442 VSUBS 0.007726f
C529 B.n443 VSUBS 0.007726f
C530 B.n444 VSUBS 0.007726f
C531 B.n445 VSUBS 0.007726f
C532 B.n446 VSUBS 0.007726f
C533 B.n447 VSUBS 0.018014f
C534 B.n448 VSUBS 0.018919f
C535 B.n449 VSUBS 0.01744f
C536 B.n450 VSUBS 0.007726f
C537 B.n451 VSUBS 0.007726f
C538 B.n452 VSUBS 0.007726f
C539 B.n453 VSUBS 0.007726f
C540 B.n454 VSUBS 0.007726f
C541 B.n455 VSUBS 0.007726f
C542 B.n456 VSUBS 0.007726f
C543 B.n457 VSUBS 0.007726f
C544 B.n458 VSUBS 0.007726f
C545 B.n459 VSUBS 0.007726f
C546 B.n460 VSUBS 0.007726f
C547 B.n461 VSUBS 0.007726f
C548 B.n462 VSUBS 0.007726f
C549 B.n463 VSUBS 0.007726f
C550 B.n464 VSUBS 0.007726f
C551 B.n465 VSUBS 0.007726f
C552 B.n466 VSUBS 0.007726f
C553 B.n467 VSUBS 0.007726f
C554 B.n468 VSUBS 0.007726f
C555 B.n469 VSUBS 0.007726f
C556 B.n470 VSUBS 0.007726f
C557 B.n471 VSUBS 0.007726f
C558 B.n472 VSUBS 0.007726f
C559 B.n473 VSUBS 0.007726f
C560 B.n474 VSUBS 0.007726f
C561 B.n475 VSUBS 0.007726f
C562 B.n476 VSUBS 0.007726f
C563 B.n477 VSUBS 0.007726f
C564 B.n478 VSUBS 0.007726f
C565 B.n479 VSUBS 0.007726f
C566 B.n480 VSUBS 0.007726f
C567 B.n481 VSUBS 0.007726f
C568 B.n482 VSUBS 0.007726f
C569 B.n483 VSUBS 0.007726f
C570 B.n484 VSUBS 0.007726f
C571 B.n485 VSUBS 0.007726f
C572 B.n486 VSUBS 0.007726f
C573 B.n487 VSUBS 0.007726f
C574 B.n488 VSUBS 0.007726f
C575 B.n489 VSUBS 0.007726f
C576 B.n490 VSUBS 0.007726f
C577 B.n491 VSUBS 0.007726f
C578 B.n492 VSUBS 0.007726f
C579 B.n493 VSUBS 0.007726f
C580 B.n494 VSUBS 0.007726f
C581 B.n495 VSUBS 0.007726f
C582 B.n496 VSUBS 0.007726f
C583 B.n497 VSUBS 0.007726f
C584 B.n498 VSUBS 0.007726f
C585 B.n499 VSUBS 0.007726f
C586 B.n500 VSUBS 0.007726f
C587 B.n501 VSUBS 0.007726f
C588 B.n502 VSUBS 0.007726f
C589 B.n503 VSUBS 0.007726f
C590 B.n504 VSUBS 0.007726f
C591 B.n505 VSUBS 0.007726f
C592 B.n506 VSUBS 0.007726f
C593 B.n507 VSUBS 0.007726f
C594 B.n508 VSUBS 0.007726f
C595 B.n509 VSUBS 0.007726f
C596 B.n510 VSUBS 0.007726f
C597 B.n511 VSUBS 0.007726f
C598 B.n512 VSUBS 0.007726f
C599 B.n513 VSUBS 0.007726f
C600 B.n514 VSUBS 0.007726f
C601 B.n515 VSUBS 0.007726f
C602 B.n516 VSUBS 0.007726f
C603 B.n517 VSUBS 0.007726f
C604 B.n518 VSUBS 0.007726f
C605 B.n519 VSUBS 0.007726f
C606 B.n520 VSUBS 0.007726f
C607 B.n521 VSUBS 0.007726f
C608 B.n522 VSUBS 0.007726f
C609 B.n523 VSUBS 0.007726f
C610 B.n524 VSUBS 0.007726f
C611 B.n525 VSUBS 0.007726f
C612 B.n526 VSUBS 0.007726f
C613 B.n527 VSUBS 0.007726f
C614 B.n528 VSUBS 0.007726f
C615 B.n529 VSUBS 0.007726f
C616 B.n530 VSUBS 0.007726f
C617 B.n531 VSUBS 0.007726f
C618 B.n532 VSUBS 0.007726f
C619 B.n533 VSUBS 0.007726f
C620 B.n534 VSUBS 0.007726f
C621 B.n535 VSUBS 0.007726f
C622 B.n536 VSUBS 0.007726f
C623 B.n537 VSUBS 0.007726f
C624 B.n538 VSUBS 0.007272f
C625 B.n539 VSUBS 0.017901f
C626 B.n540 VSUBS 0.004318f
C627 B.n541 VSUBS 0.007726f
C628 B.n542 VSUBS 0.007726f
C629 B.n543 VSUBS 0.007726f
C630 B.n544 VSUBS 0.007726f
C631 B.n545 VSUBS 0.007726f
C632 B.n546 VSUBS 0.007726f
C633 B.n547 VSUBS 0.007726f
C634 B.n548 VSUBS 0.007726f
C635 B.n549 VSUBS 0.007726f
C636 B.n550 VSUBS 0.007726f
C637 B.n551 VSUBS 0.007726f
C638 B.n552 VSUBS 0.007726f
C639 B.n553 VSUBS 0.004318f
C640 B.n554 VSUBS 0.007726f
C641 B.n555 VSUBS 0.007726f
C642 B.n556 VSUBS 0.007726f
C643 B.n557 VSUBS 0.007726f
C644 B.n558 VSUBS 0.007726f
C645 B.n559 VSUBS 0.007726f
C646 B.n560 VSUBS 0.007726f
C647 B.n561 VSUBS 0.007726f
C648 B.n562 VSUBS 0.007726f
C649 B.n563 VSUBS 0.007726f
C650 B.n564 VSUBS 0.007726f
C651 B.n565 VSUBS 0.007726f
C652 B.n566 VSUBS 0.007726f
C653 B.n567 VSUBS 0.007726f
C654 B.n568 VSUBS 0.007726f
C655 B.n569 VSUBS 0.007726f
C656 B.n570 VSUBS 0.007726f
C657 B.n571 VSUBS 0.007726f
C658 B.n572 VSUBS 0.007726f
C659 B.n573 VSUBS 0.007726f
C660 B.n574 VSUBS 0.007726f
C661 B.n575 VSUBS 0.007726f
C662 B.n576 VSUBS 0.007726f
C663 B.n577 VSUBS 0.007726f
C664 B.n578 VSUBS 0.007726f
C665 B.n579 VSUBS 0.007726f
C666 B.n580 VSUBS 0.007726f
C667 B.n581 VSUBS 0.007726f
C668 B.n582 VSUBS 0.007726f
C669 B.n583 VSUBS 0.007726f
C670 B.n584 VSUBS 0.007726f
C671 B.n585 VSUBS 0.007726f
C672 B.n586 VSUBS 0.007726f
C673 B.n587 VSUBS 0.007726f
C674 B.n588 VSUBS 0.007726f
C675 B.n589 VSUBS 0.007726f
C676 B.n590 VSUBS 0.007726f
C677 B.n591 VSUBS 0.007726f
C678 B.n592 VSUBS 0.007726f
C679 B.n593 VSUBS 0.007726f
C680 B.n594 VSUBS 0.007726f
C681 B.n595 VSUBS 0.007726f
C682 B.n596 VSUBS 0.007726f
C683 B.n597 VSUBS 0.007726f
C684 B.n598 VSUBS 0.007726f
C685 B.n599 VSUBS 0.007726f
C686 B.n600 VSUBS 0.007726f
C687 B.n601 VSUBS 0.007726f
C688 B.n602 VSUBS 0.007726f
C689 B.n603 VSUBS 0.007726f
C690 B.n604 VSUBS 0.007726f
C691 B.n605 VSUBS 0.007726f
C692 B.n606 VSUBS 0.007726f
C693 B.n607 VSUBS 0.007726f
C694 B.n608 VSUBS 0.007726f
C695 B.n609 VSUBS 0.007726f
C696 B.n610 VSUBS 0.007726f
C697 B.n611 VSUBS 0.007726f
C698 B.n612 VSUBS 0.007726f
C699 B.n613 VSUBS 0.007726f
C700 B.n614 VSUBS 0.007726f
C701 B.n615 VSUBS 0.007726f
C702 B.n616 VSUBS 0.007726f
C703 B.n617 VSUBS 0.007726f
C704 B.n618 VSUBS 0.007726f
C705 B.n619 VSUBS 0.007726f
C706 B.n620 VSUBS 0.007726f
C707 B.n621 VSUBS 0.007726f
C708 B.n622 VSUBS 0.007726f
C709 B.n623 VSUBS 0.007726f
C710 B.n624 VSUBS 0.007726f
C711 B.n625 VSUBS 0.007726f
C712 B.n626 VSUBS 0.007726f
C713 B.n627 VSUBS 0.007726f
C714 B.n628 VSUBS 0.007726f
C715 B.n629 VSUBS 0.007726f
C716 B.n630 VSUBS 0.007726f
C717 B.n631 VSUBS 0.007726f
C718 B.n632 VSUBS 0.007726f
C719 B.n633 VSUBS 0.007726f
C720 B.n634 VSUBS 0.007726f
C721 B.n635 VSUBS 0.007726f
C722 B.n636 VSUBS 0.007726f
C723 B.n637 VSUBS 0.007726f
C724 B.n638 VSUBS 0.007726f
C725 B.n639 VSUBS 0.007726f
C726 B.n640 VSUBS 0.007726f
C727 B.n641 VSUBS 0.007726f
C728 B.n642 VSUBS 0.007726f
C729 B.n643 VSUBS 0.018345f
C730 B.n644 VSUBS 0.018345f
C731 B.n645 VSUBS 0.018014f
C732 B.n646 VSUBS 0.007726f
C733 B.n647 VSUBS 0.007726f
C734 B.n648 VSUBS 0.007726f
C735 B.n649 VSUBS 0.007726f
C736 B.n650 VSUBS 0.007726f
C737 B.n651 VSUBS 0.007726f
C738 B.n652 VSUBS 0.007726f
C739 B.n653 VSUBS 0.007726f
C740 B.n654 VSUBS 0.007726f
C741 B.n655 VSUBS 0.007726f
C742 B.n656 VSUBS 0.007726f
C743 B.n657 VSUBS 0.007726f
C744 B.n658 VSUBS 0.007726f
C745 B.n659 VSUBS 0.007726f
C746 B.n660 VSUBS 0.007726f
C747 B.n661 VSUBS 0.007726f
C748 B.n662 VSUBS 0.007726f
C749 B.n663 VSUBS 0.007726f
C750 B.n664 VSUBS 0.007726f
C751 B.n665 VSUBS 0.007726f
C752 B.n666 VSUBS 0.007726f
C753 B.n667 VSUBS 0.007726f
C754 B.n668 VSUBS 0.007726f
C755 B.n669 VSUBS 0.007726f
C756 B.n670 VSUBS 0.007726f
C757 B.n671 VSUBS 0.017495f
.ends

