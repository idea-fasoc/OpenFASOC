* NGSPICE file created from diff_pair_sample_1750.ext - technology: sky130A

.subckt diff_pair_sample_1750 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=6.3453 pd=33.32 as=2.68455 ps=16.6 w=16.27 l=2.35
X1 VDD1.t2 VP.t1 VTAIL.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=2.68455 pd=16.6 as=6.3453 ps=33.32 w=16.27 l=2.35
X2 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=6.3453 pd=33.32 as=0 ps=0 w=16.27 l=2.35
X3 VDD1.t5 VP.t2 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=2.68455 pd=16.6 as=2.68455 ps=16.6 w=16.27 l=2.35
X4 VTAIL.t12 VP.t3 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=2.68455 pd=16.6 as=2.68455 ps=16.6 w=16.27 l=2.35
X5 VTAIL.t6 VN.t0 VDD2.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=6.3453 pd=33.32 as=2.68455 ps=16.6 w=16.27 l=2.35
X6 VDD1.t1 VP.t4 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=2.68455 pd=16.6 as=6.3453 ps=33.32 w=16.27 l=2.35
X7 VTAIL.t10 VP.t5 VDD1.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=2.68455 pd=16.6 as=2.68455 ps=16.6 w=16.27 l=2.35
X8 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=6.3453 pd=33.32 as=0 ps=0 w=16.27 l=2.35
X9 VTAIL.t7 VN.t1 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=2.68455 pd=16.6 as=2.68455 ps=16.6 w=16.27 l=2.35
X10 VDD1.t7 VP.t6 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=2.68455 pd=16.6 as=2.68455 ps=16.6 w=16.27 l=2.35
X11 VDD2.t5 VN.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.68455 pd=16.6 as=2.68455 ps=16.6 w=16.27 l=2.35
X12 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=6.3453 pd=33.32 as=0 ps=0 w=16.27 l=2.35
X13 VDD2.t4 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.68455 pd=16.6 as=6.3453 ps=33.32 w=16.27 l=2.35
X14 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.3453 pd=33.32 as=0 ps=0 w=16.27 l=2.35
X15 VTAIL.t2 VN.t4 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=2.68455 pd=16.6 as=2.68455 ps=16.6 w=16.27 l=2.35
X16 VTAIL.t8 VP.t7 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=6.3453 pd=33.32 as=2.68455 ps=16.6 w=16.27 l=2.35
X17 VDD2.t2 VN.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.68455 pd=16.6 as=2.68455 ps=16.6 w=16.27 l=2.35
X18 VTAIL.t1 VN.t6 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.3453 pd=33.32 as=2.68455 ps=16.6 w=16.27 l=2.35
X19 VDD2.t0 VN.t7 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.68455 pd=16.6 as=6.3453 ps=33.32 w=16.27 l=2.35
R0 VP.n15 VP.t7 198.825
R1 VP.n36 VP.t0 166.855
R2 VP.n43 VP.t2 166.855
R3 VP.n55 VP.t5 166.855
R4 VP.n63 VP.t4 166.855
R5 VP.n33 VP.t1 166.855
R6 VP.n25 VP.t3 166.855
R7 VP.n14 VP.t6 166.855
R8 VP.n16 VP.n13 161.3
R9 VP.n18 VP.n17 161.3
R10 VP.n19 VP.n12 161.3
R11 VP.n21 VP.n20 161.3
R12 VP.n22 VP.n11 161.3
R13 VP.n24 VP.n23 161.3
R14 VP.n26 VP.n10 161.3
R15 VP.n28 VP.n27 161.3
R16 VP.n29 VP.n9 161.3
R17 VP.n31 VP.n30 161.3
R18 VP.n32 VP.n8 161.3
R19 VP.n62 VP.n0 161.3
R20 VP.n61 VP.n60 161.3
R21 VP.n59 VP.n1 161.3
R22 VP.n58 VP.n57 161.3
R23 VP.n56 VP.n2 161.3
R24 VP.n54 VP.n53 161.3
R25 VP.n52 VP.n3 161.3
R26 VP.n51 VP.n50 161.3
R27 VP.n49 VP.n4 161.3
R28 VP.n48 VP.n47 161.3
R29 VP.n46 VP.n5 161.3
R30 VP.n45 VP.n44 161.3
R31 VP.n42 VP.n6 161.3
R32 VP.n41 VP.n40 161.3
R33 VP.n39 VP.n7 161.3
R34 VP.n38 VP.n37 161.3
R35 VP.n36 VP.n35 97.5443
R36 VP.n64 VP.n63 97.5443
R37 VP.n34 VP.n33 97.5443
R38 VP.n15 VP.n14 67.7723
R39 VP.n50 VP.n49 56.5193
R40 VP.n20 VP.n19 56.5193
R41 VP.n35 VP.n34 52.9693
R42 VP.n42 VP.n41 47.2923
R43 VP.n57 VP.n1 47.2923
R44 VP.n27 VP.n9 47.2923
R45 VP.n41 VP.n7 33.6945
R46 VP.n61 VP.n1 33.6945
R47 VP.n31 VP.n9 33.6945
R48 VP.n37 VP.n7 24.4675
R49 VP.n44 VP.n42 24.4675
R50 VP.n48 VP.n5 24.4675
R51 VP.n49 VP.n48 24.4675
R52 VP.n50 VP.n3 24.4675
R53 VP.n54 VP.n3 24.4675
R54 VP.n57 VP.n56 24.4675
R55 VP.n62 VP.n61 24.4675
R56 VP.n32 VP.n31 24.4675
R57 VP.n20 VP.n11 24.4675
R58 VP.n24 VP.n11 24.4675
R59 VP.n27 VP.n26 24.4675
R60 VP.n18 VP.n13 24.4675
R61 VP.n19 VP.n18 24.4675
R62 VP.n44 VP.n43 20.0634
R63 VP.n56 VP.n55 20.0634
R64 VP.n26 VP.n25 20.0634
R65 VP.n37 VP.n36 13.2127
R66 VP.n63 VP.n62 13.2127
R67 VP.n33 VP.n32 13.2127
R68 VP.n16 VP.n15 9.67836
R69 VP.n43 VP.n5 4.40456
R70 VP.n55 VP.n54 4.40456
R71 VP.n25 VP.n24 4.40456
R72 VP.n14 VP.n13 4.40456
R73 VP.n34 VP.n8 0.278367
R74 VP.n38 VP.n35 0.278367
R75 VP.n64 VP.n0 0.278367
R76 VP.n17 VP.n16 0.189894
R77 VP.n17 VP.n12 0.189894
R78 VP.n21 VP.n12 0.189894
R79 VP.n22 VP.n21 0.189894
R80 VP.n23 VP.n22 0.189894
R81 VP.n23 VP.n10 0.189894
R82 VP.n28 VP.n10 0.189894
R83 VP.n29 VP.n28 0.189894
R84 VP.n30 VP.n29 0.189894
R85 VP.n30 VP.n8 0.189894
R86 VP.n39 VP.n38 0.189894
R87 VP.n40 VP.n39 0.189894
R88 VP.n40 VP.n6 0.189894
R89 VP.n45 VP.n6 0.189894
R90 VP.n46 VP.n45 0.189894
R91 VP.n47 VP.n46 0.189894
R92 VP.n47 VP.n4 0.189894
R93 VP.n51 VP.n4 0.189894
R94 VP.n52 VP.n51 0.189894
R95 VP.n53 VP.n52 0.189894
R96 VP.n53 VP.n2 0.189894
R97 VP.n58 VP.n2 0.189894
R98 VP.n59 VP.n58 0.189894
R99 VP.n60 VP.n59 0.189894
R100 VP.n60 VP.n0 0.189894
R101 VP VP.n64 0.153454
R102 VDD1 VDD1.n0 65.6759
R103 VDD1.n3 VDD1.n2 65.5622
R104 VDD1.n3 VDD1.n1 65.5622
R105 VDD1.n5 VDD1.n4 64.4624
R106 VDD1.n5 VDD1.n3 48.7207
R107 VDD1.n4 VDD1.t4 1.21746
R108 VDD1.n4 VDD1.t2 1.21746
R109 VDD1.n0 VDD1.t6 1.21746
R110 VDD1.n0 VDD1.t7 1.21746
R111 VDD1.n2 VDD1.t0 1.21746
R112 VDD1.n2 VDD1.t1 1.21746
R113 VDD1.n1 VDD1.t3 1.21746
R114 VDD1.n1 VDD1.t5 1.21746
R115 VDD1 VDD1.n5 1.09748
R116 VTAIL.n722 VTAIL.n638 289.615
R117 VTAIL.n86 VTAIL.n2 289.615
R118 VTAIL.n176 VTAIL.n92 289.615
R119 VTAIL.n268 VTAIL.n184 289.615
R120 VTAIL.n632 VTAIL.n548 289.615
R121 VTAIL.n540 VTAIL.n456 289.615
R122 VTAIL.n450 VTAIL.n366 289.615
R123 VTAIL.n358 VTAIL.n274 289.615
R124 VTAIL.n666 VTAIL.n665 185
R125 VTAIL.n671 VTAIL.n670 185
R126 VTAIL.n673 VTAIL.n672 185
R127 VTAIL.n662 VTAIL.n661 185
R128 VTAIL.n679 VTAIL.n678 185
R129 VTAIL.n681 VTAIL.n680 185
R130 VTAIL.n658 VTAIL.n657 185
R131 VTAIL.n687 VTAIL.n686 185
R132 VTAIL.n689 VTAIL.n688 185
R133 VTAIL.n654 VTAIL.n653 185
R134 VTAIL.n695 VTAIL.n694 185
R135 VTAIL.n697 VTAIL.n696 185
R136 VTAIL.n650 VTAIL.n649 185
R137 VTAIL.n703 VTAIL.n702 185
R138 VTAIL.n705 VTAIL.n704 185
R139 VTAIL.n646 VTAIL.n645 185
R140 VTAIL.n712 VTAIL.n711 185
R141 VTAIL.n713 VTAIL.n644 185
R142 VTAIL.n715 VTAIL.n714 185
R143 VTAIL.n642 VTAIL.n641 185
R144 VTAIL.n721 VTAIL.n720 185
R145 VTAIL.n723 VTAIL.n722 185
R146 VTAIL.n30 VTAIL.n29 185
R147 VTAIL.n35 VTAIL.n34 185
R148 VTAIL.n37 VTAIL.n36 185
R149 VTAIL.n26 VTAIL.n25 185
R150 VTAIL.n43 VTAIL.n42 185
R151 VTAIL.n45 VTAIL.n44 185
R152 VTAIL.n22 VTAIL.n21 185
R153 VTAIL.n51 VTAIL.n50 185
R154 VTAIL.n53 VTAIL.n52 185
R155 VTAIL.n18 VTAIL.n17 185
R156 VTAIL.n59 VTAIL.n58 185
R157 VTAIL.n61 VTAIL.n60 185
R158 VTAIL.n14 VTAIL.n13 185
R159 VTAIL.n67 VTAIL.n66 185
R160 VTAIL.n69 VTAIL.n68 185
R161 VTAIL.n10 VTAIL.n9 185
R162 VTAIL.n76 VTAIL.n75 185
R163 VTAIL.n77 VTAIL.n8 185
R164 VTAIL.n79 VTAIL.n78 185
R165 VTAIL.n6 VTAIL.n5 185
R166 VTAIL.n85 VTAIL.n84 185
R167 VTAIL.n87 VTAIL.n86 185
R168 VTAIL.n120 VTAIL.n119 185
R169 VTAIL.n125 VTAIL.n124 185
R170 VTAIL.n127 VTAIL.n126 185
R171 VTAIL.n116 VTAIL.n115 185
R172 VTAIL.n133 VTAIL.n132 185
R173 VTAIL.n135 VTAIL.n134 185
R174 VTAIL.n112 VTAIL.n111 185
R175 VTAIL.n141 VTAIL.n140 185
R176 VTAIL.n143 VTAIL.n142 185
R177 VTAIL.n108 VTAIL.n107 185
R178 VTAIL.n149 VTAIL.n148 185
R179 VTAIL.n151 VTAIL.n150 185
R180 VTAIL.n104 VTAIL.n103 185
R181 VTAIL.n157 VTAIL.n156 185
R182 VTAIL.n159 VTAIL.n158 185
R183 VTAIL.n100 VTAIL.n99 185
R184 VTAIL.n166 VTAIL.n165 185
R185 VTAIL.n167 VTAIL.n98 185
R186 VTAIL.n169 VTAIL.n168 185
R187 VTAIL.n96 VTAIL.n95 185
R188 VTAIL.n175 VTAIL.n174 185
R189 VTAIL.n177 VTAIL.n176 185
R190 VTAIL.n212 VTAIL.n211 185
R191 VTAIL.n217 VTAIL.n216 185
R192 VTAIL.n219 VTAIL.n218 185
R193 VTAIL.n208 VTAIL.n207 185
R194 VTAIL.n225 VTAIL.n224 185
R195 VTAIL.n227 VTAIL.n226 185
R196 VTAIL.n204 VTAIL.n203 185
R197 VTAIL.n233 VTAIL.n232 185
R198 VTAIL.n235 VTAIL.n234 185
R199 VTAIL.n200 VTAIL.n199 185
R200 VTAIL.n241 VTAIL.n240 185
R201 VTAIL.n243 VTAIL.n242 185
R202 VTAIL.n196 VTAIL.n195 185
R203 VTAIL.n249 VTAIL.n248 185
R204 VTAIL.n251 VTAIL.n250 185
R205 VTAIL.n192 VTAIL.n191 185
R206 VTAIL.n258 VTAIL.n257 185
R207 VTAIL.n259 VTAIL.n190 185
R208 VTAIL.n261 VTAIL.n260 185
R209 VTAIL.n188 VTAIL.n187 185
R210 VTAIL.n267 VTAIL.n266 185
R211 VTAIL.n269 VTAIL.n268 185
R212 VTAIL.n633 VTAIL.n632 185
R213 VTAIL.n631 VTAIL.n630 185
R214 VTAIL.n552 VTAIL.n551 185
R215 VTAIL.n625 VTAIL.n624 185
R216 VTAIL.n623 VTAIL.n554 185
R217 VTAIL.n622 VTAIL.n621 185
R218 VTAIL.n557 VTAIL.n555 185
R219 VTAIL.n616 VTAIL.n615 185
R220 VTAIL.n614 VTAIL.n613 185
R221 VTAIL.n561 VTAIL.n560 185
R222 VTAIL.n608 VTAIL.n607 185
R223 VTAIL.n606 VTAIL.n605 185
R224 VTAIL.n565 VTAIL.n564 185
R225 VTAIL.n600 VTAIL.n599 185
R226 VTAIL.n598 VTAIL.n597 185
R227 VTAIL.n569 VTAIL.n568 185
R228 VTAIL.n592 VTAIL.n591 185
R229 VTAIL.n590 VTAIL.n589 185
R230 VTAIL.n573 VTAIL.n572 185
R231 VTAIL.n584 VTAIL.n583 185
R232 VTAIL.n582 VTAIL.n581 185
R233 VTAIL.n577 VTAIL.n576 185
R234 VTAIL.n541 VTAIL.n540 185
R235 VTAIL.n539 VTAIL.n538 185
R236 VTAIL.n460 VTAIL.n459 185
R237 VTAIL.n533 VTAIL.n532 185
R238 VTAIL.n531 VTAIL.n462 185
R239 VTAIL.n530 VTAIL.n529 185
R240 VTAIL.n465 VTAIL.n463 185
R241 VTAIL.n524 VTAIL.n523 185
R242 VTAIL.n522 VTAIL.n521 185
R243 VTAIL.n469 VTAIL.n468 185
R244 VTAIL.n516 VTAIL.n515 185
R245 VTAIL.n514 VTAIL.n513 185
R246 VTAIL.n473 VTAIL.n472 185
R247 VTAIL.n508 VTAIL.n507 185
R248 VTAIL.n506 VTAIL.n505 185
R249 VTAIL.n477 VTAIL.n476 185
R250 VTAIL.n500 VTAIL.n499 185
R251 VTAIL.n498 VTAIL.n497 185
R252 VTAIL.n481 VTAIL.n480 185
R253 VTAIL.n492 VTAIL.n491 185
R254 VTAIL.n490 VTAIL.n489 185
R255 VTAIL.n485 VTAIL.n484 185
R256 VTAIL.n451 VTAIL.n450 185
R257 VTAIL.n449 VTAIL.n448 185
R258 VTAIL.n370 VTAIL.n369 185
R259 VTAIL.n443 VTAIL.n442 185
R260 VTAIL.n441 VTAIL.n372 185
R261 VTAIL.n440 VTAIL.n439 185
R262 VTAIL.n375 VTAIL.n373 185
R263 VTAIL.n434 VTAIL.n433 185
R264 VTAIL.n432 VTAIL.n431 185
R265 VTAIL.n379 VTAIL.n378 185
R266 VTAIL.n426 VTAIL.n425 185
R267 VTAIL.n424 VTAIL.n423 185
R268 VTAIL.n383 VTAIL.n382 185
R269 VTAIL.n418 VTAIL.n417 185
R270 VTAIL.n416 VTAIL.n415 185
R271 VTAIL.n387 VTAIL.n386 185
R272 VTAIL.n410 VTAIL.n409 185
R273 VTAIL.n408 VTAIL.n407 185
R274 VTAIL.n391 VTAIL.n390 185
R275 VTAIL.n402 VTAIL.n401 185
R276 VTAIL.n400 VTAIL.n399 185
R277 VTAIL.n395 VTAIL.n394 185
R278 VTAIL.n359 VTAIL.n358 185
R279 VTAIL.n357 VTAIL.n356 185
R280 VTAIL.n278 VTAIL.n277 185
R281 VTAIL.n351 VTAIL.n350 185
R282 VTAIL.n349 VTAIL.n280 185
R283 VTAIL.n348 VTAIL.n347 185
R284 VTAIL.n283 VTAIL.n281 185
R285 VTAIL.n342 VTAIL.n341 185
R286 VTAIL.n340 VTAIL.n339 185
R287 VTAIL.n287 VTAIL.n286 185
R288 VTAIL.n334 VTAIL.n333 185
R289 VTAIL.n332 VTAIL.n331 185
R290 VTAIL.n291 VTAIL.n290 185
R291 VTAIL.n326 VTAIL.n325 185
R292 VTAIL.n324 VTAIL.n323 185
R293 VTAIL.n295 VTAIL.n294 185
R294 VTAIL.n318 VTAIL.n317 185
R295 VTAIL.n316 VTAIL.n315 185
R296 VTAIL.n299 VTAIL.n298 185
R297 VTAIL.n310 VTAIL.n309 185
R298 VTAIL.n308 VTAIL.n307 185
R299 VTAIL.n303 VTAIL.n302 185
R300 VTAIL.n667 VTAIL.t3 147.659
R301 VTAIL.n31 VTAIL.t1 147.659
R302 VTAIL.n121 VTAIL.t11 147.659
R303 VTAIL.n213 VTAIL.t15 147.659
R304 VTAIL.n578 VTAIL.t14 147.659
R305 VTAIL.n486 VTAIL.t8 147.659
R306 VTAIL.n396 VTAIL.t0 147.659
R307 VTAIL.n304 VTAIL.t6 147.659
R308 VTAIL.n671 VTAIL.n665 104.615
R309 VTAIL.n672 VTAIL.n671 104.615
R310 VTAIL.n672 VTAIL.n661 104.615
R311 VTAIL.n679 VTAIL.n661 104.615
R312 VTAIL.n680 VTAIL.n679 104.615
R313 VTAIL.n680 VTAIL.n657 104.615
R314 VTAIL.n687 VTAIL.n657 104.615
R315 VTAIL.n688 VTAIL.n687 104.615
R316 VTAIL.n688 VTAIL.n653 104.615
R317 VTAIL.n695 VTAIL.n653 104.615
R318 VTAIL.n696 VTAIL.n695 104.615
R319 VTAIL.n696 VTAIL.n649 104.615
R320 VTAIL.n703 VTAIL.n649 104.615
R321 VTAIL.n704 VTAIL.n703 104.615
R322 VTAIL.n704 VTAIL.n645 104.615
R323 VTAIL.n712 VTAIL.n645 104.615
R324 VTAIL.n713 VTAIL.n712 104.615
R325 VTAIL.n714 VTAIL.n713 104.615
R326 VTAIL.n714 VTAIL.n641 104.615
R327 VTAIL.n721 VTAIL.n641 104.615
R328 VTAIL.n722 VTAIL.n721 104.615
R329 VTAIL.n35 VTAIL.n29 104.615
R330 VTAIL.n36 VTAIL.n35 104.615
R331 VTAIL.n36 VTAIL.n25 104.615
R332 VTAIL.n43 VTAIL.n25 104.615
R333 VTAIL.n44 VTAIL.n43 104.615
R334 VTAIL.n44 VTAIL.n21 104.615
R335 VTAIL.n51 VTAIL.n21 104.615
R336 VTAIL.n52 VTAIL.n51 104.615
R337 VTAIL.n52 VTAIL.n17 104.615
R338 VTAIL.n59 VTAIL.n17 104.615
R339 VTAIL.n60 VTAIL.n59 104.615
R340 VTAIL.n60 VTAIL.n13 104.615
R341 VTAIL.n67 VTAIL.n13 104.615
R342 VTAIL.n68 VTAIL.n67 104.615
R343 VTAIL.n68 VTAIL.n9 104.615
R344 VTAIL.n76 VTAIL.n9 104.615
R345 VTAIL.n77 VTAIL.n76 104.615
R346 VTAIL.n78 VTAIL.n77 104.615
R347 VTAIL.n78 VTAIL.n5 104.615
R348 VTAIL.n85 VTAIL.n5 104.615
R349 VTAIL.n86 VTAIL.n85 104.615
R350 VTAIL.n125 VTAIL.n119 104.615
R351 VTAIL.n126 VTAIL.n125 104.615
R352 VTAIL.n126 VTAIL.n115 104.615
R353 VTAIL.n133 VTAIL.n115 104.615
R354 VTAIL.n134 VTAIL.n133 104.615
R355 VTAIL.n134 VTAIL.n111 104.615
R356 VTAIL.n141 VTAIL.n111 104.615
R357 VTAIL.n142 VTAIL.n141 104.615
R358 VTAIL.n142 VTAIL.n107 104.615
R359 VTAIL.n149 VTAIL.n107 104.615
R360 VTAIL.n150 VTAIL.n149 104.615
R361 VTAIL.n150 VTAIL.n103 104.615
R362 VTAIL.n157 VTAIL.n103 104.615
R363 VTAIL.n158 VTAIL.n157 104.615
R364 VTAIL.n158 VTAIL.n99 104.615
R365 VTAIL.n166 VTAIL.n99 104.615
R366 VTAIL.n167 VTAIL.n166 104.615
R367 VTAIL.n168 VTAIL.n167 104.615
R368 VTAIL.n168 VTAIL.n95 104.615
R369 VTAIL.n175 VTAIL.n95 104.615
R370 VTAIL.n176 VTAIL.n175 104.615
R371 VTAIL.n217 VTAIL.n211 104.615
R372 VTAIL.n218 VTAIL.n217 104.615
R373 VTAIL.n218 VTAIL.n207 104.615
R374 VTAIL.n225 VTAIL.n207 104.615
R375 VTAIL.n226 VTAIL.n225 104.615
R376 VTAIL.n226 VTAIL.n203 104.615
R377 VTAIL.n233 VTAIL.n203 104.615
R378 VTAIL.n234 VTAIL.n233 104.615
R379 VTAIL.n234 VTAIL.n199 104.615
R380 VTAIL.n241 VTAIL.n199 104.615
R381 VTAIL.n242 VTAIL.n241 104.615
R382 VTAIL.n242 VTAIL.n195 104.615
R383 VTAIL.n249 VTAIL.n195 104.615
R384 VTAIL.n250 VTAIL.n249 104.615
R385 VTAIL.n250 VTAIL.n191 104.615
R386 VTAIL.n258 VTAIL.n191 104.615
R387 VTAIL.n259 VTAIL.n258 104.615
R388 VTAIL.n260 VTAIL.n259 104.615
R389 VTAIL.n260 VTAIL.n187 104.615
R390 VTAIL.n267 VTAIL.n187 104.615
R391 VTAIL.n268 VTAIL.n267 104.615
R392 VTAIL.n632 VTAIL.n631 104.615
R393 VTAIL.n631 VTAIL.n551 104.615
R394 VTAIL.n624 VTAIL.n551 104.615
R395 VTAIL.n624 VTAIL.n623 104.615
R396 VTAIL.n623 VTAIL.n622 104.615
R397 VTAIL.n622 VTAIL.n555 104.615
R398 VTAIL.n615 VTAIL.n555 104.615
R399 VTAIL.n615 VTAIL.n614 104.615
R400 VTAIL.n614 VTAIL.n560 104.615
R401 VTAIL.n607 VTAIL.n560 104.615
R402 VTAIL.n607 VTAIL.n606 104.615
R403 VTAIL.n606 VTAIL.n564 104.615
R404 VTAIL.n599 VTAIL.n564 104.615
R405 VTAIL.n599 VTAIL.n598 104.615
R406 VTAIL.n598 VTAIL.n568 104.615
R407 VTAIL.n591 VTAIL.n568 104.615
R408 VTAIL.n591 VTAIL.n590 104.615
R409 VTAIL.n590 VTAIL.n572 104.615
R410 VTAIL.n583 VTAIL.n572 104.615
R411 VTAIL.n583 VTAIL.n582 104.615
R412 VTAIL.n582 VTAIL.n576 104.615
R413 VTAIL.n540 VTAIL.n539 104.615
R414 VTAIL.n539 VTAIL.n459 104.615
R415 VTAIL.n532 VTAIL.n459 104.615
R416 VTAIL.n532 VTAIL.n531 104.615
R417 VTAIL.n531 VTAIL.n530 104.615
R418 VTAIL.n530 VTAIL.n463 104.615
R419 VTAIL.n523 VTAIL.n463 104.615
R420 VTAIL.n523 VTAIL.n522 104.615
R421 VTAIL.n522 VTAIL.n468 104.615
R422 VTAIL.n515 VTAIL.n468 104.615
R423 VTAIL.n515 VTAIL.n514 104.615
R424 VTAIL.n514 VTAIL.n472 104.615
R425 VTAIL.n507 VTAIL.n472 104.615
R426 VTAIL.n507 VTAIL.n506 104.615
R427 VTAIL.n506 VTAIL.n476 104.615
R428 VTAIL.n499 VTAIL.n476 104.615
R429 VTAIL.n499 VTAIL.n498 104.615
R430 VTAIL.n498 VTAIL.n480 104.615
R431 VTAIL.n491 VTAIL.n480 104.615
R432 VTAIL.n491 VTAIL.n490 104.615
R433 VTAIL.n490 VTAIL.n484 104.615
R434 VTAIL.n450 VTAIL.n449 104.615
R435 VTAIL.n449 VTAIL.n369 104.615
R436 VTAIL.n442 VTAIL.n369 104.615
R437 VTAIL.n442 VTAIL.n441 104.615
R438 VTAIL.n441 VTAIL.n440 104.615
R439 VTAIL.n440 VTAIL.n373 104.615
R440 VTAIL.n433 VTAIL.n373 104.615
R441 VTAIL.n433 VTAIL.n432 104.615
R442 VTAIL.n432 VTAIL.n378 104.615
R443 VTAIL.n425 VTAIL.n378 104.615
R444 VTAIL.n425 VTAIL.n424 104.615
R445 VTAIL.n424 VTAIL.n382 104.615
R446 VTAIL.n417 VTAIL.n382 104.615
R447 VTAIL.n417 VTAIL.n416 104.615
R448 VTAIL.n416 VTAIL.n386 104.615
R449 VTAIL.n409 VTAIL.n386 104.615
R450 VTAIL.n409 VTAIL.n408 104.615
R451 VTAIL.n408 VTAIL.n390 104.615
R452 VTAIL.n401 VTAIL.n390 104.615
R453 VTAIL.n401 VTAIL.n400 104.615
R454 VTAIL.n400 VTAIL.n394 104.615
R455 VTAIL.n358 VTAIL.n357 104.615
R456 VTAIL.n357 VTAIL.n277 104.615
R457 VTAIL.n350 VTAIL.n277 104.615
R458 VTAIL.n350 VTAIL.n349 104.615
R459 VTAIL.n349 VTAIL.n348 104.615
R460 VTAIL.n348 VTAIL.n281 104.615
R461 VTAIL.n341 VTAIL.n281 104.615
R462 VTAIL.n341 VTAIL.n340 104.615
R463 VTAIL.n340 VTAIL.n286 104.615
R464 VTAIL.n333 VTAIL.n286 104.615
R465 VTAIL.n333 VTAIL.n332 104.615
R466 VTAIL.n332 VTAIL.n290 104.615
R467 VTAIL.n325 VTAIL.n290 104.615
R468 VTAIL.n325 VTAIL.n324 104.615
R469 VTAIL.n324 VTAIL.n294 104.615
R470 VTAIL.n317 VTAIL.n294 104.615
R471 VTAIL.n317 VTAIL.n316 104.615
R472 VTAIL.n316 VTAIL.n298 104.615
R473 VTAIL.n309 VTAIL.n298 104.615
R474 VTAIL.n309 VTAIL.n308 104.615
R475 VTAIL.n308 VTAIL.n302 104.615
R476 VTAIL.t3 VTAIL.n665 52.3082
R477 VTAIL.t1 VTAIL.n29 52.3082
R478 VTAIL.t11 VTAIL.n119 52.3082
R479 VTAIL.t15 VTAIL.n211 52.3082
R480 VTAIL.t14 VTAIL.n576 52.3082
R481 VTAIL.t8 VTAIL.n484 52.3082
R482 VTAIL.t0 VTAIL.n394 52.3082
R483 VTAIL.t6 VTAIL.n302 52.3082
R484 VTAIL.n547 VTAIL.n546 47.7838
R485 VTAIL.n365 VTAIL.n364 47.7838
R486 VTAIL.n1 VTAIL.n0 47.7836
R487 VTAIL.n183 VTAIL.n182 47.7836
R488 VTAIL.n727 VTAIL.n726 35.8702
R489 VTAIL.n91 VTAIL.n90 35.8702
R490 VTAIL.n181 VTAIL.n180 35.8702
R491 VTAIL.n273 VTAIL.n272 35.8702
R492 VTAIL.n637 VTAIL.n636 35.8702
R493 VTAIL.n545 VTAIL.n544 35.8702
R494 VTAIL.n455 VTAIL.n454 35.8702
R495 VTAIL.n363 VTAIL.n362 35.8702
R496 VTAIL.n727 VTAIL.n637 28.7031
R497 VTAIL.n363 VTAIL.n273 28.7031
R498 VTAIL.n667 VTAIL.n666 15.6677
R499 VTAIL.n31 VTAIL.n30 15.6677
R500 VTAIL.n121 VTAIL.n120 15.6677
R501 VTAIL.n213 VTAIL.n212 15.6677
R502 VTAIL.n578 VTAIL.n577 15.6677
R503 VTAIL.n486 VTAIL.n485 15.6677
R504 VTAIL.n396 VTAIL.n395 15.6677
R505 VTAIL.n304 VTAIL.n303 15.6677
R506 VTAIL.n715 VTAIL.n644 13.1884
R507 VTAIL.n79 VTAIL.n8 13.1884
R508 VTAIL.n169 VTAIL.n98 13.1884
R509 VTAIL.n261 VTAIL.n190 13.1884
R510 VTAIL.n625 VTAIL.n554 13.1884
R511 VTAIL.n533 VTAIL.n462 13.1884
R512 VTAIL.n443 VTAIL.n372 13.1884
R513 VTAIL.n351 VTAIL.n280 13.1884
R514 VTAIL.n670 VTAIL.n669 12.8005
R515 VTAIL.n711 VTAIL.n710 12.8005
R516 VTAIL.n716 VTAIL.n642 12.8005
R517 VTAIL.n34 VTAIL.n33 12.8005
R518 VTAIL.n75 VTAIL.n74 12.8005
R519 VTAIL.n80 VTAIL.n6 12.8005
R520 VTAIL.n124 VTAIL.n123 12.8005
R521 VTAIL.n165 VTAIL.n164 12.8005
R522 VTAIL.n170 VTAIL.n96 12.8005
R523 VTAIL.n216 VTAIL.n215 12.8005
R524 VTAIL.n257 VTAIL.n256 12.8005
R525 VTAIL.n262 VTAIL.n188 12.8005
R526 VTAIL.n626 VTAIL.n552 12.8005
R527 VTAIL.n621 VTAIL.n556 12.8005
R528 VTAIL.n581 VTAIL.n580 12.8005
R529 VTAIL.n534 VTAIL.n460 12.8005
R530 VTAIL.n529 VTAIL.n464 12.8005
R531 VTAIL.n489 VTAIL.n488 12.8005
R532 VTAIL.n444 VTAIL.n370 12.8005
R533 VTAIL.n439 VTAIL.n374 12.8005
R534 VTAIL.n399 VTAIL.n398 12.8005
R535 VTAIL.n352 VTAIL.n278 12.8005
R536 VTAIL.n347 VTAIL.n282 12.8005
R537 VTAIL.n307 VTAIL.n306 12.8005
R538 VTAIL.n673 VTAIL.n664 12.0247
R539 VTAIL.n709 VTAIL.n646 12.0247
R540 VTAIL.n720 VTAIL.n719 12.0247
R541 VTAIL.n37 VTAIL.n28 12.0247
R542 VTAIL.n73 VTAIL.n10 12.0247
R543 VTAIL.n84 VTAIL.n83 12.0247
R544 VTAIL.n127 VTAIL.n118 12.0247
R545 VTAIL.n163 VTAIL.n100 12.0247
R546 VTAIL.n174 VTAIL.n173 12.0247
R547 VTAIL.n219 VTAIL.n210 12.0247
R548 VTAIL.n255 VTAIL.n192 12.0247
R549 VTAIL.n266 VTAIL.n265 12.0247
R550 VTAIL.n630 VTAIL.n629 12.0247
R551 VTAIL.n620 VTAIL.n557 12.0247
R552 VTAIL.n584 VTAIL.n575 12.0247
R553 VTAIL.n538 VTAIL.n537 12.0247
R554 VTAIL.n528 VTAIL.n465 12.0247
R555 VTAIL.n492 VTAIL.n483 12.0247
R556 VTAIL.n448 VTAIL.n447 12.0247
R557 VTAIL.n438 VTAIL.n375 12.0247
R558 VTAIL.n402 VTAIL.n393 12.0247
R559 VTAIL.n356 VTAIL.n355 12.0247
R560 VTAIL.n346 VTAIL.n283 12.0247
R561 VTAIL.n310 VTAIL.n301 12.0247
R562 VTAIL.n674 VTAIL.n662 11.249
R563 VTAIL.n706 VTAIL.n705 11.249
R564 VTAIL.n723 VTAIL.n640 11.249
R565 VTAIL.n38 VTAIL.n26 11.249
R566 VTAIL.n70 VTAIL.n69 11.249
R567 VTAIL.n87 VTAIL.n4 11.249
R568 VTAIL.n128 VTAIL.n116 11.249
R569 VTAIL.n160 VTAIL.n159 11.249
R570 VTAIL.n177 VTAIL.n94 11.249
R571 VTAIL.n220 VTAIL.n208 11.249
R572 VTAIL.n252 VTAIL.n251 11.249
R573 VTAIL.n269 VTAIL.n186 11.249
R574 VTAIL.n633 VTAIL.n550 11.249
R575 VTAIL.n617 VTAIL.n616 11.249
R576 VTAIL.n585 VTAIL.n573 11.249
R577 VTAIL.n541 VTAIL.n458 11.249
R578 VTAIL.n525 VTAIL.n524 11.249
R579 VTAIL.n493 VTAIL.n481 11.249
R580 VTAIL.n451 VTAIL.n368 11.249
R581 VTAIL.n435 VTAIL.n434 11.249
R582 VTAIL.n403 VTAIL.n391 11.249
R583 VTAIL.n359 VTAIL.n276 11.249
R584 VTAIL.n343 VTAIL.n342 11.249
R585 VTAIL.n311 VTAIL.n299 11.249
R586 VTAIL.n678 VTAIL.n677 10.4732
R587 VTAIL.n702 VTAIL.n648 10.4732
R588 VTAIL.n724 VTAIL.n638 10.4732
R589 VTAIL.n42 VTAIL.n41 10.4732
R590 VTAIL.n66 VTAIL.n12 10.4732
R591 VTAIL.n88 VTAIL.n2 10.4732
R592 VTAIL.n132 VTAIL.n131 10.4732
R593 VTAIL.n156 VTAIL.n102 10.4732
R594 VTAIL.n178 VTAIL.n92 10.4732
R595 VTAIL.n224 VTAIL.n223 10.4732
R596 VTAIL.n248 VTAIL.n194 10.4732
R597 VTAIL.n270 VTAIL.n184 10.4732
R598 VTAIL.n634 VTAIL.n548 10.4732
R599 VTAIL.n613 VTAIL.n559 10.4732
R600 VTAIL.n589 VTAIL.n588 10.4732
R601 VTAIL.n542 VTAIL.n456 10.4732
R602 VTAIL.n521 VTAIL.n467 10.4732
R603 VTAIL.n497 VTAIL.n496 10.4732
R604 VTAIL.n452 VTAIL.n366 10.4732
R605 VTAIL.n431 VTAIL.n377 10.4732
R606 VTAIL.n407 VTAIL.n406 10.4732
R607 VTAIL.n360 VTAIL.n274 10.4732
R608 VTAIL.n339 VTAIL.n285 10.4732
R609 VTAIL.n315 VTAIL.n314 10.4732
R610 VTAIL.n681 VTAIL.n660 9.69747
R611 VTAIL.n701 VTAIL.n650 9.69747
R612 VTAIL.n45 VTAIL.n24 9.69747
R613 VTAIL.n65 VTAIL.n14 9.69747
R614 VTAIL.n135 VTAIL.n114 9.69747
R615 VTAIL.n155 VTAIL.n104 9.69747
R616 VTAIL.n227 VTAIL.n206 9.69747
R617 VTAIL.n247 VTAIL.n196 9.69747
R618 VTAIL.n612 VTAIL.n561 9.69747
R619 VTAIL.n592 VTAIL.n571 9.69747
R620 VTAIL.n520 VTAIL.n469 9.69747
R621 VTAIL.n500 VTAIL.n479 9.69747
R622 VTAIL.n430 VTAIL.n379 9.69747
R623 VTAIL.n410 VTAIL.n389 9.69747
R624 VTAIL.n338 VTAIL.n287 9.69747
R625 VTAIL.n318 VTAIL.n297 9.69747
R626 VTAIL.n726 VTAIL.n725 9.45567
R627 VTAIL.n90 VTAIL.n89 9.45567
R628 VTAIL.n180 VTAIL.n179 9.45567
R629 VTAIL.n272 VTAIL.n271 9.45567
R630 VTAIL.n636 VTAIL.n635 9.45567
R631 VTAIL.n544 VTAIL.n543 9.45567
R632 VTAIL.n454 VTAIL.n453 9.45567
R633 VTAIL.n362 VTAIL.n361 9.45567
R634 VTAIL.n725 VTAIL.n724 9.3005
R635 VTAIL.n640 VTAIL.n639 9.3005
R636 VTAIL.n719 VTAIL.n718 9.3005
R637 VTAIL.n717 VTAIL.n716 9.3005
R638 VTAIL.n656 VTAIL.n655 9.3005
R639 VTAIL.n685 VTAIL.n684 9.3005
R640 VTAIL.n683 VTAIL.n682 9.3005
R641 VTAIL.n660 VTAIL.n659 9.3005
R642 VTAIL.n677 VTAIL.n676 9.3005
R643 VTAIL.n675 VTAIL.n674 9.3005
R644 VTAIL.n664 VTAIL.n663 9.3005
R645 VTAIL.n669 VTAIL.n668 9.3005
R646 VTAIL.n691 VTAIL.n690 9.3005
R647 VTAIL.n693 VTAIL.n692 9.3005
R648 VTAIL.n652 VTAIL.n651 9.3005
R649 VTAIL.n699 VTAIL.n698 9.3005
R650 VTAIL.n701 VTAIL.n700 9.3005
R651 VTAIL.n648 VTAIL.n647 9.3005
R652 VTAIL.n707 VTAIL.n706 9.3005
R653 VTAIL.n709 VTAIL.n708 9.3005
R654 VTAIL.n710 VTAIL.n643 9.3005
R655 VTAIL.n89 VTAIL.n88 9.3005
R656 VTAIL.n4 VTAIL.n3 9.3005
R657 VTAIL.n83 VTAIL.n82 9.3005
R658 VTAIL.n81 VTAIL.n80 9.3005
R659 VTAIL.n20 VTAIL.n19 9.3005
R660 VTAIL.n49 VTAIL.n48 9.3005
R661 VTAIL.n47 VTAIL.n46 9.3005
R662 VTAIL.n24 VTAIL.n23 9.3005
R663 VTAIL.n41 VTAIL.n40 9.3005
R664 VTAIL.n39 VTAIL.n38 9.3005
R665 VTAIL.n28 VTAIL.n27 9.3005
R666 VTAIL.n33 VTAIL.n32 9.3005
R667 VTAIL.n55 VTAIL.n54 9.3005
R668 VTAIL.n57 VTAIL.n56 9.3005
R669 VTAIL.n16 VTAIL.n15 9.3005
R670 VTAIL.n63 VTAIL.n62 9.3005
R671 VTAIL.n65 VTAIL.n64 9.3005
R672 VTAIL.n12 VTAIL.n11 9.3005
R673 VTAIL.n71 VTAIL.n70 9.3005
R674 VTAIL.n73 VTAIL.n72 9.3005
R675 VTAIL.n74 VTAIL.n7 9.3005
R676 VTAIL.n179 VTAIL.n178 9.3005
R677 VTAIL.n94 VTAIL.n93 9.3005
R678 VTAIL.n173 VTAIL.n172 9.3005
R679 VTAIL.n171 VTAIL.n170 9.3005
R680 VTAIL.n110 VTAIL.n109 9.3005
R681 VTAIL.n139 VTAIL.n138 9.3005
R682 VTAIL.n137 VTAIL.n136 9.3005
R683 VTAIL.n114 VTAIL.n113 9.3005
R684 VTAIL.n131 VTAIL.n130 9.3005
R685 VTAIL.n129 VTAIL.n128 9.3005
R686 VTAIL.n118 VTAIL.n117 9.3005
R687 VTAIL.n123 VTAIL.n122 9.3005
R688 VTAIL.n145 VTAIL.n144 9.3005
R689 VTAIL.n147 VTAIL.n146 9.3005
R690 VTAIL.n106 VTAIL.n105 9.3005
R691 VTAIL.n153 VTAIL.n152 9.3005
R692 VTAIL.n155 VTAIL.n154 9.3005
R693 VTAIL.n102 VTAIL.n101 9.3005
R694 VTAIL.n161 VTAIL.n160 9.3005
R695 VTAIL.n163 VTAIL.n162 9.3005
R696 VTAIL.n164 VTAIL.n97 9.3005
R697 VTAIL.n271 VTAIL.n270 9.3005
R698 VTAIL.n186 VTAIL.n185 9.3005
R699 VTAIL.n265 VTAIL.n264 9.3005
R700 VTAIL.n263 VTAIL.n262 9.3005
R701 VTAIL.n202 VTAIL.n201 9.3005
R702 VTAIL.n231 VTAIL.n230 9.3005
R703 VTAIL.n229 VTAIL.n228 9.3005
R704 VTAIL.n206 VTAIL.n205 9.3005
R705 VTAIL.n223 VTAIL.n222 9.3005
R706 VTAIL.n221 VTAIL.n220 9.3005
R707 VTAIL.n210 VTAIL.n209 9.3005
R708 VTAIL.n215 VTAIL.n214 9.3005
R709 VTAIL.n237 VTAIL.n236 9.3005
R710 VTAIL.n239 VTAIL.n238 9.3005
R711 VTAIL.n198 VTAIL.n197 9.3005
R712 VTAIL.n245 VTAIL.n244 9.3005
R713 VTAIL.n247 VTAIL.n246 9.3005
R714 VTAIL.n194 VTAIL.n193 9.3005
R715 VTAIL.n253 VTAIL.n252 9.3005
R716 VTAIL.n255 VTAIL.n254 9.3005
R717 VTAIL.n256 VTAIL.n189 9.3005
R718 VTAIL.n604 VTAIL.n603 9.3005
R719 VTAIL.n563 VTAIL.n562 9.3005
R720 VTAIL.n610 VTAIL.n609 9.3005
R721 VTAIL.n612 VTAIL.n611 9.3005
R722 VTAIL.n559 VTAIL.n558 9.3005
R723 VTAIL.n618 VTAIL.n617 9.3005
R724 VTAIL.n620 VTAIL.n619 9.3005
R725 VTAIL.n556 VTAIL.n553 9.3005
R726 VTAIL.n635 VTAIL.n634 9.3005
R727 VTAIL.n550 VTAIL.n549 9.3005
R728 VTAIL.n629 VTAIL.n628 9.3005
R729 VTAIL.n627 VTAIL.n626 9.3005
R730 VTAIL.n602 VTAIL.n601 9.3005
R731 VTAIL.n567 VTAIL.n566 9.3005
R732 VTAIL.n596 VTAIL.n595 9.3005
R733 VTAIL.n594 VTAIL.n593 9.3005
R734 VTAIL.n571 VTAIL.n570 9.3005
R735 VTAIL.n588 VTAIL.n587 9.3005
R736 VTAIL.n586 VTAIL.n585 9.3005
R737 VTAIL.n575 VTAIL.n574 9.3005
R738 VTAIL.n580 VTAIL.n579 9.3005
R739 VTAIL.n512 VTAIL.n511 9.3005
R740 VTAIL.n471 VTAIL.n470 9.3005
R741 VTAIL.n518 VTAIL.n517 9.3005
R742 VTAIL.n520 VTAIL.n519 9.3005
R743 VTAIL.n467 VTAIL.n466 9.3005
R744 VTAIL.n526 VTAIL.n525 9.3005
R745 VTAIL.n528 VTAIL.n527 9.3005
R746 VTAIL.n464 VTAIL.n461 9.3005
R747 VTAIL.n543 VTAIL.n542 9.3005
R748 VTAIL.n458 VTAIL.n457 9.3005
R749 VTAIL.n537 VTAIL.n536 9.3005
R750 VTAIL.n535 VTAIL.n534 9.3005
R751 VTAIL.n510 VTAIL.n509 9.3005
R752 VTAIL.n475 VTAIL.n474 9.3005
R753 VTAIL.n504 VTAIL.n503 9.3005
R754 VTAIL.n502 VTAIL.n501 9.3005
R755 VTAIL.n479 VTAIL.n478 9.3005
R756 VTAIL.n496 VTAIL.n495 9.3005
R757 VTAIL.n494 VTAIL.n493 9.3005
R758 VTAIL.n483 VTAIL.n482 9.3005
R759 VTAIL.n488 VTAIL.n487 9.3005
R760 VTAIL.n422 VTAIL.n421 9.3005
R761 VTAIL.n381 VTAIL.n380 9.3005
R762 VTAIL.n428 VTAIL.n427 9.3005
R763 VTAIL.n430 VTAIL.n429 9.3005
R764 VTAIL.n377 VTAIL.n376 9.3005
R765 VTAIL.n436 VTAIL.n435 9.3005
R766 VTAIL.n438 VTAIL.n437 9.3005
R767 VTAIL.n374 VTAIL.n371 9.3005
R768 VTAIL.n453 VTAIL.n452 9.3005
R769 VTAIL.n368 VTAIL.n367 9.3005
R770 VTAIL.n447 VTAIL.n446 9.3005
R771 VTAIL.n445 VTAIL.n444 9.3005
R772 VTAIL.n420 VTAIL.n419 9.3005
R773 VTAIL.n385 VTAIL.n384 9.3005
R774 VTAIL.n414 VTAIL.n413 9.3005
R775 VTAIL.n412 VTAIL.n411 9.3005
R776 VTAIL.n389 VTAIL.n388 9.3005
R777 VTAIL.n406 VTAIL.n405 9.3005
R778 VTAIL.n404 VTAIL.n403 9.3005
R779 VTAIL.n393 VTAIL.n392 9.3005
R780 VTAIL.n398 VTAIL.n397 9.3005
R781 VTAIL.n330 VTAIL.n329 9.3005
R782 VTAIL.n289 VTAIL.n288 9.3005
R783 VTAIL.n336 VTAIL.n335 9.3005
R784 VTAIL.n338 VTAIL.n337 9.3005
R785 VTAIL.n285 VTAIL.n284 9.3005
R786 VTAIL.n344 VTAIL.n343 9.3005
R787 VTAIL.n346 VTAIL.n345 9.3005
R788 VTAIL.n282 VTAIL.n279 9.3005
R789 VTAIL.n361 VTAIL.n360 9.3005
R790 VTAIL.n276 VTAIL.n275 9.3005
R791 VTAIL.n355 VTAIL.n354 9.3005
R792 VTAIL.n353 VTAIL.n352 9.3005
R793 VTAIL.n328 VTAIL.n327 9.3005
R794 VTAIL.n293 VTAIL.n292 9.3005
R795 VTAIL.n322 VTAIL.n321 9.3005
R796 VTAIL.n320 VTAIL.n319 9.3005
R797 VTAIL.n297 VTAIL.n296 9.3005
R798 VTAIL.n314 VTAIL.n313 9.3005
R799 VTAIL.n312 VTAIL.n311 9.3005
R800 VTAIL.n301 VTAIL.n300 9.3005
R801 VTAIL.n306 VTAIL.n305 9.3005
R802 VTAIL.n682 VTAIL.n658 8.92171
R803 VTAIL.n698 VTAIL.n697 8.92171
R804 VTAIL.n46 VTAIL.n22 8.92171
R805 VTAIL.n62 VTAIL.n61 8.92171
R806 VTAIL.n136 VTAIL.n112 8.92171
R807 VTAIL.n152 VTAIL.n151 8.92171
R808 VTAIL.n228 VTAIL.n204 8.92171
R809 VTAIL.n244 VTAIL.n243 8.92171
R810 VTAIL.n609 VTAIL.n608 8.92171
R811 VTAIL.n593 VTAIL.n569 8.92171
R812 VTAIL.n517 VTAIL.n516 8.92171
R813 VTAIL.n501 VTAIL.n477 8.92171
R814 VTAIL.n427 VTAIL.n426 8.92171
R815 VTAIL.n411 VTAIL.n387 8.92171
R816 VTAIL.n335 VTAIL.n334 8.92171
R817 VTAIL.n319 VTAIL.n295 8.92171
R818 VTAIL.n686 VTAIL.n685 8.14595
R819 VTAIL.n694 VTAIL.n652 8.14595
R820 VTAIL.n50 VTAIL.n49 8.14595
R821 VTAIL.n58 VTAIL.n16 8.14595
R822 VTAIL.n140 VTAIL.n139 8.14595
R823 VTAIL.n148 VTAIL.n106 8.14595
R824 VTAIL.n232 VTAIL.n231 8.14595
R825 VTAIL.n240 VTAIL.n198 8.14595
R826 VTAIL.n605 VTAIL.n563 8.14595
R827 VTAIL.n597 VTAIL.n596 8.14595
R828 VTAIL.n513 VTAIL.n471 8.14595
R829 VTAIL.n505 VTAIL.n504 8.14595
R830 VTAIL.n423 VTAIL.n381 8.14595
R831 VTAIL.n415 VTAIL.n414 8.14595
R832 VTAIL.n331 VTAIL.n289 8.14595
R833 VTAIL.n323 VTAIL.n322 8.14595
R834 VTAIL.n689 VTAIL.n656 7.3702
R835 VTAIL.n693 VTAIL.n654 7.3702
R836 VTAIL.n53 VTAIL.n20 7.3702
R837 VTAIL.n57 VTAIL.n18 7.3702
R838 VTAIL.n143 VTAIL.n110 7.3702
R839 VTAIL.n147 VTAIL.n108 7.3702
R840 VTAIL.n235 VTAIL.n202 7.3702
R841 VTAIL.n239 VTAIL.n200 7.3702
R842 VTAIL.n604 VTAIL.n565 7.3702
R843 VTAIL.n600 VTAIL.n567 7.3702
R844 VTAIL.n512 VTAIL.n473 7.3702
R845 VTAIL.n508 VTAIL.n475 7.3702
R846 VTAIL.n422 VTAIL.n383 7.3702
R847 VTAIL.n418 VTAIL.n385 7.3702
R848 VTAIL.n330 VTAIL.n291 7.3702
R849 VTAIL.n326 VTAIL.n293 7.3702
R850 VTAIL.n690 VTAIL.n689 6.59444
R851 VTAIL.n690 VTAIL.n654 6.59444
R852 VTAIL.n54 VTAIL.n53 6.59444
R853 VTAIL.n54 VTAIL.n18 6.59444
R854 VTAIL.n144 VTAIL.n143 6.59444
R855 VTAIL.n144 VTAIL.n108 6.59444
R856 VTAIL.n236 VTAIL.n235 6.59444
R857 VTAIL.n236 VTAIL.n200 6.59444
R858 VTAIL.n601 VTAIL.n565 6.59444
R859 VTAIL.n601 VTAIL.n600 6.59444
R860 VTAIL.n509 VTAIL.n473 6.59444
R861 VTAIL.n509 VTAIL.n508 6.59444
R862 VTAIL.n419 VTAIL.n383 6.59444
R863 VTAIL.n419 VTAIL.n418 6.59444
R864 VTAIL.n327 VTAIL.n291 6.59444
R865 VTAIL.n327 VTAIL.n326 6.59444
R866 VTAIL.n686 VTAIL.n656 5.81868
R867 VTAIL.n694 VTAIL.n693 5.81868
R868 VTAIL.n50 VTAIL.n20 5.81868
R869 VTAIL.n58 VTAIL.n57 5.81868
R870 VTAIL.n140 VTAIL.n110 5.81868
R871 VTAIL.n148 VTAIL.n147 5.81868
R872 VTAIL.n232 VTAIL.n202 5.81868
R873 VTAIL.n240 VTAIL.n239 5.81868
R874 VTAIL.n605 VTAIL.n604 5.81868
R875 VTAIL.n597 VTAIL.n567 5.81868
R876 VTAIL.n513 VTAIL.n512 5.81868
R877 VTAIL.n505 VTAIL.n475 5.81868
R878 VTAIL.n423 VTAIL.n422 5.81868
R879 VTAIL.n415 VTAIL.n385 5.81868
R880 VTAIL.n331 VTAIL.n330 5.81868
R881 VTAIL.n323 VTAIL.n293 5.81868
R882 VTAIL.n685 VTAIL.n658 5.04292
R883 VTAIL.n697 VTAIL.n652 5.04292
R884 VTAIL.n49 VTAIL.n22 5.04292
R885 VTAIL.n61 VTAIL.n16 5.04292
R886 VTAIL.n139 VTAIL.n112 5.04292
R887 VTAIL.n151 VTAIL.n106 5.04292
R888 VTAIL.n231 VTAIL.n204 5.04292
R889 VTAIL.n243 VTAIL.n198 5.04292
R890 VTAIL.n608 VTAIL.n563 5.04292
R891 VTAIL.n596 VTAIL.n569 5.04292
R892 VTAIL.n516 VTAIL.n471 5.04292
R893 VTAIL.n504 VTAIL.n477 5.04292
R894 VTAIL.n426 VTAIL.n381 5.04292
R895 VTAIL.n414 VTAIL.n387 5.04292
R896 VTAIL.n334 VTAIL.n289 5.04292
R897 VTAIL.n322 VTAIL.n295 5.04292
R898 VTAIL.n668 VTAIL.n667 4.38563
R899 VTAIL.n32 VTAIL.n31 4.38563
R900 VTAIL.n122 VTAIL.n121 4.38563
R901 VTAIL.n214 VTAIL.n213 4.38563
R902 VTAIL.n579 VTAIL.n578 4.38563
R903 VTAIL.n487 VTAIL.n486 4.38563
R904 VTAIL.n397 VTAIL.n396 4.38563
R905 VTAIL.n305 VTAIL.n304 4.38563
R906 VTAIL.n682 VTAIL.n681 4.26717
R907 VTAIL.n698 VTAIL.n650 4.26717
R908 VTAIL.n46 VTAIL.n45 4.26717
R909 VTAIL.n62 VTAIL.n14 4.26717
R910 VTAIL.n136 VTAIL.n135 4.26717
R911 VTAIL.n152 VTAIL.n104 4.26717
R912 VTAIL.n228 VTAIL.n227 4.26717
R913 VTAIL.n244 VTAIL.n196 4.26717
R914 VTAIL.n609 VTAIL.n561 4.26717
R915 VTAIL.n593 VTAIL.n592 4.26717
R916 VTAIL.n517 VTAIL.n469 4.26717
R917 VTAIL.n501 VTAIL.n500 4.26717
R918 VTAIL.n427 VTAIL.n379 4.26717
R919 VTAIL.n411 VTAIL.n410 4.26717
R920 VTAIL.n335 VTAIL.n287 4.26717
R921 VTAIL.n319 VTAIL.n318 4.26717
R922 VTAIL.n678 VTAIL.n660 3.49141
R923 VTAIL.n702 VTAIL.n701 3.49141
R924 VTAIL.n726 VTAIL.n638 3.49141
R925 VTAIL.n42 VTAIL.n24 3.49141
R926 VTAIL.n66 VTAIL.n65 3.49141
R927 VTAIL.n90 VTAIL.n2 3.49141
R928 VTAIL.n132 VTAIL.n114 3.49141
R929 VTAIL.n156 VTAIL.n155 3.49141
R930 VTAIL.n180 VTAIL.n92 3.49141
R931 VTAIL.n224 VTAIL.n206 3.49141
R932 VTAIL.n248 VTAIL.n247 3.49141
R933 VTAIL.n272 VTAIL.n184 3.49141
R934 VTAIL.n636 VTAIL.n548 3.49141
R935 VTAIL.n613 VTAIL.n612 3.49141
R936 VTAIL.n589 VTAIL.n571 3.49141
R937 VTAIL.n544 VTAIL.n456 3.49141
R938 VTAIL.n521 VTAIL.n520 3.49141
R939 VTAIL.n497 VTAIL.n479 3.49141
R940 VTAIL.n454 VTAIL.n366 3.49141
R941 VTAIL.n431 VTAIL.n430 3.49141
R942 VTAIL.n407 VTAIL.n389 3.49141
R943 VTAIL.n362 VTAIL.n274 3.49141
R944 VTAIL.n339 VTAIL.n338 3.49141
R945 VTAIL.n315 VTAIL.n297 3.49141
R946 VTAIL.n677 VTAIL.n662 2.71565
R947 VTAIL.n705 VTAIL.n648 2.71565
R948 VTAIL.n724 VTAIL.n723 2.71565
R949 VTAIL.n41 VTAIL.n26 2.71565
R950 VTAIL.n69 VTAIL.n12 2.71565
R951 VTAIL.n88 VTAIL.n87 2.71565
R952 VTAIL.n131 VTAIL.n116 2.71565
R953 VTAIL.n159 VTAIL.n102 2.71565
R954 VTAIL.n178 VTAIL.n177 2.71565
R955 VTAIL.n223 VTAIL.n208 2.71565
R956 VTAIL.n251 VTAIL.n194 2.71565
R957 VTAIL.n270 VTAIL.n269 2.71565
R958 VTAIL.n634 VTAIL.n633 2.71565
R959 VTAIL.n616 VTAIL.n559 2.71565
R960 VTAIL.n588 VTAIL.n573 2.71565
R961 VTAIL.n542 VTAIL.n541 2.71565
R962 VTAIL.n524 VTAIL.n467 2.71565
R963 VTAIL.n496 VTAIL.n481 2.71565
R964 VTAIL.n452 VTAIL.n451 2.71565
R965 VTAIL.n434 VTAIL.n377 2.71565
R966 VTAIL.n406 VTAIL.n391 2.71565
R967 VTAIL.n360 VTAIL.n359 2.71565
R968 VTAIL.n342 VTAIL.n285 2.71565
R969 VTAIL.n314 VTAIL.n299 2.71565
R970 VTAIL.n365 VTAIL.n363 2.31084
R971 VTAIL.n455 VTAIL.n365 2.31084
R972 VTAIL.n547 VTAIL.n545 2.31084
R973 VTAIL.n637 VTAIL.n547 2.31084
R974 VTAIL.n273 VTAIL.n183 2.31084
R975 VTAIL.n183 VTAIL.n181 2.31084
R976 VTAIL.n91 VTAIL.n1 2.31084
R977 VTAIL VTAIL.n727 2.25266
R978 VTAIL.n674 VTAIL.n673 1.93989
R979 VTAIL.n706 VTAIL.n646 1.93989
R980 VTAIL.n720 VTAIL.n640 1.93989
R981 VTAIL.n38 VTAIL.n37 1.93989
R982 VTAIL.n70 VTAIL.n10 1.93989
R983 VTAIL.n84 VTAIL.n4 1.93989
R984 VTAIL.n128 VTAIL.n127 1.93989
R985 VTAIL.n160 VTAIL.n100 1.93989
R986 VTAIL.n174 VTAIL.n94 1.93989
R987 VTAIL.n220 VTAIL.n219 1.93989
R988 VTAIL.n252 VTAIL.n192 1.93989
R989 VTAIL.n266 VTAIL.n186 1.93989
R990 VTAIL.n630 VTAIL.n550 1.93989
R991 VTAIL.n617 VTAIL.n557 1.93989
R992 VTAIL.n585 VTAIL.n584 1.93989
R993 VTAIL.n538 VTAIL.n458 1.93989
R994 VTAIL.n525 VTAIL.n465 1.93989
R995 VTAIL.n493 VTAIL.n492 1.93989
R996 VTAIL.n448 VTAIL.n368 1.93989
R997 VTAIL.n435 VTAIL.n375 1.93989
R998 VTAIL.n403 VTAIL.n402 1.93989
R999 VTAIL.n356 VTAIL.n276 1.93989
R1000 VTAIL.n343 VTAIL.n283 1.93989
R1001 VTAIL.n311 VTAIL.n310 1.93989
R1002 VTAIL.n0 VTAIL.t4 1.21746
R1003 VTAIL.n0 VTAIL.t2 1.21746
R1004 VTAIL.n182 VTAIL.t13 1.21746
R1005 VTAIL.n182 VTAIL.t10 1.21746
R1006 VTAIL.n546 VTAIL.t9 1.21746
R1007 VTAIL.n546 VTAIL.t12 1.21746
R1008 VTAIL.n364 VTAIL.t5 1.21746
R1009 VTAIL.n364 VTAIL.t7 1.21746
R1010 VTAIL.n670 VTAIL.n664 1.16414
R1011 VTAIL.n711 VTAIL.n709 1.16414
R1012 VTAIL.n719 VTAIL.n642 1.16414
R1013 VTAIL.n34 VTAIL.n28 1.16414
R1014 VTAIL.n75 VTAIL.n73 1.16414
R1015 VTAIL.n83 VTAIL.n6 1.16414
R1016 VTAIL.n124 VTAIL.n118 1.16414
R1017 VTAIL.n165 VTAIL.n163 1.16414
R1018 VTAIL.n173 VTAIL.n96 1.16414
R1019 VTAIL.n216 VTAIL.n210 1.16414
R1020 VTAIL.n257 VTAIL.n255 1.16414
R1021 VTAIL.n265 VTAIL.n188 1.16414
R1022 VTAIL.n629 VTAIL.n552 1.16414
R1023 VTAIL.n621 VTAIL.n620 1.16414
R1024 VTAIL.n581 VTAIL.n575 1.16414
R1025 VTAIL.n537 VTAIL.n460 1.16414
R1026 VTAIL.n529 VTAIL.n528 1.16414
R1027 VTAIL.n489 VTAIL.n483 1.16414
R1028 VTAIL.n447 VTAIL.n370 1.16414
R1029 VTAIL.n439 VTAIL.n438 1.16414
R1030 VTAIL.n399 VTAIL.n393 1.16414
R1031 VTAIL.n355 VTAIL.n278 1.16414
R1032 VTAIL.n347 VTAIL.n346 1.16414
R1033 VTAIL.n307 VTAIL.n301 1.16414
R1034 VTAIL.n545 VTAIL.n455 0.470328
R1035 VTAIL.n181 VTAIL.n91 0.470328
R1036 VTAIL.n669 VTAIL.n666 0.388379
R1037 VTAIL.n710 VTAIL.n644 0.388379
R1038 VTAIL.n716 VTAIL.n715 0.388379
R1039 VTAIL.n33 VTAIL.n30 0.388379
R1040 VTAIL.n74 VTAIL.n8 0.388379
R1041 VTAIL.n80 VTAIL.n79 0.388379
R1042 VTAIL.n123 VTAIL.n120 0.388379
R1043 VTAIL.n164 VTAIL.n98 0.388379
R1044 VTAIL.n170 VTAIL.n169 0.388379
R1045 VTAIL.n215 VTAIL.n212 0.388379
R1046 VTAIL.n256 VTAIL.n190 0.388379
R1047 VTAIL.n262 VTAIL.n261 0.388379
R1048 VTAIL.n626 VTAIL.n625 0.388379
R1049 VTAIL.n556 VTAIL.n554 0.388379
R1050 VTAIL.n580 VTAIL.n577 0.388379
R1051 VTAIL.n534 VTAIL.n533 0.388379
R1052 VTAIL.n464 VTAIL.n462 0.388379
R1053 VTAIL.n488 VTAIL.n485 0.388379
R1054 VTAIL.n444 VTAIL.n443 0.388379
R1055 VTAIL.n374 VTAIL.n372 0.388379
R1056 VTAIL.n398 VTAIL.n395 0.388379
R1057 VTAIL.n352 VTAIL.n351 0.388379
R1058 VTAIL.n282 VTAIL.n280 0.388379
R1059 VTAIL.n306 VTAIL.n303 0.388379
R1060 VTAIL.n668 VTAIL.n663 0.155672
R1061 VTAIL.n675 VTAIL.n663 0.155672
R1062 VTAIL.n676 VTAIL.n675 0.155672
R1063 VTAIL.n676 VTAIL.n659 0.155672
R1064 VTAIL.n683 VTAIL.n659 0.155672
R1065 VTAIL.n684 VTAIL.n683 0.155672
R1066 VTAIL.n684 VTAIL.n655 0.155672
R1067 VTAIL.n691 VTAIL.n655 0.155672
R1068 VTAIL.n692 VTAIL.n691 0.155672
R1069 VTAIL.n692 VTAIL.n651 0.155672
R1070 VTAIL.n699 VTAIL.n651 0.155672
R1071 VTAIL.n700 VTAIL.n699 0.155672
R1072 VTAIL.n700 VTAIL.n647 0.155672
R1073 VTAIL.n707 VTAIL.n647 0.155672
R1074 VTAIL.n708 VTAIL.n707 0.155672
R1075 VTAIL.n708 VTAIL.n643 0.155672
R1076 VTAIL.n717 VTAIL.n643 0.155672
R1077 VTAIL.n718 VTAIL.n717 0.155672
R1078 VTAIL.n718 VTAIL.n639 0.155672
R1079 VTAIL.n725 VTAIL.n639 0.155672
R1080 VTAIL.n32 VTAIL.n27 0.155672
R1081 VTAIL.n39 VTAIL.n27 0.155672
R1082 VTAIL.n40 VTAIL.n39 0.155672
R1083 VTAIL.n40 VTAIL.n23 0.155672
R1084 VTAIL.n47 VTAIL.n23 0.155672
R1085 VTAIL.n48 VTAIL.n47 0.155672
R1086 VTAIL.n48 VTAIL.n19 0.155672
R1087 VTAIL.n55 VTAIL.n19 0.155672
R1088 VTAIL.n56 VTAIL.n55 0.155672
R1089 VTAIL.n56 VTAIL.n15 0.155672
R1090 VTAIL.n63 VTAIL.n15 0.155672
R1091 VTAIL.n64 VTAIL.n63 0.155672
R1092 VTAIL.n64 VTAIL.n11 0.155672
R1093 VTAIL.n71 VTAIL.n11 0.155672
R1094 VTAIL.n72 VTAIL.n71 0.155672
R1095 VTAIL.n72 VTAIL.n7 0.155672
R1096 VTAIL.n81 VTAIL.n7 0.155672
R1097 VTAIL.n82 VTAIL.n81 0.155672
R1098 VTAIL.n82 VTAIL.n3 0.155672
R1099 VTAIL.n89 VTAIL.n3 0.155672
R1100 VTAIL.n122 VTAIL.n117 0.155672
R1101 VTAIL.n129 VTAIL.n117 0.155672
R1102 VTAIL.n130 VTAIL.n129 0.155672
R1103 VTAIL.n130 VTAIL.n113 0.155672
R1104 VTAIL.n137 VTAIL.n113 0.155672
R1105 VTAIL.n138 VTAIL.n137 0.155672
R1106 VTAIL.n138 VTAIL.n109 0.155672
R1107 VTAIL.n145 VTAIL.n109 0.155672
R1108 VTAIL.n146 VTAIL.n145 0.155672
R1109 VTAIL.n146 VTAIL.n105 0.155672
R1110 VTAIL.n153 VTAIL.n105 0.155672
R1111 VTAIL.n154 VTAIL.n153 0.155672
R1112 VTAIL.n154 VTAIL.n101 0.155672
R1113 VTAIL.n161 VTAIL.n101 0.155672
R1114 VTAIL.n162 VTAIL.n161 0.155672
R1115 VTAIL.n162 VTAIL.n97 0.155672
R1116 VTAIL.n171 VTAIL.n97 0.155672
R1117 VTAIL.n172 VTAIL.n171 0.155672
R1118 VTAIL.n172 VTAIL.n93 0.155672
R1119 VTAIL.n179 VTAIL.n93 0.155672
R1120 VTAIL.n214 VTAIL.n209 0.155672
R1121 VTAIL.n221 VTAIL.n209 0.155672
R1122 VTAIL.n222 VTAIL.n221 0.155672
R1123 VTAIL.n222 VTAIL.n205 0.155672
R1124 VTAIL.n229 VTAIL.n205 0.155672
R1125 VTAIL.n230 VTAIL.n229 0.155672
R1126 VTAIL.n230 VTAIL.n201 0.155672
R1127 VTAIL.n237 VTAIL.n201 0.155672
R1128 VTAIL.n238 VTAIL.n237 0.155672
R1129 VTAIL.n238 VTAIL.n197 0.155672
R1130 VTAIL.n245 VTAIL.n197 0.155672
R1131 VTAIL.n246 VTAIL.n245 0.155672
R1132 VTAIL.n246 VTAIL.n193 0.155672
R1133 VTAIL.n253 VTAIL.n193 0.155672
R1134 VTAIL.n254 VTAIL.n253 0.155672
R1135 VTAIL.n254 VTAIL.n189 0.155672
R1136 VTAIL.n263 VTAIL.n189 0.155672
R1137 VTAIL.n264 VTAIL.n263 0.155672
R1138 VTAIL.n264 VTAIL.n185 0.155672
R1139 VTAIL.n271 VTAIL.n185 0.155672
R1140 VTAIL.n635 VTAIL.n549 0.155672
R1141 VTAIL.n628 VTAIL.n549 0.155672
R1142 VTAIL.n628 VTAIL.n627 0.155672
R1143 VTAIL.n627 VTAIL.n553 0.155672
R1144 VTAIL.n619 VTAIL.n553 0.155672
R1145 VTAIL.n619 VTAIL.n618 0.155672
R1146 VTAIL.n618 VTAIL.n558 0.155672
R1147 VTAIL.n611 VTAIL.n558 0.155672
R1148 VTAIL.n611 VTAIL.n610 0.155672
R1149 VTAIL.n610 VTAIL.n562 0.155672
R1150 VTAIL.n603 VTAIL.n562 0.155672
R1151 VTAIL.n603 VTAIL.n602 0.155672
R1152 VTAIL.n602 VTAIL.n566 0.155672
R1153 VTAIL.n595 VTAIL.n566 0.155672
R1154 VTAIL.n595 VTAIL.n594 0.155672
R1155 VTAIL.n594 VTAIL.n570 0.155672
R1156 VTAIL.n587 VTAIL.n570 0.155672
R1157 VTAIL.n587 VTAIL.n586 0.155672
R1158 VTAIL.n586 VTAIL.n574 0.155672
R1159 VTAIL.n579 VTAIL.n574 0.155672
R1160 VTAIL.n543 VTAIL.n457 0.155672
R1161 VTAIL.n536 VTAIL.n457 0.155672
R1162 VTAIL.n536 VTAIL.n535 0.155672
R1163 VTAIL.n535 VTAIL.n461 0.155672
R1164 VTAIL.n527 VTAIL.n461 0.155672
R1165 VTAIL.n527 VTAIL.n526 0.155672
R1166 VTAIL.n526 VTAIL.n466 0.155672
R1167 VTAIL.n519 VTAIL.n466 0.155672
R1168 VTAIL.n519 VTAIL.n518 0.155672
R1169 VTAIL.n518 VTAIL.n470 0.155672
R1170 VTAIL.n511 VTAIL.n470 0.155672
R1171 VTAIL.n511 VTAIL.n510 0.155672
R1172 VTAIL.n510 VTAIL.n474 0.155672
R1173 VTAIL.n503 VTAIL.n474 0.155672
R1174 VTAIL.n503 VTAIL.n502 0.155672
R1175 VTAIL.n502 VTAIL.n478 0.155672
R1176 VTAIL.n495 VTAIL.n478 0.155672
R1177 VTAIL.n495 VTAIL.n494 0.155672
R1178 VTAIL.n494 VTAIL.n482 0.155672
R1179 VTAIL.n487 VTAIL.n482 0.155672
R1180 VTAIL.n453 VTAIL.n367 0.155672
R1181 VTAIL.n446 VTAIL.n367 0.155672
R1182 VTAIL.n446 VTAIL.n445 0.155672
R1183 VTAIL.n445 VTAIL.n371 0.155672
R1184 VTAIL.n437 VTAIL.n371 0.155672
R1185 VTAIL.n437 VTAIL.n436 0.155672
R1186 VTAIL.n436 VTAIL.n376 0.155672
R1187 VTAIL.n429 VTAIL.n376 0.155672
R1188 VTAIL.n429 VTAIL.n428 0.155672
R1189 VTAIL.n428 VTAIL.n380 0.155672
R1190 VTAIL.n421 VTAIL.n380 0.155672
R1191 VTAIL.n421 VTAIL.n420 0.155672
R1192 VTAIL.n420 VTAIL.n384 0.155672
R1193 VTAIL.n413 VTAIL.n384 0.155672
R1194 VTAIL.n413 VTAIL.n412 0.155672
R1195 VTAIL.n412 VTAIL.n388 0.155672
R1196 VTAIL.n405 VTAIL.n388 0.155672
R1197 VTAIL.n405 VTAIL.n404 0.155672
R1198 VTAIL.n404 VTAIL.n392 0.155672
R1199 VTAIL.n397 VTAIL.n392 0.155672
R1200 VTAIL.n361 VTAIL.n275 0.155672
R1201 VTAIL.n354 VTAIL.n275 0.155672
R1202 VTAIL.n354 VTAIL.n353 0.155672
R1203 VTAIL.n353 VTAIL.n279 0.155672
R1204 VTAIL.n345 VTAIL.n279 0.155672
R1205 VTAIL.n345 VTAIL.n344 0.155672
R1206 VTAIL.n344 VTAIL.n284 0.155672
R1207 VTAIL.n337 VTAIL.n284 0.155672
R1208 VTAIL.n337 VTAIL.n336 0.155672
R1209 VTAIL.n336 VTAIL.n288 0.155672
R1210 VTAIL.n329 VTAIL.n288 0.155672
R1211 VTAIL.n329 VTAIL.n328 0.155672
R1212 VTAIL.n328 VTAIL.n292 0.155672
R1213 VTAIL.n321 VTAIL.n292 0.155672
R1214 VTAIL.n321 VTAIL.n320 0.155672
R1215 VTAIL.n320 VTAIL.n296 0.155672
R1216 VTAIL.n313 VTAIL.n296 0.155672
R1217 VTAIL.n313 VTAIL.n312 0.155672
R1218 VTAIL.n312 VTAIL.n300 0.155672
R1219 VTAIL.n305 VTAIL.n300 0.155672
R1220 VTAIL VTAIL.n1 0.0586897
R1221 B.n979 B.n978 585
R1222 B.n383 B.n147 585
R1223 B.n382 B.n381 585
R1224 B.n380 B.n379 585
R1225 B.n378 B.n377 585
R1226 B.n376 B.n375 585
R1227 B.n374 B.n373 585
R1228 B.n372 B.n371 585
R1229 B.n370 B.n369 585
R1230 B.n368 B.n367 585
R1231 B.n366 B.n365 585
R1232 B.n364 B.n363 585
R1233 B.n362 B.n361 585
R1234 B.n360 B.n359 585
R1235 B.n358 B.n357 585
R1236 B.n356 B.n355 585
R1237 B.n354 B.n353 585
R1238 B.n352 B.n351 585
R1239 B.n350 B.n349 585
R1240 B.n348 B.n347 585
R1241 B.n346 B.n345 585
R1242 B.n344 B.n343 585
R1243 B.n342 B.n341 585
R1244 B.n340 B.n339 585
R1245 B.n338 B.n337 585
R1246 B.n336 B.n335 585
R1247 B.n334 B.n333 585
R1248 B.n332 B.n331 585
R1249 B.n330 B.n329 585
R1250 B.n328 B.n327 585
R1251 B.n326 B.n325 585
R1252 B.n324 B.n323 585
R1253 B.n322 B.n321 585
R1254 B.n320 B.n319 585
R1255 B.n318 B.n317 585
R1256 B.n316 B.n315 585
R1257 B.n314 B.n313 585
R1258 B.n312 B.n311 585
R1259 B.n310 B.n309 585
R1260 B.n308 B.n307 585
R1261 B.n306 B.n305 585
R1262 B.n304 B.n303 585
R1263 B.n302 B.n301 585
R1264 B.n300 B.n299 585
R1265 B.n298 B.n297 585
R1266 B.n296 B.n295 585
R1267 B.n294 B.n293 585
R1268 B.n292 B.n291 585
R1269 B.n290 B.n289 585
R1270 B.n288 B.n287 585
R1271 B.n286 B.n285 585
R1272 B.n284 B.n283 585
R1273 B.n282 B.n281 585
R1274 B.n280 B.n279 585
R1275 B.n278 B.n277 585
R1276 B.n276 B.n275 585
R1277 B.n274 B.n273 585
R1278 B.n272 B.n271 585
R1279 B.n270 B.n269 585
R1280 B.n268 B.n267 585
R1281 B.n266 B.n265 585
R1282 B.n264 B.n263 585
R1283 B.n262 B.n261 585
R1284 B.n260 B.n259 585
R1285 B.n258 B.n257 585
R1286 B.n256 B.n255 585
R1287 B.n254 B.n253 585
R1288 B.n252 B.n251 585
R1289 B.n250 B.n249 585
R1290 B.n248 B.n247 585
R1291 B.n246 B.n245 585
R1292 B.n244 B.n243 585
R1293 B.n242 B.n241 585
R1294 B.n240 B.n239 585
R1295 B.n238 B.n237 585
R1296 B.n236 B.n235 585
R1297 B.n234 B.n233 585
R1298 B.n232 B.n231 585
R1299 B.n230 B.n229 585
R1300 B.n228 B.n227 585
R1301 B.n226 B.n225 585
R1302 B.n224 B.n223 585
R1303 B.n222 B.n221 585
R1304 B.n220 B.n219 585
R1305 B.n218 B.n217 585
R1306 B.n216 B.n215 585
R1307 B.n214 B.n213 585
R1308 B.n212 B.n211 585
R1309 B.n210 B.n209 585
R1310 B.n208 B.n207 585
R1311 B.n206 B.n205 585
R1312 B.n204 B.n203 585
R1313 B.n202 B.n201 585
R1314 B.n200 B.n199 585
R1315 B.n198 B.n197 585
R1316 B.n196 B.n195 585
R1317 B.n194 B.n193 585
R1318 B.n192 B.n191 585
R1319 B.n190 B.n189 585
R1320 B.n188 B.n187 585
R1321 B.n186 B.n185 585
R1322 B.n184 B.n183 585
R1323 B.n182 B.n181 585
R1324 B.n180 B.n179 585
R1325 B.n178 B.n177 585
R1326 B.n176 B.n175 585
R1327 B.n174 B.n173 585
R1328 B.n172 B.n171 585
R1329 B.n170 B.n169 585
R1330 B.n168 B.n167 585
R1331 B.n166 B.n165 585
R1332 B.n164 B.n163 585
R1333 B.n162 B.n161 585
R1334 B.n160 B.n159 585
R1335 B.n158 B.n157 585
R1336 B.n156 B.n155 585
R1337 B.n89 B.n88 585
R1338 B.n984 B.n983 585
R1339 B.n977 B.n148 585
R1340 B.n148 B.n86 585
R1341 B.n976 B.n85 585
R1342 B.n988 B.n85 585
R1343 B.n975 B.n84 585
R1344 B.n989 B.n84 585
R1345 B.n974 B.n83 585
R1346 B.n990 B.n83 585
R1347 B.n973 B.n972 585
R1348 B.n972 B.n79 585
R1349 B.n971 B.n78 585
R1350 B.n996 B.n78 585
R1351 B.n970 B.n77 585
R1352 B.n997 B.n77 585
R1353 B.n969 B.n76 585
R1354 B.n998 B.n76 585
R1355 B.n968 B.n967 585
R1356 B.n967 B.n72 585
R1357 B.n966 B.n71 585
R1358 B.n1004 B.n71 585
R1359 B.n965 B.n70 585
R1360 B.n1005 B.n70 585
R1361 B.n964 B.n69 585
R1362 B.n1006 B.n69 585
R1363 B.n963 B.n962 585
R1364 B.n962 B.n65 585
R1365 B.n961 B.n64 585
R1366 B.n1012 B.n64 585
R1367 B.n960 B.n63 585
R1368 B.n1013 B.n63 585
R1369 B.n959 B.n62 585
R1370 B.n1014 B.n62 585
R1371 B.n958 B.n957 585
R1372 B.n957 B.n58 585
R1373 B.n956 B.n57 585
R1374 B.n1020 B.n57 585
R1375 B.n955 B.n56 585
R1376 B.n1021 B.n56 585
R1377 B.n954 B.n55 585
R1378 B.n1022 B.n55 585
R1379 B.n953 B.n952 585
R1380 B.n952 B.n51 585
R1381 B.n951 B.n50 585
R1382 B.n1028 B.n50 585
R1383 B.n950 B.n49 585
R1384 B.n1029 B.n49 585
R1385 B.n949 B.n48 585
R1386 B.n1030 B.n48 585
R1387 B.n948 B.n947 585
R1388 B.n947 B.n44 585
R1389 B.n946 B.n43 585
R1390 B.n1036 B.n43 585
R1391 B.n945 B.n42 585
R1392 B.n1037 B.n42 585
R1393 B.n944 B.n41 585
R1394 B.n1038 B.n41 585
R1395 B.n943 B.n942 585
R1396 B.n942 B.n37 585
R1397 B.n941 B.n36 585
R1398 B.n1044 B.n36 585
R1399 B.n940 B.n35 585
R1400 B.n1045 B.n35 585
R1401 B.n939 B.n34 585
R1402 B.n1046 B.n34 585
R1403 B.n938 B.n937 585
R1404 B.n937 B.n30 585
R1405 B.n936 B.n29 585
R1406 B.n1052 B.n29 585
R1407 B.n935 B.n28 585
R1408 B.n1053 B.n28 585
R1409 B.n934 B.n27 585
R1410 B.n1054 B.n27 585
R1411 B.n933 B.n932 585
R1412 B.n932 B.n23 585
R1413 B.n931 B.n22 585
R1414 B.n1060 B.n22 585
R1415 B.n930 B.n21 585
R1416 B.n1061 B.n21 585
R1417 B.n929 B.n20 585
R1418 B.n1062 B.n20 585
R1419 B.n928 B.n927 585
R1420 B.n927 B.n16 585
R1421 B.n926 B.n15 585
R1422 B.n1068 B.n15 585
R1423 B.n925 B.n14 585
R1424 B.n1069 B.n14 585
R1425 B.n924 B.n13 585
R1426 B.n1070 B.n13 585
R1427 B.n923 B.n922 585
R1428 B.n922 B.n12 585
R1429 B.n921 B.n920 585
R1430 B.n921 B.n8 585
R1431 B.n919 B.n7 585
R1432 B.n1077 B.n7 585
R1433 B.n918 B.n6 585
R1434 B.n1078 B.n6 585
R1435 B.n917 B.n5 585
R1436 B.n1079 B.n5 585
R1437 B.n916 B.n915 585
R1438 B.n915 B.n4 585
R1439 B.n914 B.n384 585
R1440 B.n914 B.n913 585
R1441 B.n904 B.n385 585
R1442 B.n386 B.n385 585
R1443 B.n906 B.n905 585
R1444 B.n907 B.n906 585
R1445 B.n903 B.n391 585
R1446 B.n391 B.n390 585
R1447 B.n902 B.n901 585
R1448 B.n901 B.n900 585
R1449 B.n393 B.n392 585
R1450 B.n394 B.n393 585
R1451 B.n893 B.n892 585
R1452 B.n894 B.n893 585
R1453 B.n891 B.n399 585
R1454 B.n399 B.n398 585
R1455 B.n890 B.n889 585
R1456 B.n889 B.n888 585
R1457 B.n401 B.n400 585
R1458 B.n402 B.n401 585
R1459 B.n881 B.n880 585
R1460 B.n882 B.n881 585
R1461 B.n879 B.n406 585
R1462 B.n410 B.n406 585
R1463 B.n878 B.n877 585
R1464 B.n877 B.n876 585
R1465 B.n408 B.n407 585
R1466 B.n409 B.n408 585
R1467 B.n869 B.n868 585
R1468 B.n870 B.n869 585
R1469 B.n867 B.n415 585
R1470 B.n415 B.n414 585
R1471 B.n866 B.n865 585
R1472 B.n865 B.n864 585
R1473 B.n417 B.n416 585
R1474 B.n418 B.n417 585
R1475 B.n857 B.n856 585
R1476 B.n858 B.n857 585
R1477 B.n855 B.n422 585
R1478 B.n426 B.n422 585
R1479 B.n854 B.n853 585
R1480 B.n853 B.n852 585
R1481 B.n424 B.n423 585
R1482 B.n425 B.n424 585
R1483 B.n845 B.n844 585
R1484 B.n846 B.n845 585
R1485 B.n843 B.n431 585
R1486 B.n431 B.n430 585
R1487 B.n842 B.n841 585
R1488 B.n841 B.n840 585
R1489 B.n433 B.n432 585
R1490 B.n434 B.n433 585
R1491 B.n833 B.n832 585
R1492 B.n834 B.n833 585
R1493 B.n831 B.n438 585
R1494 B.n442 B.n438 585
R1495 B.n830 B.n829 585
R1496 B.n829 B.n828 585
R1497 B.n440 B.n439 585
R1498 B.n441 B.n440 585
R1499 B.n821 B.n820 585
R1500 B.n822 B.n821 585
R1501 B.n819 B.n447 585
R1502 B.n447 B.n446 585
R1503 B.n818 B.n817 585
R1504 B.n817 B.n816 585
R1505 B.n449 B.n448 585
R1506 B.n450 B.n449 585
R1507 B.n809 B.n808 585
R1508 B.n810 B.n809 585
R1509 B.n807 B.n455 585
R1510 B.n455 B.n454 585
R1511 B.n806 B.n805 585
R1512 B.n805 B.n804 585
R1513 B.n457 B.n456 585
R1514 B.n458 B.n457 585
R1515 B.n797 B.n796 585
R1516 B.n798 B.n797 585
R1517 B.n795 B.n463 585
R1518 B.n463 B.n462 585
R1519 B.n794 B.n793 585
R1520 B.n793 B.n792 585
R1521 B.n465 B.n464 585
R1522 B.n466 B.n465 585
R1523 B.n785 B.n784 585
R1524 B.n786 B.n785 585
R1525 B.n783 B.n471 585
R1526 B.n471 B.n470 585
R1527 B.n782 B.n781 585
R1528 B.n781 B.n780 585
R1529 B.n473 B.n472 585
R1530 B.n474 B.n473 585
R1531 B.n776 B.n775 585
R1532 B.n477 B.n476 585
R1533 B.n772 B.n771 585
R1534 B.n773 B.n772 585
R1535 B.n770 B.n536 585
R1536 B.n769 B.n768 585
R1537 B.n767 B.n766 585
R1538 B.n765 B.n764 585
R1539 B.n763 B.n762 585
R1540 B.n761 B.n760 585
R1541 B.n759 B.n758 585
R1542 B.n757 B.n756 585
R1543 B.n755 B.n754 585
R1544 B.n753 B.n752 585
R1545 B.n751 B.n750 585
R1546 B.n749 B.n748 585
R1547 B.n747 B.n746 585
R1548 B.n745 B.n744 585
R1549 B.n743 B.n742 585
R1550 B.n741 B.n740 585
R1551 B.n739 B.n738 585
R1552 B.n737 B.n736 585
R1553 B.n735 B.n734 585
R1554 B.n733 B.n732 585
R1555 B.n731 B.n730 585
R1556 B.n729 B.n728 585
R1557 B.n727 B.n726 585
R1558 B.n725 B.n724 585
R1559 B.n723 B.n722 585
R1560 B.n721 B.n720 585
R1561 B.n719 B.n718 585
R1562 B.n717 B.n716 585
R1563 B.n715 B.n714 585
R1564 B.n713 B.n712 585
R1565 B.n711 B.n710 585
R1566 B.n709 B.n708 585
R1567 B.n707 B.n706 585
R1568 B.n705 B.n704 585
R1569 B.n703 B.n702 585
R1570 B.n701 B.n700 585
R1571 B.n699 B.n698 585
R1572 B.n697 B.n696 585
R1573 B.n695 B.n694 585
R1574 B.n693 B.n692 585
R1575 B.n691 B.n690 585
R1576 B.n689 B.n688 585
R1577 B.n687 B.n686 585
R1578 B.n685 B.n684 585
R1579 B.n683 B.n682 585
R1580 B.n681 B.n680 585
R1581 B.n679 B.n678 585
R1582 B.n677 B.n676 585
R1583 B.n675 B.n674 585
R1584 B.n673 B.n672 585
R1585 B.n671 B.n670 585
R1586 B.n668 B.n667 585
R1587 B.n666 B.n665 585
R1588 B.n664 B.n663 585
R1589 B.n662 B.n661 585
R1590 B.n660 B.n659 585
R1591 B.n658 B.n657 585
R1592 B.n656 B.n655 585
R1593 B.n654 B.n653 585
R1594 B.n652 B.n651 585
R1595 B.n650 B.n649 585
R1596 B.n647 B.n646 585
R1597 B.n645 B.n644 585
R1598 B.n643 B.n642 585
R1599 B.n641 B.n640 585
R1600 B.n639 B.n638 585
R1601 B.n637 B.n636 585
R1602 B.n635 B.n634 585
R1603 B.n633 B.n632 585
R1604 B.n631 B.n630 585
R1605 B.n629 B.n628 585
R1606 B.n627 B.n626 585
R1607 B.n625 B.n624 585
R1608 B.n623 B.n622 585
R1609 B.n621 B.n620 585
R1610 B.n619 B.n618 585
R1611 B.n617 B.n616 585
R1612 B.n615 B.n614 585
R1613 B.n613 B.n612 585
R1614 B.n611 B.n610 585
R1615 B.n609 B.n608 585
R1616 B.n607 B.n606 585
R1617 B.n605 B.n604 585
R1618 B.n603 B.n602 585
R1619 B.n601 B.n600 585
R1620 B.n599 B.n598 585
R1621 B.n597 B.n596 585
R1622 B.n595 B.n594 585
R1623 B.n593 B.n592 585
R1624 B.n591 B.n590 585
R1625 B.n589 B.n588 585
R1626 B.n587 B.n586 585
R1627 B.n585 B.n584 585
R1628 B.n583 B.n582 585
R1629 B.n581 B.n580 585
R1630 B.n579 B.n578 585
R1631 B.n577 B.n576 585
R1632 B.n575 B.n574 585
R1633 B.n573 B.n572 585
R1634 B.n571 B.n570 585
R1635 B.n569 B.n568 585
R1636 B.n567 B.n566 585
R1637 B.n565 B.n564 585
R1638 B.n563 B.n562 585
R1639 B.n561 B.n560 585
R1640 B.n559 B.n558 585
R1641 B.n557 B.n556 585
R1642 B.n555 B.n554 585
R1643 B.n553 B.n552 585
R1644 B.n551 B.n550 585
R1645 B.n549 B.n548 585
R1646 B.n547 B.n546 585
R1647 B.n545 B.n544 585
R1648 B.n543 B.n542 585
R1649 B.n541 B.n535 585
R1650 B.n773 B.n535 585
R1651 B.n777 B.n475 585
R1652 B.n475 B.n474 585
R1653 B.n779 B.n778 585
R1654 B.n780 B.n779 585
R1655 B.n469 B.n468 585
R1656 B.n470 B.n469 585
R1657 B.n788 B.n787 585
R1658 B.n787 B.n786 585
R1659 B.n789 B.n467 585
R1660 B.n467 B.n466 585
R1661 B.n791 B.n790 585
R1662 B.n792 B.n791 585
R1663 B.n461 B.n460 585
R1664 B.n462 B.n461 585
R1665 B.n800 B.n799 585
R1666 B.n799 B.n798 585
R1667 B.n801 B.n459 585
R1668 B.n459 B.n458 585
R1669 B.n803 B.n802 585
R1670 B.n804 B.n803 585
R1671 B.n453 B.n452 585
R1672 B.n454 B.n453 585
R1673 B.n812 B.n811 585
R1674 B.n811 B.n810 585
R1675 B.n813 B.n451 585
R1676 B.n451 B.n450 585
R1677 B.n815 B.n814 585
R1678 B.n816 B.n815 585
R1679 B.n445 B.n444 585
R1680 B.n446 B.n445 585
R1681 B.n824 B.n823 585
R1682 B.n823 B.n822 585
R1683 B.n825 B.n443 585
R1684 B.n443 B.n441 585
R1685 B.n827 B.n826 585
R1686 B.n828 B.n827 585
R1687 B.n437 B.n436 585
R1688 B.n442 B.n437 585
R1689 B.n836 B.n835 585
R1690 B.n835 B.n834 585
R1691 B.n837 B.n435 585
R1692 B.n435 B.n434 585
R1693 B.n839 B.n838 585
R1694 B.n840 B.n839 585
R1695 B.n429 B.n428 585
R1696 B.n430 B.n429 585
R1697 B.n848 B.n847 585
R1698 B.n847 B.n846 585
R1699 B.n849 B.n427 585
R1700 B.n427 B.n425 585
R1701 B.n851 B.n850 585
R1702 B.n852 B.n851 585
R1703 B.n421 B.n420 585
R1704 B.n426 B.n421 585
R1705 B.n860 B.n859 585
R1706 B.n859 B.n858 585
R1707 B.n861 B.n419 585
R1708 B.n419 B.n418 585
R1709 B.n863 B.n862 585
R1710 B.n864 B.n863 585
R1711 B.n413 B.n412 585
R1712 B.n414 B.n413 585
R1713 B.n872 B.n871 585
R1714 B.n871 B.n870 585
R1715 B.n873 B.n411 585
R1716 B.n411 B.n409 585
R1717 B.n875 B.n874 585
R1718 B.n876 B.n875 585
R1719 B.n405 B.n404 585
R1720 B.n410 B.n405 585
R1721 B.n884 B.n883 585
R1722 B.n883 B.n882 585
R1723 B.n885 B.n403 585
R1724 B.n403 B.n402 585
R1725 B.n887 B.n886 585
R1726 B.n888 B.n887 585
R1727 B.n397 B.n396 585
R1728 B.n398 B.n397 585
R1729 B.n896 B.n895 585
R1730 B.n895 B.n894 585
R1731 B.n897 B.n395 585
R1732 B.n395 B.n394 585
R1733 B.n899 B.n898 585
R1734 B.n900 B.n899 585
R1735 B.n389 B.n388 585
R1736 B.n390 B.n389 585
R1737 B.n909 B.n908 585
R1738 B.n908 B.n907 585
R1739 B.n910 B.n387 585
R1740 B.n387 B.n386 585
R1741 B.n912 B.n911 585
R1742 B.n913 B.n912 585
R1743 B.n3 B.n0 585
R1744 B.n4 B.n3 585
R1745 B.n1076 B.n1 585
R1746 B.n1077 B.n1076 585
R1747 B.n1075 B.n1074 585
R1748 B.n1075 B.n8 585
R1749 B.n1073 B.n9 585
R1750 B.n12 B.n9 585
R1751 B.n1072 B.n1071 585
R1752 B.n1071 B.n1070 585
R1753 B.n11 B.n10 585
R1754 B.n1069 B.n11 585
R1755 B.n1067 B.n1066 585
R1756 B.n1068 B.n1067 585
R1757 B.n1065 B.n17 585
R1758 B.n17 B.n16 585
R1759 B.n1064 B.n1063 585
R1760 B.n1063 B.n1062 585
R1761 B.n19 B.n18 585
R1762 B.n1061 B.n19 585
R1763 B.n1059 B.n1058 585
R1764 B.n1060 B.n1059 585
R1765 B.n1057 B.n24 585
R1766 B.n24 B.n23 585
R1767 B.n1056 B.n1055 585
R1768 B.n1055 B.n1054 585
R1769 B.n26 B.n25 585
R1770 B.n1053 B.n26 585
R1771 B.n1051 B.n1050 585
R1772 B.n1052 B.n1051 585
R1773 B.n1049 B.n31 585
R1774 B.n31 B.n30 585
R1775 B.n1048 B.n1047 585
R1776 B.n1047 B.n1046 585
R1777 B.n33 B.n32 585
R1778 B.n1045 B.n33 585
R1779 B.n1043 B.n1042 585
R1780 B.n1044 B.n1043 585
R1781 B.n1041 B.n38 585
R1782 B.n38 B.n37 585
R1783 B.n1040 B.n1039 585
R1784 B.n1039 B.n1038 585
R1785 B.n40 B.n39 585
R1786 B.n1037 B.n40 585
R1787 B.n1035 B.n1034 585
R1788 B.n1036 B.n1035 585
R1789 B.n1033 B.n45 585
R1790 B.n45 B.n44 585
R1791 B.n1032 B.n1031 585
R1792 B.n1031 B.n1030 585
R1793 B.n47 B.n46 585
R1794 B.n1029 B.n47 585
R1795 B.n1027 B.n1026 585
R1796 B.n1028 B.n1027 585
R1797 B.n1025 B.n52 585
R1798 B.n52 B.n51 585
R1799 B.n1024 B.n1023 585
R1800 B.n1023 B.n1022 585
R1801 B.n54 B.n53 585
R1802 B.n1021 B.n54 585
R1803 B.n1019 B.n1018 585
R1804 B.n1020 B.n1019 585
R1805 B.n1017 B.n59 585
R1806 B.n59 B.n58 585
R1807 B.n1016 B.n1015 585
R1808 B.n1015 B.n1014 585
R1809 B.n61 B.n60 585
R1810 B.n1013 B.n61 585
R1811 B.n1011 B.n1010 585
R1812 B.n1012 B.n1011 585
R1813 B.n1009 B.n66 585
R1814 B.n66 B.n65 585
R1815 B.n1008 B.n1007 585
R1816 B.n1007 B.n1006 585
R1817 B.n68 B.n67 585
R1818 B.n1005 B.n68 585
R1819 B.n1003 B.n1002 585
R1820 B.n1004 B.n1003 585
R1821 B.n1001 B.n73 585
R1822 B.n73 B.n72 585
R1823 B.n1000 B.n999 585
R1824 B.n999 B.n998 585
R1825 B.n75 B.n74 585
R1826 B.n997 B.n75 585
R1827 B.n995 B.n994 585
R1828 B.n996 B.n995 585
R1829 B.n993 B.n80 585
R1830 B.n80 B.n79 585
R1831 B.n992 B.n991 585
R1832 B.n991 B.n990 585
R1833 B.n82 B.n81 585
R1834 B.n989 B.n82 585
R1835 B.n987 B.n986 585
R1836 B.n988 B.n987 585
R1837 B.n985 B.n87 585
R1838 B.n87 B.n86 585
R1839 B.n1080 B.n1079 585
R1840 B.n1078 B.n2 585
R1841 B.n983 B.n87 497.305
R1842 B.n979 B.n148 497.305
R1843 B.n535 B.n473 497.305
R1844 B.n775 B.n475 497.305
R1845 B.n149 B.t14 407.943
R1846 B.n539 B.t21 407.943
R1847 B.n152 B.t17 407.943
R1848 B.n537 B.t11 407.943
R1849 B.n152 B.t16 374.49
R1850 B.n149 B.t12 374.49
R1851 B.n539 B.t19 374.49
R1852 B.n537 B.t8 374.49
R1853 B.n150 B.t15 355.967
R1854 B.n540 B.t20 355.967
R1855 B.n153 B.t18 355.967
R1856 B.n538 B.t10 355.967
R1857 B.n981 B.n980 256.663
R1858 B.n981 B.n146 256.663
R1859 B.n981 B.n145 256.663
R1860 B.n981 B.n144 256.663
R1861 B.n981 B.n143 256.663
R1862 B.n981 B.n142 256.663
R1863 B.n981 B.n141 256.663
R1864 B.n981 B.n140 256.663
R1865 B.n981 B.n139 256.663
R1866 B.n981 B.n138 256.663
R1867 B.n981 B.n137 256.663
R1868 B.n981 B.n136 256.663
R1869 B.n981 B.n135 256.663
R1870 B.n981 B.n134 256.663
R1871 B.n981 B.n133 256.663
R1872 B.n981 B.n132 256.663
R1873 B.n981 B.n131 256.663
R1874 B.n981 B.n130 256.663
R1875 B.n981 B.n129 256.663
R1876 B.n981 B.n128 256.663
R1877 B.n981 B.n127 256.663
R1878 B.n981 B.n126 256.663
R1879 B.n981 B.n125 256.663
R1880 B.n981 B.n124 256.663
R1881 B.n981 B.n123 256.663
R1882 B.n981 B.n122 256.663
R1883 B.n981 B.n121 256.663
R1884 B.n981 B.n120 256.663
R1885 B.n981 B.n119 256.663
R1886 B.n981 B.n118 256.663
R1887 B.n981 B.n117 256.663
R1888 B.n981 B.n116 256.663
R1889 B.n981 B.n115 256.663
R1890 B.n981 B.n114 256.663
R1891 B.n981 B.n113 256.663
R1892 B.n981 B.n112 256.663
R1893 B.n981 B.n111 256.663
R1894 B.n981 B.n110 256.663
R1895 B.n981 B.n109 256.663
R1896 B.n981 B.n108 256.663
R1897 B.n981 B.n107 256.663
R1898 B.n981 B.n106 256.663
R1899 B.n981 B.n105 256.663
R1900 B.n981 B.n104 256.663
R1901 B.n981 B.n103 256.663
R1902 B.n981 B.n102 256.663
R1903 B.n981 B.n101 256.663
R1904 B.n981 B.n100 256.663
R1905 B.n981 B.n99 256.663
R1906 B.n981 B.n98 256.663
R1907 B.n981 B.n97 256.663
R1908 B.n981 B.n96 256.663
R1909 B.n981 B.n95 256.663
R1910 B.n981 B.n94 256.663
R1911 B.n981 B.n93 256.663
R1912 B.n981 B.n92 256.663
R1913 B.n981 B.n91 256.663
R1914 B.n981 B.n90 256.663
R1915 B.n982 B.n981 256.663
R1916 B.n774 B.n773 256.663
R1917 B.n773 B.n478 256.663
R1918 B.n773 B.n479 256.663
R1919 B.n773 B.n480 256.663
R1920 B.n773 B.n481 256.663
R1921 B.n773 B.n482 256.663
R1922 B.n773 B.n483 256.663
R1923 B.n773 B.n484 256.663
R1924 B.n773 B.n485 256.663
R1925 B.n773 B.n486 256.663
R1926 B.n773 B.n487 256.663
R1927 B.n773 B.n488 256.663
R1928 B.n773 B.n489 256.663
R1929 B.n773 B.n490 256.663
R1930 B.n773 B.n491 256.663
R1931 B.n773 B.n492 256.663
R1932 B.n773 B.n493 256.663
R1933 B.n773 B.n494 256.663
R1934 B.n773 B.n495 256.663
R1935 B.n773 B.n496 256.663
R1936 B.n773 B.n497 256.663
R1937 B.n773 B.n498 256.663
R1938 B.n773 B.n499 256.663
R1939 B.n773 B.n500 256.663
R1940 B.n773 B.n501 256.663
R1941 B.n773 B.n502 256.663
R1942 B.n773 B.n503 256.663
R1943 B.n773 B.n504 256.663
R1944 B.n773 B.n505 256.663
R1945 B.n773 B.n506 256.663
R1946 B.n773 B.n507 256.663
R1947 B.n773 B.n508 256.663
R1948 B.n773 B.n509 256.663
R1949 B.n773 B.n510 256.663
R1950 B.n773 B.n511 256.663
R1951 B.n773 B.n512 256.663
R1952 B.n773 B.n513 256.663
R1953 B.n773 B.n514 256.663
R1954 B.n773 B.n515 256.663
R1955 B.n773 B.n516 256.663
R1956 B.n773 B.n517 256.663
R1957 B.n773 B.n518 256.663
R1958 B.n773 B.n519 256.663
R1959 B.n773 B.n520 256.663
R1960 B.n773 B.n521 256.663
R1961 B.n773 B.n522 256.663
R1962 B.n773 B.n523 256.663
R1963 B.n773 B.n524 256.663
R1964 B.n773 B.n525 256.663
R1965 B.n773 B.n526 256.663
R1966 B.n773 B.n527 256.663
R1967 B.n773 B.n528 256.663
R1968 B.n773 B.n529 256.663
R1969 B.n773 B.n530 256.663
R1970 B.n773 B.n531 256.663
R1971 B.n773 B.n532 256.663
R1972 B.n773 B.n533 256.663
R1973 B.n773 B.n534 256.663
R1974 B.n1082 B.n1081 256.663
R1975 B.n155 B.n89 163.367
R1976 B.n159 B.n158 163.367
R1977 B.n163 B.n162 163.367
R1978 B.n167 B.n166 163.367
R1979 B.n171 B.n170 163.367
R1980 B.n175 B.n174 163.367
R1981 B.n179 B.n178 163.367
R1982 B.n183 B.n182 163.367
R1983 B.n187 B.n186 163.367
R1984 B.n191 B.n190 163.367
R1985 B.n195 B.n194 163.367
R1986 B.n199 B.n198 163.367
R1987 B.n203 B.n202 163.367
R1988 B.n207 B.n206 163.367
R1989 B.n211 B.n210 163.367
R1990 B.n215 B.n214 163.367
R1991 B.n219 B.n218 163.367
R1992 B.n223 B.n222 163.367
R1993 B.n227 B.n226 163.367
R1994 B.n231 B.n230 163.367
R1995 B.n235 B.n234 163.367
R1996 B.n239 B.n238 163.367
R1997 B.n243 B.n242 163.367
R1998 B.n247 B.n246 163.367
R1999 B.n251 B.n250 163.367
R2000 B.n255 B.n254 163.367
R2001 B.n259 B.n258 163.367
R2002 B.n263 B.n262 163.367
R2003 B.n267 B.n266 163.367
R2004 B.n271 B.n270 163.367
R2005 B.n275 B.n274 163.367
R2006 B.n279 B.n278 163.367
R2007 B.n283 B.n282 163.367
R2008 B.n287 B.n286 163.367
R2009 B.n291 B.n290 163.367
R2010 B.n295 B.n294 163.367
R2011 B.n299 B.n298 163.367
R2012 B.n303 B.n302 163.367
R2013 B.n307 B.n306 163.367
R2014 B.n311 B.n310 163.367
R2015 B.n315 B.n314 163.367
R2016 B.n319 B.n318 163.367
R2017 B.n323 B.n322 163.367
R2018 B.n327 B.n326 163.367
R2019 B.n331 B.n330 163.367
R2020 B.n335 B.n334 163.367
R2021 B.n339 B.n338 163.367
R2022 B.n343 B.n342 163.367
R2023 B.n347 B.n346 163.367
R2024 B.n351 B.n350 163.367
R2025 B.n355 B.n354 163.367
R2026 B.n359 B.n358 163.367
R2027 B.n363 B.n362 163.367
R2028 B.n367 B.n366 163.367
R2029 B.n371 B.n370 163.367
R2030 B.n375 B.n374 163.367
R2031 B.n379 B.n378 163.367
R2032 B.n381 B.n147 163.367
R2033 B.n781 B.n473 163.367
R2034 B.n781 B.n471 163.367
R2035 B.n785 B.n471 163.367
R2036 B.n785 B.n465 163.367
R2037 B.n793 B.n465 163.367
R2038 B.n793 B.n463 163.367
R2039 B.n797 B.n463 163.367
R2040 B.n797 B.n457 163.367
R2041 B.n805 B.n457 163.367
R2042 B.n805 B.n455 163.367
R2043 B.n809 B.n455 163.367
R2044 B.n809 B.n449 163.367
R2045 B.n817 B.n449 163.367
R2046 B.n817 B.n447 163.367
R2047 B.n821 B.n447 163.367
R2048 B.n821 B.n440 163.367
R2049 B.n829 B.n440 163.367
R2050 B.n829 B.n438 163.367
R2051 B.n833 B.n438 163.367
R2052 B.n833 B.n433 163.367
R2053 B.n841 B.n433 163.367
R2054 B.n841 B.n431 163.367
R2055 B.n845 B.n431 163.367
R2056 B.n845 B.n424 163.367
R2057 B.n853 B.n424 163.367
R2058 B.n853 B.n422 163.367
R2059 B.n857 B.n422 163.367
R2060 B.n857 B.n417 163.367
R2061 B.n865 B.n417 163.367
R2062 B.n865 B.n415 163.367
R2063 B.n869 B.n415 163.367
R2064 B.n869 B.n408 163.367
R2065 B.n877 B.n408 163.367
R2066 B.n877 B.n406 163.367
R2067 B.n881 B.n406 163.367
R2068 B.n881 B.n401 163.367
R2069 B.n889 B.n401 163.367
R2070 B.n889 B.n399 163.367
R2071 B.n893 B.n399 163.367
R2072 B.n893 B.n393 163.367
R2073 B.n901 B.n393 163.367
R2074 B.n901 B.n391 163.367
R2075 B.n906 B.n391 163.367
R2076 B.n906 B.n385 163.367
R2077 B.n914 B.n385 163.367
R2078 B.n915 B.n914 163.367
R2079 B.n915 B.n5 163.367
R2080 B.n6 B.n5 163.367
R2081 B.n7 B.n6 163.367
R2082 B.n921 B.n7 163.367
R2083 B.n922 B.n921 163.367
R2084 B.n922 B.n13 163.367
R2085 B.n14 B.n13 163.367
R2086 B.n15 B.n14 163.367
R2087 B.n927 B.n15 163.367
R2088 B.n927 B.n20 163.367
R2089 B.n21 B.n20 163.367
R2090 B.n22 B.n21 163.367
R2091 B.n932 B.n22 163.367
R2092 B.n932 B.n27 163.367
R2093 B.n28 B.n27 163.367
R2094 B.n29 B.n28 163.367
R2095 B.n937 B.n29 163.367
R2096 B.n937 B.n34 163.367
R2097 B.n35 B.n34 163.367
R2098 B.n36 B.n35 163.367
R2099 B.n942 B.n36 163.367
R2100 B.n942 B.n41 163.367
R2101 B.n42 B.n41 163.367
R2102 B.n43 B.n42 163.367
R2103 B.n947 B.n43 163.367
R2104 B.n947 B.n48 163.367
R2105 B.n49 B.n48 163.367
R2106 B.n50 B.n49 163.367
R2107 B.n952 B.n50 163.367
R2108 B.n952 B.n55 163.367
R2109 B.n56 B.n55 163.367
R2110 B.n57 B.n56 163.367
R2111 B.n957 B.n57 163.367
R2112 B.n957 B.n62 163.367
R2113 B.n63 B.n62 163.367
R2114 B.n64 B.n63 163.367
R2115 B.n962 B.n64 163.367
R2116 B.n962 B.n69 163.367
R2117 B.n70 B.n69 163.367
R2118 B.n71 B.n70 163.367
R2119 B.n967 B.n71 163.367
R2120 B.n967 B.n76 163.367
R2121 B.n77 B.n76 163.367
R2122 B.n78 B.n77 163.367
R2123 B.n972 B.n78 163.367
R2124 B.n972 B.n83 163.367
R2125 B.n84 B.n83 163.367
R2126 B.n85 B.n84 163.367
R2127 B.n148 B.n85 163.367
R2128 B.n772 B.n477 163.367
R2129 B.n772 B.n536 163.367
R2130 B.n768 B.n767 163.367
R2131 B.n764 B.n763 163.367
R2132 B.n760 B.n759 163.367
R2133 B.n756 B.n755 163.367
R2134 B.n752 B.n751 163.367
R2135 B.n748 B.n747 163.367
R2136 B.n744 B.n743 163.367
R2137 B.n740 B.n739 163.367
R2138 B.n736 B.n735 163.367
R2139 B.n732 B.n731 163.367
R2140 B.n728 B.n727 163.367
R2141 B.n724 B.n723 163.367
R2142 B.n720 B.n719 163.367
R2143 B.n716 B.n715 163.367
R2144 B.n712 B.n711 163.367
R2145 B.n708 B.n707 163.367
R2146 B.n704 B.n703 163.367
R2147 B.n700 B.n699 163.367
R2148 B.n696 B.n695 163.367
R2149 B.n692 B.n691 163.367
R2150 B.n688 B.n687 163.367
R2151 B.n684 B.n683 163.367
R2152 B.n680 B.n679 163.367
R2153 B.n676 B.n675 163.367
R2154 B.n672 B.n671 163.367
R2155 B.n667 B.n666 163.367
R2156 B.n663 B.n662 163.367
R2157 B.n659 B.n658 163.367
R2158 B.n655 B.n654 163.367
R2159 B.n651 B.n650 163.367
R2160 B.n646 B.n645 163.367
R2161 B.n642 B.n641 163.367
R2162 B.n638 B.n637 163.367
R2163 B.n634 B.n633 163.367
R2164 B.n630 B.n629 163.367
R2165 B.n626 B.n625 163.367
R2166 B.n622 B.n621 163.367
R2167 B.n618 B.n617 163.367
R2168 B.n614 B.n613 163.367
R2169 B.n610 B.n609 163.367
R2170 B.n606 B.n605 163.367
R2171 B.n602 B.n601 163.367
R2172 B.n598 B.n597 163.367
R2173 B.n594 B.n593 163.367
R2174 B.n590 B.n589 163.367
R2175 B.n586 B.n585 163.367
R2176 B.n582 B.n581 163.367
R2177 B.n578 B.n577 163.367
R2178 B.n574 B.n573 163.367
R2179 B.n570 B.n569 163.367
R2180 B.n566 B.n565 163.367
R2181 B.n562 B.n561 163.367
R2182 B.n558 B.n557 163.367
R2183 B.n554 B.n553 163.367
R2184 B.n550 B.n549 163.367
R2185 B.n546 B.n545 163.367
R2186 B.n542 B.n535 163.367
R2187 B.n779 B.n475 163.367
R2188 B.n779 B.n469 163.367
R2189 B.n787 B.n469 163.367
R2190 B.n787 B.n467 163.367
R2191 B.n791 B.n467 163.367
R2192 B.n791 B.n461 163.367
R2193 B.n799 B.n461 163.367
R2194 B.n799 B.n459 163.367
R2195 B.n803 B.n459 163.367
R2196 B.n803 B.n453 163.367
R2197 B.n811 B.n453 163.367
R2198 B.n811 B.n451 163.367
R2199 B.n815 B.n451 163.367
R2200 B.n815 B.n445 163.367
R2201 B.n823 B.n445 163.367
R2202 B.n823 B.n443 163.367
R2203 B.n827 B.n443 163.367
R2204 B.n827 B.n437 163.367
R2205 B.n835 B.n437 163.367
R2206 B.n835 B.n435 163.367
R2207 B.n839 B.n435 163.367
R2208 B.n839 B.n429 163.367
R2209 B.n847 B.n429 163.367
R2210 B.n847 B.n427 163.367
R2211 B.n851 B.n427 163.367
R2212 B.n851 B.n421 163.367
R2213 B.n859 B.n421 163.367
R2214 B.n859 B.n419 163.367
R2215 B.n863 B.n419 163.367
R2216 B.n863 B.n413 163.367
R2217 B.n871 B.n413 163.367
R2218 B.n871 B.n411 163.367
R2219 B.n875 B.n411 163.367
R2220 B.n875 B.n405 163.367
R2221 B.n883 B.n405 163.367
R2222 B.n883 B.n403 163.367
R2223 B.n887 B.n403 163.367
R2224 B.n887 B.n397 163.367
R2225 B.n895 B.n397 163.367
R2226 B.n895 B.n395 163.367
R2227 B.n899 B.n395 163.367
R2228 B.n899 B.n389 163.367
R2229 B.n908 B.n389 163.367
R2230 B.n908 B.n387 163.367
R2231 B.n912 B.n387 163.367
R2232 B.n912 B.n3 163.367
R2233 B.n1080 B.n3 163.367
R2234 B.n1076 B.n2 163.367
R2235 B.n1076 B.n1075 163.367
R2236 B.n1075 B.n9 163.367
R2237 B.n1071 B.n9 163.367
R2238 B.n1071 B.n11 163.367
R2239 B.n1067 B.n11 163.367
R2240 B.n1067 B.n17 163.367
R2241 B.n1063 B.n17 163.367
R2242 B.n1063 B.n19 163.367
R2243 B.n1059 B.n19 163.367
R2244 B.n1059 B.n24 163.367
R2245 B.n1055 B.n24 163.367
R2246 B.n1055 B.n26 163.367
R2247 B.n1051 B.n26 163.367
R2248 B.n1051 B.n31 163.367
R2249 B.n1047 B.n31 163.367
R2250 B.n1047 B.n33 163.367
R2251 B.n1043 B.n33 163.367
R2252 B.n1043 B.n38 163.367
R2253 B.n1039 B.n38 163.367
R2254 B.n1039 B.n40 163.367
R2255 B.n1035 B.n40 163.367
R2256 B.n1035 B.n45 163.367
R2257 B.n1031 B.n45 163.367
R2258 B.n1031 B.n47 163.367
R2259 B.n1027 B.n47 163.367
R2260 B.n1027 B.n52 163.367
R2261 B.n1023 B.n52 163.367
R2262 B.n1023 B.n54 163.367
R2263 B.n1019 B.n54 163.367
R2264 B.n1019 B.n59 163.367
R2265 B.n1015 B.n59 163.367
R2266 B.n1015 B.n61 163.367
R2267 B.n1011 B.n61 163.367
R2268 B.n1011 B.n66 163.367
R2269 B.n1007 B.n66 163.367
R2270 B.n1007 B.n68 163.367
R2271 B.n1003 B.n68 163.367
R2272 B.n1003 B.n73 163.367
R2273 B.n999 B.n73 163.367
R2274 B.n999 B.n75 163.367
R2275 B.n995 B.n75 163.367
R2276 B.n995 B.n80 163.367
R2277 B.n991 B.n80 163.367
R2278 B.n991 B.n82 163.367
R2279 B.n987 B.n82 163.367
R2280 B.n987 B.n87 163.367
R2281 B.n983 B.n982 71.676
R2282 B.n155 B.n90 71.676
R2283 B.n159 B.n91 71.676
R2284 B.n163 B.n92 71.676
R2285 B.n167 B.n93 71.676
R2286 B.n171 B.n94 71.676
R2287 B.n175 B.n95 71.676
R2288 B.n179 B.n96 71.676
R2289 B.n183 B.n97 71.676
R2290 B.n187 B.n98 71.676
R2291 B.n191 B.n99 71.676
R2292 B.n195 B.n100 71.676
R2293 B.n199 B.n101 71.676
R2294 B.n203 B.n102 71.676
R2295 B.n207 B.n103 71.676
R2296 B.n211 B.n104 71.676
R2297 B.n215 B.n105 71.676
R2298 B.n219 B.n106 71.676
R2299 B.n223 B.n107 71.676
R2300 B.n227 B.n108 71.676
R2301 B.n231 B.n109 71.676
R2302 B.n235 B.n110 71.676
R2303 B.n239 B.n111 71.676
R2304 B.n243 B.n112 71.676
R2305 B.n247 B.n113 71.676
R2306 B.n251 B.n114 71.676
R2307 B.n255 B.n115 71.676
R2308 B.n259 B.n116 71.676
R2309 B.n263 B.n117 71.676
R2310 B.n267 B.n118 71.676
R2311 B.n271 B.n119 71.676
R2312 B.n275 B.n120 71.676
R2313 B.n279 B.n121 71.676
R2314 B.n283 B.n122 71.676
R2315 B.n287 B.n123 71.676
R2316 B.n291 B.n124 71.676
R2317 B.n295 B.n125 71.676
R2318 B.n299 B.n126 71.676
R2319 B.n303 B.n127 71.676
R2320 B.n307 B.n128 71.676
R2321 B.n311 B.n129 71.676
R2322 B.n315 B.n130 71.676
R2323 B.n319 B.n131 71.676
R2324 B.n323 B.n132 71.676
R2325 B.n327 B.n133 71.676
R2326 B.n331 B.n134 71.676
R2327 B.n335 B.n135 71.676
R2328 B.n339 B.n136 71.676
R2329 B.n343 B.n137 71.676
R2330 B.n347 B.n138 71.676
R2331 B.n351 B.n139 71.676
R2332 B.n355 B.n140 71.676
R2333 B.n359 B.n141 71.676
R2334 B.n363 B.n142 71.676
R2335 B.n367 B.n143 71.676
R2336 B.n371 B.n144 71.676
R2337 B.n375 B.n145 71.676
R2338 B.n379 B.n146 71.676
R2339 B.n980 B.n147 71.676
R2340 B.n980 B.n979 71.676
R2341 B.n381 B.n146 71.676
R2342 B.n378 B.n145 71.676
R2343 B.n374 B.n144 71.676
R2344 B.n370 B.n143 71.676
R2345 B.n366 B.n142 71.676
R2346 B.n362 B.n141 71.676
R2347 B.n358 B.n140 71.676
R2348 B.n354 B.n139 71.676
R2349 B.n350 B.n138 71.676
R2350 B.n346 B.n137 71.676
R2351 B.n342 B.n136 71.676
R2352 B.n338 B.n135 71.676
R2353 B.n334 B.n134 71.676
R2354 B.n330 B.n133 71.676
R2355 B.n326 B.n132 71.676
R2356 B.n322 B.n131 71.676
R2357 B.n318 B.n130 71.676
R2358 B.n314 B.n129 71.676
R2359 B.n310 B.n128 71.676
R2360 B.n306 B.n127 71.676
R2361 B.n302 B.n126 71.676
R2362 B.n298 B.n125 71.676
R2363 B.n294 B.n124 71.676
R2364 B.n290 B.n123 71.676
R2365 B.n286 B.n122 71.676
R2366 B.n282 B.n121 71.676
R2367 B.n278 B.n120 71.676
R2368 B.n274 B.n119 71.676
R2369 B.n270 B.n118 71.676
R2370 B.n266 B.n117 71.676
R2371 B.n262 B.n116 71.676
R2372 B.n258 B.n115 71.676
R2373 B.n254 B.n114 71.676
R2374 B.n250 B.n113 71.676
R2375 B.n246 B.n112 71.676
R2376 B.n242 B.n111 71.676
R2377 B.n238 B.n110 71.676
R2378 B.n234 B.n109 71.676
R2379 B.n230 B.n108 71.676
R2380 B.n226 B.n107 71.676
R2381 B.n222 B.n106 71.676
R2382 B.n218 B.n105 71.676
R2383 B.n214 B.n104 71.676
R2384 B.n210 B.n103 71.676
R2385 B.n206 B.n102 71.676
R2386 B.n202 B.n101 71.676
R2387 B.n198 B.n100 71.676
R2388 B.n194 B.n99 71.676
R2389 B.n190 B.n98 71.676
R2390 B.n186 B.n97 71.676
R2391 B.n182 B.n96 71.676
R2392 B.n178 B.n95 71.676
R2393 B.n174 B.n94 71.676
R2394 B.n170 B.n93 71.676
R2395 B.n166 B.n92 71.676
R2396 B.n162 B.n91 71.676
R2397 B.n158 B.n90 71.676
R2398 B.n982 B.n89 71.676
R2399 B.n775 B.n774 71.676
R2400 B.n536 B.n478 71.676
R2401 B.n767 B.n479 71.676
R2402 B.n763 B.n480 71.676
R2403 B.n759 B.n481 71.676
R2404 B.n755 B.n482 71.676
R2405 B.n751 B.n483 71.676
R2406 B.n747 B.n484 71.676
R2407 B.n743 B.n485 71.676
R2408 B.n739 B.n486 71.676
R2409 B.n735 B.n487 71.676
R2410 B.n731 B.n488 71.676
R2411 B.n727 B.n489 71.676
R2412 B.n723 B.n490 71.676
R2413 B.n719 B.n491 71.676
R2414 B.n715 B.n492 71.676
R2415 B.n711 B.n493 71.676
R2416 B.n707 B.n494 71.676
R2417 B.n703 B.n495 71.676
R2418 B.n699 B.n496 71.676
R2419 B.n695 B.n497 71.676
R2420 B.n691 B.n498 71.676
R2421 B.n687 B.n499 71.676
R2422 B.n683 B.n500 71.676
R2423 B.n679 B.n501 71.676
R2424 B.n675 B.n502 71.676
R2425 B.n671 B.n503 71.676
R2426 B.n666 B.n504 71.676
R2427 B.n662 B.n505 71.676
R2428 B.n658 B.n506 71.676
R2429 B.n654 B.n507 71.676
R2430 B.n650 B.n508 71.676
R2431 B.n645 B.n509 71.676
R2432 B.n641 B.n510 71.676
R2433 B.n637 B.n511 71.676
R2434 B.n633 B.n512 71.676
R2435 B.n629 B.n513 71.676
R2436 B.n625 B.n514 71.676
R2437 B.n621 B.n515 71.676
R2438 B.n617 B.n516 71.676
R2439 B.n613 B.n517 71.676
R2440 B.n609 B.n518 71.676
R2441 B.n605 B.n519 71.676
R2442 B.n601 B.n520 71.676
R2443 B.n597 B.n521 71.676
R2444 B.n593 B.n522 71.676
R2445 B.n589 B.n523 71.676
R2446 B.n585 B.n524 71.676
R2447 B.n581 B.n525 71.676
R2448 B.n577 B.n526 71.676
R2449 B.n573 B.n527 71.676
R2450 B.n569 B.n528 71.676
R2451 B.n565 B.n529 71.676
R2452 B.n561 B.n530 71.676
R2453 B.n557 B.n531 71.676
R2454 B.n553 B.n532 71.676
R2455 B.n549 B.n533 71.676
R2456 B.n545 B.n534 71.676
R2457 B.n774 B.n477 71.676
R2458 B.n768 B.n478 71.676
R2459 B.n764 B.n479 71.676
R2460 B.n760 B.n480 71.676
R2461 B.n756 B.n481 71.676
R2462 B.n752 B.n482 71.676
R2463 B.n748 B.n483 71.676
R2464 B.n744 B.n484 71.676
R2465 B.n740 B.n485 71.676
R2466 B.n736 B.n486 71.676
R2467 B.n732 B.n487 71.676
R2468 B.n728 B.n488 71.676
R2469 B.n724 B.n489 71.676
R2470 B.n720 B.n490 71.676
R2471 B.n716 B.n491 71.676
R2472 B.n712 B.n492 71.676
R2473 B.n708 B.n493 71.676
R2474 B.n704 B.n494 71.676
R2475 B.n700 B.n495 71.676
R2476 B.n696 B.n496 71.676
R2477 B.n692 B.n497 71.676
R2478 B.n688 B.n498 71.676
R2479 B.n684 B.n499 71.676
R2480 B.n680 B.n500 71.676
R2481 B.n676 B.n501 71.676
R2482 B.n672 B.n502 71.676
R2483 B.n667 B.n503 71.676
R2484 B.n663 B.n504 71.676
R2485 B.n659 B.n505 71.676
R2486 B.n655 B.n506 71.676
R2487 B.n651 B.n507 71.676
R2488 B.n646 B.n508 71.676
R2489 B.n642 B.n509 71.676
R2490 B.n638 B.n510 71.676
R2491 B.n634 B.n511 71.676
R2492 B.n630 B.n512 71.676
R2493 B.n626 B.n513 71.676
R2494 B.n622 B.n514 71.676
R2495 B.n618 B.n515 71.676
R2496 B.n614 B.n516 71.676
R2497 B.n610 B.n517 71.676
R2498 B.n606 B.n518 71.676
R2499 B.n602 B.n519 71.676
R2500 B.n598 B.n520 71.676
R2501 B.n594 B.n521 71.676
R2502 B.n590 B.n522 71.676
R2503 B.n586 B.n523 71.676
R2504 B.n582 B.n524 71.676
R2505 B.n578 B.n525 71.676
R2506 B.n574 B.n526 71.676
R2507 B.n570 B.n527 71.676
R2508 B.n566 B.n528 71.676
R2509 B.n562 B.n529 71.676
R2510 B.n558 B.n530 71.676
R2511 B.n554 B.n531 71.676
R2512 B.n550 B.n532 71.676
R2513 B.n546 B.n533 71.676
R2514 B.n542 B.n534 71.676
R2515 B.n1081 B.n1080 71.676
R2516 B.n1081 B.n2 71.676
R2517 B.n773 B.n474 63.8204
R2518 B.n981 B.n86 63.8204
R2519 B.n154 B.n153 59.5399
R2520 B.n151 B.n150 59.5399
R2521 B.n648 B.n540 59.5399
R2522 B.n669 B.n538 59.5399
R2523 B.n153 B.n152 51.9763
R2524 B.n150 B.n149 51.9763
R2525 B.n540 B.n539 51.9763
R2526 B.n538 B.n537 51.9763
R2527 B.n780 B.n474 34.7185
R2528 B.n780 B.n470 34.7185
R2529 B.n786 B.n470 34.7185
R2530 B.n786 B.n466 34.7185
R2531 B.n792 B.n466 34.7185
R2532 B.n792 B.n462 34.7185
R2533 B.n798 B.n462 34.7185
R2534 B.n804 B.n458 34.7185
R2535 B.n804 B.n454 34.7185
R2536 B.n810 B.n454 34.7185
R2537 B.n810 B.n450 34.7185
R2538 B.n816 B.n450 34.7185
R2539 B.n816 B.n446 34.7185
R2540 B.n822 B.n446 34.7185
R2541 B.n822 B.n441 34.7185
R2542 B.n828 B.n441 34.7185
R2543 B.n828 B.n442 34.7185
R2544 B.n834 B.n434 34.7185
R2545 B.n840 B.n434 34.7185
R2546 B.n840 B.n430 34.7185
R2547 B.n846 B.n430 34.7185
R2548 B.n846 B.n425 34.7185
R2549 B.n852 B.n425 34.7185
R2550 B.n852 B.n426 34.7185
R2551 B.n858 B.n418 34.7185
R2552 B.n864 B.n418 34.7185
R2553 B.n864 B.n414 34.7185
R2554 B.n870 B.n414 34.7185
R2555 B.n870 B.n409 34.7185
R2556 B.n876 B.n409 34.7185
R2557 B.n876 B.n410 34.7185
R2558 B.n882 B.n402 34.7185
R2559 B.n888 B.n402 34.7185
R2560 B.n888 B.n398 34.7185
R2561 B.n894 B.n398 34.7185
R2562 B.n894 B.n394 34.7185
R2563 B.n900 B.n394 34.7185
R2564 B.n907 B.n390 34.7185
R2565 B.n907 B.n386 34.7185
R2566 B.n913 B.n386 34.7185
R2567 B.n913 B.n4 34.7185
R2568 B.n1079 B.n4 34.7185
R2569 B.n1079 B.n1078 34.7185
R2570 B.n1078 B.n1077 34.7185
R2571 B.n1077 B.n8 34.7185
R2572 B.n12 B.n8 34.7185
R2573 B.n1070 B.n12 34.7185
R2574 B.n1070 B.n1069 34.7185
R2575 B.n1068 B.n16 34.7185
R2576 B.n1062 B.n16 34.7185
R2577 B.n1062 B.n1061 34.7185
R2578 B.n1061 B.n1060 34.7185
R2579 B.n1060 B.n23 34.7185
R2580 B.n1054 B.n23 34.7185
R2581 B.n1053 B.n1052 34.7185
R2582 B.n1052 B.n30 34.7185
R2583 B.n1046 B.n30 34.7185
R2584 B.n1046 B.n1045 34.7185
R2585 B.n1045 B.n1044 34.7185
R2586 B.n1044 B.n37 34.7185
R2587 B.n1038 B.n37 34.7185
R2588 B.n1037 B.n1036 34.7185
R2589 B.n1036 B.n44 34.7185
R2590 B.n1030 B.n44 34.7185
R2591 B.n1030 B.n1029 34.7185
R2592 B.n1029 B.n1028 34.7185
R2593 B.n1028 B.n51 34.7185
R2594 B.n1022 B.n51 34.7185
R2595 B.n1021 B.n1020 34.7185
R2596 B.n1020 B.n58 34.7185
R2597 B.n1014 B.n58 34.7185
R2598 B.n1014 B.n1013 34.7185
R2599 B.n1013 B.n1012 34.7185
R2600 B.n1012 B.n65 34.7185
R2601 B.n1006 B.n65 34.7185
R2602 B.n1006 B.n1005 34.7185
R2603 B.n1005 B.n1004 34.7185
R2604 B.n1004 B.n72 34.7185
R2605 B.n998 B.n997 34.7185
R2606 B.n997 B.n996 34.7185
R2607 B.n996 B.n79 34.7185
R2608 B.n990 B.n79 34.7185
R2609 B.n990 B.n989 34.7185
R2610 B.n989 B.n988 34.7185
R2611 B.n988 B.n86 34.7185
R2612 B.n900 B.t0 33.1869
R2613 B.t1 B.n1068 33.1869
R2614 B.n777 B.n776 32.3127
R2615 B.n541 B.n472 32.3127
R2616 B.n978 B.n977 32.3127
R2617 B.n985 B.n984 32.3127
R2618 B.n882 B.t7 32.1657
R2619 B.n1054 B.t4 32.1657
R2620 B.n858 B.t5 28.0813
R2621 B.n1038 B.t2 28.0813
R2622 B.t9 B.n458 27.0601
R2623 B.t13 B.n72 27.0601
R2624 B.n834 B.t6 23.9968
R2625 B.n1022 B.t3 23.9968
R2626 B B.n1082 18.0485
R2627 B.n442 B.t6 10.7222
R2628 B.t3 B.n1021 10.7222
R2629 B.n778 B.n777 10.6151
R2630 B.n778 B.n468 10.6151
R2631 B.n788 B.n468 10.6151
R2632 B.n789 B.n788 10.6151
R2633 B.n790 B.n789 10.6151
R2634 B.n790 B.n460 10.6151
R2635 B.n800 B.n460 10.6151
R2636 B.n801 B.n800 10.6151
R2637 B.n802 B.n801 10.6151
R2638 B.n802 B.n452 10.6151
R2639 B.n812 B.n452 10.6151
R2640 B.n813 B.n812 10.6151
R2641 B.n814 B.n813 10.6151
R2642 B.n814 B.n444 10.6151
R2643 B.n824 B.n444 10.6151
R2644 B.n825 B.n824 10.6151
R2645 B.n826 B.n825 10.6151
R2646 B.n826 B.n436 10.6151
R2647 B.n836 B.n436 10.6151
R2648 B.n837 B.n836 10.6151
R2649 B.n838 B.n837 10.6151
R2650 B.n838 B.n428 10.6151
R2651 B.n848 B.n428 10.6151
R2652 B.n849 B.n848 10.6151
R2653 B.n850 B.n849 10.6151
R2654 B.n850 B.n420 10.6151
R2655 B.n860 B.n420 10.6151
R2656 B.n861 B.n860 10.6151
R2657 B.n862 B.n861 10.6151
R2658 B.n862 B.n412 10.6151
R2659 B.n872 B.n412 10.6151
R2660 B.n873 B.n872 10.6151
R2661 B.n874 B.n873 10.6151
R2662 B.n874 B.n404 10.6151
R2663 B.n884 B.n404 10.6151
R2664 B.n885 B.n884 10.6151
R2665 B.n886 B.n885 10.6151
R2666 B.n886 B.n396 10.6151
R2667 B.n896 B.n396 10.6151
R2668 B.n897 B.n896 10.6151
R2669 B.n898 B.n897 10.6151
R2670 B.n898 B.n388 10.6151
R2671 B.n909 B.n388 10.6151
R2672 B.n910 B.n909 10.6151
R2673 B.n911 B.n910 10.6151
R2674 B.n911 B.n0 10.6151
R2675 B.n776 B.n476 10.6151
R2676 B.n771 B.n476 10.6151
R2677 B.n771 B.n770 10.6151
R2678 B.n770 B.n769 10.6151
R2679 B.n769 B.n766 10.6151
R2680 B.n766 B.n765 10.6151
R2681 B.n765 B.n762 10.6151
R2682 B.n762 B.n761 10.6151
R2683 B.n761 B.n758 10.6151
R2684 B.n758 B.n757 10.6151
R2685 B.n757 B.n754 10.6151
R2686 B.n754 B.n753 10.6151
R2687 B.n753 B.n750 10.6151
R2688 B.n750 B.n749 10.6151
R2689 B.n749 B.n746 10.6151
R2690 B.n746 B.n745 10.6151
R2691 B.n745 B.n742 10.6151
R2692 B.n742 B.n741 10.6151
R2693 B.n741 B.n738 10.6151
R2694 B.n738 B.n737 10.6151
R2695 B.n737 B.n734 10.6151
R2696 B.n734 B.n733 10.6151
R2697 B.n733 B.n730 10.6151
R2698 B.n730 B.n729 10.6151
R2699 B.n729 B.n726 10.6151
R2700 B.n726 B.n725 10.6151
R2701 B.n725 B.n722 10.6151
R2702 B.n722 B.n721 10.6151
R2703 B.n721 B.n718 10.6151
R2704 B.n718 B.n717 10.6151
R2705 B.n717 B.n714 10.6151
R2706 B.n714 B.n713 10.6151
R2707 B.n713 B.n710 10.6151
R2708 B.n710 B.n709 10.6151
R2709 B.n709 B.n706 10.6151
R2710 B.n706 B.n705 10.6151
R2711 B.n705 B.n702 10.6151
R2712 B.n702 B.n701 10.6151
R2713 B.n701 B.n698 10.6151
R2714 B.n698 B.n697 10.6151
R2715 B.n697 B.n694 10.6151
R2716 B.n694 B.n693 10.6151
R2717 B.n693 B.n690 10.6151
R2718 B.n690 B.n689 10.6151
R2719 B.n689 B.n686 10.6151
R2720 B.n686 B.n685 10.6151
R2721 B.n685 B.n682 10.6151
R2722 B.n682 B.n681 10.6151
R2723 B.n681 B.n678 10.6151
R2724 B.n678 B.n677 10.6151
R2725 B.n677 B.n674 10.6151
R2726 B.n674 B.n673 10.6151
R2727 B.n673 B.n670 10.6151
R2728 B.n668 B.n665 10.6151
R2729 B.n665 B.n664 10.6151
R2730 B.n664 B.n661 10.6151
R2731 B.n661 B.n660 10.6151
R2732 B.n660 B.n657 10.6151
R2733 B.n657 B.n656 10.6151
R2734 B.n656 B.n653 10.6151
R2735 B.n653 B.n652 10.6151
R2736 B.n652 B.n649 10.6151
R2737 B.n647 B.n644 10.6151
R2738 B.n644 B.n643 10.6151
R2739 B.n643 B.n640 10.6151
R2740 B.n640 B.n639 10.6151
R2741 B.n639 B.n636 10.6151
R2742 B.n636 B.n635 10.6151
R2743 B.n635 B.n632 10.6151
R2744 B.n632 B.n631 10.6151
R2745 B.n631 B.n628 10.6151
R2746 B.n628 B.n627 10.6151
R2747 B.n627 B.n624 10.6151
R2748 B.n624 B.n623 10.6151
R2749 B.n623 B.n620 10.6151
R2750 B.n620 B.n619 10.6151
R2751 B.n619 B.n616 10.6151
R2752 B.n616 B.n615 10.6151
R2753 B.n615 B.n612 10.6151
R2754 B.n612 B.n611 10.6151
R2755 B.n611 B.n608 10.6151
R2756 B.n608 B.n607 10.6151
R2757 B.n607 B.n604 10.6151
R2758 B.n604 B.n603 10.6151
R2759 B.n603 B.n600 10.6151
R2760 B.n600 B.n599 10.6151
R2761 B.n599 B.n596 10.6151
R2762 B.n596 B.n595 10.6151
R2763 B.n595 B.n592 10.6151
R2764 B.n592 B.n591 10.6151
R2765 B.n591 B.n588 10.6151
R2766 B.n588 B.n587 10.6151
R2767 B.n587 B.n584 10.6151
R2768 B.n584 B.n583 10.6151
R2769 B.n583 B.n580 10.6151
R2770 B.n580 B.n579 10.6151
R2771 B.n579 B.n576 10.6151
R2772 B.n576 B.n575 10.6151
R2773 B.n575 B.n572 10.6151
R2774 B.n572 B.n571 10.6151
R2775 B.n571 B.n568 10.6151
R2776 B.n568 B.n567 10.6151
R2777 B.n567 B.n564 10.6151
R2778 B.n564 B.n563 10.6151
R2779 B.n563 B.n560 10.6151
R2780 B.n560 B.n559 10.6151
R2781 B.n559 B.n556 10.6151
R2782 B.n556 B.n555 10.6151
R2783 B.n555 B.n552 10.6151
R2784 B.n552 B.n551 10.6151
R2785 B.n551 B.n548 10.6151
R2786 B.n548 B.n547 10.6151
R2787 B.n547 B.n544 10.6151
R2788 B.n544 B.n543 10.6151
R2789 B.n543 B.n541 10.6151
R2790 B.n782 B.n472 10.6151
R2791 B.n783 B.n782 10.6151
R2792 B.n784 B.n783 10.6151
R2793 B.n784 B.n464 10.6151
R2794 B.n794 B.n464 10.6151
R2795 B.n795 B.n794 10.6151
R2796 B.n796 B.n795 10.6151
R2797 B.n796 B.n456 10.6151
R2798 B.n806 B.n456 10.6151
R2799 B.n807 B.n806 10.6151
R2800 B.n808 B.n807 10.6151
R2801 B.n808 B.n448 10.6151
R2802 B.n818 B.n448 10.6151
R2803 B.n819 B.n818 10.6151
R2804 B.n820 B.n819 10.6151
R2805 B.n820 B.n439 10.6151
R2806 B.n830 B.n439 10.6151
R2807 B.n831 B.n830 10.6151
R2808 B.n832 B.n831 10.6151
R2809 B.n832 B.n432 10.6151
R2810 B.n842 B.n432 10.6151
R2811 B.n843 B.n842 10.6151
R2812 B.n844 B.n843 10.6151
R2813 B.n844 B.n423 10.6151
R2814 B.n854 B.n423 10.6151
R2815 B.n855 B.n854 10.6151
R2816 B.n856 B.n855 10.6151
R2817 B.n856 B.n416 10.6151
R2818 B.n866 B.n416 10.6151
R2819 B.n867 B.n866 10.6151
R2820 B.n868 B.n867 10.6151
R2821 B.n868 B.n407 10.6151
R2822 B.n878 B.n407 10.6151
R2823 B.n879 B.n878 10.6151
R2824 B.n880 B.n879 10.6151
R2825 B.n880 B.n400 10.6151
R2826 B.n890 B.n400 10.6151
R2827 B.n891 B.n890 10.6151
R2828 B.n892 B.n891 10.6151
R2829 B.n892 B.n392 10.6151
R2830 B.n902 B.n392 10.6151
R2831 B.n903 B.n902 10.6151
R2832 B.n905 B.n903 10.6151
R2833 B.n905 B.n904 10.6151
R2834 B.n904 B.n384 10.6151
R2835 B.n916 B.n384 10.6151
R2836 B.n917 B.n916 10.6151
R2837 B.n918 B.n917 10.6151
R2838 B.n919 B.n918 10.6151
R2839 B.n920 B.n919 10.6151
R2840 B.n923 B.n920 10.6151
R2841 B.n924 B.n923 10.6151
R2842 B.n925 B.n924 10.6151
R2843 B.n926 B.n925 10.6151
R2844 B.n928 B.n926 10.6151
R2845 B.n929 B.n928 10.6151
R2846 B.n930 B.n929 10.6151
R2847 B.n931 B.n930 10.6151
R2848 B.n933 B.n931 10.6151
R2849 B.n934 B.n933 10.6151
R2850 B.n935 B.n934 10.6151
R2851 B.n936 B.n935 10.6151
R2852 B.n938 B.n936 10.6151
R2853 B.n939 B.n938 10.6151
R2854 B.n940 B.n939 10.6151
R2855 B.n941 B.n940 10.6151
R2856 B.n943 B.n941 10.6151
R2857 B.n944 B.n943 10.6151
R2858 B.n945 B.n944 10.6151
R2859 B.n946 B.n945 10.6151
R2860 B.n948 B.n946 10.6151
R2861 B.n949 B.n948 10.6151
R2862 B.n950 B.n949 10.6151
R2863 B.n951 B.n950 10.6151
R2864 B.n953 B.n951 10.6151
R2865 B.n954 B.n953 10.6151
R2866 B.n955 B.n954 10.6151
R2867 B.n956 B.n955 10.6151
R2868 B.n958 B.n956 10.6151
R2869 B.n959 B.n958 10.6151
R2870 B.n960 B.n959 10.6151
R2871 B.n961 B.n960 10.6151
R2872 B.n963 B.n961 10.6151
R2873 B.n964 B.n963 10.6151
R2874 B.n965 B.n964 10.6151
R2875 B.n966 B.n965 10.6151
R2876 B.n968 B.n966 10.6151
R2877 B.n969 B.n968 10.6151
R2878 B.n970 B.n969 10.6151
R2879 B.n971 B.n970 10.6151
R2880 B.n973 B.n971 10.6151
R2881 B.n974 B.n973 10.6151
R2882 B.n975 B.n974 10.6151
R2883 B.n976 B.n975 10.6151
R2884 B.n977 B.n976 10.6151
R2885 B.n1074 B.n1 10.6151
R2886 B.n1074 B.n1073 10.6151
R2887 B.n1073 B.n1072 10.6151
R2888 B.n1072 B.n10 10.6151
R2889 B.n1066 B.n10 10.6151
R2890 B.n1066 B.n1065 10.6151
R2891 B.n1065 B.n1064 10.6151
R2892 B.n1064 B.n18 10.6151
R2893 B.n1058 B.n18 10.6151
R2894 B.n1058 B.n1057 10.6151
R2895 B.n1057 B.n1056 10.6151
R2896 B.n1056 B.n25 10.6151
R2897 B.n1050 B.n25 10.6151
R2898 B.n1050 B.n1049 10.6151
R2899 B.n1049 B.n1048 10.6151
R2900 B.n1048 B.n32 10.6151
R2901 B.n1042 B.n32 10.6151
R2902 B.n1042 B.n1041 10.6151
R2903 B.n1041 B.n1040 10.6151
R2904 B.n1040 B.n39 10.6151
R2905 B.n1034 B.n39 10.6151
R2906 B.n1034 B.n1033 10.6151
R2907 B.n1033 B.n1032 10.6151
R2908 B.n1032 B.n46 10.6151
R2909 B.n1026 B.n46 10.6151
R2910 B.n1026 B.n1025 10.6151
R2911 B.n1025 B.n1024 10.6151
R2912 B.n1024 B.n53 10.6151
R2913 B.n1018 B.n53 10.6151
R2914 B.n1018 B.n1017 10.6151
R2915 B.n1017 B.n1016 10.6151
R2916 B.n1016 B.n60 10.6151
R2917 B.n1010 B.n60 10.6151
R2918 B.n1010 B.n1009 10.6151
R2919 B.n1009 B.n1008 10.6151
R2920 B.n1008 B.n67 10.6151
R2921 B.n1002 B.n67 10.6151
R2922 B.n1002 B.n1001 10.6151
R2923 B.n1001 B.n1000 10.6151
R2924 B.n1000 B.n74 10.6151
R2925 B.n994 B.n74 10.6151
R2926 B.n994 B.n993 10.6151
R2927 B.n993 B.n992 10.6151
R2928 B.n992 B.n81 10.6151
R2929 B.n986 B.n81 10.6151
R2930 B.n986 B.n985 10.6151
R2931 B.n984 B.n88 10.6151
R2932 B.n156 B.n88 10.6151
R2933 B.n157 B.n156 10.6151
R2934 B.n160 B.n157 10.6151
R2935 B.n161 B.n160 10.6151
R2936 B.n164 B.n161 10.6151
R2937 B.n165 B.n164 10.6151
R2938 B.n168 B.n165 10.6151
R2939 B.n169 B.n168 10.6151
R2940 B.n172 B.n169 10.6151
R2941 B.n173 B.n172 10.6151
R2942 B.n176 B.n173 10.6151
R2943 B.n177 B.n176 10.6151
R2944 B.n180 B.n177 10.6151
R2945 B.n181 B.n180 10.6151
R2946 B.n184 B.n181 10.6151
R2947 B.n185 B.n184 10.6151
R2948 B.n188 B.n185 10.6151
R2949 B.n189 B.n188 10.6151
R2950 B.n192 B.n189 10.6151
R2951 B.n193 B.n192 10.6151
R2952 B.n196 B.n193 10.6151
R2953 B.n197 B.n196 10.6151
R2954 B.n200 B.n197 10.6151
R2955 B.n201 B.n200 10.6151
R2956 B.n204 B.n201 10.6151
R2957 B.n205 B.n204 10.6151
R2958 B.n208 B.n205 10.6151
R2959 B.n209 B.n208 10.6151
R2960 B.n212 B.n209 10.6151
R2961 B.n213 B.n212 10.6151
R2962 B.n216 B.n213 10.6151
R2963 B.n217 B.n216 10.6151
R2964 B.n220 B.n217 10.6151
R2965 B.n221 B.n220 10.6151
R2966 B.n224 B.n221 10.6151
R2967 B.n225 B.n224 10.6151
R2968 B.n228 B.n225 10.6151
R2969 B.n229 B.n228 10.6151
R2970 B.n232 B.n229 10.6151
R2971 B.n233 B.n232 10.6151
R2972 B.n236 B.n233 10.6151
R2973 B.n237 B.n236 10.6151
R2974 B.n240 B.n237 10.6151
R2975 B.n241 B.n240 10.6151
R2976 B.n244 B.n241 10.6151
R2977 B.n245 B.n244 10.6151
R2978 B.n248 B.n245 10.6151
R2979 B.n249 B.n248 10.6151
R2980 B.n252 B.n249 10.6151
R2981 B.n253 B.n252 10.6151
R2982 B.n256 B.n253 10.6151
R2983 B.n257 B.n256 10.6151
R2984 B.n261 B.n260 10.6151
R2985 B.n264 B.n261 10.6151
R2986 B.n265 B.n264 10.6151
R2987 B.n268 B.n265 10.6151
R2988 B.n269 B.n268 10.6151
R2989 B.n272 B.n269 10.6151
R2990 B.n273 B.n272 10.6151
R2991 B.n276 B.n273 10.6151
R2992 B.n277 B.n276 10.6151
R2993 B.n281 B.n280 10.6151
R2994 B.n284 B.n281 10.6151
R2995 B.n285 B.n284 10.6151
R2996 B.n288 B.n285 10.6151
R2997 B.n289 B.n288 10.6151
R2998 B.n292 B.n289 10.6151
R2999 B.n293 B.n292 10.6151
R3000 B.n296 B.n293 10.6151
R3001 B.n297 B.n296 10.6151
R3002 B.n300 B.n297 10.6151
R3003 B.n301 B.n300 10.6151
R3004 B.n304 B.n301 10.6151
R3005 B.n305 B.n304 10.6151
R3006 B.n308 B.n305 10.6151
R3007 B.n309 B.n308 10.6151
R3008 B.n312 B.n309 10.6151
R3009 B.n313 B.n312 10.6151
R3010 B.n316 B.n313 10.6151
R3011 B.n317 B.n316 10.6151
R3012 B.n320 B.n317 10.6151
R3013 B.n321 B.n320 10.6151
R3014 B.n324 B.n321 10.6151
R3015 B.n325 B.n324 10.6151
R3016 B.n328 B.n325 10.6151
R3017 B.n329 B.n328 10.6151
R3018 B.n332 B.n329 10.6151
R3019 B.n333 B.n332 10.6151
R3020 B.n336 B.n333 10.6151
R3021 B.n337 B.n336 10.6151
R3022 B.n340 B.n337 10.6151
R3023 B.n341 B.n340 10.6151
R3024 B.n344 B.n341 10.6151
R3025 B.n345 B.n344 10.6151
R3026 B.n348 B.n345 10.6151
R3027 B.n349 B.n348 10.6151
R3028 B.n352 B.n349 10.6151
R3029 B.n353 B.n352 10.6151
R3030 B.n356 B.n353 10.6151
R3031 B.n357 B.n356 10.6151
R3032 B.n360 B.n357 10.6151
R3033 B.n361 B.n360 10.6151
R3034 B.n364 B.n361 10.6151
R3035 B.n365 B.n364 10.6151
R3036 B.n368 B.n365 10.6151
R3037 B.n369 B.n368 10.6151
R3038 B.n372 B.n369 10.6151
R3039 B.n373 B.n372 10.6151
R3040 B.n376 B.n373 10.6151
R3041 B.n377 B.n376 10.6151
R3042 B.n380 B.n377 10.6151
R3043 B.n382 B.n380 10.6151
R3044 B.n383 B.n382 10.6151
R3045 B.n978 B.n383 10.6151
R3046 B.n670 B.n669 9.36635
R3047 B.n648 B.n647 9.36635
R3048 B.n257 B.n154 9.36635
R3049 B.n280 B.n151 9.36635
R3050 B.n1082 B.n0 8.11757
R3051 B.n1082 B.n1 8.11757
R3052 B.n798 B.t9 7.65889
R3053 B.n998 B.t13 7.65889
R3054 B.n426 B.t5 6.63777
R3055 B.t2 B.n1037 6.63777
R3056 B.n410 B.t7 2.5533
R3057 B.t4 B.n1053 2.5533
R3058 B.t0 B.n390 1.53218
R3059 B.n1069 B.t1 1.53218
R3060 B.n669 B.n668 1.24928
R3061 B.n649 B.n648 1.24928
R3062 B.n260 B.n154 1.24928
R3063 B.n277 B.n151 1.24928
R3064 VN.n7 VN.t6 198.825
R3065 VN.n34 VN.t3 198.825
R3066 VN.n6 VN.t5 166.855
R3067 VN.n17 VN.t4 166.855
R3068 VN.n25 VN.t7 166.855
R3069 VN.n33 VN.t1 166.855
R3070 VN.n44 VN.t2 166.855
R3071 VN.n52 VN.t0 166.855
R3072 VN.n51 VN.n27 161.3
R3073 VN.n50 VN.n49 161.3
R3074 VN.n48 VN.n28 161.3
R3075 VN.n47 VN.n46 161.3
R3076 VN.n45 VN.n29 161.3
R3077 VN.n43 VN.n42 161.3
R3078 VN.n41 VN.n30 161.3
R3079 VN.n40 VN.n39 161.3
R3080 VN.n38 VN.n31 161.3
R3081 VN.n37 VN.n36 161.3
R3082 VN.n35 VN.n32 161.3
R3083 VN.n24 VN.n0 161.3
R3084 VN.n23 VN.n22 161.3
R3085 VN.n21 VN.n1 161.3
R3086 VN.n20 VN.n19 161.3
R3087 VN.n18 VN.n2 161.3
R3088 VN.n16 VN.n15 161.3
R3089 VN.n14 VN.n3 161.3
R3090 VN.n13 VN.n12 161.3
R3091 VN.n11 VN.n4 161.3
R3092 VN.n10 VN.n9 161.3
R3093 VN.n8 VN.n5 161.3
R3094 VN.n26 VN.n25 97.5443
R3095 VN.n53 VN.n52 97.5443
R3096 VN.n7 VN.n6 67.7723
R3097 VN.n34 VN.n33 67.7723
R3098 VN.n12 VN.n11 56.5193
R3099 VN.n39 VN.n38 56.5193
R3100 VN VN.n53 53.2482
R3101 VN.n19 VN.n1 47.2923
R3102 VN.n46 VN.n28 47.2923
R3103 VN.n23 VN.n1 33.6945
R3104 VN.n50 VN.n28 33.6945
R3105 VN.n10 VN.n5 24.4675
R3106 VN.n11 VN.n10 24.4675
R3107 VN.n12 VN.n3 24.4675
R3108 VN.n16 VN.n3 24.4675
R3109 VN.n19 VN.n18 24.4675
R3110 VN.n24 VN.n23 24.4675
R3111 VN.n38 VN.n37 24.4675
R3112 VN.n37 VN.n32 24.4675
R3113 VN.n46 VN.n45 24.4675
R3114 VN.n43 VN.n30 24.4675
R3115 VN.n39 VN.n30 24.4675
R3116 VN.n51 VN.n50 24.4675
R3117 VN.n18 VN.n17 20.0634
R3118 VN.n45 VN.n44 20.0634
R3119 VN.n25 VN.n24 13.2127
R3120 VN.n52 VN.n51 13.2127
R3121 VN.n35 VN.n34 9.67836
R3122 VN.n8 VN.n7 9.67836
R3123 VN.n6 VN.n5 4.40456
R3124 VN.n17 VN.n16 4.40456
R3125 VN.n33 VN.n32 4.40456
R3126 VN.n44 VN.n43 4.40456
R3127 VN.n53 VN.n27 0.278367
R3128 VN.n26 VN.n0 0.278367
R3129 VN.n49 VN.n27 0.189894
R3130 VN.n49 VN.n48 0.189894
R3131 VN.n48 VN.n47 0.189894
R3132 VN.n47 VN.n29 0.189894
R3133 VN.n42 VN.n29 0.189894
R3134 VN.n42 VN.n41 0.189894
R3135 VN.n41 VN.n40 0.189894
R3136 VN.n40 VN.n31 0.189894
R3137 VN.n36 VN.n31 0.189894
R3138 VN.n36 VN.n35 0.189894
R3139 VN.n9 VN.n8 0.189894
R3140 VN.n9 VN.n4 0.189894
R3141 VN.n13 VN.n4 0.189894
R3142 VN.n14 VN.n13 0.189894
R3143 VN.n15 VN.n14 0.189894
R3144 VN.n15 VN.n2 0.189894
R3145 VN.n20 VN.n2 0.189894
R3146 VN.n21 VN.n20 0.189894
R3147 VN.n22 VN.n21 0.189894
R3148 VN.n22 VN.n0 0.189894
R3149 VN VN.n26 0.153454
R3150 VDD2.n2 VDD2.n1 65.5622
R3151 VDD2.n2 VDD2.n0 65.5622
R3152 VDD2 VDD2.n5 65.5594
R3153 VDD2.n4 VDD2.n3 64.4626
R3154 VDD2.n4 VDD2.n2 48.1377
R3155 VDD2.n5 VDD2.t6 1.21746
R3156 VDD2.n5 VDD2.t4 1.21746
R3157 VDD2.n3 VDD2.t7 1.21746
R3158 VDD2.n3 VDD2.t5 1.21746
R3159 VDD2.n1 VDD2.t3 1.21746
R3160 VDD2.n1 VDD2.t0 1.21746
R3161 VDD2.n0 VDD2.t1 1.21746
R3162 VDD2.n0 VDD2.t2 1.21746
R3163 VDD2 VDD2.n4 1.21386
C0 VP VDD2 0.492812f
C1 VN VDD2 11.3919f
C2 VP VTAIL 11.5275f
C3 VN VTAIL 11.5134f
C4 VP VDD1 11.732401f
C5 VN VDD1 0.151019f
C6 VTAIL VDD2 9.62312f
C7 VDD1 VDD2 1.6455f
C8 VP VN 8.14819f
C9 VTAIL VDD1 9.570379f
C10 VDD2 B 5.42854f
C11 VDD1 B 5.83759f
C12 VTAIL B 12.861473f
C13 VN B 14.92179f
C14 VP B 13.4f
C15 VDD2.t1 B 0.313674f
C16 VDD2.t2 B 0.313674f
C17 VDD2.n0 B 2.85746f
C18 VDD2.t3 B 0.313674f
C19 VDD2.t0 B 0.313674f
C20 VDD2.n1 B 2.85746f
C21 VDD2.n2 B 3.31297f
C22 VDD2.t7 B 0.313674f
C23 VDD2.t5 B 0.313674f
C24 VDD2.n3 B 2.84949f
C25 VDD2.n4 B 3.10719f
C26 VDD2.t6 B 0.313674f
C27 VDD2.t4 B 0.313674f
C28 VDD2.n5 B 2.85743f
C29 VN.n0 B 0.030134f
C30 VN.t7 B 2.3989f
C31 VN.n1 B 0.019957f
C32 VN.n2 B 0.022856f
C33 VN.t4 B 2.3989f
C34 VN.n3 B 0.042598f
C35 VN.n4 B 0.022856f
C36 VN.n5 B 0.025353f
C37 VN.t6 B 2.55408f
C38 VN.t5 B 2.3989f
C39 VN.n6 B 0.89314f
C40 VN.n7 B 0.888132f
C41 VN.n8 B 0.197987f
C42 VN.n9 B 0.022856f
C43 VN.n10 B 0.042598f
C44 VN.n11 B 0.033366f
C45 VN.n12 B 0.033366f
C46 VN.n13 B 0.022856f
C47 VN.n14 B 0.022856f
C48 VN.n15 B 0.022856f
C49 VN.n16 B 0.025353f
C50 VN.n17 B 0.837391f
C51 VN.n18 B 0.038813f
C52 VN.n19 B 0.043206f
C53 VN.n20 B 0.022856f
C54 VN.n21 B 0.022856f
C55 VN.n22 B 0.022856f
C56 VN.n23 B 0.046168f
C57 VN.n24 B 0.032924f
C58 VN.n25 B 0.910348f
C59 VN.n26 B 0.033615f
C60 VN.n27 B 0.030134f
C61 VN.t0 B 2.3989f
C62 VN.n28 B 0.019957f
C63 VN.n29 B 0.022856f
C64 VN.t2 B 2.3989f
C65 VN.n30 B 0.042598f
C66 VN.n31 B 0.022856f
C67 VN.n32 B 0.025353f
C68 VN.t3 B 2.55408f
C69 VN.t1 B 2.3989f
C70 VN.n33 B 0.89314f
C71 VN.n34 B 0.888132f
C72 VN.n35 B 0.197987f
C73 VN.n36 B 0.022856f
C74 VN.n37 B 0.042598f
C75 VN.n38 B 0.033366f
C76 VN.n39 B 0.033366f
C77 VN.n40 B 0.022856f
C78 VN.n41 B 0.022856f
C79 VN.n42 B 0.022856f
C80 VN.n43 B 0.025353f
C81 VN.n44 B 0.837391f
C82 VN.n45 B 0.038813f
C83 VN.n46 B 0.043206f
C84 VN.n47 B 0.022856f
C85 VN.n48 B 0.022856f
C86 VN.n49 B 0.022856f
C87 VN.n50 B 0.046168f
C88 VN.n51 B 0.032924f
C89 VN.n52 B 0.910348f
C90 VN.n53 B 1.39101f
C91 VTAIL.t4 B 0.240532f
C92 VTAIL.t2 B 0.240532f
C93 VTAIL.n0 B 2.1335f
C94 VTAIL.n1 B 0.32016f
C95 VTAIL.n2 B 0.02718f
C96 VTAIL.n3 B 0.018708f
C97 VTAIL.n4 B 0.010053f
C98 VTAIL.n5 B 0.023762f
C99 VTAIL.n6 B 0.010644f
C100 VTAIL.n7 B 0.018708f
C101 VTAIL.n8 B 0.010349f
C102 VTAIL.n9 B 0.023762f
C103 VTAIL.n10 B 0.010644f
C104 VTAIL.n11 B 0.018708f
C105 VTAIL.n12 B 0.010053f
C106 VTAIL.n13 B 0.023762f
C107 VTAIL.n14 B 0.010644f
C108 VTAIL.n15 B 0.018708f
C109 VTAIL.n16 B 0.010053f
C110 VTAIL.n17 B 0.023762f
C111 VTAIL.n18 B 0.010644f
C112 VTAIL.n19 B 0.018708f
C113 VTAIL.n20 B 0.010053f
C114 VTAIL.n21 B 0.023762f
C115 VTAIL.n22 B 0.010644f
C116 VTAIL.n23 B 0.018708f
C117 VTAIL.n24 B 0.010053f
C118 VTAIL.n25 B 0.023762f
C119 VTAIL.n26 B 0.010644f
C120 VTAIL.n27 B 0.018708f
C121 VTAIL.n28 B 0.010053f
C122 VTAIL.n29 B 0.017821f
C123 VTAIL.n30 B 0.014037f
C124 VTAIL.t1 B 0.039262f
C125 VTAIL.n31 B 0.127976f
C126 VTAIL.n32 B 1.32607f
C127 VTAIL.n33 B 0.010053f
C128 VTAIL.n34 B 0.010644f
C129 VTAIL.n35 B 0.023762f
C130 VTAIL.n36 B 0.023762f
C131 VTAIL.n37 B 0.010644f
C132 VTAIL.n38 B 0.010053f
C133 VTAIL.n39 B 0.018708f
C134 VTAIL.n40 B 0.018708f
C135 VTAIL.n41 B 0.010053f
C136 VTAIL.n42 B 0.010644f
C137 VTAIL.n43 B 0.023762f
C138 VTAIL.n44 B 0.023762f
C139 VTAIL.n45 B 0.010644f
C140 VTAIL.n46 B 0.010053f
C141 VTAIL.n47 B 0.018708f
C142 VTAIL.n48 B 0.018708f
C143 VTAIL.n49 B 0.010053f
C144 VTAIL.n50 B 0.010644f
C145 VTAIL.n51 B 0.023762f
C146 VTAIL.n52 B 0.023762f
C147 VTAIL.n53 B 0.010644f
C148 VTAIL.n54 B 0.010053f
C149 VTAIL.n55 B 0.018708f
C150 VTAIL.n56 B 0.018708f
C151 VTAIL.n57 B 0.010053f
C152 VTAIL.n58 B 0.010644f
C153 VTAIL.n59 B 0.023762f
C154 VTAIL.n60 B 0.023762f
C155 VTAIL.n61 B 0.010644f
C156 VTAIL.n62 B 0.010053f
C157 VTAIL.n63 B 0.018708f
C158 VTAIL.n64 B 0.018708f
C159 VTAIL.n65 B 0.010053f
C160 VTAIL.n66 B 0.010644f
C161 VTAIL.n67 B 0.023762f
C162 VTAIL.n68 B 0.023762f
C163 VTAIL.n69 B 0.010644f
C164 VTAIL.n70 B 0.010053f
C165 VTAIL.n71 B 0.018708f
C166 VTAIL.n72 B 0.018708f
C167 VTAIL.n73 B 0.010053f
C168 VTAIL.n74 B 0.010053f
C169 VTAIL.n75 B 0.010644f
C170 VTAIL.n76 B 0.023762f
C171 VTAIL.n77 B 0.023762f
C172 VTAIL.n78 B 0.023762f
C173 VTAIL.n79 B 0.010349f
C174 VTAIL.n80 B 0.010053f
C175 VTAIL.n81 B 0.018708f
C176 VTAIL.n82 B 0.018708f
C177 VTAIL.n83 B 0.010053f
C178 VTAIL.n84 B 0.010644f
C179 VTAIL.n85 B 0.023762f
C180 VTAIL.n86 B 0.053002f
C181 VTAIL.n87 B 0.010644f
C182 VTAIL.n88 B 0.010053f
C183 VTAIL.n89 B 0.048099f
C184 VTAIL.n90 B 0.02996f
C185 VTAIL.n91 B 0.18632f
C186 VTAIL.n92 B 0.02718f
C187 VTAIL.n93 B 0.018708f
C188 VTAIL.n94 B 0.010053f
C189 VTAIL.n95 B 0.023762f
C190 VTAIL.n96 B 0.010644f
C191 VTAIL.n97 B 0.018708f
C192 VTAIL.n98 B 0.010349f
C193 VTAIL.n99 B 0.023762f
C194 VTAIL.n100 B 0.010644f
C195 VTAIL.n101 B 0.018708f
C196 VTAIL.n102 B 0.010053f
C197 VTAIL.n103 B 0.023762f
C198 VTAIL.n104 B 0.010644f
C199 VTAIL.n105 B 0.018708f
C200 VTAIL.n106 B 0.010053f
C201 VTAIL.n107 B 0.023762f
C202 VTAIL.n108 B 0.010644f
C203 VTAIL.n109 B 0.018708f
C204 VTAIL.n110 B 0.010053f
C205 VTAIL.n111 B 0.023762f
C206 VTAIL.n112 B 0.010644f
C207 VTAIL.n113 B 0.018708f
C208 VTAIL.n114 B 0.010053f
C209 VTAIL.n115 B 0.023762f
C210 VTAIL.n116 B 0.010644f
C211 VTAIL.n117 B 0.018708f
C212 VTAIL.n118 B 0.010053f
C213 VTAIL.n119 B 0.017821f
C214 VTAIL.n120 B 0.014037f
C215 VTAIL.t11 B 0.039262f
C216 VTAIL.n121 B 0.127976f
C217 VTAIL.n122 B 1.32607f
C218 VTAIL.n123 B 0.010053f
C219 VTAIL.n124 B 0.010644f
C220 VTAIL.n125 B 0.023762f
C221 VTAIL.n126 B 0.023762f
C222 VTAIL.n127 B 0.010644f
C223 VTAIL.n128 B 0.010053f
C224 VTAIL.n129 B 0.018708f
C225 VTAIL.n130 B 0.018708f
C226 VTAIL.n131 B 0.010053f
C227 VTAIL.n132 B 0.010644f
C228 VTAIL.n133 B 0.023762f
C229 VTAIL.n134 B 0.023762f
C230 VTAIL.n135 B 0.010644f
C231 VTAIL.n136 B 0.010053f
C232 VTAIL.n137 B 0.018708f
C233 VTAIL.n138 B 0.018708f
C234 VTAIL.n139 B 0.010053f
C235 VTAIL.n140 B 0.010644f
C236 VTAIL.n141 B 0.023762f
C237 VTAIL.n142 B 0.023762f
C238 VTAIL.n143 B 0.010644f
C239 VTAIL.n144 B 0.010053f
C240 VTAIL.n145 B 0.018708f
C241 VTAIL.n146 B 0.018708f
C242 VTAIL.n147 B 0.010053f
C243 VTAIL.n148 B 0.010644f
C244 VTAIL.n149 B 0.023762f
C245 VTAIL.n150 B 0.023762f
C246 VTAIL.n151 B 0.010644f
C247 VTAIL.n152 B 0.010053f
C248 VTAIL.n153 B 0.018708f
C249 VTAIL.n154 B 0.018708f
C250 VTAIL.n155 B 0.010053f
C251 VTAIL.n156 B 0.010644f
C252 VTAIL.n157 B 0.023762f
C253 VTAIL.n158 B 0.023762f
C254 VTAIL.n159 B 0.010644f
C255 VTAIL.n160 B 0.010053f
C256 VTAIL.n161 B 0.018708f
C257 VTAIL.n162 B 0.018708f
C258 VTAIL.n163 B 0.010053f
C259 VTAIL.n164 B 0.010053f
C260 VTAIL.n165 B 0.010644f
C261 VTAIL.n166 B 0.023762f
C262 VTAIL.n167 B 0.023762f
C263 VTAIL.n168 B 0.023762f
C264 VTAIL.n169 B 0.010349f
C265 VTAIL.n170 B 0.010053f
C266 VTAIL.n171 B 0.018708f
C267 VTAIL.n172 B 0.018708f
C268 VTAIL.n173 B 0.010053f
C269 VTAIL.n174 B 0.010644f
C270 VTAIL.n175 B 0.023762f
C271 VTAIL.n176 B 0.053002f
C272 VTAIL.n177 B 0.010644f
C273 VTAIL.n178 B 0.010053f
C274 VTAIL.n179 B 0.048099f
C275 VTAIL.n180 B 0.02996f
C276 VTAIL.n181 B 0.18632f
C277 VTAIL.t13 B 0.240532f
C278 VTAIL.t10 B 0.240532f
C279 VTAIL.n182 B 2.1335f
C280 VTAIL.n183 B 0.455924f
C281 VTAIL.n184 B 0.02718f
C282 VTAIL.n185 B 0.018708f
C283 VTAIL.n186 B 0.010053f
C284 VTAIL.n187 B 0.023762f
C285 VTAIL.n188 B 0.010644f
C286 VTAIL.n189 B 0.018708f
C287 VTAIL.n190 B 0.010349f
C288 VTAIL.n191 B 0.023762f
C289 VTAIL.n192 B 0.010644f
C290 VTAIL.n193 B 0.018708f
C291 VTAIL.n194 B 0.010053f
C292 VTAIL.n195 B 0.023762f
C293 VTAIL.n196 B 0.010644f
C294 VTAIL.n197 B 0.018708f
C295 VTAIL.n198 B 0.010053f
C296 VTAIL.n199 B 0.023762f
C297 VTAIL.n200 B 0.010644f
C298 VTAIL.n201 B 0.018708f
C299 VTAIL.n202 B 0.010053f
C300 VTAIL.n203 B 0.023762f
C301 VTAIL.n204 B 0.010644f
C302 VTAIL.n205 B 0.018708f
C303 VTAIL.n206 B 0.010053f
C304 VTAIL.n207 B 0.023762f
C305 VTAIL.n208 B 0.010644f
C306 VTAIL.n209 B 0.018708f
C307 VTAIL.n210 B 0.010053f
C308 VTAIL.n211 B 0.017821f
C309 VTAIL.n212 B 0.014037f
C310 VTAIL.t15 B 0.039262f
C311 VTAIL.n213 B 0.127976f
C312 VTAIL.n214 B 1.32607f
C313 VTAIL.n215 B 0.010053f
C314 VTAIL.n216 B 0.010644f
C315 VTAIL.n217 B 0.023762f
C316 VTAIL.n218 B 0.023762f
C317 VTAIL.n219 B 0.010644f
C318 VTAIL.n220 B 0.010053f
C319 VTAIL.n221 B 0.018708f
C320 VTAIL.n222 B 0.018708f
C321 VTAIL.n223 B 0.010053f
C322 VTAIL.n224 B 0.010644f
C323 VTAIL.n225 B 0.023762f
C324 VTAIL.n226 B 0.023762f
C325 VTAIL.n227 B 0.010644f
C326 VTAIL.n228 B 0.010053f
C327 VTAIL.n229 B 0.018708f
C328 VTAIL.n230 B 0.018708f
C329 VTAIL.n231 B 0.010053f
C330 VTAIL.n232 B 0.010644f
C331 VTAIL.n233 B 0.023762f
C332 VTAIL.n234 B 0.023762f
C333 VTAIL.n235 B 0.010644f
C334 VTAIL.n236 B 0.010053f
C335 VTAIL.n237 B 0.018708f
C336 VTAIL.n238 B 0.018708f
C337 VTAIL.n239 B 0.010053f
C338 VTAIL.n240 B 0.010644f
C339 VTAIL.n241 B 0.023762f
C340 VTAIL.n242 B 0.023762f
C341 VTAIL.n243 B 0.010644f
C342 VTAIL.n244 B 0.010053f
C343 VTAIL.n245 B 0.018708f
C344 VTAIL.n246 B 0.018708f
C345 VTAIL.n247 B 0.010053f
C346 VTAIL.n248 B 0.010644f
C347 VTAIL.n249 B 0.023762f
C348 VTAIL.n250 B 0.023762f
C349 VTAIL.n251 B 0.010644f
C350 VTAIL.n252 B 0.010053f
C351 VTAIL.n253 B 0.018708f
C352 VTAIL.n254 B 0.018708f
C353 VTAIL.n255 B 0.010053f
C354 VTAIL.n256 B 0.010053f
C355 VTAIL.n257 B 0.010644f
C356 VTAIL.n258 B 0.023762f
C357 VTAIL.n259 B 0.023762f
C358 VTAIL.n260 B 0.023762f
C359 VTAIL.n261 B 0.010349f
C360 VTAIL.n262 B 0.010053f
C361 VTAIL.n263 B 0.018708f
C362 VTAIL.n264 B 0.018708f
C363 VTAIL.n265 B 0.010053f
C364 VTAIL.n266 B 0.010644f
C365 VTAIL.n267 B 0.023762f
C366 VTAIL.n268 B 0.053002f
C367 VTAIL.n269 B 0.010644f
C368 VTAIL.n270 B 0.010053f
C369 VTAIL.n271 B 0.048099f
C370 VTAIL.n272 B 0.02996f
C371 VTAIL.n273 B 1.39691f
C372 VTAIL.n274 B 0.02718f
C373 VTAIL.n275 B 0.018708f
C374 VTAIL.n276 B 0.010053f
C375 VTAIL.n277 B 0.023762f
C376 VTAIL.n278 B 0.010644f
C377 VTAIL.n279 B 0.018708f
C378 VTAIL.n280 B 0.010349f
C379 VTAIL.n281 B 0.023762f
C380 VTAIL.n282 B 0.010053f
C381 VTAIL.n283 B 0.010644f
C382 VTAIL.n284 B 0.018708f
C383 VTAIL.n285 B 0.010053f
C384 VTAIL.n286 B 0.023762f
C385 VTAIL.n287 B 0.010644f
C386 VTAIL.n288 B 0.018708f
C387 VTAIL.n289 B 0.010053f
C388 VTAIL.n290 B 0.023762f
C389 VTAIL.n291 B 0.010644f
C390 VTAIL.n292 B 0.018708f
C391 VTAIL.n293 B 0.010053f
C392 VTAIL.n294 B 0.023762f
C393 VTAIL.n295 B 0.010644f
C394 VTAIL.n296 B 0.018708f
C395 VTAIL.n297 B 0.010053f
C396 VTAIL.n298 B 0.023762f
C397 VTAIL.n299 B 0.010644f
C398 VTAIL.n300 B 0.018708f
C399 VTAIL.n301 B 0.010053f
C400 VTAIL.n302 B 0.017821f
C401 VTAIL.n303 B 0.014037f
C402 VTAIL.t6 B 0.039262f
C403 VTAIL.n304 B 0.127976f
C404 VTAIL.n305 B 1.32607f
C405 VTAIL.n306 B 0.010053f
C406 VTAIL.n307 B 0.010644f
C407 VTAIL.n308 B 0.023762f
C408 VTAIL.n309 B 0.023762f
C409 VTAIL.n310 B 0.010644f
C410 VTAIL.n311 B 0.010053f
C411 VTAIL.n312 B 0.018708f
C412 VTAIL.n313 B 0.018708f
C413 VTAIL.n314 B 0.010053f
C414 VTAIL.n315 B 0.010644f
C415 VTAIL.n316 B 0.023762f
C416 VTAIL.n317 B 0.023762f
C417 VTAIL.n318 B 0.010644f
C418 VTAIL.n319 B 0.010053f
C419 VTAIL.n320 B 0.018708f
C420 VTAIL.n321 B 0.018708f
C421 VTAIL.n322 B 0.010053f
C422 VTAIL.n323 B 0.010644f
C423 VTAIL.n324 B 0.023762f
C424 VTAIL.n325 B 0.023762f
C425 VTAIL.n326 B 0.010644f
C426 VTAIL.n327 B 0.010053f
C427 VTAIL.n328 B 0.018708f
C428 VTAIL.n329 B 0.018708f
C429 VTAIL.n330 B 0.010053f
C430 VTAIL.n331 B 0.010644f
C431 VTAIL.n332 B 0.023762f
C432 VTAIL.n333 B 0.023762f
C433 VTAIL.n334 B 0.010644f
C434 VTAIL.n335 B 0.010053f
C435 VTAIL.n336 B 0.018708f
C436 VTAIL.n337 B 0.018708f
C437 VTAIL.n338 B 0.010053f
C438 VTAIL.n339 B 0.010644f
C439 VTAIL.n340 B 0.023762f
C440 VTAIL.n341 B 0.023762f
C441 VTAIL.n342 B 0.010644f
C442 VTAIL.n343 B 0.010053f
C443 VTAIL.n344 B 0.018708f
C444 VTAIL.n345 B 0.018708f
C445 VTAIL.n346 B 0.010053f
C446 VTAIL.n347 B 0.010644f
C447 VTAIL.n348 B 0.023762f
C448 VTAIL.n349 B 0.023762f
C449 VTAIL.n350 B 0.023762f
C450 VTAIL.n351 B 0.010349f
C451 VTAIL.n352 B 0.010053f
C452 VTAIL.n353 B 0.018708f
C453 VTAIL.n354 B 0.018708f
C454 VTAIL.n355 B 0.010053f
C455 VTAIL.n356 B 0.010644f
C456 VTAIL.n357 B 0.023762f
C457 VTAIL.n358 B 0.053002f
C458 VTAIL.n359 B 0.010644f
C459 VTAIL.n360 B 0.010053f
C460 VTAIL.n361 B 0.048099f
C461 VTAIL.n362 B 0.02996f
C462 VTAIL.n363 B 1.39691f
C463 VTAIL.t5 B 0.240532f
C464 VTAIL.t7 B 0.240532f
C465 VTAIL.n364 B 2.1335f
C466 VTAIL.n365 B 0.455915f
C467 VTAIL.n366 B 0.02718f
C468 VTAIL.n367 B 0.018708f
C469 VTAIL.n368 B 0.010053f
C470 VTAIL.n369 B 0.023762f
C471 VTAIL.n370 B 0.010644f
C472 VTAIL.n371 B 0.018708f
C473 VTAIL.n372 B 0.010349f
C474 VTAIL.n373 B 0.023762f
C475 VTAIL.n374 B 0.010053f
C476 VTAIL.n375 B 0.010644f
C477 VTAIL.n376 B 0.018708f
C478 VTAIL.n377 B 0.010053f
C479 VTAIL.n378 B 0.023762f
C480 VTAIL.n379 B 0.010644f
C481 VTAIL.n380 B 0.018708f
C482 VTAIL.n381 B 0.010053f
C483 VTAIL.n382 B 0.023762f
C484 VTAIL.n383 B 0.010644f
C485 VTAIL.n384 B 0.018708f
C486 VTAIL.n385 B 0.010053f
C487 VTAIL.n386 B 0.023762f
C488 VTAIL.n387 B 0.010644f
C489 VTAIL.n388 B 0.018708f
C490 VTAIL.n389 B 0.010053f
C491 VTAIL.n390 B 0.023762f
C492 VTAIL.n391 B 0.010644f
C493 VTAIL.n392 B 0.018708f
C494 VTAIL.n393 B 0.010053f
C495 VTAIL.n394 B 0.017821f
C496 VTAIL.n395 B 0.014037f
C497 VTAIL.t0 B 0.039262f
C498 VTAIL.n396 B 0.127976f
C499 VTAIL.n397 B 1.32607f
C500 VTAIL.n398 B 0.010053f
C501 VTAIL.n399 B 0.010644f
C502 VTAIL.n400 B 0.023762f
C503 VTAIL.n401 B 0.023762f
C504 VTAIL.n402 B 0.010644f
C505 VTAIL.n403 B 0.010053f
C506 VTAIL.n404 B 0.018708f
C507 VTAIL.n405 B 0.018708f
C508 VTAIL.n406 B 0.010053f
C509 VTAIL.n407 B 0.010644f
C510 VTAIL.n408 B 0.023762f
C511 VTAIL.n409 B 0.023762f
C512 VTAIL.n410 B 0.010644f
C513 VTAIL.n411 B 0.010053f
C514 VTAIL.n412 B 0.018708f
C515 VTAIL.n413 B 0.018708f
C516 VTAIL.n414 B 0.010053f
C517 VTAIL.n415 B 0.010644f
C518 VTAIL.n416 B 0.023762f
C519 VTAIL.n417 B 0.023762f
C520 VTAIL.n418 B 0.010644f
C521 VTAIL.n419 B 0.010053f
C522 VTAIL.n420 B 0.018708f
C523 VTAIL.n421 B 0.018708f
C524 VTAIL.n422 B 0.010053f
C525 VTAIL.n423 B 0.010644f
C526 VTAIL.n424 B 0.023762f
C527 VTAIL.n425 B 0.023762f
C528 VTAIL.n426 B 0.010644f
C529 VTAIL.n427 B 0.010053f
C530 VTAIL.n428 B 0.018708f
C531 VTAIL.n429 B 0.018708f
C532 VTAIL.n430 B 0.010053f
C533 VTAIL.n431 B 0.010644f
C534 VTAIL.n432 B 0.023762f
C535 VTAIL.n433 B 0.023762f
C536 VTAIL.n434 B 0.010644f
C537 VTAIL.n435 B 0.010053f
C538 VTAIL.n436 B 0.018708f
C539 VTAIL.n437 B 0.018708f
C540 VTAIL.n438 B 0.010053f
C541 VTAIL.n439 B 0.010644f
C542 VTAIL.n440 B 0.023762f
C543 VTAIL.n441 B 0.023762f
C544 VTAIL.n442 B 0.023762f
C545 VTAIL.n443 B 0.010349f
C546 VTAIL.n444 B 0.010053f
C547 VTAIL.n445 B 0.018708f
C548 VTAIL.n446 B 0.018708f
C549 VTAIL.n447 B 0.010053f
C550 VTAIL.n448 B 0.010644f
C551 VTAIL.n449 B 0.023762f
C552 VTAIL.n450 B 0.053002f
C553 VTAIL.n451 B 0.010644f
C554 VTAIL.n452 B 0.010053f
C555 VTAIL.n453 B 0.048099f
C556 VTAIL.n454 B 0.02996f
C557 VTAIL.n455 B 0.18632f
C558 VTAIL.n456 B 0.02718f
C559 VTAIL.n457 B 0.018708f
C560 VTAIL.n458 B 0.010053f
C561 VTAIL.n459 B 0.023762f
C562 VTAIL.n460 B 0.010644f
C563 VTAIL.n461 B 0.018708f
C564 VTAIL.n462 B 0.010349f
C565 VTAIL.n463 B 0.023762f
C566 VTAIL.n464 B 0.010053f
C567 VTAIL.n465 B 0.010644f
C568 VTAIL.n466 B 0.018708f
C569 VTAIL.n467 B 0.010053f
C570 VTAIL.n468 B 0.023762f
C571 VTAIL.n469 B 0.010644f
C572 VTAIL.n470 B 0.018708f
C573 VTAIL.n471 B 0.010053f
C574 VTAIL.n472 B 0.023762f
C575 VTAIL.n473 B 0.010644f
C576 VTAIL.n474 B 0.018708f
C577 VTAIL.n475 B 0.010053f
C578 VTAIL.n476 B 0.023762f
C579 VTAIL.n477 B 0.010644f
C580 VTAIL.n478 B 0.018708f
C581 VTAIL.n479 B 0.010053f
C582 VTAIL.n480 B 0.023762f
C583 VTAIL.n481 B 0.010644f
C584 VTAIL.n482 B 0.018708f
C585 VTAIL.n483 B 0.010053f
C586 VTAIL.n484 B 0.017821f
C587 VTAIL.n485 B 0.014037f
C588 VTAIL.t8 B 0.039262f
C589 VTAIL.n486 B 0.127976f
C590 VTAIL.n487 B 1.32607f
C591 VTAIL.n488 B 0.010053f
C592 VTAIL.n489 B 0.010644f
C593 VTAIL.n490 B 0.023762f
C594 VTAIL.n491 B 0.023762f
C595 VTAIL.n492 B 0.010644f
C596 VTAIL.n493 B 0.010053f
C597 VTAIL.n494 B 0.018708f
C598 VTAIL.n495 B 0.018708f
C599 VTAIL.n496 B 0.010053f
C600 VTAIL.n497 B 0.010644f
C601 VTAIL.n498 B 0.023762f
C602 VTAIL.n499 B 0.023762f
C603 VTAIL.n500 B 0.010644f
C604 VTAIL.n501 B 0.010053f
C605 VTAIL.n502 B 0.018708f
C606 VTAIL.n503 B 0.018708f
C607 VTAIL.n504 B 0.010053f
C608 VTAIL.n505 B 0.010644f
C609 VTAIL.n506 B 0.023762f
C610 VTAIL.n507 B 0.023762f
C611 VTAIL.n508 B 0.010644f
C612 VTAIL.n509 B 0.010053f
C613 VTAIL.n510 B 0.018708f
C614 VTAIL.n511 B 0.018708f
C615 VTAIL.n512 B 0.010053f
C616 VTAIL.n513 B 0.010644f
C617 VTAIL.n514 B 0.023762f
C618 VTAIL.n515 B 0.023762f
C619 VTAIL.n516 B 0.010644f
C620 VTAIL.n517 B 0.010053f
C621 VTAIL.n518 B 0.018708f
C622 VTAIL.n519 B 0.018708f
C623 VTAIL.n520 B 0.010053f
C624 VTAIL.n521 B 0.010644f
C625 VTAIL.n522 B 0.023762f
C626 VTAIL.n523 B 0.023762f
C627 VTAIL.n524 B 0.010644f
C628 VTAIL.n525 B 0.010053f
C629 VTAIL.n526 B 0.018708f
C630 VTAIL.n527 B 0.018708f
C631 VTAIL.n528 B 0.010053f
C632 VTAIL.n529 B 0.010644f
C633 VTAIL.n530 B 0.023762f
C634 VTAIL.n531 B 0.023762f
C635 VTAIL.n532 B 0.023762f
C636 VTAIL.n533 B 0.010349f
C637 VTAIL.n534 B 0.010053f
C638 VTAIL.n535 B 0.018708f
C639 VTAIL.n536 B 0.018708f
C640 VTAIL.n537 B 0.010053f
C641 VTAIL.n538 B 0.010644f
C642 VTAIL.n539 B 0.023762f
C643 VTAIL.n540 B 0.053002f
C644 VTAIL.n541 B 0.010644f
C645 VTAIL.n542 B 0.010053f
C646 VTAIL.n543 B 0.048099f
C647 VTAIL.n544 B 0.02996f
C648 VTAIL.n545 B 0.18632f
C649 VTAIL.t9 B 0.240532f
C650 VTAIL.t12 B 0.240532f
C651 VTAIL.n546 B 2.1335f
C652 VTAIL.n547 B 0.455915f
C653 VTAIL.n548 B 0.02718f
C654 VTAIL.n549 B 0.018708f
C655 VTAIL.n550 B 0.010053f
C656 VTAIL.n551 B 0.023762f
C657 VTAIL.n552 B 0.010644f
C658 VTAIL.n553 B 0.018708f
C659 VTAIL.n554 B 0.010349f
C660 VTAIL.n555 B 0.023762f
C661 VTAIL.n556 B 0.010053f
C662 VTAIL.n557 B 0.010644f
C663 VTAIL.n558 B 0.018708f
C664 VTAIL.n559 B 0.010053f
C665 VTAIL.n560 B 0.023762f
C666 VTAIL.n561 B 0.010644f
C667 VTAIL.n562 B 0.018708f
C668 VTAIL.n563 B 0.010053f
C669 VTAIL.n564 B 0.023762f
C670 VTAIL.n565 B 0.010644f
C671 VTAIL.n566 B 0.018708f
C672 VTAIL.n567 B 0.010053f
C673 VTAIL.n568 B 0.023762f
C674 VTAIL.n569 B 0.010644f
C675 VTAIL.n570 B 0.018708f
C676 VTAIL.n571 B 0.010053f
C677 VTAIL.n572 B 0.023762f
C678 VTAIL.n573 B 0.010644f
C679 VTAIL.n574 B 0.018708f
C680 VTAIL.n575 B 0.010053f
C681 VTAIL.n576 B 0.017821f
C682 VTAIL.n577 B 0.014037f
C683 VTAIL.t14 B 0.039262f
C684 VTAIL.n578 B 0.127976f
C685 VTAIL.n579 B 1.32607f
C686 VTAIL.n580 B 0.010053f
C687 VTAIL.n581 B 0.010644f
C688 VTAIL.n582 B 0.023762f
C689 VTAIL.n583 B 0.023762f
C690 VTAIL.n584 B 0.010644f
C691 VTAIL.n585 B 0.010053f
C692 VTAIL.n586 B 0.018708f
C693 VTAIL.n587 B 0.018708f
C694 VTAIL.n588 B 0.010053f
C695 VTAIL.n589 B 0.010644f
C696 VTAIL.n590 B 0.023762f
C697 VTAIL.n591 B 0.023762f
C698 VTAIL.n592 B 0.010644f
C699 VTAIL.n593 B 0.010053f
C700 VTAIL.n594 B 0.018708f
C701 VTAIL.n595 B 0.018708f
C702 VTAIL.n596 B 0.010053f
C703 VTAIL.n597 B 0.010644f
C704 VTAIL.n598 B 0.023762f
C705 VTAIL.n599 B 0.023762f
C706 VTAIL.n600 B 0.010644f
C707 VTAIL.n601 B 0.010053f
C708 VTAIL.n602 B 0.018708f
C709 VTAIL.n603 B 0.018708f
C710 VTAIL.n604 B 0.010053f
C711 VTAIL.n605 B 0.010644f
C712 VTAIL.n606 B 0.023762f
C713 VTAIL.n607 B 0.023762f
C714 VTAIL.n608 B 0.010644f
C715 VTAIL.n609 B 0.010053f
C716 VTAIL.n610 B 0.018708f
C717 VTAIL.n611 B 0.018708f
C718 VTAIL.n612 B 0.010053f
C719 VTAIL.n613 B 0.010644f
C720 VTAIL.n614 B 0.023762f
C721 VTAIL.n615 B 0.023762f
C722 VTAIL.n616 B 0.010644f
C723 VTAIL.n617 B 0.010053f
C724 VTAIL.n618 B 0.018708f
C725 VTAIL.n619 B 0.018708f
C726 VTAIL.n620 B 0.010053f
C727 VTAIL.n621 B 0.010644f
C728 VTAIL.n622 B 0.023762f
C729 VTAIL.n623 B 0.023762f
C730 VTAIL.n624 B 0.023762f
C731 VTAIL.n625 B 0.010349f
C732 VTAIL.n626 B 0.010053f
C733 VTAIL.n627 B 0.018708f
C734 VTAIL.n628 B 0.018708f
C735 VTAIL.n629 B 0.010053f
C736 VTAIL.n630 B 0.010644f
C737 VTAIL.n631 B 0.023762f
C738 VTAIL.n632 B 0.053002f
C739 VTAIL.n633 B 0.010644f
C740 VTAIL.n634 B 0.010053f
C741 VTAIL.n635 B 0.048099f
C742 VTAIL.n636 B 0.02996f
C743 VTAIL.n637 B 1.39691f
C744 VTAIL.n638 B 0.02718f
C745 VTAIL.n639 B 0.018708f
C746 VTAIL.n640 B 0.010053f
C747 VTAIL.n641 B 0.023762f
C748 VTAIL.n642 B 0.010644f
C749 VTAIL.n643 B 0.018708f
C750 VTAIL.n644 B 0.010349f
C751 VTAIL.n645 B 0.023762f
C752 VTAIL.n646 B 0.010644f
C753 VTAIL.n647 B 0.018708f
C754 VTAIL.n648 B 0.010053f
C755 VTAIL.n649 B 0.023762f
C756 VTAIL.n650 B 0.010644f
C757 VTAIL.n651 B 0.018708f
C758 VTAIL.n652 B 0.010053f
C759 VTAIL.n653 B 0.023762f
C760 VTAIL.n654 B 0.010644f
C761 VTAIL.n655 B 0.018708f
C762 VTAIL.n656 B 0.010053f
C763 VTAIL.n657 B 0.023762f
C764 VTAIL.n658 B 0.010644f
C765 VTAIL.n659 B 0.018708f
C766 VTAIL.n660 B 0.010053f
C767 VTAIL.n661 B 0.023762f
C768 VTAIL.n662 B 0.010644f
C769 VTAIL.n663 B 0.018708f
C770 VTAIL.n664 B 0.010053f
C771 VTAIL.n665 B 0.017821f
C772 VTAIL.n666 B 0.014037f
C773 VTAIL.t3 B 0.039262f
C774 VTAIL.n667 B 0.127976f
C775 VTAIL.n668 B 1.32607f
C776 VTAIL.n669 B 0.010053f
C777 VTAIL.n670 B 0.010644f
C778 VTAIL.n671 B 0.023762f
C779 VTAIL.n672 B 0.023762f
C780 VTAIL.n673 B 0.010644f
C781 VTAIL.n674 B 0.010053f
C782 VTAIL.n675 B 0.018708f
C783 VTAIL.n676 B 0.018708f
C784 VTAIL.n677 B 0.010053f
C785 VTAIL.n678 B 0.010644f
C786 VTAIL.n679 B 0.023762f
C787 VTAIL.n680 B 0.023762f
C788 VTAIL.n681 B 0.010644f
C789 VTAIL.n682 B 0.010053f
C790 VTAIL.n683 B 0.018708f
C791 VTAIL.n684 B 0.018708f
C792 VTAIL.n685 B 0.010053f
C793 VTAIL.n686 B 0.010644f
C794 VTAIL.n687 B 0.023762f
C795 VTAIL.n688 B 0.023762f
C796 VTAIL.n689 B 0.010644f
C797 VTAIL.n690 B 0.010053f
C798 VTAIL.n691 B 0.018708f
C799 VTAIL.n692 B 0.018708f
C800 VTAIL.n693 B 0.010053f
C801 VTAIL.n694 B 0.010644f
C802 VTAIL.n695 B 0.023762f
C803 VTAIL.n696 B 0.023762f
C804 VTAIL.n697 B 0.010644f
C805 VTAIL.n698 B 0.010053f
C806 VTAIL.n699 B 0.018708f
C807 VTAIL.n700 B 0.018708f
C808 VTAIL.n701 B 0.010053f
C809 VTAIL.n702 B 0.010644f
C810 VTAIL.n703 B 0.023762f
C811 VTAIL.n704 B 0.023762f
C812 VTAIL.n705 B 0.010644f
C813 VTAIL.n706 B 0.010053f
C814 VTAIL.n707 B 0.018708f
C815 VTAIL.n708 B 0.018708f
C816 VTAIL.n709 B 0.010053f
C817 VTAIL.n710 B 0.010053f
C818 VTAIL.n711 B 0.010644f
C819 VTAIL.n712 B 0.023762f
C820 VTAIL.n713 B 0.023762f
C821 VTAIL.n714 B 0.023762f
C822 VTAIL.n715 B 0.010349f
C823 VTAIL.n716 B 0.010053f
C824 VTAIL.n717 B 0.018708f
C825 VTAIL.n718 B 0.018708f
C826 VTAIL.n719 B 0.010053f
C827 VTAIL.n720 B 0.010644f
C828 VTAIL.n721 B 0.023762f
C829 VTAIL.n722 B 0.053002f
C830 VTAIL.n723 B 0.010644f
C831 VTAIL.n724 B 0.010053f
C832 VTAIL.n725 B 0.048099f
C833 VTAIL.n726 B 0.02996f
C834 VTAIL.n727 B 1.3934f
C835 VDD1.t6 B 0.316795f
C836 VDD1.t7 B 0.316795f
C837 VDD1.n0 B 2.88688f
C838 VDD1.t3 B 0.316795f
C839 VDD1.t5 B 0.316795f
C840 VDD1.n1 B 2.8859f
C841 VDD1.t0 B 0.316795f
C842 VDD1.t1 B 0.316795f
C843 VDD1.n2 B 2.8859f
C844 VDD1.n3 B 3.39722f
C845 VDD1.t4 B 0.316795f
C846 VDD1.t2 B 0.316795f
C847 VDD1.n4 B 2.87784f
C848 VDD1.n5 B 3.16861f
C849 VP.n0 B 0.030457f
C850 VP.t4 B 2.42463f
C851 VP.n1 B 0.020171f
C852 VP.n2 B 0.023101f
C853 VP.t5 B 2.42463f
C854 VP.n3 B 0.043055f
C855 VP.n4 B 0.023101f
C856 VP.n5 B 0.025625f
C857 VP.n6 B 0.023101f
C858 VP.n7 B 0.046663f
C859 VP.n8 B 0.030457f
C860 VP.t1 B 2.42463f
C861 VP.n9 B 0.020171f
C862 VP.n10 B 0.023101f
C863 VP.t3 B 2.42463f
C864 VP.n11 B 0.043055f
C865 VP.n12 B 0.023101f
C866 VP.n13 B 0.025625f
C867 VP.t7 B 2.58148f
C868 VP.t6 B 2.42463f
C869 VP.n14 B 0.902719f
C870 VP.n15 B 0.897657f
C871 VP.n16 B 0.200111f
C872 VP.n17 B 0.023101f
C873 VP.n18 B 0.043055f
C874 VP.n19 B 0.033724f
C875 VP.n20 B 0.033724f
C876 VP.n21 B 0.023101f
C877 VP.n22 B 0.023101f
C878 VP.n23 B 0.023101f
C879 VP.n24 B 0.025625f
C880 VP.n25 B 0.846372f
C881 VP.n26 B 0.039229f
C882 VP.n27 B 0.043669f
C883 VP.n28 B 0.023101f
C884 VP.n29 B 0.023101f
C885 VP.n30 B 0.023101f
C886 VP.n31 B 0.046663f
C887 VP.n32 B 0.033277f
C888 VP.n33 B 0.920112f
C889 VP.n34 B 1.39363f
C890 VP.n35 B 1.40931f
C891 VP.t0 B 2.42463f
C892 VP.n36 B 0.920112f
C893 VP.n37 B 0.033277f
C894 VP.n38 B 0.030457f
C895 VP.n39 B 0.023101f
C896 VP.n40 B 0.023101f
C897 VP.n41 B 0.020171f
C898 VP.n42 B 0.043669f
C899 VP.t2 B 2.42463f
C900 VP.n43 B 0.846372f
C901 VP.n44 B 0.039229f
C902 VP.n45 B 0.023101f
C903 VP.n46 B 0.023101f
C904 VP.n47 B 0.023101f
C905 VP.n48 B 0.043055f
C906 VP.n49 B 0.033724f
C907 VP.n50 B 0.033724f
C908 VP.n51 B 0.023101f
C909 VP.n52 B 0.023101f
C910 VP.n53 B 0.023101f
C911 VP.n54 B 0.025625f
C912 VP.n55 B 0.846372f
C913 VP.n56 B 0.039229f
C914 VP.n57 B 0.043669f
C915 VP.n58 B 0.023101f
C916 VP.n59 B 0.023101f
C917 VP.n60 B 0.023101f
C918 VP.n61 B 0.046663f
C919 VP.n62 B 0.033277f
C920 VP.n63 B 0.920112f
C921 VP.n64 B 0.033975f
.ends

