* NGSPICE file created from diff_pair_sample_0422.ext - technology: sky130A

.subckt diff_pair_sample_0422 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t7 w_n5170_n3504# sky130_fd_pr__pfet_01v8 ad=2.0922 pd=13.01 as=2.0922 ps=13.01 w=12.68 l=3.87
X1 VTAIL.t14 VN.t1 VDD2.t6 w_n5170_n3504# sky130_fd_pr__pfet_01v8 ad=2.0922 pd=13.01 as=2.0922 ps=13.01 w=12.68 l=3.87
X2 VTAIL.t5 VP.t0 VDD1.t7 w_n5170_n3504# sky130_fd_pr__pfet_01v8 ad=2.0922 pd=13.01 as=2.0922 ps=13.01 w=12.68 l=3.87
X3 VTAIL.t13 VN.t2 VDD2.t5 w_n5170_n3504# sky130_fd_pr__pfet_01v8 ad=4.9452 pd=26.14 as=2.0922 ps=13.01 w=12.68 l=3.87
X4 VDD1.t6 VP.t1 VTAIL.t1 w_n5170_n3504# sky130_fd_pr__pfet_01v8 ad=2.0922 pd=13.01 as=2.0922 ps=13.01 w=12.68 l=3.87
X5 B.t11 B.t9 B.t10 w_n5170_n3504# sky130_fd_pr__pfet_01v8 ad=4.9452 pd=26.14 as=0 ps=0 w=12.68 l=3.87
X6 VTAIL.t0 VP.t2 VDD1.t5 w_n5170_n3504# sky130_fd_pr__pfet_01v8 ad=4.9452 pd=26.14 as=2.0922 ps=13.01 w=12.68 l=3.87
X7 VDD2.t1 VN.t3 VTAIL.t12 w_n5170_n3504# sky130_fd_pr__pfet_01v8 ad=2.0922 pd=13.01 as=4.9452 ps=26.14 w=12.68 l=3.87
X8 VTAIL.t3 VP.t3 VDD1.t4 w_n5170_n3504# sky130_fd_pr__pfet_01v8 ad=4.9452 pd=26.14 as=2.0922 ps=13.01 w=12.68 l=3.87
X9 VDD1.t3 VP.t4 VTAIL.t4 w_n5170_n3504# sky130_fd_pr__pfet_01v8 ad=2.0922 pd=13.01 as=4.9452 ps=26.14 w=12.68 l=3.87
X10 VDD2.t0 VN.t4 VTAIL.t11 w_n5170_n3504# sky130_fd_pr__pfet_01v8 ad=2.0922 pd=13.01 as=4.9452 ps=26.14 w=12.68 l=3.87
X11 VTAIL.t10 VN.t5 VDD2.t3 w_n5170_n3504# sky130_fd_pr__pfet_01v8 ad=4.9452 pd=26.14 as=2.0922 ps=13.01 w=12.68 l=3.87
X12 B.t8 B.t6 B.t7 w_n5170_n3504# sky130_fd_pr__pfet_01v8 ad=4.9452 pd=26.14 as=0 ps=0 w=12.68 l=3.87
X13 B.t5 B.t3 B.t4 w_n5170_n3504# sky130_fd_pr__pfet_01v8 ad=4.9452 pd=26.14 as=0 ps=0 w=12.68 l=3.87
X14 VDD1.t2 VP.t5 VTAIL.t7 w_n5170_n3504# sky130_fd_pr__pfet_01v8 ad=2.0922 pd=13.01 as=4.9452 ps=26.14 w=12.68 l=3.87
X15 VTAIL.t6 VP.t6 VDD1.t1 w_n5170_n3504# sky130_fd_pr__pfet_01v8 ad=2.0922 pd=13.01 as=2.0922 ps=13.01 w=12.68 l=3.87
X16 VDD1.t0 VP.t7 VTAIL.t2 w_n5170_n3504# sky130_fd_pr__pfet_01v8 ad=2.0922 pd=13.01 as=2.0922 ps=13.01 w=12.68 l=3.87
X17 VDD2.t2 VN.t6 VTAIL.t9 w_n5170_n3504# sky130_fd_pr__pfet_01v8 ad=2.0922 pd=13.01 as=2.0922 ps=13.01 w=12.68 l=3.87
X18 B.t2 B.t0 B.t1 w_n5170_n3504# sky130_fd_pr__pfet_01v8 ad=4.9452 pd=26.14 as=0 ps=0 w=12.68 l=3.87
X19 VDD2.t4 VN.t7 VTAIL.t8 w_n5170_n3504# sky130_fd_pr__pfet_01v8 ad=2.0922 pd=13.01 as=2.0922 ps=13.01 w=12.68 l=3.87
R0 VN.n76 VN.n75 161.3
R1 VN.n74 VN.n40 161.3
R2 VN.n73 VN.n72 161.3
R3 VN.n71 VN.n41 161.3
R4 VN.n70 VN.n69 161.3
R5 VN.n68 VN.n42 161.3
R6 VN.n67 VN.n66 161.3
R7 VN.n65 VN.n43 161.3
R8 VN.n64 VN.n63 161.3
R9 VN.n61 VN.n44 161.3
R10 VN.n60 VN.n59 161.3
R11 VN.n58 VN.n45 161.3
R12 VN.n57 VN.n56 161.3
R13 VN.n55 VN.n46 161.3
R14 VN.n54 VN.n53 161.3
R15 VN.n52 VN.n47 161.3
R16 VN.n51 VN.n50 161.3
R17 VN.n37 VN.n36 161.3
R18 VN.n35 VN.n1 161.3
R19 VN.n34 VN.n33 161.3
R20 VN.n32 VN.n2 161.3
R21 VN.n31 VN.n30 161.3
R22 VN.n29 VN.n3 161.3
R23 VN.n28 VN.n27 161.3
R24 VN.n26 VN.n4 161.3
R25 VN.n25 VN.n24 161.3
R26 VN.n22 VN.n5 161.3
R27 VN.n21 VN.n20 161.3
R28 VN.n19 VN.n6 161.3
R29 VN.n18 VN.n17 161.3
R30 VN.n16 VN.n7 161.3
R31 VN.n15 VN.n14 161.3
R32 VN.n13 VN.n8 161.3
R33 VN.n12 VN.n11 161.3
R34 VN.n48 VN.t3 111.776
R35 VN.n9 VN.t5 111.776
R36 VN.n38 VN.n0 87.7864
R37 VN.n77 VN.n39 87.7864
R38 VN.n10 VN.t6 78.9638
R39 VN.n23 VN.t1 78.9638
R40 VN.n0 VN.t4 78.9638
R41 VN.n49 VN.t0 78.9638
R42 VN.n62 VN.t7 78.9638
R43 VN.n39 VN.t2 78.9638
R44 VN.n10 VN.n9 58.1068
R45 VN.n49 VN.n48 58.1068
R46 VN VN.n77 57.5815
R47 VN.n17 VN.n16 56.5617
R48 VN.n56 VN.n55 56.5617
R49 VN.n30 VN.n29 45.4209
R50 VN.n69 VN.n68 45.4209
R51 VN.n30 VN.n2 35.7332
R52 VN.n69 VN.n41 35.7332
R53 VN.n11 VN.n8 24.5923
R54 VN.n15 VN.n8 24.5923
R55 VN.n16 VN.n15 24.5923
R56 VN.n17 VN.n6 24.5923
R57 VN.n21 VN.n6 24.5923
R58 VN.n22 VN.n21 24.5923
R59 VN.n24 VN.n4 24.5923
R60 VN.n28 VN.n4 24.5923
R61 VN.n29 VN.n28 24.5923
R62 VN.n34 VN.n2 24.5923
R63 VN.n35 VN.n34 24.5923
R64 VN.n36 VN.n35 24.5923
R65 VN.n55 VN.n54 24.5923
R66 VN.n54 VN.n47 24.5923
R67 VN.n50 VN.n47 24.5923
R68 VN.n68 VN.n67 24.5923
R69 VN.n67 VN.n43 24.5923
R70 VN.n63 VN.n43 24.5923
R71 VN.n61 VN.n60 24.5923
R72 VN.n60 VN.n45 24.5923
R73 VN.n56 VN.n45 24.5923
R74 VN.n75 VN.n74 24.5923
R75 VN.n74 VN.n73 24.5923
R76 VN.n73 VN.n41 24.5923
R77 VN.n11 VN.n10 17.2148
R78 VN.n23 VN.n22 17.2148
R79 VN.n50 VN.n49 17.2148
R80 VN.n62 VN.n61 17.2148
R81 VN.n24 VN.n23 7.37805
R82 VN.n63 VN.n62 7.37805
R83 VN.n12 VN.n9 2.46316
R84 VN.n51 VN.n48 2.46316
R85 VN.n36 VN.n0 2.45968
R86 VN.n75 VN.n39 2.45968
R87 VN.n77 VN.n76 0.354861
R88 VN.n38 VN.n37 0.354861
R89 VN VN.n38 0.267071
R90 VN.n76 VN.n40 0.189894
R91 VN.n72 VN.n40 0.189894
R92 VN.n72 VN.n71 0.189894
R93 VN.n71 VN.n70 0.189894
R94 VN.n70 VN.n42 0.189894
R95 VN.n66 VN.n42 0.189894
R96 VN.n66 VN.n65 0.189894
R97 VN.n65 VN.n64 0.189894
R98 VN.n64 VN.n44 0.189894
R99 VN.n59 VN.n44 0.189894
R100 VN.n59 VN.n58 0.189894
R101 VN.n58 VN.n57 0.189894
R102 VN.n57 VN.n46 0.189894
R103 VN.n53 VN.n46 0.189894
R104 VN.n53 VN.n52 0.189894
R105 VN.n52 VN.n51 0.189894
R106 VN.n13 VN.n12 0.189894
R107 VN.n14 VN.n13 0.189894
R108 VN.n14 VN.n7 0.189894
R109 VN.n18 VN.n7 0.189894
R110 VN.n19 VN.n18 0.189894
R111 VN.n20 VN.n19 0.189894
R112 VN.n20 VN.n5 0.189894
R113 VN.n25 VN.n5 0.189894
R114 VN.n26 VN.n25 0.189894
R115 VN.n27 VN.n26 0.189894
R116 VN.n27 VN.n3 0.189894
R117 VN.n31 VN.n3 0.189894
R118 VN.n32 VN.n31 0.189894
R119 VN.n33 VN.n32 0.189894
R120 VN.n33 VN.n1 0.189894
R121 VN.n37 VN.n1 0.189894
R122 VDD2.n2 VDD2.n1 78.2886
R123 VDD2.n2 VDD2.n0 78.2886
R124 VDD2 VDD2.n5 78.2856
R125 VDD2.n4 VDD2.n3 76.5346
R126 VDD2.n4 VDD2.n2 50.9394
R127 VDD2.n5 VDD2.t7 2.56399
R128 VDD2.n5 VDD2.t1 2.56399
R129 VDD2.n3 VDD2.t5 2.56399
R130 VDD2.n3 VDD2.t4 2.56399
R131 VDD2.n1 VDD2.t6 2.56399
R132 VDD2.n1 VDD2.t0 2.56399
R133 VDD2.n0 VDD2.t3 2.56399
R134 VDD2.n0 VDD2.t2 2.56399
R135 VDD2 VDD2.n4 1.86903
R136 VTAIL.n566 VTAIL.n565 756.745
R137 VTAIL.n70 VTAIL.n69 756.745
R138 VTAIL.n140 VTAIL.n139 756.745
R139 VTAIL.n212 VTAIL.n211 756.745
R140 VTAIL.n496 VTAIL.n495 756.745
R141 VTAIL.n424 VTAIL.n423 756.745
R142 VTAIL.n354 VTAIL.n353 756.745
R143 VTAIL.n282 VTAIL.n281 756.745
R144 VTAIL.n520 VTAIL.n519 585
R145 VTAIL.n525 VTAIL.n524 585
R146 VTAIL.n527 VTAIL.n526 585
R147 VTAIL.n516 VTAIL.n515 585
R148 VTAIL.n533 VTAIL.n532 585
R149 VTAIL.n535 VTAIL.n534 585
R150 VTAIL.n512 VTAIL.n511 585
R151 VTAIL.n541 VTAIL.n540 585
R152 VTAIL.n543 VTAIL.n542 585
R153 VTAIL.n508 VTAIL.n507 585
R154 VTAIL.n549 VTAIL.n548 585
R155 VTAIL.n551 VTAIL.n550 585
R156 VTAIL.n504 VTAIL.n503 585
R157 VTAIL.n557 VTAIL.n556 585
R158 VTAIL.n559 VTAIL.n558 585
R159 VTAIL.n500 VTAIL.n499 585
R160 VTAIL.n565 VTAIL.n564 585
R161 VTAIL.n24 VTAIL.n23 585
R162 VTAIL.n29 VTAIL.n28 585
R163 VTAIL.n31 VTAIL.n30 585
R164 VTAIL.n20 VTAIL.n19 585
R165 VTAIL.n37 VTAIL.n36 585
R166 VTAIL.n39 VTAIL.n38 585
R167 VTAIL.n16 VTAIL.n15 585
R168 VTAIL.n45 VTAIL.n44 585
R169 VTAIL.n47 VTAIL.n46 585
R170 VTAIL.n12 VTAIL.n11 585
R171 VTAIL.n53 VTAIL.n52 585
R172 VTAIL.n55 VTAIL.n54 585
R173 VTAIL.n8 VTAIL.n7 585
R174 VTAIL.n61 VTAIL.n60 585
R175 VTAIL.n63 VTAIL.n62 585
R176 VTAIL.n4 VTAIL.n3 585
R177 VTAIL.n69 VTAIL.n68 585
R178 VTAIL.n94 VTAIL.n93 585
R179 VTAIL.n99 VTAIL.n98 585
R180 VTAIL.n101 VTAIL.n100 585
R181 VTAIL.n90 VTAIL.n89 585
R182 VTAIL.n107 VTAIL.n106 585
R183 VTAIL.n109 VTAIL.n108 585
R184 VTAIL.n86 VTAIL.n85 585
R185 VTAIL.n115 VTAIL.n114 585
R186 VTAIL.n117 VTAIL.n116 585
R187 VTAIL.n82 VTAIL.n81 585
R188 VTAIL.n123 VTAIL.n122 585
R189 VTAIL.n125 VTAIL.n124 585
R190 VTAIL.n78 VTAIL.n77 585
R191 VTAIL.n131 VTAIL.n130 585
R192 VTAIL.n133 VTAIL.n132 585
R193 VTAIL.n74 VTAIL.n73 585
R194 VTAIL.n139 VTAIL.n138 585
R195 VTAIL.n166 VTAIL.n165 585
R196 VTAIL.n171 VTAIL.n170 585
R197 VTAIL.n173 VTAIL.n172 585
R198 VTAIL.n162 VTAIL.n161 585
R199 VTAIL.n179 VTAIL.n178 585
R200 VTAIL.n181 VTAIL.n180 585
R201 VTAIL.n158 VTAIL.n157 585
R202 VTAIL.n187 VTAIL.n186 585
R203 VTAIL.n189 VTAIL.n188 585
R204 VTAIL.n154 VTAIL.n153 585
R205 VTAIL.n195 VTAIL.n194 585
R206 VTAIL.n197 VTAIL.n196 585
R207 VTAIL.n150 VTAIL.n149 585
R208 VTAIL.n203 VTAIL.n202 585
R209 VTAIL.n205 VTAIL.n204 585
R210 VTAIL.n146 VTAIL.n145 585
R211 VTAIL.n211 VTAIL.n210 585
R212 VTAIL.n495 VTAIL.n494 585
R213 VTAIL.n430 VTAIL.n429 585
R214 VTAIL.n489 VTAIL.n488 585
R215 VTAIL.n487 VTAIL.n486 585
R216 VTAIL.n434 VTAIL.n433 585
R217 VTAIL.n481 VTAIL.n480 585
R218 VTAIL.n479 VTAIL.n478 585
R219 VTAIL.n438 VTAIL.n437 585
R220 VTAIL.n473 VTAIL.n472 585
R221 VTAIL.n471 VTAIL.n470 585
R222 VTAIL.n442 VTAIL.n441 585
R223 VTAIL.n465 VTAIL.n464 585
R224 VTAIL.n463 VTAIL.n462 585
R225 VTAIL.n446 VTAIL.n445 585
R226 VTAIL.n457 VTAIL.n456 585
R227 VTAIL.n455 VTAIL.n454 585
R228 VTAIL.n450 VTAIL.n449 585
R229 VTAIL.n423 VTAIL.n422 585
R230 VTAIL.n358 VTAIL.n357 585
R231 VTAIL.n417 VTAIL.n416 585
R232 VTAIL.n415 VTAIL.n414 585
R233 VTAIL.n362 VTAIL.n361 585
R234 VTAIL.n409 VTAIL.n408 585
R235 VTAIL.n407 VTAIL.n406 585
R236 VTAIL.n366 VTAIL.n365 585
R237 VTAIL.n401 VTAIL.n400 585
R238 VTAIL.n399 VTAIL.n398 585
R239 VTAIL.n370 VTAIL.n369 585
R240 VTAIL.n393 VTAIL.n392 585
R241 VTAIL.n391 VTAIL.n390 585
R242 VTAIL.n374 VTAIL.n373 585
R243 VTAIL.n385 VTAIL.n384 585
R244 VTAIL.n383 VTAIL.n382 585
R245 VTAIL.n378 VTAIL.n377 585
R246 VTAIL.n353 VTAIL.n352 585
R247 VTAIL.n288 VTAIL.n287 585
R248 VTAIL.n347 VTAIL.n346 585
R249 VTAIL.n345 VTAIL.n344 585
R250 VTAIL.n292 VTAIL.n291 585
R251 VTAIL.n339 VTAIL.n338 585
R252 VTAIL.n337 VTAIL.n336 585
R253 VTAIL.n296 VTAIL.n295 585
R254 VTAIL.n331 VTAIL.n330 585
R255 VTAIL.n329 VTAIL.n328 585
R256 VTAIL.n300 VTAIL.n299 585
R257 VTAIL.n323 VTAIL.n322 585
R258 VTAIL.n321 VTAIL.n320 585
R259 VTAIL.n304 VTAIL.n303 585
R260 VTAIL.n315 VTAIL.n314 585
R261 VTAIL.n313 VTAIL.n312 585
R262 VTAIL.n308 VTAIL.n307 585
R263 VTAIL.n281 VTAIL.n280 585
R264 VTAIL.n216 VTAIL.n215 585
R265 VTAIL.n275 VTAIL.n274 585
R266 VTAIL.n273 VTAIL.n272 585
R267 VTAIL.n220 VTAIL.n219 585
R268 VTAIL.n267 VTAIL.n266 585
R269 VTAIL.n265 VTAIL.n264 585
R270 VTAIL.n224 VTAIL.n223 585
R271 VTAIL.n259 VTAIL.n258 585
R272 VTAIL.n257 VTAIL.n256 585
R273 VTAIL.n228 VTAIL.n227 585
R274 VTAIL.n251 VTAIL.n250 585
R275 VTAIL.n249 VTAIL.n248 585
R276 VTAIL.n232 VTAIL.n231 585
R277 VTAIL.n243 VTAIL.n242 585
R278 VTAIL.n241 VTAIL.n240 585
R279 VTAIL.n236 VTAIL.n235 585
R280 VTAIL.n521 VTAIL.t11 327.466
R281 VTAIL.n25 VTAIL.t10 327.466
R282 VTAIL.n95 VTAIL.t4 327.466
R283 VTAIL.n167 VTAIL.t3 327.466
R284 VTAIL.n451 VTAIL.t7 327.466
R285 VTAIL.n379 VTAIL.t0 327.466
R286 VTAIL.n309 VTAIL.t12 327.466
R287 VTAIL.n237 VTAIL.t13 327.466
R288 VTAIL.n525 VTAIL.n519 171.744
R289 VTAIL.n526 VTAIL.n525 171.744
R290 VTAIL.n526 VTAIL.n515 171.744
R291 VTAIL.n533 VTAIL.n515 171.744
R292 VTAIL.n534 VTAIL.n533 171.744
R293 VTAIL.n534 VTAIL.n511 171.744
R294 VTAIL.n541 VTAIL.n511 171.744
R295 VTAIL.n542 VTAIL.n541 171.744
R296 VTAIL.n542 VTAIL.n507 171.744
R297 VTAIL.n549 VTAIL.n507 171.744
R298 VTAIL.n550 VTAIL.n549 171.744
R299 VTAIL.n550 VTAIL.n503 171.744
R300 VTAIL.n557 VTAIL.n503 171.744
R301 VTAIL.n558 VTAIL.n557 171.744
R302 VTAIL.n558 VTAIL.n499 171.744
R303 VTAIL.n565 VTAIL.n499 171.744
R304 VTAIL.n29 VTAIL.n23 171.744
R305 VTAIL.n30 VTAIL.n29 171.744
R306 VTAIL.n30 VTAIL.n19 171.744
R307 VTAIL.n37 VTAIL.n19 171.744
R308 VTAIL.n38 VTAIL.n37 171.744
R309 VTAIL.n38 VTAIL.n15 171.744
R310 VTAIL.n45 VTAIL.n15 171.744
R311 VTAIL.n46 VTAIL.n45 171.744
R312 VTAIL.n46 VTAIL.n11 171.744
R313 VTAIL.n53 VTAIL.n11 171.744
R314 VTAIL.n54 VTAIL.n53 171.744
R315 VTAIL.n54 VTAIL.n7 171.744
R316 VTAIL.n61 VTAIL.n7 171.744
R317 VTAIL.n62 VTAIL.n61 171.744
R318 VTAIL.n62 VTAIL.n3 171.744
R319 VTAIL.n69 VTAIL.n3 171.744
R320 VTAIL.n99 VTAIL.n93 171.744
R321 VTAIL.n100 VTAIL.n99 171.744
R322 VTAIL.n100 VTAIL.n89 171.744
R323 VTAIL.n107 VTAIL.n89 171.744
R324 VTAIL.n108 VTAIL.n107 171.744
R325 VTAIL.n108 VTAIL.n85 171.744
R326 VTAIL.n115 VTAIL.n85 171.744
R327 VTAIL.n116 VTAIL.n115 171.744
R328 VTAIL.n116 VTAIL.n81 171.744
R329 VTAIL.n123 VTAIL.n81 171.744
R330 VTAIL.n124 VTAIL.n123 171.744
R331 VTAIL.n124 VTAIL.n77 171.744
R332 VTAIL.n131 VTAIL.n77 171.744
R333 VTAIL.n132 VTAIL.n131 171.744
R334 VTAIL.n132 VTAIL.n73 171.744
R335 VTAIL.n139 VTAIL.n73 171.744
R336 VTAIL.n171 VTAIL.n165 171.744
R337 VTAIL.n172 VTAIL.n171 171.744
R338 VTAIL.n172 VTAIL.n161 171.744
R339 VTAIL.n179 VTAIL.n161 171.744
R340 VTAIL.n180 VTAIL.n179 171.744
R341 VTAIL.n180 VTAIL.n157 171.744
R342 VTAIL.n187 VTAIL.n157 171.744
R343 VTAIL.n188 VTAIL.n187 171.744
R344 VTAIL.n188 VTAIL.n153 171.744
R345 VTAIL.n195 VTAIL.n153 171.744
R346 VTAIL.n196 VTAIL.n195 171.744
R347 VTAIL.n196 VTAIL.n149 171.744
R348 VTAIL.n203 VTAIL.n149 171.744
R349 VTAIL.n204 VTAIL.n203 171.744
R350 VTAIL.n204 VTAIL.n145 171.744
R351 VTAIL.n211 VTAIL.n145 171.744
R352 VTAIL.n495 VTAIL.n429 171.744
R353 VTAIL.n488 VTAIL.n429 171.744
R354 VTAIL.n488 VTAIL.n487 171.744
R355 VTAIL.n487 VTAIL.n433 171.744
R356 VTAIL.n480 VTAIL.n433 171.744
R357 VTAIL.n480 VTAIL.n479 171.744
R358 VTAIL.n479 VTAIL.n437 171.744
R359 VTAIL.n472 VTAIL.n437 171.744
R360 VTAIL.n472 VTAIL.n471 171.744
R361 VTAIL.n471 VTAIL.n441 171.744
R362 VTAIL.n464 VTAIL.n441 171.744
R363 VTAIL.n464 VTAIL.n463 171.744
R364 VTAIL.n463 VTAIL.n445 171.744
R365 VTAIL.n456 VTAIL.n445 171.744
R366 VTAIL.n456 VTAIL.n455 171.744
R367 VTAIL.n455 VTAIL.n449 171.744
R368 VTAIL.n423 VTAIL.n357 171.744
R369 VTAIL.n416 VTAIL.n357 171.744
R370 VTAIL.n416 VTAIL.n415 171.744
R371 VTAIL.n415 VTAIL.n361 171.744
R372 VTAIL.n408 VTAIL.n361 171.744
R373 VTAIL.n408 VTAIL.n407 171.744
R374 VTAIL.n407 VTAIL.n365 171.744
R375 VTAIL.n400 VTAIL.n365 171.744
R376 VTAIL.n400 VTAIL.n399 171.744
R377 VTAIL.n399 VTAIL.n369 171.744
R378 VTAIL.n392 VTAIL.n369 171.744
R379 VTAIL.n392 VTAIL.n391 171.744
R380 VTAIL.n391 VTAIL.n373 171.744
R381 VTAIL.n384 VTAIL.n373 171.744
R382 VTAIL.n384 VTAIL.n383 171.744
R383 VTAIL.n383 VTAIL.n377 171.744
R384 VTAIL.n353 VTAIL.n287 171.744
R385 VTAIL.n346 VTAIL.n287 171.744
R386 VTAIL.n346 VTAIL.n345 171.744
R387 VTAIL.n345 VTAIL.n291 171.744
R388 VTAIL.n338 VTAIL.n291 171.744
R389 VTAIL.n338 VTAIL.n337 171.744
R390 VTAIL.n337 VTAIL.n295 171.744
R391 VTAIL.n330 VTAIL.n295 171.744
R392 VTAIL.n330 VTAIL.n329 171.744
R393 VTAIL.n329 VTAIL.n299 171.744
R394 VTAIL.n322 VTAIL.n299 171.744
R395 VTAIL.n322 VTAIL.n321 171.744
R396 VTAIL.n321 VTAIL.n303 171.744
R397 VTAIL.n314 VTAIL.n303 171.744
R398 VTAIL.n314 VTAIL.n313 171.744
R399 VTAIL.n313 VTAIL.n307 171.744
R400 VTAIL.n281 VTAIL.n215 171.744
R401 VTAIL.n274 VTAIL.n215 171.744
R402 VTAIL.n274 VTAIL.n273 171.744
R403 VTAIL.n273 VTAIL.n219 171.744
R404 VTAIL.n266 VTAIL.n219 171.744
R405 VTAIL.n266 VTAIL.n265 171.744
R406 VTAIL.n265 VTAIL.n223 171.744
R407 VTAIL.n258 VTAIL.n223 171.744
R408 VTAIL.n258 VTAIL.n257 171.744
R409 VTAIL.n257 VTAIL.n227 171.744
R410 VTAIL.n250 VTAIL.n227 171.744
R411 VTAIL.n250 VTAIL.n249 171.744
R412 VTAIL.n249 VTAIL.n231 171.744
R413 VTAIL.n242 VTAIL.n231 171.744
R414 VTAIL.n242 VTAIL.n241 171.744
R415 VTAIL.n241 VTAIL.n235 171.744
R416 VTAIL.t11 VTAIL.n519 85.8723
R417 VTAIL.t10 VTAIL.n23 85.8723
R418 VTAIL.t4 VTAIL.n93 85.8723
R419 VTAIL.t3 VTAIL.n165 85.8723
R420 VTAIL.t7 VTAIL.n449 85.8723
R421 VTAIL.t0 VTAIL.n377 85.8723
R422 VTAIL.t12 VTAIL.n307 85.8723
R423 VTAIL.t13 VTAIL.n235 85.8723
R424 VTAIL.n427 VTAIL.n426 59.8558
R425 VTAIL.n285 VTAIL.n284 59.8558
R426 VTAIL.n1 VTAIL.n0 59.8548
R427 VTAIL.n143 VTAIL.n142 59.8548
R428 VTAIL.n567 VTAIL.n566 35.6763
R429 VTAIL.n71 VTAIL.n70 35.6763
R430 VTAIL.n141 VTAIL.n140 35.6763
R431 VTAIL.n213 VTAIL.n212 35.6763
R432 VTAIL.n497 VTAIL.n496 35.6763
R433 VTAIL.n425 VTAIL.n424 35.6763
R434 VTAIL.n355 VTAIL.n354 35.6763
R435 VTAIL.n283 VTAIL.n282 35.6763
R436 VTAIL.n567 VTAIL.n497 26.9186
R437 VTAIL.n283 VTAIL.n213 26.9186
R438 VTAIL.n521 VTAIL.n520 16.3895
R439 VTAIL.n25 VTAIL.n24 16.3895
R440 VTAIL.n95 VTAIL.n94 16.3895
R441 VTAIL.n167 VTAIL.n166 16.3895
R442 VTAIL.n451 VTAIL.n450 16.3895
R443 VTAIL.n379 VTAIL.n378 16.3895
R444 VTAIL.n309 VTAIL.n308 16.3895
R445 VTAIL.n237 VTAIL.n236 16.3895
R446 VTAIL.n524 VTAIL.n523 12.8005
R447 VTAIL.n564 VTAIL.n498 12.8005
R448 VTAIL.n28 VTAIL.n27 12.8005
R449 VTAIL.n68 VTAIL.n2 12.8005
R450 VTAIL.n98 VTAIL.n97 12.8005
R451 VTAIL.n138 VTAIL.n72 12.8005
R452 VTAIL.n170 VTAIL.n169 12.8005
R453 VTAIL.n210 VTAIL.n144 12.8005
R454 VTAIL.n494 VTAIL.n428 12.8005
R455 VTAIL.n454 VTAIL.n453 12.8005
R456 VTAIL.n422 VTAIL.n356 12.8005
R457 VTAIL.n382 VTAIL.n381 12.8005
R458 VTAIL.n352 VTAIL.n286 12.8005
R459 VTAIL.n312 VTAIL.n311 12.8005
R460 VTAIL.n280 VTAIL.n214 12.8005
R461 VTAIL.n240 VTAIL.n239 12.8005
R462 VTAIL.n527 VTAIL.n518 12.0247
R463 VTAIL.n563 VTAIL.n500 12.0247
R464 VTAIL.n31 VTAIL.n22 12.0247
R465 VTAIL.n67 VTAIL.n4 12.0247
R466 VTAIL.n101 VTAIL.n92 12.0247
R467 VTAIL.n137 VTAIL.n74 12.0247
R468 VTAIL.n173 VTAIL.n164 12.0247
R469 VTAIL.n209 VTAIL.n146 12.0247
R470 VTAIL.n493 VTAIL.n430 12.0247
R471 VTAIL.n457 VTAIL.n448 12.0247
R472 VTAIL.n421 VTAIL.n358 12.0247
R473 VTAIL.n385 VTAIL.n376 12.0247
R474 VTAIL.n351 VTAIL.n288 12.0247
R475 VTAIL.n315 VTAIL.n306 12.0247
R476 VTAIL.n279 VTAIL.n216 12.0247
R477 VTAIL.n243 VTAIL.n234 12.0247
R478 VTAIL.n528 VTAIL.n516 11.249
R479 VTAIL.n560 VTAIL.n559 11.249
R480 VTAIL.n32 VTAIL.n20 11.249
R481 VTAIL.n64 VTAIL.n63 11.249
R482 VTAIL.n102 VTAIL.n90 11.249
R483 VTAIL.n134 VTAIL.n133 11.249
R484 VTAIL.n174 VTAIL.n162 11.249
R485 VTAIL.n206 VTAIL.n205 11.249
R486 VTAIL.n490 VTAIL.n489 11.249
R487 VTAIL.n458 VTAIL.n446 11.249
R488 VTAIL.n418 VTAIL.n417 11.249
R489 VTAIL.n386 VTAIL.n374 11.249
R490 VTAIL.n348 VTAIL.n347 11.249
R491 VTAIL.n316 VTAIL.n304 11.249
R492 VTAIL.n276 VTAIL.n275 11.249
R493 VTAIL.n244 VTAIL.n232 11.249
R494 VTAIL.n532 VTAIL.n531 10.4732
R495 VTAIL.n556 VTAIL.n502 10.4732
R496 VTAIL.n36 VTAIL.n35 10.4732
R497 VTAIL.n60 VTAIL.n6 10.4732
R498 VTAIL.n106 VTAIL.n105 10.4732
R499 VTAIL.n130 VTAIL.n76 10.4732
R500 VTAIL.n178 VTAIL.n177 10.4732
R501 VTAIL.n202 VTAIL.n148 10.4732
R502 VTAIL.n486 VTAIL.n432 10.4732
R503 VTAIL.n462 VTAIL.n461 10.4732
R504 VTAIL.n414 VTAIL.n360 10.4732
R505 VTAIL.n390 VTAIL.n389 10.4732
R506 VTAIL.n344 VTAIL.n290 10.4732
R507 VTAIL.n320 VTAIL.n319 10.4732
R508 VTAIL.n272 VTAIL.n218 10.4732
R509 VTAIL.n248 VTAIL.n247 10.4732
R510 VTAIL.n535 VTAIL.n514 9.69747
R511 VTAIL.n555 VTAIL.n504 9.69747
R512 VTAIL.n39 VTAIL.n18 9.69747
R513 VTAIL.n59 VTAIL.n8 9.69747
R514 VTAIL.n109 VTAIL.n88 9.69747
R515 VTAIL.n129 VTAIL.n78 9.69747
R516 VTAIL.n181 VTAIL.n160 9.69747
R517 VTAIL.n201 VTAIL.n150 9.69747
R518 VTAIL.n485 VTAIL.n434 9.69747
R519 VTAIL.n465 VTAIL.n444 9.69747
R520 VTAIL.n413 VTAIL.n362 9.69747
R521 VTAIL.n393 VTAIL.n372 9.69747
R522 VTAIL.n343 VTAIL.n292 9.69747
R523 VTAIL.n323 VTAIL.n302 9.69747
R524 VTAIL.n271 VTAIL.n220 9.69747
R525 VTAIL.n251 VTAIL.n230 9.69747
R526 VTAIL.n562 VTAIL.n498 9.45567
R527 VTAIL.n66 VTAIL.n2 9.45567
R528 VTAIL.n136 VTAIL.n72 9.45567
R529 VTAIL.n208 VTAIL.n144 9.45567
R530 VTAIL.n492 VTAIL.n428 9.45567
R531 VTAIL.n420 VTAIL.n356 9.45567
R532 VTAIL.n350 VTAIL.n286 9.45567
R533 VTAIL.n278 VTAIL.n214 9.45567
R534 VTAIL.n545 VTAIL.n544 9.3005
R535 VTAIL.n547 VTAIL.n546 9.3005
R536 VTAIL.n506 VTAIL.n505 9.3005
R537 VTAIL.n553 VTAIL.n552 9.3005
R538 VTAIL.n555 VTAIL.n554 9.3005
R539 VTAIL.n502 VTAIL.n501 9.3005
R540 VTAIL.n561 VTAIL.n560 9.3005
R541 VTAIL.n563 VTAIL.n562 9.3005
R542 VTAIL.n539 VTAIL.n538 9.3005
R543 VTAIL.n537 VTAIL.n536 9.3005
R544 VTAIL.n514 VTAIL.n513 9.3005
R545 VTAIL.n531 VTAIL.n530 9.3005
R546 VTAIL.n529 VTAIL.n528 9.3005
R547 VTAIL.n518 VTAIL.n517 9.3005
R548 VTAIL.n523 VTAIL.n522 9.3005
R549 VTAIL.n510 VTAIL.n509 9.3005
R550 VTAIL.n49 VTAIL.n48 9.3005
R551 VTAIL.n51 VTAIL.n50 9.3005
R552 VTAIL.n10 VTAIL.n9 9.3005
R553 VTAIL.n57 VTAIL.n56 9.3005
R554 VTAIL.n59 VTAIL.n58 9.3005
R555 VTAIL.n6 VTAIL.n5 9.3005
R556 VTAIL.n65 VTAIL.n64 9.3005
R557 VTAIL.n67 VTAIL.n66 9.3005
R558 VTAIL.n43 VTAIL.n42 9.3005
R559 VTAIL.n41 VTAIL.n40 9.3005
R560 VTAIL.n18 VTAIL.n17 9.3005
R561 VTAIL.n35 VTAIL.n34 9.3005
R562 VTAIL.n33 VTAIL.n32 9.3005
R563 VTAIL.n22 VTAIL.n21 9.3005
R564 VTAIL.n27 VTAIL.n26 9.3005
R565 VTAIL.n14 VTAIL.n13 9.3005
R566 VTAIL.n119 VTAIL.n118 9.3005
R567 VTAIL.n121 VTAIL.n120 9.3005
R568 VTAIL.n80 VTAIL.n79 9.3005
R569 VTAIL.n127 VTAIL.n126 9.3005
R570 VTAIL.n129 VTAIL.n128 9.3005
R571 VTAIL.n76 VTAIL.n75 9.3005
R572 VTAIL.n135 VTAIL.n134 9.3005
R573 VTAIL.n137 VTAIL.n136 9.3005
R574 VTAIL.n113 VTAIL.n112 9.3005
R575 VTAIL.n111 VTAIL.n110 9.3005
R576 VTAIL.n88 VTAIL.n87 9.3005
R577 VTAIL.n105 VTAIL.n104 9.3005
R578 VTAIL.n103 VTAIL.n102 9.3005
R579 VTAIL.n92 VTAIL.n91 9.3005
R580 VTAIL.n97 VTAIL.n96 9.3005
R581 VTAIL.n84 VTAIL.n83 9.3005
R582 VTAIL.n191 VTAIL.n190 9.3005
R583 VTAIL.n193 VTAIL.n192 9.3005
R584 VTAIL.n152 VTAIL.n151 9.3005
R585 VTAIL.n199 VTAIL.n198 9.3005
R586 VTAIL.n201 VTAIL.n200 9.3005
R587 VTAIL.n148 VTAIL.n147 9.3005
R588 VTAIL.n207 VTAIL.n206 9.3005
R589 VTAIL.n209 VTAIL.n208 9.3005
R590 VTAIL.n185 VTAIL.n184 9.3005
R591 VTAIL.n183 VTAIL.n182 9.3005
R592 VTAIL.n160 VTAIL.n159 9.3005
R593 VTAIL.n177 VTAIL.n176 9.3005
R594 VTAIL.n175 VTAIL.n174 9.3005
R595 VTAIL.n164 VTAIL.n163 9.3005
R596 VTAIL.n169 VTAIL.n168 9.3005
R597 VTAIL.n156 VTAIL.n155 9.3005
R598 VTAIL.n493 VTAIL.n492 9.3005
R599 VTAIL.n491 VTAIL.n490 9.3005
R600 VTAIL.n432 VTAIL.n431 9.3005
R601 VTAIL.n485 VTAIL.n484 9.3005
R602 VTAIL.n483 VTAIL.n482 9.3005
R603 VTAIL.n436 VTAIL.n435 9.3005
R604 VTAIL.n477 VTAIL.n476 9.3005
R605 VTAIL.n475 VTAIL.n474 9.3005
R606 VTAIL.n440 VTAIL.n439 9.3005
R607 VTAIL.n469 VTAIL.n468 9.3005
R608 VTAIL.n467 VTAIL.n466 9.3005
R609 VTAIL.n444 VTAIL.n443 9.3005
R610 VTAIL.n461 VTAIL.n460 9.3005
R611 VTAIL.n459 VTAIL.n458 9.3005
R612 VTAIL.n448 VTAIL.n447 9.3005
R613 VTAIL.n453 VTAIL.n452 9.3005
R614 VTAIL.n405 VTAIL.n404 9.3005
R615 VTAIL.n364 VTAIL.n363 9.3005
R616 VTAIL.n411 VTAIL.n410 9.3005
R617 VTAIL.n413 VTAIL.n412 9.3005
R618 VTAIL.n360 VTAIL.n359 9.3005
R619 VTAIL.n419 VTAIL.n418 9.3005
R620 VTAIL.n421 VTAIL.n420 9.3005
R621 VTAIL.n403 VTAIL.n402 9.3005
R622 VTAIL.n368 VTAIL.n367 9.3005
R623 VTAIL.n397 VTAIL.n396 9.3005
R624 VTAIL.n395 VTAIL.n394 9.3005
R625 VTAIL.n372 VTAIL.n371 9.3005
R626 VTAIL.n389 VTAIL.n388 9.3005
R627 VTAIL.n387 VTAIL.n386 9.3005
R628 VTAIL.n376 VTAIL.n375 9.3005
R629 VTAIL.n381 VTAIL.n380 9.3005
R630 VTAIL.n335 VTAIL.n334 9.3005
R631 VTAIL.n294 VTAIL.n293 9.3005
R632 VTAIL.n341 VTAIL.n340 9.3005
R633 VTAIL.n343 VTAIL.n342 9.3005
R634 VTAIL.n290 VTAIL.n289 9.3005
R635 VTAIL.n349 VTAIL.n348 9.3005
R636 VTAIL.n351 VTAIL.n350 9.3005
R637 VTAIL.n333 VTAIL.n332 9.3005
R638 VTAIL.n298 VTAIL.n297 9.3005
R639 VTAIL.n327 VTAIL.n326 9.3005
R640 VTAIL.n325 VTAIL.n324 9.3005
R641 VTAIL.n302 VTAIL.n301 9.3005
R642 VTAIL.n319 VTAIL.n318 9.3005
R643 VTAIL.n317 VTAIL.n316 9.3005
R644 VTAIL.n306 VTAIL.n305 9.3005
R645 VTAIL.n311 VTAIL.n310 9.3005
R646 VTAIL.n263 VTAIL.n262 9.3005
R647 VTAIL.n222 VTAIL.n221 9.3005
R648 VTAIL.n269 VTAIL.n268 9.3005
R649 VTAIL.n271 VTAIL.n270 9.3005
R650 VTAIL.n218 VTAIL.n217 9.3005
R651 VTAIL.n277 VTAIL.n276 9.3005
R652 VTAIL.n279 VTAIL.n278 9.3005
R653 VTAIL.n261 VTAIL.n260 9.3005
R654 VTAIL.n226 VTAIL.n225 9.3005
R655 VTAIL.n255 VTAIL.n254 9.3005
R656 VTAIL.n253 VTAIL.n252 9.3005
R657 VTAIL.n230 VTAIL.n229 9.3005
R658 VTAIL.n247 VTAIL.n246 9.3005
R659 VTAIL.n245 VTAIL.n244 9.3005
R660 VTAIL.n234 VTAIL.n233 9.3005
R661 VTAIL.n239 VTAIL.n238 9.3005
R662 VTAIL.n536 VTAIL.n512 8.92171
R663 VTAIL.n552 VTAIL.n551 8.92171
R664 VTAIL.n40 VTAIL.n16 8.92171
R665 VTAIL.n56 VTAIL.n55 8.92171
R666 VTAIL.n110 VTAIL.n86 8.92171
R667 VTAIL.n126 VTAIL.n125 8.92171
R668 VTAIL.n182 VTAIL.n158 8.92171
R669 VTAIL.n198 VTAIL.n197 8.92171
R670 VTAIL.n482 VTAIL.n481 8.92171
R671 VTAIL.n466 VTAIL.n442 8.92171
R672 VTAIL.n410 VTAIL.n409 8.92171
R673 VTAIL.n394 VTAIL.n370 8.92171
R674 VTAIL.n340 VTAIL.n339 8.92171
R675 VTAIL.n324 VTAIL.n300 8.92171
R676 VTAIL.n268 VTAIL.n267 8.92171
R677 VTAIL.n252 VTAIL.n228 8.92171
R678 VTAIL.n540 VTAIL.n539 8.14595
R679 VTAIL.n548 VTAIL.n506 8.14595
R680 VTAIL.n44 VTAIL.n43 8.14595
R681 VTAIL.n52 VTAIL.n10 8.14595
R682 VTAIL.n114 VTAIL.n113 8.14595
R683 VTAIL.n122 VTAIL.n80 8.14595
R684 VTAIL.n186 VTAIL.n185 8.14595
R685 VTAIL.n194 VTAIL.n152 8.14595
R686 VTAIL.n478 VTAIL.n436 8.14595
R687 VTAIL.n470 VTAIL.n469 8.14595
R688 VTAIL.n406 VTAIL.n364 8.14595
R689 VTAIL.n398 VTAIL.n397 8.14595
R690 VTAIL.n336 VTAIL.n294 8.14595
R691 VTAIL.n328 VTAIL.n327 8.14595
R692 VTAIL.n264 VTAIL.n222 8.14595
R693 VTAIL.n256 VTAIL.n255 8.14595
R694 VTAIL.n543 VTAIL.n510 7.3702
R695 VTAIL.n547 VTAIL.n508 7.3702
R696 VTAIL.n47 VTAIL.n14 7.3702
R697 VTAIL.n51 VTAIL.n12 7.3702
R698 VTAIL.n117 VTAIL.n84 7.3702
R699 VTAIL.n121 VTAIL.n82 7.3702
R700 VTAIL.n189 VTAIL.n156 7.3702
R701 VTAIL.n193 VTAIL.n154 7.3702
R702 VTAIL.n477 VTAIL.n438 7.3702
R703 VTAIL.n473 VTAIL.n440 7.3702
R704 VTAIL.n405 VTAIL.n366 7.3702
R705 VTAIL.n401 VTAIL.n368 7.3702
R706 VTAIL.n335 VTAIL.n296 7.3702
R707 VTAIL.n331 VTAIL.n298 7.3702
R708 VTAIL.n263 VTAIL.n224 7.3702
R709 VTAIL.n259 VTAIL.n226 7.3702
R710 VTAIL.n544 VTAIL.n543 6.59444
R711 VTAIL.n544 VTAIL.n508 6.59444
R712 VTAIL.n48 VTAIL.n47 6.59444
R713 VTAIL.n48 VTAIL.n12 6.59444
R714 VTAIL.n118 VTAIL.n117 6.59444
R715 VTAIL.n118 VTAIL.n82 6.59444
R716 VTAIL.n190 VTAIL.n189 6.59444
R717 VTAIL.n190 VTAIL.n154 6.59444
R718 VTAIL.n474 VTAIL.n438 6.59444
R719 VTAIL.n474 VTAIL.n473 6.59444
R720 VTAIL.n402 VTAIL.n366 6.59444
R721 VTAIL.n402 VTAIL.n401 6.59444
R722 VTAIL.n332 VTAIL.n296 6.59444
R723 VTAIL.n332 VTAIL.n331 6.59444
R724 VTAIL.n260 VTAIL.n224 6.59444
R725 VTAIL.n260 VTAIL.n259 6.59444
R726 VTAIL.n540 VTAIL.n510 5.81868
R727 VTAIL.n548 VTAIL.n547 5.81868
R728 VTAIL.n44 VTAIL.n14 5.81868
R729 VTAIL.n52 VTAIL.n51 5.81868
R730 VTAIL.n114 VTAIL.n84 5.81868
R731 VTAIL.n122 VTAIL.n121 5.81868
R732 VTAIL.n186 VTAIL.n156 5.81868
R733 VTAIL.n194 VTAIL.n193 5.81868
R734 VTAIL.n478 VTAIL.n477 5.81868
R735 VTAIL.n470 VTAIL.n440 5.81868
R736 VTAIL.n406 VTAIL.n405 5.81868
R737 VTAIL.n398 VTAIL.n368 5.81868
R738 VTAIL.n336 VTAIL.n335 5.81868
R739 VTAIL.n328 VTAIL.n298 5.81868
R740 VTAIL.n264 VTAIL.n263 5.81868
R741 VTAIL.n256 VTAIL.n226 5.81868
R742 VTAIL.n539 VTAIL.n512 5.04292
R743 VTAIL.n551 VTAIL.n506 5.04292
R744 VTAIL.n43 VTAIL.n16 5.04292
R745 VTAIL.n55 VTAIL.n10 5.04292
R746 VTAIL.n113 VTAIL.n86 5.04292
R747 VTAIL.n125 VTAIL.n80 5.04292
R748 VTAIL.n185 VTAIL.n158 5.04292
R749 VTAIL.n197 VTAIL.n152 5.04292
R750 VTAIL.n481 VTAIL.n436 5.04292
R751 VTAIL.n469 VTAIL.n442 5.04292
R752 VTAIL.n409 VTAIL.n364 5.04292
R753 VTAIL.n397 VTAIL.n370 5.04292
R754 VTAIL.n339 VTAIL.n294 5.04292
R755 VTAIL.n327 VTAIL.n300 5.04292
R756 VTAIL.n267 VTAIL.n222 5.04292
R757 VTAIL.n255 VTAIL.n228 5.04292
R758 VTAIL.n536 VTAIL.n535 4.26717
R759 VTAIL.n552 VTAIL.n504 4.26717
R760 VTAIL.n40 VTAIL.n39 4.26717
R761 VTAIL.n56 VTAIL.n8 4.26717
R762 VTAIL.n110 VTAIL.n109 4.26717
R763 VTAIL.n126 VTAIL.n78 4.26717
R764 VTAIL.n182 VTAIL.n181 4.26717
R765 VTAIL.n198 VTAIL.n150 4.26717
R766 VTAIL.n482 VTAIL.n434 4.26717
R767 VTAIL.n466 VTAIL.n465 4.26717
R768 VTAIL.n410 VTAIL.n362 4.26717
R769 VTAIL.n394 VTAIL.n393 4.26717
R770 VTAIL.n340 VTAIL.n292 4.26717
R771 VTAIL.n324 VTAIL.n323 4.26717
R772 VTAIL.n268 VTAIL.n220 4.26717
R773 VTAIL.n252 VTAIL.n251 4.26717
R774 VTAIL.n522 VTAIL.n521 3.70982
R775 VTAIL.n26 VTAIL.n25 3.70982
R776 VTAIL.n96 VTAIL.n95 3.70982
R777 VTAIL.n168 VTAIL.n167 3.70982
R778 VTAIL.n452 VTAIL.n451 3.70982
R779 VTAIL.n380 VTAIL.n379 3.70982
R780 VTAIL.n310 VTAIL.n309 3.70982
R781 VTAIL.n238 VTAIL.n237 3.70982
R782 VTAIL.n285 VTAIL.n283 3.62119
R783 VTAIL.n355 VTAIL.n285 3.62119
R784 VTAIL.n427 VTAIL.n425 3.62119
R785 VTAIL.n497 VTAIL.n427 3.62119
R786 VTAIL.n213 VTAIL.n143 3.62119
R787 VTAIL.n143 VTAIL.n141 3.62119
R788 VTAIL.n71 VTAIL.n1 3.62119
R789 VTAIL VTAIL.n567 3.563
R790 VTAIL.n532 VTAIL.n514 3.49141
R791 VTAIL.n556 VTAIL.n555 3.49141
R792 VTAIL.n36 VTAIL.n18 3.49141
R793 VTAIL.n60 VTAIL.n59 3.49141
R794 VTAIL.n106 VTAIL.n88 3.49141
R795 VTAIL.n130 VTAIL.n129 3.49141
R796 VTAIL.n178 VTAIL.n160 3.49141
R797 VTAIL.n202 VTAIL.n201 3.49141
R798 VTAIL.n486 VTAIL.n485 3.49141
R799 VTAIL.n462 VTAIL.n444 3.49141
R800 VTAIL.n414 VTAIL.n413 3.49141
R801 VTAIL.n390 VTAIL.n372 3.49141
R802 VTAIL.n344 VTAIL.n343 3.49141
R803 VTAIL.n320 VTAIL.n302 3.49141
R804 VTAIL.n272 VTAIL.n271 3.49141
R805 VTAIL.n248 VTAIL.n230 3.49141
R806 VTAIL.n531 VTAIL.n516 2.71565
R807 VTAIL.n559 VTAIL.n502 2.71565
R808 VTAIL.n35 VTAIL.n20 2.71565
R809 VTAIL.n63 VTAIL.n6 2.71565
R810 VTAIL.n105 VTAIL.n90 2.71565
R811 VTAIL.n133 VTAIL.n76 2.71565
R812 VTAIL.n177 VTAIL.n162 2.71565
R813 VTAIL.n205 VTAIL.n148 2.71565
R814 VTAIL.n489 VTAIL.n432 2.71565
R815 VTAIL.n461 VTAIL.n446 2.71565
R816 VTAIL.n417 VTAIL.n360 2.71565
R817 VTAIL.n389 VTAIL.n374 2.71565
R818 VTAIL.n347 VTAIL.n290 2.71565
R819 VTAIL.n319 VTAIL.n304 2.71565
R820 VTAIL.n275 VTAIL.n218 2.71565
R821 VTAIL.n247 VTAIL.n232 2.71565
R822 VTAIL.n0 VTAIL.t9 2.56399
R823 VTAIL.n0 VTAIL.t14 2.56399
R824 VTAIL.n142 VTAIL.t1 2.56399
R825 VTAIL.n142 VTAIL.t6 2.56399
R826 VTAIL.n426 VTAIL.t2 2.56399
R827 VTAIL.n426 VTAIL.t5 2.56399
R828 VTAIL.n284 VTAIL.t8 2.56399
R829 VTAIL.n284 VTAIL.t15 2.56399
R830 VTAIL.n528 VTAIL.n527 1.93989
R831 VTAIL.n560 VTAIL.n500 1.93989
R832 VTAIL.n32 VTAIL.n31 1.93989
R833 VTAIL.n64 VTAIL.n4 1.93989
R834 VTAIL.n102 VTAIL.n101 1.93989
R835 VTAIL.n134 VTAIL.n74 1.93989
R836 VTAIL.n174 VTAIL.n173 1.93989
R837 VTAIL.n206 VTAIL.n146 1.93989
R838 VTAIL.n490 VTAIL.n430 1.93989
R839 VTAIL.n458 VTAIL.n457 1.93989
R840 VTAIL.n418 VTAIL.n358 1.93989
R841 VTAIL.n386 VTAIL.n385 1.93989
R842 VTAIL.n348 VTAIL.n288 1.93989
R843 VTAIL.n316 VTAIL.n315 1.93989
R844 VTAIL.n276 VTAIL.n216 1.93989
R845 VTAIL.n244 VTAIL.n243 1.93989
R846 VTAIL.n524 VTAIL.n518 1.16414
R847 VTAIL.n564 VTAIL.n563 1.16414
R848 VTAIL.n28 VTAIL.n22 1.16414
R849 VTAIL.n68 VTAIL.n67 1.16414
R850 VTAIL.n98 VTAIL.n92 1.16414
R851 VTAIL.n138 VTAIL.n137 1.16414
R852 VTAIL.n170 VTAIL.n164 1.16414
R853 VTAIL.n210 VTAIL.n209 1.16414
R854 VTAIL.n494 VTAIL.n493 1.16414
R855 VTAIL.n454 VTAIL.n448 1.16414
R856 VTAIL.n422 VTAIL.n421 1.16414
R857 VTAIL.n382 VTAIL.n376 1.16414
R858 VTAIL.n352 VTAIL.n351 1.16414
R859 VTAIL.n312 VTAIL.n306 1.16414
R860 VTAIL.n280 VTAIL.n279 1.16414
R861 VTAIL.n240 VTAIL.n234 1.16414
R862 VTAIL.n425 VTAIL.n355 0.470328
R863 VTAIL.n141 VTAIL.n71 0.470328
R864 VTAIL.n523 VTAIL.n520 0.388379
R865 VTAIL.n566 VTAIL.n498 0.388379
R866 VTAIL.n27 VTAIL.n24 0.388379
R867 VTAIL.n70 VTAIL.n2 0.388379
R868 VTAIL.n97 VTAIL.n94 0.388379
R869 VTAIL.n140 VTAIL.n72 0.388379
R870 VTAIL.n169 VTAIL.n166 0.388379
R871 VTAIL.n212 VTAIL.n144 0.388379
R872 VTAIL.n496 VTAIL.n428 0.388379
R873 VTAIL.n453 VTAIL.n450 0.388379
R874 VTAIL.n424 VTAIL.n356 0.388379
R875 VTAIL.n381 VTAIL.n378 0.388379
R876 VTAIL.n354 VTAIL.n286 0.388379
R877 VTAIL.n311 VTAIL.n308 0.388379
R878 VTAIL.n282 VTAIL.n214 0.388379
R879 VTAIL.n239 VTAIL.n236 0.388379
R880 VTAIL.n522 VTAIL.n517 0.155672
R881 VTAIL.n529 VTAIL.n517 0.155672
R882 VTAIL.n530 VTAIL.n529 0.155672
R883 VTAIL.n530 VTAIL.n513 0.155672
R884 VTAIL.n537 VTAIL.n513 0.155672
R885 VTAIL.n538 VTAIL.n537 0.155672
R886 VTAIL.n538 VTAIL.n509 0.155672
R887 VTAIL.n545 VTAIL.n509 0.155672
R888 VTAIL.n546 VTAIL.n545 0.155672
R889 VTAIL.n546 VTAIL.n505 0.155672
R890 VTAIL.n553 VTAIL.n505 0.155672
R891 VTAIL.n554 VTAIL.n553 0.155672
R892 VTAIL.n554 VTAIL.n501 0.155672
R893 VTAIL.n561 VTAIL.n501 0.155672
R894 VTAIL.n562 VTAIL.n561 0.155672
R895 VTAIL.n26 VTAIL.n21 0.155672
R896 VTAIL.n33 VTAIL.n21 0.155672
R897 VTAIL.n34 VTAIL.n33 0.155672
R898 VTAIL.n34 VTAIL.n17 0.155672
R899 VTAIL.n41 VTAIL.n17 0.155672
R900 VTAIL.n42 VTAIL.n41 0.155672
R901 VTAIL.n42 VTAIL.n13 0.155672
R902 VTAIL.n49 VTAIL.n13 0.155672
R903 VTAIL.n50 VTAIL.n49 0.155672
R904 VTAIL.n50 VTAIL.n9 0.155672
R905 VTAIL.n57 VTAIL.n9 0.155672
R906 VTAIL.n58 VTAIL.n57 0.155672
R907 VTAIL.n58 VTAIL.n5 0.155672
R908 VTAIL.n65 VTAIL.n5 0.155672
R909 VTAIL.n66 VTAIL.n65 0.155672
R910 VTAIL.n96 VTAIL.n91 0.155672
R911 VTAIL.n103 VTAIL.n91 0.155672
R912 VTAIL.n104 VTAIL.n103 0.155672
R913 VTAIL.n104 VTAIL.n87 0.155672
R914 VTAIL.n111 VTAIL.n87 0.155672
R915 VTAIL.n112 VTAIL.n111 0.155672
R916 VTAIL.n112 VTAIL.n83 0.155672
R917 VTAIL.n119 VTAIL.n83 0.155672
R918 VTAIL.n120 VTAIL.n119 0.155672
R919 VTAIL.n120 VTAIL.n79 0.155672
R920 VTAIL.n127 VTAIL.n79 0.155672
R921 VTAIL.n128 VTAIL.n127 0.155672
R922 VTAIL.n128 VTAIL.n75 0.155672
R923 VTAIL.n135 VTAIL.n75 0.155672
R924 VTAIL.n136 VTAIL.n135 0.155672
R925 VTAIL.n168 VTAIL.n163 0.155672
R926 VTAIL.n175 VTAIL.n163 0.155672
R927 VTAIL.n176 VTAIL.n175 0.155672
R928 VTAIL.n176 VTAIL.n159 0.155672
R929 VTAIL.n183 VTAIL.n159 0.155672
R930 VTAIL.n184 VTAIL.n183 0.155672
R931 VTAIL.n184 VTAIL.n155 0.155672
R932 VTAIL.n191 VTAIL.n155 0.155672
R933 VTAIL.n192 VTAIL.n191 0.155672
R934 VTAIL.n192 VTAIL.n151 0.155672
R935 VTAIL.n199 VTAIL.n151 0.155672
R936 VTAIL.n200 VTAIL.n199 0.155672
R937 VTAIL.n200 VTAIL.n147 0.155672
R938 VTAIL.n207 VTAIL.n147 0.155672
R939 VTAIL.n208 VTAIL.n207 0.155672
R940 VTAIL.n492 VTAIL.n491 0.155672
R941 VTAIL.n491 VTAIL.n431 0.155672
R942 VTAIL.n484 VTAIL.n431 0.155672
R943 VTAIL.n484 VTAIL.n483 0.155672
R944 VTAIL.n483 VTAIL.n435 0.155672
R945 VTAIL.n476 VTAIL.n435 0.155672
R946 VTAIL.n476 VTAIL.n475 0.155672
R947 VTAIL.n475 VTAIL.n439 0.155672
R948 VTAIL.n468 VTAIL.n439 0.155672
R949 VTAIL.n468 VTAIL.n467 0.155672
R950 VTAIL.n467 VTAIL.n443 0.155672
R951 VTAIL.n460 VTAIL.n443 0.155672
R952 VTAIL.n460 VTAIL.n459 0.155672
R953 VTAIL.n459 VTAIL.n447 0.155672
R954 VTAIL.n452 VTAIL.n447 0.155672
R955 VTAIL.n420 VTAIL.n419 0.155672
R956 VTAIL.n419 VTAIL.n359 0.155672
R957 VTAIL.n412 VTAIL.n359 0.155672
R958 VTAIL.n412 VTAIL.n411 0.155672
R959 VTAIL.n411 VTAIL.n363 0.155672
R960 VTAIL.n404 VTAIL.n363 0.155672
R961 VTAIL.n404 VTAIL.n403 0.155672
R962 VTAIL.n403 VTAIL.n367 0.155672
R963 VTAIL.n396 VTAIL.n367 0.155672
R964 VTAIL.n396 VTAIL.n395 0.155672
R965 VTAIL.n395 VTAIL.n371 0.155672
R966 VTAIL.n388 VTAIL.n371 0.155672
R967 VTAIL.n388 VTAIL.n387 0.155672
R968 VTAIL.n387 VTAIL.n375 0.155672
R969 VTAIL.n380 VTAIL.n375 0.155672
R970 VTAIL.n350 VTAIL.n349 0.155672
R971 VTAIL.n349 VTAIL.n289 0.155672
R972 VTAIL.n342 VTAIL.n289 0.155672
R973 VTAIL.n342 VTAIL.n341 0.155672
R974 VTAIL.n341 VTAIL.n293 0.155672
R975 VTAIL.n334 VTAIL.n293 0.155672
R976 VTAIL.n334 VTAIL.n333 0.155672
R977 VTAIL.n333 VTAIL.n297 0.155672
R978 VTAIL.n326 VTAIL.n297 0.155672
R979 VTAIL.n326 VTAIL.n325 0.155672
R980 VTAIL.n325 VTAIL.n301 0.155672
R981 VTAIL.n318 VTAIL.n301 0.155672
R982 VTAIL.n318 VTAIL.n317 0.155672
R983 VTAIL.n317 VTAIL.n305 0.155672
R984 VTAIL.n310 VTAIL.n305 0.155672
R985 VTAIL.n278 VTAIL.n277 0.155672
R986 VTAIL.n277 VTAIL.n217 0.155672
R987 VTAIL.n270 VTAIL.n217 0.155672
R988 VTAIL.n270 VTAIL.n269 0.155672
R989 VTAIL.n269 VTAIL.n221 0.155672
R990 VTAIL.n262 VTAIL.n221 0.155672
R991 VTAIL.n262 VTAIL.n261 0.155672
R992 VTAIL.n261 VTAIL.n225 0.155672
R993 VTAIL.n254 VTAIL.n225 0.155672
R994 VTAIL.n254 VTAIL.n253 0.155672
R995 VTAIL.n253 VTAIL.n229 0.155672
R996 VTAIL.n246 VTAIL.n229 0.155672
R997 VTAIL.n246 VTAIL.n245 0.155672
R998 VTAIL.n245 VTAIL.n233 0.155672
R999 VTAIL.n238 VTAIL.n233 0.155672
R1000 VTAIL VTAIL.n1 0.0586897
R1001 VP.n26 VP.n25 161.3
R1002 VP.n27 VP.n22 161.3
R1003 VP.n29 VP.n28 161.3
R1004 VP.n30 VP.n21 161.3
R1005 VP.n32 VP.n31 161.3
R1006 VP.n33 VP.n20 161.3
R1007 VP.n35 VP.n34 161.3
R1008 VP.n36 VP.n19 161.3
R1009 VP.n39 VP.n38 161.3
R1010 VP.n40 VP.n18 161.3
R1011 VP.n42 VP.n41 161.3
R1012 VP.n43 VP.n17 161.3
R1013 VP.n45 VP.n44 161.3
R1014 VP.n46 VP.n16 161.3
R1015 VP.n48 VP.n47 161.3
R1016 VP.n49 VP.n15 161.3
R1017 VP.n51 VP.n50 161.3
R1018 VP.n95 VP.n94 161.3
R1019 VP.n93 VP.n1 161.3
R1020 VP.n92 VP.n91 161.3
R1021 VP.n90 VP.n2 161.3
R1022 VP.n89 VP.n88 161.3
R1023 VP.n87 VP.n3 161.3
R1024 VP.n86 VP.n85 161.3
R1025 VP.n84 VP.n4 161.3
R1026 VP.n83 VP.n82 161.3
R1027 VP.n80 VP.n5 161.3
R1028 VP.n79 VP.n78 161.3
R1029 VP.n77 VP.n6 161.3
R1030 VP.n76 VP.n75 161.3
R1031 VP.n74 VP.n7 161.3
R1032 VP.n73 VP.n72 161.3
R1033 VP.n71 VP.n8 161.3
R1034 VP.n70 VP.n69 161.3
R1035 VP.n67 VP.n9 161.3
R1036 VP.n66 VP.n65 161.3
R1037 VP.n64 VP.n10 161.3
R1038 VP.n63 VP.n62 161.3
R1039 VP.n61 VP.n11 161.3
R1040 VP.n60 VP.n59 161.3
R1041 VP.n58 VP.n12 161.3
R1042 VP.n57 VP.n56 161.3
R1043 VP.n55 VP.n13 161.3
R1044 VP.n23 VP.t2 111.776
R1045 VP.n54 VP.n53 87.7864
R1046 VP.n96 VP.n0 87.7864
R1047 VP.n52 VP.n14 87.7864
R1048 VP.n54 VP.t3 78.9638
R1049 VP.n68 VP.t1 78.9638
R1050 VP.n81 VP.t6 78.9638
R1051 VP.n0 VP.t4 78.9638
R1052 VP.n14 VP.t5 78.9638
R1053 VP.n37 VP.t0 78.9638
R1054 VP.n24 VP.t7 78.9638
R1055 VP.n24 VP.n23 58.1068
R1056 VP.n53 VP.n52 57.4162
R1057 VP.n75 VP.n74 56.5617
R1058 VP.n31 VP.n30 56.5617
R1059 VP.n62 VP.n61 45.4209
R1060 VP.n88 VP.n87 45.4209
R1061 VP.n44 VP.n43 45.4209
R1062 VP.n61 VP.n60 35.7332
R1063 VP.n88 VP.n2 35.7332
R1064 VP.n44 VP.n16 35.7332
R1065 VP.n56 VP.n55 24.5923
R1066 VP.n56 VP.n12 24.5923
R1067 VP.n60 VP.n12 24.5923
R1068 VP.n62 VP.n10 24.5923
R1069 VP.n66 VP.n10 24.5923
R1070 VP.n67 VP.n66 24.5923
R1071 VP.n69 VP.n8 24.5923
R1072 VP.n73 VP.n8 24.5923
R1073 VP.n74 VP.n73 24.5923
R1074 VP.n75 VP.n6 24.5923
R1075 VP.n79 VP.n6 24.5923
R1076 VP.n80 VP.n79 24.5923
R1077 VP.n82 VP.n4 24.5923
R1078 VP.n86 VP.n4 24.5923
R1079 VP.n87 VP.n86 24.5923
R1080 VP.n92 VP.n2 24.5923
R1081 VP.n93 VP.n92 24.5923
R1082 VP.n94 VP.n93 24.5923
R1083 VP.n48 VP.n16 24.5923
R1084 VP.n49 VP.n48 24.5923
R1085 VP.n50 VP.n49 24.5923
R1086 VP.n31 VP.n20 24.5923
R1087 VP.n35 VP.n20 24.5923
R1088 VP.n36 VP.n35 24.5923
R1089 VP.n38 VP.n18 24.5923
R1090 VP.n42 VP.n18 24.5923
R1091 VP.n43 VP.n42 24.5923
R1092 VP.n25 VP.n22 24.5923
R1093 VP.n29 VP.n22 24.5923
R1094 VP.n30 VP.n29 24.5923
R1095 VP.n69 VP.n68 17.2148
R1096 VP.n81 VP.n80 17.2148
R1097 VP.n37 VP.n36 17.2148
R1098 VP.n25 VP.n24 17.2148
R1099 VP.n68 VP.n67 7.37805
R1100 VP.n82 VP.n81 7.37805
R1101 VP.n38 VP.n37 7.37805
R1102 VP.n26 VP.n23 2.46315
R1103 VP.n55 VP.n54 2.45968
R1104 VP.n94 VP.n0 2.45968
R1105 VP.n50 VP.n14 2.45968
R1106 VP.n52 VP.n51 0.354861
R1107 VP.n53 VP.n13 0.354861
R1108 VP.n96 VP.n95 0.354861
R1109 VP VP.n96 0.267071
R1110 VP.n27 VP.n26 0.189894
R1111 VP.n28 VP.n27 0.189894
R1112 VP.n28 VP.n21 0.189894
R1113 VP.n32 VP.n21 0.189894
R1114 VP.n33 VP.n32 0.189894
R1115 VP.n34 VP.n33 0.189894
R1116 VP.n34 VP.n19 0.189894
R1117 VP.n39 VP.n19 0.189894
R1118 VP.n40 VP.n39 0.189894
R1119 VP.n41 VP.n40 0.189894
R1120 VP.n41 VP.n17 0.189894
R1121 VP.n45 VP.n17 0.189894
R1122 VP.n46 VP.n45 0.189894
R1123 VP.n47 VP.n46 0.189894
R1124 VP.n47 VP.n15 0.189894
R1125 VP.n51 VP.n15 0.189894
R1126 VP.n57 VP.n13 0.189894
R1127 VP.n58 VP.n57 0.189894
R1128 VP.n59 VP.n58 0.189894
R1129 VP.n59 VP.n11 0.189894
R1130 VP.n63 VP.n11 0.189894
R1131 VP.n64 VP.n63 0.189894
R1132 VP.n65 VP.n64 0.189894
R1133 VP.n65 VP.n9 0.189894
R1134 VP.n70 VP.n9 0.189894
R1135 VP.n71 VP.n70 0.189894
R1136 VP.n72 VP.n71 0.189894
R1137 VP.n72 VP.n7 0.189894
R1138 VP.n76 VP.n7 0.189894
R1139 VP.n77 VP.n76 0.189894
R1140 VP.n78 VP.n77 0.189894
R1141 VP.n78 VP.n5 0.189894
R1142 VP.n83 VP.n5 0.189894
R1143 VP.n84 VP.n83 0.189894
R1144 VP.n85 VP.n84 0.189894
R1145 VP.n85 VP.n3 0.189894
R1146 VP.n89 VP.n3 0.189894
R1147 VP.n90 VP.n89 0.189894
R1148 VP.n91 VP.n90 0.189894
R1149 VP.n91 VP.n1 0.189894
R1150 VP.n95 VP.n1 0.189894
R1151 VDD1 VDD1.n0 78.4031
R1152 VDD1.n3 VDD1.n2 78.2886
R1153 VDD1.n3 VDD1.n1 78.2886
R1154 VDD1.n5 VDD1.n4 76.5335
R1155 VDD1.n5 VDD1.n3 51.5224
R1156 VDD1.n4 VDD1.t7 2.56399
R1157 VDD1.n4 VDD1.t2 2.56399
R1158 VDD1.n0 VDD1.t5 2.56399
R1159 VDD1.n0 VDD1.t0 2.56399
R1160 VDD1.n2 VDD1.t1 2.56399
R1161 VDD1.n2 VDD1.t3 2.56399
R1162 VDD1.n1 VDD1.t4 2.56399
R1163 VDD1.n1 VDD1.t6 2.56399
R1164 VDD1 VDD1.n5 1.75266
R1165 B.n710 B.n89 585
R1166 B.n712 B.n711 585
R1167 B.n713 B.n88 585
R1168 B.n715 B.n714 585
R1169 B.n716 B.n87 585
R1170 B.n718 B.n717 585
R1171 B.n719 B.n86 585
R1172 B.n721 B.n720 585
R1173 B.n722 B.n85 585
R1174 B.n724 B.n723 585
R1175 B.n725 B.n84 585
R1176 B.n727 B.n726 585
R1177 B.n728 B.n83 585
R1178 B.n730 B.n729 585
R1179 B.n731 B.n82 585
R1180 B.n733 B.n732 585
R1181 B.n734 B.n81 585
R1182 B.n736 B.n735 585
R1183 B.n737 B.n80 585
R1184 B.n739 B.n738 585
R1185 B.n740 B.n79 585
R1186 B.n742 B.n741 585
R1187 B.n743 B.n78 585
R1188 B.n745 B.n744 585
R1189 B.n746 B.n77 585
R1190 B.n748 B.n747 585
R1191 B.n749 B.n76 585
R1192 B.n751 B.n750 585
R1193 B.n752 B.n75 585
R1194 B.n754 B.n753 585
R1195 B.n755 B.n74 585
R1196 B.n757 B.n756 585
R1197 B.n758 B.n73 585
R1198 B.n760 B.n759 585
R1199 B.n761 B.n72 585
R1200 B.n763 B.n762 585
R1201 B.n764 B.n71 585
R1202 B.n766 B.n765 585
R1203 B.n767 B.n70 585
R1204 B.n769 B.n768 585
R1205 B.n770 B.n69 585
R1206 B.n772 B.n771 585
R1207 B.n773 B.n68 585
R1208 B.n775 B.n774 585
R1209 B.n777 B.n65 585
R1210 B.n779 B.n778 585
R1211 B.n780 B.n64 585
R1212 B.n782 B.n781 585
R1213 B.n783 B.n63 585
R1214 B.n785 B.n784 585
R1215 B.n786 B.n62 585
R1216 B.n788 B.n787 585
R1217 B.n789 B.n59 585
R1218 B.n792 B.n791 585
R1219 B.n793 B.n58 585
R1220 B.n795 B.n794 585
R1221 B.n796 B.n57 585
R1222 B.n798 B.n797 585
R1223 B.n799 B.n56 585
R1224 B.n801 B.n800 585
R1225 B.n802 B.n55 585
R1226 B.n804 B.n803 585
R1227 B.n805 B.n54 585
R1228 B.n807 B.n806 585
R1229 B.n808 B.n53 585
R1230 B.n810 B.n809 585
R1231 B.n811 B.n52 585
R1232 B.n813 B.n812 585
R1233 B.n814 B.n51 585
R1234 B.n816 B.n815 585
R1235 B.n817 B.n50 585
R1236 B.n819 B.n818 585
R1237 B.n820 B.n49 585
R1238 B.n822 B.n821 585
R1239 B.n823 B.n48 585
R1240 B.n825 B.n824 585
R1241 B.n826 B.n47 585
R1242 B.n828 B.n827 585
R1243 B.n829 B.n46 585
R1244 B.n831 B.n830 585
R1245 B.n832 B.n45 585
R1246 B.n834 B.n833 585
R1247 B.n835 B.n44 585
R1248 B.n837 B.n836 585
R1249 B.n838 B.n43 585
R1250 B.n840 B.n839 585
R1251 B.n841 B.n42 585
R1252 B.n843 B.n842 585
R1253 B.n844 B.n41 585
R1254 B.n846 B.n845 585
R1255 B.n847 B.n40 585
R1256 B.n849 B.n848 585
R1257 B.n850 B.n39 585
R1258 B.n852 B.n851 585
R1259 B.n853 B.n38 585
R1260 B.n855 B.n854 585
R1261 B.n856 B.n37 585
R1262 B.n709 B.n708 585
R1263 B.n707 B.n90 585
R1264 B.n706 B.n705 585
R1265 B.n704 B.n91 585
R1266 B.n703 B.n702 585
R1267 B.n701 B.n92 585
R1268 B.n700 B.n699 585
R1269 B.n698 B.n93 585
R1270 B.n697 B.n696 585
R1271 B.n695 B.n94 585
R1272 B.n694 B.n693 585
R1273 B.n692 B.n95 585
R1274 B.n691 B.n690 585
R1275 B.n689 B.n96 585
R1276 B.n688 B.n687 585
R1277 B.n686 B.n97 585
R1278 B.n685 B.n684 585
R1279 B.n683 B.n98 585
R1280 B.n682 B.n681 585
R1281 B.n680 B.n99 585
R1282 B.n679 B.n678 585
R1283 B.n677 B.n100 585
R1284 B.n676 B.n675 585
R1285 B.n674 B.n101 585
R1286 B.n673 B.n672 585
R1287 B.n671 B.n102 585
R1288 B.n670 B.n669 585
R1289 B.n668 B.n103 585
R1290 B.n667 B.n666 585
R1291 B.n665 B.n104 585
R1292 B.n664 B.n663 585
R1293 B.n662 B.n105 585
R1294 B.n661 B.n660 585
R1295 B.n659 B.n106 585
R1296 B.n658 B.n657 585
R1297 B.n656 B.n107 585
R1298 B.n655 B.n654 585
R1299 B.n653 B.n108 585
R1300 B.n652 B.n651 585
R1301 B.n650 B.n109 585
R1302 B.n649 B.n648 585
R1303 B.n647 B.n110 585
R1304 B.n646 B.n645 585
R1305 B.n644 B.n111 585
R1306 B.n643 B.n642 585
R1307 B.n641 B.n112 585
R1308 B.n640 B.n639 585
R1309 B.n638 B.n113 585
R1310 B.n637 B.n636 585
R1311 B.n635 B.n114 585
R1312 B.n634 B.n633 585
R1313 B.n632 B.n115 585
R1314 B.n631 B.n630 585
R1315 B.n629 B.n116 585
R1316 B.n628 B.n627 585
R1317 B.n626 B.n117 585
R1318 B.n625 B.n624 585
R1319 B.n623 B.n118 585
R1320 B.n622 B.n621 585
R1321 B.n620 B.n119 585
R1322 B.n619 B.n618 585
R1323 B.n617 B.n120 585
R1324 B.n616 B.n615 585
R1325 B.n614 B.n121 585
R1326 B.n613 B.n612 585
R1327 B.n611 B.n122 585
R1328 B.n610 B.n609 585
R1329 B.n608 B.n123 585
R1330 B.n607 B.n606 585
R1331 B.n605 B.n124 585
R1332 B.n604 B.n603 585
R1333 B.n602 B.n125 585
R1334 B.n601 B.n600 585
R1335 B.n599 B.n126 585
R1336 B.n598 B.n597 585
R1337 B.n596 B.n127 585
R1338 B.n595 B.n594 585
R1339 B.n593 B.n128 585
R1340 B.n592 B.n591 585
R1341 B.n590 B.n129 585
R1342 B.n589 B.n588 585
R1343 B.n587 B.n130 585
R1344 B.n586 B.n585 585
R1345 B.n584 B.n131 585
R1346 B.n583 B.n582 585
R1347 B.n581 B.n132 585
R1348 B.n580 B.n579 585
R1349 B.n578 B.n133 585
R1350 B.n577 B.n576 585
R1351 B.n575 B.n134 585
R1352 B.n574 B.n573 585
R1353 B.n572 B.n135 585
R1354 B.n571 B.n570 585
R1355 B.n569 B.n136 585
R1356 B.n568 B.n567 585
R1357 B.n566 B.n137 585
R1358 B.n565 B.n564 585
R1359 B.n563 B.n138 585
R1360 B.n562 B.n561 585
R1361 B.n560 B.n139 585
R1362 B.n559 B.n558 585
R1363 B.n557 B.n140 585
R1364 B.n556 B.n555 585
R1365 B.n554 B.n141 585
R1366 B.n553 B.n552 585
R1367 B.n551 B.n142 585
R1368 B.n550 B.n549 585
R1369 B.n548 B.n143 585
R1370 B.n547 B.n546 585
R1371 B.n545 B.n144 585
R1372 B.n544 B.n543 585
R1373 B.n542 B.n145 585
R1374 B.n541 B.n540 585
R1375 B.n539 B.n146 585
R1376 B.n538 B.n537 585
R1377 B.n536 B.n147 585
R1378 B.n535 B.n534 585
R1379 B.n533 B.n148 585
R1380 B.n532 B.n531 585
R1381 B.n530 B.n149 585
R1382 B.n529 B.n528 585
R1383 B.n527 B.n150 585
R1384 B.n526 B.n525 585
R1385 B.n524 B.n151 585
R1386 B.n523 B.n522 585
R1387 B.n521 B.n152 585
R1388 B.n520 B.n519 585
R1389 B.n518 B.n153 585
R1390 B.n517 B.n516 585
R1391 B.n515 B.n154 585
R1392 B.n514 B.n513 585
R1393 B.n512 B.n155 585
R1394 B.n511 B.n510 585
R1395 B.n509 B.n156 585
R1396 B.n508 B.n507 585
R1397 B.n506 B.n157 585
R1398 B.n505 B.n504 585
R1399 B.n503 B.n158 585
R1400 B.n502 B.n501 585
R1401 B.n500 B.n159 585
R1402 B.n499 B.n498 585
R1403 B.n352 B.n351 585
R1404 B.n353 B.n212 585
R1405 B.n355 B.n354 585
R1406 B.n356 B.n211 585
R1407 B.n358 B.n357 585
R1408 B.n359 B.n210 585
R1409 B.n361 B.n360 585
R1410 B.n362 B.n209 585
R1411 B.n364 B.n363 585
R1412 B.n365 B.n208 585
R1413 B.n367 B.n366 585
R1414 B.n368 B.n207 585
R1415 B.n370 B.n369 585
R1416 B.n371 B.n206 585
R1417 B.n373 B.n372 585
R1418 B.n374 B.n205 585
R1419 B.n376 B.n375 585
R1420 B.n377 B.n204 585
R1421 B.n379 B.n378 585
R1422 B.n380 B.n203 585
R1423 B.n382 B.n381 585
R1424 B.n383 B.n202 585
R1425 B.n385 B.n384 585
R1426 B.n386 B.n201 585
R1427 B.n388 B.n387 585
R1428 B.n389 B.n200 585
R1429 B.n391 B.n390 585
R1430 B.n392 B.n199 585
R1431 B.n394 B.n393 585
R1432 B.n395 B.n198 585
R1433 B.n397 B.n396 585
R1434 B.n398 B.n197 585
R1435 B.n400 B.n399 585
R1436 B.n401 B.n196 585
R1437 B.n403 B.n402 585
R1438 B.n404 B.n195 585
R1439 B.n406 B.n405 585
R1440 B.n407 B.n194 585
R1441 B.n409 B.n408 585
R1442 B.n410 B.n193 585
R1443 B.n412 B.n411 585
R1444 B.n413 B.n192 585
R1445 B.n415 B.n414 585
R1446 B.n416 B.n189 585
R1447 B.n419 B.n418 585
R1448 B.n420 B.n188 585
R1449 B.n422 B.n421 585
R1450 B.n423 B.n187 585
R1451 B.n425 B.n424 585
R1452 B.n426 B.n186 585
R1453 B.n428 B.n427 585
R1454 B.n429 B.n185 585
R1455 B.n431 B.n430 585
R1456 B.n433 B.n432 585
R1457 B.n434 B.n181 585
R1458 B.n436 B.n435 585
R1459 B.n437 B.n180 585
R1460 B.n439 B.n438 585
R1461 B.n440 B.n179 585
R1462 B.n442 B.n441 585
R1463 B.n443 B.n178 585
R1464 B.n445 B.n444 585
R1465 B.n446 B.n177 585
R1466 B.n448 B.n447 585
R1467 B.n449 B.n176 585
R1468 B.n451 B.n450 585
R1469 B.n452 B.n175 585
R1470 B.n454 B.n453 585
R1471 B.n455 B.n174 585
R1472 B.n457 B.n456 585
R1473 B.n458 B.n173 585
R1474 B.n460 B.n459 585
R1475 B.n461 B.n172 585
R1476 B.n463 B.n462 585
R1477 B.n464 B.n171 585
R1478 B.n466 B.n465 585
R1479 B.n467 B.n170 585
R1480 B.n469 B.n468 585
R1481 B.n470 B.n169 585
R1482 B.n472 B.n471 585
R1483 B.n473 B.n168 585
R1484 B.n475 B.n474 585
R1485 B.n476 B.n167 585
R1486 B.n478 B.n477 585
R1487 B.n479 B.n166 585
R1488 B.n481 B.n480 585
R1489 B.n482 B.n165 585
R1490 B.n484 B.n483 585
R1491 B.n485 B.n164 585
R1492 B.n487 B.n486 585
R1493 B.n488 B.n163 585
R1494 B.n490 B.n489 585
R1495 B.n491 B.n162 585
R1496 B.n493 B.n492 585
R1497 B.n494 B.n161 585
R1498 B.n496 B.n495 585
R1499 B.n497 B.n160 585
R1500 B.n350 B.n213 585
R1501 B.n349 B.n348 585
R1502 B.n347 B.n214 585
R1503 B.n346 B.n345 585
R1504 B.n344 B.n215 585
R1505 B.n343 B.n342 585
R1506 B.n341 B.n216 585
R1507 B.n340 B.n339 585
R1508 B.n338 B.n217 585
R1509 B.n337 B.n336 585
R1510 B.n335 B.n218 585
R1511 B.n334 B.n333 585
R1512 B.n332 B.n219 585
R1513 B.n331 B.n330 585
R1514 B.n329 B.n220 585
R1515 B.n328 B.n327 585
R1516 B.n326 B.n221 585
R1517 B.n325 B.n324 585
R1518 B.n323 B.n222 585
R1519 B.n322 B.n321 585
R1520 B.n320 B.n223 585
R1521 B.n319 B.n318 585
R1522 B.n317 B.n224 585
R1523 B.n316 B.n315 585
R1524 B.n314 B.n225 585
R1525 B.n313 B.n312 585
R1526 B.n311 B.n226 585
R1527 B.n310 B.n309 585
R1528 B.n308 B.n227 585
R1529 B.n307 B.n306 585
R1530 B.n305 B.n228 585
R1531 B.n304 B.n303 585
R1532 B.n302 B.n229 585
R1533 B.n301 B.n300 585
R1534 B.n299 B.n230 585
R1535 B.n298 B.n297 585
R1536 B.n296 B.n231 585
R1537 B.n295 B.n294 585
R1538 B.n293 B.n232 585
R1539 B.n292 B.n291 585
R1540 B.n290 B.n233 585
R1541 B.n289 B.n288 585
R1542 B.n287 B.n234 585
R1543 B.n286 B.n285 585
R1544 B.n284 B.n235 585
R1545 B.n283 B.n282 585
R1546 B.n281 B.n236 585
R1547 B.n280 B.n279 585
R1548 B.n278 B.n237 585
R1549 B.n277 B.n276 585
R1550 B.n275 B.n238 585
R1551 B.n274 B.n273 585
R1552 B.n272 B.n239 585
R1553 B.n271 B.n270 585
R1554 B.n269 B.n240 585
R1555 B.n268 B.n267 585
R1556 B.n266 B.n241 585
R1557 B.n265 B.n264 585
R1558 B.n263 B.n242 585
R1559 B.n262 B.n261 585
R1560 B.n260 B.n243 585
R1561 B.n259 B.n258 585
R1562 B.n257 B.n244 585
R1563 B.n256 B.n255 585
R1564 B.n254 B.n245 585
R1565 B.n253 B.n252 585
R1566 B.n251 B.n246 585
R1567 B.n250 B.n249 585
R1568 B.n248 B.n247 585
R1569 B.n2 B.n0 585
R1570 B.n961 B.n1 585
R1571 B.n960 B.n959 585
R1572 B.n958 B.n3 585
R1573 B.n957 B.n956 585
R1574 B.n955 B.n4 585
R1575 B.n954 B.n953 585
R1576 B.n952 B.n5 585
R1577 B.n951 B.n950 585
R1578 B.n949 B.n6 585
R1579 B.n948 B.n947 585
R1580 B.n946 B.n7 585
R1581 B.n945 B.n944 585
R1582 B.n943 B.n8 585
R1583 B.n942 B.n941 585
R1584 B.n940 B.n9 585
R1585 B.n939 B.n938 585
R1586 B.n937 B.n10 585
R1587 B.n936 B.n935 585
R1588 B.n934 B.n11 585
R1589 B.n933 B.n932 585
R1590 B.n931 B.n12 585
R1591 B.n930 B.n929 585
R1592 B.n928 B.n13 585
R1593 B.n927 B.n926 585
R1594 B.n925 B.n14 585
R1595 B.n924 B.n923 585
R1596 B.n922 B.n15 585
R1597 B.n921 B.n920 585
R1598 B.n919 B.n16 585
R1599 B.n918 B.n917 585
R1600 B.n916 B.n17 585
R1601 B.n915 B.n914 585
R1602 B.n913 B.n18 585
R1603 B.n912 B.n911 585
R1604 B.n910 B.n19 585
R1605 B.n909 B.n908 585
R1606 B.n907 B.n20 585
R1607 B.n906 B.n905 585
R1608 B.n904 B.n21 585
R1609 B.n903 B.n902 585
R1610 B.n901 B.n22 585
R1611 B.n900 B.n899 585
R1612 B.n898 B.n23 585
R1613 B.n897 B.n896 585
R1614 B.n895 B.n24 585
R1615 B.n894 B.n893 585
R1616 B.n892 B.n25 585
R1617 B.n891 B.n890 585
R1618 B.n889 B.n26 585
R1619 B.n888 B.n887 585
R1620 B.n886 B.n27 585
R1621 B.n885 B.n884 585
R1622 B.n883 B.n28 585
R1623 B.n882 B.n881 585
R1624 B.n880 B.n29 585
R1625 B.n879 B.n878 585
R1626 B.n877 B.n30 585
R1627 B.n876 B.n875 585
R1628 B.n874 B.n31 585
R1629 B.n873 B.n872 585
R1630 B.n871 B.n32 585
R1631 B.n870 B.n869 585
R1632 B.n868 B.n33 585
R1633 B.n867 B.n866 585
R1634 B.n865 B.n34 585
R1635 B.n864 B.n863 585
R1636 B.n862 B.n35 585
R1637 B.n861 B.n860 585
R1638 B.n859 B.n36 585
R1639 B.n858 B.n857 585
R1640 B.n963 B.n962 585
R1641 B.n182 B.t2 469.231
R1642 B.n66 B.t4 469.231
R1643 B.n190 B.t11 469.231
R1644 B.n60 B.t7 469.231
R1645 B.n352 B.n213 463.671
R1646 B.n858 B.n37 463.671
R1647 B.n498 B.n497 463.671
R1648 B.n708 B.n89 463.671
R1649 B.n183 B.t1 387.776
R1650 B.n67 B.t5 387.776
R1651 B.n191 B.t10 387.776
R1652 B.n61 B.t8 387.776
R1653 B.n182 B.t0 288.361
R1654 B.n190 B.t9 288.361
R1655 B.n60 B.t6 288.361
R1656 B.n66 B.t3 288.361
R1657 B.n348 B.n213 163.367
R1658 B.n348 B.n347 163.367
R1659 B.n347 B.n346 163.367
R1660 B.n346 B.n215 163.367
R1661 B.n342 B.n215 163.367
R1662 B.n342 B.n341 163.367
R1663 B.n341 B.n340 163.367
R1664 B.n340 B.n217 163.367
R1665 B.n336 B.n217 163.367
R1666 B.n336 B.n335 163.367
R1667 B.n335 B.n334 163.367
R1668 B.n334 B.n219 163.367
R1669 B.n330 B.n219 163.367
R1670 B.n330 B.n329 163.367
R1671 B.n329 B.n328 163.367
R1672 B.n328 B.n221 163.367
R1673 B.n324 B.n221 163.367
R1674 B.n324 B.n323 163.367
R1675 B.n323 B.n322 163.367
R1676 B.n322 B.n223 163.367
R1677 B.n318 B.n223 163.367
R1678 B.n318 B.n317 163.367
R1679 B.n317 B.n316 163.367
R1680 B.n316 B.n225 163.367
R1681 B.n312 B.n225 163.367
R1682 B.n312 B.n311 163.367
R1683 B.n311 B.n310 163.367
R1684 B.n310 B.n227 163.367
R1685 B.n306 B.n227 163.367
R1686 B.n306 B.n305 163.367
R1687 B.n305 B.n304 163.367
R1688 B.n304 B.n229 163.367
R1689 B.n300 B.n229 163.367
R1690 B.n300 B.n299 163.367
R1691 B.n299 B.n298 163.367
R1692 B.n298 B.n231 163.367
R1693 B.n294 B.n231 163.367
R1694 B.n294 B.n293 163.367
R1695 B.n293 B.n292 163.367
R1696 B.n292 B.n233 163.367
R1697 B.n288 B.n233 163.367
R1698 B.n288 B.n287 163.367
R1699 B.n287 B.n286 163.367
R1700 B.n286 B.n235 163.367
R1701 B.n282 B.n235 163.367
R1702 B.n282 B.n281 163.367
R1703 B.n281 B.n280 163.367
R1704 B.n280 B.n237 163.367
R1705 B.n276 B.n237 163.367
R1706 B.n276 B.n275 163.367
R1707 B.n275 B.n274 163.367
R1708 B.n274 B.n239 163.367
R1709 B.n270 B.n239 163.367
R1710 B.n270 B.n269 163.367
R1711 B.n269 B.n268 163.367
R1712 B.n268 B.n241 163.367
R1713 B.n264 B.n241 163.367
R1714 B.n264 B.n263 163.367
R1715 B.n263 B.n262 163.367
R1716 B.n262 B.n243 163.367
R1717 B.n258 B.n243 163.367
R1718 B.n258 B.n257 163.367
R1719 B.n257 B.n256 163.367
R1720 B.n256 B.n245 163.367
R1721 B.n252 B.n245 163.367
R1722 B.n252 B.n251 163.367
R1723 B.n251 B.n250 163.367
R1724 B.n250 B.n247 163.367
R1725 B.n247 B.n2 163.367
R1726 B.n962 B.n2 163.367
R1727 B.n962 B.n961 163.367
R1728 B.n961 B.n960 163.367
R1729 B.n960 B.n3 163.367
R1730 B.n956 B.n3 163.367
R1731 B.n956 B.n955 163.367
R1732 B.n955 B.n954 163.367
R1733 B.n954 B.n5 163.367
R1734 B.n950 B.n5 163.367
R1735 B.n950 B.n949 163.367
R1736 B.n949 B.n948 163.367
R1737 B.n948 B.n7 163.367
R1738 B.n944 B.n7 163.367
R1739 B.n944 B.n943 163.367
R1740 B.n943 B.n942 163.367
R1741 B.n942 B.n9 163.367
R1742 B.n938 B.n9 163.367
R1743 B.n938 B.n937 163.367
R1744 B.n937 B.n936 163.367
R1745 B.n936 B.n11 163.367
R1746 B.n932 B.n11 163.367
R1747 B.n932 B.n931 163.367
R1748 B.n931 B.n930 163.367
R1749 B.n930 B.n13 163.367
R1750 B.n926 B.n13 163.367
R1751 B.n926 B.n925 163.367
R1752 B.n925 B.n924 163.367
R1753 B.n924 B.n15 163.367
R1754 B.n920 B.n15 163.367
R1755 B.n920 B.n919 163.367
R1756 B.n919 B.n918 163.367
R1757 B.n918 B.n17 163.367
R1758 B.n914 B.n17 163.367
R1759 B.n914 B.n913 163.367
R1760 B.n913 B.n912 163.367
R1761 B.n912 B.n19 163.367
R1762 B.n908 B.n19 163.367
R1763 B.n908 B.n907 163.367
R1764 B.n907 B.n906 163.367
R1765 B.n906 B.n21 163.367
R1766 B.n902 B.n21 163.367
R1767 B.n902 B.n901 163.367
R1768 B.n901 B.n900 163.367
R1769 B.n900 B.n23 163.367
R1770 B.n896 B.n23 163.367
R1771 B.n896 B.n895 163.367
R1772 B.n895 B.n894 163.367
R1773 B.n894 B.n25 163.367
R1774 B.n890 B.n25 163.367
R1775 B.n890 B.n889 163.367
R1776 B.n889 B.n888 163.367
R1777 B.n888 B.n27 163.367
R1778 B.n884 B.n27 163.367
R1779 B.n884 B.n883 163.367
R1780 B.n883 B.n882 163.367
R1781 B.n882 B.n29 163.367
R1782 B.n878 B.n29 163.367
R1783 B.n878 B.n877 163.367
R1784 B.n877 B.n876 163.367
R1785 B.n876 B.n31 163.367
R1786 B.n872 B.n31 163.367
R1787 B.n872 B.n871 163.367
R1788 B.n871 B.n870 163.367
R1789 B.n870 B.n33 163.367
R1790 B.n866 B.n33 163.367
R1791 B.n866 B.n865 163.367
R1792 B.n865 B.n864 163.367
R1793 B.n864 B.n35 163.367
R1794 B.n860 B.n35 163.367
R1795 B.n860 B.n859 163.367
R1796 B.n859 B.n858 163.367
R1797 B.n353 B.n352 163.367
R1798 B.n354 B.n353 163.367
R1799 B.n354 B.n211 163.367
R1800 B.n358 B.n211 163.367
R1801 B.n359 B.n358 163.367
R1802 B.n360 B.n359 163.367
R1803 B.n360 B.n209 163.367
R1804 B.n364 B.n209 163.367
R1805 B.n365 B.n364 163.367
R1806 B.n366 B.n365 163.367
R1807 B.n366 B.n207 163.367
R1808 B.n370 B.n207 163.367
R1809 B.n371 B.n370 163.367
R1810 B.n372 B.n371 163.367
R1811 B.n372 B.n205 163.367
R1812 B.n376 B.n205 163.367
R1813 B.n377 B.n376 163.367
R1814 B.n378 B.n377 163.367
R1815 B.n378 B.n203 163.367
R1816 B.n382 B.n203 163.367
R1817 B.n383 B.n382 163.367
R1818 B.n384 B.n383 163.367
R1819 B.n384 B.n201 163.367
R1820 B.n388 B.n201 163.367
R1821 B.n389 B.n388 163.367
R1822 B.n390 B.n389 163.367
R1823 B.n390 B.n199 163.367
R1824 B.n394 B.n199 163.367
R1825 B.n395 B.n394 163.367
R1826 B.n396 B.n395 163.367
R1827 B.n396 B.n197 163.367
R1828 B.n400 B.n197 163.367
R1829 B.n401 B.n400 163.367
R1830 B.n402 B.n401 163.367
R1831 B.n402 B.n195 163.367
R1832 B.n406 B.n195 163.367
R1833 B.n407 B.n406 163.367
R1834 B.n408 B.n407 163.367
R1835 B.n408 B.n193 163.367
R1836 B.n412 B.n193 163.367
R1837 B.n413 B.n412 163.367
R1838 B.n414 B.n413 163.367
R1839 B.n414 B.n189 163.367
R1840 B.n419 B.n189 163.367
R1841 B.n420 B.n419 163.367
R1842 B.n421 B.n420 163.367
R1843 B.n421 B.n187 163.367
R1844 B.n425 B.n187 163.367
R1845 B.n426 B.n425 163.367
R1846 B.n427 B.n426 163.367
R1847 B.n427 B.n185 163.367
R1848 B.n431 B.n185 163.367
R1849 B.n432 B.n431 163.367
R1850 B.n432 B.n181 163.367
R1851 B.n436 B.n181 163.367
R1852 B.n437 B.n436 163.367
R1853 B.n438 B.n437 163.367
R1854 B.n438 B.n179 163.367
R1855 B.n442 B.n179 163.367
R1856 B.n443 B.n442 163.367
R1857 B.n444 B.n443 163.367
R1858 B.n444 B.n177 163.367
R1859 B.n448 B.n177 163.367
R1860 B.n449 B.n448 163.367
R1861 B.n450 B.n449 163.367
R1862 B.n450 B.n175 163.367
R1863 B.n454 B.n175 163.367
R1864 B.n455 B.n454 163.367
R1865 B.n456 B.n455 163.367
R1866 B.n456 B.n173 163.367
R1867 B.n460 B.n173 163.367
R1868 B.n461 B.n460 163.367
R1869 B.n462 B.n461 163.367
R1870 B.n462 B.n171 163.367
R1871 B.n466 B.n171 163.367
R1872 B.n467 B.n466 163.367
R1873 B.n468 B.n467 163.367
R1874 B.n468 B.n169 163.367
R1875 B.n472 B.n169 163.367
R1876 B.n473 B.n472 163.367
R1877 B.n474 B.n473 163.367
R1878 B.n474 B.n167 163.367
R1879 B.n478 B.n167 163.367
R1880 B.n479 B.n478 163.367
R1881 B.n480 B.n479 163.367
R1882 B.n480 B.n165 163.367
R1883 B.n484 B.n165 163.367
R1884 B.n485 B.n484 163.367
R1885 B.n486 B.n485 163.367
R1886 B.n486 B.n163 163.367
R1887 B.n490 B.n163 163.367
R1888 B.n491 B.n490 163.367
R1889 B.n492 B.n491 163.367
R1890 B.n492 B.n161 163.367
R1891 B.n496 B.n161 163.367
R1892 B.n497 B.n496 163.367
R1893 B.n498 B.n159 163.367
R1894 B.n502 B.n159 163.367
R1895 B.n503 B.n502 163.367
R1896 B.n504 B.n503 163.367
R1897 B.n504 B.n157 163.367
R1898 B.n508 B.n157 163.367
R1899 B.n509 B.n508 163.367
R1900 B.n510 B.n509 163.367
R1901 B.n510 B.n155 163.367
R1902 B.n514 B.n155 163.367
R1903 B.n515 B.n514 163.367
R1904 B.n516 B.n515 163.367
R1905 B.n516 B.n153 163.367
R1906 B.n520 B.n153 163.367
R1907 B.n521 B.n520 163.367
R1908 B.n522 B.n521 163.367
R1909 B.n522 B.n151 163.367
R1910 B.n526 B.n151 163.367
R1911 B.n527 B.n526 163.367
R1912 B.n528 B.n527 163.367
R1913 B.n528 B.n149 163.367
R1914 B.n532 B.n149 163.367
R1915 B.n533 B.n532 163.367
R1916 B.n534 B.n533 163.367
R1917 B.n534 B.n147 163.367
R1918 B.n538 B.n147 163.367
R1919 B.n539 B.n538 163.367
R1920 B.n540 B.n539 163.367
R1921 B.n540 B.n145 163.367
R1922 B.n544 B.n145 163.367
R1923 B.n545 B.n544 163.367
R1924 B.n546 B.n545 163.367
R1925 B.n546 B.n143 163.367
R1926 B.n550 B.n143 163.367
R1927 B.n551 B.n550 163.367
R1928 B.n552 B.n551 163.367
R1929 B.n552 B.n141 163.367
R1930 B.n556 B.n141 163.367
R1931 B.n557 B.n556 163.367
R1932 B.n558 B.n557 163.367
R1933 B.n558 B.n139 163.367
R1934 B.n562 B.n139 163.367
R1935 B.n563 B.n562 163.367
R1936 B.n564 B.n563 163.367
R1937 B.n564 B.n137 163.367
R1938 B.n568 B.n137 163.367
R1939 B.n569 B.n568 163.367
R1940 B.n570 B.n569 163.367
R1941 B.n570 B.n135 163.367
R1942 B.n574 B.n135 163.367
R1943 B.n575 B.n574 163.367
R1944 B.n576 B.n575 163.367
R1945 B.n576 B.n133 163.367
R1946 B.n580 B.n133 163.367
R1947 B.n581 B.n580 163.367
R1948 B.n582 B.n581 163.367
R1949 B.n582 B.n131 163.367
R1950 B.n586 B.n131 163.367
R1951 B.n587 B.n586 163.367
R1952 B.n588 B.n587 163.367
R1953 B.n588 B.n129 163.367
R1954 B.n592 B.n129 163.367
R1955 B.n593 B.n592 163.367
R1956 B.n594 B.n593 163.367
R1957 B.n594 B.n127 163.367
R1958 B.n598 B.n127 163.367
R1959 B.n599 B.n598 163.367
R1960 B.n600 B.n599 163.367
R1961 B.n600 B.n125 163.367
R1962 B.n604 B.n125 163.367
R1963 B.n605 B.n604 163.367
R1964 B.n606 B.n605 163.367
R1965 B.n606 B.n123 163.367
R1966 B.n610 B.n123 163.367
R1967 B.n611 B.n610 163.367
R1968 B.n612 B.n611 163.367
R1969 B.n612 B.n121 163.367
R1970 B.n616 B.n121 163.367
R1971 B.n617 B.n616 163.367
R1972 B.n618 B.n617 163.367
R1973 B.n618 B.n119 163.367
R1974 B.n622 B.n119 163.367
R1975 B.n623 B.n622 163.367
R1976 B.n624 B.n623 163.367
R1977 B.n624 B.n117 163.367
R1978 B.n628 B.n117 163.367
R1979 B.n629 B.n628 163.367
R1980 B.n630 B.n629 163.367
R1981 B.n630 B.n115 163.367
R1982 B.n634 B.n115 163.367
R1983 B.n635 B.n634 163.367
R1984 B.n636 B.n635 163.367
R1985 B.n636 B.n113 163.367
R1986 B.n640 B.n113 163.367
R1987 B.n641 B.n640 163.367
R1988 B.n642 B.n641 163.367
R1989 B.n642 B.n111 163.367
R1990 B.n646 B.n111 163.367
R1991 B.n647 B.n646 163.367
R1992 B.n648 B.n647 163.367
R1993 B.n648 B.n109 163.367
R1994 B.n652 B.n109 163.367
R1995 B.n653 B.n652 163.367
R1996 B.n654 B.n653 163.367
R1997 B.n654 B.n107 163.367
R1998 B.n658 B.n107 163.367
R1999 B.n659 B.n658 163.367
R2000 B.n660 B.n659 163.367
R2001 B.n660 B.n105 163.367
R2002 B.n664 B.n105 163.367
R2003 B.n665 B.n664 163.367
R2004 B.n666 B.n665 163.367
R2005 B.n666 B.n103 163.367
R2006 B.n670 B.n103 163.367
R2007 B.n671 B.n670 163.367
R2008 B.n672 B.n671 163.367
R2009 B.n672 B.n101 163.367
R2010 B.n676 B.n101 163.367
R2011 B.n677 B.n676 163.367
R2012 B.n678 B.n677 163.367
R2013 B.n678 B.n99 163.367
R2014 B.n682 B.n99 163.367
R2015 B.n683 B.n682 163.367
R2016 B.n684 B.n683 163.367
R2017 B.n684 B.n97 163.367
R2018 B.n688 B.n97 163.367
R2019 B.n689 B.n688 163.367
R2020 B.n690 B.n689 163.367
R2021 B.n690 B.n95 163.367
R2022 B.n694 B.n95 163.367
R2023 B.n695 B.n694 163.367
R2024 B.n696 B.n695 163.367
R2025 B.n696 B.n93 163.367
R2026 B.n700 B.n93 163.367
R2027 B.n701 B.n700 163.367
R2028 B.n702 B.n701 163.367
R2029 B.n702 B.n91 163.367
R2030 B.n706 B.n91 163.367
R2031 B.n707 B.n706 163.367
R2032 B.n708 B.n707 163.367
R2033 B.n854 B.n37 163.367
R2034 B.n854 B.n853 163.367
R2035 B.n853 B.n852 163.367
R2036 B.n852 B.n39 163.367
R2037 B.n848 B.n39 163.367
R2038 B.n848 B.n847 163.367
R2039 B.n847 B.n846 163.367
R2040 B.n846 B.n41 163.367
R2041 B.n842 B.n41 163.367
R2042 B.n842 B.n841 163.367
R2043 B.n841 B.n840 163.367
R2044 B.n840 B.n43 163.367
R2045 B.n836 B.n43 163.367
R2046 B.n836 B.n835 163.367
R2047 B.n835 B.n834 163.367
R2048 B.n834 B.n45 163.367
R2049 B.n830 B.n45 163.367
R2050 B.n830 B.n829 163.367
R2051 B.n829 B.n828 163.367
R2052 B.n828 B.n47 163.367
R2053 B.n824 B.n47 163.367
R2054 B.n824 B.n823 163.367
R2055 B.n823 B.n822 163.367
R2056 B.n822 B.n49 163.367
R2057 B.n818 B.n49 163.367
R2058 B.n818 B.n817 163.367
R2059 B.n817 B.n816 163.367
R2060 B.n816 B.n51 163.367
R2061 B.n812 B.n51 163.367
R2062 B.n812 B.n811 163.367
R2063 B.n811 B.n810 163.367
R2064 B.n810 B.n53 163.367
R2065 B.n806 B.n53 163.367
R2066 B.n806 B.n805 163.367
R2067 B.n805 B.n804 163.367
R2068 B.n804 B.n55 163.367
R2069 B.n800 B.n55 163.367
R2070 B.n800 B.n799 163.367
R2071 B.n799 B.n798 163.367
R2072 B.n798 B.n57 163.367
R2073 B.n794 B.n57 163.367
R2074 B.n794 B.n793 163.367
R2075 B.n793 B.n792 163.367
R2076 B.n792 B.n59 163.367
R2077 B.n787 B.n59 163.367
R2078 B.n787 B.n786 163.367
R2079 B.n786 B.n785 163.367
R2080 B.n785 B.n63 163.367
R2081 B.n781 B.n63 163.367
R2082 B.n781 B.n780 163.367
R2083 B.n780 B.n779 163.367
R2084 B.n779 B.n65 163.367
R2085 B.n774 B.n65 163.367
R2086 B.n774 B.n773 163.367
R2087 B.n773 B.n772 163.367
R2088 B.n772 B.n69 163.367
R2089 B.n768 B.n69 163.367
R2090 B.n768 B.n767 163.367
R2091 B.n767 B.n766 163.367
R2092 B.n766 B.n71 163.367
R2093 B.n762 B.n71 163.367
R2094 B.n762 B.n761 163.367
R2095 B.n761 B.n760 163.367
R2096 B.n760 B.n73 163.367
R2097 B.n756 B.n73 163.367
R2098 B.n756 B.n755 163.367
R2099 B.n755 B.n754 163.367
R2100 B.n754 B.n75 163.367
R2101 B.n750 B.n75 163.367
R2102 B.n750 B.n749 163.367
R2103 B.n749 B.n748 163.367
R2104 B.n748 B.n77 163.367
R2105 B.n744 B.n77 163.367
R2106 B.n744 B.n743 163.367
R2107 B.n743 B.n742 163.367
R2108 B.n742 B.n79 163.367
R2109 B.n738 B.n79 163.367
R2110 B.n738 B.n737 163.367
R2111 B.n737 B.n736 163.367
R2112 B.n736 B.n81 163.367
R2113 B.n732 B.n81 163.367
R2114 B.n732 B.n731 163.367
R2115 B.n731 B.n730 163.367
R2116 B.n730 B.n83 163.367
R2117 B.n726 B.n83 163.367
R2118 B.n726 B.n725 163.367
R2119 B.n725 B.n724 163.367
R2120 B.n724 B.n85 163.367
R2121 B.n720 B.n85 163.367
R2122 B.n720 B.n719 163.367
R2123 B.n719 B.n718 163.367
R2124 B.n718 B.n87 163.367
R2125 B.n714 B.n87 163.367
R2126 B.n714 B.n713 163.367
R2127 B.n713 B.n712 163.367
R2128 B.n712 B.n89 163.367
R2129 B.n183 B.n182 81.455
R2130 B.n191 B.n190 81.455
R2131 B.n61 B.n60 81.455
R2132 B.n67 B.n66 81.455
R2133 B.n184 B.n183 59.5399
R2134 B.n417 B.n191 59.5399
R2135 B.n790 B.n61 59.5399
R2136 B.n776 B.n67 59.5399
R2137 B.n857 B.n856 30.1273
R2138 B.n710 B.n709 30.1273
R2139 B.n499 B.n160 30.1273
R2140 B.n351 B.n350 30.1273
R2141 B B.n963 18.0485
R2142 B.n856 B.n855 10.6151
R2143 B.n855 B.n38 10.6151
R2144 B.n851 B.n38 10.6151
R2145 B.n851 B.n850 10.6151
R2146 B.n850 B.n849 10.6151
R2147 B.n849 B.n40 10.6151
R2148 B.n845 B.n40 10.6151
R2149 B.n845 B.n844 10.6151
R2150 B.n844 B.n843 10.6151
R2151 B.n843 B.n42 10.6151
R2152 B.n839 B.n42 10.6151
R2153 B.n839 B.n838 10.6151
R2154 B.n838 B.n837 10.6151
R2155 B.n837 B.n44 10.6151
R2156 B.n833 B.n44 10.6151
R2157 B.n833 B.n832 10.6151
R2158 B.n832 B.n831 10.6151
R2159 B.n831 B.n46 10.6151
R2160 B.n827 B.n46 10.6151
R2161 B.n827 B.n826 10.6151
R2162 B.n826 B.n825 10.6151
R2163 B.n825 B.n48 10.6151
R2164 B.n821 B.n48 10.6151
R2165 B.n821 B.n820 10.6151
R2166 B.n820 B.n819 10.6151
R2167 B.n819 B.n50 10.6151
R2168 B.n815 B.n50 10.6151
R2169 B.n815 B.n814 10.6151
R2170 B.n814 B.n813 10.6151
R2171 B.n813 B.n52 10.6151
R2172 B.n809 B.n52 10.6151
R2173 B.n809 B.n808 10.6151
R2174 B.n808 B.n807 10.6151
R2175 B.n807 B.n54 10.6151
R2176 B.n803 B.n54 10.6151
R2177 B.n803 B.n802 10.6151
R2178 B.n802 B.n801 10.6151
R2179 B.n801 B.n56 10.6151
R2180 B.n797 B.n56 10.6151
R2181 B.n797 B.n796 10.6151
R2182 B.n796 B.n795 10.6151
R2183 B.n795 B.n58 10.6151
R2184 B.n791 B.n58 10.6151
R2185 B.n789 B.n788 10.6151
R2186 B.n788 B.n62 10.6151
R2187 B.n784 B.n62 10.6151
R2188 B.n784 B.n783 10.6151
R2189 B.n783 B.n782 10.6151
R2190 B.n782 B.n64 10.6151
R2191 B.n778 B.n64 10.6151
R2192 B.n778 B.n777 10.6151
R2193 B.n775 B.n68 10.6151
R2194 B.n771 B.n68 10.6151
R2195 B.n771 B.n770 10.6151
R2196 B.n770 B.n769 10.6151
R2197 B.n769 B.n70 10.6151
R2198 B.n765 B.n70 10.6151
R2199 B.n765 B.n764 10.6151
R2200 B.n764 B.n763 10.6151
R2201 B.n763 B.n72 10.6151
R2202 B.n759 B.n72 10.6151
R2203 B.n759 B.n758 10.6151
R2204 B.n758 B.n757 10.6151
R2205 B.n757 B.n74 10.6151
R2206 B.n753 B.n74 10.6151
R2207 B.n753 B.n752 10.6151
R2208 B.n752 B.n751 10.6151
R2209 B.n751 B.n76 10.6151
R2210 B.n747 B.n76 10.6151
R2211 B.n747 B.n746 10.6151
R2212 B.n746 B.n745 10.6151
R2213 B.n745 B.n78 10.6151
R2214 B.n741 B.n78 10.6151
R2215 B.n741 B.n740 10.6151
R2216 B.n740 B.n739 10.6151
R2217 B.n739 B.n80 10.6151
R2218 B.n735 B.n80 10.6151
R2219 B.n735 B.n734 10.6151
R2220 B.n734 B.n733 10.6151
R2221 B.n733 B.n82 10.6151
R2222 B.n729 B.n82 10.6151
R2223 B.n729 B.n728 10.6151
R2224 B.n728 B.n727 10.6151
R2225 B.n727 B.n84 10.6151
R2226 B.n723 B.n84 10.6151
R2227 B.n723 B.n722 10.6151
R2228 B.n722 B.n721 10.6151
R2229 B.n721 B.n86 10.6151
R2230 B.n717 B.n86 10.6151
R2231 B.n717 B.n716 10.6151
R2232 B.n716 B.n715 10.6151
R2233 B.n715 B.n88 10.6151
R2234 B.n711 B.n88 10.6151
R2235 B.n711 B.n710 10.6151
R2236 B.n500 B.n499 10.6151
R2237 B.n501 B.n500 10.6151
R2238 B.n501 B.n158 10.6151
R2239 B.n505 B.n158 10.6151
R2240 B.n506 B.n505 10.6151
R2241 B.n507 B.n506 10.6151
R2242 B.n507 B.n156 10.6151
R2243 B.n511 B.n156 10.6151
R2244 B.n512 B.n511 10.6151
R2245 B.n513 B.n512 10.6151
R2246 B.n513 B.n154 10.6151
R2247 B.n517 B.n154 10.6151
R2248 B.n518 B.n517 10.6151
R2249 B.n519 B.n518 10.6151
R2250 B.n519 B.n152 10.6151
R2251 B.n523 B.n152 10.6151
R2252 B.n524 B.n523 10.6151
R2253 B.n525 B.n524 10.6151
R2254 B.n525 B.n150 10.6151
R2255 B.n529 B.n150 10.6151
R2256 B.n530 B.n529 10.6151
R2257 B.n531 B.n530 10.6151
R2258 B.n531 B.n148 10.6151
R2259 B.n535 B.n148 10.6151
R2260 B.n536 B.n535 10.6151
R2261 B.n537 B.n536 10.6151
R2262 B.n537 B.n146 10.6151
R2263 B.n541 B.n146 10.6151
R2264 B.n542 B.n541 10.6151
R2265 B.n543 B.n542 10.6151
R2266 B.n543 B.n144 10.6151
R2267 B.n547 B.n144 10.6151
R2268 B.n548 B.n547 10.6151
R2269 B.n549 B.n548 10.6151
R2270 B.n549 B.n142 10.6151
R2271 B.n553 B.n142 10.6151
R2272 B.n554 B.n553 10.6151
R2273 B.n555 B.n554 10.6151
R2274 B.n555 B.n140 10.6151
R2275 B.n559 B.n140 10.6151
R2276 B.n560 B.n559 10.6151
R2277 B.n561 B.n560 10.6151
R2278 B.n561 B.n138 10.6151
R2279 B.n565 B.n138 10.6151
R2280 B.n566 B.n565 10.6151
R2281 B.n567 B.n566 10.6151
R2282 B.n567 B.n136 10.6151
R2283 B.n571 B.n136 10.6151
R2284 B.n572 B.n571 10.6151
R2285 B.n573 B.n572 10.6151
R2286 B.n573 B.n134 10.6151
R2287 B.n577 B.n134 10.6151
R2288 B.n578 B.n577 10.6151
R2289 B.n579 B.n578 10.6151
R2290 B.n579 B.n132 10.6151
R2291 B.n583 B.n132 10.6151
R2292 B.n584 B.n583 10.6151
R2293 B.n585 B.n584 10.6151
R2294 B.n585 B.n130 10.6151
R2295 B.n589 B.n130 10.6151
R2296 B.n590 B.n589 10.6151
R2297 B.n591 B.n590 10.6151
R2298 B.n591 B.n128 10.6151
R2299 B.n595 B.n128 10.6151
R2300 B.n596 B.n595 10.6151
R2301 B.n597 B.n596 10.6151
R2302 B.n597 B.n126 10.6151
R2303 B.n601 B.n126 10.6151
R2304 B.n602 B.n601 10.6151
R2305 B.n603 B.n602 10.6151
R2306 B.n603 B.n124 10.6151
R2307 B.n607 B.n124 10.6151
R2308 B.n608 B.n607 10.6151
R2309 B.n609 B.n608 10.6151
R2310 B.n609 B.n122 10.6151
R2311 B.n613 B.n122 10.6151
R2312 B.n614 B.n613 10.6151
R2313 B.n615 B.n614 10.6151
R2314 B.n615 B.n120 10.6151
R2315 B.n619 B.n120 10.6151
R2316 B.n620 B.n619 10.6151
R2317 B.n621 B.n620 10.6151
R2318 B.n621 B.n118 10.6151
R2319 B.n625 B.n118 10.6151
R2320 B.n626 B.n625 10.6151
R2321 B.n627 B.n626 10.6151
R2322 B.n627 B.n116 10.6151
R2323 B.n631 B.n116 10.6151
R2324 B.n632 B.n631 10.6151
R2325 B.n633 B.n632 10.6151
R2326 B.n633 B.n114 10.6151
R2327 B.n637 B.n114 10.6151
R2328 B.n638 B.n637 10.6151
R2329 B.n639 B.n638 10.6151
R2330 B.n639 B.n112 10.6151
R2331 B.n643 B.n112 10.6151
R2332 B.n644 B.n643 10.6151
R2333 B.n645 B.n644 10.6151
R2334 B.n645 B.n110 10.6151
R2335 B.n649 B.n110 10.6151
R2336 B.n650 B.n649 10.6151
R2337 B.n651 B.n650 10.6151
R2338 B.n651 B.n108 10.6151
R2339 B.n655 B.n108 10.6151
R2340 B.n656 B.n655 10.6151
R2341 B.n657 B.n656 10.6151
R2342 B.n657 B.n106 10.6151
R2343 B.n661 B.n106 10.6151
R2344 B.n662 B.n661 10.6151
R2345 B.n663 B.n662 10.6151
R2346 B.n663 B.n104 10.6151
R2347 B.n667 B.n104 10.6151
R2348 B.n668 B.n667 10.6151
R2349 B.n669 B.n668 10.6151
R2350 B.n669 B.n102 10.6151
R2351 B.n673 B.n102 10.6151
R2352 B.n674 B.n673 10.6151
R2353 B.n675 B.n674 10.6151
R2354 B.n675 B.n100 10.6151
R2355 B.n679 B.n100 10.6151
R2356 B.n680 B.n679 10.6151
R2357 B.n681 B.n680 10.6151
R2358 B.n681 B.n98 10.6151
R2359 B.n685 B.n98 10.6151
R2360 B.n686 B.n685 10.6151
R2361 B.n687 B.n686 10.6151
R2362 B.n687 B.n96 10.6151
R2363 B.n691 B.n96 10.6151
R2364 B.n692 B.n691 10.6151
R2365 B.n693 B.n692 10.6151
R2366 B.n693 B.n94 10.6151
R2367 B.n697 B.n94 10.6151
R2368 B.n698 B.n697 10.6151
R2369 B.n699 B.n698 10.6151
R2370 B.n699 B.n92 10.6151
R2371 B.n703 B.n92 10.6151
R2372 B.n704 B.n703 10.6151
R2373 B.n705 B.n704 10.6151
R2374 B.n705 B.n90 10.6151
R2375 B.n709 B.n90 10.6151
R2376 B.n351 B.n212 10.6151
R2377 B.n355 B.n212 10.6151
R2378 B.n356 B.n355 10.6151
R2379 B.n357 B.n356 10.6151
R2380 B.n357 B.n210 10.6151
R2381 B.n361 B.n210 10.6151
R2382 B.n362 B.n361 10.6151
R2383 B.n363 B.n362 10.6151
R2384 B.n363 B.n208 10.6151
R2385 B.n367 B.n208 10.6151
R2386 B.n368 B.n367 10.6151
R2387 B.n369 B.n368 10.6151
R2388 B.n369 B.n206 10.6151
R2389 B.n373 B.n206 10.6151
R2390 B.n374 B.n373 10.6151
R2391 B.n375 B.n374 10.6151
R2392 B.n375 B.n204 10.6151
R2393 B.n379 B.n204 10.6151
R2394 B.n380 B.n379 10.6151
R2395 B.n381 B.n380 10.6151
R2396 B.n381 B.n202 10.6151
R2397 B.n385 B.n202 10.6151
R2398 B.n386 B.n385 10.6151
R2399 B.n387 B.n386 10.6151
R2400 B.n387 B.n200 10.6151
R2401 B.n391 B.n200 10.6151
R2402 B.n392 B.n391 10.6151
R2403 B.n393 B.n392 10.6151
R2404 B.n393 B.n198 10.6151
R2405 B.n397 B.n198 10.6151
R2406 B.n398 B.n397 10.6151
R2407 B.n399 B.n398 10.6151
R2408 B.n399 B.n196 10.6151
R2409 B.n403 B.n196 10.6151
R2410 B.n404 B.n403 10.6151
R2411 B.n405 B.n404 10.6151
R2412 B.n405 B.n194 10.6151
R2413 B.n409 B.n194 10.6151
R2414 B.n410 B.n409 10.6151
R2415 B.n411 B.n410 10.6151
R2416 B.n411 B.n192 10.6151
R2417 B.n415 B.n192 10.6151
R2418 B.n416 B.n415 10.6151
R2419 B.n418 B.n188 10.6151
R2420 B.n422 B.n188 10.6151
R2421 B.n423 B.n422 10.6151
R2422 B.n424 B.n423 10.6151
R2423 B.n424 B.n186 10.6151
R2424 B.n428 B.n186 10.6151
R2425 B.n429 B.n428 10.6151
R2426 B.n430 B.n429 10.6151
R2427 B.n434 B.n433 10.6151
R2428 B.n435 B.n434 10.6151
R2429 B.n435 B.n180 10.6151
R2430 B.n439 B.n180 10.6151
R2431 B.n440 B.n439 10.6151
R2432 B.n441 B.n440 10.6151
R2433 B.n441 B.n178 10.6151
R2434 B.n445 B.n178 10.6151
R2435 B.n446 B.n445 10.6151
R2436 B.n447 B.n446 10.6151
R2437 B.n447 B.n176 10.6151
R2438 B.n451 B.n176 10.6151
R2439 B.n452 B.n451 10.6151
R2440 B.n453 B.n452 10.6151
R2441 B.n453 B.n174 10.6151
R2442 B.n457 B.n174 10.6151
R2443 B.n458 B.n457 10.6151
R2444 B.n459 B.n458 10.6151
R2445 B.n459 B.n172 10.6151
R2446 B.n463 B.n172 10.6151
R2447 B.n464 B.n463 10.6151
R2448 B.n465 B.n464 10.6151
R2449 B.n465 B.n170 10.6151
R2450 B.n469 B.n170 10.6151
R2451 B.n470 B.n469 10.6151
R2452 B.n471 B.n470 10.6151
R2453 B.n471 B.n168 10.6151
R2454 B.n475 B.n168 10.6151
R2455 B.n476 B.n475 10.6151
R2456 B.n477 B.n476 10.6151
R2457 B.n477 B.n166 10.6151
R2458 B.n481 B.n166 10.6151
R2459 B.n482 B.n481 10.6151
R2460 B.n483 B.n482 10.6151
R2461 B.n483 B.n164 10.6151
R2462 B.n487 B.n164 10.6151
R2463 B.n488 B.n487 10.6151
R2464 B.n489 B.n488 10.6151
R2465 B.n489 B.n162 10.6151
R2466 B.n493 B.n162 10.6151
R2467 B.n494 B.n493 10.6151
R2468 B.n495 B.n494 10.6151
R2469 B.n495 B.n160 10.6151
R2470 B.n350 B.n349 10.6151
R2471 B.n349 B.n214 10.6151
R2472 B.n345 B.n214 10.6151
R2473 B.n345 B.n344 10.6151
R2474 B.n344 B.n343 10.6151
R2475 B.n343 B.n216 10.6151
R2476 B.n339 B.n216 10.6151
R2477 B.n339 B.n338 10.6151
R2478 B.n338 B.n337 10.6151
R2479 B.n337 B.n218 10.6151
R2480 B.n333 B.n218 10.6151
R2481 B.n333 B.n332 10.6151
R2482 B.n332 B.n331 10.6151
R2483 B.n331 B.n220 10.6151
R2484 B.n327 B.n220 10.6151
R2485 B.n327 B.n326 10.6151
R2486 B.n326 B.n325 10.6151
R2487 B.n325 B.n222 10.6151
R2488 B.n321 B.n222 10.6151
R2489 B.n321 B.n320 10.6151
R2490 B.n320 B.n319 10.6151
R2491 B.n319 B.n224 10.6151
R2492 B.n315 B.n224 10.6151
R2493 B.n315 B.n314 10.6151
R2494 B.n314 B.n313 10.6151
R2495 B.n313 B.n226 10.6151
R2496 B.n309 B.n226 10.6151
R2497 B.n309 B.n308 10.6151
R2498 B.n308 B.n307 10.6151
R2499 B.n307 B.n228 10.6151
R2500 B.n303 B.n228 10.6151
R2501 B.n303 B.n302 10.6151
R2502 B.n302 B.n301 10.6151
R2503 B.n301 B.n230 10.6151
R2504 B.n297 B.n230 10.6151
R2505 B.n297 B.n296 10.6151
R2506 B.n296 B.n295 10.6151
R2507 B.n295 B.n232 10.6151
R2508 B.n291 B.n232 10.6151
R2509 B.n291 B.n290 10.6151
R2510 B.n290 B.n289 10.6151
R2511 B.n289 B.n234 10.6151
R2512 B.n285 B.n234 10.6151
R2513 B.n285 B.n284 10.6151
R2514 B.n284 B.n283 10.6151
R2515 B.n283 B.n236 10.6151
R2516 B.n279 B.n236 10.6151
R2517 B.n279 B.n278 10.6151
R2518 B.n278 B.n277 10.6151
R2519 B.n277 B.n238 10.6151
R2520 B.n273 B.n238 10.6151
R2521 B.n273 B.n272 10.6151
R2522 B.n272 B.n271 10.6151
R2523 B.n271 B.n240 10.6151
R2524 B.n267 B.n240 10.6151
R2525 B.n267 B.n266 10.6151
R2526 B.n266 B.n265 10.6151
R2527 B.n265 B.n242 10.6151
R2528 B.n261 B.n242 10.6151
R2529 B.n261 B.n260 10.6151
R2530 B.n260 B.n259 10.6151
R2531 B.n259 B.n244 10.6151
R2532 B.n255 B.n244 10.6151
R2533 B.n255 B.n254 10.6151
R2534 B.n254 B.n253 10.6151
R2535 B.n253 B.n246 10.6151
R2536 B.n249 B.n246 10.6151
R2537 B.n249 B.n248 10.6151
R2538 B.n248 B.n0 10.6151
R2539 B.n959 B.n1 10.6151
R2540 B.n959 B.n958 10.6151
R2541 B.n958 B.n957 10.6151
R2542 B.n957 B.n4 10.6151
R2543 B.n953 B.n4 10.6151
R2544 B.n953 B.n952 10.6151
R2545 B.n952 B.n951 10.6151
R2546 B.n951 B.n6 10.6151
R2547 B.n947 B.n6 10.6151
R2548 B.n947 B.n946 10.6151
R2549 B.n946 B.n945 10.6151
R2550 B.n945 B.n8 10.6151
R2551 B.n941 B.n8 10.6151
R2552 B.n941 B.n940 10.6151
R2553 B.n940 B.n939 10.6151
R2554 B.n939 B.n10 10.6151
R2555 B.n935 B.n10 10.6151
R2556 B.n935 B.n934 10.6151
R2557 B.n934 B.n933 10.6151
R2558 B.n933 B.n12 10.6151
R2559 B.n929 B.n12 10.6151
R2560 B.n929 B.n928 10.6151
R2561 B.n928 B.n927 10.6151
R2562 B.n927 B.n14 10.6151
R2563 B.n923 B.n14 10.6151
R2564 B.n923 B.n922 10.6151
R2565 B.n922 B.n921 10.6151
R2566 B.n921 B.n16 10.6151
R2567 B.n917 B.n16 10.6151
R2568 B.n917 B.n916 10.6151
R2569 B.n916 B.n915 10.6151
R2570 B.n915 B.n18 10.6151
R2571 B.n911 B.n18 10.6151
R2572 B.n911 B.n910 10.6151
R2573 B.n910 B.n909 10.6151
R2574 B.n909 B.n20 10.6151
R2575 B.n905 B.n20 10.6151
R2576 B.n905 B.n904 10.6151
R2577 B.n904 B.n903 10.6151
R2578 B.n903 B.n22 10.6151
R2579 B.n899 B.n22 10.6151
R2580 B.n899 B.n898 10.6151
R2581 B.n898 B.n897 10.6151
R2582 B.n897 B.n24 10.6151
R2583 B.n893 B.n24 10.6151
R2584 B.n893 B.n892 10.6151
R2585 B.n892 B.n891 10.6151
R2586 B.n891 B.n26 10.6151
R2587 B.n887 B.n26 10.6151
R2588 B.n887 B.n886 10.6151
R2589 B.n886 B.n885 10.6151
R2590 B.n885 B.n28 10.6151
R2591 B.n881 B.n28 10.6151
R2592 B.n881 B.n880 10.6151
R2593 B.n880 B.n879 10.6151
R2594 B.n879 B.n30 10.6151
R2595 B.n875 B.n30 10.6151
R2596 B.n875 B.n874 10.6151
R2597 B.n874 B.n873 10.6151
R2598 B.n873 B.n32 10.6151
R2599 B.n869 B.n32 10.6151
R2600 B.n869 B.n868 10.6151
R2601 B.n868 B.n867 10.6151
R2602 B.n867 B.n34 10.6151
R2603 B.n863 B.n34 10.6151
R2604 B.n863 B.n862 10.6151
R2605 B.n862 B.n861 10.6151
R2606 B.n861 B.n36 10.6151
R2607 B.n857 B.n36 10.6151
R2608 B.n790 B.n789 6.5566
R2609 B.n777 B.n776 6.5566
R2610 B.n418 B.n417 6.5566
R2611 B.n430 B.n184 6.5566
R2612 B.n791 B.n790 4.05904
R2613 B.n776 B.n775 4.05904
R2614 B.n417 B.n416 4.05904
R2615 B.n433 B.n184 4.05904
R2616 B.n963 B.n0 2.81026
R2617 B.n963 B.n1 2.81026
C0 VP VTAIL 10.580299f
C1 B VN 1.53364f
C2 VDD2 VTAIL 8.89836f
C3 VN VTAIL 10.5662f
C4 w_n5170_n3504# VDD1 2.37569f
C5 B VTAIL 5.73437f
C6 VP w_n5170_n3504# 11.5492f
C7 w_n5170_n3504# VDD2 2.54367f
C8 w_n5170_n3504# VN 10.8743f
C9 B w_n5170_n3504# 12.249901f
C10 VP VDD1 10.284901f
C11 VDD1 VDD2 2.43488f
C12 VP VDD2 0.654872f
C13 w_n5170_n3504# VTAIL 4.47091f
C14 VDD1 VN 0.154084f
C15 B VDD1 2.05577f
C16 VP VN 9.334201f
C17 B VP 2.67181f
C18 VDD2 VN 9.78617f
C19 B VDD2 2.19176f
C20 VDD1 VTAIL 8.835429f
C21 VDD2 VSUBS 2.535111f
C22 VDD1 VSUBS 3.40512f
C23 VTAIL VSUBS 1.607949f
C24 VN VSUBS 8.46744f
C25 VP VSUBS 4.908706f
C26 B VSUBS 6.476863f
C27 w_n5170_n3504# VSUBS 0.222786p
C28 B.n0 VSUBS 0.005303f
C29 B.n1 VSUBS 0.005303f
C30 B.n2 VSUBS 0.008386f
C31 B.n3 VSUBS 0.008386f
C32 B.n4 VSUBS 0.008386f
C33 B.n5 VSUBS 0.008386f
C34 B.n6 VSUBS 0.008386f
C35 B.n7 VSUBS 0.008386f
C36 B.n8 VSUBS 0.008386f
C37 B.n9 VSUBS 0.008386f
C38 B.n10 VSUBS 0.008386f
C39 B.n11 VSUBS 0.008386f
C40 B.n12 VSUBS 0.008386f
C41 B.n13 VSUBS 0.008386f
C42 B.n14 VSUBS 0.008386f
C43 B.n15 VSUBS 0.008386f
C44 B.n16 VSUBS 0.008386f
C45 B.n17 VSUBS 0.008386f
C46 B.n18 VSUBS 0.008386f
C47 B.n19 VSUBS 0.008386f
C48 B.n20 VSUBS 0.008386f
C49 B.n21 VSUBS 0.008386f
C50 B.n22 VSUBS 0.008386f
C51 B.n23 VSUBS 0.008386f
C52 B.n24 VSUBS 0.008386f
C53 B.n25 VSUBS 0.008386f
C54 B.n26 VSUBS 0.008386f
C55 B.n27 VSUBS 0.008386f
C56 B.n28 VSUBS 0.008386f
C57 B.n29 VSUBS 0.008386f
C58 B.n30 VSUBS 0.008386f
C59 B.n31 VSUBS 0.008386f
C60 B.n32 VSUBS 0.008386f
C61 B.n33 VSUBS 0.008386f
C62 B.n34 VSUBS 0.008386f
C63 B.n35 VSUBS 0.008386f
C64 B.n36 VSUBS 0.008386f
C65 B.n37 VSUBS 0.019108f
C66 B.n38 VSUBS 0.008386f
C67 B.n39 VSUBS 0.008386f
C68 B.n40 VSUBS 0.008386f
C69 B.n41 VSUBS 0.008386f
C70 B.n42 VSUBS 0.008386f
C71 B.n43 VSUBS 0.008386f
C72 B.n44 VSUBS 0.008386f
C73 B.n45 VSUBS 0.008386f
C74 B.n46 VSUBS 0.008386f
C75 B.n47 VSUBS 0.008386f
C76 B.n48 VSUBS 0.008386f
C77 B.n49 VSUBS 0.008386f
C78 B.n50 VSUBS 0.008386f
C79 B.n51 VSUBS 0.008386f
C80 B.n52 VSUBS 0.008386f
C81 B.n53 VSUBS 0.008386f
C82 B.n54 VSUBS 0.008386f
C83 B.n55 VSUBS 0.008386f
C84 B.n56 VSUBS 0.008386f
C85 B.n57 VSUBS 0.008386f
C86 B.n58 VSUBS 0.008386f
C87 B.n59 VSUBS 0.008386f
C88 B.t8 VSUBS 0.270937f
C89 B.t7 VSUBS 0.324298f
C90 B.t6 VSUBS 2.73679f
C91 B.n60 VSUBS 0.517699f
C92 B.n61 VSUBS 0.319358f
C93 B.n62 VSUBS 0.008386f
C94 B.n63 VSUBS 0.008386f
C95 B.n64 VSUBS 0.008386f
C96 B.n65 VSUBS 0.008386f
C97 B.t5 VSUBS 0.27094f
C98 B.t4 VSUBS 0.324301f
C99 B.t3 VSUBS 2.73679f
C100 B.n66 VSUBS 0.517695f
C101 B.n67 VSUBS 0.319354f
C102 B.n68 VSUBS 0.008386f
C103 B.n69 VSUBS 0.008386f
C104 B.n70 VSUBS 0.008386f
C105 B.n71 VSUBS 0.008386f
C106 B.n72 VSUBS 0.008386f
C107 B.n73 VSUBS 0.008386f
C108 B.n74 VSUBS 0.008386f
C109 B.n75 VSUBS 0.008386f
C110 B.n76 VSUBS 0.008386f
C111 B.n77 VSUBS 0.008386f
C112 B.n78 VSUBS 0.008386f
C113 B.n79 VSUBS 0.008386f
C114 B.n80 VSUBS 0.008386f
C115 B.n81 VSUBS 0.008386f
C116 B.n82 VSUBS 0.008386f
C117 B.n83 VSUBS 0.008386f
C118 B.n84 VSUBS 0.008386f
C119 B.n85 VSUBS 0.008386f
C120 B.n86 VSUBS 0.008386f
C121 B.n87 VSUBS 0.008386f
C122 B.n88 VSUBS 0.008386f
C123 B.n89 VSUBS 0.019108f
C124 B.n90 VSUBS 0.008386f
C125 B.n91 VSUBS 0.008386f
C126 B.n92 VSUBS 0.008386f
C127 B.n93 VSUBS 0.008386f
C128 B.n94 VSUBS 0.008386f
C129 B.n95 VSUBS 0.008386f
C130 B.n96 VSUBS 0.008386f
C131 B.n97 VSUBS 0.008386f
C132 B.n98 VSUBS 0.008386f
C133 B.n99 VSUBS 0.008386f
C134 B.n100 VSUBS 0.008386f
C135 B.n101 VSUBS 0.008386f
C136 B.n102 VSUBS 0.008386f
C137 B.n103 VSUBS 0.008386f
C138 B.n104 VSUBS 0.008386f
C139 B.n105 VSUBS 0.008386f
C140 B.n106 VSUBS 0.008386f
C141 B.n107 VSUBS 0.008386f
C142 B.n108 VSUBS 0.008386f
C143 B.n109 VSUBS 0.008386f
C144 B.n110 VSUBS 0.008386f
C145 B.n111 VSUBS 0.008386f
C146 B.n112 VSUBS 0.008386f
C147 B.n113 VSUBS 0.008386f
C148 B.n114 VSUBS 0.008386f
C149 B.n115 VSUBS 0.008386f
C150 B.n116 VSUBS 0.008386f
C151 B.n117 VSUBS 0.008386f
C152 B.n118 VSUBS 0.008386f
C153 B.n119 VSUBS 0.008386f
C154 B.n120 VSUBS 0.008386f
C155 B.n121 VSUBS 0.008386f
C156 B.n122 VSUBS 0.008386f
C157 B.n123 VSUBS 0.008386f
C158 B.n124 VSUBS 0.008386f
C159 B.n125 VSUBS 0.008386f
C160 B.n126 VSUBS 0.008386f
C161 B.n127 VSUBS 0.008386f
C162 B.n128 VSUBS 0.008386f
C163 B.n129 VSUBS 0.008386f
C164 B.n130 VSUBS 0.008386f
C165 B.n131 VSUBS 0.008386f
C166 B.n132 VSUBS 0.008386f
C167 B.n133 VSUBS 0.008386f
C168 B.n134 VSUBS 0.008386f
C169 B.n135 VSUBS 0.008386f
C170 B.n136 VSUBS 0.008386f
C171 B.n137 VSUBS 0.008386f
C172 B.n138 VSUBS 0.008386f
C173 B.n139 VSUBS 0.008386f
C174 B.n140 VSUBS 0.008386f
C175 B.n141 VSUBS 0.008386f
C176 B.n142 VSUBS 0.008386f
C177 B.n143 VSUBS 0.008386f
C178 B.n144 VSUBS 0.008386f
C179 B.n145 VSUBS 0.008386f
C180 B.n146 VSUBS 0.008386f
C181 B.n147 VSUBS 0.008386f
C182 B.n148 VSUBS 0.008386f
C183 B.n149 VSUBS 0.008386f
C184 B.n150 VSUBS 0.008386f
C185 B.n151 VSUBS 0.008386f
C186 B.n152 VSUBS 0.008386f
C187 B.n153 VSUBS 0.008386f
C188 B.n154 VSUBS 0.008386f
C189 B.n155 VSUBS 0.008386f
C190 B.n156 VSUBS 0.008386f
C191 B.n157 VSUBS 0.008386f
C192 B.n158 VSUBS 0.008386f
C193 B.n159 VSUBS 0.008386f
C194 B.n160 VSUBS 0.019108f
C195 B.n161 VSUBS 0.008386f
C196 B.n162 VSUBS 0.008386f
C197 B.n163 VSUBS 0.008386f
C198 B.n164 VSUBS 0.008386f
C199 B.n165 VSUBS 0.008386f
C200 B.n166 VSUBS 0.008386f
C201 B.n167 VSUBS 0.008386f
C202 B.n168 VSUBS 0.008386f
C203 B.n169 VSUBS 0.008386f
C204 B.n170 VSUBS 0.008386f
C205 B.n171 VSUBS 0.008386f
C206 B.n172 VSUBS 0.008386f
C207 B.n173 VSUBS 0.008386f
C208 B.n174 VSUBS 0.008386f
C209 B.n175 VSUBS 0.008386f
C210 B.n176 VSUBS 0.008386f
C211 B.n177 VSUBS 0.008386f
C212 B.n178 VSUBS 0.008386f
C213 B.n179 VSUBS 0.008386f
C214 B.n180 VSUBS 0.008386f
C215 B.n181 VSUBS 0.008386f
C216 B.t1 VSUBS 0.27094f
C217 B.t2 VSUBS 0.324301f
C218 B.t0 VSUBS 2.73679f
C219 B.n182 VSUBS 0.517695f
C220 B.n183 VSUBS 0.319354f
C221 B.n184 VSUBS 0.019431f
C222 B.n185 VSUBS 0.008386f
C223 B.n186 VSUBS 0.008386f
C224 B.n187 VSUBS 0.008386f
C225 B.n188 VSUBS 0.008386f
C226 B.n189 VSUBS 0.008386f
C227 B.t10 VSUBS 0.270937f
C228 B.t11 VSUBS 0.324298f
C229 B.t9 VSUBS 2.73679f
C230 B.n190 VSUBS 0.517699f
C231 B.n191 VSUBS 0.319358f
C232 B.n192 VSUBS 0.008386f
C233 B.n193 VSUBS 0.008386f
C234 B.n194 VSUBS 0.008386f
C235 B.n195 VSUBS 0.008386f
C236 B.n196 VSUBS 0.008386f
C237 B.n197 VSUBS 0.008386f
C238 B.n198 VSUBS 0.008386f
C239 B.n199 VSUBS 0.008386f
C240 B.n200 VSUBS 0.008386f
C241 B.n201 VSUBS 0.008386f
C242 B.n202 VSUBS 0.008386f
C243 B.n203 VSUBS 0.008386f
C244 B.n204 VSUBS 0.008386f
C245 B.n205 VSUBS 0.008386f
C246 B.n206 VSUBS 0.008386f
C247 B.n207 VSUBS 0.008386f
C248 B.n208 VSUBS 0.008386f
C249 B.n209 VSUBS 0.008386f
C250 B.n210 VSUBS 0.008386f
C251 B.n211 VSUBS 0.008386f
C252 B.n212 VSUBS 0.008386f
C253 B.n213 VSUBS 0.018138f
C254 B.n214 VSUBS 0.008386f
C255 B.n215 VSUBS 0.008386f
C256 B.n216 VSUBS 0.008386f
C257 B.n217 VSUBS 0.008386f
C258 B.n218 VSUBS 0.008386f
C259 B.n219 VSUBS 0.008386f
C260 B.n220 VSUBS 0.008386f
C261 B.n221 VSUBS 0.008386f
C262 B.n222 VSUBS 0.008386f
C263 B.n223 VSUBS 0.008386f
C264 B.n224 VSUBS 0.008386f
C265 B.n225 VSUBS 0.008386f
C266 B.n226 VSUBS 0.008386f
C267 B.n227 VSUBS 0.008386f
C268 B.n228 VSUBS 0.008386f
C269 B.n229 VSUBS 0.008386f
C270 B.n230 VSUBS 0.008386f
C271 B.n231 VSUBS 0.008386f
C272 B.n232 VSUBS 0.008386f
C273 B.n233 VSUBS 0.008386f
C274 B.n234 VSUBS 0.008386f
C275 B.n235 VSUBS 0.008386f
C276 B.n236 VSUBS 0.008386f
C277 B.n237 VSUBS 0.008386f
C278 B.n238 VSUBS 0.008386f
C279 B.n239 VSUBS 0.008386f
C280 B.n240 VSUBS 0.008386f
C281 B.n241 VSUBS 0.008386f
C282 B.n242 VSUBS 0.008386f
C283 B.n243 VSUBS 0.008386f
C284 B.n244 VSUBS 0.008386f
C285 B.n245 VSUBS 0.008386f
C286 B.n246 VSUBS 0.008386f
C287 B.n247 VSUBS 0.008386f
C288 B.n248 VSUBS 0.008386f
C289 B.n249 VSUBS 0.008386f
C290 B.n250 VSUBS 0.008386f
C291 B.n251 VSUBS 0.008386f
C292 B.n252 VSUBS 0.008386f
C293 B.n253 VSUBS 0.008386f
C294 B.n254 VSUBS 0.008386f
C295 B.n255 VSUBS 0.008386f
C296 B.n256 VSUBS 0.008386f
C297 B.n257 VSUBS 0.008386f
C298 B.n258 VSUBS 0.008386f
C299 B.n259 VSUBS 0.008386f
C300 B.n260 VSUBS 0.008386f
C301 B.n261 VSUBS 0.008386f
C302 B.n262 VSUBS 0.008386f
C303 B.n263 VSUBS 0.008386f
C304 B.n264 VSUBS 0.008386f
C305 B.n265 VSUBS 0.008386f
C306 B.n266 VSUBS 0.008386f
C307 B.n267 VSUBS 0.008386f
C308 B.n268 VSUBS 0.008386f
C309 B.n269 VSUBS 0.008386f
C310 B.n270 VSUBS 0.008386f
C311 B.n271 VSUBS 0.008386f
C312 B.n272 VSUBS 0.008386f
C313 B.n273 VSUBS 0.008386f
C314 B.n274 VSUBS 0.008386f
C315 B.n275 VSUBS 0.008386f
C316 B.n276 VSUBS 0.008386f
C317 B.n277 VSUBS 0.008386f
C318 B.n278 VSUBS 0.008386f
C319 B.n279 VSUBS 0.008386f
C320 B.n280 VSUBS 0.008386f
C321 B.n281 VSUBS 0.008386f
C322 B.n282 VSUBS 0.008386f
C323 B.n283 VSUBS 0.008386f
C324 B.n284 VSUBS 0.008386f
C325 B.n285 VSUBS 0.008386f
C326 B.n286 VSUBS 0.008386f
C327 B.n287 VSUBS 0.008386f
C328 B.n288 VSUBS 0.008386f
C329 B.n289 VSUBS 0.008386f
C330 B.n290 VSUBS 0.008386f
C331 B.n291 VSUBS 0.008386f
C332 B.n292 VSUBS 0.008386f
C333 B.n293 VSUBS 0.008386f
C334 B.n294 VSUBS 0.008386f
C335 B.n295 VSUBS 0.008386f
C336 B.n296 VSUBS 0.008386f
C337 B.n297 VSUBS 0.008386f
C338 B.n298 VSUBS 0.008386f
C339 B.n299 VSUBS 0.008386f
C340 B.n300 VSUBS 0.008386f
C341 B.n301 VSUBS 0.008386f
C342 B.n302 VSUBS 0.008386f
C343 B.n303 VSUBS 0.008386f
C344 B.n304 VSUBS 0.008386f
C345 B.n305 VSUBS 0.008386f
C346 B.n306 VSUBS 0.008386f
C347 B.n307 VSUBS 0.008386f
C348 B.n308 VSUBS 0.008386f
C349 B.n309 VSUBS 0.008386f
C350 B.n310 VSUBS 0.008386f
C351 B.n311 VSUBS 0.008386f
C352 B.n312 VSUBS 0.008386f
C353 B.n313 VSUBS 0.008386f
C354 B.n314 VSUBS 0.008386f
C355 B.n315 VSUBS 0.008386f
C356 B.n316 VSUBS 0.008386f
C357 B.n317 VSUBS 0.008386f
C358 B.n318 VSUBS 0.008386f
C359 B.n319 VSUBS 0.008386f
C360 B.n320 VSUBS 0.008386f
C361 B.n321 VSUBS 0.008386f
C362 B.n322 VSUBS 0.008386f
C363 B.n323 VSUBS 0.008386f
C364 B.n324 VSUBS 0.008386f
C365 B.n325 VSUBS 0.008386f
C366 B.n326 VSUBS 0.008386f
C367 B.n327 VSUBS 0.008386f
C368 B.n328 VSUBS 0.008386f
C369 B.n329 VSUBS 0.008386f
C370 B.n330 VSUBS 0.008386f
C371 B.n331 VSUBS 0.008386f
C372 B.n332 VSUBS 0.008386f
C373 B.n333 VSUBS 0.008386f
C374 B.n334 VSUBS 0.008386f
C375 B.n335 VSUBS 0.008386f
C376 B.n336 VSUBS 0.008386f
C377 B.n337 VSUBS 0.008386f
C378 B.n338 VSUBS 0.008386f
C379 B.n339 VSUBS 0.008386f
C380 B.n340 VSUBS 0.008386f
C381 B.n341 VSUBS 0.008386f
C382 B.n342 VSUBS 0.008386f
C383 B.n343 VSUBS 0.008386f
C384 B.n344 VSUBS 0.008386f
C385 B.n345 VSUBS 0.008386f
C386 B.n346 VSUBS 0.008386f
C387 B.n347 VSUBS 0.008386f
C388 B.n348 VSUBS 0.008386f
C389 B.n349 VSUBS 0.008386f
C390 B.n350 VSUBS 0.018138f
C391 B.n351 VSUBS 0.019108f
C392 B.n352 VSUBS 0.019108f
C393 B.n353 VSUBS 0.008386f
C394 B.n354 VSUBS 0.008386f
C395 B.n355 VSUBS 0.008386f
C396 B.n356 VSUBS 0.008386f
C397 B.n357 VSUBS 0.008386f
C398 B.n358 VSUBS 0.008386f
C399 B.n359 VSUBS 0.008386f
C400 B.n360 VSUBS 0.008386f
C401 B.n361 VSUBS 0.008386f
C402 B.n362 VSUBS 0.008386f
C403 B.n363 VSUBS 0.008386f
C404 B.n364 VSUBS 0.008386f
C405 B.n365 VSUBS 0.008386f
C406 B.n366 VSUBS 0.008386f
C407 B.n367 VSUBS 0.008386f
C408 B.n368 VSUBS 0.008386f
C409 B.n369 VSUBS 0.008386f
C410 B.n370 VSUBS 0.008386f
C411 B.n371 VSUBS 0.008386f
C412 B.n372 VSUBS 0.008386f
C413 B.n373 VSUBS 0.008386f
C414 B.n374 VSUBS 0.008386f
C415 B.n375 VSUBS 0.008386f
C416 B.n376 VSUBS 0.008386f
C417 B.n377 VSUBS 0.008386f
C418 B.n378 VSUBS 0.008386f
C419 B.n379 VSUBS 0.008386f
C420 B.n380 VSUBS 0.008386f
C421 B.n381 VSUBS 0.008386f
C422 B.n382 VSUBS 0.008386f
C423 B.n383 VSUBS 0.008386f
C424 B.n384 VSUBS 0.008386f
C425 B.n385 VSUBS 0.008386f
C426 B.n386 VSUBS 0.008386f
C427 B.n387 VSUBS 0.008386f
C428 B.n388 VSUBS 0.008386f
C429 B.n389 VSUBS 0.008386f
C430 B.n390 VSUBS 0.008386f
C431 B.n391 VSUBS 0.008386f
C432 B.n392 VSUBS 0.008386f
C433 B.n393 VSUBS 0.008386f
C434 B.n394 VSUBS 0.008386f
C435 B.n395 VSUBS 0.008386f
C436 B.n396 VSUBS 0.008386f
C437 B.n397 VSUBS 0.008386f
C438 B.n398 VSUBS 0.008386f
C439 B.n399 VSUBS 0.008386f
C440 B.n400 VSUBS 0.008386f
C441 B.n401 VSUBS 0.008386f
C442 B.n402 VSUBS 0.008386f
C443 B.n403 VSUBS 0.008386f
C444 B.n404 VSUBS 0.008386f
C445 B.n405 VSUBS 0.008386f
C446 B.n406 VSUBS 0.008386f
C447 B.n407 VSUBS 0.008386f
C448 B.n408 VSUBS 0.008386f
C449 B.n409 VSUBS 0.008386f
C450 B.n410 VSUBS 0.008386f
C451 B.n411 VSUBS 0.008386f
C452 B.n412 VSUBS 0.008386f
C453 B.n413 VSUBS 0.008386f
C454 B.n414 VSUBS 0.008386f
C455 B.n415 VSUBS 0.008386f
C456 B.n416 VSUBS 0.005797f
C457 B.n417 VSUBS 0.019431f
C458 B.n418 VSUBS 0.006783f
C459 B.n419 VSUBS 0.008386f
C460 B.n420 VSUBS 0.008386f
C461 B.n421 VSUBS 0.008386f
C462 B.n422 VSUBS 0.008386f
C463 B.n423 VSUBS 0.008386f
C464 B.n424 VSUBS 0.008386f
C465 B.n425 VSUBS 0.008386f
C466 B.n426 VSUBS 0.008386f
C467 B.n427 VSUBS 0.008386f
C468 B.n428 VSUBS 0.008386f
C469 B.n429 VSUBS 0.008386f
C470 B.n430 VSUBS 0.006783f
C471 B.n431 VSUBS 0.008386f
C472 B.n432 VSUBS 0.008386f
C473 B.n433 VSUBS 0.005797f
C474 B.n434 VSUBS 0.008386f
C475 B.n435 VSUBS 0.008386f
C476 B.n436 VSUBS 0.008386f
C477 B.n437 VSUBS 0.008386f
C478 B.n438 VSUBS 0.008386f
C479 B.n439 VSUBS 0.008386f
C480 B.n440 VSUBS 0.008386f
C481 B.n441 VSUBS 0.008386f
C482 B.n442 VSUBS 0.008386f
C483 B.n443 VSUBS 0.008386f
C484 B.n444 VSUBS 0.008386f
C485 B.n445 VSUBS 0.008386f
C486 B.n446 VSUBS 0.008386f
C487 B.n447 VSUBS 0.008386f
C488 B.n448 VSUBS 0.008386f
C489 B.n449 VSUBS 0.008386f
C490 B.n450 VSUBS 0.008386f
C491 B.n451 VSUBS 0.008386f
C492 B.n452 VSUBS 0.008386f
C493 B.n453 VSUBS 0.008386f
C494 B.n454 VSUBS 0.008386f
C495 B.n455 VSUBS 0.008386f
C496 B.n456 VSUBS 0.008386f
C497 B.n457 VSUBS 0.008386f
C498 B.n458 VSUBS 0.008386f
C499 B.n459 VSUBS 0.008386f
C500 B.n460 VSUBS 0.008386f
C501 B.n461 VSUBS 0.008386f
C502 B.n462 VSUBS 0.008386f
C503 B.n463 VSUBS 0.008386f
C504 B.n464 VSUBS 0.008386f
C505 B.n465 VSUBS 0.008386f
C506 B.n466 VSUBS 0.008386f
C507 B.n467 VSUBS 0.008386f
C508 B.n468 VSUBS 0.008386f
C509 B.n469 VSUBS 0.008386f
C510 B.n470 VSUBS 0.008386f
C511 B.n471 VSUBS 0.008386f
C512 B.n472 VSUBS 0.008386f
C513 B.n473 VSUBS 0.008386f
C514 B.n474 VSUBS 0.008386f
C515 B.n475 VSUBS 0.008386f
C516 B.n476 VSUBS 0.008386f
C517 B.n477 VSUBS 0.008386f
C518 B.n478 VSUBS 0.008386f
C519 B.n479 VSUBS 0.008386f
C520 B.n480 VSUBS 0.008386f
C521 B.n481 VSUBS 0.008386f
C522 B.n482 VSUBS 0.008386f
C523 B.n483 VSUBS 0.008386f
C524 B.n484 VSUBS 0.008386f
C525 B.n485 VSUBS 0.008386f
C526 B.n486 VSUBS 0.008386f
C527 B.n487 VSUBS 0.008386f
C528 B.n488 VSUBS 0.008386f
C529 B.n489 VSUBS 0.008386f
C530 B.n490 VSUBS 0.008386f
C531 B.n491 VSUBS 0.008386f
C532 B.n492 VSUBS 0.008386f
C533 B.n493 VSUBS 0.008386f
C534 B.n494 VSUBS 0.008386f
C535 B.n495 VSUBS 0.008386f
C536 B.n496 VSUBS 0.008386f
C537 B.n497 VSUBS 0.019108f
C538 B.n498 VSUBS 0.018138f
C539 B.n499 VSUBS 0.018138f
C540 B.n500 VSUBS 0.008386f
C541 B.n501 VSUBS 0.008386f
C542 B.n502 VSUBS 0.008386f
C543 B.n503 VSUBS 0.008386f
C544 B.n504 VSUBS 0.008386f
C545 B.n505 VSUBS 0.008386f
C546 B.n506 VSUBS 0.008386f
C547 B.n507 VSUBS 0.008386f
C548 B.n508 VSUBS 0.008386f
C549 B.n509 VSUBS 0.008386f
C550 B.n510 VSUBS 0.008386f
C551 B.n511 VSUBS 0.008386f
C552 B.n512 VSUBS 0.008386f
C553 B.n513 VSUBS 0.008386f
C554 B.n514 VSUBS 0.008386f
C555 B.n515 VSUBS 0.008386f
C556 B.n516 VSUBS 0.008386f
C557 B.n517 VSUBS 0.008386f
C558 B.n518 VSUBS 0.008386f
C559 B.n519 VSUBS 0.008386f
C560 B.n520 VSUBS 0.008386f
C561 B.n521 VSUBS 0.008386f
C562 B.n522 VSUBS 0.008386f
C563 B.n523 VSUBS 0.008386f
C564 B.n524 VSUBS 0.008386f
C565 B.n525 VSUBS 0.008386f
C566 B.n526 VSUBS 0.008386f
C567 B.n527 VSUBS 0.008386f
C568 B.n528 VSUBS 0.008386f
C569 B.n529 VSUBS 0.008386f
C570 B.n530 VSUBS 0.008386f
C571 B.n531 VSUBS 0.008386f
C572 B.n532 VSUBS 0.008386f
C573 B.n533 VSUBS 0.008386f
C574 B.n534 VSUBS 0.008386f
C575 B.n535 VSUBS 0.008386f
C576 B.n536 VSUBS 0.008386f
C577 B.n537 VSUBS 0.008386f
C578 B.n538 VSUBS 0.008386f
C579 B.n539 VSUBS 0.008386f
C580 B.n540 VSUBS 0.008386f
C581 B.n541 VSUBS 0.008386f
C582 B.n542 VSUBS 0.008386f
C583 B.n543 VSUBS 0.008386f
C584 B.n544 VSUBS 0.008386f
C585 B.n545 VSUBS 0.008386f
C586 B.n546 VSUBS 0.008386f
C587 B.n547 VSUBS 0.008386f
C588 B.n548 VSUBS 0.008386f
C589 B.n549 VSUBS 0.008386f
C590 B.n550 VSUBS 0.008386f
C591 B.n551 VSUBS 0.008386f
C592 B.n552 VSUBS 0.008386f
C593 B.n553 VSUBS 0.008386f
C594 B.n554 VSUBS 0.008386f
C595 B.n555 VSUBS 0.008386f
C596 B.n556 VSUBS 0.008386f
C597 B.n557 VSUBS 0.008386f
C598 B.n558 VSUBS 0.008386f
C599 B.n559 VSUBS 0.008386f
C600 B.n560 VSUBS 0.008386f
C601 B.n561 VSUBS 0.008386f
C602 B.n562 VSUBS 0.008386f
C603 B.n563 VSUBS 0.008386f
C604 B.n564 VSUBS 0.008386f
C605 B.n565 VSUBS 0.008386f
C606 B.n566 VSUBS 0.008386f
C607 B.n567 VSUBS 0.008386f
C608 B.n568 VSUBS 0.008386f
C609 B.n569 VSUBS 0.008386f
C610 B.n570 VSUBS 0.008386f
C611 B.n571 VSUBS 0.008386f
C612 B.n572 VSUBS 0.008386f
C613 B.n573 VSUBS 0.008386f
C614 B.n574 VSUBS 0.008386f
C615 B.n575 VSUBS 0.008386f
C616 B.n576 VSUBS 0.008386f
C617 B.n577 VSUBS 0.008386f
C618 B.n578 VSUBS 0.008386f
C619 B.n579 VSUBS 0.008386f
C620 B.n580 VSUBS 0.008386f
C621 B.n581 VSUBS 0.008386f
C622 B.n582 VSUBS 0.008386f
C623 B.n583 VSUBS 0.008386f
C624 B.n584 VSUBS 0.008386f
C625 B.n585 VSUBS 0.008386f
C626 B.n586 VSUBS 0.008386f
C627 B.n587 VSUBS 0.008386f
C628 B.n588 VSUBS 0.008386f
C629 B.n589 VSUBS 0.008386f
C630 B.n590 VSUBS 0.008386f
C631 B.n591 VSUBS 0.008386f
C632 B.n592 VSUBS 0.008386f
C633 B.n593 VSUBS 0.008386f
C634 B.n594 VSUBS 0.008386f
C635 B.n595 VSUBS 0.008386f
C636 B.n596 VSUBS 0.008386f
C637 B.n597 VSUBS 0.008386f
C638 B.n598 VSUBS 0.008386f
C639 B.n599 VSUBS 0.008386f
C640 B.n600 VSUBS 0.008386f
C641 B.n601 VSUBS 0.008386f
C642 B.n602 VSUBS 0.008386f
C643 B.n603 VSUBS 0.008386f
C644 B.n604 VSUBS 0.008386f
C645 B.n605 VSUBS 0.008386f
C646 B.n606 VSUBS 0.008386f
C647 B.n607 VSUBS 0.008386f
C648 B.n608 VSUBS 0.008386f
C649 B.n609 VSUBS 0.008386f
C650 B.n610 VSUBS 0.008386f
C651 B.n611 VSUBS 0.008386f
C652 B.n612 VSUBS 0.008386f
C653 B.n613 VSUBS 0.008386f
C654 B.n614 VSUBS 0.008386f
C655 B.n615 VSUBS 0.008386f
C656 B.n616 VSUBS 0.008386f
C657 B.n617 VSUBS 0.008386f
C658 B.n618 VSUBS 0.008386f
C659 B.n619 VSUBS 0.008386f
C660 B.n620 VSUBS 0.008386f
C661 B.n621 VSUBS 0.008386f
C662 B.n622 VSUBS 0.008386f
C663 B.n623 VSUBS 0.008386f
C664 B.n624 VSUBS 0.008386f
C665 B.n625 VSUBS 0.008386f
C666 B.n626 VSUBS 0.008386f
C667 B.n627 VSUBS 0.008386f
C668 B.n628 VSUBS 0.008386f
C669 B.n629 VSUBS 0.008386f
C670 B.n630 VSUBS 0.008386f
C671 B.n631 VSUBS 0.008386f
C672 B.n632 VSUBS 0.008386f
C673 B.n633 VSUBS 0.008386f
C674 B.n634 VSUBS 0.008386f
C675 B.n635 VSUBS 0.008386f
C676 B.n636 VSUBS 0.008386f
C677 B.n637 VSUBS 0.008386f
C678 B.n638 VSUBS 0.008386f
C679 B.n639 VSUBS 0.008386f
C680 B.n640 VSUBS 0.008386f
C681 B.n641 VSUBS 0.008386f
C682 B.n642 VSUBS 0.008386f
C683 B.n643 VSUBS 0.008386f
C684 B.n644 VSUBS 0.008386f
C685 B.n645 VSUBS 0.008386f
C686 B.n646 VSUBS 0.008386f
C687 B.n647 VSUBS 0.008386f
C688 B.n648 VSUBS 0.008386f
C689 B.n649 VSUBS 0.008386f
C690 B.n650 VSUBS 0.008386f
C691 B.n651 VSUBS 0.008386f
C692 B.n652 VSUBS 0.008386f
C693 B.n653 VSUBS 0.008386f
C694 B.n654 VSUBS 0.008386f
C695 B.n655 VSUBS 0.008386f
C696 B.n656 VSUBS 0.008386f
C697 B.n657 VSUBS 0.008386f
C698 B.n658 VSUBS 0.008386f
C699 B.n659 VSUBS 0.008386f
C700 B.n660 VSUBS 0.008386f
C701 B.n661 VSUBS 0.008386f
C702 B.n662 VSUBS 0.008386f
C703 B.n663 VSUBS 0.008386f
C704 B.n664 VSUBS 0.008386f
C705 B.n665 VSUBS 0.008386f
C706 B.n666 VSUBS 0.008386f
C707 B.n667 VSUBS 0.008386f
C708 B.n668 VSUBS 0.008386f
C709 B.n669 VSUBS 0.008386f
C710 B.n670 VSUBS 0.008386f
C711 B.n671 VSUBS 0.008386f
C712 B.n672 VSUBS 0.008386f
C713 B.n673 VSUBS 0.008386f
C714 B.n674 VSUBS 0.008386f
C715 B.n675 VSUBS 0.008386f
C716 B.n676 VSUBS 0.008386f
C717 B.n677 VSUBS 0.008386f
C718 B.n678 VSUBS 0.008386f
C719 B.n679 VSUBS 0.008386f
C720 B.n680 VSUBS 0.008386f
C721 B.n681 VSUBS 0.008386f
C722 B.n682 VSUBS 0.008386f
C723 B.n683 VSUBS 0.008386f
C724 B.n684 VSUBS 0.008386f
C725 B.n685 VSUBS 0.008386f
C726 B.n686 VSUBS 0.008386f
C727 B.n687 VSUBS 0.008386f
C728 B.n688 VSUBS 0.008386f
C729 B.n689 VSUBS 0.008386f
C730 B.n690 VSUBS 0.008386f
C731 B.n691 VSUBS 0.008386f
C732 B.n692 VSUBS 0.008386f
C733 B.n693 VSUBS 0.008386f
C734 B.n694 VSUBS 0.008386f
C735 B.n695 VSUBS 0.008386f
C736 B.n696 VSUBS 0.008386f
C737 B.n697 VSUBS 0.008386f
C738 B.n698 VSUBS 0.008386f
C739 B.n699 VSUBS 0.008386f
C740 B.n700 VSUBS 0.008386f
C741 B.n701 VSUBS 0.008386f
C742 B.n702 VSUBS 0.008386f
C743 B.n703 VSUBS 0.008386f
C744 B.n704 VSUBS 0.008386f
C745 B.n705 VSUBS 0.008386f
C746 B.n706 VSUBS 0.008386f
C747 B.n707 VSUBS 0.008386f
C748 B.n708 VSUBS 0.018138f
C749 B.n709 VSUBS 0.019212f
C750 B.n710 VSUBS 0.018033f
C751 B.n711 VSUBS 0.008386f
C752 B.n712 VSUBS 0.008386f
C753 B.n713 VSUBS 0.008386f
C754 B.n714 VSUBS 0.008386f
C755 B.n715 VSUBS 0.008386f
C756 B.n716 VSUBS 0.008386f
C757 B.n717 VSUBS 0.008386f
C758 B.n718 VSUBS 0.008386f
C759 B.n719 VSUBS 0.008386f
C760 B.n720 VSUBS 0.008386f
C761 B.n721 VSUBS 0.008386f
C762 B.n722 VSUBS 0.008386f
C763 B.n723 VSUBS 0.008386f
C764 B.n724 VSUBS 0.008386f
C765 B.n725 VSUBS 0.008386f
C766 B.n726 VSUBS 0.008386f
C767 B.n727 VSUBS 0.008386f
C768 B.n728 VSUBS 0.008386f
C769 B.n729 VSUBS 0.008386f
C770 B.n730 VSUBS 0.008386f
C771 B.n731 VSUBS 0.008386f
C772 B.n732 VSUBS 0.008386f
C773 B.n733 VSUBS 0.008386f
C774 B.n734 VSUBS 0.008386f
C775 B.n735 VSUBS 0.008386f
C776 B.n736 VSUBS 0.008386f
C777 B.n737 VSUBS 0.008386f
C778 B.n738 VSUBS 0.008386f
C779 B.n739 VSUBS 0.008386f
C780 B.n740 VSUBS 0.008386f
C781 B.n741 VSUBS 0.008386f
C782 B.n742 VSUBS 0.008386f
C783 B.n743 VSUBS 0.008386f
C784 B.n744 VSUBS 0.008386f
C785 B.n745 VSUBS 0.008386f
C786 B.n746 VSUBS 0.008386f
C787 B.n747 VSUBS 0.008386f
C788 B.n748 VSUBS 0.008386f
C789 B.n749 VSUBS 0.008386f
C790 B.n750 VSUBS 0.008386f
C791 B.n751 VSUBS 0.008386f
C792 B.n752 VSUBS 0.008386f
C793 B.n753 VSUBS 0.008386f
C794 B.n754 VSUBS 0.008386f
C795 B.n755 VSUBS 0.008386f
C796 B.n756 VSUBS 0.008386f
C797 B.n757 VSUBS 0.008386f
C798 B.n758 VSUBS 0.008386f
C799 B.n759 VSUBS 0.008386f
C800 B.n760 VSUBS 0.008386f
C801 B.n761 VSUBS 0.008386f
C802 B.n762 VSUBS 0.008386f
C803 B.n763 VSUBS 0.008386f
C804 B.n764 VSUBS 0.008386f
C805 B.n765 VSUBS 0.008386f
C806 B.n766 VSUBS 0.008386f
C807 B.n767 VSUBS 0.008386f
C808 B.n768 VSUBS 0.008386f
C809 B.n769 VSUBS 0.008386f
C810 B.n770 VSUBS 0.008386f
C811 B.n771 VSUBS 0.008386f
C812 B.n772 VSUBS 0.008386f
C813 B.n773 VSUBS 0.008386f
C814 B.n774 VSUBS 0.008386f
C815 B.n775 VSUBS 0.005797f
C816 B.n776 VSUBS 0.019431f
C817 B.n777 VSUBS 0.006783f
C818 B.n778 VSUBS 0.008386f
C819 B.n779 VSUBS 0.008386f
C820 B.n780 VSUBS 0.008386f
C821 B.n781 VSUBS 0.008386f
C822 B.n782 VSUBS 0.008386f
C823 B.n783 VSUBS 0.008386f
C824 B.n784 VSUBS 0.008386f
C825 B.n785 VSUBS 0.008386f
C826 B.n786 VSUBS 0.008386f
C827 B.n787 VSUBS 0.008386f
C828 B.n788 VSUBS 0.008386f
C829 B.n789 VSUBS 0.006783f
C830 B.n790 VSUBS 0.019431f
C831 B.n791 VSUBS 0.005797f
C832 B.n792 VSUBS 0.008386f
C833 B.n793 VSUBS 0.008386f
C834 B.n794 VSUBS 0.008386f
C835 B.n795 VSUBS 0.008386f
C836 B.n796 VSUBS 0.008386f
C837 B.n797 VSUBS 0.008386f
C838 B.n798 VSUBS 0.008386f
C839 B.n799 VSUBS 0.008386f
C840 B.n800 VSUBS 0.008386f
C841 B.n801 VSUBS 0.008386f
C842 B.n802 VSUBS 0.008386f
C843 B.n803 VSUBS 0.008386f
C844 B.n804 VSUBS 0.008386f
C845 B.n805 VSUBS 0.008386f
C846 B.n806 VSUBS 0.008386f
C847 B.n807 VSUBS 0.008386f
C848 B.n808 VSUBS 0.008386f
C849 B.n809 VSUBS 0.008386f
C850 B.n810 VSUBS 0.008386f
C851 B.n811 VSUBS 0.008386f
C852 B.n812 VSUBS 0.008386f
C853 B.n813 VSUBS 0.008386f
C854 B.n814 VSUBS 0.008386f
C855 B.n815 VSUBS 0.008386f
C856 B.n816 VSUBS 0.008386f
C857 B.n817 VSUBS 0.008386f
C858 B.n818 VSUBS 0.008386f
C859 B.n819 VSUBS 0.008386f
C860 B.n820 VSUBS 0.008386f
C861 B.n821 VSUBS 0.008386f
C862 B.n822 VSUBS 0.008386f
C863 B.n823 VSUBS 0.008386f
C864 B.n824 VSUBS 0.008386f
C865 B.n825 VSUBS 0.008386f
C866 B.n826 VSUBS 0.008386f
C867 B.n827 VSUBS 0.008386f
C868 B.n828 VSUBS 0.008386f
C869 B.n829 VSUBS 0.008386f
C870 B.n830 VSUBS 0.008386f
C871 B.n831 VSUBS 0.008386f
C872 B.n832 VSUBS 0.008386f
C873 B.n833 VSUBS 0.008386f
C874 B.n834 VSUBS 0.008386f
C875 B.n835 VSUBS 0.008386f
C876 B.n836 VSUBS 0.008386f
C877 B.n837 VSUBS 0.008386f
C878 B.n838 VSUBS 0.008386f
C879 B.n839 VSUBS 0.008386f
C880 B.n840 VSUBS 0.008386f
C881 B.n841 VSUBS 0.008386f
C882 B.n842 VSUBS 0.008386f
C883 B.n843 VSUBS 0.008386f
C884 B.n844 VSUBS 0.008386f
C885 B.n845 VSUBS 0.008386f
C886 B.n846 VSUBS 0.008386f
C887 B.n847 VSUBS 0.008386f
C888 B.n848 VSUBS 0.008386f
C889 B.n849 VSUBS 0.008386f
C890 B.n850 VSUBS 0.008386f
C891 B.n851 VSUBS 0.008386f
C892 B.n852 VSUBS 0.008386f
C893 B.n853 VSUBS 0.008386f
C894 B.n854 VSUBS 0.008386f
C895 B.n855 VSUBS 0.008386f
C896 B.n856 VSUBS 0.019108f
C897 B.n857 VSUBS 0.018138f
C898 B.n858 VSUBS 0.018138f
C899 B.n859 VSUBS 0.008386f
C900 B.n860 VSUBS 0.008386f
C901 B.n861 VSUBS 0.008386f
C902 B.n862 VSUBS 0.008386f
C903 B.n863 VSUBS 0.008386f
C904 B.n864 VSUBS 0.008386f
C905 B.n865 VSUBS 0.008386f
C906 B.n866 VSUBS 0.008386f
C907 B.n867 VSUBS 0.008386f
C908 B.n868 VSUBS 0.008386f
C909 B.n869 VSUBS 0.008386f
C910 B.n870 VSUBS 0.008386f
C911 B.n871 VSUBS 0.008386f
C912 B.n872 VSUBS 0.008386f
C913 B.n873 VSUBS 0.008386f
C914 B.n874 VSUBS 0.008386f
C915 B.n875 VSUBS 0.008386f
C916 B.n876 VSUBS 0.008386f
C917 B.n877 VSUBS 0.008386f
C918 B.n878 VSUBS 0.008386f
C919 B.n879 VSUBS 0.008386f
C920 B.n880 VSUBS 0.008386f
C921 B.n881 VSUBS 0.008386f
C922 B.n882 VSUBS 0.008386f
C923 B.n883 VSUBS 0.008386f
C924 B.n884 VSUBS 0.008386f
C925 B.n885 VSUBS 0.008386f
C926 B.n886 VSUBS 0.008386f
C927 B.n887 VSUBS 0.008386f
C928 B.n888 VSUBS 0.008386f
C929 B.n889 VSUBS 0.008386f
C930 B.n890 VSUBS 0.008386f
C931 B.n891 VSUBS 0.008386f
C932 B.n892 VSUBS 0.008386f
C933 B.n893 VSUBS 0.008386f
C934 B.n894 VSUBS 0.008386f
C935 B.n895 VSUBS 0.008386f
C936 B.n896 VSUBS 0.008386f
C937 B.n897 VSUBS 0.008386f
C938 B.n898 VSUBS 0.008386f
C939 B.n899 VSUBS 0.008386f
C940 B.n900 VSUBS 0.008386f
C941 B.n901 VSUBS 0.008386f
C942 B.n902 VSUBS 0.008386f
C943 B.n903 VSUBS 0.008386f
C944 B.n904 VSUBS 0.008386f
C945 B.n905 VSUBS 0.008386f
C946 B.n906 VSUBS 0.008386f
C947 B.n907 VSUBS 0.008386f
C948 B.n908 VSUBS 0.008386f
C949 B.n909 VSUBS 0.008386f
C950 B.n910 VSUBS 0.008386f
C951 B.n911 VSUBS 0.008386f
C952 B.n912 VSUBS 0.008386f
C953 B.n913 VSUBS 0.008386f
C954 B.n914 VSUBS 0.008386f
C955 B.n915 VSUBS 0.008386f
C956 B.n916 VSUBS 0.008386f
C957 B.n917 VSUBS 0.008386f
C958 B.n918 VSUBS 0.008386f
C959 B.n919 VSUBS 0.008386f
C960 B.n920 VSUBS 0.008386f
C961 B.n921 VSUBS 0.008386f
C962 B.n922 VSUBS 0.008386f
C963 B.n923 VSUBS 0.008386f
C964 B.n924 VSUBS 0.008386f
C965 B.n925 VSUBS 0.008386f
C966 B.n926 VSUBS 0.008386f
C967 B.n927 VSUBS 0.008386f
C968 B.n928 VSUBS 0.008386f
C969 B.n929 VSUBS 0.008386f
C970 B.n930 VSUBS 0.008386f
C971 B.n931 VSUBS 0.008386f
C972 B.n932 VSUBS 0.008386f
C973 B.n933 VSUBS 0.008386f
C974 B.n934 VSUBS 0.008386f
C975 B.n935 VSUBS 0.008386f
C976 B.n936 VSUBS 0.008386f
C977 B.n937 VSUBS 0.008386f
C978 B.n938 VSUBS 0.008386f
C979 B.n939 VSUBS 0.008386f
C980 B.n940 VSUBS 0.008386f
C981 B.n941 VSUBS 0.008386f
C982 B.n942 VSUBS 0.008386f
C983 B.n943 VSUBS 0.008386f
C984 B.n944 VSUBS 0.008386f
C985 B.n945 VSUBS 0.008386f
C986 B.n946 VSUBS 0.008386f
C987 B.n947 VSUBS 0.008386f
C988 B.n948 VSUBS 0.008386f
C989 B.n949 VSUBS 0.008386f
C990 B.n950 VSUBS 0.008386f
C991 B.n951 VSUBS 0.008386f
C992 B.n952 VSUBS 0.008386f
C993 B.n953 VSUBS 0.008386f
C994 B.n954 VSUBS 0.008386f
C995 B.n955 VSUBS 0.008386f
C996 B.n956 VSUBS 0.008386f
C997 B.n957 VSUBS 0.008386f
C998 B.n958 VSUBS 0.008386f
C999 B.n959 VSUBS 0.008386f
C1000 B.n960 VSUBS 0.008386f
C1001 B.n961 VSUBS 0.008386f
C1002 B.n962 VSUBS 0.008386f
C1003 B.n963 VSUBS 0.01899f
C1004 VDD1.t5 VSUBS 0.333408f
C1005 VDD1.t0 VSUBS 0.333408f
C1006 VDD1.n0 VSUBS 2.68522f
C1007 VDD1.t4 VSUBS 0.333408f
C1008 VDD1.t6 VSUBS 0.333408f
C1009 VDD1.n1 VSUBS 2.68325f
C1010 VDD1.t1 VSUBS 0.333408f
C1011 VDD1.t3 VSUBS 0.333408f
C1012 VDD1.n2 VSUBS 2.68325f
C1013 VDD1.n3 VSUBS 6.11208f
C1014 VDD1.t7 VSUBS 0.333408f
C1015 VDD1.t2 VSUBS 0.333408f
C1016 VDD1.n4 VSUBS 2.65655f
C1017 VDD1.n5 VSUBS 4.95038f
C1018 VP.t4 VSUBS 3.39728f
C1019 VP.n0 VSUBS 1.28184f
C1020 VP.n1 VSUBS 0.025371f
C1021 VP.n2 VSUBS 0.050958f
C1022 VP.n3 VSUBS 0.025371f
C1023 VP.n4 VSUBS 0.047047f
C1024 VP.n5 VSUBS 0.025371f
C1025 VP.t6 VSUBS 3.39728f
C1026 VP.n6 VSUBS 0.047047f
C1027 VP.n7 VSUBS 0.025371f
C1028 VP.n8 VSUBS 0.047047f
C1029 VP.n9 VSUBS 0.025371f
C1030 VP.t1 VSUBS 3.39728f
C1031 VP.n10 VSUBS 0.047047f
C1032 VP.n11 VSUBS 0.025371f
C1033 VP.n12 VSUBS 0.047047f
C1034 VP.n13 VSUBS 0.040941f
C1035 VP.t3 VSUBS 3.39728f
C1036 VP.t5 VSUBS 3.39728f
C1037 VP.n14 VSUBS 1.28184f
C1038 VP.n15 VSUBS 0.025371f
C1039 VP.n16 VSUBS 0.050958f
C1040 VP.n17 VSUBS 0.025371f
C1041 VP.n18 VSUBS 0.047047f
C1042 VP.n19 VSUBS 0.025371f
C1043 VP.t0 VSUBS 3.39728f
C1044 VP.n20 VSUBS 0.047047f
C1045 VP.n21 VSUBS 0.025371f
C1046 VP.n22 VSUBS 0.047047f
C1047 VP.t2 VSUBS 3.80504f
C1048 VP.n23 VSUBS 1.21804f
C1049 VP.t7 VSUBS 3.39728f
C1050 VP.n24 VSUBS 1.28213f
C1051 VP.n25 VSUBS 0.040079f
C1052 VP.n26 VSUBS 0.328267f
C1053 VP.n27 VSUBS 0.025371f
C1054 VP.n28 VSUBS 0.025371f
C1055 VP.n29 VSUBS 0.047047f
C1056 VP.n30 VSUBS 0.03688f
C1057 VP.n31 VSUBS 0.03688f
C1058 VP.n32 VSUBS 0.025371f
C1059 VP.n33 VSUBS 0.025371f
C1060 VP.n34 VSUBS 0.025371f
C1061 VP.n35 VSUBS 0.047047f
C1062 VP.n36 VSUBS 0.040079f
C1063 VP.n37 VSUBS 1.18622f
C1064 VP.n38 VSUBS 0.030789f
C1065 VP.n39 VSUBS 0.025371f
C1066 VP.n40 VSUBS 0.025371f
C1067 VP.n41 VSUBS 0.025371f
C1068 VP.n42 VSUBS 0.047047f
C1069 VP.n43 VSUBS 0.048538f
C1070 VP.n44 VSUBS 0.021311f
C1071 VP.n45 VSUBS 0.025371f
C1072 VP.n46 VSUBS 0.025371f
C1073 VP.n47 VSUBS 0.025371f
C1074 VP.n48 VSUBS 0.047047f
C1075 VP.n49 VSUBS 0.047047f
C1076 VP.n50 VSUBS 0.026144f
C1077 VP.n51 VSUBS 0.040941f
C1078 VP.n52 VSUBS 1.76913f
C1079 VP.n53 VSUBS 1.78506f
C1080 VP.n54 VSUBS 1.28184f
C1081 VP.n55 VSUBS 0.026144f
C1082 VP.n56 VSUBS 0.047047f
C1083 VP.n57 VSUBS 0.025371f
C1084 VP.n58 VSUBS 0.025371f
C1085 VP.n59 VSUBS 0.025371f
C1086 VP.n60 VSUBS 0.050958f
C1087 VP.n61 VSUBS 0.021311f
C1088 VP.n62 VSUBS 0.048538f
C1089 VP.n63 VSUBS 0.025371f
C1090 VP.n64 VSUBS 0.025371f
C1091 VP.n65 VSUBS 0.025371f
C1092 VP.n66 VSUBS 0.047047f
C1093 VP.n67 VSUBS 0.030789f
C1094 VP.n68 VSUBS 1.18622f
C1095 VP.n69 VSUBS 0.040079f
C1096 VP.n70 VSUBS 0.025371f
C1097 VP.n71 VSUBS 0.025371f
C1098 VP.n72 VSUBS 0.025371f
C1099 VP.n73 VSUBS 0.047047f
C1100 VP.n74 VSUBS 0.03688f
C1101 VP.n75 VSUBS 0.03688f
C1102 VP.n76 VSUBS 0.025371f
C1103 VP.n77 VSUBS 0.025371f
C1104 VP.n78 VSUBS 0.025371f
C1105 VP.n79 VSUBS 0.047047f
C1106 VP.n80 VSUBS 0.040079f
C1107 VP.n81 VSUBS 1.18622f
C1108 VP.n82 VSUBS 0.030789f
C1109 VP.n83 VSUBS 0.025371f
C1110 VP.n84 VSUBS 0.025371f
C1111 VP.n85 VSUBS 0.025371f
C1112 VP.n86 VSUBS 0.047047f
C1113 VP.n87 VSUBS 0.048538f
C1114 VP.n88 VSUBS 0.021311f
C1115 VP.n89 VSUBS 0.025371f
C1116 VP.n90 VSUBS 0.025371f
C1117 VP.n91 VSUBS 0.025371f
C1118 VP.n92 VSUBS 0.047047f
C1119 VP.n93 VSUBS 0.047047f
C1120 VP.n94 VSUBS 0.026144f
C1121 VP.n95 VSUBS 0.040941f
C1122 VP.n96 VSUBS 0.079148f
C1123 VTAIL.t9 VSUBS 0.260072f
C1124 VTAIL.t14 VSUBS 0.260072f
C1125 VTAIL.n0 VSUBS 1.94307f
C1126 VTAIL.n1 VSUBS 0.869995f
C1127 VTAIL.n2 VSUBS 0.014633f
C1128 VTAIL.n3 VSUBS 0.032966f
C1129 VTAIL.n4 VSUBS 0.014767f
C1130 VTAIL.n5 VSUBS 0.025955f
C1131 VTAIL.n6 VSUBS 0.013947f
C1132 VTAIL.n7 VSUBS 0.032966f
C1133 VTAIL.n8 VSUBS 0.014767f
C1134 VTAIL.n9 VSUBS 0.025955f
C1135 VTAIL.n10 VSUBS 0.013947f
C1136 VTAIL.n11 VSUBS 0.032966f
C1137 VTAIL.n12 VSUBS 0.014767f
C1138 VTAIL.n13 VSUBS 0.025955f
C1139 VTAIL.n14 VSUBS 0.013947f
C1140 VTAIL.n15 VSUBS 0.032966f
C1141 VTAIL.n16 VSUBS 0.014767f
C1142 VTAIL.n17 VSUBS 0.025955f
C1143 VTAIL.n18 VSUBS 0.013947f
C1144 VTAIL.n19 VSUBS 0.032966f
C1145 VTAIL.n20 VSUBS 0.014767f
C1146 VTAIL.n21 VSUBS 0.025955f
C1147 VTAIL.n22 VSUBS 0.013947f
C1148 VTAIL.n23 VSUBS 0.024724f
C1149 VTAIL.n24 VSUBS 0.020971f
C1150 VTAIL.t10 VSUBS 0.070426f
C1151 VTAIL.n25 VSUBS 0.165202f
C1152 VTAIL.n26 VSUBS 1.38391f
C1153 VTAIL.n27 VSUBS 0.013947f
C1154 VTAIL.n28 VSUBS 0.014767f
C1155 VTAIL.n29 VSUBS 0.032966f
C1156 VTAIL.n30 VSUBS 0.032966f
C1157 VTAIL.n31 VSUBS 0.014767f
C1158 VTAIL.n32 VSUBS 0.013947f
C1159 VTAIL.n33 VSUBS 0.025955f
C1160 VTAIL.n34 VSUBS 0.025955f
C1161 VTAIL.n35 VSUBS 0.013947f
C1162 VTAIL.n36 VSUBS 0.014767f
C1163 VTAIL.n37 VSUBS 0.032966f
C1164 VTAIL.n38 VSUBS 0.032966f
C1165 VTAIL.n39 VSUBS 0.014767f
C1166 VTAIL.n40 VSUBS 0.013947f
C1167 VTAIL.n41 VSUBS 0.025955f
C1168 VTAIL.n42 VSUBS 0.025955f
C1169 VTAIL.n43 VSUBS 0.013947f
C1170 VTAIL.n44 VSUBS 0.014767f
C1171 VTAIL.n45 VSUBS 0.032966f
C1172 VTAIL.n46 VSUBS 0.032966f
C1173 VTAIL.n47 VSUBS 0.014767f
C1174 VTAIL.n48 VSUBS 0.013947f
C1175 VTAIL.n49 VSUBS 0.025955f
C1176 VTAIL.n50 VSUBS 0.025955f
C1177 VTAIL.n51 VSUBS 0.013947f
C1178 VTAIL.n52 VSUBS 0.014767f
C1179 VTAIL.n53 VSUBS 0.032966f
C1180 VTAIL.n54 VSUBS 0.032966f
C1181 VTAIL.n55 VSUBS 0.014767f
C1182 VTAIL.n56 VSUBS 0.013947f
C1183 VTAIL.n57 VSUBS 0.025955f
C1184 VTAIL.n58 VSUBS 0.025955f
C1185 VTAIL.n59 VSUBS 0.013947f
C1186 VTAIL.n60 VSUBS 0.014767f
C1187 VTAIL.n61 VSUBS 0.032966f
C1188 VTAIL.n62 VSUBS 0.032966f
C1189 VTAIL.n63 VSUBS 0.014767f
C1190 VTAIL.n64 VSUBS 0.013947f
C1191 VTAIL.n65 VSUBS 0.025955f
C1192 VTAIL.n66 VSUBS 0.067085f
C1193 VTAIL.n67 VSUBS 0.013947f
C1194 VTAIL.n68 VSUBS 0.014767f
C1195 VTAIL.n69 VSUBS 0.07494f
C1196 VTAIL.n70 VSUBS 0.049716f
C1197 VTAIL.n71 VSUBS 0.36788f
C1198 VTAIL.n72 VSUBS 0.014633f
C1199 VTAIL.n73 VSUBS 0.032966f
C1200 VTAIL.n74 VSUBS 0.014767f
C1201 VTAIL.n75 VSUBS 0.025955f
C1202 VTAIL.n76 VSUBS 0.013947f
C1203 VTAIL.n77 VSUBS 0.032966f
C1204 VTAIL.n78 VSUBS 0.014767f
C1205 VTAIL.n79 VSUBS 0.025955f
C1206 VTAIL.n80 VSUBS 0.013947f
C1207 VTAIL.n81 VSUBS 0.032966f
C1208 VTAIL.n82 VSUBS 0.014767f
C1209 VTAIL.n83 VSUBS 0.025955f
C1210 VTAIL.n84 VSUBS 0.013947f
C1211 VTAIL.n85 VSUBS 0.032966f
C1212 VTAIL.n86 VSUBS 0.014767f
C1213 VTAIL.n87 VSUBS 0.025955f
C1214 VTAIL.n88 VSUBS 0.013947f
C1215 VTAIL.n89 VSUBS 0.032966f
C1216 VTAIL.n90 VSUBS 0.014767f
C1217 VTAIL.n91 VSUBS 0.025955f
C1218 VTAIL.n92 VSUBS 0.013947f
C1219 VTAIL.n93 VSUBS 0.024724f
C1220 VTAIL.n94 VSUBS 0.020971f
C1221 VTAIL.t4 VSUBS 0.070426f
C1222 VTAIL.n95 VSUBS 0.165202f
C1223 VTAIL.n96 VSUBS 1.38391f
C1224 VTAIL.n97 VSUBS 0.013947f
C1225 VTAIL.n98 VSUBS 0.014767f
C1226 VTAIL.n99 VSUBS 0.032966f
C1227 VTAIL.n100 VSUBS 0.032966f
C1228 VTAIL.n101 VSUBS 0.014767f
C1229 VTAIL.n102 VSUBS 0.013947f
C1230 VTAIL.n103 VSUBS 0.025955f
C1231 VTAIL.n104 VSUBS 0.025955f
C1232 VTAIL.n105 VSUBS 0.013947f
C1233 VTAIL.n106 VSUBS 0.014767f
C1234 VTAIL.n107 VSUBS 0.032966f
C1235 VTAIL.n108 VSUBS 0.032966f
C1236 VTAIL.n109 VSUBS 0.014767f
C1237 VTAIL.n110 VSUBS 0.013947f
C1238 VTAIL.n111 VSUBS 0.025955f
C1239 VTAIL.n112 VSUBS 0.025955f
C1240 VTAIL.n113 VSUBS 0.013947f
C1241 VTAIL.n114 VSUBS 0.014767f
C1242 VTAIL.n115 VSUBS 0.032966f
C1243 VTAIL.n116 VSUBS 0.032966f
C1244 VTAIL.n117 VSUBS 0.014767f
C1245 VTAIL.n118 VSUBS 0.013947f
C1246 VTAIL.n119 VSUBS 0.025955f
C1247 VTAIL.n120 VSUBS 0.025955f
C1248 VTAIL.n121 VSUBS 0.013947f
C1249 VTAIL.n122 VSUBS 0.014767f
C1250 VTAIL.n123 VSUBS 0.032966f
C1251 VTAIL.n124 VSUBS 0.032966f
C1252 VTAIL.n125 VSUBS 0.014767f
C1253 VTAIL.n126 VSUBS 0.013947f
C1254 VTAIL.n127 VSUBS 0.025955f
C1255 VTAIL.n128 VSUBS 0.025955f
C1256 VTAIL.n129 VSUBS 0.013947f
C1257 VTAIL.n130 VSUBS 0.014767f
C1258 VTAIL.n131 VSUBS 0.032966f
C1259 VTAIL.n132 VSUBS 0.032966f
C1260 VTAIL.n133 VSUBS 0.014767f
C1261 VTAIL.n134 VSUBS 0.013947f
C1262 VTAIL.n135 VSUBS 0.025955f
C1263 VTAIL.n136 VSUBS 0.067085f
C1264 VTAIL.n137 VSUBS 0.013947f
C1265 VTAIL.n138 VSUBS 0.014767f
C1266 VTAIL.n139 VSUBS 0.07494f
C1267 VTAIL.n140 VSUBS 0.049716f
C1268 VTAIL.n141 VSUBS 0.36788f
C1269 VTAIL.t1 VSUBS 0.260072f
C1270 VTAIL.t6 VSUBS 0.260072f
C1271 VTAIL.n142 VSUBS 1.94307f
C1272 VTAIL.n143 VSUBS 1.16794f
C1273 VTAIL.n144 VSUBS 0.014633f
C1274 VTAIL.n145 VSUBS 0.032966f
C1275 VTAIL.n146 VSUBS 0.014767f
C1276 VTAIL.n147 VSUBS 0.025955f
C1277 VTAIL.n148 VSUBS 0.013947f
C1278 VTAIL.n149 VSUBS 0.032966f
C1279 VTAIL.n150 VSUBS 0.014767f
C1280 VTAIL.n151 VSUBS 0.025955f
C1281 VTAIL.n152 VSUBS 0.013947f
C1282 VTAIL.n153 VSUBS 0.032966f
C1283 VTAIL.n154 VSUBS 0.014767f
C1284 VTAIL.n155 VSUBS 0.025955f
C1285 VTAIL.n156 VSUBS 0.013947f
C1286 VTAIL.n157 VSUBS 0.032966f
C1287 VTAIL.n158 VSUBS 0.014767f
C1288 VTAIL.n159 VSUBS 0.025955f
C1289 VTAIL.n160 VSUBS 0.013947f
C1290 VTAIL.n161 VSUBS 0.032966f
C1291 VTAIL.n162 VSUBS 0.014767f
C1292 VTAIL.n163 VSUBS 0.025955f
C1293 VTAIL.n164 VSUBS 0.013947f
C1294 VTAIL.n165 VSUBS 0.024724f
C1295 VTAIL.n166 VSUBS 0.020971f
C1296 VTAIL.t3 VSUBS 0.070426f
C1297 VTAIL.n167 VSUBS 0.165202f
C1298 VTAIL.n168 VSUBS 1.38391f
C1299 VTAIL.n169 VSUBS 0.013947f
C1300 VTAIL.n170 VSUBS 0.014767f
C1301 VTAIL.n171 VSUBS 0.032966f
C1302 VTAIL.n172 VSUBS 0.032966f
C1303 VTAIL.n173 VSUBS 0.014767f
C1304 VTAIL.n174 VSUBS 0.013947f
C1305 VTAIL.n175 VSUBS 0.025955f
C1306 VTAIL.n176 VSUBS 0.025955f
C1307 VTAIL.n177 VSUBS 0.013947f
C1308 VTAIL.n178 VSUBS 0.014767f
C1309 VTAIL.n179 VSUBS 0.032966f
C1310 VTAIL.n180 VSUBS 0.032966f
C1311 VTAIL.n181 VSUBS 0.014767f
C1312 VTAIL.n182 VSUBS 0.013947f
C1313 VTAIL.n183 VSUBS 0.025955f
C1314 VTAIL.n184 VSUBS 0.025955f
C1315 VTAIL.n185 VSUBS 0.013947f
C1316 VTAIL.n186 VSUBS 0.014767f
C1317 VTAIL.n187 VSUBS 0.032966f
C1318 VTAIL.n188 VSUBS 0.032966f
C1319 VTAIL.n189 VSUBS 0.014767f
C1320 VTAIL.n190 VSUBS 0.013947f
C1321 VTAIL.n191 VSUBS 0.025955f
C1322 VTAIL.n192 VSUBS 0.025955f
C1323 VTAIL.n193 VSUBS 0.013947f
C1324 VTAIL.n194 VSUBS 0.014767f
C1325 VTAIL.n195 VSUBS 0.032966f
C1326 VTAIL.n196 VSUBS 0.032966f
C1327 VTAIL.n197 VSUBS 0.014767f
C1328 VTAIL.n198 VSUBS 0.013947f
C1329 VTAIL.n199 VSUBS 0.025955f
C1330 VTAIL.n200 VSUBS 0.025955f
C1331 VTAIL.n201 VSUBS 0.013947f
C1332 VTAIL.n202 VSUBS 0.014767f
C1333 VTAIL.n203 VSUBS 0.032966f
C1334 VTAIL.n204 VSUBS 0.032966f
C1335 VTAIL.n205 VSUBS 0.014767f
C1336 VTAIL.n206 VSUBS 0.013947f
C1337 VTAIL.n207 VSUBS 0.025955f
C1338 VTAIL.n208 VSUBS 0.067085f
C1339 VTAIL.n209 VSUBS 0.013947f
C1340 VTAIL.n210 VSUBS 0.014767f
C1341 VTAIL.n211 VSUBS 0.07494f
C1342 VTAIL.n212 VSUBS 0.049716f
C1343 VTAIL.n213 VSUBS 1.89816f
C1344 VTAIL.n214 VSUBS 0.014633f
C1345 VTAIL.n215 VSUBS 0.032966f
C1346 VTAIL.n216 VSUBS 0.014767f
C1347 VTAIL.n217 VSUBS 0.025955f
C1348 VTAIL.n218 VSUBS 0.013947f
C1349 VTAIL.n219 VSUBS 0.032966f
C1350 VTAIL.n220 VSUBS 0.014767f
C1351 VTAIL.n221 VSUBS 0.025955f
C1352 VTAIL.n222 VSUBS 0.013947f
C1353 VTAIL.n223 VSUBS 0.032966f
C1354 VTAIL.n224 VSUBS 0.014767f
C1355 VTAIL.n225 VSUBS 0.025955f
C1356 VTAIL.n226 VSUBS 0.013947f
C1357 VTAIL.n227 VSUBS 0.032966f
C1358 VTAIL.n228 VSUBS 0.014767f
C1359 VTAIL.n229 VSUBS 0.025955f
C1360 VTAIL.n230 VSUBS 0.013947f
C1361 VTAIL.n231 VSUBS 0.032966f
C1362 VTAIL.n232 VSUBS 0.014767f
C1363 VTAIL.n233 VSUBS 0.025955f
C1364 VTAIL.n234 VSUBS 0.013947f
C1365 VTAIL.n235 VSUBS 0.024724f
C1366 VTAIL.n236 VSUBS 0.020971f
C1367 VTAIL.t13 VSUBS 0.070426f
C1368 VTAIL.n237 VSUBS 0.165202f
C1369 VTAIL.n238 VSUBS 1.38391f
C1370 VTAIL.n239 VSUBS 0.013947f
C1371 VTAIL.n240 VSUBS 0.014767f
C1372 VTAIL.n241 VSUBS 0.032966f
C1373 VTAIL.n242 VSUBS 0.032966f
C1374 VTAIL.n243 VSUBS 0.014767f
C1375 VTAIL.n244 VSUBS 0.013947f
C1376 VTAIL.n245 VSUBS 0.025955f
C1377 VTAIL.n246 VSUBS 0.025955f
C1378 VTAIL.n247 VSUBS 0.013947f
C1379 VTAIL.n248 VSUBS 0.014767f
C1380 VTAIL.n249 VSUBS 0.032966f
C1381 VTAIL.n250 VSUBS 0.032966f
C1382 VTAIL.n251 VSUBS 0.014767f
C1383 VTAIL.n252 VSUBS 0.013947f
C1384 VTAIL.n253 VSUBS 0.025955f
C1385 VTAIL.n254 VSUBS 0.025955f
C1386 VTAIL.n255 VSUBS 0.013947f
C1387 VTAIL.n256 VSUBS 0.014767f
C1388 VTAIL.n257 VSUBS 0.032966f
C1389 VTAIL.n258 VSUBS 0.032966f
C1390 VTAIL.n259 VSUBS 0.014767f
C1391 VTAIL.n260 VSUBS 0.013947f
C1392 VTAIL.n261 VSUBS 0.025955f
C1393 VTAIL.n262 VSUBS 0.025955f
C1394 VTAIL.n263 VSUBS 0.013947f
C1395 VTAIL.n264 VSUBS 0.014767f
C1396 VTAIL.n265 VSUBS 0.032966f
C1397 VTAIL.n266 VSUBS 0.032966f
C1398 VTAIL.n267 VSUBS 0.014767f
C1399 VTAIL.n268 VSUBS 0.013947f
C1400 VTAIL.n269 VSUBS 0.025955f
C1401 VTAIL.n270 VSUBS 0.025955f
C1402 VTAIL.n271 VSUBS 0.013947f
C1403 VTAIL.n272 VSUBS 0.014767f
C1404 VTAIL.n273 VSUBS 0.032966f
C1405 VTAIL.n274 VSUBS 0.032966f
C1406 VTAIL.n275 VSUBS 0.014767f
C1407 VTAIL.n276 VSUBS 0.013947f
C1408 VTAIL.n277 VSUBS 0.025955f
C1409 VTAIL.n278 VSUBS 0.067085f
C1410 VTAIL.n279 VSUBS 0.013947f
C1411 VTAIL.n280 VSUBS 0.014767f
C1412 VTAIL.n281 VSUBS 0.07494f
C1413 VTAIL.n282 VSUBS 0.049716f
C1414 VTAIL.n283 VSUBS 1.89816f
C1415 VTAIL.t8 VSUBS 0.260072f
C1416 VTAIL.t15 VSUBS 0.260072f
C1417 VTAIL.n284 VSUBS 1.94308f
C1418 VTAIL.n285 VSUBS 1.16793f
C1419 VTAIL.n286 VSUBS 0.014633f
C1420 VTAIL.n287 VSUBS 0.032966f
C1421 VTAIL.n288 VSUBS 0.014767f
C1422 VTAIL.n289 VSUBS 0.025955f
C1423 VTAIL.n290 VSUBS 0.013947f
C1424 VTAIL.n291 VSUBS 0.032966f
C1425 VTAIL.n292 VSUBS 0.014767f
C1426 VTAIL.n293 VSUBS 0.025955f
C1427 VTAIL.n294 VSUBS 0.013947f
C1428 VTAIL.n295 VSUBS 0.032966f
C1429 VTAIL.n296 VSUBS 0.014767f
C1430 VTAIL.n297 VSUBS 0.025955f
C1431 VTAIL.n298 VSUBS 0.013947f
C1432 VTAIL.n299 VSUBS 0.032966f
C1433 VTAIL.n300 VSUBS 0.014767f
C1434 VTAIL.n301 VSUBS 0.025955f
C1435 VTAIL.n302 VSUBS 0.013947f
C1436 VTAIL.n303 VSUBS 0.032966f
C1437 VTAIL.n304 VSUBS 0.014767f
C1438 VTAIL.n305 VSUBS 0.025955f
C1439 VTAIL.n306 VSUBS 0.013947f
C1440 VTAIL.n307 VSUBS 0.024724f
C1441 VTAIL.n308 VSUBS 0.020971f
C1442 VTAIL.t12 VSUBS 0.070426f
C1443 VTAIL.n309 VSUBS 0.165202f
C1444 VTAIL.n310 VSUBS 1.38391f
C1445 VTAIL.n311 VSUBS 0.013947f
C1446 VTAIL.n312 VSUBS 0.014767f
C1447 VTAIL.n313 VSUBS 0.032966f
C1448 VTAIL.n314 VSUBS 0.032966f
C1449 VTAIL.n315 VSUBS 0.014767f
C1450 VTAIL.n316 VSUBS 0.013947f
C1451 VTAIL.n317 VSUBS 0.025955f
C1452 VTAIL.n318 VSUBS 0.025955f
C1453 VTAIL.n319 VSUBS 0.013947f
C1454 VTAIL.n320 VSUBS 0.014767f
C1455 VTAIL.n321 VSUBS 0.032966f
C1456 VTAIL.n322 VSUBS 0.032966f
C1457 VTAIL.n323 VSUBS 0.014767f
C1458 VTAIL.n324 VSUBS 0.013947f
C1459 VTAIL.n325 VSUBS 0.025955f
C1460 VTAIL.n326 VSUBS 0.025955f
C1461 VTAIL.n327 VSUBS 0.013947f
C1462 VTAIL.n328 VSUBS 0.014767f
C1463 VTAIL.n329 VSUBS 0.032966f
C1464 VTAIL.n330 VSUBS 0.032966f
C1465 VTAIL.n331 VSUBS 0.014767f
C1466 VTAIL.n332 VSUBS 0.013947f
C1467 VTAIL.n333 VSUBS 0.025955f
C1468 VTAIL.n334 VSUBS 0.025955f
C1469 VTAIL.n335 VSUBS 0.013947f
C1470 VTAIL.n336 VSUBS 0.014767f
C1471 VTAIL.n337 VSUBS 0.032966f
C1472 VTAIL.n338 VSUBS 0.032966f
C1473 VTAIL.n339 VSUBS 0.014767f
C1474 VTAIL.n340 VSUBS 0.013947f
C1475 VTAIL.n341 VSUBS 0.025955f
C1476 VTAIL.n342 VSUBS 0.025955f
C1477 VTAIL.n343 VSUBS 0.013947f
C1478 VTAIL.n344 VSUBS 0.014767f
C1479 VTAIL.n345 VSUBS 0.032966f
C1480 VTAIL.n346 VSUBS 0.032966f
C1481 VTAIL.n347 VSUBS 0.014767f
C1482 VTAIL.n348 VSUBS 0.013947f
C1483 VTAIL.n349 VSUBS 0.025955f
C1484 VTAIL.n350 VSUBS 0.067085f
C1485 VTAIL.n351 VSUBS 0.013947f
C1486 VTAIL.n352 VSUBS 0.014767f
C1487 VTAIL.n353 VSUBS 0.07494f
C1488 VTAIL.n354 VSUBS 0.049716f
C1489 VTAIL.n355 VSUBS 0.36788f
C1490 VTAIL.n356 VSUBS 0.014633f
C1491 VTAIL.n357 VSUBS 0.032966f
C1492 VTAIL.n358 VSUBS 0.014767f
C1493 VTAIL.n359 VSUBS 0.025955f
C1494 VTAIL.n360 VSUBS 0.013947f
C1495 VTAIL.n361 VSUBS 0.032966f
C1496 VTAIL.n362 VSUBS 0.014767f
C1497 VTAIL.n363 VSUBS 0.025955f
C1498 VTAIL.n364 VSUBS 0.013947f
C1499 VTAIL.n365 VSUBS 0.032966f
C1500 VTAIL.n366 VSUBS 0.014767f
C1501 VTAIL.n367 VSUBS 0.025955f
C1502 VTAIL.n368 VSUBS 0.013947f
C1503 VTAIL.n369 VSUBS 0.032966f
C1504 VTAIL.n370 VSUBS 0.014767f
C1505 VTAIL.n371 VSUBS 0.025955f
C1506 VTAIL.n372 VSUBS 0.013947f
C1507 VTAIL.n373 VSUBS 0.032966f
C1508 VTAIL.n374 VSUBS 0.014767f
C1509 VTAIL.n375 VSUBS 0.025955f
C1510 VTAIL.n376 VSUBS 0.013947f
C1511 VTAIL.n377 VSUBS 0.024724f
C1512 VTAIL.n378 VSUBS 0.020971f
C1513 VTAIL.t0 VSUBS 0.070426f
C1514 VTAIL.n379 VSUBS 0.165202f
C1515 VTAIL.n380 VSUBS 1.38391f
C1516 VTAIL.n381 VSUBS 0.013947f
C1517 VTAIL.n382 VSUBS 0.014767f
C1518 VTAIL.n383 VSUBS 0.032966f
C1519 VTAIL.n384 VSUBS 0.032966f
C1520 VTAIL.n385 VSUBS 0.014767f
C1521 VTAIL.n386 VSUBS 0.013947f
C1522 VTAIL.n387 VSUBS 0.025955f
C1523 VTAIL.n388 VSUBS 0.025955f
C1524 VTAIL.n389 VSUBS 0.013947f
C1525 VTAIL.n390 VSUBS 0.014767f
C1526 VTAIL.n391 VSUBS 0.032966f
C1527 VTAIL.n392 VSUBS 0.032966f
C1528 VTAIL.n393 VSUBS 0.014767f
C1529 VTAIL.n394 VSUBS 0.013947f
C1530 VTAIL.n395 VSUBS 0.025955f
C1531 VTAIL.n396 VSUBS 0.025955f
C1532 VTAIL.n397 VSUBS 0.013947f
C1533 VTAIL.n398 VSUBS 0.014767f
C1534 VTAIL.n399 VSUBS 0.032966f
C1535 VTAIL.n400 VSUBS 0.032966f
C1536 VTAIL.n401 VSUBS 0.014767f
C1537 VTAIL.n402 VSUBS 0.013947f
C1538 VTAIL.n403 VSUBS 0.025955f
C1539 VTAIL.n404 VSUBS 0.025955f
C1540 VTAIL.n405 VSUBS 0.013947f
C1541 VTAIL.n406 VSUBS 0.014767f
C1542 VTAIL.n407 VSUBS 0.032966f
C1543 VTAIL.n408 VSUBS 0.032966f
C1544 VTAIL.n409 VSUBS 0.014767f
C1545 VTAIL.n410 VSUBS 0.013947f
C1546 VTAIL.n411 VSUBS 0.025955f
C1547 VTAIL.n412 VSUBS 0.025955f
C1548 VTAIL.n413 VSUBS 0.013947f
C1549 VTAIL.n414 VSUBS 0.014767f
C1550 VTAIL.n415 VSUBS 0.032966f
C1551 VTAIL.n416 VSUBS 0.032966f
C1552 VTAIL.n417 VSUBS 0.014767f
C1553 VTAIL.n418 VSUBS 0.013947f
C1554 VTAIL.n419 VSUBS 0.025955f
C1555 VTAIL.n420 VSUBS 0.067085f
C1556 VTAIL.n421 VSUBS 0.013947f
C1557 VTAIL.n422 VSUBS 0.014767f
C1558 VTAIL.n423 VSUBS 0.07494f
C1559 VTAIL.n424 VSUBS 0.049716f
C1560 VTAIL.n425 VSUBS 0.36788f
C1561 VTAIL.t2 VSUBS 0.260072f
C1562 VTAIL.t5 VSUBS 0.260072f
C1563 VTAIL.n426 VSUBS 1.94308f
C1564 VTAIL.n427 VSUBS 1.16793f
C1565 VTAIL.n428 VSUBS 0.014633f
C1566 VTAIL.n429 VSUBS 0.032966f
C1567 VTAIL.n430 VSUBS 0.014767f
C1568 VTAIL.n431 VSUBS 0.025955f
C1569 VTAIL.n432 VSUBS 0.013947f
C1570 VTAIL.n433 VSUBS 0.032966f
C1571 VTAIL.n434 VSUBS 0.014767f
C1572 VTAIL.n435 VSUBS 0.025955f
C1573 VTAIL.n436 VSUBS 0.013947f
C1574 VTAIL.n437 VSUBS 0.032966f
C1575 VTAIL.n438 VSUBS 0.014767f
C1576 VTAIL.n439 VSUBS 0.025955f
C1577 VTAIL.n440 VSUBS 0.013947f
C1578 VTAIL.n441 VSUBS 0.032966f
C1579 VTAIL.n442 VSUBS 0.014767f
C1580 VTAIL.n443 VSUBS 0.025955f
C1581 VTAIL.n444 VSUBS 0.013947f
C1582 VTAIL.n445 VSUBS 0.032966f
C1583 VTAIL.n446 VSUBS 0.014767f
C1584 VTAIL.n447 VSUBS 0.025955f
C1585 VTAIL.n448 VSUBS 0.013947f
C1586 VTAIL.n449 VSUBS 0.024724f
C1587 VTAIL.n450 VSUBS 0.020971f
C1588 VTAIL.t7 VSUBS 0.070426f
C1589 VTAIL.n451 VSUBS 0.165202f
C1590 VTAIL.n452 VSUBS 1.38391f
C1591 VTAIL.n453 VSUBS 0.013947f
C1592 VTAIL.n454 VSUBS 0.014767f
C1593 VTAIL.n455 VSUBS 0.032966f
C1594 VTAIL.n456 VSUBS 0.032966f
C1595 VTAIL.n457 VSUBS 0.014767f
C1596 VTAIL.n458 VSUBS 0.013947f
C1597 VTAIL.n459 VSUBS 0.025955f
C1598 VTAIL.n460 VSUBS 0.025955f
C1599 VTAIL.n461 VSUBS 0.013947f
C1600 VTAIL.n462 VSUBS 0.014767f
C1601 VTAIL.n463 VSUBS 0.032966f
C1602 VTAIL.n464 VSUBS 0.032966f
C1603 VTAIL.n465 VSUBS 0.014767f
C1604 VTAIL.n466 VSUBS 0.013947f
C1605 VTAIL.n467 VSUBS 0.025955f
C1606 VTAIL.n468 VSUBS 0.025955f
C1607 VTAIL.n469 VSUBS 0.013947f
C1608 VTAIL.n470 VSUBS 0.014767f
C1609 VTAIL.n471 VSUBS 0.032966f
C1610 VTAIL.n472 VSUBS 0.032966f
C1611 VTAIL.n473 VSUBS 0.014767f
C1612 VTAIL.n474 VSUBS 0.013947f
C1613 VTAIL.n475 VSUBS 0.025955f
C1614 VTAIL.n476 VSUBS 0.025955f
C1615 VTAIL.n477 VSUBS 0.013947f
C1616 VTAIL.n478 VSUBS 0.014767f
C1617 VTAIL.n479 VSUBS 0.032966f
C1618 VTAIL.n480 VSUBS 0.032966f
C1619 VTAIL.n481 VSUBS 0.014767f
C1620 VTAIL.n482 VSUBS 0.013947f
C1621 VTAIL.n483 VSUBS 0.025955f
C1622 VTAIL.n484 VSUBS 0.025955f
C1623 VTAIL.n485 VSUBS 0.013947f
C1624 VTAIL.n486 VSUBS 0.014767f
C1625 VTAIL.n487 VSUBS 0.032966f
C1626 VTAIL.n488 VSUBS 0.032966f
C1627 VTAIL.n489 VSUBS 0.014767f
C1628 VTAIL.n490 VSUBS 0.013947f
C1629 VTAIL.n491 VSUBS 0.025955f
C1630 VTAIL.n492 VSUBS 0.067085f
C1631 VTAIL.n493 VSUBS 0.013947f
C1632 VTAIL.n494 VSUBS 0.014767f
C1633 VTAIL.n495 VSUBS 0.07494f
C1634 VTAIL.n496 VSUBS 0.049716f
C1635 VTAIL.n497 VSUBS 1.89816f
C1636 VTAIL.n498 VSUBS 0.014633f
C1637 VTAIL.n499 VSUBS 0.032966f
C1638 VTAIL.n500 VSUBS 0.014767f
C1639 VTAIL.n501 VSUBS 0.025955f
C1640 VTAIL.n502 VSUBS 0.013947f
C1641 VTAIL.n503 VSUBS 0.032966f
C1642 VTAIL.n504 VSUBS 0.014767f
C1643 VTAIL.n505 VSUBS 0.025955f
C1644 VTAIL.n506 VSUBS 0.013947f
C1645 VTAIL.n507 VSUBS 0.032966f
C1646 VTAIL.n508 VSUBS 0.014767f
C1647 VTAIL.n509 VSUBS 0.025955f
C1648 VTAIL.n510 VSUBS 0.013947f
C1649 VTAIL.n511 VSUBS 0.032966f
C1650 VTAIL.n512 VSUBS 0.014767f
C1651 VTAIL.n513 VSUBS 0.025955f
C1652 VTAIL.n514 VSUBS 0.013947f
C1653 VTAIL.n515 VSUBS 0.032966f
C1654 VTAIL.n516 VSUBS 0.014767f
C1655 VTAIL.n517 VSUBS 0.025955f
C1656 VTAIL.n518 VSUBS 0.013947f
C1657 VTAIL.n519 VSUBS 0.024724f
C1658 VTAIL.n520 VSUBS 0.020971f
C1659 VTAIL.t11 VSUBS 0.070426f
C1660 VTAIL.n521 VSUBS 0.165202f
C1661 VTAIL.n522 VSUBS 1.38391f
C1662 VTAIL.n523 VSUBS 0.013947f
C1663 VTAIL.n524 VSUBS 0.014767f
C1664 VTAIL.n525 VSUBS 0.032966f
C1665 VTAIL.n526 VSUBS 0.032966f
C1666 VTAIL.n527 VSUBS 0.014767f
C1667 VTAIL.n528 VSUBS 0.013947f
C1668 VTAIL.n529 VSUBS 0.025955f
C1669 VTAIL.n530 VSUBS 0.025955f
C1670 VTAIL.n531 VSUBS 0.013947f
C1671 VTAIL.n532 VSUBS 0.014767f
C1672 VTAIL.n533 VSUBS 0.032966f
C1673 VTAIL.n534 VSUBS 0.032966f
C1674 VTAIL.n535 VSUBS 0.014767f
C1675 VTAIL.n536 VSUBS 0.013947f
C1676 VTAIL.n537 VSUBS 0.025955f
C1677 VTAIL.n538 VSUBS 0.025955f
C1678 VTAIL.n539 VSUBS 0.013947f
C1679 VTAIL.n540 VSUBS 0.014767f
C1680 VTAIL.n541 VSUBS 0.032966f
C1681 VTAIL.n542 VSUBS 0.032966f
C1682 VTAIL.n543 VSUBS 0.014767f
C1683 VTAIL.n544 VSUBS 0.013947f
C1684 VTAIL.n545 VSUBS 0.025955f
C1685 VTAIL.n546 VSUBS 0.025955f
C1686 VTAIL.n547 VSUBS 0.013947f
C1687 VTAIL.n548 VSUBS 0.014767f
C1688 VTAIL.n549 VSUBS 0.032966f
C1689 VTAIL.n550 VSUBS 0.032966f
C1690 VTAIL.n551 VSUBS 0.014767f
C1691 VTAIL.n552 VSUBS 0.013947f
C1692 VTAIL.n553 VSUBS 0.025955f
C1693 VTAIL.n554 VSUBS 0.025955f
C1694 VTAIL.n555 VSUBS 0.013947f
C1695 VTAIL.n556 VSUBS 0.014767f
C1696 VTAIL.n557 VSUBS 0.032966f
C1697 VTAIL.n558 VSUBS 0.032966f
C1698 VTAIL.n559 VSUBS 0.014767f
C1699 VTAIL.n560 VSUBS 0.013947f
C1700 VTAIL.n561 VSUBS 0.025955f
C1701 VTAIL.n562 VSUBS 0.067085f
C1702 VTAIL.n563 VSUBS 0.013947f
C1703 VTAIL.n564 VSUBS 0.014767f
C1704 VTAIL.n565 VSUBS 0.07494f
C1705 VTAIL.n566 VSUBS 0.049716f
C1706 VTAIL.n567 VSUBS 1.89329f
C1707 VDD2.t3 VSUBS 0.332414f
C1708 VDD2.t2 VSUBS 0.332414f
C1709 VDD2.n0 VSUBS 2.67526f
C1710 VDD2.t6 VSUBS 0.332414f
C1711 VDD2.t0 VSUBS 0.332414f
C1712 VDD2.n1 VSUBS 2.67526f
C1713 VDD2.n2 VSUBS 6.02566f
C1714 VDD2.t5 VSUBS 0.332414f
C1715 VDD2.t4 VSUBS 0.332414f
C1716 VDD2.n3 VSUBS 2.64865f
C1717 VDD2.n4 VSUBS 4.89374f
C1718 VDD2.t7 VSUBS 0.332414f
C1719 VDD2.t1 VSUBS 0.332414f
C1720 VDD2.n5 VSUBS 2.67519f
C1721 VN.t4 VSUBS 3.10402f
C1722 VN.n0 VSUBS 1.1712f
C1723 VN.n1 VSUBS 0.023181f
C1724 VN.n2 VSUBS 0.046559f
C1725 VN.n3 VSUBS 0.023181f
C1726 VN.n4 VSUBS 0.042986f
C1727 VN.n5 VSUBS 0.023181f
C1728 VN.t1 VSUBS 3.10402f
C1729 VN.n6 VSUBS 0.042986f
C1730 VN.n7 VSUBS 0.023181f
C1731 VN.n8 VSUBS 0.042986f
C1732 VN.t5 VSUBS 3.47659f
C1733 VN.n9 VSUBS 1.1129f
C1734 VN.t6 VSUBS 3.10402f
C1735 VN.n10 VSUBS 1.17146f
C1736 VN.n11 VSUBS 0.03662f
C1737 VN.n12 VSUBS 0.299931f
C1738 VN.n13 VSUBS 0.023181f
C1739 VN.n14 VSUBS 0.023181f
C1740 VN.n15 VSUBS 0.042986f
C1741 VN.n16 VSUBS 0.033696f
C1742 VN.n17 VSUBS 0.033696f
C1743 VN.n18 VSUBS 0.023181f
C1744 VN.n19 VSUBS 0.023181f
C1745 VN.n20 VSUBS 0.023181f
C1746 VN.n21 VSUBS 0.042986f
C1747 VN.n22 VSUBS 0.03662f
C1748 VN.n23 VSUBS 1.08383f
C1749 VN.n24 VSUBS 0.028131f
C1750 VN.n25 VSUBS 0.023181f
C1751 VN.n26 VSUBS 0.023181f
C1752 VN.n27 VSUBS 0.023181f
C1753 VN.n28 VSUBS 0.042986f
C1754 VN.n29 VSUBS 0.044349f
C1755 VN.n30 VSUBS 0.019472f
C1756 VN.n31 VSUBS 0.023181f
C1757 VN.n32 VSUBS 0.023181f
C1758 VN.n33 VSUBS 0.023181f
C1759 VN.n34 VSUBS 0.042986f
C1760 VN.n35 VSUBS 0.042986f
C1761 VN.n36 VSUBS 0.023887f
C1762 VN.n37 VSUBS 0.037407f
C1763 VN.n38 VSUBS 0.072316f
C1764 VN.t2 VSUBS 3.10402f
C1765 VN.n39 VSUBS 1.1712f
C1766 VN.n40 VSUBS 0.023181f
C1767 VN.n41 VSUBS 0.046559f
C1768 VN.n42 VSUBS 0.023181f
C1769 VN.n43 VSUBS 0.042986f
C1770 VN.n44 VSUBS 0.023181f
C1771 VN.t7 VSUBS 3.10402f
C1772 VN.n45 VSUBS 0.042986f
C1773 VN.n46 VSUBS 0.023181f
C1774 VN.n47 VSUBS 0.042986f
C1775 VN.t3 VSUBS 3.47659f
C1776 VN.n48 VSUBS 1.1129f
C1777 VN.t0 VSUBS 3.10402f
C1778 VN.n49 VSUBS 1.17146f
C1779 VN.n50 VSUBS 0.03662f
C1780 VN.n51 VSUBS 0.299931f
C1781 VN.n52 VSUBS 0.023181f
C1782 VN.n53 VSUBS 0.023181f
C1783 VN.n54 VSUBS 0.042986f
C1784 VN.n55 VSUBS 0.033696f
C1785 VN.n56 VSUBS 0.033696f
C1786 VN.n57 VSUBS 0.023181f
C1787 VN.n58 VSUBS 0.023181f
C1788 VN.n59 VSUBS 0.023181f
C1789 VN.n60 VSUBS 0.042986f
C1790 VN.n61 VSUBS 0.03662f
C1791 VN.n62 VSUBS 1.08383f
C1792 VN.n63 VSUBS 0.028131f
C1793 VN.n64 VSUBS 0.023181f
C1794 VN.n65 VSUBS 0.023181f
C1795 VN.n66 VSUBS 0.023181f
C1796 VN.n67 VSUBS 0.042986f
C1797 VN.n68 VSUBS 0.044349f
C1798 VN.n69 VSUBS 0.019472f
C1799 VN.n70 VSUBS 0.023181f
C1800 VN.n71 VSUBS 0.023181f
C1801 VN.n72 VSUBS 0.023181f
C1802 VN.n73 VSUBS 0.042986f
C1803 VN.n74 VSUBS 0.042986f
C1804 VN.n75 VSUBS 0.023887f
C1805 VN.n76 VSUBS 0.037407f
C1806 VN.n77 VSUBS 1.62548f
.ends

