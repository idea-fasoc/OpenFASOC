* NGSPICE file created from diff_pair_sample_0823.ext - technology: sky130A

.subckt diff_pair_sample_0823 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 w_n2610_n1240# sky130_fd_pr__pfet_01v8 ad=0.5304 pd=3.5 as=0.2244 ps=1.69 w=1.36 l=1.72
X1 VDD1.t4 VP.t1 VTAIL.t10 w_n2610_n1240# sky130_fd_pr__pfet_01v8 ad=0.5304 pd=3.5 as=0.2244 ps=1.69 w=1.36 l=1.72
X2 VDD2.t5 VN.t0 VTAIL.t4 w_n2610_n1240# sky130_fd_pr__pfet_01v8 ad=0.2244 pd=1.69 as=0.5304 ps=3.5 w=1.36 l=1.72
X3 B.t11 B.t9 B.t10 w_n2610_n1240# sky130_fd_pr__pfet_01v8 ad=0.5304 pd=3.5 as=0 ps=0 w=1.36 l=1.72
X4 B.t8 B.t6 B.t7 w_n2610_n1240# sky130_fd_pr__pfet_01v8 ad=0.5304 pd=3.5 as=0 ps=0 w=1.36 l=1.72
X5 VTAIL.t7 VP.t2 VDD1.t3 w_n2610_n1240# sky130_fd_pr__pfet_01v8 ad=0.2244 pd=1.69 as=0.2244 ps=1.69 w=1.36 l=1.72
X6 VDD1.t2 VP.t3 VTAIL.t6 w_n2610_n1240# sky130_fd_pr__pfet_01v8 ad=0.2244 pd=1.69 as=0.5304 ps=3.5 w=1.36 l=1.72
X7 VDD2.t4 VN.t1 VTAIL.t5 w_n2610_n1240# sky130_fd_pr__pfet_01v8 ad=0.2244 pd=1.69 as=0.5304 ps=3.5 w=1.36 l=1.72
X8 B.t5 B.t3 B.t4 w_n2610_n1240# sky130_fd_pr__pfet_01v8 ad=0.5304 pd=3.5 as=0 ps=0 w=1.36 l=1.72
X9 VDD2.t3 VN.t2 VTAIL.t0 w_n2610_n1240# sky130_fd_pr__pfet_01v8 ad=0.5304 pd=3.5 as=0.2244 ps=1.69 w=1.36 l=1.72
X10 VTAIL.t1 VN.t3 VDD2.t2 w_n2610_n1240# sky130_fd_pr__pfet_01v8 ad=0.2244 pd=1.69 as=0.2244 ps=1.69 w=1.36 l=1.72
X11 VDD1.t1 VP.t4 VTAIL.t9 w_n2610_n1240# sky130_fd_pr__pfet_01v8 ad=0.2244 pd=1.69 as=0.5304 ps=3.5 w=1.36 l=1.72
X12 VTAIL.t11 VP.t5 VDD1.t0 w_n2610_n1240# sky130_fd_pr__pfet_01v8 ad=0.2244 pd=1.69 as=0.2244 ps=1.69 w=1.36 l=1.72
X13 B.t2 B.t0 B.t1 w_n2610_n1240# sky130_fd_pr__pfet_01v8 ad=0.5304 pd=3.5 as=0 ps=0 w=1.36 l=1.72
X14 VDD2.t1 VN.t4 VTAIL.t2 w_n2610_n1240# sky130_fd_pr__pfet_01v8 ad=0.5304 pd=3.5 as=0.2244 ps=1.69 w=1.36 l=1.72
X15 VTAIL.t3 VN.t5 VDD2.t0 w_n2610_n1240# sky130_fd_pr__pfet_01v8 ad=0.2244 pd=1.69 as=0.2244 ps=1.69 w=1.36 l=1.72
R0 VP.n18 VP.n17 183.434
R1 VP.n33 VP.n32 183.434
R2 VP.n16 VP.n15 183.434
R3 VP.n10 VP.n9 161.3
R4 VP.n11 VP.n6 161.3
R5 VP.n13 VP.n12 161.3
R6 VP.n14 VP.n5 161.3
R7 VP.n31 VP.n0 161.3
R8 VP.n30 VP.n29 161.3
R9 VP.n28 VP.n1 161.3
R10 VP.n27 VP.n26 161.3
R11 VP.n25 VP.n2 161.3
R12 VP.n24 VP.n23 161.3
R13 VP.n22 VP.n3 161.3
R14 VP.n21 VP.n20 161.3
R15 VP.n19 VP.n4 161.3
R16 VP.n7 VP.t1 52.9651
R17 VP.n8 VP.n7 44.6952
R18 VP.n20 VP.n3 42.999
R19 VP.n30 VP.n1 42.999
R20 VP.n13 VP.n6 42.999
R21 VP.n24 VP.n3 38.1551
R22 VP.n26 VP.n1 38.1551
R23 VP.n9 VP.n6 38.1551
R24 VP.n17 VP.n16 37.027
R25 VP.n20 VP.n19 24.5923
R26 VP.n25 VP.n24 24.5923
R27 VP.n26 VP.n25 24.5923
R28 VP.n31 VP.n30 24.5923
R29 VP.n14 VP.n13 24.5923
R30 VP.n9 VP.n8 24.5923
R31 VP.n25 VP.t2 19.0563
R32 VP.n18 VP.t0 19.0563
R33 VP.n32 VP.t4 19.0563
R34 VP.n8 VP.t5 19.0563
R35 VP.n15 VP.t3 19.0563
R36 VP.n10 VP.n7 12.3444
R37 VP.n19 VP.n18 2.45968
R38 VP.n32 VP.n31 2.45968
R39 VP.n15 VP.n14 2.45968
R40 VP.n11 VP.n10 0.189894
R41 VP.n12 VP.n11 0.189894
R42 VP.n12 VP.n5 0.189894
R43 VP.n16 VP.n5 0.189894
R44 VP.n17 VP.n4 0.189894
R45 VP.n21 VP.n4 0.189894
R46 VP.n22 VP.n21 0.189894
R47 VP.n23 VP.n22 0.189894
R48 VP.n23 VP.n2 0.189894
R49 VP.n27 VP.n2 0.189894
R50 VP.n28 VP.n27 0.189894
R51 VP.n29 VP.n28 0.189894
R52 VP.n29 VP.n0 0.189894
R53 VP.n33 VP.n0 0.189894
R54 VP VP.n33 0.0516364
R55 VTAIL.n7 VTAIL.t5 255.459
R56 VTAIL.n11 VTAIL.t4 255.459
R57 VTAIL.n2 VTAIL.t9 255.459
R58 VTAIL.n10 VTAIL.t6 255.459
R59 VTAIL.n9 VTAIL.n8 231.559
R60 VTAIL.n6 VTAIL.n5 231.559
R61 VTAIL.n1 VTAIL.n0 231.559
R62 VTAIL.n4 VTAIL.n3 231.559
R63 VTAIL.n0 VTAIL.t2 23.9012
R64 VTAIL.n0 VTAIL.t1 23.9012
R65 VTAIL.n3 VTAIL.t8 23.9012
R66 VTAIL.n3 VTAIL.t7 23.9012
R67 VTAIL.n8 VTAIL.t10 23.9012
R68 VTAIL.n8 VTAIL.t11 23.9012
R69 VTAIL.n5 VTAIL.t0 23.9012
R70 VTAIL.n5 VTAIL.t3 23.9012
R71 VTAIL.n6 VTAIL.n4 17.0738
R72 VTAIL.n11 VTAIL.n10 15.3065
R73 VTAIL.n7 VTAIL.n6 1.76774
R74 VTAIL.n10 VTAIL.n9 1.76774
R75 VTAIL.n4 VTAIL.n2 1.76774
R76 VTAIL.n9 VTAIL.n7 1.35395
R77 VTAIL.n2 VTAIL.n1 1.35395
R78 VTAIL VTAIL.n11 1.26774
R79 VTAIL VTAIL.n1 0.5005
R80 VDD1 VDD1.t4 273.522
R81 VDD1.n1 VDD1.t5 273.409
R82 VDD1.n1 VDD1.n0 248.624
R83 VDD1.n3 VDD1.n2 248.238
R84 VDD1.n3 VDD1.n1 32.0979
R85 VDD1.n2 VDD1.t0 23.9012
R86 VDD1.n2 VDD1.t2 23.9012
R87 VDD1.n0 VDD1.t3 23.9012
R88 VDD1.n0 VDD1.t1 23.9012
R89 VDD1 VDD1.n3 0.384121
R90 VN.n11 VN.n10 183.434
R91 VN.n23 VN.n22 183.434
R92 VN.n21 VN.n12 161.3
R93 VN.n20 VN.n19 161.3
R94 VN.n18 VN.n13 161.3
R95 VN.n17 VN.n16 161.3
R96 VN.n9 VN.n0 161.3
R97 VN.n8 VN.n7 161.3
R98 VN.n6 VN.n1 161.3
R99 VN.n5 VN.n4 161.3
R100 VN.n2 VN.t4 52.9651
R101 VN.n14 VN.t1 52.9651
R102 VN.n15 VN.n14 44.6952
R103 VN.n3 VN.n2 44.6952
R104 VN.n8 VN.n1 42.999
R105 VN.n20 VN.n13 42.999
R106 VN.n4 VN.n1 38.1551
R107 VN.n16 VN.n13 38.1551
R108 VN VN.n23 37.4077
R109 VN.n4 VN.n3 24.5923
R110 VN.n9 VN.n8 24.5923
R111 VN.n16 VN.n15 24.5923
R112 VN.n21 VN.n20 24.5923
R113 VN.n3 VN.t3 19.0563
R114 VN.n10 VN.t0 19.0563
R115 VN.n15 VN.t5 19.0563
R116 VN.n22 VN.t2 19.0563
R117 VN.n17 VN.n14 12.3444
R118 VN.n5 VN.n2 12.3444
R119 VN.n10 VN.n9 2.45968
R120 VN.n22 VN.n21 2.45968
R121 VN.n23 VN.n12 0.189894
R122 VN.n19 VN.n12 0.189894
R123 VN.n19 VN.n18 0.189894
R124 VN.n18 VN.n17 0.189894
R125 VN.n6 VN.n5 0.189894
R126 VN.n7 VN.n6 0.189894
R127 VN.n7 VN.n0 0.189894
R128 VN.n11 VN.n0 0.189894
R129 VN VN.n11 0.0516364
R130 VDD2.n1 VDD2.t1 273.409
R131 VDD2.n2 VDD2.t3 272.139
R132 VDD2.n1 VDD2.n0 248.624
R133 VDD2 VDD2.n3 248.62
R134 VDD2.n2 VDD2.n1 30.6312
R135 VDD2.n3 VDD2.t0 23.9012
R136 VDD2.n3 VDD2.t4 23.9012
R137 VDD2.n0 VDD2.t2 23.9012
R138 VDD2.n0 VDD2.t5 23.9012
R139 VDD2 VDD2.n2 1.38412
R140 B.n296 B.n37 585
R141 B.n298 B.n297 585
R142 B.n299 B.n36 585
R143 B.n301 B.n300 585
R144 B.n302 B.n35 585
R145 B.n304 B.n303 585
R146 B.n305 B.n34 585
R147 B.n307 B.n306 585
R148 B.n308 B.n33 585
R149 B.n310 B.n309 585
R150 B.n312 B.n311 585
R151 B.n313 B.n29 585
R152 B.n315 B.n314 585
R153 B.n316 B.n28 585
R154 B.n318 B.n317 585
R155 B.n319 B.n27 585
R156 B.n321 B.n320 585
R157 B.n322 B.n26 585
R158 B.n324 B.n323 585
R159 B.n325 B.n23 585
R160 B.n328 B.n327 585
R161 B.n329 B.n22 585
R162 B.n331 B.n330 585
R163 B.n332 B.n21 585
R164 B.n334 B.n333 585
R165 B.n335 B.n20 585
R166 B.n337 B.n336 585
R167 B.n338 B.n19 585
R168 B.n340 B.n339 585
R169 B.n341 B.n18 585
R170 B.n295 B.n294 585
R171 B.n293 B.n38 585
R172 B.n292 B.n291 585
R173 B.n290 B.n39 585
R174 B.n289 B.n288 585
R175 B.n287 B.n40 585
R176 B.n286 B.n285 585
R177 B.n284 B.n41 585
R178 B.n283 B.n282 585
R179 B.n281 B.n42 585
R180 B.n280 B.n279 585
R181 B.n278 B.n43 585
R182 B.n277 B.n276 585
R183 B.n275 B.n44 585
R184 B.n274 B.n273 585
R185 B.n272 B.n45 585
R186 B.n271 B.n270 585
R187 B.n269 B.n46 585
R188 B.n268 B.n267 585
R189 B.n266 B.n47 585
R190 B.n265 B.n264 585
R191 B.n263 B.n48 585
R192 B.n262 B.n261 585
R193 B.n260 B.n49 585
R194 B.n259 B.n258 585
R195 B.n257 B.n50 585
R196 B.n256 B.n255 585
R197 B.n254 B.n51 585
R198 B.n253 B.n252 585
R199 B.n251 B.n52 585
R200 B.n250 B.n249 585
R201 B.n248 B.n53 585
R202 B.n247 B.n246 585
R203 B.n245 B.n54 585
R204 B.n244 B.n243 585
R205 B.n242 B.n55 585
R206 B.n241 B.n240 585
R207 B.n239 B.n56 585
R208 B.n238 B.n237 585
R209 B.n236 B.n57 585
R210 B.n235 B.n234 585
R211 B.n233 B.n58 585
R212 B.n232 B.n231 585
R213 B.n230 B.n59 585
R214 B.n229 B.n228 585
R215 B.n227 B.n60 585
R216 B.n226 B.n225 585
R217 B.n224 B.n61 585
R218 B.n223 B.n222 585
R219 B.n221 B.n62 585
R220 B.n220 B.n219 585
R221 B.n218 B.n63 585
R222 B.n217 B.n216 585
R223 B.n215 B.n64 585
R224 B.n214 B.n213 585
R225 B.n212 B.n65 585
R226 B.n211 B.n210 585
R227 B.n209 B.n66 585
R228 B.n208 B.n207 585
R229 B.n206 B.n67 585
R230 B.n205 B.n204 585
R231 B.n203 B.n68 585
R232 B.n202 B.n201 585
R233 B.n200 B.n69 585
R234 B.n199 B.n198 585
R235 B.n152 B.n89 585
R236 B.n154 B.n153 585
R237 B.n155 B.n88 585
R238 B.n157 B.n156 585
R239 B.n158 B.n87 585
R240 B.n160 B.n159 585
R241 B.n161 B.n86 585
R242 B.n163 B.n162 585
R243 B.n164 B.n85 585
R244 B.n166 B.n165 585
R245 B.n168 B.n167 585
R246 B.n169 B.n81 585
R247 B.n171 B.n170 585
R248 B.n172 B.n80 585
R249 B.n174 B.n173 585
R250 B.n175 B.n79 585
R251 B.n177 B.n176 585
R252 B.n178 B.n78 585
R253 B.n180 B.n179 585
R254 B.n181 B.n75 585
R255 B.n184 B.n183 585
R256 B.n185 B.n74 585
R257 B.n187 B.n186 585
R258 B.n188 B.n73 585
R259 B.n190 B.n189 585
R260 B.n191 B.n72 585
R261 B.n193 B.n192 585
R262 B.n194 B.n71 585
R263 B.n196 B.n195 585
R264 B.n197 B.n70 585
R265 B.n151 B.n150 585
R266 B.n149 B.n90 585
R267 B.n148 B.n147 585
R268 B.n146 B.n91 585
R269 B.n145 B.n144 585
R270 B.n143 B.n92 585
R271 B.n142 B.n141 585
R272 B.n140 B.n93 585
R273 B.n139 B.n138 585
R274 B.n137 B.n94 585
R275 B.n136 B.n135 585
R276 B.n134 B.n95 585
R277 B.n133 B.n132 585
R278 B.n131 B.n96 585
R279 B.n130 B.n129 585
R280 B.n128 B.n97 585
R281 B.n127 B.n126 585
R282 B.n125 B.n98 585
R283 B.n124 B.n123 585
R284 B.n122 B.n99 585
R285 B.n121 B.n120 585
R286 B.n119 B.n100 585
R287 B.n118 B.n117 585
R288 B.n116 B.n101 585
R289 B.n115 B.n114 585
R290 B.n113 B.n102 585
R291 B.n112 B.n111 585
R292 B.n110 B.n103 585
R293 B.n109 B.n108 585
R294 B.n107 B.n104 585
R295 B.n106 B.n105 585
R296 B.n2 B.n0 585
R297 B.n389 B.n1 585
R298 B.n388 B.n387 585
R299 B.n386 B.n3 585
R300 B.n385 B.n384 585
R301 B.n383 B.n4 585
R302 B.n382 B.n381 585
R303 B.n380 B.n5 585
R304 B.n379 B.n378 585
R305 B.n377 B.n6 585
R306 B.n376 B.n375 585
R307 B.n374 B.n7 585
R308 B.n373 B.n372 585
R309 B.n371 B.n8 585
R310 B.n370 B.n369 585
R311 B.n368 B.n9 585
R312 B.n367 B.n366 585
R313 B.n365 B.n10 585
R314 B.n364 B.n363 585
R315 B.n362 B.n11 585
R316 B.n361 B.n360 585
R317 B.n359 B.n12 585
R318 B.n358 B.n357 585
R319 B.n356 B.n13 585
R320 B.n355 B.n354 585
R321 B.n353 B.n14 585
R322 B.n352 B.n351 585
R323 B.n350 B.n15 585
R324 B.n349 B.n348 585
R325 B.n347 B.n16 585
R326 B.n346 B.n345 585
R327 B.n344 B.n17 585
R328 B.n343 B.n342 585
R329 B.n391 B.n390 585
R330 B.n150 B.n89 554.963
R331 B.n342 B.n341 554.963
R332 B.n198 B.n197 554.963
R333 B.n294 B.n37 554.963
R334 B.n76 B.t11 288.721
R335 B.n30 B.t7 288.721
R336 B.n82 B.t2 288.721
R337 B.n24 B.t4 288.721
R338 B.n77 B.t10 248.964
R339 B.n31 B.t8 248.964
R340 B.n83 B.t1 248.963
R341 B.n25 B.t5 248.963
R342 B.n76 B.t9 225.231
R343 B.n82 B.t0 225.231
R344 B.n24 B.t3 225.231
R345 B.n30 B.t6 225.231
R346 B.n150 B.n149 163.367
R347 B.n149 B.n148 163.367
R348 B.n148 B.n91 163.367
R349 B.n144 B.n91 163.367
R350 B.n144 B.n143 163.367
R351 B.n143 B.n142 163.367
R352 B.n142 B.n93 163.367
R353 B.n138 B.n93 163.367
R354 B.n138 B.n137 163.367
R355 B.n137 B.n136 163.367
R356 B.n136 B.n95 163.367
R357 B.n132 B.n95 163.367
R358 B.n132 B.n131 163.367
R359 B.n131 B.n130 163.367
R360 B.n130 B.n97 163.367
R361 B.n126 B.n97 163.367
R362 B.n126 B.n125 163.367
R363 B.n125 B.n124 163.367
R364 B.n124 B.n99 163.367
R365 B.n120 B.n99 163.367
R366 B.n120 B.n119 163.367
R367 B.n119 B.n118 163.367
R368 B.n118 B.n101 163.367
R369 B.n114 B.n101 163.367
R370 B.n114 B.n113 163.367
R371 B.n113 B.n112 163.367
R372 B.n112 B.n103 163.367
R373 B.n108 B.n103 163.367
R374 B.n108 B.n107 163.367
R375 B.n107 B.n106 163.367
R376 B.n106 B.n2 163.367
R377 B.n390 B.n2 163.367
R378 B.n390 B.n389 163.367
R379 B.n389 B.n388 163.367
R380 B.n388 B.n3 163.367
R381 B.n384 B.n3 163.367
R382 B.n384 B.n383 163.367
R383 B.n383 B.n382 163.367
R384 B.n382 B.n5 163.367
R385 B.n378 B.n5 163.367
R386 B.n378 B.n377 163.367
R387 B.n377 B.n376 163.367
R388 B.n376 B.n7 163.367
R389 B.n372 B.n7 163.367
R390 B.n372 B.n371 163.367
R391 B.n371 B.n370 163.367
R392 B.n370 B.n9 163.367
R393 B.n366 B.n9 163.367
R394 B.n366 B.n365 163.367
R395 B.n365 B.n364 163.367
R396 B.n364 B.n11 163.367
R397 B.n360 B.n11 163.367
R398 B.n360 B.n359 163.367
R399 B.n359 B.n358 163.367
R400 B.n358 B.n13 163.367
R401 B.n354 B.n13 163.367
R402 B.n354 B.n353 163.367
R403 B.n353 B.n352 163.367
R404 B.n352 B.n15 163.367
R405 B.n348 B.n15 163.367
R406 B.n348 B.n347 163.367
R407 B.n347 B.n346 163.367
R408 B.n346 B.n17 163.367
R409 B.n342 B.n17 163.367
R410 B.n154 B.n89 163.367
R411 B.n155 B.n154 163.367
R412 B.n156 B.n155 163.367
R413 B.n156 B.n87 163.367
R414 B.n160 B.n87 163.367
R415 B.n161 B.n160 163.367
R416 B.n162 B.n161 163.367
R417 B.n162 B.n85 163.367
R418 B.n166 B.n85 163.367
R419 B.n167 B.n166 163.367
R420 B.n167 B.n81 163.367
R421 B.n171 B.n81 163.367
R422 B.n172 B.n171 163.367
R423 B.n173 B.n172 163.367
R424 B.n173 B.n79 163.367
R425 B.n177 B.n79 163.367
R426 B.n178 B.n177 163.367
R427 B.n179 B.n178 163.367
R428 B.n179 B.n75 163.367
R429 B.n184 B.n75 163.367
R430 B.n185 B.n184 163.367
R431 B.n186 B.n185 163.367
R432 B.n186 B.n73 163.367
R433 B.n190 B.n73 163.367
R434 B.n191 B.n190 163.367
R435 B.n192 B.n191 163.367
R436 B.n192 B.n71 163.367
R437 B.n196 B.n71 163.367
R438 B.n197 B.n196 163.367
R439 B.n198 B.n69 163.367
R440 B.n202 B.n69 163.367
R441 B.n203 B.n202 163.367
R442 B.n204 B.n203 163.367
R443 B.n204 B.n67 163.367
R444 B.n208 B.n67 163.367
R445 B.n209 B.n208 163.367
R446 B.n210 B.n209 163.367
R447 B.n210 B.n65 163.367
R448 B.n214 B.n65 163.367
R449 B.n215 B.n214 163.367
R450 B.n216 B.n215 163.367
R451 B.n216 B.n63 163.367
R452 B.n220 B.n63 163.367
R453 B.n221 B.n220 163.367
R454 B.n222 B.n221 163.367
R455 B.n222 B.n61 163.367
R456 B.n226 B.n61 163.367
R457 B.n227 B.n226 163.367
R458 B.n228 B.n227 163.367
R459 B.n228 B.n59 163.367
R460 B.n232 B.n59 163.367
R461 B.n233 B.n232 163.367
R462 B.n234 B.n233 163.367
R463 B.n234 B.n57 163.367
R464 B.n238 B.n57 163.367
R465 B.n239 B.n238 163.367
R466 B.n240 B.n239 163.367
R467 B.n240 B.n55 163.367
R468 B.n244 B.n55 163.367
R469 B.n245 B.n244 163.367
R470 B.n246 B.n245 163.367
R471 B.n246 B.n53 163.367
R472 B.n250 B.n53 163.367
R473 B.n251 B.n250 163.367
R474 B.n252 B.n251 163.367
R475 B.n252 B.n51 163.367
R476 B.n256 B.n51 163.367
R477 B.n257 B.n256 163.367
R478 B.n258 B.n257 163.367
R479 B.n258 B.n49 163.367
R480 B.n262 B.n49 163.367
R481 B.n263 B.n262 163.367
R482 B.n264 B.n263 163.367
R483 B.n264 B.n47 163.367
R484 B.n268 B.n47 163.367
R485 B.n269 B.n268 163.367
R486 B.n270 B.n269 163.367
R487 B.n270 B.n45 163.367
R488 B.n274 B.n45 163.367
R489 B.n275 B.n274 163.367
R490 B.n276 B.n275 163.367
R491 B.n276 B.n43 163.367
R492 B.n280 B.n43 163.367
R493 B.n281 B.n280 163.367
R494 B.n282 B.n281 163.367
R495 B.n282 B.n41 163.367
R496 B.n286 B.n41 163.367
R497 B.n287 B.n286 163.367
R498 B.n288 B.n287 163.367
R499 B.n288 B.n39 163.367
R500 B.n292 B.n39 163.367
R501 B.n293 B.n292 163.367
R502 B.n294 B.n293 163.367
R503 B.n341 B.n340 163.367
R504 B.n340 B.n19 163.367
R505 B.n336 B.n19 163.367
R506 B.n336 B.n335 163.367
R507 B.n335 B.n334 163.367
R508 B.n334 B.n21 163.367
R509 B.n330 B.n21 163.367
R510 B.n330 B.n329 163.367
R511 B.n329 B.n328 163.367
R512 B.n328 B.n23 163.367
R513 B.n323 B.n23 163.367
R514 B.n323 B.n322 163.367
R515 B.n322 B.n321 163.367
R516 B.n321 B.n27 163.367
R517 B.n317 B.n27 163.367
R518 B.n317 B.n316 163.367
R519 B.n316 B.n315 163.367
R520 B.n315 B.n29 163.367
R521 B.n311 B.n29 163.367
R522 B.n311 B.n310 163.367
R523 B.n310 B.n33 163.367
R524 B.n306 B.n33 163.367
R525 B.n306 B.n305 163.367
R526 B.n305 B.n304 163.367
R527 B.n304 B.n35 163.367
R528 B.n300 B.n35 163.367
R529 B.n300 B.n299 163.367
R530 B.n299 B.n298 163.367
R531 B.n298 B.n37 163.367
R532 B.n182 B.n77 59.5399
R533 B.n84 B.n83 59.5399
R534 B.n326 B.n25 59.5399
R535 B.n32 B.n31 59.5399
R536 B.n77 B.n76 39.7581
R537 B.n83 B.n82 39.7581
R538 B.n25 B.n24 39.7581
R539 B.n31 B.n30 39.7581
R540 B.n296 B.n295 36.059
R541 B.n343 B.n18 36.059
R542 B.n199 B.n70 36.059
R543 B.n152 B.n151 36.059
R544 B B.n391 18.0485
R545 B.n339 B.n18 10.6151
R546 B.n339 B.n338 10.6151
R547 B.n338 B.n337 10.6151
R548 B.n337 B.n20 10.6151
R549 B.n333 B.n20 10.6151
R550 B.n333 B.n332 10.6151
R551 B.n332 B.n331 10.6151
R552 B.n331 B.n22 10.6151
R553 B.n327 B.n22 10.6151
R554 B.n325 B.n324 10.6151
R555 B.n324 B.n26 10.6151
R556 B.n320 B.n26 10.6151
R557 B.n320 B.n319 10.6151
R558 B.n319 B.n318 10.6151
R559 B.n318 B.n28 10.6151
R560 B.n314 B.n28 10.6151
R561 B.n314 B.n313 10.6151
R562 B.n313 B.n312 10.6151
R563 B.n309 B.n308 10.6151
R564 B.n308 B.n307 10.6151
R565 B.n307 B.n34 10.6151
R566 B.n303 B.n34 10.6151
R567 B.n303 B.n302 10.6151
R568 B.n302 B.n301 10.6151
R569 B.n301 B.n36 10.6151
R570 B.n297 B.n36 10.6151
R571 B.n297 B.n296 10.6151
R572 B.n200 B.n199 10.6151
R573 B.n201 B.n200 10.6151
R574 B.n201 B.n68 10.6151
R575 B.n205 B.n68 10.6151
R576 B.n206 B.n205 10.6151
R577 B.n207 B.n206 10.6151
R578 B.n207 B.n66 10.6151
R579 B.n211 B.n66 10.6151
R580 B.n212 B.n211 10.6151
R581 B.n213 B.n212 10.6151
R582 B.n213 B.n64 10.6151
R583 B.n217 B.n64 10.6151
R584 B.n218 B.n217 10.6151
R585 B.n219 B.n218 10.6151
R586 B.n219 B.n62 10.6151
R587 B.n223 B.n62 10.6151
R588 B.n224 B.n223 10.6151
R589 B.n225 B.n224 10.6151
R590 B.n225 B.n60 10.6151
R591 B.n229 B.n60 10.6151
R592 B.n230 B.n229 10.6151
R593 B.n231 B.n230 10.6151
R594 B.n231 B.n58 10.6151
R595 B.n235 B.n58 10.6151
R596 B.n236 B.n235 10.6151
R597 B.n237 B.n236 10.6151
R598 B.n237 B.n56 10.6151
R599 B.n241 B.n56 10.6151
R600 B.n242 B.n241 10.6151
R601 B.n243 B.n242 10.6151
R602 B.n243 B.n54 10.6151
R603 B.n247 B.n54 10.6151
R604 B.n248 B.n247 10.6151
R605 B.n249 B.n248 10.6151
R606 B.n249 B.n52 10.6151
R607 B.n253 B.n52 10.6151
R608 B.n254 B.n253 10.6151
R609 B.n255 B.n254 10.6151
R610 B.n255 B.n50 10.6151
R611 B.n259 B.n50 10.6151
R612 B.n260 B.n259 10.6151
R613 B.n261 B.n260 10.6151
R614 B.n261 B.n48 10.6151
R615 B.n265 B.n48 10.6151
R616 B.n266 B.n265 10.6151
R617 B.n267 B.n266 10.6151
R618 B.n267 B.n46 10.6151
R619 B.n271 B.n46 10.6151
R620 B.n272 B.n271 10.6151
R621 B.n273 B.n272 10.6151
R622 B.n273 B.n44 10.6151
R623 B.n277 B.n44 10.6151
R624 B.n278 B.n277 10.6151
R625 B.n279 B.n278 10.6151
R626 B.n279 B.n42 10.6151
R627 B.n283 B.n42 10.6151
R628 B.n284 B.n283 10.6151
R629 B.n285 B.n284 10.6151
R630 B.n285 B.n40 10.6151
R631 B.n289 B.n40 10.6151
R632 B.n290 B.n289 10.6151
R633 B.n291 B.n290 10.6151
R634 B.n291 B.n38 10.6151
R635 B.n295 B.n38 10.6151
R636 B.n153 B.n152 10.6151
R637 B.n153 B.n88 10.6151
R638 B.n157 B.n88 10.6151
R639 B.n158 B.n157 10.6151
R640 B.n159 B.n158 10.6151
R641 B.n159 B.n86 10.6151
R642 B.n163 B.n86 10.6151
R643 B.n164 B.n163 10.6151
R644 B.n165 B.n164 10.6151
R645 B.n169 B.n168 10.6151
R646 B.n170 B.n169 10.6151
R647 B.n170 B.n80 10.6151
R648 B.n174 B.n80 10.6151
R649 B.n175 B.n174 10.6151
R650 B.n176 B.n175 10.6151
R651 B.n176 B.n78 10.6151
R652 B.n180 B.n78 10.6151
R653 B.n181 B.n180 10.6151
R654 B.n183 B.n74 10.6151
R655 B.n187 B.n74 10.6151
R656 B.n188 B.n187 10.6151
R657 B.n189 B.n188 10.6151
R658 B.n189 B.n72 10.6151
R659 B.n193 B.n72 10.6151
R660 B.n194 B.n193 10.6151
R661 B.n195 B.n194 10.6151
R662 B.n195 B.n70 10.6151
R663 B.n151 B.n90 10.6151
R664 B.n147 B.n90 10.6151
R665 B.n147 B.n146 10.6151
R666 B.n146 B.n145 10.6151
R667 B.n145 B.n92 10.6151
R668 B.n141 B.n92 10.6151
R669 B.n141 B.n140 10.6151
R670 B.n140 B.n139 10.6151
R671 B.n139 B.n94 10.6151
R672 B.n135 B.n94 10.6151
R673 B.n135 B.n134 10.6151
R674 B.n134 B.n133 10.6151
R675 B.n133 B.n96 10.6151
R676 B.n129 B.n96 10.6151
R677 B.n129 B.n128 10.6151
R678 B.n128 B.n127 10.6151
R679 B.n127 B.n98 10.6151
R680 B.n123 B.n98 10.6151
R681 B.n123 B.n122 10.6151
R682 B.n122 B.n121 10.6151
R683 B.n121 B.n100 10.6151
R684 B.n117 B.n100 10.6151
R685 B.n117 B.n116 10.6151
R686 B.n116 B.n115 10.6151
R687 B.n115 B.n102 10.6151
R688 B.n111 B.n102 10.6151
R689 B.n111 B.n110 10.6151
R690 B.n110 B.n109 10.6151
R691 B.n109 B.n104 10.6151
R692 B.n105 B.n104 10.6151
R693 B.n105 B.n0 10.6151
R694 B.n387 B.n1 10.6151
R695 B.n387 B.n386 10.6151
R696 B.n386 B.n385 10.6151
R697 B.n385 B.n4 10.6151
R698 B.n381 B.n4 10.6151
R699 B.n381 B.n380 10.6151
R700 B.n380 B.n379 10.6151
R701 B.n379 B.n6 10.6151
R702 B.n375 B.n6 10.6151
R703 B.n375 B.n374 10.6151
R704 B.n374 B.n373 10.6151
R705 B.n373 B.n8 10.6151
R706 B.n369 B.n8 10.6151
R707 B.n369 B.n368 10.6151
R708 B.n368 B.n367 10.6151
R709 B.n367 B.n10 10.6151
R710 B.n363 B.n10 10.6151
R711 B.n363 B.n362 10.6151
R712 B.n362 B.n361 10.6151
R713 B.n361 B.n12 10.6151
R714 B.n357 B.n12 10.6151
R715 B.n357 B.n356 10.6151
R716 B.n356 B.n355 10.6151
R717 B.n355 B.n14 10.6151
R718 B.n351 B.n14 10.6151
R719 B.n351 B.n350 10.6151
R720 B.n350 B.n349 10.6151
R721 B.n349 B.n16 10.6151
R722 B.n345 B.n16 10.6151
R723 B.n345 B.n344 10.6151
R724 B.n344 B.n343 10.6151
R725 B.n327 B.n326 9.36635
R726 B.n309 B.n32 9.36635
R727 B.n165 B.n84 9.36635
R728 B.n183 B.n182 9.36635
R729 B.n391 B.n0 2.81026
R730 B.n391 B.n1 2.81026
R731 B.n326 B.n325 1.24928
R732 B.n312 B.n32 1.24928
R733 B.n168 B.n84 1.24928
R734 B.n182 B.n181 1.24928
C0 VN VTAIL 1.6435f
C1 VDD1 VP 1.25804f
C2 VDD2 VTAIL 3.30206f
C3 VDD2 VN 1.02613f
C4 B VTAIL 0.992004f
C5 B VN 0.832334f
C6 w_n2610_n1240# VTAIL 1.30179f
C7 w_n2610_n1240# VN 4.5132f
C8 VDD2 B 1.08949f
C9 VDD2 w_n2610_n1240# 1.36546f
C10 VDD1 VTAIL 3.25483f
C11 B w_n2610_n1240# 5.50199f
C12 VP VTAIL 1.65763f
C13 VDD1 VN 0.15703f
C14 VP VN 4.10701f
C15 VDD1 VDD2 1.08724f
C16 VDD2 VP 0.391342f
C17 VDD1 B 1.03607f
C18 B VP 1.38615f
C19 VDD1 w_n2610_n1240# 1.30952f
C20 w_n2610_n1240# VP 4.84159f
C21 VDD2 VSUBS 0.824369f
C22 VDD1 VSUBS 1.171798f
C23 VTAIL VSUBS 0.352677f
C24 VN VSUBS 4.39944f
C25 VP VSUBS 1.678105f
C26 B VSUBS 2.709837f
C27 w_n2610_n1240# VSUBS 41.561604f
C28 B.n0 VSUBS 0.006075f
C29 B.n1 VSUBS 0.006075f
C30 B.n2 VSUBS 0.009607f
C31 B.n3 VSUBS 0.009607f
C32 B.n4 VSUBS 0.009607f
C33 B.n5 VSUBS 0.009607f
C34 B.n6 VSUBS 0.009607f
C35 B.n7 VSUBS 0.009607f
C36 B.n8 VSUBS 0.009607f
C37 B.n9 VSUBS 0.009607f
C38 B.n10 VSUBS 0.009607f
C39 B.n11 VSUBS 0.009607f
C40 B.n12 VSUBS 0.009607f
C41 B.n13 VSUBS 0.009607f
C42 B.n14 VSUBS 0.009607f
C43 B.n15 VSUBS 0.009607f
C44 B.n16 VSUBS 0.009607f
C45 B.n17 VSUBS 0.009607f
C46 B.n18 VSUBS 0.024608f
C47 B.n19 VSUBS 0.009607f
C48 B.n20 VSUBS 0.009607f
C49 B.n21 VSUBS 0.009607f
C50 B.n22 VSUBS 0.009607f
C51 B.n23 VSUBS 0.009607f
C52 B.t5 VSUBS 0.037406f
C53 B.t4 VSUBS 0.044453f
C54 B.t3 VSUBS 0.159911f
C55 B.n24 VSUBS 0.076249f
C56 B.n25 VSUBS 0.064877f
C57 B.n26 VSUBS 0.009607f
C58 B.n27 VSUBS 0.009607f
C59 B.n28 VSUBS 0.009607f
C60 B.n29 VSUBS 0.009607f
C61 B.t8 VSUBS 0.037406f
C62 B.t7 VSUBS 0.044453f
C63 B.t6 VSUBS 0.159911f
C64 B.n30 VSUBS 0.076249f
C65 B.n31 VSUBS 0.064877f
C66 B.n32 VSUBS 0.022259f
C67 B.n33 VSUBS 0.009607f
C68 B.n34 VSUBS 0.009607f
C69 B.n35 VSUBS 0.009607f
C70 B.n36 VSUBS 0.009607f
C71 B.n37 VSUBS 0.024608f
C72 B.n38 VSUBS 0.009607f
C73 B.n39 VSUBS 0.009607f
C74 B.n40 VSUBS 0.009607f
C75 B.n41 VSUBS 0.009607f
C76 B.n42 VSUBS 0.009607f
C77 B.n43 VSUBS 0.009607f
C78 B.n44 VSUBS 0.009607f
C79 B.n45 VSUBS 0.009607f
C80 B.n46 VSUBS 0.009607f
C81 B.n47 VSUBS 0.009607f
C82 B.n48 VSUBS 0.009607f
C83 B.n49 VSUBS 0.009607f
C84 B.n50 VSUBS 0.009607f
C85 B.n51 VSUBS 0.009607f
C86 B.n52 VSUBS 0.009607f
C87 B.n53 VSUBS 0.009607f
C88 B.n54 VSUBS 0.009607f
C89 B.n55 VSUBS 0.009607f
C90 B.n56 VSUBS 0.009607f
C91 B.n57 VSUBS 0.009607f
C92 B.n58 VSUBS 0.009607f
C93 B.n59 VSUBS 0.009607f
C94 B.n60 VSUBS 0.009607f
C95 B.n61 VSUBS 0.009607f
C96 B.n62 VSUBS 0.009607f
C97 B.n63 VSUBS 0.009607f
C98 B.n64 VSUBS 0.009607f
C99 B.n65 VSUBS 0.009607f
C100 B.n66 VSUBS 0.009607f
C101 B.n67 VSUBS 0.009607f
C102 B.n68 VSUBS 0.009607f
C103 B.n69 VSUBS 0.009607f
C104 B.n70 VSUBS 0.024608f
C105 B.n71 VSUBS 0.009607f
C106 B.n72 VSUBS 0.009607f
C107 B.n73 VSUBS 0.009607f
C108 B.n74 VSUBS 0.009607f
C109 B.n75 VSUBS 0.009607f
C110 B.t10 VSUBS 0.037406f
C111 B.t11 VSUBS 0.044453f
C112 B.t9 VSUBS 0.159911f
C113 B.n76 VSUBS 0.076249f
C114 B.n77 VSUBS 0.064877f
C115 B.n78 VSUBS 0.009607f
C116 B.n79 VSUBS 0.009607f
C117 B.n80 VSUBS 0.009607f
C118 B.n81 VSUBS 0.009607f
C119 B.t1 VSUBS 0.037406f
C120 B.t2 VSUBS 0.044453f
C121 B.t0 VSUBS 0.159911f
C122 B.n82 VSUBS 0.076249f
C123 B.n83 VSUBS 0.064877f
C124 B.n84 VSUBS 0.022259f
C125 B.n85 VSUBS 0.009607f
C126 B.n86 VSUBS 0.009607f
C127 B.n87 VSUBS 0.009607f
C128 B.n88 VSUBS 0.009607f
C129 B.n89 VSUBS 0.024608f
C130 B.n90 VSUBS 0.009607f
C131 B.n91 VSUBS 0.009607f
C132 B.n92 VSUBS 0.009607f
C133 B.n93 VSUBS 0.009607f
C134 B.n94 VSUBS 0.009607f
C135 B.n95 VSUBS 0.009607f
C136 B.n96 VSUBS 0.009607f
C137 B.n97 VSUBS 0.009607f
C138 B.n98 VSUBS 0.009607f
C139 B.n99 VSUBS 0.009607f
C140 B.n100 VSUBS 0.009607f
C141 B.n101 VSUBS 0.009607f
C142 B.n102 VSUBS 0.009607f
C143 B.n103 VSUBS 0.009607f
C144 B.n104 VSUBS 0.009607f
C145 B.n105 VSUBS 0.009607f
C146 B.n106 VSUBS 0.009607f
C147 B.n107 VSUBS 0.009607f
C148 B.n108 VSUBS 0.009607f
C149 B.n109 VSUBS 0.009607f
C150 B.n110 VSUBS 0.009607f
C151 B.n111 VSUBS 0.009607f
C152 B.n112 VSUBS 0.009607f
C153 B.n113 VSUBS 0.009607f
C154 B.n114 VSUBS 0.009607f
C155 B.n115 VSUBS 0.009607f
C156 B.n116 VSUBS 0.009607f
C157 B.n117 VSUBS 0.009607f
C158 B.n118 VSUBS 0.009607f
C159 B.n119 VSUBS 0.009607f
C160 B.n120 VSUBS 0.009607f
C161 B.n121 VSUBS 0.009607f
C162 B.n122 VSUBS 0.009607f
C163 B.n123 VSUBS 0.009607f
C164 B.n124 VSUBS 0.009607f
C165 B.n125 VSUBS 0.009607f
C166 B.n126 VSUBS 0.009607f
C167 B.n127 VSUBS 0.009607f
C168 B.n128 VSUBS 0.009607f
C169 B.n129 VSUBS 0.009607f
C170 B.n130 VSUBS 0.009607f
C171 B.n131 VSUBS 0.009607f
C172 B.n132 VSUBS 0.009607f
C173 B.n133 VSUBS 0.009607f
C174 B.n134 VSUBS 0.009607f
C175 B.n135 VSUBS 0.009607f
C176 B.n136 VSUBS 0.009607f
C177 B.n137 VSUBS 0.009607f
C178 B.n138 VSUBS 0.009607f
C179 B.n139 VSUBS 0.009607f
C180 B.n140 VSUBS 0.009607f
C181 B.n141 VSUBS 0.009607f
C182 B.n142 VSUBS 0.009607f
C183 B.n143 VSUBS 0.009607f
C184 B.n144 VSUBS 0.009607f
C185 B.n145 VSUBS 0.009607f
C186 B.n146 VSUBS 0.009607f
C187 B.n147 VSUBS 0.009607f
C188 B.n148 VSUBS 0.009607f
C189 B.n149 VSUBS 0.009607f
C190 B.n150 VSUBS 0.023429f
C191 B.n151 VSUBS 0.023429f
C192 B.n152 VSUBS 0.024608f
C193 B.n153 VSUBS 0.009607f
C194 B.n154 VSUBS 0.009607f
C195 B.n155 VSUBS 0.009607f
C196 B.n156 VSUBS 0.009607f
C197 B.n157 VSUBS 0.009607f
C198 B.n158 VSUBS 0.009607f
C199 B.n159 VSUBS 0.009607f
C200 B.n160 VSUBS 0.009607f
C201 B.n161 VSUBS 0.009607f
C202 B.n162 VSUBS 0.009607f
C203 B.n163 VSUBS 0.009607f
C204 B.n164 VSUBS 0.009607f
C205 B.n165 VSUBS 0.009042f
C206 B.n166 VSUBS 0.009607f
C207 B.n167 VSUBS 0.009607f
C208 B.n168 VSUBS 0.005369f
C209 B.n169 VSUBS 0.009607f
C210 B.n170 VSUBS 0.009607f
C211 B.n171 VSUBS 0.009607f
C212 B.n172 VSUBS 0.009607f
C213 B.n173 VSUBS 0.009607f
C214 B.n174 VSUBS 0.009607f
C215 B.n175 VSUBS 0.009607f
C216 B.n176 VSUBS 0.009607f
C217 B.n177 VSUBS 0.009607f
C218 B.n178 VSUBS 0.009607f
C219 B.n179 VSUBS 0.009607f
C220 B.n180 VSUBS 0.009607f
C221 B.n181 VSUBS 0.005369f
C222 B.n182 VSUBS 0.022259f
C223 B.n183 VSUBS 0.009042f
C224 B.n184 VSUBS 0.009607f
C225 B.n185 VSUBS 0.009607f
C226 B.n186 VSUBS 0.009607f
C227 B.n187 VSUBS 0.009607f
C228 B.n188 VSUBS 0.009607f
C229 B.n189 VSUBS 0.009607f
C230 B.n190 VSUBS 0.009607f
C231 B.n191 VSUBS 0.009607f
C232 B.n192 VSUBS 0.009607f
C233 B.n193 VSUBS 0.009607f
C234 B.n194 VSUBS 0.009607f
C235 B.n195 VSUBS 0.009607f
C236 B.n196 VSUBS 0.009607f
C237 B.n197 VSUBS 0.024608f
C238 B.n198 VSUBS 0.023429f
C239 B.n199 VSUBS 0.023429f
C240 B.n200 VSUBS 0.009607f
C241 B.n201 VSUBS 0.009607f
C242 B.n202 VSUBS 0.009607f
C243 B.n203 VSUBS 0.009607f
C244 B.n204 VSUBS 0.009607f
C245 B.n205 VSUBS 0.009607f
C246 B.n206 VSUBS 0.009607f
C247 B.n207 VSUBS 0.009607f
C248 B.n208 VSUBS 0.009607f
C249 B.n209 VSUBS 0.009607f
C250 B.n210 VSUBS 0.009607f
C251 B.n211 VSUBS 0.009607f
C252 B.n212 VSUBS 0.009607f
C253 B.n213 VSUBS 0.009607f
C254 B.n214 VSUBS 0.009607f
C255 B.n215 VSUBS 0.009607f
C256 B.n216 VSUBS 0.009607f
C257 B.n217 VSUBS 0.009607f
C258 B.n218 VSUBS 0.009607f
C259 B.n219 VSUBS 0.009607f
C260 B.n220 VSUBS 0.009607f
C261 B.n221 VSUBS 0.009607f
C262 B.n222 VSUBS 0.009607f
C263 B.n223 VSUBS 0.009607f
C264 B.n224 VSUBS 0.009607f
C265 B.n225 VSUBS 0.009607f
C266 B.n226 VSUBS 0.009607f
C267 B.n227 VSUBS 0.009607f
C268 B.n228 VSUBS 0.009607f
C269 B.n229 VSUBS 0.009607f
C270 B.n230 VSUBS 0.009607f
C271 B.n231 VSUBS 0.009607f
C272 B.n232 VSUBS 0.009607f
C273 B.n233 VSUBS 0.009607f
C274 B.n234 VSUBS 0.009607f
C275 B.n235 VSUBS 0.009607f
C276 B.n236 VSUBS 0.009607f
C277 B.n237 VSUBS 0.009607f
C278 B.n238 VSUBS 0.009607f
C279 B.n239 VSUBS 0.009607f
C280 B.n240 VSUBS 0.009607f
C281 B.n241 VSUBS 0.009607f
C282 B.n242 VSUBS 0.009607f
C283 B.n243 VSUBS 0.009607f
C284 B.n244 VSUBS 0.009607f
C285 B.n245 VSUBS 0.009607f
C286 B.n246 VSUBS 0.009607f
C287 B.n247 VSUBS 0.009607f
C288 B.n248 VSUBS 0.009607f
C289 B.n249 VSUBS 0.009607f
C290 B.n250 VSUBS 0.009607f
C291 B.n251 VSUBS 0.009607f
C292 B.n252 VSUBS 0.009607f
C293 B.n253 VSUBS 0.009607f
C294 B.n254 VSUBS 0.009607f
C295 B.n255 VSUBS 0.009607f
C296 B.n256 VSUBS 0.009607f
C297 B.n257 VSUBS 0.009607f
C298 B.n258 VSUBS 0.009607f
C299 B.n259 VSUBS 0.009607f
C300 B.n260 VSUBS 0.009607f
C301 B.n261 VSUBS 0.009607f
C302 B.n262 VSUBS 0.009607f
C303 B.n263 VSUBS 0.009607f
C304 B.n264 VSUBS 0.009607f
C305 B.n265 VSUBS 0.009607f
C306 B.n266 VSUBS 0.009607f
C307 B.n267 VSUBS 0.009607f
C308 B.n268 VSUBS 0.009607f
C309 B.n269 VSUBS 0.009607f
C310 B.n270 VSUBS 0.009607f
C311 B.n271 VSUBS 0.009607f
C312 B.n272 VSUBS 0.009607f
C313 B.n273 VSUBS 0.009607f
C314 B.n274 VSUBS 0.009607f
C315 B.n275 VSUBS 0.009607f
C316 B.n276 VSUBS 0.009607f
C317 B.n277 VSUBS 0.009607f
C318 B.n278 VSUBS 0.009607f
C319 B.n279 VSUBS 0.009607f
C320 B.n280 VSUBS 0.009607f
C321 B.n281 VSUBS 0.009607f
C322 B.n282 VSUBS 0.009607f
C323 B.n283 VSUBS 0.009607f
C324 B.n284 VSUBS 0.009607f
C325 B.n285 VSUBS 0.009607f
C326 B.n286 VSUBS 0.009607f
C327 B.n287 VSUBS 0.009607f
C328 B.n288 VSUBS 0.009607f
C329 B.n289 VSUBS 0.009607f
C330 B.n290 VSUBS 0.009607f
C331 B.n291 VSUBS 0.009607f
C332 B.n292 VSUBS 0.009607f
C333 B.n293 VSUBS 0.009607f
C334 B.n294 VSUBS 0.023429f
C335 B.n295 VSUBS 0.024457f
C336 B.n296 VSUBS 0.02358f
C337 B.n297 VSUBS 0.009607f
C338 B.n298 VSUBS 0.009607f
C339 B.n299 VSUBS 0.009607f
C340 B.n300 VSUBS 0.009607f
C341 B.n301 VSUBS 0.009607f
C342 B.n302 VSUBS 0.009607f
C343 B.n303 VSUBS 0.009607f
C344 B.n304 VSUBS 0.009607f
C345 B.n305 VSUBS 0.009607f
C346 B.n306 VSUBS 0.009607f
C347 B.n307 VSUBS 0.009607f
C348 B.n308 VSUBS 0.009607f
C349 B.n309 VSUBS 0.009042f
C350 B.n310 VSUBS 0.009607f
C351 B.n311 VSUBS 0.009607f
C352 B.n312 VSUBS 0.005369f
C353 B.n313 VSUBS 0.009607f
C354 B.n314 VSUBS 0.009607f
C355 B.n315 VSUBS 0.009607f
C356 B.n316 VSUBS 0.009607f
C357 B.n317 VSUBS 0.009607f
C358 B.n318 VSUBS 0.009607f
C359 B.n319 VSUBS 0.009607f
C360 B.n320 VSUBS 0.009607f
C361 B.n321 VSUBS 0.009607f
C362 B.n322 VSUBS 0.009607f
C363 B.n323 VSUBS 0.009607f
C364 B.n324 VSUBS 0.009607f
C365 B.n325 VSUBS 0.005369f
C366 B.n326 VSUBS 0.022259f
C367 B.n327 VSUBS 0.009042f
C368 B.n328 VSUBS 0.009607f
C369 B.n329 VSUBS 0.009607f
C370 B.n330 VSUBS 0.009607f
C371 B.n331 VSUBS 0.009607f
C372 B.n332 VSUBS 0.009607f
C373 B.n333 VSUBS 0.009607f
C374 B.n334 VSUBS 0.009607f
C375 B.n335 VSUBS 0.009607f
C376 B.n336 VSUBS 0.009607f
C377 B.n337 VSUBS 0.009607f
C378 B.n338 VSUBS 0.009607f
C379 B.n339 VSUBS 0.009607f
C380 B.n340 VSUBS 0.009607f
C381 B.n341 VSUBS 0.024608f
C382 B.n342 VSUBS 0.023429f
C383 B.n343 VSUBS 0.023429f
C384 B.n344 VSUBS 0.009607f
C385 B.n345 VSUBS 0.009607f
C386 B.n346 VSUBS 0.009607f
C387 B.n347 VSUBS 0.009607f
C388 B.n348 VSUBS 0.009607f
C389 B.n349 VSUBS 0.009607f
C390 B.n350 VSUBS 0.009607f
C391 B.n351 VSUBS 0.009607f
C392 B.n352 VSUBS 0.009607f
C393 B.n353 VSUBS 0.009607f
C394 B.n354 VSUBS 0.009607f
C395 B.n355 VSUBS 0.009607f
C396 B.n356 VSUBS 0.009607f
C397 B.n357 VSUBS 0.009607f
C398 B.n358 VSUBS 0.009607f
C399 B.n359 VSUBS 0.009607f
C400 B.n360 VSUBS 0.009607f
C401 B.n361 VSUBS 0.009607f
C402 B.n362 VSUBS 0.009607f
C403 B.n363 VSUBS 0.009607f
C404 B.n364 VSUBS 0.009607f
C405 B.n365 VSUBS 0.009607f
C406 B.n366 VSUBS 0.009607f
C407 B.n367 VSUBS 0.009607f
C408 B.n368 VSUBS 0.009607f
C409 B.n369 VSUBS 0.009607f
C410 B.n370 VSUBS 0.009607f
C411 B.n371 VSUBS 0.009607f
C412 B.n372 VSUBS 0.009607f
C413 B.n373 VSUBS 0.009607f
C414 B.n374 VSUBS 0.009607f
C415 B.n375 VSUBS 0.009607f
C416 B.n376 VSUBS 0.009607f
C417 B.n377 VSUBS 0.009607f
C418 B.n378 VSUBS 0.009607f
C419 B.n379 VSUBS 0.009607f
C420 B.n380 VSUBS 0.009607f
C421 B.n381 VSUBS 0.009607f
C422 B.n382 VSUBS 0.009607f
C423 B.n383 VSUBS 0.009607f
C424 B.n384 VSUBS 0.009607f
C425 B.n385 VSUBS 0.009607f
C426 B.n386 VSUBS 0.009607f
C427 B.n387 VSUBS 0.009607f
C428 B.n388 VSUBS 0.009607f
C429 B.n389 VSUBS 0.009607f
C430 B.n390 VSUBS 0.009607f
C431 B.n391 VSUBS 0.021754f
C432 VDD2.t1 VSUBS 0.114371f
C433 VDD2.t2 VSUBS 0.018779f
C434 VDD2.t5 VSUBS 0.018779f
C435 VDD2.n0 VSUBS 0.071575f
C436 VDD2.n1 VSUBS 1.3134f
C437 VDD2.t3 VSUBS 0.113257f
C438 VDD2.n2 VSUBS 1.16149f
C439 VDD2.t0 VSUBS 0.018779f
C440 VDD2.t4 VSUBS 0.018779f
C441 VDD2.n3 VSUBS 0.07157f
C442 VN.n0 VSUBS 0.05007f
C443 VN.t0 VSUBS 0.247786f
C444 VN.n1 VSUBS 0.04084f
C445 VN.t4 VSUBS 0.492658f
C446 VN.n2 VSUBS 0.228912f
C447 VN.t3 VSUBS 0.247786f
C448 VN.n3 VSUBS 0.287189f
C449 VN.n4 VSUBS 0.100019f
C450 VN.n5 VSUBS 0.364525f
C451 VN.n6 VSUBS 0.05007f
C452 VN.n7 VSUBS 0.05007f
C453 VN.n8 VSUBS 0.09756f
C454 VN.n9 VSUBS 0.051596f
C455 VN.n10 VSUBS 0.258662f
C456 VN.n11 VSUBS 0.052992f
C457 VN.n12 VSUBS 0.05007f
C458 VN.t2 VSUBS 0.247786f
C459 VN.n13 VSUBS 0.04084f
C460 VN.t1 VSUBS 0.492658f
C461 VN.n14 VSUBS 0.228912f
C462 VN.t5 VSUBS 0.247786f
C463 VN.n15 VSUBS 0.287189f
C464 VN.n16 VSUBS 0.100019f
C465 VN.n17 VSUBS 0.364525f
C466 VN.n18 VSUBS 0.05007f
C467 VN.n19 VSUBS 0.05007f
C468 VN.n20 VSUBS 0.09756f
C469 VN.n21 VSUBS 0.051596f
C470 VN.n22 VSUBS 0.258662f
C471 VN.n23 VSUBS 1.70584f
C472 VDD1.t4 VSUBS 0.112305f
C473 VDD1.t5 VSUBS 0.112178f
C474 VDD1.t3 VSUBS 0.018419f
C475 VDD1.t1 VSUBS 0.018419f
C476 VDD1.n0 VSUBS 0.070202f
C477 VDD1.n1 VSUBS 1.35146f
C478 VDD1.t0 VSUBS 0.018419f
C479 VDD1.t2 VSUBS 0.018419f
C480 VDD1.n2 VSUBS 0.069773f
C481 VDD1.n3 VSUBS 1.17271f
C482 VTAIL.t2 VSUBS 0.025494f
C483 VTAIL.t1 VSUBS 0.025494f
C484 VTAIL.n0 VSUBS 0.082038f
C485 VTAIL.n1 VSUBS 0.330332f
C486 VTAIL.t9 VSUBS 0.139772f
C487 VTAIL.n2 VSUBS 0.438991f
C488 VTAIL.t8 VSUBS 0.025494f
C489 VTAIL.t7 VSUBS 0.025494f
C490 VTAIL.n3 VSUBS 0.082038f
C491 VTAIL.n4 VSUBS 1.00575f
C492 VTAIL.t0 VSUBS 0.025494f
C493 VTAIL.t3 VSUBS 0.025494f
C494 VTAIL.n5 VSUBS 0.082038f
C495 VTAIL.n6 VSUBS 1.00575f
C496 VTAIL.t5 VSUBS 0.139772f
C497 VTAIL.n7 VSUBS 0.438991f
C498 VTAIL.t10 VSUBS 0.025494f
C499 VTAIL.t11 VSUBS 0.025494f
C500 VTAIL.n8 VSUBS 0.082038f
C501 VTAIL.n9 VSUBS 0.427195f
C502 VTAIL.t6 VSUBS 0.139772f
C503 VTAIL.n10 VSUBS 0.882466f
C504 VTAIL.t4 VSUBS 0.139772f
C505 VTAIL.n11 VSUBS 0.844248f
C506 VP.n0 VSUBS 0.052244f
C507 VP.t4 VSUBS 0.258545f
C508 VP.n1 VSUBS 0.042614f
C509 VP.n2 VSUBS 0.052244f
C510 VP.t2 VSUBS 0.258545f
C511 VP.n3 VSUBS 0.042614f
C512 VP.n4 VSUBS 0.052244f
C513 VP.t0 VSUBS 0.258545f
C514 VP.n5 VSUBS 0.052244f
C515 VP.t3 VSUBS 0.258545f
C516 VP.n6 VSUBS 0.042614f
C517 VP.t1 VSUBS 0.51405f
C518 VP.n7 VSUBS 0.238852f
C519 VP.t5 VSUBS 0.258545f
C520 VP.n8 VSUBS 0.29966f
C521 VP.n9 VSUBS 0.104363f
C522 VP.n10 VSUBS 0.380354f
C523 VP.n11 VSUBS 0.052244f
C524 VP.n12 VSUBS 0.052244f
C525 VP.n13 VSUBS 0.101796f
C526 VP.n14 VSUBS 0.053837f
C527 VP.n15 VSUBS 0.269894f
C528 VP.n16 VSUBS 1.74532f
C529 VP.n17 VSUBS 1.79619f
C530 VP.n18 VSUBS 0.269894f
C531 VP.n19 VSUBS 0.053837f
C532 VP.n20 VSUBS 0.101796f
C533 VP.n21 VSUBS 0.052244f
C534 VP.n22 VSUBS 0.052244f
C535 VP.n23 VSUBS 0.052244f
C536 VP.n24 VSUBS 0.104363f
C537 VP.n25 VSUBS 0.211045f
C538 VP.n26 VSUBS 0.104363f
C539 VP.n27 VSUBS 0.052244f
C540 VP.n28 VSUBS 0.052244f
C541 VP.n29 VSUBS 0.052244f
C542 VP.n30 VSUBS 0.101796f
C543 VP.n31 VSUBS 0.053837f
C544 VP.n32 VSUBS 0.269894f
C545 VP.n33 VSUBS 0.055293f
.ends

