* NGSPICE file created from diff_pair_sample_0591.ext - technology: sky130A

.subckt diff_pair_sample_0591 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=1.443 pd=8.18 as=0 ps=0 w=3.7 l=1.44
X1 VDD1.t7 VP.t0 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=0.6105 pd=4.03 as=0.6105 ps=4.03 w=3.7 l=1.44
X2 VTAIL.t2 VN.t0 VDD2.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=0.6105 pd=4.03 as=0.6105 ps=4.03 w=3.7 l=1.44
X3 VDD1.t6 VP.t1 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=0.6105 pd=4.03 as=1.443 ps=8.18 w=3.7 l=1.44
X4 VDD1.t5 VP.t2 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=0.6105 pd=4.03 as=0.6105 ps=4.03 w=3.7 l=1.44
X5 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=1.443 pd=8.18 as=0 ps=0 w=3.7 l=1.44
X6 VTAIL.t3 VN.t1 VDD2.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=0.6105 pd=4.03 as=0.6105 ps=4.03 w=3.7 l=1.44
X7 VDD2.t5 VN.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.6105 pd=4.03 as=1.443 ps=8.18 w=3.7 l=1.44
X8 VTAIL.t12 VP.t3 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=1.443 pd=8.18 as=0.6105 ps=4.03 w=3.7 l=1.44
X9 VDD1.t3 VP.t4 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=0.6105 pd=4.03 as=1.443 ps=8.18 w=3.7 l=1.44
X10 VDD2.t4 VN.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.6105 pd=4.03 as=1.443 ps=8.18 w=3.7 l=1.44
X11 VTAIL.t7 VN.t4 VDD2.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=1.443 pd=8.18 as=0.6105 ps=4.03 w=3.7 l=1.44
X12 VTAIL.t13 VP.t5 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=0.6105 pd=4.03 as=0.6105 ps=4.03 w=3.7 l=1.44
X13 VDD2.t2 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.6105 pd=4.03 as=0.6105 ps=4.03 w=3.7 l=1.44
X14 VTAIL.t14 VP.t6 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.443 pd=8.18 as=0.6105 ps=4.03 w=3.7 l=1.44
X15 VTAIL.t1 VN.t6 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.443 pd=8.18 as=0.6105 ps=4.03 w=3.7 l=1.44
X16 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=1.443 pd=8.18 as=0 ps=0 w=3.7 l=1.44
X17 VDD2.t0 VN.t7 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.6105 pd=4.03 as=0.6105 ps=4.03 w=3.7 l=1.44
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.443 pd=8.18 as=0 ps=0 w=3.7 l=1.44
X19 VTAIL.t15 VP.t7 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.6105 pd=4.03 as=0.6105 ps=4.03 w=3.7 l=1.44
R0 B.n419 B.n418 585
R1 B.n421 B.n91 585
R2 B.n424 B.n423 585
R3 B.n425 B.n90 585
R4 B.n427 B.n426 585
R5 B.n429 B.n89 585
R6 B.n432 B.n431 585
R7 B.n433 B.n88 585
R8 B.n435 B.n434 585
R9 B.n437 B.n87 585
R10 B.n440 B.n439 585
R11 B.n441 B.n86 585
R12 B.n443 B.n442 585
R13 B.n445 B.n85 585
R14 B.n448 B.n447 585
R15 B.n449 B.n81 585
R16 B.n451 B.n450 585
R17 B.n453 B.n80 585
R18 B.n456 B.n455 585
R19 B.n457 B.n79 585
R20 B.n459 B.n458 585
R21 B.n461 B.n78 585
R22 B.n464 B.n463 585
R23 B.n465 B.n77 585
R24 B.n467 B.n466 585
R25 B.n469 B.n76 585
R26 B.n472 B.n471 585
R27 B.n474 B.n73 585
R28 B.n476 B.n475 585
R29 B.n478 B.n72 585
R30 B.n481 B.n480 585
R31 B.n482 B.n71 585
R32 B.n484 B.n483 585
R33 B.n486 B.n70 585
R34 B.n489 B.n488 585
R35 B.n490 B.n69 585
R36 B.n492 B.n491 585
R37 B.n494 B.n68 585
R38 B.n497 B.n496 585
R39 B.n498 B.n67 585
R40 B.n500 B.n499 585
R41 B.n502 B.n66 585
R42 B.n505 B.n504 585
R43 B.n506 B.n65 585
R44 B.n417 B.n63 585
R45 B.n509 B.n63 585
R46 B.n416 B.n62 585
R47 B.n510 B.n62 585
R48 B.n415 B.n61 585
R49 B.n511 B.n61 585
R50 B.n414 B.n413 585
R51 B.n413 B.n57 585
R52 B.n412 B.n56 585
R53 B.n517 B.n56 585
R54 B.n411 B.n55 585
R55 B.n518 B.n55 585
R56 B.n410 B.n54 585
R57 B.n519 B.n54 585
R58 B.n409 B.n408 585
R59 B.n408 B.n50 585
R60 B.n407 B.n49 585
R61 B.n525 B.n49 585
R62 B.n406 B.n48 585
R63 B.n526 B.n48 585
R64 B.n405 B.n47 585
R65 B.n527 B.n47 585
R66 B.n404 B.n403 585
R67 B.n403 B.n43 585
R68 B.n402 B.n42 585
R69 B.n533 B.n42 585
R70 B.n401 B.n41 585
R71 B.n534 B.n41 585
R72 B.n400 B.n40 585
R73 B.n535 B.n40 585
R74 B.n399 B.n398 585
R75 B.n398 B.n36 585
R76 B.n397 B.n35 585
R77 B.n541 B.n35 585
R78 B.n396 B.n34 585
R79 B.n542 B.n34 585
R80 B.n395 B.n33 585
R81 B.n543 B.n33 585
R82 B.n394 B.n393 585
R83 B.n393 B.n32 585
R84 B.n392 B.n28 585
R85 B.n549 B.n28 585
R86 B.n391 B.n27 585
R87 B.n550 B.n27 585
R88 B.n390 B.n26 585
R89 B.n551 B.n26 585
R90 B.n389 B.n388 585
R91 B.n388 B.n22 585
R92 B.n387 B.n21 585
R93 B.n557 B.n21 585
R94 B.n386 B.n20 585
R95 B.n558 B.n20 585
R96 B.n385 B.n19 585
R97 B.n559 B.n19 585
R98 B.n384 B.n383 585
R99 B.n383 B.n15 585
R100 B.n382 B.n14 585
R101 B.n565 B.n14 585
R102 B.n381 B.n13 585
R103 B.n566 B.n13 585
R104 B.n380 B.n12 585
R105 B.n567 B.n12 585
R106 B.n379 B.n378 585
R107 B.n378 B.n8 585
R108 B.n377 B.n7 585
R109 B.n573 B.n7 585
R110 B.n376 B.n6 585
R111 B.n574 B.n6 585
R112 B.n375 B.n5 585
R113 B.n575 B.n5 585
R114 B.n374 B.n373 585
R115 B.n373 B.n4 585
R116 B.n372 B.n92 585
R117 B.n372 B.n371 585
R118 B.n362 B.n93 585
R119 B.n94 B.n93 585
R120 B.n364 B.n363 585
R121 B.n365 B.n364 585
R122 B.n361 B.n98 585
R123 B.n102 B.n98 585
R124 B.n360 B.n359 585
R125 B.n359 B.n358 585
R126 B.n100 B.n99 585
R127 B.n101 B.n100 585
R128 B.n351 B.n350 585
R129 B.n352 B.n351 585
R130 B.n349 B.n107 585
R131 B.n107 B.n106 585
R132 B.n348 B.n347 585
R133 B.n347 B.n346 585
R134 B.n109 B.n108 585
R135 B.n110 B.n109 585
R136 B.n339 B.n338 585
R137 B.n340 B.n339 585
R138 B.n337 B.n115 585
R139 B.n115 B.n114 585
R140 B.n336 B.n335 585
R141 B.n335 B.n334 585
R142 B.n117 B.n116 585
R143 B.n327 B.n117 585
R144 B.n326 B.n325 585
R145 B.n328 B.n326 585
R146 B.n324 B.n122 585
R147 B.n122 B.n121 585
R148 B.n323 B.n322 585
R149 B.n322 B.n321 585
R150 B.n124 B.n123 585
R151 B.n125 B.n124 585
R152 B.n314 B.n313 585
R153 B.n315 B.n314 585
R154 B.n312 B.n130 585
R155 B.n130 B.n129 585
R156 B.n311 B.n310 585
R157 B.n310 B.n309 585
R158 B.n132 B.n131 585
R159 B.n133 B.n132 585
R160 B.n302 B.n301 585
R161 B.n303 B.n302 585
R162 B.n300 B.n138 585
R163 B.n138 B.n137 585
R164 B.n299 B.n298 585
R165 B.n298 B.n297 585
R166 B.n140 B.n139 585
R167 B.n141 B.n140 585
R168 B.n290 B.n289 585
R169 B.n291 B.n290 585
R170 B.n288 B.n145 585
R171 B.n149 B.n145 585
R172 B.n287 B.n286 585
R173 B.n286 B.n285 585
R174 B.n147 B.n146 585
R175 B.n148 B.n147 585
R176 B.n278 B.n277 585
R177 B.n279 B.n278 585
R178 B.n276 B.n154 585
R179 B.n154 B.n153 585
R180 B.n275 B.n274 585
R181 B.n274 B.n273 585
R182 B.n270 B.n158 585
R183 B.n269 B.n268 585
R184 B.n266 B.n159 585
R185 B.n266 B.n157 585
R186 B.n265 B.n264 585
R187 B.n263 B.n262 585
R188 B.n261 B.n161 585
R189 B.n259 B.n258 585
R190 B.n257 B.n162 585
R191 B.n256 B.n255 585
R192 B.n253 B.n163 585
R193 B.n251 B.n250 585
R194 B.n249 B.n164 585
R195 B.n248 B.n247 585
R196 B.n245 B.n165 585
R197 B.n243 B.n242 585
R198 B.n241 B.n166 585
R199 B.n240 B.n239 585
R200 B.n237 B.n236 585
R201 B.n235 B.n234 585
R202 B.n233 B.n171 585
R203 B.n231 B.n230 585
R204 B.n229 B.n172 585
R205 B.n228 B.n227 585
R206 B.n225 B.n173 585
R207 B.n223 B.n222 585
R208 B.n221 B.n174 585
R209 B.n220 B.n219 585
R210 B.n217 B.n216 585
R211 B.n215 B.n214 585
R212 B.n213 B.n179 585
R213 B.n211 B.n210 585
R214 B.n209 B.n180 585
R215 B.n208 B.n207 585
R216 B.n205 B.n181 585
R217 B.n203 B.n202 585
R218 B.n201 B.n182 585
R219 B.n200 B.n199 585
R220 B.n197 B.n183 585
R221 B.n195 B.n194 585
R222 B.n193 B.n184 585
R223 B.n192 B.n191 585
R224 B.n189 B.n185 585
R225 B.n187 B.n186 585
R226 B.n156 B.n155 585
R227 B.n157 B.n156 585
R228 B.n272 B.n271 585
R229 B.n273 B.n272 585
R230 B.n152 B.n151 585
R231 B.n153 B.n152 585
R232 B.n281 B.n280 585
R233 B.n280 B.n279 585
R234 B.n282 B.n150 585
R235 B.n150 B.n148 585
R236 B.n284 B.n283 585
R237 B.n285 B.n284 585
R238 B.n144 B.n143 585
R239 B.n149 B.n144 585
R240 B.n293 B.n292 585
R241 B.n292 B.n291 585
R242 B.n294 B.n142 585
R243 B.n142 B.n141 585
R244 B.n296 B.n295 585
R245 B.n297 B.n296 585
R246 B.n136 B.n135 585
R247 B.n137 B.n136 585
R248 B.n305 B.n304 585
R249 B.n304 B.n303 585
R250 B.n306 B.n134 585
R251 B.n134 B.n133 585
R252 B.n308 B.n307 585
R253 B.n309 B.n308 585
R254 B.n128 B.n127 585
R255 B.n129 B.n128 585
R256 B.n317 B.n316 585
R257 B.n316 B.n315 585
R258 B.n318 B.n126 585
R259 B.n126 B.n125 585
R260 B.n320 B.n319 585
R261 B.n321 B.n320 585
R262 B.n120 B.n119 585
R263 B.n121 B.n120 585
R264 B.n330 B.n329 585
R265 B.n329 B.n328 585
R266 B.n331 B.n118 585
R267 B.n327 B.n118 585
R268 B.n333 B.n332 585
R269 B.n334 B.n333 585
R270 B.n113 B.n112 585
R271 B.n114 B.n113 585
R272 B.n342 B.n341 585
R273 B.n341 B.n340 585
R274 B.n343 B.n111 585
R275 B.n111 B.n110 585
R276 B.n345 B.n344 585
R277 B.n346 B.n345 585
R278 B.n105 B.n104 585
R279 B.n106 B.n105 585
R280 B.n354 B.n353 585
R281 B.n353 B.n352 585
R282 B.n355 B.n103 585
R283 B.n103 B.n101 585
R284 B.n357 B.n356 585
R285 B.n358 B.n357 585
R286 B.n97 B.n96 585
R287 B.n102 B.n97 585
R288 B.n367 B.n366 585
R289 B.n366 B.n365 585
R290 B.n368 B.n95 585
R291 B.n95 B.n94 585
R292 B.n370 B.n369 585
R293 B.n371 B.n370 585
R294 B.n2 B.n0 585
R295 B.n4 B.n2 585
R296 B.n3 B.n1 585
R297 B.n574 B.n3 585
R298 B.n572 B.n571 585
R299 B.n573 B.n572 585
R300 B.n570 B.n9 585
R301 B.n9 B.n8 585
R302 B.n569 B.n568 585
R303 B.n568 B.n567 585
R304 B.n11 B.n10 585
R305 B.n566 B.n11 585
R306 B.n564 B.n563 585
R307 B.n565 B.n564 585
R308 B.n562 B.n16 585
R309 B.n16 B.n15 585
R310 B.n561 B.n560 585
R311 B.n560 B.n559 585
R312 B.n18 B.n17 585
R313 B.n558 B.n18 585
R314 B.n556 B.n555 585
R315 B.n557 B.n556 585
R316 B.n554 B.n23 585
R317 B.n23 B.n22 585
R318 B.n553 B.n552 585
R319 B.n552 B.n551 585
R320 B.n25 B.n24 585
R321 B.n550 B.n25 585
R322 B.n548 B.n547 585
R323 B.n549 B.n548 585
R324 B.n546 B.n29 585
R325 B.n32 B.n29 585
R326 B.n545 B.n544 585
R327 B.n544 B.n543 585
R328 B.n31 B.n30 585
R329 B.n542 B.n31 585
R330 B.n540 B.n539 585
R331 B.n541 B.n540 585
R332 B.n538 B.n37 585
R333 B.n37 B.n36 585
R334 B.n537 B.n536 585
R335 B.n536 B.n535 585
R336 B.n39 B.n38 585
R337 B.n534 B.n39 585
R338 B.n532 B.n531 585
R339 B.n533 B.n532 585
R340 B.n530 B.n44 585
R341 B.n44 B.n43 585
R342 B.n529 B.n528 585
R343 B.n528 B.n527 585
R344 B.n46 B.n45 585
R345 B.n526 B.n46 585
R346 B.n524 B.n523 585
R347 B.n525 B.n524 585
R348 B.n522 B.n51 585
R349 B.n51 B.n50 585
R350 B.n521 B.n520 585
R351 B.n520 B.n519 585
R352 B.n53 B.n52 585
R353 B.n518 B.n53 585
R354 B.n516 B.n515 585
R355 B.n517 B.n516 585
R356 B.n514 B.n58 585
R357 B.n58 B.n57 585
R358 B.n513 B.n512 585
R359 B.n512 B.n511 585
R360 B.n60 B.n59 585
R361 B.n510 B.n60 585
R362 B.n508 B.n507 585
R363 B.n509 B.n508 585
R364 B.n577 B.n576 585
R365 B.n576 B.n575 585
R366 B.n272 B.n158 521.33
R367 B.n508 B.n65 521.33
R368 B.n274 B.n156 521.33
R369 B.n419 B.n63 521.33
R370 B.n175 B.t19 267.132
R371 B.n167 B.t12 267.132
R372 B.n74 B.t16 267.132
R373 B.n82 B.t8 267.132
R374 B.n420 B.n64 256.663
R375 B.n422 B.n64 256.663
R376 B.n428 B.n64 256.663
R377 B.n430 B.n64 256.663
R378 B.n436 B.n64 256.663
R379 B.n438 B.n64 256.663
R380 B.n444 B.n64 256.663
R381 B.n446 B.n64 256.663
R382 B.n452 B.n64 256.663
R383 B.n454 B.n64 256.663
R384 B.n460 B.n64 256.663
R385 B.n462 B.n64 256.663
R386 B.n468 B.n64 256.663
R387 B.n470 B.n64 256.663
R388 B.n477 B.n64 256.663
R389 B.n479 B.n64 256.663
R390 B.n485 B.n64 256.663
R391 B.n487 B.n64 256.663
R392 B.n493 B.n64 256.663
R393 B.n495 B.n64 256.663
R394 B.n501 B.n64 256.663
R395 B.n503 B.n64 256.663
R396 B.n267 B.n157 256.663
R397 B.n160 B.n157 256.663
R398 B.n260 B.n157 256.663
R399 B.n254 B.n157 256.663
R400 B.n252 B.n157 256.663
R401 B.n246 B.n157 256.663
R402 B.n244 B.n157 256.663
R403 B.n238 B.n157 256.663
R404 B.n170 B.n157 256.663
R405 B.n232 B.n157 256.663
R406 B.n226 B.n157 256.663
R407 B.n224 B.n157 256.663
R408 B.n218 B.n157 256.663
R409 B.n178 B.n157 256.663
R410 B.n212 B.n157 256.663
R411 B.n206 B.n157 256.663
R412 B.n204 B.n157 256.663
R413 B.n198 B.n157 256.663
R414 B.n196 B.n157 256.663
R415 B.n190 B.n157 256.663
R416 B.n188 B.n157 256.663
R417 B.n272 B.n152 163.367
R418 B.n280 B.n152 163.367
R419 B.n280 B.n150 163.367
R420 B.n284 B.n150 163.367
R421 B.n284 B.n144 163.367
R422 B.n292 B.n144 163.367
R423 B.n292 B.n142 163.367
R424 B.n296 B.n142 163.367
R425 B.n296 B.n136 163.367
R426 B.n304 B.n136 163.367
R427 B.n304 B.n134 163.367
R428 B.n308 B.n134 163.367
R429 B.n308 B.n128 163.367
R430 B.n316 B.n128 163.367
R431 B.n316 B.n126 163.367
R432 B.n320 B.n126 163.367
R433 B.n320 B.n120 163.367
R434 B.n329 B.n120 163.367
R435 B.n329 B.n118 163.367
R436 B.n333 B.n118 163.367
R437 B.n333 B.n113 163.367
R438 B.n341 B.n113 163.367
R439 B.n341 B.n111 163.367
R440 B.n345 B.n111 163.367
R441 B.n345 B.n105 163.367
R442 B.n353 B.n105 163.367
R443 B.n353 B.n103 163.367
R444 B.n357 B.n103 163.367
R445 B.n357 B.n97 163.367
R446 B.n366 B.n97 163.367
R447 B.n366 B.n95 163.367
R448 B.n370 B.n95 163.367
R449 B.n370 B.n2 163.367
R450 B.n576 B.n2 163.367
R451 B.n576 B.n3 163.367
R452 B.n572 B.n3 163.367
R453 B.n572 B.n9 163.367
R454 B.n568 B.n9 163.367
R455 B.n568 B.n11 163.367
R456 B.n564 B.n11 163.367
R457 B.n564 B.n16 163.367
R458 B.n560 B.n16 163.367
R459 B.n560 B.n18 163.367
R460 B.n556 B.n18 163.367
R461 B.n556 B.n23 163.367
R462 B.n552 B.n23 163.367
R463 B.n552 B.n25 163.367
R464 B.n548 B.n25 163.367
R465 B.n548 B.n29 163.367
R466 B.n544 B.n29 163.367
R467 B.n544 B.n31 163.367
R468 B.n540 B.n31 163.367
R469 B.n540 B.n37 163.367
R470 B.n536 B.n37 163.367
R471 B.n536 B.n39 163.367
R472 B.n532 B.n39 163.367
R473 B.n532 B.n44 163.367
R474 B.n528 B.n44 163.367
R475 B.n528 B.n46 163.367
R476 B.n524 B.n46 163.367
R477 B.n524 B.n51 163.367
R478 B.n520 B.n51 163.367
R479 B.n520 B.n53 163.367
R480 B.n516 B.n53 163.367
R481 B.n516 B.n58 163.367
R482 B.n512 B.n58 163.367
R483 B.n512 B.n60 163.367
R484 B.n508 B.n60 163.367
R485 B.n268 B.n266 163.367
R486 B.n266 B.n265 163.367
R487 B.n262 B.n261 163.367
R488 B.n259 B.n162 163.367
R489 B.n255 B.n253 163.367
R490 B.n251 B.n164 163.367
R491 B.n247 B.n245 163.367
R492 B.n243 B.n166 163.367
R493 B.n239 B.n237 163.367
R494 B.n234 B.n233 163.367
R495 B.n231 B.n172 163.367
R496 B.n227 B.n225 163.367
R497 B.n223 B.n174 163.367
R498 B.n219 B.n217 163.367
R499 B.n214 B.n213 163.367
R500 B.n211 B.n180 163.367
R501 B.n207 B.n205 163.367
R502 B.n203 B.n182 163.367
R503 B.n199 B.n197 163.367
R504 B.n195 B.n184 163.367
R505 B.n191 B.n189 163.367
R506 B.n187 B.n156 163.367
R507 B.n274 B.n154 163.367
R508 B.n278 B.n154 163.367
R509 B.n278 B.n147 163.367
R510 B.n286 B.n147 163.367
R511 B.n286 B.n145 163.367
R512 B.n290 B.n145 163.367
R513 B.n290 B.n140 163.367
R514 B.n298 B.n140 163.367
R515 B.n298 B.n138 163.367
R516 B.n302 B.n138 163.367
R517 B.n302 B.n132 163.367
R518 B.n310 B.n132 163.367
R519 B.n310 B.n130 163.367
R520 B.n314 B.n130 163.367
R521 B.n314 B.n124 163.367
R522 B.n322 B.n124 163.367
R523 B.n322 B.n122 163.367
R524 B.n326 B.n122 163.367
R525 B.n326 B.n117 163.367
R526 B.n335 B.n117 163.367
R527 B.n335 B.n115 163.367
R528 B.n339 B.n115 163.367
R529 B.n339 B.n109 163.367
R530 B.n347 B.n109 163.367
R531 B.n347 B.n107 163.367
R532 B.n351 B.n107 163.367
R533 B.n351 B.n100 163.367
R534 B.n359 B.n100 163.367
R535 B.n359 B.n98 163.367
R536 B.n364 B.n98 163.367
R537 B.n364 B.n93 163.367
R538 B.n372 B.n93 163.367
R539 B.n373 B.n372 163.367
R540 B.n373 B.n5 163.367
R541 B.n6 B.n5 163.367
R542 B.n7 B.n6 163.367
R543 B.n378 B.n7 163.367
R544 B.n378 B.n12 163.367
R545 B.n13 B.n12 163.367
R546 B.n14 B.n13 163.367
R547 B.n383 B.n14 163.367
R548 B.n383 B.n19 163.367
R549 B.n20 B.n19 163.367
R550 B.n21 B.n20 163.367
R551 B.n388 B.n21 163.367
R552 B.n388 B.n26 163.367
R553 B.n27 B.n26 163.367
R554 B.n28 B.n27 163.367
R555 B.n393 B.n28 163.367
R556 B.n393 B.n33 163.367
R557 B.n34 B.n33 163.367
R558 B.n35 B.n34 163.367
R559 B.n398 B.n35 163.367
R560 B.n398 B.n40 163.367
R561 B.n41 B.n40 163.367
R562 B.n42 B.n41 163.367
R563 B.n403 B.n42 163.367
R564 B.n403 B.n47 163.367
R565 B.n48 B.n47 163.367
R566 B.n49 B.n48 163.367
R567 B.n408 B.n49 163.367
R568 B.n408 B.n54 163.367
R569 B.n55 B.n54 163.367
R570 B.n56 B.n55 163.367
R571 B.n413 B.n56 163.367
R572 B.n413 B.n61 163.367
R573 B.n62 B.n61 163.367
R574 B.n63 B.n62 163.367
R575 B.n504 B.n502 163.367
R576 B.n500 B.n67 163.367
R577 B.n496 B.n494 163.367
R578 B.n492 B.n69 163.367
R579 B.n488 B.n486 163.367
R580 B.n484 B.n71 163.367
R581 B.n480 B.n478 163.367
R582 B.n476 B.n73 163.367
R583 B.n471 B.n469 163.367
R584 B.n467 B.n77 163.367
R585 B.n463 B.n461 163.367
R586 B.n459 B.n79 163.367
R587 B.n455 B.n453 163.367
R588 B.n451 B.n81 163.367
R589 B.n447 B.n445 163.367
R590 B.n443 B.n86 163.367
R591 B.n439 B.n437 163.367
R592 B.n435 B.n88 163.367
R593 B.n431 B.n429 163.367
R594 B.n427 B.n90 163.367
R595 B.n423 B.n421 163.367
R596 B.n273 B.n157 163.008
R597 B.n509 B.n64 163.008
R598 B.n175 B.t21 112.459
R599 B.n82 B.t10 112.459
R600 B.n167 B.t15 112.456
R601 B.n74 B.t17 112.456
R602 B.n273 B.n153 83.3431
R603 B.n279 B.n153 83.3431
R604 B.n279 B.n148 83.3431
R605 B.n285 B.n148 83.3431
R606 B.n285 B.n149 83.3431
R607 B.n291 B.n141 83.3431
R608 B.n297 B.n141 83.3431
R609 B.n297 B.n137 83.3431
R610 B.n303 B.n137 83.3431
R611 B.n303 B.n133 83.3431
R612 B.n309 B.n133 83.3431
R613 B.n309 B.n129 83.3431
R614 B.n315 B.n129 83.3431
R615 B.n321 B.n125 83.3431
R616 B.n321 B.n121 83.3431
R617 B.n328 B.n121 83.3431
R618 B.n328 B.n327 83.3431
R619 B.n334 B.n114 83.3431
R620 B.n340 B.n114 83.3431
R621 B.n340 B.n110 83.3431
R622 B.n346 B.n110 83.3431
R623 B.n352 B.n106 83.3431
R624 B.n352 B.n101 83.3431
R625 B.n358 B.n101 83.3431
R626 B.n358 B.n102 83.3431
R627 B.n365 B.n94 83.3431
R628 B.n371 B.n94 83.3431
R629 B.n371 B.n4 83.3431
R630 B.n575 B.n4 83.3431
R631 B.n575 B.n574 83.3431
R632 B.n574 B.n573 83.3431
R633 B.n573 B.n8 83.3431
R634 B.n567 B.n8 83.3431
R635 B.n566 B.n565 83.3431
R636 B.n565 B.n15 83.3431
R637 B.n559 B.n15 83.3431
R638 B.n559 B.n558 83.3431
R639 B.n557 B.n22 83.3431
R640 B.n551 B.n22 83.3431
R641 B.n551 B.n550 83.3431
R642 B.n550 B.n549 83.3431
R643 B.n543 B.n32 83.3431
R644 B.n543 B.n542 83.3431
R645 B.n542 B.n541 83.3431
R646 B.n541 B.n36 83.3431
R647 B.n535 B.n534 83.3431
R648 B.n534 B.n533 83.3431
R649 B.n533 B.n43 83.3431
R650 B.n527 B.n43 83.3431
R651 B.n527 B.n526 83.3431
R652 B.n526 B.n525 83.3431
R653 B.n525 B.n50 83.3431
R654 B.n519 B.n50 83.3431
R655 B.n518 B.n517 83.3431
R656 B.n517 B.n57 83.3431
R657 B.n511 B.n57 83.3431
R658 B.n511 B.n510 83.3431
R659 B.n510 B.n509 83.3431
R660 B.n176 B.t20 78.1311
R661 B.n83 B.t11 78.1311
R662 B.n168 B.t14 78.1282
R663 B.n75 B.t18 78.1282
R664 B.n267 B.n158 71.676
R665 B.n265 B.n160 71.676
R666 B.n261 B.n260 71.676
R667 B.n254 B.n162 71.676
R668 B.n253 B.n252 71.676
R669 B.n246 B.n164 71.676
R670 B.n245 B.n244 71.676
R671 B.n238 B.n166 71.676
R672 B.n237 B.n170 71.676
R673 B.n233 B.n232 71.676
R674 B.n226 B.n172 71.676
R675 B.n225 B.n224 71.676
R676 B.n218 B.n174 71.676
R677 B.n217 B.n178 71.676
R678 B.n213 B.n212 71.676
R679 B.n206 B.n180 71.676
R680 B.n205 B.n204 71.676
R681 B.n198 B.n182 71.676
R682 B.n197 B.n196 71.676
R683 B.n190 B.n184 71.676
R684 B.n189 B.n188 71.676
R685 B.n503 B.n65 71.676
R686 B.n502 B.n501 71.676
R687 B.n495 B.n67 71.676
R688 B.n494 B.n493 71.676
R689 B.n487 B.n69 71.676
R690 B.n486 B.n485 71.676
R691 B.n479 B.n71 71.676
R692 B.n478 B.n477 71.676
R693 B.n470 B.n73 71.676
R694 B.n469 B.n468 71.676
R695 B.n462 B.n77 71.676
R696 B.n461 B.n460 71.676
R697 B.n454 B.n79 71.676
R698 B.n453 B.n452 71.676
R699 B.n446 B.n81 71.676
R700 B.n445 B.n444 71.676
R701 B.n438 B.n86 71.676
R702 B.n437 B.n436 71.676
R703 B.n430 B.n88 71.676
R704 B.n429 B.n428 71.676
R705 B.n422 B.n90 71.676
R706 B.n421 B.n420 71.676
R707 B.n420 B.n419 71.676
R708 B.n423 B.n422 71.676
R709 B.n428 B.n427 71.676
R710 B.n431 B.n430 71.676
R711 B.n436 B.n435 71.676
R712 B.n439 B.n438 71.676
R713 B.n444 B.n443 71.676
R714 B.n447 B.n446 71.676
R715 B.n452 B.n451 71.676
R716 B.n455 B.n454 71.676
R717 B.n460 B.n459 71.676
R718 B.n463 B.n462 71.676
R719 B.n468 B.n467 71.676
R720 B.n471 B.n470 71.676
R721 B.n477 B.n476 71.676
R722 B.n480 B.n479 71.676
R723 B.n485 B.n484 71.676
R724 B.n488 B.n487 71.676
R725 B.n493 B.n492 71.676
R726 B.n496 B.n495 71.676
R727 B.n501 B.n500 71.676
R728 B.n504 B.n503 71.676
R729 B.n268 B.n267 71.676
R730 B.n262 B.n160 71.676
R731 B.n260 B.n259 71.676
R732 B.n255 B.n254 71.676
R733 B.n252 B.n251 71.676
R734 B.n247 B.n246 71.676
R735 B.n244 B.n243 71.676
R736 B.n239 B.n238 71.676
R737 B.n234 B.n170 71.676
R738 B.n232 B.n231 71.676
R739 B.n227 B.n226 71.676
R740 B.n224 B.n223 71.676
R741 B.n219 B.n218 71.676
R742 B.n214 B.n178 71.676
R743 B.n212 B.n211 71.676
R744 B.n207 B.n206 71.676
R745 B.n204 B.n203 71.676
R746 B.n199 B.n198 71.676
R747 B.n196 B.n195 71.676
R748 B.n191 B.n190 71.676
R749 B.n188 B.n187 71.676
R750 B.t1 B.n125 68.6356
R751 B.t5 B.n36 68.6356
R752 B.n102 B.t6 66.1843
R753 B.t7 B.n566 66.1843
R754 B.n149 B.t13 63.7331
R755 B.t9 B.n518 63.7331
R756 B.n177 B.n176 59.5399
R757 B.n169 B.n168 59.5399
R758 B.n473 B.n75 59.5399
R759 B.n84 B.n83 59.5399
R760 B.n334 B.t4 51.4768
R761 B.n549 B.t3 51.4768
R762 B.n346 B.t2 49.0256
R763 B.t0 B.n557 49.0256
R764 B.n176 B.n175 34.3278
R765 B.n168 B.n167 34.3278
R766 B.n75 B.n74 34.3278
R767 B.n83 B.n82 34.3278
R768 B.t2 B.n106 34.318
R769 B.n558 B.t0 34.318
R770 B.n507 B.n506 33.8737
R771 B.n418 B.n417 33.8737
R772 B.n275 B.n155 33.8737
R773 B.n271 B.n270 33.8737
R774 B.n327 B.t4 31.8668
R775 B.n32 B.t3 31.8668
R776 B.n291 B.t13 19.6105
R777 B.n519 B.t9 19.6105
R778 B B.n577 18.0485
R779 B.n365 B.t6 17.1593
R780 B.n567 B.t7 17.1593
R781 B.n315 B.t1 14.708
R782 B.n535 B.t5 14.708
R783 B.n506 B.n505 10.6151
R784 B.n505 B.n66 10.6151
R785 B.n499 B.n66 10.6151
R786 B.n499 B.n498 10.6151
R787 B.n498 B.n497 10.6151
R788 B.n497 B.n68 10.6151
R789 B.n491 B.n68 10.6151
R790 B.n491 B.n490 10.6151
R791 B.n490 B.n489 10.6151
R792 B.n489 B.n70 10.6151
R793 B.n483 B.n70 10.6151
R794 B.n483 B.n482 10.6151
R795 B.n482 B.n481 10.6151
R796 B.n481 B.n72 10.6151
R797 B.n475 B.n72 10.6151
R798 B.n475 B.n474 10.6151
R799 B.n472 B.n76 10.6151
R800 B.n466 B.n76 10.6151
R801 B.n466 B.n465 10.6151
R802 B.n465 B.n464 10.6151
R803 B.n464 B.n78 10.6151
R804 B.n458 B.n78 10.6151
R805 B.n458 B.n457 10.6151
R806 B.n457 B.n456 10.6151
R807 B.n456 B.n80 10.6151
R808 B.n450 B.n449 10.6151
R809 B.n449 B.n448 10.6151
R810 B.n448 B.n85 10.6151
R811 B.n442 B.n85 10.6151
R812 B.n442 B.n441 10.6151
R813 B.n441 B.n440 10.6151
R814 B.n440 B.n87 10.6151
R815 B.n434 B.n87 10.6151
R816 B.n434 B.n433 10.6151
R817 B.n433 B.n432 10.6151
R818 B.n432 B.n89 10.6151
R819 B.n426 B.n89 10.6151
R820 B.n426 B.n425 10.6151
R821 B.n425 B.n424 10.6151
R822 B.n424 B.n91 10.6151
R823 B.n418 B.n91 10.6151
R824 B.n276 B.n275 10.6151
R825 B.n277 B.n276 10.6151
R826 B.n277 B.n146 10.6151
R827 B.n287 B.n146 10.6151
R828 B.n288 B.n287 10.6151
R829 B.n289 B.n288 10.6151
R830 B.n289 B.n139 10.6151
R831 B.n299 B.n139 10.6151
R832 B.n300 B.n299 10.6151
R833 B.n301 B.n300 10.6151
R834 B.n301 B.n131 10.6151
R835 B.n311 B.n131 10.6151
R836 B.n312 B.n311 10.6151
R837 B.n313 B.n312 10.6151
R838 B.n313 B.n123 10.6151
R839 B.n323 B.n123 10.6151
R840 B.n324 B.n323 10.6151
R841 B.n325 B.n324 10.6151
R842 B.n325 B.n116 10.6151
R843 B.n336 B.n116 10.6151
R844 B.n337 B.n336 10.6151
R845 B.n338 B.n337 10.6151
R846 B.n338 B.n108 10.6151
R847 B.n348 B.n108 10.6151
R848 B.n349 B.n348 10.6151
R849 B.n350 B.n349 10.6151
R850 B.n350 B.n99 10.6151
R851 B.n360 B.n99 10.6151
R852 B.n361 B.n360 10.6151
R853 B.n363 B.n361 10.6151
R854 B.n363 B.n362 10.6151
R855 B.n362 B.n92 10.6151
R856 B.n374 B.n92 10.6151
R857 B.n375 B.n374 10.6151
R858 B.n376 B.n375 10.6151
R859 B.n377 B.n376 10.6151
R860 B.n379 B.n377 10.6151
R861 B.n380 B.n379 10.6151
R862 B.n381 B.n380 10.6151
R863 B.n382 B.n381 10.6151
R864 B.n384 B.n382 10.6151
R865 B.n385 B.n384 10.6151
R866 B.n386 B.n385 10.6151
R867 B.n387 B.n386 10.6151
R868 B.n389 B.n387 10.6151
R869 B.n390 B.n389 10.6151
R870 B.n391 B.n390 10.6151
R871 B.n392 B.n391 10.6151
R872 B.n394 B.n392 10.6151
R873 B.n395 B.n394 10.6151
R874 B.n396 B.n395 10.6151
R875 B.n397 B.n396 10.6151
R876 B.n399 B.n397 10.6151
R877 B.n400 B.n399 10.6151
R878 B.n401 B.n400 10.6151
R879 B.n402 B.n401 10.6151
R880 B.n404 B.n402 10.6151
R881 B.n405 B.n404 10.6151
R882 B.n406 B.n405 10.6151
R883 B.n407 B.n406 10.6151
R884 B.n409 B.n407 10.6151
R885 B.n410 B.n409 10.6151
R886 B.n411 B.n410 10.6151
R887 B.n412 B.n411 10.6151
R888 B.n414 B.n412 10.6151
R889 B.n415 B.n414 10.6151
R890 B.n416 B.n415 10.6151
R891 B.n417 B.n416 10.6151
R892 B.n270 B.n269 10.6151
R893 B.n269 B.n159 10.6151
R894 B.n264 B.n159 10.6151
R895 B.n264 B.n263 10.6151
R896 B.n263 B.n161 10.6151
R897 B.n258 B.n161 10.6151
R898 B.n258 B.n257 10.6151
R899 B.n257 B.n256 10.6151
R900 B.n256 B.n163 10.6151
R901 B.n250 B.n163 10.6151
R902 B.n250 B.n249 10.6151
R903 B.n249 B.n248 10.6151
R904 B.n248 B.n165 10.6151
R905 B.n242 B.n165 10.6151
R906 B.n242 B.n241 10.6151
R907 B.n241 B.n240 10.6151
R908 B.n236 B.n235 10.6151
R909 B.n235 B.n171 10.6151
R910 B.n230 B.n171 10.6151
R911 B.n230 B.n229 10.6151
R912 B.n229 B.n228 10.6151
R913 B.n228 B.n173 10.6151
R914 B.n222 B.n173 10.6151
R915 B.n222 B.n221 10.6151
R916 B.n221 B.n220 10.6151
R917 B.n216 B.n215 10.6151
R918 B.n215 B.n179 10.6151
R919 B.n210 B.n179 10.6151
R920 B.n210 B.n209 10.6151
R921 B.n209 B.n208 10.6151
R922 B.n208 B.n181 10.6151
R923 B.n202 B.n181 10.6151
R924 B.n202 B.n201 10.6151
R925 B.n201 B.n200 10.6151
R926 B.n200 B.n183 10.6151
R927 B.n194 B.n183 10.6151
R928 B.n194 B.n193 10.6151
R929 B.n193 B.n192 10.6151
R930 B.n192 B.n185 10.6151
R931 B.n186 B.n185 10.6151
R932 B.n186 B.n155 10.6151
R933 B.n271 B.n151 10.6151
R934 B.n281 B.n151 10.6151
R935 B.n282 B.n281 10.6151
R936 B.n283 B.n282 10.6151
R937 B.n283 B.n143 10.6151
R938 B.n293 B.n143 10.6151
R939 B.n294 B.n293 10.6151
R940 B.n295 B.n294 10.6151
R941 B.n295 B.n135 10.6151
R942 B.n305 B.n135 10.6151
R943 B.n306 B.n305 10.6151
R944 B.n307 B.n306 10.6151
R945 B.n307 B.n127 10.6151
R946 B.n317 B.n127 10.6151
R947 B.n318 B.n317 10.6151
R948 B.n319 B.n318 10.6151
R949 B.n319 B.n119 10.6151
R950 B.n330 B.n119 10.6151
R951 B.n331 B.n330 10.6151
R952 B.n332 B.n331 10.6151
R953 B.n332 B.n112 10.6151
R954 B.n342 B.n112 10.6151
R955 B.n343 B.n342 10.6151
R956 B.n344 B.n343 10.6151
R957 B.n344 B.n104 10.6151
R958 B.n354 B.n104 10.6151
R959 B.n355 B.n354 10.6151
R960 B.n356 B.n355 10.6151
R961 B.n356 B.n96 10.6151
R962 B.n367 B.n96 10.6151
R963 B.n368 B.n367 10.6151
R964 B.n369 B.n368 10.6151
R965 B.n369 B.n0 10.6151
R966 B.n571 B.n1 10.6151
R967 B.n571 B.n570 10.6151
R968 B.n570 B.n569 10.6151
R969 B.n569 B.n10 10.6151
R970 B.n563 B.n10 10.6151
R971 B.n563 B.n562 10.6151
R972 B.n562 B.n561 10.6151
R973 B.n561 B.n17 10.6151
R974 B.n555 B.n17 10.6151
R975 B.n555 B.n554 10.6151
R976 B.n554 B.n553 10.6151
R977 B.n553 B.n24 10.6151
R978 B.n547 B.n24 10.6151
R979 B.n547 B.n546 10.6151
R980 B.n546 B.n545 10.6151
R981 B.n545 B.n30 10.6151
R982 B.n539 B.n30 10.6151
R983 B.n539 B.n538 10.6151
R984 B.n538 B.n537 10.6151
R985 B.n537 B.n38 10.6151
R986 B.n531 B.n38 10.6151
R987 B.n531 B.n530 10.6151
R988 B.n530 B.n529 10.6151
R989 B.n529 B.n45 10.6151
R990 B.n523 B.n45 10.6151
R991 B.n523 B.n522 10.6151
R992 B.n522 B.n521 10.6151
R993 B.n521 B.n52 10.6151
R994 B.n515 B.n52 10.6151
R995 B.n515 B.n514 10.6151
R996 B.n514 B.n513 10.6151
R997 B.n513 B.n59 10.6151
R998 B.n507 B.n59 10.6151
R999 B.n474 B.n473 9.36635
R1000 B.n450 B.n84 9.36635
R1001 B.n240 B.n169 9.36635
R1002 B.n216 B.n177 9.36635
R1003 B.n577 B.n0 2.81026
R1004 B.n577 B.n1 2.81026
R1005 B.n473 B.n472 1.24928
R1006 B.n84 B.n80 1.24928
R1007 B.n236 B.n169 1.24928
R1008 B.n220 B.n177 1.24928
R1009 VP.n26 VP.n25 178.268
R1010 VP.n46 VP.n45 178.268
R1011 VP.n24 VP.n23 178.268
R1012 VP.n12 VP.n9 161.3
R1013 VP.n14 VP.n13 161.3
R1014 VP.n15 VP.n8 161.3
R1015 VP.n18 VP.n17 161.3
R1016 VP.n19 VP.n7 161.3
R1017 VP.n21 VP.n20 161.3
R1018 VP.n22 VP.n6 161.3
R1019 VP.n44 VP.n0 161.3
R1020 VP.n43 VP.n42 161.3
R1021 VP.n41 VP.n1 161.3
R1022 VP.n40 VP.n39 161.3
R1023 VP.n37 VP.n2 161.3
R1024 VP.n36 VP.n35 161.3
R1025 VP.n34 VP.n3 161.3
R1026 VP.n33 VP.n32 161.3
R1027 VP.n30 VP.n4 161.3
R1028 VP.n29 VP.n28 161.3
R1029 VP.n27 VP.n5 161.3
R1030 VP.n11 VP.t3 94.4546
R1031 VP.n25 VP.t6 61.9241
R1032 VP.n31 VP.t2 61.9241
R1033 VP.n38 VP.t7 61.9241
R1034 VP.n45 VP.t4 61.9241
R1035 VP.n23 VP.t1 61.9241
R1036 VP.n16 VP.t5 61.9241
R1037 VP.n10 VP.t0 61.9241
R1038 VP.n30 VP.n29 56.5617
R1039 VP.n43 VP.n1 56.5617
R1040 VP.n21 VP.n7 56.5617
R1041 VP.n11 VP.n10 47.4091
R1042 VP.n36 VP.n3 40.577
R1043 VP.n37 VP.n36 40.577
R1044 VP.n15 VP.n14 40.577
R1045 VP.n14 VP.n9 40.577
R1046 VP.n26 VP.n24 39.0535
R1047 VP.n29 VP.n5 24.5923
R1048 VP.n32 VP.n30 24.5923
R1049 VP.n39 VP.n1 24.5923
R1050 VP.n44 VP.n43 24.5923
R1051 VP.n22 VP.n21 24.5923
R1052 VP.n17 VP.n7 24.5923
R1053 VP.n31 VP.n3 18.9362
R1054 VP.n38 VP.n37 18.9362
R1055 VP.n16 VP.n15 18.9362
R1056 VP.n10 VP.n9 18.9362
R1057 VP.n12 VP.n11 17.9988
R1058 VP.n25 VP.n5 7.62397
R1059 VP.n45 VP.n44 7.62397
R1060 VP.n23 VP.n22 7.62397
R1061 VP.n32 VP.n31 5.65662
R1062 VP.n39 VP.n38 5.65662
R1063 VP.n17 VP.n16 5.65662
R1064 VP.n13 VP.n12 0.189894
R1065 VP.n13 VP.n8 0.189894
R1066 VP.n18 VP.n8 0.189894
R1067 VP.n19 VP.n18 0.189894
R1068 VP.n20 VP.n19 0.189894
R1069 VP.n20 VP.n6 0.189894
R1070 VP.n24 VP.n6 0.189894
R1071 VP.n27 VP.n26 0.189894
R1072 VP.n28 VP.n27 0.189894
R1073 VP.n28 VP.n4 0.189894
R1074 VP.n33 VP.n4 0.189894
R1075 VP.n34 VP.n33 0.189894
R1076 VP.n35 VP.n34 0.189894
R1077 VP.n35 VP.n2 0.189894
R1078 VP.n40 VP.n2 0.189894
R1079 VP.n41 VP.n40 0.189894
R1080 VP.n42 VP.n41 0.189894
R1081 VP.n42 VP.n0 0.189894
R1082 VP.n46 VP.n0 0.189894
R1083 VP VP.n46 0.0516364
R1084 VTAIL.n11 VTAIL.t12 68.2998
R1085 VTAIL.n10 VTAIL.t6 68.2998
R1086 VTAIL.n7 VTAIL.t1 68.2998
R1087 VTAIL.n15 VTAIL.t5 68.2997
R1088 VTAIL.n2 VTAIL.t7 68.2997
R1089 VTAIL.n3 VTAIL.t10 68.2997
R1090 VTAIL.n6 VTAIL.t14 68.2997
R1091 VTAIL.n14 VTAIL.t9 68.2997
R1092 VTAIL.n13 VTAIL.n12 62.9485
R1093 VTAIL.n9 VTAIL.n8 62.9485
R1094 VTAIL.n1 VTAIL.n0 62.9483
R1095 VTAIL.n5 VTAIL.n4 62.9483
R1096 VTAIL.n15 VTAIL.n14 17.0824
R1097 VTAIL.n7 VTAIL.n6 17.0824
R1098 VTAIL.n0 VTAIL.t0 5.35185
R1099 VTAIL.n0 VTAIL.t3 5.35185
R1100 VTAIL.n4 VTAIL.t8 5.35185
R1101 VTAIL.n4 VTAIL.t15 5.35185
R1102 VTAIL.n12 VTAIL.t11 5.35185
R1103 VTAIL.n12 VTAIL.t13 5.35185
R1104 VTAIL.n8 VTAIL.t4 5.35185
R1105 VTAIL.n8 VTAIL.t2 5.35185
R1106 VTAIL.n9 VTAIL.n7 1.52636
R1107 VTAIL.n10 VTAIL.n9 1.52636
R1108 VTAIL.n13 VTAIL.n11 1.52636
R1109 VTAIL.n14 VTAIL.n13 1.52636
R1110 VTAIL.n6 VTAIL.n5 1.52636
R1111 VTAIL.n5 VTAIL.n3 1.52636
R1112 VTAIL.n2 VTAIL.n1 1.52636
R1113 VTAIL VTAIL.n15 1.46817
R1114 VTAIL.n11 VTAIL.n10 0.470328
R1115 VTAIL.n3 VTAIL.n2 0.470328
R1116 VTAIL VTAIL.n1 0.0586897
R1117 VDD1 VDD1.n0 80.4484
R1118 VDD1.n3 VDD1.n2 80.3347
R1119 VDD1.n3 VDD1.n1 80.3347
R1120 VDD1.n5 VDD1.n4 79.6272
R1121 VDD1.n5 VDD1.n3 34.3543
R1122 VDD1.n4 VDD1.t2 5.35185
R1123 VDD1.n4 VDD1.t6 5.35185
R1124 VDD1.n0 VDD1.t4 5.35185
R1125 VDD1.n0 VDD1.t7 5.35185
R1126 VDD1.n2 VDD1.t0 5.35185
R1127 VDD1.n2 VDD1.t3 5.35185
R1128 VDD1.n1 VDD1.t1 5.35185
R1129 VDD1.n1 VDD1.t5 5.35185
R1130 VDD1 VDD1.n5 0.705241
R1131 VN.n18 VN.n17 178.268
R1132 VN.n37 VN.n36 178.268
R1133 VN.n35 VN.n19 161.3
R1134 VN.n34 VN.n33 161.3
R1135 VN.n32 VN.n20 161.3
R1136 VN.n31 VN.n30 161.3
R1137 VN.n28 VN.n21 161.3
R1138 VN.n27 VN.n26 161.3
R1139 VN.n25 VN.n22 161.3
R1140 VN.n16 VN.n0 161.3
R1141 VN.n15 VN.n14 161.3
R1142 VN.n13 VN.n1 161.3
R1143 VN.n12 VN.n11 161.3
R1144 VN.n9 VN.n2 161.3
R1145 VN.n8 VN.n7 161.3
R1146 VN.n6 VN.n3 161.3
R1147 VN.n5 VN.t4 94.4546
R1148 VN.n24 VN.t3 94.4546
R1149 VN.n4 VN.t5 61.9241
R1150 VN.n10 VN.t1 61.9241
R1151 VN.n17 VN.t2 61.9241
R1152 VN.n23 VN.t0 61.9241
R1153 VN.n29 VN.t7 61.9241
R1154 VN.n36 VN.t6 61.9241
R1155 VN.n15 VN.n1 56.5617
R1156 VN.n34 VN.n20 56.5617
R1157 VN.n5 VN.n4 47.4091
R1158 VN.n24 VN.n23 47.4091
R1159 VN.n8 VN.n3 40.577
R1160 VN.n9 VN.n8 40.577
R1161 VN.n27 VN.n22 40.577
R1162 VN.n28 VN.n27 40.577
R1163 VN VN.n37 39.4342
R1164 VN.n11 VN.n1 24.5923
R1165 VN.n16 VN.n15 24.5923
R1166 VN.n30 VN.n20 24.5923
R1167 VN.n35 VN.n34 24.5923
R1168 VN.n4 VN.n3 18.9362
R1169 VN.n10 VN.n9 18.9362
R1170 VN.n23 VN.n22 18.9362
R1171 VN.n29 VN.n28 18.9362
R1172 VN.n25 VN.n24 17.9988
R1173 VN.n6 VN.n5 17.9988
R1174 VN.n17 VN.n16 7.62397
R1175 VN.n36 VN.n35 7.62397
R1176 VN.n11 VN.n10 5.65662
R1177 VN.n30 VN.n29 5.65662
R1178 VN.n37 VN.n19 0.189894
R1179 VN.n33 VN.n19 0.189894
R1180 VN.n33 VN.n32 0.189894
R1181 VN.n32 VN.n31 0.189894
R1182 VN.n31 VN.n21 0.189894
R1183 VN.n26 VN.n21 0.189894
R1184 VN.n26 VN.n25 0.189894
R1185 VN.n7 VN.n6 0.189894
R1186 VN.n7 VN.n2 0.189894
R1187 VN.n12 VN.n2 0.189894
R1188 VN.n13 VN.n12 0.189894
R1189 VN.n14 VN.n13 0.189894
R1190 VN.n14 VN.n0 0.189894
R1191 VN.n18 VN.n0 0.189894
R1192 VN VN.n18 0.0516364
R1193 VDD2.n2 VDD2.n1 80.3347
R1194 VDD2.n2 VDD2.n0 80.3347
R1195 VDD2 VDD2.n5 80.3319
R1196 VDD2.n4 VDD2.n3 79.6273
R1197 VDD2.n4 VDD2.n2 33.7713
R1198 VDD2.n5 VDD2.t7 5.35185
R1199 VDD2.n5 VDD2.t4 5.35185
R1200 VDD2.n3 VDD2.t1 5.35185
R1201 VDD2.n3 VDD2.t0 5.35185
R1202 VDD2.n1 VDD2.t6 5.35185
R1203 VDD2.n1 VDD2.t5 5.35185
R1204 VDD2.n0 VDD2.t3 5.35185
R1205 VDD2.n0 VDD2.t2 5.35185
R1206 VDD2 VDD2.n4 0.821621
C0 VP VTAIL 3.09966f
C1 VN VP 4.71086f
C2 VN VTAIL 3.08556f
C3 VDD1 VDD2 1.1989f
C4 VP VDD2 0.401636f
C5 VTAIL VDD2 4.65806f
C6 VN VDD2 2.58824f
C7 VDD1 VP 2.83397f
C8 VDD1 VTAIL 4.61142f
C9 VDD1 VN 0.154521f
C10 VDD2 B 3.54241f
C11 VDD1 B 3.852508f
C12 VTAIL B 4.501195f
C13 VN B 10.263741f
C14 VP B 8.799721f
C15 VDD2.t3 B 0.072858f
C16 VDD2.t2 B 0.072858f
C17 VDD2.n0 B 0.566442f
C18 VDD2.t6 B 0.072858f
C19 VDD2.t5 B 0.072858f
C20 VDD2.n1 B 0.566442f
C21 VDD2.n2 B 2.07702f
C22 VDD2.t1 B 0.072858f
C23 VDD2.t0 B 0.072858f
C24 VDD2.n3 B 0.563063f
C25 VDD2.n4 B 1.87585f
C26 VDD2.t7 B 0.072858f
C27 VDD2.t4 B 0.072858f
C28 VDD2.n5 B 0.566418f
C29 VN.n0 B 0.035461f
C30 VN.t2 B 0.481791f
C31 VN.n1 B 0.053511f
C32 VN.n2 B 0.035461f
C33 VN.t1 B 0.481791f
C34 VN.n3 B 0.062641f
C35 VN.t4 B 0.598826f
C36 VN.t5 B 0.481791f
C37 VN.n4 B 0.28141f
C38 VN.n5 B 0.275481f
C39 VN.n6 B 0.221379f
C40 VN.n7 B 0.035461f
C41 VN.n8 B 0.028641f
C42 VN.n9 B 0.062641f
C43 VN.n10 B 0.208962f
C44 VN.n11 B 0.040763f
C45 VN.n12 B 0.035461f
C46 VN.n13 B 0.035461f
C47 VN.n14 B 0.035461f
C48 VN.n15 B 0.049586f
C49 VN.n16 B 0.04336f
C50 VN.n17 B 0.274043f
C51 VN.n18 B 0.034328f
C52 VN.n19 B 0.035461f
C53 VN.t6 B 0.481791f
C54 VN.n20 B 0.053511f
C55 VN.n21 B 0.035461f
C56 VN.t7 B 0.481791f
C57 VN.n22 B 0.062641f
C58 VN.t3 B 0.598826f
C59 VN.t0 B 0.481791f
C60 VN.n23 B 0.28141f
C61 VN.n24 B 0.275481f
C62 VN.n25 B 0.221379f
C63 VN.n26 B 0.035461f
C64 VN.n27 B 0.028641f
C65 VN.n28 B 0.062641f
C66 VN.n29 B 0.208962f
C67 VN.n30 B 0.040763f
C68 VN.n31 B 0.035461f
C69 VN.n32 B 0.035461f
C70 VN.n33 B 0.035461f
C71 VN.n34 B 0.049586f
C72 VN.n35 B 0.04336f
C73 VN.n36 B 0.274043f
C74 VN.n37 B 1.32271f
C75 VDD1.t4 B 0.072937f
C76 VDD1.t7 B 0.072937f
C77 VDD1.n0 B 0.567676f
C78 VDD1.t1 B 0.072937f
C79 VDD1.t5 B 0.072937f
C80 VDD1.n1 B 0.567052f
C81 VDD1.t0 B 0.072937f
C82 VDD1.t3 B 0.072937f
C83 VDD1.n2 B 0.567052f
C84 VDD1.n3 B 2.13217f
C85 VDD1.t2 B 0.072937f
C86 VDD1.t6 B 0.072937f
C87 VDD1.n4 B 0.563667f
C88 VDD1.n5 B 1.90774f
C89 VTAIL.t0 B 0.071359f
C90 VTAIL.t3 B 0.071359f
C91 VTAIL.n0 B 0.502465f
C92 VTAIL.n1 B 0.330028f
C93 VTAIL.t7 B 0.648053f
C94 VTAIL.n2 B 0.411426f
C95 VTAIL.t10 B 0.648053f
C96 VTAIL.n3 B 0.411426f
C97 VTAIL.t8 B 0.071359f
C98 VTAIL.t15 B 0.071359f
C99 VTAIL.n4 B 0.502465f
C100 VTAIL.n5 B 0.445447f
C101 VTAIL.t14 B 0.648053f
C102 VTAIL.n6 B 1.07684f
C103 VTAIL.t1 B 0.648057f
C104 VTAIL.n7 B 1.07683f
C105 VTAIL.t4 B 0.071359f
C106 VTAIL.t2 B 0.071359f
C107 VTAIL.n8 B 0.502467f
C108 VTAIL.n9 B 0.445445f
C109 VTAIL.t6 B 0.648057f
C110 VTAIL.n10 B 0.411423f
C111 VTAIL.t12 B 0.648057f
C112 VTAIL.n11 B 0.411423f
C113 VTAIL.t11 B 0.071359f
C114 VTAIL.t13 B 0.071359f
C115 VTAIL.n12 B 0.502467f
C116 VTAIL.n13 B 0.445445f
C117 VTAIL.t9 B 0.648053f
C118 VTAIL.n14 B 1.07684f
C119 VTAIL.t5 B 0.648053f
C120 VTAIL.n15 B 1.07226f
C121 VP.n0 B 0.036317f
C122 VP.t4 B 0.493421f
C123 VP.n1 B 0.054803f
C124 VP.n2 B 0.036317f
C125 VP.t7 B 0.493421f
C126 VP.n3 B 0.064153f
C127 VP.n4 B 0.036317f
C128 VP.n5 B 0.044406f
C129 VP.n6 B 0.036317f
C130 VP.t1 B 0.493421f
C131 VP.n7 B 0.054803f
C132 VP.n8 B 0.036317f
C133 VP.t5 B 0.493421f
C134 VP.n9 B 0.064153f
C135 VP.t3 B 0.613281f
C136 VP.t0 B 0.493421f
C137 VP.n10 B 0.288203f
C138 VP.n11 B 0.282132f
C139 VP.n12 B 0.226723f
C140 VP.n13 B 0.036317f
C141 VP.n14 B 0.029332f
C142 VP.n15 B 0.064153f
C143 VP.n16 B 0.214006f
C144 VP.n17 B 0.041747f
C145 VP.n18 B 0.036317f
C146 VP.n19 B 0.036317f
C147 VP.n20 B 0.036317f
C148 VP.n21 B 0.050783f
C149 VP.n22 B 0.044406f
C150 VP.n23 B 0.280659f
C151 VP.n24 B 1.33069f
C152 VP.t6 B 0.493421f
C153 VP.n25 B 0.280659f
C154 VP.n26 B 1.36421f
C155 VP.n27 B 0.036317f
C156 VP.n28 B 0.036317f
C157 VP.n29 B 0.050783f
C158 VP.n30 B 0.054803f
C159 VP.t2 B 0.493421f
C160 VP.n31 B 0.214006f
C161 VP.n32 B 0.041747f
C162 VP.n33 B 0.036317f
C163 VP.n34 B 0.036317f
C164 VP.n35 B 0.036317f
C165 VP.n36 B 0.029332f
C166 VP.n37 B 0.064153f
C167 VP.n38 B 0.214006f
C168 VP.n39 B 0.041747f
C169 VP.n40 B 0.036317f
C170 VP.n41 B 0.036317f
C171 VP.n42 B 0.036317f
C172 VP.n43 B 0.050783f
C173 VP.n44 B 0.044406f
C174 VP.n45 B 0.280659f
C175 VP.n46 B 0.035156f
.ends

