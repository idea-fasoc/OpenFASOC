* NGSPICE file created from diff_pair_sample_1666.ext - technology: sky130A

.subckt diff_pair_sample_1666 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=4.5708 pd=24.22 as=1.9338 ps=12.05 w=11.72 l=0.78
X1 VDD2.t9 VN.t0 VTAIL.t19 B.t9 sky130_fd_pr__nfet_01v8 ad=1.9338 pd=12.05 as=1.9338 ps=12.05 w=11.72 l=0.78
X2 VDD2.t8 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.9338 pd=12.05 as=1.9338 ps=12.05 w=11.72 l=0.78
X3 VTAIL.t12 VP.t1 VDD1.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9338 pd=12.05 as=1.9338 ps=12.05 w=11.72 l=0.78
X4 VDD1.t7 VP.t2 VTAIL.t14 B.t5 sky130_fd_pr__nfet_01v8 ad=1.9338 pd=12.05 as=4.5708 ps=24.22 w=11.72 l=0.78
X5 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=4.5708 pd=24.22 as=0 ps=0 w=11.72 l=0.78
X6 VDD1.t6 VP.t3 VTAIL.t16 B.t0 sky130_fd_pr__nfet_01v8 ad=4.5708 pd=24.22 as=1.9338 ps=12.05 w=11.72 l=0.78
X7 VDD1.t5 VP.t4 VTAIL.t13 B.t8 sky130_fd_pr__nfet_01v8 ad=1.9338 pd=12.05 as=4.5708 ps=24.22 w=11.72 l=0.78
X8 VTAIL.t17 VP.t5 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=1.9338 pd=12.05 as=1.9338 ps=12.05 w=11.72 l=0.78
X9 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=4.5708 pd=24.22 as=0 ps=0 w=11.72 l=0.78
X10 VDD2.t7 VN.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.9338 pd=12.05 as=4.5708 ps=24.22 w=11.72 l=0.78
X11 VDD2.t6 VN.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=4.5708 pd=24.22 as=1.9338 ps=12.05 w=11.72 l=0.78
X12 VTAIL.t7 VN.t4 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=1.9338 pd=12.05 as=1.9338 ps=12.05 w=11.72 l=0.78
X13 VDD2.t4 VN.t5 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=1.9338 pd=12.05 as=4.5708 ps=24.22 w=11.72 l=0.78
X14 VTAIL.t3 VN.t6 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9338 pd=12.05 as=1.9338 ps=12.05 w=11.72 l=0.78
X15 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=4.5708 pd=24.22 as=0 ps=0 w=11.72 l=0.78
X16 VDD1.t3 VP.t6 VTAIL.t18 B.t2 sky130_fd_pr__nfet_01v8 ad=1.9338 pd=12.05 as=1.9338 ps=12.05 w=11.72 l=0.78
X17 VTAIL.t1 VN.t7 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9338 pd=12.05 as=1.9338 ps=12.05 w=11.72 l=0.78
X18 VDD1.t2 VP.t7 VTAIL.t11 B.t9 sky130_fd_pr__nfet_01v8 ad=1.9338 pd=12.05 as=1.9338 ps=12.05 w=11.72 l=0.78
X19 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.5708 pd=24.22 as=0 ps=0 w=11.72 l=0.78
X20 VTAIL.t4 VN.t8 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9338 pd=12.05 as=1.9338 ps=12.05 w=11.72 l=0.78
X21 VTAIL.t9 VP.t8 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9338 pd=12.05 as=1.9338 ps=12.05 w=11.72 l=0.78
X22 VDD2.t0 VN.t9 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.5708 pd=24.22 as=1.9338 ps=12.05 w=11.72 l=0.78
X23 VTAIL.t15 VP.t9 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9338 pd=12.05 as=1.9338 ps=12.05 w=11.72 l=0.78
R0 VP.n6 VP.t0 435.139
R1 VP.n14 VP.t3 413.099
R2 VP.n16 VP.t8 413.099
R3 VP.n1 VP.t7 413.099
R4 VP.n20 VP.t1 413.099
R5 VP.n22 VP.t4 413.099
R6 VP.n11 VP.t2 413.099
R7 VP.n9 VP.t9 413.099
R8 VP.n8 VP.t6 413.099
R9 VP.n7 VP.t5 413.099
R10 VP.n23 VP.n22 161.3
R11 VP.n10 VP.n3 161.3
R12 VP.n12 VP.n11 161.3
R13 VP.n21 VP.n0 161.3
R14 VP.n15 VP.n2 161.3
R15 VP.n14 VP.n13 161.3
R16 VP.n8 VP.n5 80.6037
R17 VP.n9 VP.n4 80.6037
R18 VP.n20 VP.n19 80.6037
R19 VP.n18 VP.n1 80.6037
R20 VP.n17 VP.n16 80.6037
R21 VP.n16 VP.n1 48.2005
R22 VP.n20 VP.n1 48.2005
R23 VP.n9 VP.n8 48.2005
R24 VP.n8 VP.n7 48.2005
R25 VP.n13 VP.n12 42.9588
R26 VP.n16 VP.n15 36.5157
R27 VP.n21 VP.n20 36.5157
R28 VP.n10 VP.n9 36.5157
R29 VP.n6 VP.n5 31.7379
R30 VP.n7 VP.n6 16.9109
R31 VP.n15 VP.n14 11.6853
R32 VP.n22 VP.n21 11.6853
R33 VP.n11 VP.n10 11.6853
R34 VP.n5 VP.n4 0.380177
R35 VP.n18 VP.n17 0.380177
R36 VP.n19 VP.n18 0.380177
R37 VP.n4 VP.n3 0.285035
R38 VP.n17 VP.n2 0.285035
R39 VP.n19 VP.n0 0.285035
R40 VP.n12 VP.n3 0.189894
R41 VP.n13 VP.n2 0.189894
R42 VP.n23 VP.n0 0.189894
R43 VP VP.n23 0.0516364
R44 VTAIL.n11 VTAIL.t8 46.2149
R45 VTAIL.n17 VTAIL.t5 46.2147
R46 VTAIL.n2 VTAIL.t13 46.2147
R47 VTAIL.n16 VTAIL.t14 46.2147
R48 VTAIL.n15 VTAIL.n14 44.5255
R49 VTAIL.n13 VTAIL.n12 44.5255
R50 VTAIL.n10 VTAIL.n9 44.5255
R51 VTAIL.n8 VTAIL.n7 44.5255
R52 VTAIL.n19 VTAIL.n18 44.5252
R53 VTAIL.n1 VTAIL.n0 44.5252
R54 VTAIL.n4 VTAIL.n3 44.5252
R55 VTAIL.n6 VTAIL.n5 44.5252
R56 VTAIL.n8 VTAIL.n6 24.3841
R57 VTAIL.n17 VTAIL.n16 23.4272
R58 VTAIL.n18 VTAIL.t2 1.68992
R59 VTAIL.n18 VTAIL.t1 1.68992
R60 VTAIL.n0 VTAIL.t6 1.68992
R61 VTAIL.n0 VTAIL.t7 1.68992
R62 VTAIL.n3 VTAIL.t11 1.68992
R63 VTAIL.n3 VTAIL.t12 1.68992
R64 VTAIL.n5 VTAIL.t16 1.68992
R65 VTAIL.n5 VTAIL.t9 1.68992
R66 VTAIL.n14 VTAIL.t18 1.68992
R67 VTAIL.n14 VTAIL.t15 1.68992
R68 VTAIL.n12 VTAIL.t10 1.68992
R69 VTAIL.n12 VTAIL.t17 1.68992
R70 VTAIL.n9 VTAIL.t19 1.68992
R71 VTAIL.n9 VTAIL.t4 1.68992
R72 VTAIL.n7 VTAIL.t0 1.68992
R73 VTAIL.n7 VTAIL.t3 1.68992
R74 VTAIL.n10 VTAIL.n8 0.957397
R75 VTAIL.n11 VTAIL.n10 0.957397
R76 VTAIL.n15 VTAIL.n13 0.957397
R77 VTAIL.n16 VTAIL.n15 0.957397
R78 VTAIL.n6 VTAIL.n4 0.957397
R79 VTAIL.n4 VTAIL.n2 0.957397
R80 VTAIL.n19 VTAIL.n17 0.957397
R81 VTAIL.n13 VTAIL.n11 0.948776
R82 VTAIL.n2 VTAIL.n1 0.948776
R83 VTAIL VTAIL.n1 0.776362
R84 VTAIL VTAIL.n19 0.181534
R85 VDD1.n1 VDD1.t9 63.8506
R86 VDD1.n3 VDD1.t6 63.8504
R87 VDD1.n5 VDD1.n4 61.8664
R88 VDD1.n1 VDD1.n0 61.2043
R89 VDD1.n7 VDD1.n6 61.2041
R90 VDD1.n3 VDD1.n2 61.204
R91 VDD1.n7 VDD1.n5 39.4255
R92 VDD1.n6 VDD1.t0 1.68992
R93 VDD1.n6 VDD1.t7 1.68992
R94 VDD1.n0 VDD1.t4 1.68992
R95 VDD1.n0 VDD1.t3 1.68992
R96 VDD1.n4 VDD1.t8 1.68992
R97 VDD1.n4 VDD1.t5 1.68992
R98 VDD1.n2 VDD1.t1 1.68992
R99 VDD1.n2 VDD1.t2 1.68992
R100 VDD1 VDD1.n7 0.659983
R101 VDD1 VDD1.n1 0.297914
R102 VDD1.n5 VDD1.n3 0.184378
R103 B.n684 B.n683 585
R104 B.n685 B.n684 585
R105 B.n281 B.n99 585
R106 B.n280 B.n279 585
R107 B.n278 B.n277 585
R108 B.n276 B.n275 585
R109 B.n274 B.n273 585
R110 B.n272 B.n271 585
R111 B.n270 B.n269 585
R112 B.n268 B.n267 585
R113 B.n266 B.n265 585
R114 B.n264 B.n263 585
R115 B.n262 B.n261 585
R116 B.n260 B.n259 585
R117 B.n258 B.n257 585
R118 B.n256 B.n255 585
R119 B.n254 B.n253 585
R120 B.n252 B.n251 585
R121 B.n250 B.n249 585
R122 B.n248 B.n247 585
R123 B.n246 B.n245 585
R124 B.n244 B.n243 585
R125 B.n242 B.n241 585
R126 B.n240 B.n239 585
R127 B.n238 B.n237 585
R128 B.n236 B.n235 585
R129 B.n234 B.n233 585
R130 B.n232 B.n231 585
R131 B.n230 B.n229 585
R132 B.n228 B.n227 585
R133 B.n226 B.n225 585
R134 B.n224 B.n223 585
R135 B.n222 B.n221 585
R136 B.n220 B.n219 585
R137 B.n218 B.n217 585
R138 B.n216 B.n215 585
R139 B.n214 B.n213 585
R140 B.n212 B.n211 585
R141 B.n210 B.n209 585
R142 B.n208 B.n207 585
R143 B.n206 B.n205 585
R144 B.n204 B.n203 585
R145 B.n202 B.n201 585
R146 B.n200 B.n199 585
R147 B.n198 B.n197 585
R148 B.n196 B.n195 585
R149 B.n194 B.n193 585
R150 B.n192 B.n191 585
R151 B.n190 B.n189 585
R152 B.n188 B.n187 585
R153 B.n186 B.n185 585
R154 B.n183 B.n182 585
R155 B.n181 B.n180 585
R156 B.n179 B.n178 585
R157 B.n177 B.n176 585
R158 B.n175 B.n174 585
R159 B.n173 B.n172 585
R160 B.n171 B.n170 585
R161 B.n169 B.n168 585
R162 B.n167 B.n166 585
R163 B.n165 B.n164 585
R164 B.n163 B.n162 585
R165 B.n161 B.n160 585
R166 B.n159 B.n158 585
R167 B.n157 B.n156 585
R168 B.n155 B.n154 585
R169 B.n153 B.n152 585
R170 B.n151 B.n150 585
R171 B.n149 B.n148 585
R172 B.n147 B.n146 585
R173 B.n145 B.n144 585
R174 B.n143 B.n142 585
R175 B.n141 B.n140 585
R176 B.n139 B.n138 585
R177 B.n137 B.n136 585
R178 B.n135 B.n134 585
R179 B.n133 B.n132 585
R180 B.n131 B.n130 585
R181 B.n129 B.n128 585
R182 B.n127 B.n126 585
R183 B.n125 B.n124 585
R184 B.n123 B.n122 585
R185 B.n121 B.n120 585
R186 B.n119 B.n118 585
R187 B.n117 B.n116 585
R188 B.n115 B.n114 585
R189 B.n113 B.n112 585
R190 B.n111 B.n110 585
R191 B.n109 B.n108 585
R192 B.n107 B.n106 585
R193 B.n54 B.n53 585
R194 B.n688 B.n687 585
R195 B.n682 B.n100 585
R196 B.n100 B.n51 585
R197 B.n681 B.n50 585
R198 B.n692 B.n50 585
R199 B.n680 B.n49 585
R200 B.n693 B.n49 585
R201 B.n679 B.n48 585
R202 B.n694 B.n48 585
R203 B.n678 B.n677 585
R204 B.n677 B.n47 585
R205 B.n676 B.n43 585
R206 B.n700 B.n43 585
R207 B.n675 B.n42 585
R208 B.n701 B.n42 585
R209 B.n674 B.n41 585
R210 B.n702 B.n41 585
R211 B.n673 B.n672 585
R212 B.n672 B.n37 585
R213 B.n671 B.n36 585
R214 B.n708 B.n36 585
R215 B.n670 B.n35 585
R216 B.n709 B.n35 585
R217 B.n669 B.n34 585
R218 B.n710 B.n34 585
R219 B.n668 B.n667 585
R220 B.n667 B.n30 585
R221 B.n666 B.n29 585
R222 B.n716 B.n29 585
R223 B.n665 B.n28 585
R224 B.n717 B.n28 585
R225 B.n664 B.n27 585
R226 B.n718 B.n27 585
R227 B.n663 B.n662 585
R228 B.n662 B.n23 585
R229 B.n661 B.n22 585
R230 B.n724 B.n22 585
R231 B.n660 B.n21 585
R232 B.n725 B.n21 585
R233 B.n659 B.n20 585
R234 B.n726 B.n20 585
R235 B.n658 B.n657 585
R236 B.n657 B.n16 585
R237 B.n656 B.n15 585
R238 B.t7 B.n15 585
R239 B.n655 B.n14 585
R240 B.n732 B.n14 585
R241 B.n654 B.n13 585
R242 B.n733 B.n13 585
R243 B.n653 B.n652 585
R244 B.n652 B.n12 585
R245 B.n651 B.n650 585
R246 B.n651 B.n8 585
R247 B.n649 B.n7 585
R248 B.n740 B.n7 585
R249 B.n648 B.n6 585
R250 B.n741 B.n6 585
R251 B.n647 B.n5 585
R252 B.n742 B.n5 585
R253 B.n646 B.n645 585
R254 B.n645 B.n4 585
R255 B.n644 B.n282 585
R256 B.n644 B.n643 585
R257 B.n633 B.n283 585
R258 B.n636 B.n283 585
R259 B.n635 B.n634 585
R260 B.n637 B.n635 585
R261 B.n632 B.n288 585
R262 B.n288 B.n287 585
R263 B.n631 B.n630 585
R264 B.n630 B.t4 585
R265 B.n290 B.n289 585
R266 B.n291 B.n290 585
R267 B.n623 B.n622 585
R268 B.n624 B.n623 585
R269 B.n621 B.n296 585
R270 B.n296 B.n295 585
R271 B.n620 B.n619 585
R272 B.n619 B.n618 585
R273 B.n298 B.n297 585
R274 B.n299 B.n298 585
R275 B.n611 B.n610 585
R276 B.n612 B.n611 585
R277 B.n609 B.n303 585
R278 B.n307 B.n303 585
R279 B.n608 B.n607 585
R280 B.n607 B.n606 585
R281 B.n305 B.n304 585
R282 B.n306 B.n305 585
R283 B.n599 B.n598 585
R284 B.n600 B.n599 585
R285 B.n597 B.n312 585
R286 B.n312 B.n311 585
R287 B.n596 B.n595 585
R288 B.n595 B.n594 585
R289 B.n314 B.n313 585
R290 B.n315 B.n314 585
R291 B.n587 B.n586 585
R292 B.n588 B.n587 585
R293 B.n585 B.n320 585
R294 B.n320 B.n319 585
R295 B.n584 B.n583 585
R296 B.n583 B.n582 585
R297 B.n322 B.n321 585
R298 B.n575 B.n322 585
R299 B.n574 B.n573 585
R300 B.n576 B.n574 585
R301 B.n572 B.n327 585
R302 B.n327 B.n326 585
R303 B.n571 B.n570 585
R304 B.n570 B.n569 585
R305 B.n329 B.n328 585
R306 B.n330 B.n329 585
R307 B.n565 B.n564 585
R308 B.n333 B.n332 585
R309 B.n561 B.n560 585
R310 B.n562 B.n561 585
R311 B.n559 B.n378 585
R312 B.n558 B.n557 585
R313 B.n556 B.n555 585
R314 B.n554 B.n553 585
R315 B.n552 B.n551 585
R316 B.n550 B.n549 585
R317 B.n548 B.n547 585
R318 B.n546 B.n545 585
R319 B.n544 B.n543 585
R320 B.n542 B.n541 585
R321 B.n540 B.n539 585
R322 B.n538 B.n537 585
R323 B.n536 B.n535 585
R324 B.n534 B.n533 585
R325 B.n532 B.n531 585
R326 B.n530 B.n529 585
R327 B.n528 B.n527 585
R328 B.n526 B.n525 585
R329 B.n524 B.n523 585
R330 B.n522 B.n521 585
R331 B.n520 B.n519 585
R332 B.n518 B.n517 585
R333 B.n516 B.n515 585
R334 B.n514 B.n513 585
R335 B.n512 B.n511 585
R336 B.n510 B.n509 585
R337 B.n508 B.n507 585
R338 B.n506 B.n505 585
R339 B.n504 B.n503 585
R340 B.n502 B.n501 585
R341 B.n500 B.n499 585
R342 B.n498 B.n497 585
R343 B.n496 B.n495 585
R344 B.n494 B.n493 585
R345 B.n492 B.n491 585
R346 B.n490 B.n489 585
R347 B.n488 B.n487 585
R348 B.n486 B.n485 585
R349 B.n484 B.n483 585
R350 B.n482 B.n481 585
R351 B.n480 B.n479 585
R352 B.n478 B.n477 585
R353 B.n476 B.n475 585
R354 B.n474 B.n473 585
R355 B.n472 B.n471 585
R356 B.n470 B.n469 585
R357 B.n468 B.n467 585
R358 B.n465 B.n464 585
R359 B.n463 B.n462 585
R360 B.n461 B.n460 585
R361 B.n459 B.n458 585
R362 B.n457 B.n456 585
R363 B.n455 B.n454 585
R364 B.n453 B.n452 585
R365 B.n451 B.n450 585
R366 B.n449 B.n448 585
R367 B.n447 B.n446 585
R368 B.n445 B.n444 585
R369 B.n443 B.n442 585
R370 B.n441 B.n440 585
R371 B.n439 B.n438 585
R372 B.n437 B.n436 585
R373 B.n435 B.n434 585
R374 B.n433 B.n432 585
R375 B.n431 B.n430 585
R376 B.n429 B.n428 585
R377 B.n427 B.n426 585
R378 B.n425 B.n424 585
R379 B.n423 B.n422 585
R380 B.n421 B.n420 585
R381 B.n419 B.n418 585
R382 B.n417 B.n416 585
R383 B.n415 B.n414 585
R384 B.n413 B.n412 585
R385 B.n411 B.n410 585
R386 B.n409 B.n408 585
R387 B.n407 B.n406 585
R388 B.n405 B.n404 585
R389 B.n403 B.n402 585
R390 B.n401 B.n400 585
R391 B.n399 B.n398 585
R392 B.n397 B.n396 585
R393 B.n395 B.n394 585
R394 B.n393 B.n392 585
R395 B.n391 B.n390 585
R396 B.n389 B.n388 585
R397 B.n387 B.n386 585
R398 B.n385 B.n384 585
R399 B.n566 B.n331 585
R400 B.n331 B.n330 585
R401 B.n568 B.n567 585
R402 B.n569 B.n568 585
R403 B.n325 B.n324 585
R404 B.n326 B.n325 585
R405 B.n578 B.n577 585
R406 B.n577 B.n576 585
R407 B.n579 B.n323 585
R408 B.n575 B.n323 585
R409 B.n581 B.n580 585
R410 B.n582 B.n581 585
R411 B.n318 B.n317 585
R412 B.n319 B.n318 585
R413 B.n590 B.n589 585
R414 B.n589 B.n588 585
R415 B.n591 B.n316 585
R416 B.n316 B.n315 585
R417 B.n593 B.n592 585
R418 B.n594 B.n593 585
R419 B.n310 B.n309 585
R420 B.n311 B.n310 585
R421 B.n602 B.n601 585
R422 B.n601 B.n600 585
R423 B.n603 B.n308 585
R424 B.n308 B.n306 585
R425 B.n605 B.n604 585
R426 B.n606 B.n605 585
R427 B.n302 B.n301 585
R428 B.n307 B.n302 585
R429 B.n614 B.n613 585
R430 B.n613 B.n612 585
R431 B.n615 B.n300 585
R432 B.n300 B.n299 585
R433 B.n617 B.n616 585
R434 B.n618 B.n617 585
R435 B.n294 B.n293 585
R436 B.n295 B.n294 585
R437 B.n626 B.n625 585
R438 B.n625 B.n624 585
R439 B.n627 B.n292 585
R440 B.n292 B.n291 585
R441 B.n629 B.n628 585
R442 B.t4 B.n629 585
R443 B.n286 B.n285 585
R444 B.n287 B.n286 585
R445 B.n639 B.n638 585
R446 B.n638 B.n637 585
R447 B.n640 B.n284 585
R448 B.n636 B.n284 585
R449 B.n642 B.n641 585
R450 B.n643 B.n642 585
R451 B.n3 B.n0 585
R452 B.n4 B.n3 585
R453 B.n739 B.n1 585
R454 B.n740 B.n739 585
R455 B.n738 B.n737 585
R456 B.n738 B.n8 585
R457 B.n736 B.n9 585
R458 B.n12 B.n9 585
R459 B.n735 B.n734 585
R460 B.n734 B.n733 585
R461 B.n11 B.n10 585
R462 B.n732 B.n11 585
R463 B.n731 B.n730 585
R464 B.t7 B.n731 585
R465 B.n729 B.n17 585
R466 B.n17 B.n16 585
R467 B.n728 B.n727 585
R468 B.n727 B.n726 585
R469 B.n19 B.n18 585
R470 B.n725 B.n19 585
R471 B.n723 B.n722 585
R472 B.n724 B.n723 585
R473 B.n721 B.n24 585
R474 B.n24 B.n23 585
R475 B.n720 B.n719 585
R476 B.n719 B.n718 585
R477 B.n26 B.n25 585
R478 B.n717 B.n26 585
R479 B.n715 B.n714 585
R480 B.n716 B.n715 585
R481 B.n713 B.n31 585
R482 B.n31 B.n30 585
R483 B.n712 B.n711 585
R484 B.n711 B.n710 585
R485 B.n33 B.n32 585
R486 B.n709 B.n33 585
R487 B.n707 B.n706 585
R488 B.n708 B.n707 585
R489 B.n705 B.n38 585
R490 B.n38 B.n37 585
R491 B.n704 B.n703 585
R492 B.n703 B.n702 585
R493 B.n40 B.n39 585
R494 B.n701 B.n40 585
R495 B.n699 B.n698 585
R496 B.n700 B.n699 585
R497 B.n697 B.n44 585
R498 B.n47 B.n44 585
R499 B.n696 B.n695 585
R500 B.n695 B.n694 585
R501 B.n46 B.n45 585
R502 B.n693 B.n46 585
R503 B.n691 B.n690 585
R504 B.n692 B.n691 585
R505 B.n689 B.n52 585
R506 B.n52 B.n51 585
R507 B.n743 B.n742 585
R508 B.n741 B.n2 585
R509 B.n104 B.t21 564.201
R510 B.n101 B.t17 564.201
R511 B.n382 B.t10 564.201
R512 B.n379 B.t14 564.201
R513 B.n687 B.n52 545.355
R514 B.n684 B.n100 545.355
R515 B.n384 B.n329 545.355
R516 B.n564 B.n331 545.355
R517 B.n685 B.n98 256.663
R518 B.n685 B.n97 256.663
R519 B.n685 B.n96 256.663
R520 B.n685 B.n95 256.663
R521 B.n685 B.n94 256.663
R522 B.n685 B.n93 256.663
R523 B.n685 B.n92 256.663
R524 B.n685 B.n91 256.663
R525 B.n685 B.n90 256.663
R526 B.n685 B.n89 256.663
R527 B.n685 B.n88 256.663
R528 B.n685 B.n87 256.663
R529 B.n685 B.n86 256.663
R530 B.n685 B.n85 256.663
R531 B.n685 B.n84 256.663
R532 B.n685 B.n83 256.663
R533 B.n685 B.n82 256.663
R534 B.n685 B.n81 256.663
R535 B.n685 B.n80 256.663
R536 B.n685 B.n79 256.663
R537 B.n685 B.n78 256.663
R538 B.n685 B.n77 256.663
R539 B.n685 B.n76 256.663
R540 B.n685 B.n75 256.663
R541 B.n685 B.n74 256.663
R542 B.n685 B.n73 256.663
R543 B.n685 B.n72 256.663
R544 B.n685 B.n71 256.663
R545 B.n685 B.n70 256.663
R546 B.n685 B.n69 256.663
R547 B.n685 B.n68 256.663
R548 B.n685 B.n67 256.663
R549 B.n685 B.n66 256.663
R550 B.n685 B.n65 256.663
R551 B.n685 B.n64 256.663
R552 B.n685 B.n63 256.663
R553 B.n685 B.n62 256.663
R554 B.n685 B.n61 256.663
R555 B.n685 B.n60 256.663
R556 B.n685 B.n59 256.663
R557 B.n685 B.n58 256.663
R558 B.n685 B.n57 256.663
R559 B.n685 B.n56 256.663
R560 B.n685 B.n55 256.663
R561 B.n686 B.n685 256.663
R562 B.n563 B.n562 256.663
R563 B.n562 B.n334 256.663
R564 B.n562 B.n335 256.663
R565 B.n562 B.n336 256.663
R566 B.n562 B.n337 256.663
R567 B.n562 B.n338 256.663
R568 B.n562 B.n339 256.663
R569 B.n562 B.n340 256.663
R570 B.n562 B.n341 256.663
R571 B.n562 B.n342 256.663
R572 B.n562 B.n343 256.663
R573 B.n562 B.n344 256.663
R574 B.n562 B.n345 256.663
R575 B.n562 B.n346 256.663
R576 B.n562 B.n347 256.663
R577 B.n562 B.n348 256.663
R578 B.n562 B.n349 256.663
R579 B.n562 B.n350 256.663
R580 B.n562 B.n351 256.663
R581 B.n562 B.n352 256.663
R582 B.n562 B.n353 256.663
R583 B.n562 B.n354 256.663
R584 B.n562 B.n355 256.663
R585 B.n562 B.n356 256.663
R586 B.n562 B.n357 256.663
R587 B.n562 B.n358 256.663
R588 B.n562 B.n359 256.663
R589 B.n562 B.n360 256.663
R590 B.n562 B.n361 256.663
R591 B.n562 B.n362 256.663
R592 B.n562 B.n363 256.663
R593 B.n562 B.n364 256.663
R594 B.n562 B.n365 256.663
R595 B.n562 B.n366 256.663
R596 B.n562 B.n367 256.663
R597 B.n562 B.n368 256.663
R598 B.n562 B.n369 256.663
R599 B.n562 B.n370 256.663
R600 B.n562 B.n371 256.663
R601 B.n562 B.n372 256.663
R602 B.n562 B.n373 256.663
R603 B.n562 B.n374 256.663
R604 B.n562 B.n375 256.663
R605 B.n562 B.n376 256.663
R606 B.n562 B.n377 256.663
R607 B.n745 B.n744 256.663
R608 B.n106 B.n54 163.367
R609 B.n110 B.n109 163.367
R610 B.n114 B.n113 163.367
R611 B.n118 B.n117 163.367
R612 B.n122 B.n121 163.367
R613 B.n126 B.n125 163.367
R614 B.n130 B.n129 163.367
R615 B.n134 B.n133 163.367
R616 B.n138 B.n137 163.367
R617 B.n142 B.n141 163.367
R618 B.n146 B.n145 163.367
R619 B.n150 B.n149 163.367
R620 B.n154 B.n153 163.367
R621 B.n158 B.n157 163.367
R622 B.n162 B.n161 163.367
R623 B.n166 B.n165 163.367
R624 B.n170 B.n169 163.367
R625 B.n174 B.n173 163.367
R626 B.n178 B.n177 163.367
R627 B.n182 B.n181 163.367
R628 B.n187 B.n186 163.367
R629 B.n191 B.n190 163.367
R630 B.n195 B.n194 163.367
R631 B.n199 B.n198 163.367
R632 B.n203 B.n202 163.367
R633 B.n207 B.n206 163.367
R634 B.n211 B.n210 163.367
R635 B.n215 B.n214 163.367
R636 B.n219 B.n218 163.367
R637 B.n223 B.n222 163.367
R638 B.n227 B.n226 163.367
R639 B.n231 B.n230 163.367
R640 B.n235 B.n234 163.367
R641 B.n239 B.n238 163.367
R642 B.n243 B.n242 163.367
R643 B.n247 B.n246 163.367
R644 B.n251 B.n250 163.367
R645 B.n255 B.n254 163.367
R646 B.n259 B.n258 163.367
R647 B.n263 B.n262 163.367
R648 B.n267 B.n266 163.367
R649 B.n271 B.n270 163.367
R650 B.n275 B.n274 163.367
R651 B.n279 B.n278 163.367
R652 B.n684 B.n99 163.367
R653 B.n570 B.n329 163.367
R654 B.n570 B.n327 163.367
R655 B.n574 B.n327 163.367
R656 B.n574 B.n322 163.367
R657 B.n583 B.n322 163.367
R658 B.n583 B.n320 163.367
R659 B.n587 B.n320 163.367
R660 B.n587 B.n314 163.367
R661 B.n595 B.n314 163.367
R662 B.n595 B.n312 163.367
R663 B.n599 B.n312 163.367
R664 B.n599 B.n305 163.367
R665 B.n607 B.n305 163.367
R666 B.n607 B.n303 163.367
R667 B.n611 B.n303 163.367
R668 B.n611 B.n298 163.367
R669 B.n619 B.n298 163.367
R670 B.n619 B.n296 163.367
R671 B.n623 B.n296 163.367
R672 B.n623 B.n290 163.367
R673 B.n630 B.n290 163.367
R674 B.n630 B.n288 163.367
R675 B.n635 B.n288 163.367
R676 B.n635 B.n283 163.367
R677 B.n644 B.n283 163.367
R678 B.n645 B.n644 163.367
R679 B.n645 B.n5 163.367
R680 B.n6 B.n5 163.367
R681 B.n7 B.n6 163.367
R682 B.n651 B.n7 163.367
R683 B.n652 B.n651 163.367
R684 B.n652 B.n13 163.367
R685 B.n14 B.n13 163.367
R686 B.n15 B.n14 163.367
R687 B.n657 B.n15 163.367
R688 B.n657 B.n20 163.367
R689 B.n21 B.n20 163.367
R690 B.n22 B.n21 163.367
R691 B.n662 B.n22 163.367
R692 B.n662 B.n27 163.367
R693 B.n28 B.n27 163.367
R694 B.n29 B.n28 163.367
R695 B.n667 B.n29 163.367
R696 B.n667 B.n34 163.367
R697 B.n35 B.n34 163.367
R698 B.n36 B.n35 163.367
R699 B.n672 B.n36 163.367
R700 B.n672 B.n41 163.367
R701 B.n42 B.n41 163.367
R702 B.n43 B.n42 163.367
R703 B.n677 B.n43 163.367
R704 B.n677 B.n48 163.367
R705 B.n49 B.n48 163.367
R706 B.n50 B.n49 163.367
R707 B.n100 B.n50 163.367
R708 B.n561 B.n333 163.367
R709 B.n561 B.n378 163.367
R710 B.n557 B.n556 163.367
R711 B.n553 B.n552 163.367
R712 B.n549 B.n548 163.367
R713 B.n545 B.n544 163.367
R714 B.n541 B.n540 163.367
R715 B.n537 B.n536 163.367
R716 B.n533 B.n532 163.367
R717 B.n529 B.n528 163.367
R718 B.n525 B.n524 163.367
R719 B.n521 B.n520 163.367
R720 B.n517 B.n516 163.367
R721 B.n513 B.n512 163.367
R722 B.n509 B.n508 163.367
R723 B.n505 B.n504 163.367
R724 B.n501 B.n500 163.367
R725 B.n497 B.n496 163.367
R726 B.n493 B.n492 163.367
R727 B.n489 B.n488 163.367
R728 B.n485 B.n484 163.367
R729 B.n481 B.n480 163.367
R730 B.n477 B.n476 163.367
R731 B.n473 B.n472 163.367
R732 B.n469 B.n468 163.367
R733 B.n464 B.n463 163.367
R734 B.n460 B.n459 163.367
R735 B.n456 B.n455 163.367
R736 B.n452 B.n451 163.367
R737 B.n448 B.n447 163.367
R738 B.n444 B.n443 163.367
R739 B.n440 B.n439 163.367
R740 B.n436 B.n435 163.367
R741 B.n432 B.n431 163.367
R742 B.n428 B.n427 163.367
R743 B.n424 B.n423 163.367
R744 B.n420 B.n419 163.367
R745 B.n416 B.n415 163.367
R746 B.n412 B.n411 163.367
R747 B.n408 B.n407 163.367
R748 B.n404 B.n403 163.367
R749 B.n400 B.n399 163.367
R750 B.n396 B.n395 163.367
R751 B.n392 B.n391 163.367
R752 B.n388 B.n387 163.367
R753 B.n568 B.n331 163.367
R754 B.n568 B.n325 163.367
R755 B.n577 B.n325 163.367
R756 B.n577 B.n323 163.367
R757 B.n581 B.n323 163.367
R758 B.n581 B.n318 163.367
R759 B.n589 B.n318 163.367
R760 B.n589 B.n316 163.367
R761 B.n593 B.n316 163.367
R762 B.n593 B.n310 163.367
R763 B.n601 B.n310 163.367
R764 B.n601 B.n308 163.367
R765 B.n605 B.n308 163.367
R766 B.n605 B.n302 163.367
R767 B.n613 B.n302 163.367
R768 B.n613 B.n300 163.367
R769 B.n617 B.n300 163.367
R770 B.n617 B.n294 163.367
R771 B.n625 B.n294 163.367
R772 B.n625 B.n292 163.367
R773 B.n629 B.n292 163.367
R774 B.n629 B.n286 163.367
R775 B.n638 B.n286 163.367
R776 B.n638 B.n284 163.367
R777 B.n642 B.n284 163.367
R778 B.n642 B.n3 163.367
R779 B.n743 B.n3 163.367
R780 B.n739 B.n2 163.367
R781 B.n739 B.n738 163.367
R782 B.n738 B.n9 163.367
R783 B.n734 B.n9 163.367
R784 B.n734 B.n11 163.367
R785 B.n731 B.n11 163.367
R786 B.n731 B.n17 163.367
R787 B.n727 B.n17 163.367
R788 B.n727 B.n19 163.367
R789 B.n723 B.n19 163.367
R790 B.n723 B.n24 163.367
R791 B.n719 B.n24 163.367
R792 B.n719 B.n26 163.367
R793 B.n715 B.n26 163.367
R794 B.n715 B.n31 163.367
R795 B.n711 B.n31 163.367
R796 B.n711 B.n33 163.367
R797 B.n707 B.n33 163.367
R798 B.n707 B.n38 163.367
R799 B.n703 B.n38 163.367
R800 B.n703 B.n40 163.367
R801 B.n699 B.n40 163.367
R802 B.n699 B.n44 163.367
R803 B.n695 B.n44 163.367
R804 B.n695 B.n46 163.367
R805 B.n691 B.n46 163.367
R806 B.n691 B.n52 163.367
R807 B.n101 B.t19 92.4591
R808 B.n382 B.t13 92.4591
R809 B.n104 B.t22 92.4444
R810 B.n379 B.t16 92.4444
R811 B.n562 B.n330 88.6736
R812 B.n685 B.n51 88.6736
R813 B.n687 B.n686 71.676
R814 B.n106 B.n55 71.676
R815 B.n110 B.n56 71.676
R816 B.n114 B.n57 71.676
R817 B.n118 B.n58 71.676
R818 B.n122 B.n59 71.676
R819 B.n126 B.n60 71.676
R820 B.n130 B.n61 71.676
R821 B.n134 B.n62 71.676
R822 B.n138 B.n63 71.676
R823 B.n142 B.n64 71.676
R824 B.n146 B.n65 71.676
R825 B.n150 B.n66 71.676
R826 B.n154 B.n67 71.676
R827 B.n158 B.n68 71.676
R828 B.n162 B.n69 71.676
R829 B.n166 B.n70 71.676
R830 B.n170 B.n71 71.676
R831 B.n174 B.n72 71.676
R832 B.n178 B.n73 71.676
R833 B.n182 B.n74 71.676
R834 B.n187 B.n75 71.676
R835 B.n191 B.n76 71.676
R836 B.n195 B.n77 71.676
R837 B.n199 B.n78 71.676
R838 B.n203 B.n79 71.676
R839 B.n207 B.n80 71.676
R840 B.n211 B.n81 71.676
R841 B.n215 B.n82 71.676
R842 B.n219 B.n83 71.676
R843 B.n223 B.n84 71.676
R844 B.n227 B.n85 71.676
R845 B.n231 B.n86 71.676
R846 B.n235 B.n87 71.676
R847 B.n239 B.n88 71.676
R848 B.n243 B.n89 71.676
R849 B.n247 B.n90 71.676
R850 B.n251 B.n91 71.676
R851 B.n255 B.n92 71.676
R852 B.n259 B.n93 71.676
R853 B.n263 B.n94 71.676
R854 B.n267 B.n95 71.676
R855 B.n271 B.n96 71.676
R856 B.n275 B.n97 71.676
R857 B.n279 B.n98 71.676
R858 B.n99 B.n98 71.676
R859 B.n278 B.n97 71.676
R860 B.n274 B.n96 71.676
R861 B.n270 B.n95 71.676
R862 B.n266 B.n94 71.676
R863 B.n262 B.n93 71.676
R864 B.n258 B.n92 71.676
R865 B.n254 B.n91 71.676
R866 B.n250 B.n90 71.676
R867 B.n246 B.n89 71.676
R868 B.n242 B.n88 71.676
R869 B.n238 B.n87 71.676
R870 B.n234 B.n86 71.676
R871 B.n230 B.n85 71.676
R872 B.n226 B.n84 71.676
R873 B.n222 B.n83 71.676
R874 B.n218 B.n82 71.676
R875 B.n214 B.n81 71.676
R876 B.n210 B.n80 71.676
R877 B.n206 B.n79 71.676
R878 B.n202 B.n78 71.676
R879 B.n198 B.n77 71.676
R880 B.n194 B.n76 71.676
R881 B.n190 B.n75 71.676
R882 B.n186 B.n74 71.676
R883 B.n181 B.n73 71.676
R884 B.n177 B.n72 71.676
R885 B.n173 B.n71 71.676
R886 B.n169 B.n70 71.676
R887 B.n165 B.n69 71.676
R888 B.n161 B.n68 71.676
R889 B.n157 B.n67 71.676
R890 B.n153 B.n66 71.676
R891 B.n149 B.n65 71.676
R892 B.n145 B.n64 71.676
R893 B.n141 B.n63 71.676
R894 B.n137 B.n62 71.676
R895 B.n133 B.n61 71.676
R896 B.n129 B.n60 71.676
R897 B.n125 B.n59 71.676
R898 B.n121 B.n58 71.676
R899 B.n117 B.n57 71.676
R900 B.n113 B.n56 71.676
R901 B.n109 B.n55 71.676
R902 B.n686 B.n54 71.676
R903 B.n564 B.n563 71.676
R904 B.n378 B.n334 71.676
R905 B.n556 B.n335 71.676
R906 B.n552 B.n336 71.676
R907 B.n548 B.n337 71.676
R908 B.n544 B.n338 71.676
R909 B.n540 B.n339 71.676
R910 B.n536 B.n340 71.676
R911 B.n532 B.n341 71.676
R912 B.n528 B.n342 71.676
R913 B.n524 B.n343 71.676
R914 B.n520 B.n344 71.676
R915 B.n516 B.n345 71.676
R916 B.n512 B.n346 71.676
R917 B.n508 B.n347 71.676
R918 B.n504 B.n348 71.676
R919 B.n500 B.n349 71.676
R920 B.n496 B.n350 71.676
R921 B.n492 B.n351 71.676
R922 B.n488 B.n352 71.676
R923 B.n484 B.n353 71.676
R924 B.n480 B.n354 71.676
R925 B.n476 B.n355 71.676
R926 B.n472 B.n356 71.676
R927 B.n468 B.n357 71.676
R928 B.n463 B.n358 71.676
R929 B.n459 B.n359 71.676
R930 B.n455 B.n360 71.676
R931 B.n451 B.n361 71.676
R932 B.n447 B.n362 71.676
R933 B.n443 B.n363 71.676
R934 B.n439 B.n364 71.676
R935 B.n435 B.n365 71.676
R936 B.n431 B.n366 71.676
R937 B.n427 B.n367 71.676
R938 B.n423 B.n368 71.676
R939 B.n419 B.n369 71.676
R940 B.n415 B.n370 71.676
R941 B.n411 B.n371 71.676
R942 B.n407 B.n372 71.676
R943 B.n403 B.n373 71.676
R944 B.n399 B.n374 71.676
R945 B.n395 B.n375 71.676
R946 B.n391 B.n376 71.676
R947 B.n387 B.n377 71.676
R948 B.n563 B.n333 71.676
R949 B.n557 B.n334 71.676
R950 B.n553 B.n335 71.676
R951 B.n549 B.n336 71.676
R952 B.n545 B.n337 71.676
R953 B.n541 B.n338 71.676
R954 B.n537 B.n339 71.676
R955 B.n533 B.n340 71.676
R956 B.n529 B.n341 71.676
R957 B.n525 B.n342 71.676
R958 B.n521 B.n343 71.676
R959 B.n517 B.n344 71.676
R960 B.n513 B.n345 71.676
R961 B.n509 B.n346 71.676
R962 B.n505 B.n347 71.676
R963 B.n501 B.n348 71.676
R964 B.n497 B.n349 71.676
R965 B.n493 B.n350 71.676
R966 B.n489 B.n351 71.676
R967 B.n485 B.n352 71.676
R968 B.n481 B.n353 71.676
R969 B.n477 B.n354 71.676
R970 B.n473 B.n355 71.676
R971 B.n469 B.n356 71.676
R972 B.n464 B.n357 71.676
R973 B.n460 B.n358 71.676
R974 B.n456 B.n359 71.676
R975 B.n452 B.n360 71.676
R976 B.n448 B.n361 71.676
R977 B.n444 B.n362 71.676
R978 B.n440 B.n363 71.676
R979 B.n436 B.n364 71.676
R980 B.n432 B.n365 71.676
R981 B.n428 B.n366 71.676
R982 B.n424 B.n367 71.676
R983 B.n420 B.n368 71.676
R984 B.n416 B.n369 71.676
R985 B.n412 B.n370 71.676
R986 B.n408 B.n371 71.676
R987 B.n404 B.n372 71.676
R988 B.n400 B.n373 71.676
R989 B.n396 B.n374 71.676
R990 B.n392 B.n375 71.676
R991 B.n388 B.n376 71.676
R992 B.n384 B.n377 71.676
R993 B.n744 B.n743 71.676
R994 B.n744 B.n2 71.676
R995 B.n102 B.t20 70.9318
R996 B.n383 B.t12 70.9318
R997 B.n105 B.t23 70.9171
R998 B.n380 B.t15 70.9171
R999 B.n184 B.n105 59.5399
R1000 B.n103 B.n102 59.5399
R1001 B.n466 B.n383 59.5399
R1002 B.n381 B.n380 59.5399
R1003 B.n569 B.n330 44.0134
R1004 B.n569 B.n326 44.0134
R1005 B.n576 B.n326 44.0134
R1006 B.n576 B.n575 44.0134
R1007 B.n582 B.n319 44.0134
R1008 B.n588 B.n319 44.0134
R1009 B.n588 B.n315 44.0134
R1010 B.n594 B.n315 44.0134
R1011 B.n594 B.n311 44.0134
R1012 B.n600 B.n311 44.0134
R1013 B.n606 B.n306 44.0134
R1014 B.n606 B.n307 44.0134
R1015 B.n612 B.n299 44.0134
R1016 B.n618 B.n299 44.0134
R1017 B.n624 B.n295 44.0134
R1018 B.n624 B.n291 44.0134
R1019 B.t4 B.n291 44.0134
R1020 B.t4 B.n287 44.0134
R1021 B.n637 B.n287 44.0134
R1022 B.n637 B.n636 44.0134
R1023 B.n643 B.n4 44.0134
R1024 B.n742 B.n4 44.0134
R1025 B.n742 B.n741 44.0134
R1026 B.n741 B.n740 44.0134
R1027 B.n740 B.n8 44.0134
R1028 B.n733 B.n12 44.0134
R1029 B.n733 B.n732 44.0134
R1030 B.n732 B.t7 44.0134
R1031 B.t7 B.n16 44.0134
R1032 B.n726 B.n16 44.0134
R1033 B.n726 B.n725 44.0134
R1034 B.n724 B.n23 44.0134
R1035 B.n718 B.n23 44.0134
R1036 B.n717 B.n716 44.0134
R1037 B.n716 B.n30 44.0134
R1038 B.n710 B.n709 44.0134
R1039 B.n709 B.n708 44.0134
R1040 B.n708 B.n37 44.0134
R1041 B.n702 B.n37 44.0134
R1042 B.n702 B.n701 44.0134
R1043 B.n701 B.n700 44.0134
R1044 B.n694 B.n47 44.0134
R1045 B.n694 B.n693 44.0134
R1046 B.n693 B.n692 44.0134
R1047 B.n692 B.n51 44.0134
R1048 B.n683 B.n682 35.4346
R1049 B.n566 B.n565 35.4346
R1050 B.n385 B.n328 35.4346
R1051 B.n689 B.n688 35.4346
R1052 B.t0 B.n306 34.952
R1053 B.t5 B.n30 34.952
R1054 B.n575 B.t11 32.363
R1055 B.n618 B.t9 32.363
R1056 B.n643 B.t8 32.363
R1057 B.t6 B.n8 32.363
R1058 B.t2 B.n724 32.363
R1059 B.n47 B.t18 32.363
R1060 B.n612 B.t3 23.3015
R1061 B.n718 B.t1 23.3015
R1062 B.n105 B.n104 21.5278
R1063 B.n102 B.n101 21.5278
R1064 B.n383 B.n382 21.5278
R1065 B.n380 B.n379 21.5278
R1066 B.n307 B.t3 20.7125
R1067 B.t1 B.n717 20.7125
R1068 B B.n745 18.0485
R1069 B.n582 B.t11 11.651
R1070 B.t9 B.n295 11.651
R1071 B.n636 B.t8 11.651
R1072 B.n12 B.t6 11.651
R1073 B.n725 B.t2 11.651
R1074 B.n700 B.t18 11.651
R1075 B.n567 B.n566 10.6151
R1076 B.n567 B.n324 10.6151
R1077 B.n578 B.n324 10.6151
R1078 B.n579 B.n578 10.6151
R1079 B.n580 B.n579 10.6151
R1080 B.n580 B.n317 10.6151
R1081 B.n590 B.n317 10.6151
R1082 B.n591 B.n590 10.6151
R1083 B.n592 B.n591 10.6151
R1084 B.n592 B.n309 10.6151
R1085 B.n602 B.n309 10.6151
R1086 B.n603 B.n602 10.6151
R1087 B.n604 B.n603 10.6151
R1088 B.n604 B.n301 10.6151
R1089 B.n614 B.n301 10.6151
R1090 B.n615 B.n614 10.6151
R1091 B.n616 B.n615 10.6151
R1092 B.n616 B.n293 10.6151
R1093 B.n626 B.n293 10.6151
R1094 B.n627 B.n626 10.6151
R1095 B.n628 B.n627 10.6151
R1096 B.n628 B.n285 10.6151
R1097 B.n639 B.n285 10.6151
R1098 B.n640 B.n639 10.6151
R1099 B.n641 B.n640 10.6151
R1100 B.n641 B.n0 10.6151
R1101 B.n565 B.n332 10.6151
R1102 B.n560 B.n332 10.6151
R1103 B.n560 B.n559 10.6151
R1104 B.n559 B.n558 10.6151
R1105 B.n558 B.n555 10.6151
R1106 B.n555 B.n554 10.6151
R1107 B.n554 B.n551 10.6151
R1108 B.n551 B.n550 10.6151
R1109 B.n550 B.n547 10.6151
R1110 B.n547 B.n546 10.6151
R1111 B.n546 B.n543 10.6151
R1112 B.n543 B.n542 10.6151
R1113 B.n542 B.n539 10.6151
R1114 B.n539 B.n538 10.6151
R1115 B.n538 B.n535 10.6151
R1116 B.n535 B.n534 10.6151
R1117 B.n534 B.n531 10.6151
R1118 B.n531 B.n530 10.6151
R1119 B.n530 B.n527 10.6151
R1120 B.n527 B.n526 10.6151
R1121 B.n526 B.n523 10.6151
R1122 B.n523 B.n522 10.6151
R1123 B.n522 B.n519 10.6151
R1124 B.n519 B.n518 10.6151
R1125 B.n518 B.n515 10.6151
R1126 B.n515 B.n514 10.6151
R1127 B.n514 B.n511 10.6151
R1128 B.n511 B.n510 10.6151
R1129 B.n510 B.n507 10.6151
R1130 B.n507 B.n506 10.6151
R1131 B.n506 B.n503 10.6151
R1132 B.n503 B.n502 10.6151
R1133 B.n502 B.n499 10.6151
R1134 B.n499 B.n498 10.6151
R1135 B.n498 B.n495 10.6151
R1136 B.n495 B.n494 10.6151
R1137 B.n494 B.n491 10.6151
R1138 B.n491 B.n490 10.6151
R1139 B.n490 B.n487 10.6151
R1140 B.n487 B.n486 10.6151
R1141 B.n483 B.n482 10.6151
R1142 B.n482 B.n479 10.6151
R1143 B.n479 B.n478 10.6151
R1144 B.n478 B.n475 10.6151
R1145 B.n475 B.n474 10.6151
R1146 B.n474 B.n471 10.6151
R1147 B.n471 B.n470 10.6151
R1148 B.n470 B.n467 10.6151
R1149 B.n465 B.n462 10.6151
R1150 B.n462 B.n461 10.6151
R1151 B.n461 B.n458 10.6151
R1152 B.n458 B.n457 10.6151
R1153 B.n457 B.n454 10.6151
R1154 B.n454 B.n453 10.6151
R1155 B.n453 B.n450 10.6151
R1156 B.n450 B.n449 10.6151
R1157 B.n449 B.n446 10.6151
R1158 B.n446 B.n445 10.6151
R1159 B.n445 B.n442 10.6151
R1160 B.n442 B.n441 10.6151
R1161 B.n441 B.n438 10.6151
R1162 B.n438 B.n437 10.6151
R1163 B.n437 B.n434 10.6151
R1164 B.n434 B.n433 10.6151
R1165 B.n433 B.n430 10.6151
R1166 B.n430 B.n429 10.6151
R1167 B.n429 B.n426 10.6151
R1168 B.n426 B.n425 10.6151
R1169 B.n425 B.n422 10.6151
R1170 B.n422 B.n421 10.6151
R1171 B.n421 B.n418 10.6151
R1172 B.n418 B.n417 10.6151
R1173 B.n417 B.n414 10.6151
R1174 B.n414 B.n413 10.6151
R1175 B.n413 B.n410 10.6151
R1176 B.n410 B.n409 10.6151
R1177 B.n409 B.n406 10.6151
R1178 B.n406 B.n405 10.6151
R1179 B.n405 B.n402 10.6151
R1180 B.n402 B.n401 10.6151
R1181 B.n401 B.n398 10.6151
R1182 B.n398 B.n397 10.6151
R1183 B.n397 B.n394 10.6151
R1184 B.n394 B.n393 10.6151
R1185 B.n393 B.n390 10.6151
R1186 B.n390 B.n389 10.6151
R1187 B.n389 B.n386 10.6151
R1188 B.n386 B.n385 10.6151
R1189 B.n571 B.n328 10.6151
R1190 B.n572 B.n571 10.6151
R1191 B.n573 B.n572 10.6151
R1192 B.n573 B.n321 10.6151
R1193 B.n584 B.n321 10.6151
R1194 B.n585 B.n584 10.6151
R1195 B.n586 B.n585 10.6151
R1196 B.n586 B.n313 10.6151
R1197 B.n596 B.n313 10.6151
R1198 B.n597 B.n596 10.6151
R1199 B.n598 B.n597 10.6151
R1200 B.n598 B.n304 10.6151
R1201 B.n608 B.n304 10.6151
R1202 B.n609 B.n608 10.6151
R1203 B.n610 B.n609 10.6151
R1204 B.n610 B.n297 10.6151
R1205 B.n620 B.n297 10.6151
R1206 B.n621 B.n620 10.6151
R1207 B.n622 B.n621 10.6151
R1208 B.n622 B.n289 10.6151
R1209 B.n631 B.n289 10.6151
R1210 B.n632 B.n631 10.6151
R1211 B.n634 B.n632 10.6151
R1212 B.n634 B.n633 10.6151
R1213 B.n633 B.n282 10.6151
R1214 B.n646 B.n282 10.6151
R1215 B.n647 B.n646 10.6151
R1216 B.n648 B.n647 10.6151
R1217 B.n649 B.n648 10.6151
R1218 B.n650 B.n649 10.6151
R1219 B.n653 B.n650 10.6151
R1220 B.n654 B.n653 10.6151
R1221 B.n655 B.n654 10.6151
R1222 B.n656 B.n655 10.6151
R1223 B.n658 B.n656 10.6151
R1224 B.n659 B.n658 10.6151
R1225 B.n660 B.n659 10.6151
R1226 B.n661 B.n660 10.6151
R1227 B.n663 B.n661 10.6151
R1228 B.n664 B.n663 10.6151
R1229 B.n665 B.n664 10.6151
R1230 B.n666 B.n665 10.6151
R1231 B.n668 B.n666 10.6151
R1232 B.n669 B.n668 10.6151
R1233 B.n670 B.n669 10.6151
R1234 B.n671 B.n670 10.6151
R1235 B.n673 B.n671 10.6151
R1236 B.n674 B.n673 10.6151
R1237 B.n675 B.n674 10.6151
R1238 B.n676 B.n675 10.6151
R1239 B.n678 B.n676 10.6151
R1240 B.n679 B.n678 10.6151
R1241 B.n680 B.n679 10.6151
R1242 B.n681 B.n680 10.6151
R1243 B.n682 B.n681 10.6151
R1244 B.n737 B.n1 10.6151
R1245 B.n737 B.n736 10.6151
R1246 B.n736 B.n735 10.6151
R1247 B.n735 B.n10 10.6151
R1248 B.n730 B.n10 10.6151
R1249 B.n730 B.n729 10.6151
R1250 B.n729 B.n728 10.6151
R1251 B.n728 B.n18 10.6151
R1252 B.n722 B.n18 10.6151
R1253 B.n722 B.n721 10.6151
R1254 B.n721 B.n720 10.6151
R1255 B.n720 B.n25 10.6151
R1256 B.n714 B.n25 10.6151
R1257 B.n714 B.n713 10.6151
R1258 B.n713 B.n712 10.6151
R1259 B.n712 B.n32 10.6151
R1260 B.n706 B.n32 10.6151
R1261 B.n706 B.n705 10.6151
R1262 B.n705 B.n704 10.6151
R1263 B.n704 B.n39 10.6151
R1264 B.n698 B.n39 10.6151
R1265 B.n698 B.n697 10.6151
R1266 B.n697 B.n696 10.6151
R1267 B.n696 B.n45 10.6151
R1268 B.n690 B.n45 10.6151
R1269 B.n690 B.n689 10.6151
R1270 B.n688 B.n53 10.6151
R1271 B.n107 B.n53 10.6151
R1272 B.n108 B.n107 10.6151
R1273 B.n111 B.n108 10.6151
R1274 B.n112 B.n111 10.6151
R1275 B.n115 B.n112 10.6151
R1276 B.n116 B.n115 10.6151
R1277 B.n119 B.n116 10.6151
R1278 B.n120 B.n119 10.6151
R1279 B.n123 B.n120 10.6151
R1280 B.n124 B.n123 10.6151
R1281 B.n127 B.n124 10.6151
R1282 B.n128 B.n127 10.6151
R1283 B.n131 B.n128 10.6151
R1284 B.n132 B.n131 10.6151
R1285 B.n135 B.n132 10.6151
R1286 B.n136 B.n135 10.6151
R1287 B.n139 B.n136 10.6151
R1288 B.n140 B.n139 10.6151
R1289 B.n143 B.n140 10.6151
R1290 B.n144 B.n143 10.6151
R1291 B.n147 B.n144 10.6151
R1292 B.n148 B.n147 10.6151
R1293 B.n151 B.n148 10.6151
R1294 B.n152 B.n151 10.6151
R1295 B.n155 B.n152 10.6151
R1296 B.n156 B.n155 10.6151
R1297 B.n159 B.n156 10.6151
R1298 B.n160 B.n159 10.6151
R1299 B.n163 B.n160 10.6151
R1300 B.n164 B.n163 10.6151
R1301 B.n167 B.n164 10.6151
R1302 B.n168 B.n167 10.6151
R1303 B.n171 B.n168 10.6151
R1304 B.n172 B.n171 10.6151
R1305 B.n175 B.n172 10.6151
R1306 B.n176 B.n175 10.6151
R1307 B.n179 B.n176 10.6151
R1308 B.n180 B.n179 10.6151
R1309 B.n183 B.n180 10.6151
R1310 B.n188 B.n185 10.6151
R1311 B.n189 B.n188 10.6151
R1312 B.n192 B.n189 10.6151
R1313 B.n193 B.n192 10.6151
R1314 B.n196 B.n193 10.6151
R1315 B.n197 B.n196 10.6151
R1316 B.n200 B.n197 10.6151
R1317 B.n201 B.n200 10.6151
R1318 B.n205 B.n204 10.6151
R1319 B.n208 B.n205 10.6151
R1320 B.n209 B.n208 10.6151
R1321 B.n212 B.n209 10.6151
R1322 B.n213 B.n212 10.6151
R1323 B.n216 B.n213 10.6151
R1324 B.n217 B.n216 10.6151
R1325 B.n220 B.n217 10.6151
R1326 B.n221 B.n220 10.6151
R1327 B.n224 B.n221 10.6151
R1328 B.n225 B.n224 10.6151
R1329 B.n228 B.n225 10.6151
R1330 B.n229 B.n228 10.6151
R1331 B.n232 B.n229 10.6151
R1332 B.n233 B.n232 10.6151
R1333 B.n236 B.n233 10.6151
R1334 B.n237 B.n236 10.6151
R1335 B.n240 B.n237 10.6151
R1336 B.n241 B.n240 10.6151
R1337 B.n244 B.n241 10.6151
R1338 B.n245 B.n244 10.6151
R1339 B.n248 B.n245 10.6151
R1340 B.n249 B.n248 10.6151
R1341 B.n252 B.n249 10.6151
R1342 B.n253 B.n252 10.6151
R1343 B.n256 B.n253 10.6151
R1344 B.n257 B.n256 10.6151
R1345 B.n260 B.n257 10.6151
R1346 B.n261 B.n260 10.6151
R1347 B.n264 B.n261 10.6151
R1348 B.n265 B.n264 10.6151
R1349 B.n268 B.n265 10.6151
R1350 B.n269 B.n268 10.6151
R1351 B.n272 B.n269 10.6151
R1352 B.n273 B.n272 10.6151
R1353 B.n276 B.n273 10.6151
R1354 B.n277 B.n276 10.6151
R1355 B.n280 B.n277 10.6151
R1356 B.n281 B.n280 10.6151
R1357 B.n683 B.n281 10.6151
R1358 B.n600 B.t0 9.06199
R1359 B.n710 B.t5 9.06199
R1360 B.n745 B.n0 8.11757
R1361 B.n745 B.n1 8.11757
R1362 B.n483 B.n381 6.5566
R1363 B.n467 B.n466 6.5566
R1364 B.n185 B.n184 6.5566
R1365 B.n201 B.n103 6.5566
R1366 B.n486 B.n381 4.05904
R1367 B.n466 B.n465 4.05904
R1368 B.n184 B.n183 4.05904
R1369 B.n204 B.n103 4.05904
R1370 VN.n3 VN.t3 435.139
R1371 VN.n13 VN.t5 435.139
R1372 VN.n2 VN.t4 413.099
R1373 VN.n1 VN.t1 413.099
R1374 VN.n6 VN.t7 413.099
R1375 VN.n8 VN.t2 413.099
R1376 VN.n12 VN.t8 413.099
R1377 VN.n11 VN.t0 413.099
R1378 VN.n16 VN.t6 413.099
R1379 VN.n18 VN.t9 413.099
R1380 VN.n9 VN.n8 161.3
R1381 VN.n19 VN.n18 161.3
R1382 VN.n17 VN.n10 161.3
R1383 VN.n7 VN.n0 161.3
R1384 VN.n16 VN.n15 80.6037
R1385 VN.n14 VN.n11 80.6037
R1386 VN.n6 VN.n5 80.6037
R1387 VN.n4 VN.n1 80.6037
R1388 VN.n2 VN.n1 48.2005
R1389 VN.n6 VN.n1 48.2005
R1390 VN.n12 VN.n11 48.2005
R1391 VN.n16 VN.n11 48.2005
R1392 VN VN.n19 43.3395
R1393 VN.n7 VN.n6 36.5157
R1394 VN.n17 VN.n16 36.5157
R1395 VN.n14 VN.n13 31.7379
R1396 VN.n4 VN.n3 31.7379
R1397 VN.n3 VN.n2 16.9109
R1398 VN.n13 VN.n12 16.9109
R1399 VN.n8 VN.n7 11.6853
R1400 VN.n18 VN.n17 11.6853
R1401 VN.n15 VN.n14 0.380177
R1402 VN.n5 VN.n4 0.380177
R1403 VN.n15 VN.n10 0.285035
R1404 VN.n5 VN.n0 0.285035
R1405 VN.n19 VN.n10 0.189894
R1406 VN.n9 VN.n0 0.189894
R1407 VN VN.n9 0.0516364
R1408 VDD2.n1 VDD2.t6 63.8504
R1409 VDD2.n4 VDD2.t0 62.8937
R1410 VDD2.n3 VDD2.n2 61.8664
R1411 VDD2 VDD2.n7 61.8636
R1412 VDD2.n6 VDD2.n5 61.2043
R1413 VDD2.n1 VDD2.n0 61.204
R1414 VDD2.n4 VDD2.n3 38.364
R1415 VDD2.n7 VDD2.t1 1.68992
R1416 VDD2.n7 VDD2.t4 1.68992
R1417 VDD2.n5 VDD2.t3 1.68992
R1418 VDD2.n5 VDD2.t9 1.68992
R1419 VDD2.n2 VDD2.t2 1.68992
R1420 VDD2.n2 VDD2.t7 1.68992
R1421 VDD2.n0 VDD2.t5 1.68992
R1422 VDD2.n0 VDD2.t8 1.68992
R1423 VDD2.n6 VDD2.n4 0.957397
R1424 VDD2 VDD2.n6 0.297914
R1425 VDD2.n3 VDD2.n1 0.184378
C0 VN VDD1 0.148847f
C1 VN VP 5.66948f
C2 VTAIL VDD1 13.3161f
C3 VTAIL VP 6.81848f
C4 VDD2 VDD1 1.02238f
C5 VDD2 VP 0.351352f
C6 VTAIL VN 6.80391f
C7 VDD1 VP 7.11382f
C8 VN VDD2 6.91583f
C9 VTAIL VDD2 13.3513f
C10 VDD2 B 5.020462f
C11 VDD1 B 4.949712f
C12 VTAIL B 6.495539f
C13 VN B 9.77287f
C14 VP B 7.871217f
C15 VDD2.t6 B 2.53407f
C16 VDD2.t5 B 0.223092f
C17 VDD2.t8 B 0.223092f
C18 VDD2.n0 B 1.98408f
C19 VDD2.n1 B 0.633929f
C20 VDD2.t2 B 0.223092f
C21 VDD2.t7 B 0.223092f
C22 VDD2.n2 B 1.98768f
C23 VDD2.n3 B 1.8602f
C24 VDD2.t0 B 2.52887f
C25 VDD2.n4 B 2.31155f
C26 VDD2.t3 B 0.223092f
C27 VDD2.t9 B 0.223092f
C28 VDD2.n5 B 1.98408f
C29 VDD2.n6 B 0.29732f
C30 VDD2.t1 B 0.223092f
C31 VDD2.t4 B 0.223092f
C32 VDD2.n7 B 1.98765f
C33 VN.n0 B 0.054719f
C34 VN.t1 B 1.06999f
C35 VN.n1 B 0.437821f
C36 VN.t3 B 1.09169f
C37 VN.t4 B 1.06999f
C38 VN.n2 B 0.437042f
C39 VN.n3 B 0.410998f
C40 VN.n4 B 0.249158f
C41 VN.n5 B 0.068303f
C42 VN.t7 B 1.06999f
C43 VN.n6 B 0.435798f
C44 VN.n7 B 0.009305f
C45 VN.t2 B 1.06999f
C46 VN.n8 B 0.422195f
C47 VN.n9 B 0.031779f
C48 VN.n10 B 0.054719f
C49 VN.t0 B 1.06999f
C50 VN.n11 B 0.437821f
C51 VN.t6 B 1.06999f
C52 VN.t5 B 1.09169f
C53 VN.t8 B 1.06999f
C54 VN.n12 B 0.437042f
C55 VN.n13 B 0.410998f
C56 VN.n14 B 0.249158f
C57 VN.n15 B 0.068303f
C58 VN.n16 B 0.435798f
C59 VN.n17 B 0.009305f
C60 VN.t9 B 1.06999f
C61 VN.n18 B 0.422195f
C62 VN.n19 B 1.78397f
C63 VDD1.t9 B 2.53545f
C64 VDD1.t4 B 0.223213f
C65 VDD1.t3 B 0.223213f
C66 VDD1.n0 B 1.98516f
C67 VDD1.n1 B 0.640042f
C68 VDD1.t6 B 2.53545f
C69 VDD1.t1 B 0.223213f
C70 VDD1.t2 B 0.223213f
C71 VDD1.n2 B 1.98515f
C72 VDD1.n3 B 0.634272f
C73 VDD1.t8 B 0.223213f
C74 VDD1.t5 B 0.223213f
C75 VDD1.n4 B 1.98875f
C76 VDD1.n5 B 1.93716f
C77 VDD1.t0 B 0.223213f
C78 VDD1.t7 B 0.223213f
C79 VDD1.n6 B 1.98515f
C80 VDD1.n7 B 2.31341f
C81 VTAIL.t6 B 0.2354f
C82 VTAIL.t7 B 0.2354f
C83 VTAIL.n0 B 2.01631f
C84 VTAIL.n1 B 0.394887f
C85 VTAIL.t13 B 2.56974f
C86 VTAIL.n2 B 0.498286f
C87 VTAIL.t11 B 0.2354f
C88 VTAIL.t12 B 0.2354f
C89 VTAIL.n3 B 2.01631f
C90 VTAIL.n4 B 0.410419f
C91 VTAIL.t16 B 0.2354f
C92 VTAIL.t9 B 0.2354f
C93 VTAIL.n5 B 2.01631f
C94 VTAIL.n6 B 1.66152f
C95 VTAIL.t0 B 0.2354f
C96 VTAIL.t3 B 0.2354f
C97 VTAIL.n7 B 2.01632f
C98 VTAIL.n8 B 1.66151f
C99 VTAIL.t19 B 0.2354f
C100 VTAIL.t4 B 0.2354f
C101 VTAIL.n9 B 2.01632f
C102 VTAIL.n10 B 0.410413f
C103 VTAIL.t8 B 2.56975f
C104 VTAIL.n11 B 0.498279f
C105 VTAIL.t10 B 0.2354f
C106 VTAIL.t17 B 0.2354f
C107 VTAIL.n12 B 2.01632f
C108 VTAIL.n13 B 0.409707f
C109 VTAIL.t18 B 0.2354f
C110 VTAIL.t15 B 0.2354f
C111 VTAIL.n14 B 2.01632f
C112 VTAIL.n15 B 0.410413f
C113 VTAIL.t14 B 2.56974f
C114 VTAIL.n16 B 1.67172f
C115 VTAIL.t5 B 2.56974f
C116 VTAIL.n17 B 1.67172f
C117 VTAIL.t2 B 0.2354f
C118 VTAIL.t1 B 0.2354f
C119 VTAIL.n18 B 2.01631f
C120 VTAIL.n19 B 0.346877f
C121 VP.n0 B 0.055448f
C122 VP.t7 B 1.08424f
C123 VP.n1 B 0.443653f
C124 VP.n2 B 0.055448f
C125 VP.n3 B 0.055448f
C126 VP.t2 B 1.08424f
C127 VP.t9 B 1.08424f
C128 VP.n4 B 0.069212f
C129 VP.t6 B 1.08424f
C130 VP.n5 B 0.252477f
C131 VP.t5 B 1.08424f
C132 VP.t0 B 1.10623f
C133 VP.n6 B 0.416472f
C134 VP.n7 B 0.442864f
C135 VP.n8 B 0.443653f
C136 VP.n9 B 0.441603f
C137 VP.n10 B 0.009429f
C138 VP.n11 B 0.427819f
C139 VP.n12 B 1.78049f
C140 VP.n13 B 1.81517f
C141 VP.t3 B 1.08424f
C142 VP.n14 B 0.427819f
C143 VP.n15 B 0.009429f
C144 VP.t8 B 1.08424f
C145 VP.n16 B 0.441603f
C146 VP.n17 B 0.069212f
C147 VP.n18 B 0.083107f
C148 VP.n19 B 0.069212f
C149 VP.t1 B 1.08424f
C150 VP.n20 B 0.441603f
C151 VP.n21 B 0.009429f
C152 VP.t4 B 1.08424f
C153 VP.n22 B 0.427819f
C154 VP.n23 B 0.032202f
.ends

