* NGSPICE file created from diff_pair_sample_0681.ext - technology: sky130A

.subckt diff_pair_sample_0681 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t14 VN.t0 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=6.4506 pd=33.86 as=2.7291 ps=16.87 w=16.54 l=3.48
X1 B.t20 B.t18 B.t19 B.t12 sky130_fd_pr__nfet_01v8 ad=6.4506 pd=33.86 as=0 ps=0 w=16.54 l=3.48
X2 VTAIL.t15 VP.t0 VDD1.t7 B.t21 sky130_fd_pr__nfet_01v8 ad=2.7291 pd=16.87 as=2.7291 ps=16.87 w=16.54 l=3.48
X3 VDD2.t1 VN.t1 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=2.7291 pd=16.87 as=6.4506 ps=33.86 w=16.54 l=3.48
X4 VTAIL.t12 VN.t2 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=6.4506 pd=33.86 as=2.7291 ps=16.87 w=16.54 l=3.48
X5 VTAIL.t3 VP.t1 VDD1.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=6.4506 pd=33.86 as=2.7291 ps=16.87 w=16.54 l=3.48
X6 VDD2.t7 VN.t3 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=2.7291 pd=16.87 as=2.7291 ps=16.87 w=16.54 l=3.48
X7 VDD1.t5 VP.t2 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.7291 pd=16.87 as=2.7291 ps=16.87 w=16.54 l=3.48
X8 VDD2.t6 VN.t4 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=2.7291 pd=16.87 as=2.7291 ps=16.87 w=16.54 l=3.48
X9 B.t17 B.t15 B.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=6.4506 pd=33.86 as=0 ps=0 w=16.54 l=3.48
X10 VTAIL.t4 VP.t3 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.7291 pd=16.87 as=2.7291 ps=16.87 w=16.54 l=3.48
X11 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=6.4506 pd=33.86 as=0 ps=0 w=16.54 l=3.48
X12 VTAIL.t9 VN.t5 VDD2.t5 B.t21 sky130_fd_pr__nfet_01v8 ad=2.7291 pd=16.87 as=2.7291 ps=16.87 w=16.54 l=3.48
X13 VTAIL.t8 VN.t6 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.7291 pd=16.87 as=2.7291 ps=16.87 w=16.54 l=3.48
X14 VDD2.t3 VN.t7 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7291 pd=16.87 as=6.4506 ps=33.86 w=16.54 l=3.48
X15 VDD1.t3 VP.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.7291 pd=16.87 as=2.7291 ps=16.87 w=16.54 l=3.48
X16 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=6.4506 pd=33.86 as=0 ps=0 w=16.54 l=3.48
X17 VTAIL.t0 VP.t5 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=6.4506 pd=33.86 as=2.7291 ps=16.87 w=16.54 l=3.48
X18 VDD1.t1 VP.t6 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.7291 pd=16.87 as=6.4506 ps=33.86 w=16.54 l=3.48
X19 VDD1.t0 VP.t7 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7291 pd=16.87 as=6.4506 ps=33.86 w=16.54 l=3.48
R0 VN.n68 VN.n67 161.3
R1 VN.n66 VN.n36 161.3
R2 VN.n65 VN.n64 161.3
R3 VN.n63 VN.n37 161.3
R4 VN.n62 VN.n61 161.3
R5 VN.n60 VN.n38 161.3
R6 VN.n59 VN.n58 161.3
R7 VN.n57 VN.n39 161.3
R8 VN.n56 VN.n55 161.3
R9 VN.n54 VN.n40 161.3
R10 VN.n53 VN.n52 161.3
R11 VN.n51 VN.n42 161.3
R12 VN.n50 VN.n49 161.3
R13 VN.n48 VN.n43 161.3
R14 VN.n47 VN.n46 161.3
R15 VN.n33 VN.n32 161.3
R16 VN.n31 VN.n1 161.3
R17 VN.n30 VN.n29 161.3
R18 VN.n28 VN.n2 161.3
R19 VN.n27 VN.n26 161.3
R20 VN.n25 VN.n3 161.3
R21 VN.n24 VN.n23 161.3
R22 VN.n22 VN.n4 161.3
R23 VN.n21 VN.n20 161.3
R24 VN.n18 VN.n5 161.3
R25 VN.n17 VN.n16 161.3
R26 VN.n15 VN.n6 161.3
R27 VN.n14 VN.n13 161.3
R28 VN.n12 VN.n7 161.3
R29 VN.n11 VN.n10 161.3
R30 VN.n45 VN.t7 148.103
R31 VN.n9 VN.t0 148.103
R32 VN.n8 VN.t3 114.544
R33 VN.n19 VN.t5 114.544
R34 VN.n0 VN.t1 114.544
R35 VN.n44 VN.t6 114.544
R36 VN.n41 VN.t4 114.544
R37 VN.n35 VN.t2 114.544
R38 VN.n34 VN.n0 79.6711
R39 VN.n69 VN.n35 79.6711
R40 VN VN.n69 58.7103
R41 VN.n26 VN.n2 56.5617
R42 VN.n61 VN.n37 56.5617
R43 VN.n9 VN.n8 54.9348
R44 VN.n45 VN.n44 54.9348
R45 VN.n13 VN.n6 40.577
R46 VN.n17 VN.n6 40.577
R47 VN.n49 VN.n42 40.577
R48 VN.n53 VN.n42 40.577
R49 VN.n12 VN.n11 24.5923
R50 VN.n13 VN.n12 24.5923
R51 VN.n18 VN.n17 24.5923
R52 VN.n20 VN.n18 24.5923
R53 VN.n24 VN.n4 24.5923
R54 VN.n25 VN.n24 24.5923
R55 VN.n26 VN.n25 24.5923
R56 VN.n30 VN.n2 24.5923
R57 VN.n31 VN.n30 24.5923
R58 VN.n32 VN.n31 24.5923
R59 VN.n49 VN.n48 24.5923
R60 VN.n48 VN.n47 24.5923
R61 VN.n61 VN.n60 24.5923
R62 VN.n60 VN.n59 24.5923
R63 VN.n59 VN.n39 24.5923
R64 VN.n55 VN.n54 24.5923
R65 VN.n54 VN.n53 24.5923
R66 VN.n67 VN.n66 24.5923
R67 VN.n66 VN.n65 24.5923
R68 VN.n65 VN.n37 24.5923
R69 VN.n11 VN.n8 19.9199
R70 VN.n20 VN.n19 19.9199
R71 VN.n47 VN.n44 19.9199
R72 VN.n55 VN.n41 19.9199
R73 VN.n32 VN.n0 10.575
R74 VN.n67 VN.n35 10.575
R75 VN.n19 VN.n4 4.67295
R76 VN.n41 VN.n39 4.67295
R77 VN.n10 VN.n9 3.12721
R78 VN.n46 VN.n45 3.12721
R79 VN.n69 VN.n68 0.354861
R80 VN.n34 VN.n33 0.354861
R81 VN VN.n34 0.267071
R82 VN.n68 VN.n36 0.189894
R83 VN.n64 VN.n36 0.189894
R84 VN.n64 VN.n63 0.189894
R85 VN.n63 VN.n62 0.189894
R86 VN.n62 VN.n38 0.189894
R87 VN.n58 VN.n38 0.189894
R88 VN.n58 VN.n57 0.189894
R89 VN.n57 VN.n56 0.189894
R90 VN.n56 VN.n40 0.189894
R91 VN.n52 VN.n40 0.189894
R92 VN.n52 VN.n51 0.189894
R93 VN.n51 VN.n50 0.189894
R94 VN.n50 VN.n43 0.189894
R95 VN.n46 VN.n43 0.189894
R96 VN.n10 VN.n7 0.189894
R97 VN.n14 VN.n7 0.189894
R98 VN.n15 VN.n14 0.189894
R99 VN.n16 VN.n15 0.189894
R100 VN.n16 VN.n5 0.189894
R101 VN.n21 VN.n5 0.189894
R102 VN.n22 VN.n21 0.189894
R103 VN.n23 VN.n22 0.189894
R104 VN.n23 VN.n3 0.189894
R105 VN.n27 VN.n3 0.189894
R106 VN.n28 VN.n27 0.189894
R107 VN.n29 VN.n28 0.189894
R108 VN.n29 VN.n1 0.189894
R109 VN.n33 VN.n1 0.189894
R110 VDD2.n2 VDD2.n1 64.2757
R111 VDD2.n2 VDD2.n0 64.2757
R112 VDD2 VDD2.n5 64.2729
R113 VDD2.n4 VDD2.n3 62.689
R114 VDD2.n4 VDD2.n2 52.7541
R115 VDD2 VDD2.n4 1.70093
R116 VDD2.n5 VDD2.t4 1.1976
R117 VDD2.n5 VDD2.t3 1.1976
R118 VDD2.n3 VDD2.t0 1.1976
R119 VDD2.n3 VDD2.t6 1.1976
R120 VDD2.n1 VDD2.t5 1.1976
R121 VDD2.n1 VDD2.t1 1.1976
R122 VDD2.n0 VDD2.t2 1.1976
R123 VDD2.n0 VDD2.t7 1.1976
R124 VTAIL.n11 VTAIL.t0 47.2073
R125 VTAIL.n10 VTAIL.t7 47.2073
R126 VTAIL.n7 VTAIL.t12 47.2073
R127 VTAIL.n14 VTAIL.t5 47.2071
R128 VTAIL.n15 VTAIL.t13 47.2071
R129 VTAIL.n2 VTAIL.t14 47.2071
R130 VTAIL.n3 VTAIL.t1 47.2071
R131 VTAIL.n6 VTAIL.t3 47.2071
R132 VTAIL.n13 VTAIL.n12 46.0102
R133 VTAIL.n9 VTAIL.n8 46.0102
R134 VTAIL.n1 VTAIL.n0 46.01
R135 VTAIL.n5 VTAIL.n4 46.01
R136 VTAIL.n15 VTAIL.n14 29.91
R137 VTAIL.n7 VTAIL.n6 29.91
R138 VTAIL.n9 VTAIL.n7 3.28498
R139 VTAIL.n10 VTAIL.n9 3.28498
R140 VTAIL.n13 VTAIL.n11 3.28498
R141 VTAIL.n14 VTAIL.n13 3.28498
R142 VTAIL.n6 VTAIL.n5 3.28498
R143 VTAIL.n5 VTAIL.n3 3.28498
R144 VTAIL.n2 VTAIL.n1 3.28498
R145 VTAIL VTAIL.n15 3.22679
R146 VTAIL.n0 VTAIL.t11 1.1976
R147 VTAIL.n0 VTAIL.t9 1.1976
R148 VTAIL.n4 VTAIL.t2 1.1976
R149 VTAIL.n4 VTAIL.t4 1.1976
R150 VTAIL.n12 VTAIL.t6 1.1976
R151 VTAIL.n12 VTAIL.t15 1.1976
R152 VTAIL.n8 VTAIL.t10 1.1976
R153 VTAIL.n8 VTAIL.t8 1.1976
R154 VTAIL.n11 VTAIL.n10 0.470328
R155 VTAIL.n3 VTAIL.n2 0.470328
R156 VTAIL VTAIL.n1 0.0586897
R157 B.n1124 B.n1123 585
R158 B.n418 B.n177 585
R159 B.n417 B.n416 585
R160 B.n415 B.n414 585
R161 B.n413 B.n412 585
R162 B.n411 B.n410 585
R163 B.n409 B.n408 585
R164 B.n407 B.n406 585
R165 B.n405 B.n404 585
R166 B.n403 B.n402 585
R167 B.n401 B.n400 585
R168 B.n399 B.n398 585
R169 B.n397 B.n396 585
R170 B.n395 B.n394 585
R171 B.n393 B.n392 585
R172 B.n391 B.n390 585
R173 B.n389 B.n388 585
R174 B.n387 B.n386 585
R175 B.n385 B.n384 585
R176 B.n383 B.n382 585
R177 B.n381 B.n380 585
R178 B.n379 B.n378 585
R179 B.n377 B.n376 585
R180 B.n375 B.n374 585
R181 B.n373 B.n372 585
R182 B.n371 B.n370 585
R183 B.n369 B.n368 585
R184 B.n367 B.n366 585
R185 B.n365 B.n364 585
R186 B.n363 B.n362 585
R187 B.n361 B.n360 585
R188 B.n359 B.n358 585
R189 B.n357 B.n356 585
R190 B.n355 B.n354 585
R191 B.n353 B.n352 585
R192 B.n351 B.n350 585
R193 B.n349 B.n348 585
R194 B.n347 B.n346 585
R195 B.n345 B.n344 585
R196 B.n343 B.n342 585
R197 B.n341 B.n340 585
R198 B.n339 B.n338 585
R199 B.n337 B.n336 585
R200 B.n335 B.n334 585
R201 B.n333 B.n332 585
R202 B.n331 B.n330 585
R203 B.n329 B.n328 585
R204 B.n327 B.n326 585
R205 B.n325 B.n324 585
R206 B.n323 B.n322 585
R207 B.n321 B.n320 585
R208 B.n319 B.n318 585
R209 B.n317 B.n316 585
R210 B.n315 B.n314 585
R211 B.n313 B.n312 585
R212 B.n310 B.n309 585
R213 B.n308 B.n307 585
R214 B.n306 B.n305 585
R215 B.n304 B.n303 585
R216 B.n302 B.n301 585
R217 B.n300 B.n299 585
R218 B.n298 B.n297 585
R219 B.n296 B.n295 585
R220 B.n294 B.n293 585
R221 B.n292 B.n291 585
R222 B.n289 B.n288 585
R223 B.n287 B.n286 585
R224 B.n285 B.n284 585
R225 B.n283 B.n282 585
R226 B.n281 B.n280 585
R227 B.n279 B.n278 585
R228 B.n277 B.n276 585
R229 B.n275 B.n274 585
R230 B.n273 B.n272 585
R231 B.n271 B.n270 585
R232 B.n269 B.n268 585
R233 B.n267 B.n266 585
R234 B.n265 B.n264 585
R235 B.n263 B.n262 585
R236 B.n261 B.n260 585
R237 B.n259 B.n258 585
R238 B.n257 B.n256 585
R239 B.n255 B.n254 585
R240 B.n253 B.n252 585
R241 B.n251 B.n250 585
R242 B.n249 B.n248 585
R243 B.n247 B.n246 585
R244 B.n245 B.n244 585
R245 B.n243 B.n242 585
R246 B.n241 B.n240 585
R247 B.n239 B.n238 585
R248 B.n237 B.n236 585
R249 B.n235 B.n234 585
R250 B.n233 B.n232 585
R251 B.n231 B.n230 585
R252 B.n229 B.n228 585
R253 B.n227 B.n226 585
R254 B.n225 B.n224 585
R255 B.n223 B.n222 585
R256 B.n221 B.n220 585
R257 B.n219 B.n218 585
R258 B.n217 B.n216 585
R259 B.n215 B.n214 585
R260 B.n213 B.n212 585
R261 B.n211 B.n210 585
R262 B.n209 B.n208 585
R263 B.n207 B.n206 585
R264 B.n205 B.n204 585
R265 B.n203 B.n202 585
R266 B.n201 B.n200 585
R267 B.n199 B.n198 585
R268 B.n197 B.n196 585
R269 B.n195 B.n194 585
R270 B.n193 B.n192 585
R271 B.n191 B.n190 585
R272 B.n189 B.n188 585
R273 B.n187 B.n186 585
R274 B.n185 B.n184 585
R275 B.n183 B.n182 585
R276 B.n116 B.n115 585
R277 B.n1122 B.n117 585
R278 B.n1127 B.n117 585
R279 B.n1121 B.n1120 585
R280 B.n1120 B.n113 585
R281 B.n1119 B.n112 585
R282 B.n1133 B.n112 585
R283 B.n1118 B.n111 585
R284 B.n1134 B.n111 585
R285 B.n1117 B.n110 585
R286 B.n1135 B.n110 585
R287 B.n1116 B.n1115 585
R288 B.n1115 B.n106 585
R289 B.n1114 B.n105 585
R290 B.n1141 B.n105 585
R291 B.n1113 B.n104 585
R292 B.n1142 B.n104 585
R293 B.n1112 B.n103 585
R294 B.n1143 B.n103 585
R295 B.n1111 B.n1110 585
R296 B.n1110 B.n99 585
R297 B.n1109 B.n98 585
R298 B.n1149 B.n98 585
R299 B.n1108 B.n97 585
R300 B.n1150 B.n97 585
R301 B.n1107 B.n96 585
R302 B.n1151 B.n96 585
R303 B.n1106 B.n1105 585
R304 B.n1105 B.n92 585
R305 B.n1104 B.n91 585
R306 B.n1157 B.n91 585
R307 B.n1103 B.n90 585
R308 B.n1158 B.n90 585
R309 B.n1102 B.n89 585
R310 B.n1159 B.n89 585
R311 B.n1101 B.n1100 585
R312 B.n1100 B.n85 585
R313 B.n1099 B.n84 585
R314 B.n1165 B.n84 585
R315 B.n1098 B.n83 585
R316 B.n1166 B.n83 585
R317 B.n1097 B.n82 585
R318 B.n1167 B.n82 585
R319 B.n1096 B.n1095 585
R320 B.n1095 B.n78 585
R321 B.n1094 B.n77 585
R322 B.n1173 B.n77 585
R323 B.n1093 B.n76 585
R324 B.n1174 B.n76 585
R325 B.n1092 B.n75 585
R326 B.n1175 B.n75 585
R327 B.n1091 B.n1090 585
R328 B.n1090 B.n71 585
R329 B.n1089 B.n70 585
R330 B.n1181 B.n70 585
R331 B.n1088 B.n69 585
R332 B.n1182 B.n69 585
R333 B.n1087 B.n68 585
R334 B.n1183 B.n68 585
R335 B.n1086 B.n1085 585
R336 B.n1085 B.n64 585
R337 B.n1084 B.n63 585
R338 B.n1189 B.n63 585
R339 B.n1083 B.n62 585
R340 B.n1190 B.n62 585
R341 B.n1082 B.n61 585
R342 B.n1191 B.n61 585
R343 B.n1081 B.n1080 585
R344 B.n1080 B.n57 585
R345 B.n1079 B.n56 585
R346 B.n1197 B.n56 585
R347 B.n1078 B.n55 585
R348 B.n1198 B.n55 585
R349 B.n1077 B.n54 585
R350 B.n1199 B.n54 585
R351 B.n1076 B.n1075 585
R352 B.n1075 B.n50 585
R353 B.n1074 B.n49 585
R354 B.n1205 B.n49 585
R355 B.n1073 B.n48 585
R356 B.n1206 B.n48 585
R357 B.n1072 B.n47 585
R358 B.n1207 B.n47 585
R359 B.n1071 B.n1070 585
R360 B.n1070 B.n43 585
R361 B.n1069 B.n42 585
R362 B.n1213 B.n42 585
R363 B.n1068 B.n41 585
R364 B.n1214 B.n41 585
R365 B.n1067 B.n40 585
R366 B.n1215 B.n40 585
R367 B.n1066 B.n1065 585
R368 B.n1065 B.n39 585
R369 B.n1064 B.n35 585
R370 B.n1221 B.n35 585
R371 B.n1063 B.n34 585
R372 B.n1222 B.n34 585
R373 B.n1062 B.n33 585
R374 B.n1223 B.n33 585
R375 B.n1061 B.n1060 585
R376 B.n1060 B.n29 585
R377 B.n1059 B.n28 585
R378 B.n1229 B.n28 585
R379 B.n1058 B.n27 585
R380 B.n1230 B.n27 585
R381 B.n1057 B.n26 585
R382 B.n1231 B.n26 585
R383 B.n1056 B.n1055 585
R384 B.n1055 B.n22 585
R385 B.n1054 B.n21 585
R386 B.n1237 B.n21 585
R387 B.n1053 B.n20 585
R388 B.n1238 B.n20 585
R389 B.n1052 B.n19 585
R390 B.n1239 B.n19 585
R391 B.n1051 B.n1050 585
R392 B.n1050 B.n15 585
R393 B.n1049 B.n14 585
R394 B.n1245 B.n14 585
R395 B.n1048 B.n13 585
R396 B.n1246 B.n13 585
R397 B.n1047 B.n12 585
R398 B.n1247 B.n12 585
R399 B.n1046 B.n1045 585
R400 B.n1045 B.n8 585
R401 B.n1044 B.n7 585
R402 B.n1253 B.n7 585
R403 B.n1043 B.n6 585
R404 B.n1254 B.n6 585
R405 B.n1042 B.n5 585
R406 B.n1255 B.n5 585
R407 B.n1041 B.n1040 585
R408 B.n1040 B.n4 585
R409 B.n1039 B.n419 585
R410 B.n1039 B.n1038 585
R411 B.n1029 B.n420 585
R412 B.n421 B.n420 585
R413 B.n1031 B.n1030 585
R414 B.n1032 B.n1031 585
R415 B.n1028 B.n426 585
R416 B.n426 B.n425 585
R417 B.n1027 B.n1026 585
R418 B.n1026 B.n1025 585
R419 B.n428 B.n427 585
R420 B.n429 B.n428 585
R421 B.n1018 B.n1017 585
R422 B.n1019 B.n1018 585
R423 B.n1016 B.n434 585
R424 B.n434 B.n433 585
R425 B.n1015 B.n1014 585
R426 B.n1014 B.n1013 585
R427 B.n436 B.n435 585
R428 B.n437 B.n436 585
R429 B.n1006 B.n1005 585
R430 B.n1007 B.n1006 585
R431 B.n1004 B.n442 585
R432 B.n442 B.n441 585
R433 B.n1003 B.n1002 585
R434 B.n1002 B.n1001 585
R435 B.n444 B.n443 585
R436 B.n445 B.n444 585
R437 B.n994 B.n993 585
R438 B.n995 B.n994 585
R439 B.n992 B.n450 585
R440 B.n450 B.n449 585
R441 B.n991 B.n990 585
R442 B.n990 B.n989 585
R443 B.n452 B.n451 585
R444 B.n982 B.n452 585
R445 B.n981 B.n980 585
R446 B.n983 B.n981 585
R447 B.n979 B.n457 585
R448 B.n457 B.n456 585
R449 B.n978 B.n977 585
R450 B.n977 B.n976 585
R451 B.n459 B.n458 585
R452 B.n460 B.n459 585
R453 B.n969 B.n968 585
R454 B.n970 B.n969 585
R455 B.n967 B.n465 585
R456 B.n465 B.n464 585
R457 B.n966 B.n965 585
R458 B.n965 B.n964 585
R459 B.n467 B.n466 585
R460 B.n468 B.n467 585
R461 B.n957 B.n956 585
R462 B.n958 B.n957 585
R463 B.n955 B.n473 585
R464 B.n473 B.n472 585
R465 B.n954 B.n953 585
R466 B.n953 B.n952 585
R467 B.n475 B.n474 585
R468 B.n476 B.n475 585
R469 B.n945 B.n944 585
R470 B.n946 B.n945 585
R471 B.n943 B.n481 585
R472 B.n481 B.n480 585
R473 B.n942 B.n941 585
R474 B.n941 B.n940 585
R475 B.n483 B.n482 585
R476 B.n484 B.n483 585
R477 B.n933 B.n932 585
R478 B.n934 B.n933 585
R479 B.n931 B.n489 585
R480 B.n489 B.n488 585
R481 B.n930 B.n929 585
R482 B.n929 B.n928 585
R483 B.n491 B.n490 585
R484 B.n492 B.n491 585
R485 B.n921 B.n920 585
R486 B.n922 B.n921 585
R487 B.n919 B.n496 585
R488 B.n500 B.n496 585
R489 B.n918 B.n917 585
R490 B.n917 B.n916 585
R491 B.n498 B.n497 585
R492 B.n499 B.n498 585
R493 B.n909 B.n908 585
R494 B.n910 B.n909 585
R495 B.n907 B.n505 585
R496 B.n505 B.n504 585
R497 B.n906 B.n905 585
R498 B.n905 B.n904 585
R499 B.n507 B.n506 585
R500 B.n508 B.n507 585
R501 B.n897 B.n896 585
R502 B.n898 B.n897 585
R503 B.n895 B.n513 585
R504 B.n513 B.n512 585
R505 B.n894 B.n893 585
R506 B.n893 B.n892 585
R507 B.n515 B.n514 585
R508 B.n516 B.n515 585
R509 B.n885 B.n884 585
R510 B.n886 B.n885 585
R511 B.n883 B.n521 585
R512 B.n521 B.n520 585
R513 B.n882 B.n881 585
R514 B.n881 B.n880 585
R515 B.n523 B.n522 585
R516 B.n524 B.n523 585
R517 B.n873 B.n872 585
R518 B.n874 B.n873 585
R519 B.n871 B.n529 585
R520 B.n529 B.n528 585
R521 B.n870 B.n869 585
R522 B.n869 B.n868 585
R523 B.n531 B.n530 585
R524 B.n532 B.n531 585
R525 B.n861 B.n860 585
R526 B.n862 B.n861 585
R527 B.n859 B.n537 585
R528 B.n537 B.n536 585
R529 B.n858 B.n857 585
R530 B.n857 B.n856 585
R531 B.n539 B.n538 585
R532 B.n540 B.n539 585
R533 B.n849 B.n848 585
R534 B.n850 B.n849 585
R535 B.n543 B.n542 585
R536 B.n612 B.n611 585
R537 B.n613 B.n609 585
R538 B.n609 B.n544 585
R539 B.n615 B.n614 585
R540 B.n617 B.n608 585
R541 B.n620 B.n619 585
R542 B.n621 B.n607 585
R543 B.n623 B.n622 585
R544 B.n625 B.n606 585
R545 B.n628 B.n627 585
R546 B.n629 B.n605 585
R547 B.n631 B.n630 585
R548 B.n633 B.n604 585
R549 B.n636 B.n635 585
R550 B.n637 B.n603 585
R551 B.n639 B.n638 585
R552 B.n641 B.n602 585
R553 B.n644 B.n643 585
R554 B.n645 B.n601 585
R555 B.n647 B.n646 585
R556 B.n649 B.n600 585
R557 B.n652 B.n651 585
R558 B.n653 B.n599 585
R559 B.n655 B.n654 585
R560 B.n657 B.n598 585
R561 B.n660 B.n659 585
R562 B.n661 B.n597 585
R563 B.n663 B.n662 585
R564 B.n665 B.n596 585
R565 B.n668 B.n667 585
R566 B.n669 B.n595 585
R567 B.n671 B.n670 585
R568 B.n673 B.n594 585
R569 B.n676 B.n675 585
R570 B.n677 B.n593 585
R571 B.n679 B.n678 585
R572 B.n681 B.n592 585
R573 B.n684 B.n683 585
R574 B.n685 B.n591 585
R575 B.n687 B.n686 585
R576 B.n689 B.n590 585
R577 B.n692 B.n691 585
R578 B.n693 B.n589 585
R579 B.n695 B.n694 585
R580 B.n697 B.n588 585
R581 B.n700 B.n699 585
R582 B.n701 B.n587 585
R583 B.n703 B.n702 585
R584 B.n705 B.n586 585
R585 B.n708 B.n707 585
R586 B.n709 B.n585 585
R587 B.n711 B.n710 585
R588 B.n713 B.n584 585
R589 B.n716 B.n715 585
R590 B.n717 B.n581 585
R591 B.n720 B.n719 585
R592 B.n722 B.n580 585
R593 B.n725 B.n724 585
R594 B.n726 B.n579 585
R595 B.n728 B.n727 585
R596 B.n730 B.n578 585
R597 B.n733 B.n732 585
R598 B.n734 B.n577 585
R599 B.n736 B.n735 585
R600 B.n738 B.n576 585
R601 B.n741 B.n740 585
R602 B.n742 B.n572 585
R603 B.n744 B.n743 585
R604 B.n746 B.n571 585
R605 B.n749 B.n748 585
R606 B.n750 B.n570 585
R607 B.n752 B.n751 585
R608 B.n754 B.n569 585
R609 B.n757 B.n756 585
R610 B.n758 B.n568 585
R611 B.n760 B.n759 585
R612 B.n762 B.n567 585
R613 B.n765 B.n764 585
R614 B.n766 B.n566 585
R615 B.n768 B.n767 585
R616 B.n770 B.n565 585
R617 B.n773 B.n772 585
R618 B.n774 B.n564 585
R619 B.n776 B.n775 585
R620 B.n778 B.n563 585
R621 B.n781 B.n780 585
R622 B.n782 B.n562 585
R623 B.n784 B.n783 585
R624 B.n786 B.n561 585
R625 B.n789 B.n788 585
R626 B.n790 B.n560 585
R627 B.n792 B.n791 585
R628 B.n794 B.n559 585
R629 B.n797 B.n796 585
R630 B.n798 B.n558 585
R631 B.n800 B.n799 585
R632 B.n802 B.n557 585
R633 B.n805 B.n804 585
R634 B.n806 B.n556 585
R635 B.n808 B.n807 585
R636 B.n810 B.n555 585
R637 B.n813 B.n812 585
R638 B.n814 B.n554 585
R639 B.n816 B.n815 585
R640 B.n818 B.n553 585
R641 B.n821 B.n820 585
R642 B.n822 B.n552 585
R643 B.n824 B.n823 585
R644 B.n826 B.n551 585
R645 B.n829 B.n828 585
R646 B.n830 B.n550 585
R647 B.n832 B.n831 585
R648 B.n834 B.n549 585
R649 B.n837 B.n836 585
R650 B.n838 B.n548 585
R651 B.n840 B.n839 585
R652 B.n842 B.n547 585
R653 B.n843 B.n546 585
R654 B.n846 B.n845 585
R655 B.n847 B.n545 585
R656 B.n545 B.n544 585
R657 B.n852 B.n851 585
R658 B.n851 B.n850 585
R659 B.n853 B.n541 585
R660 B.n541 B.n540 585
R661 B.n855 B.n854 585
R662 B.n856 B.n855 585
R663 B.n535 B.n534 585
R664 B.n536 B.n535 585
R665 B.n864 B.n863 585
R666 B.n863 B.n862 585
R667 B.n865 B.n533 585
R668 B.n533 B.n532 585
R669 B.n867 B.n866 585
R670 B.n868 B.n867 585
R671 B.n527 B.n526 585
R672 B.n528 B.n527 585
R673 B.n876 B.n875 585
R674 B.n875 B.n874 585
R675 B.n877 B.n525 585
R676 B.n525 B.n524 585
R677 B.n879 B.n878 585
R678 B.n880 B.n879 585
R679 B.n519 B.n518 585
R680 B.n520 B.n519 585
R681 B.n888 B.n887 585
R682 B.n887 B.n886 585
R683 B.n889 B.n517 585
R684 B.n517 B.n516 585
R685 B.n891 B.n890 585
R686 B.n892 B.n891 585
R687 B.n511 B.n510 585
R688 B.n512 B.n511 585
R689 B.n900 B.n899 585
R690 B.n899 B.n898 585
R691 B.n901 B.n509 585
R692 B.n509 B.n508 585
R693 B.n903 B.n902 585
R694 B.n904 B.n903 585
R695 B.n503 B.n502 585
R696 B.n504 B.n503 585
R697 B.n912 B.n911 585
R698 B.n911 B.n910 585
R699 B.n913 B.n501 585
R700 B.n501 B.n499 585
R701 B.n915 B.n914 585
R702 B.n916 B.n915 585
R703 B.n495 B.n494 585
R704 B.n500 B.n495 585
R705 B.n924 B.n923 585
R706 B.n923 B.n922 585
R707 B.n925 B.n493 585
R708 B.n493 B.n492 585
R709 B.n927 B.n926 585
R710 B.n928 B.n927 585
R711 B.n487 B.n486 585
R712 B.n488 B.n487 585
R713 B.n936 B.n935 585
R714 B.n935 B.n934 585
R715 B.n937 B.n485 585
R716 B.n485 B.n484 585
R717 B.n939 B.n938 585
R718 B.n940 B.n939 585
R719 B.n479 B.n478 585
R720 B.n480 B.n479 585
R721 B.n948 B.n947 585
R722 B.n947 B.n946 585
R723 B.n949 B.n477 585
R724 B.n477 B.n476 585
R725 B.n951 B.n950 585
R726 B.n952 B.n951 585
R727 B.n471 B.n470 585
R728 B.n472 B.n471 585
R729 B.n960 B.n959 585
R730 B.n959 B.n958 585
R731 B.n961 B.n469 585
R732 B.n469 B.n468 585
R733 B.n963 B.n962 585
R734 B.n964 B.n963 585
R735 B.n463 B.n462 585
R736 B.n464 B.n463 585
R737 B.n972 B.n971 585
R738 B.n971 B.n970 585
R739 B.n973 B.n461 585
R740 B.n461 B.n460 585
R741 B.n975 B.n974 585
R742 B.n976 B.n975 585
R743 B.n455 B.n454 585
R744 B.n456 B.n455 585
R745 B.n985 B.n984 585
R746 B.n984 B.n983 585
R747 B.n986 B.n453 585
R748 B.n982 B.n453 585
R749 B.n988 B.n987 585
R750 B.n989 B.n988 585
R751 B.n448 B.n447 585
R752 B.n449 B.n448 585
R753 B.n997 B.n996 585
R754 B.n996 B.n995 585
R755 B.n998 B.n446 585
R756 B.n446 B.n445 585
R757 B.n1000 B.n999 585
R758 B.n1001 B.n1000 585
R759 B.n440 B.n439 585
R760 B.n441 B.n440 585
R761 B.n1009 B.n1008 585
R762 B.n1008 B.n1007 585
R763 B.n1010 B.n438 585
R764 B.n438 B.n437 585
R765 B.n1012 B.n1011 585
R766 B.n1013 B.n1012 585
R767 B.n432 B.n431 585
R768 B.n433 B.n432 585
R769 B.n1021 B.n1020 585
R770 B.n1020 B.n1019 585
R771 B.n1022 B.n430 585
R772 B.n430 B.n429 585
R773 B.n1024 B.n1023 585
R774 B.n1025 B.n1024 585
R775 B.n424 B.n423 585
R776 B.n425 B.n424 585
R777 B.n1034 B.n1033 585
R778 B.n1033 B.n1032 585
R779 B.n1035 B.n422 585
R780 B.n422 B.n421 585
R781 B.n1037 B.n1036 585
R782 B.n1038 B.n1037 585
R783 B.n2 B.n0 585
R784 B.n4 B.n2 585
R785 B.n3 B.n1 585
R786 B.n1254 B.n3 585
R787 B.n1252 B.n1251 585
R788 B.n1253 B.n1252 585
R789 B.n1250 B.n9 585
R790 B.n9 B.n8 585
R791 B.n1249 B.n1248 585
R792 B.n1248 B.n1247 585
R793 B.n11 B.n10 585
R794 B.n1246 B.n11 585
R795 B.n1244 B.n1243 585
R796 B.n1245 B.n1244 585
R797 B.n1242 B.n16 585
R798 B.n16 B.n15 585
R799 B.n1241 B.n1240 585
R800 B.n1240 B.n1239 585
R801 B.n18 B.n17 585
R802 B.n1238 B.n18 585
R803 B.n1236 B.n1235 585
R804 B.n1237 B.n1236 585
R805 B.n1234 B.n23 585
R806 B.n23 B.n22 585
R807 B.n1233 B.n1232 585
R808 B.n1232 B.n1231 585
R809 B.n25 B.n24 585
R810 B.n1230 B.n25 585
R811 B.n1228 B.n1227 585
R812 B.n1229 B.n1228 585
R813 B.n1226 B.n30 585
R814 B.n30 B.n29 585
R815 B.n1225 B.n1224 585
R816 B.n1224 B.n1223 585
R817 B.n32 B.n31 585
R818 B.n1222 B.n32 585
R819 B.n1220 B.n1219 585
R820 B.n1221 B.n1220 585
R821 B.n1218 B.n36 585
R822 B.n39 B.n36 585
R823 B.n1217 B.n1216 585
R824 B.n1216 B.n1215 585
R825 B.n38 B.n37 585
R826 B.n1214 B.n38 585
R827 B.n1212 B.n1211 585
R828 B.n1213 B.n1212 585
R829 B.n1210 B.n44 585
R830 B.n44 B.n43 585
R831 B.n1209 B.n1208 585
R832 B.n1208 B.n1207 585
R833 B.n46 B.n45 585
R834 B.n1206 B.n46 585
R835 B.n1204 B.n1203 585
R836 B.n1205 B.n1204 585
R837 B.n1202 B.n51 585
R838 B.n51 B.n50 585
R839 B.n1201 B.n1200 585
R840 B.n1200 B.n1199 585
R841 B.n53 B.n52 585
R842 B.n1198 B.n53 585
R843 B.n1196 B.n1195 585
R844 B.n1197 B.n1196 585
R845 B.n1194 B.n58 585
R846 B.n58 B.n57 585
R847 B.n1193 B.n1192 585
R848 B.n1192 B.n1191 585
R849 B.n60 B.n59 585
R850 B.n1190 B.n60 585
R851 B.n1188 B.n1187 585
R852 B.n1189 B.n1188 585
R853 B.n1186 B.n65 585
R854 B.n65 B.n64 585
R855 B.n1185 B.n1184 585
R856 B.n1184 B.n1183 585
R857 B.n67 B.n66 585
R858 B.n1182 B.n67 585
R859 B.n1180 B.n1179 585
R860 B.n1181 B.n1180 585
R861 B.n1178 B.n72 585
R862 B.n72 B.n71 585
R863 B.n1177 B.n1176 585
R864 B.n1176 B.n1175 585
R865 B.n74 B.n73 585
R866 B.n1174 B.n74 585
R867 B.n1172 B.n1171 585
R868 B.n1173 B.n1172 585
R869 B.n1170 B.n79 585
R870 B.n79 B.n78 585
R871 B.n1169 B.n1168 585
R872 B.n1168 B.n1167 585
R873 B.n81 B.n80 585
R874 B.n1166 B.n81 585
R875 B.n1164 B.n1163 585
R876 B.n1165 B.n1164 585
R877 B.n1162 B.n86 585
R878 B.n86 B.n85 585
R879 B.n1161 B.n1160 585
R880 B.n1160 B.n1159 585
R881 B.n88 B.n87 585
R882 B.n1158 B.n88 585
R883 B.n1156 B.n1155 585
R884 B.n1157 B.n1156 585
R885 B.n1154 B.n93 585
R886 B.n93 B.n92 585
R887 B.n1153 B.n1152 585
R888 B.n1152 B.n1151 585
R889 B.n95 B.n94 585
R890 B.n1150 B.n95 585
R891 B.n1148 B.n1147 585
R892 B.n1149 B.n1148 585
R893 B.n1146 B.n100 585
R894 B.n100 B.n99 585
R895 B.n1145 B.n1144 585
R896 B.n1144 B.n1143 585
R897 B.n102 B.n101 585
R898 B.n1142 B.n102 585
R899 B.n1140 B.n1139 585
R900 B.n1141 B.n1140 585
R901 B.n1138 B.n107 585
R902 B.n107 B.n106 585
R903 B.n1137 B.n1136 585
R904 B.n1136 B.n1135 585
R905 B.n109 B.n108 585
R906 B.n1134 B.n109 585
R907 B.n1132 B.n1131 585
R908 B.n1133 B.n1132 585
R909 B.n1130 B.n114 585
R910 B.n114 B.n113 585
R911 B.n1129 B.n1128 585
R912 B.n1128 B.n1127 585
R913 B.n1257 B.n1256 585
R914 B.n1256 B.n1255 585
R915 B.n851 B.n543 482.89
R916 B.n1128 B.n116 482.89
R917 B.n849 B.n545 482.89
R918 B.n1124 B.n117 482.89
R919 B.n573 B.t7 323.62
R920 B.n582 B.t15 323.62
R921 B.n180 B.t18 323.62
R922 B.n178 B.t11 323.62
R923 B.n1126 B.n1125 256.663
R924 B.n1126 B.n176 256.663
R925 B.n1126 B.n175 256.663
R926 B.n1126 B.n174 256.663
R927 B.n1126 B.n173 256.663
R928 B.n1126 B.n172 256.663
R929 B.n1126 B.n171 256.663
R930 B.n1126 B.n170 256.663
R931 B.n1126 B.n169 256.663
R932 B.n1126 B.n168 256.663
R933 B.n1126 B.n167 256.663
R934 B.n1126 B.n166 256.663
R935 B.n1126 B.n165 256.663
R936 B.n1126 B.n164 256.663
R937 B.n1126 B.n163 256.663
R938 B.n1126 B.n162 256.663
R939 B.n1126 B.n161 256.663
R940 B.n1126 B.n160 256.663
R941 B.n1126 B.n159 256.663
R942 B.n1126 B.n158 256.663
R943 B.n1126 B.n157 256.663
R944 B.n1126 B.n156 256.663
R945 B.n1126 B.n155 256.663
R946 B.n1126 B.n154 256.663
R947 B.n1126 B.n153 256.663
R948 B.n1126 B.n152 256.663
R949 B.n1126 B.n151 256.663
R950 B.n1126 B.n150 256.663
R951 B.n1126 B.n149 256.663
R952 B.n1126 B.n148 256.663
R953 B.n1126 B.n147 256.663
R954 B.n1126 B.n146 256.663
R955 B.n1126 B.n145 256.663
R956 B.n1126 B.n144 256.663
R957 B.n1126 B.n143 256.663
R958 B.n1126 B.n142 256.663
R959 B.n1126 B.n141 256.663
R960 B.n1126 B.n140 256.663
R961 B.n1126 B.n139 256.663
R962 B.n1126 B.n138 256.663
R963 B.n1126 B.n137 256.663
R964 B.n1126 B.n136 256.663
R965 B.n1126 B.n135 256.663
R966 B.n1126 B.n134 256.663
R967 B.n1126 B.n133 256.663
R968 B.n1126 B.n132 256.663
R969 B.n1126 B.n131 256.663
R970 B.n1126 B.n130 256.663
R971 B.n1126 B.n129 256.663
R972 B.n1126 B.n128 256.663
R973 B.n1126 B.n127 256.663
R974 B.n1126 B.n126 256.663
R975 B.n1126 B.n125 256.663
R976 B.n1126 B.n124 256.663
R977 B.n1126 B.n123 256.663
R978 B.n1126 B.n122 256.663
R979 B.n1126 B.n121 256.663
R980 B.n1126 B.n120 256.663
R981 B.n1126 B.n119 256.663
R982 B.n1126 B.n118 256.663
R983 B.n610 B.n544 256.663
R984 B.n616 B.n544 256.663
R985 B.n618 B.n544 256.663
R986 B.n624 B.n544 256.663
R987 B.n626 B.n544 256.663
R988 B.n632 B.n544 256.663
R989 B.n634 B.n544 256.663
R990 B.n640 B.n544 256.663
R991 B.n642 B.n544 256.663
R992 B.n648 B.n544 256.663
R993 B.n650 B.n544 256.663
R994 B.n656 B.n544 256.663
R995 B.n658 B.n544 256.663
R996 B.n664 B.n544 256.663
R997 B.n666 B.n544 256.663
R998 B.n672 B.n544 256.663
R999 B.n674 B.n544 256.663
R1000 B.n680 B.n544 256.663
R1001 B.n682 B.n544 256.663
R1002 B.n688 B.n544 256.663
R1003 B.n690 B.n544 256.663
R1004 B.n696 B.n544 256.663
R1005 B.n698 B.n544 256.663
R1006 B.n704 B.n544 256.663
R1007 B.n706 B.n544 256.663
R1008 B.n712 B.n544 256.663
R1009 B.n714 B.n544 256.663
R1010 B.n721 B.n544 256.663
R1011 B.n723 B.n544 256.663
R1012 B.n729 B.n544 256.663
R1013 B.n731 B.n544 256.663
R1014 B.n737 B.n544 256.663
R1015 B.n739 B.n544 256.663
R1016 B.n745 B.n544 256.663
R1017 B.n747 B.n544 256.663
R1018 B.n753 B.n544 256.663
R1019 B.n755 B.n544 256.663
R1020 B.n761 B.n544 256.663
R1021 B.n763 B.n544 256.663
R1022 B.n769 B.n544 256.663
R1023 B.n771 B.n544 256.663
R1024 B.n777 B.n544 256.663
R1025 B.n779 B.n544 256.663
R1026 B.n785 B.n544 256.663
R1027 B.n787 B.n544 256.663
R1028 B.n793 B.n544 256.663
R1029 B.n795 B.n544 256.663
R1030 B.n801 B.n544 256.663
R1031 B.n803 B.n544 256.663
R1032 B.n809 B.n544 256.663
R1033 B.n811 B.n544 256.663
R1034 B.n817 B.n544 256.663
R1035 B.n819 B.n544 256.663
R1036 B.n825 B.n544 256.663
R1037 B.n827 B.n544 256.663
R1038 B.n833 B.n544 256.663
R1039 B.n835 B.n544 256.663
R1040 B.n841 B.n544 256.663
R1041 B.n844 B.n544 256.663
R1042 B.n851 B.n541 163.367
R1043 B.n855 B.n541 163.367
R1044 B.n855 B.n535 163.367
R1045 B.n863 B.n535 163.367
R1046 B.n863 B.n533 163.367
R1047 B.n867 B.n533 163.367
R1048 B.n867 B.n527 163.367
R1049 B.n875 B.n527 163.367
R1050 B.n875 B.n525 163.367
R1051 B.n879 B.n525 163.367
R1052 B.n879 B.n519 163.367
R1053 B.n887 B.n519 163.367
R1054 B.n887 B.n517 163.367
R1055 B.n891 B.n517 163.367
R1056 B.n891 B.n511 163.367
R1057 B.n899 B.n511 163.367
R1058 B.n899 B.n509 163.367
R1059 B.n903 B.n509 163.367
R1060 B.n903 B.n503 163.367
R1061 B.n911 B.n503 163.367
R1062 B.n911 B.n501 163.367
R1063 B.n915 B.n501 163.367
R1064 B.n915 B.n495 163.367
R1065 B.n923 B.n495 163.367
R1066 B.n923 B.n493 163.367
R1067 B.n927 B.n493 163.367
R1068 B.n927 B.n487 163.367
R1069 B.n935 B.n487 163.367
R1070 B.n935 B.n485 163.367
R1071 B.n939 B.n485 163.367
R1072 B.n939 B.n479 163.367
R1073 B.n947 B.n479 163.367
R1074 B.n947 B.n477 163.367
R1075 B.n951 B.n477 163.367
R1076 B.n951 B.n471 163.367
R1077 B.n959 B.n471 163.367
R1078 B.n959 B.n469 163.367
R1079 B.n963 B.n469 163.367
R1080 B.n963 B.n463 163.367
R1081 B.n971 B.n463 163.367
R1082 B.n971 B.n461 163.367
R1083 B.n975 B.n461 163.367
R1084 B.n975 B.n455 163.367
R1085 B.n984 B.n455 163.367
R1086 B.n984 B.n453 163.367
R1087 B.n988 B.n453 163.367
R1088 B.n988 B.n448 163.367
R1089 B.n996 B.n448 163.367
R1090 B.n996 B.n446 163.367
R1091 B.n1000 B.n446 163.367
R1092 B.n1000 B.n440 163.367
R1093 B.n1008 B.n440 163.367
R1094 B.n1008 B.n438 163.367
R1095 B.n1012 B.n438 163.367
R1096 B.n1012 B.n432 163.367
R1097 B.n1020 B.n432 163.367
R1098 B.n1020 B.n430 163.367
R1099 B.n1024 B.n430 163.367
R1100 B.n1024 B.n424 163.367
R1101 B.n1033 B.n424 163.367
R1102 B.n1033 B.n422 163.367
R1103 B.n1037 B.n422 163.367
R1104 B.n1037 B.n2 163.367
R1105 B.n1256 B.n2 163.367
R1106 B.n1256 B.n3 163.367
R1107 B.n1252 B.n3 163.367
R1108 B.n1252 B.n9 163.367
R1109 B.n1248 B.n9 163.367
R1110 B.n1248 B.n11 163.367
R1111 B.n1244 B.n11 163.367
R1112 B.n1244 B.n16 163.367
R1113 B.n1240 B.n16 163.367
R1114 B.n1240 B.n18 163.367
R1115 B.n1236 B.n18 163.367
R1116 B.n1236 B.n23 163.367
R1117 B.n1232 B.n23 163.367
R1118 B.n1232 B.n25 163.367
R1119 B.n1228 B.n25 163.367
R1120 B.n1228 B.n30 163.367
R1121 B.n1224 B.n30 163.367
R1122 B.n1224 B.n32 163.367
R1123 B.n1220 B.n32 163.367
R1124 B.n1220 B.n36 163.367
R1125 B.n1216 B.n36 163.367
R1126 B.n1216 B.n38 163.367
R1127 B.n1212 B.n38 163.367
R1128 B.n1212 B.n44 163.367
R1129 B.n1208 B.n44 163.367
R1130 B.n1208 B.n46 163.367
R1131 B.n1204 B.n46 163.367
R1132 B.n1204 B.n51 163.367
R1133 B.n1200 B.n51 163.367
R1134 B.n1200 B.n53 163.367
R1135 B.n1196 B.n53 163.367
R1136 B.n1196 B.n58 163.367
R1137 B.n1192 B.n58 163.367
R1138 B.n1192 B.n60 163.367
R1139 B.n1188 B.n60 163.367
R1140 B.n1188 B.n65 163.367
R1141 B.n1184 B.n65 163.367
R1142 B.n1184 B.n67 163.367
R1143 B.n1180 B.n67 163.367
R1144 B.n1180 B.n72 163.367
R1145 B.n1176 B.n72 163.367
R1146 B.n1176 B.n74 163.367
R1147 B.n1172 B.n74 163.367
R1148 B.n1172 B.n79 163.367
R1149 B.n1168 B.n79 163.367
R1150 B.n1168 B.n81 163.367
R1151 B.n1164 B.n81 163.367
R1152 B.n1164 B.n86 163.367
R1153 B.n1160 B.n86 163.367
R1154 B.n1160 B.n88 163.367
R1155 B.n1156 B.n88 163.367
R1156 B.n1156 B.n93 163.367
R1157 B.n1152 B.n93 163.367
R1158 B.n1152 B.n95 163.367
R1159 B.n1148 B.n95 163.367
R1160 B.n1148 B.n100 163.367
R1161 B.n1144 B.n100 163.367
R1162 B.n1144 B.n102 163.367
R1163 B.n1140 B.n102 163.367
R1164 B.n1140 B.n107 163.367
R1165 B.n1136 B.n107 163.367
R1166 B.n1136 B.n109 163.367
R1167 B.n1132 B.n109 163.367
R1168 B.n1132 B.n114 163.367
R1169 B.n1128 B.n114 163.367
R1170 B.n611 B.n609 163.367
R1171 B.n615 B.n609 163.367
R1172 B.n619 B.n617 163.367
R1173 B.n623 B.n607 163.367
R1174 B.n627 B.n625 163.367
R1175 B.n631 B.n605 163.367
R1176 B.n635 B.n633 163.367
R1177 B.n639 B.n603 163.367
R1178 B.n643 B.n641 163.367
R1179 B.n647 B.n601 163.367
R1180 B.n651 B.n649 163.367
R1181 B.n655 B.n599 163.367
R1182 B.n659 B.n657 163.367
R1183 B.n663 B.n597 163.367
R1184 B.n667 B.n665 163.367
R1185 B.n671 B.n595 163.367
R1186 B.n675 B.n673 163.367
R1187 B.n679 B.n593 163.367
R1188 B.n683 B.n681 163.367
R1189 B.n687 B.n591 163.367
R1190 B.n691 B.n689 163.367
R1191 B.n695 B.n589 163.367
R1192 B.n699 B.n697 163.367
R1193 B.n703 B.n587 163.367
R1194 B.n707 B.n705 163.367
R1195 B.n711 B.n585 163.367
R1196 B.n715 B.n713 163.367
R1197 B.n720 B.n581 163.367
R1198 B.n724 B.n722 163.367
R1199 B.n728 B.n579 163.367
R1200 B.n732 B.n730 163.367
R1201 B.n736 B.n577 163.367
R1202 B.n740 B.n738 163.367
R1203 B.n744 B.n572 163.367
R1204 B.n748 B.n746 163.367
R1205 B.n752 B.n570 163.367
R1206 B.n756 B.n754 163.367
R1207 B.n760 B.n568 163.367
R1208 B.n764 B.n762 163.367
R1209 B.n768 B.n566 163.367
R1210 B.n772 B.n770 163.367
R1211 B.n776 B.n564 163.367
R1212 B.n780 B.n778 163.367
R1213 B.n784 B.n562 163.367
R1214 B.n788 B.n786 163.367
R1215 B.n792 B.n560 163.367
R1216 B.n796 B.n794 163.367
R1217 B.n800 B.n558 163.367
R1218 B.n804 B.n802 163.367
R1219 B.n808 B.n556 163.367
R1220 B.n812 B.n810 163.367
R1221 B.n816 B.n554 163.367
R1222 B.n820 B.n818 163.367
R1223 B.n824 B.n552 163.367
R1224 B.n828 B.n826 163.367
R1225 B.n832 B.n550 163.367
R1226 B.n836 B.n834 163.367
R1227 B.n840 B.n548 163.367
R1228 B.n843 B.n842 163.367
R1229 B.n845 B.n545 163.367
R1230 B.n849 B.n539 163.367
R1231 B.n857 B.n539 163.367
R1232 B.n857 B.n537 163.367
R1233 B.n861 B.n537 163.367
R1234 B.n861 B.n531 163.367
R1235 B.n869 B.n531 163.367
R1236 B.n869 B.n529 163.367
R1237 B.n873 B.n529 163.367
R1238 B.n873 B.n523 163.367
R1239 B.n881 B.n523 163.367
R1240 B.n881 B.n521 163.367
R1241 B.n885 B.n521 163.367
R1242 B.n885 B.n515 163.367
R1243 B.n893 B.n515 163.367
R1244 B.n893 B.n513 163.367
R1245 B.n897 B.n513 163.367
R1246 B.n897 B.n507 163.367
R1247 B.n905 B.n507 163.367
R1248 B.n905 B.n505 163.367
R1249 B.n909 B.n505 163.367
R1250 B.n909 B.n498 163.367
R1251 B.n917 B.n498 163.367
R1252 B.n917 B.n496 163.367
R1253 B.n921 B.n496 163.367
R1254 B.n921 B.n491 163.367
R1255 B.n929 B.n491 163.367
R1256 B.n929 B.n489 163.367
R1257 B.n933 B.n489 163.367
R1258 B.n933 B.n483 163.367
R1259 B.n941 B.n483 163.367
R1260 B.n941 B.n481 163.367
R1261 B.n945 B.n481 163.367
R1262 B.n945 B.n475 163.367
R1263 B.n953 B.n475 163.367
R1264 B.n953 B.n473 163.367
R1265 B.n957 B.n473 163.367
R1266 B.n957 B.n467 163.367
R1267 B.n965 B.n467 163.367
R1268 B.n965 B.n465 163.367
R1269 B.n969 B.n465 163.367
R1270 B.n969 B.n459 163.367
R1271 B.n977 B.n459 163.367
R1272 B.n977 B.n457 163.367
R1273 B.n981 B.n457 163.367
R1274 B.n981 B.n452 163.367
R1275 B.n990 B.n452 163.367
R1276 B.n990 B.n450 163.367
R1277 B.n994 B.n450 163.367
R1278 B.n994 B.n444 163.367
R1279 B.n1002 B.n444 163.367
R1280 B.n1002 B.n442 163.367
R1281 B.n1006 B.n442 163.367
R1282 B.n1006 B.n436 163.367
R1283 B.n1014 B.n436 163.367
R1284 B.n1014 B.n434 163.367
R1285 B.n1018 B.n434 163.367
R1286 B.n1018 B.n428 163.367
R1287 B.n1026 B.n428 163.367
R1288 B.n1026 B.n426 163.367
R1289 B.n1031 B.n426 163.367
R1290 B.n1031 B.n420 163.367
R1291 B.n1039 B.n420 163.367
R1292 B.n1040 B.n1039 163.367
R1293 B.n1040 B.n5 163.367
R1294 B.n6 B.n5 163.367
R1295 B.n7 B.n6 163.367
R1296 B.n1045 B.n7 163.367
R1297 B.n1045 B.n12 163.367
R1298 B.n13 B.n12 163.367
R1299 B.n14 B.n13 163.367
R1300 B.n1050 B.n14 163.367
R1301 B.n1050 B.n19 163.367
R1302 B.n20 B.n19 163.367
R1303 B.n21 B.n20 163.367
R1304 B.n1055 B.n21 163.367
R1305 B.n1055 B.n26 163.367
R1306 B.n27 B.n26 163.367
R1307 B.n28 B.n27 163.367
R1308 B.n1060 B.n28 163.367
R1309 B.n1060 B.n33 163.367
R1310 B.n34 B.n33 163.367
R1311 B.n35 B.n34 163.367
R1312 B.n1065 B.n35 163.367
R1313 B.n1065 B.n40 163.367
R1314 B.n41 B.n40 163.367
R1315 B.n42 B.n41 163.367
R1316 B.n1070 B.n42 163.367
R1317 B.n1070 B.n47 163.367
R1318 B.n48 B.n47 163.367
R1319 B.n49 B.n48 163.367
R1320 B.n1075 B.n49 163.367
R1321 B.n1075 B.n54 163.367
R1322 B.n55 B.n54 163.367
R1323 B.n56 B.n55 163.367
R1324 B.n1080 B.n56 163.367
R1325 B.n1080 B.n61 163.367
R1326 B.n62 B.n61 163.367
R1327 B.n63 B.n62 163.367
R1328 B.n1085 B.n63 163.367
R1329 B.n1085 B.n68 163.367
R1330 B.n69 B.n68 163.367
R1331 B.n70 B.n69 163.367
R1332 B.n1090 B.n70 163.367
R1333 B.n1090 B.n75 163.367
R1334 B.n76 B.n75 163.367
R1335 B.n77 B.n76 163.367
R1336 B.n1095 B.n77 163.367
R1337 B.n1095 B.n82 163.367
R1338 B.n83 B.n82 163.367
R1339 B.n84 B.n83 163.367
R1340 B.n1100 B.n84 163.367
R1341 B.n1100 B.n89 163.367
R1342 B.n90 B.n89 163.367
R1343 B.n91 B.n90 163.367
R1344 B.n1105 B.n91 163.367
R1345 B.n1105 B.n96 163.367
R1346 B.n97 B.n96 163.367
R1347 B.n98 B.n97 163.367
R1348 B.n1110 B.n98 163.367
R1349 B.n1110 B.n103 163.367
R1350 B.n104 B.n103 163.367
R1351 B.n105 B.n104 163.367
R1352 B.n1115 B.n105 163.367
R1353 B.n1115 B.n110 163.367
R1354 B.n111 B.n110 163.367
R1355 B.n112 B.n111 163.367
R1356 B.n1120 B.n112 163.367
R1357 B.n1120 B.n117 163.367
R1358 B.n184 B.n183 163.367
R1359 B.n188 B.n187 163.367
R1360 B.n192 B.n191 163.367
R1361 B.n196 B.n195 163.367
R1362 B.n200 B.n199 163.367
R1363 B.n204 B.n203 163.367
R1364 B.n208 B.n207 163.367
R1365 B.n212 B.n211 163.367
R1366 B.n216 B.n215 163.367
R1367 B.n220 B.n219 163.367
R1368 B.n224 B.n223 163.367
R1369 B.n228 B.n227 163.367
R1370 B.n232 B.n231 163.367
R1371 B.n236 B.n235 163.367
R1372 B.n240 B.n239 163.367
R1373 B.n244 B.n243 163.367
R1374 B.n248 B.n247 163.367
R1375 B.n252 B.n251 163.367
R1376 B.n256 B.n255 163.367
R1377 B.n260 B.n259 163.367
R1378 B.n264 B.n263 163.367
R1379 B.n268 B.n267 163.367
R1380 B.n272 B.n271 163.367
R1381 B.n276 B.n275 163.367
R1382 B.n280 B.n279 163.367
R1383 B.n284 B.n283 163.367
R1384 B.n288 B.n287 163.367
R1385 B.n293 B.n292 163.367
R1386 B.n297 B.n296 163.367
R1387 B.n301 B.n300 163.367
R1388 B.n305 B.n304 163.367
R1389 B.n309 B.n308 163.367
R1390 B.n314 B.n313 163.367
R1391 B.n318 B.n317 163.367
R1392 B.n322 B.n321 163.367
R1393 B.n326 B.n325 163.367
R1394 B.n330 B.n329 163.367
R1395 B.n334 B.n333 163.367
R1396 B.n338 B.n337 163.367
R1397 B.n342 B.n341 163.367
R1398 B.n346 B.n345 163.367
R1399 B.n350 B.n349 163.367
R1400 B.n354 B.n353 163.367
R1401 B.n358 B.n357 163.367
R1402 B.n362 B.n361 163.367
R1403 B.n366 B.n365 163.367
R1404 B.n370 B.n369 163.367
R1405 B.n374 B.n373 163.367
R1406 B.n378 B.n377 163.367
R1407 B.n382 B.n381 163.367
R1408 B.n386 B.n385 163.367
R1409 B.n390 B.n389 163.367
R1410 B.n394 B.n393 163.367
R1411 B.n398 B.n397 163.367
R1412 B.n402 B.n401 163.367
R1413 B.n406 B.n405 163.367
R1414 B.n410 B.n409 163.367
R1415 B.n414 B.n413 163.367
R1416 B.n416 B.n177 163.367
R1417 B.n573 B.t10 145.501
R1418 B.n178 B.t13 145.501
R1419 B.n582 B.t17 145.48
R1420 B.n180 B.t19 145.48
R1421 B.n574 B.n573 73.8914
R1422 B.n583 B.n582 73.8914
R1423 B.n181 B.n180 73.8914
R1424 B.n179 B.n178 73.8914
R1425 B.n610 B.n543 71.676
R1426 B.n616 B.n615 71.676
R1427 B.n619 B.n618 71.676
R1428 B.n624 B.n623 71.676
R1429 B.n627 B.n626 71.676
R1430 B.n632 B.n631 71.676
R1431 B.n635 B.n634 71.676
R1432 B.n640 B.n639 71.676
R1433 B.n643 B.n642 71.676
R1434 B.n648 B.n647 71.676
R1435 B.n651 B.n650 71.676
R1436 B.n656 B.n655 71.676
R1437 B.n659 B.n658 71.676
R1438 B.n664 B.n663 71.676
R1439 B.n667 B.n666 71.676
R1440 B.n672 B.n671 71.676
R1441 B.n675 B.n674 71.676
R1442 B.n680 B.n679 71.676
R1443 B.n683 B.n682 71.676
R1444 B.n688 B.n687 71.676
R1445 B.n691 B.n690 71.676
R1446 B.n696 B.n695 71.676
R1447 B.n699 B.n698 71.676
R1448 B.n704 B.n703 71.676
R1449 B.n707 B.n706 71.676
R1450 B.n712 B.n711 71.676
R1451 B.n715 B.n714 71.676
R1452 B.n721 B.n720 71.676
R1453 B.n724 B.n723 71.676
R1454 B.n729 B.n728 71.676
R1455 B.n732 B.n731 71.676
R1456 B.n737 B.n736 71.676
R1457 B.n740 B.n739 71.676
R1458 B.n745 B.n744 71.676
R1459 B.n748 B.n747 71.676
R1460 B.n753 B.n752 71.676
R1461 B.n756 B.n755 71.676
R1462 B.n761 B.n760 71.676
R1463 B.n764 B.n763 71.676
R1464 B.n769 B.n768 71.676
R1465 B.n772 B.n771 71.676
R1466 B.n777 B.n776 71.676
R1467 B.n780 B.n779 71.676
R1468 B.n785 B.n784 71.676
R1469 B.n788 B.n787 71.676
R1470 B.n793 B.n792 71.676
R1471 B.n796 B.n795 71.676
R1472 B.n801 B.n800 71.676
R1473 B.n804 B.n803 71.676
R1474 B.n809 B.n808 71.676
R1475 B.n812 B.n811 71.676
R1476 B.n817 B.n816 71.676
R1477 B.n820 B.n819 71.676
R1478 B.n825 B.n824 71.676
R1479 B.n828 B.n827 71.676
R1480 B.n833 B.n832 71.676
R1481 B.n836 B.n835 71.676
R1482 B.n841 B.n840 71.676
R1483 B.n844 B.n843 71.676
R1484 B.n118 B.n116 71.676
R1485 B.n184 B.n119 71.676
R1486 B.n188 B.n120 71.676
R1487 B.n192 B.n121 71.676
R1488 B.n196 B.n122 71.676
R1489 B.n200 B.n123 71.676
R1490 B.n204 B.n124 71.676
R1491 B.n208 B.n125 71.676
R1492 B.n212 B.n126 71.676
R1493 B.n216 B.n127 71.676
R1494 B.n220 B.n128 71.676
R1495 B.n224 B.n129 71.676
R1496 B.n228 B.n130 71.676
R1497 B.n232 B.n131 71.676
R1498 B.n236 B.n132 71.676
R1499 B.n240 B.n133 71.676
R1500 B.n244 B.n134 71.676
R1501 B.n248 B.n135 71.676
R1502 B.n252 B.n136 71.676
R1503 B.n256 B.n137 71.676
R1504 B.n260 B.n138 71.676
R1505 B.n264 B.n139 71.676
R1506 B.n268 B.n140 71.676
R1507 B.n272 B.n141 71.676
R1508 B.n276 B.n142 71.676
R1509 B.n280 B.n143 71.676
R1510 B.n284 B.n144 71.676
R1511 B.n288 B.n145 71.676
R1512 B.n293 B.n146 71.676
R1513 B.n297 B.n147 71.676
R1514 B.n301 B.n148 71.676
R1515 B.n305 B.n149 71.676
R1516 B.n309 B.n150 71.676
R1517 B.n314 B.n151 71.676
R1518 B.n318 B.n152 71.676
R1519 B.n322 B.n153 71.676
R1520 B.n326 B.n154 71.676
R1521 B.n330 B.n155 71.676
R1522 B.n334 B.n156 71.676
R1523 B.n338 B.n157 71.676
R1524 B.n342 B.n158 71.676
R1525 B.n346 B.n159 71.676
R1526 B.n350 B.n160 71.676
R1527 B.n354 B.n161 71.676
R1528 B.n358 B.n162 71.676
R1529 B.n362 B.n163 71.676
R1530 B.n366 B.n164 71.676
R1531 B.n370 B.n165 71.676
R1532 B.n374 B.n166 71.676
R1533 B.n378 B.n167 71.676
R1534 B.n382 B.n168 71.676
R1535 B.n386 B.n169 71.676
R1536 B.n390 B.n170 71.676
R1537 B.n394 B.n171 71.676
R1538 B.n398 B.n172 71.676
R1539 B.n402 B.n173 71.676
R1540 B.n406 B.n174 71.676
R1541 B.n410 B.n175 71.676
R1542 B.n414 B.n176 71.676
R1543 B.n1125 B.n177 71.676
R1544 B.n1125 B.n1124 71.676
R1545 B.n416 B.n176 71.676
R1546 B.n413 B.n175 71.676
R1547 B.n409 B.n174 71.676
R1548 B.n405 B.n173 71.676
R1549 B.n401 B.n172 71.676
R1550 B.n397 B.n171 71.676
R1551 B.n393 B.n170 71.676
R1552 B.n389 B.n169 71.676
R1553 B.n385 B.n168 71.676
R1554 B.n381 B.n167 71.676
R1555 B.n377 B.n166 71.676
R1556 B.n373 B.n165 71.676
R1557 B.n369 B.n164 71.676
R1558 B.n365 B.n163 71.676
R1559 B.n361 B.n162 71.676
R1560 B.n357 B.n161 71.676
R1561 B.n353 B.n160 71.676
R1562 B.n349 B.n159 71.676
R1563 B.n345 B.n158 71.676
R1564 B.n341 B.n157 71.676
R1565 B.n337 B.n156 71.676
R1566 B.n333 B.n155 71.676
R1567 B.n329 B.n154 71.676
R1568 B.n325 B.n153 71.676
R1569 B.n321 B.n152 71.676
R1570 B.n317 B.n151 71.676
R1571 B.n313 B.n150 71.676
R1572 B.n308 B.n149 71.676
R1573 B.n304 B.n148 71.676
R1574 B.n300 B.n147 71.676
R1575 B.n296 B.n146 71.676
R1576 B.n292 B.n145 71.676
R1577 B.n287 B.n144 71.676
R1578 B.n283 B.n143 71.676
R1579 B.n279 B.n142 71.676
R1580 B.n275 B.n141 71.676
R1581 B.n271 B.n140 71.676
R1582 B.n267 B.n139 71.676
R1583 B.n263 B.n138 71.676
R1584 B.n259 B.n137 71.676
R1585 B.n255 B.n136 71.676
R1586 B.n251 B.n135 71.676
R1587 B.n247 B.n134 71.676
R1588 B.n243 B.n133 71.676
R1589 B.n239 B.n132 71.676
R1590 B.n235 B.n131 71.676
R1591 B.n231 B.n130 71.676
R1592 B.n227 B.n129 71.676
R1593 B.n223 B.n128 71.676
R1594 B.n219 B.n127 71.676
R1595 B.n215 B.n126 71.676
R1596 B.n211 B.n125 71.676
R1597 B.n207 B.n124 71.676
R1598 B.n203 B.n123 71.676
R1599 B.n199 B.n122 71.676
R1600 B.n195 B.n121 71.676
R1601 B.n191 B.n120 71.676
R1602 B.n187 B.n119 71.676
R1603 B.n183 B.n118 71.676
R1604 B.n611 B.n610 71.676
R1605 B.n617 B.n616 71.676
R1606 B.n618 B.n607 71.676
R1607 B.n625 B.n624 71.676
R1608 B.n626 B.n605 71.676
R1609 B.n633 B.n632 71.676
R1610 B.n634 B.n603 71.676
R1611 B.n641 B.n640 71.676
R1612 B.n642 B.n601 71.676
R1613 B.n649 B.n648 71.676
R1614 B.n650 B.n599 71.676
R1615 B.n657 B.n656 71.676
R1616 B.n658 B.n597 71.676
R1617 B.n665 B.n664 71.676
R1618 B.n666 B.n595 71.676
R1619 B.n673 B.n672 71.676
R1620 B.n674 B.n593 71.676
R1621 B.n681 B.n680 71.676
R1622 B.n682 B.n591 71.676
R1623 B.n689 B.n688 71.676
R1624 B.n690 B.n589 71.676
R1625 B.n697 B.n696 71.676
R1626 B.n698 B.n587 71.676
R1627 B.n705 B.n704 71.676
R1628 B.n706 B.n585 71.676
R1629 B.n713 B.n712 71.676
R1630 B.n714 B.n581 71.676
R1631 B.n722 B.n721 71.676
R1632 B.n723 B.n579 71.676
R1633 B.n730 B.n729 71.676
R1634 B.n731 B.n577 71.676
R1635 B.n738 B.n737 71.676
R1636 B.n739 B.n572 71.676
R1637 B.n746 B.n745 71.676
R1638 B.n747 B.n570 71.676
R1639 B.n754 B.n753 71.676
R1640 B.n755 B.n568 71.676
R1641 B.n762 B.n761 71.676
R1642 B.n763 B.n566 71.676
R1643 B.n770 B.n769 71.676
R1644 B.n771 B.n564 71.676
R1645 B.n778 B.n777 71.676
R1646 B.n779 B.n562 71.676
R1647 B.n786 B.n785 71.676
R1648 B.n787 B.n560 71.676
R1649 B.n794 B.n793 71.676
R1650 B.n795 B.n558 71.676
R1651 B.n802 B.n801 71.676
R1652 B.n803 B.n556 71.676
R1653 B.n810 B.n809 71.676
R1654 B.n811 B.n554 71.676
R1655 B.n818 B.n817 71.676
R1656 B.n819 B.n552 71.676
R1657 B.n826 B.n825 71.676
R1658 B.n827 B.n550 71.676
R1659 B.n834 B.n833 71.676
R1660 B.n835 B.n548 71.676
R1661 B.n842 B.n841 71.676
R1662 B.n845 B.n844 71.676
R1663 B.n574 B.t9 71.6102
R1664 B.n179 B.t14 71.6102
R1665 B.n583 B.t16 71.5884
R1666 B.n181 B.t20 71.5884
R1667 B.n850 B.n544 67.0644
R1668 B.n1127 B.n1126 67.0644
R1669 B.n575 B.n574 59.5399
R1670 B.n718 B.n583 59.5399
R1671 B.n290 B.n181 59.5399
R1672 B.n311 B.n179 59.5399
R1673 B.n850 B.n540 34.2888
R1674 B.n856 B.n540 34.2888
R1675 B.n856 B.n536 34.2888
R1676 B.n862 B.n536 34.2888
R1677 B.n862 B.n532 34.2888
R1678 B.n868 B.n532 34.2888
R1679 B.n868 B.n528 34.2888
R1680 B.n874 B.n528 34.2888
R1681 B.n880 B.n524 34.2888
R1682 B.n880 B.n520 34.2888
R1683 B.n886 B.n520 34.2888
R1684 B.n886 B.n516 34.2888
R1685 B.n892 B.n516 34.2888
R1686 B.n892 B.n512 34.2888
R1687 B.n898 B.n512 34.2888
R1688 B.n898 B.n508 34.2888
R1689 B.n904 B.n508 34.2888
R1690 B.n904 B.n504 34.2888
R1691 B.n910 B.n504 34.2888
R1692 B.n910 B.n499 34.2888
R1693 B.n916 B.n499 34.2888
R1694 B.n916 B.n500 34.2888
R1695 B.n922 B.n492 34.2888
R1696 B.n928 B.n492 34.2888
R1697 B.n928 B.n488 34.2888
R1698 B.n934 B.n488 34.2888
R1699 B.n934 B.n484 34.2888
R1700 B.n940 B.n484 34.2888
R1701 B.n940 B.n480 34.2888
R1702 B.n946 B.n480 34.2888
R1703 B.n946 B.n476 34.2888
R1704 B.n952 B.n476 34.2888
R1705 B.n958 B.n472 34.2888
R1706 B.n958 B.n468 34.2888
R1707 B.n964 B.n468 34.2888
R1708 B.n964 B.n464 34.2888
R1709 B.n970 B.n464 34.2888
R1710 B.n970 B.n460 34.2888
R1711 B.n976 B.n460 34.2888
R1712 B.n976 B.n456 34.2888
R1713 B.n983 B.n456 34.2888
R1714 B.n983 B.n982 34.2888
R1715 B.n989 B.n449 34.2888
R1716 B.n995 B.n449 34.2888
R1717 B.n995 B.n445 34.2888
R1718 B.n1001 B.n445 34.2888
R1719 B.n1001 B.n441 34.2888
R1720 B.n1007 B.n441 34.2888
R1721 B.n1007 B.n437 34.2888
R1722 B.n1013 B.n437 34.2888
R1723 B.n1013 B.n433 34.2888
R1724 B.n1019 B.n433 34.2888
R1725 B.n1025 B.n429 34.2888
R1726 B.n1025 B.n425 34.2888
R1727 B.n1032 B.n425 34.2888
R1728 B.n1032 B.n421 34.2888
R1729 B.n1038 B.n421 34.2888
R1730 B.n1038 B.n4 34.2888
R1731 B.n1255 B.n4 34.2888
R1732 B.n1255 B.n1254 34.2888
R1733 B.n1254 B.n1253 34.2888
R1734 B.n1253 B.n8 34.2888
R1735 B.n1247 B.n8 34.2888
R1736 B.n1247 B.n1246 34.2888
R1737 B.n1246 B.n1245 34.2888
R1738 B.n1245 B.n15 34.2888
R1739 B.n1239 B.n1238 34.2888
R1740 B.n1238 B.n1237 34.2888
R1741 B.n1237 B.n22 34.2888
R1742 B.n1231 B.n22 34.2888
R1743 B.n1231 B.n1230 34.2888
R1744 B.n1230 B.n1229 34.2888
R1745 B.n1229 B.n29 34.2888
R1746 B.n1223 B.n29 34.2888
R1747 B.n1223 B.n1222 34.2888
R1748 B.n1222 B.n1221 34.2888
R1749 B.n1215 B.n39 34.2888
R1750 B.n1215 B.n1214 34.2888
R1751 B.n1214 B.n1213 34.2888
R1752 B.n1213 B.n43 34.2888
R1753 B.n1207 B.n43 34.2888
R1754 B.n1207 B.n1206 34.2888
R1755 B.n1206 B.n1205 34.2888
R1756 B.n1205 B.n50 34.2888
R1757 B.n1199 B.n50 34.2888
R1758 B.n1199 B.n1198 34.2888
R1759 B.n1197 B.n57 34.2888
R1760 B.n1191 B.n57 34.2888
R1761 B.n1191 B.n1190 34.2888
R1762 B.n1190 B.n1189 34.2888
R1763 B.n1189 B.n64 34.2888
R1764 B.n1183 B.n64 34.2888
R1765 B.n1183 B.n1182 34.2888
R1766 B.n1182 B.n1181 34.2888
R1767 B.n1181 B.n71 34.2888
R1768 B.n1175 B.n71 34.2888
R1769 B.n1174 B.n1173 34.2888
R1770 B.n1173 B.n78 34.2888
R1771 B.n1167 B.n78 34.2888
R1772 B.n1167 B.n1166 34.2888
R1773 B.n1166 B.n1165 34.2888
R1774 B.n1165 B.n85 34.2888
R1775 B.n1159 B.n85 34.2888
R1776 B.n1159 B.n1158 34.2888
R1777 B.n1158 B.n1157 34.2888
R1778 B.n1157 B.n92 34.2888
R1779 B.n1151 B.n92 34.2888
R1780 B.n1151 B.n1150 34.2888
R1781 B.n1150 B.n1149 34.2888
R1782 B.n1149 B.n99 34.2888
R1783 B.n1143 B.n1142 34.2888
R1784 B.n1142 B.n1141 34.2888
R1785 B.n1141 B.n106 34.2888
R1786 B.n1135 B.n106 34.2888
R1787 B.n1135 B.n1134 34.2888
R1788 B.n1134 B.n1133 34.2888
R1789 B.n1133 B.n113 34.2888
R1790 B.n1127 B.n113 34.2888
R1791 B.n1129 B.n115 31.3761
R1792 B.n1123 B.n1122 31.3761
R1793 B.n848 B.n847 31.3761
R1794 B.n852 B.n542 31.3761
R1795 B.n922 B.t3 28.238
R1796 B.n1175 B.t5 28.238
R1797 B.n1019 B.t1 27.2295
R1798 B.n1239 B.t0 27.2295
R1799 B.n874 B.t8 26.221
R1800 B.n1143 B.t12 26.221
R1801 B.t2 B.n472 21.1786
R1802 B.n1198 B.t21 21.1786
R1803 B.n982 B.t4 20.1701
R1804 B.n39 B.t6 20.1701
R1805 B B.n1257 18.0485
R1806 B.n989 B.t4 14.1192
R1807 B.n1221 B.t6 14.1192
R1808 B.n952 B.t2 13.1107
R1809 B.t21 B.n1197 13.1107
R1810 B.n182 B.n115 10.6151
R1811 B.n185 B.n182 10.6151
R1812 B.n186 B.n185 10.6151
R1813 B.n189 B.n186 10.6151
R1814 B.n190 B.n189 10.6151
R1815 B.n193 B.n190 10.6151
R1816 B.n194 B.n193 10.6151
R1817 B.n197 B.n194 10.6151
R1818 B.n198 B.n197 10.6151
R1819 B.n201 B.n198 10.6151
R1820 B.n202 B.n201 10.6151
R1821 B.n205 B.n202 10.6151
R1822 B.n206 B.n205 10.6151
R1823 B.n209 B.n206 10.6151
R1824 B.n210 B.n209 10.6151
R1825 B.n213 B.n210 10.6151
R1826 B.n214 B.n213 10.6151
R1827 B.n217 B.n214 10.6151
R1828 B.n218 B.n217 10.6151
R1829 B.n221 B.n218 10.6151
R1830 B.n222 B.n221 10.6151
R1831 B.n225 B.n222 10.6151
R1832 B.n226 B.n225 10.6151
R1833 B.n229 B.n226 10.6151
R1834 B.n230 B.n229 10.6151
R1835 B.n233 B.n230 10.6151
R1836 B.n234 B.n233 10.6151
R1837 B.n237 B.n234 10.6151
R1838 B.n238 B.n237 10.6151
R1839 B.n241 B.n238 10.6151
R1840 B.n242 B.n241 10.6151
R1841 B.n245 B.n242 10.6151
R1842 B.n246 B.n245 10.6151
R1843 B.n249 B.n246 10.6151
R1844 B.n250 B.n249 10.6151
R1845 B.n253 B.n250 10.6151
R1846 B.n254 B.n253 10.6151
R1847 B.n257 B.n254 10.6151
R1848 B.n258 B.n257 10.6151
R1849 B.n261 B.n258 10.6151
R1850 B.n262 B.n261 10.6151
R1851 B.n265 B.n262 10.6151
R1852 B.n266 B.n265 10.6151
R1853 B.n269 B.n266 10.6151
R1854 B.n270 B.n269 10.6151
R1855 B.n273 B.n270 10.6151
R1856 B.n274 B.n273 10.6151
R1857 B.n277 B.n274 10.6151
R1858 B.n278 B.n277 10.6151
R1859 B.n281 B.n278 10.6151
R1860 B.n282 B.n281 10.6151
R1861 B.n285 B.n282 10.6151
R1862 B.n286 B.n285 10.6151
R1863 B.n289 B.n286 10.6151
R1864 B.n294 B.n291 10.6151
R1865 B.n295 B.n294 10.6151
R1866 B.n298 B.n295 10.6151
R1867 B.n299 B.n298 10.6151
R1868 B.n302 B.n299 10.6151
R1869 B.n303 B.n302 10.6151
R1870 B.n306 B.n303 10.6151
R1871 B.n307 B.n306 10.6151
R1872 B.n310 B.n307 10.6151
R1873 B.n315 B.n312 10.6151
R1874 B.n316 B.n315 10.6151
R1875 B.n319 B.n316 10.6151
R1876 B.n320 B.n319 10.6151
R1877 B.n323 B.n320 10.6151
R1878 B.n324 B.n323 10.6151
R1879 B.n327 B.n324 10.6151
R1880 B.n328 B.n327 10.6151
R1881 B.n331 B.n328 10.6151
R1882 B.n332 B.n331 10.6151
R1883 B.n335 B.n332 10.6151
R1884 B.n336 B.n335 10.6151
R1885 B.n339 B.n336 10.6151
R1886 B.n340 B.n339 10.6151
R1887 B.n343 B.n340 10.6151
R1888 B.n344 B.n343 10.6151
R1889 B.n347 B.n344 10.6151
R1890 B.n348 B.n347 10.6151
R1891 B.n351 B.n348 10.6151
R1892 B.n352 B.n351 10.6151
R1893 B.n355 B.n352 10.6151
R1894 B.n356 B.n355 10.6151
R1895 B.n359 B.n356 10.6151
R1896 B.n360 B.n359 10.6151
R1897 B.n363 B.n360 10.6151
R1898 B.n364 B.n363 10.6151
R1899 B.n367 B.n364 10.6151
R1900 B.n368 B.n367 10.6151
R1901 B.n371 B.n368 10.6151
R1902 B.n372 B.n371 10.6151
R1903 B.n375 B.n372 10.6151
R1904 B.n376 B.n375 10.6151
R1905 B.n379 B.n376 10.6151
R1906 B.n380 B.n379 10.6151
R1907 B.n383 B.n380 10.6151
R1908 B.n384 B.n383 10.6151
R1909 B.n387 B.n384 10.6151
R1910 B.n388 B.n387 10.6151
R1911 B.n391 B.n388 10.6151
R1912 B.n392 B.n391 10.6151
R1913 B.n395 B.n392 10.6151
R1914 B.n396 B.n395 10.6151
R1915 B.n399 B.n396 10.6151
R1916 B.n400 B.n399 10.6151
R1917 B.n403 B.n400 10.6151
R1918 B.n404 B.n403 10.6151
R1919 B.n407 B.n404 10.6151
R1920 B.n408 B.n407 10.6151
R1921 B.n411 B.n408 10.6151
R1922 B.n412 B.n411 10.6151
R1923 B.n415 B.n412 10.6151
R1924 B.n417 B.n415 10.6151
R1925 B.n418 B.n417 10.6151
R1926 B.n1123 B.n418 10.6151
R1927 B.n848 B.n538 10.6151
R1928 B.n858 B.n538 10.6151
R1929 B.n859 B.n858 10.6151
R1930 B.n860 B.n859 10.6151
R1931 B.n860 B.n530 10.6151
R1932 B.n870 B.n530 10.6151
R1933 B.n871 B.n870 10.6151
R1934 B.n872 B.n871 10.6151
R1935 B.n872 B.n522 10.6151
R1936 B.n882 B.n522 10.6151
R1937 B.n883 B.n882 10.6151
R1938 B.n884 B.n883 10.6151
R1939 B.n884 B.n514 10.6151
R1940 B.n894 B.n514 10.6151
R1941 B.n895 B.n894 10.6151
R1942 B.n896 B.n895 10.6151
R1943 B.n896 B.n506 10.6151
R1944 B.n906 B.n506 10.6151
R1945 B.n907 B.n906 10.6151
R1946 B.n908 B.n907 10.6151
R1947 B.n908 B.n497 10.6151
R1948 B.n918 B.n497 10.6151
R1949 B.n919 B.n918 10.6151
R1950 B.n920 B.n919 10.6151
R1951 B.n920 B.n490 10.6151
R1952 B.n930 B.n490 10.6151
R1953 B.n931 B.n930 10.6151
R1954 B.n932 B.n931 10.6151
R1955 B.n932 B.n482 10.6151
R1956 B.n942 B.n482 10.6151
R1957 B.n943 B.n942 10.6151
R1958 B.n944 B.n943 10.6151
R1959 B.n944 B.n474 10.6151
R1960 B.n954 B.n474 10.6151
R1961 B.n955 B.n954 10.6151
R1962 B.n956 B.n955 10.6151
R1963 B.n956 B.n466 10.6151
R1964 B.n966 B.n466 10.6151
R1965 B.n967 B.n966 10.6151
R1966 B.n968 B.n967 10.6151
R1967 B.n968 B.n458 10.6151
R1968 B.n978 B.n458 10.6151
R1969 B.n979 B.n978 10.6151
R1970 B.n980 B.n979 10.6151
R1971 B.n980 B.n451 10.6151
R1972 B.n991 B.n451 10.6151
R1973 B.n992 B.n991 10.6151
R1974 B.n993 B.n992 10.6151
R1975 B.n993 B.n443 10.6151
R1976 B.n1003 B.n443 10.6151
R1977 B.n1004 B.n1003 10.6151
R1978 B.n1005 B.n1004 10.6151
R1979 B.n1005 B.n435 10.6151
R1980 B.n1015 B.n435 10.6151
R1981 B.n1016 B.n1015 10.6151
R1982 B.n1017 B.n1016 10.6151
R1983 B.n1017 B.n427 10.6151
R1984 B.n1027 B.n427 10.6151
R1985 B.n1028 B.n1027 10.6151
R1986 B.n1030 B.n1028 10.6151
R1987 B.n1030 B.n1029 10.6151
R1988 B.n1029 B.n419 10.6151
R1989 B.n1041 B.n419 10.6151
R1990 B.n1042 B.n1041 10.6151
R1991 B.n1043 B.n1042 10.6151
R1992 B.n1044 B.n1043 10.6151
R1993 B.n1046 B.n1044 10.6151
R1994 B.n1047 B.n1046 10.6151
R1995 B.n1048 B.n1047 10.6151
R1996 B.n1049 B.n1048 10.6151
R1997 B.n1051 B.n1049 10.6151
R1998 B.n1052 B.n1051 10.6151
R1999 B.n1053 B.n1052 10.6151
R2000 B.n1054 B.n1053 10.6151
R2001 B.n1056 B.n1054 10.6151
R2002 B.n1057 B.n1056 10.6151
R2003 B.n1058 B.n1057 10.6151
R2004 B.n1059 B.n1058 10.6151
R2005 B.n1061 B.n1059 10.6151
R2006 B.n1062 B.n1061 10.6151
R2007 B.n1063 B.n1062 10.6151
R2008 B.n1064 B.n1063 10.6151
R2009 B.n1066 B.n1064 10.6151
R2010 B.n1067 B.n1066 10.6151
R2011 B.n1068 B.n1067 10.6151
R2012 B.n1069 B.n1068 10.6151
R2013 B.n1071 B.n1069 10.6151
R2014 B.n1072 B.n1071 10.6151
R2015 B.n1073 B.n1072 10.6151
R2016 B.n1074 B.n1073 10.6151
R2017 B.n1076 B.n1074 10.6151
R2018 B.n1077 B.n1076 10.6151
R2019 B.n1078 B.n1077 10.6151
R2020 B.n1079 B.n1078 10.6151
R2021 B.n1081 B.n1079 10.6151
R2022 B.n1082 B.n1081 10.6151
R2023 B.n1083 B.n1082 10.6151
R2024 B.n1084 B.n1083 10.6151
R2025 B.n1086 B.n1084 10.6151
R2026 B.n1087 B.n1086 10.6151
R2027 B.n1088 B.n1087 10.6151
R2028 B.n1089 B.n1088 10.6151
R2029 B.n1091 B.n1089 10.6151
R2030 B.n1092 B.n1091 10.6151
R2031 B.n1093 B.n1092 10.6151
R2032 B.n1094 B.n1093 10.6151
R2033 B.n1096 B.n1094 10.6151
R2034 B.n1097 B.n1096 10.6151
R2035 B.n1098 B.n1097 10.6151
R2036 B.n1099 B.n1098 10.6151
R2037 B.n1101 B.n1099 10.6151
R2038 B.n1102 B.n1101 10.6151
R2039 B.n1103 B.n1102 10.6151
R2040 B.n1104 B.n1103 10.6151
R2041 B.n1106 B.n1104 10.6151
R2042 B.n1107 B.n1106 10.6151
R2043 B.n1108 B.n1107 10.6151
R2044 B.n1109 B.n1108 10.6151
R2045 B.n1111 B.n1109 10.6151
R2046 B.n1112 B.n1111 10.6151
R2047 B.n1113 B.n1112 10.6151
R2048 B.n1114 B.n1113 10.6151
R2049 B.n1116 B.n1114 10.6151
R2050 B.n1117 B.n1116 10.6151
R2051 B.n1118 B.n1117 10.6151
R2052 B.n1119 B.n1118 10.6151
R2053 B.n1121 B.n1119 10.6151
R2054 B.n1122 B.n1121 10.6151
R2055 B.n612 B.n542 10.6151
R2056 B.n613 B.n612 10.6151
R2057 B.n614 B.n613 10.6151
R2058 B.n614 B.n608 10.6151
R2059 B.n620 B.n608 10.6151
R2060 B.n621 B.n620 10.6151
R2061 B.n622 B.n621 10.6151
R2062 B.n622 B.n606 10.6151
R2063 B.n628 B.n606 10.6151
R2064 B.n629 B.n628 10.6151
R2065 B.n630 B.n629 10.6151
R2066 B.n630 B.n604 10.6151
R2067 B.n636 B.n604 10.6151
R2068 B.n637 B.n636 10.6151
R2069 B.n638 B.n637 10.6151
R2070 B.n638 B.n602 10.6151
R2071 B.n644 B.n602 10.6151
R2072 B.n645 B.n644 10.6151
R2073 B.n646 B.n645 10.6151
R2074 B.n646 B.n600 10.6151
R2075 B.n652 B.n600 10.6151
R2076 B.n653 B.n652 10.6151
R2077 B.n654 B.n653 10.6151
R2078 B.n654 B.n598 10.6151
R2079 B.n660 B.n598 10.6151
R2080 B.n661 B.n660 10.6151
R2081 B.n662 B.n661 10.6151
R2082 B.n662 B.n596 10.6151
R2083 B.n668 B.n596 10.6151
R2084 B.n669 B.n668 10.6151
R2085 B.n670 B.n669 10.6151
R2086 B.n670 B.n594 10.6151
R2087 B.n676 B.n594 10.6151
R2088 B.n677 B.n676 10.6151
R2089 B.n678 B.n677 10.6151
R2090 B.n678 B.n592 10.6151
R2091 B.n684 B.n592 10.6151
R2092 B.n685 B.n684 10.6151
R2093 B.n686 B.n685 10.6151
R2094 B.n686 B.n590 10.6151
R2095 B.n692 B.n590 10.6151
R2096 B.n693 B.n692 10.6151
R2097 B.n694 B.n693 10.6151
R2098 B.n694 B.n588 10.6151
R2099 B.n700 B.n588 10.6151
R2100 B.n701 B.n700 10.6151
R2101 B.n702 B.n701 10.6151
R2102 B.n702 B.n586 10.6151
R2103 B.n708 B.n586 10.6151
R2104 B.n709 B.n708 10.6151
R2105 B.n710 B.n709 10.6151
R2106 B.n710 B.n584 10.6151
R2107 B.n716 B.n584 10.6151
R2108 B.n717 B.n716 10.6151
R2109 B.n719 B.n580 10.6151
R2110 B.n725 B.n580 10.6151
R2111 B.n726 B.n725 10.6151
R2112 B.n727 B.n726 10.6151
R2113 B.n727 B.n578 10.6151
R2114 B.n733 B.n578 10.6151
R2115 B.n734 B.n733 10.6151
R2116 B.n735 B.n734 10.6151
R2117 B.n735 B.n576 10.6151
R2118 B.n742 B.n741 10.6151
R2119 B.n743 B.n742 10.6151
R2120 B.n743 B.n571 10.6151
R2121 B.n749 B.n571 10.6151
R2122 B.n750 B.n749 10.6151
R2123 B.n751 B.n750 10.6151
R2124 B.n751 B.n569 10.6151
R2125 B.n757 B.n569 10.6151
R2126 B.n758 B.n757 10.6151
R2127 B.n759 B.n758 10.6151
R2128 B.n759 B.n567 10.6151
R2129 B.n765 B.n567 10.6151
R2130 B.n766 B.n765 10.6151
R2131 B.n767 B.n766 10.6151
R2132 B.n767 B.n565 10.6151
R2133 B.n773 B.n565 10.6151
R2134 B.n774 B.n773 10.6151
R2135 B.n775 B.n774 10.6151
R2136 B.n775 B.n563 10.6151
R2137 B.n781 B.n563 10.6151
R2138 B.n782 B.n781 10.6151
R2139 B.n783 B.n782 10.6151
R2140 B.n783 B.n561 10.6151
R2141 B.n789 B.n561 10.6151
R2142 B.n790 B.n789 10.6151
R2143 B.n791 B.n790 10.6151
R2144 B.n791 B.n559 10.6151
R2145 B.n797 B.n559 10.6151
R2146 B.n798 B.n797 10.6151
R2147 B.n799 B.n798 10.6151
R2148 B.n799 B.n557 10.6151
R2149 B.n805 B.n557 10.6151
R2150 B.n806 B.n805 10.6151
R2151 B.n807 B.n806 10.6151
R2152 B.n807 B.n555 10.6151
R2153 B.n813 B.n555 10.6151
R2154 B.n814 B.n813 10.6151
R2155 B.n815 B.n814 10.6151
R2156 B.n815 B.n553 10.6151
R2157 B.n821 B.n553 10.6151
R2158 B.n822 B.n821 10.6151
R2159 B.n823 B.n822 10.6151
R2160 B.n823 B.n551 10.6151
R2161 B.n829 B.n551 10.6151
R2162 B.n830 B.n829 10.6151
R2163 B.n831 B.n830 10.6151
R2164 B.n831 B.n549 10.6151
R2165 B.n837 B.n549 10.6151
R2166 B.n838 B.n837 10.6151
R2167 B.n839 B.n838 10.6151
R2168 B.n839 B.n547 10.6151
R2169 B.n547 B.n546 10.6151
R2170 B.n846 B.n546 10.6151
R2171 B.n847 B.n846 10.6151
R2172 B.n853 B.n852 10.6151
R2173 B.n854 B.n853 10.6151
R2174 B.n854 B.n534 10.6151
R2175 B.n864 B.n534 10.6151
R2176 B.n865 B.n864 10.6151
R2177 B.n866 B.n865 10.6151
R2178 B.n866 B.n526 10.6151
R2179 B.n876 B.n526 10.6151
R2180 B.n877 B.n876 10.6151
R2181 B.n878 B.n877 10.6151
R2182 B.n878 B.n518 10.6151
R2183 B.n888 B.n518 10.6151
R2184 B.n889 B.n888 10.6151
R2185 B.n890 B.n889 10.6151
R2186 B.n890 B.n510 10.6151
R2187 B.n900 B.n510 10.6151
R2188 B.n901 B.n900 10.6151
R2189 B.n902 B.n901 10.6151
R2190 B.n902 B.n502 10.6151
R2191 B.n912 B.n502 10.6151
R2192 B.n913 B.n912 10.6151
R2193 B.n914 B.n913 10.6151
R2194 B.n914 B.n494 10.6151
R2195 B.n924 B.n494 10.6151
R2196 B.n925 B.n924 10.6151
R2197 B.n926 B.n925 10.6151
R2198 B.n926 B.n486 10.6151
R2199 B.n936 B.n486 10.6151
R2200 B.n937 B.n936 10.6151
R2201 B.n938 B.n937 10.6151
R2202 B.n938 B.n478 10.6151
R2203 B.n948 B.n478 10.6151
R2204 B.n949 B.n948 10.6151
R2205 B.n950 B.n949 10.6151
R2206 B.n950 B.n470 10.6151
R2207 B.n960 B.n470 10.6151
R2208 B.n961 B.n960 10.6151
R2209 B.n962 B.n961 10.6151
R2210 B.n962 B.n462 10.6151
R2211 B.n972 B.n462 10.6151
R2212 B.n973 B.n972 10.6151
R2213 B.n974 B.n973 10.6151
R2214 B.n974 B.n454 10.6151
R2215 B.n985 B.n454 10.6151
R2216 B.n986 B.n985 10.6151
R2217 B.n987 B.n986 10.6151
R2218 B.n987 B.n447 10.6151
R2219 B.n997 B.n447 10.6151
R2220 B.n998 B.n997 10.6151
R2221 B.n999 B.n998 10.6151
R2222 B.n999 B.n439 10.6151
R2223 B.n1009 B.n439 10.6151
R2224 B.n1010 B.n1009 10.6151
R2225 B.n1011 B.n1010 10.6151
R2226 B.n1011 B.n431 10.6151
R2227 B.n1021 B.n431 10.6151
R2228 B.n1022 B.n1021 10.6151
R2229 B.n1023 B.n1022 10.6151
R2230 B.n1023 B.n423 10.6151
R2231 B.n1034 B.n423 10.6151
R2232 B.n1035 B.n1034 10.6151
R2233 B.n1036 B.n1035 10.6151
R2234 B.n1036 B.n0 10.6151
R2235 B.n1251 B.n1 10.6151
R2236 B.n1251 B.n1250 10.6151
R2237 B.n1250 B.n1249 10.6151
R2238 B.n1249 B.n10 10.6151
R2239 B.n1243 B.n10 10.6151
R2240 B.n1243 B.n1242 10.6151
R2241 B.n1242 B.n1241 10.6151
R2242 B.n1241 B.n17 10.6151
R2243 B.n1235 B.n17 10.6151
R2244 B.n1235 B.n1234 10.6151
R2245 B.n1234 B.n1233 10.6151
R2246 B.n1233 B.n24 10.6151
R2247 B.n1227 B.n24 10.6151
R2248 B.n1227 B.n1226 10.6151
R2249 B.n1226 B.n1225 10.6151
R2250 B.n1225 B.n31 10.6151
R2251 B.n1219 B.n31 10.6151
R2252 B.n1219 B.n1218 10.6151
R2253 B.n1218 B.n1217 10.6151
R2254 B.n1217 B.n37 10.6151
R2255 B.n1211 B.n37 10.6151
R2256 B.n1211 B.n1210 10.6151
R2257 B.n1210 B.n1209 10.6151
R2258 B.n1209 B.n45 10.6151
R2259 B.n1203 B.n45 10.6151
R2260 B.n1203 B.n1202 10.6151
R2261 B.n1202 B.n1201 10.6151
R2262 B.n1201 B.n52 10.6151
R2263 B.n1195 B.n52 10.6151
R2264 B.n1195 B.n1194 10.6151
R2265 B.n1194 B.n1193 10.6151
R2266 B.n1193 B.n59 10.6151
R2267 B.n1187 B.n59 10.6151
R2268 B.n1187 B.n1186 10.6151
R2269 B.n1186 B.n1185 10.6151
R2270 B.n1185 B.n66 10.6151
R2271 B.n1179 B.n66 10.6151
R2272 B.n1179 B.n1178 10.6151
R2273 B.n1178 B.n1177 10.6151
R2274 B.n1177 B.n73 10.6151
R2275 B.n1171 B.n73 10.6151
R2276 B.n1171 B.n1170 10.6151
R2277 B.n1170 B.n1169 10.6151
R2278 B.n1169 B.n80 10.6151
R2279 B.n1163 B.n80 10.6151
R2280 B.n1163 B.n1162 10.6151
R2281 B.n1162 B.n1161 10.6151
R2282 B.n1161 B.n87 10.6151
R2283 B.n1155 B.n87 10.6151
R2284 B.n1155 B.n1154 10.6151
R2285 B.n1154 B.n1153 10.6151
R2286 B.n1153 B.n94 10.6151
R2287 B.n1147 B.n94 10.6151
R2288 B.n1147 B.n1146 10.6151
R2289 B.n1146 B.n1145 10.6151
R2290 B.n1145 B.n101 10.6151
R2291 B.n1139 B.n101 10.6151
R2292 B.n1139 B.n1138 10.6151
R2293 B.n1138 B.n1137 10.6151
R2294 B.n1137 B.n108 10.6151
R2295 B.n1131 B.n108 10.6151
R2296 B.n1131 B.n1130 10.6151
R2297 B.n1130 B.n1129 10.6151
R2298 B.n290 B.n289 9.36635
R2299 B.n312 B.n311 9.36635
R2300 B.n718 B.n717 9.36635
R2301 B.n741 B.n575 9.36635
R2302 B.t8 B.n524 8.06834
R2303 B.t12 B.n99 8.06834
R2304 B.t1 B.n429 7.05986
R2305 B.t0 B.n15 7.05986
R2306 B.n500 B.t3 6.05138
R2307 B.t5 B.n1174 6.05138
R2308 B.n1257 B.n0 2.81026
R2309 B.n1257 B.n1 2.81026
R2310 B.n291 B.n290 1.24928
R2311 B.n311 B.n310 1.24928
R2312 B.n719 B.n718 1.24928
R2313 B.n576 B.n575 1.24928
R2314 VP.n24 VP.n23 161.3
R2315 VP.n25 VP.n20 161.3
R2316 VP.n27 VP.n26 161.3
R2317 VP.n28 VP.n19 161.3
R2318 VP.n30 VP.n29 161.3
R2319 VP.n31 VP.n18 161.3
R2320 VP.n34 VP.n33 161.3
R2321 VP.n35 VP.n17 161.3
R2322 VP.n37 VP.n36 161.3
R2323 VP.n38 VP.n16 161.3
R2324 VP.n40 VP.n39 161.3
R2325 VP.n41 VP.n15 161.3
R2326 VP.n43 VP.n42 161.3
R2327 VP.n44 VP.n14 161.3
R2328 VP.n46 VP.n45 161.3
R2329 VP.n85 VP.n84 161.3
R2330 VP.n83 VP.n1 161.3
R2331 VP.n82 VP.n81 161.3
R2332 VP.n80 VP.n2 161.3
R2333 VP.n79 VP.n78 161.3
R2334 VP.n77 VP.n3 161.3
R2335 VP.n76 VP.n75 161.3
R2336 VP.n74 VP.n4 161.3
R2337 VP.n73 VP.n72 161.3
R2338 VP.n70 VP.n5 161.3
R2339 VP.n69 VP.n68 161.3
R2340 VP.n67 VP.n6 161.3
R2341 VP.n66 VP.n65 161.3
R2342 VP.n64 VP.n7 161.3
R2343 VP.n63 VP.n62 161.3
R2344 VP.n61 VP.n60 161.3
R2345 VP.n59 VP.n9 161.3
R2346 VP.n58 VP.n57 161.3
R2347 VP.n56 VP.n10 161.3
R2348 VP.n55 VP.n54 161.3
R2349 VP.n53 VP.n11 161.3
R2350 VP.n52 VP.n51 161.3
R2351 VP.n50 VP.n12 161.3
R2352 VP.n22 VP.t5 148.102
R2353 VP.n48 VP.t1 114.544
R2354 VP.n8 VP.t4 114.544
R2355 VP.n71 VP.t3 114.544
R2356 VP.n0 VP.t7 114.544
R2357 VP.n13 VP.t6 114.544
R2358 VP.n32 VP.t0 114.544
R2359 VP.n21 VP.t2 114.544
R2360 VP.n49 VP.n48 79.6711
R2361 VP.n86 VP.n0 79.6711
R2362 VP.n47 VP.n13 79.6711
R2363 VP.n49 VP.n47 58.545
R2364 VP.n54 VP.n10 56.5617
R2365 VP.n78 VP.n2 56.5617
R2366 VP.n39 VP.n15 56.5617
R2367 VP.n22 VP.n21 54.9348
R2368 VP.n65 VP.n6 40.577
R2369 VP.n69 VP.n6 40.577
R2370 VP.n30 VP.n19 40.577
R2371 VP.n26 VP.n19 40.577
R2372 VP.n52 VP.n12 24.5923
R2373 VP.n53 VP.n52 24.5923
R2374 VP.n54 VP.n53 24.5923
R2375 VP.n58 VP.n10 24.5923
R2376 VP.n59 VP.n58 24.5923
R2377 VP.n60 VP.n59 24.5923
R2378 VP.n64 VP.n63 24.5923
R2379 VP.n65 VP.n64 24.5923
R2380 VP.n70 VP.n69 24.5923
R2381 VP.n72 VP.n70 24.5923
R2382 VP.n76 VP.n4 24.5923
R2383 VP.n77 VP.n76 24.5923
R2384 VP.n78 VP.n77 24.5923
R2385 VP.n82 VP.n2 24.5923
R2386 VP.n83 VP.n82 24.5923
R2387 VP.n84 VP.n83 24.5923
R2388 VP.n43 VP.n15 24.5923
R2389 VP.n44 VP.n43 24.5923
R2390 VP.n45 VP.n44 24.5923
R2391 VP.n31 VP.n30 24.5923
R2392 VP.n33 VP.n31 24.5923
R2393 VP.n37 VP.n17 24.5923
R2394 VP.n38 VP.n37 24.5923
R2395 VP.n39 VP.n38 24.5923
R2396 VP.n25 VP.n24 24.5923
R2397 VP.n26 VP.n25 24.5923
R2398 VP.n63 VP.n8 19.9199
R2399 VP.n72 VP.n71 19.9199
R2400 VP.n33 VP.n32 19.9199
R2401 VP.n24 VP.n21 19.9199
R2402 VP.n48 VP.n12 10.575
R2403 VP.n84 VP.n0 10.575
R2404 VP.n45 VP.n13 10.575
R2405 VP.n60 VP.n8 4.67295
R2406 VP.n71 VP.n4 4.67295
R2407 VP.n32 VP.n17 4.67295
R2408 VP.n23 VP.n22 3.1272
R2409 VP.n47 VP.n46 0.354861
R2410 VP.n50 VP.n49 0.354861
R2411 VP.n86 VP.n85 0.354861
R2412 VP VP.n86 0.267071
R2413 VP.n23 VP.n20 0.189894
R2414 VP.n27 VP.n20 0.189894
R2415 VP.n28 VP.n27 0.189894
R2416 VP.n29 VP.n28 0.189894
R2417 VP.n29 VP.n18 0.189894
R2418 VP.n34 VP.n18 0.189894
R2419 VP.n35 VP.n34 0.189894
R2420 VP.n36 VP.n35 0.189894
R2421 VP.n36 VP.n16 0.189894
R2422 VP.n40 VP.n16 0.189894
R2423 VP.n41 VP.n40 0.189894
R2424 VP.n42 VP.n41 0.189894
R2425 VP.n42 VP.n14 0.189894
R2426 VP.n46 VP.n14 0.189894
R2427 VP.n51 VP.n50 0.189894
R2428 VP.n51 VP.n11 0.189894
R2429 VP.n55 VP.n11 0.189894
R2430 VP.n56 VP.n55 0.189894
R2431 VP.n57 VP.n56 0.189894
R2432 VP.n57 VP.n9 0.189894
R2433 VP.n61 VP.n9 0.189894
R2434 VP.n62 VP.n61 0.189894
R2435 VP.n62 VP.n7 0.189894
R2436 VP.n66 VP.n7 0.189894
R2437 VP.n67 VP.n66 0.189894
R2438 VP.n68 VP.n67 0.189894
R2439 VP.n68 VP.n5 0.189894
R2440 VP.n73 VP.n5 0.189894
R2441 VP.n74 VP.n73 0.189894
R2442 VP.n75 VP.n74 0.189894
R2443 VP.n75 VP.n3 0.189894
R2444 VP.n79 VP.n3 0.189894
R2445 VP.n80 VP.n79 0.189894
R2446 VP.n81 VP.n80 0.189894
R2447 VP.n81 VP.n1 0.189894
R2448 VP.n85 VP.n1 0.189894
R2449 VDD1 VDD1.n0 64.3895
R2450 VDD1.n3 VDD1.n2 64.2757
R2451 VDD1.n3 VDD1.n1 64.2757
R2452 VDD1.n5 VDD1.n4 62.6889
R2453 VDD1.n5 VDD1.n3 53.3371
R2454 VDD1 VDD1.n5 1.58455
R2455 VDD1.n4 VDD1.t7 1.1976
R2456 VDD1.n4 VDD1.t1 1.1976
R2457 VDD1.n0 VDD1.t2 1.1976
R2458 VDD1.n0 VDD1.t5 1.1976
R2459 VDD1.n2 VDD1.t4 1.1976
R2460 VDD1.n2 VDD1.t0 1.1976
R2461 VDD1.n1 VDD1.t6 1.1976
R2462 VDD1.n1 VDD1.t3 1.1976
C0 VTAIL VP 12.9198f
C1 VTAIL VN 12.905701f
C2 VDD2 VP 0.613781f
C3 VDD2 VN 12.4186f
C4 VDD1 VP 12.876699f
C5 VDD1 VN 0.153788f
C6 VP VN 9.57336f
C7 VTAIL VDD2 9.7917f
C8 VTAIL VDD1 9.73138f
C9 VDD1 VDD2 2.23428f
C10 VDD2 B 6.61742f
C11 VDD1 B 7.148021f
C12 VTAIL B 13.81882f
C13 VN B 19.242477f
C14 VP B 17.84803f
C15 VDD1.t2 B 0.350048f
C16 VDD1.t5 B 0.350048f
C17 VDD1.n0 B 3.19758f
C18 VDD1.t6 B 0.350048f
C19 VDD1.t3 B 0.350048f
C20 VDD1.n1 B 3.19621f
C21 VDD1.t4 B 0.350048f
C22 VDD1.t0 B 0.350048f
C23 VDD1.n2 B 3.19621f
C24 VDD1.n3 B 4.41729f
C25 VDD1.t7 B 0.350048f
C26 VDD1.t1 B 0.350048f
C27 VDD1.n4 B 3.18014f
C28 VDD1.n5 B 3.88645f
C29 VP.t7 B 2.80781f
C30 VP.n0 B 1.03972f
C31 VP.n1 B 0.017765f
C32 VP.n2 B 0.022875f
C33 VP.n3 B 0.017765f
C34 VP.n4 B 0.01977f
C35 VP.n5 B 0.017765f
C36 VP.n6 B 0.014348f
C37 VP.n7 B 0.017765f
C38 VP.t4 B 2.80781f
C39 VP.n8 B 0.97145f
C40 VP.n9 B 0.017765f
C41 VP.n10 B 0.028772f
C42 VP.n11 B 0.017765f
C43 VP.n12 B 0.023673f
C44 VP.t6 B 2.80781f
C45 VP.n13 B 1.03972f
C46 VP.n14 B 0.017765f
C47 VP.n15 B 0.022875f
C48 VP.n16 B 0.017765f
C49 VP.n17 B 0.01977f
C50 VP.n18 B 0.017765f
C51 VP.n19 B 0.014348f
C52 VP.n20 B 0.017765f
C53 VP.t2 B 2.80781f
C54 VP.n21 B 1.03763f
C55 VP.t5 B 3.05785f
C56 VP.n22 B 0.986156f
C57 VP.n23 B 0.218775f
C58 VP.n24 B 0.029853f
C59 VP.n25 B 0.032943f
C60 VP.n26 B 0.035121f
C61 VP.n27 B 0.017765f
C62 VP.n28 B 0.017765f
C63 VP.n29 B 0.017765f
C64 VP.n30 B 0.035121f
C65 VP.n31 B 0.032943f
C66 VP.t0 B 2.80781f
C67 VP.n32 B 0.97145f
C68 VP.n33 B 0.029853f
C69 VP.n34 B 0.017765f
C70 VP.n35 B 0.017765f
C71 VP.n36 B 0.017765f
C72 VP.n37 B 0.032943f
C73 VP.n38 B 0.032943f
C74 VP.n39 B 0.028772f
C75 VP.n40 B 0.017765f
C76 VP.n41 B 0.017765f
C77 VP.n42 B 0.017765f
C78 VP.n43 B 0.032943f
C79 VP.n44 B 0.032943f
C80 VP.n45 B 0.023673f
C81 VP.n46 B 0.028667f
C82 VP.n47 B 1.26287f
C83 VP.t1 B 2.80781f
C84 VP.n48 B 1.03972f
C85 VP.n49 B 1.27381f
C86 VP.n50 B 0.028667f
C87 VP.n51 B 0.017765f
C88 VP.n52 B 0.032943f
C89 VP.n53 B 0.032943f
C90 VP.n54 B 0.022875f
C91 VP.n55 B 0.017765f
C92 VP.n56 B 0.017765f
C93 VP.n57 B 0.017765f
C94 VP.n58 B 0.032943f
C95 VP.n59 B 0.032943f
C96 VP.n60 B 0.01977f
C97 VP.n61 B 0.017765f
C98 VP.n62 B 0.017765f
C99 VP.n63 B 0.029853f
C100 VP.n64 B 0.032943f
C101 VP.n65 B 0.035121f
C102 VP.n66 B 0.017765f
C103 VP.n67 B 0.017765f
C104 VP.n68 B 0.017765f
C105 VP.n69 B 0.035121f
C106 VP.n70 B 0.032943f
C107 VP.t3 B 2.80781f
C108 VP.n71 B 0.97145f
C109 VP.n72 B 0.029853f
C110 VP.n73 B 0.017765f
C111 VP.n74 B 0.017765f
C112 VP.n75 B 0.017765f
C113 VP.n76 B 0.032943f
C114 VP.n77 B 0.032943f
C115 VP.n78 B 0.028772f
C116 VP.n79 B 0.017765f
C117 VP.n80 B 0.017765f
C118 VP.n81 B 0.017765f
C119 VP.n82 B 0.032943f
C120 VP.n83 B 0.032943f
C121 VP.n84 B 0.023673f
C122 VP.n85 B 0.028667f
C123 VP.n86 B 0.047159f
C124 VTAIL.t11 B 0.251718f
C125 VTAIL.t9 B 0.251718f
C126 VTAIL.n0 B 2.23113f
C127 VTAIL.n1 B 0.394257f
C128 VTAIL.t14 B 2.85003f
C129 VTAIL.n2 B 0.487406f
C130 VTAIL.t1 B 2.85003f
C131 VTAIL.n3 B 0.487406f
C132 VTAIL.t2 B 0.251718f
C133 VTAIL.t4 B 0.251718f
C134 VTAIL.n4 B 2.23113f
C135 VTAIL.n5 B 0.594466f
C136 VTAIL.t3 B 2.85003f
C137 VTAIL.n6 B 1.8085f
C138 VTAIL.t12 B 2.85003f
C139 VTAIL.n7 B 1.8085f
C140 VTAIL.t10 B 0.251718f
C141 VTAIL.t8 B 0.251718f
C142 VTAIL.n8 B 2.23114f
C143 VTAIL.n9 B 0.594464f
C144 VTAIL.t7 B 2.85003f
C145 VTAIL.n10 B 0.487403f
C146 VTAIL.t0 B 2.85003f
C147 VTAIL.n11 B 0.487403f
C148 VTAIL.t6 B 0.251718f
C149 VTAIL.t15 B 0.251718f
C150 VTAIL.n12 B 2.23114f
C151 VTAIL.n13 B 0.594464f
C152 VTAIL.t5 B 2.85003f
C153 VTAIL.n14 B 1.8085f
C154 VTAIL.t13 B 2.85003f
C155 VTAIL.n15 B 1.80489f
C156 VDD2.t2 B 0.345781f
C157 VDD2.t7 B 0.345781f
C158 VDD2.n0 B 3.15725f
C159 VDD2.t5 B 0.345781f
C160 VDD2.t1 B 0.345781f
C161 VDD2.n1 B 3.15725f
C162 VDD2.n2 B 4.30901f
C163 VDD2.t0 B 0.345781f
C164 VDD2.t6 B 0.345781f
C165 VDD2.n3 B 3.14139f
C166 VDD2.n4 B 3.80571f
C167 VDD2.t4 B 0.345781f
C168 VDD2.t3 B 0.345781f
C169 VDD2.n5 B 3.1572f
C170 VN.t1 B 2.7662f
C171 VN.n0 B 1.02431f
C172 VN.n1 B 0.017501f
C173 VN.n2 B 0.022536f
C174 VN.n3 B 0.017501f
C175 VN.n4 B 0.019477f
C176 VN.n5 B 0.017501f
C177 VN.n6 B 0.014135f
C178 VN.n7 B 0.017501f
C179 VN.t3 B 2.7662f
C180 VN.n8 B 1.02225f
C181 VN.t0 B 3.01254f
C182 VN.n9 B 0.971542f
C183 VN.n10 B 0.215533f
C184 VN.n11 B 0.02941f
C185 VN.n12 B 0.032454f
C186 VN.n13 B 0.034601f
C187 VN.n14 B 0.017501f
C188 VN.n15 B 0.017501f
C189 VN.n16 B 0.017501f
C190 VN.n17 B 0.034601f
C191 VN.n18 B 0.032454f
C192 VN.t5 B 2.7662f
C193 VN.n19 B 0.957054f
C194 VN.n20 B 0.02941f
C195 VN.n21 B 0.017501f
C196 VN.n22 B 0.017501f
C197 VN.n23 B 0.017501f
C198 VN.n24 B 0.032454f
C199 VN.n25 B 0.032454f
C200 VN.n26 B 0.028346f
C201 VN.n27 B 0.017501f
C202 VN.n28 B 0.017501f
C203 VN.n29 B 0.017501f
C204 VN.n30 B 0.032454f
C205 VN.n31 B 0.032454f
C206 VN.n32 B 0.023322f
C207 VN.n33 B 0.028242f
C208 VN.n34 B 0.04646f
C209 VN.t2 B 2.7662f
C210 VN.n35 B 1.02431f
C211 VN.n36 B 0.017501f
C212 VN.n37 B 0.022536f
C213 VN.n38 B 0.017501f
C214 VN.n39 B 0.019477f
C215 VN.n40 B 0.017501f
C216 VN.t4 B 2.7662f
C217 VN.n41 B 0.957054f
C218 VN.n42 B 0.014135f
C219 VN.n43 B 0.017501f
C220 VN.t6 B 2.7662f
C221 VN.n44 B 1.02225f
C222 VN.t7 B 3.01254f
C223 VN.n45 B 0.971542f
C224 VN.n46 B 0.215533f
C225 VN.n47 B 0.02941f
C226 VN.n48 B 0.032454f
C227 VN.n49 B 0.034601f
C228 VN.n50 B 0.017501f
C229 VN.n51 B 0.017501f
C230 VN.n52 B 0.017501f
C231 VN.n53 B 0.034601f
C232 VN.n54 B 0.032454f
C233 VN.n55 B 0.02941f
C234 VN.n56 B 0.017501f
C235 VN.n57 B 0.017501f
C236 VN.n58 B 0.017501f
C237 VN.n59 B 0.032454f
C238 VN.n60 B 0.032454f
C239 VN.n61 B 0.028346f
C240 VN.n62 B 0.017501f
C241 VN.n63 B 0.017501f
C242 VN.n64 B 0.017501f
C243 VN.n65 B 0.032454f
C244 VN.n66 B 0.032454f
C245 VN.n67 B 0.023322f
C246 VN.n68 B 0.028242f
C247 VN.n69 B 1.25095f
.ends

