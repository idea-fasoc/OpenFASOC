* NGSPICE file created from diff_pair_sample_0837.ext - technology: sky130A

.subckt diff_pair_sample_0837 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t10 w_n4090_n2088# sky130_fd_pr__pfet_01v8 ad=0.924 pd=5.93 as=2.184 ps=11.98 w=5.6 l=2.79
X1 VTAIL.t13 VN.t1 VDD2.t6 w_n4090_n2088# sky130_fd_pr__pfet_01v8 ad=2.184 pd=11.98 as=0.924 ps=5.93 w=5.6 l=2.79
X2 VDD1.t7 VP.t0 VTAIL.t7 w_n4090_n2088# sky130_fd_pr__pfet_01v8 ad=0.924 pd=5.93 as=2.184 ps=11.98 w=5.6 l=2.79
X3 VDD2.t5 VN.t2 VTAIL.t11 w_n4090_n2088# sky130_fd_pr__pfet_01v8 ad=0.924 pd=5.93 as=0.924 ps=5.93 w=5.6 l=2.79
X4 VDD2.t4 VN.t3 VTAIL.t9 w_n4090_n2088# sky130_fd_pr__pfet_01v8 ad=0.924 pd=5.93 as=2.184 ps=11.98 w=5.6 l=2.79
X5 VDD1.t6 VP.t1 VTAIL.t3 w_n4090_n2088# sky130_fd_pr__pfet_01v8 ad=0.924 pd=5.93 as=0.924 ps=5.93 w=5.6 l=2.79
X6 VTAIL.t0 VP.t2 VDD1.t5 w_n4090_n2088# sky130_fd_pr__pfet_01v8 ad=0.924 pd=5.93 as=0.924 ps=5.93 w=5.6 l=2.79
X7 B.t11 B.t9 B.t10 w_n4090_n2088# sky130_fd_pr__pfet_01v8 ad=2.184 pd=11.98 as=0 ps=0 w=5.6 l=2.79
X8 VTAIL.t14 VN.t4 VDD2.t3 w_n4090_n2088# sky130_fd_pr__pfet_01v8 ad=0.924 pd=5.93 as=0.924 ps=5.93 w=5.6 l=2.79
X9 B.t8 B.t6 B.t7 w_n4090_n2088# sky130_fd_pr__pfet_01v8 ad=2.184 pd=11.98 as=0 ps=0 w=5.6 l=2.79
X10 VTAIL.t8 VN.t5 VDD2.t2 w_n4090_n2088# sky130_fd_pr__pfet_01v8 ad=2.184 pd=11.98 as=0.924 ps=5.93 w=5.6 l=2.79
X11 VDD1.t4 VP.t3 VTAIL.t6 w_n4090_n2088# sky130_fd_pr__pfet_01v8 ad=0.924 pd=5.93 as=2.184 ps=11.98 w=5.6 l=2.79
X12 VTAIL.t15 VN.t6 VDD2.t1 w_n4090_n2088# sky130_fd_pr__pfet_01v8 ad=0.924 pd=5.93 as=0.924 ps=5.93 w=5.6 l=2.79
X13 VDD2.t0 VN.t7 VTAIL.t12 w_n4090_n2088# sky130_fd_pr__pfet_01v8 ad=0.924 pd=5.93 as=0.924 ps=5.93 w=5.6 l=2.79
X14 VDD1.t3 VP.t4 VTAIL.t1 w_n4090_n2088# sky130_fd_pr__pfet_01v8 ad=0.924 pd=5.93 as=0.924 ps=5.93 w=5.6 l=2.79
X15 VTAIL.t5 VP.t5 VDD1.t2 w_n4090_n2088# sky130_fd_pr__pfet_01v8 ad=2.184 pd=11.98 as=0.924 ps=5.93 w=5.6 l=2.79
X16 VTAIL.t4 VP.t6 VDD1.t1 w_n4090_n2088# sky130_fd_pr__pfet_01v8 ad=0.924 pd=5.93 as=0.924 ps=5.93 w=5.6 l=2.79
X17 B.t5 B.t3 B.t4 w_n4090_n2088# sky130_fd_pr__pfet_01v8 ad=2.184 pd=11.98 as=0 ps=0 w=5.6 l=2.79
X18 B.t2 B.t0 B.t1 w_n4090_n2088# sky130_fd_pr__pfet_01v8 ad=2.184 pd=11.98 as=0 ps=0 w=5.6 l=2.79
X19 VTAIL.t2 VP.t7 VDD1.t0 w_n4090_n2088# sky130_fd_pr__pfet_01v8 ad=2.184 pd=11.98 as=0.924 ps=5.93 w=5.6 l=2.79
R0 VN.n56 VN.n55 161.3
R1 VN.n54 VN.n30 161.3
R2 VN.n53 VN.n52 161.3
R3 VN.n51 VN.n31 161.3
R4 VN.n50 VN.n49 161.3
R5 VN.n48 VN.n32 161.3
R6 VN.n46 VN.n45 161.3
R7 VN.n44 VN.n33 161.3
R8 VN.n43 VN.n42 161.3
R9 VN.n41 VN.n34 161.3
R10 VN.n40 VN.n39 161.3
R11 VN.n38 VN.n35 161.3
R12 VN.n27 VN.n26 161.3
R13 VN.n25 VN.n1 161.3
R14 VN.n24 VN.n23 161.3
R15 VN.n22 VN.n2 161.3
R16 VN.n21 VN.n20 161.3
R17 VN.n19 VN.n3 161.3
R18 VN.n17 VN.n16 161.3
R19 VN.n15 VN.n4 161.3
R20 VN.n14 VN.n13 161.3
R21 VN.n12 VN.n5 161.3
R22 VN.n11 VN.n10 161.3
R23 VN.n9 VN.n6 161.3
R24 VN.n37 VN.t3 80.293
R25 VN.n8 VN.t1 80.293
R26 VN.n28 VN.n0 69.0966
R27 VN.n57 VN.n29 69.0966
R28 VN.n8 VN.n7 58.6055
R29 VN.n37 VN.n36 58.6055
R30 VN.n13 VN.n12 56.5617
R31 VN.n42 VN.n41 56.5617
R32 VN.n24 VN.n2 53.171
R33 VN.n53 VN.n31 53.171
R34 VN.n7 VN.t7 48.3733
R35 VN.n18 VN.t4 48.3733
R36 VN.n0 VN.t0 48.3733
R37 VN.n36 VN.t6 48.3733
R38 VN.n47 VN.t2 48.3733
R39 VN.n29 VN.t5 48.3733
R40 VN VN.n57 47.1875
R41 VN.n25 VN.n24 27.983
R42 VN.n54 VN.n53 27.983
R43 VN.n11 VN.n6 24.5923
R44 VN.n12 VN.n11 24.5923
R45 VN.n13 VN.n4 24.5923
R46 VN.n17 VN.n4 24.5923
R47 VN.n20 VN.n19 24.5923
R48 VN.n20 VN.n2 24.5923
R49 VN.n26 VN.n25 24.5923
R50 VN.n41 VN.n40 24.5923
R51 VN.n40 VN.n35 24.5923
R52 VN.n49 VN.n31 24.5923
R53 VN.n49 VN.n48 24.5923
R54 VN.n46 VN.n33 24.5923
R55 VN.n42 VN.n33 24.5923
R56 VN.n55 VN.n54 24.5923
R57 VN.n26 VN.n0 21.1495
R58 VN.n55 VN.n29 21.1495
R59 VN.n7 VN.n6 15.2474
R60 VN.n18 VN.n17 15.2474
R61 VN.n36 VN.n35 15.2474
R62 VN.n47 VN.n46 15.2474
R63 VN.n19 VN.n18 9.3454
R64 VN.n48 VN.n47 9.3454
R65 VN.n38 VN.n37 5.4467
R66 VN.n9 VN.n8 5.4467
R67 VN.n57 VN.n56 0.354861
R68 VN.n28 VN.n27 0.354861
R69 VN VN.n28 0.267071
R70 VN.n56 VN.n30 0.189894
R71 VN.n52 VN.n30 0.189894
R72 VN.n52 VN.n51 0.189894
R73 VN.n51 VN.n50 0.189894
R74 VN.n50 VN.n32 0.189894
R75 VN.n45 VN.n32 0.189894
R76 VN.n45 VN.n44 0.189894
R77 VN.n44 VN.n43 0.189894
R78 VN.n43 VN.n34 0.189894
R79 VN.n39 VN.n34 0.189894
R80 VN.n39 VN.n38 0.189894
R81 VN.n10 VN.n9 0.189894
R82 VN.n10 VN.n5 0.189894
R83 VN.n14 VN.n5 0.189894
R84 VN.n15 VN.n14 0.189894
R85 VN.n16 VN.n15 0.189894
R86 VN.n16 VN.n3 0.189894
R87 VN.n21 VN.n3 0.189894
R88 VN.n22 VN.n21 0.189894
R89 VN.n23 VN.n22 0.189894
R90 VN.n23 VN.n1 0.189894
R91 VN.n27 VN.n1 0.189894
R92 VTAIL.n11 VTAIL.t2 82.9904
R93 VTAIL.n10 VTAIL.t9 82.9904
R94 VTAIL.n7 VTAIL.t8 82.9904
R95 VTAIL.n14 VTAIL.t7 82.9902
R96 VTAIL.n15 VTAIL.t10 82.9902
R97 VTAIL.n2 VTAIL.t13 82.9902
R98 VTAIL.n3 VTAIL.t6 82.9902
R99 VTAIL.n6 VTAIL.t5 82.9902
R100 VTAIL.n13 VTAIL.n12 77.186
R101 VTAIL.n9 VTAIL.n8 77.186
R102 VTAIL.n1 VTAIL.n0 77.1857
R103 VTAIL.n5 VTAIL.n4 77.1857
R104 VTAIL.n15 VTAIL.n14 19.8841
R105 VTAIL.n7 VTAIL.n6 19.8841
R106 VTAIL.n0 VTAIL.t12 5.80496
R107 VTAIL.n0 VTAIL.t14 5.80496
R108 VTAIL.n4 VTAIL.t1 5.80496
R109 VTAIL.n4 VTAIL.t0 5.80496
R110 VTAIL.n12 VTAIL.t3 5.80496
R111 VTAIL.n12 VTAIL.t4 5.80496
R112 VTAIL.n8 VTAIL.t11 5.80496
R113 VTAIL.n8 VTAIL.t15 5.80496
R114 VTAIL.n9 VTAIL.n7 2.69016
R115 VTAIL.n10 VTAIL.n9 2.69016
R116 VTAIL.n13 VTAIL.n11 2.69016
R117 VTAIL.n14 VTAIL.n13 2.69016
R118 VTAIL.n6 VTAIL.n5 2.69016
R119 VTAIL.n5 VTAIL.n3 2.69016
R120 VTAIL.n2 VTAIL.n1 2.69016
R121 VTAIL VTAIL.n15 2.63197
R122 VTAIL.n11 VTAIL.n10 0.470328
R123 VTAIL.n3 VTAIL.n2 0.470328
R124 VTAIL VTAIL.n1 0.0586897
R125 VDD2.n2 VDD2.n1 95.154
R126 VDD2.n2 VDD2.n0 95.154
R127 VDD2 VDD2.n5 95.1512
R128 VDD2.n4 VDD2.n3 93.8648
R129 VDD2.n4 VDD2.n2 40.6463
R130 VDD2.n5 VDD2.t1 5.80496
R131 VDD2.n5 VDD2.t4 5.80496
R132 VDD2.n3 VDD2.t2 5.80496
R133 VDD2.n3 VDD2.t5 5.80496
R134 VDD2.n1 VDD2.t3 5.80496
R135 VDD2.n1 VDD2.t7 5.80496
R136 VDD2.n0 VDD2.t6 5.80496
R137 VDD2.n0 VDD2.t0 5.80496
R138 VDD2 VDD2.n4 1.40352
R139 VP.n19 VP.n16 161.3
R140 VP.n21 VP.n20 161.3
R141 VP.n22 VP.n15 161.3
R142 VP.n24 VP.n23 161.3
R143 VP.n25 VP.n14 161.3
R144 VP.n27 VP.n26 161.3
R145 VP.n29 VP.n13 161.3
R146 VP.n31 VP.n30 161.3
R147 VP.n32 VP.n12 161.3
R148 VP.n34 VP.n33 161.3
R149 VP.n35 VP.n11 161.3
R150 VP.n37 VP.n36 161.3
R151 VP.n69 VP.n68 161.3
R152 VP.n67 VP.n1 161.3
R153 VP.n66 VP.n65 161.3
R154 VP.n64 VP.n2 161.3
R155 VP.n63 VP.n62 161.3
R156 VP.n61 VP.n3 161.3
R157 VP.n59 VP.n58 161.3
R158 VP.n57 VP.n4 161.3
R159 VP.n56 VP.n55 161.3
R160 VP.n54 VP.n5 161.3
R161 VP.n53 VP.n52 161.3
R162 VP.n51 VP.n6 161.3
R163 VP.n50 VP.n49 161.3
R164 VP.n47 VP.n7 161.3
R165 VP.n46 VP.n45 161.3
R166 VP.n44 VP.n8 161.3
R167 VP.n43 VP.n42 161.3
R168 VP.n41 VP.n9 161.3
R169 VP.n18 VP.t7 80.2928
R170 VP.n40 VP.n39 69.0966
R171 VP.n70 VP.n0 69.0966
R172 VP.n38 VP.n10 69.0966
R173 VP.n18 VP.n17 58.6055
R174 VP.n55 VP.n54 56.5617
R175 VP.n23 VP.n22 56.5617
R176 VP.n46 VP.n8 53.171
R177 VP.n66 VP.n2 53.171
R178 VP.n34 VP.n12 53.171
R179 VP.n40 VP.t5 48.3733
R180 VP.n48 VP.t4 48.3733
R181 VP.n60 VP.t2 48.3733
R182 VP.n0 VP.t3 48.3733
R183 VP.n10 VP.t0 48.3733
R184 VP.n28 VP.t6 48.3733
R185 VP.n17 VP.t1 48.3733
R186 VP.n39 VP.n38 47.0223
R187 VP.n42 VP.n8 27.983
R188 VP.n67 VP.n66 27.983
R189 VP.n35 VP.n34 27.983
R190 VP.n42 VP.n41 24.5923
R191 VP.n47 VP.n46 24.5923
R192 VP.n49 VP.n47 24.5923
R193 VP.n53 VP.n6 24.5923
R194 VP.n54 VP.n53 24.5923
R195 VP.n55 VP.n4 24.5923
R196 VP.n59 VP.n4 24.5923
R197 VP.n62 VP.n61 24.5923
R198 VP.n62 VP.n2 24.5923
R199 VP.n68 VP.n67 24.5923
R200 VP.n36 VP.n35 24.5923
R201 VP.n23 VP.n14 24.5923
R202 VP.n27 VP.n14 24.5923
R203 VP.n30 VP.n29 24.5923
R204 VP.n30 VP.n12 24.5923
R205 VP.n21 VP.n16 24.5923
R206 VP.n22 VP.n21 24.5923
R207 VP.n41 VP.n40 21.1495
R208 VP.n68 VP.n0 21.1495
R209 VP.n36 VP.n10 21.1495
R210 VP.n48 VP.n6 15.2474
R211 VP.n60 VP.n59 15.2474
R212 VP.n28 VP.n27 15.2474
R213 VP.n17 VP.n16 15.2474
R214 VP.n49 VP.n48 9.3454
R215 VP.n61 VP.n60 9.3454
R216 VP.n29 VP.n28 9.3454
R217 VP.n19 VP.n18 5.44666
R218 VP.n38 VP.n37 0.354861
R219 VP.n39 VP.n9 0.354861
R220 VP.n70 VP.n69 0.354861
R221 VP VP.n70 0.267071
R222 VP.n20 VP.n19 0.189894
R223 VP.n20 VP.n15 0.189894
R224 VP.n24 VP.n15 0.189894
R225 VP.n25 VP.n24 0.189894
R226 VP.n26 VP.n25 0.189894
R227 VP.n26 VP.n13 0.189894
R228 VP.n31 VP.n13 0.189894
R229 VP.n32 VP.n31 0.189894
R230 VP.n33 VP.n32 0.189894
R231 VP.n33 VP.n11 0.189894
R232 VP.n37 VP.n11 0.189894
R233 VP.n43 VP.n9 0.189894
R234 VP.n44 VP.n43 0.189894
R235 VP.n45 VP.n44 0.189894
R236 VP.n45 VP.n7 0.189894
R237 VP.n50 VP.n7 0.189894
R238 VP.n51 VP.n50 0.189894
R239 VP.n52 VP.n51 0.189894
R240 VP.n52 VP.n5 0.189894
R241 VP.n56 VP.n5 0.189894
R242 VP.n57 VP.n56 0.189894
R243 VP.n58 VP.n57 0.189894
R244 VP.n58 VP.n3 0.189894
R245 VP.n63 VP.n3 0.189894
R246 VP.n64 VP.n63 0.189894
R247 VP.n65 VP.n64 0.189894
R248 VP.n65 VP.n1 0.189894
R249 VP.n69 VP.n1 0.189894
R250 VDD1 VDD1.n0 95.2678
R251 VDD1.n3 VDD1.n2 95.154
R252 VDD1.n3 VDD1.n1 95.154
R253 VDD1.n5 VDD1.n4 93.8646
R254 VDD1.n5 VDD1.n3 41.2293
R255 VDD1.n4 VDD1.t1 5.80496
R256 VDD1.n4 VDD1.t7 5.80496
R257 VDD1.n0 VDD1.t0 5.80496
R258 VDD1.n0 VDD1.t6 5.80496
R259 VDD1.n2 VDD1.t5 5.80496
R260 VDD1.n2 VDD1.t4 5.80496
R261 VDD1.n1 VDD1.t2 5.80496
R262 VDD1.n1 VDD1.t3 5.80496
R263 VDD1 VDD1.n5 1.28714
R264 B.n502 B.n61 585
R265 B.n504 B.n503 585
R266 B.n505 B.n60 585
R267 B.n507 B.n506 585
R268 B.n508 B.n59 585
R269 B.n510 B.n509 585
R270 B.n511 B.n58 585
R271 B.n513 B.n512 585
R272 B.n514 B.n57 585
R273 B.n516 B.n515 585
R274 B.n517 B.n56 585
R275 B.n519 B.n518 585
R276 B.n520 B.n55 585
R277 B.n522 B.n521 585
R278 B.n523 B.n54 585
R279 B.n525 B.n524 585
R280 B.n526 B.n53 585
R281 B.n528 B.n527 585
R282 B.n529 B.n52 585
R283 B.n531 B.n530 585
R284 B.n532 B.n51 585
R285 B.n534 B.n533 585
R286 B.n535 B.n48 585
R287 B.n538 B.n537 585
R288 B.n539 B.n47 585
R289 B.n541 B.n540 585
R290 B.n542 B.n46 585
R291 B.n544 B.n543 585
R292 B.n545 B.n45 585
R293 B.n547 B.n546 585
R294 B.n548 B.n41 585
R295 B.n550 B.n549 585
R296 B.n551 B.n40 585
R297 B.n553 B.n552 585
R298 B.n554 B.n39 585
R299 B.n556 B.n555 585
R300 B.n557 B.n38 585
R301 B.n559 B.n558 585
R302 B.n560 B.n37 585
R303 B.n562 B.n561 585
R304 B.n563 B.n36 585
R305 B.n565 B.n564 585
R306 B.n566 B.n35 585
R307 B.n568 B.n567 585
R308 B.n569 B.n34 585
R309 B.n571 B.n570 585
R310 B.n572 B.n33 585
R311 B.n574 B.n573 585
R312 B.n575 B.n32 585
R313 B.n577 B.n576 585
R314 B.n578 B.n31 585
R315 B.n580 B.n579 585
R316 B.n581 B.n30 585
R317 B.n583 B.n582 585
R318 B.n584 B.n29 585
R319 B.n501 B.n500 585
R320 B.n499 B.n62 585
R321 B.n498 B.n497 585
R322 B.n496 B.n63 585
R323 B.n495 B.n494 585
R324 B.n493 B.n64 585
R325 B.n492 B.n491 585
R326 B.n490 B.n65 585
R327 B.n489 B.n488 585
R328 B.n487 B.n66 585
R329 B.n486 B.n485 585
R330 B.n484 B.n67 585
R331 B.n483 B.n482 585
R332 B.n481 B.n68 585
R333 B.n480 B.n479 585
R334 B.n478 B.n69 585
R335 B.n477 B.n476 585
R336 B.n475 B.n70 585
R337 B.n474 B.n473 585
R338 B.n472 B.n71 585
R339 B.n471 B.n470 585
R340 B.n469 B.n72 585
R341 B.n468 B.n467 585
R342 B.n466 B.n73 585
R343 B.n465 B.n464 585
R344 B.n463 B.n74 585
R345 B.n462 B.n461 585
R346 B.n460 B.n75 585
R347 B.n459 B.n458 585
R348 B.n457 B.n76 585
R349 B.n456 B.n455 585
R350 B.n454 B.n77 585
R351 B.n453 B.n452 585
R352 B.n451 B.n78 585
R353 B.n450 B.n449 585
R354 B.n448 B.n79 585
R355 B.n447 B.n446 585
R356 B.n445 B.n80 585
R357 B.n444 B.n443 585
R358 B.n442 B.n81 585
R359 B.n441 B.n440 585
R360 B.n439 B.n82 585
R361 B.n438 B.n437 585
R362 B.n436 B.n83 585
R363 B.n435 B.n434 585
R364 B.n433 B.n84 585
R365 B.n432 B.n431 585
R366 B.n430 B.n85 585
R367 B.n429 B.n428 585
R368 B.n427 B.n86 585
R369 B.n426 B.n425 585
R370 B.n424 B.n87 585
R371 B.n423 B.n422 585
R372 B.n421 B.n88 585
R373 B.n420 B.n419 585
R374 B.n418 B.n89 585
R375 B.n417 B.n416 585
R376 B.n415 B.n90 585
R377 B.n414 B.n413 585
R378 B.n412 B.n91 585
R379 B.n411 B.n410 585
R380 B.n409 B.n92 585
R381 B.n408 B.n407 585
R382 B.n406 B.n93 585
R383 B.n405 B.n404 585
R384 B.n403 B.n94 585
R385 B.n402 B.n401 585
R386 B.n400 B.n95 585
R387 B.n399 B.n398 585
R388 B.n397 B.n96 585
R389 B.n396 B.n395 585
R390 B.n394 B.n97 585
R391 B.n393 B.n392 585
R392 B.n391 B.n98 585
R393 B.n390 B.n389 585
R394 B.n388 B.n99 585
R395 B.n387 B.n386 585
R396 B.n385 B.n100 585
R397 B.n384 B.n383 585
R398 B.n382 B.n101 585
R399 B.n381 B.n380 585
R400 B.n379 B.n102 585
R401 B.n378 B.n377 585
R402 B.n376 B.n103 585
R403 B.n375 B.n374 585
R404 B.n373 B.n104 585
R405 B.n372 B.n371 585
R406 B.n370 B.n105 585
R407 B.n369 B.n368 585
R408 B.n367 B.n106 585
R409 B.n366 B.n365 585
R410 B.n364 B.n107 585
R411 B.n363 B.n362 585
R412 B.n361 B.n108 585
R413 B.n360 B.n359 585
R414 B.n358 B.n109 585
R415 B.n357 B.n356 585
R416 B.n355 B.n110 585
R417 B.n354 B.n353 585
R418 B.n352 B.n111 585
R419 B.n351 B.n350 585
R420 B.n349 B.n112 585
R421 B.n348 B.n347 585
R422 B.n346 B.n113 585
R423 B.n345 B.n344 585
R424 B.n343 B.n114 585
R425 B.n342 B.n341 585
R426 B.n340 B.n115 585
R427 B.n339 B.n338 585
R428 B.n252 B.n145 585
R429 B.n254 B.n253 585
R430 B.n255 B.n144 585
R431 B.n257 B.n256 585
R432 B.n258 B.n143 585
R433 B.n260 B.n259 585
R434 B.n261 B.n142 585
R435 B.n263 B.n262 585
R436 B.n264 B.n141 585
R437 B.n266 B.n265 585
R438 B.n267 B.n140 585
R439 B.n269 B.n268 585
R440 B.n270 B.n139 585
R441 B.n272 B.n271 585
R442 B.n273 B.n138 585
R443 B.n275 B.n274 585
R444 B.n276 B.n137 585
R445 B.n278 B.n277 585
R446 B.n279 B.n136 585
R447 B.n281 B.n280 585
R448 B.n282 B.n135 585
R449 B.n284 B.n283 585
R450 B.n285 B.n132 585
R451 B.n288 B.n287 585
R452 B.n289 B.n131 585
R453 B.n291 B.n290 585
R454 B.n292 B.n130 585
R455 B.n294 B.n293 585
R456 B.n295 B.n129 585
R457 B.n297 B.n296 585
R458 B.n298 B.n128 585
R459 B.n303 B.n302 585
R460 B.n304 B.n127 585
R461 B.n306 B.n305 585
R462 B.n307 B.n126 585
R463 B.n309 B.n308 585
R464 B.n310 B.n125 585
R465 B.n312 B.n311 585
R466 B.n313 B.n124 585
R467 B.n315 B.n314 585
R468 B.n316 B.n123 585
R469 B.n318 B.n317 585
R470 B.n319 B.n122 585
R471 B.n321 B.n320 585
R472 B.n322 B.n121 585
R473 B.n324 B.n323 585
R474 B.n325 B.n120 585
R475 B.n327 B.n326 585
R476 B.n328 B.n119 585
R477 B.n330 B.n329 585
R478 B.n331 B.n118 585
R479 B.n333 B.n332 585
R480 B.n334 B.n117 585
R481 B.n336 B.n335 585
R482 B.n337 B.n116 585
R483 B.n251 B.n250 585
R484 B.n249 B.n146 585
R485 B.n248 B.n247 585
R486 B.n246 B.n147 585
R487 B.n245 B.n244 585
R488 B.n243 B.n148 585
R489 B.n242 B.n241 585
R490 B.n240 B.n149 585
R491 B.n239 B.n238 585
R492 B.n237 B.n150 585
R493 B.n236 B.n235 585
R494 B.n234 B.n151 585
R495 B.n233 B.n232 585
R496 B.n231 B.n152 585
R497 B.n230 B.n229 585
R498 B.n228 B.n153 585
R499 B.n227 B.n226 585
R500 B.n225 B.n154 585
R501 B.n224 B.n223 585
R502 B.n222 B.n155 585
R503 B.n221 B.n220 585
R504 B.n219 B.n156 585
R505 B.n218 B.n217 585
R506 B.n216 B.n157 585
R507 B.n215 B.n214 585
R508 B.n213 B.n158 585
R509 B.n212 B.n211 585
R510 B.n210 B.n159 585
R511 B.n209 B.n208 585
R512 B.n207 B.n160 585
R513 B.n206 B.n205 585
R514 B.n204 B.n161 585
R515 B.n203 B.n202 585
R516 B.n201 B.n162 585
R517 B.n200 B.n199 585
R518 B.n198 B.n163 585
R519 B.n197 B.n196 585
R520 B.n195 B.n164 585
R521 B.n194 B.n193 585
R522 B.n192 B.n165 585
R523 B.n191 B.n190 585
R524 B.n189 B.n166 585
R525 B.n188 B.n187 585
R526 B.n186 B.n167 585
R527 B.n185 B.n184 585
R528 B.n183 B.n168 585
R529 B.n182 B.n181 585
R530 B.n180 B.n169 585
R531 B.n179 B.n178 585
R532 B.n177 B.n170 585
R533 B.n176 B.n175 585
R534 B.n174 B.n171 585
R535 B.n173 B.n172 585
R536 B.n2 B.n0 585
R537 B.n665 B.n1 585
R538 B.n664 B.n663 585
R539 B.n662 B.n3 585
R540 B.n661 B.n660 585
R541 B.n659 B.n4 585
R542 B.n658 B.n657 585
R543 B.n656 B.n5 585
R544 B.n655 B.n654 585
R545 B.n653 B.n6 585
R546 B.n652 B.n651 585
R547 B.n650 B.n7 585
R548 B.n649 B.n648 585
R549 B.n647 B.n8 585
R550 B.n646 B.n645 585
R551 B.n644 B.n9 585
R552 B.n643 B.n642 585
R553 B.n641 B.n10 585
R554 B.n640 B.n639 585
R555 B.n638 B.n11 585
R556 B.n637 B.n636 585
R557 B.n635 B.n12 585
R558 B.n634 B.n633 585
R559 B.n632 B.n13 585
R560 B.n631 B.n630 585
R561 B.n629 B.n14 585
R562 B.n628 B.n627 585
R563 B.n626 B.n15 585
R564 B.n625 B.n624 585
R565 B.n623 B.n16 585
R566 B.n622 B.n621 585
R567 B.n620 B.n17 585
R568 B.n619 B.n618 585
R569 B.n617 B.n18 585
R570 B.n616 B.n615 585
R571 B.n614 B.n19 585
R572 B.n613 B.n612 585
R573 B.n611 B.n20 585
R574 B.n610 B.n609 585
R575 B.n608 B.n21 585
R576 B.n607 B.n606 585
R577 B.n605 B.n22 585
R578 B.n604 B.n603 585
R579 B.n602 B.n23 585
R580 B.n601 B.n600 585
R581 B.n599 B.n24 585
R582 B.n598 B.n597 585
R583 B.n596 B.n25 585
R584 B.n595 B.n594 585
R585 B.n593 B.n26 585
R586 B.n592 B.n591 585
R587 B.n590 B.n27 585
R588 B.n589 B.n588 585
R589 B.n587 B.n28 585
R590 B.n586 B.n585 585
R591 B.n667 B.n666 585
R592 B.n252 B.n251 511.721
R593 B.n586 B.n29 511.721
R594 B.n339 B.n116 511.721
R595 B.n502 B.n501 511.721
R596 B.n299 B.t9 256.69
R597 B.n133 B.t6 256.69
R598 B.n42 B.t0 256.69
R599 B.n49 B.t3 256.69
R600 B.n299 B.t11 175.775
R601 B.n49 B.t4 175.775
R602 B.n133 B.t8 175.77
R603 B.n42 B.t1 175.77
R604 B.n251 B.n146 163.367
R605 B.n247 B.n146 163.367
R606 B.n247 B.n246 163.367
R607 B.n246 B.n245 163.367
R608 B.n245 B.n148 163.367
R609 B.n241 B.n148 163.367
R610 B.n241 B.n240 163.367
R611 B.n240 B.n239 163.367
R612 B.n239 B.n150 163.367
R613 B.n235 B.n150 163.367
R614 B.n235 B.n234 163.367
R615 B.n234 B.n233 163.367
R616 B.n233 B.n152 163.367
R617 B.n229 B.n152 163.367
R618 B.n229 B.n228 163.367
R619 B.n228 B.n227 163.367
R620 B.n227 B.n154 163.367
R621 B.n223 B.n154 163.367
R622 B.n223 B.n222 163.367
R623 B.n222 B.n221 163.367
R624 B.n221 B.n156 163.367
R625 B.n217 B.n156 163.367
R626 B.n217 B.n216 163.367
R627 B.n216 B.n215 163.367
R628 B.n215 B.n158 163.367
R629 B.n211 B.n158 163.367
R630 B.n211 B.n210 163.367
R631 B.n210 B.n209 163.367
R632 B.n209 B.n160 163.367
R633 B.n205 B.n160 163.367
R634 B.n205 B.n204 163.367
R635 B.n204 B.n203 163.367
R636 B.n203 B.n162 163.367
R637 B.n199 B.n162 163.367
R638 B.n199 B.n198 163.367
R639 B.n198 B.n197 163.367
R640 B.n197 B.n164 163.367
R641 B.n193 B.n164 163.367
R642 B.n193 B.n192 163.367
R643 B.n192 B.n191 163.367
R644 B.n191 B.n166 163.367
R645 B.n187 B.n166 163.367
R646 B.n187 B.n186 163.367
R647 B.n186 B.n185 163.367
R648 B.n185 B.n168 163.367
R649 B.n181 B.n168 163.367
R650 B.n181 B.n180 163.367
R651 B.n180 B.n179 163.367
R652 B.n179 B.n170 163.367
R653 B.n175 B.n170 163.367
R654 B.n175 B.n174 163.367
R655 B.n174 B.n173 163.367
R656 B.n173 B.n2 163.367
R657 B.n666 B.n2 163.367
R658 B.n666 B.n665 163.367
R659 B.n665 B.n664 163.367
R660 B.n664 B.n3 163.367
R661 B.n660 B.n3 163.367
R662 B.n660 B.n659 163.367
R663 B.n659 B.n658 163.367
R664 B.n658 B.n5 163.367
R665 B.n654 B.n5 163.367
R666 B.n654 B.n653 163.367
R667 B.n653 B.n652 163.367
R668 B.n652 B.n7 163.367
R669 B.n648 B.n7 163.367
R670 B.n648 B.n647 163.367
R671 B.n647 B.n646 163.367
R672 B.n646 B.n9 163.367
R673 B.n642 B.n9 163.367
R674 B.n642 B.n641 163.367
R675 B.n641 B.n640 163.367
R676 B.n640 B.n11 163.367
R677 B.n636 B.n11 163.367
R678 B.n636 B.n635 163.367
R679 B.n635 B.n634 163.367
R680 B.n634 B.n13 163.367
R681 B.n630 B.n13 163.367
R682 B.n630 B.n629 163.367
R683 B.n629 B.n628 163.367
R684 B.n628 B.n15 163.367
R685 B.n624 B.n15 163.367
R686 B.n624 B.n623 163.367
R687 B.n623 B.n622 163.367
R688 B.n622 B.n17 163.367
R689 B.n618 B.n17 163.367
R690 B.n618 B.n617 163.367
R691 B.n617 B.n616 163.367
R692 B.n616 B.n19 163.367
R693 B.n612 B.n19 163.367
R694 B.n612 B.n611 163.367
R695 B.n611 B.n610 163.367
R696 B.n610 B.n21 163.367
R697 B.n606 B.n21 163.367
R698 B.n606 B.n605 163.367
R699 B.n605 B.n604 163.367
R700 B.n604 B.n23 163.367
R701 B.n600 B.n23 163.367
R702 B.n600 B.n599 163.367
R703 B.n599 B.n598 163.367
R704 B.n598 B.n25 163.367
R705 B.n594 B.n25 163.367
R706 B.n594 B.n593 163.367
R707 B.n593 B.n592 163.367
R708 B.n592 B.n27 163.367
R709 B.n588 B.n27 163.367
R710 B.n588 B.n587 163.367
R711 B.n587 B.n586 163.367
R712 B.n253 B.n252 163.367
R713 B.n253 B.n144 163.367
R714 B.n257 B.n144 163.367
R715 B.n258 B.n257 163.367
R716 B.n259 B.n258 163.367
R717 B.n259 B.n142 163.367
R718 B.n263 B.n142 163.367
R719 B.n264 B.n263 163.367
R720 B.n265 B.n264 163.367
R721 B.n265 B.n140 163.367
R722 B.n269 B.n140 163.367
R723 B.n270 B.n269 163.367
R724 B.n271 B.n270 163.367
R725 B.n271 B.n138 163.367
R726 B.n275 B.n138 163.367
R727 B.n276 B.n275 163.367
R728 B.n277 B.n276 163.367
R729 B.n277 B.n136 163.367
R730 B.n281 B.n136 163.367
R731 B.n282 B.n281 163.367
R732 B.n283 B.n282 163.367
R733 B.n283 B.n132 163.367
R734 B.n288 B.n132 163.367
R735 B.n289 B.n288 163.367
R736 B.n290 B.n289 163.367
R737 B.n290 B.n130 163.367
R738 B.n294 B.n130 163.367
R739 B.n295 B.n294 163.367
R740 B.n296 B.n295 163.367
R741 B.n296 B.n128 163.367
R742 B.n303 B.n128 163.367
R743 B.n304 B.n303 163.367
R744 B.n305 B.n304 163.367
R745 B.n305 B.n126 163.367
R746 B.n309 B.n126 163.367
R747 B.n310 B.n309 163.367
R748 B.n311 B.n310 163.367
R749 B.n311 B.n124 163.367
R750 B.n315 B.n124 163.367
R751 B.n316 B.n315 163.367
R752 B.n317 B.n316 163.367
R753 B.n317 B.n122 163.367
R754 B.n321 B.n122 163.367
R755 B.n322 B.n321 163.367
R756 B.n323 B.n322 163.367
R757 B.n323 B.n120 163.367
R758 B.n327 B.n120 163.367
R759 B.n328 B.n327 163.367
R760 B.n329 B.n328 163.367
R761 B.n329 B.n118 163.367
R762 B.n333 B.n118 163.367
R763 B.n334 B.n333 163.367
R764 B.n335 B.n334 163.367
R765 B.n335 B.n116 163.367
R766 B.n340 B.n339 163.367
R767 B.n341 B.n340 163.367
R768 B.n341 B.n114 163.367
R769 B.n345 B.n114 163.367
R770 B.n346 B.n345 163.367
R771 B.n347 B.n346 163.367
R772 B.n347 B.n112 163.367
R773 B.n351 B.n112 163.367
R774 B.n352 B.n351 163.367
R775 B.n353 B.n352 163.367
R776 B.n353 B.n110 163.367
R777 B.n357 B.n110 163.367
R778 B.n358 B.n357 163.367
R779 B.n359 B.n358 163.367
R780 B.n359 B.n108 163.367
R781 B.n363 B.n108 163.367
R782 B.n364 B.n363 163.367
R783 B.n365 B.n364 163.367
R784 B.n365 B.n106 163.367
R785 B.n369 B.n106 163.367
R786 B.n370 B.n369 163.367
R787 B.n371 B.n370 163.367
R788 B.n371 B.n104 163.367
R789 B.n375 B.n104 163.367
R790 B.n376 B.n375 163.367
R791 B.n377 B.n376 163.367
R792 B.n377 B.n102 163.367
R793 B.n381 B.n102 163.367
R794 B.n382 B.n381 163.367
R795 B.n383 B.n382 163.367
R796 B.n383 B.n100 163.367
R797 B.n387 B.n100 163.367
R798 B.n388 B.n387 163.367
R799 B.n389 B.n388 163.367
R800 B.n389 B.n98 163.367
R801 B.n393 B.n98 163.367
R802 B.n394 B.n393 163.367
R803 B.n395 B.n394 163.367
R804 B.n395 B.n96 163.367
R805 B.n399 B.n96 163.367
R806 B.n400 B.n399 163.367
R807 B.n401 B.n400 163.367
R808 B.n401 B.n94 163.367
R809 B.n405 B.n94 163.367
R810 B.n406 B.n405 163.367
R811 B.n407 B.n406 163.367
R812 B.n407 B.n92 163.367
R813 B.n411 B.n92 163.367
R814 B.n412 B.n411 163.367
R815 B.n413 B.n412 163.367
R816 B.n413 B.n90 163.367
R817 B.n417 B.n90 163.367
R818 B.n418 B.n417 163.367
R819 B.n419 B.n418 163.367
R820 B.n419 B.n88 163.367
R821 B.n423 B.n88 163.367
R822 B.n424 B.n423 163.367
R823 B.n425 B.n424 163.367
R824 B.n425 B.n86 163.367
R825 B.n429 B.n86 163.367
R826 B.n430 B.n429 163.367
R827 B.n431 B.n430 163.367
R828 B.n431 B.n84 163.367
R829 B.n435 B.n84 163.367
R830 B.n436 B.n435 163.367
R831 B.n437 B.n436 163.367
R832 B.n437 B.n82 163.367
R833 B.n441 B.n82 163.367
R834 B.n442 B.n441 163.367
R835 B.n443 B.n442 163.367
R836 B.n443 B.n80 163.367
R837 B.n447 B.n80 163.367
R838 B.n448 B.n447 163.367
R839 B.n449 B.n448 163.367
R840 B.n449 B.n78 163.367
R841 B.n453 B.n78 163.367
R842 B.n454 B.n453 163.367
R843 B.n455 B.n454 163.367
R844 B.n455 B.n76 163.367
R845 B.n459 B.n76 163.367
R846 B.n460 B.n459 163.367
R847 B.n461 B.n460 163.367
R848 B.n461 B.n74 163.367
R849 B.n465 B.n74 163.367
R850 B.n466 B.n465 163.367
R851 B.n467 B.n466 163.367
R852 B.n467 B.n72 163.367
R853 B.n471 B.n72 163.367
R854 B.n472 B.n471 163.367
R855 B.n473 B.n472 163.367
R856 B.n473 B.n70 163.367
R857 B.n477 B.n70 163.367
R858 B.n478 B.n477 163.367
R859 B.n479 B.n478 163.367
R860 B.n479 B.n68 163.367
R861 B.n483 B.n68 163.367
R862 B.n484 B.n483 163.367
R863 B.n485 B.n484 163.367
R864 B.n485 B.n66 163.367
R865 B.n489 B.n66 163.367
R866 B.n490 B.n489 163.367
R867 B.n491 B.n490 163.367
R868 B.n491 B.n64 163.367
R869 B.n495 B.n64 163.367
R870 B.n496 B.n495 163.367
R871 B.n497 B.n496 163.367
R872 B.n497 B.n62 163.367
R873 B.n501 B.n62 163.367
R874 B.n582 B.n29 163.367
R875 B.n582 B.n581 163.367
R876 B.n581 B.n580 163.367
R877 B.n580 B.n31 163.367
R878 B.n576 B.n31 163.367
R879 B.n576 B.n575 163.367
R880 B.n575 B.n574 163.367
R881 B.n574 B.n33 163.367
R882 B.n570 B.n33 163.367
R883 B.n570 B.n569 163.367
R884 B.n569 B.n568 163.367
R885 B.n568 B.n35 163.367
R886 B.n564 B.n35 163.367
R887 B.n564 B.n563 163.367
R888 B.n563 B.n562 163.367
R889 B.n562 B.n37 163.367
R890 B.n558 B.n37 163.367
R891 B.n558 B.n557 163.367
R892 B.n557 B.n556 163.367
R893 B.n556 B.n39 163.367
R894 B.n552 B.n39 163.367
R895 B.n552 B.n551 163.367
R896 B.n551 B.n550 163.367
R897 B.n550 B.n41 163.367
R898 B.n546 B.n41 163.367
R899 B.n546 B.n545 163.367
R900 B.n545 B.n544 163.367
R901 B.n544 B.n46 163.367
R902 B.n540 B.n46 163.367
R903 B.n540 B.n539 163.367
R904 B.n539 B.n538 163.367
R905 B.n538 B.n48 163.367
R906 B.n533 B.n48 163.367
R907 B.n533 B.n532 163.367
R908 B.n532 B.n531 163.367
R909 B.n531 B.n52 163.367
R910 B.n527 B.n52 163.367
R911 B.n527 B.n526 163.367
R912 B.n526 B.n525 163.367
R913 B.n525 B.n54 163.367
R914 B.n521 B.n54 163.367
R915 B.n521 B.n520 163.367
R916 B.n520 B.n519 163.367
R917 B.n519 B.n56 163.367
R918 B.n515 B.n56 163.367
R919 B.n515 B.n514 163.367
R920 B.n514 B.n513 163.367
R921 B.n513 B.n58 163.367
R922 B.n509 B.n58 163.367
R923 B.n509 B.n508 163.367
R924 B.n508 B.n507 163.367
R925 B.n507 B.n60 163.367
R926 B.n503 B.n60 163.367
R927 B.n503 B.n502 163.367
R928 B.n300 B.t10 115.266
R929 B.n50 B.t5 115.266
R930 B.n134 B.t7 115.261
R931 B.n43 B.t2 115.261
R932 B.n300 B.n299 60.5096
R933 B.n134 B.n133 60.5096
R934 B.n43 B.n42 60.5096
R935 B.n50 B.n49 60.5096
R936 B.n301 B.n300 59.5399
R937 B.n286 B.n134 59.5399
R938 B.n44 B.n43 59.5399
R939 B.n536 B.n50 59.5399
R940 B.n585 B.n584 33.2493
R941 B.n500 B.n61 33.2493
R942 B.n338 B.n337 33.2493
R943 B.n250 B.n145 33.2493
R944 B B.n667 18.0485
R945 B.n584 B.n583 10.6151
R946 B.n583 B.n30 10.6151
R947 B.n579 B.n30 10.6151
R948 B.n579 B.n578 10.6151
R949 B.n578 B.n577 10.6151
R950 B.n577 B.n32 10.6151
R951 B.n573 B.n32 10.6151
R952 B.n573 B.n572 10.6151
R953 B.n572 B.n571 10.6151
R954 B.n571 B.n34 10.6151
R955 B.n567 B.n34 10.6151
R956 B.n567 B.n566 10.6151
R957 B.n566 B.n565 10.6151
R958 B.n565 B.n36 10.6151
R959 B.n561 B.n36 10.6151
R960 B.n561 B.n560 10.6151
R961 B.n560 B.n559 10.6151
R962 B.n559 B.n38 10.6151
R963 B.n555 B.n38 10.6151
R964 B.n555 B.n554 10.6151
R965 B.n554 B.n553 10.6151
R966 B.n553 B.n40 10.6151
R967 B.n549 B.n548 10.6151
R968 B.n548 B.n547 10.6151
R969 B.n547 B.n45 10.6151
R970 B.n543 B.n45 10.6151
R971 B.n543 B.n542 10.6151
R972 B.n542 B.n541 10.6151
R973 B.n541 B.n47 10.6151
R974 B.n537 B.n47 10.6151
R975 B.n535 B.n534 10.6151
R976 B.n534 B.n51 10.6151
R977 B.n530 B.n51 10.6151
R978 B.n530 B.n529 10.6151
R979 B.n529 B.n528 10.6151
R980 B.n528 B.n53 10.6151
R981 B.n524 B.n53 10.6151
R982 B.n524 B.n523 10.6151
R983 B.n523 B.n522 10.6151
R984 B.n522 B.n55 10.6151
R985 B.n518 B.n55 10.6151
R986 B.n518 B.n517 10.6151
R987 B.n517 B.n516 10.6151
R988 B.n516 B.n57 10.6151
R989 B.n512 B.n57 10.6151
R990 B.n512 B.n511 10.6151
R991 B.n511 B.n510 10.6151
R992 B.n510 B.n59 10.6151
R993 B.n506 B.n59 10.6151
R994 B.n506 B.n505 10.6151
R995 B.n505 B.n504 10.6151
R996 B.n504 B.n61 10.6151
R997 B.n338 B.n115 10.6151
R998 B.n342 B.n115 10.6151
R999 B.n343 B.n342 10.6151
R1000 B.n344 B.n343 10.6151
R1001 B.n344 B.n113 10.6151
R1002 B.n348 B.n113 10.6151
R1003 B.n349 B.n348 10.6151
R1004 B.n350 B.n349 10.6151
R1005 B.n350 B.n111 10.6151
R1006 B.n354 B.n111 10.6151
R1007 B.n355 B.n354 10.6151
R1008 B.n356 B.n355 10.6151
R1009 B.n356 B.n109 10.6151
R1010 B.n360 B.n109 10.6151
R1011 B.n361 B.n360 10.6151
R1012 B.n362 B.n361 10.6151
R1013 B.n362 B.n107 10.6151
R1014 B.n366 B.n107 10.6151
R1015 B.n367 B.n366 10.6151
R1016 B.n368 B.n367 10.6151
R1017 B.n368 B.n105 10.6151
R1018 B.n372 B.n105 10.6151
R1019 B.n373 B.n372 10.6151
R1020 B.n374 B.n373 10.6151
R1021 B.n374 B.n103 10.6151
R1022 B.n378 B.n103 10.6151
R1023 B.n379 B.n378 10.6151
R1024 B.n380 B.n379 10.6151
R1025 B.n380 B.n101 10.6151
R1026 B.n384 B.n101 10.6151
R1027 B.n385 B.n384 10.6151
R1028 B.n386 B.n385 10.6151
R1029 B.n386 B.n99 10.6151
R1030 B.n390 B.n99 10.6151
R1031 B.n391 B.n390 10.6151
R1032 B.n392 B.n391 10.6151
R1033 B.n392 B.n97 10.6151
R1034 B.n396 B.n97 10.6151
R1035 B.n397 B.n396 10.6151
R1036 B.n398 B.n397 10.6151
R1037 B.n398 B.n95 10.6151
R1038 B.n402 B.n95 10.6151
R1039 B.n403 B.n402 10.6151
R1040 B.n404 B.n403 10.6151
R1041 B.n404 B.n93 10.6151
R1042 B.n408 B.n93 10.6151
R1043 B.n409 B.n408 10.6151
R1044 B.n410 B.n409 10.6151
R1045 B.n410 B.n91 10.6151
R1046 B.n414 B.n91 10.6151
R1047 B.n415 B.n414 10.6151
R1048 B.n416 B.n415 10.6151
R1049 B.n416 B.n89 10.6151
R1050 B.n420 B.n89 10.6151
R1051 B.n421 B.n420 10.6151
R1052 B.n422 B.n421 10.6151
R1053 B.n422 B.n87 10.6151
R1054 B.n426 B.n87 10.6151
R1055 B.n427 B.n426 10.6151
R1056 B.n428 B.n427 10.6151
R1057 B.n428 B.n85 10.6151
R1058 B.n432 B.n85 10.6151
R1059 B.n433 B.n432 10.6151
R1060 B.n434 B.n433 10.6151
R1061 B.n434 B.n83 10.6151
R1062 B.n438 B.n83 10.6151
R1063 B.n439 B.n438 10.6151
R1064 B.n440 B.n439 10.6151
R1065 B.n440 B.n81 10.6151
R1066 B.n444 B.n81 10.6151
R1067 B.n445 B.n444 10.6151
R1068 B.n446 B.n445 10.6151
R1069 B.n446 B.n79 10.6151
R1070 B.n450 B.n79 10.6151
R1071 B.n451 B.n450 10.6151
R1072 B.n452 B.n451 10.6151
R1073 B.n452 B.n77 10.6151
R1074 B.n456 B.n77 10.6151
R1075 B.n457 B.n456 10.6151
R1076 B.n458 B.n457 10.6151
R1077 B.n458 B.n75 10.6151
R1078 B.n462 B.n75 10.6151
R1079 B.n463 B.n462 10.6151
R1080 B.n464 B.n463 10.6151
R1081 B.n464 B.n73 10.6151
R1082 B.n468 B.n73 10.6151
R1083 B.n469 B.n468 10.6151
R1084 B.n470 B.n469 10.6151
R1085 B.n470 B.n71 10.6151
R1086 B.n474 B.n71 10.6151
R1087 B.n475 B.n474 10.6151
R1088 B.n476 B.n475 10.6151
R1089 B.n476 B.n69 10.6151
R1090 B.n480 B.n69 10.6151
R1091 B.n481 B.n480 10.6151
R1092 B.n482 B.n481 10.6151
R1093 B.n482 B.n67 10.6151
R1094 B.n486 B.n67 10.6151
R1095 B.n487 B.n486 10.6151
R1096 B.n488 B.n487 10.6151
R1097 B.n488 B.n65 10.6151
R1098 B.n492 B.n65 10.6151
R1099 B.n493 B.n492 10.6151
R1100 B.n494 B.n493 10.6151
R1101 B.n494 B.n63 10.6151
R1102 B.n498 B.n63 10.6151
R1103 B.n499 B.n498 10.6151
R1104 B.n500 B.n499 10.6151
R1105 B.n254 B.n145 10.6151
R1106 B.n255 B.n254 10.6151
R1107 B.n256 B.n255 10.6151
R1108 B.n256 B.n143 10.6151
R1109 B.n260 B.n143 10.6151
R1110 B.n261 B.n260 10.6151
R1111 B.n262 B.n261 10.6151
R1112 B.n262 B.n141 10.6151
R1113 B.n266 B.n141 10.6151
R1114 B.n267 B.n266 10.6151
R1115 B.n268 B.n267 10.6151
R1116 B.n268 B.n139 10.6151
R1117 B.n272 B.n139 10.6151
R1118 B.n273 B.n272 10.6151
R1119 B.n274 B.n273 10.6151
R1120 B.n274 B.n137 10.6151
R1121 B.n278 B.n137 10.6151
R1122 B.n279 B.n278 10.6151
R1123 B.n280 B.n279 10.6151
R1124 B.n280 B.n135 10.6151
R1125 B.n284 B.n135 10.6151
R1126 B.n285 B.n284 10.6151
R1127 B.n287 B.n131 10.6151
R1128 B.n291 B.n131 10.6151
R1129 B.n292 B.n291 10.6151
R1130 B.n293 B.n292 10.6151
R1131 B.n293 B.n129 10.6151
R1132 B.n297 B.n129 10.6151
R1133 B.n298 B.n297 10.6151
R1134 B.n302 B.n298 10.6151
R1135 B.n306 B.n127 10.6151
R1136 B.n307 B.n306 10.6151
R1137 B.n308 B.n307 10.6151
R1138 B.n308 B.n125 10.6151
R1139 B.n312 B.n125 10.6151
R1140 B.n313 B.n312 10.6151
R1141 B.n314 B.n313 10.6151
R1142 B.n314 B.n123 10.6151
R1143 B.n318 B.n123 10.6151
R1144 B.n319 B.n318 10.6151
R1145 B.n320 B.n319 10.6151
R1146 B.n320 B.n121 10.6151
R1147 B.n324 B.n121 10.6151
R1148 B.n325 B.n324 10.6151
R1149 B.n326 B.n325 10.6151
R1150 B.n326 B.n119 10.6151
R1151 B.n330 B.n119 10.6151
R1152 B.n331 B.n330 10.6151
R1153 B.n332 B.n331 10.6151
R1154 B.n332 B.n117 10.6151
R1155 B.n336 B.n117 10.6151
R1156 B.n337 B.n336 10.6151
R1157 B.n250 B.n249 10.6151
R1158 B.n249 B.n248 10.6151
R1159 B.n248 B.n147 10.6151
R1160 B.n244 B.n147 10.6151
R1161 B.n244 B.n243 10.6151
R1162 B.n243 B.n242 10.6151
R1163 B.n242 B.n149 10.6151
R1164 B.n238 B.n149 10.6151
R1165 B.n238 B.n237 10.6151
R1166 B.n237 B.n236 10.6151
R1167 B.n236 B.n151 10.6151
R1168 B.n232 B.n151 10.6151
R1169 B.n232 B.n231 10.6151
R1170 B.n231 B.n230 10.6151
R1171 B.n230 B.n153 10.6151
R1172 B.n226 B.n153 10.6151
R1173 B.n226 B.n225 10.6151
R1174 B.n225 B.n224 10.6151
R1175 B.n224 B.n155 10.6151
R1176 B.n220 B.n155 10.6151
R1177 B.n220 B.n219 10.6151
R1178 B.n219 B.n218 10.6151
R1179 B.n218 B.n157 10.6151
R1180 B.n214 B.n157 10.6151
R1181 B.n214 B.n213 10.6151
R1182 B.n213 B.n212 10.6151
R1183 B.n212 B.n159 10.6151
R1184 B.n208 B.n159 10.6151
R1185 B.n208 B.n207 10.6151
R1186 B.n207 B.n206 10.6151
R1187 B.n206 B.n161 10.6151
R1188 B.n202 B.n161 10.6151
R1189 B.n202 B.n201 10.6151
R1190 B.n201 B.n200 10.6151
R1191 B.n200 B.n163 10.6151
R1192 B.n196 B.n163 10.6151
R1193 B.n196 B.n195 10.6151
R1194 B.n195 B.n194 10.6151
R1195 B.n194 B.n165 10.6151
R1196 B.n190 B.n165 10.6151
R1197 B.n190 B.n189 10.6151
R1198 B.n189 B.n188 10.6151
R1199 B.n188 B.n167 10.6151
R1200 B.n184 B.n167 10.6151
R1201 B.n184 B.n183 10.6151
R1202 B.n183 B.n182 10.6151
R1203 B.n182 B.n169 10.6151
R1204 B.n178 B.n169 10.6151
R1205 B.n178 B.n177 10.6151
R1206 B.n177 B.n176 10.6151
R1207 B.n176 B.n171 10.6151
R1208 B.n172 B.n171 10.6151
R1209 B.n172 B.n0 10.6151
R1210 B.n663 B.n1 10.6151
R1211 B.n663 B.n662 10.6151
R1212 B.n662 B.n661 10.6151
R1213 B.n661 B.n4 10.6151
R1214 B.n657 B.n4 10.6151
R1215 B.n657 B.n656 10.6151
R1216 B.n656 B.n655 10.6151
R1217 B.n655 B.n6 10.6151
R1218 B.n651 B.n6 10.6151
R1219 B.n651 B.n650 10.6151
R1220 B.n650 B.n649 10.6151
R1221 B.n649 B.n8 10.6151
R1222 B.n645 B.n8 10.6151
R1223 B.n645 B.n644 10.6151
R1224 B.n644 B.n643 10.6151
R1225 B.n643 B.n10 10.6151
R1226 B.n639 B.n10 10.6151
R1227 B.n639 B.n638 10.6151
R1228 B.n638 B.n637 10.6151
R1229 B.n637 B.n12 10.6151
R1230 B.n633 B.n12 10.6151
R1231 B.n633 B.n632 10.6151
R1232 B.n632 B.n631 10.6151
R1233 B.n631 B.n14 10.6151
R1234 B.n627 B.n14 10.6151
R1235 B.n627 B.n626 10.6151
R1236 B.n626 B.n625 10.6151
R1237 B.n625 B.n16 10.6151
R1238 B.n621 B.n16 10.6151
R1239 B.n621 B.n620 10.6151
R1240 B.n620 B.n619 10.6151
R1241 B.n619 B.n18 10.6151
R1242 B.n615 B.n18 10.6151
R1243 B.n615 B.n614 10.6151
R1244 B.n614 B.n613 10.6151
R1245 B.n613 B.n20 10.6151
R1246 B.n609 B.n20 10.6151
R1247 B.n609 B.n608 10.6151
R1248 B.n608 B.n607 10.6151
R1249 B.n607 B.n22 10.6151
R1250 B.n603 B.n22 10.6151
R1251 B.n603 B.n602 10.6151
R1252 B.n602 B.n601 10.6151
R1253 B.n601 B.n24 10.6151
R1254 B.n597 B.n24 10.6151
R1255 B.n597 B.n596 10.6151
R1256 B.n596 B.n595 10.6151
R1257 B.n595 B.n26 10.6151
R1258 B.n591 B.n26 10.6151
R1259 B.n591 B.n590 10.6151
R1260 B.n590 B.n589 10.6151
R1261 B.n589 B.n28 10.6151
R1262 B.n585 B.n28 10.6151
R1263 B.n549 B.n44 6.5566
R1264 B.n537 B.n536 6.5566
R1265 B.n287 B.n286 6.5566
R1266 B.n302 B.n301 6.5566
R1267 B.n44 B.n40 4.05904
R1268 B.n536 B.n535 4.05904
R1269 B.n286 B.n285 4.05904
R1270 B.n301 B.n127 4.05904
R1271 B.n667 B.n0 2.81026
R1272 B.n667 B.n1 2.81026
C0 VP VDD1 4.74186f
C1 VN VDD2 4.35554f
C2 VP VN 6.70839f
C3 VP VDD2 0.540193f
C4 w_n4090_n2088# VTAIL 2.79326f
C5 w_n4090_n2088# B 8.62639f
C6 VTAIL B 2.9304f
C7 w_n4090_n2088# VDD1 1.84436f
C8 VTAIL VDD1 6.05044f
C9 VDD1 B 1.5342f
C10 w_n4090_n2088# VN 8.26575f
C11 VN VTAIL 5.28966f
C12 w_n4090_n2088# VDD2 1.96689f
C13 VN B 1.19141f
C14 VTAIL VDD2 6.10613f
C15 VDD2 B 1.63637f
C16 w_n4090_n2088# VP 8.79728f
C17 VN VDD1 0.152375f
C18 VP VTAIL 5.30377f
C19 VP B 2.08344f
C20 VDD2 VDD1 1.87613f
C21 VDD2 VSUBS 1.614149f
C22 VDD1 VSUBS 2.304857f
C23 VTAIL VSUBS 0.709813f
C24 VN VSUBS 6.77079f
C25 VP VSUBS 3.368962f
C26 B VSUBS 4.53397f
C27 w_n4090_n2088# VSUBS 0.106749p
C28 B.n0 VSUBS 0.006087f
C29 B.n1 VSUBS 0.006087f
C30 B.n2 VSUBS 0.009626f
C31 B.n3 VSUBS 0.009626f
C32 B.n4 VSUBS 0.009626f
C33 B.n5 VSUBS 0.009626f
C34 B.n6 VSUBS 0.009626f
C35 B.n7 VSUBS 0.009626f
C36 B.n8 VSUBS 0.009626f
C37 B.n9 VSUBS 0.009626f
C38 B.n10 VSUBS 0.009626f
C39 B.n11 VSUBS 0.009626f
C40 B.n12 VSUBS 0.009626f
C41 B.n13 VSUBS 0.009626f
C42 B.n14 VSUBS 0.009626f
C43 B.n15 VSUBS 0.009626f
C44 B.n16 VSUBS 0.009626f
C45 B.n17 VSUBS 0.009626f
C46 B.n18 VSUBS 0.009626f
C47 B.n19 VSUBS 0.009626f
C48 B.n20 VSUBS 0.009626f
C49 B.n21 VSUBS 0.009626f
C50 B.n22 VSUBS 0.009626f
C51 B.n23 VSUBS 0.009626f
C52 B.n24 VSUBS 0.009626f
C53 B.n25 VSUBS 0.009626f
C54 B.n26 VSUBS 0.009626f
C55 B.n27 VSUBS 0.009626f
C56 B.n28 VSUBS 0.009626f
C57 B.n29 VSUBS 0.02324f
C58 B.n30 VSUBS 0.009626f
C59 B.n31 VSUBS 0.009626f
C60 B.n32 VSUBS 0.009626f
C61 B.n33 VSUBS 0.009626f
C62 B.n34 VSUBS 0.009626f
C63 B.n35 VSUBS 0.009626f
C64 B.n36 VSUBS 0.009626f
C65 B.n37 VSUBS 0.009626f
C66 B.n38 VSUBS 0.009626f
C67 B.n39 VSUBS 0.009626f
C68 B.n40 VSUBS 0.006653f
C69 B.n41 VSUBS 0.009626f
C70 B.t2 VSUBS 0.221186f
C71 B.t1 VSUBS 0.25026f
C72 B.t0 VSUBS 1.02266f
C73 B.n42 VSUBS 0.154634f
C74 B.n43 VSUBS 0.098186f
C75 B.n44 VSUBS 0.022302f
C76 B.n45 VSUBS 0.009626f
C77 B.n46 VSUBS 0.009626f
C78 B.n47 VSUBS 0.009626f
C79 B.n48 VSUBS 0.009626f
C80 B.t5 VSUBS 0.221186f
C81 B.t4 VSUBS 0.250259f
C82 B.t3 VSUBS 1.02266f
C83 B.n49 VSUBS 0.154635f
C84 B.n50 VSUBS 0.098186f
C85 B.n51 VSUBS 0.009626f
C86 B.n52 VSUBS 0.009626f
C87 B.n53 VSUBS 0.009626f
C88 B.n54 VSUBS 0.009626f
C89 B.n55 VSUBS 0.009626f
C90 B.n56 VSUBS 0.009626f
C91 B.n57 VSUBS 0.009626f
C92 B.n58 VSUBS 0.009626f
C93 B.n59 VSUBS 0.009626f
C94 B.n60 VSUBS 0.009626f
C95 B.n61 VSUBS 0.022123f
C96 B.n62 VSUBS 0.009626f
C97 B.n63 VSUBS 0.009626f
C98 B.n64 VSUBS 0.009626f
C99 B.n65 VSUBS 0.009626f
C100 B.n66 VSUBS 0.009626f
C101 B.n67 VSUBS 0.009626f
C102 B.n68 VSUBS 0.009626f
C103 B.n69 VSUBS 0.009626f
C104 B.n70 VSUBS 0.009626f
C105 B.n71 VSUBS 0.009626f
C106 B.n72 VSUBS 0.009626f
C107 B.n73 VSUBS 0.009626f
C108 B.n74 VSUBS 0.009626f
C109 B.n75 VSUBS 0.009626f
C110 B.n76 VSUBS 0.009626f
C111 B.n77 VSUBS 0.009626f
C112 B.n78 VSUBS 0.009626f
C113 B.n79 VSUBS 0.009626f
C114 B.n80 VSUBS 0.009626f
C115 B.n81 VSUBS 0.009626f
C116 B.n82 VSUBS 0.009626f
C117 B.n83 VSUBS 0.009626f
C118 B.n84 VSUBS 0.009626f
C119 B.n85 VSUBS 0.009626f
C120 B.n86 VSUBS 0.009626f
C121 B.n87 VSUBS 0.009626f
C122 B.n88 VSUBS 0.009626f
C123 B.n89 VSUBS 0.009626f
C124 B.n90 VSUBS 0.009626f
C125 B.n91 VSUBS 0.009626f
C126 B.n92 VSUBS 0.009626f
C127 B.n93 VSUBS 0.009626f
C128 B.n94 VSUBS 0.009626f
C129 B.n95 VSUBS 0.009626f
C130 B.n96 VSUBS 0.009626f
C131 B.n97 VSUBS 0.009626f
C132 B.n98 VSUBS 0.009626f
C133 B.n99 VSUBS 0.009626f
C134 B.n100 VSUBS 0.009626f
C135 B.n101 VSUBS 0.009626f
C136 B.n102 VSUBS 0.009626f
C137 B.n103 VSUBS 0.009626f
C138 B.n104 VSUBS 0.009626f
C139 B.n105 VSUBS 0.009626f
C140 B.n106 VSUBS 0.009626f
C141 B.n107 VSUBS 0.009626f
C142 B.n108 VSUBS 0.009626f
C143 B.n109 VSUBS 0.009626f
C144 B.n110 VSUBS 0.009626f
C145 B.n111 VSUBS 0.009626f
C146 B.n112 VSUBS 0.009626f
C147 B.n113 VSUBS 0.009626f
C148 B.n114 VSUBS 0.009626f
C149 B.n115 VSUBS 0.009626f
C150 B.n116 VSUBS 0.02324f
C151 B.n117 VSUBS 0.009626f
C152 B.n118 VSUBS 0.009626f
C153 B.n119 VSUBS 0.009626f
C154 B.n120 VSUBS 0.009626f
C155 B.n121 VSUBS 0.009626f
C156 B.n122 VSUBS 0.009626f
C157 B.n123 VSUBS 0.009626f
C158 B.n124 VSUBS 0.009626f
C159 B.n125 VSUBS 0.009626f
C160 B.n126 VSUBS 0.009626f
C161 B.n127 VSUBS 0.006653f
C162 B.n128 VSUBS 0.009626f
C163 B.n129 VSUBS 0.009626f
C164 B.n130 VSUBS 0.009626f
C165 B.n131 VSUBS 0.009626f
C166 B.n132 VSUBS 0.009626f
C167 B.t7 VSUBS 0.221186f
C168 B.t8 VSUBS 0.25026f
C169 B.t6 VSUBS 1.02266f
C170 B.n133 VSUBS 0.154634f
C171 B.n134 VSUBS 0.098186f
C172 B.n135 VSUBS 0.009626f
C173 B.n136 VSUBS 0.009626f
C174 B.n137 VSUBS 0.009626f
C175 B.n138 VSUBS 0.009626f
C176 B.n139 VSUBS 0.009626f
C177 B.n140 VSUBS 0.009626f
C178 B.n141 VSUBS 0.009626f
C179 B.n142 VSUBS 0.009626f
C180 B.n143 VSUBS 0.009626f
C181 B.n144 VSUBS 0.009626f
C182 B.n145 VSUBS 0.02324f
C183 B.n146 VSUBS 0.009626f
C184 B.n147 VSUBS 0.009626f
C185 B.n148 VSUBS 0.009626f
C186 B.n149 VSUBS 0.009626f
C187 B.n150 VSUBS 0.009626f
C188 B.n151 VSUBS 0.009626f
C189 B.n152 VSUBS 0.009626f
C190 B.n153 VSUBS 0.009626f
C191 B.n154 VSUBS 0.009626f
C192 B.n155 VSUBS 0.009626f
C193 B.n156 VSUBS 0.009626f
C194 B.n157 VSUBS 0.009626f
C195 B.n158 VSUBS 0.009626f
C196 B.n159 VSUBS 0.009626f
C197 B.n160 VSUBS 0.009626f
C198 B.n161 VSUBS 0.009626f
C199 B.n162 VSUBS 0.009626f
C200 B.n163 VSUBS 0.009626f
C201 B.n164 VSUBS 0.009626f
C202 B.n165 VSUBS 0.009626f
C203 B.n166 VSUBS 0.009626f
C204 B.n167 VSUBS 0.009626f
C205 B.n168 VSUBS 0.009626f
C206 B.n169 VSUBS 0.009626f
C207 B.n170 VSUBS 0.009626f
C208 B.n171 VSUBS 0.009626f
C209 B.n172 VSUBS 0.009626f
C210 B.n173 VSUBS 0.009626f
C211 B.n174 VSUBS 0.009626f
C212 B.n175 VSUBS 0.009626f
C213 B.n176 VSUBS 0.009626f
C214 B.n177 VSUBS 0.009626f
C215 B.n178 VSUBS 0.009626f
C216 B.n179 VSUBS 0.009626f
C217 B.n180 VSUBS 0.009626f
C218 B.n181 VSUBS 0.009626f
C219 B.n182 VSUBS 0.009626f
C220 B.n183 VSUBS 0.009626f
C221 B.n184 VSUBS 0.009626f
C222 B.n185 VSUBS 0.009626f
C223 B.n186 VSUBS 0.009626f
C224 B.n187 VSUBS 0.009626f
C225 B.n188 VSUBS 0.009626f
C226 B.n189 VSUBS 0.009626f
C227 B.n190 VSUBS 0.009626f
C228 B.n191 VSUBS 0.009626f
C229 B.n192 VSUBS 0.009626f
C230 B.n193 VSUBS 0.009626f
C231 B.n194 VSUBS 0.009626f
C232 B.n195 VSUBS 0.009626f
C233 B.n196 VSUBS 0.009626f
C234 B.n197 VSUBS 0.009626f
C235 B.n198 VSUBS 0.009626f
C236 B.n199 VSUBS 0.009626f
C237 B.n200 VSUBS 0.009626f
C238 B.n201 VSUBS 0.009626f
C239 B.n202 VSUBS 0.009626f
C240 B.n203 VSUBS 0.009626f
C241 B.n204 VSUBS 0.009626f
C242 B.n205 VSUBS 0.009626f
C243 B.n206 VSUBS 0.009626f
C244 B.n207 VSUBS 0.009626f
C245 B.n208 VSUBS 0.009626f
C246 B.n209 VSUBS 0.009626f
C247 B.n210 VSUBS 0.009626f
C248 B.n211 VSUBS 0.009626f
C249 B.n212 VSUBS 0.009626f
C250 B.n213 VSUBS 0.009626f
C251 B.n214 VSUBS 0.009626f
C252 B.n215 VSUBS 0.009626f
C253 B.n216 VSUBS 0.009626f
C254 B.n217 VSUBS 0.009626f
C255 B.n218 VSUBS 0.009626f
C256 B.n219 VSUBS 0.009626f
C257 B.n220 VSUBS 0.009626f
C258 B.n221 VSUBS 0.009626f
C259 B.n222 VSUBS 0.009626f
C260 B.n223 VSUBS 0.009626f
C261 B.n224 VSUBS 0.009626f
C262 B.n225 VSUBS 0.009626f
C263 B.n226 VSUBS 0.009626f
C264 B.n227 VSUBS 0.009626f
C265 B.n228 VSUBS 0.009626f
C266 B.n229 VSUBS 0.009626f
C267 B.n230 VSUBS 0.009626f
C268 B.n231 VSUBS 0.009626f
C269 B.n232 VSUBS 0.009626f
C270 B.n233 VSUBS 0.009626f
C271 B.n234 VSUBS 0.009626f
C272 B.n235 VSUBS 0.009626f
C273 B.n236 VSUBS 0.009626f
C274 B.n237 VSUBS 0.009626f
C275 B.n238 VSUBS 0.009626f
C276 B.n239 VSUBS 0.009626f
C277 B.n240 VSUBS 0.009626f
C278 B.n241 VSUBS 0.009626f
C279 B.n242 VSUBS 0.009626f
C280 B.n243 VSUBS 0.009626f
C281 B.n244 VSUBS 0.009626f
C282 B.n245 VSUBS 0.009626f
C283 B.n246 VSUBS 0.009626f
C284 B.n247 VSUBS 0.009626f
C285 B.n248 VSUBS 0.009626f
C286 B.n249 VSUBS 0.009626f
C287 B.n250 VSUBS 0.022341f
C288 B.n251 VSUBS 0.022341f
C289 B.n252 VSUBS 0.02324f
C290 B.n253 VSUBS 0.009626f
C291 B.n254 VSUBS 0.009626f
C292 B.n255 VSUBS 0.009626f
C293 B.n256 VSUBS 0.009626f
C294 B.n257 VSUBS 0.009626f
C295 B.n258 VSUBS 0.009626f
C296 B.n259 VSUBS 0.009626f
C297 B.n260 VSUBS 0.009626f
C298 B.n261 VSUBS 0.009626f
C299 B.n262 VSUBS 0.009626f
C300 B.n263 VSUBS 0.009626f
C301 B.n264 VSUBS 0.009626f
C302 B.n265 VSUBS 0.009626f
C303 B.n266 VSUBS 0.009626f
C304 B.n267 VSUBS 0.009626f
C305 B.n268 VSUBS 0.009626f
C306 B.n269 VSUBS 0.009626f
C307 B.n270 VSUBS 0.009626f
C308 B.n271 VSUBS 0.009626f
C309 B.n272 VSUBS 0.009626f
C310 B.n273 VSUBS 0.009626f
C311 B.n274 VSUBS 0.009626f
C312 B.n275 VSUBS 0.009626f
C313 B.n276 VSUBS 0.009626f
C314 B.n277 VSUBS 0.009626f
C315 B.n278 VSUBS 0.009626f
C316 B.n279 VSUBS 0.009626f
C317 B.n280 VSUBS 0.009626f
C318 B.n281 VSUBS 0.009626f
C319 B.n282 VSUBS 0.009626f
C320 B.n283 VSUBS 0.009626f
C321 B.n284 VSUBS 0.009626f
C322 B.n285 VSUBS 0.006653f
C323 B.n286 VSUBS 0.022302f
C324 B.n287 VSUBS 0.007785f
C325 B.n288 VSUBS 0.009626f
C326 B.n289 VSUBS 0.009626f
C327 B.n290 VSUBS 0.009626f
C328 B.n291 VSUBS 0.009626f
C329 B.n292 VSUBS 0.009626f
C330 B.n293 VSUBS 0.009626f
C331 B.n294 VSUBS 0.009626f
C332 B.n295 VSUBS 0.009626f
C333 B.n296 VSUBS 0.009626f
C334 B.n297 VSUBS 0.009626f
C335 B.n298 VSUBS 0.009626f
C336 B.t10 VSUBS 0.221186f
C337 B.t11 VSUBS 0.250259f
C338 B.t9 VSUBS 1.02266f
C339 B.n299 VSUBS 0.154635f
C340 B.n300 VSUBS 0.098186f
C341 B.n301 VSUBS 0.022302f
C342 B.n302 VSUBS 0.007785f
C343 B.n303 VSUBS 0.009626f
C344 B.n304 VSUBS 0.009626f
C345 B.n305 VSUBS 0.009626f
C346 B.n306 VSUBS 0.009626f
C347 B.n307 VSUBS 0.009626f
C348 B.n308 VSUBS 0.009626f
C349 B.n309 VSUBS 0.009626f
C350 B.n310 VSUBS 0.009626f
C351 B.n311 VSUBS 0.009626f
C352 B.n312 VSUBS 0.009626f
C353 B.n313 VSUBS 0.009626f
C354 B.n314 VSUBS 0.009626f
C355 B.n315 VSUBS 0.009626f
C356 B.n316 VSUBS 0.009626f
C357 B.n317 VSUBS 0.009626f
C358 B.n318 VSUBS 0.009626f
C359 B.n319 VSUBS 0.009626f
C360 B.n320 VSUBS 0.009626f
C361 B.n321 VSUBS 0.009626f
C362 B.n322 VSUBS 0.009626f
C363 B.n323 VSUBS 0.009626f
C364 B.n324 VSUBS 0.009626f
C365 B.n325 VSUBS 0.009626f
C366 B.n326 VSUBS 0.009626f
C367 B.n327 VSUBS 0.009626f
C368 B.n328 VSUBS 0.009626f
C369 B.n329 VSUBS 0.009626f
C370 B.n330 VSUBS 0.009626f
C371 B.n331 VSUBS 0.009626f
C372 B.n332 VSUBS 0.009626f
C373 B.n333 VSUBS 0.009626f
C374 B.n334 VSUBS 0.009626f
C375 B.n335 VSUBS 0.009626f
C376 B.n336 VSUBS 0.009626f
C377 B.n337 VSUBS 0.02324f
C378 B.n338 VSUBS 0.022341f
C379 B.n339 VSUBS 0.022341f
C380 B.n340 VSUBS 0.009626f
C381 B.n341 VSUBS 0.009626f
C382 B.n342 VSUBS 0.009626f
C383 B.n343 VSUBS 0.009626f
C384 B.n344 VSUBS 0.009626f
C385 B.n345 VSUBS 0.009626f
C386 B.n346 VSUBS 0.009626f
C387 B.n347 VSUBS 0.009626f
C388 B.n348 VSUBS 0.009626f
C389 B.n349 VSUBS 0.009626f
C390 B.n350 VSUBS 0.009626f
C391 B.n351 VSUBS 0.009626f
C392 B.n352 VSUBS 0.009626f
C393 B.n353 VSUBS 0.009626f
C394 B.n354 VSUBS 0.009626f
C395 B.n355 VSUBS 0.009626f
C396 B.n356 VSUBS 0.009626f
C397 B.n357 VSUBS 0.009626f
C398 B.n358 VSUBS 0.009626f
C399 B.n359 VSUBS 0.009626f
C400 B.n360 VSUBS 0.009626f
C401 B.n361 VSUBS 0.009626f
C402 B.n362 VSUBS 0.009626f
C403 B.n363 VSUBS 0.009626f
C404 B.n364 VSUBS 0.009626f
C405 B.n365 VSUBS 0.009626f
C406 B.n366 VSUBS 0.009626f
C407 B.n367 VSUBS 0.009626f
C408 B.n368 VSUBS 0.009626f
C409 B.n369 VSUBS 0.009626f
C410 B.n370 VSUBS 0.009626f
C411 B.n371 VSUBS 0.009626f
C412 B.n372 VSUBS 0.009626f
C413 B.n373 VSUBS 0.009626f
C414 B.n374 VSUBS 0.009626f
C415 B.n375 VSUBS 0.009626f
C416 B.n376 VSUBS 0.009626f
C417 B.n377 VSUBS 0.009626f
C418 B.n378 VSUBS 0.009626f
C419 B.n379 VSUBS 0.009626f
C420 B.n380 VSUBS 0.009626f
C421 B.n381 VSUBS 0.009626f
C422 B.n382 VSUBS 0.009626f
C423 B.n383 VSUBS 0.009626f
C424 B.n384 VSUBS 0.009626f
C425 B.n385 VSUBS 0.009626f
C426 B.n386 VSUBS 0.009626f
C427 B.n387 VSUBS 0.009626f
C428 B.n388 VSUBS 0.009626f
C429 B.n389 VSUBS 0.009626f
C430 B.n390 VSUBS 0.009626f
C431 B.n391 VSUBS 0.009626f
C432 B.n392 VSUBS 0.009626f
C433 B.n393 VSUBS 0.009626f
C434 B.n394 VSUBS 0.009626f
C435 B.n395 VSUBS 0.009626f
C436 B.n396 VSUBS 0.009626f
C437 B.n397 VSUBS 0.009626f
C438 B.n398 VSUBS 0.009626f
C439 B.n399 VSUBS 0.009626f
C440 B.n400 VSUBS 0.009626f
C441 B.n401 VSUBS 0.009626f
C442 B.n402 VSUBS 0.009626f
C443 B.n403 VSUBS 0.009626f
C444 B.n404 VSUBS 0.009626f
C445 B.n405 VSUBS 0.009626f
C446 B.n406 VSUBS 0.009626f
C447 B.n407 VSUBS 0.009626f
C448 B.n408 VSUBS 0.009626f
C449 B.n409 VSUBS 0.009626f
C450 B.n410 VSUBS 0.009626f
C451 B.n411 VSUBS 0.009626f
C452 B.n412 VSUBS 0.009626f
C453 B.n413 VSUBS 0.009626f
C454 B.n414 VSUBS 0.009626f
C455 B.n415 VSUBS 0.009626f
C456 B.n416 VSUBS 0.009626f
C457 B.n417 VSUBS 0.009626f
C458 B.n418 VSUBS 0.009626f
C459 B.n419 VSUBS 0.009626f
C460 B.n420 VSUBS 0.009626f
C461 B.n421 VSUBS 0.009626f
C462 B.n422 VSUBS 0.009626f
C463 B.n423 VSUBS 0.009626f
C464 B.n424 VSUBS 0.009626f
C465 B.n425 VSUBS 0.009626f
C466 B.n426 VSUBS 0.009626f
C467 B.n427 VSUBS 0.009626f
C468 B.n428 VSUBS 0.009626f
C469 B.n429 VSUBS 0.009626f
C470 B.n430 VSUBS 0.009626f
C471 B.n431 VSUBS 0.009626f
C472 B.n432 VSUBS 0.009626f
C473 B.n433 VSUBS 0.009626f
C474 B.n434 VSUBS 0.009626f
C475 B.n435 VSUBS 0.009626f
C476 B.n436 VSUBS 0.009626f
C477 B.n437 VSUBS 0.009626f
C478 B.n438 VSUBS 0.009626f
C479 B.n439 VSUBS 0.009626f
C480 B.n440 VSUBS 0.009626f
C481 B.n441 VSUBS 0.009626f
C482 B.n442 VSUBS 0.009626f
C483 B.n443 VSUBS 0.009626f
C484 B.n444 VSUBS 0.009626f
C485 B.n445 VSUBS 0.009626f
C486 B.n446 VSUBS 0.009626f
C487 B.n447 VSUBS 0.009626f
C488 B.n448 VSUBS 0.009626f
C489 B.n449 VSUBS 0.009626f
C490 B.n450 VSUBS 0.009626f
C491 B.n451 VSUBS 0.009626f
C492 B.n452 VSUBS 0.009626f
C493 B.n453 VSUBS 0.009626f
C494 B.n454 VSUBS 0.009626f
C495 B.n455 VSUBS 0.009626f
C496 B.n456 VSUBS 0.009626f
C497 B.n457 VSUBS 0.009626f
C498 B.n458 VSUBS 0.009626f
C499 B.n459 VSUBS 0.009626f
C500 B.n460 VSUBS 0.009626f
C501 B.n461 VSUBS 0.009626f
C502 B.n462 VSUBS 0.009626f
C503 B.n463 VSUBS 0.009626f
C504 B.n464 VSUBS 0.009626f
C505 B.n465 VSUBS 0.009626f
C506 B.n466 VSUBS 0.009626f
C507 B.n467 VSUBS 0.009626f
C508 B.n468 VSUBS 0.009626f
C509 B.n469 VSUBS 0.009626f
C510 B.n470 VSUBS 0.009626f
C511 B.n471 VSUBS 0.009626f
C512 B.n472 VSUBS 0.009626f
C513 B.n473 VSUBS 0.009626f
C514 B.n474 VSUBS 0.009626f
C515 B.n475 VSUBS 0.009626f
C516 B.n476 VSUBS 0.009626f
C517 B.n477 VSUBS 0.009626f
C518 B.n478 VSUBS 0.009626f
C519 B.n479 VSUBS 0.009626f
C520 B.n480 VSUBS 0.009626f
C521 B.n481 VSUBS 0.009626f
C522 B.n482 VSUBS 0.009626f
C523 B.n483 VSUBS 0.009626f
C524 B.n484 VSUBS 0.009626f
C525 B.n485 VSUBS 0.009626f
C526 B.n486 VSUBS 0.009626f
C527 B.n487 VSUBS 0.009626f
C528 B.n488 VSUBS 0.009626f
C529 B.n489 VSUBS 0.009626f
C530 B.n490 VSUBS 0.009626f
C531 B.n491 VSUBS 0.009626f
C532 B.n492 VSUBS 0.009626f
C533 B.n493 VSUBS 0.009626f
C534 B.n494 VSUBS 0.009626f
C535 B.n495 VSUBS 0.009626f
C536 B.n496 VSUBS 0.009626f
C537 B.n497 VSUBS 0.009626f
C538 B.n498 VSUBS 0.009626f
C539 B.n499 VSUBS 0.009626f
C540 B.n500 VSUBS 0.023458f
C541 B.n501 VSUBS 0.022341f
C542 B.n502 VSUBS 0.02324f
C543 B.n503 VSUBS 0.009626f
C544 B.n504 VSUBS 0.009626f
C545 B.n505 VSUBS 0.009626f
C546 B.n506 VSUBS 0.009626f
C547 B.n507 VSUBS 0.009626f
C548 B.n508 VSUBS 0.009626f
C549 B.n509 VSUBS 0.009626f
C550 B.n510 VSUBS 0.009626f
C551 B.n511 VSUBS 0.009626f
C552 B.n512 VSUBS 0.009626f
C553 B.n513 VSUBS 0.009626f
C554 B.n514 VSUBS 0.009626f
C555 B.n515 VSUBS 0.009626f
C556 B.n516 VSUBS 0.009626f
C557 B.n517 VSUBS 0.009626f
C558 B.n518 VSUBS 0.009626f
C559 B.n519 VSUBS 0.009626f
C560 B.n520 VSUBS 0.009626f
C561 B.n521 VSUBS 0.009626f
C562 B.n522 VSUBS 0.009626f
C563 B.n523 VSUBS 0.009626f
C564 B.n524 VSUBS 0.009626f
C565 B.n525 VSUBS 0.009626f
C566 B.n526 VSUBS 0.009626f
C567 B.n527 VSUBS 0.009626f
C568 B.n528 VSUBS 0.009626f
C569 B.n529 VSUBS 0.009626f
C570 B.n530 VSUBS 0.009626f
C571 B.n531 VSUBS 0.009626f
C572 B.n532 VSUBS 0.009626f
C573 B.n533 VSUBS 0.009626f
C574 B.n534 VSUBS 0.009626f
C575 B.n535 VSUBS 0.006653f
C576 B.n536 VSUBS 0.022302f
C577 B.n537 VSUBS 0.007785f
C578 B.n538 VSUBS 0.009626f
C579 B.n539 VSUBS 0.009626f
C580 B.n540 VSUBS 0.009626f
C581 B.n541 VSUBS 0.009626f
C582 B.n542 VSUBS 0.009626f
C583 B.n543 VSUBS 0.009626f
C584 B.n544 VSUBS 0.009626f
C585 B.n545 VSUBS 0.009626f
C586 B.n546 VSUBS 0.009626f
C587 B.n547 VSUBS 0.009626f
C588 B.n548 VSUBS 0.009626f
C589 B.n549 VSUBS 0.007785f
C590 B.n550 VSUBS 0.009626f
C591 B.n551 VSUBS 0.009626f
C592 B.n552 VSUBS 0.009626f
C593 B.n553 VSUBS 0.009626f
C594 B.n554 VSUBS 0.009626f
C595 B.n555 VSUBS 0.009626f
C596 B.n556 VSUBS 0.009626f
C597 B.n557 VSUBS 0.009626f
C598 B.n558 VSUBS 0.009626f
C599 B.n559 VSUBS 0.009626f
C600 B.n560 VSUBS 0.009626f
C601 B.n561 VSUBS 0.009626f
C602 B.n562 VSUBS 0.009626f
C603 B.n563 VSUBS 0.009626f
C604 B.n564 VSUBS 0.009626f
C605 B.n565 VSUBS 0.009626f
C606 B.n566 VSUBS 0.009626f
C607 B.n567 VSUBS 0.009626f
C608 B.n568 VSUBS 0.009626f
C609 B.n569 VSUBS 0.009626f
C610 B.n570 VSUBS 0.009626f
C611 B.n571 VSUBS 0.009626f
C612 B.n572 VSUBS 0.009626f
C613 B.n573 VSUBS 0.009626f
C614 B.n574 VSUBS 0.009626f
C615 B.n575 VSUBS 0.009626f
C616 B.n576 VSUBS 0.009626f
C617 B.n577 VSUBS 0.009626f
C618 B.n578 VSUBS 0.009626f
C619 B.n579 VSUBS 0.009626f
C620 B.n580 VSUBS 0.009626f
C621 B.n581 VSUBS 0.009626f
C622 B.n582 VSUBS 0.009626f
C623 B.n583 VSUBS 0.009626f
C624 B.n584 VSUBS 0.02324f
C625 B.n585 VSUBS 0.022341f
C626 B.n586 VSUBS 0.022341f
C627 B.n587 VSUBS 0.009626f
C628 B.n588 VSUBS 0.009626f
C629 B.n589 VSUBS 0.009626f
C630 B.n590 VSUBS 0.009626f
C631 B.n591 VSUBS 0.009626f
C632 B.n592 VSUBS 0.009626f
C633 B.n593 VSUBS 0.009626f
C634 B.n594 VSUBS 0.009626f
C635 B.n595 VSUBS 0.009626f
C636 B.n596 VSUBS 0.009626f
C637 B.n597 VSUBS 0.009626f
C638 B.n598 VSUBS 0.009626f
C639 B.n599 VSUBS 0.009626f
C640 B.n600 VSUBS 0.009626f
C641 B.n601 VSUBS 0.009626f
C642 B.n602 VSUBS 0.009626f
C643 B.n603 VSUBS 0.009626f
C644 B.n604 VSUBS 0.009626f
C645 B.n605 VSUBS 0.009626f
C646 B.n606 VSUBS 0.009626f
C647 B.n607 VSUBS 0.009626f
C648 B.n608 VSUBS 0.009626f
C649 B.n609 VSUBS 0.009626f
C650 B.n610 VSUBS 0.009626f
C651 B.n611 VSUBS 0.009626f
C652 B.n612 VSUBS 0.009626f
C653 B.n613 VSUBS 0.009626f
C654 B.n614 VSUBS 0.009626f
C655 B.n615 VSUBS 0.009626f
C656 B.n616 VSUBS 0.009626f
C657 B.n617 VSUBS 0.009626f
C658 B.n618 VSUBS 0.009626f
C659 B.n619 VSUBS 0.009626f
C660 B.n620 VSUBS 0.009626f
C661 B.n621 VSUBS 0.009626f
C662 B.n622 VSUBS 0.009626f
C663 B.n623 VSUBS 0.009626f
C664 B.n624 VSUBS 0.009626f
C665 B.n625 VSUBS 0.009626f
C666 B.n626 VSUBS 0.009626f
C667 B.n627 VSUBS 0.009626f
C668 B.n628 VSUBS 0.009626f
C669 B.n629 VSUBS 0.009626f
C670 B.n630 VSUBS 0.009626f
C671 B.n631 VSUBS 0.009626f
C672 B.n632 VSUBS 0.009626f
C673 B.n633 VSUBS 0.009626f
C674 B.n634 VSUBS 0.009626f
C675 B.n635 VSUBS 0.009626f
C676 B.n636 VSUBS 0.009626f
C677 B.n637 VSUBS 0.009626f
C678 B.n638 VSUBS 0.009626f
C679 B.n639 VSUBS 0.009626f
C680 B.n640 VSUBS 0.009626f
C681 B.n641 VSUBS 0.009626f
C682 B.n642 VSUBS 0.009626f
C683 B.n643 VSUBS 0.009626f
C684 B.n644 VSUBS 0.009626f
C685 B.n645 VSUBS 0.009626f
C686 B.n646 VSUBS 0.009626f
C687 B.n647 VSUBS 0.009626f
C688 B.n648 VSUBS 0.009626f
C689 B.n649 VSUBS 0.009626f
C690 B.n650 VSUBS 0.009626f
C691 B.n651 VSUBS 0.009626f
C692 B.n652 VSUBS 0.009626f
C693 B.n653 VSUBS 0.009626f
C694 B.n654 VSUBS 0.009626f
C695 B.n655 VSUBS 0.009626f
C696 B.n656 VSUBS 0.009626f
C697 B.n657 VSUBS 0.009626f
C698 B.n658 VSUBS 0.009626f
C699 B.n659 VSUBS 0.009626f
C700 B.n660 VSUBS 0.009626f
C701 B.n661 VSUBS 0.009626f
C702 B.n662 VSUBS 0.009626f
C703 B.n663 VSUBS 0.009626f
C704 B.n664 VSUBS 0.009626f
C705 B.n665 VSUBS 0.009626f
C706 B.n666 VSUBS 0.009626f
C707 B.n667 VSUBS 0.021796f
C708 VDD1.t0 VSUBS 0.109527f
C709 VDD1.t6 VSUBS 0.109527f
C710 VDD1.n0 VSUBS 0.721318f
C711 VDD1.t2 VSUBS 0.109527f
C712 VDD1.t3 VSUBS 0.109527f
C713 VDD1.n1 VSUBS 0.720339f
C714 VDD1.t5 VSUBS 0.109527f
C715 VDD1.t4 VSUBS 0.109527f
C716 VDD1.n2 VSUBS 0.720339f
C717 VDD1.n3 VSUBS 3.39835f
C718 VDD1.t1 VSUBS 0.109527f
C719 VDD1.t7 VSUBS 0.109527f
C720 VDD1.n4 VSUBS 0.71055f
C721 VDD1.n5 VSUBS 2.7182f
C722 VP.t3 VSUBS 1.68119f
C723 VP.n0 VSUBS 0.786394f
C724 VP.n1 VSUBS 0.040826f
C725 VP.n2 VSUBS 0.072092f
C726 VP.n3 VSUBS 0.040826f
C727 VP.t2 VSUBS 1.68119f
C728 VP.n4 VSUBS 0.075708f
C729 VP.n5 VSUBS 0.040826f
C730 VP.n6 VSUBS 0.061505f
C731 VP.n7 VSUBS 0.040826f
C732 VP.n8 VSUBS 0.042707f
C733 VP.n9 VSUBS 0.065882f
C734 VP.t5 VSUBS 1.68119f
C735 VP.t0 VSUBS 1.68119f
C736 VP.n10 VSUBS 0.786394f
C737 VP.n11 VSUBS 0.040826f
C738 VP.n12 VSUBS 0.072092f
C739 VP.n13 VSUBS 0.040826f
C740 VP.t6 VSUBS 1.68119f
C741 VP.n14 VSUBS 0.075708f
C742 VP.n15 VSUBS 0.040826f
C743 VP.n16 VSUBS 0.061505f
C744 VP.t7 VSUBS 2.03671f
C745 VP.t1 VSUBS 1.68119f
C746 VP.n17 VSUBS 0.761795f
C747 VP.n18 VSUBS 0.729872f
C748 VP.n19 VSUBS 0.430651f
C749 VP.n20 VSUBS 0.040826f
C750 VP.n21 VSUBS 0.075708f
C751 VP.n22 VSUBS 0.059347f
C752 VP.n23 VSUBS 0.059347f
C753 VP.n24 VSUBS 0.040826f
C754 VP.n25 VSUBS 0.040826f
C755 VP.n26 VSUBS 0.040826f
C756 VP.n27 VSUBS 0.061505f
C757 VP.n28 VSUBS 0.633241f
C758 VP.n29 VSUBS 0.052535f
C759 VP.n30 VSUBS 0.075708f
C760 VP.n31 VSUBS 0.040826f
C761 VP.n32 VSUBS 0.040826f
C762 VP.n33 VSUBS 0.040826f
C763 VP.n34 VSUBS 0.042707f
C764 VP.n35 VSUBS 0.079603f
C765 VP.n36 VSUBS 0.070476f
C766 VP.n37 VSUBS 0.065882f
C767 VP.n38 VSUBS 2.10173f
C768 VP.n39 VSUBS 2.13303f
C769 VP.n40 VSUBS 0.786394f
C770 VP.n41 VSUBS 0.070476f
C771 VP.n42 VSUBS 0.079603f
C772 VP.n43 VSUBS 0.040826f
C773 VP.n44 VSUBS 0.040826f
C774 VP.n45 VSUBS 0.040826f
C775 VP.n46 VSUBS 0.072092f
C776 VP.n47 VSUBS 0.075708f
C777 VP.t4 VSUBS 1.68119f
C778 VP.n48 VSUBS 0.633241f
C779 VP.n49 VSUBS 0.052535f
C780 VP.n50 VSUBS 0.040826f
C781 VP.n51 VSUBS 0.040826f
C782 VP.n52 VSUBS 0.040826f
C783 VP.n53 VSUBS 0.075708f
C784 VP.n54 VSUBS 0.059347f
C785 VP.n55 VSUBS 0.059347f
C786 VP.n56 VSUBS 0.040826f
C787 VP.n57 VSUBS 0.040826f
C788 VP.n58 VSUBS 0.040826f
C789 VP.n59 VSUBS 0.061505f
C790 VP.n60 VSUBS 0.633241f
C791 VP.n61 VSUBS 0.052535f
C792 VP.n62 VSUBS 0.075708f
C793 VP.n63 VSUBS 0.040826f
C794 VP.n64 VSUBS 0.040826f
C795 VP.n65 VSUBS 0.040826f
C796 VP.n66 VSUBS 0.042707f
C797 VP.n67 VSUBS 0.079603f
C798 VP.n68 VSUBS 0.070476f
C799 VP.n69 VSUBS 0.065882f
C800 VP.n70 VSUBS 0.080276f
C801 VDD2.t6 VSUBS 0.107393f
C802 VDD2.t0 VSUBS 0.107393f
C803 VDD2.n0 VSUBS 0.706308f
C804 VDD2.t3 VSUBS 0.107393f
C805 VDD2.t7 VSUBS 0.107393f
C806 VDD2.n1 VSUBS 0.706308f
C807 VDD2.n2 VSUBS 3.28154f
C808 VDD2.t2 VSUBS 0.107393f
C809 VDD2.t5 VSUBS 0.107393f
C810 VDD2.n3 VSUBS 0.696713f
C811 VDD2.n4 VSUBS 2.63534f
C812 VDD2.t1 VSUBS 0.107393f
C813 VDD2.t4 VSUBS 0.107393f
C814 VDD2.n5 VSUBS 0.706278f
C815 VTAIL.t12 VSUBS 0.133121f
C816 VTAIL.t14 VSUBS 0.133121f
C817 VTAIL.n0 VSUBS 0.761222f
C818 VTAIL.n1 VSUBS 0.807455f
C819 VTAIL.t13 VSUBS 1.05496f
C820 VTAIL.n2 VSUBS 0.916679f
C821 VTAIL.t6 VSUBS 1.05496f
C822 VTAIL.n3 VSUBS 0.916679f
C823 VTAIL.t1 VSUBS 0.133121f
C824 VTAIL.t0 VSUBS 0.133121f
C825 VTAIL.n4 VSUBS 0.761222f
C826 VTAIL.n5 VSUBS 1.06252f
C827 VTAIL.t5 VSUBS 1.05496f
C828 VTAIL.n6 VSUBS 2.00842f
C829 VTAIL.t8 VSUBS 1.05496f
C830 VTAIL.n7 VSUBS 2.00841f
C831 VTAIL.t11 VSUBS 0.133121f
C832 VTAIL.t15 VSUBS 0.133121f
C833 VTAIL.n8 VSUBS 0.761227f
C834 VTAIL.n9 VSUBS 1.06252f
C835 VTAIL.t9 VSUBS 1.05496f
C836 VTAIL.n10 VSUBS 0.916674f
C837 VTAIL.t2 VSUBS 1.05496f
C838 VTAIL.n11 VSUBS 0.916674f
C839 VTAIL.t3 VSUBS 0.133121f
C840 VTAIL.t4 VSUBS 0.133121f
C841 VTAIL.n12 VSUBS 0.761227f
C842 VTAIL.n13 VSUBS 1.06252f
C843 VTAIL.t7 VSUBS 1.05496f
C844 VTAIL.n14 VSUBS 2.00842f
C845 VTAIL.t10 VSUBS 1.05496f
C846 VTAIL.n15 VSUBS 2.00278f
C847 VN.t0 VSUBS 1.50142f
C848 VN.n0 VSUBS 0.702305f
C849 VN.n1 VSUBS 0.036461f
C850 VN.n2 VSUBS 0.064383f
C851 VN.n3 VSUBS 0.036461f
C852 VN.t4 VSUBS 1.50142f
C853 VN.n4 VSUBS 0.067613f
C854 VN.n5 VSUBS 0.036461f
C855 VN.n6 VSUBS 0.054929f
C856 VN.t7 VSUBS 1.50142f
C857 VN.n7 VSUBS 0.680336f
C858 VN.t1 VSUBS 1.81892f
C859 VN.n8 VSUBS 0.651826f
C860 VN.n9 VSUBS 0.384601f
C861 VN.n10 VSUBS 0.036461f
C862 VN.n11 VSUBS 0.067613f
C863 VN.n12 VSUBS 0.053001f
C864 VN.n13 VSUBS 0.053001f
C865 VN.n14 VSUBS 0.036461f
C866 VN.n15 VSUBS 0.036461f
C867 VN.n16 VSUBS 0.036461f
C868 VN.n17 VSUBS 0.054929f
C869 VN.n18 VSUBS 0.565529f
C870 VN.n19 VSUBS 0.046918f
C871 VN.n20 VSUBS 0.067613f
C872 VN.n21 VSUBS 0.036461f
C873 VN.n22 VSUBS 0.036461f
C874 VN.n23 VSUBS 0.036461f
C875 VN.n24 VSUBS 0.03814f
C876 VN.n25 VSUBS 0.071091f
C877 VN.n26 VSUBS 0.06294f
C878 VN.n27 VSUBS 0.058837f
C879 VN.n28 VSUBS 0.071692f
C880 VN.t5 VSUBS 1.50142f
C881 VN.n29 VSUBS 0.702305f
C882 VN.n30 VSUBS 0.036461f
C883 VN.n31 VSUBS 0.064383f
C884 VN.n32 VSUBS 0.036461f
C885 VN.t2 VSUBS 1.50142f
C886 VN.n33 VSUBS 0.067613f
C887 VN.n34 VSUBS 0.036461f
C888 VN.n35 VSUBS 0.054929f
C889 VN.t3 VSUBS 1.81892f
C890 VN.t6 VSUBS 1.50142f
C891 VN.n36 VSUBS 0.680336f
C892 VN.n37 VSUBS 0.651826f
C893 VN.n38 VSUBS 0.384601f
C894 VN.n39 VSUBS 0.036461f
C895 VN.n40 VSUBS 0.067613f
C896 VN.n41 VSUBS 0.053001f
C897 VN.n42 VSUBS 0.053001f
C898 VN.n43 VSUBS 0.036461f
C899 VN.n44 VSUBS 0.036461f
C900 VN.n45 VSUBS 0.036461f
C901 VN.n46 VSUBS 0.054929f
C902 VN.n47 VSUBS 0.565529f
C903 VN.n48 VSUBS 0.046918f
C904 VN.n49 VSUBS 0.067613f
C905 VN.n50 VSUBS 0.036461f
C906 VN.n51 VSUBS 0.036461f
C907 VN.n52 VSUBS 0.036461f
C908 VN.n53 VSUBS 0.03814f
C909 VN.n54 VSUBS 0.071091f
C910 VN.n55 VSUBS 0.06294f
C911 VN.n56 VSUBS 0.058837f
C912 VN.n57 VSUBS 1.89225f
.ends

