* NGSPICE file created from diff_pair_sample_0327.ext - technology: sky130A

.subckt diff_pair_sample_0327 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1814_n2488# sky130_fd_pr__pfet_01v8 ad=2.964 pd=15.98 as=0 ps=0 w=7.6 l=1.78
X1 VDD1.t1 VP.t0 VTAIL.t2 w_n1814_n2488# sky130_fd_pr__pfet_01v8 ad=2.964 pd=15.98 as=2.964 ps=15.98 w=7.6 l=1.78
X2 B.t8 B.t6 B.t7 w_n1814_n2488# sky130_fd_pr__pfet_01v8 ad=2.964 pd=15.98 as=0 ps=0 w=7.6 l=1.78
X3 VDD2.t1 VN.t0 VTAIL.t1 w_n1814_n2488# sky130_fd_pr__pfet_01v8 ad=2.964 pd=15.98 as=2.964 ps=15.98 w=7.6 l=1.78
X4 VDD2.t0 VN.t1 VTAIL.t0 w_n1814_n2488# sky130_fd_pr__pfet_01v8 ad=2.964 pd=15.98 as=2.964 ps=15.98 w=7.6 l=1.78
X5 VDD1.t0 VP.t1 VTAIL.t3 w_n1814_n2488# sky130_fd_pr__pfet_01v8 ad=2.964 pd=15.98 as=2.964 ps=15.98 w=7.6 l=1.78
X6 B.t5 B.t3 B.t4 w_n1814_n2488# sky130_fd_pr__pfet_01v8 ad=2.964 pd=15.98 as=0 ps=0 w=7.6 l=1.78
X7 B.t2 B.t0 B.t1 w_n1814_n2488# sky130_fd_pr__pfet_01v8 ad=2.964 pd=15.98 as=0 ps=0 w=7.6 l=1.78
R0 B.n249 B.n248 585
R1 B.n247 B.n72 585
R2 B.n246 B.n245 585
R3 B.n244 B.n73 585
R4 B.n243 B.n242 585
R5 B.n241 B.n74 585
R6 B.n240 B.n239 585
R7 B.n238 B.n75 585
R8 B.n237 B.n236 585
R9 B.n235 B.n76 585
R10 B.n234 B.n233 585
R11 B.n232 B.n77 585
R12 B.n231 B.n230 585
R13 B.n229 B.n78 585
R14 B.n228 B.n227 585
R15 B.n226 B.n79 585
R16 B.n225 B.n224 585
R17 B.n223 B.n80 585
R18 B.n222 B.n221 585
R19 B.n220 B.n81 585
R20 B.n219 B.n218 585
R21 B.n217 B.n82 585
R22 B.n216 B.n215 585
R23 B.n214 B.n83 585
R24 B.n213 B.n212 585
R25 B.n211 B.n84 585
R26 B.n210 B.n209 585
R27 B.n208 B.n85 585
R28 B.n207 B.n206 585
R29 B.n204 B.n86 585
R30 B.n203 B.n202 585
R31 B.n201 B.n89 585
R32 B.n200 B.n199 585
R33 B.n198 B.n90 585
R34 B.n197 B.n196 585
R35 B.n195 B.n91 585
R36 B.n194 B.n193 585
R37 B.n192 B.n92 585
R38 B.n190 B.n189 585
R39 B.n188 B.n95 585
R40 B.n187 B.n186 585
R41 B.n185 B.n96 585
R42 B.n184 B.n183 585
R43 B.n182 B.n97 585
R44 B.n181 B.n180 585
R45 B.n179 B.n98 585
R46 B.n178 B.n177 585
R47 B.n176 B.n99 585
R48 B.n175 B.n174 585
R49 B.n173 B.n100 585
R50 B.n172 B.n171 585
R51 B.n170 B.n101 585
R52 B.n169 B.n168 585
R53 B.n167 B.n102 585
R54 B.n166 B.n165 585
R55 B.n164 B.n103 585
R56 B.n163 B.n162 585
R57 B.n161 B.n104 585
R58 B.n160 B.n159 585
R59 B.n158 B.n105 585
R60 B.n157 B.n156 585
R61 B.n155 B.n106 585
R62 B.n154 B.n153 585
R63 B.n152 B.n107 585
R64 B.n151 B.n150 585
R65 B.n149 B.n108 585
R66 B.n148 B.n147 585
R67 B.n250 B.n71 585
R68 B.n252 B.n251 585
R69 B.n253 B.n70 585
R70 B.n255 B.n254 585
R71 B.n256 B.n69 585
R72 B.n258 B.n257 585
R73 B.n259 B.n68 585
R74 B.n261 B.n260 585
R75 B.n262 B.n67 585
R76 B.n264 B.n263 585
R77 B.n265 B.n66 585
R78 B.n267 B.n266 585
R79 B.n268 B.n65 585
R80 B.n270 B.n269 585
R81 B.n271 B.n64 585
R82 B.n273 B.n272 585
R83 B.n274 B.n63 585
R84 B.n276 B.n275 585
R85 B.n277 B.n62 585
R86 B.n279 B.n278 585
R87 B.n280 B.n61 585
R88 B.n282 B.n281 585
R89 B.n283 B.n60 585
R90 B.n285 B.n284 585
R91 B.n286 B.n59 585
R92 B.n288 B.n287 585
R93 B.n289 B.n58 585
R94 B.n291 B.n290 585
R95 B.n292 B.n57 585
R96 B.n294 B.n293 585
R97 B.n295 B.n56 585
R98 B.n297 B.n296 585
R99 B.n298 B.n55 585
R100 B.n300 B.n299 585
R101 B.n301 B.n54 585
R102 B.n303 B.n302 585
R103 B.n304 B.n53 585
R104 B.n306 B.n305 585
R105 B.n307 B.n52 585
R106 B.n309 B.n308 585
R107 B.n310 B.n51 585
R108 B.n312 B.n311 585
R109 B.n413 B.n12 585
R110 B.n412 B.n411 585
R111 B.n410 B.n13 585
R112 B.n409 B.n408 585
R113 B.n407 B.n14 585
R114 B.n406 B.n405 585
R115 B.n404 B.n15 585
R116 B.n403 B.n402 585
R117 B.n401 B.n16 585
R118 B.n400 B.n399 585
R119 B.n398 B.n17 585
R120 B.n397 B.n396 585
R121 B.n395 B.n18 585
R122 B.n394 B.n393 585
R123 B.n392 B.n19 585
R124 B.n391 B.n390 585
R125 B.n389 B.n20 585
R126 B.n388 B.n387 585
R127 B.n386 B.n21 585
R128 B.n385 B.n384 585
R129 B.n383 B.n22 585
R130 B.n382 B.n381 585
R131 B.n380 B.n23 585
R132 B.n379 B.n378 585
R133 B.n377 B.n24 585
R134 B.n376 B.n375 585
R135 B.n374 B.n25 585
R136 B.n373 B.n372 585
R137 B.n371 B.n26 585
R138 B.n370 B.n369 585
R139 B.n368 B.n27 585
R140 B.n367 B.n366 585
R141 B.n365 B.n31 585
R142 B.n364 B.n363 585
R143 B.n362 B.n32 585
R144 B.n361 B.n360 585
R145 B.n359 B.n33 585
R146 B.n358 B.n357 585
R147 B.n355 B.n34 585
R148 B.n354 B.n353 585
R149 B.n352 B.n37 585
R150 B.n351 B.n350 585
R151 B.n349 B.n38 585
R152 B.n348 B.n347 585
R153 B.n346 B.n39 585
R154 B.n345 B.n344 585
R155 B.n343 B.n40 585
R156 B.n342 B.n341 585
R157 B.n340 B.n41 585
R158 B.n339 B.n338 585
R159 B.n337 B.n42 585
R160 B.n336 B.n335 585
R161 B.n334 B.n43 585
R162 B.n333 B.n332 585
R163 B.n331 B.n44 585
R164 B.n330 B.n329 585
R165 B.n328 B.n45 585
R166 B.n327 B.n326 585
R167 B.n325 B.n46 585
R168 B.n324 B.n323 585
R169 B.n322 B.n47 585
R170 B.n321 B.n320 585
R171 B.n319 B.n48 585
R172 B.n318 B.n317 585
R173 B.n316 B.n49 585
R174 B.n315 B.n314 585
R175 B.n313 B.n50 585
R176 B.n415 B.n414 585
R177 B.n416 B.n11 585
R178 B.n418 B.n417 585
R179 B.n419 B.n10 585
R180 B.n421 B.n420 585
R181 B.n422 B.n9 585
R182 B.n424 B.n423 585
R183 B.n425 B.n8 585
R184 B.n427 B.n426 585
R185 B.n428 B.n7 585
R186 B.n430 B.n429 585
R187 B.n431 B.n6 585
R188 B.n433 B.n432 585
R189 B.n434 B.n5 585
R190 B.n436 B.n435 585
R191 B.n437 B.n4 585
R192 B.n439 B.n438 585
R193 B.n440 B.n3 585
R194 B.n442 B.n441 585
R195 B.n443 B.n0 585
R196 B.n2 B.n1 585
R197 B.n119 B.n118 585
R198 B.n121 B.n120 585
R199 B.n122 B.n117 585
R200 B.n124 B.n123 585
R201 B.n125 B.n116 585
R202 B.n127 B.n126 585
R203 B.n128 B.n115 585
R204 B.n130 B.n129 585
R205 B.n131 B.n114 585
R206 B.n133 B.n132 585
R207 B.n134 B.n113 585
R208 B.n136 B.n135 585
R209 B.n137 B.n112 585
R210 B.n139 B.n138 585
R211 B.n140 B.n111 585
R212 B.n142 B.n141 585
R213 B.n143 B.n110 585
R214 B.n145 B.n144 585
R215 B.n146 B.n109 585
R216 B.n147 B.n146 497.305
R217 B.n250 B.n249 497.305
R218 B.n311 B.n50 497.305
R219 B.n414 B.n413 497.305
R220 B.n93 B.t3 309.248
R221 B.n87 B.t6 309.248
R222 B.n35 B.t9 309.248
R223 B.n28 B.t0 309.248
R224 B.n445 B.n444 256.663
R225 B.n444 B.n443 235.042
R226 B.n444 B.n2 235.042
R227 B.n147 B.n108 163.367
R228 B.n151 B.n108 163.367
R229 B.n152 B.n151 163.367
R230 B.n153 B.n152 163.367
R231 B.n153 B.n106 163.367
R232 B.n157 B.n106 163.367
R233 B.n158 B.n157 163.367
R234 B.n159 B.n158 163.367
R235 B.n159 B.n104 163.367
R236 B.n163 B.n104 163.367
R237 B.n164 B.n163 163.367
R238 B.n165 B.n164 163.367
R239 B.n165 B.n102 163.367
R240 B.n169 B.n102 163.367
R241 B.n170 B.n169 163.367
R242 B.n171 B.n170 163.367
R243 B.n171 B.n100 163.367
R244 B.n175 B.n100 163.367
R245 B.n176 B.n175 163.367
R246 B.n177 B.n176 163.367
R247 B.n177 B.n98 163.367
R248 B.n181 B.n98 163.367
R249 B.n182 B.n181 163.367
R250 B.n183 B.n182 163.367
R251 B.n183 B.n96 163.367
R252 B.n187 B.n96 163.367
R253 B.n188 B.n187 163.367
R254 B.n189 B.n188 163.367
R255 B.n189 B.n92 163.367
R256 B.n194 B.n92 163.367
R257 B.n195 B.n194 163.367
R258 B.n196 B.n195 163.367
R259 B.n196 B.n90 163.367
R260 B.n200 B.n90 163.367
R261 B.n201 B.n200 163.367
R262 B.n202 B.n201 163.367
R263 B.n202 B.n86 163.367
R264 B.n207 B.n86 163.367
R265 B.n208 B.n207 163.367
R266 B.n209 B.n208 163.367
R267 B.n209 B.n84 163.367
R268 B.n213 B.n84 163.367
R269 B.n214 B.n213 163.367
R270 B.n215 B.n214 163.367
R271 B.n215 B.n82 163.367
R272 B.n219 B.n82 163.367
R273 B.n220 B.n219 163.367
R274 B.n221 B.n220 163.367
R275 B.n221 B.n80 163.367
R276 B.n225 B.n80 163.367
R277 B.n226 B.n225 163.367
R278 B.n227 B.n226 163.367
R279 B.n227 B.n78 163.367
R280 B.n231 B.n78 163.367
R281 B.n232 B.n231 163.367
R282 B.n233 B.n232 163.367
R283 B.n233 B.n76 163.367
R284 B.n237 B.n76 163.367
R285 B.n238 B.n237 163.367
R286 B.n239 B.n238 163.367
R287 B.n239 B.n74 163.367
R288 B.n243 B.n74 163.367
R289 B.n244 B.n243 163.367
R290 B.n245 B.n244 163.367
R291 B.n245 B.n72 163.367
R292 B.n249 B.n72 163.367
R293 B.n311 B.n310 163.367
R294 B.n310 B.n309 163.367
R295 B.n309 B.n52 163.367
R296 B.n305 B.n52 163.367
R297 B.n305 B.n304 163.367
R298 B.n304 B.n303 163.367
R299 B.n303 B.n54 163.367
R300 B.n299 B.n54 163.367
R301 B.n299 B.n298 163.367
R302 B.n298 B.n297 163.367
R303 B.n297 B.n56 163.367
R304 B.n293 B.n56 163.367
R305 B.n293 B.n292 163.367
R306 B.n292 B.n291 163.367
R307 B.n291 B.n58 163.367
R308 B.n287 B.n58 163.367
R309 B.n287 B.n286 163.367
R310 B.n286 B.n285 163.367
R311 B.n285 B.n60 163.367
R312 B.n281 B.n60 163.367
R313 B.n281 B.n280 163.367
R314 B.n280 B.n279 163.367
R315 B.n279 B.n62 163.367
R316 B.n275 B.n62 163.367
R317 B.n275 B.n274 163.367
R318 B.n274 B.n273 163.367
R319 B.n273 B.n64 163.367
R320 B.n269 B.n64 163.367
R321 B.n269 B.n268 163.367
R322 B.n268 B.n267 163.367
R323 B.n267 B.n66 163.367
R324 B.n263 B.n66 163.367
R325 B.n263 B.n262 163.367
R326 B.n262 B.n261 163.367
R327 B.n261 B.n68 163.367
R328 B.n257 B.n68 163.367
R329 B.n257 B.n256 163.367
R330 B.n256 B.n255 163.367
R331 B.n255 B.n70 163.367
R332 B.n251 B.n70 163.367
R333 B.n251 B.n250 163.367
R334 B.n413 B.n412 163.367
R335 B.n412 B.n13 163.367
R336 B.n408 B.n13 163.367
R337 B.n408 B.n407 163.367
R338 B.n407 B.n406 163.367
R339 B.n406 B.n15 163.367
R340 B.n402 B.n15 163.367
R341 B.n402 B.n401 163.367
R342 B.n401 B.n400 163.367
R343 B.n400 B.n17 163.367
R344 B.n396 B.n17 163.367
R345 B.n396 B.n395 163.367
R346 B.n395 B.n394 163.367
R347 B.n394 B.n19 163.367
R348 B.n390 B.n19 163.367
R349 B.n390 B.n389 163.367
R350 B.n389 B.n388 163.367
R351 B.n388 B.n21 163.367
R352 B.n384 B.n21 163.367
R353 B.n384 B.n383 163.367
R354 B.n383 B.n382 163.367
R355 B.n382 B.n23 163.367
R356 B.n378 B.n23 163.367
R357 B.n378 B.n377 163.367
R358 B.n377 B.n376 163.367
R359 B.n376 B.n25 163.367
R360 B.n372 B.n25 163.367
R361 B.n372 B.n371 163.367
R362 B.n371 B.n370 163.367
R363 B.n370 B.n27 163.367
R364 B.n366 B.n27 163.367
R365 B.n366 B.n365 163.367
R366 B.n365 B.n364 163.367
R367 B.n364 B.n32 163.367
R368 B.n360 B.n32 163.367
R369 B.n360 B.n359 163.367
R370 B.n359 B.n358 163.367
R371 B.n358 B.n34 163.367
R372 B.n353 B.n34 163.367
R373 B.n353 B.n352 163.367
R374 B.n352 B.n351 163.367
R375 B.n351 B.n38 163.367
R376 B.n347 B.n38 163.367
R377 B.n347 B.n346 163.367
R378 B.n346 B.n345 163.367
R379 B.n345 B.n40 163.367
R380 B.n341 B.n40 163.367
R381 B.n341 B.n340 163.367
R382 B.n340 B.n339 163.367
R383 B.n339 B.n42 163.367
R384 B.n335 B.n42 163.367
R385 B.n335 B.n334 163.367
R386 B.n334 B.n333 163.367
R387 B.n333 B.n44 163.367
R388 B.n329 B.n44 163.367
R389 B.n329 B.n328 163.367
R390 B.n328 B.n327 163.367
R391 B.n327 B.n46 163.367
R392 B.n323 B.n46 163.367
R393 B.n323 B.n322 163.367
R394 B.n322 B.n321 163.367
R395 B.n321 B.n48 163.367
R396 B.n317 B.n48 163.367
R397 B.n317 B.n316 163.367
R398 B.n316 B.n315 163.367
R399 B.n315 B.n50 163.367
R400 B.n414 B.n11 163.367
R401 B.n418 B.n11 163.367
R402 B.n419 B.n418 163.367
R403 B.n420 B.n419 163.367
R404 B.n420 B.n9 163.367
R405 B.n424 B.n9 163.367
R406 B.n425 B.n424 163.367
R407 B.n426 B.n425 163.367
R408 B.n426 B.n7 163.367
R409 B.n430 B.n7 163.367
R410 B.n431 B.n430 163.367
R411 B.n432 B.n431 163.367
R412 B.n432 B.n5 163.367
R413 B.n436 B.n5 163.367
R414 B.n437 B.n436 163.367
R415 B.n438 B.n437 163.367
R416 B.n438 B.n3 163.367
R417 B.n442 B.n3 163.367
R418 B.n443 B.n442 163.367
R419 B.n118 B.n2 163.367
R420 B.n121 B.n118 163.367
R421 B.n122 B.n121 163.367
R422 B.n123 B.n122 163.367
R423 B.n123 B.n116 163.367
R424 B.n127 B.n116 163.367
R425 B.n128 B.n127 163.367
R426 B.n129 B.n128 163.367
R427 B.n129 B.n114 163.367
R428 B.n133 B.n114 163.367
R429 B.n134 B.n133 163.367
R430 B.n135 B.n134 163.367
R431 B.n135 B.n112 163.367
R432 B.n139 B.n112 163.367
R433 B.n140 B.n139 163.367
R434 B.n141 B.n140 163.367
R435 B.n141 B.n110 163.367
R436 B.n145 B.n110 163.367
R437 B.n146 B.n145 163.367
R438 B.n87 B.t7 152.232
R439 B.n35 B.t11 152.232
R440 B.n93 B.t4 152.225
R441 B.n28 B.t2 152.225
R442 B.n88 B.t8 111.311
R443 B.n36 B.t10 111.311
R444 B.n94 B.t5 111.303
R445 B.n29 B.t1 111.303
R446 B.n191 B.n94 59.5399
R447 B.n205 B.n88 59.5399
R448 B.n356 B.n36 59.5399
R449 B.n30 B.n29 59.5399
R450 B.n94 B.n93 40.9217
R451 B.n88 B.n87 40.9217
R452 B.n36 B.n35 40.9217
R453 B.n29 B.n28 40.9217
R454 B.n415 B.n12 32.3127
R455 B.n313 B.n312 32.3127
R456 B.n248 B.n71 32.3127
R457 B.n148 B.n109 32.3127
R458 B B.n445 18.0485
R459 B.n416 B.n415 10.6151
R460 B.n417 B.n416 10.6151
R461 B.n417 B.n10 10.6151
R462 B.n421 B.n10 10.6151
R463 B.n422 B.n421 10.6151
R464 B.n423 B.n422 10.6151
R465 B.n423 B.n8 10.6151
R466 B.n427 B.n8 10.6151
R467 B.n428 B.n427 10.6151
R468 B.n429 B.n428 10.6151
R469 B.n429 B.n6 10.6151
R470 B.n433 B.n6 10.6151
R471 B.n434 B.n433 10.6151
R472 B.n435 B.n434 10.6151
R473 B.n435 B.n4 10.6151
R474 B.n439 B.n4 10.6151
R475 B.n440 B.n439 10.6151
R476 B.n441 B.n440 10.6151
R477 B.n441 B.n0 10.6151
R478 B.n411 B.n12 10.6151
R479 B.n411 B.n410 10.6151
R480 B.n410 B.n409 10.6151
R481 B.n409 B.n14 10.6151
R482 B.n405 B.n14 10.6151
R483 B.n405 B.n404 10.6151
R484 B.n404 B.n403 10.6151
R485 B.n403 B.n16 10.6151
R486 B.n399 B.n16 10.6151
R487 B.n399 B.n398 10.6151
R488 B.n398 B.n397 10.6151
R489 B.n397 B.n18 10.6151
R490 B.n393 B.n18 10.6151
R491 B.n393 B.n392 10.6151
R492 B.n392 B.n391 10.6151
R493 B.n391 B.n20 10.6151
R494 B.n387 B.n20 10.6151
R495 B.n387 B.n386 10.6151
R496 B.n386 B.n385 10.6151
R497 B.n385 B.n22 10.6151
R498 B.n381 B.n22 10.6151
R499 B.n381 B.n380 10.6151
R500 B.n380 B.n379 10.6151
R501 B.n379 B.n24 10.6151
R502 B.n375 B.n24 10.6151
R503 B.n375 B.n374 10.6151
R504 B.n374 B.n373 10.6151
R505 B.n373 B.n26 10.6151
R506 B.n369 B.n368 10.6151
R507 B.n368 B.n367 10.6151
R508 B.n367 B.n31 10.6151
R509 B.n363 B.n31 10.6151
R510 B.n363 B.n362 10.6151
R511 B.n362 B.n361 10.6151
R512 B.n361 B.n33 10.6151
R513 B.n357 B.n33 10.6151
R514 B.n355 B.n354 10.6151
R515 B.n354 B.n37 10.6151
R516 B.n350 B.n37 10.6151
R517 B.n350 B.n349 10.6151
R518 B.n349 B.n348 10.6151
R519 B.n348 B.n39 10.6151
R520 B.n344 B.n39 10.6151
R521 B.n344 B.n343 10.6151
R522 B.n343 B.n342 10.6151
R523 B.n342 B.n41 10.6151
R524 B.n338 B.n41 10.6151
R525 B.n338 B.n337 10.6151
R526 B.n337 B.n336 10.6151
R527 B.n336 B.n43 10.6151
R528 B.n332 B.n43 10.6151
R529 B.n332 B.n331 10.6151
R530 B.n331 B.n330 10.6151
R531 B.n330 B.n45 10.6151
R532 B.n326 B.n45 10.6151
R533 B.n326 B.n325 10.6151
R534 B.n325 B.n324 10.6151
R535 B.n324 B.n47 10.6151
R536 B.n320 B.n47 10.6151
R537 B.n320 B.n319 10.6151
R538 B.n319 B.n318 10.6151
R539 B.n318 B.n49 10.6151
R540 B.n314 B.n49 10.6151
R541 B.n314 B.n313 10.6151
R542 B.n312 B.n51 10.6151
R543 B.n308 B.n51 10.6151
R544 B.n308 B.n307 10.6151
R545 B.n307 B.n306 10.6151
R546 B.n306 B.n53 10.6151
R547 B.n302 B.n53 10.6151
R548 B.n302 B.n301 10.6151
R549 B.n301 B.n300 10.6151
R550 B.n300 B.n55 10.6151
R551 B.n296 B.n55 10.6151
R552 B.n296 B.n295 10.6151
R553 B.n295 B.n294 10.6151
R554 B.n294 B.n57 10.6151
R555 B.n290 B.n57 10.6151
R556 B.n290 B.n289 10.6151
R557 B.n289 B.n288 10.6151
R558 B.n288 B.n59 10.6151
R559 B.n284 B.n59 10.6151
R560 B.n284 B.n283 10.6151
R561 B.n283 B.n282 10.6151
R562 B.n282 B.n61 10.6151
R563 B.n278 B.n61 10.6151
R564 B.n278 B.n277 10.6151
R565 B.n277 B.n276 10.6151
R566 B.n276 B.n63 10.6151
R567 B.n272 B.n63 10.6151
R568 B.n272 B.n271 10.6151
R569 B.n271 B.n270 10.6151
R570 B.n270 B.n65 10.6151
R571 B.n266 B.n65 10.6151
R572 B.n266 B.n265 10.6151
R573 B.n265 B.n264 10.6151
R574 B.n264 B.n67 10.6151
R575 B.n260 B.n67 10.6151
R576 B.n260 B.n259 10.6151
R577 B.n259 B.n258 10.6151
R578 B.n258 B.n69 10.6151
R579 B.n254 B.n69 10.6151
R580 B.n254 B.n253 10.6151
R581 B.n253 B.n252 10.6151
R582 B.n252 B.n71 10.6151
R583 B.n119 B.n1 10.6151
R584 B.n120 B.n119 10.6151
R585 B.n120 B.n117 10.6151
R586 B.n124 B.n117 10.6151
R587 B.n125 B.n124 10.6151
R588 B.n126 B.n125 10.6151
R589 B.n126 B.n115 10.6151
R590 B.n130 B.n115 10.6151
R591 B.n131 B.n130 10.6151
R592 B.n132 B.n131 10.6151
R593 B.n132 B.n113 10.6151
R594 B.n136 B.n113 10.6151
R595 B.n137 B.n136 10.6151
R596 B.n138 B.n137 10.6151
R597 B.n138 B.n111 10.6151
R598 B.n142 B.n111 10.6151
R599 B.n143 B.n142 10.6151
R600 B.n144 B.n143 10.6151
R601 B.n144 B.n109 10.6151
R602 B.n149 B.n148 10.6151
R603 B.n150 B.n149 10.6151
R604 B.n150 B.n107 10.6151
R605 B.n154 B.n107 10.6151
R606 B.n155 B.n154 10.6151
R607 B.n156 B.n155 10.6151
R608 B.n156 B.n105 10.6151
R609 B.n160 B.n105 10.6151
R610 B.n161 B.n160 10.6151
R611 B.n162 B.n161 10.6151
R612 B.n162 B.n103 10.6151
R613 B.n166 B.n103 10.6151
R614 B.n167 B.n166 10.6151
R615 B.n168 B.n167 10.6151
R616 B.n168 B.n101 10.6151
R617 B.n172 B.n101 10.6151
R618 B.n173 B.n172 10.6151
R619 B.n174 B.n173 10.6151
R620 B.n174 B.n99 10.6151
R621 B.n178 B.n99 10.6151
R622 B.n179 B.n178 10.6151
R623 B.n180 B.n179 10.6151
R624 B.n180 B.n97 10.6151
R625 B.n184 B.n97 10.6151
R626 B.n185 B.n184 10.6151
R627 B.n186 B.n185 10.6151
R628 B.n186 B.n95 10.6151
R629 B.n190 B.n95 10.6151
R630 B.n193 B.n192 10.6151
R631 B.n193 B.n91 10.6151
R632 B.n197 B.n91 10.6151
R633 B.n198 B.n197 10.6151
R634 B.n199 B.n198 10.6151
R635 B.n199 B.n89 10.6151
R636 B.n203 B.n89 10.6151
R637 B.n204 B.n203 10.6151
R638 B.n206 B.n85 10.6151
R639 B.n210 B.n85 10.6151
R640 B.n211 B.n210 10.6151
R641 B.n212 B.n211 10.6151
R642 B.n212 B.n83 10.6151
R643 B.n216 B.n83 10.6151
R644 B.n217 B.n216 10.6151
R645 B.n218 B.n217 10.6151
R646 B.n218 B.n81 10.6151
R647 B.n222 B.n81 10.6151
R648 B.n223 B.n222 10.6151
R649 B.n224 B.n223 10.6151
R650 B.n224 B.n79 10.6151
R651 B.n228 B.n79 10.6151
R652 B.n229 B.n228 10.6151
R653 B.n230 B.n229 10.6151
R654 B.n230 B.n77 10.6151
R655 B.n234 B.n77 10.6151
R656 B.n235 B.n234 10.6151
R657 B.n236 B.n235 10.6151
R658 B.n236 B.n75 10.6151
R659 B.n240 B.n75 10.6151
R660 B.n241 B.n240 10.6151
R661 B.n242 B.n241 10.6151
R662 B.n242 B.n73 10.6151
R663 B.n246 B.n73 10.6151
R664 B.n247 B.n246 10.6151
R665 B.n248 B.n247 10.6151
R666 B.n445 B.n0 8.11757
R667 B.n445 B.n1 8.11757
R668 B.n369 B.n30 6.5566
R669 B.n357 B.n356 6.5566
R670 B.n192 B.n191 6.5566
R671 B.n205 B.n204 6.5566
R672 B.n30 B.n26 4.05904
R673 B.n356 B.n355 4.05904
R674 B.n191 B.n190 4.05904
R675 B.n206 B.n205 4.05904
R676 VP.n0 VP.t0 200.934
R677 VP.n0 VP.t1 161.786
R678 VP VP.n0 0.241678
R679 VTAIL.n1 VTAIL.t1 74.2414
R680 VTAIL.n3 VTAIL.t0 74.2412
R681 VTAIL.n0 VTAIL.t3 74.2412
R682 VTAIL.n2 VTAIL.t2 74.2412
R683 VTAIL.n1 VTAIL.n0 22.5565
R684 VTAIL.n3 VTAIL.n2 20.7376
R685 VTAIL.n2 VTAIL.n1 1.37981
R686 VTAIL VTAIL.n0 0.983259
R687 VTAIL VTAIL.n3 0.397052
R688 VDD1 VDD1.t0 125.749
R689 VDD1 VDD1.t1 91.4329
R690 VN VN.t0 201.125
R691 VN VN.t1 162.026
R692 VDD2.n0 VDD2.t0 124.769
R693 VDD2.n0 VDD2.t1 90.92
R694 VDD2 VDD2.n0 0.513431
C0 B VN 0.862729f
C1 VN w_n1814_n2488# 2.35406f
C2 VN VDD2 1.73285f
C3 VTAIL VN 1.53315f
C4 VN VP 4.2547f
C5 VN VDD1 0.14808f
C6 B w_n1814_n2488# 6.68944f
C7 B VDD2 1.27425f
C8 w_n1814_n2488# VDD2 1.39417f
C9 B VTAIL 2.37781f
C10 VTAIL w_n1814_n2488# 2.13038f
C11 VTAIL VDD2 3.81681f
C12 B VP 1.23642f
C13 VP w_n1814_n2488# 2.58336f
C14 B VDD1 1.25142f
C15 VP VDD2 0.29858f
C16 w_n1814_n2488# VDD1 1.37815f
C17 VDD1 VDD2 0.577199f
C18 VTAIL VP 1.54742f
C19 VTAIL VDD1 3.77141f
C20 VP VDD1 1.88129f
C21 VDD2 VSUBS 0.65421f
C22 VDD1 VSUBS 2.765716f
C23 VTAIL VSUBS 0.71908f
C24 VN VSUBS 5.22825f
C25 VP VSUBS 1.264384f
C26 B VSUBS 2.914437f
C27 w_n1814_n2488# VSUBS 56.0526f
C28 VDD2.t0 VSUBS 1.04808f
C29 VDD2.t1 VSUBS 0.801311f
C30 VDD2.n0 VSUBS 1.88572f
C31 VN.t1 VSUBS 1.52098f
C32 VN.t0 VSUBS 1.87337f
C33 VDD1.t1 VSUBS 0.792148f
C34 VDD1.t0 VSUBS 1.05027f
C35 VTAIL.t3 VSUBS 1.29939f
C36 VTAIL.n0 VSUBS 1.76638f
C37 VTAIL.t1 VSUBS 1.29939f
C38 VTAIL.n1 VSUBS 1.79789f
C39 VTAIL.t2 VSUBS 1.29939f
C40 VTAIL.n2 VSUBS 1.65333f
C41 VTAIL.t0 VSUBS 1.29939f
C42 VTAIL.n3 VSUBS 1.57522f
C43 VP.t0 VSUBS 1.93889f
C44 VP.t1 VSUBS 1.5773f
C45 VP.n0 VSUBS 3.3286f
C46 B.n0 VSUBS 0.006663f
C47 B.n1 VSUBS 0.006663f
C48 B.n2 VSUBS 0.009854f
C49 B.n3 VSUBS 0.007551f
C50 B.n4 VSUBS 0.007551f
C51 B.n5 VSUBS 0.007551f
C52 B.n6 VSUBS 0.007551f
C53 B.n7 VSUBS 0.007551f
C54 B.n8 VSUBS 0.007551f
C55 B.n9 VSUBS 0.007551f
C56 B.n10 VSUBS 0.007551f
C57 B.n11 VSUBS 0.007551f
C58 B.n12 VSUBS 0.018018f
C59 B.n13 VSUBS 0.007551f
C60 B.n14 VSUBS 0.007551f
C61 B.n15 VSUBS 0.007551f
C62 B.n16 VSUBS 0.007551f
C63 B.n17 VSUBS 0.007551f
C64 B.n18 VSUBS 0.007551f
C65 B.n19 VSUBS 0.007551f
C66 B.n20 VSUBS 0.007551f
C67 B.n21 VSUBS 0.007551f
C68 B.n22 VSUBS 0.007551f
C69 B.n23 VSUBS 0.007551f
C70 B.n24 VSUBS 0.007551f
C71 B.n25 VSUBS 0.007551f
C72 B.n26 VSUBS 0.005219f
C73 B.n27 VSUBS 0.007551f
C74 B.t1 VSUBS 0.250778f
C75 B.t2 VSUBS 0.267574f
C76 B.t0 VSUBS 0.666446f
C77 B.n28 VSUBS 0.136794f
C78 B.n29 VSUBS 0.073252f
C79 B.n30 VSUBS 0.017495f
C80 B.n31 VSUBS 0.007551f
C81 B.n32 VSUBS 0.007551f
C82 B.n33 VSUBS 0.007551f
C83 B.n34 VSUBS 0.007551f
C84 B.t10 VSUBS 0.250776f
C85 B.t11 VSUBS 0.267572f
C86 B.t9 VSUBS 0.666446f
C87 B.n35 VSUBS 0.136796f
C88 B.n36 VSUBS 0.073254f
C89 B.n37 VSUBS 0.007551f
C90 B.n38 VSUBS 0.007551f
C91 B.n39 VSUBS 0.007551f
C92 B.n40 VSUBS 0.007551f
C93 B.n41 VSUBS 0.007551f
C94 B.n42 VSUBS 0.007551f
C95 B.n43 VSUBS 0.007551f
C96 B.n44 VSUBS 0.007551f
C97 B.n45 VSUBS 0.007551f
C98 B.n46 VSUBS 0.007551f
C99 B.n47 VSUBS 0.007551f
C100 B.n48 VSUBS 0.007551f
C101 B.n49 VSUBS 0.007551f
C102 B.n50 VSUBS 0.018018f
C103 B.n51 VSUBS 0.007551f
C104 B.n52 VSUBS 0.007551f
C105 B.n53 VSUBS 0.007551f
C106 B.n54 VSUBS 0.007551f
C107 B.n55 VSUBS 0.007551f
C108 B.n56 VSUBS 0.007551f
C109 B.n57 VSUBS 0.007551f
C110 B.n58 VSUBS 0.007551f
C111 B.n59 VSUBS 0.007551f
C112 B.n60 VSUBS 0.007551f
C113 B.n61 VSUBS 0.007551f
C114 B.n62 VSUBS 0.007551f
C115 B.n63 VSUBS 0.007551f
C116 B.n64 VSUBS 0.007551f
C117 B.n65 VSUBS 0.007551f
C118 B.n66 VSUBS 0.007551f
C119 B.n67 VSUBS 0.007551f
C120 B.n68 VSUBS 0.007551f
C121 B.n69 VSUBS 0.007551f
C122 B.n70 VSUBS 0.007551f
C123 B.n71 VSUBS 0.017974f
C124 B.n72 VSUBS 0.007551f
C125 B.n73 VSUBS 0.007551f
C126 B.n74 VSUBS 0.007551f
C127 B.n75 VSUBS 0.007551f
C128 B.n76 VSUBS 0.007551f
C129 B.n77 VSUBS 0.007551f
C130 B.n78 VSUBS 0.007551f
C131 B.n79 VSUBS 0.007551f
C132 B.n80 VSUBS 0.007551f
C133 B.n81 VSUBS 0.007551f
C134 B.n82 VSUBS 0.007551f
C135 B.n83 VSUBS 0.007551f
C136 B.n84 VSUBS 0.007551f
C137 B.n85 VSUBS 0.007551f
C138 B.n86 VSUBS 0.007551f
C139 B.t8 VSUBS 0.250776f
C140 B.t7 VSUBS 0.267572f
C141 B.t6 VSUBS 0.666446f
C142 B.n87 VSUBS 0.136796f
C143 B.n88 VSUBS 0.073254f
C144 B.n89 VSUBS 0.007551f
C145 B.n90 VSUBS 0.007551f
C146 B.n91 VSUBS 0.007551f
C147 B.n92 VSUBS 0.007551f
C148 B.t5 VSUBS 0.250778f
C149 B.t4 VSUBS 0.267574f
C150 B.t3 VSUBS 0.666446f
C151 B.n93 VSUBS 0.136794f
C152 B.n94 VSUBS 0.073252f
C153 B.n95 VSUBS 0.007551f
C154 B.n96 VSUBS 0.007551f
C155 B.n97 VSUBS 0.007551f
C156 B.n98 VSUBS 0.007551f
C157 B.n99 VSUBS 0.007551f
C158 B.n100 VSUBS 0.007551f
C159 B.n101 VSUBS 0.007551f
C160 B.n102 VSUBS 0.007551f
C161 B.n103 VSUBS 0.007551f
C162 B.n104 VSUBS 0.007551f
C163 B.n105 VSUBS 0.007551f
C164 B.n106 VSUBS 0.007551f
C165 B.n107 VSUBS 0.007551f
C166 B.n108 VSUBS 0.007551f
C167 B.n109 VSUBS 0.017072f
C168 B.n110 VSUBS 0.007551f
C169 B.n111 VSUBS 0.007551f
C170 B.n112 VSUBS 0.007551f
C171 B.n113 VSUBS 0.007551f
C172 B.n114 VSUBS 0.007551f
C173 B.n115 VSUBS 0.007551f
C174 B.n116 VSUBS 0.007551f
C175 B.n117 VSUBS 0.007551f
C176 B.n118 VSUBS 0.007551f
C177 B.n119 VSUBS 0.007551f
C178 B.n120 VSUBS 0.007551f
C179 B.n121 VSUBS 0.007551f
C180 B.n122 VSUBS 0.007551f
C181 B.n123 VSUBS 0.007551f
C182 B.n124 VSUBS 0.007551f
C183 B.n125 VSUBS 0.007551f
C184 B.n126 VSUBS 0.007551f
C185 B.n127 VSUBS 0.007551f
C186 B.n128 VSUBS 0.007551f
C187 B.n129 VSUBS 0.007551f
C188 B.n130 VSUBS 0.007551f
C189 B.n131 VSUBS 0.007551f
C190 B.n132 VSUBS 0.007551f
C191 B.n133 VSUBS 0.007551f
C192 B.n134 VSUBS 0.007551f
C193 B.n135 VSUBS 0.007551f
C194 B.n136 VSUBS 0.007551f
C195 B.n137 VSUBS 0.007551f
C196 B.n138 VSUBS 0.007551f
C197 B.n139 VSUBS 0.007551f
C198 B.n140 VSUBS 0.007551f
C199 B.n141 VSUBS 0.007551f
C200 B.n142 VSUBS 0.007551f
C201 B.n143 VSUBS 0.007551f
C202 B.n144 VSUBS 0.007551f
C203 B.n145 VSUBS 0.007551f
C204 B.n146 VSUBS 0.017072f
C205 B.n147 VSUBS 0.018018f
C206 B.n148 VSUBS 0.018018f
C207 B.n149 VSUBS 0.007551f
C208 B.n150 VSUBS 0.007551f
C209 B.n151 VSUBS 0.007551f
C210 B.n152 VSUBS 0.007551f
C211 B.n153 VSUBS 0.007551f
C212 B.n154 VSUBS 0.007551f
C213 B.n155 VSUBS 0.007551f
C214 B.n156 VSUBS 0.007551f
C215 B.n157 VSUBS 0.007551f
C216 B.n158 VSUBS 0.007551f
C217 B.n159 VSUBS 0.007551f
C218 B.n160 VSUBS 0.007551f
C219 B.n161 VSUBS 0.007551f
C220 B.n162 VSUBS 0.007551f
C221 B.n163 VSUBS 0.007551f
C222 B.n164 VSUBS 0.007551f
C223 B.n165 VSUBS 0.007551f
C224 B.n166 VSUBS 0.007551f
C225 B.n167 VSUBS 0.007551f
C226 B.n168 VSUBS 0.007551f
C227 B.n169 VSUBS 0.007551f
C228 B.n170 VSUBS 0.007551f
C229 B.n171 VSUBS 0.007551f
C230 B.n172 VSUBS 0.007551f
C231 B.n173 VSUBS 0.007551f
C232 B.n174 VSUBS 0.007551f
C233 B.n175 VSUBS 0.007551f
C234 B.n176 VSUBS 0.007551f
C235 B.n177 VSUBS 0.007551f
C236 B.n178 VSUBS 0.007551f
C237 B.n179 VSUBS 0.007551f
C238 B.n180 VSUBS 0.007551f
C239 B.n181 VSUBS 0.007551f
C240 B.n182 VSUBS 0.007551f
C241 B.n183 VSUBS 0.007551f
C242 B.n184 VSUBS 0.007551f
C243 B.n185 VSUBS 0.007551f
C244 B.n186 VSUBS 0.007551f
C245 B.n187 VSUBS 0.007551f
C246 B.n188 VSUBS 0.007551f
C247 B.n189 VSUBS 0.007551f
C248 B.n190 VSUBS 0.005219f
C249 B.n191 VSUBS 0.017495f
C250 B.n192 VSUBS 0.006108f
C251 B.n193 VSUBS 0.007551f
C252 B.n194 VSUBS 0.007551f
C253 B.n195 VSUBS 0.007551f
C254 B.n196 VSUBS 0.007551f
C255 B.n197 VSUBS 0.007551f
C256 B.n198 VSUBS 0.007551f
C257 B.n199 VSUBS 0.007551f
C258 B.n200 VSUBS 0.007551f
C259 B.n201 VSUBS 0.007551f
C260 B.n202 VSUBS 0.007551f
C261 B.n203 VSUBS 0.007551f
C262 B.n204 VSUBS 0.006108f
C263 B.n205 VSUBS 0.017495f
C264 B.n206 VSUBS 0.005219f
C265 B.n207 VSUBS 0.007551f
C266 B.n208 VSUBS 0.007551f
C267 B.n209 VSUBS 0.007551f
C268 B.n210 VSUBS 0.007551f
C269 B.n211 VSUBS 0.007551f
C270 B.n212 VSUBS 0.007551f
C271 B.n213 VSUBS 0.007551f
C272 B.n214 VSUBS 0.007551f
C273 B.n215 VSUBS 0.007551f
C274 B.n216 VSUBS 0.007551f
C275 B.n217 VSUBS 0.007551f
C276 B.n218 VSUBS 0.007551f
C277 B.n219 VSUBS 0.007551f
C278 B.n220 VSUBS 0.007551f
C279 B.n221 VSUBS 0.007551f
C280 B.n222 VSUBS 0.007551f
C281 B.n223 VSUBS 0.007551f
C282 B.n224 VSUBS 0.007551f
C283 B.n225 VSUBS 0.007551f
C284 B.n226 VSUBS 0.007551f
C285 B.n227 VSUBS 0.007551f
C286 B.n228 VSUBS 0.007551f
C287 B.n229 VSUBS 0.007551f
C288 B.n230 VSUBS 0.007551f
C289 B.n231 VSUBS 0.007551f
C290 B.n232 VSUBS 0.007551f
C291 B.n233 VSUBS 0.007551f
C292 B.n234 VSUBS 0.007551f
C293 B.n235 VSUBS 0.007551f
C294 B.n236 VSUBS 0.007551f
C295 B.n237 VSUBS 0.007551f
C296 B.n238 VSUBS 0.007551f
C297 B.n239 VSUBS 0.007551f
C298 B.n240 VSUBS 0.007551f
C299 B.n241 VSUBS 0.007551f
C300 B.n242 VSUBS 0.007551f
C301 B.n243 VSUBS 0.007551f
C302 B.n244 VSUBS 0.007551f
C303 B.n245 VSUBS 0.007551f
C304 B.n246 VSUBS 0.007551f
C305 B.n247 VSUBS 0.007551f
C306 B.n248 VSUBS 0.017116f
C307 B.n249 VSUBS 0.018018f
C308 B.n250 VSUBS 0.017072f
C309 B.n251 VSUBS 0.007551f
C310 B.n252 VSUBS 0.007551f
C311 B.n253 VSUBS 0.007551f
C312 B.n254 VSUBS 0.007551f
C313 B.n255 VSUBS 0.007551f
C314 B.n256 VSUBS 0.007551f
C315 B.n257 VSUBS 0.007551f
C316 B.n258 VSUBS 0.007551f
C317 B.n259 VSUBS 0.007551f
C318 B.n260 VSUBS 0.007551f
C319 B.n261 VSUBS 0.007551f
C320 B.n262 VSUBS 0.007551f
C321 B.n263 VSUBS 0.007551f
C322 B.n264 VSUBS 0.007551f
C323 B.n265 VSUBS 0.007551f
C324 B.n266 VSUBS 0.007551f
C325 B.n267 VSUBS 0.007551f
C326 B.n268 VSUBS 0.007551f
C327 B.n269 VSUBS 0.007551f
C328 B.n270 VSUBS 0.007551f
C329 B.n271 VSUBS 0.007551f
C330 B.n272 VSUBS 0.007551f
C331 B.n273 VSUBS 0.007551f
C332 B.n274 VSUBS 0.007551f
C333 B.n275 VSUBS 0.007551f
C334 B.n276 VSUBS 0.007551f
C335 B.n277 VSUBS 0.007551f
C336 B.n278 VSUBS 0.007551f
C337 B.n279 VSUBS 0.007551f
C338 B.n280 VSUBS 0.007551f
C339 B.n281 VSUBS 0.007551f
C340 B.n282 VSUBS 0.007551f
C341 B.n283 VSUBS 0.007551f
C342 B.n284 VSUBS 0.007551f
C343 B.n285 VSUBS 0.007551f
C344 B.n286 VSUBS 0.007551f
C345 B.n287 VSUBS 0.007551f
C346 B.n288 VSUBS 0.007551f
C347 B.n289 VSUBS 0.007551f
C348 B.n290 VSUBS 0.007551f
C349 B.n291 VSUBS 0.007551f
C350 B.n292 VSUBS 0.007551f
C351 B.n293 VSUBS 0.007551f
C352 B.n294 VSUBS 0.007551f
C353 B.n295 VSUBS 0.007551f
C354 B.n296 VSUBS 0.007551f
C355 B.n297 VSUBS 0.007551f
C356 B.n298 VSUBS 0.007551f
C357 B.n299 VSUBS 0.007551f
C358 B.n300 VSUBS 0.007551f
C359 B.n301 VSUBS 0.007551f
C360 B.n302 VSUBS 0.007551f
C361 B.n303 VSUBS 0.007551f
C362 B.n304 VSUBS 0.007551f
C363 B.n305 VSUBS 0.007551f
C364 B.n306 VSUBS 0.007551f
C365 B.n307 VSUBS 0.007551f
C366 B.n308 VSUBS 0.007551f
C367 B.n309 VSUBS 0.007551f
C368 B.n310 VSUBS 0.007551f
C369 B.n311 VSUBS 0.017072f
C370 B.n312 VSUBS 0.017072f
C371 B.n313 VSUBS 0.018018f
C372 B.n314 VSUBS 0.007551f
C373 B.n315 VSUBS 0.007551f
C374 B.n316 VSUBS 0.007551f
C375 B.n317 VSUBS 0.007551f
C376 B.n318 VSUBS 0.007551f
C377 B.n319 VSUBS 0.007551f
C378 B.n320 VSUBS 0.007551f
C379 B.n321 VSUBS 0.007551f
C380 B.n322 VSUBS 0.007551f
C381 B.n323 VSUBS 0.007551f
C382 B.n324 VSUBS 0.007551f
C383 B.n325 VSUBS 0.007551f
C384 B.n326 VSUBS 0.007551f
C385 B.n327 VSUBS 0.007551f
C386 B.n328 VSUBS 0.007551f
C387 B.n329 VSUBS 0.007551f
C388 B.n330 VSUBS 0.007551f
C389 B.n331 VSUBS 0.007551f
C390 B.n332 VSUBS 0.007551f
C391 B.n333 VSUBS 0.007551f
C392 B.n334 VSUBS 0.007551f
C393 B.n335 VSUBS 0.007551f
C394 B.n336 VSUBS 0.007551f
C395 B.n337 VSUBS 0.007551f
C396 B.n338 VSUBS 0.007551f
C397 B.n339 VSUBS 0.007551f
C398 B.n340 VSUBS 0.007551f
C399 B.n341 VSUBS 0.007551f
C400 B.n342 VSUBS 0.007551f
C401 B.n343 VSUBS 0.007551f
C402 B.n344 VSUBS 0.007551f
C403 B.n345 VSUBS 0.007551f
C404 B.n346 VSUBS 0.007551f
C405 B.n347 VSUBS 0.007551f
C406 B.n348 VSUBS 0.007551f
C407 B.n349 VSUBS 0.007551f
C408 B.n350 VSUBS 0.007551f
C409 B.n351 VSUBS 0.007551f
C410 B.n352 VSUBS 0.007551f
C411 B.n353 VSUBS 0.007551f
C412 B.n354 VSUBS 0.007551f
C413 B.n355 VSUBS 0.005219f
C414 B.n356 VSUBS 0.017495f
C415 B.n357 VSUBS 0.006108f
C416 B.n358 VSUBS 0.007551f
C417 B.n359 VSUBS 0.007551f
C418 B.n360 VSUBS 0.007551f
C419 B.n361 VSUBS 0.007551f
C420 B.n362 VSUBS 0.007551f
C421 B.n363 VSUBS 0.007551f
C422 B.n364 VSUBS 0.007551f
C423 B.n365 VSUBS 0.007551f
C424 B.n366 VSUBS 0.007551f
C425 B.n367 VSUBS 0.007551f
C426 B.n368 VSUBS 0.007551f
C427 B.n369 VSUBS 0.006108f
C428 B.n370 VSUBS 0.007551f
C429 B.n371 VSUBS 0.007551f
C430 B.n372 VSUBS 0.007551f
C431 B.n373 VSUBS 0.007551f
C432 B.n374 VSUBS 0.007551f
C433 B.n375 VSUBS 0.007551f
C434 B.n376 VSUBS 0.007551f
C435 B.n377 VSUBS 0.007551f
C436 B.n378 VSUBS 0.007551f
C437 B.n379 VSUBS 0.007551f
C438 B.n380 VSUBS 0.007551f
C439 B.n381 VSUBS 0.007551f
C440 B.n382 VSUBS 0.007551f
C441 B.n383 VSUBS 0.007551f
C442 B.n384 VSUBS 0.007551f
C443 B.n385 VSUBS 0.007551f
C444 B.n386 VSUBS 0.007551f
C445 B.n387 VSUBS 0.007551f
C446 B.n388 VSUBS 0.007551f
C447 B.n389 VSUBS 0.007551f
C448 B.n390 VSUBS 0.007551f
C449 B.n391 VSUBS 0.007551f
C450 B.n392 VSUBS 0.007551f
C451 B.n393 VSUBS 0.007551f
C452 B.n394 VSUBS 0.007551f
C453 B.n395 VSUBS 0.007551f
C454 B.n396 VSUBS 0.007551f
C455 B.n397 VSUBS 0.007551f
C456 B.n398 VSUBS 0.007551f
C457 B.n399 VSUBS 0.007551f
C458 B.n400 VSUBS 0.007551f
C459 B.n401 VSUBS 0.007551f
C460 B.n402 VSUBS 0.007551f
C461 B.n403 VSUBS 0.007551f
C462 B.n404 VSUBS 0.007551f
C463 B.n405 VSUBS 0.007551f
C464 B.n406 VSUBS 0.007551f
C465 B.n407 VSUBS 0.007551f
C466 B.n408 VSUBS 0.007551f
C467 B.n409 VSUBS 0.007551f
C468 B.n410 VSUBS 0.007551f
C469 B.n411 VSUBS 0.007551f
C470 B.n412 VSUBS 0.007551f
C471 B.n413 VSUBS 0.018018f
C472 B.n414 VSUBS 0.017072f
C473 B.n415 VSUBS 0.017072f
C474 B.n416 VSUBS 0.007551f
C475 B.n417 VSUBS 0.007551f
C476 B.n418 VSUBS 0.007551f
C477 B.n419 VSUBS 0.007551f
C478 B.n420 VSUBS 0.007551f
C479 B.n421 VSUBS 0.007551f
C480 B.n422 VSUBS 0.007551f
C481 B.n423 VSUBS 0.007551f
C482 B.n424 VSUBS 0.007551f
C483 B.n425 VSUBS 0.007551f
C484 B.n426 VSUBS 0.007551f
C485 B.n427 VSUBS 0.007551f
C486 B.n428 VSUBS 0.007551f
C487 B.n429 VSUBS 0.007551f
C488 B.n430 VSUBS 0.007551f
C489 B.n431 VSUBS 0.007551f
C490 B.n432 VSUBS 0.007551f
C491 B.n433 VSUBS 0.007551f
C492 B.n434 VSUBS 0.007551f
C493 B.n435 VSUBS 0.007551f
C494 B.n436 VSUBS 0.007551f
C495 B.n437 VSUBS 0.007551f
C496 B.n438 VSUBS 0.007551f
C497 B.n439 VSUBS 0.007551f
C498 B.n440 VSUBS 0.007551f
C499 B.n441 VSUBS 0.007551f
C500 B.n442 VSUBS 0.007551f
C501 B.n443 VSUBS 0.009854f
C502 B.n444 VSUBS 0.010497f
C503 B.n445 VSUBS 0.020874f
.ends

