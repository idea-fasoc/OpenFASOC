* NGSPICE file created from diff_pair_sample_0704.ext - technology: sky130A

.subckt diff_pair_sample_0704 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t14 w_n5100_n3794# sky130_fd_pr__pfet_01v8 ad=2.33145 pd=14.46 as=2.33145 ps=14.46 w=14.13 l=3.8
X1 VTAIL.t3 VN.t0 VDD2.t7 w_n5100_n3794# sky130_fd_pr__pfet_01v8 ad=2.33145 pd=14.46 as=2.33145 ps=14.46 w=14.13 l=3.8
X2 B.t11 B.t9 B.t10 w_n5100_n3794# sky130_fd_pr__pfet_01v8 ad=5.5107 pd=29.04 as=0 ps=0 w=14.13 l=3.8
X3 B.t8 B.t6 B.t7 w_n5100_n3794# sky130_fd_pr__pfet_01v8 ad=5.5107 pd=29.04 as=0 ps=0 w=14.13 l=3.8
X4 VDD2.t6 VN.t1 VTAIL.t7 w_n5100_n3794# sky130_fd_pr__pfet_01v8 ad=2.33145 pd=14.46 as=5.5107 ps=29.04 w=14.13 l=3.8
X5 B.t5 B.t3 B.t4 w_n5100_n3794# sky130_fd_pr__pfet_01v8 ad=5.5107 pd=29.04 as=0 ps=0 w=14.13 l=3.8
X6 VDD2.t5 VN.t2 VTAIL.t2 w_n5100_n3794# sky130_fd_pr__pfet_01v8 ad=2.33145 pd=14.46 as=2.33145 ps=14.46 w=14.13 l=3.8
X7 VTAIL.t9 VP.t1 VDD1.t6 w_n5100_n3794# sky130_fd_pr__pfet_01v8 ad=5.5107 pd=29.04 as=2.33145 ps=14.46 w=14.13 l=3.8
X8 VTAIL.t5 VN.t3 VDD2.t4 w_n5100_n3794# sky130_fd_pr__pfet_01v8 ad=5.5107 pd=29.04 as=2.33145 ps=14.46 w=14.13 l=3.8
X9 VDD1.t5 VP.t2 VTAIL.t8 w_n5100_n3794# sky130_fd_pr__pfet_01v8 ad=2.33145 pd=14.46 as=2.33145 ps=14.46 w=14.13 l=3.8
X10 VTAIL.t0 VN.t4 VDD2.t3 w_n5100_n3794# sky130_fd_pr__pfet_01v8 ad=2.33145 pd=14.46 as=2.33145 ps=14.46 w=14.13 l=3.8
X11 VDD2.t2 VN.t5 VTAIL.t4 w_n5100_n3794# sky130_fd_pr__pfet_01v8 ad=2.33145 pd=14.46 as=2.33145 ps=14.46 w=14.13 l=3.8
X12 VDD1.t4 VP.t3 VTAIL.t13 w_n5100_n3794# sky130_fd_pr__pfet_01v8 ad=2.33145 pd=14.46 as=5.5107 ps=29.04 w=14.13 l=3.8
X13 B.t2 B.t0 B.t1 w_n5100_n3794# sky130_fd_pr__pfet_01v8 ad=5.5107 pd=29.04 as=0 ps=0 w=14.13 l=3.8
X14 VTAIL.t15 VP.t4 VDD1.t3 w_n5100_n3794# sky130_fd_pr__pfet_01v8 ad=2.33145 pd=14.46 as=2.33145 ps=14.46 w=14.13 l=3.8
X15 VTAIL.t12 VP.t5 VDD1.t2 w_n5100_n3794# sky130_fd_pr__pfet_01v8 ad=5.5107 pd=29.04 as=2.33145 ps=14.46 w=14.13 l=3.8
X16 VTAIL.t1 VN.t6 VDD2.t1 w_n5100_n3794# sky130_fd_pr__pfet_01v8 ad=5.5107 pd=29.04 as=2.33145 ps=14.46 w=14.13 l=3.8
X17 VTAIL.t10 VP.t6 VDD1.t1 w_n5100_n3794# sky130_fd_pr__pfet_01v8 ad=2.33145 pd=14.46 as=2.33145 ps=14.46 w=14.13 l=3.8
X18 VDD2.t0 VN.t7 VTAIL.t6 w_n5100_n3794# sky130_fd_pr__pfet_01v8 ad=2.33145 pd=14.46 as=5.5107 ps=29.04 w=14.13 l=3.8
X19 VDD1.t0 VP.t7 VTAIL.t11 w_n5100_n3794# sky130_fd_pr__pfet_01v8 ad=2.33145 pd=14.46 as=5.5107 ps=29.04 w=14.13 l=3.8
R0 VP.n23 VP.n22 161.3
R1 VP.n24 VP.n19 161.3
R2 VP.n26 VP.n25 161.3
R3 VP.n27 VP.n18 161.3
R4 VP.n29 VP.n28 161.3
R5 VP.n30 VP.n17 161.3
R6 VP.n32 VP.n31 161.3
R7 VP.n33 VP.n16 161.3
R8 VP.n36 VP.n35 161.3
R9 VP.n37 VP.n15 161.3
R10 VP.n39 VP.n38 161.3
R11 VP.n40 VP.n14 161.3
R12 VP.n42 VP.n41 161.3
R13 VP.n43 VP.n13 161.3
R14 VP.n45 VP.n44 161.3
R15 VP.n46 VP.n12 161.3
R16 VP.n88 VP.n0 161.3
R17 VP.n87 VP.n86 161.3
R18 VP.n85 VP.n1 161.3
R19 VP.n84 VP.n83 161.3
R20 VP.n82 VP.n2 161.3
R21 VP.n81 VP.n80 161.3
R22 VP.n79 VP.n3 161.3
R23 VP.n78 VP.n77 161.3
R24 VP.n75 VP.n4 161.3
R25 VP.n74 VP.n73 161.3
R26 VP.n72 VP.n5 161.3
R27 VP.n71 VP.n70 161.3
R28 VP.n69 VP.n6 161.3
R29 VP.n68 VP.n67 161.3
R30 VP.n66 VP.n7 161.3
R31 VP.n65 VP.n64 161.3
R32 VP.n62 VP.n8 161.3
R33 VP.n61 VP.n60 161.3
R34 VP.n59 VP.n9 161.3
R35 VP.n58 VP.n57 161.3
R36 VP.n56 VP.n10 161.3
R37 VP.n55 VP.n54 161.3
R38 VP.n53 VP.n11 161.3
R39 VP.n52 VP.n51 161.3
R40 VP.n20 VP.t5 121.847
R41 VP.n50 VP.t1 89.6144
R42 VP.n63 VP.t2 89.6144
R43 VP.n76 VP.t6 89.6144
R44 VP.n89 VP.t7 89.6144
R45 VP.n47 VP.t3 89.6144
R46 VP.n34 VP.t4 89.6144
R47 VP.n21 VP.t0 89.6144
R48 VP.n50 VP.n49 60.4062
R49 VP.n90 VP.n89 60.4062
R50 VP.n48 VP.n47 60.4062
R51 VP.n21 VP.n20 59.6416
R52 VP.n49 VP.n48 58.3449
R53 VP.n70 VP.n69 56.5193
R54 VP.n28 VP.n27 56.5193
R55 VP.n57 VP.n56 52.1486
R56 VP.n83 VP.n82 52.1486
R57 VP.n41 VP.n40 52.1486
R58 VP.n56 VP.n55 28.8382
R59 VP.n83 VP.n1 28.8382
R60 VP.n41 VP.n13 28.8382
R61 VP.n51 VP.n11 24.4675
R62 VP.n55 VP.n11 24.4675
R63 VP.n57 VP.n9 24.4675
R64 VP.n61 VP.n9 24.4675
R65 VP.n62 VP.n61 24.4675
R66 VP.n64 VP.n7 24.4675
R67 VP.n68 VP.n7 24.4675
R68 VP.n69 VP.n68 24.4675
R69 VP.n70 VP.n5 24.4675
R70 VP.n74 VP.n5 24.4675
R71 VP.n75 VP.n74 24.4675
R72 VP.n77 VP.n3 24.4675
R73 VP.n81 VP.n3 24.4675
R74 VP.n82 VP.n81 24.4675
R75 VP.n87 VP.n1 24.4675
R76 VP.n88 VP.n87 24.4675
R77 VP.n45 VP.n13 24.4675
R78 VP.n46 VP.n45 24.4675
R79 VP.n28 VP.n17 24.4675
R80 VP.n32 VP.n17 24.4675
R81 VP.n33 VP.n32 24.4675
R82 VP.n35 VP.n15 24.4675
R83 VP.n39 VP.n15 24.4675
R84 VP.n40 VP.n39 24.4675
R85 VP.n22 VP.n19 24.4675
R86 VP.n26 VP.n19 24.4675
R87 VP.n27 VP.n26 24.4675
R88 VP.n51 VP.n50 21.7761
R89 VP.n89 VP.n88 21.7761
R90 VP.n47 VP.n46 21.7761
R91 VP.n64 VP.n63 15.4147
R92 VP.n76 VP.n75 15.4147
R93 VP.n34 VP.n33 15.4147
R94 VP.n22 VP.n21 15.4147
R95 VP.n63 VP.n62 9.05329
R96 VP.n77 VP.n76 9.05329
R97 VP.n35 VP.n34 9.05329
R98 VP.n23 VP.n20 2.62602
R99 VP.n48 VP.n12 0.417535
R100 VP.n52 VP.n49 0.417535
R101 VP.n90 VP.n0 0.417535
R102 VP VP.n90 0.394291
R103 VP.n24 VP.n23 0.189894
R104 VP.n25 VP.n24 0.189894
R105 VP.n25 VP.n18 0.189894
R106 VP.n29 VP.n18 0.189894
R107 VP.n30 VP.n29 0.189894
R108 VP.n31 VP.n30 0.189894
R109 VP.n31 VP.n16 0.189894
R110 VP.n36 VP.n16 0.189894
R111 VP.n37 VP.n36 0.189894
R112 VP.n38 VP.n37 0.189894
R113 VP.n38 VP.n14 0.189894
R114 VP.n42 VP.n14 0.189894
R115 VP.n43 VP.n42 0.189894
R116 VP.n44 VP.n43 0.189894
R117 VP.n44 VP.n12 0.189894
R118 VP.n53 VP.n52 0.189894
R119 VP.n54 VP.n53 0.189894
R120 VP.n54 VP.n10 0.189894
R121 VP.n58 VP.n10 0.189894
R122 VP.n59 VP.n58 0.189894
R123 VP.n60 VP.n59 0.189894
R124 VP.n60 VP.n8 0.189894
R125 VP.n65 VP.n8 0.189894
R126 VP.n66 VP.n65 0.189894
R127 VP.n67 VP.n66 0.189894
R128 VP.n67 VP.n6 0.189894
R129 VP.n71 VP.n6 0.189894
R130 VP.n72 VP.n71 0.189894
R131 VP.n73 VP.n72 0.189894
R132 VP.n73 VP.n4 0.189894
R133 VP.n78 VP.n4 0.189894
R134 VP.n79 VP.n78 0.189894
R135 VP.n80 VP.n79 0.189894
R136 VP.n80 VP.n2 0.189894
R137 VP.n84 VP.n2 0.189894
R138 VP.n85 VP.n84 0.189894
R139 VP.n86 VP.n85 0.189894
R140 VP.n86 VP.n0 0.189894
R141 VTAIL.n626 VTAIL.n554 756.745
R142 VTAIL.n74 VTAIL.n2 756.745
R143 VTAIL.n152 VTAIL.n80 756.745
R144 VTAIL.n232 VTAIL.n160 756.745
R145 VTAIL.n548 VTAIL.n476 756.745
R146 VTAIL.n468 VTAIL.n396 756.745
R147 VTAIL.n390 VTAIL.n318 756.745
R148 VTAIL.n310 VTAIL.n238 756.745
R149 VTAIL.n578 VTAIL.n577 585
R150 VTAIL.n583 VTAIL.n582 585
R151 VTAIL.n585 VTAIL.n584 585
R152 VTAIL.n574 VTAIL.n573 585
R153 VTAIL.n591 VTAIL.n590 585
R154 VTAIL.n593 VTAIL.n592 585
R155 VTAIL.n570 VTAIL.n569 585
R156 VTAIL.n599 VTAIL.n598 585
R157 VTAIL.n601 VTAIL.n600 585
R158 VTAIL.n566 VTAIL.n565 585
R159 VTAIL.n607 VTAIL.n606 585
R160 VTAIL.n609 VTAIL.n608 585
R161 VTAIL.n562 VTAIL.n561 585
R162 VTAIL.n615 VTAIL.n614 585
R163 VTAIL.n617 VTAIL.n616 585
R164 VTAIL.n558 VTAIL.n557 585
R165 VTAIL.n624 VTAIL.n623 585
R166 VTAIL.n625 VTAIL.n556 585
R167 VTAIL.n627 VTAIL.n626 585
R168 VTAIL.n26 VTAIL.n25 585
R169 VTAIL.n31 VTAIL.n30 585
R170 VTAIL.n33 VTAIL.n32 585
R171 VTAIL.n22 VTAIL.n21 585
R172 VTAIL.n39 VTAIL.n38 585
R173 VTAIL.n41 VTAIL.n40 585
R174 VTAIL.n18 VTAIL.n17 585
R175 VTAIL.n47 VTAIL.n46 585
R176 VTAIL.n49 VTAIL.n48 585
R177 VTAIL.n14 VTAIL.n13 585
R178 VTAIL.n55 VTAIL.n54 585
R179 VTAIL.n57 VTAIL.n56 585
R180 VTAIL.n10 VTAIL.n9 585
R181 VTAIL.n63 VTAIL.n62 585
R182 VTAIL.n65 VTAIL.n64 585
R183 VTAIL.n6 VTAIL.n5 585
R184 VTAIL.n72 VTAIL.n71 585
R185 VTAIL.n73 VTAIL.n4 585
R186 VTAIL.n75 VTAIL.n74 585
R187 VTAIL.n104 VTAIL.n103 585
R188 VTAIL.n109 VTAIL.n108 585
R189 VTAIL.n111 VTAIL.n110 585
R190 VTAIL.n100 VTAIL.n99 585
R191 VTAIL.n117 VTAIL.n116 585
R192 VTAIL.n119 VTAIL.n118 585
R193 VTAIL.n96 VTAIL.n95 585
R194 VTAIL.n125 VTAIL.n124 585
R195 VTAIL.n127 VTAIL.n126 585
R196 VTAIL.n92 VTAIL.n91 585
R197 VTAIL.n133 VTAIL.n132 585
R198 VTAIL.n135 VTAIL.n134 585
R199 VTAIL.n88 VTAIL.n87 585
R200 VTAIL.n141 VTAIL.n140 585
R201 VTAIL.n143 VTAIL.n142 585
R202 VTAIL.n84 VTAIL.n83 585
R203 VTAIL.n150 VTAIL.n149 585
R204 VTAIL.n151 VTAIL.n82 585
R205 VTAIL.n153 VTAIL.n152 585
R206 VTAIL.n184 VTAIL.n183 585
R207 VTAIL.n189 VTAIL.n188 585
R208 VTAIL.n191 VTAIL.n190 585
R209 VTAIL.n180 VTAIL.n179 585
R210 VTAIL.n197 VTAIL.n196 585
R211 VTAIL.n199 VTAIL.n198 585
R212 VTAIL.n176 VTAIL.n175 585
R213 VTAIL.n205 VTAIL.n204 585
R214 VTAIL.n207 VTAIL.n206 585
R215 VTAIL.n172 VTAIL.n171 585
R216 VTAIL.n213 VTAIL.n212 585
R217 VTAIL.n215 VTAIL.n214 585
R218 VTAIL.n168 VTAIL.n167 585
R219 VTAIL.n221 VTAIL.n220 585
R220 VTAIL.n223 VTAIL.n222 585
R221 VTAIL.n164 VTAIL.n163 585
R222 VTAIL.n230 VTAIL.n229 585
R223 VTAIL.n231 VTAIL.n162 585
R224 VTAIL.n233 VTAIL.n232 585
R225 VTAIL.n549 VTAIL.n548 585
R226 VTAIL.n547 VTAIL.n478 585
R227 VTAIL.n546 VTAIL.n545 585
R228 VTAIL.n481 VTAIL.n479 585
R229 VTAIL.n540 VTAIL.n539 585
R230 VTAIL.n538 VTAIL.n537 585
R231 VTAIL.n485 VTAIL.n484 585
R232 VTAIL.n532 VTAIL.n531 585
R233 VTAIL.n530 VTAIL.n529 585
R234 VTAIL.n489 VTAIL.n488 585
R235 VTAIL.n524 VTAIL.n523 585
R236 VTAIL.n522 VTAIL.n521 585
R237 VTAIL.n493 VTAIL.n492 585
R238 VTAIL.n516 VTAIL.n515 585
R239 VTAIL.n514 VTAIL.n513 585
R240 VTAIL.n497 VTAIL.n496 585
R241 VTAIL.n508 VTAIL.n507 585
R242 VTAIL.n506 VTAIL.n505 585
R243 VTAIL.n501 VTAIL.n500 585
R244 VTAIL.n469 VTAIL.n468 585
R245 VTAIL.n467 VTAIL.n398 585
R246 VTAIL.n466 VTAIL.n465 585
R247 VTAIL.n401 VTAIL.n399 585
R248 VTAIL.n460 VTAIL.n459 585
R249 VTAIL.n458 VTAIL.n457 585
R250 VTAIL.n405 VTAIL.n404 585
R251 VTAIL.n452 VTAIL.n451 585
R252 VTAIL.n450 VTAIL.n449 585
R253 VTAIL.n409 VTAIL.n408 585
R254 VTAIL.n444 VTAIL.n443 585
R255 VTAIL.n442 VTAIL.n441 585
R256 VTAIL.n413 VTAIL.n412 585
R257 VTAIL.n436 VTAIL.n435 585
R258 VTAIL.n434 VTAIL.n433 585
R259 VTAIL.n417 VTAIL.n416 585
R260 VTAIL.n428 VTAIL.n427 585
R261 VTAIL.n426 VTAIL.n425 585
R262 VTAIL.n421 VTAIL.n420 585
R263 VTAIL.n391 VTAIL.n390 585
R264 VTAIL.n389 VTAIL.n320 585
R265 VTAIL.n388 VTAIL.n387 585
R266 VTAIL.n323 VTAIL.n321 585
R267 VTAIL.n382 VTAIL.n381 585
R268 VTAIL.n380 VTAIL.n379 585
R269 VTAIL.n327 VTAIL.n326 585
R270 VTAIL.n374 VTAIL.n373 585
R271 VTAIL.n372 VTAIL.n371 585
R272 VTAIL.n331 VTAIL.n330 585
R273 VTAIL.n366 VTAIL.n365 585
R274 VTAIL.n364 VTAIL.n363 585
R275 VTAIL.n335 VTAIL.n334 585
R276 VTAIL.n358 VTAIL.n357 585
R277 VTAIL.n356 VTAIL.n355 585
R278 VTAIL.n339 VTAIL.n338 585
R279 VTAIL.n350 VTAIL.n349 585
R280 VTAIL.n348 VTAIL.n347 585
R281 VTAIL.n343 VTAIL.n342 585
R282 VTAIL.n311 VTAIL.n310 585
R283 VTAIL.n309 VTAIL.n240 585
R284 VTAIL.n308 VTAIL.n307 585
R285 VTAIL.n243 VTAIL.n241 585
R286 VTAIL.n302 VTAIL.n301 585
R287 VTAIL.n300 VTAIL.n299 585
R288 VTAIL.n247 VTAIL.n246 585
R289 VTAIL.n294 VTAIL.n293 585
R290 VTAIL.n292 VTAIL.n291 585
R291 VTAIL.n251 VTAIL.n250 585
R292 VTAIL.n286 VTAIL.n285 585
R293 VTAIL.n284 VTAIL.n283 585
R294 VTAIL.n255 VTAIL.n254 585
R295 VTAIL.n278 VTAIL.n277 585
R296 VTAIL.n276 VTAIL.n275 585
R297 VTAIL.n259 VTAIL.n258 585
R298 VTAIL.n270 VTAIL.n269 585
R299 VTAIL.n268 VTAIL.n267 585
R300 VTAIL.n263 VTAIL.n262 585
R301 VTAIL.n579 VTAIL.t6 327.466
R302 VTAIL.n27 VTAIL.t5 327.466
R303 VTAIL.n105 VTAIL.t11 327.466
R304 VTAIL.n185 VTAIL.t9 327.466
R305 VTAIL.n502 VTAIL.t13 327.466
R306 VTAIL.n422 VTAIL.t12 327.466
R307 VTAIL.n344 VTAIL.t7 327.466
R308 VTAIL.n264 VTAIL.t1 327.466
R309 VTAIL.n583 VTAIL.n577 171.744
R310 VTAIL.n584 VTAIL.n583 171.744
R311 VTAIL.n584 VTAIL.n573 171.744
R312 VTAIL.n591 VTAIL.n573 171.744
R313 VTAIL.n592 VTAIL.n591 171.744
R314 VTAIL.n592 VTAIL.n569 171.744
R315 VTAIL.n599 VTAIL.n569 171.744
R316 VTAIL.n600 VTAIL.n599 171.744
R317 VTAIL.n600 VTAIL.n565 171.744
R318 VTAIL.n607 VTAIL.n565 171.744
R319 VTAIL.n608 VTAIL.n607 171.744
R320 VTAIL.n608 VTAIL.n561 171.744
R321 VTAIL.n615 VTAIL.n561 171.744
R322 VTAIL.n616 VTAIL.n615 171.744
R323 VTAIL.n616 VTAIL.n557 171.744
R324 VTAIL.n624 VTAIL.n557 171.744
R325 VTAIL.n625 VTAIL.n624 171.744
R326 VTAIL.n626 VTAIL.n625 171.744
R327 VTAIL.n31 VTAIL.n25 171.744
R328 VTAIL.n32 VTAIL.n31 171.744
R329 VTAIL.n32 VTAIL.n21 171.744
R330 VTAIL.n39 VTAIL.n21 171.744
R331 VTAIL.n40 VTAIL.n39 171.744
R332 VTAIL.n40 VTAIL.n17 171.744
R333 VTAIL.n47 VTAIL.n17 171.744
R334 VTAIL.n48 VTAIL.n47 171.744
R335 VTAIL.n48 VTAIL.n13 171.744
R336 VTAIL.n55 VTAIL.n13 171.744
R337 VTAIL.n56 VTAIL.n55 171.744
R338 VTAIL.n56 VTAIL.n9 171.744
R339 VTAIL.n63 VTAIL.n9 171.744
R340 VTAIL.n64 VTAIL.n63 171.744
R341 VTAIL.n64 VTAIL.n5 171.744
R342 VTAIL.n72 VTAIL.n5 171.744
R343 VTAIL.n73 VTAIL.n72 171.744
R344 VTAIL.n74 VTAIL.n73 171.744
R345 VTAIL.n109 VTAIL.n103 171.744
R346 VTAIL.n110 VTAIL.n109 171.744
R347 VTAIL.n110 VTAIL.n99 171.744
R348 VTAIL.n117 VTAIL.n99 171.744
R349 VTAIL.n118 VTAIL.n117 171.744
R350 VTAIL.n118 VTAIL.n95 171.744
R351 VTAIL.n125 VTAIL.n95 171.744
R352 VTAIL.n126 VTAIL.n125 171.744
R353 VTAIL.n126 VTAIL.n91 171.744
R354 VTAIL.n133 VTAIL.n91 171.744
R355 VTAIL.n134 VTAIL.n133 171.744
R356 VTAIL.n134 VTAIL.n87 171.744
R357 VTAIL.n141 VTAIL.n87 171.744
R358 VTAIL.n142 VTAIL.n141 171.744
R359 VTAIL.n142 VTAIL.n83 171.744
R360 VTAIL.n150 VTAIL.n83 171.744
R361 VTAIL.n151 VTAIL.n150 171.744
R362 VTAIL.n152 VTAIL.n151 171.744
R363 VTAIL.n189 VTAIL.n183 171.744
R364 VTAIL.n190 VTAIL.n189 171.744
R365 VTAIL.n190 VTAIL.n179 171.744
R366 VTAIL.n197 VTAIL.n179 171.744
R367 VTAIL.n198 VTAIL.n197 171.744
R368 VTAIL.n198 VTAIL.n175 171.744
R369 VTAIL.n205 VTAIL.n175 171.744
R370 VTAIL.n206 VTAIL.n205 171.744
R371 VTAIL.n206 VTAIL.n171 171.744
R372 VTAIL.n213 VTAIL.n171 171.744
R373 VTAIL.n214 VTAIL.n213 171.744
R374 VTAIL.n214 VTAIL.n167 171.744
R375 VTAIL.n221 VTAIL.n167 171.744
R376 VTAIL.n222 VTAIL.n221 171.744
R377 VTAIL.n222 VTAIL.n163 171.744
R378 VTAIL.n230 VTAIL.n163 171.744
R379 VTAIL.n231 VTAIL.n230 171.744
R380 VTAIL.n232 VTAIL.n231 171.744
R381 VTAIL.n548 VTAIL.n547 171.744
R382 VTAIL.n547 VTAIL.n546 171.744
R383 VTAIL.n546 VTAIL.n479 171.744
R384 VTAIL.n539 VTAIL.n479 171.744
R385 VTAIL.n539 VTAIL.n538 171.744
R386 VTAIL.n538 VTAIL.n484 171.744
R387 VTAIL.n531 VTAIL.n484 171.744
R388 VTAIL.n531 VTAIL.n530 171.744
R389 VTAIL.n530 VTAIL.n488 171.744
R390 VTAIL.n523 VTAIL.n488 171.744
R391 VTAIL.n523 VTAIL.n522 171.744
R392 VTAIL.n522 VTAIL.n492 171.744
R393 VTAIL.n515 VTAIL.n492 171.744
R394 VTAIL.n515 VTAIL.n514 171.744
R395 VTAIL.n514 VTAIL.n496 171.744
R396 VTAIL.n507 VTAIL.n496 171.744
R397 VTAIL.n507 VTAIL.n506 171.744
R398 VTAIL.n506 VTAIL.n500 171.744
R399 VTAIL.n468 VTAIL.n467 171.744
R400 VTAIL.n467 VTAIL.n466 171.744
R401 VTAIL.n466 VTAIL.n399 171.744
R402 VTAIL.n459 VTAIL.n399 171.744
R403 VTAIL.n459 VTAIL.n458 171.744
R404 VTAIL.n458 VTAIL.n404 171.744
R405 VTAIL.n451 VTAIL.n404 171.744
R406 VTAIL.n451 VTAIL.n450 171.744
R407 VTAIL.n450 VTAIL.n408 171.744
R408 VTAIL.n443 VTAIL.n408 171.744
R409 VTAIL.n443 VTAIL.n442 171.744
R410 VTAIL.n442 VTAIL.n412 171.744
R411 VTAIL.n435 VTAIL.n412 171.744
R412 VTAIL.n435 VTAIL.n434 171.744
R413 VTAIL.n434 VTAIL.n416 171.744
R414 VTAIL.n427 VTAIL.n416 171.744
R415 VTAIL.n427 VTAIL.n426 171.744
R416 VTAIL.n426 VTAIL.n420 171.744
R417 VTAIL.n390 VTAIL.n389 171.744
R418 VTAIL.n389 VTAIL.n388 171.744
R419 VTAIL.n388 VTAIL.n321 171.744
R420 VTAIL.n381 VTAIL.n321 171.744
R421 VTAIL.n381 VTAIL.n380 171.744
R422 VTAIL.n380 VTAIL.n326 171.744
R423 VTAIL.n373 VTAIL.n326 171.744
R424 VTAIL.n373 VTAIL.n372 171.744
R425 VTAIL.n372 VTAIL.n330 171.744
R426 VTAIL.n365 VTAIL.n330 171.744
R427 VTAIL.n365 VTAIL.n364 171.744
R428 VTAIL.n364 VTAIL.n334 171.744
R429 VTAIL.n357 VTAIL.n334 171.744
R430 VTAIL.n357 VTAIL.n356 171.744
R431 VTAIL.n356 VTAIL.n338 171.744
R432 VTAIL.n349 VTAIL.n338 171.744
R433 VTAIL.n349 VTAIL.n348 171.744
R434 VTAIL.n348 VTAIL.n342 171.744
R435 VTAIL.n310 VTAIL.n309 171.744
R436 VTAIL.n309 VTAIL.n308 171.744
R437 VTAIL.n308 VTAIL.n241 171.744
R438 VTAIL.n301 VTAIL.n241 171.744
R439 VTAIL.n301 VTAIL.n300 171.744
R440 VTAIL.n300 VTAIL.n246 171.744
R441 VTAIL.n293 VTAIL.n246 171.744
R442 VTAIL.n293 VTAIL.n292 171.744
R443 VTAIL.n292 VTAIL.n250 171.744
R444 VTAIL.n285 VTAIL.n250 171.744
R445 VTAIL.n285 VTAIL.n284 171.744
R446 VTAIL.n284 VTAIL.n254 171.744
R447 VTAIL.n277 VTAIL.n254 171.744
R448 VTAIL.n277 VTAIL.n276 171.744
R449 VTAIL.n276 VTAIL.n258 171.744
R450 VTAIL.n269 VTAIL.n258 171.744
R451 VTAIL.n269 VTAIL.n268 171.744
R452 VTAIL.n268 VTAIL.n262 171.744
R453 VTAIL.t6 VTAIL.n577 85.8723
R454 VTAIL.t5 VTAIL.n25 85.8723
R455 VTAIL.t11 VTAIL.n103 85.8723
R456 VTAIL.t9 VTAIL.n183 85.8723
R457 VTAIL.t13 VTAIL.n500 85.8723
R458 VTAIL.t12 VTAIL.n420 85.8723
R459 VTAIL.t7 VTAIL.n342 85.8723
R460 VTAIL.t1 VTAIL.n262 85.8723
R461 VTAIL.n475 VTAIL.n474 58.7283
R462 VTAIL.n317 VTAIL.n316 58.7283
R463 VTAIL.n1 VTAIL.n0 58.7281
R464 VTAIL.n159 VTAIL.n158 58.7281
R465 VTAIL.n631 VTAIL.n630 36.2581
R466 VTAIL.n79 VTAIL.n78 36.2581
R467 VTAIL.n157 VTAIL.n156 36.2581
R468 VTAIL.n237 VTAIL.n236 36.2581
R469 VTAIL.n553 VTAIL.n552 36.2581
R470 VTAIL.n473 VTAIL.n472 36.2581
R471 VTAIL.n395 VTAIL.n394 36.2581
R472 VTAIL.n315 VTAIL.n314 36.2581
R473 VTAIL.n631 VTAIL.n553 28.1083
R474 VTAIL.n315 VTAIL.n237 28.1083
R475 VTAIL.n579 VTAIL.n578 16.3895
R476 VTAIL.n27 VTAIL.n26 16.3895
R477 VTAIL.n105 VTAIL.n104 16.3895
R478 VTAIL.n185 VTAIL.n184 16.3895
R479 VTAIL.n502 VTAIL.n501 16.3895
R480 VTAIL.n422 VTAIL.n421 16.3895
R481 VTAIL.n344 VTAIL.n343 16.3895
R482 VTAIL.n264 VTAIL.n263 16.3895
R483 VTAIL.n627 VTAIL.n556 13.1884
R484 VTAIL.n75 VTAIL.n4 13.1884
R485 VTAIL.n153 VTAIL.n82 13.1884
R486 VTAIL.n233 VTAIL.n162 13.1884
R487 VTAIL.n549 VTAIL.n478 13.1884
R488 VTAIL.n469 VTAIL.n398 13.1884
R489 VTAIL.n391 VTAIL.n320 13.1884
R490 VTAIL.n311 VTAIL.n240 13.1884
R491 VTAIL.n582 VTAIL.n581 12.8005
R492 VTAIL.n623 VTAIL.n622 12.8005
R493 VTAIL.n628 VTAIL.n554 12.8005
R494 VTAIL.n30 VTAIL.n29 12.8005
R495 VTAIL.n71 VTAIL.n70 12.8005
R496 VTAIL.n76 VTAIL.n2 12.8005
R497 VTAIL.n108 VTAIL.n107 12.8005
R498 VTAIL.n149 VTAIL.n148 12.8005
R499 VTAIL.n154 VTAIL.n80 12.8005
R500 VTAIL.n188 VTAIL.n187 12.8005
R501 VTAIL.n229 VTAIL.n228 12.8005
R502 VTAIL.n234 VTAIL.n160 12.8005
R503 VTAIL.n550 VTAIL.n476 12.8005
R504 VTAIL.n545 VTAIL.n480 12.8005
R505 VTAIL.n505 VTAIL.n504 12.8005
R506 VTAIL.n470 VTAIL.n396 12.8005
R507 VTAIL.n465 VTAIL.n400 12.8005
R508 VTAIL.n425 VTAIL.n424 12.8005
R509 VTAIL.n392 VTAIL.n318 12.8005
R510 VTAIL.n387 VTAIL.n322 12.8005
R511 VTAIL.n347 VTAIL.n346 12.8005
R512 VTAIL.n312 VTAIL.n238 12.8005
R513 VTAIL.n307 VTAIL.n242 12.8005
R514 VTAIL.n267 VTAIL.n266 12.8005
R515 VTAIL.n585 VTAIL.n576 12.0247
R516 VTAIL.n621 VTAIL.n558 12.0247
R517 VTAIL.n33 VTAIL.n24 12.0247
R518 VTAIL.n69 VTAIL.n6 12.0247
R519 VTAIL.n111 VTAIL.n102 12.0247
R520 VTAIL.n147 VTAIL.n84 12.0247
R521 VTAIL.n191 VTAIL.n182 12.0247
R522 VTAIL.n227 VTAIL.n164 12.0247
R523 VTAIL.n544 VTAIL.n481 12.0247
R524 VTAIL.n508 VTAIL.n499 12.0247
R525 VTAIL.n464 VTAIL.n401 12.0247
R526 VTAIL.n428 VTAIL.n419 12.0247
R527 VTAIL.n386 VTAIL.n323 12.0247
R528 VTAIL.n350 VTAIL.n341 12.0247
R529 VTAIL.n306 VTAIL.n243 12.0247
R530 VTAIL.n270 VTAIL.n261 12.0247
R531 VTAIL.n586 VTAIL.n574 11.249
R532 VTAIL.n618 VTAIL.n617 11.249
R533 VTAIL.n34 VTAIL.n22 11.249
R534 VTAIL.n66 VTAIL.n65 11.249
R535 VTAIL.n112 VTAIL.n100 11.249
R536 VTAIL.n144 VTAIL.n143 11.249
R537 VTAIL.n192 VTAIL.n180 11.249
R538 VTAIL.n224 VTAIL.n223 11.249
R539 VTAIL.n541 VTAIL.n540 11.249
R540 VTAIL.n509 VTAIL.n497 11.249
R541 VTAIL.n461 VTAIL.n460 11.249
R542 VTAIL.n429 VTAIL.n417 11.249
R543 VTAIL.n383 VTAIL.n382 11.249
R544 VTAIL.n351 VTAIL.n339 11.249
R545 VTAIL.n303 VTAIL.n302 11.249
R546 VTAIL.n271 VTAIL.n259 11.249
R547 VTAIL.n590 VTAIL.n589 10.4732
R548 VTAIL.n614 VTAIL.n560 10.4732
R549 VTAIL.n38 VTAIL.n37 10.4732
R550 VTAIL.n62 VTAIL.n8 10.4732
R551 VTAIL.n116 VTAIL.n115 10.4732
R552 VTAIL.n140 VTAIL.n86 10.4732
R553 VTAIL.n196 VTAIL.n195 10.4732
R554 VTAIL.n220 VTAIL.n166 10.4732
R555 VTAIL.n537 VTAIL.n483 10.4732
R556 VTAIL.n513 VTAIL.n512 10.4732
R557 VTAIL.n457 VTAIL.n403 10.4732
R558 VTAIL.n433 VTAIL.n432 10.4732
R559 VTAIL.n379 VTAIL.n325 10.4732
R560 VTAIL.n355 VTAIL.n354 10.4732
R561 VTAIL.n299 VTAIL.n245 10.4732
R562 VTAIL.n275 VTAIL.n274 10.4732
R563 VTAIL.n593 VTAIL.n572 9.69747
R564 VTAIL.n613 VTAIL.n562 9.69747
R565 VTAIL.n41 VTAIL.n20 9.69747
R566 VTAIL.n61 VTAIL.n10 9.69747
R567 VTAIL.n119 VTAIL.n98 9.69747
R568 VTAIL.n139 VTAIL.n88 9.69747
R569 VTAIL.n199 VTAIL.n178 9.69747
R570 VTAIL.n219 VTAIL.n168 9.69747
R571 VTAIL.n536 VTAIL.n485 9.69747
R572 VTAIL.n516 VTAIL.n495 9.69747
R573 VTAIL.n456 VTAIL.n405 9.69747
R574 VTAIL.n436 VTAIL.n415 9.69747
R575 VTAIL.n378 VTAIL.n327 9.69747
R576 VTAIL.n358 VTAIL.n337 9.69747
R577 VTAIL.n298 VTAIL.n247 9.69747
R578 VTAIL.n278 VTAIL.n257 9.69747
R579 VTAIL.n630 VTAIL.n629 9.45567
R580 VTAIL.n78 VTAIL.n77 9.45567
R581 VTAIL.n156 VTAIL.n155 9.45567
R582 VTAIL.n236 VTAIL.n235 9.45567
R583 VTAIL.n552 VTAIL.n551 9.45567
R584 VTAIL.n472 VTAIL.n471 9.45567
R585 VTAIL.n394 VTAIL.n393 9.45567
R586 VTAIL.n314 VTAIL.n313 9.45567
R587 VTAIL.n629 VTAIL.n628 9.3005
R588 VTAIL.n568 VTAIL.n567 9.3005
R589 VTAIL.n597 VTAIL.n596 9.3005
R590 VTAIL.n595 VTAIL.n594 9.3005
R591 VTAIL.n572 VTAIL.n571 9.3005
R592 VTAIL.n589 VTAIL.n588 9.3005
R593 VTAIL.n587 VTAIL.n586 9.3005
R594 VTAIL.n576 VTAIL.n575 9.3005
R595 VTAIL.n581 VTAIL.n580 9.3005
R596 VTAIL.n603 VTAIL.n602 9.3005
R597 VTAIL.n605 VTAIL.n604 9.3005
R598 VTAIL.n564 VTAIL.n563 9.3005
R599 VTAIL.n611 VTAIL.n610 9.3005
R600 VTAIL.n613 VTAIL.n612 9.3005
R601 VTAIL.n560 VTAIL.n559 9.3005
R602 VTAIL.n619 VTAIL.n618 9.3005
R603 VTAIL.n621 VTAIL.n620 9.3005
R604 VTAIL.n622 VTAIL.n555 9.3005
R605 VTAIL.n77 VTAIL.n76 9.3005
R606 VTAIL.n16 VTAIL.n15 9.3005
R607 VTAIL.n45 VTAIL.n44 9.3005
R608 VTAIL.n43 VTAIL.n42 9.3005
R609 VTAIL.n20 VTAIL.n19 9.3005
R610 VTAIL.n37 VTAIL.n36 9.3005
R611 VTAIL.n35 VTAIL.n34 9.3005
R612 VTAIL.n24 VTAIL.n23 9.3005
R613 VTAIL.n29 VTAIL.n28 9.3005
R614 VTAIL.n51 VTAIL.n50 9.3005
R615 VTAIL.n53 VTAIL.n52 9.3005
R616 VTAIL.n12 VTAIL.n11 9.3005
R617 VTAIL.n59 VTAIL.n58 9.3005
R618 VTAIL.n61 VTAIL.n60 9.3005
R619 VTAIL.n8 VTAIL.n7 9.3005
R620 VTAIL.n67 VTAIL.n66 9.3005
R621 VTAIL.n69 VTAIL.n68 9.3005
R622 VTAIL.n70 VTAIL.n3 9.3005
R623 VTAIL.n155 VTAIL.n154 9.3005
R624 VTAIL.n94 VTAIL.n93 9.3005
R625 VTAIL.n123 VTAIL.n122 9.3005
R626 VTAIL.n121 VTAIL.n120 9.3005
R627 VTAIL.n98 VTAIL.n97 9.3005
R628 VTAIL.n115 VTAIL.n114 9.3005
R629 VTAIL.n113 VTAIL.n112 9.3005
R630 VTAIL.n102 VTAIL.n101 9.3005
R631 VTAIL.n107 VTAIL.n106 9.3005
R632 VTAIL.n129 VTAIL.n128 9.3005
R633 VTAIL.n131 VTAIL.n130 9.3005
R634 VTAIL.n90 VTAIL.n89 9.3005
R635 VTAIL.n137 VTAIL.n136 9.3005
R636 VTAIL.n139 VTAIL.n138 9.3005
R637 VTAIL.n86 VTAIL.n85 9.3005
R638 VTAIL.n145 VTAIL.n144 9.3005
R639 VTAIL.n147 VTAIL.n146 9.3005
R640 VTAIL.n148 VTAIL.n81 9.3005
R641 VTAIL.n235 VTAIL.n234 9.3005
R642 VTAIL.n174 VTAIL.n173 9.3005
R643 VTAIL.n203 VTAIL.n202 9.3005
R644 VTAIL.n201 VTAIL.n200 9.3005
R645 VTAIL.n178 VTAIL.n177 9.3005
R646 VTAIL.n195 VTAIL.n194 9.3005
R647 VTAIL.n193 VTAIL.n192 9.3005
R648 VTAIL.n182 VTAIL.n181 9.3005
R649 VTAIL.n187 VTAIL.n186 9.3005
R650 VTAIL.n209 VTAIL.n208 9.3005
R651 VTAIL.n211 VTAIL.n210 9.3005
R652 VTAIL.n170 VTAIL.n169 9.3005
R653 VTAIL.n217 VTAIL.n216 9.3005
R654 VTAIL.n219 VTAIL.n218 9.3005
R655 VTAIL.n166 VTAIL.n165 9.3005
R656 VTAIL.n225 VTAIL.n224 9.3005
R657 VTAIL.n227 VTAIL.n226 9.3005
R658 VTAIL.n228 VTAIL.n161 9.3005
R659 VTAIL.n528 VTAIL.n527 9.3005
R660 VTAIL.n487 VTAIL.n486 9.3005
R661 VTAIL.n534 VTAIL.n533 9.3005
R662 VTAIL.n536 VTAIL.n535 9.3005
R663 VTAIL.n483 VTAIL.n482 9.3005
R664 VTAIL.n542 VTAIL.n541 9.3005
R665 VTAIL.n544 VTAIL.n543 9.3005
R666 VTAIL.n480 VTAIL.n477 9.3005
R667 VTAIL.n551 VTAIL.n550 9.3005
R668 VTAIL.n526 VTAIL.n525 9.3005
R669 VTAIL.n491 VTAIL.n490 9.3005
R670 VTAIL.n520 VTAIL.n519 9.3005
R671 VTAIL.n518 VTAIL.n517 9.3005
R672 VTAIL.n495 VTAIL.n494 9.3005
R673 VTAIL.n512 VTAIL.n511 9.3005
R674 VTAIL.n510 VTAIL.n509 9.3005
R675 VTAIL.n499 VTAIL.n498 9.3005
R676 VTAIL.n504 VTAIL.n503 9.3005
R677 VTAIL.n448 VTAIL.n447 9.3005
R678 VTAIL.n407 VTAIL.n406 9.3005
R679 VTAIL.n454 VTAIL.n453 9.3005
R680 VTAIL.n456 VTAIL.n455 9.3005
R681 VTAIL.n403 VTAIL.n402 9.3005
R682 VTAIL.n462 VTAIL.n461 9.3005
R683 VTAIL.n464 VTAIL.n463 9.3005
R684 VTAIL.n400 VTAIL.n397 9.3005
R685 VTAIL.n471 VTAIL.n470 9.3005
R686 VTAIL.n446 VTAIL.n445 9.3005
R687 VTAIL.n411 VTAIL.n410 9.3005
R688 VTAIL.n440 VTAIL.n439 9.3005
R689 VTAIL.n438 VTAIL.n437 9.3005
R690 VTAIL.n415 VTAIL.n414 9.3005
R691 VTAIL.n432 VTAIL.n431 9.3005
R692 VTAIL.n430 VTAIL.n429 9.3005
R693 VTAIL.n419 VTAIL.n418 9.3005
R694 VTAIL.n424 VTAIL.n423 9.3005
R695 VTAIL.n370 VTAIL.n369 9.3005
R696 VTAIL.n329 VTAIL.n328 9.3005
R697 VTAIL.n376 VTAIL.n375 9.3005
R698 VTAIL.n378 VTAIL.n377 9.3005
R699 VTAIL.n325 VTAIL.n324 9.3005
R700 VTAIL.n384 VTAIL.n383 9.3005
R701 VTAIL.n386 VTAIL.n385 9.3005
R702 VTAIL.n322 VTAIL.n319 9.3005
R703 VTAIL.n393 VTAIL.n392 9.3005
R704 VTAIL.n368 VTAIL.n367 9.3005
R705 VTAIL.n333 VTAIL.n332 9.3005
R706 VTAIL.n362 VTAIL.n361 9.3005
R707 VTAIL.n360 VTAIL.n359 9.3005
R708 VTAIL.n337 VTAIL.n336 9.3005
R709 VTAIL.n354 VTAIL.n353 9.3005
R710 VTAIL.n352 VTAIL.n351 9.3005
R711 VTAIL.n341 VTAIL.n340 9.3005
R712 VTAIL.n346 VTAIL.n345 9.3005
R713 VTAIL.n290 VTAIL.n289 9.3005
R714 VTAIL.n249 VTAIL.n248 9.3005
R715 VTAIL.n296 VTAIL.n295 9.3005
R716 VTAIL.n298 VTAIL.n297 9.3005
R717 VTAIL.n245 VTAIL.n244 9.3005
R718 VTAIL.n304 VTAIL.n303 9.3005
R719 VTAIL.n306 VTAIL.n305 9.3005
R720 VTAIL.n242 VTAIL.n239 9.3005
R721 VTAIL.n313 VTAIL.n312 9.3005
R722 VTAIL.n288 VTAIL.n287 9.3005
R723 VTAIL.n253 VTAIL.n252 9.3005
R724 VTAIL.n282 VTAIL.n281 9.3005
R725 VTAIL.n280 VTAIL.n279 9.3005
R726 VTAIL.n257 VTAIL.n256 9.3005
R727 VTAIL.n274 VTAIL.n273 9.3005
R728 VTAIL.n272 VTAIL.n271 9.3005
R729 VTAIL.n261 VTAIL.n260 9.3005
R730 VTAIL.n266 VTAIL.n265 9.3005
R731 VTAIL.n594 VTAIL.n570 8.92171
R732 VTAIL.n610 VTAIL.n609 8.92171
R733 VTAIL.n42 VTAIL.n18 8.92171
R734 VTAIL.n58 VTAIL.n57 8.92171
R735 VTAIL.n120 VTAIL.n96 8.92171
R736 VTAIL.n136 VTAIL.n135 8.92171
R737 VTAIL.n200 VTAIL.n176 8.92171
R738 VTAIL.n216 VTAIL.n215 8.92171
R739 VTAIL.n533 VTAIL.n532 8.92171
R740 VTAIL.n517 VTAIL.n493 8.92171
R741 VTAIL.n453 VTAIL.n452 8.92171
R742 VTAIL.n437 VTAIL.n413 8.92171
R743 VTAIL.n375 VTAIL.n374 8.92171
R744 VTAIL.n359 VTAIL.n335 8.92171
R745 VTAIL.n295 VTAIL.n294 8.92171
R746 VTAIL.n279 VTAIL.n255 8.92171
R747 VTAIL.n598 VTAIL.n597 8.14595
R748 VTAIL.n606 VTAIL.n564 8.14595
R749 VTAIL.n46 VTAIL.n45 8.14595
R750 VTAIL.n54 VTAIL.n12 8.14595
R751 VTAIL.n124 VTAIL.n123 8.14595
R752 VTAIL.n132 VTAIL.n90 8.14595
R753 VTAIL.n204 VTAIL.n203 8.14595
R754 VTAIL.n212 VTAIL.n170 8.14595
R755 VTAIL.n529 VTAIL.n487 8.14595
R756 VTAIL.n521 VTAIL.n520 8.14595
R757 VTAIL.n449 VTAIL.n407 8.14595
R758 VTAIL.n441 VTAIL.n440 8.14595
R759 VTAIL.n371 VTAIL.n329 8.14595
R760 VTAIL.n363 VTAIL.n362 8.14595
R761 VTAIL.n291 VTAIL.n249 8.14595
R762 VTAIL.n283 VTAIL.n282 8.14595
R763 VTAIL.n601 VTAIL.n568 7.3702
R764 VTAIL.n605 VTAIL.n566 7.3702
R765 VTAIL.n49 VTAIL.n16 7.3702
R766 VTAIL.n53 VTAIL.n14 7.3702
R767 VTAIL.n127 VTAIL.n94 7.3702
R768 VTAIL.n131 VTAIL.n92 7.3702
R769 VTAIL.n207 VTAIL.n174 7.3702
R770 VTAIL.n211 VTAIL.n172 7.3702
R771 VTAIL.n528 VTAIL.n489 7.3702
R772 VTAIL.n524 VTAIL.n491 7.3702
R773 VTAIL.n448 VTAIL.n409 7.3702
R774 VTAIL.n444 VTAIL.n411 7.3702
R775 VTAIL.n370 VTAIL.n331 7.3702
R776 VTAIL.n366 VTAIL.n333 7.3702
R777 VTAIL.n290 VTAIL.n251 7.3702
R778 VTAIL.n286 VTAIL.n253 7.3702
R779 VTAIL.n602 VTAIL.n601 6.59444
R780 VTAIL.n602 VTAIL.n566 6.59444
R781 VTAIL.n50 VTAIL.n49 6.59444
R782 VTAIL.n50 VTAIL.n14 6.59444
R783 VTAIL.n128 VTAIL.n127 6.59444
R784 VTAIL.n128 VTAIL.n92 6.59444
R785 VTAIL.n208 VTAIL.n207 6.59444
R786 VTAIL.n208 VTAIL.n172 6.59444
R787 VTAIL.n525 VTAIL.n489 6.59444
R788 VTAIL.n525 VTAIL.n524 6.59444
R789 VTAIL.n445 VTAIL.n409 6.59444
R790 VTAIL.n445 VTAIL.n444 6.59444
R791 VTAIL.n367 VTAIL.n331 6.59444
R792 VTAIL.n367 VTAIL.n366 6.59444
R793 VTAIL.n287 VTAIL.n251 6.59444
R794 VTAIL.n287 VTAIL.n286 6.59444
R795 VTAIL.n598 VTAIL.n568 5.81868
R796 VTAIL.n606 VTAIL.n605 5.81868
R797 VTAIL.n46 VTAIL.n16 5.81868
R798 VTAIL.n54 VTAIL.n53 5.81868
R799 VTAIL.n124 VTAIL.n94 5.81868
R800 VTAIL.n132 VTAIL.n131 5.81868
R801 VTAIL.n204 VTAIL.n174 5.81868
R802 VTAIL.n212 VTAIL.n211 5.81868
R803 VTAIL.n529 VTAIL.n528 5.81868
R804 VTAIL.n521 VTAIL.n491 5.81868
R805 VTAIL.n449 VTAIL.n448 5.81868
R806 VTAIL.n441 VTAIL.n411 5.81868
R807 VTAIL.n371 VTAIL.n370 5.81868
R808 VTAIL.n363 VTAIL.n333 5.81868
R809 VTAIL.n291 VTAIL.n290 5.81868
R810 VTAIL.n283 VTAIL.n253 5.81868
R811 VTAIL.n597 VTAIL.n570 5.04292
R812 VTAIL.n609 VTAIL.n564 5.04292
R813 VTAIL.n45 VTAIL.n18 5.04292
R814 VTAIL.n57 VTAIL.n12 5.04292
R815 VTAIL.n123 VTAIL.n96 5.04292
R816 VTAIL.n135 VTAIL.n90 5.04292
R817 VTAIL.n203 VTAIL.n176 5.04292
R818 VTAIL.n215 VTAIL.n170 5.04292
R819 VTAIL.n532 VTAIL.n487 5.04292
R820 VTAIL.n520 VTAIL.n493 5.04292
R821 VTAIL.n452 VTAIL.n407 5.04292
R822 VTAIL.n440 VTAIL.n413 5.04292
R823 VTAIL.n374 VTAIL.n329 5.04292
R824 VTAIL.n362 VTAIL.n335 5.04292
R825 VTAIL.n294 VTAIL.n249 5.04292
R826 VTAIL.n282 VTAIL.n255 5.04292
R827 VTAIL.n594 VTAIL.n593 4.26717
R828 VTAIL.n610 VTAIL.n562 4.26717
R829 VTAIL.n42 VTAIL.n41 4.26717
R830 VTAIL.n58 VTAIL.n10 4.26717
R831 VTAIL.n120 VTAIL.n119 4.26717
R832 VTAIL.n136 VTAIL.n88 4.26717
R833 VTAIL.n200 VTAIL.n199 4.26717
R834 VTAIL.n216 VTAIL.n168 4.26717
R835 VTAIL.n533 VTAIL.n485 4.26717
R836 VTAIL.n517 VTAIL.n516 4.26717
R837 VTAIL.n453 VTAIL.n405 4.26717
R838 VTAIL.n437 VTAIL.n436 4.26717
R839 VTAIL.n375 VTAIL.n327 4.26717
R840 VTAIL.n359 VTAIL.n358 4.26717
R841 VTAIL.n295 VTAIL.n247 4.26717
R842 VTAIL.n279 VTAIL.n278 4.26717
R843 VTAIL.n580 VTAIL.n579 3.70982
R844 VTAIL.n28 VTAIL.n27 3.70982
R845 VTAIL.n106 VTAIL.n105 3.70982
R846 VTAIL.n186 VTAIL.n185 3.70982
R847 VTAIL.n503 VTAIL.n502 3.70982
R848 VTAIL.n423 VTAIL.n422 3.70982
R849 VTAIL.n345 VTAIL.n344 3.70982
R850 VTAIL.n265 VTAIL.n264 3.70982
R851 VTAIL.n317 VTAIL.n315 3.56084
R852 VTAIL.n395 VTAIL.n317 3.56084
R853 VTAIL.n475 VTAIL.n473 3.56084
R854 VTAIL.n553 VTAIL.n475 3.56084
R855 VTAIL.n237 VTAIL.n159 3.56084
R856 VTAIL.n159 VTAIL.n157 3.56084
R857 VTAIL.n79 VTAIL.n1 3.56084
R858 VTAIL VTAIL.n631 3.50266
R859 VTAIL.n590 VTAIL.n572 3.49141
R860 VTAIL.n614 VTAIL.n613 3.49141
R861 VTAIL.n38 VTAIL.n20 3.49141
R862 VTAIL.n62 VTAIL.n61 3.49141
R863 VTAIL.n116 VTAIL.n98 3.49141
R864 VTAIL.n140 VTAIL.n139 3.49141
R865 VTAIL.n196 VTAIL.n178 3.49141
R866 VTAIL.n220 VTAIL.n219 3.49141
R867 VTAIL.n537 VTAIL.n536 3.49141
R868 VTAIL.n513 VTAIL.n495 3.49141
R869 VTAIL.n457 VTAIL.n456 3.49141
R870 VTAIL.n433 VTAIL.n415 3.49141
R871 VTAIL.n379 VTAIL.n378 3.49141
R872 VTAIL.n355 VTAIL.n337 3.49141
R873 VTAIL.n299 VTAIL.n298 3.49141
R874 VTAIL.n275 VTAIL.n257 3.49141
R875 VTAIL.n589 VTAIL.n574 2.71565
R876 VTAIL.n617 VTAIL.n560 2.71565
R877 VTAIL.n37 VTAIL.n22 2.71565
R878 VTAIL.n65 VTAIL.n8 2.71565
R879 VTAIL.n115 VTAIL.n100 2.71565
R880 VTAIL.n143 VTAIL.n86 2.71565
R881 VTAIL.n195 VTAIL.n180 2.71565
R882 VTAIL.n223 VTAIL.n166 2.71565
R883 VTAIL.n540 VTAIL.n483 2.71565
R884 VTAIL.n512 VTAIL.n497 2.71565
R885 VTAIL.n460 VTAIL.n403 2.71565
R886 VTAIL.n432 VTAIL.n417 2.71565
R887 VTAIL.n382 VTAIL.n325 2.71565
R888 VTAIL.n354 VTAIL.n339 2.71565
R889 VTAIL.n302 VTAIL.n245 2.71565
R890 VTAIL.n274 VTAIL.n259 2.71565
R891 VTAIL.n0 VTAIL.t2 2.30092
R892 VTAIL.n0 VTAIL.t3 2.30092
R893 VTAIL.n158 VTAIL.t8 2.30092
R894 VTAIL.n158 VTAIL.t10 2.30092
R895 VTAIL.n474 VTAIL.t14 2.30092
R896 VTAIL.n474 VTAIL.t15 2.30092
R897 VTAIL.n316 VTAIL.t4 2.30092
R898 VTAIL.n316 VTAIL.t0 2.30092
R899 VTAIL.n586 VTAIL.n585 1.93989
R900 VTAIL.n618 VTAIL.n558 1.93989
R901 VTAIL.n34 VTAIL.n33 1.93989
R902 VTAIL.n66 VTAIL.n6 1.93989
R903 VTAIL.n112 VTAIL.n111 1.93989
R904 VTAIL.n144 VTAIL.n84 1.93989
R905 VTAIL.n192 VTAIL.n191 1.93989
R906 VTAIL.n224 VTAIL.n164 1.93989
R907 VTAIL.n541 VTAIL.n481 1.93989
R908 VTAIL.n509 VTAIL.n508 1.93989
R909 VTAIL.n461 VTAIL.n401 1.93989
R910 VTAIL.n429 VTAIL.n428 1.93989
R911 VTAIL.n383 VTAIL.n323 1.93989
R912 VTAIL.n351 VTAIL.n350 1.93989
R913 VTAIL.n303 VTAIL.n243 1.93989
R914 VTAIL.n271 VTAIL.n270 1.93989
R915 VTAIL.n582 VTAIL.n576 1.16414
R916 VTAIL.n623 VTAIL.n621 1.16414
R917 VTAIL.n630 VTAIL.n554 1.16414
R918 VTAIL.n30 VTAIL.n24 1.16414
R919 VTAIL.n71 VTAIL.n69 1.16414
R920 VTAIL.n78 VTAIL.n2 1.16414
R921 VTAIL.n108 VTAIL.n102 1.16414
R922 VTAIL.n149 VTAIL.n147 1.16414
R923 VTAIL.n156 VTAIL.n80 1.16414
R924 VTAIL.n188 VTAIL.n182 1.16414
R925 VTAIL.n229 VTAIL.n227 1.16414
R926 VTAIL.n236 VTAIL.n160 1.16414
R927 VTAIL.n552 VTAIL.n476 1.16414
R928 VTAIL.n545 VTAIL.n544 1.16414
R929 VTAIL.n505 VTAIL.n499 1.16414
R930 VTAIL.n472 VTAIL.n396 1.16414
R931 VTAIL.n465 VTAIL.n464 1.16414
R932 VTAIL.n425 VTAIL.n419 1.16414
R933 VTAIL.n394 VTAIL.n318 1.16414
R934 VTAIL.n387 VTAIL.n386 1.16414
R935 VTAIL.n347 VTAIL.n341 1.16414
R936 VTAIL.n314 VTAIL.n238 1.16414
R937 VTAIL.n307 VTAIL.n306 1.16414
R938 VTAIL.n267 VTAIL.n261 1.16414
R939 VTAIL.n473 VTAIL.n395 0.470328
R940 VTAIL.n157 VTAIL.n79 0.470328
R941 VTAIL.n581 VTAIL.n578 0.388379
R942 VTAIL.n622 VTAIL.n556 0.388379
R943 VTAIL.n628 VTAIL.n627 0.388379
R944 VTAIL.n29 VTAIL.n26 0.388379
R945 VTAIL.n70 VTAIL.n4 0.388379
R946 VTAIL.n76 VTAIL.n75 0.388379
R947 VTAIL.n107 VTAIL.n104 0.388379
R948 VTAIL.n148 VTAIL.n82 0.388379
R949 VTAIL.n154 VTAIL.n153 0.388379
R950 VTAIL.n187 VTAIL.n184 0.388379
R951 VTAIL.n228 VTAIL.n162 0.388379
R952 VTAIL.n234 VTAIL.n233 0.388379
R953 VTAIL.n550 VTAIL.n549 0.388379
R954 VTAIL.n480 VTAIL.n478 0.388379
R955 VTAIL.n504 VTAIL.n501 0.388379
R956 VTAIL.n470 VTAIL.n469 0.388379
R957 VTAIL.n400 VTAIL.n398 0.388379
R958 VTAIL.n424 VTAIL.n421 0.388379
R959 VTAIL.n392 VTAIL.n391 0.388379
R960 VTAIL.n322 VTAIL.n320 0.388379
R961 VTAIL.n346 VTAIL.n343 0.388379
R962 VTAIL.n312 VTAIL.n311 0.388379
R963 VTAIL.n242 VTAIL.n240 0.388379
R964 VTAIL.n266 VTAIL.n263 0.388379
R965 VTAIL.n580 VTAIL.n575 0.155672
R966 VTAIL.n587 VTAIL.n575 0.155672
R967 VTAIL.n588 VTAIL.n587 0.155672
R968 VTAIL.n588 VTAIL.n571 0.155672
R969 VTAIL.n595 VTAIL.n571 0.155672
R970 VTAIL.n596 VTAIL.n595 0.155672
R971 VTAIL.n596 VTAIL.n567 0.155672
R972 VTAIL.n603 VTAIL.n567 0.155672
R973 VTAIL.n604 VTAIL.n603 0.155672
R974 VTAIL.n604 VTAIL.n563 0.155672
R975 VTAIL.n611 VTAIL.n563 0.155672
R976 VTAIL.n612 VTAIL.n611 0.155672
R977 VTAIL.n612 VTAIL.n559 0.155672
R978 VTAIL.n619 VTAIL.n559 0.155672
R979 VTAIL.n620 VTAIL.n619 0.155672
R980 VTAIL.n620 VTAIL.n555 0.155672
R981 VTAIL.n629 VTAIL.n555 0.155672
R982 VTAIL.n28 VTAIL.n23 0.155672
R983 VTAIL.n35 VTAIL.n23 0.155672
R984 VTAIL.n36 VTAIL.n35 0.155672
R985 VTAIL.n36 VTAIL.n19 0.155672
R986 VTAIL.n43 VTAIL.n19 0.155672
R987 VTAIL.n44 VTAIL.n43 0.155672
R988 VTAIL.n44 VTAIL.n15 0.155672
R989 VTAIL.n51 VTAIL.n15 0.155672
R990 VTAIL.n52 VTAIL.n51 0.155672
R991 VTAIL.n52 VTAIL.n11 0.155672
R992 VTAIL.n59 VTAIL.n11 0.155672
R993 VTAIL.n60 VTAIL.n59 0.155672
R994 VTAIL.n60 VTAIL.n7 0.155672
R995 VTAIL.n67 VTAIL.n7 0.155672
R996 VTAIL.n68 VTAIL.n67 0.155672
R997 VTAIL.n68 VTAIL.n3 0.155672
R998 VTAIL.n77 VTAIL.n3 0.155672
R999 VTAIL.n106 VTAIL.n101 0.155672
R1000 VTAIL.n113 VTAIL.n101 0.155672
R1001 VTAIL.n114 VTAIL.n113 0.155672
R1002 VTAIL.n114 VTAIL.n97 0.155672
R1003 VTAIL.n121 VTAIL.n97 0.155672
R1004 VTAIL.n122 VTAIL.n121 0.155672
R1005 VTAIL.n122 VTAIL.n93 0.155672
R1006 VTAIL.n129 VTAIL.n93 0.155672
R1007 VTAIL.n130 VTAIL.n129 0.155672
R1008 VTAIL.n130 VTAIL.n89 0.155672
R1009 VTAIL.n137 VTAIL.n89 0.155672
R1010 VTAIL.n138 VTAIL.n137 0.155672
R1011 VTAIL.n138 VTAIL.n85 0.155672
R1012 VTAIL.n145 VTAIL.n85 0.155672
R1013 VTAIL.n146 VTAIL.n145 0.155672
R1014 VTAIL.n146 VTAIL.n81 0.155672
R1015 VTAIL.n155 VTAIL.n81 0.155672
R1016 VTAIL.n186 VTAIL.n181 0.155672
R1017 VTAIL.n193 VTAIL.n181 0.155672
R1018 VTAIL.n194 VTAIL.n193 0.155672
R1019 VTAIL.n194 VTAIL.n177 0.155672
R1020 VTAIL.n201 VTAIL.n177 0.155672
R1021 VTAIL.n202 VTAIL.n201 0.155672
R1022 VTAIL.n202 VTAIL.n173 0.155672
R1023 VTAIL.n209 VTAIL.n173 0.155672
R1024 VTAIL.n210 VTAIL.n209 0.155672
R1025 VTAIL.n210 VTAIL.n169 0.155672
R1026 VTAIL.n217 VTAIL.n169 0.155672
R1027 VTAIL.n218 VTAIL.n217 0.155672
R1028 VTAIL.n218 VTAIL.n165 0.155672
R1029 VTAIL.n225 VTAIL.n165 0.155672
R1030 VTAIL.n226 VTAIL.n225 0.155672
R1031 VTAIL.n226 VTAIL.n161 0.155672
R1032 VTAIL.n235 VTAIL.n161 0.155672
R1033 VTAIL.n551 VTAIL.n477 0.155672
R1034 VTAIL.n543 VTAIL.n477 0.155672
R1035 VTAIL.n543 VTAIL.n542 0.155672
R1036 VTAIL.n542 VTAIL.n482 0.155672
R1037 VTAIL.n535 VTAIL.n482 0.155672
R1038 VTAIL.n535 VTAIL.n534 0.155672
R1039 VTAIL.n534 VTAIL.n486 0.155672
R1040 VTAIL.n527 VTAIL.n486 0.155672
R1041 VTAIL.n527 VTAIL.n526 0.155672
R1042 VTAIL.n526 VTAIL.n490 0.155672
R1043 VTAIL.n519 VTAIL.n490 0.155672
R1044 VTAIL.n519 VTAIL.n518 0.155672
R1045 VTAIL.n518 VTAIL.n494 0.155672
R1046 VTAIL.n511 VTAIL.n494 0.155672
R1047 VTAIL.n511 VTAIL.n510 0.155672
R1048 VTAIL.n510 VTAIL.n498 0.155672
R1049 VTAIL.n503 VTAIL.n498 0.155672
R1050 VTAIL.n471 VTAIL.n397 0.155672
R1051 VTAIL.n463 VTAIL.n397 0.155672
R1052 VTAIL.n463 VTAIL.n462 0.155672
R1053 VTAIL.n462 VTAIL.n402 0.155672
R1054 VTAIL.n455 VTAIL.n402 0.155672
R1055 VTAIL.n455 VTAIL.n454 0.155672
R1056 VTAIL.n454 VTAIL.n406 0.155672
R1057 VTAIL.n447 VTAIL.n406 0.155672
R1058 VTAIL.n447 VTAIL.n446 0.155672
R1059 VTAIL.n446 VTAIL.n410 0.155672
R1060 VTAIL.n439 VTAIL.n410 0.155672
R1061 VTAIL.n439 VTAIL.n438 0.155672
R1062 VTAIL.n438 VTAIL.n414 0.155672
R1063 VTAIL.n431 VTAIL.n414 0.155672
R1064 VTAIL.n431 VTAIL.n430 0.155672
R1065 VTAIL.n430 VTAIL.n418 0.155672
R1066 VTAIL.n423 VTAIL.n418 0.155672
R1067 VTAIL.n393 VTAIL.n319 0.155672
R1068 VTAIL.n385 VTAIL.n319 0.155672
R1069 VTAIL.n385 VTAIL.n384 0.155672
R1070 VTAIL.n384 VTAIL.n324 0.155672
R1071 VTAIL.n377 VTAIL.n324 0.155672
R1072 VTAIL.n377 VTAIL.n376 0.155672
R1073 VTAIL.n376 VTAIL.n328 0.155672
R1074 VTAIL.n369 VTAIL.n328 0.155672
R1075 VTAIL.n369 VTAIL.n368 0.155672
R1076 VTAIL.n368 VTAIL.n332 0.155672
R1077 VTAIL.n361 VTAIL.n332 0.155672
R1078 VTAIL.n361 VTAIL.n360 0.155672
R1079 VTAIL.n360 VTAIL.n336 0.155672
R1080 VTAIL.n353 VTAIL.n336 0.155672
R1081 VTAIL.n353 VTAIL.n352 0.155672
R1082 VTAIL.n352 VTAIL.n340 0.155672
R1083 VTAIL.n345 VTAIL.n340 0.155672
R1084 VTAIL.n313 VTAIL.n239 0.155672
R1085 VTAIL.n305 VTAIL.n239 0.155672
R1086 VTAIL.n305 VTAIL.n304 0.155672
R1087 VTAIL.n304 VTAIL.n244 0.155672
R1088 VTAIL.n297 VTAIL.n244 0.155672
R1089 VTAIL.n297 VTAIL.n296 0.155672
R1090 VTAIL.n296 VTAIL.n248 0.155672
R1091 VTAIL.n289 VTAIL.n248 0.155672
R1092 VTAIL.n289 VTAIL.n288 0.155672
R1093 VTAIL.n288 VTAIL.n252 0.155672
R1094 VTAIL.n281 VTAIL.n252 0.155672
R1095 VTAIL.n281 VTAIL.n280 0.155672
R1096 VTAIL.n280 VTAIL.n256 0.155672
R1097 VTAIL.n273 VTAIL.n256 0.155672
R1098 VTAIL.n273 VTAIL.n272 0.155672
R1099 VTAIL.n272 VTAIL.n260 0.155672
R1100 VTAIL.n265 VTAIL.n260 0.155672
R1101 VTAIL VTAIL.n1 0.0586897
R1102 VDD1 VDD1.n0 77.2454
R1103 VDD1.n3 VDD1.n2 77.1317
R1104 VDD1.n3 VDD1.n1 77.1317
R1105 VDD1.n5 VDD1.n4 75.4068
R1106 VDD1.n5 VDD1.n3 52.5009
R1107 VDD1.n4 VDD1.t3 2.30092
R1108 VDD1.n4 VDD1.t4 2.30092
R1109 VDD1.n0 VDD1.t2 2.30092
R1110 VDD1.n0 VDD1.t7 2.30092
R1111 VDD1.n2 VDD1.t1 2.30092
R1112 VDD1.n2 VDD1.t0 2.30092
R1113 VDD1.n1 VDD1.t6 2.30092
R1114 VDD1.n1 VDD1.t5 2.30092
R1115 VDD1 VDD1.n5 1.72248
R1116 VN.n71 VN.n37 161.3
R1117 VN.n70 VN.n69 161.3
R1118 VN.n68 VN.n38 161.3
R1119 VN.n67 VN.n66 161.3
R1120 VN.n65 VN.n39 161.3
R1121 VN.n64 VN.n63 161.3
R1122 VN.n62 VN.n40 161.3
R1123 VN.n61 VN.n60 161.3
R1124 VN.n58 VN.n41 161.3
R1125 VN.n57 VN.n56 161.3
R1126 VN.n55 VN.n42 161.3
R1127 VN.n54 VN.n53 161.3
R1128 VN.n52 VN.n43 161.3
R1129 VN.n51 VN.n50 161.3
R1130 VN.n49 VN.n44 161.3
R1131 VN.n48 VN.n47 161.3
R1132 VN.n34 VN.n0 161.3
R1133 VN.n33 VN.n32 161.3
R1134 VN.n31 VN.n1 161.3
R1135 VN.n30 VN.n29 161.3
R1136 VN.n28 VN.n2 161.3
R1137 VN.n27 VN.n26 161.3
R1138 VN.n25 VN.n3 161.3
R1139 VN.n24 VN.n23 161.3
R1140 VN.n21 VN.n4 161.3
R1141 VN.n20 VN.n19 161.3
R1142 VN.n18 VN.n5 161.3
R1143 VN.n17 VN.n16 161.3
R1144 VN.n15 VN.n6 161.3
R1145 VN.n14 VN.n13 161.3
R1146 VN.n12 VN.n7 161.3
R1147 VN.n11 VN.n10 161.3
R1148 VN.n8 VN.t3 121.847
R1149 VN.n45 VN.t1 121.847
R1150 VN.n9 VN.t2 89.6144
R1151 VN.n22 VN.t0 89.6144
R1152 VN.n35 VN.t7 89.6144
R1153 VN.n46 VN.t4 89.6144
R1154 VN.n59 VN.t5 89.6144
R1155 VN.n72 VN.t6 89.6144
R1156 VN.n36 VN.n35 60.4062
R1157 VN.n73 VN.n72 60.4062
R1158 VN.n9 VN.n8 59.6416
R1159 VN.n46 VN.n45 59.6416
R1160 VN VN.n73 58.3829
R1161 VN.n16 VN.n15 56.5193
R1162 VN.n53 VN.n52 56.5193
R1163 VN.n29 VN.n28 52.1486
R1164 VN.n66 VN.n65 52.1486
R1165 VN.n29 VN.n1 28.8382
R1166 VN.n66 VN.n38 28.8382
R1167 VN.n10 VN.n7 24.4675
R1168 VN.n14 VN.n7 24.4675
R1169 VN.n15 VN.n14 24.4675
R1170 VN.n16 VN.n5 24.4675
R1171 VN.n20 VN.n5 24.4675
R1172 VN.n21 VN.n20 24.4675
R1173 VN.n23 VN.n3 24.4675
R1174 VN.n27 VN.n3 24.4675
R1175 VN.n28 VN.n27 24.4675
R1176 VN.n33 VN.n1 24.4675
R1177 VN.n34 VN.n33 24.4675
R1178 VN.n52 VN.n51 24.4675
R1179 VN.n51 VN.n44 24.4675
R1180 VN.n47 VN.n44 24.4675
R1181 VN.n65 VN.n64 24.4675
R1182 VN.n64 VN.n40 24.4675
R1183 VN.n60 VN.n40 24.4675
R1184 VN.n58 VN.n57 24.4675
R1185 VN.n57 VN.n42 24.4675
R1186 VN.n53 VN.n42 24.4675
R1187 VN.n71 VN.n70 24.4675
R1188 VN.n70 VN.n38 24.4675
R1189 VN.n35 VN.n34 21.7761
R1190 VN.n72 VN.n71 21.7761
R1191 VN.n10 VN.n9 15.4147
R1192 VN.n22 VN.n21 15.4147
R1193 VN.n47 VN.n46 15.4147
R1194 VN.n59 VN.n58 15.4147
R1195 VN.n23 VN.n22 9.05329
R1196 VN.n60 VN.n59 9.05329
R1197 VN.n48 VN.n45 2.62604
R1198 VN.n11 VN.n8 2.62604
R1199 VN.n73 VN.n37 0.417535
R1200 VN.n36 VN.n0 0.417535
R1201 VN VN.n36 0.394291
R1202 VN.n69 VN.n37 0.189894
R1203 VN.n69 VN.n68 0.189894
R1204 VN.n68 VN.n67 0.189894
R1205 VN.n67 VN.n39 0.189894
R1206 VN.n63 VN.n39 0.189894
R1207 VN.n63 VN.n62 0.189894
R1208 VN.n62 VN.n61 0.189894
R1209 VN.n61 VN.n41 0.189894
R1210 VN.n56 VN.n41 0.189894
R1211 VN.n56 VN.n55 0.189894
R1212 VN.n55 VN.n54 0.189894
R1213 VN.n54 VN.n43 0.189894
R1214 VN.n50 VN.n43 0.189894
R1215 VN.n50 VN.n49 0.189894
R1216 VN.n49 VN.n48 0.189894
R1217 VN.n12 VN.n11 0.189894
R1218 VN.n13 VN.n12 0.189894
R1219 VN.n13 VN.n6 0.189894
R1220 VN.n17 VN.n6 0.189894
R1221 VN.n18 VN.n17 0.189894
R1222 VN.n19 VN.n18 0.189894
R1223 VN.n19 VN.n4 0.189894
R1224 VN.n24 VN.n4 0.189894
R1225 VN.n25 VN.n24 0.189894
R1226 VN.n26 VN.n25 0.189894
R1227 VN.n26 VN.n2 0.189894
R1228 VN.n30 VN.n2 0.189894
R1229 VN.n31 VN.n30 0.189894
R1230 VN.n32 VN.n31 0.189894
R1231 VN.n32 VN.n0 0.189894
R1232 VDD2.n2 VDD2.n1 77.1317
R1233 VDD2.n2 VDD2.n0 77.1317
R1234 VDD2 VDD2.n5 77.1288
R1235 VDD2.n4 VDD2.n3 75.407
R1236 VDD2.n4 VDD2.n2 51.9179
R1237 VDD2.n5 VDD2.t3 2.30092
R1238 VDD2.n5 VDD2.t6 2.30092
R1239 VDD2.n3 VDD2.t1 2.30092
R1240 VDD2.n3 VDD2.t2 2.30092
R1241 VDD2.n1 VDD2.t7 2.30092
R1242 VDD2.n1 VDD2.t0 2.30092
R1243 VDD2.n0 VDD2.t4 2.30092
R1244 VDD2.n0 VDD2.t5 2.30092
R1245 VDD2 VDD2.n4 1.83886
R1246 B.n725 B.n724 585
R1247 B.n726 B.n93 585
R1248 B.n728 B.n727 585
R1249 B.n729 B.n92 585
R1250 B.n731 B.n730 585
R1251 B.n732 B.n91 585
R1252 B.n734 B.n733 585
R1253 B.n735 B.n90 585
R1254 B.n737 B.n736 585
R1255 B.n738 B.n89 585
R1256 B.n740 B.n739 585
R1257 B.n741 B.n88 585
R1258 B.n743 B.n742 585
R1259 B.n744 B.n87 585
R1260 B.n746 B.n745 585
R1261 B.n747 B.n86 585
R1262 B.n749 B.n748 585
R1263 B.n750 B.n85 585
R1264 B.n752 B.n751 585
R1265 B.n753 B.n84 585
R1266 B.n755 B.n754 585
R1267 B.n756 B.n83 585
R1268 B.n758 B.n757 585
R1269 B.n759 B.n82 585
R1270 B.n761 B.n760 585
R1271 B.n762 B.n81 585
R1272 B.n764 B.n763 585
R1273 B.n765 B.n80 585
R1274 B.n767 B.n766 585
R1275 B.n768 B.n79 585
R1276 B.n770 B.n769 585
R1277 B.n771 B.n78 585
R1278 B.n773 B.n772 585
R1279 B.n774 B.n77 585
R1280 B.n776 B.n775 585
R1281 B.n777 B.n76 585
R1282 B.n779 B.n778 585
R1283 B.n780 B.n75 585
R1284 B.n782 B.n781 585
R1285 B.n783 B.n74 585
R1286 B.n785 B.n784 585
R1287 B.n786 B.n73 585
R1288 B.n788 B.n787 585
R1289 B.n789 B.n72 585
R1290 B.n791 B.n790 585
R1291 B.n792 B.n71 585
R1292 B.n794 B.n793 585
R1293 B.n795 B.n68 585
R1294 B.n798 B.n797 585
R1295 B.n799 B.n67 585
R1296 B.n801 B.n800 585
R1297 B.n802 B.n66 585
R1298 B.n804 B.n803 585
R1299 B.n805 B.n65 585
R1300 B.n807 B.n806 585
R1301 B.n808 B.n61 585
R1302 B.n810 B.n809 585
R1303 B.n811 B.n60 585
R1304 B.n813 B.n812 585
R1305 B.n814 B.n59 585
R1306 B.n816 B.n815 585
R1307 B.n817 B.n58 585
R1308 B.n819 B.n818 585
R1309 B.n820 B.n57 585
R1310 B.n822 B.n821 585
R1311 B.n823 B.n56 585
R1312 B.n825 B.n824 585
R1313 B.n826 B.n55 585
R1314 B.n828 B.n827 585
R1315 B.n829 B.n54 585
R1316 B.n831 B.n830 585
R1317 B.n832 B.n53 585
R1318 B.n834 B.n833 585
R1319 B.n835 B.n52 585
R1320 B.n837 B.n836 585
R1321 B.n838 B.n51 585
R1322 B.n840 B.n839 585
R1323 B.n841 B.n50 585
R1324 B.n843 B.n842 585
R1325 B.n844 B.n49 585
R1326 B.n846 B.n845 585
R1327 B.n847 B.n48 585
R1328 B.n849 B.n848 585
R1329 B.n850 B.n47 585
R1330 B.n852 B.n851 585
R1331 B.n853 B.n46 585
R1332 B.n855 B.n854 585
R1333 B.n856 B.n45 585
R1334 B.n858 B.n857 585
R1335 B.n859 B.n44 585
R1336 B.n861 B.n860 585
R1337 B.n862 B.n43 585
R1338 B.n864 B.n863 585
R1339 B.n865 B.n42 585
R1340 B.n867 B.n866 585
R1341 B.n868 B.n41 585
R1342 B.n870 B.n869 585
R1343 B.n871 B.n40 585
R1344 B.n873 B.n872 585
R1345 B.n874 B.n39 585
R1346 B.n876 B.n875 585
R1347 B.n877 B.n38 585
R1348 B.n879 B.n878 585
R1349 B.n880 B.n37 585
R1350 B.n882 B.n881 585
R1351 B.n723 B.n94 585
R1352 B.n722 B.n721 585
R1353 B.n720 B.n95 585
R1354 B.n719 B.n718 585
R1355 B.n717 B.n96 585
R1356 B.n716 B.n715 585
R1357 B.n714 B.n97 585
R1358 B.n713 B.n712 585
R1359 B.n711 B.n98 585
R1360 B.n710 B.n709 585
R1361 B.n708 B.n99 585
R1362 B.n707 B.n706 585
R1363 B.n705 B.n100 585
R1364 B.n704 B.n703 585
R1365 B.n702 B.n101 585
R1366 B.n701 B.n700 585
R1367 B.n699 B.n102 585
R1368 B.n698 B.n697 585
R1369 B.n696 B.n103 585
R1370 B.n695 B.n694 585
R1371 B.n693 B.n104 585
R1372 B.n692 B.n691 585
R1373 B.n690 B.n105 585
R1374 B.n689 B.n688 585
R1375 B.n687 B.n106 585
R1376 B.n686 B.n685 585
R1377 B.n684 B.n107 585
R1378 B.n683 B.n682 585
R1379 B.n681 B.n108 585
R1380 B.n680 B.n679 585
R1381 B.n678 B.n109 585
R1382 B.n677 B.n676 585
R1383 B.n675 B.n110 585
R1384 B.n674 B.n673 585
R1385 B.n672 B.n111 585
R1386 B.n671 B.n670 585
R1387 B.n669 B.n112 585
R1388 B.n668 B.n667 585
R1389 B.n666 B.n113 585
R1390 B.n665 B.n664 585
R1391 B.n663 B.n114 585
R1392 B.n662 B.n661 585
R1393 B.n660 B.n115 585
R1394 B.n659 B.n658 585
R1395 B.n657 B.n116 585
R1396 B.n656 B.n655 585
R1397 B.n654 B.n117 585
R1398 B.n653 B.n652 585
R1399 B.n651 B.n118 585
R1400 B.n650 B.n649 585
R1401 B.n648 B.n119 585
R1402 B.n647 B.n646 585
R1403 B.n645 B.n120 585
R1404 B.n644 B.n643 585
R1405 B.n642 B.n121 585
R1406 B.n641 B.n640 585
R1407 B.n639 B.n122 585
R1408 B.n638 B.n637 585
R1409 B.n636 B.n123 585
R1410 B.n635 B.n634 585
R1411 B.n633 B.n124 585
R1412 B.n632 B.n631 585
R1413 B.n630 B.n125 585
R1414 B.n629 B.n628 585
R1415 B.n627 B.n126 585
R1416 B.n626 B.n625 585
R1417 B.n624 B.n127 585
R1418 B.n623 B.n622 585
R1419 B.n621 B.n128 585
R1420 B.n620 B.n619 585
R1421 B.n618 B.n129 585
R1422 B.n617 B.n616 585
R1423 B.n615 B.n130 585
R1424 B.n614 B.n613 585
R1425 B.n612 B.n131 585
R1426 B.n611 B.n610 585
R1427 B.n609 B.n132 585
R1428 B.n608 B.n607 585
R1429 B.n606 B.n133 585
R1430 B.n605 B.n604 585
R1431 B.n603 B.n134 585
R1432 B.n602 B.n601 585
R1433 B.n600 B.n135 585
R1434 B.n599 B.n598 585
R1435 B.n597 B.n136 585
R1436 B.n596 B.n595 585
R1437 B.n594 B.n137 585
R1438 B.n593 B.n592 585
R1439 B.n591 B.n138 585
R1440 B.n590 B.n589 585
R1441 B.n588 B.n139 585
R1442 B.n587 B.n586 585
R1443 B.n585 B.n140 585
R1444 B.n584 B.n583 585
R1445 B.n582 B.n141 585
R1446 B.n581 B.n580 585
R1447 B.n579 B.n142 585
R1448 B.n578 B.n577 585
R1449 B.n576 B.n143 585
R1450 B.n575 B.n574 585
R1451 B.n573 B.n144 585
R1452 B.n572 B.n571 585
R1453 B.n570 B.n145 585
R1454 B.n569 B.n568 585
R1455 B.n567 B.n146 585
R1456 B.n566 B.n565 585
R1457 B.n564 B.n147 585
R1458 B.n563 B.n562 585
R1459 B.n561 B.n148 585
R1460 B.n560 B.n559 585
R1461 B.n558 B.n149 585
R1462 B.n557 B.n556 585
R1463 B.n555 B.n150 585
R1464 B.n554 B.n553 585
R1465 B.n552 B.n151 585
R1466 B.n551 B.n550 585
R1467 B.n549 B.n152 585
R1468 B.n548 B.n547 585
R1469 B.n546 B.n153 585
R1470 B.n545 B.n544 585
R1471 B.n543 B.n154 585
R1472 B.n542 B.n541 585
R1473 B.n540 B.n155 585
R1474 B.n539 B.n538 585
R1475 B.n537 B.n156 585
R1476 B.n536 B.n535 585
R1477 B.n534 B.n157 585
R1478 B.n533 B.n532 585
R1479 B.n531 B.n158 585
R1480 B.n530 B.n529 585
R1481 B.n528 B.n159 585
R1482 B.n527 B.n526 585
R1483 B.n525 B.n160 585
R1484 B.n524 B.n523 585
R1485 B.n522 B.n161 585
R1486 B.n521 B.n520 585
R1487 B.n519 B.n162 585
R1488 B.n518 B.n517 585
R1489 B.n516 B.n163 585
R1490 B.n355 B.n354 585
R1491 B.n356 B.n217 585
R1492 B.n358 B.n357 585
R1493 B.n359 B.n216 585
R1494 B.n361 B.n360 585
R1495 B.n362 B.n215 585
R1496 B.n364 B.n363 585
R1497 B.n365 B.n214 585
R1498 B.n367 B.n366 585
R1499 B.n368 B.n213 585
R1500 B.n370 B.n369 585
R1501 B.n371 B.n212 585
R1502 B.n373 B.n372 585
R1503 B.n374 B.n211 585
R1504 B.n376 B.n375 585
R1505 B.n377 B.n210 585
R1506 B.n379 B.n378 585
R1507 B.n380 B.n209 585
R1508 B.n382 B.n381 585
R1509 B.n383 B.n208 585
R1510 B.n385 B.n384 585
R1511 B.n386 B.n207 585
R1512 B.n388 B.n387 585
R1513 B.n389 B.n206 585
R1514 B.n391 B.n390 585
R1515 B.n392 B.n205 585
R1516 B.n394 B.n393 585
R1517 B.n395 B.n204 585
R1518 B.n397 B.n396 585
R1519 B.n398 B.n203 585
R1520 B.n400 B.n399 585
R1521 B.n401 B.n202 585
R1522 B.n403 B.n402 585
R1523 B.n404 B.n201 585
R1524 B.n406 B.n405 585
R1525 B.n407 B.n200 585
R1526 B.n409 B.n408 585
R1527 B.n410 B.n199 585
R1528 B.n412 B.n411 585
R1529 B.n413 B.n198 585
R1530 B.n415 B.n414 585
R1531 B.n416 B.n197 585
R1532 B.n418 B.n417 585
R1533 B.n419 B.n196 585
R1534 B.n421 B.n420 585
R1535 B.n422 B.n195 585
R1536 B.n424 B.n423 585
R1537 B.n425 B.n192 585
R1538 B.n428 B.n427 585
R1539 B.n429 B.n191 585
R1540 B.n431 B.n430 585
R1541 B.n432 B.n190 585
R1542 B.n434 B.n433 585
R1543 B.n435 B.n189 585
R1544 B.n437 B.n436 585
R1545 B.n438 B.n188 585
R1546 B.n443 B.n442 585
R1547 B.n444 B.n187 585
R1548 B.n446 B.n445 585
R1549 B.n447 B.n186 585
R1550 B.n449 B.n448 585
R1551 B.n450 B.n185 585
R1552 B.n452 B.n451 585
R1553 B.n453 B.n184 585
R1554 B.n455 B.n454 585
R1555 B.n456 B.n183 585
R1556 B.n458 B.n457 585
R1557 B.n459 B.n182 585
R1558 B.n461 B.n460 585
R1559 B.n462 B.n181 585
R1560 B.n464 B.n463 585
R1561 B.n465 B.n180 585
R1562 B.n467 B.n466 585
R1563 B.n468 B.n179 585
R1564 B.n470 B.n469 585
R1565 B.n471 B.n178 585
R1566 B.n473 B.n472 585
R1567 B.n474 B.n177 585
R1568 B.n476 B.n475 585
R1569 B.n477 B.n176 585
R1570 B.n479 B.n478 585
R1571 B.n480 B.n175 585
R1572 B.n482 B.n481 585
R1573 B.n483 B.n174 585
R1574 B.n485 B.n484 585
R1575 B.n486 B.n173 585
R1576 B.n488 B.n487 585
R1577 B.n489 B.n172 585
R1578 B.n491 B.n490 585
R1579 B.n492 B.n171 585
R1580 B.n494 B.n493 585
R1581 B.n495 B.n170 585
R1582 B.n497 B.n496 585
R1583 B.n498 B.n169 585
R1584 B.n500 B.n499 585
R1585 B.n501 B.n168 585
R1586 B.n503 B.n502 585
R1587 B.n504 B.n167 585
R1588 B.n506 B.n505 585
R1589 B.n507 B.n166 585
R1590 B.n509 B.n508 585
R1591 B.n510 B.n165 585
R1592 B.n512 B.n511 585
R1593 B.n513 B.n164 585
R1594 B.n515 B.n514 585
R1595 B.n353 B.n218 585
R1596 B.n352 B.n351 585
R1597 B.n350 B.n219 585
R1598 B.n349 B.n348 585
R1599 B.n347 B.n220 585
R1600 B.n346 B.n345 585
R1601 B.n344 B.n221 585
R1602 B.n343 B.n342 585
R1603 B.n341 B.n222 585
R1604 B.n340 B.n339 585
R1605 B.n338 B.n223 585
R1606 B.n337 B.n336 585
R1607 B.n335 B.n224 585
R1608 B.n334 B.n333 585
R1609 B.n332 B.n225 585
R1610 B.n331 B.n330 585
R1611 B.n329 B.n226 585
R1612 B.n328 B.n327 585
R1613 B.n326 B.n227 585
R1614 B.n325 B.n324 585
R1615 B.n323 B.n228 585
R1616 B.n322 B.n321 585
R1617 B.n320 B.n229 585
R1618 B.n319 B.n318 585
R1619 B.n317 B.n230 585
R1620 B.n316 B.n315 585
R1621 B.n314 B.n231 585
R1622 B.n313 B.n312 585
R1623 B.n311 B.n232 585
R1624 B.n310 B.n309 585
R1625 B.n308 B.n233 585
R1626 B.n307 B.n306 585
R1627 B.n305 B.n234 585
R1628 B.n304 B.n303 585
R1629 B.n302 B.n235 585
R1630 B.n301 B.n300 585
R1631 B.n299 B.n236 585
R1632 B.n298 B.n297 585
R1633 B.n296 B.n237 585
R1634 B.n295 B.n294 585
R1635 B.n293 B.n238 585
R1636 B.n292 B.n291 585
R1637 B.n290 B.n239 585
R1638 B.n289 B.n288 585
R1639 B.n287 B.n240 585
R1640 B.n286 B.n285 585
R1641 B.n284 B.n241 585
R1642 B.n283 B.n282 585
R1643 B.n281 B.n242 585
R1644 B.n280 B.n279 585
R1645 B.n278 B.n243 585
R1646 B.n277 B.n276 585
R1647 B.n275 B.n244 585
R1648 B.n274 B.n273 585
R1649 B.n272 B.n245 585
R1650 B.n271 B.n270 585
R1651 B.n269 B.n246 585
R1652 B.n268 B.n267 585
R1653 B.n266 B.n247 585
R1654 B.n265 B.n264 585
R1655 B.n263 B.n248 585
R1656 B.n262 B.n261 585
R1657 B.n260 B.n249 585
R1658 B.n259 B.n258 585
R1659 B.n257 B.n250 585
R1660 B.n256 B.n255 585
R1661 B.n254 B.n251 585
R1662 B.n253 B.n252 585
R1663 B.n2 B.n0 585
R1664 B.n985 B.n1 585
R1665 B.n984 B.n983 585
R1666 B.n982 B.n3 585
R1667 B.n981 B.n980 585
R1668 B.n979 B.n4 585
R1669 B.n978 B.n977 585
R1670 B.n976 B.n5 585
R1671 B.n975 B.n974 585
R1672 B.n973 B.n6 585
R1673 B.n972 B.n971 585
R1674 B.n970 B.n7 585
R1675 B.n969 B.n968 585
R1676 B.n967 B.n8 585
R1677 B.n966 B.n965 585
R1678 B.n964 B.n9 585
R1679 B.n963 B.n962 585
R1680 B.n961 B.n10 585
R1681 B.n960 B.n959 585
R1682 B.n958 B.n11 585
R1683 B.n957 B.n956 585
R1684 B.n955 B.n12 585
R1685 B.n954 B.n953 585
R1686 B.n952 B.n13 585
R1687 B.n951 B.n950 585
R1688 B.n949 B.n14 585
R1689 B.n948 B.n947 585
R1690 B.n946 B.n15 585
R1691 B.n945 B.n944 585
R1692 B.n943 B.n16 585
R1693 B.n942 B.n941 585
R1694 B.n940 B.n17 585
R1695 B.n939 B.n938 585
R1696 B.n937 B.n18 585
R1697 B.n936 B.n935 585
R1698 B.n934 B.n19 585
R1699 B.n933 B.n932 585
R1700 B.n931 B.n20 585
R1701 B.n930 B.n929 585
R1702 B.n928 B.n21 585
R1703 B.n927 B.n926 585
R1704 B.n925 B.n22 585
R1705 B.n924 B.n923 585
R1706 B.n922 B.n23 585
R1707 B.n921 B.n920 585
R1708 B.n919 B.n24 585
R1709 B.n918 B.n917 585
R1710 B.n916 B.n25 585
R1711 B.n915 B.n914 585
R1712 B.n913 B.n26 585
R1713 B.n912 B.n911 585
R1714 B.n910 B.n27 585
R1715 B.n909 B.n908 585
R1716 B.n907 B.n28 585
R1717 B.n906 B.n905 585
R1718 B.n904 B.n29 585
R1719 B.n903 B.n902 585
R1720 B.n901 B.n30 585
R1721 B.n900 B.n899 585
R1722 B.n898 B.n31 585
R1723 B.n897 B.n896 585
R1724 B.n895 B.n32 585
R1725 B.n894 B.n893 585
R1726 B.n892 B.n33 585
R1727 B.n891 B.n890 585
R1728 B.n889 B.n34 585
R1729 B.n888 B.n887 585
R1730 B.n886 B.n35 585
R1731 B.n885 B.n884 585
R1732 B.n883 B.n36 585
R1733 B.n987 B.n986 585
R1734 B.n355 B.n218 502.111
R1735 B.n883 B.n882 502.111
R1736 B.n516 B.n515 502.111
R1737 B.n725 B.n94 502.111
R1738 B.n439 B.t11 494.115
R1739 B.n69 B.t1 494.115
R1740 B.n193 B.t8 494.115
R1741 B.n62 B.t4 494.115
R1742 B.n440 B.t10 414.017
R1743 B.n70 B.t2 414.017
R1744 B.n194 B.t7 414.017
R1745 B.n63 B.t5 414.017
R1746 B.n439 B.t9 298.957
R1747 B.n193 B.t6 298.957
R1748 B.n62 B.t3 298.957
R1749 B.n69 B.t0 298.957
R1750 B.n351 B.n218 163.367
R1751 B.n351 B.n350 163.367
R1752 B.n350 B.n349 163.367
R1753 B.n349 B.n220 163.367
R1754 B.n345 B.n220 163.367
R1755 B.n345 B.n344 163.367
R1756 B.n344 B.n343 163.367
R1757 B.n343 B.n222 163.367
R1758 B.n339 B.n222 163.367
R1759 B.n339 B.n338 163.367
R1760 B.n338 B.n337 163.367
R1761 B.n337 B.n224 163.367
R1762 B.n333 B.n224 163.367
R1763 B.n333 B.n332 163.367
R1764 B.n332 B.n331 163.367
R1765 B.n331 B.n226 163.367
R1766 B.n327 B.n226 163.367
R1767 B.n327 B.n326 163.367
R1768 B.n326 B.n325 163.367
R1769 B.n325 B.n228 163.367
R1770 B.n321 B.n228 163.367
R1771 B.n321 B.n320 163.367
R1772 B.n320 B.n319 163.367
R1773 B.n319 B.n230 163.367
R1774 B.n315 B.n230 163.367
R1775 B.n315 B.n314 163.367
R1776 B.n314 B.n313 163.367
R1777 B.n313 B.n232 163.367
R1778 B.n309 B.n232 163.367
R1779 B.n309 B.n308 163.367
R1780 B.n308 B.n307 163.367
R1781 B.n307 B.n234 163.367
R1782 B.n303 B.n234 163.367
R1783 B.n303 B.n302 163.367
R1784 B.n302 B.n301 163.367
R1785 B.n301 B.n236 163.367
R1786 B.n297 B.n236 163.367
R1787 B.n297 B.n296 163.367
R1788 B.n296 B.n295 163.367
R1789 B.n295 B.n238 163.367
R1790 B.n291 B.n238 163.367
R1791 B.n291 B.n290 163.367
R1792 B.n290 B.n289 163.367
R1793 B.n289 B.n240 163.367
R1794 B.n285 B.n240 163.367
R1795 B.n285 B.n284 163.367
R1796 B.n284 B.n283 163.367
R1797 B.n283 B.n242 163.367
R1798 B.n279 B.n242 163.367
R1799 B.n279 B.n278 163.367
R1800 B.n278 B.n277 163.367
R1801 B.n277 B.n244 163.367
R1802 B.n273 B.n244 163.367
R1803 B.n273 B.n272 163.367
R1804 B.n272 B.n271 163.367
R1805 B.n271 B.n246 163.367
R1806 B.n267 B.n246 163.367
R1807 B.n267 B.n266 163.367
R1808 B.n266 B.n265 163.367
R1809 B.n265 B.n248 163.367
R1810 B.n261 B.n248 163.367
R1811 B.n261 B.n260 163.367
R1812 B.n260 B.n259 163.367
R1813 B.n259 B.n250 163.367
R1814 B.n255 B.n250 163.367
R1815 B.n255 B.n254 163.367
R1816 B.n254 B.n253 163.367
R1817 B.n253 B.n2 163.367
R1818 B.n986 B.n2 163.367
R1819 B.n986 B.n985 163.367
R1820 B.n985 B.n984 163.367
R1821 B.n984 B.n3 163.367
R1822 B.n980 B.n3 163.367
R1823 B.n980 B.n979 163.367
R1824 B.n979 B.n978 163.367
R1825 B.n978 B.n5 163.367
R1826 B.n974 B.n5 163.367
R1827 B.n974 B.n973 163.367
R1828 B.n973 B.n972 163.367
R1829 B.n972 B.n7 163.367
R1830 B.n968 B.n7 163.367
R1831 B.n968 B.n967 163.367
R1832 B.n967 B.n966 163.367
R1833 B.n966 B.n9 163.367
R1834 B.n962 B.n9 163.367
R1835 B.n962 B.n961 163.367
R1836 B.n961 B.n960 163.367
R1837 B.n960 B.n11 163.367
R1838 B.n956 B.n11 163.367
R1839 B.n956 B.n955 163.367
R1840 B.n955 B.n954 163.367
R1841 B.n954 B.n13 163.367
R1842 B.n950 B.n13 163.367
R1843 B.n950 B.n949 163.367
R1844 B.n949 B.n948 163.367
R1845 B.n948 B.n15 163.367
R1846 B.n944 B.n15 163.367
R1847 B.n944 B.n943 163.367
R1848 B.n943 B.n942 163.367
R1849 B.n942 B.n17 163.367
R1850 B.n938 B.n17 163.367
R1851 B.n938 B.n937 163.367
R1852 B.n937 B.n936 163.367
R1853 B.n936 B.n19 163.367
R1854 B.n932 B.n19 163.367
R1855 B.n932 B.n931 163.367
R1856 B.n931 B.n930 163.367
R1857 B.n930 B.n21 163.367
R1858 B.n926 B.n21 163.367
R1859 B.n926 B.n925 163.367
R1860 B.n925 B.n924 163.367
R1861 B.n924 B.n23 163.367
R1862 B.n920 B.n23 163.367
R1863 B.n920 B.n919 163.367
R1864 B.n919 B.n918 163.367
R1865 B.n918 B.n25 163.367
R1866 B.n914 B.n25 163.367
R1867 B.n914 B.n913 163.367
R1868 B.n913 B.n912 163.367
R1869 B.n912 B.n27 163.367
R1870 B.n908 B.n27 163.367
R1871 B.n908 B.n907 163.367
R1872 B.n907 B.n906 163.367
R1873 B.n906 B.n29 163.367
R1874 B.n902 B.n29 163.367
R1875 B.n902 B.n901 163.367
R1876 B.n901 B.n900 163.367
R1877 B.n900 B.n31 163.367
R1878 B.n896 B.n31 163.367
R1879 B.n896 B.n895 163.367
R1880 B.n895 B.n894 163.367
R1881 B.n894 B.n33 163.367
R1882 B.n890 B.n33 163.367
R1883 B.n890 B.n889 163.367
R1884 B.n889 B.n888 163.367
R1885 B.n888 B.n35 163.367
R1886 B.n884 B.n35 163.367
R1887 B.n884 B.n883 163.367
R1888 B.n356 B.n355 163.367
R1889 B.n357 B.n356 163.367
R1890 B.n357 B.n216 163.367
R1891 B.n361 B.n216 163.367
R1892 B.n362 B.n361 163.367
R1893 B.n363 B.n362 163.367
R1894 B.n363 B.n214 163.367
R1895 B.n367 B.n214 163.367
R1896 B.n368 B.n367 163.367
R1897 B.n369 B.n368 163.367
R1898 B.n369 B.n212 163.367
R1899 B.n373 B.n212 163.367
R1900 B.n374 B.n373 163.367
R1901 B.n375 B.n374 163.367
R1902 B.n375 B.n210 163.367
R1903 B.n379 B.n210 163.367
R1904 B.n380 B.n379 163.367
R1905 B.n381 B.n380 163.367
R1906 B.n381 B.n208 163.367
R1907 B.n385 B.n208 163.367
R1908 B.n386 B.n385 163.367
R1909 B.n387 B.n386 163.367
R1910 B.n387 B.n206 163.367
R1911 B.n391 B.n206 163.367
R1912 B.n392 B.n391 163.367
R1913 B.n393 B.n392 163.367
R1914 B.n393 B.n204 163.367
R1915 B.n397 B.n204 163.367
R1916 B.n398 B.n397 163.367
R1917 B.n399 B.n398 163.367
R1918 B.n399 B.n202 163.367
R1919 B.n403 B.n202 163.367
R1920 B.n404 B.n403 163.367
R1921 B.n405 B.n404 163.367
R1922 B.n405 B.n200 163.367
R1923 B.n409 B.n200 163.367
R1924 B.n410 B.n409 163.367
R1925 B.n411 B.n410 163.367
R1926 B.n411 B.n198 163.367
R1927 B.n415 B.n198 163.367
R1928 B.n416 B.n415 163.367
R1929 B.n417 B.n416 163.367
R1930 B.n417 B.n196 163.367
R1931 B.n421 B.n196 163.367
R1932 B.n422 B.n421 163.367
R1933 B.n423 B.n422 163.367
R1934 B.n423 B.n192 163.367
R1935 B.n428 B.n192 163.367
R1936 B.n429 B.n428 163.367
R1937 B.n430 B.n429 163.367
R1938 B.n430 B.n190 163.367
R1939 B.n434 B.n190 163.367
R1940 B.n435 B.n434 163.367
R1941 B.n436 B.n435 163.367
R1942 B.n436 B.n188 163.367
R1943 B.n443 B.n188 163.367
R1944 B.n444 B.n443 163.367
R1945 B.n445 B.n444 163.367
R1946 B.n445 B.n186 163.367
R1947 B.n449 B.n186 163.367
R1948 B.n450 B.n449 163.367
R1949 B.n451 B.n450 163.367
R1950 B.n451 B.n184 163.367
R1951 B.n455 B.n184 163.367
R1952 B.n456 B.n455 163.367
R1953 B.n457 B.n456 163.367
R1954 B.n457 B.n182 163.367
R1955 B.n461 B.n182 163.367
R1956 B.n462 B.n461 163.367
R1957 B.n463 B.n462 163.367
R1958 B.n463 B.n180 163.367
R1959 B.n467 B.n180 163.367
R1960 B.n468 B.n467 163.367
R1961 B.n469 B.n468 163.367
R1962 B.n469 B.n178 163.367
R1963 B.n473 B.n178 163.367
R1964 B.n474 B.n473 163.367
R1965 B.n475 B.n474 163.367
R1966 B.n475 B.n176 163.367
R1967 B.n479 B.n176 163.367
R1968 B.n480 B.n479 163.367
R1969 B.n481 B.n480 163.367
R1970 B.n481 B.n174 163.367
R1971 B.n485 B.n174 163.367
R1972 B.n486 B.n485 163.367
R1973 B.n487 B.n486 163.367
R1974 B.n487 B.n172 163.367
R1975 B.n491 B.n172 163.367
R1976 B.n492 B.n491 163.367
R1977 B.n493 B.n492 163.367
R1978 B.n493 B.n170 163.367
R1979 B.n497 B.n170 163.367
R1980 B.n498 B.n497 163.367
R1981 B.n499 B.n498 163.367
R1982 B.n499 B.n168 163.367
R1983 B.n503 B.n168 163.367
R1984 B.n504 B.n503 163.367
R1985 B.n505 B.n504 163.367
R1986 B.n505 B.n166 163.367
R1987 B.n509 B.n166 163.367
R1988 B.n510 B.n509 163.367
R1989 B.n511 B.n510 163.367
R1990 B.n511 B.n164 163.367
R1991 B.n515 B.n164 163.367
R1992 B.n517 B.n516 163.367
R1993 B.n517 B.n162 163.367
R1994 B.n521 B.n162 163.367
R1995 B.n522 B.n521 163.367
R1996 B.n523 B.n522 163.367
R1997 B.n523 B.n160 163.367
R1998 B.n527 B.n160 163.367
R1999 B.n528 B.n527 163.367
R2000 B.n529 B.n528 163.367
R2001 B.n529 B.n158 163.367
R2002 B.n533 B.n158 163.367
R2003 B.n534 B.n533 163.367
R2004 B.n535 B.n534 163.367
R2005 B.n535 B.n156 163.367
R2006 B.n539 B.n156 163.367
R2007 B.n540 B.n539 163.367
R2008 B.n541 B.n540 163.367
R2009 B.n541 B.n154 163.367
R2010 B.n545 B.n154 163.367
R2011 B.n546 B.n545 163.367
R2012 B.n547 B.n546 163.367
R2013 B.n547 B.n152 163.367
R2014 B.n551 B.n152 163.367
R2015 B.n552 B.n551 163.367
R2016 B.n553 B.n552 163.367
R2017 B.n553 B.n150 163.367
R2018 B.n557 B.n150 163.367
R2019 B.n558 B.n557 163.367
R2020 B.n559 B.n558 163.367
R2021 B.n559 B.n148 163.367
R2022 B.n563 B.n148 163.367
R2023 B.n564 B.n563 163.367
R2024 B.n565 B.n564 163.367
R2025 B.n565 B.n146 163.367
R2026 B.n569 B.n146 163.367
R2027 B.n570 B.n569 163.367
R2028 B.n571 B.n570 163.367
R2029 B.n571 B.n144 163.367
R2030 B.n575 B.n144 163.367
R2031 B.n576 B.n575 163.367
R2032 B.n577 B.n576 163.367
R2033 B.n577 B.n142 163.367
R2034 B.n581 B.n142 163.367
R2035 B.n582 B.n581 163.367
R2036 B.n583 B.n582 163.367
R2037 B.n583 B.n140 163.367
R2038 B.n587 B.n140 163.367
R2039 B.n588 B.n587 163.367
R2040 B.n589 B.n588 163.367
R2041 B.n589 B.n138 163.367
R2042 B.n593 B.n138 163.367
R2043 B.n594 B.n593 163.367
R2044 B.n595 B.n594 163.367
R2045 B.n595 B.n136 163.367
R2046 B.n599 B.n136 163.367
R2047 B.n600 B.n599 163.367
R2048 B.n601 B.n600 163.367
R2049 B.n601 B.n134 163.367
R2050 B.n605 B.n134 163.367
R2051 B.n606 B.n605 163.367
R2052 B.n607 B.n606 163.367
R2053 B.n607 B.n132 163.367
R2054 B.n611 B.n132 163.367
R2055 B.n612 B.n611 163.367
R2056 B.n613 B.n612 163.367
R2057 B.n613 B.n130 163.367
R2058 B.n617 B.n130 163.367
R2059 B.n618 B.n617 163.367
R2060 B.n619 B.n618 163.367
R2061 B.n619 B.n128 163.367
R2062 B.n623 B.n128 163.367
R2063 B.n624 B.n623 163.367
R2064 B.n625 B.n624 163.367
R2065 B.n625 B.n126 163.367
R2066 B.n629 B.n126 163.367
R2067 B.n630 B.n629 163.367
R2068 B.n631 B.n630 163.367
R2069 B.n631 B.n124 163.367
R2070 B.n635 B.n124 163.367
R2071 B.n636 B.n635 163.367
R2072 B.n637 B.n636 163.367
R2073 B.n637 B.n122 163.367
R2074 B.n641 B.n122 163.367
R2075 B.n642 B.n641 163.367
R2076 B.n643 B.n642 163.367
R2077 B.n643 B.n120 163.367
R2078 B.n647 B.n120 163.367
R2079 B.n648 B.n647 163.367
R2080 B.n649 B.n648 163.367
R2081 B.n649 B.n118 163.367
R2082 B.n653 B.n118 163.367
R2083 B.n654 B.n653 163.367
R2084 B.n655 B.n654 163.367
R2085 B.n655 B.n116 163.367
R2086 B.n659 B.n116 163.367
R2087 B.n660 B.n659 163.367
R2088 B.n661 B.n660 163.367
R2089 B.n661 B.n114 163.367
R2090 B.n665 B.n114 163.367
R2091 B.n666 B.n665 163.367
R2092 B.n667 B.n666 163.367
R2093 B.n667 B.n112 163.367
R2094 B.n671 B.n112 163.367
R2095 B.n672 B.n671 163.367
R2096 B.n673 B.n672 163.367
R2097 B.n673 B.n110 163.367
R2098 B.n677 B.n110 163.367
R2099 B.n678 B.n677 163.367
R2100 B.n679 B.n678 163.367
R2101 B.n679 B.n108 163.367
R2102 B.n683 B.n108 163.367
R2103 B.n684 B.n683 163.367
R2104 B.n685 B.n684 163.367
R2105 B.n685 B.n106 163.367
R2106 B.n689 B.n106 163.367
R2107 B.n690 B.n689 163.367
R2108 B.n691 B.n690 163.367
R2109 B.n691 B.n104 163.367
R2110 B.n695 B.n104 163.367
R2111 B.n696 B.n695 163.367
R2112 B.n697 B.n696 163.367
R2113 B.n697 B.n102 163.367
R2114 B.n701 B.n102 163.367
R2115 B.n702 B.n701 163.367
R2116 B.n703 B.n702 163.367
R2117 B.n703 B.n100 163.367
R2118 B.n707 B.n100 163.367
R2119 B.n708 B.n707 163.367
R2120 B.n709 B.n708 163.367
R2121 B.n709 B.n98 163.367
R2122 B.n713 B.n98 163.367
R2123 B.n714 B.n713 163.367
R2124 B.n715 B.n714 163.367
R2125 B.n715 B.n96 163.367
R2126 B.n719 B.n96 163.367
R2127 B.n720 B.n719 163.367
R2128 B.n721 B.n720 163.367
R2129 B.n721 B.n94 163.367
R2130 B.n882 B.n37 163.367
R2131 B.n878 B.n37 163.367
R2132 B.n878 B.n877 163.367
R2133 B.n877 B.n876 163.367
R2134 B.n876 B.n39 163.367
R2135 B.n872 B.n39 163.367
R2136 B.n872 B.n871 163.367
R2137 B.n871 B.n870 163.367
R2138 B.n870 B.n41 163.367
R2139 B.n866 B.n41 163.367
R2140 B.n866 B.n865 163.367
R2141 B.n865 B.n864 163.367
R2142 B.n864 B.n43 163.367
R2143 B.n860 B.n43 163.367
R2144 B.n860 B.n859 163.367
R2145 B.n859 B.n858 163.367
R2146 B.n858 B.n45 163.367
R2147 B.n854 B.n45 163.367
R2148 B.n854 B.n853 163.367
R2149 B.n853 B.n852 163.367
R2150 B.n852 B.n47 163.367
R2151 B.n848 B.n47 163.367
R2152 B.n848 B.n847 163.367
R2153 B.n847 B.n846 163.367
R2154 B.n846 B.n49 163.367
R2155 B.n842 B.n49 163.367
R2156 B.n842 B.n841 163.367
R2157 B.n841 B.n840 163.367
R2158 B.n840 B.n51 163.367
R2159 B.n836 B.n51 163.367
R2160 B.n836 B.n835 163.367
R2161 B.n835 B.n834 163.367
R2162 B.n834 B.n53 163.367
R2163 B.n830 B.n53 163.367
R2164 B.n830 B.n829 163.367
R2165 B.n829 B.n828 163.367
R2166 B.n828 B.n55 163.367
R2167 B.n824 B.n55 163.367
R2168 B.n824 B.n823 163.367
R2169 B.n823 B.n822 163.367
R2170 B.n822 B.n57 163.367
R2171 B.n818 B.n57 163.367
R2172 B.n818 B.n817 163.367
R2173 B.n817 B.n816 163.367
R2174 B.n816 B.n59 163.367
R2175 B.n812 B.n59 163.367
R2176 B.n812 B.n811 163.367
R2177 B.n811 B.n810 163.367
R2178 B.n810 B.n61 163.367
R2179 B.n806 B.n61 163.367
R2180 B.n806 B.n805 163.367
R2181 B.n805 B.n804 163.367
R2182 B.n804 B.n66 163.367
R2183 B.n800 B.n66 163.367
R2184 B.n800 B.n799 163.367
R2185 B.n799 B.n798 163.367
R2186 B.n798 B.n68 163.367
R2187 B.n793 B.n68 163.367
R2188 B.n793 B.n792 163.367
R2189 B.n792 B.n791 163.367
R2190 B.n791 B.n72 163.367
R2191 B.n787 B.n72 163.367
R2192 B.n787 B.n786 163.367
R2193 B.n786 B.n785 163.367
R2194 B.n785 B.n74 163.367
R2195 B.n781 B.n74 163.367
R2196 B.n781 B.n780 163.367
R2197 B.n780 B.n779 163.367
R2198 B.n779 B.n76 163.367
R2199 B.n775 B.n76 163.367
R2200 B.n775 B.n774 163.367
R2201 B.n774 B.n773 163.367
R2202 B.n773 B.n78 163.367
R2203 B.n769 B.n78 163.367
R2204 B.n769 B.n768 163.367
R2205 B.n768 B.n767 163.367
R2206 B.n767 B.n80 163.367
R2207 B.n763 B.n80 163.367
R2208 B.n763 B.n762 163.367
R2209 B.n762 B.n761 163.367
R2210 B.n761 B.n82 163.367
R2211 B.n757 B.n82 163.367
R2212 B.n757 B.n756 163.367
R2213 B.n756 B.n755 163.367
R2214 B.n755 B.n84 163.367
R2215 B.n751 B.n84 163.367
R2216 B.n751 B.n750 163.367
R2217 B.n750 B.n749 163.367
R2218 B.n749 B.n86 163.367
R2219 B.n745 B.n86 163.367
R2220 B.n745 B.n744 163.367
R2221 B.n744 B.n743 163.367
R2222 B.n743 B.n88 163.367
R2223 B.n739 B.n88 163.367
R2224 B.n739 B.n738 163.367
R2225 B.n738 B.n737 163.367
R2226 B.n737 B.n90 163.367
R2227 B.n733 B.n90 163.367
R2228 B.n733 B.n732 163.367
R2229 B.n732 B.n731 163.367
R2230 B.n731 B.n92 163.367
R2231 B.n727 B.n92 163.367
R2232 B.n727 B.n726 163.367
R2233 B.n726 B.n725 163.367
R2234 B.n440 B.n439 80.0975
R2235 B.n194 B.n193 80.0975
R2236 B.n63 B.n62 80.0975
R2237 B.n70 B.n69 80.0975
R2238 B.n441 B.n440 59.5399
R2239 B.n426 B.n194 59.5399
R2240 B.n64 B.n63 59.5399
R2241 B.n796 B.n70 59.5399
R2242 B.n881 B.n36 32.6249
R2243 B.n724 B.n723 32.6249
R2244 B.n514 B.n163 32.6249
R2245 B.n354 B.n353 32.6249
R2246 B B.n987 18.0485
R2247 B.n881 B.n880 10.6151
R2248 B.n880 B.n879 10.6151
R2249 B.n879 B.n38 10.6151
R2250 B.n875 B.n38 10.6151
R2251 B.n875 B.n874 10.6151
R2252 B.n874 B.n873 10.6151
R2253 B.n873 B.n40 10.6151
R2254 B.n869 B.n40 10.6151
R2255 B.n869 B.n868 10.6151
R2256 B.n868 B.n867 10.6151
R2257 B.n867 B.n42 10.6151
R2258 B.n863 B.n42 10.6151
R2259 B.n863 B.n862 10.6151
R2260 B.n862 B.n861 10.6151
R2261 B.n861 B.n44 10.6151
R2262 B.n857 B.n44 10.6151
R2263 B.n857 B.n856 10.6151
R2264 B.n856 B.n855 10.6151
R2265 B.n855 B.n46 10.6151
R2266 B.n851 B.n46 10.6151
R2267 B.n851 B.n850 10.6151
R2268 B.n850 B.n849 10.6151
R2269 B.n849 B.n48 10.6151
R2270 B.n845 B.n48 10.6151
R2271 B.n845 B.n844 10.6151
R2272 B.n844 B.n843 10.6151
R2273 B.n843 B.n50 10.6151
R2274 B.n839 B.n50 10.6151
R2275 B.n839 B.n838 10.6151
R2276 B.n838 B.n837 10.6151
R2277 B.n837 B.n52 10.6151
R2278 B.n833 B.n52 10.6151
R2279 B.n833 B.n832 10.6151
R2280 B.n832 B.n831 10.6151
R2281 B.n831 B.n54 10.6151
R2282 B.n827 B.n54 10.6151
R2283 B.n827 B.n826 10.6151
R2284 B.n826 B.n825 10.6151
R2285 B.n825 B.n56 10.6151
R2286 B.n821 B.n56 10.6151
R2287 B.n821 B.n820 10.6151
R2288 B.n820 B.n819 10.6151
R2289 B.n819 B.n58 10.6151
R2290 B.n815 B.n58 10.6151
R2291 B.n815 B.n814 10.6151
R2292 B.n814 B.n813 10.6151
R2293 B.n813 B.n60 10.6151
R2294 B.n809 B.n808 10.6151
R2295 B.n808 B.n807 10.6151
R2296 B.n807 B.n65 10.6151
R2297 B.n803 B.n65 10.6151
R2298 B.n803 B.n802 10.6151
R2299 B.n802 B.n801 10.6151
R2300 B.n801 B.n67 10.6151
R2301 B.n797 B.n67 10.6151
R2302 B.n795 B.n794 10.6151
R2303 B.n794 B.n71 10.6151
R2304 B.n790 B.n71 10.6151
R2305 B.n790 B.n789 10.6151
R2306 B.n789 B.n788 10.6151
R2307 B.n788 B.n73 10.6151
R2308 B.n784 B.n73 10.6151
R2309 B.n784 B.n783 10.6151
R2310 B.n783 B.n782 10.6151
R2311 B.n782 B.n75 10.6151
R2312 B.n778 B.n75 10.6151
R2313 B.n778 B.n777 10.6151
R2314 B.n777 B.n776 10.6151
R2315 B.n776 B.n77 10.6151
R2316 B.n772 B.n77 10.6151
R2317 B.n772 B.n771 10.6151
R2318 B.n771 B.n770 10.6151
R2319 B.n770 B.n79 10.6151
R2320 B.n766 B.n79 10.6151
R2321 B.n766 B.n765 10.6151
R2322 B.n765 B.n764 10.6151
R2323 B.n764 B.n81 10.6151
R2324 B.n760 B.n81 10.6151
R2325 B.n760 B.n759 10.6151
R2326 B.n759 B.n758 10.6151
R2327 B.n758 B.n83 10.6151
R2328 B.n754 B.n83 10.6151
R2329 B.n754 B.n753 10.6151
R2330 B.n753 B.n752 10.6151
R2331 B.n752 B.n85 10.6151
R2332 B.n748 B.n85 10.6151
R2333 B.n748 B.n747 10.6151
R2334 B.n747 B.n746 10.6151
R2335 B.n746 B.n87 10.6151
R2336 B.n742 B.n87 10.6151
R2337 B.n742 B.n741 10.6151
R2338 B.n741 B.n740 10.6151
R2339 B.n740 B.n89 10.6151
R2340 B.n736 B.n89 10.6151
R2341 B.n736 B.n735 10.6151
R2342 B.n735 B.n734 10.6151
R2343 B.n734 B.n91 10.6151
R2344 B.n730 B.n91 10.6151
R2345 B.n730 B.n729 10.6151
R2346 B.n729 B.n728 10.6151
R2347 B.n728 B.n93 10.6151
R2348 B.n724 B.n93 10.6151
R2349 B.n518 B.n163 10.6151
R2350 B.n519 B.n518 10.6151
R2351 B.n520 B.n519 10.6151
R2352 B.n520 B.n161 10.6151
R2353 B.n524 B.n161 10.6151
R2354 B.n525 B.n524 10.6151
R2355 B.n526 B.n525 10.6151
R2356 B.n526 B.n159 10.6151
R2357 B.n530 B.n159 10.6151
R2358 B.n531 B.n530 10.6151
R2359 B.n532 B.n531 10.6151
R2360 B.n532 B.n157 10.6151
R2361 B.n536 B.n157 10.6151
R2362 B.n537 B.n536 10.6151
R2363 B.n538 B.n537 10.6151
R2364 B.n538 B.n155 10.6151
R2365 B.n542 B.n155 10.6151
R2366 B.n543 B.n542 10.6151
R2367 B.n544 B.n543 10.6151
R2368 B.n544 B.n153 10.6151
R2369 B.n548 B.n153 10.6151
R2370 B.n549 B.n548 10.6151
R2371 B.n550 B.n549 10.6151
R2372 B.n550 B.n151 10.6151
R2373 B.n554 B.n151 10.6151
R2374 B.n555 B.n554 10.6151
R2375 B.n556 B.n555 10.6151
R2376 B.n556 B.n149 10.6151
R2377 B.n560 B.n149 10.6151
R2378 B.n561 B.n560 10.6151
R2379 B.n562 B.n561 10.6151
R2380 B.n562 B.n147 10.6151
R2381 B.n566 B.n147 10.6151
R2382 B.n567 B.n566 10.6151
R2383 B.n568 B.n567 10.6151
R2384 B.n568 B.n145 10.6151
R2385 B.n572 B.n145 10.6151
R2386 B.n573 B.n572 10.6151
R2387 B.n574 B.n573 10.6151
R2388 B.n574 B.n143 10.6151
R2389 B.n578 B.n143 10.6151
R2390 B.n579 B.n578 10.6151
R2391 B.n580 B.n579 10.6151
R2392 B.n580 B.n141 10.6151
R2393 B.n584 B.n141 10.6151
R2394 B.n585 B.n584 10.6151
R2395 B.n586 B.n585 10.6151
R2396 B.n586 B.n139 10.6151
R2397 B.n590 B.n139 10.6151
R2398 B.n591 B.n590 10.6151
R2399 B.n592 B.n591 10.6151
R2400 B.n592 B.n137 10.6151
R2401 B.n596 B.n137 10.6151
R2402 B.n597 B.n596 10.6151
R2403 B.n598 B.n597 10.6151
R2404 B.n598 B.n135 10.6151
R2405 B.n602 B.n135 10.6151
R2406 B.n603 B.n602 10.6151
R2407 B.n604 B.n603 10.6151
R2408 B.n604 B.n133 10.6151
R2409 B.n608 B.n133 10.6151
R2410 B.n609 B.n608 10.6151
R2411 B.n610 B.n609 10.6151
R2412 B.n610 B.n131 10.6151
R2413 B.n614 B.n131 10.6151
R2414 B.n615 B.n614 10.6151
R2415 B.n616 B.n615 10.6151
R2416 B.n616 B.n129 10.6151
R2417 B.n620 B.n129 10.6151
R2418 B.n621 B.n620 10.6151
R2419 B.n622 B.n621 10.6151
R2420 B.n622 B.n127 10.6151
R2421 B.n626 B.n127 10.6151
R2422 B.n627 B.n626 10.6151
R2423 B.n628 B.n627 10.6151
R2424 B.n628 B.n125 10.6151
R2425 B.n632 B.n125 10.6151
R2426 B.n633 B.n632 10.6151
R2427 B.n634 B.n633 10.6151
R2428 B.n634 B.n123 10.6151
R2429 B.n638 B.n123 10.6151
R2430 B.n639 B.n638 10.6151
R2431 B.n640 B.n639 10.6151
R2432 B.n640 B.n121 10.6151
R2433 B.n644 B.n121 10.6151
R2434 B.n645 B.n644 10.6151
R2435 B.n646 B.n645 10.6151
R2436 B.n646 B.n119 10.6151
R2437 B.n650 B.n119 10.6151
R2438 B.n651 B.n650 10.6151
R2439 B.n652 B.n651 10.6151
R2440 B.n652 B.n117 10.6151
R2441 B.n656 B.n117 10.6151
R2442 B.n657 B.n656 10.6151
R2443 B.n658 B.n657 10.6151
R2444 B.n658 B.n115 10.6151
R2445 B.n662 B.n115 10.6151
R2446 B.n663 B.n662 10.6151
R2447 B.n664 B.n663 10.6151
R2448 B.n664 B.n113 10.6151
R2449 B.n668 B.n113 10.6151
R2450 B.n669 B.n668 10.6151
R2451 B.n670 B.n669 10.6151
R2452 B.n670 B.n111 10.6151
R2453 B.n674 B.n111 10.6151
R2454 B.n675 B.n674 10.6151
R2455 B.n676 B.n675 10.6151
R2456 B.n676 B.n109 10.6151
R2457 B.n680 B.n109 10.6151
R2458 B.n681 B.n680 10.6151
R2459 B.n682 B.n681 10.6151
R2460 B.n682 B.n107 10.6151
R2461 B.n686 B.n107 10.6151
R2462 B.n687 B.n686 10.6151
R2463 B.n688 B.n687 10.6151
R2464 B.n688 B.n105 10.6151
R2465 B.n692 B.n105 10.6151
R2466 B.n693 B.n692 10.6151
R2467 B.n694 B.n693 10.6151
R2468 B.n694 B.n103 10.6151
R2469 B.n698 B.n103 10.6151
R2470 B.n699 B.n698 10.6151
R2471 B.n700 B.n699 10.6151
R2472 B.n700 B.n101 10.6151
R2473 B.n704 B.n101 10.6151
R2474 B.n705 B.n704 10.6151
R2475 B.n706 B.n705 10.6151
R2476 B.n706 B.n99 10.6151
R2477 B.n710 B.n99 10.6151
R2478 B.n711 B.n710 10.6151
R2479 B.n712 B.n711 10.6151
R2480 B.n712 B.n97 10.6151
R2481 B.n716 B.n97 10.6151
R2482 B.n717 B.n716 10.6151
R2483 B.n718 B.n717 10.6151
R2484 B.n718 B.n95 10.6151
R2485 B.n722 B.n95 10.6151
R2486 B.n723 B.n722 10.6151
R2487 B.n354 B.n217 10.6151
R2488 B.n358 B.n217 10.6151
R2489 B.n359 B.n358 10.6151
R2490 B.n360 B.n359 10.6151
R2491 B.n360 B.n215 10.6151
R2492 B.n364 B.n215 10.6151
R2493 B.n365 B.n364 10.6151
R2494 B.n366 B.n365 10.6151
R2495 B.n366 B.n213 10.6151
R2496 B.n370 B.n213 10.6151
R2497 B.n371 B.n370 10.6151
R2498 B.n372 B.n371 10.6151
R2499 B.n372 B.n211 10.6151
R2500 B.n376 B.n211 10.6151
R2501 B.n377 B.n376 10.6151
R2502 B.n378 B.n377 10.6151
R2503 B.n378 B.n209 10.6151
R2504 B.n382 B.n209 10.6151
R2505 B.n383 B.n382 10.6151
R2506 B.n384 B.n383 10.6151
R2507 B.n384 B.n207 10.6151
R2508 B.n388 B.n207 10.6151
R2509 B.n389 B.n388 10.6151
R2510 B.n390 B.n389 10.6151
R2511 B.n390 B.n205 10.6151
R2512 B.n394 B.n205 10.6151
R2513 B.n395 B.n394 10.6151
R2514 B.n396 B.n395 10.6151
R2515 B.n396 B.n203 10.6151
R2516 B.n400 B.n203 10.6151
R2517 B.n401 B.n400 10.6151
R2518 B.n402 B.n401 10.6151
R2519 B.n402 B.n201 10.6151
R2520 B.n406 B.n201 10.6151
R2521 B.n407 B.n406 10.6151
R2522 B.n408 B.n407 10.6151
R2523 B.n408 B.n199 10.6151
R2524 B.n412 B.n199 10.6151
R2525 B.n413 B.n412 10.6151
R2526 B.n414 B.n413 10.6151
R2527 B.n414 B.n197 10.6151
R2528 B.n418 B.n197 10.6151
R2529 B.n419 B.n418 10.6151
R2530 B.n420 B.n419 10.6151
R2531 B.n420 B.n195 10.6151
R2532 B.n424 B.n195 10.6151
R2533 B.n425 B.n424 10.6151
R2534 B.n427 B.n191 10.6151
R2535 B.n431 B.n191 10.6151
R2536 B.n432 B.n431 10.6151
R2537 B.n433 B.n432 10.6151
R2538 B.n433 B.n189 10.6151
R2539 B.n437 B.n189 10.6151
R2540 B.n438 B.n437 10.6151
R2541 B.n442 B.n438 10.6151
R2542 B.n446 B.n187 10.6151
R2543 B.n447 B.n446 10.6151
R2544 B.n448 B.n447 10.6151
R2545 B.n448 B.n185 10.6151
R2546 B.n452 B.n185 10.6151
R2547 B.n453 B.n452 10.6151
R2548 B.n454 B.n453 10.6151
R2549 B.n454 B.n183 10.6151
R2550 B.n458 B.n183 10.6151
R2551 B.n459 B.n458 10.6151
R2552 B.n460 B.n459 10.6151
R2553 B.n460 B.n181 10.6151
R2554 B.n464 B.n181 10.6151
R2555 B.n465 B.n464 10.6151
R2556 B.n466 B.n465 10.6151
R2557 B.n466 B.n179 10.6151
R2558 B.n470 B.n179 10.6151
R2559 B.n471 B.n470 10.6151
R2560 B.n472 B.n471 10.6151
R2561 B.n472 B.n177 10.6151
R2562 B.n476 B.n177 10.6151
R2563 B.n477 B.n476 10.6151
R2564 B.n478 B.n477 10.6151
R2565 B.n478 B.n175 10.6151
R2566 B.n482 B.n175 10.6151
R2567 B.n483 B.n482 10.6151
R2568 B.n484 B.n483 10.6151
R2569 B.n484 B.n173 10.6151
R2570 B.n488 B.n173 10.6151
R2571 B.n489 B.n488 10.6151
R2572 B.n490 B.n489 10.6151
R2573 B.n490 B.n171 10.6151
R2574 B.n494 B.n171 10.6151
R2575 B.n495 B.n494 10.6151
R2576 B.n496 B.n495 10.6151
R2577 B.n496 B.n169 10.6151
R2578 B.n500 B.n169 10.6151
R2579 B.n501 B.n500 10.6151
R2580 B.n502 B.n501 10.6151
R2581 B.n502 B.n167 10.6151
R2582 B.n506 B.n167 10.6151
R2583 B.n507 B.n506 10.6151
R2584 B.n508 B.n507 10.6151
R2585 B.n508 B.n165 10.6151
R2586 B.n512 B.n165 10.6151
R2587 B.n513 B.n512 10.6151
R2588 B.n514 B.n513 10.6151
R2589 B.n353 B.n352 10.6151
R2590 B.n352 B.n219 10.6151
R2591 B.n348 B.n219 10.6151
R2592 B.n348 B.n347 10.6151
R2593 B.n347 B.n346 10.6151
R2594 B.n346 B.n221 10.6151
R2595 B.n342 B.n221 10.6151
R2596 B.n342 B.n341 10.6151
R2597 B.n341 B.n340 10.6151
R2598 B.n340 B.n223 10.6151
R2599 B.n336 B.n223 10.6151
R2600 B.n336 B.n335 10.6151
R2601 B.n335 B.n334 10.6151
R2602 B.n334 B.n225 10.6151
R2603 B.n330 B.n225 10.6151
R2604 B.n330 B.n329 10.6151
R2605 B.n329 B.n328 10.6151
R2606 B.n328 B.n227 10.6151
R2607 B.n324 B.n227 10.6151
R2608 B.n324 B.n323 10.6151
R2609 B.n323 B.n322 10.6151
R2610 B.n322 B.n229 10.6151
R2611 B.n318 B.n229 10.6151
R2612 B.n318 B.n317 10.6151
R2613 B.n317 B.n316 10.6151
R2614 B.n316 B.n231 10.6151
R2615 B.n312 B.n231 10.6151
R2616 B.n312 B.n311 10.6151
R2617 B.n311 B.n310 10.6151
R2618 B.n310 B.n233 10.6151
R2619 B.n306 B.n233 10.6151
R2620 B.n306 B.n305 10.6151
R2621 B.n305 B.n304 10.6151
R2622 B.n304 B.n235 10.6151
R2623 B.n300 B.n235 10.6151
R2624 B.n300 B.n299 10.6151
R2625 B.n299 B.n298 10.6151
R2626 B.n298 B.n237 10.6151
R2627 B.n294 B.n237 10.6151
R2628 B.n294 B.n293 10.6151
R2629 B.n293 B.n292 10.6151
R2630 B.n292 B.n239 10.6151
R2631 B.n288 B.n239 10.6151
R2632 B.n288 B.n287 10.6151
R2633 B.n287 B.n286 10.6151
R2634 B.n286 B.n241 10.6151
R2635 B.n282 B.n241 10.6151
R2636 B.n282 B.n281 10.6151
R2637 B.n281 B.n280 10.6151
R2638 B.n280 B.n243 10.6151
R2639 B.n276 B.n243 10.6151
R2640 B.n276 B.n275 10.6151
R2641 B.n275 B.n274 10.6151
R2642 B.n274 B.n245 10.6151
R2643 B.n270 B.n245 10.6151
R2644 B.n270 B.n269 10.6151
R2645 B.n269 B.n268 10.6151
R2646 B.n268 B.n247 10.6151
R2647 B.n264 B.n247 10.6151
R2648 B.n264 B.n263 10.6151
R2649 B.n263 B.n262 10.6151
R2650 B.n262 B.n249 10.6151
R2651 B.n258 B.n249 10.6151
R2652 B.n258 B.n257 10.6151
R2653 B.n257 B.n256 10.6151
R2654 B.n256 B.n251 10.6151
R2655 B.n252 B.n251 10.6151
R2656 B.n252 B.n0 10.6151
R2657 B.n983 B.n1 10.6151
R2658 B.n983 B.n982 10.6151
R2659 B.n982 B.n981 10.6151
R2660 B.n981 B.n4 10.6151
R2661 B.n977 B.n4 10.6151
R2662 B.n977 B.n976 10.6151
R2663 B.n976 B.n975 10.6151
R2664 B.n975 B.n6 10.6151
R2665 B.n971 B.n6 10.6151
R2666 B.n971 B.n970 10.6151
R2667 B.n970 B.n969 10.6151
R2668 B.n969 B.n8 10.6151
R2669 B.n965 B.n8 10.6151
R2670 B.n965 B.n964 10.6151
R2671 B.n964 B.n963 10.6151
R2672 B.n963 B.n10 10.6151
R2673 B.n959 B.n10 10.6151
R2674 B.n959 B.n958 10.6151
R2675 B.n958 B.n957 10.6151
R2676 B.n957 B.n12 10.6151
R2677 B.n953 B.n12 10.6151
R2678 B.n953 B.n952 10.6151
R2679 B.n952 B.n951 10.6151
R2680 B.n951 B.n14 10.6151
R2681 B.n947 B.n14 10.6151
R2682 B.n947 B.n946 10.6151
R2683 B.n946 B.n945 10.6151
R2684 B.n945 B.n16 10.6151
R2685 B.n941 B.n16 10.6151
R2686 B.n941 B.n940 10.6151
R2687 B.n940 B.n939 10.6151
R2688 B.n939 B.n18 10.6151
R2689 B.n935 B.n18 10.6151
R2690 B.n935 B.n934 10.6151
R2691 B.n934 B.n933 10.6151
R2692 B.n933 B.n20 10.6151
R2693 B.n929 B.n20 10.6151
R2694 B.n929 B.n928 10.6151
R2695 B.n928 B.n927 10.6151
R2696 B.n927 B.n22 10.6151
R2697 B.n923 B.n22 10.6151
R2698 B.n923 B.n922 10.6151
R2699 B.n922 B.n921 10.6151
R2700 B.n921 B.n24 10.6151
R2701 B.n917 B.n24 10.6151
R2702 B.n917 B.n916 10.6151
R2703 B.n916 B.n915 10.6151
R2704 B.n915 B.n26 10.6151
R2705 B.n911 B.n26 10.6151
R2706 B.n911 B.n910 10.6151
R2707 B.n910 B.n909 10.6151
R2708 B.n909 B.n28 10.6151
R2709 B.n905 B.n28 10.6151
R2710 B.n905 B.n904 10.6151
R2711 B.n904 B.n903 10.6151
R2712 B.n903 B.n30 10.6151
R2713 B.n899 B.n30 10.6151
R2714 B.n899 B.n898 10.6151
R2715 B.n898 B.n897 10.6151
R2716 B.n897 B.n32 10.6151
R2717 B.n893 B.n32 10.6151
R2718 B.n893 B.n892 10.6151
R2719 B.n892 B.n891 10.6151
R2720 B.n891 B.n34 10.6151
R2721 B.n887 B.n34 10.6151
R2722 B.n887 B.n886 10.6151
R2723 B.n886 B.n885 10.6151
R2724 B.n885 B.n36 10.6151
R2725 B.n809 B.n64 6.5566
R2726 B.n797 B.n796 6.5566
R2727 B.n427 B.n426 6.5566
R2728 B.n442 B.n441 6.5566
R2729 B.n64 B.n60 4.05904
R2730 B.n796 B.n795 4.05904
R2731 B.n426 B.n425 4.05904
R2732 B.n441 B.n187 4.05904
R2733 B.n987 B.n0 2.81026
R2734 B.n987 B.n1 2.81026
C0 VDD2 VTAIL 9.257719f
C1 B VN 1.52952f
C2 VDD1 VN 0.153868f
C3 VP VN 9.52946f
C4 VDD2 VN 10.8166f
C5 VN VTAIL 11.51f
C6 B w_n5100_n3794# 12.549299f
C7 w_n5100_n3794# VDD1 2.39667f
C8 VP w_n5100_n3794# 11.4277f
C9 w_n5100_n3794# VDD2 2.56172f
C10 w_n5100_n3794# VTAIL 4.78014f
C11 w_n5100_n3794# VN 10.7621f
C12 B VDD1 2.07339f
C13 B VP 2.65174f
C14 B VDD2 2.20717f
C15 VP VDD1 11.308f
C16 VDD1 VDD2 2.40007f
C17 VP VDD2 0.647335f
C18 B VTAIL 6.21081f
C19 VDD1 VTAIL 9.19526f
C20 VP VTAIL 11.524099f
C21 VDD2 VSUBS 2.5266f
C22 VDD1 VSUBS 3.37827f
C23 VTAIL VSUBS 1.653659f
C24 VN VSUBS 8.43016f
C25 VP VSUBS 4.910807f
C26 B VSUBS 6.521326f
C27 w_n5100_n3794# VSUBS 0.237517p
C28 B.n0 VSUBS 0.0051f
C29 B.n1 VSUBS 0.0051f
C30 B.n2 VSUBS 0.008064f
C31 B.n3 VSUBS 0.008064f
C32 B.n4 VSUBS 0.008064f
C33 B.n5 VSUBS 0.008064f
C34 B.n6 VSUBS 0.008064f
C35 B.n7 VSUBS 0.008064f
C36 B.n8 VSUBS 0.008064f
C37 B.n9 VSUBS 0.008064f
C38 B.n10 VSUBS 0.008064f
C39 B.n11 VSUBS 0.008064f
C40 B.n12 VSUBS 0.008064f
C41 B.n13 VSUBS 0.008064f
C42 B.n14 VSUBS 0.008064f
C43 B.n15 VSUBS 0.008064f
C44 B.n16 VSUBS 0.008064f
C45 B.n17 VSUBS 0.008064f
C46 B.n18 VSUBS 0.008064f
C47 B.n19 VSUBS 0.008064f
C48 B.n20 VSUBS 0.008064f
C49 B.n21 VSUBS 0.008064f
C50 B.n22 VSUBS 0.008064f
C51 B.n23 VSUBS 0.008064f
C52 B.n24 VSUBS 0.008064f
C53 B.n25 VSUBS 0.008064f
C54 B.n26 VSUBS 0.008064f
C55 B.n27 VSUBS 0.008064f
C56 B.n28 VSUBS 0.008064f
C57 B.n29 VSUBS 0.008064f
C58 B.n30 VSUBS 0.008064f
C59 B.n31 VSUBS 0.008064f
C60 B.n32 VSUBS 0.008064f
C61 B.n33 VSUBS 0.008064f
C62 B.n34 VSUBS 0.008064f
C63 B.n35 VSUBS 0.008064f
C64 B.n36 VSUBS 0.018659f
C65 B.n37 VSUBS 0.008064f
C66 B.n38 VSUBS 0.008064f
C67 B.n39 VSUBS 0.008064f
C68 B.n40 VSUBS 0.008064f
C69 B.n41 VSUBS 0.008064f
C70 B.n42 VSUBS 0.008064f
C71 B.n43 VSUBS 0.008064f
C72 B.n44 VSUBS 0.008064f
C73 B.n45 VSUBS 0.008064f
C74 B.n46 VSUBS 0.008064f
C75 B.n47 VSUBS 0.008064f
C76 B.n48 VSUBS 0.008064f
C77 B.n49 VSUBS 0.008064f
C78 B.n50 VSUBS 0.008064f
C79 B.n51 VSUBS 0.008064f
C80 B.n52 VSUBS 0.008064f
C81 B.n53 VSUBS 0.008064f
C82 B.n54 VSUBS 0.008064f
C83 B.n55 VSUBS 0.008064f
C84 B.n56 VSUBS 0.008064f
C85 B.n57 VSUBS 0.008064f
C86 B.n58 VSUBS 0.008064f
C87 B.n59 VSUBS 0.008064f
C88 B.n60 VSUBS 0.005574f
C89 B.n61 VSUBS 0.008064f
C90 B.t5 VSUBS 0.298858f
C91 B.t4 VSUBS 0.350298f
C92 B.t3 VSUBS 2.85944f
C93 B.n62 VSUBS 0.558414f
C94 B.n63 VSUBS 0.32883f
C95 B.n64 VSUBS 0.018684f
C96 B.n65 VSUBS 0.008064f
C97 B.n66 VSUBS 0.008064f
C98 B.n67 VSUBS 0.008064f
C99 B.n68 VSUBS 0.008064f
C100 B.t2 VSUBS 0.298862f
C101 B.t1 VSUBS 0.350301f
C102 B.t0 VSUBS 2.85944f
C103 B.n69 VSUBS 0.558411f
C104 B.n70 VSUBS 0.328826f
C105 B.n71 VSUBS 0.008064f
C106 B.n72 VSUBS 0.008064f
C107 B.n73 VSUBS 0.008064f
C108 B.n74 VSUBS 0.008064f
C109 B.n75 VSUBS 0.008064f
C110 B.n76 VSUBS 0.008064f
C111 B.n77 VSUBS 0.008064f
C112 B.n78 VSUBS 0.008064f
C113 B.n79 VSUBS 0.008064f
C114 B.n80 VSUBS 0.008064f
C115 B.n81 VSUBS 0.008064f
C116 B.n82 VSUBS 0.008064f
C117 B.n83 VSUBS 0.008064f
C118 B.n84 VSUBS 0.008064f
C119 B.n85 VSUBS 0.008064f
C120 B.n86 VSUBS 0.008064f
C121 B.n87 VSUBS 0.008064f
C122 B.n88 VSUBS 0.008064f
C123 B.n89 VSUBS 0.008064f
C124 B.n90 VSUBS 0.008064f
C125 B.n91 VSUBS 0.008064f
C126 B.n92 VSUBS 0.008064f
C127 B.n93 VSUBS 0.008064f
C128 B.n94 VSUBS 0.018659f
C129 B.n95 VSUBS 0.008064f
C130 B.n96 VSUBS 0.008064f
C131 B.n97 VSUBS 0.008064f
C132 B.n98 VSUBS 0.008064f
C133 B.n99 VSUBS 0.008064f
C134 B.n100 VSUBS 0.008064f
C135 B.n101 VSUBS 0.008064f
C136 B.n102 VSUBS 0.008064f
C137 B.n103 VSUBS 0.008064f
C138 B.n104 VSUBS 0.008064f
C139 B.n105 VSUBS 0.008064f
C140 B.n106 VSUBS 0.008064f
C141 B.n107 VSUBS 0.008064f
C142 B.n108 VSUBS 0.008064f
C143 B.n109 VSUBS 0.008064f
C144 B.n110 VSUBS 0.008064f
C145 B.n111 VSUBS 0.008064f
C146 B.n112 VSUBS 0.008064f
C147 B.n113 VSUBS 0.008064f
C148 B.n114 VSUBS 0.008064f
C149 B.n115 VSUBS 0.008064f
C150 B.n116 VSUBS 0.008064f
C151 B.n117 VSUBS 0.008064f
C152 B.n118 VSUBS 0.008064f
C153 B.n119 VSUBS 0.008064f
C154 B.n120 VSUBS 0.008064f
C155 B.n121 VSUBS 0.008064f
C156 B.n122 VSUBS 0.008064f
C157 B.n123 VSUBS 0.008064f
C158 B.n124 VSUBS 0.008064f
C159 B.n125 VSUBS 0.008064f
C160 B.n126 VSUBS 0.008064f
C161 B.n127 VSUBS 0.008064f
C162 B.n128 VSUBS 0.008064f
C163 B.n129 VSUBS 0.008064f
C164 B.n130 VSUBS 0.008064f
C165 B.n131 VSUBS 0.008064f
C166 B.n132 VSUBS 0.008064f
C167 B.n133 VSUBS 0.008064f
C168 B.n134 VSUBS 0.008064f
C169 B.n135 VSUBS 0.008064f
C170 B.n136 VSUBS 0.008064f
C171 B.n137 VSUBS 0.008064f
C172 B.n138 VSUBS 0.008064f
C173 B.n139 VSUBS 0.008064f
C174 B.n140 VSUBS 0.008064f
C175 B.n141 VSUBS 0.008064f
C176 B.n142 VSUBS 0.008064f
C177 B.n143 VSUBS 0.008064f
C178 B.n144 VSUBS 0.008064f
C179 B.n145 VSUBS 0.008064f
C180 B.n146 VSUBS 0.008064f
C181 B.n147 VSUBS 0.008064f
C182 B.n148 VSUBS 0.008064f
C183 B.n149 VSUBS 0.008064f
C184 B.n150 VSUBS 0.008064f
C185 B.n151 VSUBS 0.008064f
C186 B.n152 VSUBS 0.008064f
C187 B.n153 VSUBS 0.008064f
C188 B.n154 VSUBS 0.008064f
C189 B.n155 VSUBS 0.008064f
C190 B.n156 VSUBS 0.008064f
C191 B.n157 VSUBS 0.008064f
C192 B.n158 VSUBS 0.008064f
C193 B.n159 VSUBS 0.008064f
C194 B.n160 VSUBS 0.008064f
C195 B.n161 VSUBS 0.008064f
C196 B.n162 VSUBS 0.008064f
C197 B.n163 VSUBS 0.018659f
C198 B.n164 VSUBS 0.008064f
C199 B.n165 VSUBS 0.008064f
C200 B.n166 VSUBS 0.008064f
C201 B.n167 VSUBS 0.008064f
C202 B.n168 VSUBS 0.008064f
C203 B.n169 VSUBS 0.008064f
C204 B.n170 VSUBS 0.008064f
C205 B.n171 VSUBS 0.008064f
C206 B.n172 VSUBS 0.008064f
C207 B.n173 VSUBS 0.008064f
C208 B.n174 VSUBS 0.008064f
C209 B.n175 VSUBS 0.008064f
C210 B.n176 VSUBS 0.008064f
C211 B.n177 VSUBS 0.008064f
C212 B.n178 VSUBS 0.008064f
C213 B.n179 VSUBS 0.008064f
C214 B.n180 VSUBS 0.008064f
C215 B.n181 VSUBS 0.008064f
C216 B.n182 VSUBS 0.008064f
C217 B.n183 VSUBS 0.008064f
C218 B.n184 VSUBS 0.008064f
C219 B.n185 VSUBS 0.008064f
C220 B.n186 VSUBS 0.008064f
C221 B.n187 VSUBS 0.005574f
C222 B.n188 VSUBS 0.008064f
C223 B.n189 VSUBS 0.008064f
C224 B.n190 VSUBS 0.008064f
C225 B.n191 VSUBS 0.008064f
C226 B.n192 VSUBS 0.008064f
C227 B.t7 VSUBS 0.298858f
C228 B.t8 VSUBS 0.350298f
C229 B.t6 VSUBS 2.85944f
C230 B.n193 VSUBS 0.558414f
C231 B.n194 VSUBS 0.32883f
C232 B.n195 VSUBS 0.008064f
C233 B.n196 VSUBS 0.008064f
C234 B.n197 VSUBS 0.008064f
C235 B.n198 VSUBS 0.008064f
C236 B.n199 VSUBS 0.008064f
C237 B.n200 VSUBS 0.008064f
C238 B.n201 VSUBS 0.008064f
C239 B.n202 VSUBS 0.008064f
C240 B.n203 VSUBS 0.008064f
C241 B.n204 VSUBS 0.008064f
C242 B.n205 VSUBS 0.008064f
C243 B.n206 VSUBS 0.008064f
C244 B.n207 VSUBS 0.008064f
C245 B.n208 VSUBS 0.008064f
C246 B.n209 VSUBS 0.008064f
C247 B.n210 VSUBS 0.008064f
C248 B.n211 VSUBS 0.008064f
C249 B.n212 VSUBS 0.008064f
C250 B.n213 VSUBS 0.008064f
C251 B.n214 VSUBS 0.008064f
C252 B.n215 VSUBS 0.008064f
C253 B.n216 VSUBS 0.008064f
C254 B.n217 VSUBS 0.008064f
C255 B.n218 VSUBS 0.018659f
C256 B.n219 VSUBS 0.008064f
C257 B.n220 VSUBS 0.008064f
C258 B.n221 VSUBS 0.008064f
C259 B.n222 VSUBS 0.008064f
C260 B.n223 VSUBS 0.008064f
C261 B.n224 VSUBS 0.008064f
C262 B.n225 VSUBS 0.008064f
C263 B.n226 VSUBS 0.008064f
C264 B.n227 VSUBS 0.008064f
C265 B.n228 VSUBS 0.008064f
C266 B.n229 VSUBS 0.008064f
C267 B.n230 VSUBS 0.008064f
C268 B.n231 VSUBS 0.008064f
C269 B.n232 VSUBS 0.008064f
C270 B.n233 VSUBS 0.008064f
C271 B.n234 VSUBS 0.008064f
C272 B.n235 VSUBS 0.008064f
C273 B.n236 VSUBS 0.008064f
C274 B.n237 VSUBS 0.008064f
C275 B.n238 VSUBS 0.008064f
C276 B.n239 VSUBS 0.008064f
C277 B.n240 VSUBS 0.008064f
C278 B.n241 VSUBS 0.008064f
C279 B.n242 VSUBS 0.008064f
C280 B.n243 VSUBS 0.008064f
C281 B.n244 VSUBS 0.008064f
C282 B.n245 VSUBS 0.008064f
C283 B.n246 VSUBS 0.008064f
C284 B.n247 VSUBS 0.008064f
C285 B.n248 VSUBS 0.008064f
C286 B.n249 VSUBS 0.008064f
C287 B.n250 VSUBS 0.008064f
C288 B.n251 VSUBS 0.008064f
C289 B.n252 VSUBS 0.008064f
C290 B.n253 VSUBS 0.008064f
C291 B.n254 VSUBS 0.008064f
C292 B.n255 VSUBS 0.008064f
C293 B.n256 VSUBS 0.008064f
C294 B.n257 VSUBS 0.008064f
C295 B.n258 VSUBS 0.008064f
C296 B.n259 VSUBS 0.008064f
C297 B.n260 VSUBS 0.008064f
C298 B.n261 VSUBS 0.008064f
C299 B.n262 VSUBS 0.008064f
C300 B.n263 VSUBS 0.008064f
C301 B.n264 VSUBS 0.008064f
C302 B.n265 VSUBS 0.008064f
C303 B.n266 VSUBS 0.008064f
C304 B.n267 VSUBS 0.008064f
C305 B.n268 VSUBS 0.008064f
C306 B.n269 VSUBS 0.008064f
C307 B.n270 VSUBS 0.008064f
C308 B.n271 VSUBS 0.008064f
C309 B.n272 VSUBS 0.008064f
C310 B.n273 VSUBS 0.008064f
C311 B.n274 VSUBS 0.008064f
C312 B.n275 VSUBS 0.008064f
C313 B.n276 VSUBS 0.008064f
C314 B.n277 VSUBS 0.008064f
C315 B.n278 VSUBS 0.008064f
C316 B.n279 VSUBS 0.008064f
C317 B.n280 VSUBS 0.008064f
C318 B.n281 VSUBS 0.008064f
C319 B.n282 VSUBS 0.008064f
C320 B.n283 VSUBS 0.008064f
C321 B.n284 VSUBS 0.008064f
C322 B.n285 VSUBS 0.008064f
C323 B.n286 VSUBS 0.008064f
C324 B.n287 VSUBS 0.008064f
C325 B.n288 VSUBS 0.008064f
C326 B.n289 VSUBS 0.008064f
C327 B.n290 VSUBS 0.008064f
C328 B.n291 VSUBS 0.008064f
C329 B.n292 VSUBS 0.008064f
C330 B.n293 VSUBS 0.008064f
C331 B.n294 VSUBS 0.008064f
C332 B.n295 VSUBS 0.008064f
C333 B.n296 VSUBS 0.008064f
C334 B.n297 VSUBS 0.008064f
C335 B.n298 VSUBS 0.008064f
C336 B.n299 VSUBS 0.008064f
C337 B.n300 VSUBS 0.008064f
C338 B.n301 VSUBS 0.008064f
C339 B.n302 VSUBS 0.008064f
C340 B.n303 VSUBS 0.008064f
C341 B.n304 VSUBS 0.008064f
C342 B.n305 VSUBS 0.008064f
C343 B.n306 VSUBS 0.008064f
C344 B.n307 VSUBS 0.008064f
C345 B.n308 VSUBS 0.008064f
C346 B.n309 VSUBS 0.008064f
C347 B.n310 VSUBS 0.008064f
C348 B.n311 VSUBS 0.008064f
C349 B.n312 VSUBS 0.008064f
C350 B.n313 VSUBS 0.008064f
C351 B.n314 VSUBS 0.008064f
C352 B.n315 VSUBS 0.008064f
C353 B.n316 VSUBS 0.008064f
C354 B.n317 VSUBS 0.008064f
C355 B.n318 VSUBS 0.008064f
C356 B.n319 VSUBS 0.008064f
C357 B.n320 VSUBS 0.008064f
C358 B.n321 VSUBS 0.008064f
C359 B.n322 VSUBS 0.008064f
C360 B.n323 VSUBS 0.008064f
C361 B.n324 VSUBS 0.008064f
C362 B.n325 VSUBS 0.008064f
C363 B.n326 VSUBS 0.008064f
C364 B.n327 VSUBS 0.008064f
C365 B.n328 VSUBS 0.008064f
C366 B.n329 VSUBS 0.008064f
C367 B.n330 VSUBS 0.008064f
C368 B.n331 VSUBS 0.008064f
C369 B.n332 VSUBS 0.008064f
C370 B.n333 VSUBS 0.008064f
C371 B.n334 VSUBS 0.008064f
C372 B.n335 VSUBS 0.008064f
C373 B.n336 VSUBS 0.008064f
C374 B.n337 VSUBS 0.008064f
C375 B.n338 VSUBS 0.008064f
C376 B.n339 VSUBS 0.008064f
C377 B.n340 VSUBS 0.008064f
C378 B.n341 VSUBS 0.008064f
C379 B.n342 VSUBS 0.008064f
C380 B.n343 VSUBS 0.008064f
C381 B.n344 VSUBS 0.008064f
C382 B.n345 VSUBS 0.008064f
C383 B.n346 VSUBS 0.008064f
C384 B.n347 VSUBS 0.008064f
C385 B.n348 VSUBS 0.008064f
C386 B.n349 VSUBS 0.008064f
C387 B.n350 VSUBS 0.008064f
C388 B.n351 VSUBS 0.008064f
C389 B.n352 VSUBS 0.008064f
C390 B.n353 VSUBS 0.018659f
C391 B.n354 VSUBS 0.019054f
C392 B.n355 VSUBS 0.019054f
C393 B.n356 VSUBS 0.008064f
C394 B.n357 VSUBS 0.008064f
C395 B.n358 VSUBS 0.008064f
C396 B.n359 VSUBS 0.008064f
C397 B.n360 VSUBS 0.008064f
C398 B.n361 VSUBS 0.008064f
C399 B.n362 VSUBS 0.008064f
C400 B.n363 VSUBS 0.008064f
C401 B.n364 VSUBS 0.008064f
C402 B.n365 VSUBS 0.008064f
C403 B.n366 VSUBS 0.008064f
C404 B.n367 VSUBS 0.008064f
C405 B.n368 VSUBS 0.008064f
C406 B.n369 VSUBS 0.008064f
C407 B.n370 VSUBS 0.008064f
C408 B.n371 VSUBS 0.008064f
C409 B.n372 VSUBS 0.008064f
C410 B.n373 VSUBS 0.008064f
C411 B.n374 VSUBS 0.008064f
C412 B.n375 VSUBS 0.008064f
C413 B.n376 VSUBS 0.008064f
C414 B.n377 VSUBS 0.008064f
C415 B.n378 VSUBS 0.008064f
C416 B.n379 VSUBS 0.008064f
C417 B.n380 VSUBS 0.008064f
C418 B.n381 VSUBS 0.008064f
C419 B.n382 VSUBS 0.008064f
C420 B.n383 VSUBS 0.008064f
C421 B.n384 VSUBS 0.008064f
C422 B.n385 VSUBS 0.008064f
C423 B.n386 VSUBS 0.008064f
C424 B.n387 VSUBS 0.008064f
C425 B.n388 VSUBS 0.008064f
C426 B.n389 VSUBS 0.008064f
C427 B.n390 VSUBS 0.008064f
C428 B.n391 VSUBS 0.008064f
C429 B.n392 VSUBS 0.008064f
C430 B.n393 VSUBS 0.008064f
C431 B.n394 VSUBS 0.008064f
C432 B.n395 VSUBS 0.008064f
C433 B.n396 VSUBS 0.008064f
C434 B.n397 VSUBS 0.008064f
C435 B.n398 VSUBS 0.008064f
C436 B.n399 VSUBS 0.008064f
C437 B.n400 VSUBS 0.008064f
C438 B.n401 VSUBS 0.008064f
C439 B.n402 VSUBS 0.008064f
C440 B.n403 VSUBS 0.008064f
C441 B.n404 VSUBS 0.008064f
C442 B.n405 VSUBS 0.008064f
C443 B.n406 VSUBS 0.008064f
C444 B.n407 VSUBS 0.008064f
C445 B.n408 VSUBS 0.008064f
C446 B.n409 VSUBS 0.008064f
C447 B.n410 VSUBS 0.008064f
C448 B.n411 VSUBS 0.008064f
C449 B.n412 VSUBS 0.008064f
C450 B.n413 VSUBS 0.008064f
C451 B.n414 VSUBS 0.008064f
C452 B.n415 VSUBS 0.008064f
C453 B.n416 VSUBS 0.008064f
C454 B.n417 VSUBS 0.008064f
C455 B.n418 VSUBS 0.008064f
C456 B.n419 VSUBS 0.008064f
C457 B.n420 VSUBS 0.008064f
C458 B.n421 VSUBS 0.008064f
C459 B.n422 VSUBS 0.008064f
C460 B.n423 VSUBS 0.008064f
C461 B.n424 VSUBS 0.008064f
C462 B.n425 VSUBS 0.005574f
C463 B.n426 VSUBS 0.018684f
C464 B.n427 VSUBS 0.006523f
C465 B.n428 VSUBS 0.008064f
C466 B.n429 VSUBS 0.008064f
C467 B.n430 VSUBS 0.008064f
C468 B.n431 VSUBS 0.008064f
C469 B.n432 VSUBS 0.008064f
C470 B.n433 VSUBS 0.008064f
C471 B.n434 VSUBS 0.008064f
C472 B.n435 VSUBS 0.008064f
C473 B.n436 VSUBS 0.008064f
C474 B.n437 VSUBS 0.008064f
C475 B.n438 VSUBS 0.008064f
C476 B.t10 VSUBS 0.298862f
C477 B.t11 VSUBS 0.350301f
C478 B.t9 VSUBS 2.85944f
C479 B.n439 VSUBS 0.558411f
C480 B.n440 VSUBS 0.328826f
C481 B.n441 VSUBS 0.018684f
C482 B.n442 VSUBS 0.006523f
C483 B.n443 VSUBS 0.008064f
C484 B.n444 VSUBS 0.008064f
C485 B.n445 VSUBS 0.008064f
C486 B.n446 VSUBS 0.008064f
C487 B.n447 VSUBS 0.008064f
C488 B.n448 VSUBS 0.008064f
C489 B.n449 VSUBS 0.008064f
C490 B.n450 VSUBS 0.008064f
C491 B.n451 VSUBS 0.008064f
C492 B.n452 VSUBS 0.008064f
C493 B.n453 VSUBS 0.008064f
C494 B.n454 VSUBS 0.008064f
C495 B.n455 VSUBS 0.008064f
C496 B.n456 VSUBS 0.008064f
C497 B.n457 VSUBS 0.008064f
C498 B.n458 VSUBS 0.008064f
C499 B.n459 VSUBS 0.008064f
C500 B.n460 VSUBS 0.008064f
C501 B.n461 VSUBS 0.008064f
C502 B.n462 VSUBS 0.008064f
C503 B.n463 VSUBS 0.008064f
C504 B.n464 VSUBS 0.008064f
C505 B.n465 VSUBS 0.008064f
C506 B.n466 VSUBS 0.008064f
C507 B.n467 VSUBS 0.008064f
C508 B.n468 VSUBS 0.008064f
C509 B.n469 VSUBS 0.008064f
C510 B.n470 VSUBS 0.008064f
C511 B.n471 VSUBS 0.008064f
C512 B.n472 VSUBS 0.008064f
C513 B.n473 VSUBS 0.008064f
C514 B.n474 VSUBS 0.008064f
C515 B.n475 VSUBS 0.008064f
C516 B.n476 VSUBS 0.008064f
C517 B.n477 VSUBS 0.008064f
C518 B.n478 VSUBS 0.008064f
C519 B.n479 VSUBS 0.008064f
C520 B.n480 VSUBS 0.008064f
C521 B.n481 VSUBS 0.008064f
C522 B.n482 VSUBS 0.008064f
C523 B.n483 VSUBS 0.008064f
C524 B.n484 VSUBS 0.008064f
C525 B.n485 VSUBS 0.008064f
C526 B.n486 VSUBS 0.008064f
C527 B.n487 VSUBS 0.008064f
C528 B.n488 VSUBS 0.008064f
C529 B.n489 VSUBS 0.008064f
C530 B.n490 VSUBS 0.008064f
C531 B.n491 VSUBS 0.008064f
C532 B.n492 VSUBS 0.008064f
C533 B.n493 VSUBS 0.008064f
C534 B.n494 VSUBS 0.008064f
C535 B.n495 VSUBS 0.008064f
C536 B.n496 VSUBS 0.008064f
C537 B.n497 VSUBS 0.008064f
C538 B.n498 VSUBS 0.008064f
C539 B.n499 VSUBS 0.008064f
C540 B.n500 VSUBS 0.008064f
C541 B.n501 VSUBS 0.008064f
C542 B.n502 VSUBS 0.008064f
C543 B.n503 VSUBS 0.008064f
C544 B.n504 VSUBS 0.008064f
C545 B.n505 VSUBS 0.008064f
C546 B.n506 VSUBS 0.008064f
C547 B.n507 VSUBS 0.008064f
C548 B.n508 VSUBS 0.008064f
C549 B.n509 VSUBS 0.008064f
C550 B.n510 VSUBS 0.008064f
C551 B.n511 VSUBS 0.008064f
C552 B.n512 VSUBS 0.008064f
C553 B.n513 VSUBS 0.008064f
C554 B.n514 VSUBS 0.019054f
C555 B.n515 VSUBS 0.019054f
C556 B.n516 VSUBS 0.018659f
C557 B.n517 VSUBS 0.008064f
C558 B.n518 VSUBS 0.008064f
C559 B.n519 VSUBS 0.008064f
C560 B.n520 VSUBS 0.008064f
C561 B.n521 VSUBS 0.008064f
C562 B.n522 VSUBS 0.008064f
C563 B.n523 VSUBS 0.008064f
C564 B.n524 VSUBS 0.008064f
C565 B.n525 VSUBS 0.008064f
C566 B.n526 VSUBS 0.008064f
C567 B.n527 VSUBS 0.008064f
C568 B.n528 VSUBS 0.008064f
C569 B.n529 VSUBS 0.008064f
C570 B.n530 VSUBS 0.008064f
C571 B.n531 VSUBS 0.008064f
C572 B.n532 VSUBS 0.008064f
C573 B.n533 VSUBS 0.008064f
C574 B.n534 VSUBS 0.008064f
C575 B.n535 VSUBS 0.008064f
C576 B.n536 VSUBS 0.008064f
C577 B.n537 VSUBS 0.008064f
C578 B.n538 VSUBS 0.008064f
C579 B.n539 VSUBS 0.008064f
C580 B.n540 VSUBS 0.008064f
C581 B.n541 VSUBS 0.008064f
C582 B.n542 VSUBS 0.008064f
C583 B.n543 VSUBS 0.008064f
C584 B.n544 VSUBS 0.008064f
C585 B.n545 VSUBS 0.008064f
C586 B.n546 VSUBS 0.008064f
C587 B.n547 VSUBS 0.008064f
C588 B.n548 VSUBS 0.008064f
C589 B.n549 VSUBS 0.008064f
C590 B.n550 VSUBS 0.008064f
C591 B.n551 VSUBS 0.008064f
C592 B.n552 VSUBS 0.008064f
C593 B.n553 VSUBS 0.008064f
C594 B.n554 VSUBS 0.008064f
C595 B.n555 VSUBS 0.008064f
C596 B.n556 VSUBS 0.008064f
C597 B.n557 VSUBS 0.008064f
C598 B.n558 VSUBS 0.008064f
C599 B.n559 VSUBS 0.008064f
C600 B.n560 VSUBS 0.008064f
C601 B.n561 VSUBS 0.008064f
C602 B.n562 VSUBS 0.008064f
C603 B.n563 VSUBS 0.008064f
C604 B.n564 VSUBS 0.008064f
C605 B.n565 VSUBS 0.008064f
C606 B.n566 VSUBS 0.008064f
C607 B.n567 VSUBS 0.008064f
C608 B.n568 VSUBS 0.008064f
C609 B.n569 VSUBS 0.008064f
C610 B.n570 VSUBS 0.008064f
C611 B.n571 VSUBS 0.008064f
C612 B.n572 VSUBS 0.008064f
C613 B.n573 VSUBS 0.008064f
C614 B.n574 VSUBS 0.008064f
C615 B.n575 VSUBS 0.008064f
C616 B.n576 VSUBS 0.008064f
C617 B.n577 VSUBS 0.008064f
C618 B.n578 VSUBS 0.008064f
C619 B.n579 VSUBS 0.008064f
C620 B.n580 VSUBS 0.008064f
C621 B.n581 VSUBS 0.008064f
C622 B.n582 VSUBS 0.008064f
C623 B.n583 VSUBS 0.008064f
C624 B.n584 VSUBS 0.008064f
C625 B.n585 VSUBS 0.008064f
C626 B.n586 VSUBS 0.008064f
C627 B.n587 VSUBS 0.008064f
C628 B.n588 VSUBS 0.008064f
C629 B.n589 VSUBS 0.008064f
C630 B.n590 VSUBS 0.008064f
C631 B.n591 VSUBS 0.008064f
C632 B.n592 VSUBS 0.008064f
C633 B.n593 VSUBS 0.008064f
C634 B.n594 VSUBS 0.008064f
C635 B.n595 VSUBS 0.008064f
C636 B.n596 VSUBS 0.008064f
C637 B.n597 VSUBS 0.008064f
C638 B.n598 VSUBS 0.008064f
C639 B.n599 VSUBS 0.008064f
C640 B.n600 VSUBS 0.008064f
C641 B.n601 VSUBS 0.008064f
C642 B.n602 VSUBS 0.008064f
C643 B.n603 VSUBS 0.008064f
C644 B.n604 VSUBS 0.008064f
C645 B.n605 VSUBS 0.008064f
C646 B.n606 VSUBS 0.008064f
C647 B.n607 VSUBS 0.008064f
C648 B.n608 VSUBS 0.008064f
C649 B.n609 VSUBS 0.008064f
C650 B.n610 VSUBS 0.008064f
C651 B.n611 VSUBS 0.008064f
C652 B.n612 VSUBS 0.008064f
C653 B.n613 VSUBS 0.008064f
C654 B.n614 VSUBS 0.008064f
C655 B.n615 VSUBS 0.008064f
C656 B.n616 VSUBS 0.008064f
C657 B.n617 VSUBS 0.008064f
C658 B.n618 VSUBS 0.008064f
C659 B.n619 VSUBS 0.008064f
C660 B.n620 VSUBS 0.008064f
C661 B.n621 VSUBS 0.008064f
C662 B.n622 VSUBS 0.008064f
C663 B.n623 VSUBS 0.008064f
C664 B.n624 VSUBS 0.008064f
C665 B.n625 VSUBS 0.008064f
C666 B.n626 VSUBS 0.008064f
C667 B.n627 VSUBS 0.008064f
C668 B.n628 VSUBS 0.008064f
C669 B.n629 VSUBS 0.008064f
C670 B.n630 VSUBS 0.008064f
C671 B.n631 VSUBS 0.008064f
C672 B.n632 VSUBS 0.008064f
C673 B.n633 VSUBS 0.008064f
C674 B.n634 VSUBS 0.008064f
C675 B.n635 VSUBS 0.008064f
C676 B.n636 VSUBS 0.008064f
C677 B.n637 VSUBS 0.008064f
C678 B.n638 VSUBS 0.008064f
C679 B.n639 VSUBS 0.008064f
C680 B.n640 VSUBS 0.008064f
C681 B.n641 VSUBS 0.008064f
C682 B.n642 VSUBS 0.008064f
C683 B.n643 VSUBS 0.008064f
C684 B.n644 VSUBS 0.008064f
C685 B.n645 VSUBS 0.008064f
C686 B.n646 VSUBS 0.008064f
C687 B.n647 VSUBS 0.008064f
C688 B.n648 VSUBS 0.008064f
C689 B.n649 VSUBS 0.008064f
C690 B.n650 VSUBS 0.008064f
C691 B.n651 VSUBS 0.008064f
C692 B.n652 VSUBS 0.008064f
C693 B.n653 VSUBS 0.008064f
C694 B.n654 VSUBS 0.008064f
C695 B.n655 VSUBS 0.008064f
C696 B.n656 VSUBS 0.008064f
C697 B.n657 VSUBS 0.008064f
C698 B.n658 VSUBS 0.008064f
C699 B.n659 VSUBS 0.008064f
C700 B.n660 VSUBS 0.008064f
C701 B.n661 VSUBS 0.008064f
C702 B.n662 VSUBS 0.008064f
C703 B.n663 VSUBS 0.008064f
C704 B.n664 VSUBS 0.008064f
C705 B.n665 VSUBS 0.008064f
C706 B.n666 VSUBS 0.008064f
C707 B.n667 VSUBS 0.008064f
C708 B.n668 VSUBS 0.008064f
C709 B.n669 VSUBS 0.008064f
C710 B.n670 VSUBS 0.008064f
C711 B.n671 VSUBS 0.008064f
C712 B.n672 VSUBS 0.008064f
C713 B.n673 VSUBS 0.008064f
C714 B.n674 VSUBS 0.008064f
C715 B.n675 VSUBS 0.008064f
C716 B.n676 VSUBS 0.008064f
C717 B.n677 VSUBS 0.008064f
C718 B.n678 VSUBS 0.008064f
C719 B.n679 VSUBS 0.008064f
C720 B.n680 VSUBS 0.008064f
C721 B.n681 VSUBS 0.008064f
C722 B.n682 VSUBS 0.008064f
C723 B.n683 VSUBS 0.008064f
C724 B.n684 VSUBS 0.008064f
C725 B.n685 VSUBS 0.008064f
C726 B.n686 VSUBS 0.008064f
C727 B.n687 VSUBS 0.008064f
C728 B.n688 VSUBS 0.008064f
C729 B.n689 VSUBS 0.008064f
C730 B.n690 VSUBS 0.008064f
C731 B.n691 VSUBS 0.008064f
C732 B.n692 VSUBS 0.008064f
C733 B.n693 VSUBS 0.008064f
C734 B.n694 VSUBS 0.008064f
C735 B.n695 VSUBS 0.008064f
C736 B.n696 VSUBS 0.008064f
C737 B.n697 VSUBS 0.008064f
C738 B.n698 VSUBS 0.008064f
C739 B.n699 VSUBS 0.008064f
C740 B.n700 VSUBS 0.008064f
C741 B.n701 VSUBS 0.008064f
C742 B.n702 VSUBS 0.008064f
C743 B.n703 VSUBS 0.008064f
C744 B.n704 VSUBS 0.008064f
C745 B.n705 VSUBS 0.008064f
C746 B.n706 VSUBS 0.008064f
C747 B.n707 VSUBS 0.008064f
C748 B.n708 VSUBS 0.008064f
C749 B.n709 VSUBS 0.008064f
C750 B.n710 VSUBS 0.008064f
C751 B.n711 VSUBS 0.008064f
C752 B.n712 VSUBS 0.008064f
C753 B.n713 VSUBS 0.008064f
C754 B.n714 VSUBS 0.008064f
C755 B.n715 VSUBS 0.008064f
C756 B.n716 VSUBS 0.008064f
C757 B.n717 VSUBS 0.008064f
C758 B.n718 VSUBS 0.008064f
C759 B.n719 VSUBS 0.008064f
C760 B.n720 VSUBS 0.008064f
C761 B.n721 VSUBS 0.008064f
C762 B.n722 VSUBS 0.008064f
C763 B.n723 VSUBS 0.019613f
C764 B.n724 VSUBS 0.0181f
C765 B.n725 VSUBS 0.019054f
C766 B.n726 VSUBS 0.008064f
C767 B.n727 VSUBS 0.008064f
C768 B.n728 VSUBS 0.008064f
C769 B.n729 VSUBS 0.008064f
C770 B.n730 VSUBS 0.008064f
C771 B.n731 VSUBS 0.008064f
C772 B.n732 VSUBS 0.008064f
C773 B.n733 VSUBS 0.008064f
C774 B.n734 VSUBS 0.008064f
C775 B.n735 VSUBS 0.008064f
C776 B.n736 VSUBS 0.008064f
C777 B.n737 VSUBS 0.008064f
C778 B.n738 VSUBS 0.008064f
C779 B.n739 VSUBS 0.008064f
C780 B.n740 VSUBS 0.008064f
C781 B.n741 VSUBS 0.008064f
C782 B.n742 VSUBS 0.008064f
C783 B.n743 VSUBS 0.008064f
C784 B.n744 VSUBS 0.008064f
C785 B.n745 VSUBS 0.008064f
C786 B.n746 VSUBS 0.008064f
C787 B.n747 VSUBS 0.008064f
C788 B.n748 VSUBS 0.008064f
C789 B.n749 VSUBS 0.008064f
C790 B.n750 VSUBS 0.008064f
C791 B.n751 VSUBS 0.008064f
C792 B.n752 VSUBS 0.008064f
C793 B.n753 VSUBS 0.008064f
C794 B.n754 VSUBS 0.008064f
C795 B.n755 VSUBS 0.008064f
C796 B.n756 VSUBS 0.008064f
C797 B.n757 VSUBS 0.008064f
C798 B.n758 VSUBS 0.008064f
C799 B.n759 VSUBS 0.008064f
C800 B.n760 VSUBS 0.008064f
C801 B.n761 VSUBS 0.008064f
C802 B.n762 VSUBS 0.008064f
C803 B.n763 VSUBS 0.008064f
C804 B.n764 VSUBS 0.008064f
C805 B.n765 VSUBS 0.008064f
C806 B.n766 VSUBS 0.008064f
C807 B.n767 VSUBS 0.008064f
C808 B.n768 VSUBS 0.008064f
C809 B.n769 VSUBS 0.008064f
C810 B.n770 VSUBS 0.008064f
C811 B.n771 VSUBS 0.008064f
C812 B.n772 VSUBS 0.008064f
C813 B.n773 VSUBS 0.008064f
C814 B.n774 VSUBS 0.008064f
C815 B.n775 VSUBS 0.008064f
C816 B.n776 VSUBS 0.008064f
C817 B.n777 VSUBS 0.008064f
C818 B.n778 VSUBS 0.008064f
C819 B.n779 VSUBS 0.008064f
C820 B.n780 VSUBS 0.008064f
C821 B.n781 VSUBS 0.008064f
C822 B.n782 VSUBS 0.008064f
C823 B.n783 VSUBS 0.008064f
C824 B.n784 VSUBS 0.008064f
C825 B.n785 VSUBS 0.008064f
C826 B.n786 VSUBS 0.008064f
C827 B.n787 VSUBS 0.008064f
C828 B.n788 VSUBS 0.008064f
C829 B.n789 VSUBS 0.008064f
C830 B.n790 VSUBS 0.008064f
C831 B.n791 VSUBS 0.008064f
C832 B.n792 VSUBS 0.008064f
C833 B.n793 VSUBS 0.008064f
C834 B.n794 VSUBS 0.008064f
C835 B.n795 VSUBS 0.005574f
C836 B.n796 VSUBS 0.018684f
C837 B.n797 VSUBS 0.006523f
C838 B.n798 VSUBS 0.008064f
C839 B.n799 VSUBS 0.008064f
C840 B.n800 VSUBS 0.008064f
C841 B.n801 VSUBS 0.008064f
C842 B.n802 VSUBS 0.008064f
C843 B.n803 VSUBS 0.008064f
C844 B.n804 VSUBS 0.008064f
C845 B.n805 VSUBS 0.008064f
C846 B.n806 VSUBS 0.008064f
C847 B.n807 VSUBS 0.008064f
C848 B.n808 VSUBS 0.008064f
C849 B.n809 VSUBS 0.006523f
C850 B.n810 VSUBS 0.008064f
C851 B.n811 VSUBS 0.008064f
C852 B.n812 VSUBS 0.008064f
C853 B.n813 VSUBS 0.008064f
C854 B.n814 VSUBS 0.008064f
C855 B.n815 VSUBS 0.008064f
C856 B.n816 VSUBS 0.008064f
C857 B.n817 VSUBS 0.008064f
C858 B.n818 VSUBS 0.008064f
C859 B.n819 VSUBS 0.008064f
C860 B.n820 VSUBS 0.008064f
C861 B.n821 VSUBS 0.008064f
C862 B.n822 VSUBS 0.008064f
C863 B.n823 VSUBS 0.008064f
C864 B.n824 VSUBS 0.008064f
C865 B.n825 VSUBS 0.008064f
C866 B.n826 VSUBS 0.008064f
C867 B.n827 VSUBS 0.008064f
C868 B.n828 VSUBS 0.008064f
C869 B.n829 VSUBS 0.008064f
C870 B.n830 VSUBS 0.008064f
C871 B.n831 VSUBS 0.008064f
C872 B.n832 VSUBS 0.008064f
C873 B.n833 VSUBS 0.008064f
C874 B.n834 VSUBS 0.008064f
C875 B.n835 VSUBS 0.008064f
C876 B.n836 VSUBS 0.008064f
C877 B.n837 VSUBS 0.008064f
C878 B.n838 VSUBS 0.008064f
C879 B.n839 VSUBS 0.008064f
C880 B.n840 VSUBS 0.008064f
C881 B.n841 VSUBS 0.008064f
C882 B.n842 VSUBS 0.008064f
C883 B.n843 VSUBS 0.008064f
C884 B.n844 VSUBS 0.008064f
C885 B.n845 VSUBS 0.008064f
C886 B.n846 VSUBS 0.008064f
C887 B.n847 VSUBS 0.008064f
C888 B.n848 VSUBS 0.008064f
C889 B.n849 VSUBS 0.008064f
C890 B.n850 VSUBS 0.008064f
C891 B.n851 VSUBS 0.008064f
C892 B.n852 VSUBS 0.008064f
C893 B.n853 VSUBS 0.008064f
C894 B.n854 VSUBS 0.008064f
C895 B.n855 VSUBS 0.008064f
C896 B.n856 VSUBS 0.008064f
C897 B.n857 VSUBS 0.008064f
C898 B.n858 VSUBS 0.008064f
C899 B.n859 VSUBS 0.008064f
C900 B.n860 VSUBS 0.008064f
C901 B.n861 VSUBS 0.008064f
C902 B.n862 VSUBS 0.008064f
C903 B.n863 VSUBS 0.008064f
C904 B.n864 VSUBS 0.008064f
C905 B.n865 VSUBS 0.008064f
C906 B.n866 VSUBS 0.008064f
C907 B.n867 VSUBS 0.008064f
C908 B.n868 VSUBS 0.008064f
C909 B.n869 VSUBS 0.008064f
C910 B.n870 VSUBS 0.008064f
C911 B.n871 VSUBS 0.008064f
C912 B.n872 VSUBS 0.008064f
C913 B.n873 VSUBS 0.008064f
C914 B.n874 VSUBS 0.008064f
C915 B.n875 VSUBS 0.008064f
C916 B.n876 VSUBS 0.008064f
C917 B.n877 VSUBS 0.008064f
C918 B.n878 VSUBS 0.008064f
C919 B.n879 VSUBS 0.008064f
C920 B.n880 VSUBS 0.008064f
C921 B.n881 VSUBS 0.019054f
C922 B.n882 VSUBS 0.019054f
C923 B.n883 VSUBS 0.018659f
C924 B.n884 VSUBS 0.008064f
C925 B.n885 VSUBS 0.008064f
C926 B.n886 VSUBS 0.008064f
C927 B.n887 VSUBS 0.008064f
C928 B.n888 VSUBS 0.008064f
C929 B.n889 VSUBS 0.008064f
C930 B.n890 VSUBS 0.008064f
C931 B.n891 VSUBS 0.008064f
C932 B.n892 VSUBS 0.008064f
C933 B.n893 VSUBS 0.008064f
C934 B.n894 VSUBS 0.008064f
C935 B.n895 VSUBS 0.008064f
C936 B.n896 VSUBS 0.008064f
C937 B.n897 VSUBS 0.008064f
C938 B.n898 VSUBS 0.008064f
C939 B.n899 VSUBS 0.008064f
C940 B.n900 VSUBS 0.008064f
C941 B.n901 VSUBS 0.008064f
C942 B.n902 VSUBS 0.008064f
C943 B.n903 VSUBS 0.008064f
C944 B.n904 VSUBS 0.008064f
C945 B.n905 VSUBS 0.008064f
C946 B.n906 VSUBS 0.008064f
C947 B.n907 VSUBS 0.008064f
C948 B.n908 VSUBS 0.008064f
C949 B.n909 VSUBS 0.008064f
C950 B.n910 VSUBS 0.008064f
C951 B.n911 VSUBS 0.008064f
C952 B.n912 VSUBS 0.008064f
C953 B.n913 VSUBS 0.008064f
C954 B.n914 VSUBS 0.008064f
C955 B.n915 VSUBS 0.008064f
C956 B.n916 VSUBS 0.008064f
C957 B.n917 VSUBS 0.008064f
C958 B.n918 VSUBS 0.008064f
C959 B.n919 VSUBS 0.008064f
C960 B.n920 VSUBS 0.008064f
C961 B.n921 VSUBS 0.008064f
C962 B.n922 VSUBS 0.008064f
C963 B.n923 VSUBS 0.008064f
C964 B.n924 VSUBS 0.008064f
C965 B.n925 VSUBS 0.008064f
C966 B.n926 VSUBS 0.008064f
C967 B.n927 VSUBS 0.008064f
C968 B.n928 VSUBS 0.008064f
C969 B.n929 VSUBS 0.008064f
C970 B.n930 VSUBS 0.008064f
C971 B.n931 VSUBS 0.008064f
C972 B.n932 VSUBS 0.008064f
C973 B.n933 VSUBS 0.008064f
C974 B.n934 VSUBS 0.008064f
C975 B.n935 VSUBS 0.008064f
C976 B.n936 VSUBS 0.008064f
C977 B.n937 VSUBS 0.008064f
C978 B.n938 VSUBS 0.008064f
C979 B.n939 VSUBS 0.008064f
C980 B.n940 VSUBS 0.008064f
C981 B.n941 VSUBS 0.008064f
C982 B.n942 VSUBS 0.008064f
C983 B.n943 VSUBS 0.008064f
C984 B.n944 VSUBS 0.008064f
C985 B.n945 VSUBS 0.008064f
C986 B.n946 VSUBS 0.008064f
C987 B.n947 VSUBS 0.008064f
C988 B.n948 VSUBS 0.008064f
C989 B.n949 VSUBS 0.008064f
C990 B.n950 VSUBS 0.008064f
C991 B.n951 VSUBS 0.008064f
C992 B.n952 VSUBS 0.008064f
C993 B.n953 VSUBS 0.008064f
C994 B.n954 VSUBS 0.008064f
C995 B.n955 VSUBS 0.008064f
C996 B.n956 VSUBS 0.008064f
C997 B.n957 VSUBS 0.008064f
C998 B.n958 VSUBS 0.008064f
C999 B.n959 VSUBS 0.008064f
C1000 B.n960 VSUBS 0.008064f
C1001 B.n961 VSUBS 0.008064f
C1002 B.n962 VSUBS 0.008064f
C1003 B.n963 VSUBS 0.008064f
C1004 B.n964 VSUBS 0.008064f
C1005 B.n965 VSUBS 0.008064f
C1006 B.n966 VSUBS 0.008064f
C1007 B.n967 VSUBS 0.008064f
C1008 B.n968 VSUBS 0.008064f
C1009 B.n969 VSUBS 0.008064f
C1010 B.n970 VSUBS 0.008064f
C1011 B.n971 VSUBS 0.008064f
C1012 B.n972 VSUBS 0.008064f
C1013 B.n973 VSUBS 0.008064f
C1014 B.n974 VSUBS 0.008064f
C1015 B.n975 VSUBS 0.008064f
C1016 B.n976 VSUBS 0.008064f
C1017 B.n977 VSUBS 0.008064f
C1018 B.n978 VSUBS 0.008064f
C1019 B.n979 VSUBS 0.008064f
C1020 B.n980 VSUBS 0.008064f
C1021 B.n981 VSUBS 0.008064f
C1022 B.n982 VSUBS 0.008064f
C1023 B.n983 VSUBS 0.008064f
C1024 B.n984 VSUBS 0.008064f
C1025 B.n985 VSUBS 0.008064f
C1026 B.n986 VSUBS 0.008064f
C1027 B.n987 VSUBS 0.018261f
C1028 VDD2.t4 VSUBS 0.364881f
C1029 VDD2.t5 VSUBS 0.364881f
C1030 VDD2.n0 VSUBS 2.98077f
C1031 VDD2.t7 VSUBS 0.364881f
C1032 VDD2.t0 VSUBS 0.364881f
C1033 VDD2.n1 VSUBS 2.98077f
C1034 VDD2.n2 VSUBS 6.02313f
C1035 VDD2.t1 VSUBS 0.364881f
C1036 VDD2.t2 VSUBS 0.364881f
C1037 VDD2.n3 VSUBS 2.9546f
C1038 VDD2.n4 VSUBS 4.94238f
C1039 VDD2.t3 VSUBS 0.364881f
C1040 VDD2.t6 VSUBS 0.364881f
C1041 VDD2.n5 VSUBS 2.98071f
C1042 VN.n0 VSUBS 0.042385f
C1043 VN.t7 VSUBS 3.31073f
C1044 VN.n1 VSUBS 0.044572f
C1045 VN.n2 VSUBS 0.022533f
C1046 VN.n3 VSUBS 0.041996f
C1047 VN.n4 VSUBS 0.022533f
C1048 VN.t0 VSUBS 3.31073f
C1049 VN.n5 VSUBS 0.041996f
C1050 VN.n6 VSUBS 0.022533f
C1051 VN.n7 VSUBS 0.041996f
C1052 VN.t3 VSUBS 3.66167f
C1053 VN.n8 VSUBS 1.17785f
C1054 VN.t2 VSUBS 3.31073f
C1055 VN.n9 VSUBS 1.23458f
C1056 VN.n10 VSUBS 0.034324f
C1057 VN.n11 VSUBS 0.293971f
C1058 VN.n12 VSUBS 0.022533f
C1059 VN.n13 VSUBS 0.022533f
C1060 VN.n14 VSUBS 0.041996f
C1061 VN.n15 VSUBS 0.032895f
C1062 VN.n16 VSUBS 0.032895f
C1063 VN.n17 VSUBS 0.022533f
C1064 VN.n18 VSUBS 0.022533f
C1065 VN.n19 VSUBS 0.022533f
C1066 VN.n20 VSUBS 0.041996f
C1067 VN.n21 VSUBS 0.034324f
C1068 VN.n22 VSUBS 1.15097f
C1069 VN.n23 VSUBS 0.028933f
C1070 VN.n24 VSUBS 0.022533f
C1071 VN.n25 VSUBS 0.022533f
C1072 VN.n26 VSUBS 0.022533f
C1073 VN.n27 VSUBS 0.041996f
C1074 VN.n28 VSUBS 0.040454f
C1075 VN.n29 VSUBS 0.02276f
C1076 VN.n30 VSUBS 0.022533f
C1077 VN.n31 VSUBS 0.022533f
C1078 VN.n32 VSUBS 0.022533f
C1079 VN.n33 VSUBS 0.041996f
C1080 VN.n34 VSUBS 0.039715f
C1081 VN.n35 VSUBS 1.24894f
C1082 VN.n36 VSUBS 0.068167f
C1083 VN.n37 VSUBS 0.042385f
C1084 VN.t6 VSUBS 3.31073f
C1085 VN.n38 VSUBS 0.044572f
C1086 VN.n39 VSUBS 0.022533f
C1087 VN.n40 VSUBS 0.041996f
C1088 VN.n41 VSUBS 0.022533f
C1089 VN.t5 VSUBS 3.31073f
C1090 VN.n42 VSUBS 0.041996f
C1091 VN.n43 VSUBS 0.022533f
C1092 VN.n44 VSUBS 0.041996f
C1093 VN.t1 VSUBS 3.66167f
C1094 VN.n45 VSUBS 1.17785f
C1095 VN.t4 VSUBS 3.31073f
C1096 VN.n46 VSUBS 1.23458f
C1097 VN.n47 VSUBS 0.034324f
C1098 VN.n48 VSUBS 0.293971f
C1099 VN.n49 VSUBS 0.022533f
C1100 VN.n50 VSUBS 0.022533f
C1101 VN.n51 VSUBS 0.041996f
C1102 VN.n52 VSUBS 0.032895f
C1103 VN.n53 VSUBS 0.032895f
C1104 VN.n54 VSUBS 0.022533f
C1105 VN.n55 VSUBS 0.022533f
C1106 VN.n56 VSUBS 0.022533f
C1107 VN.n57 VSUBS 0.041996f
C1108 VN.n58 VSUBS 0.034324f
C1109 VN.n59 VSUBS 1.15097f
C1110 VN.n60 VSUBS 0.028933f
C1111 VN.n61 VSUBS 0.022533f
C1112 VN.n62 VSUBS 0.022533f
C1113 VN.n63 VSUBS 0.022533f
C1114 VN.n64 VSUBS 0.041996f
C1115 VN.n65 VSUBS 0.040454f
C1116 VN.n66 VSUBS 0.02276f
C1117 VN.n67 VSUBS 0.022533f
C1118 VN.n68 VSUBS 0.022533f
C1119 VN.n69 VSUBS 0.022533f
C1120 VN.n70 VSUBS 0.041996f
C1121 VN.n71 VSUBS 0.039715f
C1122 VN.n72 VSUBS 1.24894f
C1123 VN.n73 VSUBS 1.6196f
C1124 VDD1.t2 VSUBS 0.364606f
C1125 VDD1.t7 VSUBS 0.364606f
C1126 VDD1.n0 VSUBS 2.98048f
C1127 VDD1.t6 VSUBS 0.364606f
C1128 VDD1.t5 VSUBS 0.364606f
C1129 VDD1.n1 VSUBS 2.97852f
C1130 VDD1.t1 VSUBS 0.364606f
C1131 VDD1.t0 VSUBS 0.364606f
C1132 VDD1.n2 VSUBS 2.97852f
C1133 VDD1.n3 VSUBS 6.0857f
C1134 VDD1.t3 VSUBS 0.364606f
C1135 VDD1.t4 VSUBS 0.364606f
C1136 VDD1.n4 VSUBS 2.95236f
C1137 VDD1.n5 VSUBS 4.9799f
C1138 VTAIL.t2 VSUBS 0.283337f
C1139 VTAIL.t3 VSUBS 0.283337f
C1140 VTAIL.n0 VSUBS 2.16324f
C1141 VTAIL.n1 VSUBS 0.858699f
C1142 VTAIL.n2 VSUBS 0.027453f
C1143 VTAIL.n3 VSUBS 0.025375f
C1144 VTAIL.n4 VSUBS 0.014037f
C1145 VTAIL.n5 VSUBS 0.032229f
C1146 VTAIL.n6 VSUBS 0.014438f
C1147 VTAIL.n7 VSUBS 0.025375f
C1148 VTAIL.n8 VSUBS 0.013636f
C1149 VTAIL.n9 VSUBS 0.032229f
C1150 VTAIL.n10 VSUBS 0.014438f
C1151 VTAIL.n11 VSUBS 0.025375f
C1152 VTAIL.n12 VSUBS 0.013636f
C1153 VTAIL.n13 VSUBS 0.032229f
C1154 VTAIL.n14 VSUBS 0.014438f
C1155 VTAIL.n15 VSUBS 0.025375f
C1156 VTAIL.n16 VSUBS 0.013636f
C1157 VTAIL.n17 VSUBS 0.032229f
C1158 VTAIL.n18 VSUBS 0.014438f
C1159 VTAIL.n19 VSUBS 0.025375f
C1160 VTAIL.n20 VSUBS 0.013636f
C1161 VTAIL.n21 VSUBS 0.032229f
C1162 VTAIL.n22 VSUBS 0.014438f
C1163 VTAIL.n23 VSUBS 0.025375f
C1164 VTAIL.n24 VSUBS 0.013636f
C1165 VTAIL.n25 VSUBS 0.024172f
C1166 VTAIL.n26 VSUBS 0.020503f
C1167 VTAIL.t5 VSUBS 0.068942f
C1168 VTAIL.n27 VSUBS 0.172362f
C1169 VTAIL.n28 VSUBS 1.52003f
C1170 VTAIL.n29 VSUBS 0.013636f
C1171 VTAIL.n30 VSUBS 0.014438f
C1172 VTAIL.n31 VSUBS 0.032229f
C1173 VTAIL.n32 VSUBS 0.032229f
C1174 VTAIL.n33 VSUBS 0.014438f
C1175 VTAIL.n34 VSUBS 0.013636f
C1176 VTAIL.n35 VSUBS 0.025375f
C1177 VTAIL.n36 VSUBS 0.025375f
C1178 VTAIL.n37 VSUBS 0.013636f
C1179 VTAIL.n38 VSUBS 0.014438f
C1180 VTAIL.n39 VSUBS 0.032229f
C1181 VTAIL.n40 VSUBS 0.032229f
C1182 VTAIL.n41 VSUBS 0.014438f
C1183 VTAIL.n42 VSUBS 0.013636f
C1184 VTAIL.n43 VSUBS 0.025375f
C1185 VTAIL.n44 VSUBS 0.025375f
C1186 VTAIL.n45 VSUBS 0.013636f
C1187 VTAIL.n46 VSUBS 0.014438f
C1188 VTAIL.n47 VSUBS 0.032229f
C1189 VTAIL.n48 VSUBS 0.032229f
C1190 VTAIL.n49 VSUBS 0.014438f
C1191 VTAIL.n50 VSUBS 0.013636f
C1192 VTAIL.n51 VSUBS 0.025375f
C1193 VTAIL.n52 VSUBS 0.025375f
C1194 VTAIL.n53 VSUBS 0.013636f
C1195 VTAIL.n54 VSUBS 0.014438f
C1196 VTAIL.n55 VSUBS 0.032229f
C1197 VTAIL.n56 VSUBS 0.032229f
C1198 VTAIL.n57 VSUBS 0.014438f
C1199 VTAIL.n58 VSUBS 0.013636f
C1200 VTAIL.n59 VSUBS 0.025375f
C1201 VTAIL.n60 VSUBS 0.025375f
C1202 VTAIL.n61 VSUBS 0.013636f
C1203 VTAIL.n62 VSUBS 0.014438f
C1204 VTAIL.n63 VSUBS 0.032229f
C1205 VTAIL.n64 VSUBS 0.032229f
C1206 VTAIL.n65 VSUBS 0.014438f
C1207 VTAIL.n66 VSUBS 0.013636f
C1208 VTAIL.n67 VSUBS 0.025375f
C1209 VTAIL.n68 VSUBS 0.025375f
C1210 VTAIL.n69 VSUBS 0.013636f
C1211 VTAIL.n70 VSUBS 0.013636f
C1212 VTAIL.n71 VSUBS 0.014438f
C1213 VTAIL.n72 VSUBS 0.032229f
C1214 VTAIL.n73 VSUBS 0.032229f
C1215 VTAIL.n74 VSUBS 0.076563f
C1216 VTAIL.n75 VSUBS 0.014037f
C1217 VTAIL.n76 VSUBS 0.013636f
C1218 VTAIL.n77 VSUBS 0.065933f
C1219 VTAIL.n78 VSUBS 0.03865f
C1220 VTAIL.n79 VSUBS 0.355316f
C1221 VTAIL.n80 VSUBS 0.027453f
C1222 VTAIL.n81 VSUBS 0.025375f
C1223 VTAIL.n82 VSUBS 0.014037f
C1224 VTAIL.n83 VSUBS 0.032229f
C1225 VTAIL.n84 VSUBS 0.014438f
C1226 VTAIL.n85 VSUBS 0.025375f
C1227 VTAIL.n86 VSUBS 0.013636f
C1228 VTAIL.n87 VSUBS 0.032229f
C1229 VTAIL.n88 VSUBS 0.014438f
C1230 VTAIL.n89 VSUBS 0.025375f
C1231 VTAIL.n90 VSUBS 0.013636f
C1232 VTAIL.n91 VSUBS 0.032229f
C1233 VTAIL.n92 VSUBS 0.014438f
C1234 VTAIL.n93 VSUBS 0.025375f
C1235 VTAIL.n94 VSUBS 0.013636f
C1236 VTAIL.n95 VSUBS 0.032229f
C1237 VTAIL.n96 VSUBS 0.014438f
C1238 VTAIL.n97 VSUBS 0.025375f
C1239 VTAIL.n98 VSUBS 0.013636f
C1240 VTAIL.n99 VSUBS 0.032229f
C1241 VTAIL.n100 VSUBS 0.014438f
C1242 VTAIL.n101 VSUBS 0.025375f
C1243 VTAIL.n102 VSUBS 0.013636f
C1244 VTAIL.n103 VSUBS 0.024172f
C1245 VTAIL.n104 VSUBS 0.020503f
C1246 VTAIL.t11 VSUBS 0.068942f
C1247 VTAIL.n105 VSUBS 0.172362f
C1248 VTAIL.n106 VSUBS 1.52003f
C1249 VTAIL.n107 VSUBS 0.013636f
C1250 VTAIL.n108 VSUBS 0.014438f
C1251 VTAIL.n109 VSUBS 0.032229f
C1252 VTAIL.n110 VSUBS 0.032229f
C1253 VTAIL.n111 VSUBS 0.014438f
C1254 VTAIL.n112 VSUBS 0.013636f
C1255 VTAIL.n113 VSUBS 0.025375f
C1256 VTAIL.n114 VSUBS 0.025375f
C1257 VTAIL.n115 VSUBS 0.013636f
C1258 VTAIL.n116 VSUBS 0.014438f
C1259 VTAIL.n117 VSUBS 0.032229f
C1260 VTAIL.n118 VSUBS 0.032229f
C1261 VTAIL.n119 VSUBS 0.014438f
C1262 VTAIL.n120 VSUBS 0.013636f
C1263 VTAIL.n121 VSUBS 0.025375f
C1264 VTAIL.n122 VSUBS 0.025375f
C1265 VTAIL.n123 VSUBS 0.013636f
C1266 VTAIL.n124 VSUBS 0.014438f
C1267 VTAIL.n125 VSUBS 0.032229f
C1268 VTAIL.n126 VSUBS 0.032229f
C1269 VTAIL.n127 VSUBS 0.014438f
C1270 VTAIL.n128 VSUBS 0.013636f
C1271 VTAIL.n129 VSUBS 0.025375f
C1272 VTAIL.n130 VSUBS 0.025375f
C1273 VTAIL.n131 VSUBS 0.013636f
C1274 VTAIL.n132 VSUBS 0.014438f
C1275 VTAIL.n133 VSUBS 0.032229f
C1276 VTAIL.n134 VSUBS 0.032229f
C1277 VTAIL.n135 VSUBS 0.014438f
C1278 VTAIL.n136 VSUBS 0.013636f
C1279 VTAIL.n137 VSUBS 0.025375f
C1280 VTAIL.n138 VSUBS 0.025375f
C1281 VTAIL.n139 VSUBS 0.013636f
C1282 VTAIL.n140 VSUBS 0.014438f
C1283 VTAIL.n141 VSUBS 0.032229f
C1284 VTAIL.n142 VSUBS 0.032229f
C1285 VTAIL.n143 VSUBS 0.014438f
C1286 VTAIL.n144 VSUBS 0.013636f
C1287 VTAIL.n145 VSUBS 0.025375f
C1288 VTAIL.n146 VSUBS 0.025375f
C1289 VTAIL.n147 VSUBS 0.013636f
C1290 VTAIL.n148 VSUBS 0.013636f
C1291 VTAIL.n149 VSUBS 0.014438f
C1292 VTAIL.n150 VSUBS 0.032229f
C1293 VTAIL.n151 VSUBS 0.032229f
C1294 VTAIL.n152 VSUBS 0.076563f
C1295 VTAIL.n153 VSUBS 0.014037f
C1296 VTAIL.n154 VSUBS 0.013636f
C1297 VTAIL.n155 VSUBS 0.065933f
C1298 VTAIL.n156 VSUBS 0.03865f
C1299 VTAIL.n157 VSUBS 0.355316f
C1300 VTAIL.t8 VSUBS 0.283337f
C1301 VTAIL.t10 VSUBS 0.283337f
C1302 VTAIL.n158 VSUBS 2.16324f
C1303 VTAIL.n159 VSUBS 1.14505f
C1304 VTAIL.n160 VSUBS 0.027453f
C1305 VTAIL.n161 VSUBS 0.025375f
C1306 VTAIL.n162 VSUBS 0.014037f
C1307 VTAIL.n163 VSUBS 0.032229f
C1308 VTAIL.n164 VSUBS 0.014438f
C1309 VTAIL.n165 VSUBS 0.025375f
C1310 VTAIL.n166 VSUBS 0.013636f
C1311 VTAIL.n167 VSUBS 0.032229f
C1312 VTAIL.n168 VSUBS 0.014438f
C1313 VTAIL.n169 VSUBS 0.025375f
C1314 VTAIL.n170 VSUBS 0.013636f
C1315 VTAIL.n171 VSUBS 0.032229f
C1316 VTAIL.n172 VSUBS 0.014438f
C1317 VTAIL.n173 VSUBS 0.025375f
C1318 VTAIL.n174 VSUBS 0.013636f
C1319 VTAIL.n175 VSUBS 0.032229f
C1320 VTAIL.n176 VSUBS 0.014438f
C1321 VTAIL.n177 VSUBS 0.025375f
C1322 VTAIL.n178 VSUBS 0.013636f
C1323 VTAIL.n179 VSUBS 0.032229f
C1324 VTAIL.n180 VSUBS 0.014438f
C1325 VTAIL.n181 VSUBS 0.025375f
C1326 VTAIL.n182 VSUBS 0.013636f
C1327 VTAIL.n183 VSUBS 0.024172f
C1328 VTAIL.n184 VSUBS 0.020503f
C1329 VTAIL.t9 VSUBS 0.068942f
C1330 VTAIL.n185 VSUBS 0.172362f
C1331 VTAIL.n186 VSUBS 1.52003f
C1332 VTAIL.n187 VSUBS 0.013636f
C1333 VTAIL.n188 VSUBS 0.014438f
C1334 VTAIL.n189 VSUBS 0.032229f
C1335 VTAIL.n190 VSUBS 0.032229f
C1336 VTAIL.n191 VSUBS 0.014438f
C1337 VTAIL.n192 VSUBS 0.013636f
C1338 VTAIL.n193 VSUBS 0.025375f
C1339 VTAIL.n194 VSUBS 0.025375f
C1340 VTAIL.n195 VSUBS 0.013636f
C1341 VTAIL.n196 VSUBS 0.014438f
C1342 VTAIL.n197 VSUBS 0.032229f
C1343 VTAIL.n198 VSUBS 0.032229f
C1344 VTAIL.n199 VSUBS 0.014438f
C1345 VTAIL.n200 VSUBS 0.013636f
C1346 VTAIL.n201 VSUBS 0.025375f
C1347 VTAIL.n202 VSUBS 0.025375f
C1348 VTAIL.n203 VSUBS 0.013636f
C1349 VTAIL.n204 VSUBS 0.014438f
C1350 VTAIL.n205 VSUBS 0.032229f
C1351 VTAIL.n206 VSUBS 0.032229f
C1352 VTAIL.n207 VSUBS 0.014438f
C1353 VTAIL.n208 VSUBS 0.013636f
C1354 VTAIL.n209 VSUBS 0.025375f
C1355 VTAIL.n210 VSUBS 0.025375f
C1356 VTAIL.n211 VSUBS 0.013636f
C1357 VTAIL.n212 VSUBS 0.014438f
C1358 VTAIL.n213 VSUBS 0.032229f
C1359 VTAIL.n214 VSUBS 0.032229f
C1360 VTAIL.n215 VSUBS 0.014438f
C1361 VTAIL.n216 VSUBS 0.013636f
C1362 VTAIL.n217 VSUBS 0.025375f
C1363 VTAIL.n218 VSUBS 0.025375f
C1364 VTAIL.n219 VSUBS 0.013636f
C1365 VTAIL.n220 VSUBS 0.014438f
C1366 VTAIL.n221 VSUBS 0.032229f
C1367 VTAIL.n222 VSUBS 0.032229f
C1368 VTAIL.n223 VSUBS 0.014438f
C1369 VTAIL.n224 VSUBS 0.013636f
C1370 VTAIL.n225 VSUBS 0.025375f
C1371 VTAIL.n226 VSUBS 0.025375f
C1372 VTAIL.n227 VSUBS 0.013636f
C1373 VTAIL.n228 VSUBS 0.013636f
C1374 VTAIL.n229 VSUBS 0.014438f
C1375 VTAIL.n230 VSUBS 0.032229f
C1376 VTAIL.n231 VSUBS 0.032229f
C1377 VTAIL.n232 VSUBS 0.076563f
C1378 VTAIL.n233 VSUBS 0.014037f
C1379 VTAIL.n234 VSUBS 0.013636f
C1380 VTAIL.n235 VSUBS 0.065933f
C1381 VTAIL.n236 VSUBS 0.03865f
C1382 VTAIL.n237 VSUBS 1.94867f
C1383 VTAIL.n238 VSUBS 0.027453f
C1384 VTAIL.n239 VSUBS 0.025375f
C1385 VTAIL.n240 VSUBS 0.014037f
C1386 VTAIL.n241 VSUBS 0.032229f
C1387 VTAIL.n242 VSUBS 0.013636f
C1388 VTAIL.n243 VSUBS 0.014438f
C1389 VTAIL.n244 VSUBS 0.025375f
C1390 VTAIL.n245 VSUBS 0.013636f
C1391 VTAIL.n246 VSUBS 0.032229f
C1392 VTAIL.n247 VSUBS 0.014438f
C1393 VTAIL.n248 VSUBS 0.025375f
C1394 VTAIL.n249 VSUBS 0.013636f
C1395 VTAIL.n250 VSUBS 0.032229f
C1396 VTAIL.n251 VSUBS 0.014438f
C1397 VTAIL.n252 VSUBS 0.025375f
C1398 VTAIL.n253 VSUBS 0.013636f
C1399 VTAIL.n254 VSUBS 0.032229f
C1400 VTAIL.n255 VSUBS 0.014438f
C1401 VTAIL.n256 VSUBS 0.025375f
C1402 VTAIL.n257 VSUBS 0.013636f
C1403 VTAIL.n258 VSUBS 0.032229f
C1404 VTAIL.n259 VSUBS 0.014438f
C1405 VTAIL.n260 VSUBS 0.025375f
C1406 VTAIL.n261 VSUBS 0.013636f
C1407 VTAIL.n262 VSUBS 0.024172f
C1408 VTAIL.n263 VSUBS 0.020503f
C1409 VTAIL.t1 VSUBS 0.068942f
C1410 VTAIL.n264 VSUBS 0.172362f
C1411 VTAIL.n265 VSUBS 1.52003f
C1412 VTAIL.n266 VSUBS 0.013636f
C1413 VTAIL.n267 VSUBS 0.014438f
C1414 VTAIL.n268 VSUBS 0.032229f
C1415 VTAIL.n269 VSUBS 0.032229f
C1416 VTAIL.n270 VSUBS 0.014438f
C1417 VTAIL.n271 VSUBS 0.013636f
C1418 VTAIL.n272 VSUBS 0.025375f
C1419 VTAIL.n273 VSUBS 0.025375f
C1420 VTAIL.n274 VSUBS 0.013636f
C1421 VTAIL.n275 VSUBS 0.014438f
C1422 VTAIL.n276 VSUBS 0.032229f
C1423 VTAIL.n277 VSUBS 0.032229f
C1424 VTAIL.n278 VSUBS 0.014438f
C1425 VTAIL.n279 VSUBS 0.013636f
C1426 VTAIL.n280 VSUBS 0.025375f
C1427 VTAIL.n281 VSUBS 0.025375f
C1428 VTAIL.n282 VSUBS 0.013636f
C1429 VTAIL.n283 VSUBS 0.014438f
C1430 VTAIL.n284 VSUBS 0.032229f
C1431 VTAIL.n285 VSUBS 0.032229f
C1432 VTAIL.n286 VSUBS 0.014438f
C1433 VTAIL.n287 VSUBS 0.013636f
C1434 VTAIL.n288 VSUBS 0.025375f
C1435 VTAIL.n289 VSUBS 0.025375f
C1436 VTAIL.n290 VSUBS 0.013636f
C1437 VTAIL.n291 VSUBS 0.014438f
C1438 VTAIL.n292 VSUBS 0.032229f
C1439 VTAIL.n293 VSUBS 0.032229f
C1440 VTAIL.n294 VSUBS 0.014438f
C1441 VTAIL.n295 VSUBS 0.013636f
C1442 VTAIL.n296 VSUBS 0.025375f
C1443 VTAIL.n297 VSUBS 0.025375f
C1444 VTAIL.n298 VSUBS 0.013636f
C1445 VTAIL.n299 VSUBS 0.014438f
C1446 VTAIL.n300 VSUBS 0.032229f
C1447 VTAIL.n301 VSUBS 0.032229f
C1448 VTAIL.n302 VSUBS 0.014438f
C1449 VTAIL.n303 VSUBS 0.013636f
C1450 VTAIL.n304 VSUBS 0.025375f
C1451 VTAIL.n305 VSUBS 0.025375f
C1452 VTAIL.n306 VSUBS 0.013636f
C1453 VTAIL.n307 VSUBS 0.014438f
C1454 VTAIL.n308 VSUBS 0.032229f
C1455 VTAIL.n309 VSUBS 0.032229f
C1456 VTAIL.n310 VSUBS 0.076563f
C1457 VTAIL.n311 VSUBS 0.014037f
C1458 VTAIL.n312 VSUBS 0.013636f
C1459 VTAIL.n313 VSUBS 0.065933f
C1460 VTAIL.n314 VSUBS 0.03865f
C1461 VTAIL.n315 VSUBS 1.94867f
C1462 VTAIL.t4 VSUBS 0.283337f
C1463 VTAIL.t0 VSUBS 0.283337f
C1464 VTAIL.n316 VSUBS 2.16326f
C1465 VTAIL.n317 VSUBS 1.14504f
C1466 VTAIL.n318 VSUBS 0.027453f
C1467 VTAIL.n319 VSUBS 0.025375f
C1468 VTAIL.n320 VSUBS 0.014037f
C1469 VTAIL.n321 VSUBS 0.032229f
C1470 VTAIL.n322 VSUBS 0.013636f
C1471 VTAIL.n323 VSUBS 0.014438f
C1472 VTAIL.n324 VSUBS 0.025375f
C1473 VTAIL.n325 VSUBS 0.013636f
C1474 VTAIL.n326 VSUBS 0.032229f
C1475 VTAIL.n327 VSUBS 0.014438f
C1476 VTAIL.n328 VSUBS 0.025375f
C1477 VTAIL.n329 VSUBS 0.013636f
C1478 VTAIL.n330 VSUBS 0.032229f
C1479 VTAIL.n331 VSUBS 0.014438f
C1480 VTAIL.n332 VSUBS 0.025375f
C1481 VTAIL.n333 VSUBS 0.013636f
C1482 VTAIL.n334 VSUBS 0.032229f
C1483 VTAIL.n335 VSUBS 0.014438f
C1484 VTAIL.n336 VSUBS 0.025375f
C1485 VTAIL.n337 VSUBS 0.013636f
C1486 VTAIL.n338 VSUBS 0.032229f
C1487 VTAIL.n339 VSUBS 0.014438f
C1488 VTAIL.n340 VSUBS 0.025375f
C1489 VTAIL.n341 VSUBS 0.013636f
C1490 VTAIL.n342 VSUBS 0.024172f
C1491 VTAIL.n343 VSUBS 0.020503f
C1492 VTAIL.t7 VSUBS 0.068942f
C1493 VTAIL.n344 VSUBS 0.172362f
C1494 VTAIL.n345 VSUBS 1.52003f
C1495 VTAIL.n346 VSUBS 0.013636f
C1496 VTAIL.n347 VSUBS 0.014438f
C1497 VTAIL.n348 VSUBS 0.032229f
C1498 VTAIL.n349 VSUBS 0.032229f
C1499 VTAIL.n350 VSUBS 0.014438f
C1500 VTAIL.n351 VSUBS 0.013636f
C1501 VTAIL.n352 VSUBS 0.025375f
C1502 VTAIL.n353 VSUBS 0.025375f
C1503 VTAIL.n354 VSUBS 0.013636f
C1504 VTAIL.n355 VSUBS 0.014438f
C1505 VTAIL.n356 VSUBS 0.032229f
C1506 VTAIL.n357 VSUBS 0.032229f
C1507 VTAIL.n358 VSUBS 0.014438f
C1508 VTAIL.n359 VSUBS 0.013636f
C1509 VTAIL.n360 VSUBS 0.025375f
C1510 VTAIL.n361 VSUBS 0.025375f
C1511 VTAIL.n362 VSUBS 0.013636f
C1512 VTAIL.n363 VSUBS 0.014438f
C1513 VTAIL.n364 VSUBS 0.032229f
C1514 VTAIL.n365 VSUBS 0.032229f
C1515 VTAIL.n366 VSUBS 0.014438f
C1516 VTAIL.n367 VSUBS 0.013636f
C1517 VTAIL.n368 VSUBS 0.025375f
C1518 VTAIL.n369 VSUBS 0.025375f
C1519 VTAIL.n370 VSUBS 0.013636f
C1520 VTAIL.n371 VSUBS 0.014438f
C1521 VTAIL.n372 VSUBS 0.032229f
C1522 VTAIL.n373 VSUBS 0.032229f
C1523 VTAIL.n374 VSUBS 0.014438f
C1524 VTAIL.n375 VSUBS 0.013636f
C1525 VTAIL.n376 VSUBS 0.025375f
C1526 VTAIL.n377 VSUBS 0.025375f
C1527 VTAIL.n378 VSUBS 0.013636f
C1528 VTAIL.n379 VSUBS 0.014438f
C1529 VTAIL.n380 VSUBS 0.032229f
C1530 VTAIL.n381 VSUBS 0.032229f
C1531 VTAIL.n382 VSUBS 0.014438f
C1532 VTAIL.n383 VSUBS 0.013636f
C1533 VTAIL.n384 VSUBS 0.025375f
C1534 VTAIL.n385 VSUBS 0.025375f
C1535 VTAIL.n386 VSUBS 0.013636f
C1536 VTAIL.n387 VSUBS 0.014438f
C1537 VTAIL.n388 VSUBS 0.032229f
C1538 VTAIL.n389 VSUBS 0.032229f
C1539 VTAIL.n390 VSUBS 0.076563f
C1540 VTAIL.n391 VSUBS 0.014037f
C1541 VTAIL.n392 VSUBS 0.013636f
C1542 VTAIL.n393 VSUBS 0.065933f
C1543 VTAIL.n394 VSUBS 0.03865f
C1544 VTAIL.n395 VSUBS 0.355316f
C1545 VTAIL.n396 VSUBS 0.027453f
C1546 VTAIL.n397 VSUBS 0.025375f
C1547 VTAIL.n398 VSUBS 0.014037f
C1548 VTAIL.n399 VSUBS 0.032229f
C1549 VTAIL.n400 VSUBS 0.013636f
C1550 VTAIL.n401 VSUBS 0.014438f
C1551 VTAIL.n402 VSUBS 0.025375f
C1552 VTAIL.n403 VSUBS 0.013636f
C1553 VTAIL.n404 VSUBS 0.032229f
C1554 VTAIL.n405 VSUBS 0.014438f
C1555 VTAIL.n406 VSUBS 0.025375f
C1556 VTAIL.n407 VSUBS 0.013636f
C1557 VTAIL.n408 VSUBS 0.032229f
C1558 VTAIL.n409 VSUBS 0.014438f
C1559 VTAIL.n410 VSUBS 0.025375f
C1560 VTAIL.n411 VSUBS 0.013636f
C1561 VTAIL.n412 VSUBS 0.032229f
C1562 VTAIL.n413 VSUBS 0.014438f
C1563 VTAIL.n414 VSUBS 0.025375f
C1564 VTAIL.n415 VSUBS 0.013636f
C1565 VTAIL.n416 VSUBS 0.032229f
C1566 VTAIL.n417 VSUBS 0.014438f
C1567 VTAIL.n418 VSUBS 0.025375f
C1568 VTAIL.n419 VSUBS 0.013636f
C1569 VTAIL.n420 VSUBS 0.024172f
C1570 VTAIL.n421 VSUBS 0.020503f
C1571 VTAIL.t12 VSUBS 0.068942f
C1572 VTAIL.n422 VSUBS 0.172362f
C1573 VTAIL.n423 VSUBS 1.52003f
C1574 VTAIL.n424 VSUBS 0.013636f
C1575 VTAIL.n425 VSUBS 0.014438f
C1576 VTAIL.n426 VSUBS 0.032229f
C1577 VTAIL.n427 VSUBS 0.032229f
C1578 VTAIL.n428 VSUBS 0.014438f
C1579 VTAIL.n429 VSUBS 0.013636f
C1580 VTAIL.n430 VSUBS 0.025375f
C1581 VTAIL.n431 VSUBS 0.025375f
C1582 VTAIL.n432 VSUBS 0.013636f
C1583 VTAIL.n433 VSUBS 0.014438f
C1584 VTAIL.n434 VSUBS 0.032229f
C1585 VTAIL.n435 VSUBS 0.032229f
C1586 VTAIL.n436 VSUBS 0.014438f
C1587 VTAIL.n437 VSUBS 0.013636f
C1588 VTAIL.n438 VSUBS 0.025375f
C1589 VTAIL.n439 VSUBS 0.025375f
C1590 VTAIL.n440 VSUBS 0.013636f
C1591 VTAIL.n441 VSUBS 0.014438f
C1592 VTAIL.n442 VSUBS 0.032229f
C1593 VTAIL.n443 VSUBS 0.032229f
C1594 VTAIL.n444 VSUBS 0.014438f
C1595 VTAIL.n445 VSUBS 0.013636f
C1596 VTAIL.n446 VSUBS 0.025375f
C1597 VTAIL.n447 VSUBS 0.025375f
C1598 VTAIL.n448 VSUBS 0.013636f
C1599 VTAIL.n449 VSUBS 0.014438f
C1600 VTAIL.n450 VSUBS 0.032229f
C1601 VTAIL.n451 VSUBS 0.032229f
C1602 VTAIL.n452 VSUBS 0.014438f
C1603 VTAIL.n453 VSUBS 0.013636f
C1604 VTAIL.n454 VSUBS 0.025375f
C1605 VTAIL.n455 VSUBS 0.025375f
C1606 VTAIL.n456 VSUBS 0.013636f
C1607 VTAIL.n457 VSUBS 0.014438f
C1608 VTAIL.n458 VSUBS 0.032229f
C1609 VTAIL.n459 VSUBS 0.032229f
C1610 VTAIL.n460 VSUBS 0.014438f
C1611 VTAIL.n461 VSUBS 0.013636f
C1612 VTAIL.n462 VSUBS 0.025375f
C1613 VTAIL.n463 VSUBS 0.025375f
C1614 VTAIL.n464 VSUBS 0.013636f
C1615 VTAIL.n465 VSUBS 0.014438f
C1616 VTAIL.n466 VSUBS 0.032229f
C1617 VTAIL.n467 VSUBS 0.032229f
C1618 VTAIL.n468 VSUBS 0.076563f
C1619 VTAIL.n469 VSUBS 0.014037f
C1620 VTAIL.n470 VSUBS 0.013636f
C1621 VTAIL.n471 VSUBS 0.065933f
C1622 VTAIL.n472 VSUBS 0.03865f
C1623 VTAIL.n473 VSUBS 0.355316f
C1624 VTAIL.t14 VSUBS 0.283337f
C1625 VTAIL.t15 VSUBS 0.283337f
C1626 VTAIL.n474 VSUBS 2.16326f
C1627 VTAIL.n475 VSUBS 1.14504f
C1628 VTAIL.n476 VSUBS 0.027453f
C1629 VTAIL.n477 VSUBS 0.025375f
C1630 VTAIL.n478 VSUBS 0.014037f
C1631 VTAIL.n479 VSUBS 0.032229f
C1632 VTAIL.n480 VSUBS 0.013636f
C1633 VTAIL.n481 VSUBS 0.014438f
C1634 VTAIL.n482 VSUBS 0.025375f
C1635 VTAIL.n483 VSUBS 0.013636f
C1636 VTAIL.n484 VSUBS 0.032229f
C1637 VTAIL.n485 VSUBS 0.014438f
C1638 VTAIL.n486 VSUBS 0.025375f
C1639 VTAIL.n487 VSUBS 0.013636f
C1640 VTAIL.n488 VSUBS 0.032229f
C1641 VTAIL.n489 VSUBS 0.014438f
C1642 VTAIL.n490 VSUBS 0.025375f
C1643 VTAIL.n491 VSUBS 0.013636f
C1644 VTAIL.n492 VSUBS 0.032229f
C1645 VTAIL.n493 VSUBS 0.014438f
C1646 VTAIL.n494 VSUBS 0.025375f
C1647 VTAIL.n495 VSUBS 0.013636f
C1648 VTAIL.n496 VSUBS 0.032229f
C1649 VTAIL.n497 VSUBS 0.014438f
C1650 VTAIL.n498 VSUBS 0.025375f
C1651 VTAIL.n499 VSUBS 0.013636f
C1652 VTAIL.n500 VSUBS 0.024172f
C1653 VTAIL.n501 VSUBS 0.020503f
C1654 VTAIL.t13 VSUBS 0.068942f
C1655 VTAIL.n502 VSUBS 0.172362f
C1656 VTAIL.n503 VSUBS 1.52003f
C1657 VTAIL.n504 VSUBS 0.013636f
C1658 VTAIL.n505 VSUBS 0.014438f
C1659 VTAIL.n506 VSUBS 0.032229f
C1660 VTAIL.n507 VSUBS 0.032229f
C1661 VTAIL.n508 VSUBS 0.014438f
C1662 VTAIL.n509 VSUBS 0.013636f
C1663 VTAIL.n510 VSUBS 0.025375f
C1664 VTAIL.n511 VSUBS 0.025375f
C1665 VTAIL.n512 VSUBS 0.013636f
C1666 VTAIL.n513 VSUBS 0.014438f
C1667 VTAIL.n514 VSUBS 0.032229f
C1668 VTAIL.n515 VSUBS 0.032229f
C1669 VTAIL.n516 VSUBS 0.014438f
C1670 VTAIL.n517 VSUBS 0.013636f
C1671 VTAIL.n518 VSUBS 0.025375f
C1672 VTAIL.n519 VSUBS 0.025375f
C1673 VTAIL.n520 VSUBS 0.013636f
C1674 VTAIL.n521 VSUBS 0.014438f
C1675 VTAIL.n522 VSUBS 0.032229f
C1676 VTAIL.n523 VSUBS 0.032229f
C1677 VTAIL.n524 VSUBS 0.014438f
C1678 VTAIL.n525 VSUBS 0.013636f
C1679 VTAIL.n526 VSUBS 0.025375f
C1680 VTAIL.n527 VSUBS 0.025375f
C1681 VTAIL.n528 VSUBS 0.013636f
C1682 VTAIL.n529 VSUBS 0.014438f
C1683 VTAIL.n530 VSUBS 0.032229f
C1684 VTAIL.n531 VSUBS 0.032229f
C1685 VTAIL.n532 VSUBS 0.014438f
C1686 VTAIL.n533 VSUBS 0.013636f
C1687 VTAIL.n534 VSUBS 0.025375f
C1688 VTAIL.n535 VSUBS 0.025375f
C1689 VTAIL.n536 VSUBS 0.013636f
C1690 VTAIL.n537 VSUBS 0.014438f
C1691 VTAIL.n538 VSUBS 0.032229f
C1692 VTAIL.n539 VSUBS 0.032229f
C1693 VTAIL.n540 VSUBS 0.014438f
C1694 VTAIL.n541 VSUBS 0.013636f
C1695 VTAIL.n542 VSUBS 0.025375f
C1696 VTAIL.n543 VSUBS 0.025375f
C1697 VTAIL.n544 VSUBS 0.013636f
C1698 VTAIL.n545 VSUBS 0.014438f
C1699 VTAIL.n546 VSUBS 0.032229f
C1700 VTAIL.n547 VSUBS 0.032229f
C1701 VTAIL.n548 VSUBS 0.076563f
C1702 VTAIL.n549 VSUBS 0.014037f
C1703 VTAIL.n550 VSUBS 0.013636f
C1704 VTAIL.n551 VSUBS 0.065933f
C1705 VTAIL.n552 VSUBS 0.03865f
C1706 VTAIL.n553 VSUBS 1.94867f
C1707 VTAIL.n554 VSUBS 0.027453f
C1708 VTAIL.n555 VSUBS 0.025375f
C1709 VTAIL.n556 VSUBS 0.014037f
C1710 VTAIL.n557 VSUBS 0.032229f
C1711 VTAIL.n558 VSUBS 0.014438f
C1712 VTAIL.n559 VSUBS 0.025375f
C1713 VTAIL.n560 VSUBS 0.013636f
C1714 VTAIL.n561 VSUBS 0.032229f
C1715 VTAIL.n562 VSUBS 0.014438f
C1716 VTAIL.n563 VSUBS 0.025375f
C1717 VTAIL.n564 VSUBS 0.013636f
C1718 VTAIL.n565 VSUBS 0.032229f
C1719 VTAIL.n566 VSUBS 0.014438f
C1720 VTAIL.n567 VSUBS 0.025375f
C1721 VTAIL.n568 VSUBS 0.013636f
C1722 VTAIL.n569 VSUBS 0.032229f
C1723 VTAIL.n570 VSUBS 0.014438f
C1724 VTAIL.n571 VSUBS 0.025375f
C1725 VTAIL.n572 VSUBS 0.013636f
C1726 VTAIL.n573 VSUBS 0.032229f
C1727 VTAIL.n574 VSUBS 0.014438f
C1728 VTAIL.n575 VSUBS 0.025375f
C1729 VTAIL.n576 VSUBS 0.013636f
C1730 VTAIL.n577 VSUBS 0.024172f
C1731 VTAIL.n578 VSUBS 0.020503f
C1732 VTAIL.t6 VSUBS 0.068942f
C1733 VTAIL.n579 VSUBS 0.172362f
C1734 VTAIL.n580 VSUBS 1.52003f
C1735 VTAIL.n581 VSUBS 0.013636f
C1736 VTAIL.n582 VSUBS 0.014438f
C1737 VTAIL.n583 VSUBS 0.032229f
C1738 VTAIL.n584 VSUBS 0.032229f
C1739 VTAIL.n585 VSUBS 0.014438f
C1740 VTAIL.n586 VSUBS 0.013636f
C1741 VTAIL.n587 VSUBS 0.025375f
C1742 VTAIL.n588 VSUBS 0.025375f
C1743 VTAIL.n589 VSUBS 0.013636f
C1744 VTAIL.n590 VSUBS 0.014438f
C1745 VTAIL.n591 VSUBS 0.032229f
C1746 VTAIL.n592 VSUBS 0.032229f
C1747 VTAIL.n593 VSUBS 0.014438f
C1748 VTAIL.n594 VSUBS 0.013636f
C1749 VTAIL.n595 VSUBS 0.025375f
C1750 VTAIL.n596 VSUBS 0.025375f
C1751 VTAIL.n597 VSUBS 0.013636f
C1752 VTAIL.n598 VSUBS 0.014438f
C1753 VTAIL.n599 VSUBS 0.032229f
C1754 VTAIL.n600 VSUBS 0.032229f
C1755 VTAIL.n601 VSUBS 0.014438f
C1756 VTAIL.n602 VSUBS 0.013636f
C1757 VTAIL.n603 VSUBS 0.025375f
C1758 VTAIL.n604 VSUBS 0.025375f
C1759 VTAIL.n605 VSUBS 0.013636f
C1760 VTAIL.n606 VSUBS 0.014438f
C1761 VTAIL.n607 VSUBS 0.032229f
C1762 VTAIL.n608 VSUBS 0.032229f
C1763 VTAIL.n609 VSUBS 0.014438f
C1764 VTAIL.n610 VSUBS 0.013636f
C1765 VTAIL.n611 VSUBS 0.025375f
C1766 VTAIL.n612 VSUBS 0.025375f
C1767 VTAIL.n613 VSUBS 0.013636f
C1768 VTAIL.n614 VSUBS 0.014438f
C1769 VTAIL.n615 VSUBS 0.032229f
C1770 VTAIL.n616 VSUBS 0.032229f
C1771 VTAIL.n617 VSUBS 0.014438f
C1772 VTAIL.n618 VSUBS 0.013636f
C1773 VTAIL.n619 VSUBS 0.025375f
C1774 VTAIL.n620 VSUBS 0.025375f
C1775 VTAIL.n621 VSUBS 0.013636f
C1776 VTAIL.n622 VSUBS 0.013636f
C1777 VTAIL.n623 VSUBS 0.014438f
C1778 VTAIL.n624 VSUBS 0.032229f
C1779 VTAIL.n625 VSUBS 0.032229f
C1780 VTAIL.n626 VSUBS 0.076563f
C1781 VTAIL.n627 VSUBS 0.014037f
C1782 VTAIL.n628 VSUBS 0.013636f
C1783 VTAIL.n629 VSUBS 0.065933f
C1784 VTAIL.n630 VSUBS 0.03865f
C1785 VTAIL.n631 VSUBS 1.94392f
C1786 VP.n0 VSUBS 0.0462f
C1787 VP.t7 VSUBS 3.60874f
C1788 VP.n1 VSUBS 0.048584f
C1789 VP.n2 VSUBS 0.024562f
C1790 VP.n3 VSUBS 0.045777f
C1791 VP.n4 VSUBS 0.024562f
C1792 VP.t6 VSUBS 3.60874f
C1793 VP.n5 VSUBS 0.045777f
C1794 VP.n6 VSUBS 0.024562f
C1795 VP.n7 VSUBS 0.045777f
C1796 VP.n8 VSUBS 0.024562f
C1797 VP.t2 VSUBS 3.60874f
C1798 VP.n9 VSUBS 0.045777f
C1799 VP.n10 VSUBS 0.024562f
C1800 VP.n11 VSUBS 0.045777f
C1801 VP.n12 VSUBS 0.0462f
C1802 VP.t3 VSUBS 3.60874f
C1803 VP.n13 VSUBS 0.048584f
C1804 VP.n14 VSUBS 0.024562f
C1805 VP.n15 VSUBS 0.045777f
C1806 VP.n16 VSUBS 0.024562f
C1807 VP.t4 VSUBS 3.60874f
C1808 VP.n17 VSUBS 0.045777f
C1809 VP.n18 VSUBS 0.024562f
C1810 VP.n19 VSUBS 0.045777f
C1811 VP.t5 VSUBS 3.99127f
C1812 VP.n20 VSUBS 1.28388f
C1813 VP.t0 VSUBS 3.60874f
C1814 VP.n21 VSUBS 1.34571f
C1815 VP.n22 VSUBS 0.037413f
C1816 VP.n23 VSUBS 0.320433f
C1817 VP.n24 VSUBS 0.024562f
C1818 VP.n25 VSUBS 0.024562f
C1819 VP.n26 VSUBS 0.045777f
C1820 VP.n27 VSUBS 0.035856f
C1821 VP.n28 VSUBS 0.035856f
C1822 VP.n29 VSUBS 0.024562f
C1823 VP.n30 VSUBS 0.024562f
C1824 VP.n31 VSUBS 0.024562f
C1825 VP.n32 VSUBS 0.045777f
C1826 VP.n33 VSUBS 0.037413f
C1827 VP.n34 VSUBS 1.25457f
C1828 VP.n35 VSUBS 0.031537f
C1829 VP.n36 VSUBS 0.024562f
C1830 VP.n37 VSUBS 0.024562f
C1831 VP.n38 VSUBS 0.024562f
C1832 VP.n39 VSUBS 0.045777f
C1833 VP.n40 VSUBS 0.044095f
C1834 VP.n41 VSUBS 0.024809f
C1835 VP.n42 VSUBS 0.024562f
C1836 VP.n43 VSUBS 0.024562f
C1837 VP.n44 VSUBS 0.024562f
C1838 VP.n45 VSUBS 0.045777f
C1839 VP.n46 VSUBS 0.04329f
C1840 VP.n47 VSUBS 1.36136f
C1841 VP.n48 VSUBS 1.75966f
C1842 VP.n49 VSUBS 1.77479f
C1843 VP.t1 VSUBS 3.60874f
C1844 VP.n50 VSUBS 1.36136f
C1845 VP.n51 VSUBS 0.04329f
C1846 VP.n52 VSUBS 0.0462f
C1847 VP.n53 VSUBS 0.024562f
C1848 VP.n54 VSUBS 0.024562f
C1849 VP.n55 VSUBS 0.048584f
C1850 VP.n56 VSUBS 0.024809f
C1851 VP.n57 VSUBS 0.044095f
C1852 VP.n58 VSUBS 0.024562f
C1853 VP.n59 VSUBS 0.024562f
C1854 VP.n60 VSUBS 0.024562f
C1855 VP.n61 VSUBS 0.045777f
C1856 VP.n62 VSUBS 0.031537f
C1857 VP.n63 VSUBS 1.25457f
C1858 VP.n64 VSUBS 0.037413f
C1859 VP.n65 VSUBS 0.024562f
C1860 VP.n66 VSUBS 0.024562f
C1861 VP.n67 VSUBS 0.024562f
C1862 VP.n68 VSUBS 0.045777f
C1863 VP.n69 VSUBS 0.035856f
C1864 VP.n70 VSUBS 0.035856f
C1865 VP.n71 VSUBS 0.024562f
C1866 VP.n72 VSUBS 0.024562f
C1867 VP.n73 VSUBS 0.024562f
C1868 VP.n74 VSUBS 0.045777f
C1869 VP.n75 VSUBS 0.037413f
C1870 VP.n76 VSUBS 1.25457f
C1871 VP.n77 VSUBS 0.031537f
C1872 VP.n78 VSUBS 0.024562f
C1873 VP.n79 VSUBS 0.024562f
C1874 VP.n80 VSUBS 0.024562f
C1875 VP.n81 VSUBS 0.045777f
C1876 VP.n82 VSUBS 0.044095f
C1877 VP.n83 VSUBS 0.024809f
C1878 VP.n84 VSUBS 0.024562f
C1879 VP.n85 VSUBS 0.024562f
C1880 VP.n86 VSUBS 0.024562f
C1881 VP.n87 VSUBS 0.045777f
C1882 VP.n88 VSUBS 0.04329f
C1883 VP.n89 VSUBS 1.36136f
C1884 VP.n90 VSUBS 0.074302f
.ends

