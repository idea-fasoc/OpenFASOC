* NGSPICE file created from diff_pair_sample_0667.ext - technology: sky130A

.subckt diff_pair_sample_0667 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t11 w_n4700_n2366# sky130_fd_pr__pfet_01v8 ad=1.15335 pd=7.32 as=2.7261 ps=14.76 w=6.99 l=3.4
X1 VDD1.t6 VP.t1 VTAIL.t12 w_n4700_n2366# sky130_fd_pr__pfet_01v8 ad=1.15335 pd=7.32 as=1.15335 ps=7.32 w=6.99 l=3.4
X2 B.t11 B.t9 B.t10 w_n4700_n2366# sky130_fd_pr__pfet_01v8 ad=2.7261 pd=14.76 as=0 ps=0 w=6.99 l=3.4
X3 VTAIL.t2 VN.t0 VDD2.t7 w_n4700_n2366# sky130_fd_pr__pfet_01v8 ad=2.7261 pd=14.76 as=1.15335 ps=7.32 w=6.99 l=3.4
X4 VDD1.t5 VP.t2 VTAIL.t10 w_n4700_n2366# sky130_fd_pr__pfet_01v8 ad=1.15335 pd=7.32 as=2.7261 ps=14.76 w=6.99 l=3.4
X5 VTAIL.t7 VN.t1 VDD2.t6 w_n4700_n2366# sky130_fd_pr__pfet_01v8 ad=2.7261 pd=14.76 as=1.15335 ps=7.32 w=6.99 l=3.4
X6 B.t8 B.t6 B.t7 w_n4700_n2366# sky130_fd_pr__pfet_01v8 ad=2.7261 pd=14.76 as=0 ps=0 w=6.99 l=3.4
X7 VTAIL.t6 VN.t2 VDD2.t5 w_n4700_n2366# sky130_fd_pr__pfet_01v8 ad=1.15335 pd=7.32 as=1.15335 ps=7.32 w=6.99 l=3.4
X8 VTAIL.t8 VP.t3 VDD1.t4 w_n4700_n2366# sky130_fd_pr__pfet_01v8 ad=2.7261 pd=14.76 as=1.15335 ps=7.32 w=6.99 l=3.4
X9 VTAIL.t5 VN.t3 VDD2.t4 w_n4700_n2366# sky130_fd_pr__pfet_01v8 ad=1.15335 pd=7.32 as=1.15335 ps=7.32 w=6.99 l=3.4
X10 VDD2.t3 VN.t4 VTAIL.t0 w_n4700_n2366# sky130_fd_pr__pfet_01v8 ad=1.15335 pd=7.32 as=2.7261 ps=14.76 w=6.99 l=3.4
X11 VTAIL.t13 VP.t4 VDD1.t3 w_n4700_n2366# sky130_fd_pr__pfet_01v8 ad=1.15335 pd=7.32 as=1.15335 ps=7.32 w=6.99 l=3.4
X12 VDD1.t2 VP.t5 VTAIL.t9 w_n4700_n2366# sky130_fd_pr__pfet_01v8 ad=1.15335 pd=7.32 as=1.15335 ps=7.32 w=6.99 l=3.4
X13 VTAIL.t14 VP.t6 VDD1.t1 w_n4700_n2366# sky130_fd_pr__pfet_01v8 ad=1.15335 pd=7.32 as=1.15335 ps=7.32 w=6.99 l=3.4
X14 VDD2.t2 VN.t5 VTAIL.t4 w_n4700_n2366# sky130_fd_pr__pfet_01v8 ad=1.15335 pd=7.32 as=1.15335 ps=7.32 w=6.99 l=3.4
X15 B.t5 B.t3 B.t4 w_n4700_n2366# sky130_fd_pr__pfet_01v8 ad=2.7261 pd=14.76 as=0 ps=0 w=6.99 l=3.4
X16 VTAIL.t15 VP.t7 VDD1.t0 w_n4700_n2366# sky130_fd_pr__pfet_01v8 ad=2.7261 pd=14.76 as=1.15335 ps=7.32 w=6.99 l=3.4
X17 VDD2.t1 VN.t6 VTAIL.t3 w_n4700_n2366# sky130_fd_pr__pfet_01v8 ad=1.15335 pd=7.32 as=1.15335 ps=7.32 w=6.99 l=3.4
X18 B.t2 B.t0 B.t1 w_n4700_n2366# sky130_fd_pr__pfet_01v8 ad=2.7261 pd=14.76 as=0 ps=0 w=6.99 l=3.4
X19 VDD2.t0 VN.t7 VTAIL.t1 w_n4700_n2366# sky130_fd_pr__pfet_01v8 ad=1.15335 pd=7.32 as=2.7261 ps=14.76 w=6.99 l=3.4
R0 VP.n24 VP.n21 161.3
R1 VP.n26 VP.n25 161.3
R2 VP.n27 VP.n20 161.3
R3 VP.n29 VP.n28 161.3
R4 VP.n30 VP.n19 161.3
R5 VP.n32 VP.n31 161.3
R6 VP.n33 VP.n18 161.3
R7 VP.n35 VP.n34 161.3
R8 VP.n37 VP.n36 161.3
R9 VP.n38 VP.n16 161.3
R10 VP.n40 VP.n39 161.3
R11 VP.n41 VP.n15 161.3
R12 VP.n43 VP.n42 161.3
R13 VP.n44 VP.n14 161.3
R14 VP.n46 VP.n45 161.3
R15 VP.n83 VP.n82 161.3
R16 VP.n81 VP.n1 161.3
R17 VP.n80 VP.n79 161.3
R18 VP.n78 VP.n2 161.3
R19 VP.n77 VP.n76 161.3
R20 VP.n75 VP.n3 161.3
R21 VP.n74 VP.n73 161.3
R22 VP.n72 VP.n71 161.3
R23 VP.n70 VP.n5 161.3
R24 VP.n69 VP.n68 161.3
R25 VP.n67 VP.n6 161.3
R26 VP.n66 VP.n65 161.3
R27 VP.n64 VP.n7 161.3
R28 VP.n63 VP.n62 161.3
R29 VP.n61 VP.n8 161.3
R30 VP.n60 VP.n59 161.3
R31 VP.n57 VP.n9 161.3
R32 VP.n56 VP.n55 161.3
R33 VP.n54 VP.n10 161.3
R34 VP.n53 VP.n52 161.3
R35 VP.n51 VP.n11 161.3
R36 VP.n50 VP.n49 161.3
R37 VP.n23 VP.t7 82.63
R38 VP.n48 VP.n12 73.1852
R39 VP.n84 VP.n0 73.1852
R40 VP.n47 VP.n13 73.1852
R41 VP.n23 VP.n22 68.9427
R42 VP.n65 VP.n6 56.5193
R43 VP.n28 VP.n19 56.5193
R44 VP.n48 VP.n47 51.0145
R45 VP.n12 VP.t3 49.5473
R46 VP.n58 VP.t1 49.5473
R47 VP.n4 VP.t6 49.5473
R48 VP.n0 VP.t0 49.5473
R49 VP.n13 VP.t2 49.5473
R50 VP.n17 VP.t4 49.5473
R51 VP.n22 VP.t5 49.5473
R52 VP.n56 VP.n10 42.4359
R53 VP.n76 VP.n2 42.4359
R54 VP.n39 VP.n15 42.4359
R55 VP.n52 VP.n10 38.5509
R56 VP.n80 VP.n2 38.5509
R57 VP.n43 VP.n15 38.5509
R58 VP.n51 VP.n50 24.4675
R59 VP.n52 VP.n51 24.4675
R60 VP.n57 VP.n56 24.4675
R61 VP.n59 VP.n57 24.4675
R62 VP.n63 VP.n8 24.4675
R63 VP.n64 VP.n63 24.4675
R64 VP.n65 VP.n64 24.4675
R65 VP.n69 VP.n6 24.4675
R66 VP.n70 VP.n69 24.4675
R67 VP.n71 VP.n70 24.4675
R68 VP.n75 VP.n74 24.4675
R69 VP.n76 VP.n75 24.4675
R70 VP.n81 VP.n80 24.4675
R71 VP.n82 VP.n81 24.4675
R72 VP.n44 VP.n43 24.4675
R73 VP.n45 VP.n44 24.4675
R74 VP.n32 VP.n19 24.4675
R75 VP.n33 VP.n32 24.4675
R76 VP.n34 VP.n33 24.4675
R77 VP.n38 VP.n37 24.4675
R78 VP.n39 VP.n38 24.4675
R79 VP.n26 VP.n21 24.4675
R80 VP.n27 VP.n26 24.4675
R81 VP.n28 VP.n27 24.4675
R82 VP.n59 VP.n58 18.8401
R83 VP.n74 VP.n4 18.8401
R84 VP.n37 VP.n17 18.8401
R85 VP.n50 VP.n12 16.8827
R86 VP.n82 VP.n0 16.8827
R87 VP.n45 VP.n13 16.8827
R88 VP.n58 VP.n8 5.62791
R89 VP.n71 VP.n4 5.62791
R90 VP.n34 VP.n17 5.62791
R91 VP.n22 VP.n21 5.62791
R92 VP.n24 VP.n23 4.05577
R93 VP.n47 VP.n46 0.354971
R94 VP.n49 VP.n48 0.354971
R95 VP.n84 VP.n83 0.354971
R96 VP VP.n84 0.26696
R97 VP.n25 VP.n24 0.189894
R98 VP.n25 VP.n20 0.189894
R99 VP.n29 VP.n20 0.189894
R100 VP.n30 VP.n29 0.189894
R101 VP.n31 VP.n30 0.189894
R102 VP.n31 VP.n18 0.189894
R103 VP.n35 VP.n18 0.189894
R104 VP.n36 VP.n35 0.189894
R105 VP.n36 VP.n16 0.189894
R106 VP.n40 VP.n16 0.189894
R107 VP.n41 VP.n40 0.189894
R108 VP.n42 VP.n41 0.189894
R109 VP.n42 VP.n14 0.189894
R110 VP.n46 VP.n14 0.189894
R111 VP.n49 VP.n11 0.189894
R112 VP.n53 VP.n11 0.189894
R113 VP.n54 VP.n53 0.189894
R114 VP.n55 VP.n54 0.189894
R115 VP.n55 VP.n9 0.189894
R116 VP.n60 VP.n9 0.189894
R117 VP.n61 VP.n60 0.189894
R118 VP.n62 VP.n61 0.189894
R119 VP.n62 VP.n7 0.189894
R120 VP.n66 VP.n7 0.189894
R121 VP.n67 VP.n66 0.189894
R122 VP.n68 VP.n67 0.189894
R123 VP.n68 VP.n5 0.189894
R124 VP.n72 VP.n5 0.189894
R125 VP.n73 VP.n72 0.189894
R126 VP.n73 VP.n3 0.189894
R127 VP.n77 VP.n3 0.189894
R128 VP.n78 VP.n77 0.189894
R129 VP.n79 VP.n78 0.189894
R130 VP.n79 VP.n1 0.189894
R131 VP.n83 VP.n1 0.189894
R132 VTAIL.n11 VTAIL.t15 72.9921
R133 VTAIL.n10 VTAIL.t0 72.9921
R134 VTAIL.n7 VTAIL.t7 72.9921
R135 VTAIL.n15 VTAIL.t1 72.9919
R136 VTAIL.n2 VTAIL.t2 72.9919
R137 VTAIL.n3 VTAIL.t11 72.9919
R138 VTAIL.n6 VTAIL.t8 72.9919
R139 VTAIL.n14 VTAIL.t10 72.9919
R140 VTAIL.n13 VTAIL.n12 68.3419
R141 VTAIL.n9 VTAIL.n8 68.3419
R142 VTAIL.n1 VTAIL.n0 68.3418
R143 VTAIL.n5 VTAIL.n4 68.3418
R144 VTAIL.n15 VTAIL.n14 21.6083
R145 VTAIL.n7 VTAIL.n6 21.6083
R146 VTAIL.n0 VTAIL.t3 4.65071
R147 VTAIL.n0 VTAIL.t6 4.65071
R148 VTAIL.n4 VTAIL.t12 4.65071
R149 VTAIL.n4 VTAIL.t14 4.65071
R150 VTAIL.n12 VTAIL.t9 4.65071
R151 VTAIL.n12 VTAIL.t13 4.65071
R152 VTAIL.n8 VTAIL.t4 4.65071
R153 VTAIL.n8 VTAIL.t5 4.65071
R154 VTAIL.n9 VTAIL.n7 3.21602
R155 VTAIL.n10 VTAIL.n9 3.21602
R156 VTAIL.n13 VTAIL.n11 3.21602
R157 VTAIL.n14 VTAIL.n13 3.21602
R158 VTAIL.n6 VTAIL.n5 3.21602
R159 VTAIL.n5 VTAIL.n3 3.21602
R160 VTAIL.n2 VTAIL.n1 3.21602
R161 VTAIL VTAIL.n15 3.15783
R162 VTAIL.n11 VTAIL.n10 0.470328
R163 VTAIL.n3 VTAIL.n2 0.470328
R164 VTAIL VTAIL.n1 0.0586897
R165 VDD1 VDD1.n0 86.6866
R166 VDD1.n3 VDD1.n2 86.573
R167 VDD1.n3 VDD1.n1 86.573
R168 VDD1.n5 VDD1.n4 85.0205
R169 VDD1.n5 VDD1.n3 44.794
R170 VDD1.n4 VDD1.t3 4.65071
R171 VDD1.n4 VDD1.t5 4.65071
R172 VDD1.n0 VDD1.t0 4.65071
R173 VDD1.n0 VDD1.t2 4.65071
R174 VDD1.n2 VDD1.t1 4.65071
R175 VDD1.n2 VDD1.t7 4.65071
R176 VDD1.n1 VDD1.t4 4.65071
R177 VDD1.n1 VDD1.t6 4.65071
R178 VDD1 VDD1.n5 1.55007
R179 B.n580 B.n579 585
R180 B.n581 B.n68 585
R181 B.n583 B.n582 585
R182 B.n584 B.n67 585
R183 B.n586 B.n585 585
R184 B.n587 B.n66 585
R185 B.n589 B.n588 585
R186 B.n590 B.n65 585
R187 B.n592 B.n591 585
R188 B.n593 B.n64 585
R189 B.n595 B.n594 585
R190 B.n596 B.n63 585
R191 B.n598 B.n597 585
R192 B.n599 B.n62 585
R193 B.n601 B.n600 585
R194 B.n602 B.n61 585
R195 B.n604 B.n603 585
R196 B.n605 B.n60 585
R197 B.n607 B.n606 585
R198 B.n608 B.n59 585
R199 B.n610 B.n609 585
R200 B.n611 B.n58 585
R201 B.n613 B.n612 585
R202 B.n614 B.n57 585
R203 B.n616 B.n615 585
R204 B.n617 B.n56 585
R205 B.n619 B.n618 585
R206 B.n621 B.n53 585
R207 B.n623 B.n622 585
R208 B.n624 B.n52 585
R209 B.n626 B.n625 585
R210 B.n627 B.n51 585
R211 B.n629 B.n628 585
R212 B.n630 B.n50 585
R213 B.n632 B.n631 585
R214 B.n633 B.n47 585
R215 B.n636 B.n635 585
R216 B.n637 B.n46 585
R217 B.n639 B.n638 585
R218 B.n640 B.n45 585
R219 B.n642 B.n641 585
R220 B.n643 B.n44 585
R221 B.n645 B.n644 585
R222 B.n646 B.n43 585
R223 B.n648 B.n647 585
R224 B.n649 B.n42 585
R225 B.n651 B.n650 585
R226 B.n652 B.n41 585
R227 B.n654 B.n653 585
R228 B.n655 B.n40 585
R229 B.n657 B.n656 585
R230 B.n658 B.n39 585
R231 B.n660 B.n659 585
R232 B.n661 B.n38 585
R233 B.n663 B.n662 585
R234 B.n664 B.n37 585
R235 B.n666 B.n665 585
R236 B.n667 B.n36 585
R237 B.n669 B.n668 585
R238 B.n670 B.n35 585
R239 B.n672 B.n671 585
R240 B.n673 B.n34 585
R241 B.n675 B.n674 585
R242 B.n578 B.n69 585
R243 B.n577 B.n576 585
R244 B.n575 B.n70 585
R245 B.n574 B.n573 585
R246 B.n572 B.n71 585
R247 B.n571 B.n570 585
R248 B.n569 B.n72 585
R249 B.n568 B.n567 585
R250 B.n566 B.n73 585
R251 B.n565 B.n564 585
R252 B.n563 B.n74 585
R253 B.n562 B.n561 585
R254 B.n560 B.n75 585
R255 B.n559 B.n558 585
R256 B.n557 B.n76 585
R257 B.n556 B.n555 585
R258 B.n554 B.n77 585
R259 B.n553 B.n552 585
R260 B.n551 B.n78 585
R261 B.n550 B.n549 585
R262 B.n548 B.n79 585
R263 B.n547 B.n546 585
R264 B.n545 B.n80 585
R265 B.n544 B.n543 585
R266 B.n542 B.n81 585
R267 B.n541 B.n540 585
R268 B.n539 B.n82 585
R269 B.n538 B.n537 585
R270 B.n536 B.n83 585
R271 B.n535 B.n534 585
R272 B.n533 B.n84 585
R273 B.n532 B.n531 585
R274 B.n530 B.n85 585
R275 B.n529 B.n528 585
R276 B.n527 B.n86 585
R277 B.n526 B.n525 585
R278 B.n524 B.n87 585
R279 B.n523 B.n522 585
R280 B.n521 B.n88 585
R281 B.n520 B.n519 585
R282 B.n518 B.n89 585
R283 B.n517 B.n516 585
R284 B.n515 B.n90 585
R285 B.n514 B.n513 585
R286 B.n512 B.n91 585
R287 B.n511 B.n510 585
R288 B.n509 B.n92 585
R289 B.n508 B.n507 585
R290 B.n506 B.n93 585
R291 B.n505 B.n504 585
R292 B.n503 B.n94 585
R293 B.n502 B.n501 585
R294 B.n500 B.n95 585
R295 B.n499 B.n498 585
R296 B.n497 B.n96 585
R297 B.n496 B.n495 585
R298 B.n494 B.n97 585
R299 B.n493 B.n492 585
R300 B.n491 B.n98 585
R301 B.n490 B.n489 585
R302 B.n488 B.n99 585
R303 B.n487 B.n486 585
R304 B.n485 B.n100 585
R305 B.n484 B.n483 585
R306 B.n482 B.n101 585
R307 B.n481 B.n480 585
R308 B.n479 B.n102 585
R309 B.n478 B.n477 585
R310 B.n476 B.n103 585
R311 B.n475 B.n474 585
R312 B.n473 B.n104 585
R313 B.n472 B.n471 585
R314 B.n470 B.n105 585
R315 B.n469 B.n468 585
R316 B.n467 B.n106 585
R317 B.n466 B.n465 585
R318 B.n464 B.n107 585
R319 B.n463 B.n462 585
R320 B.n461 B.n108 585
R321 B.n460 B.n459 585
R322 B.n458 B.n109 585
R323 B.n457 B.n456 585
R324 B.n455 B.n110 585
R325 B.n454 B.n453 585
R326 B.n452 B.n111 585
R327 B.n451 B.n450 585
R328 B.n449 B.n112 585
R329 B.n448 B.n447 585
R330 B.n446 B.n113 585
R331 B.n445 B.n444 585
R332 B.n443 B.n114 585
R333 B.n442 B.n441 585
R334 B.n440 B.n115 585
R335 B.n439 B.n438 585
R336 B.n437 B.n116 585
R337 B.n436 B.n435 585
R338 B.n434 B.n117 585
R339 B.n433 B.n432 585
R340 B.n431 B.n118 585
R341 B.n430 B.n429 585
R342 B.n428 B.n119 585
R343 B.n427 B.n426 585
R344 B.n425 B.n120 585
R345 B.n424 B.n423 585
R346 B.n422 B.n121 585
R347 B.n421 B.n420 585
R348 B.n419 B.n122 585
R349 B.n418 B.n417 585
R350 B.n416 B.n123 585
R351 B.n415 B.n414 585
R352 B.n413 B.n124 585
R353 B.n412 B.n411 585
R354 B.n410 B.n125 585
R355 B.n409 B.n408 585
R356 B.n407 B.n126 585
R357 B.n406 B.n405 585
R358 B.n404 B.n127 585
R359 B.n403 B.n402 585
R360 B.n401 B.n128 585
R361 B.n400 B.n399 585
R362 B.n398 B.n129 585
R363 B.n397 B.n396 585
R364 B.n395 B.n130 585
R365 B.n394 B.n393 585
R366 B.n392 B.n131 585
R367 B.n391 B.n390 585
R368 B.n389 B.n132 585
R369 B.n293 B.n168 585
R370 B.n295 B.n294 585
R371 B.n296 B.n167 585
R372 B.n298 B.n297 585
R373 B.n299 B.n166 585
R374 B.n301 B.n300 585
R375 B.n302 B.n165 585
R376 B.n304 B.n303 585
R377 B.n305 B.n164 585
R378 B.n307 B.n306 585
R379 B.n308 B.n163 585
R380 B.n310 B.n309 585
R381 B.n311 B.n162 585
R382 B.n313 B.n312 585
R383 B.n314 B.n161 585
R384 B.n316 B.n315 585
R385 B.n317 B.n160 585
R386 B.n319 B.n318 585
R387 B.n320 B.n159 585
R388 B.n322 B.n321 585
R389 B.n323 B.n158 585
R390 B.n325 B.n324 585
R391 B.n326 B.n157 585
R392 B.n328 B.n327 585
R393 B.n329 B.n156 585
R394 B.n331 B.n330 585
R395 B.n332 B.n153 585
R396 B.n335 B.n334 585
R397 B.n336 B.n152 585
R398 B.n338 B.n337 585
R399 B.n339 B.n151 585
R400 B.n341 B.n340 585
R401 B.n342 B.n150 585
R402 B.n344 B.n343 585
R403 B.n345 B.n149 585
R404 B.n347 B.n346 585
R405 B.n349 B.n348 585
R406 B.n350 B.n145 585
R407 B.n352 B.n351 585
R408 B.n353 B.n144 585
R409 B.n355 B.n354 585
R410 B.n356 B.n143 585
R411 B.n358 B.n357 585
R412 B.n359 B.n142 585
R413 B.n361 B.n360 585
R414 B.n362 B.n141 585
R415 B.n364 B.n363 585
R416 B.n365 B.n140 585
R417 B.n367 B.n366 585
R418 B.n368 B.n139 585
R419 B.n370 B.n369 585
R420 B.n371 B.n138 585
R421 B.n373 B.n372 585
R422 B.n374 B.n137 585
R423 B.n376 B.n375 585
R424 B.n377 B.n136 585
R425 B.n379 B.n378 585
R426 B.n380 B.n135 585
R427 B.n382 B.n381 585
R428 B.n383 B.n134 585
R429 B.n385 B.n384 585
R430 B.n386 B.n133 585
R431 B.n388 B.n387 585
R432 B.n292 B.n291 585
R433 B.n290 B.n169 585
R434 B.n289 B.n288 585
R435 B.n287 B.n170 585
R436 B.n286 B.n285 585
R437 B.n284 B.n171 585
R438 B.n283 B.n282 585
R439 B.n281 B.n172 585
R440 B.n280 B.n279 585
R441 B.n278 B.n173 585
R442 B.n277 B.n276 585
R443 B.n275 B.n174 585
R444 B.n274 B.n273 585
R445 B.n272 B.n175 585
R446 B.n271 B.n270 585
R447 B.n269 B.n176 585
R448 B.n268 B.n267 585
R449 B.n266 B.n177 585
R450 B.n265 B.n264 585
R451 B.n263 B.n178 585
R452 B.n262 B.n261 585
R453 B.n260 B.n179 585
R454 B.n259 B.n258 585
R455 B.n257 B.n180 585
R456 B.n256 B.n255 585
R457 B.n254 B.n181 585
R458 B.n253 B.n252 585
R459 B.n251 B.n182 585
R460 B.n250 B.n249 585
R461 B.n248 B.n183 585
R462 B.n247 B.n246 585
R463 B.n245 B.n184 585
R464 B.n244 B.n243 585
R465 B.n242 B.n185 585
R466 B.n241 B.n240 585
R467 B.n239 B.n186 585
R468 B.n238 B.n237 585
R469 B.n236 B.n187 585
R470 B.n235 B.n234 585
R471 B.n233 B.n188 585
R472 B.n232 B.n231 585
R473 B.n230 B.n189 585
R474 B.n229 B.n228 585
R475 B.n227 B.n190 585
R476 B.n226 B.n225 585
R477 B.n224 B.n191 585
R478 B.n223 B.n222 585
R479 B.n221 B.n192 585
R480 B.n220 B.n219 585
R481 B.n218 B.n193 585
R482 B.n217 B.n216 585
R483 B.n215 B.n194 585
R484 B.n214 B.n213 585
R485 B.n212 B.n195 585
R486 B.n211 B.n210 585
R487 B.n209 B.n196 585
R488 B.n208 B.n207 585
R489 B.n206 B.n197 585
R490 B.n205 B.n204 585
R491 B.n203 B.n198 585
R492 B.n202 B.n201 585
R493 B.n200 B.n199 585
R494 B.n2 B.n0 585
R495 B.n769 B.n1 585
R496 B.n768 B.n767 585
R497 B.n766 B.n3 585
R498 B.n765 B.n764 585
R499 B.n763 B.n4 585
R500 B.n762 B.n761 585
R501 B.n760 B.n5 585
R502 B.n759 B.n758 585
R503 B.n757 B.n6 585
R504 B.n756 B.n755 585
R505 B.n754 B.n7 585
R506 B.n753 B.n752 585
R507 B.n751 B.n8 585
R508 B.n750 B.n749 585
R509 B.n748 B.n9 585
R510 B.n747 B.n746 585
R511 B.n745 B.n10 585
R512 B.n744 B.n743 585
R513 B.n742 B.n11 585
R514 B.n741 B.n740 585
R515 B.n739 B.n12 585
R516 B.n738 B.n737 585
R517 B.n736 B.n13 585
R518 B.n735 B.n734 585
R519 B.n733 B.n14 585
R520 B.n732 B.n731 585
R521 B.n730 B.n15 585
R522 B.n729 B.n728 585
R523 B.n727 B.n16 585
R524 B.n726 B.n725 585
R525 B.n724 B.n17 585
R526 B.n723 B.n722 585
R527 B.n721 B.n18 585
R528 B.n720 B.n719 585
R529 B.n718 B.n19 585
R530 B.n717 B.n716 585
R531 B.n715 B.n20 585
R532 B.n714 B.n713 585
R533 B.n712 B.n21 585
R534 B.n711 B.n710 585
R535 B.n709 B.n22 585
R536 B.n708 B.n707 585
R537 B.n706 B.n23 585
R538 B.n705 B.n704 585
R539 B.n703 B.n24 585
R540 B.n702 B.n701 585
R541 B.n700 B.n25 585
R542 B.n699 B.n698 585
R543 B.n697 B.n26 585
R544 B.n696 B.n695 585
R545 B.n694 B.n27 585
R546 B.n693 B.n692 585
R547 B.n691 B.n28 585
R548 B.n690 B.n689 585
R549 B.n688 B.n29 585
R550 B.n687 B.n686 585
R551 B.n685 B.n30 585
R552 B.n684 B.n683 585
R553 B.n682 B.n31 585
R554 B.n681 B.n680 585
R555 B.n679 B.n32 585
R556 B.n678 B.n677 585
R557 B.n676 B.n33 585
R558 B.n771 B.n770 585
R559 B.n293 B.n292 521.33
R560 B.n674 B.n33 521.33
R561 B.n389 B.n388 521.33
R562 B.n580 B.n69 521.33
R563 B.n146 B.t9 258.548
R564 B.n154 B.t0 258.548
R565 B.n48 B.t3 258.548
R566 B.n54 B.t6 258.548
R567 B.n146 B.t11 185.648
R568 B.n54 B.t7 185.648
R569 B.n154 B.t2 185.641
R570 B.n48 B.t4 185.641
R571 B.n292 B.n169 163.367
R572 B.n288 B.n169 163.367
R573 B.n288 B.n287 163.367
R574 B.n287 B.n286 163.367
R575 B.n286 B.n171 163.367
R576 B.n282 B.n171 163.367
R577 B.n282 B.n281 163.367
R578 B.n281 B.n280 163.367
R579 B.n280 B.n173 163.367
R580 B.n276 B.n173 163.367
R581 B.n276 B.n275 163.367
R582 B.n275 B.n274 163.367
R583 B.n274 B.n175 163.367
R584 B.n270 B.n175 163.367
R585 B.n270 B.n269 163.367
R586 B.n269 B.n268 163.367
R587 B.n268 B.n177 163.367
R588 B.n264 B.n177 163.367
R589 B.n264 B.n263 163.367
R590 B.n263 B.n262 163.367
R591 B.n262 B.n179 163.367
R592 B.n258 B.n179 163.367
R593 B.n258 B.n257 163.367
R594 B.n257 B.n256 163.367
R595 B.n256 B.n181 163.367
R596 B.n252 B.n181 163.367
R597 B.n252 B.n251 163.367
R598 B.n251 B.n250 163.367
R599 B.n250 B.n183 163.367
R600 B.n246 B.n183 163.367
R601 B.n246 B.n245 163.367
R602 B.n245 B.n244 163.367
R603 B.n244 B.n185 163.367
R604 B.n240 B.n185 163.367
R605 B.n240 B.n239 163.367
R606 B.n239 B.n238 163.367
R607 B.n238 B.n187 163.367
R608 B.n234 B.n187 163.367
R609 B.n234 B.n233 163.367
R610 B.n233 B.n232 163.367
R611 B.n232 B.n189 163.367
R612 B.n228 B.n189 163.367
R613 B.n228 B.n227 163.367
R614 B.n227 B.n226 163.367
R615 B.n226 B.n191 163.367
R616 B.n222 B.n191 163.367
R617 B.n222 B.n221 163.367
R618 B.n221 B.n220 163.367
R619 B.n220 B.n193 163.367
R620 B.n216 B.n193 163.367
R621 B.n216 B.n215 163.367
R622 B.n215 B.n214 163.367
R623 B.n214 B.n195 163.367
R624 B.n210 B.n195 163.367
R625 B.n210 B.n209 163.367
R626 B.n209 B.n208 163.367
R627 B.n208 B.n197 163.367
R628 B.n204 B.n197 163.367
R629 B.n204 B.n203 163.367
R630 B.n203 B.n202 163.367
R631 B.n202 B.n199 163.367
R632 B.n199 B.n2 163.367
R633 B.n770 B.n2 163.367
R634 B.n770 B.n769 163.367
R635 B.n769 B.n768 163.367
R636 B.n768 B.n3 163.367
R637 B.n764 B.n3 163.367
R638 B.n764 B.n763 163.367
R639 B.n763 B.n762 163.367
R640 B.n762 B.n5 163.367
R641 B.n758 B.n5 163.367
R642 B.n758 B.n757 163.367
R643 B.n757 B.n756 163.367
R644 B.n756 B.n7 163.367
R645 B.n752 B.n7 163.367
R646 B.n752 B.n751 163.367
R647 B.n751 B.n750 163.367
R648 B.n750 B.n9 163.367
R649 B.n746 B.n9 163.367
R650 B.n746 B.n745 163.367
R651 B.n745 B.n744 163.367
R652 B.n744 B.n11 163.367
R653 B.n740 B.n11 163.367
R654 B.n740 B.n739 163.367
R655 B.n739 B.n738 163.367
R656 B.n738 B.n13 163.367
R657 B.n734 B.n13 163.367
R658 B.n734 B.n733 163.367
R659 B.n733 B.n732 163.367
R660 B.n732 B.n15 163.367
R661 B.n728 B.n15 163.367
R662 B.n728 B.n727 163.367
R663 B.n727 B.n726 163.367
R664 B.n726 B.n17 163.367
R665 B.n722 B.n17 163.367
R666 B.n722 B.n721 163.367
R667 B.n721 B.n720 163.367
R668 B.n720 B.n19 163.367
R669 B.n716 B.n19 163.367
R670 B.n716 B.n715 163.367
R671 B.n715 B.n714 163.367
R672 B.n714 B.n21 163.367
R673 B.n710 B.n21 163.367
R674 B.n710 B.n709 163.367
R675 B.n709 B.n708 163.367
R676 B.n708 B.n23 163.367
R677 B.n704 B.n23 163.367
R678 B.n704 B.n703 163.367
R679 B.n703 B.n702 163.367
R680 B.n702 B.n25 163.367
R681 B.n698 B.n25 163.367
R682 B.n698 B.n697 163.367
R683 B.n697 B.n696 163.367
R684 B.n696 B.n27 163.367
R685 B.n692 B.n27 163.367
R686 B.n692 B.n691 163.367
R687 B.n691 B.n690 163.367
R688 B.n690 B.n29 163.367
R689 B.n686 B.n29 163.367
R690 B.n686 B.n685 163.367
R691 B.n685 B.n684 163.367
R692 B.n684 B.n31 163.367
R693 B.n680 B.n31 163.367
R694 B.n680 B.n679 163.367
R695 B.n679 B.n678 163.367
R696 B.n678 B.n33 163.367
R697 B.n294 B.n293 163.367
R698 B.n294 B.n167 163.367
R699 B.n298 B.n167 163.367
R700 B.n299 B.n298 163.367
R701 B.n300 B.n299 163.367
R702 B.n300 B.n165 163.367
R703 B.n304 B.n165 163.367
R704 B.n305 B.n304 163.367
R705 B.n306 B.n305 163.367
R706 B.n306 B.n163 163.367
R707 B.n310 B.n163 163.367
R708 B.n311 B.n310 163.367
R709 B.n312 B.n311 163.367
R710 B.n312 B.n161 163.367
R711 B.n316 B.n161 163.367
R712 B.n317 B.n316 163.367
R713 B.n318 B.n317 163.367
R714 B.n318 B.n159 163.367
R715 B.n322 B.n159 163.367
R716 B.n323 B.n322 163.367
R717 B.n324 B.n323 163.367
R718 B.n324 B.n157 163.367
R719 B.n328 B.n157 163.367
R720 B.n329 B.n328 163.367
R721 B.n330 B.n329 163.367
R722 B.n330 B.n153 163.367
R723 B.n335 B.n153 163.367
R724 B.n336 B.n335 163.367
R725 B.n337 B.n336 163.367
R726 B.n337 B.n151 163.367
R727 B.n341 B.n151 163.367
R728 B.n342 B.n341 163.367
R729 B.n343 B.n342 163.367
R730 B.n343 B.n149 163.367
R731 B.n347 B.n149 163.367
R732 B.n348 B.n347 163.367
R733 B.n348 B.n145 163.367
R734 B.n352 B.n145 163.367
R735 B.n353 B.n352 163.367
R736 B.n354 B.n353 163.367
R737 B.n354 B.n143 163.367
R738 B.n358 B.n143 163.367
R739 B.n359 B.n358 163.367
R740 B.n360 B.n359 163.367
R741 B.n360 B.n141 163.367
R742 B.n364 B.n141 163.367
R743 B.n365 B.n364 163.367
R744 B.n366 B.n365 163.367
R745 B.n366 B.n139 163.367
R746 B.n370 B.n139 163.367
R747 B.n371 B.n370 163.367
R748 B.n372 B.n371 163.367
R749 B.n372 B.n137 163.367
R750 B.n376 B.n137 163.367
R751 B.n377 B.n376 163.367
R752 B.n378 B.n377 163.367
R753 B.n378 B.n135 163.367
R754 B.n382 B.n135 163.367
R755 B.n383 B.n382 163.367
R756 B.n384 B.n383 163.367
R757 B.n384 B.n133 163.367
R758 B.n388 B.n133 163.367
R759 B.n390 B.n389 163.367
R760 B.n390 B.n131 163.367
R761 B.n394 B.n131 163.367
R762 B.n395 B.n394 163.367
R763 B.n396 B.n395 163.367
R764 B.n396 B.n129 163.367
R765 B.n400 B.n129 163.367
R766 B.n401 B.n400 163.367
R767 B.n402 B.n401 163.367
R768 B.n402 B.n127 163.367
R769 B.n406 B.n127 163.367
R770 B.n407 B.n406 163.367
R771 B.n408 B.n407 163.367
R772 B.n408 B.n125 163.367
R773 B.n412 B.n125 163.367
R774 B.n413 B.n412 163.367
R775 B.n414 B.n413 163.367
R776 B.n414 B.n123 163.367
R777 B.n418 B.n123 163.367
R778 B.n419 B.n418 163.367
R779 B.n420 B.n419 163.367
R780 B.n420 B.n121 163.367
R781 B.n424 B.n121 163.367
R782 B.n425 B.n424 163.367
R783 B.n426 B.n425 163.367
R784 B.n426 B.n119 163.367
R785 B.n430 B.n119 163.367
R786 B.n431 B.n430 163.367
R787 B.n432 B.n431 163.367
R788 B.n432 B.n117 163.367
R789 B.n436 B.n117 163.367
R790 B.n437 B.n436 163.367
R791 B.n438 B.n437 163.367
R792 B.n438 B.n115 163.367
R793 B.n442 B.n115 163.367
R794 B.n443 B.n442 163.367
R795 B.n444 B.n443 163.367
R796 B.n444 B.n113 163.367
R797 B.n448 B.n113 163.367
R798 B.n449 B.n448 163.367
R799 B.n450 B.n449 163.367
R800 B.n450 B.n111 163.367
R801 B.n454 B.n111 163.367
R802 B.n455 B.n454 163.367
R803 B.n456 B.n455 163.367
R804 B.n456 B.n109 163.367
R805 B.n460 B.n109 163.367
R806 B.n461 B.n460 163.367
R807 B.n462 B.n461 163.367
R808 B.n462 B.n107 163.367
R809 B.n466 B.n107 163.367
R810 B.n467 B.n466 163.367
R811 B.n468 B.n467 163.367
R812 B.n468 B.n105 163.367
R813 B.n472 B.n105 163.367
R814 B.n473 B.n472 163.367
R815 B.n474 B.n473 163.367
R816 B.n474 B.n103 163.367
R817 B.n478 B.n103 163.367
R818 B.n479 B.n478 163.367
R819 B.n480 B.n479 163.367
R820 B.n480 B.n101 163.367
R821 B.n484 B.n101 163.367
R822 B.n485 B.n484 163.367
R823 B.n486 B.n485 163.367
R824 B.n486 B.n99 163.367
R825 B.n490 B.n99 163.367
R826 B.n491 B.n490 163.367
R827 B.n492 B.n491 163.367
R828 B.n492 B.n97 163.367
R829 B.n496 B.n97 163.367
R830 B.n497 B.n496 163.367
R831 B.n498 B.n497 163.367
R832 B.n498 B.n95 163.367
R833 B.n502 B.n95 163.367
R834 B.n503 B.n502 163.367
R835 B.n504 B.n503 163.367
R836 B.n504 B.n93 163.367
R837 B.n508 B.n93 163.367
R838 B.n509 B.n508 163.367
R839 B.n510 B.n509 163.367
R840 B.n510 B.n91 163.367
R841 B.n514 B.n91 163.367
R842 B.n515 B.n514 163.367
R843 B.n516 B.n515 163.367
R844 B.n516 B.n89 163.367
R845 B.n520 B.n89 163.367
R846 B.n521 B.n520 163.367
R847 B.n522 B.n521 163.367
R848 B.n522 B.n87 163.367
R849 B.n526 B.n87 163.367
R850 B.n527 B.n526 163.367
R851 B.n528 B.n527 163.367
R852 B.n528 B.n85 163.367
R853 B.n532 B.n85 163.367
R854 B.n533 B.n532 163.367
R855 B.n534 B.n533 163.367
R856 B.n534 B.n83 163.367
R857 B.n538 B.n83 163.367
R858 B.n539 B.n538 163.367
R859 B.n540 B.n539 163.367
R860 B.n540 B.n81 163.367
R861 B.n544 B.n81 163.367
R862 B.n545 B.n544 163.367
R863 B.n546 B.n545 163.367
R864 B.n546 B.n79 163.367
R865 B.n550 B.n79 163.367
R866 B.n551 B.n550 163.367
R867 B.n552 B.n551 163.367
R868 B.n552 B.n77 163.367
R869 B.n556 B.n77 163.367
R870 B.n557 B.n556 163.367
R871 B.n558 B.n557 163.367
R872 B.n558 B.n75 163.367
R873 B.n562 B.n75 163.367
R874 B.n563 B.n562 163.367
R875 B.n564 B.n563 163.367
R876 B.n564 B.n73 163.367
R877 B.n568 B.n73 163.367
R878 B.n569 B.n568 163.367
R879 B.n570 B.n569 163.367
R880 B.n570 B.n71 163.367
R881 B.n574 B.n71 163.367
R882 B.n575 B.n574 163.367
R883 B.n576 B.n575 163.367
R884 B.n576 B.n69 163.367
R885 B.n674 B.n673 163.367
R886 B.n673 B.n672 163.367
R887 B.n672 B.n35 163.367
R888 B.n668 B.n35 163.367
R889 B.n668 B.n667 163.367
R890 B.n667 B.n666 163.367
R891 B.n666 B.n37 163.367
R892 B.n662 B.n37 163.367
R893 B.n662 B.n661 163.367
R894 B.n661 B.n660 163.367
R895 B.n660 B.n39 163.367
R896 B.n656 B.n39 163.367
R897 B.n656 B.n655 163.367
R898 B.n655 B.n654 163.367
R899 B.n654 B.n41 163.367
R900 B.n650 B.n41 163.367
R901 B.n650 B.n649 163.367
R902 B.n649 B.n648 163.367
R903 B.n648 B.n43 163.367
R904 B.n644 B.n43 163.367
R905 B.n644 B.n643 163.367
R906 B.n643 B.n642 163.367
R907 B.n642 B.n45 163.367
R908 B.n638 B.n45 163.367
R909 B.n638 B.n637 163.367
R910 B.n637 B.n636 163.367
R911 B.n636 B.n47 163.367
R912 B.n631 B.n47 163.367
R913 B.n631 B.n630 163.367
R914 B.n630 B.n629 163.367
R915 B.n629 B.n51 163.367
R916 B.n625 B.n51 163.367
R917 B.n625 B.n624 163.367
R918 B.n624 B.n623 163.367
R919 B.n623 B.n53 163.367
R920 B.n618 B.n53 163.367
R921 B.n618 B.n617 163.367
R922 B.n617 B.n616 163.367
R923 B.n616 B.n57 163.367
R924 B.n612 B.n57 163.367
R925 B.n612 B.n611 163.367
R926 B.n611 B.n610 163.367
R927 B.n610 B.n59 163.367
R928 B.n606 B.n59 163.367
R929 B.n606 B.n605 163.367
R930 B.n605 B.n604 163.367
R931 B.n604 B.n61 163.367
R932 B.n600 B.n61 163.367
R933 B.n600 B.n599 163.367
R934 B.n599 B.n598 163.367
R935 B.n598 B.n63 163.367
R936 B.n594 B.n63 163.367
R937 B.n594 B.n593 163.367
R938 B.n593 B.n592 163.367
R939 B.n592 B.n65 163.367
R940 B.n588 B.n65 163.367
R941 B.n588 B.n587 163.367
R942 B.n587 B.n586 163.367
R943 B.n586 B.n67 163.367
R944 B.n582 B.n67 163.367
R945 B.n582 B.n581 163.367
R946 B.n581 B.n580 163.367
R947 B.n147 B.t10 113.308
R948 B.n55 B.t8 113.308
R949 B.n155 B.t1 113.302
R950 B.n49 B.t5 113.302
R951 B.n147 B.n146 72.3399
R952 B.n155 B.n154 72.3399
R953 B.n49 B.n48 72.3399
R954 B.n55 B.n54 72.3399
R955 B.n148 B.n147 59.5399
R956 B.n333 B.n155 59.5399
R957 B.n634 B.n49 59.5399
R958 B.n620 B.n55 59.5399
R959 B.n676 B.n675 33.8737
R960 B.n579 B.n578 33.8737
R961 B.n387 B.n132 33.8737
R962 B.n291 B.n168 33.8737
R963 B B.n771 18.0485
R964 B.n675 B.n34 10.6151
R965 B.n671 B.n34 10.6151
R966 B.n671 B.n670 10.6151
R967 B.n670 B.n669 10.6151
R968 B.n669 B.n36 10.6151
R969 B.n665 B.n36 10.6151
R970 B.n665 B.n664 10.6151
R971 B.n664 B.n663 10.6151
R972 B.n663 B.n38 10.6151
R973 B.n659 B.n38 10.6151
R974 B.n659 B.n658 10.6151
R975 B.n658 B.n657 10.6151
R976 B.n657 B.n40 10.6151
R977 B.n653 B.n40 10.6151
R978 B.n653 B.n652 10.6151
R979 B.n652 B.n651 10.6151
R980 B.n651 B.n42 10.6151
R981 B.n647 B.n42 10.6151
R982 B.n647 B.n646 10.6151
R983 B.n646 B.n645 10.6151
R984 B.n645 B.n44 10.6151
R985 B.n641 B.n44 10.6151
R986 B.n641 B.n640 10.6151
R987 B.n640 B.n639 10.6151
R988 B.n639 B.n46 10.6151
R989 B.n635 B.n46 10.6151
R990 B.n633 B.n632 10.6151
R991 B.n632 B.n50 10.6151
R992 B.n628 B.n50 10.6151
R993 B.n628 B.n627 10.6151
R994 B.n627 B.n626 10.6151
R995 B.n626 B.n52 10.6151
R996 B.n622 B.n52 10.6151
R997 B.n622 B.n621 10.6151
R998 B.n619 B.n56 10.6151
R999 B.n615 B.n56 10.6151
R1000 B.n615 B.n614 10.6151
R1001 B.n614 B.n613 10.6151
R1002 B.n613 B.n58 10.6151
R1003 B.n609 B.n58 10.6151
R1004 B.n609 B.n608 10.6151
R1005 B.n608 B.n607 10.6151
R1006 B.n607 B.n60 10.6151
R1007 B.n603 B.n60 10.6151
R1008 B.n603 B.n602 10.6151
R1009 B.n602 B.n601 10.6151
R1010 B.n601 B.n62 10.6151
R1011 B.n597 B.n62 10.6151
R1012 B.n597 B.n596 10.6151
R1013 B.n596 B.n595 10.6151
R1014 B.n595 B.n64 10.6151
R1015 B.n591 B.n64 10.6151
R1016 B.n591 B.n590 10.6151
R1017 B.n590 B.n589 10.6151
R1018 B.n589 B.n66 10.6151
R1019 B.n585 B.n66 10.6151
R1020 B.n585 B.n584 10.6151
R1021 B.n584 B.n583 10.6151
R1022 B.n583 B.n68 10.6151
R1023 B.n579 B.n68 10.6151
R1024 B.n391 B.n132 10.6151
R1025 B.n392 B.n391 10.6151
R1026 B.n393 B.n392 10.6151
R1027 B.n393 B.n130 10.6151
R1028 B.n397 B.n130 10.6151
R1029 B.n398 B.n397 10.6151
R1030 B.n399 B.n398 10.6151
R1031 B.n399 B.n128 10.6151
R1032 B.n403 B.n128 10.6151
R1033 B.n404 B.n403 10.6151
R1034 B.n405 B.n404 10.6151
R1035 B.n405 B.n126 10.6151
R1036 B.n409 B.n126 10.6151
R1037 B.n410 B.n409 10.6151
R1038 B.n411 B.n410 10.6151
R1039 B.n411 B.n124 10.6151
R1040 B.n415 B.n124 10.6151
R1041 B.n416 B.n415 10.6151
R1042 B.n417 B.n416 10.6151
R1043 B.n417 B.n122 10.6151
R1044 B.n421 B.n122 10.6151
R1045 B.n422 B.n421 10.6151
R1046 B.n423 B.n422 10.6151
R1047 B.n423 B.n120 10.6151
R1048 B.n427 B.n120 10.6151
R1049 B.n428 B.n427 10.6151
R1050 B.n429 B.n428 10.6151
R1051 B.n429 B.n118 10.6151
R1052 B.n433 B.n118 10.6151
R1053 B.n434 B.n433 10.6151
R1054 B.n435 B.n434 10.6151
R1055 B.n435 B.n116 10.6151
R1056 B.n439 B.n116 10.6151
R1057 B.n440 B.n439 10.6151
R1058 B.n441 B.n440 10.6151
R1059 B.n441 B.n114 10.6151
R1060 B.n445 B.n114 10.6151
R1061 B.n446 B.n445 10.6151
R1062 B.n447 B.n446 10.6151
R1063 B.n447 B.n112 10.6151
R1064 B.n451 B.n112 10.6151
R1065 B.n452 B.n451 10.6151
R1066 B.n453 B.n452 10.6151
R1067 B.n453 B.n110 10.6151
R1068 B.n457 B.n110 10.6151
R1069 B.n458 B.n457 10.6151
R1070 B.n459 B.n458 10.6151
R1071 B.n459 B.n108 10.6151
R1072 B.n463 B.n108 10.6151
R1073 B.n464 B.n463 10.6151
R1074 B.n465 B.n464 10.6151
R1075 B.n465 B.n106 10.6151
R1076 B.n469 B.n106 10.6151
R1077 B.n470 B.n469 10.6151
R1078 B.n471 B.n470 10.6151
R1079 B.n471 B.n104 10.6151
R1080 B.n475 B.n104 10.6151
R1081 B.n476 B.n475 10.6151
R1082 B.n477 B.n476 10.6151
R1083 B.n477 B.n102 10.6151
R1084 B.n481 B.n102 10.6151
R1085 B.n482 B.n481 10.6151
R1086 B.n483 B.n482 10.6151
R1087 B.n483 B.n100 10.6151
R1088 B.n487 B.n100 10.6151
R1089 B.n488 B.n487 10.6151
R1090 B.n489 B.n488 10.6151
R1091 B.n489 B.n98 10.6151
R1092 B.n493 B.n98 10.6151
R1093 B.n494 B.n493 10.6151
R1094 B.n495 B.n494 10.6151
R1095 B.n495 B.n96 10.6151
R1096 B.n499 B.n96 10.6151
R1097 B.n500 B.n499 10.6151
R1098 B.n501 B.n500 10.6151
R1099 B.n501 B.n94 10.6151
R1100 B.n505 B.n94 10.6151
R1101 B.n506 B.n505 10.6151
R1102 B.n507 B.n506 10.6151
R1103 B.n507 B.n92 10.6151
R1104 B.n511 B.n92 10.6151
R1105 B.n512 B.n511 10.6151
R1106 B.n513 B.n512 10.6151
R1107 B.n513 B.n90 10.6151
R1108 B.n517 B.n90 10.6151
R1109 B.n518 B.n517 10.6151
R1110 B.n519 B.n518 10.6151
R1111 B.n519 B.n88 10.6151
R1112 B.n523 B.n88 10.6151
R1113 B.n524 B.n523 10.6151
R1114 B.n525 B.n524 10.6151
R1115 B.n525 B.n86 10.6151
R1116 B.n529 B.n86 10.6151
R1117 B.n530 B.n529 10.6151
R1118 B.n531 B.n530 10.6151
R1119 B.n531 B.n84 10.6151
R1120 B.n535 B.n84 10.6151
R1121 B.n536 B.n535 10.6151
R1122 B.n537 B.n536 10.6151
R1123 B.n537 B.n82 10.6151
R1124 B.n541 B.n82 10.6151
R1125 B.n542 B.n541 10.6151
R1126 B.n543 B.n542 10.6151
R1127 B.n543 B.n80 10.6151
R1128 B.n547 B.n80 10.6151
R1129 B.n548 B.n547 10.6151
R1130 B.n549 B.n548 10.6151
R1131 B.n549 B.n78 10.6151
R1132 B.n553 B.n78 10.6151
R1133 B.n554 B.n553 10.6151
R1134 B.n555 B.n554 10.6151
R1135 B.n555 B.n76 10.6151
R1136 B.n559 B.n76 10.6151
R1137 B.n560 B.n559 10.6151
R1138 B.n561 B.n560 10.6151
R1139 B.n561 B.n74 10.6151
R1140 B.n565 B.n74 10.6151
R1141 B.n566 B.n565 10.6151
R1142 B.n567 B.n566 10.6151
R1143 B.n567 B.n72 10.6151
R1144 B.n571 B.n72 10.6151
R1145 B.n572 B.n571 10.6151
R1146 B.n573 B.n572 10.6151
R1147 B.n573 B.n70 10.6151
R1148 B.n577 B.n70 10.6151
R1149 B.n578 B.n577 10.6151
R1150 B.n295 B.n168 10.6151
R1151 B.n296 B.n295 10.6151
R1152 B.n297 B.n296 10.6151
R1153 B.n297 B.n166 10.6151
R1154 B.n301 B.n166 10.6151
R1155 B.n302 B.n301 10.6151
R1156 B.n303 B.n302 10.6151
R1157 B.n303 B.n164 10.6151
R1158 B.n307 B.n164 10.6151
R1159 B.n308 B.n307 10.6151
R1160 B.n309 B.n308 10.6151
R1161 B.n309 B.n162 10.6151
R1162 B.n313 B.n162 10.6151
R1163 B.n314 B.n313 10.6151
R1164 B.n315 B.n314 10.6151
R1165 B.n315 B.n160 10.6151
R1166 B.n319 B.n160 10.6151
R1167 B.n320 B.n319 10.6151
R1168 B.n321 B.n320 10.6151
R1169 B.n321 B.n158 10.6151
R1170 B.n325 B.n158 10.6151
R1171 B.n326 B.n325 10.6151
R1172 B.n327 B.n326 10.6151
R1173 B.n327 B.n156 10.6151
R1174 B.n331 B.n156 10.6151
R1175 B.n332 B.n331 10.6151
R1176 B.n334 B.n152 10.6151
R1177 B.n338 B.n152 10.6151
R1178 B.n339 B.n338 10.6151
R1179 B.n340 B.n339 10.6151
R1180 B.n340 B.n150 10.6151
R1181 B.n344 B.n150 10.6151
R1182 B.n345 B.n344 10.6151
R1183 B.n346 B.n345 10.6151
R1184 B.n350 B.n349 10.6151
R1185 B.n351 B.n350 10.6151
R1186 B.n351 B.n144 10.6151
R1187 B.n355 B.n144 10.6151
R1188 B.n356 B.n355 10.6151
R1189 B.n357 B.n356 10.6151
R1190 B.n357 B.n142 10.6151
R1191 B.n361 B.n142 10.6151
R1192 B.n362 B.n361 10.6151
R1193 B.n363 B.n362 10.6151
R1194 B.n363 B.n140 10.6151
R1195 B.n367 B.n140 10.6151
R1196 B.n368 B.n367 10.6151
R1197 B.n369 B.n368 10.6151
R1198 B.n369 B.n138 10.6151
R1199 B.n373 B.n138 10.6151
R1200 B.n374 B.n373 10.6151
R1201 B.n375 B.n374 10.6151
R1202 B.n375 B.n136 10.6151
R1203 B.n379 B.n136 10.6151
R1204 B.n380 B.n379 10.6151
R1205 B.n381 B.n380 10.6151
R1206 B.n381 B.n134 10.6151
R1207 B.n385 B.n134 10.6151
R1208 B.n386 B.n385 10.6151
R1209 B.n387 B.n386 10.6151
R1210 B.n291 B.n290 10.6151
R1211 B.n290 B.n289 10.6151
R1212 B.n289 B.n170 10.6151
R1213 B.n285 B.n170 10.6151
R1214 B.n285 B.n284 10.6151
R1215 B.n284 B.n283 10.6151
R1216 B.n283 B.n172 10.6151
R1217 B.n279 B.n172 10.6151
R1218 B.n279 B.n278 10.6151
R1219 B.n278 B.n277 10.6151
R1220 B.n277 B.n174 10.6151
R1221 B.n273 B.n174 10.6151
R1222 B.n273 B.n272 10.6151
R1223 B.n272 B.n271 10.6151
R1224 B.n271 B.n176 10.6151
R1225 B.n267 B.n176 10.6151
R1226 B.n267 B.n266 10.6151
R1227 B.n266 B.n265 10.6151
R1228 B.n265 B.n178 10.6151
R1229 B.n261 B.n178 10.6151
R1230 B.n261 B.n260 10.6151
R1231 B.n260 B.n259 10.6151
R1232 B.n259 B.n180 10.6151
R1233 B.n255 B.n180 10.6151
R1234 B.n255 B.n254 10.6151
R1235 B.n254 B.n253 10.6151
R1236 B.n253 B.n182 10.6151
R1237 B.n249 B.n182 10.6151
R1238 B.n249 B.n248 10.6151
R1239 B.n248 B.n247 10.6151
R1240 B.n247 B.n184 10.6151
R1241 B.n243 B.n184 10.6151
R1242 B.n243 B.n242 10.6151
R1243 B.n242 B.n241 10.6151
R1244 B.n241 B.n186 10.6151
R1245 B.n237 B.n186 10.6151
R1246 B.n237 B.n236 10.6151
R1247 B.n236 B.n235 10.6151
R1248 B.n235 B.n188 10.6151
R1249 B.n231 B.n188 10.6151
R1250 B.n231 B.n230 10.6151
R1251 B.n230 B.n229 10.6151
R1252 B.n229 B.n190 10.6151
R1253 B.n225 B.n190 10.6151
R1254 B.n225 B.n224 10.6151
R1255 B.n224 B.n223 10.6151
R1256 B.n223 B.n192 10.6151
R1257 B.n219 B.n192 10.6151
R1258 B.n219 B.n218 10.6151
R1259 B.n218 B.n217 10.6151
R1260 B.n217 B.n194 10.6151
R1261 B.n213 B.n194 10.6151
R1262 B.n213 B.n212 10.6151
R1263 B.n212 B.n211 10.6151
R1264 B.n211 B.n196 10.6151
R1265 B.n207 B.n196 10.6151
R1266 B.n207 B.n206 10.6151
R1267 B.n206 B.n205 10.6151
R1268 B.n205 B.n198 10.6151
R1269 B.n201 B.n198 10.6151
R1270 B.n201 B.n200 10.6151
R1271 B.n200 B.n0 10.6151
R1272 B.n767 B.n1 10.6151
R1273 B.n767 B.n766 10.6151
R1274 B.n766 B.n765 10.6151
R1275 B.n765 B.n4 10.6151
R1276 B.n761 B.n4 10.6151
R1277 B.n761 B.n760 10.6151
R1278 B.n760 B.n759 10.6151
R1279 B.n759 B.n6 10.6151
R1280 B.n755 B.n6 10.6151
R1281 B.n755 B.n754 10.6151
R1282 B.n754 B.n753 10.6151
R1283 B.n753 B.n8 10.6151
R1284 B.n749 B.n8 10.6151
R1285 B.n749 B.n748 10.6151
R1286 B.n748 B.n747 10.6151
R1287 B.n747 B.n10 10.6151
R1288 B.n743 B.n10 10.6151
R1289 B.n743 B.n742 10.6151
R1290 B.n742 B.n741 10.6151
R1291 B.n741 B.n12 10.6151
R1292 B.n737 B.n12 10.6151
R1293 B.n737 B.n736 10.6151
R1294 B.n736 B.n735 10.6151
R1295 B.n735 B.n14 10.6151
R1296 B.n731 B.n14 10.6151
R1297 B.n731 B.n730 10.6151
R1298 B.n730 B.n729 10.6151
R1299 B.n729 B.n16 10.6151
R1300 B.n725 B.n16 10.6151
R1301 B.n725 B.n724 10.6151
R1302 B.n724 B.n723 10.6151
R1303 B.n723 B.n18 10.6151
R1304 B.n719 B.n18 10.6151
R1305 B.n719 B.n718 10.6151
R1306 B.n718 B.n717 10.6151
R1307 B.n717 B.n20 10.6151
R1308 B.n713 B.n20 10.6151
R1309 B.n713 B.n712 10.6151
R1310 B.n712 B.n711 10.6151
R1311 B.n711 B.n22 10.6151
R1312 B.n707 B.n22 10.6151
R1313 B.n707 B.n706 10.6151
R1314 B.n706 B.n705 10.6151
R1315 B.n705 B.n24 10.6151
R1316 B.n701 B.n24 10.6151
R1317 B.n701 B.n700 10.6151
R1318 B.n700 B.n699 10.6151
R1319 B.n699 B.n26 10.6151
R1320 B.n695 B.n26 10.6151
R1321 B.n695 B.n694 10.6151
R1322 B.n694 B.n693 10.6151
R1323 B.n693 B.n28 10.6151
R1324 B.n689 B.n28 10.6151
R1325 B.n689 B.n688 10.6151
R1326 B.n688 B.n687 10.6151
R1327 B.n687 B.n30 10.6151
R1328 B.n683 B.n30 10.6151
R1329 B.n683 B.n682 10.6151
R1330 B.n682 B.n681 10.6151
R1331 B.n681 B.n32 10.6151
R1332 B.n677 B.n32 10.6151
R1333 B.n677 B.n676 10.6151
R1334 B.n634 B.n633 6.5566
R1335 B.n621 B.n620 6.5566
R1336 B.n334 B.n333 6.5566
R1337 B.n346 B.n148 6.5566
R1338 B.n635 B.n634 4.05904
R1339 B.n620 B.n619 4.05904
R1340 B.n333 B.n332 4.05904
R1341 B.n349 B.n148 4.05904
R1342 B.n771 B.n0 2.81026
R1343 B.n771 B.n1 2.81026
R1344 VN.n68 VN.n67 161.3
R1345 VN.n66 VN.n36 161.3
R1346 VN.n65 VN.n64 161.3
R1347 VN.n63 VN.n37 161.3
R1348 VN.n62 VN.n61 161.3
R1349 VN.n60 VN.n38 161.3
R1350 VN.n59 VN.n58 161.3
R1351 VN.n57 VN.n56 161.3
R1352 VN.n55 VN.n40 161.3
R1353 VN.n54 VN.n53 161.3
R1354 VN.n52 VN.n41 161.3
R1355 VN.n51 VN.n50 161.3
R1356 VN.n49 VN.n42 161.3
R1357 VN.n48 VN.n47 161.3
R1358 VN.n46 VN.n43 161.3
R1359 VN.n33 VN.n32 161.3
R1360 VN.n31 VN.n1 161.3
R1361 VN.n30 VN.n29 161.3
R1362 VN.n28 VN.n2 161.3
R1363 VN.n27 VN.n26 161.3
R1364 VN.n25 VN.n3 161.3
R1365 VN.n24 VN.n23 161.3
R1366 VN.n22 VN.n21 161.3
R1367 VN.n20 VN.n5 161.3
R1368 VN.n19 VN.n18 161.3
R1369 VN.n17 VN.n6 161.3
R1370 VN.n16 VN.n15 161.3
R1371 VN.n14 VN.n7 161.3
R1372 VN.n13 VN.n12 161.3
R1373 VN.n11 VN.n8 161.3
R1374 VN.n45 VN.t4 82.6302
R1375 VN.n10 VN.t0 82.6302
R1376 VN.n34 VN.n0 73.1852
R1377 VN.n69 VN.n35 73.1852
R1378 VN.n10 VN.n9 68.9426
R1379 VN.n45 VN.n44 68.9426
R1380 VN.n15 VN.n6 56.5193
R1381 VN.n50 VN.n41 56.5193
R1382 VN VN.n69 51.1798
R1383 VN.n9 VN.t6 49.5473
R1384 VN.n4 VN.t2 49.5473
R1385 VN.n0 VN.t7 49.5473
R1386 VN.n44 VN.t3 49.5473
R1387 VN.n39 VN.t5 49.5473
R1388 VN.n35 VN.t1 49.5473
R1389 VN.n26 VN.n2 42.4359
R1390 VN.n61 VN.n37 42.4359
R1391 VN.n30 VN.n2 38.5509
R1392 VN.n65 VN.n37 38.5509
R1393 VN.n13 VN.n8 24.4675
R1394 VN.n14 VN.n13 24.4675
R1395 VN.n15 VN.n14 24.4675
R1396 VN.n19 VN.n6 24.4675
R1397 VN.n20 VN.n19 24.4675
R1398 VN.n21 VN.n20 24.4675
R1399 VN.n25 VN.n24 24.4675
R1400 VN.n26 VN.n25 24.4675
R1401 VN.n31 VN.n30 24.4675
R1402 VN.n32 VN.n31 24.4675
R1403 VN.n50 VN.n49 24.4675
R1404 VN.n49 VN.n48 24.4675
R1405 VN.n48 VN.n43 24.4675
R1406 VN.n61 VN.n60 24.4675
R1407 VN.n60 VN.n59 24.4675
R1408 VN.n56 VN.n55 24.4675
R1409 VN.n55 VN.n54 24.4675
R1410 VN.n54 VN.n41 24.4675
R1411 VN.n67 VN.n66 24.4675
R1412 VN.n66 VN.n65 24.4675
R1413 VN.n24 VN.n4 18.8401
R1414 VN.n59 VN.n39 18.8401
R1415 VN.n32 VN.n0 16.8827
R1416 VN.n67 VN.n35 16.8827
R1417 VN.n9 VN.n8 5.62791
R1418 VN.n21 VN.n4 5.62791
R1419 VN.n44 VN.n43 5.62791
R1420 VN.n56 VN.n39 5.62791
R1421 VN.n11 VN.n10 4.0558
R1422 VN.n46 VN.n45 4.05579
R1423 VN.n69 VN.n68 0.354971
R1424 VN.n34 VN.n33 0.354971
R1425 VN VN.n34 0.26696
R1426 VN.n68 VN.n36 0.189894
R1427 VN.n64 VN.n36 0.189894
R1428 VN.n64 VN.n63 0.189894
R1429 VN.n63 VN.n62 0.189894
R1430 VN.n62 VN.n38 0.189894
R1431 VN.n58 VN.n38 0.189894
R1432 VN.n58 VN.n57 0.189894
R1433 VN.n57 VN.n40 0.189894
R1434 VN.n53 VN.n40 0.189894
R1435 VN.n53 VN.n52 0.189894
R1436 VN.n52 VN.n51 0.189894
R1437 VN.n51 VN.n42 0.189894
R1438 VN.n47 VN.n42 0.189894
R1439 VN.n47 VN.n46 0.189894
R1440 VN.n12 VN.n11 0.189894
R1441 VN.n12 VN.n7 0.189894
R1442 VN.n16 VN.n7 0.189894
R1443 VN.n17 VN.n16 0.189894
R1444 VN.n18 VN.n17 0.189894
R1445 VN.n18 VN.n5 0.189894
R1446 VN.n22 VN.n5 0.189894
R1447 VN.n23 VN.n22 0.189894
R1448 VN.n23 VN.n3 0.189894
R1449 VN.n27 VN.n3 0.189894
R1450 VN.n28 VN.n27 0.189894
R1451 VN.n29 VN.n28 0.189894
R1452 VN.n29 VN.n1 0.189894
R1453 VN.n33 VN.n1 0.189894
R1454 VDD2.n2 VDD2.n1 86.573
R1455 VDD2.n2 VDD2.n0 86.573
R1456 VDD2 VDD2.n5 86.5701
R1457 VDD2.n4 VDD2.n3 85.0207
R1458 VDD2.n4 VDD2.n2 44.211
R1459 VDD2.n5 VDD2.t4 4.65071
R1460 VDD2.n5 VDD2.t3 4.65071
R1461 VDD2.n3 VDD2.t6 4.65071
R1462 VDD2.n3 VDD2.t2 4.65071
R1463 VDD2.n1 VDD2.t5 4.65071
R1464 VDD2.n1 VDD2.t0 4.65071
R1465 VDD2.n0 VDD2.t7 4.65071
R1466 VDD2.n0 VDD2.t1 4.65071
R1467 VDD2 VDD2.n4 1.66645
C0 w_n4700_n2366# VP 10.3037f
C1 VN VDD2 5.50789f
C2 B VDD2 1.87979f
C3 VTAIL VDD1 6.910181f
C4 VP VDD2 0.604402f
C5 w_n4700_n2366# VTAIL 3.18544f
C6 VTAIL VDD2 6.96996f
C7 VN B 1.3517f
C8 w_n4700_n2366# VDD1 2.07162f
C9 VN VP 7.71117f
C10 VP B 2.38275f
C11 VDD1 VDD2 2.1888f
C12 w_n4700_n2366# VDD2 2.21988f
C13 VTAIL VN 6.6043f
C14 VTAIL B 3.60778f
C15 VTAIL VP 6.61841f
C16 VN VDD1 0.152777f
C17 w_n4700_n2366# VN 9.69122f
C18 B VDD1 1.75859f
C19 w_n4700_n2366# B 9.939361f
C20 VP VDD1 5.95771f
C21 VDD2 VSUBS 2.195341f
C22 VDD1 VSUBS 2.99273f
C23 VTAIL VSUBS 0.810491f
C24 VN VSUBS 7.55879f
C25 VP VSUBS 4.004187f
C26 B VSUBS 5.473161f
C27 w_n4700_n2366# VSUBS 0.138349p
C28 VDD2.t7 VSUBS 0.180181f
C29 VDD2.t1 VSUBS 0.180181f
C30 VDD2.n0 VSUBS 1.25801f
C31 VDD2.t5 VSUBS 0.180181f
C32 VDD2.t0 VSUBS 0.180181f
C33 VDD2.n1 VSUBS 1.25801f
C34 VDD2.n2 VSUBS 5.05304f
C35 VDD2.t6 VSUBS 0.180181f
C36 VDD2.t2 VSUBS 0.180181f
C37 VDD2.n3 VSUBS 1.23876f
C38 VDD2.n4 VSUBS 4.00132f
C39 VDD2.t4 VSUBS 0.180181f
C40 VDD2.t3 VSUBS 0.180181f
C41 VDD2.n5 VSUBS 1.25796f
C42 VN.t7 VSUBS 1.95645f
C43 VN.n0 VSUBS 0.842475f
C44 VN.n1 VSUBS 0.030846f
C45 VN.n2 VSUBS 0.025095f
C46 VN.n3 VSUBS 0.030846f
C47 VN.t2 VSUBS 1.95645f
C48 VN.n4 VSUBS 0.713186f
C49 VN.n5 VSUBS 0.030846f
C50 VN.n6 VSUBS 0.045029f
C51 VN.n7 VSUBS 0.030846f
C52 VN.n8 VSUBS 0.035632f
C53 VN.t6 VSUBS 1.95645f
C54 VN.n9 VSUBS 0.810856f
C55 VN.t0 VSUBS 2.33302f
C56 VN.n10 VSUBS 0.773099f
C57 VN.n11 VSUBS 0.364906f
C58 VN.n12 VSUBS 0.030846f
C59 VN.n13 VSUBS 0.057488f
C60 VN.n14 VSUBS 0.057488f
C61 VN.n15 VSUBS 0.045029f
C62 VN.n16 VSUBS 0.030846f
C63 VN.n17 VSUBS 0.030846f
C64 VN.n18 VSUBS 0.030846f
C65 VN.n19 VSUBS 0.057488f
C66 VN.n20 VSUBS 0.057488f
C67 VN.n21 VSUBS 0.035632f
C68 VN.n22 VSUBS 0.030846f
C69 VN.n23 VSUBS 0.030846f
C70 VN.n24 VSUBS 0.050959f
C71 VN.n25 VSUBS 0.057488f
C72 VN.n26 VSUBS 0.060611f
C73 VN.n27 VSUBS 0.030846f
C74 VN.n28 VSUBS 0.030846f
C75 VN.n29 VSUBS 0.030846f
C76 VN.n30 VSUBS 0.061841f
C77 VN.n31 VSUBS 0.057488f
C78 VN.n32 VSUBS 0.048688f
C79 VN.n33 VSUBS 0.049784f
C80 VN.n34 VSUBS 0.072939f
C81 VN.t1 VSUBS 1.95645f
C82 VN.n35 VSUBS 0.842475f
C83 VN.n36 VSUBS 0.030846f
C84 VN.n37 VSUBS 0.025095f
C85 VN.n38 VSUBS 0.030846f
C86 VN.t5 VSUBS 1.95645f
C87 VN.n39 VSUBS 0.713186f
C88 VN.n40 VSUBS 0.030846f
C89 VN.n41 VSUBS 0.045029f
C90 VN.n42 VSUBS 0.030846f
C91 VN.n43 VSUBS 0.035632f
C92 VN.t4 VSUBS 2.33302f
C93 VN.t3 VSUBS 1.95645f
C94 VN.n44 VSUBS 0.810856f
C95 VN.n45 VSUBS 0.773099f
C96 VN.n46 VSUBS 0.364906f
C97 VN.n47 VSUBS 0.030846f
C98 VN.n48 VSUBS 0.057488f
C99 VN.n49 VSUBS 0.057488f
C100 VN.n50 VSUBS 0.045029f
C101 VN.n51 VSUBS 0.030846f
C102 VN.n52 VSUBS 0.030846f
C103 VN.n53 VSUBS 0.030846f
C104 VN.n54 VSUBS 0.057488f
C105 VN.n55 VSUBS 0.057488f
C106 VN.n56 VSUBS 0.035632f
C107 VN.n57 VSUBS 0.030846f
C108 VN.n58 VSUBS 0.030846f
C109 VN.n59 VSUBS 0.050959f
C110 VN.n60 VSUBS 0.057488f
C111 VN.n61 VSUBS 0.060611f
C112 VN.n62 VSUBS 0.030846f
C113 VN.n63 VSUBS 0.030846f
C114 VN.n64 VSUBS 0.030846f
C115 VN.n65 VSUBS 0.061841f
C116 VN.n66 VSUBS 0.057488f
C117 VN.n67 VSUBS 0.048688f
C118 VN.n68 VSUBS 0.049784f
C119 VN.n69 VSUBS 1.81886f
C120 B.n0 VSUBS 0.005542f
C121 B.n1 VSUBS 0.005542f
C122 B.n2 VSUBS 0.008764f
C123 B.n3 VSUBS 0.008764f
C124 B.n4 VSUBS 0.008764f
C125 B.n5 VSUBS 0.008764f
C126 B.n6 VSUBS 0.008764f
C127 B.n7 VSUBS 0.008764f
C128 B.n8 VSUBS 0.008764f
C129 B.n9 VSUBS 0.008764f
C130 B.n10 VSUBS 0.008764f
C131 B.n11 VSUBS 0.008764f
C132 B.n12 VSUBS 0.008764f
C133 B.n13 VSUBS 0.008764f
C134 B.n14 VSUBS 0.008764f
C135 B.n15 VSUBS 0.008764f
C136 B.n16 VSUBS 0.008764f
C137 B.n17 VSUBS 0.008764f
C138 B.n18 VSUBS 0.008764f
C139 B.n19 VSUBS 0.008764f
C140 B.n20 VSUBS 0.008764f
C141 B.n21 VSUBS 0.008764f
C142 B.n22 VSUBS 0.008764f
C143 B.n23 VSUBS 0.008764f
C144 B.n24 VSUBS 0.008764f
C145 B.n25 VSUBS 0.008764f
C146 B.n26 VSUBS 0.008764f
C147 B.n27 VSUBS 0.008764f
C148 B.n28 VSUBS 0.008764f
C149 B.n29 VSUBS 0.008764f
C150 B.n30 VSUBS 0.008764f
C151 B.n31 VSUBS 0.008764f
C152 B.n32 VSUBS 0.008764f
C153 B.n33 VSUBS 0.020704f
C154 B.n34 VSUBS 0.008764f
C155 B.n35 VSUBS 0.008764f
C156 B.n36 VSUBS 0.008764f
C157 B.n37 VSUBS 0.008764f
C158 B.n38 VSUBS 0.008764f
C159 B.n39 VSUBS 0.008764f
C160 B.n40 VSUBS 0.008764f
C161 B.n41 VSUBS 0.008764f
C162 B.n42 VSUBS 0.008764f
C163 B.n43 VSUBS 0.008764f
C164 B.n44 VSUBS 0.008764f
C165 B.n45 VSUBS 0.008764f
C166 B.n46 VSUBS 0.008764f
C167 B.n47 VSUBS 0.008764f
C168 B.t5 VSUBS 0.263566f
C169 B.t4 VSUBS 0.295055f
C170 B.t3 VSUBS 1.41555f
C171 B.n48 VSUBS 0.173495f
C172 B.n49 VSUBS 0.093307f
C173 B.n50 VSUBS 0.008764f
C174 B.n51 VSUBS 0.008764f
C175 B.n52 VSUBS 0.008764f
C176 B.n53 VSUBS 0.008764f
C177 B.t8 VSUBS 0.263565f
C178 B.t7 VSUBS 0.295053f
C179 B.t6 VSUBS 1.41555f
C180 B.n54 VSUBS 0.173497f
C181 B.n55 VSUBS 0.093309f
C182 B.n56 VSUBS 0.008764f
C183 B.n57 VSUBS 0.008764f
C184 B.n58 VSUBS 0.008764f
C185 B.n59 VSUBS 0.008764f
C186 B.n60 VSUBS 0.008764f
C187 B.n61 VSUBS 0.008764f
C188 B.n62 VSUBS 0.008764f
C189 B.n63 VSUBS 0.008764f
C190 B.n64 VSUBS 0.008764f
C191 B.n65 VSUBS 0.008764f
C192 B.n66 VSUBS 0.008764f
C193 B.n67 VSUBS 0.008764f
C194 B.n68 VSUBS 0.008764f
C195 B.n69 VSUBS 0.020704f
C196 B.n70 VSUBS 0.008764f
C197 B.n71 VSUBS 0.008764f
C198 B.n72 VSUBS 0.008764f
C199 B.n73 VSUBS 0.008764f
C200 B.n74 VSUBS 0.008764f
C201 B.n75 VSUBS 0.008764f
C202 B.n76 VSUBS 0.008764f
C203 B.n77 VSUBS 0.008764f
C204 B.n78 VSUBS 0.008764f
C205 B.n79 VSUBS 0.008764f
C206 B.n80 VSUBS 0.008764f
C207 B.n81 VSUBS 0.008764f
C208 B.n82 VSUBS 0.008764f
C209 B.n83 VSUBS 0.008764f
C210 B.n84 VSUBS 0.008764f
C211 B.n85 VSUBS 0.008764f
C212 B.n86 VSUBS 0.008764f
C213 B.n87 VSUBS 0.008764f
C214 B.n88 VSUBS 0.008764f
C215 B.n89 VSUBS 0.008764f
C216 B.n90 VSUBS 0.008764f
C217 B.n91 VSUBS 0.008764f
C218 B.n92 VSUBS 0.008764f
C219 B.n93 VSUBS 0.008764f
C220 B.n94 VSUBS 0.008764f
C221 B.n95 VSUBS 0.008764f
C222 B.n96 VSUBS 0.008764f
C223 B.n97 VSUBS 0.008764f
C224 B.n98 VSUBS 0.008764f
C225 B.n99 VSUBS 0.008764f
C226 B.n100 VSUBS 0.008764f
C227 B.n101 VSUBS 0.008764f
C228 B.n102 VSUBS 0.008764f
C229 B.n103 VSUBS 0.008764f
C230 B.n104 VSUBS 0.008764f
C231 B.n105 VSUBS 0.008764f
C232 B.n106 VSUBS 0.008764f
C233 B.n107 VSUBS 0.008764f
C234 B.n108 VSUBS 0.008764f
C235 B.n109 VSUBS 0.008764f
C236 B.n110 VSUBS 0.008764f
C237 B.n111 VSUBS 0.008764f
C238 B.n112 VSUBS 0.008764f
C239 B.n113 VSUBS 0.008764f
C240 B.n114 VSUBS 0.008764f
C241 B.n115 VSUBS 0.008764f
C242 B.n116 VSUBS 0.008764f
C243 B.n117 VSUBS 0.008764f
C244 B.n118 VSUBS 0.008764f
C245 B.n119 VSUBS 0.008764f
C246 B.n120 VSUBS 0.008764f
C247 B.n121 VSUBS 0.008764f
C248 B.n122 VSUBS 0.008764f
C249 B.n123 VSUBS 0.008764f
C250 B.n124 VSUBS 0.008764f
C251 B.n125 VSUBS 0.008764f
C252 B.n126 VSUBS 0.008764f
C253 B.n127 VSUBS 0.008764f
C254 B.n128 VSUBS 0.008764f
C255 B.n129 VSUBS 0.008764f
C256 B.n130 VSUBS 0.008764f
C257 B.n131 VSUBS 0.008764f
C258 B.n132 VSUBS 0.020704f
C259 B.n133 VSUBS 0.008764f
C260 B.n134 VSUBS 0.008764f
C261 B.n135 VSUBS 0.008764f
C262 B.n136 VSUBS 0.008764f
C263 B.n137 VSUBS 0.008764f
C264 B.n138 VSUBS 0.008764f
C265 B.n139 VSUBS 0.008764f
C266 B.n140 VSUBS 0.008764f
C267 B.n141 VSUBS 0.008764f
C268 B.n142 VSUBS 0.008764f
C269 B.n143 VSUBS 0.008764f
C270 B.n144 VSUBS 0.008764f
C271 B.n145 VSUBS 0.008764f
C272 B.t10 VSUBS 0.263565f
C273 B.t11 VSUBS 0.295053f
C274 B.t9 VSUBS 1.41555f
C275 B.n146 VSUBS 0.173497f
C276 B.n147 VSUBS 0.093309f
C277 B.n148 VSUBS 0.020306f
C278 B.n149 VSUBS 0.008764f
C279 B.n150 VSUBS 0.008764f
C280 B.n151 VSUBS 0.008764f
C281 B.n152 VSUBS 0.008764f
C282 B.n153 VSUBS 0.008764f
C283 B.t1 VSUBS 0.263566f
C284 B.t2 VSUBS 0.295055f
C285 B.t0 VSUBS 1.41555f
C286 B.n154 VSUBS 0.173495f
C287 B.n155 VSUBS 0.093307f
C288 B.n156 VSUBS 0.008764f
C289 B.n157 VSUBS 0.008764f
C290 B.n158 VSUBS 0.008764f
C291 B.n159 VSUBS 0.008764f
C292 B.n160 VSUBS 0.008764f
C293 B.n161 VSUBS 0.008764f
C294 B.n162 VSUBS 0.008764f
C295 B.n163 VSUBS 0.008764f
C296 B.n164 VSUBS 0.008764f
C297 B.n165 VSUBS 0.008764f
C298 B.n166 VSUBS 0.008764f
C299 B.n167 VSUBS 0.008764f
C300 B.n168 VSUBS 0.021313f
C301 B.n169 VSUBS 0.008764f
C302 B.n170 VSUBS 0.008764f
C303 B.n171 VSUBS 0.008764f
C304 B.n172 VSUBS 0.008764f
C305 B.n173 VSUBS 0.008764f
C306 B.n174 VSUBS 0.008764f
C307 B.n175 VSUBS 0.008764f
C308 B.n176 VSUBS 0.008764f
C309 B.n177 VSUBS 0.008764f
C310 B.n178 VSUBS 0.008764f
C311 B.n179 VSUBS 0.008764f
C312 B.n180 VSUBS 0.008764f
C313 B.n181 VSUBS 0.008764f
C314 B.n182 VSUBS 0.008764f
C315 B.n183 VSUBS 0.008764f
C316 B.n184 VSUBS 0.008764f
C317 B.n185 VSUBS 0.008764f
C318 B.n186 VSUBS 0.008764f
C319 B.n187 VSUBS 0.008764f
C320 B.n188 VSUBS 0.008764f
C321 B.n189 VSUBS 0.008764f
C322 B.n190 VSUBS 0.008764f
C323 B.n191 VSUBS 0.008764f
C324 B.n192 VSUBS 0.008764f
C325 B.n193 VSUBS 0.008764f
C326 B.n194 VSUBS 0.008764f
C327 B.n195 VSUBS 0.008764f
C328 B.n196 VSUBS 0.008764f
C329 B.n197 VSUBS 0.008764f
C330 B.n198 VSUBS 0.008764f
C331 B.n199 VSUBS 0.008764f
C332 B.n200 VSUBS 0.008764f
C333 B.n201 VSUBS 0.008764f
C334 B.n202 VSUBS 0.008764f
C335 B.n203 VSUBS 0.008764f
C336 B.n204 VSUBS 0.008764f
C337 B.n205 VSUBS 0.008764f
C338 B.n206 VSUBS 0.008764f
C339 B.n207 VSUBS 0.008764f
C340 B.n208 VSUBS 0.008764f
C341 B.n209 VSUBS 0.008764f
C342 B.n210 VSUBS 0.008764f
C343 B.n211 VSUBS 0.008764f
C344 B.n212 VSUBS 0.008764f
C345 B.n213 VSUBS 0.008764f
C346 B.n214 VSUBS 0.008764f
C347 B.n215 VSUBS 0.008764f
C348 B.n216 VSUBS 0.008764f
C349 B.n217 VSUBS 0.008764f
C350 B.n218 VSUBS 0.008764f
C351 B.n219 VSUBS 0.008764f
C352 B.n220 VSUBS 0.008764f
C353 B.n221 VSUBS 0.008764f
C354 B.n222 VSUBS 0.008764f
C355 B.n223 VSUBS 0.008764f
C356 B.n224 VSUBS 0.008764f
C357 B.n225 VSUBS 0.008764f
C358 B.n226 VSUBS 0.008764f
C359 B.n227 VSUBS 0.008764f
C360 B.n228 VSUBS 0.008764f
C361 B.n229 VSUBS 0.008764f
C362 B.n230 VSUBS 0.008764f
C363 B.n231 VSUBS 0.008764f
C364 B.n232 VSUBS 0.008764f
C365 B.n233 VSUBS 0.008764f
C366 B.n234 VSUBS 0.008764f
C367 B.n235 VSUBS 0.008764f
C368 B.n236 VSUBS 0.008764f
C369 B.n237 VSUBS 0.008764f
C370 B.n238 VSUBS 0.008764f
C371 B.n239 VSUBS 0.008764f
C372 B.n240 VSUBS 0.008764f
C373 B.n241 VSUBS 0.008764f
C374 B.n242 VSUBS 0.008764f
C375 B.n243 VSUBS 0.008764f
C376 B.n244 VSUBS 0.008764f
C377 B.n245 VSUBS 0.008764f
C378 B.n246 VSUBS 0.008764f
C379 B.n247 VSUBS 0.008764f
C380 B.n248 VSUBS 0.008764f
C381 B.n249 VSUBS 0.008764f
C382 B.n250 VSUBS 0.008764f
C383 B.n251 VSUBS 0.008764f
C384 B.n252 VSUBS 0.008764f
C385 B.n253 VSUBS 0.008764f
C386 B.n254 VSUBS 0.008764f
C387 B.n255 VSUBS 0.008764f
C388 B.n256 VSUBS 0.008764f
C389 B.n257 VSUBS 0.008764f
C390 B.n258 VSUBS 0.008764f
C391 B.n259 VSUBS 0.008764f
C392 B.n260 VSUBS 0.008764f
C393 B.n261 VSUBS 0.008764f
C394 B.n262 VSUBS 0.008764f
C395 B.n263 VSUBS 0.008764f
C396 B.n264 VSUBS 0.008764f
C397 B.n265 VSUBS 0.008764f
C398 B.n266 VSUBS 0.008764f
C399 B.n267 VSUBS 0.008764f
C400 B.n268 VSUBS 0.008764f
C401 B.n269 VSUBS 0.008764f
C402 B.n270 VSUBS 0.008764f
C403 B.n271 VSUBS 0.008764f
C404 B.n272 VSUBS 0.008764f
C405 B.n273 VSUBS 0.008764f
C406 B.n274 VSUBS 0.008764f
C407 B.n275 VSUBS 0.008764f
C408 B.n276 VSUBS 0.008764f
C409 B.n277 VSUBS 0.008764f
C410 B.n278 VSUBS 0.008764f
C411 B.n279 VSUBS 0.008764f
C412 B.n280 VSUBS 0.008764f
C413 B.n281 VSUBS 0.008764f
C414 B.n282 VSUBS 0.008764f
C415 B.n283 VSUBS 0.008764f
C416 B.n284 VSUBS 0.008764f
C417 B.n285 VSUBS 0.008764f
C418 B.n286 VSUBS 0.008764f
C419 B.n287 VSUBS 0.008764f
C420 B.n288 VSUBS 0.008764f
C421 B.n289 VSUBS 0.008764f
C422 B.n290 VSUBS 0.008764f
C423 B.n291 VSUBS 0.020704f
C424 B.n292 VSUBS 0.020704f
C425 B.n293 VSUBS 0.021313f
C426 B.n294 VSUBS 0.008764f
C427 B.n295 VSUBS 0.008764f
C428 B.n296 VSUBS 0.008764f
C429 B.n297 VSUBS 0.008764f
C430 B.n298 VSUBS 0.008764f
C431 B.n299 VSUBS 0.008764f
C432 B.n300 VSUBS 0.008764f
C433 B.n301 VSUBS 0.008764f
C434 B.n302 VSUBS 0.008764f
C435 B.n303 VSUBS 0.008764f
C436 B.n304 VSUBS 0.008764f
C437 B.n305 VSUBS 0.008764f
C438 B.n306 VSUBS 0.008764f
C439 B.n307 VSUBS 0.008764f
C440 B.n308 VSUBS 0.008764f
C441 B.n309 VSUBS 0.008764f
C442 B.n310 VSUBS 0.008764f
C443 B.n311 VSUBS 0.008764f
C444 B.n312 VSUBS 0.008764f
C445 B.n313 VSUBS 0.008764f
C446 B.n314 VSUBS 0.008764f
C447 B.n315 VSUBS 0.008764f
C448 B.n316 VSUBS 0.008764f
C449 B.n317 VSUBS 0.008764f
C450 B.n318 VSUBS 0.008764f
C451 B.n319 VSUBS 0.008764f
C452 B.n320 VSUBS 0.008764f
C453 B.n321 VSUBS 0.008764f
C454 B.n322 VSUBS 0.008764f
C455 B.n323 VSUBS 0.008764f
C456 B.n324 VSUBS 0.008764f
C457 B.n325 VSUBS 0.008764f
C458 B.n326 VSUBS 0.008764f
C459 B.n327 VSUBS 0.008764f
C460 B.n328 VSUBS 0.008764f
C461 B.n329 VSUBS 0.008764f
C462 B.n330 VSUBS 0.008764f
C463 B.n331 VSUBS 0.008764f
C464 B.n332 VSUBS 0.006058f
C465 B.n333 VSUBS 0.020306f
C466 B.n334 VSUBS 0.007089f
C467 B.n335 VSUBS 0.008764f
C468 B.n336 VSUBS 0.008764f
C469 B.n337 VSUBS 0.008764f
C470 B.n338 VSUBS 0.008764f
C471 B.n339 VSUBS 0.008764f
C472 B.n340 VSUBS 0.008764f
C473 B.n341 VSUBS 0.008764f
C474 B.n342 VSUBS 0.008764f
C475 B.n343 VSUBS 0.008764f
C476 B.n344 VSUBS 0.008764f
C477 B.n345 VSUBS 0.008764f
C478 B.n346 VSUBS 0.007089f
C479 B.n347 VSUBS 0.008764f
C480 B.n348 VSUBS 0.008764f
C481 B.n349 VSUBS 0.006058f
C482 B.n350 VSUBS 0.008764f
C483 B.n351 VSUBS 0.008764f
C484 B.n352 VSUBS 0.008764f
C485 B.n353 VSUBS 0.008764f
C486 B.n354 VSUBS 0.008764f
C487 B.n355 VSUBS 0.008764f
C488 B.n356 VSUBS 0.008764f
C489 B.n357 VSUBS 0.008764f
C490 B.n358 VSUBS 0.008764f
C491 B.n359 VSUBS 0.008764f
C492 B.n360 VSUBS 0.008764f
C493 B.n361 VSUBS 0.008764f
C494 B.n362 VSUBS 0.008764f
C495 B.n363 VSUBS 0.008764f
C496 B.n364 VSUBS 0.008764f
C497 B.n365 VSUBS 0.008764f
C498 B.n366 VSUBS 0.008764f
C499 B.n367 VSUBS 0.008764f
C500 B.n368 VSUBS 0.008764f
C501 B.n369 VSUBS 0.008764f
C502 B.n370 VSUBS 0.008764f
C503 B.n371 VSUBS 0.008764f
C504 B.n372 VSUBS 0.008764f
C505 B.n373 VSUBS 0.008764f
C506 B.n374 VSUBS 0.008764f
C507 B.n375 VSUBS 0.008764f
C508 B.n376 VSUBS 0.008764f
C509 B.n377 VSUBS 0.008764f
C510 B.n378 VSUBS 0.008764f
C511 B.n379 VSUBS 0.008764f
C512 B.n380 VSUBS 0.008764f
C513 B.n381 VSUBS 0.008764f
C514 B.n382 VSUBS 0.008764f
C515 B.n383 VSUBS 0.008764f
C516 B.n384 VSUBS 0.008764f
C517 B.n385 VSUBS 0.008764f
C518 B.n386 VSUBS 0.008764f
C519 B.n387 VSUBS 0.021313f
C520 B.n388 VSUBS 0.021313f
C521 B.n389 VSUBS 0.020704f
C522 B.n390 VSUBS 0.008764f
C523 B.n391 VSUBS 0.008764f
C524 B.n392 VSUBS 0.008764f
C525 B.n393 VSUBS 0.008764f
C526 B.n394 VSUBS 0.008764f
C527 B.n395 VSUBS 0.008764f
C528 B.n396 VSUBS 0.008764f
C529 B.n397 VSUBS 0.008764f
C530 B.n398 VSUBS 0.008764f
C531 B.n399 VSUBS 0.008764f
C532 B.n400 VSUBS 0.008764f
C533 B.n401 VSUBS 0.008764f
C534 B.n402 VSUBS 0.008764f
C535 B.n403 VSUBS 0.008764f
C536 B.n404 VSUBS 0.008764f
C537 B.n405 VSUBS 0.008764f
C538 B.n406 VSUBS 0.008764f
C539 B.n407 VSUBS 0.008764f
C540 B.n408 VSUBS 0.008764f
C541 B.n409 VSUBS 0.008764f
C542 B.n410 VSUBS 0.008764f
C543 B.n411 VSUBS 0.008764f
C544 B.n412 VSUBS 0.008764f
C545 B.n413 VSUBS 0.008764f
C546 B.n414 VSUBS 0.008764f
C547 B.n415 VSUBS 0.008764f
C548 B.n416 VSUBS 0.008764f
C549 B.n417 VSUBS 0.008764f
C550 B.n418 VSUBS 0.008764f
C551 B.n419 VSUBS 0.008764f
C552 B.n420 VSUBS 0.008764f
C553 B.n421 VSUBS 0.008764f
C554 B.n422 VSUBS 0.008764f
C555 B.n423 VSUBS 0.008764f
C556 B.n424 VSUBS 0.008764f
C557 B.n425 VSUBS 0.008764f
C558 B.n426 VSUBS 0.008764f
C559 B.n427 VSUBS 0.008764f
C560 B.n428 VSUBS 0.008764f
C561 B.n429 VSUBS 0.008764f
C562 B.n430 VSUBS 0.008764f
C563 B.n431 VSUBS 0.008764f
C564 B.n432 VSUBS 0.008764f
C565 B.n433 VSUBS 0.008764f
C566 B.n434 VSUBS 0.008764f
C567 B.n435 VSUBS 0.008764f
C568 B.n436 VSUBS 0.008764f
C569 B.n437 VSUBS 0.008764f
C570 B.n438 VSUBS 0.008764f
C571 B.n439 VSUBS 0.008764f
C572 B.n440 VSUBS 0.008764f
C573 B.n441 VSUBS 0.008764f
C574 B.n442 VSUBS 0.008764f
C575 B.n443 VSUBS 0.008764f
C576 B.n444 VSUBS 0.008764f
C577 B.n445 VSUBS 0.008764f
C578 B.n446 VSUBS 0.008764f
C579 B.n447 VSUBS 0.008764f
C580 B.n448 VSUBS 0.008764f
C581 B.n449 VSUBS 0.008764f
C582 B.n450 VSUBS 0.008764f
C583 B.n451 VSUBS 0.008764f
C584 B.n452 VSUBS 0.008764f
C585 B.n453 VSUBS 0.008764f
C586 B.n454 VSUBS 0.008764f
C587 B.n455 VSUBS 0.008764f
C588 B.n456 VSUBS 0.008764f
C589 B.n457 VSUBS 0.008764f
C590 B.n458 VSUBS 0.008764f
C591 B.n459 VSUBS 0.008764f
C592 B.n460 VSUBS 0.008764f
C593 B.n461 VSUBS 0.008764f
C594 B.n462 VSUBS 0.008764f
C595 B.n463 VSUBS 0.008764f
C596 B.n464 VSUBS 0.008764f
C597 B.n465 VSUBS 0.008764f
C598 B.n466 VSUBS 0.008764f
C599 B.n467 VSUBS 0.008764f
C600 B.n468 VSUBS 0.008764f
C601 B.n469 VSUBS 0.008764f
C602 B.n470 VSUBS 0.008764f
C603 B.n471 VSUBS 0.008764f
C604 B.n472 VSUBS 0.008764f
C605 B.n473 VSUBS 0.008764f
C606 B.n474 VSUBS 0.008764f
C607 B.n475 VSUBS 0.008764f
C608 B.n476 VSUBS 0.008764f
C609 B.n477 VSUBS 0.008764f
C610 B.n478 VSUBS 0.008764f
C611 B.n479 VSUBS 0.008764f
C612 B.n480 VSUBS 0.008764f
C613 B.n481 VSUBS 0.008764f
C614 B.n482 VSUBS 0.008764f
C615 B.n483 VSUBS 0.008764f
C616 B.n484 VSUBS 0.008764f
C617 B.n485 VSUBS 0.008764f
C618 B.n486 VSUBS 0.008764f
C619 B.n487 VSUBS 0.008764f
C620 B.n488 VSUBS 0.008764f
C621 B.n489 VSUBS 0.008764f
C622 B.n490 VSUBS 0.008764f
C623 B.n491 VSUBS 0.008764f
C624 B.n492 VSUBS 0.008764f
C625 B.n493 VSUBS 0.008764f
C626 B.n494 VSUBS 0.008764f
C627 B.n495 VSUBS 0.008764f
C628 B.n496 VSUBS 0.008764f
C629 B.n497 VSUBS 0.008764f
C630 B.n498 VSUBS 0.008764f
C631 B.n499 VSUBS 0.008764f
C632 B.n500 VSUBS 0.008764f
C633 B.n501 VSUBS 0.008764f
C634 B.n502 VSUBS 0.008764f
C635 B.n503 VSUBS 0.008764f
C636 B.n504 VSUBS 0.008764f
C637 B.n505 VSUBS 0.008764f
C638 B.n506 VSUBS 0.008764f
C639 B.n507 VSUBS 0.008764f
C640 B.n508 VSUBS 0.008764f
C641 B.n509 VSUBS 0.008764f
C642 B.n510 VSUBS 0.008764f
C643 B.n511 VSUBS 0.008764f
C644 B.n512 VSUBS 0.008764f
C645 B.n513 VSUBS 0.008764f
C646 B.n514 VSUBS 0.008764f
C647 B.n515 VSUBS 0.008764f
C648 B.n516 VSUBS 0.008764f
C649 B.n517 VSUBS 0.008764f
C650 B.n518 VSUBS 0.008764f
C651 B.n519 VSUBS 0.008764f
C652 B.n520 VSUBS 0.008764f
C653 B.n521 VSUBS 0.008764f
C654 B.n522 VSUBS 0.008764f
C655 B.n523 VSUBS 0.008764f
C656 B.n524 VSUBS 0.008764f
C657 B.n525 VSUBS 0.008764f
C658 B.n526 VSUBS 0.008764f
C659 B.n527 VSUBS 0.008764f
C660 B.n528 VSUBS 0.008764f
C661 B.n529 VSUBS 0.008764f
C662 B.n530 VSUBS 0.008764f
C663 B.n531 VSUBS 0.008764f
C664 B.n532 VSUBS 0.008764f
C665 B.n533 VSUBS 0.008764f
C666 B.n534 VSUBS 0.008764f
C667 B.n535 VSUBS 0.008764f
C668 B.n536 VSUBS 0.008764f
C669 B.n537 VSUBS 0.008764f
C670 B.n538 VSUBS 0.008764f
C671 B.n539 VSUBS 0.008764f
C672 B.n540 VSUBS 0.008764f
C673 B.n541 VSUBS 0.008764f
C674 B.n542 VSUBS 0.008764f
C675 B.n543 VSUBS 0.008764f
C676 B.n544 VSUBS 0.008764f
C677 B.n545 VSUBS 0.008764f
C678 B.n546 VSUBS 0.008764f
C679 B.n547 VSUBS 0.008764f
C680 B.n548 VSUBS 0.008764f
C681 B.n549 VSUBS 0.008764f
C682 B.n550 VSUBS 0.008764f
C683 B.n551 VSUBS 0.008764f
C684 B.n552 VSUBS 0.008764f
C685 B.n553 VSUBS 0.008764f
C686 B.n554 VSUBS 0.008764f
C687 B.n555 VSUBS 0.008764f
C688 B.n556 VSUBS 0.008764f
C689 B.n557 VSUBS 0.008764f
C690 B.n558 VSUBS 0.008764f
C691 B.n559 VSUBS 0.008764f
C692 B.n560 VSUBS 0.008764f
C693 B.n561 VSUBS 0.008764f
C694 B.n562 VSUBS 0.008764f
C695 B.n563 VSUBS 0.008764f
C696 B.n564 VSUBS 0.008764f
C697 B.n565 VSUBS 0.008764f
C698 B.n566 VSUBS 0.008764f
C699 B.n567 VSUBS 0.008764f
C700 B.n568 VSUBS 0.008764f
C701 B.n569 VSUBS 0.008764f
C702 B.n570 VSUBS 0.008764f
C703 B.n571 VSUBS 0.008764f
C704 B.n572 VSUBS 0.008764f
C705 B.n573 VSUBS 0.008764f
C706 B.n574 VSUBS 0.008764f
C707 B.n575 VSUBS 0.008764f
C708 B.n576 VSUBS 0.008764f
C709 B.n577 VSUBS 0.008764f
C710 B.n578 VSUBS 0.021702f
C711 B.n579 VSUBS 0.020314f
C712 B.n580 VSUBS 0.021313f
C713 B.n581 VSUBS 0.008764f
C714 B.n582 VSUBS 0.008764f
C715 B.n583 VSUBS 0.008764f
C716 B.n584 VSUBS 0.008764f
C717 B.n585 VSUBS 0.008764f
C718 B.n586 VSUBS 0.008764f
C719 B.n587 VSUBS 0.008764f
C720 B.n588 VSUBS 0.008764f
C721 B.n589 VSUBS 0.008764f
C722 B.n590 VSUBS 0.008764f
C723 B.n591 VSUBS 0.008764f
C724 B.n592 VSUBS 0.008764f
C725 B.n593 VSUBS 0.008764f
C726 B.n594 VSUBS 0.008764f
C727 B.n595 VSUBS 0.008764f
C728 B.n596 VSUBS 0.008764f
C729 B.n597 VSUBS 0.008764f
C730 B.n598 VSUBS 0.008764f
C731 B.n599 VSUBS 0.008764f
C732 B.n600 VSUBS 0.008764f
C733 B.n601 VSUBS 0.008764f
C734 B.n602 VSUBS 0.008764f
C735 B.n603 VSUBS 0.008764f
C736 B.n604 VSUBS 0.008764f
C737 B.n605 VSUBS 0.008764f
C738 B.n606 VSUBS 0.008764f
C739 B.n607 VSUBS 0.008764f
C740 B.n608 VSUBS 0.008764f
C741 B.n609 VSUBS 0.008764f
C742 B.n610 VSUBS 0.008764f
C743 B.n611 VSUBS 0.008764f
C744 B.n612 VSUBS 0.008764f
C745 B.n613 VSUBS 0.008764f
C746 B.n614 VSUBS 0.008764f
C747 B.n615 VSUBS 0.008764f
C748 B.n616 VSUBS 0.008764f
C749 B.n617 VSUBS 0.008764f
C750 B.n618 VSUBS 0.008764f
C751 B.n619 VSUBS 0.006058f
C752 B.n620 VSUBS 0.020306f
C753 B.n621 VSUBS 0.007089f
C754 B.n622 VSUBS 0.008764f
C755 B.n623 VSUBS 0.008764f
C756 B.n624 VSUBS 0.008764f
C757 B.n625 VSUBS 0.008764f
C758 B.n626 VSUBS 0.008764f
C759 B.n627 VSUBS 0.008764f
C760 B.n628 VSUBS 0.008764f
C761 B.n629 VSUBS 0.008764f
C762 B.n630 VSUBS 0.008764f
C763 B.n631 VSUBS 0.008764f
C764 B.n632 VSUBS 0.008764f
C765 B.n633 VSUBS 0.007089f
C766 B.n634 VSUBS 0.020306f
C767 B.n635 VSUBS 0.006058f
C768 B.n636 VSUBS 0.008764f
C769 B.n637 VSUBS 0.008764f
C770 B.n638 VSUBS 0.008764f
C771 B.n639 VSUBS 0.008764f
C772 B.n640 VSUBS 0.008764f
C773 B.n641 VSUBS 0.008764f
C774 B.n642 VSUBS 0.008764f
C775 B.n643 VSUBS 0.008764f
C776 B.n644 VSUBS 0.008764f
C777 B.n645 VSUBS 0.008764f
C778 B.n646 VSUBS 0.008764f
C779 B.n647 VSUBS 0.008764f
C780 B.n648 VSUBS 0.008764f
C781 B.n649 VSUBS 0.008764f
C782 B.n650 VSUBS 0.008764f
C783 B.n651 VSUBS 0.008764f
C784 B.n652 VSUBS 0.008764f
C785 B.n653 VSUBS 0.008764f
C786 B.n654 VSUBS 0.008764f
C787 B.n655 VSUBS 0.008764f
C788 B.n656 VSUBS 0.008764f
C789 B.n657 VSUBS 0.008764f
C790 B.n658 VSUBS 0.008764f
C791 B.n659 VSUBS 0.008764f
C792 B.n660 VSUBS 0.008764f
C793 B.n661 VSUBS 0.008764f
C794 B.n662 VSUBS 0.008764f
C795 B.n663 VSUBS 0.008764f
C796 B.n664 VSUBS 0.008764f
C797 B.n665 VSUBS 0.008764f
C798 B.n666 VSUBS 0.008764f
C799 B.n667 VSUBS 0.008764f
C800 B.n668 VSUBS 0.008764f
C801 B.n669 VSUBS 0.008764f
C802 B.n670 VSUBS 0.008764f
C803 B.n671 VSUBS 0.008764f
C804 B.n672 VSUBS 0.008764f
C805 B.n673 VSUBS 0.008764f
C806 B.n674 VSUBS 0.021313f
C807 B.n675 VSUBS 0.021313f
C808 B.n676 VSUBS 0.020704f
C809 B.n677 VSUBS 0.008764f
C810 B.n678 VSUBS 0.008764f
C811 B.n679 VSUBS 0.008764f
C812 B.n680 VSUBS 0.008764f
C813 B.n681 VSUBS 0.008764f
C814 B.n682 VSUBS 0.008764f
C815 B.n683 VSUBS 0.008764f
C816 B.n684 VSUBS 0.008764f
C817 B.n685 VSUBS 0.008764f
C818 B.n686 VSUBS 0.008764f
C819 B.n687 VSUBS 0.008764f
C820 B.n688 VSUBS 0.008764f
C821 B.n689 VSUBS 0.008764f
C822 B.n690 VSUBS 0.008764f
C823 B.n691 VSUBS 0.008764f
C824 B.n692 VSUBS 0.008764f
C825 B.n693 VSUBS 0.008764f
C826 B.n694 VSUBS 0.008764f
C827 B.n695 VSUBS 0.008764f
C828 B.n696 VSUBS 0.008764f
C829 B.n697 VSUBS 0.008764f
C830 B.n698 VSUBS 0.008764f
C831 B.n699 VSUBS 0.008764f
C832 B.n700 VSUBS 0.008764f
C833 B.n701 VSUBS 0.008764f
C834 B.n702 VSUBS 0.008764f
C835 B.n703 VSUBS 0.008764f
C836 B.n704 VSUBS 0.008764f
C837 B.n705 VSUBS 0.008764f
C838 B.n706 VSUBS 0.008764f
C839 B.n707 VSUBS 0.008764f
C840 B.n708 VSUBS 0.008764f
C841 B.n709 VSUBS 0.008764f
C842 B.n710 VSUBS 0.008764f
C843 B.n711 VSUBS 0.008764f
C844 B.n712 VSUBS 0.008764f
C845 B.n713 VSUBS 0.008764f
C846 B.n714 VSUBS 0.008764f
C847 B.n715 VSUBS 0.008764f
C848 B.n716 VSUBS 0.008764f
C849 B.n717 VSUBS 0.008764f
C850 B.n718 VSUBS 0.008764f
C851 B.n719 VSUBS 0.008764f
C852 B.n720 VSUBS 0.008764f
C853 B.n721 VSUBS 0.008764f
C854 B.n722 VSUBS 0.008764f
C855 B.n723 VSUBS 0.008764f
C856 B.n724 VSUBS 0.008764f
C857 B.n725 VSUBS 0.008764f
C858 B.n726 VSUBS 0.008764f
C859 B.n727 VSUBS 0.008764f
C860 B.n728 VSUBS 0.008764f
C861 B.n729 VSUBS 0.008764f
C862 B.n730 VSUBS 0.008764f
C863 B.n731 VSUBS 0.008764f
C864 B.n732 VSUBS 0.008764f
C865 B.n733 VSUBS 0.008764f
C866 B.n734 VSUBS 0.008764f
C867 B.n735 VSUBS 0.008764f
C868 B.n736 VSUBS 0.008764f
C869 B.n737 VSUBS 0.008764f
C870 B.n738 VSUBS 0.008764f
C871 B.n739 VSUBS 0.008764f
C872 B.n740 VSUBS 0.008764f
C873 B.n741 VSUBS 0.008764f
C874 B.n742 VSUBS 0.008764f
C875 B.n743 VSUBS 0.008764f
C876 B.n744 VSUBS 0.008764f
C877 B.n745 VSUBS 0.008764f
C878 B.n746 VSUBS 0.008764f
C879 B.n747 VSUBS 0.008764f
C880 B.n748 VSUBS 0.008764f
C881 B.n749 VSUBS 0.008764f
C882 B.n750 VSUBS 0.008764f
C883 B.n751 VSUBS 0.008764f
C884 B.n752 VSUBS 0.008764f
C885 B.n753 VSUBS 0.008764f
C886 B.n754 VSUBS 0.008764f
C887 B.n755 VSUBS 0.008764f
C888 B.n756 VSUBS 0.008764f
C889 B.n757 VSUBS 0.008764f
C890 B.n758 VSUBS 0.008764f
C891 B.n759 VSUBS 0.008764f
C892 B.n760 VSUBS 0.008764f
C893 B.n761 VSUBS 0.008764f
C894 B.n762 VSUBS 0.008764f
C895 B.n763 VSUBS 0.008764f
C896 B.n764 VSUBS 0.008764f
C897 B.n765 VSUBS 0.008764f
C898 B.n766 VSUBS 0.008764f
C899 B.n767 VSUBS 0.008764f
C900 B.n768 VSUBS 0.008764f
C901 B.n769 VSUBS 0.008764f
C902 B.n770 VSUBS 0.008764f
C903 B.n771 VSUBS 0.019845f
C904 VDD1.t0 VSUBS 0.182081f
C905 VDD1.t2 VSUBS 0.182081f
C906 VDD1.n0 VSUBS 1.2729f
C907 VDD1.t4 VSUBS 0.182081f
C908 VDD1.t6 VSUBS 0.182081f
C909 VDD1.n1 VSUBS 1.27128f
C910 VDD1.t1 VSUBS 0.182081f
C911 VDD1.t7 VSUBS 0.182081f
C912 VDD1.n2 VSUBS 1.27128f
C913 VDD1.n3 VSUBS 5.17463f
C914 VDD1.t3 VSUBS 0.182081f
C915 VDD1.t5 VSUBS 0.182081f
C916 VDD1.n4 VSUBS 1.25182f
C917 VDD1.n5 VSUBS 4.08463f
C918 VTAIL.t3 VSUBS 0.162136f
C919 VTAIL.t6 VSUBS 0.162136f
C920 VTAIL.n0 VSUBS 0.993368f
C921 VTAIL.n1 VSUBS 0.893804f
C922 VTAIL.t2 VSUBS 1.35443f
C923 VTAIL.n2 VSUBS 1.01387f
C924 VTAIL.t11 VSUBS 1.35443f
C925 VTAIL.n3 VSUBS 1.01387f
C926 VTAIL.t12 VSUBS 0.162136f
C927 VTAIL.t14 VSUBS 0.162136f
C928 VTAIL.n4 VSUBS 0.993368f
C929 VTAIL.n5 VSUBS 1.19243f
C930 VTAIL.t8 VSUBS 1.35443f
C931 VTAIL.n6 VSUBS 2.24221f
C932 VTAIL.t7 VSUBS 1.35443f
C933 VTAIL.n7 VSUBS 2.24221f
C934 VTAIL.t4 VSUBS 0.162136f
C935 VTAIL.t5 VSUBS 0.162136f
C936 VTAIL.n8 VSUBS 0.993373f
C937 VTAIL.n9 VSUBS 1.19242f
C938 VTAIL.t0 VSUBS 1.35443f
C939 VTAIL.n10 VSUBS 1.01386f
C940 VTAIL.t15 VSUBS 1.35443f
C941 VTAIL.n11 VSUBS 1.01386f
C942 VTAIL.t9 VSUBS 0.162136f
C943 VTAIL.t13 VSUBS 0.162136f
C944 VTAIL.n12 VSUBS 0.993373f
C945 VTAIL.n13 VSUBS 1.19242f
C946 VTAIL.t10 VSUBS 1.35443f
C947 VTAIL.n14 VSUBS 2.24221f
C948 VTAIL.t1 VSUBS 1.35443f
C949 VTAIL.n15 VSUBS 2.23671f
C950 VP.t0 VSUBS 2.19179f
C951 VP.n0 VSUBS 0.943816f
C952 VP.n1 VSUBS 0.034556f
C953 VP.n2 VSUBS 0.028113f
C954 VP.n3 VSUBS 0.034556f
C955 VP.t6 VSUBS 2.19179f
C956 VP.n4 VSUBS 0.798975f
C957 VP.n5 VSUBS 0.034556f
C958 VP.n6 VSUBS 0.050446f
C959 VP.n7 VSUBS 0.034556f
C960 VP.n8 VSUBS 0.039919f
C961 VP.n9 VSUBS 0.034556f
C962 VP.n10 VSUBS 0.028113f
C963 VP.n11 VSUBS 0.034556f
C964 VP.t3 VSUBS 2.19179f
C965 VP.n12 VSUBS 0.943816f
C966 VP.t2 VSUBS 2.19179f
C967 VP.n13 VSUBS 0.943816f
C968 VP.n14 VSUBS 0.034556f
C969 VP.n15 VSUBS 0.028113f
C970 VP.n16 VSUBS 0.034556f
C971 VP.t4 VSUBS 2.19179f
C972 VP.n17 VSUBS 0.798975f
C973 VP.n18 VSUBS 0.034556f
C974 VP.n19 VSUBS 0.050446f
C975 VP.n20 VSUBS 0.034556f
C976 VP.n21 VSUBS 0.039919f
C977 VP.t7 VSUBS 2.61366f
C978 VP.t5 VSUBS 2.19179f
C979 VP.n22 VSUBS 0.908394f
C980 VP.n23 VSUBS 0.866097f
C981 VP.n24 VSUBS 0.408801f
C982 VP.n25 VSUBS 0.034556f
C983 VP.n26 VSUBS 0.064404f
C984 VP.n27 VSUBS 0.064404f
C985 VP.n28 VSUBS 0.050446f
C986 VP.n29 VSUBS 0.034556f
C987 VP.n30 VSUBS 0.034556f
C988 VP.n31 VSUBS 0.034556f
C989 VP.n32 VSUBS 0.064404f
C990 VP.n33 VSUBS 0.064404f
C991 VP.n34 VSUBS 0.039919f
C992 VP.n35 VSUBS 0.034556f
C993 VP.n36 VSUBS 0.034556f
C994 VP.n37 VSUBS 0.057089f
C995 VP.n38 VSUBS 0.064404f
C996 VP.n39 VSUBS 0.067901f
C997 VP.n40 VSUBS 0.034556f
C998 VP.n41 VSUBS 0.034556f
C999 VP.n42 VSUBS 0.034556f
C1000 VP.n43 VSUBS 0.06928f
C1001 VP.n44 VSUBS 0.064404f
C1002 VP.n45 VSUBS 0.054545f
C1003 VP.n46 VSUBS 0.055773f
C1004 VP.n47 VSUBS 2.02362f
C1005 VP.n48 VSUBS 2.04797f
C1006 VP.n49 VSUBS 0.055773f
C1007 VP.n50 VSUBS 0.054545f
C1008 VP.n51 VSUBS 0.064404f
C1009 VP.n52 VSUBS 0.06928f
C1010 VP.n53 VSUBS 0.034556f
C1011 VP.n54 VSUBS 0.034556f
C1012 VP.n55 VSUBS 0.034556f
C1013 VP.n56 VSUBS 0.067901f
C1014 VP.n57 VSUBS 0.064404f
C1015 VP.t1 VSUBS 2.19179f
C1016 VP.n58 VSUBS 0.798975f
C1017 VP.n59 VSUBS 0.057089f
C1018 VP.n60 VSUBS 0.034556f
C1019 VP.n61 VSUBS 0.034556f
C1020 VP.n62 VSUBS 0.034556f
C1021 VP.n63 VSUBS 0.064404f
C1022 VP.n64 VSUBS 0.064404f
C1023 VP.n65 VSUBS 0.050446f
C1024 VP.n66 VSUBS 0.034556f
C1025 VP.n67 VSUBS 0.034556f
C1026 VP.n68 VSUBS 0.034556f
C1027 VP.n69 VSUBS 0.064404f
C1028 VP.n70 VSUBS 0.064404f
C1029 VP.n71 VSUBS 0.039919f
C1030 VP.n72 VSUBS 0.034556f
C1031 VP.n73 VSUBS 0.034556f
C1032 VP.n74 VSUBS 0.057089f
C1033 VP.n75 VSUBS 0.064404f
C1034 VP.n76 VSUBS 0.067901f
C1035 VP.n77 VSUBS 0.034556f
C1036 VP.n78 VSUBS 0.034556f
C1037 VP.n79 VSUBS 0.034556f
C1038 VP.n80 VSUBS 0.06928f
C1039 VP.n81 VSUBS 0.064404f
C1040 VP.n82 VSUBS 0.054545f
C1041 VP.n83 VSUBS 0.055773f
C1042 VP.n84 VSUBS 0.081713f
.ends

